module fake_ariane_1283_n_1963 (n_83, n_8, n_56, n_60, n_170, n_190, n_160, n_64, n_179, n_180, n_119, n_124, n_167, n_90, n_195, n_38, n_47, n_110, n_153, n_18, n_197, n_86, n_75, n_89, n_67, n_176, n_149, n_34, n_158, n_172, n_69, n_95, n_175, n_92, n_143, n_183, n_150, n_98, n_74, n_113, n_114, n_33, n_19, n_40, n_181, n_152, n_120, n_169, n_106, n_12, n_53, n_173, n_111, n_21, n_115, n_133, n_66, n_71, n_24, n_7, n_109, n_96, n_156, n_49, n_20, n_174, n_100, n_17, n_50, n_187, n_132, n_62, n_147, n_51, n_166, n_76, n_103, n_79, n_26, n_3, n_46, n_0, n_84, n_36, n_199, n_91, n_159, n_107, n_189, n_72, n_105, n_128, n_44, n_30, n_82, n_178, n_31, n_42, n_57, n_131, n_70, n_10, n_117, n_139, n_165, n_85, n_130, n_144, n_6, n_48, n_94, n_101, n_4, n_134, n_188, n_185, n_2, n_32, n_37, n_58, n_65, n_123, n_9, n_138, n_112, n_45, n_162, n_11, n_129, n_126, n_137, n_122, n_198, n_148, n_164, n_52, n_157, n_184, n_177, n_135, n_73, n_77, n_171, n_15, n_118, n_93, n_121, n_23, n_61, n_108, n_102, n_182, n_196, n_125, n_22, n_168, n_43, n_1, n_81, n_87, n_13, n_27, n_29, n_41, n_140, n_55, n_191, n_151, n_136, n_192, n_28, n_80, n_146, n_194, n_97, n_154, n_142, n_161, n_14, n_163, n_88, n_186, n_141, n_68, n_116, n_104, n_145, n_78, n_193, n_39, n_59, n_63, n_99, n_16, n_5, n_155, n_127, n_35, n_54, n_25, n_1963);

input n_83;
input n_8;
input n_56;
input n_60;
input n_170;
input n_190;
input n_160;
input n_64;
input n_179;
input n_180;
input n_119;
input n_124;
input n_167;
input n_90;
input n_195;
input n_38;
input n_47;
input n_110;
input n_153;
input n_18;
input n_197;
input n_86;
input n_75;
input n_89;
input n_67;
input n_176;
input n_149;
input n_34;
input n_158;
input n_172;
input n_69;
input n_95;
input n_175;
input n_92;
input n_143;
input n_183;
input n_150;
input n_98;
input n_74;
input n_113;
input n_114;
input n_33;
input n_19;
input n_40;
input n_181;
input n_152;
input n_120;
input n_169;
input n_106;
input n_12;
input n_53;
input n_173;
input n_111;
input n_21;
input n_115;
input n_133;
input n_66;
input n_71;
input n_24;
input n_7;
input n_109;
input n_96;
input n_156;
input n_49;
input n_20;
input n_174;
input n_100;
input n_17;
input n_50;
input n_187;
input n_132;
input n_62;
input n_147;
input n_51;
input n_166;
input n_76;
input n_103;
input n_79;
input n_26;
input n_3;
input n_46;
input n_0;
input n_84;
input n_36;
input n_199;
input n_91;
input n_159;
input n_107;
input n_189;
input n_72;
input n_105;
input n_128;
input n_44;
input n_30;
input n_82;
input n_178;
input n_31;
input n_42;
input n_57;
input n_131;
input n_70;
input n_10;
input n_117;
input n_139;
input n_165;
input n_85;
input n_130;
input n_144;
input n_6;
input n_48;
input n_94;
input n_101;
input n_4;
input n_134;
input n_188;
input n_185;
input n_2;
input n_32;
input n_37;
input n_58;
input n_65;
input n_123;
input n_9;
input n_138;
input n_112;
input n_45;
input n_162;
input n_11;
input n_129;
input n_126;
input n_137;
input n_122;
input n_198;
input n_148;
input n_164;
input n_52;
input n_157;
input n_184;
input n_177;
input n_135;
input n_73;
input n_77;
input n_171;
input n_15;
input n_118;
input n_93;
input n_121;
input n_23;
input n_61;
input n_108;
input n_102;
input n_182;
input n_196;
input n_125;
input n_22;
input n_168;
input n_43;
input n_1;
input n_81;
input n_87;
input n_13;
input n_27;
input n_29;
input n_41;
input n_140;
input n_55;
input n_191;
input n_151;
input n_136;
input n_192;
input n_28;
input n_80;
input n_146;
input n_194;
input n_97;
input n_154;
input n_142;
input n_161;
input n_14;
input n_163;
input n_88;
input n_186;
input n_141;
input n_68;
input n_116;
input n_104;
input n_145;
input n_78;
input n_193;
input n_39;
input n_59;
input n_63;
input n_99;
input n_16;
input n_5;
input n_155;
input n_127;
input n_35;
input n_54;
input n_25;

output n_1963;

wire n_913;
wire n_1681;
wire n_1486;
wire n_1507;
wire n_1938;
wire n_589;
wire n_1174;
wire n_1469;
wire n_691;
wire n_1353;
wire n_1355;
wire n_423;
wire n_1383;
wire n_603;
wire n_373;
wire n_1250;
wire n_1169;
wire n_789;
wire n_850;
wire n_1916;
wire n_610;
wire n_245;
wire n_1713;
wire n_319;
wire n_1436;
wire n_690;
wire n_416;
wire n_1109;
wire n_1430;
wire n_525;
wire n_1463;
wire n_1238;
wire n_1515;
wire n_817;
wire n_1837;
wire n_924;
wire n_781;
wire n_1566;
wire n_717;
wire n_952;
wire n_864;
wire n_1096;
wire n_1379;
wire n_1706;
wire n_524;
wire n_1214;
wire n_634;
wire n_1839;
wire n_1246;
wire n_1138;
wire n_214;
wire n_1853;
wire n_764;
wire n_1503;
wire n_462;
wire n_1196;
wire n_1181;
wire n_410;
wire n_1187;
wire n_1131;
wire n_1225;
wire n_737;
wire n_1298;
wire n_1745;
wire n_1366;
wire n_232;
wire n_568;
wire n_1088;
wire n_1424;
wire n_766;
wire n_1835;
wire n_1457;
wire n_377;
wire n_1682;
wire n_1836;
wire n_520;
wire n_870;
wire n_1453;
wire n_279;
wire n_958;
wire n_945;
wire n_813;
wire n_419;
wire n_270;
wire n_338;
wire n_995;
wire n_285;
wire n_1909;
wire n_1184;
wire n_1961;
wire n_202;
wire n_1535;
wire n_500;
wire n_665;
wire n_754;
wire n_903;
wire n_871;
wire n_1073;
wire n_239;
wire n_402;
wire n_1277;
wire n_1746;
wire n_829;
wire n_1761;
wire n_1062;
wire n_339;
wire n_738;
wire n_1690;
wire n_672;
wire n_740;
wire n_1283;
wire n_1736;
wire n_1018;
wire n_259;
wire n_953;
wire n_1364;
wire n_1888;
wire n_1224;
wire n_1425;
wire n_625;
wire n_557;
wire n_1107;
wire n_1688;
wire n_989;
wire n_242;
wire n_645;
wire n_1944;
wire n_331;
wire n_559;
wire n_267;
wire n_495;
wire n_350;
wire n_381;
wire n_795;
wire n_721;
wire n_1084;
wire n_1718;
wire n_1276;
wire n_1936;
wire n_200;
wire n_1428;
wire n_1284;
wire n_1241;
wire n_821;
wire n_561;
wire n_770;
wire n_1514;
wire n_1528;
wire n_507;
wire n_486;
wire n_901;
wire n_569;
wire n_1145;
wire n_971;
wire n_787;
wire n_1650;
wire n_1519;
wire n_1195;
wire n_1522;
wire n_518;
wire n_1207;
wire n_222;
wire n_786;
wire n_1404;
wire n_868;
wire n_1847;
wire n_1542;
wire n_1314;
wire n_1512;
wire n_1539;
wire n_884;
wire n_1851;
wire n_1415;
wire n_1034;
wire n_1652;
wire n_1676;
wire n_1085;
wire n_277;
wire n_1636;
wire n_432;
wire n_293;
wire n_823;
wire n_1900;
wire n_620;
wire n_1074;
wire n_859;
wire n_1765;
wire n_1889;
wire n_587;
wire n_693;
wire n_863;
wire n_303;
wire n_1254;
wire n_929;
wire n_352;
wire n_206;
wire n_899;
wire n_1703;
wire n_611;
wire n_1295;
wire n_1850;
wire n_365;
wire n_238;
wire n_1013;
wire n_1495;
wire n_1637;
wire n_334;
wire n_661;
wire n_1751;
wire n_300;
wire n_533;
wire n_1917;
wire n_1924;
wire n_438;
wire n_1560;
wire n_1654;
wire n_1548;
wire n_1811;
wire n_440;
wire n_273;
wire n_1396;
wire n_1230;
wire n_612;
wire n_333;
wire n_1840;
wire n_376;
wire n_512;
wire n_1597;
wire n_1771;
wire n_1544;
wire n_579;
wire n_844;
wire n_1012;
wire n_1267;
wire n_1354;
wire n_1790;
wire n_1213;
wire n_237;
wire n_780;
wire n_1918;
wire n_1021;
wire n_1443;
wire n_491;
wire n_1465;
wire n_1949;
wire n_1595;
wire n_1142;
wire n_1140;
wire n_705;
wire n_570;
wire n_260;
wire n_942;
wire n_1437;
wire n_1378;
wire n_461;
wire n_1121;
wire n_1416;
wire n_209;
wire n_490;
wire n_1461;
wire n_1391;
wire n_1947;
wire n_225;
wire n_1599;
wire n_1876;
wire n_1006;
wire n_1830;
wire n_575;
wire n_546;
wire n_503;
wire n_1112;
wire n_700;
wire n_1159;
wire n_772;
wire n_1216;
wire n_1245;
wire n_1669;
wire n_1675;
wire n_676;
wire n_1838;
wire n_1594;
wire n_680;
wire n_1935;
wire n_287;
wire n_1716;
wire n_302;
wire n_1872;
wire n_380;
wire n_1585;
wire n_1432;
wire n_249;
wire n_1108;
wire n_355;
wire n_212;
wire n_444;
wire n_851;
wire n_1590;
wire n_1351;
wire n_1274;
wire n_257;
wire n_652;
wire n_1819;
wire n_475;
wire n_947;
wire n_930;
wire n_1260;
wire n_1179;
wire n_468;
wire n_696;
wire n_1442;
wire n_482;
wire n_798;
wire n_577;
wire n_1833;
wire n_407;
wire n_1691;
wire n_916;
wire n_1386;
wire n_912;
wire n_1884;
wire n_460;
wire n_1555;
wire n_1842;
wire n_366;
wire n_762;
wire n_1253;
wire n_1468;
wire n_1661;
wire n_555;
wire n_804;
wire n_1656;
wire n_1382;
wire n_966;
wire n_992;
wire n_955;
wire n_1182;
wire n_794;
wire n_1692;
wire n_1562;
wire n_514;
wire n_418;
wire n_1376;
wire n_513;
wire n_288;
wire n_1292;
wire n_1178;
wire n_1435;
wire n_1750;
wire n_1026;
wire n_1506;
wire n_1610;
wire n_306;
wire n_203;
wire n_436;
wire n_324;
wire n_669;
wire n_931;
wire n_1491;
wire n_619;
wire n_437;
wire n_967;
wire n_274;
wire n_337;
wire n_1083;
wire n_1418;
wire n_746;
wire n_1357;
wire n_292;
wire n_1079;
wire n_1787;
wire n_1389;
wire n_615;
wire n_1139;
wire n_517;
wire n_1312;
wire n_1717;
wire n_1812;
wire n_824;
wire n_428;
wire n_892;
wire n_1880;
wire n_959;
wire n_1399;
wire n_1101;
wire n_1567;
wire n_1343;
wire n_563;
wire n_1855;
wire n_990;
wire n_1623;
wire n_1903;
wire n_867;
wire n_1226;
wire n_944;
wire n_749;
wire n_1932;
wire n_1780;
wire n_1920;
wire n_815;
wire n_542;
wire n_1340;
wire n_470;
wire n_1240;
wire n_1087;
wire n_632;
wire n_477;
wire n_650;
wire n_425;
wire n_1433;
wire n_1911;
wire n_1825;
wire n_1908;
wire n_1155;
wire n_1071;
wire n_712;
wire n_976;
wire n_909;
wire n_1392;
wire n_767;
wire n_1832;
wire n_1841;
wire n_1680;
wire n_964;
wire n_1627;
wire n_382;
wire n_489;
wire n_251;
wire n_974;
wire n_506;
wire n_1731;
wire n_799;
wire n_1147;
wire n_397;
wire n_471;
wire n_351;
wire n_965;
wire n_1914;
wire n_934;
wire n_1447;
wire n_1220;
wire n_356;
wire n_698;
wire n_1674;
wire n_307;
wire n_1209;
wire n_1020;
wire n_1563;
wire n_646;
wire n_1633;
wire n_404;
wire n_1913;
wire n_1058;
wire n_347;
wire n_1042;
wire n_1234;
wire n_479;
wire n_1578;
wire n_1455;
wire n_299;
wire n_836;
wire n_1279;
wire n_564;
wire n_205;
wire n_1029;
wire n_1247;
wire n_760;
wire n_522;
wire n_1568;
wire n_1483;
wire n_1363;
wire n_367;
wire n_1111;
wire n_970;
wire n_1689;
wire n_713;
wire n_1255;
wire n_1646;
wire n_598;
wire n_345;
wire n_1237;
wire n_927;
wire n_261;
wire n_1095;
wire n_1728;
wire n_370;
wire n_706;
wire n_286;
wire n_1401;
wire n_1419;
wire n_1531;
wire n_776;
wire n_424;
wire n_1933;
wire n_1651;
wire n_1387;
wire n_466;
wire n_1263;
wire n_346;
wire n_1817;
wire n_348;
wire n_552;
wire n_670;
wire n_1826;
wire n_379;
wire n_264;
wire n_441;
wire n_1951;
wire n_1032;
wire n_1217;
wire n_1496;
wire n_637;
wire n_1592;
wire n_327;
wire n_1259;
wire n_1177;
wire n_1231;
wire n_980;
wire n_1618;
wire n_1869;
wire n_1743;
wire n_905;
wire n_207;
wire n_720;
wire n_926;
wire n_1943;
wire n_1802;
wire n_1163;
wire n_1795;
wire n_1384;
wire n_1868;
wire n_1501;
wire n_1173;
wire n_1068;
wire n_1198;
wire n_1570;
wire n_487;
wire n_1518;
wire n_1456;
wire n_1879;
wire n_1886;
wire n_1648;
wire n_1413;
wire n_855;
wire n_808;
wire n_1365;
wire n_553;
wire n_1439;
wire n_814;
wire n_578;
wire n_1665;
wire n_1287;
wire n_405;
wire n_1611;
wire n_320;
wire n_1414;
wire n_1134;
wire n_1484;
wire n_1901;
wire n_647;
wire n_1423;
wire n_481;
wire n_600;
wire n_1053;
wire n_1609;
wire n_1939;
wire n_1906;
wire n_529;
wire n_1899;
wire n_502;
wire n_218;
wire n_1467;
wire n_247;
wire n_1828;
wire n_1798;
wire n_1304;
wire n_1608;
wire n_1744;
wire n_1105;
wire n_547;
wire n_439;
wire n_604;
wire n_677;
wire n_478;
wire n_703;
wire n_1349;
wire n_1709;
wire n_1061;
wire n_326;
wire n_681;
wire n_227;
wire n_874;
wire n_1278;
wire n_707;
wire n_983;
wire n_590;
wire n_699;
wire n_727;
wire n_301;
wire n_1726;
wire n_1945;
wire n_545;
wire n_1015;
wire n_1377;
wire n_1162;
wire n_536;
wire n_1614;
wire n_325;
wire n_1740;
wire n_1602;
wire n_688;
wire n_636;
wire n_427;
wire n_1098;
wire n_1490;
wire n_442;
wire n_777;
wire n_1553;
wire n_1080;
wire n_920;
wire n_1760;
wire n_1086;
wire n_1092;
wire n_986;
wire n_1104;
wire n_729;
wire n_887;
wire n_1122;
wire n_1205;
wire n_1408;
wire n_1693;
wire n_1132;
wire n_390;
wire n_1156;
wire n_501;
wire n_314;
wire n_1823;
wire n_1120;
wire n_1202;
wire n_627;
wire n_1188;
wire n_1498;
wire n_1371;
wire n_233;
wire n_957;
wire n_388;
wire n_1402;
wire n_1242;
wire n_1607;
wire n_1489;
wire n_1218;
wire n_321;
wire n_221;
wire n_1586;
wire n_861;
wire n_1543;
wire n_1431;
wire n_877;
wire n_1119;
wire n_1863;
wire n_1763;
wire n_1666;
wire n_1500;
wire n_616;
wire n_1055;
wire n_1395;
wire n_1346;
wire n_1189;
wire n_1089;
wire n_281;
wire n_1859;
wire n_262;
wire n_1502;
wire n_1523;
wire n_1478;
wire n_1883;
wire n_735;
wire n_297;
wire n_1005;
wire n_527;
wire n_1294;
wire n_1667;
wire n_845;
wire n_888;
wire n_1649;
wire n_1677;
wire n_1927;
wire n_1297;
wire n_551;
wire n_417;
wire n_1708;
wire n_343;
wire n_1222;
wire n_1844;
wire n_582;
wire n_1957;
wire n_1953;
wire n_755;
wire n_1097;
wire n_1219;
wire n_1711;
wire n_710;
wire n_1919;
wire n_534;
wire n_1791;
wire n_1894;
wire n_1460;
wire n_1239;
wire n_278;
wire n_560;
wire n_890;
wire n_842;
wire n_1898;
wire n_451;
wire n_745;
wire n_1741;
wire n_1572;
wire n_1907;
wire n_1793;
wire n_742;
wire n_1081;
wire n_1373;
wire n_1388;
wire n_1266;
wire n_1540;
wire n_1719;
wire n_769;
wire n_1797;
wire n_1753;
wire n_1372;
wire n_476;
wire n_832;
wire n_535;
wire n_744;
wire n_1895;
wire n_982;
wire n_1800;
wire n_915;
wire n_215;
wire n_1075;
wire n_454;
wire n_298;
wire n_1331;
wire n_1890;
wire n_1529;
wire n_1227;
wire n_655;
wire n_1734;
wire n_1860;
wire n_403;
wire n_1007;
wire n_1580;
wire n_1319;
wire n_657;
wire n_837;
wire n_812;
wire n_606;
wire n_951;
wire n_862;
wire n_1700;
wire n_659;
wire n_1332;
wire n_509;
wire n_1854;
wire n_666;
wire n_1747;
wire n_430;
wire n_1206;
wire n_1729;
wire n_722;
wire n_1508;
wire n_1532;
wire n_1171;
wire n_1030;
wire n_785;
wire n_1309;
wire n_999;
wire n_1766;
wire n_1338;
wire n_1342;
wire n_456;
wire n_1867;
wire n_852;
wire n_1394;
wire n_704;
wire n_1060;
wire n_1044;
wire n_1714;
wire n_521;
wire n_873;
wire n_1301;
wire n_1748;
wire n_1243;
wire n_1400;
wire n_342;
wire n_1466;
wire n_1527;
wire n_1513;
wire n_358;
wire n_1783;
wire n_608;
wire n_1538;
wire n_1037;
wire n_1329;
wire n_317;
wire n_1545;
wire n_1257;
wire n_1480;
wire n_1954;
wire n_1668;
wire n_1878;
wire n_1605;
wire n_1078;
wire n_266;
wire n_1897;
wire n_1161;
wire n_811;
wire n_624;
wire n_876;
wire n_791;
wire n_618;
wire n_1191;
wire n_736;
wire n_1025;
wire n_1215;
wire n_241;
wire n_1449;
wire n_687;
wire n_797;
wire n_1786;
wire n_480;
wire n_1327;
wire n_1475;
wire n_642;
wire n_211;
wire n_1804;
wire n_408;
wire n_1406;
wire n_595;
wire n_1405;
wire n_602;
wire n_1757;
wire n_592;
wire n_1499;
wire n_854;
wire n_1318;
wire n_393;
wire n_1632;
wire n_1769;
wire n_474;
wire n_1929;
wire n_1950;
wire n_805;
wire n_295;
wire n_1658;
wire n_1072;
wire n_695;
wire n_1526;
wire n_1305;
wire n_730;
wire n_386;
wire n_1596;
wire n_1281;
wire n_516;
wire n_1137;
wire n_1873;
wire n_1258;
wire n_640;
wire n_463;
wire n_1524;
wire n_1476;
wire n_1733;
wire n_1856;
wire n_943;
wire n_1118;
wire n_678;
wire n_651;
wire n_1874;
wire n_1293;
wire n_961;
wire n_469;
wire n_1046;
wire n_1807;
wire n_726;
wire n_1123;
wire n_1657;
wire n_878;
wire n_1784;
wire n_771;
wire n_1321;
wire n_752;
wire n_1488;
wire n_985;
wire n_421;
wire n_1330;
wire n_906;
wire n_1180;
wire n_1697;
wire n_283;
wire n_806;
wire n_1350;
wire n_1556;
wire n_649;
wire n_1561;
wire n_374;
wire n_1352;
wire n_1824;
wire n_643;
wire n_1492;
wire n_226;
wire n_1441;
wire n_1822;
wire n_682;
wire n_1616;
wire n_819;
wire n_586;
wire n_1324;
wire n_1429;
wire n_1778;
wire n_1776;
wire n_686;
wire n_605;
wire n_1154;
wire n_584;
wire n_1557;
wire n_1759;
wire n_1829;
wire n_1130;
wire n_1450;
wire n_349;
wire n_756;
wire n_1016;
wire n_1149;
wire n_1505;
wire n_979;
wire n_1642;
wire n_1815;
wire n_897;
wire n_949;
wire n_1493;
wire n_515;
wire n_807;
wire n_891;
wire n_885;
wire n_1659;
wire n_1864;
wire n_1887;
wire n_1208;
wire n_396;
wire n_802;
wire n_1151;
wire n_554;
wire n_960;
wire n_1256;
wire n_714;
wire n_790;
wire n_354;
wire n_725;
wire n_1577;
wire n_1448;
wire n_1009;
wire n_230;
wire n_1133;
wire n_883;
wire n_473;
wire n_1852;
wire n_801;
wire n_1286;
wire n_818;
wire n_1685;
wire n_779;
wire n_594;
wire n_1877;
wire n_1397;
wire n_1052;
wire n_272;
wire n_1333;
wire n_1306;
wire n_1849;
wire n_833;
wire n_1426;
wire n_879;
wire n_1117;
wire n_422;
wire n_1269;
wire n_1303;
wire n_1547;
wire n_1438;
wire n_1541;
wire n_597;
wire n_1047;
wire n_1472;
wire n_1593;
wire n_1050;
wire n_566;
wire n_1201;
wire n_1288;
wire n_858;
wire n_1185;
wire n_335;
wire n_1035;
wire n_1143;
wire n_344;
wire n_426;
wire n_433;
wire n_398;
wire n_210;
wire n_1090;
wire n_1367;
wire n_253;
wire n_928;
wire n_1153;
wire n_271;
wire n_465;
wire n_825;
wire n_1103;
wire n_732;
wire n_1565;
wire n_1192;
wire n_224;
wire n_894;
wire n_1380;
wire n_1624;
wire n_1801;
wire n_420;
wire n_1291;
wire n_562;
wire n_748;
wire n_510;
wire n_1045;
wire n_256;
wire n_1160;
wire n_1882;
wire n_1023;
wire n_1881;
wire n_988;
wire n_330;
wire n_914;
wire n_400;
wire n_689;
wire n_1116;
wire n_282;
wire n_328;
wire n_368;
wire n_1958;
wire n_467;
wire n_1511;
wire n_1422;
wire n_644;
wire n_1197;
wire n_276;
wire n_497;
wire n_1165;
wire n_1641;
wire n_538;
wire n_1517;
wire n_576;
wire n_843;
wire n_511;
wire n_455;
wire n_429;
wire n_588;
wire n_638;
wire n_1307;
wire n_1128;
wire n_1671;
wire n_1417;
wire n_1048;
wire n_775;
wire n_667;
wire n_1049;
wire n_869;
wire n_846;
wire n_1398;
wire n_1921;
wire n_1356;
wire n_1341;
wire n_1504;
wire n_1955;
wire n_1773;
wire n_1440;
wire n_1370;
wire n_1603;
wire n_305;
wire n_312;
wire n_728;
wire n_413;
wire n_715;
wire n_889;
wire n_1066;
wire n_1549;
wire n_935;
wire n_685;
wire n_911;
wire n_361;
wire n_623;
wire n_1712;
wire n_1403;
wire n_1065;
wire n_453;
wire n_1534;
wire n_1948;
wire n_810;
wire n_1290;
wire n_1959;
wire n_617;
wire n_543;
wire n_1362;
wire n_1559;
wire n_236;
wire n_601;
wire n_683;
wire n_565;
wire n_628;
wire n_1300;
wire n_1960;
wire n_743;
wire n_1194;
wire n_1647;
wire n_1546;
wire n_1420;
wire n_907;
wire n_1454;
wire n_660;
wire n_464;
wire n_962;
wire n_941;
wire n_1210;
wire n_847;
wire n_747;
wire n_1622;
wire n_1135;
wire n_918;
wire n_1885;
wire n_639;
wire n_452;
wire n_673;
wire n_1038;
wire n_571;
wire n_414;
wire n_1521;
wire n_1694;
wire n_1940;
wire n_284;
wire n_593;
wire n_1695;
wire n_1164;
wire n_609;
wire n_1193;
wire n_1345;
wire n_613;
wire n_1022;
wire n_1336;
wire n_1033;
wire n_1774;
wire n_409;
wire n_519;
wire n_384;
wire n_1166;
wire n_1056;
wire n_526;
wire n_1767;
wire n_1040;
wire n_674;
wire n_1158;
wire n_316;
wire n_1444;
wire n_1803;
wire n_820;
wire n_1749;
wire n_872;
wire n_1653;
wire n_254;
wire n_1157;
wire n_1584;
wire n_234;
wire n_848;
wire n_1664;
wire n_280;
wire n_629;
wire n_1739;
wire n_1814;
wire n_532;
wire n_1789;
wire n_763;
wire n_540;
wire n_216;
wire n_692;
wire n_1857;
wire n_984;
wire n_1687;
wire n_223;
wire n_1552;
wire n_750;
wire n_834;
wire n_1612;
wire n_800;
wire n_1816;
wire n_1910;
wire n_1756;
wire n_1606;
wire n_395;
wire n_621;
wire n_1587;
wire n_213;
wire n_1772;
wire n_1014;
wire n_724;
wire n_1427;
wire n_1481;
wire n_493;
wire n_1311;
wire n_1956;
wire n_1589;
wire n_1100;
wire n_585;
wire n_875;
wire n_1617;
wire n_827;
wire n_697;
wire n_622;
wire n_1626;
wire n_1962;
wire n_1335;
wire n_1715;
wire n_296;
wire n_880;
wire n_793;
wire n_1175;
wire n_751;
wire n_1027;
wire n_1070;
wire n_1621;
wire n_739;
wire n_1485;
wire n_1028;
wire n_1221;
wire n_530;
wire n_1785;
wire n_792;
wire n_1262;
wire n_1942;
wire n_580;
wire n_1579;
wire n_494;
wire n_434;
wire n_975;
wire n_229;
wire n_394;
wire n_923;
wire n_1645;
wire n_1124;
wire n_1381;
wire n_1494;
wire n_932;
wire n_1893;
wire n_1183;
wire n_1326;
wire n_1805;
wire n_981;
wire n_1110;
wire n_1758;
wire n_243;
wire n_1407;
wire n_1204;
wire n_1554;
wire n_994;
wire n_1360;
wire n_973;
wire n_268;
wire n_972;
wire n_856;
wire n_1248;
wire n_1176;
wire n_1564;
wire n_1054;
wire n_508;
wire n_1679;
wire n_1952;
wire n_1858;
wire n_353;
wire n_1678;
wire n_1482;
wire n_1361;
wire n_1601;
wire n_1057;
wire n_1834;
wire n_978;
wire n_1011;
wire n_1520;
wire n_1509;
wire n_828;
wire n_322;
wire n_1411;
wire n_1359;
wire n_558;
wire n_1721;
wire n_653;
wire n_1445;
wire n_1317;
wire n_783;
wire n_556;
wire n_1127;
wire n_1536;
wire n_1471;
wire n_1008;
wire n_332;
wire n_581;
wire n_294;
wire n_1024;
wire n_830;
wire n_987;
wire n_936;
wire n_1620;
wire n_1385;
wire n_1525;
wire n_541;
wire n_499;
wire n_1775;
wire n_788;
wire n_908;
wire n_1036;
wire n_341;
wire n_1270;
wire n_1167;
wire n_1272;
wire n_549;
wire n_591;
wire n_969;
wire n_919;
wire n_1663;
wire n_1625;
wire n_1926;
wire n_318;
wire n_1458;
wire n_679;
wire n_244;
wire n_1630;
wire n_220;
wire n_663;
wire n_1720;
wire n_443;
wire n_1412;
wire n_1738;
wire n_1550;
wire n_528;
wire n_1358;
wire n_1200;
wire n_387;
wire n_406;
wire n_826;
wire n_1922;
wire n_1735;
wire n_1788;
wire n_391;
wire n_940;
wire n_1537;
wire n_1077;
wire n_607;
wire n_956;
wire n_445;
wire n_1930;
wire n_765;
wire n_1809;
wire n_1843;
wire n_1904;
wire n_1268;
wire n_385;
wire n_917;
wire n_1271;
wire n_372;
wire n_1530;
wire n_631;
wire n_399;
wire n_1170;
wire n_1261;
wire n_702;
wire n_898;
wire n_857;
wire n_363;
wire n_1067;
wire n_968;
wire n_1235;
wire n_1323;
wire n_1462;
wire n_1937;
wire n_1064;
wire n_633;
wire n_900;
wire n_1446;
wire n_1282;
wire n_1701;
wire n_1093;
wire n_1551;
wire n_1755;
wire n_1285;
wire n_733;
wire n_761;
wire n_731;
wire n_336;
wire n_1813;
wire n_315;
wire n_311;
wire n_1452;
wire n_1573;
wire n_668;
wire n_758;
wire n_1106;
wire n_648;
wire n_784;
wire n_269;
wire n_816;
wire n_1322;
wire n_1473;
wire n_835;
wire n_446;
wire n_1076;
wire n_1348;
wire n_753;
wire n_1770;
wire n_701;
wire n_1003;
wire n_1125;
wire n_1710;
wire n_1865;
wire n_309;
wire n_1344;
wire n_1390;
wire n_401;
wire n_485;
wire n_1792;
wire n_504;
wire n_483;
wire n_435;
wire n_1141;
wire n_1629;
wire n_291;
wire n_1640;
wire n_822;
wire n_1094;
wire n_840;
wire n_1459;
wire n_1510;
wire n_1099;
wire n_839;
wire n_1754;
wire n_759;
wire n_567;
wire n_240;
wire n_369;
wire n_1727;
wire n_1575;
wire n_1848;
wire n_1892;
wire n_1172;
wire n_614;
wire n_1212;
wire n_831;
wire n_778;
wire n_1619;
wire n_323;
wire n_550;
wire n_1315;
wire n_1660;
wire n_1902;
wire n_997;
wire n_635;
wire n_694;
wire n_1643;
wire n_1320;
wire n_1113;
wire n_248;
wire n_1152;
wire n_1845;
wire n_1934;
wire n_921;
wire n_1615;
wire n_1236;
wire n_228;
wire n_1265;
wire n_1576;
wire n_1470;
wire n_671;
wire n_1533;
wire n_1806;
wire n_1409;
wire n_1148;
wire n_1588;
wire n_1684;
wire n_1673;
wire n_1334;
wire n_654;
wire n_1275;
wire n_488;
wire n_904;
wire n_505;
wire n_1696;
wire n_498;
wire n_1875;
wire n_1059;
wire n_684;
wire n_1039;
wire n_539;
wire n_1150;
wire n_977;
wire n_449;
wire n_392;
wire n_1628;
wire n_1289;
wire n_1831;
wire n_1497;
wire n_1866;
wire n_459;
wire n_1136;
wire n_1782;
wire n_458;
wire n_1190;
wire n_1600;
wire n_1144;
wire n_838;
wire n_383;
wire n_1558;
wire n_1941;
wire n_1316;
wire n_950;
wire n_1017;
wire n_711;
wire n_734;
wire n_1915;
wire n_723;
wire n_1393;
wire n_658;
wire n_630;
wire n_1369;
wire n_362;
wire n_310;
wire n_1781;
wire n_709;
wire n_809;
wire n_1686;
wire n_235;
wire n_881;
wire n_1019;
wire n_1477;
wire n_1777;
wire n_662;
wire n_641;
wire n_910;
wire n_290;
wire n_741;
wire n_939;
wire n_1410;
wire n_371;
wire n_217;
wire n_1114;
wire n_1325;
wire n_1742;
wire n_708;
wire n_308;
wire n_1223;
wire n_201;
wire n_1768;
wire n_572;
wire n_1199;
wire n_865;
wire n_1273;
wire n_1041;
wire n_993;
wire n_1862;
wire n_948;
wire n_922;
wire n_1004;
wire n_1810;
wire n_448;
wire n_1347;
wire n_860;
wire n_1043;
wire n_255;
wire n_450;
wire n_1923;
wire n_1764;
wire n_896;
wire n_1737;
wire n_1479;
wire n_1613;
wire n_902;
wire n_1031;
wire n_1723;
wire n_1638;
wire n_853;
wire n_716;
wire n_1571;
wire n_1698;
wire n_1337;
wire n_774;
wire n_1946;
wire n_933;
wire n_1779;
wire n_596;
wire n_954;
wire n_1168;
wire n_1821;
wire n_219;
wire n_1310;
wire n_231;
wire n_656;
wire n_492;
wire n_574;
wire n_252;
wire n_664;
wire n_1591;
wire n_1229;
wire n_1683;
wire n_1896;
wire n_1732;
wire n_415;
wire n_1280;
wire n_544;
wire n_1516;
wire n_1186;
wire n_1705;
wire n_599;
wire n_768;
wire n_1091;
wire n_537;
wire n_1063;
wire n_991;
wire n_389;
wire n_1724;
wire n_1670;
wire n_1707;
wire n_1799;
wire n_1126;
wire n_1846;
wire n_1912;
wire n_938;
wire n_1891;
wire n_1328;
wire n_895;
wire n_304;
wire n_1639;
wire n_583;
wire n_1302;
wire n_1000;
wire n_313;
wire n_626;
wire n_378;
wire n_1581;
wire n_1928;
wire n_946;
wire n_757;
wire n_375;
wire n_1655;
wire n_1818;
wire n_1146;
wire n_1634;
wire n_1203;
wire n_998;
wire n_1699;
wire n_1598;
wire n_472;
wire n_937;
wire n_1474;
wire n_265;
wire n_1583;
wire n_1604;
wire n_208;
wire n_1631;
wire n_1702;
wire n_275;
wire n_1794;
wire n_1375;
wire n_204;
wire n_1232;
wire n_996;
wire n_1211;
wire n_1368;
wire n_963;
wire n_1264;
wire n_1082;
wire n_1725;
wire n_496;
wire n_1827;
wire n_866;
wire n_246;
wire n_925;
wire n_1752;
wire n_1313;
wire n_1001;
wire n_1722;
wire n_1115;
wire n_1339;
wire n_1002;
wire n_1644;
wire n_1051;
wire n_719;
wire n_263;
wire n_1102;
wire n_360;
wire n_1129;
wire n_1252;
wire n_250;
wire n_1464;
wire n_1296;
wire n_773;
wire n_1010;
wire n_882;
wire n_1249;
wire n_803;
wire n_1871;
wire n_718;
wire n_329;
wire n_1434;
wire n_340;
wire n_1905;
wire n_1569;
wire n_548;
wire n_289;
wire n_523;
wire n_1662;
wire n_457;
wire n_1299;
wire n_1870;
wire n_1925;
wire n_782;
wire n_364;
wire n_258;
wire n_431;
wire n_1861;
wire n_1228;
wire n_1931;
wire n_1244;
wire n_1796;
wire n_411;
wire n_484;
wire n_849;
wire n_1820;
wire n_357;
wire n_412;
wire n_1251;
wire n_447;
wire n_1421;
wire n_1762;
wire n_1233;
wire n_1808;
wire n_1574;
wire n_1672;
wire n_1635;
wire n_1704;
wire n_893;
wire n_1582;
wire n_841;
wire n_886;
wire n_1069;
wire n_359;
wire n_1308;
wire n_573;
wire n_796;
wire n_531;
wire n_1730;
wire n_1374;
wire n_1451;
wire n_1487;
wire n_675;

BUFx6f_ASAP7_75t_L g200 ( 
.A(n_71),
.Y(n_200)
);

INVx1_ASAP7_75t_SL g201 ( 
.A(n_129),
.Y(n_201)
);

CKINVDCx5p33_ASAP7_75t_R g202 ( 
.A(n_78),
.Y(n_202)
);

CKINVDCx5p33_ASAP7_75t_R g203 ( 
.A(n_167),
.Y(n_203)
);

CKINVDCx5p33_ASAP7_75t_R g204 ( 
.A(n_182),
.Y(n_204)
);

CKINVDCx5p33_ASAP7_75t_R g205 ( 
.A(n_175),
.Y(n_205)
);

CKINVDCx5p33_ASAP7_75t_R g206 ( 
.A(n_65),
.Y(n_206)
);

CKINVDCx5p33_ASAP7_75t_R g207 ( 
.A(n_110),
.Y(n_207)
);

HB1xp67_ASAP7_75t_L g208 ( 
.A(n_93),
.Y(n_208)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_7),
.Y(n_209)
);

CKINVDCx5p33_ASAP7_75t_R g210 ( 
.A(n_166),
.Y(n_210)
);

BUFx6f_ASAP7_75t_L g211 ( 
.A(n_171),
.Y(n_211)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_176),
.Y(n_212)
);

CKINVDCx5p33_ASAP7_75t_R g213 ( 
.A(n_194),
.Y(n_213)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_179),
.Y(n_214)
);

CKINVDCx5p33_ASAP7_75t_R g215 ( 
.A(n_99),
.Y(n_215)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_139),
.Y(n_216)
);

INVx2_ASAP7_75t_L g217 ( 
.A(n_10),
.Y(n_217)
);

HB1xp67_ASAP7_75t_L g218 ( 
.A(n_149),
.Y(n_218)
);

CKINVDCx5p33_ASAP7_75t_R g219 ( 
.A(n_148),
.Y(n_219)
);

CKINVDCx5p33_ASAP7_75t_R g220 ( 
.A(n_186),
.Y(n_220)
);

CKINVDCx5p33_ASAP7_75t_R g221 ( 
.A(n_124),
.Y(n_221)
);

CKINVDCx5p33_ASAP7_75t_R g222 ( 
.A(n_188),
.Y(n_222)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_67),
.Y(n_223)
);

CKINVDCx5p33_ASAP7_75t_R g224 ( 
.A(n_191),
.Y(n_224)
);

CKINVDCx5p33_ASAP7_75t_R g225 ( 
.A(n_162),
.Y(n_225)
);

CKINVDCx5p33_ASAP7_75t_R g226 ( 
.A(n_79),
.Y(n_226)
);

INVx2_ASAP7_75t_L g227 ( 
.A(n_146),
.Y(n_227)
);

INVx1_ASAP7_75t_SL g228 ( 
.A(n_199),
.Y(n_228)
);

CKINVDCx5p33_ASAP7_75t_R g229 ( 
.A(n_31),
.Y(n_229)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_16),
.Y(n_230)
);

CKINVDCx5p33_ASAP7_75t_R g231 ( 
.A(n_43),
.Y(n_231)
);

CKINVDCx5p33_ASAP7_75t_R g232 ( 
.A(n_101),
.Y(n_232)
);

CKINVDCx5p33_ASAP7_75t_R g233 ( 
.A(n_3),
.Y(n_233)
);

CKINVDCx20_ASAP7_75t_R g234 ( 
.A(n_31),
.Y(n_234)
);

CKINVDCx5p33_ASAP7_75t_R g235 ( 
.A(n_61),
.Y(n_235)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_100),
.Y(n_236)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_75),
.Y(n_237)
);

BUFx3_ASAP7_75t_L g238 ( 
.A(n_135),
.Y(n_238)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_54),
.Y(n_239)
);

INVx2_ASAP7_75t_SL g240 ( 
.A(n_119),
.Y(n_240)
);

CKINVDCx5p33_ASAP7_75t_R g241 ( 
.A(n_80),
.Y(n_241)
);

BUFx10_ASAP7_75t_L g242 ( 
.A(n_154),
.Y(n_242)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_52),
.Y(n_243)
);

CKINVDCx5p33_ASAP7_75t_R g244 ( 
.A(n_116),
.Y(n_244)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_134),
.Y(n_245)
);

CKINVDCx5p33_ASAP7_75t_R g246 ( 
.A(n_4),
.Y(n_246)
);

CKINVDCx5p33_ASAP7_75t_R g247 ( 
.A(n_152),
.Y(n_247)
);

INVx2_ASAP7_75t_L g248 ( 
.A(n_158),
.Y(n_248)
);

BUFx6f_ASAP7_75t_L g249 ( 
.A(n_69),
.Y(n_249)
);

CKINVDCx5p33_ASAP7_75t_R g250 ( 
.A(n_133),
.Y(n_250)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_64),
.Y(n_251)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_56),
.Y(n_252)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_98),
.Y(n_253)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_72),
.Y(n_254)
);

CKINVDCx5p33_ASAP7_75t_R g255 ( 
.A(n_26),
.Y(n_255)
);

CKINVDCx5p33_ASAP7_75t_R g256 ( 
.A(n_12),
.Y(n_256)
);

CKINVDCx5p33_ASAP7_75t_R g257 ( 
.A(n_57),
.Y(n_257)
);

CKINVDCx5p33_ASAP7_75t_R g258 ( 
.A(n_1),
.Y(n_258)
);

CKINVDCx20_ASAP7_75t_R g259 ( 
.A(n_84),
.Y(n_259)
);

BUFx3_ASAP7_75t_L g260 ( 
.A(n_82),
.Y(n_260)
);

INVxp67_ASAP7_75t_SL g261 ( 
.A(n_170),
.Y(n_261)
);

CKINVDCx20_ASAP7_75t_R g262 ( 
.A(n_121),
.Y(n_262)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_144),
.Y(n_263)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_140),
.Y(n_264)
);

CKINVDCx5p33_ASAP7_75t_R g265 ( 
.A(n_26),
.Y(n_265)
);

BUFx10_ASAP7_75t_L g266 ( 
.A(n_32),
.Y(n_266)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_145),
.Y(n_267)
);

INVx2_ASAP7_75t_L g268 ( 
.A(n_181),
.Y(n_268)
);

INVx2_ASAP7_75t_L g269 ( 
.A(n_97),
.Y(n_269)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_21),
.Y(n_270)
);

CKINVDCx5p33_ASAP7_75t_R g271 ( 
.A(n_161),
.Y(n_271)
);

INVx2_ASAP7_75t_L g272 ( 
.A(n_57),
.Y(n_272)
);

CKINVDCx20_ASAP7_75t_R g273 ( 
.A(n_102),
.Y(n_273)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_128),
.Y(n_274)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_151),
.Y(n_275)
);

CKINVDCx5p33_ASAP7_75t_R g276 ( 
.A(n_147),
.Y(n_276)
);

CKINVDCx5p33_ASAP7_75t_R g277 ( 
.A(n_59),
.Y(n_277)
);

CKINVDCx5p33_ASAP7_75t_R g278 ( 
.A(n_49),
.Y(n_278)
);

BUFx10_ASAP7_75t_L g279 ( 
.A(n_174),
.Y(n_279)
);

CKINVDCx5p33_ASAP7_75t_R g280 ( 
.A(n_153),
.Y(n_280)
);

CKINVDCx5p33_ASAP7_75t_R g281 ( 
.A(n_3),
.Y(n_281)
);

CKINVDCx5p33_ASAP7_75t_R g282 ( 
.A(n_86),
.Y(n_282)
);

CKINVDCx5p33_ASAP7_75t_R g283 ( 
.A(n_160),
.Y(n_283)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_39),
.Y(n_284)
);

CKINVDCx5p33_ASAP7_75t_R g285 ( 
.A(n_6),
.Y(n_285)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_45),
.Y(n_286)
);

CKINVDCx5p33_ASAP7_75t_R g287 ( 
.A(n_185),
.Y(n_287)
);

CKINVDCx20_ASAP7_75t_R g288 ( 
.A(n_163),
.Y(n_288)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_90),
.Y(n_289)
);

CKINVDCx5p33_ASAP7_75t_R g290 ( 
.A(n_50),
.Y(n_290)
);

CKINVDCx5p33_ASAP7_75t_R g291 ( 
.A(n_107),
.Y(n_291)
);

INVx1_ASAP7_75t_SL g292 ( 
.A(n_122),
.Y(n_292)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_92),
.Y(n_293)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_156),
.Y(n_294)
);

CKINVDCx5p33_ASAP7_75t_R g295 ( 
.A(n_63),
.Y(n_295)
);

BUFx3_ASAP7_75t_L g296 ( 
.A(n_62),
.Y(n_296)
);

CKINVDCx5p33_ASAP7_75t_R g297 ( 
.A(n_89),
.Y(n_297)
);

CKINVDCx5p33_ASAP7_75t_R g298 ( 
.A(n_106),
.Y(n_298)
);

CKINVDCx5p33_ASAP7_75t_R g299 ( 
.A(n_142),
.Y(n_299)
);

CKINVDCx5p33_ASAP7_75t_R g300 ( 
.A(n_183),
.Y(n_300)
);

CKINVDCx5p33_ASAP7_75t_R g301 ( 
.A(n_16),
.Y(n_301)
);

BUFx2_ASAP7_75t_L g302 ( 
.A(n_187),
.Y(n_302)
);

CKINVDCx5p33_ASAP7_75t_R g303 ( 
.A(n_42),
.Y(n_303)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_29),
.Y(n_304)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_68),
.Y(n_305)
);

HB1xp67_ASAP7_75t_L g306 ( 
.A(n_195),
.Y(n_306)
);

CKINVDCx5p33_ASAP7_75t_R g307 ( 
.A(n_52),
.Y(n_307)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_190),
.Y(n_308)
);

CKINVDCx5p33_ASAP7_75t_R g309 ( 
.A(n_61),
.Y(n_309)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_59),
.Y(n_310)
);

CKINVDCx5p33_ASAP7_75t_R g311 ( 
.A(n_192),
.Y(n_311)
);

BUFx2_ASAP7_75t_L g312 ( 
.A(n_13),
.Y(n_312)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_35),
.Y(n_313)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_132),
.Y(n_314)
);

INVx2_ASAP7_75t_L g315 ( 
.A(n_74),
.Y(n_315)
);

CKINVDCx5p33_ASAP7_75t_R g316 ( 
.A(n_62),
.Y(n_316)
);

CKINVDCx5p33_ASAP7_75t_R g317 ( 
.A(n_96),
.Y(n_317)
);

CKINVDCx5p33_ASAP7_75t_R g318 ( 
.A(n_46),
.Y(n_318)
);

CKINVDCx5p33_ASAP7_75t_R g319 ( 
.A(n_125),
.Y(n_319)
);

CKINVDCx5p33_ASAP7_75t_R g320 ( 
.A(n_168),
.Y(n_320)
);

BUFx10_ASAP7_75t_L g321 ( 
.A(n_51),
.Y(n_321)
);

CKINVDCx5p33_ASAP7_75t_R g322 ( 
.A(n_196),
.Y(n_322)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_85),
.Y(n_323)
);

CKINVDCx5p33_ASAP7_75t_R g324 ( 
.A(n_157),
.Y(n_324)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_83),
.Y(n_325)
);

CKINVDCx5p33_ASAP7_75t_R g326 ( 
.A(n_21),
.Y(n_326)
);

CKINVDCx5p33_ASAP7_75t_R g327 ( 
.A(n_18),
.Y(n_327)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_180),
.Y(n_328)
);

CKINVDCx5p33_ASAP7_75t_R g329 ( 
.A(n_126),
.Y(n_329)
);

BUFx2_ASAP7_75t_L g330 ( 
.A(n_12),
.Y(n_330)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_77),
.Y(n_331)
);

INVx2_ASAP7_75t_SL g332 ( 
.A(n_51),
.Y(n_332)
);

CKINVDCx5p33_ASAP7_75t_R g333 ( 
.A(n_104),
.Y(n_333)
);

CKINVDCx14_ASAP7_75t_R g334 ( 
.A(n_46),
.Y(n_334)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_70),
.Y(n_335)
);

BUFx10_ASAP7_75t_L g336 ( 
.A(n_49),
.Y(n_336)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_66),
.Y(n_337)
);

CKINVDCx5p33_ASAP7_75t_R g338 ( 
.A(n_87),
.Y(n_338)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_164),
.Y(n_339)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_189),
.Y(n_340)
);

BUFx10_ASAP7_75t_L g341 ( 
.A(n_58),
.Y(n_341)
);

CKINVDCx5p33_ASAP7_75t_R g342 ( 
.A(n_136),
.Y(n_342)
);

BUFx2_ASAP7_75t_L g343 ( 
.A(n_193),
.Y(n_343)
);

INVx2_ASAP7_75t_L g344 ( 
.A(n_44),
.Y(n_344)
);

CKINVDCx5p33_ASAP7_75t_R g345 ( 
.A(n_13),
.Y(n_345)
);

CKINVDCx14_ASAP7_75t_R g346 ( 
.A(n_45),
.Y(n_346)
);

CKINVDCx5p33_ASAP7_75t_R g347 ( 
.A(n_143),
.Y(n_347)
);

CKINVDCx5p33_ASAP7_75t_R g348 ( 
.A(n_27),
.Y(n_348)
);

INVx1_ASAP7_75t_L g349 ( 
.A(n_53),
.Y(n_349)
);

INVx2_ASAP7_75t_L g350 ( 
.A(n_172),
.Y(n_350)
);

INVx1_ASAP7_75t_SL g351 ( 
.A(n_118),
.Y(n_351)
);

INVx1_ASAP7_75t_L g352 ( 
.A(n_23),
.Y(n_352)
);

INVx1_ASAP7_75t_SL g353 ( 
.A(n_17),
.Y(n_353)
);

CKINVDCx5p33_ASAP7_75t_R g354 ( 
.A(n_42),
.Y(n_354)
);

INVx1_ASAP7_75t_SL g355 ( 
.A(n_115),
.Y(n_355)
);

INVx1_ASAP7_75t_L g356 ( 
.A(n_30),
.Y(n_356)
);

INVx1_ASAP7_75t_L g357 ( 
.A(n_81),
.Y(n_357)
);

BUFx2_ASAP7_75t_SL g358 ( 
.A(n_197),
.Y(n_358)
);

CKINVDCx5p33_ASAP7_75t_R g359 ( 
.A(n_47),
.Y(n_359)
);

BUFx8_ASAP7_75t_SL g360 ( 
.A(n_159),
.Y(n_360)
);

CKINVDCx5p33_ASAP7_75t_R g361 ( 
.A(n_47),
.Y(n_361)
);

INVx1_ASAP7_75t_L g362 ( 
.A(n_112),
.Y(n_362)
);

INVx2_ASAP7_75t_L g363 ( 
.A(n_58),
.Y(n_363)
);

CKINVDCx5p33_ASAP7_75t_R g364 ( 
.A(n_120),
.Y(n_364)
);

BUFx6f_ASAP7_75t_L g365 ( 
.A(n_23),
.Y(n_365)
);

CKINVDCx5p33_ASAP7_75t_R g366 ( 
.A(n_109),
.Y(n_366)
);

INVx2_ASAP7_75t_L g367 ( 
.A(n_114),
.Y(n_367)
);

CKINVDCx5p33_ASAP7_75t_R g368 ( 
.A(n_137),
.Y(n_368)
);

CKINVDCx5p33_ASAP7_75t_R g369 ( 
.A(n_53),
.Y(n_369)
);

INVx1_ASAP7_75t_L g370 ( 
.A(n_76),
.Y(n_370)
);

INVx1_ASAP7_75t_L g371 ( 
.A(n_36),
.Y(n_371)
);

INVxp67_ASAP7_75t_L g372 ( 
.A(n_103),
.Y(n_372)
);

CKINVDCx5p33_ASAP7_75t_R g373 ( 
.A(n_1),
.Y(n_373)
);

INVx1_ASAP7_75t_L g374 ( 
.A(n_7),
.Y(n_374)
);

CKINVDCx5p33_ASAP7_75t_R g375 ( 
.A(n_0),
.Y(n_375)
);

INVx2_ASAP7_75t_L g376 ( 
.A(n_25),
.Y(n_376)
);

CKINVDCx5p33_ASAP7_75t_R g377 ( 
.A(n_5),
.Y(n_377)
);

INVx1_ASAP7_75t_L g378 ( 
.A(n_108),
.Y(n_378)
);

CKINVDCx5p33_ASAP7_75t_R g379 ( 
.A(n_24),
.Y(n_379)
);

CKINVDCx5p33_ASAP7_75t_R g380 ( 
.A(n_56),
.Y(n_380)
);

INVx1_ASAP7_75t_L g381 ( 
.A(n_105),
.Y(n_381)
);

BUFx3_ASAP7_75t_L g382 ( 
.A(n_127),
.Y(n_382)
);

CKINVDCx5p33_ASAP7_75t_R g383 ( 
.A(n_169),
.Y(n_383)
);

INVx1_ASAP7_75t_L g384 ( 
.A(n_91),
.Y(n_384)
);

CKINVDCx5p33_ASAP7_75t_R g385 ( 
.A(n_41),
.Y(n_385)
);

CKINVDCx5p33_ASAP7_75t_R g386 ( 
.A(n_184),
.Y(n_386)
);

CKINVDCx20_ASAP7_75t_R g387 ( 
.A(n_50),
.Y(n_387)
);

CKINVDCx5p33_ASAP7_75t_R g388 ( 
.A(n_55),
.Y(n_388)
);

CKINVDCx5p33_ASAP7_75t_R g389 ( 
.A(n_60),
.Y(n_389)
);

CKINVDCx20_ASAP7_75t_R g390 ( 
.A(n_4),
.Y(n_390)
);

CKINVDCx5p33_ASAP7_75t_R g391 ( 
.A(n_32),
.Y(n_391)
);

INVx1_ASAP7_75t_L g392 ( 
.A(n_10),
.Y(n_392)
);

INVx1_ASAP7_75t_L g393 ( 
.A(n_15),
.Y(n_393)
);

INVx1_ASAP7_75t_L g394 ( 
.A(n_36),
.Y(n_394)
);

CKINVDCx5p33_ASAP7_75t_R g395 ( 
.A(n_38),
.Y(n_395)
);

INVx2_ASAP7_75t_SL g396 ( 
.A(n_155),
.Y(n_396)
);

CKINVDCx20_ASAP7_75t_R g397 ( 
.A(n_113),
.Y(n_397)
);

INVx1_ASAP7_75t_L g398 ( 
.A(n_296),
.Y(n_398)
);

INVx1_ASAP7_75t_L g399 ( 
.A(n_296),
.Y(n_399)
);

INVx1_ASAP7_75t_L g400 ( 
.A(n_365),
.Y(n_400)
);

INVx1_ASAP7_75t_L g401 ( 
.A(n_365),
.Y(n_401)
);

INVx1_ASAP7_75t_L g402 ( 
.A(n_365),
.Y(n_402)
);

INVx1_ASAP7_75t_L g403 ( 
.A(n_365),
.Y(n_403)
);

INVxp33_ASAP7_75t_L g404 ( 
.A(n_312),
.Y(n_404)
);

INVx1_ASAP7_75t_L g405 ( 
.A(n_365),
.Y(n_405)
);

INVx1_ASAP7_75t_L g406 ( 
.A(n_217),
.Y(n_406)
);

CKINVDCx20_ASAP7_75t_R g407 ( 
.A(n_334),
.Y(n_407)
);

INVx1_ASAP7_75t_L g408 ( 
.A(n_217),
.Y(n_408)
);

CKINVDCx5p33_ASAP7_75t_R g409 ( 
.A(n_360),
.Y(n_409)
);

INVx2_ASAP7_75t_L g410 ( 
.A(n_238),
.Y(n_410)
);

CKINVDCx5p33_ASAP7_75t_R g411 ( 
.A(n_259),
.Y(n_411)
);

INVx1_ASAP7_75t_L g412 ( 
.A(n_272),
.Y(n_412)
);

INVx1_ASAP7_75t_L g413 ( 
.A(n_272),
.Y(n_413)
);

INVx1_ASAP7_75t_L g414 ( 
.A(n_344),
.Y(n_414)
);

CKINVDCx20_ASAP7_75t_R g415 ( 
.A(n_346),
.Y(n_415)
);

INVx1_ASAP7_75t_L g416 ( 
.A(n_344),
.Y(n_416)
);

CKINVDCx5p33_ASAP7_75t_R g417 ( 
.A(n_262),
.Y(n_417)
);

INVx1_ASAP7_75t_L g418 ( 
.A(n_363),
.Y(n_418)
);

INVx1_ASAP7_75t_L g419 ( 
.A(n_363),
.Y(n_419)
);

INVx1_ASAP7_75t_L g420 ( 
.A(n_376),
.Y(n_420)
);

CKINVDCx5p33_ASAP7_75t_R g421 ( 
.A(n_273),
.Y(n_421)
);

CKINVDCx5p33_ASAP7_75t_R g422 ( 
.A(n_288),
.Y(n_422)
);

CKINVDCx20_ASAP7_75t_R g423 ( 
.A(n_397),
.Y(n_423)
);

INVxp67_ASAP7_75t_L g424 ( 
.A(n_330),
.Y(n_424)
);

INVxp33_ASAP7_75t_SL g425 ( 
.A(n_229),
.Y(n_425)
);

INVx1_ASAP7_75t_L g426 ( 
.A(n_376),
.Y(n_426)
);

INVx1_ASAP7_75t_L g427 ( 
.A(n_227),
.Y(n_427)
);

INVx1_ASAP7_75t_L g428 ( 
.A(n_227),
.Y(n_428)
);

INVxp67_ASAP7_75t_L g429 ( 
.A(n_332),
.Y(n_429)
);

INVx1_ASAP7_75t_L g430 ( 
.A(n_248),
.Y(n_430)
);

INVxp33_ASAP7_75t_SL g431 ( 
.A(n_229),
.Y(n_431)
);

CKINVDCx5p33_ASAP7_75t_R g432 ( 
.A(n_255),
.Y(n_432)
);

INVx1_ASAP7_75t_L g433 ( 
.A(n_248),
.Y(n_433)
);

INVx1_ASAP7_75t_L g434 ( 
.A(n_268),
.Y(n_434)
);

CKINVDCx5p33_ASAP7_75t_R g435 ( 
.A(n_256),
.Y(n_435)
);

INVx1_ASAP7_75t_L g436 ( 
.A(n_268),
.Y(n_436)
);

INVxp67_ASAP7_75t_L g437 ( 
.A(n_332),
.Y(n_437)
);

CKINVDCx5p33_ASAP7_75t_R g438 ( 
.A(n_257),
.Y(n_438)
);

INVx1_ASAP7_75t_L g439 ( 
.A(n_269),
.Y(n_439)
);

INVx1_ASAP7_75t_L g440 ( 
.A(n_269),
.Y(n_440)
);

INVx1_ASAP7_75t_L g441 ( 
.A(n_315),
.Y(n_441)
);

CKINVDCx20_ASAP7_75t_R g442 ( 
.A(n_234),
.Y(n_442)
);

CKINVDCx20_ASAP7_75t_R g443 ( 
.A(n_387),
.Y(n_443)
);

BUFx2_ASAP7_75t_L g444 ( 
.A(n_231),
.Y(n_444)
);

INVx1_ASAP7_75t_L g445 ( 
.A(n_209),
.Y(n_445)
);

CKINVDCx5p33_ASAP7_75t_R g446 ( 
.A(n_258),
.Y(n_446)
);

INVx1_ASAP7_75t_L g447 ( 
.A(n_230),
.Y(n_447)
);

INVx1_ASAP7_75t_L g448 ( 
.A(n_239),
.Y(n_448)
);

INVx1_ASAP7_75t_L g449 ( 
.A(n_243),
.Y(n_449)
);

BUFx2_ASAP7_75t_L g450 ( 
.A(n_231),
.Y(n_450)
);

INVx1_ASAP7_75t_L g451 ( 
.A(n_252),
.Y(n_451)
);

CKINVDCx20_ASAP7_75t_R g452 ( 
.A(n_390),
.Y(n_452)
);

INVx1_ASAP7_75t_L g453 ( 
.A(n_315),
.Y(n_453)
);

HB1xp67_ASAP7_75t_L g454 ( 
.A(n_233),
.Y(n_454)
);

INVx2_ASAP7_75t_L g455 ( 
.A(n_238),
.Y(n_455)
);

INVxp67_ASAP7_75t_SL g456 ( 
.A(n_270),
.Y(n_456)
);

INVxp33_ASAP7_75t_L g457 ( 
.A(n_284),
.Y(n_457)
);

CKINVDCx5p33_ASAP7_75t_R g458 ( 
.A(n_265),
.Y(n_458)
);

INVx1_ASAP7_75t_L g459 ( 
.A(n_350),
.Y(n_459)
);

INVxp67_ASAP7_75t_SL g460 ( 
.A(n_286),
.Y(n_460)
);

INVx2_ASAP7_75t_L g461 ( 
.A(n_260),
.Y(n_461)
);

INVx1_ASAP7_75t_L g462 ( 
.A(n_350),
.Y(n_462)
);

INVxp67_ASAP7_75t_SL g463 ( 
.A(n_304),
.Y(n_463)
);

CKINVDCx5p33_ASAP7_75t_R g464 ( 
.A(n_277),
.Y(n_464)
);

INVx2_ASAP7_75t_L g465 ( 
.A(n_260),
.Y(n_465)
);

INVx1_ASAP7_75t_L g466 ( 
.A(n_367),
.Y(n_466)
);

INVx1_ASAP7_75t_L g467 ( 
.A(n_367),
.Y(n_467)
);

INVxp67_ASAP7_75t_L g468 ( 
.A(n_266),
.Y(n_468)
);

INVx1_ASAP7_75t_L g469 ( 
.A(n_310),
.Y(n_469)
);

INVx2_ASAP7_75t_L g470 ( 
.A(n_382),
.Y(n_470)
);

INVxp67_ASAP7_75t_SL g471 ( 
.A(n_313),
.Y(n_471)
);

CKINVDCx5p33_ASAP7_75t_R g472 ( 
.A(n_278),
.Y(n_472)
);

CKINVDCx20_ASAP7_75t_R g473 ( 
.A(n_242),
.Y(n_473)
);

INVx2_ASAP7_75t_L g474 ( 
.A(n_382),
.Y(n_474)
);

INVx1_ASAP7_75t_L g475 ( 
.A(n_349),
.Y(n_475)
);

INVx2_ASAP7_75t_L g476 ( 
.A(n_212),
.Y(n_476)
);

CKINVDCx5p33_ASAP7_75t_R g477 ( 
.A(n_281),
.Y(n_477)
);

INVx1_ASAP7_75t_L g478 ( 
.A(n_352),
.Y(n_478)
);

INVx2_ASAP7_75t_L g479 ( 
.A(n_214),
.Y(n_479)
);

INVxp67_ASAP7_75t_L g480 ( 
.A(n_266),
.Y(n_480)
);

CKINVDCx16_ASAP7_75t_R g481 ( 
.A(n_266),
.Y(n_481)
);

CKINVDCx5p33_ASAP7_75t_R g482 ( 
.A(n_285),
.Y(n_482)
);

INVx1_ASAP7_75t_L g483 ( 
.A(n_356),
.Y(n_483)
);

INVxp67_ASAP7_75t_SL g484 ( 
.A(n_371),
.Y(n_484)
);

INVx1_ASAP7_75t_L g485 ( 
.A(n_374),
.Y(n_485)
);

INVx1_ASAP7_75t_L g486 ( 
.A(n_392),
.Y(n_486)
);

INVx1_ASAP7_75t_L g487 ( 
.A(n_393),
.Y(n_487)
);

INVx1_ASAP7_75t_L g488 ( 
.A(n_394),
.Y(n_488)
);

INVx1_ASAP7_75t_L g489 ( 
.A(n_216),
.Y(n_489)
);

INVx1_ASAP7_75t_L g490 ( 
.A(n_223),
.Y(n_490)
);

CKINVDCx20_ASAP7_75t_R g491 ( 
.A(n_242),
.Y(n_491)
);

INVx1_ASAP7_75t_L g492 ( 
.A(n_236),
.Y(n_492)
);

INVxp33_ASAP7_75t_SL g493 ( 
.A(n_233),
.Y(n_493)
);

INVx1_ASAP7_75t_L g494 ( 
.A(n_237),
.Y(n_494)
);

INVx1_ASAP7_75t_L g495 ( 
.A(n_245),
.Y(n_495)
);

INVxp67_ASAP7_75t_SL g496 ( 
.A(n_208),
.Y(n_496)
);

CKINVDCx5p33_ASAP7_75t_R g497 ( 
.A(n_290),
.Y(n_497)
);

CKINVDCx16_ASAP7_75t_R g498 ( 
.A(n_321),
.Y(n_498)
);

AND2x4_ASAP7_75t_L g499 ( 
.A(n_489),
.B(n_302),
.Y(n_499)
);

INVx1_ASAP7_75t_L g500 ( 
.A(n_400),
.Y(n_500)
);

INVx2_ASAP7_75t_L g501 ( 
.A(n_400),
.Y(n_501)
);

BUFx2_ASAP7_75t_SL g502 ( 
.A(n_473),
.Y(n_502)
);

INVx1_ASAP7_75t_L g503 ( 
.A(n_401),
.Y(n_503)
);

AND2x4_ASAP7_75t_L g504 ( 
.A(n_489),
.B(n_343),
.Y(n_504)
);

AND2x2_ASAP7_75t_L g505 ( 
.A(n_457),
.B(n_321),
.Y(n_505)
);

CKINVDCx20_ASAP7_75t_R g506 ( 
.A(n_442),
.Y(n_506)
);

INVx2_ASAP7_75t_L g507 ( 
.A(n_401),
.Y(n_507)
);

BUFx6f_ASAP7_75t_L g508 ( 
.A(n_402),
.Y(n_508)
);

INVx1_ASAP7_75t_L g509 ( 
.A(n_402),
.Y(n_509)
);

BUFx3_ASAP7_75t_L g510 ( 
.A(n_410),
.Y(n_510)
);

INVx1_ASAP7_75t_L g511 ( 
.A(n_403),
.Y(n_511)
);

INVx1_ASAP7_75t_L g512 ( 
.A(n_403),
.Y(n_512)
);

NAND2x1p5_ASAP7_75t_L g513 ( 
.A(n_490),
.B(n_201),
.Y(n_513)
);

BUFx6f_ASAP7_75t_L g514 ( 
.A(n_405),
.Y(n_514)
);

INVx3_ASAP7_75t_L g515 ( 
.A(n_405),
.Y(n_515)
);

AND2x4_ASAP7_75t_L g516 ( 
.A(n_490),
.B(n_218),
.Y(n_516)
);

INVx1_ASAP7_75t_L g517 ( 
.A(n_427),
.Y(n_517)
);

AND2x4_ASAP7_75t_L g518 ( 
.A(n_492),
.B(n_306),
.Y(n_518)
);

INVx1_ASAP7_75t_L g519 ( 
.A(n_427),
.Y(n_519)
);

INVxp67_ASAP7_75t_SL g520 ( 
.A(n_410),
.Y(n_520)
);

NAND2xp5_ASAP7_75t_L g521 ( 
.A(n_455),
.B(n_251),
.Y(n_521)
);

AND2x2_ASAP7_75t_SL g522 ( 
.A(n_444),
.B(n_200),
.Y(n_522)
);

INVx3_ASAP7_75t_L g523 ( 
.A(n_476),
.Y(n_523)
);

INVx2_ASAP7_75t_L g524 ( 
.A(n_428),
.Y(n_524)
);

BUFx6f_ASAP7_75t_L g525 ( 
.A(n_428),
.Y(n_525)
);

CKINVDCx5p33_ASAP7_75t_R g526 ( 
.A(n_411),
.Y(n_526)
);

OAI22xp5_ASAP7_75t_SL g527 ( 
.A1(n_443),
.A2(n_235),
.B1(n_246),
.B2(n_395),
.Y(n_527)
);

INVxp67_ASAP7_75t_SL g528 ( 
.A(n_455),
.Y(n_528)
);

INVx1_ASAP7_75t_L g529 ( 
.A(n_430),
.Y(n_529)
);

INVx1_ASAP7_75t_L g530 ( 
.A(n_430),
.Y(n_530)
);

INVx4_ASAP7_75t_L g531 ( 
.A(n_476),
.Y(n_531)
);

INVx1_ASAP7_75t_L g532 ( 
.A(n_433),
.Y(n_532)
);

INVx2_ASAP7_75t_L g533 ( 
.A(n_433),
.Y(n_533)
);

INVx2_ASAP7_75t_L g534 ( 
.A(n_434),
.Y(n_534)
);

CKINVDCx6p67_ASAP7_75t_R g535 ( 
.A(n_407),
.Y(n_535)
);

INVx1_ASAP7_75t_L g536 ( 
.A(n_434),
.Y(n_536)
);

INVx3_ASAP7_75t_L g537 ( 
.A(n_479),
.Y(n_537)
);

AND2x2_ASAP7_75t_SL g538 ( 
.A(n_444),
.B(n_200),
.Y(n_538)
);

NAND2xp5_ASAP7_75t_L g539 ( 
.A(n_461),
.B(n_253),
.Y(n_539)
);

AND2x4_ASAP7_75t_L g540 ( 
.A(n_492),
.B(n_240),
.Y(n_540)
);

INVx2_ASAP7_75t_L g541 ( 
.A(n_436),
.Y(n_541)
);

BUFx6f_ASAP7_75t_L g542 ( 
.A(n_436),
.Y(n_542)
);

BUFx6f_ASAP7_75t_L g543 ( 
.A(n_439),
.Y(n_543)
);

AND2x4_ASAP7_75t_L g544 ( 
.A(n_494),
.B(n_240),
.Y(n_544)
);

AND2x2_ASAP7_75t_L g545 ( 
.A(n_398),
.B(n_336),
.Y(n_545)
);

AND2x4_ASAP7_75t_L g546 ( 
.A(n_494),
.B(n_396),
.Y(n_546)
);

OAI22xp5_ASAP7_75t_SL g547 ( 
.A1(n_452),
.A2(n_246),
.B1(n_235),
.B2(n_395),
.Y(n_547)
);

BUFx6f_ASAP7_75t_L g548 ( 
.A(n_439),
.Y(n_548)
);

NOR2xp33_ASAP7_75t_R g549 ( 
.A(n_409),
.B(n_250),
.Y(n_549)
);

OA21x2_ASAP7_75t_L g550 ( 
.A1(n_440),
.A2(n_263),
.B(n_254),
.Y(n_550)
);

CKINVDCx5p33_ASAP7_75t_R g551 ( 
.A(n_417),
.Y(n_551)
);

INVx1_ASAP7_75t_L g552 ( 
.A(n_440),
.Y(n_552)
);

NAND2xp5_ASAP7_75t_L g553 ( 
.A(n_461),
.B(n_465),
.Y(n_553)
);

CKINVDCx5p33_ASAP7_75t_R g554 ( 
.A(n_421),
.Y(n_554)
);

NAND2xp5_ASAP7_75t_L g555 ( 
.A(n_465),
.B(n_264),
.Y(n_555)
);

INVx1_ASAP7_75t_L g556 ( 
.A(n_441),
.Y(n_556)
);

INVx1_ASAP7_75t_L g557 ( 
.A(n_441),
.Y(n_557)
);

BUFx6f_ASAP7_75t_L g558 ( 
.A(n_453),
.Y(n_558)
);

NOR2xp33_ASAP7_75t_SL g559 ( 
.A(n_491),
.B(n_242),
.Y(n_559)
);

HB1xp67_ASAP7_75t_L g560 ( 
.A(n_432),
.Y(n_560)
);

BUFx6f_ASAP7_75t_L g561 ( 
.A(n_453),
.Y(n_561)
);

INVx1_ASAP7_75t_L g562 ( 
.A(n_459),
.Y(n_562)
);

BUFx8_ASAP7_75t_L g563 ( 
.A(n_450),
.Y(n_563)
);

BUFx6f_ASAP7_75t_L g564 ( 
.A(n_459),
.Y(n_564)
);

OR2x2_ASAP7_75t_L g565 ( 
.A(n_424),
.B(n_353),
.Y(n_565)
);

INVx1_ASAP7_75t_L g566 ( 
.A(n_462),
.Y(n_566)
);

INVx1_ASAP7_75t_L g567 ( 
.A(n_462),
.Y(n_567)
);

NOR2xp33_ASAP7_75t_L g568 ( 
.A(n_496),
.B(n_372),
.Y(n_568)
);

INVx1_ASAP7_75t_L g569 ( 
.A(n_466),
.Y(n_569)
);

INVx1_ASAP7_75t_L g570 ( 
.A(n_466),
.Y(n_570)
);

INVx2_ASAP7_75t_L g571 ( 
.A(n_467),
.Y(n_571)
);

CKINVDCx5p33_ASAP7_75t_R g572 ( 
.A(n_422),
.Y(n_572)
);

BUFx6f_ASAP7_75t_L g573 ( 
.A(n_467),
.Y(n_573)
);

INVx2_ASAP7_75t_L g574 ( 
.A(n_479),
.Y(n_574)
);

INVx2_ASAP7_75t_L g575 ( 
.A(n_470),
.Y(n_575)
);

INVx2_ASAP7_75t_L g576 ( 
.A(n_470),
.Y(n_576)
);

INVx3_ASAP7_75t_L g577 ( 
.A(n_474),
.Y(n_577)
);

BUFx2_ASAP7_75t_L g578 ( 
.A(n_450),
.Y(n_578)
);

NAND2xp5_ASAP7_75t_L g579 ( 
.A(n_474),
.B(n_267),
.Y(n_579)
);

AND2x4_ASAP7_75t_L g580 ( 
.A(n_495),
.B(n_396),
.Y(n_580)
);

AND2x2_ASAP7_75t_L g581 ( 
.A(n_522),
.B(n_495),
.Y(n_581)
);

INVx2_ASAP7_75t_SL g582 ( 
.A(n_522),
.Y(n_582)
);

INVx2_ASAP7_75t_L g583 ( 
.A(n_515),
.Y(n_583)
);

NAND2xp5_ASAP7_75t_SL g584 ( 
.A(n_522),
.B(n_538),
.Y(n_584)
);

INVx2_ASAP7_75t_L g585 ( 
.A(n_515),
.Y(n_585)
);

NOR2xp33_ASAP7_75t_L g586 ( 
.A(n_513),
.B(n_425),
.Y(n_586)
);

INVx2_ASAP7_75t_L g587 ( 
.A(n_515),
.Y(n_587)
);

BUFx3_ASAP7_75t_L g588 ( 
.A(n_510),
.Y(n_588)
);

INVx1_ASAP7_75t_L g589 ( 
.A(n_500),
.Y(n_589)
);

NAND2xp5_ASAP7_75t_L g590 ( 
.A(n_538),
.B(n_435),
.Y(n_590)
);

INVx2_ASAP7_75t_L g591 ( 
.A(n_515),
.Y(n_591)
);

INVx1_ASAP7_75t_L g592 ( 
.A(n_500),
.Y(n_592)
);

BUFx3_ASAP7_75t_L g593 ( 
.A(n_510),
.Y(n_593)
);

INVx2_ASAP7_75t_L g594 ( 
.A(n_508),
.Y(n_594)
);

CKINVDCx5p33_ASAP7_75t_R g595 ( 
.A(n_526),
.Y(n_595)
);

BUFx10_ASAP7_75t_L g596 ( 
.A(n_538),
.Y(n_596)
);

HB1xp67_ASAP7_75t_L g597 ( 
.A(n_578),
.Y(n_597)
);

NAND2xp5_ASAP7_75t_SL g598 ( 
.A(n_499),
.B(n_504),
.Y(n_598)
);

INVx2_ASAP7_75t_L g599 ( 
.A(n_508),
.Y(n_599)
);

AOI22xp33_ASAP7_75t_L g600 ( 
.A1(n_499),
.A2(n_404),
.B1(n_493),
.B2(n_431),
.Y(n_600)
);

BUFx2_ASAP7_75t_L g601 ( 
.A(n_578),
.Y(n_601)
);

INVx2_ASAP7_75t_L g602 ( 
.A(n_508),
.Y(n_602)
);

INVx3_ASAP7_75t_L g603 ( 
.A(n_508),
.Y(n_603)
);

NAND2xp5_ASAP7_75t_L g604 ( 
.A(n_520),
.B(n_438),
.Y(n_604)
);

INVx1_ASAP7_75t_L g605 ( 
.A(n_503),
.Y(n_605)
);

INVx2_ASAP7_75t_L g606 ( 
.A(n_501),
.Y(n_606)
);

INVx2_ASAP7_75t_L g607 ( 
.A(n_501),
.Y(n_607)
);

INVx2_ASAP7_75t_L g608 ( 
.A(n_507),
.Y(n_608)
);

NAND2xp5_ASAP7_75t_L g609 ( 
.A(n_528),
.B(n_446),
.Y(n_609)
);

OAI22xp5_ASAP7_75t_L g610 ( 
.A1(n_499),
.A2(n_348),
.B1(n_354),
.B2(n_345),
.Y(n_610)
);

INVx2_ASAP7_75t_L g611 ( 
.A(n_507),
.Y(n_611)
);

INVx1_ASAP7_75t_L g612 ( 
.A(n_503),
.Y(n_612)
);

INVx1_ASAP7_75t_L g613 ( 
.A(n_509),
.Y(n_613)
);

INVx2_ASAP7_75t_L g614 ( 
.A(n_525),
.Y(n_614)
);

NAND2xp5_ASAP7_75t_SL g615 ( 
.A(n_499),
.B(n_458),
.Y(n_615)
);

OAI21xp33_ASAP7_75t_SL g616 ( 
.A1(n_568),
.A2(n_545),
.B(n_505),
.Y(n_616)
);

INVx1_ASAP7_75t_L g617 ( 
.A(n_509),
.Y(n_617)
);

NAND2xp5_ASAP7_75t_SL g618 ( 
.A(n_504),
.B(n_464),
.Y(n_618)
);

INVx2_ASAP7_75t_L g619 ( 
.A(n_508),
.Y(n_619)
);

INVx2_ASAP7_75t_L g620 ( 
.A(n_508),
.Y(n_620)
);

BUFx6f_ASAP7_75t_L g621 ( 
.A(n_525),
.Y(n_621)
);

INVx2_ASAP7_75t_L g622 ( 
.A(n_514),
.Y(n_622)
);

NAND2xp5_ASAP7_75t_SL g623 ( 
.A(n_504),
.B(n_472),
.Y(n_623)
);

CKINVDCx5p33_ASAP7_75t_R g624 ( 
.A(n_551),
.Y(n_624)
);

BUFx3_ASAP7_75t_L g625 ( 
.A(n_577),
.Y(n_625)
);

INVx2_ASAP7_75t_L g626 ( 
.A(n_514),
.Y(n_626)
);

INVx3_ASAP7_75t_L g627 ( 
.A(n_514),
.Y(n_627)
);

AND2x2_ASAP7_75t_L g628 ( 
.A(n_505),
.B(n_456),
.Y(n_628)
);

INVx1_ASAP7_75t_L g629 ( 
.A(n_511),
.Y(n_629)
);

INVx2_ASAP7_75t_L g630 ( 
.A(n_514),
.Y(n_630)
);

AND2x4_ASAP7_75t_L g631 ( 
.A(n_504),
.B(n_460),
.Y(n_631)
);

INVx1_ASAP7_75t_L g632 ( 
.A(n_511),
.Y(n_632)
);

INVx4_ASAP7_75t_L g633 ( 
.A(n_550),
.Y(n_633)
);

NOR2xp33_ASAP7_75t_L g634 ( 
.A(n_513),
.B(n_477),
.Y(n_634)
);

INVx2_ASAP7_75t_L g635 ( 
.A(n_514),
.Y(n_635)
);

INVx3_ASAP7_75t_L g636 ( 
.A(n_514),
.Y(n_636)
);

INVx1_ASAP7_75t_L g637 ( 
.A(n_512),
.Y(n_637)
);

OAI22xp5_ASAP7_75t_L g638 ( 
.A1(n_513),
.A2(n_348),
.B1(n_354),
.B2(n_345),
.Y(n_638)
);

INVx2_ASAP7_75t_L g639 ( 
.A(n_525),
.Y(n_639)
);

NAND2xp5_ASAP7_75t_SL g640 ( 
.A(n_549),
.B(n_482),
.Y(n_640)
);

INVx2_ASAP7_75t_L g641 ( 
.A(n_525),
.Y(n_641)
);

INVx1_ASAP7_75t_L g642 ( 
.A(n_512),
.Y(n_642)
);

INVxp67_ASAP7_75t_L g643 ( 
.A(n_565),
.Y(n_643)
);

BUFx3_ASAP7_75t_L g644 ( 
.A(n_577),
.Y(n_644)
);

OR2x2_ASAP7_75t_L g645 ( 
.A(n_565),
.B(n_481),
.Y(n_645)
);

AOI22xp33_ASAP7_75t_L g646 ( 
.A1(n_516),
.A2(n_454),
.B1(n_471),
.B2(n_463),
.Y(n_646)
);

NAND2xp5_ASAP7_75t_SL g647 ( 
.A(n_516),
.B(n_497),
.Y(n_647)
);

INVx2_ASAP7_75t_L g648 ( 
.A(n_525),
.Y(n_648)
);

CKINVDCx5p33_ASAP7_75t_R g649 ( 
.A(n_554),
.Y(n_649)
);

CKINVDCx5p33_ASAP7_75t_R g650 ( 
.A(n_572),
.Y(n_650)
);

INVx2_ASAP7_75t_L g651 ( 
.A(n_525),
.Y(n_651)
);

INVx2_ASAP7_75t_L g652 ( 
.A(n_542),
.Y(n_652)
);

NAND2xp5_ASAP7_75t_L g653 ( 
.A(n_540),
.B(n_468),
.Y(n_653)
);

AOI22xp5_ASAP7_75t_L g654 ( 
.A1(n_516),
.A2(n_375),
.B1(n_377),
.B2(n_373),
.Y(n_654)
);

INVx2_ASAP7_75t_L g655 ( 
.A(n_542),
.Y(n_655)
);

INVx2_ASAP7_75t_L g656 ( 
.A(n_542),
.Y(n_656)
);

NAND2xp5_ASAP7_75t_L g657 ( 
.A(n_540),
.B(n_480),
.Y(n_657)
);

INVx2_ASAP7_75t_L g658 ( 
.A(n_542),
.Y(n_658)
);

NAND2xp5_ASAP7_75t_SL g659 ( 
.A(n_518),
.B(n_498),
.Y(n_659)
);

INVxp67_ASAP7_75t_SL g660 ( 
.A(n_553),
.Y(n_660)
);

INVxp33_ASAP7_75t_L g661 ( 
.A(n_527),
.Y(n_661)
);

CKINVDCx6p67_ASAP7_75t_R g662 ( 
.A(n_535),
.Y(n_662)
);

NAND2xp5_ASAP7_75t_SL g663 ( 
.A(n_518),
.B(n_202),
.Y(n_663)
);

OAI22xp33_ASAP7_75t_L g664 ( 
.A1(n_559),
.A2(n_429),
.B1(n_437),
.B2(n_379),
.Y(n_664)
);

INVx3_ASAP7_75t_L g665 ( 
.A(n_542),
.Y(n_665)
);

INVx2_ASAP7_75t_L g666 ( 
.A(n_542),
.Y(n_666)
);

CKINVDCx5p33_ASAP7_75t_R g667 ( 
.A(n_506),
.Y(n_667)
);

INVx2_ASAP7_75t_SL g668 ( 
.A(n_540),
.Y(n_668)
);

INVx2_ASAP7_75t_L g669 ( 
.A(n_543),
.Y(n_669)
);

INVx2_ASAP7_75t_L g670 ( 
.A(n_543),
.Y(n_670)
);

NOR2xp33_ASAP7_75t_L g671 ( 
.A(n_531),
.B(n_415),
.Y(n_671)
);

INVx2_ASAP7_75t_SL g672 ( 
.A(n_540),
.Y(n_672)
);

INVx1_ASAP7_75t_L g673 ( 
.A(n_543),
.Y(n_673)
);

INVx2_ASAP7_75t_L g674 ( 
.A(n_543),
.Y(n_674)
);

INVx1_ASAP7_75t_L g675 ( 
.A(n_543),
.Y(n_675)
);

NAND2xp5_ASAP7_75t_SL g676 ( 
.A(n_518),
.B(n_202),
.Y(n_676)
);

INVx2_ASAP7_75t_L g677 ( 
.A(n_543),
.Y(n_677)
);

INVx5_ASAP7_75t_L g678 ( 
.A(n_548),
.Y(n_678)
);

NAND2xp5_ASAP7_75t_SL g679 ( 
.A(n_518),
.B(n_203),
.Y(n_679)
);

INVx2_ASAP7_75t_L g680 ( 
.A(n_548),
.Y(n_680)
);

INVx2_ASAP7_75t_L g681 ( 
.A(n_548),
.Y(n_681)
);

INVx1_ASAP7_75t_L g682 ( 
.A(n_548),
.Y(n_682)
);

AOI22xp5_ASAP7_75t_L g683 ( 
.A1(n_545),
.A2(n_547),
.B1(n_546),
.B2(n_544),
.Y(n_683)
);

OAI22xp33_ASAP7_75t_L g684 ( 
.A1(n_560),
.A2(n_388),
.B1(n_389),
.B2(n_391),
.Y(n_684)
);

INVx1_ASAP7_75t_L g685 ( 
.A(n_548),
.Y(n_685)
);

NAND2xp5_ASAP7_75t_SL g686 ( 
.A(n_544),
.B(n_203),
.Y(n_686)
);

INVx2_ASAP7_75t_L g687 ( 
.A(n_548),
.Y(n_687)
);

OAI22xp33_ASAP7_75t_L g688 ( 
.A1(n_531),
.A2(n_361),
.B1(n_369),
.B2(n_359),
.Y(n_688)
);

INVx1_ASAP7_75t_L g689 ( 
.A(n_558),
.Y(n_689)
);

NOR2x1p5_ASAP7_75t_L g690 ( 
.A(n_535),
.B(n_484),
.Y(n_690)
);

INVx2_ASAP7_75t_SL g691 ( 
.A(n_544),
.Y(n_691)
);

INVx1_ASAP7_75t_L g692 ( 
.A(n_558),
.Y(n_692)
);

INVx2_ASAP7_75t_L g693 ( 
.A(n_558),
.Y(n_693)
);

INVx1_ASAP7_75t_L g694 ( 
.A(n_558),
.Y(n_694)
);

INVx1_ASAP7_75t_L g695 ( 
.A(n_558),
.Y(n_695)
);

NAND3xp33_ASAP7_75t_L g696 ( 
.A(n_531),
.B(n_361),
.C(n_359),
.Y(n_696)
);

OA22x2_ASAP7_75t_L g697 ( 
.A1(n_517),
.A2(n_399),
.B1(n_451),
.B2(n_445),
.Y(n_697)
);

INVx3_ASAP7_75t_L g698 ( 
.A(n_558),
.Y(n_698)
);

INVx4_ASAP7_75t_L g699 ( 
.A(n_550),
.Y(n_699)
);

INVx2_ASAP7_75t_SL g700 ( 
.A(n_546),
.Y(n_700)
);

OAI22xp33_ASAP7_75t_L g701 ( 
.A1(n_531),
.A2(n_385),
.B1(n_388),
.B2(n_389),
.Y(n_701)
);

NAND2xp5_ASAP7_75t_SL g702 ( 
.A(n_546),
.B(n_204),
.Y(n_702)
);

INVx1_ASAP7_75t_L g703 ( 
.A(n_561),
.Y(n_703)
);

INVx3_ASAP7_75t_L g704 ( 
.A(n_561),
.Y(n_704)
);

NOR2xp33_ASAP7_75t_L g705 ( 
.A(n_546),
.B(n_580),
.Y(n_705)
);

INVx2_ASAP7_75t_L g706 ( 
.A(n_561),
.Y(n_706)
);

INVx1_ASAP7_75t_L g707 ( 
.A(n_561),
.Y(n_707)
);

NAND3xp33_ASAP7_75t_L g708 ( 
.A(n_580),
.B(n_373),
.C(n_369),
.Y(n_708)
);

NOR2xp33_ASAP7_75t_L g709 ( 
.A(n_580),
.B(n_447),
.Y(n_709)
);

INVx2_ASAP7_75t_L g710 ( 
.A(n_561),
.Y(n_710)
);

NOR2xp33_ASAP7_75t_L g711 ( 
.A(n_580),
.B(n_521),
.Y(n_711)
);

INVx1_ASAP7_75t_L g712 ( 
.A(n_561),
.Y(n_712)
);

NAND2xp5_ASAP7_75t_SL g713 ( 
.A(n_563),
.B(n_204),
.Y(n_713)
);

INVx1_ASAP7_75t_L g714 ( 
.A(n_564),
.Y(n_714)
);

INVx2_ASAP7_75t_L g715 ( 
.A(n_564),
.Y(n_715)
);

INVx2_ASAP7_75t_L g716 ( 
.A(n_564),
.Y(n_716)
);

INVx2_ASAP7_75t_L g717 ( 
.A(n_564),
.Y(n_717)
);

INVx2_ASAP7_75t_L g718 ( 
.A(n_564),
.Y(n_718)
);

INVx1_ASAP7_75t_L g719 ( 
.A(n_564),
.Y(n_719)
);

CKINVDCx11_ASAP7_75t_R g720 ( 
.A(n_563),
.Y(n_720)
);

INVx2_ASAP7_75t_L g721 ( 
.A(n_573),
.Y(n_721)
);

BUFx2_ASAP7_75t_L g722 ( 
.A(n_563),
.Y(n_722)
);

INVx1_ASAP7_75t_L g723 ( 
.A(n_573),
.Y(n_723)
);

NOR2xp33_ASAP7_75t_L g724 ( 
.A(n_539),
.B(n_448),
.Y(n_724)
);

INVxp67_ASAP7_75t_SL g725 ( 
.A(n_577),
.Y(n_725)
);

INVx2_ASAP7_75t_L g726 ( 
.A(n_573),
.Y(n_726)
);

INVx1_ASAP7_75t_L g727 ( 
.A(n_573),
.Y(n_727)
);

INVx3_ASAP7_75t_L g728 ( 
.A(n_573),
.Y(n_728)
);

AOI22xp33_ASAP7_75t_L g729 ( 
.A1(n_550),
.A2(n_449),
.B1(n_336),
.B2(n_341),
.Y(n_729)
);

INVx2_ASAP7_75t_L g730 ( 
.A(n_573),
.Y(n_730)
);

INVx1_ASAP7_75t_L g731 ( 
.A(n_574),
.Y(n_731)
);

OAI22xp33_ASAP7_75t_L g732 ( 
.A1(n_661),
.A2(n_519),
.B1(n_529),
.B2(n_517),
.Y(n_732)
);

NAND2xp5_ASAP7_75t_L g733 ( 
.A(n_581),
.B(n_577),
.Y(n_733)
);

HB1xp67_ASAP7_75t_L g734 ( 
.A(n_631),
.Y(n_734)
);

NAND2xp5_ASAP7_75t_SL g735 ( 
.A(n_596),
.B(n_563),
.Y(n_735)
);

NAND2xp5_ASAP7_75t_L g736 ( 
.A(n_581),
.B(n_523),
.Y(n_736)
);

NAND2xp5_ASAP7_75t_SL g737 ( 
.A(n_596),
.B(n_205),
.Y(n_737)
);

OR2x2_ASAP7_75t_L g738 ( 
.A(n_643),
.B(n_502),
.Y(n_738)
);

AND2x2_ASAP7_75t_L g739 ( 
.A(n_631),
.B(n_502),
.Y(n_739)
);

NAND2xp33_ASAP7_75t_L g740 ( 
.A(n_582),
.B(n_205),
.Y(n_740)
);

OAI22xp5_ASAP7_75t_L g741 ( 
.A1(n_582),
.A2(n_377),
.B1(n_379),
.B2(n_375),
.Y(n_741)
);

INVx1_ASAP7_75t_L g742 ( 
.A(n_589),
.Y(n_742)
);

INVx2_ASAP7_75t_L g743 ( 
.A(n_625),
.Y(n_743)
);

INVx1_ASAP7_75t_L g744 ( 
.A(n_589),
.Y(n_744)
);

INVx1_ASAP7_75t_L g745 ( 
.A(n_592),
.Y(n_745)
);

NAND2xp33_ASAP7_75t_L g746 ( 
.A(n_595),
.B(n_206),
.Y(n_746)
);

NAND2xp5_ASAP7_75t_SL g747 ( 
.A(n_596),
.B(n_616),
.Y(n_747)
);

OAI22xp5_ASAP7_75t_L g748 ( 
.A1(n_584),
.A2(n_380),
.B1(n_385),
.B2(n_391),
.Y(n_748)
);

NAND2xp5_ASAP7_75t_L g749 ( 
.A(n_711),
.B(n_523),
.Y(n_749)
);

INVx1_ASAP7_75t_L g750 ( 
.A(n_592),
.Y(n_750)
);

INVx8_ASAP7_75t_L g751 ( 
.A(n_631),
.Y(n_751)
);

AO22x2_ASAP7_75t_L g752 ( 
.A1(n_598),
.A2(n_532),
.B1(n_536),
.B2(n_530),
.Y(n_752)
);

NAND2xp5_ASAP7_75t_SL g753 ( 
.A(n_596),
.B(n_206),
.Y(n_753)
);

NAND3xp33_ASAP7_75t_L g754 ( 
.A(n_600),
.B(n_380),
.C(n_303),
.Y(n_754)
);

NAND2xp5_ASAP7_75t_SL g755 ( 
.A(n_616),
.B(n_207),
.Y(n_755)
);

INVx2_ASAP7_75t_L g756 ( 
.A(n_625),
.Y(n_756)
);

NAND2xp5_ASAP7_75t_L g757 ( 
.A(n_668),
.B(n_523),
.Y(n_757)
);

AND2x2_ASAP7_75t_SL g758 ( 
.A(n_722),
.B(n_550),
.Y(n_758)
);

NOR2xp33_ASAP7_75t_L g759 ( 
.A(n_590),
.B(n_555),
.Y(n_759)
);

INVx2_ASAP7_75t_L g760 ( 
.A(n_625),
.Y(n_760)
);

NAND2xp5_ASAP7_75t_L g761 ( 
.A(n_668),
.B(n_523),
.Y(n_761)
);

INVx1_ASAP7_75t_L g762 ( 
.A(n_605),
.Y(n_762)
);

INVx2_ASAP7_75t_L g763 ( 
.A(n_644),
.Y(n_763)
);

INVx4_ASAP7_75t_L g764 ( 
.A(n_588),
.Y(n_764)
);

NAND2xp33_ASAP7_75t_SL g765 ( 
.A(n_624),
.B(n_423),
.Y(n_765)
);

NAND2xp5_ASAP7_75t_SL g766 ( 
.A(n_586),
.B(n_207),
.Y(n_766)
);

INVx1_ASAP7_75t_L g767 ( 
.A(n_605),
.Y(n_767)
);

INVx1_ASAP7_75t_L g768 ( 
.A(n_612),
.Y(n_768)
);

INVx1_ASAP7_75t_L g769 ( 
.A(n_612),
.Y(n_769)
);

BUFx5_ASAP7_75t_L g770 ( 
.A(n_673),
.Y(n_770)
);

INVx2_ASAP7_75t_L g771 ( 
.A(n_606),
.Y(n_771)
);

NAND2xp5_ASAP7_75t_SL g772 ( 
.A(n_634),
.B(n_210),
.Y(n_772)
);

INVx1_ASAP7_75t_L g773 ( 
.A(n_613),
.Y(n_773)
);

INVx2_ASAP7_75t_L g774 ( 
.A(n_606),
.Y(n_774)
);

NOR2xp33_ASAP7_75t_L g775 ( 
.A(n_604),
.B(n_609),
.Y(n_775)
);

NAND2xp5_ASAP7_75t_L g776 ( 
.A(n_672),
.B(n_537),
.Y(n_776)
);

NAND2xp5_ASAP7_75t_L g777 ( 
.A(n_672),
.B(n_537),
.Y(n_777)
);

INVx1_ASAP7_75t_L g778 ( 
.A(n_613),
.Y(n_778)
);

INVx1_ASAP7_75t_L g779 ( 
.A(n_617),
.Y(n_779)
);

BUFx6f_ASAP7_75t_L g780 ( 
.A(n_588),
.Y(n_780)
);

INVx1_ASAP7_75t_L g781 ( 
.A(n_617),
.Y(n_781)
);

INVx2_ASAP7_75t_L g782 ( 
.A(n_644),
.Y(n_782)
);

AOI22xp5_ASAP7_75t_L g783 ( 
.A1(n_691),
.A2(n_261),
.B1(n_537),
.B2(n_569),
.Y(n_783)
);

NAND2xp5_ASAP7_75t_SL g784 ( 
.A(n_631),
.B(n_691),
.Y(n_784)
);

INVx2_ASAP7_75t_L g785 ( 
.A(n_644),
.Y(n_785)
);

NAND2xp5_ASAP7_75t_SL g786 ( 
.A(n_700),
.B(n_210),
.Y(n_786)
);

BUFx6f_ASAP7_75t_L g787 ( 
.A(n_588),
.Y(n_787)
);

INVx2_ASAP7_75t_L g788 ( 
.A(n_593),
.Y(n_788)
);

BUFx6f_ASAP7_75t_SL g789 ( 
.A(n_662),
.Y(n_789)
);

NAND2xp5_ASAP7_75t_SL g790 ( 
.A(n_700),
.B(n_621),
.Y(n_790)
);

NAND2xp5_ASAP7_75t_L g791 ( 
.A(n_660),
.B(n_537),
.Y(n_791)
);

NAND2xp5_ASAP7_75t_SL g792 ( 
.A(n_621),
.B(n_213),
.Y(n_792)
);

NAND2xp5_ASAP7_75t_L g793 ( 
.A(n_705),
.B(n_724),
.Y(n_793)
);

NAND2xp5_ASAP7_75t_L g794 ( 
.A(n_628),
.B(n_575),
.Y(n_794)
);

NOR2xp33_ASAP7_75t_L g795 ( 
.A(n_663),
.B(n_579),
.Y(n_795)
);

NAND2xp5_ASAP7_75t_L g796 ( 
.A(n_628),
.B(n_575),
.Y(n_796)
);

AOI21xp5_ASAP7_75t_L g797 ( 
.A1(n_725),
.A2(n_529),
.B(n_519),
.Y(n_797)
);

INVx3_ASAP7_75t_L g798 ( 
.A(n_593),
.Y(n_798)
);

AND2x2_ASAP7_75t_L g799 ( 
.A(n_601),
.B(n_574),
.Y(n_799)
);

AOI22xp5_ASAP7_75t_L g800 ( 
.A1(n_683),
.A2(n_709),
.B1(n_676),
.B2(n_679),
.Y(n_800)
);

INVx1_ASAP7_75t_L g801 ( 
.A(n_629),
.Y(n_801)
);

NOR2xp33_ASAP7_75t_L g802 ( 
.A(n_647),
.B(n_576),
.Y(n_802)
);

INVxp67_ASAP7_75t_L g803 ( 
.A(n_601),
.Y(n_803)
);

INVxp67_ASAP7_75t_L g804 ( 
.A(n_597),
.Y(n_804)
);

AND2x2_ASAP7_75t_L g805 ( 
.A(n_645),
.B(n_469),
.Y(n_805)
);

INVx2_ASAP7_75t_L g806 ( 
.A(n_593),
.Y(n_806)
);

INVx3_ASAP7_75t_L g807 ( 
.A(n_583),
.Y(n_807)
);

AOI22xp33_ASAP7_75t_L g808 ( 
.A1(n_633),
.A2(n_571),
.B1(n_524),
.B2(n_533),
.Y(n_808)
);

INVx1_ASAP7_75t_L g809 ( 
.A(n_629),
.Y(n_809)
);

NOR2xp33_ASAP7_75t_L g810 ( 
.A(n_615),
.B(n_618),
.Y(n_810)
);

INVx1_ASAP7_75t_L g811 ( 
.A(n_632),
.Y(n_811)
);

AOI22xp33_ASAP7_75t_L g812 ( 
.A1(n_633),
.A2(n_571),
.B1(n_524),
.B2(n_533),
.Y(n_812)
);

INVx2_ASAP7_75t_L g813 ( 
.A(n_583),
.Y(n_813)
);

INVx2_ASAP7_75t_L g814 ( 
.A(n_607),
.Y(n_814)
);

BUFx3_ASAP7_75t_L g815 ( 
.A(n_649),
.Y(n_815)
);

NAND2xp5_ASAP7_75t_L g816 ( 
.A(n_653),
.B(n_530),
.Y(n_816)
);

INVx2_ASAP7_75t_L g817 ( 
.A(n_607),
.Y(n_817)
);

INVx1_ASAP7_75t_L g818 ( 
.A(n_632),
.Y(n_818)
);

NOR2xp33_ASAP7_75t_L g819 ( 
.A(n_623),
.B(n_532),
.Y(n_819)
);

INVx1_ASAP7_75t_L g820 ( 
.A(n_637),
.Y(n_820)
);

INVx3_ASAP7_75t_L g821 ( 
.A(n_583),
.Y(n_821)
);

NAND2xp5_ASAP7_75t_L g822 ( 
.A(n_657),
.B(n_536),
.Y(n_822)
);

NAND2xp5_ASAP7_75t_L g823 ( 
.A(n_646),
.B(n_552),
.Y(n_823)
);

NAND2xp5_ASAP7_75t_L g824 ( 
.A(n_729),
.B(n_552),
.Y(n_824)
);

INVx2_ASAP7_75t_SL g825 ( 
.A(n_645),
.Y(n_825)
);

NAND2xp5_ASAP7_75t_SL g826 ( 
.A(n_621),
.B(n_213),
.Y(n_826)
);

NAND2xp5_ASAP7_75t_L g827 ( 
.A(n_731),
.B(n_556),
.Y(n_827)
);

NAND2xp33_ASAP7_75t_L g828 ( 
.A(n_650),
.B(n_215),
.Y(n_828)
);

INVx1_ASAP7_75t_L g829 ( 
.A(n_637),
.Y(n_829)
);

INVxp67_ASAP7_75t_L g830 ( 
.A(n_667),
.Y(n_830)
);

INVx1_ASAP7_75t_L g831 ( 
.A(n_642),
.Y(n_831)
);

NAND2xp33_ASAP7_75t_L g832 ( 
.A(n_621),
.B(n_215),
.Y(n_832)
);

INVxp67_ASAP7_75t_L g833 ( 
.A(n_671),
.Y(n_833)
);

NOR2xp67_ASAP7_75t_L g834 ( 
.A(n_640),
.B(n_696),
.Y(n_834)
);

A2O1A1Ixp33_ASAP7_75t_L g835 ( 
.A1(n_683),
.A2(n_570),
.B(n_569),
.C(n_567),
.Y(n_835)
);

NAND2xp5_ASAP7_75t_L g836 ( 
.A(n_731),
.B(n_556),
.Y(n_836)
);

NAND2xp5_ASAP7_75t_SL g837 ( 
.A(n_621),
.B(n_219),
.Y(n_837)
);

NAND2xp33_ASAP7_75t_L g838 ( 
.A(n_621),
.B(n_219),
.Y(n_838)
);

NOR2xp67_ASAP7_75t_L g839 ( 
.A(n_713),
.B(n_557),
.Y(n_839)
);

BUFx8_ASAP7_75t_L g840 ( 
.A(n_722),
.Y(n_840)
);

NOR3xp33_ASAP7_75t_L g841 ( 
.A(n_684),
.B(n_307),
.C(n_301),
.Y(n_841)
);

NAND2xp5_ASAP7_75t_SL g842 ( 
.A(n_585),
.B(n_220),
.Y(n_842)
);

AOI22xp33_ASAP7_75t_L g843 ( 
.A1(n_633),
.A2(n_699),
.B1(n_654),
.B2(n_697),
.Y(n_843)
);

AO22x2_ASAP7_75t_L g844 ( 
.A1(n_610),
.A2(n_570),
.B1(n_567),
.B2(n_566),
.Y(n_844)
);

AND2x2_ASAP7_75t_L g845 ( 
.A(n_654),
.B(n_475),
.Y(n_845)
);

NAND2xp5_ASAP7_75t_SL g846 ( 
.A(n_585),
.B(n_220),
.Y(n_846)
);

NAND2xp5_ASAP7_75t_L g847 ( 
.A(n_585),
.B(n_557),
.Y(n_847)
);

INVx1_ASAP7_75t_L g848 ( 
.A(n_642),
.Y(n_848)
);

NAND2xp5_ASAP7_75t_L g849 ( 
.A(n_587),
.B(n_562),
.Y(n_849)
);

AND2x2_ASAP7_75t_L g850 ( 
.A(n_690),
.B(n_475),
.Y(n_850)
);

NOR2xp33_ASAP7_75t_L g851 ( 
.A(n_659),
.B(n_562),
.Y(n_851)
);

INVx2_ASAP7_75t_L g852 ( 
.A(n_587),
.Y(n_852)
);

AND2x2_ASAP7_75t_L g853 ( 
.A(n_690),
.B(n_478),
.Y(n_853)
);

NAND2xp5_ASAP7_75t_L g854 ( 
.A(n_587),
.B(n_566),
.Y(n_854)
);

INVx2_ASAP7_75t_L g855 ( 
.A(n_591),
.Y(n_855)
);

NAND2xp5_ASAP7_75t_SL g856 ( 
.A(n_591),
.B(n_221),
.Y(n_856)
);

NAND2xp5_ASAP7_75t_L g857 ( 
.A(n_591),
.B(n_608),
.Y(n_857)
);

NAND2xp5_ASAP7_75t_L g858 ( 
.A(n_608),
.B(n_534),
.Y(n_858)
);

INVx4_ASAP7_75t_L g859 ( 
.A(n_678),
.Y(n_859)
);

AND2x2_ASAP7_75t_L g860 ( 
.A(n_638),
.B(n_478),
.Y(n_860)
);

INVx2_ASAP7_75t_SL g861 ( 
.A(n_697),
.Y(n_861)
);

NAND2xp5_ASAP7_75t_L g862 ( 
.A(n_611),
.B(n_665),
.Y(n_862)
);

AOI221xp5_ASAP7_75t_L g863 ( 
.A1(n_664),
.A2(n_483),
.B1(n_485),
.B2(n_488),
.C(n_487),
.Y(n_863)
);

A2O1A1Ixp33_ASAP7_75t_L g864 ( 
.A1(n_708),
.A2(n_541),
.B(n_534),
.C(n_488),
.Y(n_864)
);

AOI22xp33_ASAP7_75t_L g865 ( 
.A1(n_633),
.A2(n_541),
.B1(n_279),
.B2(n_341),
.Y(n_865)
);

NAND2xp5_ASAP7_75t_SL g866 ( 
.A(n_665),
.B(n_221),
.Y(n_866)
);

AOI221xp5_ASAP7_75t_L g867 ( 
.A1(n_688),
.A2(n_486),
.B1(n_485),
.B2(n_483),
.C(n_487),
.Y(n_867)
);

AOI22xp5_ASAP7_75t_L g868 ( 
.A1(n_686),
.A2(n_300),
.B1(n_222),
.B2(n_386),
.Y(n_868)
);

INVx1_ASAP7_75t_L g869 ( 
.A(n_697),
.Y(n_869)
);

NOR2xp67_ASAP7_75t_L g870 ( 
.A(n_665),
.B(n_486),
.Y(n_870)
);

INVx2_ASAP7_75t_L g871 ( 
.A(n_614),
.Y(n_871)
);

INVx3_ASAP7_75t_L g872 ( 
.A(n_698),
.Y(n_872)
);

INVx1_ASAP7_75t_L g873 ( 
.A(n_673),
.Y(n_873)
);

INVxp67_ASAP7_75t_L g874 ( 
.A(n_702),
.Y(n_874)
);

BUFx6f_ASAP7_75t_SL g875 ( 
.A(n_662),
.Y(n_875)
);

INVx2_ASAP7_75t_L g876 ( 
.A(n_614),
.Y(n_876)
);

INVxp67_ASAP7_75t_L g877 ( 
.A(n_701),
.Y(n_877)
);

NAND2xp5_ASAP7_75t_L g878 ( 
.A(n_698),
.B(n_704),
.Y(n_878)
);

AOI21xp5_ASAP7_75t_L g879 ( 
.A1(n_675),
.A2(n_275),
.B(n_274),
.Y(n_879)
);

NAND2xp5_ASAP7_75t_L g880 ( 
.A(n_698),
.B(n_704),
.Y(n_880)
);

INVx1_ASAP7_75t_SL g881 ( 
.A(n_720),
.Y(n_881)
);

INVx1_ASAP7_75t_L g882 ( 
.A(n_675),
.Y(n_882)
);

NAND2xp5_ASAP7_75t_L g883 ( 
.A(n_698),
.B(n_228),
.Y(n_883)
);

NOR2xp33_ASAP7_75t_L g884 ( 
.A(n_704),
.B(n_309),
.Y(n_884)
);

NAND2xp5_ASAP7_75t_L g885 ( 
.A(n_704),
.B(n_292),
.Y(n_885)
);

NAND2xp5_ASAP7_75t_L g886 ( 
.A(n_728),
.B(n_682),
.Y(n_886)
);

NAND2xp5_ASAP7_75t_L g887 ( 
.A(n_728),
.B(n_351),
.Y(n_887)
);

NAND2xp5_ASAP7_75t_L g888 ( 
.A(n_728),
.B(n_355),
.Y(n_888)
);

NAND2xp5_ASAP7_75t_L g889 ( 
.A(n_728),
.B(n_222),
.Y(n_889)
);

AOI22xp33_ASAP7_75t_L g890 ( 
.A1(n_699),
.A2(n_279),
.B1(n_341),
.B2(n_336),
.Y(n_890)
);

INVx1_ASAP7_75t_L g891 ( 
.A(n_682),
.Y(n_891)
);

NOR2xp33_ASAP7_75t_L g892 ( 
.A(n_699),
.B(n_316),
.Y(n_892)
);

AND2x2_ASAP7_75t_L g893 ( 
.A(n_699),
.B(n_406),
.Y(n_893)
);

INVx1_ASAP7_75t_L g894 ( 
.A(n_685),
.Y(n_894)
);

NAND2xp5_ASAP7_75t_L g895 ( 
.A(n_685),
.B(n_224),
.Y(n_895)
);

INVx2_ASAP7_75t_L g896 ( 
.A(n_658),
.Y(n_896)
);

INVx1_ASAP7_75t_L g897 ( 
.A(n_689),
.Y(n_897)
);

NAND2xp5_ASAP7_75t_SL g898 ( 
.A(n_639),
.B(n_641),
.Y(n_898)
);

NAND2xp5_ASAP7_75t_L g899 ( 
.A(n_689),
.B(n_224),
.Y(n_899)
);

NAND2xp5_ASAP7_75t_SL g900 ( 
.A(n_639),
.B(n_225),
.Y(n_900)
);

NOR2xp33_ASAP7_75t_L g901 ( 
.A(n_833),
.B(n_603),
.Y(n_901)
);

CKINVDCx20_ASAP7_75t_R g902 ( 
.A(n_765),
.Y(n_902)
);

CKINVDCx5p33_ASAP7_75t_R g903 ( 
.A(n_815),
.Y(n_903)
);

BUFx3_ASAP7_75t_L g904 ( 
.A(n_815),
.Y(n_904)
);

INVx1_ASAP7_75t_L g905 ( 
.A(n_734),
.Y(n_905)
);

BUFx2_ASAP7_75t_L g906 ( 
.A(n_803),
.Y(n_906)
);

BUFx6f_ASAP7_75t_L g907 ( 
.A(n_751),
.Y(n_907)
);

NOR2xp33_ASAP7_75t_L g908 ( 
.A(n_775),
.B(n_603),
.Y(n_908)
);

NAND2xp5_ASAP7_75t_L g909 ( 
.A(n_793),
.B(n_775),
.Y(n_909)
);

NAND2xp5_ASAP7_75t_L g910 ( 
.A(n_759),
.B(n_639),
.Y(n_910)
);

BUFx6f_ASAP7_75t_L g911 ( 
.A(n_751),
.Y(n_911)
);

INVx1_ASAP7_75t_SL g912 ( 
.A(n_751),
.Y(n_912)
);

BUFx6f_ASAP7_75t_SL g913 ( 
.A(n_825),
.Y(n_913)
);

INVx2_ASAP7_75t_SL g914 ( 
.A(n_739),
.Y(n_914)
);

NOR2x1p5_ASAP7_75t_L g915 ( 
.A(n_738),
.B(n_754),
.Y(n_915)
);

INVx1_ASAP7_75t_L g916 ( 
.A(n_734),
.Y(n_916)
);

NAND2xp5_ASAP7_75t_L g917 ( 
.A(n_759),
.B(n_742),
.Y(n_917)
);

NAND2xp5_ASAP7_75t_L g918 ( 
.A(n_744),
.B(n_641),
.Y(n_918)
);

INVx1_ASAP7_75t_L g919 ( 
.A(n_745),
.Y(n_919)
);

OR2x6_ASAP7_75t_L g920 ( 
.A(n_735),
.B(n_730),
.Y(n_920)
);

AOI22xp5_ASAP7_75t_L g921 ( 
.A1(n_877),
.A2(n_692),
.B1(n_727),
.B2(n_694),
.Y(n_921)
);

NAND2xp5_ASAP7_75t_L g922 ( 
.A(n_750),
.B(n_641),
.Y(n_922)
);

AND2x2_ASAP7_75t_L g923 ( 
.A(n_805),
.B(n_406),
.Y(n_923)
);

INVx1_ASAP7_75t_L g924 ( 
.A(n_762),
.Y(n_924)
);

INVx1_ASAP7_75t_L g925 ( 
.A(n_767),
.Y(n_925)
);

HB1xp67_ASAP7_75t_L g926 ( 
.A(n_804),
.Y(n_926)
);

AOI22xp33_ASAP7_75t_L g927 ( 
.A1(n_845),
.A2(n_670),
.B1(n_658),
.B2(n_666),
.Y(n_927)
);

NOR2xp33_ASAP7_75t_L g928 ( 
.A(n_766),
.B(n_603),
.Y(n_928)
);

INVx5_ASAP7_75t_L g929 ( 
.A(n_780),
.Y(n_929)
);

OAI22xp5_ASAP7_75t_SL g930 ( 
.A1(n_810),
.A2(n_318),
.B1(n_326),
.B2(n_327),
.Y(n_930)
);

AOI22xp33_ASAP7_75t_L g931 ( 
.A1(n_755),
.A2(n_677),
.B1(n_666),
.B2(n_669),
.Y(n_931)
);

OAI22xp5_ASAP7_75t_L g932 ( 
.A1(n_835),
.A2(n_636),
.B1(n_603),
.B2(n_627),
.Y(n_932)
);

INVx5_ASAP7_75t_L g933 ( 
.A(n_780),
.Y(n_933)
);

BUFx6f_ASAP7_75t_L g934 ( 
.A(n_780),
.Y(n_934)
);

INVx2_ASAP7_75t_L g935 ( 
.A(n_807),
.Y(n_935)
);

AOI211xp5_ASAP7_75t_L g936 ( 
.A1(n_810),
.A2(n_323),
.B(n_325),
.C(n_328),
.Y(n_936)
);

INVx1_ASAP7_75t_L g937 ( 
.A(n_768),
.Y(n_937)
);

INVx2_ASAP7_75t_L g938 ( 
.A(n_807),
.Y(n_938)
);

AND2x4_ASAP7_75t_L g939 ( 
.A(n_799),
.B(n_648),
.Y(n_939)
);

BUFx6f_ASAP7_75t_L g940 ( 
.A(n_780),
.Y(n_940)
);

INVx5_ASAP7_75t_L g941 ( 
.A(n_787),
.Y(n_941)
);

NAND2xp33_ASAP7_75t_L g942 ( 
.A(n_770),
.B(n_627),
.Y(n_942)
);

NOR2xp33_ASAP7_75t_L g943 ( 
.A(n_766),
.B(n_627),
.Y(n_943)
);

INVx1_ASAP7_75t_L g944 ( 
.A(n_769),
.Y(n_944)
);

INVx3_ASAP7_75t_L g945 ( 
.A(n_787),
.Y(n_945)
);

INVxp67_ASAP7_75t_SL g946 ( 
.A(n_787),
.Y(n_946)
);

AOI22xp5_ASAP7_75t_L g947 ( 
.A1(n_747),
.A2(n_692),
.B1(n_727),
.B2(n_694),
.Y(n_947)
);

INVx2_ASAP7_75t_L g948 ( 
.A(n_821),
.Y(n_948)
);

NAND2xp5_ASAP7_75t_L g949 ( 
.A(n_773),
.B(n_648),
.Y(n_949)
);

INVx2_ASAP7_75t_L g950 ( 
.A(n_821),
.Y(n_950)
);

NAND2xp5_ASAP7_75t_L g951 ( 
.A(n_778),
.B(n_648),
.Y(n_951)
);

NAND2xp5_ASAP7_75t_L g952 ( 
.A(n_779),
.B(n_651),
.Y(n_952)
);

O2A1O1Ixp33_ASAP7_75t_L g953 ( 
.A1(n_755),
.A2(n_695),
.B(n_703),
.C(n_723),
.Y(n_953)
);

NAND2x1p5_ASAP7_75t_L g954 ( 
.A(n_764),
.B(n_678),
.Y(n_954)
);

INVx5_ASAP7_75t_L g955 ( 
.A(n_787),
.Y(n_955)
);

INVx2_ASAP7_75t_L g956 ( 
.A(n_771),
.Y(n_956)
);

AND2x4_ASAP7_75t_L g957 ( 
.A(n_784),
.B(n_651),
.Y(n_957)
);

NAND2xp5_ASAP7_75t_SL g958 ( 
.A(n_732),
.B(n_678),
.Y(n_958)
);

NOR2xp33_ASAP7_75t_L g959 ( 
.A(n_874),
.B(n_627),
.Y(n_959)
);

INVx1_ASAP7_75t_L g960 ( 
.A(n_781),
.Y(n_960)
);

AOI22xp33_ASAP7_75t_L g961 ( 
.A1(n_844),
.A2(n_669),
.B1(n_670),
.B2(n_674),
.Y(n_961)
);

INVx1_ASAP7_75t_L g962 ( 
.A(n_801),
.Y(n_962)
);

NOR2xp33_ASAP7_75t_L g963 ( 
.A(n_732),
.B(n_636),
.Y(n_963)
);

OAI21xp5_ASAP7_75t_L g964 ( 
.A1(n_892),
.A2(n_703),
.B(n_695),
.Y(n_964)
);

NOR2xp67_ASAP7_75t_L g965 ( 
.A(n_830),
.B(n_636),
.Y(n_965)
);

CKINVDCx5p33_ASAP7_75t_R g966 ( 
.A(n_789),
.Y(n_966)
);

NAND3xp33_ASAP7_75t_SL g967 ( 
.A(n_841),
.B(n_800),
.C(n_772),
.Y(n_967)
);

O2A1O1Ixp33_ASAP7_75t_L g968 ( 
.A1(n_816),
.A2(n_707),
.B(n_712),
.C(n_723),
.Y(n_968)
);

INVx1_ASAP7_75t_L g969 ( 
.A(n_809),
.Y(n_969)
);

AND2x4_ASAP7_75t_L g970 ( 
.A(n_784),
.B(n_850),
.Y(n_970)
);

AND2x6_ASAP7_75t_SL g971 ( 
.A(n_819),
.B(n_408),
.Y(n_971)
);

BUFx4f_ASAP7_75t_L g972 ( 
.A(n_853),
.Y(n_972)
);

INVx4_ASAP7_75t_L g973 ( 
.A(n_789),
.Y(n_973)
);

INVx1_ASAP7_75t_L g974 ( 
.A(n_811),
.Y(n_974)
);

BUFx8_ASAP7_75t_L g975 ( 
.A(n_875),
.Y(n_975)
);

NOR2xp33_ASAP7_75t_L g976 ( 
.A(n_772),
.B(n_636),
.Y(n_976)
);

INVx1_ASAP7_75t_L g977 ( 
.A(n_818),
.Y(n_977)
);

INVx2_ASAP7_75t_L g978 ( 
.A(n_774),
.Y(n_978)
);

BUFx3_ASAP7_75t_L g979 ( 
.A(n_840),
.Y(n_979)
);

NAND2xp5_ASAP7_75t_L g980 ( 
.A(n_820),
.B(n_651),
.Y(n_980)
);

NAND2xp5_ASAP7_75t_L g981 ( 
.A(n_829),
.B(n_652),
.Y(n_981)
);

BUFx3_ASAP7_75t_L g982 ( 
.A(n_881),
.Y(n_982)
);

INVx1_ASAP7_75t_L g983 ( 
.A(n_831),
.Y(n_983)
);

INVx2_ASAP7_75t_L g984 ( 
.A(n_814),
.Y(n_984)
);

NAND2xp5_ASAP7_75t_SL g985 ( 
.A(n_764),
.B(n_678),
.Y(n_985)
);

NAND2xp33_ASAP7_75t_L g986 ( 
.A(n_770),
.B(n_848),
.Y(n_986)
);

INVx2_ASAP7_75t_L g987 ( 
.A(n_814),
.Y(n_987)
);

INVx1_ASAP7_75t_L g988 ( 
.A(n_827),
.Y(n_988)
);

NAND2x1p5_ASAP7_75t_L g989 ( 
.A(n_747),
.B(n_678),
.Y(n_989)
);

INVx2_ASAP7_75t_SL g990 ( 
.A(n_860),
.Y(n_990)
);

INVx1_ASAP7_75t_L g991 ( 
.A(n_836),
.Y(n_991)
);

NAND2xp5_ASAP7_75t_L g992 ( 
.A(n_736),
.B(n_652),
.Y(n_992)
);

NAND2xp5_ASAP7_75t_SL g993 ( 
.A(n_834),
.B(n_678),
.Y(n_993)
);

INVx2_ASAP7_75t_SL g994 ( 
.A(n_794),
.Y(n_994)
);

NAND2xp5_ASAP7_75t_L g995 ( 
.A(n_733),
.B(n_652),
.Y(n_995)
);

NAND2xp5_ASAP7_75t_L g996 ( 
.A(n_893),
.B(n_655),
.Y(n_996)
);

INVx1_ASAP7_75t_L g997 ( 
.A(n_847),
.Y(n_997)
);

BUFx6f_ASAP7_75t_L g998 ( 
.A(n_798),
.Y(n_998)
);

INVx1_ASAP7_75t_L g999 ( 
.A(n_849),
.Y(n_999)
);

INVx2_ASAP7_75t_L g1000 ( 
.A(n_817),
.Y(n_1000)
);

INVx1_ASAP7_75t_L g1001 ( 
.A(n_854),
.Y(n_1001)
);

BUFx2_ASAP7_75t_L g1002 ( 
.A(n_844),
.Y(n_1002)
);

AOI22xp33_ASAP7_75t_L g1003 ( 
.A1(n_844),
.A2(n_680),
.B1(n_674),
.B2(n_677),
.Y(n_1003)
);

AOI22xp33_ASAP7_75t_L g1004 ( 
.A1(n_861),
.A2(n_681),
.B1(n_680),
.B2(n_687),
.Y(n_1004)
);

BUFx6f_ASAP7_75t_L g1005 ( 
.A(n_798),
.Y(n_1005)
);

NAND2xp5_ASAP7_75t_L g1006 ( 
.A(n_835),
.B(n_655),
.Y(n_1006)
);

NOR2xp33_ASAP7_75t_L g1007 ( 
.A(n_795),
.B(n_707),
.Y(n_1007)
);

AOI22xp5_ASAP7_75t_L g1008 ( 
.A1(n_851),
.A2(n_714),
.B1(n_712),
.B2(n_719),
.Y(n_1008)
);

NAND2xp5_ASAP7_75t_L g1009 ( 
.A(n_796),
.B(n_655),
.Y(n_1009)
);

NAND2xp5_ASAP7_75t_SL g1010 ( 
.A(n_819),
.B(n_656),
.Y(n_1010)
);

INVx2_ASAP7_75t_SL g1011 ( 
.A(n_869),
.Y(n_1011)
);

HB1xp67_ASAP7_75t_L g1012 ( 
.A(n_752),
.Y(n_1012)
);

INVx1_ASAP7_75t_L g1013 ( 
.A(n_813),
.Y(n_1013)
);

INVx3_ASAP7_75t_L g1014 ( 
.A(n_859),
.Y(n_1014)
);

INVx1_ASAP7_75t_L g1015 ( 
.A(n_852),
.Y(n_1015)
);

INVx3_ASAP7_75t_L g1016 ( 
.A(n_859),
.Y(n_1016)
);

NAND2xp5_ASAP7_75t_L g1017 ( 
.A(n_749),
.B(n_656),
.Y(n_1017)
);

INVx3_ASAP7_75t_L g1018 ( 
.A(n_872),
.Y(n_1018)
);

AOI21x1_ASAP7_75t_L g1019 ( 
.A1(n_898),
.A2(n_719),
.B(n_714),
.Y(n_1019)
);

AND2x2_ASAP7_75t_L g1020 ( 
.A(n_851),
.B(n_408),
.Y(n_1020)
);

INVx1_ASAP7_75t_L g1021 ( 
.A(n_855),
.Y(n_1021)
);

HB1xp67_ASAP7_75t_L g1022 ( 
.A(n_752),
.Y(n_1022)
);

INVx2_ASAP7_75t_L g1023 ( 
.A(n_896),
.Y(n_1023)
);

AND2x2_ASAP7_75t_L g1024 ( 
.A(n_863),
.B(n_412),
.Y(n_1024)
);

NAND2xp5_ASAP7_75t_SL g1025 ( 
.A(n_783),
.B(n_795),
.Y(n_1025)
);

AND2x2_ASAP7_75t_L g1026 ( 
.A(n_867),
.B(n_412),
.Y(n_1026)
);

INVx2_ASAP7_75t_L g1027 ( 
.A(n_896),
.Y(n_1027)
);

BUFx6f_ASAP7_75t_L g1028 ( 
.A(n_788),
.Y(n_1028)
);

HB1xp67_ASAP7_75t_L g1029 ( 
.A(n_752),
.Y(n_1029)
);

INVxp67_ASAP7_75t_L g1030 ( 
.A(n_802),
.Y(n_1030)
);

INVx1_ASAP7_75t_L g1031 ( 
.A(n_873),
.Y(n_1031)
);

NAND2xp5_ASAP7_75t_L g1032 ( 
.A(n_822),
.B(n_656),
.Y(n_1032)
);

AND2x6_ASAP7_75t_SL g1033 ( 
.A(n_802),
.B(n_892),
.Y(n_1033)
);

INVx1_ASAP7_75t_L g1034 ( 
.A(n_882),
.Y(n_1034)
);

AOI22xp5_ASAP7_75t_L g1035 ( 
.A1(n_737),
.A2(n_730),
.B1(n_726),
.B2(n_721),
.Y(n_1035)
);

INVx4_ASAP7_75t_L g1036 ( 
.A(n_875),
.Y(n_1036)
);

NAND2xp33_ASAP7_75t_SL g1037 ( 
.A(n_786),
.B(n_693),
.Y(n_1037)
);

INVx1_ASAP7_75t_SL g1038 ( 
.A(n_758),
.Y(n_1038)
);

OAI22xp33_ASAP7_75t_L g1039 ( 
.A1(n_741),
.A2(n_730),
.B1(n_726),
.B2(n_721),
.Y(n_1039)
);

INVx1_ASAP7_75t_L g1040 ( 
.A(n_891),
.Y(n_1040)
);

NAND2xp5_ASAP7_75t_L g1041 ( 
.A(n_843),
.B(n_693),
.Y(n_1041)
);

OAI21xp33_ASAP7_75t_L g1042 ( 
.A1(n_748),
.A2(n_226),
.B(n_225),
.Y(n_1042)
);

AO22x1_ASAP7_75t_L g1043 ( 
.A1(n_823),
.A2(n_232),
.B1(n_300),
.B2(n_247),
.Y(n_1043)
);

BUFx4f_ASAP7_75t_L g1044 ( 
.A(n_758),
.Y(n_1044)
);

NAND2xp5_ASAP7_75t_L g1045 ( 
.A(n_843),
.B(n_693),
.Y(n_1045)
);

INVx2_ASAP7_75t_SL g1046 ( 
.A(n_735),
.Y(n_1046)
);

BUFx8_ASAP7_75t_L g1047 ( 
.A(n_806),
.Y(n_1047)
);

NAND2xp5_ASAP7_75t_L g1048 ( 
.A(n_872),
.B(n_706),
.Y(n_1048)
);

NOR2xp33_ASAP7_75t_L g1049 ( 
.A(n_786),
.B(n_681),
.Y(n_1049)
);

NAND2xp5_ASAP7_75t_L g1050 ( 
.A(n_857),
.B(n_706),
.Y(n_1050)
);

AOI22xp5_ASAP7_75t_L g1051 ( 
.A1(n_737),
.A2(n_726),
.B1(n_721),
.B2(n_718),
.Y(n_1051)
);

NAND2xp5_ASAP7_75t_SL g1052 ( 
.A(n_839),
.B(n_710),
.Y(n_1052)
);

INVx3_ASAP7_75t_L g1053 ( 
.A(n_743),
.Y(n_1053)
);

INVx1_ASAP7_75t_L g1054 ( 
.A(n_894),
.Y(n_1054)
);

INVx8_ASAP7_75t_L g1055 ( 
.A(n_746),
.Y(n_1055)
);

OAI21xp5_ASAP7_75t_L g1056 ( 
.A1(n_864),
.A2(n_715),
.B(n_710),
.Y(n_1056)
);

INVx4_ASAP7_75t_L g1057 ( 
.A(n_756),
.Y(n_1057)
);

OR2x6_ASAP7_75t_L g1058 ( 
.A(n_753),
.B(n_718),
.Y(n_1058)
);

NAND2xp5_ASAP7_75t_L g1059 ( 
.A(n_797),
.B(n_710),
.Y(n_1059)
);

NOR2x1_ASAP7_75t_L g1060 ( 
.A(n_828),
.B(n_715),
.Y(n_1060)
);

NAND2xp5_ASAP7_75t_SL g1061 ( 
.A(n_753),
.B(n_715),
.Y(n_1061)
);

INVx2_ASAP7_75t_SL g1062 ( 
.A(n_842),
.Y(n_1062)
);

OAI22xp33_ASAP7_75t_L g1063 ( 
.A1(n_868),
.A2(n_718),
.B1(n_717),
.B2(n_716),
.Y(n_1063)
);

INVx1_ASAP7_75t_L g1064 ( 
.A(n_897),
.Y(n_1064)
);

INVx2_ASAP7_75t_L g1065 ( 
.A(n_871),
.Y(n_1065)
);

NAND2xp5_ASAP7_75t_SL g1066 ( 
.A(n_865),
.B(n_716),
.Y(n_1066)
);

INVx2_ASAP7_75t_SL g1067 ( 
.A(n_842),
.Y(n_1067)
);

AOI22xp33_ASAP7_75t_L g1068 ( 
.A1(n_865),
.A2(n_687),
.B1(n_717),
.B2(n_716),
.Y(n_1068)
);

INVx3_ASAP7_75t_SL g1069 ( 
.A(n_866),
.Y(n_1069)
);

CKINVDCx5p33_ASAP7_75t_R g1070 ( 
.A(n_890),
.Y(n_1070)
);

A2O1A1Ixp33_ASAP7_75t_L g1071 ( 
.A1(n_884),
.A2(n_717),
.B(n_635),
.C(n_630),
.Y(n_1071)
);

OR2x6_ASAP7_75t_L g1072 ( 
.A(n_760),
.B(n_413),
.Y(n_1072)
);

INVx2_ASAP7_75t_L g1073 ( 
.A(n_876),
.Y(n_1073)
);

INVx1_ASAP7_75t_L g1074 ( 
.A(n_757),
.Y(n_1074)
);

NAND2xp5_ASAP7_75t_L g1075 ( 
.A(n_808),
.B(n_594),
.Y(n_1075)
);

NAND2xp5_ASAP7_75t_L g1076 ( 
.A(n_808),
.B(n_594),
.Y(n_1076)
);

AND2x4_ASAP7_75t_L g1077 ( 
.A(n_763),
.B(n_413),
.Y(n_1077)
);

INVx1_ASAP7_75t_L g1078 ( 
.A(n_761),
.Y(n_1078)
);

NAND2xp33_ASAP7_75t_L g1079 ( 
.A(n_770),
.B(n_594),
.Y(n_1079)
);

HB1xp67_ASAP7_75t_L g1080 ( 
.A(n_870),
.Y(n_1080)
);

INVx3_ASAP7_75t_L g1081 ( 
.A(n_782),
.Y(n_1081)
);

INVx2_ASAP7_75t_SL g1082 ( 
.A(n_846),
.Y(n_1082)
);

AOI22xp5_ASAP7_75t_L g1083 ( 
.A1(n_740),
.A2(n_635),
.B1(n_630),
.B2(n_626),
.Y(n_1083)
);

INVx1_ASAP7_75t_L g1084 ( 
.A(n_776),
.Y(n_1084)
);

INVx3_ASAP7_75t_L g1085 ( 
.A(n_785),
.Y(n_1085)
);

NAND2xp5_ASAP7_75t_L g1086 ( 
.A(n_812),
.B(n_599),
.Y(n_1086)
);

INVx2_ASAP7_75t_SL g1087 ( 
.A(n_846),
.Y(n_1087)
);

AOI22xp33_ASAP7_75t_L g1088 ( 
.A1(n_1070),
.A2(n_890),
.B1(n_824),
.B2(n_856),
.Y(n_1088)
);

NAND2x1_ASAP7_75t_L g1089 ( 
.A(n_1014),
.B(n_599),
.Y(n_1089)
);

OAI22xp5_ASAP7_75t_L g1090 ( 
.A1(n_909),
.A2(n_884),
.B1(n_777),
.B2(n_889),
.Y(n_1090)
);

NAND2xp5_ASAP7_75t_SL g1091 ( 
.A(n_903),
.B(n_770),
.Y(n_1091)
);

NAND2xp5_ASAP7_75t_L g1092 ( 
.A(n_917),
.B(n_791),
.Y(n_1092)
);

O2A1O1Ixp33_ASAP7_75t_L g1093 ( 
.A1(n_967),
.A2(n_864),
.B(n_856),
.C(n_866),
.Y(n_1093)
);

BUFx3_ASAP7_75t_L g1094 ( 
.A(n_904),
.Y(n_1094)
);

INVx2_ASAP7_75t_L g1095 ( 
.A(n_956),
.Y(n_1095)
);

NAND2xp5_ASAP7_75t_SL g1096 ( 
.A(n_907),
.B(n_770),
.Y(n_1096)
);

INVxp67_ASAP7_75t_SL g1097 ( 
.A(n_986),
.Y(n_1097)
);

AND2x2_ASAP7_75t_L g1098 ( 
.A(n_972),
.B(n_414),
.Y(n_1098)
);

NAND2xp5_ASAP7_75t_L g1099 ( 
.A(n_917),
.B(n_812),
.Y(n_1099)
);

INVx1_ASAP7_75t_L g1100 ( 
.A(n_919),
.Y(n_1100)
);

BUFx2_ASAP7_75t_L g1101 ( 
.A(n_906),
.Y(n_1101)
);

NOR2xp33_ASAP7_75t_L g1102 ( 
.A(n_1030),
.B(n_792),
.Y(n_1102)
);

AOI21xp5_ASAP7_75t_L g1103 ( 
.A1(n_1079),
.A2(n_790),
.B(n_878),
.Y(n_1103)
);

AOI21xp5_ASAP7_75t_L g1104 ( 
.A1(n_908),
.A2(n_790),
.B(n_880),
.Y(n_1104)
);

NAND3xp33_ASAP7_75t_SL g1105 ( 
.A(n_936),
.B(n_232),
.C(n_226),
.Y(n_1105)
);

BUFx6f_ASAP7_75t_L g1106 ( 
.A(n_907),
.Y(n_1106)
);

AOI21xp5_ASAP7_75t_L g1107 ( 
.A1(n_942),
.A2(n_910),
.B(n_964),
.Y(n_1107)
);

NAND2xp5_ASAP7_75t_SL g1108 ( 
.A(n_907),
.B(n_883),
.Y(n_1108)
);

A2O1A1Ixp33_ASAP7_75t_L g1109 ( 
.A1(n_967),
.A2(n_879),
.B(n_888),
.C(n_887),
.Y(n_1109)
);

A2O1A1Ixp33_ASAP7_75t_L g1110 ( 
.A1(n_1007),
.A2(n_963),
.B(n_1030),
.C(n_1025),
.Y(n_1110)
);

NAND2xp5_ASAP7_75t_L g1111 ( 
.A(n_994),
.B(n_885),
.Y(n_1111)
);

BUFx6f_ASAP7_75t_L g1112 ( 
.A(n_911),
.Y(n_1112)
);

INVx1_ASAP7_75t_L g1113 ( 
.A(n_924),
.Y(n_1113)
);

OR2x2_ASAP7_75t_L g1114 ( 
.A(n_990),
.B(n_895),
.Y(n_1114)
);

INVx6_ASAP7_75t_L g1115 ( 
.A(n_975),
.Y(n_1115)
);

AND2x2_ASAP7_75t_L g1116 ( 
.A(n_923),
.B(n_926),
.Y(n_1116)
);

INVx2_ASAP7_75t_L g1117 ( 
.A(n_978),
.Y(n_1117)
);

NAND2xp5_ASAP7_75t_L g1118 ( 
.A(n_1020),
.B(n_858),
.Y(n_1118)
);

OAI22xp5_ASAP7_75t_L g1119 ( 
.A1(n_988),
.A2(n_991),
.B1(n_910),
.B2(n_997),
.Y(n_1119)
);

INVx1_ASAP7_75t_L g1120 ( 
.A(n_925),
.Y(n_1120)
);

AOI21xp5_ASAP7_75t_L g1121 ( 
.A1(n_964),
.A2(n_862),
.B(n_886),
.Y(n_1121)
);

NOR2xp33_ASAP7_75t_SL g1122 ( 
.A(n_979),
.B(n_279),
.Y(n_1122)
);

INVx3_ASAP7_75t_L g1123 ( 
.A(n_911),
.Y(n_1123)
);

O2A1O1Ixp33_ASAP7_75t_L g1124 ( 
.A1(n_1042),
.A2(n_837),
.B(n_826),
.C(n_792),
.Y(n_1124)
);

NOR2xp33_ASAP7_75t_L g1125 ( 
.A(n_971),
.B(n_826),
.Y(n_1125)
);

INVx3_ASAP7_75t_L g1126 ( 
.A(n_911),
.Y(n_1126)
);

NOR2xp33_ASAP7_75t_SL g1127 ( 
.A(n_973),
.B(n_241),
.Y(n_1127)
);

AND2x2_ASAP7_75t_L g1128 ( 
.A(n_970),
.B(n_416),
.Y(n_1128)
);

BUFx6f_ASAP7_75t_L g1129 ( 
.A(n_934),
.Y(n_1129)
);

NAND2xp5_ASAP7_75t_SL g1130 ( 
.A(n_912),
.B(n_899),
.Y(n_1130)
);

OAI22xp5_ASAP7_75t_L g1131 ( 
.A1(n_999),
.A2(n_837),
.B1(n_900),
.B2(n_898),
.Y(n_1131)
);

OAI22xp5_ASAP7_75t_L g1132 ( 
.A1(n_1001),
.A2(n_900),
.B1(n_635),
.B2(n_630),
.Y(n_1132)
);

NAND2xp5_ASAP7_75t_L g1133 ( 
.A(n_1026),
.B(n_599),
.Y(n_1133)
);

O2A1O1Ixp33_ASAP7_75t_L g1134 ( 
.A1(n_901),
.A2(n_838),
.B(n_832),
.C(n_370),
.Y(n_1134)
);

INVx2_ASAP7_75t_L g1135 ( 
.A(n_984),
.Y(n_1135)
);

NAND3xp33_ASAP7_75t_SL g1136 ( 
.A(n_902),
.B(n_244),
.C(n_247),
.Y(n_1136)
);

CKINVDCx5p33_ASAP7_75t_R g1137 ( 
.A(n_975),
.Y(n_1137)
);

AOI21xp5_ASAP7_75t_L g1138 ( 
.A1(n_1059),
.A2(n_626),
.B(n_622),
.Y(n_1138)
);

BUFx6f_ASAP7_75t_L g1139 ( 
.A(n_934),
.Y(n_1139)
);

NOR2xp33_ASAP7_75t_L g1140 ( 
.A(n_914),
.B(n_602),
.Y(n_1140)
);

INVxp67_ASAP7_75t_L g1141 ( 
.A(n_913),
.Y(n_1141)
);

NOR2xp33_ASAP7_75t_L g1142 ( 
.A(n_1033),
.B(n_602),
.Y(n_1142)
);

INVx1_ASAP7_75t_L g1143 ( 
.A(n_937),
.Y(n_1143)
);

NAND2xp5_ASAP7_75t_L g1144 ( 
.A(n_1024),
.B(n_602),
.Y(n_1144)
);

O2A1O1Ixp33_ASAP7_75t_L g1145 ( 
.A1(n_1031),
.A2(n_357),
.B(n_293),
.C(n_294),
.Y(n_1145)
);

AND2x4_ASAP7_75t_L g1146 ( 
.A(n_912),
.B(n_619),
.Y(n_1146)
);

AND2x2_ASAP7_75t_L g1147 ( 
.A(n_905),
.B(n_418),
.Y(n_1147)
);

NAND2xp5_ASAP7_75t_L g1148 ( 
.A(n_916),
.B(n_619),
.Y(n_1148)
);

NAND2xp33_ASAP7_75t_SL g1149 ( 
.A(n_1069),
.B(n_626),
.Y(n_1149)
);

HB1xp67_ASAP7_75t_L g1150 ( 
.A(n_913),
.Y(n_1150)
);

AOI21xp5_ASAP7_75t_L g1151 ( 
.A1(n_1059),
.A2(n_622),
.B(n_620),
.Y(n_1151)
);

CKINVDCx5p33_ASAP7_75t_R g1152 ( 
.A(n_966),
.Y(n_1152)
);

BUFx6f_ASAP7_75t_L g1153 ( 
.A(n_934),
.Y(n_1153)
);

NAND2xp5_ASAP7_75t_L g1154 ( 
.A(n_944),
.B(n_619),
.Y(n_1154)
);

AO32x1_ASAP7_75t_L g1155 ( 
.A1(n_932),
.A2(n_426),
.A3(n_420),
.B1(n_419),
.B2(n_418),
.Y(n_1155)
);

NOR3xp33_ASAP7_75t_SL g1156 ( 
.A(n_930),
.B(n_366),
.C(n_241),
.Y(n_1156)
);

INVx1_ASAP7_75t_L g1157 ( 
.A(n_960),
.Y(n_1157)
);

OR2x6_ASAP7_75t_L g1158 ( 
.A(n_1055),
.B(n_622),
.Y(n_1158)
);

O2A1O1Ixp33_ASAP7_75t_L g1159 ( 
.A1(n_1034),
.A2(n_340),
.B(n_305),
.C(n_308),
.Y(n_1159)
);

BUFx8_ASAP7_75t_L g1160 ( 
.A(n_982),
.Y(n_1160)
);

A2O1A1Ixp33_ASAP7_75t_L g1161 ( 
.A1(n_928),
.A2(n_620),
.B(n_362),
.C(n_314),
.Y(n_1161)
);

BUFx6f_ASAP7_75t_L g1162 ( 
.A(n_940),
.Y(n_1162)
);

OAI21x1_ASAP7_75t_L g1163 ( 
.A1(n_1019),
.A2(n_1056),
.B(n_932),
.Y(n_1163)
);

AOI33xp33_ASAP7_75t_L g1164 ( 
.A1(n_962),
.A2(n_426),
.A3(n_420),
.B1(n_419),
.B2(n_337),
.B3(n_339),
.Y(n_1164)
);

A2O1A1Ixp33_ASAP7_75t_SL g1165 ( 
.A1(n_976),
.A2(n_620),
.B(n_384),
.C(n_381),
.Y(n_1165)
);

INVx2_ASAP7_75t_SL g1166 ( 
.A(n_1047),
.Y(n_1166)
);

CKINVDCx5p33_ASAP7_75t_R g1167 ( 
.A(n_973),
.Y(n_1167)
);

NOR2xp67_ASAP7_75t_L g1168 ( 
.A(n_929),
.B(n_933),
.Y(n_1168)
);

INVx1_ASAP7_75t_L g1169 ( 
.A(n_969),
.Y(n_1169)
);

A2O1A1Ixp33_ASAP7_75t_L g1170 ( 
.A1(n_943),
.A2(n_289),
.B(n_331),
.C(n_378),
.Y(n_1170)
);

AND2x2_ASAP7_75t_L g1171 ( 
.A(n_1002),
.B(n_0),
.Y(n_1171)
);

INVx5_ASAP7_75t_L g1172 ( 
.A(n_1036),
.Y(n_1172)
);

INVx1_ASAP7_75t_L g1173 ( 
.A(n_974),
.Y(n_1173)
);

NAND2xp5_ASAP7_75t_SL g1174 ( 
.A(n_939),
.B(n_244),
.Y(n_1174)
);

NAND2xp5_ASAP7_75t_L g1175 ( 
.A(n_977),
.B(n_338),
.Y(n_1175)
);

INVx1_ASAP7_75t_L g1176 ( 
.A(n_983),
.Y(n_1176)
);

OAI22xp5_ASAP7_75t_L g1177 ( 
.A1(n_1040),
.A2(n_386),
.B1(n_383),
.B2(n_368),
.Y(n_1177)
);

AOI21xp5_ASAP7_75t_L g1178 ( 
.A1(n_1017),
.A2(n_335),
.B(n_271),
.Y(n_1178)
);

AOI21xp5_ASAP7_75t_L g1179 ( 
.A1(n_1017),
.A2(n_317),
.B(n_276),
.Y(n_1179)
);

NAND2xp5_ASAP7_75t_L g1180 ( 
.A(n_939),
.B(n_338),
.Y(n_1180)
);

BUFx6f_ASAP7_75t_L g1181 ( 
.A(n_940),
.Y(n_1181)
);

NOR2xp33_ASAP7_75t_SL g1182 ( 
.A(n_1036),
.B(n_342),
.Y(n_1182)
);

AOI21xp5_ASAP7_75t_L g1183 ( 
.A1(n_1032),
.A2(n_311),
.B(n_280),
.Y(n_1183)
);

NOR2xp33_ASAP7_75t_L g1184 ( 
.A(n_1055),
.B(n_342),
.Y(n_1184)
);

AOI21xp5_ASAP7_75t_L g1185 ( 
.A1(n_1032),
.A2(n_319),
.B(n_282),
.Y(n_1185)
);

BUFx6f_ASAP7_75t_L g1186 ( 
.A(n_940),
.Y(n_1186)
);

OAI22xp5_ASAP7_75t_L g1187 ( 
.A1(n_1054),
.A2(n_383),
.B1(n_368),
.B2(n_366),
.Y(n_1187)
);

NAND2xp5_ASAP7_75t_SL g1188 ( 
.A(n_929),
.B(n_347),
.Y(n_1188)
);

AOI22xp5_ASAP7_75t_L g1189 ( 
.A1(n_915),
.A2(n_364),
.B1(n_347),
.B2(n_358),
.Y(n_1189)
);

INVx1_ASAP7_75t_L g1190 ( 
.A(n_1064),
.Y(n_1190)
);

AND2x4_ASAP7_75t_L g1191 ( 
.A(n_929),
.B(n_933),
.Y(n_1191)
);

NAND2xp5_ASAP7_75t_SL g1192 ( 
.A(n_929),
.B(n_364),
.Y(n_1192)
);

OR2x6_ASAP7_75t_L g1193 ( 
.A(n_1055),
.B(n_200),
.Y(n_1193)
);

BUFx2_ASAP7_75t_SL g1194 ( 
.A(n_933),
.Y(n_1194)
);

NAND2xp5_ASAP7_75t_L g1195 ( 
.A(n_1074),
.B(n_2),
.Y(n_1195)
);

INVx3_ASAP7_75t_L g1196 ( 
.A(n_933),
.Y(n_1196)
);

INVx1_ASAP7_75t_L g1197 ( 
.A(n_1011),
.Y(n_1197)
);

BUFx3_ASAP7_75t_L g1198 ( 
.A(n_1077),
.Y(n_1198)
);

AOI21xp5_ASAP7_75t_L g1199 ( 
.A1(n_996),
.A2(n_333),
.B(n_329),
.Y(n_1199)
);

NAND2xp5_ASAP7_75t_L g1200 ( 
.A(n_1078),
.B(n_2),
.Y(n_1200)
);

NAND2xp5_ASAP7_75t_L g1201 ( 
.A(n_1084),
.B(n_5),
.Y(n_1201)
);

INVx1_ASAP7_75t_L g1202 ( 
.A(n_1077),
.Y(n_1202)
);

INVx4_ASAP7_75t_L g1203 ( 
.A(n_941),
.Y(n_1203)
);

BUFx6f_ASAP7_75t_L g1204 ( 
.A(n_941),
.Y(n_1204)
);

BUFx12f_ASAP7_75t_L g1205 ( 
.A(n_1062),
.Y(n_1205)
);

INVx5_ASAP7_75t_L g1206 ( 
.A(n_920),
.Y(n_1206)
);

O2A1O1Ixp5_ASAP7_75t_L g1207 ( 
.A1(n_1037),
.A2(n_6),
.B(n_8),
.C(n_9),
.Y(n_1207)
);

NAND2xp5_ASAP7_75t_L g1208 ( 
.A(n_959),
.B(n_8),
.Y(n_1208)
);

OAI22xp5_ASAP7_75t_L g1209 ( 
.A1(n_1044),
.A2(n_324),
.B1(n_322),
.B2(n_320),
.Y(n_1209)
);

AND2x2_ASAP7_75t_L g1210 ( 
.A(n_1072),
.B(n_9),
.Y(n_1210)
);

O2A1O1Ixp33_ASAP7_75t_L g1211 ( 
.A1(n_1067),
.A2(n_11),
.B(n_14),
.C(n_15),
.Y(n_1211)
);

AOI21xp5_ASAP7_75t_L g1212 ( 
.A1(n_996),
.A2(n_299),
.B(n_298),
.Y(n_1212)
);

AOI221xp5_ASAP7_75t_L g1213 ( 
.A1(n_1043),
.A2(n_283),
.B1(n_295),
.B2(n_291),
.C(n_287),
.Y(n_1213)
);

OAI22xp5_ASAP7_75t_L g1214 ( 
.A1(n_1044),
.A2(n_297),
.B1(n_249),
.B2(n_211),
.Y(n_1214)
);

O2A1O1Ixp33_ASAP7_75t_L g1215 ( 
.A1(n_1082),
.A2(n_11),
.B(n_17),
.C(n_18),
.Y(n_1215)
);

INVx6_ASAP7_75t_L g1216 ( 
.A(n_941),
.Y(n_1216)
);

INVx2_ASAP7_75t_SL g1217 ( 
.A(n_1087),
.Y(n_1217)
);

AOI21xp5_ASAP7_75t_L g1218 ( 
.A1(n_1050),
.A2(n_249),
.B(n_211),
.Y(n_1218)
);

BUFx6f_ASAP7_75t_L g1219 ( 
.A(n_941),
.Y(n_1219)
);

INVx3_ASAP7_75t_L g1220 ( 
.A(n_955),
.Y(n_1220)
);

CKINVDCx11_ASAP7_75t_R g1221 ( 
.A(n_1058),
.Y(n_1221)
);

OAI22xp5_ASAP7_75t_L g1222 ( 
.A1(n_918),
.A2(n_249),
.B1(n_211),
.B2(n_200),
.Y(n_1222)
);

O2A1O1Ixp33_ASAP7_75t_L g1223 ( 
.A1(n_968),
.A2(n_19),
.B(n_20),
.C(n_22),
.Y(n_1223)
);

OAI22xp5_ASAP7_75t_L g1224 ( 
.A1(n_918),
.A2(n_249),
.B1(n_211),
.B2(n_200),
.Y(n_1224)
);

INVx2_ASAP7_75t_L g1225 ( 
.A(n_987),
.Y(n_1225)
);

INVx1_ASAP7_75t_L g1226 ( 
.A(n_1013),
.Y(n_1226)
);

NAND2xp5_ASAP7_75t_L g1227 ( 
.A(n_1046),
.B(n_19),
.Y(n_1227)
);

AOI22xp5_ASAP7_75t_L g1228 ( 
.A1(n_1012),
.A2(n_211),
.B1(n_249),
.B2(n_25),
.Y(n_1228)
);

A2O1A1Ixp33_ASAP7_75t_L g1229 ( 
.A1(n_953),
.A2(n_20),
.B(n_22),
.C(n_27),
.Y(n_1229)
);

NOR2xp33_ASAP7_75t_L g1230 ( 
.A(n_1018),
.B(n_28),
.Y(n_1230)
);

OR2x6_ASAP7_75t_L g1231 ( 
.A(n_1022),
.B(n_28),
.Y(n_1231)
);

INVx5_ASAP7_75t_L g1232 ( 
.A(n_920),
.Y(n_1232)
);

O2A1O1Ixp33_ASAP7_75t_L g1233 ( 
.A1(n_968),
.A2(n_29),
.B(n_30),
.C(n_33),
.Y(n_1233)
);

NAND2xp5_ASAP7_75t_L g1234 ( 
.A(n_1038),
.B(n_33),
.Y(n_1234)
);

NOR2xp33_ASAP7_75t_L g1235 ( 
.A(n_1018),
.B(n_34),
.Y(n_1235)
);

OAI22xp5_ASAP7_75t_L g1236 ( 
.A1(n_922),
.A2(n_34),
.B1(n_35),
.B2(n_37),
.Y(n_1236)
);

NAND2xp5_ASAP7_75t_SL g1237 ( 
.A(n_955),
.B(n_38),
.Y(n_1237)
);

NAND2xp5_ASAP7_75t_L g1238 ( 
.A(n_1009),
.B(n_39),
.Y(n_1238)
);

OAI22xp5_ASAP7_75t_L g1239 ( 
.A1(n_1110),
.A2(n_1029),
.B1(n_952),
.B2(n_951),
.Y(n_1239)
);

AOI21xp5_ASAP7_75t_L g1240 ( 
.A1(n_1097),
.A2(n_1071),
.B(n_995),
.Y(n_1240)
);

NAND2xp5_ASAP7_75t_L g1241 ( 
.A(n_1116),
.B(n_965),
.Y(n_1241)
);

OR2x6_ASAP7_75t_L g1242 ( 
.A(n_1231),
.B(n_920),
.Y(n_1242)
);

NOR2xp33_ASAP7_75t_L g1243 ( 
.A(n_1125),
.B(n_1057),
.Y(n_1243)
);

AOI221xp5_ASAP7_75t_SL g1244 ( 
.A1(n_1223),
.A2(n_953),
.B1(n_1039),
.B2(n_952),
.C(n_951),
.Y(n_1244)
);

AO31x2_ASAP7_75t_L g1245 ( 
.A1(n_1107),
.A2(n_1041),
.A3(n_1045),
.B(n_1006),
.Y(n_1245)
);

NAND2xp5_ASAP7_75t_L g1246 ( 
.A(n_1128),
.B(n_1053),
.Y(n_1246)
);

OAI21x1_ASAP7_75t_L g1247 ( 
.A1(n_1138),
.A2(n_1056),
.B(n_1006),
.Y(n_1247)
);

AO21x2_ASAP7_75t_L g1248 ( 
.A1(n_1218),
.A2(n_1165),
.B(n_1163),
.Y(n_1248)
);

A2O1A1Ixp33_ASAP7_75t_L g1249 ( 
.A1(n_1102),
.A2(n_1049),
.B(n_921),
.C(n_958),
.Y(n_1249)
);

AOI21xp5_ASAP7_75t_SL g1250 ( 
.A1(n_1119),
.A2(n_1009),
.B(n_1041),
.Y(n_1250)
);

NAND2xp5_ASAP7_75t_L g1251 ( 
.A(n_1098),
.B(n_1081),
.Y(n_1251)
);

INVx1_ASAP7_75t_L g1252 ( 
.A(n_1100),
.Y(n_1252)
);

AOI21xp5_ASAP7_75t_L g1253 ( 
.A1(n_1092),
.A2(n_995),
.B(n_992),
.Y(n_1253)
);

AOI21xp5_ASAP7_75t_L g1254 ( 
.A1(n_1090),
.A2(n_980),
.B(n_949),
.Y(n_1254)
);

OAI21xp5_ASAP7_75t_L g1255 ( 
.A1(n_1099),
.A2(n_1010),
.B(n_947),
.Y(n_1255)
);

NAND2x1p5_ASAP7_75t_L g1256 ( 
.A(n_1094),
.B(n_1191),
.Y(n_1256)
);

AND2x2_ASAP7_75t_L g1257 ( 
.A(n_1171),
.B(n_957),
.Y(n_1257)
);

AOI21xp5_ASAP7_75t_L g1258 ( 
.A1(n_1121),
.A2(n_1104),
.B(n_1103),
.Y(n_1258)
);

BUFx3_ASAP7_75t_L g1259 ( 
.A(n_1160),
.Y(n_1259)
);

INVx2_ASAP7_75t_L g1260 ( 
.A(n_1117),
.Y(n_1260)
);

OAI21xp5_ASAP7_75t_L g1261 ( 
.A1(n_1109),
.A2(n_1086),
.B(n_1076),
.Y(n_1261)
);

AOI21xp5_ASAP7_75t_L g1262 ( 
.A1(n_1238),
.A2(n_980),
.B(n_949),
.Y(n_1262)
);

AOI21xp5_ASAP7_75t_L g1263 ( 
.A1(n_1118),
.A2(n_981),
.B(n_922),
.Y(n_1263)
);

NAND2xp5_ASAP7_75t_L g1264 ( 
.A(n_1198),
.B(n_1081),
.Y(n_1264)
);

INVx1_ASAP7_75t_L g1265 ( 
.A(n_1113),
.Y(n_1265)
);

AO21x1_ASAP7_75t_L g1266 ( 
.A1(n_1228),
.A2(n_1061),
.B(n_989),
.Y(n_1266)
);

AO31x2_ASAP7_75t_L g1267 ( 
.A1(n_1131),
.A2(n_1045),
.A3(n_1076),
.B(n_1075),
.Y(n_1267)
);

AO22x2_ASAP7_75t_L g1268 ( 
.A1(n_1202),
.A2(n_1021),
.B1(n_1015),
.B2(n_1027),
.Y(n_1268)
);

INVx1_ASAP7_75t_L g1269 ( 
.A(n_1120),
.Y(n_1269)
);

NAND3xp33_ASAP7_75t_L g1270 ( 
.A(n_1233),
.B(n_931),
.C(n_1008),
.Y(n_1270)
);

OAI22xp5_ASAP7_75t_L g1271 ( 
.A1(n_1189),
.A2(n_981),
.B1(n_1080),
.B2(n_927),
.Y(n_1271)
);

INVx1_ASAP7_75t_SL g1272 ( 
.A(n_1221),
.Y(n_1272)
);

OR2x6_ASAP7_75t_L g1273 ( 
.A(n_1231),
.B(n_957),
.Y(n_1273)
);

INVx1_ASAP7_75t_L g1274 ( 
.A(n_1143),
.Y(n_1274)
);

NAND2x1_ASAP7_75t_L g1275 ( 
.A(n_1203),
.B(n_945),
.Y(n_1275)
);

AND2x2_ASAP7_75t_L g1276 ( 
.A(n_1210),
.B(n_1085),
.Y(n_1276)
);

NAND2xp5_ASAP7_75t_L g1277 ( 
.A(n_1147),
.B(n_1085),
.Y(n_1277)
);

AOI21x1_ASAP7_75t_L g1278 ( 
.A1(n_1222),
.A2(n_1066),
.B(n_1086),
.Y(n_1278)
);

AOI21xp5_ASAP7_75t_L g1279 ( 
.A1(n_1124),
.A2(n_1048),
.B(n_985),
.Y(n_1279)
);

NAND2xp5_ASAP7_75t_L g1280 ( 
.A(n_1111),
.B(n_1073),
.Y(n_1280)
);

NAND2x1p5_ASAP7_75t_L g1281 ( 
.A(n_1172),
.B(n_955),
.Y(n_1281)
);

CKINVDCx20_ASAP7_75t_R g1282 ( 
.A(n_1137),
.Y(n_1282)
);

OAI21xp5_ASAP7_75t_SL g1283 ( 
.A1(n_1189),
.A2(n_1060),
.B(n_1003),
.Y(n_1283)
);

INVx1_ASAP7_75t_L g1284 ( 
.A(n_1157),
.Y(n_1284)
);

AOI21xp5_ASAP7_75t_L g1285 ( 
.A1(n_1134),
.A2(n_1048),
.B(n_1063),
.Y(n_1285)
);

AOI21xp5_ASAP7_75t_L g1286 ( 
.A1(n_1178),
.A2(n_993),
.B(n_946),
.Y(n_1286)
);

AOI21xp5_ASAP7_75t_L g1287 ( 
.A1(n_1208),
.A2(n_1016),
.B(n_1014),
.Y(n_1287)
);

OAI21x1_ASAP7_75t_L g1288 ( 
.A1(n_1132),
.A2(n_961),
.B(n_1051),
.Y(n_1288)
);

AOI21xp5_ASAP7_75t_L g1289 ( 
.A1(n_1091),
.A2(n_1016),
.B(n_1005),
.Y(n_1289)
);

OAI21x1_ASAP7_75t_SL g1290 ( 
.A1(n_1195),
.A2(n_935),
.B(n_938),
.Y(n_1290)
);

O2A1O1Ixp33_ASAP7_75t_SL g1291 ( 
.A1(n_1229),
.A2(n_1052),
.B(n_948),
.C(n_950),
.Y(n_1291)
);

AO31x2_ASAP7_75t_L g1292 ( 
.A1(n_1224),
.A2(n_1000),
.A3(n_1023),
.B(n_1065),
.Y(n_1292)
);

BUFx6f_ASAP7_75t_L g1293 ( 
.A(n_1204),
.Y(n_1293)
);

AOI21xp5_ASAP7_75t_L g1294 ( 
.A1(n_1096),
.A2(n_1005),
.B(n_998),
.Y(n_1294)
);

AOI21xp5_ASAP7_75t_SL g1295 ( 
.A1(n_1193),
.A2(n_1058),
.B(n_1028),
.Y(n_1295)
);

NAND2xp5_ASAP7_75t_L g1296 ( 
.A(n_1184),
.B(n_945),
.Y(n_1296)
);

AOI21xp5_ASAP7_75t_L g1297 ( 
.A1(n_1130),
.A2(n_1005),
.B(n_998),
.Y(n_1297)
);

O2A1O1Ixp5_ASAP7_75t_L g1298 ( 
.A1(n_1188),
.A2(n_955),
.B(n_1083),
.C(n_1035),
.Y(n_1298)
);

AOI21xp5_ASAP7_75t_L g1299 ( 
.A1(n_1089),
.A2(n_1155),
.B(n_1154),
.Y(n_1299)
);

BUFx4f_ASAP7_75t_L g1300 ( 
.A(n_1115),
.Y(n_1300)
);

NAND2xp5_ASAP7_75t_L g1301 ( 
.A(n_1169),
.B(n_1173),
.Y(n_1301)
);

OAI21xp5_ASAP7_75t_L g1302 ( 
.A1(n_1200),
.A2(n_1068),
.B(n_954),
.Y(n_1302)
);

AOI21xp5_ASAP7_75t_L g1303 ( 
.A1(n_1155),
.A2(n_998),
.B(n_954),
.Y(n_1303)
);

OAI21x1_ASAP7_75t_SL g1304 ( 
.A1(n_1201),
.A2(n_1004),
.B(n_1028),
.Y(n_1304)
);

CKINVDCx5p33_ASAP7_75t_R g1305 ( 
.A(n_1152),
.Y(n_1305)
);

INVx4_ASAP7_75t_L g1306 ( 
.A(n_1172),
.Y(n_1306)
);

NAND2xp5_ASAP7_75t_L g1307 ( 
.A(n_1176),
.B(n_1028),
.Y(n_1307)
);

OAI21x1_ASAP7_75t_L g1308 ( 
.A1(n_1108),
.A2(n_117),
.B(n_178),
.Y(n_1308)
);

OAI21x1_ASAP7_75t_L g1309 ( 
.A1(n_1196),
.A2(n_111),
.B(n_177),
.Y(n_1309)
);

OAI21x1_ASAP7_75t_L g1310 ( 
.A1(n_1196),
.A2(n_95),
.B(n_173),
.Y(n_1310)
);

AOI21xp33_ASAP7_75t_L g1311 ( 
.A1(n_1088),
.A2(n_1145),
.B(n_1159),
.Y(n_1311)
);

NAND3x1_ASAP7_75t_L g1312 ( 
.A(n_1142),
.B(n_1228),
.C(n_1227),
.Y(n_1312)
);

OAI21xp5_ASAP7_75t_L g1313 ( 
.A1(n_1161),
.A2(n_1207),
.B(n_1170),
.Y(n_1313)
);

AO32x2_ASAP7_75t_L g1314 ( 
.A1(n_1236),
.A2(n_40),
.A3(n_41),
.B1(n_43),
.B2(n_44),
.Y(n_1314)
);

OA21x2_ASAP7_75t_L g1315 ( 
.A1(n_1133),
.A2(n_1144),
.B(n_1135),
.Y(n_1315)
);

INVx1_ASAP7_75t_L g1316 ( 
.A(n_1190),
.Y(n_1316)
);

NOR2xp33_ASAP7_75t_L g1317 ( 
.A(n_1136),
.B(n_40),
.Y(n_1317)
);

AOI21xp5_ASAP7_75t_L g1318 ( 
.A1(n_1155),
.A2(n_130),
.B(n_165),
.Y(n_1318)
);

OAI21x1_ASAP7_75t_SL g1319 ( 
.A1(n_1148),
.A2(n_48),
.B(n_55),
.Y(n_1319)
);

INVx1_ASAP7_75t_L g1320 ( 
.A(n_1226),
.Y(n_1320)
);

AO31x2_ASAP7_75t_L g1321 ( 
.A1(n_1214),
.A2(n_123),
.A3(n_150),
.B(n_73),
.Y(n_1321)
);

A2O1A1Ixp33_ASAP7_75t_L g1322 ( 
.A1(n_1105),
.A2(n_48),
.B(n_60),
.C(n_88),
.Y(n_1322)
);

OR2x2_ASAP7_75t_L g1323 ( 
.A(n_1234),
.B(n_94),
.Y(n_1323)
);

AOI21x1_ASAP7_75t_L g1324 ( 
.A1(n_1179),
.A2(n_1185),
.B(n_1183),
.Y(n_1324)
);

INVx2_ASAP7_75t_L g1325 ( 
.A(n_1225),
.Y(n_1325)
);

AOI21xp5_ASAP7_75t_L g1326 ( 
.A1(n_1158),
.A2(n_131),
.B(n_138),
.Y(n_1326)
);

OR2x2_ASAP7_75t_L g1327 ( 
.A(n_1180),
.B(n_141),
.Y(n_1327)
);

BUFx6f_ASAP7_75t_L g1328 ( 
.A(n_1204),
.Y(n_1328)
);

INVx1_ASAP7_75t_SL g1329 ( 
.A(n_1146),
.Y(n_1329)
);

NOR2xp33_ASAP7_75t_L g1330 ( 
.A(n_1127),
.B(n_198),
.Y(n_1330)
);

CKINVDCx9p33_ASAP7_75t_R g1331 ( 
.A(n_1230),
.Y(n_1331)
);

NAND2xp5_ASAP7_75t_L g1332 ( 
.A(n_1217),
.B(n_1197),
.Y(n_1332)
);

AND2x2_ASAP7_75t_L g1333 ( 
.A(n_1231),
.B(n_1156),
.Y(n_1333)
);

OAI21x1_ASAP7_75t_L g1334 ( 
.A1(n_1220),
.A2(n_1168),
.B(n_1237),
.Y(n_1334)
);

AND2x4_ASAP7_75t_L g1335 ( 
.A(n_1158),
.B(n_1206),
.Y(n_1335)
);

OAI22xp5_ASAP7_75t_L g1336 ( 
.A1(n_1175),
.A2(n_1114),
.B1(n_1235),
.B2(n_1158),
.Y(n_1336)
);

AO31x2_ASAP7_75t_L g1337 ( 
.A1(n_1140),
.A2(n_1199),
.A3(n_1212),
.B(n_1209),
.Y(n_1337)
);

INVx1_ASAP7_75t_L g1338 ( 
.A(n_1164),
.Y(n_1338)
);

AOI21xp5_ASAP7_75t_L g1339 ( 
.A1(n_1168),
.A2(n_1193),
.B(n_1149),
.Y(n_1339)
);

CKINVDCx5p33_ASAP7_75t_R g1340 ( 
.A(n_1167),
.Y(n_1340)
);

INVx2_ASAP7_75t_SL g1341 ( 
.A(n_1166),
.Y(n_1341)
);

OAI21x1_ASAP7_75t_L g1342 ( 
.A1(n_1220),
.A2(n_1192),
.B(n_1123),
.Y(n_1342)
);

A2O1A1Ixp33_ASAP7_75t_L g1343 ( 
.A1(n_1211),
.A2(n_1215),
.B(n_1174),
.C(n_1146),
.Y(n_1343)
);

AND2x4_ASAP7_75t_L g1344 ( 
.A(n_1206),
.B(n_1232),
.Y(n_1344)
);

AO31x2_ASAP7_75t_L g1345 ( 
.A1(n_1177),
.A2(n_1187),
.A3(n_1203),
.B(n_1232),
.Y(n_1345)
);

OAI21x1_ASAP7_75t_L g1346 ( 
.A1(n_1123),
.A2(n_1126),
.B(n_1232),
.Y(n_1346)
);

NAND2xp5_ASAP7_75t_L g1347 ( 
.A(n_1122),
.B(n_1126),
.Y(n_1347)
);

BUFx6f_ASAP7_75t_L g1348 ( 
.A(n_1204),
.Y(n_1348)
);

INVx6_ASAP7_75t_L g1349 ( 
.A(n_1205),
.Y(n_1349)
);

INVxp67_ASAP7_75t_SL g1350 ( 
.A(n_1219),
.Y(n_1350)
);

NAND3x1_ASAP7_75t_L g1351 ( 
.A(n_1182),
.B(n_1213),
.C(n_1150),
.Y(n_1351)
);

O2A1O1Ixp33_ASAP7_75t_SL g1352 ( 
.A1(n_1141),
.A2(n_1194),
.B(n_1216),
.C(n_1219),
.Y(n_1352)
);

OAI21xp5_ASAP7_75t_L g1353 ( 
.A1(n_1193),
.A2(n_1206),
.B(n_1153),
.Y(n_1353)
);

INVx1_ASAP7_75t_L g1354 ( 
.A(n_1129),
.Y(n_1354)
);

OR2x2_ASAP7_75t_L g1355 ( 
.A(n_1106),
.B(n_1112),
.Y(n_1355)
);

NAND2xp5_ASAP7_75t_L g1356 ( 
.A(n_1106),
.B(n_1112),
.Y(n_1356)
);

OAI22xp5_ASAP7_75t_L g1357 ( 
.A1(n_1216),
.A2(n_1112),
.B1(n_1219),
.B2(n_1153),
.Y(n_1357)
);

AO21x2_ASAP7_75t_L g1358 ( 
.A1(n_1139),
.A2(n_1153),
.B(n_1162),
.Y(n_1358)
);

OAI21x1_ASAP7_75t_L g1359 ( 
.A1(n_1139),
.A2(n_1162),
.B(n_1181),
.Y(n_1359)
);

NAND2xp5_ASAP7_75t_L g1360 ( 
.A(n_1186),
.B(n_1162),
.Y(n_1360)
);

AND2x4_ASAP7_75t_L g1361 ( 
.A(n_1181),
.B(n_1186),
.Y(n_1361)
);

OAI21x1_ASAP7_75t_L g1362 ( 
.A1(n_1181),
.A2(n_1151),
.B(n_1138),
.Y(n_1362)
);

AOI21xp5_ASAP7_75t_L g1363 ( 
.A1(n_1186),
.A2(n_1097),
.B(n_986),
.Y(n_1363)
);

OAI22xp5_ASAP7_75t_L g1364 ( 
.A1(n_1110),
.A2(n_909),
.B1(n_917),
.B2(n_833),
.Y(n_1364)
);

OA21x2_ASAP7_75t_L g1365 ( 
.A1(n_1163),
.A2(n_1107),
.B(n_964),
.Y(n_1365)
);

OAI21xp5_ASAP7_75t_L g1366 ( 
.A1(n_1110),
.A2(n_909),
.B(n_1107),
.Y(n_1366)
);

AOI21xp5_ASAP7_75t_L g1367 ( 
.A1(n_1097),
.A2(n_986),
.B(n_909),
.Y(n_1367)
);

NAND2xp5_ASAP7_75t_L g1368 ( 
.A(n_1116),
.B(n_909),
.Y(n_1368)
);

AOI21x1_ASAP7_75t_L g1369 ( 
.A1(n_1107),
.A2(n_1218),
.B(n_1151),
.Y(n_1369)
);

BUFx2_ASAP7_75t_L g1370 ( 
.A(n_1101),
.Y(n_1370)
);

INVx1_ASAP7_75t_L g1371 ( 
.A(n_1100),
.Y(n_1371)
);

OAI21x1_ASAP7_75t_SL g1372 ( 
.A1(n_1119),
.A2(n_1093),
.B(n_953),
.Y(n_1372)
);

NAND2xp5_ASAP7_75t_L g1373 ( 
.A(n_1116),
.B(n_909),
.Y(n_1373)
);

AO32x2_ASAP7_75t_L g1374 ( 
.A1(n_1119),
.A2(n_1236),
.A3(n_1131),
.B1(n_1090),
.B2(n_990),
.Y(n_1374)
);

OAI21x1_ASAP7_75t_L g1375 ( 
.A1(n_1138),
.A2(n_1151),
.B(n_1163),
.Y(n_1375)
);

OAI21xp5_ASAP7_75t_L g1376 ( 
.A1(n_1110),
.A2(n_909),
.B(n_1107),
.Y(n_1376)
);

INVx1_ASAP7_75t_L g1377 ( 
.A(n_1100),
.Y(n_1377)
);

OAI22xp5_ASAP7_75t_L g1378 ( 
.A1(n_1110),
.A2(n_909),
.B1(n_917),
.B2(n_833),
.Y(n_1378)
);

AOI21xp5_ASAP7_75t_L g1379 ( 
.A1(n_1097),
.A2(n_986),
.B(n_909),
.Y(n_1379)
);

OAI21x1_ASAP7_75t_L g1380 ( 
.A1(n_1138),
.A2(n_1151),
.B(n_1163),
.Y(n_1380)
);

INVx4_ASAP7_75t_L g1381 ( 
.A(n_1172),
.Y(n_1381)
);

NAND2xp5_ASAP7_75t_L g1382 ( 
.A(n_1116),
.B(n_909),
.Y(n_1382)
);

OAI21x1_ASAP7_75t_L g1383 ( 
.A1(n_1138),
.A2(n_1151),
.B(n_1163),
.Y(n_1383)
);

INVx2_ASAP7_75t_L g1384 ( 
.A(n_1095),
.Y(n_1384)
);

NAND2xp5_ASAP7_75t_SL g1385 ( 
.A(n_1110),
.B(n_833),
.Y(n_1385)
);

OAI21x1_ASAP7_75t_L g1386 ( 
.A1(n_1138),
.A2(n_1151),
.B(n_1163),
.Y(n_1386)
);

OAI22xp5_ASAP7_75t_L g1387 ( 
.A1(n_1110),
.A2(n_909),
.B1(n_917),
.B2(n_1092),
.Y(n_1387)
);

OAI21x1_ASAP7_75t_L g1388 ( 
.A1(n_1138),
.A2(n_1151),
.B(n_1163),
.Y(n_1388)
);

NOR2xp67_ASAP7_75t_L g1389 ( 
.A(n_1203),
.B(n_929),
.Y(n_1389)
);

OAI21x1_ASAP7_75t_L g1390 ( 
.A1(n_1138),
.A2(n_1151),
.B(n_1163),
.Y(n_1390)
);

AOI22xp5_ASAP7_75t_L g1391 ( 
.A1(n_1110),
.A2(n_1070),
.B1(n_909),
.B2(n_967),
.Y(n_1391)
);

INVx1_ASAP7_75t_L g1392 ( 
.A(n_1301),
.Y(n_1392)
);

OAI21xp5_ASAP7_75t_L g1393 ( 
.A1(n_1391),
.A2(n_1378),
.B(n_1364),
.Y(n_1393)
);

BUFx2_ASAP7_75t_L g1394 ( 
.A(n_1370),
.Y(n_1394)
);

AND2x4_ASAP7_75t_L g1395 ( 
.A(n_1335),
.B(n_1344),
.Y(n_1395)
);

AOI21xp5_ASAP7_75t_L g1396 ( 
.A1(n_1367),
.A2(n_1379),
.B(n_1254),
.Y(n_1396)
);

OA21x2_ASAP7_75t_L g1397 ( 
.A1(n_1258),
.A2(n_1380),
.B(n_1375),
.Y(n_1397)
);

OAI21x1_ASAP7_75t_L g1398 ( 
.A1(n_1383),
.A2(n_1388),
.B(n_1386),
.Y(n_1398)
);

AND2x2_ASAP7_75t_L g1399 ( 
.A(n_1368),
.B(n_1373),
.Y(n_1399)
);

OAI22xp5_ASAP7_75t_L g1400 ( 
.A1(n_1391),
.A2(n_1385),
.B1(n_1387),
.B2(n_1382),
.Y(n_1400)
);

INVx1_ASAP7_75t_L g1401 ( 
.A(n_1252),
.Y(n_1401)
);

INVx1_ASAP7_75t_SL g1402 ( 
.A(n_1340),
.Y(n_1402)
);

OAI21x1_ASAP7_75t_L g1403 ( 
.A1(n_1390),
.A2(n_1369),
.B(n_1362),
.Y(n_1403)
);

BUFx12f_ASAP7_75t_L g1404 ( 
.A(n_1305),
.Y(n_1404)
);

INVx2_ASAP7_75t_L g1405 ( 
.A(n_1267),
.Y(n_1405)
);

OAI22xp5_ASAP7_75t_L g1406 ( 
.A1(n_1387),
.A2(n_1312),
.B1(n_1249),
.B2(n_1376),
.Y(n_1406)
);

AO31x2_ASAP7_75t_L g1407 ( 
.A1(n_1266),
.A2(n_1239),
.A3(n_1299),
.B(n_1262),
.Y(n_1407)
);

NAND2x1p5_ASAP7_75t_L g1408 ( 
.A(n_1344),
.B(n_1335),
.Y(n_1408)
);

NAND3xp33_ASAP7_75t_L g1409 ( 
.A(n_1317),
.B(n_1322),
.C(n_1330),
.Y(n_1409)
);

INVx2_ASAP7_75t_L g1410 ( 
.A(n_1267),
.Y(n_1410)
);

INVx1_ASAP7_75t_L g1411 ( 
.A(n_1265),
.Y(n_1411)
);

OAI21x1_ASAP7_75t_L g1412 ( 
.A1(n_1247),
.A2(n_1240),
.B(n_1278),
.Y(n_1412)
);

AND2x2_ASAP7_75t_L g1413 ( 
.A(n_1257),
.B(n_1276),
.Y(n_1413)
);

AOI22xp33_ASAP7_75t_L g1414 ( 
.A1(n_1311),
.A2(n_1242),
.B1(n_1273),
.B2(n_1239),
.Y(n_1414)
);

NAND2xp5_ASAP7_75t_L g1415 ( 
.A(n_1243),
.B(n_1280),
.Y(n_1415)
);

INVx2_ASAP7_75t_L g1416 ( 
.A(n_1245),
.Y(n_1416)
);

AOI21xp5_ASAP7_75t_L g1417 ( 
.A1(n_1253),
.A2(n_1366),
.B(n_1376),
.Y(n_1417)
);

INVx2_ASAP7_75t_L g1418 ( 
.A(n_1245),
.Y(n_1418)
);

NOR2xp67_ASAP7_75t_L g1419 ( 
.A(n_1306),
.B(n_1381),
.Y(n_1419)
);

INVx1_ASAP7_75t_L g1420 ( 
.A(n_1269),
.Y(n_1420)
);

OAI21x1_ASAP7_75t_L g1421 ( 
.A1(n_1279),
.A2(n_1303),
.B(n_1366),
.Y(n_1421)
);

HB1xp67_ASAP7_75t_L g1422 ( 
.A(n_1245),
.Y(n_1422)
);

INVx1_ASAP7_75t_L g1423 ( 
.A(n_1274),
.Y(n_1423)
);

INVx4_ASAP7_75t_SL g1424 ( 
.A(n_1242),
.Y(n_1424)
);

OAI21xp5_ASAP7_75t_L g1425 ( 
.A1(n_1270),
.A2(n_1313),
.B(n_1285),
.Y(n_1425)
);

AOI22x1_ASAP7_75t_L g1426 ( 
.A1(n_1319),
.A2(n_1372),
.B1(n_1287),
.B2(n_1363),
.Y(n_1426)
);

OAI22xp33_ASAP7_75t_L g1427 ( 
.A1(n_1242),
.A2(n_1273),
.B1(n_1338),
.B2(n_1283),
.Y(n_1427)
);

INVx1_ASAP7_75t_L g1428 ( 
.A(n_1284),
.Y(n_1428)
);

CKINVDCx16_ASAP7_75t_R g1429 ( 
.A(n_1282),
.Y(n_1429)
);

OAI21x1_ASAP7_75t_L g1430 ( 
.A1(n_1261),
.A2(n_1288),
.B(n_1304),
.Y(n_1430)
);

INVx2_ASAP7_75t_L g1431 ( 
.A(n_1315),
.Y(n_1431)
);

OA21x2_ASAP7_75t_L g1432 ( 
.A1(n_1261),
.A2(n_1244),
.B(n_1318),
.Y(n_1432)
);

OA21x2_ASAP7_75t_L g1433 ( 
.A1(n_1244),
.A2(n_1255),
.B(n_1302),
.Y(n_1433)
);

OAI21x1_ASAP7_75t_L g1434 ( 
.A1(n_1365),
.A2(n_1308),
.B(n_1324),
.Y(n_1434)
);

OAI21x1_ASAP7_75t_L g1435 ( 
.A1(n_1365),
.A2(n_1290),
.B(n_1298),
.Y(n_1435)
);

OAI21x1_ASAP7_75t_L g1436 ( 
.A1(n_1309),
.A2(n_1310),
.B(n_1286),
.Y(n_1436)
);

OAI22xp5_ASAP7_75t_L g1437 ( 
.A1(n_1270),
.A2(n_1241),
.B1(n_1336),
.B2(n_1343),
.Y(n_1437)
);

OAI21xp5_ASAP7_75t_L g1438 ( 
.A1(n_1313),
.A2(n_1263),
.B(n_1302),
.Y(n_1438)
);

AOI21xp5_ASAP7_75t_L g1439 ( 
.A1(n_1250),
.A2(n_1291),
.B(n_1248),
.Y(n_1439)
);

INVx2_ASAP7_75t_L g1440 ( 
.A(n_1260),
.Y(n_1440)
);

AOI22xp33_ASAP7_75t_L g1441 ( 
.A1(n_1273),
.A2(n_1271),
.B1(n_1277),
.B2(n_1251),
.Y(n_1441)
);

OAI21xp5_ASAP7_75t_L g1442 ( 
.A1(n_1255),
.A2(n_1351),
.B(n_1283),
.Y(n_1442)
);

AOI22xp33_ASAP7_75t_L g1443 ( 
.A1(n_1323),
.A2(n_1320),
.B1(n_1327),
.B2(n_1246),
.Y(n_1443)
);

OA21x2_ASAP7_75t_L g1444 ( 
.A1(n_1339),
.A2(n_1334),
.B(n_1289),
.Y(n_1444)
);

AOI221xp5_ASAP7_75t_L g1445 ( 
.A1(n_1316),
.A2(n_1377),
.B1(n_1371),
.B2(n_1332),
.C(n_1296),
.Y(n_1445)
);

AOI22xp33_ASAP7_75t_L g1446 ( 
.A1(n_1272),
.A2(n_1325),
.B1(n_1384),
.B2(n_1268),
.Y(n_1446)
);

OAI21x1_ASAP7_75t_L g1447 ( 
.A1(n_1326),
.A2(n_1342),
.B(n_1294),
.Y(n_1447)
);

OAI21x1_ASAP7_75t_L g1448 ( 
.A1(n_1359),
.A2(n_1353),
.B(n_1346),
.Y(n_1448)
);

OAI21x1_ASAP7_75t_L g1449 ( 
.A1(n_1353),
.A2(n_1297),
.B(n_1275),
.Y(n_1449)
);

BUFx3_ASAP7_75t_L g1450 ( 
.A(n_1256),
.Y(n_1450)
);

INVx1_ASAP7_75t_L g1451 ( 
.A(n_1268),
.Y(n_1451)
);

NOR2xp33_ASAP7_75t_L g1452 ( 
.A(n_1347),
.B(n_1307),
.Y(n_1452)
);

AOI21xp5_ASAP7_75t_L g1453 ( 
.A1(n_1248),
.A2(n_1295),
.B(n_1374),
.Y(n_1453)
);

OAI21x1_ASAP7_75t_SL g1454 ( 
.A1(n_1306),
.A2(n_1381),
.B(n_1360),
.Y(n_1454)
);

INVx2_ASAP7_75t_L g1455 ( 
.A(n_1292),
.Y(n_1455)
);

INVx4_ASAP7_75t_L g1456 ( 
.A(n_1300),
.Y(n_1456)
);

INVx2_ASAP7_75t_SL g1457 ( 
.A(n_1300),
.Y(n_1457)
);

OAI21x1_ASAP7_75t_L g1458 ( 
.A1(n_1281),
.A2(n_1357),
.B(n_1354),
.Y(n_1458)
);

OAI22xp5_ASAP7_75t_L g1459 ( 
.A1(n_1331),
.A2(n_1341),
.B1(n_1329),
.B2(n_1264),
.Y(n_1459)
);

OAI21x1_ASAP7_75t_L g1460 ( 
.A1(n_1389),
.A2(n_1356),
.B(n_1350),
.Y(n_1460)
);

AND2x4_ASAP7_75t_L g1461 ( 
.A(n_1361),
.B(n_1329),
.Y(n_1461)
);

AO21x2_ASAP7_75t_L g1462 ( 
.A1(n_1292),
.A2(n_1358),
.B(n_1374),
.Y(n_1462)
);

BUFx2_ASAP7_75t_L g1463 ( 
.A(n_1355),
.Y(n_1463)
);

AO32x2_ASAP7_75t_L g1464 ( 
.A1(n_1374),
.A2(n_1314),
.A3(n_1292),
.B1(n_1345),
.B2(n_1321),
.Y(n_1464)
);

OAI21x1_ASAP7_75t_L g1465 ( 
.A1(n_1321),
.A2(n_1337),
.B(n_1358),
.Y(n_1465)
);

AND2x2_ASAP7_75t_L g1466 ( 
.A(n_1259),
.B(n_1314),
.Y(n_1466)
);

AOI22xp5_ASAP7_75t_L g1467 ( 
.A1(n_1349),
.A2(n_1352),
.B1(n_1328),
.B2(n_1348),
.Y(n_1467)
);

OAI21x1_ASAP7_75t_L g1468 ( 
.A1(n_1321),
.A2(n_1337),
.B(n_1314),
.Y(n_1468)
);

AOI222xp33_ASAP7_75t_L g1469 ( 
.A1(n_1349),
.A2(n_1070),
.B1(n_845),
.B2(n_598),
.C1(n_616),
.C2(n_563),
.Y(n_1469)
);

OAI21x1_ASAP7_75t_SL g1470 ( 
.A1(n_1337),
.A2(n_1348),
.B(n_1391),
.Y(n_1470)
);

BUFx3_ASAP7_75t_L g1471 ( 
.A(n_1256),
.Y(n_1471)
);

AOI22xp33_ASAP7_75t_L g1472 ( 
.A1(n_1311),
.A2(n_1070),
.B1(n_1391),
.B2(n_1002),
.Y(n_1472)
);

INVx1_ASAP7_75t_L g1473 ( 
.A(n_1301),
.Y(n_1473)
);

INVx2_ASAP7_75t_L g1474 ( 
.A(n_1267),
.Y(n_1474)
);

INVx1_ASAP7_75t_L g1475 ( 
.A(n_1301),
.Y(n_1475)
);

BUFx3_ASAP7_75t_L g1476 ( 
.A(n_1256),
.Y(n_1476)
);

AND2x4_ASAP7_75t_L g1477 ( 
.A(n_1335),
.B(n_1344),
.Y(n_1477)
);

AND3x2_ASAP7_75t_L g1478 ( 
.A(n_1330),
.B(n_1002),
.C(n_722),
.Y(n_1478)
);

INVx3_ASAP7_75t_L g1479 ( 
.A(n_1293),
.Y(n_1479)
);

OAI21x1_ASAP7_75t_L g1480 ( 
.A1(n_1375),
.A2(n_1383),
.B(n_1380),
.Y(n_1480)
);

OAI21xp5_ASAP7_75t_L g1481 ( 
.A1(n_1391),
.A2(n_833),
.B(n_1110),
.Y(n_1481)
);

BUFx3_ASAP7_75t_L g1482 ( 
.A(n_1256),
.Y(n_1482)
);

INVx4_ASAP7_75t_L g1483 ( 
.A(n_1300),
.Y(n_1483)
);

INVx1_ASAP7_75t_L g1484 ( 
.A(n_1301),
.Y(n_1484)
);

AND2x4_ASAP7_75t_L g1485 ( 
.A(n_1335),
.B(n_1344),
.Y(n_1485)
);

O2A1O1Ixp33_ASAP7_75t_L g1486 ( 
.A1(n_1385),
.A2(n_833),
.B(n_1110),
.C(n_909),
.Y(n_1486)
);

OAI21xp5_ASAP7_75t_L g1487 ( 
.A1(n_1391),
.A2(n_833),
.B(n_1110),
.Y(n_1487)
);

OAI21x1_ASAP7_75t_L g1488 ( 
.A1(n_1375),
.A2(n_1383),
.B(n_1380),
.Y(n_1488)
);

OAI21xp5_ASAP7_75t_L g1489 ( 
.A1(n_1391),
.A2(n_833),
.B(n_1110),
.Y(n_1489)
);

AOI21xp5_ASAP7_75t_L g1490 ( 
.A1(n_1367),
.A2(n_1097),
.B(n_986),
.Y(n_1490)
);

AOI22xp33_ASAP7_75t_L g1491 ( 
.A1(n_1311),
.A2(n_1070),
.B1(n_1391),
.B2(n_1002),
.Y(n_1491)
);

INVx2_ASAP7_75t_L g1492 ( 
.A(n_1267),
.Y(n_1492)
);

AND2x2_ASAP7_75t_L g1493 ( 
.A(n_1368),
.B(n_1116),
.Y(n_1493)
);

INVx2_ASAP7_75t_L g1494 ( 
.A(n_1267),
.Y(n_1494)
);

NAND2x1p5_ASAP7_75t_L g1495 ( 
.A(n_1344),
.B(n_1206),
.Y(n_1495)
);

AND2x4_ASAP7_75t_L g1496 ( 
.A(n_1335),
.B(n_1344),
.Y(n_1496)
);

AND2x4_ASAP7_75t_L g1497 ( 
.A(n_1335),
.B(n_1344),
.Y(n_1497)
);

AOI21xp5_ASAP7_75t_L g1498 ( 
.A1(n_1367),
.A2(n_1097),
.B(n_986),
.Y(n_1498)
);

INVx3_ASAP7_75t_L g1499 ( 
.A(n_1293),
.Y(n_1499)
);

BUFx6f_ASAP7_75t_L g1500 ( 
.A(n_1335),
.Y(n_1500)
);

INVx1_ASAP7_75t_L g1501 ( 
.A(n_1301),
.Y(n_1501)
);

AO31x2_ASAP7_75t_L g1502 ( 
.A1(n_1266),
.A2(n_1239),
.A3(n_1299),
.B(n_1262),
.Y(n_1502)
);

OAI21x1_ASAP7_75t_L g1503 ( 
.A1(n_1375),
.A2(n_1383),
.B(n_1380),
.Y(n_1503)
);

BUFx3_ASAP7_75t_L g1504 ( 
.A(n_1256),
.Y(n_1504)
);

OAI21x1_ASAP7_75t_L g1505 ( 
.A1(n_1375),
.A2(n_1383),
.B(n_1380),
.Y(n_1505)
);

OAI21x1_ASAP7_75t_L g1506 ( 
.A1(n_1375),
.A2(n_1383),
.B(n_1380),
.Y(n_1506)
);

AND2x2_ASAP7_75t_L g1507 ( 
.A(n_1368),
.B(n_1116),
.Y(n_1507)
);

OAI21xp5_ASAP7_75t_L g1508 ( 
.A1(n_1391),
.A2(n_833),
.B(n_1110),
.Y(n_1508)
);

INVx4_ASAP7_75t_L g1509 ( 
.A(n_1300),
.Y(n_1509)
);

AND2x2_ASAP7_75t_L g1510 ( 
.A(n_1368),
.B(n_1116),
.Y(n_1510)
);

OA21x2_ASAP7_75t_L g1511 ( 
.A1(n_1258),
.A2(n_1380),
.B(n_1375),
.Y(n_1511)
);

OR2x2_ASAP7_75t_L g1512 ( 
.A(n_1368),
.B(n_1373),
.Y(n_1512)
);

INVx1_ASAP7_75t_L g1513 ( 
.A(n_1301),
.Y(n_1513)
);

INVx2_ASAP7_75t_L g1514 ( 
.A(n_1267),
.Y(n_1514)
);

INVx1_ASAP7_75t_L g1515 ( 
.A(n_1301),
.Y(n_1515)
);

OA21x2_ASAP7_75t_L g1516 ( 
.A1(n_1258),
.A2(n_1380),
.B(n_1375),
.Y(n_1516)
);

AO32x2_ASAP7_75t_L g1517 ( 
.A1(n_1239),
.A2(n_1387),
.A3(n_1336),
.B1(n_1378),
.B2(n_1364),
.Y(n_1517)
);

AO31x2_ASAP7_75t_L g1518 ( 
.A1(n_1266),
.A2(n_1239),
.A3(n_1299),
.B(n_1262),
.Y(n_1518)
);

CKINVDCx20_ASAP7_75t_R g1519 ( 
.A(n_1282),
.Y(n_1519)
);

OAI21x1_ASAP7_75t_L g1520 ( 
.A1(n_1375),
.A2(n_1383),
.B(n_1380),
.Y(n_1520)
);

AND2x4_ASAP7_75t_L g1521 ( 
.A(n_1335),
.B(n_1344),
.Y(n_1521)
);

INVx2_ASAP7_75t_L g1522 ( 
.A(n_1267),
.Y(n_1522)
);

NAND2xp5_ASAP7_75t_L g1523 ( 
.A(n_1368),
.B(n_1373),
.Y(n_1523)
);

OA21x2_ASAP7_75t_L g1524 ( 
.A1(n_1258),
.A2(n_1380),
.B(n_1375),
.Y(n_1524)
);

CKINVDCx14_ASAP7_75t_R g1525 ( 
.A(n_1282),
.Y(n_1525)
);

OAI22xp5_ASAP7_75t_L g1526 ( 
.A1(n_1391),
.A2(n_909),
.B1(n_833),
.B2(n_1110),
.Y(n_1526)
);

OR2x2_ASAP7_75t_L g1527 ( 
.A(n_1368),
.B(n_1373),
.Y(n_1527)
);

INVx4_ASAP7_75t_L g1528 ( 
.A(n_1300),
.Y(n_1528)
);

OAI21x1_ASAP7_75t_L g1529 ( 
.A1(n_1375),
.A2(n_1383),
.B(n_1380),
.Y(n_1529)
);

INVx2_ASAP7_75t_L g1530 ( 
.A(n_1267),
.Y(n_1530)
);

INVx1_ASAP7_75t_L g1531 ( 
.A(n_1301),
.Y(n_1531)
);

OAI21x1_ASAP7_75t_L g1532 ( 
.A1(n_1375),
.A2(n_1383),
.B(n_1380),
.Y(n_1532)
);

NAND2xp5_ASAP7_75t_L g1533 ( 
.A(n_1368),
.B(n_1373),
.Y(n_1533)
);

OA21x2_ASAP7_75t_L g1534 ( 
.A1(n_1258),
.A2(n_1380),
.B(n_1375),
.Y(n_1534)
);

OAI21xp5_ASAP7_75t_L g1535 ( 
.A1(n_1391),
.A2(n_833),
.B(n_1110),
.Y(n_1535)
);

OAI21xp5_ASAP7_75t_L g1536 ( 
.A1(n_1391),
.A2(n_833),
.B(n_1110),
.Y(n_1536)
);

OA21x2_ASAP7_75t_L g1537 ( 
.A1(n_1258),
.A2(n_1380),
.B(n_1375),
.Y(n_1537)
);

OAI21x1_ASAP7_75t_L g1538 ( 
.A1(n_1375),
.A2(n_1383),
.B(n_1380),
.Y(n_1538)
);

HB1xp67_ASAP7_75t_L g1539 ( 
.A(n_1245),
.Y(n_1539)
);

CKINVDCx20_ASAP7_75t_R g1540 ( 
.A(n_1282),
.Y(n_1540)
);

INVx1_ASAP7_75t_L g1541 ( 
.A(n_1301),
.Y(n_1541)
);

CKINVDCx5p33_ASAP7_75t_R g1542 ( 
.A(n_1404),
.Y(n_1542)
);

NAND2xp5_ASAP7_75t_L g1543 ( 
.A(n_1392),
.B(n_1473),
.Y(n_1543)
);

OA21x2_ASAP7_75t_L g1544 ( 
.A1(n_1439),
.A2(n_1403),
.B(n_1465),
.Y(n_1544)
);

OAI22xp5_ASAP7_75t_L g1545 ( 
.A1(n_1393),
.A2(n_1526),
.B1(n_1472),
.B2(n_1491),
.Y(n_1545)
);

HB1xp67_ASAP7_75t_L g1546 ( 
.A(n_1463),
.Y(n_1546)
);

NAND2xp5_ASAP7_75t_L g1547 ( 
.A(n_1475),
.B(n_1484),
.Y(n_1547)
);

AND2x2_ASAP7_75t_L g1548 ( 
.A(n_1413),
.B(n_1399),
.Y(n_1548)
);

OAI22xp5_ASAP7_75t_L g1549 ( 
.A1(n_1472),
.A2(n_1491),
.B1(n_1508),
.B2(n_1481),
.Y(n_1549)
);

OA22x2_ASAP7_75t_L g1550 ( 
.A1(n_1442),
.A2(n_1478),
.B1(n_1406),
.B2(n_1466),
.Y(n_1550)
);

NOR2xp33_ASAP7_75t_L g1551 ( 
.A(n_1402),
.B(n_1519),
.Y(n_1551)
);

O2A1O1Ixp33_ASAP7_75t_L g1552 ( 
.A1(n_1487),
.A2(n_1489),
.B(n_1535),
.C(n_1536),
.Y(n_1552)
);

BUFx12f_ASAP7_75t_L g1553 ( 
.A(n_1404),
.Y(n_1553)
);

INVx1_ASAP7_75t_L g1554 ( 
.A(n_1401),
.Y(n_1554)
);

A2O1A1Ixp33_ASAP7_75t_L g1555 ( 
.A1(n_1409),
.A2(n_1425),
.B(n_1486),
.C(n_1400),
.Y(n_1555)
);

OAI22xp5_ASAP7_75t_L g1556 ( 
.A1(n_1414),
.A2(n_1443),
.B1(n_1437),
.B2(n_1441),
.Y(n_1556)
);

AND2x2_ASAP7_75t_L g1557 ( 
.A(n_1493),
.B(n_1507),
.Y(n_1557)
);

OR2x2_ASAP7_75t_L g1558 ( 
.A(n_1512),
.B(n_1527),
.Y(n_1558)
);

A2O1A1Ixp33_ASAP7_75t_L g1559 ( 
.A1(n_1438),
.A2(n_1443),
.B(n_1417),
.C(n_1453),
.Y(n_1559)
);

OAI22xp5_ASAP7_75t_L g1560 ( 
.A1(n_1414),
.A2(n_1441),
.B1(n_1427),
.B2(n_1433),
.Y(n_1560)
);

AOI21xp5_ASAP7_75t_SL g1561 ( 
.A1(n_1415),
.A2(n_1459),
.B(n_1427),
.Y(n_1561)
);

AOI21xp5_ASAP7_75t_L g1562 ( 
.A1(n_1396),
.A2(n_1498),
.B(n_1490),
.Y(n_1562)
);

AND2x2_ASAP7_75t_L g1563 ( 
.A(n_1510),
.B(n_1394),
.Y(n_1563)
);

CKINVDCx20_ASAP7_75t_R g1564 ( 
.A(n_1519),
.Y(n_1564)
);

CKINVDCx5p33_ASAP7_75t_R g1565 ( 
.A(n_1540),
.Y(n_1565)
);

NAND2xp5_ASAP7_75t_L g1566 ( 
.A(n_1501),
.B(n_1513),
.Y(n_1566)
);

A2O1A1Ixp33_ASAP7_75t_SL g1567 ( 
.A1(n_1525),
.A2(n_1479),
.B(n_1499),
.C(n_1452),
.Y(n_1567)
);

NOR2xp67_ASAP7_75t_L g1568 ( 
.A(n_1467),
.B(n_1456),
.Y(n_1568)
);

OR2x2_ASAP7_75t_L g1569 ( 
.A(n_1523),
.B(n_1533),
.Y(n_1569)
);

INVx1_ASAP7_75t_L g1570 ( 
.A(n_1411),
.Y(n_1570)
);

NAND2xp5_ASAP7_75t_L g1571 ( 
.A(n_1515),
.B(n_1531),
.Y(n_1571)
);

AND2x2_ASAP7_75t_L g1572 ( 
.A(n_1452),
.B(n_1541),
.Y(n_1572)
);

OR2x2_ASAP7_75t_SL g1573 ( 
.A(n_1429),
.B(n_1420),
.Y(n_1573)
);

OR2x2_ASAP7_75t_L g1574 ( 
.A(n_1423),
.B(n_1428),
.Y(n_1574)
);

OA21x2_ASAP7_75t_L g1575 ( 
.A1(n_1403),
.A2(n_1465),
.B(n_1421),
.Y(n_1575)
);

HB1xp67_ASAP7_75t_L g1576 ( 
.A(n_1422),
.Y(n_1576)
);

AOI21xp5_ASAP7_75t_SL g1577 ( 
.A1(n_1445),
.A2(n_1482),
.B(n_1450),
.Y(n_1577)
);

HB1xp67_ASAP7_75t_L g1578 ( 
.A(n_1539),
.Y(n_1578)
);

NOR2xp33_ASAP7_75t_L g1579 ( 
.A(n_1540),
.B(n_1457),
.Y(n_1579)
);

OR2x2_ASAP7_75t_L g1580 ( 
.A(n_1433),
.B(n_1440),
.Y(n_1580)
);

OA21x2_ASAP7_75t_L g1581 ( 
.A1(n_1468),
.A2(n_1434),
.B(n_1538),
.Y(n_1581)
);

HB1xp67_ASAP7_75t_L g1582 ( 
.A(n_1539),
.Y(n_1582)
);

AND2x2_ASAP7_75t_SL g1583 ( 
.A(n_1395),
.B(n_1477),
.Y(n_1583)
);

OAI22xp5_ASAP7_75t_L g1584 ( 
.A1(n_1433),
.A2(n_1432),
.B1(n_1517),
.B2(n_1426),
.Y(n_1584)
);

OAI22xp5_ASAP7_75t_L g1585 ( 
.A1(n_1432),
.A2(n_1517),
.B1(n_1446),
.B2(n_1525),
.Y(n_1585)
);

OA21x2_ASAP7_75t_L g1586 ( 
.A1(n_1468),
.A2(n_1434),
.B(n_1538),
.Y(n_1586)
);

OAI22xp5_ASAP7_75t_L g1587 ( 
.A1(n_1432),
.A2(n_1517),
.B1(n_1446),
.B2(n_1528),
.Y(n_1587)
);

AOI21xp5_ASAP7_75t_L g1588 ( 
.A1(n_1397),
.A2(n_1524),
.B(n_1516),
.Y(n_1588)
);

AOI21xp5_ASAP7_75t_L g1589 ( 
.A1(n_1397),
.A2(n_1524),
.B(n_1516),
.Y(n_1589)
);

NAND2xp5_ASAP7_75t_L g1590 ( 
.A(n_1416),
.B(n_1418),
.Y(n_1590)
);

AOI221x1_ASAP7_75t_SL g1591 ( 
.A1(n_1517),
.A2(n_1469),
.B1(n_1419),
.B2(n_1405),
.C(n_1530),
.Y(n_1591)
);

AND2x2_ASAP7_75t_SL g1592 ( 
.A(n_1477),
.B(n_1485),
.Y(n_1592)
);

AND2x4_ASAP7_75t_L g1593 ( 
.A(n_1424),
.B(n_1497),
.Y(n_1593)
);

OA21x2_ASAP7_75t_L g1594 ( 
.A1(n_1398),
.A2(n_1480),
.B(n_1488),
.Y(n_1594)
);

AND2x4_ASAP7_75t_L g1595 ( 
.A(n_1485),
.B(n_1497),
.Y(n_1595)
);

OAI22xp5_ASAP7_75t_L g1596 ( 
.A1(n_1483),
.A2(n_1509),
.B1(n_1528),
.B2(n_1408),
.Y(n_1596)
);

AND2x4_ASAP7_75t_L g1597 ( 
.A(n_1496),
.B(n_1521),
.Y(n_1597)
);

INVx1_ASAP7_75t_L g1598 ( 
.A(n_1470),
.Y(n_1598)
);

AND2x2_ASAP7_75t_L g1599 ( 
.A(n_1496),
.B(n_1521),
.Y(n_1599)
);

OAI22xp5_ASAP7_75t_L g1600 ( 
.A1(n_1483),
.A2(n_1509),
.B1(n_1408),
.B2(n_1504),
.Y(n_1600)
);

OAI22xp5_ASAP7_75t_L g1601 ( 
.A1(n_1471),
.A2(n_1476),
.B1(n_1504),
.B2(n_1500),
.Y(n_1601)
);

O2A1O1Ixp33_ASAP7_75t_L g1602 ( 
.A1(n_1454),
.A2(n_1522),
.B(n_1474),
.C(n_1410),
.Y(n_1602)
);

AND2x2_ASAP7_75t_L g1603 ( 
.A(n_1500),
.B(n_1460),
.Y(n_1603)
);

AND2x2_ASAP7_75t_L g1604 ( 
.A(n_1458),
.B(n_1464),
.Y(n_1604)
);

A2O1A1Ixp33_ASAP7_75t_L g1605 ( 
.A1(n_1430),
.A2(n_1435),
.B(n_1514),
.C(n_1492),
.Y(n_1605)
);

AND2x2_ASAP7_75t_L g1606 ( 
.A(n_1464),
.B(n_1430),
.Y(n_1606)
);

OAI22xp5_ASAP7_75t_L g1607 ( 
.A1(n_1494),
.A2(n_1530),
.B1(n_1522),
.B2(n_1495),
.Y(n_1607)
);

INVx1_ASAP7_75t_SL g1608 ( 
.A(n_1444),
.Y(n_1608)
);

INVxp33_ASAP7_75t_L g1609 ( 
.A(n_1448),
.Y(n_1609)
);

AOI21xp5_ASAP7_75t_SL g1610 ( 
.A1(n_1444),
.A2(n_1494),
.B(n_1462),
.Y(n_1610)
);

OAI22xp5_ASAP7_75t_L g1611 ( 
.A1(n_1478),
.A2(n_1537),
.B1(n_1511),
.B2(n_1534),
.Y(n_1611)
);

CKINVDCx5p33_ASAP7_75t_R g1612 ( 
.A(n_1431),
.Y(n_1612)
);

INVxp67_ASAP7_75t_L g1613 ( 
.A(n_1448),
.Y(n_1613)
);

A2O1A1Ixp33_ASAP7_75t_L g1614 ( 
.A1(n_1435),
.A2(n_1436),
.B(n_1447),
.C(n_1449),
.Y(n_1614)
);

OA21x2_ASAP7_75t_L g1615 ( 
.A1(n_1503),
.A2(n_1506),
.B(n_1505),
.Y(n_1615)
);

OR2x2_ASAP7_75t_L g1616 ( 
.A(n_1407),
.B(n_1502),
.Y(n_1616)
);

INVx4_ASAP7_75t_SL g1617 ( 
.A(n_1407),
.Y(n_1617)
);

AOI21xp5_ASAP7_75t_SL g1618 ( 
.A1(n_1534),
.A2(n_1455),
.B(n_1464),
.Y(n_1618)
);

NAND2xp5_ASAP7_75t_L g1619 ( 
.A(n_1502),
.B(n_1518),
.Y(n_1619)
);

O2A1O1Ixp5_ASAP7_75t_L g1620 ( 
.A1(n_1502),
.A2(n_1518),
.B(n_1449),
.C(n_1412),
.Y(n_1620)
);

NOR2xp67_ASAP7_75t_R g1621 ( 
.A(n_1502),
.B(n_1518),
.Y(n_1621)
);

INVx1_ASAP7_75t_L g1622 ( 
.A(n_1412),
.Y(n_1622)
);

INVx2_ASAP7_75t_L g1623 ( 
.A(n_1436),
.Y(n_1623)
);

CKINVDCx5p33_ASAP7_75t_R g1624 ( 
.A(n_1532),
.Y(n_1624)
);

AOI21xp5_ASAP7_75t_SL g1625 ( 
.A1(n_1520),
.A2(n_1110),
.B(n_1406),
.Y(n_1625)
);

NAND2xp5_ASAP7_75t_L g1626 ( 
.A(n_1529),
.B(n_1392),
.Y(n_1626)
);

CKINVDCx5p33_ASAP7_75t_R g1627 ( 
.A(n_1404),
.Y(n_1627)
);

O2A1O1Ixp33_ASAP7_75t_L g1628 ( 
.A1(n_1526),
.A2(n_1481),
.B(n_1489),
.C(n_1487),
.Y(n_1628)
);

AOI21x1_ASAP7_75t_SL g1629 ( 
.A1(n_1466),
.A2(n_1333),
.B(n_1208),
.Y(n_1629)
);

AND2x4_ASAP7_75t_L g1630 ( 
.A(n_1424),
.B(n_1461),
.Y(n_1630)
);

AND2x2_ASAP7_75t_L g1631 ( 
.A(n_1413),
.B(n_1399),
.Y(n_1631)
);

AND2x2_ASAP7_75t_L g1632 ( 
.A(n_1413),
.B(n_1399),
.Y(n_1632)
);

HB1xp67_ASAP7_75t_L g1633 ( 
.A(n_1463),
.Y(n_1633)
);

O2A1O1Ixp33_ASAP7_75t_L g1634 ( 
.A1(n_1526),
.A2(n_1481),
.B(n_1489),
.C(n_1487),
.Y(n_1634)
);

AND2x2_ASAP7_75t_L g1635 ( 
.A(n_1413),
.B(n_1399),
.Y(n_1635)
);

INVx4_ASAP7_75t_SL g1636 ( 
.A(n_1451),
.Y(n_1636)
);

AND2x2_ASAP7_75t_L g1637 ( 
.A(n_1413),
.B(n_1399),
.Y(n_1637)
);

INVx1_ASAP7_75t_L g1638 ( 
.A(n_1401),
.Y(n_1638)
);

NAND2xp5_ASAP7_75t_L g1639 ( 
.A(n_1392),
.B(n_1473),
.Y(n_1639)
);

BUFx3_ASAP7_75t_L g1640 ( 
.A(n_1394),
.Y(n_1640)
);

AND2x4_ASAP7_75t_L g1641 ( 
.A(n_1424),
.B(n_1461),
.Y(n_1641)
);

AND2x2_ASAP7_75t_L g1642 ( 
.A(n_1413),
.B(n_1399),
.Y(n_1642)
);

A2O1A1Ixp33_ASAP7_75t_L g1643 ( 
.A1(n_1409),
.A2(n_1393),
.B(n_1442),
.C(n_1125),
.Y(n_1643)
);

AND2x2_ASAP7_75t_L g1644 ( 
.A(n_1606),
.B(n_1604),
.Y(n_1644)
);

INVx1_ASAP7_75t_L g1645 ( 
.A(n_1626),
.Y(n_1645)
);

INVx1_ASAP7_75t_L g1646 ( 
.A(n_1626),
.Y(n_1646)
);

OR2x6_ASAP7_75t_L g1647 ( 
.A(n_1618),
.B(n_1610),
.Y(n_1647)
);

INVx1_ASAP7_75t_L g1648 ( 
.A(n_1554),
.Y(n_1648)
);

INVx1_ASAP7_75t_L g1649 ( 
.A(n_1570),
.Y(n_1649)
);

NAND2xp5_ASAP7_75t_L g1650 ( 
.A(n_1559),
.B(n_1585),
.Y(n_1650)
);

HB1xp67_ASAP7_75t_L g1651 ( 
.A(n_1546),
.Y(n_1651)
);

AND2x2_ASAP7_75t_L g1652 ( 
.A(n_1638),
.B(n_1548),
.Y(n_1652)
);

OR2x6_ASAP7_75t_L g1653 ( 
.A(n_1577),
.B(n_1560),
.Y(n_1653)
);

INVx1_ASAP7_75t_L g1654 ( 
.A(n_1580),
.Y(n_1654)
);

AND2x2_ASAP7_75t_L g1655 ( 
.A(n_1631),
.B(n_1632),
.Y(n_1655)
);

AND2x2_ASAP7_75t_L g1656 ( 
.A(n_1635),
.B(n_1637),
.Y(n_1656)
);

HB1xp67_ASAP7_75t_L g1657 ( 
.A(n_1633),
.Y(n_1657)
);

AND2x2_ASAP7_75t_L g1658 ( 
.A(n_1642),
.B(n_1563),
.Y(n_1658)
);

INVx1_ASAP7_75t_L g1659 ( 
.A(n_1574),
.Y(n_1659)
);

INVx3_ASAP7_75t_L g1660 ( 
.A(n_1581),
.Y(n_1660)
);

AO21x1_ASAP7_75t_SL g1661 ( 
.A1(n_1619),
.A2(n_1616),
.B(n_1598),
.Y(n_1661)
);

NAND2x1p5_ASAP7_75t_L g1662 ( 
.A(n_1583),
.B(n_1592),
.Y(n_1662)
);

AND2x2_ASAP7_75t_L g1663 ( 
.A(n_1617),
.B(n_1557),
.Y(n_1663)
);

AOI21x1_ASAP7_75t_L g1664 ( 
.A1(n_1611),
.A2(n_1588),
.B(n_1589),
.Y(n_1664)
);

HB1xp67_ASAP7_75t_L g1665 ( 
.A(n_1576),
.Y(n_1665)
);

OR2x2_ASAP7_75t_L g1666 ( 
.A(n_1578),
.B(n_1582),
.Y(n_1666)
);

NAND2xp5_ASAP7_75t_L g1667 ( 
.A(n_1585),
.B(n_1572),
.Y(n_1667)
);

HB1xp67_ASAP7_75t_L g1668 ( 
.A(n_1640),
.Y(n_1668)
);

INVx1_ASAP7_75t_L g1669 ( 
.A(n_1543),
.Y(n_1669)
);

INVx1_ASAP7_75t_L g1670 ( 
.A(n_1543),
.Y(n_1670)
);

INVx1_ASAP7_75t_L g1671 ( 
.A(n_1547),
.Y(n_1671)
);

INVx1_ASAP7_75t_L g1672 ( 
.A(n_1547),
.Y(n_1672)
);

AO21x2_ASAP7_75t_L g1673 ( 
.A1(n_1605),
.A2(n_1584),
.B(n_1587),
.Y(n_1673)
);

INVx1_ASAP7_75t_L g1674 ( 
.A(n_1566),
.Y(n_1674)
);

INVx1_ASAP7_75t_L g1675 ( 
.A(n_1566),
.Y(n_1675)
);

BUFx2_ASAP7_75t_L g1676 ( 
.A(n_1624),
.Y(n_1676)
);

AND2x2_ASAP7_75t_L g1677 ( 
.A(n_1609),
.B(n_1613),
.Y(n_1677)
);

NOR2x1p5_ASAP7_75t_L g1678 ( 
.A(n_1553),
.B(n_1593),
.Y(n_1678)
);

HB1xp67_ASAP7_75t_L g1679 ( 
.A(n_1571),
.Y(n_1679)
);

INVx1_ASAP7_75t_L g1680 ( 
.A(n_1639),
.Y(n_1680)
);

OAI22xp5_ASAP7_75t_L g1681 ( 
.A1(n_1545),
.A2(n_1555),
.B1(n_1549),
.B2(n_1643),
.Y(n_1681)
);

OA21x2_ASAP7_75t_L g1682 ( 
.A1(n_1620),
.A2(n_1562),
.B(n_1614),
.Y(n_1682)
);

OR2x6_ASAP7_75t_L g1683 ( 
.A(n_1560),
.B(n_1593),
.Y(n_1683)
);

INVx3_ASAP7_75t_L g1684 ( 
.A(n_1586),
.Y(n_1684)
);

AO21x2_ASAP7_75t_L g1685 ( 
.A1(n_1562),
.A2(n_1549),
.B(n_1545),
.Y(n_1685)
);

AO21x2_ASAP7_75t_L g1686 ( 
.A1(n_1590),
.A2(n_1623),
.B(n_1556),
.Y(n_1686)
);

AND2x2_ASAP7_75t_L g1687 ( 
.A(n_1608),
.B(n_1612),
.Y(n_1687)
);

OAI22xp33_ASAP7_75t_L g1688 ( 
.A1(n_1550),
.A2(n_1600),
.B1(n_1568),
.B2(n_1552),
.Y(n_1688)
);

AND2x2_ASAP7_75t_L g1689 ( 
.A(n_1608),
.B(n_1603),
.Y(n_1689)
);

BUFx3_ASAP7_75t_L g1690 ( 
.A(n_1595),
.Y(n_1690)
);

INVx2_ASAP7_75t_SL g1691 ( 
.A(n_1599),
.Y(n_1691)
);

AND2x4_ASAP7_75t_L g1692 ( 
.A(n_1636),
.B(n_1597),
.Y(n_1692)
);

INVx1_ASAP7_75t_L g1693 ( 
.A(n_1602),
.Y(n_1693)
);

NOR2xp33_ASAP7_75t_L g1694 ( 
.A(n_1565),
.B(n_1564),
.Y(n_1694)
);

NAND2x1_ASAP7_75t_L g1695 ( 
.A(n_1625),
.B(n_1561),
.Y(n_1695)
);

AO21x2_ASAP7_75t_L g1696 ( 
.A1(n_1607),
.A2(n_1622),
.B(n_1628),
.Y(n_1696)
);

BUFx2_ASAP7_75t_L g1697 ( 
.A(n_1575),
.Y(n_1697)
);

INVx1_ASAP7_75t_L g1698 ( 
.A(n_1607),
.Y(n_1698)
);

AOI21xp5_ASAP7_75t_SL g1699 ( 
.A1(n_1634),
.A2(n_1600),
.B(n_1596),
.Y(n_1699)
);

AND2x2_ASAP7_75t_L g1700 ( 
.A(n_1575),
.B(n_1544),
.Y(n_1700)
);

OR2x2_ASAP7_75t_L g1701 ( 
.A(n_1667),
.B(n_1573),
.Y(n_1701)
);

INVx1_ASAP7_75t_L g1702 ( 
.A(n_1648),
.Y(n_1702)
);

INVx4_ASAP7_75t_L g1703 ( 
.A(n_1685),
.Y(n_1703)
);

OR2x6_ASAP7_75t_L g1704 ( 
.A(n_1647),
.B(n_1662),
.Y(n_1704)
);

AND2x4_ASAP7_75t_L g1705 ( 
.A(n_1692),
.B(n_1595),
.Y(n_1705)
);

OR2x2_ASAP7_75t_L g1706 ( 
.A(n_1667),
.B(n_1558),
.Y(n_1706)
);

AOI22xp5_ASAP7_75t_L g1707 ( 
.A1(n_1681),
.A2(n_1596),
.B1(n_1601),
.B2(n_1569),
.Y(n_1707)
);

HB1xp67_ASAP7_75t_L g1708 ( 
.A(n_1665),
.Y(n_1708)
);

AND2x2_ASAP7_75t_L g1709 ( 
.A(n_1644),
.B(n_1594),
.Y(n_1709)
);

AND2x2_ASAP7_75t_L g1710 ( 
.A(n_1644),
.B(n_1594),
.Y(n_1710)
);

INVx1_ASAP7_75t_L g1711 ( 
.A(n_1648),
.Y(n_1711)
);

HB1xp67_ASAP7_75t_L g1712 ( 
.A(n_1645),
.Y(n_1712)
);

INVxp67_ASAP7_75t_SL g1713 ( 
.A(n_1660),
.Y(n_1713)
);

NAND2xp5_ASAP7_75t_L g1714 ( 
.A(n_1685),
.B(n_1679),
.Y(n_1714)
);

INVx1_ASAP7_75t_L g1715 ( 
.A(n_1649),
.Y(n_1715)
);

AND2x2_ASAP7_75t_L g1716 ( 
.A(n_1673),
.B(n_1646),
.Y(n_1716)
);

INVxp67_ASAP7_75t_SL g1717 ( 
.A(n_1660),
.Y(n_1717)
);

BUFx3_ASAP7_75t_L g1718 ( 
.A(n_1695),
.Y(n_1718)
);

AND2x2_ASAP7_75t_L g1719 ( 
.A(n_1673),
.B(n_1615),
.Y(n_1719)
);

INVx1_ASAP7_75t_L g1720 ( 
.A(n_1654),
.Y(n_1720)
);

HB1xp67_ASAP7_75t_L g1721 ( 
.A(n_1666),
.Y(n_1721)
);

AND2x2_ASAP7_75t_L g1722 ( 
.A(n_1673),
.B(n_1697),
.Y(n_1722)
);

BUFx2_ASAP7_75t_L g1723 ( 
.A(n_1666),
.Y(n_1723)
);

INVxp67_ASAP7_75t_L g1724 ( 
.A(n_1661),
.Y(n_1724)
);

NAND2xp5_ASAP7_75t_L g1725 ( 
.A(n_1685),
.B(n_1621),
.Y(n_1725)
);

AND2x2_ASAP7_75t_L g1726 ( 
.A(n_1673),
.B(n_1697),
.Y(n_1726)
);

NAND2xp5_ASAP7_75t_L g1727 ( 
.A(n_1685),
.B(n_1591),
.Y(n_1727)
);

INVx2_ASAP7_75t_SL g1728 ( 
.A(n_1689),
.Y(n_1728)
);

HB1xp67_ASAP7_75t_L g1729 ( 
.A(n_1651),
.Y(n_1729)
);

INVx5_ASAP7_75t_L g1730 ( 
.A(n_1647),
.Y(n_1730)
);

NOR2xp33_ASAP7_75t_L g1731 ( 
.A(n_1668),
.B(n_1542),
.Y(n_1731)
);

AOI22xp33_ASAP7_75t_SL g1732 ( 
.A1(n_1681),
.A2(n_1630),
.B1(n_1641),
.B2(n_1629),
.Y(n_1732)
);

CKINVDCx5p33_ASAP7_75t_R g1733 ( 
.A(n_1731),
.Y(n_1733)
);

INVx1_ASAP7_75t_L g1734 ( 
.A(n_1702),
.Y(n_1734)
);

NAND2xp5_ASAP7_75t_L g1735 ( 
.A(n_1708),
.B(n_1655),
.Y(n_1735)
);

AND2x4_ASAP7_75t_L g1736 ( 
.A(n_1724),
.B(n_1690),
.Y(n_1736)
);

NAND2xp5_ASAP7_75t_L g1737 ( 
.A(n_1708),
.B(n_1655),
.Y(n_1737)
);

INVx1_ASAP7_75t_L g1738 ( 
.A(n_1711),
.Y(n_1738)
);

OAI221xp5_ASAP7_75t_L g1739 ( 
.A1(n_1727),
.A2(n_1650),
.B1(n_1653),
.B2(n_1647),
.C(n_1676),
.Y(n_1739)
);

HB1xp67_ASAP7_75t_L g1740 ( 
.A(n_1721),
.Y(n_1740)
);

OR2x6_ASAP7_75t_L g1741 ( 
.A(n_1704),
.B(n_1699),
.Y(n_1741)
);

AND2x2_ASAP7_75t_L g1742 ( 
.A(n_1728),
.B(n_1658),
.Y(n_1742)
);

BUFx2_ASAP7_75t_L g1743 ( 
.A(n_1729),
.Y(n_1743)
);

AND2x4_ASAP7_75t_L g1744 ( 
.A(n_1724),
.B(n_1690),
.Y(n_1744)
);

AOI22xp33_ASAP7_75t_L g1745 ( 
.A1(n_1727),
.A2(n_1653),
.B1(n_1688),
.B2(n_1683),
.Y(n_1745)
);

INVx1_ASAP7_75t_L g1746 ( 
.A(n_1711),
.Y(n_1746)
);

OAI21xp33_ASAP7_75t_L g1747 ( 
.A1(n_1722),
.A2(n_1677),
.B(n_1699),
.Y(n_1747)
);

HB1xp67_ASAP7_75t_L g1748 ( 
.A(n_1721),
.Y(n_1748)
);

AOI22xp33_ASAP7_75t_L g1749 ( 
.A1(n_1703),
.A2(n_1653),
.B1(n_1683),
.B2(n_1647),
.Y(n_1749)
);

OR2x2_ASAP7_75t_L g1750 ( 
.A(n_1706),
.B(n_1723),
.Y(n_1750)
);

INVx1_ASAP7_75t_L g1751 ( 
.A(n_1715),
.Y(n_1751)
);

OA21x2_ASAP7_75t_L g1752 ( 
.A1(n_1725),
.A2(n_1714),
.B(n_1719),
.Y(n_1752)
);

OAI211xp5_ASAP7_75t_L g1753 ( 
.A1(n_1703),
.A2(n_1657),
.B(n_1682),
.C(n_1567),
.Y(n_1753)
);

AOI33xp33_ASAP7_75t_L g1754 ( 
.A1(n_1722),
.A2(n_1656),
.A3(n_1652),
.B1(n_1659),
.B2(n_1700),
.B3(n_1669),
.Y(n_1754)
);

OAI22xp5_ASAP7_75t_L g1755 ( 
.A1(n_1732),
.A2(n_1683),
.B1(n_1662),
.B2(n_1676),
.Y(n_1755)
);

HB1xp67_ASAP7_75t_L g1756 ( 
.A(n_1729),
.Y(n_1756)
);

AOI22xp33_ASAP7_75t_L g1757 ( 
.A1(n_1703),
.A2(n_1693),
.B1(n_1696),
.B2(n_1686),
.Y(n_1757)
);

BUFx2_ASAP7_75t_L g1758 ( 
.A(n_1705),
.Y(n_1758)
);

AOI33xp33_ASAP7_75t_L g1759 ( 
.A1(n_1722),
.A2(n_1652),
.A3(n_1671),
.B1(n_1675),
.B2(n_1674),
.B3(n_1670),
.Y(n_1759)
);

OAI22xp5_ASAP7_75t_L g1760 ( 
.A1(n_1732),
.A2(n_1662),
.B1(n_1691),
.B2(n_1690),
.Y(n_1760)
);

AOI22xp33_ASAP7_75t_L g1761 ( 
.A1(n_1703),
.A2(n_1693),
.B1(n_1696),
.B2(n_1686),
.Y(n_1761)
);

NAND4xp25_ASAP7_75t_L g1762 ( 
.A(n_1719),
.B(n_1677),
.C(n_1694),
.D(n_1684),
.Y(n_1762)
);

AOI22xp5_ASAP7_75t_L g1763 ( 
.A1(n_1707),
.A2(n_1663),
.B1(n_1687),
.B2(n_1698),
.Y(n_1763)
);

BUFx3_ASAP7_75t_L g1764 ( 
.A(n_1718),
.Y(n_1764)
);

INVxp67_ASAP7_75t_L g1765 ( 
.A(n_1701),
.Y(n_1765)
);

OAI33xp33_ASAP7_75t_L g1766 ( 
.A1(n_1701),
.A2(n_1706),
.A3(n_1680),
.B1(n_1672),
.B2(n_1675),
.B3(n_1674),
.Y(n_1766)
);

HB1xp67_ASAP7_75t_L g1767 ( 
.A(n_1756),
.Y(n_1767)
);

AND2x2_ASAP7_75t_L g1768 ( 
.A(n_1758),
.B(n_1709),
.Y(n_1768)
);

INVx1_ASAP7_75t_L g1769 ( 
.A(n_1734),
.Y(n_1769)
);

AND2x4_ASAP7_75t_L g1770 ( 
.A(n_1764),
.B(n_1726),
.Y(n_1770)
);

OA21x2_ASAP7_75t_L g1771 ( 
.A1(n_1757),
.A2(n_1719),
.B(n_1726),
.Y(n_1771)
);

BUFx3_ASAP7_75t_L g1772 ( 
.A(n_1764),
.Y(n_1772)
);

OR2x2_ASAP7_75t_L g1773 ( 
.A(n_1750),
.B(n_1706),
.Y(n_1773)
);

INVx1_ASAP7_75t_L g1774 ( 
.A(n_1738),
.Y(n_1774)
);

AND2x6_ASAP7_75t_SL g1775 ( 
.A(n_1741),
.B(n_1551),
.Y(n_1775)
);

INVx1_ASAP7_75t_L g1776 ( 
.A(n_1746),
.Y(n_1776)
);

INVx1_ASAP7_75t_L g1777 ( 
.A(n_1751),
.Y(n_1777)
);

BUFx2_ASAP7_75t_L g1778 ( 
.A(n_1740),
.Y(n_1778)
);

OA21x2_ASAP7_75t_L g1779 ( 
.A1(n_1757),
.A2(n_1717),
.B(n_1713),
.Y(n_1779)
);

AND2x2_ASAP7_75t_L g1780 ( 
.A(n_1754),
.B(n_1709),
.Y(n_1780)
);

BUFx8_ASAP7_75t_L g1781 ( 
.A(n_1743),
.Y(n_1781)
);

HB1xp67_ASAP7_75t_L g1782 ( 
.A(n_1748),
.Y(n_1782)
);

HB1xp67_ASAP7_75t_L g1783 ( 
.A(n_1765),
.Y(n_1783)
);

INVx4_ASAP7_75t_L g1784 ( 
.A(n_1741),
.Y(n_1784)
);

NOR3xp33_ASAP7_75t_SL g1785 ( 
.A(n_1753),
.B(n_1627),
.C(n_1579),
.Y(n_1785)
);

NAND2xp5_ASAP7_75t_L g1786 ( 
.A(n_1759),
.B(n_1716),
.Y(n_1786)
);

AO21x1_ASAP7_75t_L g1787 ( 
.A1(n_1755),
.A2(n_1701),
.B(n_1716),
.Y(n_1787)
);

INVx1_ASAP7_75t_L g1788 ( 
.A(n_1759),
.Y(n_1788)
);

OAI21x1_ASAP7_75t_L g1789 ( 
.A1(n_1761),
.A2(n_1664),
.B(n_1684),
.Y(n_1789)
);

NAND2xp5_ASAP7_75t_L g1790 ( 
.A(n_1754),
.B(n_1716),
.Y(n_1790)
);

INVx1_ASAP7_75t_L g1791 ( 
.A(n_1735),
.Y(n_1791)
);

OR2x2_ASAP7_75t_L g1792 ( 
.A(n_1737),
.B(n_1720),
.Y(n_1792)
);

AND2x2_ASAP7_75t_L g1793 ( 
.A(n_1742),
.B(n_1710),
.Y(n_1793)
);

NAND2xp5_ASAP7_75t_L g1794 ( 
.A(n_1752),
.B(n_1712),
.Y(n_1794)
);

INVx2_ASAP7_75t_L g1795 ( 
.A(n_1771),
.Y(n_1795)
);

OR2x2_ASAP7_75t_L g1796 ( 
.A(n_1773),
.B(n_1762),
.Y(n_1796)
);

INVx2_ASAP7_75t_L g1797 ( 
.A(n_1771),
.Y(n_1797)
);

INVx1_ASAP7_75t_SL g1798 ( 
.A(n_1772),
.Y(n_1798)
);

OR2x2_ASAP7_75t_L g1799 ( 
.A(n_1773),
.B(n_1752),
.Y(n_1799)
);

OAI33xp33_ASAP7_75t_L g1800 ( 
.A1(n_1788),
.A2(n_1747),
.A3(n_1760),
.B1(n_1720),
.B2(n_1671),
.B3(n_1672),
.Y(n_1800)
);

INVx1_ASAP7_75t_L g1801 ( 
.A(n_1769),
.Y(n_1801)
);

AND2x2_ASAP7_75t_L g1802 ( 
.A(n_1780),
.B(n_1736),
.Y(n_1802)
);

AOI22xp5_ASAP7_75t_L g1803 ( 
.A1(n_1771),
.A2(n_1707),
.B1(n_1745),
.B2(n_1761),
.Y(n_1803)
);

INVx2_ASAP7_75t_L g1804 ( 
.A(n_1771),
.Y(n_1804)
);

OR2x2_ASAP7_75t_L g1805 ( 
.A(n_1788),
.B(n_1752),
.Y(n_1805)
);

INVx5_ASAP7_75t_L g1806 ( 
.A(n_1775),
.Y(n_1806)
);

INVx4_ASAP7_75t_L g1807 ( 
.A(n_1772),
.Y(n_1807)
);

INVx2_ASAP7_75t_L g1808 ( 
.A(n_1779),
.Y(n_1808)
);

AND2x2_ASAP7_75t_L g1809 ( 
.A(n_1772),
.B(n_1744),
.Y(n_1809)
);

INVx1_ASAP7_75t_L g1810 ( 
.A(n_1769),
.Y(n_1810)
);

AND2x2_ASAP7_75t_L g1811 ( 
.A(n_1793),
.B(n_1744),
.Y(n_1811)
);

INVx3_ASAP7_75t_L g1812 ( 
.A(n_1779),
.Y(n_1812)
);

INVx6_ASAP7_75t_L g1813 ( 
.A(n_1781),
.Y(n_1813)
);

INVx1_ASAP7_75t_SL g1814 ( 
.A(n_1783),
.Y(n_1814)
);

OR2x4_ASAP7_75t_L g1815 ( 
.A(n_1786),
.B(n_1790),
.Y(n_1815)
);

AND2x2_ASAP7_75t_SL g1816 ( 
.A(n_1779),
.B(n_1749),
.Y(n_1816)
);

NAND2xp5_ASAP7_75t_L g1817 ( 
.A(n_1791),
.B(n_1763),
.Y(n_1817)
);

INVx2_ASAP7_75t_SL g1818 ( 
.A(n_1781),
.Y(n_1818)
);

OR2x2_ASAP7_75t_L g1819 ( 
.A(n_1792),
.B(n_1712),
.Y(n_1819)
);

INVx2_ASAP7_75t_L g1820 ( 
.A(n_1779),
.Y(n_1820)
);

AOI22xp33_ASAP7_75t_SL g1821 ( 
.A1(n_1787),
.A2(n_1739),
.B1(n_1718),
.B2(n_1730),
.Y(n_1821)
);

INVxp67_ASAP7_75t_SL g1822 ( 
.A(n_1781),
.Y(n_1822)
);

INVx1_ASAP7_75t_L g1823 ( 
.A(n_1774),
.Y(n_1823)
);

INVx1_ASAP7_75t_L g1824 ( 
.A(n_1801),
.Y(n_1824)
);

NOR2xp33_ASAP7_75t_L g1825 ( 
.A(n_1813),
.B(n_1733),
.Y(n_1825)
);

INVxp67_ASAP7_75t_L g1826 ( 
.A(n_1822),
.Y(n_1826)
);

XOR2x2_ASAP7_75t_L g1827 ( 
.A(n_1803),
.B(n_1745),
.Y(n_1827)
);

AOI22xp33_ASAP7_75t_SL g1828 ( 
.A1(n_1795),
.A2(n_1789),
.B1(n_1787),
.B2(n_1784),
.Y(n_1828)
);

INVx2_ASAP7_75t_L g1829 ( 
.A(n_1812),
.Y(n_1829)
);

NAND2xp5_ASAP7_75t_L g1830 ( 
.A(n_1814),
.B(n_1791),
.Y(n_1830)
);

INVx1_ASAP7_75t_L g1831 ( 
.A(n_1801),
.Y(n_1831)
);

INVx1_ASAP7_75t_L g1832 ( 
.A(n_1810),
.Y(n_1832)
);

AND2x2_ASAP7_75t_L g1833 ( 
.A(n_1809),
.B(n_1778),
.Y(n_1833)
);

INVx2_ASAP7_75t_L g1834 ( 
.A(n_1812),
.Y(n_1834)
);

INVx1_ASAP7_75t_L g1835 ( 
.A(n_1810),
.Y(n_1835)
);

NAND2xp5_ASAP7_75t_L g1836 ( 
.A(n_1798),
.B(n_1778),
.Y(n_1836)
);

AND2x2_ASAP7_75t_L g1837 ( 
.A(n_1809),
.B(n_1782),
.Y(n_1837)
);

AOI21xp5_ASAP7_75t_L g1838 ( 
.A1(n_1800),
.A2(n_1766),
.B(n_1794),
.Y(n_1838)
);

NAND2x1_ASAP7_75t_L g1839 ( 
.A(n_1812),
.B(n_1770),
.Y(n_1839)
);

OR2x2_ASAP7_75t_L g1840 ( 
.A(n_1805),
.B(n_1767),
.Y(n_1840)
);

NAND2xp5_ASAP7_75t_L g1841 ( 
.A(n_1817),
.B(n_1776),
.Y(n_1841)
);

AND2x2_ASAP7_75t_L g1842 ( 
.A(n_1802),
.B(n_1768),
.Y(n_1842)
);

AND2x2_ASAP7_75t_L g1843 ( 
.A(n_1802),
.B(n_1768),
.Y(n_1843)
);

OR2x2_ASAP7_75t_L g1844 ( 
.A(n_1805),
.B(n_1794),
.Y(n_1844)
);

AOI221xp5_ASAP7_75t_L g1845 ( 
.A1(n_1795),
.A2(n_1797),
.B1(n_1804),
.B2(n_1803),
.C(n_1808),
.Y(n_1845)
);

NOR2xp67_ASAP7_75t_L g1846 ( 
.A(n_1806),
.B(n_1784),
.Y(n_1846)
);

INVx1_ASAP7_75t_L g1847 ( 
.A(n_1823),
.Y(n_1847)
);

AND2x2_ASAP7_75t_L g1848 ( 
.A(n_1811),
.B(n_1785),
.Y(n_1848)
);

INVx1_ASAP7_75t_L g1849 ( 
.A(n_1823),
.Y(n_1849)
);

INVx1_ASAP7_75t_SL g1850 ( 
.A(n_1813),
.Y(n_1850)
);

NAND2x1p5_ASAP7_75t_L g1851 ( 
.A(n_1806),
.B(n_1784),
.Y(n_1851)
);

INVx1_ASAP7_75t_SL g1852 ( 
.A(n_1813),
.Y(n_1852)
);

AND2x2_ASAP7_75t_L g1853 ( 
.A(n_1811),
.B(n_1776),
.Y(n_1853)
);

NAND2xp5_ASAP7_75t_L g1854 ( 
.A(n_1806),
.B(n_1777),
.Y(n_1854)
);

INVx1_ASAP7_75t_SL g1855 ( 
.A(n_1850),
.Y(n_1855)
);

NAND2xp5_ASAP7_75t_L g1856 ( 
.A(n_1838),
.B(n_1815),
.Y(n_1856)
);

NOR2xp33_ASAP7_75t_L g1857 ( 
.A(n_1852),
.B(n_1825),
.Y(n_1857)
);

BUFx12f_ASAP7_75t_L g1858 ( 
.A(n_1851),
.Y(n_1858)
);

HB1xp67_ASAP7_75t_L g1859 ( 
.A(n_1826),
.Y(n_1859)
);

INVx1_ASAP7_75t_SL g1860 ( 
.A(n_1851),
.Y(n_1860)
);

INVx2_ASAP7_75t_L g1861 ( 
.A(n_1829),
.Y(n_1861)
);

INVx2_ASAP7_75t_L g1862 ( 
.A(n_1829),
.Y(n_1862)
);

INVx1_ASAP7_75t_L g1863 ( 
.A(n_1824),
.Y(n_1863)
);

AOI21xp5_ASAP7_75t_L g1864 ( 
.A1(n_1828),
.A2(n_1806),
.B(n_1804),
.Y(n_1864)
);

OA22x2_ASAP7_75t_L g1865 ( 
.A1(n_1841),
.A2(n_1797),
.B1(n_1808),
.B2(n_1820),
.Y(n_1865)
);

INVx3_ASAP7_75t_L g1866 ( 
.A(n_1839),
.Y(n_1866)
);

INVx2_ASAP7_75t_L g1867 ( 
.A(n_1834),
.Y(n_1867)
);

OR2x2_ASAP7_75t_L g1868 ( 
.A(n_1840),
.B(n_1819),
.Y(n_1868)
);

INVx2_ASAP7_75t_L g1869 ( 
.A(n_1834),
.Y(n_1869)
);

INVx1_ASAP7_75t_L g1870 ( 
.A(n_1831),
.Y(n_1870)
);

INVx2_ASAP7_75t_L g1871 ( 
.A(n_1827),
.Y(n_1871)
);

AOI22xp33_ASAP7_75t_L g1872 ( 
.A1(n_1827),
.A2(n_1806),
.B1(n_1816),
.B2(n_1821),
.Y(n_1872)
);

HB1xp67_ASAP7_75t_L g1873 ( 
.A(n_1833),
.Y(n_1873)
);

NAND2xp5_ASAP7_75t_L g1874 ( 
.A(n_1845),
.B(n_1815),
.Y(n_1874)
);

INVx1_ASAP7_75t_L g1875 ( 
.A(n_1832),
.Y(n_1875)
);

HB1xp67_ASAP7_75t_L g1876 ( 
.A(n_1833),
.Y(n_1876)
);

INVxp67_ASAP7_75t_L g1877 ( 
.A(n_1825),
.Y(n_1877)
);

INVx3_ASAP7_75t_L g1878 ( 
.A(n_1839),
.Y(n_1878)
);

INVx2_ASAP7_75t_L g1879 ( 
.A(n_1840),
.Y(n_1879)
);

INVx3_ASAP7_75t_L g1880 ( 
.A(n_1851),
.Y(n_1880)
);

INVxp67_ASAP7_75t_L g1881 ( 
.A(n_1836),
.Y(n_1881)
);

INVx2_ASAP7_75t_L g1882 ( 
.A(n_1866),
.Y(n_1882)
);

AND2x2_ASAP7_75t_L g1883 ( 
.A(n_1873),
.B(n_1837),
.Y(n_1883)
);

NAND2xp5_ASAP7_75t_L g1884 ( 
.A(n_1876),
.B(n_1837),
.Y(n_1884)
);

INVx1_ASAP7_75t_L g1885 ( 
.A(n_1859),
.Y(n_1885)
);

AOI221xp5_ASAP7_75t_L g1886 ( 
.A1(n_1874),
.A2(n_1820),
.B1(n_1844),
.B2(n_1799),
.C(n_1806),
.Y(n_1886)
);

NAND2xp5_ASAP7_75t_L g1887 ( 
.A(n_1855),
.B(n_1853),
.Y(n_1887)
);

INVx1_ASAP7_75t_L g1888 ( 
.A(n_1879),
.Y(n_1888)
);

NOR4xp25_ASAP7_75t_L g1889 ( 
.A(n_1874),
.B(n_1856),
.C(n_1855),
.D(n_1871),
.Y(n_1889)
);

NAND2xp5_ASAP7_75t_SL g1890 ( 
.A(n_1864),
.B(n_1846),
.Y(n_1890)
);

OAI22xp5_ASAP7_75t_L g1891 ( 
.A1(n_1872),
.A2(n_1815),
.B1(n_1813),
.B2(n_1796),
.Y(n_1891)
);

OAI32xp33_ASAP7_75t_L g1892 ( 
.A1(n_1856),
.A2(n_1844),
.A3(n_1799),
.B1(n_1796),
.B2(n_1854),
.Y(n_1892)
);

AOI21xp33_ASAP7_75t_L g1893 ( 
.A1(n_1865),
.A2(n_1816),
.B(n_1835),
.Y(n_1893)
);

OAI21xp5_ASAP7_75t_L g1894 ( 
.A1(n_1864),
.A2(n_1816),
.B(n_1830),
.Y(n_1894)
);

NOR2xp33_ASAP7_75t_L g1895 ( 
.A(n_1877),
.B(n_1818),
.Y(n_1895)
);

INVx1_ASAP7_75t_L g1896 ( 
.A(n_1879),
.Y(n_1896)
);

NAND2xp5_ASAP7_75t_L g1897 ( 
.A(n_1879),
.B(n_1853),
.Y(n_1897)
);

INVxp67_ASAP7_75t_L g1898 ( 
.A(n_1857),
.Y(n_1898)
);

NAND2xp5_ASAP7_75t_L g1899 ( 
.A(n_1881),
.B(n_1842),
.Y(n_1899)
);

OAI21xp33_ASAP7_75t_SL g1900 ( 
.A1(n_1865),
.A2(n_1843),
.B(n_1842),
.Y(n_1900)
);

NAND2xp5_ASAP7_75t_L g1901 ( 
.A(n_1881),
.B(n_1843),
.Y(n_1901)
);

INVx1_ASAP7_75t_SL g1902 ( 
.A(n_1858),
.Y(n_1902)
);

NAND2xp5_ASAP7_75t_L g1903 ( 
.A(n_1868),
.B(n_1807),
.Y(n_1903)
);

INVx1_ASAP7_75t_SL g1904 ( 
.A(n_1883),
.Y(n_1904)
);

INVx1_ASAP7_75t_L g1905 ( 
.A(n_1888),
.Y(n_1905)
);

AOI22xp33_ASAP7_75t_L g1906 ( 
.A1(n_1893),
.A2(n_1871),
.B1(n_1865),
.B2(n_1861),
.Y(n_1906)
);

INVx1_ASAP7_75t_SL g1907 ( 
.A(n_1887),
.Y(n_1907)
);

NAND2xp5_ASAP7_75t_L g1908 ( 
.A(n_1889),
.B(n_1868),
.Y(n_1908)
);

INVx1_ASAP7_75t_L g1909 ( 
.A(n_1896),
.Y(n_1909)
);

INVx1_ASAP7_75t_L g1910 ( 
.A(n_1897),
.Y(n_1910)
);

HB1xp67_ASAP7_75t_L g1911 ( 
.A(n_1882),
.Y(n_1911)
);

NAND2xp5_ASAP7_75t_L g1912 ( 
.A(n_1898),
.B(n_1861),
.Y(n_1912)
);

AND2x2_ASAP7_75t_L g1913 ( 
.A(n_1898),
.B(n_1848),
.Y(n_1913)
);

NOR2xp33_ASAP7_75t_L g1914 ( 
.A(n_1902),
.B(n_1818),
.Y(n_1914)
);

INVx1_ASAP7_75t_L g1915 ( 
.A(n_1885),
.Y(n_1915)
);

INVx2_ASAP7_75t_L g1916 ( 
.A(n_1884),
.Y(n_1916)
);

INVx1_ASAP7_75t_SL g1917 ( 
.A(n_1904),
.Y(n_1917)
);

NAND2xp5_ASAP7_75t_SL g1918 ( 
.A(n_1908),
.B(n_1894),
.Y(n_1918)
);

NAND2xp5_ASAP7_75t_L g1919 ( 
.A(n_1913),
.B(n_1899),
.Y(n_1919)
);

NOR4xp25_ASAP7_75t_L g1920 ( 
.A(n_1906),
.B(n_1900),
.C(n_1890),
.D(n_1871),
.Y(n_1920)
);

AOI21xp5_ASAP7_75t_L g1921 ( 
.A1(n_1912),
.A2(n_1890),
.B(n_1892),
.Y(n_1921)
);

AOI311xp33_ASAP7_75t_L g1922 ( 
.A1(n_1915),
.A2(n_1895),
.A3(n_1891),
.B(n_1901),
.C(n_1886),
.Y(n_1922)
);

AOI211xp5_ASAP7_75t_L g1923 ( 
.A1(n_1907),
.A2(n_1860),
.B(n_1895),
.C(n_1903),
.Y(n_1923)
);

NAND2xp5_ASAP7_75t_L g1924 ( 
.A(n_1913),
.B(n_1863),
.Y(n_1924)
);

NOR3xp33_ASAP7_75t_L g1925 ( 
.A(n_1916),
.B(n_1860),
.C(n_1880),
.Y(n_1925)
);

OAI21xp33_ASAP7_75t_L g1926 ( 
.A1(n_1914),
.A2(n_1862),
.B(n_1861),
.Y(n_1926)
);

O2A1O1Ixp33_ASAP7_75t_L g1927 ( 
.A1(n_1911),
.A2(n_1880),
.B(n_1862),
.C(n_1867),
.Y(n_1927)
);

AOI21xp5_ASAP7_75t_L g1928 ( 
.A1(n_1918),
.A2(n_1905),
.B(n_1909),
.Y(n_1928)
);

OAI21xp33_ASAP7_75t_L g1929 ( 
.A1(n_1920),
.A2(n_1916),
.B(n_1910),
.Y(n_1929)
);

INVx1_ASAP7_75t_L g1930 ( 
.A(n_1924),
.Y(n_1930)
);

INVx1_ASAP7_75t_L g1931 ( 
.A(n_1917),
.Y(n_1931)
);

NAND2xp5_ASAP7_75t_L g1932 ( 
.A(n_1921),
.B(n_1910),
.Y(n_1932)
);

AOI322xp5_ASAP7_75t_L g1933 ( 
.A1(n_1926),
.A2(n_1905),
.A3(n_1862),
.B1(n_1869),
.B2(n_1867),
.C1(n_1875),
.C2(n_1870),
.Y(n_1933)
);

INVx2_ASAP7_75t_L g1934 ( 
.A(n_1919),
.Y(n_1934)
);

NAND2xp5_ASAP7_75t_L g1935 ( 
.A(n_1934),
.B(n_1925),
.Y(n_1935)
);

INVx1_ASAP7_75t_L g1936 ( 
.A(n_1931),
.Y(n_1936)
);

NAND2xp5_ASAP7_75t_L g1937 ( 
.A(n_1928),
.B(n_1923),
.Y(n_1937)
);

INVx1_ASAP7_75t_L g1938 ( 
.A(n_1930),
.Y(n_1938)
);

INVxp67_ASAP7_75t_L g1939 ( 
.A(n_1932),
.Y(n_1939)
);

INVxp67_ASAP7_75t_L g1940 ( 
.A(n_1929),
.Y(n_1940)
);

INVx1_ASAP7_75t_L g1941 ( 
.A(n_1933),
.Y(n_1941)
);

O2A1O1Ixp33_ASAP7_75t_L g1942 ( 
.A1(n_1940),
.A2(n_1927),
.B(n_1880),
.C(n_1922),
.Y(n_1942)
);

AOI21xp5_ASAP7_75t_L g1943 ( 
.A1(n_1937),
.A2(n_1880),
.B(n_1869),
.Y(n_1943)
);

INVx3_ASAP7_75t_L g1944 ( 
.A(n_1936),
.Y(n_1944)
);

NOR2xp33_ASAP7_75t_R g1945 ( 
.A(n_1938),
.B(n_1858),
.Y(n_1945)
);

HB1xp67_ASAP7_75t_L g1946 ( 
.A(n_1939),
.Y(n_1946)
);

AND2x2_ASAP7_75t_L g1947 ( 
.A(n_1946),
.B(n_1944),
.Y(n_1947)
);

BUFx2_ASAP7_75t_L g1948 ( 
.A(n_1945),
.Y(n_1948)
);

AND2x2_ASAP7_75t_SL g1949 ( 
.A(n_1942),
.B(n_1941),
.Y(n_1949)
);

INVx1_ASAP7_75t_L g1950 ( 
.A(n_1947),
.Y(n_1950)
);

NOR2xp33_ASAP7_75t_L g1951 ( 
.A(n_1950),
.B(n_1935),
.Y(n_1951)
);

INVx1_ASAP7_75t_L g1952 ( 
.A(n_1951),
.Y(n_1952)
);

AOI22xp5_ASAP7_75t_SL g1953 ( 
.A1(n_1951),
.A2(n_1948),
.B1(n_1943),
.B2(n_1949),
.Y(n_1953)
);

AOI22xp33_ASAP7_75t_L g1954 ( 
.A1(n_1952),
.A2(n_1949),
.B1(n_1869),
.B2(n_1867),
.Y(n_1954)
);

OAI22xp33_ASAP7_75t_L g1955 ( 
.A1(n_1953),
.A2(n_1858),
.B1(n_1875),
.B2(n_1870),
.Y(n_1955)
);

HB1xp67_ASAP7_75t_L g1956 ( 
.A(n_1954),
.Y(n_1956)
);

NOR2xp33_ASAP7_75t_L g1957 ( 
.A(n_1955),
.B(n_1863),
.Y(n_1957)
);

XOR2xp5_ASAP7_75t_L g1958 ( 
.A(n_1956),
.B(n_1733),
.Y(n_1958)
);

XOR2xp5_ASAP7_75t_L g1959 ( 
.A(n_1958),
.B(n_1957),
.Y(n_1959)
);

OR2x6_ASAP7_75t_L g1960 ( 
.A(n_1959),
.B(n_1807),
.Y(n_1960)
);

XNOR2xp5_ASAP7_75t_L g1961 ( 
.A(n_1960),
.B(n_1678),
.Y(n_1961)
);

AOI221xp5_ASAP7_75t_L g1962 ( 
.A1(n_1961),
.A2(n_1878),
.B1(n_1866),
.B2(n_1807),
.C(n_1847),
.Y(n_1962)
);

AOI211xp5_ASAP7_75t_L g1963 ( 
.A1(n_1962),
.A2(n_1878),
.B(n_1866),
.C(n_1849),
.Y(n_1963)
);


endmodule