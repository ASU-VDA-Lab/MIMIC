module real_jpeg_25094_n_16 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_3, n_10, n_356, n_9, n_16);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_3;
input n_10;
input n_356;
input n_9;

output n_16;

wire n_37;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_300;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_199;
wire n_95;
wire n_238;
wire n_67;
wire n_350;
wire n_235;
wire n_107;
wire n_354;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_123;
wire n_50;
wire n_186;
wire n_137;
wire n_72;
wire n_171;
wire n_151;
wire n_272;
wire n_198;
wire n_203;
wire n_23;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_326;
wire n_339;
wire n_80;
wire n_30;
wire n_332;
wire n_149;
wire n_328;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_353;
wire n_230;
wire n_128;
wire n_202;
wire n_216;
wire n_127;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_348;
wire n_252;
wire n_310;
wire n_345;
wire n_78;
wire n_288;
wire n_83;
wire n_221;
wire n_104;
wire n_153;
wire n_337;
wire n_131;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_200;
wire n_335;
wire n_214;
wire n_113;
wire n_251;
wire n_139;
wire n_33;
wire n_175;
wire n_338;
wire n_156;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_77;
wire n_219;
wire n_122;
wire n_19;
wire n_262;
wire n_334;
wire n_17;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_20;
wire n_278;
wire n_314;
wire n_103;
wire n_232;
wire n_212;
wire n_284;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_213;
wire n_25;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_341;
wire n_331;
wire n_49;
wire n_68;
wire n_146;
wire n_286;
wire n_323;
wire n_166;
wire n_176;
wire n_215;
wire n_312;
wire n_325;
wire n_307;
wire n_316;
wire n_161;
wire n_207;
wire n_237;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_140;
wire n_126;
wire n_342;
wire n_120;
wire n_155;
wire n_319;
wire n_93;
wire n_242;
wire n_142;
wire n_76;
wire n_79;
wire n_282;
wire n_147;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_18;
wire n_145;
wire n_266;
wire n_109;
wire n_148;
wire n_196;
wire n_298;
wire n_330;
wire n_333;
wire n_152;
wire n_270;
wire n_159;
wire n_347;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_336;
wire n_258;
wire n_150;
wire n_41;
wire n_74;
wire n_158;
wire n_204;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_75;
wire n_346;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_119;
wire n_283;
wire n_181;
wire n_256;
wire n_273;
wire n_253;
wire n_54;
wire n_168;
wire n_38;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_349;
wire n_292;
wire n_343;
wire n_64;
wire n_291;
wire n_236;
wire n_276;
wire n_287;
wire n_174;
wire n_255;
wire n_299;
wire n_243;
wire n_352;
wire n_56;
wire n_293;
wire n_275;
wire n_227;
wire n_229;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_45;
wire n_268;
wire n_42;
wire n_313;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_143;
wire n_351;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_303;
wire n_321;
wire n_100;
wire n_51;
wire n_205;
wire n_324;
wire n_86;
wire n_261;
wire n_70;
wire n_32;
wire n_228;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_133;
wire n_257;
wire n_344;
wire n_210;
wire n_206;
wire n_85;
wire n_96;
wire n_308;

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_0),
.Y(n_68)
);

OAI22xp5_ASAP7_75t_L g77 ( 
.A1(n_1),
.A2(n_67),
.B1(n_70),
.B2(n_78),
.Y(n_77)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_1),
.Y(n_78)
);

AOI22xp33_ASAP7_75t_L g156 ( 
.A1(n_1),
.A2(n_30),
.B1(n_33),
.B2(n_78),
.Y(n_156)
);

OAI22xp5_ASAP7_75t_L g198 ( 
.A1(n_1),
.A2(n_47),
.B1(n_48),
.B2(n_78),
.Y(n_198)
);

OAI22xp5_ASAP7_75t_L g232 ( 
.A1(n_1),
.A2(n_78),
.B1(n_93),
.B2(n_94),
.Y(n_232)
);

BUFx12f_ASAP7_75t_L g45 ( 
.A(n_2),
.Y(n_45)
);

BUFx10_ASAP7_75t_L g30 ( 
.A(n_3),
.Y(n_30)
);

INVx8_ASAP7_75t_SL g91 ( 
.A(n_4),
.Y(n_91)
);

AOI22xp33_ASAP7_75t_SL g46 ( 
.A1(n_5),
.A2(n_47),
.B1(n_48),
.B2(n_50),
.Y(n_46)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_5),
.Y(n_50)
);

OAI22xp5_ASAP7_75t_L g114 ( 
.A1(n_5),
.A2(n_30),
.B1(n_33),
.B2(n_50),
.Y(n_114)
);

AOI22xp33_ASAP7_75t_SL g267 ( 
.A1(n_5),
.A2(n_50),
.B1(n_67),
.B2(n_70),
.Y(n_267)
);

AOI22xp33_ASAP7_75t_SL g305 ( 
.A1(n_5),
.A2(n_50),
.B1(n_84),
.B2(n_94),
.Y(n_305)
);

OAI22xp33_ASAP7_75t_SL g61 ( 
.A1(n_6),
.A2(n_47),
.B1(n_48),
.B2(n_62),
.Y(n_61)
);

CKINVDCx20_ASAP7_75t_R g62 ( 
.A(n_6),
.Y(n_62)
);

OAI22xp5_ASAP7_75t_SL g110 ( 
.A1(n_6),
.A2(n_62),
.B1(n_67),
.B2(n_70),
.Y(n_110)
);

OAI22xp5_ASAP7_75t_SL g159 ( 
.A1(n_6),
.A2(n_30),
.B1(n_33),
.B2(n_62),
.Y(n_159)
);

OAI22xp5_ASAP7_75t_SL g265 ( 
.A1(n_6),
.A2(n_62),
.B1(n_84),
.B2(n_87),
.Y(n_265)
);

CKINVDCx20_ASAP7_75t_R g85 ( 
.A(n_7),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_L g130 ( 
.A(n_7),
.B(n_95),
.Y(n_130)
);

MAJIxp5_ASAP7_75t_L g143 ( 
.A(n_7),
.B(n_30),
.C(n_44),
.Y(n_143)
);

AOI22xp5_ASAP7_75t_L g146 ( 
.A1(n_7),
.A2(n_47),
.B1(n_48),
.B2(n_85),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_L g151 ( 
.A(n_7),
.B(n_76),
.Y(n_151)
);

OAI22xp5_ASAP7_75t_SL g171 ( 
.A1(n_7),
.A2(n_29),
.B1(n_172),
.B2(n_173),
.Y(n_171)
);

BUFx12f_ASAP7_75t_L g73 ( 
.A(n_8),
.Y(n_73)
);

INVx13_ASAP7_75t_L g84 ( 
.A(n_9),
.Y(n_84)
);

AOI22xp33_ASAP7_75t_L g97 ( 
.A1(n_10),
.A2(n_81),
.B1(n_93),
.B2(n_98),
.Y(n_97)
);

CKINVDCx20_ASAP7_75t_R g98 ( 
.A(n_10),
.Y(n_98)
);

OAI22xp5_ASAP7_75t_L g127 ( 
.A1(n_10),
.A2(n_67),
.B1(n_70),
.B2(n_98),
.Y(n_127)
);

AOI22xp5_ASAP7_75t_L g147 ( 
.A1(n_10),
.A2(n_47),
.B1(n_48),
.B2(n_98),
.Y(n_147)
);

AOI22xp5_ASAP7_75t_SL g172 ( 
.A1(n_10),
.A2(n_30),
.B1(n_33),
.B2(n_98),
.Y(n_172)
);

OAI22xp5_ASAP7_75t_SL g66 ( 
.A1(n_11),
.A2(n_67),
.B1(n_69),
.B2(n_70),
.Y(n_66)
);

CKINVDCx20_ASAP7_75t_R g69 ( 
.A(n_11),
.Y(n_69)
);

OAI22xp33_ASAP7_75t_SL g105 ( 
.A1(n_11),
.A2(n_69),
.B1(n_84),
.B2(n_94),
.Y(n_105)
);

AOI22xp33_ASAP7_75t_L g154 ( 
.A1(n_11),
.A2(n_47),
.B1(n_48),
.B2(n_69),
.Y(n_154)
);

AOI22xp33_ASAP7_75t_L g165 ( 
.A1(n_11),
.A2(n_30),
.B1(n_33),
.B2(n_69),
.Y(n_165)
);

BUFx12f_ASAP7_75t_L g49 ( 
.A(n_12),
.Y(n_49)
);

AOI22xp33_ASAP7_75t_L g39 ( 
.A1(n_13),
.A2(n_30),
.B1(n_33),
.B2(n_40),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_13),
.Y(n_40)
);

OAI22xp33_ASAP7_75t_SL g52 ( 
.A1(n_13),
.A2(n_40),
.B1(n_47),
.B2(n_48),
.Y(n_52)
);

OAI22xp5_ASAP7_75t_L g237 ( 
.A1(n_13),
.A2(n_40),
.B1(n_67),
.B2(n_70),
.Y(n_237)
);

OAI22xp33_ASAP7_75t_L g286 ( 
.A1(n_13),
.A2(n_40),
.B1(n_287),
.B2(n_288),
.Y(n_286)
);

AOI22xp33_ASAP7_75t_L g32 ( 
.A1(n_14),
.A2(n_30),
.B1(n_33),
.B2(n_34),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_14),
.Y(n_34)
);

AOI22xp5_ASAP7_75t_SL g244 ( 
.A1(n_14),
.A2(n_34),
.B1(n_47),
.B2(n_48),
.Y(n_244)
);

AOI22xp33_ASAP7_75t_L g296 ( 
.A1(n_14),
.A2(n_34),
.B1(n_67),
.B2(n_70),
.Y(n_296)
);

OAI22xp5_ASAP7_75t_L g324 ( 
.A1(n_14),
.A2(n_34),
.B1(n_81),
.B2(n_325),
.Y(n_324)
);

INVx6_ASAP7_75t_L g31 ( 
.A(n_15),
.Y(n_31)
);

INVx3_ASAP7_75t_L g115 ( 
.A(n_15),
.Y(n_115)
);

INVx6_ASAP7_75t_L g175 ( 
.A(n_15),
.Y(n_175)
);

MAJx2_ASAP7_75t_L g16 ( 
.A(n_17),
.B(n_349),
.C(n_354),
.Y(n_16)
);

OAI21xp5_ASAP7_75t_SL g17 ( 
.A1(n_18),
.A2(n_347),
.B(n_352),
.Y(n_17)
);

AOI21xp5_ASAP7_75t_L g18 ( 
.A1(n_19),
.A2(n_334),
.B(n_346),
.Y(n_18)
);

OAI321xp33_ASAP7_75t_L g19 ( 
.A1(n_20),
.A2(n_300),
.A3(n_327),
.B1(n_332),
.B2(n_333),
.C(n_356),
.Y(n_19)
);

AOI21xp5_ASAP7_75t_L g20 ( 
.A1(n_21),
.A2(n_273),
.B(n_299),
.Y(n_20)
);

OAI21xp5_ASAP7_75t_SL g21 ( 
.A1(n_22),
.A2(n_249),
.B(n_272),
.Y(n_21)
);

O2A1O1Ixp33_ASAP7_75t_SL g22 ( 
.A1(n_23),
.A2(n_135),
.B(n_223),
.C(n_248),
.Y(n_22)
);

AND2x2_ASAP7_75t_L g23 ( 
.A(n_24),
.B(n_119),
.Y(n_23)
);

NOR2xp33_ASAP7_75t_L g222 ( 
.A(n_24),
.B(n_119),
.Y(n_222)
);

XNOR2xp5_ASAP7_75t_L g24 ( 
.A(n_25),
.B(n_99),
.Y(n_24)
);

AOI22xp5_ASAP7_75t_L g25 ( 
.A1(n_26),
.A2(n_27),
.B1(n_56),
.B2(n_57),
.Y(n_25)
);

MAJIxp5_ASAP7_75t_L g224 ( 
.A(n_26),
.B(n_57),
.C(n_99),
.Y(n_224)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_27),
.Y(n_26)
);

XNOR2xp5_ASAP7_75t_SL g27 ( 
.A(n_28),
.B(n_41),
.Y(n_27)
);

NAND2xp5_ASAP7_75t_L g228 ( 
.A(n_28),
.B(n_41),
.Y(n_228)
);

OAI21xp5_ASAP7_75t_L g28 ( 
.A1(n_29),
.A2(n_32),
.B(n_35),
.Y(n_28)
);

OAI22xp5_ASAP7_75t_SL g112 ( 
.A1(n_29),
.A2(n_32),
.B1(n_113),
.B2(n_115),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_L g134 ( 
.A(n_29),
.B(n_39),
.Y(n_134)
);

OAI21xp5_ASAP7_75t_L g155 ( 
.A1(n_29),
.A2(n_156),
.B(n_157),
.Y(n_155)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_29),
.Y(n_163)
);

OAI22xp5_ASAP7_75t_SL g182 ( 
.A1(n_29),
.A2(n_165),
.B1(n_172),
.B2(n_178),
.Y(n_182)
);

AOI21xp5_ASAP7_75t_L g255 ( 
.A1(n_29),
.A2(n_37),
.B(n_256),
.Y(n_255)
);

NAND2xp5_ASAP7_75t_L g29 ( 
.A(n_30),
.B(n_31),
.Y(n_29)
);

INVx6_ASAP7_75t_L g33 ( 
.A(n_30),
.Y(n_33)
);

OA22x2_ASAP7_75t_L g42 ( 
.A1(n_30),
.A2(n_33),
.B1(n_43),
.B2(n_44),
.Y(n_42)
);

INVx8_ASAP7_75t_L g38 ( 
.A(n_31),
.Y(n_38)
);

INVx3_ASAP7_75t_SL g133 ( 
.A(n_31),
.Y(n_133)
);

INVx5_ASAP7_75t_L g179 ( 
.A(n_31),
.Y(n_179)
);

NOR2xp33_ASAP7_75t_L g176 ( 
.A(n_33),
.B(n_177),
.Y(n_176)
);

INVxp67_ASAP7_75t_L g35 ( 
.A(n_36),
.Y(n_35)
);

AOI21xp5_ASAP7_75t_L g192 ( 
.A1(n_36),
.A2(n_159),
.B(n_163),
.Y(n_192)
);

NOR2xp33_ASAP7_75t_L g36 ( 
.A(n_37),
.B(n_39),
.Y(n_36)
);

INVx3_ASAP7_75t_L g158 ( 
.A(n_37),
.Y(n_158)
);

INVx5_ASAP7_75t_L g37 ( 
.A(n_38),
.Y(n_37)
);

OAI21xp5_ASAP7_75t_L g41 ( 
.A1(n_42),
.A2(n_46),
.B(n_51),
.Y(n_41)
);

NAND2xp5_ASAP7_75t_L g54 ( 
.A(n_42),
.B(n_55),
.Y(n_54)
);

CKINVDCx20_ASAP7_75t_R g64 ( 
.A(n_42),
.Y(n_64)
);

OAI22xp5_ASAP7_75t_SL g145 ( 
.A1(n_42),
.A2(n_54),
.B1(n_146),
.B2(n_147),
.Y(n_145)
);

OAI22xp5_ASAP7_75t_SL g153 ( 
.A1(n_42),
.A2(n_54),
.B1(n_147),
.B2(n_154),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_SL g181 ( 
.A(n_42),
.B(n_85),
.Y(n_181)
);

OAI22xp5_ASAP7_75t_SL g243 ( 
.A1(n_42),
.A2(n_46),
.B1(n_54),
.B2(n_244),
.Y(n_243)
);

AOI21xp5_ASAP7_75t_L g310 ( 
.A1(n_42),
.A2(n_54),
.B(n_60),
.Y(n_310)
);

OAI22xp33_ASAP7_75t_L g55 ( 
.A1(n_43),
.A2(n_44),
.B1(n_47),
.B2(n_48),
.Y(n_55)
);

INVx13_ASAP7_75t_L g43 ( 
.A(n_44),
.Y(n_43)
);

BUFx24_ASAP7_75t_L g44 ( 
.A(n_45),
.Y(n_44)
);

AOI22xp5_ASAP7_75t_L g72 ( 
.A1(n_47),
.A2(n_48),
.B1(n_73),
.B2(n_74),
.Y(n_72)
);

NAND3xp33_ASAP7_75t_L g191 ( 
.A(n_47),
.B(n_67),
.C(n_74),
.Y(n_191)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_48),
.Y(n_47)
);

NAND2xp5_ASAP7_75t_L g142 ( 
.A(n_48),
.B(n_143),
.Y(n_142)
);

A2O1A1Ixp33_ASAP7_75t_L g189 ( 
.A1(n_48),
.A2(n_73),
.B(n_190),
.C(n_191),
.Y(n_189)
);

BUFx2_ASAP7_75t_L g48 ( 
.A(n_49),
.Y(n_48)
);

AND2x2_ASAP7_75t_L g292 ( 
.A(n_51),
.B(n_213),
.Y(n_292)
);

NAND2xp5_ASAP7_75t_L g51 ( 
.A(n_52),
.B(n_53),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_SL g63 ( 
.A(n_52),
.B(n_64),
.Y(n_63)
);

AOI22xp5_ASAP7_75t_L g196 ( 
.A1(n_53),
.A2(n_64),
.B1(n_197),
.B2(n_198),
.Y(n_196)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_54),
.Y(n_53)
);

OAI21xp5_ASAP7_75t_SL g59 ( 
.A1(n_54),
.A2(n_60),
.B(n_63),
.Y(n_59)
);

OAI21xp5_ASAP7_75t_SL g211 ( 
.A1(n_54),
.A2(n_212),
.B(n_213),
.Y(n_211)
);

OAI21xp5_ASAP7_75t_SL g257 ( 
.A1(n_54),
.A2(n_63),
.B(n_244),
.Y(n_257)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_57),
.Y(n_56)
);

MAJIxp5_ASAP7_75t_L g57 ( 
.A(n_58),
.B(n_65),
.C(n_79),
.Y(n_57)
);

AOI22xp5_ASAP7_75t_L g121 ( 
.A1(n_58),
.A2(n_59),
.B1(n_65),
.B2(n_122),
.Y(n_121)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_59),
.Y(n_58)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_61),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_SL g213 ( 
.A(n_61),
.B(n_64),
.Y(n_213)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_65),
.Y(n_122)
);

AOI22xp5_ASAP7_75t_L g65 ( 
.A1(n_66),
.A2(n_71),
.B1(n_76),
.B2(n_77),
.Y(n_65)
);

CKINVDCx20_ASAP7_75t_R g128 ( 
.A(n_66),
.Y(n_128)
);

INVx5_ASAP7_75t_L g70 ( 
.A(n_67),
.Y(n_70)
);

OAI22xp5_ASAP7_75t_L g75 ( 
.A1(n_67),
.A2(n_70),
.B1(n_73),
.B2(n_74),
.Y(n_75)
);

AOI22xp5_ASAP7_75t_L g89 ( 
.A1(n_67),
.A2(n_70),
.B1(n_90),
.B2(n_91),
.Y(n_89)
);

A2O1A1Ixp33_ASAP7_75t_L g116 ( 
.A1(n_67),
.A2(n_86),
.B(n_90),
.C(n_117),
.Y(n_116)
);

HAxp5_ASAP7_75t_SL g190 ( 
.A(n_67),
.B(n_85),
.CON(n_190),
.SN(n_190)
);

BUFx12f_ASAP7_75t_L g67 ( 
.A(n_68),
.Y(n_67)
);

NAND3xp33_ASAP7_75t_L g117 ( 
.A(n_70),
.B(n_91),
.C(n_94),
.Y(n_117)
);

CKINVDCx20_ASAP7_75t_R g108 ( 
.A(n_71),
.Y(n_108)
);

AOI22xp5_ASAP7_75t_L g199 ( 
.A1(n_71),
.A2(n_76),
.B1(n_127),
.B2(n_190),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_L g268 ( 
.A(n_71),
.B(n_237),
.Y(n_268)
);

AOI22xp5_ASAP7_75t_SL g293 ( 
.A1(n_71),
.A2(n_76),
.B1(n_294),
.B2(n_295),
.Y(n_293)
);

OAI21xp5_ASAP7_75t_SL g339 ( 
.A1(n_71),
.A2(n_76),
.B(n_110),
.Y(n_339)
);

AND2x2_ASAP7_75t_L g71 ( 
.A(n_72),
.B(n_75),
.Y(n_71)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_72),
.Y(n_76)
);

OAI22xp5_ASAP7_75t_L g125 ( 
.A1(n_72),
.A2(n_108),
.B1(n_126),
.B2(n_128),
.Y(n_125)
);

OAI21xp5_ASAP7_75t_L g266 ( 
.A1(n_72),
.A2(n_267),
.B(n_268),
.Y(n_266)
);

INVx5_ASAP7_75t_L g74 ( 
.A(n_73),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_SL g109 ( 
.A(n_76),
.B(n_110),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_SL g236 ( 
.A(n_76),
.B(n_237),
.Y(n_236)
);

CKINVDCx16_ASAP7_75t_R g107 ( 
.A(n_77),
.Y(n_107)
);

XNOR2xp5_ASAP7_75t_SL g120 ( 
.A(n_79),
.B(n_121),
.Y(n_120)
);

AOI22xp5_ASAP7_75t_L g79 ( 
.A1(n_80),
.A2(n_88),
.B1(n_95),
.B2(n_96),
.Y(n_79)
);

OAI21xp33_ASAP7_75t_L g80 ( 
.A1(n_81),
.A2(n_85),
.B(n_86),
.Y(n_80)
);

INVx8_ASAP7_75t_L g81 ( 
.A(n_82),
.Y(n_81)
);

INVx8_ASAP7_75t_L g82 ( 
.A(n_83),
.Y(n_82)
);

INVx6_ASAP7_75t_L g83 ( 
.A(n_84),
.Y(n_83)
);

INVx8_ASAP7_75t_L g87 ( 
.A(n_84),
.Y(n_87)
);

INVx11_ASAP7_75t_L g94 ( 
.A(n_84),
.Y(n_94)
);

INVx8_ASAP7_75t_L g287 ( 
.A(n_84),
.Y(n_287)
);

NAND2xp5_ASAP7_75t_SL g86 ( 
.A(n_85),
.B(n_87),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g177 ( 
.A(n_85),
.B(n_178),
.Y(n_177)
);

OAI22xp33_ASAP7_75t_L g92 ( 
.A1(n_87),
.A2(n_90),
.B1(n_91),
.B2(n_93),
.Y(n_92)
);

INVx11_ASAP7_75t_L g325 ( 
.A(n_87),
.Y(n_325)
);

CKINVDCx20_ASAP7_75t_R g103 ( 
.A(n_88),
.Y(n_103)
);

AOI22xp5_ASAP7_75t_L g231 ( 
.A1(n_88),
.A2(n_95),
.B1(n_105),
.B2(n_232),
.Y(n_231)
);

NAND2xp5_ASAP7_75t_L g306 ( 
.A(n_88),
.B(n_286),
.Y(n_306)
);

AOI22xp5_ASAP7_75t_L g322 ( 
.A1(n_88),
.A2(n_95),
.B1(n_323),
.B2(n_324),
.Y(n_322)
);

AOI21xp5_ASAP7_75t_L g340 ( 
.A1(n_88),
.A2(n_324),
.B(n_341),
.Y(n_340)
);

OAI21xp5_ASAP7_75t_SL g354 ( 
.A1(n_88),
.A2(n_95),
.B(n_265),
.Y(n_354)
);

AND2x2_ASAP7_75t_L g88 ( 
.A(n_89),
.B(n_92),
.Y(n_88)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_89),
.Y(n_95)
);

OAI22xp5_ASAP7_75t_SL g102 ( 
.A1(n_89),
.A2(n_97),
.B1(n_103),
.B2(n_104),
.Y(n_102)
);

OAI21xp5_ASAP7_75t_L g304 ( 
.A1(n_89),
.A2(n_305),
.B(n_306),
.Y(n_304)
);

INVx8_ASAP7_75t_L g90 ( 
.A(n_91),
.Y(n_90)
);

INVx8_ASAP7_75t_L g93 ( 
.A(n_94),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_SL g264 ( 
.A(n_95),
.B(n_265),
.Y(n_264)
);

NAND2xp5_ASAP7_75t_SL g285 ( 
.A(n_95),
.B(n_286),
.Y(n_285)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_97),
.Y(n_96)
);

OAI22xp5_ASAP7_75t_SL g99 ( 
.A1(n_100),
.A2(n_101),
.B1(n_111),
.B2(n_118),
.Y(n_99)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_101),
.Y(n_100)
);

XNOR2xp5_ASAP7_75t_SL g101 ( 
.A(n_102),
.B(n_106),
.Y(n_101)
);

MAJIxp5_ASAP7_75t_L g247 ( 
.A(n_102),
.B(n_106),
.C(n_118),
.Y(n_247)
);

OAI21xp5_ASAP7_75t_SL g262 ( 
.A1(n_103),
.A2(n_263),
.B(n_264),
.Y(n_262)
);

OAI21xp5_ASAP7_75t_SL g283 ( 
.A1(n_103),
.A2(n_284),
.B(n_285),
.Y(n_283)
);

CKINVDCx20_ASAP7_75t_R g104 ( 
.A(n_105),
.Y(n_104)
);

OAI21xp5_ASAP7_75t_L g106 ( 
.A1(n_107),
.A2(n_108),
.B(n_109),
.Y(n_106)
);

OAI21xp33_ASAP7_75t_L g234 ( 
.A1(n_108),
.A2(n_235),
.B(n_236),
.Y(n_234)
);

OAI21xp33_ASAP7_75t_L g309 ( 
.A1(n_108),
.A2(n_236),
.B(n_296),
.Y(n_309)
);

NAND2xp5_ASAP7_75t_L g321 ( 
.A(n_109),
.B(n_268),
.Y(n_321)
);

CKINVDCx20_ASAP7_75t_R g235 ( 
.A(n_110),
.Y(n_235)
);

CKINVDCx14_ASAP7_75t_R g118 ( 
.A(n_111),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_L g111 ( 
.A(n_112),
.B(n_116),
.Y(n_111)
);

XNOR2xp5_ASAP7_75t_L g123 ( 
.A(n_112),
.B(n_116),
.Y(n_123)
);

CKINVDCx20_ASAP7_75t_R g113 ( 
.A(n_114),
.Y(n_113)
);

AOI21xp5_ASAP7_75t_L g132 ( 
.A1(n_114),
.A2(n_133),
.B(n_134),
.Y(n_132)
);

MAJIxp5_ASAP7_75t_L g119 ( 
.A(n_120),
.B(n_123),
.C(n_124),
.Y(n_119)
);

XOR2xp5_ASAP7_75t_L g218 ( 
.A(n_120),
.B(n_219),
.Y(n_218)
);

XOR2xp5_ASAP7_75t_L g219 ( 
.A(n_123),
.B(n_124),
.Y(n_219)
);

MAJIxp5_ASAP7_75t_L g124 ( 
.A(n_125),
.B(n_129),
.C(n_131),
.Y(n_124)
);

XOR2xp5_ASAP7_75t_L g206 ( 
.A(n_125),
.B(n_207),
.Y(n_206)
);

CKINVDCx16_ASAP7_75t_R g126 ( 
.A(n_127),
.Y(n_126)
);

AOI22xp5_ASAP7_75t_L g207 ( 
.A1(n_129),
.A2(n_130),
.B1(n_131),
.B2(n_132),
.Y(n_207)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_130),
.Y(n_129)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_132),
.Y(n_131)
);

AOI22xp5_ASAP7_75t_L g162 ( 
.A1(n_133),
.A2(n_163),
.B1(n_164),
.B2(n_166),
.Y(n_162)
);

NOR2xp33_ASAP7_75t_SL g240 ( 
.A(n_134),
.B(n_241),
.Y(n_240)
);

NOR2xp33_ASAP7_75t_SL g135 ( 
.A(n_136),
.B(n_222),
.Y(n_135)
);

AOI21xp5_ASAP7_75t_SL g136 ( 
.A1(n_137),
.A2(n_217),
.B(n_221),
.Y(n_136)
);

OAI21xp5_ASAP7_75t_SL g137 ( 
.A1(n_138),
.A2(n_202),
.B(n_216),
.Y(n_137)
);

AOI21xp5_ASAP7_75t_SL g138 ( 
.A1(n_139),
.A2(n_186),
.B(n_201),
.Y(n_138)
);

OAI21xp5_ASAP7_75t_SL g139 ( 
.A1(n_140),
.A2(n_160),
.B(n_185),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_L g140 ( 
.A(n_141),
.B(n_148),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_L g185 ( 
.A(n_141),
.B(n_148),
.Y(n_185)
);

NOR2xp33_ASAP7_75t_L g141 ( 
.A(n_142),
.B(n_144),
.Y(n_141)
);

AOI22xp5_ASAP7_75t_L g167 ( 
.A1(n_142),
.A2(n_144),
.B1(n_145),
.B2(n_168),
.Y(n_167)
);

CKINVDCx20_ASAP7_75t_R g168 ( 
.A(n_142),
.Y(n_168)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_145),
.Y(n_144)
);

XNOR2xp5_ASAP7_75t_L g148 ( 
.A(n_149),
.B(n_155),
.Y(n_148)
);

AOI22xp5_ASAP7_75t_L g149 ( 
.A1(n_150),
.A2(n_151),
.B1(n_152),
.B2(n_153),
.Y(n_149)
);

MAJIxp5_ASAP7_75t_L g200 ( 
.A(n_150),
.B(n_153),
.C(n_155),
.Y(n_200)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_151),
.Y(n_150)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_153),
.Y(n_152)
);

INVxp67_ASAP7_75t_L g197 ( 
.A(n_154),
.Y(n_197)
);

CKINVDCx14_ASAP7_75t_R g166 ( 
.A(n_156),
.Y(n_166)
);

INVxp33_ASAP7_75t_L g241 ( 
.A(n_157),
.Y(n_241)
);

NAND2xp5_ASAP7_75t_L g157 ( 
.A(n_158),
.B(n_159),
.Y(n_157)
);

CKINVDCx20_ASAP7_75t_R g256 ( 
.A(n_159),
.Y(n_256)
);

AOI21xp5_ASAP7_75t_L g160 ( 
.A1(n_161),
.A2(n_169),
.B(n_184),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_L g161 ( 
.A(n_162),
.B(n_167),
.Y(n_161)
);

NOR2xp33_ASAP7_75t_L g184 ( 
.A(n_162),
.B(n_167),
.Y(n_184)
);

CKINVDCx16_ASAP7_75t_R g164 ( 
.A(n_165),
.Y(n_164)
);

OAI21xp5_ASAP7_75t_L g169 ( 
.A1(n_170),
.A2(n_180),
.B(n_183),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_SL g170 ( 
.A(n_171),
.B(n_176),
.Y(n_170)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_174),
.Y(n_173)
);

INVx2_ASAP7_75t_L g174 ( 
.A(n_175),
.Y(n_174)
);

INVx2_ASAP7_75t_L g178 ( 
.A(n_179),
.Y(n_178)
);

NOR2xp33_ASAP7_75t_L g180 ( 
.A(n_181),
.B(n_182),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_SL g183 ( 
.A(n_181),
.B(n_182),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_SL g186 ( 
.A(n_187),
.B(n_200),
.Y(n_186)
);

NOR2xp33_ASAP7_75t_L g201 ( 
.A(n_187),
.B(n_200),
.Y(n_201)
);

XOR2xp5_ASAP7_75t_L g187 ( 
.A(n_188),
.B(n_195),
.Y(n_187)
);

MAJIxp5_ASAP7_75t_L g203 ( 
.A(n_188),
.B(n_196),
.C(n_199),
.Y(n_203)
);

AOI22xp5_ASAP7_75t_L g188 ( 
.A1(n_189),
.A2(n_192),
.B1(n_193),
.B2(n_194),
.Y(n_188)
);

CKINVDCx14_ASAP7_75t_R g193 ( 
.A(n_189),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_L g210 ( 
.A(n_189),
.B(n_194),
.Y(n_210)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_192),
.Y(n_194)
);

XOR2xp5_ASAP7_75t_L g195 ( 
.A(n_196),
.B(n_199),
.Y(n_195)
);

CKINVDCx16_ASAP7_75t_R g212 ( 
.A(n_198),
.Y(n_212)
);

NOR2xp33_ASAP7_75t_L g202 ( 
.A(n_203),
.B(n_204),
.Y(n_202)
);

NAND2xp5_ASAP7_75t_SL g216 ( 
.A(n_203),
.B(n_204),
.Y(n_216)
);

OAI22xp5_ASAP7_75t_SL g204 ( 
.A1(n_205),
.A2(n_206),
.B1(n_208),
.B2(n_209),
.Y(n_204)
);

MAJIxp5_ASAP7_75t_L g220 ( 
.A(n_205),
.B(n_211),
.C(n_214),
.Y(n_220)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_206),
.Y(n_205)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_209),
.Y(n_208)
);

OAI22xp5_ASAP7_75t_SL g209 ( 
.A1(n_210),
.A2(n_211),
.B1(n_214),
.B2(n_215),
.Y(n_209)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_210),
.Y(n_214)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_211),
.Y(n_215)
);

NAND2xp5_ASAP7_75t_SL g217 ( 
.A(n_218),
.B(n_220),
.Y(n_217)
);

NOR2xp33_ASAP7_75t_L g221 ( 
.A(n_218),
.B(n_220),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_L g223 ( 
.A(n_224),
.B(n_225),
.Y(n_223)
);

NOR2xp33_ASAP7_75t_L g248 ( 
.A(n_224),
.B(n_225),
.Y(n_248)
);

XOR2xp5_ASAP7_75t_L g225 ( 
.A(n_226),
.B(n_247),
.Y(n_225)
);

OAI22xp5_ASAP7_75t_SL g226 ( 
.A1(n_227),
.A2(n_238),
.B1(n_245),
.B2(n_246),
.Y(n_226)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_227),
.Y(n_245)
);

XOR2xp5_ASAP7_75t_L g227 ( 
.A(n_228),
.B(n_229),
.Y(n_227)
);

MAJIxp5_ASAP7_75t_L g271 ( 
.A(n_228),
.B(n_231),
.C(n_233),
.Y(n_271)
);

AOI22xp5_ASAP7_75t_L g229 ( 
.A1(n_230),
.A2(n_231),
.B1(n_233),
.B2(n_234),
.Y(n_229)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_231),
.Y(n_230)
);

CKINVDCx20_ASAP7_75t_R g263 ( 
.A(n_232),
.Y(n_263)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_234),
.Y(n_233)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_238),
.Y(n_246)
);

MAJIxp5_ASAP7_75t_L g250 ( 
.A(n_238),
.B(n_245),
.C(n_247),
.Y(n_250)
);

AOI22xp5_ASAP7_75t_L g238 ( 
.A1(n_239),
.A2(n_240),
.B1(n_242),
.B2(n_243),
.Y(n_238)
);

NAND2xp5_ASAP7_75t_L g269 ( 
.A(n_239),
.B(n_243),
.Y(n_269)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_240),
.Y(n_239)
);

CKINVDCx14_ASAP7_75t_R g242 ( 
.A(n_243),
.Y(n_242)
);

NOR2xp33_ASAP7_75t_L g249 ( 
.A(n_250),
.B(n_251),
.Y(n_249)
);

NAND2xp5_ASAP7_75t_SL g272 ( 
.A(n_250),
.B(n_251),
.Y(n_272)
);

XNOR2xp5_ASAP7_75t_L g251 ( 
.A(n_252),
.B(n_271),
.Y(n_251)
);

XNOR2xp5_ASAP7_75t_L g252 ( 
.A(n_253),
.B(n_259),
.Y(n_252)
);

MAJIxp5_ASAP7_75t_L g274 ( 
.A(n_253),
.B(n_259),
.C(n_271),
.Y(n_274)
);

OAI22xp5_ASAP7_75t_L g253 ( 
.A1(n_254),
.A2(n_255),
.B1(n_257),
.B2(n_258),
.Y(n_253)
);

AOI22xp5_ASAP7_75t_L g281 ( 
.A1(n_254),
.A2(n_255),
.B1(n_282),
.B2(n_283),
.Y(n_281)
);

OAI21xp5_ASAP7_75t_L g314 ( 
.A1(n_254),
.A2(n_279),
.B(n_283),
.Y(n_314)
);

CKINVDCx14_ASAP7_75t_R g254 ( 
.A(n_255),
.Y(n_254)
);

NAND2xp5_ASAP7_75t_L g280 ( 
.A(n_255),
.B(n_257),
.Y(n_280)
);

CKINVDCx20_ASAP7_75t_R g258 ( 
.A(n_257),
.Y(n_258)
);

OAI22xp5_ASAP7_75t_SL g259 ( 
.A1(n_260),
.A2(n_261),
.B1(n_269),
.B2(n_270),
.Y(n_259)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_261),
.Y(n_260)
);

XNOR2xp5_ASAP7_75t_SL g261 ( 
.A(n_262),
.B(n_266),
.Y(n_261)
);

MAJIxp5_ASAP7_75t_L g298 ( 
.A(n_262),
.B(n_266),
.C(n_270),
.Y(n_298)
);

NAND2xp5_ASAP7_75t_SL g349 ( 
.A(n_264),
.B(n_306),
.Y(n_349)
);

CKINVDCx20_ASAP7_75t_R g284 ( 
.A(n_265),
.Y(n_284)
);

CKINVDCx16_ASAP7_75t_R g294 ( 
.A(n_267),
.Y(n_294)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_269),
.Y(n_270)
);

NAND2xp5_ASAP7_75t_L g273 ( 
.A(n_274),
.B(n_275),
.Y(n_273)
);

NOR2xp33_ASAP7_75t_SL g299 ( 
.A(n_274),
.B(n_275),
.Y(n_299)
);

XOR2xp5_ASAP7_75t_L g275 ( 
.A(n_276),
.B(n_298),
.Y(n_275)
);

OAI22xp5_ASAP7_75t_SL g276 ( 
.A1(n_277),
.A2(n_278),
.B1(n_290),
.B2(n_291),
.Y(n_276)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_278),
.Y(n_277)
);

MAJIxp5_ASAP7_75t_L g328 ( 
.A(n_278),
.B(n_290),
.C(n_298),
.Y(n_328)
);

AOI22xp5_ASAP7_75t_L g278 ( 
.A1(n_279),
.A2(n_280),
.B1(n_281),
.B2(n_289),
.Y(n_278)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_280),
.Y(n_279)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_281),
.Y(n_289)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_283),
.Y(n_282)
);

CKINVDCx20_ASAP7_75t_R g341 ( 
.A(n_285),
.Y(n_341)
);

INVx4_ASAP7_75t_L g288 ( 
.A(n_287),
.Y(n_288)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_291),
.Y(n_290)
);

OAI21xp5_ASAP7_75t_SL g291 ( 
.A1(n_292),
.A2(n_293),
.B(n_297),
.Y(n_291)
);

NAND2xp5_ASAP7_75t_L g297 ( 
.A(n_292),
.B(n_293),
.Y(n_297)
);

CKINVDCx20_ASAP7_75t_R g295 ( 
.A(n_296),
.Y(n_295)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_297),
.Y(n_313)
);

AOI22xp5_ASAP7_75t_L g330 ( 
.A1(n_297),
.A2(n_302),
.B1(n_313),
.B2(n_331),
.Y(n_330)
);

NOR2xp33_ASAP7_75t_L g300 ( 
.A(n_301),
.B(n_315),
.Y(n_300)
);

NAND2xp5_ASAP7_75t_L g333 ( 
.A(n_301),
.B(n_315),
.Y(n_333)
);

MAJIxp5_ASAP7_75t_L g301 ( 
.A(n_302),
.B(n_313),
.C(n_314),
.Y(n_301)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_302),
.Y(n_331)
);

AOI22xp5_ASAP7_75t_L g302 ( 
.A1(n_303),
.A2(n_304),
.B1(n_307),
.B2(n_312),
.Y(n_302)
);

AOI22xp5_ASAP7_75t_L g316 ( 
.A1(n_303),
.A2(n_304),
.B1(n_317),
.B2(n_318),
.Y(n_316)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_304),
.Y(n_303)
);

MAJIxp5_ASAP7_75t_L g326 ( 
.A(n_304),
.B(n_308),
.C(n_311),
.Y(n_326)
);

MAJIxp5_ASAP7_75t_L g335 ( 
.A(n_304),
.B(n_318),
.C(n_326),
.Y(n_335)
);

CKINVDCx20_ASAP7_75t_R g323 ( 
.A(n_305),
.Y(n_323)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_307),
.Y(n_312)
);

AOI22xp5_ASAP7_75t_L g307 ( 
.A1(n_308),
.A2(n_309),
.B1(n_310),
.B2(n_311),
.Y(n_307)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_309),
.Y(n_308)
);

CKINVDCx20_ASAP7_75t_R g311 ( 
.A(n_310),
.Y(n_311)
);

AOI22xp5_ASAP7_75t_L g319 ( 
.A1(n_310),
.A2(n_311),
.B1(n_320),
.B2(n_321),
.Y(n_319)
);

MAJIxp5_ASAP7_75t_L g345 ( 
.A(n_310),
.B(n_320),
.C(n_322),
.Y(n_345)
);

XOR2xp5_ASAP7_75t_L g329 ( 
.A(n_314),
.B(n_330),
.Y(n_329)
);

XNOR2xp5_ASAP7_75t_L g315 ( 
.A(n_316),
.B(n_326),
.Y(n_315)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_318),
.Y(n_317)
);

XOR2xp5_ASAP7_75t_L g318 ( 
.A(n_319),
.B(n_322),
.Y(n_318)
);

CKINVDCx20_ASAP7_75t_R g320 ( 
.A(n_321),
.Y(n_320)
);

NOR2xp33_ASAP7_75t_L g327 ( 
.A(n_328),
.B(n_329),
.Y(n_327)
);

NAND2xp5_ASAP7_75t_SL g332 ( 
.A(n_328),
.B(n_329),
.Y(n_332)
);

NAND2xp5_ASAP7_75t_SL g334 ( 
.A(n_335),
.B(n_336),
.Y(n_334)
);

NOR2xp33_ASAP7_75t_L g346 ( 
.A(n_335),
.B(n_336),
.Y(n_346)
);

AOI22xp5_ASAP7_75t_L g336 ( 
.A1(n_337),
.A2(n_338),
.B1(n_344),
.B2(n_345),
.Y(n_336)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_338),
.Y(n_337)
);

AOI22xp5_ASAP7_75t_L g338 ( 
.A1(n_339),
.A2(n_340),
.B1(n_342),
.B2(n_343),
.Y(n_338)
);

CKINVDCx20_ASAP7_75t_R g342 ( 
.A(n_339),
.Y(n_342)
);

CKINVDCx20_ASAP7_75t_R g343 ( 
.A(n_340),
.Y(n_343)
);

MAJIxp5_ASAP7_75t_L g351 ( 
.A(n_340),
.B(n_342),
.C(n_344),
.Y(n_351)
);

CKINVDCx16_ASAP7_75t_R g344 ( 
.A(n_345),
.Y(n_344)
);

INVxp67_ASAP7_75t_L g347 ( 
.A(n_348),
.Y(n_347)
);

NAND2xp5_ASAP7_75t_L g348 ( 
.A(n_349),
.B(n_350),
.Y(n_348)
);

CKINVDCx20_ASAP7_75t_R g353 ( 
.A(n_349),
.Y(n_353)
);

INVx1_ASAP7_75t_L g350 ( 
.A(n_351),
.Y(n_350)
);

NAND2xp5_ASAP7_75t_SL g352 ( 
.A(n_351),
.B(n_353),
.Y(n_352)
);


endmodule