module fake_jpeg_28102_n_132 (n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_132);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_132;

wire n_117;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_42;
wire n_49;
wire n_16;
wire n_76;
wire n_127;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_31;
wire n_29;
wire n_103;
wire n_50;
wire n_15;
wire n_124;
wire n_13;
wire n_57;
wire n_21;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_30;
wire n_106;
wire n_111;
wire n_44;
wire n_24;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_20;
wire n_18;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_22;
wire n_101;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_97;
wire n_36;
wire n_62;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_96;

INVx13_ASAP7_75t_L g13 ( 
.A(n_7),
.Y(n_13)
);

INVx1_ASAP7_75t_L g14 ( 
.A(n_7),
.Y(n_14)
);

INVx1_ASAP7_75t_L g15 ( 
.A(n_1),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_4),
.Y(n_16)
);

BUFx12f_ASAP7_75t_L g17 ( 
.A(n_11),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_2),
.Y(n_18)
);

NOR2xp33_ASAP7_75t_L g19 ( 
.A(n_11),
.B(n_8),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_4),
.Y(n_20)
);

BUFx3_ASAP7_75t_L g21 ( 
.A(n_2),
.Y(n_21)
);

BUFx12f_ASAP7_75t_L g22 ( 
.A(n_5),
.Y(n_22)
);

INVx1_ASAP7_75t_SL g23 ( 
.A(n_8),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_4),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_10),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_3),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_3),
.Y(n_27)
);

NOR2xp33_ASAP7_75t_L g28 ( 
.A(n_23),
.B(n_0),
.Y(n_28)
);

NOR2xp33_ASAP7_75t_L g38 ( 
.A(n_28),
.B(n_29),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_L g29 ( 
.A(n_23),
.B(n_5),
.Y(n_29)
);

OR2x2_ASAP7_75t_L g30 ( 
.A(n_17),
.B(n_0),
.Y(n_30)
);

NOR2xp33_ASAP7_75t_L g41 ( 
.A(n_30),
.B(n_33),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_17),
.Y(n_31)
);

INVx2_ASAP7_75t_L g43 ( 
.A(n_31),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_17),
.Y(n_32)
);

INVx2_ASAP7_75t_L g45 ( 
.A(n_32),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g33 ( 
.A(n_19),
.B(n_6),
.Y(n_33)
);

BUFx12f_ASAP7_75t_L g34 ( 
.A(n_17),
.Y(n_34)
);

INVx4_ASAP7_75t_L g49 ( 
.A(n_34),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g35 ( 
.A(n_22),
.B(n_6),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_35),
.B(n_36),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g36 ( 
.A(n_22),
.B(n_9),
.Y(n_36)
);

AOI22xp5_ASAP7_75t_L g37 ( 
.A1(n_28),
.A2(n_13),
.B1(n_27),
.B2(n_15),
.Y(n_37)
);

MAJIxp5_ASAP7_75t_L g64 ( 
.A(n_37),
.B(n_26),
.C(n_27),
.Y(n_64)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_34),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_39),
.B(n_42),
.Y(n_55)
);

BUFx2_ASAP7_75t_L g40 ( 
.A(n_31),
.Y(n_40)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_40),
.Y(n_61)
);

CKINVDCx16_ASAP7_75t_R g42 ( 
.A(n_30),
.Y(n_42)
);

INVx11_ASAP7_75t_L g44 ( 
.A(n_34),
.Y(n_44)
);

INVx5_ASAP7_75t_L g58 ( 
.A(n_44),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_L g46 ( 
.A(n_30),
.B(n_22),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_L g52 ( 
.A(n_46),
.B(n_48),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g47 ( 
.A(n_34),
.B(n_14),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_SL g54 ( 
.A(n_47),
.B(n_13),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_L g48 ( 
.A(n_31),
.B(n_22),
.Y(n_48)
);

AOI22xp33_ASAP7_75t_SL g51 ( 
.A1(n_49),
.A2(n_13),
.B1(n_16),
.B2(n_26),
.Y(n_51)
);

INVxp67_ASAP7_75t_L g69 ( 
.A(n_51),
.Y(n_69)
);

INVx2_ASAP7_75t_L g53 ( 
.A(n_43),
.Y(n_53)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_53),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_SL g68 ( 
.A(n_54),
.B(n_63),
.Y(n_68)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_43),
.Y(n_56)
);

INVx2_ASAP7_75t_L g80 ( 
.A(n_56),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_L g57 ( 
.A(n_46),
.B(n_16),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_L g75 ( 
.A(n_57),
.B(n_65),
.Y(n_75)
);

XOR2xp5_ASAP7_75t_L g59 ( 
.A(n_41),
.B(n_15),
.Y(n_59)
);

XOR2xp5_ASAP7_75t_L g76 ( 
.A(n_59),
.B(n_38),
.Y(n_76)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_45),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_60),
.B(n_62),
.Y(n_73)
);

INVx3_ASAP7_75t_L g62 ( 
.A(n_44),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_50),
.B(n_14),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_SL g67 ( 
.A(n_64),
.B(n_41),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_L g65 ( 
.A(n_42),
.B(n_24),
.Y(n_65)
);

OAI21xp5_ASAP7_75t_SL g66 ( 
.A1(n_55),
.A2(n_65),
.B(n_52),
.Y(n_66)
);

AOI21xp5_ASAP7_75t_L g87 ( 
.A1(n_66),
.A2(n_38),
.B(n_50),
.Y(n_87)
);

AND2x2_ASAP7_75t_L g92 ( 
.A(n_67),
.B(n_76),
.Y(n_92)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_53),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_L g86 ( 
.A(n_71),
.B(n_74),
.Y(n_86)
);

CKINVDCx20_ASAP7_75t_R g72 ( 
.A(n_56),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_SL g88 ( 
.A(n_72),
.B(n_77),
.Y(n_88)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_60),
.Y(n_74)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_61),
.Y(n_77)
);

CKINVDCx20_ASAP7_75t_R g78 ( 
.A(n_62),
.Y(n_78)
);

OR2x2_ASAP7_75t_L g84 ( 
.A(n_78),
.B(n_45),
.Y(n_84)
);

O2A1O1Ixp33_ASAP7_75t_L g79 ( 
.A1(n_52),
.A2(n_48),
.B(n_39),
.C(n_49),
.Y(n_79)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_79),
.Y(n_90)
);

OAI22xp5_ASAP7_75t_L g81 ( 
.A1(n_69),
.A2(n_64),
.B1(n_57),
.B2(n_37),
.Y(n_81)
);

OAI22xp5_ASAP7_75t_L g103 ( 
.A1(n_81),
.A2(n_74),
.B1(n_71),
.B2(n_20),
.Y(n_103)
);

INVx2_ASAP7_75t_L g82 ( 
.A(n_70),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_82),
.B(n_84),
.Y(n_93)
);

MAJIxp5_ASAP7_75t_L g83 ( 
.A(n_76),
.B(n_59),
.C(n_32),
.Y(n_83)
);

MAJIxp5_ASAP7_75t_L g94 ( 
.A(n_83),
.B(n_85),
.C(n_91),
.Y(n_94)
);

MAJIxp5_ASAP7_75t_L g85 ( 
.A(n_66),
.B(n_32),
.C(n_61),
.Y(n_85)
);

MAJIxp5_ASAP7_75t_L g101 ( 
.A(n_87),
.B(n_89),
.C(n_20),
.Y(n_101)
);

XNOR2xp5_ASAP7_75t_L g89 ( 
.A(n_75),
.B(n_18),
.Y(n_89)
);

MAJIxp5_ASAP7_75t_L g91 ( 
.A(n_75),
.B(n_25),
.C(n_40),
.Y(n_91)
);

XNOR2x2_ASAP7_75t_L g95 ( 
.A(n_90),
.B(n_79),
.Y(n_95)
);

OAI21xp5_ASAP7_75t_L g105 ( 
.A1(n_95),
.A2(n_96),
.B(n_18),
.Y(n_105)
);

NOR2xp67_ASAP7_75t_SL g96 ( 
.A(n_85),
.B(n_69),
.Y(n_96)
);

A2O1A1Ixp33_ASAP7_75t_SL g97 ( 
.A1(n_88),
.A2(n_73),
.B(n_77),
.C(n_40),
.Y(n_97)
);

INVxp67_ASAP7_75t_L g109 ( 
.A(n_97),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_91),
.B(n_84),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_SL g106 ( 
.A(n_98),
.B(n_99),
.Y(n_106)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_86),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_89),
.B(n_68),
.Y(n_100)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_100),
.Y(n_112)
);

XNOR2xp5_ASAP7_75t_L g107 ( 
.A(n_101),
.B(n_103),
.Y(n_107)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_92),
.Y(n_102)
);

AOI22xp5_ASAP7_75t_SL g110 ( 
.A1(n_102),
.A2(n_24),
.B1(n_70),
.B2(n_58),
.Y(n_110)
);

OAI22xp5_ASAP7_75t_L g104 ( 
.A1(n_95),
.A2(n_83),
.B1(n_92),
.B2(n_80),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_L g116 ( 
.A(n_104),
.B(n_110),
.Y(n_116)
);

OAI21xp5_ASAP7_75t_L g118 ( 
.A1(n_105),
.A2(n_97),
.B(n_9),
.Y(n_118)
);

XOR2xp5_ASAP7_75t_L g108 ( 
.A(n_94),
.B(n_80),
.Y(n_108)
);

MAJIxp5_ASAP7_75t_L g115 ( 
.A(n_108),
.B(n_111),
.C(n_97),
.Y(n_115)
);

MAJIxp5_ASAP7_75t_L g111 ( 
.A(n_94),
.B(n_25),
.C(n_58),
.Y(n_111)
);

XNOR2xp5_ASAP7_75t_L g113 ( 
.A(n_108),
.B(n_111),
.Y(n_113)
);

XOR2xp5_ASAP7_75t_L g121 ( 
.A(n_113),
.B(n_106),
.Y(n_121)
);

AOI21xp5_ASAP7_75t_L g114 ( 
.A1(n_109),
.A2(n_97),
.B(n_93),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_L g123 ( 
.A(n_114),
.B(n_21),
.Y(n_123)
);

MAJIxp5_ASAP7_75t_L g120 ( 
.A(n_115),
.B(n_117),
.C(n_118),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_107),
.B(n_10),
.Y(n_117)
);

INVxp33_ASAP7_75t_L g119 ( 
.A(n_116),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_L g125 ( 
.A(n_119),
.B(n_122),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_L g126 ( 
.A(n_121),
.B(n_0),
.Y(n_126)
);

AOI322xp5_ASAP7_75t_L g122 ( 
.A1(n_115),
.A2(n_109),
.A3(n_112),
.B1(n_25),
.B2(n_12),
.C1(n_21),
.C2(n_3),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_L g127 ( 
.A(n_123),
.B(n_1),
.Y(n_127)
);

OAI21xp5_ASAP7_75t_SL g124 ( 
.A1(n_119),
.A2(n_113),
.B(n_12),
.Y(n_124)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_124),
.Y(n_129)
);

MAJIxp5_ASAP7_75t_L g128 ( 
.A(n_126),
.B(n_127),
.C(n_120),
.Y(n_128)
);

XOR2xp5_ASAP7_75t_L g131 ( 
.A(n_128),
.B(n_2),
.Y(n_131)
);

OAI21xp5_ASAP7_75t_L g130 ( 
.A1(n_129),
.A2(n_125),
.B(n_1),
.Y(n_130)
);

XNOR2xp5_ASAP7_75t_L g132 ( 
.A(n_130),
.B(n_131),
.Y(n_132)
);


endmodule