module fake_netlist_6_2895_n_1085 (n_52, n_16, n_1, n_91, n_119, n_46, n_146, n_163, n_235, n_18, n_21, n_193, n_147, n_154, n_191, n_88, n_3, n_209, n_98, n_113, n_39, n_63, n_223, n_73, n_4, n_148, n_199, n_138, n_22, n_161, n_208, n_68, n_226, n_228, n_252, n_166, n_28, n_184, n_212, n_50, n_158, n_49, n_7, n_210, n_216, n_83, n_206, n_217, n_5, n_101, n_167, n_144, n_174, n_127, n_125, n_153, n_168, n_215, n_178, n_247, n_225, n_77, n_156, n_149, n_152, n_106, n_92, n_145, n_42, n_133, n_96, n_8, n_90, n_160, n_24, n_105, n_131, n_54, n_227, n_132, n_188, n_102, n_186, n_204, n_245, n_0, n_87, n_195, n_189, n_32, n_66, n_85, n_99, n_78, n_84, n_130, n_213, n_164, n_100, n_129, n_13, n_121, n_197, n_11, n_137, n_17, n_23, n_203, n_254, n_142, n_20, n_143, n_207, n_2, n_242, n_180, n_19, n_47, n_62, n_29, n_155, n_219, n_75, n_109, n_150, n_233, n_122, n_45, n_255, n_205, n_34, n_140, n_218, n_70, n_120, n_234, n_251, n_214, n_37, n_15, n_67, n_33, n_82, n_27, n_236, n_246, n_38, n_110, n_151, n_61, n_112, n_172, n_237, n_81, n_59, n_244, n_181, n_76, n_36, n_182, n_26, n_124, n_238, n_239, n_55, n_126, n_202, n_94, n_97, n_108, n_58, n_116, n_211, n_64, n_220, n_117, n_118, n_175, n_224, n_48, n_231, n_65, n_230, n_25, n_40, n_93, n_80, n_141, n_240, n_135, n_196, n_200, n_165, n_139, n_41, n_134, n_177, n_176, n_114, n_86, n_198, n_104, n_222, n_95, n_179, n_243, n_9, n_248, n_107, n_10, n_71, n_74, n_229, n_253, n_6, n_190, n_14, n_123, n_136, n_72, n_187, n_89, n_249, n_173, n_201, n_250, n_103, n_111, n_60, n_159, n_157, n_162, n_170, n_185, n_35, n_183, n_232, n_115, n_12, n_69, n_128, n_241, n_30, n_79, n_43, n_194, n_171, n_31, n_192, n_57, n_169, n_53, n_51, n_44, n_56, n_221, n_1085);

input n_52;
input n_16;
input n_1;
input n_91;
input n_119;
input n_46;
input n_146;
input n_163;
input n_235;
input n_18;
input n_21;
input n_193;
input n_147;
input n_154;
input n_191;
input n_88;
input n_3;
input n_209;
input n_98;
input n_113;
input n_39;
input n_63;
input n_223;
input n_73;
input n_4;
input n_148;
input n_199;
input n_138;
input n_22;
input n_161;
input n_208;
input n_68;
input n_226;
input n_228;
input n_252;
input n_166;
input n_28;
input n_184;
input n_212;
input n_50;
input n_158;
input n_49;
input n_7;
input n_210;
input n_216;
input n_83;
input n_206;
input n_217;
input n_5;
input n_101;
input n_167;
input n_144;
input n_174;
input n_127;
input n_125;
input n_153;
input n_168;
input n_215;
input n_178;
input n_247;
input n_225;
input n_77;
input n_156;
input n_149;
input n_152;
input n_106;
input n_92;
input n_145;
input n_42;
input n_133;
input n_96;
input n_8;
input n_90;
input n_160;
input n_24;
input n_105;
input n_131;
input n_54;
input n_227;
input n_132;
input n_188;
input n_102;
input n_186;
input n_204;
input n_245;
input n_0;
input n_87;
input n_195;
input n_189;
input n_32;
input n_66;
input n_85;
input n_99;
input n_78;
input n_84;
input n_130;
input n_213;
input n_164;
input n_100;
input n_129;
input n_13;
input n_121;
input n_197;
input n_11;
input n_137;
input n_17;
input n_23;
input n_203;
input n_254;
input n_142;
input n_20;
input n_143;
input n_207;
input n_2;
input n_242;
input n_180;
input n_19;
input n_47;
input n_62;
input n_29;
input n_155;
input n_219;
input n_75;
input n_109;
input n_150;
input n_233;
input n_122;
input n_45;
input n_255;
input n_205;
input n_34;
input n_140;
input n_218;
input n_70;
input n_120;
input n_234;
input n_251;
input n_214;
input n_37;
input n_15;
input n_67;
input n_33;
input n_82;
input n_27;
input n_236;
input n_246;
input n_38;
input n_110;
input n_151;
input n_61;
input n_112;
input n_172;
input n_237;
input n_81;
input n_59;
input n_244;
input n_181;
input n_76;
input n_36;
input n_182;
input n_26;
input n_124;
input n_238;
input n_239;
input n_55;
input n_126;
input n_202;
input n_94;
input n_97;
input n_108;
input n_58;
input n_116;
input n_211;
input n_64;
input n_220;
input n_117;
input n_118;
input n_175;
input n_224;
input n_48;
input n_231;
input n_65;
input n_230;
input n_25;
input n_40;
input n_93;
input n_80;
input n_141;
input n_240;
input n_135;
input n_196;
input n_200;
input n_165;
input n_139;
input n_41;
input n_134;
input n_177;
input n_176;
input n_114;
input n_86;
input n_198;
input n_104;
input n_222;
input n_95;
input n_179;
input n_243;
input n_9;
input n_248;
input n_107;
input n_10;
input n_71;
input n_74;
input n_229;
input n_253;
input n_6;
input n_190;
input n_14;
input n_123;
input n_136;
input n_72;
input n_187;
input n_89;
input n_249;
input n_173;
input n_201;
input n_250;
input n_103;
input n_111;
input n_60;
input n_159;
input n_157;
input n_162;
input n_170;
input n_185;
input n_35;
input n_183;
input n_232;
input n_115;
input n_12;
input n_69;
input n_128;
input n_241;
input n_30;
input n_79;
input n_43;
input n_194;
input n_171;
input n_31;
input n_192;
input n_57;
input n_169;
input n_53;
input n_51;
input n_44;
input n_56;
input n_221;

output n_1085;

wire n_992;
wire n_591;
wire n_435;
wire n_793;
wire n_326;
wire n_801;
wire n_256;
wire n_853;
wire n_440;
wire n_587;
wire n_695;
wire n_507;
wire n_968;
wire n_909;
wire n_580;
wire n_762;
wire n_1030;
wire n_881;
wire n_1008;
wire n_465;
wire n_367;
wire n_680;
wire n_760;
wire n_741;
wire n_1027;
wire n_875;
wire n_590;
wire n_625;
wire n_661;
wire n_278;
wire n_1079;
wire n_341;
wire n_362;
wire n_828;
wire n_462;
wire n_1033;
wire n_607;
wire n_671;
wire n_726;
wire n_1052;
wire n_316;
wire n_419;
wire n_304;
wire n_700;
wire n_694;
wire n_933;
wire n_740;
wire n_1038;
wire n_578;
wire n_703;
wire n_1003;
wire n_365;
wire n_978;
wire n_1061;
wire n_384;
wire n_297;
wire n_595;
wire n_627;
wire n_524;
wire n_342;
wire n_820;
wire n_1044;
wire n_951;
wire n_783;
wire n_725;
wire n_952;
wire n_999;
wire n_358;
wire n_751;
wire n_449;
wire n_749;
wire n_798;
wire n_310;
wire n_509;
wire n_368;
wire n_575;
wire n_994;
wire n_1072;
wire n_677;
wire n_969;
wire n_988;
wire n_805;
wire n_396;
wire n_495;
wire n_1065;
wire n_815;
wire n_350;
wire n_585;
wire n_732;
wire n_974;
wire n_568;
wire n_392;
wire n_840;
wire n_442;
wire n_480;
wire n_874;
wire n_724;
wire n_382;
wire n_673;
wire n_1020;
wire n_1009;
wire n_1042;
wire n_1071;
wire n_628;
wire n_1067;
wire n_883;
wire n_557;
wire n_823;
wire n_349;
wire n_643;
wire n_617;
wire n_698;
wire n_898;
wire n_1074;
wire n_1032;
wire n_845;
wire n_807;
wire n_1036;
wire n_739;
wire n_400;
wire n_284;
wire n_337;
wire n_955;
wire n_865;
wire n_893;
wire n_925;
wire n_485;
wire n_1026;
wire n_443;
wire n_892;
wire n_768;
wire n_471;
wire n_289;
wire n_935;
wire n_421;
wire n_781;
wire n_424;
wire n_789;
wire n_615;
wire n_573;
wire n_769;
wire n_320;
wire n_639;
wire n_676;
wire n_327;
wire n_794;
wire n_963;
wire n_727;
wire n_894;
wire n_369;
wire n_597;
wire n_685;
wire n_280;
wire n_287;
wire n_832;
wire n_353;
wire n_610;
wire n_555;
wire n_389;
wire n_814;
wire n_415;
wire n_830;
wire n_605;
wire n_461;
wire n_873;
wire n_383;
wire n_826;
wire n_1024;
wire n_669;
wire n_447;
wire n_872;
wire n_300;
wire n_718;
wire n_517;
wire n_1018;
wire n_747;
wire n_852;
wire n_667;
wire n_542;
wire n_847;
wire n_644;
wire n_682;
wire n_851;
wire n_621;
wire n_305;
wire n_1037;
wire n_721;
wire n_996;
wire n_750;
wire n_532;
wire n_742;
wire n_535;
wire n_691;
wire n_372;
wire n_468;
wire n_544;
wire n_901;
wire n_504;
wire n_923;
wire n_314;
wire n_378;
wire n_413;
wire n_377;
wire n_791;
wire n_510;
wire n_837;
wire n_836;
wire n_1015;
wire n_863;
wire n_375;
wire n_601;
wire n_338;
wire n_522;
wire n_948;
wire n_466;
wire n_704;
wire n_918;
wire n_748;
wire n_506;
wire n_763;
wire n_1057;
wire n_360;
wire n_977;
wire n_945;
wire n_603;
wire n_1005;
wire n_991;
wire n_957;
wire n_536;
wire n_895;
wire n_866;
wire n_622;
wire n_340;
wire n_710;
wire n_387;
wire n_452;
wire n_616;
wire n_658;
wire n_744;
wire n_971;
wire n_946;
wire n_344;
wire n_581;
wire n_428;
wire n_761;
wire n_785;
wire n_746;
wire n_609;
wire n_765;
wire n_432;
wire n_987;
wire n_641;
wire n_822;
wire n_693;
wire n_1056;
wire n_631;
wire n_516;
wire n_720;
wire n_758;
wire n_525;
wire n_842;
wire n_611;
wire n_943;
wire n_491;
wire n_878;
wire n_656;
wire n_772;
wire n_843;
wire n_989;
wire n_797;
wire n_666;
wire n_1016;
wire n_371;
wire n_795;
wire n_770;
wire n_940;
wire n_567;
wire n_899;
wire n_738;
wire n_405;
wire n_538;
wire n_1035;
wire n_294;
wire n_302;
wire n_499;
wire n_380;
wire n_838;
wire n_705;
wire n_647;
wire n_343;
wire n_886;
wire n_448;
wire n_844;
wire n_953;
wire n_1004;
wire n_1017;
wire n_494;
wire n_539;
wire n_493;
wire n_397;
wire n_1022;
wire n_1083;
wire n_614;
wire n_529;
wire n_445;
wire n_425;
wire n_684;
wire n_930;
wire n_888;
wire n_454;
wire n_638;
wire n_910;
wire n_486;
wire n_911;
wire n_381;
wire n_947;
wire n_653;
wire n_887;
wire n_752;
wire n_908;
wire n_944;
wire n_713;
wire n_648;
wire n_657;
wire n_1049;
wire n_576;
wire n_1028;
wire n_472;
wire n_270;
wire n_414;
wire n_563;
wire n_782;
wire n_976;
wire n_490;
wire n_803;
wire n_290;
wire n_809;
wire n_1043;
wire n_1011;
wire n_926;
wire n_927;
wire n_839;
wire n_986;
wire n_734;
wire n_708;
wire n_919;
wire n_1081;
wire n_402;
wire n_352;
wire n_917;
wire n_668;
wire n_478;
wire n_626;
wire n_990;
wire n_574;
wire n_779;
wire n_800;
wire n_929;
wire n_460;
wire n_1084;
wire n_907;
wire n_854;
wire n_1058;
wire n_417;
wire n_446;
wire n_498;
wire n_662;
wire n_374;
wire n_659;
wire n_709;
wire n_904;
wire n_366;
wire n_870;
wire n_777;
wire n_407;
wire n_913;
wire n_450;
wire n_808;
wire n_867;
wire n_272;
wire n_526;
wire n_921;
wire n_712;
wire n_348;
wire n_711;
wire n_579;
wire n_376;
wire n_937;
wire n_390;
wire n_473;
wire n_293;
wire n_1054;
wire n_334;
wire n_559;
wire n_370;
wire n_458;
wire n_1070;
wire n_650;
wire n_998;
wire n_1046;
wire n_717;
wire n_330;
wire n_771;
wire n_470;
wire n_475;
wire n_924;
wire n_298;
wire n_492;
wire n_972;
wire n_281;
wire n_258;
wire n_551;
wire n_699;
wire n_456;
wire n_564;
wire n_260;
wire n_265;
wire n_313;
wire n_451;
wire n_624;
wire n_824;
wire n_962;
wire n_1073;
wire n_1000;
wire n_279;
wire n_686;
wire n_796;
wire n_1041;
wire n_757;
wire n_594;
wire n_565;
wire n_719;
wire n_356;
wire n_577;
wire n_936;
wire n_552;
wire n_1062;
wire n_619;
wire n_885;
wire n_455;
wire n_896;
wire n_521;
wire n_363;
wire n_572;
wire n_912;
wire n_395;
wire n_813;
wire n_592;
wire n_745;
wire n_654;
wire n_323;
wire n_829;
wire n_606;
wire n_393;
wire n_818;
wire n_984;
wire n_411;
wire n_503;
wire n_716;
wire n_623;
wire n_1048;
wire n_884;
wire n_599;
wire n_513;
wire n_855;
wire n_776;
wire n_321;
wire n_645;
wire n_331;
wire n_916;
wire n_1078;
wire n_868;
wire n_570;
wire n_731;
wire n_859;
wire n_406;
wire n_483;
wire n_735;
wire n_934;
wire n_482;
wire n_755;
wire n_931;
wire n_1021;
wire n_474;
wire n_527;
wire n_261;
wire n_608;
wire n_683;
wire n_420;
wire n_620;
wire n_630;
wire n_394;
wire n_312;
wire n_519;
wire n_541;
wire n_512;
wire n_958;
wire n_292;
wire n_307;
wire n_469;
wire n_433;
wire n_500;
wire n_942;
wire n_792;
wire n_880;
wire n_476;
wire n_981;
wire n_714;
wire n_291;
wire n_543;
wire n_889;
wire n_357;
wire n_264;
wire n_263;
wire n_985;
wire n_589;
wire n_860;
wire n_481;
wire n_788;
wire n_819;
wire n_939;
wire n_997;
wire n_821;
wire n_325;
wire n_938;
wire n_1068;
wire n_767;
wire n_804;
wire n_329;
wire n_464;
wire n_600;
wire n_831;
wire n_802;
wire n_982;
wire n_964;
wire n_561;
wire n_477;
wire n_549;
wire n_980;
wire n_533;
wire n_954;
wire n_1075;
wire n_408;
wire n_932;
wire n_806;
wire n_864;
wire n_959;
wire n_879;
wire n_584;
wire n_399;
wire n_979;
wire n_548;
wire n_905;
wire n_282;
wire n_436;
wire n_833;
wire n_523;
wire n_707;
wire n_322;
wire n_993;
wire n_345;
wire n_409;
wire n_354;
wire n_689;
wire n_799;
wire n_505;
wire n_756;
wire n_319;
wire n_547;
wire n_537;
wire n_273;
wire n_558;
wire n_810;
wire n_635;
wire n_787;
wire n_311;
wire n_1064;
wire n_403;
wire n_1080;
wire n_723;
wire n_634;
wire n_1051;
wire n_583;
wire n_596;
wire n_966;
wire n_546;
wire n_562;
wire n_386;
wire n_764;
wire n_1039;
wire n_556;
wire n_1034;
wire n_1066;
wire n_692;
wire n_733;
wire n_754;
wire n_941;
wire n_975;
wire n_1031;
wire n_487;
wire n_550;
wire n_275;
wire n_553;
wire n_652;
wire n_849;
wire n_970;
wire n_560;
wire n_1014;
wire n_753;
wire n_642;
wire n_995;
wire n_276;
wire n_569;
wire n_441;
wire n_811;
wire n_882;
wire n_1060;
wire n_444;
wire n_586;
wire n_423;
wire n_737;
wire n_318;
wire n_303;
wire n_511;
wire n_715;
wire n_467;
wire n_306;
wire n_269;
wire n_359;
wire n_973;
wire n_346;
wire n_416;
wire n_1053;
wire n_530;
wire n_277;
wire n_520;
wire n_1029;
wire n_418;
wire n_618;
wire n_1055;
wire n_790;
wire n_582;
wire n_266;
wire n_296;
wire n_861;
wire n_674;
wire n_857;
wire n_871;
wire n_967;
wire n_775;
wire n_922;
wire n_571;
wire n_268;
wire n_271;
wire n_404;
wire n_651;
wire n_439;
wire n_518;
wire n_299;
wire n_679;
wire n_1069;
wire n_453;
wire n_612;
wire n_633;
wire n_665;
wire n_902;
wire n_333;
wire n_588;
wire n_308;
wire n_309;
wire n_914;
wire n_759;
wire n_1047;
wire n_1010;
wire n_355;
wire n_426;
wire n_317;
wire n_1040;
wire n_915;
wire n_632;
wire n_702;
wire n_431;
wire n_347;
wire n_812;
wire n_459;
wire n_502;
wire n_328;
wire n_672;
wire n_534;
wire n_488;
wire n_429;
wire n_1006;
wire n_373;
wire n_1012;
wire n_497;
wire n_285;
wire n_780;
wire n_773;
wire n_675;
wire n_920;
wire n_257;
wire n_903;
wire n_730;
wire n_655;
wire n_706;
wire n_1045;
wire n_786;
wire n_670;
wire n_286;
wire n_834;
wire n_835;
wire n_928;
wire n_690;
wire n_850;
wire n_401;
wire n_324;
wire n_766;
wire n_743;
wire n_816;
wire n_335;
wire n_430;
wire n_1002;
wire n_463;
wire n_545;
wire n_489;
wire n_877;
wire n_604;
wire n_848;
wire n_1019;
wire n_301;
wire n_274;
wire n_636;
wire n_825;
wire n_728;
wire n_681;
wire n_1063;
wire n_729;
wire n_876;
wire n_774;
wire n_412;
wire n_640;
wire n_660;
wire n_965;
wire n_267;
wire n_438;
wire n_339;
wire n_784;
wire n_315;
wire n_434;
wire n_515;
wire n_983;
wire n_288;
wire n_427;
wire n_1059;
wire n_479;
wire n_496;
wire n_598;
wire n_422;
wire n_696;
wire n_906;
wire n_688;
wire n_722;
wire n_1077;
wire n_961;
wire n_862;
wire n_869;
wire n_351;
wire n_437;
wire n_1082;
wire n_259;
wire n_540;
wire n_593;
wire n_514;
wire n_646;
wire n_528;
wire n_391;
wire n_457;
wire n_697;
wire n_687;
wire n_364;
wire n_890;
wire n_637;
wire n_385;
wire n_295;
wire n_701;
wire n_817;
wire n_950;
wire n_629;
wire n_388;
wire n_858;
wire n_262;
wire n_484;
wire n_613;
wire n_736;
wire n_900;
wire n_897;
wire n_846;
wire n_501;
wire n_841;
wire n_956;
wire n_960;
wire n_531;
wire n_827;
wire n_1001;
wire n_361;
wire n_508;
wire n_663;
wire n_856;
wire n_1050;
wire n_379;
wire n_778;
wire n_1025;
wire n_332;
wire n_891;
wire n_336;
wire n_398;
wire n_410;
wire n_566;
wire n_554;
wire n_602;
wire n_1013;
wire n_1023;
wire n_1076;
wire n_664;
wire n_949;
wire n_678;
wire n_1007;
wire n_649;
wire n_283;

INVx2_ASAP7_75t_SL g256 ( 
.A(n_146),
.Y(n_256)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_172),
.Y(n_257)
);

INVx1_ASAP7_75t_SL g258 ( 
.A(n_42),
.Y(n_258)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_226),
.Y(n_259)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_123),
.Y(n_260)
);

CKINVDCx5p33_ASAP7_75t_R g261 ( 
.A(n_248),
.Y(n_261)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_64),
.Y(n_262)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_1),
.Y(n_263)
);

BUFx2_ASAP7_75t_L g264 ( 
.A(n_133),
.Y(n_264)
);

CKINVDCx5p33_ASAP7_75t_R g265 ( 
.A(n_244),
.Y(n_265)
);

INVx1_ASAP7_75t_SL g266 ( 
.A(n_8),
.Y(n_266)
);

BUFx6f_ASAP7_75t_L g267 ( 
.A(n_26),
.Y(n_267)
);

CKINVDCx5p33_ASAP7_75t_R g268 ( 
.A(n_161),
.Y(n_268)
);

CKINVDCx5p33_ASAP7_75t_R g269 ( 
.A(n_196),
.Y(n_269)
);

HB1xp67_ASAP7_75t_L g270 ( 
.A(n_57),
.Y(n_270)
);

BUFx10_ASAP7_75t_L g271 ( 
.A(n_190),
.Y(n_271)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_135),
.Y(n_272)
);

CKINVDCx5p33_ASAP7_75t_R g273 ( 
.A(n_191),
.Y(n_273)
);

INVx1_ASAP7_75t_SL g274 ( 
.A(n_90),
.Y(n_274)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_101),
.Y(n_275)
);

BUFx2_ASAP7_75t_L g276 ( 
.A(n_50),
.Y(n_276)
);

CKINVDCx5p33_ASAP7_75t_R g277 ( 
.A(n_81),
.Y(n_277)
);

CKINVDCx5p33_ASAP7_75t_R g278 ( 
.A(n_224),
.Y(n_278)
);

CKINVDCx5p33_ASAP7_75t_R g279 ( 
.A(n_200),
.Y(n_279)
);

INVx2_ASAP7_75t_SL g280 ( 
.A(n_119),
.Y(n_280)
);

INVx2_ASAP7_75t_L g281 ( 
.A(n_70),
.Y(n_281)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_75),
.Y(n_282)
);

CKINVDCx5p33_ASAP7_75t_R g283 ( 
.A(n_227),
.Y(n_283)
);

CKINVDCx5p33_ASAP7_75t_R g284 ( 
.A(n_96),
.Y(n_284)
);

CKINVDCx5p33_ASAP7_75t_R g285 ( 
.A(n_18),
.Y(n_285)
);

CKINVDCx5p33_ASAP7_75t_R g286 ( 
.A(n_2),
.Y(n_286)
);

CKINVDCx5p33_ASAP7_75t_R g287 ( 
.A(n_234),
.Y(n_287)
);

CKINVDCx5p33_ASAP7_75t_R g288 ( 
.A(n_116),
.Y(n_288)
);

CKINVDCx5p33_ASAP7_75t_R g289 ( 
.A(n_66),
.Y(n_289)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_103),
.Y(n_290)
);

CKINVDCx5p33_ASAP7_75t_R g291 ( 
.A(n_85),
.Y(n_291)
);

INVx1_ASAP7_75t_SL g292 ( 
.A(n_149),
.Y(n_292)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_218),
.Y(n_293)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_197),
.Y(n_294)
);

CKINVDCx5p33_ASAP7_75t_R g295 ( 
.A(n_245),
.Y(n_295)
);

CKINVDCx20_ASAP7_75t_R g296 ( 
.A(n_98),
.Y(n_296)
);

CKINVDCx5p33_ASAP7_75t_R g297 ( 
.A(n_61),
.Y(n_297)
);

CKINVDCx5p33_ASAP7_75t_R g298 ( 
.A(n_233),
.Y(n_298)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_237),
.Y(n_299)
);

CKINVDCx5p33_ASAP7_75t_R g300 ( 
.A(n_79),
.Y(n_300)
);

CKINVDCx5p33_ASAP7_75t_R g301 ( 
.A(n_0),
.Y(n_301)
);

CKINVDCx5p33_ASAP7_75t_R g302 ( 
.A(n_104),
.Y(n_302)
);

CKINVDCx5p33_ASAP7_75t_R g303 ( 
.A(n_142),
.Y(n_303)
);

CKINVDCx5p33_ASAP7_75t_R g304 ( 
.A(n_219),
.Y(n_304)
);

CKINVDCx20_ASAP7_75t_R g305 ( 
.A(n_207),
.Y(n_305)
);

CKINVDCx5p33_ASAP7_75t_R g306 ( 
.A(n_131),
.Y(n_306)
);

INVx1_ASAP7_75t_SL g307 ( 
.A(n_254),
.Y(n_307)
);

CKINVDCx5p33_ASAP7_75t_R g308 ( 
.A(n_186),
.Y(n_308)
);

CKINVDCx5p33_ASAP7_75t_R g309 ( 
.A(n_19),
.Y(n_309)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_82),
.Y(n_310)
);

CKINVDCx20_ASAP7_75t_R g311 ( 
.A(n_225),
.Y(n_311)
);

CKINVDCx5p33_ASAP7_75t_R g312 ( 
.A(n_137),
.Y(n_312)
);

CKINVDCx5p33_ASAP7_75t_R g313 ( 
.A(n_220),
.Y(n_313)
);

CKINVDCx20_ASAP7_75t_R g314 ( 
.A(n_21),
.Y(n_314)
);

CKINVDCx5p33_ASAP7_75t_R g315 ( 
.A(n_148),
.Y(n_315)
);

CKINVDCx5p33_ASAP7_75t_R g316 ( 
.A(n_145),
.Y(n_316)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_121),
.Y(n_317)
);

BUFx2_ASAP7_75t_L g318 ( 
.A(n_213),
.Y(n_318)
);

CKINVDCx5p33_ASAP7_75t_R g319 ( 
.A(n_223),
.Y(n_319)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_267),
.Y(n_320)
);

INVxp67_ASAP7_75t_SL g321 ( 
.A(n_270),
.Y(n_321)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_267),
.Y(n_322)
);

CKINVDCx5p33_ASAP7_75t_R g323 ( 
.A(n_285),
.Y(n_323)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_267),
.Y(n_324)
);

CKINVDCx5p33_ASAP7_75t_R g325 ( 
.A(n_286),
.Y(n_325)
);

CKINVDCx5p33_ASAP7_75t_R g326 ( 
.A(n_301),
.Y(n_326)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_267),
.Y(n_327)
);

CKINVDCx5p33_ASAP7_75t_R g328 ( 
.A(n_309),
.Y(n_328)
);

CKINVDCx5p33_ASAP7_75t_R g329 ( 
.A(n_288),
.Y(n_329)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_263),
.Y(n_330)
);

NOR2xp33_ASAP7_75t_L g331 ( 
.A(n_264),
.B(n_0),
.Y(n_331)
);

CKINVDCx20_ASAP7_75t_R g332 ( 
.A(n_314),
.Y(n_332)
);

BUFx2_ASAP7_75t_L g333 ( 
.A(n_314),
.Y(n_333)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_257),
.Y(n_334)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_259),
.Y(n_335)
);

CKINVDCx5p33_ASAP7_75t_R g336 ( 
.A(n_261),
.Y(n_336)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_260),
.Y(n_337)
);

INVx1_ASAP7_75t_L g338 ( 
.A(n_262),
.Y(n_338)
);

CKINVDCx5p33_ASAP7_75t_R g339 ( 
.A(n_265),
.Y(n_339)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_272),
.Y(n_340)
);

CKINVDCx20_ASAP7_75t_R g341 ( 
.A(n_296),
.Y(n_341)
);

INVx1_ASAP7_75t_L g342 ( 
.A(n_275),
.Y(n_342)
);

INVx1_ASAP7_75t_L g343 ( 
.A(n_282),
.Y(n_343)
);

INVx1_ASAP7_75t_SL g344 ( 
.A(n_266),
.Y(n_344)
);

AND2x2_ASAP7_75t_L g345 ( 
.A(n_276),
.B(n_318),
.Y(n_345)
);

CKINVDCx5p33_ASAP7_75t_R g346 ( 
.A(n_268),
.Y(n_346)
);

CKINVDCx5p33_ASAP7_75t_R g347 ( 
.A(n_269),
.Y(n_347)
);

CKINVDCx5p33_ASAP7_75t_R g348 ( 
.A(n_288),
.Y(n_348)
);

INVx1_ASAP7_75t_L g349 ( 
.A(n_290),
.Y(n_349)
);

CKINVDCx5p33_ASAP7_75t_R g350 ( 
.A(n_296),
.Y(n_350)
);

CKINVDCx16_ASAP7_75t_R g351 ( 
.A(n_305),
.Y(n_351)
);

CKINVDCx20_ASAP7_75t_R g352 ( 
.A(n_305),
.Y(n_352)
);

INVx1_ASAP7_75t_L g353 ( 
.A(n_293),
.Y(n_353)
);

INVx1_ASAP7_75t_L g354 ( 
.A(n_294),
.Y(n_354)
);

NOR2xp67_ASAP7_75t_L g355 ( 
.A(n_256),
.B(n_1),
.Y(n_355)
);

INVx2_ASAP7_75t_L g356 ( 
.A(n_281),
.Y(n_356)
);

INVxp67_ASAP7_75t_SL g357 ( 
.A(n_299),
.Y(n_357)
);

CKINVDCx5p33_ASAP7_75t_R g358 ( 
.A(n_273),
.Y(n_358)
);

NAND2xp5_ASAP7_75t_L g359 ( 
.A(n_256),
.B(n_2),
.Y(n_359)
);

CKINVDCx20_ASAP7_75t_R g360 ( 
.A(n_311),
.Y(n_360)
);

INVx1_ASAP7_75t_L g361 ( 
.A(n_310),
.Y(n_361)
);

INVx1_ASAP7_75t_L g362 ( 
.A(n_317),
.Y(n_362)
);

CKINVDCx5p33_ASAP7_75t_R g363 ( 
.A(n_336),
.Y(n_363)
);

CKINVDCx5p33_ASAP7_75t_R g364 ( 
.A(n_339),
.Y(n_364)
);

INVx2_ASAP7_75t_L g365 ( 
.A(n_320),
.Y(n_365)
);

NOR2xp33_ASAP7_75t_L g366 ( 
.A(n_329),
.B(n_280),
.Y(n_366)
);

HB1xp67_ASAP7_75t_L g367 ( 
.A(n_344),
.Y(n_367)
);

CKINVDCx5p33_ASAP7_75t_R g368 ( 
.A(n_346),
.Y(n_368)
);

INVx1_ASAP7_75t_L g369 ( 
.A(n_322),
.Y(n_369)
);

INVx1_ASAP7_75t_L g370 ( 
.A(n_324),
.Y(n_370)
);

INVx2_ASAP7_75t_L g371 ( 
.A(n_327),
.Y(n_371)
);

AND2x2_ASAP7_75t_L g372 ( 
.A(n_345),
.B(n_321),
.Y(n_372)
);

INVx1_ASAP7_75t_L g373 ( 
.A(n_356),
.Y(n_373)
);

BUFx6f_ASAP7_75t_L g374 ( 
.A(n_356),
.Y(n_374)
);

NAND2xp5_ASAP7_75t_L g375 ( 
.A(n_347),
.B(n_280),
.Y(n_375)
);

INVx1_ASAP7_75t_SL g376 ( 
.A(n_350),
.Y(n_376)
);

CKINVDCx5p33_ASAP7_75t_R g377 ( 
.A(n_358),
.Y(n_377)
);

INVx1_ASAP7_75t_L g378 ( 
.A(n_334),
.Y(n_378)
);

NAND2xp5_ASAP7_75t_SL g379 ( 
.A(n_323),
.B(n_325),
.Y(n_379)
);

BUFx3_ASAP7_75t_L g380 ( 
.A(n_335),
.Y(n_380)
);

CKINVDCx5p33_ASAP7_75t_R g381 ( 
.A(n_329),
.Y(n_381)
);

CKINVDCx5p33_ASAP7_75t_R g382 ( 
.A(n_348),
.Y(n_382)
);

CKINVDCx20_ASAP7_75t_R g383 ( 
.A(n_341),
.Y(n_383)
);

CKINVDCx5p33_ASAP7_75t_R g384 ( 
.A(n_348),
.Y(n_384)
);

NAND2xp5_ASAP7_75t_L g385 ( 
.A(n_357),
.B(n_281),
.Y(n_385)
);

NAND2xp5_ASAP7_75t_L g386 ( 
.A(n_337),
.B(n_277),
.Y(n_386)
);

INVx1_ASAP7_75t_L g387 ( 
.A(n_338),
.Y(n_387)
);

CKINVDCx5p33_ASAP7_75t_R g388 ( 
.A(n_351),
.Y(n_388)
);

INVx2_ASAP7_75t_L g389 ( 
.A(n_340),
.Y(n_389)
);

INVx3_ASAP7_75t_L g390 ( 
.A(n_342),
.Y(n_390)
);

INVx1_ASAP7_75t_L g391 ( 
.A(n_343),
.Y(n_391)
);

INVx2_ASAP7_75t_L g392 ( 
.A(n_349),
.Y(n_392)
);

NOR2xp33_ASAP7_75t_R g393 ( 
.A(n_323),
.B(n_311),
.Y(n_393)
);

INVx1_ASAP7_75t_L g394 ( 
.A(n_353),
.Y(n_394)
);

INVx1_ASAP7_75t_L g395 ( 
.A(n_354),
.Y(n_395)
);

INVx3_ASAP7_75t_L g396 ( 
.A(n_361),
.Y(n_396)
);

INVx2_ASAP7_75t_L g397 ( 
.A(n_362),
.Y(n_397)
);

BUFx6f_ASAP7_75t_L g398 ( 
.A(n_330),
.Y(n_398)
);

CKINVDCx5p33_ASAP7_75t_R g399 ( 
.A(n_350),
.Y(n_399)
);

INVx2_ASAP7_75t_L g400 ( 
.A(n_359),
.Y(n_400)
);

NAND2xp5_ASAP7_75t_L g401 ( 
.A(n_325),
.B(n_278),
.Y(n_401)
);

INVx1_ASAP7_75t_L g402 ( 
.A(n_355),
.Y(n_402)
);

INVx5_ASAP7_75t_L g403 ( 
.A(n_331),
.Y(n_403)
);

NAND2xp5_ASAP7_75t_L g404 ( 
.A(n_326),
.B(n_319),
.Y(n_404)
);

CKINVDCx20_ASAP7_75t_R g405 ( 
.A(n_341),
.Y(n_405)
);

CKINVDCx5p33_ASAP7_75t_R g406 ( 
.A(n_326),
.Y(n_406)
);

INVx1_ASAP7_75t_SL g407 ( 
.A(n_360),
.Y(n_407)
);

BUFx10_ASAP7_75t_L g408 ( 
.A(n_328),
.Y(n_408)
);

HB1xp67_ASAP7_75t_L g409 ( 
.A(n_328),
.Y(n_409)
);

INVx1_ASAP7_75t_L g410 ( 
.A(n_333),
.Y(n_410)
);

BUFx6f_ASAP7_75t_L g411 ( 
.A(n_352),
.Y(n_411)
);

INVx1_ASAP7_75t_L g412 ( 
.A(n_378),
.Y(n_412)
);

INVx1_ASAP7_75t_L g413 ( 
.A(n_387),
.Y(n_413)
);

NAND2xp5_ASAP7_75t_SL g414 ( 
.A(n_403),
.B(n_279),
.Y(n_414)
);

NAND2xp5_ASAP7_75t_L g415 ( 
.A(n_400),
.B(n_258),
.Y(n_415)
);

INVx1_ASAP7_75t_L g416 ( 
.A(n_391),
.Y(n_416)
);

INVx2_ASAP7_75t_L g417 ( 
.A(n_374),
.Y(n_417)
);

INVx4_ASAP7_75t_L g418 ( 
.A(n_374),
.Y(n_418)
);

NOR2xp33_ASAP7_75t_L g419 ( 
.A(n_386),
.B(n_366),
.Y(n_419)
);

NAND2xp5_ASAP7_75t_L g420 ( 
.A(n_400),
.B(n_274),
.Y(n_420)
);

NAND2xp33_ASAP7_75t_L g421 ( 
.A(n_385),
.B(n_292),
.Y(n_421)
);

NAND2xp5_ASAP7_75t_L g422 ( 
.A(n_375),
.B(n_307),
.Y(n_422)
);

INVx2_ASAP7_75t_SL g423 ( 
.A(n_367),
.Y(n_423)
);

AND2x2_ASAP7_75t_L g424 ( 
.A(n_372),
.B(n_352),
.Y(n_424)
);

AOI22xp33_ASAP7_75t_L g425 ( 
.A1(n_403),
.A2(n_271),
.B1(n_284),
.B2(n_283),
.Y(n_425)
);

INVx2_ASAP7_75t_L g426 ( 
.A(n_374),
.Y(n_426)
);

AND2x6_ASAP7_75t_L g427 ( 
.A(n_402),
.B(n_271),
.Y(n_427)
);

CKINVDCx5p33_ASAP7_75t_R g428 ( 
.A(n_393),
.Y(n_428)
);

NAND2xp5_ASAP7_75t_SL g429 ( 
.A(n_403),
.B(n_401),
.Y(n_429)
);

AOI22xp33_ASAP7_75t_L g430 ( 
.A1(n_403),
.A2(n_271),
.B1(n_289),
.B2(n_287),
.Y(n_430)
);

AOI22xp5_ASAP7_75t_L g431 ( 
.A1(n_379),
.A2(n_295),
.B1(n_297),
.B2(n_291),
.Y(n_431)
);

BUFx6f_ASAP7_75t_L g432 ( 
.A(n_374),
.Y(n_432)
);

INVx2_ASAP7_75t_L g433 ( 
.A(n_365),
.Y(n_433)
);

BUFx4f_ASAP7_75t_L g434 ( 
.A(n_398),
.Y(n_434)
);

NAND2xp5_ASAP7_75t_L g435 ( 
.A(n_403),
.B(n_298),
.Y(n_435)
);

BUFx3_ASAP7_75t_L g436 ( 
.A(n_380),
.Y(n_436)
);

NOR2xp33_ASAP7_75t_SL g437 ( 
.A(n_363),
.B(n_360),
.Y(n_437)
);

INVx2_ASAP7_75t_L g438 ( 
.A(n_365),
.Y(n_438)
);

INVx2_ASAP7_75t_L g439 ( 
.A(n_371),
.Y(n_439)
);

NAND2xp5_ASAP7_75t_SL g440 ( 
.A(n_404),
.B(n_300),
.Y(n_440)
);

INVx1_ASAP7_75t_L g441 ( 
.A(n_394),
.Y(n_441)
);

AND2x6_ASAP7_75t_L g442 ( 
.A(n_395),
.B(n_41),
.Y(n_442)
);

INVx2_ASAP7_75t_L g443 ( 
.A(n_371),
.Y(n_443)
);

INVx3_ASAP7_75t_L g444 ( 
.A(n_398),
.Y(n_444)
);

INVx1_ASAP7_75t_L g445 ( 
.A(n_380),
.Y(n_445)
);

AOI22xp5_ASAP7_75t_L g446 ( 
.A1(n_377),
.A2(n_303),
.B1(n_304),
.B2(n_302),
.Y(n_446)
);

NAND2xp5_ASAP7_75t_SL g447 ( 
.A(n_363),
.B(n_364),
.Y(n_447)
);

BUFx6f_ASAP7_75t_L g448 ( 
.A(n_398),
.Y(n_448)
);

AND2x2_ASAP7_75t_SL g449 ( 
.A(n_409),
.B(n_411),
.Y(n_449)
);

AND2x2_ASAP7_75t_L g450 ( 
.A(n_408),
.B(n_306),
.Y(n_450)
);

INVx4_ASAP7_75t_L g451 ( 
.A(n_398),
.Y(n_451)
);

AND2x2_ASAP7_75t_L g452 ( 
.A(n_408),
.B(n_308),
.Y(n_452)
);

BUFx3_ASAP7_75t_L g453 ( 
.A(n_390),
.Y(n_453)
);

AND2x2_ASAP7_75t_L g454 ( 
.A(n_408),
.B(n_312),
.Y(n_454)
);

INVx3_ASAP7_75t_L g455 ( 
.A(n_389),
.Y(n_455)
);

INVx2_ASAP7_75t_L g456 ( 
.A(n_373),
.Y(n_456)
);

INVx1_ASAP7_75t_L g457 ( 
.A(n_389),
.Y(n_457)
);

NAND2xp33_ASAP7_75t_L g458 ( 
.A(n_390),
.B(n_313),
.Y(n_458)
);

INVx5_ASAP7_75t_L g459 ( 
.A(n_390),
.Y(n_459)
);

INVx1_ASAP7_75t_L g460 ( 
.A(n_392),
.Y(n_460)
);

NAND2xp5_ASAP7_75t_L g461 ( 
.A(n_396),
.B(n_369),
.Y(n_461)
);

AND2x2_ASAP7_75t_L g462 ( 
.A(n_364),
.B(n_315),
.Y(n_462)
);

NAND2xp5_ASAP7_75t_L g463 ( 
.A(n_396),
.B(n_316),
.Y(n_463)
);

AND2x2_ASAP7_75t_L g464 ( 
.A(n_368),
.B(n_332),
.Y(n_464)
);

INVx1_ASAP7_75t_L g465 ( 
.A(n_392),
.Y(n_465)
);

NAND3xp33_ASAP7_75t_L g466 ( 
.A(n_384),
.B(n_332),
.C(n_3),
.Y(n_466)
);

AND2x6_ASAP7_75t_L g467 ( 
.A(n_396),
.B(n_43),
.Y(n_467)
);

INVx1_ASAP7_75t_L g468 ( 
.A(n_397),
.Y(n_468)
);

INVx5_ASAP7_75t_L g469 ( 
.A(n_397),
.Y(n_469)
);

INVx1_ASAP7_75t_L g470 ( 
.A(n_370),
.Y(n_470)
);

INVx5_ASAP7_75t_L g471 ( 
.A(n_411),
.Y(n_471)
);

AND2x4_ASAP7_75t_L g472 ( 
.A(n_410),
.B(n_368),
.Y(n_472)
);

INVx1_ASAP7_75t_L g473 ( 
.A(n_381),
.Y(n_473)
);

NAND2xp5_ASAP7_75t_L g474 ( 
.A(n_382),
.B(n_44),
.Y(n_474)
);

INVx1_ASAP7_75t_L g475 ( 
.A(n_384),
.Y(n_475)
);

AND2x2_ASAP7_75t_L g476 ( 
.A(n_406),
.B(n_3),
.Y(n_476)
);

AND2x4_ASAP7_75t_L g477 ( 
.A(n_406),
.B(n_45),
.Y(n_477)
);

OR2x2_ASAP7_75t_L g478 ( 
.A(n_423),
.B(n_407),
.Y(n_478)
);

INVx1_ASAP7_75t_L g479 ( 
.A(n_412),
.Y(n_479)
);

NAND2xp5_ASAP7_75t_SL g480 ( 
.A(n_419),
.B(n_376),
.Y(n_480)
);

AND2x4_ASAP7_75t_L g481 ( 
.A(n_436),
.B(n_411),
.Y(n_481)
);

NAND2xp5_ASAP7_75t_L g482 ( 
.A(n_419),
.B(n_46),
.Y(n_482)
);

NAND2xp5_ASAP7_75t_L g483 ( 
.A(n_415),
.B(n_47),
.Y(n_483)
);

NAND2xp5_ASAP7_75t_SL g484 ( 
.A(n_422),
.B(n_399),
.Y(n_484)
);

AND2x4_ASAP7_75t_L g485 ( 
.A(n_436),
.B(n_411),
.Y(n_485)
);

NAND2xp5_ASAP7_75t_L g486 ( 
.A(n_420),
.B(n_48),
.Y(n_486)
);

INVx2_ASAP7_75t_L g487 ( 
.A(n_455),
.Y(n_487)
);

AOI22xp5_ASAP7_75t_L g488 ( 
.A1(n_421),
.A2(n_399),
.B1(n_388),
.B2(n_383),
.Y(n_488)
);

NAND3xp33_ASAP7_75t_L g489 ( 
.A(n_425),
.B(n_388),
.C(n_383),
.Y(n_489)
);

NAND2xp5_ASAP7_75t_SL g490 ( 
.A(n_425),
.B(n_405),
.Y(n_490)
);

NAND2xp5_ASAP7_75t_SL g491 ( 
.A(n_430),
.B(n_405),
.Y(n_491)
);

NAND2xp5_ASAP7_75t_SL g492 ( 
.A(n_430),
.B(n_4),
.Y(n_492)
);

OR2x2_ASAP7_75t_L g493 ( 
.A(n_424),
.B(n_4),
.Y(n_493)
);

NAND2xp33_ASAP7_75t_L g494 ( 
.A(n_427),
.B(n_49),
.Y(n_494)
);

NOR2xp67_ASAP7_75t_L g495 ( 
.A(n_428),
.B(n_51),
.Y(n_495)
);

NOR2xp33_ASAP7_75t_L g496 ( 
.A(n_440),
.B(n_5),
.Y(n_496)
);

OR2x2_ASAP7_75t_SL g497 ( 
.A(n_466),
.B(n_5),
.Y(n_497)
);

INVx1_ASAP7_75t_L g498 ( 
.A(n_413),
.Y(n_498)
);

NAND2xp5_ASAP7_75t_L g499 ( 
.A(n_453),
.B(n_52),
.Y(n_499)
);

BUFx3_ASAP7_75t_L g500 ( 
.A(n_471),
.Y(n_500)
);

NAND2xp5_ASAP7_75t_SL g501 ( 
.A(n_477),
.B(n_6),
.Y(n_501)
);

INVx2_ASAP7_75t_L g502 ( 
.A(n_455),
.Y(n_502)
);

AOI22xp33_ASAP7_75t_L g503 ( 
.A1(n_442),
.A2(n_8),
.B1(n_6),
.B2(n_7),
.Y(n_503)
);

INVx2_ASAP7_75t_L g504 ( 
.A(n_433),
.Y(n_504)
);

NOR2xp33_ASAP7_75t_L g505 ( 
.A(n_440),
.B(n_7),
.Y(n_505)
);

INVx2_ASAP7_75t_L g506 ( 
.A(n_433),
.Y(n_506)
);

NOR2xp33_ASAP7_75t_L g507 ( 
.A(n_462),
.B(n_431),
.Y(n_507)
);

INVx2_ASAP7_75t_L g508 ( 
.A(n_438),
.Y(n_508)
);

NAND2xp5_ASAP7_75t_L g509 ( 
.A(n_453),
.B(n_53),
.Y(n_509)
);

OR2x6_ASAP7_75t_L g510 ( 
.A(n_472),
.B(n_9),
.Y(n_510)
);

NOR2xp33_ASAP7_75t_L g511 ( 
.A(n_446),
.B(n_9),
.Y(n_511)
);

NOR2x1p5_ASAP7_75t_L g512 ( 
.A(n_428),
.B(n_10),
.Y(n_512)
);

INVx2_ASAP7_75t_L g513 ( 
.A(n_438),
.Y(n_513)
);

OAI22xp33_ASAP7_75t_L g514 ( 
.A1(n_474),
.A2(n_12),
.B1(n_10),
.B2(n_11),
.Y(n_514)
);

NAND2xp5_ASAP7_75t_L g515 ( 
.A(n_416),
.B(n_54),
.Y(n_515)
);

INVx1_ASAP7_75t_L g516 ( 
.A(n_441),
.Y(n_516)
);

INVx2_ASAP7_75t_L g517 ( 
.A(n_439),
.Y(n_517)
);

INVx1_ASAP7_75t_L g518 ( 
.A(n_457),
.Y(n_518)
);

HB1xp67_ASAP7_75t_L g519 ( 
.A(n_471),
.Y(n_519)
);

OR2x2_ASAP7_75t_L g520 ( 
.A(n_475),
.B(n_11),
.Y(n_520)
);

OR2x6_ASAP7_75t_L g521 ( 
.A(n_472),
.B(n_12),
.Y(n_521)
);

INVx1_ASAP7_75t_L g522 ( 
.A(n_460),
.Y(n_522)
);

NAND2xp5_ASAP7_75t_L g523 ( 
.A(n_463),
.B(n_55),
.Y(n_523)
);

INVx2_ASAP7_75t_L g524 ( 
.A(n_439),
.Y(n_524)
);

O2A1O1Ixp33_ASAP7_75t_L g525 ( 
.A1(n_421),
.A2(n_458),
.B(n_414),
.C(n_429),
.Y(n_525)
);

NAND2xp5_ASAP7_75t_L g526 ( 
.A(n_429),
.B(n_56),
.Y(n_526)
);

NAND2xp5_ASAP7_75t_L g527 ( 
.A(n_459),
.B(n_58),
.Y(n_527)
);

NAND2xp5_ASAP7_75t_L g528 ( 
.A(n_459),
.B(n_59),
.Y(n_528)
);

AOI22xp5_ASAP7_75t_L g529 ( 
.A1(n_427),
.A2(n_155),
.B1(n_253),
.B2(n_252),
.Y(n_529)
);

NAND2xp5_ASAP7_75t_L g530 ( 
.A(n_459),
.B(n_60),
.Y(n_530)
);

INVx1_ASAP7_75t_L g531 ( 
.A(n_465),
.Y(n_531)
);

AOI22xp5_ASAP7_75t_L g532 ( 
.A1(n_427),
.A2(n_445),
.B1(n_414),
.B2(n_458),
.Y(n_532)
);

HB1xp67_ASAP7_75t_L g533 ( 
.A(n_471),
.Y(n_533)
);

INVx3_ASAP7_75t_L g534 ( 
.A(n_448),
.Y(n_534)
);

INVx2_ASAP7_75t_L g535 ( 
.A(n_443),
.Y(n_535)
);

NAND2xp5_ASAP7_75t_L g536 ( 
.A(n_444),
.B(n_461),
.Y(n_536)
);

NOR2x1_ASAP7_75t_L g537 ( 
.A(n_473),
.B(n_62),
.Y(n_537)
);

AND2x4_ASAP7_75t_L g538 ( 
.A(n_471),
.B(n_63),
.Y(n_538)
);

INVx2_ASAP7_75t_SL g539 ( 
.A(n_449),
.Y(n_539)
);

NAND2xp5_ASAP7_75t_L g540 ( 
.A(n_444),
.B(n_65),
.Y(n_540)
);

NOR3xp33_ASAP7_75t_L g541 ( 
.A(n_464),
.B(n_13),
.C(n_14),
.Y(n_541)
);

NAND2xp5_ASAP7_75t_L g542 ( 
.A(n_470),
.B(n_67),
.Y(n_542)
);

NAND2xp5_ASAP7_75t_L g543 ( 
.A(n_451),
.B(n_68),
.Y(n_543)
);

NAND2xp5_ASAP7_75t_L g544 ( 
.A(n_459),
.B(n_69),
.Y(n_544)
);

AOI22xp33_ASAP7_75t_SL g545 ( 
.A1(n_449),
.A2(n_477),
.B1(n_437),
.B2(n_476),
.Y(n_545)
);

INVx2_ASAP7_75t_L g546 ( 
.A(n_443),
.Y(n_546)
);

NAND2xp5_ASAP7_75t_SL g547 ( 
.A(n_477),
.B(n_13),
.Y(n_547)
);

INVx4_ASAP7_75t_L g548 ( 
.A(n_448),
.Y(n_548)
);

INVx2_ASAP7_75t_SL g549 ( 
.A(n_450),
.Y(n_549)
);

NAND2x1p5_ASAP7_75t_L g550 ( 
.A(n_451),
.B(n_434),
.Y(n_550)
);

BUFx4f_ASAP7_75t_L g551 ( 
.A(n_481),
.Y(n_551)
);

INVx1_ASAP7_75t_L g552 ( 
.A(n_504),
.Y(n_552)
);

AOI22xp33_ASAP7_75t_L g553 ( 
.A1(n_496),
.A2(n_442),
.B1(n_467),
.B2(n_427),
.Y(n_553)
);

AOI21xp5_ASAP7_75t_L g554 ( 
.A1(n_536),
.A2(n_434),
.B(n_418),
.Y(n_554)
);

OAI22xp5_ASAP7_75t_L g555 ( 
.A1(n_482),
.A2(n_454),
.B1(n_452),
.B2(n_447),
.Y(n_555)
);

AOI22xp5_ASAP7_75t_L g556 ( 
.A1(n_507),
.A2(n_427),
.B1(n_447),
.B2(n_435),
.Y(n_556)
);

BUFx6f_ASAP7_75t_L g557 ( 
.A(n_500),
.Y(n_557)
);

AOI21xp5_ASAP7_75t_L g558 ( 
.A1(n_550),
.A2(n_482),
.B(n_525),
.Y(n_558)
);

NAND2xp5_ASAP7_75t_L g559 ( 
.A(n_479),
.B(n_468),
.Y(n_559)
);

NAND2xp5_ASAP7_75t_L g560 ( 
.A(n_498),
.B(n_456),
.Y(n_560)
);

OAI21x1_ASAP7_75t_L g561 ( 
.A1(n_540),
.A2(n_534),
.B(n_509),
.Y(n_561)
);

NAND2xp5_ASAP7_75t_SL g562 ( 
.A(n_539),
.B(n_448),
.Y(n_562)
);

INVx2_ASAP7_75t_L g563 ( 
.A(n_506),
.Y(n_563)
);

NAND2xp5_ASAP7_75t_SL g564 ( 
.A(n_545),
.B(n_448),
.Y(n_564)
);

AOI21xp5_ASAP7_75t_L g565 ( 
.A1(n_550),
.A2(n_418),
.B(n_432),
.Y(n_565)
);

NOR2xp33_ASAP7_75t_L g566 ( 
.A(n_480),
.B(n_456),
.Y(n_566)
);

O2A1O1Ixp33_ASAP7_75t_SL g567 ( 
.A1(n_492),
.A2(n_417),
.B(n_426),
.C(n_467),
.Y(n_567)
);

NOR2xp33_ASAP7_75t_L g568 ( 
.A(n_478),
.B(n_417),
.Y(n_568)
);

AOI21xp5_ASAP7_75t_L g569 ( 
.A1(n_548),
.A2(n_432),
.B(n_426),
.Y(n_569)
);

NOR2x1_ASAP7_75t_L g570 ( 
.A(n_495),
.B(n_432),
.Y(n_570)
);

NAND2xp5_ASAP7_75t_L g571 ( 
.A(n_516),
.B(n_432),
.Y(n_571)
);

INVx2_ASAP7_75t_L g572 ( 
.A(n_508),
.Y(n_572)
);

AOI21xp5_ASAP7_75t_L g573 ( 
.A1(n_548),
.A2(n_526),
.B(n_486),
.Y(n_573)
);

AOI21xp5_ASAP7_75t_L g574 ( 
.A1(n_526),
.A2(n_469),
.B(n_467),
.Y(n_574)
);

NAND2xp5_ASAP7_75t_SL g575 ( 
.A(n_549),
.B(n_481),
.Y(n_575)
);

AOI21xp5_ASAP7_75t_L g576 ( 
.A1(n_483),
.A2(n_469),
.B(n_467),
.Y(n_576)
);

INVx1_ASAP7_75t_L g577 ( 
.A(n_513),
.Y(n_577)
);

INVx2_ASAP7_75t_L g578 ( 
.A(n_517),
.Y(n_578)
);

NOR2xp33_ASAP7_75t_L g579 ( 
.A(n_484),
.B(n_469),
.Y(n_579)
);

NOR2xp33_ASAP7_75t_L g580 ( 
.A(n_490),
.B(n_469),
.Y(n_580)
);

OAI21xp5_ASAP7_75t_L g581 ( 
.A1(n_483),
.A2(n_467),
.B(n_442),
.Y(n_581)
);

AOI21xp5_ASAP7_75t_L g582 ( 
.A1(n_486),
.A2(n_442),
.B(n_72),
.Y(n_582)
);

AOI21xp5_ASAP7_75t_L g583 ( 
.A1(n_494),
.A2(n_538),
.B(n_523),
.Y(n_583)
);

INVx3_ASAP7_75t_L g584 ( 
.A(n_534),
.Y(n_584)
);

OAI22xp5_ASAP7_75t_L g585 ( 
.A1(n_532),
.A2(n_442),
.B1(n_159),
.B2(n_160),
.Y(n_585)
);

OAI22xp5_ASAP7_75t_L g586 ( 
.A1(n_503),
.A2(n_158),
.B1(n_251),
.B2(n_250),
.Y(n_586)
);

AOI21xp5_ASAP7_75t_L g587 ( 
.A1(n_538),
.A2(n_73),
.B(n_71),
.Y(n_587)
);

OAI21xp5_ASAP7_75t_L g588 ( 
.A1(n_505),
.A2(n_76),
.B(n_74),
.Y(n_588)
);

AND2x2_ASAP7_75t_L g589 ( 
.A(n_485),
.B(n_493),
.Y(n_589)
);

AND2x2_ASAP7_75t_L g590 ( 
.A(n_485),
.B(n_14),
.Y(n_590)
);

OR2x2_ASAP7_75t_L g591 ( 
.A(n_491),
.B(n_15),
.Y(n_591)
);

INVx1_ASAP7_75t_L g592 ( 
.A(n_524),
.Y(n_592)
);

O2A1O1Ixp33_ASAP7_75t_L g593 ( 
.A1(n_501),
.A2(n_15),
.B(n_16),
.C(n_17),
.Y(n_593)
);

NAND2xp5_ASAP7_75t_L g594 ( 
.A(n_518),
.B(n_16),
.Y(n_594)
);

AOI21xp5_ASAP7_75t_L g595 ( 
.A1(n_543),
.A2(n_78),
.B(n_77),
.Y(n_595)
);

AOI21xp5_ASAP7_75t_L g596 ( 
.A1(n_499),
.A2(n_83),
.B(n_80),
.Y(n_596)
);

NOR3xp33_ASAP7_75t_L g597 ( 
.A(n_489),
.B(n_511),
.C(n_488),
.Y(n_597)
);

OAI21x1_ASAP7_75t_L g598 ( 
.A1(n_535),
.A2(n_86),
.B(n_84),
.Y(n_598)
);

AOI21x1_ASAP7_75t_L g599 ( 
.A1(n_546),
.A2(n_88),
.B(n_87),
.Y(n_599)
);

AOI21xp5_ASAP7_75t_L g600 ( 
.A1(n_515),
.A2(n_542),
.B(n_502),
.Y(n_600)
);

AOI21xp5_ASAP7_75t_L g601 ( 
.A1(n_487),
.A2(n_91),
.B(n_89),
.Y(n_601)
);

AOI21xp5_ASAP7_75t_L g602 ( 
.A1(n_522),
.A2(n_93),
.B(n_92),
.Y(n_602)
);

CKINVDCx5p33_ASAP7_75t_R g603 ( 
.A(n_510),
.Y(n_603)
);

OAI22xp5_ASAP7_75t_L g604 ( 
.A1(n_547),
.A2(n_17),
.B1(n_18),
.B2(n_19),
.Y(n_604)
);

NAND2xp5_ASAP7_75t_L g605 ( 
.A(n_531),
.B(n_20),
.Y(n_605)
);

OAI22xp5_ASAP7_75t_L g606 ( 
.A1(n_497),
.A2(n_20),
.B1(n_21),
.B2(n_22),
.Y(n_606)
);

AOI22xp5_ASAP7_75t_L g607 ( 
.A1(n_537),
.A2(n_173),
.B1(n_249),
.B2(n_247),
.Y(n_607)
);

NAND2xp5_ASAP7_75t_L g608 ( 
.A(n_519),
.B(n_533),
.Y(n_608)
);

NOR2xp33_ASAP7_75t_L g609 ( 
.A(n_489),
.B(n_22),
.Y(n_609)
);

NOR2xp33_ASAP7_75t_L g610 ( 
.A(n_520),
.B(n_23),
.Y(n_610)
);

OAI21xp5_ASAP7_75t_L g611 ( 
.A1(n_529),
.A2(n_95),
.B(n_94),
.Y(n_611)
);

INVx2_ASAP7_75t_L g612 ( 
.A(n_527),
.Y(n_612)
);

NOR2xp67_ASAP7_75t_SL g613 ( 
.A(n_611),
.B(n_527),
.Y(n_613)
);

AOI21xp5_ASAP7_75t_L g614 ( 
.A1(n_583),
.A2(n_530),
.B(n_528),
.Y(n_614)
);

HB1xp67_ASAP7_75t_L g615 ( 
.A(n_589),
.Y(n_615)
);

INVx1_ASAP7_75t_L g616 ( 
.A(n_552),
.Y(n_616)
);

AO21x1_ASAP7_75t_L g617 ( 
.A1(n_555),
.A2(n_514),
.B(n_528),
.Y(n_617)
);

A2O1A1Ixp33_ASAP7_75t_L g618 ( 
.A1(n_597),
.A2(n_541),
.B(n_544),
.C(n_530),
.Y(n_618)
);

INVx2_ASAP7_75t_L g619 ( 
.A(n_563),
.Y(n_619)
);

OAI21x1_ASAP7_75t_L g620 ( 
.A1(n_561),
.A2(n_544),
.B(n_512),
.Y(n_620)
);

NAND2xp5_ASAP7_75t_L g621 ( 
.A(n_612),
.B(n_510),
.Y(n_621)
);

OAI21x1_ASAP7_75t_L g622 ( 
.A1(n_565),
.A2(n_99),
.B(n_97),
.Y(n_622)
);

O2A1O1Ixp5_ASAP7_75t_L g623 ( 
.A1(n_558),
.A2(n_521),
.B(n_510),
.C(n_176),
.Y(n_623)
);

INVx2_ASAP7_75t_L g624 ( 
.A(n_572),
.Y(n_624)
);

OAI21xp5_ASAP7_75t_L g625 ( 
.A1(n_581),
.A2(n_521),
.B(n_102),
.Y(n_625)
);

OAI22xp5_ASAP7_75t_L g626 ( 
.A1(n_553),
.A2(n_521),
.B1(n_24),
.B2(n_25),
.Y(n_626)
);

INVx1_ASAP7_75t_L g627 ( 
.A(n_577),
.Y(n_627)
);

OAI21x1_ASAP7_75t_L g628 ( 
.A1(n_600),
.A2(n_105),
.B(n_100),
.Y(n_628)
);

INVx1_ASAP7_75t_L g629 ( 
.A(n_592),
.Y(n_629)
);

AOI21x1_ASAP7_75t_L g630 ( 
.A1(n_573),
.A2(n_107),
.B(n_106),
.Y(n_630)
);

INVx3_ASAP7_75t_L g631 ( 
.A(n_584),
.Y(n_631)
);

OAI21x1_ASAP7_75t_L g632 ( 
.A1(n_574),
.A2(n_569),
.B(n_576),
.Y(n_632)
);

OAI21x1_ASAP7_75t_SL g633 ( 
.A1(n_588),
.A2(n_587),
.B(n_611),
.Y(n_633)
);

OAI21x1_ASAP7_75t_L g634 ( 
.A1(n_554),
.A2(n_109),
.B(n_108),
.Y(n_634)
);

AO22x1_ASAP7_75t_L g635 ( 
.A1(n_609),
.A2(n_23),
.B1(n_24),
.B2(n_25),
.Y(n_635)
);

A2O1A1Ixp33_ASAP7_75t_L g636 ( 
.A1(n_610),
.A2(n_26),
.B(n_27),
.C(n_28),
.Y(n_636)
);

OAI21x1_ASAP7_75t_L g637 ( 
.A1(n_598),
.A2(n_581),
.B(n_599),
.Y(n_637)
);

INVx2_ASAP7_75t_L g638 ( 
.A(n_578),
.Y(n_638)
);

AOI22xp5_ASAP7_75t_L g639 ( 
.A1(n_556),
.A2(n_181),
.B1(n_246),
.B2(n_243),
.Y(n_639)
);

OAI21x1_ASAP7_75t_L g640 ( 
.A1(n_582),
.A2(n_180),
.B(n_242),
.Y(n_640)
);

NAND2xp5_ASAP7_75t_L g641 ( 
.A(n_566),
.B(n_110),
.Y(n_641)
);

AOI21xp5_ASAP7_75t_L g642 ( 
.A1(n_567),
.A2(n_179),
.B(n_241),
.Y(n_642)
);

INVx1_ASAP7_75t_L g643 ( 
.A(n_560),
.Y(n_643)
);

OA21x2_ASAP7_75t_L g644 ( 
.A1(n_588),
.A2(n_178),
.B(n_240),
.Y(n_644)
);

NOR2xp33_ASAP7_75t_L g645 ( 
.A(n_591),
.B(n_27),
.Y(n_645)
);

AOI21xp5_ASAP7_75t_SL g646 ( 
.A1(n_585),
.A2(n_182),
.B(n_239),
.Y(n_646)
);

AND2x2_ASAP7_75t_L g647 ( 
.A(n_568),
.B(n_28),
.Y(n_647)
);

NAND2xp33_ASAP7_75t_L g648 ( 
.A(n_586),
.B(n_111),
.Y(n_648)
);

AND2x6_ASAP7_75t_L g649 ( 
.A(n_590),
.B(n_112),
.Y(n_649)
);

AO21x2_ASAP7_75t_L g650 ( 
.A1(n_564),
.A2(n_580),
.B(n_571),
.Y(n_650)
);

OAI21x1_ASAP7_75t_L g651 ( 
.A1(n_584),
.A2(n_570),
.B(n_559),
.Y(n_651)
);

AND2x4_ASAP7_75t_L g652 ( 
.A(n_575),
.B(n_113),
.Y(n_652)
);

OAI21x1_ASAP7_75t_L g653 ( 
.A1(n_596),
.A2(n_595),
.B(n_562),
.Y(n_653)
);

NAND2xp5_ASAP7_75t_L g654 ( 
.A(n_551),
.B(n_114),
.Y(n_654)
);

NAND2xp5_ASAP7_75t_L g655 ( 
.A(n_551),
.B(n_115),
.Y(n_655)
);

NAND2x1p5_ASAP7_75t_L g656 ( 
.A(n_557),
.B(n_117),
.Y(n_656)
);

AOI21xp5_ASAP7_75t_L g657 ( 
.A1(n_579),
.A2(n_185),
.B(n_238),
.Y(n_657)
);

AND2x2_ASAP7_75t_L g658 ( 
.A(n_557),
.B(n_29),
.Y(n_658)
);

BUFx3_ASAP7_75t_L g659 ( 
.A(n_557),
.Y(n_659)
);

OAI22xp5_ASAP7_75t_L g660 ( 
.A1(n_606),
.A2(n_29),
.B1(n_30),
.B2(n_31),
.Y(n_660)
);

OAI21xp5_ASAP7_75t_L g661 ( 
.A1(n_594),
.A2(n_187),
.B(n_236),
.Y(n_661)
);

OAI21x1_ASAP7_75t_L g662 ( 
.A1(n_601),
.A2(n_184),
.B(n_235),
.Y(n_662)
);

NAND2xp5_ASAP7_75t_L g663 ( 
.A(n_605),
.B(n_604),
.Y(n_663)
);

AOI21xp5_ASAP7_75t_L g664 ( 
.A1(n_602),
.A2(n_183),
.B(n_232),
.Y(n_664)
);

NOR2xp33_ASAP7_75t_L g665 ( 
.A(n_608),
.B(n_30),
.Y(n_665)
);

AND2x2_ASAP7_75t_L g666 ( 
.A(n_603),
.B(n_31),
.Y(n_666)
);

AO21x2_ASAP7_75t_L g667 ( 
.A1(n_607),
.A2(n_188),
.B(n_231),
.Y(n_667)
);

BUFx6f_ASAP7_75t_L g668 ( 
.A(n_593),
.Y(n_668)
);

INVx1_ASAP7_75t_L g669 ( 
.A(n_604),
.Y(n_669)
);

AOI21xp5_ASAP7_75t_L g670 ( 
.A1(n_606),
.A2(n_177),
.B(n_230),
.Y(n_670)
);

AND2x2_ASAP7_75t_L g671 ( 
.A(n_589),
.B(n_32),
.Y(n_671)
);

INVx3_ASAP7_75t_L g672 ( 
.A(n_584),
.Y(n_672)
);

INVx2_ASAP7_75t_L g673 ( 
.A(n_616),
.Y(n_673)
);

NOR2xp33_ASAP7_75t_L g674 ( 
.A(n_615),
.B(n_32),
.Y(n_674)
);

NAND2xp5_ASAP7_75t_L g675 ( 
.A(n_643),
.B(n_33),
.Y(n_675)
);

INVx1_ASAP7_75t_L g676 ( 
.A(n_627),
.Y(n_676)
);

BUFx6f_ASAP7_75t_L g677 ( 
.A(n_659),
.Y(n_677)
);

INVx6_ASAP7_75t_L g678 ( 
.A(n_658),
.Y(n_678)
);

NAND2xp5_ASAP7_75t_L g679 ( 
.A(n_669),
.B(n_33),
.Y(n_679)
);

AND2x4_ASAP7_75t_L g680 ( 
.A(n_652),
.B(n_629),
.Y(n_680)
);

AOI21xp33_ASAP7_75t_SL g681 ( 
.A1(n_645),
.A2(n_34),
.B(n_35),
.Y(n_681)
);

INVx1_ASAP7_75t_L g682 ( 
.A(n_619),
.Y(n_682)
);

BUFx12f_ASAP7_75t_L g683 ( 
.A(n_656),
.Y(n_683)
);

INVx1_ASAP7_75t_L g684 ( 
.A(n_624),
.Y(n_684)
);

INVx1_ASAP7_75t_L g685 ( 
.A(n_638),
.Y(n_685)
);

AOI21xp5_ASAP7_75t_L g686 ( 
.A1(n_614),
.A2(n_189),
.B(n_229),
.Y(n_686)
);

AND2x4_ASAP7_75t_L g687 ( 
.A(n_652),
.B(n_118),
.Y(n_687)
);

INVx2_ASAP7_75t_L g688 ( 
.A(n_631),
.Y(n_688)
);

INVx3_ASAP7_75t_SL g689 ( 
.A(n_666),
.Y(n_689)
);

O2A1O1Ixp33_ASAP7_75t_L g690 ( 
.A1(n_663),
.A2(n_34),
.B(n_35),
.C(n_36),
.Y(n_690)
);

INVx3_ASAP7_75t_L g691 ( 
.A(n_631),
.Y(n_691)
);

OR2x2_ASAP7_75t_L g692 ( 
.A(n_621),
.B(n_36),
.Y(n_692)
);

INVx2_ASAP7_75t_L g693 ( 
.A(n_672),
.Y(n_693)
);

AOI22xp5_ASAP7_75t_L g694 ( 
.A1(n_648),
.A2(n_37),
.B1(n_38),
.B2(n_39),
.Y(n_694)
);

BUFx6f_ASAP7_75t_SL g695 ( 
.A(n_649),
.Y(n_695)
);

INVx8_ASAP7_75t_L g696 ( 
.A(n_649),
.Y(n_696)
);

INVx5_ASAP7_75t_L g697 ( 
.A(n_649),
.Y(n_697)
);

AND2x4_ASAP7_75t_L g698 ( 
.A(n_671),
.B(n_120),
.Y(n_698)
);

AOI21xp5_ASAP7_75t_L g699 ( 
.A1(n_614),
.A2(n_193),
.B(n_228),
.Y(n_699)
);

OAI21xp33_ASAP7_75t_L g700 ( 
.A1(n_663),
.A2(n_37),
.B(n_38),
.Y(n_700)
);

AOI22xp33_ASAP7_75t_SL g701 ( 
.A1(n_626),
.A2(n_39),
.B1(n_40),
.B2(n_122),
.Y(n_701)
);

INVx2_ASAP7_75t_SL g702 ( 
.A(n_621),
.Y(n_702)
);

BUFx3_ASAP7_75t_L g703 ( 
.A(n_656),
.Y(n_703)
);

AOI21xp5_ASAP7_75t_L g704 ( 
.A1(n_633),
.A2(n_195),
.B(n_124),
.Y(n_704)
);

HB1xp67_ASAP7_75t_L g705 ( 
.A(n_672),
.Y(n_705)
);

NAND2xp5_ASAP7_75t_L g706 ( 
.A(n_647),
.B(n_40),
.Y(n_706)
);

INVx5_ASAP7_75t_L g707 ( 
.A(n_649),
.Y(n_707)
);

INVxp67_ASAP7_75t_L g708 ( 
.A(n_665),
.Y(n_708)
);

AND2x2_ASAP7_75t_L g709 ( 
.A(n_636),
.B(n_125),
.Y(n_709)
);

AOI21xp5_ASAP7_75t_L g710 ( 
.A1(n_618),
.A2(n_126),
.B(n_127),
.Y(n_710)
);

INVx5_ASAP7_75t_L g711 ( 
.A(n_668),
.Y(n_711)
);

BUFx2_ASAP7_75t_L g712 ( 
.A(n_625),
.Y(n_712)
);

INVx3_ASAP7_75t_SL g713 ( 
.A(n_668),
.Y(n_713)
);

NAND2xp5_ASAP7_75t_SL g714 ( 
.A(n_668),
.B(n_128),
.Y(n_714)
);

INVx2_ASAP7_75t_L g715 ( 
.A(n_651),
.Y(n_715)
);

INVx1_ASAP7_75t_L g716 ( 
.A(n_650),
.Y(n_716)
);

AND2x2_ASAP7_75t_L g717 ( 
.A(n_625),
.B(n_129),
.Y(n_717)
);

NAND2xp5_ASAP7_75t_L g718 ( 
.A(n_641),
.B(n_130),
.Y(n_718)
);

HB1xp67_ASAP7_75t_L g719 ( 
.A(n_626),
.Y(n_719)
);

NAND2xp5_ASAP7_75t_L g720 ( 
.A(n_641),
.B(n_132),
.Y(n_720)
);

BUFx6f_ASAP7_75t_L g721 ( 
.A(n_654),
.Y(n_721)
);

AOI21xp5_ASAP7_75t_L g722 ( 
.A1(n_653),
.A2(n_134),
.B(n_136),
.Y(n_722)
);

AND2x2_ASAP7_75t_L g723 ( 
.A(n_660),
.B(n_138),
.Y(n_723)
);

BUFx6f_ASAP7_75t_L g724 ( 
.A(n_654),
.Y(n_724)
);

AOI22xp5_ASAP7_75t_L g725 ( 
.A1(n_708),
.A2(n_613),
.B1(n_660),
.B2(n_639),
.Y(n_725)
);

BUFx12f_ASAP7_75t_L g726 ( 
.A(n_677),
.Y(n_726)
);

BUFx12f_ASAP7_75t_L g727 ( 
.A(n_677),
.Y(n_727)
);

INVx6_ASAP7_75t_L g728 ( 
.A(n_711),
.Y(n_728)
);

INVx1_ASAP7_75t_L g729 ( 
.A(n_676),
.Y(n_729)
);

INVx1_ASAP7_75t_L g730 ( 
.A(n_676),
.Y(n_730)
);

AOI22xp33_ASAP7_75t_L g731 ( 
.A1(n_719),
.A2(n_617),
.B1(n_670),
.B2(n_661),
.Y(n_731)
);

OAI22xp5_ASAP7_75t_SL g732 ( 
.A1(n_701),
.A2(n_644),
.B1(n_661),
.B2(n_635),
.Y(n_732)
);

OAI21xp5_ASAP7_75t_L g733 ( 
.A1(n_718),
.A2(n_623),
.B(n_670),
.Y(n_733)
);

INVx1_ASAP7_75t_L g734 ( 
.A(n_673),
.Y(n_734)
);

INVx6_ASAP7_75t_L g735 ( 
.A(n_711),
.Y(n_735)
);

AOI22xp33_ASAP7_75t_SL g736 ( 
.A1(n_712),
.A2(n_717),
.B1(n_709),
.B2(n_695),
.Y(n_736)
);

INVx1_ASAP7_75t_L g737 ( 
.A(n_682),
.Y(n_737)
);

AND2x2_ASAP7_75t_L g738 ( 
.A(n_680),
.B(n_655),
.Y(n_738)
);

INVx1_ASAP7_75t_L g739 ( 
.A(n_682),
.Y(n_739)
);

INVx2_ASAP7_75t_L g740 ( 
.A(n_684),
.Y(n_740)
);

INVx2_ASAP7_75t_L g741 ( 
.A(n_684),
.Y(n_741)
);

INVx1_ASAP7_75t_L g742 ( 
.A(n_685),
.Y(n_742)
);

INVx1_ASAP7_75t_L g743 ( 
.A(n_685),
.Y(n_743)
);

INVx2_ASAP7_75t_L g744 ( 
.A(n_716),
.Y(n_744)
);

INVx2_ASAP7_75t_L g745 ( 
.A(n_716),
.Y(n_745)
);

AOI22xp33_ASAP7_75t_L g746 ( 
.A1(n_700),
.A2(n_644),
.B1(n_667),
.B2(n_650),
.Y(n_746)
);

INVx2_ASAP7_75t_SL g747 ( 
.A(n_677),
.Y(n_747)
);

INVx1_ASAP7_75t_L g748 ( 
.A(n_711),
.Y(n_748)
);

INVx1_ASAP7_75t_L g749 ( 
.A(n_702),
.Y(n_749)
);

INVx1_ASAP7_75t_L g750 ( 
.A(n_705),
.Y(n_750)
);

BUFx3_ASAP7_75t_L g751 ( 
.A(n_713),
.Y(n_751)
);

AO21x2_ASAP7_75t_L g752 ( 
.A1(n_715),
.A2(n_642),
.B(n_632),
.Y(n_752)
);

INVx1_ASAP7_75t_L g753 ( 
.A(n_675),
.Y(n_753)
);

NAND2x1p5_ASAP7_75t_L g754 ( 
.A(n_697),
.B(n_707),
.Y(n_754)
);

BUFx12f_ASAP7_75t_L g755 ( 
.A(n_678),
.Y(n_755)
);

INVx1_ASAP7_75t_L g756 ( 
.A(n_679),
.Y(n_756)
);

AOI22xp33_ASAP7_75t_SL g757 ( 
.A1(n_695),
.A2(n_667),
.B1(n_655),
.B2(n_657),
.Y(n_757)
);

INVx1_ASAP7_75t_L g758 ( 
.A(n_688),
.Y(n_758)
);

INVx2_ASAP7_75t_L g759 ( 
.A(n_691),
.Y(n_759)
);

CKINVDCx5p33_ASAP7_75t_R g760 ( 
.A(n_689),
.Y(n_760)
);

INVx2_ASAP7_75t_L g761 ( 
.A(n_691),
.Y(n_761)
);

INVx1_ASAP7_75t_L g762 ( 
.A(n_693),
.Y(n_762)
);

INVx3_ASAP7_75t_L g763 ( 
.A(n_696),
.Y(n_763)
);

AOI22xp33_ASAP7_75t_L g764 ( 
.A1(n_723),
.A2(n_657),
.B1(n_664),
.B2(n_642),
.Y(n_764)
);

INVx1_ASAP7_75t_L g765 ( 
.A(n_680),
.Y(n_765)
);

INVx2_ASAP7_75t_L g766 ( 
.A(n_721),
.Y(n_766)
);

INVx2_ASAP7_75t_L g767 ( 
.A(n_721),
.Y(n_767)
);

BUFx8_ASAP7_75t_L g768 ( 
.A(n_683),
.Y(n_768)
);

CKINVDCx11_ASAP7_75t_R g769 ( 
.A(n_696),
.Y(n_769)
);

INVx1_ASAP7_75t_L g770 ( 
.A(n_692),
.Y(n_770)
);

AOI22xp33_ASAP7_75t_L g771 ( 
.A1(n_694),
.A2(n_664),
.B1(n_640),
.B2(n_662),
.Y(n_771)
);

AOI22xp33_ASAP7_75t_L g772 ( 
.A1(n_706),
.A2(n_620),
.B1(n_628),
.B2(n_634),
.Y(n_772)
);

NAND2xp5_ASAP7_75t_L g773 ( 
.A(n_687),
.B(n_646),
.Y(n_773)
);

BUFx2_ASAP7_75t_R g774 ( 
.A(n_703),
.Y(n_774)
);

INVx1_ASAP7_75t_L g775 ( 
.A(n_690),
.Y(n_775)
);

OAI22xp5_ASAP7_75t_L g776 ( 
.A1(n_697),
.A2(n_630),
.B1(n_637),
.B2(n_622),
.Y(n_776)
);

AOI22xp33_ASAP7_75t_L g777 ( 
.A1(n_687),
.A2(n_714),
.B1(n_674),
.B2(n_710),
.Y(n_777)
);

OR2x2_ASAP7_75t_L g778 ( 
.A(n_698),
.B(n_139),
.Y(n_778)
);

HB1xp67_ASAP7_75t_L g779 ( 
.A(n_721),
.Y(n_779)
);

HB1xp67_ASAP7_75t_L g780 ( 
.A(n_724),
.Y(n_780)
);

INVx1_ASAP7_75t_L g781 ( 
.A(n_724),
.Y(n_781)
);

BUFx6f_ASAP7_75t_L g782 ( 
.A(n_697),
.Y(n_782)
);

INVx2_ASAP7_75t_L g783 ( 
.A(n_724),
.Y(n_783)
);

OAI21xp5_ASAP7_75t_L g784 ( 
.A1(n_720),
.A2(n_699),
.B(n_686),
.Y(n_784)
);

OR2x2_ASAP7_75t_L g785 ( 
.A(n_698),
.B(n_140),
.Y(n_785)
);

INVx2_ASAP7_75t_L g786 ( 
.A(n_707),
.Y(n_786)
);

INVxp67_ASAP7_75t_SL g787 ( 
.A(n_750),
.Y(n_787)
);

AND2x2_ASAP7_75t_L g788 ( 
.A(n_744),
.B(n_681),
.Y(n_788)
);

INVx1_ASAP7_75t_L g789 ( 
.A(n_744),
.Y(n_789)
);

INVx2_ASAP7_75t_L g790 ( 
.A(n_745),
.Y(n_790)
);

INVx1_ASAP7_75t_L g791 ( 
.A(n_745),
.Y(n_791)
);

INVx1_ASAP7_75t_L g792 ( 
.A(n_729),
.Y(n_792)
);

INVx1_ASAP7_75t_L g793 ( 
.A(n_730),
.Y(n_793)
);

INVx1_ASAP7_75t_L g794 ( 
.A(n_740),
.Y(n_794)
);

INVx1_ASAP7_75t_L g795 ( 
.A(n_740),
.Y(n_795)
);

NAND2x1p5_ASAP7_75t_L g796 ( 
.A(n_782),
.B(n_707),
.Y(n_796)
);

INVxp67_ASAP7_75t_SL g797 ( 
.A(n_779),
.Y(n_797)
);

AO21x2_ASAP7_75t_L g798 ( 
.A1(n_784),
.A2(n_722),
.B(n_704),
.Y(n_798)
);

INVx1_ASAP7_75t_L g799 ( 
.A(n_741),
.Y(n_799)
);

INVx1_ASAP7_75t_L g800 ( 
.A(n_741),
.Y(n_800)
);

OA21x2_ASAP7_75t_L g801 ( 
.A1(n_733),
.A2(n_681),
.B(n_143),
.Y(n_801)
);

INVx1_ASAP7_75t_L g802 ( 
.A(n_737),
.Y(n_802)
);

INVx2_ASAP7_75t_L g803 ( 
.A(n_739),
.Y(n_803)
);

AND2x4_ASAP7_75t_L g804 ( 
.A(n_766),
.B(n_141),
.Y(n_804)
);

AND2x2_ASAP7_75t_L g805 ( 
.A(n_766),
.B(n_767),
.Y(n_805)
);

AND2x4_ASAP7_75t_L g806 ( 
.A(n_767),
.B(n_144),
.Y(n_806)
);

INVx2_ASAP7_75t_L g807 ( 
.A(n_742),
.Y(n_807)
);

INVx1_ASAP7_75t_L g808 ( 
.A(n_743),
.Y(n_808)
);

INVx1_ASAP7_75t_L g809 ( 
.A(n_734),
.Y(n_809)
);

NAND2xp5_ASAP7_75t_L g810 ( 
.A(n_756),
.B(n_678),
.Y(n_810)
);

INVx1_ASAP7_75t_L g811 ( 
.A(n_770),
.Y(n_811)
);

INVx2_ASAP7_75t_L g812 ( 
.A(n_752),
.Y(n_812)
);

INVx1_ASAP7_75t_L g813 ( 
.A(n_749),
.Y(n_813)
);

INVx1_ASAP7_75t_L g814 ( 
.A(n_752),
.Y(n_814)
);

HB1xp67_ASAP7_75t_L g815 ( 
.A(n_779),
.Y(n_815)
);

HB1xp67_ASAP7_75t_L g816 ( 
.A(n_780),
.Y(n_816)
);

INVx2_ASAP7_75t_L g817 ( 
.A(n_759),
.Y(n_817)
);

INVx1_ASAP7_75t_L g818 ( 
.A(n_759),
.Y(n_818)
);

INVx1_ASAP7_75t_L g819 ( 
.A(n_761),
.Y(n_819)
);

INVx1_ASAP7_75t_L g820 ( 
.A(n_761),
.Y(n_820)
);

INVx2_ASAP7_75t_L g821 ( 
.A(n_758),
.Y(n_821)
);

BUFx8_ASAP7_75t_L g822 ( 
.A(n_726),
.Y(n_822)
);

INVx1_ASAP7_75t_SL g823 ( 
.A(n_774),
.Y(n_823)
);

INVx1_ASAP7_75t_L g824 ( 
.A(n_762),
.Y(n_824)
);

OR2x2_ASAP7_75t_L g825 ( 
.A(n_753),
.B(n_255),
.Y(n_825)
);

OAI21x1_ASAP7_75t_L g826 ( 
.A1(n_776),
.A2(n_147),
.B(n_150),
.Y(n_826)
);

INVx2_ASAP7_75t_L g827 ( 
.A(n_783),
.Y(n_827)
);

OAI21x1_ASAP7_75t_L g828 ( 
.A1(n_772),
.A2(n_151),
.B(n_152),
.Y(n_828)
);

INVxp67_ASAP7_75t_L g829 ( 
.A(n_747),
.Y(n_829)
);

INVxp67_ASAP7_75t_L g830 ( 
.A(n_780),
.Y(n_830)
);

INVx2_ASAP7_75t_L g831 ( 
.A(n_783),
.Y(n_831)
);

INVx1_ASAP7_75t_L g832 ( 
.A(n_775),
.Y(n_832)
);

AND2x4_ASAP7_75t_L g833 ( 
.A(n_786),
.B(n_781),
.Y(n_833)
);

INVx2_ASAP7_75t_L g834 ( 
.A(n_786),
.Y(n_834)
);

INVx2_ASAP7_75t_L g835 ( 
.A(n_728),
.Y(n_835)
);

AND2x2_ASAP7_75t_L g836 ( 
.A(n_738),
.B(n_153),
.Y(n_836)
);

INVx2_ASAP7_75t_L g837 ( 
.A(n_728),
.Y(n_837)
);

AND2x4_ASAP7_75t_L g838 ( 
.A(n_790),
.B(n_763),
.Y(n_838)
);

INVx2_ASAP7_75t_SL g839 ( 
.A(n_815),
.Y(n_839)
);

AND2x4_ASAP7_75t_L g840 ( 
.A(n_790),
.B(n_763),
.Y(n_840)
);

OAI22xp5_ASAP7_75t_L g841 ( 
.A1(n_823),
.A2(n_736),
.B1(n_777),
.B2(n_725),
.Y(n_841)
);

INVx1_ASAP7_75t_L g842 ( 
.A(n_792),
.Y(n_842)
);

INVx1_ASAP7_75t_L g843 ( 
.A(n_792),
.Y(n_843)
);

INVx1_ASAP7_75t_L g844 ( 
.A(n_793),
.Y(n_844)
);

INVx2_ASAP7_75t_L g845 ( 
.A(n_789),
.Y(n_845)
);

AND2x4_ASAP7_75t_L g846 ( 
.A(n_789),
.B(n_748),
.Y(n_846)
);

INVx2_ASAP7_75t_L g847 ( 
.A(n_791),
.Y(n_847)
);

HB1xp67_ASAP7_75t_L g848 ( 
.A(n_816),
.Y(n_848)
);

AND2x2_ASAP7_75t_L g849 ( 
.A(n_791),
.B(n_731),
.Y(n_849)
);

AND2x2_ASAP7_75t_L g850 ( 
.A(n_793),
.B(n_731),
.Y(n_850)
);

INVx2_ASAP7_75t_L g851 ( 
.A(n_803),
.Y(n_851)
);

OR2x2_ASAP7_75t_L g852 ( 
.A(n_787),
.B(n_746),
.Y(n_852)
);

INVx2_ASAP7_75t_L g853 ( 
.A(n_803),
.Y(n_853)
);

AND2x4_ASAP7_75t_L g854 ( 
.A(n_807),
.B(n_765),
.Y(n_854)
);

INVx1_ASAP7_75t_SL g855 ( 
.A(n_810),
.Y(n_855)
);

BUFx6f_ASAP7_75t_L g856 ( 
.A(n_835),
.Y(n_856)
);

AND2x2_ASAP7_75t_L g857 ( 
.A(n_802),
.B(n_746),
.Y(n_857)
);

AND2x2_ASAP7_75t_L g858 ( 
.A(n_802),
.B(n_764),
.Y(n_858)
);

HB1xp67_ASAP7_75t_L g859 ( 
.A(n_797),
.Y(n_859)
);

INVx4_ASAP7_75t_SL g860 ( 
.A(n_788),
.Y(n_860)
);

AND2x2_ASAP7_75t_L g861 ( 
.A(n_807),
.B(n_764),
.Y(n_861)
);

INVx1_ASAP7_75t_L g862 ( 
.A(n_808),
.Y(n_862)
);

INVx2_ASAP7_75t_L g863 ( 
.A(n_794),
.Y(n_863)
);

AO31x2_ASAP7_75t_L g864 ( 
.A1(n_814),
.A2(n_732),
.A3(n_773),
.B(n_771),
.Y(n_864)
);

OA21x2_ASAP7_75t_L g865 ( 
.A1(n_814),
.A2(n_772),
.B(n_771),
.Y(n_865)
);

OR2x2_ASAP7_75t_L g866 ( 
.A(n_832),
.B(n_751),
.Y(n_866)
);

INVx1_ASAP7_75t_L g867 ( 
.A(n_794),
.Y(n_867)
);

INVx1_ASAP7_75t_L g868 ( 
.A(n_795),
.Y(n_868)
);

HB1xp67_ASAP7_75t_L g869 ( 
.A(n_830),
.Y(n_869)
);

INVx1_ASAP7_75t_L g870 ( 
.A(n_795),
.Y(n_870)
);

NOR4xp25_ASAP7_75t_L g871 ( 
.A(n_832),
.B(n_777),
.C(n_785),
.D(n_778),
.Y(n_871)
);

AND2x2_ASAP7_75t_L g872 ( 
.A(n_805),
.B(n_757),
.Y(n_872)
);

BUFx2_ASAP7_75t_L g873 ( 
.A(n_799),
.Y(n_873)
);

AND2x2_ASAP7_75t_L g874 ( 
.A(n_805),
.B(n_751),
.Y(n_874)
);

INVx2_ASAP7_75t_L g875 ( 
.A(n_799),
.Y(n_875)
);

INVx2_ASAP7_75t_L g876 ( 
.A(n_800),
.Y(n_876)
);

NAND2xp5_ASAP7_75t_L g877 ( 
.A(n_811),
.B(n_760),
.Y(n_877)
);

INVx2_ASAP7_75t_L g878 ( 
.A(n_800),
.Y(n_878)
);

AND2x4_ASAP7_75t_L g879 ( 
.A(n_834),
.B(n_782),
.Y(n_879)
);

BUFx2_ASAP7_75t_L g880 ( 
.A(n_833),
.Y(n_880)
);

AND2x2_ASAP7_75t_L g881 ( 
.A(n_788),
.B(n_782),
.Y(n_881)
);

AND2x2_ASAP7_75t_L g882 ( 
.A(n_827),
.B(n_782),
.Y(n_882)
);

INVx1_ASAP7_75t_L g883 ( 
.A(n_824),
.Y(n_883)
);

AND2x2_ASAP7_75t_L g884 ( 
.A(n_827),
.B(n_754),
.Y(n_884)
);

OR2x2_ASAP7_75t_L g885 ( 
.A(n_824),
.B(n_754),
.Y(n_885)
);

OR2x2_ASAP7_75t_L g886 ( 
.A(n_831),
.B(n_154),
.Y(n_886)
);

OR2x2_ASAP7_75t_L g887 ( 
.A(n_831),
.B(n_821),
.Y(n_887)
);

AO31x2_ASAP7_75t_L g888 ( 
.A1(n_812),
.A2(n_735),
.A3(n_728),
.B(n_162),
.Y(n_888)
);

NAND2xp5_ASAP7_75t_L g889 ( 
.A(n_813),
.B(n_735),
.Y(n_889)
);

NAND2xp5_ASAP7_75t_L g890 ( 
.A(n_821),
.B(n_809),
.Y(n_890)
);

AND2x4_ASAP7_75t_L g891 ( 
.A(n_834),
.B(n_735),
.Y(n_891)
);

AOI221xp5_ASAP7_75t_L g892 ( 
.A1(n_871),
.A2(n_829),
.B1(n_833),
.B2(n_825),
.C(n_818),
.Y(n_892)
);

OAI221xp5_ASAP7_75t_L g893 ( 
.A1(n_841),
.A2(n_877),
.B1(n_855),
.B2(n_889),
.C(n_825),
.Y(n_893)
);

AOI22xp33_ASAP7_75t_L g894 ( 
.A1(n_852),
.A2(n_801),
.B1(n_798),
.B2(n_769),
.Y(n_894)
);

AND2x2_ASAP7_75t_L g895 ( 
.A(n_857),
.B(n_801),
.Y(n_895)
);

NAND2xp5_ASAP7_75t_L g896 ( 
.A(n_848),
.B(n_818),
.Y(n_896)
);

NAND3xp33_ASAP7_75t_L g897 ( 
.A(n_852),
.B(n_801),
.C(n_836),
.Y(n_897)
);

AOI22xp33_ASAP7_75t_SL g898 ( 
.A1(n_872),
.A2(n_801),
.B1(n_826),
.B2(n_828),
.Y(n_898)
);

NAND2xp5_ASAP7_75t_L g899 ( 
.A(n_869),
.B(n_819),
.Y(n_899)
);

NAND2xp5_ASAP7_75t_SL g900 ( 
.A(n_860),
.B(n_833),
.Y(n_900)
);

NAND3xp33_ASAP7_75t_L g901 ( 
.A(n_866),
.B(n_836),
.C(n_837),
.Y(n_901)
);

OAI22xp5_ASAP7_75t_L g902 ( 
.A1(n_866),
.A2(n_796),
.B1(n_837),
.B2(n_835),
.Y(n_902)
);

NAND3xp33_ASAP7_75t_L g903 ( 
.A(n_886),
.B(n_806),
.C(n_804),
.Y(n_903)
);

NAND2xp5_ASAP7_75t_L g904 ( 
.A(n_859),
.B(n_819),
.Y(n_904)
);

INVx1_ASAP7_75t_L g905 ( 
.A(n_842),
.Y(n_905)
);

INVx1_ASAP7_75t_L g906 ( 
.A(n_843),
.Y(n_906)
);

NAND2xp5_ASAP7_75t_L g907 ( 
.A(n_839),
.B(n_890),
.Y(n_907)
);

AOI22xp5_ASAP7_75t_L g908 ( 
.A1(n_872),
.A2(n_804),
.B1(n_806),
.B2(n_798),
.Y(n_908)
);

NAND2xp5_ASAP7_75t_L g909 ( 
.A(n_839),
.B(n_820),
.Y(n_909)
);

AND2x2_ASAP7_75t_SL g910 ( 
.A(n_858),
.B(n_804),
.Y(n_910)
);

NAND2xp5_ASAP7_75t_L g911 ( 
.A(n_862),
.B(n_820),
.Y(n_911)
);

AND2x2_ASAP7_75t_L g912 ( 
.A(n_874),
.B(n_880),
.Y(n_912)
);

OAI21xp5_ASAP7_75t_SL g913 ( 
.A1(n_850),
.A2(n_858),
.B(n_796),
.Y(n_913)
);

AND2x2_ASAP7_75t_L g914 ( 
.A(n_857),
.B(n_812),
.Y(n_914)
);

NAND2xp5_ASAP7_75t_L g915 ( 
.A(n_846),
.B(n_817),
.Y(n_915)
);

AOI21xp5_ASAP7_75t_SL g916 ( 
.A1(n_886),
.A2(n_796),
.B(n_806),
.Y(n_916)
);

OAI221xp5_ASAP7_75t_SL g917 ( 
.A1(n_850),
.A2(n_817),
.B1(n_798),
.B2(n_769),
.C(n_826),
.Y(n_917)
);

OA21x2_ASAP7_75t_L g918 ( 
.A1(n_844),
.A2(n_828),
.B(n_157),
.Y(n_918)
);

NAND2xp5_ASAP7_75t_L g919 ( 
.A(n_846),
.B(n_822),
.Y(n_919)
);

NAND3xp33_ASAP7_75t_L g920 ( 
.A(n_885),
.B(n_822),
.C(n_768),
.Y(n_920)
);

AOI22xp33_ASAP7_75t_L g921 ( 
.A1(n_849),
.A2(n_822),
.B1(n_755),
.B2(n_768),
.Y(n_921)
);

AND2x2_ASAP7_75t_L g922 ( 
.A(n_860),
.B(n_156),
.Y(n_922)
);

AND2x2_ASAP7_75t_L g923 ( 
.A(n_860),
.B(n_163),
.Y(n_923)
);

AND2x2_ASAP7_75t_L g924 ( 
.A(n_874),
.B(n_881),
.Y(n_924)
);

NAND2xp5_ASAP7_75t_L g925 ( 
.A(n_846),
.B(n_854),
.Y(n_925)
);

AND2x2_ASAP7_75t_L g926 ( 
.A(n_881),
.B(n_727),
.Y(n_926)
);

OR2x2_ASAP7_75t_L g927 ( 
.A(n_895),
.B(n_873),
.Y(n_927)
);

INVx1_ASAP7_75t_L g928 ( 
.A(n_905),
.Y(n_928)
);

AND2x2_ASAP7_75t_L g929 ( 
.A(n_912),
.B(n_860),
.Y(n_929)
);

INVx2_ASAP7_75t_SL g930 ( 
.A(n_919),
.Y(n_930)
);

NAND2xp5_ASAP7_75t_L g931 ( 
.A(n_907),
.B(n_861),
.Y(n_931)
);

INVx1_ASAP7_75t_L g932 ( 
.A(n_906),
.Y(n_932)
);

NAND2xp5_ASAP7_75t_L g933 ( 
.A(n_899),
.B(n_861),
.Y(n_933)
);

OR2x2_ASAP7_75t_L g934 ( 
.A(n_925),
.B(n_887),
.Y(n_934)
);

INVx2_ASAP7_75t_L g935 ( 
.A(n_914),
.Y(n_935)
);

NOR2xp33_ASAP7_75t_L g936 ( 
.A(n_893),
.B(n_856),
.Y(n_936)
);

INVx1_ASAP7_75t_L g937 ( 
.A(n_909),
.Y(n_937)
);

AND2x2_ASAP7_75t_L g938 ( 
.A(n_924),
.B(n_873),
.Y(n_938)
);

AND2x4_ASAP7_75t_L g939 ( 
.A(n_900),
.B(n_914),
.Y(n_939)
);

INVx1_ASAP7_75t_L g940 ( 
.A(n_911),
.Y(n_940)
);

AND2x2_ASAP7_75t_L g941 ( 
.A(n_895),
.B(n_864),
.Y(n_941)
);

AND2x2_ASAP7_75t_L g942 ( 
.A(n_913),
.B(n_864),
.Y(n_942)
);

INVx3_ASAP7_75t_L g943 ( 
.A(n_918),
.Y(n_943)
);

HB1xp67_ASAP7_75t_L g944 ( 
.A(n_915),
.Y(n_944)
);

INVx2_ASAP7_75t_L g945 ( 
.A(n_896),
.Y(n_945)
);

NAND2xp5_ASAP7_75t_L g946 ( 
.A(n_904),
.B(n_849),
.Y(n_946)
);

OR2x2_ASAP7_75t_L g947 ( 
.A(n_897),
.B(n_887),
.Y(n_947)
);

AND2x2_ASAP7_75t_L g948 ( 
.A(n_910),
.B(n_864),
.Y(n_948)
);

INVx1_ASAP7_75t_L g949 ( 
.A(n_902),
.Y(n_949)
);

OR2x2_ASAP7_75t_L g950 ( 
.A(n_894),
.B(n_864),
.Y(n_950)
);

INVx1_ASAP7_75t_L g951 ( 
.A(n_900),
.Y(n_951)
);

AND2x4_ASAP7_75t_SL g952 ( 
.A(n_922),
.B(n_891),
.Y(n_952)
);

NAND2xp5_ASAP7_75t_L g953 ( 
.A(n_949),
.B(n_944),
.Y(n_953)
);

AND2x2_ASAP7_75t_L g954 ( 
.A(n_939),
.B(n_894),
.Y(n_954)
);

INVx2_ASAP7_75t_L g955 ( 
.A(n_943),
.Y(n_955)
);

AND2x2_ASAP7_75t_L g956 ( 
.A(n_939),
.B(n_910),
.Y(n_956)
);

OR2x2_ASAP7_75t_L g957 ( 
.A(n_947),
.B(n_934),
.Y(n_957)
);

AND2x2_ASAP7_75t_L g958 ( 
.A(n_929),
.B(n_939),
.Y(n_958)
);

NAND2xp33_ASAP7_75t_L g959 ( 
.A(n_950),
.B(n_922),
.Y(n_959)
);

INVx2_ASAP7_75t_L g960 ( 
.A(n_943),
.Y(n_960)
);

OA211x2_ASAP7_75t_L g961 ( 
.A1(n_936),
.A2(n_921),
.B(n_892),
.C(n_920),
.Y(n_961)
);

NAND2xp5_ASAP7_75t_L g962 ( 
.A(n_937),
.B(n_901),
.Y(n_962)
);

INVx1_ASAP7_75t_SL g963 ( 
.A(n_952),
.Y(n_963)
);

INVx2_ASAP7_75t_L g964 ( 
.A(n_943),
.Y(n_964)
);

AND2x2_ASAP7_75t_L g965 ( 
.A(n_929),
.B(n_926),
.Y(n_965)
);

INVx1_ASAP7_75t_L g966 ( 
.A(n_928),
.Y(n_966)
);

INVx1_ASAP7_75t_L g967 ( 
.A(n_932),
.Y(n_967)
);

AND2x2_ASAP7_75t_L g968 ( 
.A(n_958),
.B(n_930),
.Y(n_968)
);

OAI21xp5_ASAP7_75t_SL g969 ( 
.A1(n_954),
.A2(n_921),
.B(n_950),
.Y(n_969)
);

NOR2xp33_ASAP7_75t_L g970 ( 
.A(n_962),
.B(n_936),
.Y(n_970)
);

INVx1_ASAP7_75t_L g971 ( 
.A(n_966),
.Y(n_971)
);

INVx3_ASAP7_75t_L g972 ( 
.A(n_955),
.Y(n_972)
);

AND2x2_ASAP7_75t_L g973 ( 
.A(n_956),
.B(n_930),
.Y(n_973)
);

AND2x2_ASAP7_75t_L g974 ( 
.A(n_956),
.B(n_942),
.Y(n_974)
);

INVx1_ASAP7_75t_L g975 ( 
.A(n_967),
.Y(n_975)
);

INVx1_ASAP7_75t_L g976 ( 
.A(n_953),
.Y(n_976)
);

INVx2_ASAP7_75t_SL g977 ( 
.A(n_955),
.Y(n_977)
);

INVx1_ASAP7_75t_L g978 ( 
.A(n_957),
.Y(n_978)
);

AND2x2_ASAP7_75t_L g979 ( 
.A(n_954),
.B(n_963),
.Y(n_979)
);

AND2x2_ASAP7_75t_L g980 ( 
.A(n_979),
.B(n_965),
.Y(n_980)
);

INVx1_ASAP7_75t_SL g981 ( 
.A(n_979),
.Y(n_981)
);

INVx1_ASAP7_75t_L g982 ( 
.A(n_971),
.Y(n_982)
);

INVx1_ASAP7_75t_SL g983 ( 
.A(n_968),
.Y(n_983)
);

OR2x2_ASAP7_75t_L g984 ( 
.A(n_978),
.B(n_946),
.Y(n_984)
);

INVx4_ASAP7_75t_L g985 ( 
.A(n_972),
.Y(n_985)
);

BUFx2_ASAP7_75t_L g986 ( 
.A(n_973),
.Y(n_986)
);

OR2x2_ASAP7_75t_L g987 ( 
.A(n_976),
.B(n_931),
.Y(n_987)
);

OR2x2_ASAP7_75t_L g988 ( 
.A(n_981),
.B(n_969),
.Y(n_988)
);

AOI211xp5_ASAP7_75t_L g989 ( 
.A1(n_982),
.A2(n_970),
.B(n_959),
.C(n_961),
.Y(n_989)
);

NAND2xp5_ASAP7_75t_L g990 ( 
.A(n_980),
.B(n_970),
.Y(n_990)
);

HB1xp67_ASAP7_75t_L g991 ( 
.A(n_986),
.Y(n_991)
);

INVx1_ASAP7_75t_L g992 ( 
.A(n_984),
.Y(n_992)
);

OR2x2_ASAP7_75t_L g993 ( 
.A(n_988),
.B(n_983),
.Y(n_993)
);

NOR2xp33_ASAP7_75t_L g994 ( 
.A(n_990),
.B(n_987),
.Y(n_994)
);

NAND2xp5_ASAP7_75t_SL g995 ( 
.A(n_989),
.B(n_991),
.Y(n_995)
);

NAND2xp5_ASAP7_75t_L g996 ( 
.A(n_992),
.B(n_974),
.Y(n_996)
);

HB1xp67_ASAP7_75t_L g997 ( 
.A(n_991),
.Y(n_997)
);

AOI221xp5_ASAP7_75t_L g998 ( 
.A1(n_995),
.A2(n_959),
.B1(n_985),
.B2(n_975),
.C(n_974),
.Y(n_998)
);

OAI221xp5_ASAP7_75t_L g999 ( 
.A1(n_993),
.A2(n_985),
.B1(n_977),
.B2(n_972),
.C(n_964),
.Y(n_999)
);

XOR2xp5_ASAP7_75t_L g1000 ( 
.A(n_997),
.B(n_908),
.Y(n_1000)
);

AOI221xp5_ASAP7_75t_L g1001 ( 
.A1(n_994),
.A2(n_977),
.B1(n_972),
.B2(n_942),
.C(n_960),
.Y(n_1001)
);

AOI221xp5_ASAP7_75t_L g1002 ( 
.A1(n_996),
.A2(n_964),
.B1(n_960),
.B2(n_917),
.C(n_948),
.Y(n_1002)
);

NOR2xp33_ASAP7_75t_SL g1003 ( 
.A(n_997),
.B(n_923),
.Y(n_1003)
);

HB1xp67_ASAP7_75t_L g1004 ( 
.A(n_997),
.Y(n_1004)
);

NOR4xp25_ASAP7_75t_L g1005 ( 
.A(n_999),
.B(n_951),
.C(n_923),
.D(n_948),
.Y(n_1005)
);

NAND3xp33_ASAP7_75t_L g1006 ( 
.A(n_1004),
.B(n_898),
.C(n_918),
.Y(n_1006)
);

NAND2xp5_ASAP7_75t_L g1007 ( 
.A(n_998),
.B(n_940),
.Y(n_1007)
);

OR2x2_ASAP7_75t_L g1008 ( 
.A(n_1000),
.B(n_945),
.Y(n_1008)
);

NAND2xp5_ASAP7_75t_SL g1009 ( 
.A(n_1003),
.B(n_952),
.Y(n_1009)
);

NOR3xp33_ASAP7_75t_L g1010 ( 
.A(n_1001),
.B(n_1002),
.C(n_903),
.Y(n_1010)
);

NAND4xp25_ASAP7_75t_L g1011 ( 
.A(n_1010),
.B(n_916),
.C(n_941),
.D(n_933),
.Y(n_1011)
);

NAND4xp75_ASAP7_75t_L g1012 ( 
.A(n_1009),
.B(n_941),
.C(n_918),
.D(n_938),
.Y(n_1012)
);

NAND2xp5_ASAP7_75t_L g1013 ( 
.A(n_1005),
.B(n_945),
.Y(n_1013)
);

NOR2xp67_ASAP7_75t_L g1014 ( 
.A(n_1008),
.B(n_164),
.Y(n_1014)
);

NAND3xp33_ASAP7_75t_SL g1015 ( 
.A(n_1007),
.B(n_927),
.C(n_938),
.Y(n_1015)
);

OAI211xp5_ASAP7_75t_SL g1016 ( 
.A1(n_1006),
.A2(n_927),
.B(n_885),
.C(n_935),
.Y(n_1016)
);

NOR2x1_ASAP7_75t_L g1017 ( 
.A(n_1009),
.B(n_935),
.Y(n_1017)
);

NAND4xp25_ASAP7_75t_L g1018 ( 
.A(n_1010),
.B(n_882),
.C(n_891),
.D(n_838),
.Y(n_1018)
);

NOR2x2_ASAP7_75t_L g1019 ( 
.A(n_1012),
.B(n_851),
.Y(n_1019)
);

BUFx2_ASAP7_75t_L g1020 ( 
.A(n_1017),
.Y(n_1020)
);

INVx1_ASAP7_75t_L g1021 ( 
.A(n_1014),
.Y(n_1021)
);

AND2x2_ASAP7_75t_L g1022 ( 
.A(n_1013),
.B(n_856),
.Y(n_1022)
);

INVxp67_ASAP7_75t_SL g1023 ( 
.A(n_1018),
.Y(n_1023)
);

INVx1_ASAP7_75t_L g1024 ( 
.A(n_1015),
.Y(n_1024)
);

NAND2xp5_ASAP7_75t_L g1025 ( 
.A(n_1011),
.B(n_856),
.Y(n_1025)
);

INVx1_ASAP7_75t_L g1026 ( 
.A(n_1016),
.Y(n_1026)
);

INVx1_ASAP7_75t_L g1027 ( 
.A(n_1014),
.Y(n_1027)
);

INVx1_ASAP7_75t_L g1028 ( 
.A(n_1014),
.Y(n_1028)
);

INVx1_ASAP7_75t_L g1029 ( 
.A(n_1014),
.Y(n_1029)
);

INVx1_ASAP7_75t_L g1030 ( 
.A(n_1014),
.Y(n_1030)
);

OAI22xp33_ASAP7_75t_L g1031 ( 
.A1(n_1011),
.A2(n_856),
.B1(n_883),
.B2(n_870),
.Y(n_1031)
);

INVx1_ASAP7_75t_L g1032 ( 
.A(n_1014),
.Y(n_1032)
);

NAND2xp5_ASAP7_75t_L g1033 ( 
.A(n_1014),
.B(n_867),
.Y(n_1033)
);

NAND2xp5_ASAP7_75t_SL g1034 ( 
.A(n_1014),
.B(n_838),
.Y(n_1034)
);

INVx1_ASAP7_75t_L g1035 ( 
.A(n_1020),
.Y(n_1035)
);

AND2x2_ASAP7_75t_L g1036 ( 
.A(n_1024),
.B(n_882),
.Y(n_1036)
);

OAI221xp5_ASAP7_75t_L g1037 ( 
.A1(n_1023),
.A2(n_1026),
.B1(n_1021),
.B2(n_1032),
.C(n_1030),
.Y(n_1037)
);

AOI221xp5_ASAP7_75t_L g1038 ( 
.A1(n_1031),
.A2(n_1027),
.B1(n_1029),
.B2(n_1028),
.C(n_1022),
.Y(n_1038)
);

NAND4xp25_ASAP7_75t_L g1039 ( 
.A(n_1025),
.B(n_891),
.C(n_838),
.D(n_840),
.Y(n_1039)
);

NAND4xp25_ASAP7_75t_L g1040 ( 
.A(n_1033),
.B(n_840),
.C(n_879),
.D(n_884),
.Y(n_1040)
);

OR2x2_ASAP7_75t_L g1041 ( 
.A(n_1033),
.B(n_864),
.Y(n_1041)
);

BUFx2_ASAP7_75t_L g1042 ( 
.A(n_1019),
.Y(n_1042)
);

NAND2xp5_ASAP7_75t_SL g1043 ( 
.A(n_1034),
.B(n_840),
.Y(n_1043)
);

INVx2_ASAP7_75t_L g1044 ( 
.A(n_1020),
.Y(n_1044)
);

AND2x2_ASAP7_75t_L g1045 ( 
.A(n_1024),
.B(n_879),
.Y(n_1045)
);

INVx2_ASAP7_75t_L g1046 ( 
.A(n_1020),
.Y(n_1046)
);

NOR3xp33_ASAP7_75t_L g1047 ( 
.A(n_1021),
.B(n_884),
.C(n_879),
.Y(n_1047)
);

NAND2xp5_ASAP7_75t_L g1048 ( 
.A(n_1020),
.B(n_868),
.Y(n_1048)
);

NAND5xp2_ASAP7_75t_L g1049 ( 
.A(n_1024),
.B(n_888),
.C(n_166),
.D(n_167),
.E(n_168),
.Y(n_1049)
);

NOR2xp33_ASAP7_75t_R g1050 ( 
.A(n_1021),
.B(n_165),
.Y(n_1050)
);

NOR2xp67_ASAP7_75t_L g1051 ( 
.A(n_1021),
.B(n_169),
.Y(n_1051)
);

AND2x2_ASAP7_75t_L g1052 ( 
.A(n_1024),
.B(n_854),
.Y(n_1052)
);

OR2x2_ASAP7_75t_L g1053 ( 
.A(n_1044),
.B(n_851),
.Y(n_1053)
);

INVx1_ASAP7_75t_L g1054 ( 
.A(n_1042),
.Y(n_1054)
);

INVx1_ASAP7_75t_L g1055 ( 
.A(n_1035),
.Y(n_1055)
);

AND2x4_ASAP7_75t_L g1056 ( 
.A(n_1046),
.B(n_854),
.Y(n_1056)
);

NOR2xp67_ASAP7_75t_L g1057 ( 
.A(n_1049),
.B(n_170),
.Y(n_1057)
);

NAND4xp75_ASAP7_75t_L g1058 ( 
.A(n_1038),
.B(n_865),
.C(n_174),
.D(n_175),
.Y(n_1058)
);

NOR2x1p5_ASAP7_75t_L g1059 ( 
.A(n_1045),
.B(n_853),
.Y(n_1059)
);

INVx1_ASAP7_75t_L g1060 ( 
.A(n_1036),
.Y(n_1060)
);

INVx1_ASAP7_75t_L g1061 ( 
.A(n_1051),
.Y(n_1061)
);

NAND4xp25_ASAP7_75t_L g1062 ( 
.A(n_1037),
.B(n_853),
.C(n_876),
.D(n_875),
.Y(n_1062)
);

NAND4xp75_ASAP7_75t_L g1063 ( 
.A(n_1051),
.B(n_865),
.C(n_192),
.D(n_194),
.Y(n_1063)
);

OAI22xp5_ASAP7_75t_L g1064 ( 
.A1(n_1054),
.A2(n_1043),
.B1(n_1052),
.B2(n_1048),
.Y(n_1064)
);

INVx1_ASAP7_75t_SL g1065 ( 
.A(n_1061),
.Y(n_1065)
);

INVx1_ASAP7_75t_L g1066 ( 
.A(n_1055),
.Y(n_1066)
);

NAND4xp25_ASAP7_75t_L g1067 ( 
.A(n_1057),
.B(n_1047),
.C(n_1040),
.D(n_1041),
.Y(n_1067)
);

AOI22x1_ASAP7_75t_L g1068 ( 
.A1(n_1060),
.A2(n_1050),
.B1(n_1039),
.B2(n_199),
.Y(n_1068)
);

INVx1_ASAP7_75t_L g1069 ( 
.A(n_1053),
.Y(n_1069)
);

OAI221xp5_ASAP7_75t_L g1070 ( 
.A1(n_1065),
.A2(n_1062),
.B1(n_1058),
.B2(n_1059),
.C(n_1063),
.Y(n_1070)
);

NAND3xp33_ASAP7_75t_L g1071 ( 
.A(n_1066),
.B(n_1056),
.C(n_878),
.Y(n_1071)
);

NAND3xp33_ASAP7_75t_SL g1072 ( 
.A(n_1069),
.B(n_171),
.C(n_198),
.Y(n_1072)
);

NAND3xp33_ASAP7_75t_SL g1073 ( 
.A(n_1064),
.B(n_1068),
.C(n_1067),
.Y(n_1073)
);

AOI221xp5_ASAP7_75t_L g1074 ( 
.A1(n_1073),
.A2(n_878),
.B1(n_876),
.B2(n_875),
.C(n_863),
.Y(n_1074)
);

OAI22xp5_ASAP7_75t_L g1075 ( 
.A1(n_1070),
.A2(n_1071),
.B1(n_1072),
.B2(n_863),
.Y(n_1075)
);

AOI21x1_ASAP7_75t_L g1076 ( 
.A1(n_1075),
.A2(n_201),
.B(n_202),
.Y(n_1076)
);

AOI21xp5_ASAP7_75t_L g1077 ( 
.A1(n_1074),
.A2(n_203),
.B(n_204),
.Y(n_1077)
);

OAI22xp5_ASAP7_75t_SL g1078 ( 
.A1(n_1075),
.A2(n_888),
.B1(n_206),
.B2(n_208),
.Y(n_1078)
);

NAND2x1p5_ASAP7_75t_L g1079 ( 
.A(n_1076),
.B(n_205),
.Y(n_1079)
);

OAI21xp33_ASAP7_75t_L g1080 ( 
.A1(n_1077),
.A2(n_847),
.B(n_845),
.Y(n_1080)
);

AOI21xp5_ASAP7_75t_L g1081 ( 
.A1(n_1079),
.A2(n_1078),
.B(n_210),
.Y(n_1081)
);

INVx3_ASAP7_75t_L g1082 ( 
.A(n_1080),
.Y(n_1082)
);

AOI22xp5_ASAP7_75t_SL g1083 ( 
.A1(n_1081),
.A2(n_209),
.B1(n_211),
.B2(n_212),
.Y(n_1083)
);

AOI221xp5_ASAP7_75t_L g1084 ( 
.A1(n_1083),
.A2(n_1082),
.B1(n_215),
.B2(n_216),
.C(n_217),
.Y(n_1084)
);

AOI211xp5_ASAP7_75t_L g1085 ( 
.A1(n_1084),
.A2(n_214),
.B(n_221),
.C(n_222),
.Y(n_1085)
);


endmodule