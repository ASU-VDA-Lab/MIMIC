module real_aes_6299_n_104 (n_17, n_28, n_76, n_56, n_34, n_98, n_90, n_82, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_83, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_91, n_100, n_43, n_103, n_96, n_54, n_35, n_42, n_99, n_15, n_9, n_23, n_72, n_95, n_44, n_102, n_7, n_4, n_80, n_6, n_12, n_68, n_79, n_69, n_46, n_59, n_25, n_73, n_77, n_81, n_48, n_37, n_97, n_70, n_50, n_89, n_26, n_86, n_93, n_13, n_24, n_2, n_55, n_62, n_84, n_67, n_92, n_33, n_88, n_14, n_11, n_85, n_16, n_94, n_39, n_5, n_45, n_60, n_38, n_87, n_0, n_78, n_101, n_63, n_1, n_53, n_36, n_104);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_98;
input n_90;
input n_82;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_83;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_91;
input n_100;
input n_43;
input n_103;
input n_96;
input n_54;
input n_35;
input n_42;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_95;
input n_44;
input n_102;
input n_7;
input n_4;
input n_80;
input n_6;
input n_12;
input n_68;
input n_79;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_81;
input n_48;
input n_37;
input n_97;
input n_70;
input n_50;
input n_89;
input n_26;
input n_86;
input n_93;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_84;
input n_67;
input n_92;
input n_33;
input n_88;
input n_14;
input n_11;
input n_85;
input n_16;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_87;
input n_0;
input n_78;
input n_101;
input n_63;
input n_1;
input n_53;
input n_36;
output n_104;
wire n_480;
wire n_113;
wire n_476;
wire n_758;
wire n_599;
wire n_187;
wire n_436;
wire n_684;
wire n_257;
wire n_390;
wire n_185;
wire n_285;
wire n_624;
wire n_618;
wire n_522;
wire n_485;
wire n_222;
wire n_750;
wire n_631;
wire n_503;
wire n_287;
wire n_357;
wire n_635;
wire n_386;
wire n_673;
wire n_518;
wire n_254;
wire n_207;
wire n_665;
wire n_667;
wire n_580;
wire n_577;
wire n_469;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_759;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_718;
wire n_318;
wire n_355;
wire n_239;
wire n_669;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_761;
wire n_742;
wire n_112;
wire n_319;
wire n_364;
wire n_555;
wire n_421;
wire n_329;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_242;
wire n_169;
wire n_571;
wire n_549;
wire n_376;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_752;
wire n_448;
wire n_556;
wire n_341;
wire n_545;
wire n_593;
wire n_232;
wire n_460;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_537;
wire n_551;
wire n_320;
wire n_666;
wire n_560;
wire n_260;
wire n_660;
wire n_594;
wire n_186;
wire n_138;
wire n_696;
wire n_704;
wire n_379;
wire n_374;
wire n_453;
wire n_647;
wire n_235;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_161;
wire n_763;
wire n_189;
wire n_271;
wire n_489;
wire n_548;
wire n_427;
wire n_678;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_519;
wire n_564;
wire n_638;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_512;
wire n_395;
wire n_332;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_116;
wire n_625;
wire n_462;
wire n_289;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_716;
wire n_213;
wire n_356;
wire n_478;
wire n_584;
wire n_408;
wire n_553;
wire n_184;
wire n_578;
wire n_528;
wire n_372;
wire n_202;
wire n_495;
wire n_370;
wire n_384;
wire n_744;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_467;
wire n_327;
wire n_106;
wire n_466;
wire n_559;
wire n_636;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_726;
wire n_517;
wire n_683;
wire n_174;
wire n_570;
wire n_675;
wire n_530;
wire n_535;
wire n_732;
wire n_211;
wire n_281;
wire n_496;
wire n_693;
wire n_173;
wire n_468;
wire n_234;
wire n_755;
wire n_284;
wire n_153;
wire n_316;
wire n_532;
wire n_746;
wire n_656;
wire n_178;
wire n_409;
wire n_748;
wire n_523;
wire n_298;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_649;
wire n_651;
wire n_297;
wire n_383;
wire n_529;
wire n_119;
wire n_504;
wire n_310;
wire n_455;
wire n_725;
wire n_164;
wire n_671;
wire n_231;
wire n_547;
wire n_659;
wire n_634;
wire n_682;
wire n_454;
wire n_122;
wire n_565;
wire n_443;
wire n_760;
wire n_608;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_267;
wire n_218;
wire n_737;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_722;
wire n_745;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_331;
wire n_449;
wire n_182;
wire n_417;
wire n_754;
wire n_363;
wire n_607;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_142;
wire n_561;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_655;
wire n_654;
wire n_527;
wire n_505;
wire n_434;
wire n_502;
wire n_600;
wire n_731;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_617;
wire n_552;
wire n_402;
wire n_602;
wire n_733;
wire n_171;
wire n_658;
wire n_676;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_146;
wire n_432;
wire n_255;
wire n_226;
wire n_286;
wire n_416;
wire n_410;
wire n_120;
wire n_751;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_695;
wire n_685;
wire n_165;
wire n_361;
wire n_632;
wire n_246;
wire n_176;
wire n_412;
wire n_163;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_488;
wire n_501;
wire n_251;
wire n_642;
wire n_613;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_702;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_734;
wire n_110;
wire n_392;
wire n_562;
wire n_150;
wire n_147;
wire n_756;
wire n_288;
wire n_404;
wire n_598;
wire n_728;
wire n_713;
wire n_735;
wire n_334;
wire n_274;
wire n_160;
wire n_569;
wire n_303;
wire n_563;
wire n_188;
wire n_269;
wire n_430;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_193;
wire n_397;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_749;
wire n_663;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_707;
wire n_622;
wire n_470;
wire n_133;
wire n_494;
wire n_711;
wire n_377;
wire n_273;
wire n_723;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_265;
wire n_354;
wire n_720;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_730;
wire n_643;
wire n_747;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_148;
wire n_481;
wire n_498;
wire n_691;
wire n_765;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_233;
wire n_487;
wire n_290;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_155;
wire n_243;
wire n_692;
wire n_544;
wire n_268;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_738;
wire n_701;
wire n_309;
wire n_344;
wire n_229;
wire n_107;
wire n_482;
wire n_520;
wire n_633;
wire n_679;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_262;
wire n_630;
wire n_689;
wire n_715;
wire n_134;
wire n_349;
wire n_336;
wire n_420;
wire n_612;
wire n_195;
wire n_438;
wire n_764;
wire n_300;
wire n_252;
wire n_283;
wire n_314;
wire n_741;
wire n_753;
wire n_249;
wire n_623;
wire n_446;
wire n_721;
wire n_221;
wire n_681;
wire n_456;
wire n_156;
wire n_359;
wire n_717;
wire n_312;
wire n_183;
wire n_266;
wire n_712;
wire n_205;
wire n_433;
wire n_516;
wire n_177;
wire n_335;
wire n_313;
wire n_627;
wire n_739;
wire n_140;
wire n_418;
wire n_521;
wire n_422;
wire n_524;
wire n_219;
wire n_705;
wire n_180;
wire n_212;
wire n_575;
wire n_210;
wire n_325;
wire n_762;
wire n_338;
wire n_479;
wire n_442;
wire n_740;
wire n_371;
wire n_698;
wire n_166;
wire n_541;
wire n_224;
wire n_151;
wire n_546;
wire n_587;
wire n_639;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_724;
wire n_440;
wire n_525;
wire n_674;
wire n_644;
wire n_152;
wire n_198;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_414;
wire n_757;
wire n_123;
wire n_279;
wire n_686;
wire n_543;
wire n_497;
wire n_514;
wire n_507;
wire n_270;
wire n_614;
wire n_305;
wire n_586;
wire n_450;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_465;
wire n_473;
wire n_719;
wire n_566;
wire n_474;
wire n_170;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_168;
wire n_175;
wire n_241;
wire n_687;
wire n_729;
wire n_646;
wire n_650;
wire n_710;
wire n_105;
wire n_743;
wire n_294;
wire n_393;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_307;
wire n_500;
wire n_601;
wire n_661;
wire n_463;
wire n_396;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_143;
wire n_192;
wire n_554;
wire n_475;
wire n_264;
wire n_237;
wire n_668;
A2O1A1Ixp33_ASAP7_75t_SL g256 ( .A1(n_0), .A2(n_257), .B(n_258), .C(n_261), .Y(n_256) );
NAND2xp5_ASAP7_75t_L g262 ( .A(n_1), .B(n_245), .Y(n_262) );
INVx1_ASAP7_75t_L g109 ( .A(n_2), .Y(n_109) );
NAND2xp5_ASAP7_75t_SL g172 ( .A(n_3), .B(n_173), .Y(n_172) );
A2O1A1Ixp33_ASAP7_75t_L g550 ( .A1(n_4), .A2(n_134), .B(n_137), .C(n_551), .Y(n_550) );
AOI21xp5_ASAP7_75t_L g574 ( .A1(n_5), .A2(n_129), .B(n_575), .Y(n_574) );
AOI21xp5_ASAP7_75t_L g238 ( .A1(n_6), .A2(n_129), .B(n_239), .Y(n_238) );
NAND2xp5_ASAP7_75t_L g581 ( .A(n_7), .B(n_245), .Y(n_581) );
AO21x2_ASAP7_75t_L g200 ( .A1(n_8), .A2(n_164), .B(n_201), .Y(n_200) );
AND2x6_ASAP7_75t_L g134 ( .A(n_9), .B(n_135), .Y(n_134) );
A2O1A1Ixp33_ASAP7_75t_L g217 ( .A1(n_10), .A2(n_134), .B(n_137), .C(n_218), .Y(n_217) );
INVx1_ASAP7_75t_L g519 ( .A(n_11), .Y(n_519) );
NAND2xp5_ASAP7_75t_L g107 ( .A(n_12), .B(n_40), .Y(n_107) );
NOR2xp33_ASAP7_75t_L g458 ( .A(n_12), .B(n_40), .Y(n_458) );
AOI22xp5_ASAP7_75t_L g465 ( .A1(n_13), .A2(n_466), .B1(n_467), .B2(n_468), .Y(n_465) );
CKINVDCx20_ASAP7_75t_R g466 ( .A(n_13), .Y(n_466) );
NAND2xp5_ASAP7_75t_SL g553 ( .A(n_14), .B(n_221), .Y(n_553) );
INVx1_ASAP7_75t_L g155 ( .A(n_15), .Y(n_155) );
NAND2xp5_ASAP7_75t_SL g207 ( .A(n_16), .B(n_173), .Y(n_207) );
A2O1A1Ixp33_ASAP7_75t_L g536 ( .A1(n_17), .A2(n_174), .B(n_537), .C(n_539), .Y(n_536) );
NAND2xp5_ASAP7_75t_L g540 ( .A(n_18), .B(n_245), .Y(n_540) );
NAND2xp5_ASAP7_75t_L g510 ( .A(n_19), .B(n_149), .Y(n_510) );
A2O1A1Ixp33_ASAP7_75t_L g136 ( .A1(n_20), .A2(n_137), .B(n_140), .C(n_148), .Y(n_136) );
A2O1A1Ixp33_ASAP7_75t_L g526 ( .A1(n_21), .A2(n_209), .B(n_260), .C(n_527), .Y(n_526) );
NAND2xp5_ASAP7_75t_SL g570 ( .A(n_22), .B(n_221), .Y(n_570) );
AOI22xp5_ASAP7_75t_L g447 ( .A1(n_23), .A2(n_56), .B1(n_448), .B2(n_449), .Y(n_447) );
CKINVDCx20_ASAP7_75t_R g448 ( .A(n_23), .Y(n_448) );
NAND2xp5_ASAP7_75t_SL g492 ( .A(n_24), .B(n_221), .Y(n_492) );
CKINVDCx16_ASAP7_75t_R g566 ( .A(n_25), .Y(n_566) );
INVx1_ASAP7_75t_L g491 ( .A(n_26), .Y(n_491) );
A2O1A1Ixp33_ASAP7_75t_L g203 ( .A1(n_27), .A2(n_137), .B(n_148), .C(n_204), .Y(n_203) );
BUFx6f_ASAP7_75t_L g133 ( .A(n_28), .Y(n_133) );
CKINVDCx20_ASAP7_75t_R g549 ( .A(n_29), .Y(n_549) );
INVx1_ASAP7_75t_L g507 ( .A(n_30), .Y(n_507) );
AOI21xp5_ASAP7_75t_L g253 ( .A1(n_31), .A2(n_129), .B(n_254), .Y(n_253) );
INVx2_ASAP7_75t_L g132 ( .A(n_32), .Y(n_132) );
A2O1A1Ixp33_ASAP7_75t_L g185 ( .A1(n_33), .A2(n_177), .B(n_186), .C(n_188), .Y(n_185) );
CKINVDCx20_ASAP7_75t_R g556 ( .A(n_34), .Y(n_556) );
A2O1A1Ixp33_ASAP7_75t_L g577 ( .A1(n_35), .A2(n_260), .B(n_578), .C(n_580), .Y(n_577) );
INVxp67_ASAP7_75t_L g508 ( .A(n_36), .Y(n_508) );
NAND2xp5_ASAP7_75t_L g205 ( .A(n_37), .B(n_206), .Y(n_205) );
A2O1A1Ixp33_ASAP7_75t_L g489 ( .A1(n_38), .A2(n_137), .B(n_148), .C(n_490), .Y(n_489) );
CKINVDCx14_ASAP7_75t_R g576 ( .A(n_39), .Y(n_576) );
A2O1A1Ixp33_ASAP7_75t_L g516 ( .A1(n_41), .A2(n_261), .B(n_517), .C(n_518), .Y(n_516) );
NAND2xp5_ASAP7_75t_L g127 ( .A(n_42), .B(n_128), .Y(n_127) );
CKINVDCx20_ASAP7_75t_R g223 ( .A(n_43), .Y(n_223) );
NAND2xp5_ASAP7_75t_L g232 ( .A(n_44), .B(n_173), .Y(n_232) );
NAND2xp5_ASAP7_75t_L g202 ( .A(n_45), .B(n_129), .Y(n_202) );
CKINVDCx20_ASAP7_75t_R g494 ( .A(n_46), .Y(n_494) );
CKINVDCx20_ASAP7_75t_R g504 ( .A(n_47), .Y(n_504) );
A2O1A1Ixp33_ASAP7_75t_L g229 ( .A1(n_48), .A2(n_177), .B(n_186), .C(n_230), .Y(n_229) );
NAND2xp5_ASAP7_75t_L g459 ( .A(n_49), .B(n_460), .Y(n_459) );
INVx1_ASAP7_75t_L g259 ( .A(n_50), .Y(n_259) );
OAI22xp5_ASAP7_75t_SL g445 ( .A1(n_51), .A2(n_446), .B1(n_447), .B2(n_450), .Y(n_445) );
CKINVDCx16_ASAP7_75t_R g450 ( .A(n_51), .Y(n_450) );
AOI222xp33_ASAP7_75t_L g463 ( .A1(n_52), .A2(n_464), .B1(n_465), .B2(n_474), .C1(n_754), .C2(n_758), .Y(n_463) );
INVx1_ASAP7_75t_L g231 ( .A(n_53), .Y(n_231) );
INVx1_ASAP7_75t_L g525 ( .A(n_54), .Y(n_525) );
NAND2xp5_ASAP7_75t_L g228 ( .A(n_55), .B(n_129), .Y(n_228) );
CKINVDCx20_ASAP7_75t_R g449 ( .A(n_56), .Y(n_449) );
CKINVDCx20_ASAP7_75t_R g157 ( .A(n_57), .Y(n_157) );
CKINVDCx14_ASAP7_75t_R g515 ( .A(n_58), .Y(n_515) );
INVx1_ASAP7_75t_L g135 ( .A(n_59), .Y(n_135) );
NAND2xp5_ASAP7_75t_L g179 ( .A(n_60), .B(n_129), .Y(n_179) );
NAND2xp5_ASAP7_75t_L g244 ( .A(n_61), .B(n_245), .Y(n_244) );
A2O1A1Ixp33_ASAP7_75t_L g241 ( .A1(n_62), .A2(n_147), .B(n_170), .C(n_242), .Y(n_241) );
INVx1_ASAP7_75t_L g154 ( .A(n_63), .Y(n_154) );
OAI22xp5_ASAP7_75t_L g469 ( .A1(n_64), .A2(n_103), .B1(n_470), .B2(n_471), .Y(n_469) );
CKINVDCx20_ASAP7_75t_R g471 ( .A(n_64), .Y(n_471) );
INVx1_ASAP7_75t_SL g579 ( .A(n_65), .Y(n_579) );
CKINVDCx20_ASAP7_75t_R g115 ( .A(n_66), .Y(n_115) );
NAND2xp5_ASAP7_75t_SL g190 ( .A(n_67), .B(n_173), .Y(n_190) );
NAND2xp5_ASAP7_75t_L g529 ( .A(n_68), .B(n_245), .Y(n_529) );
NAND2xp5_ASAP7_75t_L g219 ( .A(n_69), .B(n_174), .Y(n_219) );
INVx1_ASAP7_75t_L g569 ( .A(n_70), .Y(n_569) );
CKINVDCx16_ASAP7_75t_R g255 ( .A(n_71), .Y(n_255) );
NAND2xp5_ASAP7_75t_L g141 ( .A(n_72), .B(n_142), .Y(n_141) );
A2O1A1Ixp33_ASAP7_75t_L g167 ( .A1(n_73), .A2(n_137), .B(n_168), .C(n_177), .Y(n_167) );
CKINVDCx16_ASAP7_75t_R g240 ( .A(n_74), .Y(n_240) );
INVx1_ASAP7_75t_L g112 ( .A(n_75), .Y(n_112) );
AOI21xp5_ASAP7_75t_L g513 ( .A1(n_76), .A2(n_129), .B(n_514), .Y(n_513) );
CKINVDCx20_ASAP7_75t_R g572 ( .A(n_77), .Y(n_572) );
AOI21xp5_ASAP7_75t_L g533 ( .A1(n_78), .A2(n_129), .B(n_534), .Y(n_533) );
AOI21xp5_ASAP7_75t_L g502 ( .A1(n_79), .A2(n_128), .B(n_503), .Y(n_502) );
CKINVDCx16_ASAP7_75t_R g488 ( .A(n_80), .Y(n_488) );
INVx1_ASAP7_75t_L g535 ( .A(n_81), .Y(n_535) );
NAND2xp5_ASAP7_75t_SL g144 ( .A(n_82), .B(n_145), .Y(n_144) );
CKINVDCx20_ASAP7_75t_R g194 ( .A(n_83), .Y(n_194) );
AOI21xp5_ASAP7_75t_L g523 ( .A1(n_84), .A2(n_129), .B(n_524), .Y(n_523) );
INVx1_ASAP7_75t_L g538 ( .A(n_85), .Y(n_538) );
INVx2_ASAP7_75t_L g152 ( .A(n_86), .Y(n_152) );
INVx1_ASAP7_75t_L g552 ( .A(n_87), .Y(n_552) );
CKINVDCx20_ASAP7_75t_R g181 ( .A(n_88), .Y(n_181) );
NAND2xp5_ASAP7_75t_SL g220 ( .A(n_89), .B(n_221), .Y(n_220) );
NAND3xp33_ASAP7_75t_SL g108 ( .A(n_90), .B(n_109), .C(n_110), .Y(n_108) );
OR2x2_ASAP7_75t_L g455 ( .A(n_90), .B(n_456), .Y(n_455) );
OR2x2_ASAP7_75t_L g477 ( .A(n_90), .B(n_457), .Y(n_477) );
INVx2_ASAP7_75t_L g479 ( .A(n_90), .Y(n_479) );
OAI22xp5_ASAP7_75t_SL g468 ( .A1(n_91), .A2(n_469), .B1(n_472), .B2(n_473), .Y(n_468) );
CKINVDCx20_ASAP7_75t_R g473 ( .A(n_91), .Y(n_473) );
A2O1A1Ixp33_ASAP7_75t_L g567 ( .A1(n_92), .A2(n_137), .B(n_177), .C(n_568), .Y(n_567) );
NAND2xp5_ASAP7_75t_L g184 ( .A(n_93), .B(n_129), .Y(n_184) );
INVx1_ASAP7_75t_L g189 ( .A(n_94), .Y(n_189) );
INVxp67_ASAP7_75t_L g243 ( .A(n_95), .Y(n_243) );
XNOR2xp5_ASAP7_75t_L g117 ( .A(n_96), .B(n_118), .Y(n_117) );
NAND2xp5_ASAP7_75t_L g520 ( .A(n_96), .B(n_164), .Y(n_520) );
AOI22xp5_ASAP7_75t_L g104 ( .A1(n_97), .A2(n_105), .B1(n_113), .B2(n_764), .Y(n_104) );
NAND2xp5_ASAP7_75t_L g111 ( .A(n_98), .B(n_112), .Y(n_111) );
INVx1_ASAP7_75t_L g169 ( .A(n_99), .Y(n_169) );
INVx1_ASAP7_75t_L g215 ( .A(n_100), .Y(n_215) );
INVx2_ASAP7_75t_L g528 ( .A(n_101), .Y(n_528) );
AND2x2_ASAP7_75t_L g233 ( .A(n_102), .B(n_151), .Y(n_233) );
CKINVDCx20_ASAP7_75t_R g470 ( .A(n_103), .Y(n_470) );
INVx1_ASAP7_75t_SL g105 ( .A(n_106), .Y(n_105) );
CKINVDCx12_ASAP7_75t_R g765 ( .A(n_106), .Y(n_765) );
OR2x2_ASAP7_75t_L g106 ( .A(n_107), .B(n_108), .Y(n_106) );
AND2x2_ASAP7_75t_L g457 ( .A(n_109), .B(n_458), .Y(n_457) );
INVx1_ASAP7_75t_SL g110 ( .A(n_111), .Y(n_110) );
OA21x2_ASAP7_75t_L g113 ( .A1(n_114), .A2(n_116), .B(n_462), .Y(n_113) );
INVx1_ASAP7_75t_L g114 ( .A(n_115), .Y(n_114) );
INVx2_ASAP7_75t_L g763 ( .A(n_115), .Y(n_763) );
OAI21xp5_ASAP7_75t_SL g116 ( .A1(n_117), .A2(n_452), .B(n_459), .Y(n_116) );
OAI22xp5_ASAP7_75t_SL g118 ( .A1(n_119), .A2(n_444), .B1(n_445), .B2(n_451), .Y(n_118) );
OAI22xp5_ASAP7_75t_SL g754 ( .A1(n_119), .A2(n_481), .B1(n_755), .B2(n_756), .Y(n_754) );
INVx1_ASAP7_75t_L g119 ( .A(n_120), .Y(n_119) );
BUFx2_ASAP7_75t_L g451 ( .A(n_120), .Y(n_451) );
AND3x1_ASAP7_75t_L g120 ( .A(n_121), .B(n_348), .C(n_405), .Y(n_120) );
NOR3xp33_ASAP7_75t_L g121 ( .A(n_122), .B(n_293), .C(n_329), .Y(n_121) );
OAI211xp5_ASAP7_75t_L g122 ( .A1(n_123), .A2(n_195), .B(n_247), .C(n_280), .Y(n_122) );
NAND2xp5_ASAP7_75t_L g123 ( .A(n_124), .B(n_159), .Y(n_123) );
HB1xp67_ASAP7_75t_L g124 ( .A(n_125), .Y(n_124) );
AND2x4_ASAP7_75t_L g250 ( .A(n_125), .B(n_251), .Y(n_250) );
INVx5_ASAP7_75t_L g279 ( .A(n_125), .Y(n_279) );
AND2x2_ASAP7_75t_L g352 ( .A(n_125), .B(n_268), .Y(n_352) );
AND2x2_ASAP7_75t_L g390 ( .A(n_125), .B(n_296), .Y(n_390) );
AND2x2_ASAP7_75t_L g410 ( .A(n_125), .B(n_252), .Y(n_410) );
OR2x6_ASAP7_75t_L g125 ( .A(n_126), .B(n_156), .Y(n_125) );
AOI21xp5_ASAP7_75t_SL g126 ( .A1(n_127), .A2(n_136), .B(n_149), .Y(n_126) );
BUFx2_ASAP7_75t_L g128 ( .A(n_129), .Y(n_128) );
AND2x4_ASAP7_75t_L g129 ( .A(n_130), .B(n_134), .Y(n_129) );
NAND2x1p5_ASAP7_75t_L g216 ( .A(n_130), .B(n_134), .Y(n_216) );
AND2x2_ASAP7_75t_L g130 ( .A(n_131), .B(n_133), .Y(n_130) );
INVx1_ASAP7_75t_L g147 ( .A(n_131), .Y(n_147) );
INVx1_ASAP7_75t_L g131 ( .A(n_132), .Y(n_131) );
INVx2_ASAP7_75t_L g138 ( .A(n_132), .Y(n_138) );
INVx1_ASAP7_75t_L g210 ( .A(n_132), .Y(n_210) );
INVx1_ASAP7_75t_L g139 ( .A(n_133), .Y(n_139) );
BUFx6f_ASAP7_75t_L g143 ( .A(n_133), .Y(n_143) );
INVx3_ASAP7_75t_L g174 ( .A(n_133), .Y(n_174) );
INVx1_ASAP7_75t_L g206 ( .A(n_133), .Y(n_206) );
BUFx6f_ASAP7_75t_L g221 ( .A(n_133), .Y(n_221) );
BUFx3_ASAP7_75t_L g148 ( .A(n_134), .Y(n_148) );
INVx4_ASAP7_75t_SL g178 ( .A(n_134), .Y(n_178) );
INVx5_ASAP7_75t_L g187 ( .A(n_137), .Y(n_187) );
AND2x6_ASAP7_75t_L g137 ( .A(n_138), .B(n_139), .Y(n_137) );
BUFx6f_ASAP7_75t_L g176 ( .A(n_138), .Y(n_176) );
BUFx3_ASAP7_75t_L g192 ( .A(n_138), .Y(n_192) );
AOI21xp5_ASAP7_75t_L g140 ( .A1(n_141), .A2(n_144), .B(n_146), .Y(n_140) );
INVx2_ASAP7_75t_L g145 ( .A(n_142), .Y(n_145) );
INVx2_ASAP7_75t_L g142 ( .A(n_143), .Y(n_142) );
INVx4_ASAP7_75t_L g171 ( .A(n_143), .Y(n_171) );
O2A1O1Ixp33_ASAP7_75t_L g188 ( .A1(n_145), .A2(n_189), .B(n_190), .C(n_191), .Y(n_188) );
O2A1O1Ixp33_ASAP7_75t_L g230 ( .A1(n_145), .A2(n_191), .B(n_231), .C(n_232), .Y(n_230) );
O2A1O1Ixp5_ASAP7_75t_L g551 ( .A1(n_145), .A2(n_552), .B(n_553), .C(n_554), .Y(n_551) );
O2A1O1Ixp33_ASAP7_75t_L g568 ( .A1(n_145), .A2(n_554), .B(n_569), .C(n_570), .Y(n_568) );
O2A1O1Ixp33_ASAP7_75t_L g490 ( .A1(n_146), .A2(n_173), .B(n_491), .C(n_492), .Y(n_490) );
INVx2_ASAP7_75t_L g146 ( .A(n_147), .Y(n_146) );
NAND2xp5_ASAP7_75t_SL g505 ( .A(n_147), .B(n_506), .Y(n_505) );
INVx1_ASAP7_75t_L g149 ( .A(n_150), .Y(n_149) );
NOR2xp33_ASAP7_75t_L g571 ( .A(n_150), .B(n_572), .Y(n_571) );
INVx2_ASAP7_75t_L g150 ( .A(n_151), .Y(n_150) );
INVx1_ASAP7_75t_L g158 ( .A(n_151), .Y(n_158) );
AOI21xp5_ASAP7_75t_L g183 ( .A1(n_151), .A2(n_184), .B(n_185), .Y(n_183) );
AOI21xp5_ASAP7_75t_L g227 ( .A1(n_151), .A2(n_228), .B(n_229), .Y(n_227) );
O2A1O1Ixp33_ASAP7_75t_L g487 ( .A1(n_151), .A2(n_216), .B(n_488), .C(n_489), .Y(n_487) );
OA21x2_ASAP7_75t_L g512 ( .A1(n_151), .A2(n_513), .B(n_520), .Y(n_512) );
AND2x2_ASAP7_75t_SL g151 ( .A(n_152), .B(n_153), .Y(n_151) );
AND2x2_ASAP7_75t_L g165 ( .A(n_152), .B(n_153), .Y(n_165) );
NAND2xp5_ASAP7_75t_L g153 ( .A(n_154), .B(n_155), .Y(n_153) );
NOR2xp33_ASAP7_75t_L g156 ( .A(n_157), .B(n_158), .Y(n_156) );
AO21x2_ASAP7_75t_L g547 ( .A1(n_158), .A2(n_548), .B(n_555), .Y(n_547) );
NAND2xp5_ASAP7_75t_L g282 ( .A(n_159), .B(n_283), .Y(n_282) );
AND2x2_ASAP7_75t_L g159 ( .A(n_160), .B(n_182), .Y(n_159) );
HB1xp67_ASAP7_75t_L g291 ( .A(n_160), .Y(n_291) );
AND2x2_ASAP7_75t_L g305 ( .A(n_160), .B(n_251), .Y(n_305) );
INVx1_ASAP7_75t_L g328 ( .A(n_160), .Y(n_328) );
NAND2xp5_ASAP7_75t_L g367 ( .A(n_160), .B(n_279), .Y(n_367) );
OR2x2_ASAP7_75t_L g404 ( .A(n_160), .B(n_249), .Y(n_404) );
INVx2_ASAP7_75t_L g160 ( .A(n_161), .Y(n_160) );
HB1xp67_ASAP7_75t_L g340 ( .A(n_161), .Y(n_340) );
AND2x2_ASAP7_75t_L g347 ( .A(n_161), .B(n_252), .Y(n_347) );
INVx2_ASAP7_75t_L g161 ( .A(n_162), .Y(n_161) );
AND2x2_ASAP7_75t_L g268 ( .A(n_162), .B(n_252), .Y(n_268) );
BUFx2_ASAP7_75t_L g296 ( .A(n_162), .Y(n_296) );
AO21x2_ASAP7_75t_L g162 ( .A1(n_163), .A2(n_166), .B(n_180), .Y(n_162) );
NOR2xp33_ASAP7_75t_L g180 ( .A(n_163), .B(n_181), .Y(n_180) );
NOR2xp33_ASAP7_75t_L g193 ( .A(n_163), .B(n_194), .Y(n_193) );
AO21x2_ASAP7_75t_L g213 ( .A1(n_163), .A2(n_214), .B(n_222), .Y(n_213) );
INVx3_ASAP7_75t_L g245 ( .A(n_163), .Y(n_245) );
NOR2xp33_ASAP7_75t_L g493 ( .A(n_163), .B(n_494), .Y(n_493) );
NOR2xp33_ASAP7_75t_L g555 ( .A(n_163), .B(n_556), .Y(n_555) );
AO21x2_ASAP7_75t_L g564 ( .A1(n_163), .A2(n_565), .B(n_571), .Y(n_564) );
INVx4_ASAP7_75t_L g163 ( .A(n_164), .Y(n_163) );
AOI21xp5_ASAP7_75t_L g201 ( .A1(n_164), .A2(n_202), .B(n_203), .Y(n_201) );
HB1xp67_ASAP7_75t_L g237 ( .A(n_164), .Y(n_237) );
BUFx6f_ASAP7_75t_L g164 ( .A(n_165), .Y(n_164) );
INVx1_ASAP7_75t_L g224 ( .A(n_165), .Y(n_224) );
NAND2xp5_ASAP7_75t_L g166 ( .A(n_167), .B(n_179), .Y(n_166) );
O2A1O1Ixp33_ASAP7_75t_L g168 ( .A1(n_169), .A2(n_170), .B(n_172), .C(n_175), .Y(n_168) );
INVx1_ASAP7_75t_L g170 ( .A(n_171), .Y(n_170) );
OAI22xp33_ASAP7_75t_L g506 ( .A1(n_171), .A2(n_173), .B1(n_507), .B2(n_508), .Y(n_506) );
NOR2xp33_ASAP7_75t_L g527 ( .A(n_171), .B(n_528), .Y(n_527) );
NOR2xp33_ASAP7_75t_L g537 ( .A(n_171), .B(n_538), .Y(n_537) );
NOR2xp33_ASAP7_75t_L g242 ( .A(n_173), .B(n_243), .Y(n_242) );
INVx2_ASAP7_75t_L g257 ( .A(n_173), .Y(n_257) );
INVx5_ASAP7_75t_L g173 ( .A(n_174), .Y(n_173) );
NOR2xp33_ASAP7_75t_L g518 ( .A(n_174), .B(n_519), .Y(n_518) );
HB1xp67_ASAP7_75t_L g175 ( .A(n_176), .Y(n_175) );
INVx3_ASAP7_75t_L g580 ( .A(n_176), .Y(n_580) );
INVx1_ASAP7_75t_L g177 ( .A(n_178), .Y(n_177) );
O2A1O1Ixp33_ASAP7_75t_L g239 ( .A1(n_178), .A2(n_187), .B(n_240), .C(n_241), .Y(n_239) );
O2A1O1Ixp33_ASAP7_75t_SL g254 ( .A1(n_178), .A2(n_187), .B(n_255), .C(n_256), .Y(n_254) );
O2A1O1Ixp33_ASAP7_75t_SL g503 ( .A1(n_178), .A2(n_187), .B(n_504), .C(n_505), .Y(n_503) );
O2A1O1Ixp33_ASAP7_75t_SL g514 ( .A1(n_178), .A2(n_187), .B(n_515), .C(n_516), .Y(n_514) );
O2A1O1Ixp33_ASAP7_75t_SL g524 ( .A1(n_178), .A2(n_187), .B(n_525), .C(n_526), .Y(n_524) );
O2A1O1Ixp33_ASAP7_75t_SL g534 ( .A1(n_178), .A2(n_187), .B(n_535), .C(n_536), .Y(n_534) );
O2A1O1Ixp33_ASAP7_75t_L g575 ( .A1(n_178), .A2(n_187), .B(n_576), .C(n_577), .Y(n_575) );
INVx5_ASAP7_75t_L g249 ( .A(n_182), .Y(n_249) );
BUFx2_ASAP7_75t_L g272 ( .A(n_182), .Y(n_272) );
AND2x2_ASAP7_75t_L g429 ( .A(n_182), .B(n_283), .Y(n_429) );
OR2x6_ASAP7_75t_L g182 ( .A(n_183), .B(n_193), .Y(n_182) );
INVx2_ASAP7_75t_L g186 ( .A(n_187), .Y(n_186) );
HB1xp67_ASAP7_75t_L g191 ( .A(n_192), .Y(n_191) );
INVx2_ASAP7_75t_L g261 ( .A(n_192), .Y(n_261) );
INVx1_ASAP7_75t_L g539 ( .A(n_192), .Y(n_539) );
INVx1_ASAP7_75t_L g195 ( .A(n_196), .Y(n_195) );
NAND2xp33_ASAP7_75t_L g196 ( .A(n_197), .B(n_234), .Y(n_196) );
OAI221xp5_ASAP7_75t_L g329 ( .A1(n_197), .A2(n_330), .B1(n_337), .B2(n_338), .C(n_341), .Y(n_329) );
OR2x2_ASAP7_75t_L g197 ( .A(n_198), .B(n_211), .Y(n_197) );
AND2x2_ASAP7_75t_L g235 ( .A(n_198), .B(n_236), .Y(n_235) );
NAND2xp5_ASAP7_75t_L g323 ( .A(n_198), .B(n_324), .Y(n_323) );
INVx1_ASAP7_75t_SL g198 ( .A(n_199), .Y(n_198) );
AND2x2_ASAP7_75t_L g264 ( .A(n_199), .B(n_212), .Y(n_264) );
NAND2xp5_ASAP7_75t_SL g274 ( .A(n_199), .B(n_213), .Y(n_274) );
OR2x2_ASAP7_75t_L g285 ( .A(n_199), .B(n_236), .Y(n_285) );
AND2x2_ASAP7_75t_L g288 ( .A(n_199), .B(n_276), .Y(n_288) );
AND2x2_ASAP7_75t_L g304 ( .A(n_199), .B(n_225), .Y(n_304) );
OR2x2_ASAP7_75t_L g320 ( .A(n_199), .B(n_213), .Y(n_320) );
NAND2xp5_ASAP7_75t_L g382 ( .A(n_199), .B(n_236), .Y(n_382) );
INVx2_ASAP7_75t_L g199 ( .A(n_200), .Y(n_199) );
NAND2xp5_ASAP7_75t_L g374 ( .A(n_200), .B(n_225), .Y(n_374) );
AND2x2_ASAP7_75t_L g377 ( .A(n_200), .B(n_213), .Y(n_377) );
AOI21xp5_ASAP7_75t_L g204 ( .A1(n_205), .A2(n_207), .B(n_208), .Y(n_204) );
AOI21xp5_ASAP7_75t_L g218 ( .A1(n_208), .A2(n_219), .B(n_220), .Y(n_218) );
INVx2_ASAP7_75t_L g208 ( .A(n_209), .Y(n_208) );
INVx3_ASAP7_75t_L g209 ( .A(n_210), .Y(n_209) );
OR2x2_ASAP7_75t_L g298 ( .A(n_211), .B(n_285), .Y(n_298) );
INVx2_ASAP7_75t_L g324 ( .A(n_211), .Y(n_324) );
OR2x2_ASAP7_75t_L g211 ( .A(n_212), .B(n_225), .Y(n_211) );
AND2x2_ASAP7_75t_L g246 ( .A(n_212), .B(n_226), .Y(n_246) );
NAND2xp5_ASAP7_75t_L g303 ( .A(n_212), .B(n_236), .Y(n_303) );
OR2x2_ASAP7_75t_L g314 ( .A(n_212), .B(n_226), .Y(n_314) );
NAND2xp5_ASAP7_75t_L g373 ( .A(n_212), .B(n_276), .Y(n_373) );
OAI221xp5_ASAP7_75t_L g406 ( .A1(n_212), .A2(n_407), .B1(n_409), .B2(n_411), .C(n_414), .Y(n_406) );
INVx5_ASAP7_75t_SL g212 ( .A(n_213), .Y(n_212) );
NAND2xp5_ASAP7_75t_L g345 ( .A(n_213), .B(n_236), .Y(n_345) );
OAI21xp5_ASAP7_75t_L g214 ( .A1(n_215), .A2(n_216), .B(n_217), .Y(n_214) );
OAI21xp5_ASAP7_75t_L g548 ( .A1(n_216), .A2(n_549), .B(n_550), .Y(n_548) );
OAI21xp5_ASAP7_75t_L g565 ( .A1(n_216), .A2(n_566), .B(n_567), .Y(n_565) );
INVx4_ASAP7_75t_L g260 ( .A(n_221), .Y(n_260) );
INVx2_ASAP7_75t_L g517 ( .A(n_221), .Y(n_517) );
NOR2xp33_ASAP7_75t_L g222 ( .A(n_223), .B(n_224), .Y(n_222) );
INVx2_ASAP7_75t_L g500 ( .A(n_224), .Y(n_500) );
NAND2xp5_ASAP7_75t_L g275 ( .A(n_225), .B(n_276), .Y(n_275) );
NOR2xp33_ASAP7_75t_L g286 ( .A(n_225), .B(n_287), .Y(n_286) );
AND2x2_ASAP7_75t_L g292 ( .A(n_225), .B(n_264), .Y(n_292) );
OR2x2_ASAP7_75t_L g336 ( .A(n_225), .B(n_236), .Y(n_336) );
NAND2xp5_ASAP7_75t_L g355 ( .A(n_225), .B(n_288), .Y(n_355) );
NAND2xp5_ASAP7_75t_L g380 ( .A(n_225), .B(n_381), .Y(n_380) );
AND2x2_ASAP7_75t_L g401 ( .A(n_225), .B(n_402), .Y(n_401) );
INVx5_ASAP7_75t_SL g225 ( .A(n_226), .Y(n_225) );
AND2x2_ASAP7_75t_SL g265 ( .A(n_226), .B(n_235), .Y(n_265) );
O2A1O1Ixp33_ASAP7_75t_SL g269 ( .A1(n_226), .A2(n_270), .B(n_273), .C(n_277), .Y(n_269) );
OR2x2_ASAP7_75t_L g307 ( .A(n_226), .B(n_303), .Y(n_307) );
OR2x2_ASAP7_75t_L g343 ( .A(n_226), .B(n_285), .Y(n_343) );
OAI311xp33_ASAP7_75t_L g349 ( .A1(n_226), .A2(n_288), .A3(n_350), .B1(n_353), .C1(n_360), .Y(n_349) );
AND2x2_ASAP7_75t_L g400 ( .A(n_226), .B(n_236), .Y(n_400) );
AND2x2_ASAP7_75t_L g408 ( .A(n_226), .B(n_263), .Y(n_408) );
HB1xp67_ASAP7_75t_L g426 ( .A(n_226), .Y(n_426) );
AND2x2_ASAP7_75t_L g443 ( .A(n_226), .B(n_264), .Y(n_443) );
OR2x6_ASAP7_75t_L g226 ( .A(n_227), .B(n_233), .Y(n_226) );
NAND2xp5_ASAP7_75t_L g234 ( .A(n_235), .B(n_246), .Y(n_234) );
AND2x2_ASAP7_75t_L g271 ( .A(n_235), .B(n_272), .Y(n_271) );
INVx2_ASAP7_75t_L g427 ( .A(n_235), .Y(n_427) );
AND2x2_ASAP7_75t_L g263 ( .A(n_236), .B(n_264), .Y(n_263) );
INVx3_ASAP7_75t_L g276 ( .A(n_236), .Y(n_276) );
HB1xp67_ASAP7_75t_L g319 ( .A(n_236), .Y(n_319) );
INVxp67_ASAP7_75t_L g358 ( .A(n_236), .Y(n_358) );
OA21x2_ASAP7_75t_L g236 ( .A1(n_237), .A2(n_238), .B(n_244), .Y(n_236) );
OA21x2_ASAP7_75t_L g522 ( .A1(n_237), .A2(n_523), .B(n_529), .Y(n_522) );
OA21x2_ASAP7_75t_L g532 ( .A1(n_237), .A2(n_533), .B(n_540), .Y(n_532) );
OA21x2_ASAP7_75t_L g573 ( .A1(n_237), .A2(n_574), .B(n_581), .Y(n_573) );
OA21x2_ASAP7_75t_L g252 ( .A1(n_245), .A2(n_253), .B(n_262), .Y(n_252) );
AND2x2_ASAP7_75t_L g436 ( .A(n_246), .B(n_284), .Y(n_436) );
AOI221xp5_ASAP7_75t_L g247 ( .A1(n_248), .A2(n_263), .B1(n_265), .B2(n_266), .C(n_269), .Y(n_247) );
AND2x2_ASAP7_75t_L g248 ( .A(n_249), .B(n_250), .Y(n_248) );
NAND2xp5_ASAP7_75t_L g267 ( .A(n_249), .B(n_268), .Y(n_267) );
AND2x2_ASAP7_75t_L g289 ( .A(n_249), .B(n_279), .Y(n_289) );
AND2x2_ASAP7_75t_L g297 ( .A(n_249), .B(n_251), .Y(n_297) );
OR2x2_ASAP7_75t_L g309 ( .A(n_249), .B(n_310), .Y(n_309) );
AND2x2_ASAP7_75t_L g327 ( .A(n_249), .B(n_328), .Y(n_327) );
AND2x2_ASAP7_75t_L g351 ( .A(n_249), .B(n_352), .Y(n_351) );
HB1xp67_ASAP7_75t_L g371 ( .A(n_249), .Y(n_371) );
AND2x2_ASAP7_75t_L g423 ( .A(n_249), .B(n_347), .Y(n_423) );
OAI31xp33_ASAP7_75t_L g431 ( .A1(n_249), .A2(n_300), .A3(n_399), .B(n_432), .Y(n_431) );
NAND2xp5_ASAP7_75t_L g326 ( .A(n_250), .B(n_327), .Y(n_326) );
INVx1_ASAP7_75t_SL g395 ( .A(n_250), .Y(n_395) );
NOR2xp33_ASAP7_75t_L g403 ( .A(n_250), .B(n_404), .Y(n_403) );
AND2x4_ASAP7_75t_L g283 ( .A(n_251), .B(n_279), .Y(n_283) );
INVx1_ASAP7_75t_L g370 ( .A(n_251), .Y(n_370) );
INVx2_ASAP7_75t_L g251 ( .A(n_252), .Y(n_251) );
AND2x2_ASAP7_75t_L g420 ( .A(n_252), .B(n_279), .Y(n_420) );
NOR2xp33_ASAP7_75t_L g258 ( .A(n_259), .B(n_260), .Y(n_258) );
NOR2xp33_ASAP7_75t_L g578 ( .A(n_260), .B(n_579), .Y(n_578) );
INVx2_ASAP7_75t_L g554 ( .A(n_261), .Y(n_554) );
INVx1_ASAP7_75t_SL g430 ( .A(n_263), .Y(n_430) );
NAND2xp5_ASAP7_75t_L g334 ( .A(n_264), .B(n_335), .Y(n_334) );
AOI22xp5_ASAP7_75t_L g414 ( .A1(n_265), .A2(n_377), .B1(n_415), .B2(n_418), .Y(n_414) );
INVx1_ASAP7_75t_L g266 ( .A(n_267), .Y(n_266) );
AND2x2_ASAP7_75t_L g278 ( .A(n_268), .B(n_279), .Y(n_278) );
INVx1_ASAP7_75t_L g337 ( .A(n_268), .Y(n_337) );
NAND2xp5_ASAP7_75t_L g442 ( .A(n_268), .B(n_289), .Y(n_442) );
INVx1_ASAP7_75t_SL g270 ( .A(n_271), .Y(n_270) );
AND2x2_ASAP7_75t_L g412 ( .A(n_271), .B(n_413), .Y(n_412) );
AOI21xp5_ASAP7_75t_L g330 ( .A1(n_272), .A2(n_331), .B(n_333), .Y(n_330) );
OR2x2_ASAP7_75t_L g338 ( .A(n_272), .B(n_339), .Y(n_338) );
AND2x2_ASAP7_75t_L g359 ( .A(n_272), .B(n_347), .Y(n_359) );
NAND2xp5_ASAP7_75t_L g398 ( .A(n_272), .B(n_370), .Y(n_398) );
NAND2xp5_ASAP7_75t_L g409 ( .A(n_272), .B(n_410), .Y(n_409) );
OAI221xp5_ASAP7_75t_SL g386 ( .A1(n_273), .A2(n_387), .B1(n_392), .B2(n_395), .C(n_396), .Y(n_386) );
OR2x2_ASAP7_75t_L g273 ( .A(n_274), .B(n_275), .Y(n_273) );
OR2x2_ASAP7_75t_L g363 ( .A(n_274), .B(n_336), .Y(n_363) );
INVx1_ASAP7_75t_L g402 ( .A(n_274), .Y(n_402) );
INVx2_ASAP7_75t_L g378 ( .A(n_275), .Y(n_378) );
INVx1_ASAP7_75t_L g312 ( .A(n_276), .Y(n_312) );
INVx1_ASAP7_75t_SL g277 ( .A(n_278), .Y(n_277) );
INVx2_ASAP7_75t_L g317 ( .A(n_279), .Y(n_317) );
NAND2xp5_ASAP7_75t_L g339 ( .A(n_279), .B(n_340), .Y(n_339) );
AND2x2_ASAP7_75t_L g346 ( .A(n_279), .B(n_347), .Y(n_346) );
OR2x2_ASAP7_75t_L g434 ( .A(n_279), .B(n_404), .Y(n_434) );
AOI222xp33_ASAP7_75t_L g280 ( .A1(n_281), .A2(n_284), .B1(n_286), .B2(n_289), .C1(n_290), .C2(n_292), .Y(n_280) );
INVxp67_ASAP7_75t_L g281 ( .A(n_282), .Y(n_281) );
AND2x2_ASAP7_75t_L g290 ( .A(n_283), .B(n_291), .Y(n_290) );
AOI22xp33_ASAP7_75t_L g360 ( .A1(n_283), .A2(n_333), .B1(n_361), .B2(n_362), .Y(n_360) );
NAND2xp5_ASAP7_75t_L g416 ( .A(n_283), .B(n_417), .Y(n_416) );
INVx1_ASAP7_75t_SL g284 ( .A(n_285), .Y(n_284) );
INVx1_ASAP7_75t_SL g287 ( .A(n_288), .Y(n_287) );
OAI21xp33_ASAP7_75t_SL g321 ( .A1(n_292), .A2(n_322), .B(n_325), .Y(n_321) );
OAI211xp5_ASAP7_75t_SL g293 ( .A1(n_294), .A2(n_298), .B(n_299), .C(n_321), .Y(n_293) );
INVxp67_ASAP7_75t_L g294 ( .A(n_295), .Y(n_294) );
AND2x2_ASAP7_75t_L g295 ( .A(n_296), .B(n_297), .Y(n_295) );
AOI221xp5_ASAP7_75t_L g299 ( .A1(n_297), .A2(n_300), .B1(n_305), .B2(n_306), .C(n_308), .Y(n_299) );
NAND2xp5_ASAP7_75t_L g384 ( .A(n_297), .B(n_385), .Y(n_384) );
INVxp67_ASAP7_75t_L g391 ( .A(n_297), .Y(n_391) );
INVx1_ASAP7_75t_L g300 ( .A(n_301), .Y(n_300) );
NAND2xp5_ASAP7_75t_L g301 ( .A(n_302), .B(n_304), .Y(n_301) );
AND2x2_ASAP7_75t_L g393 ( .A(n_302), .B(n_394), .Y(n_393) );
INVx1_ASAP7_75t_SL g302 ( .A(n_303), .Y(n_302) );
INVx1_ASAP7_75t_L g310 ( .A(n_305), .Y(n_310) );
AND2x2_ASAP7_75t_L g316 ( .A(n_305), .B(n_317), .Y(n_316) );
INVx1_ASAP7_75t_L g306 ( .A(n_307), .Y(n_306) );
OAI22xp5_ASAP7_75t_L g308 ( .A1(n_309), .A2(n_311), .B1(n_315), .B2(n_318), .Y(n_308) );
NAND2xp5_ASAP7_75t_L g311 ( .A(n_312), .B(n_313), .Y(n_311) );
NAND2xp5_ASAP7_75t_L g332 ( .A(n_312), .B(n_324), .Y(n_332) );
NAND2xp5_ASAP7_75t_L g357 ( .A(n_313), .B(n_358), .Y(n_357) );
INVx1_ASAP7_75t_SL g313 ( .A(n_314), .Y(n_313) );
INVx1_ASAP7_75t_L g315 ( .A(n_316), .Y(n_315) );
INVx1_ASAP7_75t_L g413 ( .A(n_317), .Y(n_413) );
AND2x2_ASAP7_75t_L g432 ( .A(n_317), .B(n_347), .Y(n_432) );
OR2x2_ASAP7_75t_L g318 ( .A(n_319), .B(n_320), .Y(n_318) );
INVx1_ASAP7_75t_L g322 ( .A(n_323), .Y(n_322) );
NAND2xp5_ASAP7_75t_L g440 ( .A(n_324), .B(n_381), .Y(n_440) );
INVx1_ASAP7_75t_L g325 ( .A(n_326), .Y(n_325) );
NOR2xp33_ASAP7_75t_L g438 ( .A(n_327), .B(n_395), .Y(n_438) );
INVx1_ASAP7_75t_L g331 ( .A(n_332), .Y(n_331) );
INVx1_ASAP7_75t_L g333 ( .A(n_334), .Y(n_333) );
INVx1_ASAP7_75t_L g335 ( .A(n_336), .Y(n_335) );
INVx1_ASAP7_75t_L g361 ( .A(n_339), .Y(n_361) );
BUFx2_ASAP7_75t_L g385 ( .A(n_340), .Y(n_385) );
OAI21xp5_ASAP7_75t_SL g341 ( .A1(n_342), .A2(n_344), .B(n_346), .Y(n_341) );
INVx1_ASAP7_75t_L g342 ( .A(n_343), .Y(n_342) );
INVx1_ASAP7_75t_L g344 ( .A(n_345), .Y(n_344) );
NOR3xp33_ASAP7_75t_L g348 ( .A(n_349), .B(n_364), .C(n_386), .Y(n_348) );
INVx1_ASAP7_75t_L g350 ( .A(n_351), .Y(n_350) );
OAI21xp5_ASAP7_75t_L g353 ( .A1(n_354), .A2(n_356), .B(n_359), .Y(n_353) );
INVx1_ASAP7_75t_L g354 ( .A(n_355), .Y(n_354) );
INVx1_ASAP7_75t_L g356 ( .A(n_357), .Y(n_356) );
INVx1_ASAP7_75t_SL g362 ( .A(n_363), .Y(n_362) );
A2O1A1Ixp33_ASAP7_75t_SL g364 ( .A1(n_365), .A2(n_368), .B(n_372), .C(n_375), .Y(n_364) );
NAND2xp5_ASAP7_75t_SL g397 ( .A(n_365), .B(n_398), .Y(n_397) );
INVx1_ASAP7_75t_L g365 ( .A(n_366), .Y(n_365) );
INVx1_ASAP7_75t_L g366 ( .A(n_367), .Y(n_366) );
INVx1_ASAP7_75t_L g368 ( .A(n_369), .Y(n_368) );
NOR2xp67_ASAP7_75t_SL g369 ( .A(n_370), .B(n_371), .Y(n_369) );
OR2x2_ASAP7_75t_L g372 ( .A(n_373), .B(n_374), .Y(n_372) );
INVx1_ASAP7_75t_SL g394 ( .A(n_374), .Y(n_394) );
OAI21xp5_ASAP7_75t_L g375 ( .A1(n_376), .A2(n_379), .B(n_383), .Y(n_375) );
AND2x4_ASAP7_75t_L g376 ( .A(n_377), .B(n_378), .Y(n_376) );
AND2x2_ASAP7_75t_L g399 ( .A(n_377), .B(n_400), .Y(n_399) );
INVx1_ASAP7_75t_L g379 ( .A(n_380), .Y(n_379) );
INVx1_ASAP7_75t_SL g381 ( .A(n_382), .Y(n_381) );
INVx1_ASAP7_75t_L g383 ( .A(n_384), .Y(n_383) );
INVx1_ASAP7_75t_L g387 ( .A(n_388), .Y(n_387) );
NOR2xp33_ASAP7_75t_L g388 ( .A(n_389), .B(n_391), .Y(n_388) );
INVx2_ASAP7_75t_L g389 ( .A(n_390), .Y(n_389) );
INVx1_ASAP7_75t_L g392 ( .A(n_393), .Y(n_392) );
AOI22xp33_ASAP7_75t_L g396 ( .A1(n_397), .A2(n_399), .B1(n_401), .B2(n_403), .Y(n_396) );
INVx2_ASAP7_75t_SL g417 ( .A(n_404), .Y(n_417) );
NOR3xp33_ASAP7_75t_L g405 ( .A(n_406), .B(n_421), .C(n_433), .Y(n_405) );
INVx1_ASAP7_75t_L g407 ( .A(n_408), .Y(n_407) );
INVxp67_ASAP7_75t_L g411 ( .A(n_412), .Y(n_411) );
INVxp67_ASAP7_75t_L g415 ( .A(n_416), .Y(n_415) );
NAND2xp5_ASAP7_75t_L g419 ( .A(n_417), .B(n_420), .Y(n_419) );
INVx1_ASAP7_75t_L g418 ( .A(n_419), .Y(n_418) );
OAI221xp5_ASAP7_75t_L g421 ( .A1(n_422), .A2(n_424), .B1(n_428), .B2(n_430), .C(n_431), .Y(n_421) );
A2O1A1Ixp33_ASAP7_75t_L g433 ( .A1(n_422), .A2(n_434), .B(n_435), .C(n_437), .Y(n_433) );
INVx1_ASAP7_75t_SL g422 ( .A(n_423), .Y(n_422) );
INVxp67_ASAP7_75t_L g424 ( .A(n_425), .Y(n_424) );
NOR2xp33_ASAP7_75t_L g425 ( .A(n_426), .B(n_427), .Y(n_425) );
INVx1_ASAP7_75t_L g428 ( .A(n_429), .Y(n_428) );
INVx1_ASAP7_75t_L g435 ( .A(n_436), .Y(n_435) );
AOI22xp5_ASAP7_75t_L g437 ( .A1(n_438), .A2(n_439), .B1(n_441), .B2(n_443), .Y(n_437) );
INVx1_ASAP7_75t_L g439 ( .A(n_440), .Y(n_439) );
INVx1_ASAP7_75t_L g441 ( .A(n_442), .Y(n_441) );
CKINVDCx20_ASAP7_75t_R g444 ( .A(n_445), .Y(n_444) );
INVx1_ASAP7_75t_L g446 ( .A(n_447), .Y(n_446) );
OAI22xp5_ASAP7_75t_L g474 ( .A1(n_451), .A2(n_475), .B1(n_478), .B2(n_480), .Y(n_474) );
INVx1_ASAP7_75t_L g452 ( .A(n_453), .Y(n_452) );
INVx1_ASAP7_75t_SL g453 ( .A(n_454), .Y(n_453) );
INVx1_ASAP7_75t_SL g454 ( .A(n_455), .Y(n_454) );
HB1xp67_ASAP7_75t_L g461 ( .A(n_455), .Y(n_461) );
NOR2x2_ASAP7_75t_L g760 ( .A(n_456), .B(n_479), .Y(n_760) );
INVx2_ASAP7_75t_L g456 ( .A(n_457), .Y(n_456) );
OR2x2_ASAP7_75t_L g478 ( .A(n_457), .B(n_479), .Y(n_478) );
NAND3xp33_ASAP7_75t_L g462 ( .A(n_459), .B(n_463), .C(n_761), .Y(n_462) );
INVx1_ASAP7_75t_L g460 ( .A(n_461), .Y(n_460) );
CKINVDCx20_ASAP7_75t_R g464 ( .A(n_465), .Y(n_464) );
INVx1_ASAP7_75t_L g467 ( .A(n_468), .Y(n_467) );
INVx1_ASAP7_75t_L g472 ( .A(n_469), .Y(n_472) );
INVx2_ASAP7_75t_L g475 ( .A(n_476), .Y(n_475) );
INVx2_ASAP7_75t_L g755 ( .A(n_476), .Y(n_755) );
INVx1_ASAP7_75t_L g476 ( .A(n_477), .Y(n_476) );
INVx1_ASAP7_75t_L g757 ( .A(n_478), .Y(n_757) );
INVx1_ASAP7_75t_SL g480 ( .A(n_481), .Y(n_480) );
OR5x1_ASAP7_75t_L g481 ( .A(n_482), .B(n_648), .C(n_712), .D(n_728), .E(n_743), .Y(n_481) );
NAND4xp25_ASAP7_75t_L g482 ( .A(n_483), .B(n_582), .C(n_609), .D(n_632), .Y(n_482) );
AOI21xp5_ASAP7_75t_L g483 ( .A1(n_484), .A2(n_530), .B(n_541), .Y(n_483) );
NOR2xp33_ASAP7_75t_L g484 ( .A(n_485), .B(n_495), .Y(n_484) );
HB1xp67_ASAP7_75t_L g485 ( .A(n_486), .Y(n_485) );
INVx3_ASAP7_75t_SL g561 ( .A(n_486), .Y(n_561) );
AND2x4_ASAP7_75t_L g595 ( .A(n_486), .B(n_584), .Y(n_595) );
OR2x2_ASAP7_75t_L g605 ( .A(n_486), .B(n_563), .Y(n_605) );
OR2x2_ASAP7_75t_L g651 ( .A(n_486), .B(n_498), .Y(n_651) );
AND2x2_ASAP7_75t_L g665 ( .A(n_486), .B(n_562), .Y(n_665) );
AND2x2_ASAP7_75t_L g708 ( .A(n_486), .B(n_598), .Y(n_708) );
AND2x2_ASAP7_75t_L g715 ( .A(n_486), .B(n_573), .Y(n_715) );
AND2x2_ASAP7_75t_L g734 ( .A(n_486), .B(n_624), .Y(n_734) );
AND2x2_ASAP7_75t_L g752 ( .A(n_486), .B(n_594), .Y(n_752) );
OR2x6_ASAP7_75t_L g486 ( .A(n_487), .B(n_493), .Y(n_486) );
INVx1_ASAP7_75t_L g717 ( .A(n_495), .Y(n_717) );
NAND2xp5_ASAP7_75t_L g495 ( .A(n_496), .B(n_511), .Y(n_495) );
AND2x2_ASAP7_75t_L g627 ( .A(n_496), .B(n_562), .Y(n_627) );
NAND2xp5_ASAP7_75t_L g646 ( .A(n_496), .B(n_647), .Y(n_646) );
AOI32xp33_ASAP7_75t_L g660 ( .A1(n_496), .A2(n_661), .A3(n_664), .B1(n_666), .B2(n_670), .Y(n_660) );
AND2x2_ASAP7_75t_L g730 ( .A(n_496), .B(n_624), .Y(n_730) );
INVx2_ASAP7_75t_L g496 ( .A(n_497), .Y(n_496) );
INVx1_ASAP7_75t_SL g497 ( .A(n_498), .Y(n_497) );
AND2x2_ASAP7_75t_L g594 ( .A(n_498), .B(n_563), .Y(n_594) );
NAND2xp5_ASAP7_75t_L g603 ( .A(n_498), .B(n_604), .Y(n_603) );
AND2x2_ASAP7_75t_L g636 ( .A(n_498), .B(n_583), .Y(n_636) );
NAND2xp5_ASAP7_75t_L g714 ( .A(n_498), .B(n_715), .Y(n_714) );
AO21x2_ASAP7_75t_L g498 ( .A1(n_499), .A2(n_501), .B(n_509), .Y(n_498) );
INVx1_ASAP7_75t_L g599 ( .A(n_499), .Y(n_599) );
INVx1_ASAP7_75t_L g499 ( .A(n_500), .Y(n_499) );
INVx1_ASAP7_75t_L g501 ( .A(n_502), .Y(n_501) );
OA21x2_ASAP7_75t_L g598 ( .A1(n_502), .A2(n_510), .B(n_599), .Y(n_598) );
INVx1_ASAP7_75t_L g509 ( .A(n_510), .Y(n_509) );
AND2x2_ASAP7_75t_L g601 ( .A(n_511), .B(n_545), .Y(n_601) );
AND2x2_ASAP7_75t_L g677 ( .A(n_511), .B(n_678), .Y(n_677) );
INVx1_ASAP7_75t_SL g749 ( .A(n_511), .Y(n_749) );
AND2x2_ASAP7_75t_L g511 ( .A(n_512), .B(n_521), .Y(n_511) );
OR2x2_ASAP7_75t_L g544 ( .A(n_512), .B(n_522), .Y(n_544) );
AND2x2_ASAP7_75t_L g558 ( .A(n_512), .B(n_559), .Y(n_558) );
NOR2xp33_ASAP7_75t_L g586 ( .A(n_512), .B(n_587), .Y(n_586) );
INVx2_ASAP7_75t_L g608 ( .A(n_512), .Y(n_608) );
AND2x2_ASAP7_75t_L g635 ( .A(n_512), .B(n_522), .Y(n_635) );
BUFx3_ASAP7_75t_L g638 ( .A(n_512), .Y(n_638) );
NAND2xp5_ASAP7_75t_L g645 ( .A(n_512), .B(n_613), .Y(n_645) );
NAND2xp5_ASAP7_75t_L g731 ( .A(n_512), .B(n_732), .Y(n_731) );
INVx2_ASAP7_75t_L g589 ( .A(n_521), .Y(n_589) );
AND2x2_ASAP7_75t_L g607 ( .A(n_521), .B(n_587), .Y(n_607) );
INVx2_ASAP7_75t_L g521 ( .A(n_522), .Y(n_521) );
AND2x2_ASAP7_75t_L g618 ( .A(n_522), .B(n_532), .Y(n_618) );
HB1xp67_ASAP7_75t_L g631 ( .A(n_522), .Y(n_631) );
INVx1_ASAP7_75t_L g530 ( .A(n_531), .Y(n_530) );
NAND2xp5_ASAP7_75t_L g688 ( .A(n_531), .B(n_638), .Y(n_688) );
HB1xp67_ASAP7_75t_L g531 ( .A(n_532), .Y(n_531) );
INVx1_ASAP7_75t_SL g559 ( .A(n_532), .Y(n_559) );
NAND3xp33_ASAP7_75t_L g606 ( .A(n_532), .B(n_607), .C(n_608), .Y(n_606) );
OR2x2_ASAP7_75t_L g614 ( .A(n_532), .B(n_587), .Y(n_614) );
AND2x2_ASAP7_75t_L g634 ( .A(n_532), .B(n_587), .Y(n_634) );
AND2x2_ASAP7_75t_L g678 ( .A(n_532), .B(n_547), .Y(n_678) );
AOI21xp5_ASAP7_75t_L g541 ( .A1(n_542), .A2(n_557), .B(n_560), .Y(n_541) );
NAND2xp5_ASAP7_75t_SL g542 ( .A(n_543), .B(n_545), .Y(n_542) );
AND2x2_ASAP7_75t_L g753 ( .A(n_543), .B(n_678), .Y(n_753) );
INVx1_ASAP7_75t_L g543 ( .A(n_544), .Y(n_543) );
OAI22xp5_ASAP7_75t_L g692 ( .A1(n_544), .A2(n_651), .B1(n_693), .B2(n_695), .Y(n_692) );
OR2x2_ASAP7_75t_L g699 ( .A(n_544), .B(n_614), .Y(n_699) );
OR2x2_ASAP7_75t_L g723 ( .A(n_544), .B(n_724), .Y(n_723) );
NOR2xp33_ASAP7_75t_L g736 ( .A(n_544), .B(n_643), .Y(n_736) );
AND2x2_ASAP7_75t_L g629 ( .A(n_545), .B(n_630), .Y(n_629) );
AOI21xp5_ASAP7_75t_L g716 ( .A1(n_545), .A2(n_702), .B(n_717), .Y(n_716) );
AOI32xp33_ASAP7_75t_L g737 ( .A1(n_545), .A2(n_627), .A3(n_738), .B1(n_740), .B2(n_741), .Y(n_737) );
OR2x2_ASAP7_75t_L g748 ( .A(n_545), .B(n_749), .Y(n_748) );
CKINVDCx16_ASAP7_75t_R g545 ( .A(n_546), .Y(n_545) );
OR2x2_ASAP7_75t_L g616 ( .A(n_546), .B(n_617), .Y(n_616) );
NAND2xp5_ASAP7_75t_L g695 ( .A(n_546), .B(n_630), .Y(n_695) );
BUFx3_ASAP7_75t_L g546 ( .A(n_547), .Y(n_546) );
INVx4_ASAP7_75t_L g587 ( .A(n_547), .Y(n_587) );
AND2x2_ASAP7_75t_L g653 ( .A(n_547), .B(n_618), .Y(n_653) );
AND3x2_ASAP7_75t_L g662 ( .A(n_547), .B(n_558), .C(n_663), .Y(n_662) );
INVx1_ASAP7_75t_L g557 ( .A(n_558), .Y(n_557) );
AND2x2_ASAP7_75t_L g588 ( .A(n_559), .B(n_589), .Y(n_588) );
HB1xp67_ASAP7_75t_L g643 ( .A(n_559), .Y(n_643) );
NAND2xp5_ASAP7_75t_L g724 ( .A(n_559), .B(n_587), .Y(n_724) );
NAND2xp5_ASAP7_75t_L g560 ( .A(n_561), .B(n_562), .Y(n_560) );
AND2x2_ASAP7_75t_L g583 ( .A(n_561), .B(n_584), .Y(n_583) );
AND2x2_ASAP7_75t_L g623 ( .A(n_561), .B(n_624), .Y(n_623) );
AND2x2_ASAP7_75t_L g641 ( .A(n_561), .B(n_573), .Y(n_641) );
AND2x2_ASAP7_75t_L g659 ( .A(n_561), .B(n_563), .Y(n_659) );
OR2x2_ASAP7_75t_L g673 ( .A(n_561), .B(n_674), .Y(n_673) );
AND2x2_ASAP7_75t_L g719 ( .A(n_561), .B(n_647), .Y(n_719) );
NAND2xp5_ASAP7_75t_L g597 ( .A(n_562), .B(n_598), .Y(n_597) );
AND2x2_ASAP7_75t_L g562 ( .A(n_563), .B(n_573), .Y(n_562) );
AND2x2_ASAP7_75t_L g620 ( .A(n_563), .B(n_598), .Y(n_620) );
OR2x2_ASAP7_75t_L g674 ( .A(n_563), .B(n_598), .Y(n_674) );
AND2x2_ASAP7_75t_L g727 ( .A(n_563), .B(n_584), .Y(n_727) );
INVx2_ASAP7_75t_SL g563 ( .A(n_564), .Y(n_563) );
BUFx2_ASAP7_75t_L g625 ( .A(n_564), .Y(n_625) );
AND2x2_ASAP7_75t_L g647 ( .A(n_564), .B(n_573), .Y(n_647) );
INVx2_ASAP7_75t_L g584 ( .A(n_573), .Y(n_584) );
INVx1_ASAP7_75t_L g604 ( .A(n_573), .Y(n_604) );
AOI211xp5_ASAP7_75t_L g582 ( .A1(n_583), .A2(n_585), .B(n_590), .C(n_602), .Y(n_582) );
NAND2xp5_ASAP7_75t_L g693 ( .A(n_583), .B(n_694), .Y(n_693) );
INVx1_ASAP7_75t_L g746 ( .A(n_583), .Y(n_746) );
AND2x2_ASAP7_75t_L g624 ( .A(n_584), .B(n_625), .Y(n_624) );
AND2x2_ASAP7_75t_L g585 ( .A(n_586), .B(n_588), .Y(n_585) );
NAND2xp5_ASAP7_75t_L g596 ( .A(n_587), .B(n_588), .Y(n_596) );
INVx1_ASAP7_75t_L g681 ( .A(n_587), .Y(n_681) );
NAND2xp5_ASAP7_75t_L g705 ( .A(n_587), .B(n_608), .Y(n_705) );
AND2x2_ASAP7_75t_L g721 ( .A(n_587), .B(n_635), .Y(n_721) );
NAND2xp5_ASAP7_75t_SL g703 ( .A(n_588), .B(n_704), .Y(n_703) );
INVx2_ASAP7_75t_L g612 ( .A(n_589), .Y(n_612) );
OAI22xp5_ASAP7_75t_L g590 ( .A1(n_591), .A2(n_596), .B1(n_597), .B2(n_600), .Y(n_590) );
INVx1_ASAP7_75t_L g591 ( .A(n_592), .Y(n_591) );
NOR2xp33_ASAP7_75t_L g592 ( .A(n_593), .B(n_595), .Y(n_592) );
NOR2xp33_ASAP7_75t_L g745 ( .A(n_593), .B(n_746), .Y(n_745) );
INVx1_ASAP7_75t_L g593 ( .A(n_594), .Y(n_593) );
NAND2xp5_ASAP7_75t_L g640 ( .A(n_594), .B(n_641), .Y(n_640) );
AND2x2_ASAP7_75t_L g619 ( .A(n_595), .B(n_620), .Y(n_619) );
AOI221xp5_ASAP7_75t_SL g684 ( .A1(n_595), .A2(n_637), .B1(n_685), .B2(n_690), .C(n_692), .Y(n_684) );
NAND2xp5_ASAP7_75t_L g691 ( .A(n_595), .B(n_658), .Y(n_691) );
INVx1_ASAP7_75t_L g751 ( .A(n_597), .Y(n_751) );
BUFx3_ASAP7_75t_L g658 ( .A(n_598), .Y(n_658) );
INVx1_ASAP7_75t_L g600 ( .A(n_601), .Y(n_600) );
AOI21xp33_ASAP7_75t_SL g602 ( .A1(n_603), .A2(n_605), .B(n_606), .Y(n_602) );
INVx1_ASAP7_75t_L g667 ( .A(n_604), .Y(n_667) );
NAND2xp5_ASAP7_75t_L g711 ( .A(n_604), .B(n_658), .Y(n_711) );
INVx1_ASAP7_75t_L g668 ( .A(n_605), .Y(n_668) );
NAND2xp5_ASAP7_75t_SL g669 ( .A(n_605), .B(n_658), .Y(n_669) );
INVxp67_ASAP7_75t_L g689 ( .A(n_607), .Y(n_689) );
AND2x2_ASAP7_75t_L g630 ( .A(n_608), .B(n_631), .Y(n_630) );
O2A1O1Ixp33_ASAP7_75t_L g609 ( .A1(n_610), .A2(n_615), .B(n_619), .C(n_621), .Y(n_609) );
INVx1_ASAP7_75t_L g610 ( .A(n_611), .Y(n_610) );
NAND2xp5_ASAP7_75t_L g611 ( .A(n_612), .B(n_613), .Y(n_611) );
INVx1_ASAP7_75t_SL g644 ( .A(n_612), .Y(n_644) );
NAND2xp5_ASAP7_75t_L g655 ( .A(n_613), .B(n_644), .Y(n_655) );
NAND2xp5_ASAP7_75t_L g686 ( .A(n_613), .B(n_635), .Y(n_686) );
INVx2_ASAP7_75t_SL g613 ( .A(n_614), .Y(n_613) );
INVx1_ASAP7_75t_L g615 ( .A(n_616), .Y(n_615) );
OAI22xp5_ASAP7_75t_L g621 ( .A1(n_616), .A2(n_622), .B1(n_626), .B2(n_628), .Y(n_621) );
INVx1_ASAP7_75t_SL g617 ( .A(n_618), .Y(n_617) );
AND2x2_ASAP7_75t_L g637 ( .A(n_618), .B(n_638), .Y(n_637) );
AND2x2_ASAP7_75t_L g682 ( .A(n_618), .B(n_683), .Y(n_682) );
OAI21xp33_ASAP7_75t_L g685 ( .A1(n_620), .A2(n_686), .B(n_687), .Y(n_685) );
INVx1_ASAP7_75t_SL g622 ( .A(n_623), .Y(n_622) );
AOI221xp5_ASAP7_75t_L g632 ( .A1(n_624), .A2(n_633), .B1(n_636), .B2(n_637), .C(n_639), .Y(n_632) );
NAND2xp5_ASAP7_75t_L g701 ( .A(n_624), .B(n_658), .Y(n_701) );
NAND2xp5_ASAP7_75t_L g707 ( .A(n_624), .B(n_708), .Y(n_707) );
INVx1_ASAP7_75t_L g626 ( .A(n_627), .Y(n_626) );
INVx1_ASAP7_75t_L g628 ( .A(n_629), .Y(n_628) );
INVx1_ASAP7_75t_L g740 ( .A(n_630), .Y(n_740) );
INVxp67_ASAP7_75t_L g663 ( .A(n_631), .Y(n_663) );
INVx1_ASAP7_75t_L g670 ( .A(n_633), .Y(n_670) );
AND2x2_ASAP7_75t_L g633 ( .A(n_634), .B(n_635), .Y(n_633) );
AND2x2_ASAP7_75t_L g709 ( .A(n_634), .B(n_638), .Y(n_709) );
INVx1_ASAP7_75t_L g683 ( .A(n_638), .Y(n_683) );
NAND2xp5_ASAP7_75t_SL g713 ( .A(n_638), .B(n_653), .Y(n_713) );
OAI32xp33_ASAP7_75t_L g639 ( .A1(n_640), .A2(n_642), .A3(n_644), .B1(n_645), .B2(n_646), .Y(n_639) );
INVx1_ASAP7_75t_L g642 ( .A(n_643), .Y(n_642) );
INVx2_ASAP7_75t_SL g652 ( .A(n_647), .Y(n_652) );
NAND2xp5_ASAP7_75t_L g696 ( .A(n_647), .B(n_679), .Y(n_696) );
NAND2xp5_ASAP7_75t_L g739 ( .A(n_647), .B(n_708), .Y(n_739) );
NAND2x1p5_ASAP7_75t_L g747 ( .A(n_647), .B(n_658), .Y(n_747) );
NAND5xp2_ASAP7_75t_L g648 ( .A(n_649), .B(n_671), .C(n_684), .D(n_696), .E(n_697), .Y(n_648) );
AOI221xp5_ASAP7_75t_L g649 ( .A1(n_650), .A2(n_653), .B1(n_654), .B2(n_656), .C(n_660), .Y(n_649) );
NOR2xp33_ASAP7_75t_L g650 ( .A(n_651), .B(n_652), .Y(n_650) );
INVx1_ASAP7_75t_L g654 ( .A(n_655), .Y(n_654) );
NAND2xp33_ASAP7_75t_SL g675 ( .A(n_655), .B(n_676), .Y(n_675) );
INVx1_ASAP7_75t_L g656 ( .A(n_657), .Y(n_656) );
NAND2xp5_ASAP7_75t_L g657 ( .A(n_658), .B(n_659), .Y(n_657) );
NAND2xp5_ASAP7_75t_L g726 ( .A(n_658), .B(n_727), .Y(n_726) );
AOI22xp33_ASAP7_75t_L g671 ( .A1(n_659), .A2(n_672), .B1(n_675), .B2(n_679), .Y(n_671) );
INVx2_ASAP7_75t_SL g661 ( .A(n_662), .Y(n_661) );
OAI211xp5_ASAP7_75t_SL g666 ( .A1(n_662), .A2(n_667), .B(n_668), .C(n_669), .Y(n_666) );
INVx1_ASAP7_75t_L g664 ( .A(n_665), .Y(n_664) );
INVx1_ASAP7_75t_L g672 ( .A(n_673), .Y(n_672) );
INVx1_ASAP7_75t_SL g694 ( .A(n_674), .Y(n_694) );
INVx1_ASAP7_75t_SL g676 ( .A(n_677), .Y(n_676) );
INVx1_ASAP7_75t_SL g679 ( .A(n_680), .Y(n_679) );
NAND2xp5_ASAP7_75t_L g680 ( .A(n_681), .B(n_682), .Y(n_680) );
NAND2xp5_ASAP7_75t_L g742 ( .A(n_683), .B(n_732), .Y(n_742) );
OR2x2_ASAP7_75t_L g687 ( .A(n_688), .B(n_689), .Y(n_687) );
INVx1_ASAP7_75t_L g690 ( .A(n_691), .Y(n_690) );
AOI222xp33_ASAP7_75t_L g697 ( .A1(n_698), .A2(n_700), .B1(n_702), .B2(n_706), .C1(n_709), .C2(n_710), .Y(n_697) );
INVx1_ASAP7_75t_L g698 ( .A(n_699), .Y(n_698) );
INVx1_ASAP7_75t_L g700 ( .A(n_701), .Y(n_700) );
INVx1_ASAP7_75t_L g702 ( .A(n_703), .Y(n_702) );
INVx1_ASAP7_75t_L g704 ( .A(n_705), .Y(n_704) );
INVx1_ASAP7_75t_L g706 ( .A(n_707), .Y(n_706) );
INVx1_ASAP7_75t_L g710 ( .A(n_711), .Y(n_710) );
OAI221xp5_ASAP7_75t_L g712 ( .A1(n_713), .A2(n_714), .B1(n_716), .B2(n_718), .C(n_720), .Y(n_712) );
INVx1_ASAP7_75t_SL g718 ( .A(n_719), .Y(n_718) );
OAI21xp33_ASAP7_75t_L g720 ( .A1(n_721), .A2(n_722), .B(n_725), .Y(n_720) );
INVx2_ASAP7_75t_L g722 ( .A(n_723), .Y(n_722) );
INVx1_ASAP7_75t_L g732 ( .A(n_724), .Y(n_732) );
INVx1_ASAP7_75t_L g725 ( .A(n_726), .Y(n_725) );
OAI221xp5_ASAP7_75t_L g728 ( .A1(n_729), .A2(n_731), .B1(n_733), .B2(n_735), .C(n_737), .Y(n_728) );
INVx1_ASAP7_75t_L g729 ( .A(n_730), .Y(n_729) );
INVx1_ASAP7_75t_SL g733 ( .A(n_734), .Y(n_733) );
INVxp67_ASAP7_75t_L g735 ( .A(n_736), .Y(n_735) );
INVx1_ASAP7_75t_L g738 ( .A(n_739), .Y(n_738) );
INVx1_ASAP7_75t_L g741 ( .A(n_742), .Y(n_741) );
A2O1A1Ixp33_ASAP7_75t_L g743 ( .A1(n_744), .A2(n_747), .B(n_748), .C(n_750), .Y(n_743) );
INVxp67_ASAP7_75t_L g744 ( .A(n_745), .Y(n_744) );
OAI21xp33_ASAP7_75t_L g750 ( .A1(n_751), .A2(n_752), .B(n_753), .Y(n_750) );
INVx2_ASAP7_75t_L g756 ( .A(n_757), .Y(n_756) );
INVx1_ASAP7_75t_SL g758 ( .A(n_759), .Y(n_758) );
INVx2_ASAP7_75t_L g759 ( .A(n_760), .Y(n_759) );
INVx1_ASAP7_75t_SL g761 ( .A(n_762), .Y(n_761) );
INVx1_ASAP7_75t_SL g762 ( .A(n_763), .Y(n_762) );
CKINVDCx20_ASAP7_75t_R g764 ( .A(n_765), .Y(n_764) );
endmodule