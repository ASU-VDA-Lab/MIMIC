module real_aes_6713_n_77 (n_17, n_28, n_76, n_56, n_34, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_43, n_54, n_35, n_42, n_15, n_9, n_23, n_72, n_44, n_7, n_4, n_6, n_12, n_68, n_69, n_46, n_59, n_25, n_73, n_48, n_37, n_70, n_50, n_26, n_13, n_24, n_2, n_55, n_62, n_67, n_33, n_14, n_11, n_16, n_39, n_5, n_45, n_60, n_38, n_0, n_63, n_1, n_53, n_36, n_77);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_43;
input n_54;
input n_35;
input n_42;
input n_15;
input n_9;
input n_23;
input n_72;
input n_44;
input n_7;
input n_4;
input n_6;
input n_12;
input n_68;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_48;
input n_37;
input n_70;
input n_50;
input n_26;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_67;
input n_33;
input n_14;
input n_11;
input n_16;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_0;
input n_63;
input n_1;
input n_53;
input n_36;
output n_77;
wire n_480;
wire n_113;
wire n_476;
wire n_187;
wire n_436;
wire n_90;
wire n_257;
wire n_390;
wire n_185;
wire n_285;
wire n_485;
wire n_222;
wire n_503;
wire n_287;
wire n_357;
wire n_386;
wire n_518;
wire n_254;
wire n_207;
wire n_469;
wire n_83;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_445;
wire n_299;
wire n_322;
wire n_328;
wire n_318;
wire n_355;
wire n_239;
wire n_100;
wire n_423;
wire n_458;
wire n_444;
wire n_112;
wire n_319;
wire n_364;
wire n_421;
wire n_329;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_242;
wire n_169;
wire n_376;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_448;
wire n_341;
wire n_232;
wire n_460;
wire n_401;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_320;
wire n_260;
wire n_97;
wire n_186;
wire n_138;
wire n_379;
wire n_374;
wire n_453;
wire n_235;
wire n_399;
wire n_378;
wire n_245;
wire n_161;
wire n_189;
wire n_271;
wire n_489;
wire n_427;
wire n_145;
wire n_415;
wire n_227;
wire n_92;
wire n_519;
wire n_510;
wire n_330;
wire n_388;
wire n_512;
wire n_395;
wire n_332;
wire n_292;
wire n_400;
wire n_116;
wire n_94;
wire n_289;
wire n_462;
wire n_280;
wire n_333;
wire n_213;
wire n_478;
wire n_356;
wire n_408;
wire n_184;
wire n_372;
wire n_202;
wire n_495;
wire n_370;
wire n_98;
wire n_384;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_82;
wire n_467;
wire n_327;
wire n_106;
wire n_466;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_517;
wire n_174;
wire n_104;
wire n_211;
wire n_281;
wire n_496;
wire n_173;
wire n_468;
wire n_234;
wire n_284;
wire n_153;
wire n_316;
wire n_178;
wire n_409;
wire n_298;
wire n_439;
wire n_506;
wire n_513;
wire n_297;
wire n_383;
wire n_119;
wire n_310;
wire n_455;
wire n_504;
wire n_164;
wire n_231;
wire n_102;
wire n_454;
wire n_122;
wire n_443;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_80;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_367;
wire n_267;
wire n_218;
wire n_204;
wire n_339;
wire n_398;
wire n_89;
wire n_277;
wire n_425;
wire n_331;
wire n_93;
wire n_182;
wire n_363;
wire n_417;
wire n_449;
wire n_323;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_142;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_368;
wire n_505;
wire n_502;
wire n_434;
wire n_250;
wire n_85;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_402;
wire n_171;
wire n_87;
wire n_78;
wire n_451;
wire n_146;
wire n_432;
wire n_255;
wire n_226;
wire n_286;
wire n_416;
wire n_410;
wire n_120;
wire n_490;
wire n_261;
wire n_238;
wire n_391;
wire n_360;
wire n_165;
wire n_361;
wire n_246;
wire n_176;
wire n_412;
wire n_163;
wire n_488;
wire n_501;
wire n_251;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_115;
wire n_96;
wire n_110;
wire n_392;
wire n_150;
wire n_147;
wire n_288;
wire n_404;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_95;
wire n_188;
wire n_269;
wire n_430;
wire n_201;
wire n_413;
wire n_471;
wire n_306;
wire n_158;
wire n_366;
wire n_346;
wire n_193;
wire n_397;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_109;
wire n_203;
wire n_470;
wire n_81;
wire n_133;
wire n_494;
wire n_377;
wire n_273;
wire n_114;
wire n_276;
wire n_295;
wire n_382;
wire n_265;
wire n_354;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_419;
wire n_217;
wire n_486;
wire n_411;
wire n_291;
wire n_148;
wire n_481;
wire n_498;
wire n_88;
wire n_159;
wire n_108;
wire n_373;
wire n_233;
wire n_487;
wire n_290;
wire n_365;
wire n_155;
wire n_243;
wire n_268;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_101;
wire n_309;
wire n_344;
wire n_229;
wire n_107;
wire n_482;
wire n_520;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_262;
wire n_134;
wire n_349;
wire n_336;
wire n_420;
wire n_195;
wire n_438;
wire n_300;
wire n_252;
wire n_283;
wire n_314;
wire n_249;
wire n_446;
wire n_221;
wire n_156;
wire n_359;
wire n_456;
wire n_312;
wire n_183;
wire n_266;
wire n_205;
wire n_433;
wire n_335;
wire n_177;
wire n_516;
wire n_313;
wire n_140;
wire n_521;
wire n_418;
wire n_422;
wire n_219;
wire n_180;
wire n_212;
wire n_210;
wire n_325;
wire n_338;
wire n_479;
wire n_442;
wire n_371;
wire n_166;
wire n_103;
wire n_224;
wire n_151;
wire n_130;
wire n_253;
wire n_459;
wire n_99;
wire n_440;
wire n_152;
wire n_198;
wire n_228;
wire n_272;
wire n_196;
wire n_347;
wire n_315;
wire n_414;
wire n_123;
wire n_279;
wire n_79;
wire n_497;
wire n_514;
wire n_270;
wire n_507;
wire n_305;
wire n_450;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_465;
wire n_473;
wire n_474;
wire n_170;
wire n_86;
wire n_375;
wire n_340;
wire n_483;
wire n_380;
wire n_394;
wire n_168;
wire n_241;
wire n_175;
wire n_105;
wire n_84;
wire n_294;
wire n_393;
wire n_258;
wire n_206;
wire n_307;
wire n_500;
wire n_463;
wire n_396;
wire n_447;
wire n_342;
wire n_348;
wire n_403;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_143;
wire n_192;
wire n_475;
wire n_264;
wire n_237;
wire n_91;
AOI22xp5_ASAP7_75t_L g79 ( .A1(n_0), .A2(n_80), .B1(n_81), .B2(n_163), .Y(n_79) );
INVx1_ASAP7_75t_L g163 ( .A(n_0), .Y(n_163) );
INVx1_ASAP7_75t_L g288 ( .A(n_1), .Y(n_288) );
AOI22xp33_ASAP7_75t_L g238 ( .A1(n_2), .A2(n_31), .B1(n_201), .B2(n_213), .Y(n_238) );
NAND2xp5_ASAP7_75t_L g277 ( .A(n_3), .B(n_244), .Y(n_277) );
INVx1_ASAP7_75t_L g185 ( .A(n_4), .Y(n_185) );
AND2x6_ASAP7_75t_L g216 ( .A(n_4), .B(n_183), .Y(n_216) );
NAND2xp5_ASAP7_75t_L g508 ( .A(n_4), .B(n_509), .Y(n_508) );
CKINVDCx20_ASAP7_75t_R g162 ( .A(n_5), .Y(n_162) );
AO22x2_ASAP7_75t_L g97 ( .A1(n_6), .A2(n_27), .B1(n_89), .B2(n_94), .Y(n_97) );
INVx1_ASAP7_75t_L g282 ( .A(n_7), .Y(n_282) );
INVx1_ASAP7_75t_L g197 ( .A(n_8), .Y(n_197) );
AOI22xp33_ASAP7_75t_SL g123 ( .A1(n_9), .A2(n_35), .B1(n_124), .B2(n_127), .Y(n_123) );
NAND2xp5_ASAP7_75t_L g204 ( .A(n_10), .B(n_205), .Y(n_204) );
NAND2xp5_ASAP7_75t_L g260 ( .A(n_11), .B(n_242), .Y(n_260) );
AO32x2_ASAP7_75t_L g236 ( .A1(n_12), .A2(n_237), .A3(n_241), .B1(n_243), .B2(n_244), .Y(n_236) );
NAND2xp5_ASAP7_75t_SL g211 ( .A(n_13), .B(n_201), .Y(n_211) );
AO22x2_ASAP7_75t_L g99 ( .A1(n_14), .A2(n_29), .B1(n_89), .B2(n_90), .Y(n_99) );
NAND2xp5_ASAP7_75t_L g290 ( .A(n_15), .B(n_242), .Y(n_290) );
AOI22xp33_ASAP7_75t_L g240 ( .A1(n_16), .A2(n_41), .B1(n_201), .B2(n_213), .Y(n_240) );
AOI22xp33_ASAP7_75t_SL g253 ( .A1(n_17), .A2(n_61), .B1(n_201), .B2(n_205), .Y(n_253) );
NAND2xp5_ASAP7_75t_SL g230 ( .A(n_18), .B(n_201), .Y(n_230) );
OAI22xp5_ASAP7_75t_SL g168 ( .A1(n_19), .A2(n_34), .B1(n_169), .B2(n_170), .Y(n_168) );
INVx1_ASAP7_75t_L g169 ( .A(n_19), .Y(n_169) );
BUFx6f_ASAP7_75t_L g209 ( .A(n_20), .Y(n_209) );
NAND2xp5_ASAP7_75t_L g302 ( .A(n_21), .B(n_193), .Y(n_302) );
XOR2xp5_ASAP7_75t_L g517 ( .A(n_22), .B(n_80), .Y(n_517) );
CKINVDCx20_ASAP7_75t_R g134 ( .A(n_23), .Y(n_134) );
NAND2xp5_ASAP7_75t_L g234 ( .A(n_24), .B(n_193), .Y(n_234) );
AOI22xp5_ASAP7_75t_SL g84 ( .A1(n_25), .A2(n_43), .B1(n_85), .B2(n_100), .Y(n_84) );
INVx2_ASAP7_75t_L g203 ( .A(n_26), .Y(n_203) );
NAND2xp5_ASAP7_75t_SL g297 ( .A(n_28), .B(n_201), .Y(n_297) );
OAI221xp5_ASAP7_75t_L g176 ( .A1(n_29), .A2(n_46), .B1(n_59), .B2(n_177), .C(n_178), .Y(n_176) );
INVxp67_ASAP7_75t_L g179 ( .A(n_29), .Y(n_179) );
NAND2xp5_ASAP7_75t_L g217 ( .A(n_30), .B(n_193), .Y(n_217) );
AOI22xp5_ASAP7_75t_L g145 ( .A1(n_32), .A2(n_56), .B1(n_146), .B2(n_150), .Y(n_145) );
AOI22xp5_ASAP7_75t_L g104 ( .A1(n_33), .A2(n_49), .B1(n_105), .B2(n_111), .Y(n_104) );
INVx1_ASAP7_75t_L g170 ( .A(n_34), .Y(n_170) );
NAND2xp5_ASAP7_75t_SL g270 ( .A(n_36), .B(n_201), .Y(n_270) );
AOI22xp33_ASAP7_75t_L g251 ( .A1(n_37), .A2(n_69), .B1(n_213), .B2(n_252), .Y(n_251) );
AOI22xp5_ASAP7_75t_L g165 ( .A1(n_38), .A2(n_166), .B1(n_167), .B2(n_168), .Y(n_165) );
INVx1_ASAP7_75t_L g166 ( .A(n_38), .Y(n_166) );
NAND2xp5_ASAP7_75t_SL g273 ( .A(n_38), .B(n_201), .Y(n_273) );
NAND2xp5_ASAP7_75t_L g284 ( .A(n_39), .B(n_201), .Y(n_284) );
NAND2xp5_ASAP7_75t_L g274 ( .A(n_40), .B(n_275), .Y(n_274) );
AOI22xp33_ASAP7_75t_SL g264 ( .A1(n_42), .A2(n_47), .B1(n_201), .B2(n_205), .Y(n_264) );
INVx1_ASAP7_75t_L g516 ( .A(n_42), .Y(n_516) );
NAND2xp5_ASAP7_75t_SL g200 ( .A(n_44), .B(n_201), .Y(n_200) );
NAND2xp5_ASAP7_75t_SL g301 ( .A(n_45), .B(n_201), .Y(n_301) );
AO22x2_ASAP7_75t_L g88 ( .A1(n_46), .A2(n_64), .B1(n_89), .B2(n_90), .Y(n_88) );
INVxp67_ASAP7_75t_L g180 ( .A(n_46), .Y(n_180) );
AOI22xp5_ASAP7_75t_SL g504 ( .A1(n_47), .A2(n_80), .B1(n_81), .B2(n_505), .Y(n_504) );
INVx1_ASAP7_75t_L g505 ( .A(n_47), .Y(n_505) );
INVx1_ASAP7_75t_L g183 ( .A(n_48), .Y(n_183) );
CKINVDCx20_ASAP7_75t_R g144 ( .A(n_50), .Y(n_144) );
CKINVDCx20_ASAP7_75t_R g157 ( .A(n_51), .Y(n_157) );
INVx1_ASAP7_75t_L g196 ( .A(n_52), .Y(n_196) );
NAND2xp5_ASAP7_75t_L g289 ( .A(n_53), .B(n_201), .Y(n_289) );
CKINVDCx20_ASAP7_75t_R g177 ( .A(n_54), .Y(n_177) );
AO32x2_ASAP7_75t_L g249 ( .A1(n_55), .A2(n_243), .A3(n_244), .B1(n_250), .B2(n_254), .Y(n_249) );
INVx1_ASAP7_75t_L g300 ( .A(n_57), .Y(n_300) );
INVx1_ASAP7_75t_L g225 ( .A(n_58), .Y(n_225) );
AO22x2_ASAP7_75t_L g93 ( .A1(n_59), .A2(n_71), .B1(n_89), .B2(n_94), .Y(n_93) );
NAND2xp5_ASAP7_75t_SL g226 ( .A(n_60), .B(n_205), .Y(n_226) );
NAND2xp5_ASAP7_75t_L g212 ( .A(n_62), .B(n_213), .Y(n_212) );
NAND2xp5_ASAP7_75t_SL g231 ( .A(n_63), .B(n_205), .Y(n_231) );
INVx2_ASAP7_75t_L g194 ( .A(n_65), .Y(n_194) );
AOI22xp5_ASAP7_75t_L g164 ( .A1(n_66), .A2(n_165), .B1(n_171), .B2(n_172), .Y(n_164) );
INVx1_ASAP7_75t_L g171 ( .A(n_66), .Y(n_171) );
AOI22xp5_ASAP7_75t_SL g113 ( .A1(n_67), .A2(n_75), .B1(n_114), .B2(n_119), .Y(n_113) );
NAND2xp5_ASAP7_75t_L g271 ( .A(n_68), .B(n_205), .Y(n_271) );
AOI22xp33_ASAP7_75t_L g263 ( .A1(n_70), .A2(n_76), .B1(n_205), .B2(n_206), .Y(n_263) );
CKINVDCx20_ASAP7_75t_R g139 ( .A(n_72), .Y(n_139) );
INVx1_ASAP7_75t_L g89 ( .A(n_73), .Y(n_89) );
INVx1_ASAP7_75t_L g91 ( .A(n_73), .Y(n_91) );
NAND2xp5_ASAP7_75t_L g298 ( .A(n_74), .B(n_205), .Y(n_298) );
AOI221xp5_ASAP7_75t_L g77 ( .A1(n_78), .A2(n_173), .B1(n_186), .B2(n_497), .C(n_503), .Y(n_77) );
XOR2xp5_ASAP7_75t_L g78 ( .A(n_79), .B(n_164), .Y(n_78) );
CKINVDCx20_ASAP7_75t_R g80 ( .A(n_81), .Y(n_80) );
HB1xp67_ASAP7_75t_L g81 ( .A(n_82), .Y(n_81) );
NAND3x1_ASAP7_75t_SL g82 ( .A(n_83), .B(n_112), .C(n_129), .Y(n_82) );
AND2x2_ASAP7_75t_L g83 ( .A(n_84), .B(n_104), .Y(n_83) );
BUFx3_ASAP7_75t_L g85 ( .A(n_86), .Y(n_85) );
AND2x2_ASAP7_75t_L g86 ( .A(n_87), .B(n_95), .Y(n_86) );
AND2x2_ASAP7_75t_L g102 ( .A(n_87), .B(n_103), .Y(n_102) );
AND2x2_ASAP7_75t_L g87 ( .A(n_88), .B(n_92), .Y(n_87) );
INVx2_ASAP7_75t_L g109 ( .A(n_88), .Y(n_109) );
NAND2xp5_ASAP7_75t_L g122 ( .A(n_88), .B(n_93), .Y(n_122) );
AND2x2_ASAP7_75t_L g138 ( .A(n_88), .B(n_97), .Y(n_138) );
INVx1_ASAP7_75t_L g90 ( .A(n_91), .Y(n_90) );
INVx1_ASAP7_75t_L g94 ( .A(n_91), .Y(n_94) );
INVx1_ASAP7_75t_L g152 ( .A(n_92), .Y(n_152) );
INVx1_ASAP7_75t_L g92 ( .A(n_93), .Y(n_92) );
INVx1_ASAP7_75t_L g110 ( .A(n_93), .Y(n_110) );
AND2x2_ASAP7_75t_L g126 ( .A(n_93), .B(n_109), .Y(n_126) );
INVx1_ASAP7_75t_L g149 ( .A(n_93), .Y(n_149) );
AND2x2_ASAP7_75t_L g107 ( .A(n_95), .B(n_108), .Y(n_107) );
AND2x4_ASAP7_75t_L g120 ( .A(n_95), .B(n_121), .Y(n_120) );
AND2x4_ASAP7_75t_L g125 ( .A(n_95), .B(n_126), .Y(n_125) );
AND2x2_ASAP7_75t_L g95 ( .A(n_96), .B(n_98), .Y(n_95) );
AND2x2_ASAP7_75t_L g103 ( .A(n_96), .B(n_99), .Y(n_103) );
OR2x2_ASAP7_75t_L g118 ( .A(n_96), .B(n_99), .Y(n_118) );
INVx2_ASAP7_75t_L g96 ( .A(n_97), .Y(n_96) );
AND2x2_ASAP7_75t_L g153 ( .A(n_97), .B(n_99), .Y(n_153) );
INVx1_ASAP7_75t_L g128 ( .A(n_98), .Y(n_128) );
AND2x2_ASAP7_75t_L g161 ( .A(n_98), .B(n_149), .Y(n_161) );
INVx2_ASAP7_75t_L g98 ( .A(n_99), .Y(n_98) );
INVx3_ASAP7_75t_L g100 ( .A(n_101), .Y(n_100) );
INVx8_ASAP7_75t_L g101 ( .A(n_102), .Y(n_101) );
AND2x4_ASAP7_75t_L g111 ( .A(n_103), .B(n_108), .Y(n_111) );
NAND2x1p5_ASAP7_75t_L g133 ( .A(n_103), .B(n_126), .Y(n_133) );
INVx3_ASAP7_75t_L g105 ( .A(n_106), .Y(n_105) );
INVx2_ASAP7_75t_L g106 ( .A(n_107), .Y(n_106) );
AND2x6_ASAP7_75t_L g116 ( .A(n_108), .B(n_117), .Y(n_116) );
AND2x6_ASAP7_75t_L g156 ( .A(n_108), .B(n_153), .Y(n_156) );
AND2x2_ASAP7_75t_L g108 ( .A(n_109), .B(n_110), .Y(n_108) );
AND2x2_ASAP7_75t_L g112 ( .A(n_113), .B(n_123), .Y(n_112) );
INVx4_ASAP7_75t_L g114 ( .A(n_115), .Y(n_114) );
INVx11_ASAP7_75t_L g115 ( .A(n_116), .Y(n_115) );
INVx2_ASAP7_75t_L g117 ( .A(n_118), .Y(n_117) );
OR2x2_ASAP7_75t_L g142 ( .A(n_118), .B(n_143), .Y(n_142) );
BUFx3_ASAP7_75t_L g119 ( .A(n_120), .Y(n_119) );
AND2x2_ASAP7_75t_L g127 ( .A(n_121), .B(n_128), .Y(n_127) );
INVx1_ASAP7_75t_L g121 ( .A(n_122), .Y(n_121) );
BUFx6f_ASAP7_75t_L g124 ( .A(n_125), .Y(n_124) );
INVx1_ASAP7_75t_L g143 ( .A(n_126), .Y(n_143) );
NAND2x1p5_ASAP7_75t_L g137 ( .A(n_128), .B(n_138), .Y(n_137) );
NOR3xp33_ASAP7_75t_L g129 ( .A(n_130), .B(n_140), .C(n_154), .Y(n_129) );
OAI22xp5_ASAP7_75t_SL g130 ( .A1(n_131), .A2(n_134), .B1(n_135), .B2(n_139), .Y(n_130) );
INVx2_ASAP7_75t_L g131 ( .A(n_132), .Y(n_131) );
INVx1_ASAP7_75t_L g132 ( .A(n_133), .Y(n_132) );
INVx3_ASAP7_75t_SL g135 ( .A(n_136), .Y(n_135) );
INVx4_ASAP7_75t_L g136 ( .A(n_137), .Y(n_136) );
AND2x4_ASAP7_75t_L g147 ( .A(n_138), .B(n_148), .Y(n_147) );
AND2x4_ASAP7_75t_L g160 ( .A(n_138), .B(n_161), .Y(n_160) );
OAI21xp5_ASAP7_75t_SL g140 ( .A1(n_141), .A2(n_144), .B(n_145), .Y(n_140) );
BUFx6f_ASAP7_75t_L g141 ( .A(n_142), .Y(n_141) );
BUFx6f_ASAP7_75t_L g146 ( .A(n_147), .Y(n_146) );
INVx1_ASAP7_75t_L g148 ( .A(n_149), .Y(n_148) );
BUFx6f_ASAP7_75t_L g150 ( .A(n_151), .Y(n_150) );
AND2x4_ASAP7_75t_L g151 ( .A(n_152), .B(n_153), .Y(n_151) );
OAI22xp5_ASAP7_75t_SL g154 ( .A1(n_155), .A2(n_157), .B1(n_158), .B2(n_162), .Y(n_154) );
INVx4_ASAP7_75t_L g155 ( .A(n_156), .Y(n_155) );
INVx2_ASAP7_75t_L g158 ( .A(n_159), .Y(n_158) );
BUFx6f_ASAP7_75t_L g159 ( .A(n_160), .Y(n_159) );
CKINVDCx20_ASAP7_75t_R g172 ( .A(n_165), .Y(n_172) );
CKINVDCx20_ASAP7_75t_R g167 ( .A(n_168), .Y(n_167) );
CKINVDCx20_ASAP7_75t_R g173 ( .A(n_174), .Y(n_173) );
CKINVDCx20_ASAP7_75t_R g174 ( .A(n_175), .Y(n_174) );
AND3x1_ASAP7_75t_SL g175 ( .A(n_176), .B(n_181), .C(n_184), .Y(n_175) );
INVxp67_ASAP7_75t_L g509 ( .A(n_176), .Y(n_509) );
NOR2xp33_ASAP7_75t_L g178 ( .A(n_179), .B(n_180), .Y(n_178) );
INVx1_ASAP7_75t_SL g510 ( .A(n_181), .Y(n_510) );
OAI21xp5_ASAP7_75t_L g512 ( .A1(n_181), .A2(n_513), .B(n_515), .Y(n_512) );
INVx1_ASAP7_75t_L g521 ( .A(n_181), .Y(n_521) );
INVx1_ASAP7_75t_L g181 ( .A(n_182), .Y(n_181) );
NAND2xp5_ASAP7_75t_SL g515 ( .A(n_182), .B(n_185), .Y(n_515) );
HB1xp67_ASAP7_75t_L g182 ( .A(n_183), .Y(n_182) );
OR2x2_ASAP7_75t_SL g520 ( .A(n_184), .B(n_521), .Y(n_520) );
CKINVDCx20_ASAP7_75t_R g184 ( .A(n_185), .Y(n_184) );
OR2x2_ASAP7_75t_L g186 ( .A(n_187), .B(n_419), .Y(n_186) );
NAND5xp2_ASAP7_75t_L g187 ( .A(n_188), .B(n_338), .C(n_353), .D(n_379), .E(n_401), .Y(n_187) );
NOR2xp33_ASAP7_75t_SL g188 ( .A(n_189), .B(n_318), .Y(n_188) );
OAI221xp5_ASAP7_75t_L g189 ( .A1(n_190), .A2(n_255), .B1(n_291), .B2(n_307), .C(n_308), .Y(n_189) );
NOR2xp33_ASAP7_75t_SL g190 ( .A(n_191), .B(n_245), .Y(n_190) );
NAND2xp5_ASAP7_75t_L g367 ( .A(n_191), .B(n_368), .Y(n_367) );
INVx1_ASAP7_75t_SL g495 ( .A(n_191), .Y(n_495) );
AND2x2_ASAP7_75t_L g191 ( .A(n_192), .B(n_218), .Y(n_191) );
INVx1_ASAP7_75t_L g335 ( .A(n_192), .Y(n_335) );
AND2x2_ASAP7_75t_L g337 ( .A(n_192), .B(n_236), .Y(n_337) );
AND2x2_ASAP7_75t_L g347 ( .A(n_192), .B(n_235), .Y(n_347) );
HB1xp67_ASAP7_75t_L g365 ( .A(n_192), .Y(n_365) );
INVx1_ASAP7_75t_L g375 ( .A(n_192), .Y(n_375) );
OR2x2_ASAP7_75t_L g413 ( .A(n_192), .B(n_312), .Y(n_413) );
INVx2_ASAP7_75t_L g463 ( .A(n_192), .Y(n_463) );
NAND2xp5_ASAP7_75t_L g480 ( .A(n_192), .B(n_311), .Y(n_480) );
OA21x2_ASAP7_75t_L g192 ( .A1(n_193), .A2(n_198), .B(n_217), .Y(n_192) );
OA21x2_ASAP7_75t_L g221 ( .A1(n_193), .A2(n_222), .B(n_234), .Y(n_221) );
INVx2_ASAP7_75t_L g254 ( .A(n_193), .Y(n_254) );
AND2x2_ASAP7_75t_SL g193 ( .A(n_194), .B(n_195), .Y(n_193) );
AND2x2_ASAP7_75t_L g242 ( .A(n_194), .B(n_195), .Y(n_242) );
NAND2xp5_ASAP7_75t_L g195 ( .A(n_196), .B(n_197), .Y(n_195) );
OAI21xp5_ASAP7_75t_L g198 ( .A1(n_199), .A2(n_210), .B(n_216), .Y(n_198) );
AOI21xp5_ASAP7_75t_L g199 ( .A1(n_200), .A2(n_204), .B(n_207), .Y(n_199) );
INVx3_ASAP7_75t_L g224 ( .A(n_201), .Y(n_224) );
BUFx6f_ASAP7_75t_L g201 ( .A(n_202), .Y(n_201) );
INVx1_ASAP7_75t_L g213 ( .A(n_202), .Y(n_213) );
BUFx3_ASAP7_75t_L g252 ( .A(n_202), .Y(n_252) );
INVx2_ASAP7_75t_L g202 ( .A(n_203), .Y(n_202) );
INVx1_ASAP7_75t_L g206 ( .A(n_203), .Y(n_206) );
INVx1_ASAP7_75t_L g276 ( .A(n_203), .Y(n_276) );
INVx2_ASAP7_75t_L g283 ( .A(n_205), .Y(n_283) );
INVx3_ASAP7_75t_L g205 ( .A(n_206), .Y(n_205) );
INVx1_ASAP7_75t_L g207 ( .A(n_208), .Y(n_207) );
INVx1_ASAP7_75t_L g208 ( .A(n_209), .Y(n_208) );
BUFx6f_ASAP7_75t_L g215 ( .A(n_209), .Y(n_215) );
INVx3_ASAP7_75t_L g228 ( .A(n_209), .Y(n_228) );
BUFx6f_ASAP7_75t_L g233 ( .A(n_209), .Y(n_233) );
AOI21xp5_ASAP7_75t_L g210 ( .A1(n_211), .A2(n_212), .B(n_214), .Y(n_210) );
O2A1O1Ixp5_ASAP7_75t_L g299 ( .A1(n_214), .A2(n_287), .B(n_300), .C(n_301), .Y(n_299) );
INVx2_ASAP7_75t_L g214 ( .A(n_215), .Y(n_214) );
OAI22xp5_ASAP7_75t_L g237 ( .A1(n_215), .A2(n_238), .B1(n_239), .B2(n_240), .Y(n_237) );
OAI22xp5_ASAP7_75t_SL g250 ( .A1(n_215), .A2(n_228), .B1(n_251), .B2(n_253), .Y(n_250) );
OAI22xp5_ASAP7_75t_L g262 ( .A1(n_215), .A2(n_239), .B1(n_263), .B2(n_264), .Y(n_262) );
OAI21xp5_ASAP7_75t_L g222 ( .A1(n_216), .A2(n_223), .B(n_229), .Y(n_222) );
BUFx3_ASAP7_75t_L g243 ( .A(n_216), .Y(n_243) );
OAI21xp5_ASAP7_75t_L g268 ( .A1(n_216), .A2(n_269), .B(n_272), .Y(n_268) );
OAI21xp5_ASAP7_75t_L g280 ( .A1(n_216), .A2(n_281), .B(n_286), .Y(n_280) );
INVx4_ASAP7_75t_SL g502 ( .A(n_216), .Y(n_502) );
NOR2xp67_ASAP7_75t_L g218 ( .A(n_219), .B(n_235), .Y(n_218) );
INVx1_ASAP7_75t_L g219 ( .A(n_220), .Y(n_219) );
HB1xp67_ASAP7_75t_L g329 ( .A(n_220), .Y(n_329) );
NAND2xp5_ASAP7_75t_L g345 ( .A(n_220), .B(n_346), .Y(n_345) );
AND2x2_ASAP7_75t_SL g395 ( .A(n_220), .B(n_335), .Y(n_395) );
INVx2_ASAP7_75t_L g220 ( .A(n_221), .Y(n_220) );
HB1xp67_ASAP7_75t_L g247 ( .A(n_221), .Y(n_247) );
INVx2_ASAP7_75t_L g312 ( .A(n_221), .Y(n_312) );
OR2x2_ASAP7_75t_L g374 ( .A(n_221), .B(n_375), .Y(n_374) );
O2A1O1Ixp5_ASAP7_75t_SL g223 ( .A1(n_224), .A2(n_225), .B(n_226), .C(n_227), .Y(n_223) );
INVx2_ASAP7_75t_L g239 ( .A(n_227), .Y(n_239) );
AOI21xp5_ASAP7_75t_L g269 ( .A1(n_227), .A2(n_270), .B(n_271), .Y(n_269) );
AOI21xp5_ASAP7_75t_L g296 ( .A1(n_227), .A2(n_297), .B(n_298), .Y(n_296) );
INVx5_ASAP7_75t_L g227 ( .A(n_228), .Y(n_227) );
AOI21xp5_ASAP7_75t_L g229 ( .A1(n_230), .A2(n_231), .B(n_232), .Y(n_229) );
INVx1_ASAP7_75t_L g285 ( .A(n_232), .Y(n_285) );
INVx4_ASAP7_75t_L g232 ( .A(n_233), .Y(n_232) );
INVx2_ASAP7_75t_L g500 ( .A(n_233), .Y(n_500) );
AND2x2_ASAP7_75t_L g313 ( .A(n_235), .B(n_249), .Y(n_313) );
AND2x2_ASAP7_75t_L g330 ( .A(n_235), .B(n_310), .Y(n_330) );
INVx2_ASAP7_75t_L g235 ( .A(n_236), .Y(n_235) );
AND2x2_ASAP7_75t_L g248 ( .A(n_236), .B(n_249), .Y(n_248) );
BUFx2_ASAP7_75t_L g333 ( .A(n_236), .Y(n_333) );
AND2x2_ASAP7_75t_L g462 ( .A(n_236), .B(n_463), .Y(n_462) );
AOI21xp5_ASAP7_75t_L g272 ( .A1(n_239), .A2(n_273), .B(n_274), .Y(n_272) );
O2A1O1Ixp33_ASAP7_75t_L g286 ( .A1(n_239), .A2(n_287), .B(n_288), .C(n_289), .Y(n_286) );
INVx2_ASAP7_75t_L g279 ( .A(n_241), .Y(n_279) );
INVx1_ASAP7_75t_L g241 ( .A(n_242), .Y(n_241) );
BUFx6f_ASAP7_75t_L g244 ( .A(n_242), .Y(n_244) );
NAND3xp33_ASAP7_75t_L g261 ( .A(n_243), .B(n_262), .C(n_265), .Y(n_261) );
OAI21xp5_ASAP7_75t_L g295 ( .A1(n_243), .A2(n_296), .B(n_299), .Y(n_295) );
INVx4_ASAP7_75t_L g265 ( .A(n_244), .Y(n_265) );
OA21x2_ASAP7_75t_L g267 ( .A1(n_244), .A2(n_268), .B(n_277), .Y(n_267) );
INVx1_ASAP7_75t_L g307 ( .A(n_245), .Y(n_307) );
AND2x2_ASAP7_75t_L g245 ( .A(n_246), .B(n_248), .Y(n_245) );
AND2x2_ASAP7_75t_L g425 ( .A(n_246), .B(n_313), .Y(n_425) );
INVx1_ASAP7_75t_L g246 ( .A(n_247), .Y(n_246) );
AND2x2_ASAP7_75t_L g426 ( .A(n_247), .B(n_337), .Y(n_426) );
O2A1O1Ixp33_ASAP7_75t_L g393 ( .A1(n_248), .A2(n_394), .B(n_396), .C(n_398), .Y(n_393) );
NAND2xp5_ASAP7_75t_L g403 ( .A(n_248), .B(n_394), .Y(n_403) );
AOI221xp5_ASAP7_75t_L g466 ( .A1(n_248), .A2(n_324), .B1(n_467), .B2(n_468), .C(n_470), .Y(n_466) );
INVx1_ASAP7_75t_L g310 ( .A(n_249), .Y(n_310) );
INVx1_ASAP7_75t_L g346 ( .A(n_249), .Y(n_346) );
BUFx6f_ASAP7_75t_L g355 ( .A(n_249), .Y(n_355) );
INVx1_ASAP7_75t_SL g255 ( .A(n_256), .Y(n_255) );
AND2x2_ASAP7_75t_L g256 ( .A(n_257), .B(n_266), .Y(n_256) );
AND2x2_ASAP7_75t_L g372 ( .A(n_257), .B(n_317), .Y(n_372) );
NAND2xp5_ASAP7_75t_L g391 ( .A(n_257), .B(n_392), .Y(n_391) );
INVx2_ASAP7_75t_L g257 ( .A(n_258), .Y(n_257) );
NOR2xp33_ASAP7_75t_L g340 ( .A(n_258), .B(n_341), .Y(n_340) );
OR2x2_ASAP7_75t_L g464 ( .A(n_258), .B(n_465), .Y(n_464) );
INVx1_ASAP7_75t_L g496 ( .A(n_258), .Y(n_496) );
INVx2_ASAP7_75t_L g258 ( .A(n_259), .Y(n_258) );
INVx3_ASAP7_75t_L g326 ( .A(n_259), .Y(n_326) );
AND2x2_ASAP7_75t_L g352 ( .A(n_259), .B(n_306), .Y(n_352) );
NOR2x1_ASAP7_75t_L g361 ( .A(n_259), .B(n_362), .Y(n_361) );
AND2x2_ASAP7_75t_L g368 ( .A(n_259), .B(n_369), .Y(n_368) );
AND2x4_ASAP7_75t_L g259 ( .A(n_260), .B(n_261), .Y(n_259) );
INVx1_ASAP7_75t_L g304 ( .A(n_260), .Y(n_304) );
AO21x1_ASAP7_75t_L g303 ( .A1(n_262), .A2(n_265), .B(n_304), .Y(n_303) );
NAND2xp5_ASAP7_75t_L g443 ( .A(n_266), .B(n_408), .Y(n_443) );
INVx1_ASAP7_75t_SL g447 ( .A(n_266), .Y(n_447) );
AND2x2_ASAP7_75t_L g266 ( .A(n_267), .B(n_278), .Y(n_266) );
INVx3_ASAP7_75t_L g306 ( .A(n_267), .Y(n_306) );
AND2x2_ASAP7_75t_L g317 ( .A(n_267), .B(n_294), .Y(n_317) );
AND2x2_ASAP7_75t_L g339 ( .A(n_267), .B(n_340), .Y(n_339) );
AND2x2_ASAP7_75t_L g384 ( .A(n_267), .B(n_378), .Y(n_384) );
NAND2xp5_ASAP7_75t_L g465 ( .A(n_267), .B(n_316), .Y(n_465) );
INVx2_ASAP7_75t_L g287 ( .A(n_275), .Y(n_287) );
INVx1_ASAP7_75t_L g275 ( .A(n_276), .Y(n_275) );
AND2x2_ASAP7_75t_L g305 ( .A(n_278), .B(n_306), .Y(n_305) );
INVx2_ASAP7_75t_L g316 ( .A(n_278), .Y(n_316) );
NAND2xp5_ASAP7_75t_L g341 ( .A(n_278), .B(n_294), .Y(n_341) );
AND2x2_ASAP7_75t_L g377 ( .A(n_278), .B(n_378), .Y(n_377) );
OA21x2_ASAP7_75t_L g278 ( .A1(n_279), .A2(n_280), .B(n_290), .Y(n_278) );
OA21x2_ASAP7_75t_L g294 ( .A1(n_279), .A2(n_295), .B(n_302), .Y(n_294) );
O2A1O1Ixp33_ASAP7_75t_L g281 ( .A1(n_282), .A2(n_283), .B(n_284), .C(n_285), .Y(n_281) );
NOR2xp33_ASAP7_75t_L g501 ( .A(n_287), .B(n_502), .Y(n_501) );
NOR2xp33_ASAP7_75t_L g513 ( .A(n_287), .B(n_514), .Y(n_513) );
INVx1_ASAP7_75t_L g291 ( .A(n_292), .Y(n_291) );
AND2x2_ASAP7_75t_L g292 ( .A(n_293), .B(n_305), .Y(n_292) );
INVx1_ASAP7_75t_L g357 ( .A(n_293), .Y(n_357) );
AND2x2_ASAP7_75t_L g399 ( .A(n_293), .B(n_400), .Y(n_399) );
NAND2xp5_ASAP7_75t_SL g405 ( .A(n_293), .B(n_320), .Y(n_405) );
AOI21xp5_ASAP7_75t_SL g479 ( .A1(n_293), .A2(n_311), .B(n_334), .Y(n_479) );
AND2x2_ASAP7_75t_L g293 ( .A(n_294), .B(n_303), .Y(n_293) );
OR2x2_ASAP7_75t_L g322 ( .A(n_294), .B(n_303), .Y(n_322) );
AND2x2_ASAP7_75t_L g369 ( .A(n_294), .B(n_306), .Y(n_369) );
INVx2_ASAP7_75t_L g378 ( .A(n_294), .Y(n_378) );
INVx1_ASAP7_75t_L g484 ( .A(n_294), .Y(n_484) );
AND2x2_ASAP7_75t_L g408 ( .A(n_303), .B(n_378), .Y(n_408) );
INVx1_ASAP7_75t_L g433 ( .A(n_303), .Y(n_433) );
AND2x2_ASAP7_75t_L g342 ( .A(n_305), .B(n_326), .Y(n_342) );
AND2x2_ASAP7_75t_L g354 ( .A(n_305), .B(n_355), .Y(n_354) );
INVx2_ASAP7_75t_SL g472 ( .A(n_305), .Y(n_472) );
INVx2_ASAP7_75t_L g362 ( .A(n_306), .Y(n_362) );
AND2x2_ASAP7_75t_L g400 ( .A(n_306), .B(n_316), .Y(n_400) );
NAND2xp5_ASAP7_75t_L g483 ( .A(n_306), .B(n_484), .Y(n_483) );
OAI21xp33_ASAP7_75t_L g308 ( .A1(n_309), .A2(n_313), .B(n_314), .Y(n_308) );
AND2x2_ASAP7_75t_L g415 ( .A(n_309), .B(n_416), .Y(n_415) );
INVx1_ASAP7_75t_L g469 ( .A(n_309), .Y(n_469) );
AND2x2_ASAP7_75t_L g309 ( .A(n_310), .B(n_311), .Y(n_309) );
INVx1_ASAP7_75t_L g389 ( .A(n_310), .Y(n_389) );
BUFx2_ASAP7_75t_L g488 ( .A(n_310), .Y(n_488) );
BUFx2_ASAP7_75t_L g359 ( .A(n_311), .Y(n_359) );
AND2x2_ASAP7_75t_L g461 ( .A(n_311), .B(n_462), .Y(n_461) );
INVx2_ASAP7_75t_L g311 ( .A(n_312), .Y(n_311) );
INVx1_ASAP7_75t_L g444 ( .A(n_312), .Y(n_444) );
AND2x4_ASAP7_75t_L g371 ( .A(n_313), .B(n_334), .Y(n_371) );
NAND2xp5_ASAP7_75t_SL g407 ( .A(n_313), .B(n_395), .Y(n_407) );
AOI32xp33_ASAP7_75t_L g331 ( .A1(n_314), .A2(n_332), .A3(n_334), .B1(n_336), .B2(n_337), .Y(n_331) );
AND2x2_ASAP7_75t_L g314 ( .A(n_315), .B(n_317), .Y(n_314) );
INVx3_ASAP7_75t_L g320 ( .A(n_315), .Y(n_320) );
OR2x2_ASAP7_75t_L g456 ( .A(n_315), .B(n_412), .Y(n_456) );
INVx2_ASAP7_75t_L g315 ( .A(n_316), .Y(n_315) );
AND2x2_ASAP7_75t_L g325 ( .A(n_316), .B(n_326), .Y(n_325) );
AND2x2_ASAP7_75t_L g432 ( .A(n_316), .B(n_433), .Y(n_432) );
AND2x2_ASAP7_75t_L g324 ( .A(n_317), .B(n_325), .Y(n_324) );
AND2x2_ASAP7_75t_L g336 ( .A(n_317), .B(n_326), .Y(n_336) );
INVx1_ASAP7_75t_L g457 ( .A(n_317), .Y(n_457) );
NAND2xp5_ASAP7_75t_L g490 ( .A(n_317), .B(n_432), .Y(n_490) );
A2O1A1Ixp33_ASAP7_75t_L g318 ( .A1(n_319), .A2(n_323), .B(n_327), .C(n_331), .Y(n_318) );
OAI322xp33_ASAP7_75t_L g427 ( .A1(n_319), .A2(n_364), .A3(n_428), .B1(n_430), .B2(n_434), .C1(n_435), .C2(n_439), .Y(n_427) );
NAND2xp5_ASAP7_75t_L g319 ( .A(n_320), .B(n_321), .Y(n_319) );
INVxp67_ASAP7_75t_L g392 ( .A(n_320), .Y(n_392) );
INVx1_ASAP7_75t_SL g321 ( .A(n_322), .Y(n_321) );
OR2x2_ASAP7_75t_L g446 ( .A(n_322), .B(n_447), .Y(n_446) );
NOR2xp33_ASAP7_75t_L g493 ( .A(n_322), .B(n_362), .Y(n_493) );
INVxp67_ASAP7_75t_L g323 ( .A(n_324), .Y(n_323) );
INVx1_ASAP7_75t_L g385 ( .A(n_325), .Y(n_385) );
OR2x2_ASAP7_75t_L g471 ( .A(n_326), .B(n_472), .Y(n_471) );
INVx1_ASAP7_75t_L g327 ( .A(n_328), .Y(n_327) );
AND2x2_ASAP7_75t_L g328 ( .A(n_329), .B(n_330), .Y(n_328) );
NAND2xp5_ASAP7_75t_L g387 ( .A(n_329), .B(n_388), .Y(n_387) );
AND2x2_ASAP7_75t_L g380 ( .A(n_330), .B(n_359), .Y(n_380) );
AND2x2_ASAP7_75t_L g451 ( .A(n_330), .B(n_364), .Y(n_451) );
NAND2xp5_ASAP7_75t_L g473 ( .A(n_330), .B(n_438), .Y(n_473) );
AOI221xp5_ASAP7_75t_L g338 ( .A1(n_332), .A2(n_339), .B1(n_342), .B2(n_343), .C(n_348), .Y(n_338) );
OR2x2_ASAP7_75t_L g349 ( .A(n_332), .B(n_345), .Y(n_349) );
AND2x2_ASAP7_75t_L g437 ( .A(n_332), .B(n_438), .Y(n_437) );
AOI32xp33_ASAP7_75t_L g476 ( .A1(n_332), .A2(n_362), .A3(n_477), .B1(n_478), .B2(n_481), .Y(n_476) );
INVx2_ASAP7_75t_L g332 ( .A(n_333), .Y(n_332) );
NAND3xp33_ASAP7_75t_L g410 ( .A(n_333), .B(n_369), .C(n_392), .Y(n_410) );
AND2x2_ASAP7_75t_L g436 ( .A(n_333), .B(n_429), .Y(n_436) );
INVxp67_ASAP7_75t_L g416 ( .A(n_334), .Y(n_416) );
BUFx3_ASAP7_75t_L g334 ( .A(n_335), .Y(n_334) );
NAND2xp5_ASAP7_75t_SL g445 ( .A(n_337), .B(n_389), .Y(n_445) );
INVx2_ASAP7_75t_L g455 ( .A(n_337), .Y(n_455) );
NOR2xp33_ASAP7_75t_L g468 ( .A(n_337), .B(n_469), .Y(n_468) );
INVx1_ASAP7_75t_L g424 ( .A(n_340), .Y(n_424) );
OR2x2_ASAP7_75t_L g350 ( .A(n_341), .B(n_351), .Y(n_350) );
NOR2xp33_ASAP7_75t_L g460 ( .A(n_343), .B(n_461), .Y(n_460) );
AND2x2_ASAP7_75t_L g343 ( .A(n_344), .B(n_347), .Y(n_343) );
INVx1_ASAP7_75t_SL g344 ( .A(n_345), .Y(n_344) );
HB1xp67_ASAP7_75t_L g429 ( .A(n_346), .Y(n_429) );
AND2x2_ASAP7_75t_L g388 ( .A(n_347), .B(n_389), .Y(n_388) );
INVx1_ASAP7_75t_L g434 ( .A(n_347), .Y(n_434) );
HB1xp67_ASAP7_75t_L g459 ( .A(n_347), .Y(n_459) );
NOR2xp33_ASAP7_75t_L g348 ( .A(n_349), .B(n_350), .Y(n_348) );
AOI21xp33_ASAP7_75t_SL g373 ( .A1(n_349), .A2(n_374), .B(n_376), .Y(n_373) );
INVx1_ASAP7_75t_L g351 ( .A(n_352), .Y(n_351) );
AND2x2_ASAP7_75t_L g467 ( .A(n_352), .B(n_377), .Y(n_467) );
AOI211xp5_ASAP7_75t_L g353 ( .A1(n_354), .A2(n_356), .B(n_366), .C(n_373), .Y(n_353) );
AND2x2_ASAP7_75t_L g397 ( .A(n_355), .B(n_365), .Y(n_397) );
INVx2_ASAP7_75t_L g412 ( .A(n_355), .Y(n_412) );
OR2x2_ASAP7_75t_L g450 ( .A(n_355), .B(n_413), .Y(n_450) );
NAND2xp5_ASAP7_75t_L g492 ( .A(n_355), .B(n_493), .Y(n_492) );
AOI211xp5_ASAP7_75t_SL g356 ( .A1(n_357), .A2(n_358), .B(n_360), .C(n_363), .Y(n_356) );
INVxp67_ASAP7_75t_L g358 ( .A(n_359), .Y(n_358) );
NAND2xp5_ASAP7_75t_L g396 ( .A(n_359), .B(n_397), .Y(n_396) );
OAI211xp5_ASAP7_75t_L g478 ( .A1(n_360), .A2(n_455), .B(n_479), .C(n_480), .Y(n_478) );
INVx1_ASAP7_75t_L g360 ( .A(n_361), .Y(n_360) );
NAND2x1p5_ASAP7_75t_L g376 ( .A(n_361), .B(n_377), .Y(n_376) );
AND2x2_ASAP7_75t_L g418 ( .A(n_362), .B(n_408), .Y(n_418) );
INVx1_ASAP7_75t_L g423 ( .A(n_362), .Y(n_423) );
INVx1_ASAP7_75t_L g363 ( .A(n_364), .Y(n_363) );
INVx1_ASAP7_75t_L g364 ( .A(n_365), .Y(n_364) );
NAND2xp5_ASAP7_75t_SL g366 ( .A(n_367), .B(n_370), .Y(n_366) );
INVxp33_ASAP7_75t_L g474 ( .A(n_368), .Y(n_474) );
AND2x2_ASAP7_75t_L g453 ( .A(n_369), .B(n_432), .Y(n_453) );
NAND2xp5_ASAP7_75t_L g370 ( .A(n_371), .B(n_372), .Y(n_370) );
AOI21xp5_ASAP7_75t_L g435 ( .A1(n_374), .A2(n_436), .B(n_437), .Y(n_435) );
OAI322xp33_ASAP7_75t_L g454 ( .A1(n_376), .A2(n_455), .A3(n_456), .B1(n_457), .B2(n_458), .C1(n_460), .C2(n_464), .Y(n_454) );
AOI221xp5_ASAP7_75t_L g379 ( .A1(n_380), .A2(n_381), .B1(n_386), .B2(n_390), .C(n_393), .Y(n_379) );
INVx2_ASAP7_75t_L g381 ( .A(n_382), .Y(n_381) );
OR2x2_ASAP7_75t_L g382 ( .A(n_383), .B(n_385), .Y(n_382) );
INVx1_ASAP7_75t_L g383 ( .A(n_384), .Y(n_383) );
AND2x2_ASAP7_75t_L g431 ( .A(n_384), .B(n_432), .Y(n_431) );
INVx1_ASAP7_75t_L g386 ( .A(n_387), .Y(n_386) );
INVx1_ASAP7_75t_L g475 ( .A(n_388), .Y(n_475) );
INVxp67_ASAP7_75t_L g390 ( .A(n_391), .Y(n_390) );
NOR2xp33_ASAP7_75t_L g477 ( .A(n_391), .B(n_411), .Y(n_477) );
INVx2_ASAP7_75t_L g394 ( .A(n_395), .Y(n_394) );
INVx1_ASAP7_75t_SL g398 ( .A(n_399), .Y(n_398) );
AND2x2_ASAP7_75t_L g440 ( .A(n_400), .B(n_408), .Y(n_440) );
AOI221xp5_ASAP7_75t_L g401 ( .A1(n_402), .A2(n_404), .B1(n_406), .B2(n_408), .C(n_409), .Y(n_401) );
INVx1_ASAP7_75t_L g402 ( .A(n_403), .Y(n_402) );
AOI221xp5_ASAP7_75t_L g420 ( .A1(n_404), .A2(n_421), .B1(n_425), .B2(n_426), .C(n_427), .Y(n_420) );
INVx1_ASAP7_75t_L g404 ( .A(n_405), .Y(n_404) );
INVxp67_ASAP7_75t_L g406 ( .A(n_407), .Y(n_406) );
NAND2xp5_ASAP7_75t_L g422 ( .A(n_408), .B(n_423), .Y(n_422) );
OAI22xp5_ASAP7_75t_L g409 ( .A1(n_410), .A2(n_411), .B1(n_414), .B2(n_417), .Y(n_409) );
OR2x2_ASAP7_75t_L g411 ( .A(n_412), .B(n_413), .Y(n_411) );
INVx2_ASAP7_75t_SL g438 ( .A(n_413), .Y(n_438) );
INVxp67_ASAP7_75t_L g414 ( .A(n_415), .Y(n_414) );
INVx1_ASAP7_75t_L g417 ( .A(n_418), .Y(n_417) );
NAND5xp2_ASAP7_75t_L g419 ( .A(n_420), .B(n_441), .C(n_466), .D(n_476), .E(n_486), .Y(n_419) );
NAND2xp5_ASAP7_75t_SL g421 ( .A(n_422), .B(n_424), .Y(n_421) );
NOR4xp25_ASAP7_75t_L g494 ( .A(n_423), .B(n_429), .C(n_495), .D(n_496), .Y(n_494) );
AOI221xp5_ASAP7_75t_L g486 ( .A1(n_426), .A2(n_487), .B1(n_489), .B2(n_491), .C(n_494), .Y(n_486) );
INVx1_ASAP7_75t_L g428 ( .A(n_429), .Y(n_428) );
INVx1_ASAP7_75t_L g430 ( .A(n_431), .Y(n_430) );
INVx1_ASAP7_75t_L g485 ( .A(n_432), .Y(n_485) );
OAI322xp33_ASAP7_75t_L g442 ( .A1(n_436), .A2(n_443), .A3(n_444), .B1(n_445), .B2(n_446), .C1(n_448), .C2(n_452), .Y(n_442) );
INVx1_ASAP7_75t_SL g439 ( .A(n_440), .Y(n_439) );
NOR2xp33_ASAP7_75t_L g441 ( .A(n_442), .B(n_454), .Y(n_441) );
NOR2xp33_ASAP7_75t_L g448 ( .A(n_449), .B(n_451), .Y(n_448) );
INVx2_ASAP7_75t_L g449 ( .A(n_450), .Y(n_449) );
INVx1_ASAP7_75t_L g452 ( .A(n_453), .Y(n_452) );
INVx1_ASAP7_75t_L g458 ( .A(n_459), .Y(n_458) );
AND2x2_ASAP7_75t_L g487 ( .A(n_462), .B(n_488), .Y(n_487) );
OAI22xp33_ASAP7_75t_L g470 ( .A1(n_471), .A2(n_473), .B1(n_474), .B2(n_475), .Y(n_470) );
INVx1_ASAP7_75t_L g481 ( .A(n_482), .Y(n_481) );
OR2x2_ASAP7_75t_L g482 ( .A(n_483), .B(n_485), .Y(n_482) );
INVx1_ASAP7_75t_L g489 ( .A(n_490), .Y(n_489) );
INVxp67_ASAP7_75t_L g491 ( .A(n_492), .Y(n_491) );
AND2x2_ASAP7_75t_L g497 ( .A(n_498), .B(n_501), .Y(n_497) );
INVx1_ASAP7_75t_L g514 ( .A(n_498), .Y(n_514) );
HB1xp67_ASAP7_75t_L g498 ( .A(n_499), .Y(n_498) );
INVx2_ASAP7_75t_L g499 ( .A(n_500), .Y(n_499) );
OAI322xp33_ASAP7_75t_L g503 ( .A1(n_504), .A2(n_506), .A3(n_510), .B1(n_511), .B2(n_516), .C1(n_517), .C2(n_518), .Y(n_503) );
CKINVDCx20_ASAP7_75t_R g506 ( .A(n_507), .Y(n_506) );
CKINVDCx20_ASAP7_75t_R g507 ( .A(n_508), .Y(n_507) );
CKINVDCx20_ASAP7_75t_R g511 ( .A(n_512), .Y(n_511) );
CKINVDCx20_ASAP7_75t_R g518 ( .A(n_519), .Y(n_518) );
CKINVDCx20_ASAP7_75t_R g519 ( .A(n_520), .Y(n_519) );
endmodule