module fake_jpeg_11700_n_76 (n_3, n_2, n_1, n_0, n_4, n_8, n_6, n_5, n_7, n_76);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_8;
input n_6;
input n_5;
input n_7;

output n_76;

wire n_13;
wire n_21;
wire n_57;
wire n_53;
wire n_33;
wire n_54;
wire n_61;
wire n_45;
wire n_10;
wire n_23;
wire n_69;
wire n_27;
wire n_64;
wire n_55;
wire n_22;
wire n_51;
wire n_47;
wire n_14;
wire n_40;
wire n_73;
wire n_19;
wire n_20;
wire n_18;
wire n_59;
wire n_35;
wire n_48;
wire n_71;
wire n_52;
wire n_68;
wire n_46;
wire n_58;
wire n_41;
wire n_60;
wire n_63;
wire n_65;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_16;
wire n_49;
wire n_72;
wire n_24;
wire n_28;
wire n_38;
wire n_26;
wire n_44;
wire n_9;
wire n_36;
wire n_74;
wire n_11;
wire n_62;
wire n_25;
wire n_17;
wire n_31;
wire n_56;
wire n_67;
wire n_75;
wire n_29;
wire n_43;
wire n_37;
wire n_50;
wire n_12;
wire n_32;
wire n_70;
wire n_15;
wire n_66;

CKINVDCx20_ASAP7_75t_R g9 ( 
.A(n_2),
.Y(n_9)
);

BUFx12f_ASAP7_75t_L g10 ( 
.A(n_7),
.Y(n_10)
);

INVx1_ASAP7_75t_SL g11 ( 
.A(n_6),
.Y(n_11)
);

CKINVDCx20_ASAP7_75t_R g12 ( 
.A(n_1),
.Y(n_12)
);

INVx2_ASAP7_75t_L g13 ( 
.A(n_1),
.Y(n_13)
);

CKINVDCx20_ASAP7_75t_R g14 ( 
.A(n_1),
.Y(n_14)
);

BUFx12_ASAP7_75t_L g15 ( 
.A(n_2),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_5),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_8),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_7),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_0),
.Y(n_19)
);

INVx2_ASAP7_75t_L g20 ( 
.A(n_13),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_20),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_10),
.Y(n_21)
);

CKINVDCx6p67_ASAP7_75t_R g37 ( 
.A(n_21),
.Y(n_37)
);

INVx2_ASAP7_75t_L g22 ( 
.A(n_13),
.Y(n_22)
);

NAND2xp5_ASAP7_75t_SL g39 ( 
.A(n_22),
.B(n_24),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_15),
.Y(n_23)
);

NOR2xp33_ASAP7_75t_L g30 ( 
.A(n_23),
.B(n_25),
.Y(n_30)
);

NOR2xp33_ASAP7_75t_L g24 ( 
.A(n_17),
.B(n_4),
.Y(n_24)
);

OR2x2_ASAP7_75t_L g25 ( 
.A(n_11),
.B(n_0),
.Y(n_25)
);

INVx2_ASAP7_75t_L g26 ( 
.A(n_10),
.Y(n_26)
);

NAND2xp5_ASAP7_75t_L g29 ( 
.A(n_26),
.B(n_10),
.Y(n_29)
);

NOR2xp33_ASAP7_75t_L g27 ( 
.A(n_16),
.B(n_4),
.Y(n_27)
);

NOR2xp33_ASAP7_75t_L g33 ( 
.A(n_27),
.B(n_28),
.Y(n_33)
);

INVx2_ASAP7_75t_L g28 ( 
.A(n_10),
.Y(n_28)
);

AND2x2_ASAP7_75t_L g43 ( 
.A(n_29),
.B(n_11),
.Y(n_43)
);

NAND2xp5_ASAP7_75t_L g31 ( 
.A(n_20),
.B(n_19),
.Y(n_31)
);

NAND2xp5_ASAP7_75t_L g44 ( 
.A(n_31),
.B(n_36),
.Y(n_44)
);

BUFx24_ASAP7_75t_SL g32 ( 
.A(n_25),
.Y(n_32)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_32),
.B(n_38),
.Y(n_50)
);

AOI22xp33_ASAP7_75t_L g35 ( 
.A1(n_22),
.A2(n_19),
.B1(n_14),
.B2(n_12),
.Y(n_35)
);

OAI22xp5_ASAP7_75t_SL g45 ( 
.A1(n_35),
.A2(n_40),
.B1(n_9),
.B2(n_15),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g36 ( 
.A(n_26),
.B(n_18),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g38 ( 
.A(n_21),
.B(n_18),
.Y(n_38)
);

AOI22xp33_ASAP7_75t_L g40 ( 
.A1(n_20),
.A2(n_9),
.B1(n_14),
.B2(n_12),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g41 ( 
.A(n_24),
.B(n_16),
.Y(n_41)
);

INVxp67_ASAP7_75t_L g47 ( 
.A(n_41),
.Y(n_47)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_34),
.Y(n_42)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_42),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_SL g53 ( 
.A(n_43),
.B(n_45),
.Y(n_53)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_31),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_SL g54 ( 
.A(n_46),
.B(n_51),
.Y(n_54)
);

HB1xp67_ASAP7_75t_L g48 ( 
.A(n_34),
.Y(n_48)
);

HB1xp67_ASAP7_75t_L g58 ( 
.A(n_48),
.Y(n_58)
);

XNOR2xp5_ASAP7_75t_L g49 ( 
.A(n_39),
.B(n_15),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_SL g56 ( 
.A(n_49),
.B(n_52),
.Y(n_56)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_33),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_L g52 ( 
.A(n_29),
.B(n_0),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_SL g57 ( 
.A(n_44),
.B(n_30),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_SL g63 ( 
.A(n_57),
.B(n_47),
.Y(n_63)
);

AOI22xp5_ASAP7_75t_L g59 ( 
.A1(n_45),
.A2(n_37),
.B1(n_15),
.B2(n_3),
.Y(n_59)
);

OAI22xp5_ASAP7_75t_L g61 ( 
.A1(n_59),
.A2(n_47),
.B1(n_50),
.B2(n_37),
.Y(n_61)
);

NOR3xp33_ASAP7_75t_L g60 ( 
.A(n_53),
.B(n_43),
.C(n_52),
.Y(n_60)
);

BUFx2_ASAP7_75t_L g65 ( 
.A(n_60),
.Y(n_65)
);

XOR2xp5_ASAP7_75t_L g67 ( 
.A(n_61),
.B(n_64),
.Y(n_67)
);

XNOR2xp5_ASAP7_75t_SL g62 ( 
.A(n_56),
.B(n_49),
.Y(n_62)
);

XNOR2xp5_ASAP7_75t_SL g68 ( 
.A(n_62),
.B(n_63),
.Y(n_68)
);

XNOR2xp5_ASAP7_75t_SL g64 ( 
.A(n_54),
.B(n_43),
.Y(n_64)
);

OAI21xp33_ASAP7_75t_SL g66 ( 
.A1(n_60),
.A2(n_59),
.B(n_58),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_L g69 ( 
.A(n_66),
.B(n_55),
.Y(n_69)
);

MAJIxp5_ASAP7_75t_L g71 ( 
.A(n_69),
.B(n_70),
.C(n_67),
.Y(n_71)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_66),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_SL g73 ( 
.A(n_71),
.B(n_72),
.Y(n_73)
);

MAJIxp5_ASAP7_75t_L g72 ( 
.A(n_70),
.B(n_68),
.C(n_65),
.Y(n_72)
);

MAJIxp5_ASAP7_75t_L g74 ( 
.A(n_73),
.B(n_55),
.C(n_5),
.Y(n_74)
);

OAI21xp5_ASAP7_75t_SL g75 ( 
.A1(n_74),
.A2(n_6),
.B(n_8),
.Y(n_75)
);

XOR2xp5_ASAP7_75t_L g76 ( 
.A(n_75),
.B(n_2),
.Y(n_76)
);


endmodule