module fake_jpeg_22253_n_44 (n_13, n_1, n_10, n_6, n_14, n_19, n_18, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_44);

input n_13;
input n_1;
input n_10;
input n_6;
input n_14;
input n_19;
input n_18;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_44;

wire n_21;
wire n_33;
wire n_23;
wire n_27;
wire n_22;
wire n_40;
wire n_20;
wire n_35;
wire n_41;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_24;
wire n_28;
wire n_38;
wire n_26;
wire n_36;
wire n_25;
wire n_31;
wire n_29;
wire n_37;
wire n_43;
wire n_32;

INVx5_ASAP7_75t_L g20 ( 
.A(n_13),
.Y(n_20)
);

BUFx10_ASAP7_75t_L g21 ( 
.A(n_15),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_1),
.Y(n_22)
);

INVx4_ASAP7_75t_L g23 ( 
.A(n_19),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_16),
.Y(n_24)
);

AOI21xp33_ASAP7_75t_L g25 ( 
.A1(n_21),
.A2(n_0),
.B(n_1),
.Y(n_25)
);

OAI22xp5_ASAP7_75t_SL g34 ( 
.A1(n_25),
.A2(n_27),
.B1(n_4),
.B2(n_5),
.Y(n_34)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_23),
.Y(n_26)
);

NOR2xp33_ASAP7_75t_L g30 ( 
.A(n_26),
.B(n_29),
.Y(n_30)
);

AOI22xp5_ASAP7_75t_SL g27 ( 
.A1(n_22),
.A2(n_0),
.B1(n_2),
.B2(n_3),
.Y(n_27)
);

NAND2xp5_ASAP7_75t_SL g28 ( 
.A(n_22),
.B(n_2),
.Y(n_28)
);

NAND2xp5_ASAP7_75t_L g31 ( 
.A(n_28),
.B(n_4),
.Y(n_31)
);

NOR2xp33_ASAP7_75t_L g29 ( 
.A(n_23),
.B(n_3),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_31),
.Y(n_37)
);

AOI22xp5_ASAP7_75t_L g32 ( 
.A1(n_27),
.A2(n_20),
.B1(n_24),
.B2(n_21),
.Y(n_32)
);

OAI22xp5_ASAP7_75t_SL g36 ( 
.A1(n_32),
.A2(n_33),
.B1(n_35),
.B2(n_21),
.Y(n_36)
);

OAI22xp5_ASAP7_75t_SL g33 ( 
.A1(n_25),
.A2(n_20),
.B1(n_24),
.B2(n_12),
.Y(n_33)
);

XNOR2xp5_ASAP7_75t_L g38 ( 
.A(n_34),
.B(n_5),
.Y(n_38)
);

OAI22xp5_ASAP7_75t_SL g35 ( 
.A1(n_25),
.A2(n_24),
.B1(n_14),
.B2(n_7),
.Y(n_35)
);

AOI22xp5_ASAP7_75t_SL g40 ( 
.A1(n_36),
.A2(n_30),
.B1(n_21),
.B2(n_6),
.Y(n_40)
);

OAI22xp5_ASAP7_75t_SL g39 ( 
.A1(n_38),
.A2(n_32),
.B1(n_37),
.B2(n_33),
.Y(n_39)
);

NOR2xp67_ASAP7_75t_L g41 ( 
.A(n_39),
.B(n_40),
.Y(n_41)
);

A2O1A1Ixp33_ASAP7_75t_L g42 ( 
.A1(n_41),
.A2(n_38),
.B(n_6),
.C(n_9),
.Y(n_42)
);

AOI21xp5_ASAP7_75t_SL g43 ( 
.A1(n_42),
.A2(n_8),
.B(n_10),
.Y(n_43)
);

OAI22xp5_ASAP7_75t_SL g44 ( 
.A1(n_43),
.A2(n_11),
.B1(n_17),
.B2(n_18),
.Y(n_44)
);


endmodule