module fake_jpeg_9119_n_252 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_252);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_252;

wire n_159;
wire n_117;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_84;
wire n_59;
wire n_98;
wire n_251;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_223;
wire n_234;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_44;
wire n_24;
wire n_143;
wire n_202;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_217;
wire n_216;
wire n_184;
wire n_53;
wire n_91;
wire n_54;
wire n_93;
wire n_33;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_118;
wire n_140;
wire n_82;
wire n_128;
wire n_100;
wire n_96;

INVx1_ASAP7_75t_L g17 ( 
.A(n_11),
.Y(n_17)
);

BUFx12f_ASAP7_75t_L g18 ( 
.A(n_5),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_14),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_12),
.Y(n_20)
);

BUFx12_ASAP7_75t_L g21 ( 
.A(n_4),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_10),
.Y(n_22)
);

BUFx16f_ASAP7_75t_L g23 ( 
.A(n_14),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_16),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_4),
.Y(n_25)
);

INVx11_ASAP7_75t_L g26 ( 
.A(n_0),
.Y(n_26)
);

BUFx3_ASAP7_75t_L g27 ( 
.A(n_15),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_4),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_0),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_1),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_8),
.Y(n_31)
);

INVx11_ASAP7_75t_SL g32 ( 
.A(n_6),
.Y(n_32)
);

INVx11_ASAP7_75t_SL g33 ( 
.A(n_1),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_7),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_L g35 ( 
.A(n_25),
.B(n_0),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_SL g55 ( 
.A(n_35),
.B(n_36),
.Y(n_55)
);

OR2x2_ASAP7_75t_L g36 ( 
.A(n_25),
.B(n_1),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_18),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_37),
.Y(n_48)
);

INVx5_ASAP7_75t_L g38 ( 
.A(n_23),
.Y(n_38)
);

INVx2_ASAP7_75t_L g52 ( 
.A(n_38),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_18),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_39),
.Y(n_49)
);

BUFx12f_ASAP7_75t_L g40 ( 
.A(n_23),
.Y(n_40)
);

INVx4_ASAP7_75t_L g65 ( 
.A(n_40),
.Y(n_65)
);

AOI22xp33_ASAP7_75t_SL g41 ( 
.A1(n_26),
.A2(n_2),
.B1(n_3),
.B2(n_5),
.Y(n_41)
);

OAI22xp33_ASAP7_75t_SL g56 ( 
.A1(n_41),
.A2(n_17),
.B1(n_29),
.B2(n_30),
.Y(n_56)
);

BUFx5_ASAP7_75t_L g42 ( 
.A(n_23),
.Y(n_42)
);

BUFx3_ASAP7_75t_L g51 ( 
.A(n_42),
.Y(n_51)
);

INVx3_ASAP7_75t_L g43 ( 
.A(n_22),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g47 ( 
.A(n_43),
.B(n_44),
.Y(n_47)
);

INVx6_ASAP7_75t_SL g44 ( 
.A(n_23),
.Y(n_44)
);

INVx4_ASAP7_75t_SL g45 ( 
.A(n_23),
.Y(n_45)
);

OR2x2_ASAP7_75t_L g57 ( 
.A(n_45),
.B(n_21),
.Y(n_57)
);

AOI22xp33_ASAP7_75t_SL g46 ( 
.A1(n_43),
.A2(n_26),
.B1(n_17),
.B2(n_29),
.Y(n_46)
);

AOI22xp33_ASAP7_75t_SL g70 ( 
.A1(n_46),
.A2(n_56),
.B1(n_62),
.B2(n_67),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_SL g50 ( 
.A(n_36),
.B(n_17),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_SL g98 ( 
.A(n_50),
.B(n_66),
.Y(n_98)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_40),
.Y(n_53)
);

INVx6_ASAP7_75t_L g100 ( 
.A(n_53),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_L g54 ( 
.A(n_36),
.B(n_18),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_L g75 ( 
.A(n_54),
.B(n_58),
.Y(n_75)
);

BUFx2_ASAP7_75t_SL g72 ( 
.A(n_57),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_L g58 ( 
.A(n_35),
.B(n_18),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_40),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g76 ( 
.A(n_59),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_L g60 ( 
.A(n_37),
.B(n_18),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_L g77 ( 
.A(n_60),
.B(n_64),
.Y(n_77)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_40),
.Y(n_61)
);

INVx5_ASAP7_75t_L g69 ( 
.A(n_61),
.Y(n_69)
);

AOI22xp33_ASAP7_75t_SL g62 ( 
.A1(n_43),
.A2(n_26),
.B1(n_30),
.B2(n_29),
.Y(n_62)
);

INVx2_ASAP7_75t_L g63 ( 
.A(n_38),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_63),
.B(n_40),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_L g64 ( 
.A(n_37),
.B(n_18),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_38),
.B(n_30),
.Y(n_66)
);

AOI22xp33_ASAP7_75t_SL g67 ( 
.A1(n_45),
.A2(n_34),
.B1(n_25),
.B2(n_19),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_SL g68 ( 
.A(n_41),
.B(n_31),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_SL g99 ( 
.A(n_68),
.B(n_2),
.Y(n_99)
);

OAI21xp5_ASAP7_75t_SL g71 ( 
.A1(n_54),
.A2(n_42),
.B(n_44),
.Y(n_71)
);

MAJIxp5_ASAP7_75t_L g124 ( 
.A(n_71),
.B(n_87),
.C(n_32),
.Y(n_124)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_73),
.Y(n_105)
);

CKINVDCx16_ASAP7_75t_R g74 ( 
.A(n_66),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_74),
.B(n_82),
.Y(n_102)
);

INVxp67_ASAP7_75t_L g78 ( 
.A(n_47),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_SL g103 ( 
.A(n_78),
.B(n_80),
.Y(n_103)
);

AOI22xp33_ASAP7_75t_L g79 ( 
.A1(n_68),
.A2(n_34),
.B1(n_19),
.B2(n_31),
.Y(n_79)
);

OAI22xp5_ASAP7_75t_SL g121 ( 
.A1(n_79),
.A2(n_85),
.B1(n_94),
.B2(n_96),
.Y(n_121)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_47),
.Y(n_80)
);

OAI21xp33_ASAP7_75t_L g81 ( 
.A1(n_50),
.A2(n_42),
.B(n_3),
.Y(n_81)
);

OAI21xp5_ASAP7_75t_L g113 ( 
.A1(n_81),
.A2(n_99),
.B(n_2),
.Y(n_113)
);

INVx2_ASAP7_75t_L g82 ( 
.A(n_48),
.Y(n_82)
);

AOI22xp33_ASAP7_75t_SL g83 ( 
.A1(n_52),
.A2(n_34),
.B1(n_45),
.B2(n_28),
.Y(n_83)
);

INVxp67_ASAP7_75t_L g104 ( 
.A(n_83),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_58),
.B(n_28),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_SL g114 ( 
.A(n_84),
.B(n_86),
.Y(n_114)
);

AOI22xp33_ASAP7_75t_L g85 ( 
.A1(n_60),
.A2(n_24),
.B1(n_20),
.B2(n_45),
.Y(n_85)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_64),
.Y(n_86)
);

XNOR2xp5_ASAP7_75t_L g87 ( 
.A(n_55),
.B(n_57),
.Y(n_87)
);

AOI22xp33_ASAP7_75t_SL g88 ( 
.A1(n_52),
.A2(n_24),
.B1(n_20),
.B2(n_22),
.Y(n_88)
);

CKINVDCx16_ASAP7_75t_R g108 ( 
.A(n_88),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_63),
.B(n_21),
.Y(n_89)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_89),
.Y(n_110)
);

INVx5_ASAP7_75t_L g90 ( 
.A(n_48),
.Y(n_90)
);

INVx2_ASAP7_75t_L g126 ( 
.A(n_90),
.Y(n_126)
);

INVxp67_ASAP7_75t_L g91 ( 
.A(n_51),
.Y(n_91)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_91),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_65),
.B(n_21),
.Y(n_92)
);

CKINVDCx20_ASAP7_75t_R g107 ( 
.A(n_92),
.Y(n_107)
);

OA22x2_ASAP7_75t_L g93 ( 
.A1(n_57),
.A2(n_39),
.B1(n_22),
.B2(n_27),
.Y(n_93)
);

AOI22xp5_ASAP7_75t_L g122 ( 
.A1(n_93),
.A2(n_49),
.B1(n_33),
.B2(n_32),
.Y(n_122)
);

AOI22xp5_ASAP7_75t_L g94 ( 
.A1(n_55),
.A2(n_22),
.B1(n_27),
.B2(n_39),
.Y(n_94)
);

CKINVDCx16_ASAP7_75t_R g95 ( 
.A(n_51),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_SL g115 ( 
.A(n_95),
.B(n_97),
.Y(n_115)
);

AOI22xp5_ASAP7_75t_L g96 ( 
.A1(n_65),
.A2(n_27),
.B1(n_21),
.B2(n_33),
.Y(n_96)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_48),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g101 ( 
.A(n_77),
.B(n_61),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_L g131 ( 
.A(n_101),
.B(n_112),
.Y(n_131)
);

XNOR2xp5_ASAP7_75t_SL g106 ( 
.A(n_75),
.B(n_87),
.Y(n_106)
);

MAJIxp5_ASAP7_75t_L g134 ( 
.A(n_106),
.B(n_118),
.C(n_123),
.Y(n_134)
);

AOI32xp33_ASAP7_75t_L g109 ( 
.A1(n_72),
.A2(n_75),
.A3(n_77),
.B1(n_71),
.B2(n_70),
.Y(n_109)
);

OAI21xp5_ASAP7_75t_SL g136 ( 
.A1(n_109),
.A2(n_93),
.B(n_91),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_L g112 ( 
.A(n_86),
.B(n_61),
.Y(n_112)
);

NOR3xp33_ASAP7_75t_L g143 ( 
.A(n_113),
.B(n_6),
.C(n_7),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_L g116 ( 
.A(n_74),
.B(n_59),
.Y(n_116)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_116),
.Y(n_130)
);

INVx3_ASAP7_75t_L g117 ( 
.A(n_76),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_L g132 ( 
.A(n_117),
.B(n_119),
.Y(n_132)
);

XOR2xp5_ASAP7_75t_L g118 ( 
.A(n_94),
.B(n_21),
.Y(n_118)
);

INVx2_ASAP7_75t_L g119 ( 
.A(n_90),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_L g120 ( 
.A(n_98),
.B(n_59),
.Y(n_120)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_120),
.Y(n_137)
);

OAI22xp5_ASAP7_75t_L g135 ( 
.A1(n_122),
.A2(n_96),
.B1(n_69),
.B2(n_97),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_L g123 ( 
.A(n_98),
.B(n_53),
.Y(n_123)
);

AND2x2_ASAP7_75t_L g145 ( 
.A(n_124),
.B(n_7),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_L g125 ( 
.A(n_99),
.B(n_53),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_L g138 ( 
.A(n_125),
.B(n_95),
.Y(n_138)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_102),
.Y(n_127)
);

AOI22xp33_ASAP7_75t_SL g154 ( 
.A1(n_127),
.A2(n_133),
.B1(n_141),
.B2(n_144),
.Y(n_154)
);

OAI22xp5_ASAP7_75t_SL g128 ( 
.A1(n_109),
.A2(n_78),
.B1(n_80),
.B2(n_93),
.Y(n_128)
);

OAI22xp5_ASAP7_75t_SL g170 ( 
.A1(n_128),
.A2(n_140),
.B1(n_142),
.B2(n_150),
.Y(n_170)
);

INVxp67_ASAP7_75t_L g129 ( 
.A(n_115),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_SL g163 ( 
.A(n_129),
.B(n_147),
.Y(n_163)
);

AOI22xp33_ASAP7_75t_SL g133 ( 
.A1(n_108),
.A2(n_69),
.B1(n_100),
.B2(n_82),
.Y(n_133)
);

CKINVDCx14_ASAP7_75t_R g169 ( 
.A(n_135),
.Y(n_169)
);

MAJIxp5_ASAP7_75t_L g164 ( 
.A(n_136),
.B(n_128),
.C(n_139),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_L g157 ( 
.A(n_138),
.B(n_114),
.Y(n_157)
);

AOI21xp5_ASAP7_75t_L g139 ( 
.A1(n_104),
.A2(n_93),
.B(n_100),
.Y(n_139)
);

OAI21xp5_ASAP7_75t_SL g155 ( 
.A1(n_139),
.A2(n_145),
.B(n_149),
.Y(n_155)
);

AO21x2_ASAP7_75t_L g140 ( 
.A1(n_108),
.A2(n_49),
.B(n_76),
.Y(n_140)
);

AOI22xp33_ASAP7_75t_SL g141 ( 
.A1(n_119),
.A2(n_3),
.B1(n_5),
.B2(n_6),
.Y(n_141)
);

AOI22xp5_ASAP7_75t_L g142 ( 
.A1(n_121),
.A2(n_49),
.B1(n_76),
.B2(n_8),
.Y(n_142)
);

NOR3xp33_ASAP7_75t_L g158 ( 
.A(n_143),
.B(n_148),
.C(n_113),
.Y(n_158)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_112),
.Y(n_144)
);

CKINVDCx16_ASAP7_75t_R g146 ( 
.A(n_115),
.Y(n_146)
);

INVxp67_ASAP7_75t_L g160 ( 
.A(n_146),
.Y(n_160)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_116),
.Y(n_147)
);

NAND3xp33_ASAP7_75t_L g148 ( 
.A(n_120),
.B(n_123),
.C(n_125),
.Y(n_148)
);

OAI21x1_ASAP7_75t_R g149 ( 
.A1(n_126),
.A2(n_16),
.B(n_9),
.Y(n_149)
);

AOI22xp5_ASAP7_75t_L g150 ( 
.A1(n_121),
.A2(n_8),
.B1(n_9),
.B2(n_10),
.Y(n_150)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_103),
.Y(n_151)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_151),
.Y(n_156)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_101),
.Y(n_152)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_152),
.Y(n_161)
);

INVxp67_ASAP7_75t_L g153 ( 
.A(n_122),
.Y(n_153)
);

OAI21xp5_ASAP7_75t_SL g168 ( 
.A1(n_153),
.A2(n_104),
.B(n_111),
.Y(n_168)
);

CKINVDCx16_ASAP7_75t_R g192 ( 
.A(n_157),
.Y(n_192)
);

NOR2xp33_ASAP7_75t_L g180 ( 
.A(n_158),
.B(n_168),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_L g159 ( 
.A(n_131),
.B(n_124),
.Y(n_159)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_159),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_L g162 ( 
.A(n_131),
.B(n_118),
.Y(n_162)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_162),
.Y(n_184)
);

OAI21xp5_ASAP7_75t_L g182 ( 
.A1(n_164),
.A2(n_174),
.B(n_134),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_L g165 ( 
.A(n_137),
.B(n_130),
.Y(n_165)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_165),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_L g166 ( 
.A(n_137),
.B(n_106),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_L g178 ( 
.A(n_166),
.B(n_172),
.Y(n_178)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_132),
.Y(n_167)
);

NOR2xp33_ASAP7_75t_L g194 ( 
.A(n_167),
.B(n_171),
.Y(n_194)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_142),
.Y(n_171)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_140),
.Y(n_172)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_140),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_L g187 ( 
.A(n_173),
.B(n_175),
.Y(n_187)
);

XOR2x1_ASAP7_75t_L g174 ( 
.A(n_136),
.B(n_140),
.Y(n_174)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_140),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_L g176 ( 
.A(n_130),
.B(n_129),
.Y(n_176)
);

NOR2xp33_ASAP7_75t_L g188 ( 
.A(n_176),
.B(n_105),
.Y(n_188)
);

INVxp67_ASAP7_75t_L g177 ( 
.A(n_149),
.Y(n_177)
);

INVx1_ASAP7_75t_SL g190 ( 
.A(n_177),
.Y(n_190)
);

MAJIxp5_ASAP7_75t_L g181 ( 
.A(n_166),
.B(n_134),
.C(n_107),
.Y(n_181)
);

XOR2xp5_ASAP7_75t_L g209 ( 
.A(n_181),
.B(n_186),
.Y(n_209)
);

OAI21xp5_ASAP7_75t_SL g205 ( 
.A1(n_182),
.A2(n_170),
.B(n_155),
.Y(n_205)
);

BUFx3_ASAP7_75t_L g183 ( 
.A(n_174),
.Y(n_183)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_183),
.Y(n_211)
);

OAI22xp5_ASAP7_75t_SL g185 ( 
.A1(n_172),
.A2(n_150),
.B1(n_153),
.B2(n_107),
.Y(n_185)
);

AOI22xp5_ASAP7_75t_L g206 ( 
.A1(n_185),
.A2(n_161),
.B1(n_167),
.B2(n_156),
.Y(n_206)
);

MAJIxp5_ASAP7_75t_L g186 ( 
.A(n_162),
.B(n_159),
.C(n_164),
.Y(n_186)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_188),
.Y(n_207)
);

AOI22xp5_ASAP7_75t_L g191 ( 
.A1(n_170),
.A2(n_105),
.B1(n_145),
.B2(n_126),
.Y(n_191)
);

OAI22xp5_ASAP7_75t_L g197 ( 
.A1(n_191),
.A2(n_171),
.B1(n_175),
.B2(n_173),
.Y(n_197)
);

INVxp67_ASAP7_75t_L g193 ( 
.A(n_154),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_SL g204 ( 
.A(n_193),
.B(n_168),
.Y(n_204)
);

MAJIxp5_ASAP7_75t_L g195 ( 
.A(n_165),
.B(n_110),
.C(n_145),
.Y(n_195)
);

NOR2xp33_ASAP7_75t_L g199 ( 
.A(n_195),
.B(n_196),
.Y(n_199)
);

AOI322xp5_ASAP7_75t_L g196 ( 
.A1(n_174),
.A2(n_110),
.A3(n_149),
.B1(n_111),
.B2(n_117),
.C1(n_13),
.C2(n_14),
.Y(n_196)
);

NAND2xp5_ASAP7_75t_L g216 ( 
.A(n_197),
.B(n_201),
.Y(n_216)
);

NAND2xp5_ASAP7_75t_L g198 ( 
.A(n_189),
.B(n_176),
.Y(n_198)
);

CKINVDCx20_ASAP7_75t_R g214 ( 
.A(n_198),
.Y(n_214)
);

OAI22xp5_ASAP7_75t_L g200 ( 
.A1(n_193),
.A2(n_169),
.B1(n_160),
.B2(n_163),
.Y(n_200)
);

OAI22xp5_ASAP7_75t_L g223 ( 
.A1(n_200),
.A2(n_204),
.B1(n_179),
.B2(n_161),
.Y(n_223)
);

INVxp67_ASAP7_75t_L g201 ( 
.A(n_194),
.Y(n_201)
);

XNOR2xp5_ASAP7_75t_SL g202 ( 
.A(n_182),
.B(n_155),
.Y(n_202)
);

XNOR2xp5_ASAP7_75t_L g219 ( 
.A(n_202),
.B(n_208),
.Y(n_219)
);

OAI21xp5_ASAP7_75t_L g203 ( 
.A1(n_178),
.A2(n_163),
.B(n_169),
.Y(n_203)
);

OAI21xp5_ASAP7_75t_L g221 ( 
.A1(n_203),
.A2(n_194),
.B(n_180),
.Y(n_221)
);

AO21x1_ASAP7_75t_L g218 ( 
.A1(n_205),
.A2(n_183),
.B(n_187),
.Y(n_218)
);

OAI22xp5_ASAP7_75t_SL g217 ( 
.A1(n_206),
.A2(n_187),
.B1(n_189),
.B2(n_191),
.Y(n_217)
);

XNOR2xp5_ASAP7_75t_SL g208 ( 
.A(n_178),
.B(n_157),
.Y(n_208)
);

NOR2xp33_ASAP7_75t_SL g210 ( 
.A(n_192),
.B(n_156),
.Y(n_210)
);

NOR2xp33_ASAP7_75t_L g212 ( 
.A(n_210),
.B(n_192),
.Y(n_212)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_212),
.Y(n_230)
);

MAJIxp5_ASAP7_75t_L g213 ( 
.A(n_209),
.B(n_186),
.C(n_181),
.Y(n_213)
);

MAJIxp5_ASAP7_75t_L g227 ( 
.A(n_213),
.B(n_220),
.C(n_205),
.Y(n_227)
);

INVx5_ASAP7_75t_L g215 ( 
.A(n_211),
.Y(n_215)
);

NOR2xp33_ASAP7_75t_SL g226 ( 
.A(n_215),
.B(n_222),
.Y(n_226)
);

AOI22xp5_ASAP7_75t_L g224 ( 
.A1(n_217),
.A2(n_208),
.B1(n_201),
.B2(n_185),
.Y(n_224)
);

AOI21xp5_ASAP7_75t_L g228 ( 
.A1(n_218),
.A2(n_221),
.B(n_223),
.Y(n_228)
);

MAJIxp5_ASAP7_75t_L g220 ( 
.A(n_209),
.B(n_179),
.C(n_184),
.Y(n_220)
);

NOR2xp33_ASAP7_75t_L g222 ( 
.A(n_207),
.B(n_190),
.Y(n_222)
);

NAND2xp5_ASAP7_75t_SL g233 ( 
.A(n_224),
.B(n_218),
.Y(n_233)
);

XNOR2xp5_ASAP7_75t_L g225 ( 
.A(n_213),
.B(n_202),
.Y(n_225)
);

MAJIxp5_ASAP7_75t_L g234 ( 
.A(n_225),
.B(n_227),
.C(n_229),
.Y(n_234)
);

XNOR2xp5_ASAP7_75t_L g229 ( 
.A(n_220),
.B(n_203),
.Y(n_229)
);

AOI21xp5_ASAP7_75t_L g231 ( 
.A1(n_221),
.A2(n_198),
.B(n_199),
.Y(n_231)
);

OAI21xp5_ASAP7_75t_SL g236 ( 
.A1(n_231),
.A2(n_216),
.B(n_217),
.Y(n_236)
);

XNOR2xp5_ASAP7_75t_L g232 ( 
.A(n_219),
.B(n_206),
.Y(n_232)
);

NAND2xp5_ASAP7_75t_L g235 ( 
.A(n_232),
.B(n_216),
.Y(n_235)
);

A2O1A1Ixp33_ASAP7_75t_SL g241 ( 
.A1(n_233),
.A2(n_232),
.B(n_229),
.C(n_227),
.Y(n_241)
);

XNOR2xp5_ASAP7_75t_L g240 ( 
.A(n_235),
.B(n_237),
.Y(n_240)
);

MAJIxp5_ASAP7_75t_L g243 ( 
.A(n_236),
.B(n_184),
.C(n_10),
.Y(n_243)
);

NAND2xp5_ASAP7_75t_L g237 ( 
.A(n_226),
.B(n_215),
.Y(n_237)
);

NAND2xp5_ASAP7_75t_L g238 ( 
.A(n_230),
.B(n_214),
.Y(n_238)
);

OAI21xp5_ASAP7_75t_SL g244 ( 
.A1(n_238),
.A2(n_9),
.B(n_11),
.Y(n_244)
);

AOI31xp33_ASAP7_75t_L g239 ( 
.A1(n_228),
.A2(n_158),
.A3(n_195),
.B(n_219),
.Y(n_239)
);

AOI21x1_ASAP7_75t_L g242 ( 
.A1(n_239),
.A2(n_225),
.B(n_190),
.Y(n_242)
);

OR2x2_ASAP7_75t_L g247 ( 
.A(n_241),
.B(n_243),
.Y(n_247)
);

AOI21x1_ASAP7_75t_L g245 ( 
.A1(n_242),
.A2(n_244),
.B(n_11),
.Y(n_245)
);

OAI22xp5_ASAP7_75t_SL g249 ( 
.A1(n_245),
.A2(n_246),
.B1(n_12),
.B2(n_13),
.Y(n_249)
);

O2A1O1Ixp33_ASAP7_75t_SL g246 ( 
.A1(n_240),
.A2(n_234),
.B(n_13),
.C(n_15),
.Y(n_246)
);

NOR2xp33_ASAP7_75t_L g248 ( 
.A(n_247),
.B(n_234),
.Y(n_248)
);

AOI21xp5_ASAP7_75t_L g250 ( 
.A1(n_248),
.A2(n_249),
.B(n_241),
.Y(n_250)
);

OAI22xp5_ASAP7_75t_SL g251 ( 
.A1(n_250),
.A2(n_249),
.B1(n_15),
.B2(n_16),
.Y(n_251)
);

XNOR2xp5_ASAP7_75t_SL g252 ( 
.A(n_251),
.B(n_12),
.Y(n_252)
);


endmodule