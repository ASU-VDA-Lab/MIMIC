module fake_jpeg_26083_n_152 (n_13, n_21, n_33, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_40, n_19, n_18, n_20, n_35, n_41, n_4, n_34, n_30, n_39, n_42, n_16, n_3, n_0, n_24, n_28, n_38, n_26, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_43, n_12, n_32, n_8, n_15, n_7, n_152);

input n_13;
input n_21;
input n_33;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_42;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_43;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_152;

wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_147;
wire n_73;
wire n_84;
wire n_59;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_49;
wire n_76;
wire n_127;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_103;
wire n_50;
wire n_150;
wire n_124;
wire n_141;
wire n_57;
wire n_119;
wire n_69;
wire n_83;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_106;
wire n_111;
wire n_44;
wire n_143;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_78;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_91;
wire n_54;
wire n_93;
wire n_138;
wire n_101;
wire n_48;
wire n_149;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_135;
wire n_62;
wire n_120;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_17),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_29),
.Y(n_45)
);

INVx2_ASAP7_75t_L g46 ( 
.A(n_23),
.Y(n_46)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_28),
.Y(n_47)
);

INVx1_ASAP7_75t_SL g48 ( 
.A(n_35),
.Y(n_48)
);

BUFx12f_ASAP7_75t_L g49 ( 
.A(n_20),
.Y(n_49)
);

CKINVDCx14_ASAP7_75t_R g50 ( 
.A(n_3),
.Y(n_50)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_9),
.Y(n_51)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_16),
.Y(n_52)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_13),
.Y(n_53)
);

INVx4_ASAP7_75t_L g54 ( 
.A(n_40),
.Y(n_54)
);

CKINVDCx20_ASAP7_75t_R g55 ( 
.A(n_42),
.Y(n_55)
);

INVx13_ASAP7_75t_L g56 ( 
.A(n_9),
.Y(n_56)
);

BUFx2_ASAP7_75t_L g57 ( 
.A(n_1),
.Y(n_57)
);

CKINVDCx20_ASAP7_75t_R g58 ( 
.A(n_5),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_26),
.Y(n_59)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_38),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_6),
.Y(n_61)
);

INVx4_ASAP7_75t_L g62 ( 
.A(n_6),
.Y(n_62)
);

BUFx3_ASAP7_75t_L g63 ( 
.A(n_34),
.Y(n_63)
);

BUFx5_ASAP7_75t_L g64 ( 
.A(n_39),
.Y(n_64)
);

BUFx10_ASAP7_75t_L g65 ( 
.A(n_31),
.Y(n_65)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_7),
.Y(n_66)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_15),
.Y(n_67)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_3),
.Y(n_68)
);

AOI22xp5_ASAP7_75t_L g69 ( 
.A1(n_46),
.A2(n_22),
.B1(n_43),
.B2(n_41),
.Y(n_69)
);

AOI22xp5_ASAP7_75t_L g86 ( 
.A1(n_69),
.A2(n_50),
.B1(n_56),
.B2(n_48),
.Y(n_86)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_57),
.Y(n_70)
);

INVx2_ASAP7_75t_L g76 ( 
.A(n_70),
.Y(n_76)
);

INVx8_ASAP7_75t_L g71 ( 
.A(n_65),
.Y(n_71)
);

INVx5_ASAP7_75t_L g80 ( 
.A(n_71),
.Y(n_80)
);

INVx4_ASAP7_75t_SL g72 ( 
.A(n_49),
.Y(n_72)
);

BUFx16f_ASAP7_75t_L g84 ( 
.A(n_72),
.Y(n_84)
);

CKINVDCx20_ASAP7_75t_R g73 ( 
.A(n_44),
.Y(n_73)
);

OR2x2_ASAP7_75t_L g87 ( 
.A(n_73),
.B(n_75),
.Y(n_87)
);

INVx11_ASAP7_75t_L g74 ( 
.A(n_49),
.Y(n_74)
);

INVx2_ASAP7_75t_L g88 ( 
.A(n_74),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_L g75 ( 
.A(n_65),
.B(n_0),
.Y(n_75)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_71),
.Y(n_77)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_77),
.Y(n_93)
);

BUFx6f_ASAP7_75t_L g78 ( 
.A(n_74),
.Y(n_78)
);

INVx2_ASAP7_75t_L g90 ( 
.A(n_78),
.Y(n_90)
);

AOI22xp33_ASAP7_75t_L g79 ( 
.A1(n_70),
.A2(n_60),
.B1(n_54),
.B2(n_62),
.Y(n_79)
);

OAI22xp5_ASAP7_75t_L g91 ( 
.A1(n_79),
.A2(n_65),
.B1(n_57),
.B2(n_61),
.Y(n_91)
);

BUFx6f_ASAP7_75t_L g81 ( 
.A(n_72),
.Y(n_81)
);

INVx2_ASAP7_75t_L g92 ( 
.A(n_81),
.Y(n_92)
);

INVx3_ASAP7_75t_L g82 ( 
.A(n_75),
.Y(n_82)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_82),
.Y(n_95)
);

BUFx6f_ASAP7_75t_L g83 ( 
.A(n_69),
.Y(n_83)
);

INVx2_ASAP7_75t_L g96 ( 
.A(n_83),
.Y(n_96)
);

BUFx6f_ASAP7_75t_L g85 ( 
.A(n_71),
.Y(n_85)
);

INVx2_ASAP7_75t_L g101 ( 
.A(n_85),
.Y(n_101)
);

OAI22xp5_ASAP7_75t_SL g94 ( 
.A1(n_86),
.A2(n_68),
.B1(n_58),
.B2(n_51),
.Y(n_94)
);

AOI22xp5_ASAP7_75t_SL g89 ( 
.A1(n_79),
.A2(n_50),
.B1(n_56),
.B2(n_66),
.Y(n_89)
);

AND2x2_ASAP7_75t_L g106 ( 
.A(n_89),
.B(n_91),
.Y(n_106)
);

OAI22xp5_ASAP7_75t_SL g108 ( 
.A1(n_94),
.A2(n_98),
.B1(n_53),
.B2(n_88),
.Y(n_108)
);

INVx5_ASAP7_75t_L g97 ( 
.A(n_84),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_97),
.B(n_100),
.Y(n_103)
);

AOI22xp33_ASAP7_75t_SL g98 ( 
.A1(n_80),
.A2(n_49),
.B1(n_45),
.B2(n_47),
.Y(n_98)
);

MAJIxp5_ASAP7_75t_L g99 ( 
.A(n_76),
.B(n_59),
.C(n_67),
.Y(n_99)
);

MAJIxp5_ASAP7_75t_L g104 ( 
.A(n_99),
.B(n_61),
.C(n_59),
.Y(n_104)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_87),
.Y(n_100)
);

INVx2_ASAP7_75t_L g102 ( 
.A(n_90),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_L g123 ( 
.A(n_102),
.B(n_109),
.Y(n_123)
);

AND2x2_ASAP7_75t_L g116 ( 
.A(n_104),
.B(n_108),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_95),
.B(n_55),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_L g114 ( 
.A(n_105),
.B(n_107),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g107 ( 
.A(n_96),
.B(n_52),
.Y(n_107)
);

INVx1_ASAP7_75t_SL g109 ( 
.A(n_97),
.Y(n_109)
);

AOI22xp33_ASAP7_75t_L g110 ( 
.A1(n_101),
.A2(n_85),
.B1(n_63),
.B2(n_78),
.Y(n_110)
);

OAI22xp5_ASAP7_75t_L g119 ( 
.A1(n_110),
.A2(n_2),
.B1(n_4),
.B2(n_5),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_93),
.B(n_0),
.Y(n_111)
);

CKINVDCx14_ASAP7_75t_R g117 ( 
.A(n_111),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_L g112 ( 
.A(n_99),
.B(n_98),
.Y(n_112)
);

MAJIxp5_ASAP7_75t_L g121 ( 
.A(n_112),
.B(n_25),
.C(n_37),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_SL g113 ( 
.A(n_92),
.B(n_84),
.Y(n_113)
);

OAI21xp5_ASAP7_75t_SL g118 ( 
.A1(n_113),
.A2(n_1),
.B(n_2),
.Y(n_118)
);

HAxp5_ASAP7_75t_SL g115 ( 
.A(n_106),
.B(n_64),
.CON(n_115),
.SN(n_115)
);

OAI21xp5_ASAP7_75t_L g129 ( 
.A1(n_115),
.A2(n_118),
.B(n_120),
.Y(n_129)
);

OAI22xp5_ASAP7_75t_L g132 ( 
.A1(n_119),
.A2(n_122),
.B1(n_10),
.B2(n_12),
.Y(n_132)
);

OAI21xp5_ASAP7_75t_L g120 ( 
.A1(n_106),
.A2(n_4),
.B(n_7),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_SL g124 ( 
.A(n_121),
.B(n_30),
.Y(n_124)
);

AOI22xp33_ASAP7_75t_SL g122 ( 
.A1(n_110),
.A2(n_24),
.B1(n_36),
.B2(n_11),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_L g140 ( 
.A(n_124),
.B(n_125),
.Y(n_140)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_123),
.Y(n_125)
);

AOI22xp5_ASAP7_75t_SL g126 ( 
.A1(n_116),
.A2(n_109),
.B1(n_103),
.B2(n_8),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_L g136 ( 
.A(n_126),
.B(n_127),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_SL g127 ( 
.A(n_114),
.B(n_8),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_SL g128 ( 
.A(n_117),
.B(n_10),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_L g139 ( 
.A(n_128),
.B(n_131),
.Y(n_139)
);

CKINVDCx20_ASAP7_75t_R g130 ( 
.A(n_116),
.Y(n_130)
);

CKINVDCx20_ASAP7_75t_R g137 ( 
.A(n_130),
.Y(n_137)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_115),
.Y(n_131)
);

CKINVDCx20_ASAP7_75t_R g141 ( 
.A(n_132),
.Y(n_141)
);

CKINVDCx20_ASAP7_75t_R g133 ( 
.A(n_122),
.Y(n_133)
);

XOR2xp5_ASAP7_75t_L g138 ( 
.A(n_133),
.B(n_134),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_SL g134 ( 
.A(n_114),
.B(n_14),
.Y(n_134)
);

OAI21xp5_ASAP7_75t_L g135 ( 
.A1(n_116),
.A2(n_18),
.B(n_19),
.Y(n_135)
);

XOR2xp5_ASAP7_75t_L g142 ( 
.A(n_138),
.B(n_135),
.Y(n_142)
);

AOI22xp5_ASAP7_75t_L g144 ( 
.A1(n_142),
.A2(n_143),
.B1(n_136),
.B2(n_139),
.Y(n_144)
);

CKINVDCx20_ASAP7_75t_R g143 ( 
.A(n_137),
.Y(n_143)
);

NAND4xp25_ASAP7_75t_L g145 ( 
.A(n_144),
.B(n_138),
.C(n_141),
.D(n_126),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_L g146 ( 
.A(n_145),
.B(n_135),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_SL g147 ( 
.A(n_146),
.B(n_140),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_L g148 ( 
.A(n_147),
.B(n_129),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_L g149 ( 
.A(n_148),
.B(n_21),
.Y(n_149)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_149),
.Y(n_150)
);

OAI21xp5_ASAP7_75t_L g151 ( 
.A1(n_150),
.A2(n_27),
.B(n_32),
.Y(n_151)
);

XOR2xp5_ASAP7_75t_L g152 ( 
.A(n_151),
.B(n_33),
.Y(n_152)
);


endmodule