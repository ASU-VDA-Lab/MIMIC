module real_jpeg_32801_n_18 (n_17, n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_16, n_3, n_10, n_9, n_18);

input n_17;
input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_16;
input n_3;
input n_10;
input n_9;

output n_18;

wire n_384;
wire n_37;
wire n_430;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_460;
wire n_300;
wire n_415;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_271;
wire n_47;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_446;
wire n_199;
wire n_95;
wire n_441;
wire n_238;
wire n_67;
wire n_350;
wire n_235;
wire n_107;
wire n_369;
wire n_376;
wire n_354;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_355;
wire n_123;
wire n_463;
wire n_425;
wire n_455;
wire n_462;
wire n_50;
wire n_409;
wire n_186;
wire n_137;
wire n_72;
wire n_440;
wire n_171;
wire n_151;
wire n_272;
wire n_461;
wire n_198;
wire n_203;
wire n_23;
wire n_362;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_339;
wire n_326;
wire n_80;
wire n_30;
wire n_328;
wire n_149;
wire n_332;
wire n_366;
wire n_456;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_353;
wire n_453;
wire n_230;
wire n_417;
wire n_428;
wire n_128;
wire n_216;
wire n_202;
wire n_367;
wire n_127;
wire n_356;
wire n_365;
wire n_464;
wire n_423;
wire n_36;
wire n_102;
wire n_81;
wire n_101;
wire n_422;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_348;
wire n_252;
wire n_363;
wire n_310;
wire n_345;
wire n_83;
wire n_78;
wire n_288;
wire n_221;
wire n_393;
wire n_104;
wire n_153;
wire n_443;
wire n_337;
wire n_131;
wire n_439;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_378;
wire n_200;
wire n_432;
wire n_465;
wire n_335;
wire n_214;
wire n_113;
wire n_251;
wire n_459;
wire n_139;
wire n_33;
wire n_175;
wire n_338;
wire n_156;
wire n_387;
wire n_434;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_390;
wire n_77;
wire n_399;
wire n_219;
wire n_372;
wire n_122;
wire n_19;
wire n_262;
wire n_334;
wire n_383;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_426;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_371;
wire n_410;
wire n_421;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_411;
wire n_382;
wire n_20;
wire n_278;
wire n_314;
wire n_103;
wire n_232;
wire n_448;
wire n_212;
wire n_284;
wire n_402;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_452;
wire n_213;
wire n_25;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_407;
wire n_419;
wire n_386;
wire n_341;
wire n_331;
wire n_49;
wire n_68;
wire n_395;
wire n_146;
wire n_286;
wire n_215;
wire n_176;
wire n_166;
wire n_323;
wire n_312;
wire n_325;
wire n_307;
wire n_316;
wire n_161;
wire n_207;
wire n_431;
wire n_420;
wire n_357;
wire n_237;
wire n_445;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_380;
wire n_414;
wire n_140;
wire n_126;
wire n_342;
wire n_120;
wire n_155;
wire n_412;
wire n_405;
wire n_319;
wire n_93;
wire n_242;
wire n_142;
wire n_397;
wire n_76;
wire n_403;
wire n_79;
wire n_282;
wire n_147;
wire n_359;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_449;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_145;
wire n_266;
wire n_377;
wire n_109;
wire n_391;
wire n_427;
wire n_401;
wire n_148;
wire n_373;
wire n_396;
wire n_392;
wire n_196;
wire n_375;
wire n_298;
wire n_330;
wire n_450;
wire n_333;
wire n_152;
wire n_270;
wire n_159;
wire n_429;
wire n_347;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_336;
wire n_258;
wire n_458;
wire n_150;
wire n_41;
wire n_74;
wire n_404;
wire n_158;
wire n_204;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_413;
wire n_75;
wire n_346;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_457;
wire n_119;
wire n_283;
wire n_358;
wire n_181;
wire n_256;
wire n_273;
wire n_253;
wire n_54;
wire n_168;
wire n_38;
wire n_442;
wire n_385;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_349;
wire n_418;
wire n_343;
wire n_292;
wire n_64;
wire n_291;
wire n_236;
wire n_370;
wire n_276;
wire n_374;
wire n_287;
wire n_388;
wire n_174;
wire n_400;
wire n_255;
wire n_243;
wire n_299;
wire n_352;
wire n_56;
wire n_293;
wire n_275;
wire n_381;
wire n_227;
wire n_229;
wire n_454;
wire n_379;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_444;
wire n_360;
wire n_398;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_451;
wire n_45;
wire n_437;
wire n_268;
wire n_42;
wire n_313;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_416;
wire n_143;
wire n_351;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_406;
wire n_303;
wire n_321;
wire n_100;
wire n_368;
wire n_51;
wire n_205;
wire n_361;
wire n_324;
wire n_86;
wire n_261;
wire n_70;
wire n_435;
wire n_32;
wire n_228;
wire n_389;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_438;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_394;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_436;
wire n_169;
wire n_88;
wire n_167;
wire n_295;
wire n_424;
wire n_133;
wire n_447;
wire n_257;
wire n_344;
wire n_210;
wire n_206;
wire n_408;
wire n_85;
wire n_96;
wire n_308;
wire n_433;
wire n_364;

NAND2x1p5_ASAP7_75t_L g32 ( 
.A(n_0),
.B(n_33),
.Y(n_32)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_0),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_SL g249 ( 
.A(n_0),
.B(n_250),
.Y(n_249)
);

NAND2x1_ASAP7_75t_L g264 ( 
.A(n_0),
.B(n_265),
.Y(n_264)
);

NAND2xp33_ASAP7_75t_R g270 ( 
.A(n_0),
.B(n_271),
.Y(n_270)
);

NAND2xp5_ASAP7_75t_L g314 ( 
.A(n_0),
.B(n_315),
.Y(n_314)
);

AND2x4_ASAP7_75t_L g334 ( 
.A(n_0),
.B(n_102),
.Y(n_334)
);

NAND2xp5_ASAP7_75t_L g342 ( 
.A(n_0),
.B(n_343),
.Y(n_342)
);

NAND2xp5_ASAP7_75t_L g365 ( 
.A(n_0),
.B(n_262),
.Y(n_365)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_1),
.Y(n_37)
);

INVx2_ASAP7_75t_L g89 ( 
.A(n_1),
.Y(n_89)
);

BUFx3_ASAP7_75t_L g263 ( 
.A(n_1),
.Y(n_263)
);

BUFx12f_ASAP7_75t_L g306 ( 
.A(n_1),
.Y(n_306)
);

AND2x4_ASAP7_75t_L g35 ( 
.A(n_2),
.B(n_36),
.Y(n_35)
);

AND2x2_ASAP7_75t_L g66 ( 
.A(n_2),
.B(n_67),
.Y(n_66)
);

AND2x2_ASAP7_75t_L g114 ( 
.A(n_2),
.B(n_115),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_SL g126 ( 
.A(n_2),
.B(n_127),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_L g152 ( 
.A(n_2),
.B(n_153),
.Y(n_152)
);

NAND2x1p5_ASAP7_75t_L g223 ( 
.A(n_2),
.B(n_130),
.Y(n_223)
);

NAND2xp5_ASAP7_75t_SL g439 ( 
.A(n_2),
.B(n_440),
.Y(n_439)
);

AND2x2_ASAP7_75t_SL g57 ( 
.A(n_3),
.B(n_58),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_L g71 ( 
.A(n_3),
.B(n_72),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_L g94 ( 
.A(n_3),
.B(n_95),
.Y(n_94)
);

NAND2x1_ASAP7_75t_L g142 ( 
.A(n_3),
.B(n_143),
.Y(n_142)
);

AND2x2_ASAP7_75t_L g245 ( 
.A(n_3),
.B(n_246),
.Y(n_245)
);

INVxp67_ASAP7_75t_L g308 ( 
.A(n_3),
.Y(n_308)
);

NAND2xp5_ASAP7_75t_L g319 ( 
.A(n_3),
.B(n_320),
.Y(n_319)
);

NAND2xp5_ASAP7_75t_L g347 ( 
.A(n_3),
.B(n_348),
.Y(n_347)
);

CKINVDCx5p33_ASAP7_75t_R g20 ( 
.A(n_4),
.Y(n_20)
);

NAND2xp5_ASAP7_75t_L g61 ( 
.A(n_5),
.B(n_62),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_L g156 ( 
.A(n_5),
.B(n_157),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_SL g241 ( 
.A(n_5),
.B(n_242),
.Y(n_241)
);

NAND2xp5_ASAP7_75t_L g323 ( 
.A(n_5),
.B(n_324),
.Y(n_323)
);

NAND2xp5_ASAP7_75t_L g336 ( 
.A(n_5),
.B(n_337),
.Y(n_336)
);

NAND2xp5_ASAP7_75t_L g357 ( 
.A(n_5),
.B(n_358),
.Y(n_357)
);

NAND2xp5_ASAP7_75t_L g361 ( 
.A(n_5),
.B(n_362),
.Y(n_361)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_6),
.Y(n_34)
);

BUFx3_ASAP7_75t_L g160 ( 
.A(n_6),
.Y(n_160)
);

BUFx3_ASAP7_75t_L g212 ( 
.A(n_6),
.Y(n_212)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_7),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g189 ( 
.A(n_7),
.Y(n_189)
);

INVx4_ASAP7_75t_L g51 ( 
.A(n_8),
.Y(n_51)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_8),
.Y(n_68)
);

BUFx6f_ASAP7_75t_L g291 ( 
.A(n_8),
.Y(n_291)
);

BUFx6f_ASAP7_75t_L g310 ( 
.A(n_8),
.Y(n_310)
);

AND2x2_ASAP7_75t_L g48 ( 
.A(n_9),
.B(n_49),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_L g100 ( 
.A(n_9),
.B(n_101),
.Y(n_100)
);

NAND2x1_ASAP7_75t_L g172 ( 
.A(n_9),
.B(n_173),
.Y(n_172)
);

AND2x2_ASAP7_75t_L g185 ( 
.A(n_9),
.B(n_186),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_L g192 ( 
.A(n_9),
.B(n_186),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_SL g261 ( 
.A(n_9),
.B(n_262),
.Y(n_261)
);

NAND2xp5_ASAP7_75t_SL g450 ( 
.A(n_9),
.B(n_451),
.Y(n_450)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_10),
.Y(n_22)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_11),
.Y(n_56)
);

BUFx3_ASAP7_75t_L g77 ( 
.A(n_11),
.Y(n_77)
);

BUFx6f_ASAP7_75t_L g128 ( 
.A(n_11),
.Y(n_128)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_12),
.Y(n_64)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_12),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g40 ( 
.A(n_13),
.B(n_41),
.Y(n_40)
);

AND2x2_ASAP7_75t_L g53 ( 
.A(n_13),
.B(n_54),
.Y(n_53)
);

AND2x2_ASAP7_75t_SL g79 ( 
.A(n_13),
.B(n_80),
.Y(n_79)
);

AND2x2_ASAP7_75t_L g110 ( 
.A(n_13),
.B(n_111),
.Y(n_110)
);

AND2x4_ASAP7_75t_L g133 ( 
.A(n_13),
.B(n_134),
.Y(n_133)
);

AND2x4_ASAP7_75t_L g190 ( 
.A(n_13),
.B(n_191),
.Y(n_190)
);

AND2x2_ASAP7_75t_L g219 ( 
.A(n_13),
.B(n_67),
.Y(n_219)
);

AND2x2_ASAP7_75t_SL g428 ( 
.A(n_13),
.B(n_429),
.Y(n_428)
);

INVx2_ASAP7_75t_L g82 ( 
.A(n_14),
.Y(n_82)
);

INVx4_ASAP7_75t_L g155 ( 
.A(n_14),
.Y(n_155)
);

INVxp67_ASAP7_75t_L g86 ( 
.A(n_15),
.Y(n_86)
);

AND2x2_ASAP7_75t_L g139 ( 
.A(n_15),
.B(n_140),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_L g221 ( 
.A(n_15),
.B(n_222),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_SL g269 ( 
.A(n_15),
.B(n_262),
.Y(n_269)
);

NAND2xp5_ASAP7_75t_L g435 ( 
.A(n_15),
.B(n_436),
.Y(n_435)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_16),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g137 ( 
.A(n_16),
.Y(n_137)
);

INVx2_ASAP7_75t_L g244 ( 
.A(n_16),
.Y(n_244)
);

BUFx6f_ASAP7_75t_L g453 ( 
.A(n_16),
.Y(n_453)
);

NAND2xp5_ASAP7_75t_SL g75 ( 
.A(n_17),
.B(n_76),
.Y(n_75)
);

NAND2x1_ASAP7_75t_L g129 ( 
.A(n_17),
.B(n_130),
.Y(n_129)
);

AND2x2_ASAP7_75t_L g149 ( 
.A(n_17),
.B(n_150),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_L g175 ( 
.A(n_17),
.B(n_176),
.Y(n_175)
);

AND2x4_ASAP7_75t_SL g210 ( 
.A(n_17),
.B(n_211),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_SL g284 ( 
.A(n_17),
.B(n_285),
.Y(n_284)
);

NAND2xp5_ASAP7_75t_SL g288 ( 
.A(n_17),
.B(n_289),
.Y(n_288)
);

INVxp67_ASAP7_75t_L g304 ( 
.A(n_17),
.Y(n_304)
);

OAI211xp5_ASAP7_75t_L g18 ( 
.A1(n_19),
.A2(n_21),
.B(n_23),
.C(n_463),
.Y(n_18)
);

NOR2xp33_ASAP7_75t_L g21 ( 
.A(n_19),
.B(n_22),
.Y(n_21)
);

CKINVDCx5p33_ASAP7_75t_R g19 ( 
.A(n_20),
.Y(n_19)
);

NOR2xp33_ASAP7_75t_L g414 ( 
.A(n_21),
.B(n_415),
.Y(n_414)
);

INVx1_ASAP7_75t_L g464 ( 
.A(n_21),
.Y(n_464)
);

OAI21xp33_ASAP7_75t_L g23 ( 
.A1(n_24),
.A2(n_411),
.B(n_414),
.Y(n_23)
);

NOR2xp33_ASAP7_75t_L g24 ( 
.A(n_25),
.B(n_226),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_26),
.Y(n_25)
);

A2O1A1Ixp33_ASAP7_75t_R g465 ( 
.A1(n_26),
.A2(n_227),
.B(n_388),
.C(n_407),
.Y(n_465)
);

NAND2xp5_ASAP7_75t_L g26 ( 
.A(n_27),
.B(n_178),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_28),
.Y(n_27)
);

NAND2xp5_ASAP7_75t_L g413 ( 
.A(n_28),
.B(n_179),
.Y(n_413)
);

MAJIxp5_ASAP7_75t_L g28 ( 
.A(n_29),
.B(n_105),
.C(n_145),
.Y(n_28)
);

XNOR2xp5_ASAP7_75t_L g405 ( 
.A(n_29),
.B(n_406),
.Y(n_405)
);

MAJIxp5_ASAP7_75t_L g29 ( 
.A(n_30),
.B(n_46),
.C(n_83),
.Y(n_29)
);

XOR2xp5_ASAP7_75t_L g402 ( 
.A(n_30),
.B(n_84),
.Y(n_402)
);

OAI22xp5_ASAP7_75t_SL g30 ( 
.A1(n_31),
.A2(n_38),
.B1(n_44),
.B2(n_45),
.Y(n_30)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_31),
.Y(n_44)
);

XNOR2xp5_ASAP7_75t_SL g31 ( 
.A(n_32),
.B(n_35),
.Y(n_31)
);

MAJIxp5_ASAP7_75t_L g168 ( 
.A(n_32),
.B(n_35),
.C(n_169),
.Y(n_168)
);

INVx2_ASAP7_75t_SL g430 ( 
.A(n_33),
.Y(n_430)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_34),
.Y(n_33)
);

INVx6_ASAP7_75t_L g144 ( 
.A(n_34),
.Y(n_144)
);

AND2x2_ASAP7_75t_L g260 ( 
.A(n_35),
.B(n_219),
.Y(n_260)
);

OAI21x1_ASAP7_75t_L g292 ( 
.A1(n_35),
.A2(n_218),
.B(n_293),
.Y(n_292)
);

NAND2xp5_ASAP7_75t_L g293 ( 
.A(n_35),
.B(n_294),
.Y(n_293)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_37),
.Y(n_36)
);

HB1xp67_ASAP7_75t_L g38 ( 
.A(n_39),
.Y(n_38)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_39),
.Y(n_45)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_40),
.Y(n_39)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_40),
.Y(n_169)
);

INVxp67_ASAP7_75t_L g41 ( 
.A(n_42),
.Y(n_41)
);

INVx5_ASAP7_75t_L g150 ( 
.A(n_42),
.Y(n_150)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_43),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g74 ( 
.A(n_43),
.Y(n_74)
);

XOR2x2_ASAP7_75t_SL g401 ( 
.A(n_46),
.B(n_402),
.Y(n_401)
);

MAJIxp5_ASAP7_75t_L g46 ( 
.A(n_47),
.B(n_60),
.C(n_69),
.Y(n_46)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_47),
.Y(n_255)
);

XNOR2xp5_ASAP7_75t_SL g47 ( 
.A(n_48),
.B(n_52),
.Y(n_47)
);

MAJIxp5_ASAP7_75t_L g161 ( 
.A(n_48),
.B(n_53),
.C(n_57),
.Y(n_161)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_50),
.Y(n_49)
);

INVx2_ASAP7_75t_L g50 ( 
.A(n_51),
.Y(n_50)
);

INVx2_ASAP7_75t_L g123 ( 
.A(n_51),
.Y(n_123)
);

XOR2xp5_ASAP7_75t_L g52 ( 
.A(n_53),
.B(n_57),
.Y(n_52)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_55),
.Y(n_54)
);

INVx2_ASAP7_75t_L g338 ( 
.A(n_55),
.Y(n_338)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_56),
.Y(n_55)
);

BUFx5_ASAP7_75t_L g247 ( 
.A(n_56),
.Y(n_247)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_59),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g130 ( 
.A(n_59),
.Y(n_130)
);

XNOR2xp5_ASAP7_75t_L g254 ( 
.A(n_60),
.B(n_70),
.Y(n_254)
);

OR2x2_ASAP7_75t_L g60 ( 
.A(n_61),
.B(n_65),
.Y(n_60)
);

OAI22xp5_ASAP7_75t_SL g237 ( 
.A1(n_61),
.A2(n_65),
.B1(n_66),
.B2(n_238),
.Y(n_237)
);

INVxp67_ASAP7_75t_L g238 ( 
.A(n_61),
.Y(n_238)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_63),
.Y(n_62)
);

INVx2_ASAP7_75t_L g176 ( 
.A(n_63),
.Y(n_176)
);

INVx2_ASAP7_75t_L g63 ( 
.A(n_64),
.Y(n_63)
);

BUFx6f_ASAP7_75t_L g92 ( 
.A(n_64),
.Y(n_92)
);

BUFx6f_ASAP7_75t_L g191 ( 
.A(n_64),
.Y(n_191)
);

BUFx3_ASAP7_75t_L g440 ( 
.A(n_64),
.Y(n_440)
);

AOI22xp5_ASAP7_75t_L g109 ( 
.A1(n_65),
.A2(n_66),
.B1(n_110),
.B2(n_112),
.Y(n_109)
);

INVx1_ASAP7_75t_SL g65 ( 
.A(n_66),
.Y(n_65)
);

MAJIxp5_ASAP7_75t_L g183 ( 
.A(n_66),
.B(n_110),
.C(n_114),
.Y(n_183)
);

INVx2_ASAP7_75t_L g67 ( 
.A(n_68),
.Y(n_67)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_70),
.Y(n_69)
);

MAJIxp5_ASAP7_75t_L g70 ( 
.A(n_71),
.B(n_75),
.C(n_78),
.Y(n_70)
);

AOI22xp5_ASAP7_75t_L g234 ( 
.A1(n_71),
.A2(n_78),
.B1(n_79),
.B2(n_235),
.Y(n_234)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_71),
.Y(n_235)
);

HB1xp67_ASAP7_75t_L g72 ( 
.A(n_73),
.Y(n_72)
);

INVx2_ASAP7_75t_L g73 ( 
.A(n_74),
.Y(n_73)
);

INVx2_ASAP7_75t_L g115 ( 
.A(n_74),
.Y(n_115)
);

INVx4_ASAP7_75t_L g326 ( 
.A(n_74),
.Y(n_326)
);

INVx1_ASAP7_75t_L g436 ( 
.A(n_74),
.Y(n_436)
);

XNOR2xp5_ASAP7_75t_L g233 ( 
.A(n_75),
.B(n_234),
.Y(n_233)
);

BUFx6f_ASAP7_75t_L g76 ( 
.A(n_77),
.Y(n_76)
);

OAI22xp5_ASAP7_75t_SL g424 ( 
.A1(n_78),
.A2(n_79),
.B1(n_425),
.B2(n_426),
.Y(n_424)
);

INVx2_ASAP7_75t_L g78 ( 
.A(n_79),
.Y(n_78)
);

HB1xp67_ASAP7_75t_L g285 ( 
.A(n_80),
.Y(n_285)
);

INVx4_ASAP7_75t_L g80 ( 
.A(n_81),
.Y(n_80)
);

INVx4_ASAP7_75t_L g102 ( 
.A(n_81),
.Y(n_102)
);

BUFx6f_ASAP7_75t_L g81 ( 
.A(n_82),
.Y(n_81)
);

BUFx6f_ASAP7_75t_L g141 ( 
.A(n_82),
.Y(n_141)
);

HB1xp67_ASAP7_75t_L g83 ( 
.A(n_84),
.Y(n_83)
);

XNOR2xp5_ASAP7_75t_L g84 ( 
.A(n_85),
.B(n_93),
.Y(n_84)
);

MAJIxp5_ASAP7_75t_L g166 ( 
.A(n_85),
.B(n_103),
.C(n_104),
.Y(n_166)
);

OAI21xp5_ASAP7_75t_L g268 ( 
.A1(n_85),
.A2(n_269),
.B(n_270),
.Y(n_268)
);

OAI22xp5_ASAP7_75t_L g85 ( 
.A1(n_86),
.A2(n_87),
.B1(n_90),
.B2(n_91),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g121 ( 
.A(n_86),
.B(n_122),
.Y(n_121)
);

INVx2_ASAP7_75t_SL g87 ( 
.A(n_88),
.Y(n_87)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_89),
.Y(n_88)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_89),
.Y(n_111)
);

INVx2_ASAP7_75t_L g271 ( 
.A(n_91),
.Y(n_271)
);

INVx2_ASAP7_75t_L g91 ( 
.A(n_92),
.Y(n_91)
);

OAI22xp5_ASAP7_75t_L g93 ( 
.A1(n_94),
.A2(n_100),
.B1(n_103),
.B2(n_104),
.Y(n_93)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_94),
.Y(n_104)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_96),
.Y(n_95)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_97),
.Y(n_96)
);

INVx5_ASAP7_75t_L g97 ( 
.A(n_98),
.Y(n_97)
);

BUFx6f_ASAP7_75t_L g98 ( 
.A(n_99),
.Y(n_98)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_100),
.Y(n_103)
);

BUFx2_ASAP7_75t_L g101 ( 
.A(n_102),
.Y(n_101)
);

HB1xp67_ASAP7_75t_L g105 ( 
.A(n_106),
.Y(n_105)
);

XNOR2xp5_ASAP7_75t_L g406 ( 
.A(n_106),
.B(n_146),
.Y(n_406)
);

XOR2xp5_ASAP7_75t_L g106 ( 
.A(n_107),
.B(n_117),
.Y(n_106)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_108),
.Y(n_107)
);

MAJIxp5_ASAP7_75t_L g199 ( 
.A(n_108),
.B(n_118),
.C(n_131),
.Y(n_199)
);

OAI22xp5_ASAP7_75t_L g108 ( 
.A1(n_109),
.A2(n_113),
.B1(n_114),
.B2(n_116),
.Y(n_108)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_109),
.Y(n_116)
);

INVx2_ASAP7_75t_L g112 ( 
.A(n_110),
.Y(n_112)
);

AOI22xp5_ASAP7_75t_L g208 ( 
.A1(n_110),
.A2(n_112),
.B1(n_209),
.B2(n_210),
.Y(n_208)
);

AND2x2_ASAP7_75t_L g286 ( 
.A(n_110),
.B(n_287),
.Y(n_286)
);

XNOR2xp5_ASAP7_75t_L g312 ( 
.A(n_110),
.B(n_288),
.Y(n_312)
);

MAJIxp5_ASAP7_75t_L g446 ( 
.A(n_112),
.B(n_209),
.C(n_447),
.Y(n_446)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_114),
.Y(n_113)
);

OAI22xp5_ASAP7_75t_L g117 ( 
.A1(n_118),
.A2(n_119),
.B1(n_131),
.B2(n_132),
.Y(n_117)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_119),
.Y(n_118)
);

MAJIxp5_ASAP7_75t_L g119 ( 
.A(n_120),
.B(n_124),
.C(n_129),
.Y(n_119)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_121),
.Y(n_120)
);

XOR2x2_ASAP7_75t_L g162 ( 
.A(n_121),
.B(n_163),
.Y(n_162)
);

INVx2_ASAP7_75t_L g364 ( 
.A(n_122),
.Y(n_364)
);

INVx4_ASAP7_75t_L g122 ( 
.A(n_123),
.Y(n_122)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_125),
.Y(n_124)
);

AOI22xp5_ASAP7_75t_L g163 ( 
.A1(n_125),
.A2(n_126),
.B1(n_129),
.B2(n_164),
.Y(n_163)
);

OAI22xp5_ASAP7_75t_L g437 ( 
.A1(n_125),
.A2(n_438),
.B1(n_439),
.B2(n_441),
.Y(n_437)
);

INVx1_ASAP7_75t_L g441 ( 
.A(n_125),
.Y(n_441)
);

INVx2_ASAP7_75t_L g125 ( 
.A(n_126),
.Y(n_125)
);

BUFx6f_ASAP7_75t_L g127 ( 
.A(n_128),
.Y(n_127)
);

INVx2_ASAP7_75t_L g174 ( 
.A(n_128),
.Y(n_174)
);

BUFx6f_ASAP7_75t_L g222 ( 
.A(n_128),
.Y(n_222)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_129),
.Y(n_164)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_132),
.Y(n_131)
);

XNOR2xp5_ASAP7_75t_L g132 ( 
.A(n_133),
.B(n_138),
.Y(n_132)
);

OAI22x1_ASAP7_75t_L g214 ( 
.A1(n_133),
.A2(n_142),
.B1(n_215),
.B2(n_216),
.Y(n_214)
);

INVx3_ASAP7_75t_L g134 ( 
.A(n_135),
.Y(n_134)
);

INVx2_ASAP7_75t_L g135 ( 
.A(n_136),
.Y(n_135)
);

BUFx6f_ASAP7_75t_L g136 ( 
.A(n_137),
.Y(n_136)
);

XNOR2x1_ASAP7_75t_L g138 ( 
.A(n_139),
.B(n_142),
.Y(n_138)
);

AND2x2_ASAP7_75t_L g215 ( 
.A(n_139),
.B(n_142),
.Y(n_215)
);

HB1xp67_ASAP7_75t_L g216 ( 
.A(n_139),
.Y(n_216)
);

INVx6_ASAP7_75t_L g140 ( 
.A(n_141),
.Y(n_140)
);

INVx3_ASAP7_75t_L g322 ( 
.A(n_141),
.Y(n_322)
);

INVx2_ASAP7_75t_L g143 ( 
.A(n_144),
.Y(n_143)
);

HB1xp67_ASAP7_75t_L g145 ( 
.A(n_146),
.Y(n_145)
);

XOR2xp5_ASAP7_75t_L g146 ( 
.A(n_147),
.B(n_165),
.Y(n_146)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_147),
.Y(n_202)
);

MAJIxp5_ASAP7_75t_L g147 ( 
.A(n_148),
.B(n_161),
.C(n_162),
.Y(n_147)
);

XNOR2xp5_ASAP7_75t_L g400 ( 
.A(n_148),
.B(n_162),
.Y(n_400)
);

MAJIxp5_ASAP7_75t_L g148 ( 
.A(n_149),
.B(n_151),
.C(n_156),
.Y(n_148)
);

XNOR2x1_ASAP7_75t_L g273 ( 
.A(n_149),
.B(n_207),
.Y(n_273)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_152),
.Y(n_151)
);

BUFx2_ASAP7_75t_L g207 ( 
.A(n_152),
.Y(n_207)
);

INVx1_ASAP7_75t_L g447 ( 
.A(n_152),
.Y(n_447)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_154),
.Y(n_153)
);

BUFx6f_ASAP7_75t_L g154 ( 
.A(n_155),
.Y(n_154)
);

INVx4_ASAP7_75t_L g359 ( 
.A(n_155),
.Y(n_359)
);

XOR2xp5_ASAP7_75t_SL g272 ( 
.A(n_156),
.B(n_273),
.Y(n_272)
);

INVx3_ASAP7_75t_L g157 ( 
.A(n_158),
.Y(n_157)
);

INVx6_ASAP7_75t_L g158 ( 
.A(n_159),
.Y(n_158)
);

BUFx6f_ASAP7_75t_L g159 ( 
.A(n_160),
.Y(n_159)
);

INVx1_ASAP7_75t_L g399 ( 
.A(n_161),
.Y(n_399)
);

XNOR2xp5_ASAP7_75t_L g165 ( 
.A(n_166),
.B(n_167),
.Y(n_165)
);

HB1xp67_ASAP7_75t_L g204 ( 
.A(n_166),
.Y(n_204)
);

BUFx2_ASAP7_75t_SL g203 ( 
.A(n_167),
.Y(n_203)
);

XNOR2x1_ASAP7_75t_L g167 ( 
.A(n_168),
.B(n_170),
.Y(n_167)
);

INVxp67_ASAP7_75t_SL g195 ( 
.A(n_168),
.Y(n_195)
);

AOI22xp5_ASAP7_75t_L g170 ( 
.A1(n_171),
.A2(n_172),
.B1(n_175),
.B2(n_177),
.Y(n_170)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_172),
.Y(n_171)
);

INVx1_ASAP7_75t_SL g196 ( 
.A(n_172),
.Y(n_196)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_174),
.Y(n_173)
);

INVx4_ASAP7_75t_L g317 ( 
.A(n_174),
.Y(n_317)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_175),
.Y(n_177)
);

HB1xp67_ASAP7_75t_L g198 ( 
.A(n_175),
.Y(n_198)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_179),
.Y(n_178)
);

XOR2xp5_ASAP7_75t_L g179 ( 
.A(n_180),
.B(n_200),
.Y(n_179)
);

MAJx2_ASAP7_75t_L g418 ( 
.A(n_180),
.B(n_419),
.C(n_420),
.Y(n_418)
);

XOR2xp5_ASAP7_75t_L g180 ( 
.A(n_181),
.B(n_199),
.Y(n_180)
);

XNOR2xp5_ASAP7_75t_L g181 ( 
.A(n_182),
.B(n_194),
.Y(n_181)
);

INVx1_ASAP7_75t_L g461 ( 
.A(n_182),
.Y(n_461)
);

XNOR2xp5_ASAP7_75t_SL g182 ( 
.A(n_183),
.B(n_184),
.Y(n_182)
);

A2O1A1Ixp33_ASAP7_75t_L g454 ( 
.A1(n_183),
.A2(n_190),
.B(n_455),
.C(n_456),
.Y(n_454)
);

AOI22xp5_ASAP7_75t_L g184 ( 
.A1(n_185),
.A2(n_190),
.B1(n_192),
.B2(n_193),
.Y(n_184)
);

INVxp67_ASAP7_75t_L g455 ( 
.A(n_185),
.Y(n_455)
);

NAND2xp5_ASAP7_75t_L g456 ( 
.A(n_185),
.B(n_193),
.Y(n_456)
);

INVx2_ASAP7_75t_L g186 ( 
.A(n_187),
.Y(n_186)
);

INVx3_ASAP7_75t_L g187 ( 
.A(n_188),
.Y(n_187)
);

BUFx6f_ASAP7_75t_L g188 ( 
.A(n_189),
.Y(n_188)
);

BUFx3_ASAP7_75t_L g252 ( 
.A(n_189),
.Y(n_252)
);

INVx2_ASAP7_75t_L g193 ( 
.A(n_190),
.Y(n_193)
);

OAI22xp5_ASAP7_75t_L g448 ( 
.A1(n_190),
.A2(n_193),
.B1(n_449),
.B2(n_450),
.Y(n_448)
);

MAJx2_ASAP7_75t_L g460 ( 
.A(n_194),
.B(n_199),
.C(n_461),
.Y(n_460)
);

MAJx2_ASAP7_75t_L g194 ( 
.A(n_195),
.B(n_196),
.C(n_197),
.Y(n_194)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_198),
.Y(n_197)
);

XNOR2xp5_ASAP7_75t_L g200 ( 
.A(n_201),
.B(n_205),
.Y(n_200)
);

MAJIxp5_ASAP7_75t_L g201 ( 
.A(n_202),
.B(n_203),
.C(n_204),
.Y(n_201)
);

MAJIxp5_ASAP7_75t_L g419 ( 
.A(n_202),
.B(n_203),
.C(n_204),
.Y(n_419)
);

INVx1_ASAP7_75t_L g420 ( 
.A(n_205),
.Y(n_420)
);

XOR2x2_ASAP7_75t_L g205 ( 
.A(n_206),
.B(n_213),
.Y(n_205)
);

MAJx2_ASAP7_75t_L g458 ( 
.A(n_206),
.B(n_214),
.C(n_217),
.Y(n_458)
);

XNOR2xp5_ASAP7_75t_L g206 ( 
.A(n_207),
.B(n_208),
.Y(n_206)
);

INVx2_ASAP7_75t_L g209 ( 
.A(n_210),
.Y(n_209)
);

BUFx3_ASAP7_75t_L g211 ( 
.A(n_212),
.Y(n_211)
);

XOR2xp5_ASAP7_75t_L g213 ( 
.A(n_214),
.B(n_217),
.Y(n_213)
);

XNOR2x1_ASAP7_75t_L g217 ( 
.A(n_218),
.B(n_220),
.Y(n_217)
);

AOI22xp5_ASAP7_75t_L g426 ( 
.A1(n_218),
.A2(n_219),
.B1(n_427),
.B2(n_428),
.Y(n_426)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_219),
.Y(n_218)
);

INVx1_ASAP7_75t_SL g294 ( 
.A(n_219),
.Y(n_294)
);

MAJIxp5_ASAP7_75t_L g433 ( 
.A(n_219),
.B(n_224),
.C(n_225),
.Y(n_433)
);

OAI22xp5_ASAP7_75t_L g220 ( 
.A1(n_221),
.A2(n_223),
.B1(n_224),
.B2(n_225),
.Y(n_220)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_221),
.Y(n_224)
);

INVx2_ASAP7_75t_L g225 ( 
.A(n_223),
.Y(n_225)
);

AOI21xp5_ASAP7_75t_SL g226 ( 
.A1(n_227),
.A2(n_388),
.B(n_407),
.Y(n_226)
);

HB1xp67_ASAP7_75t_L g227 ( 
.A(n_228),
.Y(n_227)
);

OAI21xp5_ASAP7_75t_L g228 ( 
.A1(n_229),
.A2(n_295),
.B(n_386),
.Y(n_228)
);

AND2x2_ASAP7_75t_L g229 ( 
.A(n_230),
.B(n_274),
.Y(n_229)
);

INVx1_ASAP7_75t_L g387 ( 
.A(n_230),
.Y(n_387)
);

XNOR2xp5_ASAP7_75t_L g230 ( 
.A(n_231),
.B(n_256),
.Y(n_230)
);

XOR2xp5_ASAP7_75t_L g231 ( 
.A(n_232),
.B(n_253),
.Y(n_231)
);

HB1xp67_ASAP7_75t_L g394 ( 
.A(n_232),
.Y(n_394)
);

MAJIxp5_ASAP7_75t_L g232 ( 
.A(n_233),
.B(n_236),
.C(n_239),
.Y(n_232)
);

XNOR2xp5_ASAP7_75t_SL g276 ( 
.A(n_233),
.B(n_277),
.Y(n_276)
);

AOI22xp5_ASAP7_75t_L g277 ( 
.A1(n_236),
.A2(n_237),
.B1(n_239),
.B2(n_278),
.Y(n_277)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_237),
.Y(n_236)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_239),
.Y(n_278)
);

MAJIxp5_ASAP7_75t_L g239 ( 
.A(n_240),
.B(n_245),
.C(n_248),
.Y(n_239)
);

OAI22xp5_ASAP7_75t_L g378 ( 
.A1(n_240),
.A2(n_241),
.B1(n_248),
.B2(n_249),
.Y(n_378)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_241),
.Y(n_240)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_243),
.Y(n_242)
);

BUFx5_ASAP7_75t_L g243 ( 
.A(n_244),
.Y(n_243)
);

BUFx6f_ASAP7_75t_L g267 ( 
.A(n_244),
.Y(n_267)
);

XNOR2xp5_ASAP7_75t_L g377 ( 
.A(n_245),
.B(n_378),
.Y(n_377)
);

INVx2_ASAP7_75t_L g246 ( 
.A(n_247),
.Y(n_246)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_249),
.Y(n_248)
);

INVx5_ASAP7_75t_L g250 ( 
.A(n_251),
.Y(n_250)
);

INVx5_ASAP7_75t_L g251 ( 
.A(n_252),
.Y(n_251)
);

INVx1_ASAP7_75t_L g393 ( 
.A(n_253),
.Y(n_393)
);

XNOR2x1_ASAP7_75t_L g253 ( 
.A(n_254),
.B(n_255),
.Y(n_253)
);

INVx1_ASAP7_75t_L g392 ( 
.A(n_256),
.Y(n_392)
);

XOR2xp5_ASAP7_75t_L g256 ( 
.A(n_257),
.B(n_272),
.Y(n_256)
);

XNOR2xp5_ASAP7_75t_L g257 ( 
.A(n_258),
.B(n_268),
.Y(n_257)
);

MAJx2_ASAP7_75t_L g397 ( 
.A(n_258),
.B(n_268),
.C(n_272),
.Y(n_397)
);

MAJIxp5_ASAP7_75t_L g258 ( 
.A(n_259),
.B(n_261),
.C(n_264),
.Y(n_258)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_260),
.Y(n_259)
);

XNOR2xp5_ASAP7_75t_SL g280 ( 
.A(n_260),
.B(n_281),
.Y(n_280)
);

XNOR2xp5_ASAP7_75t_L g281 ( 
.A(n_261),
.B(n_264),
.Y(n_281)
);

BUFx6f_ASAP7_75t_L g262 ( 
.A(n_263),
.Y(n_262)
);

BUFx2_ASAP7_75t_L g265 ( 
.A(n_266),
.Y(n_265)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_267),
.Y(n_266)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_275),
.Y(n_274)
);

NAND2xp5_ASAP7_75t_L g386 ( 
.A(n_275),
.B(n_387),
.Y(n_386)
);

MAJIxp5_ASAP7_75t_L g275 ( 
.A(n_276),
.B(n_279),
.C(n_282),
.Y(n_275)
);

XNOR2xp5_ASAP7_75t_L g381 ( 
.A(n_276),
.B(n_382),
.Y(n_381)
);

AOI22xp5_ASAP7_75t_L g382 ( 
.A1(n_279),
.A2(n_280),
.B1(n_282),
.B2(n_383),
.Y(n_382)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_280),
.Y(n_279)
);

INVx1_ASAP7_75t_L g383 ( 
.A(n_282),
.Y(n_383)
);

MAJIxp5_ASAP7_75t_L g282 ( 
.A(n_283),
.B(n_286),
.C(n_292),
.Y(n_282)
);

OAI22xp5_ASAP7_75t_L g373 ( 
.A1(n_283),
.A2(n_284),
.B1(n_292),
.B2(n_374),
.Y(n_373)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_284),
.Y(n_283)
);

XNOR2xp5_ASAP7_75t_L g372 ( 
.A(n_286),
.B(n_373),
.Y(n_372)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_288),
.Y(n_287)
);

INVx2_ASAP7_75t_L g289 ( 
.A(n_290),
.Y(n_289)
);

INVx2_ASAP7_75t_L g290 ( 
.A(n_291),
.Y(n_290)
);

INVxp67_ASAP7_75t_SL g374 ( 
.A(n_292),
.Y(n_374)
);

AOI21xp5_ASAP7_75t_L g295 ( 
.A1(n_296),
.A2(n_380),
.B(n_385),
.Y(n_295)
);

OAI21xp5_ASAP7_75t_L g296 ( 
.A1(n_297),
.A2(n_369),
.B(n_379),
.Y(n_296)
);

AOI21x1_ASAP7_75t_L g297 ( 
.A1(n_298),
.A2(n_339),
.B(n_368),
.Y(n_297)
);

NAND2xp5_ASAP7_75t_L g298 ( 
.A(n_299),
.B(n_331),
.Y(n_298)
);

OAI22xp33_ASAP7_75t_L g299 ( 
.A1(n_300),
.A2(n_313),
.B1(n_329),
.B2(n_330),
.Y(n_299)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_300),
.Y(n_329)
);

AOI221xp5_ASAP7_75t_L g368 ( 
.A1(n_300),
.A2(n_313),
.B1(n_329),
.B2(n_330),
.C(n_331),
.Y(n_368)
);

AOI22xp5_ASAP7_75t_L g300 ( 
.A1(n_301),
.A2(n_302),
.B1(n_311),
.B2(n_312),
.Y(n_300)
);

MAJIxp5_ASAP7_75t_L g370 ( 
.A(n_301),
.B(n_312),
.C(n_330),
.Y(n_370)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_302),
.Y(n_301)
);

NAND2xp5_ASAP7_75t_L g302 ( 
.A(n_303),
.B(n_307),
.Y(n_302)
);

XNOR2xp5_ASAP7_75t_L g333 ( 
.A(n_303),
.B(n_307),
.Y(n_333)
);

NOR2xp33_ASAP7_75t_L g303 ( 
.A(n_304),
.B(n_305),
.Y(n_303)
);

INVx8_ASAP7_75t_L g305 ( 
.A(n_306),
.Y(n_305)
);

INVx8_ASAP7_75t_L g349 ( 
.A(n_306),
.Y(n_349)
);

NOR2xp33_ASAP7_75t_L g307 ( 
.A(n_308),
.B(n_309),
.Y(n_307)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_310),
.Y(n_309)
);

INVx6_ASAP7_75t_L g346 ( 
.A(n_310),
.Y(n_346)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_312),
.Y(n_311)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_313),
.Y(n_330)
);

XNOR2xp5_ASAP7_75t_L g313 ( 
.A(n_314),
.B(n_318),
.Y(n_313)
);

MAJIxp5_ASAP7_75t_L g376 ( 
.A(n_314),
.B(n_319),
.C(n_323),
.Y(n_376)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_316),
.Y(n_315)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_317),
.Y(n_316)
);

OAI22xp5_ASAP7_75t_L g318 ( 
.A1(n_319),
.A2(n_323),
.B1(n_327),
.B2(n_328),
.Y(n_318)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_319),
.Y(n_327)
);

INVx2_ASAP7_75t_L g320 ( 
.A(n_321),
.Y(n_320)
);

INVx2_ASAP7_75t_L g321 ( 
.A(n_322),
.Y(n_321)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_323),
.Y(n_328)
);

INVx2_ASAP7_75t_SL g324 ( 
.A(n_325),
.Y(n_324)
);

INVx3_ASAP7_75t_L g325 ( 
.A(n_326),
.Y(n_325)
);

MAJIxp5_ASAP7_75t_L g331 ( 
.A(n_332),
.B(n_334),
.C(n_335),
.Y(n_331)
);

OAI22xp5_ASAP7_75t_SL g350 ( 
.A1(n_332),
.A2(n_333),
.B1(n_351),
.B2(n_352),
.Y(n_350)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_333),
.Y(n_332)
);

OAI22xp5_ASAP7_75t_SL g352 ( 
.A1(n_334),
.A2(n_335),
.B1(n_336),
.B2(n_353),
.Y(n_352)
);

CKINVDCx12_ASAP7_75t_R g353 ( 
.A(n_334),
.Y(n_353)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_336),
.Y(n_335)
);

BUFx6f_ASAP7_75t_L g337 ( 
.A(n_338),
.Y(n_337)
);

OAI21xp5_ASAP7_75t_L g339 ( 
.A1(n_340),
.A2(n_354),
.B(n_367),
.Y(n_339)
);

NOR2xp33_ASAP7_75t_L g340 ( 
.A(n_341),
.B(n_350),
.Y(n_340)
);

NAND2xp5_ASAP7_75t_L g367 ( 
.A(n_341),
.B(n_350),
.Y(n_367)
);

NOR2xp33_ASAP7_75t_L g341 ( 
.A(n_342),
.B(n_347),
.Y(n_341)
);

XNOR2xp5_ASAP7_75t_L g356 ( 
.A(n_342),
.B(n_347),
.Y(n_356)
);

INVx3_ASAP7_75t_L g343 ( 
.A(n_344),
.Y(n_343)
);

INVx2_ASAP7_75t_L g344 ( 
.A(n_345),
.Y(n_344)
);

INVx2_ASAP7_75t_L g345 ( 
.A(n_346),
.Y(n_345)
);

INVx5_ASAP7_75t_L g348 ( 
.A(n_349),
.Y(n_348)
);

INVx1_ASAP7_75t_L g351 ( 
.A(n_352),
.Y(n_351)
);

AOI21xp5_ASAP7_75t_L g354 ( 
.A1(n_355),
.A2(n_360),
.B(n_366),
.Y(n_354)
);

NAND2xp5_ASAP7_75t_SL g355 ( 
.A(n_356),
.B(n_357),
.Y(n_355)
);

NOR2xp33_ASAP7_75t_L g366 ( 
.A(n_356),
.B(n_357),
.Y(n_366)
);

BUFx3_ASAP7_75t_L g358 ( 
.A(n_359),
.Y(n_358)
);

NOR2xp33_ASAP7_75t_L g360 ( 
.A(n_361),
.B(n_365),
.Y(n_360)
);

INVx2_ASAP7_75t_L g362 ( 
.A(n_363),
.Y(n_362)
);

INVx2_ASAP7_75t_L g363 ( 
.A(n_364),
.Y(n_363)
);

AND2x2_ASAP7_75t_L g369 ( 
.A(n_370),
.B(n_371),
.Y(n_369)
);

OR2x2_ASAP7_75t_L g379 ( 
.A(n_370),
.B(n_371),
.Y(n_379)
);

XOR2xp5_ASAP7_75t_L g371 ( 
.A(n_372),
.B(n_375),
.Y(n_371)
);

MAJIxp5_ASAP7_75t_L g384 ( 
.A(n_372),
.B(n_376),
.C(n_377),
.Y(n_384)
);

XNOR2xp5_ASAP7_75t_L g375 ( 
.A(n_376),
.B(n_377),
.Y(n_375)
);

NAND2xp5_ASAP7_75t_SL g380 ( 
.A(n_381),
.B(n_384),
.Y(n_380)
);

NOR2xp67_ASAP7_75t_SL g385 ( 
.A(n_381),
.B(n_384),
.Y(n_385)
);

HB1xp67_ASAP7_75t_L g388 ( 
.A(n_389),
.Y(n_388)
);

NOR2x1_ASAP7_75t_L g389 ( 
.A(n_390),
.B(n_403),
.Y(n_389)
);

NOR2xp67_ASAP7_75t_L g390 ( 
.A(n_391),
.B(n_395),
.Y(n_390)
);

NAND2xp5_ASAP7_75t_L g409 ( 
.A(n_391),
.B(n_395),
.Y(n_409)
);

MAJx2_ASAP7_75t_L g391 ( 
.A(n_392),
.B(n_393),
.C(n_394),
.Y(n_391)
);

XNOR2x1_ASAP7_75t_L g395 ( 
.A(n_396),
.B(n_401),
.Y(n_395)
);

XNOR2xp5_ASAP7_75t_L g396 ( 
.A(n_397),
.B(n_398),
.Y(n_396)
);

MAJIxp5_ASAP7_75t_L g404 ( 
.A(n_397),
.B(n_398),
.C(n_401),
.Y(n_404)
);

XNOR2x2_ASAP7_75t_L g398 ( 
.A(n_399),
.B(n_400),
.Y(n_398)
);

OAI21xp5_ASAP7_75t_L g408 ( 
.A1(n_403),
.A2(n_409),
.B(n_410),
.Y(n_408)
);

AND2x2_ASAP7_75t_L g403 ( 
.A(n_404),
.B(n_405),
.Y(n_403)
);

OR2x2_ASAP7_75t_L g410 ( 
.A(n_404),
.B(n_405),
.Y(n_410)
);

HB1xp67_ASAP7_75t_L g407 ( 
.A(n_408),
.Y(n_407)
);

INVx1_ASAP7_75t_L g411 ( 
.A(n_412),
.Y(n_411)
);

NAND4xp25_ASAP7_75t_SL g463 ( 
.A(n_412),
.B(n_415),
.C(n_464),
.D(n_465),
.Y(n_463)
);

HB1xp67_ASAP7_75t_L g412 ( 
.A(n_413),
.Y(n_412)
);

OR2x2_ASAP7_75t_L g415 ( 
.A(n_416),
.B(n_462),
.Y(n_415)
);

INVxp33_ASAP7_75t_L g416 ( 
.A(n_417),
.Y(n_416)
);

NAND2xp5_ASAP7_75t_L g417 ( 
.A(n_418),
.B(n_421),
.Y(n_417)
);

NOR2xp67_ASAP7_75t_L g462 ( 
.A(n_418),
.B(n_421),
.Y(n_462)
);

XNOR2x1_ASAP7_75t_L g421 ( 
.A(n_422),
.B(n_460),
.Y(n_421)
);

XNOR2x1_ASAP7_75t_L g422 ( 
.A(n_423),
.B(n_443),
.Y(n_422)
);

XOR2x2_ASAP7_75t_L g423 ( 
.A(n_424),
.B(n_431),
.Y(n_423)
);

INVx1_ASAP7_75t_L g425 ( 
.A(n_426),
.Y(n_425)
);

INVx1_ASAP7_75t_L g427 ( 
.A(n_428),
.Y(n_427)
);

INVx1_ASAP7_75t_L g429 ( 
.A(n_430),
.Y(n_429)
);

OAI22xp5_ASAP7_75t_L g431 ( 
.A1(n_432),
.A2(n_433),
.B1(n_434),
.B2(n_442),
.Y(n_431)
);

INVx1_ASAP7_75t_L g432 ( 
.A(n_433),
.Y(n_432)
);

INVx1_ASAP7_75t_L g442 ( 
.A(n_434),
.Y(n_442)
);

XNOR2x1_ASAP7_75t_L g434 ( 
.A(n_435),
.B(n_437),
.Y(n_434)
);

INVx1_ASAP7_75t_L g438 ( 
.A(n_439),
.Y(n_438)
);

OAI22x1_ASAP7_75t_L g443 ( 
.A1(n_444),
.A2(n_457),
.B1(n_458),
.B2(n_459),
.Y(n_443)
);

INVx2_ASAP7_75t_L g459 ( 
.A(n_444),
.Y(n_459)
);

XNOR2x1_ASAP7_75t_L g444 ( 
.A(n_445),
.B(n_454),
.Y(n_444)
);

XNOR2xp5_ASAP7_75t_L g445 ( 
.A(n_446),
.B(n_448),
.Y(n_445)
);

INVx1_ASAP7_75t_L g449 ( 
.A(n_450),
.Y(n_449)
);

INVx2_ASAP7_75t_L g451 ( 
.A(n_452),
.Y(n_451)
);

INVx8_ASAP7_75t_L g452 ( 
.A(n_453),
.Y(n_452)
);

INVx1_ASAP7_75t_L g457 ( 
.A(n_458),
.Y(n_457)
);


endmodule