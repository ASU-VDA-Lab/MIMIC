module fake_jpeg_17270_n_394 (n_13, n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_394);

input n_13;
input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_394;

wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_385;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_340;
wire n_381;
wire n_377;
wire n_291;
wire n_236;
wire n_15;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_370;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_327;
wire n_122;
wire n_75;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_39;
wire n_371;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_382;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_14;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_352;
wire n_350;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_389;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_384;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_360;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_378;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_379;
wire n_114;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_356;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_375;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_391;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

BUFx6f_ASAP7_75t_L g14 ( 
.A(n_4),
.Y(n_14)
);

BUFx6f_ASAP7_75t_L g15 ( 
.A(n_13),
.Y(n_15)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_13),
.Y(n_16)
);

INVx2_ASAP7_75t_L g17 ( 
.A(n_12),
.Y(n_17)
);

CKINVDCx16_ASAP7_75t_R g18 ( 
.A(n_12),
.Y(n_18)
);

CKINVDCx14_ASAP7_75t_R g19 ( 
.A(n_13),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_12),
.Y(n_20)
);

BUFx12f_ASAP7_75t_L g21 ( 
.A(n_8),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_11),
.Y(n_22)
);

INVx6_ASAP7_75t_L g23 ( 
.A(n_5),
.Y(n_23)
);

BUFx10_ASAP7_75t_L g24 ( 
.A(n_4),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_10),
.Y(n_25)
);

NOR2xp33_ASAP7_75t_L g26 ( 
.A(n_12),
.B(n_8),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_9),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_11),
.Y(n_28)
);

BUFx12f_ASAP7_75t_L g29 ( 
.A(n_7),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_1),
.Y(n_30)
);

BUFx12f_ASAP7_75t_L g31 ( 
.A(n_0),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_3),
.Y(n_32)
);

INVx2_ASAP7_75t_L g33 ( 
.A(n_10),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_13),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_0),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_9),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_3),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_14),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g101 ( 
.A(n_38),
.Y(n_101)
);

INVx5_ASAP7_75t_L g39 ( 
.A(n_23),
.Y(n_39)
);

INVx3_ASAP7_75t_L g72 ( 
.A(n_39),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_L g40 ( 
.A(n_26),
.B(n_0),
.Y(n_40)
);

AND2x2_ASAP7_75t_L g100 ( 
.A(n_40),
.B(n_47),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g41 ( 
.A(n_26),
.B(n_0),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_SL g73 ( 
.A(n_41),
.B(n_53),
.Y(n_73)
);

INVx8_ASAP7_75t_L g42 ( 
.A(n_23),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g104 ( 
.A(n_42),
.Y(n_104)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_14),
.Y(n_43)
);

INVx3_ASAP7_75t_L g85 ( 
.A(n_43),
.Y(n_85)
);

INVx2_ASAP7_75t_L g44 ( 
.A(n_17),
.Y(n_44)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_44),
.Y(n_69)
);

INVx11_ASAP7_75t_L g45 ( 
.A(n_14),
.Y(n_45)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_45),
.Y(n_84)
);

INVx6_ASAP7_75t_L g46 ( 
.A(n_29),
.Y(n_46)
);

INVx2_ASAP7_75t_L g74 ( 
.A(n_46),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_L g47 ( 
.A(n_16),
.B(n_1),
.Y(n_47)
);

INVx5_ASAP7_75t_L g48 ( 
.A(n_23),
.Y(n_48)
);

INVx3_ASAP7_75t_L g86 ( 
.A(n_48),
.Y(n_86)
);

INVx11_ASAP7_75t_L g49 ( 
.A(n_15),
.Y(n_49)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_49),
.Y(n_112)
);

INVx11_ASAP7_75t_L g50 ( 
.A(n_15),
.Y(n_50)
);

INVx2_ASAP7_75t_L g76 ( 
.A(n_50),
.Y(n_76)
);

INVx11_ASAP7_75t_L g51 ( 
.A(n_15),
.Y(n_51)
);

INVx2_ASAP7_75t_L g88 ( 
.A(n_51),
.Y(n_88)
);

INVx6_ASAP7_75t_L g52 ( 
.A(n_29),
.Y(n_52)
);

INVx2_ASAP7_75t_L g95 ( 
.A(n_52),
.Y(n_95)
);

OR2x2_ASAP7_75t_L g53 ( 
.A(n_18),
.B(n_1),
.Y(n_53)
);

INVx3_ASAP7_75t_L g54 ( 
.A(n_17),
.Y(n_54)
);

INVx3_ASAP7_75t_L g90 ( 
.A(n_54),
.Y(n_90)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_33),
.Y(n_55)
);

CKINVDCx16_ASAP7_75t_R g68 ( 
.A(n_55),
.Y(n_68)
);

INVx8_ASAP7_75t_L g56 ( 
.A(n_29),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_56),
.B(n_57),
.Y(n_82)
);

INVx8_ASAP7_75t_L g57 ( 
.A(n_29),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_19),
.B(n_1),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_L g75 ( 
.A(n_58),
.B(n_63),
.Y(n_75)
);

BUFx5_ASAP7_75t_L g59 ( 
.A(n_24),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_59),
.B(n_61),
.Y(n_97)
);

INVx3_ASAP7_75t_L g60 ( 
.A(n_33),
.Y(n_60)
);

INVx3_ASAP7_75t_L g91 ( 
.A(n_60),
.Y(n_91)
);

CKINVDCx20_ASAP7_75t_R g61 ( 
.A(n_16),
.Y(n_61)
);

BUFx3_ASAP7_75t_L g62 ( 
.A(n_24),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_62),
.B(n_24),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_19),
.B(n_2),
.Y(n_63)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_20),
.Y(n_64)
);

INVx3_ASAP7_75t_L g113 ( 
.A(n_64),
.Y(n_113)
);

AND2x2_ASAP7_75t_SL g65 ( 
.A(n_22),
.B(n_2),
.Y(n_65)
);

MAJIxp5_ASAP7_75t_L g98 ( 
.A(n_65),
.B(n_31),
.C(n_29),
.Y(n_98)
);

INVx11_ASAP7_75t_L g66 ( 
.A(n_20),
.Y(n_66)
);

INVx2_ASAP7_75t_L g96 ( 
.A(n_66),
.Y(n_96)
);

BUFx3_ASAP7_75t_L g67 ( 
.A(n_38),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g129 ( 
.A(n_67),
.B(n_114),
.Y(n_129)
);

AOI22xp33_ASAP7_75t_L g70 ( 
.A1(n_45),
.A2(n_18),
.B1(n_36),
.B2(n_30),
.Y(n_70)
);

OAI22xp5_ASAP7_75t_L g139 ( 
.A1(n_70),
.A2(n_78),
.B1(n_92),
.B2(n_103),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_SL g71 ( 
.A(n_61),
.B(n_36),
.Y(n_71)
);

AND2x2_ASAP7_75t_L g125 ( 
.A(n_71),
.B(n_80),
.Y(n_125)
);

OAI22xp5_ASAP7_75t_L g77 ( 
.A1(n_47),
.A2(n_37),
.B1(n_30),
.B2(n_28),
.Y(n_77)
);

AOI22xp5_ASAP7_75t_L g118 ( 
.A1(n_77),
.A2(n_81),
.B1(n_102),
.B2(n_5),
.Y(n_118)
);

AOI22xp33_ASAP7_75t_L g78 ( 
.A1(n_45),
.A2(n_37),
.B1(n_27),
.B2(n_28),
.Y(n_78)
);

AND2x2_ASAP7_75t_SL g79 ( 
.A(n_55),
.B(n_34),
.Y(n_79)
);

OAI21xp5_ASAP7_75t_SL g138 ( 
.A1(n_79),
.A2(n_108),
.B(n_21),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_L g80 ( 
.A(n_65),
.B(n_34),
.Y(n_80)
);

OAI22xp5_ASAP7_75t_L g81 ( 
.A1(n_42),
.A2(n_39),
.B1(n_48),
.B2(n_50),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_SL g83 ( 
.A(n_65),
.B(n_27),
.Y(n_83)
);

AND2x2_ASAP7_75t_L g167 ( 
.A(n_83),
.B(n_89),
.Y(n_167)
);

OR2x2_ASAP7_75t_L g87 ( 
.A(n_40),
.B(n_32),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_SL g147 ( 
.A(n_87),
.B(n_110),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_SL g89 ( 
.A(n_65),
.B(n_32),
.Y(n_89)
);

OAI22xp33_ASAP7_75t_SL g92 ( 
.A1(n_66),
.A2(n_35),
.B1(n_20),
.B2(n_25),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_L g93 ( 
.A(n_53),
.B(n_22),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_L g119 ( 
.A(n_93),
.B(n_94),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_L g94 ( 
.A(n_53),
.B(n_21),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_L g120 ( 
.A(n_98),
.B(n_111),
.Y(n_120)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_99),
.Y(n_127)
);

OAI22xp5_ASAP7_75t_L g102 ( 
.A1(n_42),
.A2(n_35),
.B1(n_25),
.B2(n_24),
.Y(n_102)
);

AOI22xp33_ASAP7_75t_L g103 ( 
.A1(n_49),
.A2(n_66),
.B1(n_50),
.B2(n_51),
.Y(n_103)
);

AOI22xp33_ASAP7_75t_SL g105 ( 
.A1(n_49),
.A2(n_25),
.B1(n_35),
.B2(n_4),
.Y(n_105)
);

AOI22xp33_ASAP7_75t_SL g126 ( 
.A1(n_105),
.A2(n_117),
.B1(n_46),
.B2(n_52),
.Y(n_126)
);

INVx2_ASAP7_75t_L g106 ( 
.A(n_44),
.Y(n_106)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_106),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_41),
.B(n_24),
.Y(n_107)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_107),
.Y(n_131)
);

AND2x2_ASAP7_75t_L g108 ( 
.A(n_54),
.B(n_2),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_58),
.B(n_2),
.Y(n_109)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_109),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_63),
.B(n_3),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_62),
.B(n_3),
.Y(n_111)
);

BUFx3_ASAP7_75t_L g114 ( 
.A(n_38),
.Y(n_114)
);

INVx1_ASAP7_75t_SL g115 ( 
.A(n_43),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_L g158 ( 
.A(n_115),
.B(n_5),
.Y(n_158)
);

INVx3_ASAP7_75t_L g116 ( 
.A(n_60),
.Y(n_116)
);

INVx3_ASAP7_75t_L g146 ( 
.A(n_116),
.Y(n_146)
);

AOI22xp33_ASAP7_75t_SL g117 ( 
.A1(n_51),
.A2(n_4),
.B1(n_5),
.B2(n_6),
.Y(n_117)
);

AOI22xp33_ASAP7_75t_L g179 ( 
.A1(n_118),
.A2(n_151),
.B1(n_86),
.B2(n_72),
.Y(n_179)
);

INVx2_ASAP7_75t_L g121 ( 
.A(n_106),
.Y(n_121)
);

INVx2_ASAP7_75t_L g205 ( 
.A(n_121),
.Y(n_205)
);

INVx2_ASAP7_75t_L g122 ( 
.A(n_69),
.Y(n_122)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_122),
.Y(n_189)
);

INVx2_ASAP7_75t_L g123 ( 
.A(n_74),
.Y(n_123)
);

INVx2_ASAP7_75t_L g211 ( 
.A(n_123),
.Y(n_211)
);

AOI22xp33_ASAP7_75t_L g124 ( 
.A1(n_102),
.A2(n_52),
.B1(n_46),
.B2(n_56),
.Y(n_124)
);

OAI22xp5_ASAP7_75t_SL g172 ( 
.A1(n_124),
.A2(n_165),
.B1(n_86),
.B2(n_72),
.Y(n_172)
);

AOI22xp33_ASAP7_75t_SL g188 ( 
.A1(n_126),
.A2(n_132),
.B1(n_90),
.B2(n_91),
.Y(n_188)
);

BUFx3_ASAP7_75t_L g130 ( 
.A(n_104),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_L g206 ( 
.A(n_130),
.B(n_145),
.Y(n_206)
);

AOI22xp33_ASAP7_75t_SL g132 ( 
.A1(n_85),
.A2(n_56),
.B1(n_57),
.B2(n_7),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_L g133 ( 
.A(n_100),
.B(n_21),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_SL g173 ( 
.A(n_133),
.B(n_152),
.Y(n_173)
);

BUFx12f_ASAP7_75t_L g134 ( 
.A(n_101),
.Y(n_134)
);

INVx5_ASAP7_75t_L g196 ( 
.A(n_134),
.Y(n_196)
);

INVx6_ASAP7_75t_L g135 ( 
.A(n_101),
.Y(n_135)
);

INVx8_ASAP7_75t_L g174 ( 
.A(n_135),
.Y(n_174)
);

INVx2_ASAP7_75t_L g136 ( 
.A(n_74),
.Y(n_136)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_136),
.Y(n_198)
);

OAI32xp33_ASAP7_75t_L g137 ( 
.A1(n_80),
.A2(n_64),
.A3(n_43),
.B1(n_62),
.B2(n_59),
.Y(n_137)
);

CKINVDCx14_ASAP7_75t_R g195 ( 
.A(n_137),
.Y(n_195)
);

AO21x1_ASAP7_75t_L g175 ( 
.A1(n_138),
.A2(n_154),
.B(n_75),
.Y(n_175)
);

AOI22xp5_ASAP7_75t_L g140 ( 
.A1(n_100),
.A2(n_57),
.B1(n_64),
.B2(n_7),
.Y(n_140)
);

OAI22xp5_ASAP7_75t_L g200 ( 
.A1(n_140),
.A2(n_112),
.B1(n_10),
.B2(n_11),
.Y(n_200)
);

AND2x2_ASAP7_75t_SL g142 ( 
.A(n_94),
.B(n_31),
.Y(n_142)
);

OAI21xp5_ASAP7_75t_SL g190 ( 
.A1(n_142),
.A2(n_108),
.B(n_68),
.Y(n_190)
);

BUFx6f_ASAP7_75t_L g143 ( 
.A(n_85),
.Y(n_143)
);

INVx3_ASAP7_75t_L g194 ( 
.A(n_143),
.Y(n_194)
);

BUFx6f_ASAP7_75t_L g144 ( 
.A(n_113),
.Y(n_144)
);

CKINVDCx20_ASAP7_75t_R g177 ( 
.A(n_144),
.Y(n_177)
);

BUFx6f_ASAP7_75t_L g145 ( 
.A(n_113),
.Y(n_145)
);

INVx2_ASAP7_75t_L g148 ( 
.A(n_95),
.Y(n_148)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_148),
.Y(n_208)
);

BUFx2_ASAP7_75t_L g149 ( 
.A(n_76),
.Y(n_149)
);

NOR2xp33_ASAP7_75t_L g171 ( 
.A(n_149),
.B(n_150),
.Y(n_171)
);

INVx4_ASAP7_75t_L g150 ( 
.A(n_69),
.Y(n_150)
);

OAI22xp33_ASAP7_75t_SL g151 ( 
.A1(n_115),
.A2(n_31),
.B1(n_21),
.B2(n_7),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_SL g152 ( 
.A(n_100),
.B(n_31),
.Y(n_152)
);

INVx2_ASAP7_75t_L g153 ( 
.A(n_95),
.Y(n_153)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_153),
.Y(n_213)
);

OR2x2_ASAP7_75t_SL g154 ( 
.A(n_87),
.B(n_31),
.Y(n_154)
);

INVx2_ASAP7_75t_L g155 ( 
.A(n_76),
.Y(n_155)
);

INVxp67_ASAP7_75t_L g187 ( 
.A(n_155),
.Y(n_187)
);

BUFx6f_ASAP7_75t_L g156 ( 
.A(n_104),
.Y(n_156)
);

INVxp67_ASAP7_75t_L g197 ( 
.A(n_156),
.Y(n_197)
);

INVx2_ASAP7_75t_L g157 ( 
.A(n_88),
.Y(n_157)
);

NOR2xp33_ASAP7_75t_L g178 ( 
.A(n_157),
.B(n_159),
.Y(n_178)
);

CKINVDCx16_ASAP7_75t_R g202 ( 
.A(n_158),
.Y(n_202)
);

NOR2xp33_ASAP7_75t_L g159 ( 
.A(n_97),
.B(n_6),
.Y(n_159)
);

NOR2xp33_ASAP7_75t_L g160 ( 
.A(n_75),
.B(n_79),
.Y(n_160)
);

NOR2xp33_ASAP7_75t_L g180 ( 
.A(n_160),
.B(n_161),
.Y(n_180)
);

INVx2_ASAP7_75t_L g161 ( 
.A(n_88),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_L g162 ( 
.A(n_93),
.B(n_6),
.Y(n_162)
);

NOR2xp33_ASAP7_75t_SL g186 ( 
.A(n_162),
.B(n_166),
.Y(n_186)
);

HB1xp67_ASAP7_75t_L g163 ( 
.A(n_84),
.Y(n_163)
);

NOR2xp33_ASAP7_75t_L g183 ( 
.A(n_163),
.B(n_164),
.Y(n_183)
);

INVx3_ASAP7_75t_L g164 ( 
.A(n_90),
.Y(n_164)
);

AOI22xp33_ASAP7_75t_L g165 ( 
.A1(n_81),
.A2(n_6),
.B1(n_8),
.B2(n_9),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_L g166 ( 
.A(n_73),
.B(n_8),
.Y(n_166)
);

INVx2_ASAP7_75t_L g168 ( 
.A(n_96),
.Y(n_168)
);

NOR2xp33_ASAP7_75t_L g185 ( 
.A(n_168),
.B(n_114),
.Y(n_185)
);

NOR2x1_ASAP7_75t_L g169 ( 
.A(n_154),
.B(n_73),
.Y(n_169)
);

OAI21xp5_ASAP7_75t_L g249 ( 
.A1(n_169),
.A2(n_182),
.B(n_214),
.Y(n_249)
);

NAND2xp5_ASAP7_75t_L g170 ( 
.A(n_142),
.B(n_119),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_L g220 ( 
.A(n_170),
.B(n_176),
.Y(n_220)
);

AOI22xp33_ASAP7_75t_L g230 ( 
.A1(n_172),
.A2(n_179),
.B1(n_174),
.B2(n_194),
.Y(n_230)
);

NOR2xp33_ASAP7_75t_SL g234 ( 
.A(n_175),
.B(n_191),
.Y(n_234)
);

NAND2xp5_ASAP7_75t_L g176 ( 
.A(n_142),
.B(n_79),
.Y(n_176)
);

AOI22xp5_ASAP7_75t_L g181 ( 
.A1(n_120),
.A2(n_139),
.B1(n_137),
.B2(n_118),
.Y(n_181)
);

OAI22xp5_ASAP7_75t_L g246 ( 
.A1(n_181),
.A2(n_188),
.B1(n_199),
.B2(n_201),
.Y(n_246)
);

NAND2xp33_ASAP7_75t_SL g182 ( 
.A(n_150),
.B(n_98),
.Y(n_182)
);

XNOR2xp5_ASAP7_75t_L g184 ( 
.A(n_140),
.B(n_82),
.Y(n_184)
);

XNOR2xp5_ASAP7_75t_SL g237 ( 
.A(n_184),
.B(n_190),
.Y(n_237)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_185),
.Y(n_227)
);

NOR2xp33_ASAP7_75t_L g191 ( 
.A(n_147),
.B(n_91),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_L g192 ( 
.A(n_125),
.B(n_108),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_L g224 ( 
.A(n_192),
.B(n_207),
.Y(n_224)
);

NOR2xp33_ASAP7_75t_L g193 ( 
.A(n_141),
.B(n_116),
.Y(n_193)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_193),
.Y(n_236)
);

AOI22xp5_ASAP7_75t_L g199 ( 
.A1(n_125),
.A2(n_84),
.B1(n_112),
.B2(n_96),
.Y(n_199)
);

AOI22xp5_ASAP7_75t_L g219 ( 
.A1(n_200),
.A2(n_135),
.B1(n_156),
.B2(n_144),
.Y(n_219)
);

AOI22xp5_ASAP7_75t_L g201 ( 
.A1(n_167),
.A2(n_67),
.B1(n_10),
.B2(n_11),
.Y(n_201)
);

NOR2xp33_ASAP7_75t_L g203 ( 
.A(n_131),
.B(n_9),
.Y(n_203)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_203),
.Y(n_239)
);

NOR2xp33_ASAP7_75t_L g204 ( 
.A(n_127),
.B(n_122),
.Y(n_204)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_204),
.Y(n_242)
);

NAND2xp5_ASAP7_75t_SL g207 ( 
.A(n_167),
.B(n_128),
.Y(n_207)
);

NOR2xp33_ASAP7_75t_L g209 ( 
.A(n_146),
.B(n_164),
.Y(n_209)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_209),
.Y(n_245)
);

XOR2xp5_ASAP7_75t_L g210 ( 
.A(n_124),
.B(n_165),
.Y(n_210)
);

MAJx2_ASAP7_75t_L g243 ( 
.A(n_210),
.B(n_175),
.C(n_173),
.Y(n_243)
);

NAND2xp5_ASAP7_75t_L g212 ( 
.A(n_146),
.B(n_168),
.Y(n_212)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_212),
.Y(n_256)
);

OAI21xp33_ASAP7_75t_SL g214 ( 
.A1(n_126),
.A2(n_151),
.B(n_132),
.Y(n_214)
);

NOR2xp33_ASAP7_75t_L g215 ( 
.A(n_149),
.B(n_129),
.Y(n_215)
);

NOR2xp33_ASAP7_75t_L g216 ( 
.A(n_215),
.B(n_143),
.Y(n_216)
);

NOR2xp33_ASAP7_75t_SL g259 ( 
.A(n_216),
.B(n_236),
.Y(n_259)
);

INVx2_ASAP7_75t_L g217 ( 
.A(n_205),
.Y(n_217)
);

INVxp67_ASAP7_75t_L g262 ( 
.A(n_217),
.Y(n_262)
);

CKINVDCx20_ASAP7_75t_R g218 ( 
.A(n_198),
.Y(n_218)
);

NAND2xp5_ASAP7_75t_SL g268 ( 
.A(n_218),
.B(n_221),
.Y(n_268)
);

OAI22xp5_ASAP7_75t_L g283 ( 
.A1(n_219),
.A2(n_228),
.B1(n_230),
.B2(n_238),
.Y(n_283)
);

CKINVDCx20_ASAP7_75t_R g221 ( 
.A(n_198),
.Y(n_221)
);

CKINVDCx20_ASAP7_75t_R g222 ( 
.A(n_208),
.Y(n_222)
);

NAND2xp5_ASAP7_75t_SL g274 ( 
.A(n_222),
.B(n_231),
.Y(n_274)
);

AOI21xp5_ASAP7_75t_L g223 ( 
.A1(n_195),
.A2(n_134),
.B(n_130),
.Y(n_223)
);

OAI21xp5_ASAP7_75t_SL g270 ( 
.A1(n_223),
.A2(n_225),
.B(n_226),
.Y(n_270)
);

AND2x2_ASAP7_75t_L g225 ( 
.A(n_176),
.B(n_145),
.Y(n_225)
);

OR2x2_ASAP7_75t_SL g226 ( 
.A(n_169),
.B(n_134),
.Y(n_226)
);

AOI22xp5_ASAP7_75t_L g228 ( 
.A1(n_181),
.A2(n_210),
.B1(n_182),
.B2(n_200),
.Y(n_228)
);

INVx3_ASAP7_75t_L g229 ( 
.A(n_194),
.Y(n_229)
);

NOR2xp33_ASAP7_75t_L g288 ( 
.A(n_229),
.B(n_232),
.Y(n_288)
);

CKINVDCx16_ASAP7_75t_R g231 ( 
.A(n_212),
.Y(n_231)
);

BUFx3_ASAP7_75t_L g232 ( 
.A(n_196),
.Y(n_232)
);

NOR2xp33_ASAP7_75t_L g233 ( 
.A(n_204),
.B(n_193),
.Y(n_233)
);

NAND2xp5_ASAP7_75t_SL g277 ( 
.A(n_233),
.B(n_240),
.Y(n_277)
);

AOI21xp5_ASAP7_75t_L g235 ( 
.A1(n_190),
.A2(n_184),
.B(n_215),
.Y(n_235)
);

OAI21xp5_ASAP7_75t_SL g273 ( 
.A1(n_235),
.A2(n_243),
.B(n_250),
.Y(n_273)
);

AOI22xp5_ASAP7_75t_L g238 ( 
.A1(n_170),
.A2(n_172),
.B1(n_169),
.B2(n_192),
.Y(n_238)
);

INVxp67_ASAP7_75t_L g240 ( 
.A(n_206),
.Y(n_240)
);

OAI22xp5_ASAP7_75t_SL g241 ( 
.A1(n_199),
.A2(n_175),
.B1(n_207),
.B2(n_180),
.Y(n_241)
);

OAI22xp5_ASAP7_75t_SL g258 ( 
.A1(n_241),
.A2(n_255),
.B1(n_202),
.B2(n_174),
.Y(n_258)
);

CKINVDCx20_ASAP7_75t_R g244 ( 
.A(n_208),
.Y(n_244)
);

NAND2xp5_ASAP7_75t_SL g278 ( 
.A(n_244),
.B(n_248),
.Y(n_278)
);

INVx2_ASAP7_75t_L g247 ( 
.A(n_205),
.Y(n_247)
);

CKINVDCx20_ASAP7_75t_R g263 ( 
.A(n_247),
.Y(n_263)
);

CKINVDCx20_ASAP7_75t_R g248 ( 
.A(n_213),
.Y(n_248)
);

AOI32xp33_ASAP7_75t_L g250 ( 
.A1(n_180),
.A2(n_191),
.A3(n_178),
.B1(n_173),
.B2(n_183),
.Y(n_250)
);

NOR2xp33_ASAP7_75t_L g251 ( 
.A(n_178),
.B(n_209),
.Y(n_251)
);

CKINVDCx20_ASAP7_75t_R g279 ( 
.A(n_251),
.Y(n_279)
);

AOI21xp5_ASAP7_75t_L g252 ( 
.A1(n_183),
.A2(n_185),
.B(n_171),
.Y(n_252)
);

AOI22xp33_ASAP7_75t_SL g276 ( 
.A1(n_252),
.A2(n_227),
.B1(n_245),
.B2(n_242),
.Y(n_276)
);

CKINVDCx16_ASAP7_75t_R g253 ( 
.A(n_171),
.Y(n_253)
);

BUFx24_ASAP7_75t_SL g267 ( 
.A(n_253),
.Y(n_267)
);

BUFx3_ASAP7_75t_L g254 ( 
.A(n_196),
.Y(n_254)
);

CKINVDCx20_ASAP7_75t_R g286 ( 
.A(n_254),
.Y(n_286)
);

AOI22xp5_ASAP7_75t_L g255 ( 
.A1(n_202),
.A2(n_174),
.B1(n_189),
.B2(n_177),
.Y(n_255)
);

XNOR2xp5_ASAP7_75t_L g257 ( 
.A(n_237),
.B(n_201),
.Y(n_257)
);

MAJIxp5_ASAP7_75t_L g292 ( 
.A(n_257),
.B(n_269),
.C(n_272),
.Y(n_292)
);

NOR2xp33_ASAP7_75t_L g311 ( 
.A(n_258),
.B(n_287),
.Y(n_311)
);

NAND2xp5_ASAP7_75t_SL g306 ( 
.A(n_259),
.B(n_261),
.Y(n_306)
);

NAND2xp5_ASAP7_75t_L g260 ( 
.A(n_256),
.B(n_186),
.Y(n_260)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_260),
.Y(n_298)
);

NOR2xp33_ASAP7_75t_SL g261 ( 
.A(n_234),
.B(n_186),
.Y(n_261)
);

AOI22xp5_ASAP7_75t_L g264 ( 
.A1(n_246),
.A2(n_187),
.B1(n_177),
.B2(n_197),
.Y(n_264)
);

OAI22xp5_ASAP7_75t_SL g313 ( 
.A1(n_264),
.A2(n_284),
.B1(n_289),
.B2(n_271),
.Y(n_313)
);

NAND2xp5_ASAP7_75t_L g265 ( 
.A(n_256),
.B(n_203),
.Y(n_265)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_265),
.Y(n_305)
);

NAND2xp5_ASAP7_75t_L g266 ( 
.A(n_220),
.B(n_189),
.Y(n_266)
);

NAND2xp5_ASAP7_75t_L g297 ( 
.A(n_266),
.B(n_280),
.Y(n_297)
);

MAJIxp5_ASAP7_75t_L g269 ( 
.A(n_237),
.B(n_235),
.C(n_249),
.Y(n_269)
);

AOI22xp5_ASAP7_75t_SL g271 ( 
.A1(n_225),
.A2(n_211),
.B1(n_213),
.B2(n_226),
.Y(n_271)
);

OAI21xp5_ASAP7_75t_L g295 ( 
.A1(n_271),
.A2(n_290),
.B(n_274),
.Y(n_295)
);

XOR2xp5_ASAP7_75t_L g272 ( 
.A(n_249),
.B(n_211),
.Y(n_272)
);

XOR2xp5_ASAP7_75t_L g275 ( 
.A(n_228),
.B(n_241),
.Y(n_275)
);

MAJIxp5_ASAP7_75t_L g302 ( 
.A(n_275),
.B(n_282),
.C(n_287),
.Y(n_302)
);

OAI21xp5_ASAP7_75t_SL g299 ( 
.A1(n_276),
.A2(n_270),
.B(n_285),
.Y(n_299)
);

NAND2xp5_ASAP7_75t_L g280 ( 
.A(n_220),
.B(n_238),
.Y(n_280)
);

MAJx2_ASAP7_75t_L g281 ( 
.A(n_243),
.B(n_234),
.C(n_224),
.Y(n_281)
);

XNOR2xp5_ASAP7_75t_L g291 ( 
.A(n_281),
.B(n_222),
.Y(n_291)
);

XOR2xp5_ASAP7_75t_L g282 ( 
.A(n_224),
.B(n_225),
.Y(n_282)
);

AOI22xp5_ASAP7_75t_L g284 ( 
.A1(n_223),
.A2(n_227),
.B1(n_245),
.B2(n_242),
.Y(n_284)
);

NAND2xp5_ASAP7_75t_L g285 ( 
.A(n_236),
.B(n_252),
.Y(n_285)
);

NAND2xp5_ASAP7_75t_L g300 ( 
.A(n_285),
.B(n_258),
.Y(n_300)
);

XNOR2xp5_ASAP7_75t_L g287 ( 
.A(n_255),
.B(n_219),
.Y(n_287)
);

OAI22xp5_ASAP7_75t_SL g289 ( 
.A1(n_240),
.A2(n_239),
.B1(n_218),
.B2(n_221),
.Y(n_289)
);

OAI22x1_ASAP7_75t_SL g290 ( 
.A1(n_239),
.A2(n_254),
.B1(n_232),
.B2(n_229),
.Y(n_290)
);

AOI22xp5_ASAP7_75t_L g293 ( 
.A1(n_290),
.A2(n_244),
.B1(n_248),
.B2(n_247),
.Y(n_293)
);

XNOR2xp5_ASAP7_75t_SL g322 ( 
.A(n_291),
.B(n_292),
.Y(n_322)
);

OAI21xp5_ASAP7_75t_SL g337 ( 
.A1(n_293),
.A2(n_299),
.B(n_309),
.Y(n_337)
);

OR2x2_ASAP7_75t_L g294 ( 
.A(n_284),
.B(n_217),
.Y(n_294)
);

OAI21xp5_ASAP7_75t_L g323 ( 
.A1(n_294),
.A2(n_295),
.B(n_316),
.Y(n_323)
);

BUFx2_ASAP7_75t_L g296 ( 
.A(n_262),
.Y(n_296)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_296),
.Y(n_334)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_300),
.Y(n_335)
);

NAND2xp5_ASAP7_75t_L g301 ( 
.A(n_266),
.B(n_260),
.Y(n_301)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_301),
.Y(n_321)
);

CKINVDCx16_ASAP7_75t_R g303 ( 
.A(n_268),
.Y(n_303)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_303),
.Y(n_326)
);

NAND2xp5_ASAP7_75t_L g304 ( 
.A(n_265),
.B(n_289),
.Y(n_304)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_304),
.Y(n_329)
);

NAND2xp5_ASAP7_75t_L g307 ( 
.A(n_261),
.B(n_280),
.Y(n_307)
);

INVx1_ASAP7_75t_L g338 ( 
.A(n_307),
.Y(n_338)
);

INVxp67_ASAP7_75t_L g308 ( 
.A(n_288),
.Y(n_308)
);

AOI22xp5_ASAP7_75t_SL g339 ( 
.A1(n_308),
.A2(n_310),
.B1(n_303),
.B2(n_309),
.Y(n_339)
);

CKINVDCx20_ASAP7_75t_R g309 ( 
.A(n_278),
.Y(n_309)
);

CKINVDCx16_ASAP7_75t_R g310 ( 
.A(n_259),
.Y(n_310)
);

NOR2xp33_ASAP7_75t_SL g327 ( 
.A(n_310),
.B(n_314),
.Y(n_327)
);

AOI22xp5_ASAP7_75t_L g333 ( 
.A1(n_311),
.A2(n_317),
.B1(n_316),
.B2(n_298),
.Y(n_333)
);

MAJIxp5_ASAP7_75t_L g312 ( 
.A(n_269),
.B(n_282),
.C(n_273),
.Y(n_312)
);

MAJIxp5_ASAP7_75t_L g320 ( 
.A(n_312),
.B(n_315),
.C(n_292),
.Y(n_320)
);

XNOR2xp5_ASAP7_75t_L g340 ( 
.A(n_313),
.B(n_318),
.Y(n_340)
);

NOR2xp33_ASAP7_75t_L g314 ( 
.A(n_286),
.B(n_279),
.Y(n_314)
);

MAJIxp5_ASAP7_75t_L g315 ( 
.A(n_273),
.B(n_272),
.C(n_275),
.Y(n_315)
);

AND2x2_ASAP7_75t_L g316 ( 
.A(n_264),
.B(n_283),
.Y(n_316)
);

OAI22xp33_ASAP7_75t_SL g317 ( 
.A1(n_279),
.A2(n_270),
.B1(n_286),
.B2(n_277),
.Y(n_317)
);

NOR2xp33_ASAP7_75t_L g318 ( 
.A(n_262),
.B(n_263),
.Y(n_318)
);

OAI22xp5_ASAP7_75t_SL g319 ( 
.A1(n_281),
.A2(n_257),
.B1(n_263),
.B2(n_267),
.Y(n_319)
);

OAI22xp5_ASAP7_75t_SL g330 ( 
.A1(n_319),
.A2(n_307),
.B1(n_298),
.B2(n_300),
.Y(n_330)
);

XOR2xp5_ASAP7_75t_L g349 ( 
.A(n_320),
.B(n_322),
.Y(n_349)
);

MAJIxp5_ASAP7_75t_L g324 ( 
.A(n_312),
.B(n_315),
.C(n_302),
.Y(n_324)
);

MAJIxp5_ASAP7_75t_L g358 ( 
.A(n_324),
.B(n_328),
.C(n_331),
.Y(n_358)
);

XOR2xp5_ASAP7_75t_L g325 ( 
.A(n_302),
.B(n_291),
.Y(n_325)
);

XOR2xp5_ASAP7_75t_L g354 ( 
.A(n_325),
.B(n_336),
.Y(n_354)
);

MAJIxp5_ASAP7_75t_L g328 ( 
.A(n_299),
.B(n_297),
.C(n_319),
.Y(n_328)
);

NAND2xp5_ASAP7_75t_SL g346 ( 
.A(n_330),
.B(n_296),
.Y(n_346)
);

MAJIxp5_ASAP7_75t_L g331 ( 
.A(n_297),
.B(n_305),
.C(n_301),
.Y(n_331)
);

OAI21xp5_ASAP7_75t_L g332 ( 
.A1(n_294),
.A2(n_295),
.B(n_304),
.Y(n_332)
);

AOI21xp5_ASAP7_75t_L g350 ( 
.A1(n_332),
.A2(n_323),
.B(n_337),
.Y(n_350)
);

OAI22xp5_ASAP7_75t_L g343 ( 
.A1(n_333),
.A2(n_293),
.B1(n_305),
.B2(n_308),
.Y(n_343)
);

XOR2xp5_ASAP7_75t_L g336 ( 
.A(n_313),
.B(n_316),
.Y(n_336)
);

NAND2xp5_ASAP7_75t_L g348 ( 
.A(n_339),
.B(n_296),
.Y(n_348)
);

XNOR2xp5_ASAP7_75t_SL g341 ( 
.A(n_306),
.B(n_294),
.Y(n_341)
);

XOR2xp5_ASAP7_75t_L g359 ( 
.A(n_341),
.B(n_332),
.Y(n_359)
);

INVx1_ASAP7_75t_L g342 ( 
.A(n_327),
.Y(n_342)
);

INVx1_ASAP7_75t_L g360 ( 
.A(n_342),
.Y(n_360)
);

INVxp67_ASAP7_75t_L g361 ( 
.A(n_343),
.Y(n_361)
);

HB1xp67_ASAP7_75t_L g344 ( 
.A(n_334),
.Y(n_344)
);

XNOR2xp5_ASAP7_75t_L g365 ( 
.A(n_344),
.B(n_355),
.Y(n_365)
);

INVx1_ASAP7_75t_L g345 ( 
.A(n_326),
.Y(n_345)
);

NAND2xp5_ASAP7_75t_L g363 ( 
.A(n_345),
.B(n_346),
.Y(n_363)
);

INVx1_ASAP7_75t_L g347 ( 
.A(n_335),
.Y(n_347)
);

NAND2xp5_ASAP7_75t_L g370 ( 
.A(n_347),
.B(n_352),
.Y(n_370)
);

OAI21xp5_ASAP7_75t_L g362 ( 
.A1(n_348),
.A2(n_350),
.B(n_323),
.Y(n_362)
);

AOI22xp5_ASAP7_75t_L g351 ( 
.A1(n_335),
.A2(n_329),
.B1(n_338),
.B2(n_336),
.Y(n_351)
);

OAI22xp5_ASAP7_75t_L g364 ( 
.A1(n_351),
.A2(n_333),
.B1(n_340),
.B2(n_337),
.Y(n_364)
);

INVx1_ASAP7_75t_L g352 ( 
.A(n_339),
.Y(n_352)
);

INVx1_ASAP7_75t_L g353 ( 
.A(n_334),
.Y(n_353)
);

NOR2xp33_ASAP7_75t_SL g369 ( 
.A(n_353),
.B(n_356),
.Y(n_369)
);

NAND2xp5_ASAP7_75t_L g355 ( 
.A(n_331),
.B(n_321),
.Y(n_355)
);

INVx1_ASAP7_75t_L g356 ( 
.A(n_341),
.Y(n_356)
);

HB1xp67_ASAP7_75t_L g357 ( 
.A(n_328),
.Y(n_357)
);

CKINVDCx5p33_ASAP7_75t_R g371 ( 
.A(n_357),
.Y(n_371)
);

MAJIxp5_ASAP7_75t_L g367 ( 
.A(n_359),
.B(n_320),
.C(n_324),
.Y(n_367)
);

INVx1_ASAP7_75t_L g373 ( 
.A(n_362),
.Y(n_373)
);

INVx1_ASAP7_75t_L g374 ( 
.A(n_364),
.Y(n_374)
);

BUFx24_ASAP7_75t_SL g366 ( 
.A(n_355),
.Y(n_366)
);

NOR2xp33_ASAP7_75t_SL g376 ( 
.A(n_366),
.B(n_372),
.Y(n_376)
);

NAND2xp5_ASAP7_75t_L g375 ( 
.A(n_367),
.B(n_368),
.Y(n_375)
);

MAJIxp5_ASAP7_75t_L g368 ( 
.A(n_358),
.B(n_325),
.C(n_322),
.Y(n_368)
);

MAJIxp5_ASAP7_75t_L g372 ( 
.A(n_358),
.B(n_340),
.C(n_330),
.Y(n_372)
);

AOI22xp5_ASAP7_75t_SL g377 ( 
.A1(n_361),
.A2(n_350),
.B1(n_347),
.B2(n_359),
.Y(n_377)
);

OR2x2_ASAP7_75t_L g381 ( 
.A(n_377),
.B(n_378),
.Y(n_381)
);

AOI22xp5_ASAP7_75t_SL g378 ( 
.A1(n_361),
.A2(n_348),
.B1(n_354),
.B2(n_345),
.Y(n_378)
);

NAND2xp5_ASAP7_75t_L g379 ( 
.A(n_371),
.B(n_363),
.Y(n_379)
);

INVx1_ASAP7_75t_L g380 ( 
.A(n_379),
.Y(n_380)
);

INVx1_ASAP7_75t_L g382 ( 
.A(n_379),
.Y(n_382)
);

AOI21xp5_ASAP7_75t_L g385 ( 
.A1(n_382),
.A2(n_383),
.B(n_365),
.Y(n_385)
);

OAI21xp5_ASAP7_75t_L g383 ( 
.A1(n_373),
.A2(n_372),
.B(n_360),
.Y(n_383)
);

MAJIxp5_ASAP7_75t_L g384 ( 
.A(n_380),
.B(n_375),
.C(n_376),
.Y(n_384)
);

OR2x2_ASAP7_75t_L g388 ( 
.A(n_384),
.B(n_386),
.Y(n_388)
);

AOI22xp33_ASAP7_75t_L g387 ( 
.A1(n_385),
.A2(n_381),
.B1(n_367),
.B2(n_378),
.Y(n_387)
);

MAJIxp5_ASAP7_75t_L g386 ( 
.A(n_381),
.B(n_371),
.C(n_374),
.Y(n_386)
);

MAJIxp5_ASAP7_75t_L g389 ( 
.A(n_387),
.B(n_377),
.C(n_368),
.Y(n_389)
);

INVx1_ASAP7_75t_L g390 ( 
.A(n_389),
.Y(n_390)
);

NAND2xp5_ASAP7_75t_L g391 ( 
.A(n_390),
.B(n_388),
.Y(n_391)
);

AOI311xp33_ASAP7_75t_L g392 ( 
.A1(n_391),
.A2(n_369),
.A3(n_370),
.B(n_351),
.C(n_349),
.Y(n_392)
);

NAND2xp5_ASAP7_75t_SL g393 ( 
.A(n_392),
.B(n_354),
.Y(n_393)
);

XNOR2xp5_ASAP7_75t_L g394 ( 
.A(n_393),
.B(n_349),
.Y(n_394)
);


endmodule