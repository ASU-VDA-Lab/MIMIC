module fake_jpeg_5671_n_181 (n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_181);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_181;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_14;
wire n_73;
wire n_152;
wire n_19;
wire n_84;
wire n_59;
wire n_98;
wire n_178;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_13;
wire n_175;
wire n_21;
wire n_57;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_44;
wire n_24;
wire n_143;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_121;
wire n_130;
wire n_99;
wire n_70;
wire n_177;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_161;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_176;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_36;
wire n_62;
wire n_167;
wire n_174;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_140;
wire n_82;
wire n_128;
wire n_118;
wire n_96;

INVx1_ASAP7_75t_L g13 ( 
.A(n_9),
.Y(n_13)
);

CKINVDCx20_ASAP7_75t_R g14 ( 
.A(n_3),
.Y(n_14)
);

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_4),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_6),
.Y(n_16)
);

BUFx5_ASAP7_75t_L g17 ( 
.A(n_12),
.Y(n_17)
);

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_12),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_4),
.Y(n_19)
);

BUFx16f_ASAP7_75t_L g20 ( 
.A(n_11),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_11),
.Y(n_21)
);

BUFx5_ASAP7_75t_L g22 ( 
.A(n_5),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_10),
.Y(n_23)
);

CKINVDCx16_ASAP7_75t_R g24 ( 
.A(n_11),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_6),
.Y(n_25)
);

NOR2xp33_ASAP7_75t_L g26 ( 
.A(n_13),
.B(n_0),
.Y(n_26)
);

NOR2xp33_ASAP7_75t_L g39 ( 
.A(n_26),
.B(n_28),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_20),
.Y(n_27)
);

INVx11_ASAP7_75t_L g44 ( 
.A(n_27),
.Y(n_44)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_20),
.Y(n_28)
);

INVx8_ASAP7_75t_L g29 ( 
.A(n_20),
.Y(n_29)
);

INVx8_ASAP7_75t_L g50 ( 
.A(n_29),
.Y(n_50)
);

INVx11_ASAP7_75t_L g30 ( 
.A(n_19),
.Y(n_30)
);

NOR2xp33_ASAP7_75t_L g46 ( 
.A(n_30),
.B(n_32),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_20),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_31),
.Y(n_38)
);

INVx6_ASAP7_75t_L g32 ( 
.A(n_20),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_22),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_L g47 ( 
.A(n_33),
.B(n_34),
.Y(n_47)
);

INVx2_ASAP7_75t_L g34 ( 
.A(n_17),
.Y(n_34)
);

INVx2_ASAP7_75t_L g35 ( 
.A(n_17),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_35),
.B(n_18),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_L g36 ( 
.A(n_26),
.B(n_13),
.Y(n_36)
);

NAND2xp5_ASAP7_75t_L g58 ( 
.A(n_36),
.B(n_25),
.Y(n_58)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_34),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_37),
.B(n_40),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_SL g40 ( 
.A(n_32),
.B(n_13),
.Y(n_40)
);

OAI22xp5_ASAP7_75t_L g41 ( 
.A1(n_30),
.A2(n_16),
.B1(n_15),
.B2(n_21),
.Y(n_41)
);

AOI22xp33_ASAP7_75t_L g51 ( 
.A1(n_41),
.A2(n_16),
.B1(n_14),
.B2(n_23),
.Y(n_51)
);

AOI22xp33_ASAP7_75t_SL g42 ( 
.A1(n_30),
.A2(n_17),
.B1(n_16),
.B2(n_15),
.Y(n_42)
);

INVxp67_ASAP7_75t_L g54 ( 
.A(n_42),
.Y(n_54)
);

OR2x2_ASAP7_75t_L g43 ( 
.A(n_34),
.B(n_15),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g57 ( 
.A(n_43),
.B(n_49),
.Y(n_57)
);

NOR2x1_ASAP7_75t_L g45 ( 
.A(n_35),
.B(n_22),
.Y(n_45)
);

A2O1A1Ixp33_ASAP7_75t_L g62 ( 
.A1(n_45),
.A2(n_23),
.B(n_21),
.C(n_14),
.Y(n_62)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_48),
.Y(n_61)
);

INVx3_ASAP7_75t_L g49 ( 
.A(n_35),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_51),
.B(n_53),
.Y(n_74)
);

BUFx2_ASAP7_75t_L g52 ( 
.A(n_45),
.Y(n_52)
);

INVx3_ASAP7_75t_L g79 ( 
.A(n_52),
.Y(n_79)
);

INVx2_ASAP7_75t_SL g53 ( 
.A(n_45),
.Y(n_53)
);

INVx3_ASAP7_75t_L g56 ( 
.A(n_45),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_56),
.B(n_60),
.Y(n_77)
);

AND2x2_ASAP7_75t_L g78 ( 
.A(n_58),
.B(n_43),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_36),
.B(n_25),
.Y(n_59)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_59),
.Y(n_70)
);

INVx3_ASAP7_75t_L g60 ( 
.A(n_49),
.Y(n_60)
);

NOR2x1_ASAP7_75t_R g80 ( 
.A(n_62),
.B(n_43),
.Y(n_80)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_41),
.Y(n_63)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_63),
.Y(n_72)
);

INVx4_ASAP7_75t_L g64 ( 
.A(n_38),
.Y(n_64)
);

AOI22xp33_ASAP7_75t_SL g82 ( 
.A1(n_64),
.A2(n_65),
.B1(n_66),
.B2(n_44),
.Y(n_82)
);

AOI22xp33_ASAP7_75t_L g65 ( 
.A1(n_49),
.A2(n_22),
.B1(n_25),
.B2(n_32),
.Y(n_65)
);

INVx2_ASAP7_75t_SL g66 ( 
.A(n_38),
.Y(n_66)
);

AOI22xp5_ASAP7_75t_L g67 ( 
.A1(n_63),
.A2(n_37),
.B1(n_48),
.B2(n_40),
.Y(n_67)
);

MAJIxp5_ASAP7_75t_L g85 ( 
.A(n_67),
.B(n_73),
.C(n_75),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_L g68 ( 
.A(n_57),
.B(n_39),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_SL g86 ( 
.A(n_68),
.B(n_78),
.Y(n_86)
);

INVx2_ASAP7_75t_L g69 ( 
.A(n_60),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_69),
.B(n_66),
.Y(n_84)
);

OAI21xp5_ASAP7_75t_SL g71 ( 
.A1(n_57),
.A2(n_47),
.B(n_46),
.Y(n_71)
);

AOI21xp5_ASAP7_75t_L g93 ( 
.A1(n_71),
.A2(n_76),
.B(n_62),
.Y(n_93)
);

AOI22xp5_ASAP7_75t_L g73 ( 
.A1(n_54),
.A2(n_47),
.B1(n_46),
.B2(n_50),
.Y(n_73)
);

MAJIxp5_ASAP7_75t_L g75 ( 
.A(n_61),
.B(n_28),
.C(n_39),
.Y(n_75)
);

OAI21xp5_ASAP7_75t_SL g76 ( 
.A1(n_54),
.A2(n_28),
.B(n_43),
.Y(n_76)
);

OAI21xp5_ASAP7_75t_L g94 ( 
.A1(n_80),
.A2(n_53),
.B(n_52),
.Y(n_94)
);

INVxp67_ASAP7_75t_L g81 ( 
.A(n_55),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_SL g98 ( 
.A(n_81),
.B(n_32),
.Y(n_98)
);

INVxp67_ASAP7_75t_L g91 ( 
.A(n_82),
.Y(n_91)
);

AND2x2_ASAP7_75t_L g83 ( 
.A(n_68),
.B(n_58),
.Y(n_83)
);

AOI21xp5_ASAP7_75t_L g112 ( 
.A1(n_83),
.A2(n_94),
.B(n_96),
.Y(n_112)
);

CKINVDCx20_ASAP7_75t_R g113 ( 
.A(n_84),
.Y(n_113)
);

INVx2_ASAP7_75t_L g87 ( 
.A(n_69),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_87),
.B(n_92),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_79),
.B(n_61),
.Y(n_88)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_88),
.Y(n_99)
);

MAJIxp5_ASAP7_75t_L g89 ( 
.A(n_75),
.B(n_55),
.C(n_59),
.Y(n_89)
);

MAJIxp5_ASAP7_75t_L g104 ( 
.A(n_89),
.B(n_90),
.C(n_72),
.Y(n_104)
);

MAJIxp5_ASAP7_75t_L g90 ( 
.A(n_76),
.B(n_50),
.C(n_52),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_SL g92 ( 
.A(n_70),
.B(n_78),
.Y(n_92)
);

OAI21xp5_ASAP7_75t_L g101 ( 
.A1(n_93),
.A2(n_81),
.B(n_78),
.Y(n_101)
);

CKINVDCx20_ASAP7_75t_R g95 ( 
.A(n_77),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_95),
.B(n_97),
.Y(n_105)
);

AO22x1_ASAP7_75t_L g96 ( 
.A1(n_80),
.A2(n_53),
.B1(n_56),
.B2(n_42),
.Y(n_96)
);

CKINVDCx20_ASAP7_75t_R g97 ( 
.A(n_67),
.Y(n_97)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_98),
.Y(n_103)
);

XNOR2xp5_ASAP7_75t_L g116 ( 
.A(n_101),
.B(n_93),
.Y(n_116)
);

AOI322xp5_ASAP7_75t_L g102 ( 
.A1(n_96),
.A2(n_72),
.A3(n_74),
.B1(n_73),
.B2(n_71),
.C1(n_79),
.C2(n_44),
.Y(n_102)
);

AOI322xp5_ASAP7_75t_L g124 ( 
.A1(n_102),
.A2(n_33),
.A3(n_18),
.B1(n_31),
.B2(n_27),
.C1(n_19),
.C2(n_6),
.Y(n_124)
);

MAJIxp5_ASAP7_75t_L g120 ( 
.A(n_104),
.B(n_85),
.C(n_90),
.Y(n_120)
);

OAI22xp5_ASAP7_75t_SL g106 ( 
.A1(n_97),
.A2(n_50),
.B1(n_44),
.B2(n_29),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g127 ( 
.A(n_106),
.B(n_111),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_L g107 ( 
.A(n_83),
.B(n_66),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_L g115 ( 
.A(n_107),
.B(n_108),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_L g108 ( 
.A(n_83),
.B(n_0),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_L g109 ( 
.A(n_86),
.B(n_0),
.Y(n_109)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_109),
.Y(n_118)
);

AOI22xp5_ASAP7_75t_L g110 ( 
.A1(n_85),
.A2(n_29),
.B1(n_33),
.B2(n_38),
.Y(n_110)
);

OAI22xp5_ASAP7_75t_L g122 ( 
.A1(n_110),
.A2(n_91),
.B1(n_95),
.B2(n_87),
.Y(n_122)
);

OAI22xp5_ASAP7_75t_SL g111 ( 
.A1(n_96),
.A2(n_29),
.B1(n_64),
.B2(n_38),
.Y(n_111)
);

AOI22xp5_ASAP7_75t_SL g114 ( 
.A1(n_91),
.A2(n_24),
.B1(n_18),
.B2(n_19),
.Y(n_114)
);

INVxp67_ASAP7_75t_L g126 ( 
.A(n_114),
.Y(n_126)
);

XOR2xp5_ASAP7_75t_L g133 ( 
.A(n_116),
.B(n_120),
.Y(n_133)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_105),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_L g131 ( 
.A(n_117),
.B(n_125),
.Y(n_131)
);

HB1xp67_ASAP7_75t_L g119 ( 
.A(n_113),
.Y(n_119)
);

INVxp67_ASAP7_75t_L g135 ( 
.A(n_119),
.Y(n_135)
);

XNOR2xp5_ASAP7_75t_L g121 ( 
.A(n_112),
.B(n_89),
.Y(n_121)
);

XOR2xp5_ASAP7_75t_L g138 ( 
.A(n_121),
.B(n_101),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_SL g132 ( 
.A(n_122),
.B(n_123),
.Y(n_132)
);

OAI22xp5_ASAP7_75t_L g123 ( 
.A1(n_102),
.A2(n_94),
.B1(n_24),
.B2(n_33),
.Y(n_123)
);

XNOR2xp5_ASAP7_75t_SL g130 ( 
.A(n_124),
.B(n_111),
.Y(n_130)
);

OA21x2_ASAP7_75t_L g125 ( 
.A1(n_107),
.A2(n_19),
.B(n_27),
.Y(n_125)
);

CKINVDCx20_ASAP7_75t_R g128 ( 
.A(n_113),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_L g136 ( 
.A(n_128),
.B(n_129),
.Y(n_136)
);

CKINVDCx16_ASAP7_75t_R g129 ( 
.A(n_105),
.Y(n_129)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_130),
.Y(n_149)
);

XNOR2xp5_ASAP7_75t_SL g134 ( 
.A(n_116),
.B(n_112),
.Y(n_134)
);

XNOR2xp5_ASAP7_75t_L g151 ( 
.A(n_134),
.B(n_138),
.Y(n_151)
);

OAI21xp5_ASAP7_75t_SL g137 ( 
.A1(n_120),
.A2(n_104),
.B(n_100),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_L g142 ( 
.A(n_137),
.B(n_139),
.Y(n_142)
);

NOR3xp33_ASAP7_75t_SL g139 ( 
.A(n_121),
.B(n_108),
.C(n_110),
.Y(n_139)
);

XOR2xp5_ASAP7_75t_L g140 ( 
.A(n_115),
.B(n_100),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_L g146 ( 
.A(n_140),
.B(n_141),
.Y(n_146)
);

OAI21xp5_ASAP7_75t_SL g141 ( 
.A1(n_115),
.A2(n_109),
.B(n_103),
.Y(n_141)
);

AOI22xp5_ASAP7_75t_L g143 ( 
.A1(n_132),
.A2(n_127),
.B1(n_126),
.B2(n_106),
.Y(n_143)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_143),
.Y(n_153)
);

OAI21x1_ASAP7_75t_L g144 ( 
.A1(n_139),
.A2(n_125),
.B(n_126),
.Y(n_144)
);

OAI21xp5_ASAP7_75t_L g152 ( 
.A1(n_144),
.A2(n_114),
.B(n_118),
.Y(n_152)
);

OAI22xp5_ASAP7_75t_L g145 ( 
.A1(n_136),
.A2(n_131),
.B1(n_135),
.B2(n_134),
.Y(n_145)
);

AOI22xp5_ASAP7_75t_L g156 ( 
.A1(n_145),
.A2(n_147),
.B1(n_146),
.B2(n_149),
.Y(n_156)
);

OAI22xp5_ASAP7_75t_SL g147 ( 
.A1(n_133),
.A2(n_125),
.B1(n_103),
.B2(n_118),
.Y(n_147)
);

BUFx6f_ASAP7_75t_L g148 ( 
.A(n_135),
.Y(n_148)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_148),
.Y(n_157)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_130),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_L g154 ( 
.A(n_150),
.B(n_99),
.Y(n_154)
);

FAx1_ASAP7_75t_SL g165 ( 
.A(n_152),
.B(n_156),
.CI(n_155),
.CON(n_165),
.SN(n_165)
);

MAJIxp5_ASAP7_75t_L g161 ( 
.A(n_154),
.B(n_155),
.C(n_18),
.Y(n_161)
);

MAJIxp5_ASAP7_75t_L g155 ( 
.A(n_142),
.B(n_99),
.C(n_31),
.Y(n_155)
);

AOI21xp5_ASAP7_75t_L g158 ( 
.A1(n_147),
.A2(n_148),
.B(n_143),
.Y(n_158)
);

OAI21xp5_ASAP7_75t_SL g162 ( 
.A1(n_158),
.A2(n_160),
.B(n_1),
.Y(n_162)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_151),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_SL g164 ( 
.A(n_159),
.B(n_1),
.Y(n_164)
);

OAI21xp5_ASAP7_75t_L g160 ( 
.A1(n_151),
.A2(n_1),
.B(n_2),
.Y(n_160)
);

MAJIxp5_ASAP7_75t_L g168 ( 
.A(n_161),
.B(n_162),
.C(n_163),
.Y(n_168)
);

NAND4xp25_ASAP7_75t_SL g163 ( 
.A(n_157),
.B(n_31),
.C(n_27),
.D(n_3),
.Y(n_163)
);

OAI21xp5_ASAP7_75t_L g171 ( 
.A1(n_164),
.A2(n_166),
.B(n_5),
.Y(n_171)
);

MAJx2_ASAP7_75t_L g170 ( 
.A(n_165),
.B(n_4),
.C(n_5),
.Y(n_170)
);

INVxp67_ASAP7_75t_L g166 ( 
.A(n_160),
.Y(n_166)
);

MAJIxp5_ASAP7_75t_L g167 ( 
.A(n_153),
.B(n_2),
.C(n_3),
.Y(n_167)
);

AND2x2_ASAP7_75t_L g169 ( 
.A(n_167),
.B(n_2),
.Y(n_169)
);

NOR2xp33_ASAP7_75t_SL g175 ( 
.A(n_169),
.B(n_7),
.Y(n_175)
);

OAI22xp5_ASAP7_75t_L g173 ( 
.A1(n_170),
.A2(n_165),
.B1(n_8),
.B2(n_9),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_L g174 ( 
.A(n_171),
.B(n_7),
.Y(n_174)
);

OAI22xp5_ASAP7_75t_SL g172 ( 
.A1(n_166),
.A2(n_7),
.B1(n_8),
.B2(n_9),
.Y(n_172)
);

NOR2xp33_ASAP7_75t_L g176 ( 
.A(n_172),
.B(n_8),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_SL g177 ( 
.A(n_173),
.B(n_175),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_L g178 ( 
.A(n_174),
.B(n_176),
.Y(n_178)
);

OAI21xp5_ASAP7_75t_SL g179 ( 
.A1(n_177),
.A2(n_168),
.B(n_172),
.Y(n_179)
);

MAJIxp5_ASAP7_75t_L g180 ( 
.A(n_179),
.B(n_178),
.C(n_10),
.Y(n_180)
);

XOR2xp5_ASAP7_75t_L g181 ( 
.A(n_180),
.B(n_10),
.Y(n_181)
);


endmodule