module fake_jpeg_27930_n_313 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_313);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_313;

wire n_253;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_51;
wire n_84;
wire n_59;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_20;
wire n_18;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_208;
wire n_308;
wire n_297;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_1),
.Y(n_16)
);

NOR2xp33_ASAP7_75t_L g17 ( 
.A(n_7),
.B(n_13),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_8),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_12),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_14),
.Y(n_20)
);

CKINVDCx16_ASAP7_75t_R g21 ( 
.A(n_15),
.Y(n_21)
);

INVxp67_ASAP7_75t_L g22 ( 
.A(n_5),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_2),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_10),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_13),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_9),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_1),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_15),
.Y(n_28)
);

BUFx8_ASAP7_75t_L g29 ( 
.A(n_8),
.Y(n_29)
);

INVx6_ASAP7_75t_SL g30 ( 
.A(n_4),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_12),
.Y(n_31)
);

INVx4_ASAP7_75t_L g32 ( 
.A(n_4),
.Y(n_32)
);

BUFx5_ASAP7_75t_L g33 ( 
.A(n_4),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_7),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_9),
.Y(n_35)
);

INVx4_ASAP7_75t_L g36 ( 
.A(n_19),
.Y(n_36)
);

INVx2_ASAP7_75t_L g46 ( 
.A(n_36),
.Y(n_46)
);

INVx2_ASAP7_75t_L g37 ( 
.A(n_32),
.Y(n_37)
);

BUFx24_ASAP7_75t_L g59 ( 
.A(n_37),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_32),
.Y(n_38)
);

INVx6_ASAP7_75t_L g55 ( 
.A(n_38),
.Y(n_55)
);

INVx3_ASAP7_75t_L g39 ( 
.A(n_19),
.Y(n_39)
);

INVx6_ASAP7_75t_L g66 ( 
.A(n_39),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g40 ( 
.A(n_17),
.B(n_8),
.Y(n_40)
);

AND2x2_ASAP7_75t_L g69 ( 
.A(n_40),
.B(n_45),
.Y(n_69)
);

INVx3_ASAP7_75t_L g41 ( 
.A(n_19),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_41),
.Y(n_63)
);

HB1xp67_ASAP7_75t_L g42 ( 
.A(n_29),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_42),
.Y(n_51)
);

INVx2_ASAP7_75t_L g43 ( 
.A(n_32),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_43),
.Y(n_67)
);

INVx3_ASAP7_75t_L g44 ( 
.A(n_19),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g47 ( 
.A(n_44),
.B(n_35),
.Y(n_47)
);

NAND2xp5_ASAP7_75t_SL g45 ( 
.A(n_17),
.B(n_0),
.Y(n_45)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_47),
.Y(n_79)
);

BUFx12f_ASAP7_75t_L g48 ( 
.A(n_38),
.Y(n_48)
);

BUFx3_ASAP7_75t_L g99 ( 
.A(n_48),
.Y(n_99)
);

OAI22xp33_ASAP7_75t_L g49 ( 
.A1(n_44),
.A2(n_35),
.B1(n_20),
.B2(n_26),
.Y(n_49)
);

OAI22xp5_ASAP7_75t_L g77 ( 
.A1(n_49),
.A2(n_54),
.B1(n_30),
.B2(n_21),
.Y(n_77)
);

INVx2_ASAP7_75t_SL g50 ( 
.A(n_38),
.Y(n_50)
);

INVx1_ASAP7_75t_SL g78 ( 
.A(n_50),
.Y(n_78)
);

OAI22xp5_ASAP7_75t_L g52 ( 
.A1(n_45),
.A2(n_34),
.B1(n_31),
.B2(n_18),
.Y(n_52)
);

AOI22xp5_ASAP7_75t_L g101 ( 
.A1(n_52),
.A2(n_26),
.B1(n_29),
.B2(n_10),
.Y(n_101)
);

AOI22xp33_ASAP7_75t_SL g53 ( 
.A1(n_36),
.A2(n_18),
.B1(n_28),
.B2(n_31),
.Y(n_53)
);

AOI22xp33_ASAP7_75t_SL g70 ( 
.A1(n_53),
.A2(n_24),
.B1(n_25),
.B2(n_28),
.Y(n_70)
);

AOI22xp5_ASAP7_75t_L g54 ( 
.A1(n_39),
.A2(n_30),
.B1(n_22),
.B2(n_23),
.Y(n_54)
);

BUFx12_ASAP7_75t_L g56 ( 
.A(n_42),
.Y(n_56)
);

INVx4_ASAP7_75t_L g94 ( 
.A(n_56),
.Y(n_94)
);

INVx8_ASAP7_75t_L g57 ( 
.A(n_36),
.Y(n_57)
);

INVx3_ASAP7_75t_L g97 ( 
.A(n_57),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_SL g58 ( 
.A(n_40),
.B(n_34),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_SL g73 ( 
.A(n_58),
.B(n_28),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_37),
.B(n_18),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_60),
.B(n_61),
.Y(n_72)
);

INVx3_ASAP7_75t_L g61 ( 
.A(n_43),
.Y(n_61)
);

INVx5_ASAP7_75t_L g62 ( 
.A(n_39),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_62),
.B(n_64),
.Y(n_82)
);

INVx3_ASAP7_75t_L g64 ( 
.A(n_41),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_L g65 ( 
.A(n_41),
.B(n_23),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_L g83 ( 
.A(n_65),
.B(n_68),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g68 ( 
.A(n_45),
.B(n_23),
.Y(n_68)
);

CKINVDCx16_ASAP7_75t_R g121 ( 
.A(n_70),
.Y(n_121)
);

INVx2_ASAP7_75t_L g71 ( 
.A(n_67),
.Y(n_71)
);

INVx2_ASAP7_75t_L g139 ( 
.A(n_71),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_SL g134 ( 
.A(n_73),
.B(n_75),
.Y(n_134)
);

AND2x2_ASAP7_75t_SL g74 ( 
.A(n_51),
.B(n_35),
.Y(n_74)
);

MAJIxp5_ASAP7_75t_L g113 ( 
.A(n_74),
.B(n_86),
.C(n_95),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_SL g75 ( 
.A(n_69),
.B(n_16),
.Y(n_75)
);

INVxp67_ASAP7_75t_L g76 ( 
.A(n_54),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g112 ( 
.A(n_76),
.B(n_80),
.Y(n_112)
);

AOI22xp5_ASAP7_75t_L g116 ( 
.A1(n_77),
.A2(n_88),
.B1(n_33),
.B2(n_1),
.Y(n_116)
);

CKINVDCx20_ASAP7_75t_R g80 ( 
.A(n_65),
.Y(n_80)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_57),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g123 ( 
.A(n_81),
.B(n_89),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_L g84 ( 
.A(n_68),
.B(n_27),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g119 ( 
.A(n_84),
.B(n_87),
.Y(n_119)
);

AOI22xp33_ASAP7_75t_SL g85 ( 
.A1(n_62),
.A2(n_16),
.B1(n_27),
.B2(n_25),
.Y(n_85)
);

OAI22xp33_ASAP7_75t_SL g135 ( 
.A1(n_85),
.A2(n_90),
.B1(n_103),
.B2(n_0),
.Y(n_135)
);

MAJIxp5_ASAP7_75t_L g86 ( 
.A(n_69),
.B(n_35),
.C(n_20),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_L g87 ( 
.A(n_69),
.B(n_20),
.Y(n_87)
);

OAI22xp5_ASAP7_75t_L g88 ( 
.A1(n_55),
.A2(n_30),
.B1(n_25),
.B2(n_24),
.Y(n_88)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_61),
.Y(n_89)
);

AOI22xp33_ASAP7_75t_SL g90 ( 
.A1(n_55),
.A2(n_24),
.B1(n_29),
.B2(n_26),
.Y(n_90)
);

INVx2_ASAP7_75t_L g91 ( 
.A(n_67),
.Y(n_91)
);

BUFx2_ASAP7_75t_SL g137 ( 
.A(n_91),
.Y(n_137)
);

XNOR2xp5_ASAP7_75t_SL g92 ( 
.A(n_51),
.B(n_29),
.Y(n_92)
);

XOR2xp5_ASAP7_75t_L g136 ( 
.A(n_92),
.B(n_3),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_L g93 ( 
.A(n_46),
.B(n_20),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_L g120 ( 
.A(n_93),
.B(n_104),
.Y(n_120)
);

AND2x2_ASAP7_75t_L g95 ( 
.A(n_49),
.B(n_26),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_59),
.B(n_21),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_96),
.B(n_98),
.Y(n_117)
);

INVxp67_ASAP7_75t_L g98 ( 
.A(n_56),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_SL g100 ( 
.A(n_59),
.B(n_10),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_SL g118 ( 
.A(n_100),
.B(n_101),
.Y(n_118)
);

OA22x2_ASAP7_75t_SL g102 ( 
.A1(n_66),
.A2(n_29),
.B1(n_33),
.B2(n_2),
.Y(n_102)
);

AND2x2_ASAP7_75t_L g114 ( 
.A(n_102),
.B(n_106),
.Y(n_114)
);

AOI22xp33_ASAP7_75t_SL g103 ( 
.A1(n_66),
.A2(n_7),
.B1(n_15),
.B2(n_14),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_L g104 ( 
.A(n_46),
.B(n_0),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_59),
.B(n_14),
.Y(n_105)
);

CKINVDCx20_ASAP7_75t_R g138 ( 
.A(n_105),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_SL g106 ( 
.A(n_56),
.B(n_11),
.Y(n_106)
);

INVx2_ASAP7_75t_L g107 ( 
.A(n_48),
.Y(n_107)
);

INVx1_ASAP7_75t_SL g127 ( 
.A(n_107),
.Y(n_127)
);

AOI22xp33_ASAP7_75t_L g108 ( 
.A1(n_64),
.A2(n_33),
.B1(n_13),
.B2(n_12),
.Y(n_108)
);

AOI22xp33_ASAP7_75t_L g122 ( 
.A1(n_108),
.A2(n_11),
.B1(n_9),
.B2(n_2),
.Y(n_122)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_59),
.Y(n_109)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_109),
.Y(n_115)
);

OAI22xp33_ASAP7_75t_L g110 ( 
.A1(n_76),
.A2(n_50),
.B1(n_63),
.B2(n_48),
.Y(n_110)
);

AOI22xp33_ASAP7_75t_L g157 ( 
.A1(n_110),
.A2(n_116),
.B1(n_122),
.B2(n_135),
.Y(n_157)
);

O2A1O1Ixp33_ASAP7_75t_L g111 ( 
.A1(n_102),
.A2(n_50),
.B(n_63),
.C(n_48),
.Y(n_111)
);

OA21x2_ASAP7_75t_L g158 ( 
.A1(n_111),
.A2(n_109),
.B(n_88),
.Y(n_158)
);

AOI22xp5_ASAP7_75t_L g124 ( 
.A1(n_95),
.A2(n_11),
.B1(n_1),
.B2(n_2),
.Y(n_124)
);

OAI22xp5_ASAP7_75t_SL g143 ( 
.A1(n_124),
.A2(n_84),
.B1(n_101),
.B2(n_83),
.Y(n_143)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_93),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_L g149 ( 
.A(n_125),
.B(n_128),
.Y(n_149)
);

AND2x2_ASAP7_75t_L g126 ( 
.A(n_80),
.B(n_6),
.Y(n_126)
);

AOI21xp5_ASAP7_75t_L g142 ( 
.A1(n_126),
.A2(n_131),
.B(n_100),
.Y(n_142)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_82),
.Y(n_128)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_72),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_L g160 ( 
.A(n_129),
.B(n_130),
.Y(n_160)
);

INVx1_ASAP7_75t_SL g130 ( 
.A(n_99),
.Y(n_130)
);

NAND2xp33_ASAP7_75t_SL g131 ( 
.A(n_92),
.B(n_0),
.Y(n_131)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_104),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_L g169 ( 
.A(n_132),
.B(n_133),
.Y(n_169)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_102),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_L g146 ( 
.A(n_136),
.B(n_86),
.Y(n_146)
);

AOI22xp5_ASAP7_75t_L g140 ( 
.A1(n_133),
.A2(n_95),
.B1(n_77),
.B2(n_74),
.Y(n_140)
);

OAI22xp5_ASAP7_75t_SL g184 ( 
.A1(n_140),
.A2(n_141),
.B1(n_162),
.B2(n_163),
.Y(n_184)
);

AOI22xp5_ASAP7_75t_L g141 ( 
.A1(n_121),
.A2(n_74),
.B1(n_79),
.B2(n_83),
.Y(n_141)
);

OAI21xp5_ASAP7_75t_SL g189 ( 
.A1(n_142),
.A2(n_144),
.B(n_155),
.Y(n_189)
);

AOI22xp5_ASAP7_75t_L g187 ( 
.A1(n_143),
.A2(n_150),
.B1(n_167),
.B2(n_126),
.Y(n_187)
);

AOI21xp5_ASAP7_75t_L g144 ( 
.A1(n_121),
.A2(n_81),
.B(n_102),
.Y(n_144)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_123),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_L g172 ( 
.A(n_145),
.B(n_147),
.Y(n_172)
);

XOR2xp5_ASAP7_75t_L g177 ( 
.A(n_146),
.B(n_136),
.Y(n_177)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_123),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_L g148 ( 
.A(n_120),
.B(n_87),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_L g197 ( 
.A(n_148),
.B(n_153),
.Y(n_197)
);

OAI22xp5_ASAP7_75t_SL g150 ( 
.A1(n_125),
.A2(n_79),
.B1(n_89),
.B2(n_91),
.Y(n_150)
);

CKINVDCx16_ASAP7_75t_R g151 ( 
.A(n_112),
.Y(n_151)
);

NOR2xp33_ASAP7_75t_L g179 ( 
.A(n_151),
.B(n_152),
.Y(n_179)
);

INVxp67_ASAP7_75t_L g152 ( 
.A(n_117),
.Y(n_152)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_137),
.Y(n_153)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_112),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_L g201 ( 
.A(n_154),
.B(n_161),
.Y(n_201)
);

CKINVDCx14_ASAP7_75t_R g155 ( 
.A(n_114),
.Y(n_155)
);

INVxp67_ASAP7_75t_L g156 ( 
.A(n_114),
.Y(n_156)
);

NOR2xp33_ASAP7_75t_L g186 ( 
.A(n_156),
.B(n_166),
.Y(n_186)
);

OA22x2_ASAP7_75t_L g183 ( 
.A1(n_158),
.A2(n_163),
.B1(n_144),
.B2(n_151),
.Y(n_183)
);

INVx4_ASAP7_75t_L g159 ( 
.A(n_127),
.Y(n_159)
);

INVx2_ASAP7_75t_L g190 ( 
.A(n_159),
.Y(n_190)
);

NOR2xp33_ASAP7_75t_SL g161 ( 
.A(n_119),
.B(n_73),
.Y(n_161)
);

AOI22xp5_ASAP7_75t_L g162 ( 
.A1(n_114),
.A2(n_71),
.B1(n_97),
.B2(n_78),
.Y(n_162)
);

AOI22xp5_ASAP7_75t_L g163 ( 
.A1(n_111),
.A2(n_97),
.B1(n_78),
.B2(n_107),
.Y(n_163)
);

AOI22xp5_ASAP7_75t_L g164 ( 
.A1(n_118),
.A2(n_98),
.B1(n_94),
.B2(n_99),
.Y(n_164)
);

OAI22xp5_ASAP7_75t_L g175 ( 
.A1(n_164),
.A2(n_118),
.B1(n_113),
.B2(n_124),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_L g165 ( 
.A(n_120),
.B(n_94),
.Y(n_165)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_165),
.Y(n_180)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_115),
.Y(n_166)
);

OAI22xp5_ASAP7_75t_SL g167 ( 
.A1(n_116),
.A2(n_3),
.B1(n_4),
.B2(n_5),
.Y(n_167)
);

NOR2xp33_ASAP7_75t_SL g168 ( 
.A(n_119),
.B(n_3),
.Y(n_168)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_168),
.Y(n_176)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_115),
.Y(n_170)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_170),
.Y(n_181)
);

CKINVDCx20_ASAP7_75t_R g171 ( 
.A(n_138),
.Y(n_171)
);

CKINVDCx20_ASAP7_75t_R g174 ( 
.A(n_171),
.Y(n_174)
);

INVxp67_ASAP7_75t_L g173 ( 
.A(n_160),
.Y(n_173)
);

NOR2xp33_ASAP7_75t_L g205 ( 
.A(n_173),
.B(n_178),
.Y(n_205)
);

AOI22xp5_ASAP7_75t_L g221 ( 
.A1(n_175),
.A2(n_199),
.B1(n_161),
.B2(n_126),
.Y(n_221)
);

XNOR2xp5_ASAP7_75t_L g219 ( 
.A(n_177),
.B(n_187),
.Y(n_219)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_160),
.Y(n_178)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_149),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_SL g211 ( 
.A(n_182),
.B(n_185),
.Y(n_211)
);

CKINVDCx14_ASAP7_75t_R g203 ( 
.A(n_183),
.Y(n_203)
);

NAND3xp33_ASAP7_75t_L g185 ( 
.A(n_171),
.B(n_134),
.C(n_131),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_L g216 ( 
.A(n_187),
.B(n_188),
.Y(n_216)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_165),
.Y(n_188)
);

INVx2_ASAP7_75t_SL g191 ( 
.A(n_159),
.Y(n_191)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_191),
.Y(n_212)
);

CKINVDCx12_ASAP7_75t_R g192 ( 
.A(n_149),
.Y(n_192)
);

INVxp67_ASAP7_75t_L g215 ( 
.A(n_192),
.Y(n_215)
);

INVxp67_ASAP7_75t_L g193 ( 
.A(n_164),
.Y(n_193)
);

OAI21xp5_ASAP7_75t_SL g207 ( 
.A1(n_193),
.A2(n_154),
.B(n_153),
.Y(n_207)
);

INVx4_ASAP7_75t_L g194 ( 
.A(n_159),
.Y(n_194)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_194),
.Y(n_222)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_150),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_L g217 ( 
.A(n_195),
.B(n_196),
.Y(n_217)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_169),
.Y(n_196)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_169),
.Y(n_198)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_198),
.Y(n_223)
);

OAI22xp5_ASAP7_75t_L g199 ( 
.A1(n_157),
.A2(n_129),
.B1(n_113),
.B2(n_128),
.Y(n_199)
);

CKINVDCx20_ASAP7_75t_R g200 ( 
.A(n_166),
.Y(n_200)
);

CKINVDCx20_ASAP7_75t_R g206 ( 
.A(n_200),
.Y(n_206)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_162),
.Y(n_202)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_202),
.Y(n_228)
);

MAJIxp5_ASAP7_75t_L g204 ( 
.A(n_177),
.B(n_146),
.C(n_155),
.Y(n_204)
);

MAJIxp5_ASAP7_75t_L g235 ( 
.A(n_204),
.B(n_197),
.C(n_186),
.Y(n_235)
);

CKINVDCx14_ASAP7_75t_R g236 ( 
.A(n_207),
.Y(n_236)
);

OAI22xp5_ASAP7_75t_SL g208 ( 
.A1(n_202),
.A2(n_140),
.B1(n_158),
.B2(n_141),
.Y(n_208)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_208),
.Y(n_234)
);

CKINVDCx20_ASAP7_75t_R g209 ( 
.A(n_174),
.Y(n_209)
);

CKINVDCx20_ASAP7_75t_R g239 ( 
.A(n_209),
.Y(n_239)
);

OAI21xp5_ASAP7_75t_L g210 ( 
.A1(n_189),
.A2(n_158),
.B(n_142),
.Y(n_210)
);

CKINVDCx14_ASAP7_75t_R g248 ( 
.A(n_210),
.Y(n_248)
);

BUFx24_ASAP7_75t_SL g213 ( 
.A(n_201),
.Y(n_213)
);

NOR2xp33_ASAP7_75t_L g232 ( 
.A(n_213),
.B(n_224),
.Y(n_232)
);

OAI22xp5_ASAP7_75t_SL g214 ( 
.A1(n_180),
.A2(n_158),
.B1(n_170),
.B2(n_148),
.Y(n_214)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_214),
.Y(n_237)
);

OAI21xp5_ASAP7_75t_SL g218 ( 
.A1(n_189),
.A2(n_147),
.B(n_145),
.Y(n_218)
);

INVxp67_ASAP7_75t_L g247 ( 
.A(n_218),
.Y(n_247)
);

XOR2xp5_ASAP7_75t_L g240 ( 
.A(n_219),
.B(n_184),
.Y(n_240)
);

OAI22xp5_ASAP7_75t_L g220 ( 
.A1(n_180),
.A2(n_167),
.B1(n_132),
.B2(n_143),
.Y(n_220)
);

OAI22xp5_ASAP7_75t_L g231 ( 
.A1(n_220),
.A2(n_227),
.B1(n_198),
.B2(n_193),
.Y(n_231)
);

XNOR2xp5_ASAP7_75t_L g249 ( 
.A(n_221),
.B(n_176),
.Y(n_249)
);

AOI21xp5_ASAP7_75t_L g224 ( 
.A1(n_183),
.A2(n_127),
.B(n_130),
.Y(n_224)
);

CKINVDCx14_ASAP7_75t_R g225 ( 
.A(n_172),
.Y(n_225)
);

NOR2xp33_ASAP7_75t_L g233 ( 
.A(n_225),
.B(n_226),
.Y(n_233)
);

CKINVDCx16_ASAP7_75t_R g226 ( 
.A(n_172),
.Y(n_226)
);

AOI22xp5_ASAP7_75t_L g227 ( 
.A1(n_184),
.A2(n_168),
.B1(n_138),
.B2(n_139),
.Y(n_227)
);

NAND2xp5_ASAP7_75t_L g229 ( 
.A(n_226),
.B(n_201),
.Y(n_229)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_229),
.Y(n_255)
);

AND2x6_ASAP7_75t_L g230 ( 
.A(n_218),
.B(n_183),
.Y(n_230)
);

NOR2xp33_ASAP7_75t_L g264 ( 
.A(n_230),
.B(n_245),
.Y(n_264)
);

AOI22xp5_ASAP7_75t_L g253 ( 
.A1(n_231),
.A2(n_208),
.B1(n_203),
.B2(n_220),
.Y(n_253)
);

XOR2xp5_ASAP7_75t_L g250 ( 
.A(n_235),
.B(n_240),
.Y(n_250)
);

MAJIxp5_ASAP7_75t_L g238 ( 
.A(n_219),
.B(n_188),
.C(n_197),
.Y(n_238)
);

MAJIxp5_ASAP7_75t_L g252 ( 
.A(n_238),
.B(n_244),
.C(n_246),
.Y(n_252)
);

NAND2xp5_ASAP7_75t_L g241 ( 
.A(n_223),
.B(n_205),
.Y(n_241)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_241),
.Y(n_257)
);

NAND2xp5_ASAP7_75t_L g242 ( 
.A(n_223),
.B(n_173),
.Y(n_242)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_242),
.Y(n_258)
);

NAND2xp5_ASAP7_75t_L g243 ( 
.A(n_217),
.B(n_214),
.Y(n_243)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_243),
.Y(n_261)
);

MAJIxp5_ASAP7_75t_L g244 ( 
.A(n_204),
.B(n_179),
.C(n_181),
.Y(n_244)
);

NOR2xp33_ASAP7_75t_SL g245 ( 
.A(n_211),
.B(n_134),
.Y(n_245)
);

MAJIxp5_ASAP7_75t_L g246 ( 
.A(n_221),
.B(n_181),
.C(n_183),
.Y(n_246)
);

XNOR2xp5_ASAP7_75t_L g251 ( 
.A(n_249),
.B(n_240),
.Y(n_251)
);

XNOR2xp5_ASAP7_75t_L g276 ( 
.A(n_251),
.B(n_227),
.Y(n_276)
);

CKINVDCx16_ASAP7_75t_R g267 ( 
.A(n_253),
.Y(n_267)
);

MAJIxp5_ASAP7_75t_L g254 ( 
.A(n_244),
.B(n_216),
.C(n_207),
.Y(n_254)
);

MAJIxp5_ASAP7_75t_L g269 ( 
.A(n_254),
.B(n_256),
.C(n_260),
.Y(n_269)
);

MAJIxp5_ASAP7_75t_L g256 ( 
.A(n_235),
.B(n_216),
.C(n_210),
.Y(n_256)
);

NAND2xp5_ASAP7_75t_L g259 ( 
.A(n_233),
.B(n_229),
.Y(n_259)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_259),
.Y(n_272)
);

MAJIxp5_ASAP7_75t_L g260 ( 
.A(n_238),
.B(n_224),
.C(n_217),
.Y(n_260)
);

NAND2xp5_ASAP7_75t_L g262 ( 
.A(n_242),
.B(n_206),
.Y(n_262)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_262),
.Y(n_279)
);

AOI21xp5_ASAP7_75t_L g263 ( 
.A1(n_247),
.A2(n_228),
.B(n_209),
.Y(n_263)
);

INVxp67_ASAP7_75t_L g277 ( 
.A(n_263),
.Y(n_277)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_241),
.Y(n_265)
);

NAND2xp5_ASAP7_75t_L g280 ( 
.A(n_265),
.B(n_266),
.Y(n_280)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_243),
.Y(n_266)
);

XOR2xp5_ASAP7_75t_L g268 ( 
.A(n_250),
.B(n_246),
.Y(n_268)
);

XOR2xp5_ASAP7_75t_L g281 ( 
.A(n_268),
.B(n_273),
.Y(n_281)
);

MAJIxp5_ASAP7_75t_L g270 ( 
.A(n_252),
.B(n_250),
.C(n_254),
.Y(n_270)
);

MAJIxp5_ASAP7_75t_L g286 ( 
.A(n_270),
.B(n_276),
.C(n_256),
.Y(n_286)
);

XNOR2xp5_ASAP7_75t_L g271 ( 
.A(n_251),
.B(n_249),
.Y(n_271)
);

NAND2xp5_ASAP7_75t_SL g284 ( 
.A(n_271),
.B(n_274),
.Y(n_284)
);

XOR2xp5_ASAP7_75t_L g273 ( 
.A(n_252),
.B(n_230),
.Y(n_273)
);

AOI21xp5_ASAP7_75t_L g274 ( 
.A1(n_264),
.A2(n_247),
.B(n_211),
.Y(n_274)
);

NOR2xp33_ASAP7_75t_L g275 ( 
.A(n_263),
.B(n_239),
.Y(n_275)
);

CKINVDCx20_ASAP7_75t_R g290 ( 
.A(n_275),
.Y(n_290)
);

AOI22xp5_ASAP7_75t_L g278 ( 
.A1(n_257),
.A2(n_234),
.B1(n_236),
.B2(n_237),
.Y(n_278)
);

OAI22xp5_ASAP7_75t_L g285 ( 
.A1(n_278),
.A2(n_253),
.B1(n_237),
.B2(n_234),
.Y(n_285)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_280),
.Y(n_282)
);

NAND2xp5_ASAP7_75t_L g299 ( 
.A(n_282),
.B(n_283),
.Y(n_299)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_279),
.Y(n_283)
);

XNOR2xp5_ASAP7_75t_L g292 ( 
.A(n_285),
.B(n_291),
.Y(n_292)
);

MAJx2_ASAP7_75t_L g297 ( 
.A(n_286),
.B(n_215),
.C(n_222),
.Y(n_297)
);

MAJIxp5_ASAP7_75t_L g287 ( 
.A(n_270),
.B(n_260),
.C(n_262),
.Y(n_287)
);

MAJIxp5_ASAP7_75t_L g296 ( 
.A(n_287),
.B(n_269),
.C(n_222),
.Y(n_296)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_273),
.Y(n_288)
);

AOI21xp5_ASAP7_75t_L g295 ( 
.A1(n_288),
.A2(n_268),
.B(n_269),
.Y(n_295)
);

AOI21xp5_ASAP7_75t_L g289 ( 
.A1(n_277),
.A2(n_248),
.B(n_258),
.Y(n_289)
);

OAI21xp5_ASAP7_75t_SL g294 ( 
.A1(n_289),
.A2(n_277),
.B(n_272),
.Y(n_294)
);

AOI322xp5_ASAP7_75t_L g291 ( 
.A1(n_267),
.A2(n_232),
.A3(n_206),
.B1(n_259),
.B2(n_228),
.C1(n_255),
.C2(n_261),
.Y(n_291)
);

XNOR2xp5_ASAP7_75t_L g293 ( 
.A(n_286),
.B(n_276),
.Y(n_293)
);

NOR2xp33_ASAP7_75t_L g302 ( 
.A(n_293),
.B(n_295),
.Y(n_302)
);

AOI322xp5_ASAP7_75t_L g301 ( 
.A1(n_294),
.A2(n_290),
.A3(n_284),
.B1(n_289),
.B2(n_288),
.C1(n_283),
.C2(n_281),
.Y(n_301)
);

MAJIxp5_ASAP7_75t_L g303 ( 
.A(n_296),
.B(n_297),
.C(n_298),
.Y(n_303)
);

MAJIxp5_ASAP7_75t_L g298 ( 
.A(n_287),
.B(n_212),
.C(n_194),
.Y(n_298)
);

NOR2xp33_ASAP7_75t_SL g300 ( 
.A(n_296),
.B(n_282),
.Y(n_300)
);

OAI21xp5_ASAP7_75t_SL g307 ( 
.A1(n_300),
.A2(n_304),
.B(n_191),
.Y(n_307)
);

OAI22xp5_ASAP7_75t_L g305 ( 
.A1(n_301),
.A2(n_298),
.B1(n_299),
.B2(n_297),
.Y(n_305)
);

NOR2xp33_ASAP7_75t_L g304 ( 
.A(n_292),
.B(n_190),
.Y(n_304)
);

NOR2xp33_ASAP7_75t_SL g308 ( 
.A(n_305),
.B(n_306),
.Y(n_308)
);

OAI22xp5_ASAP7_75t_L g306 ( 
.A1(n_303),
.A2(n_281),
.B1(n_212),
.B2(n_191),
.Y(n_306)
);

NOR2xp67_ASAP7_75t_SL g309 ( 
.A(n_307),
.B(n_303),
.Y(n_309)
);

MAJIxp5_ASAP7_75t_L g310 ( 
.A(n_309),
.B(n_302),
.C(n_190),
.Y(n_310)
);

OAI321xp33_ASAP7_75t_L g311 ( 
.A1(n_310),
.A2(n_308),
.A3(n_139),
.B1(n_6),
.B2(n_5),
.C(n_3),
.Y(n_311)
);

NAND2xp5_ASAP7_75t_L g312 ( 
.A(n_311),
.B(n_5),
.Y(n_312)
);

XNOR2xp5_ASAP7_75t_L g313 ( 
.A(n_312),
.B(n_6),
.Y(n_313)
);


endmodule