module fake_jpeg_31327_n_545 (n_13, n_1, n_10, n_6, n_14, n_18, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_545);

input n_13;
input n_1;
input n_10;
input n_6;
input n_14;
input n_18;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_545;

wire n_529;
wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_525;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_519;
wire n_276;
wire n_143;
wire n_431;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_513;
wire n_283;
wire n_107;
wire n_490;
wire n_517;
wire n_479;
wire n_415;
wire n_543;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_542;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_48;
wire n_465;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_221;
wire n_256;
wire n_454;
wire n_540;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_508;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_544;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_530;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_474;
wire n_539;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_511;
wire n_486;
wire n_305;
wire n_161;
wire n_441;
wire n_342;
wire n_101;
wire n_226;
wire n_509;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_510;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_536;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_537;
wire n_110;
wire n_531;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_523;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_533;
wire n_296;
wire n_384;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_491;
wire n_24;
wire n_526;
wire n_467;
wire n_269;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_473;
wire n_45;
wire n_520;
wire n_476;
wire n_337;
wire n_317;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_481;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_522;
wire n_333;
wire n_518;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_302;
wire n_216;
wire n_528;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_199;
wire n_260;
wire n_413;
wire n_275;
wire n_494;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_492;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_515;
wire n_347;
wire n_521;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_538;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_534;
wire n_472;
wire n_279;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_484;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_469;
wire n_111;
wire n_197;
wire n_396;
wire n_375;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_527;
wire n_482;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_512;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_516;
wire n_183;
wire n_409;
wire n_532;
wire n_249;
wire n_412;
wire n_217;
wire n_471;
wire n_541;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_535;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_524;
wire n_402;
wire n_504;
wire n_438;
wire n_475;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_514;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

CKINVDCx16_ASAP7_75t_R g19 ( 
.A(n_17),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_2),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_16),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_14),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_2),
.Y(n_23)
);

INVx6_ASAP7_75t_L g24 ( 
.A(n_13),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_16),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_8),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_0),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_5),
.Y(n_28)
);

BUFx12f_ASAP7_75t_L g29 ( 
.A(n_3),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_14),
.Y(n_30)
);

BUFx5_ASAP7_75t_L g31 ( 
.A(n_6),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_17),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_8),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_15),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_6),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_6),
.Y(n_36)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_1),
.Y(n_37)
);

BUFx3_ASAP7_75t_L g38 ( 
.A(n_1),
.Y(n_38)
);

BUFx5_ASAP7_75t_L g39 ( 
.A(n_15),
.Y(n_39)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_14),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_15),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_8),
.Y(n_42)
);

INVx13_ASAP7_75t_L g43 ( 
.A(n_15),
.Y(n_43)
);

INVx13_ASAP7_75t_L g44 ( 
.A(n_13),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_10),
.Y(n_45)
);

BUFx12f_ASAP7_75t_L g46 ( 
.A(n_11),
.Y(n_46)
);

CKINVDCx16_ASAP7_75t_R g47 ( 
.A(n_4),
.Y(n_47)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_13),
.Y(n_48)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_0),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_4),
.Y(n_50)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_18),
.Y(n_51)
);

BUFx3_ASAP7_75t_L g52 ( 
.A(n_31),
.Y(n_52)
);

INVx5_ASAP7_75t_L g126 ( 
.A(n_52),
.Y(n_126)
);

BUFx2_ASAP7_75t_L g53 ( 
.A(n_31),
.Y(n_53)
);

INVx3_ASAP7_75t_L g108 ( 
.A(n_53),
.Y(n_108)
);

BUFx3_ASAP7_75t_L g54 ( 
.A(n_31),
.Y(n_54)
);

INVx5_ASAP7_75t_L g133 ( 
.A(n_54),
.Y(n_133)
);

INVx2_ASAP7_75t_L g55 ( 
.A(n_24),
.Y(n_55)
);

INVx2_ASAP7_75t_L g106 ( 
.A(n_55),
.Y(n_106)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_24),
.Y(n_56)
);

INVx2_ASAP7_75t_L g119 ( 
.A(n_56),
.Y(n_119)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_27),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g124 ( 
.A(n_57),
.Y(n_124)
);

INVx8_ASAP7_75t_L g58 ( 
.A(n_39),
.Y(n_58)
);

INVx5_ASAP7_75t_L g137 ( 
.A(n_58),
.Y(n_137)
);

INVx6_ASAP7_75t_L g59 ( 
.A(n_27),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g127 ( 
.A(n_59),
.Y(n_127)
);

INVx11_ASAP7_75t_L g60 ( 
.A(n_27),
.Y(n_60)
);

INVx5_ASAP7_75t_L g147 ( 
.A(n_60),
.Y(n_147)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_24),
.Y(n_61)
);

INVx2_ASAP7_75t_L g131 ( 
.A(n_61),
.Y(n_131)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_27),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g130 ( 
.A(n_62),
.Y(n_130)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_28),
.Y(n_63)
);

BUFx6f_ASAP7_75t_L g138 ( 
.A(n_63),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_L g64 ( 
.A(n_25),
.B(n_18),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_L g139 ( 
.A(n_64),
.B(n_85),
.Y(n_139)
);

INVx2_ASAP7_75t_L g65 ( 
.A(n_21),
.Y(n_65)
);

INVx2_ASAP7_75t_L g132 ( 
.A(n_65),
.Y(n_132)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_21),
.Y(n_66)
);

INVx2_ASAP7_75t_L g143 ( 
.A(n_66),
.Y(n_143)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_28),
.Y(n_67)
);

BUFx6f_ASAP7_75t_L g146 ( 
.A(n_67),
.Y(n_146)
);

BUFx12f_ASAP7_75t_L g68 ( 
.A(n_43),
.Y(n_68)
);

INVx3_ASAP7_75t_L g112 ( 
.A(n_68),
.Y(n_112)
);

CKINVDCx20_ASAP7_75t_R g69 ( 
.A(n_38),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_69),
.B(n_78),
.Y(n_107)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_21),
.Y(n_70)
);

INVx2_ASAP7_75t_L g149 ( 
.A(n_70),
.Y(n_149)
);

INVx4_ASAP7_75t_L g71 ( 
.A(n_39),
.Y(n_71)
);

INVx4_ASAP7_75t_SL g123 ( 
.A(n_71),
.Y(n_123)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_37),
.Y(n_72)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_72),
.Y(n_105)
);

INVx4_ASAP7_75t_L g73 ( 
.A(n_39),
.Y(n_73)
);

INVx4_ASAP7_75t_L g104 ( 
.A(n_73),
.Y(n_104)
);

INVx6_ASAP7_75t_L g74 ( 
.A(n_28),
.Y(n_74)
);

BUFx6f_ASAP7_75t_L g148 ( 
.A(n_74),
.Y(n_148)
);

BUFx6f_ASAP7_75t_L g75 ( 
.A(n_28),
.Y(n_75)
);

INVx6_ASAP7_75t_L g110 ( 
.A(n_75),
.Y(n_110)
);

BUFx12f_ASAP7_75t_L g76 ( 
.A(n_43),
.Y(n_76)
);

INVx3_ASAP7_75t_L g154 ( 
.A(n_76),
.Y(n_154)
);

INVx3_ASAP7_75t_L g77 ( 
.A(n_38),
.Y(n_77)
);

INVx4_ASAP7_75t_L g111 ( 
.A(n_77),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_SL g78 ( 
.A(n_25),
.B(n_18),
.Y(n_78)
);

INVx2_ASAP7_75t_L g79 ( 
.A(n_21),
.Y(n_79)
);

INVx2_ASAP7_75t_L g153 ( 
.A(n_79),
.Y(n_153)
);

BUFx6f_ASAP7_75t_L g80 ( 
.A(n_30),
.Y(n_80)
);

INVx5_ASAP7_75t_L g162 ( 
.A(n_80),
.Y(n_162)
);

INVx8_ASAP7_75t_L g81 ( 
.A(n_30),
.Y(n_81)
);

BUFx3_ASAP7_75t_L g156 ( 
.A(n_81),
.Y(n_156)
);

BUFx6f_ASAP7_75t_L g82 ( 
.A(n_30),
.Y(n_82)
);

INVx4_ASAP7_75t_L g134 ( 
.A(n_82),
.Y(n_134)
);

BUFx3_ASAP7_75t_L g83 ( 
.A(n_38),
.Y(n_83)
);

INVx4_ASAP7_75t_L g145 ( 
.A(n_83),
.Y(n_145)
);

INVx6_ASAP7_75t_L g84 ( 
.A(n_30),
.Y(n_84)
);

INVx2_ASAP7_75t_L g155 ( 
.A(n_84),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_SL g85 ( 
.A(n_51),
.B(n_17),
.Y(n_85)
);

BUFx5_ASAP7_75t_L g86 ( 
.A(n_29),
.Y(n_86)
);

BUFx10_ASAP7_75t_L g113 ( 
.A(n_86),
.Y(n_113)
);

BUFx5_ASAP7_75t_L g87 ( 
.A(n_29),
.Y(n_87)
);

AND2x2_ASAP7_75t_L g128 ( 
.A(n_87),
.B(n_96),
.Y(n_128)
);

BUFx6f_ASAP7_75t_L g88 ( 
.A(n_36),
.Y(n_88)
);

INVx2_ASAP7_75t_L g161 ( 
.A(n_88),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_51),
.B(n_16),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g164 ( 
.A(n_89),
.B(n_91),
.Y(n_164)
);

INVx2_ASAP7_75t_L g90 ( 
.A(n_32),
.Y(n_90)
);

INVx2_ASAP7_75t_L g165 ( 
.A(n_90),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_L g91 ( 
.A(n_22),
.B(n_0),
.Y(n_91)
);

INVx6_ASAP7_75t_L g92 ( 
.A(n_36),
.Y(n_92)
);

INVx2_ASAP7_75t_L g166 ( 
.A(n_92),
.Y(n_166)
);

BUFx6f_ASAP7_75t_L g93 ( 
.A(n_36),
.Y(n_93)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_93),
.Y(n_109)
);

INVx2_ASAP7_75t_L g94 ( 
.A(n_32),
.Y(n_94)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_94),
.Y(n_115)
);

BUFx6f_ASAP7_75t_L g95 ( 
.A(n_36),
.Y(n_95)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_95),
.Y(n_120)
);

BUFx5_ASAP7_75t_L g96 ( 
.A(n_29),
.Y(n_96)
);

INVx2_ASAP7_75t_L g97 ( 
.A(n_32),
.Y(n_97)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_97),
.Y(n_122)
);

INVx2_ASAP7_75t_L g98 ( 
.A(n_32),
.Y(n_98)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_98),
.Y(n_135)
);

INVx6_ASAP7_75t_L g99 ( 
.A(n_41),
.Y(n_99)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_99),
.Y(n_136)
);

INVx3_ASAP7_75t_L g100 ( 
.A(n_29),
.Y(n_100)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_100),
.Y(n_142)
);

AOI22xp33_ASAP7_75t_L g101 ( 
.A1(n_41),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_101)
);

OAI22xp5_ASAP7_75t_L g141 ( 
.A1(n_101),
.A2(n_47),
.B1(n_48),
.B2(n_35),
.Y(n_141)
);

BUFx6f_ASAP7_75t_L g102 ( 
.A(n_41),
.Y(n_102)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_102),
.Y(n_144)
);

HAxp5_ASAP7_75t_SL g103 ( 
.A(n_47),
.B(n_1),
.CON(n_103),
.SN(n_103)
);

AND2x2_ASAP7_75t_L g160 ( 
.A(n_103),
.B(n_20),
.Y(n_160)
);

NOR2xp33_ASAP7_75t_L g114 ( 
.A(n_68),
.B(n_19),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g181 ( 
.A(n_114),
.B(n_118),
.Y(n_181)
);

MAJIxp5_ASAP7_75t_L g116 ( 
.A(n_83),
.B(n_37),
.C(n_19),
.Y(n_116)
);

MAJIxp5_ASAP7_75t_L g218 ( 
.A(n_116),
.B(n_44),
.C(n_4),
.Y(n_218)
);

AOI21xp33_ASAP7_75t_SL g117 ( 
.A1(n_103),
.A2(n_29),
.B(n_46),
.Y(n_117)
);

AND2x2_ASAP7_75t_L g169 ( 
.A(n_117),
.B(n_121),
.Y(n_169)
);

NOR2xp33_ASAP7_75t_L g118 ( 
.A(n_68),
.B(n_50),
.Y(n_118)
);

NAND2x1_ASAP7_75t_L g121 ( 
.A(n_101),
.B(n_43),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_L g125 ( 
.A(n_76),
.B(n_50),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_L g182 ( 
.A(n_125),
.B(n_152),
.Y(n_182)
);

AOI22xp33_ASAP7_75t_SL g129 ( 
.A1(n_53),
.A2(n_29),
.B1(n_46),
.B2(n_41),
.Y(n_129)
);

OAI22xp5_ASAP7_75t_L g173 ( 
.A1(n_129),
.A2(n_140),
.B1(n_163),
.B2(n_74),
.Y(n_173)
);

AOI22xp33_ASAP7_75t_SL g140 ( 
.A1(n_81),
.A2(n_46),
.B1(n_42),
.B2(n_48),
.Y(n_140)
);

AOI22xp5_ASAP7_75t_L g201 ( 
.A1(n_141),
.A2(n_157),
.B1(n_23),
.B2(n_22),
.Y(n_201)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_60),
.Y(n_150)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_150),
.Y(n_193)
);

NAND2xp33_ASAP7_75t_SL g151 ( 
.A(n_73),
.B(n_48),
.Y(n_151)
);

OR2x2_ASAP7_75t_L g189 ( 
.A(n_151),
.B(n_159),
.Y(n_189)
);

NOR2xp33_ASAP7_75t_L g152 ( 
.A(n_76),
.B(n_49),
.Y(n_152)
);

OAI22xp5_ASAP7_75t_L g157 ( 
.A1(n_57),
.A2(n_49),
.B1(n_45),
.B2(n_34),
.Y(n_157)
);

NOR2xp33_ASAP7_75t_L g158 ( 
.A(n_52),
.B(n_45),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_L g212 ( 
.A(n_158),
.B(n_2),
.Y(n_212)
);

AOI21xp33_ASAP7_75t_L g159 ( 
.A1(n_54),
.A2(n_20),
.B(n_26),
.Y(n_159)
);

AND2x2_ASAP7_75t_L g206 ( 
.A(n_160),
.B(n_88),
.Y(n_206)
);

AOI22xp33_ASAP7_75t_SL g163 ( 
.A1(n_58),
.A2(n_46),
.B1(n_42),
.B2(n_40),
.Y(n_163)
);

INVx6_ASAP7_75t_L g167 ( 
.A(n_124),
.Y(n_167)
);

BUFx2_ASAP7_75t_L g241 ( 
.A(n_167),
.Y(n_241)
);

AOI22xp33_ASAP7_75t_SL g168 ( 
.A1(n_121),
.A2(n_46),
.B1(n_42),
.B2(n_40),
.Y(n_168)
);

INVxp67_ASAP7_75t_L g279 ( 
.A(n_168),
.Y(n_279)
);

INVx11_ASAP7_75t_L g170 ( 
.A(n_137),
.Y(n_170)
);

BUFx6f_ASAP7_75t_L g238 ( 
.A(n_170),
.Y(n_238)
);

INVx2_ASAP7_75t_L g171 ( 
.A(n_132),
.Y(n_171)
);

INVx2_ASAP7_75t_L g245 ( 
.A(n_171),
.Y(n_245)
);

AND2x2_ASAP7_75t_SL g172 ( 
.A(n_164),
.B(n_59),
.Y(n_172)
);

AND2x2_ASAP7_75t_L g277 ( 
.A(n_172),
.B(n_173),
.Y(n_277)
);

BUFx3_ASAP7_75t_L g174 ( 
.A(n_154),
.Y(n_174)
);

INVx4_ASAP7_75t_L g258 ( 
.A(n_174),
.Y(n_258)
);

AOI22xp33_ASAP7_75t_SL g175 ( 
.A1(n_123),
.A2(n_46),
.B1(n_42),
.B2(n_40),
.Y(n_175)
);

AOI22xp33_ASAP7_75t_SL g243 ( 
.A1(n_175),
.A2(n_177),
.B1(n_196),
.B2(n_200),
.Y(n_243)
);

NAND2xp5_ASAP7_75t_SL g176 ( 
.A(n_139),
.B(n_34),
.Y(n_176)
);

NOR2xp33_ASAP7_75t_L g251 ( 
.A(n_176),
.B(n_188),
.Y(n_251)
);

AOI22xp33_ASAP7_75t_SL g177 ( 
.A1(n_123),
.A2(n_33),
.B1(n_20),
.B2(n_26),
.Y(n_177)
);

BUFx6f_ASAP7_75t_L g178 ( 
.A(n_124),
.Y(n_178)
);

BUFx6f_ASAP7_75t_L g262 ( 
.A(n_178),
.Y(n_262)
);

INVx2_ASAP7_75t_L g179 ( 
.A(n_106),
.Y(n_179)
);

INVx2_ASAP7_75t_L g255 ( 
.A(n_179),
.Y(n_255)
);

INVx6_ASAP7_75t_L g180 ( 
.A(n_130),
.Y(n_180)
);

INVx6_ASAP7_75t_L g260 ( 
.A(n_180),
.Y(n_260)
);

INVx2_ASAP7_75t_L g183 ( 
.A(n_119),
.Y(n_183)
);

INVx2_ASAP7_75t_L g257 ( 
.A(n_183),
.Y(n_257)
);

BUFx2_ASAP7_75t_L g184 ( 
.A(n_145),
.Y(n_184)
);

CKINVDCx20_ASAP7_75t_R g233 ( 
.A(n_184),
.Y(n_233)
);

BUFx8_ASAP7_75t_L g185 ( 
.A(n_156),
.Y(n_185)
);

INVx8_ASAP7_75t_L g230 ( 
.A(n_185),
.Y(n_230)
);

INVx2_ASAP7_75t_L g186 ( 
.A(n_143),
.Y(n_186)
);

INVx4_ASAP7_75t_L g269 ( 
.A(n_186),
.Y(n_269)
);

INVxp33_ASAP7_75t_L g187 ( 
.A(n_113),
.Y(n_187)
);

INVx13_ASAP7_75t_L g228 ( 
.A(n_187),
.Y(n_228)
);

CKINVDCx16_ASAP7_75t_R g188 ( 
.A(n_128),
.Y(n_188)
);

BUFx6f_ASAP7_75t_L g190 ( 
.A(n_130),
.Y(n_190)
);

INVx8_ASAP7_75t_L g234 ( 
.A(n_190),
.Y(n_234)
);

INVx3_ASAP7_75t_L g191 ( 
.A(n_154),
.Y(n_191)
);

INVx8_ASAP7_75t_L g247 ( 
.A(n_191),
.Y(n_247)
);

INVx2_ASAP7_75t_L g192 ( 
.A(n_131),
.Y(n_192)
);

HB1xp67_ASAP7_75t_L g271 ( 
.A(n_192),
.Y(n_271)
);

INVxp67_ASAP7_75t_L g194 ( 
.A(n_128),
.Y(n_194)
);

NOR2xp33_ASAP7_75t_L g276 ( 
.A(n_194),
.B(n_195),
.Y(n_276)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_105),
.Y(n_195)
);

AOI22xp33_ASAP7_75t_SL g196 ( 
.A1(n_111),
.A2(n_35),
.B1(n_26),
.B2(n_33),
.Y(n_196)
);

INVx8_ASAP7_75t_L g197 ( 
.A(n_112),
.Y(n_197)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_197),
.Y(n_235)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_115),
.Y(n_198)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_198),
.Y(n_237)
);

BUFx6f_ASAP7_75t_L g199 ( 
.A(n_138),
.Y(n_199)
);

BUFx12f_ASAP7_75t_L g275 ( 
.A(n_199),
.Y(n_275)
);

AOI22xp33_ASAP7_75t_SL g200 ( 
.A1(n_111),
.A2(n_35),
.B1(n_33),
.B2(n_23),
.Y(n_200)
);

OAI22xp5_ASAP7_75t_SL g236 ( 
.A1(n_201),
.A2(n_203),
.B1(n_223),
.B2(n_140),
.Y(n_236)
);

NOR2xp33_ASAP7_75t_L g202 ( 
.A(n_107),
.B(n_44),
.Y(n_202)
);

NOR2xp33_ASAP7_75t_L g229 ( 
.A(n_202),
.B(n_207),
.Y(n_229)
);

OAI22xp5_ASAP7_75t_SL g203 ( 
.A1(n_129),
.A2(n_84),
.B1(n_99),
.B2(n_92),
.Y(n_203)
);

INVx2_ASAP7_75t_L g204 ( 
.A(n_149),
.Y(n_204)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_204),
.Y(n_248)
);

AOI22xp33_ASAP7_75t_SL g205 ( 
.A1(n_126),
.A2(n_102),
.B1(n_95),
.B2(n_93),
.Y(n_205)
);

AOI22xp33_ASAP7_75t_SL g264 ( 
.A1(n_205),
.A2(n_208),
.B1(n_220),
.B2(n_225),
.Y(n_264)
);

XNOR2xp5_ASAP7_75t_SL g240 ( 
.A(n_206),
.B(n_218),
.Y(n_240)
);

BUFx4f_ASAP7_75t_SL g207 ( 
.A(n_126),
.Y(n_207)
);

AOI22xp33_ASAP7_75t_SL g208 ( 
.A1(n_133),
.A2(n_82),
.B1(n_80),
.B2(n_75),
.Y(n_208)
);

BUFx6f_ASAP7_75t_L g209 ( 
.A(n_138),
.Y(n_209)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_209),
.Y(n_256)
);

A2O1A1O1Ixp25_ASAP7_75t_L g210 ( 
.A1(n_160),
.A2(n_44),
.B(n_43),
.C(n_62),
.D(n_67),
.Y(n_210)
);

NOR2xp33_ASAP7_75t_L g231 ( 
.A(n_210),
.B(n_212),
.Y(n_231)
);

INVx4_ASAP7_75t_L g211 ( 
.A(n_104),
.Y(n_211)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_211),
.Y(n_261)
);

HB1xp67_ASAP7_75t_L g213 ( 
.A(n_142),
.Y(n_213)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_213),
.Y(n_265)
);

OAI21xp33_ASAP7_75t_L g214 ( 
.A1(n_145),
.A2(n_104),
.B(n_122),
.Y(n_214)
);

OAI21xp5_ASAP7_75t_L g263 ( 
.A1(n_214),
.A2(n_113),
.B(n_147),
.Y(n_263)
);

NOR2xp33_ASAP7_75t_L g215 ( 
.A(n_108),
.B(n_44),
.Y(n_215)
);

NOR2xp33_ASAP7_75t_L g246 ( 
.A(n_215),
.B(n_221),
.Y(n_246)
);

AOI22xp5_ASAP7_75t_L g216 ( 
.A1(n_135),
.A2(n_63),
.B1(n_4),
.B2(n_5),
.Y(n_216)
);

OAI22xp5_ASAP7_75t_L g239 ( 
.A1(n_216),
.A2(n_110),
.B1(n_120),
.B2(n_134),
.Y(n_239)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_136),
.Y(n_217)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_217),
.Y(n_266)
);

BUFx6f_ASAP7_75t_L g219 ( 
.A(n_146),
.Y(n_219)
);

INVx2_ASAP7_75t_SL g278 ( 
.A(n_219),
.Y(n_278)
);

AOI22xp33_ASAP7_75t_SL g220 ( 
.A1(n_133),
.A2(n_3),
.B1(n_5),
.B2(n_6),
.Y(n_220)
);

BUFx3_ASAP7_75t_L g221 ( 
.A(n_137),
.Y(n_221)
);

INVx2_ASAP7_75t_L g222 ( 
.A(n_153),
.Y(n_222)
);

NOR2xp33_ASAP7_75t_L g249 ( 
.A(n_222),
.B(n_224),
.Y(n_249)
);

OA22x2_ASAP7_75t_L g223 ( 
.A1(n_163),
.A2(n_3),
.B1(n_5),
.B2(n_7),
.Y(n_223)
);

INVx2_ASAP7_75t_L g224 ( 
.A(n_165),
.Y(n_224)
);

AOI22xp33_ASAP7_75t_SL g225 ( 
.A1(n_134),
.A2(n_3),
.B1(n_7),
.B2(n_8),
.Y(n_225)
);

INVx2_ASAP7_75t_L g226 ( 
.A(n_155),
.Y(n_226)
);

NOR2xp33_ASAP7_75t_L g250 ( 
.A(n_226),
.B(n_227),
.Y(n_250)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_109),
.Y(n_227)
);

NAND2xp5_ASAP7_75t_L g232 ( 
.A(n_172),
.B(n_144),
.Y(n_232)
);

NAND2xp5_ASAP7_75t_L g280 ( 
.A(n_232),
.B(n_206),
.Y(n_280)
);

AOI22xp5_ASAP7_75t_L g290 ( 
.A1(n_236),
.A2(n_239),
.B1(n_242),
.B2(n_253),
.Y(n_290)
);

OAI22xp5_ASAP7_75t_SL g242 ( 
.A1(n_189),
.A2(n_166),
.B1(n_161),
.B2(n_148),
.Y(n_242)
);

AOI22xp33_ASAP7_75t_L g244 ( 
.A1(n_201),
.A2(n_162),
.B1(n_110),
.B2(n_148),
.Y(n_244)
);

OAI22xp5_ASAP7_75t_SL g301 ( 
.A1(n_244),
.A2(n_259),
.B1(n_279),
.B2(n_264),
.Y(n_301)
);

NOR2xp33_ASAP7_75t_L g252 ( 
.A(n_182),
.B(n_156),
.Y(n_252)
);

NOR2xp33_ASAP7_75t_SL g295 ( 
.A(n_252),
.B(n_270),
.Y(n_295)
);

OAI22xp5_ASAP7_75t_SL g253 ( 
.A1(n_189),
.A2(n_127),
.B1(n_146),
.B2(n_162),
.Y(n_253)
);

NOR2xp33_ASAP7_75t_SL g254 ( 
.A(n_181),
.B(n_7),
.Y(n_254)
);

NAND2xp5_ASAP7_75t_SL g289 ( 
.A(n_254),
.B(n_268),
.Y(n_289)
);

AOI22xp33_ASAP7_75t_L g259 ( 
.A1(n_169),
.A2(n_127),
.B1(n_147),
.B2(n_113),
.Y(n_259)
);

AND2x2_ASAP7_75t_L g298 ( 
.A(n_263),
.B(n_223),
.Y(n_298)
);

OAI22xp5_ASAP7_75t_L g267 ( 
.A1(n_172),
.A2(n_169),
.B1(n_216),
.B2(n_206),
.Y(n_267)
);

AOI22xp5_ASAP7_75t_L g300 ( 
.A1(n_267),
.A2(n_273),
.B1(n_223),
.B2(n_180),
.Y(n_300)
);

NOR2xp33_ASAP7_75t_SL g268 ( 
.A(n_194),
.B(n_7),
.Y(n_268)
);

NOR2xp33_ASAP7_75t_L g270 ( 
.A(n_193),
.B(n_218),
.Y(n_270)
);

NOR2xp33_ASAP7_75t_L g272 ( 
.A(n_191),
.B(n_9),
.Y(n_272)
);

NOR2xp33_ASAP7_75t_SL g310 ( 
.A(n_272),
.B(n_185),
.Y(n_310)
);

OAI22xp5_ASAP7_75t_SL g273 ( 
.A1(n_169),
.A2(n_9),
.B1(n_10),
.B2(n_11),
.Y(n_273)
);

AOI22xp33_ASAP7_75t_SL g274 ( 
.A1(n_223),
.A2(n_9),
.B1(n_10),
.B2(n_11),
.Y(n_274)
);

INVxp67_ASAP7_75t_L g287 ( 
.A(n_274),
.Y(n_287)
);

NAND2xp5_ASAP7_75t_L g336 ( 
.A(n_280),
.B(n_286),
.Y(n_336)
);

AND2x2_ASAP7_75t_SL g281 ( 
.A(n_232),
.B(n_214),
.Y(n_281)
);

INVxp67_ASAP7_75t_L g349 ( 
.A(n_281),
.Y(n_349)
);

NOR2xp33_ASAP7_75t_L g282 ( 
.A(n_254),
.B(n_197),
.Y(n_282)
);

CKINVDCx14_ASAP7_75t_R g351 ( 
.A(n_282),
.Y(n_351)
);

CKINVDCx16_ASAP7_75t_R g283 ( 
.A(n_229),
.Y(n_283)
);

NOR2xp33_ASAP7_75t_L g339 ( 
.A(n_283),
.B(n_284),
.Y(n_339)
);

NOR2xp33_ASAP7_75t_L g284 ( 
.A(n_276),
.B(n_174),
.Y(n_284)
);

OAI21xp5_ASAP7_75t_SL g285 ( 
.A1(n_277),
.A2(n_267),
.B(n_243),
.Y(n_285)
);

OAI21xp5_ASAP7_75t_SL g365 ( 
.A1(n_285),
.A2(n_298),
.B(n_304),
.Y(n_365)
);

NAND2xp5_ASAP7_75t_L g286 ( 
.A(n_277),
.B(n_171),
.Y(n_286)
);

INVxp67_ASAP7_75t_L g288 ( 
.A(n_263),
.Y(n_288)
);

NOR2xp33_ASAP7_75t_L g345 ( 
.A(n_288),
.B(n_299),
.Y(n_345)
);

MAJIxp5_ASAP7_75t_L g291 ( 
.A(n_240),
.B(n_277),
.C(n_231),
.Y(n_291)
);

MAJIxp5_ASAP7_75t_L g331 ( 
.A(n_291),
.B(n_308),
.C(n_293),
.Y(n_331)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_266),
.Y(n_292)
);

INVx1_ASAP7_75t_L g343 ( 
.A(n_292),
.Y(n_343)
);

FAx1_ASAP7_75t_SL g293 ( 
.A(n_240),
.B(n_210),
.CI(n_203),
.CON(n_293),
.SN(n_293)
);

NOR2xp33_ASAP7_75t_SL g347 ( 
.A(n_293),
.B(n_310),
.Y(n_347)
);

NAND2xp5_ASAP7_75t_L g294 ( 
.A(n_273),
.B(n_186),
.Y(n_294)
);

NAND2xp5_ASAP7_75t_L g348 ( 
.A(n_294),
.B(n_297),
.Y(n_348)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_248),
.Y(n_296)
);

NAND2xp5_ASAP7_75t_SL g330 ( 
.A(n_296),
.B(n_305),
.Y(n_330)
);

NAND2xp5_ASAP7_75t_L g297 ( 
.A(n_236),
.B(n_204),
.Y(n_297)
);

INVxp67_ASAP7_75t_L g299 ( 
.A(n_246),
.Y(n_299)
);

NAND2xp5_ASAP7_75t_L g353 ( 
.A(n_300),
.B(n_315),
.Y(n_353)
);

AOI22xp5_ASAP7_75t_L g338 ( 
.A1(n_301),
.A2(n_314),
.B1(n_241),
.B2(n_230),
.Y(n_338)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_266),
.Y(n_302)
);

NOR2xp33_ASAP7_75t_L g354 ( 
.A(n_302),
.B(n_306),
.Y(n_354)
);

AOI22xp33_ASAP7_75t_SL g303 ( 
.A1(n_279),
.A2(n_184),
.B1(n_221),
.B2(n_211),
.Y(n_303)
);

INVxp67_ASAP7_75t_L g362 ( 
.A(n_303),
.Y(n_362)
);

AOI22xp33_ASAP7_75t_SL g304 ( 
.A1(n_230),
.A2(n_167),
.B1(n_178),
.B2(n_219),
.Y(n_304)
);

NAND2xp5_ASAP7_75t_SL g305 ( 
.A(n_251),
.B(n_224),
.Y(n_305)
);

NOR2xp33_ASAP7_75t_L g306 ( 
.A(n_276),
.B(n_187),
.Y(n_306)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_237),
.Y(n_307)
);

CKINVDCx20_ASAP7_75t_R g333 ( 
.A(n_307),
.Y(n_333)
);

XOR2xp5_ASAP7_75t_L g308 ( 
.A(n_242),
.B(n_207),
.Y(n_308)
);

INVx3_ASAP7_75t_L g309 ( 
.A(n_275),
.Y(n_309)
);

INVxp33_ASAP7_75t_L g341 ( 
.A(n_309),
.Y(n_341)
);

CKINVDCx20_ASAP7_75t_R g311 ( 
.A(n_249),
.Y(n_311)
);

CKINVDCx20_ASAP7_75t_R g364 ( 
.A(n_311),
.Y(n_364)
);

INVx4_ASAP7_75t_L g312 ( 
.A(n_230),
.Y(n_312)
);

CKINVDCx20_ASAP7_75t_R g367 ( 
.A(n_312),
.Y(n_367)
);

INVx3_ASAP7_75t_L g313 ( 
.A(n_275),
.Y(n_313)
);

CKINVDCx20_ASAP7_75t_R g368 ( 
.A(n_313),
.Y(n_368)
);

OAI22xp5_ASAP7_75t_SL g314 ( 
.A1(n_253),
.A2(n_226),
.B1(n_209),
.B2(n_199),
.Y(n_314)
);

BUFx12f_ASAP7_75t_L g315 ( 
.A(n_228),
.Y(n_315)
);

NAND2xp5_ASAP7_75t_L g316 ( 
.A(n_268),
.B(n_250),
.Y(n_316)
);

NAND2xp5_ASAP7_75t_L g358 ( 
.A(n_316),
.B(n_318),
.Y(n_358)
);

AOI22xp5_ASAP7_75t_L g317 ( 
.A1(n_239),
.A2(n_190),
.B1(n_170),
.B2(n_207),
.Y(n_317)
);

OAI22xp5_ASAP7_75t_SL g328 ( 
.A1(n_317),
.A2(n_321),
.B1(n_323),
.B2(n_278),
.Y(n_328)
);

INVx2_ASAP7_75t_L g318 ( 
.A(n_245),
.Y(n_318)
);

NAND2xp5_ASAP7_75t_L g319 ( 
.A(n_237),
.B(n_185),
.Y(n_319)
);

NAND2xp5_ASAP7_75t_L g363 ( 
.A(n_319),
.B(n_322),
.Y(n_363)
);

AOI22xp5_ASAP7_75t_SL g320 ( 
.A1(n_235),
.A2(n_9),
.B1(n_10),
.B2(n_11),
.Y(n_320)
);

AOI32xp33_ASAP7_75t_L g361 ( 
.A1(n_320),
.A2(n_258),
.A3(n_12),
.B1(n_247),
.B2(n_238),
.Y(n_361)
);

AOI22xp5_ASAP7_75t_L g321 ( 
.A1(n_251),
.A2(n_12),
.B1(n_13),
.B2(n_14),
.Y(n_321)
);

INVx3_ASAP7_75t_L g322 ( 
.A(n_275),
.Y(n_322)
);

AOI22xp5_ASAP7_75t_L g323 ( 
.A1(n_265),
.A2(n_12),
.B1(n_248),
.B2(n_235),
.Y(n_323)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_265),
.Y(n_324)
);

NAND2xp5_ASAP7_75t_SL g335 ( 
.A(n_324),
.B(n_325),
.Y(n_335)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_245),
.Y(n_325)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_271),
.Y(n_326)
);

NAND2xp5_ASAP7_75t_SL g337 ( 
.A(n_326),
.B(n_233),
.Y(n_337)
);

INVx3_ASAP7_75t_L g327 ( 
.A(n_275),
.Y(n_327)
);

NAND2xp5_ASAP7_75t_L g369 ( 
.A(n_327),
.B(n_12),
.Y(n_369)
);

AOI22xp5_ASAP7_75t_L g375 ( 
.A1(n_328),
.A2(n_329),
.B1(n_332),
.B2(n_334),
.Y(n_375)
);

OAI22xp5_ASAP7_75t_SL g329 ( 
.A1(n_297),
.A2(n_278),
.B1(n_256),
.B2(n_260),
.Y(n_329)
);

XOR2xp5_ASAP7_75t_L g389 ( 
.A(n_331),
.B(n_346),
.Y(n_389)
);

OAI22xp5_ASAP7_75t_L g332 ( 
.A1(n_290),
.A2(n_256),
.B1(n_278),
.B2(n_260),
.Y(n_332)
);

OAI22xp5_ASAP7_75t_SL g334 ( 
.A1(n_290),
.A2(n_260),
.B1(n_241),
.B2(n_234),
.Y(n_334)
);

INVxp67_ASAP7_75t_L g402 ( 
.A(n_337),
.Y(n_402)
);

AOI22xp33_ASAP7_75t_L g373 ( 
.A1(n_338),
.A2(n_344),
.B1(n_350),
.B2(n_359),
.Y(n_373)
);

XNOR2xp5_ASAP7_75t_L g340 ( 
.A(n_291),
.B(n_261),
.Y(n_340)
);

MAJIxp5_ASAP7_75t_L g391 ( 
.A(n_340),
.B(n_356),
.C(n_322),
.Y(n_391)
);

AOI21xp5_ASAP7_75t_SL g342 ( 
.A1(n_288),
.A2(n_261),
.B(n_228),
.Y(n_342)
);

OAI21xp5_ASAP7_75t_SL g379 ( 
.A1(n_342),
.A2(n_325),
.B(n_323),
.Y(n_379)
);

OAI22xp5_ASAP7_75t_L g344 ( 
.A1(n_300),
.A2(n_241),
.B1(n_234),
.B2(n_262),
.Y(n_344)
);

MAJx2_ASAP7_75t_L g346 ( 
.A(n_285),
.B(n_228),
.C(n_233),
.Y(n_346)
);

OAI22xp5_ASAP7_75t_L g350 ( 
.A1(n_298),
.A2(n_286),
.B1(n_287),
.B2(n_281),
.Y(n_350)
);

AOI22xp5_ASAP7_75t_L g352 ( 
.A1(n_301),
.A2(n_269),
.B1(n_234),
.B2(n_262),
.Y(n_352)
);

OAI22xp5_ASAP7_75t_L g378 ( 
.A1(n_352),
.A2(n_357),
.B1(n_360),
.B2(n_338),
.Y(n_378)
);

OAI22xp5_ASAP7_75t_SL g355 ( 
.A1(n_287),
.A2(n_293),
.B1(n_298),
.B2(n_294),
.Y(n_355)
);

NAND2xp5_ASAP7_75t_L g376 ( 
.A(n_355),
.B(n_366),
.Y(n_376)
);

MAJIxp5_ASAP7_75t_L g356 ( 
.A(n_295),
.B(n_257),
.C(n_255),
.Y(n_356)
);

AOI22xp5_ASAP7_75t_L g357 ( 
.A1(n_308),
.A2(n_269),
.B1(n_262),
.B2(n_257),
.Y(n_357)
);

OAI22xp5_ASAP7_75t_L g359 ( 
.A1(n_281),
.A2(n_255),
.B1(n_247),
.B2(n_238),
.Y(n_359)
);

OAI22xp5_ASAP7_75t_L g360 ( 
.A1(n_317),
.A2(n_247),
.B1(n_238),
.B2(n_258),
.Y(n_360)
);

OAI21xp33_ASAP7_75t_SL g372 ( 
.A1(n_361),
.A2(n_320),
.B(n_280),
.Y(n_372)
);

OAI22xp33_ASAP7_75t_SL g366 ( 
.A1(n_299),
.A2(n_314),
.B1(n_316),
.B2(n_312),
.Y(n_366)
);

CKINVDCx20_ASAP7_75t_R g382 ( 
.A(n_369),
.Y(n_382)
);

INVx1_ASAP7_75t_L g370 ( 
.A(n_343),
.Y(n_370)
);

INVx1_ASAP7_75t_L g415 ( 
.A(n_370),
.Y(n_415)
);

NOR2xp33_ASAP7_75t_L g371 ( 
.A(n_364),
.B(n_319),
.Y(n_371)
);

INVxp33_ASAP7_75t_L g409 ( 
.A(n_371),
.Y(n_409)
);

AOI22xp5_ASAP7_75t_L g433 ( 
.A1(n_372),
.A2(n_378),
.B1(n_400),
.B2(n_398),
.Y(n_433)
);

INVx1_ASAP7_75t_L g374 ( 
.A(n_343),
.Y(n_374)
);

INVx1_ASAP7_75t_L g427 ( 
.A(n_374),
.Y(n_427)
);

NOR2xp33_ASAP7_75t_L g377 ( 
.A(n_364),
.B(n_296),
.Y(n_377)
);

CKINVDCx20_ASAP7_75t_R g428 ( 
.A(n_377),
.Y(n_428)
);

AOI21xp5_ASAP7_75t_L g417 ( 
.A1(n_379),
.A2(n_387),
.B(n_329),
.Y(n_417)
);

INVx1_ASAP7_75t_L g380 ( 
.A(n_335),
.Y(n_380)
);

INVx1_ASAP7_75t_L g429 ( 
.A(n_380),
.Y(n_429)
);

OAI21xp5_ASAP7_75t_L g381 ( 
.A1(n_349),
.A2(n_289),
.B(n_321),
.Y(n_381)
);

OAI21xp5_ASAP7_75t_L g432 ( 
.A1(n_381),
.A2(n_371),
.B(n_377),
.Y(n_432)
);

NAND2xp5_ASAP7_75t_L g383 ( 
.A(n_330),
.B(n_318),
.Y(n_383)
);

INVx1_ASAP7_75t_L g435 ( 
.A(n_383),
.Y(n_435)
);

NAND2xp5_ASAP7_75t_L g384 ( 
.A(n_330),
.B(n_315),
.Y(n_384)
);

NAND2xp5_ASAP7_75t_L g414 ( 
.A(n_384),
.B(n_385),
.Y(n_414)
);

NAND2xp5_ASAP7_75t_L g385 ( 
.A(n_358),
.B(n_315),
.Y(n_385)
);

NAND2xp5_ASAP7_75t_L g386 ( 
.A(n_358),
.B(n_315),
.Y(n_386)
);

NAND2xp5_ASAP7_75t_SL g413 ( 
.A(n_386),
.B(n_388),
.Y(n_413)
);

NAND2x1_ASAP7_75t_SL g387 ( 
.A(n_350),
.B(n_342),
.Y(n_387)
);

NAND2xp5_ASAP7_75t_L g388 ( 
.A(n_348),
.B(n_309),
.Y(n_388)
);

XOR2xp5_ASAP7_75t_L g390 ( 
.A(n_331),
.B(n_313),
.Y(n_390)
);

MAJIxp5_ASAP7_75t_L g419 ( 
.A(n_390),
.B(n_391),
.C(n_393),
.Y(n_419)
);

INVx1_ASAP7_75t_L g392 ( 
.A(n_335),
.Y(n_392)
);

CKINVDCx16_ASAP7_75t_R g407 ( 
.A(n_392),
.Y(n_407)
);

MAJIxp5_ASAP7_75t_L g393 ( 
.A(n_340),
.B(n_327),
.C(n_336),
.Y(n_393)
);

CKINVDCx20_ASAP7_75t_R g394 ( 
.A(n_363),
.Y(n_394)
);

CKINVDCx5p33_ASAP7_75t_R g405 ( 
.A(n_394),
.Y(n_405)
);

AOI22xp33_ASAP7_75t_SL g395 ( 
.A1(n_351),
.A2(n_362),
.B1(n_367),
.B2(n_368),
.Y(n_395)
);

OAI22xp5_ASAP7_75t_SL g406 ( 
.A1(n_395),
.A2(n_352),
.B1(n_353),
.B2(n_357),
.Y(n_406)
);

XOR2xp5_ASAP7_75t_L g396 ( 
.A(n_355),
.B(n_336),
.Y(n_396)
);

MAJIxp5_ASAP7_75t_L g422 ( 
.A(n_396),
.B(n_367),
.C(n_328),
.Y(n_422)
);

NAND2xp5_ASAP7_75t_L g397 ( 
.A(n_348),
.B(n_363),
.Y(n_397)
);

NAND2xp5_ASAP7_75t_SL g423 ( 
.A(n_397),
.B(n_399),
.Y(n_423)
);

INVx1_ASAP7_75t_L g398 ( 
.A(n_337),
.Y(n_398)
);

INVxp67_ASAP7_75t_L g431 ( 
.A(n_398),
.Y(n_431)
);

NAND2xp5_ASAP7_75t_L g399 ( 
.A(n_354),
.B(n_345),
.Y(n_399)
);

INVx1_ASAP7_75t_L g400 ( 
.A(n_359),
.Y(n_400)
);

NOR2xp33_ASAP7_75t_L g411 ( 
.A(n_400),
.B(n_401),
.Y(n_411)
);

INVx1_ASAP7_75t_L g401 ( 
.A(n_369),
.Y(n_401)
);

INVx1_ASAP7_75t_L g403 ( 
.A(n_339),
.Y(n_403)
);

NOR2xp33_ASAP7_75t_L g421 ( 
.A(n_403),
.B(n_333),
.Y(n_421)
);

OR2x2_ASAP7_75t_L g404 ( 
.A(n_333),
.B(n_342),
.Y(n_404)
);

OR2x2_ASAP7_75t_L g430 ( 
.A(n_404),
.B(n_394),
.Y(n_430)
);

AOI22xp5_ASAP7_75t_L g460 ( 
.A1(n_406),
.A2(n_408),
.B1(n_372),
.B2(n_370),
.Y(n_460)
);

OAI22xp5_ASAP7_75t_SL g408 ( 
.A1(n_373),
.A2(n_353),
.B1(n_365),
.B2(n_344),
.Y(n_408)
);

FAx1_ASAP7_75t_SL g410 ( 
.A(n_396),
.B(n_347),
.CI(n_346),
.CON(n_410),
.SN(n_410)
);

NOR2xp33_ASAP7_75t_SL g451 ( 
.A(n_410),
.B(n_381),
.Y(n_451)
);

AOI22xp5_ASAP7_75t_SL g412 ( 
.A1(n_378),
.A2(n_332),
.B1(n_365),
.B2(n_334),
.Y(n_412)
);

AND2x2_ASAP7_75t_L g455 ( 
.A(n_412),
.B(n_375),
.Y(n_455)
);

XOR2xp5_ASAP7_75t_L g416 ( 
.A(n_389),
.B(n_346),
.Y(n_416)
);

XOR2xp5_ASAP7_75t_L g456 ( 
.A(n_416),
.B(n_418),
.Y(n_456)
);

OAI21xp5_ASAP7_75t_L g444 ( 
.A1(n_417),
.A2(n_434),
.B(n_386),
.Y(n_444)
);

XOR2xp5_ASAP7_75t_L g418 ( 
.A(n_389),
.B(n_356),
.Y(n_418)
);

XOR2xp5_ASAP7_75t_L g420 ( 
.A(n_393),
.B(n_347),
.Y(n_420)
);

XOR2xp5_ASAP7_75t_L g458 ( 
.A(n_420),
.B(n_422),
.Y(n_458)
);

NAND2xp5_ASAP7_75t_SL g437 ( 
.A(n_421),
.B(n_402),
.Y(n_437)
);

MAJIxp5_ASAP7_75t_L g424 ( 
.A(n_390),
.B(n_368),
.C(n_360),
.Y(n_424)
);

MAJIxp5_ASAP7_75t_L g440 ( 
.A(n_424),
.B(n_425),
.C(n_376),
.Y(n_440)
);

XOR2xp5_ASAP7_75t_L g425 ( 
.A(n_391),
.B(n_361),
.Y(n_425)
);

XNOR2x2_ASAP7_75t_L g426 ( 
.A(n_387),
.B(n_341),
.Y(n_426)
);

AO21x1_ASAP7_75t_L g442 ( 
.A1(n_426),
.A2(n_432),
.B(n_404),
.Y(n_442)
);

INVx1_ASAP7_75t_L g443 ( 
.A(n_430),
.Y(n_443)
);

OAI22xp5_ASAP7_75t_L g448 ( 
.A1(n_433),
.A2(n_375),
.B1(n_373),
.B2(n_395),
.Y(n_448)
);

AOI21xp5_ASAP7_75t_L g434 ( 
.A1(n_387),
.A2(n_404),
.B(n_379),
.Y(n_434)
);

NAND2xp5_ASAP7_75t_L g436 ( 
.A(n_428),
.B(n_392),
.Y(n_436)
);

INVx1_ASAP7_75t_L g468 ( 
.A(n_436),
.Y(n_468)
);

INVx1_ASAP7_75t_L g469 ( 
.A(n_437),
.Y(n_469)
);

NAND2xp5_ASAP7_75t_L g438 ( 
.A(n_428),
.B(n_380),
.Y(n_438)
);

INVx1_ASAP7_75t_L g483 ( 
.A(n_438),
.Y(n_483)
);

NAND2xp5_ASAP7_75t_L g439 ( 
.A(n_430),
.B(n_397),
.Y(n_439)
);

NAND2xp5_ASAP7_75t_L g484 ( 
.A(n_439),
.B(n_441),
.Y(n_484)
);

XOR2xp5_ASAP7_75t_L g474 ( 
.A(n_440),
.B(n_406),
.Y(n_474)
);

INVx2_ASAP7_75t_L g441 ( 
.A(n_430),
.Y(n_441)
);

AOI21xp5_ASAP7_75t_L g470 ( 
.A1(n_442),
.A2(n_444),
.B(n_445),
.Y(n_470)
);

OAI21xp5_ASAP7_75t_L g445 ( 
.A1(n_434),
.A2(n_376),
.B(n_385),
.Y(n_445)
);

MAJIxp5_ASAP7_75t_L g446 ( 
.A(n_419),
.B(n_401),
.C(n_382),
.Y(n_446)
);

MAJIxp5_ASAP7_75t_L g463 ( 
.A(n_446),
.B(n_457),
.C(n_461),
.Y(n_463)
);

NOR2xp33_ASAP7_75t_L g447 ( 
.A(n_409),
.B(n_399),
.Y(n_447)
);

CKINVDCx16_ASAP7_75t_R g472 ( 
.A(n_447),
.Y(n_472)
);

AOI22xp5_ASAP7_75t_L g477 ( 
.A1(n_448),
.A2(n_455),
.B1(n_408),
.B2(n_417),
.Y(n_477)
);

INVx1_ASAP7_75t_L g449 ( 
.A(n_414),
.Y(n_449)
);

NOR2xp33_ASAP7_75t_L g464 ( 
.A(n_449),
.B(n_450),
.Y(n_464)
);

NAND2xp5_ASAP7_75t_L g450 ( 
.A(n_431),
.B(n_382),
.Y(n_450)
);

NOR2xp33_ASAP7_75t_L g481 ( 
.A(n_451),
.B(n_452),
.Y(n_481)
);

NAND2xp5_ASAP7_75t_L g452 ( 
.A(n_431),
.B(n_423),
.Y(n_452)
);

NAND2xp5_ASAP7_75t_L g453 ( 
.A(n_413),
.B(n_383),
.Y(n_453)
);

HB1xp67_ASAP7_75t_L g475 ( 
.A(n_453),
.Y(n_475)
);

NAND2xp5_ASAP7_75t_L g454 ( 
.A(n_429),
.B(n_414),
.Y(n_454)
);

XNOR2xp5_ASAP7_75t_L g467 ( 
.A(n_454),
.B(n_459),
.Y(n_467)
);

MAJIxp5_ASAP7_75t_L g457 ( 
.A(n_419),
.B(n_384),
.C(n_388),
.Y(n_457)
);

XNOR2xp5_ASAP7_75t_L g459 ( 
.A(n_418),
.B(n_403),
.Y(n_459)
);

OAI22xp5_ASAP7_75t_SL g473 ( 
.A1(n_460),
.A2(n_412),
.B1(n_433),
.B2(n_411),
.Y(n_473)
);

MAJIxp5_ASAP7_75t_L g461 ( 
.A(n_416),
.B(n_374),
.C(n_420),
.Y(n_461)
);

NAND2x1_ASAP7_75t_L g462 ( 
.A(n_426),
.B(n_405),
.Y(n_462)
);

XOR2x2_ASAP7_75t_L g465 ( 
.A(n_462),
.B(n_426),
.Y(n_465)
);

XNOR2xp5_ASAP7_75t_L g486 ( 
.A(n_465),
.B(n_482),
.Y(n_486)
);

MAJIxp5_ASAP7_75t_L g466 ( 
.A(n_458),
.B(n_424),
.C(n_422),
.Y(n_466)
);

MAJIxp5_ASAP7_75t_L g489 ( 
.A(n_466),
.B(n_471),
.C(n_478),
.Y(n_489)
);

MAJIxp5_ASAP7_75t_L g471 ( 
.A(n_458),
.B(n_425),
.C(n_432),
.Y(n_471)
);

AOI22xp5_ASAP7_75t_SL g485 ( 
.A1(n_473),
.A2(n_455),
.B1(n_441),
.B2(n_460),
.Y(n_485)
);

XOR2xp5_ASAP7_75t_L g491 ( 
.A(n_474),
.B(n_476),
.Y(n_491)
);

XNOR2xp5_ASAP7_75t_SL g476 ( 
.A(n_456),
.B(n_410),
.Y(n_476)
);

OAI22xp5_ASAP7_75t_SL g488 ( 
.A1(n_477),
.A2(n_444),
.B1(n_445),
.B2(n_443),
.Y(n_488)
);

MAJIxp5_ASAP7_75t_L g478 ( 
.A(n_446),
.B(n_410),
.C(n_429),
.Y(n_478)
);

MAJIxp5_ASAP7_75t_L g479 ( 
.A(n_456),
.B(n_435),
.C(n_407),
.Y(n_479)
);

MAJIxp5_ASAP7_75t_L g495 ( 
.A(n_479),
.B(n_438),
.C(n_452),
.Y(n_495)
);

NOR2xp33_ASAP7_75t_SL g480 ( 
.A(n_436),
.B(n_415),
.Y(n_480)
);

NOR2xp33_ASAP7_75t_L g494 ( 
.A(n_480),
.B(n_405),
.Y(n_494)
);

XNOR2xp5_ASAP7_75t_L g482 ( 
.A(n_440),
.B(n_435),
.Y(n_482)
);

OAI22xp5_ASAP7_75t_SL g504 ( 
.A1(n_485),
.A2(n_477),
.B1(n_481),
.B2(n_464),
.Y(n_504)
);

XNOR2xp5_ASAP7_75t_L g487 ( 
.A(n_466),
.B(n_459),
.Y(n_487)
);

NOR2xp33_ASAP7_75t_L g510 ( 
.A(n_487),
.B(n_490),
.Y(n_510)
);

AOI22xp5_ASAP7_75t_L g502 ( 
.A1(n_488),
.A2(n_499),
.B1(n_500),
.B2(n_443),
.Y(n_502)
);

XNOR2xp5_ASAP7_75t_L g490 ( 
.A(n_471),
.B(n_457),
.Y(n_490)
);

INVx1_ASAP7_75t_L g492 ( 
.A(n_484),
.Y(n_492)
);

INVx1_ASAP7_75t_L g503 ( 
.A(n_492),
.Y(n_503)
);

XNOR2xp5_ASAP7_75t_L g493 ( 
.A(n_463),
.B(n_461),
.Y(n_493)
);

XNOR2xp5_ASAP7_75t_L g514 ( 
.A(n_493),
.B(n_495),
.Y(n_514)
);

CKINVDCx20_ASAP7_75t_R g515 ( 
.A(n_494),
.Y(n_515)
);

MAJIxp5_ASAP7_75t_L g496 ( 
.A(n_463),
.B(n_455),
.C(n_450),
.Y(n_496)
);

MAJIxp5_ASAP7_75t_L g511 ( 
.A(n_496),
.B(n_501),
.C(n_482),
.Y(n_511)
);

BUFx24_ASAP7_75t_SL g497 ( 
.A(n_469),
.Y(n_497)
);

OAI21xp5_ASAP7_75t_SL g508 ( 
.A1(n_497),
.A2(n_451),
.B(n_475),
.Y(n_508)
);

XOR2xp5_ASAP7_75t_L g498 ( 
.A(n_474),
.B(n_442),
.Y(n_498)
);

XOR2xp5_ASAP7_75t_L g505 ( 
.A(n_498),
.B(n_470),
.Y(n_505)
);

INVx1_ASAP7_75t_L g499 ( 
.A(n_468),
.Y(n_499)
);

INVx1_ASAP7_75t_L g500 ( 
.A(n_483),
.Y(n_500)
);

XNOR2xp5_ASAP7_75t_L g501 ( 
.A(n_467),
.B(n_454),
.Y(n_501)
);

CKINVDCx20_ASAP7_75t_R g517 ( 
.A(n_502),
.Y(n_517)
);

AOI22xp5_ASAP7_75t_SL g516 ( 
.A1(n_504),
.A2(n_462),
.B1(n_472),
.B2(n_498),
.Y(n_516)
);

XOR2xp5_ASAP7_75t_L g525 ( 
.A(n_505),
.B(n_506),
.Y(n_525)
);

MAJx2_ASAP7_75t_L g506 ( 
.A(n_496),
.B(n_478),
.C(n_479),
.Y(n_506)
);

XOR2xp5_ASAP7_75t_L g507 ( 
.A(n_491),
.B(n_467),
.Y(n_507)
);

MAJIxp5_ASAP7_75t_L g524 ( 
.A(n_507),
.B(n_512),
.C(n_513),
.Y(n_524)
);

NOR2xp33_ASAP7_75t_L g520 ( 
.A(n_508),
.B(n_511),
.Y(n_520)
);

OAI22xp5_ASAP7_75t_SL g509 ( 
.A1(n_485),
.A2(n_449),
.B1(n_439),
.B2(n_462),
.Y(n_509)
);

AOI22xp5_ASAP7_75t_L g518 ( 
.A1(n_509),
.A2(n_486),
.B1(n_427),
.B2(n_415),
.Y(n_518)
);

MAJIxp5_ASAP7_75t_L g512 ( 
.A(n_489),
.B(n_473),
.C(n_476),
.Y(n_512)
);

XOR2xp5_ASAP7_75t_L g513 ( 
.A(n_491),
.B(n_465),
.Y(n_513)
);

NAND2xp5_ASAP7_75t_L g529 ( 
.A(n_516),
.B(n_519),
.Y(n_529)
);

NAND2xp5_ASAP7_75t_SL g527 ( 
.A(n_518),
.B(n_523),
.Y(n_527)
);

OAI22xp5_ASAP7_75t_L g519 ( 
.A1(n_515),
.A2(n_495),
.B1(n_453),
.B2(n_489),
.Y(n_519)
);

NOR2xp33_ASAP7_75t_L g521 ( 
.A(n_514),
.B(n_427),
.Y(n_521)
);

NAND2xp5_ASAP7_75t_L g530 ( 
.A(n_521),
.B(n_507),
.Y(n_530)
);

OAI21xp5_ASAP7_75t_SL g522 ( 
.A1(n_510),
.A2(n_512),
.B(n_511),
.Y(n_522)
);

NAND2xp5_ASAP7_75t_SL g528 ( 
.A(n_522),
.B(n_514),
.Y(n_528)
);

AOI21xp5_ASAP7_75t_L g523 ( 
.A1(n_504),
.A2(n_509),
.B(n_502),
.Y(n_523)
);

BUFx6f_ASAP7_75t_L g526 ( 
.A(n_520),
.Y(n_526)
);

INVx1_ASAP7_75t_L g532 ( 
.A(n_526),
.Y(n_532)
);

INVx1_ASAP7_75t_L g533 ( 
.A(n_528),
.Y(n_533)
);

INVx1_ASAP7_75t_L g535 ( 
.A(n_530),
.Y(n_535)
);

NAND2xp5_ASAP7_75t_L g531 ( 
.A(n_517),
.B(n_503),
.Y(n_531)
);

NOR2xp33_ASAP7_75t_L g534 ( 
.A(n_531),
.B(n_518),
.Y(n_534)
);

INVx1_ASAP7_75t_L g537 ( 
.A(n_534),
.Y(n_537)
);

XOR2xp5_ASAP7_75t_L g536 ( 
.A(n_532),
.B(n_524),
.Y(n_536)
);

INVx1_ASAP7_75t_L g539 ( 
.A(n_536),
.Y(n_539)
);

MAJIxp5_ASAP7_75t_L g538 ( 
.A(n_537),
.B(n_533),
.C(n_535),
.Y(n_538)
);

A2O1A1O1Ixp25_ASAP7_75t_L g540 ( 
.A1(n_538),
.A2(n_529),
.B(n_527),
.C(n_525),
.D(n_524),
.Y(n_540)
);

NAND2xp5_ASAP7_75t_L g541 ( 
.A(n_540),
.B(n_525),
.Y(n_541)
);

OAI21xp5_ASAP7_75t_L g542 ( 
.A1(n_541),
.A2(n_539),
.B(n_523),
.Y(n_542)
);

MAJIxp5_ASAP7_75t_L g543 ( 
.A(n_542),
.B(n_527),
.C(n_506),
.Y(n_543)
);

FAx1_ASAP7_75t_SL g544 ( 
.A(n_543),
.B(n_505),
.CI(n_513),
.CON(n_544),
.SN(n_544)
);

XNOR2xp5_ASAP7_75t_L g545 ( 
.A(n_544),
.B(n_516),
.Y(n_545)
);


endmodule