module fake_ariane_1718_n_1702 (n_83, n_8, n_56, n_60, n_64, n_119, n_124, n_90, n_38, n_47, n_110, n_153, n_18, n_86, n_75, n_89, n_67, n_149, n_34, n_69, n_95, n_92, n_143, n_150, n_98, n_74, n_113, n_114, n_33, n_19, n_40, n_152, n_120, n_106, n_12, n_53, n_111, n_21, n_115, n_133, n_66, n_71, n_24, n_7, n_109, n_96, n_49, n_20, n_100, n_17, n_50, n_132, n_62, n_147, n_51, n_76, n_103, n_79, n_26, n_3, n_46, n_0, n_84, n_36, n_91, n_107, n_72, n_105, n_128, n_44, n_30, n_82, n_31, n_42, n_57, n_131, n_70, n_10, n_117, n_139, n_85, n_130, n_144, n_6, n_48, n_94, n_101, n_4, n_134, n_2, n_32, n_37, n_58, n_65, n_123, n_9, n_138, n_112, n_45, n_11, n_129, n_126, n_137, n_122, n_148, n_52, n_135, n_73, n_77, n_15, n_118, n_93, n_121, n_23, n_61, n_108, n_102, n_125, n_22, n_43, n_1, n_81, n_87, n_13, n_27, n_29, n_41, n_140, n_55, n_151, n_136, n_28, n_80, n_146, n_97, n_154, n_142, n_14, n_88, n_141, n_68, n_116, n_104, n_145, n_78, n_39, n_59, n_63, n_99, n_16, n_5, n_127, n_35, n_54, n_25, n_1702);

input n_83;
input n_8;
input n_56;
input n_60;
input n_64;
input n_119;
input n_124;
input n_90;
input n_38;
input n_47;
input n_110;
input n_153;
input n_18;
input n_86;
input n_75;
input n_89;
input n_67;
input n_149;
input n_34;
input n_69;
input n_95;
input n_92;
input n_143;
input n_150;
input n_98;
input n_74;
input n_113;
input n_114;
input n_33;
input n_19;
input n_40;
input n_152;
input n_120;
input n_106;
input n_12;
input n_53;
input n_111;
input n_21;
input n_115;
input n_133;
input n_66;
input n_71;
input n_24;
input n_7;
input n_109;
input n_96;
input n_49;
input n_20;
input n_100;
input n_17;
input n_50;
input n_132;
input n_62;
input n_147;
input n_51;
input n_76;
input n_103;
input n_79;
input n_26;
input n_3;
input n_46;
input n_0;
input n_84;
input n_36;
input n_91;
input n_107;
input n_72;
input n_105;
input n_128;
input n_44;
input n_30;
input n_82;
input n_31;
input n_42;
input n_57;
input n_131;
input n_70;
input n_10;
input n_117;
input n_139;
input n_85;
input n_130;
input n_144;
input n_6;
input n_48;
input n_94;
input n_101;
input n_4;
input n_134;
input n_2;
input n_32;
input n_37;
input n_58;
input n_65;
input n_123;
input n_9;
input n_138;
input n_112;
input n_45;
input n_11;
input n_129;
input n_126;
input n_137;
input n_122;
input n_148;
input n_52;
input n_135;
input n_73;
input n_77;
input n_15;
input n_118;
input n_93;
input n_121;
input n_23;
input n_61;
input n_108;
input n_102;
input n_125;
input n_22;
input n_43;
input n_1;
input n_81;
input n_87;
input n_13;
input n_27;
input n_29;
input n_41;
input n_140;
input n_55;
input n_151;
input n_136;
input n_28;
input n_80;
input n_146;
input n_97;
input n_154;
input n_142;
input n_14;
input n_88;
input n_141;
input n_68;
input n_116;
input n_104;
input n_145;
input n_78;
input n_39;
input n_59;
input n_63;
input n_99;
input n_16;
input n_5;
input n_127;
input n_35;
input n_54;
input n_25;

output n_1702;

wire n_913;
wire n_1681;
wire n_1507;
wire n_1486;
wire n_589;
wire n_1174;
wire n_1469;
wire n_691;
wire n_1353;
wire n_1355;
wire n_423;
wire n_1383;
wire n_603;
wire n_373;
wire n_1250;
wire n_1169;
wire n_789;
wire n_850;
wire n_610;
wire n_245;
wire n_319;
wire n_1436;
wire n_690;
wire n_416;
wire n_1109;
wire n_1430;
wire n_525;
wire n_187;
wire n_1463;
wire n_1238;
wire n_1515;
wire n_817;
wire n_924;
wire n_781;
wire n_1566;
wire n_189;
wire n_717;
wire n_952;
wire n_864;
wire n_1096;
wire n_1379;
wire n_524;
wire n_1214;
wire n_634;
wire n_1246;
wire n_1138;
wire n_214;
wire n_764;
wire n_1503;
wire n_462;
wire n_1196;
wire n_1181;
wire n_410;
wire n_1187;
wire n_1131;
wire n_1225;
wire n_737;
wire n_1298;
wire n_1366;
wire n_232;
wire n_568;
wire n_1088;
wire n_1424;
wire n_766;
wire n_1457;
wire n_377;
wire n_1682;
wire n_520;
wire n_870;
wire n_1453;
wire n_279;
wire n_945;
wire n_958;
wire n_813;
wire n_419;
wire n_270;
wire n_338;
wire n_995;
wire n_285;
wire n_1184;
wire n_202;
wire n_1535;
wire n_500;
wire n_665;
wire n_754;
wire n_903;
wire n_871;
wire n_1073;
wire n_239;
wire n_402;
wire n_1277;
wire n_829;
wire n_1062;
wire n_339;
wire n_738;
wire n_1690;
wire n_672;
wire n_740;
wire n_1283;
wire n_167;
wire n_1018;
wire n_259;
wire n_953;
wire n_1364;
wire n_1224;
wire n_1425;
wire n_625;
wire n_557;
wire n_1107;
wire n_1688;
wire n_989;
wire n_242;
wire n_645;
wire n_331;
wire n_559;
wire n_267;
wire n_495;
wire n_350;
wire n_381;
wire n_795;
wire n_721;
wire n_1084;
wire n_1276;
wire n_200;
wire n_1428;
wire n_1284;
wire n_1241;
wire n_821;
wire n_561;
wire n_770;
wire n_1514;
wire n_1528;
wire n_507;
wire n_486;
wire n_901;
wire n_569;
wire n_1145;
wire n_971;
wire n_787;
wire n_1650;
wire n_1519;
wire n_1195;
wire n_1522;
wire n_518;
wire n_1207;
wire n_222;
wire n_786;
wire n_1404;
wire n_868;
wire n_1542;
wire n_1314;
wire n_1512;
wire n_1539;
wire n_884;
wire n_1415;
wire n_1034;
wire n_1652;
wire n_1676;
wire n_1085;
wire n_277;
wire n_1636;
wire n_432;
wire n_293;
wire n_823;
wire n_620;
wire n_1074;
wire n_859;
wire n_587;
wire n_693;
wire n_863;
wire n_303;
wire n_1254;
wire n_929;
wire n_206;
wire n_352;
wire n_899;
wire n_611;
wire n_1295;
wire n_365;
wire n_238;
wire n_1013;
wire n_1495;
wire n_1637;
wire n_334;
wire n_192;
wire n_661;
wire n_300;
wire n_533;
wire n_438;
wire n_1654;
wire n_1560;
wire n_1548;
wire n_440;
wire n_273;
wire n_1396;
wire n_1230;
wire n_612;
wire n_333;
wire n_376;
wire n_512;
wire n_1597;
wire n_1544;
wire n_579;
wire n_844;
wire n_1012;
wire n_1267;
wire n_1354;
wire n_1213;
wire n_237;
wire n_780;
wire n_1021;
wire n_1443;
wire n_491;
wire n_1465;
wire n_1595;
wire n_1142;
wire n_1140;
wire n_705;
wire n_570;
wire n_260;
wire n_942;
wire n_1437;
wire n_1378;
wire n_461;
wire n_1121;
wire n_1416;
wire n_490;
wire n_209;
wire n_1461;
wire n_1391;
wire n_225;
wire n_1599;
wire n_1006;
wire n_575;
wire n_546;
wire n_503;
wire n_1112;
wire n_700;
wire n_1159;
wire n_772;
wire n_1216;
wire n_1245;
wire n_1669;
wire n_1675;
wire n_676;
wire n_1594;
wire n_680;
wire n_287;
wire n_302;
wire n_380;
wire n_1585;
wire n_1432;
wire n_249;
wire n_1108;
wire n_355;
wire n_212;
wire n_444;
wire n_851;
wire n_1590;
wire n_1351;
wire n_1274;
wire n_257;
wire n_652;
wire n_475;
wire n_947;
wire n_930;
wire n_1260;
wire n_1179;
wire n_468;
wire n_182;
wire n_696;
wire n_1442;
wire n_482;
wire n_798;
wire n_577;
wire n_407;
wire n_1691;
wire n_916;
wire n_1386;
wire n_912;
wire n_460;
wire n_1555;
wire n_366;
wire n_762;
wire n_1253;
wire n_1468;
wire n_1661;
wire n_555;
wire n_804;
wire n_1656;
wire n_1382;
wire n_992;
wire n_966;
wire n_955;
wire n_1182;
wire n_794;
wire n_1692;
wire n_1562;
wire n_514;
wire n_418;
wire n_1376;
wire n_513;
wire n_288;
wire n_179;
wire n_1292;
wire n_1178;
wire n_1435;
wire n_1026;
wire n_1506;
wire n_1610;
wire n_306;
wire n_203;
wire n_436;
wire n_324;
wire n_669;
wire n_931;
wire n_1491;
wire n_619;
wire n_337;
wire n_437;
wire n_274;
wire n_1083;
wire n_967;
wire n_1418;
wire n_746;
wire n_1357;
wire n_292;
wire n_1079;
wire n_1389;
wire n_615;
wire n_1139;
wire n_517;
wire n_1312;
wire n_824;
wire n_428;
wire n_159;
wire n_892;
wire n_959;
wire n_1399;
wire n_1101;
wire n_1567;
wire n_1343;
wire n_563;
wire n_990;
wire n_1623;
wire n_867;
wire n_1226;
wire n_944;
wire n_749;
wire n_815;
wire n_542;
wire n_1340;
wire n_470;
wire n_1240;
wire n_1087;
wire n_632;
wire n_477;
wire n_650;
wire n_425;
wire n_1433;
wire n_1155;
wire n_1071;
wire n_712;
wire n_976;
wire n_909;
wire n_1392;
wire n_767;
wire n_1680;
wire n_964;
wire n_1627;
wire n_382;
wire n_489;
wire n_251;
wire n_974;
wire n_506;
wire n_799;
wire n_1147;
wire n_397;
wire n_471;
wire n_351;
wire n_965;
wire n_155;
wire n_934;
wire n_1447;
wire n_1220;
wire n_356;
wire n_698;
wire n_1674;
wire n_307;
wire n_1209;
wire n_1020;
wire n_1563;
wire n_646;
wire n_1633;
wire n_404;
wire n_172;
wire n_1058;
wire n_347;
wire n_1042;
wire n_183;
wire n_1234;
wire n_479;
wire n_1578;
wire n_1455;
wire n_299;
wire n_836;
wire n_1279;
wire n_564;
wire n_205;
wire n_1029;
wire n_1247;
wire n_760;
wire n_522;
wire n_1568;
wire n_1483;
wire n_1363;
wire n_367;
wire n_1111;
wire n_970;
wire n_1689;
wire n_713;
wire n_1255;
wire n_1646;
wire n_598;
wire n_345;
wire n_1237;
wire n_927;
wire n_261;
wire n_1095;
wire n_370;
wire n_706;
wire n_286;
wire n_1401;
wire n_1419;
wire n_1531;
wire n_776;
wire n_424;
wire n_1651;
wire n_1387;
wire n_466;
wire n_1263;
wire n_346;
wire n_348;
wire n_552;
wire n_670;
wire n_379;
wire n_162;
wire n_264;
wire n_441;
wire n_1032;
wire n_1217;
wire n_1496;
wire n_637;
wire n_1592;
wire n_327;
wire n_1259;
wire n_1177;
wire n_1231;
wire n_980;
wire n_1618;
wire n_905;
wire n_207;
wire n_720;
wire n_926;
wire n_194;
wire n_1163;
wire n_186;
wire n_1384;
wire n_1501;
wire n_1173;
wire n_1068;
wire n_1198;
wire n_1570;
wire n_487;
wire n_1518;
wire n_1456;
wire n_1648;
wire n_1413;
wire n_855;
wire n_158;
wire n_808;
wire n_1365;
wire n_553;
wire n_1439;
wire n_814;
wire n_578;
wire n_1665;
wire n_1287;
wire n_405;
wire n_1611;
wire n_320;
wire n_1414;
wire n_1134;
wire n_1484;
wire n_647;
wire n_1423;
wire n_481;
wire n_600;
wire n_1053;
wire n_1609;
wire n_529;
wire n_502;
wire n_218;
wire n_1467;
wire n_247;
wire n_1304;
wire n_1608;
wire n_1105;
wire n_547;
wire n_439;
wire n_604;
wire n_677;
wire n_478;
wire n_703;
wire n_1349;
wire n_1061;
wire n_326;
wire n_681;
wire n_227;
wire n_874;
wire n_1278;
wire n_707;
wire n_983;
wire n_590;
wire n_727;
wire n_699;
wire n_301;
wire n_545;
wire n_1015;
wire n_1377;
wire n_1162;
wire n_536;
wire n_1614;
wire n_325;
wire n_1602;
wire n_688;
wire n_636;
wire n_427;
wire n_1098;
wire n_1490;
wire n_442;
wire n_777;
wire n_1553;
wire n_1080;
wire n_920;
wire n_1086;
wire n_1092;
wire n_986;
wire n_1104;
wire n_729;
wire n_887;
wire n_1122;
wire n_1205;
wire n_1408;
wire n_163;
wire n_1693;
wire n_1132;
wire n_390;
wire n_1156;
wire n_501;
wire n_314;
wire n_1120;
wire n_1202;
wire n_627;
wire n_1188;
wire n_1498;
wire n_1371;
wire n_233;
wire n_957;
wire n_388;
wire n_1402;
wire n_1242;
wire n_1607;
wire n_1489;
wire n_1218;
wire n_221;
wire n_321;
wire n_1586;
wire n_861;
wire n_1543;
wire n_1431;
wire n_877;
wire n_1119;
wire n_1666;
wire n_1500;
wire n_616;
wire n_1055;
wire n_1395;
wire n_1346;
wire n_1189;
wire n_1089;
wire n_281;
wire n_262;
wire n_1502;
wire n_1523;
wire n_1478;
wire n_735;
wire n_297;
wire n_1005;
wire n_527;
wire n_1294;
wire n_1667;
wire n_845;
wire n_888;
wire n_1649;
wire n_1677;
wire n_1297;
wire n_178;
wire n_551;
wire n_417;
wire n_343;
wire n_1222;
wire n_582;
wire n_755;
wire n_1097;
wire n_1219;
wire n_710;
wire n_534;
wire n_1460;
wire n_1239;
wire n_278;
wire n_560;
wire n_890;
wire n_842;
wire n_451;
wire n_745;
wire n_1572;
wire n_742;
wire n_1081;
wire n_1373;
wire n_1388;
wire n_1266;
wire n_1540;
wire n_769;
wire n_1372;
wire n_476;
wire n_832;
wire n_535;
wire n_744;
wire n_982;
wire n_915;
wire n_215;
wire n_1075;
wire n_454;
wire n_298;
wire n_1331;
wire n_1529;
wire n_1227;
wire n_655;
wire n_403;
wire n_1007;
wire n_1580;
wire n_1319;
wire n_657;
wire n_837;
wire n_812;
wire n_606;
wire n_951;
wire n_862;
wire n_1700;
wire n_659;
wire n_1332;
wire n_509;
wire n_666;
wire n_430;
wire n_1206;
wire n_722;
wire n_1508;
wire n_1532;
wire n_1171;
wire n_1030;
wire n_785;
wire n_1309;
wire n_999;
wire n_1338;
wire n_1342;
wire n_456;
wire n_852;
wire n_1394;
wire n_704;
wire n_1060;
wire n_1044;
wire n_521;
wire n_873;
wire n_1301;
wire n_1243;
wire n_1400;
wire n_342;
wire n_1466;
wire n_1513;
wire n_1527;
wire n_358;
wire n_608;
wire n_1538;
wire n_1037;
wire n_1329;
wire n_317;
wire n_1545;
wire n_1257;
wire n_1480;
wire n_1668;
wire n_1605;
wire n_1078;
wire n_266;
wire n_157;
wire n_1161;
wire n_811;
wire n_624;
wire n_791;
wire n_876;
wire n_618;
wire n_1191;
wire n_736;
wire n_1025;
wire n_1215;
wire n_241;
wire n_1449;
wire n_687;
wire n_797;
wire n_480;
wire n_1327;
wire n_1475;
wire n_211;
wire n_642;
wire n_408;
wire n_1406;
wire n_595;
wire n_1405;
wire n_602;
wire n_592;
wire n_1499;
wire n_854;
wire n_1318;
wire n_393;
wire n_1632;
wire n_474;
wire n_805;
wire n_295;
wire n_1658;
wire n_190;
wire n_1072;
wire n_695;
wire n_1526;
wire n_1305;
wire n_180;
wire n_730;
wire n_386;
wire n_1596;
wire n_1281;
wire n_516;
wire n_1137;
wire n_1258;
wire n_197;
wire n_640;
wire n_463;
wire n_1476;
wire n_1524;
wire n_943;
wire n_1118;
wire n_678;
wire n_651;
wire n_1293;
wire n_961;
wire n_469;
wire n_1046;
wire n_726;
wire n_1123;
wire n_1657;
wire n_878;
wire n_771;
wire n_1321;
wire n_752;
wire n_1488;
wire n_985;
wire n_421;
wire n_1330;
wire n_906;
wire n_1180;
wire n_1697;
wire n_283;
wire n_806;
wire n_1350;
wire n_1556;
wire n_649;
wire n_1561;
wire n_374;
wire n_1352;
wire n_643;
wire n_1492;
wire n_226;
wire n_1441;
wire n_682;
wire n_1616;
wire n_819;
wire n_586;
wire n_1324;
wire n_1429;
wire n_686;
wire n_605;
wire n_1154;
wire n_584;
wire n_1557;
wire n_1130;
wire n_1450;
wire n_349;
wire n_756;
wire n_1016;
wire n_1149;
wire n_1505;
wire n_979;
wire n_1642;
wire n_897;
wire n_949;
wire n_1493;
wire n_515;
wire n_807;
wire n_891;
wire n_885;
wire n_1659;
wire n_198;
wire n_1208;
wire n_396;
wire n_802;
wire n_1151;
wire n_554;
wire n_960;
wire n_1256;
wire n_714;
wire n_790;
wire n_354;
wire n_725;
wire n_1577;
wire n_1448;
wire n_1009;
wire n_230;
wire n_1133;
wire n_883;
wire n_473;
wire n_801;
wire n_1286;
wire n_818;
wire n_1685;
wire n_779;
wire n_594;
wire n_1397;
wire n_1052;
wire n_272;
wire n_1333;
wire n_1306;
wire n_833;
wire n_1426;
wire n_879;
wire n_1117;
wire n_422;
wire n_1269;
wire n_1303;
wire n_1547;
wire n_1438;
wire n_1541;
wire n_597;
wire n_1047;
wire n_1472;
wire n_1593;
wire n_1050;
wire n_566;
wire n_169;
wire n_1201;
wire n_1288;
wire n_173;
wire n_858;
wire n_1185;
wire n_335;
wire n_1035;
wire n_1143;
wire n_344;
wire n_426;
wire n_433;
wire n_398;
wire n_210;
wire n_1090;
wire n_1367;
wire n_253;
wire n_166;
wire n_928;
wire n_1153;
wire n_271;
wire n_465;
wire n_825;
wire n_1103;
wire n_732;
wire n_1565;
wire n_1192;
wire n_224;
wire n_894;
wire n_1380;
wire n_1624;
wire n_420;
wire n_1291;
wire n_562;
wire n_748;
wire n_510;
wire n_1045;
wire n_256;
wire n_1160;
wire n_1023;
wire n_988;
wire n_330;
wire n_914;
wire n_400;
wire n_689;
wire n_1116;
wire n_282;
wire n_328;
wire n_368;
wire n_467;
wire n_1511;
wire n_1422;
wire n_644;
wire n_1197;
wire n_276;
wire n_497;
wire n_1165;
wire n_1641;
wire n_168;
wire n_538;
wire n_1517;
wire n_576;
wire n_843;
wire n_511;
wire n_455;
wire n_429;
wire n_588;
wire n_638;
wire n_1307;
wire n_1128;
wire n_1671;
wire n_1417;
wire n_1048;
wire n_775;
wire n_667;
wire n_1049;
wire n_869;
wire n_846;
wire n_1398;
wire n_1356;
wire n_1341;
wire n_1504;
wire n_1440;
wire n_1370;
wire n_1603;
wire n_305;
wire n_312;
wire n_728;
wire n_413;
wire n_715;
wire n_889;
wire n_1066;
wire n_1549;
wire n_935;
wire n_685;
wire n_911;
wire n_361;
wire n_623;
wire n_1403;
wire n_1065;
wire n_453;
wire n_1534;
wire n_810;
wire n_1290;
wire n_181;
wire n_617;
wire n_543;
wire n_1362;
wire n_1559;
wire n_236;
wire n_683;
wire n_601;
wire n_565;
wire n_628;
wire n_1300;
wire n_743;
wire n_1194;
wire n_1647;
wire n_1546;
wire n_1420;
wire n_907;
wire n_1454;
wire n_660;
wire n_464;
wire n_962;
wire n_941;
wire n_1210;
wire n_847;
wire n_747;
wire n_1622;
wire n_1135;
wire n_918;
wire n_639;
wire n_452;
wire n_673;
wire n_1038;
wire n_414;
wire n_571;
wire n_1521;
wire n_1694;
wire n_284;
wire n_593;
wire n_1695;
wire n_1164;
wire n_609;
wire n_1193;
wire n_1345;
wire n_613;
wire n_1022;
wire n_1336;
wire n_1033;
wire n_409;
wire n_171;
wire n_519;
wire n_384;
wire n_1166;
wire n_1056;
wire n_526;
wire n_1040;
wire n_674;
wire n_1158;
wire n_316;
wire n_1444;
wire n_820;
wire n_872;
wire n_1653;
wire n_254;
wire n_1157;
wire n_1584;
wire n_234;
wire n_848;
wire n_1664;
wire n_280;
wire n_629;
wire n_161;
wire n_532;
wire n_763;
wire n_540;
wire n_216;
wire n_692;
wire n_984;
wire n_1687;
wire n_223;
wire n_1552;
wire n_750;
wire n_834;
wire n_1612;
wire n_800;
wire n_1606;
wire n_395;
wire n_621;
wire n_1587;
wire n_213;
wire n_1014;
wire n_724;
wire n_1427;
wire n_1481;
wire n_493;
wire n_1311;
wire n_1589;
wire n_1100;
wire n_585;
wire n_875;
wire n_1617;
wire n_827;
wire n_697;
wire n_622;
wire n_1626;
wire n_1335;
wire n_296;
wire n_880;
wire n_793;
wire n_1175;
wire n_751;
wire n_1027;
wire n_1070;
wire n_1621;
wire n_739;
wire n_1485;
wire n_1028;
wire n_1221;
wire n_530;
wire n_792;
wire n_1262;
wire n_580;
wire n_1579;
wire n_494;
wire n_434;
wire n_975;
wire n_229;
wire n_394;
wire n_923;
wire n_1645;
wire n_1124;
wire n_1381;
wire n_1494;
wire n_932;
wire n_1183;
wire n_1326;
wire n_981;
wire n_1110;
wire n_243;
wire n_1407;
wire n_185;
wire n_1204;
wire n_1554;
wire n_994;
wire n_1360;
wire n_973;
wire n_268;
wire n_972;
wire n_164;
wire n_184;
wire n_856;
wire n_1248;
wire n_1176;
wire n_1564;
wire n_1054;
wire n_508;
wire n_1679;
wire n_353;
wire n_1678;
wire n_1482;
wire n_1361;
wire n_1601;
wire n_1057;
wire n_191;
wire n_978;
wire n_1011;
wire n_1520;
wire n_1509;
wire n_828;
wire n_322;
wire n_1411;
wire n_1359;
wire n_558;
wire n_653;
wire n_1445;
wire n_1317;
wire n_783;
wire n_556;
wire n_1127;
wire n_170;
wire n_1536;
wire n_1471;
wire n_160;
wire n_1008;
wire n_332;
wire n_581;
wire n_294;
wire n_1024;
wire n_830;
wire n_176;
wire n_987;
wire n_936;
wire n_1620;
wire n_1385;
wire n_1525;
wire n_541;
wire n_499;
wire n_788;
wire n_908;
wire n_1036;
wire n_341;
wire n_1270;
wire n_1167;
wire n_1272;
wire n_549;
wire n_591;
wire n_969;
wire n_919;
wire n_1663;
wire n_1625;
wire n_318;
wire n_1458;
wire n_244;
wire n_679;
wire n_1630;
wire n_220;
wire n_663;
wire n_443;
wire n_1412;
wire n_1550;
wire n_528;
wire n_1358;
wire n_1200;
wire n_387;
wire n_406;
wire n_826;
wire n_391;
wire n_940;
wire n_1537;
wire n_1077;
wire n_607;
wire n_956;
wire n_445;
wire n_765;
wire n_1268;
wire n_385;
wire n_917;
wire n_1271;
wire n_372;
wire n_1530;
wire n_631;
wire n_399;
wire n_1170;
wire n_1261;
wire n_702;
wire n_898;
wire n_857;
wire n_363;
wire n_1067;
wire n_968;
wire n_1235;
wire n_1323;
wire n_1462;
wire n_1064;
wire n_633;
wire n_900;
wire n_1446;
wire n_1282;
wire n_1701;
wire n_1093;
wire n_1551;
wire n_1285;
wire n_193;
wire n_733;
wire n_761;
wire n_731;
wire n_336;
wire n_315;
wire n_311;
wire n_1452;
wire n_1573;
wire n_668;
wire n_758;
wire n_1106;
wire n_648;
wire n_784;
wire n_269;
wire n_816;
wire n_1322;
wire n_1473;
wire n_835;
wire n_446;
wire n_1076;
wire n_1348;
wire n_753;
wire n_701;
wire n_1003;
wire n_1125;
wire n_309;
wire n_1344;
wire n_1390;
wire n_401;
wire n_485;
wire n_504;
wire n_483;
wire n_435;
wire n_1141;
wire n_1629;
wire n_291;
wire n_1640;
wire n_822;
wire n_1094;
wire n_840;
wire n_1459;
wire n_1510;
wire n_1099;
wire n_839;
wire n_759;
wire n_567;
wire n_240;
wire n_369;
wire n_1575;
wire n_1172;
wire n_614;
wire n_1212;
wire n_831;
wire n_778;
wire n_1619;
wire n_188;
wire n_323;
wire n_550;
wire n_1315;
wire n_1660;
wire n_997;
wire n_635;
wire n_694;
wire n_1643;
wire n_1320;
wire n_1113;
wire n_248;
wire n_1152;
wire n_921;
wire n_1615;
wire n_1236;
wire n_228;
wire n_1265;
wire n_1576;
wire n_1470;
wire n_671;
wire n_1533;
wire n_1409;
wire n_1148;
wire n_1588;
wire n_1684;
wire n_1673;
wire n_1334;
wire n_654;
wire n_1275;
wire n_488;
wire n_904;
wire n_505;
wire n_1696;
wire n_498;
wire n_1059;
wire n_684;
wire n_1039;
wire n_539;
wire n_1150;
wire n_977;
wire n_449;
wire n_392;
wire n_1628;
wire n_1289;
wire n_1497;
wire n_459;
wire n_1136;
wire n_458;
wire n_1190;
wire n_1600;
wire n_1144;
wire n_383;
wire n_838;
wire n_1558;
wire n_1316;
wire n_175;
wire n_950;
wire n_1017;
wire n_711;
wire n_734;
wire n_723;
wire n_1393;
wire n_658;
wire n_630;
wire n_1369;
wire n_362;
wire n_310;
wire n_709;
wire n_809;
wire n_1686;
wire n_235;
wire n_881;
wire n_1019;
wire n_1477;
wire n_662;
wire n_641;
wire n_910;
wire n_290;
wire n_741;
wire n_939;
wire n_1410;
wire n_371;
wire n_199;
wire n_217;
wire n_1114;
wire n_1325;
wire n_708;
wire n_308;
wire n_1223;
wire n_201;
wire n_572;
wire n_1199;
wire n_865;
wire n_1273;
wire n_1041;
wire n_993;
wire n_948;
wire n_922;
wire n_1004;
wire n_448;
wire n_1347;
wire n_860;
wire n_1043;
wire n_255;
wire n_450;
wire n_896;
wire n_1479;
wire n_1613;
wire n_902;
wire n_1031;
wire n_1638;
wire n_853;
wire n_716;
wire n_1571;
wire n_1698;
wire n_196;
wire n_1337;
wire n_774;
wire n_933;
wire n_596;
wire n_954;
wire n_1168;
wire n_219;
wire n_1310;
wire n_231;
wire n_656;
wire n_492;
wire n_574;
wire n_252;
wire n_664;
wire n_1591;
wire n_1229;
wire n_1683;
wire n_415;
wire n_1280;
wire n_544;
wire n_1516;
wire n_1186;
wire n_599;
wire n_768;
wire n_1091;
wire n_537;
wire n_1063;
wire n_991;
wire n_389;
wire n_1670;
wire n_1126;
wire n_195;
wire n_938;
wire n_1328;
wire n_895;
wire n_304;
wire n_1639;
wire n_583;
wire n_1302;
wire n_1000;
wire n_313;
wire n_626;
wire n_378;
wire n_1581;
wire n_946;
wire n_757;
wire n_375;
wire n_1655;
wire n_1146;
wire n_1634;
wire n_1203;
wire n_998;
wire n_1699;
wire n_1598;
wire n_472;
wire n_937;
wire n_1474;
wire n_265;
wire n_1583;
wire n_1604;
wire n_208;
wire n_1631;
wire n_156;
wire n_174;
wire n_275;
wire n_1375;
wire n_204;
wire n_1232;
wire n_996;
wire n_1211;
wire n_1368;
wire n_963;
wire n_1264;
wire n_1082;
wire n_496;
wire n_866;
wire n_246;
wire n_925;
wire n_1313;
wire n_1001;
wire n_1115;
wire n_1339;
wire n_1002;
wire n_1644;
wire n_1051;
wire n_719;
wire n_263;
wire n_1102;
wire n_360;
wire n_1129;
wire n_1252;
wire n_250;
wire n_1464;
wire n_1296;
wire n_773;
wire n_165;
wire n_1010;
wire n_882;
wire n_1249;
wire n_803;
wire n_329;
wire n_718;
wire n_1434;
wire n_340;
wire n_1569;
wire n_548;
wire n_289;
wire n_523;
wire n_1662;
wire n_457;
wire n_1299;
wire n_177;
wire n_782;
wire n_364;
wire n_258;
wire n_431;
wire n_1228;
wire n_1244;
wire n_411;
wire n_484;
wire n_849;
wire n_357;
wire n_412;
wire n_1251;
wire n_447;
wire n_1421;
wire n_1233;
wire n_1574;
wire n_1672;
wire n_1635;
wire n_893;
wire n_1582;
wire n_841;
wire n_886;
wire n_1069;
wire n_359;
wire n_1308;
wire n_573;
wire n_796;
wire n_531;
wire n_1374;
wire n_1451;
wire n_1487;
wire n_675;

BUFx6f_ASAP7_75t_L g155 ( 
.A(n_10),
.Y(n_155)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_55),
.Y(n_156)
);

CKINVDCx5p33_ASAP7_75t_R g157 ( 
.A(n_37),
.Y(n_157)
);

CKINVDCx14_ASAP7_75t_R g158 ( 
.A(n_78),
.Y(n_158)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_148),
.Y(n_159)
);

CKINVDCx5p33_ASAP7_75t_R g160 ( 
.A(n_64),
.Y(n_160)
);

BUFx6f_ASAP7_75t_L g161 ( 
.A(n_59),
.Y(n_161)
);

CKINVDCx20_ASAP7_75t_R g162 ( 
.A(n_112),
.Y(n_162)
);

CKINVDCx20_ASAP7_75t_R g163 ( 
.A(n_45),
.Y(n_163)
);

CKINVDCx5p33_ASAP7_75t_R g164 ( 
.A(n_66),
.Y(n_164)
);

CKINVDCx5p33_ASAP7_75t_R g165 ( 
.A(n_128),
.Y(n_165)
);

CKINVDCx5p33_ASAP7_75t_R g166 ( 
.A(n_56),
.Y(n_166)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_139),
.Y(n_167)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_61),
.Y(n_168)
);

CKINVDCx20_ASAP7_75t_R g169 ( 
.A(n_36),
.Y(n_169)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_40),
.Y(n_170)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_53),
.Y(n_171)
);

CKINVDCx5p33_ASAP7_75t_R g172 ( 
.A(n_48),
.Y(n_172)
);

CKINVDCx20_ASAP7_75t_R g173 ( 
.A(n_142),
.Y(n_173)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_11),
.Y(n_174)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_141),
.Y(n_175)
);

CKINVDCx5p33_ASAP7_75t_R g176 ( 
.A(n_14),
.Y(n_176)
);

CKINVDCx5p33_ASAP7_75t_R g177 ( 
.A(n_14),
.Y(n_177)
);

CKINVDCx5p33_ASAP7_75t_R g178 ( 
.A(n_140),
.Y(n_178)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_100),
.Y(n_179)
);

BUFx8_ASAP7_75t_SL g180 ( 
.A(n_117),
.Y(n_180)
);

CKINVDCx5p33_ASAP7_75t_R g181 ( 
.A(n_133),
.Y(n_181)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_96),
.Y(n_182)
);

CKINVDCx16_ASAP7_75t_R g183 ( 
.A(n_134),
.Y(n_183)
);

CKINVDCx5p33_ASAP7_75t_R g184 ( 
.A(n_67),
.Y(n_184)
);

CKINVDCx5p33_ASAP7_75t_R g185 ( 
.A(n_22),
.Y(n_185)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_54),
.Y(n_186)
);

CKINVDCx5p33_ASAP7_75t_R g187 ( 
.A(n_39),
.Y(n_187)
);

CKINVDCx5p33_ASAP7_75t_R g188 ( 
.A(n_49),
.Y(n_188)
);

BUFx3_ASAP7_75t_L g189 ( 
.A(n_52),
.Y(n_189)
);

CKINVDCx5p33_ASAP7_75t_R g190 ( 
.A(n_104),
.Y(n_190)
);

CKINVDCx5p33_ASAP7_75t_R g191 ( 
.A(n_41),
.Y(n_191)
);

CKINVDCx5p33_ASAP7_75t_R g192 ( 
.A(n_48),
.Y(n_192)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_9),
.Y(n_193)
);

INVx1_ASAP7_75t_SL g194 ( 
.A(n_82),
.Y(n_194)
);

CKINVDCx16_ASAP7_75t_R g195 ( 
.A(n_103),
.Y(n_195)
);

CKINVDCx5p33_ASAP7_75t_R g196 ( 
.A(n_81),
.Y(n_196)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_76),
.Y(n_197)
);

CKINVDCx5p33_ASAP7_75t_R g198 ( 
.A(n_146),
.Y(n_198)
);

CKINVDCx5p33_ASAP7_75t_R g199 ( 
.A(n_68),
.Y(n_199)
);

INVx2_ASAP7_75t_L g200 ( 
.A(n_147),
.Y(n_200)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_75),
.Y(n_201)
);

CKINVDCx5p33_ASAP7_75t_R g202 ( 
.A(n_92),
.Y(n_202)
);

CKINVDCx5p33_ASAP7_75t_R g203 ( 
.A(n_85),
.Y(n_203)
);

CKINVDCx14_ASAP7_75t_R g204 ( 
.A(n_10),
.Y(n_204)
);

CKINVDCx5p33_ASAP7_75t_R g205 ( 
.A(n_44),
.Y(n_205)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_24),
.Y(n_206)
);

INVx1_ASAP7_75t_SL g207 ( 
.A(n_62),
.Y(n_207)
);

CKINVDCx5p33_ASAP7_75t_R g208 ( 
.A(n_136),
.Y(n_208)
);

CKINVDCx5p33_ASAP7_75t_R g209 ( 
.A(n_151),
.Y(n_209)
);

INVx2_ASAP7_75t_L g210 ( 
.A(n_113),
.Y(n_210)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_114),
.Y(n_211)
);

CKINVDCx20_ASAP7_75t_R g212 ( 
.A(n_57),
.Y(n_212)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_109),
.Y(n_213)
);

CKINVDCx5p33_ASAP7_75t_R g214 ( 
.A(n_18),
.Y(n_214)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_2),
.Y(n_215)
);

BUFx6f_ASAP7_75t_L g216 ( 
.A(n_77),
.Y(n_216)
);

CKINVDCx5p33_ASAP7_75t_R g217 ( 
.A(n_46),
.Y(n_217)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_135),
.Y(n_218)
);

CKINVDCx20_ASAP7_75t_R g219 ( 
.A(n_99),
.Y(n_219)
);

BUFx2_ASAP7_75t_L g220 ( 
.A(n_31),
.Y(n_220)
);

CKINVDCx20_ASAP7_75t_R g221 ( 
.A(n_123),
.Y(n_221)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_138),
.Y(n_222)
);

INVx2_ASAP7_75t_L g223 ( 
.A(n_152),
.Y(n_223)
);

CKINVDCx5p33_ASAP7_75t_R g224 ( 
.A(n_50),
.Y(n_224)
);

CKINVDCx5p33_ASAP7_75t_R g225 ( 
.A(n_11),
.Y(n_225)
);

CKINVDCx5p33_ASAP7_75t_R g226 ( 
.A(n_130),
.Y(n_226)
);

INVx2_ASAP7_75t_L g227 ( 
.A(n_49),
.Y(n_227)
);

CKINVDCx5p33_ASAP7_75t_R g228 ( 
.A(n_63),
.Y(n_228)
);

CKINVDCx5p33_ASAP7_75t_R g229 ( 
.A(n_116),
.Y(n_229)
);

CKINVDCx5p33_ASAP7_75t_R g230 ( 
.A(n_86),
.Y(n_230)
);

BUFx2_ASAP7_75t_L g231 ( 
.A(n_33),
.Y(n_231)
);

CKINVDCx20_ASAP7_75t_R g232 ( 
.A(n_46),
.Y(n_232)
);

CKINVDCx16_ASAP7_75t_R g233 ( 
.A(n_73),
.Y(n_233)
);

CKINVDCx5p33_ASAP7_75t_R g234 ( 
.A(n_38),
.Y(n_234)
);

CKINVDCx5p33_ASAP7_75t_R g235 ( 
.A(n_9),
.Y(n_235)
);

CKINVDCx5p33_ASAP7_75t_R g236 ( 
.A(n_127),
.Y(n_236)
);

CKINVDCx5p33_ASAP7_75t_R g237 ( 
.A(n_44),
.Y(n_237)
);

CKINVDCx5p33_ASAP7_75t_R g238 ( 
.A(n_17),
.Y(n_238)
);

CKINVDCx5p33_ASAP7_75t_R g239 ( 
.A(n_90),
.Y(n_239)
);

INVx2_ASAP7_75t_L g240 ( 
.A(n_21),
.Y(n_240)
);

CKINVDCx5p33_ASAP7_75t_R g241 ( 
.A(n_153),
.Y(n_241)
);

CKINVDCx5p33_ASAP7_75t_R g242 ( 
.A(n_97),
.Y(n_242)
);

CKINVDCx5p33_ASAP7_75t_R g243 ( 
.A(n_58),
.Y(n_243)
);

CKINVDCx5p33_ASAP7_75t_R g244 ( 
.A(n_0),
.Y(n_244)
);

CKINVDCx20_ASAP7_75t_R g245 ( 
.A(n_51),
.Y(n_245)
);

CKINVDCx5p33_ASAP7_75t_R g246 ( 
.A(n_27),
.Y(n_246)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_34),
.Y(n_247)
);

CKINVDCx5p33_ASAP7_75t_R g248 ( 
.A(n_20),
.Y(n_248)
);

CKINVDCx5p33_ASAP7_75t_R g249 ( 
.A(n_84),
.Y(n_249)
);

CKINVDCx5p33_ASAP7_75t_R g250 ( 
.A(n_50),
.Y(n_250)
);

CKINVDCx20_ASAP7_75t_R g251 ( 
.A(n_105),
.Y(n_251)
);

CKINVDCx5p33_ASAP7_75t_R g252 ( 
.A(n_15),
.Y(n_252)
);

BUFx5_ASAP7_75t_L g253 ( 
.A(n_65),
.Y(n_253)
);

INVx2_ASAP7_75t_L g254 ( 
.A(n_129),
.Y(n_254)
);

CKINVDCx5p33_ASAP7_75t_R g255 ( 
.A(n_149),
.Y(n_255)
);

CKINVDCx5p33_ASAP7_75t_R g256 ( 
.A(n_32),
.Y(n_256)
);

BUFx10_ASAP7_75t_L g257 ( 
.A(n_0),
.Y(n_257)
);

CKINVDCx5p33_ASAP7_75t_R g258 ( 
.A(n_19),
.Y(n_258)
);

CKINVDCx5p33_ASAP7_75t_R g259 ( 
.A(n_91),
.Y(n_259)
);

INVx2_ASAP7_75t_L g260 ( 
.A(n_60),
.Y(n_260)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_89),
.Y(n_261)
);

CKINVDCx5p33_ASAP7_75t_R g262 ( 
.A(n_45),
.Y(n_262)
);

INVx3_ASAP7_75t_L g263 ( 
.A(n_98),
.Y(n_263)
);

CKINVDCx5p33_ASAP7_75t_R g264 ( 
.A(n_111),
.Y(n_264)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_3),
.Y(n_265)
);

CKINVDCx5p33_ASAP7_75t_R g266 ( 
.A(n_1),
.Y(n_266)
);

CKINVDCx5p33_ASAP7_75t_R g267 ( 
.A(n_34),
.Y(n_267)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_110),
.Y(n_268)
);

CKINVDCx5p33_ASAP7_75t_R g269 ( 
.A(n_28),
.Y(n_269)
);

CKINVDCx5p33_ASAP7_75t_R g270 ( 
.A(n_33),
.Y(n_270)
);

BUFx5_ASAP7_75t_L g271 ( 
.A(n_52),
.Y(n_271)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_4),
.Y(n_272)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_41),
.Y(n_273)
);

INVx2_ASAP7_75t_L g274 ( 
.A(n_79),
.Y(n_274)
);

BUFx3_ASAP7_75t_L g275 ( 
.A(n_131),
.Y(n_275)
);

CKINVDCx5p33_ASAP7_75t_R g276 ( 
.A(n_118),
.Y(n_276)
);

CKINVDCx5p33_ASAP7_75t_R g277 ( 
.A(n_51),
.Y(n_277)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_40),
.Y(n_278)
);

CKINVDCx5p33_ASAP7_75t_R g279 ( 
.A(n_74),
.Y(n_279)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_93),
.Y(n_280)
);

CKINVDCx14_ASAP7_75t_R g281 ( 
.A(n_3),
.Y(n_281)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_35),
.Y(n_282)
);

BUFx6f_ASAP7_75t_L g283 ( 
.A(n_126),
.Y(n_283)
);

CKINVDCx5p33_ASAP7_75t_R g284 ( 
.A(n_16),
.Y(n_284)
);

CKINVDCx5p33_ASAP7_75t_R g285 ( 
.A(n_20),
.Y(n_285)
);

CKINVDCx5p33_ASAP7_75t_R g286 ( 
.A(n_54),
.Y(n_286)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_101),
.Y(n_287)
);

CKINVDCx5p33_ASAP7_75t_R g288 ( 
.A(n_30),
.Y(n_288)
);

CKINVDCx5p33_ASAP7_75t_R g289 ( 
.A(n_12),
.Y(n_289)
);

INVx2_ASAP7_75t_SL g290 ( 
.A(n_38),
.Y(n_290)
);

CKINVDCx5p33_ASAP7_75t_R g291 ( 
.A(n_27),
.Y(n_291)
);

CKINVDCx5p33_ASAP7_75t_R g292 ( 
.A(n_72),
.Y(n_292)
);

CKINVDCx5p33_ASAP7_75t_R g293 ( 
.A(n_21),
.Y(n_293)
);

CKINVDCx5p33_ASAP7_75t_R g294 ( 
.A(n_29),
.Y(n_294)
);

CKINVDCx5p33_ASAP7_75t_R g295 ( 
.A(n_32),
.Y(n_295)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_8),
.Y(n_296)
);

CKINVDCx5p33_ASAP7_75t_R g297 ( 
.A(n_83),
.Y(n_297)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_55),
.Y(n_298)
);

CKINVDCx20_ASAP7_75t_R g299 ( 
.A(n_144),
.Y(n_299)
);

CKINVDCx5p33_ASAP7_75t_R g300 ( 
.A(n_39),
.Y(n_300)
);

INVx2_ASAP7_75t_L g301 ( 
.A(n_71),
.Y(n_301)
);

CKINVDCx5p33_ASAP7_75t_R g302 ( 
.A(n_42),
.Y(n_302)
);

CKINVDCx5p33_ASAP7_75t_R g303 ( 
.A(n_15),
.Y(n_303)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_150),
.Y(n_304)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_31),
.Y(n_305)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_29),
.Y(n_306)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_47),
.Y(n_307)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_119),
.Y(n_308)
);

INVxp67_ASAP7_75t_SL g309 ( 
.A(n_189),
.Y(n_309)
);

CKINVDCx5p33_ASAP7_75t_R g310 ( 
.A(n_180),
.Y(n_310)
);

NOR2xp33_ASAP7_75t_L g311 ( 
.A(n_204),
.B(n_281),
.Y(n_311)
);

CKINVDCx20_ASAP7_75t_R g312 ( 
.A(n_162),
.Y(n_312)
);

INVxp67_ASAP7_75t_L g313 ( 
.A(n_220),
.Y(n_313)
);

NAND2xp5_ASAP7_75t_L g314 ( 
.A(n_271),
.B(n_1),
.Y(n_314)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_271),
.Y(n_315)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_271),
.Y(n_316)
);

CKINVDCx5p33_ASAP7_75t_R g317 ( 
.A(n_173),
.Y(n_317)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_271),
.Y(n_318)
);

NOR2xp67_ASAP7_75t_L g319 ( 
.A(n_290),
.B(n_2),
.Y(n_319)
);

INVx2_ASAP7_75t_L g320 ( 
.A(n_271),
.Y(n_320)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_271),
.Y(n_321)
);

CKINVDCx20_ASAP7_75t_R g322 ( 
.A(n_212),
.Y(n_322)
);

INVxp67_ASAP7_75t_L g323 ( 
.A(n_231),
.Y(n_323)
);

CKINVDCx20_ASAP7_75t_R g324 ( 
.A(n_219),
.Y(n_324)
);

CKINVDCx20_ASAP7_75t_R g325 ( 
.A(n_221),
.Y(n_325)
);

CKINVDCx5p33_ASAP7_75t_R g326 ( 
.A(n_251),
.Y(n_326)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_271),
.Y(n_327)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_271),
.Y(n_328)
);

CKINVDCx5p33_ASAP7_75t_R g329 ( 
.A(n_299),
.Y(n_329)
);

INVxp67_ASAP7_75t_SL g330 ( 
.A(n_189),
.Y(n_330)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_155),
.Y(n_331)
);

CKINVDCx20_ASAP7_75t_R g332 ( 
.A(n_163),
.Y(n_332)
);

CKINVDCx20_ASAP7_75t_R g333 ( 
.A(n_169),
.Y(n_333)
);

CKINVDCx5p33_ASAP7_75t_R g334 ( 
.A(n_185),
.Y(n_334)
);

CKINVDCx5p33_ASAP7_75t_R g335 ( 
.A(n_187),
.Y(n_335)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_155),
.Y(n_336)
);

CKINVDCx20_ASAP7_75t_R g337 ( 
.A(n_232),
.Y(n_337)
);

INVx1_ASAP7_75t_L g338 ( 
.A(n_155),
.Y(n_338)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_155),
.Y(n_339)
);

CKINVDCx20_ASAP7_75t_R g340 ( 
.A(n_245),
.Y(n_340)
);

CKINVDCx5p33_ASAP7_75t_R g341 ( 
.A(n_188),
.Y(n_341)
);

INVx1_ASAP7_75t_L g342 ( 
.A(n_155),
.Y(n_342)
);

CKINVDCx5p33_ASAP7_75t_R g343 ( 
.A(n_191),
.Y(n_343)
);

CKINVDCx20_ASAP7_75t_R g344 ( 
.A(n_183),
.Y(n_344)
);

CKINVDCx20_ASAP7_75t_R g345 ( 
.A(n_195),
.Y(n_345)
);

INVxp67_ASAP7_75t_SL g346 ( 
.A(n_227),
.Y(n_346)
);

CKINVDCx20_ASAP7_75t_R g347 ( 
.A(n_233),
.Y(n_347)
);

NOR2xp33_ASAP7_75t_L g348 ( 
.A(n_263),
.B(n_4),
.Y(n_348)
);

INVx1_ASAP7_75t_L g349 ( 
.A(n_227),
.Y(n_349)
);

CKINVDCx20_ASAP7_75t_R g350 ( 
.A(n_158),
.Y(n_350)
);

INVx1_ASAP7_75t_L g351 ( 
.A(n_240),
.Y(n_351)
);

INVx1_ASAP7_75t_L g352 ( 
.A(n_240),
.Y(n_352)
);

CKINVDCx5p33_ASAP7_75t_R g353 ( 
.A(n_192),
.Y(n_353)
);

CKINVDCx20_ASAP7_75t_R g354 ( 
.A(n_275),
.Y(n_354)
);

CKINVDCx20_ASAP7_75t_R g355 ( 
.A(n_275),
.Y(n_355)
);

INVx1_ASAP7_75t_L g356 ( 
.A(n_200),
.Y(n_356)
);

INVx1_ASAP7_75t_L g357 ( 
.A(n_200),
.Y(n_357)
);

CKINVDCx5p33_ASAP7_75t_R g358 ( 
.A(n_205),
.Y(n_358)
);

INVx1_ASAP7_75t_L g359 ( 
.A(n_156),
.Y(n_359)
);

INVxp33_ASAP7_75t_L g360 ( 
.A(n_170),
.Y(n_360)
);

CKINVDCx5p33_ASAP7_75t_R g361 ( 
.A(n_214),
.Y(n_361)
);

INVx1_ASAP7_75t_L g362 ( 
.A(n_171),
.Y(n_362)
);

CKINVDCx5p33_ASAP7_75t_R g363 ( 
.A(n_217),
.Y(n_363)
);

CKINVDCx5p33_ASAP7_75t_R g364 ( 
.A(n_224),
.Y(n_364)
);

INVx1_ASAP7_75t_L g365 ( 
.A(n_210),
.Y(n_365)
);

CKINVDCx5p33_ASAP7_75t_R g366 ( 
.A(n_225),
.Y(n_366)
);

INVx3_ASAP7_75t_L g367 ( 
.A(n_174),
.Y(n_367)
);

INVxp67_ASAP7_75t_L g368 ( 
.A(n_290),
.Y(n_368)
);

INVx1_ASAP7_75t_L g369 ( 
.A(n_210),
.Y(n_369)
);

INVx1_ASAP7_75t_L g370 ( 
.A(n_223),
.Y(n_370)
);

INVx1_ASAP7_75t_L g371 ( 
.A(n_223),
.Y(n_371)
);

INVx1_ASAP7_75t_L g372 ( 
.A(n_254),
.Y(n_372)
);

INVx1_ASAP7_75t_L g373 ( 
.A(n_254),
.Y(n_373)
);

INVx3_ASAP7_75t_L g374 ( 
.A(n_186),
.Y(n_374)
);

INVxp33_ASAP7_75t_SL g375 ( 
.A(n_157),
.Y(n_375)
);

INVxp67_ASAP7_75t_L g376 ( 
.A(n_257),
.Y(n_376)
);

INVxp33_ASAP7_75t_SL g377 ( 
.A(n_157),
.Y(n_377)
);

INVx1_ASAP7_75t_L g378 ( 
.A(n_260),
.Y(n_378)
);

INVx1_ASAP7_75t_L g379 ( 
.A(n_260),
.Y(n_379)
);

NAND2xp5_ASAP7_75t_L g380 ( 
.A(n_315),
.B(n_159),
.Y(n_380)
);

NAND2xp5_ASAP7_75t_L g381 ( 
.A(n_315),
.B(n_167),
.Y(n_381)
);

INVxp33_ASAP7_75t_SL g382 ( 
.A(n_310),
.Y(n_382)
);

INVx1_ASAP7_75t_L g383 ( 
.A(n_316),
.Y(n_383)
);

INVx1_ASAP7_75t_L g384 ( 
.A(n_316),
.Y(n_384)
);

HB1xp67_ASAP7_75t_L g385 ( 
.A(n_313),
.Y(n_385)
);

HB1xp67_ASAP7_75t_L g386 ( 
.A(n_323),
.Y(n_386)
);

INVx2_ASAP7_75t_L g387 ( 
.A(n_320),
.Y(n_387)
);

INVx3_ASAP7_75t_L g388 ( 
.A(n_320),
.Y(n_388)
);

BUFx6f_ASAP7_75t_L g389 ( 
.A(n_318),
.Y(n_389)
);

INVx2_ASAP7_75t_L g390 ( 
.A(n_318),
.Y(n_390)
);

BUFx6f_ASAP7_75t_L g391 ( 
.A(n_321),
.Y(n_391)
);

NOR2xp33_ASAP7_75t_L g392 ( 
.A(n_311),
.B(n_263),
.Y(n_392)
);

CKINVDCx20_ASAP7_75t_R g393 ( 
.A(n_332),
.Y(n_393)
);

INVx1_ASAP7_75t_L g394 ( 
.A(n_321),
.Y(n_394)
);

BUFx6f_ASAP7_75t_L g395 ( 
.A(n_327),
.Y(n_395)
);

INVx1_ASAP7_75t_L g396 ( 
.A(n_327),
.Y(n_396)
);

INVx1_ASAP7_75t_L g397 ( 
.A(n_328),
.Y(n_397)
);

BUFx6f_ASAP7_75t_L g398 ( 
.A(n_328),
.Y(n_398)
);

BUFx6f_ASAP7_75t_L g399 ( 
.A(n_331),
.Y(n_399)
);

INVx1_ASAP7_75t_L g400 ( 
.A(n_314),
.Y(n_400)
);

HB1xp67_ASAP7_75t_L g401 ( 
.A(n_334),
.Y(n_401)
);

INVx2_ASAP7_75t_L g402 ( 
.A(n_331),
.Y(n_402)
);

INVxp67_ASAP7_75t_L g403 ( 
.A(n_309),
.Y(n_403)
);

NOR2xp33_ASAP7_75t_L g404 ( 
.A(n_330),
.B(n_263),
.Y(n_404)
);

AND2x2_ASAP7_75t_L g405 ( 
.A(n_346),
.B(n_193),
.Y(n_405)
);

AND2x2_ASAP7_75t_L g406 ( 
.A(n_360),
.B(n_206),
.Y(n_406)
);

AND2x2_ASAP7_75t_L g407 ( 
.A(n_367),
.B(n_215),
.Y(n_407)
);

INVx2_ASAP7_75t_L g408 ( 
.A(n_336),
.Y(n_408)
);

BUFx3_ASAP7_75t_L g409 ( 
.A(n_356),
.Y(n_409)
);

BUFx6f_ASAP7_75t_L g410 ( 
.A(n_336),
.Y(n_410)
);

INVx1_ASAP7_75t_L g411 ( 
.A(n_338),
.Y(n_411)
);

INVx2_ASAP7_75t_L g412 ( 
.A(n_338),
.Y(n_412)
);

AND2x4_ASAP7_75t_L g413 ( 
.A(n_356),
.B(n_247),
.Y(n_413)
);

OAI22xp5_ASAP7_75t_SL g414 ( 
.A1(n_333),
.A2(n_177),
.B1(n_176),
.B2(n_172),
.Y(n_414)
);

INVx1_ASAP7_75t_L g415 ( 
.A(n_339),
.Y(n_415)
);

BUFx6f_ASAP7_75t_L g416 ( 
.A(n_339),
.Y(n_416)
);

NAND2xp5_ASAP7_75t_L g417 ( 
.A(n_357),
.B(n_168),
.Y(n_417)
);

AND2x2_ASAP7_75t_L g418 ( 
.A(n_367),
.B(n_265),
.Y(n_418)
);

INVx1_ASAP7_75t_L g419 ( 
.A(n_342),
.Y(n_419)
);

NAND2xp5_ASAP7_75t_L g420 ( 
.A(n_357),
.B(n_175),
.Y(n_420)
);

AND2x2_ASAP7_75t_L g421 ( 
.A(n_367),
.B(n_272),
.Y(n_421)
);

AND2x2_ASAP7_75t_L g422 ( 
.A(n_374),
.B(n_365),
.Y(n_422)
);

NAND2xp5_ASAP7_75t_L g423 ( 
.A(n_365),
.B(n_179),
.Y(n_423)
);

INVx2_ASAP7_75t_L g424 ( 
.A(n_342),
.Y(n_424)
);

OAI22xp5_ASAP7_75t_SL g425 ( 
.A1(n_337),
.A2(n_172),
.B1(n_258),
.B2(n_176),
.Y(n_425)
);

INVx1_ASAP7_75t_L g426 ( 
.A(n_369),
.Y(n_426)
);

INVx2_ASAP7_75t_L g427 ( 
.A(n_369),
.Y(n_427)
);

INVx2_ASAP7_75t_L g428 ( 
.A(n_379),
.Y(n_428)
);

INVx1_ASAP7_75t_SL g429 ( 
.A(n_317),
.Y(n_429)
);

AND2x2_ASAP7_75t_L g430 ( 
.A(n_374),
.B(n_273),
.Y(n_430)
);

INVx1_ASAP7_75t_L g431 ( 
.A(n_370),
.Y(n_431)
);

AND3x2_ASAP7_75t_L g432 ( 
.A(n_376),
.B(n_301),
.C(n_274),
.Y(n_432)
);

NAND2xp5_ASAP7_75t_L g433 ( 
.A(n_370),
.B(n_371),
.Y(n_433)
);

INVx2_ASAP7_75t_L g434 ( 
.A(n_371),
.Y(n_434)
);

INVx2_ASAP7_75t_L g435 ( 
.A(n_379),
.Y(n_435)
);

NAND2xp5_ASAP7_75t_L g436 ( 
.A(n_372),
.B(n_182),
.Y(n_436)
);

INVx1_ASAP7_75t_L g437 ( 
.A(n_372),
.Y(n_437)
);

INVx1_ASAP7_75t_L g438 ( 
.A(n_373),
.Y(n_438)
);

INVx3_ASAP7_75t_L g439 ( 
.A(n_373),
.Y(n_439)
);

NOR2xp33_ASAP7_75t_SL g440 ( 
.A(n_350),
.B(n_257),
.Y(n_440)
);

AND2x4_ASAP7_75t_L g441 ( 
.A(n_378),
.B(n_278),
.Y(n_441)
);

INVx1_ASAP7_75t_L g442 ( 
.A(n_378),
.Y(n_442)
);

OAI22xp5_ASAP7_75t_SL g443 ( 
.A1(n_340),
.A2(n_267),
.B1(n_177),
.B2(n_258),
.Y(n_443)
);

INVx1_ASAP7_75t_L g444 ( 
.A(n_348),
.Y(n_444)
);

INVx2_ASAP7_75t_L g445 ( 
.A(n_390),
.Y(n_445)
);

INVx2_ASAP7_75t_L g446 ( 
.A(n_390),
.Y(n_446)
);

AOI22xp33_ASAP7_75t_L g447 ( 
.A1(n_406),
.A2(n_319),
.B1(n_375),
.B2(n_377),
.Y(n_447)
);

AND2x2_ASAP7_75t_L g448 ( 
.A(n_422),
.B(n_374),
.Y(n_448)
);

OAI22xp5_ASAP7_75t_L g449 ( 
.A1(n_444),
.A2(n_288),
.B1(n_262),
.B2(n_266),
.Y(n_449)
);

INVx4_ASAP7_75t_L g450 ( 
.A(n_389),
.Y(n_450)
);

CKINVDCx5p33_ASAP7_75t_R g451 ( 
.A(n_382),
.Y(n_451)
);

AOI22xp33_ASAP7_75t_L g452 ( 
.A1(n_406),
.A2(n_354),
.B1(n_355),
.B2(n_282),
.Y(n_452)
);

INVx2_ASAP7_75t_SL g453 ( 
.A(n_406),
.Y(n_453)
);

INVx1_ASAP7_75t_L g454 ( 
.A(n_390),
.Y(n_454)
);

NAND2xp5_ASAP7_75t_L g455 ( 
.A(n_392),
.B(n_335),
.Y(n_455)
);

AOI22xp5_ASAP7_75t_L g456 ( 
.A1(n_414),
.A2(n_284),
.B1(n_262),
.B2(n_266),
.Y(n_456)
);

AND2x2_ASAP7_75t_L g457 ( 
.A(n_422),
.B(n_368),
.Y(n_457)
);

NAND2xp5_ASAP7_75t_L g458 ( 
.A(n_392),
.B(n_341),
.Y(n_458)
);

INVx2_ASAP7_75t_L g459 ( 
.A(n_390),
.Y(n_459)
);

NAND2xp5_ASAP7_75t_L g460 ( 
.A(n_400),
.B(n_343),
.Y(n_460)
);

NAND2xp5_ASAP7_75t_L g461 ( 
.A(n_400),
.B(n_353),
.Y(n_461)
);

NOR2xp33_ASAP7_75t_L g462 ( 
.A(n_403),
.B(n_358),
.Y(n_462)
);

INVx2_ASAP7_75t_L g463 ( 
.A(n_387),
.Y(n_463)
);

BUFx2_ASAP7_75t_L g464 ( 
.A(n_385),
.Y(n_464)
);

OR2x6_ASAP7_75t_L g465 ( 
.A(n_413),
.B(n_359),
.Y(n_465)
);

INVx1_ASAP7_75t_L g466 ( 
.A(n_411),
.Y(n_466)
);

NOR2x1p5_ASAP7_75t_L g467 ( 
.A(n_382),
.B(n_361),
.Y(n_467)
);

INVx4_ASAP7_75t_L g468 ( 
.A(n_389),
.Y(n_468)
);

INVx2_ASAP7_75t_L g469 ( 
.A(n_387),
.Y(n_469)
);

NAND2xp5_ASAP7_75t_SL g470 ( 
.A(n_401),
.B(n_363),
.Y(n_470)
);

AOI22xp33_ASAP7_75t_L g471 ( 
.A1(n_413),
.A2(n_298),
.B1(n_296),
.B2(n_305),
.Y(n_471)
);

NAND2xp5_ASAP7_75t_SL g472 ( 
.A(n_401),
.B(n_364),
.Y(n_472)
);

BUFx10_ASAP7_75t_L g473 ( 
.A(n_404),
.Y(n_473)
);

INVx3_ASAP7_75t_L g474 ( 
.A(n_389),
.Y(n_474)
);

NOR2xp33_ASAP7_75t_L g475 ( 
.A(n_403),
.B(n_366),
.Y(n_475)
);

INVx3_ASAP7_75t_L g476 ( 
.A(n_389),
.Y(n_476)
);

INVx1_ASAP7_75t_L g477 ( 
.A(n_411),
.Y(n_477)
);

CKINVDCx5p33_ASAP7_75t_R g478 ( 
.A(n_429),
.Y(n_478)
);

INVx2_ASAP7_75t_L g479 ( 
.A(n_387),
.Y(n_479)
);

INVx1_ASAP7_75t_L g480 ( 
.A(n_411),
.Y(n_480)
);

INVx1_ASAP7_75t_L g481 ( 
.A(n_415),
.Y(n_481)
);

INVx2_ASAP7_75t_L g482 ( 
.A(n_387),
.Y(n_482)
);

NAND2xp5_ASAP7_75t_L g483 ( 
.A(n_400),
.B(n_362),
.Y(n_483)
);

INVx1_ASAP7_75t_L g484 ( 
.A(n_415),
.Y(n_484)
);

AND2x2_ASAP7_75t_L g485 ( 
.A(n_422),
.B(n_349),
.Y(n_485)
);

NOR2xp33_ASAP7_75t_L g486 ( 
.A(n_444),
.B(n_344),
.Y(n_486)
);

INVx2_ASAP7_75t_L g487 ( 
.A(n_388),
.Y(n_487)
);

OR2x2_ASAP7_75t_L g488 ( 
.A(n_385),
.B(n_326),
.Y(n_488)
);

XOR2xp5_ASAP7_75t_L g489 ( 
.A(n_393),
.B(n_312),
.Y(n_489)
);

NAND2xp5_ASAP7_75t_SL g490 ( 
.A(n_404),
.B(n_329),
.Y(n_490)
);

NAND2xp5_ASAP7_75t_L g491 ( 
.A(n_444),
.B(n_194),
.Y(n_491)
);

INVx2_ASAP7_75t_L g492 ( 
.A(n_388),
.Y(n_492)
);

INVx3_ASAP7_75t_L g493 ( 
.A(n_389),
.Y(n_493)
);

NAND2xp33_ASAP7_75t_L g494 ( 
.A(n_389),
.B(n_253),
.Y(n_494)
);

BUFx6f_ASAP7_75t_L g495 ( 
.A(n_389),
.Y(n_495)
);

INVx1_ASAP7_75t_SL g496 ( 
.A(n_429),
.Y(n_496)
);

NAND2xp5_ASAP7_75t_SL g497 ( 
.A(n_405),
.B(n_160),
.Y(n_497)
);

INVx1_ASAP7_75t_L g498 ( 
.A(n_415),
.Y(n_498)
);

INVx1_ASAP7_75t_L g499 ( 
.A(n_419),
.Y(n_499)
);

INVx4_ASAP7_75t_L g500 ( 
.A(n_389),
.Y(n_500)
);

AOI22xp33_ASAP7_75t_L g501 ( 
.A1(n_413),
.A2(n_306),
.B1(n_307),
.B2(n_257),
.Y(n_501)
);

NOR2xp33_ASAP7_75t_SL g502 ( 
.A(n_440),
.B(n_345),
.Y(n_502)
);

AND2x6_ASAP7_75t_L g503 ( 
.A(n_388),
.B(n_274),
.Y(n_503)
);

AND2x2_ASAP7_75t_L g504 ( 
.A(n_407),
.B(n_349),
.Y(n_504)
);

INVx1_ASAP7_75t_L g505 ( 
.A(n_419),
.Y(n_505)
);

NAND2xp5_ASAP7_75t_L g506 ( 
.A(n_383),
.B(n_384),
.Y(n_506)
);

INVx1_ASAP7_75t_L g507 ( 
.A(n_419),
.Y(n_507)
);

BUFx10_ASAP7_75t_L g508 ( 
.A(n_432),
.Y(n_508)
);

NOR2xp33_ASAP7_75t_L g509 ( 
.A(n_383),
.B(n_347),
.Y(n_509)
);

NAND2xp5_ASAP7_75t_L g510 ( 
.A(n_384),
.B(n_207),
.Y(n_510)
);

INVx2_ASAP7_75t_L g511 ( 
.A(n_388),
.Y(n_511)
);

INVx1_ASAP7_75t_L g512 ( 
.A(n_384),
.Y(n_512)
);

INVx2_ASAP7_75t_L g513 ( 
.A(n_388),
.Y(n_513)
);

INVx1_ASAP7_75t_L g514 ( 
.A(n_394),
.Y(n_514)
);

NOR2xp33_ASAP7_75t_L g515 ( 
.A(n_394),
.B(n_322),
.Y(n_515)
);

INVx2_ASAP7_75t_L g516 ( 
.A(n_402),
.Y(n_516)
);

NAND2xp5_ASAP7_75t_L g517 ( 
.A(n_394),
.B(n_160),
.Y(n_517)
);

NOR2xp33_ASAP7_75t_L g518 ( 
.A(n_396),
.B(n_324),
.Y(n_518)
);

INVx4_ASAP7_75t_L g519 ( 
.A(n_389),
.Y(n_519)
);

NOR2x1p5_ASAP7_75t_L g520 ( 
.A(n_405),
.B(n_267),
.Y(n_520)
);

NAND2xp5_ASAP7_75t_L g521 ( 
.A(n_396),
.B(n_164),
.Y(n_521)
);

INVx4_ASAP7_75t_L g522 ( 
.A(n_391),
.Y(n_522)
);

INVx2_ASAP7_75t_SL g523 ( 
.A(n_386),
.Y(n_523)
);

INVx3_ASAP7_75t_L g524 ( 
.A(n_391),
.Y(n_524)
);

INVx1_ASAP7_75t_L g525 ( 
.A(n_396),
.Y(n_525)
);

INVx2_ASAP7_75t_SL g526 ( 
.A(n_386),
.Y(n_526)
);

BUFx6f_ASAP7_75t_SL g527 ( 
.A(n_413),
.Y(n_527)
);

CKINVDCx5p33_ASAP7_75t_R g528 ( 
.A(n_393),
.Y(n_528)
);

INVx1_ASAP7_75t_L g529 ( 
.A(n_397),
.Y(n_529)
);

INVx1_ASAP7_75t_SL g530 ( 
.A(n_414),
.Y(n_530)
);

INVxp67_ASAP7_75t_L g531 ( 
.A(n_440),
.Y(n_531)
);

NAND2xp5_ASAP7_75t_SL g532 ( 
.A(n_405),
.B(n_164),
.Y(n_532)
);

INVx2_ASAP7_75t_L g533 ( 
.A(n_402),
.Y(n_533)
);

INVx3_ASAP7_75t_L g534 ( 
.A(n_391),
.Y(n_534)
);

OAI22xp5_ASAP7_75t_L g535 ( 
.A1(n_397),
.A2(n_269),
.B1(n_270),
.B2(n_277),
.Y(n_535)
);

AOI22xp33_ASAP7_75t_L g536 ( 
.A1(n_413),
.A2(n_352),
.B1(n_351),
.B2(n_234),
.Y(n_536)
);

OR2x2_ASAP7_75t_L g537 ( 
.A(n_425),
.B(n_269),
.Y(n_537)
);

INVx4_ASAP7_75t_L g538 ( 
.A(n_391),
.Y(n_538)
);

NAND2xp5_ASAP7_75t_SL g539 ( 
.A(n_441),
.B(n_165),
.Y(n_539)
);

INVx2_ASAP7_75t_L g540 ( 
.A(n_402),
.Y(n_540)
);

INVx2_ASAP7_75t_L g541 ( 
.A(n_402),
.Y(n_541)
);

NOR2xp33_ASAP7_75t_L g542 ( 
.A(n_397),
.B(n_325),
.Y(n_542)
);

NAND2xp5_ASAP7_75t_SL g543 ( 
.A(n_441),
.B(n_165),
.Y(n_543)
);

INVx1_ASAP7_75t_L g544 ( 
.A(n_427),
.Y(n_544)
);

NAND2xp5_ASAP7_75t_SL g545 ( 
.A(n_441),
.B(n_166),
.Y(n_545)
);

NAND2xp5_ASAP7_75t_L g546 ( 
.A(n_409),
.B(n_166),
.Y(n_546)
);

NAND2xp5_ASAP7_75t_SL g547 ( 
.A(n_441),
.B(n_178),
.Y(n_547)
);

AND2x2_ASAP7_75t_L g548 ( 
.A(n_407),
.B(n_270),
.Y(n_548)
);

INVx2_ASAP7_75t_L g549 ( 
.A(n_408),
.Y(n_549)
);

INVx3_ASAP7_75t_L g550 ( 
.A(n_391),
.Y(n_550)
);

BUFx6f_ASAP7_75t_L g551 ( 
.A(n_391),
.Y(n_551)
);

NAND2xp5_ASAP7_75t_SL g552 ( 
.A(n_441),
.B(n_178),
.Y(n_552)
);

NOR2xp33_ASAP7_75t_SL g553 ( 
.A(n_443),
.B(n_277),
.Y(n_553)
);

NOR2xp33_ASAP7_75t_L g554 ( 
.A(n_437),
.B(n_197),
.Y(n_554)
);

INVx4_ASAP7_75t_L g555 ( 
.A(n_391),
.Y(n_555)
);

AND2x2_ASAP7_75t_L g556 ( 
.A(n_407),
.B(n_284),
.Y(n_556)
);

NOR2xp33_ASAP7_75t_L g557 ( 
.A(n_437),
.B(n_201),
.Y(n_557)
);

NAND2xp33_ASAP7_75t_L g558 ( 
.A(n_391),
.B(n_253),
.Y(n_558)
);

INVx3_ASAP7_75t_L g559 ( 
.A(n_391),
.Y(n_559)
);

INVx1_ASAP7_75t_L g560 ( 
.A(n_427),
.Y(n_560)
);

INVx1_ASAP7_75t_SL g561 ( 
.A(n_425),
.Y(n_561)
);

BUFx6f_ASAP7_75t_L g562 ( 
.A(n_395),
.Y(n_562)
);

INVx2_ASAP7_75t_L g563 ( 
.A(n_408),
.Y(n_563)
);

BUFx2_ASAP7_75t_L g564 ( 
.A(n_443),
.Y(n_564)
);

NAND2xp5_ASAP7_75t_L g565 ( 
.A(n_409),
.B(n_181),
.Y(n_565)
);

NOR2xp33_ASAP7_75t_L g566 ( 
.A(n_426),
.B(n_211),
.Y(n_566)
);

INVx1_ASAP7_75t_L g567 ( 
.A(n_427),
.Y(n_567)
);

AND2x2_ASAP7_75t_L g568 ( 
.A(n_418),
.B(n_285),
.Y(n_568)
);

AO22x2_ASAP7_75t_L g569 ( 
.A1(n_441),
.A2(n_308),
.B1(n_304),
.B2(n_218),
.Y(n_569)
);

INVxp67_ASAP7_75t_SL g570 ( 
.A(n_395),
.Y(n_570)
);

INVx2_ASAP7_75t_L g571 ( 
.A(n_408),
.Y(n_571)
);

NAND2xp5_ASAP7_75t_SL g572 ( 
.A(n_418),
.B(n_181),
.Y(n_572)
);

INVx3_ASAP7_75t_L g573 ( 
.A(n_395),
.Y(n_573)
);

INVx1_ASAP7_75t_L g574 ( 
.A(n_427),
.Y(n_574)
);

INVx2_ASAP7_75t_L g575 ( 
.A(n_408),
.Y(n_575)
);

INVx1_ASAP7_75t_L g576 ( 
.A(n_428),
.Y(n_576)
);

NOR2xp33_ASAP7_75t_L g577 ( 
.A(n_426),
.B(n_213),
.Y(n_577)
);

BUFx6f_ASAP7_75t_L g578 ( 
.A(n_395),
.Y(n_578)
);

INVx2_ASAP7_75t_L g579 ( 
.A(n_412),
.Y(n_579)
);

NAND2xp5_ASAP7_75t_L g580 ( 
.A(n_409),
.B(n_259),
.Y(n_580)
);

NAND2xp5_ASAP7_75t_L g581 ( 
.A(n_409),
.B(n_259),
.Y(n_581)
);

INVx2_ASAP7_75t_SL g582 ( 
.A(n_432),
.Y(n_582)
);

INVx4_ASAP7_75t_L g583 ( 
.A(n_395),
.Y(n_583)
);

INVx1_ASAP7_75t_L g584 ( 
.A(n_428),
.Y(n_584)
);

INVx2_ASAP7_75t_L g585 ( 
.A(n_412),
.Y(n_585)
);

CKINVDCx20_ASAP7_75t_R g586 ( 
.A(n_418),
.Y(n_586)
);

OR2x6_ASAP7_75t_L g587 ( 
.A(n_417),
.B(n_222),
.Y(n_587)
);

INVx1_ASAP7_75t_L g588 ( 
.A(n_428),
.Y(n_588)
);

INVx2_ASAP7_75t_L g589 ( 
.A(n_412),
.Y(n_589)
);

INVx1_ASAP7_75t_L g590 ( 
.A(n_428),
.Y(n_590)
);

OAI22xp33_ASAP7_75t_L g591 ( 
.A1(n_417),
.A2(n_303),
.B1(n_302),
.B2(n_285),
.Y(n_591)
);

AND2x2_ASAP7_75t_L g592 ( 
.A(n_496),
.B(n_421),
.Y(n_592)
);

INVx2_ASAP7_75t_SL g593 ( 
.A(n_478),
.Y(n_593)
);

NOR2xp33_ASAP7_75t_L g594 ( 
.A(n_455),
.B(n_380),
.Y(n_594)
);

NAND2xp5_ASAP7_75t_SL g595 ( 
.A(n_462),
.B(n_380),
.Y(n_595)
);

O2A1O1Ixp33_ASAP7_75t_L g596 ( 
.A1(n_491),
.A2(n_381),
.B(n_439),
.C(n_438),
.Y(n_596)
);

NAND2xp33_ASAP7_75t_SL g597 ( 
.A(n_467),
.B(n_421),
.Y(n_597)
);

NAND2xp5_ASAP7_75t_L g598 ( 
.A(n_458),
.B(n_439),
.Y(n_598)
);

NAND2xp5_ASAP7_75t_SL g599 ( 
.A(n_473),
.B(n_395),
.Y(n_599)
);

NAND2xp5_ASAP7_75t_SL g600 ( 
.A(n_473),
.B(n_395),
.Y(n_600)
);

NAND2xp5_ASAP7_75t_L g601 ( 
.A(n_475),
.B(n_439),
.Y(n_601)
);

AND2x4_ASAP7_75t_L g602 ( 
.A(n_453),
.B(n_421),
.Y(n_602)
);

NAND2xp5_ASAP7_75t_SL g603 ( 
.A(n_473),
.B(n_395),
.Y(n_603)
);

INVx2_ASAP7_75t_L g604 ( 
.A(n_463),
.Y(n_604)
);

INVx2_ASAP7_75t_L g605 ( 
.A(n_463),
.Y(n_605)
);

NOR2xp33_ASAP7_75t_L g606 ( 
.A(n_473),
.B(n_460),
.Y(n_606)
);

BUFx8_ASAP7_75t_L g607 ( 
.A(n_464),
.Y(n_607)
);

NOR2xp33_ASAP7_75t_L g608 ( 
.A(n_461),
.B(n_381),
.Y(n_608)
);

AOI22xp5_ASAP7_75t_L g609 ( 
.A1(n_587),
.A2(n_430),
.B1(n_439),
.B2(n_438),
.Y(n_609)
);

OR2x2_ASAP7_75t_L g610 ( 
.A(n_464),
.B(n_430),
.Y(n_610)
);

NOR2xp33_ASAP7_75t_L g611 ( 
.A(n_490),
.B(n_439),
.Y(n_611)
);

AOI22xp33_ASAP7_75t_L g612 ( 
.A1(n_569),
.A2(n_435),
.B1(n_434),
.B2(n_426),
.Y(n_612)
);

INVx2_ASAP7_75t_L g613 ( 
.A(n_469),
.Y(n_613)
);

NAND2xp5_ASAP7_75t_L g614 ( 
.A(n_448),
.B(n_430),
.Y(n_614)
);

AND2x2_ASAP7_75t_L g615 ( 
.A(n_523),
.B(n_431),
.Y(n_615)
);

NOR2xp33_ASAP7_75t_L g616 ( 
.A(n_453),
.B(n_395),
.Y(n_616)
);

NAND2xp5_ASAP7_75t_SL g617 ( 
.A(n_495),
.B(n_398),
.Y(n_617)
);

NAND2xp5_ASAP7_75t_L g618 ( 
.A(n_448),
.B(n_431),
.Y(n_618)
);

INVx2_ASAP7_75t_L g619 ( 
.A(n_469),
.Y(n_619)
);

NAND2xp5_ASAP7_75t_L g620 ( 
.A(n_504),
.B(n_431),
.Y(n_620)
);

NAND2xp5_ASAP7_75t_L g621 ( 
.A(n_504),
.B(n_438),
.Y(n_621)
);

AOI22xp5_ASAP7_75t_L g622 ( 
.A1(n_587),
.A2(n_442),
.B1(n_264),
.B2(n_276),
.Y(n_622)
);

INVx1_ASAP7_75t_L g623 ( 
.A(n_466),
.Y(n_623)
);

O2A1O1Ixp33_ASAP7_75t_L g624 ( 
.A1(n_483),
.A2(n_442),
.B(n_436),
.C(n_420),
.Y(n_624)
);

AO221x1_ASAP7_75t_L g625 ( 
.A1(n_564),
.A2(n_161),
.B1(n_216),
.B2(n_283),
.C(n_268),
.Y(n_625)
);

NAND2xp5_ASAP7_75t_SL g626 ( 
.A(n_495),
.B(n_398),
.Y(n_626)
);

NAND2xp5_ASAP7_75t_L g627 ( 
.A(n_485),
.B(n_442),
.Y(n_627)
);

NOR2xp33_ASAP7_75t_L g628 ( 
.A(n_497),
.B(n_398),
.Y(n_628)
);

NAND2xp5_ASAP7_75t_L g629 ( 
.A(n_485),
.B(n_434),
.Y(n_629)
);

NAND2xp5_ASAP7_75t_SL g630 ( 
.A(n_523),
.B(n_264),
.Y(n_630)
);

INVx2_ASAP7_75t_L g631 ( 
.A(n_479),
.Y(n_631)
);

AOI22xp5_ASAP7_75t_L g632 ( 
.A1(n_587),
.A2(n_276),
.B1(n_279),
.B2(n_436),
.Y(n_632)
);

CKINVDCx5p33_ASAP7_75t_R g633 ( 
.A(n_451),
.Y(n_633)
);

INVx2_ASAP7_75t_L g634 ( 
.A(n_479),
.Y(n_634)
);

INVx2_ASAP7_75t_L g635 ( 
.A(n_482),
.Y(n_635)
);

NAND2xp5_ASAP7_75t_SL g636 ( 
.A(n_495),
.B(n_398),
.Y(n_636)
);

BUFx3_ASAP7_75t_L g637 ( 
.A(n_528),
.Y(n_637)
);

NAND2xp5_ASAP7_75t_L g638 ( 
.A(n_510),
.B(n_434),
.Y(n_638)
);

NAND2xp5_ASAP7_75t_L g639 ( 
.A(n_587),
.B(n_434),
.Y(n_639)
);

O2A1O1Ixp5_ASAP7_75t_L g640 ( 
.A1(n_570),
.A2(n_420),
.B(n_423),
.C(n_435),
.Y(n_640)
);

NAND2xp5_ASAP7_75t_SL g641 ( 
.A(n_495),
.B(n_398),
.Y(n_641)
);

NOR2xp33_ASAP7_75t_L g642 ( 
.A(n_532),
.B(n_398),
.Y(n_642)
);

NAND2xp5_ASAP7_75t_L g643 ( 
.A(n_587),
.B(n_435),
.Y(n_643)
);

NOR2xp67_ASAP7_75t_SL g644 ( 
.A(n_548),
.B(n_286),
.Y(n_644)
);

INVx2_ASAP7_75t_L g645 ( 
.A(n_482),
.Y(n_645)
);

AOI22xp5_ASAP7_75t_L g646 ( 
.A1(n_527),
.A2(n_279),
.B1(n_287),
.B2(n_280),
.Y(n_646)
);

NAND2xp5_ASAP7_75t_L g647 ( 
.A(n_548),
.B(n_435),
.Y(n_647)
);

INVx2_ASAP7_75t_L g648 ( 
.A(n_445),
.Y(n_648)
);

NAND2xp5_ASAP7_75t_L g649 ( 
.A(n_556),
.B(n_433),
.Y(n_649)
);

NAND2xp5_ASAP7_75t_L g650 ( 
.A(n_556),
.B(n_433),
.Y(n_650)
);

INVxp67_ASAP7_75t_L g651 ( 
.A(n_489),
.Y(n_651)
);

NOR2xp33_ASAP7_75t_L g652 ( 
.A(n_572),
.B(n_398),
.Y(n_652)
);

AOI22xp5_ASAP7_75t_L g653 ( 
.A1(n_527),
.A2(n_569),
.B1(n_486),
.B2(n_465),
.Y(n_653)
);

NAND2xp5_ASAP7_75t_L g654 ( 
.A(n_568),
.B(n_457),
.Y(n_654)
);

INVxp67_ASAP7_75t_L g655 ( 
.A(n_489),
.Y(n_655)
);

NAND2xp5_ASAP7_75t_SL g656 ( 
.A(n_526),
.B(n_286),
.Y(n_656)
);

NAND2xp5_ASAP7_75t_SL g657 ( 
.A(n_495),
.B(n_398),
.Y(n_657)
);

INVx3_ASAP7_75t_L g658 ( 
.A(n_527),
.Y(n_658)
);

INVx2_ASAP7_75t_L g659 ( 
.A(n_445),
.Y(n_659)
);

AND2x2_ASAP7_75t_L g660 ( 
.A(n_457),
.B(n_288),
.Y(n_660)
);

INVx1_ASAP7_75t_L g661 ( 
.A(n_466),
.Y(n_661)
);

INVx2_ASAP7_75t_L g662 ( 
.A(n_446),
.Y(n_662)
);

NAND2xp5_ASAP7_75t_L g663 ( 
.A(n_568),
.B(n_398),
.Y(n_663)
);

INVx1_ASAP7_75t_L g664 ( 
.A(n_477),
.Y(n_664)
);

INVx8_ASAP7_75t_L g665 ( 
.A(n_465),
.Y(n_665)
);

NAND2xp5_ASAP7_75t_L g666 ( 
.A(n_465),
.B(n_412),
.Y(n_666)
);

INVx4_ASAP7_75t_L g667 ( 
.A(n_465),
.Y(n_667)
);

NAND2xp33_ASAP7_75t_L g668 ( 
.A(n_551),
.B(n_235),
.Y(n_668)
);

AOI22xp33_ASAP7_75t_L g669 ( 
.A1(n_569),
.A2(n_424),
.B1(n_291),
.B2(n_289),
.Y(n_669)
);

OAI22xp33_ASAP7_75t_L g670 ( 
.A1(n_553),
.A2(n_289),
.B1(n_291),
.B2(n_302),
.Y(n_670)
);

OR2x2_ASAP7_75t_L g671 ( 
.A(n_488),
.B(n_303),
.Y(n_671)
);

O2A1O1Ixp5_ASAP7_75t_L g672 ( 
.A1(n_539),
.A2(n_261),
.B(n_424),
.C(n_238),
.Y(n_672)
);

NOR2xp33_ASAP7_75t_L g673 ( 
.A(n_543),
.B(n_237),
.Y(n_673)
);

NAND2xp5_ASAP7_75t_L g674 ( 
.A(n_465),
.B(n_424),
.Y(n_674)
);

INVx1_ASAP7_75t_L g675 ( 
.A(n_480),
.Y(n_675)
);

NAND2xp5_ASAP7_75t_SL g676 ( 
.A(n_551),
.B(n_399),
.Y(n_676)
);

NAND2xp5_ASAP7_75t_L g677 ( 
.A(n_517),
.B(n_424),
.Y(n_677)
);

INVx2_ASAP7_75t_SL g678 ( 
.A(n_488),
.Y(n_678)
);

AND2x4_ASAP7_75t_L g679 ( 
.A(n_582),
.B(n_244),
.Y(n_679)
);

NAND2xp5_ASAP7_75t_L g680 ( 
.A(n_521),
.B(n_246),
.Y(n_680)
);

NAND2xp33_ASAP7_75t_L g681 ( 
.A(n_551),
.B(n_248),
.Y(n_681)
);

AND2x2_ASAP7_75t_L g682 ( 
.A(n_515),
.B(n_250),
.Y(n_682)
);

INVxp67_ASAP7_75t_L g683 ( 
.A(n_518),
.Y(n_683)
);

INVx2_ASAP7_75t_L g684 ( 
.A(n_446),
.Y(n_684)
);

NAND2xp5_ASAP7_75t_L g685 ( 
.A(n_512),
.B(n_252),
.Y(n_685)
);

INVx2_ASAP7_75t_L g686 ( 
.A(n_459),
.Y(n_686)
);

OAI22xp33_ASAP7_75t_L g687 ( 
.A1(n_456),
.A2(n_256),
.B1(n_293),
.B2(n_294),
.Y(n_687)
);

NAND2xp5_ASAP7_75t_L g688 ( 
.A(n_512),
.B(n_295),
.Y(n_688)
);

INVxp67_ASAP7_75t_L g689 ( 
.A(n_542),
.Y(n_689)
);

AOI22xp33_ASAP7_75t_L g690 ( 
.A1(n_569),
.A2(n_416),
.B1(n_410),
.B2(n_399),
.Y(n_690)
);

INVx1_ASAP7_75t_L g691 ( 
.A(n_480),
.Y(n_691)
);

INVx8_ASAP7_75t_L g692 ( 
.A(n_503),
.Y(n_692)
);

INVxp33_ASAP7_75t_L g693 ( 
.A(n_509),
.Y(n_693)
);

A2O1A1Ixp33_ASAP7_75t_L g694 ( 
.A1(n_514),
.A2(n_300),
.B(n_410),
.C(n_399),
.Y(n_694)
);

NAND2xp5_ASAP7_75t_L g695 ( 
.A(n_514),
.B(n_184),
.Y(n_695)
);

BUFx6f_ASAP7_75t_L g696 ( 
.A(n_551),
.Y(n_696)
);

NAND2xp5_ASAP7_75t_L g697 ( 
.A(n_525),
.B(n_190),
.Y(n_697)
);

HB1xp67_ASAP7_75t_L g698 ( 
.A(n_528),
.Y(n_698)
);

O2A1O1Ixp33_ASAP7_75t_L g699 ( 
.A1(n_506),
.A2(n_5),
.B(n_6),
.C(n_7),
.Y(n_699)
);

NAND2xp5_ASAP7_75t_L g700 ( 
.A(n_525),
.B(n_196),
.Y(n_700)
);

OAI22xp5_ASAP7_75t_SL g701 ( 
.A1(n_564),
.A2(n_230),
.B1(n_198),
.B2(n_199),
.Y(n_701)
);

NAND2xp5_ASAP7_75t_SL g702 ( 
.A(n_447),
.B(n_202),
.Y(n_702)
);

BUFx6f_ASAP7_75t_L g703 ( 
.A(n_551),
.Y(n_703)
);

INVxp67_ASAP7_75t_SL g704 ( 
.A(n_562),
.Y(n_704)
);

NOR2xp33_ASAP7_75t_L g705 ( 
.A(n_545),
.B(n_5),
.Y(n_705)
);

NAND2xp5_ASAP7_75t_L g706 ( 
.A(n_529),
.B(n_203),
.Y(n_706)
);

INVx2_ASAP7_75t_L g707 ( 
.A(n_459),
.Y(n_707)
);

NOR2xp33_ASAP7_75t_L g708 ( 
.A(n_547),
.B(n_6),
.Y(n_708)
);

INVx3_ASAP7_75t_L g709 ( 
.A(n_529),
.Y(n_709)
);

NAND2xp5_ASAP7_75t_SL g710 ( 
.A(n_562),
.B(n_578),
.Y(n_710)
);

NOR3xp33_ASAP7_75t_L g711 ( 
.A(n_470),
.B(n_472),
.C(n_456),
.Y(n_711)
);

NAND2xp33_ASAP7_75t_L g712 ( 
.A(n_562),
.B(n_253),
.Y(n_712)
);

NAND2xp5_ASAP7_75t_L g713 ( 
.A(n_487),
.B(n_208),
.Y(n_713)
);

NOR2xp33_ASAP7_75t_L g714 ( 
.A(n_552),
.B(n_7),
.Y(n_714)
);

INVxp67_ASAP7_75t_L g715 ( 
.A(n_502),
.Y(n_715)
);

NAND2xp5_ASAP7_75t_SL g716 ( 
.A(n_562),
.B(n_578),
.Y(n_716)
);

BUFx6f_ASAP7_75t_SL g717 ( 
.A(n_508),
.Y(n_717)
);

INVx1_ASAP7_75t_L g718 ( 
.A(n_481),
.Y(n_718)
);

AOI221xp5_ASAP7_75t_L g719 ( 
.A1(n_530),
.A2(n_242),
.B1(n_209),
.B2(n_226),
.C(n_297),
.Y(n_719)
);

OR2x2_ASAP7_75t_L g720 ( 
.A(n_452),
.B(n_8),
.Y(n_720)
);

INVx2_ASAP7_75t_SL g721 ( 
.A(n_508),
.Y(n_721)
);

NOR2xp33_ASAP7_75t_L g722 ( 
.A(n_531),
.B(n_12),
.Y(n_722)
);

NOR2xp33_ASAP7_75t_L g723 ( 
.A(n_582),
.B(n_546),
.Y(n_723)
);

NAND2xp5_ASAP7_75t_L g724 ( 
.A(n_487),
.B(n_249),
.Y(n_724)
);

INVx2_ASAP7_75t_L g725 ( 
.A(n_516),
.Y(n_725)
);

BUFx3_ASAP7_75t_L g726 ( 
.A(n_586),
.Y(n_726)
);

NAND2xp5_ASAP7_75t_L g727 ( 
.A(n_492),
.B(n_243),
.Y(n_727)
);

BUFx8_ASAP7_75t_L g728 ( 
.A(n_537),
.Y(n_728)
);

NAND2xp5_ASAP7_75t_SL g729 ( 
.A(n_562),
.B(n_416),
.Y(n_729)
);

OAI22xp5_ASAP7_75t_L g730 ( 
.A1(n_520),
.A2(n_241),
.B1(n_228),
.B2(n_229),
.Y(n_730)
);

INVx3_ASAP7_75t_L g731 ( 
.A(n_492),
.Y(n_731)
);

CKINVDCx11_ASAP7_75t_R g732 ( 
.A(n_561),
.Y(n_732)
);

INVx1_ASAP7_75t_SL g733 ( 
.A(n_537),
.Y(n_733)
);

AOI22xp5_ASAP7_75t_L g734 ( 
.A1(n_520),
.A2(n_255),
.B1(n_236),
.B2(n_239),
.Y(n_734)
);

INVx2_ASAP7_75t_L g735 ( 
.A(n_516),
.Y(n_735)
);

NAND2xp5_ASAP7_75t_L g736 ( 
.A(n_511),
.B(n_292),
.Y(n_736)
);

NOR2xp33_ASAP7_75t_L g737 ( 
.A(n_565),
.B(n_13),
.Y(n_737)
);

NAND2xp5_ASAP7_75t_SL g738 ( 
.A(n_578),
.B(n_416),
.Y(n_738)
);

NAND2xp5_ASAP7_75t_L g739 ( 
.A(n_511),
.B(n_410),
.Y(n_739)
);

INVx2_ASAP7_75t_L g740 ( 
.A(n_533),
.Y(n_740)
);

NAND2xp5_ASAP7_75t_SL g741 ( 
.A(n_578),
.B(n_416),
.Y(n_741)
);

AOI22xp33_ASAP7_75t_L g742 ( 
.A1(n_503),
.A2(n_416),
.B1(n_410),
.B2(n_399),
.Y(n_742)
);

NAND2xp5_ASAP7_75t_SL g743 ( 
.A(n_578),
.B(n_416),
.Y(n_743)
);

NOR2xp33_ASAP7_75t_L g744 ( 
.A(n_580),
.B(n_13),
.Y(n_744)
);

BUFx6f_ASAP7_75t_L g745 ( 
.A(n_474),
.Y(n_745)
);

A2O1A1Ixp33_ASAP7_75t_L g746 ( 
.A1(n_566),
.A2(n_416),
.B(n_410),
.C(n_399),
.Y(n_746)
);

INVx1_ASAP7_75t_L g747 ( 
.A(n_481),
.Y(n_747)
);

NAND2xp5_ASAP7_75t_L g748 ( 
.A(n_513),
.B(n_416),
.Y(n_748)
);

OR2x2_ASAP7_75t_L g749 ( 
.A(n_449),
.B(n_16),
.Y(n_749)
);

INVx1_ASAP7_75t_L g750 ( 
.A(n_484),
.Y(n_750)
);

BUFx6f_ASAP7_75t_L g751 ( 
.A(n_474),
.Y(n_751)
);

OR2x6_ASAP7_75t_L g752 ( 
.A(n_467),
.B(n_283),
.Y(n_752)
);

NAND2xp5_ASAP7_75t_L g753 ( 
.A(n_513),
.B(n_410),
.Y(n_753)
);

BUFx4f_ASAP7_75t_L g754 ( 
.A(n_503),
.Y(n_754)
);

OR2x2_ASAP7_75t_L g755 ( 
.A(n_535),
.B(n_17),
.Y(n_755)
);

AND2x2_ASAP7_75t_L g756 ( 
.A(n_508),
.B(n_18),
.Y(n_756)
);

AOI22xp5_ASAP7_75t_L g757 ( 
.A1(n_581),
.A2(n_416),
.B1(n_410),
.B2(n_399),
.Y(n_757)
);

NAND2xp5_ASAP7_75t_L g758 ( 
.A(n_554),
.B(n_410),
.Y(n_758)
);

NOR2xp33_ASAP7_75t_L g759 ( 
.A(n_450),
.B(n_19),
.Y(n_759)
);

OR2x2_ASAP7_75t_L g760 ( 
.A(n_591),
.B(n_22),
.Y(n_760)
);

INVx1_ASAP7_75t_L g761 ( 
.A(n_623),
.Y(n_761)
);

INVx2_ASAP7_75t_L g762 ( 
.A(n_604),
.Y(n_762)
);

OAI21xp5_ASAP7_75t_L g763 ( 
.A1(n_640),
.A2(n_454),
.B(n_484),
.Y(n_763)
);

AOI21xp5_ASAP7_75t_L g764 ( 
.A1(n_598),
.A2(n_468),
.B(n_555),
.Y(n_764)
);

NAND2xp5_ASAP7_75t_L g765 ( 
.A(n_608),
.B(n_536),
.Y(n_765)
);

NAND2xp5_ASAP7_75t_SL g766 ( 
.A(n_667),
.B(n_450),
.Y(n_766)
);

OR2x2_ASAP7_75t_SL g767 ( 
.A(n_720),
.B(n_501),
.Y(n_767)
);

AOI21xp5_ASAP7_75t_L g768 ( 
.A1(n_710),
.A2(n_716),
.B(n_594),
.Y(n_768)
);

AOI21xp5_ASAP7_75t_L g769 ( 
.A1(n_710),
.A2(n_555),
.B(n_468),
.Y(n_769)
);

NOR3xp33_ASAP7_75t_L g770 ( 
.A(n_683),
.B(n_557),
.C(n_577),
.Y(n_770)
);

INVx1_ASAP7_75t_L g771 ( 
.A(n_661),
.Y(n_771)
);

AOI21xp5_ASAP7_75t_L g772 ( 
.A1(n_716),
.A2(n_468),
.B(n_583),
.Y(n_772)
);

AOI21xp5_ASAP7_75t_L g773 ( 
.A1(n_594),
.A2(n_522),
.B(n_583),
.Y(n_773)
);

NAND2xp5_ASAP7_75t_L g774 ( 
.A(n_608),
.B(n_471),
.Y(n_774)
);

AOI22xp5_ASAP7_75t_L g775 ( 
.A1(n_689),
.A2(n_503),
.B1(n_507),
.B2(n_505),
.Y(n_775)
);

AOI21xp5_ASAP7_75t_L g776 ( 
.A1(n_599),
.A2(n_522),
.B(n_583),
.Y(n_776)
);

NOR2xp33_ASAP7_75t_SL g777 ( 
.A(n_633),
.B(n_508),
.Y(n_777)
);

AOI21xp5_ASAP7_75t_L g778 ( 
.A1(n_599),
.A2(n_555),
.B(n_538),
.Y(n_778)
);

AOI21xp5_ASAP7_75t_L g779 ( 
.A1(n_600),
.A2(n_500),
.B(n_519),
.Y(n_779)
);

NAND2xp5_ASAP7_75t_L g780 ( 
.A(n_606),
.B(n_454),
.Y(n_780)
);

INVx1_ASAP7_75t_L g781 ( 
.A(n_664),
.Y(n_781)
);

NAND2xp5_ASAP7_75t_L g782 ( 
.A(n_606),
.B(n_544),
.Y(n_782)
);

BUFx4f_ASAP7_75t_L g783 ( 
.A(n_665),
.Y(n_783)
);

NAND2xp5_ASAP7_75t_L g784 ( 
.A(n_615),
.B(n_544),
.Y(n_784)
);

OAI21xp33_ASAP7_75t_L g785 ( 
.A1(n_682),
.A2(n_505),
.B(n_498),
.Y(n_785)
);

NAND2xp5_ASAP7_75t_L g786 ( 
.A(n_592),
.B(n_560),
.Y(n_786)
);

NOR2xp67_ASAP7_75t_L g787 ( 
.A(n_593),
.B(n_590),
.Y(n_787)
);

NOR2xp33_ASAP7_75t_L g788 ( 
.A(n_693),
.B(n_500),
.Y(n_788)
);

AOI21xp5_ASAP7_75t_L g789 ( 
.A1(n_600),
.A2(n_538),
.B(n_522),
.Y(n_789)
);

NAND2xp5_ASAP7_75t_L g790 ( 
.A(n_602),
.B(n_560),
.Y(n_790)
);

INVx2_ASAP7_75t_SL g791 ( 
.A(n_607),
.Y(n_791)
);

NAND2xp5_ASAP7_75t_SL g792 ( 
.A(n_667),
.B(n_500),
.Y(n_792)
);

OAI321xp33_ASAP7_75t_L g793 ( 
.A1(n_670),
.A2(n_590),
.A3(n_567),
.B1(n_588),
.B2(n_574),
.C(n_584),
.Y(n_793)
);

NAND2xp5_ASAP7_75t_L g794 ( 
.A(n_602),
.B(n_567),
.Y(n_794)
);

NAND2xp5_ASAP7_75t_SL g795 ( 
.A(n_709),
.B(n_519),
.Y(n_795)
);

INVx1_ASAP7_75t_L g796 ( 
.A(n_675),
.Y(n_796)
);

NAND2xp5_ASAP7_75t_L g797 ( 
.A(n_649),
.B(n_650),
.Y(n_797)
);

INVx2_ASAP7_75t_L g798 ( 
.A(n_605),
.Y(n_798)
);

NAND2xp5_ASAP7_75t_L g799 ( 
.A(n_595),
.B(n_574),
.Y(n_799)
);

INVx1_ASAP7_75t_L g800 ( 
.A(n_691),
.Y(n_800)
);

AO21x1_ASAP7_75t_L g801 ( 
.A1(n_737),
.A2(n_507),
.B(n_499),
.Y(n_801)
);

AOI21xp5_ASAP7_75t_L g802 ( 
.A1(n_603),
.A2(n_538),
.B(n_519),
.Y(n_802)
);

NOR2xp33_ASAP7_75t_L g803 ( 
.A(n_654),
.B(n_474),
.Y(n_803)
);

AOI21x1_ASAP7_75t_L g804 ( 
.A1(n_617),
.A2(n_498),
.B(n_499),
.Y(n_804)
);

AO21x1_ASAP7_75t_L g805 ( 
.A1(n_737),
.A2(n_588),
.B(n_584),
.Y(n_805)
);

NOR3xp33_ASAP7_75t_L g806 ( 
.A(n_687),
.B(n_576),
.C(n_494),
.Y(n_806)
);

AND2x4_ASAP7_75t_L g807 ( 
.A(n_721),
.B(n_576),
.Y(n_807)
);

HB1xp67_ASAP7_75t_L g808 ( 
.A(n_665),
.Y(n_808)
);

NAND2xp5_ASAP7_75t_L g809 ( 
.A(n_614),
.B(n_589),
.Y(n_809)
);

AOI21xp5_ASAP7_75t_L g810 ( 
.A1(n_603),
.A2(n_534),
.B(n_476),
.Y(n_810)
);

CKINVDCx10_ASAP7_75t_R g811 ( 
.A(n_717),
.Y(n_811)
);

INVx1_ASAP7_75t_L g812 ( 
.A(n_718),
.Y(n_812)
);

BUFx6f_ASAP7_75t_L g813 ( 
.A(n_665),
.Y(n_813)
);

AOI21xp5_ASAP7_75t_L g814 ( 
.A1(n_601),
.A2(n_534),
.B(n_476),
.Y(n_814)
);

BUFx2_ASAP7_75t_L g815 ( 
.A(n_607),
.Y(n_815)
);

NAND2xp5_ASAP7_75t_L g816 ( 
.A(n_723),
.B(n_589),
.Y(n_816)
);

NAND2xp5_ASAP7_75t_L g817 ( 
.A(n_723),
.B(n_585),
.Y(n_817)
);

NOR2xp67_ASAP7_75t_L g818 ( 
.A(n_715),
.B(n_585),
.Y(n_818)
);

NAND2xp5_ASAP7_75t_L g819 ( 
.A(n_660),
.B(n_647),
.Y(n_819)
);

NOR2xp33_ASAP7_75t_L g820 ( 
.A(n_733),
.B(n_476),
.Y(n_820)
);

NOR2x2_ASAP7_75t_L g821 ( 
.A(n_752),
.B(n_579),
.Y(n_821)
);

INVx3_ASAP7_75t_L g822 ( 
.A(n_709),
.Y(n_822)
);

AOI21xp5_ASAP7_75t_L g823 ( 
.A1(n_704),
.A2(n_534),
.B(n_493),
.Y(n_823)
);

BUFx12f_ASAP7_75t_L g824 ( 
.A(n_732),
.Y(n_824)
);

AOI21xp5_ASAP7_75t_L g825 ( 
.A1(n_677),
.A2(n_493),
.B(n_573),
.Y(n_825)
);

INVx2_ASAP7_75t_L g826 ( 
.A(n_613),
.Y(n_826)
);

OAI21xp5_ASAP7_75t_L g827 ( 
.A1(n_746),
.A2(n_493),
.B(n_524),
.Y(n_827)
);

HB1xp67_ASAP7_75t_L g828 ( 
.A(n_726),
.Y(n_828)
);

AOI21xp5_ASAP7_75t_L g829 ( 
.A1(n_617),
.A2(n_524),
.B(n_573),
.Y(n_829)
);

NAND2xp5_ASAP7_75t_L g830 ( 
.A(n_620),
.B(n_579),
.Y(n_830)
);

BUFx12f_ASAP7_75t_L g831 ( 
.A(n_728),
.Y(n_831)
);

AOI21xp33_ASAP7_75t_L g832 ( 
.A1(n_673),
.A2(n_575),
.B(n_533),
.Y(n_832)
);

INVxp67_ASAP7_75t_L g833 ( 
.A(n_678),
.Y(n_833)
);

NAND2xp5_ASAP7_75t_L g834 ( 
.A(n_621),
.B(n_575),
.Y(n_834)
);

BUFx6f_ASAP7_75t_L g835 ( 
.A(n_696),
.Y(n_835)
);

BUFx2_ASAP7_75t_L g836 ( 
.A(n_637),
.Y(n_836)
);

INVx2_ASAP7_75t_L g837 ( 
.A(n_619),
.Y(n_837)
);

NAND2xp5_ASAP7_75t_L g838 ( 
.A(n_627),
.B(n_549),
.Y(n_838)
);

NAND2xp5_ASAP7_75t_L g839 ( 
.A(n_722),
.B(n_549),
.Y(n_839)
);

NAND2xp5_ASAP7_75t_L g840 ( 
.A(n_722),
.B(n_540),
.Y(n_840)
);

INVx1_ASAP7_75t_L g841 ( 
.A(n_747),
.Y(n_841)
);

INVx1_ASAP7_75t_L g842 ( 
.A(n_750),
.Y(n_842)
);

AOI22xp5_ASAP7_75t_L g843 ( 
.A1(n_711),
.A2(n_503),
.B1(n_524),
.B2(n_573),
.Y(n_843)
);

AOI21xp5_ASAP7_75t_L g844 ( 
.A1(n_626),
.A2(n_550),
.B(n_559),
.Y(n_844)
);

AOI21xp5_ASAP7_75t_L g845 ( 
.A1(n_626),
.A2(n_550),
.B(n_559),
.Y(n_845)
);

AOI21x1_ASAP7_75t_L g846 ( 
.A1(n_636),
.A2(n_657),
.B(n_641),
.Y(n_846)
);

CKINVDCx20_ASAP7_75t_R g847 ( 
.A(n_728),
.Y(n_847)
);

A2O1A1Ixp33_ASAP7_75t_L g848 ( 
.A1(n_705),
.A2(n_571),
.B(n_563),
.C(n_540),
.Y(n_848)
);

NAND2xp5_ASAP7_75t_L g849 ( 
.A(n_618),
.B(n_571),
.Y(n_849)
);

AOI21xp5_ASAP7_75t_L g850 ( 
.A1(n_636),
.A2(n_559),
.B(n_550),
.Y(n_850)
);

NAND2xp5_ASAP7_75t_L g851 ( 
.A(n_680),
.B(n_563),
.Y(n_851)
);

AOI21xp5_ASAP7_75t_L g852 ( 
.A1(n_641),
.A2(n_558),
.B(n_494),
.Y(n_852)
);

NAND2xp5_ASAP7_75t_SL g853 ( 
.A(n_754),
.B(n_541),
.Y(n_853)
);

NAND2xp5_ASAP7_75t_L g854 ( 
.A(n_609),
.B(n_541),
.Y(n_854)
);

NOR2x2_ASAP7_75t_L g855 ( 
.A(n_752),
.B(n_23),
.Y(n_855)
);

NAND2xp5_ASAP7_75t_L g856 ( 
.A(n_629),
.B(n_503),
.Y(n_856)
);

O2A1O1Ixp33_ASAP7_75t_SL g857 ( 
.A1(n_663),
.A2(n_503),
.B(n_558),
.C(n_25),
.Y(n_857)
);

OAI21xp5_ASAP7_75t_L g858 ( 
.A1(n_616),
.A2(n_410),
.B(n_399),
.Y(n_858)
);

OAI321xp33_ASAP7_75t_L g859 ( 
.A1(n_670),
.A2(n_399),
.A3(n_283),
.B1(n_216),
.B2(n_161),
.C(n_28),
.Y(n_859)
);

AOI21xp5_ASAP7_75t_L g860 ( 
.A1(n_657),
.A2(n_729),
.B(n_676),
.Y(n_860)
);

INVx2_ASAP7_75t_L g861 ( 
.A(n_631),
.Y(n_861)
);

AOI21x1_ASAP7_75t_L g862 ( 
.A1(n_676),
.A2(n_399),
.B(n_253),
.Y(n_862)
);

NAND2xp5_ASAP7_75t_L g863 ( 
.A(n_611),
.B(n_23),
.Y(n_863)
);

NAND2xp5_ASAP7_75t_L g864 ( 
.A(n_611),
.B(n_24),
.Y(n_864)
);

AOI21xp5_ASAP7_75t_L g865 ( 
.A1(n_729),
.A2(n_283),
.B(n_216),
.Y(n_865)
);

NAND2xp5_ASAP7_75t_L g866 ( 
.A(n_610),
.B(n_685),
.Y(n_866)
);

A2O1A1Ixp33_ASAP7_75t_L g867 ( 
.A1(n_705),
.A2(n_216),
.B(n_161),
.C(n_283),
.Y(n_867)
);

NAND2xp5_ASAP7_75t_SL g868 ( 
.A(n_754),
.B(n_253),
.Y(n_868)
);

AND2x4_ASAP7_75t_L g869 ( 
.A(n_658),
.B(n_25),
.Y(n_869)
);

BUFx4f_ASAP7_75t_L g870 ( 
.A(n_658),
.Y(n_870)
);

INVx2_ASAP7_75t_L g871 ( 
.A(n_634),
.Y(n_871)
);

INVx3_ASAP7_75t_L g872 ( 
.A(n_692),
.Y(n_872)
);

OAI21xp5_ASAP7_75t_L g873 ( 
.A1(n_616),
.A2(n_253),
.B(n_216),
.Y(n_873)
);

NAND2xp5_ASAP7_75t_L g874 ( 
.A(n_688),
.B(n_26),
.Y(n_874)
);

INVx1_ASAP7_75t_SL g875 ( 
.A(n_698),
.Y(n_875)
);

AOI21xp5_ASAP7_75t_L g876 ( 
.A1(n_738),
.A2(n_161),
.B(n_253),
.Y(n_876)
);

INVx1_ASAP7_75t_L g877 ( 
.A(n_639),
.Y(n_877)
);

NAND2xp5_ASAP7_75t_L g878 ( 
.A(n_756),
.B(n_26),
.Y(n_878)
);

AOI21xp5_ASAP7_75t_L g879 ( 
.A1(n_738),
.A2(n_161),
.B(n_253),
.Y(n_879)
);

O2A1O1Ixp33_ASAP7_75t_L g880 ( 
.A1(n_687),
.A2(n_30),
.B(n_35),
.C(n_36),
.Y(n_880)
);

INVx5_ASAP7_75t_L g881 ( 
.A(n_692),
.Y(n_881)
);

AOI21xp5_ASAP7_75t_L g882 ( 
.A1(n_741),
.A2(n_106),
.B(n_145),
.Y(n_882)
);

AOI21xp5_ASAP7_75t_L g883 ( 
.A1(n_741),
.A2(n_102),
.B(n_143),
.Y(n_883)
);

BUFx2_ASAP7_75t_L g884 ( 
.A(n_698),
.Y(n_884)
);

NAND2xp5_ASAP7_75t_L g885 ( 
.A(n_638),
.B(n_37),
.Y(n_885)
);

AOI21xp5_ASAP7_75t_L g886 ( 
.A1(n_743),
.A2(n_95),
.B(n_137),
.Y(n_886)
);

NAND2xp5_ASAP7_75t_L g887 ( 
.A(n_632),
.B(n_42),
.Y(n_887)
);

AOI21xp5_ASAP7_75t_L g888 ( 
.A1(n_743),
.A2(n_107),
.B(n_132),
.Y(n_888)
);

O2A1O1Ixp33_ASAP7_75t_L g889 ( 
.A1(n_760),
.A2(n_43),
.B(n_47),
.C(n_53),
.Y(n_889)
);

INVx2_ASAP7_75t_SL g890 ( 
.A(n_679),
.Y(n_890)
);

AOI22xp5_ASAP7_75t_L g891 ( 
.A1(n_653),
.A2(n_43),
.B1(n_69),
.B2(n_70),
.Y(n_891)
);

NAND2xp5_ASAP7_75t_SL g892 ( 
.A(n_745),
.B(n_80),
.Y(n_892)
);

NOR2xp67_ASAP7_75t_L g893 ( 
.A(n_734),
.B(n_87),
.Y(n_893)
);

NAND2xp5_ASAP7_75t_L g894 ( 
.A(n_673),
.B(n_88),
.Y(n_894)
);

NAND2xp5_ASAP7_75t_L g895 ( 
.A(n_708),
.B(n_94),
.Y(n_895)
);

AOI21xp5_ASAP7_75t_L g896 ( 
.A1(n_739),
.A2(n_748),
.B(n_753),
.Y(n_896)
);

INVx1_ASAP7_75t_L g897 ( 
.A(n_643),
.Y(n_897)
);

HB1xp67_ASAP7_75t_L g898 ( 
.A(n_666),
.Y(n_898)
);

AOI21xp5_ASAP7_75t_L g899 ( 
.A1(n_596),
.A2(n_108),
.B(n_115),
.Y(n_899)
);

HB1xp67_ASAP7_75t_L g900 ( 
.A(n_674),
.Y(n_900)
);

AOI21xp5_ASAP7_75t_L g901 ( 
.A1(n_758),
.A2(n_120),
.B(n_121),
.Y(n_901)
);

AOI21xp5_ASAP7_75t_L g902 ( 
.A1(n_652),
.A2(n_122),
.B(n_124),
.Y(n_902)
);

INVx1_ASAP7_75t_SL g903 ( 
.A(n_671),
.Y(n_903)
);

O2A1O1Ixp33_ASAP7_75t_L g904 ( 
.A1(n_749),
.A2(n_755),
.B(n_708),
.C(n_714),
.Y(n_904)
);

AOI21xp5_ASAP7_75t_L g905 ( 
.A1(n_652),
.A2(n_125),
.B(n_154),
.Y(n_905)
);

AOI21xp5_ASAP7_75t_L g906 ( 
.A1(n_695),
.A2(n_697),
.B(n_706),
.Y(n_906)
);

AOI21xp5_ASAP7_75t_L g907 ( 
.A1(n_700),
.A2(n_624),
.B(n_751),
.Y(n_907)
);

INVx1_ASAP7_75t_L g908 ( 
.A(n_648),
.Y(n_908)
);

AOI21xp5_ASAP7_75t_L g909 ( 
.A1(n_745),
.A2(n_751),
.B(n_731),
.Y(n_909)
);

OAI21xp33_ASAP7_75t_L g910 ( 
.A1(n_744),
.A2(n_714),
.B(n_622),
.Y(n_910)
);

AOI22xp33_ASAP7_75t_L g911 ( 
.A1(n_669),
.A2(n_690),
.B1(n_612),
.B2(n_701),
.Y(n_911)
);

NAND2xp5_ASAP7_75t_L g912 ( 
.A(n_644),
.B(n_744),
.Y(n_912)
);

OR2x2_ASAP7_75t_SL g913 ( 
.A(n_651),
.B(n_655),
.Y(n_913)
);

NAND2xp5_ASAP7_75t_L g914 ( 
.A(n_719),
.B(n_669),
.Y(n_914)
);

NAND2xp5_ASAP7_75t_L g915 ( 
.A(n_628),
.B(n_642),
.Y(n_915)
);

A2O1A1Ixp33_ASAP7_75t_L g916 ( 
.A1(n_759),
.A2(n_642),
.B(n_628),
.C(n_597),
.Y(n_916)
);

OAI21xp5_ASAP7_75t_L g917 ( 
.A1(n_757),
.A2(n_694),
.B(n_740),
.Y(n_917)
);

BUFx4f_ASAP7_75t_L g918 ( 
.A(n_752),
.Y(n_918)
);

HB1xp67_ASAP7_75t_L g919 ( 
.A(n_731),
.Y(n_919)
);

INVx1_ASAP7_75t_L g920 ( 
.A(n_659),
.Y(n_920)
);

OAI21xp5_ASAP7_75t_L g921 ( 
.A1(n_662),
.A2(n_707),
.B(n_686),
.Y(n_921)
);

NOR2xp33_ASAP7_75t_L g922 ( 
.A(n_656),
.B(n_630),
.Y(n_922)
);

AOI22xp5_ASAP7_75t_L g923 ( 
.A1(n_646),
.A2(n_690),
.B1(n_759),
.B2(n_702),
.Y(n_923)
);

AOI21xp5_ASAP7_75t_L g924 ( 
.A1(n_745),
.A2(n_751),
.B(n_736),
.Y(n_924)
);

NAND2xp5_ASAP7_75t_L g925 ( 
.A(n_612),
.B(n_735),
.Y(n_925)
);

AOI21xp5_ASAP7_75t_L g926 ( 
.A1(n_745),
.A2(n_751),
.B(n_727),
.Y(n_926)
);

NOR2xp33_ASAP7_75t_L g927 ( 
.A(n_717),
.B(n_730),
.Y(n_927)
);

AND2x2_ASAP7_75t_L g928 ( 
.A(n_684),
.B(n_725),
.Y(n_928)
);

AOI21xp5_ASAP7_75t_L g929 ( 
.A1(n_713),
.A2(n_724),
.B(n_696),
.Y(n_929)
);

NAND2xp5_ASAP7_75t_SL g930 ( 
.A(n_696),
.B(n_703),
.Y(n_930)
);

INVx3_ASAP7_75t_L g931 ( 
.A(n_692),
.Y(n_931)
);

NOR2xp33_ASAP7_75t_L g932 ( 
.A(n_635),
.B(n_645),
.Y(n_932)
);

NAND2xp5_ASAP7_75t_L g933 ( 
.A(n_696),
.B(n_703),
.Y(n_933)
);

NAND2xp5_ASAP7_75t_L g934 ( 
.A(n_703),
.B(n_625),
.Y(n_934)
);

HB1xp67_ASAP7_75t_L g935 ( 
.A(n_703),
.Y(n_935)
);

NAND2xp5_ASAP7_75t_L g936 ( 
.A(n_742),
.B(n_668),
.Y(n_936)
);

INVxp67_ASAP7_75t_SL g937 ( 
.A(n_742),
.Y(n_937)
);

NOR2xp33_ASAP7_75t_L g938 ( 
.A(n_681),
.B(n_712),
.Y(n_938)
);

NAND2xp5_ASAP7_75t_SL g939 ( 
.A(n_672),
.B(n_699),
.Y(n_939)
);

NAND2xp5_ASAP7_75t_L g940 ( 
.A(n_608),
.B(n_594),
.Y(n_940)
);

NAND2xp5_ASAP7_75t_L g941 ( 
.A(n_608),
.B(n_594),
.Y(n_941)
);

INVx1_ASAP7_75t_L g942 ( 
.A(n_623),
.Y(n_942)
);

AOI21xp5_ASAP7_75t_L g943 ( 
.A1(n_598),
.A2(n_716),
.B(n_710),
.Y(n_943)
);

NOR2xp33_ASAP7_75t_L g944 ( 
.A(n_683),
.B(n_689),
.Y(n_944)
);

AOI21xp5_ASAP7_75t_L g945 ( 
.A1(n_598),
.A2(n_716),
.B(n_710),
.Y(n_945)
);

INVx2_ASAP7_75t_L g946 ( 
.A(n_762),
.Y(n_946)
);

CKINVDCx8_ASAP7_75t_R g947 ( 
.A(n_811),
.Y(n_947)
);

OR2x6_ASAP7_75t_L g948 ( 
.A(n_813),
.B(n_791),
.Y(n_948)
);

AND2x2_ASAP7_75t_L g949 ( 
.A(n_944),
.B(n_903),
.Y(n_949)
);

OAI22xp5_ASAP7_75t_L g950 ( 
.A1(n_940),
.A2(n_941),
.B1(n_797),
.B2(n_910),
.Y(n_950)
);

NAND2xp5_ASAP7_75t_L g951 ( 
.A(n_944),
.B(n_774),
.Y(n_951)
);

OAI22x1_ASAP7_75t_L g952 ( 
.A1(n_891),
.A2(n_914),
.B1(n_923),
.B2(n_927),
.Y(n_952)
);

INVx5_ASAP7_75t_L g953 ( 
.A(n_813),
.Y(n_953)
);

NOR2xp33_ASAP7_75t_L g954 ( 
.A(n_875),
.B(n_777),
.Y(n_954)
);

NOR2xp33_ASAP7_75t_SL g955 ( 
.A(n_831),
.B(n_847),
.Y(n_955)
);

NAND2xp5_ASAP7_75t_SL g956 ( 
.A(n_918),
.B(n_833),
.Y(n_956)
);

AND2x2_ASAP7_75t_L g957 ( 
.A(n_884),
.B(n_890),
.Y(n_957)
);

INVx2_ASAP7_75t_L g958 ( 
.A(n_798),
.Y(n_958)
);

AOI22xp33_ASAP7_75t_SL g959 ( 
.A1(n_765),
.A2(n_937),
.B1(n_887),
.B2(n_767),
.Y(n_959)
);

A2O1A1Ixp33_ASAP7_75t_L g960 ( 
.A1(n_904),
.A2(n_916),
.B(n_770),
.C(n_895),
.Y(n_960)
);

BUFx12f_ASAP7_75t_L g961 ( 
.A(n_824),
.Y(n_961)
);

INVx1_ASAP7_75t_L g962 ( 
.A(n_761),
.Y(n_962)
);

BUFx2_ASAP7_75t_L g963 ( 
.A(n_836),
.Y(n_963)
);

OA22x2_ASAP7_75t_L g964 ( 
.A1(n_828),
.A2(n_866),
.B1(n_819),
.B2(n_878),
.Y(n_964)
);

NAND2xp5_ASAP7_75t_SL g965 ( 
.A(n_918),
.B(n_788),
.Y(n_965)
);

A2O1A1Ixp33_ASAP7_75t_SL g966 ( 
.A1(n_770),
.A2(n_803),
.B(n_912),
.C(n_906),
.Y(n_966)
);

HB1xp67_ASAP7_75t_L g967 ( 
.A(n_898),
.Y(n_967)
);

AND2x4_ASAP7_75t_L g968 ( 
.A(n_808),
.B(n_813),
.Y(n_968)
);

INVx2_ASAP7_75t_L g969 ( 
.A(n_826),
.Y(n_969)
);

AOI21xp5_ASAP7_75t_L g970 ( 
.A1(n_780),
.A2(n_782),
.B(n_768),
.Y(n_970)
);

INVx1_ASAP7_75t_L g971 ( 
.A(n_771),
.Y(n_971)
);

AOI22xp5_ASAP7_75t_L g972 ( 
.A1(n_911),
.A2(n_820),
.B1(n_927),
.B2(n_788),
.Y(n_972)
);

NOR2xp33_ASAP7_75t_L g973 ( 
.A(n_898),
.B(n_900),
.Y(n_973)
);

NAND2xp5_ASAP7_75t_L g974 ( 
.A(n_900),
.B(n_786),
.Y(n_974)
);

INVx4_ASAP7_75t_L g975 ( 
.A(n_813),
.Y(n_975)
);

OAI22xp5_ASAP7_75t_L g976 ( 
.A1(n_911),
.A2(n_784),
.B1(n_785),
.B2(n_822),
.Y(n_976)
);

OAI22xp5_ASAP7_75t_SL g977 ( 
.A1(n_913),
.A2(n_815),
.B1(n_922),
.B2(n_828),
.Y(n_977)
);

AOI21xp5_ASAP7_75t_L g978 ( 
.A1(n_907),
.A2(n_945),
.B(n_943),
.Y(n_978)
);

NAND2xp5_ASAP7_75t_L g979 ( 
.A(n_820),
.B(n_877),
.Y(n_979)
);

NOR2xp33_ASAP7_75t_L g980 ( 
.A(n_922),
.B(n_808),
.Y(n_980)
);

NOR2xp33_ASAP7_75t_L g981 ( 
.A(n_897),
.B(n_781),
.Y(n_981)
);

BUFx3_ASAP7_75t_L g982 ( 
.A(n_783),
.Y(n_982)
);

NOR2xp33_ASAP7_75t_SL g983 ( 
.A(n_783),
.B(n_870),
.Y(n_983)
);

INVx2_ASAP7_75t_L g984 ( 
.A(n_837),
.Y(n_984)
);

BUFx12f_ASAP7_75t_L g985 ( 
.A(n_869),
.Y(n_985)
);

INVx2_ASAP7_75t_L g986 ( 
.A(n_861),
.Y(n_986)
);

BUFx6f_ASAP7_75t_L g987 ( 
.A(n_835),
.Y(n_987)
);

AOI21xp5_ASAP7_75t_L g988 ( 
.A1(n_773),
.A2(n_929),
.B(n_915),
.Y(n_988)
);

INVx1_ASAP7_75t_L g989 ( 
.A(n_796),
.Y(n_989)
);

AOI21xp5_ASAP7_75t_L g990 ( 
.A1(n_896),
.A2(n_851),
.B(n_814),
.Y(n_990)
);

OAI21xp5_ASAP7_75t_L g991 ( 
.A1(n_803),
.A2(n_856),
.B(n_860),
.Y(n_991)
);

O2A1O1Ixp5_ASAP7_75t_L g992 ( 
.A1(n_801),
.A2(n_939),
.B(n_805),
.C(n_864),
.Y(n_992)
);

INVx1_ASAP7_75t_L g993 ( 
.A(n_800),
.Y(n_993)
);

NOR2xp67_ASAP7_75t_SL g994 ( 
.A(n_859),
.B(n_881),
.Y(n_994)
);

BUFx6f_ASAP7_75t_L g995 ( 
.A(n_835),
.Y(n_995)
);

O2A1O1Ixp33_ASAP7_75t_L g996 ( 
.A1(n_880),
.A2(n_889),
.B(n_863),
.C(n_874),
.Y(n_996)
);

NAND2xp5_ASAP7_75t_SL g997 ( 
.A(n_822),
.B(n_793),
.Y(n_997)
);

INVxp67_ASAP7_75t_L g998 ( 
.A(n_919),
.Y(n_998)
);

AOI33xp33_ASAP7_75t_L g999 ( 
.A1(n_812),
.A2(n_942),
.A3(n_841),
.B1(n_842),
.B2(n_869),
.B3(n_857),
.Y(n_999)
);

A2O1A1Ixp33_ASAP7_75t_L g1000 ( 
.A1(n_894),
.A2(n_893),
.B(n_873),
.C(n_806),
.Y(n_1000)
);

INVx1_ASAP7_75t_L g1001 ( 
.A(n_908),
.Y(n_1001)
);

BUFx2_ASAP7_75t_L g1002 ( 
.A(n_855),
.Y(n_1002)
);

AOI21xp5_ASAP7_75t_L g1003 ( 
.A1(n_849),
.A2(n_764),
.B(n_838),
.Y(n_1003)
);

AOI21xp5_ASAP7_75t_L g1004 ( 
.A1(n_830),
.A2(n_834),
.B(n_825),
.Y(n_1004)
);

NAND2xp5_ASAP7_75t_L g1005 ( 
.A(n_790),
.B(n_794),
.Y(n_1005)
);

INVx2_ASAP7_75t_L g1006 ( 
.A(n_871),
.Y(n_1006)
);

NAND2xp5_ASAP7_75t_L g1007 ( 
.A(n_807),
.B(n_925),
.Y(n_1007)
);

OAI21x1_ASAP7_75t_L g1008 ( 
.A1(n_862),
.A2(n_804),
.B(n_763),
.Y(n_1008)
);

NAND2xp5_ASAP7_75t_L g1009 ( 
.A(n_807),
.B(n_787),
.Y(n_1009)
);

AOI21xp5_ASAP7_75t_L g1010 ( 
.A1(n_839),
.A2(n_840),
.B(n_858),
.Y(n_1010)
);

OAI22xp5_ASAP7_75t_L g1011 ( 
.A1(n_775),
.A2(n_937),
.B1(n_809),
.B2(n_799),
.Y(n_1011)
);

AOI21xp5_ASAP7_75t_L g1012 ( 
.A1(n_776),
.A2(n_802),
.B(n_789),
.Y(n_1012)
);

INVx3_ASAP7_75t_L g1013 ( 
.A(n_881),
.Y(n_1013)
);

CKINVDCx5p33_ASAP7_75t_R g1014 ( 
.A(n_935),
.Y(n_1014)
);

INVx2_ASAP7_75t_L g1015 ( 
.A(n_928),
.Y(n_1015)
);

NOR2xp33_ASAP7_75t_L g1016 ( 
.A(n_816),
.B(n_817),
.Y(n_1016)
);

AOI21xp5_ASAP7_75t_L g1017 ( 
.A1(n_778),
.A2(n_779),
.B(n_924),
.Y(n_1017)
);

BUFx3_ASAP7_75t_L g1018 ( 
.A(n_835),
.Y(n_1018)
);

NAND3xp33_ASAP7_75t_L g1019 ( 
.A(n_806),
.B(n_885),
.C(n_843),
.Y(n_1019)
);

NOR3xp33_ASAP7_75t_SL g1020 ( 
.A(n_939),
.B(n_795),
.C(n_899),
.Y(n_1020)
);

INVx1_ASAP7_75t_SL g1021 ( 
.A(n_821),
.Y(n_1021)
);

AND2x2_ASAP7_75t_L g1022 ( 
.A(n_818),
.B(n_920),
.Y(n_1022)
);

BUFx4f_ASAP7_75t_L g1023 ( 
.A(n_835),
.Y(n_1023)
);

AOI21xp5_ASAP7_75t_L g1024 ( 
.A1(n_926),
.A2(n_769),
.B(n_772),
.Y(n_1024)
);

AOI22xp5_ASAP7_75t_L g1025 ( 
.A1(n_934),
.A2(n_854),
.B1(n_792),
.B2(n_766),
.Y(n_1025)
);

OAI22xp33_ASAP7_75t_L g1026 ( 
.A1(n_936),
.A2(n_881),
.B1(n_935),
.B2(n_905),
.Y(n_1026)
);

INVx2_ASAP7_75t_L g1027 ( 
.A(n_846),
.Y(n_1027)
);

INVxp67_ASAP7_75t_SL g1028 ( 
.A(n_933),
.Y(n_1028)
);

BUFx4f_ASAP7_75t_L g1029 ( 
.A(n_872),
.Y(n_1029)
);

AND2x4_ASAP7_75t_L g1030 ( 
.A(n_872),
.B(n_931),
.Y(n_1030)
);

NOR2xp33_ASAP7_75t_L g1031 ( 
.A(n_795),
.B(n_932),
.Y(n_1031)
);

INVx1_ASAP7_75t_L g1032 ( 
.A(n_921),
.Y(n_1032)
);

INVx2_ASAP7_75t_L g1033 ( 
.A(n_930),
.Y(n_1033)
);

AOI21xp5_ASAP7_75t_L g1034 ( 
.A1(n_810),
.A2(n_827),
.B(n_845),
.Y(n_1034)
);

INVx1_ASAP7_75t_L g1035 ( 
.A(n_848),
.Y(n_1035)
);

OAI22xp5_ASAP7_75t_L g1036 ( 
.A1(n_938),
.A2(n_931),
.B1(n_792),
.B2(n_766),
.Y(n_1036)
);

NAND2xp5_ASAP7_75t_L g1037 ( 
.A(n_909),
.B(n_832),
.Y(n_1037)
);

BUFx8_ASAP7_75t_L g1038 ( 
.A(n_930),
.Y(n_1038)
);

HB1xp67_ASAP7_75t_L g1039 ( 
.A(n_853),
.Y(n_1039)
);

NAND2xp5_ASAP7_75t_L g1040 ( 
.A(n_938),
.B(n_853),
.Y(n_1040)
);

OAI22xp5_ASAP7_75t_L g1041 ( 
.A1(n_829),
.A2(n_844),
.B1(n_850),
.B2(n_823),
.Y(n_1041)
);

OA21x2_ASAP7_75t_L g1042 ( 
.A1(n_917),
.A2(n_867),
.B(n_876),
.Y(n_1042)
);

NAND2xp5_ASAP7_75t_L g1043 ( 
.A(n_868),
.B(n_852),
.Y(n_1043)
);

BUFx4f_ASAP7_75t_L g1044 ( 
.A(n_892),
.Y(n_1044)
);

AOI21xp5_ASAP7_75t_L g1045 ( 
.A1(n_868),
.A2(n_901),
.B(n_902),
.Y(n_1045)
);

INVx2_ASAP7_75t_L g1046 ( 
.A(n_892),
.Y(n_1046)
);

AND2x2_ASAP7_75t_L g1047 ( 
.A(n_879),
.B(n_865),
.Y(n_1047)
);

OAI22xp5_ASAP7_75t_L g1048 ( 
.A1(n_882),
.A2(n_883),
.B1(n_886),
.B2(n_888),
.Y(n_1048)
);

AOI21xp5_ASAP7_75t_L g1049 ( 
.A1(n_940),
.A2(n_941),
.B(n_906),
.Y(n_1049)
);

OAI22xp5_ASAP7_75t_L g1050 ( 
.A1(n_940),
.A2(n_941),
.B1(n_797),
.B2(n_594),
.Y(n_1050)
);

BUFx12f_ASAP7_75t_L g1051 ( 
.A(n_831),
.Y(n_1051)
);

AOI22xp5_ASAP7_75t_L g1052 ( 
.A1(n_940),
.A2(n_941),
.B1(n_564),
.B2(n_478),
.Y(n_1052)
);

OR2x6_ASAP7_75t_L g1053 ( 
.A(n_813),
.B(n_665),
.Y(n_1053)
);

BUFx12f_ASAP7_75t_L g1054 ( 
.A(n_831),
.Y(n_1054)
);

NAND2xp5_ASAP7_75t_SL g1055 ( 
.A(n_944),
.B(n_593),
.Y(n_1055)
);

HB1xp67_ASAP7_75t_L g1056 ( 
.A(n_898),
.Y(n_1056)
);

AND2x2_ASAP7_75t_L g1057 ( 
.A(n_944),
.B(n_733),
.Y(n_1057)
);

OAI21x1_ASAP7_75t_L g1058 ( 
.A1(n_862),
.A2(n_896),
.B(n_943),
.Y(n_1058)
);

OAI21x1_ASAP7_75t_L g1059 ( 
.A1(n_862),
.A2(n_896),
.B(n_943),
.Y(n_1059)
);

AOI22xp33_ASAP7_75t_L g1060 ( 
.A1(n_914),
.A2(n_911),
.B1(n_669),
.B2(n_910),
.Y(n_1060)
);

NAND3xp33_ASAP7_75t_SL g1061 ( 
.A(n_940),
.B(n_941),
.C(n_910),
.Y(n_1061)
);

AND2x4_ASAP7_75t_L g1062 ( 
.A(n_808),
.B(n_813),
.Y(n_1062)
);

OAI22xp5_ASAP7_75t_L g1063 ( 
.A1(n_940),
.A2(n_941),
.B1(n_797),
.B2(n_594),
.Y(n_1063)
);

OR2x2_ASAP7_75t_L g1064 ( 
.A(n_903),
.B(n_496),
.Y(n_1064)
);

NOR2xp67_ASAP7_75t_SL g1065 ( 
.A(n_836),
.B(n_451),
.Y(n_1065)
);

OAI22xp5_ASAP7_75t_L g1066 ( 
.A1(n_940),
.A2(n_941),
.B1(n_797),
.B2(n_594),
.Y(n_1066)
);

NAND2xp5_ASAP7_75t_L g1067 ( 
.A(n_940),
.B(n_941),
.Y(n_1067)
);

INVx2_ASAP7_75t_L g1068 ( 
.A(n_762),
.Y(n_1068)
);

BUFx3_ASAP7_75t_L g1069 ( 
.A(n_836),
.Y(n_1069)
);

BUFx2_ASAP7_75t_L g1070 ( 
.A(n_884),
.Y(n_1070)
);

BUFx6f_ASAP7_75t_L g1071 ( 
.A(n_813),
.Y(n_1071)
);

NAND2xp33_ASAP7_75t_SL g1072 ( 
.A(n_940),
.B(n_941),
.Y(n_1072)
);

NOR2xp33_ASAP7_75t_SL g1073 ( 
.A(n_831),
.B(n_496),
.Y(n_1073)
);

AOI21xp5_ASAP7_75t_L g1074 ( 
.A1(n_940),
.A2(n_941),
.B(n_906),
.Y(n_1074)
);

INVx1_ASAP7_75t_L g1075 ( 
.A(n_761),
.Y(n_1075)
);

INVx2_ASAP7_75t_L g1076 ( 
.A(n_762),
.Y(n_1076)
);

OAI22xp5_ASAP7_75t_L g1077 ( 
.A1(n_940),
.A2(n_941),
.B1(n_797),
.B2(n_594),
.Y(n_1077)
);

AOI21xp5_ASAP7_75t_L g1078 ( 
.A1(n_940),
.A2(n_941),
.B(n_906),
.Y(n_1078)
);

NAND2xp5_ASAP7_75t_L g1079 ( 
.A(n_940),
.B(n_941),
.Y(n_1079)
);

AOI21xp5_ASAP7_75t_L g1080 ( 
.A1(n_940),
.A2(n_941),
.B(n_906),
.Y(n_1080)
);

BUFx6f_ASAP7_75t_L g1081 ( 
.A(n_813),
.Y(n_1081)
);

BUFx12f_ASAP7_75t_L g1082 ( 
.A(n_831),
.Y(n_1082)
);

AOI22xp33_ASAP7_75t_L g1083 ( 
.A1(n_914),
.A2(n_911),
.B1(n_669),
.B2(n_910),
.Y(n_1083)
);

NAND2xp5_ASAP7_75t_SL g1084 ( 
.A(n_944),
.B(n_593),
.Y(n_1084)
);

AND2x2_ASAP7_75t_L g1085 ( 
.A(n_944),
.B(n_733),
.Y(n_1085)
);

AND2x4_ASAP7_75t_L g1086 ( 
.A(n_808),
.B(n_813),
.Y(n_1086)
);

BUFx2_ASAP7_75t_L g1087 ( 
.A(n_884),
.Y(n_1087)
);

INVx3_ASAP7_75t_L g1088 ( 
.A(n_813),
.Y(n_1088)
);

OA21x2_ASAP7_75t_L g1089 ( 
.A1(n_992),
.A2(n_978),
.B(n_988),
.Y(n_1089)
);

O2A1O1Ixp33_ASAP7_75t_L g1090 ( 
.A1(n_960),
.A2(n_1063),
.B(n_1050),
.C(n_1077),
.Y(n_1090)
);

NAND2x1p5_ASAP7_75t_L g1091 ( 
.A(n_953),
.B(n_1023),
.Y(n_1091)
);

AO31x2_ASAP7_75t_L g1092 ( 
.A1(n_1000),
.A2(n_990),
.A3(n_1027),
.B(n_952),
.Y(n_1092)
);

OAI21x1_ASAP7_75t_L g1093 ( 
.A1(n_1012),
.A2(n_1059),
.B(n_1058),
.Y(n_1093)
);

A2O1A1Ixp33_ASAP7_75t_L g1094 ( 
.A1(n_1066),
.A2(n_996),
.B(n_1072),
.C(n_1052),
.Y(n_1094)
);

OAI21x1_ASAP7_75t_L g1095 ( 
.A1(n_1012),
.A2(n_1024),
.B(n_1017),
.Y(n_1095)
);

AOI21x1_ASAP7_75t_L g1096 ( 
.A1(n_970),
.A2(n_1034),
.B(n_1024),
.Y(n_1096)
);

NOR2xp33_ASAP7_75t_SL g1097 ( 
.A(n_994),
.B(n_985),
.Y(n_1097)
);

CKINVDCx16_ASAP7_75t_R g1098 ( 
.A(n_955),
.Y(n_1098)
);

OA21x2_ASAP7_75t_L g1099 ( 
.A1(n_992),
.A2(n_978),
.B(n_988),
.Y(n_1099)
);

AOI21xp5_ASAP7_75t_L g1100 ( 
.A1(n_1049),
.A2(n_1080),
.B(n_1078),
.Y(n_1100)
);

O2A1O1Ixp33_ASAP7_75t_L g1101 ( 
.A1(n_950),
.A2(n_1061),
.B(n_1067),
.C(n_1079),
.Y(n_1101)
);

NOR2xp67_ASAP7_75t_L g1102 ( 
.A(n_1064),
.B(n_954),
.Y(n_1102)
);

OAI21x1_ASAP7_75t_L g1103 ( 
.A1(n_1017),
.A2(n_1034),
.B(n_1008),
.Y(n_1103)
);

AOI21xp5_ASAP7_75t_L g1104 ( 
.A1(n_1049),
.A2(n_1078),
.B(n_1074),
.Y(n_1104)
);

O2A1O1Ixp33_ASAP7_75t_L g1105 ( 
.A1(n_1061),
.A2(n_951),
.B(n_996),
.C(n_966),
.Y(n_1105)
);

AND2x2_ASAP7_75t_L g1106 ( 
.A(n_1057),
.B(n_1085),
.Y(n_1106)
);

OAI22xp5_ASAP7_75t_L g1107 ( 
.A1(n_1060),
.A2(n_1083),
.B1(n_972),
.B2(n_1016),
.Y(n_1107)
);

AOI21xp5_ASAP7_75t_L g1108 ( 
.A1(n_1074),
.A2(n_1080),
.B(n_970),
.Y(n_1108)
);

AO31x2_ASAP7_75t_L g1109 ( 
.A1(n_990),
.A2(n_1041),
.A3(n_1004),
.B(n_1037),
.Y(n_1109)
);

BUFx3_ASAP7_75t_L g1110 ( 
.A(n_1069),
.Y(n_1110)
);

NAND2xp5_ASAP7_75t_L g1111 ( 
.A(n_1016),
.B(n_1060),
.Y(n_1111)
);

AOI21xp5_ASAP7_75t_L g1112 ( 
.A1(n_1026),
.A2(n_1003),
.B(n_1004),
.Y(n_1112)
);

OAI22xp5_ASAP7_75t_L g1113 ( 
.A1(n_1083),
.A2(n_959),
.B1(n_1019),
.B2(n_1044),
.Y(n_1113)
);

INVx2_ASAP7_75t_L g1114 ( 
.A(n_1015),
.Y(n_1114)
);

BUFx2_ASAP7_75t_L g1115 ( 
.A(n_963),
.Y(n_1115)
);

NAND2xp5_ASAP7_75t_L g1116 ( 
.A(n_949),
.B(n_973),
.Y(n_1116)
);

INVx1_ASAP7_75t_L g1117 ( 
.A(n_962),
.Y(n_1117)
);

NAND3xp33_ASAP7_75t_L g1118 ( 
.A(n_959),
.B(n_999),
.C(n_1020),
.Y(n_1118)
);

OAI21xp5_ASAP7_75t_L g1119 ( 
.A1(n_1010),
.A2(n_991),
.B(n_1011),
.Y(n_1119)
);

OAI21x1_ASAP7_75t_L g1120 ( 
.A1(n_1045),
.A2(n_1003),
.B(n_1043),
.Y(n_1120)
);

INVx1_ASAP7_75t_L g1121 ( 
.A(n_971),
.Y(n_1121)
);

CKINVDCx11_ASAP7_75t_R g1122 ( 
.A(n_947),
.Y(n_1122)
);

OAI21xp5_ASAP7_75t_L g1123 ( 
.A1(n_1010),
.A2(n_997),
.B(n_976),
.Y(n_1123)
);

NAND2xp5_ASAP7_75t_L g1124 ( 
.A(n_973),
.B(n_967),
.Y(n_1124)
);

NAND3xp33_ASAP7_75t_L g1125 ( 
.A(n_1020),
.B(n_1031),
.C(n_1025),
.Y(n_1125)
);

CKINVDCx20_ASAP7_75t_R g1126 ( 
.A(n_961),
.Y(n_1126)
);

CKINVDCx20_ASAP7_75t_R g1127 ( 
.A(n_1051),
.Y(n_1127)
);

INVx3_ASAP7_75t_L g1128 ( 
.A(n_1023),
.Y(n_1128)
);

INVx3_ASAP7_75t_L g1129 ( 
.A(n_1029),
.Y(n_1129)
);

OAI21xp5_ASAP7_75t_L g1130 ( 
.A1(n_1044),
.A2(n_1040),
.B(n_1035),
.Y(n_1130)
);

OAI21x1_ASAP7_75t_L g1131 ( 
.A1(n_1045),
.A2(n_1048),
.B(n_1047),
.Y(n_1131)
);

AO21x2_ASAP7_75t_L g1132 ( 
.A1(n_1032),
.A2(n_1046),
.B(n_1028),
.Y(n_1132)
);

NAND2xp5_ASAP7_75t_L g1133 ( 
.A(n_967),
.B(n_1056),
.Y(n_1133)
);

O2A1O1Ixp33_ASAP7_75t_L g1134 ( 
.A1(n_1055),
.A2(n_1084),
.B(n_998),
.C(n_1009),
.Y(n_1134)
);

INVx1_ASAP7_75t_L g1135 ( 
.A(n_989),
.Y(n_1135)
);

AOI21xp5_ASAP7_75t_L g1136 ( 
.A1(n_1036),
.A2(n_979),
.B(n_965),
.Y(n_1136)
);

NAND2xp5_ASAP7_75t_L g1137 ( 
.A(n_1056),
.B(n_981),
.Y(n_1137)
);

OR2x6_ASAP7_75t_L g1138 ( 
.A(n_1053),
.B(n_948),
.Y(n_1138)
);

AND2x2_ASAP7_75t_L g1139 ( 
.A(n_1070),
.B(n_1087),
.Y(n_1139)
);

NAND2xp5_ASAP7_75t_L g1140 ( 
.A(n_974),
.B(n_980),
.Y(n_1140)
);

AOI221xp5_ASAP7_75t_L g1141 ( 
.A1(n_993),
.A2(n_1075),
.B1(n_957),
.B2(n_1002),
.C(n_977),
.Y(n_1141)
);

INVxp67_ASAP7_75t_SL g1142 ( 
.A(n_998),
.Y(n_1142)
);

BUFx12f_ASAP7_75t_L g1143 ( 
.A(n_1054),
.Y(n_1143)
);

AOI21xp5_ASAP7_75t_SL g1144 ( 
.A1(n_1007),
.A2(n_1005),
.B(n_1028),
.Y(n_1144)
);

BUFx2_ASAP7_75t_R g1145 ( 
.A(n_982),
.Y(n_1145)
);

BUFx3_ASAP7_75t_L g1146 ( 
.A(n_1082),
.Y(n_1146)
);

A2O1A1Ixp33_ASAP7_75t_L g1147 ( 
.A1(n_1022),
.A2(n_1039),
.B(n_1033),
.C(n_1029),
.Y(n_1147)
);

BUFx10_ASAP7_75t_L g1148 ( 
.A(n_1014),
.Y(n_1148)
);

AOI21xp5_ASAP7_75t_L g1149 ( 
.A1(n_1042),
.A2(n_1030),
.B(n_1039),
.Y(n_1149)
);

AND2x2_ASAP7_75t_L g1150 ( 
.A(n_1021),
.B(n_948),
.Y(n_1150)
);

NAND2xp5_ASAP7_75t_L g1151 ( 
.A(n_1065),
.B(n_1086),
.Y(n_1151)
);

NAND2xp5_ASAP7_75t_SL g1152 ( 
.A(n_953),
.B(n_983),
.Y(n_1152)
);

OAI21xp5_ASAP7_75t_L g1153 ( 
.A1(n_964),
.A2(n_1030),
.B(n_1001),
.Y(n_1153)
);

OAI21xp5_ASAP7_75t_L g1154 ( 
.A1(n_964),
.A2(n_946),
.B(n_1076),
.Y(n_1154)
);

INVx3_ASAP7_75t_SL g1155 ( 
.A(n_948),
.Y(n_1155)
);

OAI21x1_ASAP7_75t_L g1156 ( 
.A1(n_1013),
.A2(n_1088),
.B(n_1006),
.Y(n_1156)
);

INVx1_ASAP7_75t_L g1157 ( 
.A(n_958),
.Y(n_1157)
);

INVx1_ASAP7_75t_L g1158 ( 
.A(n_969),
.Y(n_1158)
);

INVx1_ASAP7_75t_L g1159 ( 
.A(n_984),
.Y(n_1159)
);

OAI21x1_ASAP7_75t_L g1160 ( 
.A1(n_1013),
.A2(n_1088),
.B(n_1068),
.Y(n_1160)
);

O2A1O1Ixp5_ASAP7_75t_L g1161 ( 
.A1(n_956),
.A2(n_975),
.B(n_968),
.C(n_1086),
.Y(n_1161)
);

NAND2xp5_ASAP7_75t_L g1162 ( 
.A(n_968),
.B(n_1062),
.Y(n_1162)
);

OAI21x1_ASAP7_75t_L g1163 ( 
.A1(n_986),
.A2(n_1038),
.B(n_987),
.Y(n_1163)
);

NAND3xp33_ASAP7_75t_L g1164 ( 
.A(n_1038),
.B(n_987),
.C(n_995),
.Y(n_1164)
);

A2O1A1Ixp33_ASAP7_75t_L g1165 ( 
.A1(n_1018),
.A2(n_1062),
.B(n_1081),
.C(n_1071),
.Y(n_1165)
);

AOI221x1_ASAP7_75t_L g1166 ( 
.A1(n_987),
.A2(n_995),
.B1(n_975),
.B2(n_1071),
.C(n_1081),
.Y(n_1166)
);

AO31x2_ASAP7_75t_L g1167 ( 
.A1(n_995),
.A2(n_1053),
.A3(n_953),
.B(n_1071),
.Y(n_1167)
);

OAI21x1_ASAP7_75t_L g1168 ( 
.A1(n_953),
.A2(n_1053),
.B(n_1073),
.Y(n_1168)
);

INVx2_ASAP7_75t_L g1169 ( 
.A(n_1015),
.Y(n_1169)
);

BUFx8_ASAP7_75t_L g1170 ( 
.A(n_961),
.Y(n_1170)
);

OAI22xp5_ASAP7_75t_L g1171 ( 
.A1(n_1050),
.A2(n_940),
.B1(n_941),
.B2(n_1063),
.Y(n_1171)
);

NAND2xp5_ASAP7_75t_L g1172 ( 
.A(n_1067),
.B(n_940),
.Y(n_1172)
);

BUFx6f_ASAP7_75t_L g1173 ( 
.A(n_1023),
.Y(n_1173)
);

AO31x2_ASAP7_75t_L g1174 ( 
.A1(n_1000),
.A2(n_801),
.A3(n_805),
.B(n_990),
.Y(n_1174)
);

INVx2_ASAP7_75t_L g1175 ( 
.A(n_1015),
.Y(n_1175)
);

OAI22xp5_ASAP7_75t_L g1176 ( 
.A1(n_1050),
.A2(n_940),
.B1(n_941),
.B2(n_1063),
.Y(n_1176)
);

OAI21xp5_ASAP7_75t_L g1177 ( 
.A1(n_1050),
.A2(n_941),
.B(n_940),
.Y(n_1177)
);

AO21x2_ASAP7_75t_L g1178 ( 
.A1(n_990),
.A2(n_801),
.B(n_1000),
.Y(n_1178)
);

AOI21xp5_ASAP7_75t_L g1179 ( 
.A1(n_1049),
.A2(n_941),
.B(n_940),
.Y(n_1179)
);

O2A1O1Ixp33_ASAP7_75t_L g1180 ( 
.A1(n_960),
.A2(n_689),
.B(n_683),
.C(n_940),
.Y(n_1180)
);

AOI21xp5_ASAP7_75t_L g1181 ( 
.A1(n_1049),
.A2(n_941),
.B(n_940),
.Y(n_1181)
);

NOR2xp33_ASAP7_75t_L g1182 ( 
.A(n_1052),
.B(n_693),
.Y(n_1182)
);

INVx4_ASAP7_75t_L g1183 ( 
.A(n_1023),
.Y(n_1183)
);

AO31x2_ASAP7_75t_L g1184 ( 
.A1(n_1000),
.A2(n_801),
.A3(n_805),
.B(n_990),
.Y(n_1184)
);

OAI21x1_ASAP7_75t_L g1185 ( 
.A1(n_1012),
.A2(n_1059),
.B(n_1058),
.Y(n_1185)
);

A2O1A1Ixp33_ASAP7_75t_L g1186 ( 
.A1(n_1050),
.A2(n_940),
.B(n_941),
.C(n_910),
.Y(n_1186)
);

INVx1_ASAP7_75t_L g1187 ( 
.A(n_962),
.Y(n_1187)
);

AO32x2_ASAP7_75t_L g1188 ( 
.A1(n_950),
.A2(n_976),
.A3(n_1011),
.B1(n_1063),
.B2(n_1050),
.Y(n_1188)
);

INVxp67_ASAP7_75t_SL g1189 ( 
.A(n_973),
.Y(n_1189)
);

OAI21x1_ASAP7_75t_L g1190 ( 
.A1(n_1012),
.A2(n_1059),
.B(n_1058),
.Y(n_1190)
);

AND2x2_ASAP7_75t_L g1191 ( 
.A(n_1057),
.B(n_1085),
.Y(n_1191)
);

INVx2_ASAP7_75t_L g1192 ( 
.A(n_1015),
.Y(n_1192)
);

AOI21xp5_ASAP7_75t_L g1193 ( 
.A1(n_1049),
.A2(n_941),
.B(n_940),
.Y(n_1193)
);

OAI22xp5_ASAP7_75t_L g1194 ( 
.A1(n_1050),
.A2(n_940),
.B1(n_941),
.B2(n_1063),
.Y(n_1194)
);

CKINVDCx11_ASAP7_75t_R g1195 ( 
.A(n_947),
.Y(n_1195)
);

AOI21xp5_ASAP7_75t_L g1196 ( 
.A1(n_1049),
.A2(n_941),
.B(n_940),
.Y(n_1196)
);

O2A1O1Ixp5_ASAP7_75t_SL g1197 ( 
.A1(n_1041),
.A2(n_444),
.B(n_939),
.C(n_357),
.Y(n_1197)
);

CKINVDCx5p33_ASAP7_75t_R g1198 ( 
.A(n_947),
.Y(n_1198)
);

AOI21xp5_ASAP7_75t_L g1199 ( 
.A1(n_1049),
.A2(n_941),
.B(n_940),
.Y(n_1199)
);

INVx1_ASAP7_75t_L g1200 ( 
.A(n_962),
.Y(n_1200)
);

O2A1O1Ixp33_ASAP7_75t_L g1201 ( 
.A1(n_960),
.A2(n_689),
.B(n_683),
.C(n_940),
.Y(n_1201)
);

AOI21xp5_ASAP7_75t_L g1202 ( 
.A1(n_1049),
.A2(n_941),
.B(n_940),
.Y(n_1202)
);

NOR2xp33_ASAP7_75t_SL g1203 ( 
.A(n_994),
.B(n_918),
.Y(n_1203)
);

AOI21xp5_ASAP7_75t_L g1204 ( 
.A1(n_1049),
.A2(n_941),
.B(n_940),
.Y(n_1204)
);

INVx1_ASAP7_75t_L g1205 ( 
.A(n_962),
.Y(n_1205)
);

NAND2xp5_ASAP7_75t_L g1206 ( 
.A(n_1067),
.B(n_940),
.Y(n_1206)
);

AOI21xp5_ASAP7_75t_L g1207 ( 
.A1(n_1049),
.A2(n_941),
.B(n_940),
.Y(n_1207)
);

NAND2x1_ASAP7_75t_L g1208 ( 
.A(n_1013),
.B(n_1030),
.Y(n_1208)
);

INVx1_ASAP7_75t_L g1209 ( 
.A(n_962),
.Y(n_1209)
);

OAI22xp5_ASAP7_75t_L g1210 ( 
.A1(n_1050),
.A2(n_940),
.B1(n_941),
.B2(n_1063),
.Y(n_1210)
);

AOI221xp5_ASAP7_75t_SL g1211 ( 
.A1(n_960),
.A2(n_910),
.B1(n_950),
.B2(n_940),
.C(n_941),
.Y(n_1211)
);

OAI21x1_ASAP7_75t_L g1212 ( 
.A1(n_1012),
.A2(n_1059),
.B(n_1058),
.Y(n_1212)
);

BUFx6f_ASAP7_75t_L g1213 ( 
.A(n_1023),
.Y(n_1213)
);

AOI221xp5_ASAP7_75t_SL g1214 ( 
.A1(n_960),
.A2(n_910),
.B1(n_950),
.B2(n_940),
.C(n_941),
.Y(n_1214)
);

A2O1A1Ixp33_ASAP7_75t_L g1215 ( 
.A1(n_1050),
.A2(n_940),
.B(n_941),
.C(n_910),
.Y(n_1215)
);

AOI221x1_ASAP7_75t_L g1216 ( 
.A1(n_952),
.A2(n_910),
.B1(n_960),
.B2(n_1000),
.C(n_1061),
.Y(n_1216)
);

INVx5_ASAP7_75t_L g1217 ( 
.A(n_1053),
.Y(n_1217)
);

OA21x2_ASAP7_75t_L g1218 ( 
.A1(n_992),
.A2(n_978),
.B(n_988),
.Y(n_1218)
);

AO31x2_ASAP7_75t_L g1219 ( 
.A1(n_1000),
.A2(n_801),
.A3(n_805),
.B(n_990),
.Y(n_1219)
);

INVx1_ASAP7_75t_L g1220 ( 
.A(n_962),
.Y(n_1220)
);

NAND3xp33_ASAP7_75t_L g1221 ( 
.A(n_960),
.B(n_941),
.C(n_940),
.Y(n_1221)
);

OAI21x1_ASAP7_75t_L g1222 ( 
.A1(n_1012),
.A2(n_1059),
.B(n_1058),
.Y(n_1222)
);

AO31x2_ASAP7_75t_L g1223 ( 
.A1(n_1000),
.A2(n_801),
.A3(n_805),
.B(n_990),
.Y(n_1223)
);

BUFx2_ASAP7_75t_L g1224 ( 
.A(n_1069),
.Y(n_1224)
);

BUFx12f_ASAP7_75t_L g1225 ( 
.A(n_961),
.Y(n_1225)
);

AOI22xp33_ASAP7_75t_L g1226 ( 
.A1(n_1107),
.A2(n_1113),
.B1(n_1111),
.B2(n_1182),
.Y(n_1226)
);

AOI22xp33_ASAP7_75t_L g1227 ( 
.A1(n_1107),
.A2(n_1113),
.B1(n_1111),
.B2(n_1118),
.Y(n_1227)
);

INVx2_ASAP7_75t_L g1228 ( 
.A(n_1132),
.Y(n_1228)
);

AOI22xp33_ASAP7_75t_L g1229 ( 
.A1(n_1118),
.A2(n_1221),
.B1(n_1176),
.B2(n_1210),
.Y(n_1229)
);

INVx1_ASAP7_75t_L g1230 ( 
.A(n_1117),
.Y(n_1230)
);

NAND2xp5_ASAP7_75t_L g1231 ( 
.A(n_1140),
.B(n_1172),
.Y(n_1231)
);

AOI22xp33_ASAP7_75t_L g1232 ( 
.A1(n_1221),
.A2(n_1176),
.B1(n_1194),
.B2(n_1210),
.Y(n_1232)
);

OAI221xp5_ASAP7_75t_L g1233 ( 
.A1(n_1177),
.A2(n_1215),
.B1(n_1186),
.B2(n_1094),
.C(n_1194),
.Y(n_1233)
);

OAI22xp5_ASAP7_75t_L g1234 ( 
.A1(n_1171),
.A2(n_1177),
.B1(n_1125),
.B2(n_1090),
.Y(n_1234)
);

AOI22xp5_ASAP7_75t_SL g1235 ( 
.A1(n_1098),
.A2(n_1127),
.B1(n_1126),
.B2(n_1191),
.Y(n_1235)
);

BUFx4f_ASAP7_75t_L g1236 ( 
.A(n_1091),
.Y(n_1236)
);

AOI22xp5_ASAP7_75t_L g1237 ( 
.A1(n_1097),
.A2(n_1141),
.B1(n_1171),
.B2(n_1189),
.Y(n_1237)
);

OAI22xp33_ASAP7_75t_L g1238 ( 
.A1(n_1097),
.A2(n_1203),
.B1(n_1206),
.B2(n_1216),
.Y(n_1238)
);

INVx1_ASAP7_75t_SL g1239 ( 
.A(n_1110),
.Y(n_1239)
);

BUFx4f_ASAP7_75t_L g1240 ( 
.A(n_1091),
.Y(n_1240)
);

INVx1_ASAP7_75t_L g1241 ( 
.A(n_1121),
.Y(n_1241)
);

INVx1_ASAP7_75t_L g1242 ( 
.A(n_1135),
.Y(n_1242)
);

CKINVDCx20_ASAP7_75t_R g1243 ( 
.A(n_1122),
.Y(n_1243)
);

AOI22xp33_ASAP7_75t_L g1244 ( 
.A1(n_1114),
.A2(n_1175),
.B1(n_1169),
.B2(n_1192),
.Y(n_1244)
);

HB1xp67_ASAP7_75t_L g1245 ( 
.A(n_1133),
.Y(n_1245)
);

BUFx3_ASAP7_75t_L g1246 ( 
.A(n_1224),
.Y(n_1246)
);

INVx1_ASAP7_75t_L g1247 ( 
.A(n_1187),
.Y(n_1247)
);

CKINVDCx20_ASAP7_75t_R g1248 ( 
.A(n_1195),
.Y(n_1248)
);

AND2x2_ASAP7_75t_L g1249 ( 
.A(n_1106),
.B(n_1116),
.Y(n_1249)
);

INVx3_ASAP7_75t_L g1250 ( 
.A(n_1092),
.Y(n_1250)
);

NAND2xp5_ASAP7_75t_L g1251 ( 
.A(n_1124),
.B(n_1137),
.Y(n_1251)
);

AOI22xp33_ASAP7_75t_SL g1252 ( 
.A1(n_1203),
.A2(n_1125),
.B1(n_1123),
.B2(n_1153),
.Y(n_1252)
);

NAND2xp5_ASAP7_75t_L g1253 ( 
.A(n_1101),
.B(n_1180),
.Y(n_1253)
);

AOI22xp33_ASAP7_75t_L g1254 ( 
.A1(n_1154),
.A2(n_1102),
.B1(n_1153),
.B2(n_1159),
.Y(n_1254)
);

AOI22xp33_ASAP7_75t_L g1255 ( 
.A1(n_1154),
.A2(n_1158),
.B1(n_1157),
.B2(n_1130),
.Y(n_1255)
);

BUFx4_ASAP7_75t_R g1256 ( 
.A(n_1148),
.Y(n_1256)
);

BUFx4_ASAP7_75t_R g1257 ( 
.A(n_1146),
.Y(n_1257)
);

BUFx8_ASAP7_75t_L g1258 ( 
.A(n_1225),
.Y(n_1258)
);

INVx1_ASAP7_75t_L g1259 ( 
.A(n_1200),
.Y(n_1259)
);

INVx1_ASAP7_75t_L g1260 ( 
.A(n_1205),
.Y(n_1260)
);

INVx1_ASAP7_75t_L g1261 ( 
.A(n_1209),
.Y(n_1261)
);

INVx1_ASAP7_75t_L g1262 ( 
.A(n_1220),
.Y(n_1262)
);

CKINVDCx20_ASAP7_75t_R g1263 ( 
.A(n_1170),
.Y(n_1263)
);

AOI22xp33_ASAP7_75t_L g1264 ( 
.A1(n_1130),
.A2(n_1150),
.B1(n_1123),
.B2(n_1136),
.Y(n_1264)
);

AOI22xp33_ASAP7_75t_L g1265 ( 
.A1(n_1217),
.A2(n_1138),
.B1(n_1142),
.B2(n_1162),
.Y(n_1265)
);

INVx6_ASAP7_75t_L g1266 ( 
.A(n_1173),
.Y(n_1266)
);

INVx8_ASAP7_75t_L g1267 ( 
.A(n_1138),
.Y(n_1267)
);

OAI21xp5_ASAP7_75t_SL g1268 ( 
.A1(n_1201),
.A2(n_1105),
.B(n_1119),
.Y(n_1268)
);

AOI22xp33_ASAP7_75t_SL g1269 ( 
.A1(n_1119),
.A2(n_1168),
.B1(n_1164),
.B2(n_1188),
.Y(n_1269)
);

INVx1_ASAP7_75t_L g1270 ( 
.A(n_1134),
.Y(n_1270)
);

CKINVDCx11_ASAP7_75t_R g1271 ( 
.A(n_1143),
.Y(n_1271)
);

INVx1_ASAP7_75t_L g1272 ( 
.A(n_1188),
.Y(n_1272)
);

INVx1_ASAP7_75t_L g1273 ( 
.A(n_1188),
.Y(n_1273)
);

BUFx2_ASAP7_75t_L g1274 ( 
.A(n_1115),
.Y(n_1274)
);

AOI22xp33_ASAP7_75t_L g1275 ( 
.A1(n_1138),
.A2(n_1139),
.B1(n_1155),
.B2(n_1164),
.Y(n_1275)
);

NAND2xp5_ASAP7_75t_L g1276 ( 
.A(n_1211),
.B(n_1214),
.Y(n_1276)
);

INVx2_ASAP7_75t_L g1277 ( 
.A(n_1109),
.Y(n_1277)
);

INVx2_ASAP7_75t_L g1278 ( 
.A(n_1156),
.Y(n_1278)
);

BUFx2_ASAP7_75t_SL g1279 ( 
.A(n_1129),
.Y(n_1279)
);

OAI22xp5_ASAP7_75t_L g1280 ( 
.A1(n_1151),
.A2(n_1196),
.B1(n_1181),
.B2(n_1179),
.Y(n_1280)
);

CKINVDCx11_ASAP7_75t_R g1281 ( 
.A(n_1170),
.Y(n_1281)
);

INVx6_ASAP7_75t_L g1282 ( 
.A(n_1173),
.Y(n_1282)
);

BUFx3_ASAP7_75t_L g1283 ( 
.A(n_1173),
.Y(n_1283)
);

CKINVDCx11_ASAP7_75t_R g1284 ( 
.A(n_1198),
.Y(n_1284)
);

INVx1_ASAP7_75t_L g1285 ( 
.A(n_1160),
.Y(n_1285)
);

INVx1_ASAP7_75t_L g1286 ( 
.A(n_1167),
.Y(n_1286)
);

AND2x2_ASAP7_75t_L g1287 ( 
.A(n_1211),
.B(n_1214),
.Y(n_1287)
);

INVx1_ASAP7_75t_L g1288 ( 
.A(n_1167),
.Y(n_1288)
);

BUFx6f_ASAP7_75t_L g1289 ( 
.A(n_1213),
.Y(n_1289)
);

AND2x2_ASAP7_75t_L g1290 ( 
.A(n_1149),
.B(n_1223),
.Y(n_1290)
);

INVxp67_ASAP7_75t_L g1291 ( 
.A(n_1145),
.Y(n_1291)
);

INVx3_ASAP7_75t_L g1292 ( 
.A(n_1178),
.Y(n_1292)
);

AOI22xp33_ASAP7_75t_SL g1293 ( 
.A1(n_1178),
.A2(n_1163),
.B1(n_1193),
.B2(n_1204),
.Y(n_1293)
);

OAI22xp33_ASAP7_75t_L g1294 ( 
.A1(n_1183),
.A2(n_1129),
.B1(n_1213),
.B2(n_1199),
.Y(n_1294)
);

BUFx2_ASAP7_75t_L g1295 ( 
.A(n_1213),
.Y(n_1295)
);

CKINVDCx11_ASAP7_75t_R g1296 ( 
.A(n_1183),
.Y(n_1296)
);

CKINVDCx10_ASAP7_75t_R g1297 ( 
.A(n_1161),
.Y(n_1297)
);

AOI21xp5_ASAP7_75t_SL g1298 ( 
.A1(n_1147),
.A2(n_1152),
.B(n_1165),
.Y(n_1298)
);

BUFx8_ASAP7_75t_SL g1299 ( 
.A(n_1128),
.Y(n_1299)
);

INVx1_ASAP7_75t_SL g1300 ( 
.A(n_1128),
.Y(n_1300)
);

INVx6_ASAP7_75t_L g1301 ( 
.A(n_1166),
.Y(n_1301)
);

CKINVDCx11_ASAP7_75t_R g1302 ( 
.A(n_1208),
.Y(n_1302)
);

AOI22xp33_ASAP7_75t_L g1303 ( 
.A1(n_1202),
.A2(n_1207),
.B1(n_1144),
.B2(n_1112),
.Y(n_1303)
);

INVx1_ASAP7_75t_L g1304 ( 
.A(n_1096),
.Y(n_1304)
);

OAI22xp33_ASAP7_75t_L g1305 ( 
.A1(n_1100),
.A2(n_1104),
.B1(n_1108),
.B2(n_1218),
.Y(n_1305)
);

CKINVDCx6p67_ASAP7_75t_R g1306 ( 
.A(n_1197),
.Y(n_1306)
);

AOI22xp33_ASAP7_75t_L g1307 ( 
.A1(n_1089),
.A2(n_1099),
.B1(n_1218),
.B2(n_1131),
.Y(n_1307)
);

AND2x2_ASAP7_75t_L g1308 ( 
.A(n_1174),
.B(n_1223),
.Y(n_1308)
);

OAI22xp33_ASAP7_75t_L g1309 ( 
.A1(n_1089),
.A2(n_1099),
.B1(n_1223),
.B2(n_1184),
.Y(n_1309)
);

AOI22xp33_ASAP7_75t_L g1310 ( 
.A1(n_1120),
.A2(n_1103),
.B1(n_1095),
.B2(n_1222),
.Y(n_1310)
);

BUFx6f_ASAP7_75t_L g1311 ( 
.A(n_1093),
.Y(n_1311)
);

AOI22xp33_ASAP7_75t_L g1312 ( 
.A1(n_1185),
.A2(n_1190),
.B1(n_1212),
.B2(n_1184),
.Y(n_1312)
);

AOI22xp33_ASAP7_75t_L g1313 ( 
.A1(n_1219),
.A2(n_1107),
.B1(n_564),
.B2(n_489),
.Y(n_1313)
);

INVx1_ASAP7_75t_L g1314 ( 
.A(n_1117),
.Y(n_1314)
);

INVx1_ASAP7_75t_L g1315 ( 
.A(n_1117),
.Y(n_1315)
);

INVx1_ASAP7_75t_L g1316 ( 
.A(n_1117),
.Y(n_1316)
);

BUFx3_ASAP7_75t_L g1317 ( 
.A(n_1110),
.Y(n_1317)
);

AOI22xp5_ASAP7_75t_L g1318 ( 
.A1(n_1182),
.A2(n_478),
.B1(n_553),
.B2(n_1052),
.Y(n_1318)
);

CKINVDCx11_ASAP7_75t_R g1319 ( 
.A(n_1122),
.Y(n_1319)
);

INVx2_ASAP7_75t_L g1320 ( 
.A(n_1132),
.Y(n_1320)
);

OAI22xp5_ASAP7_75t_L g1321 ( 
.A1(n_1171),
.A2(n_941),
.B1(n_940),
.B2(n_1052),
.Y(n_1321)
);

CKINVDCx5p33_ASAP7_75t_R g1322 ( 
.A(n_1122),
.Y(n_1322)
);

INVx6_ASAP7_75t_L g1323 ( 
.A(n_1217),
.Y(n_1323)
);

INVx1_ASAP7_75t_L g1324 ( 
.A(n_1117),
.Y(n_1324)
);

BUFx4f_ASAP7_75t_SL g1325 ( 
.A(n_1225),
.Y(n_1325)
);

HB1xp67_ASAP7_75t_L g1326 ( 
.A(n_1133),
.Y(n_1326)
);

INVxp67_ASAP7_75t_SL g1327 ( 
.A(n_1133),
.Y(n_1327)
);

OAI21xp5_ASAP7_75t_SL g1328 ( 
.A1(n_1090),
.A2(n_1094),
.B(n_1052),
.Y(n_1328)
);

BUFx8_ASAP7_75t_SL g1329 ( 
.A(n_1198),
.Y(n_1329)
);

HB1xp67_ASAP7_75t_L g1330 ( 
.A(n_1133),
.Y(n_1330)
);

OAI21xp5_ASAP7_75t_SL g1331 ( 
.A1(n_1090),
.A2(n_1094),
.B(n_1052),
.Y(n_1331)
);

BUFx3_ASAP7_75t_L g1332 ( 
.A(n_1110),
.Y(n_1332)
);

BUFx8_ASAP7_75t_L g1333 ( 
.A(n_1225),
.Y(n_1333)
);

OAI22xp33_ASAP7_75t_L g1334 ( 
.A1(n_1113),
.A2(n_553),
.B1(n_1052),
.B2(n_941),
.Y(n_1334)
);

OAI22xp33_ASAP7_75t_L g1335 ( 
.A1(n_1113),
.A2(n_553),
.B1(n_1052),
.B2(n_941),
.Y(n_1335)
);

INVx3_ASAP7_75t_SL g1336 ( 
.A(n_1198),
.Y(n_1336)
);

OAI21x1_ASAP7_75t_L g1337 ( 
.A1(n_1307),
.A2(n_1303),
.B(n_1310),
.Y(n_1337)
);

NAND2xp5_ASAP7_75t_L g1338 ( 
.A(n_1327),
.B(n_1251),
.Y(n_1338)
);

INVx1_ASAP7_75t_L g1339 ( 
.A(n_1308),
.Y(n_1339)
);

AND2x2_ASAP7_75t_L g1340 ( 
.A(n_1272),
.B(n_1273),
.Y(n_1340)
);

OAI21x1_ASAP7_75t_L g1341 ( 
.A1(n_1280),
.A2(n_1292),
.B(n_1312),
.Y(n_1341)
);

OAI21xp5_ASAP7_75t_L g1342 ( 
.A1(n_1328),
.A2(n_1331),
.B(n_1234),
.Y(n_1342)
);

OAI21x1_ASAP7_75t_L g1343 ( 
.A1(n_1292),
.A2(n_1304),
.B(n_1277),
.Y(n_1343)
);

INVx1_ASAP7_75t_L g1344 ( 
.A(n_1308),
.Y(n_1344)
);

INVx1_ASAP7_75t_L g1345 ( 
.A(n_1285),
.Y(n_1345)
);

OAI22xp33_ASAP7_75t_L g1346 ( 
.A1(n_1318),
.A2(n_1237),
.B1(n_1335),
.B2(n_1334),
.Y(n_1346)
);

NAND2xp5_ASAP7_75t_L g1347 ( 
.A(n_1245),
.B(n_1326),
.Y(n_1347)
);

NAND2xp5_ASAP7_75t_L g1348 ( 
.A(n_1330),
.B(n_1232),
.Y(n_1348)
);

AND2x2_ASAP7_75t_L g1349 ( 
.A(n_1230),
.B(n_1241),
.Y(n_1349)
);

BUFx2_ASAP7_75t_L g1350 ( 
.A(n_1250),
.Y(n_1350)
);

CKINVDCx20_ASAP7_75t_R g1351 ( 
.A(n_1243),
.Y(n_1351)
);

HB1xp67_ASAP7_75t_L g1352 ( 
.A(n_1274),
.Y(n_1352)
);

BUFx3_ASAP7_75t_L g1353 ( 
.A(n_1301),
.Y(n_1353)
);

HB1xp67_ASAP7_75t_L g1354 ( 
.A(n_1246),
.Y(n_1354)
);

INVx1_ASAP7_75t_L g1355 ( 
.A(n_1242),
.Y(n_1355)
);

INVx2_ASAP7_75t_SL g1356 ( 
.A(n_1301),
.Y(n_1356)
);

BUFx4f_ASAP7_75t_L g1357 ( 
.A(n_1267),
.Y(n_1357)
);

INVx2_ASAP7_75t_L g1358 ( 
.A(n_1278),
.Y(n_1358)
);

NAND2xp5_ASAP7_75t_L g1359 ( 
.A(n_1226),
.B(n_1287),
.Y(n_1359)
);

INVxp33_ASAP7_75t_L g1360 ( 
.A(n_1235),
.Y(n_1360)
);

INVx1_ASAP7_75t_SL g1361 ( 
.A(n_1301),
.Y(n_1361)
);

OAI21x1_ASAP7_75t_L g1362 ( 
.A1(n_1290),
.A2(n_1320),
.B(n_1228),
.Y(n_1362)
);

AOI22xp33_ASAP7_75t_L g1363 ( 
.A1(n_1313),
.A2(n_1227),
.B1(n_1238),
.B2(n_1252),
.Y(n_1363)
);

NAND2xp5_ASAP7_75t_L g1364 ( 
.A(n_1287),
.B(n_1229),
.Y(n_1364)
);

HB1xp67_ASAP7_75t_L g1365 ( 
.A(n_1246),
.Y(n_1365)
);

INVxp67_ASAP7_75t_L g1366 ( 
.A(n_1249),
.Y(n_1366)
);

INVx1_ASAP7_75t_L g1367 ( 
.A(n_1247),
.Y(n_1367)
);

INVx1_ASAP7_75t_L g1368 ( 
.A(n_1259),
.Y(n_1368)
);

AND2x2_ASAP7_75t_L g1369 ( 
.A(n_1260),
.B(n_1261),
.Y(n_1369)
);

INVx1_ASAP7_75t_L g1370 ( 
.A(n_1262),
.Y(n_1370)
);

INVx1_ASAP7_75t_L g1371 ( 
.A(n_1314),
.Y(n_1371)
);

AND2x2_ASAP7_75t_L g1372 ( 
.A(n_1315),
.B(n_1316),
.Y(n_1372)
);

INVx1_ASAP7_75t_L g1373 ( 
.A(n_1324),
.Y(n_1373)
);

BUFx2_ASAP7_75t_L g1374 ( 
.A(n_1311),
.Y(n_1374)
);

AOI21x1_ASAP7_75t_L g1375 ( 
.A1(n_1253),
.A2(n_1276),
.B(n_1270),
.Y(n_1375)
);

OR2x6_ASAP7_75t_L g1376 ( 
.A(n_1267),
.B(n_1298),
.Y(n_1376)
);

AOI22xp33_ASAP7_75t_L g1377 ( 
.A1(n_1321),
.A2(n_1254),
.B1(n_1233),
.B2(n_1255),
.Y(n_1377)
);

INVx2_ASAP7_75t_SL g1378 ( 
.A(n_1317),
.Y(n_1378)
);

AND2x2_ASAP7_75t_L g1379 ( 
.A(n_1269),
.B(n_1264),
.Y(n_1379)
);

HB1xp67_ASAP7_75t_L g1380 ( 
.A(n_1300),
.Y(n_1380)
);

NAND2xp5_ASAP7_75t_L g1381 ( 
.A(n_1268),
.B(n_1231),
.Y(n_1381)
);

BUFx2_ASAP7_75t_L g1382 ( 
.A(n_1286),
.Y(n_1382)
);

AND2x2_ASAP7_75t_L g1383 ( 
.A(n_1288),
.B(n_1293),
.Y(n_1383)
);

HB1xp67_ASAP7_75t_L g1384 ( 
.A(n_1332),
.Y(n_1384)
);

AOI21xp5_ASAP7_75t_L g1385 ( 
.A1(n_1305),
.A2(n_1309),
.B(n_1294),
.Y(n_1385)
);

CKINVDCx5p33_ASAP7_75t_R g1386 ( 
.A(n_1281),
.Y(n_1386)
);

INVx1_ASAP7_75t_L g1387 ( 
.A(n_1306),
.Y(n_1387)
);

INVx1_ASAP7_75t_L g1388 ( 
.A(n_1306),
.Y(n_1388)
);

OA21x2_ASAP7_75t_L g1389 ( 
.A1(n_1265),
.A2(n_1244),
.B(n_1275),
.Y(n_1389)
);

INVx1_ASAP7_75t_SL g1390 ( 
.A(n_1297),
.Y(n_1390)
);

NAND2xp5_ASAP7_75t_L g1391 ( 
.A(n_1279),
.B(n_1289),
.Y(n_1391)
);

OA21x2_ASAP7_75t_L g1392 ( 
.A1(n_1295),
.A2(n_1323),
.B(n_1291),
.Y(n_1392)
);

AND2x2_ASAP7_75t_L g1393 ( 
.A(n_1332),
.B(n_1239),
.Y(n_1393)
);

INVx4_ASAP7_75t_L g1394 ( 
.A(n_1257),
.Y(n_1394)
);

AND2x4_ASAP7_75t_L g1395 ( 
.A(n_1283),
.B(n_1257),
.Y(n_1395)
);

INVx2_ASAP7_75t_L g1396 ( 
.A(n_1302),
.Y(n_1396)
);

INVx2_ASAP7_75t_L g1397 ( 
.A(n_1302),
.Y(n_1397)
);

HB1xp67_ASAP7_75t_L g1398 ( 
.A(n_1256),
.Y(n_1398)
);

AOI211xp5_ASAP7_75t_L g1399 ( 
.A1(n_1342),
.A2(n_1336),
.B(n_1322),
.C(n_1256),
.Y(n_1399)
);

INVx1_ASAP7_75t_L g1400 ( 
.A(n_1355),
.Y(n_1400)
);

INVx1_ASAP7_75t_L g1401 ( 
.A(n_1355),
.Y(n_1401)
);

OAI21x1_ASAP7_75t_SL g1402 ( 
.A1(n_1342),
.A2(n_1281),
.B(n_1296),
.Y(n_1402)
);

OR2x2_ASAP7_75t_L g1403 ( 
.A(n_1347),
.B(n_1322),
.Y(n_1403)
);

NAND2xp5_ASAP7_75t_L g1404 ( 
.A(n_1381),
.B(n_1299),
.Y(n_1404)
);

HB1xp67_ASAP7_75t_L g1405 ( 
.A(n_1352),
.Y(n_1405)
);

OAI21xp5_ASAP7_75t_L g1406 ( 
.A1(n_1346),
.A2(n_1236),
.B(n_1240),
.Y(n_1406)
);

OR2x2_ASAP7_75t_L g1407 ( 
.A(n_1347),
.B(n_1299),
.Y(n_1407)
);

NAND2xp5_ASAP7_75t_L g1408 ( 
.A(n_1381),
.B(n_1338),
.Y(n_1408)
);

OAI21x1_ASAP7_75t_SL g1409 ( 
.A1(n_1394),
.A2(n_1296),
.B(n_1333),
.Y(n_1409)
);

AND2x4_ASAP7_75t_SL g1410 ( 
.A(n_1394),
.B(n_1263),
.Y(n_1410)
);

AND2x2_ASAP7_75t_L g1411 ( 
.A(n_1340),
.B(n_1349),
.Y(n_1411)
);

OAI21xp5_ASAP7_75t_L g1412 ( 
.A1(n_1375),
.A2(n_1263),
.B(n_1243),
.Y(n_1412)
);

NAND4xp25_ASAP7_75t_L g1413 ( 
.A(n_1364),
.B(n_1319),
.C(n_1284),
.D(n_1325),
.Y(n_1413)
);

AOI22xp33_ASAP7_75t_L g1414 ( 
.A1(n_1379),
.A2(n_1271),
.B1(n_1266),
.B2(n_1282),
.Y(n_1414)
);

NAND2xp5_ASAP7_75t_L g1415 ( 
.A(n_1380),
.B(n_1258),
.Y(n_1415)
);

OA21x2_ASAP7_75t_L g1416 ( 
.A1(n_1341),
.A2(n_1258),
.B(n_1333),
.Y(n_1416)
);

AND2x4_ASAP7_75t_L g1417 ( 
.A(n_1353),
.B(n_1248),
.Y(n_1417)
);

AOI211xp5_ASAP7_75t_L g1418 ( 
.A1(n_1359),
.A2(n_1271),
.B(n_1319),
.C(n_1258),
.Y(n_1418)
);

AND2x4_ASAP7_75t_L g1419 ( 
.A(n_1353),
.B(n_1248),
.Y(n_1419)
);

NOR2xp33_ASAP7_75t_L g1420 ( 
.A(n_1351),
.B(n_1284),
.Y(n_1420)
);

AND2x4_ASAP7_75t_L g1421 ( 
.A(n_1353),
.B(n_1329),
.Y(n_1421)
);

AND2x2_ASAP7_75t_L g1422 ( 
.A(n_1349),
.B(n_1329),
.Y(n_1422)
);

OAI21xp5_ASAP7_75t_L g1423 ( 
.A1(n_1375),
.A2(n_1377),
.B(n_1363),
.Y(n_1423)
);

INVx1_ASAP7_75t_L g1424 ( 
.A(n_1367),
.Y(n_1424)
);

AND2x2_ASAP7_75t_L g1425 ( 
.A(n_1369),
.B(n_1372),
.Y(n_1425)
);

OAI21xp5_ASAP7_75t_L g1426 ( 
.A1(n_1364),
.A2(n_1379),
.B(n_1359),
.Y(n_1426)
);

AO32x2_ASAP7_75t_L g1427 ( 
.A1(n_1356),
.A2(n_1378),
.A3(n_1394),
.B1(n_1344),
.B2(n_1339),
.Y(n_1427)
);

AOI21xp5_ASAP7_75t_L g1428 ( 
.A1(n_1385),
.A2(n_1348),
.B(n_1376),
.Y(n_1428)
);

O2A1O1Ixp33_ASAP7_75t_SL g1429 ( 
.A1(n_1398),
.A2(n_1348),
.B(n_1397),
.C(n_1396),
.Y(n_1429)
);

AND2x2_ASAP7_75t_L g1430 ( 
.A(n_1369),
.B(n_1372),
.Y(n_1430)
);

OAI21x1_ASAP7_75t_L g1431 ( 
.A1(n_1337),
.A2(n_1385),
.B(n_1343),
.Y(n_1431)
);

BUFx3_ASAP7_75t_L g1432 ( 
.A(n_1395),
.Y(n_1432)
);

AOI21xp5_ASAP7_75t_L g1433 ( 
.A1(n_1376),
.A2(n_1388),
.B(n_1387),
.Y(n_1433)
);

BUFx2_ASAP7_75t_L g1434 ( 
.A(n_1374),
.Y(n_1434)
);

HB1xp67_ASAP7_75t_L g1435 ( 
.A(n_1354),
.Y(n_1435)
);

AND2x2_ASAP7_75t_L g1436 ( 
.A(n_1368),
.B(n_1370),
.Y(n_1436)
);

O2A1O1Ixp33_ASAP7_75t_SL g1437 ( 
.A1(n_1396),
.A2(n_1397),
.B(n_1365),
.C(n_1384),
.Y(n_1437)
);

OR2x2_ASAP7_75t_L g1438 ( 
.A(n_1344),
.B(n_1370),
.Y(n_1438)
);

OR2x6_ASAP7_75t_L g1439 ( 
.A(n_1392),
.B(n_1383),
.Y(n_1439)
);

OAI21xp5_ASAP7_75t_L g1440 ( 
.A1(n_1387),
.A2(n_1388),
.B(n_1337),
.Y(n_1440)
);

AND2x2_ASAP7_75t_L g1441 ( 
.A(n_1371),
.B(n_1373),
.Y(n_1441)
);

AO32x2_ASAP7_75t_L g1442 ( 
.A1(n_1382),
.A2(n_1361),
.A3(n_1392),
.B1(n_1366),
.B2(n_1362),
.Y(n_1442)
);

NAND2xp5_ASAP7_75t_L g1443 ( 
.A(n_1408),
.B(n_1345),
.Y(n_1443)
);

BUFx2_ASAP7_75t_L g1444 ( 
.A(n_1427),
.Y(n_1444)
);

NOR2xp33_ASAP7_75t_L g1445 ( 
.A(n_1413),
.B(n_1386),
.Y(n_1445)
);

AND2x2_ASAP7_75t_L g1446 ( 
.A(n_1411),
.B(n_1425),
.Y(n_1446)
);

AND2x2_ASAP7_75t_L g1447 ( 
.A(n_1425),
.B(n_1350),
.Y(n_1447)
);

BUFx2_ASAP7_75t_L g1448 ( 
.A(n_1427),
.Y(n_1448)
);

AOI22xp33_ASAP7_75t_SL g1449 ( 
.A1(n_1423),
.A2(n_1390),
.B1(n_1389),
.B2(n_1395),
.Y(n_1449)
);

INVx1_ASAP7_75t_L g1450 ( 
.A(n_1438),
.Y(n_1450)
);

INVx1_ASAP7_75t_L g1451 ( 
.A(n_1438),
.Y(n_1451)
);

NOR2x1p5_ASAP7_75t_L g1452 ( 
.A(n_1432),
.B(n_1395),
.Y(n_1452)
);

INVx1_ASAP7_75t_L g1453 ( 
.A(n_1400),
.Y(n_1453)
);

HB1xp67_ASAP7_75t_L g1454 ( 
.A(n_1405),
.Y(n_1454)
);

AOI22xp33_ASAP7_75t_L g1455 ( 
.A1(n_1426),
.A2(n_1389),
.B1(n_1360),
.B2(n_1390),
.Y(n_1455)
);

HB1xp67_ASAP7_75t_L g1456 ( 
.A(n_1435),
.Y(n_1456)
);

OR2x2_ASAP7_75t_L g1457 ( 
.A(n_1430),
.B(n_1382),
.Y(n_1457)
);

INVx4_ASAP7_75t_L g1458 ( 
.A(n_1421),
.Y(n_1458)
);

INVx1_ASAP7_75t_L g1459 ( 
.A(n_1401),
.Y(n_1459)
);

BUFx2_ASAP7_75t_L g1460 ( 
.A(n_1427),
.Y(n_1460)
);

AND2x2_ASAP7_75t_L g1461 ( 
.A(n_1427),
.B(n_1436),
.Y(n_1461)
);

BUFx2_ASAP7_75t_L g1462 ( 
.A(n_1427),
.Y(n_1462)
);

HB1xp67_ASAP7_75t_L g1463 ( 
.A(n_1434),
.Y(n_1463)
);

BUFx6f_ASAP7_75t_L g1464 ( 
.A(n_1431),
.Y(n_1464)
);

OAI22xp5_ASAP7_75t_L g1465 ( 
.A1(n_1399),
.A2(n_1357),
.B1(n_1391),
.B2(n_1393),
.Y(n_1465)
);

INVx1_ASAP7_75t_SL g1466 ( 
.A(n_1407),
.Y(n_1466)
);

NAND2xp5_ASAP7_75t_L g1467 ( 
.A(n_1441),
.B(n_1343),
.Y(n_1467)
);

INVx1_ASAP7_75t_L g1468 ( 
.A(n_1453),
.Y(n_1468)
);

BUFx2_ASAP7_75t_L g1469 ( 
.A(n_1444),
.Y(n_1469)
);

INVx1_ASAP7_75t_L g1470 ( 
.A(n_1453),
.Y(n_1470)
);

INVx1_ASAP7_75t_L g1471 ( 
.A(n_1459),
.Y(n_1471)
);

INVxp67_ASAP7_75t_SL g1472 ( 
.A(n_1463),
.Y(n_1472)
);

AND2x2_ASAP7_75t_L g1473 ( 
.A(n_1461),
.B(n_1440),
.Y(n_1473)
);

OAI31xp33_ASAP7_75t_L g1474 ( 
.A1(n_1455),
.A2(n_1428),
.A3(n_1429),
.B(n_1410),
.Y(n_1474)
);

NAND2xp5_ASAP7_75t_L g1475 ( 
.A(n_1443),
.B(n_1424),
.Y(n_1475)
);

AND2x2_ASAP7_75t_L g1476 ( 
.A(n_1461),
.B(n_1416),
.Y(n_1476)
);

BUFx6f_ASAP7_75t_L g1477 ( 
.A(n_1464),
.Y(n_1477)
);

INVx4_ASAP7_75t_L g1478 ( 
.A(n_1458),
.Y(n_1478)
);

OAI221xp5_ASAP7_75t_L g1479 ( 
.A1(n_1449),
.A2(n_1412),
.B1(n_1414),
.B2(n_1418),
.C(n_1429),
.Y(n_1479)
);

AO21x2_ASAP7_75t_L g1480 ( 
.A1(n_1467),
.A2(n_1431),
.B(n_1358),
.Y(n_1480)
);

AND2x2_ASAP7_75t_L g1481 ( 
.A(n_1461),
.B(n_1444),
.Y(n_1481)
);

INVxp67_ASAP7_75t_SL g1482 ( 
.A(n_1463),
.Y(n_1482)
);

AOI22xp33_ASAP7_75t_L g1483 ( 
.A1(n_1449),
.A2(n_1389),
.B1(n_1406),
.B2(n_1439),
.Y(n_1483)
);

INVx1_ASAP7_75t_L g1484 ( 
.A(n_1467),
.Y(n_1484)
);

INVx1_ASAP7_75t_L g1485 ( 
.A(n_1450),
.Y(n_1485)
);

AND2x2_ASAP7_75t_L g1486 ( 
.A(n_1448),
.B(n_1416),
.Y(n_1486)
);

AND2x2_ASAP7_75t_L g1487 ( 
.A(n_1448),
.B(n_1416),
.Y(n_1487)
);

AND2x2_ASAP7_75t_L g1488 ( 
.A(n_1460),
.B(n_1442),
.Y(n_1488)
);

NOR3xp33_ASAP7_75t_SL g1489 ( 
.A(n_1445),
.B(n_1420),
.C(n_1404),
.Y(n_1489)
);

AND2x2_ASAP7_75t_L g1490 ( 
.A(n_1460),
.B(n_1442),
.Y(n_1490)
);

AND2x2_ASAP7_75t_L g1491 ( 
.A(n_1462),
.B(n_1442),
.Y(n_1491)
);

AOI21x1_ASAP7_75t_L g1492 ( 
.A1(n_1462),
.A2(n_1433),
.B(n_1402),
.Y(n_1492)
);

OR2x6_ASAP7_75t_L g1493 ( 
.A(n_1452),
.B(n_1439),
.Y(n_1493)
);

AND2x2_ASAP7_75t_L g1494 ( 
.A(n_1446),
.B(n_1442),
.Y(n_1494)
);

AND2x2_ASAP7_75t_L g1495 ( 
.A(n_1446),
.B(n_1442),
.Y(n_1495)
);

INVx2_ASAP7_75t_L g1496 ( 
.A(n_1480),
.Y(n_1496)
);

INVx1_ASAP7_75t_L g1497 ( 
.A(n_1468),
.Y(n_1497)
);

AND2x2_ASAP7_75t_L g1498 ( 
.A(n_1494),
.B(n_1446),
.Y(n_1498)
);

OR2x2_ASAP7_75t_L g1499 ( 
.A(n_1484),
.B(n_1457),
.Y(n_1499)
);

NAND2xp5_ASAP7_75t_L g1500 ( 
.A(n_1484),
.B(n_1451),
.Y(n_1500)
);

INVx2_ASAP7_75t_L g1501 ( 
.A(n_1480),
.Y(n_1501)
);

BUFx2_ASAP7_75t_L g1502 ( 
.A(n_1469),
.Y(n_1502)
);

OR2x2_ASAP7_75t_L g1503 ( 
.A(n_1484),
.B(n_1457),
.Y(n_1503)
);

INVx2_ASAP7_75t_L g1504 ( 
.A(n_1480),
.Y(n_1504)
);

OR2x2_ASAP7_75t_L g1505 ( 
.A(n_1469),
.B(n_1451),
.Y(n_1505)
);

BUFx3_ASAP7_75t_L g1506 ( 
.A(n_1477),
.Y(n_1506)
);

AND2x2_ASAP7_75t_L g1507 ( 
.A(n_1494),
.B(n_1447),
.Y(n_1507)
);

AND2x4_ASAP7_75t_L g1508 ( 
.A(n_1493),
.B(n_1458),
.Y(n_1508)
);

AND2x2_ASAP7_75t_L g1509 ( 
.A(n_1495),
.B(n_1466),
.Y(n_1509)
);

INVx1_ASAP7_75t_L g1510 ( 
.A(n_1468),
.Y(n_1510)
);

INVx2_ASAP7_75t_L g1511 ( 
.A(n_1480),
.Y(n_1511)
);

OR2x2_ASAP7_75t_L g1512 ( 
.A(n_1469),
.B(n_1456),
.Y(n_1512)
);

INVx1_ASAP7_75t_L g1513 ( 
.A(n_1468),
.Y(n_1513)
);

AND2x2_ASAP7_75t_L g1514 ( 
.A(n_1495),
.B(n_1466),
.Y(n_1514)
);

INVx1_ASAP7_75t_L g1515 ( 
.A(n_1470),
.Y(n_1515)
);

OR2x2_ASAP7_75t_L g1516 ( 
.A(n_1495),
.B(n_1456),
.Y(n_1516)
);

NAND2xp5_ASAP7_75t_L g1517 ( 
.A(n_1470),
.B(n_1471),
.Y(n_1517)
);

INVx2_ASAP7_75t_L g1518 ( 
.A(n_1480),
.Y(n_1518)
);

INVx1_ASAP7_75t_SL g1519 ( 
.A(n_1475),
.Y(n_1519)
);

NAND2xp5_ASAP7_75t_L g1520 ( 
.A(n_1470),
.B(n_1454),
.Y(n_1520)
);

INVx1_ASAP7_75t_L g1521 ( 
.A(n_1471),
.Y(n_1521)
);

AND2x2_ASAP7_75t_L g1522 ( 
.A(n_1476),
.B(n_1481),
.Y(n_1522)
);

OR2x2_ASAP7_75t_L g1523 ( 
.A(n_1481),
.B(n_1454),
.Y(n_1523)
);

INVxp33_ASAP7_75t_L g1524 ( 
.A(n_1474),
.Y(n_1524)
);

HB1xp67_ASAP7_75t_L g1525 ( 
.A(n_1471),
.Y(n_1525)
);

AND2x2_ASAP7_75t_L g1526 ( 
.A(n_1476),
.B(n_1481),
.Y(n_1526)
);

NOR4xp25_ASAP7_75t_SL g1527 ( 
.A(n_1479),
.B(n_1437),
.C(n_1409),
.D(n_1402),
.Y(n_1527)
);

INVx1_ASAP7_75t_SL g1528 ( 
.A(n_1475),
.Y(n_1528)
);

INVx1_ASAP7_75t_L g1529 ( 
.A(n_1525),
.Y(n_1529)
);

OR2x2_ASAP7_75t_L g1530 ( 
.A(n_1523),
.B(n_1481),
.Y(n_1530)
);

INVx1_ASAP7_75t_L g1531 ( 
.A(n_1525),
.Y(n_1531)
);

INVx1_ASAP7_75t_L g1532 ( 
.A(n_1497),
.Y(n_1532)
);

OR2x2_ASAP7_75t_L g1533 ( 
.A(n_1523),
.B(n_1485),
.Y(n_1533)
);

NAND2xp5_ASAP7_75t_L g1534 ( 
.A(n_1519),
.B(n_1473),
.Y(n_1534)
);

INVx1_ASAP7_75t_L g1535 ( 
.A(n_1497),
.Y(n_1535)
);

INVx1_ASAP7_75t_L g1536 ( 
.A(n_1513),
.Y(n_1536)
);

INVxp67_ASAP7_75t_L g1537 ( 
.A(n_1512),
.Y(n_1537)
);

INVx2_ASAP7_75t_L g1538 ( 
.A(n_1502),
.Y(n_1538)
);

HB1xp67_ASAP7_75t_L g1539 ( 
.A(n_1502),
.Y(n_1539)
);

INVx3_ASAP7_75t_R g1540 ( 
.A(n_1502),
.Y(n_1540)
);

INVx1_ASAP7_75t_L g1541 ( 
.A(n_1513),
.Y(n_1541)
);

INVx1_ASAP7_75t_L g1542 ( 
.A(n_1510),
.Y(n_1542)
);

INVx3_ASAP7_75t_L g1543 ( 
.A(n_1508),
.Y(n_1543)
);

INVx3_ASAP7_75t_L g1544 ( 
.A(n_1508),
.Y(n_1544)
);

NAND2xp5_ASAP7_75t_L g1545 ( 
.A(n_1528),
.B(n_1473),
.Y(n_1545)
);

INVx1_ASAP7_75t_L g1546 ( 
.A(n_1510),
.Y(n_1546)
);

INVx1_ASAP7_75t_L g1547 ( 
.A(n_1510),
.Y(n_1547)
);

AOI211xp5_ASAP7_75t_SL g1548 ( 
.A1(n_1524),
.A2(n_1479),
.B(n_1465),
.C(n_1437),
.Y(n_1548)
);

NAND2x1_ASAP7_75t_L g1549 ( 
.A(n_1508),
.B(n_1478),
.Y(n_1549)
);

INVx1_ASAP7_75t_SL g1550 ( 
.A(n_1512),
.Y(n_1550)
);

NOR2xp33_ASAP7_75t_L g1551 ( 
.A(n_1524),
.B(n_1407),
.Y(n_1551)
);

INVx1_ASAP7_75t_L g1552 ( 
.A(n_1515),
.Y(n_1552)
);

AND2x2_ASAP7_75t_L g1553 ( 
.A(n_1498),
.B(n_1473),
.Y(n_1553)
);

INVx1_ASAP7_75t_L g1554 ( 
.A(n_1515),
.Y(n_1554)
);

INVx1_ASAP7_75t_L g1555 ( 
.A(n_1515),
.Y(n_1555)
);

INVx2_ASAP7_75t_L g1556 ( 
.A(n_1505),
.Y(n_1556)
);

NOR2xp33_ASAP7_75t_L g1557 ( 
.A(n_1519),
.B(n_1458),
.Y(n_1557)
);

BUFx2_ASAP7_75t_SL g1558 ( 
.A(n_1509),
.Y(n_1558)
);

NAND2xp5_ASAP7_75t_L g1559 ( 
.A(n_1528),
.B(n_1473),
.Y(n_1559)
);

INVx1_ASAP7_75t_L g1560 ( 
.A(n_1521),
.Y(n_1560)
);

AND2x4_ASAP7_75t_L g1561 ( 
.A(n_1508),
.B(n_1493),
.Y(n_1561)
);

INVx1_ASAP7_75t_L g1562 ( 
.A(n_1521),
.Y(n_1562)
);

AND2x2_ASAP7_75t_L g1563 ( 
.A(n_1498),
.B(n_1476),
.Y(n_1563)
);

INVx1_ASAP7_75t_L g1564 ( 
.A(n_1521),
.Y(n_1564)
);

INVx3_ASAP7_75t_L g1565 ( 
.A(n_1508),
.Y(n_1565)
);

INVx2_ASAP7_75t_SL g1566 ( 
.A(n_1523),
.Y(n_1566)
);

INVx1_ASAP7_75t_L g1567 ( 
.A(n_1517),
.Y(n_1567)
);

NAND3xp33_ASAP7_75t_L g1568 ( 
.A(n_1527),
.B(n_1474),
.C(n_1488),
.Y(n_1568)
);

NOR2xp33_ASAP7_75t_L g1569 ( 
.A(n_1512),
.B(n_1422),
.Y(n_1569)
);

INVx1_ASAP7_75t_L g1570 ( 
.A(n_1517),
.Y(n_1570)
);

INVx1_ASAP7_75t_L g1571 ( 
.A(n_1532),
.Y(n_1571)
);

OR2x2_ASAP7_75t_L g1572 ( 
.A(n_1550),
.B(n_1516),
.Y(n_1572)
);

AND2x2_ASAP7_75t_L g1573 ( 
.A(n_1553),
.B(n_1498),
.Y(n_1573)
);

NAND2xp5_ASAP7_75t_L g1574 ( 
.A(n_1551),
.B(n_1509),
.Y(n_1574)
);

AND2x2_ASAP7_75t_L g1575 ( 
.A(n_1553),
.B(n_1558),
.Y(n_1575)
);

INVx2_ASAP7_75t_SL g1576 ( 
.A(n_1538),
.Y(n_1576)
);

AND2x2_ASAP7_75t_L g1577 ( 
.A(n_1566),
.B(n_1522),
.Y(n_1577)
);

NAND2xp5_ASAP7_75t_L g1578 ( 
.A(n_1551),
.B(n_1509),
.Y(n_1578)
);

OR2x2_ASAP7_75t_L g1579 ( 
.A(n_1530),
.B(n_1516),
.Y(n_1579)
);

NAND2xp5_ASAP7_75t_L g1580 ( 
.A(n_1569),
.B(n_1514),
.Y(n_1580)
);

INVx1_ASAP7_75t_L g1581 ( 
.A(n_1535),
.Y(n_1581)
);

AND2x2_ASAP7_75t_L g1582 ( 
.A(n_1566),
.B(n_1522),
.Y(n_1582)
);

AND2x4_ASAP7_75t_L g1583 ( 
.A(n_1538),
.B(n_1508),
.Y(n_1583)
);

NOR2xp33_ASAP7_75t_L g1584 ( 
.A(n_1569),
.B(n_1422),
.Y(n_1584)
);

OR2x2_ASAP7_75t_L g1585 ( 
.A(n_1530),
.B(n_1516),
.Y(n_1585)
);

AND2x2_ASAP7_75t_L g1586 ( 
.A(n_1563),
.B(n_1522),
.Y(n_1586)
);

OR2x2_ASAP7_75t_L g1587 ( 
.A(n_1534),
.B(n_1499),
.Y(n_1587)
);

INVx1_ASAP7_75t_L g1588 ( 
.A(n_1536),
.Y(n_1588)
);

NAND2xp5_ASAP7_75t_L g1589 ( 
.A(n_1548),
.B(n_1514),
.Y(n_1589)
);

INVx1_ASAP7_75t_L g1590 ( 
.A(n_1541),
.Y(n_1590)
);

OR2x2_ASAP7_75t_L g1591 ( 
.A(n_1545),
.B(n_1559),
.Y(n_1591)
);

AND2x2_ASAP7_75t_L g1592 ( 
.A(n_1563),
.B(n_1526),
.Y(n_1592)
);

OR2x6_ASAP7_75t_L g1593 ( 
.A(n_1568),
.B(n_1409),
.Y(n_1593)
);

NAND2xp5_ASAP7_75t_L g1594 ( 
.A(n_1537),
.B(n_1514),
.Y(n_1594)
);

NAND2xp5_ASAP7_75t_L g1595 ( 
.A(n_1539),
.B(n_1488),
.Y(n_1595)
);

INVx1_ASAP7_75t_L g1596 ( 
.A(n_1529),
.Y(n_1596)
);

INVx1_ASAP7_75t_L g1597 ( 
.A(n_1531),
.Y(n_1597)
);

OAI22xp5_ASAP7_75t_L g1598 ( 
.A1(n_1543),
.A2(n_1527),
.B1(n_1483),
.B2(n_1526),
.Y(n_1598)
);

AND2x4_ASAP7_75t_L g1599 ( 
.A(n_1561),
.B(n_1526),
.Y(n_1599)
);

OR2x2_ASAP7_75t_L g1600 ( 
.A(n_1556),
.B(n_1499),
.Y(n_1600)
);

INVx1_ASAP7_75t_L g1601 ( 
.A(n_1542),
.Y(n_1601)
);

AND2x2_ASAP7_75t_L g1602 ( 
.A(n_1543),
.B(n_1507),
.Y(n_1602)
);

NAND2xp5_ASAP7_75t_L g1603 ( 
.A(n_1556),
.B(n_1488),
.Y(n_1603)
);

INVx1_ASAP7_75t_SL g1604 ( 
.A(n_1549),
.Y(n_1604)
);

AND2x2_ASAP7_75t_L g1605 ( 
.A(n_1543),
.B(n_1544),
.Y(n_1605)
);

NAND2xp5_ASAP7_75t_L g1606 ( 
.A(n_1584),
.B(n_1567),
.Y(n_1606)
);

INVx1_ASAP7_75t_L g1607 ( 
.A(n_1601),
.Y(n_1607)
);

NOR3xp33_ASAP7_75t_L g1608 ( 
.A(n_1589),
.B(n_1565),
.C(n_1544),
.Y(n_1608)
);

AND2x2_ASAP7_75t_L g1609 ( 
.A(n_1575),
.B(n_1557),
.Y(n_1609)
);

OAI21xp33_ASAP7_75t_L g1610 ( 
.A1(n_1574),
.A2(n_1557),
.B(n_1570),
.Y(n_1610)
);

OAI31xp33_ASAP7_75t_L g1611 ( 
.A1(n_1598),
.A2(n_1491),
.A3(n_1490),
.B(n_1488),
.Y(n_1611)
);

INVx1_ASAP7_75t_L g1612 ( 
.A(n_1571),
.Y(n_1612)
);

INVx1_ASAP7_75t_L g1613 ( 
.A(n_1581),
.Y(n_1613)
);

NAND2xp5_ASAP7_75t_L g1614 ( 
.A(n_1584),
.B(n_1507),
.Y(n_1614)
);

INVx1_ASAP7_75t_L g1615 ( 
.A(n_1588),
.Y(n_1615)
);

INVx1_ASAP7_75t_SL g1616 ( 
.A(n_1593),
.Y(n_1616)
);

NAND2x1_ASAP7_75t_SL g1617 ( 
.A(n_1575),
.B(n_1544),
.Y(n_1617)
);

AND2x2_ASAP7_75t_L g1618 ( 
.A(n_1599),
.B(n_1565),
.Y(n_1618)
);

INVx1_ASAP7_75t_L g1619 ( 
.A(n_1590),
.Y(n_1619)
);

NAND2xp5_ASAP7_75t_L g1620 ( 
.A(n_1576),
.B(n_1507),
.Y(n_1620)
);

AOI22xp5_ASAP7_75t_L g1621 ( 
.A1(n_1578),
.A2(n_1491),
.B1(n_1490),
.B2(n_1483),
.Y(n_1621)
);

NAND2xp33_ASAP7_75t_L g1622 ( 
.A(n_1576),
.B(n_1489),
.Y(n_1622)
);

INVx1_ASAP7_75t_L g1623 ( 
.A(n_1596),
.Y(n_1623)
);

OAI321xp33_ASAP7_75t_L g1624 ( 
.A1(n_1593),
.A2(n_1492),
.A3(n_1491),
.B1(n_1490),
.B2(n_1501),
.C(n_1496),
.Y(n_1624)
);

AND2x2_ASAP7_75t_L g1625 ( 
.A(n_1599),
.B(n_1565),
.Y(n_1625)
);

OR2x2_ASAP7_75t_L g1626 ( 
.A(n_1572),
.B(n_1533),
.Y(n_1626)
);

AND2x2_ASAP7_75t_L g1627 ( 
.A(n_1599),
.B(n_1549),
.Y(n_1627)
);

INVx1_ASAP7_75t_L g1628 ( 
.A(n_1597),
.Y(n_1628)
);

INVx1_ASAP7_75t_SL g1629 ( 
.A(n_1593),
.Y(n_1629)
);

INVx1_ASAP7_75t_L g1630 ( 
.A(n_1600),
.Y(n_1630)
);

AOI322xp5_ASAP7_75t_L g1631 ( 
.A1(n_1621),
.A2(n_1490),
.A3(n_1491),
.B1(n_1603),
.B2(n_1580),
.C1(n_1595),
.C2(n_1594),
.Y(n_1631)
);

AOI21xp5_ASAP7_75t_L g1632 ( 
.A1(n_1622),
.A2(n_1593),
.B(n_1604),
.Y(n_1632)
);

AND2x2_ASAP7_75t_L g1633 ( 
.A(n_1609),
.B(n_1573),
.Y(n_1633)
);

OAI222xp33_ASAP7_75t_L g1634 ( 
.A1(n_1616),
.A2(n_1572),
.B1(n_1591),
.B2(n_1579),
.C1(n_1585),
.C2(n_1587),
.Y(n_1634)
);

AOI22xp5_ASAP7_75t_L g1635 ( 
.A1(n_1622),
.A2(n_1487),
.B1(n_1486),
.B2(n_1583),
.Y(n_1635)
);

OAI22xp33_ASAP7_75t_L g1636 ( 
.A1(n_1624),
.A2(n_1585),
.B1(n_1579),
.B2(n_1493),
.Y(n_1636)
);

INVx1_ASAP7_75t_L g1637 ( 
.A(n_1626),
.Y(n_1637)
);

INVxp67_ASAP7_75t_L g1638 ( 
.A(n_1629),
.Y(n_1638)
);

AOI221x1_ASAP7_75t_L g1639 ( 
.A1(n_1608),
.A2(n_1583),
.B1(n_1605),
.B2(n_1555),
.C(n_1552),
.Y(n_1639)
);

NOR2xp33_ASAP7_75t_L g1640 ( 
.A(n_1606),
.B(n_1540),
.Y(n_1640)
);

AND2x2_ASAP7_75t_L g1641 ( 
.A(n_1609),
.B(n_1573),
.Y(n_1641)
);

INVx1_ASAP7_75t_SL g1642 ( 
.A(n_1617),
.Y(n_1642)
);

AOI22xp5_ASAP7_75t_L g1643 ( 
.A1(n_1630),
.A2(n_1620),
.B1(n_1610),
.B2(n_1618),
.Y(n_1643)
);

AOI22xp5_ASAP7_75t_L g1644 ( 
.A1(n_1618),
.A2(n_1486),
.B1(n_1487),
.B2(n_1583),
.Y(n_1644)
);

INVx1_ASAP7_75t_L g1645 ( 
.A(n_1626),
.Y(n_1645)
);

AND2x2_ASAP7_75t_L g1646 ( 
.A(n_1625),
.B(n_1577),
.Y(n_1646)
);

NAND2xp5_ASAP7_75t_L g1647 ( 
.A(n_1613),
.B(n_1577),
.Y(n_1647)
);

AOI21xp33_ASAP7_75t_SL g1648 ( 
.A1(n_1611),
.A2(n_1582),
.B(n_1605),
.Y(n_1648)
);

NAND2xp5_ASAP7_75t_L g1649 ( 
.A(n_1613),
.B(n_1582),
.Y(n_1649)
);

AOI22xp33_ASAP7_75t_L g1650 ( 
.A1(n_1636),
.A2(n_1474),
.B1(n_1496),
.B2(n_1518),
.Y(n_1650)
);

OR2x2_ASAP7_75t_L g1651 ( 
.A(n_1637),
.B(n_1614),
.Y(n_1651)
);

OAI21xp5_ASAP7_75t_L g1652 ( 
.A1(n_1639),
.A2(n_1617),
.B(n_1625),
.Y(n_1652)
);

AOI22xp5_ASAP7_75t_L g1653 ( 
.A1(n_1640),
.A2(n_1628),
.B1(n_1623),
.B2(n_1615),
.Y(n_1653)
);

AOI22xp5_ASAP7_75t_L g1654 ( 
.A1(n_1635),
.A2(n_1487),
.B1(n_1486),
.B2(n_1612),
.Y(n_1654)
);

INVxp67_ASAP7_75t_L g1655 ( 
.A(n_1645),
.Y(n_1655)
);

OR2x2_ASAP7_75t_L g1656 ( 
.A(n_1647),
.B(n_1619),
.Y(n_1656)
);

AND2x2_ASAP7_75t_L g1657 ( 
.A(n_1633),
.B(n_1627),
.Y(n_1657)
);

AOI322xp5_ASAP7_75t_L g1658 ( 
.A1(n_1638),
.A2(n_1607),
.A3(n_1486),
.B1(n_1487),
.B2(n_1518),
.C1(n_1501),
.C2(n_1511),
.Y(n_1658)
);

OAI21xp33_ASAP7_75t_L g1659 ( 
.A1(n_1641),
.A2(n_1627),
.B(n_1602),
.Y(n_1659)
);

INVx1_ASAP7_75t_L g1660 ( 
.A(n_1647),
.Y(n_1660)
);

AND2x2_ASAP7_75t_L g1661 ( 
.A(n_1646),
.B(n_1586),
.Y(n_1661)
);

NOR2xp33_ASAP7_75t_SL g1662 ( 
.A(n_1657),
.B(n_1634),
.Y(n_1662)
);

INVxp33_ASAP7_75t_L g1663 ( 
.A(n_1652),
.Y(n_1663)
);

NOR2x1_ASAP7_75t_L g1664 ( 
.A(n_1660),
.B(n_1642),
.Y(n_1664)
);

NOR4xp25_ASAP7_75t_L g1665 ( 
.A(n_1655),
.B(n_1649),
.C(n_1540),
.D(n_1602),
.Y(n_1665)
);

INVx1_ASAP7_75t_L g1666 ( 
.A(n_1661),
.Y(n_1666)
);

NAND4xp25_ASAP7_75t_L g1667 ( 
.A(n_1653),
.B(n_1632),
.C(n_1643),
.D(n_1649),
.Y(n_1667)
);

NOR2x1_ASAP7_75t_L g1668 ( 
.A(n_1656),
.B(n_1415),
.Y(n_1668)
);

OAI21xp33_ASAP7_75t_L g1669 ( 
.A1(n_1659),
.A2(n_1631),
.B(n_1648),
.Y(n_1669)
);

NOR2xp33_ASAP7_75t_L g1670 ( 
.A(n_1651),
.B(n_1653),
.Y(n_1670)
);

NAND2xp5_ASAP7_75t_SL g1671 ( 
.A(n_1662),
.B(n_1665),
.Y(n_1671)
);

AOI211xp5_ASAP7_75t_L g1672 ( 
.A1(n_1663),
.A2(n_1654),
.B(n_1644),
.C(n_1592),
.Y(n_1672)
);

AOI22xp5_ASAP7_75t_L g1673 ( 
.A1(n_1670),
.A2(n_1650),
.B1(n_1561),
.B2(n_1592),
.Y(n_1673)
);

OAI221xp5_ASAP7_75t_L g1674 ( 
.A1(n_1664),
.A2(n_1658),
.B1(n_1511),
.B2(n_1518),
.C(n_1501),
.Y(n_1674)
);

NOR3xp33_ASAP7_75t_L g1675 ( 
.A(n_1667),
.B(n_1501),
.C(n_1496),
.Y(n_1675)
);

CKINVDCx20_ASAP7_75t_R g1676 ( 
.A(n_1671),
.Y(n_1676)
);

NAND4xp75_ASAP7_75t_L g1677 ( 
.A(n_1673),
.B(n_1666),
.C(n_1668),
.D(n_1669),
.Y(n_1677)
);

NOR3xp33_ASAP7_75t_L g1678 ( 
.A(n_1674),
.B(n_1504),
.C(n_1496),
.Y(n_1678)
);

NAND2xp33_ASAP7_75t_L g1679 ( 
.A(n_1675),
.B(n_1489),
.Y(n_1679)
);

NOR4xp75_ASAP7_75t_SL g1680 ( 
.A(n_1672),
.B(n_1520),
.C(n_1465),
.D(n_1500),
.Y(n_1680)
);

NAND2xp33_ASAP7_75t_L g1681 ( 
.A(n_1671),
.B(n_1586),
.Y(n_1681)
);

AND2x4_ASAP7_75t_L g1682 ( 
.A(n_1676),
.B(n_1403),
.Y(n_1682)
);

NOR2x1_ASAP7_75t_L g1683 ( 
.A(n_1677),
.B(n_1546),
.Y(n_1683)
);

INVxp67_ASAP7_75t_L g1684 ( 
.A(n_1681),
.Y(n_1684)
);

NAND4xp75_ASAP7_75t_L g1685 ( 
.A(n_1680),
.B(n_1679),
.C(n_1678),
.D(n_1393),
.Y(n_1685)
);

INVxp67_ASAP7_75t_L g1686 ( 
.A(n_1681),
.Y(n_1686)
);

OAI211xp5_ASAP7_75t_L g1687 ( 
.A1(n_1684),
.A2(n_1506),
.B(n_1562),
.C(n_1564),
.Y(n_1687)
);

AOI22xp5_ASAP7_75t_L g1688 ( 
.A1(n_1686),
.A2(n_1561),
.B1(n_1419),
.B2(n_1417),
.Y(n_1688)
);

NAND3x1_ASAP7_75t_L g1689 ( 
.A(n_1683),
.B(n_1554),
.C(n_1547),
.Y(n_1689)
);

NAND2xp5_ASAP7_75t_L g1690 ( 
.A(n_1688),
.B(n_1682),
.Y(n_1690)
);

AOI22xp5_ASAP7_75t_L g1691 ( 
.A1(n_1690),
.A2(n_1685),
.B1(n_1689),
.B2(n_1687),
.Y(n_1691)
);

OAI22xp5_ASAP7_75t_L g1692 ( 
.A1(n_1691),
.A2(n_1533),
.B1(n_1560),
.B2(n_1505),
.Y(n_1692)
);

AND2x4_ASAP7_75t_L g1693 ( 
.A(n_1692),
.B(n_1403),
.Y(n_1693)
);

AOI21xp5_ASAP7_75t_L g1694 ( 
.A1(n_1693),
.A2(n_1511),
.B(n_1504),
.Y(n_1694)
);

AO21x2_ASAP7_75t_L g1695 ( 
.A1(n_1694),
.A2(n_1511),
.B(n_1504),
.Y(n_1695)
);

INVx1_ASAP7_75t_L g1696 ( 
.A(n_1694),
.Y(n_1696)
);

OAI321xp33_ASAP7_75t_L g1697 ( 
.A1(n_1696),
.A2(n_1518),
.A3(n_1504),
.B1(n_1520),
.B2(n_1492),
.C(n_1505),
.Y(n_1697)
);

OAI21xp5_ASAP7_75t_L g1698 ( 
.A1(n_1695),
.A2(n_1419),
.B(n_1417),
.Y(n_1698)
);

OAI22xp5_ASAP7_75t_L g1699 ( 
.A1(n_1698),
.A2(n_1695),
.B1(n_1506),
.B2(n_1503),
.Y(n_1699)
);

INVx1_ASAP7_75t_L g1700 ( 
.A(n_1697),
.Y(n_1700)
);

OAI221xp5_ASAP7_75t_R g1701 ( 
.A1(n_1700),
.A2(n_1506),
.B1(n_1482),
.B2(n_1472),
.C(n_1503),
.Y(n_1701)
);

AOI211xp5_ASAP7_75t_L g1702 ( 
.A1(n_1701),
.A2(n_1699),
.B(n_1419),
.C(n_1417),
.Y(n_1702)
);


endmodule