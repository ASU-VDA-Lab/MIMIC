module fake_aes_7609_n_676 (n_117, n_44, n_133, n_149, n_81, n_69, n_22, n_57, n_88, n_52, n_26, n_50, n_33, n_102, n_73, n_49, n_119, n_141, n_115, n_97, n_80, n_167, n_107, n_158, n_60, n_114, n_121, n_41, n_35, n_94, n_65, n_171, n_125, n_9, n_161, n_10, n_177, n_130, n_103, n_19, n_87, n_137, n_180, n_104, n_160, n_98, n_74, n_154, n_7, n_29, n_165, n_146, n_45, n_85, n_181, n_101, n_62, n_36, n_47, n_37, n_34, n_5, n_23, n_8, n_91, n_108, n_116, n_155, n_139, n_16, n_13, n_169, n_152, n_113, n_95, n_124, n_156, n_128, n_120, n_129, n_70, n_17, n_63, n_14, n_71, n_90, n_56, n_135, n_42, n_24, n_78, n_6, n_4, n_127, n_170, n_40, n_111, n_157, n_79, n_38, n_64, n_142, n_184, n_46, n_31, n_58, n_122, n_138, n_126, n_178, n_118, n_32, n_0, n_179, n_84, n_131, n_112, n_55, n_12, n_86, n_143, n_182, n_166, n_162, n_75, n_163, n_105, n_159, n_174, n_72, n_136, n_43, n_76, n_89, n_176, n_68, n_144, n_27, n_53, n_183, n_67, n_77, n_20, n_2, n_147, n_54, n_148, n_123, n_83, n_172, n_28, n_48, n_100, n_92, n_11, n_25, n_30, n_59, n_150, n_168, n_3, n_18, n_110, n_66, n_134, n_1, n_164, n_82, n_106, n_175, n_15, n_173, n_145, n_153, n_61, n_21, n_99, n_109, n_93, n_132, n_151, n_51, n_140, n_96, n_39, n_676);
input n_117;
input n_44;
input n_133;
input n_149;
input n_81;
input n_69;
input n_22;
input n_57;
input n_88;
input n_52;
input n_26;
input n_50;
input n_33;
input n_102;
input n_73;
input n_49;
input n_119;
input n_141;
input n_115;
input n_97;
input n_80;
input n_167;
input n_107;
input n_158;
input n_60;
input n_114;
input n_121;
input n_41;
input n_35;
input n_94;
input n_65;
input n_171;
input n_125;
input n_9;
input n_161;
input n_10;
input n_177;
input n_130;
input n_103;
input n_19;
input n_87;
input n_137;
input n_180;
input n_104;
input n_160;
input n_98;
input n_74;
input n_154;
input n_7;
input n_29;
input n_165;
input n_146;
input n_45;
input n_85;
input n_181;
input n_101;
input n_62;
input n_36;
input n_47;
input n_37;
input n_34;
input n_5;
input n_23;
input n_8;
input n_91;
input n_108;
input n_116;
input n_155;
input n_139;
input n_16;
input n_13;
input n_169;
input n_152;
input n_113;
input n_95;
input n_124;
input n_156;
input n_128;
input n_120;
input n_129;
input n_70;
input n_17;
input n_63;
input n_14;
input n_71;
input n_90;
input n_56;
input n_135;
input n_42;
input n_24;
input n_78;
input n_6;
input n_4;
input n_127;
input n_170;
input n_40;
input n_111;
input n_157;
input n_79;
input n_38;
input n_64;
input n_142;
input n_184;
input n_46;
input n_31;
input n_58;
input n_122;
input n_138;
input n_126;
input n_178;
input n_118;
input n_32;
input n_0;
input n_179;
input n_84;
input n_131;
input n_112;
input n_55;
input n_12;
input n_86;
input n_143;
input n_182;
input n_166;
input n_162;
input n_75;
input n_163;
input n_105;
input n_159;
input n_174;
input n_72;
input n_136;
input n_43;
input n_76;
input n_89;
input n_176;
input n_68;
input n_144;
input n_27;
input n_53;
input n_183;
input n_67;
input n_77;
input n_20;
input n_2;
input n_147;
input n_54;
input n_148;
input n_123;
input n_83;
input n_172;
input n_28;
input n_48;
input n_100;
input n_92;
input n_11;
input n_25;
input n_30;
input n_59;
input n_150;
input n_168;
input n_3;
input n_18;
input n_110;
input n_66;
input n_134;
input n_1;
input n_164;
input n_82;
input n_106;
input n_175;
input n_15;
input n_173;
input n_145;
input n_153;
input n_61;
input n_21;
input n_99;
input n_109;
input n_93;
input n_132;
input n_151;
input n_51;
input n_140;
input n_96;
input n_39;
output n_676;
wire n_663;
wire n_361;
wire n_513;
wire n_185;
wire n_603;
wire n_604;
wire n_590;
wire n_407;
wire n_646;
wire n_284;
wire n_278;
wire n_500;
wire n_607;
wire n_431;
wire n_484;
wire n_496;
wire n_667;
wire n_189;
wire n_311;
wire n_292;
wire n_309;
wire n_612;
wire n_328;
wire n_655;
wire n_468;
wire n_523;
wire n_229;
wire n_336;
wire n_464;
wire n_448;
wire n_645;
wire n_348;
wire n_252;
wire n_637;
wire n_353;
wire n_564;
wire n_528;
wire n_206;
wire n_288;
wire n_383;
wire n_661;
wire n_672;
wire n_532;
wire n_627;
wire n_544;
wire n_400;
wire n_296;
wire n_202;
wire n_386;
wire n_432;
wire n_659;
wire n_232;
wire n_462;
wire n_316;
wire n_545;
wire n_211;
wire n_334;
wire n_389;
wire n_548;
wire n_436;
wire n_588;
wire n_275;
wire n_463;
wire n_205;
wire n_330;
wire n_587;
wire n_662;
wire n_387;
wire n_434;
wire n_384;
wire n_227;
wire n_476;
wire n_617;
wire n_231;
wire n_452;
wire n_518;
wire n_547;
wire n_298;
wire n_628;
wire n_411;
wire n_598;
wire n_489;
wire n_199;
wire n_351;
wire n_401;
wire n_305;
wire n_461;
wire n_599;
wire n_228;
wire n_345;
wire n_360;
wire n_236;
wire n_340;
wire n_481;
wire n_443;
wire n_373;
wire n_576;
wire n_301;
wire n_222;
wire n_234;
wire n_465;
wire n_609;
wire n_636;
wire n_366;
wire n_596;
wire n_286;
wire n_190;
wire n_246;
wire n_321;
wire n_572;
wire n_324;
wire n_392;
wire n_668;
wire n_652;
wire n_279;
wire n_303;
wire n_437;
wire n_512;
wire n_326;
wire n_289;
wire n_333;
wire n_249;
wire n_642;
wire n_586;
wire n_671;
wire n_244;
wire n_563;
wire n_540;
wire n_638;
wire n_517;
wire n_560;
wire n_479;
wire n_623;
wire n_593;
wire n_554;
wire n_447;
wire n_608;
wire n_567;
wire n_196;
wire n_580;
wire n_192;
wire n_502;
wire n_543;
wire n_312;
wire n_455;
wire n_529;
wire n_630;
wire n_511;
wire n_277;
wire n_467;
wire n_647;
wire n_367;
wire n_644;
wire n_250;
wire n_314;
wire n_237;
wire n_255;
wire n_426;
wire n_624;
wire n_230;
wire n_209;
wire n_274;
wire n_282;
wire n_319;
wire n_499;
wire n_417;
wire n_241;
wire n_575;
wire n_238;
wire n_318;
wire n_471;
wire n_632;
wire n_293;
wire n_506;
wire n_533;
wire n_393;
wire n_247;
wire n_490;
wire n_648;
wire n_613;
wire n_381;
wire n_550;
wire n_304;
wire n_399;
wire n_665;
wire n_571;
wire n_294;
wire n_459;
wire n_313;
wire n_210;
wire n_322;
wire n_310;
wire n_191;
wire n_307;
wire n_634;
wire n_610;
wire n_474;
wire n_354;
wire n_402;
wire n_413;
wire n_391;
wire n_427;
wire n_460;
wire n_478;
wire n_243;
wire n_235;
wire n_415;
wire n_394;
wire n_482;
wire n_442;
wire n_331;
wire n_485;
wire n_352;
wire n_619;
wire n_268;
wire n_501;
wire n_248;
wire n_299;
wire n_338;
wire n_519;
wire n_256;
wire n_551;
wire n_404;
wire n_369;
wire n_509;
wire n_651;
wire n_674;
wire n_329;
wire n_251;
wire n_635;
wire n_525;
wire n_218;
wire n_507;
wire n_605;
wire n_611;
wire n_633;
wire n_271;
wire n_626;
wire n_302;
wire n_466;
wire n_270;
wire n_362;
wire n_259;
wire n_308;
wire n_546;
wire n_412;
wire n_664;
wire n_207;
wire n_565;
wire n_224;
wire n_219;
wire n_475;
wire n_578;
wire n_542;
wire n_537;
wire n_214;
wire n_204;
wire n_660;
wire n_430;
wire n_450;
wire n_579;
wire n_403;
wire n_557;
wire n_516;
wire n_254;
wire n_549;
wire n_622;
wire n_262;
wire n_556;
wire n_239;
wire n_439;
wire n_601;
wire n_379;
wire n_641;
wire n_614;
wire n_527;
wire n_526;
wire n_276;
wire n_649;
wire n_320;
wire n_285;
wire n_195;
wire n_446;
wire n_420;
wire n_423;
wire n_342;
wire n_621;
wire n_666;
wire n_370;
wire n_589;
wire n_643;
wire n_574;
wire n_217;
wire n_388;
wire n_454;
wire n_193;
wire n_273;
wire n_505;
wire n_390;
wire n_514;
wire n_486;
wire n_568;
wire n_357;
wire n_245;
wire n_653;
wire n_260;
wire n_539;
wire n_197;
wire n_201;
wire n_591;
wire n_317;
wire n_416;
wire n_374;
wire n_536;
wire n_265;
wire n_264;
wire n_522;
wire n_200;
wire n_208;
wire n_573;
wire n_673;
wire n_669;
wire n_616;
wire n_365;
wire n_541;
wire n_315;
wire n_363;
wire n_409;
wire n_295;
wire n_654;
wire n_263;
wire n_495;
wire n_186;
wire n_364;
wire n_428;
wire n_566;
wire n_376;
wire n_639;
wire n_552;
wire n_344;
wire n_503;
wire n_283;
wire n_520;
wire n_435;
wire n_216;
wire n_577;
wire n_615;
wire n_212;
wire n_472;
wire n_419;
wire n_396;
wire n_477;
wire n_508;
wire n_570;
wire n_398;
wire n_445;
wire n_656;
wire n_438;
wire n_640;
wire n_429;
wire n_488;
wire n_233;
wire n_440;
wire n_553;
wire n_422;
wire n_327;
wire n_325;
wire n_349;
wire n_498;
wire n_597;
wire n_225;
wire n_535;
wire n_530;
wire n_220;
wire n_358;
wire n_267;
wire n_221;
wire n_456;
wire n_203;
wire n_449;
wire n_300;
wire n_524;
wire n_584;
wire n_497;
wire n_339;
wire n_657;
wire n_583;
wire n_620;
wire n_240;
wire n_378;
wire n_582;
wire n_359;
wire n_346;
wire n_441;
wire n_561;
wire n_335;
wire n_272;
wire n_594;
wire n_534;
wire n_531;
wire n_397;
wire n_306;
wire n_215;
wire n_242;
wire n_602;
wire n_198;
wire n_424;
wire n_629;
wire n_569;
wire n_297;
wire n_410;
wire n_188;
wire n_377;
wire n_510;
wire n_343;
wire n_675;
wire n_291;
wire n_504;
wire n_458;
wire n_581;
wire n_418;
wire n_493;
wire n_555;
wire n_380;
wire n_618;
wire n_356;
wire n_281;
wire n_341;
wire n_470;
wire n_600;
wire n_187;
wire n_375;
wire n_451;
wire n_487;
wire n_371;
wire n_323;
wire n_473;
wire n_347;
wire n_558;
wire n_258;
wire n_253;
wire n_515;
wire n_670;
wire n_266;
wire n_213;
wire n_538;
wire n_492;
wire n_592;
wire n_368;
wire n_355;
wire n_226;
wire n_382;
wire n_337;
wire n_658;
wire n_444;
wire n_521;
wire n_625;
wire n_650;
wire n_469;
wire n_585;
wire n_457;
wire n_595;
wire n_223;
wire n_494;
wire n_559;
wire n_480;
wire n_372;
wire n_453;
wire n_631;
wire n_194;
wire n_287;
wire n_261;
wire n_606;
wire n_425;
wire n_332;
wire n_414;
wire n_562;
wire n_350;
wire n_433;
wire n_421;
wire n_483;
wire n_408;
wire n_290;
wire n_405;
wire n_280;
wire n_395;
wire n_406;
wire n_491;
wire n_385;
wire n_257;
wire n_269;
CKINVDCx16_ASAP7_75t_R g185 ( .A(n_67), .Y(n_185) );
CKINVDCx5p33_ASAP7_75t_R g186 ( .A(n_133), .Y(n_186) );
BUFx10_ASAP7_75t_L g187 ( .A(n_125), .Y(n_187) );
HB1xp67_ASAP7_75t_L g188 ( .A(n_101), .Y(n_188) );
CKINVDCx5p33_ASAP7_75t_R g189 ( .A(n_20), .Y(n_189) );
INVx1_ASAP7_75t_L g190 ( .A(n_160), .Y(n_190) );
INVx1_ASAP7_75t_L g191 ( .A(n_70), .Y(n_191) );
CKINVDCx20_ASAP7_75t_R g192 ( .A(n_162), .Y(n_192) );
BUFx3_ASAP7_75t_L g193 ( .A(n_74), .Y(n_193) );
CKINVDCx5p33_ASAP7_75t_R g194 ( .A(n_179), .Y(n_194) );
CKINVDCx5p33_ASAP7_75t_R g195 ( .A(n_137), .Y(n_195) );
BUFx3_ASAP7_75t_L g196 ( .A(n_151), .Y(n_196) );
INVx1_ASAP7_75t_SL g197 ( .A(n_128), .Y(n_197) );
INVx1_ASAP7_75t_L g198 ( .A(n_167), .Y(n_198) );
INVx1_ASAP7_75t_L g199 ( .A(n_127), .Y(n_199) );
BUFx3_ASAP7_75t_L g200 ( .A(n_184), .Y(n_200) );
NAND2xp5_ASAP7_75t_L g201 ( .A(n_178), .B(n_95), .Y(n_201) );
INVxp67_ASAP7_75t_SL g202 ( .A(n_148), .Y(n_202) );
INVx1_ASAP7_75t_L g203 ( .A(n_9), .Y(n_203) );
CKINVDCx20_ASAP7_75t_R g204 ( .A(n_5), .Y(n_204) );
INVx1_ASAP7_75t_L g205 ( .A(n_159), .Y(n_205) );
BUFx6f_ASAP7_75t_L g206 ( .A(n_103), .Y(n_206) );
INVx1_ASAP7_75t_SL g207 ( .A(n_113), .Y(n_207) );
INVx1_ASAP7_75t_L g208 ( .A(n_41), .Y(n_208) );
CKINVDCx5p33_ASAP7_75t_R g209 ( .A(n_12), .Y(n_209) );
INVx1_ASAP7_75t_L g210 ( .A(n_3), .Y(n_210) );
INVx1_ASAP7_75t_L g211 ( .A(n_172), .Y(n_211) );
INVx1_ASAP7_75t_L g212 ( .A(n_98), .Y(n_212) );
INVx1_ASAP7_75t_SL g213 ( .A(n_153), .Y(n_213) );
INVx1_ASAP7_75t_L g214 ( .A(n_163), .Y(n_214) );
INVx1_ASAP7_75t_L g215 ( .A(n_106), .Y(n_215) );
HB1xp67_ASAP7_75t_L g216 ( .A(n_72), .Y(n_216) );
INVx1_ASAP7_75t_L g217 ( .A(n_89), .Y(n_217) );
BUFx6f_ASAP7_75t_L g218 ( .A(n_29), .Y(n_218) );
INVx1_ASAP7_75t_L g219 ( .A(n_123), .Y(n_219) );
INVx1_ASAP7_75t_L g220 ( .A(n_3), .Y(n_220) );
CKINVDCx5p33_ASAP7_75t_R g221 ( .A(n_136), .Y(n_221) );
INVx1_ASAP7_75t_L g222 ( .A(n_154), .Y(n_222) );
INVx1_ASAP7_75t_L g223 ( .A(n_114), .Y(n_223) );
INVx1_ASAP7_75t_SL g224 ( .A(n_36), .Y(n_224) );
INVx2_ASAP7_75t_L g225 ( .A(n_177), .Y(n_225) );
BUFx10_ASAP7_75t_L g226 ( .A(n_42), .Y(n_226) );
INVx1_ASAP7_75t_L g227 ( .A(n_66), .Y(n_227) );
INVx1_ASAP7_75t_L g228 ( .A(n_9), .Y(n_228) );
INVx2_ASAP7_75t_L g229 ( .A(n_116), .Y(n_229) );
INVx1_ASAP7_75t_L g230 ( .A(n_149), .Y(n_230) );
INVx1_ASAP7_75t_L g231 ( .A(n_156), .Y(n_231) );
BUFx2_ASAP7_75t_SL g232 ( .A(n_171), .Y(n_232) );
INVx1_ASAP7_75t_L g233 ( .A(n_5), .Y(n_233) );
BUFx3_ASAP7_75t_L g234 ( .A(n_51), .Y(n_234) );
CKINVDCx5p33_ASAP7_75t_R g235 ( .A(n_34), .Y(n_235) );
BUFx3_ASAP7_75t_L g236 ( .A(n_173), .Y(n_236) );
INVx1_ASAP7_75t_L g237 ( .A(n_180), .Y(n_237) );
CKINVDCx5p33_ASAP7_75t_R g238 ( .A(n_24), .Y(n_238) );
CKINVDCx5p33_ASAP7_75t_R g239 ( .A(n_37), .Y(n_239) );
CKINVDCx5p33_ASAP7_75t_R g240 ( .A(n_13), .Y(n_240) );
INVxp67_ASAP7_75t_L g241 ( .A(n_166), .Y(n_241) );
INVx2_ASAP7_75t_L g242 ( .A(n_126), .Y(n_242) );
CKINVDCx5p33_ASAP7_75t_R g243 ( .A(n_97), .Y(n_243) );
INVxp33_ASAP7_75t_SL g244 ( .A(n_16), .Y(n_244) );
INVx1_ASAP7_75t_L g245 ( .A(n_19), .Y(n_245) );
INVx1_ASAP7_75t_L g246 ( .A(n_124), .Y(n_246) );
INVx1_ASAP7_75t_L g247 ( .A(n_119), .Y(n_247) );
INVx1_ASAP7_75t_L g248 ( .A(n_183), .Y(n_248) );
CKINVDCx14_ASAP7_75t_R g249 ( .A(n_31), .Y(n_249) );
INVx1_ASAP7_75t_L g250 ( .A(n_158), .Y(n_250) );
BUFx3_ASAP7_75t_L g251 ( .A(n_142), .Y(n_251) );
INVx1_ASAP7_75t_L g252 ( .A(n_155), .Y(n_252) );
INVx1_ASAP7_75t_L g253 ( .A(n_32), .Y(n_253) );
INVx1_ASAP7_75t_L g254 ( .A(n_147), .Y(n_254) );
CKINVDCx20_ASAP7_75t_R g255 ( .A(n_30), .Y(n_255) );
INVx1_ASAP7_75t_L g256 ( .A(n_26), .Y(n_256) );
CKINVDCx20_ASAP7_75t_R g257 ( .A(n_8), .Y(n_257) );
INVx2_ASAP7_75t_L g258 ( .A(n_129), .Y(n_258) );
HB1xp67_ASAP7_75t_L g259 ( .A(n_65), .Y(n_259) );
CKINVDCx16_ASAP7_75t_R g260 ( .A(n_115), .Y(n_260) );
INVx1_ASAP7_75t_L g261 ( .A(n_68), .Y(n_261) );
INVx1_ASAP7_75t_L g262 ( .A(n_39), .Y(n_262) );
INVx1_ASAP7_75t_L g263 ( .A(n_157), .Y(n_263) );
CKINVDCx20_ASAP7_75t_R g264 ( .A(n_170), .Y(n_264) );
INVx1_ASAP7_75t_L g265 ( .A(n_20), .Y(n_265) );
NOR2xp67_ASAP7_75t_L g266 ( .A(n_109), .B(n_87), .Y(n_266) );
CKINVDCx20_ASAP7_75t_R g267 ( .A(n_1), .Y(n_267) );
CKINVDCx20_ASAP7_75t_R g268 ( .A(n_46), .Y(n_268) );
INVx1_ASAP7_75t_L g269 ( .A(n_161), .Y(n_269) );
CKINVDCx20_ASAP7_75t_R g270 ( .A(n_182), .Y(n_270) );
INVx1_ASAP7_75t_L g271 ( .A(n_41), .Y(n_271) );
BUFx6f_ASAP7_75t_L g272 ( .A(n_84), .Y(n_272) );
CKINVDCx5p33_ASAP7_75t_R g273 ( .A(n_55), .Y(n_273) );
BUFx5_ASAP7_75t_L g274 ( .A(n_11), .Y(n_274) );
INVx1_ASAP7_75t_L g275 ( .A(n_34), .Y(n_275) );
CKINVDCx5p33_ASAP7_75t_R g276 ( .A(n_85), .Y(n_276) );
BUFx6f_ASAP7_75t_L g277 ( .A(n_92), .Y(n_277) );
INVxp67_ASAP7_75t_SL g278 ( .A(n_77), .Y(n_278) );
CKINVDCx14_ASAP7_75t_R g279 ( .A(n_168), .Y(n_279) );
INVx1_ASAP7_75t_L g280 ( .A(n_48), .Y(n_280) );
CKINVDCx5p33_ASAP7_75t_R g281 ( .A(n_169), .Y(n_281) );
CKINVDCx20_ASAP7_75t_R g282 ( .A(n_40), .Y(n_282) );
INVx2_ASAP7_75t_L g283 ( .A(n_25), .Y(n_283) );
BUFx3_ASAP7_75t_L g284 ( .A(n_120), .Y(n_284) );
INVx1_ASAP7_75t_L g285 ( .A(n_82), .Y(n_285) );
CKINVDCx5p33_ASAP7_75t_R g286 ( .A(n_181), .Y(n_286) );
BUFx2_ASAP7_75t_L g287 ( .A(n_146), .Y(n_287) );
INVxp67_ASAP7_75t_L g288 ( .A(n_150), .Y(n_288) );
INVx1_ASAP7_75t_L g289 ( .A(n_175), .Y(n_289) );
INVx2_ASAP7_75t_L g290 ( .A(n_206), .Y(n_290) );
BUFx6f_ASAP7_75t_L g291 ( .A(n_206), .Y(n_291) );
BUFx6f_ASAP7_75t_L g292 ( .A(n_206), .Y(n_292) );
AND2x6_ASAP7_75t_L g293 ( .A(n_193), .B(n_60), .Y(n_293) );
INVx2_ASAP7_75t_L g294 ( .A(n_206), .Y(n_294) );
CKINVDCx5p33_ASAP7_75t_R g295 ( .A(n_185), .Y(n_295) );
BUFx6f_ASAP7_75t_L g296 ( .A(n_272), .Y(n_296) );
AND2x4_ASAP7_75t_SL g297 ( .A(n_187), .B(n_61), .Y(n_297) );
AND2x6_ASAP7_75t_L g298 ( .A(n_193), .B(n_62), .Y(n_298) );
NOR2x1_ASAP7_75t_L g299 ( .A(n_234), .B(n_0), .Y(n_299) );
HB1xp67_ASAP7_75t_L g300 ( .A(n_249), .Y(n_300) );
INVx2_ASAP7_75t_L g301 ( .A(n_272), .Y(n_301) );
INVx1_ASAP7_75t_L g302 ( .A(n_274), .Y(n_302) );
BUFx6f_ASAP7_75t_L g303 ( .A(n_272), .Y(n_303) );
OAI21x1_ASAP7_75t_L g304 ( .A1(n_225), .A2(n_64), .B(n_63), .Y(n_304) );
INVx2_ASAP7_75t_L g305 ( .A(n_277), .Y(n_305) );
BUFx2_ASAP7_75t_L g306 ( .A(n_234), .Y(n_306) );
AOI22xp5_ASAP7_75t_L g307 ( .A1(n_244), .A2(n_1), .B1(n_2), .B2(n_4), .Y(n_307) );
AOI22xp5_ASAP7_75t_SL g308 ( .A1(n_204), .A2(n_2), .B1(n_4), .B2(n_6), .Y(n_308) );
NAND2xp5_ASAP7_75t_L g309 ( .A(n_287), .B(n_6), .Y(n_309) );
BUFx3_ASAP7_75t_L g310 ( .A(n_196), .Y(n_310) );
OA21x2_ASAP7_75t_L g311 ( .A1(n_225), .A2(n_71), .B(n_69), .Y(n_311) );
NOR2xp33_ASAP7_75t_L g312 ( .A(n_188), .B(n_216), .Y(n_312) );
INVx1_ASAP7_75t_L g313 ( .A(n_274), .Y(n_313) );
INVx1_ASAP7_75t_L g314 ( .A(n_274), .Y(n_314) );
INVx1_ASAP7_75t_L g315 ( .A(n_274), .Y(n_315) );
AND2x2_ASAP7_75t_L g316 ( .A(n_279), .B(n_7), .Y(n_316) );
BUFx6f_ASAP7_75t_L g317 ( .A(n_277), .Y(n_317) );
BUFx3_ASAP7_75t_L g318 ( .A(n_196), .Y(n_318) );
INVx1_ASAP7_75t_SL g319 ( .A(n_189), .Y(n_319) );
AND2x2_ASAP7_75t_R g320 ( .A(n_204), .B(n_7), .Y(n_320) );
XNOR2xp5_ASAP7_75t_L g321 ( .A(n_308), .B(n_255), .Y(n_321) );
BUFx3_ASAP7_75t_L g322 ( .A(n_310), .Y(n_322) );
INVx2_ASAP7_75t_SL g323 ( .A(n_310), .Y(n_323) );
BUFx3_ASAP7_75t_L g324 ( .A(n_310), .Y(n_324) );
BUFx3_ASAP7_75t_L g325 ( .A(n_318), .Y(n_325) );
INVx3_ASAP7_75t_L g326 ( .A(n_302), .Y(n_326) );
AND2x2_ASAP7_75t_L g327 ( .A(n_306), .B(n_279), .Y(n_327) );
NAND2xp5_ASAP7_75t_SL g328 ( .A(n_300), .B(n_260), .Y(n_328) );
INVx2_ASAP7_75t_L g329 ( .A(n_291), .Y(n_329) );
AND2x6_ASAP7_75t_L g330 ( .A(n_316), .B(n_200), .Y(n_330) );
BUFx2_ASAP7_75t_L g331 ( .A(n_316), .Y(n_331) );
AOI22xp33_ASAP7_75t_L g332 ( .A1(n_313), .A2(n_208), .B1(n_210), .B2(n_203), .Y(n_332) );
INVx2_ASAP7_75t_L g333 ( .A(n_291), .Y(n_333) );
HB1xp67_ASAP7_75t_L g334 ( .A(n_319), .Y(n_334) );
INVx1_ASAP7_75t_L g335 ( .A(n_313), .Y(n_335) );
INVx3_ASAP7_75t_L g336 ( .A(n_314), .Y(n_336) );
NAND2xp5_ASAP7_75t_L g337 ( .A(n_318), .B(n_259), .Y(n_337) );
NOR2xp33_ASAP7_75t_L g338 ( .A(n_312), .B(n_241), .Y(n_338) );
NAND2xp5_ASAP7_75t_L g339 ( .A(n_314), .B(n_229), .Y(n_339) );
BUFx10_ASAP7_75t_L g340 ( .A(n_297), .Y(n_340) );
BUFx6f_ASAP7_75t_L g341 ( .A(n_291), .Y(n_341) );
INVx4_ASAP7_75t_L g342 ( .A(n_293), .Y(n_342) );
NOR2xp33_ASAP7_75t_L g343 ( .A(n_309), .B(n_288), .Y(n_343) );
INVx3_ASAP7_75t_L g344 ( .A(n_315), .Y(n_344) );
OR2x2_ASAP7_75t_L g345 ( .A(n_295), .B(n_189), .Y(n_345) );
NAND3xp33_ASAP7_75t_L g346 ( .A(n_315), .B(n_289), .C(n_191), .Y(n_346) );
INVx4_ASAP7_75t_L g347 ( .A(n_293), .Y(n_347) );
NAND2xp5_ASAP7_75t_SL g348 ( .A(n_297), .B(n_187), .Y(n_348) );
BUFx6f_ASAP7_75t_L g349 ( .A(n_292), .Y(n_349) );
OR2x6_ASAP7_75t_L g350 ( .A(n_299), .B(n_232), .Y(n_350) );
INVx2_ASAP7_75t_L g351 ( .A(n_292), .Y(n_351) );
INVx2_ASAP7_75t_L g352 ( .A(n_292), .Y(n_352) );
INVx1_ASAP7_75t_L g353 ( .A(n_290), .Y(n_353) );
INVx2_ASAP7_75t_L g354 ( .A(n_292), .Y(n_354) );
AND2x6_ASAP7_75t_L g355 ( .A(n_307), .B(n_200), .Y(n_355) );
NAND2xp5_ASAP7_75t_L g356 ( .A(n_337), .B(n_186), .Y(n_356) );
BUFx12f_ASAP7_75t_L g357 ( .A(n_340), .Y(n_357) );
INVx1_ASAP7_75t_L g358 ( .A(n_339), .Y(n_358) );
OR2x6_ASAP7_75t_L g359 ( .A(n_327), .B(n_304), .Y(n_359) );
INVx1_ASAP7_75t_SL g360 ( .A(n_334), .Y(n_360) );
OAI22xp5_ASAP7_75t_SL g361 ( .A1(n_321), .A2(n_257), .B1(n_267), .B2(n_255), .Y(n_361) );
NAND2xp5_ASAP7_75t_L g362 ( .A(n_327), .B(n_194), .Y(n_362) );
NAND2xp5_ASAP7_75t_L g363 ( .A(n_343), .B(n_195), .Y(n_363) );
NAND2xp5_ASAP7_75t_L g364 ( .A(n_331), .B(n_195), .Y(n_364) );
INVx1_ASAP7_75t_L g365 ( .A(n_339), .Y(n_365) );
NOR2xp33_ASAP7_75t_L g366 ( .A(n_328), .B(n_221), .Y(n_366) );
NAND2xp5_ASAP7_75t_L g367 ( .A(n_338), .B(n_243), .Y(n_367) );
INVx2_ASAP7_75t_L g368 ( .A(n_353), .Y(n_368) );
INVx2_ASAP7_75t_L g369 ( .A(n_353), .Y(n_369) );
NAND2xp5_ASAP7_75t_L g370 ( .A(n_330), .B(n_286), .Y(n_370) );
NAND2xp5_ASAP7_75t_L g371 ( .A(n_330), .B(n_286), .Y(n_371) );
INVx2_ASAP7_75t_L g372 ( .A(n_322), .Y(n_372) );
AOI22xp5_ASAP7_75t_L g373 ( .A1(n_355), .A2(n_330), .B1(n_348), .B2(n_350), .Y(n_373) );
CKINVDCx5p33_ASAP7_75t_R g374 ( .A(n_340), .Y(n_374) );
INVx2_ASAP7_75t_L g375 ( .A(n_322), .Y(n_375) );
INVx2_ASAP7_75t_SL g376 ( .A(n_340), .Y(n_376) );
CKINVDCx5p33_ASAP7_75t_R g377 ( .A(n_321), .Y(n_377) );
INVx2_ASAP7_75t_L g378 ( .A(n_322), .Y(n_378) );
CKINVDCx5p33_ASAP7_75t_R g379 ( .A(n_345), .Y(n_379) );
OAI22xp33_ASAP7_75t_L g380 ( .A1(n_350), .A2(n_257), .B1(n_268), .B2(n_267), .Y(n_380) );
INVx2_ASAP7_75t_L g381 ( .A(n_324), .Y(n_381) );
INVx2_ASAP7_75t_L g382 ( .A(n_324), .Y(n_382) );
BUFx3_ASAP7_75t_L g383 ( .A(n_324), .Y(n_383) );
BUFx3_ASAP7_75t_L g384 ( .A(n_325), .Y(n_384) );
INVx2_ASAP7_75t_L g385 ( .A(n_325), .Y(n_385) );
INVx2_ASAP7_75t_L g386 ( .A(n_325), .Y(n_386) );
NAND2xp5_ASAP7_75t_L g387 ( .A(n_332), .B(n_276), .Y(n_387) );
CKINVDCx5p33_ASAP7_75t_R g388 ( .A(n_355), .Y(n_388) );
AO22x1_ASAP7_75t_L g389 ( .A1(n_355), .A2(n_298), .B1(n_293), .B2(n_202), .Y(n_389) );
BUFx6f_ASAP7_75t_L g390 ( .A(n_342), .Y(n_390) );
INVx2_ASAP7_75t_L g391 ( .A(n_323), .Y(n_391) );
INVx1_ASAP7_75t_L g392 ( .A(n_350), .Y(n_392) );
NAND2xp5_ASAP7_75t_SL g393 ( .A(n_347), .B(n_281), .Y(n_393) );
INVx1_ASAP7_75t_L g394 ( .A(n_350), .Y(n_394) );
INVx3_ASAP7_75t_L g395 ( .A(n_350), .Y(n_395) );
INVx2_ASAP7_75t_L g396 ( .A(n_323), .Y(n_396) );
NAND2xp5_ASAP7_75t_SL g397 ( .A(n_347), .B(n_197), .Y(n_397) );
NAND2xp5_ASAP7_75t_SL g398 ( .A(n_347), .B(n_207), .Y(n_398) );
BUFx6f_ASAP7_75t_SL g399 ( .A(n_355), .Y(n_399) );
NAND2xp5_ASAP7_75t_L g400 ( .A(n_332), .B(n_274), .Y(n_400) );
AOI22xp33_ASAP7_75t_L g401 ( .A1(n_355), .A2(n_298), .B1(n_228), .B2(n_233), .Y(n_401) );
NAND2xp5_ASAP7_75t_L g402 ( .A(n_326), .B(n_274), .Y(n_402) );
BUFx6f_ASAP7_75t_L g403 ( .A(n_390), .Y(n_403) );
AOI22xp5_ASAP7_75t_L g404 ( .A1(n_360), .A2(n_192), .B1(n_270), .B2(n_264), .Y(n_404) );
AOI21x1_ASAP7_75t_L g405 ( .A1(n_389), .A2(n_335), .B(n_311), .Y(n_405) );
INVx1_ASAP7_75t_SL g406 ( .A(n_358), .Y(n_406) );
OAI22xp5_ASAP7_75t_L g407 ( .A1(n_365), .A2(n_270), .B1(n_264), .B2(n_346), .Y(n_407) );
OAI22xp5_ASAP7_75t_L g408 ( .A1(n_365), .A2(n_282), .B1(n_268), .B2(n_308), .Y(n_408) );
O2A1O1Ixp5_ASAP7_75t_L g409 ( .A1(n_389), .A2(n_336), .B(n_344), .C(n_278), .Y(n_409) );
OR2x6_ASAP7_75t_L g410 ( .A(n_357), .B(n_320), .Y(n_410) );
AOI22xp33_ASAP7_75t_SL g411 ( .A1(n_379), .A2(n_226), .B1(n_235), .B2(n_209), .Y(n_411) );
HB1xp67_ASAP7_75t_L g412 ( .A(n_357), .Y(n_412) );
OAI22xp5_ASAP7_75t_L g413 ( .A1(n_388), .A2(n_245), .B1(n_253), .B2(n_220), .Y(n_413) );
OAI22xp5_ASAP7_75t_SL g414 ( .A1(n_361), .A2(n_238), .B1(n_240), .B2(n_239), .Y(n_414) );
INVx4_ASAP7_75t_SL g415 ( .A(n_399), .Y(n_415) );
OR2x2_ASAP7_75t_L g416 ( .A(n_380), .B(n_224), .Y(n_416) );
A2O1A1Ixp33_ASAP7_75t_L g417 ( .A1(n_400), .A2(n_344), .B(n_262), .C(n_265), .Y(n_417) );
INVx4_ASAP7_75t_L g418 ( .A(n_374), .Y(n_418) );
NAND2xp5_ASAP7_75t_SL g419 ( .A(n_374), .B(n_213), .Y(n_419) );
OAI22xp5_ASAP7_75t_L g420 ( .A1(n_388), .A2(n_271), .B1(n_275), .B2(n_256), .Y(n_420) );
BUFx6f_ASAP7_75t_L g421 ( .A(n_390), .Y(n_421) );
NAND2xp5_ASAP7_75t_L g422 ( .A(n_356), .B(n_273), .Y(n_422) );
INVx1_ASAP7_75t_L g423 ( .A(n_402), .Y(n_423) );
INVx2_ASAP7_75t_L g424 ( .A(n_372), .Y(n_424) );
NAND2xp5_ASAP7_75t_L g425 ( .A(n_362), .B(n_280), .Y(n_425) );
AOI21xp5_ASAP7_75t_L g426 ( .A1(n_359), .A2(n_201), .B(n_198), .Y(n_426) );
A2O1A1Ixp33_ASAP7_75t_L g427 ( .A1(n_373), .A2(n_283), .B(n_199), .C(n_205), .Y(n_427) );
NAND2xp5_ASAP7_75t_SL g428 ( .A(n_376), .B(n_190), .Y(n_428) );
A2O1A1Ixp33_ASAP7_75t_L g429 ( .A1(n_395), .A2(n_212), .B(n_214), .C(n_211), .Y(n_429) );
A2O1A1Ixp33_ASAP7_75t_L g430 ( .A1(n_395), .A2(n_217), .B(n_219), .C(n_215), .Y(n_430) );
NAND2xp5_ASAP7_75t_L g431 ( .A(n_363), .B(n_298), .Y(n_431) );
INVx2_ASAP7_75t_SL g432 ( .A(n_392), .Y(n_432) );
INVx2_ASAP7_75t_L g433 ( .A(n_372), .Y(n_433) );
AOI22xp33_ASAP7_75t_L g434 ( .A1(n_399), .A2(n_298), .B1(n_218), .B2(n_223), .Y(n_434) );
O2A1O1Ixp33_ASAP7_75t_L g435 ( .A1(n_364), .A2(n_222), .B(n_230), .C(n_227), .Y(n_435) );
BUFx6f_ASAP7_75t_L g436 ( .A(n_390), .Y(n_436) );
NOR2xp33_ASAP7_75t_L g437 ( .A(n_366), .B(n_231), .Y(n_437) );
AOI21xp5_ASAP7_75t_L g438 ( .A1(n_359), .A2(n_398), .B(n_397), .Y(n_438) );
NAND2xp5_ASAP7_75t_SL g439 ( .A(n_376), .B(n_237), .Y(n_439) );
BUFx3_ASAP7_75t_L g440 ( .A(n_394), .Y(n_440) );
NOR3xp33_ASAP7_75t_SL g441 ( .A(n_377), .B(n_247), .C(n_246), .Y(n_441) );
OAI22xp5_ASAP7_75t_L g442 ( .A1(n_399), .A2(n_248), .B1(n_252), .B2(n_250), .Y(n_442) );
NOR2xp33_ASAP7_75t_L g443 ( .A(n_367), .B(n_254), .Y(n_443) );
INVx2_ASAP7_75t_L g444 ( .A(n_375), .Y(n_444) );
BUFx6f_ASAP7_75t_SL g445 ( .A(n_383), .Y(n_445) );
O2A1O1Ixp33_ASAP7_75t_L g446 ( .A1(n_387), .A2(n_263), .B(n_269), .C(n_261), .Y(n_446) );
AND2x2_ASAP7_75t_L g447 ( .A(n_368), .B(n_10), .Y(n_447) );
HB1xp67_ASAP7_75t_L g448 ( .A(n_370), .Y(n_448) );
BUFx12f_ASAP7_75t_L g449 ( .A(n_390), .Y(n_449) );
OAI22xp5_ASAP7_75t_L g450 ( .A1(n_401), .A2(n_285), .B1(n_229), .B2(n_242), .Y(n_450) );
BUFx6f_ASAP7_75t_L g451 ( .A(n_383), .Y(n_451) );
NOR2xp33_ASAP7_75t_L g452 ( .A(n_371), .B(n_10), .Y(n_452) );
INVx4_ASAP7_75t_L g453 ( .A(n_384), .Y(n_453) );
NAND2xp5_ASAP7_75t_L g454 ( .A(n_369), .B(n_236), .Y(n_454) );
INVx2_ASAP7_75t_L g455 ( .A(n_378), .Y(n_455) );
A2O1A1Ixp33_ASAP7_75t_L g456 ( .A1(n_378), .A2(n_258), .B(n_266), .C(n_236), .Y(n_456) );
INVx4_ASAP7_75t_L g457 ( .A(n_381), .Y(n_457) );
INVx1_ASAP7_75t_L g458 ( .A(n_382), .Y(n_458) );
INVx5_ASAP7_75t_L g459 ( .A(n_382), .Y(n_459) );
OAI22xp5_ASAP7_75t_L g460 ( .A1(n_385), .A2(n_284), .B1(n_251), .B2(n_294), .Y(n_460) );
NOR2xp33_ASAP7_75t_L g461 ( .A(n_393), .B(n_14), .Y(n_461) );
NAND2xp5_ASAP7_75t_L g462 ( .A(n_385), .B(n_14), .Y(n_462) );
NAND2xp33_ASAP7_75t_R g463 ( .A(n_386), .B(n_15), .Y(n_463) );
A2O1A1Ixp33_ASAP7_75t_L g464 ( .A1(n_391), .A2(n_305), .B(n_290), .C(n_301), .Y(n_464) );
A2O1A1Ixp33_ASAP7_75t_L g465 ( .A1(n_391), .A2(n_305), .B(n_290), .C(n_301), .Y(n_465) );
OA21x2_ASAP7_75t_L g466 ( .A1(n_396), .A2(n_333), .B(n_329), .Y(n_466) );
BUFx4f_ASAP7_75t_SL g467 ( .A(n_396), .Y(n_467) );
CKINVDCx20_ASAP7_75t_R g468 ( .A(n_360), .Y(n_468) );
AOI21xp5_ASAP7_75t_L g469 ( .A1(n_431), .A2(n_354), .B(n_333), .Y(n_469) );
O2A1O1Ixp33_ASAP7_75t_L g470 ( .A1(n_429), .A2(n_354), .B(n_352), .C(n_351), .Y(n_470) );
O2A1O1Ixp33_ASAP7_75t_L g471 ( .A1(n_430), .A2(n_354), .B(n_352), .C(n_351), .Y(n_471) );
BUFx2_ASAP7_75t_L g472 ( .A(n_468), .Y(n_472) );
AOI22xp33_ASAP7_75t_L g473 ( .A1(n_408), .A2(n_317), .B1(n_303), .B2(n_296), .Y(n_473) );
A2O1A1Ixp33_ASAP7_75t_L g474 ( .A1(n_443), .A2(n_317), .B(n_303), .C(n_296), .Y(n_474) );
O2A1O1Ixp33_ASAP7_75t_L g475 ( .A1(n_417), .A2(n_17), .B(n_18), .C(n_19), .Y(n_475) );
INVx1_ASAP7_75t_L g476 ( .A(n_447), .Y(n_476) );
INVx5_ASAP7_75t_L g477 ( .A(n_449), .Y(n_477) );
BUFx6f_ASAP7_75t_L g478 ( .A(n_403), .Y(n_478) );
INVx3_ASAP7_75t_L g479 ( .A(n_453), .Y(n_479) );
OAI21xp5_ASAP7_75t_L g480 ( .A1(n_409), .A2(n_317), .B(n_75), .Y(n_480) );
AO31x2_ASAP7_75t_L g481 ( .A1(n_456), .A2(n_317), .A3(n_349), .B(n_341), .Y(n_481) );
INVx4_ASAP7_75t_L g482 ( .A(n_418), .Y(n_482) );
A2O1A1Ixp33_ASAP7_75t_L g483 ( .A1(n_435), .A2(n_349), .B(n_341), .C(n_21), .Y(n_483) );
AO31x2_ASAP7_75t_L g484 ( .A1(n_427), .A2(n_349), .A3(n_341), .B(n_22), .Y(n_484) );
A2O1A1Ixp33_ASAP7_75t_L g485 ( .A1(n_446), .A2(n_349), .B(n_341), .C(n_22), .Y(n_485) );
OAI21x1_ASAP7_75t_L g486 ( .A1(n_405), .A2(n_76), .B(n_73), .Y(n_486) );
AOI22xp33_ASAP7_75t_L g487 ( .A1(n_410), .A2(n_349), .B1(n_341), .B2(n_23), .Y(n_487) );
HB1xp67_ASAP7_75t_L g488 ( .A(n_463), .Y(n_488) );
BUFx6f_ASAP7_75t_L g489 ( .A(n_403), .Y(n_489) );
AO32x2_ASAP7_75t_L g490 ( .A1(n_442), .A2(n_25), .A3(n_26), .B1(n_27), .B2(n_28), .Y(n_490) );
AO31x2_ASAP7_75t_L g491 ( .A1(n_426), .A2(n_27), .A3(n_28), .B(n_30), .Y(n_491) );
A2O1A1Ixp33_ASAP7_75t_L g492 ( .A1(n_437), .A2(n_33), .B(n_35), .C(n_36), .Y(n_492) );
A2O1A1Ixp33_ASAP7_75t_L g493 ( .A1(n_452), .A2(n_38), .B(n_39), .C(n_40), .Y(n_493) );
AO32x2_ASAP7_75t_L g494 ( .A1(n_442), .A2(n_42), .A3(n_43), .B1(n_44), .B2(n_45), .Y(n_494) );
BUFx3_ASAP7_75t_L g495 ( .A(n_412), .Y(n_495) );
AO32x2_ASAP7_75t_L g496 ( .A1(n_450), .A2(n_47), .A3(n_48), .B1(n_49), .B2(n_50), .Y(n_496) );
INVx2_ASAP7_75t_L g497 ( .A(n_424), .Y(n_497) );
A2O1A1Ixp33_ASAP7_75t_L g498 ( .A1(n_461), .A2(n_49), .B(n_50), .C(n_51), .Y(n_498) );
AOI221x1_ASAP7_75t_L g499 ( .A1(n_438), .A2(n_52), .B1(n_53), .B2(n_54), .C(n_56), .Y(n_499) );
INVx1_ASAP7_75t_L g500 ( .A(n_423), .Y(n_500) );
INVx2_ASAP7_75t_SL g501 ( .A(n_467), .Y(n_501) );
INVx1_ASAP7_75t_SL g502 ( .A(n_416), .Y(n_502) );
AO31x2_ASAP7_75t_L g503 ( .A1(n_460), .A2(n_57), .A3(n_58), .B(n_59), .Y(n_503) );
OR2x2_ASAP7_75t_L g504 ( .A(n_425), .B(n_78), .Y(n_504) );
OA21x2_ASAP7_75t_L g505 ( .A1(n_464), .A2(n_79), .B(n_80), .Y(n_505) );
INVxp67_ASAP7_75t_SL g506 ( .A(n_451), .Y(n_506) );
AO31x2_ASAP7_75t_L g507 ( .A1(n_460), .A2(n_81), .A3(n_83), .B(n_86), .Y(n_507) );
NAND2xp5_ASAP7_75t_L g508 ( .A(n_422), .B(n_88), .Y(n_508) );
OAI21x1_ASAP7_75t_L g509 ( .A1(n_466), .A2(n_90), .B(n_91), .Y(n_509) );
BUFx10_ASAP7_75t_L g510 ( .A(n_445), .Y(n_510) );
INVxp67_ASAP7_75t_L g511 ( .A(n_413), .Y(n_511) );
AO31x2_ASAP7_75t_L g512 ( .A1(n_450), .A2(n_93), .A3(n_94), .B(n_96), .Y(n_512) );
INVx1_ASAP7_75t_L g513 ( .A(n_458), .Y(n_513) );
OAI21x1_ASAP7_75t_L g514 ( .A1(n_466), .A2(n_99), .B(n_100), .Y(n_514) );
OAI21x1_ASAP7_75t_L g515 ( .A1(n_462), .A2(n_102), .B(n_104), .Y(n_515) );
INVx1_ASAP7_75t_L g516 ( .A(n_440), .Y(n_516) );
O2A1O1Ixp33_ASAP7_75t_L g517 ( .A1(n_420), .A2(n_105), .B(n_107), .C(n_108), .Y(n_517) );
BUFx6f_ASAP7_75t_L g518 ( .A(n_403), .Y(n_518) );
HB1xp67_ASAP7_75t_L g519 ( .A(n_451), .Y(n_519) );
AOI21xp5_ASAP7_75t_L g520 ( .A1(n_428), .A2(n_110), .B(n_111), .Y(n_520) );
INVx1_ASAP7_75t_L g521 ( .A(n_454), .Y(n_521) );
O2A1O1Ixp33_ASAP7_75t_SL g522 ( .A1(n_465), .A2(n_112), .B(n_117), .C(n_118), .Y(n_522) );
AND2x4_ASAP7_75t_L g523 ( .A(n_415), .B(n_432), .Y(n_523) );
AOI21xp5_ASAP7_75t_L g524 ( .A1(n_439), .A2(n_121), .B(n_122), .Y(n_524) );
AOI22xp33_ASAP7_75t_L g525 ( .A1(n_448), .A2(n_130), .B1(n_131), .B2(n_132), .Y(n_525) );
AND2x4_ASAP7_75t_L g526 ( .A(n_415), .B(n_134), .Y(n_526) );
INVx2_ASAP7_75t_L g527 ( .A(n_433), .Y(n_527) );
O2A1O1Ixp33_ASAP7_75t_L g528 ( .A1(n_419), .A2(n_135), .B(n_138), .C(n_139), .Y(n_528) );
BUFx2_ASAP7_75t_L g529 ( .A(n_421), .Y(n_529) );
OR2x6_ASAP7_75t_L g530 ( .A(n_421), .B(n_140), .Y(n_530) );
NOR2xp33_ASAP7_75t_SL g531 ( .A(n_436), .B(n_141), .Y(n_531) );
A2O1A1Ixp33_ASAP7_75t_SL g532 ( .A1(n_434), .A2(n_143), .B(n_144), .C(n_145), .Y(n_532) );
OR2x6_ASAP7_75t_L g533 ( .A(n_530), .B(n_436), .Y(n_533) );
OAI21xp5_ASAP7_75t_L g534 ( .A1(n_480), .A2(n_455), .B(n_444), .Y(n_534) );
AOI21xp5_ASAP7_75t_L g535 ( .A1(n_508), .A2(n_457), .B(n_459), .Y(n_535) );
BUFx8_ASAP7_75t_L g536 ( .A(n_472), .Y(n_536) );
CKINVDCx11_ASAP7_75t_R g537 ( .A(n_510), .Y(n_537) );
OR2x6_ASAP7_75t_L g538 ( .A(n_482), .B(n_152), .Y(n_538) );
INVx4_ASAP7_75t_L g539 ( .A(n_477), .Y(n_539) );
OAI21xp5_ASAP7_75t_L g540 ( .A1(n_476), .A2(n_164), .B(n_165), .Y(n_540) );
AOI21xp5_ASAP7_75t_L g541 ( .A1(n_469), .A2(n_174), .B(n_176), .Y(n_541) );
OAI22xp5_ASAP7_75t_L g542 ( .A1(n_513), .A2(n_473), .B1(n_504), .B2(n_487), .Y(n_542) );
INVx3_ASAP7_75t_L g543 ( .A(n_482), .Y(n_543) );
OA21x2_ASAP7_75t_L g544 ( .A1(n_486), .A2(n_514), .B(n_509), .Y(n_544) );
OA21x2_ASAP7_75t_L g545 ( .A1(n_515), .A2(n_499), .B(n_474), .Y(n_545) );
BUFx6f_ASAP7_75t_L g546 ( .A(n_478), .Y(n_546) );
OAI21xp5_ASAP7_75t_L g547 ( .A1(n_485), .A2(n_483), .B(n_521), .Y(n_547) );
INVx2_ASAP7_75t_L g548 ( .A(n_497), .Y(n_548) );
INVx2_ASAP7_75t_L g549 ( .A(n_527), .Y(n_549) );
INVx2_ASAP7_75t_L g550 ( .A(n_481), .Y(n_550) );
INVx2_ASAP7_75t_L g551 ( .A(n_481), .Y(n_551) );
OAI21xp5_ASAP7_75t_L g552 ( .A1(n_470), .A2(n_471), .B(n_475), .Y(n_552) );
INVx1_ASAP7_75t_SL g553 ( .A(n_529), .Y(n_553) );
OR2x6_ASAP7_75t_L g554 ( .A(n_501), .B(n_526), .Y(n_554) );
NAND2xp5_ASAP7_75t_L g555 ( .A(n_516), .B(n_479), .Y(n_555) );
NAND2xp5_ASAP7_75t_L g556 ( .A(n_479), .B(n_519), .Y(n_556) );
NAND2xp5_ASAP7_75t_L g557 ( .A(n_523), .B(n_492), .Y(n_557) );
CKINVDCx11_ASAP7_75t_R g558 ( .A(n_495), .Y(n_558) );
BUFx8_ASAP7_75t_L g559 ( .A(n_490), .Y(n_559) );
A2O1A1Ixp33_ASAP7_75t_L g560 ( .A1(n_517), .A2(n_493), .B(n_498), .C(n_528), .Y(n_560) );
NAND2xp5_ASAP7_75t_L g561 ( .A(n_506), .B(n_491), .Y(n_561) );
OA21x2_ASAP7_75t_L g562 ( .A1(n_525), .A2(n_524), .B(n_520), .Y(n_562) );
AOI21xp5_ASAP7_75t_L g563 ( .A1(n_532), .A2(n_522), .B(n_505), .Y(n_563) );
NAND2xp5_ASAP7_75t_L g564 ( .A(n_503), .B(n_489), .Y(n_564) );
OAI22xp33_ASAP7_75t_L g565 ( .A1(n_531), .A2(n_518), .B1(n_494), .B2(n_505), .Y(n_565) );
AOI21xp5_ASAP7_75t_L g566 ( .A1(n_518), .A2(n_512), .B(n_507), .Y(n_566) );
OAI22xp33_ASAP7_75t_L g567 ( .A1(n_518), .A2(n_496), .B1(n_503), .B2(n_512), .Y(n_567) );
AOI21xp5_ASAP7_75t_L g568 ( .A1(n_512), .A2(n_507), .B(n_484), .Y(n_568) );
OR2x2_ASAP7_75t_L g569 ( .A(n_484), .B(n_507), .Y(n_569) );
OAI21xp5_ASAP7_75t_L g570 ( .A1(n_484), .A2(n_409), .B(n_417), .Y(n_570) );
INVx2_ASAP7_75t_L g571 ( .A(n_500), .Y(n_571) );
AOI22xp33_ASAP7_75t_SL g572 ( .A1(n_488), .A2(n_468), .B1(n_408), .B2(n_361), .Y(n_572) );
OAI22xp33_ASAP7_75t_L g573 ( .A1(n_511), .A2(n_404), .B1(n_407), .B2(n_410), .Y(n_573) );
OAI221xp5_ASAP7_75t_L g574 ( .A1(n_502), .A2(n_360), .B1(n_441), .B2(n_408), .C(n_411), .Y(n_574) );
NAND2x1_ASAP7_75t_L g575 ( .A(n_530), .B(n_526), .Y(n_575) );
INVx2_ASAP7_75t_L g576 ( .A(n_500), .Y(n_576) );
NAND2xp5_ASAP7_75t_L g577 ( .A(n_511), .B(n_406), .Y(n_577) );
NAND2xp5_ASAP7_75t_L g578 ( .A(n_511), .B(n_406), .Y(n_578) );
AO21x2_ASAP7_75t_L g579 ( .A1(n_568), .A2(n_567), .B(n_566), .Y(n_579) );
OAI222xp33_ASAP7_75t_L g580 ( .A1(n_554), .A2(n_538), .B1(n_573), .B2(n_572), .C1(n_575), .C2(n_574), .Y(n_580) );
AND2x2_ASAP7_75t_L g581 ( .A(n_571), .B(n_576), .Y(n_581) );
OR2x2_ASAP7_75t_L g582 ( .A(n_577), .B(n_578), .Y(n_582) );
AND2x2_ASAP7_75t_L g583 ( .A(n_548), .B(n_549), .Y(n_583) );
AO21x2_ASAP7_75t_L g584 ( .A1(n_565), .A2(n_564), .B(n_563), .Y(n_584) );
INVx2_ASAP7_75t_L g585 ( .A(n_551), .Y(n_585) );
INVx6_ASAP7_75t_L g586 ( .A(n_539), .Y(n_586) );
OAI21xp5_ASAP7_75t_L g587 ( .A1(n_560), .A2(n_542), .B(n_547), .Y(n_587) );
AOI21xp5_ASAP7_75t_SL g588 ( .A1(n_538), .A2(n_533), .B(n_554), .Y(n_588) );
INVx3_ASAP7_75t_L g589 ( .A(n_533), .Y(n_589) );
AND2x4_ASAP7_75t_L g590 ( .A(n_546), .B(n_557), .Y(n_590) );
AND2x4_ASAP7_75t_L g591 ( .A(n_543), .B(n_540), .Y(n_591) );
INVxp67_ASAP7_75t_SL g592 ( .A(n_556), .Y(n_592) );
OA21x2_ASAP7_75t_L g593 ( .A1(n_569), .A2(n_561), .B(n_534), .Y(n_593) );
INVx1_ASAP7_75t_L g594 ( .A(n_559), .Y(n_594) );
INVx1_ASAP7_75t_L g595 ( .A(n_559), .Y(n_595) );
AND2x4_ASAP7_75t_L g596 ( .A(n_556), .B(n_553), .Y(n_596) );
AND2x4_ASAP7_75t_L g597 ( .A(n_555), .B(n_570), .Y(n_597) );
BUFx3_ASAP7_75t_L g598 ( .A(n_558), .Y(n_598) );
INVx1_ASAP7_75t_L g599 ( .A(n_545), .Y(n_599) );
INVx5_ASAP7_75t_L g600 ( .A(n_537), .Y(n_600) );
AND2x4_ASAP7_75t_L g601 ( .A(n_552), .B(n_535), .Y(n_601) );
INVx4_ASAP7_75t_L g602 ( .A(n_544), .Y(n_602) );
OAI332xp33_ASAP7_75t_L g603 ( .A1(n_536), .A2(n_408), .A3(n_361), .B1(n_574), .B2(n_502), .B3(n_380), .C1(n_414), .C2(n_573), .Y(n_603) );
AO21x2_ASAP7_75t_L g604 ( .A1(n_541), .A2(n_562), .B(n_536), .Y(n_604) );
INVx2_ASAP7_75t_L g605 ( .A(n_550), .Y(n_605) );
INVx3_ASAP7_75t_L g606 ( .A(n_533), .Y(n_606) );
OA21x2_ASAP7_75t_L g607 ( .A1(n_568), .A2(n_566), .B(n_564), .Y(n_607) );
AND2x2_ASAP7_75t_L g608 ( .A(n_571), .B(n_576), .Y(n_608) );
OA21x2_ASAP7_75t_L g609 ( .A1(n_568), .A2(n_566), .B(n_564), .Y(n_609) );
AND2x4_ASAP7_75t_L g610 ( .A(n_554), .B(n_538), .Y(n_610) );
AND2x2_ASAP7_75t_L g611 ( .A(n_597), .B(n_581), .Y(n_611) );
OR2x2_ASAP7_75t_SL g612 ( .A(n_594), .B(n_595), .Y(n_612) );
AND2x4_ASAP7_75t_L g613 ( .A(n_610), .B(n_594), .Y(n_613) );
OR2x2_ASAP7_75t_L g614 ( .A(n_592), .B(n_595), .Y(n_614) );
CKINVDCx8_ASAP7_75t_R g615 ( .A(n_600), .Y(n_615) );
AND2x2_ASAP7_75t_L g616 ( .A(n_608), .B(n_587), .Y(n_616) );
INVx3_ASAP7_75t_L g617 ( .A(n_591), .Y(n_617) );
INVx1_ASAP7_75t_L g618 ( .A(n_585), .Y(n_618) );
INVx1_ASAP7_75t_L g619 ( .A(n_585), .Y(n_619) );
INVx1_ASAP7_75t_L g620 ( .A(n_605), .Y(n_620) );
NOR2x1_ASAP7_75t_L g621 ( .A(n_588), .B(n_598), .Y(n_621) );
INVx4_ASAP7_75t_L g622 ( .A(n_586), .Y(n_622) );
OR2x2_ASAP7_75t_L g623 ( .A(n_582), .B(n_596), .Y(n_623) );
BUFx3_ASAP7_75t_L g624 ( .A(n_586), .Y(n_624) );
NAND2xp5_ASAP7_75t_L g625 ( .A(n_583), .B(n_603), .Y(n_625) );
INVx3_ASAP7_75t_L g626 ( .A(n_591), .Y(n_626) );
INVx2_ASAP7_75t_L g627 ( .A(n_602), .Y(n_627) );
INVx4_ASAP7_75t_L g628 ( .A(n_589), .Y(n_628) );
AND2x2_ASAP7_75t_L g629 ( .A(n_601), .B(n_593), .Y(n_629) );
INVx1_ASAP7_75t_L g630 ( .A(n_599), .Y(n_630) );
INVx4_ASAP7_75t_L g631 ( .A(n_589), .Y(n_631) );
INVx1_ASAP7_75t_L g632 ( .A(n_630), .Y(n_632) );
AND2x2_ASAP7_75t_L g633 ( .A(n_611), .B(n_609), .Y(n_633) );
OR2x2_ASAP7_75t_L g634 ( .A(n_623), .B(n_609), .Y(n_634) );
AND2x4_ASAP7_75t_L g635 ( .A(n_617), .B(n_579), .Y(n_635) );
OR2x2_ASAP7_75t_L g636 ( .A(n_623), .B(n_607), .Y(n_636) );
AND2x2_ASAP7_75t_L g637 ( .A(n_629), .B(n_607), .Y(n_637) );
AND2x4_ASAP7_75t_L g638 ( .A(n_617), .B(n_579), .Y(n_638) );
AND2x4_ASAP7_75t_L g639 ( .A(n_617), .B(n_579), .Y(n_639) );
INVx1_ASAP7_75t_L g640 ( .A(n_618), .Y(n_640) );
INVx1_ASAP7_75t_L g641 ( .A(n_619), .Y(n_641) );
AND2x2_ASAP7_75t_L g642 ( .A(n_616), .B(n_590), .Y(n_642) );
CKINVDCx16_ASAP7_75t_R g643 ( .A(n_621), .Y(n_643) );
AND2x4_ASAP7_75t_SL g644 ( .A(n_622), .B(n_606), .Y(n_644) );
AND2x6_ASAP7_75t_SL g645 ( .A(n_625), .B(n_580), .Y(n_645) );
BUFx3_ASAP7_75t_L g646 ( .A(n_624), .Y(n_646) );
INVx1_ASAP7_75t_L g647 ( .A(n_619), .Y(n_647) );
INVx1_ASAP7_75t_L g648 ( .A(n_620), .Y(n_648) );
OR2x2_ASAP7_75t_L g649 ( .A(n_614), .B(n_584), .Y(n_649) );
AND2x4_ASAP7_75t_L g650 ( .A(n_626), .B(n_604), .Y(n_650) );
NAND2xp5_ASAP7_75t_SL g651 ( .A(n_643), .B(n_622), .Y(n_651) );
INVx1_ASAP7_75t_L g652 ( .A(n_632), .Y(n_652) );
INVx1_ASAP7_75t_L g653 ( .A(n_640), .Y(n_653) );
AND2x2_ASAP7_75t_L g654 ( .A(n_633), .B(n_627), .Y(n_654) );
INVx1_ASAP7_75t_L g655 ( .A(n_641), .Y(n_655) );
INVx1_ASAP7_75t_L g656 ( .A(n_641), .Y(n_656) );
INVx1_ASAP7_75t_L g657 ( .A(n_647), .Y(n_657) );
INVx1_ASAP7_75t_L g658 ( .A(n_648), .Y(n_658) );
NAND2x1_ASAP7_75t_L g659 ( .A(n_654), .B(n_650), .Y(n_659) );
INVx1_ASAP7_75t_L g660 ( .A(n_652), .Y(n_660) );
BUFx2_ASAP7_75t_L g661 ( .A(n_654), .Y(n_661) );
NAND2xp5_ASAP7_75t_SL g662 ( .A(n_651), .B(n_615), .Y(n_662) );
AND2x2_ASAP7_75t_L g663 ( .A(n_661), .B(n_637), .Y(n_663) );
INVx1_ASAP7_75t_L g664 ( .A(n_660), .Y(n_664) );
INVxp67_ASAP7_75t_SL g665 ( .A(n_659), .Y(n_665) );
AOI21xp5_ASAP7_75t_L g666 ( .A1(n_665), .A2(n_659), .B(n_662), .Y(n_666) );
OAI22xp5_ASAP7_75t_L g667 ( .A1(n_666), .A2(n_663), .B1(n_612), .B2(n_664), .Y(n_667) );
AOI211xp5_ASAP7_75t_L g668 ( .A1(n_667), .A2(n_613), .B(n_646), .C(n_645), .Y(n_668) );
AND2x2_ASAP7_75t_L g669 ( .A(n_668), .B(n_642), .Y(n_669) );
NOR2xp67_ASAP7_75t_L g670 ( .A(n_669), .B(n_628), .Y(n_670) );
OAI22xp5_ASAP7_75t_L g671 ( .A1(n_670), .A2(n_649), .B1(n_636), .B2(n_634), .Y(n_671) );
AOI22xp5_ASAP7_75t_L g672 ( .A1(n_671), .A2(n_644), .B1(n_638), .B2(n_635), .Y(n_672) );
AOI222xp33_ASAP7_75t_L g673 ( .A1(n_672), .A2(n_644), .B1(n_658), .B2(n_656), .C1(n_655), .C2(n_653), .Y(n_673) );
NAND2xp5_ASAP7_75t_L g674 ( .A(n_673), .B(n_657), .Y(n_674) );
INVx3_ASAP7_75t_L g675 ( .A(n_674), .Y(n_675) );
AOI222xp33_ASAP7_75t_L g676 ( .A1(n_675), .A2(n_631), .B1(n_650), .B2(n_635), .C1(n_638), .C2(n_639), .Y(n_676) );
endmodule