module fake_jpeg_11800_n_379 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_379);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_379;

wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_340;
wire n_377;
wire n_291;
wire n_236;
wire n_15;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_256;
wire n_221;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_370;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_368;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_39;
wire n_371;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_352;
wire n_350;
wire n_367;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_360;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_378;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_356;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_375;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVx3_ASAP7_75t_L g15 ( 
.A(n_14),
.Y(n_15)
);

BUFx10_ASAP7_75t_L g16 ( 
.A(n_2),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_9),
.Y(n_17)
);

INVx11_ASAP7_75t_L g18 ( 
.A(n_14),
.Y(n_18)
);

INVx8_ASAP7_75t_L g19 ( 
.A(n_2),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_2),
.Y(n_20)
);

BUFx3_ASAP7_75t_L g21 ( 
.A(n_12),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_2),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_8),
.Y(n_23)
);

BUFx12f_ASAP7_75t_L g24 ( 
.A(n_8),
.Y(n_24)
);

BUFx6f_ASAP7_75t_SL g25 ( 
.A(n_1),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_14),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_5),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_5),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_10),
.Y(n_29)
);

BUFx10_ASAP7_75t_L g30 ( 
.A(n_10),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_8),
.Y(n_31)
);

INVx2_ASAP7_75t_L g32 ( 
.A(n_13),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_3),
.Y(n_33)
);

BUFx5_ASAP7_75t_L g34 ( 
.A(n_9),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_17),
.Y(n_35)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_35),
.Y(n_63)
);

BUFx3_ASAP7_75t_L g36 ( 
.A(n_24),
.Y(n_36)
);

BUFx12f_ASAP7_75t_L g70 ( 
.A(n_36),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g37 ( 
.A(n_32),
.B(n_13),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_SL g80 ( 
.A(n_37),
.B(n_45),
.Y(n_80)
);

NAND2xp67_ASAP7_75t_L g38 ( 
.A(n_16),
.B(n_0),
.Y(n_38)
);

AND2x2_ASAP7_75t_L g88 ( 
.A(n_38),
.B(n_16),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_SL g39 ( 
.A(n_32),
.B(n_0),
.Y(n_39)
);

NAND2xp5_ASAP7_75t_L g81 ( 
.A(n_39),
.B(n_51),
.Y(n_81)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_17),
.Y(n_40)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_40),
.Y(n_78)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_28),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g74 ( 
.A(n_41),
.Y(n_74)
);

INVx5_ASAP7_75t_L g42 ( 
.A(n_19),
.Y(n_42)
);

INVx5_ASAP7_75t_L g67 ( 
.A(n_42),
.Y(n_67)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_17),
.Y(n_43)
);

INVx2_ASAP7_75t_L g68 ( 
.A(n_43),
.Y(n_68)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_28),
.Y(n_44)
);

INVx6_ASAP7_75t_L g62 ( 
.A(n_44),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g45 ( 
.A(n_32),
.B(n_13),
.Y(n_45)
);

INVx4_ASAP7_75t_L g46 ( 
.A(n_24),
.Y(n_46)
);

INVx3_ASAP7_75t_L g69 ( 
.A(n_46),
.Y(n_69)
);

INVx4_ASAP7_75t_L g47 ( 
.A(n_24),
.Y(n_47)
);

INVx3_ASAP7_75t_L g71 ( 
.A(n_47),
.Y(n_71)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_27),
.Y(n_48)
);

INVx2_ASAP7_75t_L g73 ( 
.A(n_48),
.Y(n_73)
);

INVx3_ASAP7_75t_L g49 ( 
.A(n_21),
.Y(n_49)
);

INVx3_ASAP7_75t_L g82 ( 
.A(n_49),
.Y(n_82)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_28),
.Y(n_50)
);

INVx5_ASAP7_75t_L g76 ( 
.A(n_50),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_L g51 ( 
.A(n_15),
.B(n_0),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_28),
.Y(n_52)
);

BUFx3_ASAP7_75t_L g66 ( 
.A(n_52),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_33),
.Y(n_53)
);

INVx3_ASAP7_75t_L g86 ( 
.A(n_53),
.Y(n_86)
);

INVx3_ASAP7_75t_L g54 ( 
.A(n_21),
.Y(n_54)
);

INVx2_ASAP7_75t_L g75 ( 
.A(n_54),
.Y(n_75)
);

INVx2_ASAP7_75t_L g55 ( 
.A(n_24),
.Y(n_55)
);

INVx2_ASAP7_75t_L g77 ( 
.A(n_55),
.Y(n_77)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_27),
.Y(n_56)
);

INVx2_ASAP7_75t_L g83 ( 
.A(n_56),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g57 ( 
.A(n_15),
.B(n_0),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_L g84 ( 
.A(n_57),
.B(n_1),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_37),
.B(n_15),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_58),
.B(n_59),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_45),
.B(n_20),
.Y(n_59)
);

OAI22xp5_ASAP7_75t_L g60 ( 
.A1(n_39),
.A2(n_26),
.B1(n_33),
.B2(n_21),
.Y(n_60)
);

AOI22xp5_ASAP7_75t_L g109 ( 
.A1(n_60),
.A2(n_72),
.B1(n_79),
.B2(n_16),
.Y(n_109)
);

CKINVDCx14_ASAP7_75t_R g61 ( 
.A(n_51),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g123 ( 
.A(n_61),
.B(n_64),
.Y(n_123)
);

CKINVDCx14_ASAP7_75t_R g64 ( 
.A(n_57),
.Y(n_64)
);

AOI22xp33_ASAP7_75t_SL g65 ( 
.A1(n_35),
.A2(n_19),
.B1(n_21),
.B2(n_25),
.Y(n_65)
);

AOI22xp33_ASAP7_75t_SL g96 ( 
.A1(n_65),
.A2(n_30),
.B1(n_16),
.B2(n_25),
.Y(n_96)
);

OAI22xp5_ASAP7_75t_L g72 ( 
.A1(n_41),
.A2(n_26),
.B1(n_33),
.B2(n_31),
.Y(n_72)
);

OAI22xp33_ASAP7_75t_L g79 ( 
.A1(n_41),
.A2(n_33),
.B1(n_25),
.B2(n_16),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_84),
.B(n_31),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_40),
.B(n_23),
.Y(n_85)
);

INVxp67_ASAP7_75t_L g90 ( 
.A(n_85),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_43),
.B(n_23),
.Y(n_87)
);

INVxp67_ASAP7_75t_L g113 ( 
.A(n_87),
.Y(n_113)
);

AND2x2_ASAP7_75t_L g93 ( 
.A(n_88),
.B(n_46),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_SL g132 ( 
.A(n_89),
.B(n_20),
.Y(n_132)
);

BUFx3_ASAP7_75t_L g91 ( 
.A(n_70),
.Y(n_91)
);

INVx4_ASAP7_75t_L g131 ( 
.A(n_91),
.Y(n_131)
);

CKINVDCx14_ASAP7_75t_R g92 ( 
.A(n_80),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g139 ( 
.A(n_92),
.B(n_97),
.Y(n_139)
);

AND2x2_ASAP7_75t_L g140 ( 
.A(n_93),
.B(n_118),
.Y(n_140)
);

INVx2_ASAP7_75t_L g94 ( 
.A(n_77),
.Y(n_94)
);

INVx2_ASAP7_75t_L g141 ( 
.A(n_94),
.Y(n_141)
);

OAI22xp5_ASAP7_75t_SL g95 ( 
.A1(n_81),
.A2(n_50),
.B1(n_53),
.B2(n_52),
.Y(n_95)
);

AOI22xp5_ASAP7_75t_L g125 ( 
.A1(n_95),
.A2(n_102),
.B1(n_117),
.B2(n_120),
.Y(n_125)
);

AOI22xp33_ASAP7_75t_SL g146 ( 
.A1(n_96),
.A2(n_36),
.B1(n_30),
.B2(n_16),
.Y(n_146)
);

CKINVDCx14_ASAP7_75t_R g97 ( 
.A(n_70),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g98 ( 
.A(n_81),
.B(n_38),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g133 ( 
.A(n_98),
.B(n_105),
.Y(n_133)
);

INVx2_ASAP7_75t_L g99 ( 
.A(n_77),
.Y(n_99)
);

INVx1_ASAP7_75t_SL g154 ( 
.A(n_99),
.Y(n_154)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_63),
.Y(n_101)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_101),
.Y(n_126)
);

OAI22xp5_ASAP7_75t_SL g102 ( 
.A1(n_84),
.A2(n_50),
.B1(n_53),
.B2(n_52),
.Y(n_102)
);

INVx1_ASAP7_75t_SL g103 ( 
.A(n_63),
.Y(n_103)
);

CKINVDCx14_ASAP7_75t_R g142 ( 
.A(n_103),
.Y(n_142)
);

HB1xp67_ASAP7_75t_L g104 ( 
.A(n_75),
.Y(n_104)
);

CKINVDCx16_ASAP7_75t_R g130 ( 
.A(n_104),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_L g105 ( 
.A(n_78),
.B(n_56),
.Y(n_105)
);

CKINVDCx20_ASAP7_75t_R g106 ( 
.A(n_78),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g151 ( 
.A(n_106),
.B(n_114),
.Y(n_151)
);

AOI22xp33_ASAP7_75t_L g107 ( 
.A1(n_79),
.A2(n_48),
.B1(n_44),
.B2(n_23),
.Y(n_107)
);

OAI22xp5_ASAP7_75t_L g129 ( 
.A1(n_107),
.A2(n_109),
.B1(n_86),
.B2(n_76),
.Y(n_129)
);

AOI22xp5_ASAP7_75t_SL g108 ( 
.A1(n_88),
.A2(n_54),
.B1(n_49),
.B2(n_18),
.Y(n_108)
);

CKINVDCx16_ASAP7_75t_R g137 ( 
.A(n_108),
.Y(n_137)
);

BUFx3_ASAP7_75t_L g110 ( 
.A(n_70),
.Y(n_110)
);

BUFx6f_ASAP7_75t_L g138 ( 
.A(n_110),
.Y(n_138)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_68),
.Y(n_111)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_111),
.Y(n_135)
);

BUFx3_ASAP7_75t_L g112 ( 
.A(n_70),
.Y(n_112)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_112),
.Y(n_145)
);

INVxp67_ASAP7_75t_L g114 ( 
.A(n_88),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g115 ( 
.A(n_68),
.B(n_55),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_L g134 ( 
.A(n_115),
.B(n_75),
.Y(n_134)
);

INVx4_ASAP7_75t_L g116 ( 
.A(n_69),
.Y(n_116)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_116),
.Y(n_148)
);

OAI22xp5_ASAP7_75t_SL g117 ( 
.A1(n_73),
.A2(n_44),
.B1(n_42),
.B2(n_26),
.Y(n_117)
);

INVx4_ASAP7_75t_SL g118 ( 
.A(n_74),
.Y(n_118)
);

BUFx2_ASAP7_75t_L g119 ( 
.A(n_76),
.Y(n_119)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_119),
.Y(n_156)
);

OAI22xp5_ASAP7_75t_L g120 ( 
.A1(n_62),
.A2(n_26),
.B1(n_30),
.B2(n_16),
.Y(n_120)
);

OAI22xp5_ASAP7_75t_SL g121 ( 
.A1(n_73),
.A2(n_47),
.B1(n_46),
.B2(n_36),
.Y(n_121)
);

AOI22xp5_ASAP7_75t_L g153 ( 
.A1(n_121),
.A2(n_30),
.B1(n_19),
.B2(n_18),
.Y(n_153)
);

INVx4_ASAP7_75t_L g122 ( 
.A(n_69),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_L g152 ( 
.A(n_122),
.B(n_71),
.Y(n_152)
);

AND2x2_ASAP7_75t_L g124 ( 
.A(n_83),
.B(n_47),
.Y(n_124)
);

CKINVDCx16_ASAP7_75t_R g150 ( 
.A(n_124),
.Y(n_150)
);

AOI21xp5_ASAP7_75t_L g127 ( 
.A1(n_114),
.A2(n_83),
.B(n_67),
.Y(n_127)
);

AOI21xp5_ASAP7_75t_L g170 ( 
.A1(n_127),
.A2(n_122),
.B(n_116),
.Y(n_170)
);

OAI22xp5_ASAP7_75t_SL g128 ( 
.A1(n_109),
.A2(n_86),
.B1(n_62),
.B2(n_74),
.Y(n_128)
);

AOI22xp5_ASAP7_75t_L g181 ( 
.A1(n_128),
.A2(n_129),
.B1(n_147),
.B2(n_149),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_SL g169 ( 
.A(n_132),
.B(n_143),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_L g179 ( 
.A(n_134),
.B(n_144),
.Y(n_179)
);

OAI21xp5_ASAP7_75t_L g136 ( 
.A1(n_105),
.A2(n_20),
.B(n_22),
.Y(n_136)
);

OAI21xp5_ASAP7_75t_L g183 ( 
.A1(n_136),
.A2(n_30),
.B(n_29),
.Y(n_183)
);

CKINVDCx20_ASAP7_75t_R g143 ( 
.A(n_124),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_L g144 ( 
.A(n_98),
.B(n_89),
.Y(n_144)
);

AOI22xp33_ASAP7_75t_SL g180 ( 
.A1(n_146),
.A2(n_119),
.B1(n_121),
.B2(n_30),
.Y(n_180)
);

OAI22xp5_ASAP7_75t_SL g147 ( 
.A1(n_108),
.A2(n_82),
.B1(n_66),
.B2(n_67),
.Y(n_147)
);

OAI22xp5_ASAP7_75t_SL g149 ( 
.A1(n_123),
.A2(n_82),
.B1(n_66),
.B2(n_71),
.Y(n_149)
);

HB1xp67_ASAP7_75t_L g168 ( 
.A(n_152),
.Y(n_168)
);

OA22x2_ASAP7_75t_L g164 ( 
.A1(n_153),
.A2(n_22),
.B1(n_111),
.B2(n_103),
.Y(n_164)
);

AOI22xp33_ASAP7_75t_L g155 ( 
.A1(n_117),
.A2(n_31),
.B1(n_22),
.B2(n_27),
.Y(n_155)
);

OAI22xp5_ASAP7_75t_L g193 ( 
.A1(n_155),
.A2(n_34),
.B1(n_3),
.B2(n_4),
.Y(n_193)
);

OAI22xp5_ASAP7_75t_L g157 ( 
.A1(n_100),
.A2(n_30),
.B1(n_19),
.B2(n_18),
.Y(n_157)
);

AOI22xp5_ASAP7_75t_L g190 ( 
.A1(n_157),
.A2(n_112),
.B1(n_91),
.B2(n_24),
.Y(n_190)
);

NOR2xp33_ASAP7_75t_SL g158 ( 
.A(n_139),
.B(n_100),
.Y(n_158)
);

NOR2xp33_ASAP7_75t_L g209 ( 
.A(n_158),
.B(n_172),
.Y(n_209)
);

BUFx3_ASAP7_75t_L g159 ( 
.A(n_138),
.Y(n_159)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_159),
.Y(n_208)
);

AO21x2_ASAP7_75t_L g160 ( 
.A1(n_136),
.A2(n_115),
.B(n_101),
.Y(n_160)
);

OAI22xp5_ASAP7_75t_L g222 ( 
.A1(n_160),
.A2(n_1),
.B1(n_3),
.B2(n_4),
.Y(n_222)
);

MAJIxp5_ASAP7_75t_L g161 ( 
.A(n_133),
.B(n_93),
.C(n_113),
.Y(n_161)
);

MAJIxp5_ASAP7_75t_L g194 ( 
.A(n_161),
.B(n_162),
.C(n_167),
.Y(n_194)
);

MAJIxp5_ASAP7_75t_L g162 ( 
.A(n_133),
.B(n_93),
.C(n_113),
.Y(n_162)
);

OAI22xp5_ASAP7_75t_SL g163 ( 
.A1(n_125),
.A2(n_106),
.B1(n_95),
.B2(n_90),
.Y(n_163)
);

AOI22xp5_ASAP7_75t_L g198 ( 
.A1(n_163),
.A2(n_166),
.B1(n_186),
.B2(n_193),
.Y(n_198)
);

AND2x2_ASAP7_75t_L g227 ( 
.A(n_164),
.B(n_174),
.Y(n_227)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_126),
.Y(n_165)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_165),
.Y(n_217)
);

OAI22xp5_ASAP7_75t_SL g166 ( 
.A1(n_125),
.A2(n_90),
.B1(n_102),
.B2(n_120),
.Y(n_166)
);

XOR2xp5_ASAP7_75t_L g167 ( 
.A(n_144),
.B(n_124),
.Y(n_167)
);

OAI21xp5_ASAP7_75t_SL g210 ( 
.A1(n_170),
.A2(n_182),
.B(n_148),
.Y(n_210)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_126),
.Y(n_171)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_171),
.Y(n_223)
);

CKINVDCx20_ASAP7_75t_R g172 ( 
.A(n_152),
.Y(n_172)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_135),
.Y(n_173)
);

INVxp67_ASAP7_75t_L g196 ( 
.A(n_173),
.Y(n_196)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_135),
.Y(n_174)
);

NOR2x1_ASAP7_75t_L g175 ( 
.A(n_149),
.B(n_140),
.Y(n_175)
);

INVxp67_ASAP7_75t_L g214 ( 
.A(n_175),
.Y(n_214)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_141),
.Y(n_176)
);

INVxp67_ASAP7_75t_L g221 ( 
.A(n_176),
.Y(n_221)
);

INVx13_ASAP7_75t_L g177 ( 
.A(n_131),
.Y(n_177)
);

CKINVDCx14_ASAP7_75t_R g197 ( 
.A(n_177),
.Y(n_197)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_141),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_L g199 ( 
.A(n_178),
.B(n_189),
.Y(n_199)
);

AOI22xp33_ASAP7_75t_SL g216 ( 
.A1(n_180),
.A2(n_138),
.B1(n_34),
.B2(n_4),
.Y(n_216)
);

AND2x2_ASAP7_75t_L g182 ( 
.A(n_140),
.B(n_99),
.Y(n_182)
);

AOI21xp5_ASAP7_75t_SL g200 ( 
.A1(n_183),
.A2(n_151),
.B(n_139),
.Y(n_200)
);

XOR2xp5_ASAP7_75t_L g184 ( 
.A(n_151),
.B(n_94),
.Y(n_184)
);

MAJIxp5_ASAP7_75t_L g195 ( 
.A(n_184),
.B(n_127),
.C(n_150),
.Y(n_195)
);

XNOR2x1_ASAP7_75t_L g185 ( 
.A(n_140),
.B(n_118),
.Y(n_185)
);

XNOR2xp5_ASAP7_75t_L g204 ( 
.A(n_185),
.B(n_182),
.Y(n_204)
);

OAI22xp5_ASAP7_75t_SL g186 ( 
.A1(n_137),
.A2(n_119),
.B1(n_24),
.B2(n_29),
.Y(n_186)
);

INVx11_ASAP7_75t_L g187 ( 
.A(n_142),
.Y(n_187)
);

CKINVDCx16_ASAP7_75t_R g202 ( 
.A(n_187),
.Y(n_202)
);

AOI22xp33_ASAP7_75t_L g188 ( 
.A1(n_128),
.A2(n_29),
.B1(n_118),
.B2(n_110),
.Y(n_188)
);

AOI22xp33_ASAP7_75t_L g226 ( 
.A1(n_188),
.A2(n_6),
.B1(n_7),
.B2(n_8),
.Y(n_226)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_134),
.Y(n_189)
);

OAI22xp5_ASAP7_75t_SL g205 ( 
.A1(n_190),
.A2(n_150),
.B1(n_153),
.B2(n_156),
.Y(n_205)
);

NAND2xp5_ASAP7_75t_SL g191 ( 
.A(n_132),
.B(n_1),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_L g211 ( 
.A(n_191),
.B(n_192),
.Y(n_211)
);

INVx1_ASAP7_75t_SL g192 ( 
.A(n_154),
.Y(n_192)
);

MAJIxp5_ASAP7_75t_L g245 ( 
.A(n_195),
.B(n_204),
.C(n_161),
.Y(n_245)
);

OAI21xp5_ASAP7_75t_SL g246 ( 
.A1(n_200),
.A2(n_213),
.B(n_225),
.Y(n_246)
);

AOI21xp5_ASAP7_75t_L g201 ( 
.A1(n_170),
.A2(n_143),
.B(n_137),
.Y(n_201)
);

AOI21xp5_ASAP7_75t_L g239 ( 
.A1(n_201),
.A2(n_210),
.B(n_216),
.Y(n_239)
);

OAI21xp5_ASAP7_75t_L g203 ( 
.A1(n_175),
.A2(n_142),
.B(n_147),
.Y(n_203)
);

OAI21xp5_ASAP7_75t_L g243 ( 
.A1(n_203),
.A2(n_219),
.B(n_224),
.Y(n_243)
);

AOI22xp5_ASAP7_75t_L g247 ( 
.A1(n_205),
.A2(n_207),
.B1(n_222),
.B2(n_186),
.Y(n_247)
);

AOI22xp5_ASAP7_75t_L g206 ( 
.A1(n_163),
.A2(n_129),
.B1(n_157),
.B2(n_156),
.Y(n_206)
);

OAI22xp5_ASAP7_75t_SL g255 ( 
.A1(n_206),
.A2(n_212),
.B1(n_218),
.B2(n_178),
.Y(n_255)
);

OAI22xp5_ASAP7_75t_SL g207 ( 
.A1(n_189),
.A2(n_154),
.B1(n_148),
.B2(n_130),
.Y(n_207)
);

AOI22xp5_ASAP7_75t_L g212 ( 
.A1(n_166),
.A2(n_130),
.B1(n_145),
.B2(n_131),
.Y(n_212)
);

OA21x2_ASAP7_75t_L g213 ( 
.A1(n_181),
.A2(n_145),
.B(n_131),
.Y(n_213)
);

NAND2xp5_ASAP7_75t_L g215 ( 
.A(n_179),
.B(n_138),
.Y(n_215)
);

NAND2xp5_ASAP7_75t_L g234 ( 
.A(n_215),
.B(n_228),
.Y(n_234)
);

AOI22xp5_ASAP7_75t_L g218 ( 
.A1(n_184),
.A2(n_34),
.B1(n_3),
.B2(n_4),
.Y(n_218)
);

OAI21xp5_ASAP7_75t_L g219 ( 
.A1(n_168),
.A2(n_183),
.B(n_179),
.Y(n_219)
);

CKINVDCx20_ASAP7_75t_R g220 ( 
.A(n_187),
.Y(n_220)
);

NOR2xp33_ASAP7_75t_L g237 ( 
.A(n_220),
.B(n_192),
.Y(n_237)
);

OAI21xp5_ASAP7_75t_L g224 ( 
.A1(n_169),
.A2(n_5),
.B(n_6),
.Y(n_224)
);

AOI21xp5_ASAP7_75t_L g225 ( 
.A1(n_160),
.A2(n_5),
.B(n_6),
.Y(n_225)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_226),
.Y(n_232)
);

NAND2xp5_ASAP7_75t_L g228 ( 
.A(n_160),
.B(n_6),
.Y(n_228)
);

OAI21xp33_ASAP7_75t_L g229 ( 
.A1(n_211),
.A2(n_182),
.B(n_185),
.Y(n_229)
);

OAI21xp5_ASAP7_75t_SL g275 ( 
.A1(n_229),
.A2(n_259),
.B(n_202),
.Y(n_275)
);

CKINVDCx14_ASAP7_75t_R g230 ( 
.A(n_227),
.Y(n_230)
);

NAND2xp5_ASAP7_75t_L g281 ( 
.A(n_230),
.B(n_237),
.Y(n_281)
);

NOR2xp33_ASAP7_75t_SL g231 ( 
.A(n_209),
.B(n_162),
.Y(n_231)
);

NAND2xp5_ASAP7_75t_SL g265 ( 
.A(n_231),
.B(n_244),
.Y(n_265)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_215),
.Y(n_233)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_233),
.Y(n_262)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_223),
.Y(n_235)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_235),
.Y(n_276)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_223),
.Y(n_236)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_236),
.Y(n_285)
);

OAI22xp5_ASAP7_75t_L g238 ( 
.A1(n_198),
.A2(n_181),
.B1(n_160),
.B2(n_190),
.Y(n_238)
);

AOI22xp5_ASAP7_75t_L g264 ( 
.A1(n_238),
.A2(n_255),
.B1(n_213),
.B2(n_203),
.Y(n_264)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_217),
.Y(n_240)
);

INVxp67_ASAP7_75t_L g273 ( 
.A(n_240),
.Y(n_273)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_217),
.Y(n_241)
);

HB1xp67_ASAP7_75t_L g261 ( 
.A(n_241),
.Y(n_261)
);

CKINVDCx20_ASAP7_75t_R g242 ( 
.A(n_199),
.Y(n_242)
);

NOR2xp33_ASAP7_75t_L g267 ( 
.A(n_242),
.B(n_248),
.Y(n_267)
);

NAND2xp5_ASAP7_75t_SL g244 ( 
.A(n_211),
.B(n_167),
.Y(n_244)
);

MAJIxp5_ASAP7_75t_L g260 ( 
.A(n_245),
.B(n_251),
.C(n_194),
.Y(n_260)
);

OAI22xp5_ASAP7_75t_L g283 ( 
.A1(n_247),
.A2(n_256),
.B1(n_257),
.B2(n_258),
.Y(n_283)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_199),
.Y(n_248)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_196),
.Y(n_249)
);

NOR2xp33_ASAP7_75t_L g274 ( 
.A(n_249),
.B(n_250),
.Y(n_274)
);

CKINVDCx20_ASAP7_75t_R g250 ( 
.A(n_207),
.Y(n_250)
);

MAJIxp5_ASAP7_75t_L g251 ( 
.A(n_194),
.B(n_171),
.C(n_174),
.Y(n_251)
);

NAND2xp5_ASAP7_75t_L g252 ( 
.A(n_227),
.B(n_160),
.Y(n_252)
);

CKINVDCx20_ASAP7_75t_R g269 ( 
.A(n_252),
.Y(n_269)
);

OAI21xp5_ASAP7_75t_L g253 ( 
.A1(n_214),
.A2(n_201),
.B(n_200),
.Y(n_253)
);

OAI21xp5_ASAP7_75t_L g272 ( 
.A1(n_253),
.A2(n_225),
.B(n_224),
.Y(n_272)
);

CKINVDCx20_ASAP7_75t_R g254 ( 
.A(n_227),
.Y(n_254)
);

CKINVDCx20_ASAP7_75t_R g278 ( 
.A(n_254),
.Y(n_278)
);

NOR2xp33_ASAP7_75t_L g256 ( 
.A(n_220),
.B(n_176),
.Y(n_256)
);

NAND2xp5_ASAP7_75t_L g257 ( 
.A(n_228),
.B(n_164),
.Y(n_257)
);

NOR2xp33_ASAP7_75t_L g258 ( 
.A(n_196),
.B(n_164),
.Y(n_258)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_221),
.Y(n_259)
);

MAJIxp5_ASAP7_75t_L g295 ( 
.A(n_260),
.B(n_263),
.C(n_266),
.Y(n_295)
);

MAJIxp5_ASAP7_75t_L g263 ( 
.A(n_251),
.B(n_195),
.C(n_204),
.Y(n_263)
);

OAI22xp5_ASAP7_75t_SL g304 ( 
.A1(n_264),
.A2(n_280),
.B1(n_274),
.B2(n_262),
.Y(n_304)
);

MAJIxp5_ASAP7_75t_L g266 ( 
.A(n_245),
.B(n_214),
.C(n_219),
.Y(n_266)
);

MAJIxp5_ASAP7_75t_L g268 ( 
.A(n_244),
.B(n_210),
.C(n_212),
.Y(n_268)
);

MAJIxp5_ASAP7_75t_L g306 ( 
.A(n_268),
.B(n_271),
.C(n_286),
.Y(n_306)
);

XNOR2xp5_ASAP7_75t_SL g270 ( 
.A(n_248),
.B(n_198),
.Y(n_270)
);

XOR2xp5_ASAP7_75t_L g289 ( 
.A(n_270),
.B(n_275),
.Y(n_289)
);

MAJIxp5_ASAP7_75t_L g271 ( 
.A(n_253),
.B(n_242),
.C(n_254),
.Y(n_271)
);

NOR3xp33_ASAP7_75t_L g303 ( 
.A(n_272),
.B(n_257),
.C(n_234),
.Y(n_303)
);

XNOR2xp5_ASAP7_75t_L g277 ( 
.A(n_243),
.B(n_218),
.Y(n_277)
);

XOR2xp5_ASAP7_75t_L g291 ( 
.A(n_277),
.B(n_284),
.Y(n_291)
);

MAJx2_ASAP7_75t_L g279 ( 
.A(n_231),
.B(n_205),
.C(n_222),
.Y(n_279)
);

XNOR2xp5_ASAP7_75t_L g294 ( 
.A(n_279),
.B(n_246),
.Y(n_294)
);

AOI22xp5_ASAP7_75t_L g280 ( 
.A1(n_238),
.A2(n_213),
.B1(n_206),
.B2(n_221),
.Y(n_280)
);

OAI22xp5_ASAP7_75t_SL g282 ( 
.A1(n_250),
.A2(n_164),
.B1(n_208),
.B2(n_159),
.Y(n_282)
);

AOI22xp5_ASAP7_75t_L g296 ( 
.A1(n_282),
.A2(n_255),
.B1(n_230),
.B2(n_259),
.Y(n_296)
);

XNOR2xp5_ASAP7_75t_L g284 ( 
.A(n_243),
.B(n_208),
.Y(n_284)
);

MAJIxp5_ASAP7_75t_L g286 ( 
.A(n_252),
.B(n_177),
.C(n_197),
.Y(n_286)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_261),
.Y(n_287)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_287),
.Y(n_312)
);

NOR2xp33_ASAP7_75t_SL g288 ( 
.A(n_265),
.B(n_249),
.Y(n_288)
);

NOR2xp33_ASAP7_75t_SL g317 ( 
.A(n_288),
.B(n_298),
.Y(n_317)
);

OAI22xp5_ASAP7_75t_L g290 ( 
.A1(n_280),
.A2(n_247),
.B1(n_258),
.B2(n_232),
.Y(n_290)
);

HB1xp67_ASAP7_75t_L g322 ( 
.A(n_290),
.Y(n_322)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_267),
.Y(n_292)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_292),
.Y(n_313)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_276),
.Y(n_293)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_293),
.Y(n_315)
);

XNOR2xp5_ASAP7_75t_L g311 ( 
.A(n_294),
.B(n_297),
.Y(n_311)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_296),
.Y(n_323)
);

XNOR2xp5_ASAP7_75t_L g297 ( 
.A(n_260),
.B(n_266),
.Y(n_297)
);

NAND2xp5_ASAP7_75t_SL g298 ( 
.A(n_271),
.B(n_237),
.Y(n_298)
);

OAI21xp5_ASAP7_75t_SL g299 ( 
.A1(n_278),
.A2(n_239),
.B(n_246),
.Y(n_299)
);

AOI21xp5_ASAP7_75t_SL g316 ( 
.A1(n_299),
.A2(n_303),
.B(n_272),
.Y(n_316)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_285),
.Y(n_300)
);

AOI22xp33_ASAP7_75t_L g321 ( 
.A1(n_300),
.A2(n_307),
.B1(n_273),
.B2(n_235),
.Y(n_321)
);

XOR2xp5_ASAP7_75t_L g301 ( 
.A(n_263),
.B(n_233),
.Y(n_301)
);

XOR2xp5_ASAP7_75t_L g319 ( 
.A(n_301),
.B(n_302),
.Y(n_319)
);

XOR2xp5_ASAP7_75t_L g302 ( 
.A(n_268),
.B(n_234),
.Y(n_302)
);

AOI22xp5_ASAP7_75t_L g310 ( 
.A1(n_304),
.A2(n_282),
.B1(n_281),
.B2(n_269),
.Y(n_310)
);

AOI22xp5_ASAP7_75t_L g305 ( 
.A1(n_283),
.A2(n_232),
.B1(n_239),
.B2(n_236),
.Y(n_305)
);

NAND2xp5_ASAP7_75t_L g325 ( 
.A(n_305),
.B(n_264),
.Y(n_325)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_273),
.Y(n_307)
);

NOR2xp33_ASAP7_75t_L g308 ( 
.A(n_270),
.B(n_241),
.Y(n_308)
);

NOR2xp33_ASAP7_75t_SL g320 ( 
.A(n_308),
.B(n_309),
.Y(n_320)
);

NOR2xp33_ASAP7_75t_L g309 ( 
.A(n_277),
.B(n_240),
.Y(n_309)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_310),
.Y(n_330)
);

NOR2xp33_ASAP7_75t_L g314 ( 
.A(n_301),
.B(n_302),
.Y(n_314)
);

NAND2xp5_ASAP7_75t_L g328 ( 
.A(n_314),
.B(n_318),
.Y(n_328)
);

XOR2xp5_ASAP7_75t_L g334 ( 
.A(n_316),
.B(n_294),
.Y(n_334)
);

NOR2xp33_ASAP7_75t_L g318 ( 
.A(n_297),
.B(n_284),
.Y(n_318)
);

NAND2xp5_ASAP7_75t_L g337 ( 
.A(n_321),
.B(n_324),
.Y(n_337)
);

BUFx12_ASAP7_75t_L g324 ( 
.A(n_299),
.Y(n_324)
);

NAND2xp5_ASAP7_75t_L g339 ( 
.A(n_325),
.B(n_327),
.Y(n_339)
);

OAI21xp5_ASAP7_75t_SL g326 ( 
.A1(n_305),
.A2(n_286),
.B(n_279),
.Y(n_326)
);

AOI21xp5_ASAP7_75t_L g335 ( 
.A1(n_326),
.A2(n_289),
.B(n_291),
.Y(n_335)
);

INVxp67_ASAP7_75t_SL g327 ( 
.A(n_307),
.Y(n_327)
);

NOR2xp33_ASAP7_75t_L g329 ( 
.A(n_317),
.B(n_304),
.Y(n_329)
);

NAND2xp5_ASAP7_75t_SL g344 ( 
.A(n_329),
.B(n_331),
.Y(n_344)
);

NOR2xp33_ASAP7_75t_L g331 ( 
.A(n_320),
.B(n_306),
.Y(n_331)
);

MAJIxp5_ASAP7_75t_L g332 ( 
.A(n_319),
.B(n_295),
.C(n_306),
.Y(n_332)
);

MAJIxp5_ASAP7_75t_L g353 ( 
.A(n_332),
.B(n_336),
.C(n_342),
.Y(n_353)
);

NOR2xp33_ASAP7_75t_L g333 ( 
.A(n_313),
.B(n_295),
.Y(n_333)
);

INVx1_ASAP7_75t_L g343 ( 
.A(n_333),
.Y(n_343)
);

AND2x2_ASAP7_75t_L g352 ( 
.A(n_334),
.B(n_340),
.Y(n_352)
);

OAI22xp5_ASAP7_75t_SL g345 ( 
.A1(n_335),
.A2(n_341),
.B1(n_316),
.B2(n_310),
.Y(n_345)
);

MAJIxp5_ASAP7_75t_L g336 ( 
.A(n_319),
.B(n_291),
.C(n_289),
.Y(n_336)
);

NOR2xp33_ASAP7_75t_L g338 ( 
.A(n_313),
.B(n_296),
.Y(n_338)
);

CKINVDCx20_ASAP7_75t_R g350 ( 
.A(n_338),
.Y(n_350)
);

AOI21xp5_ASAP7_75t_L g340 ( 
.A1(n_326),
.A2(n_256),
.B(n_9),
.Y(n_340)
);

AOI22xp5_ASAP7_75t_L g341 ( 
.A1(n_322),
.A2(n_12),
.B1(n_9),
.B2(n_10),
.Y(n_341)
);

MAJIxp5_ASAP7_75t_L g342 ( 
.A(n_311),
.B(n_7),
.C(n_10),
.Y(n_342)
);

AOI22xp5_ASAP7_75t_L g361 ( 
.A1(n_345),
.A2(n_11),
.B1(n_12),
.B2(n_352),
.Y(n_361)
);

AOI22xp33_ASAP7_75t_L g346 ( 
.A1(n_330),
.A2(n_315),
.B1(n_312),
.B2(n_323),
.Y(n_346)
);

NAND2xp5_ASAP7_75t_L g359 ( 
.A(n_346),
.B(n_347),
.Y(n_359)
);

AOI22xp33_ASAP7_75t_L g347 ( 
.A1(n_339),
.A2(n_315),
.B1(n_323),
.B2(n_324),
.Y(n_347)
);

AOI22xp5_ASAP7_75t_L g348 ( 
.A1(n_337),
.A2(n_325),
.B1(n_334),
.B2(n_324),
.Y(n_348)
);

NAND2xp5_ASAP7_75t_L g362 ( 
.A(n_348),
.B(n_349),
.Y(n_362)
);

NOR2xp33_ASAP7_75t_L g349 ( 
.A(n_328),
.B(n_311),
.Y(n_349)
);

NOR2xp33_ASAP7_75t_L g351 ( 
.A(n_332),
.B(n_7),
.Y(n_351)
);

NOR2xp33_ASAP7_75t_SL g363 ( 
.A(n_351),
.B(n_12),
.Y(n_363)
);

MAJIxp5_ASAP7_75t_L g354 ( 
.A(n_336),
.B(n_7),
.C(n_11),
.Y(n_354)
);

NAND2xp5_ASAP7_75t_SL g358 ( 
.A(n_354),
.B(n_11),
.Y(n_358)
);

NOR2xp33_ASAP7_75t_L g355 ( 
.A(n_350),
.B(n_341),
.Y(n_355)
);

NAND2xp5_ASAP7_75t_L g364 ( 
.A(n_355),
.B(n_357),
.Y(n_364)
);

XOR2xp5_ASAP7_75t_L g356 ( 
.A(n_345),
.B(n_335),
.Y(n_356)
);

XNOR2xp5_ASAP7_75t_L g366 ( 
.A(n_356),
.B(n_348),
.Y(n_366)
);

OAI21xp5_ASAP7_75t_L g357 ( 
.A1(n_352),
.A2(n_340),
.B(n_342),
.Y(n_357)
);

INVx1_ASAP7_75t_L g365 ( 
.A(n_358),
.Y(n_365)
);

NAND2xp5_ASAP7_75t_SL g360 ( 
.A(n_343),
.B(n_11),
.Y(n_360)
);

NOR2xp33_ASAP7_75t_L g368 ( 
.A(n_360),
.B(n_363),
.Y(n_368)
);

XOR2xp5_ASAP7_75t_L g367 ( 
.A(n_361),
.B(n_352),
.Y(n_367)
);

INVx1_ASAP7_75t_L g370 ( 
.A(n_366),
.Y(n_370)
);

INVx1_ASAP7_75t_L g372 ( 
.A(n_367),
.Y(n_372)
);

NOR2xp67_ASAP7_75t_SL g369 ( 
.A(n_356),
.B(n_353),
.Y(n_369)
);

INVxp67_ASAP7_75t_L g373 ( 
.A(n_369),
.Y(n_373)
);

XOR2xp5_ASAP7_75t_L g371 ( 
.A(n_364),
.B(n_353),
.Y(n_371)
);

OAI21xp5_ASAP7_75t_SL g374 ( 
.A1(n_371),
.A2(n_344),
.B(n_362),
.Y(n_374)
);

OAI22xp5_ASAP7_75t_L g376 ( 
.A1(n_374),
.A2(n_375),
.B1(n_370),
.B2(n_372),
.Y(n_376)
);

OAI21xp5_ASAP7_75t_L g375 ( 
.A1(n_373),
.A2(n_359),
.B(n_357),
.Y(n_375)
);

MAJIxp5_ASAP7_75t_L g377 ( 
.A(n_376),
.B(n_365),
.C(n_354),
.Y(n_377)
);

OAI21x1_ASAP7_75t_L g378 ( 
.A1(n_377),
.A2(n_368),
.B(n_369),
.Y(n_378)
);

BUFx24_ASAP7_75t_SL g379 ( 
.A(n_378),
.Y(n_379)
);


endmodule