module fake_jpeg_684_n_528 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_528);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_528;

wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_525;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_16;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_519;
wire n_276;
wire n_143;
wire n_17;
wire n_431;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_513;
wire n_283;
wire n_107;
wire n_490;
wire n_517;
wire n_415;
wire n_479;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_48;
wire n_465;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_256;
wire n_221;
wire n_454;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_508;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_474;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_511;
wire n_305;
wire n_161;
wire n_441;
wire n_342;
wire n_101;
wire n_226;
wire n_509;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_510;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_523;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_296;
wire n_384;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_491;
wire n_24;
wire n_526;
wire n_467;
wire n_269;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_473;
wire n_45;
wire n_520;
wire n_476;
wire n_337;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_481;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_522;
wire n_333;
wire n_518;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_199;
wire n_260;
wire n_413;
wire n_275;
wire n_494;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_492;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_515;
wire n_347;
wire n_521;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_472;
wire n_279;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_484;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_469;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_527;
wire n_482;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_512;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_516;
wire n_183;
wire n_409;
wire n_249;
wire n_412;
wire n_217;
wire n_471;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_524;
wire n_402;
wire n_504;
wire n_438;
wire n_475;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_514;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

BUFx12f_ASAP7_75t_L g16 ( 
.A(n_4),
.Y(n_16)
);

INVx2_ASAP7_75t_L g17 ( 
.A(n_10),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_2),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_3),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_1),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_8),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_11),
.Y(n_22)
);

INVx6_ASAP7_75t_L g23 ( 
.A(n_14),
.Y(n_23)
);

BUFx3_ASAP7_75t_L g24 ( 
.A(n_11),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_0),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_12),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_11),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_1),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_4),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_9),
.Y(n_30)
);

BUFx24_ASAP7_75t_L g31 ( 
.A(n_5),
.Y(n_31)
);

INVx11_ASAP7_75t_L g32 ( 
.A(n_1),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_3),
.Y(n_33)
);

INVx3_ASAP7_75t_L g34 ( 
.A(n_1),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_10),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_14),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_14),
.Y(n_37)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_6),
.Y(n_38)
);

INVx8_ASAP7_75t_L g39 ( 
.A(n_4),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_0),
.Y(n_40)
);

INVx13_ASAP7_75t_L g41 ( 
.A(n_2),
.Y(n_41)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_8),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_13),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_12),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_37),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g136 ( 
.A(n_45),
.Y(n_136)
);

INVx4_ASAP7_75t_L g46 ( 
.A(n_34),
.Y(n_46)
);

INVx3_ASAP7_75t_L g101 ( 
.A(n_46),
.Y(n_101)
);

INVx2_ASAP7_75t_L g47 ( 
.A(n_17),
.Y(n_47)
);

INVx2_ASAP7_75t_L g97 ( 
.A(n_47),
.Y(n_97)
);

BUFx3_ASAP7_75t_L g48 ( 
.A(n_24),
.Y(n_48)
);

BUFx3_ASAP7_75t_L g113 ( 
.A(n_48),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_L g49 ( 
.A(n_17),
.B(n_34),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_L g115 ( 
.A(n_49),
.B(n_55),
.Y(n_115)
);

INVx5_ASAP7_75t_L g50 ( 
.A(n_39),
.Y(n_50)
);

BUFx3_ASAP7_75t_L g137 ( 
.A(n_50),
.Y(n_137)
);

BUFx5_ASAP7_75t_L g51 ( 
.A(n_17),
.Y(n_51)
);

INVx2_ASAP7_75t_SL g125 ( 
.A(n_51),
.Y(n_125)
);

INVx4_ASAP7_75t_L g52 ( 
.A(n_34),
.Y(n_52)
);

INVx3_ASAP7_75t_L g124 ( 
.A(n_52),
.Y(n_124)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_34),
.Y(n_53)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_53),
.Y(n_103)
);

INVx11_ASAP7_75t_L g54 ( 
.A(n_16),
.Y(n_54)
);

INVx4_ASAP7_75t_L g107 ( 
.A(n_54),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_36),
.B(n_15),
.Y(n_55)
);

INVx6_ASAP7_75t_L g56 ( 
.A(n_37),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g141 ( 
.A(n_56),
.Y(n_141)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_37),
.Y(n_57)
);

INVx3_ASAP7_75t_SL g118 ( 
.A(n_57),
.Y(n_118)
);

INVx6_ASAP7_75t_L g58 ( 
.A(n_37),
.Y(n_58)
);

BUFx2_ASAP7_75t_L g145 ( 
.A(n_58),
.Y(n_145)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_37),
.Y(n_59)
);

INVx8_ASAP7_75t_L g120 ( 
.A(n_59),
.Y(n_120)
);

INVx8_ASAP7_75t_L g60 ( 
.A(n_16),
.Y(n_60)
);

INVx3_ASAP7_75t_L g105 ( 
.A(n_60),
.Y(n_105)
);

BUFx24_ASAP7_75t_L g61 ( 
.A(n_31),
.Y(n_61)
);

INVx8_ASAP7_75t_L g121 ( 
.A(n_61),
.Y(n_121)
);

BUFx5_ASAP7_75t_L g62 ( 
.A(n_31),
.Y(n_62)
);

INVx4_ASAP7_75t_L g129 ( 
.A(n_62),
.Y(n_129)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_43),
.Y(n_63)
);

INVx3_ASAP7_75t_L g111 ( 
.A(n_63),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_36),
.B(n_15),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_L g122 ( 
.A(n_64),
.B(n_65),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_L g65 ( 
.A(n_36),
.B(n_15),
.Y(n_65)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_43),
.Y(n_66)
);

INVx3_ASAP7_75t_L g123 ( 
.A(n_66),
.Y(n_123)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_43),
.Y(n_67)
);

INVx3_ASAP7_75t_L g126 ( 
.A(n_67),
.Y(n_126)
);

INVx3_ASAP7_75t_L g68 ( 
.A(n_24),
.Y(n_68)
);

HB1xp67_ASAP7_75t_L g128 ( 
.A(n_68),
.Y(n_128)
);

INVx2_ASAP7_75t_L g69 ( 
.A(n_16),
.Y(n_69)
);

INVx2_ASAP7_75t_L g98 ( 
.A(n_69),
.Y(n_98)
);

BUFx5_ASAP7_75t_L g70 ( 
.A(n_31),
.Y(n_70)
);

INVx4_ASAP7_75t_L g139 ( 
.A(n_70),
.Y(n_139)
);

INVx4_ASAP7_75t_SL g71 ( 
.A(n_16),
.Y(n_71)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_71),
.Y(n_116)
);

INVx6_ASAP7_75t_L g72 ( 
.A(n_43),
.Y(n_72)
);

INVx2_ASAP7_75t_L g99 ( 
.A(n_72),
.Y(n_99)
);

INVx3_ASAP7_75t_L g73 ( 
.A(n_24),
.Y(n_73)
);

INVx3_ASAP7_75t_L g135 ( 
.A(n_73),
.Y(n_135)
);

INVx5_ASAP7_75t_L g74 ( 
.A(n_39),
.Y(n_74)
);

INVx4_ASAP7_75t_L g140 ( 
.A(n_74),
.Y(n_140)
);

INVx4_ASAP7_75t_L g75 ( 
.A(n_24),
.Y(n_75)
);

INVx3_ASAP7_75t_L g148 ( 
.A(n_75),
.Y(n_148)
);

BUFx6f_ASAP7_75t_L g76 ( 
.A(n_43),
.Y(n_76)
);

INVx3_ASAP7_75t_L g149 ( 
.A(n_76),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_L g77 ( 
.A(n_18),
.B(n_15),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_L g130 ( 
.A(n_77),
.B(n_94),
.Y(n_130)
);

BUFx12f_ASAP7_75t_L g78 ( 
.A(n_39),
.Y(n_78)
);

INVx4_ASAP7_75t_L g152 ( 
.A(n_78),
.Y(n_152)
);

BUFx6f_ASAP7_75t_L g79 ( 
.A(n_44),
.Y(n_79)
);

INVx2_ASAP7_75t_L g106 ( 
.A(n_79),
.Y(n_106)
);

BUFx5_ASAP7_75t_L g80 ( 
.A(n_31),
.Y(n_80)
);

INVx2_ASAP7_75t_L g109 ( 
.A(n_80),
.Y(n_109)
);

BUFx6f_ASAP7_75t_L g81 ( 
.A(n_44),
.Y(n_81)
);

INVx2_ASAP7_75t_L g110 ( 
.A(n_81),
.Y(n_110)
);

INVx4_ASAP7_75t_SL g82 ( 
.A(n_16),
.Y(n_82)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_82),
.Y(n_117)
);

BUFx3_ASAP7_75t_L g83 ( 
.A(n_39),
.Y(n_83)
);

INVx2_ASAP7_75t_L g112 ( 
.A(n_83),
.Y(n_112)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_23),
.Y(n_84)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_84),
.Y(n_138)
);

INVx2_ASAP7_75t_L g85 ( 
.A(n_16),
.Y(n_85)
);

INVx2_ASAP7_75t_L g153 ( 
.A(n_85),
.Y(n_153)
);

BUFx12f_ASAP7_75t_L g86 ( 
.A(n_44),
.Y(n_86)
);

AND2x2_ASAP7_75t_L g104 ( 
.A(n_86),
.B(n_91),
.Y(n_104)
);

BUFx5_ASAP7_75t_L g87 ( 
.A(n_31),
.Y(n_87)
);

INVx2_ASAP7_75t_L g155 ( 
.A(n_87),
.Y(n_155)
);

INVx2_ASAP7_75t_L g88 ( 
.A(n_16),
.Y(n_88)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_88),
.Y(n_143)
);

INVx2_ASAP7_75t_L g89 ( 
.A(n_22),
.Y(n_89)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_89),
.Y(n_146)
);

INVx4_ASAP7_75t_SL g90 ( 
.A(n_44),
.Y(n_90)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_90),
.Y(n_156)
);

INVx8_ASAP7_75t_L g91 ( 
.A(n_22),
.Y(n_91)
);

BUFx6f_ASAP7_75t_L g92 ( 
.A(n_44),
.Y(n_92)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_92),
.Y(n_150)
);

BUFx2_ASAP7_75t_L g93 ( 
.A(n_22),
.Y(n_93)
);

AND2x2_ASAP7_75t_L g133 ( 
.A(n_93),
.B(n_96),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_23),
.B(n_14),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_23),
.B(n_13),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g147 ( 
.A(n_95),
.B(n_18),
.Y(n_147)
);

INVx2_ASAP7_75t_L g96 ( 
.A(n_22),
.Y(n_96)
);

AOI22xp33_ASAP7_75t_SL g100 ( 
.A1(n_71),
.A2(n_32),
.B1(n_20),
.B2(n_40),
.Y(n_100)
);

OA22x2_ASAP7_75t_L g158 ( 
.A1(n_100),
.A2(n_108),
.B1(n_132),
.B2(n_144),
.Y(n_158)
);

AOI22xp5_ASAP7_75t_L g102 ( 
.A1(n_45),
.A2(n_79),
.B1(n_92),
.B2(n_57),
.Y(n_102)
);

OAI22xp5_ASAP7_75t_L g160 ( 
.A1(n_102),
.A2(n_114),
.B1(n_30),
.B2(n_29),
.Y(n_160)
);

AOI22xp33_ASAP7_75t_SL g108 ( 
.A1(n_82),
.A2(n_32),
.B1(n_20),
.B2(n_40),
.Y(n_108)
);

AOI22xp33_ASAP7_75t_L g114 ( 
.A1(n_59),
.A2(n_40),
.B1(n_22),
.B2(n_20),
.Y(n_114)
);

OAI21xp33_ASAP7_75t_L g119 ( 
.A1(n_73),
.A2(n_19),
.B(n_18),
.Y(n_119)
);

OAI21xp33_ASAP7_75t_L g168 ( 
.A1(n_119),
.A2(n_61),
.B(n_31),
.Y(n_168)
);

CKINVDCx20_ASAP7_75t_R g127 ( 
.A(n_93),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_L g181 ( 
.A(n_127),
.B(n_142),
.Y(n_181)
);

NOR2xp33_ASAP7_75t_L g131 ( 
.A(n_46),
.B(n_23),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g173 ( 
.A(n_131),
.B(n_134),
.Y(n_173)
);

AOI22xp33_ASAP7_75t_SL g132 ( 
.A1(n_90),
.A2(n_32),
.B1(n_20),
.B2(n_40),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_L g134 ( 
.A(n_52),
.B(n_26),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_L g142 ( 
.A(n_48),
.B(n_26),
.Y(n_142)
);

AOI22xp33_ASAP7_75t_SL g144 ( 
.A1(n_83),
.A2(n_32),
.B1(n_40),
.B2(n_33),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_SL g165 ( 
.A(n_147),
.B(n_151),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_L g151 ( 
.A(n_75),
.B(n_19),
.Y(n_151)
);

OAI22xp33_ASAP7_75t_SL g154 ( 
.A1(n_63),
.A2(n_19),
.B1(n_33),
.B2(n_30),
.Y(n_154)
);

AOI22xp5_ASAP7_75t_L g159 ( 
.A1(n_154),
.A2(n_29),
.B1(n_30),
.B2(n_33),
.Y(n_159)
);

NOR2x1_ASAP7_75t_R g157 ( 
.A(n_115),
.B(n_119),
.Y(n_157)
);

CKINVDCx14_ASAP7_75t_R g216 ( 
.A(n_157),
.Y(n_216)
);

AOI22xp5_ASAP7_75t_L g205 ( 
.A1(n_159),
.A2(n_188),
.B1(n_196),
.B2(n_25),
.Y(n_205)
);

AOI22xp33_ASAP7_75t_SL g207 ( 
.A1(n_160),
.A2(n_194),
.B1(n_195),
.B2(n_198),
.Y(n_207)
);

INVx2_ASAP7_75t_L g161 ( 
.A(n_99),
.Y(n_161)
);

BUFx2_ASAP7_75t_L g209 ( 
.A(n_161),
.Y(n_209)
);

AOI22xp33_ASAP7_75t_L g162 ( 
.A1(n_154),
.A2(n_29),
.B1(n_81),
.B2(n_76),
.Y(n_162)
);

OAI22xp5_ASAP7_75t_L g203 ( 
.A1(n_162),
.A2(n_132),
.B1(n_118),
.B2(n_27),
.Y(n_203)
);

INVx2_ASAP7_75t_L g163 ( 
.A(n_106),
.Y(n_163)
);

INVx2_ASAP7_75t_L g210 ( 
.A(n_163),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_L g164 ( 
.A(n_130),
.B(n_28),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_SL g235 ( 
.A(n_164),
.B(n_201),
.Y(n_235)
);

MAJIxp5_ASAP7_75t_L g166 ( 
.A(n_103),
.B(n_67),
.C(n_66),
.Y(n_166)
);

AND2x2_ASAP7_75t_L g211 ( 
.A(n_166),
.B(n_175),
.Y(n_211)
);

INVx4_ASAP7_75t_L g167 ( 
.A(n_105),
.Y(n_167)
);

INVx4_ASAP7_75t_L g220 ( 
.A(n_167),
.Y(n_220)
);

CKINVDCx16_ASAP7_75t_R g223 ( 
.A(n_168),
.Y(n_223)
);

OAI22xp33_ASAP7_75t_SL g169 ( 
.A1(n_114),
.A2(n_54),
.B1(n_26),
.B2(n_61),
.Y(n_169)
);

AOI22xp5_ASAP7_75t_SL g233 ( 
.A1(n_169),
.A2(n_199),
.B1(n_202),
.B2(n_139),
.Y(n_233)
);

INVx2_ASAP7_75t_L g170 ( 
.A(n_110),
.Y(n_170)
);

INVx2_ASAP7_75t_L g225 ( 
.A(n_170),
.Y(n_225)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_138),
.Y(n_171)
);

INVx1_ASAP7_75t_SL g232 ( 
.A(n_171),
.Y(n_232)
);

INVx3_ASAP7_75t_SL g172 ( 
.A(n_121),
.Y(n_172)
);

INVx2_ASAP7_75t_L g227 ( 
.A(n_172),
.Y(n_227)
);

NAND2xp5_ASAP7_75t_SL g174 ( 
.A(n_122),
.B(n_50),
.Y(n_174)
);

NOR2xp33_ASAP7_75t_L g212 ( 
.A(n_174),
.B(n_182),
.Y(n_212)
);

AOI22xp5_ASAP7_75t_SL g175 ( 
.A1(n_112),
.A2(n_74),
.B1(n_21),
.B2(n_38),
.Y(n_175)
);

INVx4_ASAP7_75t_L g176 ( 
.A(n_105),
.Y(n_176)
);

INVx5_ASAP7_75t_L g221 ( 
.A(n_176),
.Y(n_221)
);

BUFx6f_ASAP7_75t_L g177 ( 
.A(n_136),
.Y(n_177)
);

BUFx6f_ASAP7_75t_L g224 ( 
.A(n_177),
.Y(n_224)
);

AND2x2_ASAP7_75t_L g178 ( 
.A(n_116),
.B(n_60),
.Y(n_178)
);

AND2x2_ASAP7_75t_L g215 ( 
.A(n_178),
.B(n_197),
.Y(n_215)
);

INVx3_ASAP7_75t_L g179 ( 
.A(n_156),
.Y(n_179)
);

INVx2_ASAP7_75t_L g228 ( 
.A(n_179),
.Y(n_228)
);

INVx4_ASAP7_75t_L g180 ( 
.A(n_140),
.Y(n_180)
);

INVx2_ASAP7_75t_L g234 ( 
.A(n_180),
.Y(n_234)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_117),
.Y(n_182)
);

BUFx8_ASAP7_75t_L g183 ( 
.A(n_121),
.Y(n_183)
);

CKINVDCx20_ASAP7_75t_R g208 ( 
.A(n_183),
.Y(n_208)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_146),
.Y(n_184)
);

NOR2xp33_ASAP7_75t_L g222 ( 
.A(n_184),
.B(n_187),
.Y(n_222)
);

INVx3_ASAP7_75t_L g185 ( 
.A(n_140),
.Y(n_185)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_185),
.Y(n_204)
);

NAND2x1_ASAP7_75t_SL g186 ( 
.A(n_129),
.B(n_21),
.Y(n_186)
);

NAND2x1_ASAP7_75t_L g213 ( 
.A(n_186),
.B(n_200),
.Y(n_213)
);

INVx13_ASAP7_75t_L g187 ( 
.A(n_125),
.Y(n_187)
);

OAI22xp5_ASAP7_75t_L g188 ( 
.A1(n_144),
.A2(n_72),
.B1(n_58),
.B2(n_56),
.Y(n_188)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_143),
.Y(n_189)
);

NOR2xp33_ASAP7_75t_L g231 ( 
.A(n_189),
.B(n_192),
.Y(n_231)
);

HB1xp67_ASAP7_75t_L g190 ( 
.A(n_135),
.Y(n_190)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_190),
.Y(n_219)
);

INVx4_ASAP7_75t_L g191 ( 
.A(n_152),
.Y(n_191)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_191),
.Y(n_226)
);

NOR2x1_ASAP7_75t_L g192 ( 
.A(n_97),
.B(n_78),
.Y(n_192)
);

BUFx2_ASAP7_75t_SL g193 ( 
.A(n_109),
.Y(n_193)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_193),
.Y(n_230)
);

BUFx6f_ASAP7_75t_L g194 ( 
.A(n_136),
.Y(n_194)
);

BUFx6f_ASAP7_75t_L g195 ( 
.A(n_141),
.Y(n_195)
);

OAI22xp33_ASAP7_75t_L g196 ( 
.A1(n_100),
.A2(n_91),
.B1(n_38),
.B2(n_35),
.Y(n_196)
);

INVx2_ASAP7_75t_L g197 ( 
.A(n_98),
.Y(n_197)
);

INVxp67_ASAP7_75t_SL g198 ( 
.A(n_155),
.Y(n_198)
);

INVx8_ASAP7_75t_L g199 ( 
.A(n_141),
.Y(n_199)
);

AND2x2_ASAP7_75t_L g200 ( 
.A(n_133),
.B(n_78),
.Y(n_200)
);

NOR2xp33_ASAP7_75t_L g201 ( 
.A(n_128),
.B(n_86),
.Y(n_201)
);

NAND2xp33_ASAP7_75t_L g202 ( 
.A(n_108),
.B(n_28),
.Y(n_202)
);

AOI22xp33_ASAP7_75t_L g246 ( 
.A1(n_203),
.A2(n_158),
.B1(n_107),
.B2(n_177),
.Y(n_246)
);

OA22x2_ASAP7_75t_L g256 ( 
.A1(n_205),
.A2(n_236),
.B1(n_107),
.B2(n_183),
.Y(n_256)
);

OAI22xp5_ASAP7_75t_SL g206 ( 
.A1(n_157),
.A2(n_150),
.B1(n_126),
.B2(n_149),
.Y(n_206)
);

AOI22xp5_ASAP7_75t_L g240 ( 
.A1(n_206),
.A2(n_214),
.B1(n_200),
.B2(n_178),
.Y(n_240)
);

OAI22xp5_ASAP7_75t_SL g214 ( 
.A1(n_165),
.A2(n_126),
.B1(n_149),
.B2(n_111),
.Y(n_214)
);

A2O1A1Ixp33_ASAP7_75t_L g217 ( 
.A1(n_168),
.A2(n_133),
.B(n_153),
.C(n_104),
.Y(n_217)
);

NAND2xp5_ASAP7_75t_L g254 ( 
.A(n_217),
.B(n_125),
.Y(n_254)
);

AOI22xp5_ASAP7_75t_L g218 ( 
.A1(n_159),
.A2(n_111),
.B1(n_123),
.B2(n_118),
.Y(n_218)
);

OAI22xp5_ASAP7_75t_L g247 ( 
.A1(n_218),
.A2(n_163),
.B1(n_170),
.B2(n_161),
.Y(n_247)
);

OAI22xp33_ASAP7_75t_SL g229 ( 
.A1(n_173),
.A2(n_123),
.B1(n_145),
.B2(n_137),
.Y(n_229)
);

AOI22xp5_ASAP7_75t_SL g263 ( 
.A1(n_229),
.A2(n_172),
.B1(n_152),
.B2(n_137),
.Y(n_263)
);

AND2x2_ASAP7_75t_L g243 ( 
.A(n_233),
.B(n_186),
.Y(n_243)
);

AOI22xp33_ASAP7_75t_L g236 ( 
.A1(n_196),
.A2(n_145),
.B1(n_135),
.B2(n_101),
.Y(n_236)
);

INVx2_ASAP7_75t_L g237 ( 
.A(n_227),
.Y(n_237)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_237),
.Y(n_267)
);

NOR2xp33_ASAP7_75t_SL g238 ( 
.A(n_212),
.B(n_164),
.Y(n_238)
);

NAND2xp5_ASAP7_75t_SL g277 ( 
.A(n_238),
.B(n_245),
.Y(n_277)
);

AOI22xp33_ASAP7_75t_SL g239 ( 
.A1(n_203),
.A2(n_158),
.B1(n_129),
.B2(n_139),
.Y(n_239)
);

INVxp67_ASAP7_75t_L g268 ( 
.A(n_239),
.Y(n_268)
);

AOI22xp5_ASAP7_75t_L g273 ( 
.A1(n_240),
.A2(n_244),
.B1(n_247),
.B2(n_250),
.Y(n_273)
);

OAI22xp5_ASAP7_75t_SL g241 ( 
.A1(n_205),
.A2(n_158),
.B1(n_175),
.B2(n_181),
.Y(n_241)
);

AOI22xp5_ASAP7_75t_L g287 ( 
.A1(n_241),
.A2(n_213),
.B1(n_208),
.B2(n_227),
.Y(n_287)
);

CKINVDCx14_ASAP7_75t_R g242 ( 
.A(n_231),
.Y(n_242)
);

NAND2xp5_ASAP7_75t_L g276 ( 
.A(n_242),
.B(n_257),
.Y(n_276)
);

OR2x2_ASAP7_75t_L g282 ( 
.A(n_243),
.B(n_263),
.Y(n_282)
);

OAI22xp5_ASAP7_75t_SL g244 ( 
.A1(n_216),
.A2(n_158),
.B1(n_200),
.B2(n_192),
.Y(n_244)
);

NOR2xp33_ASAP7_75t_SL g245 ( 
.A(n_212),
.B(n_179),
.Y(n_245)
);

OAI22xp5_ASAP7_75t_L g281 ( 
.A1(n_246),
.A2(n_249),
.B1(n_265),
.B2(n_218),
.Y(n_281)
);

CKINVDCx16_ASAP7_75t_R g248 ( 
.A(n_215),
.Y(n_248)
);

NOR2xp33_ASAP7_75t_L g272 ( 
.A(n_248),
.B(n_258),
.Y(n_272)
);

AOI22xp5_ASAP7_75t_L g249 ( 
.A1(n_211),
.A2(n_166),
.B1(n_178),
.B2(n_197),
.Y(n_249)
);

OAI22xp5_ASAP7_75t_SL g250 ( 
.A1(n_216),
.A2(n_195),
.B1(n_120),
.B2(n_104),
.Y(n_250)
);

AND2x2_ASAP7_75t_L g251 ( 
.A(n_217),
.B(n_167),
.Y(n_251)
);

OAI21xp33_ASAP7_75t_L g285 ( 
.A1(n_251),
.A2(n_254),
.B(n_213),
.Y(n_285)
);

INVx5_ASAP7_75t_L g252 ( 
.A(n_224),
.Y(n_252)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_252),
.Y(n_283)
);

MAJIxp5_ASAP7_75t_L g253 ( 
.A(n_223),
.B(n_148),
.C(n_185),
.Y(n_253)
);

XNOR2xp5_ASAP7_75t_L g271 ( 
.A(n_253),
.B(n_255),
.Y(n_271)
);

MAJIxp5_ASAP7_75t_L g255 ( 
.A(n_223),
.B(n_148),
.C(n_176),
.Y(n_255)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_256),
.Y(n_288)
);

NAND2xp5_ASAP7_75t_L g257 ( 
.A(n_235),
.B(n_180),
.Y(n_257)
);

CKINVDCx16_ASAP7_75t_R g258 ( 
.A(n_215),
.Y(n_258)
);

CKINVDCx20_ASAP7_75t_R g259 ( 
.A(n_209),
.Y(n_259)
);

NOR2xp33_ASAP7_75t_L g274 ( 
.A(n_259),
.B(n_262),
.Y(n_274)
);

NOR2xp33_ASAP7_75t_L g260 ( 
.A(n_232),
.B(n_191),
.Y(n_260)
);

NAND2xp5_ASAP7_75t_L g290 ( 
.A(n_260),
.B(n_261),
.Y(n_290)
);

NOR2xp33_ASAP7_75t_L g261 ( 
.A(n_232),
.B(n_124),
.Y(n_261)
);

CKINVDCx20_ASAP7_75t_R g262 ( 
.A(n_209),
.Y(n_262)
);

OAI22xp5_ASAP7_75t_L g264 ( 
.A1(n_211),
.A2(n_233),
.B1(n_207),
.B2(n_236),
.Y(n_264)
);

AOI22xp5_ASAP7_75t_L g275 ( 
.A1(n_264),
.A2(n_211),
.B1(n_217),
.B2(n_206),
.Y(n_275)
);

AOI22xp5_ASAP7_75t_L g265 ( 
.A1(n_211),
.A2(n_120),
.B1(n_199),
.B2(n_194),
.Y(n_265)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_232),
.Y(n_266)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_266),
.Y(n_291)
);

AOI21xp5_ASAP7_75t_L g269 ( 
.A1(n_254),
.A2(n_243),
.B(n_251),
.Y(n_269)
);

AOI21xp5_ASAP7_75t_L g299 ( 
.A1(n_269),
.A2(n_284),
.B(n_251),
.Y(n_299)
);

OAI22xp5_ASAP7_75t_SL g270 ( 
.A1(n_246),
.A2(n_239),
.B1(n_249),
.B2(n_241),
.Y(n_270)
);

AOI22xp5_ASAP7_75t_L g305 ( 
.A1(n_270),
.A2(n_281),
.B1(n_287),
.B2(n_289),
.Y(n_305)
);

OAI22x1_ASAP7_75t_L g319 ( 
.A1(n_275),
.A2(n_265),
.B1(n_240),
.B2(n_263),
.Y(n_319)
);

CKINVDCx20_ASAP7_75t_R g278 ( 
.A(n_260),
.Y(n_278)
);

NAND2xp5_ASAP7_75t_L g303 ( 
.A(n_278),
.B(n_279),
.Y(n_303)
);

CKINVDCx20_ASAP7_75t_R g279 ( 
.A(n_245),
.Y(n_279)
);

OAI32xp33_ASAP7_75t_L g280 ( 
.A1(n_257),
.A2(n_231),
.A3(n_215),
.B1(n_235),
.B2(n_222),
.Y(n_280)
);

INVxp67_ASAP7_75t_L g298 ( 
.A(n_280),
.Y(n_298)
);

AOI21xp5_ASAP7_75t_L g284 ( 
.A1(n_243),
.A2(n_213),
.B(n_208),
.Y(n_284)
);

OAI21xp5_ASAP7_75t_L g320 ( 
.A1(n_285),
.A2(n_293),
.B(n_255),
.Y(n_320)
);

OAI32xp33_ASAP7_75t_L g286 ( 
.A1(n_238),
.A2(n_215),
.A3(n_222),
.B1(n_229),
.B2(n_214),
.Y(n_286)
);

INVxp67_ASAP7_75t_L g302 ( 
.A(n_286),
.Y(n_302)
);

OAI22xp5_ASAP7_75t_L g289 ( 
.A1(n_249),
.A2(n_213),
.B1(n_224),
.B2(n_219),
.Y(n_289)
);

OAI22xp5_ASAP7_75t_SL g292 ( 
.A1(n_241),
.A2(n_224),
.B1(n_219),
.B2(n_204),
.Y(n_292)
);

AOI22xp5_ASAP7_75t_L g316 ( 
.A1(n_292),
.A2(n_265),
.B1(n_240),
.B2(n_261),
.Y(n_316)
);

AOI21xp5_ASAP7_75t_SL g293 ( 
.A1(n_243),
.A2(n_183),
.B(n_230),
.Y(n_293)
);

NAND2xp5_ASAP7_75t_SL g294 ( 
.A(n_248),
.B(n_204),
.Y(n_294)
);

NAND2xp5_ASAP7_75t_SL g313 ( 
.A(n_294),
.B(n_250),
.Y(n_313)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_266),
.Y(n_295)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_295),
.Y(n_308)
);

AOI22xp5_ASAP7_75t_L g296 ( 
.A1(n_264),
.A2(n_220),
.B1(n_221),
.B2(n_209),
.Y(n_296)
);

OAI22xp5_ASAP7_75t_SL g321 ( 
.A1(n_296),
.A2(n_263),
.B1(n_262),
.B2(n_259),
.Y(n_321)
);

CKINVDCx20_ASAP7_75t_R g297 ( 
.A(n_274),
.Y(n_297)
);

NAND2xp5_ASAP7_75t_SL g335 ( 
.A(n_297),
.B(n_300),
.Y(n_335)
);

OAI21xp5_ASAP7_75t_L g349 ( 
.A1(n_299),
.A2(n_320),
.B(n_329),
.Y(n_349)
);

NOR2xp33_ASAP7_75t_L g300 ( 
.A(n_279),
.B(n_242),
.Y(n_300)
);

AOI21xp5_ASAP7_75t_L g301 ( 
.A1(n_269),
.A2(n_251),
.B(n_244),
.Y(n_301)
);

AOI21xp5_ASAP7_75t_L g354 ( 
.A1(n_301),
.A2(n_187),
.B(n_221),
.Y(n_354)
);

MAJIxp5_ASAP7_75t_L g304 ( 
.A(n_271),
.B(n_258),
.C(n_253),
.Y(n_304)
);

MAJIxp5_ASAP7_75t_L g357 ( 
.A(n_304),
.B(n_306),
.C(n_327),
.Y(n_357)
);

MAJIxp5_ASAP7_75t_L g306 ( 
.A(n_271),
.B(n_272),
.C(n_284),
.Y(n_306)
);

INVxp33_ASAP7_75t_L g307 ( 
.A(n_277),
.Y(n_307)
);

NOR2xp33_ASAP7_75t_L g351 ( 
.A(n_307),
.B(n_312),
.Y(n_351)
);

INVx3_ASAP7_75t_L g309 ( 
.A(n_283),
.Y(n_309)
);

INVxp67_ASAP7_75t_L g337 ( 
.A(n_309),
.Y(n_337)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_267),
.Y(n_310)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_310),
.Y(n_331)
);

INVx2_ASAP7_75t_L g311 ( 
.A(n_267),
.Y(n_311)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_311),
.Y(n_333)
);

INVxp33_ASAP7_75t_L g312 ( 
.A(n_277),
.Y(n_312)
);

CKINVDCx16_ASAP7_75t_R g336 ( 
.A(n_313),
.Y(n_336)
);

CKINVDCx20_ASAP7_75t_R g314 ( 
.A(n_274),
.Y(n_314)
);

CKINVDCx20_ASAP7_75t_R g356 ( 
.A(n_314),
.Y(n_356)
);

XNOR2xp5_ASAP7_75t_L g315 ( 
.A(n_271),
.B(n_253),
.Y(n_315)
);

XOR2xp5_ASAP7_75t_L g332 ( 
.A(n_315),
.B(n_317),
.Y(n_332)
);

OAI22xp5_ASAP7_75t_L g338 ( 
.A1(n_316),
.A2(n_288),
.B1(n_273),
.B2(n_287),
.Y(n_338)
);

XNOR2xp5_ASAP7_75t_L g317 ( 
.A(n_272),
.B(n_255),
.Y(n_317)
);

BUFx6f_ASAP7_75t_L g318 ( 
.A(n_283),
.Y(n_318)
);

INVx1_ASAP7_75t_L g348 ( 
.A(n_318),
.Y(n_348)
);

OA21x2_ASAP7_75t_L g350 ( 
.A1(n_319),
.A2(n_234),
.B(n_230),
.Y(n_350)
);

AOI22xp5_ASAP7_75t_L g330 ( 
.A1(n_321),
.A2(n_323),
.B1(n_288),
.B2(n_281),
.Y(n_330)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_291),
.Y(n_322)
);

INVx1_ASAP7_75t_L g360 ( 
.A(n_322),
.Y(n_360)
);

OAI22xp5_ASAP7_75t_SL g323 ( 
.A1(n_275),
.A2(n_256),
.B1(n_252),
.B2(n_237),
.Y(n_323)
);

NOR2xp33_ASAP7_75t_L g324 ( 
.A(n_276),
.B(n_226),
.Y(n_324)
);

NAND2xp5_ASAP7_75t_SL g345 ( 
.A(n_324),
.B(n_325),
.Y(n_345)
);

CKINVDCx20_ASAP7_75t_R g325 ( 
.A(n_276),
.Y(n_325)
);

AOI22xp5_ASAP7_75t_L g326 ( 
.A1(n_270),
.A2(n_256),
.B1(n_247),
.B2(n_252),
.Y(n_326)
);

OAI22xp5_ASAP7_75t_SL g358 ( 
.A1(n_326),
.A2(n_328),
.B1(n_113),
.B2(n_86),
.Y(n_358)
);

XOR2xp5_ASAP7_75t_L g327 ( 
.A(n_285),
.B(n_256),
.Y(n_327)
);

AOI22xp5_ASAP7_75t_L g328 ( 
.A1(n_292),
.A2(n_256),
.B1(n_220),
.B2(n_228),
.Y(n_328)
);

OAI32xp33_ASAP7_75t_L g329 ( 
.A1(n_280),
.A2(n_256),
.A3(n_210),
.B1(n_225),
.B2(n_226),
.Y(n_329)
);

OAI22xp5_ASAP7_75t_L g372 ( 
.A1(n_330),
.A2(n_340),
.B1(n_341),
.B2(n_342),
.Y(n_372)
);

XNOR2xp5_ASAP7_75t_L g334 ( 
.A(n_306),
.B(n_287),
.Y(n_334)
);

XOR2xp5_ASAP7_75t_L g369 ( 
.A(n_334),
.B(n_346),
.Y(n_369)
);

AOI22xp5_ASAP7_75t_L g364 ( 
.A1(n_338),
.A2(n_339),
.B1(n_358),
.B2(n_319),
.Y(n_364)
);

OAI22x1_ASAP7_75t_SL g339 ( 
.A1(n_302),
.A2(n_273),
.B1(n_296),
.B2(n_268),
.Y(n_339)
);

OAI22xp5_ASAP7_75t_L g340 ( 
.A1(n_305),
.A2(n_282),
.B1(n_296),
.B2(n_289),
.Y(n_340)
);

AOI22xp5_ASAP7_75t_L g341 ( 
.A1(n_323),
.A2(n_282),
.B1(n_278),
.B2(n_294),
.Y(n_341)
);

AOI22xp5_ASAP7_75t_L g342 ( 
.A1(n_302),
.A2(n_282),
.B1(n_290),
.B2(n_291),
.Y(n_342)
);

AOI22xp5_ASAP7_75t_L g343 ( 
.A1(n_305),
.A2(n_290),
.B1(n_295),
.B2(n_286),
.Y(n_343)
);

OAI22xp5_ASAP7_75t_L g383 ( 
.A1(n_343),
.A2(n_344),
.B1(n_350),
.B2(n_355),
.Y(n_383)
);

OAI22xp5_ASAP7_75t_L g344 ( 
.A1(n_326),
.A2(n_293),
.B1(n_220),
.B2(n_221),
.Y(n_344)
);

XOR2xp5_ASAP7_75t_L g346 ( 
.A(n_315),
.B(n_293),
.Y(n_346)
);

XNOR2xp5_ASAP7_75t_SL g347 ( 
.A(n_304),
.B(n_228),
.Y(n_347)
);

XNOR2xp5_ASAP7_75t_SL g366 ( 
.A(n_347),
.B(n_301),
.Y(n_366)
);

OAI21xp5_ASAP7_75t_L g352 ( 
.A1(n_299),
.A2(n_234),
.B(n_225),
.Y(n_352)
);

NOR2xp33_ASAP7_75t_L g385 ( 
.A(n_352),
.B(n_321),
.Y(n_385)
);

NAND2xp5_ASAP7_75t_SL g353 ( 
.A(n_298),
.B(n_210),
.Y(n_353)
);

NAND2xp5_ASAP7_75t_SL g367 ( 
.A(n_353),
.B(n_303),
.Y(n_367)
);

OAI22xp5_ASAP7_75t_SL g388 ( 
.A1(n_354),
.A2(n_359),
.B1(n_328),
.B2(n_318),
.Y(n_388)
);

OAI22xp5_ASAP7_75t_L g355 ( 
.A1(n_325),
.A2(n_113),
.B1(n_35),
.B2(n_42),
.Y(n_355)
);

AOI22xp5_ASAP7_75t_L g359 ( 
.A1(n_298),
.A2(n_42),
.B1(n_38),
.B2(n_35),
.Y(n_359)
);

INVx1_ASAP7_75t_L g361 ( 
.A(n_303),
.Y(n_361)
);

INVx1_ASAP7_75t_L g368 ( 
.A(n_361),
.Y(n_368)
);

INVx2_ASAP7_75t_L g362 ( 
.A(n_348),
.Y(n_362)
);

INVx1_ASAP7_75t_L g405 ( 
.A(n_362),
.Y(n_405)
);

MAJIxp5_ASAP7_75t_L g363 ( 
.A(n_357),
.B(n_317),
.C(n_320),
.Y(n_363)
);

MAJIxp5_ASAP7_75t_L g395 ( 
.A(n_363),
.B(n_370),
.C(n_377),
.Y(n_395)
);

OAI22xp5_ASAP7_75t_L g397 ( 
.A1(n_364),
.A2(n_330),
.B1(n_341),
.B2(n_383),
.Y(n_397)
);

INVx1_ASAP7_75t_L g365 ( 
.A(n_361),
.Y(n_365)
);

INVx1_ASAP7_75t_L g392 ( 
.A(n_365),
.Y(n_392)
);

XNOR2xp5_ASAP7_75t_L g404 ( 
.A(n_366),
.B(n_373),
.Y(n_404)
);

AOI22xp33_ASAP7_75t_L g410 ( 
.A1(n_367),
.A2(n_376),
.B1(n_381),
.B2(n_384),
.Y(n_410)
);

MAJIxp5_ASAP7_75t_L g370 ( 
.A(n_357),
.B(n_314),
.C(n_327),
.Y(n_370)
);

INVx1_ASAP7_75t_L g371 ( 
.A(n_345),
.Y(n_371)
);

INVx1_ASAP7_75t_L g394 ( 
.A(n_371),
.Y(n_394)
);

XNOR2xp5_ASAP7_75t_L g373 ( 
.A(n_332),
.B(n_316),
.Y(n_373)
);

INVx1_ASAP7_75t_L g374 ( 
.A(n_331),
.Y(n_374)
);

INVx1_ASAP7_75t_L g418 ( 
.A(n_374),
.Y(n_418)
);

INVx1_ASAP7_75t_L g375 ( 
.A(n_331),
.Y(n_375)
);

INVx1_ASAP7_75t_L g419 ( 
.A(n_375),
.Y(n_419)
);

INVx1_ASAP7_75t_L g376 ( 
.A(n_360),
.Y(n_376)
);

MAJIxp5_ASAP7_75t_L g377 ( 
.A(n_332),
.B(n_308),
.C(n_322),
.Y(n_377)
);

NAND2xp5_ASAP7_75t_SL g378 ( 
.A(n_335),
.B(n_336),
.Y(n_378)
);

NAND2xp5_ASAP7_75t_SL g399 ( 
.A(n_378),
.B(n_359),
.Y(n_399)
);

MAJIxp5_ASAP7_75t_L g379 ( 
.A(n_347),
.B(n_334),
.C(n_346),
.Y(n_379)
);

MAJIxp5_ASAP7_75t_L g409 ( 
.A(n_379),
.B(n_380),
.C(n_382),
.Y(n_409)
);

MAJIxp5_ASAP7_75t_L g380 ( 
.A(n_338),
.B(n_342),
.C(n_349),
.Y(n_380)
);

CKINVDCx20_ASAP7_75t_R g381 ( 
.A(n_351),
.Y(n_381)
);

MAJIxp5_ASAP7_75t_L g382 ( 
.A(n_349),
.B(n_308),
.C(n_310),
.Y(n_382)
);

INVx1_ASAP7_75t_L g384 ( 
.A(n_360),
.Y(n_384)
);

NAND2xp5_ASAP7_75t_L g393 ( 
.A(n_385),
.B(n_336),
.Y(n_393)
);

INVx1_ASAP7_75t_L g386 ( 
.A(n_355),
.Y(n_386)
);

NOR2xp33_ASAP7_75t_L g414 ( 
.A(n_386),
.B(n_389),
.Y(n_414)
);

MAJIxp5_ASAP7_75t_L g387 ( 
.A(n_356),
.B(n_311),
.C(n_309),
.Y(n_387)
);

MAJIxp5_ASAP7_75t_L g412 ( 
.A(n_387),
.B(n_390),
.C(n_391),
.Y(n_412)
);

AND2x2_ASAP7_75t_L g413 ( 
.A(n_388),
.B(n_13),
.Y(n_413)
);

INVx1_ASAP7_75t_L g389 ( 
.A(n_333),
.Y(n_389)
);

MAJIxp5_ASAP7_75t_L g390 ( 
.A(n_356),
.B(n_329),
.C(n_42),
.Y(n_390)
);

MAJIxp5_ASAP7_75t_L g391 ( 
.A(n_343),
.B(n_28),
.C(n_27),
.Y(n_391)
);

CKINVDCx5p33_ASAP7_75t_R g427 ( 
.A(n_393),
.Y(n_427)
);

NAND2xp5_ASAP7_75t_L g396 ( 
.A(n_387),
.B(n_337),
.Y(n_396)
);

INVx1_ASAP7_75t_L g424 ( 
.A(n_396),
.Y(n_424)
);

AOI22xp5_ASAP7_75t_L g420 ( 
.A1(n_397),
.A2(n_388),
.B1(n_391),
.B2(n_373),
.Y(n_420)
);

AOI22xp5_ASAP7_75t_L g398 ( 
.A1(n_372),
.A2(n_339),
.B1(n_340),
.B2(n_350),
.Y(n_398)
);

OAI22xp5_ASAP7_75t_L g423 ( 
.A1(n_398),
.A2(n_407),
.B1(n_416),
.B2(n_374),
.Y(n_423)
);

NOR2xp33_ASAP7_75t_SL g421 ( 
.A(n_399),
.B(n_376),
.Y(n_421)
);

XOR2xp5_ASAP7_75t_L g400 ( 
.A(n_369),
.B(n_350),
.Y(n_400)
);

XNOR2xp5_ASAP7_75t_L g430 ( 
.A(n_400),
.B(n_402),
.Y(n_430)
);

XNOR2x1_ASAP7_75t_L g401 ( 
.A(n_366),
.B(n_354),
.Y(n_401)
);

XNOR2xp5_ASAP7_75t_SL g444 ( 
.A(n_401),
.B(n_4),
.Y(n_444)
);

XOR2xp5_ASAP7_75t_L g402 ( 
.A(n_369),
.B(n_352),
.Y(n_402)
);

NAND2xp5_ASAP7_75t_L g403 ( 
.A(n_371),
.B(n_337),
.Y(n_403)
);

INVx1_ASAP7_75t_L g425 ( 
.A(n_403),
.Y(n_425)
);

CKINVDCx16_ASAP7_75t_R g406 ( 
.A(n_382),
.Y(n_406)
);

NOR2xp33_ASAP7_75t_L g434 ( 
.A(n_406),
.B(n_12),
.Y(n_434)
);

AOI21xp5_ASAP7_75t_L g407 ( 
.A1(n_380),
.A2(n_344),
.B(n_358),
.Y(n_407)
);

OAI21xp5_ASAP7_75t_SL g408 ( 
.A1(n_364),
.A2(n_333),
.B(n_348),
.Y(n_408)
);

AOI21xp5_ASAP7_75t_SL g443 ( 
.A1(n_408),
.A2(n_0),
.B(n_3),
.Y(n_443)
);

AOI22xp5_ASAP7_75t_SL g411 ( 
.A1(n_365),
.A2(n_27),
.B1(n_25),
.B2(n_21),
.Y(n_411)
);

OAI22xp5_ASAP7_75t_SL g438 ( 
.A1(n_411),
.A2(n_41),
.B1(n_2),
.B2(n_3),
.Y(n_438)
);

INVx1_ASAP7_75t_L g426 ( 
.A(n_413),
.Y(n_426)
);

MAJIxp5_ASAP7_75t_L g415 ( 
.A(n_370),
.B(n_25),
.C(n_41),
.Y(n_415)
);

MAJIxp5_ASAP7_75t_L g429 ( 
.A(n_415),
.B(n_363),
.C(n_379),
.Y(n_429)
);

AOI22xp5_ASAP7_75t_L g416 ( 
.A1(n_368),
.A2(n_13),
.B1(n_12),
.B2(n_2),
.Y(n_416)
);

NAND2xp5_ASAP7_75t_L g417 ( 
.A(n_390),
.B(n_377),
.Y(n_417)
);

INVx1_ASAP7_75t_L g436 ( 
.A(n_417),
.Y(n_436)
);

OAI22xp5_ASAP7_75t_SL g456 ( 
.A1(n_420),
.A2(n_398),
.B1(n_413),
.B2(n_410),
.Y(n_456)
);

NAND2xp5_ASAP7_75t_SL g455 ( 
.A(n_421),
.B(n_438),
.Y(n_455)
);

NAND2xp5_ASAP7_75t_L g422 ( 
.A(n_403),
.B(n_375),
.Y(n_422)
);

INVx1_ASAP7_75t_L g449 ( 
.A(n_422),
.Y(n_449)
);

HB1xp67_ASAP7_75t_L g451 ( 
.A(n_423),
.Y(n_451)
);

BUFx24_ASAP7_75t_SL g428 ( 
.A(n_394),
.Y(n_428)
);

NAND2xp5_ASAP7_75t_SL g454 ( 
.A(n_428),
.B(n_431),
.Y(n_454)
);

XOR2xp5_ASAP7_75t_L g448 ( 
.A(n_429),
.B(n_444),
.Y(n_448)
);

MAJIxp5_ASAP7_75t_L g431 ( 
.A(n_395),
.B(n_409),
.C(n_417),
.Y(n_431)
);

NAND2xp5_ASAP7_75t_L g432 ( 
.A(n_405),
.B(n_362),
.Y(n_432)
);

INVx1_ASAP7_75t_L g460 ( 
.A(n_432),
.Y(n_460)
);

CKINVDCx16_ASAP7_75t_R g433 ( 
.A(n_393),
.Y(n_433)
);

INVx1_ASAP7_75t_L g461 ( 
.A(n_433),
.Y(n_461)
);

NOR2xp33_ASAP7_75t_SL g445 ( 
.A(n_434),
.B(n_427),
.Y(n_445)
);

NAND2xp5_ASAP7_75t_L g435 ( 
.A(n_405),
.B(n_0),
.Y(n_435)
);

CKINVDCx20_ASAP7_75t_R g453 ( 
.A(n_435),
.Y(n_453)
);

MAJIxp5_ASAP7_75t_L g437 ( 
.A(n_395),
.B(n_41),
.C(n_1),
.Y(n_437)
);

MAJIxp5_ASAP7_75t_L g450 ( 
.A(n_437),
.B(n_440),
.C(n_442),
.Y(n_450)
);

INVx1_ASAP7_75t_L g439 ( 
.A(n_416),
.Y(n_439)
);

NAND2xp5_ASAP7_75t_L g457 ( 
.A(n_439),
.B(n_441),
.Y(n_457)
);

MAJIxp5_ASAP7_75t_L g440 ( 
.A(n_409),
.B(n_41),
.C(n_2),
.Y(n_440)
);

INVx1_ASAP7_75t_L g441 ( 
.A(n_418),
.Y(n_441)
);

MAJIxp5_ASAP7_75t_L g442 ( 
.A(n_412),
.B(n_0),
.C(n_3),
.Y(n_442)
);

OAI21xp5_ASAP7_75t_L g459 ( 
.A1(n_443),
.A2(n_438),
.B(n_418),
.Y(n_459)
);

NAND2xp5_ASAP7_75t_L g477 ( 
.A(n_445),
.B(n_452),
.Y(n_477)
);

AOI21xp5_ASAP7_75t_L g446 ( 
.A1(n_425),
.A2(n_401),
.B(n_408),
.Y(n_446)
);

AOI21xp5_ASAP7_75t_L g478 ( 
.A1(n_446),
.A2(n_462),
.B(n_5),
.Y(n_478)
);

NOR2xp33_ASAP7_75t_SL g447 ( 
.A(n_436),
.B(n_414),
.Y(n_447)
);

OAI21x1_ASAP7_75t_L g474 ( 
.A1(n_447),
.A2(n_5),
.B(n_6),
.Y(n_474)
);

MAJIxp5_ASAP7_75t_L g452 ( 
.A(n_431),
.B(n_396),
.C(n_407),
.Y(n_452)
);

AOI22xp5_ASAP7_75t_L g465 ( 
.A1(n_456),
.A2(n_458),
.B1(n_426),
.B2(n_446),
.Y(n_465)
);

OAI22xp5_ASAP7_75t_SL g458 ( 
.A1(n_420),
.A2(n_413),
.B1(n_392),
.B2(n_419),
.Y(n_458)
);

INVx1_ASAP7_75t_L g467 ( 
.A(n_459),
.Y(n_467)
);

OAI21xp5_ASAP7_75t_SL g462 ( 
.A1(n_424),
.A2(n_400),
.B(n_419),
.Y(n_462)
);

XOR2xp5_ASAP7_75t_L g463 ( 
.A(n_430),
.B(n_402),
.Y(n_463)
);

NOR2xp33_ASAP7_75t_L g473 ( 
.A(n_463),
.B(n_4),
.Y(n_473)
);

MAJIxp5_ASAP7_75t_L g464 ( 
.A(n_429),
.B(n_412),
.C(n_404),
.Y(n_464)
);

NAND2xp5_ASAP7_75t_L g481 ( 
.A(n_464),
.B(n_7),
.Y(n_481)
);

OR2x2_ASAP7_75t_L g484 ( 
.A(n_465),
.B(n_468),
.Y(n_484)
);

AOI22xp5_ASAP7_75t_L g466 ( 
.A1(n_451),
.A2(n_426),
.B1(n_422),
.B2(n_427),
.Y(n_466)
);

OAI22xp5_ASAP7_75t_SL g489 ( 
.A1(n_466),
.A2(n_470),
.B1(n_471),
.B2(n_476),
.Y(n_489)
);

AOI21xp5_ASAP7_75t_L g468 ( 
.A1(n_454),
.A2(n_440),
.B(n_437),
.Y(n_468)
);

AOI21x1_ASAP7_75t_L g469 ( 
.A1(n_461),
.A2(n_432),
.B(n_415),
.Y(n_469)
);

OAI21xp5_ASAP7_75t_SL g491 ( 
.A1(n_469),
.A2(n_449),
.B(n_460),
.Y(n_491)
);

AOI22xp5_ASAP7_75t_L g470 ( 
.A1(n_456),
.A2(n_430),
.B1(n_435),
.B2(n_404),
.Y(n_470)
);

AOI22xp5_ASAP7_75t_L g471 ( 
.A1(n_458),
.A2(n_444),
.B1(n_442),
.B2(n_443),
.Y(n_471)
);

NOR2xp67_ASAP7_75t_SL g472 ( 
.A(n_464),
.B(n_411),
.Y(n_472)
);

AOI21x1_ASAP7_75t_L g486 ( 
.A1(n_472),
.A2(n_474),
.B(n_475),
.Y(n_486)
);

NOR2xp33_ASAP7_75t_SL g493 ( 
.A(n_473),
.B(n_450),
.Y(n_493)
);

OAI21xp5_ASAP7_75t_L g475 ( 
.A1(n_462),
.A2(n_5),
.B(n_6),
.Y(n_475)
);

AOI22xp5_ASAP7_75t_L g476 ( 
.A1(n_449),
.A2(n_5),
.B1(n_6),
.B2(n_7),
.Y(n_476)
);

XOR2xp5_ASAP7_75t_L g485 ( 
.A(n_478),
.B(n_459),
.Y(n_485)
);

NOR2xp33_ASAP7_75t_L g479 ( 
.A(n_452),
.B(n_6),
.Y(n_479)
);

NAND2xp5_ASAP7_75t_L g487 ( 
.A(n_479),
.B(n_480),
.Y(n_487)
);

NOR2xp33_ASAP7_75t_L g480 ( 
.A(n_447),
.B(n_11),
.Y(n_480)
);

NAND2xp5_ASAP7_75t_L g495 ( 
.A(n_481),
.B(n_7),
.Y(n_495)
);

NOR2xp33_ASAP7_75t_L g482 ( 
.A(n_477),
.B(n_445),
.Y(n_482)
);

NAND2xp5_ASAP7_75t_L g497 ( 
.A(n_482),
.B(n_483),
.Y(n_497)
);

NOR2xp33_ASAP7_75t_L g483 ( 
.A(n_465),
.B(n_461),
.Y(n_483)
);

NAND2xp5_ASAP7_75t_L g498 ( 
.A(n_485),
.B(n_488),
.Y(n_498)
);

XOR2xp5_ASAP7_75t_L g488 ( 
.A(n_470),
.B(n_463),
.Y(n_488)
);

XOR2xp5_ASAP7_75t_L g490 ( 
.A(n_466),
.B(n_448),
.Y(n_490)
);

INVxp67_ASAP7_75t_L g504 ( 
.A(n_490),
.Y(n_504)
);

AOI21xp5_ASAP7_75t_SL g502 ( 
.A1(n_491),
.A2(n_455),
.B(n_453),
.Y(n_502)
);

NOR2xp33_ASAP7_75t_L g492 ( 
.A(n_467),
.B(n_457),
.Y(n_492)
);

NOR2xp33_ASAP7_75t_SL g505 ( 
.A(n_492),
.B(n_494),
.Y(n_505)
);

CKINVDCx20_ASAP7_75t_R g500 ( 
.A(n_493),
.Y(n_500)
);

NOR2xp33_ASAP7_75t_L g494 ( 
.A(n_478),
.B(n_457),
.Y(n_494)
);

CKINVDCx20_ASAP7_75t_R g507 ( 
.A(n_495),
.Y(n_507)
);

XOR2xp5_ASAP7_75t_L g496 ( 
.A(n_471),
.B(n_448),
.Y(n_496)
);

NOR2xp33_ASAP7_75t_L g508 ( 
.A(n_496),
.B(n_8),
.Y(n_508)
);

OAI321xp33_ASAP7_75t_L g499 ( 
.A1(n_484),
.A2(n_460),
.A3(n_453),
.B1(n_455),
.B2(n_475),
.C(n_476),
.Y(n_499)
);

AOI21xp5_ASAP7_75t_L g511 ( 
.A1(n_499),
.A2(n_501),
.B(n_506),
.Y(n_511)
);

NOR2xp67_ASAP7_75t_SL g501 ( 
.A(n_490),
.B(n_450),
.Y(n_501)
);

OAI21xp5_ASAP7_75t_L g512 ( 
.A1(n_502),
.A2(n_489),
.B(n_485),
.Y(n_512)
);

NAND3xp33_ASAP7_75t_L g503 ( 
.A(n_484),
.B(n_7),
.C(n_8),
.Y(n_503)
);

CKINVDCx20_ASAP7_75t_R g509 ( 
.A(n_503),
.Y(n_509)
);

OAI21xp5_ASAP7_75t_SL g506 ( 
.A1(n_486),
.A2(n_7),
.B(n_8),
.Y(n_506)
);

INVx1_ASAP7_75t_L g510 ( 
.A(n_508),
.Y(n_510)
);

AOI21xp5_ASAP7_75t_L g519 ( 
.A1(n_512),
.A2(n_513),
.B(n_514),
.Y(n_519)
);

AOI21xp5_ASAP7_75t_L g513 ( 
.A1(n_497),
.A2(n_496),
.B(n_488),
.Y(n_513)
);

AOI21xp5_ASAP7_75t_L g514 ( 
.A1(n_505),
.A2(n_487),
.B(n_10),
.Y(n_514)
);

AOI21xp5_ASAP7_75t_L g515 ( 
.A1(n_500),
.A2(n_9),
.B(n_10),
.Y(n_515)
);

OAI21xp5_ASAP7_75t_SL g518 ( 
.A1(n_515),
.A2(n_507),
.B(n_10),
.Y(n_518)
);

AND2x2_ASAP7_75t_L g516 ( 
.A(n_504),
.B(n_9),
.Y(n_516)
);

XNOR2xp5_ASAP7_75t_L g520 ( 
.A(n_516),
.B(n_9),
.Y(n_520)
);

MAJIxp5_ASAP7_75t_L g517 ( 
.A(n_511),
.B(n_498),
.C(n_508),
.Y(n_517)
);

NAND2xp5_ASAP7_75t_SL g522 ( 
.A(n_517),
.B(n_518),
.Y(n_522)
);

HB1xp67_ASAP7_75t_L g524 ( 
.A(n_520),
.Y(n_524)
);

OAI21xp5_ASAP7_75t_SL g521 ( 
.A1(n_509),
.A2(n_9),
.B(n_11),
.Y(n_521)
);

BUFx24_ASAP7_75t_SL g523 ( 
.A(n_521),
.Y(n_523)
);

BUFx24_ASAP7_75t_SL g525 ( 
.A(n_523),
.Y(n_525)
);

OAI21xp5_ASAP7_75t_L g527 ( 
.A1(n_525),
.A2(n_526),
.B(n_524),
.Y(n_527)
);

AOI21xp5_ASAP7_75t_SL g526 ( 
.A1(n_522),
.A2(n_519),
.B(n_510),
.Y(n_526)
);

BUFx24_ASAP7_75t_SL g528 ( 
.A(n_527),
.Y(n_528)
);


endmodule