module fake_jpeg_13512_n_472 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_472);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_472;

wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_377;
wire n_291;
wire n_236;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_17;
wire n_431;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_415;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_48;
wire n_465;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_221;
wire n_256;
wire n_454;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_429;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_305;
wire n_161;
wire n_441;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_352;
wire n_350;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_389;
wire n_457;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_384;
wire n_168;
wire n_459;
wire n_274;
wire n_24;
wire n_467;
wire n_269;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_145;
wire n_18;
wire n_20;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_344;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_199;
wire n_260;
wire n_413;
wire n_275;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_379;
wire n_114;
wire n_444;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_469;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_183;
wire n_409;
wire n_249;
wire n_412;
wire n_217;
wire n_471;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_391;
wire n_209;
wire n_22;
wire n_138;
wire n_402;
wire n_438;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

BUFx6f_ASAP7_75t_L g16 ( 
.A(n_0),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_13),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_4),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_3),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_9),
.Y(n_20)
);

BUFx2_ASAP7_75t_L g21 ( 
.A(n_3),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_2),
.Y(n_22)
);

BUFx24_ASAP7_75t_L g23 ( 
.A(n_9),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_6),
.Y(n_24)
);

INVx2_ASAP7_75t_L g25 ( 
.A(n_13),
.Y(n_25)
);

BUFx12f_ASAP7_75t_L g26 ( 
.A(n_9),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_10),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_3),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_7),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_9),
.Y(n_30)
);

INVx4_ASAP7_75t_L g31 ( 
.A(n_2),
.Y(n_31)
);

INVx8_ASAP7_75t_L g32 ( 
.A(n_13),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_4),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_1),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_2),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_1),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_0),
.Y(n_37)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_6),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_4),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_14),
.Y(n_40)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_2),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g42 ( 
.A(n_2),
.B(n_8),
.Y(n_42)
);

BUFx8_ASAP7_75t_L g43 ( 
.A(n_10),
.Y(n_43)
);

INVx6_ASAP7_75t_SL g44 ( 
.A(n_4),
.Y(n_44)
);

INVx8_ASAP7_75t_L g45 ( 
.A(n_44),
.Y(n_45)
);

INVx5_ASAP7_75t_L g112 ( 
.A(n_45),
.Y(n_112)
);

BUFx5_ASAP7_75t_L g46 ( 
.A(n_44),
.Y(n_46)
);

BUFx3_ASAP7_75t_L g104 ( 
.A(n_46),
.Y(n_104)
);

HAxp5_ASAP7_75t_SL g47 ( 
.A(n_44),
.B(n_0),
.CON(n_47),
.SN(n_47)
);

AND2x2_ASAP7_75t_L g97 ( 
.A(n_47),
.B(n_82),
.Y(n_97)
);

INVx6_ASAP7_75t_L g48 ( 
.A(n_40),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g100 ( 
.A(n_48),
.Y(n_100)
);

BUFx3_ASAP7_75t_L g49 ( 
.A(n_26),
.Y(n_49)
);

BUFx3_ASAP7_75t_L g127 ( 
.A(n_49),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_42),
.B(n_8),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_SL g116 ( 
.A(n_50),
.B(n_67),
.Y(n_116)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_16),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g139 ( 
.A(n_51),
.Y(n_139)
);

INVx3_ASAP7_75t_L g52 ( 
.A(n_43),
.Y(n_52)
);

HB1xp67_ASAP7_75t_L g129 ( 
.A(n_52),
.Y(n_129)
);

INVx2_ASAP7_75t_L g53 ( 
.A(n_25),
.Y(n_53)
);

INVx2_ASAP7_75t_L g95 ( 
.A(n_53),
.Y(n_95)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_16),
.Y(n_54)
);

INVx6_ASAP7_75t_L g105 ( 
.A(n_54),
.Y(n_105)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_16),
.Y(n_55)
);

INVx4_ASAP7_75t_L g113 ( 
.A(n_55),
.Y(n_113)
);

INVx3_ASAP7_75t_L g56 ( 
.A(n_43),
.Y(n_56)
);

INVx1_ASAP7_75t_SL g131 ( 
.A(n_56),
.Y(n_131)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_25),
.Y(n_57)
);

INVx2_ASAP7_75t_L g98 ( 
.A(n_57),
.Y(n_98)
);

INVx4_ASAP7_75t_L g58 ( 
.A(n_31),
.Y(n_58)
);

INVx3_ASAP7_75t_L g109 ( 
.A(n_58),
.Y(n_109)
);

BUFx3_ASAP7_75t_L g59 ( 
.A(n_26),
.Y(n_59)
);

INVx4_ASAP7_75t_L g123 ( 
.A(n_59),
.Y(n_123)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_16),
.Y(n_60)
);

INVx3_ASAP7_75t_L g111 ( 
.A(n_60),
.Y(n_111)
);

INVx3_ASAP7_75t_L g61 ( 
.A(n_43),
.Y(n_61)
);

INVx3_ASAP7_75t_L g122 ( 
.A(n_61),
.Y(n_122)
);

INVx3_ASAP7_75t_L g62 ( 
.A(n_43),
.Y(n_62)
);

INVx3_ASAP7_75t_L g137 ( 
.A(n_62),
.Y(n_137)
);

BUFx3_ASAP7_75t_L g63 ( 
.A(n_26),
.Y(n_63)
);

INVx3_ASAP7_75t_L g143 ( 
.A(n_63),
.Y(n_143)
);

BUFx3_ASAP7_75t_L g64 ( 
.A(n_26),
.Y(n_64)
);

INVx2_ASAP7_75t_L g107 ( 
.A(n_64),
.Y(n_107)
);

INVx3_ASAP7_75t_L g65 ( 
.A(n_43),
.Y(n_65)
);

INVx2_ASAP7_75t_L g115 ( 
.A(n_65),
.Y(n_115)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_25),
.Y(n_66)
);

INVx2_ASAP7_75t_L g121 ( 
.A(n_66),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_42),
.B(n_8),
.Y(n_67)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_22),
.Y(n_68)
);

INVx2_ASAP7_75t_L g94 ( 
.A(n_68),
.Y(n_94)
);

INVx6_ASAP7_75t_L g69 ( 
.A(n_40),
.Y(n_69)
);

INVx2_ASAP7_75t_L g108 ( 
.A(n_69),
.Y(n_108)
);

BUFx3_ASAP7_75t_L g70 ( 
.A(n_26),
.Y(n_70)
);

INVx2_ASAP7_75t_L g133 ( 
.A(n_70),
.Y(n_133)
);

BUFx6f_ASAP7_75t_L g71 ( 
.A(n_22),
.Y(n_71)
);

INVx2_ASAP7_75t_L g114 ( 
.A(n_71),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_34),
.B(n_8),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_72),
.B(n_83),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_L g73 ( 
.A(n_34),
.B(n_15),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_L g102 ( 
.A(n_73),
.B(n_86),
.Y(n_102)
);

BUFx3_ASAP7_75t_L g74 ( 
.A(n_26),
.Y(n_74)
);

INVx2_ASAP7_75t_L g134 ( 
.A(n_74),
.Y(n_134)
);

INVx11_ASAP7_75t_L g75 ( 
.A(n_23),
.Y(n_75)
);

INVx2_ASAP7_75t_L g135 ( 
.A(n_75),
.Y(n_135)
);

BUFx6f_ASAP7_75t_L g76 ( 
.A(n_22),
.Y(n_76)
);

INVx2_ASAP7_75t_L g141 ( 
.A(n_76),
.Y(n_141)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_21),
.Y(n_77)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_77),
.Y(n_99)
);

INVx3_ASAP7_75t_L g78 ( 
.A(n_43),
.Y(n_78)
);

INVx2_ASAP7_75t_L g142 ( 
.A(n_78),
.Y(n_142)
);

BUFx6f_ASAP7_75t_L g79 ( 
.A(n_22),
.Y(n_79)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_79),
.Y(n_120)
);

INVx2_ASAP7_75t_L g80 ( 
.A(n_31),
.Y(n_80)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_80),
.Y(n_125)
);

INVx4_ASAP7_75t_L g81 ( 
.A(n_31),
.Y(n_81)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_81),
.Y(n_130)
);

INVx4_ASAP7_75t_L g82 ( 
.A(n_32),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_27),
.B(n_7),
.Y(n_83)
);

BUFx12f_ASAP7_75t_L g84 ( 
.A(n_23),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_84),
.B(n_85),
.Y(n_124)
);

INVx5_ASAP7_75t_L g85 ( 
.A(n_32),
.Y(n_85)
);

BUFx6f_ASAP7_75t_L g86 ( 
.A(n_36),
.Y(n_86)
);

BUFx6f_ASAP7_75t_L g87 ( 
.A(n_36),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_L g117 ( 
.A(n_87),
.B(n_89),
.Y(n_117)
);

BUFx2_ASAP7_75t_L g88 ( 
.A(n_32),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g132 ( 
.A(n_88),
.B(n_92),
.Y(n_132)
);

BUFx6f_ASAP7_75t_L g89 ( 
.A(n_36),
.Y(n_89)
);

BUFx6f_ASAP7_75t_L g90 ( 
.A(n_36),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_L g140 ( 
.A(n_90),
.B(n_91),
.Y(n_140)
);

INVx6_ASAP7_75t_L g91 ( 
.A(n_40),
.Y(n_91)
);

BUFx6f_ASAP7_75t_L g92 ( 
.A(n_37),
.Y(n_92)
);

MAJIxp5_ASAP7_75t_L g93 ( 
.A(n_50),
.B(n_21),
.C(n_40),
.Y(n_93)
);

MAJIxp5_ASAP7_75t_L g185 ( 
.A(n_93),
.B(n_145),
.C(n_35),
.Y(n_185)
);

AOI22xp33_ASAP7_75t_SL g96 ( 
.A1(n_47),
.A2(n_32),
.B1(n_21),
.B2(n_23),
.Y(n_96)
);

AOI22xp33_ASAP7_75t_SL g157 ( 
.A1(n_96),
.A2(n_101),
.B1(n_119),
.B2(n_128),
.Y(n_157)
);

AOI22xp33_ASAP7_75t_SL g101 ( 
.A1(n_84),
.A2(n_21),
.B1(n_23),
.B2(n_37),
.Y(n_101)
);

OA22x2_ASAP7_75t_SL g103 ( 
.A1(n_67),
.A2(n_23),
.B1(n_39),
.B2(n_28),
.Y(n_103)
);

A2O1A1Ixp33_ASAP7_75t_L g163 ( 
.A1(n_103),
.A2(n_38),
.B(n_33),
.C(n_35),
.Y(n_163)
);

OAI22xp33_ASAP7_75t_L g106 ( 
.A1(n_48),
.A2(n_37),
.B1(n_23),
.B2(n_39),
.Y(n_106)
);

AOI22xp5_ASAP7_75t_L g174 ( 
.A1(n_106),
.A2(n_126),
.B1(n_41),
.B2(n_38),
.Y(n_174)
);

AOI22xp33_ASAP7_75t_L g118 ( 
.A1(n_83),
.A2(n_27),
.B1(n_37),
.B2(n_39),
.Y(n_118)
);

OAI22xp5_ASAP7_75t_L g153 ( 
.A1(n_118),
.A2(n_136),
.B1(n_18),
.B2(n_19),
.Y(n_153)
);

AOI22xp33_ASAP7_75t_SL g119 ( 
.A1(n_88),
.A2(n_27),
.B1(n_30),
.B2(n_29),
.Y(n_119)
);

OAI22xp5_ASAP7_75t_L g126 ( 
.A1(n_72),
.A2(n_28),
.B1(n_18),
.B2(n_19),
.Y(n_126)
);

AOI22xp33_ASAP7_75t_SL g128 ( 
.A1(n_45),
.A2(n_17),
.B1(n_20),
.B2(n_29),
.Y(n_128)
);

AOI22xp33_ASAP7_75t_SL g136 ( 
.A1(n_69),
.A2(n_17),
.B1(n_20),
.B2(n_29),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_L g138 ( 
.A(n_91),
.B(n_28),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_L g164 ( 
.A(n_138),
.B(n_144),
.Y(n_164)
);

NOR2xp33_ASAP7_75t_L g144 ( 
.A(n_51),
.B(n_18),
.Y(n_144)
);

MAJIxp5_ASAP7_75t_L g145 ( 
.A(n_54),
.B(n_17),
.C(n_20),
.Y(n_145)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_99),
.Y(n_146)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_146),
.Y(n_191)
);

CKINVDCx20_ASAP7_75t_R g147 ( 
.A(n_129),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_L g200 ( 
.A(n_147),
.B(n_149),
.Y(n_200)
);

OAI22xp5_ASAP7_75t_SL g148 ( 
.A1(n_93),
.A2(n_92),
.B1(n_90),
.B2(n_89),
.Y(n_148)
);

AOI22xp5_ASAP7_75t_L g211 ( 
.A1(n_148),
.A2(n_153),
.B1(n_171),
.B2(n_190),
.Y(n_211)
);

OAI32xp33_ASAP7_75t_L g149 ( 
.A1(n_102),
.A2(n_71),
.A3(n_86),
.B1(n_79),
.B2(n_76),
.Y(n_149)
);

INVx2_ASAP7_75t_L g150 ( 
.A(n_108),
.Y(n_150)
);

INVx2_ASAP7_75t_L g205 ( 
.A(n_150),
.Y(n_205)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_132),
.Y(n_151)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_151),
.Y(n_193)
);

INVx2_ASAP7_75t_L g152 ( 
.A(n_108),
.Y(n_152)
);

INVx3_ASAP7_75t_L g192 ( 
.A(n_152),
.Y(n_192)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_120),
.Y(n_154)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_154),
.Y(n_198)
);

INVx2_ASAP7_75t_L g155 ( 
.A(n_94),
.Y(n_155)
);

INVx3_ASAP7_75t_L g212 ( 
.A(n_155),
.Y(n_212)
);

INVx3_ASAP7_75t_L g156 ( 
.A(n_112),
.Y(n_156)
);

BUFx6f_ASAP7_75t_L g194 ( 
.A(n_156),
.Y(n_194)
);

CKINVDCx20_ASAP7_75t_R g158 ( 
.A(n_124),
.Y(n_158)
);

NOR2xp33_ASAP7_75t_L g218 ( 
.A(n_158),
.B(n_159),
.Y(n_218)
);

INVx2_ASAP7_75t_L g159 ( 
.A(n_94),
.Y(n_159)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_111),
.Y(n_160)
);

AND2x2_ASAP7_75t_L g202 ( 
.A(n_160),
.B(n_168),
.Y(n_202)
);

AOI21xp33_ASAP7_75t_L g161 ( 
.A1(n_110),
.A2(n_19),
.B(n_30),
.Y(n_161)
);

NOR2xp33_ASAP7_75t_SL g223 ( 
.A(n_161),
.B(n_177),
.Y(n_223)
);

XOR2xp5_ASAP7_75t_L g162 ( 
.A(n_97),
.B(n_125),
.Y(n_162)
);

MAJIxp5_ASAP7_75t_L g217 ( 
.A(n_162),
.B(n_179),
.C(n_185),
.Y(n_217)
);

NAND2xp5_ASAP7_75t_L g203 ( 
.A(n_163),
.B(n_178),
.Y(n_203)
);

INVx5_ASAP7_75t_L g165 ( 
.A(n_112),
.Y(n_165)
);

INVx13_ASAP7_75t_L g206 ( 
.A(n_165),
.Y(n_206)
);

INVx2_ASAP7_75t_SL g166 ( 
.A(n_122),
.Y(n_166)
);

BUFx24_ASAP7_75t_L g201 ( 
.A(n_166),
.Y(n_201)
);

INVx3_ASAP7_75t_L g167 ( 
.A(n_104),
.Y(n_167)
);

NOR2xp33_ASAP7_75t_L g219 ( 
.A(n_167),
.B(n_169),
.Y(n_219)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_111),
.Y(n_168)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_142),
.Y(n_169)
);

OAI21xp33_ASAP7_75t_L g170 ( 
.A1(n_97),
.A2(n_14),
.B(n_15),
.Y(n_170)
);

CKINVDCx16_ASAP7_75t_R g195 ( 
.A(n_170),
.Y(n_195)
);

OAI22xp33_ASAP7_75t_SL g171 ( 
.A1(n_103),
.A2(n_87),
.B1(n_68),
.B2(n_60),
.Y(n_171)
);

INVx4_ASAP7_75t_L g172 ( 
.A(n_143),
.Y(n_172)
);

CKINVDCx16_ASAP7_75t_R g214 ( 
.A(n_172),
.Y(n_214)
);

BUFx3_ASAP7_75t_L g173 ( 
.A(n_104),
.Y(n_173)
);

CKINVDCx16_ASAP7_75t_R g225 ( 
.A(n_173),
.Y(n_225)
);

OAI22xp5_ASAP7_75t_L g199 ( 
.A1(n_174),
.A2(n_181),
.B1(n_33),
.B2(n_105),
.Y(n_199)
);

INVx2_ASAP7_75t_L g175 ( 
.A(n_114),
.Y(n_175)
);

CKINVDCx20_ASAP7_75t_R g196 ( 
.A(n_175),
.Y(n_196)
);

INVx3_ASAP7_75t_L g176 ( 
.A(n_143),
.Y(n_176)
);

CKINVDCx20_ASAP7_75t_R g216 ( 
.A(n_176),
.Y(n_216)
);

NOR2xp33_ASAP7_75t_L g177 ( 
.A(n_116),
.B(n_30),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_L g178 ( 
.A(n_145),
.B(n_24),
.Y(n_178)
);

AND2x2_ASAP7_75t_L g179 ( 
.A(n_97),
.B(n_24),
.Y(n_179)
);

INVx2_ASAP7_75t_L g180 ( 
.A(n_114),
.Y(n_180)
);

AOI22xp33_ASAP7_75t_SL g222 ( 
.A1(n_180),
.A2(n_183),
.B1(n_187),
.B2(n_189),
.Y(n_222)
);

AOI22xp5_ASAP7_75t_L g181 ( 
.A1(n_106),
.A2(n_55),
.B1(n_41),
.B2(n_38),
.Y(n_181)
);

NOR2xp33_ASAP7_75t_L g182 ( 
.A(n_130),
.B(n_41),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_SL g215 ( 
.A(n_182),
.B(n_184),
.Y(n_215)
);

BUFx2_ASAP7_75t_L g183 ( 
.A(n_123),
.Y(n_183)
);

NOR2xp33_ASAP7_75t_L g184 ( 
.A(n_95),
.B(n_121),
.Y(n_184)
);

AND2x2_ASAP7_75t_L g186 ( 
.A(n_98),
.B(n_142),
.Y(n_186)
);

OAI21xp5_ASAP7_75t_SL g208 ( 
.A1(n_186),
.A2(n_131),
.B(n_115),
.Y(n_208)
);

BUFx10_ASAP7_75t_L g187 ( 
.A(n_127),
.Y(n_187)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_113),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_L g204 ( 
.A(n_188),
.B(n_113),
.Y(n_204)
);

INVx2_ASAP7_75t_L g189 ( 
.A(n_141),
.Y(n_189)
);

OAI22xp5_ASAP7_75t_L g190 ( 
.A1(n_103),
.A2(n_35),
.B1(n_33),
.B2(n_24),
.Y(n_190)
);

XOR2xp5_ASAP7_75t_L g197 ( 
.A(n_162),
.B(n_140),
.Y(n_197)
);

MAJIxp5_ASAP7_75t_L g246 ( 
.A(n_197),
.B(n_176),
.C(n_107),
.Y(n_246)
);

AOI22xp5_ASAP7_75t_L g233 ( 
.A1(n_199),
.A2(n_207),
.B1(n_220),
.B2(n_131),
.Y(n_233)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_204),
.Y(n_236)
);

OAI22xp5_ASAP7_75t_SL g207 ( 
.A1(n_185),
.A2(n_117),
.B1(n_141),
.B2(n_100),
.Y(n_207)
);

NAND2xp33_ASAP7_75t_SL g234 ( 
.A(n_208),
.B(n_166),
.Y(n_234)
);

AOI22xp33_ASAP7_75t_SL g209 ( 
.A1(n_151),
.A2(n_123),
.B1(n_127),
.B2(n_122),
.Y(n_209)
);

BUFx8_ASAP7_75t_L g230 ( 
.A(n_209),
.Y(n_230)
);

NAND2xp5_ASAP7_75t_L g210 ( 
.A(n_178),
.B(n_164),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_L g231 ( 
.A(n_210),
.B(n_221),
.Y(n_231)
);

AOI22xp33_ASAP7_75t_L g213 ( 
.A1(n_148),
.A2(n_105),
.B1(n_139),
.B2(n_100),
.Y(n_213)
);

OAI22xp5_ASAP7_75t_L g229 ( 
.A1(n_213),
.A2(n_224),
.B1(n_209),
.B2(n_222),
.Y(n_229)
);

OAI22xp5_ASAP7_75t_SL g220 ( 
.A1(n_157),
.A2(n_139),
.B1(n_137),
.B2(n_109),
.Y(n_220)
);

NAND2xp5_ASAP7_75t_L g221 ( 
.A(n_163),
.B(n_134),
.Y(n_221)
);

AOI22xp33_ASAP7_75t_SL g224 ( 
.A1(n_158),
.A2(n_137),
.B1(n_134),
.B2(n_133),
.Y(n_224)
);

OAI21xp5_ASAP7_75t_L g226 ( 
.A1(n_203),
.A2(n_221),
.B(n_223),
.Y(n_226)
);

OAI21xp5_ASAP7_75t_L g270 ( 
.A1(n_226),
.A2(n_228),
.B(n_241),
.Y(n_270)
);

OAI22xp5_ASAP7_75t_SL g227 ( 
.A1(n_200),
.A2(n_174),
.B1(n_149),
.B2(n_181),
.Y(n_227)
);

AOI22xp5_ASAP7_75t_L g258 ( 
.A1(n_227),
.A2(n_235),
.B1(n_238),
.B2(n_240),
.Y(n_258)
);

OAI21xp5_ASAP7_75t_L g228 ( 
.A1(n_203),
.A2(n_179),
.B(n_146),
.Y(n_228)
);

AND2x2_ASAP7_75t_L g282 ( 
.A(n_229),
.B(n_234),
.Y(n_282)
);

NAND2xp5_ASAP7_75t_L g232 ( 
.A(n_210),
.B(n_179),
.Y(n_232)
);

NAND2xp5_ASAP7_75t_L g267 ( 
.A(n_232),
.B(n_239),
.Y(n_267)
);

OAI22xp5_ASAP7_75t_L g266 ( 
.A1(n_233),
.A2(n_247),
.B1(n_196),
.B2(n_201),
.Y(n_266)
);

OAI22xp5_ASAP7_75t_L g235 ( 
.A1(n_211),
.A2(n_154),
.B1(n_156),
.B2(n_160),
.Y(n_235)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_191),
.Y(n_237)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_237),
.Y(n_265)
);

OAI22xp5_ASAP7_75t_SL g238 ( 
.A1(n_200),
.A2(n_168),
.B1(n_188),
.B2(n_152),
.Y(n_238)
);

NAND2xp5_ASAP7_75t_L g239 ( 
.A(n_207),
.B(n_186),
.Y(n_239)
);

OAI22xp5_ASAP7_75t_SL g240 ( 
.A1(n_211),
.A2(n_213),
.B1(n_217),
.B2(n_215),
.Y(n_240)
);

AOI21xp5_ASAP7_75t_SL g241 ( 
.A1(n_223),
.A2(n_187),
.B(n_186),
.Y(n_241)
);

OAI21xp5_ASAP7_75t_L g242 ( 
.A1(n_218),
.A2(n_167),
.B(n_169),
.Y(n_242)
);

AOI21xp5_ASAP7_75t_L g261 ( 
.A1(n_242),
.A2(n_208),
.B(n_202),
.Y(n_261)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_191),
.Y(n_243)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_243),
.Y(n_269)
);

OAI22xp5_ASAP7_75t_SL g244 ( 
.A1(n_217),
.A2(n_150),
.B1(n_166),
.B2(n_175),
.Y(n_244)
);

AOI22xp5_ASAP7_75t_L g277 ( 
.A1(n_244),
.A2(n_253),
.B1(n_229),
.B2(n_235),
.Y(n_277)
);

NAND2xp5_ASAP7_75t_L g245 ( 
.A(n_197),
.B(n_189),
.Y(n_245)
);

XNOR2xp5_ASAP7_75t_L g280 ( 
.A(n_245),
.B(n_246),
.Y(n_280)
);

AOI22xp5_ASAP7_75t_L g247 ( 
.A1(n_199),
.A2(n_155),
.B1(n_180),
.B2(n_159),
.Y(n_247)
);

XNOR2xp5_ASAP7_75t_SL g248 ( 
.A(n_215),
.B(n_187),
.Y(n_248)
);

XOR2xp5_ASAP7_75t_L g257 ( 
.A(n_248),
.B(n_252),
.Y(n_257)
);

INVx4_ASAP7_75t_L g249 ( 
.A(n_194),
.Y(n_249)
);

INVx2_ASAP7_75t_L g286 ( 
.A(n_249),
.Y(n_286)
);

CKINVDCx20_ASAP7_75t_R g250 ( 
.A(n_202),
.Y(n_250)
);

NOR2xp33_ASAP7_75t_L g264 ( 
.A(n_250),
.B(n_256),
.Y(n_264)
);

O2A1O1Ixp33_ASAP7_75t_L g251 ( 
.A1(n_201),
.A2(n_187),
.B(n_165),
.C(n_135),
.Y(n_251)
);

OAI21xp33_ASAP7_75t_SL g274 ( 
.A1(n_251),
.A2(n_201),
.B(n_205),
.Y(n_274)
);

XOR2xp5_ASAP7_75t_L g252 ( 
.A(n_218),
.B(n_172),
.Y(n_252)
);

OAI22xp5_ASAP7_75t_SL g253 ( 
.A1(n_195),
.A2(n_193),
.B1(n_224),
.B2(n_220),
.Y(n_253)
);

A2O1A1O1Ixp25_ASAP7_75t_L g254 ( 
.A1(n_195),
.A2(n_183),
.B(n_173),
.C(n_109),
.D(n_135),
.Y(n_254)
);

INVxp67_ASAP7_75t_L g272 ( 
.A(n_254),
.Y(n_272)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_198),
.Y(n_255)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_255),
.Y(n_276)
);

NOR2xp33_ASAP7_75t_L g256 ( 
.A(n_193),
.B(n_7),
.Y(n_256)
);

OAI22xp5_ASAP7_75t_SL g259 ( 
.A1(n_233),
.A2(n_204),
.B1(n_219),
.B2(n_198),
.Y(n_259)
);

AOI22xp5_ASAP7_75t_L g298 ( 
.A1(n_259),
.A2(n_260),
.B1(n_266),
.B2(n_271),
.Y(n_298)
);

OAI22xp5_ASAP7_75t_SL g260 ( 
.A1(n_231),
.A2(n_219),
.B1(n_216),
.B2(n_194),
.Y(n_260)
);

OAI21xp5_ASAP7_75t_SL g297 ( 
.A1(n_261),
.A2(n_278),
.B(n_281),
.Y(n_297)
);

XOR2xp5_ASAP7_75t_L g262 ( 
.A(n_231),
.B(n_202),
.Y(n_262)
);

MAJIxp5_ASAP7_75t_L g288 ( 
.A(n_262),
.B(n_268),
.C(n_248),
.Y(n_288)
);

CKINVDCx20_ASAP7_75t_R g263 ( 
.A(n_256),
.Y(n_263)
);

NOR2xp33_ASAP7_75t_L g293 ( 
.A(n_263),
.B(n_275),
.Y(n_293)
);

XOR2xp5_ASAP7_75t_L g268 ( 
.A(n_226),
.B(n_202),
.Y(n_268)
);

OAI22xp5_ASAP7_75t_SL g271 ( 
.A1(n_239),
.A2(n_216),
.B1(n_194),
.B2(n_196),
.Y(n_271)
);

INVxp67_ASAP7_75t_L g273 ( 
.A(n_241),
.Y(n_273)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_273),
.Y(n_311)
);

AOI22xp5_ASAP7_75t_L g310 ( 
.A1(n_274),
.A2(n_251),
.B1(n_230),
.B2(n_254),
.Y(n_310)
);

CKINVDCx16_ASAP7_75t_R g275 ( 
.A(n_242),
.Y(n_275)
);

OAI22xp5_ASAP7_75t_L g300 ( 
.A1(n_277),
.A2(n_279),
.B1(n_236),
.B2(n_247),
.Y(n_300)
);

AOI22xp5_ASAP7_75t_SL g278 ( 
.A1(n_253),
.A2(n_225),
.B1(n_214),
.B2(n_201),
.Y(n_278)
);

AOI22xp5_ASAP7_75t_L g279 ( 
.A1(n_227),
.A2(n_214),
.B1(n_212),
.B2(n_192),
.Y(n_279)
);

AOI22x1_ASAP7_75t_SL g281 ( 
.A1(n_238),
.A2(n_201),
.B1(n_225),
.B2(n_206),
.Y(n_281)
);

AOI21xp5_ASAP7_75t_L g283 ( 
.A1(n_234),
.A2(n_192),
.B(n_206),
.Y(n_283)
);

OAI21xp5_ASAP7_75t_SL g313 ( 
.A1(n_283),
.A2(n_285),
.B(n_251),
.Y(n_313)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_237),
.Y(n_284)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_284),
.Y(n_290)
);

AOI21xp5_ASAP7_75t_L g285 ( 
.A1(n_230),
.A2(n_192),
.B(n_206),
.Y(n_285)
);

INVx2_ASAP7_75t_L g287 ( 
.A(n_265),
.Y(n_287)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_287),
.Y(n_318)
);

MAJIxp5_ASAP7_75t_L g323 ( 
.A(n_288),
.B(n_294),
.C(n_296),
.Y(n_323)
);

XNOR2xp5_ASAP7_75t_L g289 ( 
.A(n_280),
.B(n_246),
.Y(n_289)
);

MAJIxp5_ASAP7_75t_L g341 ( 
.A(n_289),
.B(n_295),
.C(n_301),
.Y(n_341)
);

OAI22xp5_ASAP7_75t_SL g291 ( 
.A1(n_258),
.A2(n_236),
.B1(n_240),
.B2(n_241),
.Y(n_291)
);

AOI22xp5_ASAP7_75t_L g332 ( 
.A1(n_291),
.A2(n_300),
.B1(n_304),
.B2(n_316),
.Y(n_332)
);

BUFx3_ASAP7_75t_L g292 ( 
.A(n_286),
.Y(n_292)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_292),
.Y(n_320)
);

XNOR2xp5_ASAP7_75t_SL g294 ( 
.A(n_280),
.B(n_232),
.Y(n_294)
);

MAJIxp5_ASAP7_75t_L g295 ( 
.A(n_257),
.B(n_268),
.C(n_262),
.Y(n_295)
);

XNOR2xp5_ASAP7_75t_SL g296 ( 
.A(n_257),
.B(n_267),
.Y(n_296)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_265),
.Y(n_299)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_299),
.Y(n_324)
);

MAJIxp5_ASAP7_75t_L g301 ( 
.A(n_270),
.B(n_245),
.C(n_267),
.Y(n_301)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_269),
.Y(n_302)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_302),
.Y(n_334)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_269),
.Y(n_303)
);

NAND2xp5_ASAP7_75t_L g328 ( 
.A(n_303),
.B(n_305),
.Y(n_328)
);

OAI22xp5_ASAP7_75t_SL g304 ( 
.A1(n_258),
.A2(n_228),
.B1(n_250),
.B2(n_230),
.Y(n_304)
);

NAND2xp5_ASAP7_75t_L g305 ( 
.A(n_263),
.B(n_252),
.Y(n_305)
);

INVxp67_ASAP7_75t_L g306 ( 
.A(n_283),
.Y(n_306)
);

NAND2xp5_ASAP7_75t_L g342 ( 
.A(n_306),
.B(n_315),
.Y(n_342)
);

MAJIxp5_ASAP7_75t_L g307 ( 
.A(n_270),
.B(n_244),
.C(n_255),
.Y(n_307)
);

MAJIxp5_ASAP7_75t_L g344 ( 
.A(n_307),
.B(n_10),
.C(n_14),
.Y(n_344)
);

CKINVDCx20_ASAP7_75t_R g308 ( 
.A(n_264),
.Y(n_308)
);

NOR2xp33_ASAP7_75t_SL g333 ( 
.A(n_308),
.B(n_309),
.Y(n_333)
);

NOR2xp33_ASAP7_75t_L g309 ( 
.A(n_264),
.B(n_243),
.Y(n_309)
);

AOI21xp5_ASAP7_75t_L g325 ( 
.A1(n_310),
.A2(n_313),
.B(n_297),
.Y(n_325)
);

XOR2xp5_ASAP7_75t_L g312 ( 
.A(n_259),
.B(n_254),
.Y(n_312)
);

MAJIxp5_ASAP7_75t_L g343 ( 
.A(n_312),
.B(n_317),
.C(n_7),
.Y(n_343)
);

AOI22xp5_ASAP7_75t_L g314 ( 
.A1(n_272),
.A2(n_230),
.B1(n_249),
.B2(n_212),
.Y(n_314)
);

OAI22xp5_ASAP7_75t_SL g337 ( 
.A1(n_314),
.A2(n_279),
.B1(n_261),
.B2(n_274),
.Y(n_337)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_276),
.Y(n_315)
);

OAI22xp5_ASAP7_75t_SL g316 ( 
.A1(n_277),
.A2(n_249),
.B1(n_212),
.B2(n_205),
.Y(n_316)
);

XOR2x2_ASAP7_75t_L g317 ( 
.A(n_282),
.B(n_260),
.Y(n_317)
);

FAx1_ASAP7_75t_SL g319 ( 
.A(n_301),
.B(n_288),
.CI(n_295),
.CON(n_319),
.SN(n_319)
);

NOR2xp33_ASAP7_75t_L g353 ( 
.A(n_319),
.B(n_321),
.Y(n_353)
);

CKINVDCx20_ASAP7_75t_R g321 ( 
.A(n_293),
.Y(n_321)
);

INVxp67_ASAP7_75t_L g322 ( 
.A(n_304),
.Y(n_322)
);

INVx1_ASAP7_75t_L g350 ( 
.A(n_322),
.Y(n_350)
);

OAI21xp5_ASAP7_75t_SL g364 ( 
.A1(n_325),
.A2(n_326),
.B(n_329),
.Y(n_364)
);

AOI21xp5_ASAP7_75t_L g326 ( 
.A1(n_306),
.A2(n_282),
.B(n_285),
.Y(n_326)
);

CKINVDCx20_ASAP7_75t_R g327 ( 
.A(n_287),
.Y(n_327)
);

NOR2xp33_ASAP7_75t_L g368 ( 
.A(n_327),
.B(n_330),
.Y(n_368)
);

AOI22xp5_ASAP7_75t_SL g329 ( 
.A1(n_311),
.A2(n_282),
.B1(n_275),
.B2(n_271),
.Y(n_329)
);

CKINVDCx20_ASAP7_75t_R g330 ( 
.A(n_290),
.Y(n_330)
);

CKINVDCx20_ASAP7_75t_R g331 ( 
.A(n_290),
.Y(n_331)
);

NAND2xp5_ASAP7_75t_SL g347 ( 
.A(n_331),
.B(n_336),
.Y(n_347)
);

AOI21xp5_ASAP7_75t_L g335 ( 
.A1(n_297),
.A2(n_278),
.B(n_281),
.Y(n_335)
);

OAI21xp5_ASAP7_75t_L g371 ( 
.A1(n_335),
.A2(n_346),
.B(n_11),
.Y(n_371)
);

NOR3xp33_ASAP7_75t_SL g336 ( 
.A(n_305),
.B(n_276),
.C(n_284),
.Y(n_336)
);

AOI22xp5_ASAP7_75t_L g349 ( 
.A1(n_337),
.A2(n_317),
.B1(n_312),
.B2(n_316),
.Y(n_349)
);

CKINVDCx20_ASAP7_75t_R g338 ( 
.A(n_299),
.Y(n_338)
);

NAND2xp5_ASAP7_75t_SL g357 ( 
.A(n_338),
.B(n_340),
.Y(n_357)
);

AOI22xp5_ASAP7_75t_L g339 ( 
.A1(n_291),
.A2(n_266),
.B1(n_281),
.B2(n_286),
.Y(n_339)
);

OAI22xp5_ASAP7_75t_SL g370 ( 
.A1(n_339),
.A2(n_3),
.B1(n_4),
.B2(n_5),
.Y(n_370)
);

CKINVDCx20_ASAP7_75t_R g340 ( 
.A(n_302),
.Y(n_340)
);

XOR2xp5_ASAP7_75t_L g358 ( 
.A(n_343),
.B(n_315),
.Y(n_358)
);

MAJIxp5_ASAP7_75t_L g348 ( 
.A(n_344),
.B(n_294),
.C(n_307),
.Y(n_348)
);

BUFx24_ASAP7_75t_SL g345 ( 
.A(n_289),
.Y(n_345)
);

INVx1_ASAP7_75t_L g360 ( 
.A(n_345),
.Y(n_360)
);

OAI21xp5_ASAP7_75t_L g346 ( 
.A1(n_313),
.A2(n_10),
.B(n_14),
.Y(n_346)
);

NAND2xp5_ASAP7_75t_L g376 ( 
.A(n_348),
.B(n_355),
.Y(n_376)
);

OAI22xp5_ASAP7_75t_SL g378 ( 
.A1(n_349),
.A2(n_369),
.B1(n_329),
.B2(n_339),
.Y(n_378)
);

INVx2_ASAP7_75t_SL g351 ( 
.A(n_318),
.Y(n_351)
);

INVx1_ASAP7_75t_L g381 ( 
.A(n_351),
.Y(n_381)
);

MAJIxp5_ASAP7_75t_L g352 ( 
.A(n_341),
.B(n_296),
.C(n_298),
.Y(n_352)
);

MAJIxp5_ASAP7_75t_L g374 ( 
.A(n_352),
.B(n_365),
.C(n_344),
.Y(n_374)
);

XNOR2xp5_ASAP7_75t_L g354 ( 
.A(n_341),
.B(n_323),
.Y(n_354)
);

XNOR2xp5_ASAP7_75t_L g373 ( 
.A(n_354),
.B(n_319),
.Y(n_373)
);

BUFx2_ASAP7_75t_L g355 ( 
.A(n_320),
.Y(n_355)
);

OAI22xp5_ASAP7_75t_L g356 ( 
.A1(n_321),
.A2(n_298),
.B1(n_310),
.B2(n_314),
.Y(n_356)
);

INVx1_ASAP7_75t_L g386 ( 
.A(n_356),
.Y(n_386)
);

NAND2xp5_ASAP7_75t_SL g375 ( 
.A(n_358),
.B(n_366),
.Y(n_375)
);

XOR2xp5_ASAP7_75t_L g359 ( 
.A(n_341),
.B(n_303),
.Y(n_359)
);

XOR2xp5_ASAP7_75t_L g377 ( 
.A(n_359),
.B(n_367),
.Y(n_377)
);

AO21x2_ASAP7_75t_L g361 ( 
.A1(n_342),
.A2(n_292),
.B(n_1),
.Y(n_361)
);

OAI22xp5_ASAP7_75t_L g389 ( 
.A1(n_361),
.A2(n_372),
.B1(n_340),
.B2(n_331),
.Y(n_389)
);

INVx1_ASAP7_75t_L g362 ( 
.A(n_328),
.Y(n_362)
);

INVx1_ASAP7_75t_L g390 ( 
.A(n_362),
.Y(n_390)
);

OAI22xp5_ASAP7_75t_L g363 ( 
.A1(n_332),
.A2(n_15),
.B1(n_13),
.B2(n_12),
.Y(n_363)
);

INVx1_ASAP7_75t_L g394 ( 
.A(n_363),
.Y(n_394)
);

MAJIxp5_ASAP7_75t_L g365 ( 
.A(n_323),
.B(n_0),
.C(n_1),
.Y(n_365)
);

INVx1_ASAP7_75t_L g366 ( 
.A(n_333),
.Y(n_366)
);

XOR2xp5_ASAP7_75t_L g367 ( 
.A(n_328),
.B(n_12),
.Y(n_367)
);

AOI22xp5_ASAP7_75t_L g369 ( 
.A1(n_337),
.A2(n_0),
.B1(n_1),
.B2(n_3),
.Y(n_369)
);

AOI22xp5_ASAP7_75t_L g384 ( 
.A1(n_370),
.A2(n_324),
.B1(n_334),
.B2(n_338),
.Y(n_384)
);

OAI21xp5_ASAP7_75t_L g391 ( 
.A1(n_371),
.A2(n_346),
.B(n_330),
.Y(n_391)
);

INVx1_ASAP7_75t_L g372 ( 
.A(n_324),
.Y(n_372)
);

MAJIxp5_ASAP7_75t_L g406 ( 
.A(n_373),
.B(n_380),
.C(n_382),
.Y(n_406)
);

XNOR2xp5_ASAP7_75t_L g405 ( 
.A(n_374),
.B(n_379),
.Y(n_405)
);

AOI22xp5_ASAP7_75t_L g399 ( 
.A1(n_378),
.A2(n_370),
.B1(n_349),
.B2(n_351),
.Y(n_399)
);

XNOR2xp5_ASAP7_75t_L g379 ( 
.A(n_354),
.B(n_343),
.Y(n_379)
);

MAJIxp5_ASAP7_75t_L g380 ( 
.A(n_359),
.B(n_344),
.C(n_325),
.Y(n_380)
);

MAJIxp5_ASAP7_75t_L g382 ( 
.A(n_352),
.B(n_319),
.C(n_342),
.Y(n_382)
);

XOR2xp5_ASAP7_75t_L g383 ( 
.A(n_348),
.B(n_332),
.Y(n_383)
);

NOR2xp67_ASAP7_75t_SL g396 ( 
.A(n_383),
.B(n_388),
.Y(n_396)
);

INVx1_ASAP7_75t_L g397 ( 
.A(n_384),
.Y(n_397)
);

NOR2x1_ASAP7_75t_L g385 ( 
.A(n_362),
.B(n_333),
.Y(n_385)
);

INVx1_ASAP7_75t_L g403 ( 
.A(n_385),
.Y(n_403)
);

MAJIxp5_ASAP7_75t_L g387 ( 
.A(n_358),
.B(n_319),
.C(n_335),
.Y(n_387)
);

MAJIxp5_ASAP7_75t_L g412 ( 
.A(n_387),
.B(n_392),
.C(n_365),
.Y(n_412)
);

XOR2xp5_ASAP7_75t_L g388 ( 
.A(n_364),
.B(n_326),
.Y(n_388)
);

INVx1_ASAP7_75t_L g400 ( 
.A(n_389),
.Y(n_400)
);

INVx1_ASAP7_75t_L g404 ( 
.A(n_391),
.Y(n_404)
);

MAJIxp5_ASAP7_75t_L g392 ( 
.A(n_353),
.B(n_327),
.C(n_318),
.Y(n_392)
);

XOR2xp5_ASAP7_75t_L g393 ( 
.A(n_364),
.B(n_336),
.Y(n_393)
);

XNOR2xp5_ASAP7_75t_L g414 ( 
.A(n_393),
.B(n_369),
.Y(n_414)
);

OAI22xp5_ASAP7_75t_SL g395 ( 
.A1(n_350),
.A2(n_334),
.B1(n_336),
.B2(n_320),
.Y(n_395)
);

INVx1_ASAP7_75t_L g408 ( 
.A(n_395),
.Y(n_408)
);

AOI21xp33_ASAP7_75t_L g398 ( 
.A1(n_376),
.A2(n_347),
.B(n_368),
.Y(n_398)
);

NOR2xp33_ASAP7_75t_SL g417 ( 
.A(n_398),
.B(n_379),
.Y(n_417)
);

INVx1_ASAP7_75t_L g418 ( 
.A(n_399),
.Y(n_418)
);

NAND2xp5_ASAP7_75t_L g401 ( 
.A(n_384),
.B(n_357),
.Y(n_401)
);

INVx1_ASAP7_75t_L g419 ( 
.A(n_401),
.Y(n_419)
);

OAI22xp5_ASAP7_75t_SL g402 ( 
.A1(n_386),
.A2(n_390),
.B1(n_392),
.B2(n_387),
.Y(n_402)
);

INVx1_ASAP7_75t_L g429 ( 
.A(n_402),
.Y(n_429)
);

CKINVDCx14_ASAP7_75t_R g407 ( 
.A(n_375),
.Y(n_407)
);

INVxp67_ASAP7_75t_SL g428 ( 
.A(n_407),
.Y(n_428)
);

INVx1_ASAP7_75t_L g409 ( 
.A(n_385),
.Y(n_409)
);

INVx1_ASAP7_75t_L g430 ( 
.A(n_409),
.Y(n_430)
);

AOI21xp5_ASAP7_75t_L g410 ( 
.A1(n_393),
.A2(n_371),
.B(n_351),
.Y(n_410)
);

AOI21xp5_ASAP7_75t_L g420 ( 
.A1(n_410),
.A2(n_414),
.B(n_391),
.Y(n_420)
);

INVx1_ASAP7_75t_L g411 ( 
.A(n_381),
.Y(n_411)
);

INVx1_ASAP7_75t_L g422 ( 
.A(n_411),
.Y(n_422)
);

MAJIxp5_ASAP7_75t_L g415 ( 
.A(n_412),
.B(n_380),
.C(n_374),
.Y(n_415)
);

FAx1_ASAP7_75t_SL g413 ( 
.A(n_382),
.B(n_367),
.CI(n_361),
.CON(n_413),
.SN(n_413)
);

AO21x1_ASAP7_75t_L g426 ( 
.A1(n_413),
.A2(n_361),
.B(n_394),
.Y(n_426)
);

NAND2xp5_ASAP7_75t_L g440 ( 
.A(n_415),
.B(n_416),
.Y(n_440)
);

MAJIxp5_ASAP7_75t_L g416 ( 
.A(n_405),
.B(n_383),
.C(n_373),
.Y(n_416)
);

NOR2xp33_ASAP7_75t_SL g432 ( 
.A(n_417),
.B(n_427),
.Y(n_432)
);

XOR2xp5_ASAP7_75t_L g436 ( 
.A(n_420),
.B(n_414),
.Y(n_436)
);

MAJIxp5_ASAP7_75t_L g421 ( 
.A(n_405),
.B(n_377),
.C(n_388),
.Y(n_421)
);

NAND2xp5_ASAP7_75t_L g443 ( 
.A(n_421),
.B(n_423),
.Y(n_443)
);

MAJIxp5_ASAP7_75t_L g423 ( 
.A(n_412),
.B(n_406),
.C(n_402),
.Y(n_423)
);

AOI21xp5_ASAP7_75t_L g424 ( 
.A1(n_403),
.A2(n_378),
.B(n_372),
.Y(n_424)
);

OAI21xp5_ASAP7_75t_L g431 ( 
.A1(n_424),
.A2(n_401),
.B(n_410),
.Y(n_431)
);

MAJIxp5_ASAP7_75t_L g425 ( 
.A(n_406),
.B(n_377),
.C(n_355),
.Y(n_425)
);

MAJIxp5_ASAP7_75t_L g442 ( 
.A(n_425),
.B(n_5),
.C(n_6),
.Y(n_442)
);

OAI22xp5_ASAP7_75t_SL g433 ( 
.A1(n_426),
.A2(n_400),
.B1(n_397),
.B2(n_404),
.Y(n_433)
);

NOR2xp33_ASAP7_75t_SL g427 ( 
.A(n_404),
.B(n_360),
.Y(n_427)
);

INVx1_ASAP7_75t_L g454 ( 
.A(n_431),
.Y(n_454)
);

NAND2xp5_ASAP7_75t_L g448 ( 
.A(n_433),
.B(n_434),
.Y(n_448)
);

NOR2xp33_ASAP7_75t_L g434 ( 
.A(n_423),
.B(n_408),
.Y(n_434)
);

OAI22xp5_ASAP7_75t_SL g435 ( 
.A1(n_429),
.A2(n_397),
.B1(n_400),
.B2(n_399),
.Y(n_435)
);

NAND2xp5_ASAP7_75t_L g451 ( 
.A(n_435),
.B(n_438),
.Y(n_451)
);

XNOR2xp5_ASAP7_75t_SL g445 ( 
.A(n_436),
.B(n_419),
.Y(n_445)
);

NOR2xp33_ASAP7_75t_SL g437 ( 
.A(n_430),
.B(n_396),
.Y(n_437)
);

NAND2xp5_ASAP7_75t_SL g452 ( 
.A(n_437),
.B(n_442),
.Y(n_452)
);

XNOR2xp5_ASAP7_75t_L g438 ( 
.A(n_425),
.B(n_413),
.Y(n_438)
);

OAI22xp5_ASAP7_75t_L g439 ( 
.A1(n_428),
.A2(n_361),
.B1(n_413),
.B2(n_11),
.Y(n_439)
);

NAND2xp5_ASAP7_75t_L g455 ( 
.A(n_439),
.B(n_441),
.Y(n_455)
);

NOR2xp33_ASAP7_75t_L g441 ( 
.A(n_418),
.B(n_361),
.Y(n_441)
);

NOR2xp33_ASAP7_75t_L g444 ( 
.A(n_418),
.B(n_15),
.Y(n_444)
);

NOR2xp33_ASAP7_75t_L g446 ( 
.A(n_444),
.B(n_422),
.Y(n_446)
);

XOR2xp5_ASAP7_75t_L g461 ( 
.A(n_445),
.B(n_431),
.Y(n_461)
);

NOR2xp33_ASAP7_75t_L g458 ( 
.A(n_446),
.B(n_442),
.Y(n_458)
);

NOR2xp33_ASAP7_75t_L g447 ( 
.A(n_440),
.B(n_432),
.Y(n_447)
);

NOR2xp33_ASAP7_75t_SL g456 ( 
.A(n_447),
.B(n_453),
.Y(n_456)
);

OAI21xp5_ASAP7_75t_SL g449 ( 
.A1(n_443),
.A2(n_415),
.B(n_416),
.Y(n_449)
);

AOI21xp5_ASAP7_75t_L g460 ( 
.A1(n_449),
.A2(n_450),
.B(n_438),
.Y(n_460)
);

MAJIxp5_ASAP7_75t_L g450 ( 
.A(n_436),
.B(n_421),
.C(n_424),
.Y(n_450)
);

NOR2xp33_ASAP7_75t_L g453 ( 
.A(n_435),
.B(n_422),
.Y(n_453)
);

INVxp67_ASAP7_75t_L g457 ( 
.A(n_450),
.Y(n_457)
);

AO21x1_ASAP7_75t_L g463 ( 
.A1(n_457),
.A2(n_458),
.B(n_462),
.Y(n_463)
);

NOR2xp33_ASAP7_75t_L g459 ( 
.A(n_452),
.B(n_433),
.Y(n_459)
);

AOI21xp5_ASAP7_75t_L g464 ( 
.A1(n_459),
.A2(n_460),
.B(n_461),
.Y(n_464)
);

OAI21xp5_ASAP7_75t_L g462 ( 
.A1(n_454),
.A2(n_420),
.B(n_426),
.Y(n_462)
);

MAJIxp5_ASAP7_75t_L g465 ( 
.A(n_457),
.B(n_451),
.C(n_448),
.Y(n_465)
);

OAI21xp5_ASAP7_75t_L g467 ( 
.A1(n_465),
.A2(n_466),
.B(n_11),
.Y(n_467)
);

OAI21xp5_ASAP7_75t_SL g466 ( 
.A1(n_456),
.A2(n_455),
.B(n_445),
.Y(n_466)
);

MAJIxp5_ASAP7_75t_L g469 ( 
.A(n_467),
.B(n_468),
.C(n_463),
.Y(n_469)
);

OAI21xp5_ASAP7_75t_SL g468 ( 
.A1(n_464),
.A2(n_11),
.B(n_12),
.Y(n_468)
);

OAI21xp5_ASAP7_75t_L g470 ( 
.A1(n_469),
.A2(n_12),
.B(n_5),
.Y(n_470)
);

OAI22xp33_ASAP7_75t_R g471 ( 
.A1(n_470),
.A2(n_5),
.B1(n_6),
.B2(n_403),
.Y(n_471)
);

XOR2xp5_ASAP7_75t_L g472 ( 
.A(n_471),
.B(n_5),
.Y(n_472)
);


endmodule