module fake_netlist_6_1697_n_1228 (n_52, n_16, n_1, n_91, n_119, n_46, n_146, n_163, n_18, n_21, n_147, n_154, n_88, n_3, n_98, n_113, n_39, n_63, n_73, n_4, n_148, n_138, n_22, n_161, n_68, n_166, n_28, n_50, n_158, n_49, n_7, n_83, n_5, n_101, n_167, n_144, n_174, n_127, n_125, n_153, n_168, n_77, n_156, n_149, n_152, n_106, n_92, n_145, n_42, n_133, n_96, n_8, n_90, n_160, n_24, n_105, n_131, n_54, n_132, n_102, n_0, n_87, n_32, n_66, n_85, n_99, n_78, n_84, n_130, n_164, n_100, n_129, n_13, n_121, n_11, n_137, n_17, n_23, n_142, n_20, n_143, n_2, n_19, n_47, n_62, n_29, n_155, n_75, n_109, n_150, n_122, n_45, n_34, n_140, n_70, n_120, n_37, n_15, n_67, n_33, n_82, n_27, n_38, n_110, n_151, n_61, n_112, n_172, n_81, n_59, n_76, n_36, n_26, n_124, n_55, n_126, n_94, n_97, n_108, n_58, n_116, n_64, n_117, n_118, n_175, n_48, n_65, n_25, n_40, n_93, n_80, n_141, n_135, n_165, n_139, n_41, n_134, n_114, n_86, n_104, n_95, n_9, n_107, n_10, n_71, n_74, n_6, n_14, n_123, n_136, n_72, n_89, n_173, n_103, n_111, n_60, n_159, n_157, n_162, n_170, n_35, n_115, n_12, n_69, n_128, n_30, n_79, n_43, n_171, n_31, n_57, n_169, n_53, n_51, n_44, n_56, n_1228);

input n_52;
input n_16;
input n_1;
input n_91;
input n_119;
input n_46;
input n_146;
input n_163;
input n_18;
input n_21;
input n_147;
input n_154;
input n_88;
input n_3;
input n_98;
input n_113;
input n_39;
input n_63;
input n_73;
input n_4;
input n_148;
input n_138;
input n_22;
input n_161;
input n_68;
input n_166;
input n_28;
input n_50;
input n_158;
input n_49;
input n_7;
input n_83;
input n_5;
input n_101;
input n_167;
input n_144;
input n_174;
input n_127;
input n_125;
input n_153;
input n_168;
input n_77;
input n_156;
input n_149;
input n_152;
input n_106;
input n_92;
input n_145;
input n_42;
input n_133;
input n_96;
input n_8;
input n_90;
input n_160;
input n_24;
input n_105;
input n_131;
input n_54;
input n_132;
input n_102;
input n_0;
input n_87;
input n_32;
input n_66;
input n_85;
input n_99;
input n_78;
input n_84;
input n_130;
input n_164;
input n_100;
input n_129;
input n_13;
input n_121;
input n_11;
input n_137;
input n_17;
input n_23;
input n_142;
input n_20;
input n_143;
input n_2;
input n_19;
input n_47;
input n_62;
input n_29;
input n_155;
input n_75;
input n_109;
input n_150;
input n_122;
input n_45;
input n_34;
input n_140;
input n_70;
input n_120;
input n_37;
input n_15;
input n_67;
input n_33;
input n_82;
input n_27;
input n_38;
input n_110;
input n_151;
input n_61;
input n_112;
input n_172;
input n_81;
input n_59;
input n_76;
input n_36;
input n_26;
input n_124;
input n_55;
input n_126;
input n_94;
input n_97;
input n_108;
input n_58;
input n_116;
input n_64;
input n_117;
input n_118;
input n_175;
input n_48;
input n_65;
input n_25;
input n_40;
input n_93;
input n_80;
input n_141;
input n_135;
input n_165;
input n_139;
input n_41;
input n_134;
input n_114;
input n_86;
input n_104;
input n_95;
input n_9;
input n_107;
input n_10;
input n_71;
input n_74;
input n_6;
input n_14;
input n_123;
input n_136;
input n_72;
input n_89;
input n_173;
input n_103;
input n_111;
input n_60;
input n_159;
input n_157;
input n_162;
input n_170;
input n_35;
input n_115;
input n_12;
input n_69;
input n_128;
input n_30;
input n_79;
input n_43;
input n_171;
input n_31;
input n_57;
input n_169;
input n_53;
input n_51;
input n_44;
input n_56;

output n_1228;

wire n_992;
wire n_591;
wire n_435;
wire n_1115;
wire n_793;
wire n_326;
wire n_801;
wire n_256;
wire n_853;
wire n_440;
wire n_587;
wire n_695;
wire n_507;
wire n_968;
wire n_909;
wire n_580;
wire n_762;
wire n_1030;
wire n_1202;
wire n_881;
wire n_1199;
wire n_875;
wire n_465;
wire n_367;
wire n_680;
wire n_760;
wire n_741;
wire n_209;
wire n_1027;
wire n_1008;
wire n_590;
wire n_625;
wire n_661;
wire n_1189;
wire n_223;
wire n_278;
wire n_1079;
wire n_341;
wire n_362;
wire n_1212;
wire n_226;
wire n_828;
wire n_462;
wire n_208;
wire n_607;
wire n_671;
wire n_726;
wire n_1033;
wire n_316;
wire n_419;
wire n_304;
wire n_212;
wire n_700;
wire n_694;
wire n_1103;
wire n_933;
wire n_740;
wire n_1038;
wire n_578;
wire n_703;
wire n_1003;
wire n_365;
wire n_978;
wire n_1061;
wire n_384;
wire n_297;
wire n_595;
wire n_627;
wire n_1203;
wire n_524;
wire n_342;
wire n_820;
wire n_1044;
wire n_951;
wire n_783;
wire n_725;
wire n_952;
wire n_999;
wire n_358;
wire n_1217;
wire n_751;
wire n_449;
wire n_749;
wire n_1208;
wire n_798;
wire n_188;
wire n_1164;
wire n_310;
wire n_509;
wire n_186;
wire n_245;
wire n_1209;
wire n_368;
wire n_575;
wire n_994;
wire n_1072;
wire n_677;
wire n_969;
wire n_988;
wire n_805;
wire n_1151;
wire n_396;
wire n_495;
wire n_1065;
wire n_815;
wire n_350;
wire n_1100;
wire n_1214;
wire n_585;
wire n_732;
wire n_974;
wire n_568;
wire n_392;
wire n_840;
wire n_442;
wire n_480;
wire n_874;
wire n_724;
wire n_1128;
wire n_382;
wire n_673;
wire n_1020;
wire n_180;
wire n_1009;
wire n_1042;
wire n_1071;
wire n_628;
wire n_1067;
wire n_1204;
wire n_1160;
wire n_883;
wire n_557;
wire n_823;
wire n_1132;
wire n_349;
wire n_643;
wire n_233;
wire n_698;
wire n_617;
wire n_898;
wire n_1074;
wire n_1032;
wire n_845;
wire n_255;
wire n_807;
wire n_1036;
wire n_739;
wire n_284;
wire n_400;
wire n_955;
wire n_337;
wire n_865;
wire n_1138;
wire n_893;
wire n_214;
wire n_925;
wire n_1099;
wire n_1101;
wire n_485;
wire n_1026;
wire n_443;
wire n_246;
wire n_892;
wire n_768;
wire n_1097;
wire n_471;
wire n_289;
wire n_935;
wire n_1192;
wire n_421;
wire n_781;
wire n_424;
wire n_789;
wire n_615;
wire n_1130;
wire n_181;
wire n_1127;
wire n_182;
wire n_238;
wire n_1095;
wire n_573;
wire n_769;
wire n_202;
wire n_320;
wire n_639;
wire n_963;
wire n_676;
wire n_327;
wire n_794;
wire n_727;
wire n_894;
wire n_369;
wire n_1120;
wire n_597;
wire n_685;
wire n_280;
wire n_287;
wire n_832;
wire n_353;
wire n_1187;
wire n_610;
wire n_555;
wire n_389;
wire n_814;
wire n_415;
wire n_830;
wire n_605;
wire n_230;
wire n_461;
wire n_873;
wire n_383;
wire n_826;
wire n_1024;
wire n_669;
wire n_200;
wire n_447;
wire n_872;
wire n_176;
wire n_1139;
wire n_198;
wire n_300;
wire n_179;
wire n_248;
wire n_222;
wire n_718;
wire n_1018;
wire n_517;
wire n_1172;
wire n_747;
wire n_852;
wire n_667;
wire n_229;
wire n_542;
wire n_847;
wire n_644;
wire n_682;
wire n_851;
wire n_1105;
wire n_1206;
wire n_621;
wire n_305;
wire n_1037;
wire n_721;
wire n_996;
wire n_750;
wire n_532;
wire n_742;
wire n_535;
wire n_691;
wire n_250;
wire n_372;
wire n_468;
wire n_544;
wire n_901;
wire n_923;
wire n_504;
wire n_1078;
wire n_314;
wire n_1140;
wire n_378;
wire n_413;
wire n_1196;
wire n_377;
wire n_791;
wire n_183;
wire n_510;
wire n_837;
wire n_836;
wire n_1015;
wire n_863;
wire n_375;
wire n_601;
wire n_338;
wire n_522;
wire n_948;
wire n_466;
wire n_704;
wire n_918;
wire n_748;
wire n_506;
wire n_1114;
wire n_1147;
wire n_763;
wire n_1057;
wire n_360;
wire n_945;
wire n_977;
wire n_603;
wire n_1005;
wire n_991;
wire n_957;
wire n_235;
wire n_1143;
wire n_536;
wire n_895;
wire n_1126;
wire n_866;
wire n_1227;
wire n_622;
wire n_191;
wire n_340;
wire n_710;
wire n_1108;
wire n_387;
wire n_1182;
wire n_452;
wire n_658;
wire n_616;
wire n_744;
wire n_971;
wire n_946;
wire n_1119;
wire n_344;
wire n_581;
wire n_428;
wire n_785;
wire n_761;
wire n_746;
wire n_1205;
wire n_609;
wire n_765;
wire n_432;
wire n_987;
wire n_641;
wire n_822;
wire n_693;
wire n_1056;
wire n_631;
wire n_516;
wire n_720;
wire n_758;
wire n_842;
wire n_525;
wire n_1163;
wire n_1173;
wire n_1116;
wire n_1180;
wire n_611;
wire n_943;
wire n_1168;
wire n_491;
wire n_1219;
wire n_1216;
wire n_843;
wire n_772;
wire n_656;
wire n_989;
wire n_1174;
wire n_797;
wire n_666;
wire n_1016;
wire n_371;
wire n_795;
wire n_770;
wire n_940;
wire n_1221;
wire n_567;
wire n_899;
wire n_189;
wire n_738;
wire n_405;
wire n_213;
wire n_538;
wire n_1035;
wire n_294;
wire n_302;
wire n_499;
wire n_380;
wire n_838;
wire n_705;
wire n_647;
wire n_197;
wire n_1106;
wire n_886;
wire n_343;
wire n_844;
wire n_448;
wire n_953;
wire n_1017;
wire n_1004;
wire n_1094;
wire n_1176;
wire n_1190;
wire n_494;
wire n_539;
wire n_493;
wire n_397;
wire n_1022;
wire n_1083;
wire n_614;
wire n_529;
wire n_445;
wire n_425;
wire n_684;
wire n_930;
wire n_888;
wire n_1112;
wire n_454;
wire n_218;
wire n_1213;
wire n_638;
wire n_234;
wire n_1181;
wire n_910;
wire n_1211;
wire n_911;
wire n_947;
wire n_381;
wire n_486;
wire n_236;
wire n_653;
wire n_887;
wire n_1117;
wire n_1087;
wire n_752;
wire n_908;
wire n_944;
wire n_713;
wire n_648;
wire n_657;
wire n_1049;
wire n_576;
wire n_1028;
wire n_472;
wire n_270;
wire n_239;
wire n_414;
wire n_563;
wire n_782;
wire n_976;
wire n_490;
wire n_803;
wire n_290;
wire n_220;
wire n_809;
wire n_1043;
wire n_1011;
wire n_224;
wire n_926;
wire n_927;
wire n_1215;
wire n_986;
wire n_839;
wire n_734;
wire n_1088;
wire n_708;
wire n_196;
wire n_919;
wire n_1081;
wire n_402;
wire n_352;
wire n_917;
wire n_668;
wire n_478;
wire n_626;
wire n_990;
wire n_574;
wire n_800;
wire n_779;
wire n_1084;
wire n_929;
wire n_460;
wire n_1171;
wire n_1104;
wire n_907;
wire n_854;
wire n_1058;
wire n_417;
wire n_446;
wire n_498;
wire n_662;
wire n_1122;
wire n_870;
wire n_374;
wire n_659;
wire n_709;
wire n_904;
wire n_366;
wire n_1152;
wire n_777;
wire n_407;
wire n_913;
wire n_450;
wire n_808;
wire n_867;
wire n_272;
wire n_526;
wire n_1109;
wire n_921;
wire n_185;
wire n_712;
wire n_1183;
wire n_348;
wire n_711;
wire n_579;
wire n_376;
wire n_937;
wire n_390;
wire n_473;
wire n_1193;
wire n_1148;
wire n_293;
wire n_1054;
wire n_334;
wire n_559;
wire n_370;
wire n_1161;
wire n_458;
wire n_1070;
wire n_1085;
wire n_232;
wire n_650;
wire n_998;
wire n_1046;
wire n_717;
wire n_1145;
wire n_330;
wire n_771;
wire n_1121;
wire n_470;
wire n_475;
wire n_924;
wire n_1102;
wire n_298;
wire n_492;
wire n_972;
wire n_281;
wire n_258;
wire n_551;
wire n_699;
wire n_456;
wire n_1149;
wire n_564;
wire n_1178;
wire n_260;
wire n_265;
wire n_313;
wire n_451;
wire n_624;
wire n_1184;
wire n_824;
wire n_962;
wire n_1073;
wire n_1000;
wire n_279;
wire n_686;
wire n_796;
wire n_1041;
wire n_252;
wire n_757;
wire n_228;
wire n_565;
wire n_594;
wire n_719;
wire n_1195;
wire n_356;
wire n_577;
wire n_936;
wire n_184;
wire n_552;
wire n_1186;
wire n_1062;
wire n_619;
wire n_885;
wire n_455;
wire n_216;
wire n_896;
wire n_521;
wire n_363;
wire n_572;
wire n_912;
wire n_395;
wire n_813;
wire n_592;
wire n_1090;
wire n_745;
wire n_654;
wire n_323;
wire n_829;
wire n_1156;
wire n_606;
wire n_393;
wire n_818;
wire n_984;
wire n_411;
wire n_1142;
wire n_503;
wire n_716;
wire n_623;
wire n_1048;
wire n_1123;
wire n_884;
wire n_1201;
wire n_599;
wire n_1222;
wire n_513;
wire n_776;
wire n_321;
wire n_645;
wire n_331;
wire n_916;
wire n_227;
wire n_868;
wire n_570;
wire n_731;
wire n_859;
wire n_406;
wire n_735;
wire n_483;
wire n_204;
wire n_482;
wire n_934;
wire n_755;
wire n_931;
wire n_1021;
wire n_474;
wire n_527;
wire n_261;
wire n_608;
wire n_620;
wire n_420;
wire n_683;
wire n_630;
wire n_312;
wire n_394;
wire n_878;
wire n_519;
wire n_541;
wire n_512;
wire n_958;
wire n_292;
wire n_307;
wire n_469;
wire n_1137;
wire n_433;
wire n_500;
wire n_1218;
wire n_942;
wire n_792;
wire n_880;
wire n_476;
wire n_981;
wire n_714;
wire n_291;
wire n_219;
wire n_543;
wire n_1144;
wire n_889;
wire n_357;
wire n_264;
wire n_263;
wire n_985;
wire n_589;
wire n_860;
wire n_481;
wire n_1162;
wire n_1225;
wire n_788;
wire n_819;
wire n_939;
wire n_997;
wire n_821;
wire n_325;
wire n_938;
wire n_1068;
wire n_767;
wire n_804;
wire n_329;
wire n_464;
wire n_600;
wire n_831;
wire n_802;
wire n_964;
wire n_982;
wire n_561;
wire n_477;
wire n_549;
wire n_980;
wire n_533;
wire n_954;
wire n_1075;
wire n_408;
wire n_932;
wire n_806;
wire n_864;
wire n_879;
wire n_959;
wire n_1198;
wire n_237;
wire n_584;
wire n_1110;
wire n_244;
wire n_399;
wire n_243;
wire n_979;
wire n_548;
wire n_905;
wire n_282;
wire n_436;
wire n_833;
wire n_211;
wire n_523;
wire n_707;
wire n_322;
wire n_993;
wire n_345;
wire n_409;
wire n_231;
wire n_354;
wire n_689;
wire n_799;
wire n_505;
wire n_240;
wire n_1155;
wire n_756;
wire n_319;
wire n_547;
wire n_537;
wire n_273;
wire n_558;
wire n_810;
wire n_1133;
wire n_635;
wire n_787;
wire n_1194;
wire n_311;
wire n_1064;
wire n_403;
wire n_1080;
wire n_723;
wire n_253;
wire n_634;
wire n_1051;
wire n_583;
wire n_596;
wire n_966;
wire n_546;
wire n_562;
wire n_1141;
wire n_1146;
wire n_249;
wire n_386;
wire n_201;
wire n_764;
wire n_1039;
wire n_1220;
wire n_556;
wire n_1034;
wire n_1086;
wire n_1066;
wire n_692;
wire n_733;
wire n_1158;
wire n_754;
wire n_1136;
wire n_941;
wire n_975;
wire n_1031;
wire n_487;
wire n_550;
wire n_241;
wire n_1125;
wire n_275;
wire n_553;
wire n_652;
wire n_849;
wire n_970;
wire n_1107;
wire n_560;
wire n_1014;
wire n_753;
wire n_642;
wire n_995;
wire n_276;
wire n_1159;
wire n_569;
wire n_1092;
wire n_441;
wire n_221;
wire n_882;
wire n_811;
wire n_1060;
wire n_444;
wire n_586;
wire n_423;
wire n_737;
wire n_318;
wire n_1207;
wire n_1111;
wire n_303;
wire n_1223;
wire n_511;
wire n_715;
wire n_467;
wire n_306;
wire n_269;
wire n_193;
wire n_359;
wire n_973;
wire n_346;
wire n_1053;
wire n_416;
wire n_530;
wire n_277;
wire n_520;
wire n_1029;
wire n_418;
wire n_1093;
wire n_618;
wire n_1055;
wire n_790;
wire n_582;
wire n_199;
wire n_1167;
wire n_266;
wire n_296;
wire n_861;
wire n_674;
wire n_857;
wire n_871;
wire n_967;
wire n_775;
wire n_922;
wire n_571;
wire n_268;
wire n_271;
wire n_404;
wire n_651;
wire n_439;
wire n_1153;
wire n_1210;
wire n_217;
wire n_518;
wire n_299;
wire n_210;
wire n_206;
wire n_679;
wire n_1069;
wire n_1185;
wire n_453;
wire n_612;
wire n_633;
wire n_1170;
wire n_665;
wire n_902;
wire n_333;
wire n_588;
wire n_215;
wire n_178;
wire n_247;
wire n_225;
wire n_308;
wire n_309;
wire n_914;
wire n_759;
wire n_1047;
wire n_1010;
wire n_355;
wire n_1165;
wire n_426;
wire n_317;
wire n_1040;
wire n_915;
wire n_632;
wire n_702;
wire n_1166;
wire n_431;
wire n_347;
wire n_812;
wire n_459;
wire n_1131;
wire n_1052;
wire n_502;
wire n_1175;
wire n_328;
wire n_672;
wire n_534;
wire n_488;
wire n_429;
wire n_1006;
wire n_373;
wire n_1012;
wire n_497;
wire n_195;
wire n_285;
wire n_780;
wire n_773;
wire n_675;
wire n_903;
wire n_257;
wire n_920;
wire n_730;
wire n_655;
wire n_706;
wire n_1045;
wire n_786;
wire n_670;
wire n_286;
wire n_203;
wire n_1224;
wire n_254;
wire n_207;
wire n_834;
wire n_242;
wire n_835;
wire n_928;
wire n_690;
wire n_850;
wire n_1135;
wire n_1089;
wire n_1169;
wire n_1179;
wire n_401;
wire n_324;
wire n_743;
wire n_816;
wire n_766;
wire n_1157;
wire n_335;
wire n_430;
wire n_1002;
wire n_463;
wire n_1188;
wire n_545;
wire n_489;
wire n_877;
wire n_205;
wire n_604;
wire n_848;
wire n_251;
wire n_1019;
wire n_301;
wire n_274;
wire n_636;
wire n_825;
wire n_728;
wire n_681;
wire n_1096;
wire n_1063;
wire n_1226;
wire n_729;
wire n_1091;
wire n_876;
wire n_774;
wire n_412;
wire n_640;
wire n_660;
wire n_965;
wire n_267;
wire n_438;
wire n_1124;
wire n_339;
wire n_784;
wire n_315;
wire n_515;
wire n_434;
wire n_983;
wire n_288;
wire n_427;
wire n_1200;
wire n_1059;
wire n_1197;
wire n_479;
wire n_496;
wire n_598;
wire n_422;
wire n_696;
wire n_906;
wire n_688;
wire n_722;
wire n_1077;
wire n_961;
wire n_862;
wire n_869;
wire n_351;
wire n_1154;
wire n_437;
wire n_1082;
wire n_259;
wire n_177;
wire n_1113;
wire n_540;
wire n_593;
wire n_514;
wire n_646;
wire n_528;
wire n_391;
wire n_457;
wire n_1098;
wire n_697;
wire n_687;
wire n_364;
wire n_890;
wire n_637;
wire n_295;
wire n_385;
wire n_701;
wire n_817;
wire n_950;
wire n_629;
wire n_388;
wire n_190;
wire n_858;
wire n_262;
wire n_484;
wire n_613;
wire n_736;
wire n_187;
wire n_897;
wire n_900;
wire n_846;
wire n_501;
wire n_841;
wire n_956;
wire n_960;
wire n_531;
wire n_827;
wire n_1001;
wire n_508;
wire n_361;
wire n_663;
wire n_856;
wire n_1050;
wire n_379;
wire n_778;
wire n_1025;
wire n_1134;
wire n_1177;
wire n_332;
wire n_891;
wire n_336;
wire n_1150;
wire n_398;
wire n_410;
wire n_1129;
wire n_1191;
wire n_566;
wire n_554;
wire n_602;
wire n_1013;
wire n_1023;
wire n_1076;
wire n_1118;
wire n_664;
wire n_194;
wire n_949;
wire n_678;
wire n_192;
wire n_1007;
wire n_649;
wire n_855;
wire n_283;

INVx1_ASAP7_75t_L g176 ( 
.A(n_77),
.Y(n_176)
);

INVxp33_ASAP7_75t_R g177 ( 
.A(n_13),
.Y(n_177)
);

CKINVDCx20_ASAP7_75t_R g178 ( 
.A(n_84),
.Y(n_178)
);

CKINVDCx5p33_ASAP7_75t_R g179 ( 
.A(n_122),
.Y(n_179)
);

BUFx6f_ASAP7_75t_L g180 ( 
.A(n_164),
.Y(n_180)
);

CKINVDCx5p33_ASAP7_75t_R g181 ( 
.A(n_18),
.Y(n_181)
);

CKINVDCx5p33_ASAP7_75t_R g182 ( 
.A(n_70),
.Y(n_182)
);

INVx1_ASAP7_75t_SL g183 ( 
.A(n_79),
.Y(n_183)
);

CKINVDCx5p33_ASAP7_75t_R g184 ( 
.A(n_114),
.Y(n_184)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_68),
.Y(n_185)
);

CKINVDCx5p33_ASAP7_75t_R g186 ( 
.A(n_119),
.Y(n_186)
);

CKINVDCx5p33_ASAP7_75t_R g187 ( 
.A(n_92),
.Y(n_187)
);

CKINVDCx5p33_ASAP7_75t_R g188 ( 
.A(n_161),
.Y(n_188)
);

CKINVDCx5p33_ASAP7_75t_R g189 ( 
.A(n_73),
.Y(n_189)
);

CKINVDCx20_ASAP7_75t_R g190 ( 
.A(n_110),
.Y(n_190)
);

CKINVDCx5p33_ASAP7_75t_R g191 ( 
.A(n_4),
.Y(n_191)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_15),
.Y(n_192)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_6),
.Y(n_193)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_102),
.Y(n_194)
);

CKINVDCx5p33_ASAP7_75t_R g195 ( 
.A(n_26),
.Y(n_195)
);

CKINVDCx5p33_ASAP7_75t_R g196 ( 
.A(n_100),
.Y(n_196)
);

INVxp67_ASAP7_75t_L g197 ( 
.A(n_168),
.Y(n_197)
);

CKINVDCx5p33_ASAP7_75t_R g198 ( 
.A(n_160),
.Y(n_198)
);

BUFx3_ASAP7_75t_L g199 ( 
.A(n_156),
.Y(n_199)
);

CKINVDCx5p33_ASAP7_75t_R g200 ( 
.A(n_170),
.Y(n_200)
);

CKINVDCx5p33_ASAP7_75t_R g201 ( 
.A(n_32),
.Y(n_201)
);

CKINVDCx5p33_ASAP7_75t_R g202 ( 
.A(n_36),
.Y(n_202)
);

CKINVDCx5p33_ASAP7_75t_R g203 ( 
.A(n_3),
.Y(n_203)
);

INVx2_ASAP7_75t_L g204 ( 
.A(n_104),
.Y(n_204)
);

CKINVDCx5p33_ASAP7_75t_R g205 ( 
.A(n_45),
.Y(n_205)
);

CKINVDCx5p33_ASAP7_75t_R g206 ( 
.A(n_171),
.Y(n_206)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_18),
.Y(n_207)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_134),
.Y(n_208)
);

CKINVDCx5p33_ASAP7_75t_R g209 ( 
.A(n_32),
.Y(n_209)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_91),
.Y(n_210)
);

CKINVDCx20_ASAP7_75t_R g211 ( 
.A(n_155),
.Y(n_211)
);

CKINVDCx5p33_ASAP7_75t_R g212 ( 
.A(n_116),
.Y(n_212)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_106),
.Y(n_213)
);

CKINVDCx5p33_ASAP7_75t_R g214 ( 
.A(n_175),
.Y(n_214)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_19),
.Y(n_215)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_173),
.Y(n_216)
);

INVx2_ASAP7_75t_L g217 ( 
.A(n_103),
.Y(n_217)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_123),
.Y(n_218)
);

CKINVDCx20_ASAP7_75t_R g219 ( 
.A(n_17),
.Y(n_219)
);

CKINVDCx5p33_ASAP7_75t_R g220 ( 
.A(n_85),
.Y(n_220)
);

BUFx10_ASAP7_75t_L g221 ( 
.A(n_14),
.Y(n_221)
);

CKINVDCx20_ASAP7_75t_R g222 ( 
.A(n_46),
.Y(n_222)
);

CKINVDCx5p33_ASAP7_75t_R g223 ( 
.A(n_55),
.Y(n_223)
);

BUFx3_ASAP7_75t_L g224 ( 
.A(n_76),
.Y(n_224)
);

CKINVDCx5p33_ASAP7_75t_R g225 ( 
.A(n_34),
.Y(n_225)
);

CKINVDCx5p33_ASAP7_75t_R g226 ( 
.A(n_174),
.Y(n_226)
);

CKINVDCx5p33_ASAP7_75t_R g227 ( 
.A(n_152),
.Y(n_227)
);

BUFx5_ASAP7_75t_L g228 ( 
.A(n_31),
.Y(n_228)
);

CKINVDCx5p33_ASAP7_75t_R g229 ( 
.A(n_145),
.Y(n_229)
);

CKINVDCx5p33_ASAP7_75t_R g230 ( 
.A(n_20),
.Y(n_230)
);

INVxp67_ASAP7_75t_L g231 ( 
.A(n_25),
.Y(n_231)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_22),
.Y(n_232)
);

BUFx2_ASAP7_75t_L g233 ( 
.A(n_99),
.Y(n_233)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_228),
.Y(n_234)
);

CKINVDCx5p33_ASAP7_75t_R g235 ( 
.A(n_179),
.Y(n_235)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_228),
.Y(n_236)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_228),
.Y(n_237)
);

CKINVDCx5p33_ASAP7_75t_R g238 ( 
.A(n_182),
.Y(n_238)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_228),
.Y(n_239)
);

CKINVDCx5p33_ASAP7_75t_R g240 ( 
.A(n_184),
.Y(n_240)
);

CKINVDCx16_ASAP7_75t_R g241 ( 
.A(n_221),
.Y(n_241)
);

CKINVDCx5p33_ASAP7_75t_R g242 ( 
.A(n_186),
.Y(n_242)
);

CKINVDCx5p33_ASAP7_75t_R g243 ( 
.A(n_187),
.Y(n_243)
);

BUFx8_ASAP7_75t_SL g244 ( 
.A(n_219),
.Y(n_244)
);

BUFx2_ASAP7_75t_L g245 ( 
.A(n_181),
.Y(n_245)
);

CKINVDCx5p33_ASAP7_75t_R g246 ( 
.A(n_188),
.Y(n_246)
);

CKINVDCx5p33_ASAP7_75t_R g247 ( 
.A(n_189),
.Y(n_247)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_228),
.Y(n_248)
);

CKINVDCx5p33_ASAP7_75t_R g249 ( 
.A(n_196),
.Y(n_249)
);

INVx2_ASAP7_75t_L g250 ( 
.A(n_228),
.Y(n_250)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_228),
.Y(n_251)
);

CKINVDCx5p33_ASAP7_75t_R g252 ( 
.A(n_198),
.Y(n_252)
);

HB1xp67_ASAP7_75t_L g253 ( 
.A(n_181),
.Y(n_253)
);

CKINVDCx5p33_ASAP7_75t_R g254 ( 
.A(n_200),
.Y(n_254)
);

CKINVDCx14_ASAP7_75t_R g255 ( 
.A(n_233),
.Y(n_255)
);

CKINVDCx5p33_ASAP7_75t_R g256 ( 
.A(n_205),
.Y(n_256)
);

CKINVDCx5p33_ASAP7_75t_R g257 ( 
.A(n_206),
.Y(n_257)
);

CKINVDCx5p33_ASAP7_75t_R g258 ( 
.A(n_212),
.Y(n_258)
);

CKINVDCx5p33_ASAP7_75t_R g259 ( 
.A(n_214),
.Y(n_259)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_232),
.Y(n_260)
);

BUFx3_ASAP7_75t_L g261 ( 
.A(n_199),
.Y(n_261)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_192),
.Y(n_262)
);

CKINVDCx5p33_ASAP7_75t_R g263 ( 
.A(n_220),
.Y(n_263)
);

CKINVDCx5p33_ASAP7_75t_R g264 ( 
.A(n_235),
.Y(n_264)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_234),
.Y(n_265)
);

CKINVDCx5p33_ASAP7_75t_R g266 ( 
.A(n_238),
.Y(n_266)
);

CKINVDCx5p33_ASAP7_75t_R g267 ( 
.A(n_240),
.Y(n_267)
);

CKINVDCx5p33_ASAP7_75t_R g268 ( 
.A(n_242),
.Y(n_268)
);

CKINVDCx20_ASAP7_75t_R g269 ( 
.A(n_244),
.Y(n_269)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_234),
.Y(n_270)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_236),
.Y(n_271)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_236),
.Y(n_272)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_237),
.Y(n_273)
);

INVx2_ASAP7_75t_L g274 ( 
.A(n_250),
.Y(n_274)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_237),
.Y(n_275)
);

BUFx6f_ASAP7_75t_L g276 ( 
.A(n_250),
.Y(n_276)
);

BUFx3_ASAP7_75t_L g277 ( 
.A(n_261),
.Y(n_277)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_239),
.Y(n_278)
);

CKINVDCx5p33_ASAP7_75t_R g279 ( 
.A(n_243),
.Y(n_279)
);

INVx1_ASAP7_75t_SL g280 ( 
.A(n_244),
.Y(n_280)
);

CKINVDCx5p33_ASAP7_75t_R g281 ( 
.A(n_246),
.Y(n_281)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_239),
.Y(n_282)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_248),
.Y(n_283)
);

BUFx6f_ASAP7_75t_L g284 ( 
.A(n_250),
.Y(n_284)
);

CKINVDCx20_ASAP7_75t_R g285 ( 
.A(n_241),
.Y(n_285)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_248),
.Y(n_286)
);

CKINVDCx5p33_ASAP7_75t_R g287 ( 
.A(n_247),
.Y(n_287)
);

BUFx10_ASAP7_75t_L g288 ( 
.A(n_249),
.Y(n_288)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_251),
.Y(n_289)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_251),
.Y(n_290)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_260),
.Y(n_291)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_260),
.Y(n_292)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_262),
.Y(n_293)
);

CKINVDCx16_ASAP7_75t_R g294 ( 
.A(n_241),
.Y(n_294)
);

CKINVDCx5p33_ASAP7_75t_R g295 ( 
.A(n_252),
.Y(n_295)
);

NOR2xp67_ASAP7_75t_L g296 ( 
.A(n_263),
.B(n_197),
.Y(n_296)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_262),
.Y(n_297)
);

CKINVDCx5p33_ASAP7_75t_R g298 ( 
.A(n_254),
.Y(n_298)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_261),
.Y(n_299)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_261),
.Y(n_300)
);

CKINVDCx20_ASAP7_75t_R g301 ( 
.A(n_255),
.Y(n_301)
);

CKINVDCx16_ASAP7_75t_R g302 ( 
.A(n_255),
.Y(n_302)
);

CKINVDCx20_ASAP7_75t_R g303 ( 
.A(n_245),
.Y(n_303)
);

CKINVDCx20_ASAP7_75t_R g304 ( 
.A(n_245),
.Y(n_304)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_256),
.Y(n_305)
);

CKINVDCx5p33_ASAP7_75t_R g306 ( 
.A(n_257),
.Y(n_306)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_258),
.Y(n_307)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_259),
.Y(n_308)
);

CKINVDCx5p33_ASAP7_75t_R g309 ( 
.A(n_253),
.Y(n_309)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_253),
.Y(n_310)
);

CKINVDCx5p33_ASAP7_75t_R g311 ( 
.A(n_235),
.Y(n_311)
);

INVx2_ASAP7_75t_L g312 ( 
.A(n_250),
.Y(n_312)
);

INVxp67_ASAP7_75t_L g313 ( 
.A(n_253),
.Y(n_313)
);

CKINVDCx20_ASAP7_75t_R g314 ( 
.A(n_244),
.Y(n_314)
);

CKINVDCx5p33_ASAP7_75t_R g315 ( 
.A(n_235),
.Y(n_315)
);

INVxp67_ASAP7_75t_SL g316 ( 
.A(n_276),
.Y(n_316)
);

INVxp67_ASAP7_75t_SL g317 ( 
.A(n_276),
.Y(n_317)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_265),
.Y(n_318)
);

INVx2_ASAP7_75t_L g319 ( 
.A(n_274),
.Y(n_319)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_270),
.Y(n_320)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_271),
.Y(n_321)
);

CKINVDCx5p33_ASAP7_75t_R g322 ( 
.A(n_266),
.Y(n_322)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_272),
.Y(n_323)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_273),
.Y(n_324)
);

CKINVDCx5p33_ASAP7_75t_R g325 ( 
.A(n_267),
.Y(n_325)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_275),
.Y(n_326)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_278),
.Y(n_327)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_282),
.Y(n_328)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_283),
.Y(n_329)
);

CKINVDCx5p33_ASAP7_75t_R g330 ( 
.A(n_268),
.Y(n_330)
);

CKINVDCx20_ASAP7_75t_R g331 ( 
.A(n_301),
.Y(n_331)
);

INVxp33_ASAP7_75t_SL g332 ( 
.A(n_264),
.Y(n_332)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_286),
.Y(n_333)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_289),
.Y(n_334)
);

INVx1_ASAP7_75t_SL g335 ( 
.A(n_303),
.Y(n_335)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_290),
.Y(n_336)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_291),
.Y(n_337)
);

INVx2_ASAP7_75t_L g338 ( 
.A(n_312),
.Y(n_338)
);

INVxp33_ASAP7_75t_SL g339 ( 
.A(n_264),
.Y(n_339)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_312),
.Y(n_340)
);

CKINVDCx5p33_ASAP7_75t_R g341 ( 
.A(n_279),
.Y(n_341)
);

CKINVDCx5p33_ASAP7_75t_R g342 ( 
.A(n_281),
.Y(n_342)
);

INVxp67_ASAP7_75t_SL g343 ( 
.A(n_276),
.Y(n_343)
);

INVx1_ASAP7_75t_L g344 ( 
.A(n_276),
.Y(n_344)
);

INVx1_ASAP7_75t_L g345 ( 
.A(n_292),
.Y(n_345)
);

CKINVDCx5p33_ASAP7_75t_R g346 ( 
.A(n_287),
.Y(n_346)
);

INVxp67_ASAP7_75t_SL g347 ( 
.A(n_284),
.Y(n_347)
);

INVx1_ASAP7_75t_L g348 ( 
.A(n_284),
.Y(n_348)
);

INVx1_ASAP7_75t_L g349 ( 
.A(n_284),
.Y(n_349)
);

INVxp67_ASAP7_75t_L g350 ( 
.A(n_310),
.Y(n_350)
);

INVxp33_ASAP7_75t_L g351 ( 
.A(n_299),
.Y(n_351)
);

INVx1_ASAP7_75t_L g352 ( 
.A(n_284),
.Y(n_352)
);

INVx1_ASAP7_75t_L g353 ( 
.A(n_293),
.Y(n_353)
);

CKINVDCx5p33_ASAP7_75t_R g354 ( 
.A(n_295),
.Y(n_354)
);

CKINVDCx20_ASAP7_75t_R g355 ( 
.A(n_301),
.Y(n_355)
);

INVx1_ASAP7_75t_L g356 ( 
.A(n_297),
.Y(n_356)
);

INVxp33_ASAP7_75t_L g357 ( 
.A(n_300),
.Y(n_357)
);

CKINVDCx16_ASAP7_75t_R g358 ( 
.A(n_302),
.Y(n_358)
);

INVx1_ASAP7_75t_L g359 ( 
.A(n_277),
.Y(n_359)
);

CKINVDCx5p33_ASAP7_75t_R g360 ( 
.A(n_298),
.Y(n_360)
);

CKINVDCx5p33_ASAP7_75t_R g361 ( 
.A(n_306),
.Y(n_361)
);

INVx1_ASAP7_75t_L g362 ( 
.A(n_277),
.Y(n_362)
);

INVx1_ASAP7_75t_L g363 ( 
.A(n_305),
.Y(n_363)
);

BUFx3_ASAP7_75t_L g364 ( 
.A(n_307),
.Y(n_364)
);

CKINVDCx5p33_ASAP7_75t_R g365 ( 
.A(n_322),
.Y(n_365)
);

CKINVDCx20_ASAP7_75t_R g366 ( 
.A(n_331),
.Y(n_366)
);

CKINVDCx16_ASAP7_75t_R g367 ( 
.A(n_358),
.Y(n_367)
);

INVx1_ASAP7_75t_L g368 ( 
.A(n_353),
.Y(n_368)
);

INVxp67_ASAP7_75t_SL g369 ( 
.A(n_344),
.Y(n_369)
);

CKINVDCx16_ASAP7_75t_R g370 ( 
.A(n_355),
.Y(n_370)
);

INVx1_ASAP7_75t_L g371 ( 
.A(n_353),
.Y(n_371)
);

INVx1_ASAP7_75t_L g372 ( 
.A(n_356),
.Y(n_372)
);

NOR2xp67_ASAP7_75t_L g373 ( 
.A(n_325),
.B(n_311),
.Y(n_373)
);

INVx1_ASAP7_75t_L g374 ( 
.A(n_356),
.Y(n_374)
);

INVx1_ASAP7_75t_L g375 ( 
.A(n_337),
.Y(n_375)
);

CKINVDCx5p33_ASAP7_75t_R g376 ( 
.A(n_330),
.Y(n_376)
);

INVx2_ASAP7_75t_L g377 ( 
.A(n_319),
.Y(n_377)
);

CKINVDCx20_ASAP7_75t_R g378 ( 
.A(n_335),
.Y(n_378)
);

INVx1_ASAP7_75t_L g379 ( 
.A(n_345),
.Y(n_379)
);

CKINVDCx20_ASAP7_75t_R g380 ( 
.A(n_341),
.Y(n_380)
);

INVx1_ASAP7_75t_L g381 ( 
.A(n_318),
.Y(n_381)
);

INVx1_ASAP7_75t_L g382 ( 
.A(n_318),
.Y(n_382)
);

INVxp67_ASAP7_75t_L g383 ( 
.A(n_363),
.Y(n_383)
);

INVxp33_ASAP7_75t_SL g384 ( 
.A(n_342),
.Y(n_384)
);

INVx1_ASAP7_75t_L g385 ( 
.A(n_320),
.Y(n_385)
);

INVx1_ASAP7_75t_L g386 ( 
.A(n_320),
.Y(n_386)
);

INVx1_ASAP7_75t_L g387 ( 
.A(n_321),
.Y(n_387)
);

INVx1_ASAP7_75t_L g388 ( 
.A(n_321),
.Y(n_388)
);

CKINVDCx5p33_ASAP7_75t_R g389 ( 
.A(n_346),
.Y(n_389)
);

CKINVDCx20_ASAP7_75t_R g390 ( 
.A(n_354),
.Y(n_390)
);

INVx1_ASAP7_75t_L g391 ( 
.A(n_323),
.Y(n_391)
);

INVx1_ASAP7_75t_L g392 ( 
.A(n_323),
.Y(n_392)
);

INVx1_ASAP7_75t_L g393 ( 
.A(n_324),
.Y(n_393)
);

INVx1_ASAP7_75t_L g394 ( 
.A(n_324),
.Y(n_394)
);

INVx1_ASAP7_75t_L g395 ( 
.A(n_326),
.Y(n_395)
);

CKINVDCx20_ASAP7_75t_R g396 ( 
.A(n_360),
.Y(n_396)
);

INVx1_ASAP7_75t_L g397 ( 
.A(n_326),
.Y(n_397)
);

CKINVDCx20_ASAP7_75t_R g398 ( 
.A(n_361),
.Y(n_398)
);

CKINVDCx20_ASAP7_75t_R g399 ( 
.A(n_364),
.Y(n_399)
);

CKINVDCx20_ASAP7_75t_R g400 ( 
.A(n_364),
.Y(n_400)
);

CKINVDCx20_ASAP7_75t_R g401 ( 
.A(n_350),
.Y(n_401)
);

INVx1_ASAP7_75t_L g402 ( 
.A(n_327),
.Y(n_402)
);

CKINVDCx5p33_ASAP7_75t_R g403 ( 
.A(n_332),
.Y(n_403)
);

INVxp67_ASAP7_75t_SL g404 ( 
.A(n_344),
.Y(n_404)
);

NOR2xp67_ASAP7_75t_L g405 ( 
.A(n_363),
.B(n_311),
.Y(n_405)
);

INVxp33_ASAP7_75t_L g406 ( 
.A(n_351),
.Y(n_406)
);

CKINVDCx5p33_ASAP7_75t_R g407 ( 
.A(n_339),
.Y(n_407)
);

CKINVDCx5p33_ASAP7_75t_R g408 ( 
.A(n_359),
.Y(n_408)
);

CKINVDCx20_ASAP7_75t_R g409 ( 
.A(n_359),
.Y(n_409)
);

INVx1_ASAP7_75t_L g410 ( 
.A(n_377),
.Y(n_410)
);

BUFx6f_ASAP7_75t_L g411 ( 
.A(n_368),
.Y(n_411)
);

OAI22xp5_ASAP7_75t_L g412 ( 
.A1(n_383),
.A2(n_371),
.B1(n_374),
.B2(n_372),
.Y(n_412)
);

INVx2_ASAP7_75t_L g413 ( 
.A(n_381),
.Y(n_413)
);

NAND2xp5_ASAP7_75t_L g414 ( 
.A(n_382),
.B(n_328),
.Y(n_414)
);

INVx1_ASAP7_75t_L g415 ( 
.A(n_385),
.Y(n_415)
);

INVx2_ASAP7_75t_L g416 ( 
.A(n_386),
.Y(n_416)
);

NAND2xp5_ASAP7_75t_L g417 ( 
.A(n_387),
.B(n_328),
.Y(n_417)
);

INVx2_ASAP7_75t_L g418 ( 
.A(n_388),
.Y(n_418)
);

BUFx3_ASAP7_75t_L g419 ( 
.A(n_380),
.Y(n_419)
);

INVx3_ASAP7_75t_L g420 ( 
.A(n_391),
.Y(n_420)
);

CKINVDCx11_ASAP7_75t_R g421 ( 
.A(n_366),
.Y(n_421)
);

INVx1_ASAP7_75t_L g422 ( 
.A(n_392),
.Y(n_422)
);

OAI22xp5_ASAP7_75t_L g423 ( 
.A1(n_393),
.A2(n_333),
.B1(n_334),
.B2(n_329),
.Y(n_423)
);

OAI22x1_ASAP7_75t_L g424 ( 
.A1(n_408),
.A2(n_309),
.B1(n_313),
.B2(n_280),
.Y(n_424)
);

INVx2_ASAP7_75t_L g425 ( 
.A(n_394),
.Y(n_425)
);

CKINVDCx5p33_ASAP7_75t_R g426 ( 
.A(n_365),
.Y(n_426)
);

INVx2_ASAP7_75t_L g427 ( 
.A(n_395),
.Y(n_427)
);

INVx2_ASAP7_75t_L g428 ( 
.A(n_397),
.Y(n_428)
);

INVx1_ASAP7_75t_L g429 ( 
.A(n_402),
.Y(n_429)
);

INVx1_ASAP7_75t_L g430 ( 
.A(n_375),
.Y(n_430)
);

INVx2_ASAP7_75t_L g431 ( 
.A(n_379),
.Y(n_431)
);

AND2x4_ASAP7_75t_L g432 ( 
.A(n_405),
.B(n_362),
.Y(n_432)
);

INVx1_ASAP7_75t_L g433 ( 
.A(n_369),
.Y(n_433)
);

NOR2x1_ASAP7_75t_L g434 ( 
.A(n_373),
.B(n_308),
.Y(n_434)
);

INVx3_ASAP7_75t_L g435 ( 
.A(n_404),
.Y(n_435)
);

AOI22x1_ASAP7_75t_SL g436 ( 
.A1(n_380),
.A2(n_269),
.B1(n_314),
.B2(n_219),
.Y(n_436)
);

BUFx6f_ASAP7_75t_L g437 ( 
.A(n_376),
.Y(n_437)
);

INVx2_ASAP7_75t_L g438 ( 
.A(n_409),
.Y(n_438)
);

CKINVDCx5p33_ASAP7_75t_R g439 ( 
.A(n_389),
.Y(n_439)
);

AND2x2_ASAP7_75t_L g440 ( 
.A(n_406),
.B(n_362),
.Y(n_440)
);

NAND2xp5_ASAP7_75t_L g441 ( 
.A(n_409),
.B(n_329),
.Y(n_441)
);

AND2x4_ASAP7_75t_L g442 ( 
.A(n_399),
.B(n_333),
.Y(n_442)
);

INVx1_ASAP7_75t_L g443 ( 
.A(n_399),
.Y(n_443)
);

INVx2_ASAP7_75t_L g444 ( 
.A(n_401),
.Y(n_444)
);

NAND2xp5_ASAP7_75t_L g445 ( 
.A(n_384),
.B(n_334),
.Y(n_445)
);

INVx3_ASAP7_75t_L g446 ( 
.A(n_367),
.Y(n_446)
);

BUFx12f_ASAP7_75t_L g447 ( 
.A(n_403),
.Y(n_447)
);

AND2x4_ASAP7_75t_L g448 ( 
.A(n_400),
.B(n_336),
.Y(n_448)
);

OA21x2_ASAP7_75t_L g449 ( 
.A1(n_407),
.A2(n_349),
.B(n_348),
.Y(n_449)
);

AND2x2_ASAP7_75t_L g450 ( 
.A(n_400),
.B(n_309),
.Y(n_450)
);

INVx2_ASAP7_75t_L g451 ( 
.A(n_401),
.Y(n_451)
);

INVx1_ASAP7_75t_L g452 ( 
.A(n_378),
.Y(n_452)
);

INVx6_ASAP7_75t_L g453 ( 
.A(n_370),
.Y(n_453)
);

INVx1_ASAP7_75t_L g454 ( 
.A(n_378),
.Y(n_454)
);

INVx2_ASAP7_75t_L g455 ( 
.A(n_390),
.Y(n_455)
);

HB1xp67_ASAP7_75t_L g456 ( 
.A(n_366),
.Y(n_456)
);

INVx2_ASAP7_75t_L g457 ( 
.A(n_390),
.Y(n_457)
);

INVx2_ASAP7_75t_L g458 ( 
.A(n_396),
.Y(n_458)
);

BUFx2_ASAP7_75t_L g459 ( 
.A(n_396),
.Y(n_459)
);

BUFx6f_ASAP7_75t_L g460 ( 
.A(n_398),
.Y(n_460)
);

BUFx6f_ASAP7_75t_L g461 ( 
.A(n_398),
.Y(n_461)
);

BUFx3_ASAP7_75t_L g462 ( 
.A(n_380),
.Y(n_462)
);

INVx4_ASAP7_75t_L g463 ( 
.A(n_377),
.Y(n_463)
);

BUFx2_ASAP7_75t_L g464 ( 
.A(n_399),
.Y(n_464)
);

INVx1_ASAP7_75t_L g465 ( 
.A(n_368),
.Y(n_465)
);

INVx1_ASAP7_75t_L g466 ( 
.A(n_368),
.Y(n_466)
);

OAI22xp5_ASAP7_75t_SL g467 ( 
.A1(n_366),
.A2(n_314),
.B1(n_269),
.B2(n_285),
.Y(n_467)
);

HB1xp67_ASAP7_75t_L g468 ( 
.A(n_409),
.Y(n_468)
);

CKINVDCx8_ASAP7_75t_R g469 ( 
.A(n_367),
.Y(n_469)
);

OAI21x1_ASAP7_75t_L g470 ( 
.A1(n_377),
.A2(n_349),
.B(n_348),
.Y(n_470)
);

AND2x4_ASAP7_75t_L g471 ( 
.A(n_375),
.B(n_336),
.Y(n_471)
);

BUFx6f_ASAP7_75t_L g472 ( 
.A(n_368),
.Y(n_472)
);

AND2x2_ASAP7_75t_L g473 ( 
.A(n_383),
.B(n_357),
.Y(n_473)
);

CKINVDCx20_ASAP7_75t_R g474 ( 
.A(n_366),
.Y(n_474)
);

BUFx3_ASAP7_75t_L g475 ( 
.A(n_380),
.Y(n_475)
);

AND2x2_ASAP7_75t_L g476 ( 
.A(n_383),
.B(n_288),
.Y(n_476)
);

INVx2_ASAP7_75t_L g477 ( 
.A(n_377),
.Y(n_477)
);

NAND2xp5_ASAP7_75t_L g478 ( 
.A(n_383),
.B(n_296),
.Y(n_478)
);

INVx2_ASAP7_75t_SL g479 ( 
.A(n_408),
.Y(n_479)
);

AOI22xp5_ASAP7_75t_L g480 ( 
.A1(n_383),
.A2(n_315),
.B1(n_352),
.B2(n_222),
.Y(n_480)
);

BUFx6f_ASAP7_75t_L g481 ( 
.A(n_368),
.Y(n_481)
);

INVx2_ASAP7_75t_L g482 ( 
.A(n_377),
.Y(n_482)
);

BUFx6f_ASAP7_75t_L g483 ( 
.A(n_368),
.Y(n_483)
);

BUFx6f_ASAP7_75t_L g484 ( 
.A(n_368),
.Y(n_484)
);

BUFx6f_ASAP7_75t_L g485 ( 
.A(n_368),
.Y(n_485)
);

AND2x4_ASAP7_75t_L g486 ( 
.A(n_375),
.B(n_352),
.Y(n_486)
);

NAND2xp5_ASAP7_75t_L g487 ( 
.A(n_383),
.B(n_315),
.Y(n_487)
);

NOR2xp33_ASAP7_75t_L g488 ( 
.A(n_406),
.B(n_303),
.Y(n_488)
);

AND2x4_ASAP7_75t_L g489 ( 
.A(n_375),
.B(n_347),
.Y(n_489)
);

BUFx6f_ASAP7_75t_L g490 ( 
.A(n_368),
.Y(n_490)
);

NAND2xp5_ASAP7_75t_L g491 ( 
.A(n_383),
.B(n_316),
.Y(n_491)
);

INVx1_ASAP7_75t_L g492 ( 
.A(n_377),
.Y(n_492)
);

NAND2xp5_ASAP7_75t_SL g493 ( 
.A(n_405),
.B(n_288),
.Y(n_493)
);

BUFx2_ASAP7_75t_L g494 ( 
.A(n_399),
.Y(n_494)
);

NAND2xp5_ASAP7_75t_L g495 ( 
.A(n_435),
.B(n_288),
.Y(n_495)
);

AND2x4_ASAP7_75t_L g496 ( 
.A(n_471),
.B(n_317),
.Y(n_496)
);

AND2x2_ASAP7_75t_L g497 ( 
.A(n_413),
.B(n_294),
.Y(n_497)
);

INVx1_ASAP7_75t_L g498 ( 
.A(n_410),
.Y(n_498)
);

INVx3_ASAP7_75t_L g499 ( 
.A(n_463),
.Y(n_499)
);

INVx2_ASAP7_75t_L g500 ( 
.A(n_477),
.Y(n_500)
);

INVx2_ASAP7_75t_L g501 ( 
.A(n_477),
.Y(n_501)
);

BUFx6f_ASAP7_75t_L g502 ( 
.A(n_411),
.Y(n_502)
);

BUFx8_ASAP7_75t_L g503 ( 
.A(n_437),
.Y(n_503)
);

BUFx6f_ASAP7_75t_L g504 ( 
.A(n_411),
.Y(n_504)
);

INVx2_ASAP7_75t_L g505 ( 
.A(n_482),
.Y(n_505)
);

NAND2xp5_ASAP7_75t_L g506 ( 
.A(n_435),
.B(n_340),
.Y(n_506)
);

CKINVDCx5p33_ASAP7_75t_R g507 ( 
.A(n_426),
.Y(n_507)
);

INVx3_ASAP7_75t_L g508 ( 
.A(n_463),
.Y(n_508)
);

AND2x4_ASAP7_75t_L g509 ( 
.A(n_471),
.B(n_413),
.Y(n_509)
);

OAI22xp5_ASAP7_75t_SL g510 ( 
.A1(n_467),
.A2(n_304),
.B1(n_285),
.B2(n_178),
.Y(n_510)
);

AND2x4_ASAP7_75t_L g511 ( 
.A(n_471),
.B(n_343),
.Y(n_511)
);

AND2x2_ASAP7_75t_L g512 ( 
.A(n_416),
.B(n_418),
.Y(n_512)
);

INVx1_ASAP7_75t_L g513 ( 
.A(n_492),
.Y(n_513)
);

NAND2xp5_ASAP7_75t_SL g514 ( 
.A(n_445),
.B(n_178),
.Y(n_514)
);

OR2x2_ASAP7_75t_L g515 ( 
.A(n_452),
.B(n_304),
.Y(n_515)
);

INVxp67_ASAP7_75t_L g516 ( 
.A(n_441),
.Y(n_516)
);

INVx1_ASAP7_75t_L g517 ( 
.A(n_492),
.Y(n_517)
);

AND3x2_ASAP7_75t_L g518 ( 
.A(n_459),
.B(n_231),
.C(n_177),
.Y(n_518)
);

HB1xp67_ASAP7_75t_L g519 ( 
.A(n_442),
.Y(n_519)
);

NOR2xp33_ASAP7_75t_L g520 ( 
.A(n_487),
.B(n_190),
.Y(n_520)
);

BUFx6f_ASAP7_75t_L g521 ( 
.A(n_411),
.Y(n_521)
);

AND2x2_ASAP7_75t_L g522 ( 
.A(n_416),
.B(n_418),
.Y(n_522)
);

INVxp67_ASAP7_75t_L g523 ( 
.A(n_440),
.Y(n_523)
);

NOR2xp33_ASAP7_75t_L g524 ( 
.A(n_479),
.B(n_190),
.Y(n_524)
);

AND2x4_ASAP7_75t_L g525 ( 
.A(n_425),
.B(n_427),
.Y(n_525)
);

BUFx2_ASAP7_75t_L g526 ( 
.A(n_442),
.Y(n_526)
);

BUFx3_ASAP7_75t_L g527 ( 
.A(n_437),
.Y(n_527)
);

INVx2_ASAP7_75t_L g528 ( 
.A(n_470),
.Y(n_528)
);

HB1xp67_ASAP7_75t_L g529 ( 
.A(n_442),
.Y(n_529)
);

AND2x2_ASAP7_75t_L g530 ( 
.A(n_427),
.B(n_428),
.Y(n_530)
);

NOR2xp33_ASAP7_75t_SL g531 ( 
.A(n_426),
.B(n_211),
.Y(n_531)
);

INVx3_ASAP7_75t_L g532 ( 
.A(n_472),
.Y(n_532)
);

OAI22xp33_ASAP7_75t_L g533 ( 
.A1(n_531),
.A2(n_480),
.B1(n_479),
.B2(n_431),
.Y(n_533)
);

OR2x2_ASAP7_75t_L g534 ( 
.A(n_515),
.B(n_444),
.Y(n_534)
);

AND2x2_ASAP7_75t_L g535 ( 
.A(n_526),
.B(n_473),
.Y(n_535)
);

AND2x2_ASAP7_75t_L g536 ( 
.A(n_526),
.B(n_473),
.Y(n_536)
);

AND2x2_ASAP7_75t_L g537 ( 
.A(n_516),
.B(n_440),
.Y(n_537)
);

INVx2_ASAP7_75t_L g538 ( 
.A(n_500),
.Y(n_538)
);

AND2x2_ASAP7_75t_L g539 ( 
.A(n_519),
.B(n_450),
.Y(n_539)
);

AOI22xp5_ASAP7_75t_L g540 ( 
.A1(n_520),
.A2(n_488),
.B1(n_450),
.B2(n_439),
.Y(n_540)
);

INVxp33_ASAP7_75t_L g541 ( 
.A(n_524),
.Y(n_541)
);

AND2x2_ASAP7_75t_L g542 ( 
.A(n_529),
.B(n_448),
.Y(n_542)
);

AOI22xp5_ASAP7_75t_L g543 ( 
.A1(n_514),
.A2(n_439),
.B1(n_476),
.B2(n_443),
.Y(n_543)
);

AND2x2_ASAP7_75t_L g544 ( 
.A(n_497),
.B(n_448),
.Y(n_544)
);

OAI22xp5_ASAP7_75t_SL g545 ( 
.A1(n_510),
.A2(n_474),
.B1(n_457),
.B2(n_458),
.Y(n_545)
);

AOI22xp5_ASAP7_75t_L g546 ( 
.A1(n_497),
.A2(n_476),
.B1(n_444),
.B2(n_451),
.Y(n_546)
);

OR2x6_ASAP7_75t_L g547 ( 
.A(n_527),
.B(n_437),
.Y(n_547)
);

AOI22xp5_ASAP7_75t_L g548 ( 
.A1(n_510),
.A2(n_451),
.B1(n_448),
.B2(n_454),
.Y(n_548)
);

BUFx10_ASAP7_75t_L g549 ( 
.A(n_507),
.Y(n_549)
);

OAI22xp33_ASAP7_75t_L g550 ( 
.A1(n_523),
.A2(n_431),
.B1(n_428),
.B2(n_414),
.Y(n_550)
);

INVx1_ASAP7_75t_L g551 ( 
.A(n_512),
.Y(n_551)
);

OAI22xp33_ASAP7_75t_L g552 ( 
.A1(n_495),
.A2(n_417),
.B1(n_422),
.B2(n_415),
.Y(n_552)
);

OAI22xp5_ASAP7_75t_SL g553 ( 
.A1(n_515),
.A2(n_474),
.B1(n_455),
.B2(n_458),
.Y(n_553)
);

AOI22xp5_ASAP7_75t_L g554 ( 
.A1(n_509),
.A2(n_455),
.B1(n_457),
.B2(n_437),
.Y(n_554)
);

AND2x2_ASAP7_75t_L g555 ( 
.A(n_509),
.B(n_438),
.Y(n_555)
);

AOI22xp5_ASAP7_75t_L g556 ( 
.A1(n_509),
.A2(n_437),
.B1(n_446),
.B2(n_438),
.Y(n_556)
);

AND2x2_ASAP7_75t_L g557 ( 
.A(n_509),
.B(n_464),
.Y(n_557)
);

INVx2_ASAP7_75t_L g558 ( 
.A(n_500),
.Y(n_558)
);

NOR2xp33_ASAP7_75t_L g559 ( 
.A(n_525),
.B(n_468),
.Y(n_559)
);

INVx1_ASAP7_75t_L g560 ( 
.A(n_512),
.Y(n_560)
);

AND2x2_ASAP7_75t_L g561 ( 
.A(n_527),
.B(n_464),
.Y(n_561)
);

OAI22xp33_ASAP7_75t_L g562 ( 
.A1(n_527),
.A2(n_429),
.B1(n_466),
.B2(n_465),
.Y(n_562)
);

INVx2_ASAP7_75t_L g563 ( 
.A(n_501),
.Y(n_563)
);

INVx2_ASAP7_75t_L g564 ( 
.A(n_501),
.Y(n_564)
);

AO22x2_ASAP7_75t_L g565 ( 
.A1(n_528),
.A2(n_412),
.B1(n_436),
.B2(n_433),
.Y(n_565)
);

AO22x2_ASAP7_75t_L g566 ( 
.A1(n_528),
.A2(n_436),
.B1(n_433),
.B2(n_423),
.Y(n_566)
);

INVx2_ASAP7_75t_L g567 ( 
.A(n_505),
.Y(n_567)
);

OR2x2_ASAP7_75t_L g568 ( 
.A(n_522),
.B(n_494),
.Y(n_568)
);

INVx2_ASAP7_75t_SL g569 ( 
.A(n_503),
.Y(n_569)
);

OAI22xp33_ASAP7_75t_L g570 ( 
.A1(n_499),
.A2(n_430),
.B1(n_481),
.B2(n_472),
.Y(n_570)
);

CKINVDCx5p33_ASAP7_75t_R g571 ( 
.A(n_503),
.Y(n_571)
);

BUFx10_ASAP7_75t_L g572 ( 
.A(n_496),
.Y(n_572)
);

AO22x2_ASAP7_75t_L g573 ( 
.A1(n_528),
.A2(n_446),
.B1(n_420),
.B2(n_493),
.Y(n_573)
);

NAND2xp5_ASAP7_75t_SL g574 ( 
.A(n_552),
.B(n_499),
.Y(n_574)
);

INVx1_ASAP7_75t_L g575 ( 
.A(n_538),
.Y(n_575)
);

NAND2xp5_ASAP7_75t_SL g576 ( 
.A(n_552),
.B(n_570),
.Y(n_576)
);

OAI22xp5_ASAP7_75t_L g577 ( 
.A1(n_540),
.A2(n_469),
.B1(n_453),
.B2(n_494),
.Y(n_577)
);

CKINVDCx5p33_ASAP7_75t_R g578 ( 
.A(n_549),
.Y(n_578)
);

NAND2xp5_ASAP7_75t_L g579 ( 
.A(n_537),
.B(n_522),
.Y(n_579)
);

NAND2xp5_ASAP7_75t_L g580 ( 
.A(n_535),
.B(n_530),
.Y(n_580)
);

INVx1_ASAP7_75t_L g581 ( 
.A(n_538),
.Y(n_581)
);

NAND2xp5_ASAP7_75t_SL g582 ( 
.A(n_570),
.B(n_499),
.Y(n_582)
);

INVx1_ASAP7_75t_L g583 ( 
.A(n_558),
.Y(n_583)
);

BUFx3_ASAP7_75t_L g584 ( 
.A(n_547),
.Y(n_584)
);

INVx2_ASAP7_75t_L g585 ( 
.A(n_558),
.Y(n_585)
);

INVx3_ASAP7_75t_L g586 ( 
.A(n_572),
.Y(n_586)
);

AO21x2_ASAP7_75t_L g587 ( 
.A1(n_550),
.A2(n_470),
.B(n_506),
.Y(n_587)
);

INVx4_ASAP7_75t_L g588 ( 
.A(n_547),
.Y(n_588)
);

NAND2xp5_ASAP7_75t_L g589 ( 
.A(n_536),
.B(n_530),
.Y(n_589)
);

CKINVDCx5p33_ASAP7_75t_R g590 ( 
.A(n_549),
.Y(n_590)
);

BUFx8_ASAP7_75t_SL g591 ( 
.A(n_571),
.Y(n_591)
);

INVx1_ASAP7_75t_L g592 ( 
.A(n_563),
.Y(n_592)
);

NAND2xp5_ASAP7_75t_L g593 ( 
.A(n_544),
.B(n_568),
.Y(n_593)
);

NAND2xp5_ASAP7_75t_SL g594 ( 
.A(n_533),
.B(n_550),
.Y(n_594)
);

INVx1_ASAP7_75t_L g595 ( 
.A(n_563),
.Y(n_595)
);

INVx1_ASAP7_75t_L g596 ( 
.A(n_564),
.Y(n_596)
);

NAND2xp5_ASAP7_75t_L g597 ( 
.A(n_555),
.B(n_525),
.Y(n_597)
);

NAND2xp5_ASAP7_75t_L g598 ( 
.A(n_534),
.B(n_525),
.Y(n_598)
);

INVx2_ASAP7_75t_L g599 ( 
.A(n_564),
.Y(n_599)
);

NAND2xp33_ASAP7_75t_L g600 ( 
.A(n_571),
.B(n_502),
.Y(n_600)
);

BUFx6f_ASAP7_75t_L g601 ( 
.A(n_547),
.Y(n_601)
);

INVx2_ASAP7_75t_L g602 ( 
.A(n_567),
.Y(n_602)
);

NAND2xp5_ASAP7_75t_SL g603 ( 
.A(n_533),
.B(n_499),
.Y(n_603)
);

INVx1_ASAP7_75t_SL g604 ( 
.A(n_539),
.Y(n_604)
);

INVx5_ASAP7_75t_L g605 ( 
.A(n_572),
.Y(n_605)
);

INVx1_ASAP7_75t_L g606 ( 
.A(n_567),
.Y(n_606)
);

CKINVDCx20_ASAP7_75t_R g607 ( 
.A(n_545),
.Y(n_607)
);

NAND3xp33_ASAP7_75t_L g608 ( 
.A(n_543),
.B(n_478),
.C(n_434),
.Y(n_608)
);

NAND2xp5_ASAP7_75t_L g609 ( 
.A(n_559),
.B(n_525),
.Y(n_609)
);

INVx2_ASAP7_75t_SL g610 ( 
.A(n_561),
.Y(n_610)
);

INVx2_ASAP7_75t_L g611 ( 
.A(n_551),
.Y(n_611)
);

NOR2xp33_ASAP7_75t_L g612 ( 
.A(n_541),
.B(n_546),
.Y(n_612)
);

NAND2xp33_ASAP7_75t_R g613 ( 
.A(n_559),
.B(n_446),
.Y(n_613)
);

INVx2_ASAP7_75t_SL g614 ( 
.A(n_557),
.Y(n_614)
);

BUFx6f_ASAP7_75t_L g615 ( 
.A(n_569),
.Y(n_615)
);

INVx4_ASAP7_75t_L g616 ( 
.A(n_572),
.Y(n_616)
);

NAND2xp5_ASAP7_75t_SL g617 ( 
.A(n_562),
.B(n_508),
.Y(n_617)
);

BUFx10_ASAP7_75t_L g618 ( 
.A(n_560),
.Y(n_618)
);

INVx2_ASAP7_75t_L g619 ( 
.A(n_573),
.Y(n_619)
);

INVx2_ASAP7_75t_SL g620 ( 
.A(n_542),
.Y(n_620)
);

INVx2_ASAP7_75t_L g621 ( 
.A(n_573),
.Y(n_621)
);

AND2x2_ASAP7_75t_L g622 ( 
.A(n_541),
.B(n_459),
.Y(n_622)
);

INVx2_ASAP7_75t_L g623 ( 
.A(n_573),
.Y(n_623)
);

INVx2_ASAP7_75t_SL g624 ( 
.A(n_554),
.Y(n_624)
);

INVx8_ASAP7_75t_L g625 ( 
.A(n_562),
.Y(n_625)
);

INVx1_ASAP7_75t_L g626 ( 
.A(n_556),
.Y(n_626)
);

INVx2_ASAP7_75t_SL g627 ( 
.A(n_565),
.Y(n_627)
);

INVx2_ASAP7_75t_L g628 ( 
.A(n_565),
.Y(n_628)
);

INVx3_ASAP7_75t_L g629 ( 
.A(n_565),
.Y(n_629)
);

NAND2xp5_ASAP7_75t_SL g630 ( 
.A(n_548),
.B(n_508),
.Y(n_630)
);

BUFx3_ASAP7_75t_L g631 ( 
.A(n_553),
.Y(n_631)
);

CKINVDCx16_ASAP7_75t_R g632 ( 
.A(n_566),
.Y(n_632)
);

INVx1_ASAP7_75t_L g633 ( 
.A(n_566),
.Y(n_633)
);

INVx2_ASAP7_75t_L g634 ( 
.A(n_566),
.Y(n_634)
);

INVx4_ASAP7_75t_L g635 ( 
.A(n_547),
.Y(n_635)
);

NAND2xp5_ASAP7_75t_SL g636 ( 
.A(n_552),
.B(n_508),
.Y(n_636)
);

INVx2_ASAP7_75t_L g637 ( 
.A(n_538),
.Y(n_637)
);

INVx3_ASAP7_75t_L g638 ( 
.A(n_572),
.Y(n_638)
);

INVx2_ASAP7_75t_L g639 ( 
.A(n_538),
.Y(n_639)
);

INVx1_ASAP7_75t_L g640 ( 
.A(n_538),
.Y(n_640)
);

INVx1_ASAP7_75t_L g641 ( 
.A(n_538),
.Y(n_641)
);

AOI22xp33_ASAP7_75t_L g642 ( 
.A1(n_566),
.A2(n_221),
.B1(n_424),
.B2(n_453),
.Y(n_642)
);

INVx3_ASAP7_75t_L g643 ( 
.A(n_572),
.Y(n_643)
);

INVx3_ASAP7_75t_L g644 ( 
.A(n_572),
.Y(n_644)
);

INVx1_ASAP7_75t_L g645 ( 
.A(n_538),
.Y(n_645)
);

INVx2_ASAP7_75t_L g646 ( 
.A(n_538),
.Y(n_646)
);

OAI22xp5_ASAP7_75t_SL g647 ( 
.A1(n_545),
.A2(n_469),
.B1(n_461),
.B2(n_460),
.Y(n_647)
);

AOI22xp33_ASAP7_75t_L g648 ( 
.A1(n_566),
.A2(n_221),
.B1(n_424),
.B2(n_453),
.Y(n_648)
);

HB1xp67_ASAP7_75t_L g649 ( 
.A(n_568),
.Y(n_649)
);

INVx1_ASAP7_75t_L g650 ( 
.A(n_538),
.Y(n_650)
);

AND2x6_ASAP7_75t_L g651 ( 
.A(n_551),
.B(n_502),
.Y(n_651)
);

AND2x6_ASAP7_75t_L g652 ( 
.A(n_551),
.B(n_502),
.Y(n_652)
);

INVx1_ASAP7_75t_L g653 ( 
.A(n_538),
.Y(n_653)
);

NAND2xp5_ASAP7_75t_SL g654 ( 
.A(n_552),
.B(n_508),
.Y(n_654)
);

INVx1_ASAP7_75t_L g655 ( 
.A(n_538),
.Y(n_655)
);

INVx2_ASAP7_75t_L g656 ( 
.A(n_538),
.Y(n_656)
);

NAND2xp5_ASAP7_75t_L g657 ( 
.A(n_537),
.B(n_432),
.Y(n_657)
);

INVx2_ASAP7_75t_SL g658 ( 
.A(n_549),
.Y(n_658)
);

INVx1_ASAP7_75t_L g659 ( 
.A(n_538),
.Y(n_659)
);

INVx1_ASAP7_75t_L g660 ( 
.A(n_611),
.Y(n_660)
);

INVx3_ASAP7_75t_L g661 ( 
.A(n_601),
.Y(n_661)
);

AND2x2_ASAP7_75t_L g662 ( 
.A(n_610),
.B(n_460),
.Y(n_662)
);

INVx4_ASAP7_75t_SL g663 ( 
.A(n_651),
.Y(n_663)
);

INVx1_ASAP7_75t_L g664 ( 
.A(n_611),
.Y(n_664)
);

INVx1_ASAP7_75t_L g665 ( 
.A(n_575),
.Y(n_665)
);

NAND2xp5_ASAP7_75t_L g666 ( 
.A(n_649),
.B(n_456),
.Y(n_666)
);

HB1xp67_ASAP7_75t_L g667 ( 
.A(n_619),
.Y(n_667)
);

NAND2xp5_ASAP7_75t_L g668 ( 
.A(n_598),
.B(n_593),
.Y(n_668)
);

NAND2xp5_ASAP7_75t_L g669 ( 
.A(n_580),
.B(n_503),
.Y(n_669)
);

INVx1_ASAP7_75t_L g670 ( 
.A(n_581),
.Y(n_670)
);

INVx1_ASAP7_75t_L g671 ( 
.A(n_583),
.Y(n_671)
);

INVx1_ASAP7_75t_L g672 ( 
.A(n_592),
.Y(n_672)
);

AND2x4_ASAP7_75t_L g673 ( 
.A(n_588),
.B(n_532),
.Y(n_673)
);

INVx1_ASAP7_75t_L g674 ( 
.A(n_595),
.Y(n_674)
);

NAND2xp5_ASAP7_75t_L g675 ( 
.A(n_589),
.B(n_503),
.Y(n_675)
);

INVx3_ASAP7_75t_L g676 ( 
.A(n_601),
.Y(n_676)
);

HB1xp67_ASAP7_75t_L g677 ( 
.A(n_619),
.Y(n_677)
);

INVx1_ASAP7_75t_L g678 ( 
.A(n_596),
.Y(n_678)
);

INVx2_ASAP7_75t_L g679 ( 
.A(n_585),
.Y(n_679)
);

BUFx2_ASAP7_75t_L g680 ( 
.A(n_584),
.Y(n_680)
);

AND2x4_ASAP7_75t_L g681 ( 
.A(n_588),
.B(n_532),
.Y(n_681)
);

INVx2_ASAP7_75t_L g682 ( 
.A(n_585),
.Y(n_682)
);

OAI22xp5_ASAP7_75t_L g683 ( 
.A1(n_631),
.A2(n_461),
.B1(n_460),
.B2(n_453),
.Y(n_683)
);

INVx2_ASAP7_75t_L g684 ( 
.A(n_599),
.Y(n_684)
);

NAND2xp5_ASAP7_75t_L g685 ( 
.A(n_579),
.B(n_460),
.Y(n_685)
);

INVx2_ASAP7_75t_L g686 ( 
.A(n_599),
.Y(n_686)
);

INVxp33_ASAP7_75t_SL g687 ( 
.A(n_578),
.Y(n_687)
);

NAND2xp5_ASAP7_75t_L g688 ( 
.A(n_609),
.B(n_460),
.Y(n_688)
);

INVx1_ASAP7_75t_L g689 ( 
.A(n_606),
.Y(n_689)
);

CKINVDCx5p33_ASAP7_75t_R g690 ( 
.A(n_591),
.Y(n_690)
);

NAND2xp5_ASAP7_75t_SL g691 ( 
.A(n_608),
.B(n_472),
.Y(n_691)
);

BUFx2_ASAP7_75t_L g692 ( 
.A(n_584),
.Y(n_692)
);

BUFx6f_ASAP7_75t_L g693 ( 
.A(n_601),
.Y(n_693)
);

INVx3_ASAP7_75t_L g694 ( 
.A(n_601),
.Y(n_694)
);

AND2x2_ASAP7_75t_L g695 ( 
.A(n_614),
.B(n_461),
.Y(n_695)
);

NAND2xp5_ASAP7_75t_SL g696 ( 
.A(n_576),
.B(n_472),
.Y(n_696)
);

INVx4_ASAP7_75t_L g697 ( 
.A(n_578),
.Y(n_697)
);

BUFx6f_ASAP7_75t_L g698 ( 
.A(n_615),
.Y(n_698)
);

INVx1_ASAP7_75t_L g699 ( 
.A(n_640),
.Y(n_699)
);

NOR2xp33_ASAP7_75t_L g700 ( 
.A(n_612),
.B(n_481),
.Y(n_700)
);

INVxp67_ASAP7_75t_L g701 ( 
.A(n_612),
.Y(n_701)
);

NAND2xp5_ASAP7_75t_SL g702 ( 
.A(n_576),
.B(n_481),
.Y(n_702)
);

INVx3_ASAP7_75t_L g703 ( 
.A(n_588),
.Y(n_703)
);

AND2x4_ASAP7_75t_L g704 ( 
.A(n_635),
.B(n_532),
.Y(n_704)
);

NOR2xp33_ASAP7_75t_L g705 ( 
.A(n_657),
.B(n_481),
.Y(n_705)
);

NAND2xp5_ASAP7_75t_L g706 ( 
.A(n_604),
.B(n_461),
.Y(n_706)
);

INVx2_ASAP7_75t_SL g707 ( 
.A(n_658),
.Y(n_707)
);

INVx4_ASAP7_75t_L g708 ( 
.A(n_590),
.Y(n_708)
);

INVx2_ASAP7_75t_L g709 ( 
.A(n_602),
.Y(n_709)
);

INVx1_ASAP7_75t_L g710 ( 
.A(n_641),
.Y(n_710)
);

INVx2_ASAP7_75t_L g711 ( 
.A(n_602),
.Y(n_711)
);

INVx2_ASAP7_75t_L g712 ( 
.A(n_637),
.Y(n_712)
);

AND2x2_ASAP7_75t_SL g713 ( 
.A(n_632),
.B(n_461),
.Y(n_713)
);

AND2x2_ASAP7_75t_L g714 ( 
.A(n_620),
.B(n_449),
.Y(n_714)
);

INVx4_ASAP7_75t_L g715 ( 
.A(n_590),
.Y(n_715)
);

CKINVDCx6p67_ASAP7_75t_R g716 ( 
.A(n_622),
.Y(n_716)
);

INVx2_ASAP7_75t_L g717 ( 
.A(n_637),
.Y(n_717)
);

AND2x4_ASAP7_75t_L g718 ( 
.A(n_635),
.B(n_532),
.Y(n_718)
);

NOR2xp33_ASAP7_75t_L g719 ( 
.A(n_624),
.B(n_631),
.Y(n_719)
);

INVx3_ASAP7_75t_L g720 ( 
.A(n_635),
.Y(n_720)
);

AND2x2_ASAP7_75t_L g721 ( 
.A(n_597),
.B(n_449),
.Y(n_721)
);

NOR2xp33_ASAP7_75t_SL g722 ( 
.A(n_591),
.B(n_447),
.Y(n_722)
);

BUFx6f_ASAP7_75t_L g723 ( 
.A(n_615),
.Y(n_723)
);

NAND2xp5_ASAP7_75t_L g724 ( 
.A(n_626),
.B(n_419),
.Y(n_724)
);

OAI22xp5_ASAP7_75t_L g725 ( 
.A1(n_607),
.A2(n_462),
.B1(n_475),
.B2(n_419),
.Y(n_725)
);

INVx1_ASAP7_75t_L g726 ( 
.A(n_645),
.Y(n_726)
);

BUFx6f_ASAP7_75t_L g727 ( 
.A(n_615),
.Y(n_727)
);

INVx1_ASAP7_75t_L g728 ( 
.A(n_650),
.Y(n_728)
);

BUFx6f_ASAP7_75t_L g729 ( 
.A(n_618),
.Y(n_729)
);

AOI22xp33_ASAP7_75t_L g730 ( 
.A1(n_594),
.A2(n_193),
.B1(n_215),
.B2(n_207),
.Y(n_730)
);

INVx2_ASAP7_75t_L g731 ( 
.A(n_639),
.Y(n_731)
);

AND2x6_ASAP7_75t_L g732 ( 
.A(n_634),
.B(n_502),
.Y(n_732)
);

INVx5_ASAP7_75t_L g733 ( 
.A(n_651),
.Y(n_733)
);

AND2x2_ASAP7_75t_L g734 ( 
.A(n_628),
.B(n_449),
.Y(n_734)
);

INVx1_ASAP7_75t_L g735 ( 
.A(n_653),
.Y(n_735)
);

AND2x4_ASAP7_75t_L g736 ( 
.A(n_586),
.B(n_638),
.Y(n_736)
);

INVx2_ASAP7_75t_L g737 ( 
.A(n_639),
.Y(n_737)
);

NAND2xp5_ASAP7_75t_L g738 ( 
.A(n_594),
.B(n_577),
.Y(n_738)
);

INVx4_ASAP7_75t_L g739 ( 
.A(n_605),
.Y(n_739)
);

NOR2xp33_ASAP7_75t_R g740 ( 
.A(n_613),
.B(n_421),
.Y(n_740)
);

INVx3_ASAP7_75t_L g741 ( 
.A(n_618),
.Y(n_741)
);

BUFx6f_ASAP7_75t_L g742 ( 
.A(n_618),
.Y(n_742)
);

NAND2xp5_ASAP7_75t_SL g743 ( 
.A(n_574),
.B(n_481),
.Y(n_743)
);

INVx3_ASAP7_75t_L g744 ( 
.A(n_616),
.Y(n_744)
);

NAND2xp5_ASAP7_75t_L g745 ( 
.A(n_655),
.B(n_462),
.Y(n_745)
);

NAND2xp5_ASAP7_75t_L g746 ( 
.A(n_701),
.B(n_668),
.Y(n_746)
);

INVx1_ASAP7_75t_L g747 ( 
.A(n_667),
.Y(n_747)
);

NOR2xp33_ASAP7_75t_L g748 ( 
.A(n_701),
.B(n_633),
.Y(n_748)
);

INVx2_ASAP7_75t_L g749 ( 
.A(n_660),
.Y(n_749)
);

INVx2_ASAP7_75t_L g750 ( 
.A(n_664),
.Y(n_750)
);

INVxp67_ASAP7_75t_L g751 ( 
.A(n_666),
.Y(n_751)
);

INVx2_ASAP7_75t_L g752 ( 
.A(n_665),
.Y(n_752)
);

NAND3xp33_ASAP7_75t_L g753 ( 
.A(n_730),
.B(n_648),
.C(n_642),
.Y(n_753)
);

INVx2_ASAP7_75t_L g754 ( 
.A(n_670),
.Y(n_754)
);

INVx1_ASAP7_75t_L g755 ( 
.A(n_667),
.Y(n_755)
);

INVx8_ASAP7_75t_L g756 ( 
.A(n_690),
.Y(n_756)
);

INVx2_ASAP7_75t_L g757 ( 
.A(n_671),
.Y(n_757)
);

AOI22xp5_ASAP7_75t_L g758 ( 
.A1(n_738),
.A2(n_647),
.B1(n_607),
.B2(n_625),
.Y(n_758)
);

NAND2xp5_ASAP7_75t_L g759 ( 
.A(n_688),
.B(n_628),
.Y(n_759)
);

INVx2_ASAP7_75t_L g760 ( 
.A(n_672),
.Y(n_760)
);

NAND2xp5_ASAP7_75t_L g761 ( 
.A(n_685),
.B(n_634),
.Y(n_761)
);

NAND2xp5_ASAP7_75t_L g762 ( 
.A(n_721),
.B(n_627),
.Y(n_762)
);

OR2x6_ASAP7_75t_L g763 ( 
.A(n_743),
.B(n_625),
.Y(n_763)
);

BUFx3_ASAP7_75t_L g764 ( 
.A(n_698),
.Y(n_764)
);

NAND2xp5_ASAP7_75t_SL g765 ( 
.A(n_740),
.B(n_625),
.Y(n_765)
);

OR2x6_ASAP7_75t_L g766 ( 
.A(n_743),
.B(n_621),
.Y(n_766)
);

INVx2_ASAP7_75t_L g767 ( 
.A(n_674),
.Y(n_767)
);

NAND2xp5_ASAP7_75t_L g768 ( 
.A(n_706),
.B(n_629),
.Y(n_768)
);

NAND2xp5_ASAP7_75t_L g769 ( 
.A(n_700),
.B(n_629),
.Y(n_769)
);

AND2x2_ASAP7_75t_L g770 ( 
.A(n_662),
.B(n_621),
.Y(n_770)
);

INVx2_ASAP7_75t_L g771 ( 
.A(n_678),
.Y(n_771)
);

INVx2_ASAP7_75t_L g772 ( 
.A(n_689),
.Y(n_772)
);

AOI21x1_ASAP7_75t_L g773 ( 
.A1(n_691),
.A2(n_636),
.B(n_574),
.Y(n_773)
);

AOI22xp5_ASAP7_75t_L g774 ( 
.A1(n_730),
.A2(n_642),
.B1(n_648),
.B2(n_613),
.Y(n_774)
);

NOR2xp33_ASAP7_75t_L g775 ( 
.A(n_700),
.B(n_630),
.Y(n_775)
);

INVx2_ASAP7_75t_L g776 ( 
.A(n_699),
.Y(n_776)
);

NAND2xp5_ASAP7_75t_L g777 ( 
.A(n_710),
.B(n_726),
.Y(n_777)
);

INVx1_ASAP7_75t_L g778 ( 
.A(n_677),
.Y(n_778)
);

INVx2_ASAP7_75t_L g779 ( 
.A(n_728),
.Y(n_779)
);

INVxp33_ASAP7_75t_L g780 ( 
.A(n_740),
.Y(n_780)
);

AO221x1_ASAP7_75t_L g781 ( 
.A1(n_729),
.A2(n_623),
.B1(n_643),
.B2(n_586),
.C(n_638),
.Y(n_781)
);

OA21x2_ASAP7_75t_L g782 ( 
.A1(n_691),
.A2(n_623),
.B(n_636),
.Y(n_782)
);

INVx2_ASAP7_75t_L g783 ( 
.A(n_735),
.Y(n_783)
);

NOR2xp33_ASAP7_75t_L g784 ( 
.A(n_669),
.B(n_630),
.Y(n_784)
);

INVx1_ASAP7_75t_L g785 ( 
.A(n_677),
.Y(n_785)
);

NOR2xp33_ASAP7_75t_L g786 ( 
.A(n_675),
.B(n_603),
.Y(n_786)
);

NAND2xp5_ASAP7_75t_SL g787 ( 
.A(n_713),
.B(n_654),
.Y(n_787)
);

NAND2xp5_ASAP7_75t_L g788 ( 
.A(n_724),
.B(n_603),
.Y(n_788)
);

NAND2xp5_ASAP7_75t_L g789 ( 
.A(n_745),
.B(n_659),
.Y(n_789)
);

NAND2xp5_ASAP7_75t_L g790 ( 
.A(n_705),
.B(n_646),
.Y(n_790)
);

INVx2_ASAP7_75t_L g791 ( 
.A(n_679),
.Y(n_791)
);

AND2x2_ASAP7_75t_L g792 ( 
.A(n_695),
.B(n_643),
.Y(n_792)
);

NAND2x1_ASAP7_75t_L g793 ( 
.A(n_744),
.B(n_651),
.Y(n_793)
);

INVx1_ASAP7_75t_L g794 ( 
.A(n_679),
.Y(n_794)
);

INVx1_ASAP7_75t_L g795 ( 
.A(n_682),
.Y(n_795)
);

INVx2_ASAP7_75t_SL g796 ( 
.A(n_707),
.Y(n_796)
);

INVx1_ASAP7_75t_L g797 ( 
.A(n_682),
.Y(n_797)
);

NOR3xp33_ASAP7_75t_L g798 ( 
.A(n_683),
.B(n_719),
.C(n_725),
.Y(n_798)
);

NOR2xp33_ASAP7_75t_L g799 ( 
.A(n_719),
.B(n_654),
.Y(n_799)
);

NAND2xp5_ASAP7_75t_SL g800 ( 
.A(n_713),
.B(n_605),
.Y(n_800)
);

INVx2_ASAP7_75t_SL g801 ( 
.A(n_698),
.Y(n_801)
);

NOR2xp33_ASAP7_75t_L g802 ( 
.A(n_696),
.B(n_617),
.Y(n_802)
);

NAND2xp5_ASAP7_75t_L g803 ( 
.A(n_705),
.B(n_646),
.Y(n_803)
);

AND2x4_ASAP7_75t_L g804 ( 
.A(n_663),
.B(n_605),
.Y(n_804)
);

NAND2xp5_ASAP7_75t_L g805 ( 
.A(n_680),
.B(n_656),
.Y(n_805)
);

INVx2_ASAP7_75t_L g806 ( 
.A(n_684),
.Y(n_806)
);

NAND2xp5_ASAP7_75t_L g807 ( 
.A(n_692),
.B(n_656),
.Y(n_807)
);

AND2x2_ASAP7_75t_L g808 ( 
.A(n_716),
.B(n_644),
.Y(n_808)
);

INVx1_ASAP7_75t_L g809 ( 
.A(n_684),
.Y(n_809)
);

INVx2_ASAP7_75t_L g810 ( 
.A(n_686),
.Y(n_810)
);

INVx1_ASAP7_75t_L g811 ( 
.A(n_686),
.Y(n_811)
);

INVx1_ASAP7_75t_L g812 ( 
.A(n_709),
.Y(n_812)
);

NAND2xp5_ASAP7_75t_L g813 ( 
.A(n_736),
.B(n_617),
.Y(n_813)
);

NOR2xp33_ASAP7_75t_L g814 ( 
.A(n_696),
.B(n_582),
.Y(n_814)
);

BUFx3_ASAP7_75t_L g815 ( 
.A(n_698),
.Y(n_815)
);

HB1xp67_ASAP7_75t_L g816 ( 
.A(n_736),
.Y(n_816)
);

AOI221x1_ASAP7_75t_L g817 ( 
.A1(n_661),
.A2(n_217),
.B1(n_204),
.B2(n_185),
.C(n_194),
.Y(n_817)
);

INVx2_ASAP7_75t_L g818 ( 
.A(n_709),
.Y(n_818)
);

INVx2_ASAP7_75t_L g819 ( 
.A(n_711),
.Y(n_819)
);

NAND2xp5_ASAP7_75t_SL g820 ( 
.A(n_798),
.B(n_697),
.Y(n_820)
);

INVx1_ASAP7_75t_L g821 ( 
.A(n_752),
.Y(n_821)
);

NAND2xp5_ASAP7_75t_L g822 ( 
.A(n_751),
.B(n_702),
.Y(n_822)
);

INVxp67_ASAP7_75t_SL g823 ( 
.A(n_747),
.Y(n_823)
);

NAND2xp5_ASAP7_75t_L g824 ( 
.A(n_746),
.B(n_702),
.Y(n_824)
);

NAND2xp5_ASAP7_75t_L g825 ( 
.A(n_784),
.B(n_736),
.Y(n_825)
);

AND2x2_ASAP7_75t_L g826 ( 
.A(n_816),
.B(n_697),
.Y(n_826)
);

NOR2x1p5_ASAP7_75t_L g827 ( 
.A(n_788),
.B(n_690),
.Y(n_827)
);

NAND2xp5_ASAP7_75t_SL g828 ( 
.A(n_799),
.B(n_708),
.Y(n_828)
);

INVx1_ASAP7_75t_L g829 ( 
.A(n_752),
.Y(n_829)
);

NOR2xp33_ASAP7_75t_R g830 ( 
.A(n_756),
.B(n_421),
.Y(n_830)
);

NAND2xp5_ASAP7_75t_L g831 ( 
.A(n_784),
.B(n_734),
.Y(n_831)
);

NAND2xp5_ASAP7_75t_L g832 ( 
.A(n_786),
.B(n_714),
.Y(n_832)
);

AND2x2_ASAP7_75t_L g833 ( 
.A(n_808),
.B(n_708),
.Y(n_833)
);

NAND2xp5_ASAP7_75t_SL g834 ( 
.A(n_799),
.B(n_715),
.Y(n_834)
);

BUFx6f_ASAP7_75t_L g835 ( 
.A(n_764),
.Y(n_835)
);

NOR2xp33_ASAP7_75t_L g836 ( 
.A(n_775),
.B(n_661),
.Y(n_836)
);

NAND2xp5_ASAP7_75t_SL g837 ( 
.A(n_780),
.B(n_775),
.Y(n_837)
);

NOR2xp33_ASAP7_75t_L g838 ( 
.A(n_780),
.B(n_715),
.Y(n_838)
);

NAND2xp5_ASAP7_75t_L g839 ( 
.A(n_786),
.B(n_711),
.Y(n_839)
);

NAND2xp5_ASAP7_75t_SL g840 ( 
.A(n_765),
.B(n_729),
.Y(n_840)
);

NAND2xp5_ASAP7_75t_L g841 ( 
.A(n_748),
.B(n_814),
.Y(n_841)
);

NAND2xp5_ASAP7_75t_L g842 ( 
.A(n_748),
.B(n_712),
.Y(n_842)
);

INVx1_ASAP7_75t_L g843 ( 
.A(n_754),
.Y(n_843)
);

AOI22xp33_ASAP7_75t_L g844 ( 
.A1(n_753),
.A2(n_199),
.B1(n_224),
.B2(n_217),
.Y(n_844)
);

OR2x2_ASAP7_75t_L g845 ( 
.A(n_762),
.B(n_712),
.Y(n_845)
);

INVx1_ASAP7_75t_L g846 ( 
.A(n_754),
.Y(n_846)
);

AND2x4_ASAP7_75t_SL g847 ( 
.A(n_804),
.B(n_698),
.Y(n_847)
);

O2A1O1Ixp5_ASAP7_75t_L g848 ( 
.A1(n_787),
.A2(n_582),
.B(n_739),
.C(n_720),
.Y(n_848)
);

HB1xp67_ASAP7_75t_L g849 ( 
.A(n_755),
.Y(n_849)
);

AOI22xp33_ASAP7_75t_L g850 ( 
.A1(n_774),
.A2(n_758),
.B1(n_814),
.B2(n_802),
.Y(n_850)
);

NAND2xp5_ASAP7_75t_L g851 ( 
.A(n_802),
.B(n_717),
.Y(n_851)
);

INVx3_ASAP7_75t_L g852 ( 
.A(n_764),
.Y(n_852)
);

OR2x2_ASAP7_75t_L g853 ( 
.A(n_778),
.B(n_717),
.Y(n_853)
);

OAI22xp5_ASAP7_75t_L g854 ( 
.A1(n_765),
.A2(n_687),
.B1(n_733),
.B2(n_694),
.Y(n_854)
);

NAND2xp5_ASAP7_75t_SL g855 ( 
.A(n_804),
.B(n_729),
.Y(n_855)
);

INVx2_ASAP7_75t_L g856 ( 
.A(n_757),
.Y(n_856)
);

OAI221xp5_ASAP7_75t_L g857 ( 
.A1(n_796),
.A2(n_475),
.B1(n_722),
.B2(n_225),
.C(n_191),
.Y(n_857)
);

AO221x1_ASAP7_75t_L g858 ( 
.A1(n_785),
.A2(n_742),
.B1(n_729),
.B2(n_693),
.C(n_741),
.Y(n_858)
);

OAI22xp33_ASAP7_75t_L g859 ( 
.A1(n_787),
.A2(n_733),
.B1(n_687),
.B2(n_605),
.Y(n_859)
);

NAND2xp5_ASAP7_75t_L g860 ( 
.A(n_790),
.B(n_731),
.Y(n_860)
);

NAND2xp5_ASAP7_75t_L g861 ( 
.A(n_803),
.B(n_731),
.Y(n_861)
);

AND2x2_ASAP7_75t_L g862 ( 
.A(n_770),
.B(n_676),
.Y(n_862)
);

NAND2xp5_ASAP7_75t_L g863 ( 
.A(n_761),
.B(n_737),
.Y(n_863)
);

NOR2xp33_ASAP7_75t_L g864 ( 
.A(n_789),
.B(n_723),
.Y(n_864)
);

AND2x2_ASAP7_75t_L g865 ( 
.A(n_792),
.B(n_769),
.Y(n_865)
);

NOR2xp33_ASAP7_75t_L g866 ( 
.A(n_756),
.B(n_723),
.Y(n_866)
);

HB1xp67_ASAP7_75t_L g867 ( 
.A(n_819),
.Y(n_867)
);

NOR2xp33_ASAP7_75t_SL g868 ( 
.A(n_756),
.B(n_447),
.Y(n_868)
);

NAND2xp5_ASAP7_75t_L g869 ( 
.A(n_759),
.B(n_737),
.Y(n_869)
);

NOR2xp33_ASAP7_75t_L g870 ( 
.A(n_813),
.B(n_694),
.Y(n_870)
);

INVx1_ASAP7_75t_L g871 ( 
.A(n_757),
.Y(n_871)
);

BUFx3_ASAP7_75t_L g872 ( 
.A(n_815),
.Y(n_872)
);

NAND2xp5_ASAP7_75t_L g873 ( 
.A(n_805),
.B(n_741),
.Y(n_873)
);

AND2x6_ASAP7_75t_SL g874 ( 
.A(n_768),
.B(n_518),
.Y(n_874)
);

NAND2xp5_ASAP7_75t_SL g875 ( 
.A(n_804),
.B(n_742),
.Y(n_875)
);

INVx2_ASAP7_75t_L g876 ( 
.A(n_760),
.Y(n_876)
);

INVx4_ASAP7_75t_L g877 ( 
.A(n_815),
.Y(n_877)
);

NAND2xp5_ASAP7_75t_L g878 ( 
.A(n_807),
.B(n_703),
.Y(n_878)
);

NAND2xp5_ASAP7_75t_L g879 ( 
.A(n_760),
.B(n_703),
.Y(n_879)
);

AND2x2_ASAP7_75t_L g880 ( 
.A(n_767),
.B(n_771),
.Y(n_880)
);

NAND2xp5_ASAP7_75t_SL g881 ( 
.A(n_800),
.B(n_742),
.Y(n_881)
);

INVxp67_ASAP7_75t_L g882 ( 
.A(n_777),
.Y(n_882)
);

NOR2xp33_ASAP7_75t_L g883 ( 
.A(n_801),
.B(n_723),
.Y(n_883)
);

OR2x6_ASAP7_75t_L g884 ( 
.A(n_763),
.B(n_739),
.Y(n_884)
);

NAND2xp5_ASAP7_75t_L g885 ( 
.A(n_767),
.B(n_720),
.Y(n_885)
);

NOR2xp67_ASAP7_75t_L g886 ( 
.A(n_771),
.B(n_733),
.Y(n_886)
);

NOR3xp33_ASAP7_75t_L g887 ( 
.A(n_800),
.B(n_600),
.C(n_744),
.Y(n_887)
);

NAND2xp5_ASAP7_75t_L g888 ( 
.A(n_772),
.B(n_693),
.Y(n_888)
);

INVx2_ASAP7_75t_L g889 ( 
.A(n_772),
.Y(n_889)
);

NAND2xp5_ASAP7_75t_L g890 ( 
.A(n_776),
.B(n_693),
.Y(n_890)
);

INVx1_ASAP7_75t_L g891 ( 
.A(n_776),
.Y(n_891)
);

AOI22xp33_ASAP7_75t_L g892 ( 
.A1(n_763),
.A2(n_224),
.B1(n_204),
.B2(n_222),
.Y(n_892)
);

NOR2xp33_ASAP7_75t_L g893 ( 
.A(n_779),
.B(n_723),
.Y(n_893)
);

NAND2xp5_ASAP7_75t_L g894 ( 
.A(n_779),
.B(n_693),
.Y(n_894)
);

NAND2xp5_ASAP7_75t_SL g895 ( 
.A(n_783),
.B(n_742),
.Y(n_895)
);

INVx2_ASAP7_75t_L g896 ( 
.A(n_783),
.Y(n_896)
);

AOI21xp5_ASAP7_75t_L g897 ( 
.A1(n_817),
.A2(n_600),
.B(n_733),
.Y(n_897)
);

NAND2x1p5_ASAP7_75t_L g898 ( 
.A(n_886),
.B(n_793),
.Y(n_898)
);

NAND2xp5_ASAP7_75t_L g899 ( 
.A(n_882),
.B(n_841),
.Y(n_899)
);

INVx1_ASAP7_75t_L g900 ( 
.A(n_867),
.Y(n_900)
);

INVx1_ASAP7_75t_L g901 ( 
.A(n_867),
.Y(n_901)
);

INVx2_ASAP7_75t_L g902 ( 
.A(n_880),
.Y(n_902)
);

NAND2x1p5_ASAP7_75t_L g903 ( 
.A(n_877),
.B(n_773),
.Y(n_903)
);

INVx1_ASAP7_75t_L g904 ( 
.A(n_849),
.Y(n_904)
);

NAND2xp5_ASAP7_75t_L g905 ( 
.A(n_882),
.B(n_749),
.Y(n_905)
);

BUFx3_ASAP7_75t_L g906 ( 
.A(n_833),
.Y(n_906)
);

INVx1_ASAP7_75t_L g907 ( 
.A(n_849),
.Y(n_907)
);

NAND2x1p5_ASAP7_75t_L g908 ( 
.A(n_877),
.B(n_782),
.Y(n_908)
);

INVx1_ASAP7_75t_L g909 ( 
.A(n_821),
.Y(n_909)
);

INVx1_ASAP7_75t_L g910 ( 
.A(n_829),
.Y(n_910)
);

NAND2x1p5_ASAP7_75t_L g911 ( 
.A(n_881),
.B(n_782),
.Y(n_911)
);

NAND2x1p5_ASAP7_75t_L g912 ( 
.A(n_840),
.B(n_782),
.Y(n_912)
);

BUFx8_ASAP7_75t_L g913 ( 
.A(n_830),
.Y(n_913)
);

AND2x4_ASAP7_75t_L g914 ( 
.A(n_884),
.B(n_749),
.Y(n_914)
);

INVx2_ASAP7_75t_L g915 ( 
.A(n_843),
.Y(n_915)
);

INVx1_ASAP7_75t_L g916 ( 
.A(n_846),
.Y(n_916)
);

NOR2xp33_ASAP7_75t_R g917 ( 
.A(n_868),
.B(n_727),
.Y(n_917)
);

INVx1_ASAP7_75t_L g918 ( 
.A(n_871),
.Y(n_918)
);

AO22x2_ASAP7_75t_L g919 ( 
.A1(n_823),
.A2(n_750),
.B1(n_795),
.B2(n_794),
.Y(n_919)
);

INVx1_ASAP7_75t_L g920 ( 
.A(n_891),
.Y(n_920)
);

INVx2_ASAP7_75t_L g921 ( 
.A(n_856),
.Y(n_921)
);

INVx1_ASAP7_75t_L g922 ( 
.A(n_823),
.Y(n_922)
);

INVx1_ASAP7_75t_L g923 ( 
.A(n_876),
.Y(n_923)
);

INVx1_ASAP7_75t_L g924 ( 
.A(n_889),
.Y(n_924)
);

INVx1_ASAP7_75t_L g925 ( 
.A(n_896),
.Y(n_925)
);

AO22x2_ASAP7_75t_L g926 ( 
.A1(n_854),
.A2(n_750),
.B1(n_809),
.B2(n_797),
.Y(n_926)
);

AO22x2_ASAP7_75t_L g927 ( 
.A1(n_828),
.A2(n_812),
.B1(n_811),
.B2(n_791),
.Y(n_927)
);

INVx1_ASAP7_75t_L g928 ( 
.A(n_853),
.Y(n_928)
);

AOI22xp5_ASAP7_75t_L g929 ( 
.A1(n_850),
.A2(n_763),
.B1(n_681),
.B2(n_718),
.Y(n_929)
);

INVxp67_ASAP7_75t_L g930 ( 
.A(n_837),
.Y(n_930)
);

INVx2_ASAP7_75t_L g931 ( 
.A(n_852),
.Y(n_931)
);

NAND2xp5_ASAP7_75t_L g932 ( 
.A(n_839),
.B(n_791),
.Y(n_932)
);

INVx2_ASAP7_75t_L g933 ( 
.A(n_852),
.Y(n_933)
);

INVx1_ASAP7_75t_L g934 ( 
.A(n_845),
.Y(n_934)
);

AND2x2_ASAP7_75t_L g935 ( 
.A(n_865),
.B(n_806),
.Y(n_935)
);

NAND2xp5_ASAP7_75t_L g936 ( 
.A(n_851),
.B(n_806),
.Y(n_936)
);

AO22x2_ASAP7_75t_L g937 ( 
.A1(n_834),
.A2(n_810),
.B1(n_819),
.B2(n_818),
.Y(n_937)
);

AO22x2_ASAP7_75t_L g938 ( 
.A1(n_822),
.A2(n_820),
.B1(n_895),
.B2(n_875),
.Y(n_938)
);

NOR2xp33_ASAP7_75t_L g939 ( 
.A(n_838),
.B(n_727),
.Y(n_939)
);

INVx1_ASAP7_75t_L g940 ( 
.A(n_860),
.Y(n_940)
);

AO22x2_ASAP7_75t_L g941 ( 
.A1(n_855),
.A2(n_810),
.B1(n_818),
.B2(n_663),
.Y(n_941)
);

NAND2xp5_ASAP7_75t_L g942 ( 
.A(n_824),
.B(n_832),
.Y(n_942)
);

INVx1_ASAP7_75t_L g943 ( 
.A(n_888),
.Y(n_943)
);

NOR2xp67_ASAP7_75t_L g944 ( 
.A(n_825),
.B(n_727),
.Y(n_944)
);

INVx1_ASAP7_75t_L g945 ( 
.A(n_890),
.Y(n_945)
);

INVx1_ASAP7_75t_L g946 ( 
.A(n_861),
.Y(n_946)
);

AO22x2_ASAP7_75t_L g947 ( 
.A1(n_879),
.A2(n_663),
.B1(n_681),
.B2(n_673),
.Y(n_947)
);

OR2x2_ASAP7_75t_L g948 ( 
.A(n_831),
.B(n_766),
.Y(n_948)
);

AND2x2_ASAP7_75t_L g949 ( 
.A(n_826),
.B(n_766),
.Y(n_949)
);

INVx2_ASAP7_75t_L g950 ( 
.A(n_835),
.Y(n_950)
);

AND2x4_ASAP7_75t_L g951 ( 
.A(n_884),
.B(n_766),
.Y(n_951)
);

INVx1_ASAP7_75t_L g952 ( 
.A(n_842),
.Y(n_952)
);

INVxp67_ASAP7_75t_L g953 ( 
.A(n_836),
.Y(n_953)
);

A2O1A1Ixp33_ASAP7_75t_L g954 ( 
.A1(n_930),
.A2(n_850),
.B(n_892),
.C(n_848),
.Y(n_954)
);

AND2x2_ASAP7_75t_L g955 ( 
.A(n_906),
.B(n_862),
.Y(n_955)
);

INVx1_ASAP7_75t_L g956 ( 
.A(n_904),
.Y(n_956)
);

INVx2_ASAP7_75t_SL g957 ( 
.A(n_950),
.Y(n_957)
);

O2A1O1Ixp33_ASAP7_75t_L g958 ( 
.A1(n_899),
.A2(n_892),
.B(n_844),
.C(n_859),
.Y(n_958)
);

NOR2xp33_ASAP7_75t_L g959 ( 
.A(n_913),
.B(n_953),
.Y(n_959)
);

INVx1_ASAP7_75t_L g960 ( 
.A(n_907),
.Y(n_960)
);

NAND2xp5_ASAP7_75t_L g961 ( 
.A(n_952),
.B(n_836),
.Y(n_961)
);

AOI22xp5_ASAP7_75t_L g962 ( 
.A1(n_929),
.A2(n_859),
.B1(n_844),
.B2(n_884),
.Y(n_962)
);

NAND2xp5_ASAP7_75t_SL g963 ( 
.A(n_917),
.B(n_848),
.Y(n_963)
);

AOI21xp5_ASAP7_75t_L g964 ( 
.A1(n_938),
.A2(n_897),
.B(n_887),
.Y(n_964)
);

NOR2xp67_ASAP7_75t_L g965 ( 
.A(n_900),
.B(n_866),
.Y(n_965)
);

AOI21xp5_ASAP7_75t_L g966 ( 
.A1(n_938),
.A2(n_887),
.B(n_858),
.Y(n_966)
);

HB1xp67_ASAP7_75t_L g967 ( 
.A(n_922),
.Y(n_967)
);

AO21x1_ASAP7_75t_L g968 ( 
.A1(n_908),
.A2(n_870),
.B(n_864),
.Y(n_968)
);

INVx2_ASAP7_75t_L g969 ( 
.A(n_919),
.Y(n_969)
);

AOI21xp5_ASAP7_75t_L g970 ( 
.A1(n_947),
.A2(n_781),
.B(n_878),
.Y(n_970)
);

NAND2xp5_ASAP7_75t_L g971 ( 
.A(n_952),
.B(n_942),
.Y(n_971)
);

BUFx2_ASAP7_75t_L g972 ( 
.A(n_898),
.Y(n_972)
);

AO21x1_ASAP7_75t_L g973 ( 
.A1(n_911),
.A2(n_870),
.B(n_893),
.Y(n_973)
);

NAND2xp5_ASAP7_75t_L g974 ( 
.A(n_943),
.B(n_873),
.Y(n_974)
);

AND2x2_ASAP7_75t_L g975 ( 
.A(n_949),
.B(n_872),
.Y(n_975)
);

NAND2xp5_ASAP7_75t_L g976 ( 
.A(n_945),
.B(n_885),
.Y(n_976)
);

INVxp67_ASAP7_75t_L g977 ( 
.A(n_905),
.Y(n_977)
);

BUFx6f_ASAP7_75t_L g978 ( 
.A(n_903),
.Y(n_978)
);

AOI21xp5_ASAP7_75t_L g979 ( 
.A1(n_947),
.A2(n_857),
.B(n_863),
.Y(n_979)
);

NAND2xp5_ASAP7_75t_SL g980 ( 
.A(n_913),
.B(n_835),
.Y(n_980)
);

NAND2xp5_ASAP7_75t_L g981 ( 
.A(n_940),
.B(n_894),
.Y(n_981)
);

AOI21xp33_ASAP7_75t_L g982 ( 
.A1(n_926),
.A2(n_883),
.B(n_869),
.Y(n_982)
);

NOR2xp33_ASAP7_75t_SL g983 ( 
.A(n_951),
.B(n_835),
.Y(n_983)
);

NOR3xp33_ASAP7_75t_L g984 ( 
.A(n_939),
.B(n_208),
.C(n_176),
.Y(n_984)
);

CKINVDCx5p33_ASAP7_75t_R g985 ( 
.A(n_931),
.Y(n_985)
);

O2A1O1Ixp33_ASAP7_75t_L g986 ( 
.A1(n_912),
.A2(n_827),
.B(n_210),
.C(n_216),
.Y(n_986)
);

AOI21xp5_ASAP7_75t_L g987 ( 
.A1(n_941),
.A2(n_847),
.B(n_681),
.Y(n_987)
);

NAND2xp5_ASAP7_75t_L g988 ( 
.A(n_940),
.B(n_835),
.Y(n_988)
);

AOI21xp5_ASAP7_75t_L g989 ( 
.A1(n_941),
.A2(n_718),
.B(n_673),
.Y(n_989)
);

AOI22xp33_ASAP7_75t_L g990 ( 
.A1(n_951),
.A2(n_732),
.B1(n_718),
.B2(n_673),
.Y(n_990)
);

NAND2xp5_ASAP7_75t_L g991 ( 
.A(n_946),
.B(n_874),
.Y(n_991)
);

OAI22xp5_ASAP7_75t_L g992 ( 
.A1(n_948),
.A2(n_944),
.B1(n_927),
.B2(n_926),
.Y(n_992)
);

HB1xp67_ASAP7_75t_L g993 ( 
.A(n_927),
.Y(n_993)
);

AOI21xp5_ASAP7_75t_L g994 ( 
.A1(n_937),
.A2(n_919),
.B(n_936),
.Y(n_994)
);

AOI21xp5_ASAP7_75t_L g995 ( 
.A1(n_937),
.A2(n_704),
.B(n_644),
.Y(n_995)
);

AOI21xp5_ASAP7_75t_L g996 ( 
.A1(n_932),
.A2(n_704),
.B(n_616),
.Y(n_996)
);

INVx2_ASAP7_75t_L g997 ( 
.A(n_915),
.Y(n_997)
);

INVx3_ASAP7_75t_L g998 ( 
.A(n_914),
.Y(n_998)
);

NOR2xp33_ASAP7_75t_L g999 ( 
.A(n_934),
.B(n_213),
.Y(n_999)
);

NOR2xp33_ASAP7_75t_L g1000 ( 
.A(n_928),
.B(n_218),
.Y(n_1000)
);

AOI21xp5_ASAP7_75t_L g1001 ( 
.A1(n_946),
.A2(n_616),
.B(n_211),
.Y(n_1001)
);

INVx1_ASAP7_75t_L g1002 ( 
.A(n_909),
.Y(n_1002)
);

O2A1O1Ixp5_ASAP7_75t_L g1003 ( 
.A1(n_914),
.A2(n_432),
.B(n_732),
.C(n_498),
.Y(n_1003)
);

NAND2xp5_ASAP7_75t_L g1004 ( 
.A(n_935),
.B(n_732),
.Y(n_1004)
);

AOI22xp5_ASAP7_75t_L g1005 ( 
.A1(n_933),
.A2(n_732),
.B1(n_652),
.B2(n_651),
.Y(n_1005)
);

INVx2_ASAP7_75t_SL g1006 ( 
.A(n_902),
.Y(n_1006)
);

AOI22xp5_ASAP7_75t_L g1007 ( 
.A1(n_910),
.A2(n_732),
.B1(n_652),
.B2(n_651),
.Y(n_1007)
);

NAND2xp5_ASAP7_75t_L g1008 ( 
.A(n_923),
.B(n_587),
.Y(n_1008)
);

AO21x1_ASAP7_75t_L g1009 ( 
.A1(n_916),
.A2(n_0),
.B(n_1),
.Y(n_1009)
);

NAND2xp5_ASAP7_75t_L g1010 ( 
.A(n_924),
.B(n_587),
.Y(n_1010)
);

HB1xp67_ASAP7_75t_L g1011 ( 
.A(n_900),
.Y(n_1011)
);

OAI21xp5_ASAP7_75t_L g1012 ( 
.A1(n_918),
.A2(n_652),
.B(n_201),
.Y(n_1012)
);

AOI21xp5_ASAP7_75t_L g1013 ( 
.A1(n_920),
.A2(n_432),
.B(n_183),
.Y(n_1013)
);

NAND2xp5_ASAP7_75t_L g1014 ( 
.A(n_925),
.B(n_652),
.Y(n_1014)
);

INVx4_ASAP7_75t_L g1015 ( 
.A(n_921),
.Y(n_1015)
);

AOI21xp5_ASAP7_75t_L g1016 ( 
.A1(n_901),
.A2(n_925),
.B(n_180),
.Y(n_1016)
);

NAND2x1p5_ASAP7_75t_L g1017 ( 
.A(n_901),
.B(n_502),
.Y(n_1017)
);

NOR2xp33_ASAP7_75t_L g1018 ( 
.A(n_913),
.B(n_195),
.Y(n_1018)
);

AO22x1_ASAP7_75t_L g1019 ( 
.A1(n_993),
.A2(n_652),
.B1(n_202),
.B2(n_209),
.Y(n_1019)
);

INVx1_ASAP7_75t_L g1020 ( 
.A(n_1002),
.Y(n_1020)
);

NAND2xp33_ASAP7_75t_SL g1021 ( 
.A(n_963),
.B(n_203),
.Y(n_1021)
);

INVx1_ASAP7_75t_L g1022 ( 
.A(n_1011),
.Y(n_1022)
);

AO22x1_ASAP7_75t_L g1023 ( 
.A1(n_959),
.A2(n_230),
.B1(n_180),
.B2(n_521),
.Y(n_1023)
);

CKINVDCx5p33_ASAP7_75t_R g1024 ( 
.A(n_1018),
.Y(n_1024)
);

BUFx2_ASAP7_75t_L g1025 ( 
.A(n_972),
.Y(n_1025)
);

NAND2xp5_ASAP7_75t_L g1026 ( 
.A(n_979),
.B(n_991),
.Y(n_1026)
);

INVx2_ASAP7_75t_L g1027 ( 
.A(n_969),
.Y(n_1027)
);

HB1xp67_ASAP7_75t_L g1028 ( 
.A(n_967),
.Y(n_1028)
);

INVx3_ASAP7_75t_L g1029 ( 
.A(n_1015),
.Y(n_1029)
);

NAND2xp5_ASAP7_75t_L g1030 ( 
.A(n_977),
.B(n_0),
.Y(n_1030)
);

OAI21xp33_ASAP7_75t_SL g1031 ( 
.A1(n_964),
.A2(n_965),
.B(n_980),
.Y(n_1031)
);

NAND2xp5_ASAP7_75t_SL g1032 ( 
.A(n_954),
.B(n_180),
.Y(n_1032)
);

INVx3_ASAP7_75t_L g1033 ( 
.A(n_1015),
.Y(n_1033)
);

NAND2xp5_ASAP7_75t_L g1034 ( 
.A(n_971),
.B(n_1),
.Y(n_1034)
);

OR2x6_ASAP7_75t_L g1035 ( 
.A(n_966),
.B(n_504),
.Y(n_1035)
);

BUFx3_ASAP7_75t_L g1036 ( 
.A(n_978),
.Y(n_1036)
);

NAND3xp33_ASAP7_75t_L g1037 ( 
.A(n_1032),
.B(n_1001),
.C(n_958),
.Y(n_1037)
);

INVx5_ASAP7_75t_L g1038 ( 
.A(n_1029),
.Y(n_1038)
);

AOI21xp5_ASAP7_75t_L g1039 ( 
.A1(n_1032),
.A2(n_986),
.B(n_1013),
.Y(n_1039)
);

AOI21xp5_ASAP7_75t_L g1040 ( 
.A1(n_1021),
.A2(n_1016),
.B(n_973),
.Y(n_1040)
);

BUFx6f_ASAP7_75t_L g1041 ( 
.A(n_1024),
.Y(n_1041)
);

NOR2x1_ASAP7_75t_L g1042 ( 
.A(n_1036),
.B(n_992),
.Y(n_1042)
);

BUFx2_ASAP7_75t_L g1043 ( 
.A(n_1025),
.Y(n_1043)
);

O2A1O1Ixp33_ASAP7_75t_L g1044 ( 
.A1(n_1026),
.A2(n_1031),
.B(n_1030),
.C(n_1034),
.Y(n_1044)
);

OAI22xp5_ASAP7_75t_L g1045 ( 
.A1(n_1035),
.A2(n_962),
.B1(n_990),
.B2(n_1007),
.Y(n_1045)
);

O2A1O1Ixp33_ASAP7_75t_L g1046 ( 
.A1(n_1035),
.A2(n_992),
.B(n_1009),
.C(n_984),
.Y(n_1046)
);

NAND2xp5_ASAP7_75t_L g1047 ( 
.A(n_1022),
.B(n_999),
.Y(n_1047)
);

OAI22xp5_ASAP7_75t_L g1048 ( 
.A1(n_1035),
.A2(n_970),
.B1(n_1005),
.B2(n_961),
.Y(n_1048)
);

OAI22xp5_ASAP7_75t_L g1049 ( 
.A1(n_1035),
.A2(n_987),
.B1(n_985),
.B2(n_978),
.Y(n_1049)
);

A2O1A1Ixp33_ASAP7_75t_L g1050 ( 
.A1(n_1021),
.A2(n_994),
.B(n_1000),
.C(n_1012),
.Y(n_1050)
);

AOI21x1_ASAP7_75t_L g1051 ( 
.A1(n_1023),
.A2(n_968),
.B(n_988),
.Y(n_1051)
);

OAI21xp5_ASAP7_75t_L g1052 ( 
.A1(n_1028),
.A2(n_1012),
.B(n_996),
.Y(n_1052)
);

INVx2_ASAP7_75t_L g1053 ( 
.A(n_1036),
.Y(n_1053)
);

A2O1A1Ixp33_ASAP7_75t_SL g1054 ( 
.A1(n_1027),
.A2(n_982),
.B(n_983),
.C(n_995),
.Y(n_1054)
);

O2A1O1Ixp33_ASAP7_75t_L g1055 ( 
.A1(n_1027),
.A2(n_1014),
.B(n_956),
.C(n_960),
.Y(n_1055)
);

AOI21xp5_ASAP7_75t_L g1056 ( 
.A1(n_1019),
.A2(n_983),
.B(n_974),
.Y(n_1056)
);

NOR2xp67_ASAP7_75t_SL g1057 ( 
.A(n_1024),
.B(n_978),
.Y(n_1057)
);

NOR2xp33_ASAP7_75t_L g1058 ( 
.A(n_1020),
.B(n_976),
.Y(n_1058)
);

AOI21xp5_ASAP7_75t_L g1059 ( 
.A1(n_1029),
.A2(n_1010),
.B(n_1008),
.Y(n_1059)
);

AOI21xp5_ASAP7_75t_L g1060 ( 
.A1(n_1029),
.A2(n_989),
.B(n_981),
.Y(n_1060)
);

OA22x2_ASAP7_75t_L g1061 ( 
.A1(n_1033),
.A2(n_998),
.B1(n_957),
.B2(n_1006),
.Y(n_1061)
);

OAI21x1_ASAP7_75t_L g1062 ( 
.A1(n_1042),
.A2(n_1033),
.B(n_998),
.Y(n_1062)
);

NAND2x1p5_ASAP7_75t_L g1063 ( 
.A(n_1057),
.B(n_1033),
.Y(n_1063)
);

BUFx2_ASAP7_75t_L g1064 ( 
.A(n_1043),
.Y(n_1064)
);

OAI21x1_ASAP7_75t_L g1065 ( 
.A1(n_1061),
.A2(n_1017),
.B(n_997),
.Y(n_1065)
);

AOI21xp5_ASAP7_75t_L g1066 ( 
.A1(n_1050),
.A2(n_1003),
.B(n_1017),
.Y(n_1066)
);

AO31x2_ASAP7_75t_L g1067 ( 
.A1(n_1053),
.A2(n_1004),
.A3(n_517),
.B(n_513),
.Y(n_1067)
);

AOI21x1_ASAP7_75t_L g1068 ( 
.A1(n_1051),
.A2(n_975),
.B(n_955),
.Y(n_1068)
);

BUFx6f_ASAP7_75t_L g1069 ( 
.A(n_1062),
.Y(n_1069)
);

INVx2_ASAP7_75t_SL g1070 ( 
.A(n_1064),
.Y(n_1070)
);

BUFx3_ASAP7_75t_L g1071 ( 
.A(n_1063),
.Y(n_1071)
);

AND2x2_ASAP7_75t_L g1072 ( 
.A(n_1071),
.B(n_1041),
.Y(n_1072)
);

NAND2xp33_ASAP7_75t_SL g1073 ( 
.A(n_1070),
.B(n_1041),
.Y(n_1073)
);

O2A1O1Ixp33_ASAP7_75t_L g1074 ( 
.A1(n_1070),
.A2(n_1054),
.B(n_1046),
.C(n_1037),
.Y(n_1074)
);

OA21x2_ASAP7_75t_L g1075 ( 
.A1(n_1072),
.A2(n_1068),
.B(n_1065),
.Y(n_1075)
);

INVx1_ASAP7_75t_L g1076 ( 
.A(n_1074),
.Y(n_1076)
);

BUFx2_ASAP7_75t_L g1077 ( 
.A(n_1075),
.Y(n_1077)
);

AOI22xp33_ASAP7_75t_SL g1078 ( 
.A1(n_1076),
.A2(n_1069),
.B1(n_1071),
.B2(n_1040),
.Y(n_1078)
);

OA21x2_ASAP7_75t_L g1079 ( 
.A1(n_1077),
.A2(n_1076),
.B(n_1068),
.Y(n_1079)
);

BUFx2_ASAP7_75t_SL g1080 ( 
.A(n_1078),
.Y(n_1080)
);

AND2x2_ASAP7_75t_L g1081 ( 
.A(n_1080),
.B(n_1038),
.Y(n_1081)
);

OAI22xp5_ASAP7_75t_L g1082 ( 
.A1(n_1079),
.A2(n_1069),
.B1(n_1044),
.B2(n_1038),
.Y(n_1082)
);

AOI22xp5_ASAP7_75t_L g1083 ( 
.A1(n_1081),
.A2(n_1073),
.B1(n_1079),
.B2(n_1069),
.Y(n_1083)
);

OAI21xp5_ASAP7_75t_SL g1084 ( 
.A1(n_1082),
.A2(n_1069),
.B(n_1039),
.Y(n_1084)
);

CKINVDCx10_ASAP7_75t_R g1085 ( 
.A(n_1083),
.Y(n_1085)
);

AOI221xp5_ASAP7_75t_L g1086 ( 
.A1(n_1084),
.A2(n_1069),
.B1(n_1066),
.B2(n_1048),
.C(n_1052),
.Y(n_1086)
);

NOR2xp33_ASAP7_75t_L g1087 ( 
.A(n_1085),
.B(n_1075),
.Y(n_1087)
);

OAI21xp5_ASAP7_75t_L g1088 ( 
.A1(n_1086),
.A2(n_1075),
.B(n_1047),
.Y(n_1088)
);

INVx2_ASAP7_75t_SL g1089 ( 
.A(n_1085),
.Y(n_1089)
);

INVx2_ASAP7_75t_SL g1090 ( 
.A(n_1089),
.Y(n_1090)
);

INVx2_ASAP7_75t_SL g1091 ( 
.A(n_1087),
.Y(n_1091)
);

AND2x4_ASAP7_75t_SL g1092 ( 
.A(n_1088),
.B(n_1058),
.Y(n_1092)
);

INVx1_ASAP7_75t_L g1093 ( 
.A(n_1090),
.Y(n_1093)
);

AND2x2_ASAP7_75t_L g1094 ( 
.A(n_1092),
.B(n_1075),
.Y(n_1094)
);

BUFx2_ASAP7_75t_L g1095 ( 
.A(n_1094),
.Y(n_1095)
);

INVx2_ASAP7_75t_L g1096 ( 
.A(n_1093),
.Y(n_1096)
);

AOI22xp5_ASAP7_75t_L g1097 ( 
.A1(n_1096),
.A2(n_1091),
.B1(n_1049),
.B2(n_1060),
.Y(n_1097)
);

OAI22xp33_ASAP7_75t_L g1098 ( 
.A1(n_1095),
.A2(n_1056),
.B1(n_1059),
.B2(n_1045),
.Y(n_1098)
);

INVx2_ASAP7_75t_L g1099 ( 
.A(n_1097),
.Y(n_1099)
);

HB1xp67_ASAP7_75t_L g1100 ( 
.A(n_1098),
.Y(n_1100)
);

AND2x4_ASAP7_75t_L g1101 ( 
.A(n_1099),
.B(n_1067),
.Y(n_1101)
);

AOI22xp33_ASAP7_75t_L g1102 ( 
.A1(n_1100),
.A2(n_180),
.B1(n_223),
.B2(n_226),
.Y(n_1102)
);

AND2x4_ASAP7_75t_SL g1103 ( 
.A(n_1102),
.B(n_489),
.Y(n_1103)
);

INVx1_ASAP7_75t_SL g1104 ( 
.A(n_1101),
.Y(n_1104)
);

OAI22xp5_ASAP7_75t_L g1105 ( 
.A1(n_1104),
.A2(n_1103),
.B1(n_1055),
.B2(n_227),
.Y(n_1105)
);

INVx2_ASAP7_75t_L g1106 ( 
.A(n_1103),
.Y(n_1106)
);

AND2x2_ASAP7_75t_L g1107 ( 
.A(n_1104),
.B(n_1067),
.Y(n_1107)
);

INVx2_ASAP7_75t_SL g1108 ( 
.A(n_1107),
.Y(n_1108)
);

INVxp67_ASAP7_75t_SL g1109 ( 
.A(n_1106),
.Y(n_1109)
);

NAND2xp5_ASAP7_75t_SL g1110 ( 
.A(n_1105),
.B(n_229),
.Y(n_1110)
);

OAI322xp33_ASAP7_75t_L g1111 ( 
.A1(n_1108),
.A2(n_2),
.A3(n_3),
.B1(n_4),
.B2(n_5),
.C1(n_6),
.C2(n_7),
.Y(n_1111)
);

AND2x4_ASAP7_75t_L g1112 ( 
.A(n_1109),
.B(n_1067),
.Y(n_1112)
);

INVx1_ASAP7_75t_SL g1113 ( 
.A(n_1111),
.Y(n_1113)
);

AOI221xp5_ASAP7_75t_L g1114 ( 
.A1(n_1112),
.A2(n_1110),
.B1(n_5),
.B2(n_7),
.C(n_8),
.Y(n_1114)
);

INVx1_ASAP7_75t_L g1115 ( 
.A(n_1113),
.Y(n_1115)
);

INVx1_ASAP7_75t_L g1116 ( 
.A(n_1114),
.Y(n_1116)
);

OR2x2_ASAP7_75t_L g1117 ( 
.A(n_1115),
.B(n_2),
.Y(n_1117)
);

BUFx3_ASAP7_75t_L g1118 ( 
.A(n_1116),
.Y(n_1118)
);

NAND2xp5_ASAP7_75t_L g1119 ( 
.A(n_1118),
.B(n_8),
.Y(n_1119)
);

AOI321xp33_ASAP7_75t_L g1120 ( 
.A1(n_1117),
.A2(n_9),
.A3(n_10),
.B1(n_11),
.B2(n_12),
.C(n_13),
.Y(n_1120)
);

INVx1_ASAP7_75t_L g1121 ( 
.A(n_1120),
.Y(n_1121)
);

OAI22xp5_ASAP7_75t_L g1122 ( 
.A1(n_1119),
.A2(n_9),
.B1(n_10),
.B2(n_11),
.Y(n_1122)
);

XNOR2xp5_ASAP7_75t_L g1123 ( 
.A(n_1121),
.B(n_12),
.Y(n_1123)
);

INVxp67_ASAP7_75t_L g1124 ( 
.A(n_1122),
.Y(n_1124)
);

INVx1_ASAP7_75t_L g1125 ( 
.A(n_1121),
.Y(n_1125)
);

XNOR2x1_ASAP7_75t_L g1126 ( 
.A(n_1125),
.B(n_14),
.Y(n_1126)
);

NOR2xp33_ASAP7_75t_L g1127 ( 
.A(n_1124),
.B(n_15),
.Y(n_1127)
);

AOI22xp33_ASAP7_75t_L g1128 ( 
.A1(n_1123),
.A2(n_16),
.B1(n_17),
.B2(n_19),
.Y(n_1128)
);

INVx1_ASAP7_75t_L g1129 ( 
.A(n_1126),
.Y(n_1129)
);

INVx1_ASAP7_75t_L g1130 ( 
.A(n_1128),
.Y(n_1130)
);

AND2x2_ASAP7_75t_L g1131 ( 
.A(n_1130),
.B(n_1127),
.Y(n_1131)
);

INVx1_ASAP7_75t_L g1132 ( 
.A(n_1129),
.Y(n_1132)
);

NOR2x1_ASAP7_75t_L g1133 ( 
.A(n_1132),
.B(n_338),
.Y(n_1133)
);

NOR2xp33_ASAP7_75t_SL g1134 ( 
.A(n_1131),
.B(n_16),
.Y(n_1134)
);

OAI21xp33_ASAP7_75t_L g1135 ( 
.A1(n_1133),
.A2(n_20),
.B(n_21),
.Y(n_1135)
);

AOI21xp33_ASAP7_75t_SL g1136 ( 
.A1(n_1134),
.A2(n_21),
.B(n_22),
.Y(n_1136)
);

NAND2xp5_ASAP7_75t_L g1137 ( 
.A(n_1136),
.B(n_23),
.Y(n_1137)
);

NOR2xp33_ASAP7_75t_L g1138 ( 
.A(n_1135),
.B(n_23),
.Y(n_1138)
);

INVx2_ASAP7_75t_L g1139 ( 
.A(n_1137),
.Y(n_1139)
);

INVx1_ASAP7_75t_L g1140 ( 
.A(n_1138),
.Y(n_1140)
);

AOI211xp5_ASAP7_75t_L g1141 ( 
.A1(n_1140),
.A2(n_24),
.B(n_25),
.C(n_26),
.Y(n_1141)
);

NAND3xp33_ASAP7_75t_SL g1142 ( 
.A(n_1139),
.B(n_24),
.C(n_27),
.Y(n_1142)
);

AOI211xp5_ASAP7_75t_L g1143 ( 
.A1(n_1140),
.A2(n_27),
.B(n_28),
.C(n_29),
.Y(n_1143)
);

INVx1_ASAP7_75t_L g1144 ( 
.A(n_1142),
.Y(n_1144)
);

OA22x2_ASAP7_75t_L g1145 ( 
.A1(n_1141),
.A2(n_28),
.B1(n_29),
.B2(n_30),
.Y(n_1145)
);

AOI221xp5_ASAP7_75t_L g1146 ( 
.A1(n_1143),
.A2(n_30),
.B1(n_31),
.B2(n_33),
.C(n_34),
.Y(n_1146)
);

OAI22xp5_ASAP7_75t_L g1147 ( 
.A1(n_1144),
.A2(n_33),
.B1(n_35),
.B2(n_36),
.Y(n_1147)
);

OAI21xp33_ASAP7_75t_L g1148 ( 
.A1(n_1145),
.A2(n_35),
.B(n_37),
.Y(n_1148)
);

NAND2xp5_ASAP7_75t_SL g1149 ( 
.A(n_1148),
.B(n_1146),
.Y(n_1149)
);

INVx1_ASAP7_75t_L g1150 ( 
.A(n_1147),
.Y(n_1150)
);

NOR3xp33_ASAP7_75t_L g1151 ( 
.A(n_1150),
.B(n_37),
.C(n_38),
.Y(n_1151)
);

AND2x4_ASAP7_75t_L g1152 ( 
.A(n_1149),
.B(n_38),
.Y(n_1152)
);

NOR3xp33_ASAP7_75t_L g1153 ( 
.A(n_1151),
.B(n_39),
.C(n_40),
.Y(n_1153)
);

NAND3xp33_ASAP7_75t_L g1154 ( 
.A(n_1152),
.B(n_491),
.C(n_41),
.Y(n_1154)
);

OR2x2_ASAP7_75t_L g1155 ( 
.A(n_1153),
.B(n_42),
.Y(n_1155)
);

INVx1_ASAP7_75t_L g1156 ( 
.A(n_1154),
.Y(n_1156)
);

OAI22xp33_ASAP7_75t_L g1157 ( 
.A1(n_1156),
.A2(n_43),
.B1(n_44),
.B2(n_47),
.Y(n_1157)
);

NAND2x1p5_ASAP7_75t_L g1158 ( 
.A(n_1155),
.B(n_486),
.Y(n_1158)
);

AND2x2_ASAP7_75t_L g1159 ( 
.A(n_1158),
.B(n_48),
.Y(n_1159)
);

OAI222xp33_ASAP7_75t_L g1160 ( 
.A1(n_1157),
.A2(n_49),
.B1(n_50),
.B2(n_51),
.C1(n_52),
.C2(n_53),
.Y(n_1160)
);

OAI221xp5_ASAP7_75t_L g1161 ( 
.A1(n_1158),
.A2(n_54),
.B1(n_56),
.B2(n_57),
.C(n_58),
.Y(n_1161)
);

OA22x2_ASAP7_75t_L g1162 ( 
.A1(n_1159),
.A2(n_59),
.B1(n_60),
.B2(n_61),
.Y(n_1162)
);

HB1xp67_ASAP7_75t_L g1163 ( 
.A(n_1160),
.Y(n_1163)
);

HB1xp67_ASAP7_75t_L g1164 ( 
.A(n_1161),
.Y(n_1164)
);

AOI221xp5_ASAP7_75t_L g1165 ( 
.A1(n_1163),
.A2(n_486),
.B1(n_489),
.B2(n_64),
.C(n_65),
.Y(n_1165)
);

AOI22xp33_ASAP7_75t_L g1166 ( 
.A1(n_1164),
.A2(n_1162),
.B1(n_486),
.B2(n_489),
.Y(n_1166)
);

INVx2_ASAP7_75t_L g1167 ( 
.A(n_1166),
.Y(n_1167)
);

INVx1_ASAP7_75t_L g1168 ( 
.A(n_1165),
.Y(n_1168)
);

INVx1_ASAP7_75t_SL g1169 ( 
.A(n_1168),
.Y(n_1169)
);

INVx1_ASAP7_75t_L g1170 ( 
.A(n_1167),
.Y(n_1170)
);

NAND2xp5_ASAP7_75t_L g1171 ( 
.A(n_1170),
.B(n_62),
.Y(n_1171)
);

AOI22xp5_ASAP7_75t_L g1172 ( 
.A1(n_1169),
.A2(n_496),
.B1(n_511),
.B2(n_484),
.Y(n_1172)
);

AOI22xp33_ASAP7_75t_L g1173 ( 
.A1(n_1171),
.A2(n_490),
.B1(n_485),
.B2(n_484),
.Y(n_1173)
);

OAI22xp5_ASAP7_75t_L g1174 ( 
.A1(n_1172),
.A2(n_511),
.B1(n_496),
.B2(n_490),
.Y(n_1174)
);

XNOR2x1_ASAP7_75t_L g1175 ( 
.A(n_1174),
.B(n_63),
.Y(n_1175)
);

NAND3xp33_ASAP7_75t_L g1176 ( 
.A(n_1173),
.B(n_66),
.C(n_67),
.Y(n_1176)
);

INVx2_ASAP7_75t_L g1177 ( 
.A(n_1175),
.Y(n_1177)
);

AO21x2_ASAP7_75t_L g1178 ( 
.A1(n_1176),
.A2(n_69),
.B(n_71),
.Y(n_1178)
);

INVx1_ASAP7_75t_L g1179 ( 
.A(n_1175),
.Y(n_1179)
);

INVx1_ASAP7_75t_L g1180 ( 
.A(n_1175),
.Y(n_1180)
);

AOI221xp5_ASAP7_75t_L g1181 ( 
.A1(n_1179),
.A2(n_72),
.B1(n_74),
.B2(n_75),
.C(n_78),
.Y(n_1181)
);

OAI21xp5_ASAP7_75t_L g1182 ( 
.A1(n_1180),
.A2(n_511),
.B(n_496),
.Y(n_1182)
);

AOI22xp5_ASAP7_75t_L g1183 ( 
.A1(n_1177),
.A2(n_511),
.B1(n_490),
.B2(n_485),
.Y(n_1183)
);

OR2x2_ASAP7_75t_SL g1184 ( 
.A(n_1178),
.B(n_80),
.Y(n_1184)
);

INVx2_ASAP7_75t_L g1185 ( 
.A(n_1184),
.Y(n_1185)
);

INVx1_ASAP7_75t_L g1186 ( 
.A(n_1182),
.Y(n_1186)
);

CKINVDCx20_ASAP7_75t_R g1187 ( 
.A(n_1181),
.Y(n_1187)
);

AOI22xp5_ASAP7_75t_L g1188 ( 
.A1(n_1187),
.A2(n_1183),
.B1(n_490),
.B2(n_485),
.Y(n_1188)
);

OAI21xp5_ASAP7_75t_SL g1189 ( 
.A1(n_1185),
.A2(n_81),
.B(n_82),
.Y(n_1189)
);

OAI21xp5_ASAP7_75t_L g1190 ( 
.A1(n_1186),
.A2(n_83),
.B(n_86),
.Y(n_1190)
);

AOI22xp5_ASAP7_75t_L g1191 ( 
.A1(n_1187),
.A2(n_490),
.B1(n_485),
.B2(n_484),
.Y(n_1191)
);

OAI21xp5_ASAP7_75t_L g1192 ( 
.A1(n_1187),
.A2(n_87),
.B(n_88),
.Y(n_1192)
);

OAI21xp5_ASAP7_75t_L g1193 ( 
.A1(n_1187),
.A2(n_89),
.B(n_90),
.Y(n_1193)
);

INVx1_ASAP7_75t_L g1194 ( 
.A(n_1187),
.Y(n_1194)
);

OA21x2_ASAP7_75t_L g1195 ( 
.A1(n_1185),
.A2(n_93),
.B(n_94),
.Y(n_1195)
);

OA22x2_ASAP7_75t_L g1196 ( 
.A1(n_1185),
.A2(n_95),
.B1(n_96),
.B2(n_97),
.Y(n_1196)
);

AOI21xp5_ASAP7_75t_L g1197 ( 
.A1(n_1187),
.A2(n_98),
.B(n_101),
.Y(n_1197)
);

AOI22xp5_ASAP7_75t_L g1198 ( 
.A1(n_1187),
.A2(n_485),
.B1(n_484),
.B2(n_483),
.Y(n_1198)
);

NOR2xp33_ASAP7_75t_L g1199 ( 
.A(n_1187),
.B(n_105),
.Y(n_1199)
);

NAND2xp5_ASAP7_75t_L g1200 ( 
.A(n_1194),
.B(n_107),
.Y(n_1200)
);

NAND4xp25_ASAP7_75t_L g1201 ( 
.A(n_1197),
.B(n_108),
.C(n_109),
.D(n_111),
.Y(n_1201)
);

XNOR2xp5_ASAP7_75t_L g1202 ( 
.A(n_1195),
.B(n_112),
.Y(n_1202)
);

OAI22xp5_ASAP7_75t_L g1203 ( 
.A1(n_1188),
.A2(n_113),
.B1(n_115),
.B2(n_117),
.Y(n_1203)
);

OAI22xp5_ASAP7_75t_SL g1204 ( 
.A1(n_1199),
.A2(n_118),
.B1(n_120),
.B2(n_121),
.Y(n_1204)
);

AOI22xp33_ASAP7_75t_L g1205 ( 
.A1(n_1196),
.A2(n_124),
.B1(n_125),
.B2(n_126),
.Y(n_1205)
);

XNOR2xp5_ASAP7_75t_L g1206 ( 
.A(n_1189),
.B(n_127),
.Y(n_1206)
);

XNOR2xp5_ASAP7_75t_L g1207 ( 
.A(n_1190),
.B(n_128),
.Y(n_1207)
);

XNOR2xp5_ASAP7_75t_L g1208 ( 
.A(n_1192),
.B(n_129),
.Y(n_1208)
);

INVx2_ASAP7_75t_L g1209 ( 
.A(n_1202),
.Y(n_1209)
);

AOI21xp5_ASAP7_75t_L g1210 ( 
.A1(n_1206),
.A2(n_1207),
.B(n_1208),
.Y(n_1210)
);

OR2x2_ASAP7_75t_L g1211 ( 
.A(n_1205),
.B(n_1201),
.Y(n_1211)
);

NAND2xp5_ASAP7_75t_L g1212 ( 
.A(n_1204),
.B(n_1193),
.Y(n_1212)
);

AOI21xp5_ASAP7_75t_L g1213 ( 
.A1(n_1200),
.A2(n_1198),
.B(n_1191),
.Y(n_1213)
);

AOI221xp5_ASAP7_75t_L g1214 ( 
.A1(n_1203),
.A2(n_130),
.B1(n_131),
.B2(n_132),
.C(n_133),
.Y(n_1214)
);

AOI222xp33_ASAP7_75t_L g1215 ( 
.A1(n_1202),
.A2(n_135),
.B1(n_136),
.B2(n_137),
.C1(n_138),
.C2(n_139),
.Y(n_1215)
);

OAI21xp5_ASAP7_75t_L g1216 ( 
.A1(n_1212),
.A2(n_140),
.B(n_141),
.Y(n_1216)
);

OAI21xp5_ASAP7_75t_L g1217 ( 
.A1(n_1210),
.A2(n_142),
.B(n_143),
.Y(n_1217)
);

NAND3xp33_ASAP7_75t_L g1218 ( 
.A(n_1209),
.B(n_144),
.C(n_146),
.Y(n_1218)
);

AOI222xp33_ASAP7_75t_SL g1219 ( 
.A1(n_1217),
.A2(n_1211),
.B1(n_1213),
.B2(n_1214),
.C1(n_1215),
.C2(n_151),
.Y(n_1219)
);

NAND2xp5_ASAP7_75t_L g1220 ( 
.A(n_1219),
.B(n_1218),
.Y(n_1220)
);

INVx1_ASAP7_75t_L g1221 ( 
.A(n_1220),
.Y(n_1221)
);

INVx1_ASAP7_75t_L g1222 ( 
.A(n_1221),
.Y(n_1222)
);

OR2x6_ASAP7_75t_L g1223 ( 
.A(n_1222),
.B(n_1216),
.Y(n_1223)
);

OAI221xp5_ASAP7_75t_R g1224 ( 
.A1(n_1223),
.A2(n_147),
.B1(n_148),
.B2(n_149),
.C(n_150),
.Y(n_1224)
);

AOI22xp5_ASAP7_75t_L g1225 ( 
.A1(n_1224),
.A2(n_153),
.B1(n_154),
.B2(n_157),
.Y(n_1225)
);

AOI22xp33_ASAP7_75t_L g1226 ( 
.A1(n_1225),
.A2(n_158),
.B1(n_159),
.B2(n_162),
.Y(n_1226)
);

AOI211xp5_ASAP7_75t_L g1227 ( 
.A1(n_1226),
.A2(n_163),
.B(n_165),
.C(n_166),
.Y(n_1227)
);

AOI211xp5_ASAP7_75t_L g1228 ( 
.A1(n_1227),
.A2(n_167),
.B(n_169),
.C(n_172),
.Y(n_1228)
);


endmodule