module fake_jpeg_2632_n_550 (n_13, n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_550);

input n_13;
input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_550;

wire n_529;
wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_525;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_16;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_15;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_519;
wire n_276;
wire n_143;
wire n_17;
wire n_431;
wire n_102;
wire n_549;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_172;
wire n_547;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_513;
wire n_283;
wire n_107;
wire n_490;
wire n_517;
wire n_415;
wire n_479;
wire n_543;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_542;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_48;
wire n_465;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_256;
wire n_221;
wire n_454;
wire n_540;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_508;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_544;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_530;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_298;
wire n_106;
wire n_545;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_474;
wire n_539;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_511;
wire n_305;
wire n_161;
wire n_441;
wire n_342;
wire n_101;
wire n_226;
wire n_509;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_510;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_536;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_14;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_537;
wire n_110;
wire n_531;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_523;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_533;
wire n_296;
wire n_384;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_491;
wire n_24;
wire n_526;
wire n_467;
wire n_269;
wire n_546;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_473;
wire n_45;
wire n_520;
wire n_476;
wire n_337;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_344;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_481;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_522;
wire n_333;
wire n_518;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_302;
wire n_216;
wire n_528;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_199;
wire n_260;
wire n_413;
wire n_275;
wire n_494;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_492;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_515;
wire n_347;
wire n_521;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_538;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_534;
wire n_472;
wire n_279;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_484;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_469;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_527;
wire n_482;
wire n_58;
wire n_41;
wire n_266;
wire n_548;
wire n_72;
wire n_512;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_516;
wire n_183;
wire n_409;
wire n_532;
wire n_412;
wire n_249;
wire n_217;
wire n_471;
wire n_541;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_535;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_524;
wire n_402;
wire n_504;
wire n_438;
wire n_475;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_514;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

BUFx5_ASAP7_75t_L g14 ( 
.A(n_10),
.Y(n_14)
);

INVx1_ASAP7_75t_L g15 ( 
.A(n_8),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_9),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_6),
.Y(n_17)
);

INVx11_ASAP7_75t_L g18 ( 
.A(n_2),
.Y(n_18)
);

INVx2_ASAP7_75t_SL g19 ( 
.A(n_7),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_9),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_3),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_13),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_1),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_9),
.Y(n_24)
);

BUFx3_ASAP7_75t_L g25 ( 
.A(n_9),
.Y(n_25)
);

BUFx5_ASAP7_75t_L g26 ( 
.A(n_0),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_12),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_0),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_5),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_13),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_6),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_10),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_7),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_13),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_7),
.Y(n_35)
);

INVx2_ASAP7_75t_L g36 ( 
.A(n_13),
.Y(n_36)
);

INVxp67_ASAP7_75t_L g37 ( 
.A(n_0),
.Y(n_37)
);

INVx8_ASAP7_75t_L g38 ( 
.A(n_5),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_13),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_11),
.Y(n_40)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_4),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_4),
.Y(n_42)
);

BUFx5_ASAP7_75t_L g43 ( 
.A(n_2),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_0),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_5),
.Y(n_45)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_6),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_SL g47 ( 
.A(n_21),
.B(n_0),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g134 ( 
.A(n_47),
.B(n_77),
.Y(n_134)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_22),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g108 ( 
.A(n_48),
.Y(n_108)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_22),
.Y(n_49)
);

INVx6_ASAP7_75t_L g116 ( 
.A(n_49),
.Y(n_116)
);

INVx5_ASAP7_75t_L g50 ( 
.A(n_38),
.Y(n_50)
);

BUFx3_ASAP7_75t_L g155 ( 
.A(n_50),
.Y(n_155)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_22),
.Y(n_51)
);

INVx6_ASAP7_75t_L g145 ( 
.A(n_51),
.Y(n_145)
);

INVx3_ASAP7_75t_L g52 ( 
.A(n_25),
.Y(n_52)
);

INVx2_ASAP7_75t_SL g110 ( 
.A(n_52),
.Y(n_110)
);

INVx8_ASAP7_75t_L g53 ( 
.A(n_22),
.Y(n_53)
);

BUFx2_ASAP7_75t_L g114 ( 
.A(n_53),
.Y(n_114)
);

BUFx3_ASAP7_75t_L g54 ( 
.A(n_25),
.Y(n_54)
);

BUFx2_ASAP7_75t_L g126 ( 
.A(n_54),
.Y(n_126)
);

INVx13_ASAP7_75t_L g55 ( 
.A(n_37),
.Y(n_55)
);

INVx1_ASAP7_75t_SL g136 ( 
.A(n_55),
.Y(n_136)
);

INVx3_ASAP7_75t_L g56 ( 
.A(n_25),
.Y(n_56)
);

INVx2_ASAP7_75t_SL g123 ( 
.A(n_56),
.Y(n_123)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_36),
.Y(n_57)
);

INVx2_ASAP7_75t_L g120 ( 
.A(n_57),
.Y(n_120)
);

INVx11_ASAP7_75t_L g58 ( 
.A(n_26),
.Y(n_58)
);

INVx4_ASAP7_75t_L g109 ( 
.A(n_58),
.Y(n_109)
);

INVx2_ASAP7_75t_L g59 ( 
.A(n_36),
.Y(n_59)
);

INVx2_ASAP7_75t_L g125 ( 
.A(n_59),
.Y(n_125)
);

INVx3_ASAP7_75t_L g60 ( 
.A(n_38),
.Y(n_60)
);

INVx2_ASAP7_75t_SL g156 ( 
.A(n_60),
.Y(n_156)
);

INVx6_ASAP7_75t_L g61 ( 
.A(n_44),
.Y(n_61)
);

INVx3_ASAP7_75t_SL g107 ( 
.A(n_61),
.Y(n_107)
);

INVx3_ASAP7_75t_L g62 ( 
.A(n_38),
.Y(n_62)
);

INVx3_ASAP7_75t_L g119 ( 
.A(n_62),
.Y(n_119)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_23),
.Y(n_63)
);

INVx6_ASAP7_75t_L g148 ( 
.A(n_63),
.Y(n_148)
);

INVx11_ASAP7_75t_L g64 ( 
.A(n_26),
.Y(n_64)
);

INVx4_ASAP7_75t_L g127 ( 
.A(n_64),
.Y(n_127)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_23),
.Y(n_65)
);

INVx3_ASAP7_75t_SL g140 ( 
.A(n_65),
.Y(n_140)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_36),
.Y(n_66)
);

INVx2_ASAP7_75t_L g130 ( 
.A(n_66),
.Y(n_130)
);

INVx2_ASAP7_75t_L g67 ( 
.A(n_44),
.Y(n_67)
);

INVx2_ASAP7_75t_L g131 ( 
.A(n_67),
.Y(n_131)
);

INVx5_ASAP7_75t_L g68 ( 
.A(n_38),
.Y(n_68)
);

INVx4_ASAP7_75t_L g137 ( 
.A(n_68),
.Y(n_137)
);

INVx3_ASAP7_75t_L g69 ( 
.A(n_44),
.Y(n_69)
);

INVx3_ASAP7_75t_L g133 ( 
.A(n_69),
.Y(n_133)
);

INVx5_ASAP7_75t_L g70 ( 
.A(n_44),
.Y(n_70)
);

INVx4_ASAP7_75t_L g160 ( 
.A(n_70),
.Y(n_160)
);

INVx2_ASAP7_75t_L g71 ( 
.A(n_26),
.Y(n_71)
);

INVx2_ASAP7_75t_L g132 ( 
.A(n_71),
.Y(n_132)
);

INVx5_ASAP7_75t_L g72 ( 
.A(n_23),
.Y(n_72)
);

INVx4_ASAP7_75t_L g104 ( 
.A(n_72),
.Y(n_104)
);

BUFx6f_ASAP7_75t_L g73 ( 
.A(n_23),
.Y(n_73)
);

INVx3_ASAP7_75t_SL g153 ( 
.A(n_73),
.Y(n_153)
);

BUFx6f_ASAP7_75t_L g74 ( 
.A(n_31),
.Y(n_74)
);

INVx8_ASAP7_75t_L g111 ( 
.A(n_74),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_21),
.B(n_0),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_L g105 ( 
.A(n_75),
.B(n_89),
.Y(n_105)
);

INVx6_ASAP7_75t_L g76 ( 
.A(n_31),
.Y(n_76)
);

INVx8_ASAP7_75t_L g135 ( 
.A(n_76),
.Y(n_135)
);

CKINVDCx16_ASAP7_75t_R g77 ( 
.A(n_31),
.Y(n_77)
);

BUFx6f_ASAP7_75t_L g78 ( 
.A(n_31),
.Y(n_78)
);

INVx8_ASAP7_75t_L g167 ( 
.A(n_78),
.Y(n_167)
);

BUFx3_ASAP7_75t_L g79 ( 
.A(n_34),
.Y(n_79)
);

INVx5_ASAP7_75t_L g112 ( 
.A(n_79),
.Y(n_112)
);

BUFx3_ASAP7_75t_L g80 ( 
.A(n_34),
.Y(n_80)
);

INVx5_ASAP7_75t_L g122 ( 
.A(n_80),
.Y(n_122)
);

BUFx6f_ASAP7_75t_L g81 ( 
.A(n_34),
.Y(n_81)
);

BUFx12f_ASAP7_75t_L g157 ( 
.A(n_81),
.Y(n_157)
);

INVx2_ASAP7_75t_L g82 ( 
.A(n_34),
.Y(n_82)
);

INVx2_ASAP7_75t_L g150 ( 
.A(n_82),
.Y(n_150)
);

INVx2_ASAP7_75t_SL g83 ( 
.A(n_19),
.Y(n_83)
);

INVx4_ASAP7_75t_L g113 ( 
.A(n_83),
.Y(n_113)
);

INVx2_ASAP7_75t_L g84 ( 
.A(n_40),
.Y(n_84)
);

INVx2_ASAP7_75t_L g151 ( 
.A(n_84),
.Y(n_151)
);

INVx4_ASAP7_75t_L g85 ( 
.A(n_14),
.Y(n_85)
);

INVx3_ASAP7_75t_L g143 ( 
.A(n_85),
.Y(n_143)
);

BUFx3_ASAP7_75t_L g86 ( 
.A(n_40),
.Y(n_86)
);

INVx5_ASAP7_75t_L g124 ( 
.A(n_86),
.Y(n_124)
);

INVx3_ASAP7_75t_L g87 ( 
.A(n_40),
.Y(n_87)
);

INVx3_ASAP7_75t_L g152 ( 
.A(n_87),
.Y(n_152)
);

INVx8_ASAP7_75t_L g88 ( 
.A(n_40),
.Y(n_88)
);

INVx5_ASAP7_75t_L g158 ( 
.A(n_88),
.Y(n_158)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_28),
.B(n_1),
.Y(n_89)
);

INVx2_ASAP7_75t_L g90 ( 
.A(n_42),
.Y(n_90)
);

INVx2_ASAP7_75t_L g154 ( 
.A(n_90),
.Y(n_154)
);

INVx3_ASAP7_75t_L g91 ( 
.A(n_42),
.Y(n_91)
);

INVx3_ASAP7_75t_L g165 ( 
.A(n_91),
.Y(n_165)
);

BUFx6f_ASAP7_75t_L g92 ( 
.A(n_42),
.Y(n_92)
);

INVx5_ASAP7_75t_L g163 ( 
.A(n_92),
.Y(n_163)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_28),
.B(n_39),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_L g118 ( 
.A(n_93),
.B(n_94),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_SL g94 ( 
.A(n_28),
.B(n_1),
.Y(n_94)
);

INVx2_ASAP7_75t_L g95 ( 
.A(n_42),
.Y(n_95)
);

INVx2_ASAP7_75t_L g161 ( 
.A(n_95),
.Y(n_161)
);

INVx2_ASAP7_75t_L g96 ( 
.A(n_14),
.Y(n_96)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_96),
.Y(n_115)
);

INVx11_ASAP7_75t_L g97 ( 
.A(n_14),
.Y(n_97)
);

INVx4_ASAP7_75t_L g117 ( 
.A(n_97),
.Y(n_117)
);

INVx3_ASAP7_75t_L g98 ( 
.A(n_15),
.Y(n_98)
);

INVx4_ASAP7_75t_L g166 ( 
.A(n_98),
.Y(n_166)
);

BUFx6f_ASAP7_75t_L g99 ( 
.A(n_15),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g144 ( 
.A(n_99),
.B(n_101),
.Y(n_144)
);

INVx8_ASAP7_75t_L g100 ( 
.A(n_43),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g164 ( 
.A(n_100),
.B(n_102),
.Y(n_164)
);

BUFx6f_ASAP7_75t_L g101 ( 
.A(n_15),
.Y(n_101)
);

BUFx12_ASAP7_75t_L g102 ( 
.A(n_43),
.Y(n_102)
);

AOI21xp5_ASAP7_75t_L g103 ( 
.A1(n_85),
.A2(n_83),
.B(n_19),
.Y(n_103)
);

AOI21xp5_ASAP7_75t_L g203 ( 
.A1(n_103),
.A2(n_46),
.B(n_33),
.Y(n_203)
);

AOI22xp33_ASAP7_75t_SL g106 ( 
.A1(n_97),
.A2(n_19),
.B1(n_18),
.B2(n_39),
.Y(n_106)
);

OA22x2_ASAP7_75t_L g175 ( 
.A1(n_106),
.A2(n_129),
.B1(n_162),
.B2(n_30),
.Y(n_175)
);

OAI22xp5_ASAP7_75t_SL g121 ( 
.A1(n_76),
.A2(n_39),
.B1(n_45),
.B2(n_20),
.Y(n_121)
);

AOI22xp5_ASAP7_75t_SL g213 ( 
.A1(n_121),
.A2(n_146),
.B1(n_159),
.B2(n_27),
.Y(n_213)
);

AOI22xp33_ASAP7_75t_L g128 ( 
.A1(n_48),
.A2(n_19),
.B1(n_45),
.B2(n_35),
.Y(n_128)
);

OAI22xp5_ASAP7_75t_L g197 ( 
.A1(n_128),
.A2(n_139),
.B1(n_142),
.B2(n_149),
.Y(n_197)
);

AOI22xp33_ASAP7_75t_SL g129 ( 
.A1(n_58),
.A2(n_18),
.B1(n_45),
.B2(n_35),
.Y(n_129)
);

OAI21xp5_ASAP7_75t_L g138 ( 
.A1(n_54),
.A2(n_17),
.B(n_35),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_L g182 ( 
.A(n_138),
.B(n_30),
.Y(n_182)
);

OAI22xp5_ASAP7_75t_L g139 ( 
.A1(n_61),
.A2(n_65),
.B1(n_49),
.B2(n_73),
.Y(n_139)
);

OR2x2_ASAP7_75t_L g141 ( 
.A(n_55),
.B(n_41),
.Y(n_141)
);

CKINVDCx14_ASAP7_75t_R g190 ( 
.A(n_141),
.Y(n_190)
);

AOI22xp5_ASAP7_75t_L g142 ( 
.A1(n_51),
.A2(n_16),
.B1(n_29),
.B2(n_24),
.Y(n_142)
);

OAI22xp5_ASAP7_75t_SL g146 ( 
.A1(n_63),
.A2(n_16),
.B1(n_29),
.B2(n_24),
.Y(n_146)
);

OR2x2_ASAP7_75t_L g147 ( 
.A(n_99),
.B(n_41),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_SL g194 ( 
.A(n_147),
.B(n_46),
.Y(n_194)
);

AOI22xp33_ASAP7_75t_L g149 ( 
.A1(n_74),
.A2(n_16),
.B1(n_29),
.B2(n_24),
.Y(n_149)
);

OAI22xp33_ASAP7_75t_SL g159 ( 
.A1(n_78),
.A2(n_17),
.B1(n_20),
.B2(n_18),
.Y(n_159)
);

AOI22xp33_ASAP7_75t_SL g162 ( 
.A1(n_64),
.A2(n_17),
.B1(n_20),
.B2(n_41),
.Y(n_162)
);

OAI22xp5_ASAP7_75t_SL g168 ( 
.A1(n_149),
.A2(n_92),
.B1(n_81),
.B2(n_79),
.Y(n_168)
);

OAI22xp5_ASAP7_75t_L g237 ( 
.A1(n_168),
.A2(n_198),
.B1(n_214),
.B2(n_216),
.Y(n_237)
);

AND2x2_ASAP7_75t_SL g169 ( 
.A(n_144),
.B(n_70),
.Y(n_169)
);

NOR2xp33_ASAP7_75t_L g217 ( 
.A(n_169),
.B(n_173),
.Y(n_217)
);

INVx3_ASAP7_75t_L g170 ( 
.A(n_113),
.Y(n_170)
);

INVx3_ASAP7_75t_L g220 ( 
.A(n_170),
.Y(n_220)
);

NAND2xp33_ASAP7_75t_SL g171 ( 
.A(n_147),
.B(n_101),
.Y(n_171)
);

OR2x2_ASAP7_75t_L g225 ( 
.A(n_171),
.B(n_174),
.Y(n_225)
);

INVx3_ASAP7_75t_L g172 ( 
.A(n_160),
.Y(n_172)
);

INVx3_ASAP7_75t_L g240 ( 
.A(n_172),
.Y(n_240)
);

CKINVDCx16_ASAP7_75t_R g173 ( 
.A(n_141),
.Y(n_173)
);

INVx5_ASAP7_75t_SL g174 ( 
.A(n_136),
.Y(n_174)
);

OA22x2_ASAP7_75t_L g247 ( 
.A1(n_175),
.A2(n_186),
.B1(n_213),
.B2(n_145),
.Y(n_247)
);

INVx8_ASAP7_75t_L g176 ( 
.A(n_157),
.Y(n_176)
);

BUFx3_ASAP7_75t_L g228 ( 
.A(n_176),
.Y(n_228)
);

CKINVDCx20_ASAP7_75t_R g177 ( 
.A(n_114),
.Y(n_177)
);

NOR2xp33_ASAP7_75t_SL g218 ( 
.A(n_177),
.B(n_185),
.Y(n_218)
);

INVx3_ASAP7_75t_L g178 ( 
.A(n_160),
.Y(n_178)
);

INVx2_ASAP7_75t_SL g245 ( 
.A(n_178),
.Y(n_245)
);

BUFx12f_ASAP7_75t_L g179 ( 
.A(n_143),
.Y(n_179)
);

INVx11_ASAP7_75t_L g224 ( 
.A(n_179),
.Y(n_224)
);

CKINVDCx16_ASAP7_75t_R g180 ( 
.A(n_164),
.Y(n_180)
);

NOR2xp33_ASAP7_75t_L g229 ( 
.A(n_180),
.B(n_193),
.Y(n_229)
);

INVx2_ASAP7_75t_L g181 ( 
.A(n_131),
.Y(n_181)
);

INVx2_ASAP7_75t_L g246 ( 
.A(n_181),
.Y(n_246)
);

NAND3xp33_ASAP7_75t_L g235 ( 
.A(n_182),
.B(n_194),
.C(n_206),
.Y(n_235)
);

INVx2_ASAP7_75t_L g183 ( 
.A(n_150),
.Y(n_183)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_183),
.Y(n_223)
);

INVx4_ASAP7_75t_L g184 ( 
.A(n_137),
.Y(n_184)
);

BUFx6f_ASAP7_75t_L g219 ( 
.A(n_184),
.Y(n_219)
);

CKINVDCx20_ASAP7_75t_R g185 ( 
.A(n_114),
.Y(n_185)
);

AO22x2_ASAP7_75t_L g186 ( 
.A1(n_128),
.A2(n_72),
.B1(n_50),
.B2(n_68),
.Y(n_186)
);

BUFx12f_ASAP7_75t_L g187 ( 
.A(n_111),
.Y(n_187)
);

BUFx6f_ASAP7_75t_L g221 ( 
.A(n_187),
.Y(n_221)
);

INVx5_ASAP7_75t_L g188 ( 
.A(n_111),
.Y(n_188)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_188),
.Y(n_244)
);

INVx8_ASAP7_75t_L g189 ( 
.A(n_157),
.Y(n_189)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_189),
.Y(n_254)
);

OAI22xp33_ASAP7_75t_SL g191 ( 
.A1(n_134),
.A2(n_80),
.B1(n_86),
.B2(n_30),
.Y(n_191)
);

AOI22xp33_ASAP7_75t_L g234 ( 
.A1(n_191),
.A2(n_140),
.B1(n_153),
.B2(n_163),
.Y(n_234)
);

BUFx2_ASAP7_75t_L g192 ( 
.A(n_126),
.Y(n_192)
);

CKINVDCx20_ASAP7_75t_R g222 ( 
.A(n_192),
.Y(n_222)
);

INVx2_ASAP7_75t_L g193 ( 
.A(n_151),
.Y(n_193)
);

INVx2_ASAP7_75t_L g195 ( 
.A(n_154),
.Y(n_195)
);

NOR2xp33_ASAP7_75t_L g242 ( 
.A(n_195),
.B(n_199),
.Y(n_242)
);

INVx6_ASAP7_75t_L g196 ( 
.A(n_108),
.Y(n_196)
);

CKINVDCx20_ASAP7_75t_R g248 ( 
.A(n_196),
.Y(n_248)
);

AOI22xp33_ASAP7_75t_SL g198 ( 
.A1(n_105),
.A2(n_46),
.B1(n_32),
.B2(n_33),
.Y(n_198)
);

INVx3_ASAP7_75t_L g199 ( 
.A(n_104),
.Y(n_199)
);

INVx5_ASAP7_75t_L g200 ( 
.A(n_167),
.Y(n_200)
);

CKINVDCx20_ASAP7_75t_R g251 ( 
.A(n_200),
.Y(n_251)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_159),
.Y(n_201)
);

OR2x2_ASAP7_75t_L g239 ( 
.A(n_201),
.B(n_205),
.Y(n_239)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_110),
.Y(n_202)
);

NOR2xp33_ASAP7_75t_L g243 ( 
.A(n_202),
.B(n_204),
.Y(n_243)
);

AOI21xp5_ASAP7_75t_L g236 ( 
.A1(n_203),
.A2(n_127),
.B(n_109),
.Y(n_236)
);

INVx2_ASAP7_75t_L g204 ( 
.A(n_161),
.Y(n_204)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_133),
.Y(n_205)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_107),
.Y(n_206)
);

BUFx6f_ASAP7_75t_L g207 ( 
.A(n_108),
.Y(n_207)
);

BUFx12_ASAP7_75t_L g249 ( 
.A(n_207),
.Y(n_249)
);

NAND2xp5_ASAP7_75t_L g208 ( 
.A(n_118),
.B(n_33),
.Y(n_208)
);

NAND2xp5_ASAP7_75t_L g230 ( 
.A(n_208),
.B(n_212),
.Y(n_230)
);

AND2x2_ASAP7_75t_L g209 ( 
.A(n_166),
.B(n_32),
.Y(n_209)
);

NOR2xp33_ASAP7_75t_SL g232 ( 
.A(n_209),
.B(n_210),
.Y(n_232)
);

CKINVDCx20_ASAP7_75t_R g210 ( 
.A(n_126),
.Y(n_210)
);

NOR2xp33_ASAP7_75t_SL g211 ( 
.A(n_115),
.B(n_32),
.Y(n_211)
);

NAND2xp5_ASAP7_75t_SL g233 ( 
.A(n_211),
.B(n_208),
.Y(n_233)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_110),
.Y(n_212)
);

OAI22xp5_ASAP7_75t_L g214 ( 
.A1(n_162),
.A2(n_129),
.B1(n_106),
.B2(n_116),
.Y(n_214)
);

NAND2xp5_ASAP7_75t_L g215 ( 
.A(n_120),
.B(n_27),
.Y(n_215)
);

NAND2xp5_ASAP7_75t_L g231 ( 
.A(n_215),
.B(n_123),
.Y(n_231)
);

AOI22xp33_ASAP7_75t_SL g216 ( 
.A1(n_123),
.A2(n_27),
.B1(n_100),
.B2(n_156),
.Y(n_216)
);

OA22x2_ASAP7_75t_SL g226 ( 
.A1(n_171),
.A2(n_107),
.B1(n_156),
.B2(n_140),
.Y(n_226)
);

CKINVDCx20_ASAP7_75t_R g261 ( 
.A(n_226),
.Y(n_261)
);

OAI22xp5_ASAP7_75t_SL g227 ( 
.A1(n_201),
.A2(n_119),
.B1(n_125),
.B2(n_130),
.Y(n_227)
);

AOI22xp5_ASAP7_75t_L g280 ( 
.A1(n_227),
.A2(n_241),
.B1(n_250),
.B2(n_252),
.Y(n_280)
);

NAND2xp5_ASAP7_75t_SL g273 ( 
.A(n_231),
.B(n_186),
.Y(n_273)
);

NOR2xp33_ASAP7_75t_SL g267 ( 
.A(n_233),
.B(n_209),
.Y(n_267)
);

OR2x2_ASAP7_75t_L g275 ( 
.A(n_234),
.B(n_236),
.Y(n_275)
);

NAND2xp5_ASAP7_75t_L g238 ( 
.A(n_215),
.B(n_132),
.Y(n_238)
);

NAND2xp5_ASAP7_75t_L g266 ( 
.A(n_238),
.B(n_253),
.Y(n_266)
);

OAI22xp5_ASAP7_75t_L g241 ( 
.A1(n_197),
.A2(n_148),
.B1(n_116),
.B2(n_145),
.Y(n_241)
);

AOI22xp33_ASAP7_75t_SL g260 ( 
.A1(n_247),
.A2(n_175),
.B1(n_168),
.B2(n_186),
.Y(n_260)
);

OAI22xp5_ASAP7_75t_L g250 ( 
.A1(n_213),
.A2(n_148),
.B1(n_135),
.B2(n_167),
.Y(n_250)
);

OAI22xp5_ASAP7_75t_SL g252 ( 
.A1(n_169),
.A2(n_165),
.B1(n_152),
.B2(n_153),
.Y(n_252)
);

NAND2xp5_ASAP7_75t_L g253 ( 
.A(n_169),
.B(n_158),
.Y(n_253)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_242),
.Y(n_255)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_255),
.Y(n_288)
);

INVx2_ASAP7_75t_L g256 ( 
.A(n_245),
.Y(n_256)
);

INVx1_ASAP7_75t_SL g304 ( 
.A(n_256),
.Y(n_304)
);

NAND2xp5_ASAP7_75t_L g257 ( 
.A(n_238),
.B(n_203),
.Y(n_257)
);

NAND2xp5_ASAP7_75t_L g307 ( 
.A(n_257),
.B(n_268),
.Y(n_307)
);

NOR2xp33_ASAP7_75t_L g258 ( 
.A(n_229),
.B(n_190),
.Y(n_258)
);

NOR2xp33_ASAP7_75t_SL g316 ( 
.A(n_258),
.B(n_259),
.Y(n_316)
);

NOR2xp33_ASAP7_75t_L g259 ( 
.A(n_229),
.B(n_205),
.Y(n_259)
);

OAI22xp5_ASAP7_75t_SL g294 ( 
.A1(n_260),
.A2(n_247),
.B1(n_225),
.B2(n_239),
.Y(n_294)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_242),
.Y(n_262)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_262),
.Y(n_306)
);

OAI22xp5_ASAP7_75t_SL g263 ( 
.A1(n_239),
.A2(n_175),
.B1(n_186),
.B2(n_135),
.Y(n_263)
);

AOI22xp5_ASAP7_75t_L g300 ( 
.A1(n_263),
.A2(n_270),
.B1(n_261),
.B2(n_275),
.Y(n_300)
);

CKINVDCx20_ASAP7_75t_R g264 ( 
.A(n_218),
.Y(n_264)
);

NOR2xp33_ASAP7_75t_L g293 ( 
.A(n_264),
.B(n_269),
.Y(n_293)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_243),
.Y(n_265)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_265),
.Y(n_310)
);

NAND2xp5_ASAP7_75t_SL g286 ( 
.A(n_267),
.B(n_273),
.Y(n_286)
);

NOR2xp33_ASAP7_75t_L g268 ( 
.A(n_218),
.B(n_170),
.Y(n_268)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_243),
.Y(n_269)
);

OAI21xp5_ASAP7_75t_L g270 ( 
.A1(n_236),
.A2(n_175),
.B(n_209),
.Y(n_270)
);

OAI21xp5_ASAP7_75t_L g298 ( 
.A1(n_270),
.A2(n_283),
.B(n_285),
.Y(n_298)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_223),
.Y(n_271)
);

NOR2xp33_ASAP7_75t_L g296 ( 
.A(n_271),
.B(n_276),
.Y(n_296)
);

NAND2xp5_ASAP7_75t_L g272 ( 
.A(n_230),
.B(n_183),
.Y(n_272)
);

NAND2xp5_ASAP7_75t_L g315 ( 
.A(n_272),
.B(n_274),
.Y(n_315)
);

NAND2xp5_ASAP7_75t_SL g274 ( 
.A(n_230),
.B(n_181),
.Y(n_274)
);

CKINVDCx20_ASAP7_75t_R g276 ( 
.A(n_239),
.Y(n_276)
);

NOR2xp33_ASAP7_75t_L g277 ( 
.A(n_235),
.B(n_204),
.Y(n_277)
);

NOR2xp33_ASAP7_75t_L g303 ( 
.A(n_277),
.B(n_279),
.Y(n_303)
);

OAI32xp33_ASAP7_75t_L g278 ( 
.A1(n_231),
.A2(n_206),
.A3(n_195),
.B1(n_193),
.B2(n_188),
.Y(n_278)
);

INVxp67_ASAP7_75t_L g291 ( 
.A(n_278),
.Y(n_291)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_223),
.Y(n_279)
);

AOI22xp33_ASAP7_75t_SL g281 ( 
.A1(n_237),
.A2(n_192),
.B1(n_187),
.B2(n_200),
.Y(n_281)
);

OAI22x1_ASAP7_75t_L g289 ( 
.A1(n_281),
.A2(n_226),
.B1(n_187),
.B2(n_244),
.Y(n_289)
);

MAJIxp5_ASAP7_75t_L g282 ( 
.A(n_217),
.B(n_184),
.C(n_172),
.Y(n_282)
);

MAJIxp5_ASAP7_75t_L g301 ( 
.A(n_282),
.B(n_284),
.C(n_252),
.Y(n_301)
);

AOI21xp5_ASAP7_75t_SL g283 ( 
.A1(n_217),
.A2(n_174),
.B(n_102),
.Y(n_283)
);

XNOR2xp5_ASAP7_75t_L g284 ( 
.A(n_233),
.B(n_178),
.Y(n_284)
);

NOR2xp33_ASAP7_75t_L g285 ( 
.A(n_235),
.B(n_199),
.Y(n_285)
);

XNOR2xp5_ASAP7_75t_L g287 ( 
.A(n_284),
.B(n_253),
.Y(n_287)
);

XNOR2xp5_ASAP7_75t_SL g337 ( 
.A(n_287),
.B(n_299),
.Y(n_337)
);

AOI22xp5_ASAP7_75t_L g327 ( 
.A1(n_289),
.A2(n_294),
.B1(n_295),
.B2(n_300),
.Y(n_327)
);

CKINVDCx20_ASAP7_75t_R g290 ( 
.A(n_268),
.Y(n_290)
);

NOR2xp33_ASAP7_75t_L g318 ( 
.A(n_290),
.B(n_305),
.Y(n_318)
);

XOR2xp5_ASAP7_75t_L g292 ( 
.A(n_284),
.B(n_266),
.Y(n_292)
);

MAJIxp5_ASAP7_75t_L g328 ( 
.A(n_292),
.B(n_308),
.C(n_255),
.Y(n_328)
);

OAI22xp5_ASAP7_75t_SL g295 ( 
.A1(n_260),
.A2(n_247),
.B1(n_225),
.B2(n_241),
.Y(n_295)
);

AOI21xp5_ASAP7_75t_L g297 ( 
.A1(n_270),
.A2(n_225),
.B(n_237),
.Y(n_297)
);

AOI21xp5_ASAP7_75t_L g344 ( 
.A1(n_297),
.A2(n_245),
.B(n_254),
.Y(n_344)
);

XNOR2xp5_ASAP7_75t_L g299 ( 
.A(n_267),
.B(n_232),
.Y(n_299)
);

XOR2xp5_ASAP7_75t_L g347 ( 
.A(n_301),
.B(n_287),
.Y(n_347)
);

OAI22xp5_ASAP7_75t_SL g302 ( 
.A1(n_261),
.A2(n_247),
.B1(n_250),
.B2(n_226),
.Y(n_302)
);

AOI22xp5_ASAP7_75t_L g330 ( 
.A1(n_302),
.A2(n_309),
.B1(n_312),
.B2(n_313),
.Y(n_330)
);

CKINVDCx20_ASAP7_75t_R g305 ( 
.A(n_259),
.Y(n_305)
);

XNOR2xp5_ASAP7_75t_L g308 ( 
.A(n_266),
.B(n_272),
.Y(n_308)
);

OAI22xp5_ASAP7_75t_SL g309 ( 
.A1(n_257),
.A2(n_247),
.B1(n_226),
.B2(n_227),
.Y(n_309)
);

A2O1A1Ixp33_ASAP7_75t_L g311 ( 
.A1(n_257),
.A2(n_232),
.B(n_251),
.C(n_222),
.Y(n_311)
);

NAND2xp5_ASAP7_75t_L g326 ( 
.A(n_311),
.B(n_263),
.Y(n_326)
);

OAI22xp5_ASAP7_75t_SL g312 ( 
.A1(n_273),
.A2(n_248),
.B1(n_251),
.B2(n_196),
.Y(n_312)
);

OAI22xp5_ASAP7_75t_SL g313 ( 
.A1(n_275),
.A2(n_248),
.B1(n_244),
.B2(n_207),
.Y(n_313)
);

OAI22xp5_ASAP7_75t_SL g314 ( 
.A1(n_275),
.A2(n_245),
.B1(n_222),
.B2(n_240),
.Y(n_314)
);

AOI22xp5_ASAP7_75t_L g348 ( 
.A1(n_314),
.A2(n_302),
.B1(n_309),
.B2(n_313),
.Y(n_348)
);

OAI21xp5_ASAP7_75t_L g317 ( 
.A1(n_276),
.A2(n_245),
.B(n_254),
.Y(n_317)
);

OAI21xp5_ASAP7_75t_SL g319 ( 
.A1(n_317),
.A2(n_283),
.B(n_275),
.Y(n_319)
);

OAI21xp5_ASAP7_75t_SL g351 ( 
.A1(n_319),
.A2(n_320),
.B(n_321),
.Y(n_351)
);

OAI21xp5_ASAP7_75t_SL g320 ( 
.A1(n_298),
.A2(n_283),
.B(n_285),
.Y(n_320)
);

AOI21xp5_ASAP7_75t_SL g321 ( 
.A1(n_298),
.A2(n_277),
.B(n_258),
.Y(n_321)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_288),
.Y(n_322)
);

INVx1_ASAP7_75t_L g362 ( 
.A(n_322),
.Y(n_362)
);

INVx2_ASAP7_75t_L g323 ( 
.A(n_288),
.Y(n_323)
);

INVx2_ASAP7_75t_L g364 ( 
.A(n_323),
.Y(n_364)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_306),
.Y(n_324)
);

INVx1_ASAP7_75t_L g353 ( 
.A(n_324),
.Y(n_353)
);

INVxp33_ASAP7_75t_L g325 ( 
.A(n_293),
.Y(n_325)
);

NOR2xp33_ASAP7_75t_L g365 ( 
.A(n_325),
.B(n_316),
.Y(n_365)
);

OAI21xp5_ASAP7_75t_L g358 ( 
.A1(n_326),
.A2(n_341),
.B(n_344),
.Y(n_358)
);

XNOR2xp5_ASAP7_75t_L g360 ( 
.A(n_328),
.B(n_299),
.Y(n_360)
);

XNOR2xp5_ASAP7_75t_L g329 ( 
.A(n_292),
.B(n_282),
.Y(n_329)
);

MAJIxp5_ASAP7_75t_L g359 ( 
.A(n_329),
.B(n_347),
.C(n_286),
.Y(n_359)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_306),
.Y(n_331)
);

INVx1_ASAP7_75t_L g354 ( 
.A(n_331),
.Y(n_354)
);

AOI22x1_ASAP7_75t_SL g332 ( 
.A1(n_294),
.A2(n_263),
.B1(n_262),
.B2(n_269),
.Y(n_332)
);

OAI22xp5_ASAP7_75t_L g355 ( 
.A1(n_332),
.A2(n_345),
.B1(n_348),
.B2(n_317),
.Y(n_355)
);

AND2x2_ASAP7_75t_L g333 ( 
.A(n_297),
.B(n_278),
.Y(n_333)
);

AND2x2_ASAP7_75t_L g383 ( 
.A(n_333),
.B(n_220),
.Y(n_383)
);

OAI22xp5_ASAP7_75t_SL g334 ( 
.A1(n_300),
.A2(n_280),
.B1(n_281),
.B2(n_265),
.Y(n_334)
);

AOI22xp5_ASAP7_75t_L g357 ( 
.A1(n_334),
.A2(n_335),
.B1(n_339),
.B2(n_311),
.Y(n_357)
);

OAI22xp5_ASAP7_75t_SL g335 ( 
.A1(n_291),
.A2(n_280),
.B1(n_264),
.B2(n_274),
.Y(n_335)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_310),
.Y(n_336)
);

INVx1_ASAP7_75t_L g361 ( 
.A(n_336),
.Y(n_361)
);

CKINVDCx20_ASAP7_75t_R g338 ( 
.A(n_293),
.Y(n_338)
);

NAND2xp5_ASAP7_75t_L g356 ( 
.A(n_338),
.B(n_305),
.Y(n_356)
);

OAI22xp5_ASAP7_75t_SL g339 ( 
.A1(n_307),
.A2(n_280),
.B1(n_278),
.B2(n_282),
.Y(n_339)
);

NAND2xp5_ASAP7_75t_L g340 ( 
.A(n_296),
.B(n_279),
.Y(n_340)
);

INVx1_ASAP7_75t_L g363 ( 
.A(n_340),
.Y(n_363)
);

OAI21xp5_ASAP7_75t_L g341 ( 
.A1(n_311),
.A2(n_271),
.B(n_256),
.Y(n_341)
);

NAND2xp5_ASAP7_75t_L g342 ( 
.A(n_296),
.B(n_256),
.Y(n_342)
);

INVx1_ASAP7_75t_L g366 ( 
.A(n_342),
.Y(n_366)
);

INVx1_ASAP7_75t_L g343 ( 
.A(n_310),
.Y(n_343)
);

INVx1_ASAP7_75t_L g367 ( 
.A(n_343),
.Y(n_367)
);

OAI22xp5_ASAP7_75t_L g345 ( 
.A1(n_301),
.A2(n_228),
.B1(n_240),
.B2(n_221),
.Y(n_345)
);

INVx1_ASAP7_75t_L g346 ( 
.A(n_312),
.Y(n_346)
);

INVx1_ASAP7_75t_L g368 ( 
.A(n_346),
.Y(n_368)
);

NOR2xp33_ASAP7_75t_L g349 ( 
.A(n_316),
.B(n_240),
.Y(n_349)
);

NAND2xp5_ASAP7_75t_SL g371 ( 
.A(n_349),
.B(n_314),
.Y(n_371)
);

INVx1_ASAP7_75t_L g350 ( 
.A(n_315),
.Y(n_350)
);

INVx1_ASAP7_75t_L g369 ( 
.A(n_350),
.Y(n_369)
);

AOI22xp5_ASAP7_75t_SL g352 ( 
.A1(n_334),
.A2(n_295),
.B1(n_289),
.B2(n_290),
.Y(n_352)
);

OAI22xp5_ASAP7_75t_L g401 ( 
.A1(n_352),
.A2(n_357),
.B1(n_372),
.B2(n_333),
.Y(n_401)
);

AOI22xp5_ASAP7_75t_L g410 ( 
.A1(n_355),
.A2(n_374),
.B1(n_379),
.B2(n_221),
.Y(n_410)
);

INVx1_ASAP7_75t_L g384 ( 
.A(n_356),
.Y(n_384)
);

MAJIxp5_ASAP7_75t_L g387 ( 
.A(n_359),
.B(n_370),
.C(n_321),
.Y(n_387)
);

XOR2xp5_ASAP7_75t_L g414 ( 
.A(n_360),
.B(n_376),
.Y(n_414)
);

INVx1_ASAP7_75t_L g389 ( 
.A(n_365),
.Y(n_389)
);

MAJIxp5_ASAP7_75t_L g370 ( 
.A(n_347),
.B(n_308),
.C(n_307),
.Y(n_370)
);

INVx1_ASAP7_75t_L g405 ( 
.A(n_371),
.Y(n_405)
);

AOI22xp5_ASAP7_75t_L g372 ( 
.A1(n_335),
.A2(n_286),
.B1(n_289),
.B2(n_303),
.Y(n_372)
);

CKINVDCx20_ASAP7_75t_R g373 ( 
.A(n_340),
.Y(n_373)
);

NAND2xp5_ASAP7_75t_SL g406 ( 
.A(n_373),
.B(n_377),
.Y(n_406)
);

OAI22xp5_ASAP7_75t_SL g374 ( 
.A1(n_348),
.A2(n_330),
.B1(n_327),
.B2(n_346),
.Y(n_374)
);

NAND2xp5_ASAP7_75t_L g375 ( 
.A(n_338),
.B(n_315),
.Y(n_375)
);

INVx1_ASAP7_75t_L g413 ( 
.A(n_375),
.Y(n_413)
);

XNOR2xp5_ASAP7_75t_SL g376 ( 
.A(n_337),
.B(n_303),
.Y(n_376)
);

CKINVDCx20_ASAP7_75t_R g377 ( 
.A(n_318),
.Y(n_377)
);

INVx2_ASAP7_75t_L g378 ( 
.A(n_323),
.Y(n_378)
);

INVx2_ASAP7_75t_L g396 ( 
.A(n_378),
.Y(n_396)
);

OAI22xp5_ASAP7_75t_SL g379 ( 
.A1(n_330),
.A2(n_304),
.B1(n_221),
.B2(n_228),
.Y(n_379)
);

INVx1_ASAP7_75t_L g380 ( 
.A(n_322),
.Y(n_380)
);

BUFx2_ASAP7_75t_L g398 ( 
.A(n_380),
.Y(n_398)
);

NAND2xp5_ASAP7_75t_L g381 ( 
.A(n_318),
.B(n_304),
.Y(n_381)
);

NAND2xp5_ASAP7_75t_L g388 ( 
.A(n_381),
.B(n_382),
.Y(n_388)
);

NAND2xp5_ASAP7_75t_L g382 ( 
.A(n_350),
.B(n_304),
.Y(n_382)
);

OAI21xp5_ASAP7_75t_L g395 ( 
.A1(n_383),
.A2(n_344),
.B(n_319),
.Y(n_395)
);

CKINVDCx20_ASAP7_75t_R g385 ( 
.A(n_382),
.Y(n_385)
);

NAND2xp5_ASAP7_75t_L g417 ( 
.A(n_385),
.B(n_391),
.Y(n_417)
);

INVxp67_ASAP7_75t_L g386 ( 
.A(n_383),
.Y(n_386)
);

INVx1_ASAP7_75t_L g415 ( 
.A(n_386),
.Y(n_415)
);

XNOR2xp5_ASAP7_75t_L g421 ( 
.A(n_387),
.B(n_402),
.Y(n_421)
);

MAJIxp5_ASAP7_75t_L g390 ( 
.A(n_359),
.B(n_329),
.C(n_328),
.Y(n_390)
);

MAJIxp5_ASAP7_75t_L g424 ( 
.A(n_390),
.B(n_392),
.C(n_351),
.Y(n_424)
);

NOR2xp33_ASAP7_75t_L g391 ( 
.A(n_370),
.B(n_349),
.Y(n_391)
);

MAJIxp5_ASAP7_75t_L g392 ( 
.A(n_360),
.B(n_337),
.C(n_345),
.Y(n_392)
);

AOI21xp5_ASAP7_75t_L g393 ( 
.A1(n_358),
.A2(n_341),
.B(n_326),
.Y(n_393)
);

INVxp67_ASAP7_75t_L g416 ( 
.A(n_393),
.Y(n_416)
);

CKINVDCx20_ASAP7_75t_R g394 ( 
.A(n_381),
.Y(n_394)
);

NAND2xp5_ASAP7_75t_L g420 ( 
.A(n_394),
.B(n_395),
.Y(n_420)
);

NOR2xp33_ASAP7_75t_L g397 ( 
.A(n_356),
.B(n_363),
.Y(n_397)
);

NAND2xp5_ASAP7_75t_L g436 ( 
.A(n_397),
.B(n_403),
.Y(n_436)
);

OAI22xp5_ASAP7_75t_SL g399 ( 
.A1(n_357),
.A2(n_327),
.B1(n_333),
.B2(n_332),
.Y(n_399)
);

AOI22xp5_ASAP7_75t_L g418 ( 
.A1(n_399),
.A2(n_401),
.B1(n_374),
.B2(n_368),
.Y(n_418)
);

BUFx12_ASAP7_75t_L g400 ( 
.A(n_364),
.Y(n_400)
);

CKINVDCx20_ASAP7_75t_R g419 ( 
.A(n_400),
.Y(n_419)
);

XNOR2xp5_ASAP7_75t_L g402 ( 
.A(n_376),
.B(n_320),
.Y(n_402)
);

CKINVDCx20_ASAP7_75t_R g403 ( 
.A(n_375),
.Y(n_403)
);

OAI21xp5_ASAP7_75t_L g404 ( 
.A1(n_358),
.A2(n_339),
.B(n_342),
.Y(n_404)
);

NAND2xp5_ASAP7_75t_L g440 ( 
.A(n_404),
.B(n_407),
.Y(n_440)
);

NOR2xp33_ASAP7_75t_L g407 ( 
.A(n_363),
.B(n_343),
.Y(n_407)
);

OAI22xp5_ASAP7_75t_L g408 ( 
.A1(n_352),
.A2(n_336),
.B1(n_331),
.B2(n_324),
.Y(n_408)
);

OAI22xp5_ASAP7_75t_L g430 ( 
.A1(n_408),
.A2(n_410),
.B1(n_412),
.B2(n_361),
.Y(n_430)
);

O2A1O1Ixp33_ASAP7_75t_L g409 ( 
.A1(n_368),
.A2(n_228),
.B(n_246),
.C(n_224),
.Y(n_409)
);

INVx1_ASAP7_75t_L g435 ( 
.A(n_409),
.Y(n_435)
);

NOR2xp33_ASAP7_75t_L g411 ( 
.A(n_369),
.B(n_372),
.Y(n_411)
);

NOR2xp33_ASAP7_75t_L g425 ( 
.A(n_411),
.B(n_364),
.Y(n_425)
);

CKINVDCx20_ASAP7_75t_R g412 ( 
.A(n_383),
.Y(n_412)
);

OAI22xp5_ASAP7_75t_SL g460 ( 
.A1(n_418),
.A2(n_388),
.B1(n_396),
.B2(n_409),
.Y(n_460)
);

XNOR2xp5_ASAP7_75t_L g422 ( 
.A(n_390),
.B(n_351),
.Y(n_422)
);

XNOR2xp5_ASAP7_75t_L g453 ( 
.A(n_422),
.B(n_424),
.Y(n_453)
);

OAI22xp5_ASAP7_75t_SL g423 ( 
.A1(n_389),
.A2(n_369),
.B1(n_366),
.B2(n_380),
.Y(n_423)
);

HB1xp67_ASAP7_75t_L g455 ( 
.A(n_423),
.Y(n_455)
);

INVxp67_ASAP7_75t_L g442 ( 
.A(n_425),
.Y(n_442)
);

FAx1_ASAP7_75t_SL g426 ( 
.A(n_399),
.B(n_402),
.CI(n_404),
.CON(n_426),
.SN(n_426)
);

NAND2xp5_ASAP7_75t_L g446 ( 
.A(n_426),
.B(n_394),
.Y(n_446)
);

XNOR2xp5_ASAP7_75t_L g427 ( 
.A(n_387),
.B(n_366),
.Y(n_427)
);

XNOR2xp5_ASAP7_75t_L g462 ( 
.A(n_427),
.B(n_400),
.Y(n_462)
);

AOI22xp5_ASAP7_75t_L g428 ( 
.A1(n_384),
.A2(n_379),
.B1(n_353),
.B2(n_367),
.Y(n_428)
);

OAI22xp5_ASAP7_75t_L g461 ( 
.A1(n_428),
.A2(n_439),
.B1(n_396),
.B2(n_224),
.Y(n_461)
);

MAJIxp5_ASAP7_75t_L g429 ( 
.A(n_392),
.B(n_378),
.C(n_367),
.Y(n_429)
);

NAND2xp5_ASAP7_75t_SL g457 ( 
.A(n_429),
.B(n_431),
.Y(n_457)
);

AOI22xp5_ASAP7_75t_L g452 ( 
.A1(n_430),
.A2(n_438),
.B1(n_398),
.B2(n_413),
.Y(n_452)
);

MAJIxp5_ASAP7_75t_L g431 ( 
.A(n_414),
.B(n_361),
.C(n_354),
.Y(n_431)
);

NOR2xp33_ASAP7_75t_L g432 ( 
.A(n_389),
.B(n_362),
.Y(n_432)
);

INVx1_ASAP7_75t_L g448 ( 
.A(n_432),
.Y(n_448)
);

MAJIxp5_ASAP7_75t_L g433 ( 
.A(n_414),
.B(n_354),
.C(n_353),
.Y(n_433)
);

MAJIxp5_ASAP7_75t_L g444 ( 
.A(n_433),
.B(n_434),
.C(n_437),
.Y(n_444)
);

MAJIxp5_ASAP7_75t_L g434 ( 
.A(n_393),
.B(n_219),
.C(n_246),
.Y(n_434)
);

MAJIxp5_ASAP7_75t_L g437 ( 
.A(n_384),
.B(n_219),
.C(n_220),
.Y(n_437)
);

OAI22xp5_ASAP7_75t_SL g438 ( 
.A1(n_410),
.A2(n_220),
.B1(n_219),
.B2(n_189),
.Y(n_438)
);

AOI22xp5_ASAP7_75t_L g439 ( 
.A1(n_408),
.A2(n_176),
.B1(n_137),
.B2(n_112),
.Y(n_439)
);

MAJIxp5_ASAP7_75t_L g441 ( 
.A(n_395),
.B(n_155),
.C(n_109),
.Y(n_441)
);

MAJIxp5_ASAP7_75t_L g449 ( 
.A(n_441),
.B(n_398),
.C(n_386),
.Y(n_449)
);

NOR2xp33_ASAP7_75t_L g443 ( 
.A(n_427),
.B(n_406),
.Y(n_443)
);

NAND2xp5_ASAP7_75t_L g477 ( 
.A(n_443),
.B(n_445),
.Y(n_477)
);

NOR2xp33_ASAP7_75t_L g445 ( 
.A(n_429),
.B(n_405),
.Y(n_445)
);

OAI21xp5_ASAP7_75t_L g469 ( 
.A1(n_446),
.A2(n_416),
.B(n_421),
.Y(n_469)
);

NAND2xp5_ASAP7_75t_L g447 ( 
.A(n_417),
.B(n_403),
.Y(n_447)
);

INVx1_ASAP7_75t_L g468 ( 
.A(n_447),
.Y(n_468)
);

XNOR2xp5_ASAP7_75t_L g484 ( 
.A(n_449),
.B(n_462),
.Y(n_484)
);

CKINVDCx20_ASAP7_75t_R g450 ( 
.A(n_436),
.Y(n_450)
);

NOR2xp33_ASAP7_75t_L g483 ( 
.A(n_450),
.B(n_456),
.Y(n_483)
);

MAJIxp5_ASAP7_75t_L g451 ( 
.A(n_422),
.B(n_412),
.C(n_385),
.Y(n_451)
);

MAJIxp5_ASAP7_75t_L g465 ( 
.A(n_451),
.B(n_454),
.C(n_458),
.Y(n_465)
);

OAI22xp5_ASAP7_75t_L g466 ( 
.A1(n_452),
.A2(n_418),
.B1(n_451),
.B2(n_428),
.Y(n_466)
);

MAJIxp5_ASAP7_75t_L g454 ( 
.A(n_424),
.B(n_405),
.C(n_413),
.Y(n_454)
);

CKINVDCx20_ASAP7_75t_R g456 ( 
.A(n_420),
.Y(n_456)
);

MAJIxp5_ASAP7_75t_L g458 ( 
.A(n_431),
.B(n_388),
.C(n_398),
.Y(n_458)
);

INVx1_ASAP7_75t_L g459 ( 
.A(n_415),
.Y(n_459)
);

INVx1_ASAP7_75t_L g478 ( 
.A(n_459),
.Y(n_478)
);

AOI22xp5_ASAP7_75t_L g470 ( 
.A1(n_460),
.A2(n_461),
.B1(n_438),
.B2(n_435),
.Y(n_470)
);

CKINVDCx16_ASAP7_75t_R g463 ( 
.A(n_440),
.Y(n_463)
);

INVxp67_ASAP7_75t_SL g476 ( 
.A(n_463),
.Y(n_476)
);

XOR2xp5_ASAP7_75t_L g464 ( 
.A(n_433),
.B(n_400),
.Y(n_464)
);

XOR2xp5_ASAP7_75t_L g481 ( 
.A(n_464),
.B(n_224),
.Y(n_481)
);

INVx1_ASAP7_75t_L g488 ( 
.A(n_466),
.Y(n_488)
);

MAJIxp5_ASAP7_75t_L g467 ( 
.A(n_453),
.B(n_421),
.C(n_416),
.Y(n_467)
);

XNOR2xp5_ASAP7_75t_L g498 ( 
.A(n_467),
.B(n_471),
.Y(n_498)
);

INVx1_ASAP7_75t_L g489 ( 
.A(n_469),
.Y(n_489)
);

OAI22xp33_ASAP7_75t_L g500 ( 
.A1(n_470),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_500)
);

MAJIxp5_ASAP7_75t_L g471 ( 
.A(n_453),
.B(n_434),
.C(n_437),
.Y(n_471)
);

MAJIxp5_ASAP7_75t_L g472 ( 
.A(n_457),
.B(n_441),
.C(n_419),
.Y(n_472)
);

MAJIxp5_ASAP7_75t_L g486 ( 
.A(n_472),
.B(n_474),
.C(n_482),
.Y(n_486)
);

AOI21xp5_ASAP7_75t_L g473 ( 
.A1(n_454),
.A2(n_426),
.B(n_439),
.Y(n_473)
);

AOI21xp5_ASAP7_75t_L g497 ( 
.A1(n_473),
.A2(n_479),
.B(n_249),
.Y(n_497)
);

MAJIxp5_ASAP7_75t_L g474 ( 
.A(n_464),
.B(n_426),
.C(n_400),
.Y(n_474)
);

AOI22xp5_ASAP7_75t_L g475 ( 
.A1(n_455),
.A2(n_124),
.B1(n_122),
.B2(n_53),
.Y(n_475)
);

OAI22xp5_ASAP7_75t_L g491 ( 
.A1(n_475),
.A2(n_442),
.B1(n_470),
.B2(n_452),
.Y(n_491)
);

AOI21xp5_ASAP7_75t_L g479 ( 
.A1(n_446),
.A2(n_127),
.B(n_117),
.Y(n_479)
);

OAI22xp5_ASAP7_75t_SL g480 ( 
.A1(n_447),
.A2(n_155),
.B1(n_179),
.B2(n_157),
.Y(n_480)
);

XNOR2xp5_ASAP7_75t_L g493 ( 
.A(n_480),
.B(n_481),
.Y(n_493)
);

MAJIxp5_ASAP7_75t_L g482 ( 
.A(n_444),
.B(n_249),
.C(n_88),
.Y(n_482)
);

MAJIxp5_ASAP7_75t_L g485 ( 
.A(n_444),
.B(n_249),
.C(n_179),
.Y(n_485)
);

MAJIxp5_ASAP7_75t_L g487 ( 
.A(n_485),
.B(n_458),
.C(n_462),
.Y(n_487)
);

XOR2xp5_ASAP7_75t_L g513 ( 
.A(n_487),
.B(n_497),
.Y(n_513)
);

NOR2xp33_ASAP7_75t_L g490 ( 
.A(n_465),
.B(n_448),
.Y(n_490)
);

NAND2xp5_ASAP7_75t_L g507 ( 
.A(n_490),
.B(n_492),
.Y(n_507)
);

AOI22xp5_ASAP7_75t_L g508 ( 
.A1(n_491),
.A2(n_500),
.B1(n_480),
.B2(n_478),
.Y(n_508)
);

MAJIxp5_ASAP7_75t_L g492 ( 
.A(n_465),
.B(n_449),
.C(n_460),
.Y(n_492)
);

NOR2xp33_ASAP7_75t_L g494 ( 
.A(n_472),
.B(n_442),
.Y(n_494)
);

NAND2xp5_ASAP7_75t_L g517 ( 
.A(n_494),
.B(n_495),
.Y(n_517)
);

MAJIxp5_ASAP7_75t_L g495 ( 
.A(n_484),
.B(n_467),
.C(n_471),
.Y(n_495)
);

NOR2xp33_ASAP7_75t_L g496 ( 
.A(n_484),
.B(n_249),
.Y(n_496)
);

NAND2xp5_ASAP7_75t_SL g518 ( 
.A(n_496),
.B(n_499),
.Y(n_518)
);

MAJIxp5_ASAP7_75t_L g499 ( 
.A(n_474),
.B(n_102),
.C(n_43),
.Y(n_499)
);

NOR2xp33_ASAP7_75t_L g501 ( 
.A(n_477),
.B(n_1),
.Y(n_501)
);

AOI21xp5_ASAP7_75t_L g515 ( 
.A1(n_501),
.A2(n_502),
.B(n_4),
.Y(n_515)
);

NOR2xp33_ASAP7_75t_L g502 ( 
.A(n_483),
.B(n_12),
.Y(n_502)
);

MAJIxp5_ASAP7_75t_L g503 ( 
.A(n_481),
.B(n_2),
.C(n_3),
.Y(n_503)
);

XOR2xp5_ASAP7_75t_L g514 ( 
.A(n_503),
.B(n_4),
.Y(n_514)
);

NOR2xp33_ASAP7_75t_L g504 ( 
.A(n_495),
.B(n_476),
.Y(n_504)
);

OR2x2_ASAP7_75t_L g522 ( 
.A(n_504),
.B(n_506),
.Y(n_522)
);

AOI31xp67_ASAP7_75t_SL g505 ( 
.A1(n_492),
.A2(n_469),
.A3(n_486),
.B(n_468),
.Y(n_505)
);

INVx1_ASAP7_75t_L g523 ( 
.A(n_505),
.Y(n_523)
);

MAJIxp5_ASAP7_75t_L g506 ( 
.A(n_498),
.B(n_482),
.C(n_485),
.Y(n_506)
);

NAND2xp5_ASAP7_75t_L g519 ( 
.A(n_508),
.B(n_510),
.Y(n_519)
);

XOR2xp5_ASAP7_75t_L g509 ( 
.A(n_487),
.B(n_475),
.Y(n_509)
);

HB1xp67_ASAP7_75t_L g525 ( 
.A(n_509),
.Y(n_525)
);

XOR2xp5_ASAP7_75t_L g510 ( 
.A(n_486),
.B(n_2),
.Y(n_510)
);

FAx1_ASAP7_75t_L g511 ( 
.A(n_489),
.B(n_3),
.CI(n_4),
.CON(n_511),
.SN(n_511)
);

AOI21xp5_ASAP7_75t_SL g524 ( 
.A1(n_511),
.A2(n_493),
.B(n_503),
.Y(n_524)
);

NOR2xp33_ASAP7_75t_L g512 ( 
.A(n_488),
.B(n_3),
.Y(n_512)
);

NAND2xp5_ASAP7_75t_L g520 ( 
.A(n_512),
.B(n_514),
.Y(n_520)
);

NAND2xp5_ASAP7_75t_L g528 ( 
.A(n_515),
.B(n_516),
.Y(n_528)
);

INVx1_ASAP7_75t_SL g516 ( 
.A(n_493),
.Y(n_516)
);

MAJIxp5_ASAP7_75t_L g521 ( 
.A(n_517),
.B(n_507),
.C(n_513),
.Y(n_521)
);

NAND2xp5_ASAP7_75t_L g533 ( 
.A(n_521),
.B(n_526),
.Y(n_533)
);

NOR2xp33_ASAP7_75t_L g531 ( 
.A(n_524),
.B(n_5),
.Y(n_531)
);

NOR2xp33_ASAP7_75t_L g526 ( 
.A(n_516),
.B(n_509),
.Y(n_526)
);

OAI21xp33_ASAP7_75t_L g527 ( 
.A1(n_518),
.A2(n_499),
.B(n_500),
.Y(n_527)
);

NAND2xp5_ASAP7_75t_L g537 ( 
.A(n_527),
.B(n_8),
.Y(n_537)
);

OAI22xp5_ASAP7_75t_L g529 ( 
.A1(n_511),
.A2(n_5),
.B1(n_6),
.B2(n_7),
.Y(n_529)
);

AOI22xp5_ASAP7_75t_SL g534 ( 
.A1(n_529),
.A2(n_12),
.B1(n_7),
.B2(n_8),
.Y(n_534)
);

AOI21x1_ASAP7_75t_L g530 ( 
.A1(n_523),
.A2(n_511),
.B(n_510),
.Y(n_530)
);

AOI21xp5_ASAP7_75t_L g539 ( 
.A1(n_530),
.A2(n_529),
.B(n_9),
.Y(n_539)
);

NOR2xp67_ASAP7_75t_SL g542 ( 
.A(n_531),
.B(n_535),
.Y(n_542)
);

INVx6_ASAP7_75t_L g532 ( 
.A(n_522),
.Y(n_532)
);

HB1xp67_ASAP7_75t_L g538 ( 
.A(n_532),
.Y(n_538)
);

OAI21xp5_ASAP7_75t_L g541 ( 
.A1(n_534),
.A2(n_536),
.B(n_10),
.Y(n_541)
);

MAJIxp5_ASAP7_75t_L g535 ( 
.A(n_525),
.B(n_6),
.C(n_8),
.Y(n_535)
);

MAJIxp5_ASAP7_75t_L g536 ( 
.A(n_519),
.B(n_528),
.C(n_520),
.Y(n_536)
);

A2O1A1Ixp33_ASAP7_75t_SL g540 ( 
.A1(n_537),
.A2(n_8),
.B(n_10),
.C(n_11),
.Y(n_540)
);

AO21x1_ASAP7_75t_L g544 ( 
.A1(n_539),
.A2(n_531),
.B(n_533),
.Y(n_544)
);

OR2x2_ASAP7_75t_L g543 ( 
.A(n_540),
.B(n_541),
.Y(n_543)
);

NOR2xp33_ASAP7_75t_L g546 ( 
.A(n_544),
.B(n_545),
.Y(n_546)
);

MAJIxp5_ASAP7_75t_L g545 ( 
.A(n_538),
.B(n_532),
.C(n_11),
.Y(n_545)
);

OAI21xp5_ASAP7_75t_L g547 ( 
.A1(n_546),
.A2(n_542),
.B(n_543),
.Y(n_547)
);

OAI21xp5_ASAP7_75t_L g548 ( 
.A1(n_547),
.A2(n_10),
.B(n_11),
.Y(n_548)
);

NAND2xp5_ASAP7_75t_L g549 ( 
.A(n_548),
.B(n_11),
.Y(n_549)
);

MAJIxp5_ASAP7_75t_L g550 ( 
.A(n_549),
.B(n_12),
.C(n_529),
.Y(n_550)
);


endmodule