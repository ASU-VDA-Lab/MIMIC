module real_jpeg_15573_n_17 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_16, n_3, n_10, n_9, n_17);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_16;
input n_3;
input n_10;
input n_9;

output n_17;

wire n_384;
wire n_37;
wire n_430;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_300;
wire n_415;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_446;
wire n_199;
wire n_95;
wire n_441;
wire n_238;
wire n_67;
wire n_350;
wire n_235;
wire n_107;
wire n_369;
wire n_376;
wire n_354;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_355;
wire n_123;
wire n_425;
wire n_50;
wire n_409;
wire n_186;
wire n_137;
wire n_72;
wire n_440;
wire n_171;
wire n_151;
wire n_272;
wire n_203;
wire n_198;
wire n_23;
wire n_362;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_326;
wire n_339;
wire n_80;
wire n_30;
wire n_328;
wire n_149;
wire n_332;
wire n_366;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_353;
wire n_453;
wire n_230;
wire n_417;
wire n_428;
wire n_216;
wire n_128;
wire n_202;
wire n_367;
wire n_127;
wire n_356;
wire n_365;
wire n_423;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_422;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_348;
wire n_252;
wire n_363;
wire n_310;
wire n_345;
wire n_83;
wire n_78;
wire n_288;
wire n_221;
wire n_393;
wire n_104;
wire n_153;
wire n_443;
wire n_337;
wire n_131;
wire n_439;
wire n_322;
wire n_87;
wire n_40;
wire n_378;
wire n_98;
wire n_200;
wire n_432;
wire n_335;
wire n_214;
wire n_113;
wire n_251;
wire n_139;
wire n_33;
wire n_175;
wire n_338;
wire n_156;
wire n_387;
wire n_434;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_390;
wire n_77;
wire n_399;
wire n_219;
wire n_372;
wire n_122;
wire n_19;
wire n_262;
wire n_334;
wire n_383;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_426;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_371;
wire n_410;
wire n_421;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_411;
wire n_382;
wire n_20;
wire n_278;
wire n_314;
wire n_103;
wire n_232;
wire n_448;
wire n_212;
wire n_284;
wire n_402;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_452;
wire n_213;
wire n_25;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_407;
wire n_419;
wire n_386;
wire n_341;
wire n_331;
wire n_49;
wire n_68;
wire n_395;
wire n_146;
wire n_286;
wire n_166;
wire n_176;
wire n_215;
wire n_323;
wire n_312;
wire n_325;
wire n_307;
wire n_316;
wire n_161;
wire n_207;
wire n_431;
wire n_420;
wire n_357;
wire n_237;
wire n_445;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_380;
wire n_414;
wire n_140;
wire n_126;
wire n_342;
wire n_120;
wire n_155;
wire n_412;
wire n_405;
wire n_319;
wire n_93;
wire n_242;
wire n_142;
wire n_397;
wire n_76;
wire n_403;
wire n_79;
wire n_282;
wire n_147;
wire n_359;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_449;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_145;
wire n_18;
wire n_266;
wire n_377;
wire n_109;
wire n_391;
wire n_427;
wire n_401;
wire n_148;
wire n_373;
wire n_396;
wire n_392;
wire n_375;
wire n_196;
wire n_330;
wire n_298;
wire n_333;
wire n_450;
wire n_152;
wire n_270;
wire n_159;
wire n_429;
wire n_347;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_336;
wire n_258;
wire n_150;
wire n_41;
wire n_74;
wire n_404;
wire n_158;
wire n_204;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_413;
wire n_75;
wire n_346;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_119;
wire n_283;
wire n_181;
wire n_358;
wire n_256;
wire n_253;
wire n_273;
wire n_54;
wire n_168;
wire n_38;
wire n_442;
wire n_385;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_349;
wire n_418;
wire n_292;
wire n_343;
wire n_64;
wire n_291;
wire n_236;
wire n_370;
wire n_276;
wire n_374;
wire n_287;
wire n_400;
wire n_174;
wire n_388;
wire n_255;
wire n_243;
wire n_299;
wire n_352;
wire n_56;
wire n_293;
wire n_275;
wire n_381;
wire n_227;
wire n_229;
wire n_379;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_444;
wire n_360;
wire n_398;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_451;
wire n_45;
wire n_437;
wire n_313;
wire n_42;
wire n_268;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_416;
wire n_143;
wire n_351;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_406;
wire n_303;
wire n_321;
wire n_100;
wire n_368;
wire n_51;
wire n_205;
wire n_361;
wire n_324;
wire n_86;
wire n_261;
wire n_70;
wire n_435;
wire n_32;
wire n_228;
wire n_389;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_438;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_394;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_436;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_424;
wire n_133;
wire n_257;
wire n_447;
wire n_344;
wire n_210;
wire n_206;
wire n_408;
wire n_85;
wire n_96;
wire n_308;
wire n_433;
wire n_364;

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_0),
.Y(n_57)
);

BUFx3_ASAP7_75t_L g73 ( 
.A(n_0),
.Y(n_73)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_0),
.Y(n_131)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_0),
.Y(n_187)
);

AND2x2_ASAP7_75t_L g28 ( 
.A(n_1),
.B(n_29),
.Y(n_28)
);

NAND2xp5_ASAP7_75t_SL g55 ( 
.A(n_1),
.B(n_56),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_L g104 ( 
.A(n_1),
.B(n_105),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_SL g124 ( 
.A(n_1),
.B(n_125),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_SL g176 ( 
.A(n_1),
.B(n_177),
.Y(n_176)
);

AND2x2_ASAP7_75t_L g232 ( 
.A(n_1),
.B(n_233),
.Y(n_232)
);

INVxp33_ASAP7_75t_L g269 ( 
.A(n_1),
.Y(n_269)
);

AND2x2_ASAP7_75t_L g323 ( 
.A(n_1),
.B(n_208),
.Y(n_323)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_2),
.Y(n_68)
);

BUFx6f_ASAP7_75t_L g233 ( 
.A(n_2),
.Y(n_233)
);

BUFx6f_ASAP7_75t_L g236 ( 
.A(n_2),
.Y(n_236)
);

BUFx5_ASAP7_75t_L g278 ( 
.A(n_2),
.Y(n_278)
);

INVx1_ASAP7_75t_L g366 ( 
.A(n_2),
.Y(n_366)
);

NAND2xp5_ASAP7_75t_SL g64 ( 
.A(n_3),
.B(n_65),
.Y(n_64)
);

AND2x2_ASAP7_75t_L g81 ( 
.A(n_3),
.B(n_82),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g111 ( 
.A(n_3),
.B(n_112),
.Y(n_111)
);

AND2x2_ASAP7_75t_L g136 ( 
.A(n_3),
.B(n_137),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_L g184 ( 
.A(n_3),
.B(n_185),
.Y(n_184)
);

BUFx5_ASAP7_75t_L g38 ( 
.A(n_4),
.Y(n_38)
);

INVx2_ASAP7_75t_L g140 ( 
.A(n_4),
.Y(n_140)
);

BUFx3_ASAP7_75t_L g210 ( 
.A(n_4),
.Y(n_210)
);

BUFx5_ASAP7_75t_L g317 ( 
.A(n_4),
.Y(n_317)
);

NAND2xp5_ASAP7_75t_SL g228 ( 
.A(n_5),
.B(n_229),
.Y(n_228)
);

NAND2xp5_ASAP7_75t_L g325 ( 
.A(n_5),
.B(n_326),
.Y(n_325)
);

NAND2xp5_ASAP7_75t_SL g344 ( 
.A(n_5),
.B(n_312),
.Y(n_344)
);

NAND2xp5_ASAP7_75t_L g360 ( 
.A(n_5),
.B(n_361),
.Y(n_360)
);

NAND2xp5_ASAP7_75t_L g410 ( 
.A(n_5),
.B(n_411),
.Y(n_410)
);

NAND2xp5_ASAP7_75t_SL g414 ( 
.A(n_5),
.B(n_415),
.Y(n_414)
);

NAND2xp5_ASAP7_75t_SL g420 ( 
.A(n_5),
.B(n_421),
.Y(n_420)
);

INVx1_ASAP7_75t_SL g34 ( 
.A(n_6),
.Y(n_34)
);

AND2x2_ASAP7_75t_L g37 ( 
.A(n_6),
.B(n_38),
.Y(n_37)
);

AND2x2_ASAP7_75t_L g161 ( 
.A(n_6),
.B(n_162),
.Y(n_161)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_7),
.Y(n_54)
);

INVx3_ASAP7_75t_L g78 ( 
.A(n_7),
.Y(n_78)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_7),
.Y(n_115)
);

BUFx5_ASAP7_75t_L g162 ( 
.A(n_7),
.Y(n_162)
);

BUFx6f_ASAP7_75t_L g281 ( 
.A(n_7),
.Y(n_281)
);

BUFx3_ASAP7_75t_L g346 ( 
.A(n_7),
.Y(n_346)
);

NAND2xp5_ASAP7_75t_SL g80 ( 
.A(n_8),
.B(n_59),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_SL g122 ( 
.A(n_8),
.B(n_123),
.Y(n_122)
);

AOI22xp5_ASAP7_75t_SL g205 ( 
.A1(n_8),
.A2(n_11),
.B1(n_206),
.B2(n_211),
.Y(n_205)
);

AND2x2_ASAP7_75t_L g274 ( 
.A(n_8),
.B(n_275),
.Y(n_274)
);

AND2x2_ASAP7_75t_L g310 ( 
.A(n_8),
.B(n_311),
.Y(n_310)
);

NAND2xp5_ASAP7_75t_SL g345 ( 
.A(n_8),
.B(n_346),
.Y(n_345)
);

NAND2xp5_ASAP7_75t_L g363 ( 
.A(n_8),
.B(n_364),
.Y(n_363)
);

AND2x2_ASAP7_75t_L g369 ( 
.A(n_8),
.B(n_370),
.Y(n_369)
);

NAND2xp5_ASAP7_75t_L g401 ( 
.A(n_8),
.B(n_402),
.Y(n_401)
);

NAND2xp5_ASAP7_75t_L g47 ( 
.A(n_9),
.B(n_48),
.Y(n_47)
);

NAND2xp5_ASAP7_75t_SL g58 ( 
.A(n_9),
.B(n_59),
.Y(n_58)
);

AND2x2_ASAP7_75t_L g216 ( 
.A(n_9),
.B(n_217),
.Y(n_216)
);

NAND2xp5_ASAP7_75t_L g237 ( 
.A(n_9),
.B(n_238),
.Y(n_237)
);

AND2x2_ASAP7_75t_L g279 ( 
.A(n_9),
.B(n_280),
.Y(n_279)
);

AND2x2_ASAP7_75t_L g374 ( 
.A(n_9),
.B(n_375),
.Y(n_374)
);

NAND2xp5_ASAP7_75t_L g377 ( 
.A(n_9),
.B(n_378),
.Y(n_377)
);

NAND2xp5_ASAP7_75t_SL g394 ( 
.A(n_9),
.B(n_395),
.Y(n_394)
);

NAND2xp5_ASAP7_75t_L g51 ( 
.A(n_10),
.B(n_52),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_L g70 ( 
.A(n_10),
.B(n_71),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_SL g91 ( 
.A(n_10),
.B(n_92),
.Y(n_91)
);

INVxp33_ASAP7_75t_L g165 ( 
.A(n_10),
.Y(n_165)
);

AND2x2_ASAP7_75t_L g219 ( 
.A(n_10),
.B(n_220),
.Y(n_219)
);

AND2x4_ASAP7_75t_SL g235 ( 
.A(n_10),
.B(n_236),
.Y(n_235)
);

AND2x2_ASAP7_75t_SL g272 ( 
.A(n_10),
.B(n_137),
.Y(n_272)
);

NAND2xp5_ASAP7_75t_SL g74 ( 
.A(n_11),
.B(n_75),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_L g108 ( 
.A(n_11),
.B(n_109),
.Y(n_108)
);

AND2x2_ASAP7_75t_L g141 ( 
.A(n_11),
.B(n_142),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_SL g144 ( 
.A(n_11),
.B(n_145),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_L g180 ( 
.A(n_11),
.B(n_181),
.Y(n_180)
);

CKINVDCx16_ASAP7_75t_R g314 ( 
.A(n_11),
.Y(n_314)
);

INVx6_ASAP7_75t_L g42 ( 
.A(n_12),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_12),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g168 ( 
.A(n_12),
.Y(n_168)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_13),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g95 ( 
.A(n_13),
.Y(n_95)
);

BUFx4f_ASAP7_75t_L g36 ( 
.A(n_14),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g223 ( 
.A(n_14),
.Y(n_223)
);

BUFx12f_ASAP7_75t_L g271 ( 
.A(n_14),
.Y(n_271)
);

INVx2_ASAP7_75t_L g373 ( 
.A(n_14),
.Y(n_373)
);

NAND2x1_ASAP7_75t_L g26 ( 
.A(n_15),
.B(n_27),
.Y(n_26)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_15),
.Y(n_40)
);

AND2x2_ASAP7_75t_SL g128 ( 
.A(n_15),
.B(n_129),
.Y(n_128)
);

AND2x2_ASAP7_75t_SL g147 ( 
.A(n_15),
.B(n_148),
.Y(n_147)
);

AND2x2_ASAP7_75t_L g226 ( 
.A(n_15),
.B(n_227),
.Y(n_226)
);

AND2x2_ASAP7_75t_L g277 ( 
.A(n_15),
.B(n_278),
.Y(n_277)
);

AND2x2_ASAP7_75t_L g320 ( 
.A(n_15),
.B(n_321),
.Y(n_320)
);

AND2x2_ASAP7_75t_L g380 ( 
.A(n_15),
.B(n_381),
.Y(n_380)
);

BUFx8_ASAP7_75t_L g27 ( 
.A(n_16),
.Y(n_27)
);

BUFx3_ASAP7_75t_L g60 ( 
.A(n_16),
.Y(n_60)
);

INVx2_ASAP7_75t_L g231 ( 
.A(n_16),
.Y(n_231)
);

XOR2xp5_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_194),
.Y(n_17)
);

NAND2xp5_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_192),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_20),
.Y(n_19)
);

NOR2xp67_ASAP7_75t_SL g20 ( 
.A(n_21),
.B(n_154),
.Y(n_20)
);

AND2x2_ASAP7_75t_L g193 ( 
.A(n_21),
.B(n_154),
.Y(n_193)
);

MAJIxp5_ASAP7_75t_L g21 ( 
.A(n_22),
.B(n_89),
.C(n_116),
.Y(n_21)
);

XNOR2xp5_ASAP7_75t_L g290 ( 
.A(n_22),
.B(n_89),
.Y(n_290)
);

XNOR2xp5_ASAP7_75t_L g22 ( 
.A(n_23),
.B(n_62),
.Y(n_22)
);

XNOR2xp5_ASAP7_75t_L g23 ( 
.A(n_24),
.B(n_45),
.Y(n_23)
);

MAJIxp5_ASAP7_75t_L g155 ( 
.A(n_24),
.B(n_45),
.C(n_156),
.Y(n_155)
);

AOI22xp5_ASAP7_75t_L g24 ( 
.A1(n_25),
.A2(n_32),
.B1(n_43),
.B2(n_44),
.Y(n_24)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_25),
.Y(n_43)
);

XOR2xp5_ASAP7_75t_L g25 ( 
.A(n_26),
.B(n_28),
.Y(n_25)
);

MAJIxp5_ASAP7_75t_L g135 ( 
.A(n_26),
.B(n_136),
.C(n_141),
.Y(n_135)
);

MAJx2_ASAP7_75t_L g174 ( 
.A(n_26),
.B(n_28),
.C(n_44),
.Y(n_174)
);

XNOR2xp5_ASAP7_75t_L g202 ( 
.A(n_26),
.B(n_203),
.Y(n_202)
);

INVx2_ASAP7_75t_L g178 ( 
.A(n_27),
.Y(n_178)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_28),
.Y(n_61)
);

OAI22xp5_ASAP7_75t_SL g152 ( 
.A1(n_28),
.A2(n_58),
.B1(n_61),
.B2(n_153),
.Y(n_152)
);

INVx6_ASAP7_75t_L g29 ( 
.A(n_30),
.Y(n_29)
);

INVx4_ASAP7_75t_L g30 ( 
.A(n_31),
.Y(n_30)
);

INVx3_ASAP7_75t_L g240 ( 
.A(n_31),
.Y(n_240)
);

INVx1_ASAP7_75t_SL g44 ( 
.A(n_32),
.Y(n_44)
);

MAJx2_ASAP7_75t_L g32 ( 
.A(n_33),
.B(n_37),
.C(n_39),
.Y(n_32)
);

OAI22xp5_ASAP7_75t_SL g86 ( 
.A1(n_33),
.A2(n_37),
.B1(n_87),
.B2(n_88),
.Y(n_86)
);

INVx1_ASAP7_75t_SL g88 ( 
.A(n_33),
.Y(n_88)
);

AOI22xp33_ASAP7_75t_L g96 ( 
.A1(n_33),
.A2(n_88),
.B1(n_97),
.B2(n_98),
.Y(n_96)
);

OR2x2_ASAP7_75t_L g33 ( 
.A(n_34),
.B(n_35),
.Y(n_33)
);

OR2x2_ASAP7_75t_L g98 ( 
.A(n_34),
.B(n_99),
.Y(n_98)
);

INVx2_ASAP7_75t_L g82 ( 
.A(n_35),
.Y(n_82)
);

INVx1_ASAP7_75t_L g421 ( 
.A(n_35),
.Y(n_421)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_36),
.Y(n_35)
);

INVx2_ASAP7_75t_L g143 ( 
.A(n_36),
.Y(n_143)
);

MAJIxp5_ASAP7_75t_L g79 ( 
.A(n_37),
.B(n_80),
.C(n_81),
.Y(n_79)
);

INVx1_ASAP7_75t_SL g87 ( 
.A(n_37),
.Y(n_87)
);

AOI22xp5_ASAP7_75t_SL g119 ( 
.A1(n_37),
.A2(n_81),
.B1(n_87),
.B2(n_120),
.Y(n_119)
);

BUFx3_ASAP7_75t_L g375 ( 
.A(n_38),
.Y(n_375)
);

INVx3_ASAP7_75t_L g403 ( 
.A(n_38),
.Y(n_403)
);

AOI22xp5_ASAP7_75t_L g83 ( 
.A1(n_39),
.A2(n_84),
.B1(n_85),
.B2(n_86),
.Y(n_83)
);

INVx1_ASAP7_75t_SL g84 ( 
.A(n_39),
.Y(n_84)
);

AOI22xp5_ASAP7_75t_L g265 ( 
.A1(n_39),
.A2(n_84),
.B1(n_219),
.B2(n_266),
.Y(n_265)
);

OR2x2_ASAP7_75t_L g39 ( 
.A(n_40),
.B(n_41),
.Y(n_39)
);

INVx2_ASAP7_75t_L g326 ( 
.A(n_41),
.Y(n_326)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_42),
.Y(n_41)
);

INVx4_ASAP7_75t_L g123 ( 
.A(n_42),
.Y(n_123)
);

MAJIxp5_ASAP7_75t_L g45 ( 
.A(n_46),
.B(n_58),
.C(n_61),
.Y(n_45)
);

XNOR2xp5_ASAP7_75t_L g151 ( 
.A(n_46),
.B(n_152),
.Y(n_151)
);

MAJIxp5_ASAP7_75t_L g46 ( 
.A(n_47),
.B(n_51),
.C(n_55),
.Y(n_46)
);

XNOR2xp5_ASAP7_75t_L g133 ( 
.A(n_47),
.B(n_55),
.Y(n_133)
);

INVx4_ASAP7_75t_L g48 ( 
.A(n_49),
.Y(n_48)
);

INVx6_ASAP7_75t_L g49 ( 
.A(n_50),
.Y(n_49)
);

INVx4_ASAP7_75t_L g106 ( 
.A(n_50),
.Y(n_106)
);

XOR2xp5_ASAP7_75t_L g132 ( 
.A(n_51),
.B(n_133),
.Y(n_132)
);

INVx5_ASAP7_75t_L g52 ( 
.A(n_53),
.Y(n_52)
);

INVx2_ASAP7_75t_L g53 ( 
.A(n_54),
.Y(n_53)
);

INVx6_ASAP7_75t_L g110 ( 
.A(n_56),
.Y(n_110)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_57),
.Y(n_56)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_58),
.Y(n_153)
);

BUFx12f_ASAP7_75t_L g59 ( 
.A(n_60),
.Y(n_59)
);

INVxp67_ASAP7_75t_L g156 ( 
.A(n_62),
.Y(n_156)
);

MAJIxp5_ASAP7_75t_L g62 ( 
.A(n_63),
.B(n_79),
.C(n_83),
.Y(n_62)
);

XNOR2xp5_ASAP7_75t_L g250 ( 
.A(n_63),
.B(n_79),
.Y(n_250)
);

XNOR2xp5_ASAP7_75t_L g63 ( 
.A(n_64),
.B(n_69),
.Y(n_63)
);

MAJIxp5_ASAP7_75t_L g102 ( 
.A(n_64),
.B(n_70),
.C(n_74),
.Y(n_102)
);

HB1xp67_ASAP7_75t_L g65 ( 
.A(n_66),
.Y(n_65)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_67),
.Y(n_66)
);

INVx4_ASAP7_75t_L g145 ( 
.A(n_67),
.Y(n_145)
);

BUFx3_ASAP7_75t_L g67 ( 
.A(n_68),
.Y(n_67)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_68),
.Y(n_100)
);

XNOR2xp5_ASAP7_75t_L g69 ( 
.A(n_70),
.B(n_74),
.Y(n_69)
);

INVx2_ASAP7_75t_L g71 ( 
.A(n_72),
.Y(n_71)
);

INVx2_ASAP7_75t_L g72 ( 
.A(n_73),
.Y(n_72)
);

INVx1_ASAP7_75t_L g362 ( 
.A(n_73),
.Y(n_362)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_76),
.Y(n_75)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_77),
.Y(n_76)
);

INVx2_ASAP7_75t_L g77 ( 
.A(n_78),
.Y(n_77)
);

BUFx3_ASAP7_75t_L g126 ( 
.A(n_78),
.Y(n_126)
);

XNOR2x1_ASAP7_75t_L g118 ( 
.A(n_80),
.B(n_119),
.Y(n_118)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_81),
.Y(n_120)
);

XOR2xp5_ASAP7_75t_L g249 ( 
.A(n_83),
.B(n_250),
.Y(n_249)
);

MAJx2_ASAP7_75t_L g215 ( 
.A(n_84),
.B(n_216),
.C(n_219),
.Y(n_215)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_86),
.Y(n_85)
);

MAJIxp5_ASAP7_75t_L g170 ( 
.A(n_88),
.B(n_91),
.C(n_98),
.Y(n_170)
);

XNOR2xp5_ASAP7_75t_L g89 ( 
.A(n_90),
.B(n_101),
.Y(n_89)
);

MAJIxp5_ASAP7_75t_L g189 ( 
.A(n_90),
.B(n_102),
.C(n_103),
.Y(n_189)
);

XOR2xp5_ASAP7_75t_L g90 ( 
.A(n_91),
.B(n_96),
.Y(n_90)
);

INVx2_ASAP7_75t_L g92 ( 
.A(n_93),
.Y(n_92)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_94),
.Y(n_93)
);

INVx4_ASAP7_75t_L g182 ( 
.A(n_94),
.Y(n_182)
);

INVx2_ASAP7_75t_L g214 ( 
.A(n_94),
.Y(n_214)
);

BUFx6f_ASAP7_75t_L g94 ( 
.A(n_95),
.Y(n_94)
);

INVx2_ASAP7_75t_L g150 ( 
.A(n_95),
.Y(n_150)
);

AOI22xp5_ASAP7_75t_L g160 ( 
.A1(n_97),
.A2(n_98),
.B1(n_161),
.B2(n_163),
.Y(n_160)
);

INVx1_ASAP7_75t_SL g97 ( 
.A(n_98),
.Y(n_97)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_100),
.Y(n_99)
);

XNOR2xp5_ASAP7_75t_L g101 ( 
.A(n_102),
.B(n_103),
.Y(n_101)
);

XOR2xp5_ASAP7_75t_L g103 ( 
.A(n_104),
.B(n_107),
.Y(n_103)
);

MAJIxp5_ASAP7_75t_L g171 ( 
.A(n_104),
.B(n_108),
.C(n_111),
.Y(n_171)
);

INVx2_ASAP7_75t_L g105 ( 
.A(n_106),
.Y(n_105)
);

XNOR2xp5_ASAP7_75t_L g107 ( 
.A(n_108),
.B(n_111),
.Y(n_107)
);

INVx8_ASAP7_75t_L g109 ( 
.A(n_110),
.Y(n_109)
);

INVx2_ASAP7_75t_L g112 ( 
.A(n_113),
.Y(n_112)
);

INVx2_ASAP7_75t_L g113 ( 
.A(n_114),
.Y(n_113)
);

INVx2_ASAP7_75t_L g114 ( 
.A(n_115),
.Y(n_114)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_115),
.Y(n_227)
);

XOR2xp5_ASAP7_75t_L g289 ( 
.A(n_116),
.B(n_290),
.Y(n_289)
);

MAJIxp5_ASAP7_75t_L g116 ( 
.A(n_117),
.B(n_134),
.C(n_151),
.Y(n_116)
);

XNOR2xp5_ASAP7_75t_SL g247 ( 
.A(n_117),
.B(n_248),
.Y(n_247)
);

MAJIxp5_ASAP7_75t_L g117 ( 
.A(n_118),
.B(n_121),
.C(n_132),
.Y(n_117)
);

XNOR2xp5_ASAP7_75t_L g259 ( 
.A(n_118),
.B(n_121),
.Y(n_259)
);

MAJIxp5_ASAP7_75t_L g121 ( 
.A(n_122),
.B(n_124),
.C(n_127),
.Y(n_121)
);

AOI22xp5_ASAP7_75t_L g286 ( 
.A1(n_122),
.A2(n_127),
.B1(n_128),
.B2(n_287),
.Y(n_286)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_122),
.Y(n_287)
);

XOR2xp5_ASAP7_75t_L g285 ( 
.A(n_124),
.B(n_286),
.Y(n_285)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_126),
.Y(n_125)
);

INVxp67_ASAP7_75t_SL g411 ( 
.A(n_126),
.Y(n_411)
);

MAJIxp5_ASAP7_75t_L g343 ( 
.A(n_127),
.B(n_344),
.C(n_345),
.Y(n_343)
);

AOI22xp5_ASAP7_75t_L g388 ( 
.A1(n_127),
.A2(n_128),
.B1(n_344),
.B2(n_389),
.Y(n_388)
);

INVx2_ASAP7_75t_L g127 ( 
.A(n_128),
.Y(n_127)
);

INVx4_ASAP7_75t_L g129 ( 
.A(n_130),
.Y(n_129)
);

INVx2_ASAP7_75t_L g218 ( 
.A(n_130),
.Y(n_218)
);

BUFx3_ASAP7_75t_L g130 ( 
.A(n_131),
.Y(n_130)
);

BUFx3_ASAP7_75t_L g276 ( 
.A(n_131),
.Y(n_276)
);

XNOR2x1_ASAP7_75t_SL g258 ( 
.A(n_132),
.B(n_259),
.Y(n_258)
);

XNOR2xp5_ASAP7_75t_L g248 ( 
.A(n_134),
.B(n_151),
.Y(n_248)
);

MAJx2_ASAP7_75t_L g134 ( 
.A(n_135),
.B(n_144),
.C(n_146),
.Y(n_134)
);

XNOR2xp5_ASAP7_75t_L g243 ( 
.A(n_135),
.B(n_244),
.Y(n_243)
);

XNOR2xp5_ASAP7_75t_L g203 ( 
.A(n_136),
.B(n_141),
.Y(n_203)
);

INVx2_ASAP7_75t_L g137 ( 
.A(n_138),
.Y(n_137)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_139),
.Y(n_138)
);

INVx2_ASAP7_75t_L g139 ( 
.A(n_140),
.Y(n_139)
);

INVx3_ASAP7_75t_L g381 ( 
.A(n_140),
.Y(n_381)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_143),
.Y(n_142)
);

AOI22xp5_ASAP7_75t_L g244 ( 
.A1(n_144),
.A2(n_146),
.B1(n_147),
.B2(n_245),
.Y(n_244)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_144),
.Y(n_245)
);

AOI22xp5_ASAP7_75t_L g437 ( 
.A1(n_146),
.A2(n_147),
.B1(n_324),
.B2(n_325),
.Y(n_437)
);

INVx2_ASAP7_75t_SL g146 ( 
.A(n_147),
.Y(n_146)
);

MAJIxp5_ASAP7_75t_L g318 ( 
.A(n_147),
.B(n_319),
.C(n_324),
.Y(n_318)
);

INVx4_ASAP7_75t_L g148 ( 
.A(n_149),
.Y(n_148)
);

BUFx6f_ASAP7_75t_L g149 ( 
.A(n_150),
.Y(n_149)
);

XOR2xp5_ASAP7_75t_L g154 ( 
.A(n_155),
.B(n_157),
.Y(n_154)
);

AOI22xp5_ASAP7_75t_L g157 ( 
.A1(n_158),
.A2(n_172),
.B1(n_190),
.B2(n_191),
.Y(n_157)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_158),
.Y(n_190)
);

XNOR2xp5_ASAP7_75t_L g158 ( 
.A(n_159),
.B(n_169),
.Y(n_158)
);

XNOR2xp5_ASAP7_75t_SL g159 ( 
.A(n_160),
.B(n_164),
.Y(n_159)
);

INVx1_ASAP7_75t_SL g163 ( 
.A(n_161),
.Y(n_163)
);

NOR2xp33_ASAP7_75t_L g164 ( 
.A(n_165),
.B(n_166),
.Y(n_164)
);

HB1xp67_ASAP7_75t_L g166 ( 
.A(n_167),
.Y(n_166)
);

INVx3_ASAP7_75t_L g167 ( 
.A(n_168),
.Y(n_167)
);

XNOR2xp5_ASAP7_75t_L g169 ( 
.A(n_170),
.B(n_171),
.Y(n_169)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_172),
.Y(n_191)
);

XNOR2xp5_ASAP7_75t_L g172 ( 
.A(n_173),
.B(n_189),
.Y(n_172)
);

XNOR2xp5_ASAP7_75t_L g173 ( 
.A(n_174),
.B(n_175),
.Y(n_173)
);

XNOR2xp5_ASAP7_75t_L g175 ( 
.A(n_176),
.B(n_179),
.Y(n_175)
);

INVx2_ASAP7_75t_L g177 ( 
.A(n_178),
.Y(n_177)
);

AOI22xp5_ASAP7_75t_L g179 ( 
.A1(n_180),
.A2(n_183),
.B1(n_184),
.B2(n_188),
.Y(n_179)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_180),
.Y(n_188)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_182),
.Y(n_181)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_184),
.Y(n_183)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_186),
.Y(n_185)
);

BUFx6f_ASAP7_75t_L g186 ( 
.A(n_187),
.Y(n_186)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_193),
.Y(n_192)
);

HB1xp67_ASAP7_75t_L g194 ( 
.A(n_195),
.Y(n_194)
);

AO21x2_ASAP7_75t_L g195 ( 
.A1(n_196),
.A2(n_294),
.B(n_451),
.Y(n_195)
);

NOR2xp33_ASAP7_75t_L g196 ( 
.A(n_197),
.B(n_288),
.Y(n_196)
);

AND2x2_ASAP7_75t_SL g197 ( 
.A(n_198),
.B(n_253),
.Y(n_197)
);

OR2x2_ASAP7_75t_L g452 ( 
.A(n_198),
.B(n_253),
.Y(n_452)
);

XNOR2xp5_ASAP7_75t_L g198 ( 
.A(n_199),
.B(n_246),
.Y(n_198)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_199),
.Y(n_292)
);

MAJIxp5_ASAP7_75t_L g199 ( 
.A(n_200),
.B(n_224),
.C(n_241),
.Y(n_199)
);

INVxp33_ASAP7_75t_SL g200 ( 
.A(n_201),
.Y(n_200)
);

XNOR2xp5_ASAP7_75t_L g255 ( 
.A(n_201),
.B(n_256),
.Y(n_255)
);

MAJIxp5_ASAP7_75t_L g201 ( 
.A(n_202),
.B(n_204),
.C(n_215),
.Y(n_201)
);

XNOR2xp5_ASAP7_75t_L g328 ( 
.A(n_202),
.B(n_329),
.Y(n_328)
);

AOI22xp5_ASAP7_75t_SL g329 ( 
.A1(n_204),
.A2(n_205),
.B1(n_215),
.B2(n_330),
.Y(n_329)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_205),
.Y(n_204)
);

AOI21xp5_ASAP7_75t_L g309 ( 
.A1(n_205),
.A2(n_310),
.B(n_313),
.Y(n_309)
);

INVx3_ASAP7_75t_L g206 ( 
.A(n_207),
.Y(n_206)
);

INVx5_ASAP7_75t_L g207 ( 
.A(n_208),
.Y(n_207)
);

INVx4_ASAP7_75t_L g208 ( 
.A(n_209),
.Y(n_208)
);

INVx3_ASAP7_75t_L g209 ( 
.A(n_210),
.Y(n_209)
);

INVx2_ASAP7_75t_L g211 ( 
.A(n_212),
.Y(n_211)
);

INVx2_ASAP7_75t_L g212 ( 
.A(n_213),
.Y(n_212)
);

INVx2_ASAP7_75t_L g213 ( 
.A(n_214),
.Y(n_213)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_215),
.Y(n_330)
);

XNOR2xp5_ASAP7_75t_L g264 ( 
.A(n_216),
.B(n_265),
.Y(n_264)
);

HB1xp67_ASAP7_75t_L g217 ( 
.A(n_218),
.Y(n_217)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_219),
.Y(n_266)
);

BUFx2_ASAP7_75t_SL g220 ( 
.A(n_221),
.Y(n_220)
);

INVx2_ASAP7_75t_L g221 ( 
.A(n_222),
.Y(n_221)
);

INVx2_ASAP7_75t_L g222 ( 
.A(n_223),
.Y(n_222)
);

AOI22xp5_ASAP7_75t_SL g256 ( 
.A1(n_224),
.A2(n_242),
.B1(n_243),
.B2(n_257),
.Y(n_256)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_224),
.Y(n_257)
);

MAJIxp5_ASAP7_75t_L g224 ( 
.A(n_225),
.B(n_234),
.C(n_237),
.Y(n_224)
);

XOR2xp5_ASAP7_75t_L g282 ( 
.A(n_225),
.B(n_283),
.Y(n_282)
);

MAJIxp5_ASAP7_75t_L g225 ( 
.A(n_226),
.B(n_228),
.C(n_232),
.Y(n_225)
);

AOI22xp5_ASAP7_75t_L g306 ( 
.A1(n_226),
.A2(n_232),
.B1(n_307),
.B2(n_308),
.Y(n_306)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_226),
.Y(n_307)
);

XNOR2xp5_ASAP7_75t_L g358 ( 
.A(n_226),
.B(n_359),
.Y(n_358)
);

XOR2xp5_ASAP7_75t_L g305 ( 
.A(n_228),
.B(n_306),
.Y(n_305)
);

INVx4_ASAP7_75t_L g229 ( 
.A(n_230),
.Y(n_229)
);

BUFx6f_ASAP7_75t_L g230 ( 
.A(n_231),
.Y(n_230)
);

CKINVDCx16_ASAP7_75t_R g308 ( 
.A(n_232),
.Y(n_308)
);

INVx6_ASAP7_75t_L g416 ( 
.A(n_233),
.Y(n_416)
);

AOI22xp5_ASAP7_75t_L g283 ( 
.A1(n_234),
.A2(n_235),
.B1(n_237),
.B2(n_284),
.Y(n_283)
);

CKINVDCx14_ASAP7_75t_R g234 ( 
.A(n_235),
.Y(n_234)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_237),
.Y(n_284)
);

BUFx2_ASAP7_75t_L g238 ( 
.A(n_239),
.Y(n_238)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_240),
.Y(n_239)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_240),
.Y(n_312)
);

HB1xp67_ASAP7_75t_L g241 ( 
.A(n_242),
.Y(n_241)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_243),
.Y(n_242)
);

AOI22xp5_ASAP7_75t_SL g246 ( 
.A1(n_247),
.A2(n_249),
.B1(n_251),
.B2(n_252),
.Y(n_246)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_247),
.Y(n_251)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_249),
.Y(n_252)
);

HB1xp67_ASAP7_75t_L g293 ( 
.A(n_249),
.Y(n_293)
);

MAJIxp5_ASAP7_75t_L g291 ( 
.A(n_251),
.B(n_292),
.C(n_293),
.Y(n_291)
);

MAJIxp5_ASAP7_75t_L g253 ( 
.A(n_254),
.B(n_258),
.C(n_260),
.Y(n_253)
);

AOI22xp5_ASAP7_75t_SL g298 ( 
.A1(n_254),
.A2(n_255),
.B1(n_258),
.B2(n_299),
.Y(n_298)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_255),
.Y(n_254)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_258),
.Y(n_299)
);

INVxp67_ASAP7_75t_SL g260 ( 
.A(n_261),
.Y(n_260)
);

XNOR2xp5_ASAP7_75t_L g297 ( 
.A(n_261),
.B(n_298),
.Y(n_297)
);

MAJIxp5_ASAP7_75t_L g261 ( 
.A(n_262),
.B(n_282),
.C(n_285),
.Y(n_261)
);

XNOR2xp5_ASAP7_75t_L g302 ( 
.A(n_262),
.B(n_303),
.Y(n_302)
);

MAJIxp5_ASAP7_75t_L g262 ( 
.A(n_263),
.B(n_267),
.C(n_273),
.Y(n_262)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_264),
.Y(n_263)
);

XNOR2x1_ASAP7_75t_L g349 ( 
.A(n_264),
.B(n_350),
.Y(n_349)
);

XNOR2xp5_ASAP7_75t_L g350 ( 
.A(n_267),
.B(n_273),
.Y(n_350)
);

NAND2xp5_ASAP7_75t_L g267 ( 
.A(n_268),
.B(n_272),
.Y(n_267)
);

XOR2xp5_ASAP7_75t_L g348 ( 
.A(n_268),
.B(n_272),
.Y(n_348)
);

NOR2xp33_ASAP7_75t_L g268 ( 
.A(n_269),
.B(n_270),
.Y(n_268)
);

INVx4_ASAP7_75t_L g270 ( 
.A(n_271),
.Y(n_270)
);

INVx5_ASAP7_75t_L g322 ( 
.A(n_271),
.Y(n_322)
);

INVx3_ASAP7_75t_L g379 ( 
.A(n_271),
.Y(n_379)
);

MAJIxp5_ASAP7_75t_L g273 ( 
.A(n_274),
.B(n_277),
.C(n_279),
.Y(n_273)
);

AOI22xp5_ASAP7_75t_SL g339 ( 
.A1(n_274),
.A2(n_277),
.B1(n_340),
.B2(n_341),
.Y(n_339)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_274),
.Y(n_340)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_276),
.Y(n_275)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_277),
.Y(n_341)
);

OAI22xp5_ASAP7_75t_SL g408 ( 
.A1(n_277),
.A2(n_341),
.B1(n_409),
.B2(n_410),
.Y(n_408)
);

MAJIxp5_ASAP7_75t_L g428 ( 
.A(n_277),
.B(n_405),
.C(n_409),
.Y(n_428)
);

BUFx2_ASAP7_75t_L g395 ( 
.A(n_278),
.Y(n_395)
);

XOR2xp5_ASAP7_75t_SL g338 ( 
.A(n_279),
.B(n_339),
.Y(n_338)
);

BUFx6f_ASAP7_75t_L g280 ( 
.A(n_281),
.Y(n_280)
);

XNOR2xp5_ASAP7_75t_L g303 ( 
.A(n_282),
.B(n_285),
.Y(n_303)
);

OAI21xp5_ASAP7_75t_L g451 ( 
.A1(n_288),
.A2(n_452),
.B(n_453),
.Y(n_451)
);

AND2x2_ASAP7_75t_SL g288 ( 
.A(n_289),
.B(n_291),
.Y(n_288)
);

OR2x2_ASAP7_75t_L g453 ( 
.A(n_289),
.B(n_291),
.Y(n_453)
);

NAND2xp5_ASAP7_75t_L g294 ( 
.A(n_295),
.B(n_351),
.Y(n_294)
);

MAJIxp5_ASAP7_75t_L g295 ( 
.A(n_296),
.B(n_300),
.C(n_331),
.Y(n_295)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_297),
.Y(n_296)
);

NAND2xp5_ASAP7_75t_L g450 ( 
.A(n_297),
.B(n_301),
.Y(n_450)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_301),
.Y(n_300)
);

MAJIxp5_ASAP7_75t_L g301 ( 
.A(n_302),
.B(n_304),
.C(n_327),
.Y(n_301)
);

XOR2xp5_ASAP7_75t_L g332 ( 
.A(n_302),
.B(n_333),
.Y(n_332)
);

XNOR2xp5_ASAP7_75t_L g333 ( 
.A(n_304),
.B(n_328),
.Y(n_333)
);

MAJIxp5_ASAP7_75t_L g304 ( 
.A(n_305),
.B(n_309),
.C(n_318),
.Y(n_304)
);

XNOR2xp5_ASAP7_75t_L g336 ( 
.A(n_305),
.B(n_309),
.Y(n_336)
);

MAJIxp5_ASAP7_75t_L g386 ( 
.A(n_307),
.B(n_360),
.C(n_363),
.Y(n_386)
);

BUFx2_ASAP7_75t_L g311 ( 
.A(n_312),
.Y(n_311)
);

NOR2xp33_ASAP7_75t_L g313 ( 
.A(n_314),
.B(n_315),
.Y(n_313)
);

INVx6_ASAP7_75t_L g315 ( 
.A(n_316),
.Y(n_315)
);

BUFx12f_ASAP7_75t_L g316 ( 
.A(n_317),
.Y(n_316)
);

XOR2xp5_ASAP7_75t_L g335 ( 
.A(n_318),
.B(n_336),
.Y(n_335)
);

XNOR2xp5_ASAP7_75t_SL g436 ( 
.A(n_319),
.B(n_437),
.Y(n_436)
);

AND2x2_ASAP7_75t_L g319 ( 
.A(n_320),
.B(n_323),
.Y(n_319)
);

XNOR2x1_ASAP7_75t_SL g393 ( 
.A(n_320),
.B(n_323),
.Y(n_393)
);

INVx1_ASAP7_75t_L g400 ( 
.A(n_320),
.Y(n_400)
);

AOI22xp5_ASAP7_75t_L g417 ( 
.A1(n_320),
.A2(n_400),
.B1(n_401),
.B2(n_418),
.Y(n_417)
);

INVx2_ASAP7_75t_L g321 ( 
.A(n_322),
.Y(n_321)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_325),
.Y(n_324)
);

HB1xp67_ASAP7_75t_L g327 ( 
.A(n_328),
.Y(n_327)
);

NOR2xp67_ASAP7_75t_SL g331 ( 
.A(n_332),
.B(n_334),
.Y(n_331)
);

NAND2xp5_ASAP7_75t_L g352 ( 
.A(n_332),
.B(n_334),
.Y(n_352)
);

MAJIxp5_ASAP7_75t_L g334 ( 
.A(n_335),
.B(n_337),
.C(n_349),
.Y(n_334)
);

XNOR2xp5_ASAP7_75t_L g446 ( 
.A(n_335),
.B(n_447),
.Y(n_446)
);

XNOR2xp5_ASAP7_75t_L g447 ( 
.A(n_337),
.B(n_349),
.Y(n_447)
);

MAJIxp5_ASAP7_75t_L g337 ( 
.A(n_338),
.B(n_342),
.C(n_347),
.Y(n_337)
);

XOR2xp5_ASAP7_75t_L g441 ( 
.A(n_338),
.B(n_442),
.Y(n_441)
);

INVx1_ASAP7_75t_L g342 ( 
.A(n_343),
.Y(n_342)
);

XNOR2xp5_ASAP7_75t_L g442 ( 
.A(n_343),
.B(n_348),
.Y(n_442)
);

INVx1_ASAP7_75t_L g389 ( 
.A(n_344),
.Y(n_389)
);

XOR2x1_ASAP7_75t_L g387 ( 
.A(n_345),
.B(n_388),
.Y(n_387)
);

INVx1_ASAP7_75t_L g347 ( 
.A(n_348),
.Y(n_347)
);

NAND3xp33_ASAP7_75t_L g351 ( 
.A(n_352),
.B(n_353),
.C(n_450),
.Y(n_351)
);

OAI21xp5_ASAP7_75t_SL g353 ( 
.A1(n_354),
.A2(n_445),
.B(n_449),
.Y(n_353)
);

AOI21xp5_ASAP7_75t_L g354 ( 
.A1(n_355),
.A2(n_431),
.B(n_444),
.Y(n_354)
);

OAI21x1_ASAP7_75t_L g355 ( 
.A1(n_356),
.A2(n_396),
.B(n_430),
.Y(n_355)
);

AND2x2_ASAP7_75t_L g356 ( 
.A(n_357),
.B(n_384),
.Y(n_356)
);

OR2x2_ASAP7_75t_L g430 ( 
.A(n_357),
.B(n_384),
.Y(n_430)
);

MAJIxp5_ASAP7_75t_L g357 ( 
.A(n_358),
.B(n_367),
.C(n_376),
.Y(n_357)
);

XOR2xp5_ASAP7_75t_L g425 ( 
.A(n_358),
.B(n_426),
.Y(n_425)
);

XNOR2xp5_ASAP7_75t_L g359 ( 
.A(n_360),
.B(n_363),
.Y(n_359)
);

INVx2_ASAP7_75t_L g361 ( 
.A(n_362),
.Y(n_361)
);

INVx3_ASAP7_75t_L g364 ( 
.A(n_365),
.Y(n_364)
);

BUFx6f_ASAP7_75t_L g365 ( 
.A(n_366),
.Y(n_365)
);

AOI22xp5_ASAP7_75t_L g426 ( 
.A1(n_367),
.A2(n_368),
.B1(n_376),
.B2(n_427),
.Y(n_426)
);

INVx1_ASAP7_75t_L g367 ( 
.A(n_368),
.Y(n_367)
);

NAND2xp5_ASAP7_75t_L g368 ( 
.A(n_369),
.B(n_374),
.Y(n_368)
);

XNOR2xp5_ASAP7_75t_SL g406 ( 
.A(n_369),
.B(n_374),
.Y(n_406)
);

BUFx6f_ASAP7_75t_L g370 ( 
.A(n_371),
.Y(n_370)
);

INVx4_ASAP7_75t_L g371 ( 
.A(n_372),
.Y(n_371)
);

BUFx6f_ASAP7_75t_L g372 ( 
.A(n_373),
.Y(n_372)
);

INVx1_ASAP7_75t_L g427 ( 
.A(n_376),
.Y(n_427)
);

AO22x1_ASAP7_75t_SL g376 ( 
.A1(n_377),
.A2(n_380),
.B1(n_382),
.B2(n_383),
.Y(n_376)
);

INVx1_ASAP7_75t_L g382 ( 
.A(n_377),
.Y(n_382)
);

INVx4_ASAP7_75t_L g378 ( 
.A(n_379),
.Y(n_378)
);

INVx1_ASAP7_75t_SL g383 ( 
.A(n_380),
.Y(n_383)
);

NAND2xp5_ASAP7_75t_L g391 ( 
.A(n_380),
.B(n_382),
.Y(n_391)
);

NOR2xp33_ASAP7_75t_L g419 ( 
.A(n_383),
.B(n_420),
.Y(n_419)
);

XOR2xp5_ASAP7_75t_L g384 ( 
.A(n_385),
.B(n_390),
.Y(n_384)
);

XNOR2xp5_ASAP7_75t_L g385 ( 
.A(n_386),
.B(n_387),
.Y(n_385)
);

MAJIxp5_ASAP7_75t_L g443 ( 
.A(n_386),
.B(n_387),
.C(n_390),
.Y(n_443)
);

XOR2xp5_ASAP7_75t_L g390 ( 
.A(n_391),
.B(n_392),
.Y(n_390)
);

MAJx2_ASAP7_75t_L g439 ( 
.A(n_391),
.B(n_393),
.C(n_394),
.Y(n_439)
);

XNOR2xp5_ASAP7_75t_L g392 ( 
.A(n_393),
.B(n_394),
.Y(n_392)
);

AOI21xp5_ASAP7_75t_L g396 ( 
.A1(n_397),
.A2(n_424),
.B(n_429),
.Y(n_396)
);

OAI21xp5_ASAP7_75t_SL g397 ( 
.A1(n_398),
.A2(n_412),
.B(n_423),
.Y(n_397)
);

NOR2xp33_ASAP7_75t_L g398 ( 
.A(n_399),
.B(n_404),
.Y(n_398)
);

NAND2xp5_ASAP7_75t_L g423 ( 
.A(n_399),
.B(n_404),
.Y(n_423)
);

NOR2xp33_ASAP7_75t_SL g399 ( 
.A(n_400),
.B(n_401),
.Y(n_399)
);

INVx1_ASAP7_75t_L g418 ( 
.A(n_401),
.Y(n_418)
);

INVx1_ASAP7_75t_L g402 ( 
.A(n_403),
.Y(n_402)
);

OAI22xp5_ASAP7_75t_SL g404 ( 
.A1(n_405),
.A2(n_406),
.B1(n_407),
.B2(n_408),
.Y(n_404)
);

INVx1_ASAP7_75t_L g405 ( 
.A(n_406),
.Y(n_405)
);

INVx1_ASAP7_75t_L g407 ( 
.A(n_408),
.Y(n_407)
);

INVx1_ASAP7_75t_L g409 ( 
.A(n_410),
.Y(n_409)
);

AOI21xp5_ASAP7_75t_L g412 ( 
.A1(n_413),
.A2(n_419),
.B(n_422),
.Y(n_412)
);

NAND2xp5_ASAP7_75t_L g413 ( 
.A(n_414),
.B(n_417),
.Y(n_413)
);

NOR2xp33_ASAP7_75t_L g422 ( 
.A(n_414),
.B(n_417),
.Y(n_422)
);

INVx4_ASAP7_75t_L g415 ( 
.A(n_416),
.Y(n_415)
);

NAND2xp5_ASAP7_75t_SL g424 ( 
.A(n_425),
.B(n_428),
.Y(n_424)
);

NOR2xp33_ASAP7_75t_L g429 ( 
.A(n_425),
.B(n_428),
.Y(n_429)
);

NAND2xp5_ASAP7_75t_SL g431 ( 
.A(n_432),
.B(n_443),
.Y(n_431)
);

NOR2xp67_ASAP7_75t_SL g444 ( 
.A(n_432),
.B(n_443),
.Y(n_444)
);

AOI22xp5_ASAP7_75t_L g432 ( 
.A1(n_433),
.A2(n_434),
.B1(n_440),
.B2(n_441),
.Y(n_432)
);

INVx1_ASAP7_75t_L g433 ( 
.A(n_434),
.Y(n_433)
);

AOI22xp5_ASAP7_75t_L g434 ( 
.A1(n_435),
.A2(n_436),
.B1(n_438),
.B2(n_439),
.Y(n_434)
);

MAJIxp5_ASAP7_75t_L g448 ( 
.A(n_435),
.B(n_439),
.C(n_440),
.Y(n_448)
);

INVx1_ASAP7_75t_L g435 ( 
.A(n_436),
.Y(n_435)
);

INVx1_ASAP7_75t_L g438 ( 
.A(n_439),
.Y(n_438)
);

INVx1_ASAP7_75t_L g440 ( 
.A(n_441),
.Y(n_440)
);

NOR2xp33_ASAP7_75t_L g445 ( 
.A(n_446),
.B(n_448),
.Y(n_445)
);

NAND2xp5_ASAP7_75t_L g449 ( 
.A(n_446),
.B(n_448),
.Y(n_449)
);


endmodule