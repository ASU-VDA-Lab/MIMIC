module real_jpeg_20186_n_12 (n_5, n_4, n_8, n_0, n_319, n_1, n_11, n_2, n_6, n_7, n_3, n_10, n_9, n_12);

input n_5;
input n_4;
input n_8;
input n_0;
input n_319;
input n_1;
input n_11;
input n_2;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_12;

wire n_37;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_300;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_13;
wire n_199;
wire n_95;
wire n_238;
wire n_67;
wire n_235;
wire n_107;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_123;
wire n_50;
wire n_186;
wire n_137;
wire n_72;
wire n_171;
wire n_151;
wire n_272;
wire n_198;
wire n_203;
wire n_23;
wire n_71;
wire n_61;
wire n_99;
wire n_80;
wire n_30;
wire n_149;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_230;
wire n_128;
wire n_202;
wire n_216;
wire n_127;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_108;
wire n_233;
wire n_73;
wire n_252;
wire n_310;
wire n_78;
wire n_83;
wire n_288;
wire n_221;
wire n_104;
wire n_153;
wire n_131;
wire n_87;
wire n_40;
wire n_98;
wire n_200;
wire n_214;
wire n_113;
wire n_251;
wire n_139;
wire n_33;
wire n_175;
wire n_156;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_77;
wire n_219;
wire n_122;
wire n_19;
wire n_262;
wire n_17;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_20;
wire n_278;
wire n_314;
wire n_103;
wire n_232;
wire n_212;
wire n_284;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_213;
wire n_25;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_49;
wire n_68;
wire n_146;
wire n_286;
wire n_166;
wire n_176;
wire n_215;
wire n_312;
wire n_307;
wire n_316;
wire n_161;
wire n_207;
wire n_237;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_140;
wire n_126;
wire n_120;
wire n_155;
wire n_93;
wire n_242;
wire n_142;
wire n_76;
wire n_79;
wire n_282;
wire n_147;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_18;
wire n_145;
wire n_266;
wire n_109;
wire n_148;
wire n_196;
wire n_298;
wire n_152;
wire n_270;
wire n_159;
wire n_183;
wire n_248;
wire n_192;
wire n_90;
wire n_258;
wire n_150;
wire n_41;
wire n_74;
wire n_158;
wire n_204;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_75;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_119;
wire n_283;
wire n_181;
wire n_256;
wire n_253;
wire n_273;
wire n_16;
wire n_54;
wire n_168;
wire n_38;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_292;
wire n_64;
wire n_291;
wire n_236;
wire n_276;
wire n_287;
wire n_174;
wire n_255;
wire n_243;
wire n_299;
wire n_56;
wire n_293;
wire n_275;
wire n_227;
wire n_229;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_45;
wire n_268;
wire n_42;
wire n_313;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_143;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_303;
wire n_100;
wire n_51;
wire n_14;
wire n_205;
wire n_261;
wire n_86;
wire n_70;
wire n_32;
wire n_228;
wire n_15;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_133;
wire n_257;
wire n_210;
wire n_206;
wire n_85;
wire n_96;
wire n_308;

AOI22xp5_ASAP7_75t_L g118 ( 
.A1(n_0),
.A2(n_20),
.B1(n_21),
.B2(n_119),
.Y(n_118)
);

CKINVDCx20_ASAP7_75t_R g119 ( 
.A(n_0),
.Y(n_119)
);

OAI22xp33_ASAP7_75t_SL g123 ( 
.A1(n_0),
.A2(n_24),
.B1(n_25),
.B2(n_119),
.Y(n_123)
);

OAI22xp5_ASAP7_75t_SL g170 ( 
.A1(n_0),
.A2(n_45),
.B1(n_47),
.B2(n_119),
.Y(n_170)
);

OAI22xp33_ASAP7_75t_SL g178 ( 
.A1(n_0),
.A2(n_39),
.B1(n_40),
.B2(n_119),
.Y(n_178)
);

AOI22xp33_ASAP7_75t_SL g19 ( 
.A1(n_1),
.A2(n_20),
.B1(n_21),
.B2(n_22),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_1),
.Y(n_22)
);

AOI22xp33_ASAP7_75t_L g79 ( 
.A1(n_1),
.A2(n_22),
.B1(n_24),
.B2(n_25),
.Y(n_79)
);

AOI22xp33_ASAP7_75t_SL g107 ( 
.A1(n_1),
.A2(n_22),
.B1(n_45),
.B2(n_47),
.Y(n_107)
);

AOI22xp33_ASAP7_75t_SL g251 ( 
.A1(n_1),
.A2(n_22),
.B1(n_39),
.B2(n_40),
.Y(n_251)
);

OAI22xp33_ASAP7_75t_SL g50 ( 
.A1(n_2),
.A2(n_39),
.B1(n_40),
.B2(n_51),
.Y(n_50)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_2),
.Y(n_51)
);

OAI22xp5_ASAP7_75t_SL g58 ( 
.A1(n_2),
.A2(n_24),
.B1(n_25),
.B2(n_51),
.Y(n_58)
);

AOI21xp5_ASAP7_75t_L g74 ( 
.A1(n_2),
.A2(n_20),
.B(n_75),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_2),
.B(n_20),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_L g155 ( 
.A(n_2),
.B(n_70),
.Y(n_155)
);

AOI22xp33_ASAP7_75t_SL g160 ( 
.A1(n_2),
.A2(n_45),
.B1(n_47),
.B2(n_51),
.Y(n_160)
);

AOI21xp33_ASAP7_75t_L g174 ( 
.A1(n_2),
.A2(n_10),
.B(n_45),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_L g195 ( 
.A(n_2),
.B(n_54),
.Y(n_195)
);

O2A1O1Ixp33_ASAP7_75t_L g208 ( 
.A1(n_2),
.A2(n_24),
.B(n_56),
.C(n_209),
.Y(n_208)
);

AOI22xp5_ASAP7_75t_L g32 ( 
.A1(n_3),
.A2(n_20),
.B1(n_21),
.B2(n_33),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_3),
.Y(n_33)
);

AOI22xp33_ASAP7_75t_L g64 ( 
.A1(n_3),
.A2(n_24),
.B1(n_25),
.B2(n_33),
.Y(n_64)
);

OAI22xp5_ASAP7_75t_SL g109 ( 
.A1(n_3),
.A2(n_33),
.B1(n_45),
.B2(n_47),
.Y(n_109)
);

OAI22xp33_ASAP7_75t_SL g113 ( 
.A1(n_3),
.A2(n_33),
.B1(n_39),
.B2(n_40),
.Y(n_113)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_4),
.Y(n_20)
);

INVx6_ASAP7_75t_L g106 ( 
.A(n_5),
.Y(n_106)
);

INVx8_ASAP7_75t_L g144 ( 
.A(n_5),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_L g169 ( 
.A(n_5),
.B(n_170),
.Y(n_169)
);

BUFx12_ASAP7_75t_L g45 ( 
.A(n_6),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_7),
.Y(n_25)
);

INVx13_ASAP7_75t_L g57 ( 
.A(n_8),
.Y(n_57)
);

AOI22xp5_ASAP7_75t_L g23 ( 
.A1(n_9),
.A2(n_24),
.B1(n_25),
.B2(n_26),
.Y(n_23)
);

INVx13_ASAP7_75t_L g26 ( 
.A(n_9),
.Y(n_26)
);

NOR2xp33_ASAP7_75t_L g31 ( 
.A(n_9),
.B(n_20),
.Y(n_31)
);

O2A1O1Ixp33_ASAP7_75t_L g38 ( 
.A1(n_10),
.A2(n_39),
.B(n_43),
.C(n_44),
.Y(n_38)
);

NAND2xp5_ASAP7_75t_SL g43 ( 
.A(n_10),
.B(n_39),
.Y(n_43)
);

OAI22xp5_ASAP7_75t_L g44 ( 
.A1(n_10),
.A2(n_45),
.B1(n_46),
.B2(n_47),
.Y(n_44)
);

INVx6_ASAP7_75t_SL g46 ( 
.A(n_10),
.Y(n_46)
);

INVx11_ASAP7_75t_SL g42 ( 
.A(n_11),
.Y(n_42)
);

XOR2xp5_ASAP7_75t_L g12 ( 
.A(n_13),
.B(n_96),
.Y(n_12)
);

NAND2xp5_ASAP7_75t_SL g13 ( 
.A(n_14),
.B(n_94),
.Y(n_13)
);

NAND2xp5_ASAP7_75t_SL g14 ( 
.A(n_15),
.B(n_81),
.Y(n_14)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_15),
.B(n_81),
.Y(n_95)
);

MAJIxp5_ASAP7_75t_L g15 ( 
.A(n_16),
.B(n_68),
.C(n_76),
.Y(n_15)
);

OAI22xp5_ASAP7_75t_SL g311 ( 
.A1(n_16),
.A2(n_17),
.B1(n_68),
.B2(n_305),
.Y(n_311)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_17),
.Y(n_16)
);

AOI22xp5_ASAP7_75t_L g17 ( 
.A1(n_18),
.A2(n_34),
.B1(n_35),
.B2(n_67),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g67 ( 
.A(n_18),
.Y(n_67)
);

OAI21xp5_ASAP7_75t_L g18 ( 
.A1(n_19),
.A2(n_23),
.B(n_27),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g86 ( 
.A(n_19),
.Y(n_86)
);

INVx4_ASAP7_75t_L g21 ( 
.A(n_20),
.Y(n_21)
);

A2O1A1Ixp33_ASAP7_75t_L g29 ( 
.A1(n_20),
.A2(n_23),
.B(n_30),
.C(n_31),
.Y(n_29)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_23),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_23),
.B(n_118),
.Y(n_117)
);

AOI21xp5_ASAP7_75t_L g294 ( 
.A1(n_23),
.A2(n_29),
.B(n_74),
.Y(n_294)
);

A2O1A1Ixp33_ASAP7_75t_L g61 ( 
.A1(n_24),
.A2(n_55),
.B(n_56),
.C(n_62),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_24),
.B(n_56),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g139 ( 
.A(n_24),
.B(n_26),
.Y(n_139)
);

INVx4_ASAP7_75t_SL g24 ( 
.A(n_25),
.Y(n_24)
);

OAI22xp5_ASAP7_75t_SL g138 ( 
.A1(n_25),
.A2(n_139),
.B1(n_140),
.B2(n_141),
.Y(n_138)
);

INVx4_ASAP7_75t_L g30 ( 
.A(n_26),
.Y(n_30)
);

CKINVDCx16_ASAP7_75t_R g27 ( 
.A(n_28),
.Y(n_27)
);

NOR2xp33_ASAP7_75t_L g256 ( 
.A(n_28),
.B(n_117),
.Y(n_256)
);

NOR2xp33_ASAP7_75t_L g28 ( 
.A(n_29),
.B(n_32),
.Y(n_28)
);

NOR2xp33_ASAP7_75t_SL g73 ( 
.A(n_29),
.B(n_74),
.Y(n_73)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_29),
.Y(n_85)
);

CKINVDCx16_ASAP7_75t_R g141 ( 
.A(n_31),
.Y(n_141)
);

CKINVDCx20_ASAP7_75t_R g71 ( 
.A(n_32),
.Y(n_71)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_35),
.Y(n_34)
);

OAI22xp5_ASAP7_75t_SL g35 ( 
.A1(n_36),
.A2(n_52),
.B1(n_65),
.B2(n_66),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g65 ( 
.A(n_36),
.Y(n_65)
);

MAJIxp5_ASAP7_75t_L g92 ( 
.A(n_36),
.B(n_66),
.C(n_67),
.Y(n_92)
);

OAI22xp5_ASAP7_75t_L g150 ( 
.A1(n_36),
.A2(n_65),
.B1(n_120),
.B2(n_121),
.Y(n_150)
);

OAI22xp5_ASAP7_75t_SL g307 ( 
.A1(n_36),
.A2(n_65),
.B1(n_77),
.B2(n_308),
.Y(n_307)
);

AOI21xp5_ASAP7_75t_SL g36 ( 
.A1(n_37),
.A2(n_48),
.B(n_49),
.Y(n_36)
);

OAI21xp5_ASAP7_75t_SL g277 ( 
.A1(n_37),
.A2(n_112),
.B(n_251),
.Y(n_277)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_38),
.Y(n_37)
);

NAND2xp5_ASAP7_75t_L g114 ( 
.A(n_38),
.B(n_50),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_SL g198 ( 
.A(n_38),
.B(n_178),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_L g214 ( 
.A(n_38),
.B(n_113),
.Y(n_214)
);

AOI22xp5_ASAP7_75t_L g55 ( 
.A1(n_39),
.A2(n_40),
.B1(n_56),
.B2(n_57),
.Y(n_55)
);

OAI21xp33_ASAP7_75t_L g209 ( 
.A1(n_39),
.A2(n_51),
.B(n_57),
.Y(n_209)
);

INVx11_ASAP7_75t_L g39 ( 
.A(n_40),
.Y(n_39)
);

A2O1A1Ixp33_ASAP7_75t_L g173 ( 
.A1(n_40),
.A2(n_46),
.B(n_51),
.C(n_174),
.Y(n_173)
);

BUFx10_ASAP7_75t_L g40 ( 
.A(n_41),
.Y(n_40)
);

INVx11_ASAP7_75t_L g41 ( 
.A(n_42),
.Y(n_41)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_44),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_SL g112 ( 
.A(n_44),
.B(n_113),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_SL g177 ( 
.A(n_44),
.B(n_178),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_L g231 ( 
.A(n_44),
.B(n_50),
.Y(n_231)
);

CKINVDCx16_ASAP7_75t_R g47 ( 
.A(n_45),
.Y(n_47)
);

NAND2xp5_ASAP7_75t_L g105 ( 
.A(n_45),
.B(n_106),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g186 ( 
.A(n_47),
.B(n_187),
.Y(n_186)
);

NOR2xp33_ASAP7_75t_L g181 ( 
.A(n_48),
.B(n_51),
.Y(n_181)
);

OAI21xp5_ASAP7_75t_L g250 ( 
.A1(n_48),
.A2(n_214),
.B(n_251),
.Y(n_250)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_50),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g187 ( 
.A(n_51),
.B(n_144),
.Y(n_187)
);

CKINVDCx20_ASAP7_75t_R g66 ( 
.A(n_52),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_L g52 ( 
.A(n_53),
.B(n_59),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_L g130 ( 
.A(n_53),
.B(n_131),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_L g53 ( 
.A(n_54),
.B(n_58),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_L g122 ( 
.A(n_54),
.B(n_123),
.Y(n_122)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_55),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_SL g80 ( 
.A(n_55),
.B(n_64),
.Y(n_80)
);

AOI21xp5_ASAP7_75t_L g88 ( 
.A1(n_55),
.A2(n_61),
.B(n_89),
.Y(n_88)
);

OAI21xp5_ASAP7_75t_SL g288 ( 
.A1(n_55),
.A2(n_59),
.B(n_79),
.Y(n_288)
);

INVx11_ASAP7_75t_L g56 ( 
.A(n_57),
.Y(n_56)
);

CKINVDCx16_ASAP7_75t_R g89 ( 
.A(n_58),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g217 ( 
.A(n_58),
.B(n_60),
.Y(n_217)
);

NAND2xp5_ASAP7_75t_L g121 ( 
.A(n_59),
.B(n_122),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_SL g59 ( 
.A(n_60),
.B(n_63),
.Y(n_59)
);

AOI21xp5_ASAP7_75t_L g77 ( 
.A1(n_60),
.A2(n_78),
.B(n_80),
.Y(n_77)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_61),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_SL g132 ( 
.A(n_61),
.B(n_133),
.Y(n_132)
);

CKINVDCx14_ASAP7_75t_R g63 ( 
.A(n_64),
.Y(n_63)
);

MAJIxp5_ASAP7_75t_L g76 ( 
.A(n_65),
.B(n_68),
.C(n_77),
.Y(n_76)
);

MAJIxp5_ASAP7_75t_L g115 ( 
.A(n_65),
.B(n_116),
.C(n_120),
.Y(n_115)
);

AOI22xp5_ASAP7_75t_L g304 ( 
.A1(n_68),
.A2(n_305),
.B1(n_306),
.B2(n_307),
.Y(n_304)
);

CKINVDCx20_ASAP7_75t_R g305 ( 
.A(n_68),
.Y(n_305)
);

NAND2xp5_ASAP7_75t_L g68 ( 
.A(n_69),
.B(n_72),
.Y(n_68)
);

CKINVDCx20_ASAP7_75t_R g87 ( 
.A(n_69),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_69),
.B(n_128),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_L g69 ( 
.A(n_70),
.B(n_71),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_SL g270 ( 
.A(n_70),
.B(n_271),
.Y(n_270)
);

CKINVDCx16_ASAP7_75t_R g72 ( 
.A(n_73),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g116 ( 
.A(n_73),
.B(n_117),
.Y(n_116)
);

INVxp67_ASAP7_75t_L g271 ( 
.A(n_74),
.Y(n_271)
);

CKINVDCx14_ASAP7_75t_R g140 ( 
.A(n_75),
.Y(n_140)
);

XOR2xp5_ASAP7_75t_L g310 ( 
.A(n_76),
.B(n_311),
.Y(n_310)
);

CKINVDCx20_ASAP7_75t_R g308 ( 
.A(n_77),
.Y(n_308)
);

CKINVDCx20_ASAP7_75t_R g78 ( 
.A(n_79),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g154 ( 
.A(n_80),
.B(n_132),
.Y(n_154)
);

INVxp67_ASAP7_75t_L g273 ( 
.A(n_80),
.Y(n_273)
);

AOI22xp5_ASAP7_75t_L g81 ( 
.A1(n_82),
.A2(n_91),
.B1(n_92),
.B2(n_93),
.Y(n_81)
);

CKINVDCx20_ASAP7_75t_R g93 ( 
.A(n_82),
.Y(n_93)
);

OAI22xp5_ASAP7_75t_SL g82 ( 
.A1(n_83),
.A2(n_84),
.B1(n_88),
.B2(n_90),
.Y(n_82)
);

CKINVDCx20_ASAP7_75t_R g83 ( 
.A(n_84),
.Y(n_83)
);

AOI21xp5_ASAP7_75t_L g84 ( 
.A1(n_85),
.A2(n_86),
.B(n_87),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_SL g128 ( 
.A(n_85),
.B(n_129),
.Y(n_128)
);

CKINVDCx20_ASAP7_75t_R g90 ( 
.A(n_88),
.Y(n_90)
);

OAI22xp5_ASAP7_75t_SL g254 ( 
.A1(n_88),
.A2(n_90),
.B1(n_255),
.B2(n_256),
.Y(n_254)
);

MAJIxp5_ASAP7_75t_L g279 ( 
.A(n_90),
.B(n_253),
.C(n_256),
.Y(n_279)
);

CKINVDCx20_ASAP7_75t_R g91 ( 
.A(n_92),
.Y(n_91)
);

INVxp67_ASAP7_75t_L g94 ( 
.A(n_95),
.Y(n_94)
);

OAI321xp33_ASAP7_75t_L g96 ( 
.A1(n_97),
.A2(n_302),
.A3(n_312),
.B1(n_315),
.B2(n_316),
.C(n_319),
.Y(n_96)
);

AOI21xp5_ASAP7_75t_L g97 ( 
.A1(n_98),
.A2(n_281),
.B(n_301),
.Y(n_97)
);

OAI21xp5_ASAP7_75t_SL g98 ( 
.A1(n_99),
.A2(n_260),
.B(n_280),
.Y(n_98)
);

O2A1O1Ixp33_ASAP7_75t_SL g99 ( 
.A1(n_100),
.A2(n_161),
.B(n_243),
.C(n_259),
.Y(n_99)
);

AND2x2_ASAP7_75t_L g100 ( 
.A(n_101),
.B(n_148),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g242 ( 
.A(n_101),
.B(n_148),
.Y(n_242)
);

XOR2xp5_ASAP7_75t_L g101 ( 
.A(n_102),
.B(n_124),
.Y(n_101)
);

XOR2xp5_ASAP7_75t_L g102 ( 
.A(n_103),
.B(n_115),
.Y(n_102)
);

MAJIxp5_ASAP7_75t_L g244 ( 
.A(n_103),
.B(n_115),
.C(n_124),
.Y(n_244)
);

XOR2xp5_ASAP7_75t_L g103 ( 
.A(n_104),
.B(n_111),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_L g253 ( 
.A(n_104),
.B(n_111),
.Y(n_253)
);

OAI21xp5_ASAP7_75t_L g104 ( 
.A1(n_105),
.A2(n_107),
.B(n_108),
.Y(n_104)
);

CKINVDCx20_ASAP7_75t_R g146 ( 
.A(n_105),
.Y(n_146)
);

AOI21xp5_ASAP7_75t_L g207 ( 
.A1(n_105),
.A2(n_144),
.B(n_160),
.Y(n_207)
);

INVx5_ASAP7_75t_L g110 ( 
.A(n_106),
.Y(n_110)
);

OAI21xp5_ASAP7_75t_L g143 ( 
.A1(n_107),
.A2(n_144),
.B(n_145),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_L g157 ( 
.A(n_108),
.B(n_158),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_L g182 ( 
.A(n_108),
.B(n_183),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_SL g108 ( 
.A(n_109),
.B(n_110),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_L g145 ( 
.A(n_109),
.B(n_146),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_SL g200 ( 
.A(n_110),
.B(n_159),
.Y(n_200)
);

NAND2xp5_ASAP7_75t_L g111 ( 
.A(n_112),
.B(n_114),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_L g197 ( 
.A(n_112),
.B(n_198),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_L g176 ( 
.A(n_114),
.B(n_177),
.Y(n_176)
);

XOR2xp5_ASAP7_75t_L g149 ( 
.A(n_116),
.B(n_150),
.Y(n_149)
);

CKINVDCx20_ASAP7_75t_R g129 ( 
.A(n_118),
.Y(n_129)
);

CKINVDCx20_ASAP7_75t_R g120 ( 
.A(n_121),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_L g216 ( 
.A(n_122),
.B(n_217),
.Y(n_216)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_123),
.Y(n_133)
);

OAI22xp5_ASAP7_75t_SL g124 ( 
.A1(n_125),
.A2(n_135),
.B1(n_136),
.B2(n_147),
.Y(n_124)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_125),
.Y(n_147)
);

OAI22xp5_ASAP7_75t_SL g125 ( 
.A1(n_126),
.A2(n_127),
.B1(n_130),
.B2(n_134),
.Y(n_125)
);

MAJIxp5_ASAP7_75t_L g257 ( 
.A(n_126),
.B(n_134),
.C(n_135),
.Y(n_257)
);

CKINVDCx20_ASAP7_75t_R g126 ( 
.A(n_127),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_L g269 ( 
.A(n_128),
.B(n_270),
.Y(n_269)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_130),
.Y(n_134)
);

CKINVDCx14_ASAP7_75t_R g131 ( 
.A(n_132),
.Y(n_131)
);

CKINVDCx14_ASAP7_75t_R g135 ( 
.A(n_136),
.Y(n_135)
);

NOR2x1_ASAP7_75t_R g136 ( 
.A(n_137),
.B(n_142),
.Y(n_136)
);

AOI22xp5_ASAP7_75t_L g151 ( 
.A1(n_137),
.A2(n_138),
.B1(n_142),
.B2(n_143),
.Y(n_151)
);

CKINVDCx20_ASAP7_75t_R g137 ( 
.A(n_138),
.Y(n_137)
);

CKINVDCx20_ASAP7_75t_R g142 ( 
.A(n_143),
.Y(n_142)
);

AND2x2_ASAP7_75t_L g168 ( 
.A(n_145),
.B(n_169),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_L g249 ( 
.A(n_145),
.B(n_200),
.Y(n_249)
);

NAND2xp5_ASAP7_75t_SL g158 ( 
.A(n_146),
.B(n_159),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_L g183 ( 
.A(n_146),
.B(n_170),
.Y(n_183)
);

MAJIxp5_ASAP7_75t_L g148 ( 
.A(n_149),
.B(n_151),
.C(n_152),
.Y(n_148)
);

XOR2xp5_ASAP7_75t_L g238 ( 
.A(n_149),
.B(n_239),
.Y(n_238)
);

OAI22xp5_ASAP7_75t_SL g239 ( 
.A1(n_151),
.A2(n_152),
.B1(n_153),
.B2(n_240),
.Y(n_239)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_151),
.Y(n_240)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_153),
.Y(n_152)
);

MAJIxp5_ASAP7_75t_L g153 ( 
.A(n_154),
.B(n_155),
.C(n_156),
.Y(n_153)
);

XNOR2xp5_ASAP7_75t_SL g225 ( 
.A(n_154),
.B(n_226),
.Y(n_225)
);

AOI22xp5_ASAP7_75t_L g226 ( 
.A1(n_155),
.A2(n_156),
.B1(n_157),
.B2(n_227),
.Y(n_226)
);

CKINVDCx20_ASAP7_75t_R g227 ( 
.A(n_155),
.Y(n_227)
);

CKINVDCx20_ASAP7_75t_R g156 ( 
.A(n_157),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_L g185 ( 
.A(n_158),
.B(n_169),
.Y(n_185)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_160),
.Y(n_159)
);

NOR2xp33_ASAP7_75t_SL g161 ( 
.A(n_162),
.B(n_242),
.Y(n_161)
);

AOI21xp5_ASAP7_75t_L g162 ( 
.A1(n_163),
.A2(n_236),
.B(n_241),
.Y(n_162)
);

OAI21xp5_ASAP7_75t_SL g163 ( 
.A1(n_164),
.A2(n_221),
.B(n_235),
.Y(n_163)
);

AOI21xp5_ASAP7_75t_L g164 ( 
.A1(n_165),
.A2(n_202),
.B(n_220),
.Y(n_164)
);

OAI21xp5_ASAP7_75t_SL g165 ( 
.A1(n_166),
.A2(n_190),
.B(n_201),
.Y(n_165)
);

AOI21xp5_ASAP7_75t_L g166 ( 
.A1(n_167),
.A2(n_179),
.B(n_189),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_L g167 ( 
.A(n_168),
.B(n_171),
.Y(n_167)
);

NOR2xp33_ASAP7_75t_L g189 ( 
.A(n_168),
.B(n_171),
.Y(n_189)
);

AOI22xp5_ASAP7_75t_L g171 ( 
.A1(n_172),
.A2(n_173),
.B1(n_175),
.B2(n_176),
.Y(n_171)
);

CKINVDCx20_ASAP7_75t_R g172 ( 
.A(n_173),
.Y(n_172)
);

NOR2xp33_ASAP7_75t_SL g191 ( 
.A(n_173),
.B(n_175),
.Y(n_191)
);

CKINVDCx20_ASAP7_75t_R g175 ( 
.A(n_176),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_L g213 ( 
.A(n_177),
.B(n_214),
.Y(n_213)
);

OAI21xp5_ASAP7_75t_SL g179 ( 
.A1(n_180),
.A2(n_184),
.B(n_188),
.Y(n_179)
);

NOR2xp33_ASAP7_75t_L g180 ( 
.A(n_181),
.B(n_182),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_L g188 ( 
.A(n_181),
.B(n_182),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_L g199 ( 
.A(n_183),
.B(n_200),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_SL g184 ( 
.A(n_185),
.B(n_186),
.Y(n_184)
);

NOR2xp33_ASAP7_75t_L g190 ( 
.A(n_191),
.B(n_192),
.Y(n_190)
);

NAND2xp5_ASAP7_75t_L g201 ( 
.A(n_191),
.B(n_192),
.Y(n_201)
);

XNOR2xp5_ASAP7_75t_L g192 ( 
.A(n_193),
.B(n_199),
.Y(n_192)
);

AOI22xp5_ASAP7_75t_L g193 ( 
.A1(n_194),
.A2(n_195),
.B1(n_196),
.B2(n_197),
.Y(n_193)
);

MAJIxp5_ASAP7_75t_L g203 ( 
.A(n_194),
.B(n_197),
.C(n_199),
.Y(n_203)
);

CKINVDCx20_ASAP7_75t_R g194 ( 
.A(n_195),
.Y(n_194)
);

CKINVDCx20_ASAP7_75t_R g196 ( 
.A(n_197),
.Y(n_196)
);

NAND2xp5_ASAP7_75t_L g230 ( 
.A(n_198),
.B(n_231),
.Y(n_230)
);

NAND2xp5_ASAP7_75t_L g202 ( 
.A(n_203),
.B(n_204),
.Y(n_202)
);

NOR2xp33_ASAP7_75t_L g220 ( 
.A(n_203),
.B(n_204),
.Y(n_220)
);

AOI22xp5_ASAP7_75t_L g204 ( 
.A1(n_205),
.A2(n_211),
.B1(n_212),
.B2(n_219),
.Y(n_204)
);

CKINVDCx20_ASAP7_75t_R g219 ( 
.A(n_205),
.Y(n_219)
);

OAI22xp5_ASAP7_75t_SL g205 ( 
.A1(n_206),
.A2(n_207),
.B1(n_208),
.B2(n_210),
.Y(n_205)
);

OAI22xp5_ASAP7_75t_L g276 ( 
.A1(n_206),
.A2(n_207),
.B1(n_277),
.B2(n_278),
.Y(n_276)
);

OAI22xp5_ASAP7_75t_L g292 ( 
.A1(n_206),
.A2(n_207),
.B1(n_293),
.B2(n_294),
.Y(n_292)
);

OAI21xp5_ASAP7_75t_L g309 ( 
.A1(n_206),
.A2(n_294),
.B(n_296),
.Y(n_309)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_207),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_L g232 ( 
.A(n_207),
.B(n_208),
.Y(n_232)
);

NAND2xp5_ASAP7_75t_L g291 ( 
.A(n_207),
.B(n_277),
.Y(n_291)
);

INVxp67_ASAP7_75t_L g210 ( 
.A(n_208),
.Y(n_210)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_212),
.Y(n_211)
);

OAI22xp5_ASAP7_75t_SL g212 ( 
.A1(n_213),
.A2(n_215),
.B1(n_216),
.B2(n_218),
.Y(n_212)
);

CKINVDCx20_ASAP7_75t_R g218 ( 
.A(n_213),
.Y(n_218)
);

NAND2xp5_ASAP7_75t_L g287 ( 
.A(n_214),
.B(n_231),
.Y(n_287)
);

MAJIxp5_ASAP7_75t_L g222 ( 
.A(n_215),
.B(n_218),
.C(n_219),
.Y(n_222)
);

CKINVDCx20_ASAP7_75t_R g215 ( 
.A(n_216),
.Y(n_215)
);

NAND2xp5_ASAP7_75t_L g272 ( 
.A(n_217),
.B(n_273),
.Y(n_272)
);

NOR2xp33_ASAP7_75t_L g221 ( 
.A(n_222),
.B(n_223),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_SL g235 ( 
.A(n_222),
.B(n_223),
.Y(n_235)
);

OAI22xp5_ASAP7_75t_SL g223 ( 
.A1(n_224),
.A2(n_225),
.B1(n_228),
.B2(n_229),
.Y(n_223)
);

MAJIxp5_ASAP7_75t_L g237 ( 
.A(n_224),
.B(n_230),
.C(n_234),
.Y(n_237)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_225),
.Y(n_224)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_229),
.Y(n_228)
);

OAI22xp5_ASAP7_75t_SL g229 ( 
.A1(n_230),
.A2(n_232),
.B1(n_233),
.B2(n_234),
.Y(n_229)
);

CKINVDCx20_ASAP7_75t_R g233 ( 
.A(n_230),
.Y(n_233)
);

CKINVDCx20_ASAP7_75t_R g234 ( 
.A(n_232),
.Y(n_234)
);

NAND2xp5_ASAP7_75t_L g236 ( 
.A(n_237),
.B(n_238),
.Y(n_236)
);

NOR2xp33_ASAP7_75t_SL g241 ( 
.A(n_237),
.B(n_238),
.Y(n_241)
);

NAND2xp5_ASAP7_75t_L g243 ( 
.A(n_244),
.B(n_245),
.Y(n_243)
);

NOR2xp33_ASAP7_75t_SL g259 ( 
.A(n_244),
.B(n_245),
.Y(n_259)
);

AOI22xp5_ASAP7_75t_SL g245 ( 
.A1(n_246),
.A2(n_247),
.B1(n_257),
.B2(n_258),
.Y(n_245)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_247),
.Y(n_246)
);

XOR2xp5_ASAP7_75t_L g247 ( 
.A(n_248),
.B(n_252),
.Y(n_247)
);

MAJIxp5_ASAP7_75t_L g261 ( 
.A(n_248),
.B(n_252),
.C(n_258),
.Y(n_261)
);

XNOR2xp5_ASAP7_75t_L g248 ( 
.A(n_249),
.B(n_250),
.Y(n_248)
);

NAND2xp5_ASAP7_75t_L g266 ( 
.A(n_249),
.B(n_250),
.Y(n_266)
);

XOR2xp5_ASAP7_75t_L g252 ( 
.A(n_253),
.B(n_254),
.Y(n_252)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_256),
.Y(n_255)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_257),
.Y(n_258)
);

NOR2xp33_ASAP7_75t_L g260 ( 
.A(n_261),
.B(n_262),
.Y(n_260)
);

NAND2xp5_ASAP7_75t_SL g280 ( 
.A(n_261),
.B(n_262),
.Y(n_280)
);

XOR2xp5_ASAP7_75t_L g262 ( 
.A(n_263),
.B(n_279),
.Y(n_262)
);

OAI22xp5_ASAP7_75t_SL g263 ( 
.A1(n_264),
.A2(n_265),
.B1(n_275),
.B2(n_276),
.Y(n_263)
);

MAJIxp5_ASAP7_75t_L g282 ( 
.A(n_264),
.B(n_276),
.C(n_279),
.Y(n_282)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_265),
.Y(n_264)
);

XOR2xp5_ASAP7_75t_L g265 ( 
.A(n_266),
.B(n_267),
.Y(n_265)
);

MAJIxp5_ASAP7_75t_L g299 ( 
.A(n_266),
.B(n_268),
.C(n_274),
.Y(n_299)
);

OAI22xp5_ASAP7_75t_SL g267 ( 
.A1(n_268),
.A2(n_269),
.B1(n_272),
.B2(n_274),
.Y(n_267)
);

CKINVDCx20_ASAP7_75t_R g268 ( 
.A(n_269),
.Y(n_268)
);

CKINVDCx20_ASAP7_75t_R g274 ( 
.A(n_272),
.Y(n_274)
);

CKINVDCx16_ASAP7_75t_R g275 ( 
.A(n_276),
.Y(n_275)
);

CKINVDCx20_ASAP7_75t_R g278 ( 
.A(n_277),
.Y(n_278)
);

NAND2xp5_ASAP7_75t_L g281 ( 
.A(n_282),
.B(n_283),
.Y(n_281)
);

NOR2xp33_ASAP7_75t_SL g301 ( 
.A(n_282),
.B(n_283),
.Y(n_301)
);

AOI22xp33_ASAP7_75t_SL g283 ( 
.A1(n_284),
.A2(n_285),
.B1(n_299),
.B2(n_300),
.Y(n_283)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_285),
.Y(n_284)
);

OAI22xp5_ASAP7_75t_L g285 ( 
.A1(n_286),
.A2(n_290),
.B1(n_297),
.B2(n_298),
.Y(n_285)
);

CKINVDCx20_ASAP7_75t_R g297 ( 
.A(n_286),
.Y(n_297)
);

MAJIxp5_ASAP7_75t_L g313 ( 
.A(n_286),
.B(n_298),
.C(n_300),
.Y(n_313)
);

AOI21xp5_ASAP7_75t_L g286 ( 
.A1(n_287),
.A2(n_288),
.B(n_289),
.Y(n_286)
);

NOR2xp33_ASAP7_75t_L g289 ( 
.A(n_287),
.B(n_288),
.Y(n_289)
);

MAJIxp5_ASAP7_75t_L g303 ( 
.A(n_289),
.B(n_304),
.C(n_309),
.Y(n_303)
);

FAx1_ASAP7_75t_SL g314 ( 
.A(n_289),
.B(n_304),
.CI(n_309),
.CON(n_314),
.SN(n_314)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_290),
.Y(n_298)
);

OAI22xp5_ASAP7_75t_SL g290 ( 
.A1(n_291),
.A2(n_292),
.B1(n_295),
.B2(n_296),
.Y(n_290)
);

CKINVDCx20_ASAP7_75t_R g296 ( 
.A(n_291),
.Y(n_296)
);

CKINVDCx20_ASAP7_75t_R g295 ( 
.A(n_292),
.Y(n_295)
);

CKINVDCx20_ASAP7_75t_R g293 ( 
.A(n_294),
.Y(n_293)
);

CKINVDCx20_ASAP7_75t_R g300 ( 
.A(n_299),
.Y(n_300)
);

NOR2xp33_ASAP7_75t_L g302 ( 
.A(n_303),
.B(n_310),
.Y(n_302)
);

NAND2xp5_ASAP7_75t_L g316 ( 
.A(n_303),
.B(n_310),
.Y(n_316)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_307),
.Y(n_306)
);

NOR2xp33_ASAP7_75t_L g312 ( 
.A(n_313),
.B(n_314),
.Y(n_312)
);

NAND2xp5_ASAP7_75t_SL g315 ( 
.A(n_313),
.B(n_314),
.Y(n_315)
);

BUFx24_ASAP7_75t_SL g318 ( 
.A(n_314),
.Y(n_318)
);


endmodule