module real_aes_3623_n_360 (n_76, n_113, n_187, n_90, n_257, n_65, n_74, n_185, n_285, n_30, n_222, n_61, n_20, n_287, n_357, n_64, n_254, n_207, n_10, n_83, n_181, n_124, n_191, n_209, n_299, n_322, n_328, n_19, n_40, n_318, n_355, n_239, n_100, n_54, n_112, n_319, n_35, n_42, n_329, n_132, n_131, n_144, n_169, n_242, n_308, n_172, n_341, n_232, n_6, n_69, n_317, n_353, n_321, n_73, n_320, n_77, n_260, n_37, n_97, n_186, n_138, n_26, n_235, n_245, n_161, n_189, n_271, n_2, n_145, n_227, n_92, n_330, n_332, n_292, n_116, n_94, n_289, n_280, n_333, n_213, n_356, n_184, n_28, n_202, n_56, n_34, n_98, n_121, n_352, n_125, n_216, n_82, n_327, n_47, n_106, n_32, n_263, n_230, n_51, n_248, n_301, n_27, n_343, n_174, n_18, n_104, n_211, n_281, n_173, n_234, n_284, n_153, n_316, n_75, n_178, n_298, n_49, n_43, n_297, n_9, n_119, n_310, n_164, n_231, n_44, n_102, n_122, n_141, n_128, n_111, n_167, n_80, n_179, n_12, n_68, n_129, n_345, n_304, n_311, n_324, n_25, n_278, n_236, n_267, n_218, n_48, n_204, n_339, n_89, n_277, n_331, n_93, n_182, n_323, n_199, n_350, n_142, n_223, n_67, n_250, n_85, n_45, n_5, n_244, n_118, n_139, n_87, n_171, n_78, n_146, n_17, n_226, n_255, n_286, n_120, n_261, n_238, n_58, n_165, n_246, n_176, n_163, n_29, n_52, n_251, n_220, n_197, n_296, n_3, n_41, n_256, n_71, n_302, n_351, n_126, n_200, n_115, n_96, n_110, n_150, n_147, n_288, n_23, n_334, n_274, n_160, n_303, n_95, n_188, n_269, n_201, n_306, n_158, n_4, n_346, n_193, n_293, n_162, n_358, n_275, n_214, n_46, n_109, n_59, n_203, n_81, n_133, n_273, n_114, n_276, n_295, n_265, n_354, n_154, n_127, n_326, n_24, n_217, n_55, n_62, n_291, n_148, n_88, n_159, n_11, n_108, n_60, n_233, n_290, n_155, n_243, n_268, n_136, n_157, n_282, n_101, n_309, n_344, n_229, n_107, n_33, n_53, n_36, n_149, n_190, n_262, n_134, n_349, n_336, n_195, n_300, n_252, n_283, n_314, n_249, n_221, n_156, n_359, n_57, n_66, n_21, n_31, n_8, n_312, n_183, n_266, n_205, n_335, n_177, n_313, n_22, n_140, n_219, n_180, n_212, n_210, n_325, n_338, n_103, n_166, n_224, n_151, n_130, n_253, n_99, n_15, n_72, n_152, n_198, n_7, n_228, n_272, n_196, n_347, n_315, n_123, n_279, n_79, n_270, n_305, n_117, n_208, n_215, n_135, n_70, n_50, n_170, n_86, n_340, n_13, n_168, n_175, n_241, n_105, n_84, n_294, n_258, n_206, n_307, n_342, n_348, n_14, n_194, n_137, n_225, n_16, n_39, n_337, n_247, n_240, n_38, n_259, n_143, n_192, n_0, n_264, n_63, n_1, n_237, n_91, n_360);
input n_76;
input n_113;
input n_187;
input n_90;
input n_257;
input n_65;
input n_74;
input n_185;
input n_285;
input n_30;
input n_222;
input n_61;
input n_20;
input n_287;
input n_357;
input n_64;
input n_254;
input n_207;
input n_10;
input n_83;
input n_181;
input n_124;
input n_191;
input n_209;
input n_299;
input n_322;
input n_328;
input n_19;
input n_40;
input n_318;
input n_355;
input n_239;
input n_100;
input n_54;
input n_112;
input n_319;
input n_35;
input n_42;
input n_329;
input n_132;
input n_131;
input n_144;
input n_169;
input n_242;
input n_308;
input n_172;
input n_341;
input n_232;
input n_6;
input n_69;
input n_317;
input n_353;
input n_321;
input n_73;
input n_320;
input n_77;
input n_260;
input n_37;
input n_97;
input n_186;
input n_138;
input n_26;
input n_235;
input n_245;
input n_161;
input n_189;
input n_271;
input n_2;
input n_145;
input n_227;
input n_92;
input n_330;
input n_332;
input n_292;
input n_116;
input n_94;
input n_289;
input n_280;
input n_333;
input n_213;
input n_356;
input n_184;
input n_28;
input n_202;
input n_56;
input n_34;
input n_98;
input n_121;
input n_352;
input n_125;
input n_216;
input n_82;
input n_327;
input n_47;
input n_106;
input n_32;
input n_263;
input n_230;
input n_51;
input n_248;
input n_301;
input n_27;
input n_343;
input n_174;
input n_18;
input n_104;
input n_211;
input n_281;
input n_173;
input n_234;
input n_284;
input n_153;
input n_316;
input n_75;
input n_178;
input n_298;
input n_49;
input n_43;
input n_297;
input n_9;
input n_119;
input n_310;
input n_164;
input n_231;
input n_44;
input n_102;
input n_122;
input n_141;
input n_128;
input n_111;
input n_167;
input n_80;
input n_179;
input n_12;
input n_68;
input n_129;
input n_345;
input n_304;
input n_311;
input n_324;
input n_25;
input n_278;
input n_236;
input n_267;
input n_218;
input n_48;
input n_204;
input n_339;
input n_89;
input n_277;
input n_331;
input n_93;
input n_182;
input n_323;
input n_199;
input n_350;
input n_142;
input n_223;
input n_67;
input n_250;
input n_85;
input n_45;
input n_5;
input n_244;
input n_118;
input n_139;
input n_87;
input n_171;
input n_78;
input n_146;
input n_17;
input n_226;
input n_255;
input n_286;
input n_120;
input n_261;
input n_238;
input n_58;
input n_165;
input n_246;
input n_176;
input n_163;
input n_29;
input n_52;
input n_251;
input n_220;
input n_197;
input n_296;
input n_3;
input n_41;
input n_256;
input n_71;
input n_302;
input n_351;
input n_126;
input n_200;
input n_115;
input n_96;
input n_110;
input n_150;
input n_147;
input n_288;
input n_23;
input n_334;
input n_274;
input n_160;
input n_303;
input n_95;
input n_188;
input n_269;
input n_201;
input n_306;
input n_158;
input n_4;
input n_346;
input n_193;
input n_293;
input n_162;
input n_358;
input n_275;
input n_214;
input n_46;
input n_109;
input n_59;
input n_203;
input n_81;
input n_133;
input n_273;
input n_114;
input n_276;
input n_295;
input n_265;
input n_354;
input n_154;
input n_127;
input n_326;
input n_24;
input n_217;
input n_55;
input n_62;
input n_291;
input n_148;
input n_88;
input n_159;
input n_11;
input n_108;
input n_60;
input n_233;
input n_290;
input n_155;
input n_243;
input n_268;
input n_136;
input n_157;
input n_282;
input n_101;
input n_309;
input n_344;
input n_229;
input n_107;
input n_33;
input n_53;
input n_36;
input n_149;
input n_190;
input n_262;
input n_134;
input n_349;
input n_336;
input n_195;
input n_300;
input n_252;
input n_283;
input n_314;
input n_249;
input n_221;
input n_156;
input n_359;
input n_57;
input n_66;
input n_21;
input n_31;
input n_8;
input n_312;
input n_183;
input n_266;
input n_205;
input n_335;
input n_177;
input n_313;
input n_22;
input n_140;
input n_219;
input n_180;
input n_212;
input n_210;
input n_325;
input n_338;
input n_103;
input n_166;
input n_224;
input n_151;
input n_130;
input n_253;
input n_99;
input n_15;
input n_72;
input n_152;
input n_198;
input n_7;
input n_228;
input n_272;
input n_196;
input n_347;
input n_315;
input n_123;
input n_279;
input n_79;
input n_270;
input n_305;
input n_117;
input n_208;
input n_215;
input n_135;
input n_70;
input n_50;
input n_170;
input n_86;
input n_340;
input n_13;
input n_168;
input n_175;
input n_241;
input n_105;
input n_84;
input n_294;
input n_258;
input n_206;
input n_307;
input n_342;
input n_348;
input n_14;
input n_194;
input n_137;
input n_225;
input n_16;
input n_39;
input n_337;
input n_247;
input n_240;
input n_38;
input n_259;
input n_143;
input n_192;
input n_0;
input n_264;
input n_63;
input n_1;
input n_237;
input n_91;
output n_360;
wire n_480;
wire n_1177;
wire n_1073;
wire n_476;
wire n_758;
wire n_887;
wire n_436;
wire n_599;
wire n_684;
wire n_1066;
wire n_390;
wire n_1178;
wire n_1096;
wire n_821;
wire n_830;
wire n_624;
wire n_1018;
wire n_980;
wire n_800;
wire n_618;
wire n_778;
wire n_1205;
wire n_1106;
wire n_522;
wire n_1092;
wire n_838;
wire n_933;
wire n_1170;
wire n_485;
wire n_822;
wire n_846;
wire n_750;
wire n_631;
wire n_977;
wire n_943;
wire n_503;
wire n_905;
wire n_386;
wire n_635;
wire n_673;
wire n_1192;
wire n_518;
wire n_792;
wire n_878;
wire n_1067;
wire n_665;
wire n_991;
wire n_667;
wire n_1114;
wire n_1004;
wire n_580;
wire n_577;
wire n_469;
wire n_987;
wire n_362;
wire n_759;
wire n_979;
wire n_445;
wire n_1065;
wire n_596;
wire n_592;
wire n_540;
wire n_1064;
wire n_1075;
wire n_1197;
wire n_657;
wire n_900;
wire n_718;
wire n_841;
wire n_1129;
wire n_669;
wire n_1091;
wire n_423;
wire n_458;
wire n_1200;
wire n_444;
wire n_736;
wire n_761;
wire n_742;
wire n_364;
wire n_555;
wire n_421;
wire n_766;
wire n_852;
wire n_1113;
wire n_974;
wire n_857;
wire n_919;
wire n_1089;
wire n_1122;
wire n_461;
wire n_1047;
wire n_1016;
wire n_908;
wire n_376;
wire n_549;
wire n_571;
wire n_694;
wire n_491;
wire n_894;
wire n_923;
wire n_1034;
wire n_1123;
wire n_952;
wire n_429;
wire n_1110;
wire n_752;
wire n_448;
wire n_545;
wire n_556;
wire n_1137;
wire n_593;
wire n_460;
wire n_937;
wire n_989;
wire n_773;
wire n_401;
wire n_538;
wire n_431;
wire n_1044;
wire n_963;
wire n_865;
wire n_551;
wire n_537;
wire n_666;
wire n_884;
wire n_560;
wire n_660;
wire n_1094;
wire n_814;
wire n_944;
wire n_886;
wire n_856;
wire n_594;
wire n_1146;
wire n_983;
wire n_767;
wire n_696;
wire n_889;
wire n_955;
wire n_1147;
wire n_975;
wire n_704;
wire n_941;
wire n_453;
wire n_374;
wire n_379;
wire n_647;
wire n_932;
wire n_399;
wire n_948;
wire n_700;
wire n_1021;
wire n_677;
wire n_958;
wire n_1046;
wire n_378;
wire n_591;
wire n_775;
wire n_763;
wire n_1093;
wire n_1109;
wire n_870;
wire n_961;
wire n_489;
wire n_427;
wire n_548;
wire n_678;
wire n_415;
wire n_572;
wire n_519;
wire n_564;
wire n_638;
wire n_815;
wire n_1116;
wire n_573;
wire n_510;
wire n_1140;
wire n_1099;
wire n_709;
wire n_786;
wire n_388;
wire n_512;
wire n_395;
wire n_795;
wire n_626;
wire n_816;
wire n_400;
wire n_539;
wire n_625;
wire n_953;
wire n_462;
wire n_615;
wire n_1118;
wire n_990;
wire n_550;
wire n_966;
wire n_1160;
wire n_1108;
wire n_670;
wire n_818;
wire n_716;
wire n_918;
wire n_478;
wire n_883;
wire n_584;
wire n_896;
wire n_408;
wire n_553;
wire n_372;
wire n_994;
wire n_528;
wire n_578;
wire n_495;
wire n_892;
wire n_1078;
wire n_370;
wire n_1072;
wire n_384;
wire n_938;
wire n_744;
wire n_1128;
wire n_935;
wire n_824;
wire n_1098;
wire n_467;
wire n_875;
wire n_951;
wire n_1199;
wire n_774;
wire n_992;
wire n_813;
wire n_1213;
wire n_981;
wire n_791;
wire n_976;
wire n_466;
wire n_559;
wire n_636;
wire n_872;
wire n_1182;
wire n_906;
wire n_477;
wire n_515;
wire n_984;
wire n_1019;
wire n_680;
wire n_595;
wire n_1086;
wire n_369;
wire n_726;
wire n_1070;
wire n_1189;
wire n_1180;
wire n_517;
wire n_683;
wire n_931;
wire n_780;
wire n_840;
wire n_570;
wire n_675;
wire n_904;
wire n_920;
wire n_530;
wire n_835;
wire n_535;
wire n_732;
wire n_1117;
wire n_834;
wire n_882;
wire n_784;
wire n_496;
wire n_1210;
wire n_693;
wire n_962;
wire n_1082;
wire n_468;
wire n_746;
wire n_532;
wire n_656;
wire n_755;
wire n_1025;
wire n_1168;
wire n_1148;
wire n_409;
wire n_860;
wire n_748;
wire n_781;
wire n_523;
wire n_909;
wire n_996;
wire n_439;
wire n_1062;
wire n_576;
wire n_924;
wire n_956;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_1049;
wire n_796;
wire n_874;
wire n_1152;
wire n_801;
wire n_1126;
wire n_383;
wire n_529;
wire n_1115;
wire n_455;
wire n_504;
wire n_725;
wire n_960;
wire n_671;
wire n_973;
wire n_1081;
wire n_1084;
wire n_547;
wire n_659;
wire n_634;
wire n_682;
wire n_903;
wire n_454;
wire n_812;
wire n_782;
wire n_443;
wire n_565;
wire n_817;
wire n_760;
wire n_608;
wire n_925;
wire n_534;
wire n_708;
wire n_1029;
wire n_1020;
wire n_457;
wire n_885;
wire n_1121;
wire n_1207;
wire n_1059;
wire n_950;
wire n_381;
wire n_993;
wire n_493;
wire n_664;
wire n_367;
wire n_819;
wire n_1196;
wire n_737;
wire n_1013;
wire n_1017;
wire n_581;
wire n_610;
wire n_936;
wire n_1035;
wire n_620;
wire n_582;
wire n_641;
wire n_1063;
wire n_1135;
wire n_828;
wire n_808;
wire n_770;
wire n_940;
wire n_722;
wire n_745;
wire n_867;
wire n_398;
wire n_1193;
wire n_1100;
wire n_1167;
wire n_688;
wire n_1174;
wire n_425;
wire n_609;
wire n_1042;
wire n_879;
wire n_449;
wire n_417;
wire n_363;
wire n_607;
wire n_754;
wire n_1006;
wire n_690;
wire n_629;
wire n_1053;
wire n_1198;
wire n_499;
wire n_508;
wire n_1142;
wire n_1141;
wire n_706;
wire n_901;
wire n_561;
wire n_947;
wire n_970;
wire n_876;
wire n_437;
wire n_1112;
wire n_428;
wire n_405;
wire n_1149;
wire n_621;
wire n_368;
wire n_783;
wire n_1107;
wire n_1012;
wire n_655;
wire n_654;
wire n_502;
wire n_434;
wire n_505;
wire n_527;
wire n_769;
wire n_600;
wire n_731;
wire n_964;
wire n_1212;
wire n_605;
wire n_1054;
wire n_672;
wire n_567;
wire n_916;
wire n_406;
wire n_1050;
wire n_426;
wire n_1134;
wire n_602;
wire n_552;
wire n_402;
wire n_617;
wire n_733;
wire n_658;
wire n_676;
wire n_986;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_880;
wire n_432;
wire n_1031;
wire n_1037;
wire n_1131;
wire n_1103;
wire n_1008;
wire n_807;
wire n_1011;
wire n_416;
wire n_790;
wire n_895;
wire n_832;
wire n_410;
wire n_799;
wire n_805;
wire n_751;
wire n_490;
wire n_913;
wire n_999;
wire n_619;
wire n_391;
wire n_1095;
wire n_1060;
wire n_859;
wire n_695;
wire n_1181;
wire n_685;
wire n_881;
wire n_1154;
wire n_1080;
wire n_361;
wire n_917;
wire n_632;
wire n_768;
wire n_412;
wire n_542;
wire n_645;
wire n_1145;
wire n_557;
wire n_714;
wire n_777;
wire n_985;
wire n_1077;
wire n_488;
wire n_501;
wire n_1041;
wire n_1111;
wire n_910;
wire n_869;
wire n_613;
wire n_642;
wire n_387;
wire n_1125;
wire n_957;
wire n_995;
wire n_1124;
wire n_702;
wire n_954;
wire n_969;
wire n_912;
wire n_1009;
wire n_1007;
wire n_1202;
wire n_464;
wire n_1163;
wire n_945;
wire n_604;
wire n_734;
wire n_898;
wire n_848;
wire n_392;
wire n_562;
wire n_1022;
wire n_404;
wire n_598;
wire n_713;
wire n_735;
wire n_728;
wire n_756;
wire n_1179;
wire n_1201;
wire n_569;
wire n_997;
wire n_563;
wire n_1203;
wire n_785;
wire n_1171;
wire n_891;
wire n_430;
wire n_568;
wire n_413;
wire n_471;
wire n_902;
wire n_1105;
wire n_1157;
wire n_1158;
wire n_1132;
wire n_853;
wire n_810;
wire n_843;
wire n_1079;
wire n_579;
wire n_1033;
wire n_699;
wire n_533;
wire n_1028;
wire n_1014;
wire n_1000;
wire n_1003;
wire n_1187;
wire n_366;
wire n_727;
wire n_1083;
wire n_649;
wire n_385;
wire n_397;
wire n_663;
wire n_749;
wire n_588;
wire n_536;
wire n_914;
wire n_707;
wire n_622;
wire n_470;
wire n_851;
wire n_915;
wire n_1002;
wire n_1155;
wire n_934;
wire n_1165;
wire n_494;
wire n_1001;
wire n_711;
wire n_864;
wire n_1027;
wire n_1169;
wire n_377;
wire n_1058;
wire n_1139;
wire n_927;
wire n_1038;
wire n_965;
wire n_723;
wire n_662;
wire n_1085;
wire n_382;
wire n_845;
wire n_850;
wire n_1043;
wire n_1136;
wire n_720;
wire n_968;
wire n_972;
wire n_435;
wire n_1127;
wire n_1026;
wire n_511;
wire n_484;
wire n_893;
wire n_492;
wire n_1068;
wire n_509;
wire n_407;
wire n_419;
wire n_730;
wire n_1023;
wire n_643;
wire n_747;
wire n_1204;
wire n_486;
wire n_930;
wire n_1209;
wire n_1057;
wire n_411;
wire n_697;
wire n_978;
wire n_847;
wire n_907;
wire n_779;
wire n_481;
wire n_498;
wire n_691;
wire n_765;
wire n_826;
wire n_648;
wire n_373;
wire n_589;
wire n_628;
wire n_939;
wire n_1005;
wire n_487;
wire n_831;
wire n_653;
wire n_365;
wire n_526;
wire n_637;
wire n_899;
wire n_928;
wire n_692;
wire n_544;
wire n_789;
wire n_1087;
wire n_1051;
wire n_1194;
wire n_389;
wire n_738;
wire n_701;
wire n_827;
wire n_809;
wire n_482;
wire n_633;
wire n_520;
wire n_922;
wire n_679;
wire n_926;
wire n_942;
wire n_1048;
wire n_472;
wire n_1120;
wire n_971;
wire n_866;
wire n_452;
wire n_787;
wire n_1052;
wire n_1071;
wire n_630;
wire n_1214;
wire n_806;
wire n_689;
wire n_820;
wire n_1097;
wire n_959;
wire n_715;
wire n_1208;
wire n_946;
wire n_420;
wire n_612;
wire n_858;
wire n_873;
wire n_1130;
wire n_438;
wire n_764;
wire n_794;
wire n_741;
wire n_753;
wire n_1188;
wire n_623;
wire n_1032;
wire n_446;
wire n_721;
wire n_681;
wire n_982;
wire n_456;
wire n_717;
wire n_1090;
wire n_1133;
wire n_1164;
wire n_712;
wire n_1183;
wire n_433;
wire n_516;
wire n_627;
wire n_739;
wire n_418;
wire n_521;
wire n_422;
wire n_771;
wire n_524;
wire n_861;
wire n_1162;
wire n_705;
wire n_1191;
wire n_1206;
wire n_1195;
wire n_575;
wire n_762;
wire n_479;
wire n_442;
wire n_825;
wire n_740;
wire n_371;
wire n_698;
wire n_541;
wire n_839;
wire n_639;
wire n_546;
wire n_587;
wire n_1186;
wire n_1010;
wire n_811;
wire n_1015;
wire n_459;
wire n_558;
wire n_1172;
wire n_863;
wire n_998;
wire n_1175;
wire n_724;
wire n_440;
wire n_525;
wire n_1074;
wire n_644;
wire n_674;
wire n_836;
wire n_888;
wire n_793;
wire n_1150;
wire n_1184;
wire n_1166;
wire n_1056;
wire n_583;
wire n_833;
wire n_414;
wire n_757;
wire n_1161;
wire n_929;
wire n_1143;
wire n_686;
wire n_776;
wire n_1190;
wire n_1138;
wire n_803;
wire n_890;
wire n_543;
wire n_497;
wire n_514;
wire n_507;
wire n_949;
wire n_614;
wire n_586;
wire n_911;
wire n_772;
wire n_450;
wire n_788;
wire n_441;
wire n_585;
wire n_465;
wire n_473;
wire n_967;
wire n_566;
wire n_719;
wire n_837;
wire n_1045;
wire n_871;
wire n_474;
wire n_1156;
wire n_1159;
wire n_829;
wire n_1030;
wire n_988;
wire n_1088;
wire n_1055;
wire n_921;
wire n_375;
wire n_597;
wire n_640;
wire n_483;
wire n_611;
wire n_1176;
wire n_1151;
wire n_380;
wire n_1036;
wire n_394;
wire n_687;
wire n_729;
wire n_844;
wire n_646;
wire n_650;
wire n_710;
wire n_743;
wire n_823;
wire n_393;
wire n_652;
wire n_703;
wire n_1040;
wire n_500;
wire n_601;
wire n_1101;
wire n_661;
wire n_463;
wire n_1076;
wire n_396;
wire n_804;
wire n_1102;
wire n_447;
wire n_1185;
wire n_1211;
wire n_1173;
wire n_603;
wire n_854;
wire n_403;
wire n_424;
wire n_877;
wire n_802;
wire n_868;
wire n_1039;
wire n_1119;
wire n_574;
wire n_1069;
wire n_1024;
wire n_842;
wire n_1104;
wire n_1144;
wire n_849;
wire n_1061;
wire n_554;
wire n_475;
wire n_897;
wire n_1153;
wire n_855;
wire n_798;
wire n_668;
wire n_797;
wire n_862;
AOI22xp33_ASAP7_75t_L g903 ( .A1(n_0), .A2(n_254), .B1(n_633), .B2(n_634), .Y(n_903) );
AOI22xp33_ASAP7_75t_L g955 ( .A1(n_1), .A2(n_344), .B1(n_506), .B2(n_507), .Y(n_955) );
AOI22xp33_ASAP7_75t_L g803 ( .A1(n_2), .A2(n_78), .B1(n_519), .B2(n_658), .Y(n_803) );
AOI22xp33_ASAP7_75t_L g902 ( .A1(n_3), .A2(n_183), .B1(n_682), .B2(n_683), .Y(n_902) );
AOI22xp5_ASAP7_75t_L g484 ( .A1(n_4), .A2(n_190), .B1(n_485), .B2(n_486), .Y(n_484) );
AOI22xp33_ASAP7_75t_L g505 ( .A1(n_5), .A2(n_144), .B1(n_506), .B2(n_507), .Y(n_505) );
AOI22xp33_ASAP7_75t_L g681 ( .A1(n_6), .A2(n_306), .B1(n_682), .B2(n_683), .Y(n_681) );
AOI22xp33_ASAP7_75t_L g882 ( .A1(n_7), .A2(n_157), .B1(n_606), .B2(n_774), .Y(n_882) );
INVx1_ASAP7_75t_L g850 ( .A(n_8), .Y(n_850) );
AOI22xp33_ASAP7_75t_L g515 ( .A1(n_9), .A2(n_320), .B1(n_434), .B2(n_516), .Y(n_515) );
AOI22xp5_ASAP7_75t_L g528 ( .A1(n_10), .A2(n_290), .B1(n_529), .B2(n_530), .Y(n_528) );
AOI22xp33_ASAP7_75t_L g775 ( .A1(n_11), .A2(n_27), .B1(n_557), .B2(n_614), .Y(n_775) );
AOI22xp33_ASAP7_75t_L g656 ( .A1(n_12), .A2(n_108), .B1(n_435), .B2(n_485), .Y(n_656) );
NAND2xp5_ASAP7_75t_SL g401 ( .A(n_13), .B(n_389), .Y(n_401) );
AOI22xp33_ASAP7_75t_L g660 ( .A1(n_14), .A2(n_187), .B1(n_530), .B2(n_661), .Y(n_660) );
CKINVDCx20_ASAP7_75t_R g884 ( .A(n_15), .Y(n_884) );
AOI22xp5_ASAP7_75t_L g966 ( .A1(n_16), .A2(n_326), .B1(n_967), .B2(n_971), .Y(n_966) );
AOI22xp33_ASAP7_75t_L g842 ( .A1(n_17), .A2(n_236), .B1(n_506), .B2(n_507), .Y(n_842) );
AOI22xp33_ASAP7_75t_L g603 ( .A1(n_18), .A2(n_160), .B1(n_551), .B2(n_604), .Y(n_603) );
AOI22xp5_ASAP7_75t_L g637 ( .A1(n_19), .A2(n_196), .B1(n_509), .B2(n_510), .Y(n_637) );
NAND2xp5_ASAP7_75t_L g785 ( .A(n_20), .B(n_786), .Y(n_785) );
BUFx6f_ASAP7_75t_L g389 ( .A(n_21), .Y(n_389) );
AOI22xp33_ASAP7_75t_L g445 ( .A1(n_22), .A2(n_324), .B1(n_446), .B2(n_449), .Y(n_445) );
AOI22xp5_ASAP7_75t_L g784 ( .A1(n_23), .A2(n_68), .B1(n_572), .B2(n_595), .Y(n_784) );
AOI22xp5_ASAP7_75t_L g525 ( .A1(n_24), .A2(n_143), .B1(n_383), .B2(n_526), .Y(n_525) );
AOI21xp5_ASAP7_75t_L g807 ( .A1(n_25), .A2(n_808), .B(n_809), .Y(n_807) );
AOI22xp33_ASAP7_75t_L g707 ( .A1(n_26), .A2(n_38), .B1(n_708), .B2(n_709), .Y(n_707) );
AOI22xp33_ASAP7_75t_L g799 ( .A1(n_28), .A2(n_137), .B1(n_524), .B2(n_800), .Y(n_799) );
AOI22xp33_ASAP7_75t_L g573 ( .A1(n_29), .A2(n_211), .B1(n_574), .B2(n_575), .Y(n_573) );
INVx1_ASAP7_75t_L g770 ( .A(n_30), .Y(n_770) );
INVx1_ASAP7_75t_L g564 ( .A(n_31), .Y(n_564) );
AOI22xp33_ASAP7_75t_L g949 ( .A1(n_32), .A2(n_199), .B1(n_503), .B2(n_628), .Y(n_949) );
AOI22xp33_ASAP7_75t_L g943 ( .A1(n_33), .A2(n_100), .B1(n_510), .B2(n_634), .Y(n_943) );
AOI22xp33_ASAP7_75t_L g612 ( .A1(n_34), .A2(n_195), .B1(n_613), .B2(n_614), .Y(n_612) );
AOI22xp33_ASAP7_75t_L g508 ( .A1(n_35), .A2(n_357), .B1(n_509), .B2(n_510), .Y(n_508) );
XOR2x2_ASAP7_75t_L g623 ( .A(n_36), .B(n_624), .Y(n_623) );
AOI22xp33_ASAP7_75t_SL g899 ( .A1(n_37), .A2(n_347), .B1(n_446), .B2(n_503), .Y(n_899) );
AOI22xp33_ASAP7_75t_L g753 ( .A1(n_39), .A2(n_142), .B1(n_440), .B2(n_516), .Y(n_753) );
INVx1_ASAP7_75t_L g825 ( .A(n_40), .Y(n_825) );
AOI22xp33_ASAP7_75t_L g452 ( .A1(n_41), .A2(n_148), .B1(n_453), .B2(n_455), .Y(n_452) );
AOI22xp33_ASAP7_75t_L g919 ( .A1(n_42), .A2(n_129), .B1(n_530), .B2(n_661), .Y(n_919) );
AOI22xp5_ASAP7_75t_L g797 ( .A1(n_43), .A2(n_93), .B1(n_602), .B2(n_798), .Y(n_797) );
AOI22xp33_ASAP7_75t_L g752 ( .A1(n_44), .A2(n_154), .B1(n_438), .B2(n_549), .Y(n_752) );
AOI22xp33_ASAP7_75t_L g821 ( .A1(n_45), .A2(n_165), .B1(n_424), .B2(n_523), .Y(n_821) );
AOI22xp33_ASAP7_75t_L g941 ( .A1(n_46), .A2(n_105), .B1(n_506), .B2(n_507), .Y(n_941) );
AOI22xp33_ASAP7_75t_L g954 ( .A1(n_47), .A2(n_225), .B1(n_682), .B2(n_683), .Y(n_954) );
AOI22xp33_ASAP7_75t_L g550 ( .A1(n_48), .A2(n_177), .B1(n_551), .B2(n_552), .Y(n_550) );
AOI22xp33_ASAP7_75t_L g951 ( .A1(n_49), .A2(n_249), .B1(n_598), .B2(n_639), .Y(n_951) );
OA22x2_ASAP7_75t_L g395 ( .A1(n_50), .A2(n_152), .B1(n_389), .B2(n_393), .Y(n_395) );
INVx1_ASAP7_75t_L g415 ( .A(n_50), .Y(n_415) );
AOI22xp33_ASAP7_75t_L g818 ( .A1(n_51), .A2(n_296), .B1(n_383), .B2(n_408), .Y(n_818) );
XNOR2x1_ASAP7_75t_L g794 ( .A(n_52), .B(n_795), .Y(n_794) );
AOI22xp33_ASAP7_75t_L g733 ( .A1(n_53), .A2(n_61), .B1(n_734), .B2(n_735), .Y(n_733) );
AOI22xp33_ASAP7_75t_L g1097 ( .A1(n_54), .A2(n_201), .B1(n_994), .B2(n_1007), .Y(n_1097) );
AOI22xp33_ASAP7_75t_L g641 ( .A1(n_55), .A2(n_58), .B1(n_506), .B2(n_507), .Y(n_641) );
AOI22xp5_ASAP7_75t_L g635 ( .A1(n_56), .A2(n_286), .B1(n_485), .B2(n_486), .Y(n_635) );
AOI22xp33_ASAP7_75t_L g531 ( .A1(n_57), .A2(n_343), .B1(n_532), .B2(n_533), .Y(n_531) );
AOI22xp33_ASAP7_75t_L g437 ( .A1(n_59), .A2(n_252), .B1(n_438), .B2(n_440), .Y(n_437) );
AOI22xp33_ASAP7_75t_L g1016 ( .A1(n_60), .A2(n_180), .B1(n_974), .B2(n_977), .Y(n_1016) );
AOI22xp33_ASAP7_75t_L g640 ( .A1(n_62), .A2(n_245), .B1(n_500), .B2(n_502), .Y(n_640) );
AOI22xp33_ASAP7_75t_L g1197 ( .A1(n_63), .A2(n_289), .B1(n_506), .B2(n_507), .Y(n_1197) );
AOI22xp33_ASAP7_75t_L g428 ( .A1(n_64), .A2(n_255), .B1(n_429), .B2(n_434), .Y(n_428) );
INVx1_ASAP7_75t_L g744 ( .A(n_65), .Y(n_744) );
AOI22xp33_ASAP7_75t_L g925 ( .A1(n_66), .A2(n_104), .B1(n_429), .B2(n_486), .Y(n_925) );
AOI22xp33_ASAP7_75t_L g1195 ( .A1(n_67), .A2(n_257), .B1(n_509), .B2(n_510), .Y(n_1195) );
AOI221xp5_ASAP7_75t_L g625 ( .A1(n_69), .A2(n_173), .B1(n_626), .B2(n_627), .C(n_629), .Y(n_625) );
NOR2xp33_ASAP7_75t_L g370 ( .A(n_70), .B(n_167), .Y(n_370) );
INVx1_ASAP7_75t_L g392 ( .A(n_70), .Y(n_392) );
OAI21xp33_ASAP7_75t_L g416 ( .A1(n_70), .A2(n_152), .B(n_417), .Y(n_416) );
AOI21xp33_ASAP7_75t_L g781 ( .A1(n_71), .A2(n_574), .B(n_782), .Y(n_781) );
AO221x2_ASAP7_75t_L g992 ( .A1(n_72), .A2(n_327), .B1(n_974), .B2(n_981), .C(n_993), .Y(n_992) );
AOI221xp5_ASAP7_75t_L g664 ( .A1(n_73), .A2(n_299), .B1(n_476), .B2(n_574), .C(n_665), .Y(n_664) );
AOI22xp33_ASAP7_75t_L g904 ( .A1(n_74), .A2(n_338), .B1(n_506), .B2(n_507), .Y(n_904) );
AOI22xp33_ASAP7_75t_L g501 ( .A1(n_75), .A2(n_287), .B1(n_502), .B2(n_503), .Y(n_501) );
AOI22xp33_ASAP7_75t_L g601 ( .A1(n_76), .A2(n_138), .B1(n_526), .B2(n_602), .Y(n_601) );
AOI22xp33_ASAP7_75t_L g776 ( .A1(n_77), .A2(n_267), .B1(n_551), .B2(n_552), .Y(n_776) );
INVx1_ASAP7_75t_L g1193 ( .A(n_79), .Y(n_1193) );
AOI22xp5_ASAP7_75t_L g924 ( .A1(n_80), .A2(n_171), .B1(n_602), .B2(n_654), .Y(n_924) );
AOI22xp33_ASAP7_75t_L g596 ( .A1(n_81), .A2(n_145), .B1(n_597), .B2(n_598), .Y(n_596) );
AOI22xp33_ASAP7_75t_SL g777 ( .A1(n_82), .A2(n_202), .B1(n_526), .B2(n_602), .Y(n_777) );
AOI22xp33_ASAP7_75t_L g569 ( .A1(n_83), .A2(n_318), .B1(n_570), .B2(n_572), .Y(n_569) );
INVx1_ASAP7_75t_L g468 ( .A(n_84), .Y(n_468) );
AOI22xp5_ASAP7_75t_L g987 ( .A1(n_85), .A2(n_315), .B1(n_977), .B2(n_988), .Y(n_987) );
AOI22xp33_ASAP7_75t_L g711 ( .A1(n_86), .A2(n_122), .B1(n_613), .B2(n_614), .Y(n_711) );
AOI22xp33_ASAP7_75t_L g1006 ( .A1(n_87), .A2(n_331), .B1(n_967), .B2(n_1007), .Y(n_1006) );
NAND2xp5_ASAP7_75t_L g827 ( .A(n_88), .B(n_828), .Y(n_827) );
NAND2xp5_ASAP7_75t_L g750 ( .A(n_89), .B(n_533), .Y(n_750) );
AND2x4_ASAP7_75t_L g970 ( .A(n_90), .B(n_266), .Y(n_970) );
INVx1_ASAP7_75t_L g976 ( .A(n_90), .Y(n_976) );
HB1xp67_ASAP7_75t_L g1213 ( .A(n_90), .Y(n_1213) );
AOI22xp33_ASAP7_75t_L g901 ( .A1(n_91), .A2(n_302), .B1(n_509), .B2(n_510), .Y(n_901) );
AOI22xp33_ASAP7_75t_L g756 ( .A1(n_92), .A2(n_232), .B1(n_526), .B2(n_757), .Y(n_756) );
AOI22xp33_ASAP7_75t_L g875 ( .A1(n_94), .A2(n_194), .B1(n_598), .B2(n_676), .Y(n_875) );
INVx1_ASAP7_75t_L g540 ( .A(n_95), .Y(n_540) );
AO22x1_ASAP7_75t_L g993 ( .A1(n_95), .A2(n_179), .B1(n_971), .B2(n_994), .Y(n_993) );
AOI22xp33_ASAP7_75t_L g802 ( .A1(n_96), .A2(n_209), .B1(n_516), .B2(n_604), .Y(n_802) );
CKINVDCx20_ASAP7_75t_R g726 ( .A(n_97), .Y(n_726) );
AOI22xp5_ASAP7_75t_L g773 ( .A1(n_98), .A2(n_99), .B1(n_554), .B2(n_774), .Y(n_773) );
AOI22xp33_ASAP7_75t_L g499 ( .A1(n_101), .A2(n_185), .B1(n_465), .B2(n_500), .Y(n_499) );
AOI22xp5_ASAP7_75t_L g990 ( .A1(n_102), .A2(n_131), .B1(n_983), .B2(n_991), .Y(n_990) );
AOI221xp5_ASAP7_75t_L g534 ( .A1(n_103), .A2(n_106), .B1(n_493), .B2(n_535), .C(n_536), .Y(n_534) );
AOI21xp5_ASAP7_75t_L g823 ( .A1(n_107), .A2(n_639), .B(n_824), .Y(n_823) );
XNOR2x1_ASAP7_75t_L g739 ( .A(n_109), .B(n_740), .Y(n_739) );
AOI21xp5_ASAP7_75t_L g492 ( .A1(n_110), .A2(n_493), .B(n_496), .Y(n_492) );
AOI22xp33_ASAP7_75t_L g942 ( .A1(n_111), .A2(n_307), .B1(n_639), .B2(n_682), .Y(n_942) );
NAND2xp5_ASAP7_75t_L g917 ( .A(n_112), .B(n_918), .Y(n_917) );
AOI21xp5_ASAP7_75t_L g560 ( .A1(n_113), .A2(n_561), .B(n_563), .Y(n_560) );
AOI22xp33_ASAP7_75t_L g806 ( .A1(n_114), .A2(n_191), .B1(n_530), .B2(n_661), .Y(n_806) );
AOI22xp5_ASAP7_75t_L g879 ( .A1(n_115), .A2(n_140), .B1(n_880), .B2(n_881), .Y(n_879) );
AOI22xp33_ASAP7_75t_L g1190 ( .A1(n_116), .A2(n_166), .B1(n_500), .B2(n_503), .Y(n_1190) );
INVx1_ASAP7_75t_L g537 ( .A(n_117), .Y(n_537) );
AOI22xp33_ASAP7_75t_L g382 ( .A1(n_118), .A2(n_132), .B1(n_383), .B2(n_408), .Y(n_382) );
INVx1_ASAP7_75t_L g969 ( .A(n_119), .Y(n_969) );
AND2x4_ASAP7_75t_L g972 ( .A(n_119), .B(n_366), .Y(n_972) );
INVx1_ASAP7_75t_SL g989 ( .A(n_119), .Y(n_989) );
AOI22xp33_ASAP7_75t_L g674 ( .A1(n_120), .A2(n_253), .B1(n_465), .B2(n_530), .Y(n_674) );
XNOR2x2_ASAP7_75t_SL g834 ( .A(n_121), .B(n_835), .Y(n_834) );
AOI22xp33_ASAP7_75t_L g877 ( .A1(n_123), .A2(n_272), .B1(n_552), .B2(n_878), .Y(n_877) );
INVx1_ASAP7_75t_L g686 ( .A(n_124), .Y(n_686) );
AOI22xp33_ASAP7_75t_L g1015 ( .A1(n_125), .A2(n_149), .B1(n_967), .B2(n_971), .Y(n_1015) );
NAND2xp5_ASAP7_75t_L g475 ( .A(n_126), .B(n_476), .Y(n_475) );
AOI22xp33_ASAP7_75t_L g926 ( .A1(n_127), .A2(n_261), .B1(n_440), .B2(n_519), .Y(n_926) );
AOI22xp33_ASAP7_75t_L g1189 ( .A1(n_128), .A2(n_342), .B1(n_502), .B2(n_639), .Y(n_1189) );
AOI221xp5_ASAP7_75t_L g853 ( .A1(n_130), .A2(n_350), .B1(n_627), .B2(n_854), .C(n_855), .Y(n_853) );
XNOR2x1_ASAP7_75t_L g481 ( .A(n_131), .B(n_482), .Y(n_481) );
OAI22x1_ASAP7_75t_L g583 ( .A1(n_133), .A2(n_584), .B1(n_620), .B2(n_621), .Y(n_583) );
NAND3xp33_ASAP7_75t_SL g620 ( .A(n_133), .B(n_600), .C(n_615), .Y(n_620) );
INVx1_ASAP7_75t_L g490 ( .A(n_134), .Y(n_490) );
AOI22xp33_ASAP7_75t_L g684 ( .A1(n_135), .A2(n_164), .B1(n_633), .B2(n_634), .Y(n_684) );
AOI22xp5_ASAP7_75t_L g678 ( .A1(n_136), .A2(n_348), .B1(n_506), .B2(n_507), .Y(n_678) );
AOI21xp5_ASAP7_75t_L g920 ( .A1(n_139), .A2(n_574), .B(n_921), .Y(n_920) );
INVx1_ASAP7_75t_L g845 ( .A(n_141), .Y(n_845) );
INVx1_ASAP7_75t_L g666 ( .A(n_146), .Y(n_666) );
AOI22xp33_ASAP7_75t_L g662 ( .A1(n_147), .A2(n_221), .B1(n_575), .B2(n_663), .Y(n_662) );
INVx1_ASAP7_75t_L g577 ( .A(n_149), .Y(n_577) );
AOI22xp5_ASAP7_75t_L g679 ( .A1(n_150), .A2(n_334), .B1(n_509), .B2(n_510), .Y(n_679) );
INVx1_ASAP7_75t_L g407 ( .A(n_151), .Y(n_407) );
NAND2xp5_ASAP7_75t_L g460 ( .A(n_151), .B(n_206), .Y(n_460) );
NAND2xp5_ASAP7_75t_L g474 ( .A(n_151), .B(n_413), .Y(n_474) );
NOR2xp33_ASAP7_75t_L g369 ( .A(n_152), .B(n_274), .Y(n_369) );
AOI22xp33_ASAP7_75t_L g1094 ( .A1(n_153), .A2(n_217), .B1(n_1004), .B2(n_1095), .Y(n_1094) );
INVx1_ASAP7_75t_L g783 ( .A(n_155), .Y(n_783) );
AOI22xp5_ASAP7_75t_L g829 ( .A1(n_156), .A2(n_270), .B1(n_529), .B2(n_830), .Y(n_829) );
OAI22xp5_ASAP7_75t_L g1205 ( .A1(n_158), .A2(n_1186), .B1(n_1206), .B2(n_1207), .Y(n_1205) );
CKINVDCx5p33_ASAP7_75t_R g1206 ( .A(n_158), .Y(n_1206) );
AOI22xp5_ASAP7_75t_L g522 ( .A1(n_159), .A2(n_233), .B1(n_523), .B2(n_524), .Y(n_522) );
AOI221xp5_ASAP7_75t_L g758 ( .A1(n_161), .A2(n_168), .B1(n_535), .B2(n_759), .C(n_761), .Y(n_758) );
INVx1_ASAP7_75t_L g922 ( .A(n_162), .Y(n_922) );
AOI21xp5_ASAP7_75t_L g892 ( .A1(n_163), .A2(n_562), .B(n_893), .Y(n_892) );
NAND2xp5_ASAP7_75t_L g399 ( .A(n_167), .B(n_400), .Y(n_399) );
AOI22xp33_ASAP7_75t_L g837 ( .A1(n_169), .A2(n_200), .B1(n_438), .B2(n_440), .Y(n_837) );
AOI22xp33_ASAP7_75t_L g956 ( .A1(n_170), .A2(n_251), .B1(n_633), .B2(n_634), .Y(n_956) );
AOI22xp33_ASAP7_75t_L g927 ( .A1(n_172), .A2(n_358), .B1(n_523), .B2(n_524), .Y(n_927) );
AOI22xp33_ASAP7_75t_L g755 ( .A1(n_174), .A2(n_359), .B1(n_524), .B2(n_554), .Y(n_755) );
AO22x2_ASAP7_75t_L g886 ( .A1(n_175), .A2(n_887), .B1(n_905), .B2(n_906), .Y(n_886) );
INVxp67_ASAP7_75t_SL g905 ( .A(n_175), .Y(n_905) );
INVx1_ASAP7_75t_L g497 ( .A(n_176), .Y(n_497) );
AOI22xp5_ASAP7_75t_L g592 ( .A1(n_178), .A2(n_239), .B1(n_593), .B2(n_595), .Y(n_592) );
INVx1_ASAP7_75t_L g810 ( .A(n_181), .Y(n_810) );
AOI22xp33_ASAP7_75t_L g518 ( .A1(n_182), .A2(n_288), .B1(n_519), .B2(n_520), .Y(n_518) );
NAND2xp5_ASAP7_75t_L g847 ( .A(n_184), .B(n_812), .Y(n_847) );
NAND2xp5_ASAP7_75t_L g813 ( .A(n_186), .B(n_814), .Y(n_813) );
AOI22xp33_ASAP7_75t_L g916 ( .A1(n_188), .A2(n_336), .B1(n_529), .B2(n_663), .Y(n_916) );
AOI22xp33_ASAP7_75t_L g652 ( .A1(n_189), .A2(n_193), .B1(n_653), .B2(n_654), .Y(n_652) );
AOI21xp33_ASAP7_75t_L g464 ( .A1(n_192), .A2(n_465), .B(n_467), .Y(n_464) );
XNOR2x1_ASAP7_75t_L g815 ( .A(n_197), .B(n_816), .Y(n_815) );
BUFx2_ASAP7_75t_L g895 ( .A(n_198), .Y(n_895) );
INVx1_ASAP7_75t_L g762 ( .A(n_203), .Y(n_762) );
AOI22xp5_ASAP7_75t_L g487 ( .A1(n_204), .A2(n_333), .B1(n_438), .B2(n_488), .Y(n_487) );
AOI22xp5_ASAP7_75t_L g980 ( .A1(n_205), .A2(n_226), .B1(n_974), .B2(n_981), .Y(n_980) );
INVx1_ASAP7_75t_L g390 ( .A(n_206), .Y(n_390) );
AOI22xp33_ASAP7_75t_L g556 ( .A1(n_207), .A2(n_244), .B1(n_557), .B2(n_558), .Y(n_556) );
AOI22xp33_ASAP7_75t_L g418 ( .A1(n_208), .A2(n_321), .B1(n_419), .B2(n_424), .Y(n_418) );
NAND2xp5_ASAP7_75t_L g587 ( .A(n_210), .B(n_588), .Y(n_587) );
AOI22xp33_ASAP7_75t_L g712 ( .A1(n_212), .A2(n_355), .B1(n_555), .B2(n_606), .Y(n_712) );
AOI22xp33_ASAP7_75t_L g998 ( .A1(n_213), .A2(n_301), .B1(n_974), .B2(n_977), .Y(n_998) );
AOI22xp33_ASAP7_75t_L g553 ( .A1(n_214), .A2(n_243), .B1(n_554), .B2(n_555), .Y(n_553) );
XNOR2x1_ASAP7_75t_L g930 ( .A(n_215), .B(n_931), .Y(n_930) );
AOI22xp33_ASAP7_75t_L g787 ( .A1(n_216), .A2(n_330), .B1(n_597), .B2(n_788), .Y(n_787) );
AOI22xp33_ASAP7_75t_L g805 ( .A1(n_218), .A2(n_328), .B1(n_529), .B2(n_532), .Y(n_805) );
AOI22xp5_ASAP7_75t_L g973 ( .A1(n_219), .A2(n_260), .B1(n_974), .B2(n_977), .Y(n_973) );
AOI22xp33_ASAP7_75t_L g657 ( .A1(n_220), .A2(n_300), .B1(n_519), .B2(n_658), .Y(n_657) );
AOI22xp5_ASAP7_75t_L g675 ( .A1(n_222), .A2(n_231), .B1(n_453), .B2(n_676), .Y(n_675) );
NAND2xp5_ASAP7_75t_L g933 ( .A(n_223), .B(n_562), .Y(n_933) );
CKINVDCx20_ASAP7_75t_R g720 ( .A(n_224), .Y(n_720) );
AOI22xp33_ASAP7_75t_L g819 ( .A1(n_227), .A2(n_311), .B1(n_429), .B2(n_434), .Y(n_819) );
AOI22xp33_ASAP7_75t_L g1003 ( .A1(n_228), .A2(n_298), .B1(n_974), .B2(n_1004), .Y(n_1003) );
OR2x2_ASAP7_75t_L g443 ( .A(n_229), .B(n_444), .Y(n_443) );
INVxp67_ASAP7_75t_L g480 ( .A(n_229), .Y(n_480) );
AOI22xp33_ASAP7_75t_L g997 ( .A1(n_229), .A2(n_294), .B1(n_971), .B2(n_994), .Y(n_997) );
AOI22xp33_ASAP7_75t_L g883 ( .A1(n_230), .A2(n_284), .B1(n_520), .B2(n_551), .Y(n_883) );
AOI22xp5_ASAP7_75t_L g632 ( .A1(n_234), .A2(n_256), .B1(n_633), .B2(n_634), .Y(n_632) );
AOI22xp33_ASAP7_75t_L g841 ( .A1(n_235), .A2(n_283), .B1(n_682), .B2(n_683), .Y(n_841) );
NAND2xp5_ASAP7_75t_SL g950 ( .A(n_237), .B(n_590), .Y(n_950) );
AOI22xp5_ASAP7_75t_L g982 ( .A1(n_238), .A2(n_323), .B1(n_967), .B2(n_983), .Y(n_982) );
AOI22xp5_ASAP7_75t_L g651 ( .A1(n_240), .A2(n_241), .B1(n_523), .B2(n_555), .Y(n_651) );
AOI22xp33_ASAP7_75t_L g870 ( .A1(n_242), .A2(n_303), .B1(n_574), .B2(n_871), .Y(n_870) );
CKINVDCx20_ASAP7_75t_R g730 ( .A(n_246), .Y(n_730) );
AOI22xp33_ASAP7_75t_L g935 ( .A1(n_247), .A2(n_279), .B1(n_500), .B2(n_502), .Y(n_935) );
AOI22xp33_ASAP7_75t_L g820 ( .A1(n_248), .A2(n_280), .B1(n_438), .B2(n_440), .Y(n_820) );
AOI22xp33_ASAP7_75t_L g838 ( .A1(n_250), .A2(n_341), .B1(n_653), .B2(n_839), .Y(n_838) );
AOI22xp33_ASAP7_75t_L g948 ( .A1(n_258), .A2(n_269), .B1(n_500), .B2(n_502), .Y(n_948) );
NAND2xp5_ASAP7_75t_L g566 ( .A(n_259), .B(n_567), .Y(n_566) );
AOI22xp33_ASAP7_75t_L g867 ( .A1(n_262), .A2(n_354), .B1(n_868), .B2(n_869), .Y(n_867) );
AOI22xp33_ASAP7_75t_L g940 ( .A1(n_263), .A2(n_291), .B1(n_633), .B2(n_683), .Y(n_940) );
INVx1_ASAP7_75t_L g852 ( .A(n_264), .Y(n_852) );
AOI22x1_ASAP7_75t_L g647 ( .A1(n_265), .A2(n_648), .B1(n_649), .B2(n_667), .Y(n_647) );
INVx1_ASAP7_75t_L g667 ( .A(n_265), .Y(n_667) );
HB1xp67_ASAP7_75t_L g371 ( .A(n_266), .Y(n_371) );
AND2x4_ASAP7_75t_L g975 ( .A(n_266), .B(n_976), .Y(n_975) );
AOI22xp33_ASAP7_75t_L g1198 ( .A1(n_268), .A2(n_295), .B1(n_633), .B2(n_634), .Y(n_1198) );
INVx1_ASAP7_75t_L g746 ( .A(n_271), .Y(n_746) );
AOI22xp33_ASAP7_75t_L g638 ( .A1(n_273), .A2(n_314), .B1(n_503), .B2(n_639), .Y(n_638) );
INVx1_ASAP7_75t_L g405 ( .A(n_274), .Y(n_405) );
INVxp67_ASAP7_75t_L g463 ( .A(n_274), .Y(n_463) );
AOI21xp33_ASAP7_75t_SL g889 ( .A1(n_275), .A2(n_465), .B(n_890), .Y(n_889) );
INVx1_ASAP7_75t_L g630 ( .A(n_276), .Y(n_630) );
INVx1_ASAP7_75t_L g691 ( .A(n_277), .Y(n_691) );
INVx1_ASAP7_75t_L g945 ( .A(n_278), .Y(n_945) );
AOI22xp5_ASAP7_75t_SL g615 ( .A1(n_281), .A2(n_325), .B1(n_616), .B2(n_618), .Y(n_615) );
AOI22xp33_ASAP7_75t_L g1196 ( .A1(n_282), .A2(n_297), .B1(n_682), .B2(n_683), .Y(n_1196) );
INVx2_ASAP7_75t_L g366 ( .A(n_285), .Y(n_366) );
AOI22xp5_ASAP7_75t_L g934 ( .A1(n_292), .A2(n_293), .B1(n_503), .B2(n_509), .Y(n_934) );
INVx1_ASAP7_75t_L g856 ( .A(n_304), .Y(n_856) );
INVx1_ASAP7_75t_L g891 ( .A(n_305), .Y(n_891) );
AOI21xp33_ASAP7_75t_L g936 ( .A1(n_308), .A2(n_628), .B(n_937), .Y(n_936) );
INVx1_ASAP7_75t_L g938 ( .A(n_309), .Y(n_938) );
INVx1_ASAP7_75t_L g748 ( .A(n_310), .Y(n_748) );
NAND2xp5_ASAP7_75t_L g872 ( .A(n_312), .B(n_873), .Y(n_872) );
AOI22xp5_ASAP7_75t_L g605 ( .A1(n_313), .A2(n_349), .B1(n_606), .B2(n_608), .Y(n_605) );
AOI22xp33_ASAP7_75t_L g826 ( .A1(n_316), .A2(n_332), .B1(n_446), .B2(n_530), .Y(n_826) );
INVx1_ASAP7_75t_L g913 ( .A(n_317), .Y(n_913) );
CKINVDCx20_ASAP7_75t_R g724 ( .A(n_319), .Y(n_724) );
AOI22xp33_ASAP7_75t_L g953 ( .A1(n_322), .A2(n_353), .B1(n_509), .B2(n_510), .Y(n_953) );
INVx1_ASAP7_75t_L g1185 ( .A(n_323), .Y(n_1185) );
AOI22xp33_ASAP7_75t_L g1204 ( .A1(n_323), .A2(n_1205), .B1(n_1208), .B2(n_1210), .Y(n_1204) );
XNOR2x2_ASAP7_75t_L g705 ( .A(n_326), .B(n_706), .Y(n_705) );
AOI22xp33_ASAP7_75t_L g713 ( .A1(n_329), .A2(n_346), .B1(n_551), .B2(n_552), .Y(n_713) );
INVx1_ASAP7_75t_L g692 ( .A(n_335), .Y(n_692) );
BUFx2_ASAP7_75t_L g897 ( .A(n_337), .Y(n_897) );
NAND2xp5_ASAP7_75t_L g1188 ( .A(n_339), .B(n_590), .Y(n_1188) );
AOI22xp33_ASAP7_75t_L g548 ( .A1(n_340), .A2(n_356), .B1(n_526), .B2(n_549), .Y(n_548) );
AOI21xp5_ASAP7_75t_L g689 ( .A1(n_345), .A2(n_495), .B(n_690), .Y(n_689) );
AOI21xp33_ASAP7_75t_L g1191 ( .A1(n_351), .A2(n_628), .B(n_1192), .Y(n_1191) );
CKINVDCx20_ASAP7_75t_R g716 ( .A(n_352), .Y(n_716) );
AOI21xp5_ASAP7_75t_L g360 ( .A1(n_361), .A2(n_372), .B(n_959), .Y(n_360) );
INVx1_ASAP7_75t_L g361 ( .A(n_362), .Y(n_361) );
BUFx4_ASAP7_75t_SL g362 ( .A(n_363), .Y(n_362) );
NAND3xp33_ASAP7_75t_L g363 ( .A(n_364), .B(n_367), .C(n_371), .Y(n_363) );
AND2x2_ASAP7_75t_L g1201 ( .A(n_364), .B(n_1202), .Y(n_1201) );
AND2x2_ASAP7_75t_L g1209 ( .A(n_364), .B(n_1203), .Y(n_1209) );
AOI21xp5_ASAP7_75t_L g1214 ( .A1(n_364), .A2(n_371), .B(n_989), .Y(n_1214) );
INVx1_ASAP7_75t_L g364 ( .A(n_365), .Y(n_364) );
AO21x1_ASAP7_75t_L g1211 ( .A1(n_365), .A2(n_1212), .B(n_1214), .Y(n_1211) );
HB1xp67_ASAP7_75t_L g365 ( .A(n_366), .Y(n_365) );
AND2x2_ASAP7_75t_L g968 ( .A(n_366), .B(n_969), .Y(n_968) );
AND3x4_ASAP7_75t_L g988 ( .A(n_366), .B(n_975), .C(n_989), .Y(n_988) );
NOR2xp33_ASAP7_75t_L g1202 ( .A(n_367), .B(n_1203), .Y(n_1202) );
HB1xp67_ASAP7_75t_L g367 ( .A(n_368), .Y(n_367) );
AO21x2_ASAP7_75t_L g471 ( .A1(n_368), .A2(n_472), .B(n_473), .Y(n_471) );
NAND2xp5_ASAP7_75t_L g368 ( .A(n_369), .B(n_370), .Y(n_368) );
INVx1_ASAP7_75t_L g1203 ( .A(n_371), .Y(n_1203) );
OAI22xp5_ASAP7_75t_L g372 ( .A1(n_373), .A2(n_374), .B1(n_699), .B2(n_700), .Y(n_372) );
INVx1_ASAP7_75t_L g373 ( .A(n_374), .Y(n_373) );
OA22x2_ASAP7_75t_L g374 ( .A1(n_375), .A2(n_376), .B1(n_579), .B2(n_580), .Y(n_374) );
INVx1_ASAP7_75t_L g375 ( .A(n_376), .Y(n_375) );
XNOR2xp5_ASAP7_75t_L g376 ( .A(n_377), .B(n_543), .Y(n_376) );
AO22x2_ASAP7_75t_L g377 ( .A1(n_378), .A2(n_511), .B1(n_541), .B2(n_542), .Y(n_377) );
INVx2_ASAP7_75t_L g542 ( .A(n_378), .Y(n_542) );
XNOR2x1_ASAP7_75t_L g378 ( .A(n_379), .B(n_481), .Y(n_378) );
OAI22x1_ASAP7_75t_L g379 ( .A1(n_380), .A2(n_443), .B1(n_479), .B2(n_480), .Y(n_379) );
HB1xp67_ASAP7_75t_L g380 ( .A(n_381), .Y(n_380) );
NOR2xp33_ASAP7_75t_L g479 ( .A(n_381), .B(n_444), .Y(n_479) );
NAND4xp25_ASAP7_75t_L g381 ( .A(n_382), .B(n_418), .C(n_428), .D(n_437), .Y(n_381) );
BUFx3_ASAP7_75t_L g881 ( .A(n_383), .Y(n_881) );
BUFx6f_ASAP7_75t_L g383 ( .A(n_384), .Y(n_383) );
BUFx6f_ASAP7_75t_L g549 ( .A(n_384), .Y(n_549) );
BUFx6f_ASAP7_75t_L g602 ( .A(n_384), .Y(n_602) );
BUFx6f_ASAP7_75t_L g653 ( .A(n_384), .Y(n_653) );
AND2x4_ASAP7_75t_L g384 ( .A(n_385), .B(n_396), .Y(n_384) );
AND2x4_ASAP7_75t_L g421 ( .A(n_385), .B(n_422), .Y(n_421) );
AND2x2_ASAP7_75t_L g425 ( .A(n_385), .B(n_426), .Y(n_425) );
AND2x4_ASAP7_75t_L g439 ( .A(n_385), .B(n_432), .Y(n_439) );
AND2x4_ASAP7_75t_L g506 ( .A(n_385), .B(n_422), .Y(n_506) );
AND2x4_ASAP7_75t_L g507 ( .A(n_385), .B(n_426), .Y(n_507) );
AND2x4_ASAP7_75t_L g509 ( .A(n_385), .B(n_436), .Y(n_509) );
AND2x4_ASAP7_75t_L g633 ( .A(n_385), .B(n_432), .Y(n_633) );
AND2x4_ASAP7_75t_L g385 ( .A(n_386), .B(n_394), .Y(n_385) );
AND2x2_ASAP7_75t_L g448 ( .A(n_386), .B(n_395), .Y(n_448) );
INVx1_ASAP7_75t_L g386 ( .A(n_387), .Y(n_386) );
AND2x2_ASAP7_75t_L g431 ( .A(n_387), .B(n_395), .Y(n_431) );
NAND2xp5_ASAP7_75t_L g387 ( .A(n_388), .B(n_391), .Y(n_387) );
NAND2xp33_ASAP7_75t_L g388 ( .A(n_389), .B(n_390), .Y(n_388) );
INVx2_ASAP7_75t_L g393 ( .A(n_389), .Y(n_393) );
INVx3_ASAP7_75t_L g400 ( .A(n_389), .Y(n_400) );
NAND2xp33_ASAP7_75t_L g406 ( .A(n_389), .B(n_407), .Y(n_406) );
INVx1_ASAP7_75t_L g417 ( .A(n_389), .Y(n_417) );
HB1xp67_ASAP7_75t_L g459 ( .A(n_389), .Y(n_459) );
NAND2xp5_ASAP7_75t_L g414 ( .A(n_390), .B(n_415), .Y(n_414) );
NAND2xp5_ASAP7_75t_L g391 ( .A(n_392), .B(n_393), .Y(n_391) );
OAI21xp5_ASAP7_75t_L g462 ( .A1(n_392), .A2(n_417), .B(n_463), .Y(n_462) );
INVx1_ASAP7_75t_L g394 ( .A(n_395), .Y(n_394) );
AND2x2_ASAP7_75t_L g461 ( .A(n_395), .B(n_462), .Y(n_461) );
AND2x4_ASAP7_75t_L g410 ( .A(n_396), .B(n_411), .Y(n_410) );
AND2x4_ASAP7_75t_L g510 ( .A(n_396), .B(n_411), .Y(n_510) );
AND2x4_ASAP7_75t_L g683 ( .A(n_396), .B(n_431), .Y(n_683) );
INVx2_ASAP7_75t_L g396 ( .A(n_397), .Y(n_396) );
INVx2_ASAP7_75t_L g436 ( .A(n_397), .Y(n_436) );
OR2x2_ASAP7_75t_L g397 ( .A(n_398), .B(n_402), .Y(n_397) );
AND2x4_ASAP7_75t_L g422 ( .A(n_398), .B(n_423), .Y(n_422) );
INVx2_ASAP7_75t_L g427 ( .A(n_398), .Y(n_427) );
AND2x4_ASAP7_75t_L g432 ( .A(n_398), .B(n_433), .Y(n_432) );
AND2x2_ASAP7_75t_L g457 ( .A(n_398), .B(n_458), .Y(n_457) );
AND2x4_ASAP7_75t_L g398 ( .A(n_399), .B(n_401), .Y(n_398) );
NAND2xp5_ASAP7_75t_L g404 ( .A(n_400), .B(n_405), .Y(n_404) );
INVxp67_ASAP7_75t_L g413 ( .A(n_400), .Y(n_413) );
NAND3xp33_ASAP7_75t_L g473 ( .A(n_401), .B(n_412), .C(n_474), .Y(n_473) );
INVx1_ASAP7_75t_L g433 ( .A(n_402), .Y(n_433) );
INVx1_ASAP7_75t_L g402 ( .A(n_403), .Y(n_402) );
INVx1_ASAP7_75t_L g423 ( .A(n_403), .Y(n_423) );
AND2x2_ASAP7_75t_L g403 ( .A(n_404), .B(n_406), .Y(n_403) );
HB1xp67_ASAP7_75t_L g709 ( .A(n_408), .Y(n_709) );
INVx5_ASAP7_75t_L g408 ( .A(n_409), .Y(n_408) );
INVx2_ASAP7_75t_L g654 ( .A(n_409), .Y(n_654) );
INVx1_ASAP7_75t_L g798 ( .A(n_409), .Y(n_798) );
INVx3_ASAP7_75t_L g839 ( .A(n_409), .Y(n_839) );
INVx1_ASAP7_75t_L g878 ( .A(n_409), .Y(n_878) );
INVx6_ASAP7_75t_L g409 ( .A(n_410), .Y(n_409) );
BUFx12f_ASAP7_75t_L g526 ( .A(n_410), .Y(n_526) );
AND2x4_ASAP7_75t_L g442 ( .A(n_411), .B(n_432), .Y(n_442) );
AND2x4_ASAP7_75t_L g451 ( .A(n_411), .B(n_426), .Y(n_451) );
AND2x4_ASAP7_75t_L g503 ( .A(n_411), .B(n_426), .Y(n_503) );
AND2x4_ASAP7_75t_L g634 ( .A(n_411), .B(n_432), .Y(n_634) );
AND2x2_ASAP7_75t_L g411 ( .A(n_412), .B(n_416), .Y(n_411) );
NAND2xp5_ASAP7_75t_L g412 ( .A(n_413), .B(n_414), .Y(n_412) );
INVx1_ASAP7_75t_L g419 ( .A(n_420), .Y(n_419) );
INVx2_ASAP7_75t_L g607 ( .A(n_420), .Y(n_607) );
INVx1_ASAP7_75t_L g800 ( .A(n_420), .Y(n_800) );
INVx3_ASAP7_75t_L g420 ( .A(n_421), .Y(n_420) );
BUFx12f_ASAP7_75t_L g523 ( .A(n_421), .Y(n_523) );
BUFx6f_ASAP7_75t_L g554 ( .A(n_421), .Y(n_554) );
AND2x2_ASAP7_75t_L g454 ( .A(n_422), .B(n_431), .Y(n_454) );
AND2x4_ASAP7_75t_L g466 ( .A(n_422), .B(n_448), .Y(n_466) );
AND2x4_ASAP7_75t_L g502 ( .A(n_422), .B(n_431), .Y(n_502) );
AND2x4_ASAP7_75t_L g639 ( .A(n_422), .B(n_448), .Y(n_639) );
AND2x4_ASAP7_75t_L g426 ( .A(n_423), .B(n_427), .Y(n_426) );
BUFx3_ASAP7_75t_L g424 ( .A(n_425), .Y(n_424) );
BUFx6f_ASAP7_75t_L g524 ( .A(n_425), .Y(n_524) );
BUFx5_ASAP7_75t_L g555 ( .A(n_425), .Y(n_555) );
INVx1_ASAP7_75t_L g611 ( .A(n_425), .Y(n_611) );
AND2x4_ASAP7_75t_L g447 ( .A(n_426), .B(n_448), .Y(n_447) );
AND2x2_ASAP7_75t_L g478 ( .A(n_426), .B(n_431), .Y(n_478) );
AND2x2_ASAP7_75t_L g495 ( .A(n_426), .B(n_431), .Y(n_495) );
AND2x2_ASAP7_75t_L g628 ( .A(n_426), .B(n_448), .Y(n_628) );
BUFx4f_ASAP7_75t_L g429 ( .A(n_430), .Y(n_429) );
BUFx6f_ASAP7_75t_L g485 ( .A(n_430), .Y(n_485) );
AND2x2_ASAP7_75t_L g430 ( .A(n_431), .B(n_432), .Y(n_430) );
AND2x4_ASAP7_75t_L g435 ( .A(n_431), .B(n_436), .Y(n_435) );
AND2x2_ASAP7_75t_L g517 ( .A(n_431), .B(n_432), .Y(n_517) );
AND2x4_ASAP7_75t_L g682 ( .A(n_431), .B(n_432), .Y(n_682) );
BUFx6f_ASAP7_75t_L g434 ( .A(n_435), .Y(n_434) );
BUFx6f_ASAP7_75t_L g486 ( .A(n_435), .Y(n_486) );
BUFx3_ASAP7_75t_L g552 ( .A(n_435), .Y(n_552) );
BUFx6f_ASAP7_75t_L g604 ( .A(n_435), .Y(n_604) );
BUFx12f_ASAP7_75t_L g757 ( .A(n_435), .Y(n_757) );
BUFx12f_ASAP7_75t_L g613 ( .A(n_438), .Y(n_613) );
BUFx6f_ASAP7_75t_L g880 ( .A(n_438), .Y(n_880) );
BUFx12f_ASAP7_75t_L g438 ( .A(n_439), .Y(n_438) );
BUFx6f_ASAP7_75t_L g519 ( .A(n_439), .Y(n_519) );
BUFx6f_ASAP7_75t_L g557 ( .A(n_439), .Y(n_557) );
INVx2_ASAP7_75t_L g440 ( .A(n_441), .Y(n_440) );
INVx1_ASAP7_75t_L g488 ( .A(n_441), .Y(n_488) );
INVx4_ASAP7_75t_L g520 ( .A(n_441), .Y(n_520) );
INVx1_ASAP7_75t_L g558 ( .A(n_441), .Y(n_558) );
INVx4_ASAP7_75t_L g614 ( .A(n_441), .Y(n_614) );
INVx4_ASAP7_75t_L g658 ( .A(n_441), .Y(n_658) );
INVx8_ASAP7_75t_L g441 ( .A(n_442), .Y(n_441) );
NAND4xp25_ASAP7_75t_L g444 ( .A(n_445), .B(n_452), .C(n_464), .D(n_475), .Y(n_444) );
INVx2_ASAP7_75t_L g491 ( .A(n_446), .Y(n_491) );
BUFx3_ASAP7_75t_L g868 ( .A(n_446), .Y(n_868) );
BUFx6f_ASAP7_75t_L g446 ( .A(n_447), .Y(n_446) );
BUFx3_ASAP7_75t_L g535 ( .A(n_447), .Y(n_535) );
INVx2_ASAP7_75t_L g571 ( .A(n_447), .Y(n_571) );
BUFx6f_ASAP7_75t_L g661 ( .A(n_447), .Y(n_661) );
BUFx8_ASAP7_75t_SL g688 ( .A(n_447), .Y(n_688) );
INVx2_ASAP7_75t_L g449 ( .A(n_450), .Y(n_449) );
INVx3_ASAP7_75t_L g450 ( .A(n_451), .Y(n_450) );
BUFx6f_ASAP7_75t_L g530 ( .A(n_451), .Y(n_530) );
BUFx6f_ASAP7_75t_L g572 ( .A(n_451), .Y(n_572) );
INVx3_ASAP7_75t_L g743 ( .A(n_453), .Y(n_743) );
BUFx6f_ASAP7_75t_L g453 ( .A(n_454), .Y(n_453) );
BUFx3_ASAP7_75t_L g529 ( .A(n_454), .Y(n_529) );
INVx2_ASAP7_75t_L g576 ( .A(n_454), .Y(n_576) );
BUFx2_ASAP7_75t_L g455 ( .A(n_456), .Y(n_455) );
BUFx4f_ASAP7_75t_L g533 ( .A(n_456), .Y(n_533) );
INVx5_ASAP7_75t_L g565 ( .A(n_456), .Y(n_565) );
BUFx2_ASAP7_75t_L g830 ( .A(n_456), .Y(n_830) );
AND2x4_ASAP7_75t_L g456 ( .A(n_457), .B(n_461), .Y(n_456) );
AND2x2_ASAP7_75t_L g500 ( .A(n_457), .B(n_461), .Y(n_500) );
AND2x4_ASAP7_75t_L g812 ( .A(n_457), .B(n_461), .Y(n_812) );
NAND2xp5_ASAP7_75t_L g458 ( .A(n_459), .B(n_460), .Y(n_458) );
INVx1_ASAP7_75t_L g472 ( .A(n_459), .Y(n_472) );
INVx2_ASAP7_75t_L g619 ( .A(n_465), .Y(n_619) );
BUFx3_ASAP7_75t_L g465 ( .A(n_466), .Y(n_465) );
BUFx3_ASAP7_75t_L g532 ( .A(n_466), .Y(n_532) );
BUFx6f_ASAP7_75t_L g574 ( .A(n_466), .Y(n_574) );
INVx1_ASAP7_75t_L g719 ( .A(n_466), .Y(n_719) );
NOR2xp33_ASAP7_75t_L g467 ( .A(n_468), .B(n_469), .Y(n_467) );
NOR2xp33_ASAP7_75t_L g496 ( .A(n_469), .B(n_497), .Y(n_496) );
INVx1_ASAP7_75t_L g814 ( .A(n_469), .Y(n_814) );
NOR2xp33_ASAP7_75t_L g824 ( .A(n_469), .B(n_825), .Y(n_824) );
NOR2xp33_ASAP7_75t_L g855 ( .A(n_469), .B(n_856), .Y(n_855) );
BUFx6f_ASAP7_75t_L g469 ( .A(n_470), .Y(n_469) );
BUFx6f_ASAP7_75t_L g568 ( .A(n_470), .Y(n_568) );
BUFx6f_ASAP7_75t_L g470 ( .A(n_471), .Y(n_470) );
INVx3_ASAP7_75t_L g539 ( .A(n_471), .Y(n_539) );
INVx2_ASAP7_75t_L g476 ( .A(n_477), .Y(n_476) );
INVx2_ASAP7_75t_L g626 ( .A(n_477), .Y(n_626) );
INVx3_ASAP7_75t_SL g732 ( .A(n_477), .Y(n_732) );
INVx2_ASAP7_75t_L g828 ( .A(n_477), .Y(n_828) );
INVx2_ASAP7_75t_L g918 ( .A(n_477), .Y(n_918) );
INVx3_ASAP7_75t_L g477 ( .A(n_478), .Y(n_477) );
BUFx3_ASAP7_75t_L g562 ( .A(n_478), .Y(n_562) );
INVx2_ASAP7_75t_L g591 ( .A(n_478), .Y(n_591) );
INVx1_ASAP7_75t_L g578 ( .A(n_481), .Y(n_578) );
NAND4xp75_ASAP7_75t_L g482 ( .A(n_483), .B(n_489), .C(n_498), .D(n_504), .Y(n_482) );
AND2x2_ASAP7_75t_L g483 ( .A(n_484), .B(n_487), .Y(n_483) );
OA21x2_ASAP7_75t_L g489 ( .A1(n_490), .A2(n_491), .B(n_492), .Y(n_489) );
INVx2_ASAP7_75t_L g493 ( .A(n_494), .Y(n_493) );
INVx2_ASAP7_75t_L g494 ( .A(n_495), .Y(n_494) );
HB1xp67_ASAP7_75t_L g854 ( .A(n_495), .Y(n_854) );
AND2x2_ASAP7_75t_L g498 ( .A(n_499), .B(n_501), .Y(n_498) );
INVx1_ASAP7_75t_L g849 ( .A(n_502), .Y(n_849) );
INVx2_ASAP7_75t_L g898 ( .A(n_502), .Y(n_898) );
INVx2_ASAP7_75t_L g851 ( .A(n_503), .Y(n_851) );
AND2x2_ASAP7_75t_L g504 ( .A(n_505), .B(n_508), .Y(n_504) );
BUFx3_ASAP7_75t_L g511 ( .A(n_512), .Y(n_511) );
INVx1_ASAP7_75t_L g541 ( .A(n_512), .Y(n_541) );
XNOR2x1_ASAP7_75t_L g512 ( .A(n_513), .B(n_540), .Y(n_512) );
NAND4xp75_ASAP7_75t_L g513 ( .A(n_514), .B(n_521), .C(n_527), .D(n_534), .Y(n_513) );
AND2x2_ASAP7_75t_L g514 ( .A(n_515), .B(n_518), .Y(n_514) );
BUFx6f_ASAP7_75t_L g516 ( .A(n_517), .Y(n_516) );
BUFx8_ASAP7_75t_L g551 ( .A(n_517), .Y(n_551) );
AND2x2_ASAP7_75t_L g521 ( .A(n_522), .B(n_525), .Y(n_521) );
AND2x2_ASAP7_75t_L g527 ( .A(n_528), .B(n_531), .Y(n_527) );
INVx2_ASAP7_75t_L g617 ( .A(n_529), .Y(n_617) );
BUFx3_ASAP7_75t_L g728 ( .A(n_530), .Y(n_728) );
INVx3_ASAP7_75t_L g745 ( .A(n_530), .Y(n_745) );
INVx2_ASAP7_75t_L g725 ( .A(n_535), .Y(n_725) );
NOR2xp33_ASAP7_75t_L g536 ( .A(n_537), .B(n_538), .Y(n_536) );
NOR2xp33_ASAP7_75t_L g690 ( .A(n_538), .B(n_691), .Y(n_690) );
INVx4_ASAP7_75t_L g735 ( .A(n_538), .Y(n_735) );
NOR2xp33_ASAP7_75t_L g782 ( .A(n_538), .B(n_783), .Y(n_782) );
NOR2xp33_ASAP7_75t_L g890 ( .A(n_538), .B(n_891), .Y(n_890) );
INVx3_ASAP7_75t_L g538 ( .A(n_539), .Y(n_538) );
INVx4_ASAP7_75t_L g599 ( .A(n_539), .Y(n_599) );
INVx1_ASAP7_75t_L g543 ( .A(n_544), .Y(n_543) );
XNOR2xp5_ASAP7_75t_L g544 ( .A(n_545), .B(n_578), .Y(n_544) );
XNOR2x1_ASAP7_75t_L g545 ( .A(n_546), .B(n_577), .Y(n_545) );
OR2x2_ASAP7_75t_L g546 ( .A(n_547), .B(n_559), .Y(n_546) );
NAND4xp25_ASAP7_75t_SL g547 ( .A(n_548), .B(n_550), .C(n_553), .D(n_556), .Y(n_547) );
BUFx3_ASAP7_75t_L g708 ( .A(n_549), .Y(n_708) );
NAND3xp33_ASAP7_75t_L g559 ( .A(n_560), .B(n_569), .C(n_573), .Y(n_559) );
BUFx3_ASAP7_75t_L g561 ( .A(n_562), .Y(n_561) );
INVx1_ASAP7_75t_L g874 ( .A(n_562), .Y(n_874) );
OAI21xp5_ASAP7_75t_L g563 ( .A1(n_564), .A2(n_565), .B(n_566), .Y(n_563) );
INVx2_ASAP7_75t_L g597 ( .A(n_565), .Y(n_597) );
INVx2_ASAP7_75t_L g663 ( .A(n_565), .Y(n_663) );
INVx3_ASAP7_75t_L g676 ( .A(n_565), .Y(n_676) );
INVx2_ASAP7_75t_L g734 ( .A(n_565), .Y(n_734) );
INVx2_ASAP7_75t_L g567 ( .A(n_568), .Y(n_567) );
NOR2xp33_ASAP7_75t_L g921 ( .A(n_568), .B(n_922), .Y(n_921) );
INVx2_ASAP7_75t_L g570 ( .A(n_571), .Y(n_570) );
INVx3_ASAP7_75t_L g595 ( .A(n_571), .Y(n_595) );
INVx4_ASAP7_75t_L g594 ( .A(n_572), .Y(n_594) );
BUFx3_ASAP7_75t_L g869 ( .A(n_572), .Y(n_869) );
INVx4_ASAP7_75t_L g749 ( .A(n_574), .Y(n_749) );
BUFx3_ASAP7_75t_L g722 ( .A(n_575), .Y(n_722) );
INVx2_ASAP7_75t_L g575 ( .A(n_576), .Y(n_575) );
BUFx6f_ASAP7_75t_L g789 ( .A(n_576), .Y(n_789) );
INVx1_ASAP7_75t_L g579 ( .A(n_580), .Y(n_579) );
AOI22xp33_ASAP7_75t_SL g580 ( .A1(n_581), .A2(n_643), .B1(n_696), .B2(n_697), .Y(n_580) );
INVx2_ASAP7_75t_L g696 ( .A(n_581), .Y(n_696) );
AO22x2_ASAP7_75t_L g581 ( .A1(n_582), .A2(n_583), .B1(n_622), .B2(n_642), .Y(n_581) );
INVx2_ASAP7_75t_L g582 ( .A(n_583), .Y(n_582) );
INVx1_ASAP7_75t_L g584 ( .A(n_585), .Y(n_584) );
NAND3xp33_ASAP7_75t_L g585 ( .A(n_586), .B(n_600), .C(n_615), .Y(n_585) );
INVx1_ASAP7_75t_L g621 ( .A(n_586), .Y(n_621) );
AND3x2_ASAP7_75t_L g586 ( .A(n_587), .B(n_592), .C(n_596), .Y(n_586) );
INVxp67_ASAP7_75t_L g588 ( .A(n_589), .Y(n_588) );
INVx1_ASAP7_75t_L g589 ( .A(n_590), .Y(n_589) );
INVx2_ASAP7_75t_L g590 ( .A(n_591), .Y(n_590) );
BUFx6f_ASAP7_75t_L g760 ( .A(n_591), .Y(n_760) );
INVx1_ASAP7_75t_L g593 ( .A(n_594), .Y(n_593) );
INVx1_ASAP7_75t_L g598 ( .A(n_599), .Y(n_598) );
NOR2xp33_ASAP7_75t_L g629 ( .A(n_599), .B(n_630), .Y(n_629) );
NOR2xp33_ASAP7_75t_L g665 ( .A(n_599), .B(n_666), .Y(n_665) );
INVx4_ASAP7_75t_L g764 ( .A(n_599), .Y(n_764) );
NOR2xp33_ASAP7_75t_L g937 ( .A(n_599), .B(n_938), .Y(n_937) );
NOR2xp33_ASAP7_75t_L g1192 ( .A(n_599), .B(n_1193), .Y(n_1192) );
AND4x1_ASAP7_75t_L g600 ( .A(n_601), .B(n_603), .C(n_605), .D(n_612), .Y(n_600) );
BUFx4f_ASAP7_75t_L g606 ( .A(n_607), .Y(n_606) );
INVx1_ASAP7_75t_L g608 ( .A(n_609), .Y(n_608) );
INVx1_ASAP7_75t_L g609 ( .A(n_610), .Y(n_609) );
BUFx6f_ASAP7_75t_L g774 ( .A(n_610), .Y(n_774) );
INVx2_ASAP7_75t_L g610 ( .A(n_611), .Y(n_610) );
INVx2_ASAP7_75t_L g616 ( .A(n_617), .Y(n_616) );
INVx2_ASAP7_75t_L g618 ( .A(n_619), .Y(n_618) );
INVx1_ASAP7_75t_L g622 ( .A(n_623), .Y(n_622) );
HB1xp67_ASAP7_75t_L g642 ( .A(n_623), .Y(n_642) );
AO22x2_ASAP7_75t_L g645 ( .A1(n_623), .A2(n_646), .B1(n_647), .B2(n_668), .Y(n_645) );
INVx1_ASAP7_75t_L g668 ( .A(n_623), .Y(n_668) );
NAND3x1_ASAP7_75t_L g624 ( .A(n_625), .B(n_631), .C(n_636), .Y(n_624) );
HB1xp67_ASAP7_75t_L g786 ( .A(n_626), .Y(n_786) );
HB1xp67_ASAP7_75t_L g627 ( .A(n_628), .Y(n_627) );
AND2x2_ASAP7_75t_L g631 ( .A(n_632), .B(n_635), .Y(n_631) );
AND4x1_ASAP7_75t_L g636 ( .A(n_637), .B(n_638), .C(n_640), .D(n_641), .Y(n_636) );
INVx2_ASAP7_75t_L g846 ( .A(n_639), .Y(n_846) );
OAI21xp5_ASAP7_75t_L g643 ( .A1(n_644), .A2(n_669), .B(n_693), .Y(n_643) );
AOI22x1_ASAP7_75t_SL g697 ( .A1(n_644), .A2(n_670), .B1(n_694), .B2(n_698), .Y(n_697) );
INVx1_ASAP7_75t_L g644 ( .A(n_645), .Y(n_644) );
INVx2_ASAP7_75t_L g695 ( .A(n_645), .Y(n_695) );
INVx2_ASAP7_75t_L g646 ( .A(n_647), .Y(n_646) );
INVx2_ASAP7_75t_L g648 ( .A(n_649), .Y(n_648) );
NAND4xp75_ASAP7_75t_L g649 ( .A(n_650), .B(n_655), .C(n_659), .D(n_664), .Y(n_649) );
AND2x2_ASAP7_75t_L g650 ( .A(n_651), .B(n_652), .Y(n_650) );
AND2x2_ASAP7_75t_L g655 ( .A(n_656), .B(n_657), .Y(n_655) );
AND2x2_ASAP7_75t_L g659 ( .A(n_660), .B(n_662), .Y(n_659) );
INVx1_ASAP7_75t_L g669 ( .A(n_670), .Y(n_669) );
INVx1_ASAP7_75t_L g670 ( .A(n_671), .Y(n_670) );
HB1xp67_ASAP7_75t_L g694 ( .A(n_671), .Y(n_694) );
XOR2x2_ASAP7_75t_L g671 ( .A(n_672), .B(n_692), .Y(n_671) );
NOR4xp75_ASAP7_75t_L g672 ( .A(n_673), .B(n_677), .C(n_680), .D(n_685), .Y(n_672) );
NAND2xp5_ASAP7_75t_L g673 ( .A(n_674), .B(n_675), .Y(n_673) );
NAND2xp5_ASAP7_75t_L g677 ( .A(n_678), .B(n_679), .Y(n_677) );
NAND2xp5_ASAP7_75t_SL g680 ( .A(n_681), .B(n_684), .Y(n_680) );
OAI21x1_ASAP7_75t_SL g685 ( .A1(n_686), .A2(n_687), .B(n_689), .Y(n_685) );
INVx1_ASAP7_75t_L g687 ( .A(n_688), .Y(n_687) );
NAND2xp5_ASAP7_75t_L g693 ( .A(n_694), .B(n_695), .Y(n_693) );
INVx2_ASAP7_75t_L g698 ( .A(n_695), .Y(n_698) );
INVx1_ASAP7_75t_L g699 ( .A(n_700), .Y(n_699) );
XNOR2xp5_ASAP7_75t_L g700 ( .A(n_701), .B(n_861), .Y(n_700) );
AOI22xp5_ASAP7_75t_L g701 ( .A1(n_702), .A2(n_790), .B1(n_859), .B2(n_860), .Y(n_701) );
INVx1_ASAP7_75t_L g859 ( .A(n_702), .Y(n_859) );
XNOR2xp5_ASAP7_75t_L g702 ( .A(n_703), .B(n_766), .Y(n_702) );
OAI22xp5_ASAP7_75t_L g703 ( .A1(n_704), .A2(n_705), .B1(n_736), .B2(n_765), .Y(n_703) );
INVx3_ASAP7_75t_L g704 ( .A(n_705), .Y(n_704) );
NAND3xp33_ASAP7_75t_SL g706 ( .A(n_707), .B(n_710), .C(n_714), .Y(n_706) );
AND3x1_ASAP7_75t_L g710 ( .A(n_711), .B(n_712), .C(n_713), .Y(n_710) );
NOR3xp33_ASAP7_75t_L g714 ( .A(n_715), .B(n_723), .C(n_729), .Y(n_714) );
OAI22xp5_ASAP7_75t_L g715 ( .A1(n_716), .A2(n_717), .B1(n_720), .B2(n_721), .Y(n_715) );
INVx2_ASAP7_75t_L g717 ( .A(n_718), .Y(n_717) );
INVx2_ASAP7_75t_L g718 ( .A(n_719), .Y(n_718) );
INVxp67_ASAP7_75t_L g721 ( .A(n_722), .Y(n_721) );
OAI22xp5_ASAP7_75t_L g723 ( .A1(n_724), .A2(n_725), .B1(n_726), .B2(n_727), .Y(n_723) );
INVx1_ASAP7_75t_L g727 ( .A(n_728), .Y(n_727) );
OAI21xp33_ASAP7_75t_L g729 ( .A1(n_730), .A2(n_731), .B(n_733), .Y(n_729) );
INVx1_ASAP7_75t_L g731 ( .A(n_732), .Y(n_731) );
INVx1_ASAP7_75t_L g736 ( .A(n_737), .Y(n_736) );
INVx1_ASAP7_75t_L g737 ( .A(n_738), .Y(n_737) );
INVx1_ASAP7_75t_L g765 ( .A(n_738), .Y(n_765) );
INVx2_ASAP7_75t_L g738 ( .A(n_739), .Y(n_738) );
NAND4xp75_ASAP7_75t_L g740 ( .A(n_741), .B(n_751), .C(n_754), .D(n_758), .Y(n_740) );
NOR2xp67_ASAP7_75t_L g741 ( .A(n_742), .B(n_747), .Y(n_741) );
OAI22xp5_ASAP7_75t_L g742 ( .A1(n_743), .A2(n_744), .B1(n_745), .B2(n_746), .Y(n_742) );
OAI21xp5_ASAP7_75t_L g747 ( .A1(n_748), .A2(n_749), .B(n_750), .Y(n_747) );
AND2x2_ASAP7_75t_L g751 ( .A(n_752), .B(n_753), .Y(n_751) );
AND2x2_ASAP7_75t_L g754 ( .A(n_755), .B(n_756), .Y(n_754) );
INVx2_ASAP7_75t_L g759 ( .A(n_760), .Y(n_759) );
INVx2_ASAP7_75t_L g808 ( .A(n_760), .Y(n_808) );
NOR2xp33_ASAP7_75t_L g761 ( .A(n_762), .B(n_763), .Y(n_761) );
INVx2_ASAP7_75t_L g763 ( .A(n_764), .Y(n_763) );
INVx1_ASAP7_75t_SL g766 ( .A(n_767), .Y(n_766) );
INVx1_ASAP7_75t_L g767 ( .A(n_768), .Y(n_767) );
INVx2_ASAP7_75t_SL g768 ( .A(n_769), .Y(n_768) );
XNOR2x1_ASAP7_75t_L g769 ( .A(n_770), .B(n_771), .Y(n_769) );
NOR2x1_ASAP7_75t_L g771 ( .A(n_772), .B(n_778), .Y(n_771) );
NAND4xp25_ASAP7_75t_L g772 ( .A(n_773), .B(n_775), .C(n_776), .D(n_777), .Y(n_772) );
NAND3xp33_ASAP7_75t_L g778 ( .A(n_779), .B(n_785), .C(n_787), .Y(n_778) );
INVx1_ASAP7_75t_L g779 ( .A(n_780), .Y(n_779) );
NAND2xp5_ASAP7_75t_L g780 ( .A(n_781), .B(n_784), .Y(n_780) );
INVx2_ASAP7_75t_L g788 ( .A(n_789), .Y(n_788) );
INVx2_ASAP7_75t_L g871 ( .A(n_789), .Y(n_871) );
INVx2_ASAP7_75t_L g790 ( .A(n_791), .Y(n_790) );
BUFx3_ASAP7_75t_L g860 ( .A(n_791), .Y(n_860) );
OAI22x1_ASAP7_75t_L g791 ( .A1(n_792), .A2(n_832), .B1(n_857), .B2(n_858), .Y(n_791) );
INVx2_ASAP7_75t_L g857 ( .A(n_792), .Y(n_857) );
OA22x2_ASAP7_75t_L g792 ( .A1(n_793), .A2(n_794), .B1(n_815), .B2(n_831), .Y(n_792) );
INVx1_ASAP7_75t_L g793 ( .A(n_794), .Y(n_793) );
NAND4xp75_ASAP7_75t_L g795 ( .A(n_796), .B(n_801), .C(n_804), .D(n_807), .Y(n_795) );
AND2x2_ASAP7_75t_L g796 ( .A(n_797), .B(n_799), .Y(n_796) );
AND2x2_ASAP7_75t_L g801 ( .A(n_802), .B(n_803), .Y(n_801) );
AND2x2_ASAP7_75t_L g804 ( .A(n_805), .B(n_806), .Y(n_804) );
OAI21xp5_ASAP7_75t_L g809 ( .A1(n_810), .A2(n_811), .B(n_813), .Y(n_809) );
OAI22xp5_ASAP7_75t_L g893 ( .A1(n_811), .A2(n_894), .B1(n_896), .B2(n_898), .Y(n_893) );
INVx4_ASAP7_75t_L g811 ( .A(n_812), .Y(n_811) );
INVx2_ASAP7_75t_L g831 ( .A(n_815), .Y(n_831) );
NOR2x1_ASAP7_75t_L g816 ( .A(n_817), .B(n_822), .Y(n_816) );
NAND4xp25_ASAP7_75t_L g817 ( .A(n_818), .B(n_819), .C(n_820), .D(n_821), .Y(n_817) );
NAND4xp25_ASAP7_75t_SL g822 ( .A(n_823), .B(n_826), .C(n_827), .D(n_829), .Y(n_822) );
INVx1_ASAP7_75t_L g832 ( .A(n_833), .Y(n_832) );
INVx2_ASAP7_75t_L g833 ( .A(n_834), .Y(n_833) );
INVx1_ASAP7_75t_L g858 ( .A(n_834), .Y(n_858) );
NAND4xp75_ASAP7_75t_L g835 ( .A(n_836), .B(n_840), .C(n_843), .D(n_853), .Y(n_835) );
AND2x2_ASAP7_75t_L g836 ( .A(n_837), .B(n_838), .Y(n_836) );
AND2x2_ASAP7_75t_L g840 ( .A(n_841), .B(n_842), .Y(n_840) );
NOR2xp33_ASAP7_75t_L g843 ( .A(n_844), .B(n_848), .Y(n_843) );
OAI21xp33_ASAP7_75t_L g844 ( .A1(n_845), .A2(n_846), .B(n_847), .Y(n_844) );
OAI22xp5_ASAP7_75t_L g848 ( .A1(n_849), .A2(n_850), .B1(n_851), .B2(n_852), .Y(n_848) );
OAI22xp33_ASAP7_75t_L g861 ( .A1(n_862), .A2(n_863), .B1(n_909), .B2(n_958), .Y(n_861) );
INVx1_ASAP7_75t_L g862 ( .A(n_863), .Y(n_862) );
OA22x2_ASAP7_75t_L g863 ( .A1(n_864), .A2(n_885), .B1(n_907), .B2(n_908), .Y(n_863) );
INVx1_ASAP7_75t_L g907 ( .A(n_864), .Y(n_907) );
XOR2x2_ASAP7_75t_L g864 ( .A(n_865), .B(n_884), .Y(n_864) );
NOR2x1_ASAP7_75t_L g865 ( .A(n_866), .B(n_876), .Y(n_865) );
NAND4xp25_ASAP7_75t_L g866 ( .A(n_867), .B(n_870), .C(n_872), .D(n_875), .Y(n_866) );
INVx2_ASAP7_75t_L g873 ( .A(n_874), .Y(n_873) );
NAND4xp25_ASAP7_75t_L g876 ( .A(n_877), .B(n_879), .C(n_882), .D(n_883), .Y(n_876) );
INVx1_ASAP7_75t_L g908 ( .A(n_885), .Y(n_908) );
INVx1_ASAP7_75t_L g885 ( .A(n_886), .Y(n_885) );
INVx1_ASAP7_75t_L g906 ( .A(n_887), .Y(n_906) );
NOR2x1_ASAP7_75t_L g887 ( .A(n_888), .B(n_900), .Y(n_887) );
NAND3xp33_ASAP7_75t_L g888 ( .A(n_889), .B(n_892), .C(n_899), .Y(n_888) );
CKINVDCx16_ASAP7_75t_R g894 ( .A(n_895), .Y(n_894) );
CKINVDCx9p33_ASAP7_75t_R g896 ( .A(n_897), .Y(n_896) );
NAND4xp25_ASAP7_75t_L g900 ( .A(n_901), .B(n_902), .C(n_903), .D(n_904), .Y(n_900) );
INVx1_ASAP7_75t_L g958 ( .A(n_909), .Y(n_958) );
INVx1_ASAP7_75t_L g909 ( .A(n_910), .Y(n_909) );
XOR2x2_ASAP7_75t_L g910 ( .A(n_911), .B(n_928), .Y(n_910) );
HB1xp67_ASAP7_75t_L g911 ( .A(n_912), .Y(n_911) );
XNOR2xp5_ASAP7_75t_L g912 ( .A(n_913), .B(n_914), .Y(n_912) );
NOR2xp67_ASAP7_75t_L g914 ( .A(n_915), .B(n_923), .Y(n_914) );
NAND4xp25_ASAP7_75t_L g915 ( .A(n_916), .B(n_917), .C(n_919), .D(n_920), .Y(n_915) );
NAND4xp25_ASAP7_75t_SL g923 ( .A(n_924), .B(n_925), .C(n_926), .D(n_927), .Y(n_923) );
OA22x2_ASAP7_75t_L g928 ( .A1(n_929), .A2(n_930), .B1(n_944), .B2(n_957), .Y(n_928) );
INVx1_ASAP7_75t_L g929 ( .A(n_930), .Y(n_929) );
OR2x2_ASAP7_75t_L g931 ( .A(n_932), .B(n_939), .Y(n_931) );
NAND4xp25_ASAP7_75t_L g932 ( .A(n_933), .B(n_934), .C(n_935), .D(n_936), .Y(n_932) );
NAND4xp25_ASAP7_75t_L g939 ( .A(n_940), .B(n_941), .C(n_942), .D(n_943), .Y(n_939) );
XNOR2xp5_ASAP7_75t_L g944 ( .A(n_945), .B(n_946), .Y(n_944) );
XOR2xp5_ASAP7_75t_L g957 ( .A(n_945), .B(n_946), .Y(n_957) );
OR2x2_ASAP7_75t_L g946 ( .A(n_947), .B(n_952), .Y(n_946) );
NAND4xp25_ASAP7_75t_L g947 ( .A(n_948), .B(n_949), .C(n_950), .D(n_951), .Y(n_947) );
NAND4xp25_ASAP7_75t_L g952 ( .A(n_953), .B(n_954), .C(n_955), .D(n_956), .Y(n_952) );
OAI221xp5_ASAP7_75t_L g959 ( .A1(n_960), .A2(n_1180), .B1(n_1182), .B2(n_1199), .C(n_1204), .Y(n_959) );
AOI211xp5_ASAP7_75t_L g960 ( .A1(n_961), .A2(n_1091), .B(n_1098), .C(n_1147), .Y(n_960) );
NAND5xp2_ASAP7_75t_L g961 ( .A(n_962), .B(n_1036), .C(n_1061), .D(n_1073), .E(n_1078), .Y(n_961) );
AOI211xp5_ASAP7_75t_SL g962 ( .A1(n_963), .A2(n_995), .B(n_999), .C(n_1028), .Y(n_962) );
AND2x2_ASAP7_75t_L g963 ( .A(n_964), .B(n_978), .Y(n_963) );
NOR2xp33_ASAP7_75t_L g1030 ( .A(n_964), .B(n_1027), .Y(n_1030) );
NAND2xp5_ASAP7_75t_L g1077 ( .A(n_964), .B(n_1035), .Y(n_1077) );
AND2x2_ASAP7_75t_L g1079 ( .A(n_964), .B(n_1080), .Y(n_1079) );
NOR2xp33_ASAP7_75t_L g1131 ( .A(n_964), .B(n_1132), .Y(n_1131) );
NOR2xp33_ASAP7_75t_L g1164 ( .A(n_964), .B(n_1165), .Y(n_1164) );
INVx2_ASAP7_75t_L g964 ( .A(n_965), .Y(n_964) );
INVx3_ASAP7_75t_L g1022 ( .A(n_965), .Y(n_1022) );
AND2x2_ASAP7_75t_L g1060 ( .A(n_965), .B(n_1043), .Y(n_1060) );
NAND2xp5_ASAP7_75t_L g1068 ( .A(n_965), .B(n_1001), .Y(n_1068) );
INVx2_ASAP7_75t_L g1101 ( .A(n_965), .Y(n_1101) );
NAND2xp5_ASAP7_75t_L g1110 ( .A(n_965), .B(n_1072), .Y(n_1110) );
NOR3xp33_ASAP7_75t_L g1157 ( .A(n_965), .B(n_1025), .C(n_1093), .Y(n_1157) );
NOR2xp33_ASAP7_75t_L g1179 ( .A(n_965), .B(n_1083), .Y(n_1179) );
AND2x2_ASAP7_75t_L g965 ( .A(n_966), .B(n_973), .Y(n_965) );
AND2x2_ASAP7_75t_L g967 ( .A(n_968), .B(n_970), .Y(n_967) );
AND2x4_ASAP7_75t_L g974 ( .A(n_968), .B(n_975), .Y(n_974) );
AND2x2_ASAP7_75t_L g991 ( .A(n_968), .B(n_970), .Y(n_991) );
AND2x4_ASAP7_75t_L g994 ( .A(n_968), .B(n_970), .Y(n_994) );
AND2x2_ASAP7_75t_L g971 ( .A(n_970), .B(n_972), .Y(n_971) );
AND2x2_ASAP7_75t_L g983 ( .A(n_970), .B(n_972), .Y(n_983) );
AND2x4_ASAP7_75t_L g1007 ( .A(n_970), .B(n_972), .Y(n_1007) );
AND2x4_ASAP7_75t_L g977 ( .A(n_972), .B(n_975), .Y(n_977) );
AND2x4_ASAP7_75t_L g981 ( .A(n_972), .B(n_975), .Y(n_981) );
INVx3_ASAP7_75t_L g1096 ( .A(n_974), .Y(n_1096) );
INVx2_ASAP7_75t_SL g1005 ( .A(n_977), .Y(n_1005) );
NAND2xp5_ASAP7_75t_L g1115 ( .A(n_978), .B(n_1033), .Y(n_1115) );
AND2x2_ASAP7_75t_L g978 ( .A(n_979), .B(n_984), .Y(n_978) );
AND2x2_ASAP7_75t_L g1020 ( .A(n_979), .B(n_1021), .Y(n_1020) );
AND2x2_ASAP7_75t_L g1035 ( .A(n_979), .B(n_1024), .Y(n_1035) );
AND2x2_ASAP7_75t_L g1037 ( .A(n_979), .B(n_1038), .Y(n_1037) );
CKINVDCx6p67_ASAP7_75t_R g1043 ( .A(n_979), .Y(n_1043) );
AOI32xp33_ASAP7_75t_L g1078 ( .A1(n_979), .A2(n_1079), .A3(n_1081), .B1(n_1084), .B2(n_1088), .Y(n_1078) );
NOR2xp33_ASAP7_75t_L g1090 ( .A(n_979), .B(n_985), .Y(n_1090) );
AND2x2_ASAP7_75t_L g1102 ( .A(n_979), .B(n_1018), .Y(n_1102) );
NAND2xp5_ASAP7_75t_L g1120 ( .A(n_979), .B(n_1025), .Y(n_1120) );
AND2x2_ASAP7_75t_L g1140 ( .A(n_979), .B(n_986), .Y(n_1140) );
AND2x2_ASAP7_75t_L g979 ( .A(n_980), .B(n_982), .Y(n_979) );
NAND2xp5_ASAP7_75t_L g1064 ( .A(n_984), .B(n_1020), .Y(n_1064) );
INVx1_ASAP7_75t_L g1083 ( .A(n_984), .Y(n_1083) );
AND2x2_ASAP7_75t_L g1106 ( .A(n_984), .B(n_1043), .Y(n_1106) );
AND2x2_ASAP7_75t_L g1114 ( .A(n_984), .B(n_1060), .Y(n_1114) );
AND2x2_ASAP7_75t_L g984 ( .A(n_985), .B(n_992), .Y(n_984) );
OAI221xp5_ASAP7_75t_L g1152 ( .A1(n_985), .A2(n_1033), .B1(n_1128), .B2(n_1153), .C(n_1154), .Y(n_1152) );
NAND2xp5_ASAP7_75t_L g1165 ( .A(n_985), .B(n_1043), .Y(n_1165) );
INVx1_ASAP7_75t_L g985 ( .A(n_986), .Y(n_985) );
OR2x2_ASAP7_75t_L g1019 ( .A(n_986), .B(n_992), .Y(n_1019) );
AND2x2_ASAP7_75t_L g1024 ( .A(n_986), .B(n_1025), .Y(n_1024) );
AND2x2_ASAP7_75t_L g1039 ( .A(n_986), .B(n_992), .Y(n_1039) );
AND2x2_ASAP7_75t_L g986 ( .A(n_987), .B(n_990), .Y(n_986) );
INVx1_ASAP7_75t_L g1025 ( .A(n_992), .Y(n_1025) );
NAND2xp5_ASAP7_75t_L g1049 ( .A(n_992), .B(n_1020), .Y(n_1049) );
AND2x2_ASAP7_75t_L g1137 ( .A(n_992), .B(n_1043), .Y(n_1137) );
BUFx2_ASAP7_75t_L g1181 ( .A(n_994), .Y(n_1181) );
INVxp67_ASAP7_75t_L g1008 ( .A(n_995), .Y(n_1008) );
OR2x2_ASAP7_75t_L g1048 ( .A(n_995), .B(n_1014), .Y(n_1048) );
OR2x2_ASAP7_75t_L g1053 ( .A(n_995), .B(n_1013), .Y(n_1053) );
AND2x2_ASAP7_75t_L g1072 ( .A(n_995), .B(n_1014), .Y(n_1072) );
INVx2_ASAP7_75t_L g1076 ( .A(n_995), .Y(n_1076) );
AND2x2_ASAP7_75t_L g1087 ( .A(n_995), .B(n_1001), .Y(n_1087) );
INVx2_ASAP7_75t_L g995 ( .A(n_996), .Y(n_995) );
OR2x2_ASAP7_75t_L g1027 ( .A(n_996), .B(n_1014), .Y(n_1027) );
AND2x2_ASAP7_75t_L g1044 ( .A(n_996), .B(n_1002), .Y(n_1044) );
NAND2xp5_ASAP7_75t_L g996 ( .A(n_997), .B(n_998), .Y(n_996) );
OAI21xp33_ASAP7_75t_L g999 ( .A1(n_1000), .A2(n_1009), .B(n_1023), .Y(n_999) );
INVx1_ASAP7_75t_L g1135 ( .A(n_1000), .Y(n_1135) );
AOI21xp33_ASAP7_75t_SL g1167 ( .A1(n_1000), .A2(n_1150), .B(n_1168), .Y(n_1167) );
OR2x2_ASAP7_75t_L g1000 ( .A(n_1001), .B(n_1008), .Y(n_1000) );
NOR2xp33_ASAP7_75t_L g1026 ( .A(n_1001), .B(n_1027), .Y(n_1026) );
AND2x2_ASAP7_75t_L g1032 ( .A(n_1001), .B(n_1033), .Y(n_1032) );
NAND2xp5_ASAP7_75t_L g1046 ( .A(n_1001), .B(n_1047), .Y(n_1046) );
NAND2xp5_ASAP7_75t_L g1075 ( .A(n_1001), .B(n_1076), .Y(n_1075) );
AOI32xp33_ASAP7_75t_L g1125 ( .A1(n_1001), .A2(n_1079), .A3(n_1126), .B1(n_1127), .B2(n_1129), .Y(n_1125) );
INVx2_ASAP7_75t_L g1151 ( .A(n_1001), .Y(n_1151) );
INVx4_ASAP7_75t_L g1001 ( .A(n_1002), .Y(n_1001) );
NAND2xp5_ASAP7_75t_L g1066 ( .A(n_1002), .B(n_1011), .Y(n_1066) );
NOR2xp33_ASAP7_75t_L g1146 ( .A(n_1002), .B(n_1093), .Y(n_1146) );
AND2x2_ASAP7_75t_L g1158 ( .A(n_1002), .B(n_1080), .Y(n_1158) );
NOR2xp33_ASAP7_75t_L g1160 ( .A(n_1002), .B(n_1053), .Y(n_1160) );
AND2x2_ASAP7_75t_L g1166 ( .A(n_1002), .B(n_1033), .Y(n_1166) );
AND2x2_ASAP7_75t_L g1002 ( .A(n_1003), .B(n_1006), .Y(n_1002) );
INVx2_ASAP7_75t_L g1004 ( .A(n_1005), .Y(n_1004) );
INVx1_ASAP7_75t_L g1129 ( .A(n_1008), .Y(n_1129) );
NAND2xp5_ASAP7_75t_L g1009 ( .A(n_1010), .B(n_1017), .Y(n_1009) );
NOR2xp33_ASAP7_75t_L g1040 ( .A(n_1010), .B(n_1041), .Y(n_1040) );
INVx2_ASAP7_75t_L g1010 ( .A(n_1011), .Y(n_1010) );
INVx1_ASAP7_75t_L g1011 ( .A(n_1012), .Y(n_1011) );
INVx1_ASAP7_75t_L g1058 ( .A(n_1012), .Y(n_1058) );
INVx1_ASAP7_75t_L g1012 ( .A(n_1013), .Y(n_1012) );
INVx2_ASAP7_75t_L g1033 ( .A(n_1013), .Y(n_1033) );
INVx4_ASAP7_75t_L g1013 ( .A(n_1014), .Y(n_1013) );
NAND2xp5_ASAP7_75t_L g1170 ( .A(n_1014), .B(n_1101), .Y(n_1170) );
AND2x2_ASAP7_75t_L g1014 ( .A(n_1015), .B(n_1016), .Y(n_1014) );
NAND2xp5_ASAP7_75t_L g1123 ( .A(n_1017), .B(n_1124), .Y(n_1123) );
AND2x2_ASAP7_75t_L g1017 ( .A(n_1018), .B(n_1020), .Y(n_1017) );
AND2x2_ASAP7_75t_L g1042 ( .A(n_1018), .B(n_1043), .Y(n_1042) );
AND2x2_ASAP7_75t_L g1059 ( .A(n_1018), .B(n_1060), .Y(n_1059) );
INVx1_ASAP7_75t_L g1018 ( .A(n_1019), .Y(n_1018) );
NOR2x1_ASAP7_75t_L g1070 ( .A(n_1019), .B(n_1021), .Y(n_1070) );
NAND2xp5_ASAP7_75t_L g1128 ( .A(n_1020), .B(n_1039), .Y(n_1128) );
NOR2x1_ASAP7_75t_L g1062 ( .A(n_1021), .B(n_1052), .Y(n_1062) );
A2O1A1Ixp33_ASAP7_75t_L g1104 ( .A1(n_1021), .A2(n_1027), .B(n_1105), .C(n_1107), .Y(n_1104) );
AOI221xp5_ASAP7_75t_L g1111 ( .A1(n_1021), .A2(n_1087), .B1(n_1112), .B2(n_1117), .C(n_1122), .Y(n_1111) );
NAND2xp5_ASAP7_75t_L g1153 ( .A(n_1021), .B(n_1047), .Y(n_1153) );
INVx3_ASAP7_75t_L g1021 ( .A(n_1022), .Y(n_1021) );
AND2x2_ASAP7_75t_L g1038 ( .A(n_1022), .B(n_1039), .Y(n_1038) );
NAND2xp5_ASAP7_75t_L g1089 ( .A(n_1022), .B(n_1090), .Y(n_1089) );
AND2x2_ASAP7_75t_L g1141 ( .A(n_1022), .B(n_1047), .Y(n_1141) );
NAND2xp5_ASAP7_75t_L g1023 ( .A(n_1024), .B(n_1026), .Y(n_1023) );
NAND2xp5_ASAP7_75t_L g1052 ( .A(n_1024), .B(n_1043), .Y(n_1052) );
INVx1_ASAP7_75t_L g1082 ( .A(n_1024), .Y(n_1082) );
O2A1O1Ixp33_ASAP7_75t_L g1067 ( .A1(n_1025), .A2(n_1068), .B(n_1069), .C(n_1071), .Y(n_1067) );
NAND2xp5_ASAP7_75t_L g1109 ( .A(n_1025), .B(n_1043), .Y(n_1109) );
INVx1_ASAP7_75t_L g1155 ( .A(n_1027), .Y(n_1155) );
AOI21xp33_ASAP7_75t_SL g1176 ( .A1(n_1027), .A2(n_1177), .B(n_1178), .Y(n_1176) );
AOI21xp33_ASAP7_75t_L g1028 ( .A1(n_1029), .A2(n_1031), .B(n_1034), .Y(n_1028) );
INVx1_ASAP7_75t_L g1029 ( .A(n_1030), .Y(n_1029) );
INVx1_ASAP7_75t_L g1031 ( .A(n_1032), .Y(n_1031) );
AOI22xp5_ASAP7_75t_L g1159 ( .A1(n_1032), .A2(n_1051), .B1(n_1062), .B2(n_1160), .Y(n_1159) );
AOI32xp33_ASAP7_75t_L g1142 ( .A1(n_1033), .A2(n_1064), .A3(n_1105), .B1(n_1143), .B2(n_1144), .Y(n_1142) );
NAND2xp5_ASAP7_75t_L g1163 ( .A(n_1033), .B(n_1164), .Y(n_1163) );
NAND2xp5_ASAP7_75t_L g1119 ( .A(n_1034), .B(n_1105), .Y(n_1119) );
INVx1_ASAP7_75t_L g1034 ( .A(n_1035), .Y(n_1034) );
O2A1O1Ixp33_ASAP7_75t_L g1036 ( .A1(n_1037), .A2(n_1040), .B(n_1044), .C(n_1045), .Y(n_1036) );
INVx1_ASAP7_75t_L g1132 ( .A(n_1039), .Y(n_1132) );
NAND2xp5_ASAP7_75t_L g1175 ( .A(n_1039), .B(n_1060), .Y(n_1175) );
INVx1_ASAP7_75t_L g1041 ( .A(n_1042), .Y(n_1041) );
NAND2xp5_ASAP7_75t_L g1069 ( .A(n_1043), .B(n_1070), .Y(n_1069) );
A2O1A1Ixp33_ASAP7_75t_SL g1130 ( .A1(n_1044), .A2(n_1092), .B(n_1131), .C(n_1133), .Y(n_1130) );
OAI221xp5_ASAP7_75t_L g1045 ( .A1(n_1046), .A2(n_1049), .B1(n_1050), .B2(n_1053), .C(n_1054), .Y(n_1045) );
INVx1_ASAP7_75t_L g1047 ( .A(n_1048), .Y(n_1047) );
INVx2_ASAP7_75t_L g1050 ( .A(n_1051), .Y(n_1050) );
NAND2xp5_ASAP7_75t_L g1107 ( .A(n_1051), .B(n_1072), .Y(n_1107) );
INVx1_ASAP7_75t_L g1051 ( .A(n_1052), .Y(n_1051) );
INVx1_ASAP7_75t_L g1080 ( .A(n_1053), .Y(n_1080) );
OAI22xp5_ASAP7_75t_L g1117 ( .A1(n_1053), .A2(n_1118), .B1(n_1120), .B2(n_1121), .Y(n_1117) );
NAND2xp5_ASAP7_75t_L g1054 ( .A(n_1055), .B(n_1059), .Y(n_1054) );
HB1xp67_ASAP7_75t_L g1055 ( .A(n_1056), .Y(n_1055) );
NAND2xp5_ASAP7_75t_L g1113 ( .A(n_1056), .B(n_1114), .Y(n_1113) );
NOR2xp33_ASAP7_75t_L g1127 ( .A(n_1056), .B(n_1128), .Y(n_1127) );
HB1xp67_ASAP7_75t_L g1173 ( .A(n_1056), .Y(n_1173) );
INVx1_ASAP7_75t_L g1056 ( .A(n_1057), .Y(n_1056) );
INVx1_ASAP7_75t_L g1086 ( .A(n_1057), .Y(n_1086) );
INVx1_ASAP7_75t_L g1057 ( .A(n_1058), .Y(n_1057) );
HB1xp67_ASAP7_75t_L g1124 ( .A(n_1058), .Y(n_1124) );
INVx1_ASAP7_75t_L g1177 ( .A(n_1059), .Y(n_1177) );
O2A1O1Ixp33_ASAP7_75t_L g1061 ( .A1(n_1062), .A2(n_1063), .B(n_1065), .C(n_1067), .Y(n_1061) );
INVx1_ASAP7_75t_L g1063 ( .A(n_1064), .Y(n_1063) );
INVx1_ASAP7_75t_L g1065 ( .A(n_1066), .Y(n_1065) );
INVx1_ASAP7_75t_L g1143 ( .A(n_1070), .Y(n_1143) );
INVx1_ASAP7_75t_L g1071 ( .A(n_1072), .Y(n_1071) );
INVx1_ASAP7_75t_L g1073 ( .A(n_1074), .Y(n_1073) );
NOR2xp33_ASAP7_75t_L g1074 ( .A(n_1075), .B(n_1077), .Y(n_1074) );
INVx3_ASAP7_75t_SL g1103 ( .A(n_1076), .Y(n_1103) );
NAND2xp5_ASAP7_75t_L g1121 ( .A(n_1076), .B(n_1092), .Y(n_1121) );
AND2x2_ASAP7_75t_L g1081 ( .A(n_1082), .B(n_1083), .Y(n_1081) );
INVx1_ASAP7_75t_L g1084 ( .A(n_1085), .Y(n_1084) );
NAND2xp5_ASAP7_75t_L g1085 ( .A(n_1086), .B(n_1087), .Y(n_1085) );
HB1xp67_ASAP7_75t_L g1145 ( .A(n_1086), .Y(n_1145) );
INVxp33_ASAP7_75t_SL g1088 ( .A(n_1089), .Y(n_1088) );
OAI211xp5_ASAP7_75t_L g1098 ( .A1(n_1091), .A2(n_1099), .B(n_1111), .C(n_1138), .Y(n_1098) );
INVx2_ASAP7_75t_L g1091 ( .A(n_1092), .Y(n_1091) );
NAND2xp5_ASAP7_75t_L g1150 ( .A(n_1092), .B(n_1151), .Y(n_1150) );
CKINVDCx5p33_ASAP7_75t_R g1092 ( .A(n_1093), .Y(n_1092) );
AND2x2_ASAP7_75t_L g1093 ( .A(n_1094), .B(n_1097), .Y(n_1093) );
INVx1_ASAP7_75t_L g1095 ( .A(n_1096), .Y(n_1095) );
AOI211xp5_ASAP7_75t_L g1099 ( .A1(n_1100), .A2(n_1103), .B(n_1104), .C(n_1108), .Y(n_1099) );
INVx1_ASAP7_75t_L g1116 ( .A(n_1100), .Y(n_1116) );
AOI22xp33_ASAP7_75t_L g1148 ( .A1(n_1100), .A2(n_1149), .B1(n_1152), .B2(n_1155), .Y(n_1148) );
OAI31xp33_ASAP7_75t_L g1156 ( .A1(n_1100), .A2(n_1106), .A3(n_1157), .B(n_1158), .Y(n_1156) );
AND2x2_ASAP7_75t_L g1100 ( .A(n_1101), .B(n_1102), .Y(n_1100) );
AND2x2_ASAP7_75t_L g1136 ( .A(n_1101), .B(n_1137), .Y(n_1136) );
INVx1_ASAP7_75t_L g1154 ( .A(n_1102), .Y(n_1154) );
OAI211xp5_ASAP7_75t_SL g1122 ( .A1(n_1103), .A2(n_1123), .B(n_1125), .C(n_1130), .Y(n_1122) );
INVx1_ASAP7_75t_L g1105 ( .A(n_1106), .Y(n_1105) );
NOR2xp33_ASAP7_75t_L g1108 ( .A(n_1109), .B(n_1110), .Y(n_1108) );
INVx1_ASAP7_75t_L g1126 ( .A(n_1109), .Y(n_1126) );
NAND3xp33_ASAP7_75t_L g1112 ( .A(n_1113), .B(n_1115), .C(n_1116), .Y(n_1112) );
AOI221xp5_ASAP7_75t_L g1161 ( .A1(n_1114), .A2(n_1149), .B1(n_1162), .B2(n_1166), .C(n_1167), .Y(n_1161) );
INVx1_ASAP7_75t_L g1118 ( .A(n_1119), .Y(n_1118) );
INVxp67_ASAP7_75t_SL g1133 ( .A(n_1134), .Y(n_1133) );
NAND2xp5_ASAP7_75t_L g1134 ( .A(n_1135), .B(n_1136), .Y(n_1134) );
A2O1A1Ixp33_ASAP7_75t_SL g1138 ( .A1(n_1139), .A2(n_1141), .B(n_1142), .C(n_1146), .Y(n_1138) );
INVx1_ASAP7_75t_L g1139 ( .A(n_1140), .Y(n_1139) );
NAND2xp5_ASAP7_75t_L g1168 ( .A(n_1140), .B(n_1169), .Y(n_1168) );
HB1xp67_ASAP7_75t_L g1144 ( .A(n_1145), .Y(n_1144) );
NAND5xp2_ASAP7_75t_L g1147 ( .A(n_1148), .B(n_1156), .C(n_1159), .D(n_1161), .E(n_1171), .Y(n_1147) );
INVx1_ASAP7_75t_L g1149 ( .A(n_1150), .Y(n_1149) );
A2O1A1Ixp33_ASAP7_75t_L g1171 ( .A1(n_1151), .A2(n_1172), .B(n_1174), .C(n_1176), .Y(n_1171) );
INVxp67_ASAP7_75t_SL g1162 ( .A(n_1163), .Y(n_1162) );
INVx1_ASAP7_75t_L g1169 ( .A(n_1170), .Y(n_1169) );
HB1xp67_ASAP7_75t_L g1172 ( .A(n_1173), .Y(n_1172) );
INVx1_ASAP7_75t_L g1174 ( .A(n_1175), .Y(n_1174) );
INVx1_ASAP7_75t_L g1178 ( .A(n_1179), .Y(n_1178) );
CKINVDCx5p33_ASAP7_75t_R g1180 ( .A(n_1181), .Y(n_1180) );
INVx3_ASAP7_75t_L g1182 ( .A(n_1183), .Y(n_1182) );
BUFx3_ASAP7_75t_L g1183 ( .A(n_1184), .Y(n_1183) );
XNOR2x1_ASAP7_75t_L g1184 ( .A(n_1185), .B(n_1186), .Y(n_1184) );
INVx1_ASAP7_75t_L g1207 ( .A(n_1186), .Y(n_1207) );
OR2x2_ASAP7_75t_L g1186 ( .A(n_1187), .B(n_1194), .Y(n_1186) );
NAND4xp25_ASAP7_75t_L g1187 ( .A(n_1188), .B(n_1189), .C(n_1190), .D(n_1191), .Y(n_1187) );
NAND4xp25_ASAP7_75t_L g1194 ( .A(n_1195), .B(n_1196), .C(n_1197), .D(n_1198), .Y(n_1194) );
INVx1_ASAP7_75t_L g1199 ( .A(n_1200), .Y(n_1199) );
HB1xp67_ASAP7_75t_L g1200 ( .A(n_1201), .Y(n_1200) );
HB1xp67_ASAP7_75t_L g1208 ( .A(n_1209), .Y(n_1208) );
BUFx3_ASAP7_75t_L g1210 ( .A(n_1211), .Y(n_1210) );
CKINVDCx5p33_ASAP7_75t_R g1212 ( .A(n_1213), .Y(n_1212) );
endmodule