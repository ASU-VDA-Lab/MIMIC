module fake_jpeg_12339_n_130 (n_13, n_21, n_33, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_19, n_18, n_20, n_35, n_4, n_34, n_30, n_39, n_16, n_3, n_0, n_24, n_28, n_38, n_26, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_12, n_32, n_8, n_15, n_7, n_130);

input n_13;
input n_21;
input n_33;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_35;
input n_4;
input n_34;
input n_30;
input n_39;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_130;

wire n_117;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_73;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_42;
wire n_49;
wire n_76;
wire n_127;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_103;
wire n_50;
wire n_124;
wire n_57;
wire n_119;
wire n_69;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_106;
wire n_111;
wire n_44;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_121;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_56;
wire n_79;
wire n_67;
wire n_53;
wire n_54;
wire n_91;
wire n_93;
wire n_101;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_97;
wire n_62;
wire n_120;
wire n_43;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_96;

BUFx3_ASAP7_75t_L g40 ( 
.A(n_28),
.Y(n_40)
);

BUFx16f_ASAP7_75t_L g41 ( 
.A(n_30),
.Y(n_41)
);

BUFx3_ASAP7_75t_L g42 ( 
.A(n_3),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_8),
.Y(n_43)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_33),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_20),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_3),
.Y(n_46)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_34),
.Y(n_47)
);

INVx4_ASAP7_75t_L g48 ( 
.A(n_26),
.Y(n_48)
);

BUFx3_ASAP7_75t_L g49 ( 
.A(n_38),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_0),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_SL g51 ( 
.A(n_37),
.B(n_25),
.Y(n_51)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_19),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_12),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_9),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_10),
.Y(n_55)
);

INVx4_ASAP7_75t_SL g56 ( 
.A(n_41),
.Y(n_56)
);

CKINVDCx14_ASAP7_75t_R g73 ( 
.A(n_56),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g57 ( 
.A(n_50),
.B(n_0),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_SL g75 ( 
.A(n_57),
.B(n_43),
.Y(n_75)
);

INVx11_ASAP7_75t_L g58 ( 
.A(n_41),
.Y(n_58)
);

BUFx12f_ASAP7_75t_L g70 ( 
.A(n_58),
.Y(n_70)
);

BUFx12f_ASAP7_75t_L g59 ( 
.A(n_40),
.Y(n_59)
);

INVxp67_ASAP7_75t_L g68 ( 
.A(n_59),
.Y(n_68)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_47),
.Y(n_60)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_60),
.Y(n_71)
);

INVx8_ASAP7_75t_L g61 ( 
.A(n_53),
.Y(n_61)
);

AOI22xp33_ASAP7_75t_SL g72 ( 
.A1(n_61),
.A2(n_49),
.B1(n_48),
.B2(n_42),
.Y(n_72)
);

INVx5_ASAP7_75t_L g62 ( 
.A(n_48),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_62),
.B(n_63),
.Y(n_67)
);

BUFx12f_ASAP7_75t_L g63 ( 
.A(n_40),
.Y(n_63)
);

INVx2_ASAP7_75t_L g64 ( 
.A(n_54),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_64),
.B(n_65),
.Y(n_78)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_53),
.Y(n_65)
);

MAJIxp5_ASAP7_75t_L g66 ( 
.A(n_58),
.B(n_47),
.C(n_51),
.Y(n_66)
);

MAJIxp5_ASAP7_75t_L g92 ( 
.A(n_66),
.B(n_72),
.C(n_68),
.Y(n_92)
);

OAI22xp5_ASAP7_75t_L g69 ( 
.A1(n_65),
.A2(n_55),
.B1(n_54),
.B2(n_42),
.Y(n_69)
);

AOI22xp5_ASAP7_75t_L g84 ( 
.A1(n_69),
.A2(n_77),
.B1(n_63),
.B2(n_59),
.Y(n_84)
);

A2O1A1Ixp33_ASAP7_75t_SL g89 ( 
.A1(n_72),
.A2(n_16),
.B(n_36),
.C(n_35),
.Y(n_89)
);

CKINVDCx20_ASAP7_75t_R g74 ( 
.A(n_56),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_74),
.B(n_75),
.Y(n_80)
);

AOI22xp5_ASAP7_75t_SL g76 ( 
.A1(n_62),
.A2(n_55),
.B1(n_43),
.B2(n_46),
.Y(n_76)
);

OAI21xp5_ASAP7_75t_SL g82 ( 
.A1(n_76),
.A2(n_41),
.B(n_63),
.Y(n_82)
);

AOI22xp33_ASAP7_75t_L g77 ( 
.A1(n_61),
.A2(n_46),
.B1(n_45),
.B2(n_49),
.Y(n_77)
);

CKINVDCx20_ASAP7_75t_R g79 ( 
.A(n_59),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_L g86 ( 
.A(n_79),
.B(n_17),
.Y(n_86)
);

AOI22xp33_ASAP7_75t_L g81 ( 
.A1(n_77),
.A2(n_45),
.B1(n_52),
.B2(n_44),
.Y(n_81)
);

OAI22xp5_ASAP7_75t_SL g101 ( 
.A1(n_81),
.A2(n_84),
.B1(n_6),
.B2(n_7),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_SL g97 ( 
.A(n_82),
.B(n_90),
.Y(n_97)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_71),
.Y(n_83)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_83),
.Y(n_102)
);

INVx3_ASAP7_75t_L g85 ( 
.A(n_70),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_L g96 ( 
.A(n_85),
.B(n_87),
.Y(n_96)
);

CKINVDCx14_ASAP7_75t_R g108 ( 
.A(n_86),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_L g87 ( 
.A(n_78),
.B(n_1),
.Y(n_87)
);

INVx1_ASAP7_75t_SL g88 ( 
.A(n_70),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_L g98 ( 
.A(n_88),
.B(n_91),
.Y(n_98)
);

AOI22xp5_ASAP7_75t_L g109 ( 
.A1(n_89),
.A2(n_23),
.B1(n_14),
.B2(n_15),
.Y(n_109)
);

CKINVDCx16_ASAP7_75t_R g90 ( 
.A(n_73),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_L g91 ( 
.A(n_67),
.B(n_1),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_L g103 ( 
.A(n_92),
.B(n_93),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_SL g93 ( 
.A(n_70),
.B(n_2),
.Y(n_93)
);

BUFx3_ASAP7_75t_L g94 ( 
.A(n_68),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_L g110 ( 
.A(n_94),
.B(n_11),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_SL g95 ( 
.A(n_75),
.B(n_2),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g104 ( 
.A(n_95),
.B(n_7),
.Y(n_104)
);

OAI21xp5_ASAP7_75t_L g99 ( 
.A1(n_80),
.A2(n_4),
.B(n_5),
.Y(n_99)
);

INVxp67_ASAP7_75t_SL g114 ( 
.A(n_99),
.Y(n_114)
);

AOI22xp33_ASAP7_75t_L g100 ( 
.A1(n_81),
.A2(n_4),
.B1(n_5),
.B2(n_6),
.Y(n_100)
);

OAI22xp5_ASAP7_75t_L g117 ( 
.A1(n_100),
.A2(n_109),
.B1(n_27),
.B2(n_31),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_SL g111 ( 
.A(n_101),
.B(n_104),
.Y(n_111)
);

AOI21xp5_ASAP7_75t_SL g105 ( 
.A1(n_89),
.A2(n_8),
.B(n_9),
.Y(n_105)
);

O2A1O1Ixp33_ASAP7_75t_L g112 ( 
.A1(n_105),
.A2(n_106),
.B(n_18),
.C(n_21),
.Y(n_112)
);

A2O1A1Ixp33_ASAP7_75t_L g106 ( 
.A1(n_89),
.A2(n_10),
.B(n_11),
.C(n_13),
.Y(n_106)
);

XOR2xp5_ASAP7_75t_L g107 ( 
.A(n_94),
.B(n_24),
.Y(n_107)
);

XNOR2xp5_ASAP7_75t_SL g116 ( 
.A(n_107),
.B(n_22),
.Y(n_116)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_110),
.Y(n_115)
);

XNOR2xp5_ASAP7_75t_L g122 ( 
.A(n_112),
.B(n_113),
.Y(n_122)
);

OAI22xp5_ASAP7_75t_SL g113 ( 
.A1(n_103),
.A2(n_88),
.B1(n_85),
.B2(n_29),
.Y(n_113)
);

MAJIxp5_ASAP7_75t_L g119 ( 
.A(n_116),
.B(n_117),
.C(n_105),
.Y(n_119)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_102),
.Y(n_118)
);

MAJIxp5_ASAP7_75t_L g121 ( 
.A(n_118),
.B(n_107),
.C(n_97),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_L g123 ( 
.A(n_119),
.B(n_120),
.Y(n_123)
);

MAJIxp5_ASAP7_75t_L g120 ( 
.A(n_116),
.B(n_98),
.C(n_96),
.Y(n_120)
);

AOI21xp5_ASAP7_75t_L g124 ( 
.A1(n_121),
.A2(n_115),
.B(n_99),
.Y(n_124)
);

OAI22xp5_ASAP7_75t_SL g125 ( 
.A1(n_124),
.A2(n_114),
.B1(n_109),
.B2(n_100),
.Y(n_125)
);

INVxp67_ASAP7_75t_L g126 ( 
.A(n_125),
.Y(n_126)
);

NAND4xp25_ASAP7_75t_SL g127 ( 
.A(n_126),
.B(n_108),
.C(n_114),
.D(n_112),
.Y(n_127)
);

XNOR2xp5_ASAP7_75t_L g128 ( 
.A(n_127),
.B(n_122),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_L g129 ( 
.A(n_128),
.B(n_123),
.Y(n_129)
);

A2O1A1O1Ixp25_ASAP7_75t_L g130 ( 
.A1(n_129),
.A2(n_111),
.B(n_106),
.C(n_39),
.D(n_32),
.Y(n_130)
);


endmodule