module fake_jpeg_20774_n_52 (n_13, n_21, n_1, n_10, n_6, n_14, n_19, n_18, n_20, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_52);

input n_13;
input n_21;
input n_1;
input n_10;
input n_6;
input n_14;
input n_19;
input n_18;
input n_20;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_52;

wire n_33;
wire n_45;
wire n_23;
wire n_27;
wire n_22;
wire n_47;
wire n_51;
wire n_40;
wire n_48;
wire n_35;
wire n_46;
wire n_41;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_49;
wire n_24;
wire n_28;
wire n_38;
wire n_26;
wire n_44;
wire n_36;
wire n_31;
wire n_25;
wire n_29;
wire n_37;
wire n_43;
wire n_50;
wire n_32;

INVx6_ASAP7_75t_L g22 ( 
.A(n_13),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_0),
.Y(n_23)
);

BUFx12f_ASAP7_75t_L g24 ( 
.A(n_10),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_17),
.Y(n_25)
);

NAND2xp5_ASAP7_75t_L g26 ( 
.A(n_19),
.B(n_5),
.Y(n_26)
);

BUFx8_ASAP7_75t_L g27 ( 
.A(n_4),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_11),
.Y(n_28)
);

NAND2xp5_ASAP7_75t_L g29 ( 
.A(n_26),
.B(n_0),
.Y(n_29)
);

NAND2xp5_ASAP7_75t_SL g38 ( 
.A(n_29),
.B(n_32),
.Y(n_38)
);

BUFx12f_ASAP7_75t_L g30 ( 
.A(n_27),
.Y(n_30)
);

NOR2xp33_ASAP7_75t_L g35 ( 
.A(n_30),
.B(n_33),
.Y(n_35)
);

AOI22xp33_ASAP7_75t_SL g31 ( 
.A1(n_22),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_31)
);

CKINVDCx14_ASAP7_75t_R g39 ( 
.A(n_31),
.Y(n_39)
);

AND2x2_ASAP7_75t_SL g32 ( 
.A(n_26),
.B(n_12),
.Y(n_32)
);

INVx2_ASAP7_75t_L g33 ( 
.A(n_24),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_L g34 ( 
.A(n_23),
.B(n_28),
.Y(n_34)
);

CKINVDCx16_ASAP7_75t_R g40 ( 
.A(n_34),
.Y(n_40)
);

OAI21xp5_ASAP7_75t_L g36 ( 
.A1(n_32),
.A2(n_24),
.B(n_27),
.Y(n_36)
);

XNOR2xp5_ASAP7_75t_L g42 ( 
.A(n_36),
.B(n_25),
.Y(n_42)
);

MAJIxp5_ASAP7_75t_SL g37 ( 
.A(n_30),
.B(n_1),
.C(n_2),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_SL g41 ( 
.A(n_37),
.B(n_3),
.Y(n_41)
);

INVxp67_ASAP7_75t_L g45 ( 
.A(n_41),
.Y(n_45)
);

XOR2xp5_ASAP7_75t_L g46 ( 
.A(n_42),
.B(n_43),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g43 ( 
.A(n_38),
.B(n_6),
.Y(n_43)
);

XOR2x2_ASAP7_75t_L g44 ( 
.A(n_36),
.B(n_7),
.Y(n_44)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_46),
.Y(n_47)
);

AO21x1_ASAP7_75t_L g48 ( 
.A1(n_47),
.A2(n_44),
.B(n_43),
.Y(n_48)
);

OAI22xp5_ASAP7_75t_L g49 ( 
.A1(n_48),
.A2(n_45),
.B1(n_39),
.B2(n_40),
.Y(n_49)
);

AOI322xp5_ASAP7_75t_L g50 ( 
.A1(n_49),
.A2(n_35),
.A3(n_9),
.B1(n_14),
.B2(n_15),
.C1(n_8),
.C2(n_18),
.Y(n_50)
);

AOI21xp5_ASAP7_75t_L g51 ( 
.A1(n_50),
.A2(n_16),
.B(n_20),
.Y(n_51)
);

NOR2x1_ASAP7_75t_L g52 ( 
.A(n_51),
.B(n_21),
.Y(n_52)
);


endmodule