module fake_jpeg_10357_n_337 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_337);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_337;

wire n_253;
wire n_330;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_265;
wire n_192;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_11),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_10),
.Y(n_17)
);

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_7),
.Y(n_18)
);

INVx3_ASAP7_75t_L g19 ( 
.A(n_7),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_11),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_3),
.Y(n_21)
);

HB1xp67_ASAP7_75t_L g22 ( 
.A(n_0),
.Y(n_22)
);

BUFx3_ASAP7_75t_L g23 ( 
.A(n_2),
.Y(n_23)
);

INVx2_ASAP7_75t_L g24 ( 
.A(n_6),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_14),
.Y(n_25)
);

INVx8_ASAP7_75t_L g26 ( 
.A(n_15),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_12),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_7),
.Y(n_28)
);

BUFx12f_ASAP7_75t_L g29 ( 
.A(n_12),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_7),
.Y(n_30)
);

BUFx5_ASAP7_75t_L g31 ( 
.A(n_13),
.Y(n_31)
);

BUFx12f_ASAP7_75t_L g32 ( 
.A(n_2),
.Y(n_32)
);

BUFx12f_ASAP7_75t_L g33 ( 
.A(n_10),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_14),
.Y(n_34)
);

BUFx12f_ASAP7_75t_L g35 ( 
.A(n_1),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_32),
.Y(n_36)
);

INVx6_ASAP7_75t_L g59 ( 
.A(n_36),
.Y(n_59)
);

INVx8_ASAP7_75t_L g37 ( 
.A(n_31),
.Y(n_37)
);

INVx11_ASAP7_75t_L g58 ( 
.A(n_37),
.Y(n_58)
);

BUFx12f_ASAP7_75t_L g38 ( 
.A(n_31),
.Y(n_38)
);

INVx4_ASAP7_75t_L g51 ( 
.A(n_38),
.Y(n_51)
);

HB1xp67_ASAP7_75t_L g39 ( 
.A(n_23),
.Y(n_39)
);

INVx2_ASAP7_75t_L g49 ( 
.A(n_39),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_L g40 ( 
.A(n_30),
.B(n_0),
.Y(n_40)
);

NAND2xp5_ASAP7_75t_L g56 ( 
.A(n_40),
.B(n_21),
.Y(n_56)
);

INVx3_ASAP7_75t_L g41 ( 
.A(n_25),
.Y(n_41)
);

INVx4_ASAP7_75t_L g53 ( 
.A(n_41),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_35),
.Y(n_42)
);

INVx3_ASAP7_75t_SL g61 ( 
.A(n_42),
.Y(n_61)
);

AOI22xp5_ASAP7_75t_L g43 ( 
.A1(n_24),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_43)
);

OAI22xp5_ASAP7_75t_L g65 ( 
.A1(n_43),
.A2(n_26),
.B1(n_28),
.B2(n_19),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g44 ( 
.A(n_16),
.B(n_15),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_44),
.B(n_47),
.Y(n_67)
);

INVx5_ASAP7_75t_L g45 ( 
.A(n_23),
.Y(n_45)
);

INVx5_ASAP7_75t_L g66 ( 
.A(n_45),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_32),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_46),
.Y(n_48)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_17),
.Y(n_47)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_40),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_50),
.B(n_52),
.Y(n_83)
);

OR2x2_ASAP7_75t_L g52 ( 
.A(n_44),
.B(n_27),
.Y(n_52)
);

INVx2_ASAP7_75t_L g54 ( 
.A(n_39),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_54),
.B(n_55),
.Y(n_84)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_47),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_SL g80 ( 
.A(n_56),
.B(n_63),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_L g57 ( 
.A(n_43),
.B(n_24),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_L g77 ( 
.A(n_57),
.B(n_64),
.Y(n_77)
);

INVx4_ASAP7_75t_L g60 ( 
.A(n_41),
.Y(n_60)
);

INVx8_ASAP7_75t_L g106 ( 
.A(n_60),
.Y(n_106)
);

AOI22xp33_ASAP7_75t_SL g62 ( 
.A1(n_41),
.A2(n_26),
.B1(n_19),
.B2(n_17),
.Y(n_62)
);

AOI22xp33_ASAP7_75t_SL g85 ( 
.A1(n_62),
.A2(n_26),
.B1(n_45),
.B2(n_37),
.Y(n_85)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_43),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_L g64 ( 
.A(n_42),
.B(n_21),
.Y(n_64)
);

AOI22xp5_ASAP7_75t_L g110 ( 
.A1(n_65),
.A2(n_29),
.B1(n_33),
.B2(n_32),
.Y(n_110)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_38),
.Y(n_68)
);

BUFx6f_ASAP7_75t_L g103 ( 
.A(n_68),
.Y(n_103)
);

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_38),
.Y(n_69)
);

BUFx2_ASAP7_75t_L g73 ( 
.A(n_69),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_L g70 ( 
.A(n_42),
.B(n_28),
.Y(n_70)
);

AOI21xp33_ASAP7_75t_L g92 ( 
.A1(n_70),
.A2(n_30),
.B(n_20),
.Y(n_92)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_42),
.Y(n_71)
);

AND2x2_ASAP7_75t_L g88 ( 
.A(n_71),
.B(n_72),
.Y(n_88)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_36),
.Y(n_72)
);

INVx2_ASAP7_75t_L g74 ( 
.A(n_66),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g121 ( 
.A(n_74),
.B(n_78),
.Y(n_121)
);

OAI22xp5_ASAP7_75t_L g75 ( 
.A1(n_63),
.A2(n_57),
.B1(n_65),
.B2(n_50),
.Y(n_75)
);

OAI22xp5_ASAP7_75t_SL g131 ( 
.A1(n_75),
.A2(n_90),
.B1(n_91),
.B2(n_94),
.Y(n_131)
);

INVxp67_ASAP7_75t_L g76 ( 
.A(n_61),
.Y(n_76)
);

INVxp67_ASAP7_75t_L g113 ( 
.A(n_76),
.Y(n_113)
);

CKINVDCx20_ASAP7_75t_R g78 ( 
.A(n_59),
.Y(n_78)
);

INVxp67_ASAP7_75t_L g79 ( 
.A(n_61),
.Y(n_79)
);

INVxp67_ASAP7_75t_L g120 ( 
.A(n_79),
.Y(n_120)
);

CKINVDCx20_ASAP7_75t_R g81 ( 
.A(n_59),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_81),
.B(n_48),
.Y(n_127)
);

BUFx3_ASAP7_75t_L g82 ( 
.A(n_61),
.Y(n_82)
);

INVx3_ASAP7_75t_L g132 ( 
.A(n_82),
.Y(n_132)
);

OAI22xp33_ASAP7_75t_SL g141 ( 
.A1(n_85),
.A2(n_9),
.B1(n_14),
.B2(n_13),
.Y(n_141)
);

INVxp67_ASAP7_75t_L g86 ( 
.A(n_64),
.Y(n_86)
);

INVxp67_ASAP7_75t_L g136 ( 
.A(n_86),
.Y(n_136)
);

BUFx12f_ASAP7_75t_L g87 ( 
.A(n_68),
.Y(n_87)
);

INVx3_ASAP7_75t_L g135 ( 
.A(n_87),
.Y(n_135)
);

AND2x2_ASAP7_75t_L g89 ( 
.A(n_55),
.B(n_22),
.Y(n_89)
);

AOI21xp5_ASAP7_75t_L g122 ( 
.A1(n_89),
.A2(n_29),
.B(n_52),
.Y(n_122)
);

OAI22xp5_ASAP7_75t_L g90 ( 
.A1(n_56),
.A2(n_45),
.B1(n_37),
.B2(n_16),
.Y(n_90)
);

AOI22xp33_ASAP7_75t_L g91 ( 
.A1(n_53),
.A2(n_60),
.B1(n_66),
.B2(n_27),
.Y(n_91)
);

OAI21xp5_ASAP7_75t_SL g117 ( 
.A1(n_92),
.A2(n_52),
.B(n_29),
.Y(n_117)
);

INVx2_ASAP7_75t_L g93 ( 
.A(n_58),
.Y(n_93)
);

INVx3_ASAP7_75t_SL g119 ( 
.A(n_93),
.Y(n_119)
);

AOI22xp5_ASAP7_75t_SL g94 ( 
.A1(n_58),
.A2(n_20),
.B1(n_22),
.B2(n_25),
.Y(n_94)
);

AOI22xp5_ASAP7_75t_SL g95 ( 
.A1(n_59),
.A2(n_25),
.B1(n_34),
.B2(n_23),
.Y(n_95)
);

OAI21xp5_ASAP7_75t_L g133 ( 
.A1(n_95),
.A2(n_38),
.B(n_69),
.Y(n_133)
);

INVx2_ASAP7_75t_L g96 ( 
.A(n_49),
.Y(n_96)
);

CKINVDCx16_ASAP7_75t_R g116 ( 
.A(n_96),
.Y(n_116)
);

OAI22xp5_ASAP7_75t_L g97 ( 
.A1(n_53),
.A2(n_18),
.B1(n_34),
.B2(n_35),
.Y(n_97)
);

AOI22xp5_ASAP7_75t_L g112 ( 
.A1(n_97),
.A2(n_100),
.B1(n_101),
.B2(n_102),
.Y(n_112)
);

INVx2_ASAP7_75t_L g98 ( 
.A(n_49),
.Y(n_98)
);

CKINVDCx16_ASAP7_75t_R g130 ( 
.A(n_98),
.Y(n_130)
);

INVx2_ASAP7_75t_L g99 ( 
.A(n_54),
.Y(n_99)
);

CKINVDCx20_ASAP7_75t_R g124 ( 
.A(n_99),
.Y(n_124)
);

OAI22xp5_ASAP7_75t_L g100 ( 
.A1(n_70),
.A2(n_18),
.B1(n_34),
.B2(n_35),
.Y(n_100)
);

OAI22xp5_ASAP7_75t_L g101 ( 
.A1(n_67),
.A2(n_18),
.B1(n_32),
.B2(n_35),
.Y(n_101)
);

OAI22xp5_ASAP7_75t_L g102 ( 
.A1(n_67),
.A2(n_35),
.B1(n_32),
.B2(n_29),
.Y(n_102)
);

CKINVDCx16_ASAP7_75t_R g104 ( 
.A(n_68),
.Y(n_104)
);

AOI22xp33_ASAP7_75t_SL g128 ( 
.A1(n_104),
.A2(n_107),
.B1(n_109),
.B2(n_9),
.Y(n_128)
);

INVx2_ASAP7_75t_L g105 ( 
.A(n_48),
.Y(n_105)
);

CKINVDCx20_ASAP7_75t_R g126 ( 
.A(n_105),
.Y(n_126)
);

AOI22xp33_ASAP7_75t_SL g107 ( 
.A1(n_51),
.A2(n_11),
.B1(n_9),
.B2(n_10),
.Y(n_107)
);

INVx2_ASAP7_75t_L g108 ( 
.A(n_48),
.Y(n_108)
);

CKINVDCx20_ASAP7_75t_R g137 ( 
.A(n_108),
.Y(n_137)
);

INVx1_ASAP7_75t_SL g109 ( 
.A(n_51),
.Y(n_109)
);

AOI22xp33_ASAP7_75t_L g138 ( 
.A1(n_110),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_138)
);

INVxp67_ASAP7_75t_L g111 ( 
.A(n_69),
.Y(n_111)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_111),
.Y(n_118)
);

AND2x2_ASAP7_75t_L g114 ( 
.A(n_80),
.B(n_71),
.Y(n_114)
);

OAI21xp5_ASAP7_75t_SL g174 ( 
.A1(n_114),
.A2(n_122),
.B(n_123),
.Y(n_174)
);

AOI22xp5_ASAP7_75t_L g115 ( 
.A1(n_75),
.A2(n_72),
.B1(n_46),
.B2(n_36),
.Y(n_115)
);

OAI22xp5_ASAP7_75t_SL g143 ( 
.A1(n_115),
.A2(n_140),
.B1(n_94),
.B2(n_95),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_SL g146 ( 
.A(n_117),
.B(n_90),
.Y(n_146)
);

AOI21xp5_ASAP7_75t_SL g123 ( 
.A1(n_89),
.A2(n_29),
.B(n_33),
.Y(n_123)
);

OAI21xp5_ASAP7_75t_SL g125 ( 
.A1(n_80),
.A2(n_46),
.B(n_33),
.Y(n_125)
);

MAJIxp5_ASAP7_75t_L g152 ( 
.A(n_125),
.B(n_129),
.C(n_102),
.Y(n_152)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_127),
.Y(n_150)
);

AOI22xp33_ASAP7_75t_L g148 ( 
.A1(n_128),
.A2(n_133),
.B1(n_74),
.B2(n_93),
.Y(n_148)
);

OAI21xp5_ASAP7_75t_SL g129 ( 
.A1(n_77),
.A2(n_33),
.B(n_38),
.Y(n_129)
);

OR2x2_ASAP7_75t_L g134 ( 
.A(n_83),
.B(n_0),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_L g154 ( 
.A(n_134),
.B(n_139),
.Y(n_154)
);

OAI22xp5_ASAP7_75t_L g172 ( 
.A1(n_138),
.A2(n_108),
.B1(n_105),
.B2(n_12),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_L g139 ( 
.A(n_77),
.B(n_1),
.Y(n_139)
);

AOI22xp5_ASAP7_75t_L g140 ( 
.A1(n_110),
.A2(n_3),
.B1(n_4),
.B2(n_5),
.Y(n_140)
);

AOI22xp5_ASAP7_75t_SL g165 ( 
.A1(n_141),
.A2(n_106),
.B1(n_15),
.B2(n_13),
.Y(n_165)
);

OR2x2_ASAP7_75t_L g142 ( 
.A(n_115),
.B(n_83),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_L g175 ( 
.A(n_142),
.B(n_159),
.Y(n_175)
);

AOI22xp5_ASAP7_75t_L g191 ( 
.A1(n_143),
.A2(n_145),
.B1(n_155),
.B2(n_164),
.Y(n_191)
);

OAI21xp5_ASAP7_75t_L g144 ( 
.A1(n_122),
.A2(n_84),
.B(n_89),
.Y(n_144)
);

OAI21xp5_ASAP7_75t_SL g176 ( 
.A1(n_144),
.A2(n_123),
.B(n_131),
.Y(n_176)
);

OAI22xp5_ASAP7_75t_SL g145 ( 
.A1(n_112),
.A2(n_92),
.B1(n_81),
.B2(n_78),
.Y(n_145)
);

OAI21xp5_ASAP7_75t_L g197 ( 
.A1(n_146),
.A2(n_152),
.B(n_137),
.Y(n_197)
);

NOR2xp33_ASAP7_75t_SL g147 ( 
.A(n_134),
.B(n_84),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_SL g203 ( 
.A(n_147),
.B(n_149),
.Y(n_203)
);

OAI22xp5_ASAP7_75t_L g181 ( 
.A1(n_148),
.A2(n_128),
.B1(n_133),
.B2(n_140),
.Y(n_181)
);

CKINVDCx20_ASAP7_75t_R g149 ( 
.A(n_121),
.Y(n_149)
);

NOR2xp33_ASAP7_75t_L g151 ( 
.A(n_121),
.B(n_96),
.Y(n_151)
);

CKINVDCx16_ASAP7_75t_R g200 ( 
.A(n_151),
.Y(n_200)
);

NOR2xp33_ASAP7_75t_L g153 ( 
.A(n_134),
.B(n_98),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_SL g204 ( 
.A(n_153),
.B(n_157),
.Y(n_204)
);

OAI22xp5_ASAP7_75t_SL g155 ( 
.A1(n_112),
.A2(n_100),
.B1(n_106),
.B2(n_101),
.Y(n_155)
);

MAJIxp5_ASAP7_75t_L g156 ( 
.A(n_129),
.B(n_109),
.C(n_97),
.Y(n_156)
);

MAJIxp5_ASAP7_75t_L g190 ( 
.A(n_156),
.B(n_118),
.C(n_130),
.Y(n_190)
);

NOR2xp33_ASAP7_75t_L g157 ( 
.A(n_127),
.B(n_139),
.Y(n_157)
);

NOR2xp33_ASAP7_75t_L g158 ( 
.A(n_115),
.B(n_99),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_SL g206 ( 
.A(n_158),
.B(n_160),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_L g159 ( 
.A(n_114),
.B(n_88),
.Y(n_159)
);

CKINVDCx20_ASAP7_75t_R g160 ( 
.A(n_119),
.Y(n_160)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_119),
.Y(n_161)
);

NOR2xp33_ASAP7_75t_L g186 ( 
.A(n_161),
.B(n_162),
.Y(n_186)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_119),
.Y(n_162)
);

A2O1A1Ixp33_ASAP7_75t_L g163 ( 
.A1(n_117),
.A2(n_88),
.B(n_82),
.C(n_5),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_L g179 ( 
.A(n_163),
.B(n_166),
.Y(n_179)
);

OAI22xp5_ASAP7_75t_SL g164 ( 
.A1(n_112),
.A2(n_106),
.B1(n_88),
.B2(n_104),
.Y(n_164)
);

NOR2xp33_ASAP7_75t_L g187 ( 
.A(n_165),
.B(n_167),
.Y(n_187)
);

NOR2xp33_ASAP7_75t_L g166 ( 
.A(n_124),
.B(n_87),
.Y(n_166)
);

INVx4_ASAP7_75t_L g167 ( 
.A(n_135),
.Y(n_167)
);

NOR2xp33_ASAP7_75t_L g168 ( 
.A(n_124),
.B(n_118),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_L g182 ( 
.A(n_168),
.B(n_171),
.Y(n_182)
);

NOR3xp33_ASAP7_75t_SL g169 ( 
.A(n_123),
.B(n_73),
.C(n_87),
.Y(n_169)
);

NOR2xp33_ASAP7_75t_L g189 ( 
.A(n_169),
.B(n_170),
.Y(n_189)
);

INVx4_ASAP7_75t_L g170 ( 
.A(n_135),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_SL g171 ( 
.A(n_114),
.B(n_3),
.Y(n_171)
);

AOI22xp5_ASAP7_75t_L g194 ( 
.A1(n_172),
.A2(n_132),
.B1(n_113),
.B2(n_120),
.Y(n_194)
);

CKINVDCx20_ASAP7_75t_R g173 ( 
.A(n_119),
.Y(n_173)
);

NOR2xp33_ASAP7_75t_L g195 ( 
.A(n_173),
.B(n_160),
.Y(n_195)
);

XNOR2xp5_ASAP7_75t_SL g214 ( 
.A(n_176),
.B(n_180),
.Y(n_214)
);

OAI22xp5_ASAP7_75t_SL g177 ( 
.A1(n_146),
.A2(n_133),
.B1(n_140),
.B2(n_138),
.Y(n_177)
);

AOI22xp5_ASAP7_75t_L g215 ( 
.A1(n_177),
.A2(n_181),
.B1(n_192),
.B2(n_143),
.Y(n_215)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_151),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_SL g222 ( 
.A(n_178),
.B(n_184),
.Y(n_222)
);

XNOR2xp5_ASAP7_75t_L g180 ( 
.A(n_174),
.B(n_152),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_L g183 ( 
.A(n_157),
.B(n_114),
.Y(n_183)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_183),
.Y(n_218)
);

INVxp67_ASAP7_75t_L g184 ( 
.A(n_166),
.Y(n_184)
);

XOR2xp5_ASAP7_75t_L g185 ( 
.A(n_174),
.B(n_125),
.Y(n_185)
);

XOR2xp5_ASAP7_75t_L g216 ( 
.A(n_185),
.B(n_196),
.Y(n_216)
);

OAI22xp5_ASAP7_75t_L g188 ( 
.A1(n_156),
.A2(n_131),
.B1(n_136),
.B2(n_132),
.Y(n_188)
);

OAI22xp5_ASAP7_75t_SL g232 ( 
.A1(n_188),
.A2(n_194),
.B1(n_208),
.B2(n_163),
.Y(n_232)
);

XNOR2xp5_ASAP7_75t_L g217 ( 
.A(n_190),
.B(n_197),
.Y(n_217)
);

OAI22xp5_ASAP7_75t_SL g192 ( 
.A1(n_158),
.A2(n_132),
.B1(n_141),
.B2(n_116),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_L g193 ( 
.A(n_150),
.B(n_130),
.Y(n_193)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_193),
.Y(n_220)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_195),
.Y(n_224)
);

XOR2xp5_ASAP7_75t_L g196 ( 
.A(n_144),
.B(n_116),
.Y(n_196)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_168),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_SL g234 ( 
.A(n_198),
.B(n_205),
.Y(n_234)
);

XNOR2xp5_ASAP7_75t_L g199 ( 
.A(n_159),
.B(n_137),
.Y(n_199)
);

XNOR2xp5_ASAP7_75t_L g227 ( 
.A(n_199),
.B(n_202),
.Y(n_227)
);

NOR2xp33_ASAP7_75t_L g201 ( 
.A(n_167),
.B(n_135),
.Y(n_201)
);

NOR2xp33_ASAP7_75t_SL g230 ( 
.A(n_201),
.B(n_207),
.Y(n_230)
);

XOR2xp5_ASAP7_75t_L g202 ( 
.A(n_145),
.B(n_171),
.Y(n_202)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_164),
.Y(n_205)
);

NOR2xp33_ASAP7_75t_L g207 ( 
.A(n_167),
.B(n_170),
.Y(n_207)
);

OAI22xp5_ASAP7_75t_L g208 ( 
.A1(n_150),
.A2(n_126),
.B1(n_103),
.B2(n_73),
.Y(n_208)
);

INVx1_ASAP7_75t_SL g209 ( 
.A(n_193),
.Y(n_209)
);

AOI22xp33_ASAP7_75t_SL g237 ( 
.A1(n_209),
.A2(n_212),
.B1(n_218),
.B2(n_225),
.Y(n_237)
);

CKINVDCx20_ASAP7_75t_R g210 ( 
.A(n_186),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_SL g240 ( 
.A(n_210),
.B(n_213),
.Y(n_240)
);

NAND2xp5_ASAP7_75t_L g211 ( 
.A(n_203),
.B(n_154),
.Y(n_211)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_211),
.Y(n_250)
);

INVx1_ASAP7_75t_SL g212 ( 
.A(n_179),
.Y(n_212)
);

CKINVDCx20_ASAP7_75t_R g213 ( 
.A(n_208),
.Y(n_213)
);

OAI22xp5_ASAP7_75t_SL g246 ( 
.A1(n_215),
.A2(n_221),
.B1(n_191),
.B2(n_197),
.Y(n_246)
);

AOI22xp5_ASAP7_75t_SL g219 ( 
.A1(n_205),
.A2(n_169),
.B1(n_149),
.B2(n_163),
.Y(n_219)
);

OAI21xp5_ASAP7_75t_L g260 ( 
.A1(n_219),
.A2(n_4),
.B(n_5),
.Y(n_260)
);

AOI22xp5_ASAP7_75t_L g221 ( 
.A1(n_177),
.A2(n_155),
.B1(n_142),
.B2(n_147),
.Y(n_221)
);

NOR2xp33_ASAP7_75t_L g223 ( 
.A(n_198),
.B(n_170),
.Y(n_223)
);

NOR2xp33_ASAP7_75t_SL g244 ( 
.A(n_223),
.B(n_226),
.Y(n_244)
);

CKINVDCx20_ASAP7_75t_R g225 ( 
.A(n_206),
.Y(n_225)
);

NAND2xp5_ASAP7_75t_L g238 ( 
.A(n_225),
.B(n_229),
.Y(n_238)
);

NOR2xp33_ASAP7_75t_L g226 ( 
.A(n_178),
.B(n_142),
.Y(n_226)
);

NOR2xp33_ASAP7_75t_L g228 ( 
.A(n_192),
.B(n_173),
.Y(n_228)
);

CKINVDCx16_ASAP7_75t_R g245 ( 
.A(n_228),
.Y(n_245)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_204),
.Y(n_229)
);

NAND2xp5_ASAP7_75t_L g231 ( 
.A(n_183),
.B(n_154),
.Y(n_231)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_231),
.Y(n_251)
);

AOI22xp5_ASAP7_75t_L g242 ( 
.A1(n_232),
.A2(n_189),
.B1(n_181),
.B2(n_187),
.Y(n_242)
);

NOR2xp33_ASAP7_75t_L g233 ( 
.A(n_200),
.B(n_162),
.Y(n_233)
);

INVxp67_ASAP7_75t_L g259 ( 
.A(n_233),
.Y(n_259)
);

NAND2xp5_ASAP7_75t_SL g235 ( 
.A(n_184),
.B(n_161),
.Y(n_235)
);

CKINVDCx20_ASAP7_75t_R g241 ( 
.A(n_235),
.Y(n_241)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_175),
.Y(n_236)
);

NAND2xp5_ASAP7_75t_L g239 ( 
.A(n_236),
.B(n_175),
.Y(n_239)
);

OAI22xp5_ASAP7_75t_L g262 ( 
.A1(n_237),
.A2(n_242),
.B1(n_243),
.B2(n_253),
.Y(n_262)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_239),
.Y(n_265)
);

AOI22xp5_ASAP7_75t_SL g243 ( 
.A1(n_213),
.A2(n_185),
.B1(n_176),
.B2(n_188),
.Y(n_243)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_246),
.Y(n_272)
);

OAI22xp5_ASAP7_75t_L g247 ( 
.A1(n_215),
.A2(n_191),
.B1(n_194),
.B2(n_179),
.Y(n_247)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_247),
.Y(n_274)
);

XOR2xp5_ASAP7_75t_L g248 ( 
.A(n_216),
.B(n_180),
.Y(n_248)
);

XOR2xp5_ASAP7_75t_L g267 ( 
.A(n_248),
.B(n_260),
.Y(n_267)
);

NAND2xp5_ASAP7_75t_L g249 ( 
.A(n_211),
.B(n_199),
.Y(n_249)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_249),
.Y(n_275)
);

OAI22xp5_ASAP7_75t_L g252 ( 
.A1(n_234),
.A2(n_190),
.B1(n_165),
.B2(n_182),
.Y(n_252)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_252),
.Y(n_279)
);

AOI22xp5_ASAP7_75t_L g253 ( 
.A1(n_232),
.A2(n_196),
.B1(n_202),
.B2(n_153),
.Y(n_253)
);

NAND2xp5_ASAP7_75t_L g254 ( 
.A(n_209),
.B(n_182),
.Y(n_254)
);

NAND2xp5_ASAP7_75t_L g268 ( 
.A(n_254),
.B(n_255),
.Y(n_268)
);

AOI22xp5_ASAP7_75t_L g255 ( 
.A1(n_212),
.A2(n_172),
.B1(n_126),
.B2(n_103),
.Y(n_255)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_222),
.Y(n_256)
);

NAND2xp5_ASAP7_75t_L g280 ( 
.A(n_256),
.B(n_258),
.Y(n_280)
);

XNOR2xp5_ASAP7_75t_L g257 ( 
.A(n_214),
.B(n_73),
.Y(n_257)
);

MAJIxp5_ASAP7_75t_L g263 ( 
.A(n_257),
.B(n_214),
.C(n_216),
.Y(n_263)
);

CKINVDCx20_ASAP7_75t_R g258 ( 
.A(n_230),
.Y(n_258)
);

NOR2xp33_ASAP7_75t_SL g261 ( 
.A(n_258),
.B(n_229),
.Y(n_261)
);

NAND2xp5_ASAP7_75t_SL g296 ( 
.A(n_261),
.B(n_277),
.Y(n_296)
);

XOR2xp5_ASAP7_75t_L g294 ( 
.A(n_263),
.B(n_271),
.Y(n_294)
);

MAJIxp5_ASAP7_75t_L g264 ( 
.A(n_248),
.B(n_217),
.C(n_227),
.Y(n_264)
);

MAJIxp5_ASAP7_75t_L g284 ( 
.A(n_264),
.B(n_266),
.C(n_273),
.Y(n_284)
);

MAJIxp5_ASAP7_75t_L g266 ( 
.A(n_257),
.B(n_217),
.C(n_227),
.Y(n_266)
);

INVx2_ASAP7_75t_SL g269 ( 
.A(n_259),
.Y(n_269)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_269),
.Y(n_286)
);

NOR2xp33_ASAP7_75t_L g270 ( 
.A(n_244),
.B(n_224),
.Y(n_270)
);

CKINVDCx14_ASAP7_75t_R g292 ( 
.A(n_270),
.Y(n_292)
);

XNOR2xp5_ASAP7_75t_L g271 ( 
.A(n_243),
.B(n_221),
.Y(n_271)
);

MAJIxp5_ASAP7_75t_L g273 ( 
.A(n_253),
.B(n_249),
.C(n_246),
.Y(n_273)
);

MAJIxp5_ASAP7_75t_L g276 ( 
.A(n_238),
.B(n_220),
.C(n_218),
.Y(n_276)
);

MAJIxp5_ASAP7_75t_L g291 ( 
.A(n_276),
.B(n_278),
.C(n_4),
.Y(n_291)
);

NAND2xp5_ASAP7_75t_SL g277 ( 
.A(n_259),
.B(n_224),
.Y(n_277)
);

MAJIxp5_ASAP7_75t_L g278 ( 
.A(n_238),
.B(n_220),
.C(n_231),
.Y(n_278)
);

AOI21xp5_ASAP7_75t_L g281 ( 
.A1(n_272),
.A2(n_245),
.B(n_240),
.Y(n_281)
);

INVxp67_ASAP7_75t_L g301 ( 
.A(n_281),
.Y(n_301)
);

NAND2xp5_ASAP7_75t_L g282 ( 
.A(n_280),
.B(n_250),
.Y(n_282)
);

CKINVDCx20_ASAP7_75t_R g299 ( 
.A(n_282),
.Y(n_299)
);

AOI22xp5_ASAP7_75t_L g283 ( 
.A1(n_274),
.A2(n_251),
.B1(n_250),
.B2(n_236),
.Y(n_283)
);

AOI22xp5_ASAP7_75t_L g309 ( 
.A1(n_283),
.A2(n_288),
.B1(n_289),
.B2(n_293),
.Y(n_309)
);

AOI21xp5_ASAP7_75t_L g285 ( 
.A1(n_268),
.A2(n_241),
.B(n_239),
.Y(n_285)
);

NOR2xp33_ASAP7_75t_L g308 ( 
.A(n_285),
.B(n_8),
.Y(n_308)
);

NAND2xp5_ASAP7_75t_L g287 ( 
.A(n_280),
.B(n_241),
.Y(n_287)
);

CKINVDCx20_ASAP7_75t_R g304 ( 
.A(n_287),
.Y(n_304)
);

OAI22xp5_ASAP7_75t_SL g288 ( 
.A1(n_279),
.A2(n_242),
.B1(n_251),
.B2(n_255),
.Y(n_288)
);

OAI22xp5_ASAP7_75t_SL g289 ( 
.A1(n_268),
.A2(n_219),
.B1(n_254),
.B2(n_256),
.Y(n_289)
);

OR2x2_ASAP7_75t_L g290 ( 
.A(n_265),
.B(n_260),
.Y(n_290)
);

NAND2xp5_ASAP7_75t_L g310 ( 
.A(n_290),
.B(n_295),
.Y(n_310)
);

MAJIxp5_ASAP7_75t_L g297 ( 
.A(n_291),
.B(n_275),
.C(n_267),
.Y(n_297)
);

OAI22xp5_ASAP7_75t_SL g293 ( 
.A1(n_276),
.A2(n_103),
.B1(n_87),
.B2(n_6),
.Y(n_293)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_278),
.Y(n_295)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_297),
.Y(n_313)
);

XNOR2xp5_ASAP7_75t_L g298 ( 
.A(n_284),
.B(n_273),
.Y(n_298)
);

MAJIxp5_ASAP7_75t_L g311 ( 
.A(n_298),
.B(n_303),
.C(n_305),
.Y(n_311)
);

NAND2xp5_ASAP7_75t_SL g300 ( 
.A(n_292),
.B(n_271),
.Y(n_300)
);

NAND2xp5_ASAP7_75t_SL g319 ( 
.A(n_300),
.B(n_306),
.Y(n_319)
);

XOR2xp5_ASAP7_75t_L g302 ( 
.A(n_294),
.B(n_264),
.Y(n_302)
);

XOR2xp5_ASAP7_75t_L g312 ( 
.A(n_302),
.B(n_294),
.Y(n_312)
);

MAJIxp5_ASAP7_75t_L g303 ( 
.A(n_284),
.B(n_266),
.C(n_263),
.Y(n_303)
);

MAJIxp5_ASAP7_75t_L g305 ( 
.A(n_295),
.B(n_267),
.C(n_262),
.Y(n_305)
);

AOI322xp5_ASAP7_75t_SL g306 ( 
.A1(n_289),
.A2(n_4),
.A3(n_5),
.B1(n_6),
.B2(n_8),
.C1(n_269),
.C2(n_296),
.Y(n_306)
);

MAJIxp5_ASAP7_75t_L g307 ( 
.A(n_291),
.B(n_6),
.C(n_8),
.Y(n_307)
);

MAJIxp5_ASAP7_75t_L g318 ( 
.A(n_307),
.B(n_287),
.C(n_293),
.Y(n_318)
);

OR2x2_ASAP7_75t_L g317 ( 
.A(n_308),
.B(n_8),
.Y(n_317)
);

MAJIxp5_ASAP7_75t_L g324 ( 
.A(n_312),
.B(n_314),
.C(n_320),
.Y(n_324)
);

XOR2xp5_ASAP7_75t_L g314 ( 
.A(n_302),
.B(n_288),
.Y(n_314)
);

AND2x2_ASAP7_75t_L g315 ( 
.A(n_305),
.B(n_286),
.Y(n_315)
);

AOI322xp5_ASAP7_75t_L g327 ( 
.A1(n_315),
.A2(n_310),
.A3(n_282),
.B1(n_297),
.B2(n_309),
.C1(n_290),
.C2(n_283),
.Y(n_327)
);

XNOR2xp5_ASAP7_75t_L g316 ( 
.A(n_298),
.B(n_281),
.Y(n_316)
);

NOR2xp33_ASAP7_75t_L g322 ( 
.A(n_316),
.B(n_317),
.Y(n_322)
);

NOR2xp33_ASAP7_75t_L g323 ( 
.A(n_318),
.B(n_307),
.Y(n_323)
);

OAI21xp5_ASAP7_75t_SL g320 ( 
.A1(n_301),
.A2(n_286),
.B(n_285),
.Y(n_320)
);

INVxp67_ASAP7_75t_L g321 ( 
.A(n_315),
.Y(n_321)
);

NAND2xp5_ASAP7_75t_L g329 ( 
.A(n_321),
.B(n_323),
.Y(n_329)
);

INVxp67_ASAP7_75t_L g325 ( 
.A(n_319),
.Y(n_325)
);

NAND2xp5_ASAP7_75t_L g330 ( 
.A(n_325),
.B(n_326),
.Y(n_330)
);

AOI22xp5_ASAP7_75t_L g326 ( 
.A1(n_313),
.A2(n_301),
.B1(n_304),
.B2(n_299),
.Y(n_326)
);

XNOR2xp5_ASAP7_75t_L g328 ( 
.A(n_327),
.B(n_314),
.Y(n_328)
);

OAI21xp33_ASAP7_75t_L g333 ( 
.A1(n_328),
.A2(n_331),
.B(n_311),
.Y(n_333)
);

NAND2xp5_ASAP7_75t_L g331 ( 
.A(n_322),
.B(n_317),
.Y(n_331)
);

OAI21xp5_ASAP7_75t_SL g332 ( 
.A1(n_329),
.A2(n_321),
.B(n_324),
.Y(n_332)
);

AOI21xp5_ASAP7_75t_SL g334 ( 
.A1(n_332),
.A2(n_333),
.B(n_330),
.Y(n_334)
);

XOR2xp5_ASAP7_75t_L g335 ( 
.A(n_334),
.B(n_328),
.Y(n_335)
);

AOI22xp5_ASAP7_75t_L g336 ( 
.A1(n_335),
.A2(n_312),
.B1(n_303),
.B2(n_290),
.Y(n_336)
);

INVxp67_ASAP7_75t_L g337 ( 
.A(n_336),
.Y(n_337)
);


endmodule