module fake_aes_8373_n_25 (n_11, n_1, n_2, n_12, n_6, n_4, n_3, n_9, n_5, n_7, n_10, n_8, n_0, n_25);
input n_11;
input n_1;
input n_2;
input n_12;
input n_6;
input n_4;
input n_3;
input n_9;
input n_5;
input n_7;
input n_10;
input n_8;
input n_0;
output n_25;
wire n_20;
wire n_23;
wire n_22;
wire n_16;
wire n_13;
wire n_18;
wire n_17;
wire n_14;
wire n_15;
wire n_24;
wire n_19;
wire n_21;
CKINVDCx5p33_ASAP7_75t_R g13 ( .A(n_6), .Y(n_13) );
INVx1_ASAP7_75t_L g14 ( .A(n_2), .Y(n_14) );
CKINVDCx5p33_ASAP7_75t_R g15 ( .A(n_3), .Y(n_15) );
CKINVDCx5p33_ASAP7_75t_R g16 ( .A(n_0), .Y(n_16) );
AOI21xp5_ASAP7_75t_L g17 ( .A1(n_14), .A2(n_8), .B(n_11), .Y(n_17) );
AOI21xp5_ASAP7_75t_L g18 ( .A1(n_14), .A2(n_7), .B(n_10), .Y(n_18) );
INVx1_ASAP7_75t_L g19 ( .A(n_17), .Y(n_19) );
OA21x2_ASAP7_75t_L g20 ( .A1(n_19), .A2(n_18), .B(n_15), .Y(n_20) );
AOI22xp5_ASAP7_75t_L g21 ( .A1(n_20), .A2(n_16), .B1(n_13), .B2(n_0), .Y(n_21) );
AND3x4_ASAP7_75t_L g22 ( .A(n_21), .B(n_1), .C(n_4), .Y(n_22) );
AND2x2_ASAP7_75t_L g23 ( .A(n_22), .B(n_1), .Y(n_23) );
CKINVDCx20_ASAP7_75t_R g24 ( .A(n_23), .Y(n_24) );
AOI22xp5_ASAP7_75t_L g25 ( .A1(n_24), .A2(n_5), .B1(n_9), .B2(n_12), .Y(n_25) );
endmodule