module fake_jpeg_12945_n_337 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_337);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_337;

wire n_253;
wire n_330;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_256;
wire n_221;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_13),
.Y(n_16)
);

BUFx12f_ASAP7_75t_L g17 ( 
.A(n_14),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_13),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_0),
.Y(n_19)
);

BUFx12f_ASAP7_75t_L g20 ( 
.A(n_3),
.Y(n_20)
);

BUFx12f_ASAP7_75t_L g21 ( 
.A(n_11),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_15),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_8),
.Y(n_23)
);

INVx4_ASAP7_75t_L g24 ( 
.A(n_15),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_6),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_12),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_9),
.Y(n_27)
);

BUFx12f_ASAP7_75t_L g28 ( 
.A(n_2),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_10),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_8),
.Y(n_30)
);

INVx2_ASAP7_75t_L g31 ( 
.A(n_13),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_4),
.Y(n_32)
);

HB1xp67_ASAP7_75t_L g33 ( 
.A(n_15),
.Y(n_33)
);

INVxp67_ASAP7_75t_L g34 ( 
.A(n_6),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_5),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g36 ( 
.A(n_16),
.B(n_0),
.Y(n_36)
);

NAND2xp5_ASAP7_75t_SL g74 ( 
.A(n_36),
.B(n_38),
.Y(n_74)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_28),
.Y(n_37)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_37),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g38 ( 
.A(n_16),
.B(n_0),
.Y(n_38)
);

BUFx8_ASAP7_75t_L g39 ( 
.A(n_28),
.Y(n_39)
);

INVx3_ASAP7_75t_L g59 ( 
.A(n_39),
.Y(n_59)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_33),
.Y(n_40)
);

NAND2xp5_ASAP7_75t_L g75 ( 
.A(n_40),
.B(n_46),
.Y(n_75)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_23),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_41),
.Y(n_65)
);

INVx8_ASAP7_75t_L g42 ( 
.A(n_23),
.Y(n_42)
);

INVx3_ASAP7_75t_L g61 ( 
.A(n_42),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g43 ( 
.A(n_18),
.B(n_14),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_43),
.B(n_47),
.Y(n_60)
);

INVx2_ASAP7_75t_L g44 ( 
.A(n_28),
.Y(n_44)
);

INVx2_ASAP7_75t_L g49 ( 
.A(n_44),
.Y(n_49)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_28),
.Y(n_45)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_45),
.Y(n_50)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_33),
.Y(n_46)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_18),
.Y(n_47)
);

CKINVDCx16_ASAP7_75t_R g51 ( 
.A(n_39),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_51),
.B(n_52),
.Y(n_79)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_37),
.Y(n_52)
);

AOI22xp33_ASAP7_75t_SL g53 ( 
.A1(n_40),
.A2(n_24),
.B1(n_34),
.B2(n_32),
.Y(n_53)
);

AOI22xp33_ASAP7_75t_SL g100 ( 
.A1(n_53),
.A2(n_57),
.B1(n_17),
.B2(n_21),
.Y(n_100)
);

INVx11_ASAP7_75t_L g54 ( 
.A(n_39),
.Y(n_54)
);

BUFx12f_ASAP7_75t_L g86 ( 
.A(n_54),
.Y(n_86)
);

INVx2_ASAP7_75t_L g55 ( 
.A(n_44),
.Y(n_55)
);

INVx2_ASAP7_75t_L g81 ( 
.A(n_55),
.Y(n_81)
);

NAND2xp67_ASAP7_75t_SL g56 ( 
.A(n_36),
.B(n_24),
.Y(n_56)
);

OAI21xp33_ASAP7_75t_L g98 ( 
.A1(n_56),
.A2(n_29),
.B(n_35),
.Y(n_98)
);

AOI22xp33_ASAP7_75t_SL g57 ( 
.A1(n_40),
.A2(n_24),
.B1(n_32),
.B2(n_23),
.Y(n_57)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_44),
.Y(n_58)
);

INVx2_ASAP7_75t_L g108 ( 
.A(n_58),
.Y(n_108)
);

INVx4_ASAP7_75t_L g62 ( 
.A(n_42),
.Y(n_62)
);

INVx4_ASAP7_75t_L g76 ( 
.A(n_62),
.Y(n_76)
);

INVx2_ASAP7_75t_L g63 ( 
.A(n_37),
.Y(n_63)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_63),
.Y(n_78)
);

INVx2_ASAP7_75t_L g64 ( 
.A(n_45),
.Y(n_64)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_64),
.Y(n_88)
);

INVx4_ASAP7_75t_L g66 ( 
.A(n_42),
.Y(n_66)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_66),
.Y(n_93)
);

AOI22xp33_ASAP7_75t_L g67 ( 
.A1(n_46),
.A2(n_31),
.B1(n_26),
.B2(n_35),
.Y(n_67)
);

OAI22xp33_ASAP7_75t_L g103 ( 
.A1(n_67),
.A2(n_25),
.B1(n_30),
.B2(n_27),
.Y(n_103)
);

INVx2_ASAP7_75t_L g68 ( 
.A(n_45),
.Y(n_68)
);

BUFx3_ASAP7_75t_L g104 ( 
.A(n_68),
.Y(n_104)
);

INVx2_ASAP7_75t_L g69 ( 
.A(n_41),
.Y(n_69)
);

AND2x2_ASAP7_75t_L g95 ( 
.A(n_69),
.B(n_70),
.Y(n_95)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_41),
.Y(n_70)
);

INVx3_ASAP7_75t_L g71 ( 
.A(n_39),
.Y(n_71)
);

INVx6_ASAP7_75t_L g83 ( 
.A(n_71),
.Y(n_83)
);

INVx2_ASAP7_75t_L g72 ( 
.A(n_41),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_72),
.B(n_73),
.Y(n_82)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_36),
.Y(n_73)
);

CKINVDCx20_ASAP7_75t_R g77 ( 
.A(n_75),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_77),
.B(n_80),
.Y(n_117)
);

CKINVDCx20_ASAP7_75t_R g80 ( 
.A(n_54),
.Y(n_80)
);

AOI22xp5_ASAP7_75t_SL g84 ( 
.A1(n_56),
.A2(n_46),
.B1(n_22),
.B2(n_31),
.Y(n_84)
);

OAI21xp5_ASAP7_75t_SL g121 ( 
.A1(n_84),
.A2(n_91),
.B(n_97),
.Y(n_121)
);

INVxp67_ASAP7_75t_L g85 ( 
.A(n_48),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g127 ( 
.A(n_85),
.B(n_94),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_L g87 ( 
.A(n_74),
.B(n_38),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_L g114 ( 
.A(n_87),
.B(n_92),
.Y(n_114)
);

AOI22xp5_ASAP7_75t_L g89 ( 
.A1(n_69),
.A2(n_41),
.B1(n_42),
.B2(n_70),
.Y(n_89)
);

OAI22xp5_ASAP7_75t_L g125 ( 
.A1(n_89),
.A2(n_101),
.B1(n_102),
.B2(n_105),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_SL g90 ( 
.A(n_60),
.B(n_38),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_SL g116 ( 
.A(n_90),
.B(n_99),
.Y(n_116)
);

OR2x2_ASAP7_75t_L g91 ( 
.A(n_59),
.B(n_19),
.Y(n_91)
);

AO22x1_ASAP7_75t_SL g92 ( 
.A1(n_68),
.A2(n_39),
.B1(n_27),
.B2(n_19),
.Y(n_92)
);

CKINVDCx20_ASAP7_75t_R g94 ( 
.A(n_50),
.Y(n_94)
);

AO22x2_ASAP7_75t_SL g96 ( 
.A1(n_49),
.A2(n_39),
.B1(n_47),
.B2(n_43),
.Y(n_96)
);

AOI22xp33_ASAP7_75t_L g119 ( 
.A1(n_96),
.A2(n_61),
.B1(n_66),
.B2(n_28),
.Y(n_119)
);

NOR2xp67_ASAP7_75t_L g97 ( 
.A(n_49),
.B(n_47),
.Y(n_97)
);

AND2x2_ASAP7_75t_L g128 ( 
.A(n_98),
.B(n_103),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_55),
.B(n_29),
.Y(n_99)
);

INVxp67_ASAP7_75t_L g111 ( 
.A(n_100),
.Y(n_111)
);

OAI22xp5_ASAP7_75t_L g101 ( 
.A1(n_72),
.A2(n_26),
.B1(n_30),
.B2(n_32),
.Y(n_101)
);

OAI22xp5_ASAP7_75t_L g102 ( 
.A1(n_65),
.A2(n_26),
.B1(n_30),
.B2(n_22),
.Y(n_102)
);

OAI22xp5_ASAP7_75t_L g105 ( 
.A1(n_65),
.A2(n_25),
.B1(n_17),
.B2(n_21),
.Y(n_105)
);

CKINVDCx16_ASAP7_75t_R g106 ( 
.A(n_59),
.Y(n_106)
);

INVxp67_ASAP7_75t_L g120 ( 
.A(n_106),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_58),
.B(n_17),
.Y(n_107)
);

INVxp67_ASAP7_75t_L g124 ( 
.A(n_107),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_71),
.B(n_17),
.Y(n_109)
);

CKINVDCx20_ASAP7_75t_R g129 ( 
.A(n_109),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_L g110 ( 
.A(n_62),
.B(n_0),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_L g136 ( 
.A(n_110),
.B(n_1),
.Y(n_136)
);

BUFx2_ASAP7_75t_L g112 ( 
.A(n_76),
.Y(n_112)
);

INVx2_ASAP7_75t_L g150 ( 
.A(n_112),
.Y(n_150)
);

BUFx2_ASAP7_75t_L g113 ( 
.A(n_76),
.Y(n_113)
);

INVx2_ASAP7_75t_L g161 ( 
.A(n_113),
.Y(n_161)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_95),
.Y(n_115)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_115),
.Y(n_144)
);

INVx3_ASAP7_75t_L g118 ( 
.A(n_83),
.Y(n_118)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_118),
.Y(n_157)
);

OAI22xp5_ASAP7_75t_L g149 ( 
.A1(n_119),
.A2(n_80),
.B1(n_91),
.B2(n_89),
.Y(n_149)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_95),
.Y(n_122)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_122),
.Y(n_158)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_95),
.Y(n_123)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_123),
.Y(n_168)
);

INVx2_ASAP7_75t_L g126 ( 
.A(n_81),
.Y(n_126)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_126),
.Y(n_174)
);

MAJIxp5_ASAP7_75t_L g130 ( 
.A(n_77),
.B(n_61),
.C(n_21),
.Y(n_130)
);

MAJIxp5_ASAP7_75t_L g147 ( 
.A(n_130),
.B(n_137),
.C(n_91),
.Y(n_147)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_78),
.Y(n_131)
);

INVxp67_ASAP7_75t_L g152 ( 
.A(n_131),
.Y(n_152)
);

INVx3_ASAP7_75t_L g132 ( 
.A(n_83),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_L g141 ( 
.A(n_132),
.B(n_133),
.Y(n_141)
);

INVx2_ASAP7_75t_L g133 ( 
.A(n_81),
.Y(n_133)
);

AOI21xp5_ASAP7_75t_SL g134 ( 
.A1(n_96),
.A2(n_1),
.B(n_2),
.Y(n_134)
);

INVxp67_ASAP7_75t_L g169 ( 
.A(n_134),
.Y(n_169)
);

OAI22xp5_ASAP7_75t_L g135 ( 
.A1(n_96),
.A2(n_21),
.B1(n_20),
.B2(n_14),
.Y(n_135)
);

AOI22xp5_ASAP7_75t_L g142 ( 
.A1(n_135),
.A2(n_140),
.B1(n_105),
.B2(n_102),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_SL g145 ( 
.A(n_136),
.B(n_139),
.Y(n_145)
);

MAJIxp5_ASAP7_75t_L g137 ( 
.A(n_87),
.B(n_82),
.C(n_90),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_L g138 ( 
.A(n_94),
.B(n_1),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_L g160 ( 
.A(n_138),
.B(n_1),
.Y(n_160)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_78),
.Y(n_139)
);

OAI22xp33_ASAP7_75t_SL g140 ( 
.A1(n_96),
.A2(n_20),
.B1(n_12),
.B2(n_11),
.Y(n_140)
);

OA22x2_ASAP7_75t_L g200 ( 
.A1(n_142),
.A2(n_158),
.B1(n_144),
.B2(n_168),
.Y(n_200)
);

NOR2xp33_ASAP7_75t_L g143 ( 
.A(n_129),
.B(n_79),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_SL g177 ( 
.A(n_143),
.B(n_154),
.Y(n_177)
);

NOR2xp33_ASAP7_75t_SL g146 ( 
.A(n_116),
.B(n_84),
.Y(n_146)
);

OR2x2_ASAP7_75t_L g184 ( 
.A(n_146),
.B(n_159),
.Y(n_184)
);

XNOR2x1_ASAP7_75t_L g202 ( 
.A(n_147),
.B(n_148),
.Y(n_202)
);

XNOR2xp5_ASAP7_75t_L g148 ( 
.A(n_137),
.B(n_110),
.Y(n_148)
);

AND2x2_ASAP7_75t_L g188 ( 
.A(n_149),
.B(n_118),
.Y(n_188)
);

XNOR2xp5_ASAP7_75t_L g151 ( 
.A(n_114),
.B(n_130),
.Y(n_151)
);

MAJIxp5_ASAP7_75t_L g206 ( 
.A(n_151),
.B(n_162),
.C(n_167),
.Y(n_206)
);

AOI21xp5_ASAP7_75t_L g153 ( 
.A1(n_114),
.A2(n_97),
.B(n_85),
.Y(n_153)
);

AOI21xp5_ASAP7_75t_L g203 ( 
.A1(n_153),
.A2(n_86),
.B(n_20),
.Y(n_203)
);

NOR2xp33_ASAP7_75t_L g154 ( 
.A(n_129),
.B(n_88),
.Y(n_154)
);

NOR2xp33_ASAP7_75t_L g155 ( 
.A(n_117),
.B(n_88),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_SL g181 ( 
.A(n_155),
.B(n_163),
.Y(n_181)
);

AOI22xp5_ASAP7_75t_L g156 ( 
.A1(n_125),
.A2(n_101),
.B1(n_92),
.B2(n_104),
.Y(n_156)
);

OAI22xp5_ASAP7_75t_SL g175 ( 
.A1(n_156),
.A2(n_134),
.B1(n_122),
.B2(n_123),
.Y(n_175)
);

CKINVDCx14_ASAP7_75t_R g159 ( 
.A(n_127),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_L g186 ( 
.A(n_160),
.B(n_164),
.Y(n_186)
);

XOR2xp5_ASAP7_75t_L g162 ( 
.A(n_136),
.B(n_93),
.Y(n_162)
);

NOR2xp33_ASAP7_75t_L g163 ( 
.A(n_124),
.B(n_104),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_L g164 ( 
.A(n_138),
.B(n_121),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_SL g165 ( 
.A(n_124),
.B(n_108),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_SL g190 ( 
.A(n_165),
.B(n_173),
.Y(n_190)
);

OAI22xp5_ASAP7_75t_L g166 ( 
.A1(n_111),
.A2(n_92),
.B1(n_108),
.B2(n_93),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_L g191 ( 
.A(n_166),
.B(n_170),
.Y(n_191)
);

MAJIxp5_ASAP7_75t_L g167 ( 
.A(n_115),
.B(n_92),
.C(n_106),
.Y(n_167)
);

OAI22xp5_ASAP7_75t_L g170 ( 
.A1(n_111),
.A2(n_83),
.B1(n_20),
.B2(n_86),
.Y(n_170)
);

CKINVDCx20_ASAP7_75t_R g171 ( 
.A(n_126),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_L g196 ( 
.A(n_171),
.B(n_172),
.Y(n_196)
);

CKINVDCx20_ASAP7_75t_R g172 ( 
.A(n_133),
.Y(n_172)
);

CKINVDCx16_ASAP7_75t_R g173 ( 
.A(n_128),
.Y(n_173)
);

AOI22xp5_ASAP7_75t_L g218 ( 
.A1(n_175),
.A2(n_180),
.B1(n_188),
.B2(n_192),
.Y(n_218)
);

XOR2xp5_ASAP7_75t_L g176 ( 
.A(n_151),
.B(n_121),
.Y(n_176)
);

MAJIxp5_ASAP7_75t_L g236 ( 
.A(n_176),
.B(n_193),
.C(n_5),
.Y(n_236)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_174),
.Y(n_178)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_178),
.Y(n_211)
);

AOI22xp33_ASAP7_75t_L g179 ( 
.A1(n_173),
.A2(n_128),
.B1(n_131),
.B2(n_139),
.Y(n_179)
);

INVxp67_ASAP7_75t_SL g212 ( 
.A(n_179),
.Y(n_212)
);

OAI22xp5_ASAP7_75t_SL g180 ( 
.A1(n_156),
.A2(n_128),
.B1(n_120),
.B2(n_132),
.Y(n_180)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_174),
.Y(n_182)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_182),
.Y(n_215)
);

CKINVDCx20_ASAP7_75t_R g183 ( 
.A(n_141),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_SL g209 ( 
.A(n_183),
.B(n_187),
.Y(n_209)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_157),
.Y(n_185)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_185),
.Y(n_216)
);

CKINVDCx20_ASAP7_75t_R g187 ( 
.A(n_171),
.Y(n_187)
);

INVxp67_ASAP7_75t_L g189 ( 
.A(n_167),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_L g213 ( 
.A(n_189),
.B(n_197),
.Y(n_213)
);

OAI22xp5_ASAP7_75t_SL g192 ( 
.A1(n_142),
.A2(n_120),
.B1(n_113),
.B2(n_112),
.Y(n_192)
);

XNOR2xp5_ASAP7_75t_L g193 ( 
.A(n_148),
.B(n_113),
.Y(n_193)
);

OAI21xp5_ASAP7_75t_L g194 ( 
.A1(n_169),
.A2(n_112),
.B(n_86),
.Y(n_194)
);

OAI21xp5_ASAP7_75t_L g222 ( 
.A1(n_194),
.A2(n_205),
.B(n_161),
.Y(n_222)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_157),
.Y(n_195)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_195),
.Y(n_231)
);

CKINVDCx20_ASAP7_75t_R g197 ( 
.A(n_172),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_SL g198 ( 
.A(n_145),
.B(n_12),
.Y(n_198)
);

NOR2xp33_ASAP7_75t_SL g219 ( 
.A(n_198),
.B(n_160),
.Y(n_219)
);

CKINVDCx20_ASAP7_75t_R g199 ( 
.A(n_166),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_L g225 ( 
.A(n_199),
.B(n_200),
.Y(n_225)
);

AOI22xp33_ASAP7_75t_L g201 ( 
.A1(n_169),
.A2(n_86),
.B1(n_11),
.B2(n_10),
.Y(n_201)
);

OAI22xp33_ASAP7_75t_L g220 ( 
.A1(n_201),
.A2(n_161),
.B1(n_150),
.B2(n_149),
.Y(n_220)
);

OAI21xp5_ASAP7_75t_SL g214 ( 
.A1(n_203),
.A2(n_158),
.B(n_168),
.Y(n_214)
);

OAI22xp5_ASAP7_75t_SL g204 ( 
.A1(n_153),
.A2(n_10),
.B1(n_3),
.B2(n_4),
.Y(n_204)
);

AOI22xp5_ASAP7_75t_L g232 ( 
.A1(n_204),
.A2(n_175),
.B1(n_205),
.B2(n_192),
.Y(n_232)
);

OAI21xp5_ASAP7_75t_L g205 ( 
.A1(n_164),
.A2(n_2),
.B(n_3),
.Y(n_205)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_152),
.Y(n_207)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_207),
.Y(n_210)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_152),
.Y(n_208)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_208),
.Y(n_221)
);

OAI21xp5_ASAP7_75t_SL g253 ( 
.A1(n_214),
.A2(n_223),
.B(n_226),
.Y(n_253)
);

A2O1A1Ixp33_ASAP7_75t_L g217 ( 
.A1(n_184),
.A2(n_147),
.B(n_144),
.C(n_146),
.Y(n_217)
);

NAND2xp5_ASAP7_75t_L g238 ( 
.A(n_217),
.B(n_222),
.Y(n_238)
);

NAND2xp5_ASAP7_75t_SL g244 ( 
.A(n_219),
.B(n_227),
.Y(n_244)
);

OAI22xp5_ASAP7_75t_L g243 ( 
.A1(n_220),
.A2(n_232),
.B1(n_199),
.B2(n_191),
.Y(n_243)
);

A2O1A1Ixp33_ASAP7_75t_SL g223 ( 
.A1(n_203),
.A2(n_170),
.B(n_150),
.C(n_162),
.Y(n_223)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_196),
.Y(n_224)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_224),
.Y(n_239)
);

OAI21xp5_ASAP7_75t_L g226 ( 
.A1(n_184),
.A2(n_189),
.B(n_190),
.Y(n_226)
);

OAI21xp5_ASAP7_75t_SL g227 ( 
.A1(n_188),
.A2(n_2),
.B(n_3),
.Y(n_227)
);

XNOR2xp5_ASAP7_75t_L g228 ( 
.A(n_206),
.B(n_4),
.Y(n_228)
);

MAJIxp5_ASAP7_75t_L g257 ( 
.A(n_228),
.B(n_233),
.C(n_236),
.Y(n_257)
);

NAND2xp5_ASAP7_75t_SL g229 ( 
.A(n_177),
.B(n_4),
.Y(n_229)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_229),
.Y(n_241)
);

OAI21xp5_ASAP7_75t_SL g230 ( 
.A1(n_188),
.A2(n_5),
.B(n_6),
.Y(n_230)
);

XNOR2xp5_ASAP7_75t_L g245 ( 
.A(n_230),
.B(n_204),
.Y(n_245)
);

XNOR2xp5_ASAP7_75t_L g233 ( 
.A(n_206),
.B(n_202),
.Y(n_233)
);

CKINVDCx20_ASAP7_75t_R g234 ( 
.A(n_196),
.Y(n_234)
);

CKINVDCx20_ASAP7_75t_R g252 ( 
.A(n_234),
.Y(n_252)
);

AOI21xp5_ASAP7_75t_L g235 ( 
.A1(n_194),
.A2(n_5),
.B(n_6),
.Y(n_235)
);

OAI22xp5_ASAP7_75t_SL g237 ( 
.A1(n_235),
.A2(n_197),
.B1(n_207),
.B2(n_208),
.Y(n_237)
);

AOI22xp5_ASAP7_75t_L g263 ( 
.A1(n_237),
.A2(n_243),
.B1(n_256),
.B2(n_258),
.Y(n_263)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_216),
.Y(n_240)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_240),
.Y(n_268)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_231),
.Y(n_242)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_242),
.Y(n_272)
);

XNOR2xp5_ASAP7_75t_L g267 ( 
.A(n_245),
.B(n_260),
.Y(n_267)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_209),
.Y(n_246)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_246),
.Y(n_275)
);

AOI22xp5_ASAP7_75t_L g247 ( 
.A1(n_224),
.A2(n_180),
.B1(n_191),
.B2(n_176),
.Y(n_247)
);

OAI22xp5_ASAP7_75t_SL g261 ( 
.A1(n_247),
.A2(n_249),
.B1(n_218),
.B2(n_212),
.Y(n_261)
);

OAI22xp5_ASAP7_75t_L g248 ( 
.A1(n_232),
.A2(n_181),
.B1(n_186),
.B2(n_200),
.Y(n_248)
);

CKINVDCx16_ASAP7_75t_R g270 ( 
.A(n_248),
.Y(n_270)
);

AOI22xp5_ASAP7_75t_L g249 ( 
.A1(n_225),
.A2(n_200),
.B1(n_186),
.B2(n_195),
.Y(n_249)
);

XNOR2xp5_ASAP7_75t_L g250 ( 
.A(n_233),
.B(n_202),
.Y(n_250)
);

MAJIxp5_ASAP7_75t_L g269 ( 
.A(n_250),
.B(n_251),
.C(n_254),
.Y(n_269)
);

XOR2xp5_ASAP7_75t_L g251 ( 
.A(n_226),
.B(n_193),
.Y(n_251)
);

XNOR2xp5_ASAP7_75t_L g254 ( 
.A(n_213),
.B(n_236),
.Y(n_254)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_210),
.Y(n_255)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_255),
.Y(n_279)
);

OAI22xp5_ASAP7_75t_SL g256 ( 
.A1(n_225),
.A2(n_200),
.B1(n_185),
.B2(n_178),
.Y(n_256)
);

OAI22xp5_ASAP7_75t_SL g258 ( 
.A1(n_218),
.A2(n_182),
.B1(n_8),
.B2(n_9),
.Y(n_258)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_210),
.Y(n_259)
);

NOR2xp33_ASAP7_75t_L g262 ( 
.A(n_259),
.B(n_221),
.Y(n_262)
);

MAJIxp5_ASAP7_75t_L g260 ( 
.A(n_213),
.B(n_7),
.C(n_8),
.Y(n_260)
);

NOR2xp33_ASAP7_75t_L g286 ( 
.A(n_261),
.B(n_274),
.Y(n_286)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_262),
.Y(n_282)
);

CKINVDCx20_ASAP7_75t_R g264 ( 
.A(n_252),
.Y(n_264)
);

NAND2xp5_ASAP7_75t_SL g281 ( 
.A(n_264),
.B(n_273),
.Y(n_281)
);

AOI22xp5_ASAP7_75t_L g265 ( 
.A1(n_256),
.A2(n_220),
.B1(n_222),
.B2(n_221),
.Y(n_265)
);

OAI22xp5_ASAP7_75t_L g283 ( 
.A1(n_265),
.A2(n_280),
.B1(n_247),
.B2(n_223),
.Y(n_283)
);

INVx1_ASAP7_75t_SL g266 ( 
.A(n_240),
.Y(n_266)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_266),
.Y(n_285)
);

OAI22xp5_ASAP7_75t_SL g271 ( 
.A1(n_249),
.A2(n_217),
.B1(n_223),
.B2(n_235),
.Y(n_271)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_271),
.Y(n_288)
);

NOR2xp33_ASAP7_75t_L g273 ( 
.A(n_254),
.B(n_228),
.Y(n_273)
);

FAx1_ASAP7_75t_SL g274 ( 
.A(n_238),
.B(n_214),
.CI(n_223),
.CON(n_274),
.SN(n_274)
);

CKINVDCx20_ASAP7_75t_R g276 ( 
.A(n_237),
.Y(n_276)
);

NOR2xp33_ASAP7_75t_L g289 ( 
.A(n_276),
.B(n_277),
.Y(n_289)
);

NOR2xp33_ASAP7_75t_L g277 ( 
.A(n_244),
.B(n_241),
.Y(n_277)
);

NAND2xp5_ASAP7_75t_L g278 ( 
.A(n_239),
.B(n_211),
.Y(n_278)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_278),
.Y(n_294)
);

AOI22xp5_ASAP7_75t_L g280 ( 
.A1(n_238),
.A2(n_223),
.B1(n_215),
.B2(n_227),
.Y(n_280)
);

AND2x2_ASAP7_75t_L g297 ( 
.A(n_283),
.B(n_261),
.Y(n_297)
);

OAI21xp5_ASAP7_75t_SL g284 ( 
.A1(n_280),
.A2(n_253),
.B(n_242),
.Y(n_284)
);

OR2x2_ASAP7_75t_L g301 ( 
.A(n_284),
.B(n_293),
.Y(n_301)
);

OAI21xp5_ASAP7_75t_L g287 ( 
.A1(n_271),
.A2(n_253),
.B(n_258),
.Y(n_287)
);

AOI21xp5_ASAP7_75t_SL g304 ( 
.A1(n_287),
.A2(n_284),
.B(n_288),
.Y(n_304)
);

AOI21xp5_ASAP7_75t_L g290 ( 
.A1(n_265),
.A2(n_251),
.B(n_250),
.Y(n_290)
);

AOI21xp5_ASAP7_75t_L g299 ( 
.A1(n_290),
.A2(n_263),
.B(n_270),
.Y(n_299)
);

MAJIxp5_ASAP7_75t_L g291 ( 
.A(n_269),
.B(n_257),
.C(n_260),
.Y(n_291)
);

NAND2xp5_ASAP7_75t_L g305 ( 
.A(n_291),
.B(n_295),
.Y(n_305)
);

XOR2xp5_ASAP7_75t_L g292 ( 
.A(n_269),
.B(n_257),
.Y(n_292)
);

MAJIxp5_ASAP7_75t_L g306 ( 
.A(n_292),
.B(n_263),
.C(n_278),
.Y(n_306)
);

OAI21xp5_ASAP7_75t_SL g293 ( 
.A1(n_274),
.A2(n_245),
.B(n_230),
.Y(n_293)
);

MAJIxp5_ASAP7_75t_L g295 ( 
.A(n_267),
.B(n_7),
.C(n_9),
.Y(n_295)
);

MAJIxp5_ASAP7_75t_L g296 ( 
.A(n_267),
.B(n_7),
.C(n_9),
.Y(n_296)
);

NAND2xp5_ASAP7_75t_L g309 ( 
.A(n_296),
.B(n_275),
.Y(n_309)
);

AOI22xp5_ASAP7_75t_SL g314 ( 
.A1(n_297),
.A2(n_288),
.B1(n_287),
.B2(n_274),
.Y(n_314)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_281),
.Y(n_298)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_298),
.Y(n_313)
);

AOI21x1_ASAP7_75t_L g318 ( 
.A1(n_299),
.A2(n_268),
.B(n_272),
.Y(n_318)
);

NOR2xp33_ASAP7_75t_L g300 ( 
.A(n_282),
.B(n_275),
.Y(n_300)
);

AOI21xp5_ASAP7_75t_L g311 ( 
.A1(n_300),
.A2(n_294),
.B(n_279),
.Y(n_311)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_285),
.Y(n_302)
);

NOR2xp33_ASAP7_75t_L g315 ( 
.A(n_302),
.B(n_303),
.Y(n_315)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_285),
.Y(n_303)
);

OAI22xp5_ASAP7_75t_SL g317 ( 
.A1(n_304),
.A2(n_290),
.B1(n_293),
.B2(n_272),
.Y(n_317)
);

MAJIxp5_ASAP7_75t_L g319 ( 
.A(n_306),
.B(n_291),
.C(n_292),
.Y(n_319)
);

AND2x2_ASAP7_75t_L g307 ( 
.A(n_289),
.B(n_266),
.Y(n_307)
);

AND2x2_ASAP7_75t_L g312 ( 
.A(n_307),
.B(n_300),
.Y(n_312)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_294),
.Y(n_308)
);

NOR2xp33_ASAP7_75t_SL g310 ( 
.A(n_308),
.B(n_309),
.Y(n_310)
);

AOI21x1_ASAP7_75t_L g325 ( 
.A1(n_311),
.A2(n_295),
.B(n_296),
.Y(n_325)
);

NAND2xp5_ASAP7_75t_L g320 ( 
.A(n_312),
.B(n_314),
.Y(n_320)
);

AOI22xp5_ASAP7_75t_L g316 ( 
.A1(n_297),
.A2(n_307),
.B1(n_286),
.B2(n_301),
.Y(n_316)
);

NAND2xp5_ASAP7_75t_L g321 ( 
.A(n_316),
.B(n_317),
.Y(n_321)
);

MAJIxp5_ASAP7_75t_L g324 ( 
.A(n_318),
.B(n_319),
.C(n_301),
.Y(n_324)
);

NOR2xp33_ASAP7_75t_L g322 ( 
.A(n_310),
.B(n_279),
.Y(n_322)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_322),
.Y(n_329)
);

NOR2xp33_ASAP7_75t_SL g323 ( 
.A(n_313),
.B(n_305),
.Y(n_323)
);

NOR2xp33_ASAP7_75t_SL g328 ( 
.A(n_323),
.B(n_326),
.Y(n_328)
);

NAND2xp5_ASAP7_75t_L g330 ( 
.A(n_324),
.B(n_325),
.Y(n_330)
);

AOI21xp5_ASAP7_75t_L g326 ( 
.A1(n_312),
.A2(n_268),
.B(n_7),
.Y(n_326)
);

NOR2xp33_ASAP7_75t_L g327 ( 
.A(n_322),
.B(n_316),
.Y(n_327)
);

INVxp67_ASAP7_75t_L g332 ( 
.A(n_327),
.Y(n_332)
);

NAND2xp33_ASAP7_75t_R g331 ( 
.A(n_330),
.B(n_329),
.Y(n_331)
);

O2A1O1Ixp33_ASAP7_75t_SL g333 ( 
.A1(n_331),
.A2(n_332),
.B(n_321),
.C(n_320),
.Y(n_333)
);

AOI21xp5_ASAP7_75t_L g334 ( 
.A1(n_333),
.A2(n_319),
.B(n_315),
.Y(n_334)
);

BUFx24_ASAP7_75t_SL g335 ( 
.A(n_334),
.Y(n_335)
);

MAJIxp5_ASAP7_75t_L g336 ( 
.A(n_335),
.B(n_314),
.C(n_317),
.Y(n_336)
);

NOR2xp33_ASAP7_75t_SL g337 ( 
.A(n_336),
.B(n_328),
.Y(n_337)
);


endmodule