module fake_jpeg_2893_n_148 (n_13, n_21, n_33, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_19, n_18, n_20, n_35, n_4, n_34, n_30, n_16, n_3, n_0, n_24, n_28, n_38, n_26, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_12, n_32, n_8, n_15, n_7, n_148);

input n_13;
input n_21;
input n_33;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_35;
input n_4;
input n_34;
input n_30;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_148;

wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_147;
wire n_73;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_49;
wire n_76;
wire n_127;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_103;
wire n_50;
wire n_124;
wire n_141;
wire n_57;
wire n_119;
wire n_69;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_106;
wire n_111;
wire n_44;
wire n_143;
wire n_75;
wire n_122;
wire n_121;
wire n_99;
wire n_102;
wire n_130;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_78;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_54;
wire n_91;
wire n_93;
wire n_138;
wire n_101;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_97;
wire n_135;
wire n_62;
wire n_120;
wire n_43;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

INVx1_ASAP7_75t_L g39 ( 
.A(n_33),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_16),
.Y(n_40)
);

BUFx12f_ASAP7_75t_L g41 ( 
.A(n_0),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_28),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_3),
.Y(n_43)
);

INVx8_ASAP7_75t_L g44 ( 
.A(n_30),
.Y(n_44)
);

BUFx3_ASAP7_75t_L g45 ( 
.A(n_20),
.Y(n_45)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_32),
.Y(n_46)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_13),
.Y(n_47)
);

BUFx3_ASAP7_75t_L g48 ( 
.A(n_7),
.Y(n_48)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_37),
.Y(n_49)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_29),
.Y(n_50)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_21),
.Y(n_51)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_26),
.Y(n_52)
);

BUFx16f_ASAP7_75t_L g53 ( 
.A(n_24),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_43),
.Y(n_54)
);

INVx2_ASAP7_75t_L g68 ( 
.A(n_54),
.Y(n_68)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_39),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_55),
.B(n_58),
.Y(n_61)
);

BUFx12f_ASAP7_75t_L g56 ( 
.A(n_53),
.Y(n_56)
);

INVx3_ASAP7_75t_L g65 ( 
.A(n_56),
.Y(n_65)
);

BUFx5_ASAP7_75t_L g57 ( 
.A(n_53),
.Y(n_57)
);

INVx3_ASAP7_75t_L g71 ( 
.A(n_57),
.Y(n_71)
);

BUFx3_ASAP7_75t_L g58 ( 
.A(n_53),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_SL g59 ( 
.A(n_47),
.B(n_0),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_59),
.B(n_60),
.Y(n_63)
);

INVx4_ASAP7_75t_L g60 ( 
.A(n_41),
.Y(n_60)
);

OAI22xp33_ASAP7_75t_L g62 ( 
.A1(n_54),
.A2(n_43),
.B1(n_40),
.B2(n_51),
.Y(n_62)
);

OAI22xp5_ASAP7_75t_SL g79 ( 
.A1(n_62),
.A2(n_67),
.B1(n_69),
.B2(n_56),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_SL g64 ( 
.A(n_59),
.B(n_40),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_SL g84 ( 
.A(n_64),
.B(n_49),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g66 ( 
.A(n_55),
.B(n_50),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_L g77 ( 
.A(n_66),
.B(n_70),
.Y(n_77)
);

AOI22xp33_ASAP7_75t_SL g67 ( 
.A1(n_60),
.A2(n_48),
.B1(n_41),
.B2(n_56),
.Y(n_67)
);

AOI22xp5_ASAP7_75t_L g69 ( 
.A1(n_54),
.A2(n_39),
.B1(n_50),
.B2(n_46),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_56),
.B(n_46),
.Y(n_70)
);

MAJIxp5_ASAP7_75t_L g72 ( 
.A(n_66),
.B(n_42),
.C(n_52),
.Y(n_72)
);

AND2x2_ASAP7_75t_L g88 ( 
.A(n_72),
.B(n_75),
.Y(n_88)
);

INVx5_ASAP7_75t_L g73 ( 
.A(n_65),
.Y(n_73)
);

BUFx2_ASAP7_75t_L g90 ( 
.A(n_73),
.Y(n_90)
);

INVx2_ASAP7_75t_SL g74 ( 
.A(n_65),
.Y(n_74)
);

INVx2_ASAP7_75t_L g95 ( 
.A(n_74),
.Y(n_95)
);

MAJIxp5_ASAP7_75t_L g75 ( 
.A(n_61),
.B(n_58),
.C(n_45),
.Y(n_75)
);

INVx4_ASAP7_75t_L g76 ( 
.A(n_71),
.Y(n_76)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_76),
.Y(n_89)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_61),
.Y(n_78)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_78),
.Y(n_93)
);

INVxp67_ASAP7_75t_L g94 ( 
.A(n_79),
.Y(n_94)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_70),
.Y(n_80)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_80),
.Y(n_100)
);

CKINVDCx20_ASAP7_75t_R g81 ( 
.A(n_64),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_SL g92 ( 
.A(n_81),
.B(n_82),
.Y(n_92)
);

XNOR2xp5_ASAP7_75t_L g82 ( 
.A(n_63),
.B(n_41),
.Y(n_82)
);

INVx3_ASAP7_75t_L g83 ( 
.A(n_71),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g98 ( 
.A(n_83),
.B(n_57),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_SL g97 ( 
.A(n_84),
.B(n_1),
.Y(n_97)
);

INVx5_ASAP7_75t_L g85 ( 
.A(n_68),
.Y(n_85)
);

CKINVDCx20_ASAP7_75t_R g96 ( 
.A(n_85),
.Y(n_96)
);

OR2x2_ASAP7_75t_L g86 ( 
.A(n_77),
.B(n_69),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_SL g103 ( 
.A(n_86),
.B(n_38),
.Y(n_103)
);

AOI22xp5_ASAP7_75t_L g87 ( 
.A1(n_75),
.A2(n_68),
.B1(n_63),
.B2(n_48),
.Y(n_87)
);

AOI22xp5_ASAP7_75t_L g112 ( 
.A1(n_87),
.A2(n_91),
.B1(n_27),
.B2(n_25),
.Y(n_112)
);

OAI22xp5_ASAP7_75t_L g91 ( 
.A1(n_85),
.A2(n_45),
.B1(n_44),
.B2(n_83),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_SL g111 ( 
.A(n_97),
.B(n_31),
.Y(n_111)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_98),
.Y(n_102)
);

AND2x2_ASAP7_75t_SL g99 ( 
.A(n_76),
.B(n_44),
.Y(n_99)
);

MAJIxp5_ASAP7_75t_L g101 ( 
.A(n_99),
.B(n_74),
.C(n_73),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_L g118 ( 
.A(n_101),
.B(n_103),
.Y(n_118)
);

AOI22xp5_ASAP7_75t_L g104 ( 
.A1(n_94),
.A2(n_36),
.B1(n_35),
.B2(n_34),
.Y(n_104)
);

OAI22xp5_ASAP7_75t_SL g119 ( 
.A1(n_104),
.A2(n_99),
.B1(n_96),
.B2(n_95),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_93),
.B(n_1),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_L g125 ( 
.A(n_105),
.B(n_106),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_L g106 ( 
.A(n_100),
.B(n_2),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_L g107 ( 
.A(n_86),
.B(n_2),
.Y(n_107)
);

AOI322xp5_ASAP7_75t_SL g128 ( 
.A1(n_107),
.A2(n_108),
.A3(n_109),
.B1(n_110),
.B2(n_111),
.C1(n_116),
.C2(n_7),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_SL g108 ( 
.A(n_92),
.B(n_3),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_L g109 ( 
.A(n_88),
.B(n_4),
.Y(n_109)
);

CKINVDCx20_ASAP7_75t_R g110 ( 
.A(n_90),
.Y(n_110)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_112),
.Y(n_117)
);

XNOR2xp5_ASAP7_75t_SL g113 ( 
.A(n_88),
.B(n_23),
.Y(n_113)
);

XOR2xp5_ASAP7_75t_L g122 ( 
.A(n_113),
.B(n_5),
.Y(n_122)
);

BUFx2_ASAP7_75t_L g114 ( 
.A(n_90),
.Y(n_114)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_114),
.Y(n_120)
);

OAI21xp33_ASAP7_75t_L g115 ( 
.A1(n_94),
.A2(n_22),
.B(n_19),
.Y(n_115)
);

OAI21xp5_ASAP7_75t_L g123 ( 
.A1(n_115),
.A2(n_17),
.B(n_15),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_L g116 ( 
.A(n_89),
.B(n_4),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_L g131 ( 
.A(n_119),
.B(n_126),
.Y(n_131)
);

MAJIxp5_ASAP7_75t_L g121 ( 
.A(n_113),
.B(n_87),
.C(n_99),
.Y(n_121)
);

MAJIxp5_ASAP7_75t_L g130 ( 
.A(n_121),
.B(n_122),
.C(n_124),
.Y(n_130)
);

INVxp67_ASAP7_75t_L g133 ( 
.A(n_123),
.Y(n_133)
);

MAJIxp5_ASAP7_75t_L g124 ( 
.A(n_102),
.B(n_18),
.C(n_6),
.Y(n_124)
);

CKINVDCx20_ASAP7_75t_R g126 ( 
.A(n_114),
.Y(n_126)
);

AOI21xp5_ASAP7_75t_L g127 ( 
.A1(n_115),
.A2(n_5),
.B(n_6),
.Y(n_127)
);

OAI21xp5_ASAP7_75t_L g129 ( 
.A1(n_127),
.A2(n_104),
.B(n_101),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_L g132 ( 
.A(n_128),
.B(n_123),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_SL g135 ( 
.A(n_129),
.B(n_132),
.Y(n_135)
);

CKINVDCx20_ASAP7_75t_R g134 ( 
.A(n_125),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_SL g137 ( 
.A(n_134),
.B(n_117),
.Y(n_137)
);

OAI21xp5_ASAP7_75t_L g136 ( 
.A1(n_133),
.A2(n_118),
.B(n_121),
.Y(n_136)
);

MAJIxp5_ASAP7_75t_L g140 ( 
.A(n_136),
.B(n_133),
.C(n_131),
.Y(n_140)
);

XNOR2xp5_ASAP7_75t_L g139 ( 
.A(n_137),
.B(n_138),
.Y(n_139)
);

OAI322xp33_ASAP7_75t_L g138 ( 
.A1(n_130),
.A2(n_122),
.A3(n_119),
.B1(n_120),
.B2(n_124),
.C1(n_12),
.C2(n_8),
.Y(n_138)
);

OAI21xp5_ASAP7_75t_L g141 ( 
.A1(n_140),
.A2(n_135),
.B(n_9),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_SL g142 ( 
.A(n_141),
.B(n_139),
.Y(n_142)
);

AOI21xp5_ASAP7_75t_L g143 ( 
.A1(n_142),
.A2(n_14),
.B(n_9),
.Y(n_143)
);

NOR2xp33_ASAP7_75t_L g144 ( 
.A(n_143),
.B(n_8),
.Y(n_144)
);

OAI21xp5_ASAP7_75t_SL g145 ( 
.A1(n_144),
.A2(n_14),
.B(n_11),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_SL g146 ( 
.A(n_145),
.B(n_10),
.Y(n_146)
);

OAI311xp33_ASAP7_75t_L g147 ( 
.A1(n_146),
.A2(n_10),
.A3(n_11),
.B1(n_12),
.C1(n_13),
.Y(n_147)
);

BUFx24_ASAP7_75t_SL g148 ( 
.A(n_147),
.Y(n_148)
);


endmodule