module fake_jpeg_10879_n_393 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_393);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_393;

wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_385;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_340;
wire n_381;
wire n_377;
wire n_291;
wire n_236;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_265;
wire n_192;
wire n_115;
wire n_270;
wire n_387;
wire n_256;
wire n_221;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_370;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_39;
wire n_371;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_382;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_352;
wire n_350;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_389;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_384;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_360;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_378;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_379;
wire n_114;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_356;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_375;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_391;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

BUFx12f_ASAP7_75t_L g16 ( 
.A(n_9),
.Y(n_16)
);

CKINVDCx16_ASAP7_75t_R g17 ( 
.A(n_1),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_14),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_5),
.Y(n_19)
);

INVx3_ASAP7_75t_L g20 ( 
.A(n_2),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_5),
.Y(n_21)
);

INVx11_ASAP7_75t_L g22 ( 
.A(n_14),
.Y(n_22)
);

BUFx12f_ASAP7_75t_L g23 ( 
.A(n_1),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_3),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_15),
.Y(n_25)
);

INVx13_ASAP7_75t_L g26 ( 
.A(n_12),
.Y(n_26)
);

BUFx12f_ASAP7_75t_L g27 ( 
.A(n_10),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_15),
.Y(n_28)
);

INVx8_ASAP7_75t_L g29 ( 
.A(n_12),
.Y(n_29)
);

INVx2_ASAP7_75t_L g30 ( 
.A(n_9),
.Y(n_30)
);

INVx6_ASAP7_75t_L g31 ( 
.A(n_11),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_4),
.Y(n_32)
);

BUFx5_ASAP7_75t_L g33 ( 
.A(n_1),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_13),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_6),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_8),
.Y(n_36)
);

BUFx3_ASAP7_75t_L g37 ( 
.A(n_7),
.Y(n_37)
);

INVx8_ASAP7_75t_L g38 ( 
.A(n_15),
.Y(n_38)
);

INVx5_ASAP7_75t_L g39 ( 
.A(n_3),
.Y(n_39)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_13),
.Y(n_40)
);

INVx11_ASAP7_75t_L g41 ( 
.A(n_0),
.Y(n_41)
);

INVx8_ASAP7_75t_L g42 ( 
.A(n_3),
.Y(n_42)
);

CKINVDCx14_ASAP7_75t_R g43 ( 
.A(n_1),
.Y(n_43)
);

INVxp33_ASAP7_75t_L g44 ( 
.A(n_7),
.Y(n_44)
);

AND2x2_ASAP7_75t_L g45 ( 
.A(n_30),
.B(n_0),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_45),
.B(n_54),
.Y(n_103)
);

INVx11_ASAP7_75t_L g46 ( 
.A(n_22),
.Y(n_46)
);

BUFx10_ASAP7_75t_L g125 ( 
.A(n_46),
.Y(n_125)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_21),
.Y(n_47)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_47),
.Y(n_94)
);

INVx11_ASAP7_75t_L g48 ( 
.A(n_22),
.Y(n_48)
);

CKINVDCx6p67_ASAP7_75t_R g112 ( 
.A(n_48),
.Y(n_112)
);

INVx2_ASAP7_75t_L g49 ( 
.A(n_30),
.Y(n_49)
);

INVx2_ASAP7_75t_L g92 ( 
.A(n_49),
.Y(n_92)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_24),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g100 ( 
.A(n_50),
.Y(n_100)
);

INVx5_ASAP7_75t_L g51 ( 
.A(n_39),
.Y(n_51)
);

INVx5_ASAP7_75t_L g99 ( 
.A(n_51),
.Y(n_99)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_22),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g113 ( 
.A(n_52),
.B(n_58),
.Y(n_113)
);

INVx2_ASAP7_75t_SL g53 ( 
.A(n_23),
.Y(n_53)
);

BUFx3_ASAP7_75t_L g96 ( 
.A(n_53),
.Y(n_96)
);

BUFx4f_ASAP7_75t_SL g54 ( 
.A(n_33),
.Y(n_54)
);

AOI21xp33_ASAP7_75t_SL g55 ( 
.A1(n_41),
.A2(n_0),
.B(n_2),
.Y(n_55)
);

AOI21xp33_ASAP7_75t_L g91 ( 
.A1(n_55),
.A2(n_80),
.B(n_81),
.Y(n_91)
);

INVx2_ASAP7_75t_SL g56 ( 
.A(n_23),
.Y(n_56)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_56),
.Y(n_124)
);

INVx3_ASAP7_75t_L g57 ( 
.A(n_37),
.Y(n_57)
);

INVx3_ASAP7_75t_L g111 ( 
.A(n_57),
.Y(n_111)
);

CKINVDCx20_ASAP7_75t_R g58 ( 
.A(n_41),
.Y(n_58)
);

INVx8_ASAP7_75t_L g59 ( 
.A(n_33),
.Y(n_59)
);

INVx3_ASAP7_75t_L g119 ( 
.A(n_59),
.Y(n_119)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_23),
.Y(n_60)
);

INVx2_ASAP7_75t_L g93 ( 
.A(n_60),
.Y(n_93)
);

BUFx3_ASAP7_75t_L g61 ( 
.A(n_16),
.Y(n_61)
);

INVx4_ASAP7_75t_L g106 ( 
.A(n_61),
.Y(n_106)
);

BUFx4f_ASAP7_75t_L g62 ( 
.A(n_41),
.Y(n_62)
);

INVx3_ASAP7_75t_L g129 ( 
.A(n_62),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_SL g63 ( 
.A(n_44),
.B(n_0),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_63),
.B(n_64),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_25),
.B(n_2),
.Y(n_64)
);

INVx2_ASAP7_75t_L g65 ( 
.A(n_23),
.Y(n_65)
);

INVx2_ASAP7_75t_L g102 ( 
.A(n_65),
.Y(n_102)
);

INVx3_ASAP7_75t_L g66 ( 
.A(n_37),
.Y(n_66)
);

INVx4_ASAP7_75t_L g110 ( 
.A(n_66),
.Y(n_110)
);

CKINVDCx20_ASAP7_75t_R g67 ( 
.A(n_18),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g114 ( 
.A(n_67),
.B(n_72),
.Y(n_114)
);

INVx2_ASAP7_75t_L g68 ( 
.A(n_23),
.Y(n_68)
);

INVx2_ASAP7_75t_L g120 ( 
.A(n_68),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_25),
.B(n_2),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_69),
.B(n_71),
.Y(n_108)
);

BUFx6f_ASAP7_75t_L g70 ( 
.A(n_24),
.Y(n_70)
);

INVx6_ASAP7_75t_L g115 ( 
.A(n_70),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_18),
.B(n_3),
.Y(n_71)
);

CKINVDCx20_ASAP7_75t_R g72 ( 
.A(n_19),
.Y(n_72)
);

CKINVDCx20_ASAP7_75t_R g73 ( 
.A(n_19),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_73),
.B(n_75),
.Y(n_109)
);

INVx2_ASAP7_75t_L g74 ( 
.A(n_27),
.Y(n_74)
);

INVx2_ASAP7_75t_L g126 ( 
.A(n_74),
.Y(n_126)
);

INVx6_ASAP7_75t_SL g75 ( 
.A(n_26),
.Y(n_75)
);

INVx4_ASAP7_75t_SL g76 ( 
.A(n_26),
.Y(n_76)
);

AND2x2_ASAP7_75t_L g95 ( 
.A(n_76),
.B(n_78),
.Y(n_95)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_21),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g118 ( 
.A(n_77),
.B(n_79),
.Y(n_118)
);

INVx2_ASAP7_75t_L g78 ( 
.A(n_27),
.Y(n_78)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_32),
.Y(n_79)
);

INVx11_ASAP7_75t_L g80 ( 
.A(n_26),
.Y(n_80)
);

INVx11_ASAP7_75t_L g81 ( 
.A(n_17),
.Y(n_81)
);

CKINVDCx20_ASAP7_75t_R g82 ( 
.A(n_35),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g121 ( 
.A(n_82),
.B(n_84),
.Y(n_121)
);

INVx3_ASAP7_75t_L g83 ( 
.A(n_37),
.Y(n_83)
);

AND2x2_ASAP7_75t_L g101 ( 
.A(n_83),
.B(n_27),
.Y(n_101)
);

CKINVDCx20_ASAP7_75t_R g84 ( 
.A(n_35),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_SL g85 ( 
.A(n_67),
.B(n_17),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_SL g156 ( 
.A(n_85),
.B(n_90),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_SL g86 ( 
.A(n_45),
.B(n_32),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_SL g137 ( 
.A(n_86),
.B(n_117),
.Y(n_137)
);

AOI22xp33_ASAP7_75t_SL g87 ( 
.A1(n_59),
.A2(n_42),
.B1(n_29),
.B2(n_20),
.Y(n_87)
);

AOI22xp33_ASAP7_75t_SL g147 ( 
.A1(n_87),
.A2(n_88),
.B1(n_122),
.B2(n_132),
.Y(n_147)
);

AOI22xp33_ASAP7_75t_SL g88 ( 
.A1(n_59),
.A2(n_42),
.B1(n_29),
.B2(n_20),
.Y(n_88)
);

AOI22xp33_ASAP7_75t_L g89 ( 
.A1(n_63),
.A2(n_31),
.B1(n_28),
.B2(n_24),
.Y(n_89)
);

OAI22xp5_ASAP7_75t_L g146 ( 
.A1(n_89),
.A2(n_97),
.B1(n_107),
.B2(n_130),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_SL g90 ( 
.A(n_72),
.B(n_84),
.Y(n_90)
);

AOI22xp33_ASAP7_75t_L g97 ( 
.A1(n_45),
.A2(n_31),
.B1(n_28),
.B2(n_36),
.Y(n_97)
);

OAI21xp5_ASAP7_75t_L g98 ( 
.A1(n_55),
.A2(n_43),
.B(n_40),
.Y(n_98)
);

OAI21xp5_ASAP7_75t_L g150 ( 
.A1(n_98),
.A2(n_131),
.B(n_58),
.Y(n_150)
);

AND2x2_ASAP7_75t_L g135 ( 
.A(n_101),
.B(n_76),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_L g105 ( 
.A(n_47),
.B(n_40),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_L g176 ( 
.A(n_105),
.B(n_116),
.Y(n_176)
);

AOI22xp33_ASAP7_75t_L g107 ( 
.A1(n_73),
.A2(n_31),
.B1(n_28),
.B2(n_36),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_L g116 ( 
.A(n_77),
.B(n_34),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_L g117 ( 
.A(n_79),
.B(n_34),
.Y(n_117)
);

AOI22xp33_ASAP7_75t_SL g122 ( 
.A1(n_53),
.A2(n_29),
.B1(n_42),
.B2(n_38),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_L g123 ( 
.A(n_49),
.B(n_27),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_SL g169 ( 
.A(n_123),
.B(n_128),
.Y(n_169)
);

OAI22xp5_ASAP7_75t_L g127 ( 
.A1(n_50),
.A2(n_36),
.B1(n_38),
.B2(n_39),
.Y(n_127)
);

AOI22xp5_ASAP7_75t_L g157 ( 
.A1(n_127),
.A2(n_46),
.B1(n_54),
.B2(n_62),
.Y(n_157)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_82),
.B(n_43),
.Y(n_128)
);

AOI22xp33_ASAP7_75t_L g130 ( 
.A1(n_50),
.A2(n_38),
.B1(n_27),
.B2(n_39),
.Y(n_130)
);

AOI22xp5_ASAP7_75t_SL g131 ( 
.A1(n_57),
.A2(n_16),
.B1(n_5),
.B2(n_6),
.Y(n_131)
);

AOI22xp33_ASAP7_75t_SL g132 ( 
.A1(n_53),
.A2(n_16),
.B1(n_5),
.B2(n_6),
.Y(n_132)
);

NAND3xp33_ASAP7_75t_L g133 ( 
.A(n_104),
.B(n_75),
.C(n_81),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_L g185 ( 
.A(n_133),
.B(n_143),
.Y(n_185)
);

AOI22xp33_ASAP7_75t_L g134 ( 
.A1(n_94),
.A2(n_70),
.B1(n_66),
.B2(n_83),
.Y(n_134)
);

OAI22xp5_ASAP7_75t_L g187 ( 
.A1(n_134),
.A2(n_157),
.B1(n_119),
.B2(n_110),
.Y(n_187)
);

CKINVDCx16_ASAP7_75t_R g199 ( 
.A(n_135),
.Y(n_199)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_94),
.Y(n_136)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_136),
.Y(n_188)
);

NOR2xp33_ASAP7_75t_L g138 ( 
.A(n_90),
.B(n_56),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_SL g180 ( 
.A(n_138),
.B(n_149),
.Y(n_180)
);

INVx4_ASAP7_75t_SL g139 ( 
.A(n_124),
.Y(n_139)
);

INVx13_ASAP7_75t_L g211 ( 
.A(n_139),
.Y(n_211)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_124),
.Y(n_140)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_140),
.Y(n_193)
);

BUFx6f_ASAP7_75t_L g141 ( 
.A(n_100),
.Y(n_141)
);

INVx4_ASAP7_75t_L g207 ( 
.A(n_141),
.Y(n_207)
);

AND2x2_ASAP7_75t_L g142 ( 
.A(n_103),
.B(n_76),
.Y(n_142)
);

MAJIxp5_ASAP7_75t_L g182 ( 
.A(n_142),
.B(n_144),
.C(n_166),
.Y(n_182)
);

NAND3xp33_ASAP7_75t_L g143 ( 
.A(n_104),
.B(n_80),
.C(n_6),
.Y(n_143)
);

MAJIxp5_ASAP7_75t_L g144 ( 
.A(n_123),
.B(n_78),
.C(n_74),
.Y(n_144)
);

AOI22xp5_ASAP7_75t_SL g145 ( 
.A1(n_105),
.A2(n_61),
.B1(n_51),
.B2(n_56),
.Y(n_145)
);

OAI21xp5_ASAP7_75t_L g183 ( 
.A1(n_145),
.A2(n_160),
.B(n_101),
.Y(n_183)
);

CKINVDCx14_ASAP7_75t_R g148 ( 
.A(n_109),
.Y(n_148)
);

NOR2xp33_ASAP7_75t_L g192 ( 
.A(n_148),
.B(n_158),
.Y(n_192)
);

NOR2xp33_ASAP7_75t_L g149 ( 
.A(n_114),
.B(n_60),
.Y(n_149)
);

AOI21xp5_ASAP7_75t_L g184 ( 
.A1(n_150),
.A2(n_128),
.B(n_101),
.Y(n_184)
);

INVx6_ASAP7_75t_L g151 ( 
.A(n_100),
.Y(n_151)
);

INVx2_ASAP7_75t_L g186 ( 
.A(n_151),
.Y(n_186)
);

NOR2xp33_ASAP7_75t_L g152 ( 
.A(n_85),
.B(n_109),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_SL g190 ( 
.A(n_152),
.B(n_173),
.Y(n_190)
);

OAI22xp5_ASAP7_75t_SL g153 ( 
.A1(n_98),
.A2(n_70),
.B1(n_68),
.B2(n_65),
.Y(n_153)
);

AOI22xp5_ASAP7_75t_L g203 ( 
.A1(n_153),
.A2(n_155),
.B1(n_168),
.B2(n_175),
.Y(n_203)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_118),
.Y(n_154)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_154),
.Y(n_200)
);

OAI22xp5_ASAP7_75t_SL g155 ( 
.A1(n_103),
.A2(n_52),
.B1(n_16),
.B2(n_48),
.Y(n_155)
);

NAND3xp33_ASAP7_75t_L g158 ( 
.A(n_108),
.B(n_4),
.C(n_7),
.Y(n_158)
);

INVx3_ASAP7_75t_L g159 ( 
.A(n_96),
.Y(n_159)
);

HB1xp67_ASAP7_75t_L g214 ( 
.A(n_159),
.Y(n_214)
);

O2A1O1Ixp33_ASAP7_75t_L g160 ( 
.A1(n_91),
.A2(n_54),
.B(n_62),
.C(n_8),
.Y(n_160)
);

BUFx6f_ASAP7_75t_L g161 ( 
.A(n_100),
.Y(n_161)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_161),
.Y(n_201)
);

INVx13_ASAP7_75t_L g162 ( 
.A(n_95),
.Y(n_162)
);

CKINVDCx20_ASAP7_75t_R g191 ( 
.A(n_162),
.Y(n_191)
);

AO22x1_ASAP7_75t_SL g163 ( 
.A1(n_92),
.A2(n_54),
.B1(n_62),
.B2(n_8),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_L g197 ( 
.A(n_163),
.B(n_99),
.Y(n_197)
);

INVx8_ASAP7_75t_L g164 ( 
.A(n_115),
.Y(n_164)
);

INVxp67_ASAP7_75t_L g196 ( 
.A(n_164),
.Y(n_196)
);

BUFx2_ASAP7_75t_L g165 ( 
.A(n_129),
.Y(n_165)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_165),
.Y(n_217)
);

AND2x2_ASAP7_75t_L g166 ( 
.A(n_86),
.B(n_95),
.Y(n_166)
);

INVx2_ASAP7_75t_L g167 ( 
.A(n_92),
.Y(n_167)
);

NOR2xp33_ASAP7_75t_L g206 ( 
.A(n_167),
.B(n_170),
.Y(n_206)
);

OAI22xp5_ASAP7_75t_SL g168 ( 
.A1(n_116),
.A2(n_14),
.B1(n_7),
.B2(n_8),
.Y(n_168)
);

INVx4_ASAP7_75t_L g170 ( 
.A(n_96),
.Y(n_170)
);

AND2x2_ASAP7_75t_L g171 ( 
.A(n_95),
.B(n_14),
.Y(n_171)
);

MAJIxp5_ASAP7_75t_L g189 ( 
.A(n_171),
.B(n_102),
.C(n_126),
.Y(n_189)
);

BUFx6f_ASAP7_75t_L g172 ( 
.A(n_115),
.Y(n_172)
);

NOR2xp33_ASAP7_75t_L g209 ( 
.A(n_172),
.B(n_112),
.Y(n_209)
);

NOR2xp33_ASAP7_75t_L g173 ( 
.A(n_121),
.B(n_4),
.Y(n_173)
);

NOR2xp33_ASAP7_75t_L g174 ( 
.A(n_121),
.B(n_4),
.Y(n_174)
);

NOR2xp33_ASAP7_75t_SL g210 ( 
.A(n_174),
.B(n_9),
.Y(n_210)
);

OAI22xp5_ASAP7_75t_L g175 ( 
.A1(n_117),
.A2(n_9),
.B1(n_10),
.B2(n_11),
.Y(n_175)
);

INVx3_ASAP7_75t_SL g177 ( 
.A(n_115),
.Y(n_177)
);

INVxp67_ASAP7_75t_L g198 ( 
.A(n_177),
.Y(n_198)
);

OAI22xp5_ASAP7_75t_SL g178 ( 
.A1(n_131),
.A2(n_118),
.B1(n_108),
.B2(n_113),
.Y(n_178)
);

AOI22xp5_ASAP7_75t_L g205 ( 
.A1(n_178),
.A2(n_106),
.B1(n_99),
.B2(n_93),
.Y(n_205)
);

AOI22xp33_ASAP7_75t_L g179 ( 
.A1(n_153),
.A2(n_111),
.B1(n_129),
.B2(n_110),
.Y(n_179)
);

OAI21xp33_ASAP7_75t_SL g252 ( 
.A1(n_179),
.A2(n_184),
.B(n_197),
.Y(n_252)
);

AND2x2_ASAP7_75t_SL g181 ( 
.A(n_144),
.B(n_126),
.Y(n_181)
);

AND2x2_ASAP7_75t_L g221 ( 
.A(n_181),
.B(n_183),
.Y(n_221)
);

AOI22xp5_ASAP7_75t_L g224 ( 
.A1(n_187),
.A2(n_195),
.B1(n_204),
.B2(n_208),
.Y(n_224)
);

XNOR2xp5_ASAP7_75t_L g222 ( 
.A(n_189),
.B(n_212),
.Y(n_222)
);

CKINVDCx20_ASAP7_75t_R g194 ( 
.A(n_139),
.Y(n_194)
);

NOR2xp33_ASAP7_75t_L g220 ( 
.A(n_194),
.B(n_205),
.Y(n_220)
);

OAI22xp5_ASAP7_75t_L g195 ( 
.A1(n_176),
.A2(n_127),
.B1(n_111),
.B2(n_119),
.Y(n_195)
);

AND2x4_ASAP7_75t_SL g202 ( 
.A(n_162),
.B(n_120),
.Y(n_202)
);

INVx1_ASAP7_75t_SL g228 ( 
.A(n_202),
.Y(n_228)
);

OAI22xp5_ASAP7_75t_L g204 ( 
.A1(n_176),
.A2(n_120),
.B1(n_102),
.B2(n_93),
.Y(n_204)
);

OAI22xp5_ASAP7_75t_SL g208 ( 
.A1(n_150),
.A2(n_112),
.B1(n_125),
.B2(n_106),
.Y(n_208)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_209),
.Y(n_233)
);

NOR2xp33_ASAP7_75t_SL g247 ( 
.A(n_210),
.B(n_139),
.Y(n_247)
);

MAJIxp5_ASAP7_75t_L g212 ( 
.A(n_169),
.B(n_125),
.C(n_112),
.Y(n_212)
);

AOI22xp5_ASAP7_75t_L g213 ( 
.A1(n_146),
.A2(n_160),
.B1(n_178),
.B2(n_155),
.Y(n_213)
);

OAI22xp5_ASAP7_75t_L g240 ( 
.A1(n_213),
.A2(n_177),
.B1(n_167),
.B2(n_151),
.Y(n_240)
);

NAND2xp5_ASAP7_75t_L g215 ( 
.A(n_154),
.B(n_10),
.Y(n_215)
);

NAND2xp5_ASAP7_75t_L g241 ( 
.A(n_215),
.B(n_11),
.Y(n_241)
);

OAI32xp33_ASAP7_75t_L g216 ( 
.A1(n_137),
.A2(n_125),
.A3(n_112),
.B1(n_12),
.B2(n_13),
.Y(n_216)
);

NOR2xp33_ASAP7_75t_L g242 ( 
.A(n_216),
.B(n_218),
.Y(n_242)
);

OAI32xp33_ASAP7_75t_L g218 ( 
.A1(n_156),
.A2(n_125),
.A3(n_11),
.B1(n_12),
.B2(n_13),
.Y(n_218)
);

AND2x6_ASAP7_75t_L g219 ( 
.A(n_156),
.B(n_10),
.Y(n_219)
);

AOI21xp33_ASAP7_75t_L g225 ( 
.A1(n_219),
.A2(n_175),
.B(n_166),
.Y(n_225)
);

CKINVDCx20_ASAP7_75t_R g223 ( 
.A(n_214),
.Y(n_223)
);

NOR2xp33_ASAP7_75t_L g271 ( 
.A(n_223),
.B(n_229),
.Y(n_271)
);

AOI21xp5_ASAP7_75t_SL g255 ( 
.A1(n_225),
.A2(n_184),
.B(n_182),
.Y(n_255)
);

INVx2_ASAP7_75t_L g226 ( 
.A(n_186),
.Y(n_226)
);

INVx1_ASAP7_75t_SL g280 ( 
.A(n_226),
.Y(n_280)
);

AOI22xp5_ASAP7_75t_L g227 ( 
.A1(n_197),
.A2(n_146),
.B1(n_166),
.B2(n_168),
.Y(n_227)
);

OAI22xp5_ASAP7_75t_L g282 ( 
.A1(n_227),
.A2(n_230),
.B1(n_232),
.B2(n_185),
.Y(n_282)
);

CKINVDCx20_ASAP7_75t_R g229 ( 
.A(n_206),
.Y(n_229)
);

AOI22xp5_ASAP7_75t_L g230 ( 
.A1(n_183),
.A2(n_136),
.B1(n_147),
.B2(n_142),
.Y(n_230)
);

CKINVDCx20_ASAP7_75t_R g231 ( 
.A(n_206),
.Y(n_231)
);

NAND2xp5_ASAP7_75t_L g262 ( 
.A(n_231),
.B(n_234),
.Y(n_262)
);

AOI22xp5_ASAP7_75t_L g232 ( 
.A1(n_195),
.A2(n_142),
.B1(n_171),
.B2(n_163),
.Y(n_232)
);

CKINVDCx20_ASAP7_75t_R g234 ( 
.A(n_204),
.Y(n_234)
);

OAI22xp5_ASAP7_75t_SL g235 ( 
.A1(n_213),
.A2(n_157),
.B1(n_145),
.B2(n_163),
.Y(n_235)
);

AOI22xp5_ASAP7_75t_L g254 ( 
.A1(n_235),
.A2(n_240),
.B1(n_187),
.B2(n_252),
.Y(n_254)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_188),
.Y(n_236)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_236),
.Y(n_260)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_188),
.Y(n_237)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_237),
.Y(n_261)
);

OAI21xp33_ASAP7_75t_L g238 ( 
.A1(n_191),
.A2(n_171),
.B(n_135),
.Y(n_238)
);

INVxp67_ASAP7_75t_L g268 ( 
.A(n_238),
.Y(n_268)
);

AOI22xp33_ASAP7_75t_L g239 ( 
.A1(n_191),
.A2(n_135),
.B1(n_140),
.B2(n_164),
.Y(n_239)
);

OA22x2_ASAP7_75t_L g275 ( 
.A1(n_239),
.A2(n_245),
.B1(n_194),
.B2(n_217),
.Y(n_275)
);

NAND2xp5_ASAP7_75t_SL g270 ( 
.A(n_241),
.B(n_247),
.Y(n_270)
);

NAND2xp5_ASAP7_75t_L g243 ( 
.A(n_181),
.B(n_172),
.Y(n_243)
);

NAND2xp5_ASAP7_75t_L g266 ( 
.A(n_243),
.B(n_246),
.Y(n_266)
);

AOI22xp33_ASAP7_75t_SL g244 ( 
.A1(n_208),
.A2(n_159),
.B1(n_170),
.B2(n_177),
.Y(n_244)
);

INVxp67_ASAP7_75t_L g272 ( 
.A(n_244),
.Y(n_272)
);

AOI22xp33_ASAP7_75t_L g245 ( 
.A1(n_200),
.A2(n_165),
.B1(n_141),
.B2(n_161),
.Y(n_245)
);

NAND2xp5_ASAP7_75t_L g246 ( 
.A(n_181),
.B(n_165),
.Y(n_246)
);

HB1xp67_ASAP7_75t_L g248 ( 
.A(n_217),
.Y(n_248)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_248),
.Y(n_263)
);

NOR2xp33_ASAP7_75t_L g249 ( 
.A(n_190),
.B(n_180),
.Y(n_249)
);

NAND2xp5_ASAP7_75t_L g267 ( 
.A(n_249),
.B(n_250),
.Y(n_267)
);

INVx2_ASAP7_75t_L g250 ( 
.A(n_186),
.Y(n_250)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_193),
.Y(n_251)
);

NAND2xp5_ASAP7_75t_L g269 ( 
.A(n_251),
.B(n_253),
.Y(n_269)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_193),
.Y(n_253)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_254),
.Y(n_291)
);

OAI21xp5_ASAP7_75t_SL g286 ( 
.A1(n_255),
.A2(n_256),
.B(n_243),
.Y(n_286)
);

AOI22xp5_ASAP7_75t_SL g256 ( 
.A1(n_235),
.A2(n_180),
.B1(n_182),
.B2(n_212),
.Y(n_256)
);

AOI22xp5_ASAP7_75t_L g257 ( 
.A1(n_240),
.A2(n_181),
.B1(n_200),
.B2(n_203),
.Y(n_257)
);

AOI22xp5_ASAP7_75t_L g300 ( 
.A1(n_257),
.A2(n_259),
.B1(n_264),
.B2(n_276),
.Y(n_300)
);

XNOR2xp5_ASAP7_75t_L g258 ( 
.A(n_222),
.B(n_189),
.Y(n_258)
);

XNOR2xp5_ASAP7_75t_SL g294 ( 
.A(n_258),
.B(n_224),
.Y(n_294)
);

OAI22xp5_ASAP7_75t_SL g259 ( 
.A1(n_227),
.A2(n_203),
.B1(n_205),
.B2(n_199),
.Y(n_259)
);

AOI22xp5_ASAP7_75t_L g264 ( 
.A1(n_234),
.A2(n_221),
.B1(n_233),
.B2(n_246),
.Y(n_264)
);

OAI21xp5_ASAP7_75t_SL g265 ( 
.A1(n_230),
.A2(n_199),
.B(n_185),
.Y(n_265)
);

OAI21xp5_ASAP7_75t_L g298 ( 
.A1(n_265),
.A2(n_283),
.B(n_220),
.Y(n_298)
);

BUFx10_ASAP7_75t_L g273 ( 
.A(n_223),
.Y(n_273)
);

BUFx12_ASAP7_75t_L g306 ( 
.A(n_273),
.Y(n_306)
);

AOI22x1_ASAP7_75t_L g274 ( 
.A1(n_221),
.A2(n_216),
.B1(n_218),
.B2(n_219),
.Y(n_274)
);

CKINVDCx16_ASAP7_75t_R g287 ( 
.A(n_274),
.Y(n_287)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_275),
.Y(n_292)
);

OAI22xp5_ASAP7_75t_SL g276 ( 
.A1(n_224),
.A2(n_219),
.B1(n_190),
.B2(n_215),
.Y(n_276)
);

AOI22xp5_ASAP7_75t_L g277 ( 
.A1(n_221),
.A2(n_202),
.B1(n_196),
.B2(n_201),
.Y(n_277)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_277),
.Y(n_295)
);

CKINVDCx20_ASAP7_75t_R g278 ( 
.A(n_249),
.Y(n_278)
);

NOR2xp33_ASAP7_75t_L g285 ( 
.A(n_278),
.B(n_281),
.Y(n_285)
);

NAND2xp5_ASAP7_75t_L g279 ( 
.A(n_229),
.B(n_202),
.Y(n_279)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_279),
.Y(n_299)
);

NAND2xp5_ASAP7_75t_L g281 ( 
.A(n_231),
.B(n_233),
.Y(n_281)
);

NAND2xp5_ASAP7_75t_SL g289 ( 
.A(n_281),
.B(n_253),
.Y(n_289)
);

AO21x1_ASAP7_75t_L g284 ( 
.A1(n_282),
.A2(n_232),
.B(n_242),
.Y(n_284)
);

OAI21xp5_ASAP7_75t_L g283 ( 
.A1(n_228),
.A2(n_192),
.B(n_202),
.Y(n_283)
);

OAI22xp5_ASAP7_75t_L g321 ( 
.A1(n_284),
.A2(n_301),
.B1(n_307),
.B2(n_283),
.Y(n_321)
);

NAND3xp33_ASAP7_75t_L g319 ( 
.A(n_285),
.B(n_286),
.C(n_304),
.Y(n_319)
);

INVx4_ASAP7_75t_L g288 ( 
.A(n_273),
.Y(n_288)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_288),
.Y(n_310)
);

NAND2xp5_ASAP7_75t_L g318 ( 
.A(n_289),
.B(n_297),
.Y(n_318)
);

MAJIxp5_ASAP7_75t_L g290 ( 
.A(n_258),
.B(n_222),
.C(n_256),
.Y(n_290)
);

MAJIxp5_ASAP7_75t_L g320 ( 
.A(n_290),
.B(n_293),
.C(n_296),
.Y(n_320)
);

MAJIxp5_ASAP7_75t_L g293 ( 
.A(n_255),
.B(n_264),
.C(n_282),
.Y(n_293)
);

XNOR2xp5_ASAP7_75t_SL g314 ( 
.A(n_294),
.B(n_308),
.Y(n_314)
);

MAJIxp5_ASAP7_75t_L g296 ( 
.A(n_268),
.B(n_228),
.C(n_251),
.Y(n_296)
);

CKINVDCx20_ASAP7_75t_R g297 ( 
.A(n_269),
.Y(n_297)
);

MAJIxp5_ASAP7_75t_L g325 ( 
.A(n_298),
.B(n_303),
.C(n_305),
.Y(n_325)
);

AOI22xp5_ASAP7_75t_SL g301 ( 
.A1(n_268),
.A2(n_247),
.B1(n_242),
.B2(n_225),
.Y(n_301)
);

CKINVDCx20_ASAP7_75t_R g302 ( 
.A(n_269),
.Y(n_302)
);

CKINVDCx20_ASAP7_75t_R g328 ( 
.A(n_302),
.Y(n_328)
);

MAJIxp5_ASAP7_75t_L g303 ( 
.A(n_265),
.B(n_236),
.C(n_237),
.Y(n_303)
);

NOR2xp33_ASAP7_75t_L g304 ( 
.A(n_278),
.B(n_210),
.Y(n_304)
);

XOR2xp5_ASAP7_75t_L g305 ( 
.A(n_262),
.B(n_220),
.Y(n_305)
);

NOR2xp33_ASAP7_75t_SL g307 ( 
.A(n_270),
.B(n_192),
.Y(n_307)
);

XOR2xp5_ASAP7_75t_L g308 ( 
.A(n_262),
.B(n_241),
.Y(n_308)
);

OAI22xp5_ASAP7_75t_SL g309 ( 
.A1(n_284),
.A2(n_254),
.B1(n_257),
.B2(n_272),
.Y(n_309)
);

AOI22xp5_ASAP7_75t_L g336 ( 
.A1(n_309),
.A2(n_328),
.B1(n_312),
.B2(n_323),
.Y(n_336)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_305),
.Y(n_311)
);

NAND2xp5_ASAP7_75t_L g332 ( 
.A(n_311),
.B(n_312),
.Y(n_332)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_299),
.Y(n_312)
);

AOI22xp5_ASAP7_75t_L g313 ( 
.A1(n_291),
.A2(n_259),
.B1(n_276),
.B2(n_272),
.Y(n_313)
);

OAI22xp5_ASAP7_75t_L g333 ( 
.A1(n_313),
.A2(n_315),
.B1(n_316),
.B2(n_322),
.Y(n_333)
);

AOI22xp5_ASAP7_75t_L g315 ( 
.A1(n_291),
.A2(n_266),
.B1(n_267),
.B2(n_279),
.Y(n_315)
);

AOI22xp5_ASAP7_75t_L g316 ( 
.A1(n_295),
.A2(n_292),
.B1(n_287),
.B2(n_293),
.Y(n_316)
);

AOI22xp5_ASAP7_75t_SL g317 ( 
.A1(n_295),
.A2(n_292),
.B1(n_303),
.B2(n_296),
.Y(n_317)
);

OAI21xp5_ASAP7_75t_SL g338 ( 
.A1(n_317),
.A2(n_300),
.B(n_286),
.Y(n_338)
);

AOI22xp5_ASAP7_75t_SL g331 ( 
.A1(n_321),
.A2(n_298),
.B1(n_301),
.B2(n_290),
.Y(n_331)
);

AOI22xp5_ASAP7_75t_L g322 ( 
.A1(n_287),
.A2(n_266),
.B1(n_267),
.B2(n_274),
.Y(n_322)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_299),
.Y(n_323)
);

AOI22xp33_ASAP7_75t_SL g337 ( 
.A1(n_323),
.A2(n_327),
.B1(n_280),
.B2(n_263),
.Y(n_337)
);

OAI22xp5_ASAP7_75t_L g324 ( 
.A1(n_284),
.A2(n_271),
.B1(n_274),
.B2(n_277),
.Y(n_324)
);

NAND2xp5_ASAP7_75t_SL g340 ( 
.A(n_324),
.B(n_209),
.Y(n_340)
);

AOI22xp5_ASAP7_75t_L g326 ( 
.A1(n_297),
.A2(n_273),
.B1(n_261),
.B2(n_260),
.Y(n_326)
);

OAI22xp5_ASAP7_75t_L g339 ( 
.A1(n_326),
.A2(n_329),
.B1(n_263),
.B2(n_300),
.Y(n_339)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_288),
.Y(n_327)
);

AOI22xp5_ASAP7_75t_L g329 ( 
.A1(n_302),
.A2(n_273),
.B1(n_261),
.B2(n_260),
.Y(n_329)
);

NOR2xp33_ASAP7_75t_L g330 ( 
.A(n_311),
.B(n_307),
.Y(n_330)
);

NAND2xp5_ASAP7_75t_L g357 ( 
.A(n_330),
.B(n_334),
.Y(n_357)
);

AOI21xp5_ASAP7_75t_L g350 ( 
.A1(n_331),
.A2(n_337),
.B(n_338),
.Y(n_350)
);

NOR2xp33_ASAP7_75t_L g334 ( 
.A(n_319),
.B(n_308),
.Y(n_334)
);

NOR2xp33_ASAP7_75t_L g335 ( 
.A(n_316),
.B(n_294),
.Y(n_335)
);

NAND2xp5_ASAP7_75t_L g359 ( 
.A(n_335),
.B(n_336),
.Y(n_359)
);

INVx1_ASAP7_75t_L g352 ( 
.A(n_339),
.Y(n_352)
);

NOR2xp33_ASAP7_75t_L g354 ( 
.A(n_340),
.B(n_344),
.Y(n_354)
);

NAND2xp5_ASAP7_75t_SL g341 ( 
.A(n_325),
.B(n_280),
.Y(n_341)
);

NAND2xp5_ASAP7_75t_SL g348 ( 
.A(n_341),
.B(n_342),
.Y(n_348)
);

OAI22xp5_ASAP7_75t_L g342 ( 
.A1(n_315),
.A2(n_275),
.B1(n_306),
.B2(n_201),
.Y(n_342)
);

AOI21xp5_ASAP7_75t_L g343 ( 
.A1(n_317),
.A2(n_306),
.B(n_275),
.Y(n_343)
);

AOI21xp5_ASAP7_75t_L g349 ( 
.A1(n_343),
.A2(n_313),
.B(n_326),
.Y(n_349)
);

CKINVDCx20_ASAP7_75t_R g344 ( 
.A(n_318),
.Y(n_344)
);

XOR2xp5_ASAP7_75t_L g345 ( 
.A(n_314),
.B(n_306),
.Y(n_345)
);

XNOR2xp5_ASAP7_75t_SL g353 ( 
.A(n_345),
.B(n_314),
.Y(n_353)
);

XNOR2xp5_ASAP7_75t_L g346 ( 
.A(n_325),
.B(n_226),
.Y(n_346)
);

XNOR2xp5_ASAP7_75t_L g351 ( 
.A(n_346),
.B(n_329),
.Y(n_351)
);

FAx1_ASAP7_75t_SL g347 ( 
.A(n_332),
.B(n_320),
.CI(n_318),
.CON(n_347),
.SN(n_347)
);

NOR2xp33_ASAP7_75t_L g361 ( 
.A(n_347),
.B(n_355),
.Y(n_361)
);

OAI21xp5_ASAP7_75t_SL g366 ( 
.A1(n_349),
.A2(n_356),
.B(n_358),
.Y(n_366)
);

XOR2xp5_ASAP7_75t_L g369 ( 
.A(n_351),
.B(n_353),
.Y(n_369)
);

XNOR2xp5_ASAP7_75t_L g355 ( 
.A(n_346),
.B(n_320),
.Y(n_355)
);

AOI21xp5_ASAP7_75t_L g356 ( 
.A1(n_338),
.A2(n_322),
.B(n_327),
.Y(n_356)
);

AOI21xp5_ASAP7_75t_L g358 ( 
.A1(n_343),
.A2(n_310),
.B(n_306),
.Y(n_358)
);

OAI22xp5_ASAP7_75t_SL g360 ( 
.A1(n_352),
.A2(n_336),
.B1(n_331),
.B2(n_350),
.Y(n_360)
);

AOI22xp5_ASAP7_75t_L g371 ( 
.A1(n_360),
.A2(n_347),
.B1(n_353),
.B2(n_250),
.Y(n_371)
);

MAJIxp5_ASAP7_75t_L g362 ( 
.A(n_355),
.B(n_345),
.C(n_333),
.Y(n_362)
);

NAND2xp5_ASAP7_75t_L g376 ( 
.A(n_362),
.B(n_363),
.Y(n_376)
);

OAI21x1_ASAP7_75t_L g363 ( 
.A1(n_359),
.A2(n_332),
.B(n_344),
.Y(n_363)
);

NAND2xp5_ASAP7_75t_L g364 ( 
.A(n_354),
.B(n_339),
.Y(n_364)
);

OAI21xp5_ASAP7_75t_L g370 ( 
.A1(n_364),
.A2(n_349),
.B(n_310),
.Y(n_370)
);

MAJIxp5_ASAP7_75t_L g365 ( 
.A(n_351),
.B(n_333),
.C(n_309),
.Y(n_365)
);

NOR2xp33_ASAP7_75t_L g375 ( 
.A(n_365),
.B(n_368),
.Y(n_375)
);

CKINVDCx20_ASAP7_75t_R g367 ( 
.A(n_348),
.Y(n_367)
);

AOI21xp5_ASAP7_75t_L g373 ( 
.A1(n_367),
.A2(n_207),
.B(n_211),
.Y(n_373)
);

FAx1_ASAP7_75t_SL g368 ( 
.A(n_357),
.B(n_342),
.CI(n_275),
.CON(n_368),
.SN(n_368)
);

INVx1_ASAP7_75t_L g381 ( 
.A(n_370),
.Y(n_381)
);

XNOR2xp5_ASAP7_75t_L g383 ( 
.A(n_371),
.B(n_372),
.Y(n_383)
);

AOI21xp5_ASAP7_75t_SL g372 ( 
.A1(n_366),
.A2(n_198),
.B(n_211),
.Y(n_372)
);

CKINVDCx20_ASAP7_75t_R g384 ( 
.A(n_373),
.Y(n_384)
);

NOR2xp33_ASAP7_75t_SL g374 ( 
.A(n_361),
.B(n_207),
.Y(n_374)
);

NOR2x1_ASAP7_75t_L g382 ( 
.A(n_374),
.B(n_364),
.Y(n_382)
);

XNOR2xp5_ASAP7_75t_L g377 ( 
.A(n_362),
.B(n_211),
.Y(n_377)
);

MAJIxp5_ASAP7_75t_L g380 ( 
.A(n_377),
.B(n_378),
.C(n_369),
.Y(n_380)
);

XOR2xp5_ASAP7_75t_L g378 ( 
.A(n_369),
.B(n_366),
.Y(n_378)
);

XNOR2x2_ASAP7_75t_SL g379 ( 
.A(n_378),
.B(n_363),
.Y(n_379)
);

INVx1_ASAP7_75t_L g386 ( 
.A(n_379),
.Y(n_386)
);

NAND2xp5_ASAP7_75t_SL g385 ( 
.A(n_380),
.B(n_382),
.Y(n_385)
);

AOI322xp5_ASAP7_75t_L g387 ( 
.A1(n_381),
.A2(n_375),
.A3(n_367),
.B1(n_360),
.B2(n_376),
.C1(n_368),
.C2(n_372),
.Y(n_387)
);

INVxp67_ASAP7_75t_L g390 ( 
.A(n_387),
.Y(n_390)
);

A2O1A1O1Ixp25_ASAP7_75t_L g388 ( 
.A1(n_379),
.A2(n_365),
.B(n_368),
.C(n_377),
.D(n_380),
.Y(n_388)
);

OAI21xp5_ASAP7_75t_L g389 ( 
.A1(n_388),
.A2(n_385),
.B(n_386),
.Y(n_389)
);

OAI21xp5_ASAP7_75t_L g391 ( 
.A1(n_389),
.A2(n_390),
.B(n_382),
.Y(n_391)
);

NAND2xp5_ASAP7_75t_SL g392 ( 
.A(n_391),
.B(n_384),
.Y(n_392)
);

XOR2xp5_ASAP7_75t_L g393 ( 
.A(n_392),
.B(n_383),
.Y(n_393)
);


endmodule