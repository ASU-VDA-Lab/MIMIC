module fake_jpeg_30051_n_123 (n_13, n_21, n_33, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_40, n_19, n_18, n_20, n_35, n_4, n_34, n_30, n_39, n_16, n_3, n_0, n_24, n_28, n_38, n_26, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_12, n_32, n_8, n_15, n_7, n_123);

input n_13;
input n_21;
input n_33;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_4;
input n_34;
input n_30;
input n_39;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_123;

wire n_117;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_73;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_42;
wire n_49;
wire n_76;
wire n_88;
wire n_116;
wire n_114;
wire n_74;
wire n_103;
wire n_50;
wire n_57;
wire n_119;
wire n_69;
wire n_83;
wire n_71;
wire n_80;
wire n_81;
wire n_109;
wire n_113;
wire n_106;
wire n_111;
wire n_44;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_121;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_56;
wire n_79;
wire n_67;
wire n_53;
wire n_54;
wire n_93;
wire n_91;
wire n_101;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_112;
wire n_95;
wire n_97;
wire n_62;
wire n_120;
wire n_43;
wire n_100;
wire n_118;
wire n_82;
wire n_96;

NAND2xp5_ASAP7_75t_L g41 ( 
.A(n_4),
.B(n_26),
.Y(n_41)
);

BUFx12f_ASAP7_75t_L g42 ( 
.A(n_30),
.Y(n_42)
);

INVx3_ASAP7_75t_L g43 ( 
.A(n_9),
.Y(n_43)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_19),
.Y(n_44)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_27),
.Y(n_45)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_12),
.Y(n_46)
);

INVx13_ASAP7_75t_L g47 ( 
.A(n_23),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_7),
.B(n_25),
.Y(n_48)
);

BUFx6f_ASAP7_75t_SL g49 ( 
.A(n_2),
.Y(n_49)
);

INVx5_ASAP7_75t_L g50 ( 
.A(n_18),
.Y(n_50)
);

INVx6_ASAP7_75t_SL g51 ( 
.A(n_39),
.Y(n_51)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_15),
.Y(n_52)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_17),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_41),
.B(n_44),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_54),
.B(n_42),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_L g55 ( 
.A(n_48),
.B(n_0),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_L g68 ( 
.A(n_55),
.B(n_58),
.Y(n_68)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_49),
.Y(n_56)
);

INVx3_ASAP7_75t_L g66 ( 
.A(n_56),
.Y(n_66)
);

BUFx12f_ASAP7_75t_L g57 ( 
.A(n_47),
.Y(n_57)
);

INVx3_ASAP7_75t_L g73 ( 
.A(n_57),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_L g58 ( 
.A(n_42),
.B(n_0),
.Y(n_58)
);

BUFx4f_ASAP7_75t_SL g59 ( 
.A(n_47),
.Y(n_59)
);

INVx13_ASAP7_75t_L g74 ( 
.A(n_59),
.Y(n_74)
);

AOI22xp33_ASAP7_75t_SL g60 ( 
.A1(n_42),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_60)
);

AOI22xp33_ASAP7_75t_SL g71 ( 
.A1(n_60),
.A2(n_50),
.B1(n_43),
.B2(n_51),
.Y(n_71)
);

INVx4_ASAP7_75t_L g61 ( 
.A(n_49),
.Y(n_61)
);

BUFx2_ASAP7_75t_L g62 ( 
.A(n_61),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_63),
.B(n_67),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_59),
.B(n_53),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_SL g78 ( 
.A(n_64),
.B(n_65),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_SL g65 ( 
.A(n_57),
.B(n_52),
.Y(n_65)
);

OR2x2_ASAP7_75t_L g67 ( 
.A(n_57),
.B(n_1),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_L g69 ( 
.A(n_59),
.B(n_45),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_L g77 ( 
.A(n_69),
.B(n_70),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_61),
.B(n_46),
.Y(n_70)
);

OAI22xp5_ASAP7_75t_SL g82 ( 
.A1(n_71),
.A2(n_4),
.B1(n_5),
.B2(n_6),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_60),
.B(n_43),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_L g79 ( 
.A(n_72),
.B(n_3),
.Y(n_79)
);

AOI22xp5_ASAP7_75t_L g75 ( 
.A1(n_66),
.A2(n_50),
.B1(n_51),
.B2(n_24),
.Y(n_75)
);

AOI22xp5_ASAP7_75t_L g104 ( 
.A1(n_75),
.A2(n_82),
.B1(n_84),
.B2(n_29),
.Y(n_104)
);

OAI21xp5_ASAP7_75t_L g96 ( 
.A1(n_79),
.A2(n_14),
.B(n_16),
.Y(n_96)
);

CKINVDCx16_ASAP7_75t_R g80 ( 
.A(n_67),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_80),
.B(n_75),
.Y(n_101)
);

INVx6_ASAP7_75t_SL g81 ( 
.A(n_74),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g93 ( 
.A(n_81),
.B(n_88),
.Y(n_93)
);

HB1xp67_ASAP7_75t_L g83 ( 
.A(n_66),
.Y(n_83)
);

INVx2_ASAP7_75t_L g90 ( 
.A(n_83),
.Y(n_90)
);

AOI22xp5_ASAP7_75t_L g84 ( 
.A1(n_71),
.A2(n_5),
.B1(n_6),
.B2(n_7),
.Y(n_84)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_62),
.Y(n_85)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_85),
.Y(n_92)
);

BUFx3_ASAP7_75t_L g86 ( 
.A(n_73),
.Y(n_86)
);

BUFx3_ASAP7_75t_L g91 ( 
.A(n_86),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_68),
.B(n_8),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_SL g98 ( 
.A(n_87),
.B(n_89),
.Y(n_98)
);

BUFx24_ASAP7_75t_L g88 ( 
.A(n_74),
.Y(n_88)
);

CKINVDCx14_ASAP7_75t_R g103 ( 
.A(n_88),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_73),
.B(n_10),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g112 ( 
.A(n_93),
.B(n_100),
.Y(n_112)
);

MAJIxp5_ASAP7_75t_SL g94 ( 
.A(n_76),
.B(n_11),
.C(n_13),
.Y(n_94)
);

MAJIxp5_ASAP7_75t_SL g111 ( 
.A(n_94),
.B(n_35),
.C(n_36),
.Y(n_111)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_83),
.Y(n_95)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_95),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_SL g106 ( 
.A(n_96),
.B(n_31),
.Y(n_106)
);

MAJIxp5_ASAP7_75t_L g97 ( 
.A(n_77),
.B(n_20),
.C(n_21),
.Y(n_97)
);

XNOR2xp5_ASAP7_75t_L g107 ( 
.A(n_97),
.B(n_99),
.Y(n_107)
);

MAJIxp5_ASAP7_75t_L g99 ( 
.A(n_78),
.B(n_22),
.C(n_28),
.Y(n_99)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_86),
.Y(n_100)
);

XNOR2xp5_ASAP7_75t_L g108 ( 
.A(n_101),
.B(n_102),
.Y(n_108)
);

XOR2xp5_ASAP7_75t_L g102 ( 
.A(n_88),
.B(n_62),
.Y(n_102)
);

OAI22xp5_ASAP7_75t_L g109 ( 
.A1(n_104),
.A2(n_32),
.B1(n_33),
.B2(n_34),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_SL g105 ( 
.A(n_98),
.B(n_101),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_L g113 ( 
.A(n_105),
.B(n_106),
.Y(n_113)
);

XOR2xp5_ASAP7_75t_L g115 ( 
.A(n_109),
.B(n_111),
.Y(n_115)
);

MAJIxp5_ASAP7_75t_L g114 ( 
.A(n_108),
.B(n_92),
.C(n_90),
.Y(n_114)
);

XNOR2xp5_ASAP7_75t_L g117 ( 
.A(n_114),
.B(n_116),
.Y(n_117)
);

MAJIxp5_ASAP7_75t_L g116 ( 
.A(n_107),
.B(n_91),
.C(n_103),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_SL g118 ( 
.A(n_113),
.B(n_112),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_L g119 ( 
.A(n_118),
.B(n_112),
.Y(n_119)
);

AOI21xp5_ASAP7_75t_L g120 ( 
.A1(n_119),
.A2(n_110),
.B(n_117),
.Y(n_120)
);

OAI31xp33_ASAP7_75t_L g121 ( 
.A1(n_120),
.A2(n_115),
.A3(n_103),
.B(n_91),
.Y(n_121)
);

OAI21xp5_ASAP7_75t_L g122 ( 
.A1(n_121),
.A2(n_37),
.B(n_38),
.Y(n_122)
);

XNOR2xp5_ASAP7_75t_L g123 ( 
.A(n_122),
.B(n_40),
.Y(n_123)
);


endmodule