module fake_jpeg_13325_n_574 (n_13, n_1, n_10, n_6, n_14, n_18, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_574);

input n_13;
input n_1;
input n_10;
input n_6;
input n_14;
input n_18;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_574;

wire n_529;
wire n_390;
wire n_552;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_525;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_519;
wire n_276;
wire n_143;
wire n_431;
wire n_102;
wire n_549;
wire n_196;
wire n_66;
wire n_374;
wire n_566;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_172;
wire n_547;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_513;
wire n_283;
wire n_107;
wire n_490;
wire n_517;
wire n_415;
wire n_479;
wire n_543;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_542;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_559;
wire n_48;
wire n_465;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_221;
wire n_256;
wire n_454;
wire n_540;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_571;
wire n_82;
wire n_155;
wire n_508;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_569;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_544;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_530;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_557;
wire n_408;
wire n_80;
wire n_562;
wire n_204;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_298;
wire n_106;
wire n_545;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_474;
wire n_539;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_511;
wire n_305;
wire n_161;
wire n_441;
wire n_555;
wire n_342;
wire n_101;
wire n_226;
wire n_509;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_573;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_560;
wire n_190;
wire n_510;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_536;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_537;
wire n_110;
wire n_531;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_570;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_352;
wire n_350;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_554;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_523;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_533;
wire n_296;
wire n_384;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_491;
wire n_24;
wire n_526;
wire n_467;
wire n_269;
wire n_572;
wire n_546;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_473;
wire n_45;
wire n_520;
wire n_476;
wire n_337;
wire n_317;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_481;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_522;
wire n_333;
wire n_518;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_565;
wire n_302;
wire n_216;
wire n_528;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_199;
wire n_260;
wire n_550;
wire n_413;
wire n_275;
wire n_494;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_551;
wire n_36;
wire n_62;
wire n_492;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_567;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_515;
wire n_347;
wire n_521;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_538;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_534;
wire n_472;
wire n_279;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_484;
wire n_568;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_469;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_553;
wire n_257;
wire n_61;
wire n_173;
wire n_561;
wire n_244;
wire n_232;
wire n_527;
wire n_482;
wire n_58;
wire n_41;
wire n_266;
wire n_548;
wire n_72;
wire n_512;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_516;
wire n_183;
wire n_409;
wire n_532;
wire n_249;
wire n_412;
wire n_217;
wire n_471;
wire n_541;
wire n_53;
wire n_372;
wire n_558;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_535;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_556;
wire n_524;
wire n_402;
wire n_563;
wire n_504;
wire n_438;
wire n_475;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_514;
wire n_564;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_0),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_15),
.Y(n_20)
);

BUFx5_ASAP7_75t_L g21 ( 
.A(n_17),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_12),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_18),
.Y(n_23)
);

INVx6_ASAP7_75t_L g24 ( 
.A(n_3),
.Y(n_24)
);

BUFx3_ASAP7_75t_L g25 ( 
.A(n_13),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_13),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_13),
.Y(n_27)
);

BUFx4f_ASAP7_75t_L g28 ( 
.A(n_11),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_8),
.Y(n_29)
);

INVxp33_ASAP7_75t_L g30 ( 
.A(n_10),
.Y(n_30)
);

BUFx3_ASAP7_75t_L g31 ( 
.A(n_1),
.Y(n_31)
);

INVx11_ASAP7_75t_SL g32 ( 
.A(n_1),
.Y(n_32)
);

INVx5_ASAP7_75t_L g33 ( 
.A(n_1),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_0),
.Y(n_34)
);

BUFx5_ASAP7_75t_L g35 ( 
.A(n_13),
.Y(n_35)
);

BUFx10_ASAP7_75t_L g36 ( 
.A(n_1),
.Y(n_36)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_3),
.Y(n_37)
);

BUFx3_ASAP7_75t_L g38 ( 
.A(n_17),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_4),
.Y(n_39)
);

BUFx12f_ASAP7_75t_L g40 ( 
.A(n_10),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g41 ( 
.A(n_3),
.B(n_17),
.Y(n_41)
);

INVx3_ASAP7_75t_L g42 ( 
.A(n_5),
.Y(n_42)
);

INVx6_ASAP7_75t_L g43 ( 
.A(n_18),
.Y(n_43)
);

INVx8_ASAP7_75t_L g44 ( 
.A(n_0),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_0),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_3),
.Y(n_46)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_7),
.Y(n_47)
);

BUFx3_ASAP7_75t_L g48 ( 
.A(n_15),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g49 ( 
.A(n_7),
.B(n_6),
.Y(n_49)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_14),
.Y(n_50)
);

BUFx3_ASAP7_75t_L g51 ( 
.A(n_8),
.Y(n_51)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_7),
.Y(n_52)
);

BUFx3_ASAP7_75t_L g53 ( 
.A(n_35),
.Y(n_53)
);

INVx5_ASAP7_75t_L g116 ( 
.A(n_53),
.Y(n_116)
);

INVx3_ASAP7_75t_L g54 ( 
.A(n_21),
.Y(n_54)
);

INVx3_ASAP7_75t_L g127 ( 
.A(n_54),
.Y(n_127)
);

BUFx4f_ASAP7_75t_SL g55 ( 
.A(n_21),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g118 ( 
.A(n_55),
.Y(n_118)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_19),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g137 ( 
.A(n_56),
.Y(n_137)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_20),
.Y(n_57)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_57),
.Y(n_129)
);

INVx6_ASAP7_75t_L g58 ( 
.A(n_19),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g138 ( 
.A(n_58),
.Y(n_138)
);

INVx2_ASAP7_75t_L g59 ( 
.A(n_28),
.Y(n_59)
);

INVx2_ASAP7_75t_L g110 ( 
.A(n_59),
.Y(n_110)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_28),
.Y(n_60)
);

INVx2_ASAP7_75t_L g113 ( 
.A(n_60),
.Y(n_113)
);

BUFx3_ASAP7_75t_L g61 ( 
.A(n_35),
.Y(n_61)
);

INVx5_ASAP7_75t_L g122 ( 
.A(n_61),
.Y(n_122)
);

HB1xp67_ASAP7_75t_L g62 ( 
.A(n_42),
.Y(n_62)
);

HB1xp67_ASAP7_75t_L g141 ( 
.A(n_62),
.Y(n_141)
);

INVx4_ASAP7_75t_SL g63 ( 
.A(n_36),
.Y(n_63)
);

INVx2_ASAP7_75t_SL g145 ( 
.A(n_63),
.Y(n_145)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_19),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g142 ( 
.A(n_64),
.Y(n_142)
);

INVx11_ASAP7_75t_L g65 ( 
.A(n_36),
.Y(n_65)
);

INVx8_ASAP7_75t_L g119 ( 
.A(n_65),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_41),
.B(n_18),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_SL g135 ( 
.A(n_66),
.B(n_78),
.Y(n_135)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_27),
.Y(n_67)
);

BUFx6f_ASAP7_75t_L g159 ( 
.A(n_67),
.Y(n_159)
);

INVx2_ASAP7_75t_L g68 ( 
.A(n_28),
.Y(n_68)
);

INVx2_ASAP7_75t_L g123 ( 
.A(n_68),
.Y(n_123)
);

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_27),
.Y(n_69)
);

BUFx6f_ASAP7_75t_L g163 ( 
.A(n_69),
.Y(n_163)
);

BUFx6f_ASAP7_75t_L g70 ( 
.A(n_27),
.Y(n_70)
);

INVx6_ASAP7_75t_L g108 ( 
.A(n_70),
.Y(n_108)
);

BUFx12f_ASAP7_75t_L g71 ( 
.A(n_21),
.Y(n_71)
);

INVx4_ASAP7_75t_L g109 ( 
.A(n_71),
.Y(n_109)
);

INVx3_ASAP7_75t_SL g72 ( 
.A(n_36),
.Y(n_72)
);

INVx2_ASAP7_75t_L g125 ( 
.A(n_72),
.Y(n_125)
);

INVx11_ASAP7_75t_L g73 ( 
.A(n_36),
.Y(n_73)
);

INVx8_ASAP7_75t_L g161 ( 
.A(n_73),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_L g74 ( 
.A(n_41),
.B(n_16),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_L g120 ( 
.A(n_74),
.B(n_91),
.Y(n_120)
);

INVx8_ASAP7_75t_L g75 ( 
.A(n_29),
.Y(n_75)
);

BUFx2_ASAP7_75t_L g131 ( 
.A(n_75),
.Y(n_131)
);

BUFx6f_ASAP7_75t_L g76 ( 
.A(n_29),
.Y(n_76)
);

INVx6_ASAP7_75t_L g156 ( 
.A(n_76),
.Y(n_156)
);

INVx11_ASAP7_75t_L g77 ( 
.A(n_36),
.Y(n_77)
);

INVxp67_ASAP7_75t_L g146 ( 
.A(n_77),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_49),
.B(n_2),
.Y(n_78)
);

BUFx6f_ASAP7_75t_L g79 ( 
.A(n_29),
.Y(n_79)
);

INVx4_ASAP7_75t_L g126 ( 
.A(n_79),
.Y(n_126)
);

BUFx12f_ASAP7_75t_L g80 ( 
.A(n_25),
.Y(n_80)
);

INVx4_ASAP7_75t_L g134 ( 
.A(n_80),
.Y(n_134)
);

BUFx5_ASAP7_75t_L g81 ( 
.A(n_46),
.Y(n_81)
);

INVx4_ASAP7_75t_L g164 ( 
.A(n_81),
.Y(n_164)
);

INVx3_ASAP7_75t_L g82 ( 
.A(n_25),
.Y(n_82)
);

INVx3_ASAP7_75t_L g157 ( 
.A(n_82),
.Y(n_157)
);

INVx3_ASAP7_75t_L g83 ( 
.A(n_38),
.Y(n_83)
);

INVx3_ASAP7_75t_L g115 ( 
.A(n_83),
.Y(n_115)
);

AND2x2_ASAP7_75t_L g84 ( 
.A(n_49),
.B(n_2),
.Y(n_84)
);

AOI21xp33_ASAP7_75t_L g128 ( 
.A1(n_84),
.A2(n_52),
.B(n_50),
.Y(n_128)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_20),
.Y(n_85)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_85),
.Y(n_154)
);

BUFx3_ASAP7_75t_L g86 ( 
.A(n_40),
.Y(n_86)
);

INVx3_ASAP7_75t_L g117 ( 
.A(n_86),
.Y(n_117)
);

BUFx6f_ASAP7_75t_L g87 ( 
.A(n_46),
.Y(n_87)
);

INVx3_ASAP7_75t_L g130 ( 
.A(n_87),
.Y(n_130)
);

BUFx6f_ASAP7_75t_L g88 ( 
.A(n_46),
.Y(n_88)
);

INVx3_ASAP7_75t_L g155 ( 
.A(n_88),
.Y(n_155)
);

BUFx3_ASAP7_75t_L g89 ( 
.A(n_40),
.Y(n_89)
);

INVx2_ASAP7_75t_L g139 ( 
.A(n_89),
.Y(n_139)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_22),
.Y(n_90)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_90),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_SL g91 ( 
.A(n_38),
.B(n_39),
.Y(n_91)
);

INVx2_ASAP7_75t_L g92 ( 
.A(n_28),
.Y(n_92)
);

INVx2_ASAP7_75t_L g143 ( 
.A(n_92),
.Y(n_143)
);

INVx6_ASAP7_75t_L g93 ( 
.A(n_24),
.Y(n_93)
);

INVx2_ASAP7_75t_L g144 ( 
.A(n_93),
.Y(n_144)
);

INVx3_ASAP7_75t_L g94 ( 
.A(n_38),
.Y(n_94)
);

INVx2_ASAP7_75t_L g172 ( 
.A(n_94),
.Y(n_172)
);

INVx3_ASAP7_75t_L g95 ( 
.A(n_25),
.Y(n_95)
);

INVx2_ASAP7_75t_L g147 ( 
.A(n_95),
.Y(n_147)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_22),
.Y(n_96)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_96),
.Y(n_168)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_30),
.B(n_2),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_SL g152 ( 
.A(n_97),
.B(n_33),
.Y(n_152)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_26),
.Y(n_98)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_98),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_39),
.B(n_16),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g124 ( 
.A(n_99),
.B(n_106),
.Y(n_124)
);

OR2x2_ASAP7_75t_L g100 ( 
.A(n_26),
.B(n_2),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g112 ( 
.A(n_100),
.B(n_104),
.Y(n_112)
);

INVx4_ASAP7_75t_L g101 ( 
.A(n_40),
.Y(n_101)
);

INVx2_ASAP7_75t_L g148 ( 
.A(n_101),
.Y(n_148)
);

BUFx6f_ASAP7_75t_L g102 ( 
.A(n_44),
.Y(n_102)
);

INVx2_ASAP7_75t_L g150 ( 
.A(n_102),
.Y(n_150)
);

INVx6_ASAP7_75t_L g103 ( 
.A(n_24),
.Y(n_103)
);

INVx2_ASAP7_75t_L g160 ( 
.A(n_103),
.Y(n_160)
);

CKINVDCx20_ASAP7_75t_R g104 ( 
.A(n_32),
.Y(n_104)
);

BUFx3_ASAP7_75t_L g105 ( 
.A(n_40),
.Y(n_105)
);

INVx2_ASAP7_75t_L g162 ( 
.A(n_105),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_L g106 ( 
.A(n_45),
.B(n_4),
.Y(n_106)
);

BUFx6f_ASAP7_75t_L g107 ( 
.A(n_44),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_L g132 ( 
.A(n_107),
.B(n_44),
.Y(n_132)
);

CKINVDCx20_ASAP7_75t_R g111 ( 
.A(n_100),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_L g180 ( 
.A(n_111),
.B(n_136),
.Y(n_180)
);

NOR2xp33_ASAP7_75t_L g114 ( 
.A(n_84),
.B(n_45),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_SL g199 ( 
.A(n_114),
.B(n_121),
.Y(n_199)
);

NOR2xp33_ASAP7_75t_L g121 ( 
.A(n_55),
.B(n_71),
.Y(n_121)
);

AND2x2_ASAP7_75t_L g179 ( 
.A(n_128),
.B(n_132),
.Y(n_179)
);

NOR2xp33_ASAP7_75t_L g133 ( 
.A(n_55),
.B(n_52),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_SL g218 ( 
.A(n_133),
.B(n_140),
.Y(n_218)
);

CKINVDCx20_ASAP7_75t_R g136 ( 
.A(n_65),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_L g140 ( 
.A(n_71),
.B(n_50),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_L g149 ( 
.A(n_101),
.B(n_34),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_L g194 ( 
.A(n_149),
.B(n_153),
.Y(n_194)
);

AOI22xp33_ASAP7_75t_SL g151 ( 
.A1(n_53),
.A2(n_42),
.B1(n_33),
.B2(n_31),
.Y(n_151)
);

AOI22xp33_ASAP7_75t_SL g184 ( 
.A1(n_151),
.A2(n_61),
.B1(n_75),
.B2(n_89),
.Y(n_184)
);

AND2x2_ASAP7_75t_L g192 ( 
.A(n_152),
.B(n_63),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_SL g153 ( 
.A(n_82),
.B(n_47),
.Y(n_153)
);

OAI22xp33_ASAP7_75t_L g158 ( 
.A1(n_58),
.A2(n_24),
.B1(n_42),
.B2(n_43),
.Y(n_158)
);

OAI22xp5_ASAP7_75t_SL g183 ( 
.A1(n_158),
.A2(n_167),
.B1(n_69),
.B2(n_56),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_L g165 ( 
.A(n_93),
.B(n_37),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_L g196 ( 
.A(n_165),
.B(n_169),
.Y(n_196)
);

OAI22xp5_ASAP7_75t_L g167 ( 
.A1(n_103),
.A2(n_43),
.B1(n_23),
.B2(n_51),
.Y(n_167)
);

NOR2xp33_ASAP7_75t_L g169 ( 
.A(n_80),
.B(n_37),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_SL g170 ( 
.A(n_80),
.B(n_34),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_L g200 ( 
.A(n_170),
.B(n_86),
.Y(n_200)
);

INVx3_ASAP7_75t_L g173 ( 
.A(n_118),
.Y(n_173)
);

INVx3_ASAP7_75t_L g279 ( 
.A(n_173),
.Y(n_279)
);

BUFx3_ASAP7_75t_L g174 ( 
.A(n_118),
.Y(n_174)
);

INVx5_ASAP7_75t_L g277 ( 
.A(n_174),
.Y(n_277)
);

INVx5_ASAP7_75t_L g175 ( 
.A(n_134),
.Y(n_175)
);

INVx3_ASAP7_75t_L g287 ( 
.A(n_175),
.Y(n_287)
);

INVx5_ASAP7_75t_L g176 ( 
.A(n_134),
.Y(n_176)
);

BUFx6f_ASAP7_75t_L g273 ( 
.A(n_176),
.Y(n_273)
);

INVx2_ASAP7_75t_L g177 ( 
.A(n_110),
.Y(n_177)
);

INVx2_ASAP7_75t_L g256 ( 
.A(n_177),
.Y(n_256)
);

MAJIxp5_ASAP7_75t_L g178 ( 
.A(n_129),
.B(n_72),
.C(n_77),
.Y(n_178)
);

AND2x2_ASAP7_75t_L g260 ( 
.A(n_178),
.B(n_192),
.Y(n_260)
);

OR2x2_ASAP7_75t_L g181 ( 
.A(n_124),
.B(n_47),
.Y(n_181)
);

NOR2xp33_ASAP7_75t_L g251 ( 
.A(n_181),
.B(n_182),
.Y(n_251)
);

CKINVDCx20_ASAP7_75t_R g182 ( 
.A(n_141),
.Y(n_182)
);

AOI22xp5_ASAP7_75t_L g280 ( 
.A1(n_183),
.A2(n_195),
.B1(n_9),
.B2(n_10),
.Y(n_280)
);

INVxp67_ASAP7_75t_L g262 ( 
.A(n_184),
.Y(n_262)
);

INVx2_ASAP7_75t_L g185 ( 
.A(n_113),
.Y(n_185)
);

INVx2_ASAP7_75t_L g285 ( 
.A(n_185),
.Y(n_285)
);

BUFx6f_ASAP7_75t_L g186 ( 
.A(n_137),
.Y(n_186)
);

INVx6_ASAP7_75t_L g247 ( 
.A(n_186),
.Y(n_247)
);

BUFx2_ASAP7_75t_L g187 ( 
.A(n_116),
.Y(n_187)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_187),
.Y(n_254)
);

INVx2_ASAP7_75t_SL g188 ( 
.A(n_117),
.Y(n_188)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_188),
.Y(n_264)
);

INVx4_ASAP7_75t_L g189 ( 
.A(n_117),
.Y(n_189)
);

INVx6_ASAP7_75t_L g259 ( 
.A(n_189),
.Y(n_259)
);

INVx2_ASAP7_75t_L g190 ( 
.A(n_123),
.Y(n_190)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_190),
.Y(n_268)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_154),
.Y(n_191)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_191),
.Y(n_272)
);

BUFx6f_ASAP7_75t_L g193 ( 
.A(n_137),
.Y(n_193)
);

INVx8_ASAP7_75t_L g240 ( 
.A(n_193),
.Y(n_240)
);

OAI22xp5_ASAP7_75t_SL g195 ( 
.A1(n_151),
.A2(n_70),
.B1(n_64),
.B2(n_67),
.Y(n_195)
);

NOR2xp33_ASAP7_75t_L g197 ( 
.A(n_112),
.B(n_105),
.Y(n_197)
);

NOR2xp33_ASAP7_75t_L g252 ( 
.A(n_197),
.B(n_200),
.Y(n_252)
);

INVx1_ASAP7_75t_SL g198 ( 
.A(n_125),
.Y(n_198)
);

AND2x2_ASAP7_75t_L g266 ( 
.A(n_198),
.B(n_211),
.Y(n_266)
);

AND2x2_ASAP7_75t_L g201 ( 
.A(n_120),
.B(n_73),
.Y(n_201)
);

CKINVDCx14_ASAP7_75t_R g286 ( 
.A(n_201),
.Y(n_286)
);

INVx3_ASAP7_75t_L g202 ( 
.A(n_116),
.Y(n_202)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_202),
.Y(n_275)
);

INVx3_ASAP7_75t_L g203 ( 
.A(n_122),
.Y(n_203)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_203),
.Y(n_288)
);

NAND2xp5_ASAP7_75t_L g204 ( 
.A(n_135),
.B(n_43),
.Y(n_204)
);

NOR2xp33_ASAP7_75t_L g261 ( 
.A(n_204),
.B(n_205),
.Y(n_261)
);

INVx2_ASAP7_75t_L g205 ( 
.A(n_143),
.Y(n_205)
);

INVx4_ASAP7_75t_L g206 ( 
.A(n_109),
.Y(n_206)
);

CKINVDCx16_ASAP7_75t_R g267 ( 
.A(n_206),
.Y(n_267)
);

A2O1A1Ixp33_ASAP7_75t_L g207 ( 
.A1(n_166),
.A2(n_40),
.B(n_48),
.C(n_31),
.Y(n_207)
);

A2O1A1Ixp33_ASAP7_75t_L g241 ( 
.A1(n_207),
.A2(n_161),
.B(n_126),
.C(n_155),
.Y(n_241)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_168),
.Y(n_208)
);

NOR2xp33_ASAP7_75t_L g265 ( 
.A(n_208),
.B(n_209),
.Y(n_265)
);

NAND2xp5_ASAP7_75t_L g209 ( 
.A(n_171),
.B(n_23),
.Y(n_209)
);

NOR2xp33_ASAP7_75t_L g210 ( 
.A(n_127),
.B(n_23),
.Y(n_210)
);

NOR2xp33_ASAP7_75t_L g281 ( 
.A(n_210),
.B(n_213),
.Y(n_281)
);

INVx2_ASAP7_75t_L g211 ( 
.A(n_144),
.Y(n_211)
);

AND2x2_ASAP7_75t_L g212 ( 
.A(n_145),
.B(n_33),
.Y(n_212)
);

AND2x2_ASAP7_75t_L g270 ( 
.A(n_212),
.B(n_217),
.Y(n_270)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_145),
.Y(n_213)
);

INVxp67_ASAP7_75t_L g214 ( 
.A(n_119),
.Y(n_214)
);

NOR2xp33_ASAP7_75t_L g284 ( 
.A(n_214),
.B(n_216),
.Y(n_284)
);

AOI21xp5_ASAP7_75t_L g215 ( 
.A1(n_146),
.A2(n_51),
.B(n_48),
.Y(n_215)
);

AOI21xp5_ASAP7_75t_L g239 ( 
.A1(n_215),
.A2(n_146),
.B(n_164),
.Y(n_239)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_172),
.Y(n_216)
);

INVx4_ASAP7_75t_L g217 ( 
.A(n_109),
.Y(n_217)
);

INVx2_ASAP7_75t_L g219 ( 
.A(n_160),
.Y(n_219)
);

AND2x2_ASAP7_75t_L g283 ( 
.A(n_219),
.B(n_221),
.Y(n_283)
);

AOI211xp5_ASAP7_75t_SL g220 ( 
.A1(n_158),
.A2(n_107),
.B(n_102),
.C(n_88),
.Y(n_220)
);

AOI22xp5_ASAP7_75t_SL g269 ( 
.A1(n_220),
.A2(n_225),
.B1(n_227),
.B2(n_233),
.Y(n_269)
);

AND2x2_ASAP7_75t_L g221 ( 
.A(n_148),
.B(n_51),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_L g222 ( 
.A(n_147),
.B(n_4),
.Y(n_222)
);

NAND2xp5_ASAP7_75t_L g236 ( 
.A(n_222),
.B(n_5),
.Y(n_236)
);

INVx2_ASAP7_75t_L g223 ( 
.A(n_157),
.Y(n_223)
);

INVx2_ASAP7_75t_R g238 ( 
.A(n_223),
.Y(n_238)
);

INVx2_ASAP7_75t_L g224 ( 
.A(n_130),
.Y(n_224)
);

CKINVDCx20_ASAP7_75t_R g244 ( 
.A(n_224),
.Y(n_244)
);

MAJIxp5_ASAP7_75t_L g225 ( 
.A(n_115),
.B(n_139),
.C(n_162),
.Y(n_225)
);

AOI22xp33_ASAP7_75t_SL g226 ( 
.A1(n_122),
.A2(n_48),
.B1(n_31),
.B2(n_76),
.Y(n_226)
);

AOI22xp33_ASAP7_75t_SL g237 ( 
.A1(n_226),
.A2(n_231),
.B1(n_234),
.B2(n_235),
.Y(n_237)
);

MAJIxp5_ASAP7_75t_L g227 ( 
.A(n_115),
.B(n_87),
.C(n_79),
.Y(n_227)
);

BUFx16f_ASAP7_75t_L g228 ( 
.A(n_131),
.Y(n_228)
);

CKINVDCx20_ASAP7_75t_R g258 ( 
.A(n_228),
.Y(n_258)
);

INVx2_ASAP7_75t_L g229 ( 
.A(n_130),
.Y(n_229)
);

CKINVDCx20_ASAP7_75t_R g282 ( 
.A(n_229),
.Y(n_282)
);

BUFx3_ASAP7_75t_L g230 ( 
.A(n_131),
.Y(n_230)
);

INVxp33_ASAP7_75t_L g250 ( 
.A(n_230),
.Y(n_250)
);

BUFx2_ASAP7_75t_L g231 ( 
.A(n_164),
.Y(n_231)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_150),
.Y(n_232)
);

OR2x2_ASAP7_75t_L g263 ( 
.A(n_232),
.B(n_6),
.Y(n_263)
);

AND2x2_ASAP7_75t_L g233 ( 
.A(n_119),
.B(n_4),
.Y(n_233)
);

BUFx6f_ASAP7_75t_L g234 ( 
.A(n_142),
.Y(n_234)
);

INVxp67_ASAP7_75t_L g235 ( 
.A(n_161),
.Y(n_235)
);

NAND2xp5_ASAP7_75t_SL g300 ( 
.A(n_236),
.B(n_271),
.Y(n_300)
);

OAI21xp5_ASAP7_75t_SL g313 ( 
.A1(n_239),
.A2(n_228),
.B(n_202),
.Y(n_313)
);

AOI21xp5_ASAP7_75t_L g293 ( 
.A1(n_241),
.A2(n_242),
.B(n_249),
.Y(n_293)
);

NAND2x1_ASAP7_75t_SL g242 ( 
.A(n_178),
.B(n_155),
.Y(n_242)
);

AOI22xp33_ASAP7_75t_SL g243 ( 
.A1(n_195),
.A2(n_126),
.B1(n_156),
.B2(n_108),
.Y(n_243)
);

INVxp67_ASAP7_75t_L g307 ( 
.A(n_243),
.Y(n_307)
);

NAND2xp5_ASAP7_75t_L g245 ( 
.A(n_194),
.B(n_156),
.Y(n_245)
);

NAND2xp5_ASAP7_75t_L g316 ( 
.A(n_245),
.B(n_248),
.Y(n_316)
);

OAI22xp5_ASAP7_75t_SL g246 ( 
.A1(n_184),
.A2(n_138),
.B1(n_108),
.B2(n_142),
.Y(n_246)
);

AOI22xp5_ASAP7_75t_L g299 ( 
.A1(n_246),
.A2(n_253),
.B1(n_255),
.B2(n_198),
.Y(n_299)
);

NAND2xp5_ASAP7_75t_L g248 ( 
.A(n_196),
.B(n_138),
.Y(n_248)
);

OAI21xp5_ASAP7_75t_L g249 ( 
.A1(n_179),
.A2(n_163),
.B(n_159),
.Y(n_249)
);

OAI22xp5_ASAP7_75t_L g253 ( 
.A1(n_220),
.A2(n_163),
.B1(n_159),
.B2(n_7),
.Y(n_253)
);

OAI22xp5_ASAP7_75t_SL g255 ( 
.A1(n_181),
.A2(n_5),
.B1(n_6),
.B2(n_8),
.Y(n_255)
);

AOI21xp5_ASAP7_75t_L g257 ( 
.A1(n_215),
.A2(n_5),
.B(n_6),
.Y(n_257)
);

AOI21xp5_ASAP7_75t_L g295 ( 
.A1(n_257),
.A2(n_207),
.B(n_233),
.Y(n_295)
);

INVxp67_ASAP7_75t_L g327 ( 
.A(n_263),
.Y(n_327)
);

NAND2xp5_ASAP7_75t_L g271 ( 
.A(n_179),
.B(n_201),
.Y(n_271)
);

NAND2xp5_ASAP7_75t_L g274 ( 
.A(n_218),
.B(n_8),
.Y(n_274)
);

NAND2xp5_ASAP7_75t_SL g301 ( 
.A(n_274),
.B(n_276),
.Y(n_301)
);

NAND2xp5_ASAP7_75t_L g276 ( 
.A(n_192),
.B(n_9),
.Y(n_276)
);

NAND2xp5_ASAP7_75t_L g278 ( 
.A(n_180),
.B(n_9),
.Y(n_278)
);

NAND2xp5_ASAP7_75t_SL g304 ( 
.A(n_278),
.B(n_9),
.Y(n_304)
);

OAI22xp5_ASAP7_75t_SL g292 ( 
.A1(n_280),
.A2(n_226),
.B1(n_234),
.B2(n_186),
.Y(n_292)
);

INVx2_ASAP7_75t_L g289 ( 
.A(n_264),
.Y(n_289)
);

INVx2_ASAP7_75t_L g359 ( 
.A(n_289),
.Y(n_359)
);

CKINVDCx20_ASAP7_75t_R g290 ( 
.A(n_266),
.Y(n_290)
);

NOR2xp33_ASAP7_75t_L g343 ( 
.A(n_290),
.B(n_308),
.Y(n_343)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_266),
.Y(n_291)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_291),
.Y(n_341)
);

AOI22xp5_ASAP7_75t_L g354 ( 
.A1(n_292),
.A2(n_320),
.B1(n_270),
.B2(n_283),
.Y(n_354)
);

NOR2xp33_ASAP7_75t_L g294 ( 
.A(n_265),
.B(n_199),
.Y(n_294)
);

NAND2xp5_ASAP7_75t_SL g346 ( 
.A(n_294),
.B(n_296),
.Y(n_346)
);

OAI21xp5_ASAP7_75t_SL g338 ( 
.A1(n_295),
.A2(n_305),
.B(n_257),
.Y(n_338)
);

NOR2xp33_ASAP7_75t_L g296 ( 
.A(n_274),
.B(n_225),
.Y(n_296)
);

AOI22xp33_ASAP7_75t_SL g297 ( 
.A1(n_262),
.A2(n_183),
.B1(n_187),
.B2(n_231),
.Y(n_297)
);

INVxp67_ASAP7_75t_L g350 ( 
.A(n_297),
.Y(n_350)
);

AND2x4_ASAP7_75t_SL g298 ( 
.A(n_242),
.B(n_211),
.Y(n_298)
);

AND2x2_ASAP7_75t_L g375 ( 
.A(n_298),
.B(n_303),
.Y(n_375)
);

OAI22xp5_ASAP7_75t_L g368 ( 
.A1(n_299),
.A2(n_310),
.B1(n_254),
.B2(n_244),
.Y(n_368)
);

XOR2xp5_ASAP7_75t_L g302 ( 
.A(n_271),
.B(n_221),
.Y(n_302)
);

MAJIxp5_ASAP7_75t_L g347 ( 
.A(n_302),
.B(n_321),
.C(n_325),
.Y(n_347)
);

AND2x2_ASAP7_75t_L g303 ( 
.A(n_260),
.B(n_212),
.Y(n_303)
);

NAND2xp5_ASAP7_75t_SL g371 ( 
.A(n_304),
.B(n_306),
.Y(n_371)
);

AOI22xp5_ASAP7_75t_SL g305 ( 
.A1(n_262),
.A2(n_286),
.B1(n_260),
.B2(n_246),
.Y(n_305)
);

NOR2xp33_ASAP7_75t_L g306 ( 
.A(n_248),
.B(n_188),
.Y(n_306)
);

CKINVDCx20_ASAP7_75t_R g308 ( 
.A(n_266),
.Y(n_308)
);

NAND2xp5_ASAP7_75t_SL g309 ( 
.A(n_261),
.B(n_227),
.Y(n_309)
);

NAND2xp5_ASAP7_75t_L g348 ( 
.A(n_309),
.B(n_312),
.Y(n_348)
);

AOI22xp5_ASAP7_75t_L g310 ( 
.A1(n_253),
.A2(n_224),
.B1(n_193),
.B2(n_189),
.Y(n_310)
);

AOI21xp5_ASAP7_75t_L g311 ( 
.A1(n_239),
.A2(n_235),
.B(n_214),
.Y(n_311)
);

AOI21xp5_ASAP7_75t_L g339 ( 
.A1(n_311),
.A2(n_313),
.B(n_249),
.Y(n_339)
);

NAND2xp5_ASAP7_75t_SL g312 ( 
.A(n_245),
.B(n_217),
.Y(n_312)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_264),
.Y(n_314)
);

INVx1_ASAP7_75t_L g342 ( 
.A(n_314),
.Y(n_342)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_272),
.Y(n_315)
);

INVx1_ASAP7_75t_L g345 ( 
.A(n_315),
.Y(n_345)
);

CKINVDCx20_ASAP7_75t_R g317 ( 
.A(n_284),
.Y(n_317)
);

NOR2xp33_ASAP7_75t_L g352 ( 
.A(n_317),
.B(n_326),
.Y(n_352)
);

OAI22xp33_ASAP7_75t_SL g318 ( 
.A1(n_269),
.A2(n_173),
.B1(n_203),
.B2(n_230),
.Y(n_318)
);

AOI22xp5_ASAP7_75t_SL g355 ( 
.A1(n_318),
.A2(n_283),
.B1(n_279),
.B2(n_288),
.Y(n_355)
);

HB1xp67_ASAP7_75t_L g319 ( 
.A(n_259),
.Y(n_319)
);

INVx1_ASAP7_75t_L g349 ( 
.A(n_319),
.Y(n_349)
);

OAI22xp5_ASAP7_75t_SL g320 ( 
.A1(n_269),
.A2(n_174),
.B1(n_206),
.B2(n_176),
.Y(n_320)
);

XOR2xp5_ASAP7_75t_L g321 ( 
.A(n_260),
.B(n_175),
.Y(n_321)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_272),
.Y(n_322)
);

INVx1_ASAP7_75t_L g351 ( 
.A(n_322),
.Y(n_351)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_268),
.Y(n_323)
);

INVx1_ASAP7_75t_L g366 ( 
.A(n_323),
.Y(n_366)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_268),
.Y(n_324)
);

INVx1_ASAP7_75t_L g376 ( 
.A(n_324),
.Y(n_376)
);

MAJIxp5_ASAP7_75t_L g325 ( 
.A(n_252),
.B(n_228),
.C(n_11),
.Y(n_325)
);

CKINVDCx20_ASAP7_75t_R g326 ( 
.A(n_281),
.Y(n_326)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_256),
.Y(n_328)
);

BUFx2_ASAP7_75t_L g367 ( 
.A(n_328),
.Y(n_367)
);

NAND2xp5_ASAP7_75t_SL g329 ( 
.A(n_236),
.B(n_10),
.Y(n_329)
);

NAND2xp5_ASAP7_75t_L g370 ( 
.A(n_329),
.B(n_330),
.Y(n_370)
);

NOR2xp33_ASAP7_75t_L g330 ( 
.A(n_251),
.B(n_11),
.Y(n_330)
);

INVx2_ASAP7_75t_L g331 ( 
.A(n_275),
.Y(n_331)
);

NAND2xp5_ASAP7_75t_L g372 ( 
.A(n_331),
.B(n_333),
.Y(n_372)
);

CKINVDCx20_ASAP7_75t_R g332 ( 
.A(n_270),
.Y(n_332)
);

NOR2xp33_ASAP7_75t_L g362 ( 
.A(n_332),
.B(n_336),
.Y(n_362)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_256),
.Y(n_333)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_285),
.Y(n_334)
);

NAND2xp5_ASAP7_75t_L g377 ( 
.A(n_334),
.B(n_335),
.Y(n_377)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_285),
.Y(n_335)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_275),
.Y(n_336)
);

OAI32xp33_ASAP7_75t_L g337 ( 
.A1(n_241),
.A2(n_11),
.A3(n_12),
.B1(n_14),
.B2(n_15),
.Y(n_337)
);

XOR2xp5_ASAP7_75t_L g340 ( 
.A(n_337),
.B(n_255),
.Y(n_340)
);

INVxp67_ASAP7_75t_L g409 ( 
.A(n_338),
.Y(n_409)
);

AOI21xp5_ASAP7_75t_L g386 ( 
.A1(n_339),
.A2(n_353),
.B(n_357),
.Y(n_386)
);

NAND2xp5_ASAP7_75t_SL g398 ( 
.A(n_340),
.B(n_325),
.Y(n_398)
);

OAI22xp5_ASAP7_75t_SL g344 ( 
.A1(n_293),
.A2(n_280),
.B1(n_242),
.B2(n_237),
.Y(n_344)
);

AOI22xp5_ASAP7_75t_L g387 ( 
.A1(n_344),
.A2(n_356),
.B1(n_368),
.B2(n_378),
.Y(n_387)
);

OAI21xp5_ASAP7_75t_SL g353 ( 
.A1(n_293),
.A2(n_270),
.B(n_276),
.Y(n_353)
);

OAI22xp33_ASAP7_75t_SL g393 ( 
.A1(n_354),
.A2(n_355),
.B1(n_307),
.B2(n_310),
.Y(n_393)
);

OAI22xp5_ASAP7_75t_SL g356 ( 
.A1(n_305),
.A2(n_263),
.B1(n_278),
.B2(n_288),
.Y(n_356)
);

AOI21xp5_ASAP7_75t_L g357 ( 
.A1(n_311),
.A2(n_263),
.B(n_258),
.Y(n_357)
);

MAJIxp5_ASAP7_75t_L g358 ( 
.A(n_321),
.B(n_283),
.C(n_282),
.Y(n_358)
);

MAJIxp5_ASAP7_75t_L g383 ( 
.A(n_358),
.B(n_363),
.C(n_373),
.Y(n_383)
);

AOI22xp5_ASAP7_75t_L g360 ( 
.A1(n_320),
.A2(n_279),
.B1(n_247),
.B2(n_240),
.Y(n_360)
);

OAI22xp5_ASAP7_75t_SL g394 ( 
.A1(n_360),
.A2(n_336),
.B1(n_314),
.B2(n_322),
.Y(n_394)
);

CKINVDCx20_ASAP7_75t_R g361 ( 
.A(n_312),
.Y(n_361)
);

NOR2xp33_ASAP7_75t_L g417 ( 
.A(n_361),
.B(n_365),
.Y(n_417)
);

XOR2xp5_ASAP7_75t_L g363 ( 
.A(n_302),
.B(n_254),
.Y(n_363)
);

AOI22xp33_ASAP7_75t_L g364 ( 
.A1(n_292),
.A2(n_240),
.B1(n_259),
.B2(n_244),
.Y(n_364)
);

INVxp67_ASAP7_75t_SL g412 ( 
.A(n_364),
.Y(n_412)
);

CKINVDCx20_ASAP7_75t_R g365 ( 
.A(n_306),
.Y(n_365)
);

CKINVDCx20_ASAP7_75t_R g369 ( 
.A(n_298),
.Y(n_369)
);

INVx13_ASAP7_75t_L g396 ( 
.A(n_369),
.Y(n_396)
);

XOR2xp5_ASAP7_75t_L g373 ( 
.A(n_296),
.B(n_282),
.Y(n_373)
);

BUFx24_ASAP7_75t_SL g374 ( 
.A(n_294),
.Y(n_374)
);

BUFx24_ASAP7_75t_SL g381 ( 
.A(n_374),
.Y(n_381)
);

OAI22xp5_ASAP7_75t_SL g378 ( 
.A1(n_299),
.A2(n_247),
.B1(n_267),
.B2(n_277),
.Y(n_378)
);

OAI21xp5_ASAP7_75t_L g379 ( 
.A1(n_295),
.A2(n_250),
.B(n_258),
.Y(n_379)
);

OAI21xp5_ASAP7_75t_L g389 ( 
.A1(n_379),
.A2(n_313),
.B(n_327),
.Y(n_389)
);

XOR2xp5_ASAP7_75t_L g380 ( 
.A(n_316),
.B(n_238),
.Y(n_380)
);

MAJIxp5_ASAP7_75t_L g392 ( 
.A(n_380),
.B(n_347),
.C(n_303),
.Y(n_392)
);

NAND2xp5_ASAP7_75t_L g382 ( 
.A(n_365),
.B(n_316),
.Y(n_382)
);

NAND2xp5_ASAP7_75t_L g427 ( 
.A(n_382),
.B(n_384),
.Y(n_427)
);

NAND2xp5_ASAP7_75t_L g384 ( 
.A(n_361),
.B(n_300),
.Y(n_384)
);

INVx1_ASAP7_75t_L g385 ( 
.A(n_377),
.Y(n_385)
);

INVx1_ASAP7_75t_L g424 ( 
.A(n_385),
.Y(n_424)
);

HB1xp67_ASAP7_75t_L g388 ( 
.A(n_349),
.Y(n_388)
);

INVx1_ASAP7_75t_L g425 ( 
.A(n_388),
.Y(n_425)
);

OAI21xp5_ASAP7_75t_L g418 ( 
.A1(n_389),
.A2(n_399),
.B(n_414),
.Y(n_418)
);

XNOR2x1_ASAP7_75t_L g390 ( 
.A(n_347),
.B(n_298),
.Y(n_390)
);

XNOR2xp5_ASAP7_75t_SL g426 ( 
.A(n_390),
.B(n_375),
.Y(n_426)
);

CKINVDCx14_ASAP7_75t_R g391 ( 
.A(n_352),
.Y(n_391)
);

CKINVDCx14_ASAP7_75t_R g445 ( 
.A(n_391),
.Y(n_445)
);

XOR2xp5_ASAP7_75t_L g441 ( 
.A(n_392),
.B(n_345),
.Y(n_441)
);

AOI22xp5_ASAP7_75t_L g420 ( 
.A1(n_393),
.A2(n_394),
.B1(n_397),
.B2(n_415),
.Y(n_420)
);

AOI22xp5_ASAP7_75t_L g395 ( 
.A1(n_344),
.A2(n_303),
.B1(n_298),
.B2(n_332),
.Y(n_395)
);

OAI22xp5_ASAP7_75t_L g428 ( 
.A1(n_395),
.A2(n_343),
.B1(n_341),
.B2(n_375),
.Y(n_428)
);

OAI22xp5_ASAP7_75t_SL g397 ( 
.A1(n_354),
.A2(n_309),
.B1(n_300),
.B2(n_308),
.Y(n_397)
);

OAI21x1_ASAP7_75t_SL g435 ( 
.A1(n_398),
.A2(n_413),
.B(n_370),
.Y(n_435)
);

AOI21xp5_ASAP7_75t_L g399 ( 
.A1(n_339),
.A2(n_290),
.B(n_291),
.Y(n_399)
);

INVx1_ASAP7_75t_L g400 ( 
.A(n_377),
.Y(n_400)
);

INVx1_ASAP7_75t_L g432 ( 
.A(n_400),
.Y(n_432)
);

INVx1_ASAP7_75t_L g401 ( 
.A(n_342),
.Y(n_401)
);

INVx1_ASAP7_75t_L g442 ( 
.A(n_401),
.Y(n_442)
);

INVx1_ASAP7_75t_L g402 ( 
.A(n_342),
.Y(n_402)
);

INVx2_ASAP7_75t_L g449 ( 
.A(n_402),
.Y(n_449)
);

INVx1_ASAP7_75t_L g403 ( 
.A(n_372),
.Y(n_403)
);

INVxp67_ASAP7_75t_L g429 ( 
.A(n_403),
.Y(n_429)
);

INVx2_ASAP7_75t_L g404 ( 
.A(n_359),
.Y(n_404)
);

NOR2xp33_ASAP7_75t_L g439 ( 
.A(n_404),
.B(n_411),
.Y(n_439)
);

OA22x2_ASAP7_75t_L g405 ( 
.A1(n_369),
.A2(n_337),
.B1(n_317),
.B2(n_289),
.Y(n_405)
);

AO22x2_ASAP7_75t_L g422 ( 
.A1(n_405),
.A2(n_341),
.B1(n_355),
.B2(n_368),
.Y(n_422)
);

MAJIxp5_ASAP7_75t_L g406 ( 
.A(n_363),
.B(n_326),
.C(n_301),
.Y(n_406)
);

MAJIxp5_ASAP7_75t_L g419 ( 
.A(n_406),
.B(n_373),
.C(n_358),
.Y(n_419)
);

CKINVDCx16_ASAP7_75t_R g407 ( 
.A(n_362),
.Y(n_407)
);

NAND2xp5_ASAP7_75t_SL g440 ( 
.A(n_407),
.B(n_349),
.Y(n_440)
);

OAI21xp5_ASAP7_75t_L g408 ( 
.A1(n_357),
.A2(n_330),
.B(n_324),
.Y(n_408)
);

AOI21xp5_ASAP7_75t_L g434 ( 
.A1(n_408),
.A2(n_353),
.B(n_371),
.Y(n_434)
);

NOR2xp33_ASAP7_75t_SL g410 ( 
.A(n_370),
.B(n_346),
.Y(n_410)
);

NOR2xp33_ASAP7_75t_SL g437 ( 
.A(n_410),
.B(n_351),
.Y(n_437)
);

INVx2_ASAP7_75t_L g411 ( 
.A(n_359),
.Y(n_411)
);

NAND2xp5_ASAP7_75t_L g413 ( 
.A(n_372),
.B(n_329),
.Y(n_413)
);

AOI21xp5_ASAP7_75t_L g414 ( 
.A1(n_379),
.A2(n_315),
.B(n_331),
.Y(n_414)
);

OAI22xp5_ASAP7_75t_SL g415 ( 
.A1(n_348),
.A2(n_301),
.B1(n_323),
.B2(n_304),
.Y(n_415)
);

AOI21xp5_ASAP7_75t_L g416 ( 
.A1(n_338),
.A2(n_287),
.B(n_277),
.Y(n_416)
);

OAI21xp5_ASAP7_75t_L g421 ( 
.A1(n_416),
.A2(n_350),
.B(n_375),
.Y(n_421)
);

MAJIxp5_ASAP7_75t_L g452 ( 
.A(n_419),
.B(n_441),
.C(n_443),
.Y(n_452)
);

INVxp67_ASAP7_75t_L g453 ( 
.A(n_421),
.Y(n_453)
);

INVx1_ASAP7_75t_SL g476 ( 
.A(n_422),
.Y(n_476)
);

AOI22xp5_ASAP7_75t_L g423 ( 
.A1(n_397),
.A2(n_350),
.B1(n_378),
.B2(n_340),
.Y(n_423)
);

OAI22xp5_ASAP7_75t_SL g454 ( 
.A1(n_423),
.A2(n_430),
.B1(n_433),
.B2(n_416),
.Y(n_454)
);

XNOR2xp5_ASAP7_75t_SL g470 ( 
.A(n_426),
.B(n_435),
.Y(n_470)
);

AOI22xp5_ASAP7_75t_L g463 ( 
.A1(n_428),
.A2(n_438),
.B1(n_446),
.B2(n_450),
.Y(n_463)
);

AOI22xp5_ASAP7_75t_L g430 ( 
.A1(n_385),
.A2(n_400),
.B1(n_403),
.B2(n_412),
.Y(n_430)
);

XNOR2xp5_ASAP7_75t_L g431 ( 
.A(n_383),
.B(n_392),
.Y(n_431)
);

XOR2xp5_ASAP7_75t_L g461 ( 
.A(n_431),
.B(n_436),
.Y(n_461)
);

AOI22xp5_ASAP7_75t_L g433 ( 
.A1(n_409),
.A2(n_348),
.B1(n_356),
.B2(n_380),
.Y(n_433)
);

OAI21xp5_ASAP7_75t_SL g466 ( 
.A1(n_434),
.A2(n_409),
.B(n_384),
.Y(n_466)
);

XNOR2xp5_ASAP7_75t_SL g436 ( 
.A(n_383),
.B(n_351),
.Y(n_436)
);

NOR2xp33_ASAP7_75t_SL g462 ( 
.A(n_437),
.B(n_407),
.Y(n_462)
);

OAI22xp5_ASAP7_75t_SL g438 ( 
.A1(n_387),
.A2(n_360),
.B1(n_345),
.B2(n_376),
.Y(n_438)
);

INVx1_ASAP7_75t_L g455 ( 
.A(n_440),
.Y(n_455)
);

XNOR2xp5_ASAP7_75t_L g443 ( 
.A(n_390),
.B(n_376),
.Y(n_443)
);

NOR2x1p5_ASAP7_75t_SL g444 ( 
.A(n_395),
.B(n_366),
.Y(n_444)
);

NAND2xp5_ASAP7_75t_L g451 ( 
.A(n_444),
.B(n_414),
.Y(n_451)
);

OAI22xp5_ASAP7_75t_SL g446 ( 
.A1(n_387),
.A2(n_366),
.B1(n_367),
.B2(n_335),
.Y(n_446)
);

XNOR2xp5_ASAP7_75t_SL g447 ( 
.A(n_406),
.B(n_334),
.Y(n_447)
);

MAJIxp5_ASAP7_75t_L g478 ( 
.A(n_447),
.B(n_448),
.C(n_401),
.Y(n_478)
);

MAJIxp5_ASAP7_75t_L g448 ( 
.A(n_399),
.B(n_333),
.C(n_328),
.Y(n_448)
);

OAI22xp5_ASAP7_75t_SL g450 ( 
.A1(n_386),
.A2(n_367),
.B1(n_273),
.B2(n_287),
.Y(n_450)
);

NAND2xp5_ASAP7_75t_L g487 ( 
.A(n_451),
.B(n_456),
.Y(n_487)
);

AOI22xp5_ASAP7_75t_L g481 ( 
.A1(n_454),
.A2(n_474),
.B1(n_479),
.B2(n_446),
.Y(n_481)
);

AO22x2_ASAP7_75t_L g456 ( 
.A1(n_418),
.A2(n_389),
.B1(n_386),
.B2(n_408),
.Y(n_456)
);

INVx1_ASAP7_75t_L g457 ( 
.A(n_449),
.Y(n_457)
);

INVx1_ASAP7_75t_L g485 ( 
.A(n_457),
.Y(n_485)
);

INVx1_ASAP7_75t_L g458 ( 
.A(n_442),
.Y(n_458)
);

INVx1_ASAP7_75t_L g497 ( 
.A(n_458),
.Y(n_497)
);

CKINVDCx20_ASAP7_75t_R g459 ( 
.A(n_439),
.Y(n_459)
);

NAND2xp5_ASAP7_75t_L g489 ( 
.A(n_459),
.B(n_460),
.Y(n_489)
);

INVx1_ASAP7_75t_L g460 ( 
.A(n_430),
.Y(n_460)
);

OAI22xp5_ASAP7_75t_L g491 ( 
.A1(n_462),
.A2(n_469),
.B1(n_472),
.B2(n_473),
.Y(n_491)
);

INVx1_ASAP7_75t_L g464 ( 
.A(n_427),
.Y(n_464)
);

NAND2xp5_ASAP7_75t_L g500 ( 
.A(n_464),
.B(n_467),
.Y(n_500)
);

AND2x2_ASAP7_75t_L g465 ( 
.A(n_421),
.B(n_417),
.Y(n_465)
);

NAND2x1_ASAP7_75t_L g493 ( 
.A(n_465),
.B(n_471),
.Y(n_493)
);

AOI21xp5_ASAP7_75t_L g490 ( 
.A1(n_466),
.A2(n_475),
.B(n_477),
.Y(n_490)
);

INVx1_ASAP7_75t_L g467 ( 
.A(n_424),
.Y(n_467)
);

NAND2xp5_ASAP7_75t_L g468 ( 
.A(n_429),
.B(n_382),
.Y(n_468)
);

CKINVDCx20_ASAP7_75t_R g494 ( 
.A(n_468),
.Y(n_494)
);

INVx1_ASAP7_75t_L g469 ( 
.A(n_425),
.Y(n_469)
);

NAND2xp5_ASAP7_75t_L g471 ( 
.A(n_429),
.B(n_413),
.Y(n_471)
);

AOI22xp5_ASAP7_75t_L g472 ( 
.A1(n_438),
.A2(n_394),
.B1(n_415),
.B2(n_410),
.Y(n_472)
);

INVx1_ASAP7_75t_L g473 ( 
.A(n_432),
.Y(n_473)
);

INVx8_ASAP7_75t_L g474 ( 
.A(n_445),
.Y(n_474)
);

CKINVDCx20_ASAP7_75t_R g475 ( 
.A(n_448),
.Y(n_475)
);

AND2x2_ASAP7_75t_L g477 ( 
.A(n_418),
.B(n_405),
.Y(n_477)
);

XNOR2xp5_ASAP7_75t_SL g488 ( 
.A(n_478),
.B(n_436),
.Y(n_488)
);

CKINVDCx20_ASAP7_75t_R g479 ( 
.A(n_450),
.Y(n_479)
);

MAJIxp5_ASAP7_75t_L g480 ( 
.A(n_452),
.B(n_441),
.C(n_431),
.Y(n_480)
);

MAJIxp5_ASAP7_75t_L g506 ( 
.A(n_480),
.B(n_492),
.C(n_496),
.Y(n_506)
);

INVx1_ASAP7_75t_L g505 ( 
.A(n_481),
.Y(n_505)
);

FAx1_ASAP7_75t_SL g482 ( 
.A(n_468),
.B(n_426),
.CI(n_433),
.CON(n_482),
.SN(n_482)
);

XNOR2xp5_ASAP7_75t_L g509 ( 
.A(n_482),
.B(n_501),
.Y(n_509)
);

AOI22xp5_ASAP7_75t_L g483 ( 
.A1(n_454),
.A2(n_444),
.B1(n_423),
.B2(n_422),
.Y(n_483)
);

OAI22xp5_ASAP7_75t_SL g518 ( 
.A1(n_483),
.A2(n_484),
.B1(n_486),
.B2(n_498),
.Y(n_518)
);

AOI22xp5_ASAP7_75t_L g484 ( 
.A1(n_476),
.A2(n_422),
.B1(n_420),
.B2(n_419),
.Y(n_484)
);

AOI22xp5_ASAP7_75t_L g486 ( 
.A1(n_476),
.A2(n_422),
.B1(n_420),
.B2(n_405),
.Y(n_486)
);

XNOR2xp5_ASAP7_75t_L g507 ( 
.A(n_488),
.B(n_466),
.Y(n_507)
);

MAJIxp5_ASAP7_75t_L g492 ( 
.A(n_452),
.B(n_447),
.C(n_443),
.Y(n_492)
);

XNOR2xp5_ASAP7_75t_SL g495 ( 
.A(n_470),
.B(n_396),
.Y(n_495)
);

XNOR2xp5_ASAP7_75t_SL g513 ( 
.A(n_495),
.B(n_499),
.Y(n_513)
);

MAJIxp5_ASAP7_75t_L g496 ( 
.A(n_461),
.B(n_405),
.C(n_396),
.Y(n_496)
);

AOI22xp5_ASAP7_75t_L g498 ( 
.A1(n_460),
.A2(n_402),
.B1(n_396),
.B2(n_411),
.Y(n_498)
);

XNOR2xp5_ASAP7_75t_SL g499 ( 
.A(n_470),
.B(n_367),
.Y(n_499)
);

XNOR2xp5_ASAP7_75t_SL g501 ( 
.A(n_461),
.B(n_238),
.Y(n_501)
);

MAJIxp5_ASAP7_75t_L g502 ( 
.A(n_478),
.B(n_404),
.C(n_273),
.Y(n_502)
);

MAJIxp5_ASAP7_75t_L g511 ( 
.A(n_502),
.B(n_480),
.C(n_496),
.Y(n_511)
);

AOI22xp5_ASAP7_75t_L g503 ( 
.A1(n_477),
.A2(n_273),
.B1(n_238),
.B2(n_381),
.Y(n_503)
);

XOR2xp5_ASAP7_75t_L g504 ( 
.A(n_503),
.B(n_472),
.Y(n_504)
);

XNOR2xp5_ASAP7_75t_L g526 ( 
.A(n_504),
.B(n_508),
.Y(n_526)
);

XOR2xp5_ASAP7_75t_L g538 ( 
.A(n_507),
.B(n_456),
.Y(n_538)
);

XOR2xp5_ASAP7_75t_L g508 ( 
.A(n_484),
.B(n_465),
.Y(n_508)
);

INVx6_ASAP7_75t_L g510 ( 
.A(n_491),
.Y(n_510)
);

INVx1_ASAP7_75t_L g533 ( 
.A(n_510),
.Y(n_533)
);

MAJIxp5_ASAP7_75t_L g524 ( 
.A(n_511),
.B(n_481),
.C(n_499),
.Y(n_524)
);

INVx1_ASAP7_75t_L g512 ( 
.A(n_500),
.Y(n_512)
);

NOR2xp33_ASAP7_75t_L g523 ( 
.A(n_512),
.B(n_517),
.Y(n_523)
);

XOR2xp5_ASAP7_75t_L g514 ( 
.A(n_492),
.B(n_465),
.Y(n_514)
);

XNOR2xp5_ASAP7_75t_L g529 ( 
.A(n_514),
.B(n_521),
.Y(n_529)
);

MAJIxp5_ASAP7_75t_L g515 ( 
.A(n_502),
.B(n_488),
.C(n_490),
.Y(n_515)
);

NAND2xp5_ASAP7_75t_SL g532 ( 
.A(n_515),
.B(n_516),
.Y(n_532)
);

XNOR2xp5_ASAP7_75t_L g516 ( 
.A(n_490),
.B(n_455),
.Y(n_516)
);

INVx11_ASAP7_75t_L g517 ( 
.A(n_494),
.Y(n_517)
);

AOI22xp5_ASAP7_75t_L g519 ( 
.A1(n_489),
.A2(n_464),
.B1(n_474),
.B2(n_467),
.Y(n_519)
);

OAI22xp5_ASAP7_75t_L g534 ( 
.A1(n_519),
.A2(n_463),
.B1(n_498),
.B2(n_471),
.Y(n_534)
);

XNOR2xp5_ASAP7_75t_L g520 ( 
.A(n_495),
.B(n_477),
.Y(n_520)
);

NOR2xp33_ASAP7_75t_SL g536 ( 
.A(n_520),
.B(n_522),
.Y(n_536)
);

XOR2xp5_ASAP7_75t_L g521 ( 
.A(n_501),
.B(n_453),
.Y(n_521)
);

INVx1_ASAP7_75t_L g522 ( 
.A(n_497),
.Y(n_522)
);

NAND2xp5_ASAP7_75t_L g545 ( 
.A(n_524),
.B(n_527),
.Y(n_545)
);

AOI21xp5_ASAP7_75t_L g525 ( 
.A1(n_517),
.A2(n_453),
.B(n_487),
.Y(n_525)
);

OAI21xp5_ASAP7_75t_SL g550 ( 
.A1(n_525),
.A2(n_533),
.B(n_524),
.Y(n_550)
);

OAI22xp5_ASAP7_75t_SL g527 ( 
.A1(n_505),
.A2(n_486),
.B1(n_483),
.B2(n_510),
.Y(n_527)
);

OAI21xp33_ASAP7_75t_L g528 ( 
.A1(n_507),
.A2(n_487),
.B(n_482),
.Y(n_528)
);

NOR3xp33_ASAP7_75t_L g549 ( 
.A(n_528),
.B(n_537),
.C(n_12),
.Y(n_549)
);

OAI22xp5_ASAP7_75t_SL g530 ( 
.A1(n_518),
.A2(n_463),
.B1(n_503),
.B2(n_451),
.Y(n_530)
);

XNOR2xp5_ASAP7_75t_L g542 ( 
.A(n_530),
.B(n_531),
.Y(n_542)
);

OAI21xp5_ASAP7_75t_SL g531 ( 
.A1(n_515),
.A2(n_493),
.B(n_456),
.Y(n_531)
);

XNOR2xp5_ASAP7_75t_L g543 ( 
.A(n_534),
.B(n_526),
.Y(n_543)
);

MAJIxp5_ASAP7_75t_L g535 ( 
.A(n_511),
.B(n_493),
.C(n_482),
.Y(n_535)
);

MAJIxp5_ASAP7_75t_L g539 ( 
.A(n_535),
.B(n_506),
.C(n_508),
.Y(n_539)
);

NOR2xp33_ASAP7_75t_SL g537 ( 
.A(n_514),
.B(n_485),
.Y(n_537)
);

XOR2xp5_ASAP7_75t_L g546 ( 
.A(n_538),
.B(n_513),
.Y(n_546)
);

AOI21xp5_ASAP7_75t_L g553 ( 
.A1(n_539),
.A2(n_540),
.B(n_541),
.Y(n_553)
);

NOR2xp33_ASAP7_75t_L g540 ( 
.A(n_536),
.B(n_504),
.Y(n_540)
);

MAJIxp5_ASAP7_75t_L g541 ( 
.A(n_526),
.B(n_506),
.C(n_513),
.Y(n_541)
);

XNOR2x1_ASAP7_75t_L g557 ( 
.A(n_543),
.B(n_546),
.Y(n_557)
);

NOR2xp33_ASAP7_75t_L g544 ( 
.A(n_532),
.B(n_458),
.Y(n_544)
);

NOR2xp33_ASAP7_75t_L g556 ( 
.A(n_544),
.B(n_547),
.Y(n_556)
);

OAI22xp5_ASAP7_75t_SL g547 ( 
.A1(n_533),
.A2(n_456),
.B1(n_509),
.B2(n_521),
.Y(n_547)
);

NOR2xp33_ASAP7_75t_SL g548 ( 
.A(n_523),
.B(n_535),
.Y(n_548)
);

NOR2x1_ASAP7_75t_L g555 ( 
.A(n_548),
.B(n_549),
.Y(n_555)
);

XNOR2xp5_ASAP7_75t_L g551 ( 
.A(n_550),
.B(n_531),
.Y(n_551)
);

INVx1_ASAP7_75t_L g562 ( 
.A(n_551),
.Y(n_562)
);

OAI22xp5_ASAP7_75t_SL g552 ( 
.A1(n_545),
.A2(n_525),
.B1(n_527),
.B2(n_530),
.Y(n_552)
);

INVxp33_ASAP7_75t_SL g560 ( 
.A(n_552),
.Y(n_560)
);

MAJIxp5_ASAP7_75t_L g554 ( 
.A(n_539),
.B(n_529),
.C(n_538),
.Y(n_554)
);

AND2x2_ASAP7_75t_L g559 ( 
.A(n_554),
.B(n_558),
.Y(n_559)
);

MAJIxp5_ASAP7_75t_L g558 ( 
.A(n_543),
.B(n_529),
.C(n_14),
.Y(n_558)
);

INVxp67_ASAP7_75t_L g561 ( 
.A(n_554),
.Y(n_561)
);

MAJIxp5_ASAP7_75t_L g565 ( 
.A(n_561),
.B(n_557),
.C(n_551),
.Y(n_565)
);

XNOR2xp5_ASAP7_75t_L g563 ( 
.A(n_557),
.B(n_541),
.Y(n_563)
);

AND2x2_ASAP7_75t_L g566 ( 
.A(n_563),
.B(n_542),
.Y(n_566)
);

OAI21xp5_ASAP7_75t_SL g564 ( 
.A1(n_562),
.A2(n_553),
.B(n_556),
.Y(n_564)
);

MAJIxp5_ASAP7_75t_L g567 ( 
.A(n_564),
.B(n_565),
.C(n_566),
.Y(n_567)
);

MAJIxp5_ASAP7_75t_L g568 ( 
.A(n_565),
.B(n_560),
.C(n_559),
.Y(n_568)
);

MAJIxp5_ASAP7_75t_L g569 ( 
.A(n_568),
.B(n_542),
.C(n_558),
.Y(n_569)
);

BUFx24_ASAP7_75t_SL g570 ( 
.A(n_569),
.Y(n_570)
);

MAJIxp5_ASAP7_75t_L g571 ( 
.A(n_570),
.B(n_567),
.C(n_555),
.Y(n_571)
);

MAJIxp5_ASAP7_75t_L g572 ( 
.A(n_571),
.B(n_555),
.C(n_546),
.Y(n_572)
);

AOI21xp5_ASAP7_75t_SL g573 ( 
.A1(n_572),
.A2(n_12),
.B(n_14),
.Y(n_573)
);

OA21x2_ASAP7_75t_L g574 ( 
.A1(n_573),
.A2(n_15),
.B(n_16),
.Y(n_574)
);


endmodule