module fake_netlist_6_4247_n_2152 (n_52, n_16, n_1, n_91, n_119, n_46, n_146, n_163, n_18, n_21, n_193, n_147, n_154, n_191, n_88, n_3, n_209, n_98, n_113, n_39, n_63, n_73, n_4, n_148, n_199, n_138, n_22, n_161, n_208, n_68, n_166, n_28, n_184, n_212, n_50, n_158, n_49, n_7, n_210, n_83, n_206, n_5, n_101, n_167, n_144, n_174, n_127, n_125, n_153, n_168, n_178, n_77, n_156, n_149, n_152, n_106, n_92, n_145, n_42, n_133, n_96, n_8, n_90, n_160, n_24, n_105, n_131, n_54, n_132, n_188, n_102, n_186, n_204, n_0, n_87, n_195, n_189, n_32, n_66, n_85, n_99, n_78, n_84, n_130, n_213, n_164, n_100, n_129, n_13, n_121, n_197, n_11, n_137, n_17, n_23, n_203, n_142, n_20, n_143, n_207, n_2, n_180, n_19, n_47, n_62, n_29, n_155, n_75, n_109, n_150, n_122, n_45, n_205, n_34, n_140, n_70, n_120, n_37, n_15, n_67, n_33, n_82, n_27, n_38, n_110, n_151, n_61, n_112, n_172, n_81, n_59, n_181, n_76, n_36, n_182, n_26, n_124, n_55, n_126, n_202, n_94, n_97, n_108, n_58, n_116, n_211, n_64, n_117, n_118, n_175, n_48, n_65, n_25, n_40, n_93, n_80, n_141, n_135, n_196, n_200, n_165, n_139, n_41, n_134, n_177, n_176, n_114, n_86, n_198, n_104, n_95, n_179, n_9, n_107, n_10, n_71, n_74, n_6, n_190, n_14, n_123, n_136, n_72, n_187, n_89, n_173, n_201, n_103, n_111, n_60, n_159, n_157, n_162, n_170, n_185, n_35, n_183, n_115, n_12, n_69, n_128, n_30, n_79, n_43, n_194, n_171, n_31, n_192, n_57, n_169, n_53, n_51, n_44, n_56, n_2152);

input n_52;
input n_16;
input n_1;
input n_91;
input n_119;
input n_46;
input n_146;
input n_163;
input n_18;
input n_21;
input n_193;
input n_147;
input n_154;
input n_191;
input n_88;
input n_3;
input n_209;
input n_98;
input n_113;
input n_39;
input n_63;
input n_73;
input n_4;
input n_148;
input n_199;
input n_138;
input n_22;
input n_161;
input n_208;
input n_68;
input n_166;
input n_28;
input n_184;
input n_212;
input n_50;
input n_158;
input n_49;
input n_7;
input n_210;
input n_83;
input n_206;
input n_5;
input n_101;
input n_167;
input n_144;
input n_174;
input n_127;
input n_125;
input n_153;
input n_168;
input n_178;
input n_77;
input n_156;
input n_149;
input n_152;
input n_106;
input n_92;
input n_145;
input n_42;
input n_133;
input n_96;
input n_8;
input n_90;
input n_160;
input n_24;
input n_105;
input n_131;
input n_54;
input n_132;
input n_188;
input n_102;
input n_186;
input n_204;
input n_0;
input n_87;
input n_195;
input n_189;
input n_32;
input n_66;
input n_85;
input n_99;
input n_78;
input n_84;
input n_130;
input n_213;
input n_164;
input n_100;
input n_129;
input n_13;
input n_121;
input n_197;
input n_11;
input n_137;
input n_17;
input n_23;
input n_203;
input n_142;
input n_20;
input n_143;
input n_207;
input n_2;
input n_180;
input n_19;
input n_47;
input n_62;
input n_29;
input n_155;
input n_75;
input n_109;
input n_150;
input n_122;
input n_45;
input n_205;
input n_34;
input n_140;
input n_70;
input n_120;
input n_37;
input n_15;
input n_67;
input n_33;
input n_82;
input n_27;
input n_38;
input n_110;
input n_151;
input n_61;
input n_112;
input n_172;
input n_81;
input n_59;
input n_181;
input n_76;
input n_36;
input n_182;
input n_26;
input n_124;
input n_55;
input n_126;
input n_202;
input n_94;
input n_97;
input n_108;
input n_58;
input n_116;
input n_211;
input n_64;
input n_117;
input n_118;
input n_175;
input n_48;
input n_65;
input n_25;
input n_40;
input n_93;
input n_80;
input n_141;
input n_135;
input n_196;
input n_200;
input n_165;
input n_139;
input n_41;
input n_134;
input n_177;
input n_176;
input n_114;
input n_86;
input n_198;
input n_104;
input n_95;
input n_179;
input n_9;
input n_107;
input n_10;
input n_71;
input n_74;
input n_6;
input n_190;
input n_14;
input n_123;
input n_136;
input n_72;
input n_187;
input n_89;
input n_173;
input n_201;
input n_103;
input n_111;
input n_60;
input n_159;
input n_157;
input n_162;
input n_170;
input n_185;
input n_35;
input n_183;
input n_115;
input n_12;
input n_69;
input n_128;
input n_30;
input n_79;
input n_43;
input n_194;
input n_171;
input n_31;
input n_192;
input n_57;
input n_169;
input n_53;
input n_51;
input n_44;
input n_56;

output n_2152;

wire n_992;
wire n_1671;
wire n_801;
wire n_1613;
wire n_1234;
wire n_1458;
wire n_1199;
wire n_1674;
wire n_741;
wire n_1027;
wire n_1351;
wire n_625;
wire n_1189;
wire n_223;
wire n_1212;
wire n_226;
wire n_726;
wire n_700;
wire n_1307;
wire n_2003;
wire n_1038;
wire n_578;
wire n_1581;
wire n_1003;
wire n_365;
wire n_1237;
wire n_1061;
wire n_1357;
wire n_1853;
wire n_783;
wire n_1738;
wire n_798;
wire n_1575;
wire n_1854;
wire n_1923;
wire n_509;
wire n_1342;
wire n_245;
wire n_1209;
wire n_1348;
wire n_1387;
wire n_677;
wire n_1708;
wire n_805;
wire n_1151;
wire n_396;
wire n_1739;
wire n_350;
wire n_2051;
wire n_1380;
wire n_442;
wire n_480;
wire n_1402;
wire n_1688;
wire n_1691;
wire n_1975;
wire n_1009;
wire n_1743;
wire n_1930;
wire n_1160;
wire n_883;
wire n_1238;
wire n_1991;
wire n_1724;
wire n_1032;
wire n_1247;
wire n_1547;
wire n_1553;
wire n_893;
wire n_1099;
wire n_1264;
wire n_1192;
wire n_471;
wire n_1844;
wire n_424;
wire n_1700;
wire n_1555;
wire n_1415;
wire n_1370;
wire n_1786;
wire n_369;
wire n_287;
wire n_415;
wire n_830;
wire n_230;
wire n_461;
wire n_873;
wire n_383;
wire n_1285;
wire n_1371;
wire n_1985;
wire n_447;
wire n_1803;
wire n_1172;
wire n_852;
wire n_229;
wire n_1590;
wire n_1532;
wire n_1393;
wire n_1517;
wire n_1867;
wire n_1704;
wire n_1078;
wire n_250;
wire n_544;
wire n_1711;
wire n_1140;
wire n_1444;
wire n_1670;
wire n_1603;
wire n_1579;
wire n_1263;
wire n_2019;
wire n_836;
wire n_375;
wire n_2074;
wire n_522;
wire n_2129;
wire n_1261;
wire n_945;
wire n_1649;
wire n_2018;
wire n_2094;
wire n_1903;
wire n_1511;
wire n_1143;
wire n_1422;
wire n_1232;
wire n_1772;
wire n_1572;
wire n_658;
wire n_616;
wire n_1874;
wire n_1119;
wire n_2013;
wire n_428;
wire n_1433;
wire n_1902;
wire n_1842;
wire n_1620;
wire n_2044;
wire n_1954;
wire n_1735;
wire n_1541;
wire n_1300;
wire n_641;
wire n_822;
wire n_693;
wire n_1313;
wire n_1056;
wire n_758;
wire n_516;
wire n_1455;
wire n_1163;
wire n_1180;
wire n_943;
wire n_1798;
wire n_1550;
wire n_491;
wire n_1591;
wire n_772;
wire n_1344;
wire n_666;
wire n_371;
wire n_940;
wire n_770;
wire n_567;
wire n_1781;
wire n_1971;
wire n_2058;
wire n_2090;
wire n_405;
wire n_538;
wire n_2004;
wire n_1106;
wire n_886;
wire n_1471;
wire n_343;
wire n_953;
wire n_1094;
wire n_1345;
wire n_1820;
wire n_494;
wire n_539;
wire n_493;
wire n_2108;
wire n_454;
wire n_1421;
wire n_1936;
wire n_638;
wire n_1404;
wire n_1211;
wire n_2124;
wire n_381;
wire n_887;
wire n_1660;
wire n_1961;
wire n_1280;
wire n_713;
wire n_1400;
wire n_1467;
wire n_976;
wire n_224;
wire n_1445;
wire n_1526;
wire n_1560;
wire n_734;
wire n_1088;
wire n_1894;
wire n_1231;
wire n_1978;
wire n_2085;
wire n_917;
wire n_574;
wire n_907;
wire n_1446;
wire n_659;
wire n_1815;
wire n_407;
wire n_913;
wire n_1658;
wire n_808;
wire n_867;
wire n_1230;
wire n_473;
wire n_1193;
wire n_1967;
wire n_1054;
wire n_559;
wire n_1333;
wire n_1648;
wire n_1911;
wire n_1956;
wire n_1644;
wire n_2011;
wire n_1558;
wire n_1732;
wire n_281;
wire n_551;
wire n_699;
wire n_1986;
wire n_564;
wire n_451;
wire n_824;
wire n_279;
wire n_686;
wire n_757;
wire n_594;
wire n_1641;
wire n_2113;
wire n_1918;
wire n_577;
wire n_1843;
wire n_619;
wire n_1367;
wire n_1336;
wire n_521;
wire n_572;
wire n_813;
wire n_395;
wire n_2080;
wire n_1909;
wire n_1481;
wire n_323;
wire n_606;
wire n_1441;
wire n_818;
wire n_1123;
wire n_1309;
wire n_2104;
wire n_513;
wire n_645;
wire n_1381;
wire n_331;
wire n_1699;
wire n_916;
wire n_2093;
wire n_483;
wire n_1970;
wire n_608;
wire n_261;
wire n_2101;
wire n_630;
wire n_2059;
wire n_541;
wire n_512;
wire n_2073;
wire n_433;
wire n_792;
wire n_476;
wire n_1328;
wire n_1957;
wire n_219;
wire n_1907;
wire n_264;
wire n_263;
wire n_1162;
wire n_860;
wire n_1530;
wire n_788;
wire n_939;
wire n_1543;
wire n_821;
wire n_938;
wire n_1302;
wire n_1068;
wire n_1599;
wire n_329;
wire n_982;
wire n_549;
wire n_1762;
wire n_1910;
wire n_1075;
wire n_408;
wire n_932;
wire n_237;
wire n_1876;
wire n_1895;
wire n_2123;
wire n_1697;
wire n_2143;
wire n_243;
wire n_979;
wire n_1873;
wire n_905;
wire n_1866;
wire n_1680;
wire n_322;
wire n_993;
wire n_689;
wire n_2031;
wire n_354;
wire n_2130;
wire n_1330;
wire n_1413;
wire n_1605;
wire n_1988;
wire n_1278;
wire n_547;
wire n_558;
wire n_1064;
wire n_1396;
wire n_634;
wire n_966;
wire n_764;
wire n_1663;
wire n_2009;
wire n_692;
wire n_733;
wire n_1793;
wire n_1233;
wire n_1289;
wire n_487;
wire n_241;
wire n_2068;
wire n_1107;
wire n_1014;
wire n_1290;
wire n_1703;
wire n_882;
wire n_2072;
wire n_1354;
wire n_586;
wire n_423;
wire n_1875;
wire n_1865;
wire n_1701;
wire n_318;
wire n_1111;
wire n_1713;
wire n_715;
wire n_1251;
wire n_1265;
wire n_1726;
wire n_1950;
wire n_530;
wire n_1563;
wire n_1912;
wire n_277;
wire n_1982;
wire n_618;
wire n_1297;
wire n_1662;
wire n_1312;
wire n_1167;
wire n_1359;
wire n_674;
wire n_871;
wire n_922;
wire n_268;
wire n_1335;
wire n_1760;
wire n_1927;
wire n_2028;
wire n_1069;
wire n_1664;
wire n_1722;
wire n_612;
wire n_247;
wire n_1165;
wire n_355;
wire n_702;
wire n_347;
wire n_2008;
wire n_1926;
wire n_1175;
wire n_328;
wire n_1386;
wire n_1896;
wire n_429;
wire n_1747;
wire n_1012;
wire n_780;
wire n_675;
wire n_903;
wire n_1540;
wire n_1977;
wire n_1802;
wire n_1504;
wire n_286;
wire n_254;
wire n_1655;
wire n_242;
wire n_835;
wire n_928;
wire n_1214;
wire n_850;
wire n_690;
wire n_1801;
wire n_1886;
wire n_2092;
wire n_1654;
wire n_816;
wire n_1157;
wire n_1750;
wire n_1462;
wire n_1188;
wire n_1752;
wire n_877;
wire n_1813;
wire n_604;
wire n_825;
wire n_728;
wire n_1063;
wire n_1588;
wire n_267;
wire n_1124;
wire n_1624;
wire n_515;
wire n_2096;
wire n_1965;
wire n_598;
wire n_696;
wire n_1515;
wire n_961;
wire n_437;
wire n_1082;
wire n_1317;
wire n_593;
wire n_514;
wire n_697;
wire n_687;
wire n_890;
wire n_637;
wire n_701;
wire n_295;
wire n_950;
wire n_388;
wire n_484;
wire n_2036;
wire n_1709;
wire n_1825;
wire n_1796;
wire n_1757;
wire n_1792;
wire n_891;
wire n_2067;
wire n_2136;
wire n_2082;
wire n_1412;
wire n_949;
wire n_1630;
wire n_678;
wire n_283;
wire n_2075;
wire n_1987;
wire n_507;
wire n_968;
wire n_909;
wire n_1369;
wire n_881;
wire n_1008;
wire n_760;
wire n_1546;
wire n_590;
wire n_362;
wire n_462;
wire n_1033;
wire n_1052;
wire n_1296;
wire n_1990;
wire n_304;
wire n_694;
wire n_2150;
wire n_1294;
wire n_1420;
wire n_1634;
wire n_2078;
wire n_297;
wire n_627;
wire n_595;
wire n_1767;
wire n_1779;
wire n_524;
wire n_1465;
wire n_342;
wire n_1858;
wire n_1044;
wire n_2133;
wire n_1712;
wire n_1391;
wire n_449;
wire n_1523;
wire n_1208;
wire n_1164;
wire n_1295;
wire n_1627;
wire n_1072;
wire n_1527;
wire n_1495;
wire n_1438;
wire n_495;
wire n_815;
wire n_1100;
wire n_585;
wire n_1487;
wire n_840;
wire n_874;
wire n_1756;
wire n_1128;
wire n_673;
wire n_382;
wire n_1969;
wire n_1071;
wire n_1067;
wire n_1565;
wire n_1493;
wire n_2145;
wire n_1968;
wire n_898;
wire n_255;
wire n_284;
wire n_1952;
wire n_865;
wire n_925;
wire n_1932;
wire n_1101;
wire n_1026;
wire n_1880;
wire n_289;
wire n_1364;
wire n_615;
wire n_1249;
wire n_1293;
wire n_1127;
wire n_1512;
wire n_2151;
wire n_1451;
wire n_320;
wire n_639;
wire n_963;
wire n_794;
wire n_727;
wire n_894;
wire n_1839;
wire n_685;
wire n_1765;
wire n_353;
wire n_605;
wire n_1514;
wire n_1863;
wire n_826;
wire n_1646;
wire n_872;
wire n_1139;
wire n_1714;
wire n_718;
wire n_1018;
wire n_1521;
wire n_1366;
wire n_542;
wire n_847;
wire n_644;
wire n_682;
wire n_851;
wire n_305;
wire n_996;
wire n_532;
wire n_1308;
wire n_2089;
wire n_1376;
wire n_1513;
wire n_413;
wire n_791;
wire n_1913;
wire n_510;
wire n_837;
wire n_2097;
wire n_1488;
wire n_1808;
wire n_948;
wire n_704;
wire n_2148;
wire n_977;
wire n_1005;
wire n_1947;
wire n_536;
wire n_1788;
wire n_1999;
wire n_622;
wire n_1469;
wire n_2060;
wire n_1838;
wire n_1835;
wire n_1766;
wire n_1776;
wire n_1959;
wire n_2002;
wire n_581;
wire n_2138;
wire n_765;
wire n_432;
wire n_987;
wire n_1492;
wire n_1340;
wire n_1771;
wire n_631;
wire n_720;
wire n_842;
wire n_1707;
wire n_1432;
wire n_843;
wire n_656;
wire n_989;
wire n_1277;
wire n_797;
wire n_1473;
wire n_1723;
wire n_1246;
wire n_1878;
wire n_899;
wire n_738;
wire n_2012;
wire n_1304;
wire n_1035;
wire n_294;
wire n_499;
wire n_1426;
wire n_705;
wire n_1004;
wire n_1176;
wire n_2134;
wire n_1529;
wire n_1022;
wire n_614;
wire n_529;
wire n_2069;
wire n_425;
wire n_684;
wire n_1431;
wire n_1615;
wire n_1474;
wire n_1571;
wire n_1809;
wire n_1577;
wire n_1181;
wire n_2119;
wire n_1822;
wire n_486;
wire n_947;
wire n_1117;
wire n_1087;
wire n_1448;
wire n_1992;
wire n_648;
wire n_657;
wire n_1049;
wire n_2057;
wire n_2103;
wire n_1666;
wire n_1505;
wire n_803;
wire n_290;
wire n_1717;
wire n_926;
wire n_1817;
wire n_927;
wire n_1849;
wire n_919;
wire n_1698;
wire n_478;
wire n_929;
wire n_1228;
wire n_417;
wire n_446;
wire n_1568;
wire n_1490;
wire n_777;
wire n_1299;
wire n_272;
wire n_526;
wire n_1183;
wire n_1436;
wire n_1384;
wire n_293;
wire n_458;
wire n_1070;
wire n_998;
wire n_717;
wire n_1665;
wire n_1383;
wire n_1178;
wire n_2127;
wire n_1424;
wire n_1073;
wire n_1000;
wire n_796;
wire n_252;
wire n_1195;
wire n_2137;
wire n_1626;
wire n_1507;
wire n_552;
wire n_1358;
wire n_1811;
wire n_1388;
wire n_216;
wire n_912;
wire n_1857;
wire n_1519;
wire n_2144;
wire n_745;
wire n_1284;
wire n_1604;
wire n_1142;
wire n_716;
wire n_1475;
wire n_623;
wire n_1048;
wire n_1201;
wire n_1398;
wire n_884;
wire n_1774;
wire n_1395;
wire n_2110;
wire n_731;
wire n_1502;
wire n_1659;
wire n_1955;
wire n_755;
wire n_931;
wire n_1021;
wire n_811;
wire n_527;
wire n_683;
wire n_1207;
wire n_474;
wire n_312;
wire n_1791;
wire n_1368;
wire n_1418;
wire n_958;
wire n_292;
wire n_1250;
wire n_1137;
wire n_1897;
wire n_2064;
wire n_880;
wire n_2053;
wire n_2121;
wire n_889;
wire n_1478;
wire n_589;
wire n_1310;
wire n_819;
wire n_1363;
wire n_1334;
wire n_1942;
wire n_1966;
wire n_767;
wire n_1314;
wire n_600;
wire n_964;
wire n_831;
wire n_1837;
wire n_477;
wire n_954;
wire n_864;
wire n_1110;
wire n_1410;
wire n_399;
wire n_1440;
wire n_2132;
wire n_2063;
wire n_1382;
wire n_1534;
wire n_1564;
wire n_1736;
wire n_1483;
wire n_1834;
wire n_1372;
wire n_231;
wire n_1457;
wire n_505;
wire n_1719;
wire n_319;
wire n_1339;
wire n_1787;
wire n_537;
wire n_1993;
wire n_1427;
wire n_311;
wire n_1466;
wire n_403;
wire n_1919;
wire n_1080;
wire n_723;
wire n_1877;
wire n_596;
wire n_546;
wire n_562;
wire n_1141;
wire n_1268;
wire n_386;
wire n_1939;
wire n_2030;
wire n_1769;
wire n_1220;
wire n_1893;
wire n_556;
wire n_1755;
wire n_1602;
wire n_1136;
wire n_2025;
wire n_1125;
wire n_970;
wire n_1980;
wire n_642;
wire n_995;
wire n_276;
wire n_1159;
wire n_1092;
wire n_441;
wire n_221;
wire n_1060;
wire n_1951;
wire n_444;
wire n_1252;
wire n_1784;
wire n_1223;
wire n_303;
wire n_511;
wire n_1286;
wire n_1773;
wire n_1775;
wire n_2115;
wire n_1053;
wire n_416;
wire n_1681;
wire n_520;
wire n_1093;
wire n_418;
wire n_1783;
wire n_1533;
wire n_1597;
wire n_266;
wire n_296;
wire n_775;
wire n_651;
wire n_1153;
wire n_439;
wire n_1618;
wire n_217;
wire n_518;
wire n_1531;
wire n_1185;
wire n_453;
wire n_215;
wire n_1745;
wire n_914;
wire n_759;
wire n_1831;
wire n_426;
wire n_317;
wire n_1653;
wire n_1679;
wire n_1625;
wire n_1453;
wire n_2146;
wire n_2131;
wire n_488;
wire n_497;
wire n_773;
wire n_1901;
wire n_920;
wire n_1374;
wire n_1315;
wire n_1647;
wire n_1224;
wire n_1614;
wire n_1459;
wire n_1892;
wire n_1933;
wire n_1135;
wire n_1169;
wire n_1179;
wire n_401;
wire n_324;
wire n_1617;
wire n_335;
wire n_1470;
wire n_463;
wire n_1243;
wire n_848;
wire n_301;
wire n_274;
wire n_1096;
wire n_1091;
wire n_1917;
wire n_2000;
wire n_1580;
wire n_1425;
wire n_1881;
wire n_1267;
wire n_1281;
wire n_1806;
wire n_983;
wire n_2023;
wire n_427;
wire n_1520;
wire n_496;
wire n_906;
wire n_1390;
wire n_688;
wire n_1077;
wire n_1733;
wire n_1419;
wire n_351;
wire n_259;
wire n_1731;
wire n_2087;
wire n_1855;
wire n_1636;
wire n_1437;
wire n_2135;
wire n_1645;
wire n_1832;
wire n_385;
wire n_1687;
wire n_1439;
wire n_1323;
wire n_858;
wire n_2049;
wire n_1331;
wire n_736;
wire n_613;
wire n_501;
wire n_956;
wire n_960;
wire n_663;
wire n_856;
wire n_2100;
wire n_379;
wire n_778;
wire n_1668;
wire n_1134;
wire n_410;
wire n_1129;
wire n_554;
wire n_602;
wire n_1696;
wire n_1995;
wire n_1594;
wire n_664;
wire n_1869;
wire n_1764;
wire n_1429;
wire n_1610;
wire n_1889;
wire n_435;
wire n_1905;
wire n_2016;
wire n_793;
wire n_326;
wire n_587;
wire n_1593;
wire n_580;
wire n_762;
wire n_1202;
wire n_1030;
wire n_1937;
wire n_465;
wire n_1790;
wire n_1778;
wire n_1635;
wire n_1079;
wire n_341;
wire n_1744;
wire n_828;
wire n_2139;
wire n_2142;
wire n_607;
wire n_316;
wire n_419;
wire n_1551;
wire n_1103;
wire n_1203;
wire n_820;
wire n_951;
wire n_725;
wire n_952;
wire n_999;
wire n_358;
wire n_1254;
wire n_575;
wire n_368;
wire n_994;
wire n_1508;
wire n_732;
wire n_974;
wire n_392;
wire n_724;
wire n_1934;
wire n_1020;
wire n_1042;
wire n_628;
wire n_1273;
wire n_1434;
wire n_1573;
wire n_1728;
wire n_557;
wire n_1871;
wire n_349;
wire n_617;
wire n_845;
wire n_807;
wire n_1036;
wire n_1138;
wire n_1661;
wire n_1275;
wire n_485;
wire n_1549;
wire n_443;
wire n_1510;
wire n_892;
wire n_768;
wire n_421;
wire n_1468;
wire n_1859;
wire n_2102;
wire n_238;
wire n_1095;
wire n_2024;
wire n_1595;
wire n_1718;
wire n_1749;
wire n_1683;
wire n_1916;
wire n_597;
wire n_280;
wire n_1270;
wire n_1187;
wire n_610;
wire n_1403;
wire n_1669;
wire n_1852;
wire n_1024;
wire n_1768;
wire n_1847;
wire n_2052;
wire n_248;
wire n_517;
wire n_1667;
wire n_667;
wire n_1206;
wire n_621;
wire n_1037;
wire n_1397;
wire n_1279;
wire n_1115;
wire n_750;
wire n_901;
wire n_1499;
wire n_468;
wire n_923;
wire n_504;
wire n_1409;
wire n_1841;
wire n_1639;
wire n_1623;
wire n_1015;
wire n_1503;
wire n_466;
wire n_1057;
wire n_603;
wire n_991;
wire n_1657;
wire n_235;
wire n_1126;
wire n_1997;
wire n_340;
wire n_710;
wire n_1108;
wire n_1818;
wire n_1182;
wire n_1298;
wire n_2088;
wire n_1611;
wire n_785;
wire n_746;
wire n_609;
wire n_1601;
wire n_1960;
wire n_2061;
wire n_1686;
wire n_1356;
wire n_1589;
wire n_1740;
wire n_1497;
wire n_1168;
wire n_1216;
wire n_1943;
wire n_1320;
wire n_1430;
wire n_1316;
wire n_1287;
wire n_1452;
wire n_1622;
wire n_1586;
wire n_302;
wire n_1694;
wire n_380;
wire n_1535;
wire n_1596;
wire n_1190;
wire n_1734;
wire n_397;
wire n_1983;
wire n_1938;
wire n_1262;
wire n_218;
wire n_1891;
wire n_1213;
wire n_1350;
wire n_1673;
wire n_1715;
wire n_1443;
wire n_1272;
wire n_239;
wire n_2037;
wire n_782;
wire n_1539;
wire n_490;
wire n_220;
wire n_809;
wire n_1043;
wire n_1797;
wire n_1608;
wire n_986;
wire n_2120;
wire n_1472;
wire n_2050;
wire n_1081;
wire n_402;
wire n_1870;
wire n_352;
wire n_1692;
wire n_800;
wire n_1084;
wire n_1171;
wire n_460;
wire n_1827;
wire n_1361;
wire n_1864;
wire n_2006;
wire n_1491;
wire n_662;
wire n_374;
wire n_1152;
wire n_1840;
wire n_1705;
wire n_450;
wire n_1684;
wire n_921;
wire n_1346;
wire n_711;
wire n_1642;
wire n_579;
wire n_1352;
wire n_937;
wire n_1682;
wire n_2017;
wire n_370;
wire n_1695;
wire n_1828;
wire n_2046;
wire n_650;
wire n_1046;
wire n_1940;
wire n_1979;
wire n_1145;
wire n_330;
wire n_1121;
wire n_1102;
wire n_1963;
wire n_972;
wire n_1405;
wire n_258;
wire n_1406;
wire n_456;
wire n_1332;
wire n_260;
wire n_313;
wire n_624;
wire n_962;
wire n_1041;
wire n_565;
wire n_356;
wire n_1569;
wire n_936;
wire n_1883;
wire n_1288;
wire n_1186;
wire n_1062;
wire n_885;
wire n_896;
wire n_2084;
wire n_654;
wire n_411;
wire n_1222;
wire n_599;
wire n_776;
wire n_321;
wire n_1823;
wire n_227;
wire n_1974;
wire n_1720;
wire n_482;
wire n_934;
wire n_1637;
wire n_1407;
wire n_1795;
wire n_420;
wire n_1341;
wire n_394;
wire n_1456;
wire n_1845;
wire n_1489;
wire n_942;
wire n_1524;
wire n_543;
wire n_1964;
wire n_1920;
wire n_2099;
wire n_1496;
wire n_1271;
wire n_1545;
wire n_2007;
wire n_2039;
wire n_1946;
wire n_1355;
wire n_1225;
wire n_1544;
wire n_1485;
wire n_325;
wire n_1640;
wire n_804;
wire n_464;
wire n_1846;
wire n_533;
wire n_806;
wire n_879;
wire n_959;
wire n_584;
wire n_2141;
wire n_244;
wire n_1343;
wire n_1522;
wire n_548;
wire n_1782;
wire n_282;
wire n_1676;
wire n_833;
wire n_1830;
wire n_1567;
wire n_523;
wire n_1319;
wire n_707;
wire n_345;
wire n_1900;
wire n_799;
wire n_1548;
wire n_1155;
wire n_273;
wire n_1633;
wire n_787;
wire n_1416;
wire n_1528;
wire n_1146;
wire n_2021;
wire n_2114;
wire n_1086;
wire n_1066;
wire n_1948;
wire n_2125;
wire n_2026;
wire n_1282;
wire n_550;
wire n_275;
wire n_652;
wire n_560;
wire n_1906;
wire n_1484;
wire n_1241;
wire n_1321;
wire n_1672;
wire n_569;
wire n_1758;
wire n_1925;
wire n_737;
wire n_1318;
wire n_1914;
wire n_1235;
wire n_1229;
wire n_306;
wire n_1292;
wire n_1373;
wire n_346;
wire n_1029;
wire n_1447;
wire n_2056;
wire n_790;
wire n_1706;
wire n_1498;
wire n_1210;
wire n_299;
wire n_1248;
wire n_1556;
wire n_902;
wire n_333;
wire n_1047;
wire n_1984;
wire n_1385;
wire n_431;
wire n_459;
wire n_1269;
wire n_1931;
wire n_2083;
wire n_502;
wire n_672;
wire n_1257;
wire n_1751;
wire n_285;
wire n_1375;
wire n_1941;
wire n_2128;
wire n_655;
wire n_706;
wire n_1045;
wire n_1650;
wire n_786;
wire n_1962;
wire n_1236;
wire n_1794;
wire n_1559;
wire n_1725;
wire n_1928;
wire n_1872;
wire n_834;
wire n_743;
wire n_766;
wire n_430;
wire n_1746;
wire n_1325;
wire n_1002;
wire n_1741;
wire n_1949;
wire n_545;
wire n_489;
wire n_1804;
wire n_1727;
wire n_251;
wire n_1019;
wire n_636;
wire n_2054;
wire n_729;
wire n_876;
wire n_774;
wire n_1337;
wire n_660;
wire n_2062;
wire n_2041;
wire n_438;
wire n_1477;
wire n_1360;
wire n_1860;
wire n_1904;
wire n_1200;
wire n_2070;
wire n_479;
wire n_1607;
wire n_1353;
wire n_1777;
wire n_1908;
wire n_1454;
wire n_2126;
wire n_869;
wire n_1154;
wire n_1113;
wire n_1600;
wire n_646;
wire n_528;
wire n_391;
wire n_1098;
wire n_1329;
wire n_2045;
wire n_817;
wire n_262;
wire n_897;
wire n_846;
wire n_2066;
wire n_841;
wire n_1476;
wire n_1001;
wire n_508;
wire n_1800;
wire n_1050;
wire n_1411;
wire n_1463;
wire n_1177;
wire n_332;
wire n_1150;
wire n_1742;
wire n_1562;
wire n_1690;
wire n_398;
wire n_1191;
wire n_1826;
wire n_566;
wire n_1023;
wire n_1882;
wire n_1076;
wire n_1118;
wire n_1007;
wire n_1807;
wire n_1929;
wire n_1378;
wire n_855;
wire n_1592;
wire n_1759;
wire n_1814;
wire n_1631;
wire n_591;
wire n_1377;
wire n_1879;
wire n_256;
wire n_853;
wire n_440;
wire n_695;
wire n_1542;
wire n_875;
wire n_680;
wire n_367;
wire n_1678;
wire n_661;
wire n_1716;
wire n_278;
wire n_1256;
wire n_671;
wire n_1953;
wire n_933;
wire n_740;
wire n_703;
wire n_978;
wire n_384;
wire n_1976;
wire n_1291;
wire n_1217;
wire n_751;
wire n_749;
wire n_1824;
wire n_310;
wire n_1628;
wire n_1324;
wire n_1399;
wire n_2122;
wire n_2109;
wire n_1435;
wire n_969;
wire n_988;
wire n_2140;
wire n_1065;
wire n_1401;
wire n_1255;
wire n_568;
wire n_1516;
wire n_1536;
wire n_2029;
wire n_1204;
wire n_823;
wire n_1132;
wire n_643;
wire n_233;
wire n_698;
wire n_1074;
wire n_1394;
wire n_1327;
wire n_1326;
wire n_739;
wire n_400;
wire n_955;
wire n_337;
wire n_1379;
wire n_214;
wire n_246;
wire n_1338;
wire n_1097;
wire n_935;
wire n_781;
wire n_789;
wire n_1554;
wire n_1130;
wire n_1810;
wire n_573;
wire n_769;
wire n_676;
wire n_327;
wire n_1120;
wire n_832;
wire n_1583;
wire n_1730;
wire n_555;
wire n_389;
wire n_814;
wire n_1643;
wire n_2020;
wire n_1729;
wire n_669;
wire n_2048;
wire n_300;
wire n_222;
wire n_2005;
wire n_747;
wire n_1389;
wire n_1105;
wire n_721;
wire n_1461;
wire n_742;
wire n_535;
wire n_691;
wire n_372;
wire n_2076;
wire n_314;
wire n_1408;
wire n_378;
wire n_1196;
wire n_377;
wire n_1598;
wire n_863;
wire n_601;
wire n_338;
wire n_1283;
wire n_918;
wire n_748;
wire n_506;
wire n_1114;
wire n_1785;
wire n_763;
wire n_1147;
wire n_1848;
wire n_360;
wire n_1754;
wire n_2149;
wire n_1506;
wire n_1652;
wire n_1812;
wire n_957;
wire n_1994;
wire n_895;
wire n_866;
wire n_1227;
wire n_387;
wire n_452;
wire n_744;
wire n_971;
wire n_946;
wire n_344;
wire n_761;
wire n_1303;
wire n_1205;
wire n_1258;
wire n_1392;
wire n_1173;
wire n_1924;
wire n_525;
wire n_1677;
wire n_1116;
wire n_611;
wire n_1570;
wire n_1702;
wire n_1219;
wire n_1780;
wire n_1689;
wire n_1174;
wire n_1944;
wire n_1016;
wire n_1347;
wire n_795;
wire n_1501;
wire n_1221;
wire n_1245;
wire n_838;
wire n_647;
wire n_844;
wire n_448;
wire n_1017;
wire n_2117;
wire n_1083;
wire n_445;
wire n_1561;
wire n_930;
wire n_888;
wire n_1112;
wire n_2081;
wire n_234;
wire n_2022;
wire n_1945;
wire n_910;
wire n_1656;
wire n_1721;
wire n_1460;
wire n_911;
wire n_2112;
wire n_1464;
wire n_236;
wire n_653;
wire n_1737;
wire n_1414;
wire n_752;
wire n_908;
wire n_944;
wire n_2034;
wire n_576;
wire n_1028;
wire n_2106;
wire n_472;
wire n_270;
wire n_414;
wire n_1922;
wire n_563;
wire n_2032;
wire n_1011;
wire n_1566;
wire n_1215;
wire n_839;
wire n_708;
wire n_1973;
wire n_668;
wire n_626;
wire n_990;
wire n_1500;
wire n_779;
wire n_1537;
wire n_1821;
wire n_1104;
wire n_854;
wire n_1058;
wire n_498;
wire n_1122;
wire n_870;
wire n_904;
wire n_1253;
wire n_709;
wire n_1266;
wire n_366;
wire n_1509;
wire n_1693;
wire n_1109;
wire n_712;
wire n_348;
wire n_1276;
wire n_376;
wire n_2015;
wire n_2118;
wire n_2111;
wire n_390;
wire n_1148;
wire n_334;
wire n_1989;
wire n_1161;
wire n_1085;
wire n_232;
wire n_2014;
wire n_2042;
wire n_1239;
wire n_771;
wire n_1584;
wire n_470;
wire n_475;
wire n_924;
wire n_298;
wire n_1582;
wire n_492;
wire n_1149;
wire n_265;
wire n_1184;
wire n_228;
wire n_719;
wire n_1972;
wire n_1525;
wire n_455;
wire n_1585;
wire n_1851;
wire n_363;
wire n_1799;
wire n_1090;
wire n_2147;
wire n_592;
wire n_1816;
wire n_1518;
wire n_829;
wire n_1156;
wire n_1362;
wire n_393;
wire n_984;
wire n_1829;
wire n_503;
wire n_2035;
wire n_1450;
wire n_1638;
wire n_868;
wire n_570;
wire n_859;
wire n_2033;
wire n_406;
wire n_735;
wire n_1789;
wire n_1770;
wire n_878;
wire n_620;
wire n_519;
wire n_307;
wire n_469;
wire n_1218;
wire n_500;
wire n_1482;
wire n_981;
wire n_714;
wire n_1349;
wire n_291;
wire n_1144;
wire n_2071;
wire n_357;
wire n_985;
wire n_481;
wire n_997;
wire n_1710;
wire n_1301;
wire n_802;
wire n_561;
wire n_980;
wire n_1306;
wire n_2010;
wire n_1651;
wire n_1198;
wire n_2047;
wire n_2095;
wire n_1609;
wire n_436;
wire n_409;
wire n_1244;
wire n_1685;
wire n_1763;
wire n_1998;
wire n_1574;
wire n_240;
wire n_756;
wire n_1619;
wire n_1981;
wire n_1606;
wire n_810;
wire n_1133;
wire n_635;
wire n_1194;
wire n_1051;
wire n_253;
wire n_1552;
wire n_583;
wire n_1996;
wire n_249;
wire n_1039;
wire n_1442;
wire n_1034;
wire n_2043;
wire n_1480;
wire n_1158;
wire n_754;
wire n_941;
wire n_975;
wire n_1031;
wire n_1305;
wire n_553;
wire n_849;
wire n_753;
wire n_1753;
wire n_467;
wire n_269;
wire n_359;
wire n_973;
wire n_1921;
wire n_1479;
wire n_1055;
wire n_1675;
wire n_582;
wire n_2065;
wire n_861;
wire n_857;
wire n_967;
wire n_571;
wire n_271;
wire n_404;
wire n_2001;
wire n_2107;
wire n_1884;
wire n_2040;
wire n_679;
wire n_633;
wire n_1170;
wire n_665;
wire n_1629;
wire n_588;
wire n_225;
wire n_1260;
wire n_308;
wire n_309;
wire n_2055;
wire n_1819;
wire n_1010;
wire n_1040;
wire n_915;
wire n_632;
wire n_1166;
wire n_2038;
wire n_812;
wire n_1131;
wire n_1761;
wire n_534;
wire n_1578;
wire n_1006;
wire n_1861;
wire n_373;
wire n_1632;
wire n_1890;
wire n_1805;
wire n_257;
wire n_1557;
wire n_1888;
wire n_1833;
wire n_730;
wire n_1311;
wire n_1494;
wire n_670;
wire n_1850;
wire n_1898;
wire n_1868;
wire n_2079;
wire n_1089;
wire n_1887;
wire n_1587;
wire n_1365;
wire n_1417;
wire n_1242;
wire n_2086;
wire n_1836;
wire n_681;
wire n_1226;
wire n_1274;
wire n_1486;
wire n_412;
wire n_640;
wire n_1322;
wire n_965;
wire n_1899;
wire n_1428;
wire n_1616;
wire n_1576;
wire n_1856;
wire n_1862;
wire n_1958;
wire n_2077;
wire n_339;
wire n_784;
wire n_315;
wire n_434;
wire n_288;
wire n_1059;
wire n_1197;
wire n_422;
wire n_722;
wire n_862;
wire n_2105;
wire n_2098;
wire n_540;
wire n_1423;
wire n_1935;
wire n_2027;
wire n_457;
wire n_2091;
wire n_364;
wire n_1915;
wire n_629;
wire n_1621;
wire n_1748;
wire n_900;
wire n_1449;
wire n_531;
wire n_827;
wire n_361;
wire n_1025;
wire n_2116;
wire n_336;
wire n_1885;
wire n_1013;
wire n_1259;
wire n_1538;
wire n_649;
wire n_1612;
wire n_1240;

INVx1_ASAP7_75t_L g214 ( 
.A(n_37),
.Y(n_214)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_131),
.Y(n_215)
);

CKINVDCx5p33_ASAP7_75t_R g216 ( 
.A(n_197),
.Y(n_216)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_133),
.Y(n_217)
);

CKINVDCx5p33_ASAP7_75t_R g218 ( 
.A(n_180),
.Y(n_218)
);

INVxp33_ASAP7_75t_R g219 ( 
.A(n_193),
.Y(n_219)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_81),
.Y(n_220)
);

CKINVDCx20_ASAP7_75t_R g221 ( 
.A(n_54),
.Y(n_221)
);

CKINVDCx5p33_ASAP7_75t_R g222 ( 
.A(n_202),
.Y(n_222)
);

CKINVDCx5p33_ASAP7_75t_R g223 ( 
.A(n_200),
.Y(n_223)
);

CKINVDCx5p33_ASAP7_75t_R g224 ( 
.A(n_112),
.Y(n_224)
);

CKINVDCx5p33_ASAP7_75t_R g225 ( 
.A(n_140),
.Y(n_225)
);

CKINVDCx5p33_ASAP7_75t_R g226 ( 
.A(n_156),
.Y(n_226)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_3),
.Y(n_227)
);

BUFx10_ASAP7_75t_L g228 ( 
.A(n_172),
.Y(n_228)
);

INVxp67_ASAP7_75t_L g229 ( 
.A(n_1),
.Y(n_229)
);

BUFx3_ASAP7_75t_L g230 ( 
.A(n_12),
.Y(n_230)
);

CKINVDCx5p33_ASAP7_75t_R g231 ( 
.A(n_33),
.Y(n_231)
);

CKINVDCx5p33_ASAP7_75t_R g232 ( 
.A(n_62),
.Y(n_232)
);

INVx2_ASAP7_75t_L g233 ( 
.A(n_129),
.Y(n_233)
);

INVx2_ASAP7_75t_L g234 ( 
.A(n_132),
.Y(n_234)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_146),
.Y(n_235)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_136),
.Y(n_236)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_69),
.Y(n_237)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_89),
.Y(n_238)
);

CKINVDCx5p33_ASAP7_75t_R g239 ( 
.A(n_155),
.Y(n_239)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_141),
.Y(n_240)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_51),
.Y(n_241)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_107),
.Y(n_242)
);

CKINVDCx20_ASAP7_75t_R g243 ( 
.A(n_38),
.Y(n_243)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_17),
.Y(n_244)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_61),
.Y(n_245)
);

INVx2_ASAP7_75t_L g246 ( 
.A(n_8),
.Y(n_246)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_12),
.Y(n_247)
);

CKINVDCx5p33_ASAP7_75t_R g248 ( 
.A(n_99),
.Y(n_248)
);

INVx2_ASAP7_75t_SL g249 ( 
.A(n_210),
.Y(n_249)
);

CKINVDCx5p33_ASAP7_75t_R g250 ( 
.A(n_186),
.Y(n_250)
);

CKINVDCx5p33_ASAP7_75t_R g251 ( 
.A(n_40),
.Y(n_251)
);

INVx2_ASAP7_75t_L g252 ( 
.A(n_106),
.Y(n_252)
);

CKINVDCx5p33_ASAP7_75t_R g253 ( 
.A(n_113),
.Y(n_253)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_167),
.Y(n_254)
);

INVx2_ASAP7_75t_L g255 ( 
.A(n_46),
.Y(n_255)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_189),
.Y(n_256)
);

CKINVDCx14_ASAP7_75t_R g257 ( 
.A(n_58),
.Y(n_257)
);

BUFx2_ASAP7_75t_L g258 ( 
.A(n_123),
.Y(n_258)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_194),
.Y(n_259)
);

CKINVDCx20_ASAP7_75t_R g260 ( 
.A(n_80),
.Y(n_260)
);

BUFx3_ASAP7_75t_L g261 ( 
.A(n_86),
.Y(n_261)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_23),
.Y(n_262)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_183),
.Y(n_263)
);

INVx2_ASAP7_75t_SL g264 ( 
.A(n_42),
.Y(n_264)
);

CKINVDCx5p33_ASAP7_75t_R g265 ( 
.A(n_101),
.Y(n_265)
);

CKINVDCx5p33_ASAP7_75t_R g266 ( 
.A(n_173),
.Y(n_266)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_147),
.Y(n_267)
);

INVx1_ASAP7_75t_SL g268 ( 
.A(n_57),
.Y(n_268)
);

CKINVDCx5p33_ASAP7_75t_R g269 ( 
.A(n_62),
.Y(n_269)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_50),
.Y(n_270)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_162),
.Y(n_271)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_23),
.Y(n_272)
);

CKINVDCx5p33_ASAP7_75t_R g273 ( 
.A(n_100),
.Y(n_273)
);

CKINVDCx5p33_ASAP7_75t_R g274 ( 
.A(n_198),
.Y(n_274)
);

CKINVDCx5p33_ASAP7_75t_R g275 ( 
.A(n_204),
.Y(n_275)
);

CKINVDCx5p33_ASAP7_75t_R g276 ( 
.A(n_72),
.Y(n_276)
);

CKINVDCx5p33_ASAP7_75t_R g277 ( 
.A(n_60),
.Y(n_277)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_67),
.Y(n_278)
);

CKINVDCx5p33_ASAP7_75t_R g279 ( 
.A(n_150),
.Y(n_279)
);

CKINVDCx5p33_ASAP7_75t_R g280 ( 
.A(n_175),
.Y(n_280)
);

CKINVDCx5p33_ASAP7_75t_R g281 ( 
.A(n_68),
.Y(n_281)
);

CKINVDCx5p33_ASAP7_75t_R g282 ( 
.A(n_134),
.Y(n_282)
);

CKINVDCx5p33_ASAP7_75t_R g283 ( 
.A(n_30),
.Y(n_283)
);

CKINVDCx5p33_ASAP7_75t_R g284 ( 
.A(n_108),
.Y(n_284)
);

CKINVDCx20_ASAP7_75t_R g285 ( 
.A(n_58),
.Y(n_285)
);

CKINVDCx5p33_ASAP7_75t_R g286 ( 
.A(n_35),
.Y(n_286)
);

CKINVDCx5p33_ASAP7_75t_R g287 ( 
.A(n_28),
.Y(n_287)
);

CKINVDCx5p33_ASAP7_75t_R g288 ( 
.A(n_195),
.Y(n_288)
);

CKINVDCx5p33_ASAP7_75t_R g289 ( 
.A(n_91),
.Y(n_289)
);

INVx2_ASAP7_75t_L g290 ( 
.A(n_213),
.Y(n_290)
);

CKINVDCx5p33_ASAP7_75t_R g291 ( 
.A(n_109),
.Y(n_291)
);

CKINVDCx16_ASAP7_75t_R g292 ( 
.A(n_40),
.Y(n_292)
);

INVx2_ASAP7_75t_L g293 ( 
.A(n_35),
.Y(n_293)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_168),
.Y(n_294)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_121),
.Y(n_295)
);

INVx1_ASAP7_75t_SL g296 ( 
.A(n_161),
.Y(n_296)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_78),
.Y(n_297)
);

CKINVDCx5p33_ASAP7_75t_R g298 ( 
.A(n_98),
.Y(n_298)
);

INVx2_ASAP7_75t_L g299 ( 
.A(n_24),
.Y(n_299)
);

CKINVDCx5p33_ASAP7_75t_R g300 ( 
.A(n_10),
.Y(n_300)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_64),
.Y(n_301)
);

BUFx6f_ASAP7_75t_L g302 ( 
.A(n_116),
.Y(n_302)
);

CKINVDCx5p33_ASAP7_75t_R g303 ( 
.A(n_19),
.Y(n_303)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_144),
.Y(n_304)
);

CKINVDCx5p33_ASAP7_75t_R g305 ( 
.A(n_56),
.Y(n_305)
);

CKINVDCx5p33_ASAP7_75t_R g306 ( 
.A(n_69),
.Y(n_306)
);

CKINVDCx5p33_ASAP7_75t_R g307 ( 
.A(n_88),
.Y(n_307)
);

CKINVDCx5p33_ASAP7_75t_R g308 ( 
.A(n_38),
.Y(n_308)
);

CKINVDCx5p33_ASAP7_75t_R g309 ( 
.A(n_96),
.Y(n_309)
);

CKINVDCx5p33_ASAP7_75t_R g310 ( 
.A(n_203),
.Y(n_310)
);

CKINVDCx5p33_ASAP7_75t_R g311 ( 
.A(n_205),
.Y(n_311)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_115),
.Y(n_312)
);

CKINVDCx5p33_ASAP7_75t_R g313 ( 
.A(n_178),
.Y(n_313)
);

CKINVDCx5p33_ASAP7_75t_R g314 ( 
.A(n_78),
.Y(n_314)
);

CKINVDCx20_ASAP7_75t_R g315 ( 
.A(n_4),
.Y(n_315)
);

CKINVDCx5p33_ASAP7_75t_R g316 ( 
.A(n_138),
.Y(n_316)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_66),
.Y(n_317)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_93),
.Y(n_318)
);

BUFx10_ASAP7_75t_L g319 ( 
.A(n_212),
.Y(n_319)
);

CKINVDCx5p33_ASAP7_75t_R g320 ( 
.A(n_184),
.Y(n_320)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_137),
.Y(n_321)
);

CKINVDCx5p33_ASAP7_75t_R g322 ( 
.A(n_7),
.Y(n_322)
);

BUFx3_ASAP7_75t_L g323 ( 
.A(n_148),
.Y(n_323)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_79),
.Y(n_324)
);

INVxp67_ASAP7_75t_L g325 ( 
.A(n_102),
.Y(n_325)
);

CKINVDCx5p33_ASAP7_75t_R g326 ( 
.A(n_3),
.Y(n_326)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_43),
.Y(n_327)
);

CKINVDCx5p33_ASAP7_75t_R g328 ( 
.A(n_84),
.Y(n_328)
);

CKINVDCx5p33_ASAP7_75t_R g329 ( 
.A(n_207),
.Y(n_329)
);

CKINVDCx5p33_ASAP7_75t_R g330 ( 
.A(n_166),
.Y(n_330)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_55),
.Y(n_331)
);

CKINVDCx5p33_ASAP7_75t_R g332 ( 
.A(n_61),
.Y(n_332)
);

CKINVDCx5p33_ASAP7_75t_R g333 ( 
.A(n_92),
.Y(n_333)
);

CKINVDCx5p33_ASAP7_75t_R g334 ( 
.A(n_5),
.Y(n_334)
);

CKINVDCx5p33_ASAP7_75t_R g335 ( 
.A(n_145),
.Y(n_335)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_190),
.Y(n_336)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_110),
.Y(n_337)
);

INVx1_ASAP7_75t_L g338 ( 
.A(n_152),
.Y(n_338)
);

CKINVDCx5p33_ASAP7_75t_R g339 ( 
.A(n_171),
.Y(n_339)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_55),
.Y(n_340)
);

CKINVDCx5p33_ASAP7_75t_R g341 ( 
.A(n_185),
.Y(n_341)
);

INVx1_ASAP7_75t_L g342 ( 
.A(n_47),
.Y(n_342)
);

INVx1_ASAP7_75t_L g343 ( 
.A(n_52),
.Y(n_343)
);

CKINVDCx5p33_ASAP7_75t_R g344 ( 
.A(n_105),
.Y(n_344)
);

CKINVDCx5p33_ASAP7_75t_R g345 ( 
.A(n_66),
.Y(n_345)
);

CKINVDCx14_ASAP7_75t_R g346 ( 
.A(n_71),
.Y(n_346)
);

CKINVDCx5p33_ASAP7_75t_R g347 ( 
.A(n_122),
.Y(n_347)
);

INVx1_ASAP7_75t_L g348 ( 
.A(n_6),
.Y(n_348)
);

INVx1_ASAP7_75t_L g349 ( 
.A(n_83),
.Y(n_349)
);

CKINVDCx5p33_ASAP7_75t_R g350 ( 
.A(n_157),
.Y(n_350)
);

CKINVDCx5p33_ASAP7_75t_R g351 ( 
.A(n_25),
.Y(n_351)
);

INVx1_ASAP7_75t_L g352 ( 
.A(n_36),
.Y(n_352)
);

CKINVDCx5p33_ASAP7_75t_R g353 ( 
.A(n_165),
.Y(n_353)
);

CKINVDCx5p33_ASAP7_75t_R g354 ( 
.A(n_30),
.Y(n_354)
);

CKINVDCx5p33_ASAP7_75t_R g355 ( 
.A(n_176),
.Y(n_355)
);

INVx1_ASAP7_75t_L g356 ( 
.A(n_159),
.Y(n_356)
);

BUFx6f_ASAP7_75t_L g357 ( 
.A(n_127),
.Y(n_357)
);

INVx1_ASAP7_75t_L g358 ( 
.A(n_63),
.Y(n_358)
);

INVxp67_ASAP7_75t_L g359 ( 
.A(n_142),
.Y(n_359)
);

CKINVDCx5p33_ASAP7_75t_R g360 ( 
.A(n_103),
.Y(n_360)
);

CKINVDCx5p33_ASAP7_75t_R g361 ( 
.A(n_47),
.Y(n_361)
);

INVx1_ASAP7_75t_L g362 ( 
.A(n_14),
.Y(n_362)
);

CKINVDCx20_ASAP7_75t_R g363 ( 
.A(n_206),
.Y(n_363)
);

INVx2_ASAP7_75t_SL g364 ( 
.A(n_4),
.Y(n_364)
);

CKINVDCx5p33_ASAP7_75t_R g365 ( 
.A(n_196),
.Y(n_365)
);

CKINVDCx5p33_ASAP7_75t_R g366 ( 
.A(n_187),
.Y(n_366)
);

CKINVDCx5p33_ASAP7_75t_R g367 ( 
.A(n_53),
.Y(n_367)
);

INVx1_ASAP7_75t_L g368 ( 
.A(n_117),
.Y(n_368)
);

CKINVDCx5p33_ASAP7_75t_R g369 ( 
.A(n_87),
.Y(n_369)
);

CKINVDCx20_ASAP7_75t_R g370 ( 
.A(n_54),
.Y(n_370)
);

CKINVDCx5p33_ASAP7_75t_R g371 ( 
.A(n_22),
.Y(n_371)
);

INVx1_ASAP7_75t_L g372 ( 
.A(n_8),
.Y(n_372)
);

CKINVDCx5p33_ASAP7_75t_R g373 ( 
.A(n_11),
.Y(n_373)
);

INVx2_ASAP7_75t_L g374 ( 
.A(n_73),
.Y(n_374)
);

INVx1_ASAP7_75t_L g375 ( 
.A(n_130),
.Y(n_375)
);

CKINVDCx5p33_ASAP7_75t_R g376 ( 
.A(n_83),
.Y(n_376)
);

CKINVDCx5p33_ASAP7_75t_R g377 ( 
.A(n_85),
.Y(n_377)
);

BUFx2_ASAP7_75t_SL g378 ( 
.A(n_151),
.Y(n_378)
);

CKINVDCx5p33_ASAP7_75t_R g379 ( 
.A(n_125),
.Y(n_379)
);

INVx1_ASAP7_75t_L g380 ( 
.A(n_160),
.Y(n_380)
);

CKINVDCx5p33_ASAP7_75t_R g381 ( 
.A(n_120),
.Y(n_381)
);

CKINVDCx5p33_ASAP7_75t_R g382 ( 
.A(n_26),
.Y(n_382)
);

CKINVDCx20_ASAP7_75t_R g383 ( 
.A(n_43),
.Y(n_383)
);

CKINVDCx5p33_ASAP7_75t_R g384 ( 
.A(n_53),
.Y(n_384)
);

CKINVDCx5p33_ASAP7_75t_R g385 ( 
.A(n_111),
.Y(n_385)
);

INVx1_ASAP7_75t_SL g386 ( 
.A(n_164),
.Y(n_386)
);

BUFx3_ASAP7_75t_L g387 ( 
.A(n_26),
.Y(n_387)
);

INVx1_ASAP7_75t_SL g388 ( 
.A(n_71),
.Y(n_388)
);

CKINVDCx5p33_ASAP7_75t_R g389 ( 
.A(n_191),
.Y(n_389)
);

INVx1_ASAP7_75t_L g390 ( 
.A(n_9),
.Y(n_390)
);

INVx1_ASAP7_75t_L g391 ( 
.A(n_39),
.Y(n_391)
);

INVx1_ASAP7_75t_L g392 ( 
.A(n_31),
.Y(n_392)
);

CKINVDCx5p33_ASAP7_75t_R g393 ( 
.A(n_177),
.Y(n_393)
);

HB1xp67_ASAP7_75t_L g394 ( 
.A(n_1),
.Y(n_394)
);

INVx1_ASAP7_75t_L g395 ( 
.A(n_135),
.Y(n_395)
);

CKINVDCx5p33_ASAP7_75t_R g396 ( 
.A(n_163),
.Y(n_396)
);

BUFx6f_ASAP7_75t_L g397 ( 
.A(n_65),
.Y(n_397)
);

CKINVDCx5p33_ASAP7_75t_R g398 ( 
.A(n_208),
.Y(n_398)
);

CKINVDCx5p33_ASAP7_75t_R g399 ( 
.A(n_37),
.Y(n_399)
);

CKINVDCx5p33_ASAP7_75t_R g400 ( 
.A(n_42),
.Y(n_400)
);

INVx2_ASAP7_75t_L g401 ( 
.A(n_192),
.Y(n_401)
);

CKINVDCx5p33_ASAP7_75t_R g402 ( 
.A(n_79),
.Y(n_402)
);

CKINVDCx5p33_ASAP7_75t_R g403 ( 
.A(n_36),
.Y(n_403)
);

INVx1_ASAP7_75t_L g404 ( 
.A(n_49),
.Y(n_404)
);

CKINVDCx20_ASAP7_75t_R g405 ( 
.A(n_52),
.Y(n_405)
);

INVx1_ASAP7_75t_L g406 ( 
.A(n_80),
.Y(n_406)
);

INVx1_ASAP7_75t_SL g407 ( 
.A(n_21),
.Y(n_407)
);

CKINVDCx5p33_ASAP7_75t_R g408 ( 
.A(n_97),
.Y(n_408)
);

CKINVDCx5p33_ASAP7_75t_R g409 ( 
.A(n_14),
.Y(n_409)
);

CKINVDCx5p33_ASAP7_75t_R g410 ( 
.A(n_119),
.Y(n_410)
);

CKINVDCx5p33_ASAP7_75t_R g411 ( 
.A(n_2),
.Y(n_411)
);

BUFx3_ASAP7_75t_L g412 ( 
.A(n_22),
.Y(n_412)
);

INVx1_ASAP7_75t_L g413 ( 
.A(n_50),
.Y(n_413)
);

BUFx6f_ASAP7_75t_L g414 ( 
.A(n_16),
.Y(n_414)
);

CKINVDCx5p33_ASAP7_75t_R g415 ( 
.A(n_60),
.Y(n_415)
);

CKINVDCx16_ASAP7_75t_R g416 ( 
.A(n_67),
.Y(n_416)
);

CKINVDCx5p33_ASAP7_75t_R g417 ( 
.A(n_170),
.Y(n_417)
);

CKINVDCx5p33_ASAP7_75t_R g418 ( 
.A(n_21),
.Y(n_418)
);

CKINVDCx5p33_ASAP7_75t_R g419 ( 
.A(n_59),
.Y(n_419)
);

CKINVDCx5p33_ASAP7_75t_R g420 ( 
.A(n_27),
.Y(n_420)
);

CKINVDCx14_ASAP7_75t_R g421 ( 
.A(n_73),
.Y(n_421)
);

CKINVDCx5p33_ASAP7_75t_R g422 ( 
.A(n_139),
.Y(n_422)
);

CKINVDCx20_ASAP7_75t_R g423 ( 
.A(n_363),
.Y(n_423)
);

CKINVDCx5p33_ASAP7_75t_R g424 ( 
.A(n_216),
.Y(n_424)
);

INVx1_ASAP7_75t_L g425 ( 
.A(n_397),
.Y(n_425)
);

INVx1_ASAP7_75t_L g426 ( 
.A(n_397),
.Y(n_426)
);

INVx1_ASAP7_75t_L g427 ( 
.A(n_397),
.Y(n_427)
);

INVx1_ASAP7_75t_SL g428 ( 
.A(n_221),
.Y(n_428)
);

CKINVDCx5p33_ASAP7_75t_R g429 ( 
.A(n_218),
.Y(n_429)
);

INVx1_ASAP7_75t_L g430 ( 
.A(n_397),
.Y(n_430)
);

INVx1_ASAP7_75t_L g431 ( 
.A(n_397),
.Y(n_431)
);

NOR2xp33_ASAP7_75t_L g432 ( 
.A(n_258),
.B(n_0),
.Y(n_432)
);

CKINVDCx5p33_ASAP7_75t_R g433 ( 
.A(n_222),
.Y(n_433)
);

INVxp33_ASAP7_75t_L g434 ( 
.A(n_394),
.Y(n_434)
);

INVxp33_ASAP7_75t_SL g435 ( 
.A(n_231),
.Y(n_435)
);

CKINVDCx5p33_ASAP7_75t_R g436 ( 
.A(n_223),
.Y(n_436)
);

INVx1_ASAP7_75t_L g437 ( 
.A(n_397),
.Y(n_437)
);

INVx1_ASAP7_75t_SL g438 ( 
.A(n_243),
.Y(n_438)
);

INVxp67_ASAP7_75t_L g439 ( 
.A(n_214),
.Y(n_439)
);

INVx1_ASAP7_75t_L g440 ( 
.A(n_414),
.Y(n_440)
);

INVx1_ASAP7_75t_L g441 ( 
.A(n_414),
.Y(n_441)
);

CKINVDCx20_ASAP7_75t_R g442 ( 
.A(n_257),
.Y(n_442)
);

CKINVDCx5p33_ASAP7_75t_R g443 ( 
.A(n_224),
.Y(n_443)
);

INVx2_ASAP7_75t_L g444 ( 
.A(n_302),
.Y(n_444)
);

INVx1_ASAP7_75t_L g445 ( 
.A(n_414),
.Y(n_445)
);

CKINVDCx5p33_ASAP7_75t_R g446 ( 
.A(n_225),
.Y(n_446)
);

NOR2xp67_ASAP7_75t_L g447 ( 
.A(n_264),
.B(n_0),
.Y(n_447)
);

INVx1_ASAP7_75t_L g448 ( 
.A(n_414),
.Y(n_448)
);

CKINVDCx16_ASAP7_75t_R g449 ( 
.A(n_346),
.Y(n_449)
);

INVx1_ASAP7_75t_L g450 ( 
.A(n_414),
.Y(n_450)
);

INVx1_ASAP7_75t_L g451 ( 
.A(n_414),
.Y(n_451)
);

CKINVDCx20_ASAP7_75t_R g452 ( 
.A(n_421),
.Y(n_452)
);

INVx1_ASAP7_75t_L g453 ( 
.A(n_246),
.Y(n_453)
);

CKINVDCx20_ASAP7_75t_R g454 ( 
.A(n_226),
.Y(n_454)
);

CKINVDCx5p33_ASAP7_75t_R g455 ( 
.A(n_239),
.Y(n_455)
);

CKINVDCx20_ASAP7_75t_R g456 ( 
.A(n_248),
.Y(n_456)
);

HB1xp67_ASAP7_75t_L g457 ( 
.A(n_292),
.Y(n_457)
);

INVx1_ASAP7_75t_L g458 ( 
.A(n_246),
.Y(n_458)
);

CKINVDCx5p33_ASAP7_75t_R g459 ( 
.A(n_250),
.Y(n_459)
);

CKINVDCx5p33_ASAP7_75t_R g460 ( 
.A(n_253),
.Y(n_460)
);

CKINVDCx5p33_ASAP7_75t_R g461 ( 
.A(n_265),
.Y(n_461)
);

INVx1_ASAP7_75t_L g462 ( 
.A(n_255),
.Y(n_462)
);

INVxp67_ASAP7_75t_SL g463 ( 
.A(n_258),
.Y(n_463)
);

INVxp67_ASAP7_75t_SL g464 ( 
.A(n_261),
.Y(n_464)
);

HB1xp67_ASAP7_75t_L g465 ( 
.A(n_292),
.Y(n_465)
);

CKINVDCx5p33_ASAP7_75t_R g466 ( 
.A(n_266),
.Y(n_466)
);

INVx1_ASAP7_75t_L g467 ( 
.A(n_255),
.Y(n_467)
);

NOR2xp33_ASAP7_75t_L g468 ( 
.A(n_249),
.B(n_2),
.Y(n_468)
);

INVx1_ASAP7_75t_L g469 ( 
.A(n_293),
.Y(n_469)
);

NOR2xp33_ASAP7_75t_L g470 ( 
.A(n_249),
.B(n_5),
.Y(n_470)
);

INVx1_ASAP7_75t_L g471 ( 
.A(n_293),
.Y(n_471)
);

INVx1_ASAP7_75t_L g472 ( 
.A(n_299),
.Y(n_472)
);

CKINVDCx5p33_ASAP7_75t_R g473 ( 
.A(n_273),
.Y(n_473)
);

INVx1_ASAP7_75t_L g474 ( 
.A(n_299),
.Y(n_474)
);

CKINVDCx16_ASAP7_75t_R g475 ( 
.A(n_416),
.Y(n_475)
);

INVx1_ASAP7_75t_L g476 ( 
.A(n_374),
.Y(n_476)
);

NOR2xp33_ASAP7_75t_R g477 ( 
.A(n_274),
.B(n_90),
.Y(n_477)
);

CKINVDCx5p33_ASAP7_75t_R g478 ( 
.A(n_275),
.Y(n_478)
);

INVx1_ASAP7_75t_L g479 ( 
.A(n_374),
.Y(n_479)
);

INVx1_ASAP7_75t_L g480 ( 
.A(n_230),
.Y(n_480)
);

NOR2xp33_ASAP7_75t_L g481 ( 
.A(n_215),
.B(n_6),
.Y(n_481)
);

INVxp67_ASAP7_75t_L g482 ( 
.A(n_214),
.Y(n_482)
);

NAND2xp5_ASAP7_75t_L g483 ( 
.A(n_233),
.B(n_7),
.Y(n_483)
);

CKINVDCx20_ASAP7_75t_R g484 ( 
.A(n_279),
.Y(n_484)
);

INVxp67_ASAP7_75t_SL g485 ( 
.A(n_261),
.Y(n_485)
);

INVxp33_ASAP7_75t_SL g486 ( 
.A(n_232),
.Y(n_486)
);

INVx1_ASAP7_75t_L g487 ( 
.A(n_230),
.Y(n_487)
);

CKINVDCx5p33_ASAP7_75t_R g488 ( 
.A(n_280),
.Y(n_488)
);

CKINVDCx5p33_ASAP7_75t_R g489 ( 
.A(n_282),
.Y(n_489)
);

INVx1_ASAP7_75t_L g490 ( 
.A(n_230),
.Y(n_490)
);

NOR2xp33_ASAP7_75t_L g491 ( 
.A(n_215),
.B(n_217),
.Y(n_491)
);

NOR2xp33_ASAP7_75t_L g492 ( 
.A(n_217),
.B(n_9),
.Y(n_492)
);

NOR2xp33_ASAP7_75t_L g493 ( 
.A(n_235),
.B(n_10),
.Y(n_493)
);

CKINVDCx5p33_ASAP7_75t_R g494 ( 
.A(n_284),
.Y(n_494)
);

CKINVDCx5p33_ASAP7_75t_R g495 ( 
.A(n_288),
.Y(n_495)
);

BUFx3_ASAP7_75t_L g496 ( 
.A(n_323),
.Y(n_496)
);

CKINVDCx20_ASAP7_75t_R g497 ( 
.A(n_289),
.Y(n_497)
);

INVx1_ASAP7_75t_L g498 ( 
.A(n_387),
.Y(n_498)
);

INVx1_ASAP7_75t_L g499 ( 
.A(n_387),
.Y(n_499)
);

INVx1_ASAP7_75t_L g500 ( 
.A(n_387),
.Y(n_500)
);

INVx1_ASAP7_75t_L g501 ( 
.A(n_412),
.Y(n_501)
);

CKINVDCx5p33_ASAP7_75t_R g502 ( 
.A(n_291),
.Y(n_502)
);

INVx1_ASAP7_75t_L g503 ( 
.A(n_412),
.Y(n_503)
);

AND2x2_ASAP7_75t_L g504 ( 
.A(n_412),
.B(n_416),
.Y(n_504)
);

CKINVDCx20_ASAP7_75t_R g505 ( 
.A(n_298),
.Y(n_505)
);

CKINVDCx5p33_ASAP7_75t_R g506 ( 
.A(n_307),
.Y(n_506)
);

HB1xp67_ASAP7_75t_L g507 ( 
.A(n_251),
.Y(n_507)
);

INVx1_ASAP7_75t_L g508 ( 
.A(n_220),
.Y(n_508)
);

INVx1_ASAP7_75t_L g509 ( 
.A(n_220),
.Y(n_509)
);

INVx2_ASAP7_75t_L g510 ( 
.A(n_302),
.Y(n_510)
);

BUFx10_ASAP7_75t_L g511 ( 
.A(n_302),
.Y(n_511)
);

INVx1_ASAP7_75t_L g512 ( 
.A(n_227),
.Y(n_512)
);

NAND2xp5_ASAP7_75t_L g513 ( 
.A(n_233),
.B(n_11),
.Y(n_513)
);

INVx1_ASAP7_75t_L g514 ( 
.A(n_227),
.Y(n_514)
);

INVxp67_ASAP7_75t_L g515 ( 
.A(n_237),
.Y(n_515)
);

NOR2xp67_ASAP7_75t_L g516 ( 
.A(n_264),
.B(n_13),
.Y(n_516)
);

CKINVDCx5p33_ASAP7_75t_R g517 ( 
.A(n_309),
.Y(n_517)
);

BUFx3_ASAP7_75t_L g518 ( 
.A(n_323),
.Y(n_518)
);

NOR2xp33_ASAP7_75t_L g519 ( 
.A(n_235),
.B(n_13),
.Y(n_519)
);

INVx1_ASAP7_75t_L g520 ( 
.A(n_237),
.Y(n_520)
);

INVx1_ASAP7_75t_L g521 ( 
.A(n_241),
.Y(n_521)
);

CKINVDCx20_ASAP7_75t_R g522 ( 
.A(n_310),
.Y(n_522)
);

CKINVDCx16_ASAP7_75t_R g523 ( 
.A(n_228),
.Y(n_523)
);

NOR2xp33_ASAP7_75t_L g524 ( 
.A(n_236),
.B(n_238),
.Y(n_524)
);

INVxp67_ASAP7_75t_SL g525 ( 
.A(n_325),
.Y(n_525)
);

CKINVDCx5p33_ASAP7_75t_R g526 ( 
.A(n_311),
.Y(n_526)
);

INVx1_ASAP7_75t_L g527 ( 
.A(n_241),
.Y(n_527)
);

INVxp67_ASAP7_75t_SL g528 ( 
.A(n_359),
.Y(n_528)
);

CKINVDCx20_ASAP7_75t_R g529 ( 
.A(n_313),
.Y(n_529)
);

NOR2xp33_ASAP7_75t_L g530 ( 
.A(n_236),
.B(n_15),
.Y(n_530)
);

INVx1_ASAP7_75t_SL g531 ( 
.A(n_260),
.Y(n_531)
);

BUFx6f_ASAP7_75t_L g532 ( 
.A(n_444),
.Y(n_532)
);

INVx2_ASAP7_75t_L g533 ( 
.A(n_444),
.Y(n_533)
);

INVx2_ASAP7_75t_L g534 ( 
.A(n_444),
.Y(n_534)
);

AND2x4_ASAP7_75t_L g535 ( 
.A(n_425),
.B(n_234),
.Y(n_535)
);

AND2x2_ASAP7_75t_L g536 ( 
.A(n_480),
.B(n_238),
.Y(n_536)
);

AND2x2_ASAP7_75t_L g537 ( 
.A(n_480),
.B(n_487),
.Y(n_537)
);

INVx3_ASAP7_75t_L g538 ( 
.A(n_510),
.Y(n_538)
);

OA21x2_ASAP7_75t_L g539 ( 
.A1(n_425),
.A2(n_245),
.B(n_244),
.Y(n_539)
);

INVx3_ASAP7_75t_L g540 ( 
.A(n_510),
.Y(n_540)
);

AND2x2_ASAP7_75t_L g541 ( 
.A(n_487),
.B(n_240),
.Y(n_541)
);

INVx1_ASAP7_75t_L g542 ( 
.A(n_426),
.Y(n_542)
);

INVx1_ASAP7_75t_L g543 ( 
.A(n_426),
.Y(n_543)
);

BUFx6f_ASAP7_75t_L g544 ( 
.A(n_510),
.Y(n_544)
);

AND2x4_ASAP7_75t_L g545 ( 
.A(n_427),
.B(n_430),
.Y(n_545)
);

NAND2xp5_ASAP7_75t_L g546 ( 
.A(n_491),
.B(n_316),
.Y(n_546)
);

CKINVDCx11_ASAP7_75t_R g547 ( 
.A(n_442),
.Y(n_547)
);

AND2x4_ASAP7_75t_L g548 ( 
.A(n_427),
.B(n_234),
.Y(n_548)
);

OA21x2_ASAP7_75t_L g549 ( 
.A1(n_430),
.A2(n_245),
.B(n_244),
.Y(n_549)
);

INVx3_ASAP7_75t_L g550 ( 
.A(n_511),
.Y(n_550)
);

INVx2_ASAP7_75t_L g551 ( 
.A(n_431),
.Y(n_551)
);

INVx1_ASAP7_75t_L g552 ( 
.A(n_431),
.Y(n_552)
);

AND2x2_ASAP7_75t_L g553 ( 
.A(n_490),
.B(n_240),
.Y(n_553)
);

BUFx3_ASAP7_75t_L g554 ( 
.A(n_511),
.Y(n_554)
);

AND2x6_ASAP7_75t_L g555 ( 
.A(n_437),
.B(n_302),
.Y(n_555)
);

INVx3_ASAP7_75t_L g556 ( 
.A(n_511),
.Y(n_556)
);

AND2x4_ASAP7_75t_L g557 ( 
.A(n_437),
.B(n_252),
.Y(n_557)
);

BUFx2_ASAP7_75t_L g558 ( 
.A(n_504),
.Y(n_558)
);

INVx1_ASAP7_75t_L g559 ( 
.A(n_440),
.Y(n_559)
);

NAND2xp5_ASAP7_75t_L g560 ( 
.A(n_524),
.B(n_422),
.Y(n_560)
);

INVx1_ASAP7_75t_L g561 ( 
.A(n_440),
.Y(n_561)
);

NAND2xp5_ASAP7_75t_L g562 ( 
.A(n_464),
.B(n_320),
.Y(n_562)
);

INVx1_ASAP7_75t_L g563 ( 
.A(n_441),
.Y(n_563)
);

INVx2_ASAP7_75t_L g564 ( 
.A(n_441),
.Y(n_564)
);

CKINVDCx20_ASAP7_75t_R g565 ( 
.A(n_452),
.Y(n_565)
);

INVx2_ASAP7_75t_SL g566 ( 
.A(n_511),
.Y(n_566)
);

BUFx2_ASAP7_75t_L g567 ( 
.A(n_504),
.Y(n_567)
);

INVx1_ASAP7_75t_L g568 ( 
.A(n_445),
.Y(n_568)
);

OAI22xp5_ASAP7_75t_L g569 ( 
.A1(n_432),
.A2(n_285),
.B1(n_370),
.B2(n_315),
.Y(n_569)
);

INVx1_ASAP7_75t_L g570 ( 
.A(n_445),
.Y(n_570)
);

INVx1_ASAP7_75t_L g571 ( 
.A(n_448),
.Y(n_571)
);

INVx2_ASAP7_75t_L g572 ( 
.A(n_448),
.Y(n_572)
);

AND2x4_ASAP7_75t_L g573 ( 
.A(n_450),
.B(n_252),
.Y(n_573)
);

HB1xp67_ASAP7_75t_L g574 ( 
.A(n_457),
.Y(n_574)
);

OAI22xp5_ASAP7_75t_L g575 ( 
.A1(n_475),
.A2(n_405),
.B1(n_383),
.B2(n_268),
.Y(n_575)
);

NAND2xp5_ASAP7_75t_SL g576 ( 
.A(n_449),
.B(n_228),
.Y(n_576)
);

INVx2_ASAP7_75t_L g577 ( 
.A(n_450),
.Y(n_577)
);

CKINVDCx20_ASAP7_75t_R g578 ( 
.A(n_423),
.Y(n_578)
);

BUFx6f_ASAP7_75t_L g579 ( 
.A(n_451),
.Y(n_579)
);

INVx3_ASAP7_75t_L g580 ( 
.A(n_451),
.Y(n_580)
);

INVx1_ASAP7_75t_L g581 ( 
.A(n_508),
.Y(n_581)
);

INVx2_ASAP7_75t_L g582 ( 
.A(n_453),
.Y(n_582)
);

AND2x4_ASAP7_75t_L g583 ( 
.A(n_496),
.B(n_290),
.Y(n_583)
);

INVx1_ASAP7_75t_L g584 ( 
.A(n_508),
.Y(n_584)
);

INVx3_ASAP7_75t_L g585 ( 
.A(n_453),
.Y(n_585)
);

INVx2_ASAP7_75t_L g586 ( 
.A(n_458),
.Y(n_586)
);

AND2x2_ASAP7_75t_L g587 ( 
.A(n_490),
.B(n_242),
.Y(n_587)
);

NAND2xp5_ASAP7_75t_L g588 ( 
.A(n_485),
.B(n_328),
.Y(n_588)
);

INVx3_ASAP7_75t_L g589 ( 
.A(n_458),
.Y(n_589)
);

INVx2_ASAP7_75t_L g590 ( 
.A(n_462),
.Y(n_590)
);

INVx1_ASAP7_75t_L g591 ( 
.A(n_509),
.Y(n_591)
);

AND2x4_ASAP7_75t_L g592 ( 
.A(n_496),
.B(n_290),
.Y(n_592)
);

BUFx6f_ASAP7_75t_L g593 ( 
.A(n_462),
.Y(n_593)
);

AND2x4_ASAP7_75t_L g594 ( 
.A(n_496),
.B(n_401),
.Y(n_594)
);

INVx1_ASAP7_75t_L g595 ( 
.A(n_509),
.Y(n_595)
);

INVx2_ASAP7_75t_L g596 ( 
.A(n_467),
.Y(n_596)
);

AND2x4_ASAP7_75t_L g597 ( 
.A(n_518),
.B(n_401),
.Y(n_597)
);

NAND2x1p5_ASAP7_75t_L g598 ( 
.A(n_481),
.B(n_302),
.Y(n_598)
);

INVx1_ASAP7_75t_L g599 ( 
.A(n_512),
.Y(n_599)
);

INVx1_ASAP7_75t_L g600 ( 
.A(n_512),
.Y(n_600)
);

NAND2xp5_ASAP7_75t_L g601 ( 
.A(n_468),
.B(n_329),
.Y(n_601)
);

OR2x2_ASAP7_75t_L g602 ( 
.A(n_449),
.B(n_364),
.Y(n_602)
);

NAND2xp5_ASAP7_75t_L g603 ( 
.A(n_470),
.B(n_330),
.Y(n_603)
);

BUFx6f_ASAP7_75t_L g604 ( 
.A(n_467),
.Y(n_604)
);

INVx2_ASAP7_75t_L g605 ( 
.A(n_469),
.Y(n_605)
);

INVx5_ASAP7_75t_L g606 ( 
.A(n_518),
.Y(n_606)
);

BUFx6f_ASAP7_75t_L g607 ( 
.A(n_469),
.Y(n_607)
);

AND2x6_ASAP7_75t_L g608 ( 
.A(n_492),
.B(n_302),
.Y(n_608)
);

NAND2xp5_ASAP7_75t_L g609 ( 
.A(n_498),
.B(n_333),
.Y(n_609)
);

INVx2_ASAP7_75t_L g610 ( 
.A(n_471),
.Y(n_610)
);

INVx1_ASAP7_75t_L g611 ( 
.A(n_514),
.Y(n_611)
);

AND2x4_ASAP7_75t_L g612 ( 
.A(n_518),
.B(n_242),
.Y(n_612)
);

INVx1_ASAP7_75t_L g613 ( 
.A(n_514),
.Y(n_613)
);

AND2x4_ASAP7_75t_L g614 ( 
.A(n_498),
.B(n_254),
.Y(n_614)
);

INVx1_ASAP7_75t_L g615 ( 
.A(n_520),
.Y(n_615)
);

BUFx6f_ASAP7_75t_L g616 ( 
.A(n_471),
.Y(n_616)
);

INVx1_ASAP7_75t_L g617 ( 
.A(n_520),
.Y(n_617)
);

INVx1_ASAP7_75t_L g618 ( 
.A(n_521),
.Y(n_618)
);

INVx2_ASAP7_75t_L g619 ( 
.A(n_545),
.Y(n_619)
);

INVx2_ASAP7_75t_SL g620 ( 
.A(n_558),
.Y(n_620)
);

INVx2_ASAP7_75t_L g621 ( 
.A(n_545),
.Y(n_621)
);

NAND2xp5_ASAP7_75t_SL g622 ( 
.A(n_558),
.B(n_523),
.Y(n_622)
);

NAND2xp5_ASAP7_75t_SL g623 ( 
.A(n_558),
.B(n_523),
.Y(n_623)
);

INVx2_ASAP7_75t_L g624 ( 
.A(n_545),
.Y(n_624)
);

NOR2xp33_ASAP7_75t_L g625 ( 
.A(n_546),
.B(n_435),
.Y(n_625)
);

INVx1_ASAP7_75t_L g626 ( 
.A(n_539),
.Y(n_626)
);

INVx1_ASAP7_75t_L g627 ( 
.A(n_539),
.Y(n_627)
);

INVx3_ASAP7_75t_L g628 ( 
.A(n_532),
.Y(n_628)
);

BUFx6f_ASAP7_75t_L g629 ( 
.A(n_532),
.Y(n_629)
);

INVxp33_ASAP7_75t_L g630 ( 
.A(n_574),
.Y(n_630)
);

BUFx3_ASAP7_75t_L g631 ( 
.A(n_539),
.Y(n_631)
);

OR2x2_ASAP7_75t_L g632 ( 
.A(n_602),
.B(n_475),
.Y(n_632)
);

AND2x2_ASAP7_75t_L g633 ( 
.A(n_567),
.B(n_499),
.Y(n_633)
);

INVx1_ASAP7_75t_L g634 ( 
.A(n_539),
.Y(n_634)
);

INVx1_ASAP7_75t_L g635 ( 
.A(n_539),
.Y(n_635)
);

NAND2xp5_ASAP7_75t_L g636 ( 
.A(n_566),
.B(n_546),
.Y(n_636)
);

INVx1_ASAP7_75t_L g637 ( 
.A(n_539),
.Y(n_637)
);

HB1xp67_ASAP7_75t_L g638 ( 
.A(n_574),
.Y(n_638)
);

HB1xp67_ASAP7_75t_SL g639 ( 
.A(n_575),
.Y(n_639)
);

AOI22xp33_ASAP7_75t_L g640 ( 
.A1(n_608),
.A2(n_463),
.B1(n_519),
.B2(n_493),
.Y(n_640)
);

NAND2xp5_ASAP7_75t_SL g641 ( 
.A(n_567),
.B(n_424),
.Y(n_641)
);

NOR2xp33_ASAP7_75t_L g642 ( 
.A(n_560),
.B(n_486),
.Y(n_642)
);

INVx2_ASAP7_75t_L g643 ( 
.A(n_545),
.Y(n_643)
);

OR2x2_ASAP7_75t_L g644 ( 
.A(n_602),
.B(n_428),
.Y(n_644)
);

AND2x2_ASAP7_75t_L g645 ( 
.A(n_567),
.B(n_499),
.Y(n_645)
);

INVx1_ASAP7_75t_L g646 ( 
.A(n_549),
.Y(n_646)
);

NAND2xp5_ASAP7_75t_L g647 ( 
.A(n_566),
.B(n_429),
.Y(n_647)
);

NAND2xp5_ASAP7_75t_L g648 ( 
.A(n_566),
.B(n_433),
.Y(n_648)
);

NAND2xp5_ASAP7_75t_L g649 ( 
.A(n_560),
.B(n_436),
.Y(n_649)
);

NAND3xp33_ASAP7_75t_L g650 ( 
.A(n_536),
.B(n_530),
.C(n_513),
.Y(n_650)
);

INVx3_ASAP7_75t_L g651 ( 
.A(n_532),
.Y(n_651)
);

INVx4_ASAP7_75t_L g652 ( 
.A(n_550),
.Y(n_652)
);

NAND2xp5_ASAP7_75t_SL g653 ( 
.A(n_602),
.B(n_443),
.Y(n_653)
);

INVx3_ASAP7_75t_L g654 ( 
.A(n_532),
.Y(n_654)
);

INVx1_ASAP7_75t_L g655 ( 
.A(n_549),
.Y(n_655)
);

INVx1_ASAP7_75t_L g656 ( 
.A(n_549),
.Y(n_656)
);

INVx2_ASAP7_75t_L g657 ( 
.A(n_545),
.Y(n_657)
);

NOR2xp33_ASAP7_75t_L g658 ( 
.A(n_562),
.B(n_446),
.Y(n_658)
);

INVxp33_ASAP7_75t_L g659 ( 
.A(n_569),
.Y(n_659)
);

INVx1_ASAP7_75t_L g660 ( 
.A(n_549),
.Y(n_660)
);

NOR2xp33_ASAP7_75t_L g661 ( 
.A(n_562),
.B(n_455),
.Y(n_661)
);

BUFx4f_ASAP7_75t_L g662 ( 
.A(n_549),
.Y(n_662)
);

INVx2_ASAP7_75t_SL g663 ( 
.A(n_588),
.Y(n_663)
);

INVx1_ASAP7_75t_L g664 ( 
.A(n_549),
.Y(n_664)
);

HB1xp67_ASAP7_75t_L g665 ( 
.A(n_588),
.Y(n_665)
);

INVx2_ASAP7_75t_L g666 ( 
.A(n_551),
.Y(n_666)
);

INVx2_ASAP7_75t_L g667 ( 
.A(n_551),
.Y(n_667)
);

INVx2_ASAP7_75t_L g668 ( 
.A(n_551),
.Y(n_668)
);

NAND2xp5_ASAP7_75t_SL g669 ( 
.A(n_576),
.B(n_459),
.Y(n_669)
);

NOR2x1p5_ASAP7_75t_L g670 ( 
.A(n_601),
.B(n_247),
.Y(n_670)
);

INVx2_ASAP7_75t_L g671 ( 
.A(n_564),
.Y(n_671)
);

INVx2_ASAP7_75t_L g672 ( 
.A(n_564),
.Y(n_672)
);

BUFx3_ASAP7_75t_L g673 ( 
.A(n_606),
.Y(n_673)
);

NAND2xp33_ASAP7_75t_R g674 ( 
.A(n_601),
.B(n_460),
.Y(n_674)
);

INVx1_ASAP7_75t_L g675 ( 
.A(n_537),
.Y(n_675)
);

BUFx3_ASAP7_75t_L g676 ( 
.A(n_606),
.Y(n_676)
);

OR2x2_ASAP7_75t_L g677 ( 
.A(n_609),
.B(n_438),
.Y(n_677)
);

INVx2_ASAP7_75t_L g678 ( 
.A(n_564),
.Y(n_678)
);

INVx2_ASAP7_75t_L g679 ( 
.A(n_572),
.Y(n_679)
);

AOI22xp33_ASAP7_75t_L g680 ( 
.A1(n_608),
.A2(n_483),
.B1(n_528),
.B2(n_525),
.Y(n_680)
);

BUFx3_ASAP7_75t_L g681 ( 
.A(n_606),
.Y(n_681)
);

AND2x2_ASAP7_75t_L g682 ( 
.A(n_537),
.B(n_500),
.Y(n_682)
);

INVx2_ASAP7_75t_L g683 ( 
.A(n_572),
.Y(n_683)
);

AOI22xp33_ASAP7_75t_L g684 ( 
.A1(n_608),
.A2(n_447),
.B1(n_516),
.B2(n_364),
.Y(n_684)
);

INVx1_ASAP7_75t_L g685 ( 
.A(n_537),
.Y(n_685)
);

INVx5_ASAP7_75t_L g686 ( 
.A(n_555),
.Y(n_686)
);

INVx2_ASAP7_75t_L g687 ( 
.A(n_572),
.Y(n_687)
);

BUFx4f_ASAP7_75t_L g688 ( 
.A(n_608),
.Y(n_688)
);

INVx2_ASAP7_75t_L g689 ( 
.A(n_577),
.Y(n_689)
);

INVx2_ASAP7_75t_L g690 ( 
.A(n_577),
.Y(n_690)
);

INVx3_ASAP7_75t_L g691 ( 
.A(n_532),
.Y(n_691)
);

INVx2_ASAP7_75t_L g692 ( 
.A(n_577),
.Y(n_692)
);

INVx1_ASAP7_75t_L g693 ( 
.A(n_542),
.Y(n_693)
);

INVx2_ASAP7_75t_L g694 ( 
.A(n_542),
.Y(n_694)
);

BUFx6f_ASAP7_75t_SL g695 ( 
.A(n_612),
.Y(n_695)
);

NOR2xp33_ASAP7_75t_L g696 ( 
.A(n_603),
.B(n_461),
.Y(n_696)
);

INVx1_ASAP7_75t_L g697 ( 
.A(n_543),
.Y(n_697)
);

INVx5_ASAP7_75t_L g698 ( 
.A(n_555),
.Y(n_698)
);

INVx1_ASAP7_75t_L g699 ( 
.A(n_543),
.Y(n_699)
);

BUFx3_ASAP7_75t_L g700 ( 
.A(n_606),
.Y(n_700)
);

INVx1_ASAP7_75t_L g701 ( 
.A(n_552),
.Y(n_701)
);

NOR2xp33_ASAP7_75t_L g702 ( 
.A(n_603),
.B(n_466),
.Y(n_702)
);

AOI22xp33_ASAP7_75t_L g703 ( 
.A1(n_608),
.A2(n_447),
.B1(n_516),
.B2(n_465),
.Y(n_703)
);

INVx1_ASAP7_75t_L g704 ( 
.A(n_552),
.Y(n_704)
);

NAND2xp5_ASAP7_75t_SL g705 ( 
.A(n_576),
.B(n_473),
.Y(n_705)
);

NAND3xp33_ASAP7_75t_L g706 ( 
.A(n_536),
.B(n_501),
.C(n_500),
.Y(n_706)
);

BUFx6f_ASAP7_75t_L g707 ( 
.A(n_532),
.Y(n_707)
);

NAND2xp5_ASAP7_75t_SL g708 ( 
.A(n_609),
.B(n_478),
.Y(n_708)
);

AOI22xp33_ASAP7_75t_L g709 ( 
.A1(n_608),
.A2(n_434),
.B1(n_262),
.B2(n_270),
.Y(n_709)
);

AND2x6_ASAP7_75t_L g710 ( 
.A(n_550),
.B(n_357),
.Y(n_710)
);

INVxp67_ASAP7_75t_L g711 ( 
.A(n_569),
.Y(n_711)
);

CKINVDCx5p33_ASAP7_75t_R g712 ( 
.A(n_547),
.Y(n_712)
);

INVx2_ASAP7_75t_L g713 ( 
.A(n_559),
.Y(n_713)
);

NAND2xp5_ASAP7_75t_L g714 ( 
.A(n_550),
.B(n_488),
.Y(n_714)
);

OR2x6_ASAP7_75t_L g715 ( 
.A(n_612),
.B(n_378),
.Y(n_715)
);

INVx1_ASAP7_75t_L g716 ( 
.A(n_559),
.Y(n_716)
);

INVx2_ASAP7_75t_L g717 ( 
.A(n_561),
.Y(n_717)
);

INVx2_ASAP7_75t_L g718 ( 
.A(n_561),
.Y(n_718)
);

INVx3_ASAP7_75t_L g719 ( 
.A(n_532),
.Y(n_719)
);

INVx4_ASAP7_75t_L g720 ( 
.A(n_550),
.Y(n_720)
);

INVx2_ASAP7_75t_L g721 ( 
.A(n_563),
.Y(n_721)
);

NAND2xp5_ASAP7_75t_SL g722 ( 
.A(n_612),
.B(n_489),
.Y(n_722)
);

BUFx10_ASAP7_75t_L g723 ( 
.A(n_612),
.Y(n_723)
);

NAND2xp5_ASAP7_75t_L g724 ( 
.A(n_550),
.B(n_494),
.Y(n_724)
);

NAND2xp5_ASAP7_75t_SL g725 ( 
.A(n_612),
.B(n_495),
.Y(n_725)
);

INVx1_ASAP7_75t_L g726 ( 
.A(n_563),
.Y(n_726)
);

INVxp67_ASAP7_75t_L g727 ( 
.A(n_575),
.Y(n_727)
);

INVx1_ASAP7_75t_L g728 ( 
.A(n_568),
.Y(n_728)
);

NAND3xp33_ASAP7_75t_L g729 ( 
.A(n_536),
.B(n_503),
.C(n_501),
.Y(n_729)
);

INVx1_ASAP7_75t_L g730 ( 
.A(n_568),
.Y(n_730)
);

INVx3_ASAP7_75t_L g731 ( 
.A(n_532),
.Y(n_731)
);

NOR2x1p5_ASAP7_75t_L g732 ( 
.A(n_581),
.B(n_247),
.Y(n_732)
);

INVx1_ASAP7_75t_L g733 ( 
.A(n_570),
.Y(n_733)
);

INVx1_ASAP7_75t_L g734 ( 
.A(n_570),
.Y(n_734)
);

INVx1_ASAP7_75t_L g735 ( 
.A(n_571),
.Y(n_735)
);

NAND2xp33_ASAP7_75t_L g736 ( 
.A(n_608),
.B(n_502),
.Y(n_736)
);

NOR2xp33_ASAP7_75t_L g737 ( 
.A(n_556),
.B(n_506),
.Y(n_737)
);

INVx1_ASAP7_75t_L g738 ( 
.A(n_571),
.Y(n_738)
);

INVx2_ASAP7_75t_L g739 ( 
.A(n_533),
.Y(n_739)
);

INVx1_ASAP7_75t_L g740 ( 
.A(n_535),
.Y(n_740)
);

OR2x6_ASAP7_75t_L g741 ( 
.A(n_583),
.B(n_378),
.Y(n_741)
);

AND2x6_ASAP7_75t_L g742 ( 
.A(n_556),
.B(n_357),
.Y(n_742)
);

INVxp67_ASAP7_75t_L g743 ( 
.A(n_541),
.Y(n_743)
);

INVx1_ASAP7_75t_L g744 ( 
.A(n_535),
.Y(n_744)
);

INVx1_ASAP7_75t_L g745 ( 
.A(n_535),
.Y(n_745)
);

INVx2_ASAP7_75t_SL g746 ( 
.A(n_583),
.Y(n_746)
);

AOI22xp33_ASAP7_75t_L g747 ( 
.A1(n_608),
.A2(n_270),
.B1(n_272),
.B2(n_262),
.Y(n_747)
);

INVx1_ASAP7_75t_L g748 ( 
.A(n_535),
.Y(n_748)
);

INVx2_ASAP7_75t_SL g749 ( 
.A(n_583),
.Y(n_749)
);

BUFx6f_ASAP7_75t_L g750 ( 
.A(n_544),
.Y(n_750)
);

INVx1_ASAP7_75t_L g751 ( 
.A(n_535),
.Y(n_751)
);

AND2x6_ASAP7_75t_L g752 ( 
.A(n_556),
.B(n_357),
.Y(n_752)
);

INVx3_ASAP7_75t_L g753 ( 
.A(n_544),
.Y(n_753)
);

BUFx3_ASAP7_75t_L g754 ( 
.A(n_606),
.Y(n_754)
);

INVx1_ASAP7_75t_L g755 ( 
.A(n_548),
.Y(n_755)
);

AOI22xp33_ASAP7_75t_L g756 ( 
.A1(n_608),
.A2(n_278),
.B1(n_297),
.B2(n_272),
.Y(n_756)
);

INVx2_ASAP7_75t_L g757 ( 
.A(n_533),
.Y(n_757)
);

HB1xp67_ASAP7_75t_L g758 ( 
.A(n_541),
.Y(n_758)
);

INVx1_ASAP7_75t_L g759 ( 
.A(n_548),
.Y(n_759)
);

NOR2xp33_ASAP7_75t_L g760 ( 
.A(n_556),
.B(n_517),
.Y(n_760)
);

OR2x6_ASAP7_75t_L g761 ( 
.A(n_583),
.B(n_254),
.Y(n_761)
);

INVx2_ASAP7_75t_L g762 ( 
.A(n_533),
.Y(n_762)
);

NAND2xp5_ASAP7_75t_SL g763 ( 
.A(n_583),
.B(n_526),
.Y(n_763)
);

OAI22x1_ASAP7_75t_L g764 ( 
.A1(n_598),
.A2(n_531),
.B1(n_407),
.B2(n_388),
.Y(n_764)
);

INVx2_ASAP7_75t_L g765 ( 
.A(n_534),
.Y(n_765)
);

AND2x6_ASAP7_75t_L g766 ( 
.A(n_556),
.B(n_357),
.Y(n_766)
);

INVx1_ASAP7_75t_L g767 ( 
.A(n_548),
.Y(n_767)
);

NOR2xp33_ASAP7_75t_L g768 ( 
.A(n_598),
.B(n_454),
.Y(n_768)
);

INVx1_ASAP7_75t_L g769 ( 
.A(n_548),
.Y(n_769)
);

INVx2_ASAP7_75t_L g770 ( 
.A(n_534),
.Y(n_770)
);

CKINVDCx5p33_ASAP7_75t_R g771 ( 
.A(n_547),
.Y(n_771)
);

INVx2_ASAP7_75t_L g772 ( 
.A(n_694),
.Y(n_772)
);

INVx1_ASAP7_75t_L g773 ( 
.A(n_675),
.Y(n_773)
);

INVx8_ASAP7_75t_L g774 ( 
.A(n_695),
.Y(n_774)
);

NAND2xp5_ASAP7_75t_L g775 ( 
.A(n_663),
.B(n_608),
.Y(n_775)
);

AND2x6_ASAP7_75t_L g776 ( 
.A(n_631),
.B(n_256),
.Y(n_776)
);

NAND2xp5_ASAP7_75t_SL g777 ( 
.A(n_663),
.B(n_554),
.Y(n_777)
);

INVx2_ASAP7_75t_L g778 ( 
.A(n_694),
.Y(n_778)
);

AOI221xp5_ASAP7_75t_L g779 ( 
.A1(n_659),
.A2(n_229),
.B1(n_439),
.B2(n_482),
.C(n_515),
.Y(n_779)
);

NAND2xp5_ASAP7_75t_L g780 ( 
.A(n_696),
.B(n_598),
.Y(n_780)
);

NOR2xp33_ASAP7_75t_L g781 ( 
.A(n_625),
.B(n_456),
.Y(n_781)
);

INVx2_ASAP7_75t_L g782 ( 
.A(n_713),
.Y(n_782)
);

NAND2xp5_ASAP7_75t_L g783 ( 
.A(n_702),
.B(n_598),
.Y(n_783)
);

NAND2xp5_ASAP7_75t_L g784 ( 
.A(n_636),
.B(n_592),
.Y(n_784)
);

NAND2xp5_ASAP7_75t_L g785 ( 
.A(n_658),
.B(n_592),
.Y(n_785)
);

NAND2xp5_ASAP7_75t_SL g786 ( 
.A(n_688),
.B(n_554),
.Y(n_786)
);

NAND2xp5_ASAP7_75t_L g787 ( 
.A(n_661),
.B(n_592),
.Y(n_787)
);

NOR2xp33_ASAP7_75t_L g788 ( 
.A(n_642),
.B(n_484),
.Y(n_788)
);

NAND2xp5_ASAP7_75t_L g789 ( 
.A(n_665),
.B(n_592),
.Y(n_789)
);

HB1xp67_ASAP7_75t_L g790 ( 
.A(n_638),
.Y(n_790)
);

AND2x2_ASAP7_75t_L g791 ( 
.A(n_620),
.B(n_758),
.Y(n_791)
);

NAND2xp5_ASAP7_75t_L g792 ( 
.A(n_737),
.B(n_592),
.Y(n_792)
);

INVx1_ASAP7_75t_L g793 ( 
.A(n_675),
.Y(n_793)
);

AND2x6_ASAP7_75t_SL g794 ( 
.A(n_768),
.B(n_278),
.Y(n_794)
);

NAND2xp5_ASAP7_75t_L g795 ( 
.A(n_760),
.B(n_594),
.Y(n_795)
);

BUFx6f_ASAP7_75t_L g796 ( 
.A(n_723),
.Y(n_796)
);

NOR2x1p5_ASAP7_75t_L g797 ( 
.A(n_644),
.B(n_219),
.Y(n_797)
);

NOR2xp33_ASAP7_75t_L g798 ( 
.A(n_649),
.B(n_497),
.Y(n_798)
);

NAND2xp5_ASAP7_75t_L g799 ( 
.A(n_743),
.B(n_594),
.Y(n_799)
);

INVx1_ASAP7_75t_L g800 ( 
.A(n_685),
.Y(n_800)
);

NAND2xp5_ASAP7_75t_L g801 ( 
.A(n_685),
.B(n_594),
.Y(n_801)
);

CKINVDCx5p33_ASAP7_75t_R g802 ( 
.A(n_712),
.Y(n_802)
);

INVx1_ASAP7_75t_L g803 ( 
.A(n_746),
.Y(n_803)
);

NOR3xp33_ASAP7_75t_L g804 ( 
.A(n_622),
.B(n_623),
.C(n_653),
.Y(n_804)
);

INVx1_ASAP7_75t_L g805 ( 
.A(n_746),
.Y(n_805)
);

INVx1_ASAP7_75t_L g806 ( 
.A(n_749),
.Y(n_806)
);

AO221x1_ASAP7_75t_L g807 ( 
.A1(n_764),
.A2(n_357),
.B1(n_342),
.B2(n_340),
.C(n_297),
.Y(n_807)
);

AOI22xp33_ASAP7_75t_L g808 ( 
.A1(n_631),
.A2(n_614),
.B1(n_597),
.B2(n_594),
.Y(n_808)
);

OR2x2_ASAP7_75t_L g809 ( 
.A(n_644),
.B(n_507),
.Y(n_809)
);

NAND2xp5_ASAP7_75t_SL g810 ( 
.A(n_688),
.B(n_554),
.Y(n_810)
);

NAND2xp33_ASAP7_75t_L g811 ( 
.A(n_626),
.B(n_357),
.Y(n_811)
);

NAND2xp5_ASAP7_75t_L g812 ( 
.A(n_749),
.B(n_594),
.Y(n_812)
);

INVx1_ASAP7_75t_L g813 ( 
.A(n_740),
.Y(n_813)
);

AOI22xp5_ASAP7_75t_L g814 ( 
.A1(n_674),
.A2(n_522),
.B1(n_529),
.B2(n_505),
.Y(n_814)
);

NAND2xp5_ASAP7_75t_L g815 ( 
.A(n_714),
.B(n_597),
.Y(n_815)
);

INVx1_ASAP7_75t_L g816 ( 
.A(n_740),
.Y(n_816)
);

NOR2xp33_ASAP7_75t_L g817 ( 
.A(n_677),
.B(n_578),
.Y(n_817)
);

INVxp67_ASAP7_75t_L g818 ( 
.A(n_677),
.Y(n_818)
);

INVx1_ASAP7_75t_L g819 ( 
.A(n_744),
.Y(n_819)
);

INVx2_ASAP7_75t_L g820 ( 
.A(n_713),
.Y(n_820)
);

NAND2xp5_ASAP7_75t_L g821 ( 
.A(n_724),
.B(n_597),
.Y(n_821)
);

NAND2xp5_ASAP7_75t_SL g822 ( 
.A(n_688),
.B(n_554),
.Y(n_822)
);

BUFx3_ASAP7_75t_L g823 ( 
.A(n_682),
.Y(n_823)
);

INVx2_ASAP7_75t_L g824 ( 
.A(n_717),
.Y(n_824)
);

AOI22xp33_ASAP7_75t_L g825 ( 
.A1(n_631),
.A2(n_614),
.B1(n_597),
.B2(n_548),
.Y(n_825)
);

INVx2_ASAP7_75t_L g826 ( 
.A(n_717),
.Y(n_826)
);

AND2x2_ASAP7_75t_L g827 ( 
.A(n_620),
.B(n_633),
.Y(n_827)
);

NAND2xp5_ASAP7_75t_L g828 ( 
.A(n_652),
.B(n_720),
.Y(n_828)
);

NAND2xp5_ASAP7_75t_L g829 ( 
.A(n_652),
.B(n_597),
.Y(n_829)
);

NAND2xp5_ASAP7_75t_L g830 ( 
.A(n_652),
.B(n_614),
.Y(n_830)
);

OAI22xp5_ASAP7_75t_L g831 ( 
.A1(n_703),
.A2(n_256),
.B1(n_263),
.B2(n_259),
.Y(n_831)
);

INVx2_ASAP7_75t_L g832 ( 
.A(n_718),
.Y(n_832)
);

INVx1_ASAP7_75t_L g833 ( 
.A(n_744),
.Y(n_833)
);

NAND2xp5_ASAP7_75t_L g834 ( 
.A(n_652),
.B(n_614),
.Y(n_834)
);

AOI22xp33_ASAP7_75t_L g835 ( 
.A1(n_650),
.A2(n_614),
.B1(n_573),
.B2(n_557),
.Y(n_835)
);

INVx1_ASAP7_75t_L g836 ( 
.A(n_745),
.Y(n_836)
);

BUFx8_ASAP7_75t_L g837 ( 
.A(n_632),
.Y(n_837)
);

NAND2xp5_ASAP7_75t_SL g838 ( 
.A(n_662),
.B(n_606),
.Y(n_838)
);

NAND2xp5_ASAP7_75t_SL g839 ( 
.A(n_662),
.B(n_606),
.Y(n_839)
);

INVx1_ASAP7_75t_L g840 ( 
.A(n_745),
.Y(n_840)
);

INVxp67_ASAP7_75t_SL g841 ( 
.A(n_626),
.Y(n_841)
);

NAND2xp5_ASAP7_75t_L g842 ( 
.A(n_720),
.B(n_541),
.Y(n_842)
);

NOR2xp33_ASAP7_75t_L g843 ( 
.A(n_708),
.B(n_578),
.Y(n_843)
);

AOI221xp5_ASAP7_75t_L g844 ( 
.A1(n_711),
.A2(n_342),
.B1(n_301),
.B2(n_317),
.C(n_324),
.Y(n_844)
);

AOI22xp33_ASAP7_75t_L g845 ( 
.A1(n_650),
.A2(n_557),
.B1(n_573),
.B2(n_553),
.Y(n_845)
);

INVx2_ASAP7_75t_SL g846 ( 
.A(n_670),
.Y(n_846)
);

AND2x4_ASAP7_75t_L g847 ( 
.A(n_732),
.B(n_553),
.Y(n_847)
);

INVx2_ASAP7_75t_L g848 ( 
.A(n_718),
.Y(n_848)
);

NAND2xp5_ASAP7_75t_SL g849 ( 
.A(n_662),
.B(n_606),
.Y(n_849)
);

NAND2xp5_ASAP7_75t_L g850 ( 
.A(n_720),
.B(n_619),
.Y(n_850)
);

INVx3_ASAP7_75t_L g851 ( 
.A(n_619),
.Y(n_851)
);

INVx1_ASAP7_75t_L g852 ( 
.A(n_748),
.Y(n_852)
);

BUFx6f_ASAP7_75t_L g853 ( 
.A(n_723),
.Y(n_853)
);

AOI22xp33_ASAP7_75t_L g854 ( 
.A1(n_640),
.A2(n_557),
.B1(n_573),
.B2(n_553),
.Y(n_854)
);

NOR3xp33_ASAP7_75t_SL g855 ( 
.A(n_641),
.B(n_276),
.C(n_269),
.Y(n_855)
);

NAND2xp5_ASAP7_75t_SL g856 ( 
.A(n_720),
.B(n_557),
.Y(n_856)
);

INVx1_ASAP7_75t_L g857 ( 
.A(n_748),
.Y(n_857)
);

CKINVDCx5p33_ASAP7_75t_R g858 ( 
.A(n_712),
.Y(n_858)
);

NAND2xp5_ASAP7_75t_L g859 ( 
.A(n_621),
.B(n_624),
.Y(n_859)
);

OR2x6_ASAP7_75t_L g860 ( 
.A(n_761),
.B(n_587),
.Y(n_860)
);

NAND3xp33_ASAP7_75t_L g861 ( 
.A(n_633),
.B(n_587),
.C(n_281),
.Y(n_861)
);

NAND2xp5_ASAP7_75t_L g862 ( 
.A(n_621),
.B(n_587),
.Y(n_862)
);

NAND2xp5_ASAP7_75t_SL g863 ( 
.A(n_624),
.B(n_557),
.Y(n_863)
);

INVx1_ASAP7_75t_L g864 ( 
.A(n_751),
.Y(n_864)
);

INVx2_ASAP7_75t_L g865 ( 
.A(n_721),
.Y(n_865)
);

OAI22xp33_ASAP7_75t_L g866 ( 
.A1(n_632),
.A2(n_259),
.B1(n_267),
.B2(n_263),
.Y(n_866)
);

OR2x2_ASAP7_75t_L g867 ( 
.A(n_630),
.B(n_503),
.Y(n_867)
);

NAND2xp5_ASAP7_75t_L g868 ( 
.A(n_643),
.B(n_573),
.Y(n_868)
);

INVx1_ASAP7_75t_L g869 ( 
.A(n_755),
.Y(n_869)
);

INVx2_ASAP7_75t_L g870 ( 
.A(n_721),
.Y(n_870)
);

AOI22xp5_ASAP7_75t_L g871 ( 
.A1(n_670),
.A2(n_386),
.B1(n_296),
.B2(n_339),
.Y(n_871)
);

NAND2xp5_ASAP7_75t_L g872 ( 
.A(n_643),
.B(n_573),
.Y(n_872)
);

A2O1A1Ixp33_ASAP7_75t_L g873 ( 
.A1(n_627),
.A2(n_317),
.B(n_324),
.C(n_301),
.Y(n_873)
);

INVx1_ASAP7_75t_L g874 ( 
.A(n_755),
.Y(n_874)
);

NAND2xp5_ASAP7_75t_SL g875 ( 
.A(n_657),
.B(n_335),
.Y(n_875)
);

NAND2xp5_ASAP7_75t_SL g876 ( 
.A(n_657),
.B(n_341),
.Y(n_876)
);

NAND2xp5_ASAP7_75t_L g877 ( 
.A(n_682),
.B(n_585),
.Y(n_877)
);

NAND2xp5_ASAP7_75t_L g878 ( 
.A(n_627),
.B(n_585),
.Y(n_878)
);

NOR2xp33_ASAP7_75t_L g879 ( 
.A(n_647),
.B(n_565),
.Y(n_879)
);

INVx4_ASAP7_75t_L g880 ( 
.A(n_723),
.Y(n_880)
);

BUFx3_ASAP7_75t_L g881 ( 
.A(n_759),
.Y(n_881)
);

INVx1_ASAP7_75t_L g882 ( 
.A(n_759),
.Y(n_882)
);

INVx2_ASAP7_75t_L g883 ( 
.A(n_693),
.Y(n_883)
);

NAND2xp5_ASAP7_75t_SL g884 ( 
.A(n_634),
.B(n_344),
.Y(n_884)
);

NAND2xp5_ASAP7_75t_L g885 ( 
.A(n_634),
.B(n_585),
.Y(n_885)
);

INVx2_ASAP7_75t_L g886 ( 
.A(n_693),
.Y(n_886)
);

NOR2xp33_ASAP7_75t_L g887 ( 
.A(n_648),
.B(n_565),
.Y(n_887)
);

INVx1_ASAP7_75t_L g888 ( 
.A(n_767),
.Y(n_888)
);

NOR2xp33_ASAP7_75t_L g889 ( 
.A(n_669),
.B(n_277),
.Y(n_889)
);

INVx1_ASAP7_75t_L g890 ( 
.A(n_767),
.Y(n_890)
);

NAND2xp5_ASAP7_75t_L g891 ( 
.A(n_635),
.B(n_585),
.Y(n_891)
);

NAND2xp5_ASAP7_75t_L g892 ( 
.A(n_635),
.B(n_585),
.Y(n_892)
);

NAND2xp5_ASAP7_75t_L g893 ( 
.A(n_637),
.B(n_589),
.Y(n_893)
);

NAND2xp5_ASAP7_75t_L g894 ( 
.A(n_637),
.B(n_589),
.Y(n_894)
);

INVx1_ASAP7_75t_L g895 ( 
.A(n_769),
.Y(n_895)
);

BUFx2_ASAP7_75t_L g896 ( 
.A(n_727),
.Y(n_896)
);

CKINVDCx5p33_ASAP7_75t_R g897 ( 
.A(n_771),
.Y(n_897)
);

A2O1A1Ixp33_ASAP7_75t_L g898 ( 
.A1(n_646),
.A2(n_392),
.B(n_327),
.C(n_331),
.Y(n_898)
);

AOI22xp5_ASAP7_75t_L g899 ( 
.A1(n_680),
.A2(n_393),
.B1(n_381),
.B2(n_385),
.Y(n_899)
);

INVx1_ASAP7_75t_L g900 ( 
.A(n_769),
.Y(n_900)
);

NAND2xp5_ASAP7_75t_L g901 ( 
.A(n_646),
.B(n_589),
.Y(n_901)
);

NAND2xp5_ASAP7_75t_SL g902 ( 
.A(n_655),
.B(n_347),
.Y(n_902)
);

INVx1_ASAP7_75t_L g903 ( 
.A(n_697),
.Y(n_903)
);

NAND3xp33_ASAP7_75t_L g904 ( 
.A(n_645),
.B(n_286),
.C(n_283),
.Y(n_904)
);

INVx2_ASAP7_75t_L g905 ( 
.A(n_697),
.Y(n_905)
);

NAND2xp5_ASAP7_75t_L g906 ( 
.A(n_655),
.B(n_589),
.Y(n_906)
);

NAND2xp5_ASAP7_75t_SL g907 ( 
.A(n_656),
.B(n_350),
.Y(n_907)
);

INVx2_ASAP7_75t_SL g908 ( 
.A(n_732),
.Y(n_908)
);

AND2x2_ASAP7_75t_L g909 ( 
.A(n_645),
.B(n_581),
.Y(n_909)
);

INVx1_ASAP7_75t_L g910 ( 
.A(n_699),
.Y(n_910)
);

OR2x2_ASAP7_75t_SL g911 ( 
.A(n_639),
.B(n_327),
.Y(n_911)
);

AOI22xp5_ASAP7_75t_L g912 ( 
.A1(n_705),
.A2(n_389),
.B1(n_355),
.B2(n_360),
.Y(n_912)
);

NAND2xp5_ASAP7_75t_SL g913 ( 
.A(n_656),
.B(n_353),
.Y(n_913)
);

NAND2xp5_ASAP7_75t_L g914 ( 
.A(n_660),
.B(n_589),
.Y(n_914)
);

NOR2x1p5_ASAP7_75t_L g915 ( 
.A(n_771),
.B(n_287),
.Y(n_915)
);

INVx1_ASAP7_75t_L g916 ( 
.A(n_699),
.Y(n_916)
);

AOI22xp33_ASAP7_75t_L g917 ( 
.A1(n_660),
.A2(n_338),
.B1(n_356),
.B2(n_337),
.Y(n_917)
);

NOR2xp33_ASAP7_75t_L g918 ( 
.A(n_763),
.B(n_300),
.Y(n_918)
);

NAND2xp5_ASAP7_75t_SL g919 ( 
.A(n_664),
.B(n_365),
.Y(n_919)
);

INVx1_ASAP7_75t_L g920 ( 
.A(n_701),
.Y(n_920)
);

NAND2xp5_ASAP7_75t_L g921 ( 
.A(n_664),
.B(n_580),
.Y(n_921)
);

NAND2xp5_ASAP7_75t_L g922 ( 
.A(n_701),
.B(n_580),
.Y(n_922)
);

AOI22xp5_ASAP7_75t_L g923 ( 
.A1(n_722),
.A2(n_366),
.B1(n_417),
.B2(n_410),
.Y(n_923)
);

INVx2_ASAP7_75t_L g924 ( 
.A(n_704),
.Y(n_924)
);

BUFx6f_ASAP7_75t_SL g925 ( 
.A(n_761),
.Y(n_925)
);

NOR2xp33_ASAP7_75t_L g926 ( 
.A(n_725),
.B(n_303),
.Y(n_926)
);

AOI22xp33_ASAP7_75t_L g927 ( 
.A1(n_747),
.A2(n_337),
.B1(n_356),
.B2(n_338),
.Y(n_927)
);

NAND2x1_ASAP7_75t_L g928 ( 
.A(n_710),
.B(n_555),
.Y(n_928)
);

NAND2xp33_ASAP7_75t_L g929 ( 
.A(n_684),
.B(n_555),
.Y(n_929)
);

NAND2xp5_ASAP7_75t_SL g930 ( 
.A(n_723),
.B(n_369),
.Y(n_930)
);

NOR2xp33_ASAP7_75t_L g931 ( 
.A(n_704),
.B(n_305),
.Y(n_931)
);

INVxp67_ASAP7_75t_L g932 ( 
.A(n_764),
.Y(n_932)
);

INVx1_ASAP7_75t_L g933 ( 
.A(n_716),
.Y(n_933)
);

NAND2xp5_ASAP7_75t_L g934 ( 
.A(n_716),
.B(n_580),
.Y(n_934)
);

NAND2xp5_ASAP7_75t_L g935 ( 
.A(n_726),
.B(n_580),
.Y(n_935)
);

INVx1_ASAP7_75t_L g936 ( 
.A(n_726),
.Y(n_936)
);

NAND2xp5_ASAP7_75t_SL g937 ( 
.A(n_709),
.B(n_377),
.Y(n_937)
);

NAND2xp5_ASAP7_75t_SL g938 ( 
.A(n_686),
.B(n_379),
.Y(n_938)
);

NAND2xp5_ASAP7_75t_L g939 ( 
.A(n_728),
.B(n_580),
.Y(n_939)
);

NAND2xp5_ASAP7_75t_L g940 ( 
.A(n_728),
.B(n_593),
.Y(n_940)
);

NAND2xp5_ASAP7_75t_L g941 ( 
.A(n_730),
.B(n_593),
.Y(n_941)
);

NAND2xp5_ASAP7_75t_L g942 ( 
.A(n_730),
.B(n_593),
.Y(n_942)
);

AOI21xp5_ASAP7_75t_L g943 ( 
.A1(n_856),
.A2(n_736),
.B(n_741),
.Y(n_943)
);

NAND2xp5_ASAP7_75t_L g944 ( 
.A(n_780),
.B(n_783),
.Y(n_944)
);

NAND2xp5_ASAP7_75t_L g945 ( 
.A(n_785),
.B(n_733),
.Y(n_945)
);

BUFx3_ASAP7_75t_L g946 ( 
.A(n_837),
.Y(n_946)
);

AND2x2_ASAP7_75t_L g947 ( 
.A(n_827),
.B(n_761),
.Y(n_947)
);

NAND2xp5_ASAP7_75t_L g948 ( 
.A(n_787),
.B(n_733),
.Y(n_948)
);

O2A1O1Ixp5_ASAP7_75t_L g949 ( 
.A1(n_884),
.A2(n_735),
.B(n_738),
.C(n_734),
.Y(n_949)
);

AOI21xp5_ASAP7_75t_L g950 ( 
.A1(n_856),
.A2(n_741),
.B(n_715),
.Y(n_950)
);

AOI21xp5_ASAP7_75t_L g951 ( 
.A1(n_829),
.A2(n_741),
.B(n_715),
.Y(n_951)
);

NAND2xp5_ASAP7_75t_L g952 ( 
.A(n_773),
.B(n_734),
.Y(n_952)
);

BUFx3_ASAP7_75t_L g953 ( 
.A(n_774),
.Y(n_953)
);

AOI21xp5_ASAP7_75t_L g954 ( 
.A1(n_792),
.A2(n_741),
.B(n_715),
.Y(n_954)
);

NAND2xp33_ASAP7_75t_L g955 ( 
.A(n_796),
.B(n_710),
.Y(n_955)
);

AOI21xp5_ASAP7_75t_L g956 ( 
.A1(n_795),
.A2(n_741),
.B(n_715),
.Y(n_956)
);

INVxp67_ASAP7_75t_L g957 ( 
.A(n_790),
.Y(n_957)
);

AOI21xp5_ASAP7_75t_L g958 ( 
.A1(n_830),
.A2(n_715),
.B(n_676),
.Y(n_958)
);

AOI21xp5_ASAP7_75t_L g959 ( 
.A1(n_834),
.A2(n_676),
.B(n_673),
.Y(n_959)
);

OAI22xp5_ASAP7_75t_L g960 ( 
.A1(n_841),
.A2(n_756),
.B1(n_695),
.B2(n_729),
.Y(n_960)
);

INVx1_ASAP7_75t_L g961 ( 
.A(n_881),
.Y(n_961)
);

INVx3_ASAP7_75t_L g962 ( 
.A(n_881),
.Y(n_962)
);

NAND2xp5_ASAP7_75t_L g963 ( 
.A(n_793),
.B(n_735),
.Y(n_963)
);

INVx2_ASAP7_75t_L g964 ( 
.A(n_851),
.Y(n_964)
);

NAND2xp5_ASAP7_75t_L g965 ( 
.A(n_800),
.B(n_738),
.Y(n_965)
);

NOR2xp33_ASAP7_75t_R g966 ( 
.A(n_802),
.B(n_695),
.Y(n_966)
);

NOR2xp33_ASAP7_75t_L g967 ( 
.A(n_818),
.B(n_706),
.Y(n_967)
);

INVx4_ASAP7_75t_L g968 ( 
.A(n_774),
.Y(n_968)
);

AOI21xp5_ASAP7_75t_L g969 ( 
.A1(n_842),
.A2(n_676),
.B(n_673),
.Y(n_969)
);

NAND2xp5_ASAP7_75t_L g970 ( 
.A(n_909),
.B(n_706),
.Y(n_970)
);

AOI21xp5_ASAP7_75t_L g971 ( 
.A1(n_850),
.A2(n_681),
.B(n_673),
.Y(n_971)
);

NAND2xp33_ASAP7_75t_L g972 ( 
.A(n_796),
.B(n_710),
.Y(n_972)
);

OAI21xp5_ASAP7_75t_L g973 ( 
.A1(n_884),
.A2(n_729),
.B(n_651),
.Y(n_973)
);

A2O1A1Ixp33_ASAP7_75t_L g974 ( 
.A1(n_781),
.A2(n_413),
.B(n_372),
.C(n_406),
.Y(n_974)
);

INVx2_ASAP7_75t_L g975 ( 
.A(n_883),
.Y(n_975)
);

AOI21xp5_ASAP7_75t_L g976 ( 
.A1(n_828),
.A2(n_700),
.B(n_681),
.Y(n_976)
);

INVx2_ASAP7_75t_L g977 ( 
.A(n_883),
.Y(n_977)
);

NOR2xp67_ASAP7_75t_L g978 ( 
.A(n_814),
.B(n_584),
.Y(n_978)
);

NAND2xp5_ASAP7_75t_L g979 ( 
.A(n_789),
.B(n_784),
.Y(n_979)
);

AND2x2_ASAP7_75t_SL g980 ( 
.A(n_788),
.B(n_267),
.Y(n_980)
);

HB1xp67_ASAP7_75t_L g981 ( 
.A(n_791),
.Y(n_981)
);

INVx4_ASAP7_75t_L g982 ( 
.A(n_774),
.Y(n_982)
);

INVx2_ASAP7_75t_SL g983 ( 
.A(n_867),
.Y(n_983)
);

NOR2xp33_ASAP7_75t_L g984 ( 
.A(n_896),
.B(n_761),
.Y(n_984)
);

INVx1_ASAP7_75t_L g985 ( 
.A(n_813),
.Y(n_985)
);

NAND2xp5_ASAP7_75t_L g986 ( 
.A(n_903),
.B(n_761),
.Y(n_986)
);

INVx3_ASAP7_75t_L g987 ( 
.A(n_823),
.Y(n_987)
);

INVx3_ASAP7_75t_L g988 ( 
.A(n_823),
.Y(n_988)
);

NOR2xp33_ASAP7_75t_L g989 ( 
.A(n_798),
.B(n_306),
.Y(n_989)
);

AOI21xp5_ASAP7_75t_L g990 ( 
.A1(n_786),
.A2(n_700),
.B(n_681),
.Y(n_990)
);

INVxp67_ASAP7_75t_L g991 ( 
.A(n_809),
.Y(n_991)
);

NAND2xp5_ASAP7_75t_L g992 ( 
.A(n_910),
.B(n_916),
.Y(n_992)
);

INVx11_ASAP7_75t_L g993 ( 
.A(n_837),
.Y(n_993)
);

AOI21xp5_ASAP7_75t_L g994 ( 
.A1(n_786),
.A2(n_754),
.B(n_700),
.Y(n_994)
);

O2A1O1Ixp33_ASAP7_75t_L g995 ( 
.A1(n_873),
.A2(n_898),
.B(n_831),
.C(n_799),
.Y(n_995)
);

AOI21xp5_ASAP7_75t_L g996 ( 
.A1(n_810),
.A2(n_822),
.B(n_821),
.Y(n_996)
);

AOI21xp5_ASAP7_75t_L g997 ( 
.A1(n_810),
.A2(n_754),
.B(n_698),
.Y(n_997)
);

AOI22xp33_ASAP7_75t_L g998 ( 
.A1(n_776),
.A2(n_349),
.B1(n_362),
.B2(n_358),
.Y(n_998)
);

A2O1A1Ixp33_ASAP7_75t_L g999 ( 
.A1(n_844),
.A2(n_413),
.B(n_372),
.C(n_406),
.Y(n_999)
);

AO21x1_ASAP7_75t_L g1000 ( 
.A1(n_902),
.A2(n_294),
.B(n_271),
.Y(n_1000)
);

BUFx4f_ASAP7_75t_L g1001 ( 
.A(n_774),
.Y(n_1001)
);

BUFx6f_ASAP7_75t_L g1002 ( 
.A(n_796),
.Y(n_1002)
);

NAND2xp5_ASAP7_75t_L g1003 ( 
.A(n_920),
.B(n_628),
.Y(n_1003)
);

BUFx8_ASAP7_75t_L g1004 ( 
.A(n_925),
.Y(n_1004)
);

INVx1_ASAP7_75t_SL g1005 ( 
.A(n_911),
.Y(n_1005)
);

NAND2xp5_ASAP7_75t_L g1006 ( 
.A(n_933),
.B(n_628),
.Y(n_1006)
);

A2O1A1Ixp33_ASAP7_75t_L g1007 ( 
.A1(n_926),
.A2(n_889),
.B(n_898),
.C(n_873),
.Y(n_1007)
);

INVx2_ASAP7_75t_SL g1008 ( 
.A(n_846),
.Y(n_1008)
);

NAND2xp5_ASAP7_75t_L g1009 ( 
.A(n_936),
.B(n_628),
.Y(n_1009)
);

AND2x2_ASAP7_75t_SL g1010 ( 
.A(n_811),
.B(n_271),
.Y(n_1010)
);

CKINVDCx5p33_ASAP7_75t_R g1011 ( 
.A(n_802),
.Y(n_1011)
);

INVx1_ASAP7_75t_L g1012 ( 
.A(n_816),
.Y(n_1012)
);

INVx2_ASAP7_75t_L g1013 ( 
.A(n_886),
.Y(n_1013)
);

AO21x1_ASAP7_75t_L g1014 ( 
.A1(n_902),
.A2(n_295),
.B(n_294),
.Y(n_1014)
);

NAND2xp5_ASAP7_75t_L g1015 ( 
.A(n_886),
.B(n_628),
.Y(n_1015)
);

NAND2xp5_ASAP7_75t_L g1016 ( 
.A(n_905),
.B(n_651),
.Y(n_1016)
);

AOI21xp5_ASAP7_75t_L g1017 ( 
.A1(n_822),
.A2(n_815),
.B(n_811),
.Y(n_1017)
);

INVx1_ASAP7_75t_L g1018 ( 
.A(n_819),
.Y(n_1018)
);

NOR3xp33_ASAP7_75t_L g1019 ( 
.A(n_817),
.B(n_591),
.C(n_584),
.Y(n_1019)
);

NAND2xp5_ASAP7_75t_L g1020 ( 
.A(n_905),
.B(n_651),
.Y(n_1020)
);

INVx2_ASAP7_75t_L g1021 ( 
.A(n_924),
.Y(n_1021)
);

AOI21xp5_ASAP7_75t_L g1022 ( 
.A1(n_859),
.A2(n_754),
.B(n_698),
.Y(n_1022)
);

AOI22xp5_ASAP7_75t_L g1023 ( 
.A1(n_804),
.A2(n_752),
.B1(n_766),
.B2(n_742),
.Y(n_1023)
);

NOR2xp33_ASAP7_75t_L g1024 ( 
.A(n_932),
.B(n_308),
.Y(n_1024)
);

INVxp67_ASAP7_75t_L g1025 ( 
.A(n_918),
.Y(n_1025)
);

O2A1O1Ixp33_ASAP7_75t_L g1026 ( 
.A1(n_801),
.A2(n_368),
.B(n_395),
.C(n_312),
.Y(n_1026)
);

NAND2xp5_ASAP7_75t_L g1027 ( 
.A(n_924),
.B(n_651),
.Y(n_1027)
);

NAND2xp5_ASAP7_75t_SL g1028 ( 
.A(n_796),
.B(n_686),
.Y(n_1028)
);

AND2x2_ASAP7_75t_L g1029 ( 
.A(n_779),
.B(n_591),
.Y(n_1029)
);

AOI21xp5_ASAP7_75t_L g1030 ( 
.A1(n_812),
.A2(n_698),
.B(n_686),
.Y(n_1030)
);

AND2x2_ASAP7_75t_SL g1031 ( 
.A(n_880),
.B(n_295),
.Y(n_1031)
);

INVx1_ASAP7_75t_L g1032 ( 
.A(n_833),
.Y(n_1032)
);

OAI22xp5_ASAP7_75t_L g1033 ( 
.A1(n_775),
.A2(n_304),
.B1(n_312),
.B2(n_318),
.Y(n_1033)
);

OAI21xp33_ASAP7_75t_L g1034 ( 
.A1(n_931),
.A2(n_322),
.B(n_314),
.Y(n_1034)
);

NAND2xp5_ASAP7_75t_L g1035 ( 
.A(n_836),
.B(n_654),
.Y(n_1035)
);

NAND2xp5_ASAP7_75t_L g1036 ( 
.A(n_840),
.B(n_654),
.Y(n_1036)
);

BUFx6f_ASAP7_75t_L g1037 ( 
.A(n_853),
.Y(n_1037)
);

AOI21xp5_ASAP7_75t_L g1038 ( 
.A1(n_862),
.A2(n_698),
.B(n_686),
.Y(n_1038)
);

NAND2xp5_ASAP7_75t_SL g1039 ( 
.A(n_853),
.B(n_686),
.Y(n_1039)
);

BUFx12f_ASAP7_75t_L g1040 ( 
.A(n_837),
.Y(n_1040)
);

BUFx3_ASAP7_75t_L g1041 ( 
.A(n_847),
.Y(n_1041)
);

INVx1_ASAP7_75t_SL g1042 ( 
.A(n_858),
.Y(n_1042)
);

INVxp67_ASAP7_75t_L g1043 ( 
.A(n_904),
.Y(n_1043)
);

NAND2xp5_ASAP7_75t_L g1044 ( 
.A(n_852),
.B(n_654),
.Y(n_1044)
);

BUFx4f_ASAP7_75t_L g1045 ( 
.A(n_847),
.Y(n_1045)
);

NOR2xp33_ASAP7_75t_R g1046 ( 
.A(n_858),
.B(n_396),
.Y(n_1046)
);

O2A1O1Ixp33_ASAP7_75t_SL g1047 ( 
.A1(n_907),
.A2(n_395),
.B(n_321),
.C(n_318),
.Y(n_1047)
);

NAND2xp5_ASAP7_75t_SL g1048 ( 
.A(n_853),
.B(n_877),
.Y(n_1048)
);

AOI21x1_ASAP7_75t_L g1049 ( 
.A1(n_838),
.A2(n_667),
.B(n_666),
.Y(n_1049)
);

INVx3_ASAP7_75t_L g1050 ( 
.A(n_772),
.Y(n_1050)
);

AOI21xp5_ASAP7_75t_L g1051 ( 
.A1(n_868),
.A2(n_698),
.B(n_686),
.Y(n_1051)
);

AOI21xp5_ASAP7_75t_L g1052 ( 
.A1(n_872),
.A2(n_698),
.B(n_629),
.Y(n_1052)
);

AOI21xp5_ASAP7_75t_L g1053 ( 
.A1(n_808),
.A2(n_707),
.B(n_629),
.Y(n_1053)
);

NOR2xp67_ASAP7_75t_L g1054 ( 
.A(n_861),
.B(n_595),
.Y(n_1054)
);

NOR2xp67_ASAP7_75t_L g1055 ( 
.A(n_912),
.B(n_595),
.Y(n_1055)
);

INVxp67_ASAP7_75t_SL g1056 ( 
.A(n_853),
.Y(n_1056)
);

AND2x2_ASAP7_75t_L g1057 ( 
.A(n_879),
.B(n_887),
.Y(n_1057)
);

NOR2xp33_ASAP7_75t_L g1058 ( 
.A(n_794),
.B(n_326),
.Y(n_1058)
);

NAND2xp5_ASAP7_75t_L g1059 ( 
.A(n_857),
.B(n_654),
.Y(n_1059)
);

AOI21x1_ASAP7_75t_L g1060 ( 
.A1(n_838),
.A2(n_667),
.B(n_666),
.Y(n_1060)
);

NAND2xp5_ASAP7_75t_L g1061 ( 
.A(n_864),
.B(n_691),
.Y(n_1061)
);

NAND2xp5_ASAP7_75t_L g1062 ( 
.A(n_869),
.B(n_874),
.Y(n_1062)
);

AOI21xp5_ASAP7_75t_L g1063 ( 
.A1(n_839),
.A2(n_707),
.B(n_629),
.Y(n_1063)
);

AOI21xp5_ASAP7_75t_L g1064 ( 
.A1(n_839),
.A2(n_707),
.B(n_629),
.Y(n_1064)
);

O2A1O1Ixp33_ASAP7_75t_L g1065 ( 
.A1(n_866),
.A2(n_336),
.B(n_368),
.C(n_375),
.Y(n_1065)
);

NAND2xp5_ASAP7_75t_L g1066 ( 
.A(n_882),
.B(n_691),
.Y(n_1066)
);

INVx1_ASAP7_75t_L g1067 ( 
.A(n_888),
.Y(n_1067)
);

AOI21xp5_ASAP7_75t_L g1068 ( 
.A1(n_849),
.A2(n_707),
.B(n_629),
.Y(n_1068)
);

NOR2xp33_ASAP7_75t_L g1069 ( 
.A(n_843),
.B(n_332),
.Y(n_1069)
);

AOI21xp5_ASAP7_75t_L g1070 ( 
.A1(n_849),
.A2(n_750),
.B(n_707),
.Y(n_1070)
);

AOI33xp33_ASAP7_75t_L g1071 ( 
.A1(n_908),
.A2(n_521),
.A3(n_527),
.B1(n_349),
.B2(n_404),
.B3(n_392),
.Y(n_1071)
);

NOR2xp33_ASAP7_75t_L g1072 ( 
.A(n_847),
.B(n_334),
.Y(n_1072)
);

AOI21xp5_ASAP7_75t_L g1073 ( 
.A1(n_825),
.A2(n_750),
.B(n_719),
.Y(n_1073)
);

O2A1O1Ixp33_ASAP7_75t_L g1074 ( 
.A1(n_907),
.A2(n_304),
.B(n_321),
.C(n_336),
.Y(n_1074)
);

INVx2_ASAP7_75t_L g1075 ( 
.A(n_772),
.Y(n_1075)
);

BUFx6f_ASAP7_75t_L g1076 ( 
.A(n_860),
.Y(n_1076)
);

AOI21xp5_ASAP7_75t_L g1077 ( 
.A1(n_863),
.A2(n_750),
.B(n_719),
.Y(n_1077)
);

NAND2xp5_ASAP7_75t_L g1078 ( 
.A(n_890),
.B(n_691),
.Y(n_1078)
);

NAND2xp5_ASAP7_75t_L g1079 ( 
.A(n_895),
.B(n_691),
.Y(n_1079)
);

NOR2xp33_ASAP7_75t_R g1080 ( 
.A(n_897),
.B(n_398),
.Y(n_1080)
);

NAND2xp5_ASAP7_75t_L g1081 ( 
.A(n_900),
.B(n_719),
.Y(n_1081)
);

NAND2xp5_ASAP7_75t_L g1082 ( 
.A(n_803),
.B(n_719),
.Y(n_1082)
);

INVx1_ASAP7_75t_L g1083 ( 
.A(n_778),
.Y(n_1083)
);

BUFx6f_ASAP7_75t_L g1084 ( 
.A(n_860),
.Y(n_1084)
);

INVx2_ASAP7_75t_L g1085 ( 
.A(n_778),
.Y(n_1085)
);

INVx1_ASAP7_75t_L g1086 ( 
.A(n_782),
.Y(n_1086)
);

AOI21xp5_ASAP7_75t_L g1087 ( 
.A1(n_863),
.A2(n_750),
.B(n_731),
.Y(n_1087)
);

NAND2xp5_ASAP7_75t_L g1088 ( 
.A(n_805),
.B(n_731),
.Y(n_1088)
);

INVx3_ASAP7_75t_L g1089 ( 
.A(n_820),
.Y(n_1089)
);

NAND2xp5_ASAP7_75t_L g1090 ( 
.A(n_806),
.B(n_731),
.Y(n_1090)
);

OAI21xp5_ASAP7_75t_L g1091 ( 
.A1(n_913),
.A2(n_753),
.B(n_742),
.Y(n_1091)
);

NOR2xp33_ASAP7_75t_L g1092 ( 
.A(n_871),
.B(n_345),
.Y(n_1092)
);

NOR2xp33_ASAP7_75t_L g1093 ( 
.A(n_777),
.B(n_875),
.Y(n_1093)
);

O2A1O1Ixp33_ASAP7_75t_L g1094 ( 
.A1(n_913),
.A2(n_380),
.B(n_375),
.C(n_613),
.Y(n_1094)
);

NOR2xp33_ASAP7_75t_L g1095 ( 
.A(n_875),
.B(n_351),
.Y(n_1095)
);

OAI22xp33_ASAP7_75t_L g1096 ( 
.A1(n_860),
.A2(n_380),
.B1(n_331),
.B2(n_340),
.Y(n_1096)
);

A2O1A1Ixp33_ASAP7_75t_L g1097 ( 
.A1(n_878),
.A2(n_343),
.B(n_348),
.C(n_352),
.Y(n_1097)
);

BUFx8_ASAP7_75t_SL g1098 ( 
.A(n_897),
.Y(n_1098)
);

AND2x2_ASAP7_75t_L g1099 ( 
.A(n_797),
.B(n_599),
.Y(n_1099)
);

BUFx2_ASAP7_75t_L g1100 ( 
.A(n_860),
.Y(n_1100)
);

A2O1A1Ixp33_ASAP7_75t_L g1101 ( 
.A1(n_885),
.A2(n_343),
.B(n_348),
.C(n_352),
.Y(n_1101)
);

INVx1_ASAP7_75t_L g1102 ( 
.A(n_820),
.Y(n_1102)
);

AOI21xp5_ASAP7_75t_L g1103 ( 
.A1(n_891),
.A2(n_750),
.B(n_753),
.Y(n_1103)
);

AOI21xp5_ASAP7_75t_L g1104 ( 
.A1(n_892),
.A2(n_753),
.B(n_671),
.Y(n_1104)
);

A2O1A1Ixp33_ASAP7_75t_L g1105 ( 
.A1(n_893),
.A2(n_358),
.B(n_362),
.C(n_390),
.Y(n_1105)
);

AOI21xp5_ASAP7_75t_L g1106 ( 
.A1(n_894),
.A2(n_906),
.B(n_901),
.Y(n_1106)
);

CKINVDCx8_ASAP7_75t_R g1107 ( 
.A(n_776),
.Y(n_1107)
);

AOI22xp5_ASAP7_75t_L g1108 ( 
.A1(n_876),
.A2(n_766),
.B1(n_710),
.B2(n_742),
.Y(n_1108)
);

NAND2xp5_ASAP7_75t_L g1109 ( 
.A(n_917),
.B(n_753),
.Y(n_1109)
);

NAND2xp5_ASAP7_75t_SL g1110 ( 
.A(n_880),
.B(n_668),
.Y(n_1110)
);

AOI21xp5_ASAP7_75t_L g1111 ( 
.A1(n_914),
.A2(n_671),
.B(n_668),
.Y(n_1111)
);

AOI21x1_ASAP7_75t_L g1112 ( 
.A1(n_919),
.A2(n_678),
.B(n_672),
.Y(n_1112)
);

O2A1O1Ixp33_ASAP7_75t_L g1113 ( 
.A1(n_919),
.A2(n_600),
.B(n_599),
.C(n_611),
.Y(n_1113)
);

O2A1O1Ixp33_ASAP7_75t_L g1114 ( 
.A1(n_937),
.A2(n_600),
.B(n_611),
.C(n_613),
.Y(n_1114)
);

INVx2_ASAP7_75t_SL g1115 ( 
.A(n_915),
.Y(n_1115)
);

NAND2xp5_ASAP7_75t_SL g1116 ( 
.A(n_880),
.B(n_672),
.Y(n_1116)
);

NAND2xp5_ASAP7_75t_L g1117 ( 
.A(n_854),
.B(n_678),
.Y(n_1117)
);

BUFx2_ASAP7_75t_L g1118 ( 
.A(n_855),
.Y(n_1118)
);

INVx1_ASAP7_75t_L g1119 ( 
.A(n_824),
.Y(n_1119)
);

AOI21xp5_ASAP7_75t_L g1120 ( 
.A1(n_921),
.A2(n_687),
.B(n_679),
.Y(n_1120)
);

NAND2xp5_ASAP7_75t_SL g1121 ( 
.A(n_824),
.B(n_679),
.Y(n_1121)
);

NAND2xp5_ASAP7_75t_L g1122 ( 
.A(n_826),
.B(n_683),
.Y(n_1122)
);

O2A1O1Ixp33_ASAP7_75t_L g1123 ( 
.A1(n_937),
.A2(n_618),
.B(n_617),
.C(n_615),
.Y(n_1123)
);

NAND2xp5_ASAP7_75t_L g1124 ( 
.A(n_826),
.B(n_683),
.Y(n_1124)
);

NOR2xp33_ASAP7_75t_L g1125 ( 
.A(n_876),
.B(n_354),
.Y(n_1125)
);

AOI21xp5_ASAP7_75t_L g1126 ( 
.A1(n_929),
.A2(n_689),
.B(n_690),
.Y(n_1126)
);

INVx1_ASAP7_75t_L g1127 ( 
.A(n_832),
.Y(n_1127)
);

AOI21xp5_ASAP7_75t_L g1128 ( 
.A1(n_929),
.A2(n_689),
.B(n_690),
.Y(n_1128)
);

NAND2xp5_ASAP7_75t_L g1129 ( 
.A(n_832),
.B(n_687),
.Y(n_1129)
);

AOI21xp5_ASAP7_75t_L g1130 ( 
.A1(n_930),
.A2(n_692),
.B(n_757),
.Y(n_1130)
);

INVx1_ASAP7_75t_L g1131 ( 
.A(n_848),
.Y(n_1131)
);

NAND2xp5_ASAP7_75t_SL g1132 ( 
.A(n_980),
.B(n_848),
.Y(n_1132)
);

O2A1O1Ixp33_ASAP7_75t_L g1133 ( 
.A1(n_989),
.A2(n_930),
.B(n_922),
.C(n_934),
.Y(n_1133)
);

AOI21xp5_ASAP7_75t_L g1134 ( 
.A1(n_943),
.A2(n_938),
.B(n_845),
.Y(n_1134)
);

A2O1A1Ixp33_ASAP7_75t_L g1135 ( 
.A1(n_989),
.A2(n_899),
.B(n_835),
.C(n_939),
.Y(n_1135)
);

INVx3_ASAP7_75t_L g1136 ( 
.A(n_1002),
.Y(n_1136)
);

BUFx12f_ASAP7_75t_L g1137 ( 
.A(n_1040),
.Y(n_1137)
);

INVx1_ASAP7_75t_L g1138 ( 
.A(n_975),
.Y(n_1138)
);

BUFx8_ASAP7_75t_L g1139 ( 
.A(n_946),
.Y(n_1139)
);

AND2x4_ASAP7_75t_L g1140 ( 
.A(n_1041),
.B(n_865),
.Y(n_1140)
);

NAND2xp5_ASAP7_75t_L g1141 ( 
.A(n_944),
.B(n_776),
.Y(n_1141)
);

NAND3xp33_ASAP7_75t_SL g1142 ( 
.A(n_1069),
.B(n_923),
.C(n_477),
.Y(n_1142)
);

NAND2xp5_ASAP7_75t_L g1143 ( 
.A(n_1057),
.B(n_776),
.Y(n_1143)
);

NOR2xp33_ASAP7_75t_L g1144 ( 
.A(n_980),
.B(n_865),
.Y(n_1144)
);

NOR2xp33_ASAP7_75t_L g1145 ( 
.A(n_1025),
.B(n_870),
.Y(n_1145)
);

INVx1_ASAP7_75t_L g1146 ( 
.A(n_977),
.Y(n_1146)
);

NOR2xp33_ASAP7_75t_L g1147 ( 
.A(n_991),
.B(n_870),
.Y(n_1147)
);

OR2x6_ASAP7_75t_L g1148 ( 
.A(n_1076),
.B(n_928),
.Y(n_1148)
);

NAND2xp5_ASAP7_75t_L g1149 ( 
.A(n_979),
.B(n_776),
.Y(n_1149)
);

NAND2xp5_ASAP7_75t_SL g1150 ( 
.A(n_987),
.B(n_935),
.Y(n_1150)
);

INVx1_ASAP7_75t_L g1151 ( 
.A(n_1013),
.Y(n_1151)
);

NAND2xp5_ASAP7_75t_SL g1152 ( 
.A(n_962),
.B(n_940),
.Y(n_1152)
);

OAI21xp5_ASAP7_75t_L g1153 ( 
.A1(n_1007),
.A2(n_942),
.B(n_941),
.Y(n_1153)
);

HB1xp67_ASAP7_75t_L g1154 ( 
.A(n_981),
.Y(n_1154)
);

AOI21xp5_ASAP7_75t_L g1155 ( 
.A1(n_1017),
.A2(n_938),
.B(n_927),
.Y(n_1155)
);

INVx2_ASAP7_75t_L g1156 ( 
.A(n_1050),
.Y(n_1156)
);

INVx3_ASAP7_75t_L g1157 ( 
.A(n_1002),
.Y(n_1157)
);

AOI21xp5_ASAP7_75t_L g1158 ( 
.A1(n_950),
.A2(n_692),
.B(n_739),
.Y(n_1158)
);

INVx2_ASAP7_75t_L g1159 ( 
.A(n_1089),
.Y(n_1159)
);

INVx6_ASAP7_75t_L g1160 ( 
.A(n_968),
.Y(n_1160)
);

A2O1A1Ixp33_ASAP7_75t_L g1161 ( 
.A1(n_1069),
.A2(n_404),
.B(n_391),
.C(n_390),
.Y(n_1161)
);

NOR2xp33_ASAP7_75t_L g1162 ( 
.A(n_1005),
.B(n_925),
.Y(n_1162)
);

NOR2xp33_ASAP7_75t_L g1163 ( 
.A(n_983),
.B(n_361),
.Y(n_1163)
);

BUFx8_ASAP7_75t_L g1164 ( 
.A(n_1115),
.Y(n_1164)
);

AOI21xp5_ASAP7_75t_L g1165 ( 
.A1(n_996),
.A2(n_739),
.B(n_770),
.Y(n_1165)
);

NAND2xp5_ASAP7_75t_SL g1166 ( 
.A(n_987),
.B(n_408),
.Y(n_1166)
);

OAI21xp5_ASAP7_75t_L g1167 ( 
.A1(n_1007),
.A2(n_710),
.B(n_742),
.Y(n_1167)
);

NAND2xp5_ASAP7_75t_SL g1168 ( 
.A(n_988),
.B(n_228),
.Y(n_1168)
);

OAI21x1_ASAP7_75t_L g1169 ( 
.A1(n_1049),
.A2(n_757),
.B(n_770),
.Y(n_1169)
);

NAND2xp5_ASAP7_75t_L g1170 ( 
.A(n_967),
.B(n_807),
.Y(n_1170)
);

NAND2xp5_ASAP7_75t_L g1171 ( 
.A(n_967),
.B(n_615),
.Y(n_1171)
);

NAND2xp5_ASAP7_75t_L g1172 ( 
.A(n_988),
.B(n_617),
.Y(n_1172)
);

AOI21x1_ASAP7_75t_L g1173 ( 
.A1(n_1110),
.A2(n_765),
.B(n_762),
.Y(n_1173)
);

NAND2xp5_ASAP7_75t_L g1174 ( 
.A(n_970),
.B(n_618),
.Y(n_1174)
);

INVx1_ASAP7_75t_L g1175 ( 
.A(n_1021),
.Y(n_1175)
);

BUFx2_ASAP7_75t_L g1176 ( 
.A(n_957),
.Y(n_1176)
);

OAI21x1_ASAP7_75t_L g1177 ( 
.A1(n_1060),
.A2(n_765),
.B(n_762),
.Y(n_1177)
);

NOR2xp33_ASAP7_75t_L g1178 ( 
.A(n_1043),
.B(n_367),
.Y(n_1178)
);

A2O1A1Ixp33_ASAP7_75t_SL g1179 ( 
.A1(n_1093),
.A2(n_596),
.B(n_605),
.C(n_586),
.Y(n_1179)
);

OAI22xp5_ASAP7_75t_L g1180 ( 
.A1(n_1010),
.A2(n_384),
.B1(n_371),
.B2(n_373),
.Y(n_1180)
);

BUFx3_ASAP7_75t_L g1181 ( 
.A(n_1098),
.Y(n_1181)
);

BUFx4f_ASAP7_75t_L g1182 ( 
.A(n_1076),
.Y(n_1182)
);

INVx1_ASAP7_75t_L g1183 ( 
.A(n_985),
.Y(n_1183)
);

NOR2xp33_ASAP7_75t_L g1184 ( 
.A(n_984),
.B(n_376),
.Y(n_1184)
);

AND2x4_ASAP7_75t_L g1185 ( 
.A(n_1041),
.B(n_1100),
.Y(n_1185)
);

NAND2xp5_ASAP7_75t_SL g1186 ( 
.A(n_1045),
.B(n_228),
.Y(n_1186)
);

AOI21xp5_ASAP7_75t_L g1187 ( 
.A1(n_954),
.A2(n_538),
.B(n_540),
.Y(n_1187)
);

OAI22xp5_ASAP7_75t_L g1188 ( 
.A1(n_1010),
.A2(n_402),
.B1(n_382),
.B2(n_419),
.Y(n_1188)
);

AOI21xp5_ASAP7_75t_L g1189 ( 
.A1(n_956),
.A2(n_538),
.B(n_540),
.Y(n_1189)
);

AOI21xp5_ASAP7_75t_L g1190 ( 
.A1(n_951),
.A2(n_538),
.B(n_540),
.Y(n_1190)
);

BUFx2_ASAP7_75t_L g1191 ( 
.A(n_1011),
.Y(n_1191)
);

HB1xp67_ASAP7_75t_L g1192 ( 
.A(n_962),
.Y(n_1192)
);

BUFx2_ASAP7_75t_L g1193 ( 
.A(n_966),
.Y(n_1193)
);

AND2x2_ASAP7_75t_L g1194 ( 
.A(n_1029),
.B(n_527),
.Y(n_1194)
);

AOI22xp5_ASAP7_75t_L g1195 ( 
.A1(n_984),
.A2(n_766),
.B1(n_752),
.B2(n_742),
.Y(n_1195)
);

O2A1O1Ixp33_ASAP7_75t_SL g1196 ( 
.A1(n_1048),
.A2(n_391),
.B(n_472),
.C(n_474),
.Y(n_1196)
);

NAND2xp5_ASAP7_75t_L g1197 ( 
.A(n_1012),
.B(n_1018),
.Y(n_1197)
);

AOI21xp5_ASAP7_75t_L g1198 ( 
.A1(n_945),
.A2(n_538),
.B(n_540),
.Y(n_1198)
);

OAI22xp5_ASAP7_75t_L g1199 ( 
.A1(n_1093),
.A2(n_411),
.B1(n_399),
.B2(n_400),
.Y(n_1199)
);

CKINVDCx5p33_ASAP7_75t_R g1200 ( 
.A(n_993),
.Y(n_1200)
);

AOI21xp5_ASAP7_75t_L g1201 ( 
.A1(n_948),
.A2(n_538),
.B(n_540),
.Y(n_1201)
);

OAI22x1_ASAP7_75t_L g1202 ( 
.A1(n_1092),
.A2(n_403),
.B1(n_409),
.B2(n_415),
.Y(n_1202)
);

OAI22xp5_ASAP7_75t_L g1203 ( 
.A1(n_1062),
.A2(n_418),
.B1(n_420),
.B2(n_596),
.Y(n_1203)
);

INVx2_ASAP7_75t_L g1204 ( 
.A(n_1075),
.Y(n_1204)
);

AOI21xp5_ASAP7_75t_L g1205 ( 
.A1(n_958),
.A2(n_544),
.B(n_752),
.Y(n_1205)
);

NAND2xp5_ASAP7_75t_L g1206 ( 
.A(n_1032),
.B(n_710),
.Y(n_1206)
);

NOR2xp33_ASAP7_75t_L g1207 ( 
.A(n_992),
.B(n_15),
.Y(n_1207)
);

AOI21xp5_ASAP7_75t_L g1208 ( 
.A1(n_1053),
.A2(n_544),
.B(n_752),
.Y(n_1208)
);

OAI22xp5_ASAP7_75t_L g1209 ( 
.A1(n_1031),
.A2(n_596),
.B1(n_582),
.B2(n_586),
.Y(n_1209)
);

INVx2_ASAP7_75t_L g1210 ( 
.A(n_1085),
.Y(n_1210)
);

OAI21xp5_ASAP7_75t_L g1211 ( 
.A1(n_949),
.A2(n_766),
.B(n_752),
.Y(n_1211)
);

OAI22xp5_ASAP7_75t_L g1212 ( 
.A1(n_1031),
.A2(n_596),
.B1(n_582),
.B2(n_586),
.Y(n_1212)
);

AOI21xp5_ASAP7_75t_L g1213 ( 
.A1(n_1117),
.A2(n_544),
.B(n_752),
.Y(n_1213)
);

NOR2xp33_ASAP7_75t_L g1214 ( 
.A(n_961),
.B(n_16),
.Y(n_1214)
);

BUFx6f_ASAP7_75t_L g1215 ( 
.A(n_1002),
.Y(n_1215)
);

AND2x2_ASAP7_75t_L g1216 ( 
.A(n_947),
.B(n_472),
.Y(n_1216)
);

NAND2x1p5_ASAP7_75t_L g1217 ( 
.A(n_1002),
.B(n_582),
.Y(n_1217)
);

NOR2xp33_ASAP7_75t_L g1218 ( 
.A(n_1067),
.B(n_17),
.Y(n_1218)
);

AOI22xp5_ASAP7_75t_L g1219 ( 
.A1(n_1095),
.A2(n_766),
.B1(n_752),
.B2(n_742),
.Y(n_1219)
);

O2A1O1Ixp33_ASAP7_75t_L g1220 ( 
.A1(n_974),
.A2(n_474),
.B(n_476),
.C(n_479),
.Y(n_1220)
);

OAI21x1_ASAP7_75t_L g1221 ( 
.A1(n_1104),
.A2(n_590),
.B(n_605),
.Y(n_1221)
);

CKINVDCx20_ASAP7_75t_R g1222 ( 
.A(n_966),
.Y(n_1222)
);

OAI22xp5_ASAP7_75t_L g1223 ( 
.A1(n_1107),
.A2(n_605),
.B1(n_590),
.B2(n_610),
.Y(n_1223)
);

A2O1A1Ixp33_ASAP7_75t_L g1224 ( 
.A1(n_1095),
.A2(n_610),
.B(n_590),
.C(n_479),
.Y(n_1224)
);

AND2x4_ASAP7_75t_L g1225 ( 
.A(n_953),
.B(n_476),
.Y(n_1225)
);

INVx1_ASAP7_75t_L g1226 ( 
.A(n_1083),
.Y(n_1226)
);

INVx1_ASAP7_75t_L g1227 ( 
.A(n_1086),
.Y(n_1227)
);

NAND2xp5_ASAP7_75t_L g1228 ( 
.A(n_952),
.B(n_710),
.Y(n_1228)
);

NAND2xp5_ASAP7_75t_SL g1229 ( 
.A(n_1045),
.B(n_319),
.Y(n_1229)
);

A2O1A1Ixp33_ASAP7_75t_L g1230 ( 
.A1(n_1125),
.A2(n_610),
.B(n_534),
.C(n_616),
.Y(n_1230)
);

BUFx3_ASAP7_75t_L g1231 ( 
.A(n_1004),
.Y(n_1231)
);

INVx1_ASAP7_75t_L g1232 ( 
.A(n_1102),
.Y(n_1232)
);

A2O1A1Ixp33_ASAP7_75t_L g1233 ( 
.A1(n_1125),
.A2(n_604),
.B(n_593),
.C(n_616),
.Y(n_1233)
);

INVx3_ASAP7_75t_L g1234 ( 
.A(n_1037),
.Y(n_1234)
);

NOR2xp33_ASAP7_75t_L g1235 ( 
.A(n_1092),
.B(n_18),
.Y(n_1235)
);

AOI21xp5_ASAP7_75t_L g1236 ( 
.A1(n_1106),
.A2(n_544),
.B(n_742),
.Y(n_1236)
);

AND2x4_ASAP7_75t_L g1237 ( 
.A(n_953),
.B(n_94),
.Y(n_1237)
);

A2O1A1Ixp33_ASAP7_75t_L g1238 ( 
.A1(n_995),
.A2(n_593),
.B(n_616),
.C(n_607),
.Y(n_1238)
);

INVx3_ASAP7_75t_L g1239 ( 
.A(n_1037),
.Y(n_1239)
);

CKINVDCx5p33_ASAP7_75t_R g1240 ( 
.A(n_1046),
.Y(n_1240)
);

INVx1_ASAP7_75t_L g1241 ( 
.A(n_1119),
.Y(n_1241)
);

INVx2_ASAP7_75t_L g1242 ( 
.A(n_964),
.Y(n_1242)
);

NAND2xp5_ASAP7_75t_L g1243 ( 
.A(n_963),
.B(n_766),
.Y(n_1243)
);

AOI22xp5_ASAP7_75t_L g1244 ( 
.A1(n_1099),
.A2(n_766),
.B1(n_319),
.B2(n_607),
.Y(n_1244)
);

INVx4_ASAP7_75t_L g1245 ( 
.A(n_1037),
.Y(n_1245)
);

A2O1A1Ixp33_ASAP7_75t_L g1246 ( 
.A1(n_1072),
.A2(n_1074),
.B(n_1034),
.C(n_1054),
.Y(n_1246)
);

BUFx8_ASAP7_75t_L g1247 ( 
.A(n_1118),
.Y(n_1247)
);

AND2x2_ASAP7_75t_L g1248 ( 
.A(n_1072),
.B(n_319),
.Y(n_1248)
);

NAND2xp5_ASAP7_75t_SL g1249 ( 
.A(n_1037),
.B(n_319),
.Y(n_1249)
);

INVx4_ASAP7_75t_L g1250 ( 
.A(n_968),
.Y(n_1250)
);

AO21x1_ASAP7_75t_L g1251 ( 
.A1(n_1048),
.A2(n_18),
.B(n_19),
.Y(n_1251)
);

NAND2x2_ASAP7_75t_L g1252 ( 
.A(n_1008),
.B(n_20),
.Y(n_1252)
);

OAI22xp5_ASAP7_75t_L g1253 ( 
.A1(n_1109),
.A2(n_616),
.B1(n_607),
.B2(n_604),
.Y(n_1253)
);

O2A1O1Ixp5_ASAP7_75t_L g1254 ( 
.A1(n_1000),
.A2(n_616),
.B(n_607),
.C(n_604),
.Y(n_1254)
);

OAI21x1_ASAP7_75t_L g1255 ( 
.A1(n_1103),
.A2(n_544),
.B(n_95),
.Y(n_1255)
);

AND2x2_ASAP7_75t_L g1256 ( 
.A(n_1019),
.B(n_616),
.Y(n_1256)
);

AOI221xp5_ASAP7_75t_L g1257 ( 
.A1(n_1058),
.A2(n_616),
.B1(n_607),
.B2(n_604),
.C(n_593),
.Y(n_1257)
);

AO21x1_ASAP7_75t_L g1258 ( 
.A1(n_1094),
.A2(n_20),
.B(n_24),
.Y(n_1258)
);

NAND2xp5_ASAP7_75t_L g1259 ( 
.A(n_965),
.B(n_616),
.Y(n_1259)
);

NAND2xp5_ASAP7_75t_L g1260 ( 
.A(n_1056),
.B(n_607),
.Y(n_1260)
);

NAND3xp33_ASAP7_75t_SL g1261 ( 
.A(n_974),
.B(n_25),
.C(n_27),
.Y(n_1261)
);

AOI21xp5_ASAP7_75t_L g1262 ( 
.A1(n_1073),
.A2(n_544),
.B(n_579),
.Y(n_1262)
);

NAND2xp5_ASAP7_75t_SL g1263 ( 
.A(n_1076),
.B(n_607),
.Y(n_1263)
);

NAND2xp5_ASAP7_75t_SL g1264 ( 
.A(n_978),
.B(n_607),
.Y(n_1264)
);

AOI21xp5_ASAP7_75t_L g1265 ( 
.A1(n_1110),
.A2(n_579),
.B(n_593),
.Y(n_1265)
);

OAI22xp5_ASAP7_75t_L g1266 ( 
.A1(n_986),
.A2(n_604),
.B1(n_593),
.B2(n_579),
.Y(n_1266)
);

A2O1A1Ixp33_ASAP7_75t_SL g1267 ( 
.A1(n_973),
.A2(n_604),
.B(n_555),
.C(n_169),
.Y(n_1267)
);

BUFx3_ASAP7_75t_L g1268 ( 
.A(n_1042),
.Y(n_1268)
);

NOR2xp33_ASAP7_75t_L g1269 ( 
.A(n_1024),
.B(n_28),
.Y(n_1269)
);

AOI21xp5_ASAP7_75t_L g1270 ( 
.A1(n_1116),
.A2(n_579),
.B(n_604),
.Y(n_1270)
);

AOI21xp5_ASAP7_75t_L g1271 ( 
.A1(n_1116),
.A2(n_579),
.B(n_604),
.Y(n_1271)
);

NAND2xp5_ASAP7_75t_L g1272 ( 
.A(n_998),
.B(n_579),
.Y(n_1272)
);

AOI21xp5_ASAP7_75t_L g1273 ( 
.A1(n_1063),
.A2(n_579),
.B(n_555),
.Y(n_1273)
);

NOR2xp33_ASAP7_75t_L g1274 ( 
.A(n_1024),
.B(n_29),
.Y(n_1274)
);

NAND2xp5_ASAP7_75t_L g1275 ( 
.A(n_998),
.B(n_579),
.Y(n_1275)
);

BUFx6f_ASAP7_75t_L g1276 ( 
.A(n_1076),
.Y(n_1276)
);

INVx2_ASAP7_75t_L g1277 ( 
.A(n_1127),
.Y(n_1277)
);

O2A1O1Ixp33_ASAP7_75t_L g1278 ( 
.A1(n_1065),
.A2(n_29),
.B(n_31),
.C(n_32),
.Y(n_1278)
);

INVx1_ASAP7_75t_L g1279 ( 
.A(n_1131),
.Y(n_1279)
);

INVx1_ASAP7_75t_L g1280 ( 
.A(n_1122),
.Y(n_1280)
);

AOI21xp5_ASAP7_75t_L g1281 ( 
.A1(n_1064),
.A2(n_555),
.B(n_211),
.Y(n_1281)
);

NOR2xp33_ASAP7_75t_R g1282 ( 
.A(n_1001),
.B(n_209),
.Y(n_1282)
);

NAND2xp5_ASAP7_75t_L g1283 ( 
.A(n_1055),
.B(n_32),
.Y(n_1283)
);

NAND2xp5_ASAP7_75t_SL g1284 ( 
.A(n_1084),
.B(n_201),
.Y(n_1284)
);

NAND2xp5_ASAP7_75t_SL g1285 ( 
.A(n_1084),
.B(n_199),
.Y(n_1285)
);

AOI21xp5_ASAP7_75t_L g1286 ( 
.A1(n_1068),
.A2(n_555),
.B(n_188),
.Y(n_1286)
);

AOI21xp5_ASAP7_75t_L g1287 ( 
.A1(n_1070),
.A2(n_555),
.B(n_182),
.Y(n_1287)
);

NAND2xp5_ASAP7_75t_L g1288 ( 
.A(n_1071),
.B(n_33),
.Y(n_1288)
);

NAND3xp33_ASAP7_75t_SL g1289 ( 
.A(n_1058),
.B(n_34),
.C(n_39),
.Y(n_1289)
);

AND2x4_ASAP7_75t_L g1290 ( 
.A(n_1084),
.B(n_181),
.Y(n_1290)
);

NOR2xp33_ASAP7_75t_L g1291 ( 
.A(n_1235),
.B(n_1096),
.Y(n_1291)
);

BUFx2_ASAP7_75t_L g1292 ( 
.A(n_1268),
.Y(n_1292)
);

AOI21xp5_ASAP7_75t_L g1293 ( 
.A1(n_1134),
.A2(n_1155),
.B(n_1141),
.Y(n_1293)
);

AOI21xp5_ASAP7_75t_L g1294 ( 
.A1(n_1149),
.A2(n_955),
.B(n_972),
.Y(n_1294)
);

AOI21xp5_ASAP7_75t_L g1295 ( 
.A1(n_1135),
.A2(n_1133),
.B(n_1238),
.Y(n_1295)
);

OAI21xp5_ASAP7_75t_L g1296 ( 
.A1(n_1170),
.A2(n_960),
.B(n_1128),
.Y(n_1296)
);

AO31x2_ASAP7_75t_L g1297 ( 
.A1(n_1233),
.A2(n_1014),
.A3(n_1033),
.B(n_1101),
.Y(n_1297)
);

CKINVDCx20_ASAP7_75t_R g1298 ( 
.A(n_1222),
.Y(n_1298)
);

OAI21xp5_ASAP7_75t_L g1299 ( 
.A1(n_1246),
.A2(n_1126),
.B(n_1130),
.Y(n_1299)
);

AO31x2_ASAP7_75t_L g1300 ( 
.A1(n_1230),
.A2(n_1101),
.A3(n_1105),
.B(n_1097),
.Y(n_1300)
);

OAI21x1_ASAP7_75t_L g1301 ( 
.A1(n_1173),
.A2(n_1112),
.B(n_1120),
.Y(n_1301)
);

BUFx6f_ASAP7_75t_L g1302 ( 
.A(n_1215),
.Y(n_1302)
);

OAI21x1_ASAP7_75t_L g1303 ( 
.A1(n_1221),
.A2(n_1111),
.B(n_1077),
.Y(n_1303)
);

BUFx2_ASAP7_75t_L g1304 ( 
.A(n_1176),
.Y(n_1304)
);

AOI21xp5_ASAP7_75t_L g1305 ( 
.A1(n_1153),
.A2(n_1039),
.B(n_1028),
.Y(n_1305)
);

AND2x4_ASAP7_75t_L g1306 ( 
.A(n_1185),
.B(n_1084),
.Y(n_1306)
);

OAI21x1_ASAP7_75t_L g1307 ( 
.A1(n_1158),
.A2(n_1087),
.B(n_1016),
.Y(n_1307)
);

INVx1_ASAP7_75t_L g1308 ( 
.A(n_1183),
.Y(n_1308)
);

AOI21xp5_ASAP7_75t_L g1309 ( 
.A1(n_1143),
.A2(n_1039),
.B(n_1028),
.Y(n_1309)
);

NOR2xp33_ASAP7_75t_SL g1310 ( 
.A(n_1235),
.B(n_982),
.Y(n_1310)
);

INVx2_ASAP7_75t_SL g1311 ( 
.A(n_1191),
.Y(n_1311)
);

AOI21xp5_ASAP7_75t_L g1312 ( 
.A1(n_1132),
.A2(n_1091),
.B(n_1052),
.Y(n_1312)
);

INVx1_ASAP7_75t_L g1313 ( 
.A(n_1197),
.Y(n_1313)
);

A2O1A1Ixp33_ASAP7_75t_L g1314 ( 
.A1(n_1269),
.A2(n_1113),
.B(n_1123),
.C(n_1114),
.Y(n_1314)
);

NAND2xp5_ASAP7_75t_SL g1315 ( 
.A(n_1184),
.B(n_1046),
.Y(n_1315)
);

INVx1_ASAP7_75t_L g1316 ( 
.A(n_1226),
.Y(n_1316)
);

NAND2xp5_ASAP7_75t_L g1317 ( 
.A(n_1194),
.B(n_1071),
.Y(n_1317)
);

AO31x2_ASAP7_75t_L g1318 ( 
.A1(n_1258),
.A2(n_1097),
.A3(n_1105),
.B(n_1061),
.Y(n_1318)
);

BUFx3_ASAP7_75t_L g1319 ( 
.A(n_1164),
.Y(n_1319)
);

A2O1A1Ixp33_ASAP7_75t_L g1320 ( 
.A1(n_1269),
.A2(n_1026),
.B(n_999),
.C(n_1001),
.Y(n_1320)
);

NAND2xp5_ASAP7_75t_SL g1321 ( 
.A(n_1184),
.B(n_1178),
.Y(n_1321)
);

AOI21xp5_ASAP7_75t_SL g1322 ( 
.A1(n_1237),
.A2(n_982),
.B(n_1059),
.Y(n_1322)
);

OAI22xp33_ASAP7_75t_L g1323 ( 
.A1(n_1274),
.A2(n_1096),
.B1(n_1023),
.B2(n_1108),
.Y(n_1323)
);

NOR2xp33_ASAP7_75t_L g1324 ( 
.A(n_1178),
.B(n_1003),
.Y(n_1324)
);

BUFx3_ASAP7_75t_L g1325 ( 
.A(n_1164),
.Y(n_1325)
);

AOI221x1_ASAP7_75t_L g1326 ( 
.A1(n_1274),
.A2(n_1261),
.B1(n_1289),
.B2(n_1142),
.C(n_1202),
.Y(n_1326)
);

NAND2xp5_ASAP7_75t_L g1327 ( 
.A(n_1171),
.B(n_1145),
.Y(n_1327)
);

OR2x6_ASAP7_75t_L g1328 ( 
.A(n_1193),
.B(n_1006),
.Y(n_1328)
);

BUFx3_ASAP7_75t_L g1329 ( 
.A(n_1139),
.Y(n_1329)
);

BUFx12f_ASAP7_75t_L g1330 ( 
.A(n_1137),
.Y(n_1330)
);

AOI21xp5_ASAP7_75t_L g1331 ( 
.A1(n_1259),
.A2(n_959),
.B(n_976),
.Y(n_1331)
);

OAI21x1_ASAP7_75t_L g1332 ( 
.A1(n_1169),
.A2(n_1027),
.B(n_1015),
.Y(n_1332)
);

AOI21xp5_ASAP7_75t_L g1333 ( 
.A1(n_1174),
.A2(n_969),
.B(n_1020),
.Y(n_1333)
);

AOI21xp5_ASAP7_75t_L g1334 ( 
.A1(n_1236),
.A2(n_990),
.B(n_994),
.Y(n_1334)
);

AOI21xp5_ASAP7_75t_L g1335 ( 
.A1(n_1167),
.A2(n_971),
.B(n_997),
.Y(n_1335)
);

NOR2xp67_ASAP7_75t_L g1336 ( 
.A(n_1240),
.B(n_1009),
.Y(n_1336)
);

AOI21xp5_ASAP7_75t_L g1337 ( 
.A1(n_1165),
.A2(n_1129),
.B(n_1124),
.Y(n_1337)
);

OAI21x1_ASAP7_75t_L g1338 ( 
.A1(n_1177),
.A2(n_1078),
.B(n_1035),
.Y(n_1338)
);

O2A1O1Ixp33_ASAP7_75t_SL g1339 ( 
.A1(n_1142),
.A2(n_999),
.B(n_1081),
.C(n_1036),
.Y(n_1339)
);

NAND2xp5_ASAP7_75t_L g1340 ( 
.A(n_1145),
.B(n_1080),
.Y(n_1340)
);

AOI21xp5_ASAP7_75t_L g1341 ( 
.A1(n_1228),
.A2(n_1079),
.B(n_1066),
.Y(n_1341)
);

OAI21xp5_ASAP7_75t_L g1342 ( 
.A1(n_1144),
.A2(n_1090),
.B(n_1088),
.Y(n_1342)
);

INVx1_ASAP7_75t_L g1343 ( 
.A(n_1280),
.Y(n_1343)
);

NAND2xp5_ASAP7_75t_SL g1344 ( 
.A(n_1248),
.B(n_1080),
.Y(n_1344)
);

INVx2_ASAP7_75t_L g1345 ( 
.A(n_1277),
.Y(n_1345)
);

O2A1O1Ixp33_ASAP7_75t_L g1346 ( 
.A1(n_1289),
.A2(n_1047),
.B(n_1044),
.C(n_1082),
.Y(n_1346)
);

OAI21x1_ASAP7_75t_L g1347 ( 
.A1(n_1262),
.A2(n_1121),
.B(n_1022),
.Y(n_1347)
);

OAI22x1_ASAP7_75t_L g1348 ( 
.A1(n_1207),
.A2(n_1047),
.B1(n_41),
.B2(n_44),
.Y(n_1348)
);

INVx1_ASAP7_75t_L g1349 ( 
.A(n_1227),
.Y(n_1349)
);

NAND2xp5_ASAP7_75t_L g1350 ( 
.A(n_1216),
.B(n_1038),
.Y(n_1350)
);

OAI22xp5_ASAP7_75t_L g1351 ( 
.A1(n_1144),
.A2(n_1030),
.B1(n_1051),
.B2(n_44),
.Y(n_1351)
);

AND2x4_ASAP7_75t_L g1352 ( 
.A(n_1185),
.B(n_179),
.Y(n_1352)
);

A2O1A1Ixp33_ASAP7_75t_L g1353 ( 
.A1(n_1207),
.A2(n_34),
.B(n_41),
.C(n_45),
.Y(n_1353)
);

AOI22xp33_ASAP7_75t_L g1354 ( 
.A1(n_1283),
.A2(n_555),
.B1(n_46),
.B2(n_48),
.Y(n_1354)
);

AOI31xp67_ASAP7_75t_L g1355 ( 
.A1(n_1263),
.A2(n_174),
.A3(n_158),
.B(n_154),
.Y(n_1355)
);

A2O1A1Ixp33_ASAP7_75t_L g1356 ( 
.A1(n_1161),
.A2(n_45),
.B(n_48),
.C(n_49),
.Y(n_1356)
);

INVx1_ASAP7_75t_L g1357 ( 
.A(n_1232),
.Y(n_1357)
);

AOI221xp5_ASAP7_75t_SL g1358 ( 
.A1(n_1180),
.A2(n_51),
.B1(n_56),
.B2(n_57),
.C(n_59),
.Y(n_1358)
);

NAND2xp5_ASAP7_75t_L g1359 ( 
.A(n_1147),
.B(n_63),
.Y(n_1359)
);

AO21x1_ASAP7_75t_L g1360 ( 
.A1(n_1263),
.A2(n_64),
.B(n_65),
.Y(n_1360)
);

INVx1_ASAP7_75t_L g1361 ( 
.A(n_1241),
.Y(n_1361)
);

INVx2_ASAP7_75t_L g1362 ( 
.A(n_1204),
.Y(n_1362)
);

AOI21xp5_ASAP7_75t_L g1363 ( 
.A1(n_1243),
.A2(n_104),
.B(n_149),
.Y(n_1363)
);

NAND2xp5_ASAP7_75t_SL g1364 ( 
.A(n_1147),
.B(n_1154),
.Y(n_1364)
);

AO31x2_ASAP7_75t_L g1365 ( 
.A1(n_1251),
.A2(n_68),
.A3(n_70),
.B(n_72),
.Y(n_1365)
);

AOI21xp5_ASAP7_75t_L g1366 ( 
.A1(n_1152),
.A2(n_114),
.B(n_143),
.Y(n_1366)
);

AOI21xp5_ASAP7_75t_L g1367 ( 
.A1(n_1152),
.A2(n_153),
.B(n_128),
.Y(n_1367)
);

BUFx2_ASAP7_75t_L g1368 ( 
.A(n_1154),
.Y(n_1368)
);

AO32x2_ASAP7_75t_L g1369 ( 
.A1(n_1253),
.A2(n_70),
.A3(n_74),
.B1(n_75),
.B2(n_76),
.Y(n_1369)
);

NAND2x1p5_ASAP7_75t_L g1370 ( 
.A(n_1250),
.B(n_124),
.Y(n_1370)
);

AO32x2_ASAP7_75t_L g1371 ( 
.A1(n_1209),
.A2(n_74),
.A3(n_75),
.B1(n_76),
.B2(n_77),
.Y(n_1371)
);

INVx1_ASAP7_75t_L g1372 ( 
.A(n_1279),
.Y(n_1372)
);

BUFx2_ASAP7_75t_L g1373 ( 
.A(n_1225),
.Y(n_1373)
);

CKINVDCx5p33_ASAP7_75t_R g1374 ( 
.A(n_1181),
.Y(n_1374)
);

INVx1_ASAP7_75t_L g1375 ( 
.A(n_1210),
.Y(n_1375)
);

AND2x6_ASAP7_75t_SL g1376 ( 
.A(n_1162),
.B(n_77),
.Y(n_1376)
);

OAI21x1_ASAP7_75t_L g1377 ( 
.A1(n_1255),
.A2(n_118),
.B(n_126),
.Y(n_1377)
);

AO32x2_ASAP7_75t_L g1378 ( 
.A1(n_1212),
.A2(n_1266),
.A3(n_1199),
.B1(n_1203),
.B2(n_1188),
.Y(n_1378)
);

OAI21x1_ASAP7_75t_L g1379 ( 
.A1(n_1190),
.A2(n_81),
.B(n_82),
.Y(n_1379)
);

INVx4_ASAP7_75t_L g1380 ( 
.A(n_1160),
.Y(n_1380)
);

AOI221x1_ASAP7_75t_L g1381 ( 
.A1(n_1261),
.A2(n_82),
.B1(n_1288),
.B2(n_1205),
.C(n_1189),
.Y(n_1381)
);

AO31x2_ASAP7_75t_L g1382 ( 
.A1(n_1224),
.A2(n_1187),
.A3(n_1213),
.B(n_1208),
.Y(n_1382)
);

AOI21xp5_ASAP7_75t_L g1383 ( 
.A1(n_1260),
.A2(n_1150),
.B(n_1264),
.Y(n_1383)
);

AOI21xp5_ASAP7_75t_L g1384 ( 
.A1(n_1211),
.A2(n_1267),
.B(n_1172),
.Y(n_1384)
);

OAI21xp5_ASAP7_75t_L g1385 ( 
.A1(n_1272),
.A2(n_1275),
.B(n_1256),
.Y(n_1385)
);

NAND2xp5_ASAP7_75t_L g1386 ( 
.A(n_1218),
.B(n_1192),
.Y(n_1386)
);

OAI21x1_ASAP7_75t_L g1387 ( 
.A1(n_1265),
.A2(n_1271),
.B(n_1270),
.Y(n_1387)
);

INVx1_ASAP7_75t_SL g1388 ( 
.A(n_1225),
.Y(n_1388)
);

AND2x6_ASAP7_75t_L g1389 ( 
.A(n_1290),
.B(n_1276),
.Y(n_1389)
);

BUFx3_ASAP7_75t_L g1390 ( 
.A(n_1139),
.Y(n_1390)
);

INVx2_ASAP7_75t_L g1391 ( 
.A(n_1138),
.Y(n_1391)
);

AOI221x1_ASAP7_75t_L g1392 ( 
.A1(n_1218),
.A2(n_1214),
.B1(n_1281),
.B2(n_1287),
.C(n_1286),
.Y(n_1392)
);

A2O1A1Ixp33_ASAP7_75t_L g1393 ( 
.A1(n_1278),
.A2(n_1214),
.B(n_1163),
.C(n_1249),
.Y(n_1393)
);

OAI21x1_ASAP7_75t_SL g1394 ( 
.A1(n_1250),
.A2(n_1220),
.B(n_1206),
.Y(n_1394)
);

AOI21xp5_ASAP7_75t_L g1395 ( 
.A1(n_1267),
.A2(n_1166),
.B(n_1179),
.Y(n_1395)
);

AOI21xp5_ASAP7_75t_L g1396 ( 
.A1(n_1179),
.A2(n_1285),
.B(n_1182),
.Y(n_1396)
);

INVx4_ASAP7_75t_L g1397 ( 
.A(n_1160),
.Y(n_1397)
);

OAI21x1_ASAP7_75t_L g1398 ( 
.A1(n_1273),
.A2(n_1217),
.B(n_1198),
.Y(n_1398)
);

OAI21xp5_ASAP7_75t_SL g1399 ( 
.A1(n_1162),
.A2(n_1163),
.B(n_1229),
.Y(n_1399)
);

INVx5_ASAP7_75t_L g1400 ( 
.A(n_1215),
.Y(n_1400)
);

BUFx10_ASAP7_75t_L g1401 ( 
.A(n_1200),
.Y(n_1401)
);

NAND2xp5_ASAP7_75t_L g1402 ( 
.A(n_1192),
.B(n_1140),
.Y(n_1402)
);

NAND2xp5_ASAP7_75t_L g1403 ( 
.A(n_1140),
.B(n_1146),
.Y(n_1403)
);

INVx3_ASAP7_75t_L g1404 ( 
.A(n_1276),
.Y(n_1404)
);

INVx2_ASAP7_75t_L g1405 ( 
.A(n_1151),
.Y(n_1405)
);

AO31x2_ASAP7_75t_L g1406 ( 
.A1(n_1223),
.A2(n_1201),
.A3(n_1175),
.B(n_1242),
.Y(n_1406)
);

AOI21xp5_ASAP7_75t_L g1407 ( 
.A1(n_1285),
.A2(n_1182),
.B(n_1249),
.Y(n_1407)
);

O2A1O1Ixp33_ASAP7_75t_SL g1408 ( 
.A1(n_1284),
.A2(n_1186),
.B(n_1168),
.C(n_1219),
.Y(n_1408)
);

AO31x2_ASAP7_75t_L g1409 ( 
.A1(n_1156),
.A2(n_1159),
.A3(n_1254),
.B(n_1245),
.Y(n_1409)
);

AOI21xp5_ASAP7_75t_L g1410 ( 
.A1(n_1148),
.A2(n_1290),
.B(n_1254),
.Y(n_1410)
);

AOI21xp5_ASAP7_75t_L g1411 ( 
.A1(n_1148),
.A2(n_1237),
.B(n_1217),
.Y(n_1411)
);

AOI21xp5_ASAP7_75t_L g1412 ( 
.A1(n_1148),
.A2(n_1215),
.B(n_1257),
.Y(n_1412)
);

OAI21x1_ASAP7_75t_L g1413 ( 
.A1(n_1136),
.A2(n_1157),
.B(n_1239),
.Y(n_1413)
);

NAND3xp33_ASAP7_75t_L g1414 ( 
.A(n_1247),
.B(n_1244),
.C(n_1196),
.Y(n_1414)
);

OAI21x1_ASAP7_75t_L g1415 ( 
.A1(n_1136),
.A2(n_1157),
.B(n_1239),
.Y(n_1415)
);

AOI21xp5_ASAP7_75t_L g1416 ( 
.A1(n_1215),
.A2(n_1245),
.B(n_1234),
.Y(n_1416)
);

AO31x2_ASAP7_75t_L g1417 ( 
.A1(n_1195),
.A2(n_1252),
.A3(n_1276),
.B(n_1234),
.Y(n_1417)
);

NAND2xp33_ASAP7_75t_SL g1418 ( 
.A(n_1282),
.B(n_1276),
.Y(n_1418)
);

BUFx2_ASAP7_75t_SL g1419 ( 
.A(n_1231),
.Y(n_1419)
);

NOR2xp33_ASAP7_75t_SL g1420 ( 
.A(n_1247),
.B(n_1160),
.Y(n_1420)
);

INVx3_ASAP7_75t_L g1421 ( 
.A(n_1282),
.Y(n_1421)
);

NAND3xp33_ASAP7_75t_SL g1422 ( 
.A(n_1252),
.B(n_788),
.C(n_781),
.Y(n_1422)
);

AOI22xp5_ASAP7_75t_L g1423 ( 
.A1(n_1235),
.A2(n_788),
.B1(n_781),
.B2(n_980),
.Y(n_1423)
);

OAI21xp5_ASAP7_75t_L g1424 ( 
.A1(n_1135),
.A2(n_1007),
.B(n_980),
.Y(n_1424)
);

AO31x2_ASAP7_75t_L g1425 ( 
.A1(n_1238),
.A2(n_1233),
.A3(n_1000),
.B(n_1014),
.Y(n_1425)
);

AO31x2_ASAP7_75t_L g1426 ( 
.A1(n_1238),
.A2(n_1233),
.A3(n_1000),
.B(n_1014),
.Y(n_1426)
);

O2A1O1Ixp33_ASAP7_75t_SL g1427 ( 
.A1(n_1246),
.A2(n_1007),
.B(n_1135),
.C(n_1235),
.Y(n_1427)
);

INVx1_ASAP7_75t_L g1428 ( 
.A(n_1183),
.Y(n_1428)
);

INVx1_ASAP7_75t_L g1429 ( 
.A(n_1183),
.Y(n_1429)
);

OAI21x1_ASAP7_75t_L g1430 ( 
.A1(n_1173),
.A2(n_1221),
.B(n_1158),
.Y(n_1430)
);

AOI221xp5_ASAP7_75t_L g1431 ( 
.A1(n_1235),
.A2(n_659),
.B1(n_711),
.B2(n_1274),
.C(n_1269),
.Y(n_1431)
);

NAND2xp5_ASAP7_75t_L g1432 ( 
.A(n_1194),
.B(n_1057),
.Y(n_1432)
);

NAND2xp5_ASAP7_75t_L g1433 ( 
.A(n_1194),
.B(n_1057),
.Y(n_1433)
);

AO31x2_ASAP7_75t_L g1434 ( 
.A1(n_1238),
.A2(n_1233),
.A3(n_1000),
.B(n_1014),
.Y(n_1434)
);

BUFx5_ASAP7_75t_L g1435 ( 
.A(n_1290),
.Y(n_1435)
);

OAI21x1_ASAP7_75t_L g1436 ( 
.A1(n_1173),
.A2(n_1221),
.B(n_1158),
.Y(n_1436)
);

AO32x2_ASAP7_75t_L g1437 ( 
.A1(n_1253),
.A2(n_1033),
.A3(n_831),
.B1(n_1212),
.B2(n_1209),
.Y(n_1437)
);

OAI21x1_ASAP7_75t_L g1438 ( 
.A1(n_1173),
.A2(n_1221),
.B(n_1158),
.Y(n_1438)
);

NAND3x1_ASAP7_75t_L g1439 ( 
.A(n_1235),
.B(n_788),
.C(n_781),
.Y(n_1439)
);

OR2x6_ASAP7_75t_L g1440 ( 
.A(n_1191),
.B(n_774),
.Y(n_1440)
);

AOI21xp5_ASAP7_75t_L g1441 ( 
.A1(n_1134),
.A2(n_720),
.B(n_652),
.Y(n_1441)
);

AND2x4_ASAP7_75t_L g1442 ( 
.A(n_1185),
.B(n_1041),
.Y(n_1442)
);

AOI22xp5_ASAP7_75t_L g1443 ( 
.A1(n_1235),
.A2(n_788),
.B1(n_781),
.B2(n_980),
.Y(n_1443)
);

AO32x2_ASAP7_75t_L g1444 ( 
.A1(n_1253),
.A2(n_1033),
.A3(n_831),
.B1(n_1212),
.B2(n_1209),
.Y(n_1444)
);

NAND2xp5_ASAP7_75t_L g1445 ( 
.A(n_1194),
.B(n_1057),
.Y(n_1445)
);

AO31x2_ASAP7_75t_L g1446 ( 
.A1(n_1238),
.A2(n_1233),
.A3(n_1000),
.B(n_1014),
.Y(n_1446)
);

BUFx8_ASAP7_75t_L g1447 ( 
.A(n_1137),
.Y(n_1447)
);

AOI22xp5_ASAP7_75t_L g1448 ( 
.A1(n_1235),
.A2(n_788),
.B1(n_781),
.B2(n_980),
.Y(n_1448)
);

AOI22xp5_ASAP7_75t_L g1449 ( 
.A1(n_1235),
.A2(n_788),
.B1(n_781),
.B2(n_980),
.Y(n_1449)
);

INVx2_ASAP7_75t_SL g1450 ( 
.A(n_1268),
.Y(n_1450)
);

O2A1O1Ixp33_ASAP7_75t_SL g1451 ( 
.A1(n_1246),
.A2(n_1007),
.B(n_1135),
.C(n_1235),
.Y(n_1451)
);

OAI21xp5_ASAP7_75t_L g1452 ( 
.A1(n_1135),
.A2(n_1007),
.B(n_980),
.Y(n_1452)
);

OAI21x1_ASAP7_75t_L g1453 ( 
.A1(n_1173),
.A2(n_1221),
.B(n_1158),
.Y(n_1453)
);

AO21x1_ASAP7_75t_L g1454 ( 
.A1(n_1235),
.A2(n_1274),
.B(n_1269),
.Y(n_1454)
);

NAND3xp33_ASAP7_75t_L g1455 ( 
.A(n_1235),
.B(n_788),
.C(n_781),
.Y(n_1455)
);

NAND2xp5_ASAP7_75t_L g1456 ( 
.A(n_1194),
.B(n_1057),
.Y(n_1456)
);

BUFx6f_ASAP7_75t_L g1457 ( 
.A(n_1215),
.Y(n_1457)
);

OAI21xp5_ASAP7_75t_L g1458 ( 
.A1(n_1135),
.A2(n_1007),
.B(n_980),
.Y(n_1458)
);

AOI21xp5_ASAP7_75t_L g1459 ( 
.A1(n_1134),
.A2(n_720),
.B(n_652),
.Y(n_1459)
);

OAI22xp33_ASAP7_75t_L g1460 ( 
.A1(n_1423),
.A2(n_1443),
.B1(n_1448),
.B2(n_1449),
.Y(n_1460)
);

BUFx2_ASAP7_75t_SL g1461 ( 
.A(n_1450),
.Y(n_1461)
);

BUFx4f_ASAP7_75t_L g1462 ( 
.A(n_1330),
.Y(n_1462)
);

OAI22xp33_ASAP7_75t_L g1463 ( 
.A1(n_1455),
.A2(n_1291),
.B1(n_1431),
.B2(n_1424),
.Y(n_1463)
);

INVx1_ASAP7_75t_SL g1464 ( 
.A(n_1304),
.Y(n_1464)
);

AOI22xp33_ASAP7_75t_SL g1465 ( 
.A1(n_1452),
.A2(n_1458),
.B1(n_1310),
.B2(n_1439),
.Y(n_1465)
);

OAI22xp33_ASAP7_75t_L g1466 ( 
.A1(n_1326),
.A2(n_1321),
.B1(n_1456),
.B2(n_1432),
.Y(n_1466)
);

NAND2x1p5_ASAP7_75t_L g1467 ( 
.A(n_1400),
.B(n_1380),
.Y(n_1467)
);

AND2x2_ASAP7_75t_L g1468 ( 
.A(n_1433),
.B(n_1445),
.Y(n_1468)
);

CKINVDCx11_ASAP7_75t_R g1469 ( 
.A(n_1401),
.Y(n_1469)
);

INVx2_ASAP7_75t_L g1470 ( 
.A(n_1349),
.Y(n_1470)
);

BUFx3_ASAP7_75t_L g1471 ( 
.A(n_1292),
.Y(n_1471)
);

INVx1_ASAP7_75t_L g1472 ( 
.A(n_1428),
.Y(n_1472)
);

BUFx4f_ASAP7_75t_SL g1473 ( 
.A(n_1447),
.Y(n_1473)
);

AOI22xp5_ASAP7_75t_L g1474 ( 
.A1(n_1315),
.A2(n_1454),
.B1(n_1422),
.B2(n_1399),
.Y(n_1474)
);

AOI22xp5_ASAP7_75t_L g1475 ( 
.A1(n_1344),
.A2(n_1340),
.B1(n_1324),
.B2(n_1336),
.Y(n_1475)
);

INVx1_ASAP7_75t_L g1476 ( 
.A(n_1429),
.Y(n_1476)
);

INVx1_ASAP7_75t_L g1477 ( 
.A(n_1349),
.Y(n_1477)
);

OAI22xp5_ASAP7_75t_L g1478 ( 
.A1(n_1393),
.A2(n_1327),
.B1(n_1386),
.B2(n_1313),
.Y(n_1478)
);

HB1xp67_ASAP7_75t_L g1479 ( 
.A(n_1368),
.Y(n_1479)
);

INVx1_ASAP7_75t_L g1480 ( 
.A(n_1357),
.Y(n_1480)
);

OAI22xp5_ASAP7_75t_L g1481 ( 
.A1(n_1343),
.A2(n_1421),
.B1(n_1388),
.B2(n_1328),
.Y(n_1481)
);

INVx2_ASAP7_75t_L g1482 ( 
.A(n_1361),
.Y(n_1482)
);

CKINVDCx20_ASAP7_75t_R g1483 ( 
.A(n_1298),
.Y(n_1483)
);

INVx1_ASAP7_75t_SL g1484 ( 
.A(n_1311),
.Y(n_1484)
);

BUFx10_ASAP7_75t_L g1485 ( 
.A(n_1374),
.Y(n_1485)
);

OAI22xp33_ASAP7_75t_SL g1486 ( 
.A1(n_1359),
.A2(n_1364),
.B1(n_1343),
.B2(n_1328),
.Y(n_1486)
);

AOI22xp33_ASAP7_75t_L g1487 ( 
.A1(n_1348),
.A2(n_1296),
.B1(n_1323),
.B2(n_1317),
.Y(n_1487)
);

AOI22xp33_ASAP7_75t_L g1488 ( 
.A1(n_1360),
.A2(n_1354),
.B1(n_1295),
.B2(n_1385),
.Y(n_1488)
);

AOI22xp33_ASAP7_75t_L g1489 ( 
.A1(n_1391),
.A2(n_1405),
.B1(n_1345),
.B2(n_1435),
.Y(n_1489)
);

CKINVDCx5p33_ASAP7_75t_R g1490 ( 
.A(n_1447),
.Y(n_1490)
);

BUFx2_ASAP7_75t_SL g1491 ( 
.A(n_1380),
.Y(n_1491)
);

AOI22xp5_ASAP7_75t_L g1492 ( 
.A1(n_1421),
.A2(n_1352),
.B1(n_1420),
.B2(n_1373),
.Y(n_1492)
);

INVx1_ASAP7_75t_L g1493 ( 
.A(n_1372),
.Y(n_1493)
);

INVx5_ASAP7_75t_L g1494 ( 
.A(n_1400),
.Y(n_1494)
);

INVx1_ASAP7_75t_L g1495 ( 
.A(n_1316),
.Y(n_1495)
);

CKINVDCx5p33_ASAP7_75t_R g1496 ( 
.A(n_1401),
.Y(n_1496)
);

INVx1_ASAP7_75t_L g1497 ( 
.A(n_1375),
.Y(n_1497)
);

CKINVDCx11_ASAP7_75t_R g1498 ( 
.A(n_1329),
.Y(n_1498)
);

INVx8_ASAP7_75t_L g1499 ( 
.A(n_1389),
.Y(n_1499)
);

CKINVDCx11_ASAP7_75t_R g1500 ( 
.A(n_1390),
.Y(n_1500)
);

BUFx3_ASAP7_75t_L g1501 ( 
.A(n_1306),
.Y(n_1501)
);

NAND2x1_ASAP7_75t_L g1502 ( 
.A(n_1322),
.B(n_1389),
.Y(n_1502)
);

HB1xp67_ASAP7_75t_L g1503 ( 
.A(n_1409),
.Y(n_1503)
);

BUFx2_ASAP7_75t_L g1504 ( 
.A(n_1442),
.Y(n_1504)
);

OAI22xp5_ASAP7_75t_L g1505 ( 
.A1(n_1320),
.A2(n_1314),
.B1(n_1411),
.B2(n_1440),
.Y(n_1505)
);

AOI22xp33_ASAP7_75t_L g1506 ( 
.A1(n_1435),
.A2(n_1375),
.B1(n_1414),
.B2(n_1362),
.Y(n_1506)
);

INVx2_ASAP7_75t_SL g1507 ( 
.A(n_1319),
.Y(n_1507)
);

AOI22xp33_ASAP7_75t_SL g1508 ( 
.A1(n_1435),
.A2(n_1389),
.B1(n_1352),
.B2(n_1407),
.Y(n_1508)
);

INVx1_ASAP7_75t_SL g1509 ( 
.A(n_1442),
.Y(n_1509)
);

CKINVDCx8_ASAP7_75t_R g1510 ( 
.A(n_1419),
.Y(n_1510)
);

INVx6_ASAP7_75t_L g1511 ( 
.A(n_1397),
.Y(n_1511)
);

OAI22xp33_ASAP7_75t_L g1512 ( 
.A1(n_1381),
.A2(n_1403),
.B1(n_1402),
.B2(n_1440),
.Y(n_1512)
);

INVx1_ASAP7_75t_L g1513 ( 
.A(n_1404),
.Y(n_1513)
);

BUFx10_ASAP7_75t_L g1514 ( 
.A(n_1376),
.Y(n_1514)
);

AOI22xp5_ASAP7_75t_L g1515 ( 
.A1(n_1435),
.A2(n_1451),
.B1(n_1427),
.B2(n_1306),
.Y(n_1515)
);

INVx6_ASAP7_75t_L g1516 ( 
.A(n_1397),
.Y(n_1516)
);

CKINVDCx11_ASAP7_75t_R g1517 ( 
.A(n_1325),
.Y(n_1517)
);

INVx6_ASAP7_75t_L g1518 ( 
.A(n_1302),
.Y(n_1518)
);

AND2x2_ASAP7_75t_L g1519 ( 
.A(n_1353),
.B(n_1417),
.Y(n_1519)
);

OAI22xp5_ASAP7_75t_L g1520 ( 
.A1(n_1412),
.A2(n_1410),
.B1(n_1396),
.B2(n_1350),
.Y(n_1520)
);

BUFx6f_ASAP7_75t_L g1521 ( 
.A(n_1302),
.Y(n_1521)
);

OAI22xp33_ASAP7_75t_SL g1522 ( 
.A1(n_1370),
.A2(n_1366),
.B1(n_1367),
.B2(n_1351),
.Y(n_1522)
);

INVx2_ASAP7_75t_L g1523 ( 
.A(n_1406),
.Y(n_1523)
);

CKINVDCx6p67_ASAP7_75t_R g1524 ( 
.A(n_1302),
.Y(n_1524)
);

OAI22xp33_ASAP7_75t_L g1525 ( 
.A1(n_1392),
.A2(n_1358),
.B1(n_1371),
.B2(n_1342),
.Y(n_1525)
);

INVx2_ASAP7_75t_L g1526 ( 
.A(n_1406),
.Y(n_1526)
);

BUFx4_ASAP7_75t_R g1527 ( 
.A(n_1435),
.Y(n_1527)
);

OAI22xp5_ASAP7_75t_L g1528 ( 
.A1(n_1305),
.A2(n_1356),
.B1(n_1384),
.B2(n_1346),
.Y(n_1528)
);

INVx1_ASAP7_75t_L g1529 ( 
.A(n_1413),
.Y(n_1529)
);

OAI22xp33_ASAP7_75t_L g1530 ( 
.A1(n_1371),
.A2(n_1299),
.B1(n_1369),
.B2(n_1383),
.Y(n_1530)
);

BUFx2_ASAP7_75t_L g1531 ( 
.A(n_1457),
.Y(n_1531)
);

AOI22xp33_ASAP7_75t_L g1532 ( 
.A1(n_1418),
.A2(n_1379),
.B1(n_1363),
.B2(n_1312),
.Y(n_1532)
);

OAI22xp5_ASAP7_75t_L g1533 ( 
.A1(n_1395),
.A2(n_1294),
.B1(n_1309),
.B2(n_1335),
.Y(n_1533)
);

AOI22xp33_ASAP7_75t_SL g1534 ( 
.A1(n_1394),
.A2(n_1371),
.B1(n_1377),
.B2(n_1408),
.Y(n_1534)
);

AOI22xp33_ASAP7_75t_L g1535 ( 
.A1(n_1333),
.A2(n_1293),
.B1(n_1341),
.B2(n_1369),
.Y(n_1535)
);

AOI22xp33_ASAP7_75t_SL g1536 ( 
.A1(n_1369),
.A2(n_1378),
.B1(n_1457),
.B2(n_1334),
.Y(n_1536)
);

BUFx12f_ASAP7_75t_L g1537 ( 
.A(n_1457),
.Y(n_1537)
);

INVx4_ASAP7_75t_L g1538 ( 
.A(n_1416),
.Y(n_1538)
);

AOI22xp33_ASAP7_75t_L g1539 ( 
.A1(n_1337),
.A2(n_1331),
.B1(n_1378),
.B2(n_1398),
.Y(n_1539)
);

INVx1_ASAP7_75t_L g1540 ( 
.A(n_1415),
.Y(n_1540)
);

INVx1_ASAP7_75t_SL g1541 ( 
.A(n_1417),
.Y(n_1541)
);

AOI22xp33_ASAP7_75t_L g1542 ( 
.A1(n_1378),
.A2(n_1347),
.B1(n_1307),
.B2(n_1338),
.Y(n_1542)
);

OAI22xp5_ASAP7_75t_L g1543 ( 
.A1(n_1441),
.A2(n_1459),
.B1(n_1444),
.B2(n_1437),
.Y(n_1543)
);

INVx1_ASAP7_75t_L g1544 ( 
.A(n_1365),
.Y(n_1544)
);

INVx1_ASAP7_75t_L g1545 ( 
.A(n_1365),
.Y(n_1545)
);

BUFx2_ASAP7_75t_L g1546 ( 
.A(n_1417),
.Y(n_1546)
);

CKINVDCx20_ASAP7_75t_R g1547 ( 
.A(n_1339),
.Y(n_1547)
);

INVxp67_ASAP7_75t_SL g1548 ( 
.A(n_1387),
.Y(n_1548)
);

AOI22xp33_ASAP7_75t_L g1549 ( 
.A1(n_1332),
.A2(n_1301),
.B1(n_1365),
.B2(n_1303),
.Y(n_1549)
);

OAI22xp5_ASAP7_75t_L g1550 ( 
.A1(n_1437),
.A2(n_1444),
.B1(n_1318),
.B2(n_1425),
.Y(n_1550)
);

AOI22xp33_ASAP7_75t_SL g1551 ( 
.A1(n_1437),
.A2(n_1444),
.B1(n_1355),
.B2(n_1300),
.Y(n_1551)
);

INVx1_ASAP7_75t_SL g1552 ( 
.A(n_1430),
.Y(n_1552)
);

AOI22xp33_ASAP7_75t_L g1553 ( 
.A1(n_1436),
.A2(n_1453),
.B1(n_1438),
.B2(n_1300),
.Y(n_1553)
);

AND2x2_ASAP7_75t_L g1554 ( 
.A(n_1318),
.B(n_1300),
.Y(n_1554)
);

AOI22xp33_ASAP7_75t_SL g1555 ( 
.A1(n_1297),
.A2(n_1425),
.B1(n_1426),
.B2(n_1434),
.Y(n_1555)
);

INVx1_ASAP7_75t_L g1556 ( 
.A(n_1382),
.Y(n_1556)
);

CKINVDCx6p67_ASAP7_75t_R g1557 ( 
.A(n_1297),
.Y(n_1557)
);

INVx2_ASAP7_75t_L g1558 ( 
.A(n_1382),
.Y(n_1558)
);

BUFx2_ASAP7_75t_L g1559 ( 
.A(n_1425),
.Y(n_1559)
);

INVx2_ASAP7_75t_L g1560 ( 
.A(n_1426),
.Y(n_1560)
);

BUFx12f_ASAP7_75t_L g1561 ( 
.A(n_1297),
.Y(n_1561)
);

OAI22xp5_ASAP7_75t_SL g1562 ( 
.A1(n_1426),
.A2(n_1443),
.B1(n_1448),
.B2(n_1423),
.Y(n_1562)
);

OAI22xp5_ASAP7_75t_L g1563 ( 
.A1(n_1434),
.A2(n_1443),
.B1(n_1448),
.B2(n_1423),
.Y(n_1563)
);

INVx1_ASAP7_75t_L g1564 ( 
.A(n_1434),
.Y(n_1564)
);

INVxp67_ASAP7_75t_SL g1565 ( 
.A(n_1446),
.Y(n_1565)
);

BUFx2_ASAP7_75t_L g1566 ( 
.A(n_1446),
.Y(n_1566)
);

INVx6_ASAP7_75t_L g1567 ( 
.A(n_1446),
.Y(n_1567)
);

NAND2xp5_ASAP7_75t_L g1568 ( 
.A(n_1432),
.B(n_1433),
.Y(n_1568)
);

AOI22xp33_ASAP7_75t_L g1569 ( 
.A1(n_1291),
.A2(n_980),
.B1(n_1431),
.B2(n_1235),
.Y(n_1569)
);

INVx1_ASAP7_75t_L g1570 ( 
.A(n_1308),
.Y(n_1570)
);

CKINVDCx20_ASAP7_75t_R g1571 ( 
.A(n_1298),
.Y(n_1571)
);

BUFx3_ASAP7_75t_L g1572 ( 
.A(n_1292),
.Y(n_1572)
);

INVx3_ASAP7_75t_L g1573 ( 
.A(n_1380),
.Y(n_1573)
);

CKINVDCx11_ASAP7_75t_R g1574 ( 
.A(n_1330),
.Y(n_1574)
);

AOI22xp33_ASAP7_75t_L g1575 ( 
.A1(n_1291),
.A2(n_980),
.B1(n_1431),
.B2(n_1235),
.Y(n_1575)
);

BUFx3_ASAP7_75t_L g1576 ( 
.A(n_1292),
.Y(n_1576)
);

BUFx10_ASAP7_75t_L g1577 ( 
.A(n_1374),
.Y(n_1577)
);

BUFx12f_ASAP7_75t_L g1578 ( 
.A(n_1447),
.Y(n_1578)
);

AOI22xp33_ASAP7_75t_L g1579 ( 
.A1(n_1291),
.A2(n_980),
.B1(n_1431),
.B2(n_1235),
.Y(n_1579)
);

INVx6_ASAP7_75t_L g1580 ( 
.A(n_1380),
.Y(n_1580)
);

OAI22xp5_ASAP7_75t_L g1581 ( 
.A1(n_1423),
.A2(n_1448),
.B1(n_1449),
.B2(n_1443),
.Y(n_1581)
);

INVx1_ASAP7_75t_L g1582 ( 
.A(n_1308),
.Y(n_1582)
);

INVx1_ASAP7_75t_SL g1583 ( 
.A(n_1304),
.Y(n_1583)
);

CKINVDCx11_ASAP7_75t_R g1584 ( 
.A(n_1330),
.Y(n_1584)
);

OAI22xp5_ASAP7_75t_L g1585 ( 
.A1(n_1423),
.A2(n_1448),
.B1(n_1449),
.B2(n_1443),
.Y(n_1585)
);

INVx1_ASAP7_75t_L g1586 ( 
.A(n_1308),
.Y(n_1586)
);

INVx1_ASAP7_75t_L g1587 ( 
.A(n_1308),
.Y(n_1587)
);

AOI22xp33_ASAP7_75t_L g1588 ( 
.A1(n_1291),
.A2(n_980),
.B1(n_1431),
.B2(n_1235),
.Y(n_1588)
);

BUFx4_ASAP7_75t_SL g1589 ( 
.A(n_1329),
.Y(n_1589)
);

CKINVDCx6p67_ASAP7_75t_R g1590 ( 
.A(n_1330),
.Y(n_1590)
);

AOI22xp33_ASAP7_75t_L g1591 ( 
.A1(n_1291),
.A2(n_980),
.B1(n_1431),
.B2(n_1235),
.Y(n_1591)
);

INVx2_ASAP7_75t_L g1592 ( 
.A(n_1349),
.Y(n_1592)
);

NAND2xp5_ASAP7_75t_L g1593 ( 
.A(n_1432),
.B(n_1433),
.Y(n_1593)
);

INVx2_ASAP7_75t_L g1594 ( 
.A(n_1349),
.Y(n_1594)
);

AOI22xp33_ASAP7_75t_L g1595 ( 
.A1(n_1291),
.A2(n_980),
.B1(n_1431),
.B2(n_1235),
.Y(n_1595)
);

CKINVDCx5p33_ASAP7_75t_R g1596 ( 
.A(n_1298),
.Y(n_1596)
);

CKINVDCx11_ASAP7_75t_R g1597 ( 
.A(n_1330),
.Y(n_1597)
);

INVx1_ASAP7_75t_L g1598 ( 
.A(n_1308),
.Y(n_1598)
);

BUFx4_ASAP7_75t_R g1599 ( 
.A(n_1435),
.Y(n_1599)
);

INVx1_ASAP7_75t_L g1600 ( 
.A(n_1308),
.Y(n_1600)
);

AOI22xp33_ASAP7_75t_SL g1601 ( 
.A1(n_1455),
.A2(n_980),
.B1(n_1235),
.B2(n_781),
.Y(n_1601)
);

AOI22xp33_ASAP7_75t_SL g1602 ( 
.A1(n_1455),
.A2(n_980),
.B1(n_1235),
.B2(n_781),
.Y(n_1602)
);

CKINVDCx6p67_ASAP7_75t_R g1603 ( 
.A(n_1330),
.Y(n_1603)
);

CKINVDCx11_ASAP7_75t_R g1604 ( 
.A(n_1330),
.Y(n_1604)
);

NAND2x1p5_ASAP7_75t_L g1605 ( 
.A(n_1400),
.B(n_1002),
.Y(n_1605)
);

INVx1_ASAP7_75t_L g1606 ( 
.A(n_1308),
.Y(n_1606)
);

INVx6_ASAP7_75t_L g1607 ( 
.A(n_1380),
.Y(n_1607)
);

NAND2xp5_ASAP7_75t_L g1608 ( 
.A(n_1432),
.B(n_1433),
.Y(n_1608)
);

AOI22xp33_ASAP7_75t_L g1609 ( 
.A1(n_1291),
.A2(n_980),
.B1(n_1431),
.B2(n_1235),
.Y(n_1609)
);

BUFx3_ASAP7_75t_L g1610 ( 
.A(n_1292),
.Y(n_1610)
);

AOI22xp33_ASAP7_75t_L g1611 ( 
.A1(n_1291),
.A2(n_980),
.B1(n_1431),
.B2(n_1235),
.Y(n_1611)
);

OAI22xp5_ASAP7_75t_L g1612 ( 
.A1(n_1423),
.A2(n_1448),
.B1(n_1449),
.B2(n_1443),
.Y(n_1612)
);

INVx1_ASAP7_75t_L g1613 ( 
.A(n_1308),
.Y(n_1613)
);

INVx1_ASAP7_75t_SL g1614 ( 
.A(n_1304),
.Y(n_1614)
);

BUFx2_ASAP7_75t_L g1615 ( 
.A(n_1304),
.Y(n_1615)
);

INVx1_ASAP7_75t_L g1616 ( 
.A(n_1308),
.Y(n_1616)
);

OAI21x1_ASAP7_75t_L g1617 ( 
.A1(n_1533),
.A2(n_1549),
.B(n_1553),
.Y(n_1617)
);

BUFx2_ASAP7_75t_L g1618 ( 
.A(n_1561),
.Y(n_1618)
);

CKINVDCx5p33_ASAP7_75t_R g1619 ( 
.A(n_1596),
.Y(n_1619)
);

OAI21x1_ASAP7_75t_L g1620 ( 
.A1(n_1549),
.A2(n_1553),
.B(n_1542),
.Y(n_1620)
);

INVx2_ASAP7_75t_SL g1621 ( 
.A(n_1479),
.Y(n_1621)
);

O2A1O1Ixp33_ASAP7_75t_L g1622 ( 
.A1(n_1463),
.A2(n_1581),
.B(n_1612),
.C(n_1585),
.Y(n_1622)
);

BUFx3_ASAP7_75t_L g1623 ( 
.A(n_1499),
.Y(n_1623)
);

AND2x2_ASAP7_75t_L g1624 ( 
.A(n_1554),
.B(n_1470),
.Y(n_1624)
);

INVx1_ASAP7_75t_L g1625 ( 
.A(n_1544),
.Y(n_1625)
);

AND2x4_ASAP7_75t_L g1626 ( 
.A(n_1529),
.B(n_1540),
.Y(n_1626)
);

NAND2x1p5_ASAP7_75t_L g1627 ( 
.A(n_1502),
.B(n_1494),
.Y(n_1627)
);

INVx1_ASAP7_75t_L g1628 ( 
.A(n_1545),
.Y(n_1628)
);

INVx2_ASAP7_75t_L g1629 ( 
.A(n_1482),
.Y(n_1629)
);

O2A1O1Ixp5_ASAP7_75t_L g1630 ( 
.A1(n_1463),
.A2(n_1460),
.B(n_1525),
.C(n_1528),
.Y(n_1630)
);

OAI21x1_ASAP7_75t_L g1631 ( 
.A1(n_1542),
.A2(n_1539),
.B(n_1520),
.Y(n_1631)
);

BUFx6f_ASAP7_75t_L g1632 ( 
.A(n_1499),
.Y(n_1632)
);

AO21x1_ASAP7_75t_L g1633 ( 
.A1(n_1460),
.A2(n_1525),
.B(n_1530),
.Y(n_1633)
);

OAI21x1_ASAP7_75t_L g1634 ( 
.A1(n_1539),
.A2(n_1535),
.B(n_1532),
.Y(n_1634)
);

INVx3_ASAP7_75t_L g1635 ( 
.A(n_1567),
.Y(n_1635)
);

HB1xp67_ASAP7_75t_L g1636 ( 
.A(n_1479),
.Y(n_1636)
);

BUFx3_ASAP7_75t_L g1637 ( 
.A(n_1499),
.Y(n_1637)
);

BUFx6f_ASAP7_75t_L g1638 ( 
.A(n_1494),
.Y(n_1638)
);

BUFx2_ASAP7_75t_L g1639 ( 
.A(n_1546),
.Y(n_1639)
);

INVxp67_ASAP7_75t_L g1640 ( 
.A(n_1615),
.Y(n_1640)
);

INVx3_ASAP7_75t_SL g1641 ( 
.A(n_1496),
.Y(n_1641)
);

INVx3_ASAP7_75t_L g1642 ( 
.A(n_1567),
.Y(n_1642)
);

O2A1O1Ixp33_ASAP7_75t_SL g1643 ( 
.A1(n_1466),
.A2(n_1478),
.B(n_1512),
.C(n_1530),
.Y(n_1643)
);

NOR2x1_ASAP7_75t_SL g1644 ( 
.A(n_1505),
.B(n_1494),
.Y(n_1644)
);

OAI21x1_ASAP7_75t_L g1645 ( 
.A1(n_1535),
.A2(n_1532),
.B(n_1558),
.Y(n_1645)
);

OR2x2_ASAP7_75t_L g1646 ( 
.A(n_1556),
.B(n_1559),
.Y(n_1646)
);

INVx1_ASAP7_75t_L g1647 ( 
.A(n_1564),
.Y(n_1647)
);

INVx1_ASAP7_75t_L g1648 ( 
.A(n_1503),
.Y(n_1648)
);

AND2x4_ASAP7_75t_L g1649 ( 
.A(n_1592),
.B(n_1594),
.Y(n_1649)
);

CKINVDCx5p33_ASAP7_75t_R g1650 ( 
.A(n_1469),
.Y(n_1650)
);

INVx4_ASAP7_75t_L g1651 ( 
.A(n_1527),
.Y(n_1651)
);

INVx5_ASAP7_75t_L g1652 ( 
.A(n_1567),
.Y(n_1652)
);

OAI21x1_ASAP7_75t_L g1653 ( 
.A1(n_1558),
.A2(n_1526),
.B(n_1523),
.Y(n_1653)
);

INVx2_ASAP7_75t_L g1654 ( 
.A(n_1477),
.Y(n_1654)
);

CKINVDCx6p67_ASAP7_75t_R g1655 ( 
.A(n_1578),
.Y(n_1655)
);

AND2x4_ASAP7_75t_L g1656 ( 
.A(n_1519),
.B(n_1538),
.Y(n_1656)
);

INVx4_ASAP7_75t_L g1657 ( 
.A(n_1527),
.Y(n_1657)
);

INVx2_ASAP7_75t_L g1658 ( 
.A(n_1480),
.Y(n_1658)
);

AOI22xp33_ASAP7_75t_L g1659 ( 
.A1(n_1569),
.A2(n_1611),
.B1(n_1595),
.B2(n_1575),
.Y(n_1659)
);

NOR2xp33_ASAP7_75t_L g1660 ( 
.A(n_1475),
.B(n_1468),
.Y(n_1660)
);

INVx3_ASAP7_75t_L g1661 ( 
.A(n_1560),
.Y(n_1661)
);

HB1xp67_ASAP7_75t_L g1662 ( 
.A(n_1481),
.Y(n_1662)
);

AOI22xp5_ASAP7_75t_L g1663 ( 
.A1(n_1569),
.A2(n_1595),
.B1(n_1588),
.B2(n_1591),
.Y(n_1663)
);

CKINVDCx5p33_ASAP7_75t_R g1664 ( 
.A(n_1483),
.Y(n_1664)
);

AND2x2_ASAP7_75t_L g1665 ( 
.A(n_1493),
.B(n_1541),
.Y(n_1665)
);

AOI22xp33_ASAP7_75t_SL g1666 ( 
.A1(n_1562),
.A2(n_1563),
.B1(n_1547),
.B2(n_1601),
.Y(n_1666)
);

INVx1_ASAP7_75t_L g1667 ( 
.A(n_1566),
.Y(n_1667)
);

AND2x4_ASAP7_75t_L g1668 ( 
.A(n_1538),
.B(n_1515),
.Y(n_1668)
);

AND2x2_ASAP7_75t_L g1669 ( 
.A(n_1536),
.B(n_1557),
.Y(n_1669)
);

INVx1_ASAP7_75t_L g1670 ( 
.A(n_1565),
.Y(n_1670)
);

INVx2_ASAP7_75t_L g1671 ( 
.A(n_1497),
.Y(n_1671)
);

INVx1_ASAP7_75t_L g1672 ( 
.A(n_1472),
.Y(n_1672)
);

AOI21xp5_ASAP7_75t_L g1673 ( 
.A1(n_1522),
.A2(n_1602),
.B(n_1543),
.Y(n_1673)
);

INVx2_ASAP7_75t_SL g1674 ( 
.A(n_1494),
.Y(n_1674)
);

INVx1_ASAP7_75t_L g1675 ( 
.A(n_1476),
.Y(n_1675)
);

OAI21xp5_ASAP7_75t_L g1676 ( 
.A1(n_1575),
.A2(n_1611),
.B(n_1579),
.Y(n_1676)
);

BUFx2_ASAP7_75t_L g1677 ( 
.A(n_1471),
.Y(n_1677)
);

INVx1_ASAP7_75t_L g1678 ( 
.A(n_1495),
.Y(n_1678)
);

INVx1_ASAP7_75t_L g1679 ( 
.A(n_1570),
.Y(n_1679)
);

OAI22xp5_ASAP7_75t_L g1680 ( 
.A1(n_1579),
.A2(n_1588),
.B1(n_1609),
.B2(n_1591),
.Y(n_1680)
);

BUFx2_ASAP7_75t_L g1681 ( 
.A(n_1471),
.Y(n_1681)
);

O2A1O1Ixp5_ASAP7_75t_L g1682 ( 
.A1(n_1466),
.A2(n_1512),
.B(n_1550),
.C(n_1548),
.Y(n_1682)
);

INVx1_ASAP7_75t_L g1683 ( 
.A(n_1582),
.Y(n_1683)
);

OAI21xp5_ASAP7_75t_L g1684 ( 
.A1(n_1609),
.A2(n_1474),
.B(n_1465),
.Y(n_1684)
);

INVx1_ASAP7_75t_L g1685 ( 
.A(n_1586),
.Y(n_1685)
);

AO21x2_ASAP7_75t_L g1686 ( 
.A1(n_1587),
.A2(n_1616),
.B(n_1613),
.Y(n_1686)
);

AND2x2_ASAP7_75t_L g1687 ( 
.A(n_1487),
.B(n_1555),
.Y(n_1687)
);

INVxp67_ASAP7_75t_L g1688 ( 
.A(n_1572),
.Y(n_1688)
);

BUFx3_ASAP7_75t_L g1689 ( 
.A(n_1572),
.Y(n_1689)
);

OAI21x1_ASAP7_75t_L g1690 ( 
.A1(n_1489),
.A2(n_1488),
.B(n_1506),
.Y(n_1690)
);

INVx1_ASAP7_75t_L g1691 ( 
.A(n_1598),
.Y(n_1691)
);

INVx2_ASAP7_75t_L g1692 ( 
.A(n_1600),
.Y(n_1692)
);

INVx1_ASAP7_75t_L g1693 ( 
.A(n_1606),
.Y(n_1693)
);

INVx3_ASAP7_75t_L g1694 ( 
.A(n_1552),
.Y(n_1694)
);

OAI21xp5_ASAP7_75t_L g1695 ( 
.A1(n_1488),
.A2(n_1487),
.B(n_1608),
.Y(n_1695)
);

NAND2xp5_ASAP7_75t_L g1696 ( 
.A(n_1568),
.B(n_1593),
.Y(n_1696)
);

INVx1_ASAP7_75t_L g1697 ( 
.A(n_1551),
.Y(n_1697)
);

AND2x2_ASAP7_75t_L g1698 ( 
.A(n_1534),
.B(n_1513),
.Y(n_1698)
);

INVx2_ASAP7_75t_L g1699 ( 
.A(n_1599),
.Y(n_1699)
);

OA21x2_ASAP7_75t_L g1700 ( 
.A1(n_1489),
.A2(n_1506),
.B(n_1492),
.Y(n_1700)
);

AND2x2_ASAP7_75t_L g1701 ( 
.A(n_1501),
.B(n_1504),
.Y(n_1701)
);

INVx1_ASAP7_75t_L g1702 ( 
.A(n_1486),
.Y(n_1702)
);

INVx1_ASAP7_75t_L g1703 ( 
.A(n_1508),
.Y(n_1703)
);

NAND2xp5_ASAP7_75t_L g1704 ( 
.A(n_1614),
.B(n_1583),
.Y(n_1704)
);

OA21x2_ASAP7_75t_L g1705 ( 
.A1(n_1531),
.A2(n_1509),
.B(n_1464),
.Y(n_1705)
);

OAI21x1_ASAP7_75t_L g1706 ( 
.A1(n_1605),
.A2(n_1467),
.B(n_1573),
.Y(n_1706)
);

OAI21xp5_ASAP7_75t_L g1707 ( 
.A1(n_1484),
.A2(n_1467),
.B(n_1573),
.Y(n_1707)
);

NAND2xp5_ASAP7_75t_L g1708 ( 
.A(n_1576),
.B(n_1610),
.Y(n_1708)
);

NAND2xp5_ASAP7_75t_L g1709 ( 
.A(n_1610),
.B(n_1571),
.Y(n_1709)
);

INVx1_ASAP7_75t_L g1710 ( 
.A(n_1521),
.Y(n_1710)
);

AND2x2_ASAP7_75t_L g1711 ( 
.A(n_1524),
.B(n_1518),
.Y(n_1711)
);

INVx1_ASAP7_75t_L g1712 ( 
.A(n_1518),
.Y(n_1712)
);

AND2x2_ASAP7_75t_L g1713 ( 
.A(n_1461),
.B(n_1514),
.Y(n_1713)
);

INVx4_ASAP7_75t_L g1714 ( 
.A(n_1511),
.Y(n_1714)
);

INVx1_ASAP7_75t_L g1715 ( 
.A(n_1491),
.Y(n_1715)
);

INVx2_ASAP7_75t_L g1716 ( 
.A(n_1511),
.Y(n_1716)
);

AOI22xp33_ASAP7_75t_L g1717 ( 
.A1(n_1514),
.A2(n_1507),
.B1(n_1462),
.B2(n_1473),
.Y(n_1717)
);

AND2x2_ASAP7_75t_L g1718 ( 
.A(n_1537),
.B(n_1607),
.Y(n_1718)
);

BUFx2_ASAP7_75t_L g1719 ( 
.A(n_1511),
.Y(n_1719)
);

INVx1_ASAP7_75t_L g1720 ( 
.A(n_1516),
.Y(n_1720)
);

INVx1_ASAP7_75t_L g1721 ( 
.A(n_1516),
.Y(n_1721)
);

BUFx4f_ASAP7_75t_L g1722 ( 
.A(n_1580),
.Y(n_1722)
);

HB1xp67_ASAP7_75t_L g1723 ( 
.A(n_1580),
.Y(n_1723)
);

INVx2_ASAP7_75t_L g1724 ( 
.A(n_1580),
.Y(n_1724)
);

INVx2_ASAP7_75t_L g1725 ( 
.A(n_1607),
.Y(n_1725)
);

BUFx3_ASAP7_75t_L g1726 ( 
.A(n_1510),
.Y(n_1726)
);

INVx1_ASAP7_75t_SL g1727 ( 
.A(n_1485),
.Y(n_1727)
);

OAI21xp5_ASAP7_75t_L g1728 ( 
.A1(n_1630),
.A2(n_1462),
.B(n_1490),
.Y(n_1728)
);

HB1xp67_ASAP7_75t_L g1729 ( 
.A(n_1705),
.Y(n_1729)
);

O2A1O1Ixp33_ASAP7_75t_L g1730 ( 
.A1(n_1680),
.A2(n_1589),
.B(n_1473),
.C(n_1590),
.Y(n_1730)
);

NAND4xp25_ASAP7_75t_L g1731 ( 
.A(n_1622),
.B(n_1659),
.C(n_1684),
.D(n_1660),
.Y(n_1731)
);

AND2x2_ASAP7_75t_L g1732 ( 
.A(n_1701),
.B(n_1485),
.Y(n_1732)
);

AND2x4_ASAP7_75t_L g1733 ( 
.A(n_1651),
.B(n_1657),
.Y(n_1733)
);

OR2x6_ASAP7_75t_L g1734 ( 
.A(n_1651),
.B(n_1603),
.Y(n_1734)
);

OAI21xp5_ASAP7_75t_L g1735 ( 
.A1(n_1673),
.A2(n_1577),
.B(n_1517),
.Y(n_1735)
);

CKINVDCx5p33_ASAP7_75t_R g1736 ( 
.A(n_1664),
.Y(n_1736)
);

AND2x2_ASAP7_75t_L g1737 ( 
.A(n_1702),
.B(n_1577),
.Y(n_1737)
);

A2O1A1Ixp33_ASAP7_75t_L g1738 ( 
.A1(n_1676),
.A2(n_1498),
.B(n_1500),
.C(n_1574),
.Y(n_1738)
);

INVx1_ASAP7_75t_L g1739 ( 
.A(n_1686),
.Y(n_1739)
);

INVx1_ASAP7_75t_L g1740 ( 
.A(n_1686),
.Y(n_1740)
);

OAI21xp33_ASAP7_75t_L g1741 ( 
.A1(n_1666),
.A2(n_1584),
.B(n_1597),
.Y(n_1741)
);

A2O1A1Ixp33_ASAP7_75t_SL g1742 ( 
.A1(n_1695),
.A2(n_1707),
.B(n_1663),
.C(n_1715),
.Y(n_1742)
);

NAND2xp5_ASAP7_75t_L g1743 ( 
.A(n_1624),
.B(n_1604),
.Y(n_1743)
);

AND2x2_ASAP7_75t_L g1744 ( 
.A(n_1677),
.B(n_1681),
.Y(n_1744)
);

NAND2xp5_ASAP7_75t_L g1745 ( 
.A(n_1624),
.B(n_1686),
.Y(n_1745)
);

OAI21xp5_ASAP7_75t_L g1746 ( 
.A1(n_1663),
.A2(n_1682),
.B(n_1643),
.Y(n_1746)
);

OAI211xp5_ASAP7_75t_L g1747 ( 
.A1(n_1696),
.A2(n_1687),
.B(n_1703),
.C(n_1662),
.Y(n_1747)
);

BUFx4f_ASAP7_75t_L g1748 ( 
.A(n_1655),
.Y(n_1748)
);

AOI22xp5_ASAP7_75t_L g1749 ( 
.A1(n_1703),
.A2(n_1687),
.B1(n_1633),
.B2(n_1713),
.Y(n_1749)
);

NAND2xp33_ASAP7_75t_L g1750 ( 
.A(n_1650),
.B(n_1727),
.Y(n_1750)
);

BUFx3_ASAP7_75t_L g1751 ( 
.A(n_1726),
.Y(n_1751)
);

AND2x4_ASAP7_75t_L g1752 ( 
.A(n_1651),
.B(n_1657),
.Y(n_1752)
);

AO21x1_ASAP7_75t_L g1753 ( 
.A1(n_1715),
.A2(n_1698),
.B(n_1672),
.Y(n_1753)
);

AND2x4_ASAP7_75t_L g1754 ( 
.A(n_1651),
.B(n_1657),
.Y(n_1754)
);

AND2x2_ASAP7_75t_L g1755 ( 
.A(n_1621),
.B(n_1636),
.Y(n_1755)
);

NOR2xp33_ASAP7_75t_SL g1756 ( 
.A(n_1619),
.B(n_1641),
.Y(n_1756)
);

BUFx6f_ASAP7_75t_L g1757 ( 
.A(n_1722),
.Y(n_1757)
);

A2O1A1Ixp33_ASAP7_75t_L g1758 ( 
.A1(n_1690),
.A2(n_1634),
.B(n_1631),
.C(n_1722),
.Y(n_1758)
);

A2O1A1Ixp33_ASAP7_75t_L g1759 ( 
.A1(n_1690),
.A2(n_1634),
.B(n_1631),
.C(n_1722),
.Y(n_1759)
);

BUFx2_ASAP7_75t_L g1760 ( 
.A(n_1689),
.Y(n_1760)
);

OR2x2_ASAP7_75t_L g1761 ( 
.A(n_1692),
.B(n_1705),
.Y(n_1761)
);

INVxp67_ASAP7_75t_L g1762 ( 
.A(n_1705),
.Y(n_1762)
);

INVxp67_ASAP7_75t_L g1763 ( 
.A(n_1705),
.Y(n_1763)
);

OAI22xp5_ASAP7_75t_L g1764 ( 
.A1(n_1657),
.A2(n_1697),
.B1(n_1640),
.B2(n_1699),
.Y(n_1764)
);

HB1xp67_ASAP7_75t_L g1765 ( 
.A(n_1648),
.Y(n_1765)
);

A2O1A1Ixp33_ASAP7_75t_L g1766 ( 
.A1(n_1668),
.A2(n_1726),
.B(n_1617),
.C(n_1669),
.Y(n_1766)
);

AOI21x1_ASAP7_75t_L g1767 ( 
.A1(n_1618),
.A2(n_1633),
.B(n_1670),
.Y(n_1767)
);

HB1xp67_ASAP7_75t_L g1768 ( 
.A(n_1648),
.Y(n_1768)
);

OAI21x1_ASAP7_75t_L g1769 ( 
.A1(n_1617),
.A2(n_1645),
.B(n_1653),
.Y(n_1769)
);

INVx1_ASAP7_75t_SL g1770 ( 
.A(n_1704),
.Y(n_1770)
);

OAI21xp5_ASAP7_75t_L g1771 ( 
.A1(n_1645),
.A2(n_1668),
.B(n_1700),
.Y(n_1771)
);

O2A1O1Ixp33_ASAP7_75t_L g1772 ( 
.A1(n_1688),
.A2(n_1708),
.B(n_1713),
.C(n_1641),
.Y(n_1772)
);

OAI21x1_ASAP7_75t_L g1773 ( 
.A1(n_1653),
.A2(n_1620),
.B(n_1627),
.Y(n_1773)
);

OR2x2_ASAP7_75t_L g1774 ( 
.A(n_1675),
.B(n_1678),
.Y(n_1774)
);

AND2x2_ASAP7_75t_L g1775 ( 
.A(n_1656),
.B(n_1669),
.Y(n_1775)
);

CKINVDCx5p33_ASAP7_75t_R g1776 ( 
.A(n_1655),
.Y(n_1776)
);

OR2x2_ASAP7_75t_L g1777 ( 
.A(n_1678),
.B(n_1679),
.Y(n_1777)
);

AOI221xp5_ASAP7_75t_L g1778 ( 
.A1(n_1697),
.A2(n_1685),
.B1(n_1679),
.B2(n_1683),
.C(n_1691),
.Y(n_1778)
);

OR2x2_ASAP7_75t_L g1779 ( 
.A(n_1683),
.B(n_1685),
.Y(n_1779)
);

NAND2xp5_ASAP7_75t_L g1780 ( 
.A(n_1654),
.B(n_1658),
.Y(n_1780)
);

AND2x4_ASAP7_75t_SL g1781 ( 
.A(n_1714),
.B(n_1718),
.Y(n_1781)
);

AO32x2_ASAP7_75t_L g1782 ( 
.A1(n_1674),
.A2(n_1639),
.A3(n_1714),
.B1(n_1646),
.B2(n_1667),
.Y(n_1782)
);

OAI22xp5_ASAP7_75t_L g1783 ( 
.A1(n_1726),
.A2(n_1717),
.B1(n_1700),
.B2(n_1652),
.Y(n_1783)
);

OR2x2_ASAP7_75t_L g1784 ( 
.A(n_1693),
.B(n_1646),
.Y(n_1784)
);

A2O1A1Ixp33_ASAP7_75t_L g1785 ( 
.A1(n_1668),
.A2(n_1618),
.B(n_1620),
.C(n_1637),
.Y(n_1785)
);

OR2x2_ASAP7_75t_L g1786 ( 
.A(n_1693),
.B(n_1665),
.Y(n_1786)
);

A2O1A1Ixp33_ASAP7_75t_L g1787 ( 
.A1(n_1668),
.A2(n_1652),
.B(n_1698),
.C(n_1623),
.Y(n_1787)
);

A2O1A1Ixp33_ASAP7_75t_L g1788 ( 
.A1(n_1623),
.A2(n_1637),
.B(n_1652),
.C(n_1706),
.Y(n_1788)
);

AND2x2_ASAP7_75t_L g1789 ( 
.A(n_1649),
.B(n_1710),
.Y(n_1789)
);

OAI22xp33_ASAP7_75t_L g1790 ( 
.A1(n_1700),
.A2(n_1641),
.B1(n_1652),
.B2(n_1632),
.Y(n_1790)
);

OR2x6_ASAP7_75t_L g1791 ( 
.A(n_1627),
.B(n_1635),
.Y(n_1791)
);

AND2x6_ASAP7_75t_L g1792 ( 
.A(n_1632),
.B(n_1623),
.Y(n_1792)
);

OAI22xp5_ASAP7_75t_L g1793 ( 
.A1(n_1700),
.A2(n_1652),
.B1(n_1637),
.B2(n_1671),
.Y(n_1793)
);

BUFx3_ASAP7_75t_L g1794 ( 
.A(n_1709),
.Y(n_1794)
);

INVx1_ASAP7_75t_L g1795 ( 
.A(n_1647),
.Y(n_1795)
);

NOR2xp33_ASAP7_75t_L g1796 ( 
.A(n_1720),
.B(n_1721),
.Y(n_1796)
);

NAND2xp5_ASAP7_75t_L g1797 ( 
.A(n_1649),
.B(n_1629),
.Y(n_1797)
);

AND2x2_ASAP7_75t_L g1798 ( 
.A(n_1771),
.B(n_1626),
.Y(n_1798)
);

HB1xp67_ASAP7_75t_L g1799 ( 
.A(n_1729),
.Y(n_1799)
);

AND2x4_ASAP7_75t_L g1800 ( 
.A(n_1773),
.B(n_1626),
.Y(n_1800)
);

AND2x2_ASAP7_75t_L g1801 ( 
.A(n_1771),
.B(n_1626),
.Y(n_1801)
);

INVx1_ASAP7_75t_L g1802 ( 
.A(n_1765),
.Y(n_1802)
);

OR2x2_ASAP7_75t_L g1803 ( 
.A(n_1745),
.B(n_1761),
.Y(n_1803)
);

INVx1_ASAP7_75t_L g1804 ( 
.A(n_1765),
.Y(n_1804)
);

INVx1_ASAP7_75t_L g1805 ( 
.A(n_1768),
.Y(n_1805)
);

INVx1_ASAP7_75t_L g1806 ( 
.A(n_1768),
.Y(n_1806)
);

INVx2_ASAP7_75t_L g1807 ( 
.A(n_1795),
.Y(n_1807)
);

AOI21x1_ASAP7_75t_L g1808 ( 
.A1(n_1767),
.A2(n_1628),
.B(n_1625),
.Y(n_1808)
);

AND2x2_ASAP7_75t_L g1809 ( 
.A(n_1782),
.B(n_1626),
.Y(n_1809)
);

NAND2xp5_ASAP7_75t_L g1810 ( 
.A(n_1745),
.B(n_1625),
.Y(n_1810)
);

BUFx2_ASAP7_75t_L g1811 ( 
.A(n_1782),
.Y(n_1811)
);

AND2x2_ASAP7_75t_L g1812 ( 
.A(n_1782),
.B(n_1661),
.Y(n_1812)
);

BUFx6f_ASAP7_75t_L g1813 ( 
.A(n_1769),
.Y(n_1813)
);

AND2x2_ASAP7_75t_L g1814 ( 
.A(n_1782),
.B(n_1661),
.Y(n_1814)
);

NAND2xp5_ASAP7_75t_SL g1815 ( 
.A(n_1735),
.B(n_1728),
.Y(n_1815)
);

OAI22xp5_ASAP7_75t_L g1816 ( 
.A1(n_1746),
.A2(n_1667),
.B1(n_1638),
.B2(n_1632),
.Y(n_1816)
);

AOI22xp33_ASAP7_75t_L g1817 ( 
.A1(n_1731),
.A2(n_1719),
.B1(n_1725),
.B2(n_1716),
.Y(n_1817)
);

INVxp67_ASAP7_75t_L g1818 ( 
.A(n_1729),
.Y(n_1818)
);

INVx2_ASAP7_75t_SL g1819 ( 
.A(n_1791),
.Y(n_1819)
);

HB1xp67_ASAP7_75t_L g1820 ( 
.A(n_1762),
.Y(n_1820)
);

BUFx2_ASAP7_75t_L g1821 ( 
.A(n_1762),
.Y(n_1821)
);

INVxp67_ASAP7_75t_SL g1822 ( 
.A(n_1763),
.Y(n_1822)
);

BUFx2_ASAP7_75t_L g1823 ( 
.A(n_1763),
.Y(n_1823)
);

BUFx2_ASAP7_75t_L g1824 ( 
.A(n_1760),
.Y(n_1824)
);

NOR2xp67_ASAP7_75t_L g1825 ( 
.A(n_1747),
.B(n_1694),
.Y(n_1825)
);

OR2x2_ASAP7_75t_L g1826 ( 
.A(n_1784),
.B(n_1786),
.Y(n_1826)
);

HB1xp67_ASAP7_75t_L g1827 ( 
.A(n_1755),
.Y(n_1827)
);

OAI22xp5_ASAP7_75t_L g1828 ( 
.A1(n_1746),
.A2(n_1638),
.B1(n_1632),
.B2(n_1670),
.Y(n_1828)
);

HB1xp67_ASAP7_75t_L g1829 ( 
.A(n_1739),
.Y(n_1829)
);

AOI22xp33_ASAP7_75t_L g1830 ( 
.A1(n_1735),
.A2(n_1725),
.B1(n_1716),
.B2(n_1724),
.Y(n_1830)
);

INVx4_ASAP7_75t_L g1831 ( 
.A(n_1734),
.Y(n_1831)
);

INVx1_ASAP7_75t_L g1832 ( 
.A(n_1774),
.Y(n_1832)
);

HB1xp67_ASAP7_75t_L g1833 ( 
.A(n_1740),
.Y(n_1833)
);

INVx1_ASAP7_75t_L g1834 ( 
.A(n_1777),
.Y(n_1834)
);

BUFx6f_ASAP7_75t_L g1835 ( 
.A(n_1791),
.Y(n_1835)
);

BUFx3_ASAP7_75t_L g1836 ( 
.A(n_1781),
.Y(n_1836)
);

INVx1_ASAP7_75t_L g1837 ( 
.A(n_1779),
.Y(n_1837)
);

INVx1_ASAP7_75t_L g1838 ( 
.A(n_1780),
.Y(n_1838)
);

AOI22xp33_ASAP7_75t_L g1839 ( 
.A1(n_1741),
.A2(n_1724),
.B1(n_1635),
.B2(n_1642),
.Y(n_1839)
);

BUFx6f_ASAP7_75t_L g1840 ( 
.A(n_1792),
.Y(n_1840)
);

AND2x2_ASAP7_75t_L g1841 ( 
.A(n_1758),
.B(n_1661),
.Y(n_1841)
);

AOI22xp33_ASAP7_75t_SL g1842 ( 
.A1(n_1747),
.A2(n_1644),
.B1(n_1638),
.B2(n_1627),
.Y(n_1842)
);

AOI22xp33_ASAP7_75t_L g1843 ( 
.A1(n_1728),
.A2(n_1642),
.B1(n_1632),
.B2(n_1721),
.Y(n_1843)
);

BUFx2_ASAP7_75t_L g1844 ( 
.A(n_1788),
.Y(n_1844)
);

INVx1_ASAP7_75t_L g1845 ( 
.A(n_1802),
.Y(n_1845)
);

HB1xp67_ASAP7_75t_L g1846 ( 
.A(n_1824),
.Y(n_1846)
);

BUFx3_ASAP7_75t_L g1847 ( 
.A(n_1840),
.Y(n_1847)
);

INVxp67_ASAP7_75t_L g1848 ( 
.A(n_1827),
.Y(n_1848)
);

OAI222xp33_ASAP7_75t_L g1849 ( 
.A1(n_1815),
.A2(n_1749),
.B1(n_1734),
.B2(n_1783),
.C1(n_1772),
.C2(n_1764),
.Y(n_1849)
);

INVx1_ASAP7_75t_L g1850 ( 
.A(n_1802),
.Y(n_1850)
);

AOI22xp33_ASAP7_75t_L g1851 ( 
.A1(n_1844),
.A2(n_1737),
.B1(n_1783),
.B2(n_1734),
.Y(n_1851)
);

INVx2_ASAP7_75t_SL g1852 ( 
.A(n_1824),
.Y(n_1852)
);

INVx1_ASAP7_75t_L g1853 ( 
.A(n_1804),
.Y(n_1853)
);

INVx1_ASAP7_75t_L g1854 ( 
.A(n_1804),
.Y(n_1854)
);

INVxp67_ASAP7_75t_SL g1855 ( 
.A(n_1825),
.Y(n_1855)
);

INVx1_ASAP7_75t_L g1856 ( 
.A(n_1805),
.Y(n_1856)
);

AND2x4_ASAP7_75t_L g1857 ( 
.A(n_1800),
.B(n_1785),
.Y(n_1857)
);

INVxp67_ASAP7_75t_L g1858 ( 
.A(n_1832),
.Y(n_1858)
);

AND2x4_ASAP7_75t_L g1859 ( 
.A(n_1800),
.B(n_1787),
.Y(n_1859)
);

AND2x2_ASAP7_75t_L g1860 ( 
.A(n_1809),
.B(n_1775),
.Y(n_1860)
);

INVx1_ASAP7_75t_L g1861 ( 
.A(n_1805),
.Y(n_1861)
);

INVx2_ASAP7_75t_L g1862 ( 
.A(n_1807),
.Y(n_1862)
);

OR2x2_ASAP7_75t_L g1863 ( 
.A(n_1803),
.B(n_1797),
.Y(n_1863)
);

NAND3xp33_ASAP7_75t_L g1864 ( 
.A(n_1844),
.B(n_1742),
.C(n_1730),
.Y(n_1864)
);

AOI22xp33_ASAP7_75t_L g1865 ( 
.A1(n_1830),
.A2(n_1754),
.B1(n_1752),
.B2(n_1733),
.Y(n_1865)
);

AND2x4_ASAP7_75t_L g1866 ( 
.A(n_1800),
.B(n_1787),
.Y(n_1866)
);

NAND2xp5_ASAP7_75t_L g1867 ( 
.A(n_1838),
.B(n_1770),
.Y(n_1867)
);

INVx1_ASAP7_75t_L g1868 ( 
.A(n_1806),
.Y(n_1868)
);

HB1xp67_ASAP7_75t_L g1869 ( 
.A(n_1821),
.Y(n_1869)
);

INVx1_ASAP7_75t_L g1870 ( 
.A(n_1806),
.Y(n_1870)
);

AND2x2_ASAP7_75t_L g1871 ( 
.A(n_1809),
.B(n_1744),
.Y(n_1871)
);

BUFx3_ASAP7_75t_L g1872 ( 
.A(n_1840),
.Y(n_1872)
);

NOR2x1_ASAP7_75t_L g1873 ( 
.A(n_1825),
.B(n_1790),
.Y(n_1873)
);

INVx1_ASAP7_75t_L g1874 ( 
.A(n_1829),
.Y(n_1874)
);

AND2x2_ASAP7_75t_L g1875 ( 
.A(n_1809),
.B(n_1798),
.Y(n_1875)
);

INVx1_ASAP7_75t_SL g1876 ( 
.A(n_1826),
.Y(n_1876)
);

INVx1_ASAP7_75t_L g1877 ( 
.A(n_1829),
.Y(n_1877)
);

BUFx3_ASAP7_75t_L g1878 ( 
.A(n_1840),
.Y(n_1878)
);

NAND3xp33_ASAP7_75t_SL g1879 ( 
.A(n_1842),
.B(n_1772),
.C(n_1730),
.Y(n_1879)
);

BUFx3_ASAP7_75t_L g1880 ( 
.A(n_1840),
.Y(n_1880)
);

AND2x2_ASAP7_75t_L g1881 ( 
.A(n_1798),
.B(n_1801),
.Y(n_1881)
);

AO21x2_ASAP7_75t_L g1882 ( 
.A1(n_1808),
.A2(n_1790),
.B(n_1759),
.Y(n_1882)
);

HB1xp67_ASAP7_75t_L g1883 ( 
.A(n_1821),
.Y(n_1883)
);

OR2x2_ASAP7_75t_L g1884 ( 
.A(n_1826),
.B(n_1797),
.Y(n_1884)
);

OR2x2_ASAP7_75t_L g1885 ( 
.A(n_1823),
.B(n_1820),
.Y(n_1885)
);

HB1xp67_ASAP7_75t_L g1886 ( 
.A(n_1823),
.Y(n_1886)
);

AOI22xp33_ASAP7_75t_L g1887 ( 
.A1(n_1842),
.A2(n_1752),
.B1(n_1754),
.B2(n_1733),
.Y(n_1887)
);

INVx1_ASAP7_75t_L g1888 ( 
.A(n_1833),
.Y(n_1888)
);

AND2x4_ASAP7_75t_L g1889 ( 
.A(n_1800),
.B(n_1766),
.Y(n_1889)
);

AOI211xp5_ASAP7_75t_L g1890 ( 
.A1(n_1816),
.A2(n_1742),
.B(n_1738),
.C(n_1753),
.Y(n_1890)
);

AOI221xp5_ASAP7_75t_SL g1891 ( 
.A1(n_1828),
.A2(n_1793),
.B1(n_1778),
.B2(n_1764),
.C(n_1750),
.Y(n_1891)
);

AND2x2_ASAP7_75t_L g1892 ( 
.A(n_1801),
.B(n_1789),
.Y(n_1892)
);

INVxp67_ASAP7_75t_SL g1893 ( 
.A(n_1820),
.Y(n_1893)
);

INVx1_ASAP7_75t_L g1894 ( 
.A(n_1833),
.Y(n_1894)
);

NAND4xp25_ASAP7_75t_L g1895 ( 
.A(n_1817),
.B(n_1743),
.C(n_1756),
.D(n_1796),
.Y(n_1895)
);

NOR2xp33_ASAP7_75t_L g1896 ( 
.A(n_1895),
.B(n_1776),
.Y(n_1896)
);

AND2x2_ASAP7_75t_L g1897 ( 
.A(n_1875),
.B(n_1881),
.Y(n_1897)
);

NAND2xp5_ASAP7_75t_L g1898 ( 
.A(n_1858),
.B(n_1832),
.Y(n_1898)
);

NAND2xp5_ASAP7_75t_SL g1899 ( 
.A(n_1890),
.B(n_1831),
.Y(n_1899)
);

NAND2xp5_ASAP7_75t_L g1900 ( 
.A(n_1893),
.B(n_1834),
.Y(n_1900)
);

NAND2xp5_ASAP7_75t_L g1901 ( 
.A(n_1845),
.B(n_1834),
.Y(n_1901)
);

INVx1_ASAP7_75t_L g1902 ( 
.A(n_1845),
.Y(n_1902)
);

AND2x2_ASAP7_75t_L g1903 ( 
.A(n_1875),
.B(n_1811),
.Y(n_1903)
);

NAND2xp5_ASAP7_75t_L g1904 ( 
.A(n_1850),
.B(n_1837),
.Y(n_1904)
);

INVx1_ASAP7_75t_L g1905 ( 
.A(n_1850),
.Y(n_1905)
);

AND2x2_ASAP7_75t_L g1906 ( 
.A(n_1881),
.B(n_1811),
.Y(n_1906)
);

AND2x4_ASAP7_75t_L g1907 ( 
.A(n_1859),
.B(n_1800),
.Y(n_1907)
);

AND2x2_ASAP7_75t_L g1908 ( 
.A(n_1860),
.B(n_1812),
.Y(n_1908)
);

AND2x2_ASAP7_75t_L g1909 ( 
.A(n_1860),
.B(n_1812),
.Y(n_1909)
);

HB1xp67_ASAP7_75t_L g1910 ( 
.A(n_1869),
.Y(n_1910)
);

AND2x4_ASAP7_75t_L g1911 ( 
.A(n_1859),
.B(n_1840),
.Y(n_1911)
);

INVx1_ASAP7_75t_L g1912 ( 
.A(n_1853),
.Y(n_1912)
);

INVx1_ASAP7_75t_L g1913 ( 
.A(n_1853),
.Y(n_1913)
);

INVx1_ASAP7_75t_L g1914 ( 
.A(n_1854),
.Y(n_1914)
);

NOR2xp33_ASAP7_75t_L g1915 ( 
.A(n_1895),
.B(n_1743),
.Y(n_1915)
);

NOR2xp67_ASAP7_75t_L g1916 ( 
.A(n_1864),
.B(n_1818),
.Y(n_1916)
);

INVx1_ASAP7_75t_L g1917 ( 
.A(n_1854),
.Y(n_1917)
);

AND2x2_ASAP7_75t_L g1918 ( 
.A(n_1859),
.B(n_1812),
.Y(n_1918)
);

HB1xp67_ASAP7_75t_L g1919 ( 
.A(n_1883),
.Y(n_1919)
);

HB1xp67_ASAP7_75t_L g1920 ( 
.A(n_1886),
.Y(n_1920)
);

OR2x2_ASAP7_75t_L g1921 ( 
.A(n_1885),
.B(n_1810),
.Y(n_1921)
);

INVx1_ASAP7_75t_L g1922 ( 
.A(n_1856),
.Y(n_1922)
);

NAND2xp5_ASAP7_75t_L g1923 ( 
.A(n_1856),
.B(n_1837),
.Y(n_1923)
);

INVx1_ASAP7_75t_SL g1924 ( 
.A(n_1846),
.Y(n_1924)
);

AND2x2_ASAP7_75t_L g1925 ( 
.A(n_1859),
.B(n_1814),
.Y(n_1925)
);

NOR2xp33_ASAP7_75t_L g1926 ( 
.A(n_1864),
.B(n_1748),
.Y(n_1926)
);

INVx2_ASAP7_75t_L g1927 ( 
.A(n_1862),
.Y(n_1927)
);

OR2x2_ASAP7_75t_L g1928 ( 
.A(n_1885),
.B(n_1810),
.Y(n_1928)
);

NAND2xp5_ASAP7_75t_L g1929 ( 
.A(n_1861),
.B(n_1822),
.Y(n_1929)
);

INVx3_ASAP7_75t_L g1930 ( 
.A(n_1866),
.Y(n_1930)
);

NAND2xp5_ASAP7_75t_L g1931 ( 
.A(n_1861),
.B(n_1822),
.Y(n_1931)
);

AND2x2_ASAP7_75t_L g1932 ( 
.A(n_1866),
.B(n_1814),
.Y(n_1932)
);

INVx2_ASAP7_75t_L g1933 ( 
.A(n_1862),
.Y(n_1933)
);

INVx2_ASAP7_75t_L g1934 ( 
.A(n_1862),
.Y(n_1934)
);

AND2x4_ASAP7_75t_L g1935 ( 
.A(n_1866),
.B(n_1840),
.Y(n_1935)
);

NOR2xp67_ASAP7_75t_L g1936 ( 
.A(n_1866),
.B(n_1818),
.Y(n_1936)
);

INVx1_ASAP7_75t_L g1937 ( 
.A(n_1868),
.Y(n_1937)
);

AOI22xp33_ASAP7_75t_L g1938 ( 
.A1(n_1879),
.A2(n_1831),
.B1(n_1835),
.B2(n_1839),
.Y(n_1938)
);

AND2x2_ASAP7_75t_L g1939 ( 
.A(n_1871),
.B(n_1814),
.Y(n_1939)
);

NAND2xp5_ASAP7_75t_L g1940 ( 
.A(n_1868),
.B(n_1799),
.Y(n_1940)
);

NAND2xp5_ASAP7_75t_L g1941 ( 
.A(n_1870),
.B(n_1874),
.Y(n_1941)
);

AND2x2_ASAP7_75t_L g1942 ( 
.A(n_1871),
.B(n_1841),
.Y(n_1942)
);

NOR2xp33_ASAP7_75t_L g1943 ( 
.A(n_1896),
.B(n_1748),
.Y(n_1943)
);

INVx1_ASAP7_75t_L g1944 ( 
.A(n_1902),
.Y(n_1944)
);

AND2x2_ASAP7_75t_L g1945 ( 
.A(n_1911),
.B(n_1889),
.Y(n_1945)
);

AND2x2_ASAP7_75t_L g1946 ( 
.A(n_1911),
.B(n_1889),
.Y(n_1946)
);

INVx1_ASAP7_75t_L g1947 ( 
.A(n_1902),
.Y(n_1947)
);

NAND2xp33_ASAP7_75t_SL g1948 ( 
.A(n_1899),
.B(n_1840),
.Y(n_1948)
);

INVx1_ASAP7_75t_L g1949 ( 
.A(n_1905),
.Y(n_1949)
);

INVx1_ASAP7_75t_L g1950 ( 
.A(n_1905),
.Y(n_1950)
);

INVx1_ASAP7_75t_L g1951 ( 
.A(n_1912),
.Y(n_1951)
);

OR2x2_ASAP7_75t_L g1952 ( 
.A(n_1921),
.B(n_1876),
.Y(n_1952)
);

NAND2xp5_ASAP7_75t_L g1953 ( 
.A(n_1915),
.B(n_1848),
.Y(n_1953)
);

AND2x2_ASAP7_75t_L g1954 ( 
.A(n_1911),
.B(n_1889),
.Y(n_1954)
);

INVx1_ASAP7_75t_L g1955 ( 
.A(n_1912),
.Y(n_1955)
);

INVx2_ASAP7_75t_L g1956 ( 
.A(n_1927),
.Y(n_1956)
);

OR2x2_ASAP7_75t_L g1957 ( 
.A(n_1921),
.B(n_1884),
.Y(n_1957)
);

NAND2xp5_ASAP7_75t_L g1958 ( 
.A(n_1916),
.B(n_1867),
.Y(n_1958)
);

OR2x2_ASAP7_75t_L g1959 ( 
.A(n_1928),
.B(n_1884),
.Y(n_1959)
);

INVx1_ASAP7_75t_SL g1960 ( 
.A(n_1924),
.Y(n_1960)
);

INVxp67_ASAP7_75t_SL g1961 ( 
.A(n_1916),
.Y(n_1961)
);

OR2x2_ASAP7_75t_L g1962 ( 
.A(n_1928),
.B(n_1863),
.Y(n_1962)
);

AND2x2_ASAP7_75t_L g1963 ( 
.A(n_1911),
.B(n_1889),
.Y(n_1963)
);

BUFx2_ASAP7_75t_L g1964 ( 
.A(n_1911),
.Y(n_1964)
);

INVx1_ASAP7_75t_L g1965 ( 
.A(n_1913),
.Y(n_1965)
);

HB1xp67_ASAP7_75t_L g1966 ( 
.A(n_1919),
.Y(n_1966)
);

NAND2xp5_ASAP7_75t_L g1967 ( 
.A(n_1924),
.B(n_1891),
.Y(n_1967)
);

NAND2xp5_ASAP7_75t_L g1968 ( 
.A(n_1938),
.B(n_1891),
.Y(n_1968)
);

AOI22xp33_ASAP7_75t_L g1969 ( 
.A1(n_1926),
.A2(n_1873),
.B1(n_1851),
.B2(n_1857),
.Y(n_1969)
);

INVx1_ASAP7_75t_L g1970 ( 
.A(n_1913),
.Y(n_1970)
);

NOR2x1_ASAP7_75t_L g1971 ( 
.A(n_1936),
.B(n_1873),
.Y(n_1971)
);

INVx1_ASAP7_75t_L g1972 ( 
.A(n_1914),
.Y(n_1972)
);

INVx2_ASAP7_75t_L g1973 ( 
.A(n_1927),
.Y(n_1973)
);

AND2x4_ASAP7_75t_SL g1974 ( 
.A(n_1935),
.B(n_1831),
.Y(n_1974)
);

AND2x2_ASAP7_75t_L g1975 ( 
.A(n_1935),
.B(n_1857),
.Y(n_1975)
);

INVx1_ASAP7_75t_L g1976 ( 
.A(n_1914),
.Y(n_1976)
);

AND2x2_ASAP7_75t_L g1977 ( 
.A(n_1935),
.B(n_1857),
.Y(n_1977)
);

INVx1_ASAP7_75t_L g1978 ( 
.A(n_1917),
.Y(n_1978)
);

OR2x2_ASAP7_75t_L g1979 ( 
.A(n_1929),
.B(n_1931),
.Y(n_1979)
);

OR2x2_ASAP7_75t_L g1980 ( 
.A(n_1929),
.B(n_1863),
.Y(n_1980)
);

NAND2xp5_ASAP7_75t_L g1981 ( 
.A(n_1898),
.B(n_1855),
.Y(n_1981)
);

AND2x4_ASAP7_75t_L g1982 ( 
.A(n_1935),
.B(n_1857),
.Y(n_1982)
);

NAND2xp5_ASAP7_75t_L g1983 ( 
.A(n_1898),
.B(n_1892),
.Y(n_1983)
);

INVx2_ASAP7_75t_L g1984 ( 
.A(n_1927),
.Y(n_1984)
);

AND2x2_ASAP7_75t_L g1985 ( 
.A(n_1935),
.B(n_1847),
.Y(n_1985)
);

INVx1_ASAP7_75t_L g1986 ( 
.A(n_1917),
.Y(n_1986)
);

NAND2x1p5_ASAP7_75t_L g1987 ( 
.A(n_1936),
.B(n_1847),
.Y(n_1987)
);

AND2x2_ASAP7_75t_L g1988 ( 
.A(n_1942),
.B(n_1847),
.Y(n_1988)
);

INVx1_ASAP7_75t_L g1989 ( 
.A(n_1922),
.Y(n_1989)
);

AND2x4_ASAP7_75t_L g1990 ( 
.A(n_1971),
.B(n_1930),
.Y(n_1990)
);

NAND2xp5_ASAP7_75t_L g1991 ( 
.A(n_1960),
.B(n_1942),
.Y(n_1991)
);

OR2x2_ASAP7_75t_L g1992 ( 
.A(n_1979),
.B(n_1941),
.Y(n_1992)
);

AOI22xp5_ASAP7_75t_L g1993 ( 
.A1(n_1948),
.A2(n_1968),
.B1(n_1961),
.B2(n_1967),
.Y(n_1993)
);

INVx1_ASAP7_75t_L g1994 ( 
.A(n_1944),
.Y(n_1994)
);

INVx1_ASAP7_75t_L g1995 ( 
.A(n_1944),
.Y(n_1995)
);

INVx1_ASAP7_75t_L g1996 ( 
.A(n_1947),
.Y(n_1996)
);

AND2x2_ASAP7_75t_L g1997 ( 
.A(n_1985),
.B(n_1930),
.Y(n_1997)
);

INVx1_ASAP7_75t_L g1998 ( 
.A(n_1947),
.Y(n_1998)
);

INVx1_ASAP7_75t_L g1999 ( 
.A(n_1949),
.Y(n_1999)
);

NAND2xp5_ASAP7_75t_L g2000 ( 
.A(n_1953),
.B(n_1942),
.Y(n_2000)
);

OAI21xp33_ASAP7_75t_L g2001 ( 
.A1(n_1969),
.A2(n_1890),
.B(n_1887),
.Y(n_2001)
);

NAND2xp5_ASAP7_75t_L g2002 ( 
.A(n_1958),
.B(n_1910),
.Y(n_2002)
);

NAND2xp5_ASAP7_75t_L g2003 ( 
.A(n_1985),
.B(n_1919),
.Y(n_2003)
);

INVx1_ASAP7_75t_L g2004 ( 
.A(n_1949),
.Y(n_2004)
);

NAND2xp5_ASAP7_75t_L g2005 ( 
.A(n_1981),
.B(n_1920),
.Y(n_2005)
);

INVx1_ASAP7_75t_SL g2006 ( 
.A(n_1964),
.Y(n_2006)
);

INVx1_ASAP7_75t_L g2007 ( 
.A(n_1950),
.Y(n_2007)
);

AND2x2_ASAP7_75t_L g2008 ( 
.A(n_1988),
.B(n_1930),
.Y(n_2008)
);

NAND2xp5_ASAP7_75t_SL g2009 ( 
.A(n_1987),
.B(n_1930),
.Y(n_2009)
);

NAND2xp5_ASAP7_75t_L g2010 ( 
.A(n_1964),
.B(n_1920),
.Y(n_2010)
);

OR2x2_ASAP7_75t_L g2011 ( 
.A(n_1979),
.B(n_1941),
.Y(n_2011)
);

AND2x2_ASAP7_75t_L g2012 ( 
.A(n_1988),
.B(n_1918),
.Y(n_2012)
);

AOI21xp5_ASAP7_75t_L g2013 ( 
.A1(n_1943),
.A2(n_1849),
.B(n_1882),
.Y(n_2013)
);

NOR2x1_ASAP7_75t_L g2014 ( 
.A(n_1982),
.B(n_1872),
.Y(n_2014)
);

INVx2_ASAP7_75t_L g2015 ( 
.A(n_1987),
.Y(n_2015)
);

NAND2xp5_ASAP7_75t_L g2016 ( 
.A(n_1966),
.B(n_1897),
.Y(n_2016)
);

NAND2xp5_ASAP7_75t_L g2017 ( 
.A(n_1983),
.B(n_1897),
.Y(n_2017)
);

NOR2xp67_ASAP7_75t_SL g2018 ( 
.A(n_1952),
.B(n_1831),
.Y(n_2018)
);

INVx2_ASAP7_75t_SL g2019 ( 
.A(n_1974),
.Y(n_2019)
);

AND2x2_ASAP7_75t_L g2020 ( 
.A(n_1945),
.B(n_1918),
.Y(n_2020)
);

NOR2xp67_ASAP7_75t_L g2021 ( 
.A(n_1982),
.B(n_1907),
.Y(n_2021)
);

OR2x2_ASAP7_75t_L g2022 ( 
.A(n_1952),
.B(n_1900),
.Y(n_2022)
);

NAND2xp5_ASAP7_75t_L g2023 ( 
.A(n_1975),
.B(n_1897),
.Y(n_2023)
);

INVx2_ASAP7_75t_SL g2024 ( 
.A(n_1974),
.Y(n_2024)
);

INVx1_ASAP7_75t_L g2025 ( 
.A(n_1950),
.Y(n_2025)
);

OR2x2_ASAP7_75t_L g2026 ( 
.A(n_1980),
.B(n_1900),
.Y(n_2026)
);

NOR2xp33_ASAP7_75t_L g2027 ( 
.A(n_1982),
.B(n_1736),
.Y(n_2027)
);

AND2x2_ASAP7_75t_L g2028 ( 
.A(n_1945),
.B(n_1918),
.Y(n_2028)
);

OA21x2_ASAP7_75t_L g2029 ( 
.A1(n_2009),
.A2(n_1973),
.B(n_1956),
.Y(n_2029)
);

INVx1_ASAP7_75t_L g2030 ( 
.A(n_1994),
.Y(n_2030)
);

INVx1_ASAP7_75t_L g2031 ( 
.A(n_1995),
.Y(n_2031)
);

AOI21xp5_ASAP7_75t_L g2032 ( 
.A1(n_2013),
.A2(n_1987),
.B(n_1882),
.Y(n_2032)
);

AND2x2_ASAP7_75t_L g2033 ( 
.A(n_2012),
.B(n_1975),
.Y(n_2033)
);

OR2x2_ASAP7_75t_L g2034 ( 
.A(n_1991),
.B(n_1980),
.Y(n_2034)
);

NAND2xp5_ASAP7_75t_L g2035 ( 
.A(n_2001),
.B(n_1977),
.Y(n_2035)
);

INVx2_ASAP7_75t_SL g2036 ( 
.A(n_2014),
.Y(n_2036)
);

OAI321xp33_ASAP7_75t_L g2037 ( 
.A1(n_1993),
.A2(n_1977),
.A3(n_1954),
.B1(n_1963),
.B2(n_1946),
.C(n_1816),
.Y(n_2037)
);

AOI22xp5_ASAP7_75t_L g2038 ( 
.A1(n_2019),
.A2(n_1954),
.B1(n_1946),
.B2(n_1963),
.Y(n_2038)
);

AOI211xp5_ASAP7_75t_L g2039 ( 
.A1(n_2009),
.A2(n_1828),
.B(n_1872),
.C(n_1878),
.Y(n_2039)
);

OAI221xp5_ASAP7_75t_SL g2040 ( 
.A1(n_2002),
.A2(n_1843),
.B1(n_1962),
.B2(n_1959),
.C(n_1957),
.Y(n_2040)
);

OAI22xp5_ASAP7_75t_L g2041 ( 
.A1(n_2021),
.A2(n_1880),
.B1(n_1878),
.B2(n_1872),
.Y(n_2041)
);

AOI222xp33_ASAP7_75t_L g2042 ( 
.A1(n_2005),
.A2(n_1903),
.B1(n_1906),
.B2(n_1925),
.C1(n_1932),
.C2(n_1989),
.Y(n_2042)
);

INVx1_ASAP7_75t_SL g2043 ( 
.A(n_2006),
.Y(n_2043)
);

A2O1A1Ixp33_ASAP7_75t_L g2044 ( 
.A1(n_2027),
.A2(n_1990),
.B(n_2018),
.C(n_2019),
.Y(n_2044)
);

INVx2_ASAP7_75t_L g2045 ( 
.A(n_2012),
.Y(n_2045)
);

INVx1_ASAP7_75t_L g2046 ( 
.A(n_1996),
.Y(n_2046)
);

INVx1_ASAP7_75t_L g2047 ( 
.A(n_1998),
.Y(n_2047)
);

NAND2x1_ASAP7_75t_L g2048 ( 
.A(n_1990),
.B(n_1925),
.Y(n_2048)
);

INVx1_ASAP7_75t_L g2049 ( 
.A(n_1999),
.Y(n_2049)
);

OR4x1_ASAP7_75t_L g2050 ( 
.A(n_2024),
.B(n_1986),
.C(n_1978),
.D(n_1976),
.Y(n_2050)
);

INVx1_ASAP7_75t_SL g2051 ( 
.A(n_2024),
.Y(n_2051)
);

INVxp33_ASAP7_75t_L g2052 ( 
.A(n_2027),
.Y(n_2052)
);

AOI211xp5_ASAP7_75t_L g2053 ( 
.A1(n_1990),
.A2(n_2015),
.B(n_2010),
.C(n_2003),
.Y(n_2053)
);

NOR2xp33_ASAP7_75t_L g2054 ( 
.A(n_2000),
.B(n_1962),
.Y(n_2054)
);

AOI22xp5_ASAP7_75t_L g2055 ( 
.A1(n_2016),
.A2(n_1882),
.B1(n_1907),
.B2(n_1880),
.Y(n_2055)
);

O2A1O1Ixp33_ASAP7_75t_SL g2056 ( 
.A1(n_2015),
.A2(n_1852),
.B(n_1955),
.C(n_1986),
.Y(n_2056)
);

INVx1_ASAP7_75t_L g2057 ( 
.A(n_2004),
.Y(n_2057)
);

AND2x2_ASAP7_75t_L g2058 ( 
.A(n_2033),
.B(n_2020),
.Y(n_2058)
);

AOI321xp33_ASAP7_75t_L g2059 ( 
.A1(n_2053),
.A2(n_1997),
.A3(n_2028),
.B1(n_2020),
.B2(n_2023),
.C(n_2008),
.Y(n_2059)
);

AND2x2_ASAP7_75t_L g2060 ( 
.A(n_2051),
.B(n_2028),
.Y(n_2060)
);

INVxp67_ASAP7_75t_SL g2061 ( 
.A(n_2036),
.Y(n_2061)
);

INVx1_ASAP7_75t_L g2062 ( 
.A(n_2030),
.Y(n_2062)
);

INVxp67_ASAP7_75t_L g2063 ( 
.A(n_2035),
.Y(n_2063)
);

INVxp67_ASAP7_75t_L g2064 ( 
.A(n_2043),
.Y(n_2064)
);

AOI21xp33_ASAP7_75t_L g2065 ( 
.A1(n_2052),
.A2(n_2022),
.B(n_2026),
.Y(n_2065)
);

INVx1_ASAP7_75t_L g2066 ( 
.A(n_2057),
.Y(n_2066)
);

AOI222xp33_ASAP7_75t_L g2067 ( 
.A1(n_2037),
.A2(n_2008),
.B1(n_1997),
.B2(n_2025),
.C1(n_2007),
.C2(n_2017),
.Y(n_2067)
);

AOI221xp5_ASAP7_75t_L g2068 ( 
.A1(n_2040),
.A2(n_2011),
.B1(n_1992),
.B2(n_1970),
.C(n_1978),
.Y(n_2068)
);

NOR2xp33_ASAP7_75t_L g2069 ( 
.A(n_2044),
.B(n_1992),
.Y(n_2069)
);

NAND2xp5_ASAP7_75t_L g2070 ( 
.A(n_2054),
.B(n_2011),
.Y(n_2070)
);

NOR2xp33_ASAP7_75t_L g2071 ( 
.A(n_2044),
.B(n_1957),
.Y(n_2071)
);

OR2x2_ASAP7_75t_L g2072 ( 
.A(n_2034),
.B(n_1959),
.Y(n_2072)
);

INVx1_ASAP7_75t_L g2073 ( 
.A(n_2031),
.Y(n_2073)
);

AND2x2_ASAP7_75t_L g2074 ( 
.A(n_2045),
.B(n_1907),
.Y(n_2074)
);

HB1xp67_ASAP7_75t_L g2075 ( 
.A(n_2029),
.Y(n_2075)
);

OR2x2_ASAP7_75t_L g2076 ( 
.A(n_2054),
.B(n_1951),
.Y(n_2076)
);

OAI31xp33_ASAP7_75t_SL g2077 ( 
.A1(n_2041),
.A2(n_2050),
.A3(n_2040),
.B(n_2032),
.Y(n_2077)
);

OAI22xp33_ASAP7_75t_L g2078 ( 
.A1(n_2032),
.A2(n_1878),
.B1(n_1880),
.B2(n_1835),
.Y(n_2078)
);

INVx2_ASAP7_75t_L g2079 ( 
.A(n_2048),
.Y(n_2079)
);

INVx1_ASAP7_75t_L g2080 ( 
.A(n_2046),
.Y(n_2080)
);

INVx1_ASAP7_75t_L g2081 ( 
.A(n_2075),
.Y(n_2081)
);

INVx2_ASAP7_75t_SL g2082 ( 
.A(n_2060),
.Y(n_2082)
);

INVx1_ASAP7_75t_L g2083 ( 
.A(n_2060),
.Y(n_2083)
);

XNOR2xp5_ASAP7_75t_L g2084 ( 
.A(n_2064),
.B(n_2038),
.Y(n_2084)
);

NOR2xp33_ASAP7_75t_L g2085 ( 
.A(n_2063),
.B(n_2047),
.Y(n_2085)
);

INVx2_ASAP7_75t_L g2086 ( 
.A(n_2058),
.Y(n_2086)
);

AND2x2_ASAP7_75t_L g2087 ( 
.A(n_2058),
.B(n_2039),
.Y(n_2087)
);

NAND2x1_ASAP7_75t_L g2088 ( 
.A(n_2079),
.B(n_2029),
.Y(n_2088)
);

INVx1_ASAP7_75t_L g2089 ( 
.A(n_2072),
.Y(n_2089)
);

INVx1_ASAP7_75t_L g2090 ( 
.A(n_2072),
.Y(n_2090)
);

AOI22xp5_ASAP7_75t_L g2091 ( 
.A1(n_2071),
.A2(n_2042),
.B1(n_2055),
.B2(n_2049),
.Y(n_2091)
);

AOI221xp5_ASAP7_75t_L g2092 ( 
.A1(n_2069),
.A2(n_2056),
.B1(n_1965),
.B2(n_1976),
.C(n_1951),
.Y(n_2092)
);

AOI21xp33_ASAP7_75t_L g2093 ( 
.A1(n_2077),
.A2(n_1973),
.B(n_1956),
.Y(n_2093)
);

INVx1_ASAP7_75t_L g2094 ( 
.A(n_2062),
.Y(n_2094)
);

INVx1_ASAP7_75t_L g2095 ( 
.A(n_2062),
.Y(n_2095)
);

NOR2x1_ASAP7_75t_L g2096 ( 
.A(n_2080),
.B(n_2066),
.Y(n_2096)
);

INVx2_ASAP7_75t_L g2097 ( 
.A(n_2082),
.Y(n_2097)
);

NOR3xp33_ASAP7_75t_L g2098 ( 
.A(n_2085),
.B(n_2061),
.C(n_2065),
.Y(n_2098)
);

OAI21xp5_ASAP7_75t_L g2099 ( 
.A1(n_2096),
.A2(n_2091),
.B(n_2084),
.Y(n_2099)
);

INVx1_ASAP7_75t_L g2100 ( 
.A(n_2083),
.Y(n_2100)
);

NAND3xp33_ASAP7_75t_L g2101 ( 
.A(n_2092),
.B(n_2059),
.C(n_2067),
.Y(n_2101)
);

NOR4xp25_ASAP7_75t_L g2102 ( 
.A(n_2081),
.B(n_2073),
.C(n_2080),
.D(n_2070),
.Y(n_2102)
);

AND3x1_ASAP7_75t_L g2103 ( 
.A(n_2086),
.B(n_2079),
.C(n_2068),
.Y(n_2103)
);

INVx1_ASAP7_75t_L g2104 ( 
.A(n_2089),
.Y(n_2104)
);

NOR2xp33_ASAP7_75t_L g2105 ( 
.A(n_2090),
.B(n_2076),
.Y(n_2105)
);

OAI311xp33_ASAP7_75t_L g2106 ( 
.A1(n_2092),
.A2(n_2076),
.A3(n_2074),
.B1(n_2078),
.C1(n_2056),
.Y(n_2106)
);

INVx2_ASAP7_75t_L g2107 ( 
.A(n_2088),
.Y(n_2107)
);

BUFx6f_ASAP7_75t_L g2108 ( 
.A(n_2094),
.Y(n_2108)
);

NAND2xp5_ASAP7_75t_L g2109 ( 
.A(n_2085),
.B(n_2074),
.Y(n_2109)
);

NAND2xp33_ASAP7_75t_L g2110 ( 
.A(n_2087),
.B(n_1955),
.Y(n_2110)
);

OAI211xp5_ASAP7_75t_L g2111 ( 
.A1(n_2093),
.A2(n_1751),
.B(n_1972),
.C(n_1965),
.Y(n_2111)
);

OAI211xp5_ASAP7_75t_L g2112 ( 
.A1(n_2099),
.A2(n_2093),
.B(n_2095),
.C(n_1972),
.Y(n_2112)
);

NAND3xp33_ASAP7_75t_L g2113 ( 
.A(n_2099),
.B(n_1984),
.C(n_1712),
.Y(n_2113)
);

NAND3xp33_ASAP7_75t_SL g2114 ( 
.A(n_2101),
.B(n_1865),
.C(n_1732),
.Y(n_2114)
);

AND5x1_ASAP7_75t_L g2115 ( 
.A(n_2106),
.B(n_1796),
.C(n_1984),
.D(n_1907),
.E(n_1925),
.Y(n_2115)
);

NAND2xp5_ASAP7_75t_SL g2116 ( 
.A(n_2103),
.B(n_1907),
.Y(n_2116)
);

NOR4xp75_ASAP7_75t_L g2117 ( 
.A(n_2109),
.B(n_1931),
.C(n_1932),
.D(n_1940),
.Y(n_2117)
);

OAI221xp5_ASAP7_75t_L g2118 ( 
.A1(n_2098),
.A2(n_1794),
.B1(n_1852),
.B2(n_1932),
.C(n_1940),
.Y(n_2118)
);

AOI21xp33_ASAP7_75t_SL g2119 ( 
.A1(n_2105),
.A2(n_1718),
.B(n_1906),
.Y(n_2119)
);

A2O1A1Ixp33_ASAP7_75t_L g2120 ( 
.A1(n_2111),
.A2(n_1903),
.B(n_1906),
.C(n_1937),
.Y(n_2120)
);

AOI22xp5_ASAP7_75t_L g2121 ( 
.A1(n_2114),
.A2(n_2110),
.B1(n_2097),
.B2(n_2109),
.Y(n_2121)
);

AOI22xp5_ASAP7_75t_L g2122 ( 
.A1(n_2116),
.A2(n_2104),
.B1(n_2100),
.B2(n_2107),
.Y(n_2122)
);

AOI221xp5_ASAP7_75t_L g2123 ( 
.A1(n_2112),
.A2(n_2102),
.B1(n_2108),
.B2(n_1922),
.C(n_1937),
.Y(n_2123)
);

OAI211xp5_ASAP7_75t_SL g2124 ( 
.A1(n_2118),
.A2(n_2113),
.B(n_2120),
.C(n_2115),
.Y(n_2124)
);

AOI322xp5_ASAP7_75t_L g2125 ( 
.A1(n_2117),
.A2(n_2108),
.A3(n_1903),
.B1(n_1939),
.B2(n_1908),
.C1(n_1909),
.C2(n_1799),
.Y(n_2125)
);

OAI211xp5_ASAP7_75t_L g2126 ( 
.A1(n_2119),
.A2(n_2108),
.B(n_1923),
.C(n_1901),
.Y(n_2126)
);

AOI211xp5_ASAP7_75t_L g2127 ( 
.A1(n_2112),
.A2(n_1835),
.B(n_1757),
.C(n_1793),
.Y(n_2127)
);

XNOR2x1_ASAP7_75t_L g2128 ( 
.A(n_2113),
.B(n_1711),
.Y(n_2128)
);

INVx1_ASAP7_75t_L g2129 ( 
.A(n_2122),
.Y(n_2129)
);

CKINVDCx6p67_ASAP7_75t_R g2130 ( 
.A(n_2121),
.Y(n_2130)
);

AND5x1_ASAP7_75t_L g2131 ( 
.A(n_2125),
.B(n_1835),
.C(n_1792),
.D(n_1819),
.E(n_1836),
.Y(n_2131)
);

INVx2_ASAP7_75t_SL g2132 ( 
.A(n_2128),
.Y(n_2132)
);

INVx3_ASAP7_75t_L g2133 ( 
.A(n_2126),
.Y(n_2133)
);

INVxp67_ASAP7_75t_SL g2134 ( 
.A(n_2123),
.Y(n_2134)
);

AOI211x1_ASAP7_75t_L g2135 ( 
.A1(n_2129),
.A2(n_2124),
.B(n_2127),
.C(n_1904),
.Y(n_2135)
);

OR2x6_ASAP7_75t_L g2136 ( 
.A(n_2132),
.B(n_1757),
.Y(n_2136)
);

INVx2_ASAP7_75t_L g2137 ( 
.A(n_2133),
.Y(n_2137)
);

NAND3xp33_ASAP7_75t_L g2138 ( 
.A(n_2133),
.B(n_1813),
.C(n_1901),
.Y(n_2138)
);

OAI22xp33_ASAP7_75t_L g2139 ( 
.A1(n_2137),
.A2(n_2130),
.B1(n_2134),
.B2(n_2136),
.Y(n_2139)
);

OAI211xp5_ASAP7_75t_L g2140 ( 
.A1(n_2135),
.A2(n_2134),
.B(n_2130),
.C(n_2131),
.Y(n_2140)
);

INVx1_ASAP7_75t_L g2141 ( 
.A(n_2139),
.Y(n_2141)
);

XNOR2xp5_ASAP7_75t_L g2142 ( 
.A(n_2141),
.B(n_2140),
.Y(n_2142)
);

OAI22x1_ASAP7_75t_L g2143 ( 
.A1(n_2141),
.A2(n_2138),
.B1(n_1933),
.B2(n_1934),
.Y(n_2143)
);

OAI22xp5_ASAP7_75t_L g2144 ( 
.A1(n_2142),
.A2(n_1934),
.B1(n_1933),
.B2(n_1904),
.Y(n_2144)
);

OAI22xp5_ASAP7_75t_SL g2145 ( 
.A1(n_2143),
.A2(n_1757),
.B1(n_1638),
.B2(n_1723),
.Y(n_2145)
);

AOI21xp5_ASAP7_75t_L g2146 ( 
.A1(n_2145),
.A2(n_1923),
.B(n_1934),
.Y(n_2146)
);

AOI22xp33_ASAP7_75t_L g2147 ( 
.A1(n_2144),
.A2(n_1933),
.B1(n_1888),
.B2(n_1874),
.Y(n_2147)
);

OAI21xp5_ASAP7_75t_L g2148 ( 
.A1(n_2146),
.A2(n_1908),
.B(n_1909),
.Y(n_2148)
);

OAI222xp33_ASAP7_75t_L g2149 ( 
.A1(n_2148),
.A2(n_2147),
.B1(n_1888),
.B2(n_1877),
.C1(n_1894),
.C2(n_1870),
.Y(n_2149)
);

INVx1_ASAP7_75t_L g2150 ( 
.A(n_2149),
.Y(n_2150)
);

AOI221xp5_ASAP7_75t_L g2151 ( 
.A1(n_2150),
.A2(n_1877),
.B1(n_1894),
.B2(n_1909),
.C(n_1908),
.Y(n_2151)
);

AOI211xp5_ASAP7_75t_L g2152 ( 
.A1(n_2151),
.A2(n_1711),
.B(n_1638),
.C(n_1674),
.Y(n_2152)
);


endmodule