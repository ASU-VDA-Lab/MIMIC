module fake_jpeg_20494_n_153 (n_13, n_21, n_33, n_1, n_45, n_10, n_23, n_27, n_6, n_22, n_14, n_40, n_19, n_18, n_20, n_35, n_46, n_41, n_4, n_34, n_30, n_39, n_42, n_16, n_3, n_0, n_24, n_28, n_38, n_26, n_44, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_43, n_12, n_32, n_8, n_15, n_7, n_153);

input n_13;
input n_21;
input n_33;
input n_1;
input n_45;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_46;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_42;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_44;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_43;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_153;

wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_147;
wire n_73;
wire n_152;
wire n_84;
wire n_59;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_49;
wire n_76;
wire n_127;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_103;
wire n_50;
wire n_150;
wire n_124;
wire n_141;
wire n_57;
wire n_119;
wire n_69;
wire n_83;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_106;
wire n_111;
wire n_143;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_77;
wire n_136;
wire n_61;
wire n_139;
wire n_78;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_91;
wire n_54;
wire n_93;
wire n_138;
wire n_101;
wire n_48;
wire n_149;
wire n_87;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_135;
wire n_62;
wire n_120;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_3),
.Y(n_47)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_37),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_15),
.Y(n_49)
);

BUFx2_ASAP7_75t_L g50 ( 
.A(n_29),
.Y(n_50)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_45),
.Y(n_51)
);

INVx8_ASAP7_75t_L g52 ( 
.A(n_30),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_33),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_39),
.Y(n_54)
);

INVx6_ASAP7_75t_L g55 ( 
.A(n_25),
.Y(n_55)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_38),
.Y(n_56)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_36),
.Y(n_57)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_44),
.Y(n_58)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_14),
.Y(n_59)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_5),
.Y(n_60)
);

BUFx12f_ASAP7_75t_L g61 ( 
.A(n_16),
.Y(n_61)
);

CKINVDCx20_ASAP7_75t_R g62 ( 
.A(n_34),
.Y(n_62)
);

INVx3_ASAP7_75t_L g63 ( 
.A(n_31),
.Y(n_63)
);

CKINVDCx20_ASAP7_75t_R g64 ( 
.A(n_23),
.Y(n_64)
);

INVx13_ASAP7_75t_L g65 ( 
.A(n_6),
.Y(n_65)
);

CKINVDCx20_ASAP7_75t_R g66 ( 
.A(n_1),
.Y(n_66)
);

BUFx5_ASAP7_75t_L g67 ( 
.A(n_4),
.Y(n_67)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_46),
.Y(n_68)
);

BUFx3_ASAP7_75t_L g69 ( 
.A(n_11),
.Y(n_69)
);

CKINVDCx14_ASAP7_75t_R g70 ( 
.A(n_41),
.Y(n_70)
);

CKINVDCx20_ASAP7_75t_R g71 ( 
.A(n_0),
.Y(n_71)
);

BUFx6f_ASAP7_75t_L g72 ( 
.A(n_8),
.Y(n_72)
);

BUFx5_ASAP7_75t_L g73 ( 
.A(n_19),
.Y(n_73)
);

INVx2_ASAP7_75t_R g74 ( 
.A(n_40),
.Y(n_74)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_42),
.Y(n_75)
);

BUFx3_ASAP7_75t_L g76 ( 
.A(n_61),
.Y(n_76)
);

INVx3_ASAP7_75t_SL g93 ( 
.A(n_76),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_65),
.B(n_0),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_77),
.B(n_79),
.Y(n_92)
);

BUFx6f_ASAP7_75t_L g78 ( 
.A(n_49),
.Y(n_78)
);

BUFx6f_ASAP7_75t_L g89 ( 
.A(n_78),
.Y(n_89)
);

CKINVDCx20_ASAP7_75t_R g79 ( 
.A(n_56),
.Y(n_79)
);

INVx3_ASAP7_75t_L g80 ( 
.A(n_61),
.Y(n_80)
);

INVx2_ASAP7_75t_SL g91 ( 
.A(n_80),
.Y(n_91)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_57),
.Y(n_81)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_81),
.Y(n_86)
);

BUFx12f_ASAP7_75t_L g82 ( 
.A(n_69),
.Y(n_82)
);

INVx4_ASAP7_75t_L g87 ( 
.A(n_82),
.Y(n_87)
);

NAND2x1_ASAP7_75t_SL g83 ( 
.A(n_74),
.B(n_1),
.Y(n_83)
);

OR2x2_ASAP7_75t_L g90 ( 
.A(n_83),
.B(n_74),
.Y(n_90)
);

AOI22xp33_ASAP7_75t_L g84 ( 
.A1(n_78),
.A2(n_55),
.B1(n_58),
.B2(n_63),
.Y(n_84)
);

AOI22xp5_ASAP7_75t_L g101 ( 
.A1(n_84),
.A2(n_85),
.B1(n_71),
.B2(n_60),
.Y(n_101)
);

OAI22xp5_ASAP7_75t_SL g85 ( 
.A1(n_83),
.A2(n_52),
.B1(n_70),
.B2(n_75),
.Y(n_85)
);

INVx4_ASAP7_75t_L g88 ( 
.A(n_82),
.Y(n_88)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_88),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_90),
.B(n_50),
.Y(n_105)
);

INVx3_ASAP7_75t_L g94 ( 
.A(n_82),
.Y(n_94)
);

INVx2_ASAP7_75t_L g96 ( 
.A(n_94),
.Y(n_96)
);

CKINVDCx20_ASAP7_75t_R g95 ( 
.A(n_86),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_SL g109 ( 
.A(n_95),
.B(n_97),
.Y(n_109)
);

CKINVDCx20_ASAP7_75t_R g97 ( 
.A(n_92),
.Y(n_97)
);

OAI22xp5_ASAP7_75t_L g98 ( 
.A1(n_84),
.A2(n_70),
.B1(n_59),
.B2(n_62),
.Y(n_98)
);

AOI22xp5_ASAP7_75t_L g122 ( 
.A1(n_98),
.A2(n_2),
.B1(n_4),
.B2(n_5),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_SL g99 ( 
.A(n_92),
.B(n_66),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_SL g115 ( 
.A(n_99),
.B(n_48),
.Y(n_115)
);

INVx8_ASAP7_75t_L g100 ( 
.A(n_89),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g118 ( 
.A(n_100),
.B(n_107),
.Y(n_118)
);

OAI22xp5_ASAP7_75t_SL g116 ( 
.A1(n_101),
.A2(n_91),
.B1(n_50),
.B2(n_72),
.Y(n_116)
);

MAJIxp5_ASAP7_75t_L g102 ( 
.A(n_87),
.B(n_54),
.C(n_53),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_L g112 ( 
.A(n_102),
.B(n_103),
.Y(n_112)
);

INVx2_ASAP7_75t_R g103 ( 
.A(n_93),
.Y(n_103)
);

OAI21xp5_ASAP7_75t_SL g117 ( 
.A1(n_105),
.A2(n_73),
.B(n_67),
.Y(n_117)
);

MAJIxp5_ASAP7_75t_L g106 ( 
.A(n_93),
.B(n_54),
.C(n_53),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_L g113 ( 
.A(n_106),
.B(n_76),
.Y(n_113)
);

INVx2_ASAP7_75t_L g107 ( 
.A(n_89),
.Y(n_107)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_104),
.Y(n_108)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_108),
.Y(n_124)
);

CKINVDCx20_ASAP7_75t_R g110 ( 
.A(n_103),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_SL g131 ( 
.A(n_110),
.B(n_113),
.Y(n_131)
);

INVx2_ASAP7_75t_L g111 ( 
.A(n_96),
.Y(n_111)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_111),
.Y(n_125)
);

OAI22xp5_ASAP7_75t_L g114 ( 
.A1(n_106),
.A2(n_91),
.B1(n_64),
.B2(n_51),
.Y(n_114)
);

AOI22xp5_ASAP7_75t_L g132 ( 
.A1(n_114),
.A2(n_116),
.B1(n_9),
.B2(n_12),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_L g133 ( 
.A(n_115),
.B(n_117),
.Y(n_133)
);

OAI21xp5_ASAP7_75t_L g119 ( 
.A1(n_102),
.A2(n_72),
.B(n_68),
.Y(n_119)
);

MAJIxp5_ASAP7_75t_L g129 ( 
.A(n_119),
.B(n_120),
.C(n_123),
.Y(n_129)
);

OAI21xp33_ASAP7_75t_L g120 ( 
.A1(n_100),
.A2(n_2),
.B(n_3),
.Y(n_120)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_104),
.Y(n_121)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_121),
.Y(n_134)
);

OAI22xp5_ASAP7_75t_SL g127 ( 
.A1(n_122),
.A2(n_6),
.B1(n_7),
.B2(n_8),
.Y(n_127)
);

AND2x6_ASAP7_75t_L g123 ( 
.A(n_101),
.B(n_24),
.Y(n_123)
);

OAI22xp5_ASAP7_75t_SL g126 ( 
.A1(n_112),
.A2(n_68),
.B1(n_49),
.B2(n_47),
.Y(n_126)
);

OAI22xp5_ASAP7_75t_SL g138 ( 
.A1(n_126),
.A2(n_130),
.B1(n_132),
.B2(n_120),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_L g137 ( 
.A(n_127),
.B(n_119),
.Y(n_137)
);

CKINVDCx20_ASAP7_75t_R g128 ( 
.A(n_109),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_L g136 ( 
.A(n_128),
.B(n_123),
.Y(n_136)
);

OAI22xp5_ASAP7_75t_SL g130 ( 
.A1(n_122),
.A2(n_7),
.B1(n_9),
.B2(n_10),
.Y(n_130)
);

INVx1_ASAP7_75t_SL g135 ( 
.A(n_124),
.Y(n_135)
);

CKINVDCx16_ASAP7_75t_R g142 ( 
.A(n_135),
.Y(n_142)
);

AOI22xp5_ASAP7_75t_L g141 ( 
.A1(n_136),
.A2(n_137),
.B1(n_138),
.B2(n_139),
.Y(n_141)
);

MAJIxp5_ASAP7_75t_L g139 ( 
.A(n_131),
.B(n_118),
.C(n_17),
.Y(n_139)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_134),
.Y(n_140)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_141),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_SL g144 ( 
.A(n_143),
.B(n_129),
.Y(n_144)
);

XOR2xp5_ASAP7_75t_L g145 ( 
.A(n_144),
.B(n_129),
.Y(n_145)
);

MAJIxp5_ASAP7_75t_L g146 ( 
.A(n_145),
.B(n_136),
.C(n_133),
.Y(n_146)
);

AOI21x1_ASAP7_75t_L g147 ( 
.A1(n_146),
.A2(n_142),
.B(n_140),
.Y(n_147)
);

MAJIxp5_ASAP7_75t_L g148 ( 
.A(n_147),
.B(n_125),
.C(n_132),
.Y(n_148)
);

AOI322xp5_ASAP7_75t_L g149 ( 
.A1(n_148),
.A2(n_126),
.A3(n_18),
.B1(n_20),
.B2(n_21),
.C1(n_22),
.C2(n_26),
.Y(n_149)
);

AOI21x1_ASAP7_75t_L g150 ( 
.A1(n_149),
.A2(n_13),
.B(n_27),
.Y(n_150)
);

MAJIxp5_ASAP7_75t_L g151 ( 
.A(n_150),
.B(n_28),
.C(n_32),
.Y(n_151)
);

XNOR2xp5_ASAP7_75t_L g152 ( 
.A(n_151),
.B(n_35),
.Y(n_152)
);

XOR2xp5_ASAP7_75t_L g153 ( 
.A(n_152),
.B(n_43),
.Y(n_153)
);


endmodule