module real_jpeg_15937_n_18 (n_17, n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_16, n_3, n_10, n_9, n_18);

input n_17;
input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_16;
input n_3;
input n_10;
input n_9;

output n_18;

wire n_384;
wire n_37;
wire n_430;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_300;
wire n_415;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_199;
wire n_95;
wire n_238;
wire n_67;
wire n_350;
wire n_235;
wire n_107;
wire n_369;
wire n_376;
wire n_354;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_355;
wire n_123;
wire n_425;
wire n_50;
wire n_409;
wire n_186;
wire n_137;
wire n_72;
wire n_171;
wire n_151;
wire n_272;
wire n_198;
wire n_203;
wire n_23;
wire n_362;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_326;
wire n_339;
wire n_80;
wire n_30;
wire n_332;
wire n_149;
wire n_328;
wire n_366;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_353;
wire n_230;
wire n_417;
wire n_428;
wire n_216;
wire n_128;
wire n_202;
wire n_367;
wire n_127;
wire n_356;
wire n_365;
wire n_423;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_422;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_348;
wire n_252;
wire n_363;
wire n_310;
wire n_345;
wire n_83;
wire n_78;
wire n_288;
wire n_221;
wire n_393;
wire n_104;
wire n_153;
wire n_337;
wire n_131;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_378;
wire n_200;
wire n_432;
wire n_335;
wire n_214;
wire n_113;
wire n_251;
wire n_139;
wire n_33;
wire n_175;
wire n_338;
wire n_156;
wire n_387;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_390;
wire n_77;
wire n_399;
wire n_219;
wire n_372;
wire n_122;
wire n_19;
wire n_262;
wire n_334;
wire n_383;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_426;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_371;
wire n_410;
wire n_421;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_382;
wire n_411;
wire n_20;
wire n_278;
wire n_314;
wire n_103;
wire n_232;
wire n_212;
wire n_284;
wire n_402;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_213;
wire n_25;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_407;
wire n_419;
wire n_386;
wire n_341;
wire n_331;
wire n_49;
wire n_68;
wire n_395;
wire n_146;
wire n_286;
wire n_166;
wire n_215;
wire n_176;
wire n_323;
wire n_312;
wire n_325;
wire n_307;
wire n_316;
wire n_161;
wire n_207;
wire n_431;
wire n_420;
wire n_357;
wire n_237;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_380;
wire n_414;
wire n_140;
wire n_126;
wire n_342;
wire n_120;
wire n_155;
wire n_412;
wire n_405;
wire n_319;
wire n_93;
wire n_242;
wire n_142;
wire n_397;
wire n_76;
wire n_403;
wire n_79;
wire n_282;
wire n_147;
wire n_359;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_145;
wire n_266;
wire n_377;
wire n_109;
wire n_391;
wire n_427;
wire n_401;
wire n_148;
wire n_373;
wire n_396;
wire n_392;
wire n_196;
wire n_375;
wire n_330;
wire n_298;
wire n_333;
wire n_152;
wire n_270;
wire n_159;
wire n_429;
wire n_347;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_336;
wire n_258;
wire n_150;
wire n_41;
wire n_74;
wire n_404;
wire n_158;
wire n_204;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_413;
wire n_75;
wire n_346;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_119;
wire n_283;
wire n_181;
wire n_358;
wire n_256;
wire n_273;
wire n_253;
wire n_54;
wire n_168;
wire n_38;
wire n_385;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_349;
wire n_418;
wire n_292;
wire n_343;
wire n_64;
wire n_291;
wire n_236;
wire n_370;
wire n_276;
wire n_374;
wire n_287;
wire n_388;
wire n_174;
wire n_400;
wire n_255;
wire n_299;
wire n_243;
wire n_352;
wire n_56;
wire n_293;
wire n_275;
wire n_381;
wire n_227;
wire n_229;
wire n_379;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_360;
wire n_398;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_45;
wire n_268;
wire n_42;
wire n_313;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_416;
wire n_143;
wire n_351;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_406;
wire n_303;
wire n_321;
wire n_100;
wire n_368;
wire n_51;
wire n_205;
wire n_361;
wire n_261;
wire n_86;
wire n_324;
wire n_70;
wire n_32;
wire n_228;
wire n_389;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_394;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_424;
wire n_133;
wire n_257;
wire n_344;
wire n_210;
wire n_206;
wire n_408;
wire n_85;
wire n_96;
wire n_308;
wire n_364;

AOI21xp5_ASAP7_75t_L g18 ( 
.A1(n_0),
.A2(n_19),
.B(n_431),
.Y(n_18)
);

NOR2xp33_ASAP7_75t_L g431 ( 
.A(n_0),
.B(n_432),
.Y(n_431)
);

AND2x2_ASAP7_75t_L g36 ( 
.A(n_1),
.B(n_37),
.Y(n_36)
);

AND2x2_ASAP7_75t_L g92 ( 
.A(n_1),
.B(n_93),
.Y(n_92)
);

AND2x2_ASAP7_75t_L g111 ( 
.A(n_1),
.B(n_112),
.Y(n_111)
);

AND2x2_ASAP7_75t_L g121 ( 
.A(n_1),
.B(n_122),
.Y(n_121)
);

AND2x2_ASAP7_75t_L g133 ( 
.A(n_1),
.B(n_134),
.Y(n_133)
);

AND2x2_ASAP7_75t_L g185 ( 
.A(n_1),
.B(n_186),
.Y(n_185)
);

AND2x2_ASAP7_75t_L g422 ( 
.A(n_1),
.B(n_423),
.Y(n_422)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_2),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g113 ( 
.A(n_2),
.Y(n_113)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_2),
.Y(n_131)
);

BUFx3_ASAP7_75t_L g153 ( 
.A(n_2),
.Y(n_153)
);

BUFx5_ASAP7_75t_L g73 ( 
.A(n_3),
.Y(n_73)
);

BUFx6f_ASAP7_75t_L g81 ( 
.A(n_3),
.Y(n_81)
);

BUFx6f_ASAP7_75t_L g94 ( 
.A(n_3),
.Y(n_94)
);

BUFx6f_ASAP7_75t_L g282 ( 
.A(n_3),
.Y(n_282)
);

AND2x2_ASAP7_75t_SL g55 ( 
.A(n_4),
.B(n_56),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_L g82 ( 
.A(n_4),
.B(n_83),
.Y(n_82)
);

AND2x2_ASAP7_75t_L g108 ( 
.A(n_4),
.B(n_109),
.Y(n_108)
);

AND2x2_ASAP7_75t_SL g154 ( 
.A(n_4),
.B(n_155),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_SL g182 ( 
.A(n_4),
.B(n_183),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_L g279 ( 
.A(n_4),
.B(n_280),
.Y(n_279)
);

NAND2xp5_ASAP7_75t_SL g284 ( 
.A(n_4),
.B(n_285),
.Y(n_284)
);

NAND2xp5_ASAP7_75t_L g307 ( 
.A(n_4),
.B(n_149),
.Y(n_307)
);

AOI22xp5_ASAP7_75t_SL g40 ( 
.A1(n_5),
.A2(n_11),
.B1(n_41),
.B2(n_44),
.Y(n_40)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_5),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_L g136 ( 
.A(n_5),
.B(n_137),
.Y(n_136)
);

AND2x2_ASAP7_75t_SL g152 ( 
.A(n_5),
.B(n_153),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_L g298 ( 
.A(n_5),
.B(n_299),
.Y(n_298)
);

NAND2xp5_ASAP7_75t_L g309 ( 
.A(n_5),
.B(n_310),
.Y(n_309)
);

NAND2xp5_ASAP7_75t_SL g340 ( 
.A(n_5),
.B(n_341),
.Y(n_340)
);

NAND2xp5_ASAP7_75t_SL g88 ( 
.A(n_6),
.B(n_89),
.Y(n_88)
);

AND2x2_ASAP7_75t_L g240 ( 
.A(n_6),
.B(n_241),
.Y(n_240)
);

NAND2xp5_ASAP7_75t_L g251 ( 
.A(n_6),
.B(n_252),
.Y(n_251)
);

NAND2xp5_ASAP7_75t_L g293 ( 
.A(n_6),
.B(n_294),
.Y(n_293)
);

NAND2xp5_ASAP7_75t_L g327 ( 
.A(n_6),
.B(n_303),
.Y(n_327)
);

NAND2xp5_ASAP7_75t_SL g349 ( 
.A(n_6),
.B(n_350),
.Y(n_349)
);

NAND2xp5_ASAP7_75t_SL g354 ( 
.A(n_6),
.B(n_355),
.Y(n_354)
);

INVx1_ASAP7_75t_L g432 ( 
.A(n_7),
.Y(n_432)
);

BUFx5_ASAP7_75t_L g37 ( 
.A(n_8),
.Y(n_37)
);

BUFx5_ASAP7_75t_L g43 ( 
.A(n_8),
.Y(n_43)
);

INVx2_ASAP7_75t_L g150 ( 
.A(n_8),
.Y(n_150)
);

BUFx3_ASAP7_75t_L g265 ( 
.A(n_8),
.Y(n_265)
);

NAND2x1p5_ASAP7_75t_L g68 ( 
.A(n_9),
.B(n_69),
.Y(n_68)
);

AND2x2_ASAP7_75t_L g85 ( 
.A(n_9),
.B(n_86),
.Y(n_85)
);

AND2x2_ASAP7_75t_L g124 ( 
.A(n_9),
.B(n_43),
.Y(n_124)
);

AND2x2_ASAP7_75t_L g128 ( 
.A(n_9),
.B(n_129),
.Y(n_128)
);

AND2x2_ASAP7_75t_L g158 ( 
.A(n_9),
.B(n_73),
.Y(n_158)
);

AND2x2_ASAP7_75t_L g193 ( 
.A(n_9),
.B(n_194),
.Y(n_193)
);

AND2x2_ASAP7_75t_L g198 ( 
.A(n_9),
.B(n_199),
.Y(n_198)
);

AND2x2_ASAP7_75t_L g406 ( 
.A(n_9),
.B(n_29),
.Y(n_406)
);

BUFx6f_ASAP7_75t_L g87 ( 
.A(n_10),
.Y(n_87)
);

BUFx3_ASAP7_75t_L g106 ( 
.A(n_10),
.Y(n_106)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_10),
.Y(n_135)
);

INVx3_ASAP7_75t_L g157 ( 
.A(n_10),
.Y(n_157)
);

INVx2_ASAP7_75t_L g212 ( 
.A(n_10),
.Y(n_212)
);

BUFx3_ASAP7_75t_L g239 ( 
.A(n_10),
.Y(n_239)
);

AND2x2_ASAP7_75t_L g32 ( 
.A(n_11),
.B(n_33),
.Y(n_32)
);

NAND2xp5_ASAP7_75t_L g72 ( 
.A(n_11),
.B(n_73),
.Y(n_72)
);

AND2x2_ASAP7_75t_L g209 ( 
.A(n_11),
.B(n_210),
.Y(n_209)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_11),
.Y(n_262)
);

NAND2xp5_ASAP7_75t_SL g425 ( 
.A(n_11),
.B(n_426),
.Y(n_425)
);

AND2x2_ASAP7_75t_L g51 ( 
.A(n_12),
.B(n_52),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_L g78 ( 
.A(n_12),
.B(n_79),
.Y(n_78)
);

AND2x2_ASAP7_75t_L g103 ( 
.A(n_12),
.B(n_104),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_L g147 ( 
.A(n_12),
.B(n_148),
.Y(n_147)
);

AND2x2_ASAP7_75t_L g207 ( 
.A(n_12),
.B(n_208),
.Y(n_207)
);

INVx1_ASAP7_75t_L g415 ( 
.A(n_12),
.Y(n_415)
);

NAND2xp5_ASAP7_75t_SL g28 ( 
.A(n_13),
.B(n_29),
.Y(n_28)
);

AND2x2_ASAP7_75t_L g60 ( 
.A(n_13),
.B(n_61),
.Y(n_60)
);

AND2x2_ASAP7_75t_L g233 ( 
.A(n_13),
.B(n_234),
.Y(n_233)
);

NAND2xp5_ASAP7_75t_L g248 ( 
.A(n_13),
.B(n_249),
.Y(n_248)
);

NAND2xp5_ASAP7_75t_L g301 ( 
.A(n_13),
.B(n_302),
.Y(n_301)
);

AND2x2_ASAP7_75t_L g328 ( 
.A(n_13),
.B(n_93),
.Y(n_328)
);

NAND2xp5_ASAP7_75t_L g336 ( 
.A(n_13),
.B(n_337),
.Y(n_336)
);

NAND2xp5_ASAP7_75t_SL g359 ( 
.A(n_13),
.B(n_341),
.Y(n_359)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_14),
.Y(n_63)
);

INVx6_ASAP7_75t_L g110 ( 
.A(n_14),
.Y(n_110)
);

BUFx6f_ASAP7_75t_L g196 ( 
.A(n_14),
.Y(n_196)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_15),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g70 ( 
.A(n_15),
.Y(n_70)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_16),
.Y(n_35)
);

BUFx12f_ASAP7_75t_L g54 ( 
.A(n_16),
.Y(n_54)
);

BUFx8_ASAP7_75t_L g29 ( 
.A(n_17),
.Y(n_29)
);

INVx2_ASAP7_75t_L g91 ( 
.A(n_17),
.Y(n_91)
);

XOR2xp5_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_392),
.Y(n_19)
);

OAI21xp5_ASAP7_75t_L g20 ( 
.A1(n_21),
.A2(n_216),
.B(n_389),
.Y(n_20)
);

INVxp67_ASAP7_75t_L g21 ( 
.A(n_22),
.Y(n_21)
);

NAND2xp5_ASAP7_75t_L g22 ( 
.A(n_23),
.B(n_167),
.Y(n_22)
);

NOR2xp33_ASAP7_75t_L g391 ( 
.A(n_23),
.B(n_167),
.Y(n_391)
);

MAJIxp5_ASAP7_75t_L g23 ( 
.A(n_24),
.B(n_100),
.C(n_140),
.Y(n_23)
);

OAI22xp5_ASAP7_75t_SL g384 ( 
.A1(n_24),
.A2(n_25),
.B1(n_101),
.B2(n_385),
.Y(n_384)
);

INVx1_ASAP7_75t_SL g24 ( 
.A(n_25),
.Y(n_24)
);

XNOR2xp5_ASAP7_75t_L g25 ( 
.A(n_26),
.B(n_64),
.Y(n_25)
);

INVxp67_ASAP7_75t_L g169 ( 
.A(n_26),
.Y(n_169)
);

MAJIxp5_ASAP7_75t_L g26 ( 
.A(n_27),
.B(n_39),
.C(n_49),
.Y(n_26)
);

XNOR2xp5_ASAP7_75t_L g378 ( 
.A(n_27),
.B(n_379),
.Y(n_378)
);

XNOR2xp5_ASAP7_75t_L g27 ( 
.A(n_28),
.B(n_30),
.Y(n_27)
);

MAJIxp5_ASAP7_75t_L g75 ( 
.A(n_28),
.B(n_32),
.C(n_36),
.Y(n_75)
);

INVx2_ASAP7_75t_L g118 ( 
.A(n_29),
.Y(n_118)
);

AOI22xp5_ASAP7_75t_L g30 ( 
.A1(n_31),
.A2(n_32),
.B1(n_36),
.B2(n_38),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_32),
.Y(n_31)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_34),
.Y(n_33)
);

INVx2_ASAP7_75t_L g358 ( 
.A(n_34),
.Y(n_358)
);

INVx2_ASAP7_75t_L g34 ( 
.A(n_35),
.Y(n_34)
);

INVx2_ASAP7_75t_L g200 ( 
.A(n_35),
.Y(n_200)
);

INVx1_ASAP7_75t_SL g38 ( 
.A(n_36),
.Y(n_38)
);

AND2x2_ASAP7_75t_L g246 ( 
.A(n_36),
.B(n_198),
.Y(n_246)
);

XNOR2xp5_ASAP7_75t_L g277 ( 
.A(n_38),
.B(n_198),
.Y(n_277)
);

AOI22xp33_ASAP7_75t_SL g379 ( 
.A1(n_39),
.A2(n_40),
.B1(n_49),
.B2(n_50),
.Y(n_379)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_40),
.Y(n_39)
);

AOI21xp5_ASAP7_75t_L g255 ( 
.A1(n_40),
.A2(n_256),
.B(n_261),
.Y(n_255)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_42),
.Y(n_41)
);

INVx3_ASAP7_75t_L g42 ( 
.A(n_43),
.Y(n_42)
);

INVx3_ASAP7_75t_L g44 ( 
.A(n_45),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_46),
.Y(n_45)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_46),
.Y(n_249)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_47),
.Y(n_46)
);

INVx2_ASAP7_75t_L g47 ( 
.A(n_48),
.Y(n_47)
);

BUFx5_ASAP7_75t_L g83 ( 
.A(n_48),
.Y(n_83)
);

BUFx6f_ASAP7_75t_L g243 ( 
.A(n_48),
.Y(n_243)
);

BUFx6f_ASAP7_75t_L g260 ( 
.A(n_48),
.Y(n_260)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_50),
.Y(n_49)
);

MAJIxp5_ASAP7_75t_L g50 ( 
.A(n_51),
.B(n_55),
.C(n_60),
.Y(n_50)
);

XNOR2xp5_ASAP7_75t_L g143 ( 
.A(n_51),
.B(n_60),
.Y(n_143)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_53),
.Y(n_52)
);

INVx3_ASAP7_75t_L g339 ( 
.A(n_53),
.Y(n_339)
);

INVx5_ASAP7_75t_L g53 ( 
.A(n_54),
.Y(n_53)
);

INVx2_ASAP7_75t_SL g123 ( 
.A(n_54),
.Y(n_123)
);

BUFx6f_ASAP7_75t_L g285 ( 
.A(n_54),
.Y(n_285)
);

INVx3_ASAP7_75t_L g311 ( 
.A(n_54),
.Y(n_311)
);

XNOR2xp5_ASAP7_75t_L g142 ( 
.A(n_55),
.B(n_143),
.Y(n_142)
);

HB1xp67_ASAP7_75t_L g56 ( 
.A(n_57),
.Y(n_56)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_58),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_59),
.Y(n_58)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_62),
.Y(n_61)
);

INVx3_ASAP7_75t_L g62 ( 
.A(n_63),
.Y(n_62)
);

INVx4_ASAP7_75t_L g253 ( 
.A(n_63),
.Y(n_253)
);

AOI22xp5_ASAP7_75t_SL g64 ( 
.A1(n_65),
.A2(n_77),
.B1(n_98),
.B2(n_99),
.Y(n_64)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_65),
.Y(n_98)
);

AOI22xp5_ASAP7_75t_SL g65 ( 
.A1(n_66),
.A2(n_67),
.B1(n_75),
.B2(n_76),
.Y(n_65)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_67),
.Y(n_66)
);

AOI22xp5_ASAP7_75t_L g67 ( 
.A1(n_68),
.A2(n_71),
.B1(n_72),
.B2(n_74),
.Y(n_67)
);

INVx2_ASAP7_75t_L g74 ( 
.A(n_68),
.Y(n_74)
);

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_70),
.Y(n_69)
);

INVx4_ASAP7_75t_L g187 ( 
.A(n_70),
.Y(n_187)
);

INVx1_ASAP7_75t_L g418 ( 
.A(n_70),
.Y(n_418)
);

MAJIxp5_ASAP7_75t_L g178 ( 
.A(n_71),
.B(n_74),
.C(n_76),
.Y(n_178)
);

INVx1_ASAP7_75t_SL g71 ( 
.A(n_72),
.Y(n_71)
);

INVx2_ASAP7_75t_L g300 ( 
.A(n_73),
.Y(n_300)
);

INVx2_ASAP7_75t_SL g351 ( 
.A(n_73),
.Y(n_351)
);

INVx1_ASAP7_75t_SL g76 ( 
.A(n_75),
.Y(n_76)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_77),
.Y(n_99)
);

HB1xp67_ASAP7_75t_L g170 ( 
.A(n_77),
.Y(n_170)
);

A2O1A1Ixp33_ASAP7_75t_L g77 ( 
.A1(n_78),
.A2(n_82),
.B(n_84),
.C(n_95),
.Y(n_77)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_78),
.Y(n_96)
);

AOI22xp5_ASAP7_75t_L g166 ( 
.A1(n_78),
.A2(n_82),
.B1(n_96),
.B2(n_97),
.Y(n_166)
);

INVx4_ASAP7_75t_L g79 ( 
.A(n_80),
.Y(n_79)
);

INVx8_ASAP7_75t_L g80 ( 
.A(n_81),
.Y(n_80)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_82),
.Y(n_97)
);

XOR2xp5_ASAP7_75t_L g165 ( 
.A(n_84),
.B(n_166),
.Y(n_165)
);

MAJIxp5_ASAP7_75t_L g84 ( 
.A(n_85),
.B(n_88),
.C(n_92),
.Y(n_84)
);

AOI22xp5_ASAP7_75t_L g267 ( 
.A1(n_85),
.A2(n_92),
.B1(n_268),
.B2(n_269),
.Y(n_267)
);

INVx1_ASAP7_75t_SL g268 ( 
.A(n_85),
.Y(n_268)
);

BUFx6f_ASAP7_75t_L g86 ( 
.A(n_87),
.Y(n_86)
);

XOR2xp5_ASAP7_75t_L g266 ( 
.A(n_88),
.B(n_267),
.Y(n_266)
);

INVx4_ASAP7_75t_L g89 ( 
.A(n_90),
.Y(n_89)
);

INVx8_ASAP7_75t_L g183 ( 
.A(n_90),
.Y(n_183)
);

BUFx6f_ASAP7_75t_L g90 ( 
.A(n_91),
.Y(n_90)
);

XNOR2xp5_ASAP7_75t_L g204 ( 
.A(n_92),
.B(n_205),
.Y(n_204)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_92),
.Y(n_269)
);

BUFx6f_ASAP7_75t_L g93 ( 
.A(n_94),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_L g95 ( 
.A(n_96),
.B(n_97),
.Y(n_95)
);

HB1xp67_ASAP7_75t_L g171 ( 
.A(n_98),
.Y(n_171)
);

HB1xp67_ASAP7_75t_L g100 ( 
.A(n_101),
.Y(n_100)
);

INVx1_ASAP7_75t_L g385 ( 
.A(n_101),
.Y(n_385)
);

XNOR2xp5_ASAP7_75t_L g101 ( 
.A(n_102),
.B(n_114),
.Y(n_101)
);

MAJIxp5_ASAP7_75t_L g175 ( 
.A(n_102),
.B(n_126),
.C(n_138),
.Y(n_175)
);

XNOR2xp5_ASAP7_75t_L g102 ( 
.A(n_103),
.B(n_107),
.Y(n_102)
);

MAJx2_ASAP7_75t_L g188 ( 
.A(n_103),
.B(n_108),
.C(n_111),
.Y(n_188)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_105),
.Y(n_104)
);

INVx2_ASAP7_75t_L g105 ( 
.A(n_106),
.Y(n_105)
);

XNOR2xp5_ASAP7_75t_SL g107 ( 
.A(n_108),
.B(n_111),
.Y(n_107)
);

INVx2_ASAP7_75t_L g109 ( 
.A(n_110),
.Y(n_109)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_110),
.Y(n_137)
);

BUFx6f_ASAP7_75t_L g112 ( 
.A(n_113),
.Y(n_112)
);

BUFx6f_ASAP7_75t_L g208 ( 
.A(n_113),
.Y(n_208)
);

BUFx6f_ASAP7_75t_L g236 ( 
.A(n_113),
.Y(n_236)
);

AOI22xp5_ASAP7_75t_SL g114 ( 
.A1(n_115),
.A2(n_126),
.B1(n_138),
.B2(n_139),
.Y(n_114)
);

INVx2_ASAP7_75t_L g138 ( 
.A(n_115),
.Y(n_138)
);

XNOR2x1_ASAP7_75t_L g115 ( 
.A(n_116),
.B(n_119),
.Y(n_115)
);

MAJIxp5_ASAP7_75t_L g203 ( 
.A(n_116),
.B(n_120),
.C(n_125),
.Y(n_203)
);

NOR2xp33_ASAP7_75t_SL g116 ( 
.A(n_117),
.B(n_118),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_L g237 ( 
.A(n_117),
.B(n_238),
.Y(n_237)
);

NOR2xp33_ASAP7_75t_L g256 ( 
.A(n_117),
.B(n_257),
.Y(n_256)
);

AOI22xp5_ASAP7_75t_SL g119 ( 
.A1(n_120),
.A2(n_121),
.B1(n_124),
.B2(n_125),
.Y(n_119)
);

OAI22xp5_ASAP7_75t_SL g231 ( 
.A1(n_120),
.A2(n_121),
.B1(n_146),
.B2(n_147),
.Y(n_231)
);

INVx2_ASAP7_75t_L g120 ( 
.A(n_121),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_L g145 ( 
.A(n_121),
.B(n_146),
.Y(n_145)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_123),
.Y(n_122)
);

INVx1_ASAP7_75t_SL g125 ( 
.A(n_124),
.Y(n_125)
);

AOI22xp5_ASAP7_75t_L g197 ( 
.A1(n_124),
.A2(n_125),
.B1(n_198),
.B2(n_201),
.Y(n_197)
);

XNOR2xp5_ASAP7_75t_L g313 ( 
.A(n_124),
.B(n_284),
.Y(n_313)
);

NOR2xp33_ASAP7_75t_L g283 ( 
.A(n_125),
.B(n_284),
.Y(n_283)
);

MAJIxp5_ASAP7_75t_L g407 ( 
.A(n_125),
.B(n_193),
.C(n_198),
.Y(n_407)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_126),
.Y(n_139)
);

MAJIxp5_ASAP7_75t_L g126 ( 
.A(n_127),
.B(n_132),
.C(n_136),
.Y(n_126)
);

AOI22xp33_ASAP7_75t_SL g162 ( 
.A1(n_127),
.A2(n_128),
.B1(n_136),
.B2(n_163),
.Y(n_162)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_128),
.Y(n_127)
);

BUFx6f_ASAP7_75t_L g129 ( 
.A(n_130),
.Y(n_129)
);

INVx2_ASAP7_75t_L g130 ( 
.A(n_131),
.Y(n_130)
);

BUFx3_ASAP7_75t_L g297 ( 
.A(n_131),
.Y(n_297)
);

OAI22xp5_ASAP7_75t_SL g160 ( 
.A1(n_132),
.A2(n_133),
.B1(n_161),
.B2(n_162),
.Y(n_160)
);

AOI22xp5_ASAP7_75t_SL g424 ( 
.A1(n_132),
.A2(n_133),
.B1(n_425),
.B2(n_428),
.Y(n_424)
);

INVx1_ASAP7_75t_SL g132 ( 
.A(n_133),
.Y(n_132)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_135),
.Y(n_134)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_136),
.Y(n_163)
);

XNOR2xp5_ASAP7_75t_L g383 ( 
.A(n_140),
.B(n_384),
.Y(n_383)
);

MAJIxp5_ASAP7_75t_L g140 ( 
.A(n_141),
.B(n_159),
.C(n_164),
.Y(n_140)
);

XOR2xp5_ASAP7_75t_L g375 ( 
.A(n_141),
.B(n_376),
.Y(n_375)
);

MAJIxp5_ASAP7_75t_L g141 ( 
.A(n_142),
.B(n_144),
.C(n_151),
.Y(n_141)
);

XNOR2xp5_ASAP7_75t_SL g222 ( 
.A(n_142),
.B(n_223),
.Y(n_222)
);

AOI22xp5_ASAP7_75t_L g223 ( 
.A1(n_144),
.A2(n_145),
.B1(n_151),
.B2(n_224),
.Y(n_223)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_145),
.Y(n_144)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_147),
.Y(n_146)
);

BUFx3_ASAP7_75t_L g148 ( 
.A(n_149),
.Y(n_148)
);

INVx3_ASAP7_75t_L g149 ( 
.A(n_150),
.Y(n_149)
);

INVx2_ASAP7_75t_L g343 ( 
.A(n_150),
.Y(n_343)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_151),
.Y(n_224)
);

MAJx2_ASAP7_75t_L g151 ( 
.A(n_152),
.B(n_154),
.C(n_158),
.Y(n_151)
);

AOI22xp5_ASAP7_75t_L g228 ( 
.A1(n_152),
.A2(n_158),
.B1(n_229),
.B2(n_230),
.Y(n_228)
);

CKINVDCx14_ASAP7_75t_R g229 ( 
.A(n_152),
.Y(n_229)
);

XNOR2xp5_ASAP7_75t_L g227 ( 
.A(n_154),
.B(n_228),
.Y(n_227)
);

BUFx3_ASAP7_75t_L g155 ( 
.A(n_156),
.Y(n_155)
);

INVx2_ASAP7_75t_L g156 ( 
.A(n_157),
.Y(n_156)
);

BUFx3_ASAP7_75t_L g304 ( 
.A(n_157),
.Y(n_304)
);

INVx1_ASAP7_75t_SL g230 ( 
.A(n_158),
.Y(n_230)
);

AOI22xp5_ASAP7_75t_L g413 ( 
.A1(n_158),
.A2(n_198),
.B1(n_201),
.B2(n_230),
.Y(n_413)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_160),
.Y(n_159)
);

XNOR2xp5_ASAP7_75t_L g376 ( 
.A(n_160),
.B(n_165),
.Y(n_376)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_162),
.Y(n_161)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_165),
.Y(n_164)
);

XNOR2xp5_ASAP7_75t_L g167 ( 
.A(n_168),
.B(n_172),
.Y(n_167)
);

INVx1_ASAP7_75t_L g395 ( 
.A(n_168),
.Y(n_395)
);

MAJIxp5_ASAP7_75t_L g168 ( 
.A(n_169),
.B(n_170),
.C(n_171),
.Y(n_168)
);

AOI22xp5_ASAP7_75t_SL g172 ( 
.A1(n_173),
.A2(n_191),
.B1(n_214),
.B2(n_215),
.Y(n_172)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_173),
.Y(n_214)
);

AOI22xp5_ASAP7_75t_L g173 ( 
.A1(n_174),
.A2(n_175),
.B1(n_176),
.B2(n_190),
.Y(n_173)
);

MAJIxp5_ASAP7_75t_L g397 ( 
.A(n_174),
.B(n_177),
.C(n_189),
.Y(n_397)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_175),
.Y(n_174)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_176),
.Y(n_190)
);

AOI22xp5_ASAP7_75t_L g176 ( 
.A1(n_177),
.A2(n_178),
.B1(n_179),
.B2(n_189),
.Y(n_176)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_178),
.Y(n_177)
);

INVx1_ASAP7_75t_SL g189 ( 
.A(n_179),
.Y(n_189)
);

XNOR2xp5_ASAP7_75t_L g179 ( 
.A(n_180),
.B(n_188),
.Y(n_179)
);

OAI22xp5_ASAP7_75t_L g180 ( 
.A1(n_181),
.A2(n_182),
.B1(n_184),
.B2(n_185),
.Y(n_180)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_182),
.Y(n_181)
);

MAJx2_ASAP7_75t_L g403 ( 
.A(n_182),
.B(n_184),
.C(n_188),
.Y(n_403)
);

INVx2_ASAP7_75t_SL g184 ( 
.A(n_185),
.Y(n_184)
);

XNOR2xp5_ASAP7_75t_L g405 ( 
.A(n_185),
.B(n_406),
.Y(n_405)
);

INVx6_ASAP7_75t_L g186 ( 
.A(n_187),
.Y(n_186)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_191),
.Y(n_215)
);

MAJIxp5_ASAP7_75t_L g394 ( 
.A(n_191),
.B(n_214),
.C(n_395),
.Y(n_394)
);

XNOR2xp5_ASAP7_75t_L g191 ( 
.A(n_192),
.B(n_202),
.Y(n_191)
);

MAJIxp5_ASAP7_75t_L g401 ( 
.A(n_192),
.B(n_203),
.C(n_204),
.Y(n_401)
);

XNOR2xp5_ASAP7_75t_L g192 ( 
.A(n_193),
.B(n_197),
.Y(n_192)
);

INVx4_ASAP7_75t_L g194 ( 
.A(n_195),
.Y(n_194)
);

INVx6_ASAP7_75t_L g195 ( 
.A(n_196),
.Y(n_195)
);

HB1xp67_ASAP7_75t_L g423 ( 
.A(n_196),
.Y(n_423)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_198),
.Y(n_201)
);

INVx5_ASAP7_75t_L g199 ( 
.A(n_200),
.Y(n_199)
);

XNOR2xp5_ASAP7_75t_L g202 ( 
.A(n_203),
.B(n_204),
.Y(n_202)
);

AOI22xp5_ASAP7_75t_L g205 ( 
.A1(n_206),
.A2(n_207),
.B1(n_209),
.B2(n_213),
.Y(n_205)
);

MAJIxp5_ASAP7_75t_L g420 ( 
.A(n_206),
.B(n_213),
.C(n_269),
.Y(n_420)
);

CKINVDCx16_ASAP7_75t_R g206 ( 
.A(n_207),
.Y(n_206)
);

INVx5_ASAP7_75t_L g427 ( 
.A(n_208),
.Y(n_427)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_209),
.Y(n_213)
);

INVx6_ASAP7_75t_L g210 ( 
.A(n_211),
.Y(n_210)
);

BUFx6f_ASAP7_75t_L g211 ( 
.A(n_212),
.Y(n_211)
);

AOI21xp5_ASAP7_75t_R g216 ( 
.A1(n_217),
.A2(n_371),
.B(n_386),
.Y(n_216)
);

OAI21x1_ASAP7_75t_SL g217 ( 
.A1(n_218),
.A2(n_286),
.B(n_370),
.Y(n_217)
);

NOR2xp67_ASAP7_75t_SL g218 ( 
.A(n_219),
.B(n_270),
.Y(n_218)
);

NAND2xp5_ASAP7_75t_SL g370 ( 
.A(n_219),
.B(n_270),
.Y(n_370)
);

XOR2xp5_ASAP7_75t_L g219 ( 
.A(n_220),
.B(n_244),
.Y(n_219)
);

AOI22xp5_ASAP7_75t_L g220 ( 
.A1(n_221),
.A2(n_222),
.B1(n_225),
.B2(n_226),
.Y(n_220)
);

MAJIxp5_ASAP7_75t_L g373 ( 
.A(n_221),
.B(n_226),
.C(n_244),
.Y(n_373)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_222),
.Y(n_221)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_226),
.Y(n_225)
);

MAJIxp5_ASAP7_75t_L g226 ( 
.A(n_227),
.B(n_231),
.C(n_232),
.Y(n_226)
);

XNOR2xp5_ASAP7_75t_L g272 ( 
.A(n_227),
.B(n_273),
.Y(n_272)
);

XNOR2xp5_ASAP7_75t_L g273 ( 
.A(n_231),
.B(n_232),
.Y(n_273)
);

MAJx2_ASAP7_75t_L g232 ( 
.A(n_233),
.B(n_237),
.C(n_240),
.Y(n_232)
);

XNOR2xp5_ASAP7_75t_L g318 ( 
.A(n_233),
.B(n_240),
.Y(n_318)
);

INVx3_ASAP7_75t_L g234 ( 
.A(n_235),
.Y(n_234)
);

INVx2_ASAP7_75t_L g235 ( 
.A(n_236),
.Y(n_235)
);

XNOR2xp5_ASAP7_75t_L g317 ( 
.A(n_237),
.B(n_318),
.Y(n_317)
);

INVx5_ASAP7_75t_L g238 ( 
.A(n_239),
.Y(n_238)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_242),
.Y(n_241)
);

INVx2_ASAP7_75t_L g242 ( 
.A(n_243),
.Y(n_242)
);

XNOR2xp5_ASAP7_75t_SL g244 ( 
.A(n_245),
.B(n_254),
.Y(n_244)
);

MAJIxp5_ASAP7_75t_L g380 ( 
.A(n_245),
.B(n_255),
.C(n_266),
.Y(n_380)
);

MAJIxp5_ASAP7_75t_L g245 ( 
.A(n_246),
.B(n_247),
.C(n_250),
.Y(n_245)
);

XOR2xp5_ASAP7_75t_L g274 ( 
.A(n_246),
.B(n_275),
.Y(n_274)
);

AOI22xp5_ASAP7_75t_L g275 ( 
.A1(n_247),
.A2(n_248),
.B1(n_250),
.B2(n_251),
.Y(n_275)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_248),
.Y(n_247)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_251),
.Y(n_250)
);

INVx4_ASAP7_75t_L g252 ( 
.A(n_253),
.Y(n_252)
);

XNOR2xp5_ASAP7_75t_L g254 ( 
.A(n_255),
.B(n_266),
.Y(n_254)
);

INVx2_ASAP7_75t_L g257 ( 
.A(n_258),
.Y(n_257)
);

BUFx3_ASAP7_75t_L g258 ( 
.A(n_259),
.Y(n_258)
);

BUFx6f_ASAP7_75t_L g259 ( 
.A(n_260),
.Y(n_259)
);

NOR2xp33_ASAP7_75t_L g261 ( 
.A(n_262),
.B(n_263),
.Y(n_261)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_264),
.Y(n_263)
);

BUFx3_ASAP7_75t_L g264 ( 
.A(n_265),
.Y(n_264)
);

MAJIxp5_ASAP7_75t_L g270 ( 
.A(n_271),
.B(n_274),
.C(n_276),
.Y(n_270)
);

AOI22xp5_ASAP7_75t_SL g366 ( 
.A1(n_271),
.A2(n_272),
.B1(n_367),
.B2(n_368),
.Y(n_366)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_272),
.Y(n_271)
);

XNOR2xp5_ASAP7_75t_SL g368 ( 
.A(n_274),
.B(n_276),
.Y(n_368)
);

MAJIxp5_ASAP7_75t_L g276 ( 
.A(n_277),
.B(n_278),
.C(n_283),
.Y(n_276)
);

AOI22xp5_ASAP7_75t_L g320 ( 
.A1(n_277),
.A2(n_278),
.B1(n_279),
.B2(n_321),
.Y(n_320)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_277),
.Y(n_321)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_279),
.Y(n_278)
);

INVx4_ASAP7_75t_L g280 ( 
.A(n_281),
.Y(n_280)
);

INVx6_ASAP7_75t_L g281 ( 
.A(n_282),
.Y(n_281)
);

XNOR2xp5_ASAP7_75t_SL g319 ( 
.A(n_283),
.B(n_320),
.Y(n_319)
);

AOI21x1_ASAP7_75t_SL g286 ( 
.A1(n_287),
.A2(n_364),
.B(n_369),
.Y(n_286)
);

OAI21xp5_ASAP7_75t_L g287 ( 
.A1(n_288),
.A2(n_322),
.B(n_363),
.Y(n_287)
);

NOR2xp33_ASAP7_75t_L g288 ( 
.A(n_289),
.B(n_314),
.Y(n_288)
);

NAND2xp5_ASAP7_75t_SL g363 ( 
.A(n_289),
.B(n_314),
.Y(n_363)
);

MAJIxp5_ASAP7_75t_L g289 ( 
.A(n_290),
.B(n_305),
.C(n_312),
.Y(n_289)
);

AOI22xp33_ASAP7_75t_SL g329 ( 
.A1(n_290),
.A2(n_291),
.B1(n_330),
.B2(n_332),
.Y(n_329)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_291),
.Y(n_290)
);

XOR2xp5_ASAP7_75t_L g291 ( 
.A(n_292),
.B(n_301),
.Y(n_291)
);

XNOR2xp5_ASAP7_75t_L g292 ( 
.A(n_293),
.B(n_298),
.Y(n_292)
);

MAJIxp5_ASAP7_75t_L g316 ( 
.A(n_293),
.B(n_298),
.C(n_301),
.Y(n_316)
);

INVx2_ASAP7_75t_L g294 ( 
.A(n_295),
.Y(n_294)
);

INVx2_ASAP7_75t_L g295 ( 
.A(n_296),
.Y(n_295)
);

INVx2_ASAP7_75t_L g296 ( 
.A(n_297),
.Y(n_296)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_300),
.Y(n_299)
);

BUFx3_ASAP7_75t_L g302 ( 
.A(n_303),
.Y(n_302)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_304),
.Y(n_303)
);

AOI22xp5_ASAP7_75t_L g330 ( 
.A1(n_305),
.A2(n_312),
.B1(n_313),
.B2(n_331),
.Y(n_330)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_305),
.Y(n_331)
);

NAND2xp5_ASAP7_75t_L g305 ( 
.A(n_306),
.B(n_308),
.Y(n_305)
);

OAI22xp5_ASAP7_75t_SL g325 ( 
.A1(n_306),
.A2(n_307),
.B1(n_308),
.B2(n_309),
.Y(n_325)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_307),
.Y(n_306)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_309),
.Y(n_308)
);

INVx4_ASAP7_75t_L g310 ( 
.A(n_311),
.Y(n_310)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_313),
.Y(n_312)
);

XNOR2xp5_ASAP7_75t_L g314 ( 
.A(n_315),
.B(n_319),
.Y(n_314)
);

XNOR2xp5_ASAP7_75t_L g315 ( 
.A(n_316),
.B(n_317),
.Y(n_315)
);

MAJIxp5_ASAP7_75t_L g365 ( 
.A(n_316),
.B(n_317),
.C(n_319),
.Y(n_365)
);

AOI21xp5_ASAP7_75t_L g322 ( 
.A1(n_323),
.A2(n_333),
.B(n_362),
.Y(n_322)
);

NAND2xp5_ASAP7_75t_L g323 ( 
.A(n_324),
.B(n_329),
.Y(n_323)
);

NOR2xp33_ASAP7_75t_SL g362 ( 
.A(n_324),
.B(n_329),
.Y(n_362)
);

MAJIxp5_ASAP7_75t_L g324 ( 
.A(n_325),
.B(n_326),
.C(n_328),
.Y(n_324)
);

XOR2xp5_ASAP7_75t_L g344 ( 
.A(n_325),
.B(n_345),
.Y(n_344)
);

OAI22xp5_ASAP7_75t_SL g345 ( 
.A1(n_326),
.A2(n_327),
.B1(n_328),
.B2(n_346),
.Y(n_345)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_327),
.Y(n_326)
);

CKINVDCx16_ASAP7_75t_R g346 ( 
.A(n_328),
.Y(n_346)
);

INVxp67_ASAP7_75t_SL g332 ( 
.A(n_330),
.Y(n_332)
);

OAI21xp5_ASAP7_75t_SL g333 ( 
.A1(n_334),
.A2(n_347),
.B(n_361),
.Y(n_333)
);

NOR2xp33_ASAP7_75t_L g334 ( 
.A(n_335),
.B(n_344),
.Y(n_334)
);

NAND2xp5_ASAP7_75t_SL g361 ( 
.A(n_335),
.B(n_344),
.Y(n_361)
);

NOR2xp33_ASAP7_75t_L g335 ( 
.A(n_336),
.B(n_340),
.Y(n_335)
);

XNOR2xp5_ASAP7_75t_L g352 ( 
.A(n_336),
.B(n_340),
.Y(n_352)
);

INVx2_ASAP7_75t_L g337 ( 
.A(n_338),
.Y(n_337)
);

INVx1_ASAP7_75t_L g338 ( 
.A(n_339),
.Y(n_338)
);

INVx2_ASAP7_75t_L g341 ( 
.A(n_342),
.Y(n_341)
);

INVx1_ASAP7_75t_L g342 ( 
.A(n_343),
.Y(n_342)
);

AOI21xp5_ASAP7_75t_L g347 ( 
.A1(n_348),
.A2(n_353),
.B(n_360),
.Y(n_347)
);

NAND2xp5_ASAP7_75t_L g348 ( 
.A(n_349),
.B(n_352),
.Y(n_348)
);

NOR2xp33_ASAP7_75t_SL g360 ( 
.A(n_349),
.B(n_352),
.Y(n_360)
);

INVx1_ASAP7_75t_L g350 ( 
.A(n_351),
.Y(n_350)
);

NOR2xp33_ASAP7_75t_L g353 ( 
.A(n_354),
.B(n_359),
.Y(n_353)
);

INVx2_ASAP7_75t_L g355 ( 
.A(n_356),
.Y(n_355)
);

BUFx2_ASAP7_75t_L g356 ( 
.A(n_357),
.Y(n_356)
);

INVx1_ASAP7_75t_L g357 ( 
.A(n_358),
.Y(n_357)
);

NAND2xp5_ASAP7_75t_L g364 ( 
.A(n_365),
.B(n_366),
.Y(n_364)
);

NOR2xp33_ASAP7_75t_SL g369 ( 
.A(n_365),
.B(n_366),
.Y(n_369)
);

INVx1_ASAP7_75t_L g367 ( 
.A(n_368),
.Y(n_367)
);

NOR2x1_ASAP7_75t_L g371 ( 
.A(n_372),
.B(n_381),
.Y(n_371)
);

NOR2xp33_ASAP7_75t_L g372 ( 
.A(n_373),
.B(n_374),
.Y(n_372)
);

NAND2xp5_ASAP7_75t_L g387 ( 
.A(n_373),
.B(n_374),
.Y(n_387)
);

XNOR2xp5_ASAP7_75t_L g374 ( 
.A(n_375),
.B(n_377),
.Y(n_374)
);

MAJIxp5_ASAP7_75t_L g382 ( 
.A(n_375),
.B(n_378),
.C(n_380),
.Y(n_382)
);

XNOR2xp5_ASAP7_75t_L g377 ( 
.A(n_378),
.B(n_380),
.Y(n_377)
);

OAI21x1_ASAP7_75t_L g386 ( 
.A1(n_381),
.A2(n_387),
.B(n_388),
.Y(n_386)
);

AND2x2_ASAP7_75t_L g381 ( 
.A(n_382),
.B(n_383),
.Y(n_381)
);

OR2x2_ASAP7_75t_L g388 ( 
.A(n_382),
.B(n_383),
.Y(n_388)
);

INVx1_ASAP7_75t_L g389 ( 
.A(n_390),
.Y(n_389)
);

HB1xp67_ASAP7_75t_L g390 ( 
.A(n_391),
.Y(n_390)
);

NOR2xp33_ASAP7_75t_L g392 ( 
.A(n_393),
.B(n_429),
.Y(n_392)
);

NOR2xp33_ASAP7_75t_L g393 ( 
.A(n_394),
.B(n_396),
.Y(n_393)
);

NAND2xp5_ASAP7_75t_L g430 ( 
.A(n_394),
.B(n_396),
.Y(n_430)
);

XNOR2xp5_ASAP7_75t_L g396 ( 
.A(n_397),
.B(n_398),
.Y(n_396)
);

XNOR2xp5_ASAP7_75t_L g398 ( 
.A(n_399),
.B(n_411),
.Y(n_398)
);

AOI22xp5_ASAP7_75t_L g399 ( 
.A1(n_400),
.A2(n_401),
.B1(n_402),
.B2(n_410),
.Y(n_399)
);

INVx1_ASAP7_75t_SL g400 ( 
.A(n_401),
.Y(n_400)
);

INVx1_ASAP7_75t_L g410 ( 
.A(n_402),
.Y(n_410)
);

XNOR2xp5_ASAP7_75t_SL g402 ( 
.A(n_403),
.B(n_404),
.Y(n_402)
);

AO22x1_ASAP7_75t_SL g404 ( 
.A1(n_405),
.A2(n_407),
.B1(n_408),
.B2(n_409),
.Y(n_404)
);

INVx1_ASAP7_75t_L g408 ( 
.A(n_405),
.Y(n_408)
);

INVx1_ASAP7_75t_SL g409 ( 
.A(n_407),
.Y(n_409)
);

XOR2xp5_ASAP7_75t_L g411 ( 
.A(n_412),
.B(n_419),
.Y(n_411)
);

XNOR2xp5_ASAP7_75t_SL g412 ( 
.A(n_413),
.B(n_414),
.Y(n_412)
);

NOR2xp33_ASAP7_75t_L g414 ( 
.A(n_415),
.B(n_416),
.Y(n_414)
);

INVx2_ASAP7_75t_L g416 ( 
.A(n_417),
.Y(n_416)
);

INVx2_ASAP7_75t_SL g417 ( 
.A(n_418),
.Y(n_417)
);

XNOR2xp5_ASAP7_75t_L g419 ( 
.A(n_420),
.B(n_421),
.Y(n_419)
);

XNOR2xp5_ASAP7_75t_L g421 ( 
.A(n_422),
.B(n_424),
.Y(n_421)
);

INVx1_ASAP7_75t_L g428 ( 
.A(n_425),
.Y(n_428)
);

INVx5_ASAP7_75t_L g426 ( 
.A(n_427),
.Y(n_426)
);

INVxp33_ASAP7_75t_L g429 ( 
.A(n_430),
.Y(n_429)
);


endmodule