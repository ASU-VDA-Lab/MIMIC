module fake_netlist_5_943_n_853 (n_137, n_91, n_82, n_122, n_142, n_10, n_140, n_24, n_124, n_86, n_136, n_146, n_143, n_83, n_132, n_61, n_90, n_127, n_75, n_101, n_65, n_78, n_74, n_144, n_114, n_57, n_96, n_37, n_111, n_108, n_129, n_31, n_13, n_66, n_98, n_60, n_155, n_152, n_16, n_43, n_107, n_0, n_58, n_9, n_69, n_18, n_116, n_42, n_22, n_1, n_45, n_117, n_46, n_21, n_94, n_113, n_38, n_123, n_139, n_105, n_80, n_4, n_125, n_35, n_128, n_73, n_17, n_92, n_19, n_149, n_120, n_135, n_30, n_5, n_33, n_126, n_14, n_84, n_23, n_130, n_29, n_79, n_131, n_151, n_47, n_25, n_53, n_8, n_44, n_40, n_34, n_100, n_62, n_138, n_148, n_71, n_154, n_109, n_112, n_85, n_95, n_119, n_59, n_26, n_133, n_55, n_99, n_2, n_3, n_49, n_20, n_6, n_39, n_54, n_147, n_12, n_67, n_121, n_36, n_76, n_87, n_150, n_27, n_64, n_77, n_102, n_106, n_81, n_118, n_28, n_89, n_70, n_115, n_68, n_93, n_72, n_134, n_32, n_41, n_104, n_103, n_56, n_51, n_63, n_97, n_141, n_11, n_153, n_7, n_15, n_145, n_48, n_50, n_52, n_88, n_110, n_853);

input n_137;
input n_91;
input n_82;
input n_122;
input n_142;
input n_10;
input n_140;
input n_24;
input n_124;
input n_86;
input n_136;
input n_146;
input n_143;
input n_83;
input n_132;
input n_61;
input n_90;
input n_127;
input n_75;
input n_101;
input n_65;
input n_78;
input n_74;
input n_144;
input n_114;
input n_57;
input n_96;
input n_37;
input n_111;
input n_108;
input n_129;
input n_31;
input n_13;
input n_66;
input n_98;
input n_60;
input n_155;
input n_152;
input n_16;
input n_43;
input n_107;
input n_0;
input n_58;
input n_9;
input n_69;
input n_18;
input n_116;
input n_42;
input n_22;
input n_1;
input n_45;
input n_117;
input n_46;
input n_21;
input n_94;
input n_113;
input n_38;
input n_123;
input n_139;
input n_105;
input n_80;
input n_4;
input n_125;
input n_35;
input n_128;
input n_73;
input n_17;
input n_92;
input n_19;
input n_149;
input n_120;
input n_135;
input n_30;
input n_5;
input n_33;
input n_126;
input n_14;
input n_84;
input n_23;
input n_130;
input n_29;
input n_79;
input n_131;
input n_151;
input n_47;
input n_25;
input n_53;
input n_8;
input n_44;
input n_40;
input n_34;
input n_100;
input n_62;
input n_138;
input n_148;
input n_71;
input n_154;
input n_109;
input n_112;
input n_85;
input n_95;
input n_119;
input n_59;
input n_26;
input n_133;
input n_55;
input n_99;
input n_2;
input n_3;
input n_49;
input n_20;
input n_6;
input n_39;
input n_54;
input n_147;
input n_12;
input n_67;
input n_121;
input n_36;
input n_76;
input n_87;
input n_150;
input n_27;
input n_64;
input n_77;
input n_102;
input n_106;
input n_81;
input n_118;
input n_28;
input n_89;
input n_70;
input n_115;
input n_68;
input n_93;
input n_72;
input n_134;
input n_32;
input n_41;
input n_104;
input n_103;
input n_56;
input n_51;
input n_63;
input n_97;
input n_141;
input n_11;
input n_153;
input n_7;
input n_15;
input n_145;
input n_48;
input n_50;
input n_52;
input n_88;
input n_110;

output n_853;

wire n_676;
wire n_294;
wire n_431;
wire n_318;
wire n_380;
wire n_419;
wire n_653;
wire n_611;
wire n_444;
wire n_642;
wire n_469;
wire n_615;
wire n_851;
wire n_194;
wire n_316;
wire n_785;
wire n_389;
wire n_843;
wire n_549;
wire n_684;
wire n_850;
wire n_418;
wire n_248;
wire n_315;
wire n_268;
wire n_523;
wire n_451;
wire n_532;
wire n_705;
wire n_619;
wire n_408;
wire n_678;
wire n_664;
wire n_376;
wire n_697;
wire n_503;
wire n_235;
wire n_226;
wire n_605;
wire n_776;
wire n_667;
wire n_515;
wire n_790;
wire n_353;
wire n_351;
wire n_367;
wire n_620;
wire n_643;
wire n_452;
wire n_397;
wire n_493;
wire n_525;
wire n_703;
wire n_698;
wire n_483;
wire n_544;
wire n_683;
wire n_780;
wire n_649;
wire n_552;
wire n_547;
wire n_721;
wire n_841;
wire n_467;
wire n_564;
wire n_802;
wire n_423;
wire n_840;
wire n_284;
wire n_501;
wire n_245;
wire n_823;
wire n_725;
wire n_280;
wire n_744;
wire n_590;
wire n_629;
wire n_672;
wire n_378;
wire n_551;
wire n_762;
wire n_581;
wire n_688;
wire n_382;
wire n_554;
wire n_800;
wire n_254;
wire n_690;
wire n_583;
wire n_671;
wire n_718;
wire n_819;
wire n_302;
wire n_265;
wire n_526;
wire n_719;
wire n_372;
wire n_293;
wire n_443;
wire n_244;
wire n_677;
wire n_173;
wire n_821;
wire n_198;
wire n_714;
wire n_447;
wire n_247;
wire n_314;
wire n_368;
wire n_433;
wire n_604;
wire n_321;
wire n_292;
wire n_625;
wire n_753;
wire n_621;
wire n_455;
wire n_674;
wire n_417;
wire n_612;
wire n_212;
wire n_385;
wire n_516;
wire n_498;
wire n_788;
wire n_507;
wire n_497;
wire n_689;
wire n_738;
wire n_606;
wire n_559;
wire n_275;
wire n_640;
wire n_252;
wire n_624;
wire n_825;
wire n_295;
wire n_330;
wire n_508;
wire n_739;
wire n_506;
wire n_737;
wire n_610;
wire n_692;
wire n_755;
wire n_509;
wire n_568;
wire n_373;
wire n_820;
wire n_757;
wire n_307;
wire n_633;
wire n_439;
wire n_530;
wire n_556;
wire n_209;
wire n_259;
wire n_448;
wire n_758;
wire n_668;
wire n_733;
wire n_375;
wire n_301;
wire n_828;
wire n_779;
wire n_576;
wire n_804;
wire n_186;
wire n_537;
wire n_191;
wire n_587;
wire n_659;
wire n_492;
wire n_792;
wire n_563;
wire n_171;
wire n_756;
wire n_524;
wire n_399;
wire n_341;
wire n_204;
wire n_394;
wire n_250;
wire n_579;
wire n_741;
wire n_548;
wire n_543;
wire n_260;
wire n_812;
wire n_842;
wire n_298;
wire n_650;
wire n_320;
wire n_694;
wire n_518;
wire n_505;
wire n_286;
wire n_282;
wire n_752;
wire n_331;
wire n_406;
wire n_519;
wire n_470;
wire n_782;
wire n_325;
wire n_449;
wire n_724;
wire n_546;
wire n_760;
wire n_658;
wire n_281;
wire n_240;
wire n_381;
wire n_189;
wire n_220;
wire n_291;
wire n_231;
wire n_257;
wire n_390;
wire n_731;
wire n_456;
wire n_371;
wire n_481;
wire n_535;
wire n_709;
wire n_540;
wire n_317;
wire n_618;
wire n_323;
wire n_569;
wire n_769;
wire n_195;
wire n_356;
wire n_227;
wire n_592;
wire n_271;
wire n_831;
wire n_826;
wire n_335;
wire n_654;
wire n_370;
wire n_167;
wire n_234;
wire n_343;
wire n_379;
wire n_308;
wire n_428;
wire n_267;
wire n_514;
wire n_457;
wire n_570;
wire n_833;
wire n_297;
wire n_156;
wire n_603;
wire n_225;
wire n_377;
wire n_751;
wire n_484;
wire n_775;
wire n_219;
wire n_442;
wire n_157;
wire n_814;
wire n_192;
wire n_636;
wire n_786;
wire n_600;
wire n_660;
wire n_223;
wire n_392;
wire n_158;
wire n_655;
wire n_704;
wire n_787;
wire n_264;
wire n_669;
wire n_472;
wire n_742;
wire n_750;
wire n_454;
wire n_387;
wire n_771;
wire n_374;
wire n_163;
wire n_276;
wire n_339;
wire n_183;
wire n_243;
wire n_185;
wire n_398;
wire n_396;
wire n_635;
wire n_347;
wire n_763;
wire n_169;
wire n_550;
wire n_522;
wire n_696;
wire n_255;
wire n_215;
wire n_350;
wire n_196;
wire n_798;
wire n_662;
wire n_459;
wire n_646;
wire n_211;
wire n_218;
wire n_400;
wire n_181;
wire n_436;
wire n_290;
wire n_580;
wire n_221;
wire n_178;
wire n_622;
wire n_723;
wire n_386;
wire n_578;
wire n_287;
wire n_344;
wire n_848;
wire n_555;
wire n_783;
wire n_473;
wire n_422;
wire n_475;
wire n_777;
wire n_661;
wire n_682;
wire n_415;
wire n_485;
wire n_496;
wire n_355;
wire n_849;
wire n_486;
wire n_670;
wire n_816;
wire n_336;
wire n_681;
wire n_584;
wire n_591;
wire n_521;
wire n_614;
wire n_663;
wire n_845;
wire n_430;
wire n_337;
wire n_313;
wire n_631;
wire n_673;
wire n_837;
wire n_479;
wire n_528;
wire n_510;
wire n_216;
wire n_680;
wire n_168;
wire n_395;
wire n_164;
wire n_432;
wire n_553;
wire n_727;
wire n_839;
wire n_311;
wire n_813;
wire n_830;
wire n_773;
wire n_208;
wire n_743;
wire n_214;
wire n_328;
wire n_801;
wire n_299;
wire n_303;
wire n_369;
wire n_675;
wire n_296;
wire n_613;
wire n_241;
wire n_637;
wire n_357;
wire n_598;
wire n_685;
wire n_608;
wire n_184;
wire n_446;
wire n_445;
wire n_829;
wire n_749;
wire n_772;
wire n_691;
wire n_717;
wire n_165;
wire n_468;
wire n_499;
wire n_213;
wire n_342;
wire n_482;
wire n_517;
wire n_588;
wire n_361;
wire n_464;
wire n_789;
wire n_363;
wire n_413;
wire n_402;
wire n_734;
wire n_638;
wire n_700;
wire n_197;
wire n_796;
wire n_573;
wire n_236;
wire n_388;
wire n_761;
wire n_249;
wire n_740;
wire n_304;
wire n_329;
wire n_203;
wire n_274;
wire n_577;
wire n_384;
wire n_582;
wire n_460;
wire n_277;
wire n_477;
wire n_338;
wire n_571;
wire n_461;
wire n_333;
wire n_693;
wire n_309;
wire n_512;
wire n_836;
wire n_462;
wire n_322;
wire n_567;
wire n_258;
wire n_652;
wire n_778;
wire n_306;
wire n_722;
wire n_458;
wire n_288;
wire n_770;
wire n_188;
wire n_190;
wire n_844;
wire n_201;
wire n_263;
wire n_471;
wire n_609;
wire n_852;
wire n_224;
wire n_228;
wire n_283;
wire n_383;
wire n_711;
wire n_781;
wire n_834;
wire n_474;
wire n_765;
wire n_542;
wire n_488;
wire n_463;
wire n_595;
wire n_736;
wire n_502;
wire n_239;
wire n_466;
wire n_420;
wire n_630;
wire n_489;
wire n_632;
wire n_699;
wire n_617;
wire n_310;
wire n_593;
wire n_504;
wire n_511;
wire n_748;
wire n_586;
wire n_846;
wire n_465;
wire n_838;
wire n_358;
wire n_362;
wire n_170;
wire n_332;
wire n_161;
wire n_273;
wire n_585;
wire n_349;
wire n_270;
wire n_616;
wire n_230;
wire n_601;
wire n_279;
wire n_253;
wire n_261;
wire n_174;
wire n_289;
wire n_745;
wire n_627;
wire n_767;
wire n_172;
wire n_206;
wire n_217;
wire n_440;
wire n_726;
wire n_478;
wire n_793;
wire n_545;
wire n_441;
wire n_450;
wire n_648;
wire n_312;
wire n_476;
wire n_818;
wire n_429;
wire n_534;
wire n_345;
wire n_210;
wire n_494;
wire n_641;
wire n_628;
wire n_365;
wire n_774;
wire n_729;
wire n_730;
wire n_176;
wire n_557;
wire n_182;
wire n_354;
wire n_575;
wire n_607;
wire n_480;
wire n_647;
wire n_237;
wire n_425;
wire n_513;
wire n_407;
wire n_527;
wire n_710;
wire n_707;
wire n_795;
wire n_832;
wire n_695;
wire n_180;
wire n_560;
wire n_656;
wire n_340;
wire n_207;
wire n_561;
wire n_346;
wire n_393;
wire n_229;
wire n_495;
wire n_487;
wire n_602;
wire n_665;
wire n_574;
wire n_437;
wire n_177;
wire n_403;
wire n_453;
wire n_421;
wire n_720;
wire n_623;
wire n_405;
wire n_824;
wire n_359;
wire n_490;
wire n_805;
wire n_326;
wire n_794;
wire n_768;
wire n_233;
wire n_404;
wire n_686;
wire n_205;
wire n_366;
wire n_572;
wire n_712;
wire n_754;
wire n_847;
wire n_815;
wire n_246;
wire n_596;
wire n_179;
wire n_410;
wire n_558;
wire n_708;
wire n_269;
wire n_529;
wire n_735;
wire n_702;
wire n_285;
wire n_822;
wire n_412;
wire n_232;
wire n_679;
wire n_327;
wire n_657;
wire n_644;
wire n_728;
wire n_202;
wire n_266;
wire n_272;
wire n_491;
wire n_427;
wire n_791;
wire n_732;
wire n_193;
wire n_251;
wire n_352;
wire n_160;
wire n_566;
wire n_565;
wire n_426;
wire n_520;
wire n_808;
wire n_409;
wire n_797;
wire n_589;
wire n_716;
wire n_597;
wire n_500;
wire n_562;
wire n_300;
wire n_651;
wire n_435;
wire n_809;
wire n_159;
wire n_334;
wire n_599;
wire n_766;
wire n_811;
wire n_541;
wire n_807;
wire n_391;
wire n_701;
wire n_434;
wire n_645;
wire n_539;
wire n_835;
wire n_175;
wire n_538;
wire n_666;
wire n_262;
wire n_803;
wire n_238;
wire n_639;
wire n_799;
wire n_687;
wire n_715;
wire n_411;
wire n_414;
wire n_319;
wire n_364;
wire n_536;
wire n_531;
wire n_242;
wire n_817;
wire n_360;
wire n_594;
wire n_764;
wire n_200;
wire n_162;
wire n_759;
wire n_222;
wire n_438;
wire n_806;
wire n_713;
wire n_324;
wire n_810;
wire n_634;
wire n_416;
wire n_199;
wire n_827;
wire n_187;
wire n_401;
wire n_348;
wire n_166;
wire n_626;
wire n_424;
wire n_706;
wire n_746;
wire n_256;
wire n_305;
wire n_533;
wire n_747;
wire n_278;
wire n_784;

CKINVDCx20_ASAP7_75t_R g156 ( 
.A(n_115),
.Y(n_156)
);

CKINVDCx5p33_ASAP7_75t_R g157 ( 
.A(n_4),
.Y(n_157)
);

CKINVDCx5p33_ASAP7_75t_R g158 ( 
.A(n_100),
.Y(n_158)
);

CKINVDCx5p33_ASAP7_75t_R g159 ( 
.A(n_9),
.Y(n_159)
);

BUFx6f_ASAP7_75t_L g160 ( 
.A(n_12),
.Y(n_160)
);

CKINVDCx5p33_ASAP7_75t_R g161 ( 
.A(n_68),
.Y(n_161)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_94),
.Y(n_162)
);

CKINVDCx5p33_ASAP7_75t_R g163 ( 
.A(n_40),
.Y(n_163)
);

CKINVDCx5p33_ASAP7_75t_R g164 ( 
.A(n_126),
.Y(n_164)
);

CKINVDCx5p33_ASAP7_75t_R g165 ( 
.A(n_18),
.Y(n_165)
);

CKINVDCx5p33_ASAP7_75t_R g166 ( 
.A(n_143),
.Y(n_166)
);

CKINVDCx5p33_ASAP7_75t_R g167 ( 
.A(n_75),
.Y(n_167)
);

BUFx10_ASAP7_75t_L g168 ( 
.A(n_107),
.Y(n_168)
);

CKINVDCx5p33_ASAP7_75t_R g169 ( 
.A(n_24),
.Y(n_169)
);

BUFx3_ASAP7_75t_L g170 ( 
.A(n_117),
.Y(n_170)
);

INVx2_ASAP7_75t_L g171 ( 
.A(n_137),
.Y(n_171)
);

CKINVDCx5p33_ASAP7_75t_R g172 ( 
.A(n_47),
.Y(n_172)
);

CKINVDCx20_ASAP7_75t_R g173 ( 
.A(n_32),
.Y(n_173)
);

CKINVDCx5p33_ASAP7_75t_R g174 ( 
.A(n_28),
.Y(n_174)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_87),
.Y(n_175)
);

CKINVDCx5p33_ASAP7_75t_R g176 ( 
.A(n_13),
.Y(n_176)
);

CKINVDCx20_ASAP7_75t_R g177 ( 
.A(n_13),
.Y(n_177)
);

BUFx3_ASAP7_75t_L g178 ( 
.A(n_73),
.Y(n_178)
);

CKINVDCx5p33_ASAP7_75t_R g179 ( 
.A(n_64),
.Y(n_179)
);

BUFx3_ASAP7_75t_L g180 ( 
.A(n_140),
.Y(n_180)
);

INVx2_ASAP7_75t_L g181 ( 
.A(n_95),
.Y(n_181)
);

CKINVDCx5p33_ASAP7_75t_R g182 ( 
.A(n_45),
.Y(n_182)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_130),
.Y(n_183)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_89),
.Y(n_184)
);

CKINVDCx20_ASAP7_75t_R g185 ( 
.A(n_26),
.Y(n_185)
);

CKINVDCx5p33_ASAP7_75t_R g186 ( 
.A(n_144),
.Y(n_186)
);

INVx2_ASAP7_75t_L g187 ( 
.A(n_12),
.Y(n_187)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_113),
.Y(n_188)
);

BUFx5_ASAP7_75t_L g189 ( 
.A(n_76),
.Y(n_189)
);

CKINVDCx5p33_ASAP7_75t_R g190 ( 
.A(n_91),
.Y(n_190)
);

CKINVDCx20_ASAP7_75t_R g191 ( 
.A(n_61),
.Y(n_191)
);

CKINVDCx5p33_ASAP7_75t_R g192 ( 
.A(n_41),
.Y(n_192)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_79),
.Y(n_193)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_17),
.Y(n_194)
);

CKINVDCx5p33_ASAP7_75t_R g195 ( 
.A(n_29),
.Y(n_195)
);

CKINVDCx5p33_ASAP7_75t_R g196 ( 
.A(n_1),
.Y(n_196)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_112),
.Y(n_197)
);

CKINVDCx20_ASAP7_75t_R g198 ( 
.A(n_124),
.Y(n_198)
);

BUFx3_ASAP7_75t_L g199 ( 
.A(n_109),
.Y(n_199)
);

CKINVDCx5p33_ASAP7_75t_R g200 ( 
.A(n_141),
.Y(n_200)
);

CKINVDCx5p33_ASAP7_75t_R g201 ( 
.A(n_56),
.Y(n_201)
);

CKINVDCx5p33_ASAP7_75t_R g202 ( 
.A(n_103),
.Y(n_202)
);

CKINVDCx5p33_ASAP7_75t_R g203 ( 
.A(n_88),
.Y(n_203)
);

CKINVDCx5p33_ASAP7_75t_R g204 ( 
.A(n_23),
.Y(n_204)
);

CKINVDCx5p33_ASAP7_75t_R g205 ( 
.A(n_136),
.Y(n_205)
);

CKINVDCx5p33_ASAP7_75t_R g206 ( 
.A(n_84),
.Y(n_206)
);

CKINVDCx5p33_ASAP7_75t_R g207 ( 
.A(n_128),
.Y(n_207)
);

BUFx10_ASAP7_75t_L g208 ( 
.A(n_69),
.Y(n_208)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_133),
.Y(n_209)
);

INVx1_ASAP7_75t_SL g210 ( 
.A(n_120),
.Y(n_210)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_118),
.Y(n_211)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_60),
.Y(n_212)
);

CKINVDCx5p33_ASAP7_75t_R g213 ( 
.A(n_58),
.Y(n_213)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_129),
.Y(n_214)
);

CKINVDCx5p33_ASAP7_75t_R g215 ( 
.A(n_7),
.Y(n_215)
);

INVx1_ASAP7_75t_SL g216 ( 
.A(n_122),
.Y(n_216)
);

CKINVDCx5p33_ASAP7_75t_R g217 ( 
.A(n_48),
.Y(n_217)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_127),
.Y(n_218)
);

CKINVDCx5p33_ASAP7_75t_R g219 ( 
.A(n_92),
.Y(n_219)
);

CKINVDCx5p33_ASAP7_75t_R g220 ( 
.A(n_110),
.Y(n_220)
);

BUFx8_ASAP7_75t_SL g221 ( 
.A(n_131),
.Y(n_221)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_132),
.Y(n_222)
);

HB1xp67_ASAP7_75t_L g223 ( 
.A(n_34),
.Y(n_223)
);

CKINVDCx5p33_ASAP7_75t_R g224 ( 
.A(n_49),
.Y(n_224)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_22),
.Y(n_225)
);

CKINVDCx5p33_ASAP7_75t_R g226 ( 
.A(n_125),
.Y(n_226)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_42),
.Y(n_227)
);

CKINVDCx20_ASAP7_75t_R g228 ( 
.A(n_156),
.Y(n_228)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_160),
.Y(n_229)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_160),
.Y(n_230)
);

CKINVDCx5p33_ASAP7_75t_R g231 ( 
.A(n_157),
.Y(n_231)
);

CKINVDCx20_ASAP7_75t_R g232 ( 
.A(n_173),
.Y(n_232)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_160),
.Y(n_233)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_160),
.Y(n_234)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_194),
.Y(n_235)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_225),
.Y(n_236)
);

INVxp67_ASAP7_75t_SL g237 ( 
.A(n_223),
.Y(n_237)
);

INVxp67_ASAP7_75t_SL g238 ( 
.A(n_170),
.Y(n_238)
);

HB1xp67_ASAP7_75t_L g239 ( 
.A(n_159),
.Y(n_239)
);

INVxp33_ASAP7_75t_SL g240 ( 
.A(n_165),
.Y(n_240)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_187),
.Y(n_241)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_187),
.Y(n_242)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_170),
.Y(n_243)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_178),
.Y(n_244)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_178),
.Y(n_245)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_180),
.Y(n_246)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_180),
.Y(n_247)
);

CKINVDCx5p33_ASAP7_75t_R g248 ( 
.A(n_169),
.Y(n_248)
);

INVxp33_ASAP7_75t_SL g249 ( 
.A(n_176),
.Y(n_249)
);

CKINVDCx5p33_ASAP7_75t_R g250 ( 
.A(n_196),
.Y(n_250)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_199),
.Y(n_251)
);

INVxp33_ASAP7_75t_SL g252 ( 
.A(n_204),
.Y(n_252)
);

CKINVDCx20_ASAP7_75t_R g253 ( 
.A(n_191),
.Y(n_253)
);

CKINVDCx5p33_ASAP7_75t_R g254 ( 
.A(n_215),
.Y(n_254)
);

HB1xp67_ASAP7_75t_L g255 ( 
.A(n_177),
.Y(n_255)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_171),
.Y(n_256)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_199),
.Y(n_257)
);

INVxp33_ASAP7_75t_SL g258 ( 
.A(n_158),
.Y(n_258)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_162),
.Y(n_259)
);

INVxp67_ASAP7_75t_L g260 ( 
.A(n_221),
.Y(n_260)
);

CKINVDCx20_ASAP7_75t_R g261 ( 
.A(n_198),
.Y(n_261)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_175),
.Y(n_262)
);

INVxp33_ASAP7_75t_SL g263 ( 
.A(n_161),
.Y(n_263)
);

CKINVDCx5p33_ASAP7_75t_R g264 ( 
.A(n_221),
.Y(n_264)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_171),
.Y(n_265)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_183),
.Y(n_266)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_184),
.Y(n_267)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_188),
.Y(n_268)
);

INVxp67_ASAP7_75t_SL g269 ( 
.A(n_193),
.Y(n_269)
);

INVx2_ASAP7_75t_L g270 ( 
.A(n_189),
.Y(n_270)
);

INVxp67_ASAP7_75t_SL g271 ( 
.A(n_197),
.Y(n_271)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_181),
.Y(n_272)
);

INVx2_ASAP7_75t_L g273 ( 
.A(n_270),
.Y(n_273)
);

NAND2xp5_ASAP7_75t_L g274 ( 
.A(n_238),
.B(n_181),
.Y(n_274)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_229),
.Y(n_275)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_230),
.Y(n_276)
);

INVx4_ASAP7_75t_L g277 ( 
.A(n_270),
.Y(n_277)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_233),
.Y(n_278)
);

AND2x2_ASAP7_75t_L g279 ( 
.A(n_243),
.B(n_168),
.Y(n_279)
);

NAND2xp5_ASAP7_75t_L g280 ( 
.A(n_269),
.B(n_271),
.Y(n_280)
);

INVx2_ASAP7_75t_L g281 ( 
.A(n_234),
.Y(n_281)
);

CKINVDCx5p33_ASAP7_75t_R g282 ( 
.A(n_264),
.Y(n_282)
);

CKINVDCx5p33_ASAP7_75t_R g283 ( 
.A(n_264),
.Y(n_283)
);

CKINVDCx5p33_ASAP7_75t_R g284 ( 
.A(n_258),
.Y(n_284)
);

INVx2_ASAP7_75t_L g285 ( 
.A(n_256),
.Y(n_285)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_272),
.Y(n_286)
);

INVxp67_ASAP7_75t_L g287 ( 
.A(n_239),
.Y(n_287)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_256),
.Y(n_288)
);

INVx6_ASAP7_75t_L g289 ( 
.A(n_259),
.Y(n_289)
);

NAND2xp5_ASAP7_75t_L g290 ( 
.A(n_237),
.B(n_258),
.Y(n_290)
);

INVx2_ASAP7_75t_L g291 ( 
.A(n_265),
.Y(n_291)
);

CKINVDCx5p33_ASAP7_75t_R g292 ( 
.A(n_263),
.Y(n_292)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_265),
.Y(n_293)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_272),
.Y(n_294)
);

HB1xp67_ASAP7_75t_L g295 ( 
.A(n_231),
.Y(n_295)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_241),
.Y(n_296)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_241),
.Y(n_297)
);

INVx2_ASAP7_75t_L g298 ( 
.A(n_242),
.Y(n_298)
);

INVx2_ASAP7_75t_L g299 ( 
.A(n_242),
.Y(n_299)
);

NAND2xp5_ASAP7_75t_L g300 ( 
.A(n_263),
.B(n_209),
.Y(n_300)
);

INVx2_ASAP7_75t_L g301 ( 
.A(n_262),
.Y(n_301)
);

NAND2xp5_ASAP7_75t_L g302 ( 
.A(n_244),
.B(n_211),
.Y(n_302)
);

NAND2xp5_ASAP7_75t_L g303 ( 
.A(n_245),
.B(n_212),
.Y(n_303)
);

INVx2_ASAP7_75t_L g304 ( 
.A(n_266),
.Y(n_304)
);

CKINVDCx6p67_ASAP7_75t_R g305 ( 
.A(n_228),
.Y(n_305)
);

INVx2_ASAP7_75t_L g306 ( 
.A(n_267),
.Y(n_306)
);

INVx2_ASAP7_75t_L g307 ( 
.A(n_268),
.Y(n_307)
);

BUFx6f_ASAP7_75t_L g308 ( 
.A(n_235),
.Y(n_308)
);

AND2x4_ASAP7_75t_L g309 ( 
.A(n_246),
.B(n_214),
.Y(n_309)
);

HB1xp67_ASAP7_75t_L g310 ( 
.A(n_231),
.Y(n_310)
);

INVx2_ASAP7_75t_L g311 ( 
.A(n_236),
.Y(n_311)
);

XNOR2xp5_ASAP7_75t_L g312 ( 
.A(n_255),
.B(n_185),
.Y(n_312)
);

CKINVDCx16_ASAP7_75t_R g313 ( 
.A(n_232),
.Y(n_313)
);

NAND2xp5_ASAP7_75t_L g314 ( 
.A(n_247),
.B(n_218),
.Y(n_314)
);

HB1xp67_ASAP7_75t_L g315 ( 
.A(n_248),
.Y(n_315)
);

INVx3_ASAP7_75t_L g316 ( 
.A(n_251),
.Y(n_316)
);

AND2x2_ASAP7_75t_L g317 ( 
.A(n_257),
.B(n_168),
.Y(n_317)
);

BUFx6f_ASAP7_75t_L g318 ( 
.A(n_248),
.Y(n_318)
);

CKINVDCx5p33_ASAP7_75t_R g319 ( 
.A(n_250),
.Y(n_319)
);

NOR2xp33_ASAP7_75t_L g320 ( 
.A(n_240),
.B(n_210),
.Y(n_320)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_250),
.Y(n_321)
);

HB1xp67_ASAP7_75t_L g322 ( 
.A(n_254),
.Y(n_322)
);

INVx2_ASAP7_75t_L g323 ( 
.A(n_273),
.Y(n_323)
);

BUFx2_ASAP7_75t_L g324 ( 
.A(n_287),
.Y(n_324)
);

NAND2xp5_ASAP7_75t_SL g325 ( 
.A(n_320),
.B(n_240),
.Y(n_325)
);

INVxp67_ASAP7_75t_SL g326 ( 
.A(n_273),
.Y(n_326)
);

INVx3_ASAP7_75t_L g327 ( 
.A(n_277),
.Y(n_327)
);

INVx2_ASAP7_75t_L g328 ( 
.A(n_273),
.Y(n_328)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_277),
.Y(n_329)
);

AOI22xp33_ASAP7_75t_L g330 ( 
.A1(n_309),
.A2(n_252),
.B1(n_249),
.B2(n_222),
.Y(n_330)
);

INVx3_ASAP7_75t_L g331 ( 
.A(n_277),
.Y(n_331)
);

BUFx3_ASAP7_75t_L g332 ( 
.A(n_309),
.Y(n_332)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_277),
.Y(n_333)
);

AOI22xp33_ASAP7_75t_L g334 ( 
.A1(n_309),
.A2(n_252),
.B1(n_249),
.B2(n_227),
.Y(n_334)
);

INVx3_ASAP7_75t_L g335 ( 
.A(n_308),
.Y(n_335)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_308),
.Y(n_336)
);

NAND2xp5_ASAP7_75t_L g337 ( 
.A(n_280),
.B(n_254),
.Y(n_337)
);

INVx2_ASAP7_75t_L g338 ( 
.A(n_281),
.Y(n_338)
);

NAND3xp33_ASAP7_75t_L g339 ( 
.A(n_274),
.B(n_260),
.C(n_164),
.Y(n_339)
);

INVx2_ASAP7_75t_L g340 ( 
.A(n_281),
.Y(n_340)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_308),
.Y(n_341)
);

BUFx10_ASAP7_75t_L g342 ( 
.A(n_282),
.Y(n_342)
);

NAND2xp5_ASAP7_75t_SL g343 ( 
.A(n_318),
.B(n_168),
.Y(n_343)
);

AND2x6_ASAP7_75t_L g344 ( 
.A(n_321),
.B(n_216),
.Y(n_344)
);

INVx3_ASAP7_75t_L g345 ( 
.A(n_308),
.Y(n_345)
);

NAND2xp5_ASAP7_75t_L g346 ( 
.A(n_300),
.B(n_163),
.Y(n_346)
);

INVx4_ASAP7_75t_L g347 ( 
.A(n_308),
.Y(n_347)
);

OAI22xp33_ASAP7_75t_SL g348 ( 
.A1(n_290),
.A2(n_166),
.B1(n_167),
.B2(n_172),
.Y(n_348)
);

INVx2_ASAP7_75t_L g349 ( 
.A(n_281),
.Y(n_349)
);

NAND2xp33_ASAP7_75t_SL g350 ( 
.A(n_321),
.B(n_318),
.Y(n_350)
);

NAND3xp33_ASAP7_75t_L g351 ( 
.A(n_302),
.B(n_179),
.C(n_174),
.Y(n_351)
);

NAND2xp5_ASAP7_75t_L g352 ( 
.A(n_316),
.B(n_182),
.Y(n_352)
);

INVx2_ASAP7_75t_L g353 ( 
.A(n_291),
.Y(n_353)
);

INVx2_ASAP7_75t_L g354 ( 
.A(n_291),
.Y(n_354)
);

NOR2xp33_ASAP7_75t_L g355 ( 
.A(n_318),
.B(n_261),
.Y(n_355)
);

NAND2xp5_ASAP7_75t_SL g356 ( 
.A(n_318),
.B(n_284),
.Y(n_356)
);

OR2x2_ASAP7_75t_L g357 ( 
.A(n_279),
.B(n_186),
.Y(n_357)
);

AOI22xp33_ASAP7_75t_L g358 ( 
.A1(n_309),
.A2(n_189),
.B1(n_208),
.B2(n_224),
.Y(n_358)
);

NAND3xp33_ASAP7_75t_L g359 ( 
.A(n_303),
.B(n_192),
.C(n_190),
.Y(n_359)
);

INVx2_ASAP7_75t_L g360 ( 
.A(n_291),
.Y(n_360)
);

NAND3xp33_ASAP7_75t_L g361 ( 
.A(n_314),
.B(n_200),
.C(n_195),
.Y(n_361)
);

INVx1_ASAP7_75t_L g362 ( 
.A(n_308),
.Y(n_362)
);

NOR2xp33_ASAP7_75t_L g363 ( 
.A(n_318),
.B(n_253),
.Y(n_363)
);

NAND2xp5_ASAP7_75t_L g364 ( 
.A(n_316),
.B(n_201),
.Y(n_364)
);

INVx2_ASAP7_75t_L g365 ( 
.A(n_298),
.Y(n_365)
);

NAND2xp5_ASAP7_75t_L g366 ( 
.A(n_316),
.B(n_202),
.Y(n_366)
);

INVx2_ASAP7_75t_L g367 ( 
.A(n_298),
.Y(n_367)
);

INVx1_ASAP7_75t_L g368 ( 
.A(n_307),
.Y(n_368)
);

NAND2xp5_ASAP7_75t_L g369 ( 
.A(n_316),
.B(n_301),
.Y(n_369)
);

INVx1_ASAP7_75t_L g370 ( 
.A(n_307),
.Y(n_370)
);

NAND2xp5_ASAP7_75t_L g371 ( 
.A(n_301),
.B(n_203),
.Y(n_371)
);

INVx1_ASAP7_75t_L g372 ( 
.A(n_307),
.Y(n_372)
);

INVx1_ASAP7_75t_L g373 ( 
.A(n_275),
.Y(n_373)
);

BUFx3_ASAP7_75t_L g374 ( 
.A(n_289),
.Y(n_374)
);

INVx2_ASAP7_75t_L g375 ( 
.A(n_298),
.Y(n_375)
);

NAND2xp5_ASAP7_75t_SL g376 ( 
.A(n_318),
.B(n_208),
.Y(n_376)
);

NOR2xp33_ASAP7_75t_L g377 ( 
.A(n_319),
.B(n_292),
.Y(n_377)
);

CKINVDCx5p33_ASAP7_75t_R g378 ( 
.A(n_305),
.Y(n_378)
);

NAND2xp5_ASAP7_75t_L g379 ( 
.A(n_304),
.B(n_205),
.Y(n_379)
);

INVx1_ASAP7_75t_L g380 ( 
.A(n_275),
.Y(n_380)
);

AOI22xp33_ASAP7_75t_L g381 ( 
.A1(n_279),
.A2(n_189),
.B1(n_208),
.B2(n_219),
.Y(n_381)
);

INVx1_ASAP7_75t_L g382 ( 
.A(n_276),
.Y(n_382)
);

NAND2xp5_ASAP7_75t_L g383 ( 
.A(n_304),
.B(n_206),
.Y(n_383)
);

AND2x2_ASAP7_75t_L g384 ( 
.A(n_317),
.B(n_207),
.Y(n_384)
);

INVx1_ASAP7_75t_L g385 ( 
.A(n_276),
.Y(n_385)
);

INVx2_ASAP7_75t_L g386 ( 
.A(n_285),
.Y(n_386)
);

INVx2_ASAP7_75t_L g387 ( 
.A(n_285),
.Y(n_387)
);

INVx1_ASAP7_75t_L g388 ( 
.A(n_278),
.Y(n_388)
);

INVx1_ASAP7_75t_L g389 ( 
.A(n_373),
.Y(n_389)
);

INVxp67_ASAP7_75t_L g390 ( 
.A(n_324),
.Y(n_390)
);

AOI22xp5_ASAP7_75t_L g391 ( 
.A1(n_350),
.A2(n_322),
.B1(n_295),
.B2(n_315),
.Y(n_391)
);

NAND2xp5_ASAP7_75t_L g392 ( 
.A(n_327),
.B(n_317),
.Y(n_392)
);

INVx1_ASAP7_75t_L g393 ( 
.A(n_373),
.Y(n_393)
);

NOR2xp33_ASAP7_75t_L g394 ( 
.A(n_337),
.B(n_310),
.Y(n_394)
);

INVx1_ASAP7_75t_L g395 ( 
.A(n_380),
.Y(n_395)
);

INVx1_ASAP7_75t_L g396 ( 
.A(n_380),
.Y(n_396)
);

NAND2xp5_ASAP7_75t_L g397 ( 
.A(n_327),
.B(n_306),
.Y(n_397)
);

NAND2xp5_ASAP7_75t_L g398 ( 
.A(n_327),
.B(n_306),
.Y(n_398)
);

INVx2_ASAP7_75t_L g399 ( 
.A(n_386),
.Y(n_399)
);

NOR2xp33_ASAP7_75t_L g400 ( 
.A(n_325),
.B(n_283),
.Y(n_400)
);

INVx2_ASAP7_75t_L g401 ( 
.A(n_386),
.Y(n_401)
);

INVxp67_ASAP7_75t_L g402 ( 
.A(n_324),
.Y(n_402)
);

INVx2_ASAP7_75t_L g403 ( 
.A(n_387),
.Y(n_403)
);

NAND2x1p5_ASAP7_75t_L g404 ( 
.A(n_332),
.B(n_286),
.Y(n_404)
);

NAND2xp5_ASAP7_75t_L g405 ( 
.A(n_331),
.B(n_289),
.Y(n_405)
);

NAND2xp5_ASAP7_75t_L g406 ( 
.A(n_331),
.B(n_289),
.Y(n_406)
);

NAND2xp5_ASAP7_75t_L g407 ( 
.A(n_331),
.B(n_289),
.Y(n_407)
);

INVx2_ASAP7_75t_L g408 ( 
.A(n_387),
.Y(n_408)
);

INVx1_ASAP7_75t_L g409 ( 
.A(n_382),
.Y(n_409)
);

INVx1_ASAP7_75t_L g410 ( 
.A(n_382),
.Y(n_410)
);

AOI22xp5_ASAP7_75t_L g411 ( 
.A1(n_344),
.A2(n_213),
.B1(n_217),
.B2(n_220),
.Y(n_411)
);

INVxp33_ASAP7_75t_L g412 ( 
.A(n_377),
.Y(n_412)
);

INVx1_ASAP7_75t_L g413 ( 
.A(n_385),
.Y(n_413)
);

NAND2xp5_ASAP7_75t_L g414 ( 
.A(n_329),
.B(n_286),
.Y(n_414)
);

NAND2xp5_ASAP7_75t_L g415 ( 
.A(n_329),
.B(n_333),
.Y(n_415)
);

AOI21xp5_ASAP7_75t_L g416 ( 
.A1(n_333),
.A2(n_311),
.B(n_293),
.Y(n_416)
);

INVx2_ASAP7_75t_L g417 ( 
.A(n_323),
.Y(n_417)
);

NAND2xp5_ASAP7_75t_L g418 ( 
.A(n_332),
.B(n_288),
.Y(n_418)
);

NAND2xp5_ASAP7_75t_SL g419 ( 
.A(n_348),
.B(n_226),
.Y(n_419)
);

NAND2xp5_ASAP7_75t_L g420 ( 
.A(n_326),
.B(n_288),
.Y(n_420)
);

CKINVDCx5p33_ASAP7_75t_R g421 ( 
.A(n_378),
.Y(n_421)
);

NAND2xp5_ASAP7_75t_L g422 ( 
.A(n_346),
.B(n_293),
.Y(n_422)
);

NAND2xp5_ASAP7_75t_SL g423 ( 
.A(n_348),
.B(n_189),
.Y(n_423)
);

AOI22xp5_ASAP7_75t_L g424 ( 
.A1(n_344),
.A2(n_311),
.B1(n_278),
.B2(n_294),
.Y(n_424)
);

INVx2_ASAP7_75t_L g425 ( 
.A(n_323),
.Y(n_425)
);

INVx1_ASAP7_75t_L g426 ( 
.A(n_385),
.Y(n_426)
);

INVx1_ASAP7_75t_L g427 ( 
.A(n_388),
.Y(n_427)
);

NAND2xp5_ASAP7_75t_L g428 ( 
.A(n_352),
.B(n_294),
.Y(n_428)
);

HB1xp67_ASAP7_75t_L g429 ( 
.A(n_384),
.Y(n_429)
);

NAND2xp5_ASAP7_75t_SL g430 ( 
.A(n_384),
.B(n_357),
.Y(n_430)
);

NAND2xp5_ASAP7_75t_L g431 ( 
.A(n_364),
.B(n_311),
.Y(n_431)
);

AOI22xp33_ASAP7_75t_L g432 ( 
.A1(n_344),
.A2(n_189),
.B1(n_297),
.B2(n_296),
.Y(n_432)
);

NOR2xp33_ASAP7_75t_L g433 ( 
.A(n_343),
.B(n_296),
.Y(n_433)
);

AOI22xp33_ASAP7_75t_L g434 ( 
.A1(n_344),
.A2(n_189),
.B1(n_297),
.B2(n_299),
.Y(n_434)
);

INVx2_ASAP7_75t_SL g435 ( 
.A(n_357),
.Y(n_435)
);

NAND2xp5_ASAP7_75t_L g436 ( 
.A(n_366),
.B(n_299),
.Y(n_436)
);

INVx2_ASAP7_75t_SL g437 ( 
.A(n_388),
.Y(n_437)
);

INVxp67_ASAP7_75t_L g438 ( 
.A(n_355),
.Y(n_438)
);

INVx1_ASAP7_75t_L g439 ( 
.A(n_369),
.Y(n_439)
);

NAND2xp33_ASAP7_75t_L g440 ( 
.A(n_344),
.B(n_189),
.Y(n_440)
);

NAND2xp5_ASAP7_75t_SL g441 ( 
.A(n_381),
.B(n_313),
.Y(n_441)
);

AND2x4_ASAP7_75t_L g442 ( 
.A(n_374),
.B(n_30),
.Y(n_442)
);

NAND2xp5_ASAP7_75t_SL g443 ( 
.A(n_351),
.B(n_313),
.Y(n_443)
);

NAND2xp5_ASAP7_75t_L g444 ( 
.A(n_344),
.B(n_31),
.Y(n_444)
);

NAND2xp5_ASAP7_75t_L g445 ( 
.A(n_344),
.B(n_33),
.Y(n_445)
);

BUFx6f_ASAP7_75t_SL g446 ( 
.A(n_342),
.Y(n_446)
);

NOR2xp67_ASAP7_75t_L g447 ( 
.A(n_351),
.B(n_312),
.Y(n_447)
);

NAND2xp5_ASAP7_75t_L g448 ( 
.A(n_371),
.B(n_35),
.Y(n_448)
);

OAI22xp5_ASAP7_75t_L g449 ( 
.A1(n_358),
.A2(n_305),
.B1(n_312),
.B2(n_86),
.Y(n_449)
);

NOR2xp33_ASAP7_75t_L g450 ( 
.A(n_376),
.B(n_339),
.Y(n_450)
);

NAND2xp5_ASAP7_75t_L g451 ( 
.A(n_379),
.B(n_36),
.Y(n_451)
);

HB1xp67_ASAP7_75t_L g452 ( 
.A(n_363),
.Y(n_452)
);

BUFx12f_ASAP7_75t_SL g453 ( 
.A(n_378),
.Y(n_453)
);

INVx2_ASAP7_75t_L g454 ( 
.A(n_328),
.Y(n_454)
);

NAND2xp5_ASAP7_75t_SL g455 ( 
.A(n_359),
.B(n_361),
.Y(n_455)
);

INVx1_ASAP7_75t_SL g456 ( 
.A(n_435),
.Y(n_456)
);

NAND2xp5_ASAP7_75t_SL g457 ( 
.A(n_392),
.B(n_356),
.Y(n_457)
);

AOI22xp5_ASAP7_75t_L g458 ( 
.A1(n_394),
.A2(n_359),
.B1(n_361),
.B2(n_383),
.Y(n_458)
);

AO21x1_ASAP7_75t_L g459 ( 
.A1(n_455),
.A2(n_341),
.B(n_336),
.Y(n_459)
);

INVx1_ASAP7_75t_L g460 ( 
.A(n_389),
.Y(n_460)
);

NAND2xp5_ASAP7_75t_SL g461 ( 
.A(n_438),
.B(n_374),
.Y(n_461)
);

NAND2xp5_ASAP7_75t_L g462 ( 
.A(n_422),
.B(n_330),
.Y(n_462)
);

BUFx3_ASAP7_75t_L g463 ( 
.A(n_442),
.Y(n_463)
);

INVx1_ASAP7_75t_L g464 ( 
.A(n_393),
.Y(n_464)
);

INVx1_ASAP7_75t_L g465 ( 
.A(n_395),
.Y(n_465)
);

INVx1_ASAP7_75t_L g466 ( 
.A(n_396),
.Y(n_466)
);

NAND2xp5_ASAP7_75t_L g467 ( 
.A(n_439),
.B(n_334),
.Y(n_467)
);

INVx2_ASAP7_75t_SL g468 ( 
.A(n_437),
.Y(n_468)
);

OAI22xp5_ASAP7_75t_L g469 ( 
.A1(n_394),
.A2(n_372),
.B1(n_370),
.B2(n_368),
.Y(n_469)
);

AND2x4_ASAP7_75t_L g470 ( 
.A(n_442),
.B(n_368),
.Y(n_470)
);

AOI22xp5_ASAP7_75t_L g471 ( 
.A1(n_450),
.A2(n_372),
.B1(n_370),
.B2(n_341),
.Y(n_471)
);

NAND2xp5_ASAP7_75t_L g472 ( 
.A(n_409),
.B(n_335),
.Y(n_472)
);

INVx1_ASAP7_75t_L g473 ( 
.A(n_410),
.Y(n_473)
);

INVx1_ASAP7_75t_L g474 ( 
.A(n_413),
.Y(n_474)
);

AOI22xp33_ASAP7_75t_L g475 ( 
.A1(n_455),
.A2(n_336),
.B1(n_362),
.B2(n_365),
.Y(n_475)
);

INVx1_ASAP7_75t_SL g476 ( 
.A(n_429),
.Y(n_476)
);

CKINVDCx5p33_ASAP7_75t_R g477 ( 
.A(n_421),
.Y(n_477)
);

NOR2xp33_ASAP7_75t_L g478 ( 
.A(n_412),
.B(n_452),
.Y(n_478)
);

BUFx3_ASAP7_75t_L g479 ( 
.A(n_404),
.Y(n_479)
);

NAND2xp5_ASAP7_75t_L g480 ( 
.A(n_426),
.B(n_335),
.Y(n_480)
);

INVx2_ASAP7_75t_L g481 ( 
.A(n_399),
.Y(n_481)
);

INVx3_ASAP7_75t_L g482 ( 
.A(n_399),
.Y(n_482)
);

AOI22xp33_ASAP7_75t_L g483 ( 
.A1(n_423),
.A2(n_362),
.B1(n_375),
.B2(n_365),
.Y(n_483)
);

INVx2_ASAP7_75t_SL g484 ( 
.A(n_430),
.Y(n_484)
);

OR2x6_ASAP7_75t_L g485 ( 
.A(n_404),
.B(n_347),
.Y(n_485)
);

INVx2_ASAP7_75t_SL g486 ( 
.A(n_418),
.Y(n_486)
);

INVx1_ASAP7_75t_L g487 ( 
.A(n_427),
.Y(n_487)
);

CKINVDCx5p33_ASAP7_75t_R g488 ( 
.A(n_446),
.Y(n_488)
);

BUFx2_ASAP7_75t_L g489 ( 
.A(n_390),
.Y(n_489)
);

INVx3_ASAP7_75t_L g490 ( 
.A(n_401),
.Y(n_490)
);

NOR2xp33_ASAP7_75t_L g491 ( 
.A(n_402),
.B(n_342),
.Y(n_491)
);

INVx2_ASAP7_75t_L g492 ( 
.A(n_401),
.Y(n_492)
);

AOI22xp5_ASAP7_75t_L g493 ( 
.A1(n_450),
.A2(n_335),
.B1(n_345),
.B2(n_347),
.Y(n_493)
);

NAND2xp5_ASAP7_75t_SL g494 ( 
.A(n_448),
.B(n_342),
.Y(n_494)
);

INVx2_ASAP7_75t_L g495 ( 
.A(n_403),
.Y(n_495)
);

AND2x4_ASAP7_75t_SL g496 ( 
.A(n_391),
.B(n_347),
.Y(n_496)
);

INVxp67_ASAP7_75t_L g497 ( 
.A(n_400),
.Y(n_497)
);

INVx2_ASAP7_75t_L g498 ( 
.A(n_403),
.Y(n_498)
);

A2O1A1Ixp33_ASAP7_75t_L g499 ( 
.A1(n_433),
.A2(n_375),
.B(n_367),
.C(n_360),
.Y(n_499)
);

BUFx2_ASAP7_75t_L g500 ( 
.A(n_453),
.Y(n_500)
);

NAND2xp5_ASAP7_75t_L g501 ( 
.A(n_428),
.B(n_345),
.Y(n_501)
);

INVx2_ASAP7_75t_SL g502 ( 
.A(n_419),
.Y(n_502)
);

NAND2xp5_ASAP7_75t_L g503 ( 
.A(n_486),
.B(n_433),
.Y(n_503)
);

A2O1A1Ixp33_ASAP7_75t_L g504 ( 
.A1(n_462),
.A2(n_400),
.B(n_449),
.C(n_447),
.Y(n_504)
);

A2O1A1Ixp33_ASAP7_75t_L g505 ( 
.A1(n_467),
.A2(n_440),
.B(n_431),
.C(n_411),
.Y(n_505)
);

AOI21x1_ASAP7_75t_L g506 ( 
.A1(n_457),
.A2(n_415),
.B(n_414),
.Y(n_506)
);

AOI21xp5_ASAP7_75t_L g507 ( 
.A1(n_501),
.A2(n_406),
.B(n_405),
.Y(n_507)
);

NAND2xp5_ASAP7_75t_SL g508 ( 
.A(n_497),
.B(n_441),
.Y(n_508)
);

NOR2xp33_ASAP7_75t_L g509 ( 
.A(n_478),
.B(n_476),
.Y(n_509)
);

AOI21xp5_ASAP7_75t_L g510 ( 
.A1(n_485),
.A2(n_407),
.B(n_398),
.Y(n_510)
);

INVx1_ASAP7_75t_L g511 ( 
.A(n_460),
.Y(n_511)
);

AOI21xp5_ASAP7_75t_L g512 ( 
.A1(n_485),
.A2(n_397),
.B(n_436),
.Y(n_512)
);

CKINVDCx5p33_ASAP7_75t_R g513 ( 
.A(n_477),
.Y(n_513)
);

BUFx2_ASAP7_75t_L g514 ( 
.A(n_489),
.Y(n_514)
);

NAND2xp5_ASAP7_75t_L g515 ( 
.A(n_486),
.B(n_420),
.Y(n_515)
);

AOI21xp5_ASAP7_75t_L g516 ( 
.A1(n_485),
.A2(n_451),
.B(n_445),
.Y(n_516)
);

NAND2xp5_ASAP7_75t_SL g517 ( 
.A(n_468),
.B(n_443),
.Y(n_517)
);

AOI21xp5_ASAP7_75t_L g518 ( 
.A1(n_485),
.A2(n_444),
.B(n_434),
.Y(n_518)
);

INVx2_ASAP7_75t_L g519 ( 
.A(n_482),
.Y(n_519)
);

AOI21xp5_ASAP7_75t_L g520 ( 
.A1(n_470),
.A2(n_457),
.B(n_472),
.Y(n_520)
);

BUFx12f_ASAP7_75t_L g521 ( 
.A(n_500),
.Y(n_521)
);

NAND2xp5_ASAP7_75t_SL g522 ( 
.A(n_468),
.B(n_443),
.Y(n_522)
);

NAND2xp33_ASAP7_75t_R g523 ( 
.A(n_477),
.B(n_408),
.Y(n_523)
);

NAND2xp5_ASAP7_75t_L g524 ( 
.A(n_464),
.B(n_408),
.Y(n_524)
);

NOR2xp33_ASAP7_75t_SL g525 ( 
.A(n_488),
.B(n_446),
.Y(n_525)
);

AOI21xp5_ASAP7_75t_L g526 ( 
.A1(n_470),
.A2(n_434),
.B(n_432),
.Y(n_526)
);

AOI21xp5_ASAP7_75t_L g527 ( 
.A1(n_470),
.A2(n_432),
.B(n_416),
.Y(n_527)
);

BUFx6f_ASAP7_75t_L g528 ( 
.A(n_479),
.Y(n_528)
);

CKINVDCx5p33_ASAP7_75t_R g529 ( 
.A(n_488),
.Y(n_529)
);

AND2x2_ASAP7_75t_L g530 ( 
.A(n_456),
.B(n_424),
.Y(n_530)
);

BUFx3_ASAP7_75t_L g531 ( 
.A(n_463),
.Y(n_531)
);

NAND2xp5_ASAP7_75t_SL g532 ( 
.A(n_458),
.B(n_417),
.Y(n_532)
);

AOI21xp5_ASAP7_75t_L g533 ( 
.A1(n_480),
.A2(n_454),
.B(n_425),
.Y(n_533)
);

INVx2_ASAP7_75t_L g534 ( 
.A(n_482),
.Y(n_534)
);

NAND2xp5_ASAP7_75t_L g535 ( 
.A(n_465),
.B(n_417),
.Y(n_535)
);

AOI22xp5_ASAP7_75t_L g536 ( 
.A1(n_484),
.A2(n_423),
.B1(n_345),
.B2(n_454),
.Y(n_536)
);

NAND2x1p5_ASAP7_75t_L g537 ( 
.A(n_479),
.B(n_425),
.Y(n_537)
);

INVx2_ASAP7_75t_SL g538 ( 
.A(n_502),
.Y(n_538)
);

NAND2xp5_ASAP7_75t_SL g539 ( 
.A(n_463),
.B(n_353),
.Y(n_539)
);

AO31x2_ASAP7_75t_L g540 ( 
.A1(n_518),
.A2(n_459),
.A3(n_499),
.B(n_469),
.Y(n_540)
);

INVx1_ASAP7_75t_L g541 ( 
.A(n_511),
.Y(n_541)
);

INVx6_ASAP7_75t_L g542 ( 
.A(n_521),
.Y(n_542)
);

OAI21x1_ASAP7_75t_L g543 ( 
.A1(n_510),
.A2(n_483),
.B(n_475),
.Y(n_543)
);

OAI21xp5_ASAP7_75t_L g544 ( 
.A1(n_505),
.A2(n_499),
.B(n_471),
.Y(n_544)
);

INVx2_ASAP7_75t_L g545 ( 
.A(n_519),
.Y(n_545)
);

AND2x4_ASAP7_75t_L g546 ( 
.A(n_531),
.B(n_466),
.Y(n_546)
);

OR2x2_ASAP7_75t_L g547 ( 
.A(n_514),
.B(n_461),
.Y(n_547)
);

INVx1_ASAP7_75t_L g548 ( 
.A(n_524),
.Y(n_548)
);

NOR2xp33_ASAP7_75t_SL g549 ( 
.A(n_513),
.B(n_491),
.Y(n_549)
);

NAND2xp5_ASAP7_75t_SL g550 ( 
.A(n_509),
.B(n_473),
.Y(n_550)
);

INVxp67_ASAP7_75t_SL g551 ( 
.A(n_523),
.Y(n_551)
);

INVx2_ASAP7_75t_SL g552 ( 
.A(n_528),
.Y(n_552)
);

NAND2xp5_ASAP7_75t_SL g553 ( 
.A(n_509),
.B(n_504),
.Y(n_553)
);

AO31x2_ASAP7_75t_L g554 ( 
.A1(n_516),
.A2(n_498),
.A3(n_481),
.B(n_495),
.Y(n_554)
);

AOI21x1_ASAP7_75t_L g555 ( 
.A1(n_532),
.A2(n_494),
.B(n_461),
.Y(n_555)
);

NAND2xp5_ASAP7_75t_L g556 ( 
.A(n_503),
.B(n_474),
.Y(n_556)
);

OAI22xp5_ASAP7_75t_L g557 ( 
.A1(n_526),
.A2(n_487),
.B1(n_496),
.B2(n_494),
.Y(n_557)
);

NAND2xp5_ASAP7_75t_L g558 ( 
.A(n_515),
.B(n_496),
.Y(n_558)
);

BUFx4_ASAP7_75t_SL g559 ( 
.A(n_529),
.Y(n_559)
);

AND2x2_ASAP7_75t_L g560 ( 
.A(n_530),
.B(n_481),
.Y(n_560)
);

NAND2xp5_ASAP7_75t_L g561 ( 
.A(n_508),
.B(n_492),
.Y(n_561)
);

A2O1A1Ixp33_ASAP7_75t_L g562 ( 
.A1(n_520),
.A2(n_493),
.B(n_490),
.C(n_482),
.Y(n_562)
);

NAND2x1_ASAP7_75t_L g563 ( 
.A(n_534),
.B(n_490),
.Y(n_563)
);

AO21x2_ASAP7_75t_L g564 ( 
.A1(n_532),
.A2(n_512),
.B(n_507),
.Y(n_564)
);

NOR2xp33_ASAP7_75t_L g565 ( 
.A(n_517),
.B(n_492),
.Y(n_565)
);

NAND3xp33_ASAP7_75t_L g566 ( 
.A(n_522),
.B(n_498),
.C(n_495),
.Y(n_566)
);

OAI21xp5_ASAP7_75t_L g567 ( 
.A1(n_527),
.A2(n_490),
.B(n_367),
.Y(n_567)
);

AOI21xp5_ASAP7_75t_L g568 ( 
.A1(n_533),
.A2(n_328),
.B(n_354),
.Y(n_568)
);

NOR4xp25_ASAP7_75t_L g569 ( 
.A(n_539),
.B(n_349),
.C(n_340),
.D(n_338),
.Y(n_569)
);

OAI21xp5_ASAP7_75t_L g570 ( 
.A1(n_506),
.A2(n_360),
.B(n_354),
.Y(n_570)
);

NAND2xp5_ASAP7_75t_L g571 ( 
.A(n_538),
.B(n_353),
.Y(n_571)
);

NAND2xp5_ASAP7_75t_L g572 ( 
.A(n_535),
.B(n_528),
.Y(n_572)
);

NAND2xp5_ASAP7_75t_L g573 ( 
.A(n_528),
.B(n_338),
.Y(n_573)
);

NAND2x1p5_ASAP7_75t_L g574 ( 
.A(n_553),
.B(n_528),
.Y(n_574)
);

O2A1O1Ixp5_ASAP7_75t_L g575 ( 
.A1(n_544),
.A2(n_539),
.B(n_523),
.C(n_349),
.Y(n_575)
);

AO21x2_ASAP7_75t_L g576 ( 
.A1(n_544),
.A2(n_536),
.B(n_340),
.Y(n_576)
);

OAI21x1_ASAP7_75t_L g577 ( 
.A1(n_570),
.A2(n_537),
.B(n_525),
.Y(n_577)
);

AOI22xp33_ASAP7_75t_L g578 ( 
.A1(n_551),
.A2(n_537),
.B1(n_1),
.B2(n_2),
.Y(n_578)
);

OAI21xp5_ASAP7_75t_L g579 ( 
.A1(n_557),
.A2(n_0),
.B(n_2),
.Y(n_579)
);

OAI21xp33_ASAP7_75t_SL g580 ( 
.A1(n_548),
.A2(n_90),
.B(n_154),
.Y(n_580)
);

INVx3_ASAP7_75t_L g581 ( 
.A(n_554),
.Y(n_581)
);

AND2x2_ASAP7_75t_L g582 ( 
.A(n_560),
.B(n_37),
.Y(n_582)
);

OAI21x1_ASAP7_75t_SL g583 ( 
.A1(n_555),
.A2(n_85),
.B(n_153),
.Y(n_583)
);

AO21x2_ASAP7_75t_L g584 ( 
.A1(n_564),
.A2(n_83),
.B(n_152),
.Y(n_584)
);

OAI21x1_ASAP7_75t_L g585 ( 
.A1(n_570),
.A2(n_82),
.B(n_151),
.Y(n_585)
);

OAI21x1_ASAP7_75t_L g586 ( 
.A1(n_567),
.A2(n_81),
.B(n_150),
.Y(n_586)
);

A2O1A1Ixp33_ASAP7_75t_L g587 ( 
.A1(n_557),
.A2(n_0),
.B(n_3),
.C(n_4),
.Y(n_587)
);

OA21x2_ASAP7_75t_L g588 ( 
.A1(n_543),
.A2(n_3),
.B(n_5),
.Y(n_588)
);

AO21x2_ASAP7_75t_L g589 ( 
.A1(n_564),
.A2(n_96),
.B(n_149),
.Y(n_589)
);

AO31x2_ASAP7_75t_L g590 ( 
.A1(n_562),
.A2(n_5),
.A3(n_6),
.B(n_7),
.Y(n_590)
);

OAI21x1_ASAP7_75t_L g591 ( 
.A1(n_567),
.A2(n_97),
.B(n_148),
.Y(n_591)
);

OAI21xp5_ASAP7_75t_L g592 ( 
.A1(n_558),
.A2(n_6),
.B(n_8),
.Y(n_592)
);

OAI21x1_ASAP7_75t_L g593 ( 
.A1(n_568),
.A2(n_93),
.B(n_147),
.Y(n_593)
);

INVx1_ASAP7_75t_L g594 ( 
.A(n_541),
.Y(n_594)
);

INVx2_ASAP7_75t_SL g595 ( 
.A(n_552),
.Y(n_595)
);

AND2x4_ASAP7_75t_L g596 ( 
.A(n_545),
.B(n_38),
.Y(n_596)
);

NAND2xp5_ASAP7_75t_L g597 ( 
.A(n_556),
.B(n_8),
.Y(n_597)
);

OAI21xp5_ASAP7_75t_L g598 ( 
.A1(n_550),
.A2(n_9),
.B(n_10),
.Y(n_598)
);

AOI21x1_ASAP7_75t_L g599 ( 
.A1(n_566),
.A2(n_99),
.B(n_146),
.Y(n_599)
);

INVx1_ASAP7_75t_L g600 ( 
.A(n_561),
.Y(n_600)
);

OAI21xp5_ASAP7_75t_L g601 ( 
.A1(n_565),
.A2(n_10),
.B(n_11),
.Y(n_601)
);

INVx2_ASAP7_75t_L g602 ( 
.A(n_554),
.Y(n_602)
);

INVx1_ASAP7_75t_L g603 ( 
.A(n_572),
.Y(n_603)
);

XNOR2xp5_ASAP7_75t_L g604 ( 
.A(n_546),
.B(n_11),
.Y(n_604)
);

OAI21xp5_ASAP7_75t_L g605 ( 
.A1(n_571),
.A2(n_14),
.B(n_15),
.Y(n_605)
);

OAI21x1_ASAP7_75t_L g606 ( 
.A1(n_563),
.A2(n_101),
.B(n_145),
.Y(n_606)
);

AO31x2_ASAP7_75t_L g607 ( 
.A1(n_569),
.A2(n_14),
.A3(n_15),
.B(n_16),
.Y(n_607)
);

INVx1_ASAP7_75t_L g608 ( 
.A(n_573),
.Y(n_608)
);

AOI21x1_ASAP7_75t_L g609 ( 
.A1(n_573),
.A2(n_102),
.B(n_142),
.Y(n_609)
);

AOI21x1_ASAP7_75t_L g610 ( 
.A1(n_554),
.A2(n_98),
.B(n_139),
.Y(n_610)
);

O2A1O1Ixp33_ASAP7_75t_L g611 ( 
.A1(n_547),
.A2(n_16),
.B(n_17),
.C(n_18),
.Y(n_611)
);

OA21x2_ASAP7_75t_L g612 ( 
.A1(n_540),
.A2(n_19),
.B(n_20),
.Y(n_612)
);

HB1xp67_ASAP7_75t_L g613 ( 
.A(n_603),
.Y(n_613)
);

AND2x4_ASAP7_75t_SL g614 ( 
.A(n_596),
.B(n_546),
.Y(n_614)
);

INVx2_ASAP7_75t_L g615 ( 
.A(n_602),
.Y(n_615)
);

OR2x2_ASAP7_75t_L g616 ( 
.A(n_590),
.B(n_540),
.Y(n_616)
);

INVx2_ASAP7_75t_L g617 ( 
.A(n_602),
.Y(n_617)
);

AND2x4_ASAP7_75t_SL g618 ( 
.A(n_596),
.B(n_559),
.Y(n_618)
);

AOI21xp5_ASAP7_75t_SL g619 ( 
.A1(n_579),
.A2(n_587),
.B(n_601),
.Y(n_619)
);

O2A1O1Ixp33_ASAP7_75t_L g620 ( 
.A1(n_587),
.A2(n_549),
.B(n_540),
.C(n_21),
.Y(n_620)
);

AOI21xp5_ASAP7_75t_L g621 ( 
.A1(n_575),
.A2(n_105),
.B(n_155),
.Y(n_621)
);

INVx2_ASAP7_75t_L g622 ( 
.A(n_581),
.Y(n_622)
);

INVx1_ASAP7_75t_L g623 ( 
.A(n_581),
.Y(n_623)
);

AOI21xp5_ASAP7_75t_L g624 ( 
.A1(n_576),
.A2(n_104),
.B(n_138),
.Y(n_624)
);

AND2x4_ASAP7_75t_L g625 ( 
.A(n_594),
.B(n_39),
.Y(n_625)
);

AOI221x1_ASAP7_75t_SL g626 ( 
.A1(n_597),
.A2(n_604),
.B1(n_600),
.B2(n_611),
.C(n_598),
.Y(n_626)
);

INVx1_ASAP7_75t_L g627 ( 
.A(n_581),
.Y(n_627)
);

AND2x2_ASAP7_75t_L g628 ( 
.A(n_590),
.B(n_608),
.Y(n_628)
);

AND2x2_ASAP7_75t_L g629 ( 
.A(n_590),
.B(n_19),
.Y(n_629)
);

OA21x2_ASAP7_75t_L g630 ( 
.A1(n_610),
.A2(n_20),
.B(n_21),
.Y(n_630)
);

INVx2_ASAP7_75t_SL g631 ( 
.A(n_574),
.Y(n_631)
);

AND2x2_ASAP7_75t_L g632 ( 
.A(n_590),
.B(n_612),
.Y(n_632)
);

OAI22xp5_ASAP7_75t_L g633 ( 
.A1(n_578),
.A2(n_542),
.B1(n_23),
.B2(n_24),
.Y(n_633)
);

AND2x4_ASAP7_75t_L g634 ( 
.A(n_596),
.B(n_111),
.Y(n_634)
);

BUFx6f_ASAP7_75t_L g635 ( 
.A(n_574),
.Y(n_635)
);

AND2x2_ASAP7_75t_L g636 ( 
.A(n_590),
.B(n_22),
.Y(n_636)
);

INVx1_ASAP7_75t_L g637 ( 
.A(n_612),
.Y(n_637)
);

INVx1_ASAP7_75t_SL g638 ( 
.A(n_604),
.Y(n_638)
);

AOI21x1_ASAP7_75t_SL g639 ( 
.A1(n_582),
.A2(n_542),
.B(n_26),
.Y(n_639)
);

AOI21xp5_ASAP7_75t_L g640 ( 
.A1(n_576),
.A2(n_114),
.B(n_135),
.Y(n_640)
);

NAND2xp5_ASAP7_75t_L g641 ( 
.A(n_582),
.B(n_542),
.Y(n_641)
);

OAI22xp5_ASAP7_75t_L g642 ( 
.A1(n_574),
.A2(n_25),
.B1(n_27),
.B2(n_43),
.Y(n_642)
);

INVx1_ASAP7_75t_SL g643 ( 
.A(n_595),
.Y(n_643)
);

O2A1O1Ixp5_ASAP7_75t_L g644 ( 
.A1(n_592),
.A2(n_605),
.B(n_599),
.C(n_609),
.Y(n_644)
);

OA21x2_ASAP7_75t_L g645 ( 
.A1(n_610),
.A2(n_25),
.B(n_27),
.Y(n_645)
);

AND2x2_ASAP7_75t_L g646 ( 
.A(n_612),
.B(n_134),
.Y(n_646)
);

AND2x4_ASAP7_75t_L g647 ( 
.A(n_577),
.B(n_44),
.Y(n_647)
);

BUFx6f_ASAP7_75t_L g648 ( 
.A(n_577),
.Y(n_648)
);

OA21x2_ASAP7_75t_L g649 ( 
.A1(n_585),
.A2(n_46),
.B(n_50),
.Y(n_649)
);

AND2x4_ASAP7_75t_L g650 ( 
.A(n_595),
.B(n_591),
.Y(n_650)
);

INVx1_ASAP7_75t_L g651 ( 
.A(n_628),
.Y(n_651)
);

INVx2_ASAP7_75t_L g652 ( 
.A(n_615),
.Y(n_652)
);

INVx2_ASAP7_75t_L g653 ( 
.A(n_617),
.Y(n_653)
);

OR2x2_ASAP7_75t_L g654 ( 
.A(n_616),
.B(n_607),
.Y(n_654)
);

INVx1_ASAP7_75t_L g655 ( 
.A(n_628),
.Y(n_655)
);

OAI21xp5_ASAP7_75t_L g656 ( 
.A1(n_644),
.A2(n_580),
.B(n_591),
.Y(n_656)
);

INVx3_ASAP7_75t_L g657 ( 
.A(n_635),
.Y(n_657)
);

BUFx6f_ASAP7_75t_L g658 ( 
.A(n_635),
.Y(n_658)
);

AND2x4_ASAP7_75t_L g659 ( 
.A(n_631),
.B(n_607),
.Y(n_659)
);

HB1xp67_ASAP7_75t_L g660 ( 
.A(n_613),
.Y(n_660)
);

INVx1_ASAP7_75t_L g661 ( 
.A(n_637),
.Y(n_661)
);

OA21x2_ASAP7_75t_L g662 ( 
.A1(n_637),
.A2(n_585),
.B(n_586),
.Y(n_662)
);

INVx2_ASAP7_75t_L g663 ( 
.A(n_617),
.Y(n_663)
);

INVx1_ASAP7_75t_L g664 ( 
.A(n_629),
.Y(n_664)
);

INVx1_ASAP7_75t_L g665 ( 
.A(n_623),
.Y(n_665)
);

INVx4_ASAP7_75t_SL g666 ( 
.A(n_629),
.Y(n_666)
);

NOR2xp33_ASAP7_75t_L g667 ( 
.A(n_641),
.B(n_51),
.Y(n_667)
);

INVx1_ASAP7_75t_L g668 ( 
.A(n_623),
.Y(n_668)
);

AND2x2_ASAP7_75t_L g669 ( 
.A(n_636),
.B(n_607),
.Y(n_669)
);

INVx1_ASAP7_75t_L g670 ( 
.A(n_627),
.Y(n_670)
);

INVx1_ASAP7_75t_L g671 ( 
.A(n_636),
.Y(n_671)
);

INVx2_ASAP7_75t_L g672 ( 
.A(n_635),
.Y(n_672)
);

INVx1_ASAP7_75t_L g673 ( 
.A(n_631),
.Y(n_673)
);

AND2x4_ASAP7_75t_L g674 ( 
.A(n_650),
.B(n_607),
.Y(n_674)
);

AND2x2_ASAP7_75t_L g675 ( 
.A(n_632),
.B(n_607),
.Y(n_675)
);

OR2x2_ASAP7_75t_L g676 ( 
.A(n_616),
.B(n_588),
.Y(n_676)
);

OR2x6_ASAP7_75t_L g677 ( 
.A(n_619),
.B(n_586),
.Y(n_677)
);

CKINVDCx20_ASAP7_75t_R g678 ( 
.A(n_638),
.Y(n_678)
);

AND2x2_ASAP7_75t_L g679 ( 
.A(n_632),
.B(n_588),
.Y(n_679)
);

NAND2xp5_ASAP7_75t_L g680 ( 
.A(n_626),
.B(n_588),
.Y(n_680)
);

INVx1_ASAP7_75t_L g681 ( 
.A(n_661),
.Y(n_681)
);

INVx2_ASAP7_75t_SL g682 ( 
.A(n_658),
.Y(n_682)
);

NOR2x1_ASAP7_75t_L g683 ( 
.A(n_673),
.B(n_619),
.Y(n_683)
);

AND2x2_ASAP7_75t_L g684 ( 
.A(n_666),
.B(n_622),
.Y(n_684)
);

AND2x2_ASAP7_75t_L g685 ( 
.A(n_666),
.B(n_622),
.Y(n_685)
);

AND2x2_ASAP7_75t_L g686 ( 
.A(n_666),
.B(n_627),
.Y(n_686)
);

BUFx2_ASAP7_75t_L g687 ( 
.A(n_651),
.Y(n_687)
);

BUFx6f_ASAP7_75t_L g688 ( 
.A(n_658),
.Y(n_688)
);

INVx2_ASAP7_75t_L g689 ( 
.A(n_661),
.Y(n_689)
);

INVx2_ASAP7_75t_L g690 ( 
.A(n_665),
.Y(n_690)
);

AND2x2_ASAP7_75t_L g691 ( 
.A(n_666),
.B(n_648),
.Y(n_691)
);

INVx1_ASAP7_75t_L g692 ( 
.A(n_651),
.Y(n_692)
);

AOI211xp5_ASAP7_75t_L g693 ( 
.A1(n_680),
.A2(n_642),
.B(n_633),
.C(n_620),
.Y(n_693)
);

AND2x2_ASAP7_75t_L g694 ( 
.A(n_664),
.B(n_648),
.Y(n_694)
);

INVx2_ASAP7_75t_L g695 ( 
.A(n_665),
.Y(n_695)
);

INVx1_ASAP7_75t_L g696 ( 
.A(n_655),
.Y(n_696)
);

INVx1_ASAP7_75t_L g697 ( 
.A(n_655),
.Y(n_697)
);

OR2x2_ASAP7_75t_L g698 ( 
.A(n_671),
.B(n_648),
.Y(n_698)
);

NOR2xp33_ASAP7_75t_L g699 ( 
.A(n_667),
.B(n_618),
.Y(n_699)
);

INVx2_ASAP7_75t_L g700 ( 
.A(n_668),
.Y(n_700)
);

INVx1_ASAP7_75t_L g701 ( 
.A(n_668),
.Y(n_701)
);

BUFx2_ASAP7_75t_L g702 ( 
.A(n_658),
.Y(n_702)
);

INVx2_ASAP7_75t_L g703 ( 
.A(n_670),
.Y(n_703)
);

AOI21xp5_ASAP7_75t_L g704 ( 
.A1(n_693),
.A2(n_656),
.B(n_677),
.Y(n_704)
);

AND2x2_ASAP7_75t_L g705 ( 
.A(n_694),
.B(n_669),
.Y(n_705)
);

OR2x2_ASAP7_75t_L g706 ( 
.A(n_687),
.B(n_654),
.Y(n_706)
);

OAI221xp5_ASAP7_75t_L g707 ( 
.A1(n_683),
.A2(n_677),
.B1(n_669),
.B2(n_660),
.C(n_654),
.Y(n_707)
);

INVx1_ASAP7_75t_L g708 ( 
.A(n_681),
.Y(n_708)
);

INVx3_ASAP7_75t_L g709 ( 
.A(n_688),
.Y(n_709)
);

NAND3xp33_ASAP7_75t_L g710 ( 
.A(n_683),
.B(n_677),
.C(n_624),
.Y(n_710)
);

BUFx2_ASAP7_75t_L g711 ( 
.A(n_702),
.Y(n_711)
);

AND2x4_ASAP7_75t_L g712 ( 
.A(n_691),
.B(n_672),
.Y(n_712)
);

AND2x2_ASAP7_75t_L g713 ( 
.A(n_694),
.B(n_675),
.Y(n_713)
);

NAND2xp5_ASAP7_75t_L g714 ( 
.A(n_698),
.B(n_675),
.Y(n_714)
);

BUFx3_ASAP7_75t_L g715 ( 
.A(n_702),
.Y(n_715)
);

INVx1_ASAP7_75t_L g716 ( 
.A(n_681),
.Y(n_716)
);

OAI22xp5_ASAP7_75t_L g717 ( 
.A1(n_699),
.A2(n_677),
.B1(n_618),
.B2(n_625),
.Y(n_717)
);

OAI21x1_ASAP7_75t_L g718 ( 
.A1(n_689),
.A2(n_676),
.B(n_662),
.Y(n_718)
);

AND2x6_ASAP7_75t_SL g719 ( 
.A(n_691),
.B(n_678),
.Y(n_719)
);

BUFx3_ASAP7_75t_L g720 ( 
.A(n_709),
.Y(n_720)
);

INVx4_ASAP7_75t_L g721 ( 
.A(n_719),
.Y(n_721)
);

INVx1_ASAP7_75t_L g722 ( 
.A(n_716),
.Y(n_722)
);

BUFx3_ASAP7_75t_L g723 ( 
.A(n_709),
.Y(n_723)
);

BUFx2_ASAP7_75t_L g724 ( 
.A(n_711),
.Y(n_724)
);

INVx3_ASAP7_75t_L g725 ( 
.A(n_718),
.Y(n_725)
);

INVx1_ASAP7_75t_L g726 ( 
.A(n_716),
.Y(n_726)
);

INVx2_ASAP7_75t_L g727 ( 
.A(n_718),
.Y(n_727)
);

BUFx2_ASAP7_75t_L g728 ( 
.A(n_711),
.Y(n_728)
);

NAND2xp5_ASAP7_75t_L g729 ( 
.A(n_704),
.B(n_698),
.Y(n_729)
);

OR2x2_ASAP7_75t_L g730 ( 
.A(n_706),
.B(n_687),
.Y(n_730)
);

INVx1_ASAP7_75t_L g731 ( 
.A(n_708),
.Y(n_731)
);

INVx2_ASAP7_75t_SL g732 ( 
.A(n_715),
.Y(n_732)
);

INVx1_ASAP7_75t_L g733 ( 
.A(n_706),
.Y(n_733)
);

NAND2xp5_ASAP7_75t_L g734 ( 
.A(n_733),
.B(n_705),
.Y(n_734)
);

AND2x2_ASAP7_75t_L g735 ( 
.A(n_721),
.B(n_705),
.Y(n_735)
);

AND2x2_ASAP7_75t_L g736 ( 
.A(n_721),
.B(n_713),
.Y(n_736)
);

AND2x2_ASAP7_75t_L g737 ( 
.A(n_721),
.B(n_713),
.Y(n_737)
);

INVx2_ASAP7_75t_SL g738 ( 
.A(n_732),
.Y(n_738)
);

NAND2xp5_ASAP7_75t_L g739 ( 
.A(n_729),
.B(n_714),
.Y(n_739)
);

NAND2xp5_ASAP7_75t_SL g740 ( 
.A(n_721),
.B(n_710),
.Y(n_740)
);

AND2x2_ASAP7_75t_L g741 ( 
.A(n_732),
.B(n_712),
.Y(n_741)
);

AND2x2_ASAP7_75t_L g742 ( 
.A(n_723),
.B(n_712),
.Y(n_742)
);

NAND2xp5_ASAP7_75t_L g743 ( 
.A(n_733),
.B(n_692),
.Y(n_743)
);

AOI22xp5_ASAP7_75t_L g744 ( 
.A1(n_740),
.A2(n_736),
.B1(n_735),
.B2(n_737),
.Y(n_744)
);

NAND2xp5_ASAP7_75t_L g745 ( 
.A(n_739),
.B(n_724),
.Y(n_745)
);

INVx2_ASAP7_75t_L g746 ( 
.A(n_742),
.Y(n_746)
);

INVx1_ASAP7_75t_SL g747 ( 
.A(n_738),
.Y(n_747)
);

AND2x2_ASAP7_75t_L g748 ( 
.A(n_741),
.B(n_723),
.Y(n_748)
);

AOI21xp5_ASAP7_75t_L g749 ( 
.A1(n_743),
.A2(n_707),
.B(n_734),
.Y(n_749)
);

AND2x2_ASAP7_75t_L g750 ( 
.A(n_748),
.B(n_734),
.Y(n_750)
);

OAI22xp5_ASAP7_75t_L g751 ( 
.A1(n_744),
.A2(n_728),
.B1(n_724),
.B2(n_717),
.Y(n_751)
);

HB1xp67_ASAP7_75t_L g752 ( 
.A(n_747),
.Y(n_752)
);

NOR2x1p5_ASAP7_75t_L g753 ( 
.A(n_745),
.B(n_720),
.Y(n_753)
);

INVx1_ASAP7_75t_L g754 ( 
.A(n_746),
.Y(n_754)
);

AOI22xp33_ASAP7_75t_L g755 ( 
.A1(n_751),
.A2(n_749),
.B1(n_727),
.B2(n_720),
.Y(n_755)
);

O2A1O1Ixp5_ASAP7_75t_L g756 ( 
.A1(n_754),
.A2(n_727),
.B(n_725),
.C(n_743),
.Y(n_756)
);

OAI21xp33_ASAP7_75t_SL g757 ( 
.A1(n_753),
.A2(n_725),
.B(n_730),
.Y(n_757)
);

AOI31xp33_ASAP7_75t_L g758 ( 
.A1(n_752),
.A2(n_750),
.A3(n_643),
.B(n_730),
.Y(n_758)
);

A2O1A1Ixp33_ASAP7_75t_L g759 ( 
.A1(n_752),
.A2(n_728),
.B(n_725),
.C(n_720),
.Y(n_759)
);

AOI21xp33_ASAP7_75t_SL g760 ( 
.A1(n_752),
.A2(n_709),
.B(n_625),
.Y(n_760)
);

OAI21xp33_ASAP7_75t_L g761 ( 
.A1(n_752),
.A2(n_725),
.B(n_731),
.Y(n_761)
);

NAND2xp5_ASAP7_75t_L g762 ( 
.A(n_752),
.B(n_731),
.Y(n_762)
);

AND2x4_ASAP7_75t_L g763 ( 
.A(n_762),
.B(n_722),
.Y(n_763)
);

AND2x2_ASAP7_75t_L g764 ( 
.A(n_755),
.B(n_712),
.Y(n_764)
);

INVx1_ASAP7_75t_L g765 ( 
.A(n_758),
.Y(n_765)
);

NAND2xp5_ASAP7_75t_L g766 ( 
.A(n_760),
.B(n_759),
.Y(n_766)
);

INVx2_ASAP7_75t_L g767 ( 
.A(n_756),
.Y(n_767)
);

AOI22xp5_ASAP7_75t_L g768 ( 
.A1(n_757),
.A2(n_761),
.B1(n_678),
.B2(n_722),
.Y(n_768)
);

CKINVDCx20_ASAP7_75t_R g769 ( 
.A(n_762),
.Y(n_769)
);

OAI211xp5_ASAP7_75t_SL g770 ( 
.A1(n_765),
.A2(n_640),
.B(n_726),
.C(n_621),
.Y(n_770)
);

OAI221xp5_ASAP7_75t_L g771 ( 
.A1(n_768),
.A2(n_715),
.B1(n_726),
.B2(n_682),
.C(n_688),
.Y(n_771)
);

NAND4xp25_ASAP7_75t_SL g772 ( 
.A(n_766),
.B(n_686),
.C(n_684),
.D(n_685),
.Y(n_772)
);

NAND4xp75_ASAP7_75t_L g773 ( 
.A(n_767),
.B(n_646),
.C(n_645),
.D(n_630),
.Y(n_773)
);

OAI22xp5_ASAP7_75t_L g774 ( 
.A1(n_769),
.A2(n_692),
.B1(n_696),
.B2(n_697),
.Y(n_774)
);

AOI211xp5_ASAP7_75t_L g775 ( 
.A1(n_771),
.A2(n_764),
.B(n_763),
.C(n_625),
.Y(n_775)
);

OAI211xp5_ASAP7_75t_L g776 ( 
.A1(n_770),
.A2(n_772),
.B(n_774),
.C(n_773),
.Y(n_776)
);

OAI221xp5_ASAP7_75t_L g777 ( 
.A1(n_771),
.A2(n_763),
.B1(n_682),
.B2(n_688),
.C(n_672),
.Y(n_777)
);

OAI22xp5_ASAP7_75t_SL g778 ( 
.A1(n_771),
.A2(n_634),
.B1(n_630),
.B2(n_645),
.Y(n_778)
);

OAI221xp5_ASAP7_75t_L g779 ( 
.A1(n_771),
.A2(n_688),
.B1(n_657),
.B2(n_630),
.C(n_645),
.Y(n_779)
);

AND2x2_ASAP7_75t_L g780 ( 
.A(n_775),
.B(n_686),
.Y(n_780)
);

INVx1_ASAP7_75t_SL g781 ( 
.A(n_778),
.Y(n_781)
);

NAND2xp5_ASAP7_75t_L g782 ( 
.A(n_776),
.B(n_696),
.Y(n_782)
);

NAND2xp5_ASAP7_75t_SL g783 ( 
.A(n_777),
.B(n_688),
.Y(n_783)
);

OAI21xp33_ASAP7_75t_SL g784 ( 
.A1(n_779),
.A2(n_684),
.B(n_685),
.Y(n_784)
);

OAI211xp5_ASAP7_75t_SL g785 ( 
.A1(n_781),
.A2(n_639),
.B(n_657),
.C(n_676),
.Y(n_785)
);

AOI22xp5_ASAP7_75t_L g786 ( 
.A1(n_780),
.A2(n_634),
.B1(n_647),
.B2(n_658),
.Y(n_786)
);

BUFx2_ASAP7_75t_L g787 ( 
.A(n_782),
.Y(n_787)
);

INVx1_ASAP7_75t_L g788 ( 
.A(n_783),
.Y(n_788)
);

INVx1_ASAP7_75t_L g789 ( 
.A(n_784),
.Y(n_789)
);

INVx2_ASAP7_75t_L g790 ( 
.A(n_780),
.Y(n_790)
);

HB1xp67_ASAP7_75t_L g791 ( 
.A(n_789),
.Y(n_791)
);

NOR3xp33_ASAP7_75t_L g792 ( 
.A(n_787),
.B(n_790),
.C(n_788),
.Y(n_792)
);

NAND4xp75_ASAP7_75t_L g793 ( 
.A(n_786),
.B(n_646),
.C(n_645),
.D(n_630),
.Y(n_793)
);

NAND3xp33_ASAP7_75t_L g794 ( 
.A(n_785),
.B(n_647),
.C(n_634),
.Y(n_794)
);

NOR4xp75_ASAP7_75t_SL g795 ( 
.A(n_789),
.B(n_583),
.C(n_584),
.D(n_589),
.Y(n_795)
);

INVx4_ASAP7_75t_L g796 ( 
.A(n_787),
.Y(n_796)
);

AOI221xp5_ASAP7_75t_L g797 ( 
.A1(n_789),
.A2(n_647),
.B1(n_583),
.B2(n_674),
.C(n_584),
.Y(n_797)
);

NOR2x1_ASAP7_75t_L g798 ( 
.A(n_796),
.B(n_584),
.Y(n_798)
);

INVx2_ASAP7_75t_L g799 ( 
.A(n_791),
.Y(n_799)
);

NOR4xp25_ASAP7_75t_L g800 ( 
.A(n_792),
.B(n_697),
.C(n_701),
.D(n_657),
.Y(n_800)
);

AND2x4_ASAP7_75t_L g801 ( 
.A(n_794),
.B(n_614),
.Y(n_801)
);

NAND2xp5_ASAP7_75t_L g802 ( 
.A(n_797),
.B(n_701),
.Y(n_802)
);

AND3x4_ASAP7_75t_L g803 ( 
.A(n_795),
.B(n_674),
.C(n_650),
.Y(n_803)
);

NOR3xp33_ASAP7_75t_L g804 ( 
.A(n_793),
.B(n_606),
.C(n_593),
.Y(n_804)
);

AND2x4_ASAP7_75t_L g805 ( 
.A(n_792),
.B(n_614),
.Y(n_805)
);

AND2x2_ASAP7_75t_L g806 ( 
.A(n_791),
.B(n_658),
.Y(n_806)
);

AND2x4_ASAP7_75t_L g807 ( 
.A(n_799),
.B(n_805),
.Y(n_807)
);

OAI322xp33_ASAP7_75t_L g808 ( 
.A1(n_806),
.A2(n_802),
.A3(n_800),
.B1(n_803),
.B2(n_801),
.C1(n_804),
.C2(n_798),
.Y(n_808)
);

OAI221xp5_ASAP7_75t_L g809 ( 
.A1(n_799),
.A2(n_649),
.B1(n_648),
.B2(n_695),
.C(n_690),
.Y(n_809)
);

AOI22xp5_ASAP7_75t_L g810 ( 
.A1(n_805),
.A2(n_674),
.B1(n_589),
.B2(n_649),
.Y(n_810)
);

OAI22xp5_ASAP7_75t_L g811 ( 
.A1(n_799),
.A2(n_689),
.B1(n_700),
.B2(n_695),
.Y(n_811)
);

OAI22xp33_ASAP7_75t_L g812 ( 
.A1(n_799),
.A2(n_649),
.B1(n_635),
.B2(n_648),
.Y(n_812)
);

OAI221xp5_ASAP7_75t_SL g813 ( 
.A1(n_799),
.A2(n_679),
.B1(n_700),
.B2(n_690),
.C(n_703),
.Y(n_813)
);

NAND3xp33_ASAP7_75t_SL g814 ( 
.A(n_799),
.B(n_52),
.C(n_53),
.Y(n_814)
);

INVx1_ASAP7_75t_L g815 ( 
.A(n_799),
.Y(n_815)
);

AND2x2_ASAP7_75t_L g816 ( 
.A(n_799),
.B(n_703),
.Y(n_816)
);

AOI221xp5_ASAP7_75t_L g817 ( 
.A1(n_799),
.A2(n_589),
.B1(n_650),
.B2(n_679),
.C(n_635),
.Y(n_817)
);

OAI22xp5_ASAP7_75t_SL g818 ( 
.A1(n_815),
.A2(n_649),
.B1(n_659),
.B2(n_662),
.Y(n_818)
);

INVxp67_ASAP7_75t_SL g819 ( 
.A(n_807),
.Y(n_819)
);

INVx2_ASAP7_75t_L g820 ( 
.A(n_816),
.Y(n_820)
);

HB1xp67_ASAP7_75t_L g821 ( 
.A(n_814),
.Y(n_821)
);

OAI22xp5_ASAP7_75t_L g822 ( 
.A1(n_813),
.A2(n_659),
.B1(n_670),
.B2(n_662),
.Y(n_822)
);

AOI22xp33_ASAP7_75t_SL g823 ( 
.A1(n_811),
.A2(n_659),
.B1(n_606),
.B2(n_593),
.Y(n_823)
);

NOR2xp33_ASAP7_75t_L g824 ( 
.A(n_808),
.B(n_54),
.Y(n_824)
);

NAND2xp5_ASAP7_75t_L g825 ( 
.A(n_817),
.B(n_55),
.Y(n_825)
);

OR2x2_ASAP7_75t_L g826 ( 
.A(n_810),
.B(n_662),
.Y(n_826)
);

AOI21xp5_ASAP7_75t_L g827 ( 
.A1(n_809),
.A2(n_576),
.B(n_59),
.Y(n_827)
);

AO22x2_ASAP7_75t_L g828 ( 
.A1(n_812),
.A2(n_57),
.B1(n_62),
.B2(n_63),
.Y(n_828)
);

OAI21xp5_ASAP7_75t_SL g829 ( 
.A1(n_815),
.A2(n_65),
.B(n_66),
.Y(n_829)
);

INVx1_ASAP7_75t_L g830 ( 
.A(n_815),
.Y(n_830)
);

OAI22xp5_ASAP7_75t_L g831 ( 
.A1(n_819),
.A2(n_830),
.B1(n_824),
.B2(n_821),
.Y(n_831)
);

INVx3_ASAP7_75t_SL g832 ( 
.A(n_820),
.Y(n_832)
);

AOI21xp33_ASAP7_75t_SL g833 ( 
.A1(n_825),
.A2(n_67),
.B(n_70),
.Y(n_833)
);

NOR2xp67_ASAP7_75t_L g834 ( 
.A(n_829),
.B(n_71),
.Y(n_834)
);

INVx2_ASAP7_75t_L g835 ( 
.A(n_828),
.Y(n_835)
);

OAI22xp5_ASAP7_75t_L g836 ( 
.A1(n_828),
.A2(n_663),
.B1(n_653),
.B2(n_652),
.Y(n_836)
);

INVx1_ASAP7_75t_L g837 ( 
.A(n_827),
.Y(n_837)
);

INVx1_ASAP7_75t_L g838 ( 
.A(n_826),
.Y(n_838)
);

OAI22xp5_ASAP7_75t_L g839 ( 
.A1(n_832),
.A2(n_822),
.B1(n_818),
.B2(n_823),
.Y(n_839)
);

INVx1_ASAP7_75t_L g840 ( 
.A(n_835),
.Y(n_840)
);

NAND2xp5_ASAP7_75t_L g841 ( 
.A(n_834),
.B(n_72),
.Y(n_841)
);

XNOR2xp5_ASAP7_75t_L g842 ( 
.A(n_831),
.B(n_74),
.Y(n_842)
);

INVx2_ASAP7_75t_L g843 ( 
.A(n_837),
.Y(n_843)
);

BUFx2_ASAP7_75t_L g844 ( 
.A(n_838),
.Y(n_844)
);

INVx1_ASAP7_75t_L g845 ( 
.A(n_833),
.Y(n_845)
);

NAND2xp5_ASAP7_75t_L g846 ( 
.A(n_844),
.B(n_836),
.Y(n_846)
);

INVx1_ASAP7_75t_SL g847 ( 
.A(n_841),
.Y(n_847)
);

CKINVDCx20_ASAP7_75t_R g848 ( 
.A(n_845),
.Y(n_848)
);

AOI21xp5_ASAP7_75t_L g849 ( 
.A1(n_846),
.A2(n_842),
.B(n_840),
.Y(n_849)
);

AOI22x1_ASAP7_75t_L g850 ( 
.A1(n_849),
.A2(n_843),
.B1(n_847),
.B2(n_848),
.Y(n_850)
);

AOI22x1_ASAP7_75t_L g851 ( 
.A1(n_850),
.A2(n_839),
.B1(n_78),
.B2(n_80),
.Y(n_851)
);

AOI221xp5_ASAP7_75t_L g852 ( 
.A1(n_851),
.A2(n_77),
.B1(n_106),
.B2(n_108),
.C(n_116),
.Y(n_852)
);

AOI211xp5_ASAP7_75t_L g853 ( 
.A1(n_852),
.A2(n_119),
.B(n_121),
.C(n_123),
.Y(n_853)
);


endmodule