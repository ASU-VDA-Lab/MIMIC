module fake_jpeg_20340_n_77 (n_3, n_2, n_1, n_0, n_4, n_8, n_6, n_5, n_7, n_77);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_8;
input n_6;
input n_5;
input n_7;

output n_77;

wire n_10;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_59;
wire n_65;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_28;
wire n_38;
wire n_26;
wire n_74;
wire n_31;
wire n_29;
wire n_50;
wire n_15;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_69;
wire n_27;
wire n_40;
wire n_71;
wire n_30;
wire n_24;
wire n_44;
wire n_17;
wire n_25;
wire n_75;
wire n_37;
wire n_70;
wire n_66;
wire n_61;
wire n_45;
wire n_18;
wire n_20;
wire n_68;
wire n_52;
wire n_58;
wire n_41;
wire n_60;
wire n_63;
wire n_34;
wire n_39;
wire n_72;
wire n_11;
wire n_56;
wire n_12;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_22;
wire n_35;
wire n_48;
wire n_46;
wire n_9;
wire n_36;
wire n_62;
wire n_43;
wire n_32;

NOR2xp33_ASAP7_75t_L g9 ( 
.A(n_4),
.B(n_0),
.Y(n_9)
);

CKINVDCx20_ASAP7_75t_R g10 ( 
.A(n_1),
.Y(n_10)
);

BUFx12_ASAP7_75t_L g11 ( 
.A(n_1),
.Y(n_11)
);

BUFx12f_ASAP7_75t_L g12 ( 
.A(n_3),
.Y(n_12)
);

BUFx12_ASAP7_75t_L g13 ( 
.A(n_2),
.Y(n_13)
);

CKINVDCx20_ASAP7_75t_R g14 ( 
.A(n_1),
.Y(n_14)
);

BUFx4f_ASAP7_75t_L g15 ( 
.A(n_5),
.Y(n_15)
);

BUFx12f_ASAP7_75t_L g16 ( 
.A(n_3),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_2),
.Y(n_17)
);

AND2x2_ASAP7_75t_L g18 ( 
.A(n_12),
.B(n_0),
.Y(n_18)
);

AND2x2_ASAP7_75t_L g25 ( 
.A(n_18),
.B(n_16),
.Y(n_25)
);

INVx8_ASAP7_75t_L g19 ( 
.A(n_12),
.Y(n_19)
);

INVx5_ASAP7_75t_L g29 ( 
.A(n_19),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_12),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_20),
.Y(n_28)
);

INVx5_ASAP7_75t_L g21 ( 
.A(n_16),
.Y(n_21)
);

NOR2xp33_ASAP7_75t_L g27 ( 
.A(n_21),
.B(n_22),
.Y(n_27)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_17),
.Y(n_22)
);

INVx2_ASAP7_75t_L g23 ( 
.A(n_15),
.Y(n_23)
);

BUFx12f_ASAP7_75t_L g26 ( 
.A(n_23),
.Y(n_26)
);

NAND2xp5_ASAP7_75t_L g24 ( 
.A(n_18),
.B(n_15),
.Y(n_24)
);

XNOR2xp5_ASAP7_75t_L g30 ( 
.A(n_24),
.B(n_18),
.Y(n_30)
);

AND2x2_ASAP7_75t_L g37 ( 
.A(n_25),
.B(n_16),
.Y(n_37)
);

AND2x2_ASAP7_75t_L g44 ( 
.A(n_30),
.B(n_31),
.Y(n_44)
);

INVx2_ASAP7_75t_R g31 ( 
.A(n_27),
.Y(n_31)
);

NOR2xp33_ASAP7_75t_L g32 ( 
.A(n_24),
.B(n_9),
.Y(n_32)
);

NAND2xp5_ASAP7_75t_L g47 ( 
.A(n_32),
.B(n_37),
.Y(n_47)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_28),
.Y(n_33)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_33),
.Y(n_48)
);

AOI22xp5_ASAP7_75t_L g34 ( 
.A1(n_25),
.A2(n_23),
.B1(n_22),
.B2(n_19),
.Y(n_34)
);

OAI22xp5_ASAP7_75t_SL g46 ( 
.A1(n_34),
.A2(n_36),
.B1(n_14),
.B2(n_20),
.Y(n_46)
);

INVx2_ASAP7_75t_SL g35 ( 
.A(n_29),
.Y(n_35)
);

BUFx5_ASAP7_75t_L g43 ( 
.A(n_35),
.Y(n_43)
);

AOI22xp5_ASAP7_75t_L g36 ( 
.A1(n_26),
.A2(n_19),
.B1(n_21),
.B2(n_17),
.Y(n_36)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_28),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_SL g45 ( 
.A(n_38),
.B(n_39),
.Y(n_45)
);

INVx2_ASAP7_75t_L g39 ( 
.A(n_26),
.Y(n_39)
);

XOR2xp5_ASAP7_75t_SL g40 ( 
.A(n_30),
.B(n_37),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_40),
.B(n_41),
.Y(n_56)
);

OR2x4_ASAP7_75t_L g41 ( 
.A(n_31),
.B(n_26),
.Y(n_41)
);

AOI22xp5_ASAP7_75t_L g42 ( 
.A1(n_34),
.A2(n_21),
.B1(n_29),
.B2(n_10),
.Y(n_42)
);

NAND2xp5_ASAP7_75t_L g50 ( 
.A(n_42),
.B(n_46),
.Y(n_50)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_48),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_L g59 ( 
.A(n_49),
.B(n_52),
.Y(n_59)
);

MAJIxp5_ASAP7_75t_L g51 ( 
.A(n_40),
.B(n_36),
.C(n_20),
.Y(n_51)
);

MAJIxp5_ASAP7_75t_L g57 ( 
.A(n_51),
.B(n_41),
.C(n_47),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_L g52 ( 
.A(n_44),
.B(n_15),
.Y(n_52)
);

INVxp67_ASAP7_75t_L g53 ( 
.A(n_45),
.Y(n_53)
);

INVxp67_ASAP7_75t_L g61 ( 
.A(n_53),
.Y(n_61)
);

CKINVDCx16_ASAP7_75t_R g54 ( 
.A(n_42),
.Y(n_54)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_54),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_L g55 ( 
.A(n_44),
.B(n_0),
.Y(n_55)
);

OAI321xp33_ASAP7_75t_L g58 ( 
.A1(n_55),
.A2(n_13),
.A3(n_11),
.B1(n_43),
.B2(n_6),
.C(n_7),
.Y(n_58)
);

XOR2xp5_ASAP7_75t_L g66 ( 
.A(n_57),
.B(n_11),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_58),
.B(n_51),
.Y(n_64)
);

AOI22xp5_ASAP7_75t_L g60 ( 
.A1(n_50),
.A2(n_35),
.B1(n_43),
.B2(n_2),
.Y(n_60)
);

AOI22xp5_ASAP7_75t_L g63 ( 
.A1(n_60),
.A2(n_53),
.B1(n_56),
.B2(n_6),
.Y(n_63)
);

CKINVDCx16_ASAP7_75t_R g68 ( 
.A(n_63),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_SL g69 ( 
.A(n_64),
.B(n_65),
.Y(n_69)
);

CKINVDCx20_ASAP7_75t_R g65 ( 
.A(n_59),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_L g67 ( 
.A(n_66),
.B(n_61),
.Y(n_67)
);

OAI21xp5_ASAP7_75t_L g71 ( 
.A1(n_67),
.A2(n_61),
.B(n_66),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_69),
.B(n_62),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_SL g73 ( 
.A(n_70),
.B(n_4),
.Y(n_73)
);

MAJIxp5_ASAP7_75t_L g72 ( 
.A(n_71),
.B(n_67),
.C(n_68),
.Y(n_72)
);

AOI21xp5_ASAP7_75t_L g74 ( 
.A1(n_72),
.A2(n_73),
.B(n_5),
.Y(n_74)
);

AOI21xp5_ASAP7_75t_L g75 ( 
.A1(n_74),
.A2(n_7),
.B(n_8),
.Y(n_75)
);

AOI22xp5_ASAP7_75t_L g76 ( 
.A1(n_75),
.A2(n_8),
.B1(n_13),
.B2(n_11),
.Y(n_76)
);

XOR2xp5_ASAP7_75t_L g77 ( 
.A(n_76),
.B(n_13),
.Y(n_77)
);


endmodule