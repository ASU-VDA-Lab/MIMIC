module fake_netlist_6_1216_n_1777 (n_52, n_16, n_1, n_91, n_119, n_46, n_146, n_163, n_18, n_21, n_147, n_154, n_88, n_3, n_98, n_113, n_39, n_63, n_73, n_4, n_148, n_138, n_22, n_161, n_68, n_28, n_50, n_158, n_49, n_7, n_83, n_5, n_101, n_144, n_127, n_125, n_153, n_77, n_156, n_149, n_152, n_106, n_92, n_145, n_42, n_133, n_96, n_8, n_90, n_160, n_24, n_105, n_131, n_54, n_132, n_102, n_0, n_87, n_32, n_66, n_85, n_99, n_78, n_84, n_130, n_164, n_100, n_129, n_13, n_121, n_11, n_137, n_17, n_23, n_142, n_20, n_143, n_2, n_19, n_47, n_62, n_29, n_155, n_75, n_109, n_150, n_122, n_45, n_34, n_140, n_70, n_120, n_37, n_15, n_67, n_33, n_82, n_27, n_38, n_110, n_151, n_61, n_112, n_81, n_59, n_76, n_36, n_26, n_124, n_55, n_126, n_94, n_97, n_108, n_58, n_116, n_64, n_117, n_118, n_48, n_65, n_25, n_40, n_93, n_80, n_141, n_135, n_139, n_41, n_134, n_114, n_86, n_104, n_95, n_9, n_107, n_10, n_71, n_74, n_6, n_14, n_123, n_136, n_72, n_89, n_103, n_111, n_60, n_159, n_157, n_162, n_35, n_115, n_12, n_69, n_128, n_30, n_79, n_43, n_31, n_57, n_53, n_51, n_44, n_56, n_1777);

input n_52;
input n_16;
input n_1;
input n_91;
input n_119;
input n_46;
input n_146;
input n_163;
input n_18;
input n_21;
input n_147;
input n_154;
input n_88;
input n_3;
input n_98;
input n_113;
input n_39;
input n_63;
input n_73;
input n_4;
input n_148;
input n_138;
input n_22;
input n_161;
input n_68;
input n_28;
input n_50;
input n_158;
input n_49;
input n_7;
input n_83;
input n_5;
input n_101;
input n_144;
input n_127;
input n_125;
input n_153;
input n_77;
input n_156;
input n_149;
input n_152;
input n_106;
input n_92;
input n_145;
input n_42;
input n_133;
input n_96;
input n_8;
input n_90;
input n_160;
input n_24;
input n_105;
input n_131;
input n_54;
input n_132;
input n_102;
input n_0;
input n_87;
input n_32;
input n_66;
input n_85;
input n_99;
input n_78;
input n_84;
input n_130;
input n_164;
input n_100;
input n_129;
input n_13;
input n_121;
input n_11;
input n_137;
input n_17;
input n_23;
input n_142;
input n_20;
input n_143;
input n_2;
input n_19;
input n_47;
input n_62;
input n_29;
input n_155;
input n_75;
input n_109;
input n_150;
input n_122;
input n_45;
input n_34;
input n_140;
input n_70;
input n_120;
input n_37;
input n_15;
input n_67;
input n_33;
input n_82;
input n_27;
input n_38;
input n_110;
input n_151;
input n_61;
input n_112;
input n_81;
input n_59;
input n_76;
input n_36;
input n_26;
input n_124;
input n_55;
input n_126;
input n_94;
input n_97;
input n_108;
input n_58;
input n_116;
input n_64;
input n_117;
input n_118;
input n_48;
input n_65;
input n_25;
input n_40;
input n_93;
input n_80;
input n_141;
input n_135;
input n_139;
input n_41;
input n_134;
input n_114;
input n_86;
input n_104;
input n_95;
input n_9;
input n_107;
input n_10;
input n_71;
input n_74;
input n_6;
input n_14;
input n_123;
input n_136;
input n_72;
input n_89;
input n_103;
input n_111;
input n_60;
input n_159;
input n_157;
input n_162;
input n_35;
input n_115;
input n_12;
input n_69;
input n_128;
input n_30;
input n_79;
input n_43;
input n_31;
input n_57;
input n_53;
input n_51;
input n_44;
input n_56;

output n_1777;

wire n_992;
wire n_1671;
wire n_801;
wire n_1613;
wire n_1234;
wire n_1458;
wire n_1199;
wire n_1674;
wire n_741;
wire n_1027;
wire n_1351;
wire n_625;
wire n_1189;
wire n_223;
wire n_1212;
wire n_226;
wire n_208;
wire n_726;
wire n_212;
wire n_700;
wire n_1307;
wire n_1038;
wire n_578;
wire n_1581;
wire n_1003;
wire n_365;
wire n_168;
wire n_1237;
wire n_1061;
wire n_1357;
wire n_783;
wire n_1738;
wire n_798;
wire n_188;
wire n_1575;
wire n_509;
wire n_1342;
wire n_245;
wire n_1209;
wire n_1348;
wire n_1387;
wire n_677;
wire n_1708;
wire n_805;
wire n_1151;
wire n_396;
wire n_1739;
wire n_350;
wire n_1380;
wire n_442;
wire n_480;
wire n_1402;
wire n_1691;
wire n_1688;
wire n_1009;
wire n_1743;
wire n_1160;
wire n_883;
wire n_1238;
wire n_1724;
wire n_1032;
wire n_1247;
wire n_1547;
wire n_1553;
wire n_893;
wire n_1099;
wire n_1264;
wire n_1192;
wire n_471;
wire n_424;
wire n_1700;
wire n_1555;
wire n_1415;
wire n_1370;
wire n_369;
wire n_287;
wire n_415;
wire n_830;
wire n_230;
wire n_461;
wire n_873;
wire n_383;
wire n_1285;
wire n_1371;
wire n_200;
wire n_447;
wire n_1172;
wire n_852;
wire n_229;
wire n_1590;
wire n_1532;
wire n_1393;
wire n_1517;
wire n_1704;
wire n_1078;
wire n_250;
wire n_544;
wire n_1711;
wire n_1140;
wire n_1444;
wire n_1670;
wire n_1603;
wire n_1579;
wire n_1263;
wire n_836;
wire n_375;
wire n_522;
wire n_1261;
wire n_945;
wire n_1649;
wire n_1511;
wire n_1143;
wire n_1422;
wire n_1232;
wire n_1772;
wire n_1572;
wire n_658;
wire n_616;
wire n_1119;
wire n_428;
wire n_1433;
wire n_1620;
wire n_1735;
wire n_1541;
wire n_1300;
wire n_641;
wire n_822;
wire n_693;
wire n_1313;
wire n_1056;
wire n_758;
wire n_516;
wire n_1455;
wire n_1163;
wire n_1180;
wire n_943;
wire n_1550;
wire n_491;
wire n_1591;
wire n_772;
wire n_1344;
wire n_666;
wire n_371;
wire n_940;
wire n_770;
wire n_567;
wire n_405;
wire n_213;
wire n_538;
wire n_1106;
wire n_886;
wire n_1471;
wire n_343;
wire n_953;
wire n_1094;
wire n_1345;
wire n_494;
wire n_539;
wire n_493;
wire n_454;
wire n_1421;
wire n_638;
wire n_1404;
wire n_1211;
wire n_381;
wire n_887;
wire n_1660;
wire n_1280;
wire n_713;
wire n_1400;
wire n_1467;
wire n_976;
wire n_224;
wire n_1445;
wire n_1526;
wire n_1560;
wire n_734;
wire n_1088;
wire n_196;
wire n_1231;
wire n_917;
wire n_574;
wire n_907;
wire n_1446;
wire n_659;
wire n_407;
wire n_913;
wire n_1658;
wire n_808;
wire n_867;
wire n_1230;
wire n_473;
wire n_1193;
wire n_1054;
wire n_559;
wire n_1333;
wire n_1648;
wire n_1644;
wire n_1558;
wire n_1732;
wire n_281;
wire n_551;
wire n_699;
wire n_564;
wire n_451;
wire n_824;
wire n_279;
wire n_686;
wire n_757;
wire n_594;
wire n_1641;
wire n_577;
wire n_166;
wire n_619;
wire n_1367;
wire n_1336;
wire n_521;
wire n_572;
wire n_395;
wire n_813;
wire n_1481;
wire n_323;
wire n_606;
wire n_1441;
wire n_818;
wire n_1123;
wire n_1309;
wire n_513;
wire n_645;
wire n_1381;
wire n_331;
wire n_1699;
wire n_916;
wire n_483;
wire n_608;
wire n_261;
wire n_630;
wire n_541;
wire n_512;
wire n_433;
wire n_792;
wire n_476;
wire n_1328;
wire n_219;
wire n_264;
wire n_263;
wire n_1162;
wire n_860;
wire n_1530;
wire n_788;
wire n_939;
wire n_1543;
wire n_821;
wire n_938;
wire n_1302;
wire n_1068;
wire n_1599;
wire n_329;
wire n_982;
wire n_549;
wire n_1762;
wire n_1075;
wire n_408;
wire n_932;
wire n_237;
wire n_1697;
wire n_243;
wire n_979;
wire n_905;
wire n_1680;
wire n_175;
wire n_322;
wire n_993;
wire n_689;
wire n_354;
wire n_1330;
wire n_1413;
wire n_1605;
wire n_1278;
wire n_547;
wire n_558;
wire n_1064;
wire n_1396;
wire n_634;
wire n_966;
wire n_764;
wire n_1663;
wire n_692;
wire n_733;
wire n_1233;
wire n_1289;
wire n_487;
wire n_241;
wire n_1107;
wire n_1014;
wire n_1290;
wire n_1703;
wire n_882;
wire n_1354;
wire n_586;
wire n_423;
wire n_1701;
wire n_318;
wire n_1111;
wire n_1713;
wire n_715;
wire n_1251;
wire n_1265;
wire n_1726;
wire n_530;
wire n_1563;
wire n_277;
wire n_618;
wire n_1297;
wire n_1662;
wire n_1312;
wire n_199;
wire n_1167;
wire n_1359;
wire n_674;
wire n_871;
wire n_922;
wire n_268;
wire n_1335;
wire n_1760;
wire n_210;
wire n_1069;
wire n_1664;
wire n_1722;
wire n_612;
wire n_178;
wire n_247;
wire n_1165;
wire n_355;
wire n_702;
wire n_347;
wire n_1175;
wire n_328;
wire n_1386;
wire n_429;
wire n_1747;
wire n_1012;
wire n_195;
wire n_780;
wire n_675;
wire n_903;
wire n_1540;
wire n_1504;
wire n_286;
wire n_254;
wire n_1655;
wire n_242;
wire n_835;
wire n_928;
wire n_1214;
wire n_690;
wire n_850;
wire n_1654;
wire n_816;
wire n_1157;
wire n_1750;
wire n_1462;
wire n_1188;
wire n_1752;
wire n_877;
wire n_604;
wire n_825;
wire n_728;
wire n_1063;
wire n_1588;
wire n_267;
wire n_1124;
wire n_1624;
wire n_515;
wire n_598;
wire n_696;
wire n_1515;
wire n_961;
wire n_437;
wire n_1082;
wire n_1317;
wire n_593;
wire n_514;
wire n_697;
wire n_687;
wire n_890;
wire n_637;
wire n_295;
wire n_701;
wire n_950;
wire n_388;
wire n_190;
wire n_484;
wire n_1709;
wire n_1757;
wire n_170;
wire n_891;
wire n_1412;
wire n_949;
wire n_1630;
wire n_678;
wire n_283;
wire n_507;
wire n_968;
wire n_909;
wire n_1369;
wire n_881;
wire n_1008;
wire n_760;
wire n_1546;
wire n_590;
wire n_362;
wire n_462;
wire n_1033;
wire n_1052;
wire n_1296;
wire n_304;
wire n_694;
wire n_1294;
wire n_1420;
wire n_1634;
wire n_297;
wire n_595;
wire n_627;
wire n_1767;
wire n_524;
wire n_1465;
wire n_342;
wire n_1044;
wire n_1712;
wire n_1391;
wire n_449;
wire n_1523;
wire n_1208;
wire n_1164;
wire n_1295;
wire n_1627;
wire n_1072;
wire n_1527;
wire n_1495;
wire n_1438;
wire n_495;
wire n_815;
wire n_1100;
wire n_585;
wire n_1487;
wire n_840;
wire n_874;
wire n_1756;
wire n_1128;
wire n_382;
wire n_673;
wire n_1071;
wire n_1067;
wire n_1565;
wire n_1493;
wire n_898;
wire n_255;
wire n_284;
wire n_865;
wire n_925;
wire n_1101;
wire n_1026;
wire n_289;
wire n_1364;
wire n_615;
wire n_1249;
wire n_1293;
wire n_1127;
wire n_1512;
wire n_1451;
wire n_320;
wire n_639;
wire n_963;
wire n_794;
wire n_727;
wire n_894;
wire n_685;
wire n_1765;
wire n_353;
wire n_605;
wire n_1514;
wire n_826;
wire n_1646;
wire n_872;
wire n_1139;
wire n_1714;
wire n_718;
wire n_1018;
wire n_1521;
wire n_1366;
wire n_542;
wire n_847;
wire n_644;
wire n_682;
wire n_851;
wire n_305;
wire n_996;
wire n_532;
wire n_173;
wire n_1308;
wire n_1376;
wire n_1513;
wire n_413;
wire n_791;
wire n_510;
wire n_837;
wire n_1488;
wire n_948;
wire n_704;
wire n_977;
wire n_1005;
wire n_536;
wire n_622;
wire n_1469;
wire n_1766;
wire n_1776;
wire n_581;
wire n_765;
wire n_432;
wire n_987;
wire n_1492;
wire n_1340;
wire n_1771;
wire n_631;
wire n_720;
wire n_842;
wire n_1707;
wire n_1432;
wire n_843;
wire n_656;
wire n_989;
wire n_1277;
wire n_797;
wire n_1473;
wire n_1723;
wire n_1246;
wire n_899;
wire n_189;
wire n_738;
wire n_1304;
wire n_1035;
wire n_294;
wire n_499;
wire n_1426;
wire n_705;
wire n_1004;
wire n_1176;
wire n_1529;
wire n_1022;
wire n_614;
wire n_529;
wire n_425;
wire n_684;
wire n_1431;
wire n_1615;
wire n_1474;
wire n_1571;
wire n_1577;
wire n_1181;
wire n_486;
wire n_947;
wire n_1117;
wire n_1087;
wire n_1448;
wire n_648;
wire n_657;
wire n_1049;
wire n_1666;
wire n_1505;
wire n_803;
wire n_290;
wire n_1717;
wire n_926;
wire n_927;
wire n_919;
wire n_1698;
wire n_478;
wire n_929;
wire n_1228;
wire n_417;
wire n_446;
wire n_1568;
wire n_1490;
wire n_777;
wire n_1299;
wire n_272;
wire n_526;
wire n_1183;
wire n_1436;
wire n_1384;
wire n_293;
wire n_458;
wire n_1070;
wire n_998;
wire n_717;
wire n_1665;
wire n_1383;
wire n_1178;
wire n_1424;
wire n_1073;
wire n_1000;
wire n_796;
wire n_252;
wire n_1195;
wire n_1626;
wire n_1507;
wire n_184;
wire n_552;
wire n_1358;
wire n_1388;
wire n_216;
wire n_912;
wire n_1519;
wire n_745;
wire n_1284;
wire n_1604;
wire n_1142;
wire n_716;
wire n_1475;
wire n_623;
wire n_1048;
wire n_1201;
wire n_1398;
wire n_884;
wire n_1774;
wire n_1395;
wire n_731;
wire n_1502;
wire n_1659;
wire n_755;
wire n_931;
wire n_1021;
wire n_474;
wire n_527;
wire n_683;
wire n_811;
wire n_1207;
wire n_312;
wire n_1368;
wire n_1418;
wire n_958;
wire n_292;
wire n_1250;
wire n_1137;
wire n_880;
wire n_889;
wire n_1478;
wire n_589;
wire n_1310;
wire n_819;
wire n_1363;
wire n_1334;
wire n_767;
wire n_1314;
wire n_600;
wire n_964;
wire n_831;
wire n_477;
wire n_954;
wire n_864;
wire n_1110;
wire n_1410;
wire n_399;
wire n_1440;
wire n_1382;
wire n_1534;
wire n_1564;
wire n_1736;
wire n_211;
wire n_1483;
wire n_1372;
wire n_231;
wire n_1457;
wire n_505;
wire n_1719;
wire n_319;
wire n_1339;
wire n_537;
wire n_1427;
wire n_311;
wire n_1466;
wire n_403;
wire n_1080;
wire n_723;
wire n_596;
wire n_546;
wire n_562;
wire n_1141;
wire n_1268;
wire n_386;
wire n_1769;
wire n_1220;
wire n_556;
wire n_1755;
wire n_1602;
wire n_1136;
wire n_1125;
wire n_970;
wire n_642;
wire n_995;
wire n_276;
wire n_1159;
wire n_1092;
wire n_441;
wire n_221;
wire n_1060;
wire n_444;
wire n_1252;
wire n_1223;
wire n_303;
wire n_511;
wire n_193;
wire n_1286;
wire n_1773;
wire n_1775;
wire n_1053;
wire n_416;
wire n_1681;
wire n_520;
wire n_418;
wire n_1093;
wire n_1533;
wire n_1597;
wire n_266;
wire n_296;
wire n_775;
wire n_651;
wire n_1153;
wire n_439;
wire n_1618;
wire n_217;
wire n_518;
wire n_1531;
wire n_1185;
wire n_453;
wire n_215;
wire n_1745;
wire n_914;
wire n_759;
wire n_426;
wire n_317;
wire n_1653;
wire n_1679;
wire n_1625;
wire n_1453;
wire n_488;
wire n_497;
wire n_773;
wire n_920;
wire n_1374;
wire n_1315;
wire n_1647;
wire n_1224;
wire n_1614;
wire n_1459;
wire n_1135;
wire n_1169;
wire n_1179;
wire n_401;
wire n_324;
wire n_1617;
wire n_335;
wire n_1470;
wire n_463;
wire n_1243;
wire n_848;
wire n_301;
wire n_274;
wire n_1096;
wire n_1091;
wire n_1580;
wire n_1425;
wire n_1267;
wire n_1281;
wire n_983;
wire n_427;
wire n_1520;
wire n_496;
wire n_906;
wire n_1390;
wire n_688;
wire n_1077;
wire n_1733;
wire n_1419;
wire n_351;
wire n_259;
wire n_1731;
wire n_177;
wire n_1636;
wire n_1437;
wire n_1645;
wire n_385;
wire n_1687;
wire n_1439;
wire n_1323;
wire n_858;
wire n_1331;
wire n_736;
wire n_613;
wire n_501;
wire n_956;
wire n_960;
wire n_663;
wire n_856;
wire n_379;
wire n_778;
wire n_1668;
wire n_1134;
wire n_410;
wire n_1129;
wire n_554;
wire n_602;
wire n_1696;
wire n_1594;
wire n_664;
wire n_171;
wire n_1764;
wire n_169;
wire n_1429;
wire n_1610;
wire n_435;
wire n_793;
wire n_326;
wire n_587;
wire n_1593;
wire n_580;
wire n_762;
wire n_1030;
wire n_1202;
wire n_465;
wire n_1635;
wire n_1079;
wire n_341;
wire n_1744;
wire n_828;
wire n_607;
wire n_316;
wire n_419;
wire n_1551;
wire n_1103;
wire n_1203;
wire n_820;
wire n_951;
wire n_725;
wire n_952;
wire n_999;
wire n_358;
wire n_1254;
wire n_186;
wire n_368;
wire n_575;
wire n_994;
wire n_1508;
wire n_732;
wire n_974;
wire n_392;
wire n_724;
wire n_1020;
wire n_1042;
wire n_628;
wire n_1273;
wire n_1434;
wire n_1573;
wire n_1728;
wire n_557;
wire n_349;
wire n_617;
wire n_845;
wire n_807;
wire n_1036;
wire n_1138;
wire n_1661;
wire n_1275;
wire n_485;
wire n_1549;
wire n_443;
wire n_1510;
wire n_892;
wire n_768;
wire n_421;
wire n_1468;
wire n_238;
wire n_1095;
wire n_1595;
wire n_202;
wire n_1718;
wire n_1749;
wire n_1683;
wire n_597;
wire n_280;
wire n_1270;
wire n_1187;
wire n_610;
wire n_1403;
wire n_1669;
wire n_1024;
wire n_1768;
wire n_198;
wire n_179;
wire n_248;
wire n_517;
wire n_1667;
wire n_667;
wire n_1206;
wire n_621;
wire n_1037;
wire n_1397;
wire n_1279;
wire n_1115;
wire n_750;
wire n_901;
wire n_1499;
wire n_468;
wire n_923;
wire n_504;
wire n_1409;
wire n_1639;
wire n_1623;
wire n_183;
wire n_1015;
wire n_1503;
wire n_466;
wire n_1057;
wire n_603;
wire n_991;
wire n_1657;
wire n_235;
wire n_1126;
wire n_340;
wire n_710;
wire n_1108;
wire n_1182;
wire n_1298;
wire n_1611;
wire n_785;
wire n_746;
wire n_609;
wire n_1601;
wire n_1686;
wire n_167;
wire n_1356;
wire n_1589;
wire n_1740;
wire n_1497;
wire n_1168;
wire n_1216;
wire n_1320;
wire n_1430;
wire n_1316;
wire n_1287;
wire n_1452;
wire n_1622;
wire n_1586;
wire n_302;
wire n_1694;
wire n_380;
wire n_1535;
wire n_1596;
wire n_1190;
wire n_1734;
wire n_397;
wire n_1262;
wire n_218;
wire n_1213;
wire n_1350;
wire n_1673;
wire n_1715;
wire n_172;
wire n_1443;
wire n_1272;
wire n_239;
wire n_782;
wire n_1539;
wire n_490;
wire n_220;
wire n_809;
wire n_1043;
wire n_1608;
wire n_986;
wire n_1472;
wire n_1081;
wire n_402;
wire n_352;
wire n_1692;
wire n_800;
wire n_1084;
wire n_1171;
wire n_460;
wire n_1361;
wire n_1491;
wire n_662;
wire n_374;
wire n_1152;
wire n_1705;
wire n_450;
wire n_1684;
wire n_921;
wire n_1346;
wire n_711;
wire n_1642;
wire n_579;
wire n_1352;
wire n_937;
wire n_1682;
wire n_370;
wire n_1695;
wire n_650;
wire n_1046;
wire n_1145;
wire n_330;
wire n_1121;
wire n_1102;
wire n_972;
wire n_1405;
wire n_258;
wire n_1406;
wire n_456;
wire n_1332;
wire n_260;
wire n_313;
wire n_624;
wire n_962;
wire n_1041;
wire n_565;
wire n_356;
wire n_1569;
wire n_936;
wire n_1288;
wire n_1186;
wire n_1062;
wire n_885;
wire n_896;
wire n_654;
wire n_411;
wire n_1222;
wire n_599;
wire n_776;
wire n_321;
wire n_227;
wire n_1720;
wire n_204;
wire n_482;
wire n_934;
wire n_1637;
wire n_1407;
wire n_420;
wire n_1341;
wire n_394;
wire n_1456;
wire n_1489;
wire n_942;
wire n_1524;
wire n_543;
wire n_1496;
wire n_1271;
wire n_1545;
wire n_1355;
wire n_1225;
wire n_1544;
wire n_1485;
wire n_325;
wire n_1640;
wire n_804;
wire n_464;
wire n_533;
wire n_806;
wire n_959;
wire n_879;
wire n_584;
wire n_244;
wire n_1343;
wire n_1522;
wire n_548;
wire n_282;
wire n_1676;
wire n_833;
wire n_1567;
wire n_523;
wire n_1319;
wire n_707;
wire n_345;
wire n_799;
wire n_1548;
wire n_1155;
wire n_273;
wire n_1633;
wire n_787;
wire n_1416;
wire n_1528;
wire n_1146;
wire n_1086;
wire n_1066;
wire n_1282;
wire n_550;
wire n_275;
wire n_652;
wire n_560;
wire n_1484;
wire n_1241;
wire n_1321;
wire n_1672;
wire n_569;
wire n_1758;
wire n_737;
wire n_1318;
wire n_1235;
wire n_1229;
wire n_306;
wire n_1292;
wire n_1373;
wire n_346;
wire n_1029;
wire n_1447;
wire n_790;
wire n_1706;
wire n_1498;
wire n_1210;
wire n_299;
wire n_1248;
wire n_1556;
wire n_902;
wire n_333;
wire n_1047;
wire n_1385;
wire n_431;
wire n_459;
wire n_1269;
wire n_502;
wire n_672;
wire n_1257;
wire n_1751;
wire n_285;
wire n_1375;
wire n_655;
wire n_706;
wire n_1045;
wire n_1650;
wire n_786;
wire n_1236;
wire n_1559;
wire n_1725;
wire n_834;
wire n_743;
wire n_766;
wire n_430;
wire n_1741;
wire n_1325;
wire n_1002;
wire n_1746;
wire n_545;
wire n_489;
wire n_1727;
wire n_251;
wire n_1019;
wire n_636;
wire n_729;
wire n_876;
wire n_774;
wire n_1337;
wire n_660;
wire n_438;
wire n_1477;
wire n_1360;
wire n_1200;
wire n_479;
wire n_1607;
wire n_1353;
wire n_1454;
wire n_869;
wire n_1154;
wire n_1113;
wire n_1600;
wire n_646;
wire n_528;
wire n_391;
wire n_1098;
wire n_1329;
wire n_817;
wire n_262;
wire n_187;
wire n_897;
wire n_846;
wire n_841;
wire n_1476;
wire n_1001;
wire n_508;
wire n_1050;
wire n_1411;
wire n_1463;
wire n_1177;
wire n_332;
wire n_1150;
wire n_1742;
wire n_1562;
wire n_1690;
wire n_398;
wire n_1191;
wire n_566;
wire n_1023;
wire n_1118;
wire n_1076;
wire n_194;
wire n_1007;
wire n_1378;
wire n_855;
wire n_1592;
wire n_1759;
wire n_1631;
wire n_591;
wire n_1377;
wire n_256;
wire n_853;
wire n_440;
wire n_695;
wire n_1542;
wire n_875;
wire n_209;
wire n_367;
wire n_680;
wire n_1678;
wire n_661;
wire n_1716;
wire n_278;
wire n_1256;
wire n_671;
wire n_933;
wire n_740;
wire n_703;
wire n_978;
wire n_384;
wire n_1291;
wire n_1217;
wire n_751;
wire n_749;
wire n_310;
wire n_1628;
wire n_1324;
wire n_1399;
wire n_1435;
wire n_969;
wire n_988;
wire n_1065;
wire n_1401;
wire n_1255;
wire n_568;
wire n_1516;
wire n_1536;
wire n_180;
wire n_1204;
wire n_823;
wire n_1132;
wire n_643;
wire n_233;
wire n_698;
wire n_1074;
wire n_1394;
wire n_1327;
wire n_1326;
wire n_739;
wire n_400;
wire n_955;
wire n_337;
wire n_1379;
wire n_214;
wire n_246;
wire n_1338;
wire n_1097;
wire n_935;
wire n_781;
wire n_789;
wire n_1554;
wire n_1130;
wire n_181;
wire n_182;
wire n_573;
wire n_769;
wire n_676;
wire n_327;
wire n_1120;
wire n_832;
wire n_1583;
wire n_1730;
wire n_555;
wire n_389;
wire n_814;
wire n_1643;
wire n_1729;
wire n_669;
wire n_176;
wire n_300;
wire n_222;
wire n_747;
wire n_1389;
wire n_1105;
wire n_721;
wire n_1461;
wire n_742;
wire n_535;
wire n_691;
wire n_372;
wire n_314;
wire n_1408;
wire n_378;
wire n_1196;
wire n_377;
wire n_1598;
wire n_863;
wire n_601;
wire n_338;
wire n_1283;
wire n_918;
wire n_748;
wire n_506;
wire n_1114;
wire n_763;
wire n_1147;
wire n_360;
wire n_1754;
wire n_1506;
wire n_1652;
wire n_957;
wire n_895;
wire n_866;
wire n_1227;
wire n_191;
wire n_387;
wire n_452;
wire n_744;
wire n_971;
wire n_946;
wire n_344;
wire n_761;
wire n_1303;
wire n_1205;
wire n_1258;
wire n_1392;
wire n_174;
wire n_1173;
wire n_525;
wire n_1677;
wire n_1116;
wire n_611;
wire n_1570;
wire n_1702;
wire n_1219;
wire n_1689;
wire n_1174;
wire n_1016;
wire n_1347;
wire n_795;
wire n_1501;
wire n_1221;
wire n_1245;
wire n_838;
wire n_647;
wire n_197;
wire n_844;
wire n_448;
wire n_1017;
wire n_1083;
wire n_445;
wire n_1561;
wire n_930;
wire n_888;
wire n_1112;
wire n_234;
wire n_910;
wire n_1656;
wire n_1721;
wire n_1460;
wire n_911;
wire n_1464;
wire n_236;
wire n_653;
wire n_1737;
wire n_1414;
wire n_752;
wire n_908;
wire n_944;
wire n_576;
wire n_1028;
wire n_472;
wire n_270;
wire n_414;
wire n_563;
wire n_1011;
wire n_1566;
wire n_1215;
wire n_839;
wire n_708;
wire n_668;
wire n_626;
wire n_990;
wire n_1500;
wire n_779;
wire n_1537;
wire n_1104;
wire n_854;
wire n_1058;
wire n_498;
wire n_1122;
wire n_870;
wire n_904;
wire n_1253;
wire n_709;
wire n_1266;
wire n_366;
wire n_1509;
wire n_1693;
wire n_1109;
wire n_185;
wire n_712;
wire n_348;
wire n_1276;
wire n_376;
wire n_390;
wire n_1148;
wire n_334;
wire n_1161;
wire n_1085;
wire n_232;
wire n_1239;
wire n_771;
wire n_1584;
wire n_470;
wire n_475;
wire n_924;
wire n_298;
wire n_1582;
wire n_492;
wire n_1149;
wire n_265;
wire n_1184;
wire n_228;
wire n_719;
wire n_1525;
wire n_455;
wire n_1585;
wire n_363;
wire n_1090;
wire n_592;
wire n_1518;
wire n_829;
wire n_1156;
wire n_1362;
wire n_393;
wire n_984;
wire n_503;
wire n_1450;
wire n_1638;
wire n_868;
wire n_570;
wire n_859;
wire n_406;
wire n_735;
wire n_1770;
wire n_878;
wire n_620;
wire n_519;
wire n_307;
wire n_469;
wire n_1218;
wire n_500;
wire n_1482;
wire n_981;
wire n_714;
wire n_1349;
wire n_291;
wire n_1144;
wire n_357;
wire n_985;
wire n_481;
wire n_997;
wire n_1710;
wire n_1301;
wire n_802;
wire n_561;
wire n_980;
wire n_1306;
wire n_1651;
wire n_1198;
wire n_1609;
wire n_436;
wire n_409;
wire n_1244;
wire n_1685;
wire n_1763;
wire n_1574;
wire n_240;
wire n_756;
wire n_1619;
wire n_1606;
wire n_810;
wire n_1133;
wire n_635;
wire n_1194;
wire n_1051;
wire n_253;
wire n_1552;
wire n_583;
wire n_249;
wire n_201;
wire n_1039;
wire n_1442;
wire n_1034;
wire n_1480;
wire n_1158;
wire n_754;
wire n_941;
wire n_975;
wire n_1031;
wire n_1305;
wire n_553;
wire n_849;
wire n_753;
wire n_1753;
wire n_467;
wire n_269;
wire n_359;
wire n_973;
wire n_1479;
wire n_1055;
wire n_1675;
wire n_582;
wire n_861;
wire n_857;
wire n_967;
wire n_571;
wire n_404;
wire n_271;
wire n_206;
wire n_679;
wire n_633;
wire n_1170;
wire n_665;
wire n_1629;
wire n_588;
wire n_225;
wire n_1260;
wire n_308;
wire n_309;
wire n_1010;
wire n_1040;
wire n_915;
wire n_632;
wire n_1166;
wire n_812;
wire n_1131;
wire n_1761;
wire n_534;
wire n_1578;
wire n_1006;
wire n_373;
wire n_1632;
wire n_257;
wire n_1557;
wire n_730;
wire n_1311;
wire n_1494;
wire n_670;
wire n_203;
wire n_207;
wire n_1089;
wire n_1587;
wire n_1365;
wire n_1417;
wire n_205;
wire n_1242;
wire n_681;
wire n_1226;
wire n_1274;
wire n_1486;
wire n_412;
wire n_640;
wire n_1322;
wire n_965;
wire n_1428;
wire n_1616;
wire n_1576;
wire n_339;
wire n_784;
wire n_434;
wire n_315;
wire n_288;
wire n_1059;
wire n_1197;
wire n_422;
wire n_722;
wire n_862;
wire n_165;
wire n_540;
wire n_1423;
wire n_457;
wire n_364;
wire n_629;
wire n_1621;
wire n_1748;
wire n_900;
wire n_1449;
wire n_531;
wire n_827;
wire n_361;
wire n_1025;
wire n_336;
wire n_1013;
wire n_1259;
wire n_192;
wire n_1538;
wire n_649;
wire n_1612;
wire n_1240;

CKINVDCx5p33_ASAP7_75t_R g165 ( 
.A(n_88),
.Y(n_165)
);

CKINVDCx5p33_ASAP7_75t_R g166 ( 
.A(n_12),
.Y(n_166)
);

CKINVDCx20_ASAP7_75t_R g167 ( 
.A(n_35),
.Y(n_167)
);

CKINVDCx5p33_ASAP7_75t_R g168 ( 
.A(n_153),
.Y(n_168)
);

CKINVDCx5p33_ASAP7_75t_R g169 ( 
.A(n_111),
.Y(n_169)
);

CKINVDCx5p33_ASAP7_75t_R g170 ( 
.A(n_25),
.Y(n_170)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_147),
.Y(n_171)
);

CKINVDCx5p33_ASAP7_75t_R g172 ( 
.A(n_96),
.Y(n_172)
);

BUFx10_ASAP7_75t_L g173 ( 
.A(n_140),
.Y(n_173)
);

CKINVDCx5p33_ASAP7_75t_R g174 ( 
.A(n_80),
.Y(n_174)
);

INVx2_ASAP7_75t_L g175 ( 
.A(n_123),
.Y(n_175)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_47),
.Y(n_176)
);

CKINVDCx5p33_ASAP7_75t_R g177 ( 
.A(n_128),
.Y(n_177)
);

CKINVDCx5p33_ASAP7_75t_R g178 ( 
.A(n_15),
.Y(n_178)
);

INVx2_ASAP7_75t_L g179 ( 
.A(n_79),
.Y(n_179)
);

CKINVDCx20_ASAP7_75t_R g180 ( 
.A(n_28),
.Y(n_180)
);

BUFx2_ASAP7_75t_L g181 ( 
.A(n_120),
.Y(n_181)
);

CKINVDCx5p33_ASAP7_75t_R g182 ( 
.A(n_110),
.Y(n_182)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_61),
.Y(n_183)
);

CKINVDCx20_ASAP7_75t_R g184 ( 
.A(n_95),
.Y(n_184)
);

CKINVDCx5p33_ASAP7_75t_R g185 ( 
.A(n_17),
.Y(n_185)
);

CKINVDCx20_ASAP7_75t_R g186 ( 
.A(n_17),
.Y(n_186)
);

INVx2_ASAP7_75t_L g187 ( 
.A(n_69),
.Y(n_187)
);

CKINVDCx5p33_ASAP7_75t_R g188 ( 
.A(n_85),
.Y(n_188)
);

INVx3_ASAP7_75t_L g189 ( 
.A(n_102),
.Y(n_189)
);

CKINVDCx5p33_ASAP7_75t_R g190 ( 
.A(n_118),
.Y(n_190)
);

BUFx10_ASAP7_75t_L g191 ( 
.A(n_86),
.Y(n_191)
);

CKINVDCx5p33_ASAP7_75t_R g192 ( 
.A(n_100),
.Y(n_192)
);

BUFx6f_ASAP7_75t_L g193 ( 
.A(n_93),
.Y(n_193)
);

CKINVDCx20_ASAP7_75t_R g194 ( 
.A(n_139),
.Y(n_194)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_114),
.Y(n_195)
);

CKINVDCx5p33_ASAP7_75t_R g196 ( 
.A(n_48),
.Y(n_196)
);

CKINVDCx5p33_ASAP7_75t_R g197 ( 
.A(n_129),
.Y(n_197)
);

CKINVDCx5p33_ASAP7_75t_R g198 ( 
.A(n_98),
.Y(n_198)
);

CKINVDCx5p33_ASAP7_75t_R g199 ( 
.A(n_40),
.Y(n_199)
);

INVx2_ASAP7_75t_SL g200 ( 
.A(n_58),
.Y(n_200)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_99),
.Y(n_201)
);

CKINVDCx5p33_ASAP7_75t_R g202 ( 
.A(n_119),
.Y(n_202)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_62),
.Y(n_203)
);

CKINVDCx5p33_ASAP7_75t_R g204 ( 
.A(n_50),
.Y(n_204)
);

CKINVDCx5p33_ASAP7_75t_R g205 ( 
.A(n_149),
.Y(n_205)
);

INVx2_ASAP7_75t_L g206 ( 
.A(n_37),
.Y(n_206)
);

CKINVDCx5p33_ASAP7_75t_R g207 ( 
.A(n_145),
.Y(n_207)
);

BUFx10_ASAP7_75t_L g208 ( 
.A(n_55),
.Y(n_208)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_0),
.Y(n_209)
);

CKINVDCx5p33_ASAP7_75t_R g210 ( 
.A(n_154),
.Y(n_210)
);

INVx1_ASAP7_75t_SL g211 ( 
.A(n_142),
.Y(n_211)
);

CKINVDCx5p33_ASAP7_75t_R g212 ( 
.A(n_104),
.Y(n_212)
);

INVx2_ASAP7_75t_SL g213 ( 
.A(n_109),
.Y(n_213)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_13),
.Y(n_214)
);

INVxp67_ASAP7_75t_L g215 ( 
.A(n_108),
.Y(n_215)
);

INVx1_ASAP7_75t_SL g216 ( 
.A(n_53),
.Y(n_216)
);

CKINVDCx5p33_ASAP7_75t_R g217 ( 
.A(n_103),
.Y(n_217)
);

CKINVDCx20_ASAP7_75t_R g218 ( 
.A(n_20),
.Y(n_218)
);

CKINVDCx5p33_ASAP7_75t_R g219 ( 
.A(n_126),
.Y(n_219)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_64),
.Y(n_220)
);

CKINVDCx5p33_ASAP7_75t_R g221 ( 
.A(n_151),
.Y(n_221)
);

CKINVDCx20_ASAP7_75t_R g222 ( 
.A(n_162),
.Y(n_222)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_65),
.Y(n_223)
);

CKINVDCx5p33_ASAP7_75t_R g224 ( 
.A(n_20),
.Y(n_224)
);

CKINVDCx5p33_ASAP7_75t_R g225 ( 
.A(n_60),
.Y(n_225)
);

CKINVDCx5p33_ASAP7_75t_R g226 ( 
.A(n_57),
.Y(n_226)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_157),
.Y(n_227)
);

INVx2_ASAP7_75t_L g228 ( 
.A(n_49),
.Y(n_228)
);

INVx1_ASAP7_75t_SL g229 ( 
.A(n_138),
.Y(n_229)
);

CKINVDCx5p33_ASAP7_75t_R g230 ( 
.A(n_161),
.Y(n_230)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_94),
.Y(n_231)
);

CKINVDCx5p33_ASAP7_75t_R g232 ( 
.A(n_34),
.Y(n_232)
);

CKINVDCx5p33_ASAP7_75t_R g233 ( 
.A(n_7),
.Y(n_233)
);

BUFx6f_ASAP7_75t_L g234 ( 
.A(n_113),
.Y(n_234)
);

INVx2_ASAP7_75t_L g235 ( 
.A(n_38),
.Y(n_235)
);

CKINVDCx5p33_ASAP7_75t_R g236 ( 
.A(n_57),
.Y(n_236)
);

CKINVDCx20_ASAP7_75t_R g237 ( 
.A(n_15),
.Y(n_237)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_116),
.Y(n_238)
);

CKINVDCx5p33_ASAP7_75t_R g239 ( 
.A(n_23),
.Y(n_239)
);

INVx2_ASAP7_75t_SL g240 ( 
.A(n_40),
.Y(n_240)
);

CKINVDCx5p33_ASAP7_75t_R g241 ( 
.A(n_54),
.Y(n_241)
);

CKINVDCx5p33_ASAP7_75t_R g242 ( 
.A(n_107),
.Y(n_242)
);

CKINVDCx5p33_ASAP7_75t_R g243 ( 
.A(n_38),
.Y(n_243)
);

INVx2_ASAP7_75t_SL g244 ( 
.A(n_91),
.Y(n_244)
);

CKINVDCx5p33_ASAP7_75t_R g245 ( 
.A(n_81),
.Y(n_245)
);

CKINVDCx5p33_ASAP7_75t_R g246 ( 
.A(n_31),
.Y(n_246)
);

CKINVDCx5p33_ASAP7_75t_R g247 ( 
.A(n_30),
.Y(n_247)
);

CKINVDCx5p33_ASAP7_75t_R g248 ( 
.A(n_67),
.Y(n_248)
);

CKINVDCx5p33_ASAP7_75t_R g249 ( 
.A(n_158),
.Y(n_249)
);

CKINVDCx5p33_ASAP7_75t_R g250 ( 
.A(n_132),
.Y(n_250)
);

BUFx6f_ASAP7_75t_L g251 ( 
.A(n_55),
.Y(n_251)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_97),
.Y(n_252)
);

BUFx6f_ASAP7_75t_L g253 ( 
.A(n_121),
.Y(n_253)
);

CKINVDCx5p33_ASAP7_75t_R g254 ( 
.A(n_35),
.Y(n_254)
);

CKINVDCx5p33_ASAP7_75t_R g255 ( 
.A(n_136),
.Y(n_255)
);

BUFx6f_ASAP7_75t_L g256 ( 
.A(n_152),
.Y(n_256)
);

CKINVDCx5p33_ASAP7_75t_R g257 ( 
.A(n_163),
.Y(n_257)
);

BUFx6f_ASAP7_75t_L g258 ( 
.A(n_6),
.Y(n_258)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_46),
.Y(n_259)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_53),
.Y(n_260)
);

CKINVDCx5p33_ASAP7_75t_R g261 ( 
.A(n_44),
.Y(n_261)
);

CKINVDCx5p33_ASAP7_75t_R g262 ( 
.A(n_50),
.Y(n_262)
);

CKINVDCx20_ASAP7_75t_R g263 ( 
.A(n_33),
.Y(n_263)
);

INVx2_ASAP7_75t_L g264 ( 
.A(n_90),
.Y(n_264)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_135),
.Y(n_265)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_27),
.Y(n_266)
);

CKINVDCx5p33_ASAP7_75t_R g267 ( 
.A(n_7),
.Y(n_267)
);

CKINVDCx20_ASAP7_75t_R g268 ( 
.A(n_141),
.Y(n_268)
);

CKINVDCx5p33_ASAP7_75t_R g269 ( 
.A(n_45),
.Y(n_269)
);

CKINVDCx5p33_ASAP7_75t_R g270 ( 
.A(n_73),
.Y(n_270)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_56),
.Y(n_271)
);

CKINVDCx5p33_ASAP7_75t_R g272 ( 
.A(n_87),
.Y(n_272)
);

INVx2_ASAP7_75t_L g273 ( 
.A(n_58),
.Y(n_273)
);

CKINVDCx5p33_ASAP7_75t_R g274 ( 
.A(n_8),
.Y(n_274)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_34),
.Y(n_275)
);

CKINVDCx5p33_ASAP7_75t_R g276 ( 
.A(n_125),
.Y(n_276)
);

CKINVDCx5p33_ASAP7_75t_R g277 ( 
.A(n_48),
.Y(n_277)
);

CKINVDCx5p33_ASAP7_75t_R g278 ( 
.A(n_41),
.Y(n_278)
);

CKINVDCx5p33_ASAP7_75t_R g279 ( 
.A(n_49),
.Y(n_279)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_122),
.Y(n_280)
);

CKINVDCx5p33_ASAP7_75t_R g281 ( 
.A(n_60),
.Y(n_281)
);

CKINVDCx5p33_ASAP7_75t_R g282 ( 
.A(n_33),
.Y(n_282)
);

CKINVDCx5p33_ASAP7_75t_R g283 ( 
.A(n_43),
.Y(n_283)
);

CKINVDCx5p33_ASAP7_75t_R g284 ( 
.A(n_54),
.Y(n_284)
);

INVxp67_ASAP7_75t_L g285 ( 
.A(n_37),
.Y(n_285)
);

CKINVDCx5p33_ASAP7_75t_R g286 ( 
.A(n_22),
.Y(n_286)
);

CKINVDCx5p33_ASAP7_75t_R g287 ( 
.A(n_2),
.Y(n_287)
);

BUFx3_ASAP7_75t_L g288 ( 
.A(n_74),
.Y(n_288)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_59),
.Y(n_289)
);

CKINVDCx20_ASAP7_75t_R g290 ( 
.A(n_89),
.Y(n_290)
);

CKINVDCx5p33_ASAP7_75t_R g291 ( 
.A(n_21),
.Y(n_291)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_82),
.Y(n_292)
);

CKINVDCx5p33_ASAP7_75t_R g293 ( 
.A(n_24),
.Y(n_293)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_144),
.Y(n_294)
);

INVx2_ASAP7_75t_L g295 ( 
.A(n_150),
.Y(n_295)
);

CKINVDCx20_ASAP7_75t_R g296 ( 
.A(n_0),
.Y(n_296)
);

CKINVDCx5p33_ASAP7_75t_R g297 ( 
.A(n_130),
.Y(n_297)
);

CKINVDCx5p33_ASAP7_75t_R g298 ( 
.A(n_156),
.Y(n_298)
);

BUFx3_ASAP7_75t_L g299 ( 
.A(n_164),
.Y(n_299)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_13),
.Y(n_300)
);

CKINVDCx5p33_ASAP7_75t_R g301 ( 
.A(n_47),
.Y(n_301)
);

CKINVDCx20_ASAP7_75t_R g302 ( 
.A(n_36),
.Y(n_302)
);

CKINVDCx5p33_ASAP7_75t_R g303 ( 
.A(n_36),
.Y(n_303)
);

BUFx2_ASAP7_75t_L g304 ( 
.A(n_52),
.Y(n_304)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_78),
.Y(n_305)
);

CKINVDCx5p33_ASAP7_75t_R g306 ( 
.A(n_4),
.Y(n_306)
);

INVx1_ASAP7_75t_SL g307 ( 
.A(n_3),
.Y(n_307)
);

CKINVDCx5p33_ASAP7_75t_R g308 ( 
.A(n_29),
.Y(n_308)
);

INVx2_ASAP7_75t_L g309 ( 
.A(n_28),
.Y(n_309)
);

CKINVDCx5p33_ASAP7_75t_R g310 ( 
.A(n_148),
.Y(n_310)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_41),
.Y(n_311)
);

CKINVDCx5p33_ASAP7_75t_R g312 ( 
.A(n_24),
.Y(n_312)
);

CKINVDCx5p33_ASAP7_75t_R g313 ( 
.A(n_52),
.Y(n_313)
);

BUFx6f_ASAP7_75t_L g314 ( 
.A(n_155),
.Y(n_314)
);

CKINVDCx5p33_ASAP7_75t_R g315 ( 
.A(n_4),
.Y(n_315)
);

CKINVDCx5p33_ASAP7_75t_R g316 ( 
.A(n_106),
.Y(n_316)
);

INVx2_ASAP7_75t_L g317 ( 
.A(n_9),
.Y(n_317)
);

CKINVDCx5p33_ASAP7_75t_R g318 ( 
.A(n_76),
.Y(n_318)
);

CKINVDCx5p33_ASAP7_75t_R g319 ( 
.A(n_12),
.Y(n_319)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_56),
.Y(n_320)
);

INVx2_ASAP7_75t_L g321 ( 
.A(n_18),
.Y(n_321)
);

CKINVDCx5p33_ASAP7_75t_R g322 ( 
.A(n_61),
.Y(n_322)
);

CKINVDCx5p33_ASAP7_75t_R g323 ( 
.A(n_105),
.Y(n_323)
);

CKINVDCx14_ASAP7_75t_R g324 ( 
.A(n_44),
.Y(n_324)
);

CKINVDCx5p33_ASAP7_75t_R g325 ( 
.A(n_112),
.Y(n_325)
);

CKINVDCx5p33_ASAP7_75t_R g326 ( 
.A(n_146),
.Y(n_326)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_77),
.Y(n_327)
);

CKINVDCx20_ASAP7_75t_R g328 ( 
.A(n_184),
.Y(n_328)
);

CKINVDCx5p33_ASAP7_75t_R g329 ( 
.A(n_165),
.Y(n_329)
);

BUFx2_ASAP7_75t_L g330 ( 
.A(n_304),
.Y(n_330)
);

BUFx6f_ASAP7_75t_SL g331 ( 
.A(n_173),
.Y(n_331)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_251),
.Y(n_332)
);

CKINVDCx5p33_ASAP7_75t_R g333 ( 
.A(n_168),
.Y(n_333)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_251),
.Y(n_334)
);

CKINVDCx20_ASAP7_75t_R g335 ( 
.A(n_194),
.Y(n_335)
);

CKINVDCx16_ASAP7_75t_R g336 ( 
.A(n_324),
.Y(n_336)
);

INVxp67_ASAP7_75t_L g337 ( 
.A(n_304),
.Y(n_337)
);

CKINVDCx5p33_ASAP7_75t_R g338 ( 
.A(n_169),
.Y(n_338)
);

CKINVDCx5p33_ASAP7_75t_R g339 ( 
.A(n_172),
.Y(n_339)
);

CKINVDCx20_ASAP7_75t_R g340 ( 
.A(n_222),
.Y(n_340)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_251),
.Y(n_341)
);

CKINVDCx5p33_ASAP7_75t_R g342 ( 
.A(n_174),
.Y(n_342)
);

CKINVDCx5p33_ASAP7_75t_R g343 ( 
.A(n_177),
.Y(n_343)
);

CKINVDCx20_ASAP7_75t_R g344 ( 
.A(n_268),
.Y(n_344)
);

BUFx6f_ASAP7_75t_SL g345 ( 
.A(n_173),
.Y(n_345)
);

CKINVDCx5p33_ASAP7_75t_R g346 ( 
.A(n_182),
.Y(n_346)
);

INVxp67_ASAP7_75t_L g347 ( 
.A(n_176),
.Y(n_347)
);

INVx1_ASAP7_75t_L g348 ( 
.A(n_251),
.Y(n_348)
);

CKINVDCx16_ASAP7_75t_R g349 ( 
.A(n_208),
.Y(n_349)
);

INVx1_ASAP7_75t_SL g350 ( 
.A(n_167),
.Y(n_350)
);

INVx1_ASAP7_75t_L g351 ( 
.A(n_251),
.Y(n_351)
);

CKINVDCx20_ASAP7_75t_R g352 ( 
.A(n_290),
.Y(n_352)
);

INVxp67_ASAP7_75t_L g353 ( 
.A(n_176),
.Y(n_353)
);

INVx1_ASAP7_75t_L g354 ( 
.A(n_258),
.Y(n_354)
);

INVx1_ASAP7_75t_L g355 ( 
.A(n_258),
.Y(n_355)
);

INVx2_ASAP7_75t_L g356 ( 
.A(n_258),
.Y(n_356)
);

NOR2xp33_ASAP7_75t_L g357 ( 
.A(n_181),
.B(n_1),
.Y(n_357)
);

CKINVDCx5p33_ASAP7_75t_R g358 ( 
.A(n_188),
.Y(n_358)
);

INVxp67_ASAP7_75t_SL g359 ( 
.A(n_181),
.Y(n_359)
);

CKINVDCx5p33_ASAP7_75t_R g360 ( 
.A(n_190),
.Y(n_360)
);

CKINVDCx5p33_ASAP7_75t_R g361 ( 
.A(n_192),
.Y(n_361)
);

CKINVDCx5p33_ASAP7_75t_R g362 ( 
.A(n_197),
.Y(n_362)
);

CKINVDCx20_ASAP7_75t_R g363 ( 
.A(n_198),
.Y(n_363)
);

CKINVDCx5p33_ASAP7_75t_R g364 ( 
.A(n_202),
.Y(n_364)
);

INVx1_ASAP7_75t_L g365 ( 
.A(n_258),
.Y(n_365)
);

CKINVDCx5p33_ASAP7_75t_R g366 ( 
.A(n_205),
.Y(n_366)
);

CKINVDCx20_ASAP7_75t_R g367 ( 
.A(n_207),
.Y(n_367)
);

BUFx3_ASAP7_75t_L g368 ( 
.A(n_288),
.Y(n_368)
);

NAND2xp5_ASAP7_75t_L g369 ( 
.A(n_213),
.B(n_1),
.Y(n_369)
);

INVx1_ASAP7_75t_L g370 ( 
.A(n_258),
.Y(n_370)
);

INVx1_ASAP7_75t_L g371 ( 
.A(n_206),
.Y(n_371)
);

CKINVDCx20_ASAP7_75t_R g372 ( 
.A(n_210),
.Y(n_372)
);

CKINVDCx20_ASAP7_75t_R g373 ( 
.A(n_212),
.Y(n_373)
);

CKINVDCx5p33_ASAP7_75t_R g374 ( 
.A(n_217),
.Y(n_374)
);

INVx1_ASAP7_75t_L g375 ( 
.A(n_206),
.Y(n_375)
);

NOR2xp67_ASAP7_75t_L g376 ( 
.A(n_189),
.B(n_2),
.Y(n_376)
);

CKINVDCx5p33_ASAP7_75t_R g377 ( 
.A(n_219),
.Y(n_377)
);

INVx1_ASAP7_75t_L g378 ( 
.A(n_228),
.Y(n_378)
);

CKINVDCx16_ASAP7_75t_R g379 ( 
.A(n_208),
.Y(n_379)
);

INVx1_ASAP7_75t_L g380 ( 
.A(n_228),
.Y(n_380)
);

INVx1_ASAP7_75t_L g381 ( 
.A(n_235),
.Y(n_381)
);

INVx1_ASAP7_75t_L g382 ( 
.A(n_235),
.Y(n_382)
);

XNOR2xp5_ASAP7_75t_L g383 ( 
.A(n_180),
.B(n_186),
.Y(n_383)
);

HB1xp67_ASAP7_75t_L g384 ( 
.A(n_166),
.Y(n_384)
);

HB1xp67_ASAP7_75t_L g385 ( 
.A(n_170),
.Y(n_385)
);

INVx1_ASAP7_75t_L g386 ( 
.A(n_273),
.Y(n_386)
);

CKINVDCx16_ASAP7_75t_R g387 ( 
.A(n_208),
.Y(n_387)
);

NOR2xp33_ASAP7_75t_L g388 ( 
.A(n_213),
.B(n_3),
.Y(n_388)
);

INVx1_ASAP7_75t_L g389 ( 
.A(n_273),
.Y(n_389)
);

NAND2xp33_ASAP7_75t_R g390 ( 
.A(n_189),
.B(n_5),
.Y(n_390)
);

NOR2xp33_ASAP7_75t_R g391 ( 
.A(n_221),
.B(n_101),
.Y(n_391)
);

CKINVDCx20_ASAP7_75t_R g392 ( 
.A(n_230),
.Y(n_392)
);

INVx1_ASAP7_75t_L g393 ( 
.A(n_309),
.Y(n_393)
);

INVx1_ASAP7_75t_L g394 ( 
.A(n_309),
.Y(n_394)
);

CKINVDCx20_ASAP7_75t_R g395 ( 
.A(n_242),
.Y(n_395)
);

CKINVDCx5p33_ASAP7_75t_R g396 ( 
.A(n_245),
.Y(n_396)
);

INVx1_ASAP7_75t_L g397 ( 
.A(n_317),
.Y(n_397)
);

INVx1_ASAP7_75t_L g398 ( 
.A(n_317),
.Y(n_398)
);

INVx1_ASAP7_75t_L g399 ( 
.A(n_321),
.Y(n_399)
);

CKINVDCx5p33_ASAP7_75t_R g400 ( 
.A(n_248),
.Y(n_400)
);

CKINVDCx5p33_ASAP7_75t_R g401 ( 
.A(n_249),
.Y(n_401)
);

CKINVDCx20_ASAP7_75t_R g402 ( 
.A(n_250),
.Y(n_402)
);

CKINVDCx20_ASAP7_75t_R g403 ( 
.A(n_255),
.Y(n_403)
);

INVx1_ASAP7_75t_L g404 ( 
.A(n_321),
.Y(n_404)
);

CKINVDCx5p33_ASAP7_75t_R g405 ( 
.A(n_257),
.Y(n_405)
);

BUFx6f_ASAP7_75t_L g406 ( 
.A(n_356),
.Y(n_406)
);

BUFx6f_ASAP7_75t_L g407 ( 
.A(n_356),
.Y(n_407)
);

INVx2_ASAP7_75t_L g408 ( 
.A(n_332),
.Y(n_408)
);

AND2x6_ASAP7_75t_L g409 ( 
.A(n_332),
.B(n_189),
.Y(n_409)
);

NAND2xp5_ASAP7_75t_L g410 ( 
.A(n_388),
.B(n_244),
.Y(n_410)
);

INVx1_ASAP7_75t_L g411 ( 
.A(n_334),
.Y(n_411)
);

INVxp67_ASAP7_75t_L g412 ( 
.A(n_384),
.Y(n_412)
);

BUFx6f_ASAP7_75t_L g413 ( 
.A(n_334),
.Y(n_413)
);

INVx1_ASAP7_75t_L g414 ( 
.A(n_341),
.Y(n_414)
);

BUFx6f_ASAP7_75t_L g415 ( 
.A(n_341),
.Y(n_415)
);

BUFx6f_ASAP7_75t_L g416 ( 
.A(n_348),
.Y(n_416)
);

INVx2_ASAP7_75t_L g417 ( 
.A(n_348),
.Y(n_417)
);

INVx2_ASAP7_75t_L g418 ( 
.A(n_351),
.Y(n_418)
);

NAND2xp5_ASAP7_75t_L g419 ( 
.A(n_351),
.B(n_354),
.Y(n_419)
);

INVx1_ASAP7_75t_L g420 ( 
.A(n_354),
.Y(n_420)
);

INVx1_ASAP7_75t_L g421 ( 
.A(n_355),
.Y(n_421)
);

BUFx6f_ASAP7_75t_L g422 ( 
.A(n_355),
.Y(n_422)
);

AND3x1_ASAP7_75t_L g423 ( 
.A(n_357),
.B(n_369),
.C(n_240),
.Y(n_423)
);

INVx1_ASAP7_75t_L g424 ( 
.A(n_365),
.Y(n_424)
);

INVxp67_ASAP7_75t_L g425 ( 
.A(n_385),
.Y(n_425)
);

INVx1_ASAP7_75t_L g426 ( 
.A(n_365),
.Y(n_426)
);

INVx2_ASAP7_75t_L g427 ( 
.A(n_370),
.Y(n_427)
);

INVx3_ASAP7_75t_L g428 ( 
.A(n_370),
.Y(n_428)
);

INVx1_ASAP7_75t_L g429 ( 
.A(n_371),
.Y(n_429)
);

NAND2xp33_ASAP7_75t_L g430 ( 
.A(n_391),
.B(n_200),
.Y(n_430)
);

INVx1_ASAP7_75t_L g431 ( 
.A(n_371),
.Y(n_431)
);

INVx2_ASAP7_75t_L g432 ( 
.A(n_375),
.Y(n_432)
);

INVx1_ASAP7_75t_L g433 ( 
.A(n_375),
.Y(n_433)
);

INVx2_ASAP7_75t_L g434 ( 
.A(n_378),
.Y(n_434)
);

BUFx6f_ASAP7_75t_L g435 ( 
.A(n_378),
.Y(n_435)
);

INVx1_ASAP7_75t_L g436 ( 
.A(n_380),
.Y(n_436)
);

NAND2xp5_ASAP7_75t_L g437 ( 
.A(n_368),
.B(n_244),
.Y(n_437)
);

INVx1_ASAP7_75t_L g438 ( 
.A(n_380),
.Y(n_438)
);

BUFx6f_ASAP7_75t_L g439 ( 
.A(n_381),
.Y(n_439)
);

AND2x2_ASAP7_75t_L g440 ( 
.A(n_368),
.B(n_288),
.Y(n_440)
);

NAND2xp5_ASAP7_75t_SL g441 ( 
.A(n_376),
.B(n_173),
.Y(n_441)
);

AND2x2_ASAP7_75t_L g442 ( 
.A(n_359),
.B(n_381),
.Y(n_442)
);

NAND2xp5_ASAP7_75t_L g443 ( 
.A(n_347),
.B(n_270),
.Y(n_443)
);

INVxp67_ASAP7_75t_L g444 ( 
.A(n_330),
.Y(n_444)
);

INVx1_ASAP7_75t_L g445 ( 
.A(n_382),
.Y(n_445)
);

NAND2xp5_ASAP7_75t_L g446 ( 
.A(n_353),
.B(n_272),
.Y(n_446)
);

INVx2_ASAP7_75t_L g447 ( 
.A(n_382),
.Y(n_447)
);

INVx2_ASAP7_75t_L g448 ( 
.A(n_386),
.Y(n_448)
);

AND2x4_ASAP7_75t_L g449 ( 
.A(n_386),
.B(n_189),
.Y(n_449)
);

INVx1_ASAP7_75t_L g450 ( 
.A(n_389),
.Y(n_450)
);

BUFx6f_ASAP7_75t_L g451 ( 
.A(n_389),
.Y(n_451)
);

AND2x4_ASAP7_75t_L g452 ( 
.A(n_393),
.B(n_288),
.Y(n_452)
);

NAND2xp5_ASAP7_75t_L g453 ( 
.A(n_393),
.B(n_276),
.Y(n_453)
);

INVx2_ASAP7_75t_L g454 ( 
.A(n_394),
.Y(n_454)
);

INVx1_ASAP7_75t_L g455 ( 
.A(n_394),
.Y(n_455)
);

INVx1_ASAP7_75t_L g456 ( 
.A(n_397),
.Y(n_456)
);

AND2x2_ASAP7_75t_L g457 ( 
.A(n_397),
.B(n_299),
.Y(n_457)
);

INVx3_ASAP7_75t_L g458 ( 
.A(n_398),
.Y(n_458)
);

CKINVDCx5p33_ASAP7_75t_R g459 ( 
.A(n_329),
.Y(n_459)
);

INVx1_ASAP7_75t_L g460 ( 
.A(n_398),
.Y(n_460)
);

INVx1_ASAP7_75t_L g461 ( 
.A(n_399),
.Y(n_461)
);

BUFx8_ASAP7_75t_L g462 ( 
.A(n_331),
.Y(n_462)
);

AND2x2_ASAP7_75t_L g463 ( 
.A(n_399),
.B(n_299),
.Y(n_463)
);

INVx2_ASAP7_75t_L g464 ( 
.A(n_404),
.Y(n_464)
);

INVx2_ASAP7_75t_L g465 ( 
.A(n_404),
.Y(n_465)
);

INVx1_ASAP7_75t_L g466 ( 
.A(n_333),
.Y(n_466)
);

NOR2xp33_ASAP7_75t_L g467 ( 
.A(n_337),
.B(n_215),
.Y(n_467)
);

INVx2_ASAP7_75t_L g468 ( 
.A(n_338),
.Y(n_468)
);

AND2x2_ASAP7_75t_L g469 ( 
.A(n_336),
.B(n_299),
.Y(n_469)
);

NAND2xp33_ASAP7_75t_L g470 ( 
.A(n_390),
.B(n_200),
.Y(n_470)
);

INVx2_ASAP7_75t_L g471 ( 
.A(n_339),
.Y(n_471)
);

HB1xp67_ASAP7_75t_L g472 ( 
.A(n_330),
.Y(n_472)
);

INVx3_ASAP7_75t_L g473 ( 
.A(n_342),
.Y(n_473)
);

HB1xp67_ASAP7_75t_L g474 ( 
.A(n_350),
.Y(n_474)
);

INVx2_ASAP7_75t_L g475 ( 
.A(n_343),
.Y(n_475)
);

INVx2_ASAP7_75t_L g476 ( 
.A(n_346),
.Y(n_476)
);

INVx2_ASAP7_75t_L g477 ( 
.A(n_358),
.Y(n_477)
);

NAND2xp5_ASAP7_75t_L g478 ( 
.A(n_360),
.B(n_297),
.Y(n_478)
);

INVx1_ASAP7_75t_L g479 ( 
.A(n_361),
.Y(n_479)
);

AOI22xp33_ASAP7_75t_L g480 ( 
.A1(n_410),
.A2(n_240),
.B1(n_260),
.B2(n_259),
.Y(n_480)
);

INVx6_ASAP7_75t_L g481 ( 
.A(n_452),
.Y(n_481)
);

INVx3_ASAP7_75t_L g482 ( 
.A(n_406),
.Y(n_482)
);

INVxp67_ASAP7_75t_SL g483 ( 
.A(n_437),
.Y(n_483)
);

AND2x6_ASAP7_75t_L g484 ( 
.A(n_468),
.B(n_179),
.Y(n_484)
);

INVx1_ASAP7_75t_L g485 ( 
.A(n_414),
.Y(n_485)
);

INVx1_ASAP7_75t_L g486 ( 
.A(n_414),
.Y(n_486)
);

BUFx4f_ASAP7_75t_L g487 ( 
.A(n_409),
.Y(n_487)
);

NOR2xp33_ASAP7_75t_L g488 ( 
.A(n_466),
.B(n_362),
.Y(n_488)
);

CKINVDCx5p33_ASAP7_75t_R g489 ( 
.A(n_459),
.Y(n_489)
);

INVx4_ASAP7_75t_L g490 ( 
.A(n_409),
.Y(n_490)
);

NAND2xp5_ASAP7_75t_L g491 ( 
.A(n_410),
.B(n_364),
.Y(n_491)
);

NAND2xp5_ASAP7_75t_L g492 ( 
.A(n_478),
.B(n_366),
.Y(n_492)
);

INVx3_ASAP7_75t_L g493 ( 
.A(n_406),
.Y(n_493)
);

NAND2xp5_ASAP7_75t_L g494 ( 
.A(n_478),
.B(n_374),
.Y(n_494)
);

BUFx6f_ASAP7_75t_L g495 ( 
.A(n_406),
.Y(n_495)
);

AOI22xp33_ASAP7_75t_L g496 ( 
.A1(n_442),
.A2(n_470),
.B1(n_467),
.B2(n_452),
.Y(n_496)
);

BUFx6f_ASAP7_75t_L g497 ( 
.A(n_406),
.Y(n_497)
);

AND2x4_ASAP7_75t_L g498 ( 
.A(n_452),
.B(n_171),
.Y(n_498)
);

NAND2xp5_ASAP7_75t_L g499 ( 
.A(n_468),
.B(n_377),
.Y(n_499)
);

INVx2_ASAP7_75t_L g500 ( 
.A(n_408),
.Y(n_500)
);

NAND2xp5_ASAP7_75t_SL g501 ( 
.A(n_468),
.B(n_396),
.Y(n_501)
);

CKINVDCx5p33_ASAP7_75t_R g502 ( 
.A(n_474),
.Y(n_502)
);

OR2x2_ASAP7_75t_L g503 ( 
.A(n_472),
.B(n_387),
.Y(n_503)
);

INVx1_ASAP7_75t_L g504 ( 
.A(n_426),
.Y(n_504)
);

AND2x4_ASAP7_75t_L g505 ( 
.A(n_452),
.B(n_171),
.Y(n_505)
);

NAND2xp33_ASAP7_75t_R g506 ( 
.A(n_469),
.B(n_400),
.Y(n_506)
);

NAND2xp5_ASAP7_75t_L g507 ( 
.A(n_468),
.B(n_401),
.Y(n_507)
);

INVx5_ASAP7_75t_L g508 ( 
.A(n_409),
.Y(n_508)
);

BUFx3_ASAP7_75t_L g509 ( 
.A(n_440),
.Y(n_509)
);

BUFx6f_ASAP7_75t_L g510 ( 
.A(n_406),
.Y(n_510)
);

INVx1_ASAP7_75t_L g511 ( 
.A(n_426),
.Y(n_511)
);

NAND3xp33_ASAP7_75t_L g512 ( 
.A(n_467),
.B(n_405),
.C(n_185),
.Y(n_512)
);

BUFx3_ASAP7_75t_L g513 ( 
.A(n_440),
.Y(n_513)
);

BUFx3_ASAP7_75t_L g514 ( 
.A(n_440),
.Y(n_514)
);

INVx2_ASAP7_75t_L g515 ( 
.A(n_408),
.Y(n_515)
);

NAND2xp5_ASAP7_75t_SL g516 ( 
.A(n_471),
.B(n_387),
.Y(n_516)
);

INVx2_ASAP7_75t_L g517 ( 
.A(n_417),
.Y(n_517)
);

INVx1_ASAP7_75t_L g518 ( 
.A(n_419),
.Y(n_518)
);

NOR2x1_ASAP7_75t_L g519 ( 
.A(n_473),
.B(n_195),
.Y(n_519)
);

INVx2_ASAP7_75t_L g520 ( 
.A(n_417),
.Y(n_520)
);

INVx2_ASAP7_75t_L g521 ( 
.A(n_417),
.Y(n_521)
);

INVx2_ASAP7_75t_L g522 ( 
.A(n_417),
.Y(n_522)
);

BUFx3_ASAP7_75t_L g523 ( 
.A(n_452),
.Y(n_523)
);

NAND2xp5_ASAP7_75t_SL g524 ( 
.A(n_471),
.B(n_349),
.Y(n_524)
);

INVx1_ASAP7_75t_L g525 ( 
.A(n_419),
.Y(n_525)
);

NAND2xp5_ASAP7_75t_L g526 ( 
.A(n_471),
.B(n_211),
.Y(n_526)
);

NAND2xp5_ASAP7_75t_SL g527 ( 
.A(n_471),
.B(n_379),
.Y(n_527)
);

AOI22xp33_ASAP7_75t_L g528 ( 
.A1(n_442),
.A2(n_300),
.B1(n_289),
.B2(n_275),
.Y(n_528)
);

INVx2_ASAP7_75t_SL g529 ( 
.A(n_469),
.Y(n_529)
);

BUFx10_ASAP7_75t_L g530 ( 
.A(n_466),
.Y(n_530)
);

AOI22xp33_ASAP7_75t_L g531 ( 
.A1(n_442),
.A2(n_300),
.B1(n_289),
.B2(n_275),
.Y(n_531)
);

BUFx10_ASAP7_75t_L g532 ( 
.A(n_466),
.Y(n_532)
);

NOR2xp33_ASAP7_75t_L g533 ( 
.A(n_479),
.B(n_363),
.Y(n_533)
);

INVx1_ASAP7_75t_L g534 ( 
.A(n_411),
.Y(n_534)
);

INVx2_ASAP7_75t_SL g535 ( 
.A(n_469),
.Y(n_535)
);

OR2x2_ASAP7_75t_L g536 ( 
.A(n_472),
.B(n_383),
.Y(n_536)
);

AND2x4_ASAP7_75t_L g537 ( 
.A(n_452),
.B(n_195),
.Y(n_537)
);

OAI22xp5_ASAP7_75t_L g538 ( 
.A1(n_479),
.A2(n_403),
.B1(n_402),
.B2(n_395),
.Y(n_538)
);

INVx2_ASAP7_75t_L g539 ( 
.A(n_418),
.Y(n_539)
);

INVx4_ASAP7_75t_L g540 ( 
.A(n_409),
.Y(n_540)
);

INVx2_ASAP7_75t_L g541 ( 
.A(n_418),
.Y(n_541)
);

AND2x4_ASAP7_75t_L g542 ( 
.A(n_449),
.B(n_201),
.Y(n_542)
);

BUFx8_ASAP7_75t_SL g543 ( 
.A(n_473),
.Y(n_543)
);

INVx2_ASAP7_75t_L g544 ( 
.A(n_418),
.Y(n_544)
);

AOI22xp33_ASAP7_75t_L g545 ( 
.A1(n_470),
.A2(n_260),
.B1(n_209),
.B2(n_311),
.Y(n_545)
);

NAND2xp5_ASAP7_75t_SL g546 ( 
.A(n_475),
.B(n_367),
.Y(n_546)
);

INVx2_ASAP7_75t_L g547 ( 
.A(n_418),
.Y(n_547)
);

NAND2xp5_ASAP7_75t_L g548 ( 
.A(n_475),
.B(n_229),
.Y(n_548)
);

INVx2_ASAP7_75t_L g549 ( 
.A(n_427),
.Y(n_549)
);

INVx2_ASAP7_75t_L g550 ( 
.A(n_427),
.Y(n_550)
);

NAND2xp5_ASAP7_75t_SL g551 ( 
.A(n_475),
.B(n_372),
.Y(n_551)
);

AOI22xp33_ASAP7_75t_L g552 ( 
.A1(n_441),
.A2(n_214),
.B1(n_209),
.B2(n_311),
.Y(n_552)
);

NAND2xp5_ASAP7_75t_L g553 ( 
.A(n_475),
.B(n_298),
.Y(n_553)
);

INVx2_ASAP7_75t_SL g554 ( 
.A(n_474),
.Y(n_554)
);

INVx1_ASAP7_75t_L g555 ( 
.A(n_411),
.Y(n_555)
);

BUFx6f_ASAP7_75t_L g556 ( 
.A(n_406),
.Y(n_556)
);

NAND2xp5_ASAP7_75t_SL g557 ( 
.A(n_476),
.B(n_373),
.Y(n_557)
);

NAND2xp33_ASAP7_75t_L g558 ( 
.A(n_409),
.B(n_193),
.Y(n_558)
);

INVx1_ASAP7_75t_L g559 ( 
.A(n_411),
.Y(n_559)
);

BUFx3_ASAP7_75t_L g560 ( 
.A(n_457),
.Y(n_560)
);

INVx1_ASAP7_75t_L g561 ( 
.A(n_420),
.Y(n_561)
);

CKINVDCx20_ASAP7_75t_R g562 ( 
.A(n_462),
.Y(n_562)
);

NAND2xp5_ASAP7_75t_L g563 ( 
.A(n_476),
.B(n_310),
.Y(n_563)
);

NAND2xp5_ASAP7_75t_SL g564 ( 
.A(n_476),
.B(n_392),
.Y(n_564)
);

INVx2_ASAP7_75t_SL g565 ( 
.A(n_443),
.Y(n_565)
);

AND2x6_ASAP7_75t_L g566 ( 
.A(n_476),
.B(n_179),
.Y(n_566)
);

INVx3_ASAP7_75t_L g567 ( 
.A(n_406),
.Y(n_567)
);

AND2x2_ASAP7_75t_L g568 ( 
.A(n_457),
.B(n_463),
.Y(n_568)
);

INVx3_ASAP7_75t_L g569 ( 
.A(n_406),
.Y(n_569)
);

AOI22xp33_ASAP7_75t_L g570 ( 
.A1(n_441),
.A2(n_266),
.B1(n_271),
.B2(n_320),
.Y(n_570)
);

NAND2xp5_ASAP7_75t_L g571 ( 
.A(n_477),
.B(n_316),
.Y(n_571)
);

INVx1_ASAP7_75t_L g572 ( 
.A(n_420),
.Y(n_572)
);

OAI22xp33_ASAP7_75t_L g573 ( 
.A1(n_412),
.A2(n_216),
.B1(n_307),
.B2(n_262),
.Y(n_573)
);

INVx1_ASAP7_75t_L g574 ( 
.A(n_420),
.Y(n_574)
);

INVx2_ASAP7_75t_L g575 ( 
.A(n_427),
.Y(n_575)
);

AOI22xp5_ASAP7_75t_L g576 ( 
.A1(n_423),
.A2(n_237),
.B1(n_263),
.B2(n_218),
.Y(n_576)
);

INVxp67_ASAP7_75t_SL g577 ( 
.A(n_437),
.Y(n_577)
);

BUFx10_ASAP7_75t_L g578 ( 
.A(n_479),
.Y(n_578)
);

NOR3xp33_ASAP7_75t_L g579 ( 
.A(n_444),
.B(n_425),
.C(n_412),
.Y(n_579)
);

BUFx6f_ASAP7_75t_L g580 ( 
.A(n_406),
.Y(n_580)
);

NAND2xp5_ASAP7_75t_SL g581 ( 
.A(n_477),
.B(n_173),
.Y(n_581)
);

INVx1_ASAP7_75t_L g582 ( 
.A(n_421),
.Y(n_582)
);

INVx1_ASAP7_75t_L g583 ( 
.A(n_421),
.Y(n_583)
);

INVx1_ASAP7_75t_L g584 ( 
.A(n_421),
.Y(n_584)
);

INVx4_ASAP7_75t_L g585 ( 
.A(n_409),
.Y(n_585)
);

INVx2_ASAP7_75t_L g586 ( 
.A(n_427),
.Y(n_586)
);

AOI22xp33_ASAP7_75t_L g587 ( 
.A1(n_449),
.A2(n_183),
.B1(n_214),
.B2(n_320),
.Y(n_587)
);

INVx1_ASAP7_75t_L g588 ( 
.A(n_424),
.Y(n_588)
);

BUFx3_ASAP7_75t_L g589 ( 
.A(n_457),
.Y(n_589)
);

INVx1_ASAP7_75t_L g590 ( 
.A(n_424),
.Y(n_590)
);

BUFx3_ASAP7_75t_L g591 ( 
.A(n_463),
.Y(n_591)
);

NAND2xp5_ASAP7_75t_L g592 ( 
.A(n_477),
.B(n_318),
.Y(n_592)
);

INVx2_ASAP7_75t_L g593 ( 
.A(n_424),
.Y(n_593)
);

AND2x2_ASAP7_75t_L g594 ( 
.A(n_463),
.B(n_201),
.Y(n_594)
);

INVx1_ASAP7_75t_L g595 ( 
.A(n_428),
.Y(n_595)
);

AO21x2_ASAP7_75t_L g596 ( 
.A1(n_443),
.A2(n_446),
.B(n_453),
.Y(n_596)
);

NAND2xp5_ASAP7_75t_SL g597 ( 
.A(n_477),
.B(n_191),
.Y(n_597)
);

INVx2_ASAP7_75t_L g598 ( 
.A(n_432),
.Y(n_598)
);

AND2x6_ASAP7_75t_L g599 ( 
.A(n_473),
.B(n_179),
.Y(n_599)
);

OR2x2_ASAP7_75t_L g600 ( 
.A(n_444),
.B(n_446),
.Y(n_600)
);

AOI22xp33_ASAP7_75t_L g601 ( 
.A1(n_449),
.A2(n_271),
.B1(n_183),
.B2(n_259),
.Y(n_601)
);

NAND2xp5_ASAP7_75t_SL g602 ( 
.A(n_425),
.B(n_191),
.Y(n_602)
);

NOR2xp33_ASAP7_75t_SL g603 ( 
.A(n_462),
.B(n_328),
.Y(n_603)
);

INVx4_ASAP7_75t_L g604 ( 
.A(n_409),
.Y(n_604)
);

INVx1_ASAP7_75t_L g605 ( 
.A(n_428),
.Y(n_605)
);

AND2x6_ASAP7_75t_L g606 ( 
.A(n_473),
.B(n_264),
.Y(n_606)
);

AOI22xp5_ASAP7_75t_L g607 ( 
.A1(n_423),
.A2(n_296),
.B1(n_302),
.B2(n_239),
.Y(n_607)
);

INVx1_ASAP7_75t_L g608 ( 
.A(n_428),
.Y(n_608)
);

BUFx6f_ASAP7_75t_L g609 ( 
.A(n_407),
.Y(n_609)
);

BUFx10_ASAP7_75t_L g610 ( 
.A(n_449),
.Y(n_610)
);

NOR2xp33_ASAP7_75t_L g611 ( 
.A(n_473),
.B(n_453),
.Y(n_611)
);

AND2x2_ASAP7_75t_L g612 ( 
.A(n_429),
.B(n_203),
.Y(n_612)
);

INVx2_ASAP7_75t_L g613 ( 
.A(n_432),
.Y(n_613)
);

AND2x6_ASAP7_75t_L g614 ( 
.A(n_449),
.B(n_264),
.Y(n_614)
);

INVx2_ASAP7_75t_L g615 ( 
.A(n_432),
.Y(n_615)
);

INVx1_ASAP7_75t_L g616 ( 
.A(n_428),
.Y(n_616)
);

INVx2_ASAP7_75t_L g617 ( 
.A(n_432),
.Y(n_617)
);

AO21x2_ASAP7_75t_L g618 ( 
.A1(n_430),
.A2(n_294),
.B(n_252),
.Y(n_618)
);

INVx2_ASAP7_75t_L g619 ( 
.A(n_434),
.Y(n_619)
);

INVx2_ASAP7_75t_L g620 ( 
.A(n_434),
.Y(n_620)
);

OAI22xp5_ASAP7_75t_L g621 ( 
.A1(n_449),
.A2(n_285),
.B1(n_278),
.B2(n_277),
.Y(n_621)
);

NOR2xp33_ASAP7_75t_L g622 ( 
.A(n_430),
.B(n_331),
.Y(n_622)
);

INVx1_ASAP7_75t_L g623 ( 
.A(n_428),
.Y(n_623)
);

NAND2xp5_ASAP7_75t_L g624 ( 
.A(n_458),
.B(n_323),
.Y(n_624)
);

INVx2_ASAP7_75t_L g625 ( 
.A(n_434),
.Y(n_625)
);

AOI22xp5_ASAP7_75t_L g626 ( 
.A1(n_409),
.A2(n_247),
.B1(n_261),
.B2(n_254),
.Y(n_626)
);

AND3x2_ASAP7_75t_L g627 ( 
.A(n_429),
.B(n_264),
.C(n_175),
.Y(n_627)
);

INVx1_ASAP7_75t_L g628 ( 
.A(n_455),
.Y(n_628)
);

NAND2xp5_ASAP7_75t_SL g629 ( 
.A(n_487),
.B(n_193),
.Y(n_629)
);

NOR2xp33_ASAP7_75t_L g630 ( 
.A(n_565),
.B(n_331),
.Y(n_630)
);

NOR2xp67_ASAP7_75t_L g631 ( 
.A(n_554),
.B(n_455),
.Y(n_631)
);

INVx1_ASAP7_75t_L g632 ( 
.A(n_523),
.Y(n_632)
);

OR2x2_ASAP7_75t_L g633 ( 
.A(n_554),
.B(n_383),
.Y(n_633)
);

INVx1_ASAP7_75t_L g634 ( 
.A(n_523),
.Y(n_634)
);

INVx1_ASAP7_75t_L g635 ( 
.A(n_509),
.Y(n_635)
);

INVx1_ASAP7_75t_L g636 ( 
.A(n_509),
.Y(n_636)
);

INVx1_ASAP7_75t_L g637 ( 
.A(n_513),
.Y(n_637)
);

OR2x2_ASAP7_75t_L g638 ( 
.A(n_600),
.B(n_178),
.Y(n_638)
);

NAND2xp5_ASAP7_75t_L g639 ( 
.A(n_483),
.B(n_458),
.Y(n_639)
);

NAND2xp5_ASAP7_75t_L g640 ( 
.A(n_577),
.B(n_458),
.Y(n_640)
);

OA21x2_ASAP7_75t_L g641 ( 
.A1(n_595),
.A2(n_220),
.B(n_203),
.Y(n_641)
);

NAND2xp5_ASAP7_75t_L g642 ( 
.A(n_611),
.B(n_458),
.Y(n_642)
);

INVx1_ASAP7_75t_L g643 ( 
.A(n_513),
.Y(n_643)
);

INVx1_ASAP7_75t_L g644 ( 
.A(n_514),
.Y(n_644)
);

NOR2xp67_ASAP7_75t_L g645 ( 
.A(n_512),
.B(n_456),
.Y(n_645)
);

NAND2xp5_ASAP7_75t_L g646 ( 
.A(n_565),
.B(n_458),
.Y(n_646)
);

INVx1_ASAP7_75t_L g647 ( 
.A(n_514),
.Y(n_647)
);

INVx1_ASAP7_75t_SL g648 ( 
.A(n_502),
.Y(n_648)
);

BUFx3_ASAP7_75t_L g649 ( 
.A(n_543),
.Y(n_649)
);

NAND2xp33_ASAP7_75t_L g650 ( 
.A(n_599),
.B(n_325),
.Y(n_650)
);

INVx3_ASAP7_75t_L g651 ( 
.A(n_481),
.Y(n_651)
);

NOR2xp33_ASAP7_75t_L g652 ( 
.A(n_600),
.B(n_345),
.Y(n_652)
);

AOI22xp5_ASAP7_75t_L g653 ( 
.A1(n_529),
.A2(n_340),
.B1(n_352),
.B2(n_344),
.Y(n_653)
);

NAND2xp5_ASAP7_75t_SL g654 ( 
.A(n_487),
.B(n_193),
.Y(n_654)
);

NAND2xp5_ASAP7_75t_SL g655 ( 
.A(n_487),
.B(n_193),
.Y(n_655)
);

NAND2xp5_ASAP7_75t_L g656 ( 
.A(n_518),
.B(n_462),
.Y(n_656)
);

AND2x4_ASAP7_75t_L g657 ( 
.A(n_560),
.B(n_456),
.Y(n_657)
);

INVx2_ASAP7_75t_SL g658 ( 
.A(n_502),
.Y(n_658)
);

NAND2xp5_ASAP7_75t_L g659 ( 
.A(n_518),
.B(n_462),
.Y(n_659)
);

INVx2_ASAP7_75t_SL g660 ( 
.A(n_503),
.Y(n_660)
);

OAI22xp5_ASAP7_75t_L g661 ( 
.A1(n_496),
.A2(n_335),
.B1(n_295),
.B2(n_175),
.Y(n_661)
);

INVx1_ASAP7_75t_L g662 ( 
.A(n_560),
.Y(n_662)
);

NAND2xp5_ASAP7_75t_L g663 ( 
.A(n_525),
.B(n_462),
.Y(n_663)
);

OAI22xp5_ASAP7_75t_SL g664 ( 
.A1(n_576),
.A2(n_236),
.B1(n_233),
.B2(n_232),
.Y(n_664)
);

INVx1_ASAP7_75t_L g665 ( 
.A(n_589),
.Y(n_665)
);

INVx8_ASAP7_75t_L g666 ( 
.A(n_599),
.Y(n_666)
);

INVxp67_ASAP7_75t_L g667 ( 
.A(n_568),
.Y(n_667)
);

NAND2xp5_ASAP7_75t_SL g668 ( 
.A(n_529),
.B(n_462),
.Y(n_668)
);

NOR2xp33_ASAP7_75t_L g669 ( 
.A(n_491),
.B(n_345),
.Y(n_669)
);

OR2x2_ASAP7_75t_L g670 ( 
.A(n_503),
.B(n_196),
.Y(n_670)
);

INVxp67_ASAP7_75t_SL g671 ( 
.A(n_568),
.Y(n_671)
);

NAND2xp5_ASAP7_75t_L g672 ( 
.A(n_525),
.B(n_409),
.Y(n_672)
);

INVx1_ASAP7_75t_L g673 ( 
.A(n_589),
.Y(n_673)
);

NAND2xp5_ASAP7_75t_L g674 ( 
.A(n_591),
.B(n_409),
.Y(n_674)
);

NAND2xp5_ASAP7_75t_SL g675 ( 
.A(n_535),
.B(n_326),
.Y(n_675)
);

OR2x6_ASAP7_75t_L g676 ( 
.A(n_535),
.B(n_266),
.Y(n_676)
);

AND2x4_ASAP7_75t_L g677 ( 
.A(n_591),
.B(n_460),
.Y(n_677)
);

INVx2_ASAP7_75t_L g678 ( 
.A(n_500),
.Y(n_678)
);

INVx2_ASAP7_75t_L g679 ( 
.A(n_500),
.Y(n_679)
);

NOR2xp33_ASAP7_75t_L g680 ( 
.A(n_526),
.B(n_548),
.Y(n_680)
);

OAI22xp5_ASAP7_75t_L g681 ( 
.A1(n_492),
.A2(n_187),
.B1(n_295),
.B2(n_220),
.Y(n_681)
);

AOI22xp5_ASAP7_75t_L g682 ( 
.A1(n_596),
.A2(n_409),
.B1(n_345),
.B2(n_227),
.Y(n_682)
);

OR2x2_ASAP7_75t_L g683 ( 
.A(n_536),
.B(n_199),
.Y(n_683)
);

INVx1_ASAP7_75t_L g684 ( 
.A(n_628),
.Y(n_684)
);

AOI22xp33_ASAP7_75t_L g685 ( 
.A1(n_599),
.A2(n_280),
.B1(n_265),
.B2(n_292),
.Y(n_685)
);

OR2x6_ASAP7_75t_L g686 ( 
.A(n_538),
.B(n_223),
.Y(n_686)
);

OR2x2_ASAP7_75t_L g687 ( 
.A(n_536),
.B(n_204),
.Y(n_687)
);

AOI22xp5_ASAP7_75t_L g688 ( 
.A1(n_596),
.A2(n_294),
.B1(n_223),
.B2(n_227),
.Y(n_688)
);

NAND2xp5_ASAP7_75t_L g689 ( 
.A(n_596),
.B(n_231),
.Y(n_689)
);

AO22x2_ASAP7_75t_L g690 ( 
.A1(n_602),
.A2(n_238),
.B1(n_231),
.B2(n_252),
.Y(n_690)
);

BUFx4f_ASAP7_75t_L g691 ( 
.A(n_599),
.Y(n_691)
);

NOR2xp33_ASAP7_75t_L g692 ( 
.A(n_488),
.B(n_499),
.Y(n_692)
);

AND2x2_ASAP7_75t_L g693 ( 
.A(n_533),
.B(n_460),
.Y(n_693)
);

INVx2_ASAP7_75t_L g694 ( 
.A(n_515),
.Y(n_694)
);

INVx2_ASAP7_75t_L g695 ( 
.A(n_515),
.Y(n_695)
);

AOI22xp5_ASAP7_75t_L g696 ( 
.A1(n_516),
.A2(n_238),
.B1(n_265),
.B2(n_280),
.Y(n_696)
);

INVx2_ASAP7_75t_SL g697 ( 
.A(n_594),
.Y(n_697)
);

NOR2xp33_ASAP7_75t_L g698 ( 
.A(n_507),
.B(n_224),
.Y(n_698)
);

NOR2xp33_ASAP7_75t_SL g699 ( 
.A(n_489),
.B(n_191),
.Y(n_699)
);

NAND2xp5_ASAP7_75t_L g700 ( 
.A(n_494),
.B(n_292),
.Y(n_700)
);

INVx3_ASAP7_75t_L g701 ( 
.A(n_481),
.Y(n_701)
);

NOR2xp33_ASAP7_75t_L g702 ( 
.A(n_501),
.B(n_225),
.Y(n_702)
);

AND2x2_ASAP7_75t_L g703 ( 
.A(n_530),
.B(n_208),
.Y(n_703)
);

AOI22xp5_ASAP7_75t_L g704 ( 
.A1(n_579),
.A2(n_305),
.B1(n_327),
.B2(n_187),
.Y(n_704)
);

INVx2_ASAP7_75t_SL g705 ( 
.A(n_594),
.Y(n_705)
);

NAND2xp5_ASAP7_75t_SL g706 ( 
.A(n_508),
.B(n_193),
.Y(n_706)
);

NAND2xp5_ASAP7_75t_L g707 ( 
.A(n_628),
.B(n_305),
.Y(n_707)
);

NAND2xp5_ASAP7_75t_L g708 ( 
.A(n_498),
.B(n_327),
.Y(n_708)
);

INVx1_ASAP7_75t_L g709 ( 
.A(n_485),
.Y(n_709)
);

NAND2xp5_ASAP7_75t_L g710 ( 
.A(n_498),
.B(n_435),
.Y(n_710)
);

BUFx6f_ASAP7_75t_L g711 ( 
.A(n_610),
.Y(n_711)
);

INVx1_ASAP7_75t_L g712 ( 
.A(n_485),
.Y(n_712)
);

NAND2xp5_ASAP7_75t_L g713 ( 
.A(n_498),
.B(n_435),
.Y(n_713)
);

OA22x2_ASAP7_75t_L g714 ( 
.A1(n_607),
.A2(n_306),
.B1(n_226),
.B2(n_274),
.Y(n_714)
);

INVx2_ASAP7_75t_SL g715 ( 
.A(n_530),
.Y(n_715)
);

NAND2xp5_ASAP7_75t_SL g716 ( 
.A(n_508),
.B(n_234),
.Y(n_716)
);

NAND2xp5_ASAP7_75t_L g717 ( 
.A(n_498),
.B(n_435),
.Y(n_717)
);

NAND2xp5_ASAP7_75t_SL g718 ( 
.A(n_508),
.B(n_234),
.Y(n_718)
);

INVx1_ASAP7_75t_L g719 ( 
.A(n_486),
.Y(n_719)
);

NOR2xp33_ASAP7_75t_L g720 ( 
.A(n_553),
.B(n_241),
.Y(n_720)
);

NAND2xp33_ASAP7_75t_L g721 ( 
.A(n_599),
.B(n_234),
.Y(n_721)
);

AOI22xp5_ASAP7_75t_L g722 ( 
.A1(n_506),
.A2(n_433),
.B1(n_461),
.B2(n_450),
.Y(n_722)
);

NAND2xp5_ASAP7_75t_L g723 ( 
.A(n_505),
.B(n_435),
.Y(n_723)
);

INVx1_ASAP7_75t_L g724 ( 
.A(n_486),
.Y(n_724)
);

INVx2_ASAP7_75t_L g725 ( 
.A(n_517),
.Y(n_725)
);

INVx1_ASAP7_75t_L g726 ( 
.A(n_504),
.Y(n_726)
);

INVx1_ASAP7_75t_L g727 ( 
.A(n_504),
.Y(n_727)
);

NAND2xp5_ASAP7_75t_SL g728 ( 
.A(n_530),
.B(n_191),
.Y(n_728)
);

INVx2_ASAP7_75t_L g729 ( 
.A(n_517),
.Y(n_729)
);

AOI22xp33_ASAP7_75t_L g730 ( 
.A1(n_599),
.A2(n_234),
.B1(n_253),
.B2(n_314),
.Y(n_730)
);

NOR2xp33_ASAP7_75t_L g731 ( 
.A(n_563),
.B(n_571),
.Y(n_731)
);

BUFx5_ASAP7_75t_L g732 ( 
.A(n_614),
.Y(n_732)
);

NAND2xp5_ASAP7_75t_L g733 ( 
.A(n_505),
.B(n_435),
.Y(n_733)
);

BUFx6f_ASAP7_75t_L g734 ( 
.A(n_610),
.Y(n_734)
);

NOR2xp33_ASAP7_75t_L g735 ( 
.A(n_592),
.B(n_243),
.Y(n_735)
);

OR2x2_ASAP7_75t_L g736 ( 
.A(n_524),
.B(n_246),
.Y(n_736)
);

NAND2xp5_ASAP7_75t_L g737 ( 
.A(n_505),
.B(n_537),
.Y(n_737)
);

AND2x2_ASAP7_75t_L g738 ( 
.A(n_532),
.B(n_429),
.Y(n_738)
);

NAND2xp5_ASAP7_75t_L g739 ( 
.A(n_505),
.B(n_435),
.Y(n_739)
);

INVxp33_ASAP7_75t_L g740 ( 
.A(n_621),
.Y(n_740)
);

INVx3_ASAP7_75t_L g741 ( 
.A(n_481),
.Y(n_741)
);

AND2x4_ASAP7_75t_L g742 ( 
.A(n_542),
.B(n_431),
.Y(n_742)
);

AND2x2_ASAP7_75t_L g743 ( 
.A(n_532),
.B(n_578),
.Y(n_743)
);

INVx1_ASAP7_75t_L g744 ( 
.A(n_511),
.Y(n_744)
);

INVx2_ASAP7_75t_L g745 ( 
.A(n_520),
.Y(n_745)
);

NAND2xp5_ASAP7_75t_SL g746 ( 
.A(n_508),
.B(n_490),
.Y(n_746)
);

NAND2xp33_ASAP7_75t_L g747 ( 
.A(n_599),
.B(n_234),
.Y(n_747)
);

INVx4_ASAP7_75t_L g748 ( 
.A(n_481),
.Y(n_748)
);

AOI22xp5_ASAP7_75t_L g749 ( 
.A1(n_581),
.A2(n_450),
.B1(n_445),
.B2(n_461),
.Y(n_749)
);

NOR2xp33_ASAP7_75t_SL g750 ( 
.A(n_489),
.B(n_267),
.Y(n_750)
);

NAND2xp5_ASAP7_75t_SL g751 ( 
.A(n_508),
.B(n_253),
.Y(n_751)
);

AND2x4_ASAP7_75t_L g752 ( 
.A(n_542),
.B(n_431),
.Y(n_752)
);

NOR2xp33_ASAP7_75t_L g753 ( 
.A(n_527),
.B(n_269),
.Y(n_753)
);

NOR2xp33_ASAP7_75t_L g754 ( 
.A(n_597),
.B(n_532),
.Y(n_754)
);

NAND2xp5_ASAP7_75t_L g755 ( 
.A(n_537),
.B(n_435),
.Y(n_755)
);

INVx1_ASAP7_75t_L g756 ( 
.A(n_511),
.Y(n_756)
);

BUFx6f_ASAP7_75t_L g757 ( 
.A(n_610),
.Y(n_757)
);

INVx2_ASAP7_75t_L g758 ( 
.A(n_520),
.Y(n_758)
);

AOI22xp33_ASAP7_75t_L g759 ( 
.A1(n_606),
.A2(n_531),
.B1(n_528),
.B2(n_614),
.Y(n_759)
);

NAND2xp5_ASAP7_75t_L g760 ( 
.A(n_537),
.B(n_519),
.Y(n_760)
);

AND2x2_ASAP7_75t_L g761 ( 
.A(n_578),
.B(n_431),
.Y(n_761)
);

INVx2_ASAP7_75t_L g762 ( 
.A(n_521),
.Y(n_762)
);

INVx1_ASAP7_75t_L g763 ( 
.A(n_534),
.Y(n_763)
);

BUFx6f_ASAP7_75t_SL g764 ( 
.A(n_578),
.Y(n_764)
);

NAND2xp5_ASAP7_75t_SL g765 ( 
.A(n_508),
.B(n_490),
.Y(n_765)
);

INVx2_ASAP7_75t_SL g766 ( 
.A(n_542),
.Y(n_766)
);

NOR2xp33_ASAP7_75t_L g767 ( 
.A(n_546),
.B(n_279),
.Y(n_767)
);

INVx2_ASAP7_75t_L g768 ( 
.A(n_521),
.Y(n_768)
);

NAND2xp5_ASAP7_75t_L g769 ( 
.A(n_537),
.B(n_435),
.Y(n_769)
);

NAND2xp5_ASAP7_75t_SL g770 ( 
.A(n_622),
.B(n_253),
.Y(n_770)
);

INVx3_ASAP7_75t_L g771 ( 
.A(n_542),
.Y(n_771)
);

BUFx6f_ASAP7_75t_SL g772 ( 
.A(n_484),
.Y(n_772)
);

A2O1A1Ixp33_ASAP7_75t_L g773 ( 
.A1(n_519),
.A2(n_436),
.B(n_438),
.C(n_461),
.Y(n_773)
);

NAND2xp5_ASAP7_75t_SL g774 ( 
.A(n_626),
.B(n_253),
.Y(n_774)
);

NOR2xp33_ASAP7_75t_L g775 ( 
.A(n_551),
.B(n_281),
.Y(n_775)
);

BUFx6f_ASAP7_75t_L g776 ( 
.A(n_614),
.Y(n_776)
);

AOI22xp33_ASAP7_75t_L g777 ( 
.A1(n_606),
.A2(n_253),
.B1(n_256),
.B2(n_314),
.Y(n_777)
);

NAND2xp5_ASAP7_75t_SL g778 ( 
.A(n_626),
.B(n_256),
.Y(n_778)
);

OAI22xp5_ASAP7_75t_L g779 ( 
.A1(n_545),
.A2(n_256),
.B1(n_314),
.B2(n_283),
.Y(n_779)
);

CKINVDCx5p33_ASAP7_75t_R g780 ( 
.A(n_562),
.Y(n_780)
);

AOI22xp5_ASAP7_75t_L g781 ( 
.A1(n_557),
.A2(n_433),
.B1(n_436),
.B2(n_450),
.Y(n_781)
);

NAND2xp5_ASAP7_75t_L g782 ( 
.A(n_555),
.B(n_435),
.Y(n_782)
);

AND2x2_ASAP7_75t_L g783 ( 
.A(n_564),
.B(n_433),
.Y(n_783)
);

NAND2xp5_ASAP7_75t_SL g784 ( 
.A(n_490),
.B(n_540),
.Y(n_784)
);

AOI22xp33_ASAP7_75t_L g785 ( 
.A1(n_606),
.A2(n_256),
.B1(n_314),
.B2(n_436),
.Y(n_785)
);

NOR2xp33_ASAP7_75t_L g786 ( 
.A(n_573),
.B(n_282),
.Y(n_786)
);

AOI22xp5_ASAP7_75t_L g787 ( 
.A1(n_606),
.A2(n_438),
.B1(n_445),
.B2(n_256),
.Y(n_787)
);

NAND2xp5_ASAP7_75t_SL g788 ( 
.A(n_540),
.B(n_314),
.Y(n_788)
);

AOI22xp33_ASAP7_75t_L g789 ( 
.A1(n_606),
.A2(n_438),
.B1(n_445),
.B2(n_287),
.Y(n_789)
);

INVx2_ASAP7_75t_L g790 ( 
.A(n_522),
.Y(n_790)
);

NAND2xp5_ASAP7_75t_L g791 ( 
.A(n_555),
.B(n_559),
.Y(n_791)
);

NAND2xp5_ASAP7_75t_SL g792 ( 
.A(n_540),
.B(n_439),
.Y(n_792)
);

NAND2xp5_ASAP7_75t_SL g793 ( 
.A(n_585),
.B(n_439),
.Y(n_793)
);

A2O1A1Ixp33_ASAP7_75t_L g794 ( 
.A1(n_559),
.A2(n_465),
.B(n_464),
.C(n_454),
.Y(n_794)
);

AND2x2_ASAP7_75t_L g795 ( 
.A(n_480),
.B(n_284),
.Y(n_795)
);

O2A1O1Ixp5_ASAP7_75t_L g796 ( 
.A1(n_561),
.A2(n_465),
.B(n_464),
.C(n_454),
.Y(n_796)
);

AOI21xp5_ASAP7_75t_L g797 ( 
.A1(n_784),
.A2(n_604),
.B(n_585),
.Y(n_797)
);

NOR2xp33_ASAP7_75t_L g798 ( 
.A(n_692),
.B(n_576),
.Y(n_798)
);

AOI21xp33_ASAP7_75t_L g799 ( 
.A1(n_692),
.A2(n_607),
.B(n_603),
.Y(n_799)
);

BUFx4f_ASAP7_75t_L g800 ( 
.A(n_715),
.Y(n_800)
);

AOI21x1_ASAP7_75t_L g801 ( 
.A1(n_788),
.A2(n_624),
.B(n_561),
.Y(n_801)
);

NOR2x1_ASAP7_75t_L g802 ( 
.A(n_743),
.B(n_618),
.Y(n_802)
);

OAI21xp33_ASAP7_75t_L g803 ( 
.A1(n_786),
.A2(n_552),
.B(n_570),
.Y(n_803)
);

HB1xp67_ASAP7_75t_L g804 ( 
.A(n_667),
.Y(n_804)
);

NAND2xp5_ASAP7_75t_L g805 ( 
.A(n_680),
.B(n_618),
.Y(n_805)
);

NOR2xp33_ASAP7_75t_L g806 ( 
.A(n_667),
.B(n_572),
.Y(n_806)
);

AO21x1_ASAP7_75t_L g807 ( 
.A1(n_774),
.A2(n_778),
.B(n_689),
.Y(n_807)
);

INVx2_ASAP7_75t_L g808 ( 
.A(n_657),
.Y(n_808)
);

AOI21xp5_ASAP7_75t_L g809 ( 
.A1(n_784),
.A2(n_604),
.B(n_585),
.Y(n_809)
);

NAND2xp5_ASAP7_75t_L g810 ( 
.A(n_680),
.B(n_618),
.Y(n_810)
);

INVx2_ASAP7_75t_L g811 ( 
.A(n_657),
.Y(n_811)
);

AOI21xp5_ASAP7_75t_L g812 ( 
.A1(n_760),
.A2(n_604),
.B(n_558),
.Y(n_812)
);

AOI21xp5_ASAP7_75t_L g813 ( 
.A1(n_691),
.A2(n_558),
.B(n_495),
.Y(n_813)
);

NOR2xp33_ASAP7_75t_L g814 ( 
.A(n_671),
.B(n_572),
.Y(n_814)
);

NAND2xp5_ASAP7_75t_L g815 ( 
.A(n_671),
.B(n_574),
.Y(n_815)
);

AOI22xp33_ASAP7_75t_L g816 ( 
.A1(n_661),
.A2(n_606),
.B1(n_484),
.B2(n_566),
.Y(n_816)
);

OAI21xp5_ASAP7_75t_L g817 ( 
.A1(n_672),
.A2(n_595),
.B(n_605),
.Y(n_817)
);

OAI21xp5_ASAP7_75t_L g818 ( 
.A1(n_688),
.A2(n_642),
.B(n_682),
.Y(n_818)
);

AOI21xp5_ASAP7_75t_L g819 ( 
.A1(n_691),
.A2(n_497),
.B(n_495),
.Y(n_819)
);

NAND2xp5_ASAP7_75t_L g820 ( 
.A(n_697),
.B(n_574),
.Y(n_820)
);

O2A1O1Ixp5_ASAP7_75t_L g821 ( 
.A1(n_770),
.A2(n_584),
.B(n_583),
.C(n_582),
.Y(n_821)
);

INVx2_ASAP7_75t_L g822 ( 
.A(n_677),
.Y(n_822)
);

NOR2xp33_ASAP7_75t_L g823 ( 
.A(n_740),
.B(n_582),
.Y(n_823)
);

BUFx6f_ASAP7_75t_L g824 ( 
.A(n_776),
.Y(n_824)
);

AOI21xp5_ASAP7_75t_L g825 ( 
.A1(n_746),
.A2(n_497),
.B(n_580),
.Y(n_825)
);

BUFx4f_ASAP7_75t_L g826 ( 
.A(n_660),
.Y(n_826)
);

INVx1_ASAP7_75t_L g827 ( 
.A(n_677),
.Y(n_827)
);

NAND2xp5_ASAP7_75t_SL g828 ( 
.A(n_732),
.B(n_731),
.Y(n_828)
);

HB1xp67_ASAP7_75t_L g829 ( 
.A(n_676),
.Y(n_829)
);

AOI21xp5_ASAP7_75t_L g830 ( 
.A1(n_746),
.A2(n_497),
.B(n_580),
.Y(n_830)
);

OAI21xp33_ASAP7_75t_L g831 ( 
.A1(n_786),
.A2(n_601),
.B(n_587),
.Y(n_831)
);

NOR2x1_ASAP7_75t_L g832 ( 
.A(n_754),
.B(n_583),
.Y(n_832)
);

A2O1A1Ixp33_ASAP7_75t_L g833 ( 
.A1(n_731),
.A2(n_612),
.B(n_584),
.C(n_590),
.Y(n_833)
);

OAI22xp5_ASAP7_75t_L g834 ( 
.A1(n_759),
.A2(n_590),
.B1(n_588),
.B2(n_623),
.Y(n_834)
);

O2A1O1Ixp5_ASAP7_75t_L g835 ( 
.A1(n_629),
.A2(n_654),
.B(n_655),
.C(n_788),
.Y(n_835)
);

OR2x2_ASAP7_75t_L g836 ( 
.A(n_648),
.B(n_612),
.Y(n_836)
);

NOR2xp67_ASAP7_75t_L g837 ( 
.A(n_658),
.B(n_588),
.Y(n_837)
);

NAND2xp5_ASAP7_75t_L g838 ( 
.A(n_705),
.B(n_606),
.Y(n_838)
);

NOR2xp33_ASAP7_75t_L g839 ( 
.A(n_693),
.B(n_605),
.Y(n_839)
);

AO21x1_ASAP7_75t_L g840 ( 
.A1(n_629),
.A2(n_608),
.B(n_623),
.Y(n_840)
);

OAI22xp33_ASAP7_75t_L g841 ( 
.A1(n_686),
.A2(n_303),
.B1(n_301),
.B2(n_293),
.Y(n_841)
);

BUFx6f_ASAP7_75t_L g842 ( 
.A(n_776),
.Y(n_842)
);

INVx1_ASAP7_75t_L g843 ( 
.A(n_763),
.Y(n_843)
);

OAI21xp5_ASAP7_75t_L g844 ( 
.A1(n_674),
.A2(n_608),
.B(n_616),
.Y(n_844)
);

AND2x2_ASAP7_75t_L g845 ( 
.A(n_703),
.B(n_286),
.Y(n_845)
);

AO21x2_ASAP7_75t_L g846 ( 
.A1(n_654),
.A2(n_593),
.B(n_616),
.Y(n_846)
);

OAI21xp5_ASAP7_75t_L g847 ( 
.A1(n_796),
.A2(n_593),
.B(n_614),
.Y(n_847)
);

INVx1_ASAP7_75t_SL g848 ( 
.A(n_633),
.Y(n_848)
);

NOR2x1p5_ASAP7_75t_L g849 ( 
.A(n_649),
.B(n_291),
.Y(n_849)
);

NAND2xp5_ASAP7_75t_L g850 ( 
.A(n_698),
.B(n_484),
.Y(n_850)
);

AND2x2_ASAP7_75t_L g851 ( 
.A(n_638),
.B(n_308),
.Y(n_851)
);

INVx8_ASAP7_75t_L g852 ( 
.A(n_676),
.Y(n_852)
);

OR2x2_ASAP7_75t_L g853 ( 
.A(n_683),
.B(n_312),
.Y(n_853)
);

NAND2xp5_ASAP7_75t_L g854 ( 
.A(n_698),
.B(n_484),
.Y(n_854)
);

AOI21xp5_ASAP7_75t_L g855 ( 
.A1(n_765),
.A2(n_609),
.B(n_510),
.Y(n_855)
);

AOI21xp5_ASAP7_75t_L g856 ( 
.A1(n_765),
.A2(n_609),
.B(n_510),
.Y(n_856)
);

INVx1_ASAP7_75t_L g857 ( 
.A(n_662),
.Y(n_857)
);

OAI22xp5_ASAP7_75t_L g858 ( 
.A1(n_759),
.A2(n_569),
.B1(n_493),
.B2(n_482),
.Y(n_858)
);

AOI21xp5_ASAP7_75t_L g859 ( 
.A1(n_737),
.A2(n_609),
.B(n_510),
.Y(n_859)
);

NOR2xp33_ASAP7_75t_L g860 ( 
.A(n_687),
.B(n_313),
.Y(n_860)
);

NAND2xp5_ASAP7_75t_SL g861 ( 
.A(n_732),
.B(n_495),
.Y(n_861)
);

INVx1_ASAP7_75t_L g862 ( 
.A(n_665),
.Y(n_862)
);

NAND2xp5_ASAP7_75t_L g863 ( 
.A(n_738),
.B(n_484),
.Y(n_863)
);

O2A1O1Ixp5_ASAP7_75t_L g864 ( 
.A1(n_655),
.A2(n_567),
.B(n_482),
.C(n_493),
.Y(n_864)
);

NAND2xp5_ASAP7_75t_SL g865 ( 
.A(n_732),
.B(n_495),
.Y(n_865)
);

AO21x1_ASAP7_75t_L g866 ( 
.A1(n_681),
.A2(n_598),
.B(n_625),
.Y(n_866)
);

INVx2_ASAP7_75t_L g867 ( 
.A(n_673),
.Y(n_867)
);

OAI22xp5_ASAP7_75t_L g868 ( 
.A1(n_656),
.A2(n_569),
.B1(n_493),
.B2(n_482),
.Y(n_868)
);

AOI21xp5_ASAP7_75t_L g869 ( 
.A1(n_792),
.A2(n_495),
.B(n_556),
.Y(n_869)
);

NAND2xp5_ASAP7_75t_SL g870 ( 
.A(n_732),
.B(n_497),
.Y(n_870)
);

AND2x2_ASAP7_75t_L g871 ( 
.A(n_783),
.B(n_315),
.Y(n_871)
);

NAND2xp5_ASAP7_75t_L g872 ( 
.A(n_761),
.B(n_484),
.Y(n_872)
);

OR2x2_ASAP7_75t_SL g873 ( 
.A(n_736),
.B(n_319),
.Y(n_873)
);

AND2x4_ASAP7_75t_L g874 ( 
.A(n_635),
.B(n_614),
.Y(n_874)
);

INVx2_ASAP7_75t_L g875 ( 
.A(n_636),
.Y(n_875)
);

INVx2_ASAP7_75t_L g876 ( 
.A(n_637),
.Y(n_876)
);

AOI21xp5_ASAP7_75t_L g877 ( 
.A1(n_792),
.A2(n_497),
.B(n_580),
.Y(n_877)
);

NOR2xp33_ASAP7_75t_L g878 ( 
.A(n_643),
.B(n_322),
.Y(n_878)
);

NOR2xp33_ASAP7_75t_L g879 ( 
.A(n_644),
.B(n_647),
.Y(n_879)
);

O2A1O1Ixp33_ASAP7_75t_L g880 ( 
.A1(n_779),
.A2(n_598),
.B(n_625),
.C(n_620),
.Y(n_880)
);

NAND2xp5_ASAP7_75t_L g881 ( 
.A(n_720),
.B(n_484),
.Y(n_881)
);

A2O1A1Ixp33_ASAP7_75t_L g882 ( 
.A1(n_767),
.A2(n_613),
.B(n_620),
.C(n_619),
.Y(n_882)
);

OAI21xp5_ASAP7_75t_L g883 ( 
.A1(n_796),
.A2(n_614),
.B(n_619),
.Y(n_883)
);

AO21x1_ASAP7_75t_L g884 ( 
.A1(n_668),
.A2(n_613),
.B(n_617),
.Y(n_884)
);

AND2x6_ASAP7_75t_L g885 ( 
.A(n_776),
.B(n_711),
.Y(n_885)
);

AOI21xp5_ASAP7_75t_L g886 ( 
.A1(n_793),
.A2(n_609),
.B(n_580),
.Y(n_886)
);

AOI21xp5_ASAP7_75t_L g887 ( 
.A1(n_793),
.A2(n_609),
.B(n_580),
.Y(n_887)
);

NAND2xp5_ASAP7_75t_L g888 ( 
.A(n_720),
.B(n_566),
.Y(n_888)
);

NOR2xp33_ASAP7_75t_L g889 ( 
.A(n_700),
.B(n_567),
.Y(n_889)
);

OAI21xp5_ASAP7_75t_L g890 ( 
.A1(n_646),
.A2(n_614),
.B(n_617),
.Y(n_890)
);

AND2x2_ASAP7_75t_L g891 ( 
.A(n_631),
.B(n_434),
.Y(n_891)
);

AOI22xp5_ASAP7_75t_L g892 ( 
.A1(n_735),
.A2(n_566),
.B1(n_567),
.B2(n_569),
.Y(n_892)
);

AOI21xp5_ASAP7_75t_L g893 ( 
.A1(n_639),
.A2(n_510),
.B(n_556),
.Y(n_893)
);

A2O1A1Ixp33_ASAP7_75t_L g894 ( 
.A1(n_767),
.A2(n_615),
.B(n_447),
.C(n_448),
.Y(n_894)
);

INVx1_ASAP7_75t_SL g895 ( 
.A(n_653),
.Y(n_895)
);

NOR2xp33_ASAP7_75t_L g896 ( 
.A(n_670),
.B(n_615),
.Y(n_896)
);

NOR2xp33_ASAP7_75t_L g897 ( 
.A(n_754),
.B(n_522),
.Y(n_897)
);

NAND2xp5_ASAP7_75t_SL g898 ( 
.A(n_732),
.B(n_510),
.Y(n_898)
);

INVx1_ASAP7_75t_L g899 ( 
.A(n_742),
.Y(n_899)
);

NAND2xp5_ASAP7_75t_SL g900 ( 
.A(n_732),
.B(n_556),
.Y(n_900)
);

O2A1O1Ixp33_ASAP7_75t_L g901 ( 
.A1(n_708),
.A2(n_544),
.B(n_586),
.C(n_575),
.Y(n_901)
);

INVxp33_ASAP7_75t_L g902 ( 
.A(n_775),
.Y(n_902)
);

AOI21xp5_ASAP7_75t_L g903 ( 
.A1(n_640),
.A2(n_556),
.B(n_586),
.Y(n_903)
);

AOI21xp5_ASAP7_75t_L g904 ( 
.A1(n_748),
.A2(n_556),
.B(n_575),
.Y(n_904)
);

AOI21xp5_ASAP7_75t_L g905 ( 
.A1(n_748),
.A2(n_539),
.B(n_550),
.Y(n_905)
);

NAND3xp33_ASAP7_75t_L g906 ( 
.A(n_775),
.B(n_627),
.C(n_454),
.Y(n_906)
);

AOI21xp5_ASAP7_75t_L g907 ( 
.A1(n_721),
.A2(n_550),
.B(n_549),
.Y(n_907)
);

INVx1_ASAP7_75t_SL g908 ( 
.A(n_750),
.Y(n_908)
);

INVx1_ASAP7_75t_L g909 ( 
.A(n_742),
.Y(n_909)
);

AO22x1_ASAP7_75t_L g910 ( 
.A1(n_702),
.A2(n_566),
.B1(n_447),
.B2(n_465),
.Y(n_910)
);

AND2x4_ASAP7_75t_L g911 ( 
.A(n_766),
.B(n_771),
.Y(n_911)
);

INVxp67_ASAP7_75t_L g912 ( 
.A(n_753),
.Y(n_912)
);

AOI21xp5_ASAP7_75t_L g913 ( 
.A1(n_747),
.A2(n_549),
.B(n_547),
.Y(n_913)
);

AND2x2_ASAP7_75t_L g914 ( 
.A(n_652),
.B(n_447),
.Y(n_914)
);

AOI21xp5_ASAP7_75t_L g915 ( 
.A1(n_710),
.A2(n_547),
.B(n_544),
.Y(n_915)
);

AOI21xp5_ASAP7_75t_L g916 ( 
.A1(n_713),
.A2(n_541),
.B(n_539),
.Y(n_916)
);

O2A1O1Ixp33_ASAP7_75t_L g917 ( 
.A1(n_707),
.A2(n_541),
.B(n_465),
.C(n_464),
.Y(n_917)
);

INVx1_ASAP7_75t_L g918 ( 
.A(n_752),
.Y(n_918)
);

NAND2xp33_ASAP7_75t_L g919 ( 
.A(n_711),
.B(n_566),
.Y(n_919)
);

NOR2xp67_ASAP7_75t_L g920 ( 
.A(n_630),
.B(n_70),
.Y(n_920)
);

NAND2xp5_ASAP7_75t_L g921 ( 
.A(n_735),
.B(n_566),
.Y(n_921)
);

INVx2_ASAP7_75t_L g922 ( 
.A(n_752),
.Y(n_922)
);

CKINVDCx5p33_ASAP7_75t_R g923 ( 
.A(n_780),
.Y(n_923)
);

AND2x2_ASAP7_75t_L g924 ( 
.A(n_652),
.B(n_464),
.Y(n_924)
);

AOI21xp5_ASAP7_75t_L g925 ( 
.A1(n_717),
.A2(n_407),
.B(n_454),
.Y(n_925)
);

AOI21xp5_ASAP7_75t_L g926 ( 
.A1(n_723),
.A2(n_739),
.B(n_733),
.Y(n_926)
);

AOI21xp5_ASAP7_75t_L g927 ( 
.A1(n_755),
.A2(n_407),
.B(n_447),
.Y(n_927)
);

NAND2xp5_ASAP7_75t_L g928 ( 
.A(n_684),
.B(n_566),
.Y(n_928)
);

AOI21xp5_ASAP7_75t_L g929 ( 
.A1(n_769),
.A2(n_666),
.B(n_789),
.Y(n_929)
);

AOI21x1_ASAP7_75t_L g930 ( 
.A1(n_791),
.A2(n_448),
.B(n_407),
.Y(n_930)
);

INVxp67_ASAP7_75t_L g931 ( 
.A(n_753),
.Y(n_931)
);

NAND2xp5_ASAP7_75t_L g932 ( 
.A(n_709),
.B(n_448),
.Y(n_932)
);

AOI21xp5_ASAP7_75t_L g933 ( 
.A1(n_666),
.A2(n_407),
.B(n_448),
.Y(n_933)
);

NOR2xp33_ASAP7_75t_L g934 ( 
.A(n_712),
.B(n_5),
.Y(n_934)
);

AOI22xp33_ASAP7_75t_L g935 ( 
.A1(n_685),
.A2(n_439),
.B1(n_451),
.B2(n_407),
.Y(n_935)
);

INVx4_ASAP7_75t_L g936 ( 
.A(n_711),
.Y(n_936)
);

AOI21x1_ASAP7_75t_L g937 ( 
.A1(n_782),
.A2(n_407),
.B(n_422),
.Y(n_937)
);

NAND2xp5_ASAP7_75t_SL g938 ( 
.A(n_711),
.B(n_451),
.Y(n_938)
);

AOI21xp5_ASAP7_75t_L g939 ( 
.A1(n_666),
.A2(n_789),
.B(n_701),
.Y(n_939)
);

NOR2xp33_ASAP7_75t_L g940 ( 
.A(n_719),
.B(n_6),
.Y(n_940)
);

AOI21xp5_ASAP7_75t_L g941 ( 
.A1(n_651),
.A2(n_407),
.B(n_422),
.Y(n_941)
);

CKINVDCx11_ASAP7_75t_R g942 ( 
.A(n_686),
.Y(n_942)
);

BUFx2_ASAP7_75t_L g943 ( 
.A(n_676),
.Y(n_943)
);

AOI21xp5_ASAP7_75t_L g944 ( 
.A1(n_651),
.A2(n_407),
.B(n_422),
.Y(n_944)
);

NAND2xp5_ASAP7_75t_L g945 ( 
.A(n_724),
.B(n_451),
.Y(n_945)
);

BUFx6f_ASAP7_75t_L g946 ( 
.A(n_776),
.Y(n_946)
);

BUFx2_ASAP7_75t_L g947 ( 
.A(n_686),
.Y(n_947)
);

INVx1_ASAP7_75t_L g948 ( 
.A(n_726),
.Y(n_948)
);

NAND2xp5_ASAP7_75t_L g949 ( 
.A(n_727),
.B(n_451),
.Y(n_949)
);

AOI21x1_ASAP7_75t_L g950 ( 
.A1(n_706),
.A2(n_422),
.B(n_416),
.Y(n_950)
);

AOI21xp5_ASAP7_75t_L g951 ( 
.A1(n_701),
.A2(n_422),
.B(n_416),
.Y(n_951)
);

AOI21x1_ASAP7_75t_L g952 ( 
.A1(n_706),
.A2(n_422),
.B(n_416),
.Y(n_952)
);

NAND2xp5_ASAP7_75t_SL g953 ( 
.A(n_734),
.B(n_451),
.Y(n_953)
);

NAND2xp5_ASAP7_75t_L g954 ( 
.A(n_744),
.B(n_451),
.Y(n_954)
);

AOI21xp5_ASAP7_75t_L g955 ( 
.A1(n_741),
.A2(n_771),
.B(n_650),
.Y(n_955)
);

NOR2xp33_ASAP7_75t_L g956 ( 
.A(n_756),
.B(n_702),
.Y(n_956)
);

NAND2xp5_ASAP7_75t_L g957 ( 
.A(n_669),
.B(n_451),
.Y(n_957)
);

AOI21xp5_ASAP7_75t_L g958 ( 
.A1(n_741),
.A2(n_422),
.B(n_416),
.Y(n_958)
);

OAI321xp33_ASAP7_75t_L g959 ( 
.A1(n_664),
.A2(n_451),
.A3(n_439),
.B1(n_10),
.B2(n_11),
.C(n_14),
.Y(n_959)
);

INVx1_ASAP7_75t_SL g960 ( 
.A(n_714),
.Y(n_960)
);

BUFx12f_ASAP7_75t_L g961 ( 
.A(n_795),
.Y(n_961)
);

A2O1A1Ixp33_ASAP7_75t_L g962 ( 
.A1(n_696),
.A2(n_451),
.B(n_439),
.C(n_422),
.Y(n_962)
);

NAND2xp33_ASAP7_75t_L g963 ( 
.A(n_734),
.B(n_439),
.Y(n_963)
);

AND2x2_ASAP7_75t_L g964 ( 
.A(n_630),
.B(n_439),
.Y(n_964)
);

OR2x2_ASAP7_75t_L g965 ( 
.A(n_675),
.B(n_8),
.Y(n_965)
);

NAND2xp5_ASAP7_75t_L g966 ( 
.A(n_669),
.B(n_439),
.Y(n_966)
);

AOI21xp33_ASAP7_75t_L g967 ( 
.A1(n_659),
.A2(n_663),
.B(n_714),
.Y(n_967)
);

INVx1_ASAP7_75t_L g968 ( 
.A(n_632),
.Y(n_968)
);

NAND2xp5_ASAP7_75t_L g969 ( 
.A(n_722),
.B(n_439),
.Y(n_969)
);

OAI21xp5_ASAP7_75t_L g970 ( 
.A1(n_773),
.A2(n_422),
.B(n_416),
.Y(n_970)
);

O2A1O1Ixp33_ASAP7_75t_L g971 ( 
.A1(n_634),
.A2(n_9),
.B(n_10),
.C(n_11),
.Y(n_971)
);

NAND2xp5_ASAP7_75t_SL g972 ( 
.A(n_734),
.B(n_416),
.Y(n_972)
);

AND2x2_ASAP7_75t_L g973 ( 
.A(n_699),
.B(n_14),
.Y(n_973)
);

INVx3_ASAP7_75t_L g974 ( 
.A(n_734),
.Y(n_974)
);

BUFx2_ASAP7_75t_L g975 ( 
.A(n_690),
.Y(n_975)
);

OAI21xp5_ASAP7_75t_L g976 ( 
.A1(n_678),
.A2(n_416),
.B(n_415),
.Y(n_976)
);

AOI21xp5_ASAP7_75t_L g977 ( 
.A1(n_785),
.A2(n_416),
.B(n_415),
.Y(n_977)
);

INVx1_ASAP7_75t_L g978 ( 
.A(n_679),
.Y(n_978)
);

AOI22xp5_ASAP7_75t_L g979 ( 
.A1(n_645),
.A2(n_416),
.B1(n_415),
.B2(n_413),
.Y(n_979)
);

AOI21xp5_ASAP7_75t_L g980 ( 
.A1(n_785),
.A2(n_415),
.B(n_413),
.Y(n_980)
);

INVx1_ASAP7_75t_L g981 ( 
.A(n_694),
.Y(n_981)
);

INVx1_ASAP7_75t_L g982 ( 
.A(n_695),
.Y(n_982)
);

NAND2xp5_ASAP7_75t_L g983 ( 
.A(n_781),
.B(n_415),
.Y(n_983)
);

NAND2xp5_ASAP7_75t_L g984 ( 
.A(n_757),
.B(n_415),
.Y(n_984)
);

AND2x4_ASAP7_75t_L g985 ( 
.A(n_808),
.B(n_811),
.Y(n_985)
);

OR2x2_ASAP7_75t_L g986 ( 
.A(n_848),
.B(n_728),
.Y(n_986)
);

NOR2xp33_ASAP7_75t_L g987 ( 
.A(n_902),
.B(n_764),
.Y(n_987)
);

NAND2x1p5_ASAP7_75t_L g988 ( 
.A(n_936),
.B(n_757),
.Y(n_988)
);

NOR2xp33_ASAP7_75t_L g989 ( 
.A(n_912),
.B(n_764),
.Y(n_989)
);

CKINVDCx20_ASAP7_75t_R g990 ( 
.A(n_923),
.Y(n_990)
);

INVx4_ASAP7_75t_L g991 ( 
.A(n_824),
.Y(n_991)
);

AND2x2_ASAP7_75t_L g992 ( 
.A(n_871),
.B(n_690),
.Y(n_992)
);

AOI21xp5_ASAP7_75t_L g993 ( 
.A1(n_797),
.A2(n_757),
.B(n_777),
.Y(n_993)
);

AND2x2_ASAP7_75t_SL g994 ( 
.A(n_798),
.B(n_730),
.Y(n_994)
);

OAI22xp5_ASAP7_75t_L g995 ( 
.A1(n_798),
.A2(n_777),
.B1(n_730),
.B2(n_685),
.Y(n_995)
);

NAND2xp33_ASAP7_75t_L g996 ( 
.A(n_885),
.B(n_757),
.Y(n_996)
);

NOR2xp33_ASAP7_75t_L g997 ( 
.A(n_931),
.B(n_704),
.Y(n_997)
);

NAND2xp5_ASAP7_75t_SL g998 ( 
.A(n_956),
.B(n_749),
.Y(n_998)
);

AOI22xp33_ASAP7_75t_L g999 ( 
.A1(n_803),
.A2(n_690),
.B1(n_772),
.B2(n_745),
.Y(n_999)
);

AND2x4_ASAP7_75t_L g1000 ( 
.A(n_822),
.B(n_758),
.Y(n_1000)
);

AND2x2_ASAP7_75t_L g1001 ( 
.A(n_836),
.B(n_641),
.Y(n_1001)
);

INVx3_ASAP7_75t_SL g1002 ( 
.A(n_908),
.Y(n_1002)
);

AOI21xp5_ASAP7_75t_L g1003 ( 
.A1(n_809),
.A2(n_718),
.B(n_751),
.Y(n_1003)
);

NAND2xp5_ASAP7_75t_L g1004 ( 
.A(n_956),
.B(n_729),
.Y(n_1004)
);

INVxp67_ASAP7_75t_L g1005 ( 
.A(n_860),
.Y(n_1005)
);

INVx1_ASAP7_75t_L g1006 ( 
.A(n_804),
.Y(n_1006)
);

AOI221xp5_ASAP7_75t_L g1007 ( 
.A1(n_799),
.A2(n_841),
.B1(n_831),
.B2(n_860),
.C(n_959),
.Y(n_1007)
);

A2O1A1Ixp33_ASAP7_75t_L g1008 ( 
.A1(n_823),
.A2(n_818),
.B(n_967),
.C(n_896),
.Y(n_1008)
);

O2A1O1Ixp33_ASAP7_75t_L g1009 ( 
.A1(n_841),
.A2(n_794),
.B(n_751),
.C(n_718),
.Y(n_1009)
);

OAI21x1_ASAP7_75t_L g1010 ( 
.A1(n_937),
.A2(n_790),
.B(n_725),
.Y(n_1010)
);

HB1xp67_ASAP7_75t_L g1011 ( 
.A(n_804),
.Y(n_1011)
);

INVx1_ASAP7_75t_L g1012 ( 
.A(n_948),
.Y(n_1012)
);

INVx6_ASAP7_75t_L g1013 ( 
.A(n_936),
.Y(n_1013)
);

NOR2xp33_ASAP7_75t_L g1014 ( 
.A(n_895),
.B(n_768),
.Y(n_1014)
);

O2A1O1Ixp33_ASAP7_75t_L g1015 ( 
.A1(n_823),
.A2(n_716),
.B(n_762),
.C(n_641),
.Y(n_1015)
);

NAND2xp5_ASAP7_75t_L g1016 ( 
.A(n_839),
.B(n_641),
.Y(n_1016)
);

AOI21xp5_ASAP7_75t_L g1017 ( 
.A1(n_939),
.A2(n_716),
.B(n_787),
.Y(n_1017)
);

NAND2xp5_ASAP7_75t_L g1018 ( 
.A(n_839),
.B(n_413),
.Y(n_1018)
);

O2A1O1Ixp5_ASAP7_75t_L g1019 ( 
.A1(n_866),
.A2(n_772),
.B(n_66),
.C(n_68),
.Y(n_1019)
);

NAND2xp5_ASAP7_75t_L g1020 ( 
.A(n_814),
.B(n_415),
.Y(n_1020)
);

OR2x6_ASAP7_75t_SL g1021 ( 
.A(n_965),
.B(n_16),
.Y(n_1021)
);

INVx4_ASAP7_75t_L g1022 ( 
.A(n_824),
.Y(n_1022)
);

AOI22xp5_ASAP7_75t_L g1023 ( 
.A1(n_827),
.A2(n_415),
.B1(n_413),
.B2(n_63),
.Y(n_1023)
);

AOI21xp5_ASAP7_75t_L g1024 ( 
.A1(n_828),
.A2(n_415),
.B(n_413),
.Y(n_1024)
);

OAI22xp5_ASAP7_75t_L g1025 ( 
.A1(n_814),
.A2(n_413),
.B1(n_18),
.B2(n_19),
.Y(n_1025)
);

O2A1O1Ixp33_ASAP7_75t_SL g1026 ( 
.A1(n_828),
.A2(n_160),
.B(n_159),
.C(n_143),
.Y(n_1026)
);

AOI22xp5_ASAP7_75t_L g1027 ( 
.A1(n_845),
.A2(n_413),
.B1(n_137),
.B2(n_134),
.Y(n_1027)
);

INVx1_ASAP7_75t_SL g1028 ( 
.A(n_960),
.Y(n_1028)
);

NAND2xp5_ASAP7_75t_SL g1029 ( 
.A(n_922),
.B(n_413),
.Y(n_1029)
);

NOR2xp33_ASAP7_75t_L g1030 ( 
.A(n_943),
.B(n_16),
.Y(n_1030)
);

OAI21x1_ASAP7_75t_L g1031 ( 
.A1(n_930),
.A2(n_115),
.B(n_133),
.Y(n_1031)
);

INVx4_ASAP7_75t_L g1032 ( 
.A(n_824),
.Y(n_1032)
);

INVxp67_ASAP7_75t_L g1033 ( 
.A(n_853),
.Y(n_1033)
);

AOI21xp5_ASAP7_75t_L g1034 ( 
.A1(n_955),
.A2(n_413),
.B(n_131),
.Y(n_1034)
);

NAND2xp5_ASAP7_75t_L g1035 ( 
.A(n_806),
.B(n_21),
.Y(n_1035)
);

BUFx8_ASAP7_75t_L g1036 ( 
.A(n_961),
.Y(n_1036)
);

NAND2xp5_ASAP7_75t_L g1037 ( 
.A(n_806),
.B(n_22),
.Y(n_1037)
);

HB1xp67_ASAP7_75t_L g1038 ( 
.A(n_829),
.Y(n_1038)
);

AND2x2_ASAP7_75t_L g1039 ( 
.A(n_851),
.B(n_23),
.Y(n_1039)
);

AND2x4_ASAP7_75t_SL g1040 ( 
.A(n_974),
.B(n_127),
.Y(n_1040)
);

INVx1_ASAP7_75t_L g1041 ( 
.A(n_843),
.Y(n_1041)
);

AOI22xp33_ASAP7_75t_SL g1042 ( 
.A1(n_973),
.A2(n_25),
.B1(n_26),
.B2(n_27),
.Y(n_1042)
);

AOI21xp5_ASAP7_75t_L g1043 ( 
.A1(n_812),
.A2(n_124),
.B(n_117),
.Y(n_1043)
);

OAI22xp5_ASAP7_75t_L g1044 ( 
.A1(n_815),
.A2(n_26),
.B1(n_29),
.B2(n_30),
.Y(n_1044)
);

O2A1O1Ixp33_ASAP7_75t_SL g1045 ( 
.A1(n_833),
.A2(n_92),
.B(n_84),
.C(n_83),
.Y(n_1045)
);

NAND2xp5_ASAP7_75t_L g1046 ( 
.A(n_896),
.B(n_31),
.Y(n_1046)
);

OAI22x1_ASAP7_75t_L g1047 ( 
.A1(n_947),
.A2(n_32),
.B1(n_39),
.B2(n_42),
.Y(n_1047)
);

NOR2xp33_ASAP7_75t_L g1048 ( 
.A(n_867),
.B(n_32),
.Y(n_1048)
);

NAND2xp5_ASAP7_75t_L g1049 ( 
.A(n_805),
.B(n_39),
.Y(n_1049)
);

NAND2xp5_ASAP7_75t_L g1050 ( 
.A(n_810),
.B(n_42),
.Y(n_1050)
);

INVx6_ASAP7_75t_L g1051 ( 
.A(n_852),
.Y(n_1051)
);

AOI21xp5_ASAP7_75t_L g1052 ( 
.A1(n_929),
.A2(n_75),
.B(n_72),
.Y(n_1052)
);

AOI22xp33_ASAP7_75t_L g1053 ( 
.A1(n_975),
.A2(n_43),
.B1(n_45),
.B2(n_46),
.Y(n_1053)
);

NAND2xp5_ASAP7_75t_L g1054 ( 
.A(n_897),
.B(n_71),
.Y(n_1054)
);

OAI22xp5_ASAP7_75t_L g1055 ( 
.A1(n_833),
.A2(n_51),
.B1(n_59),
.B2(n_834),
.Y(n_1055)
);

OAI22xp5_ASAP7_75t_L g1056 ( 
.A1(n_816),
.A2(n_51),
.B1(n_940),
.B2(n_934),
.Y(n_1056)
);

NAND2xp5_ASAP7_75t_L g1057 ( 
.A(n_820),
.B(n_879),
.Y(n_1057)
);

AOI21x1_ASAP7_75t_L g1058 ( 
.A1(n_938),
.A2(n_953),
.B(n_801),
.Y(n_1058)
);

INVx4_ASAP7_75t_L g1059 ( 
.A(n_824),
.Y(n_1059)
);

NAND2xp5_ASAP7_75t_SL g1060 ( 
.A(n_911),
.B(n_837),
.Y(n_1060)
);

NAND2xp5_ASAP7_75t_L g1061 ( 
.A(n_879),
.B(n_897),
.Y(n_1061)
);

NAND2xp5_ASAP7_75t_L g1062 ( 
.A(n_832),
.B(n_934),
.Y(n_1062)
);

INVx2_ASAP7_75t_L g1063 ( 
.A(n_875),
.Y(n_1063)
);

OAI21xp5_ASAP7_75t_L g1064 ( 
.A1(n_926),
.A2(n_835),
.B(n_882),
.Y(n_1064)
);

CKINVDCx8_ASAP7_75t_R g1065 ( 
.A(n_852),
.Y(n_1065)
);

NAND2xp5_ASAP7_75t_L g1066 ( 
.A(n_940),
.B(n_914),
.Y(n_1066)
);

NAND2xp5_ASAP7_75t_L g1067 ( 
.A(n_924),
.B(n_889),
.Y(n_1067)
);

INVx4_ASAP7_75t_L g1068 ( 
.A(n_842),
.Y(n_1068)
);

BUFx3_ASAP7_75t_L g1069 ( 
.A(n_826),
.Y(n_1069)
);

NAND2xp5_ASAP7_75t_L g1070 ( 
.A(n_889),
.B(n_891),
.Y(n_1070)
);

NOR2xp33_ASAP7_75t_L g1071 ( 
.A(n_876),
.B(n_857),
.Y(n_1071)
);

NAND2xp33_ASAP7_75t_L g1072 ( 
.A(n_885),
.B(n_842),
.Y(n_1072)
);

INVx4_ASAP7_75t_L g1073 ( 
.A(n_842),
.Y(n_1073)
);

AOI22xp33_ASAP7_75t_L g1074 ( 
.A1(n_899),
.A2(n_909),
.B1(n_918),
.B2(n_911),
.Y(n_1074)
);

OAI22xp5_ASAP7_75t_L g1075 ( 
.A1(n_816),
.A2(n_873),
.B1(n_842),
.B2(n_946),
.Y(n_1075)
);

NAND2x1p5_ASAP7_75t_L g1076 ( 
.A(n_974),
.B(n_946),
.Y(n_1076)
);

NOR2xp67_ASAP7_75t_L g1077 ( 
.A(n_906),
.B(n_878),
.Y(n_1077)
);

NOR2xp33_ASAP7_75t_L g1078 ( 
.A(n_862),
.B(n_878),
.Y(n_1078)
);

O2A1O1Ixp33_ASAP7_75t_L g1079 ( 
.A1(n_971),
.A2(n_968),
.B(n_894),
.C(n_882),
.Y(n_1079)
);

AOI22xp5_ASAP7_75t_L g1080 ( 
.A1(n_874),
.A2(n_802),
.B1(n_920),
.B2(n_863),
.Y(n_1080)
);

OAI22xp5_ASAP7_75t_L g1081 ( 
.A1(n_946),
.A2(n_872),
.B1(n_921),
.B2(n_888),
.Y(n_1081)
);

AND2x6_ASAP7_75t_L g1082 ( 
.A(n_946),
.B(n_874),
.Y(n_1082)
);

AOI21xp5_ASAP7_75t_L g1083 ( 
.A1(n_861),
.A2(n_898),
.B(n_865),
.Y(n_1083)
);

AOI21xp5_ASAP7_75t_L g1084 ( 
.A1(n_861),
.A2(n_870),
.B(n_865),
.Y(n_1084)
);

BUFx4f_ASAP7_75t_L g1085 ( 
.A(n_852),
.Y(n_1085)
);

A2O1A1Ixp33_ASAP7_75t_L g1086 ( 
.A1(n_850),
.A2(n_854),
.B(n_881),
.C(n_838),
.Y(n_1086)
);

AOI21xp5_ASAP7_75t_L g1087 ( 
.A1(n_870),
.A2(n_900),
.B(n_898),
.Y(n_1087)
);

AOI22xp5_ASAP7_75t_L g1088 ( 
.A1(n_807),
.A2(n_964),
.B1(n_982),
.B2(n_981),
.Y(n_1088)
);

OAI21xp33_ASAP7_75t_SL g1089 ( 
.A1(n_847),
.A2(n_900),
.B(n_844),
.Y(n_1089)
);

INVx2_ASAP7_75t_L g1090 ( 
.A(n_978),
.Y(n_1090)
);

HB1xp67_ASAP7_75t_L g1091 ( 
.A(n_826),
.Y(n_1091)
);

AOI22xp33_ASAP7_75t_L g1092 ( 
.A1(n_928),
.A2(n_969),
.B1(n_840),
.B2(n_932),
.Y(n_1092)
);

AOI22xp33_ASAP7_75t_L g1093 ( 
.A1(n_884),
.A2(n_890),
.B1(n_846),
.B2(n_983),
.Y(n_1093)
);

BUFx4f_ASAP7_75t_L g1094 ( 
.A(n_885),
.Y(n_1094)
);

INVxp67_ASAP7_75t_L g1095 ( 
.A(n_849),
.Y(n_1095)
);

INVx3_ASAP7_75t_L g1096 ( 
.A(n_885),
.Y(n_1096)
);

AO32x2_ASAP7_75t_L g1097 ( 
.A1(n_868),
.A2(n_858),
.A3(n_894),
.B1(n_846),
.B2(n_821),
.Y(n_1097)
);

NOR2xp33_ASAP7_75t_L g1098 ( 
.A(n_800),
.B(n_942),
.Y(n_1098)
);

INVx4_ASAP7_75t_L g1099 ( 
.A(n_885),
.Y(n_1099)
);

NAND2xp5_ASAP7_75t_L g1100 ( 
.A(n_817),
.B(n_957),
.Y(n_1100)
);

OAI22xp5_ASAP7_75t_L g1101 ( 
.A1(n_892),
.A2(n_962),
.B1(n_813),
.B2(n_800),
.Y(n_1101)
);

CKINVDCx5p33_ASAP7_75t_R g1102 ( 
.A(n_966),
.Y(n_1102)
);

O2A1O1Ixp33_ASAP7_75t_L g1103 ( 
.A1(n_962),
.A2(n_949),
.B(n_954),
.C(n_945),
.Y(n_1103)
);

INVx1_ASAP7_75t_SL g1104 ( 
.A(n_938),
.Y(n_1104)
);

NAND2xp5_ASAP7_75t_SL g1105 ( 
.A(n_859),
.B(n_953),
.Y(n_1105)
);

INVx1_ASAP7_75t_L g1106 ( 
.A(n_880),
.Y(n_1106)
);

NAND2xp5_ASAP7_75t_L g1107 ( 
.A(n_893),
.B(n_903),
.Y(n_1107)
);

AOI22xp33_ASAP7_75t_L g1108 ( 
.A1(n_883),
.A2(n_972),
.B1(n_919),
.B2(n_916),
.Y(n_1108)
);

AOI22xp5_ASAP7_75t_L g1109 ( 
.A1(n_972),
.A2(n_963),
.B1(n_910),
.B2(n_979),
.Y(n_1109)
);

NAND2xp5_ASAP7_75t_SL g1110 ( 
.A(n_984),
.B(n_877),
.Y(n_1110)
);

INVx1_ASAP7_75t_L g1111 ( 
.A(n_901),
.Y(n_1111)
);

NAND2xp5_ASAP7_75t_L g1112 ( 
.A(n_915),
.B(n_925),
.Y(n_1112)
);

O2A1O1Ixp33_ASAP7_75t_L g1113 ( 
.A1(n_917),
.A2(n_864),
.B(n_970),
.C(n_976),
.Y(n_1113)
);

A2O1A1Ixp33_ASAP7_75t_L g1114 ( 
.A1(n_927),
.A2(n_887),
.B(n_886),
.C(n_869),
.Y(n_1114)
);

INVx2_ASAP7_75t_L g1115 ( 
.A(n_950),
.Y(n_1115)
);

OAI21xp33_ASAP7_75t_L g1116 ( 
.A1(n_935),
.A2(n_977),
.B(n_980),
.Y(n_1116)
);

O2A1O1Ixp33_ASAP7_75t_L g1117 ( 
.A1(n_907),
.A2(n_913),
.B(n_905),
.C(n_904),
.Y(n_1117)
);

NAND2xp5_ASAP7_75t_L g1118 ( 
.A(n_825),
.B(n_830),
.Y(n_1118)
);

AOI21xp5_ASAP7_75t_L g1119 ( 
.A1(n_819),
.A2(n_855),
.B(n_856),
.Y(n_1119)
);

NAND2xp5_ASAP7_75t_L g1120 ( 
.A(n_951),
.B(n_958),
.Y(n_1120)
);

INVx3_ASAP7_75t_L g1121 ( 
.A(n_952),
.Y(n_1121)
);

AND2x2_ASAP7_75t_L g1122 ( 
.A(n_935),
.B(n_941),
.Y(n_1122)
);

NAND2xp5_ASAP7_75t_SL g1123 ( 
.A(n_933),
.B(n_944),
.Y(n_1123)
);

INVx1_ASAP7_75t_L g1124 ( 
.A(n_804),
.Y(n_1124)
);

HB1xp67_ASAP7_75t_L g1125 ( 
.A(n_804),
.Y(n_1125)
);

NAND2xp5_ASAP7_75t_SL g1126 ( 
.A(n_912),
.B(n_931),
.Y(n_1126)
);

OAI21xp5_ASAP7_75t_L g1127 ( 
.A1(n_926),
.A2(n_818),
.B(n_835),
.Y(n_1127)
);

AND2x4_ASAP7_75t_L g1128 ( 
.A(n_808),
.B(n_811),
.Y(n_1128)
);

NOR2xp33_ASAP7_75t_L g1129 ( 
.A(n_902),
.B(n_912),
.Y(n_1129)
);

AOI21xp5_ASAP7_75t_L g1130 ( 
.A1(n_797),
.A2(n_784),
.B(n_691),
.Y(n_1130)
);

OAI21xp5_ASAP7_75t_L g1131 ( 
.A1(n_926),
.A2(n_818),
.B(n_835),
.Y(n_1131)
);

NAND2x1p5_ASAP7_75t_L g1132 ( 
.A(n_936),
.B(n_974),
.Y(n_1132)
);

NOR2xp33_ASAP7_75t_L g1133 ( 
.A(n_902),
.B(n_912),
.Y(n_1133)
);

O2A1O1Ixp33_ASAP7_75t_L g1134 ( 
.A1(n_1005),
.A2(n_1056),
.B(n_998),
.C(n_1008),
.Y(n_1134)
);

OAI21x1_ASAP7_75t_L g1135 ( 
.A1(n_1010),
.A2(n_1119),
.B(n_1117),
.Y(n_1135)
);

A2O1A1Ixp33_ASAP7_75t_L g1136 ( 
.A1(n_1007),
.A2(n_997),
.B(n_1077),
.C(n_995),
.Y(n_1136)
);

OAI21x1_ASAP7_75t_L g1137 ( 
.A1(n_1024),
.A2(n_1107),
.B(n_1058),
.Y(n_1137)
);

O2A1O1Ixp33_ASAP7_75t_L g1138 ( 
.A1(n_1056),
.A2(n_1126),
.B(n_1055),
.C(n_1062),
.Y(n_1138)
);

AOI21xp5_ASAP7_75t_L g1139 ( 
.A1(n_1130),
.A2(n_993),
.B(n_1127),
.Y(n_1139)
);

O2A1O1Ixp5_ASAP7_75t_SL g1140 ( 
.A1(n_1025),
.A2(n_1055),
.B(n_1044),
.C(n_1105),
.Y(n_1140)
);

NAND2xp5_ASAP7_75t_SL g1141 ( 
.A(n_1129),
.B(n_1133),
.Y(n_1141)
);

OAI21xp5_ASAP7_75t_L g1142 ( 
.A1(n_1089),
.A2(n_1086),
.B(n_1127),
.Y(n_1142)
);

AND2x4_ASAP7_75t_L g1143 ( 
.A(n_985),
.B(n_1128),
.Y(n_1143)
);

CKINVDCx8_ASAP7_75t_R g1144 ( 
.A(n_1098),
.Y(n_1144)
);

AO31x2_ASAP7_75t_L g1145 ( 
.A1(n_1101),
.A2(n_1114),
.A3(n_1081),
.B(n_1107),
.Y(n_1145)
);

NAND2xp5_ASAP7_75t_L g1146 ( 
.A(n_1061),
.B(n_1057),
.Y(n_1146)
);

AO31x2_ASAP7_75t_L g1147 ( 
.A1(n_1101),
.A2(n_1081),
.A3(n_1100),
.B(n_1016),
.Y(n_1147)
);

OR2x6_ASAP7_75t_L g1148 ( 
.A(n_1051),
.B(n_1013),
.Y(n_1148)
);

AOI21xp5_ASAP7_75t_L g1149 ( 
.A1(n_1131),
.A2(n_996),
.B(n_1100),
.Y(n_1149)
);

AOI221xp5_ASAP7_75t_L g1150 ( 
.A1(n_1025),
.A2(n_1044),
.B1(n_1078),
.B2(n_1033),
.C(n_995),
.Y(n_1150)
);

NAND2xp5_ASAP7_75t_SL g1151 ( 
.A(n_986),
.B(n_1014),
.Y(n_1151)
);

INVx1_ASAP7_75t_L g1152 ( 
.A(n_1041),
.Y(n_1152)
);

CKINVDCx11_ASAP7_75t_R g1153 ( 
.A(n_990),
.Y(n_1153)
);

AOI221x1_ASAP7_75t_L g1154 ( 
.A1(n_1131),
.A2(n_1064),
.B1(n_1052),
.B2(n_1050),
.C(n_1049),
.Y(n_1154)
);

AO31x2_ASAP7_75t_L g1155 ( 
.A1(n_1111),
.A2(n_1118),
.A3(n_1112),
.B(n_1054),
.Y(n_1155)
);

AOI21xp5_ASAP7_75t_L g1156 ( 
.A1(n_1067),
.A2(n_1070),
.B(n_1064),
.Y(n_1156)
);

NAND2xp5_ASAP7_75t_L g1157 ( 
.A(n_1066),
.B(n_994),
.Y(n_1157)
);

O2A1O1Ixp33_ASAP7_75t_SL g1158 ( 
.A1(n_1054),
.A2(n_1035),
.B(n_1037),
.C(n_1075),
.Y(n_1158)
);

AOI21xp5_ASAP7_75t_L g1159 ( 
.A1(n_1067),
.A2(n_1070),
.B(n_1123),
.Y(n_1159)
);

AOI221x1_ASAP7_75t_L g1160 ( 
.A1(n_1046),
.A2(n_1075),
.B1(n_1017),
.B2(n_1034),
.C(n_1116),
.Y(n_1160)
);

HB1xp67_ASAP7_75t_L g1161 ( 
.A(n_1011),
.Y(n_1161)
);

AOI22xp5_ASAP7_75t_L g1162 ( 
.A1(n_992),
.A2(n_1048),
.B1(n_1039),
.B2(n_1071),
.Y(n_1162)
);

INVx2_ASAP7_75t_L g1163 ( 
.A(n_1090),
.Y(n_1163)
);

A2O1A1Ixp33_ASAP7_75t_L g1164 ( 
.A1(n_1079),
.A2(n_1027),
.B(n_1080),
.C(n_1009),
.Y(n_1164)
);

OAI21x1_ASAP7_75t_L g1165 ( 
.A1(n_1083),
.A2(n_1084),
.B(n_1087),
.Y(n_1165)
);

AOI21xp5_ASAP7_75t_L g1166 ( 
.A1(n_1120),
.A2(n_1110),
.B(n_1072),
.Y(n_1166)
);

AOI21x1_ASAP7_75t_SL g1167 ( 
.A1(n_1004),
.A2(n_1020),
.B(n_1122),
.Y(n_1167)
);

AO31x2_ASAP7_75t_L g1168 ( 
.A1(n_1106),
.A2(n_1018),
.A3(n_1115),
.B(n_1003),
.Y(n_1168)
);

OAI22xp33_ASAP7_75t_L g1169 ( 
.A1(n_1021),
.A2(n_1028),
.B1(n_1102),
.B2(n_1091),
.Y(n_1169)
);

AOI21x1_ASAP7_75t_L g1170 ( 
.A1(n_1043),
.A2(n_1029),
.B(n_1001),
.Y(n_1170)
);

AOI21xp5_ASAP7_75t_L g1171 ( 
.A1(n_1113),
.A2(n_1108),
.B(n_1103),
.Y(n_1171)
);

NOR2x1_ASAP7_75t_L g1172 ( 
.A(n_1069),
.B(n_1124),
.Y(n_1172)
);

AOI21xp5_ASAP7_75t_L g1173 ( 
.A1(n_1015),
.A2(n_1094),
.B(n_1093),
.Y(n_1173)
);

AOI21xp5_ASAP7_75t_L g1174 ( 
.A1(n_1094),
.A2(n_1092),
.B(n_1109),
.Y(n_1174)
);

OR2x2_ASAP7_75t_L g1175 ( 
.A(n_1125),
.B(n_1006),
.Y(n_1175)
);

BUFx6f_ASAP7_75t_L g1176 ( 
.A(n_1051),
.Y(n_1176)
);

INVxp67_ASAP7_75t_L g1177 ( 
.A(n_1038),
.Y(n_1177)
);

AO22x2_ASAP7_75t_L g1178 ( 
.A1(n_1104),
.A2(n_1060),
.B1(n_1063),
.B2(n_1047),
.Y(n_1178)
);

A2O1A1Ixp33_ASAP7_75t_L g1179 ( 
.A1(n_1019),
.A2(n_1088),
.B(n_999),
.C(n_1023),
.Y(n_1179)
);

NAND2x1_ASAP7_75t_L g1180 ( 
.A(n_1099),
.B(n_1013),
.Y(n_1180)
);

AOI21xp5_ASAP7_75t_L g1181 ( 
.A1(n_1099),
.A2(n_988),
.B(n_1045),
.Y(n_1181)
);

A2O1A1Ixp33_ASAP7_75t_L g1182 ( 
.A1(n_1074),
.A2(n_989),
.B(n_987),
.C(n_1128),
.Y(n_1182)
);

AO21x1_ASAP7_75t_L g1183 ( 
.A1(n_1031),
.A2(n_1076),
.B(n_988),
.Y(n_1183)
);

AOI21xp5_ASAP7_75t_L g1184 ( 
.A1(n_1121),
.A2(n_1026),
.B(n_1096),
.Y(n_1184)
);

AO31x2_ASAP7_75t_L g1185 ( 
.A1(n_1097),
.A2(n_991),
.A3(n_1068),
.B(n_1073),
.Y(n_1185)
);

INVxp67_ASAP7_75t_SL g1186 ( 
.A(n_1076),
.Y(n_1186)
);

AO21x1_ASAP7_75t_L g1187 ( 
.A1(n_991),
.A2(n_1032),
.B(n_1068),
.Y(n_1187)
);

BUFx12f_ASAP7_75t_L g1188 ( 
.A(n_1036),
.Y(n_1188)
);

NOR4xp25_ASAP7_75t_L g1189 ( 
.A(n_1053),
.B(n_1030),
.C(n_1042),
.D(n_1095),
.Y(n_1189)
);

NAND2xp5_ASAP7_75t_L g1190 ( 
.A(n_1000),
.B(n_1082),
.Y(n_1190)
);

NAND2xp5_ASAP7_75t_SL g1191 ( 
.A(n_1085),
.B(n_1000),
.Y(n_1191)
);

NAND2xp5_ASAP7_75t_L g1192 ( 
.A(n_1082),
.B(n_1040),
.Y(n_1192)
);

AOI21xp5_ASAP7_75t_SL g1193 ( 
.A1(n_1022),
.A2(n_1032),
.B(n_1073),
.Y(n_1193)
);

INVx1_ASAP7_75t_L g1194 ( 
.A(n_1132),
.Y(n_1194)
);

AO31x2_ASAP7_75t_L g1195 ( 
.A1(n_1097),
.A2(n_1022),
.A3(n_1059),
.B(n_1121),
.Y(n_1195)
);

OR2x6_ASAP7_75t_L g1196 ( 
.A(n_1051),
.B(n_1013),
.Y(n_1196)
);

OAI21x1_ASAP7_75t_L g1197 ( 
.A1(n_1096),
.A2(n_1132),
.B(n_1059),
.Y(n_1197)
);

INVx1_ASAP7_75t_L g1198 ( 
.A(n_1082),
.Y(n_1198)
);

OAI21x1_ASAP7_75t_L g1199 ( 
.A1(n_1036),
.A2(n_1010),
.B(n_1119),
.Y(n_1199)
);

OAI21xp5_ASAP7_75t_L g1200 ( 
.A1(n_1008),
.A2(n_1089),
.B(n_1086),
.Y(n_1200)
);

NOR2x1_ASAP7_75t_R g1201 ( 
.A(n_1069),
.B(n_489),
.Y(n_1201)
);

OA21x2_ASAP7_75t_L g1202 ( 
.A1(n_1064),
.A2(n_1131),
.B(n_1127),
.Y(n_1202)
);

AO21x2_ASAP7_75t_L g1203 ( 
.A1(n_1127),
.A2(n_1131),
.B(n_1064),
.Y(n_1203)
);

NAND2xp5_ASAP7_75t_L g1204 ( 
.A(n_1061),
.B(n_692),
.Y(n_1204)
);

HB1xp67_ASAP7_75t_L g1205 ( 
.A(n_1011),
.Y(n_1205)
);

NAND2xp5_ASAP7_75t_L g1206 ( 
.A(n_1061),
.B(n_692),
.Y(n_1206)
);

OAI21x1_ASAP7_75t_L g1207 ( 
.A1(n_1010),
.A2(n_1119),
.B(n_930),
.Y(n_1207)
);

OAI22xp5_ASAP7_75t_L g1208 ( 
.A1(n_1061),
.A2(n_692),
.B1(n_994),
.B2(n_798),
.Y(n_1208)
);

OAI21xp5_ASAP7_75t_L g1209 ( 
.A1(n_1008),
.A2(n_1089),
.B(n_1086),
.Y(n_1209)
);

BUFx6f_ASAP7_75t_L g1210 ( 
.A(n_1051),
.Y(n_1210)
);

INVx1_ASAP7_75t_L g1211 ( 
.A(n_1012),
.Y(n_1211)
);

AOI21xp5_ASAP7_75t_L g1212 ( 
.A1(n_1130),
.A2(n_691),
.B(n_993),
.Y(n_1212)
);

AOI21xp5_ASAP7_75t_L g1213 ( 
.A1(n_1130),
.A2(n_691),
.B(n_993),
.Y(n_1213)
);

OAI22xp5_ASAP7_75t_L g1214 ( 
.A1(n_1061),
.A2(n_692),
.B1(n_994),
.B2(n_798),
.Y(n_1214)
);

AO21x1_ASAP7_75t_L g1215 ( 
.A1(n_1055),
.A2(n_1056),
.B(n_998),
.Y(n_1215)
);

OAI21x1_ASAP7_75t_L g1216 ( 
.A1(n_1010),
.A2(n_1119),
.B(n_930),
.Y(n_1216)
);

OA21x2_ASAP7_75t_L g1217 ( 
.A1(n_1064),
.A2(n_1131),
.B(n_1127),
.Y(n_1217)
);

AOI21xp5_ASAP7_75t_L g1218 ( 
.A1(n_1130),
.A2(n_691),
.B(n_993),
.Y(n_1218)
);

AND2x2_ASAP7_75t_L g1219 ( 
.A(n_992),
.B(n_693),
.Y(n_1219)
);

AOI21xp5_ASAP7_75t_L g1220 ( 
.A1(n_1130),
.A2(n_691),
.B(n_993),
.Y(n_1220)
);

AND2x4_ASAP7_75t_L g1221 ( 
.A(n_985),
.B(n_1128),
.Y(n_1221)
);

AOI21xp5_ASAP7_75t_L g1222 ( 
.A1(n_1130),
.A2(n_691),
.B(n_993),
.Y(n_1222)
);

OAI21x1_ASAP7_75t_L g1223 ( 
.A1(n_1010),
.A2(n_1119),
.B(n_930),
.Y(n_1223)
);

HB1xp67_ASAP7_75t_L g1224 ( 
.A(n_1011),
.Y(n_1224)
);

AO31x2_ASAP7_75t_L g1225 ( 
.A1(n_1008),
.A2(n_866),
.A3(n_833),
.B(n_807),
.Y(n_1225)
);

O2A1O1Ixp33_ASAP7_75t_L g1226 ( 
.A1(n_1005),
.A2(n_799),
.B(n_798),
.C(n_912),
.Y(n_1226)
);

NAND2xp5_ASAP7_75t_SL g1227 ( 
.A(n_1005),
.B(n_902),
.Y(n_1227)
);

BUFx2_ASAP7_75t_L g1228 ( 
.A(n_1002),
.Y(n_1228)
);

OAI21x1_ASAP7_75t_L g1229 ( 
.A1(n_1010),
.A2(n_1119),
.B(n_930),
.Y(n_1229)
);

OAI22xp5_ASAP7_75t_L g1230 ( 
.A1(n_994),
.A2(n_995),
.B1(n_798),
.B2(n_1061),
.Y(n_1230)
);

INVx1_ASAP7_75t_L g1231 ( 
.A(n_1012),
.Y(n_1231)
);

AO21x1_ASAP7_75t_L g1232 ( 
.A1(n_1055),
.A2(n_1056),
.B(n_998),
.Y(n_1232)
);

OAI22xp5_ASAP7_75t_L g1233 ( 
.A1(n_1061),
.A2(n_692),
.B1(n_994),
.B2(n_798),
.Y(n_1233)
);

AOI21xp5_ASAP7_75t_SL g1234 ( 
.A1(n_1008),
.A2(n_995),
.B(n_734),
.Y(n_1234)
);

AOI21xp5_ASAP7_75t_L g1235 ( 
.A1(n_1130),
.A2(n_691),
.B(n_993),
.Y(n_1235)
);

INVx2_ASAP7_75t_SL g1236 ( 
.A(n_1069),
.Y(n_1236)
);

BUFx8_ASAP7_75t_SL g1237 ( 
.A(n_990),
.Y(n_1237)
);

OR2x2_ASAP7_75t_L g1238 ( 
.A(n_1005),
.B(n_848),
.Y(n_1238)
);

OAI21xp5_ASAP7_75t_L g1239 ( 
.A1(n_1008),
.A2(n_1089),
.B(n_1086),
.Y(n_1239)
);

AO31x2_ASAP7_75t_L g1240 ( 
.A1(n_1008),
.A2(n_866),
.A3(n_833),
.B(n_807),
.Y(n_1240)
);

BUFx3_ASAP7_75t_L g1241 ( 
.A(n_990),
.Y(n_1241)
);

AND2x2_ASAP7_75t_L g1242 ( 
.A(n_992),
.B(n_693),
.Y(n_1242)
);

BUFx2_ASAP7_75t_L g1243 ( 
.A(n_1002),
.Y(n_1243)
);

INVx3_ASAP7_75t_L g1244 ( 
.A(n_1099),
.Y(n_1244)
);

AO21x2_ASAP7_75t_L g1245 ( 
.A1(n_1127),
.A2(n_1131),
.B(n_1064),
.Y(n_1245)
);

A2O1A1Ixp33_ASAP7_75t_L g1246 ( 
.A1(n_1007),
.A2(n_692),
.B(n_798),
.C(n_799),
.Y(n_1246)
);

AO31x2_ASAP7_75t_L g1247 ( 
.A1(n_1008),
.A2(n_866),
.A3(n_833),
.B(n_807),
.Y(n_1247)
);

OAI21x1_ASAP7_75t_L g1248 ( 
.A1(n_1010),
.A2(n_1119),
.B(n_930),
.Y(n_1248)
);

AOI21xp5_ASAP7_75t_L g1249 ( 
.A1(n_1130),
.A2(n_691),
.B(n_993),
.Y(n_1249)
);

INVxp67_ASAP7_75t_L g1250 ( 
.A(n_1038),
.Y(n_1250)
);

OAI21x1_ASAP7_75t_L g1251 ( 
.A1(n_1010),
.A2(n_1119),
.B(n_930),
.Y(n_1251)
);

OAI22xp5_ASAP7_75t_L g1252 ( 
.A1(n_1061),
.A2(n_692),
.B1(n_994),
.B2(n_798),
.Y(n_1252)
);

CKINVDCx11_ASAP7_75t_R g1253 ( 
.A(n_990),
.Y(n_1253)
);

AOI21xp5_ASAP7_75t_L g1254 ( 
.A1(n_1130),
.A2(n_691),
.B(n_993),
.Y(n_1254)
);

INVx2_ASAP7_75t_L g1255 ( 
.A(n_1012),
.Y(n_1255)
);

AOI21xp5_ASAP7_75t_L g1256 ( 
.A1(n_1130),
.A2(n_691),
.B(n_993),
.Y(n_1256)
);

NAND2xp5_ASAP7_75t_L g1257 ( 
.A(n_1061),
.B(n_692),
.Y(n_1257)
);

NAND2xp5_ASAP7_75t_SL g1258 ( 
.A(n_1005),
.B(n_902),
.Y(n_1258)
);

OAI22x1_ASAP7_75t_L g1259 ( 
.A1(n_1005),
.A2(n_798),
.B1(n_576),
.B2(n_607),
.Y(n_1259)
);

OAI21xp5_ASAP7_75t_L g1260 ( 
.A1(n_1008),
.A2(n_1089),
.B(n_1086),
.Y(n_1260)
);

OAI21x1_ASAP7_75t_L g1261 ( 
.A1(n_1010),
.A2(n_1119),
.B(n_930),
.Y(n_1261)
);

INVx2_ASAP7_75t_SL g1262 ( 
.A(n_1069),
.Y(n_1262)
);

OAI22x1_ASAP7_75t_L g1263 ( 
.A1(n_1005),
.A2(n_798),
.B1(n_576),
.B2(n_607),
.Y(n_1263)
);

INVx1_ASAP7_75t_L g1264 ( 
.A(n_1012),
.Y(n_1264)
);

OR2x2_ASAP7_75t_L g1265 ( 
.A(n_1005),
.B(n_848),
.Y(n_1265)
);

A2O1A1Ixp33_ASAP7_75t_L g1266 ( 
.A1(n_1007),
.A2(n_692),
.B(n_798),
.C(n_799),
.Y(n_1266)
);

INVx1_ASAP7_75t_L g1267 ( 
.A(n_1012),
.Y(n_1267)
);

BUFx2_ASAP7_75t_R g1268 ( 
.A(n_1065),
.Y(n_1268)
);

OAI21xp5_ASAP7_75t_L g1269 ( 
.A1(n_1008),
.A2(n_1089),
.B(n_1086),
.Y(n_1269)
);

NAND3xp33_ASAP7_75t_L g1270 ( 
.A(n_1007),
.B(n_692),
.C(n_798),
.Y(n_1270)
);

INVx1_ASAP7_75t_L g1271 ( 
.A(n_1255),
.Y(n_1271)
);

AOI22xp33_ASAP7_75t_SL g1272 ( 
.A1(n_1270),
.A2(n_1233),
.B1(n_1252),
.B2(n_1208),
.Y(n_1272)
);

INVx3_ASAP7_75t_L g1273 ( 
.A(n_1180),
.Y(n_1273)
);

INVx2_ASAP7_75t_L g1274 ( 
.A(n_1163),
.Y(n_1274)
);

INVx2_ASAP7_75t_SL g1275 ( 
.A(n_1175),
.Y(n_1275)
);

INVx6_ASAP7_75t_L g1276 ( 
.A(n_1148),
.Y(n_1276)
);

BUFx10_ASAP7_75t_L g1277 ( 
.A(n_1176),
.Y(n_1277)
);

INVx6_ASAP7_75t_L g1278 ( 
.A(n_1148),
.Y(n_1278)
);

INVx2_ASAP7_75t_L g1279 ( 
.A(n_1152),
.Y(n_1279)
);

CKINVDCx14_ASAP7_75t_R g1280 ( 
.A(n_1153),
.Y(n_1280)
);

AOI22xp33_ASAP7_75t_L g1281 ( 
.A1(n_1215),
.A2(n_1232),
.B1(n_1214),
.B2(n_1230),
.Y(n_1281)
);

AOI22xp33_ASAP7_75t_L g1282 ( 
.A1(n_1230),
.A2(n_1150),
.B1(n_1263),
.B2(n_1259),
.Y(n_1282)
);

BUFx10_ASAP7_75t_L g1283 ( 
.A(n_1176),
.Y(n_1283)
);

INVx1_ASAP7_75t_SL g1284 ( 
.A(n_1238),
.Y(n_1284)
);

CKINVDCx5p33_ASAP7_75t_R g1285 ( 
.A(n_1237),
.Y(n_1285)
);

BUFx12f_ASAP7_75t_L g1286 ( 
.A(n_1253),
.Y(n_1286)
);

INVx1_ASAP7_75t_SL g1287 ( 
.A(n_1265),
.Y(n_1287)
);

INVx2_ASAP7_75t_L g1288 ( 
.A(n_1211),
.Y(n_1288)
);

OAI21xp33_ASAP7_75t_L g1289 ( 
.A1(n_1246),
.A2(n_1266),
.B(n_1162),
.Y(n_1289)
);

AOI22xp33_ASAP7_75t_SL g1290 ( 
.A1(n_1257),
.A2(n_1178),
.B1(n_1269),
.B2(n_1200),
.Y(n_1290)
);

AOI22xp33_ASAP7_75t_L g1291 ( 
.A1(n_1157),
.A2(n_1162),
.B1(n_1219),
.B2(n_1242),
.Y(n_1291)
);

CKINVDCx11_ASAP7_75t_R g1292 ( 
.A(n_1188),
.Y(n_1292)
);

INVx4_ASAP7_75t_L g1293 ( 
.A(n_1148),
.Y(n_1293)
);

BUFx2_ASAP7_75t_L g1294 ( 
.A(n_1205),
.Y(n_1294)
);

CKINVDCx20_ASAP7_75t_R g1295 ( 
.A(n_1241),
.Y(n_1295)
);

AOI22xp33_ASAP7_75t_L g1296 ( 
.A1(n_1146),
.A2(n_1178),
.B1(n_1151),
.B2(n_1239),
.Y(n_1296)
);

INVx1_ASAP7_75t_L g1297 ( 
.A(n_1231),
.Y(n_1297)
);

INVx6_ASAP7_75t_L g1298 ( 
.A(n_1196),
.Y(n_1298)
);

CKINVDCx11_ASAP7_75t_R g1299 ( 
.A(n_1144),
.Y(n_1299)
);

CKINVDCx8_ASAP7_75t_R g1300 ( 
.A(n_1228),
.Y(n_1300)
);

OAI22xp5_ASAP7_75t_L g1301 ( 
.A1(n_1136),
.A2(n_1141),
.B1(n_1182),
.B2(n_1227),
.Y(n_1301)
);

OAI21xp33_ASAP7_75t_SL g1302 ( 
.A1(n_1140),
.A2(n_1234),
.B(n_1174),
.Y(n_1302)
);

INVx2_ASAP7_75t_L g1303 ( 
.A(n_1264),
.Y(n_1303)
);

AOI22xp33_ASAP7_75t_L g1304 ( 
.A1(n_1200),
.A2(n_1269),
.B1(n_1209),
.B2(n_1239),
.Y(n_1304)
);

AOI22xp33_ASAP7_75t_L g1305 ( 
.A1(n_1209),
.A2(n_1260),
.B1(n_1169),
.B2(n_1245),
.Y(n_1305)
);

INVx2_ASAP7_75t_L g1306 ( 
.A(n_1267),
.Y(n_1306)
);

AOI22xp5_ASAP7_75t_L g1307 ( 
.A1(n_1258),
.A2(n_1143),
.B1(n_1221),
.B2(n_1191),
.Y(n_1307)
);

AOI22xp33_ASAP7_75t_L g1308 ( 
.A1(n_1260),
.A2(n_1203),
.B1(n_1245),
.B2(n_1171),
.Y(n_1308)
);

OAI21xp5_ASAP7_75t_SL g1309 ( 
.A1(n_1138),
.A2(n_1226),
.B(n_1134),
.Y(n_1309)
);

BUFx2_ASAP7_75t_L g1310 ( 
.A(n_1224),
.Y(n_1310)
);

INVx6_ASAP7_75t_L g1311 ( 
.A(n_1196),
.Y(n_1311)
);

AOI22xp33_ASAP7_75t_L g1312 ( 
.A1(n_1203),
.A2(n_1142),
.B1(n_1217),
.B2(n_1202),
.Y(n_1312)
);

AOI22xp5_ASAP7_75t_L g1313 ( 
.A1(n_1143),
.A2(n_1221),
.B1(n_1189),
.B2(n_1243),
.Y(n_1313)
);

CKINVDCx11_ASAP7_75t_R g1314 ( 
.A(n_1176),
.Y(n_1314)
);

INVx6_ASAP7_75t_L g1315 ( 
.A(n_1210),
.Y(n_1315)
);

BUFx10_ASAP7_75t_L g1316 ( 
.A(n_1210),
.Y(n_1316)
);

OAI22xp33_ASAP7_75t_L g1317 ( 
.A1(n_1142),
.A2(n_1173),
.B1(n_1189),
.B2(n_1160),
.Y(n_1317)
);

AOI22xp33_ASAP7_75t_L g1318 ( 
.A1(n_1202),
.A2(n_1217),
.B1(n_1156),
.B2(n_1159),
.Y(n_1318)
);

OAI22xp5_ASAP7_75t_L g1319 ( 
.A1(n_1164),
.A2(n_1179),
.B1(n_1250),
.B2(n_1177),
.Y(n_1319)
);

INVx5_ASAP7_75t_L g1320 ( 
.A(n_1244),
.Y(n_1320)
);

INVx2_ASAP7_75t_SL g1321 ( 
.A(n_1236),
.Y(n_1321)
);

INVx6_ASAP7_75t_L g1322 ( 
.A(n_1210),
.Y(n_1322)
);

INVx6_ASAP7_75t_L g1323 ( 
.A(n_1268),
.Y(n_1323)
);

BUFx3_ASAP7_75t_L g1324 ( 
.A(n_1262),
.Y(n_1324)
);

AOI22xp5_ASAP7_75t_L g1325 ( 
.A1(n_1172),
.A2(n_1190),
.B1(n_1192),
.B2(n_1158),
.Y(n_1325)
);

BUFx8_ASAP7_75t_L g1326 ( 
.A(n_1194),
.Y(n_1326)
);

AOI22xp33_ASAP7_75t_L g1327 ( 
.A1(n_1139),
.A2(n_1149),
.B1(n_1166),
.B2(n_1198),
.Y(n_1327)
);

INVx1_ASAP7_75t_L g1328 ( 
.A(n_1186),
.Y(n_1328)
);

INVx1_ASAP7_75t_L g1329 ( 
.A(n_1185),
.Y(n_1329)
);

CKINVDCx11_ASAP7_75t_R g1330 ( 
.A(n_1201),
.Y(n_1330)
);

CKINVDCx6p67_ASAP7_75t_R g1331 ( 
.A(n_1201),
.Y(n_1331)
);

BUFx2_ASAP7_75t_SL g1332 ( 
.A(n_1187),
.Y(n_1332)
);

AOI22xp33_ASAP7_75t_L g1333 ( 
.A1(n_1212),
.A2(n_1222),
.B1(n_1220),
.B2(n_1256),
.Y(n_1333)
);

OAI21xp5_ASAP7_75t_SL g1334 ( 
.A1(n_1154),
.A2(n_1235),
.B(n_1254),
.Y(n_1334)
);

BUFx12f_ASAP7_75t_L g1335 ( 
.A(n_1193),
.Y(n_1335)
);

INVx3_ASAP7_75t_L g1336 ( 
.A(n_1197),
.Y(n_1336)
);

BUFx10_ASAP7_75t_L g1337 ( 
.A(n_1167),
.Y(n_1337)
);

AOI22xp33_ASAP7_75t_SL g1338 ( 
.A1(n_1181),
.A2(n_1213),
.B1(n_1249),
.B2(n_1218),
.Y(n_1338)
);

AOI22xp33_ASAP7_75t_SL g1339 ( 
.A1(n_1165),
.A2(n_1145),
.B1(n_1147),
.B2(n_1184),
.Y(n_1339)
);

AOI22xp33_ASAP7_75t_SL g1340 ( 
.A1(n_1145),
.A2(n_1147),
.B1(n_1199),
.B2(n_1137),
.Y(n_1340)
);

INVx1_ASAP7_75t_L g1341 ( 
.A(n_1168),
.Y(n_1341)
);

INVx1_ASAP7_75t_SL g1342 ( 
.A(n_1135),
.Y(n_1342)
);

CKINVDCx20_ASAP7_75t_R g1343 ( 
.A(n_1183),
.Y(n_1343)
);

INVx1_ASAP7_75t_L g1344 ( 
.A(n_1168),
.Y(n_1344)
);

AOI22xp33_ASAP7_75t_L g1345 ( 
.A1(n_1207),
.A2(n_1223),
.B1(n_1251),
.B2(n_1248),
.Y(n_1345)
);

OAI22xp5_ASAP7_75t_L g1346 ( 
.A1(n_1170),
.A2(n_1145),
.B1(n_1147),
.B2(n_1155),
.Y(n_1346)
);

CKINVDCx20_ASAP7_75t_R g1347 ( 
.A(n_1195),
.Y(n_1347)
);

BUFx4f_ASAP7_75t_SL g1348 ( 
.A(n_1155),
.Y(n_1348)
);

BUFx6f_ASAP7_75t_L g1349 ( 
.A(n_1216),
.Y(n_1349)
);

INVx6_ASAP7_75t_L g1350 ( 
.A(n_1225),
.Y(n_1350)
);

INVx8_ASAP7_75t_L g1351 ( 
.A(n_1229),
.Y(n_1351)
);

CKINVDCx11_ASAP7_75t_R g1352 ( 
.A(n_1240),
.Y(n_1352)
);

BUFx12f_ASAP7_75t_L g1353 ( 
.A(n_1247),
.Y(n_1353)
);

OAI22xp5_ASAP7_75t_L g1354 ( 
.A1(n_1247),
.A2(n_798),
.B1(n_1270),
.B2(n_1206),
.Y(n_1354)
);

CKINVDCx12_ASAP7_75t_R g1355 ( 
.A(n_1247),
.Y(n_1355)
);

NOR2x1_ASAP7_75t_SL g1356 ( 
.A(n_1261),
.B(n_1148),
.Y(n_1356)
);

AOI22xp33_ASAP7_75t_L g1357 ( 
.A1(n_1270),
.A2(n_798),
.B1(n_1232),
.B2(n_1215),
.Y(n_1357)
);

AND2x2_ASAP7_75t_L g1358 ( 
.A(n_1219),
.B(n_1242),
.Y(n_1358)
);

BUFx6f_ASAP7_75t_L g1359 ( 
.A(n_1148),
.Y(n_1359)
);

INVx1_ASAP7_75t_L g1360 ( 
.A(n_1255),
.Y(n_1360)
);

BUFx2_ASAP7_75t_L g1361 ( 
.A(n_1161),
.Y(n_1361)
);

OAI22xp5_ASAP7_75t_L g1362 ( 
.A1(n_1270),
.A2(n_798),
.B1(n_1206),
.B2(n_1204),
.Y(n_1362)
);

CKINVDCx5p33_ASAP7_75t_R g1363 ( 
.A(n_1237),
.Y(n_1363)
);

BUFx12f_ASAP7_75t_L g1364 ( 
.A(n_1153),
.Y(n_1364)
);

AOI22xp33_ASAP7_75t_SL g1365 ( 
.A1(n_1270),
.A2(n_994),
.B1(n_798),
.B2(n_995),
.Y(n_1365)
);

AND2x2_ASAP7_75t_L g1366 ( 
.A(n_1219),
.B(n_1242),
.Y(n_1366)
);

BUFx4f_ASAP7_75t_SL g1367 ( 
.A(n_1188),
.Y(n_1367)
);

AOI22xp33_ASAP7_75t_SL g1368 ( 
.A1(n_1270),
.A2(n_994),
.B1(n_798),
.B2(n_995),
.Y(n_1368)
);

INVx6_ASAP7_75t_L g1369 ( 
.A(n_1148),
.Y(n_1369)
);

AOI22xp33_ASAP7_75t_L g1370 ( 
.A1(n_1270),
.A2(n_798),
.B1(n_1232),
.B2(n_1215),
.Y(n_1370)
);

BUFx2_ASAP7_75t_L g1371 ( 
.A(n_1161),
.Y(n_1371)
);

CKINVDCx20_ASAP7_75t_R g1372 ( 
.A(n_1237),
.Y(n_1372)
);

INVx1_ASAP7_75t_L g1373 ( 
.A(n_1255),
.Y(n_1373)
);

OAI22xp5_ASAP7_75t_L g1374 ( 
.A1(n_1270),
.A2(n_798),
.B1(n_1206),
.B2(n_1204),
.Y(n_1374)
);

CKINVDCx6p67_ASAP7_75t_R g1375 ( 
.A(n_1153),
.Y(n_1375)
);

INVx2_ASAP7_75t_R g1376 ( 
.A(n_1194),
.Y(n_1376)
);

NAND2x1p5_ASAP7_75t_L g1377 ( 
.A(n_1244),
.B(n_1094),
.Y(n_1377)
);

INVx4_ASAP7_75t_L g1378 ( 
.A(n_1148),
.Y(n_1378)
);

AND2x4_ASAP7_75t_L g1379 ( 
.A(n_1356),
.B(n_1336),
.Y(n_1379)
);

AND2x2_ASAP7_75t_L g1380 ( 
.A(n_1282),
.B(n_1304),
.Y(n_1380)
);

INVx2_ASAP7_75t_SL g1381 ( 
.A(n_1276),
.Y(n_1381)
);

AND2x2_ASAP7_75t_L g1382 ( 
.A(n_1282),
.B(n_1304),
.Y(n_1382)
);

BUFx6f_ASAP7_75t_L g1383 ( 
.A(n_1349),
.Y(n_1383)
);

AOI21xp5_ASAP7_75t_L g1384 ( 
.A1(n_1317),
.A2(n_1333),
.B(n_1302),
.Y(n_1384)
);

OA21x2_ASAP7_75t_L g1385 ( 
.A1(n_1334),
.A2(n_1344),
.B(n_1341),
.Y(n_1385)
);

BUFx2_ASAP7_75t_L g1386 ( 
.A(n_1353),
.Y(n_1386)
);

HB1xp67_ASAP7_75t_L g1387 ( 
.A(n_1294),
.Y(n_1387)
);

INVx1_ASAP7_75t_L g1388 ( 
.A(n_1329),
.Y(n_1388)
);

NOR2xp33_ASAP7_75t_L g1389 ( 
.A(n_1284),
.B(n_1287),
.Y(n_1389)
);

OAI21x1_ASAP7_75t_L g1390 ( 
.A1(n_1345),
.A2(n_1333),
.B(n_1327),
.Y(n_1390)
);

INVx3_ASAP7_75t_L g1391 ( 
.A(n_1351),
.Y(n_1391)
);

CKINVDCx20_ASAP7_75t_R g1392 ( 
.A(n_1372),
.Y(n_1392)
);

INVx1_ASAP7_75t_L g1393 ( 
.A(n_1355),
.Y(n_1393)
);

OR2x6_ASAP7_75t_L g1394 ( 
.A(n_1351),
.B(n_1350),
.Y(n_1394)
);

OR2x2_ASAP7_75t_L g1395 ( 
.A(n_1308),
.B(n_1312),
.Y(n_1395)
);

AO21x2_ASAP7_75t_L g1396 ( 
.A1(n_1317),
.A2(n_1346),
.B(n_1309),
.Y(n_1396)
);

OAI21x1_ASAP7_75t_L g1397 ( 
.A1(n_1345),
.A2(n_1327),
.B(n_1318),
.Y(n_1397)
);

INVx1_ASAP7_75t_L g1398 ( 
.A(n_1348),
.Y(n_1398)
);

BUFx12f_ASAP7_75t_L g1399 ( 
.A(n_1292),
.Y(n_1399)
);

OAI21x1_ASAP7_75t_L g1400 ( 
.A1(n_1318),
.A2(n_1312),
.B(n_1308),
.Y(n_1400)
);

AND2x2_ASAP7_75t_L g1401 ( 
.A(n_1290),
.B(n_1272),
.Y(n_1401)
);

AND2x2_ASAP7_75t_L g1402 ( 
.A(n_1290),
.B(n_1272),
.Y(n_1402)
);

INVx2_ASAP7_75t_L g1403 ( 
.A(n_1342),
.Y(n_1403)
);

AOI22xp33_ASAP7_75t_L g1404 ( 
.A1(n_1365),
.A2(n_1368),
.B1(n_1289),
.B2(n_1301),
.Y(n_1404)
);

OAI21x1_ASAP7_75t_L g1405 ( 
.A1(n_1354),
.A2(n_1370),
.B(n_1357),
.Y(n_1405)
);

AND2x2_ASAP7_75t_L g1406 ( 
.A(n_1305),
.B(n_1281),
.Y(n_1406)
);

AND2x2_ASAP7_75t_L g1407 ( 
.A(n_1305),
.B(n_1281),
.Y(n_1407)
);

BUFx2_ASAP7_75t_SL g1408 ( 
.A(n_1320),
.Y(n_1408)
);

INVx1_ASAP7_75t_L g1409 ( 
.A(n_1297),
.Y(n_1409)
);

BUFx2_ASAP7_75t_R g1410 ( 
.A(n_1285),
.Y(n_1410)
);

NAND2xp5_ASAP7_75t_L g1411 ( 
.A(n_1362),
.B(n_1374),
.Y(n_1411)
);

CKINVDCx20_ASAP7_75t_R g1412 ( 
.A(n_1372),
.Y(n_1412)
);

AND2x2_ASAP7_75t_L g1413 ( 
.A(n_1365),
.B(n_1368),
.Y(n_1413)
);

OAI21x1_ASAP7_75t_L g1414 ( 
.A1(n_1357),
.A2(n_1370),
.B(n_1296),
.Y(n_1414)
);

INVx1_ASAP7_75t_L g1415 ( 
.A(n_1347),
.Y(n_1415)
);

INVx1_ASAP7_75t_L g1416 ( 
.A(n_1347),
.Y(n_1416)
);

INVx2_ASAP7_75t_L g1417 ( 
.A(n_1352),
.Y(n_1417)
);

AO21x2_ASAP7_75t_L g1418 ( 
.A1(n_1325),
.A2(n_1319),
.B(n_1338),
.Y(n_1418)
);

INVx1_ASAP7_75t_L g1419 ( 
.A(n_1279),
.Y(n_1419)
);

INVxp33_ASAP7_75t_L g1420 ( 
.A(n_1358),
.Y(n_1420)
);

HB1xp67_ASAP7_75t_L g1421 ( 
.A(n_1310),
.Y(n_1421)
);

OR2x6_ASAP7_75t_L g1422 ( 
.A(n_1332),
.B(n_1335),
.Y(n_1422)
);

INVx2_ASAP7_75t_SL g1423 ( 
.A(n_1276),
.Y(n_1423)
);

NAND2xp5_ASAP7_75t_L g1424 ( 
.A(n_1296),
.B(n_1291),
.Y(n_1424)
);

OR2x2_ASAP7_75t_L g1425 ( 
.A(n_1291),
.B(n_1366),
.Y(n_1425)
);

INVx1_ASAP7_75t_L g1426 ( 
.A(n_1288),
.Y(n_1426)
);

INVx2_ASAP7_75t_SL g1427 ( 
.A(n_1278),
.Y(n_1427)
);

BUFx12f_ASAP7_75t_L g1428 ( 
.A(n_1292),
.Y(n_1428)
);

CKINVDCx16_ASAP7_75t_R g1429 ( 
.A(n_1286),
.Y(n_1429)
);

AO21x1_ASAP7_75t_SL g1430 ( 
.A1(n_1313),
.A2(n_1328),
.B(n_1271),
.Y(n_1430)
);

OA21x2_ASAP7_75t_L g1431 ( 
.A1(n_1303),
.A2(n_1306),
.B(n_1360),
.Y(n_1431)
);

INVx2_ASAP7_75t_L g1432 ( 
.A(n_1373),
.Y(n_1432)
);

INVx1_ASAP7_75t_L g1433 ( 
.A(n_1376),
.Y(n_1433)
);

INVx1_ASAP7_75t_L g1434 ( 
.A(n_1339),
.Y(n_1434)
);

INVx1_ASAP7_75t_L g1435 ( 
.A(n_1339),
.Y(n_1435)
);

INVx3_ASAP7_75t_L g1436 ( 
.A(n_1337),
.Y(n_1436)
);

INVx1_ASAP7_75t_L g1437 ( 
.A(n_1340),
.Y(n_1437)
);

INVx1_ASAP7_75t_L g1438 ( 
.A(n_1340),
.Y(n_1438)
);

HB1xp67_ASAP7_75t_L g1439 ( 
.A(n_1361),
.Y(n_1439)
);

INVxp33_ASAP7_75t_L g1440 ( 
.A(n_1299),
.Y(n_1440)
);

INVx4_ASAP7_75t_L g1441 ( 
.A(n_1320),
.Y(n_1441)
);

INVxp67_ASAP7_75t_L g1442 ( 
.A(n_1371),
.Y(n_1442)
);

INVx2_ASAP7_75t_L g1443 ( 
.A(n_1337),
.Y(n_1443)
);

INVx1_ASAP7_75t_L g1444 ( 
.A(n_1343),
.Y(n_1444)
);

AO21x2_ASAP7_75t_L g1445 ( 
.A1(n_1338),
.A2(n_1274),
.B(n_1343),
.Y(n_1445)
);

AO32x2_ASAP7_75t_L g1446 ( 
.A1(n_1381),
.A2(n_1275),
.A3(n_1378),
.B1(n_1293),
.B2(n_1321),
.Y(n_1446)
);

AND2x2_ASAP7_75t_L g1447 ( 
.A(n_1415),
.B(n_1307),
.Y(n_1447)
);

OA21x2_ASAP7_75t_L g1448 ( 
.A1(n_1384),
.A2(n_1320),
.B(n_1377),
.Y(n_1448)
);

INVxp67_ASAP7_75t_L g1449 ( 
.A(n_1389),
.Y(n_1449)
);

AND2x2_ASAP7_75t_L g1450 ( 
.A(n_1416),
.B(n_1359),
.Y(n_1450)
);

OR2x2_ASAP7_75t_L g1451 ( 
.A(n_1416),
.B(n_1375),
.Y(n_1451)
);

INVx2_ASAP7_75t_L g1452 ( 
.A(n_1431),
.Y(n_1452)
);

OR2x6_ASAP7_75t_L g1453 ( 
.A(n_1394),
.B(n_1298),
.Y(n_1453)
);

AO21x2_ASAP7_75t_L g1454 ( 
.A1(n_1397),
.A2(n_1369),
.B(n_1278),
.Y(n_1454)
);

OAI22xp5_ASAP7_75t_L g1455 ( 
.A1(n_1404),
.A2(n_1300),
.B1(n_1323),
.B2(n_1311),
.Y(n_1455)
);

INVxp67_ASAP7_75t_L g1456 ( 
.A(n_1387),
.Y(n_1456)
);

OR2x2_ASAP7_75t_L g1457 ( 
.A(n_1425),
.B(n_1359),
.Y(n_1457)
);

OAI21xp5_ASAP7_75t_L g1458 ( 
.A1(n_1411),
.A2(n_1377),
.B(n_1273),
.Y(n_1458)
);

INVx3_ASAP7_75t_L g1459 ( 
.A(n_1383),
.Y(n_1459)
);

NOR2xp33_ASAP7_75t_L g1460 ( 
.A(n_1401),
.B(n_1369),
.Y(n_1460)
);

HB1xp67_ASAP7_75t_L g1461 ( 
.A(n_1385),
.Y(n_1461)
);

OA21x2_ASAP7_75t_L g1462 ( 
.A1(n_1397),
.A2(n_1311),
.B(n_1273),
.Y(n_1462)
);

AOI22xp5_ASAP7_75t_L g1463 ( 
.A1(n_1401),
.A2(n_1295),
.B1(n_1331),
.B2(n_1280),
.Y(n_1463)
);

A2O1A1Ixp33_ASAP7_75t_L g1464 ( 
.A1(n_1402),
.A2(n_1280),
.B(n_1324),
.C(n_1326),
.Y(n_1464)
);

A2O1A1Ixp33_ASAP7_75t_L g1465 ( 
.A1(n_1402),
.A2(n_1295),
.B(n_1363),
.C(n_1330),
.Y(n_1465)
);

AND2x2_ASAP7_75t_L g1466 ( 
.A(n_1417),
.B(n_1323),
.Y(n_1466)
);

AND2x2_ASAP7_75t_L g1467 ( 
.A(n_1417),
.B(n_1420),
.Y(n_1467)
);

A2O1A1Ixp33_ASAP7_75t_L g1468 ( 
.A1(n_1414),
.A2(n_1330),
.B(n_1323),
.C(n_1314),
.Y(n_1468)
);

NOR2xp33_ASAP7_75t_L g1469 ( 
.A(n_1380),
.B(n_1299),
.Y(n_1469)
);

OAI22xp5_ASAP7_75t_L g1470 ( 
.A1(n_1444),
.A2(n_1413),
.B1(n_1424),
.B2(n_1417),
.Y(n_1470)
);

AND2x4_ASAP7_75t_L g1471 ( 
.A(n_1393),
.B(n_1314),
.Y(n_1471)
);

NAND2xp5_ASAP7_75t_L g1472 ( 
.A(n_1421),
.B(n_1315),
.Y(n_1472)
);

AND2x2_ASAP7_75t_L g1473 ( 
.A(n_1444),
.B(n_1315),
.Y(n_1473)
);

AO21x1_ASAP7_75t_L g1474 ( 
.A1(n_1424),
.A2(n_1322),
.B(n_1283),
.Y(n_1474)
);

OAI21xp5_ASAP7_75t_L g1475 ( 
.A1(n_1405),
.A2(n_1364),
.B(n_1283),
.Y(n_1475)
);

AOI21xp5_ASAP7_75t_L g1476 ( 
.A1(n_1418),
.A2(n_1277),
.B(n_1316),
.Y(n_1476)
);

OAI21xp5_ASAP7_75t_L g1477 ( 
.A1(n_1405),
.A2(n_1277),
.B(n_1316),
.Y(n_1477)
);

NOR2xp33_ASAP7_75t_L g1478 ( 
.A(n_1380),
.B(n_1322),
.Y(n_1478)
);

NAND2xp5_ASAP7_75t_L g1479 ( 
.A(n_1439),
.B(n_1367),
.Y(n_1479)
);

AND2x2_ASAP7_75t_L g1480 ( 
.A(n_1386),
.B(n_1430),
.Y(n_1480)
);

HB1xp67_ASAP7_75t_L g1481 ( 
.A(n_1385),
.Y(n_1481)
);

INVxp67_ASAP7_75t_SL g1482 ( 
.A(n_1403),
.Y(n_1482)
);

AO21x2_ASAP7_75t_L g1483 ( 
.A1(n_1390),
.A2(n_1418),
.B(n_1400),
.Y(n_1483)
);

AOI21xp5_ASAP7_75t_L g1484 ( 
.A1(n_1418),
.A2(n_1367),
.B(n_1396),
.Y(n_1484)
);

INVx2_ASAP7_75t_L g1485 ( 
.A(n_1409),
.Y(n_1485)
);

NOR2x1_ASAP7_75t_SL g1486 ( 
.A(n_1418),
.B(n_1422),
.Y(n_1486)
);

OR2x6_ASAP7_75t_L g1487 ( 
.A(n_1394),
.B(n_1408),
.Y(n_1487)
);

AND2x2_ASAP7_75t_L g1488 ( 
.A(n_1386),
.B(n_1413),
.Y(n_1488)
);

AND2x2_ASAP7_75t_L g1489 ( 
.A(n_1419),
.B(n_1426),
.Y(n_1489)
);

AND2x4_ASAP7_75t_L g1490 ( 
.A(n_1394),
.B(n_1391),
.Y(n_1490)
);

CKINVDCx20_ASAP7_75t_R g1491 ( 
.A(n_1392),
.Y(n_1491)
);

O2A1O1Ixp33_ASAP7_75t_L g1492 ( 
.A1(n_1382),
.A2(n_1407),
.B(n_1406),
.C(n_1442),
.Y(n_1492)
);

AO32x2_ASAP7_75t_L g1493 ( 
.A1(n_1423),
.A2(n_1427),
.A3(n_1441),
.B1(n_1396),
.B2(n_1445),
.Y(n_1493)
);

HB1xp67_ASAP7_75t_L g1494 ( 
.A(n_1385),
.Y(n_1494)
);

NOR2x1_ASAP7_75t_SL g1495 ( 
.A(n_1422),
.B(n_1445),
.Y(n_1495)
);

A2O1A1Ixp33_ASAP7_75t_L g1496 ( 
.A1(n_1414),
.A2(n_1407),
.B(n_1406),
.C(n_1382),
.Y(n_1496)
);

INVx1_ASAP7_75t_SL g1497 ( 
.A(n_1410),
.Y(n_1497)
);

CKINVDCx11_ASAP7_75t_R g1498 ( 
.A(n_1399),
.Y(n_1498)
);

OAI21x1_ASAP7_75t_L g1499 ( 
.A1(n_1390),
.A2(n_1400),
.B(n_1391),
.Y(n_1499)
);

INVx4_ASAP7_75t_L g1500 ( 
.A(n_1422),
.Y(n_1500)
);

OAI22xp5_ASAP7_75t_L g1501 ( 
.A1(n_1465),
.A2(n_1422),
.B1(n_1443),
.B2(n_1436),
.Y(n_1501)
);

AND2x2_ASAP7_75t_L g1502 ( 
.A(n_1493),
.B(n_1488),
.Y(n_1502)
);

AND2x2_ASAP7_75t_L g1503 ( 
.A(n_1493),
.B(n_1437),
.Y(n_1503)
);

INVx1_ASAP7_75t_L g1504 ( 
.A(n_1485),
.Y(n_1504)
);

AND2x4_ASAP7_75t_L g1505 ( 
.A(n_1487),
.B(n_1490),
.Y(n_1505)
);

OR2x2_ASAP7_75t_L g1506 ( 
.A(n_1482),
.B(n_1437),
.Y(n_1506)
);

AND2x2_ASAP7_75t_L g1507 ( 
.A(n_1493),
.B(n_1438),
.Y(n_1507)
);

AND2x4_ASAP7_75t_L g1508 ( 
.A(n_1487),
.B(n_1379),
.Y(n_1508)
);

NAND3xp33_ASAP7_75t_L g1509 ( 
.A(n_1484),
.B(n_1443),
.C(n_1438),
.Y(n_1509)
);

AND2x2_ASAP7_75t_L g1510 ( 
.A(n_1493),
.B(n_1445),
.Y(n_1510)
);

AND2x2_ASAP7_75t_L g1511 ( 
.A(n_1495),
.B(n_1445),
.Y(n_1511)
);

OR2x2_ASAP7_75t_L g1512 ( 
.A(n_1483),
.B(n_1396),
.Y(n_1512)
);

INVx2_ASAP7_75t_L g1513 ( 
.A(n_1452),
.Y(n_1513)
);

HB1xp67_ASAP7_75t_L g1514 ( 
.A(n_1456),
.Y(n_1514)
);

AND2x2_ASAP7_75t_L g1515 ( 
.A(n_1467),
.B(n_1434),
.Y(n_1515)
);

OAI22xp5_ASAP7_75t_L g1516 ( 
.A1(n_1465),
.A2(n_1422),
.B1(n_1443),
.B2(n_1436),
.Y(n_1516)
);

OR2x2_ASAP7_75t_L g1517 ( 
.A(n_1483),
.B(n_1396),
.Y(n_1517)
);

INVx1_ASAP7_75t_L g1518 ( 
.A(n_1452),
.Y(n_1518)
);

INVx3_ASAP7_75t_L g1519 ( 
.A(n_1459),
.Y(n_1519)
);

AND2x4_ASAP7_75t_L g1520 ( 
.A(n_1487),
.B(n_1379),
.Y(n_1520)
);

OR2x2_ASAP7_75t_L g1521 ( 
.A(n_1496),
.B(n_1395),
.Y(n_1521)
);

OR2x2_ASAP7_75t_L g1522 ( 
.A(n_1496),
.B(n_1395),
.Y(n_1522)
);

OR2x2_ASAP7_75t_L g1523 ( 
.A(n_1461),
.B(n_1385),
.Y(n_1523)
);

AND2x2_ASAP7_75t_L g1524 ( 
.A(n_1450),
.B(n_1434),
.Y(n_1524)
);

AND2x2_ASAP7_75t_L g1525 ( 
.A(n_1457),
.B(n_1435),
.Y(n_1525)
);

AND2x2_ASAP7_75t_L g1526 ( 
.A(n_1486),
.B(n_1435),
.Y(n_1526)
);

INVx1_ASAP7_75t_L g1527 ( 
.A(n_1489),
.Y(n_1527)
);

NAND2xp5_ASAP7_75t_L g1528 ( 
.A(n_1470),
.B(n_1432),
.Y(n_1528)
);

AND2x2_ASAP7_75t_L g1529 ( 
.A(n_1490),
.B(n_1433),
.Y(n_1529)
);

AND2x2_ASAP7_75t_L g1530 ( 
.A(n_1490),
.B(n_1433),
.Y(n_1530)
);

INVx1_ASAP7_75t_L g1531 ( 
.A(n_1446),
.Y(n_1531)
);

INVx3_ASAP7_75t_L g1532 ( 
.A(n_1513),
.Y(n_1532)
);

INVx1_ASAP7_75t_L g1533 ( 
.A(n_1504),
.Y(n_1533)
);

NAND2xp5_ASAP7_75t_L g1534 ( 
.A(n_1503),
.B(n_1461),
.Y(n_1534)
);

OAI221xp5_ASAP7_75t_L g1535 ( 
.A1(n_1521),
.A2(n_1468),
.B1(n_1464),
.B2(n_1463),
.C(n_1492),
.Y(n_1535)
);

INVx1_ASAP7_75t_L g1536 ( 
.A(n_1504),
.Y(n_1536)
);

HB1xp67_ASAP7_75t_L g1537 ( 
.A(n_1506),
.Y(n_1537)
);

NAND3xp33_ASAP7_75t_L g1538 ( 
.A(n_1509),
.B(n_1522),
.C(n_1521),
.Y(n_1538)
);

OAI221xp5_ASAP7_75t_L g1539 ( 
.A1(n_1522),
.A2(n_1468),
.B1(n_1464),
.B2(n_1475),
.C(n_1455),
.Y(n_1539)
);

HB1xp67_ASAP7_75t_L g1540 ( 
.A(n_1506),
.Y(n_1540)
);

NAND2xp5_ASAP7_75t_L g1541 ( 
.A(n_1503),
.B(n_1481),
.Y(n_1541)
);

AND2x4_ASAP7_75t_L g1542 ( 
.A(n_1508),
.B(n_1500),
.Y(n_1542)
);

HB1xp67_ASAP7_75t_L g1543 ( 
.A(n_1514),
.Y(n_1543)
);

NAND2xp5_ASAP7_75t_L g1544 ( 
.A(n_1507),
.B(n_1481),
.Y(n_1544)
);

OAI22xp5_ASAP7_75t_L g1545 ( 
.A1(n_1510),
.A2(n_1469),
.B1(n_1460),
.B2(n_1449),
.Y(n_1545)
);

HB1xp67_ASAP7_75t_L g1546 ( 
.A(n_1518),
.Y(n_1546)
);

OR2x2_ASAP7_75t_L g1547 ( 
.A(n_1502),
.B(n_1494),
.Y(n_1547)
);

AND2x2_ASAP7_75t_L g1548 ( 
.A(n_1502),
.B(n_1462),
.Y(n_1548)
);

INVxp67_ASAP7_75t_SL g1549 ( 
.A(n_1523),
.Y(n_1549)
);

NAND3xp33_ASAP7_75t_L g1550 ( 
.A(n_1512),
.B(n_1469),
.C(n_1477),
.Y(n_1550)
);

AOI221xp5_ASAP7_75t_L g1551 ( 
.A1(n_1510),
.A2(n_1460),
.B1(n_1478),
.B2(n_1447),
.C(n_1494),
.Y(n_1551)
);

NAND2xp5_ASAP7_75t_L g1552 ( 
.A(n_1507),
.B(n_1388),
.Y(n_1552)
);

AND2x2_ASAP7_75t_L g1553 ( 
.A(n_1529),
.B(n_1462),
.Y(n_1553)
);

INVx2_ASAP7_75t_L g1554 ( 
.A(n_1518),
.Y(n_1554)
);

NOR2x1_ASAP7_75t_L g1555 ( 
.A(n_1523),
.B(n_1448),
.Y(n_1555)
);

BUFx6f_ASAP7_75t_L g1556 ( 
.A(n_1519),
.Y(n_1556)
);

NAND2xp5_ASAP7_75t_L g1557 ( 
.A(n_1526),
.B(n_1388),
.Y(n_1557)
);

INVxp67_ASAP7_75t_L g1558 ( 
.A(n_1526),
.Y(n_1558)
);

AND2x2_ASAP7_75t_L g1559 ( 
.A(n_1529),
.B(n_1462),
.Y(n_1559)
);

AND2x2_ASAP7_75t_L g1560 ( 
.A(n_1530),
.B(n_1454),
.Y(n_1560)
);

OR2x6_ASAP7_75t_L g1561 ( 
.A(n_1505),
.B(n_1453),
.Y(n_1561)
);

AND2x2_ASAP7_75t_L g1562 ( 
.A(n_1530),
.B(n_1454),
.Y(n_1562)
);

CKINVDCx16_ASAP7_75t_R g1563 ( 
.A(n_1505),
.Y(n_1563)
);

OR2x2_ASAP7_75t_L g1564 ( 
.A(n_1531),
.B(n_1499),
.Y(n_1564)
);

AND2x2_ASAP7_75t_L g1565 ( 
.A(n_1525),
.B(n_1499),
.Y(n_1565)
);

INVx2_ASAP7_75t_L g1566 ( 
.A(n_1532),
.Y(n_1566)
);

OR2x2_ASAP7_75t_L g1567 ( 
.A(n_1534),
.B(n_1512),
.Y(n_1567)
);

INVx1_ASAP7_75t_L g1568 ( 
.A(n_1533),
.Y(n_1568)
);

AND2x2_ASAP7_75t_L g1569 ( 
.A(n_1548),
.B(n_1511),
.Y(n_1569)
);

HB1xp67_ASAP7_75t_L g1570 ( 
.A(n_1546),
.Y(n_1570)
);

INVx3_ASAP7_75t_L g1571 ( 
.A(n_1556),
.Y(n_1571)
);

INVx2_ASAP7_75t_L g1572 ( 
.A(n_1532),
.Y(n_1572)
);

AOI22xp5_ASAP7_75t_L g1573 ( 
.A1(n_1535),
.A2(n_1501),
.B1(n_1516),
.B2(n_1474),
.Y(n_1573)
);

AND2x2_ASAP7_75t_L g1574 ( 
.A(n_1548),
.B(n_1511),
.Y(n_1574)
);

OR2x2_ASAP7_75t_L g1575 ( 
.A(n_1534),
.B(n_1517),
.Y(n_1575)
);

AND2x2_ASAP7_75t_L g1576 ( 
.A(n_1553),
.B(n_1515),
.Y(n_1576)
);

AND2x2_ASAP7_75t_L g1577 ( 
.A(n_1553),
.B(n_1515),
.Y(n_1577)
);

OR2x2_ASAP7_75t_L g1578 ( 
.A(n_1541),
.B(n_1528),
.Y(n_1578)
);

INVx1_ASAP7_75t_L g1579 ( 
.A(n_1533),
.Y(n_1579)
);

AND2x4_ASAP7_75t_L g1580 ( 
.A(n_1555),
.B(n_1508),
.Y(n_1580)
);

OR2x2_ASAP7_75t_L g1581 ( 
.A(n_1541),
.B(n_1517),
.Y(n_1581)
);

AND2x2_ASAP7_75t_L g1582 ( 
.A(n_1559),
.B(n_1558),
.Y(n_1582)
);

INVx1_ASAP7_75t_SL g1583 ( 
.A(n_1543),
.Y(n_1583)
);

NAND2xp33_ASAP7_75t_L g1584 ( 
.A(n_1538),
.B(n_1497),
.Y(n_1584)
);

AND2x2_ASAP7_75t_L g1585 ( 
.A(n_1558),
.B(n_1508),
.Y(n_1585)
);

NAND2x1_ASAP7_75t_L g1586 ( 
.A(n_1555),
.B(n_1520),
.Y(n_1586)
);

NAND2xp5_ASAP7_75t_L g1587 ( 
.A(n_1549),
.B(n_1557),
.Y(n_1587)
);

NAND2xp5_ASAP7_75t_L g1588 ( 
.A(n_1557),
.B(n_1527),
.Y(n_1588)
);

AND2x2_ASAP7_75t_SL g1589 ( 
.A(n_1563),
.B(n_1448),
.Y(n_1589)
);

INVx1_ASAP7_75t_L g1590 ( 
.A(n_1536),
.Y(n_1590)
);

INVx2_ASAP7_75t_SL g1591 ( 
.A(n_1556),
.Y(n_1591)
);

BUFx2_ASAP7_75t_L g1592 ( 
.A(n_1563),
.Y(n_1592)
);

HB1xp67_ASAP7_75t_L g1593 ( 
.A(n_1546),
.Y(n_1593)
);

NAND2xp5_ASAP7_75t_L g1594 ( 
.A(n_1538),
.B(n_1525),
.Y(n_1594)
);

OR2x2_ASAP7_75t_L g1595 ( 
.A(n_1544),
.B(n_1547),
.Y(n_1595)
);

AND2x4_ASAP7_75t_L g1596 ( 
.A(n_1542),
.B(n_1520),
.Y(n_1596)
);

AND2x2_ASAP7_75t_L g1597 ( 
.A(n_1565),
.B(n_1520),
.Y(n_1597)
);

AND2x2_ASAP7_75t_L g1598 ( 
.A(n_1565),
.B(n_1520),
.Y(n_1598)
);

NAND2xp5_ASAP7_75t_SL g1599 ( 
.A(n_1550),
.B(n_1505),
.Y(n_1599)
);

OR2x2_ASAP7_75t_L g1600 ( 
.A(n_1578),
.B(n_1564),
.Y(n_1600)
);

OR2x2_ASAP7_75t_L g1601 ( 
.A(n_1578),
.B(n_1594),
.Y(n_1601)
);

AND2x2_ASAP7_75t_L g1602 ( 
.A(n_1592),
.B(n_1542),
.Y(n_1602)
);

INVx2_ASAP7_75t_L g1603 ( 
.A(n_1566),
.Y(n_1603)
);

OR2x2_ASAP7_75t_L g1604 ( 
.A(n_1594),
.B(n_1564),
.Y(n_1604)
);

AND2x2_ASAP7_75t_L g1605 ( 
.A(n_1592),
.B(n_1542),
.Y(n_1605)
);

INVx1_ASAP7_75t_L g1606 ( 
.A(n_1568),
.Y(n_1606)
);

AND2x2_ASAP7_75t_L g1607 ( 
.A(n_1596),
.B(n_1542),
.Y(n_1607)
);

INVx1_ASAP7_75t_L g1608 ( 
.A(n_1568),
.Y(n_1608)
);

INVx2_ASAP7_75t_L g1609 ( 
.A(n_1566),
.Y(n_1609)
);

OR2x2_ASAP7_75t_L g1610 ( 
.A(n_1587),
.B(n_1547),
.Y(n_1610)
);

INVxp33_ASAP7_75t_SL g1611 ( 
.A(n_1583),
.Y(n_1611)
);

INVx1_ASAP7_75t_L g1612 ( 
.A(n_1579),
.Y(n_1612)
);

OR2x2_ASAP7_75t_L g1613 ( 
.A(n_1587),
.B(n_1552),
.Y(n_1613)
);

OAI222xp33_ASAP7_75t_L g1614 ( 
.A1(n_1573),
.A2(n_1535),
.B1(n_1539),
.B2(n_1545),
.C1(n_1561),
.C2(n_1451),
.Y(n_1614)
);

INVx1_ASAP7_75t_L g1615 ( 
.A(n_1579),
.Y(n_1615)
);

INVx1_ASAP7_75t_L g1616 ( 
.A(n_1590),
.Y(n_1616)
);

INVx1_ASAP7_75t_L g1617 ( 
.A(n_1590),
.Y(n_1617)
);

NAND2xp5_ASAP7_75t_L g1618 ( 
.A(n_1583),
.B(n_1551),
.Y(n_1618)
);

NAND2xp5_ASAP7_75t_L g1619 ( 
.A(n_1588),
.B(n_1551),
.Y(n_1619)
);

AND2x2_ASAP7_75t_L g1620 ( 
.A(n_1596),
.B(n_1560),
.Y(n_1620)
);

NAND2xp5_ASAP7_75t_L g1621 ( 
.A(n_1588),
.B(n_1545),
.Y(n_1621)
);

AND2x2_ASAP7_75t_L g1622 ( 
.A(n_1596),
.B(n_1560),
.Y(n_1622)
);

NOR2x1p5_ASAP7_75t_SL g1623 ( 
.A(n_1566),
.B(n_1554),
.Y(n_1623)
);

HB1xp67_ASAP7_75t_L g1624 ( 
.A(n_1570),
.Y(n_1624)
);

INVx2_ASAP7_75t_L g1625 ( 
.A(n_1572),
.Y(n_1625)
);

OR2x2_ASAP7_75t_L g1626 ( 
.A(n_1595),
.B(n_1567),
.Y(n_1626)
);

NAND2xp5_ASAP7_75t_L g1627 ( 
.A(n_1584),
.B(n_1537),
.Y(n_1627)
);

INVx2_ASAP7_75t_SL g1628 ( 
.A(n_1586),
.Y(n_1628)
);

OR2x2_ASAP7_75t_L g1629 ( 
.A(n_1595),
.B(n_1552),
.Y(n_1629)
);

AND2x2_ASAP7_75t_L g1630 ( 
.A(n_1596),
.B(n_1562),
.Y(n_1630)
);

OAI32xp33_ASAP7_75t_L g1631 ( 
.A1(n_1599),
.A2(n_1550),
.A3(n_1539),
.B1(n_1540),
.B2(n_1440),
.Y(n_1631)
);

INVx2_ASAP7_75t_L g1632 ( 
.A(n_1572),
.Y(n_1632)
);

AOI211xp5_ASAP7_75t_SL g1633 ( 
.A1(n_1573),
.A2(n_1476),
.B(n_1480),
.C(n_1398),
.Y(n_1633)
);

INVx1_ASAP7_75t_L g1634 ( 
.A(n_1570),
.Y(n_1634)
);

INVx1_ASAP7_75t_L g1635 ( 
.A(n_1593),
.Y(n_1635)
);

AND2x2_ASAP7_75t_L g1636 ( 
.A(n_1596),
.B(n_1562),
.Y(n_1636)
);

INVx1_ASAP7_75t_L g1637 ( 
.A(n_1593),
.Y(n_1637)
);

AOI32xp33_ASAP7_75t_L g1638 ( 
.A1(n_1582),
.A2(n_1471),
.A3(n_1466),
.B1(n_1478),
.B2(n_1473),
.Y(n_1638)
);

NAND2x1p5_ASAP7_75t_L g1639 ( 
.A(n_1586),
.B(n_1448),
.Y(n_1639)
);

AND2x2_ASAP7_75t_L g1640 ( 
.A(n_1597),
.B(n_1598),
.Y(n_1640)
);

INVx2_ASAP7_75t_L g1641 ( 
.A(n_1572),
.Y(n_1641)
);

NAND2xp5_ASAP7_75t_L g1642 ( 
.A(n_1576),
.B(n_1524),
.Y(n_1642)
);

OR2x2_ASAP7_75t_L g1643 ( 
.A(n_1601),
.B(n_1567),
.Y(n_1643)
);

INVx1_ASAP7_75t_L g1644 ( 
.A(n_1606),
.Y(n_1644)
);

INVx1_ASAP7_75t_L g1645 ( 
.A(n_1606),
.Y(n_1645)
);

NOR2x1_ASAP7_75t_L g1646 ( 
.A(n_1618),
.B(n_1491),
.Y(n_1646)
);

AND2x2_ASAP7_75t_L g1647 ( 
.A(n_1640),
.B(n_1597),
.Y(n_1647)
);

NAND2xp5_ASAP7_75t_L g1648 ( 
.A(n_1611),
.B(n_1576),
.Y(n_1648)
);

NOR2x1p5_ASAP7_75t_L g1649 ( 
.A(n_1627),
.B(n_1399),
.Y(n_1649)
);

NAND2xp5_ASAP7_75t_L g1650 ( 
.A(n_1638),
.B(n_1576),
.Y(n_1650)
);

NAND2xp5_ASAP7_75t_L g1651 ( 
.A(n_1638),
.B(n_1577),
.Y(n_1651)
);

AND2x2_ASAP7_75t_L g1652 ( 
.A(n_1640),
.B(n_1597),
.Y(n_1652)
);

INVx1_ASAP7_75t_SL g1653 ( 
.A(n_1602),
.Y(n_1653)
);

INVx2_ASAP7_75t_L g1654 ( 
.A(n_1625),
.Y(n_1654)
);

AND2x2_ASAP7_75t_L g1655 ( 
.A(n_1602),
.B(n_1598),
.Y(n_1655)
);

OR2x2_ASAP7_75t_L g1656 ( 
.A(n_1601),
.B(n_1567),
.Y(n_1656)
);

OR2x2_ASAP7_75t_L g1657 ( 
.A(n_1626),
.B(n_1575),
.Y(n_1657)
);

INVx1_ASAP7_75t_L g1658 ( 
.A(n_1608),
.Y(n_1658)
);

AND2x2_ASAP7_75t_L g1659 ( 
.A(n_1605),
.B(n_1598),
.Y(n_1659)
);

NAND2xp5_ASAP7_75t_L g1660 ( 
.A(n_1619),
.B(n_1577),
.Y(n_1660)
);

AND2x4_ASAP7_75t_L g1661 ( 
.A(n_1628),
.B(n_1580),
.Y(n_1661)
);

AND2x4_ASAP7_75t_L g1662 ( 
.A(n_1628),
.B(n_1580),
.Y(n_1662)
);

INVxp67_ASAP7_75t_L g1663 ( 
.A(n_1624),
.Y(n_1663)
);

CKINVDCx16_ASAP7_75t_R g1664 ( 
.A(n_1605),
.Y(n_1664)
);

INVx1_ASAP7_75t_L g1665 ( 
.A(n_1608),
.Y(n_1665)
);

INVx1_ASAP7_75t_L g1666 ( 
.A(n_1612),
.Y(n_1666)
);

OR2x2_ASAP7_75t_L g1667 ( 
.A(n_1626),
.B(n_1575),
.Y(n_1667)
);

INVx1_ASAP7_75t_L g1668 ( 
.A(n_1612),
.Y(n_1668)
);

OR2x2_ASAP7_75t_L g1669 ( 
.A(n_1613),
.B(n_1629),
.Y(n_1669)
);

NAND2xp5_ASAP7_75t_L g1670 ( 
.A(n_1633),
.B(n_1577),
.Y(n_1670)
);

AND2x2_ASAP7_75t_L g1671 ( 
.A(n_1607),
.B(n_1589),
.Y(n_1671)
);

NAND2xp5_ASAP7_75t_L g1672 ( 
.A(n_1621),
.B(n_1582),
.Y(n_1672)
);

AND2x2_ASAP7_75t_L g1673 ( 
.A(n_1607),
.B(n_1589),
.Y(n_1673)
);

INVx1_ASAP7_75t_SL g1674 ( 
.A(n_1610),
.Y(n_1674)
);

NAND2xp5_ASAP7_75t_L g1675 ( 
.A(n_1642),
.B(n_1582),
.Y(n_1675)
);

INVx1_ASAP7_75t_L g1676 ( 
.A(n_1615),
.Y(n_1676)
);

INVx1_ASAP7_75t_L g1677 ( 
.A(n_1615),
.Y(n_1677)
);

OR2x2_ASAP7_75t_L g1678 ( 
.A(n_1613),
.B(n_1575),
.Y(n_1678)
);

NAND2xp5_ASAP7_75t_L g1679 ( 
.A(n_1663),
.B(n_1631),
.Y(n_1679)
);

INVx1_ASAP7_75t_L g1680 ( 
.A(n_1658),
.Y(n_1680)
);

INVxp67_ASAP7_75t_L g1681 ( 
.A(n_1646),
.Y(n_1681)
);

NAND2xp5_ASAP7_75t_L g1682 ( 
.A(n_1653),
.B(n_1631),
.Y(n_1682)
);

AOI22xp5_ASAP7_75t_L g1683 ( 
.A1(n_1664),
.A2(n_1589),
.B1(n_1580),
.B2(n_1637),
.Y(n_1683)
);

INVx1_ASAP7_75t_L g1684 ( 
.A(n_1658),
.Y(n_1684)
);

OAI22xp5_ASAP7_75t_L g1685 ( 
.A1(n_1670),
.A2(n_1639),
.B1(n_1561),
.B2(n_1580),
.Y(n_1685)
);

INVx2_ASAP7_75t_L g1686 ( 
.A(n_1655),
.Y(n_1686)
);

INVx1_ASAP7_75t_L g1687 ( 
.A(n_1644),
.Y(n_1687)
);

INVx1_ASAP7_75t_L g1688 ( 
.A(n_1645),
.Y(n_1688)
);

NAND2xp5_ASAP7_75t_L g1689 ( 
.A(n_1648),
.B(n_1620),
.Y(n_1689)
);

OAI211xp5_ASAP7_75t_L g1690 ( 
.A1(n_1650),
.A2(n_1637),
.B(n_1635),
.C(n_1634),
.Y(n_1690)
);

AOI22xp5_ASAP7_75t_L g1691 ( 
.A1(n_1649),
.A2(n_1580),
.B1(n_1634),
.B2(n_1635),
.Y(n_1691)
);

INVx1_ASAP7_75t_L g1692 ( 
.A(n_1665),
.Y(n_1692)
);

AND2x2_ASAP7_75t_L g1693 ( 
.A(n_1655),
.B(n_1620),
.Y(n_1693)
);

INVx1_ASAP7_75t_L g1694 ( 
.A(n_1666),
.Y(n_1694)
);

INVx1_ASAP7_75t_L g1695 ( 
.A(n_1668),
.Y(n_1695)
);

INVx1_ASAP7_75t_SL g1696 ( 
.A(n_1674),
.Y(n_1696)
);

XNOR2x1_ASAP7_75t_L g1697 ( 
.A(n_1672),
.B(n_1471),
.Y(n_1697)
);

INVx1_ASAP7_75t_L g1698 ( 
.A(n_1676),
.Y(n_1698)
);

INVx1_ASAP7_75t_L g1699 ( 
.A(n_1677),
.Y(n_1699)
);

OAI22xp5_ASAP7_75t_L g1700 ( 
.A1(n_1651),
.A2(n_1639),
.B1(n_1561),
.B2(n_1614),
.Y(n_1700)
);

INVxp67_ASAP7_75t_L g1701 ( 
.A(n_1660),
.Y(n_1701)
);

INVx1_ASAP7_75t_SL g1702 ( 
.A(n_1669),
.Y(n_1702)
);

OAI32xp33_ASAP7_75t_L g1703 ( 
.A1(n_1643),
.A2(n_1639),
.A3(n_1604),
.B1(n_1610),
.B2(n_1600),
.Y(n_1703)
);

AND2x2_ASAP7_75t_L g1704 ( 
.A(n_1659),
.B(n_1622),
.Y(n_1704)
);

INVx1_ASAP7_75t_L g1705 ( 
.A(n_1684),
.Y(n_1705)
);

AOI21xp33_ASAP7_75t_SL g1706 ( 
.A1(n_1681),
.A2(n_1429),
.B(n_1669),
.Y(n_1706)
);

INVx2_ASAP7_75t_L g1707 ( 
.A(n_1693),
.Y(n_1707)
);

AOI221xp5_ASAP7_75t_L g1708 ( 
.A1(n_1679),
.A2(n_1673),
.B1(n_1671),
.B2(n_1643),
.C(n_1656),
.Y(n_1708)
);

NAND2xp5_ASAP7_75t_L g1709 ( 
.A(n_1696),
.B(n_1659),
.Y(n_1709)
);

OA21x2_ASAP7_75t_L g1710 ( 
.A1(n_1690),
.A2(n_1654),
.B(n_1661),
.Y(n_1710)
);

INVx1_ASAP7_75t_L g1711 ( 
.A(n_1684),
.Y(n_1711)
);

NAND4xp25_ASAP7_75t_SL g1712 ( 
.A(n_1682),
.B(n_1673),
.C(n_1671),
.D(n_1675),
.Y(n_1712)
);

INVx1_ASAP7_75t_L g1713 ( 
.A(n_1680),
.Y(n_1713)
);

INVx1_ASAP7_75t_L g1714 ( 
.A(n_1702),
.Y(n_1714)
);

NOR2x1_ASAP7_75t_L g1715 ( 
.A(n_1697),
.B(n_1412),
.Y(n_1715)
);

OAI31xp33_ASAP7_75t_L g1716 ( 
.A1(n_1700),
.A2(n_1662),
.A3(n_1661),
.B(n_1656),
.Y(n_1716)
);

NAND2xp33_ASAP7_75t_L g1717 ( 
.A(n_1691),
.B(n_1657),
.Y(n_1717)
);

INVx3_ASAP7_75t_SL g1718 ( 
.A(n_1697),
.Y(n_1718)
);

AOI222xp33_ASAP7_75t_L g1719 ( 
.A1(n_1701),
.A2(n_1623),
.B1(n_1661),
.B2(n_1662),
.C1(n_1647),
.C2(n_1652),
.Y(n_1719)
);

AOI21xp33_ASAP7_75t_L g1720 ( 
.A1(n_1703),
.A2(n_1667),
.B(n_1657),
.Y(n_1720)
);

A2O1A1Ixp33_ASAP7_75t_L g1721 ( 
.A1(n_1683),
.A2(n_1623),
.B(n_1667),
.C(n_1662),
.Y(n_1721)
);

AND2x2_ASAP7_75t_L g1722 ( 
.A(n_1686),
.B(n_1647),
.Y(n_1722)
);

AOI322xp5_ASAP7_75t_L g1723 ( 
.A1(n_1686),
.A2(n_1652),
.A3(n_1630),
.B1(n_1622),
.B2(n_1636),
.C1(n_1569),
.C2(n_1574),
.Y(n_1723)
);

NOR2xp33_ASAP7_75t_L g1724 ( 
.A(n_1689),
.B(n_1498),
.Y(n_1724)
);

NAND2xp5_ASAP7_75t_L g1725 ( 
.A(n_1714),
.B(n_1687),
.Y(n_1725)
);

NAND2xp5_ASAP7_75t_L g1726 ( 
.A(n_1708),
.B(n_1693),
.Y(n_1726)
);

INVxp67_ASAP7_75t_L g1727 ( 
.A(n_1724),
.Y(n_1727)
);

INVx1_ASAP7_75t_L g1728 ( 
.A(n_1707),
.Y(n_1728)
);

AOI221xp5_ASAP7_75t_L g1729 ( 
.A1(n_1720),
.A2(n_1703),
.B1(n_1685),
.B2(n_1699),
.C(n_1698),
.Y(n_1729)
);

INVx1_ASAP7_75t_L g1730 ( 
.A(n_1705),
.Y(n_1730)
);

INVx1_ASAP7_75t_L g1731 ( 
.A(n_1711),
.Y(n_1731)
);

OAI32xp33_ASAP7_75t_L g1732 ( 
.A1(n_1709),
.A2(n_1695),
.A3(n_1694),
.B1(n_1692),
.B2(n_1688),
.Y(n_1732)
);

AND2x2_ASAP7_75t_L g1733 ( 
.A(n_1722),
.B(n_1704),
.Y(n_1733)
);

INVx1_ASAP7_75t_L g1734 ( 
.A(n_1713),
.Y(n_1734)
);

NAND2xp5_ASAP7_75t_L g1735 ( 
.A(n_1718),
.B(n_1704),
.Y(n_1735)
);

INVx2_ASAP7_75t_L g1736 ( 
.A(n_1733),
.Y(n_1736)
);

AOI21xp5_ASAP7_75t_L g1737 ( 
.A1(n_1729),
.A2(n_1717),
.B(n_1710),
.Y(n_1737)
);

AOI22xp5_ASAP7_75t_L g1738 ( 
.A1(n_1726),
.A2(n_1718),
.B1(n_1712),
.B2(n_1715),
.Y(n_1738)
);

NAND5xp2_ASAP7_75t_L g1739 ( 
.A(n_1735),
.B(n_1716),
.C(n_1724),
.D(n_1719),
.E(n_1721),
.Y(n_1739)
);

NOR2xp33_ASAP7_75t_L g1740 ( 
.A(n_1727),
.B(n_1706),
.Y(n_1740)
);

NAND2xp5_ASAP7_75t_L g1741 ( 
.A(n_1728),
.B(n_1725),
.Y(n_1741)
);

INVx2_ASAP7_75t_L g1742 ( 
.A(n_1730),
.Y(n_1742)
);

NOR3xp33_ASAP7_75t_L g1743 ( 
.A(n_1725),
.B(n_1721),
.C(n_1429),
.Y(n_1743)
);

INVx1_ASAP7_75t_L g1744 ( 
.A(n_1731),
.Y(n_1744)
);

NAND2xp5_ASAP7_75t_SL g1745 ( 
.A(n_1734),
.B(n_1723),
.Y(n_1745)
);

NAND5xp2_ASAP7_75t_L g1746 ( 
.A(n_1738),
.B(n_1732),
.C(n_1710),
.D(n_1498),
.E(n_1479),
.Y(n_1746)
);

OAI31xp33_ASAP7_75t_L g1747 ( 
.A1(n_1737),
.A2(n_1710),
.A3(n_1678),
.B(n_1604),
.Y(n_1747)
);

INVx1_ASAP7_75t_L g1748 ( 
.A(n_1736),
.Y(n_1748)
);

OAI321xp33_ASAP7_75t_L g1749 ( 
.A1(n_1745),
.A2(n_1678),
.A3(n_1654),
.B1(n_1600),
.B2(n_1636),
.C(n_1630),
.Y(n_1749)
);

A2O1A1Ixp33_ASAP7_75t_L g1750 ( 
.A1(n_1743),
.A2(n_1491),
.B(n_1471),
.C(n_1591),
.Y(n_1750)
);

OAI22xp33_ASAP7_75t_SL g1751 ( 
.A1(n_1748),
.A2(n_1741),
.B1(n_1740),
.B2(n_1744),
.Y(n_1751)
);

A2O1A1Ixp33_ASAP7_75t_L g1752 ( 
.A1(n_1747),
.A2(n_1742),
.B(n_1739),
.C(n_1591),
.Y(n_1752)
);

NAND3xp33_ASAP7_75t_SL g1753 ( 
.A(n_1750),
.B(n_1739),
.C(n_1746),
.Y(n_1753)
);

OAI21xp5_ASAP7_75t_L g1754 ( 
.A1(n_1750),
.A2(n_1617),
.B(n_1616),
.Y(n_1754)
);

AOI22xp5_ASAP7_75t_L g1755 ( 
.A1(n_1749),
.A2(n_1428),
.B1(n_1399),
.B2(n_1591),
.Y(n_1755)
);

INVx1_ASAP7_75t_L g1756 ( 
.A(n_1748),
.Y(n_1756)
);

INVx1_ASAP7_75t_SL g1757 ( 
.A(n_1755),
.Y(n_1757)
);

NOR3xp33_ASAP7_75t_L g1758 ( 
.A(n_1753),
.B(n_1428),
.C(n_1472),
.Y(n_1758)
);

NAND4xp75_ASAP7_75t_L g1759 ( 
.A(n_1756),
.B(n_1428),
.C(n_1616),
.D(n_1617),
.Y(n_1759)
);

INVx1_ASAP7_75t_L g1760 ( 
.A(n_1751),
.Y(n_1760)
);

NOR2x1_ASAP7_75t_L g1761 ( 
.A(n_1752),
.B(n_1571),
.Y(n_1761)
);

AND2x4_ASAP7_75t_L g1762 ( 
.A(n_1758),
.B(n_1754),
.Y(n_1762)
);

NOR3xp33_ASAP7_75t_L g1763 ( 
.A(n_1760),
.B(n_1571),
.C(n_1500),
.Y(n_1763)
);

AND4x1_ASAP7_75t_L g1764 ( 
.A(n_1761),
.B(n_1585),
.C(n_1458),
.D(n_1569),
.Y(n_1764)
);

INVx1_ASAP7_75t_L g1765 ( 
.A(n_1762),
.Y(n_1765)
);

INVx1_ASAP7_75t_L g1766 ( 
.A(n_1765),
.Y(n_1766)
);

NOR2x1_ASAP7_75t_L g1767 ( 
.A(n_1766),
.B(n_1759),
.Y(n_1767)
);

AOI21xp5_ASAP7_75t_L g1768 ( 
.A1(n_1766),
.A2(n_1757),
.B(n_1763),
.Y(n_1768)
);

AOI22xp5_ASAP7_75t_L g1769 ( 
.A1(n_1767),
.A2(n_1764),
.B1(n_1571),
.B2(n_1632),
.Y(n_1769)
);

CKINVDCx20_ASAP7_75t_R g1770 ( 
.A(n_1768),
.Y(n_1770)
);

AOI22xp33_ASAP7_75t_L g1771 ( 
.A1(n_1770),
.A2(n_1641),
.B1(n_1632),
.B2(n_1625),
.Y(n_1771)
);

NAND2xp5_ASAP7_75t_L g1772 ( 
.A(n_1769),
.B(n_1603),
.Y(n_1772)
);

AOI21xp5_ASAP7_75t_L g1773 ( 
.A1(n_1772),
.A2(n_1632),
.B(n_1625),
.Y(n_1773)
);

OAI21xp5_ASAP7_75t_L g1774 ( 
.A1(n_1773),
.A2(n_1771),
.B(n_1641),
.Y(n_1774)
);

INVx1_ASAP7_75t_L g1775 ( 
.A(n_1774),
.Y(n_1775)
);

OAI221xp5_ASAP7_75t_R g1776 ( 
.A1(n_1775),
.A2(n_1641),
.B1(n_1609),
.B2(n_1603),
.C(n_1571),
.Y(n_1776)
);

AOI211xp5_ASAP7_75t_L g1777 ( 
.A1(n_1776),
.A2(n_1609),
.B(n_1629),
.C(n_1581),
.Y(n_1777)
);


endmodule