module fake_netlist_6_1710_n_1723 (n_52, n_16, n_1, n_91, n_119, n_46, n_146, n_18, n_21, n_147, n_88, n_3, n_98, n_113, n_39, n_63, n_73, n_4, n_148, n_138, n_22, n_68, n_28, n_50, n_49, n_7, n_83, n_5, n_101, n_144, n_127, n_125, n_153, n_77, n_149, n_152, n_106, n_92, n_145, n_42, n_133, n_96, n_8, n_90, n_24, n_105, n_131, n_54, n_132, n_102, n_0, n_87, n_32, n_66, n_85, n_99, n_78, n_84, n_130, n_100, n_129, n_13, n_121, n_11, n_137, n_17, n_23, n_142, n_20, n_143, n_2, n_19, n_47, n_62, n_29, n_75, n_109, n_150, n_122, n_45, n_34, n_140, n_70, n_120, n_37, n_15, n_67, n_33, n_82, n_27, n_38, n_110, n_151, n_61, n_112, n_81, n_59, n_76, n_36, n_26, n_124, n_55, n_126, n_94, n_97, n_108, n_58, n_116, n_64, n_117, n_118, n_48, n_65, n_25, n_40, n_93, n_80, n_141, n_135, n_139, n_41, n_134, n_114, n_86, n_104, n_95, n_9, n_107, n_10, n_71, n_74, n_6, n_14, n_123, n_136, n_72, n_89, n_103, n_111, n_60, n_35, n_115, n_12, n_69, n_128, n_30, n_79, n_43, n_31, n_57, n_53, n_51, n_44, n_56, n_1723);

input n_52;
input n_16;
input n_1;
input n_91;
input n_119;
input n_46;
input n_146;
input n_18;
input n_21;
input n_147;
input n_88;
input n_3;
input n_98;
input n_113;
input n_39;
input n_63;
input n_73;
input n_4;
input n_148;
input n_138;
input n_22;
input n_68;
input n_28;
input n_50;
input n_49;
input n_7;
input n_83;
input n_5;
input n_101;
input n_144;
input n_127;
input n_125;
input n_153;
input n_77;
input n_149;
input n_152;
input n_106;
input n_92;
input n_145;
input n_42;
input n_133;
input n_96;
input n_8;
input n_90;
input n_24;
input n_105;
input n_131;
input n_54;
input n_132;
input n_102;
input n_0;
input n_87;
input n_32;
input n_66;
input n_85;
input n_99;
input n_78;
input n_84;
input n_130;
input n_100;
input n_129;
input n_13;
input n_121;
input n_11;
input n_137;
input n_17;
input n_23;
input n_142;
input n_20;
input n_143;
input n_2;
input n_19;
input n_47;
input n_62;
input n_29;
input n_75;
input n_109;
input n_150;
input n_122;
input n_45;
input n_34;
input n_140;
input n_70;
input n_120;
input n_37;
input n_15;
input n_67;
input n_33;
input n_82;
input n_27;
input n_38;
input n_110;
input n_151;
input n_61;
input n_112;
input n_81;
input n_59;
input n_76;
input n_36;
input n_26;
input n_124;
input n_55;
input n_126;
input n_94;
input n_97;
input n_108;
input n_58;
input n_116;
input n_64;
input n_117;
input n_118;
input n_48;
input n_65;
input n_25;
input n_40;
input n_93;
input n_80;
input n_141;
input n_135;
input n_139;
input n_41;
input n_134;
input n_114;
input n_86;
input n_104;
input n_95;
input n_9;
input n_107;
input n_10;
input n_71;
input n_74;
input n_6;
input n_14;
input n_123;
input n_136;
input n_72;
input n_89;
input n_103;
input n_111;
input n_60;
input n_35;
input n_115;
input n_12;
input n_69;
input n_128;
input n_30;
input n_79;
input n_43;
input n_31;
input n_57;
input n_53;
input n_51;
input n_44;
input n_56;

output n_1723;

wire n_992;
wire n_1671;
wire n_801;
wire n_1613;
wire n_1234;
wire n_1458;
wire n_1199;
wire n_1674;
wire n_741;
wire n_1027;
wire n_1351;
wire n_625;
wire n_1189;
wire n_223;
wire n_1212;
wire n_226;
wire n_208;
wire n_726;
wire n_212;
wire n_700;
wire n_1307;
wire n_1038;
wire n_578;
wire n_1581;
wire n_1003;
wire n_365;
wire n_168;
wire n_1237;
wire n_1061;
wire n_1357;
wire n_783;
wire n_798;
wire n_188;
wire n_1575;
wire n_509;
wire n_1342;
wire n_245;
wire n_1209;
wire n_1348;
wire n_1387;
wire n_677;
wire n_1708;
wire n_805;
wire n_1151;
wire n_396;
wire n_350;
wire n_1380;
wire n_442;
wire n_480;
wire n_1402;
wire n_1688;
wire n_1691;
wire n_1009;
wire n_1160;
wire n_883;
wire n_1238;
wire n_1032;
wire n_1247;
wire n_1547;
wire n_1553;
wire n_893;
wire n_1099;
wire n_1264;
wire n_1192;
wire n_471;
wire n_424;
wire n_1700;
wire n_1555;
wire n_1415;
wire n_1370;
wire n_369;
wire n_287;
wire n_415;
wire n_830;
wire n_230;
wire n_461;
wire n_873;
wire n_383;
wire n_1285;
wire n_1371;
wire n_200;
wire n_447;
wire n_1172;
wire n_852;
wire n_229;
wire n_1590;
wire n_1532;
wire n_1393;
wire n_1517;
wire n_1704;
wire n_1078;
wire n_250;
wire n_544;
wire n_1711;
wire n_1140;
wire n_1444;
wire n_1670;
wire n_1603;
wire n_1579;
wire n_1263;
wire n_836;
wire n_375;
wire n_522;
wire n_1261;
wire n_945;
wire n_1649;
wire n_1511;
wire n_1143;
wire n_1422;
wire n_1232;
wire n_1572;
wire n_616;
wire n_658;
wire n_1119;
wire n_428;
wire n_1433;
wire n_1620;
wire n_1541;
wire n_1300;
wire n_641;
wire n_822;
wire n_693;
wire n_1313;
wire n_1056;
wire n_758;
wire n_516;
wire n_1455;
wire n_1163;
wire n_1180;
wire n_943;
wire n_1550;
wire n_491;
wire n_1591;
wire n_772;
wire n_1344;
wire n_666;
wire n_371;
wire n_940;
wire n_770;
wire n_567;
wire n_405;
wire n_213;
wire n_538;
wire n_1106;
wire n_886;
wire n_1471;
wire n_343;
wire n_953;
wire n_1094;
wire n_1345;
wire n_494;
wire n_539;
wire n_493;
wire n_155;
wire n_454;
wire n_1421;
wire n_638;
wire n_1404;
wire n_1211;
wire n_381;
wire n_887;
wire n_1660;
wire n_1280;
wire n_713;
wire n_1400;
wire n_1467;
wire n_976;
wire n_224;
wire n_1445;
wire n_1526;
wire n_1560;
wire n_734;
wire n_1088;
wire n_196;
wire n_1231;
wire n_917;
wire n_574;
wire n_907;
wire n_1446;
wire n_659;
wire n_407;
wire n_913;
wire n_1658;
wire n_808;
wire n_867;
wire n_1230;
wire n_473;
wire n_1193;
wire n_1054;
wire n_559;
wire n_1333;
wire n_1648;
wire n_163;
wire n_1644;
wire n_1558;
wire n_281;
wire n_551;
wire n_699;
wire n_564;
wire n_451;
wire n_824;
wire n_279;
wire n_686;
wire n_757;
wire n_594;
wire n_1641;
wire n_577;
wire n_166;
wire n_619;
wire n_1367;
wire n_1336;
wire n_521;
wire n_572;
wire n_395;
wire n_813;
wire n_1481;
wire n_323;
wire n_606;
wire n_1441;
wire n_818;
wire n_1123;
wire n_1309;
wire n_513;
wire n_645;
wire n_1381;
wire n_331;
wire n_1699;
wire n_916;
wire n_483;
wire n_608;
wire n_261;
wire n_630;
wire n_541;
wire n_512;
wire n_433;
wire n_792;
wire n_476;
wire n_1328;
wire n_219;
wire n_264;
wire n_263;
wire n_1162;
wire n_860;
wire n_1530;
wire n_788;
wire n_939;
wire n_1543;
wire n_821;
wire n_938;
wire n_1302;
wire n_1068;
wire n_1599;
wire n_329;
wire n_982;
wire n_549;
wire n_1075;
wire n_408;
wire n_932;
wire n_237;
wire n_1697;
wire n_243;
wire n_979;
wire n_905;
wire n_1680;
wire n_175;
wire n_322;
wire n_993;
wire n_689;
wire n_354;
wire n_1330;
wire n_1413;
wire n_1605;
wire n_1278;
wire n_547;
wire n_558;
wire n_1064;
wire n_1396;
wire n_634;
wire n_966;
wire n_764;
wire n_1663;
wire n_692;
wire n_733;
wire n_1233;
wire n_1289;
wire n_487;
wire n_241;
wire n_1107;
wire n_1014;
wire n_1290;
wire n_1703;
wire n_882;
wire n_1354;
wire n_586;
wire n_423;
wire n_1701;
wire n_318;
wire n_1111;
wire n_1713;
wire n_715;
wire n_1251;
wire n_1265;
wire n_530;
wire n_1563;
wire n_277;
wire n_618;
wire n_1297;
wire n_1662;
wire n_1312;
wire n_199;
wire n_1167;
wire n_1359;
wire n_674;
wire n_871;
wire n_922;
wire n_1335;
wire n_268;
wire n_210;
wire n_1069;
wire n_1664;
wire n_1722;
wire n_612;
wire n_178;
wire n_247;
wire n_1165;
wire n_355;
wire n_702;
wire n_347;
wire n_1175;
wire n_328;
wire n_1386;
wire n_429;
wire n_1012;
wire n_195;
wire n_780;
wire n_675;
wire n_903;
wire n_1540;
wire n_1504;
wire n_286;
wire n_254;
wire n_1655;
wire n_242;
wire n_928;
wire n_835;
wire n_1214;
wire n_690;
wire n_850;
wire n_1654;
wire n_816;
wire n_1157;
wire n_1462;
wire n_1188;
wire n_877;
wire n_604;
wire n_825;
wire n_728;
wire n_1063;
wire n_1588;
wire n_267;
wire n_1124;
wire n_1624;
wire n_515;
wire n_598;
wire n_696;
wire n_1515;
wire n_961;
wire n_437;
wire n_1082;
wire n_1317;
wire n_593;
wire n_514;
wire n_697;
wire n_687;
wire n_890;
wire n_637;
wire n_295;
wire n_701;
wire n_950;
wire n_388;
wire n_190;
wire n_484;
wire n_1709;
wire n_170;
wire n_891;
wire n_1412;
wire n_949;
wire n_1630;
wire n_678;
wire n_283;
wire n_507;
wire n_968;
wire n_909;
wire n_1369;
wire n_881;
wire n_1008;
wire n_760;
wire n_1546;
wire n_590;
wire n_362;
wire n_161;
wire n_462;
wire n_1052;
wire n_1033;
wire n_1296;
wire n_304;
wire n_694;
wire n_1294;
wire n_1420;
wire n_1634;
wire n_297;
wire n_627;
wire n_595;
wire n_524;
wire n_1465;
wire n_342;
wire n_1044;
wire n_1712;
wire n_1391;
wire n_449;
wire n_1523;
wire n_1208;
wire n_1164;
wire n_1295;
wire n_1627;
wire n_1072;
wire n_1527;
wire n_1495;
wire n_1438;
wire n_495;
wire n_815;
wire n_1100;
wire n_585;
wire n_1487;
wire n_840;
wire n_874;
wire n_1128;
wire n_382;
wire n_673;
wire n_1071;
wire n_1067;
wire n_1565;
wire n_1493;
wire n_898;
wire n_255;
wire n_284;
wire n_865;
wire n_925;
wire n_1101;
wire n_1026;
wire n_289;
wire n_1364;
wire n_615;
wire n_1249;
wire n_1293;
wire n_1127;
wire n_1512;
wire n_1451;
wire n_320;
wire n_639;
wire n_963;
wire n_794;
wire n_727;
wire n_894;
wire n_685;
wire n_353;
wire n_605;
wire n_1514;
wire n_826;
wire n_1646;
wire n_872;
wire n_1139;
wire n_1714;
wire n_718;
wire n_1018;
wire n_1521;
wire n_1366;
wire n_542;
wire n_847;
wire n_644;
wire n_682;
wire n_851;
wire n_305;
wire n_996;
wire n_532;
wire n_173;
wire n_1308;
wire n_1376;
wire n_1513;
wire n_413;
wire n_791;
wire n_510;
wire n_837;
wire n_1488;
wire n_948;
wire n_704;
wire n_977;
wire n_1005;
wire n_536;
wire n_622;
wire n_1469;
wire n_581;
wire n_765;
wire n_432;
wire n_987;
wire n_1492;
wire n_1340;
wire n_631;
wire n_720;
wire n_842;
wire n_1707;
wire n_1432;
wire n_156;
wire n_843;
wire n_656;
wire n_989;
wire n_1277;
wire n_797;
wire n_1473;
wire n_1246;
wire n_899;
wire n_189;
wire n_738;
wire n_1304;
wire n_1035;
wire n_294;
wire n_499;
wire n_1426;
wire n_705;
wire n_1004;
wire n_1176;
wire n_1529;
wire n_1022;
wire n_614;
wire n_529;
wire n_425;
wire n_684;
wire n_1431;
wire n_1615;
wire n_1474;
wire n_1571;
wire n_1577;
wire n_1181;
wire n_486;
wire n_947;
wire n_1117;
wire n_1087;
wire n_1448;
wire n_648;
wire n_657;
wire n_1049;
wire n_1666;
wire n_1505;
wire n_803;
wire n_290;
wire n_1717;
wire n_926;
wire n_927;
wire n_919;
wire n_1698;
wire n_478;
wire n_929;
wire n_1228;
wire n_417;
wire n_446;
wire n_1568;
wire n_1490;
wire n_777;
wire n_1299;
wire n_272;
wire n_526;
wire n_1183;
wire n_1436;
wire n_1384;
wire n_293;
wire n_458;
wire n_1070;
wire n_998;
wire n_717;
wire n_1665;
wire n_154;
wire n_1383;
wire n_1178;
wire n_1424;
wire n_1073;
wire n_1000;
wire n_796;
wire n_252;
wire n_1195;
wire n_1626;
wire n_1507;
wire n_184;
wire n_552;
wire n_1358;
wire n_1388;
wire n_216;
wire n_912;
wire n_1519;
wire n_745;
wire n_1284;
wire n_1604;
wire n_1142;
wire n_716;
wire n_1475;
wire n_623;
wire n_1048;
wire n_1201;
wire n_1398;
wire n_884;
wire n_1395;
wire n_731;
wire n_1502;
wire n_1659;
wire n_755;
wire n_931;
wire n_1021;
wire n_474;
wire n_527;
wire n_683;
wire n_811;
wire n_1207;
wire n_312;
wire n_1368;
wire n_1418;
wire n_958;
wire n_292;
wire n_1250;
wire n_1137;
wire n_880;
wire n_889;
wire n_1478;
wire n_589;
wire n_1310;
wire n_819;
wire n_1363;
wire n_1334;
wire n_767;
wire n_1314;
wire n_600;
wire n_964;
wire n_831;
wire n_477;
wire n_954;
wire n_864;
wire n_1110;
wire n_1410;
wire n_399;
wire n_1440;
wire n_1382;
wire n_1534;
wire n_1564;
wire n_211;
wire n_1483;
wire n_1372;
wire n_231;
wire n_1457;
wire n_505;
wire n_1719;
wire n_319;
wire n_1339;
wire n_537;
wire n_1427;
wire n_311;
wire n_1466;
wire n_403;
wire n_1080;
wire n_723;
wire n_596;
wire n_546;
wire n_562;
wire n_1141;
wire n_1268;
wire n_386;
wire n_1220;
wire n_556;
wire n_162;
wire n_1602;
wire n_1136;
wire n_1125;
wire n_970;
wire n_642;
wire n_995;
wire n_276;
wire n_1159;
wire n_1092;
wire n_441;
wire n_221;
wire n_1060;
wire n_444;
wire n_1252;
wire n_1223;
wire n_303;
wire n_511;
wire n_193;
wire n_1286;
wire n_1053;
wire n_416;
wire n_1681;
wire n_520;
wire n_418;
wire n_1093;
wire n_1533;
wire n_1597;
wire n_266;
wire n_296;
wire n_775;
wire n_651;
wire n_1153;
wire n_439;
wire n_1618;
wire n_217;
wire n_518;
wire n_1531;
wire n_1185;
wire n_453;
wire n_215;
wire n_914;
wire n_759;
wire n_426;
wire n_317;
wire n_1653;
wire n_1679;
wire n_1625;
wire n_1453;
wire n_488;
wire n_497;
wire n_773;
wire n_920;
wire n_1374;
wire n_1315;
wire n_1647;
wire n_1224;
wire n_1614;
wire n_1459;
wire n_1135;
wire n_1169;
wire n_1179;
wire n_401;
wire n_324;
wire n_1617;
wire n_335;
wire n_1470;
wire n_463;
wire n_1243;
wire n_848;
wire n_301;
wire n_274;
wire n_1096;
wire n_1091;
wire n_1580;
wire n_1425;
wire n_1267;
wire n_1281;
wire n_983;
wire n_427;
wire n_1520;
wire n_496;
wire n_906;
wire n_1390;
wire n_688;
wire n_1077;
wire n_1419;
wire n_351;
wire n_259;
wire n_177;
wire n_1636;
wire n_1437;
wire n_1645;
wire n_385;
wire n_1687;
wire n_1439;
wire n_1323;
wire n_858;
wire n_1331;
wire n_613;
wire n_736;
wire n_501;
wire n_956;
wire n_960;
wire n_663;
wire n_856;
wire n_379;
wire n_778;
wire n_1668;
wire n_1134;
wire n_410;
wire n_1129;
wire n_554;
wire n_602;
wire n_1696;
wire n_1594;
wire n_664;
wire n_171;
wire n_169;
wire n_1429;
wire n_1610;
wire n_435;
wire n_793;
wire n_326;
wire n_587;
wire n_1593;
wire n_580;
wire n_762;
wire n_1030;
wire n_1202;
wire n_465;
wire n_1635;
wire n_1079;
wire n_341;
wire n_828;
wire n_607;
wire n_316;
wire n_419;
wire n_1551;
wire n_1103;
wire n_1203;
wire n_820;
wire n_951;
wire n_725;
wire n_952;
wire n_999;
wire n_358;
wire n_1254;
wire n_160;
wire n_186;
wire n_368;
wire n_575;
wire n_994;
wire n_1508;
wire n_732;
wire n_974;
wire n_392;
wire n_724;
wire n_1020;
wire n_1042;
wire n_628;
wire n_1273;
wire n_1434;
wire n_1573;
wire n_557;
wire n_349;
wire n_617;
wire n_845;
wire n_807;
wire n_1036;
wire n_1138;
wire n_1661;
wire n_1275;
wire n_485;
wire n_1549;
wire n_443;
wire n_1510;
wire n_892;
wire n_768;
wire n_421;
wire n_1468;
wire n_238;
wire n_1095;
wire n_1595;
wire n_202;
wire n_1718;
wire n_1683;
wire n_597;
wire n_280;
wire n_1270;
wire n_1187;
wire n_610;
wire n_1403;
wire n_1669;
wire n_1024;
wire n_198;
wire n_179;
wire n_248;
wire n_517;
wire n_1667;
wire n_667;
wire n_1206;
wire n_621;
wire n_1037;
wire n_1397;
wire n_1279;
wire n_1115;
wire n_750;
wire n_901;
wire n_1499;
wire n_468;
wire n_923;
wire n_504;
wire n_1409;
wire n_1639;
wire n_1623;
wire n_183;
wire n_1015;
wire n_1503;
wire n_466;
wire n_1057;
wire n_603;
wire n_991;
wire n_1657;
wire n_235;
wire n_1126;
wire n_340;
wire n_710;
wire n_1108;
wire n_1182;
wire n_1298;
wire n_1611;
wire n_785;
wire n_746;
wire n_609;
wire n_1601;
wire n_1686;
wire n_167;
wire n_1356;
wire n_1589;
wire n_1497;
wire n_1168;
wire n_1216;
wire n_1320;
wire n_1430;
wire n_1316;
wire n_1287;
wire n_1452;
wire n_1622;
wire n_1586;
wire n_302;
wire n_1694;
wire n_380;
wire n_1535;
wire n_1596;
wire n_1190;
wire n_397;
wire n_1262;
wire n_218;
wire n_1213;
wire n_1350;
wire n_1673;
wire n_1715;
wire n_172;
wire n_1443;
wire n_1272;
wire n_239;
wire n_782;
wire n_1539;
wire n_490;
wire n_220;
wire n_809;
wire n_1043;
wire n_1608;
wire n_986;
wire n_1472;
wire n_1081;
wire n_402;
wire n_352;
wire n_1692;
wire n_800;
wire n_1084;
wire n_1171;
wire n_460;
wire n_1361;
wire n_1491;
wire n_662;
wire n_374;
wire n_1152;
wire n_1705;
wire n_450;
wire n_1684;
wire n_921;
wire n_1346;
wire n_711;
wire n_1642;
wire n_579;
wire n_1352;
wire n_937;
wire n_1682;
wire n_370;
wire n_1695;
wire n_650;
wire n_1046;
wire n_1145;
wire n_330;
wire n_1121;
wire n_1102;
wire n_972;
wire n_1405;
wire n_258;
wire n_1406;
wire n_456;
wire n_1332;
wire n_260;
wire n_313;
wire n_624;
wire n_962;
wire n_1041;
wire n_565;
wire n_356;
wire n_1569;
wire n_936;
wire n_1288;
wire n_1186;
wire n_1062;
wire n_885;
wire n_896;
wire n_654;
wire n_411;
wire n_1222;
wire n_599;
wire n_776;
wire n_321;
wire n_227;
wire n_1720;
wire n_204;
wire n_482;
wire n_934;
wire n_1637;
wire n_1407;
wire n_420;
wire n_1341;
wire n_394;
wire n_1456;
wire n_1489;
wire n_164;
wire n_942;
wire n_1524;
wire n_543;
wire n_1496;
wire n_1271;
wire n_1545;
wire n_1355;
wire n_1225;
wire n_1544;
wire n_1485;
wire n_325;
wire n_1640;
wire n_804;
wire n_464;
wire n_533;
wire n_806;
wire n_879;
wire n_959;
wire n_584;
wire n_244;
wire n_1343;
wire n_1522;
wire n_548;
wire n_282;
wire n_1676;
wire n_833;
wire n_1567;
wire n_523;
wire n_1319;
wire n_707;
wire n_345;
wire n_799;
wire n_1548;
wire n_1155;
wire n_273;
wire n_1633;
wire n_787;
wire n_1416;
wire n_1528;
wire n_1146;
wire n_159;
wire n_1086;
wire n_1066;
wire n_157;
wire n_1282;
wire n_550;
wire n_275;
wire n_652;
wire n_560;
wire n_1484;
wire n_1241;
wire n_1321;
wire n_1672;
wire n_569;
wire n_737;
wire n_1318;
wire n_1235;
wire n_1229;
wire n_306;
wire n_1292;
wire n_1373;
wire n_346;
wire n_1029;
wire n_1447;
wire n_790;
wire n_1706;
wire n_1498;
wire n_1210;
wire n_299;
wire n_1248;
wire n_1556;
wire n_902;
wire n_333;
wire n_1047;
wire n_1385;
wire n_431;
wire n_459;
wire n_1269;
wire n_502;
wire n_672;
wire n_1257;
wire n_285;
wire n_1375;
wire n_655;
wire n_706;
wire n_1045;
wire n_1650;
wire n_786;
wire n_1236;
wire n_1559;
wire n_834;
wire n_743;
wire n_766;
wire n_430;
wire n_1325;
wire n_1002;
wire n_545;
wire n_489;
wire n_251;
wire n_1019;
wire n_636;
wire n_729;
wire n_876;
wire n_774;
wire n_1337;
wire n_660;
wire n_438;
wire n_1477;
wire n_1360;
wire n_1200;
wire n_479;
wire n_1607;
wire n_1353;
wire n_1454;
wire n_869;
wire n_1154;
wire n_1113;
wire n_1600;
wire n_646;
wire n_528;
wire n_391;
wire n_1098;
wire n_1329;
wire n_817;
wire n_262;
wire n_187;
wire n_897;
wire n_846;
wire n_841;
wire n_1476;
wire n_1001;
wire n_508;
wire n_1050;
wire n_1411;
wire n_1463;
wire n_1177;
wire n_332;
wire n_1150;
wire n_1562;
wire n_1690;
wire n_398;
wire n_1191;
wire n_566;
wire n_1023;
wire n_1076;
wire n_1118;
wire n_194;
wire n_1007;
wire n_1378;
wire n_855;
wire n_1592;
wire n_1631;
wire n_591;
wire n_1377;
wire n_256;
wire n_853;
wire n_440;
wire n_695;
wire n_1542;
wire n_875;
wire n_209;
wire n_367;
wire n_680;
wire n_1678;
wire n_661;
wire n_1716;
wire n_278;
wire n_1256;
wire n_671;
wire n_933;
wire n_740;
wire n_703;
wire n_978;
wire n_384;
wire n_1291;
wire n_1217;
wire n_751;
wire n_749;
wire n_310;
wire n_1628;
wire n_1324;
wire n_1399;
wire n_1435;
wire n_969;
wire n_988;
wire n_1065;
wire n_1401;
wire n_1255;
wire n_568;
wire n_1516;
wire n_1536;
wire n_180;
wire n_1204;
wire n_823;
wire n_1132;
wire n_643;
wire n_233;
wire n_698;
wire n_1074;
wire n_1394;
wire n_1327;
wire n_1326;
wire n_739;
wire n_400;
wire n_955;
wire n_337;
wire n_1379;
wire n_214;
wire n_246;
wire n_1338;
wire n_1097;
wire n_935;
wire n_781;
wire n_789;
wire n_1554;
wire n_1130;
wire n_181;
wire n_182;
wire n_573;
wire n_769;
wire n_676;
wire n_327;
wire n_1120;
wire n_832;
wire n_1583;
wire n_555;
wire n_389;
wire n_814;
wire n_1643;
wire n_669;
wire n_176;
wire n_300;
wire n_222;
wire n_747;
wire n_1389;
wire n_1105;
wire n_721;
wire n_1461;
wire n_742;
wire n_535;
wire n_691;
wire n_372;
wire n_314;
wire n_1408;
wire n_378;
wire n_1196;
wire n_377;
wire n_1598;
wire n_863;
wire n_601;
wire n_338;
wire n_1283;
wire n_918;
wire n_748;
wire n_506;
wire n_1114;
wire n_763;
wire n_1147;
wire n_360;
wire n_1506;
wire n_1652;
wire n_957;
wire n_895;
wire n_866;
wire n_1227;
wire n_191;
wire n_387;
wire n_452;
wire n_744;
wire n_971;
wire n_946;
wire n_344;
wire n_761;
wire n_1303;
wire n_1205;
wire n_1258;
wire n_1392;
wire n_174;
wire n_1173;
wire n_525;
wire n_1677;
wire n_1116;
wire n_611;
wire n_1702;
wire n_1570;
wire n_1219;
wire n_1689;
wire n_1174;
wire n_1016;
wire n_1347;
wire n_795;
wire n_1501;
wire n_1221;
wire n_1245;
wire n_838;
wire n_647;
wire n_197;
wire n_844;
wire n_448;
wire n_1017;
wire n_1083;
wire n_445;
wire n_1561;
wire n_930;
wire n_888;
wire n_1112;
wire n_234;
wire n_910;
wire n_1656;
wire n_1721;
wire n_1460;
wire n_911;
wire n_1464;
wire n_236;
wire n_653;
wire n_1414;
wire n_752;
wire n_908;
wire n_944;
wire n_576;
wire n_1028;
wire n_472;
wire n_270;
wire n_414;
wire n_563;
wire n_1011;
wire n_1566;
wire n_1215;
wire n_839;
wire n_708;
wire n_668;
wire n_626;
wire n_990;
wire n_1500;
wire n_779;
wire n_1537;
wire n_1104;
wire n_854;
wire n_1058;
wire n_498;
wire n_1122;
wire n_870;
wire n_904;
wire n_1253;
wire n_709;
wire n_1266;
wire n_366;
wire n_1509;
wire n_1693;
wire n_1109;
wire n_185;
wire n_712;
wire n_348;
wire n_1276;
wire n_376;
wire n_390;
wire n_1148;
wire n_334;
wire n_1161;
wire n_1085;
wire n_232;
wire n_1239;
wire n_771;
wire n_1584;
wire n_470;
wire n_475;
wire n_924;
wire n_298;
wire n_1582;
wire n_492;
wire n_1149;
wire n_265;
wire n_1184;
wire n_228;
wire n_719;
wire n_1525;
wire n_455;
wire n_1585;
wire n_363;
wire n_1090;
wire n_592;
wire n_1518;
wire n_829;
wire n_1156;
wire n_1362;
wire n_393;
wire n_984;
wire n_503;
wire n_1450;
wire n_1638;
wire n_868;
wire n_570;
wire n_859;
wire n_406;
wire n_735;
wire n_878;
wire n_620;
wire n_519;
wire n_307;
wire n_469;
wire n_1218;
wire n_500;
wire n_1482;
wire n_981;
wire n_714;
wire n_1349;
wire n_291;
wire n_1144;
wire n_357;
wire n_985;
wire n_481;
wire n_997;
wire n_1710;
wire n_1301;
wire n_802;
wire n_561;
wire n_980;
wire n_1306;
wire n_1651;
wire n_1198;
wire n_1609;
wire n_436;
wire n_409;
wire n_1244;
wire n_1685;
wire n_1574;
wire n_240;
wire n_756;
wire n_1619;
wire n_1606;
wire n_810;
wire n_1133;
wire n_635;
wire n_1194;
wire n_1051;
wire n_253;
wire n_1552;
wire n_583;
wire n_249;
wire n_201;
wire n_1039;
wire n_1442;
wire n_1034;
wire n_1480;
wire n_1158;
wire n_754;
wire n_941;
wire n_975;
wire n_1031;
wire n_1305;
wire n_553;
wire n_849;
wire n_753;
wire n_467;
wire n_269;
wire n_359;
wire n_973;
wire n_1479;
wire n_1055;
wire n_1675;
wire n_582;
wire n_861;
wire n_857;
wire n_967;
wire n_571;
wire n_404;
wire n_271;
wire n_158;
wire n_206;
wire n_679;
wire n_633;
wire n_1170;
wire n_665;
wire n_1629;
wire n_588;
wire n_225;
wire n_1260;
wire n_308;
wire n_309;
wire n_1010;
wire n_1040;
wire n_915;
wire n_632;
wire n_1166;
wire n_812;
wire n_1131;
wire n_534;
wire n_1578;
wire n_1006;
wire n_373;
wire n_1632;
wire n_257;
wire n_1557;
wire n_730;
wire n_1311;
wire n_1494;
wire n_670;
wire n_203;
wire n_207;
wire n_1089;
wire n_1587;
wire n_1365;
wire n_1417;
wire n_205;
wire n_1242;
wire n_681;
wire n_1226;
wire n_1274;
wire n_1486;
wire n_412;
wire n_640;
wire n_1322;
wire n_965;
wire n_1428;
wire n_1616;
wire n_1576;
wire n_339;
wire n_784;
wire n_315;
wire n_434;
wire n_288;
wire n_1059;
wire n_1197;
wire n_422;
wire n_722;
wire n_862;
wire n_165;
wire n_540;
wire n_1423;
wire n_457;
wire n_364;
wire n_629;
wire n_1621;
wire n_900;
wire n_1449;
wire n_531;
wire n_827;
wire n_361;
wire n_1025;
wire n_336;
wire n_1013;
wire n_1259;
wire n_192;
wire n_1538;
wire n_649;
wire n_1612;
wire n_1240;

BUFx3_ASAP7_75t_L g154 ( 
.A(n_82),
.Y(n_154)
);

CKINVDCx5p33_ASAP7_75t_R g155 ( 
.A(n_58),
.Y(n_155)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_104),
.Y(n_156)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_69),
.Y(n_157)
);

CKINVDCx5p33_ASAP7_75t_R g158 ( 
.A(n_129),
.Y(n_158)
);

CKINVDCx20_ASAP7_75t_R g159 ( 
.A(n_56),
.Y(n_159)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_49),
.Y(n_160)
);

CKINVDCx5p33_ASAP7_75t_R g161 ( 
.A(n_88),
.Y(n_161)
);

CKINVDCx5p33_ASAP7_75t_R g162 ( 
.A(n_143),
.Y(n_162)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_123),
.Y(n_163)
);

INVx2_ASAP7_75t_L g164 ( 
.A(n_134),
.Y(n_164)
);

HB1xp67_ASAP7_75t_L g165 ( 
.A(n_11),
.Y(n_165)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_8),
.Y(n_166)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_30),
.Y(n_167)
);

HB1xp67_ASAP7_75t_L g168 ( 
.A(n_13),
.Y(n_168)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_107),
.Y(n_169)
);

CKINVDCx5p33_ASAP7_75t_R g170 ( 
.A(n_109),
.Y(n_170)
);

CKINVDCx5p33_ASAP7_75t_R g171 ( 
.A(n_138),
.Y(n_171)
);

INVx1_ASAP7_75t_SL g172 ( 
.A(n_14),
.Y(n_172)
);

CKINVDCx20_ASAP7_75t_R g173 ( 
.A(n_117),
.Y(n_173)
);

CKINVDCx5p33_ASAP7_75t_R g174 ( 
.A(n_38),
.Y(n_174)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_137),
.Y(n_175)
);

BUFx2_ASAP7_75t_L g176 ( 
.A(n_95),
.Y(n_176)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_111),
.Y(n_177)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_26),
.Y(n_178)
);

CKINVDCx5p33_ASAP7_75t_R g179 ( 
.A(n_103),
.Y(n_179)
);

CKINVDCx5p33_ASAP7_75t_R g180 ( 
.A(n_67),
.Y(n_180)
);

CKINVDCx5p33_ASAP7_75t_R g181 ( 
.A(n_93),
.Y(n_181)
);

INVx1_ASAP7_75t_SL g182 ( 
.A(n_28),
.Y(n_182)
);

CKINVDCx5p33_ASAP7_75t_R g183 ( 
.A(n_80),
.Y(n_183)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_46),
.Y(n_184)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_91),
.Y(n_185)
);

CKINVDCx5p33_ASAP7_75t_R g186 ( 
.A(n_83),
.Y(n_186)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_114),
.Y(n_187)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_124),
.Y(n_188)
);

CKINVDCx5p33_ASAP7_75t_R g189 ( 
.A(n_85),
.Y(n_189)
);

CKINVDCx14_ASAP7_75t_R g190 ( 
.A(n_57),
.Y(n_190)
);

BUFx10_ASAP7_75t_L g191 ( 
.A(n_130),
.Y(n_191)
);

CKINVDCx20_ASAP7_75t_R g192 ( 
.A(n_79),
.Y(n_192)
);

BUFx10_ASAP7_75t_L g193 ( 
.A(n_92),
.Y(n_193)
);

CKINVDCx5p33_ASAP7_75t_R g194 ( 
.A(n_151),
.Y(n_194)
);

INVx2_ASAP7_75t_L g195 ( 
.A(n_121),
.Y(n_195)
);

CKINVDCx5p33_ASAP7_75t_R g196 ( 
.A(n_41),
.Y(n_196)
);

CKINVDCx20_ASAP7_75t_R g197 ( 
.A(n_36),
.Y(n_197)
);

CKINVDCx5p33_ASAP7_75t_R g198 ( 
.A(n_96),
.Y(n_198)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_144),
.Y(n_199)
);

CKINVDCx20_ASAP7_75t_R g200 ( 
.A(n_55),
.Y(n_200)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_122),
.Y(n_201)
);

CKINVDCx20_ASAP7_75t_R g202 ( 
.A(n_27),
.Y(n_202)
);

CKINVDCx5p33_ASAP7_75t_R g203 ( 
.A(n_11),
.Y(n_203)
);

CKINVDCx5p33_ASAP7_75t_R g204 ( 
.A(n_61),
.Y(n_204)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_22),
.Y(n_205)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_86),
.Y(n_206)
);

BUFx8_ASAP7_75t_SL g207 ( 
.A(n_102),
.Y(n_207)
);

CKINVDCx5p33_ASAP7_75t_R g208 ( 
.A(n_145),
.Y(n_208)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_136),
.Y(n_209)
);

INVx1_ASAP7_75t_SL g210 ( 
.A(n_24),
.Y(n_210)
);

CKINVDCx14_ASAP7_75t_R g211 ( 
.A(n_127),
.Y(n_211)
);

CKINVDCx5p33_ASAP7_75t_R g212 ( 
.A(n_106),
.Y(n_212)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_77),
.Y(n_213)
);

CKINVDCx5p33_ASAP7_75t_R g214 ( 
.A(n_62),
.Y(n_214)
);

CKINVDCx5p33_ASAP7_75t_R g215 ( 
.A(n_52),
.Y(n_215)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_45),
.Y(n_216)
);

CKINVDCx5p33_ASAP7_75t_R g217 ( 
.A(n_32),
.Y(n_217)
);

CKINVDCx5p33_ASAP7_75t_R g218 ( 
.A(n_75),
.Y(n_218)
);

CKINVDCx5p33_ASAP7_75t_R g219 ( 
.A(n_12),
.Y(n_219)
);

CKINVDCx5p33_ASAP7_75t_R g220 ( 
.A(n_46),
.Y(n_220)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_63),
.Y(n_221)
);

CKINVDCx5p33_ASAP7_75t_R g222 ( 
.A(n_149),
.Y(n_222)
);

INVx2_ASAP7_75t_L g223 ( 
.A(n_34),
.Y(n_223)
);

CKINVDCx5p33_ASAP7_75t_R g224 ( 
.A(n_44),
.Y(n_224)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_21),
.Y(n_225)
);

CKINVDCx5p33_ASAP7_75t_R g226 ( 
.A(n_6),
.Y(n_226)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_66),
.Y(n_227)
);

CKINVDCx5p33_ASAP7_75t_R g228 ( 
.A(n_110),
.Y(n_228)
);

CKINVDCx5p33_ASAP7_75t_R g229 ( 
.A(n_24),
.Y(n_229)
);

CKINVDCx20_ASAP7_75t_R g230 ( 
.A(n_27),
.Y(n_230)
);

INVx2_ASAP7_75t_L g231 ( 
.A(n_19),
.Y(n_231)
);

INVx2_ASAP7_75t_SL g232 ( 
.A(n_148),
.Y(n_232)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_97),
.Y(n_233)
);

CKINVDCx5p33_ASAP7_75t_R g234 ( 
.A(n_10),
.Y(n_234)
);

CKINVDCx5p33_ASAP7_75t_R g235 ( 
.A(n_101),
.Y(n_235)
);

CKINVDCx5p33_ASAP7_75t_R g236 ( 
.A(n_94),
.Y(n_236)
);

CKINVDCx5p33_ASAP7_75t_R g237 ( 
.A(n_8),
.Y(n_237)
);

CKINVDCx5p33_ASAP7_75t_R g238 ( 
.A(n_112),
.Y(n_238)
);

CKINVDCx5p33_ASAP7_75t_R g239 ( 
.A(n_133),
.Y(n_239)
);

CKINVDCx5p33_ASAP7_75t_R g240 ( 
.A(n_98),
.Y(n_240)
);

CKINVDCx5p33_ASAP7_75t_R g241 ( 
.A(n_125),
.Y(n_241)
);

CKINVDCx5p33_ASAP7_75t_R g242 ( 
.A(n_54),
.Y(n_242)
);

INVx2_ASAP7_75t_L g243 ( 
.A(n_50),
.Y(n_243)
);

CKINVDCx5p33_ASAP7_75t_R g244 ( 
.A(n_65),
.Y(n_244)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_30),
.Y(n_245)
);

CKINVDCx5p33_ASAP7_75t_R g246 ( 
.A(n_135),
.Y(n_246)
);

INVx1_ASAP7_75t_SL g247 ( 
.A(n_29),
.Y(n_247)
);

HB1xp67_ASAP7_75t_L g248 ( 
.A(n_18),
.Y(n_248)
);

BUFx8_ASAP7_75t_SL g249 ( 
.A(n_19),
.Y(n_249)
);

BUFx6f_ASAP7_75t_L g250 ( 
.A(n_41),
.Y(n_250)
);

CKINVDCx5p33_ASAP7_75t_R g251 ( 
.A(n_141),
.Y(n_251)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_87),
.Y(n_252)
);

CKINVDCx5p33_ASAP7_75t_R g253 ( 
.A(n_147),
.Y(n_253)
);

CKINVDCx5p33_ASAP7_75t_R g254 ( 
.A(n_5),
.Y(n_254)
);

INVx1_ASAP7_75t_SL g255 ( 
.A(n_84),
.Y(n_255)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_13),
.Y(n_256)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_150),
.Y(n_257)
);

CKINVDCx5p33_ASAP7_75t_R g258 ( 
.A(n_16),
.Y(n_258)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_38),
.Y(n_259)
);

CKINVDCx5p33_ASAP7_75t_R g260 ( 
.A(n_72),
.Y(n_260)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_139),
.Y(n_261)
);

CKINVDCx5p33_ASAP7_75t_R g262 ( 
.A(n_32),
.Y(n_262)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_22),
.Y(n_263)
);

CKINVDCx5p33_ASAP7_75t_R g264 ( 
.A(n_113),
.Y(n_264)
);

HB1xp67_ASAP7_75t_L g265 ( 
.A(n_105),
.Y(n_265)
);

CKINVDCx5p33_ASAP7_75t_R g266 ( 
.A(n_146),
.Y(n_266)
);

INVx2_ASAP7_75t_SL g267 ( 
.A(n_49),
.Y(n_267)
);

INVx1_ASAP7_75t_SL g268 ( 
.A(n_64),
.Y(n_268)
);

CKINVDCx5p33_ASAP7_75t_R g269 ( 
.A(n_7),
.Y(n_269)
);

CKINVDCx5p33_ASAP7_75t_R g270 ( 
.A(n_18),
.Y(n_270)
);

CKINVDCx5p33_ASAP7_75t_R g271 ( 
.A(n_71),
.Y(n_271)
);

BUFx2_ASAP7_75t_L g272 ( 
.A(n_53),
.Y(n_272)
);

CKINVDCx5p33_ASAP7_75t_R g273 ( 
.A(n_59),
.Y(n_273)
);

HB1xp67_ASAP7_75t_L g274 ( 
.A(n_12),
.Y(n_274)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_23),
.Y(n_275)
);

INVx2_ASAP7_75t_L g276 ( 
.A(n_10),
.Y(n_276)
);

CKINVDCx5p33_ASAP7_75t_R g277 ( 
.A(n_17),
.Y(n_277)
);

INVx2_ASAP7_75t_L g278 ( 
.A(n_100),
.Y(n_278)
);

CKINVDCx5p33_ASAP7_75t_R g279 ( 
.A(n_118),
.Y(n_279)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_76),
.Y(n_280)
);

CKINVDCx5p33_ASAP7_75t_R g281 ( 
.A(n_39),
.Y(n_281)
);

BUFx3_ASAP7_75t_L g282 ( 
.A(n_126),
.Y(n_282)
);

CKINVDCx5p33_ASAP7_75t_R g283 ( 
.A(n_4),
.Y(n_283)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_7),
.Y(n_284)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_6),
.Y(n_285)
);

CKINVDCx5p33_ASAP7_75t_R g286 ( 
.A(n_9),
.Y(n_286)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_1),
.Y(n_287)
);

HB1xp67_ASAP7_75t_L g288 ( 
.A(n_153),
.Y(n_288)
);

CKINVDCx5p33_ASAP7_75t_R g289 ( 
.A(n_115),
.Y(n_289)
);

INVx2_ASAP7_75t_L g290 ( 
.A(n_20),
.Y(n_290)
);

CKINVDCx20_ASAP7_75t_R g291 ( 
.A(n_40),
.Y(n_291)
);

INVx2_ASAP7_75t_SL g292 ( 
.A(n_14),
.Y(n_292)
);

CKINVDCx5p33_ASAP7_75t_R g293 ( 
.A(n_4),
.Y(n_293)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_81),
.Y(n_294)
);

CKINVDCx5p33_ASAP7_75t_R g295 ( 
.A(n_48),
.Y(n_295)
);

CKINVDCx5p33_ASAP7_75t_R g296 ( 
.A(n_68),
.Y(n_296)
);

CKINVDCx5p33_ASAP7_75t_R g297 ( 
.A(n_1),
.Y(n_297)
);

CKINVDCx5p33_ASAP7_75t_R g298 ( 
.A(n_152),
.Y(n_298)
);

CKINVDCx5p33_ASAP7_75t_R g299 ( 
.A(n_20),
.Y(n_299)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_37),
.Y(n_300)
);

CKINVDCx16_ASAP7_75t_R g301 ( 
.A(n_31),
.Y(n_301)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_131),
.Y(n_302)
);

BUFx2_ASAP7_75t_L g303 ( 
.A(n_33),
.Y(n_303)
);

CKINVDCx5p33_ASAP7_75t_R g304 ( 
.A(n_21),
.Y(n_304)
);

CKINVDCx5p33_ASAP7_75t_R g305 ( 
.A(n_16),
.Y(n_305)
);

CKINVDCx5p33_ASAP7_75t_R g306 ( 
.A(n_116),
.Y(n_306)
);

CKINVDCx20_ASAP7_75t_R g307 ( 
.A(n_159),
.Y(n_307)
);

CKINVDCx20_ASAP7_75t_R g308 ( 
.A(n_173),
.Y(n_308)
);

CKINVDCx5p33_ASAP7_75t_R g309 ( 
.A(n_207),
.Y(n_309)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_250),
.Y(n_310)
);

INVxp67_ASAP7_75t_SL g311 ( 
.A(n_265),
.Y(n_311)
);

BUFx3_ASAP7_75t_L g312 ( 
.A(n_154),
.Y(n_312)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_250),
.Y(n_313)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_250),
.Y(n_314)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_250),
.Y(n_315)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_250),
.Y(n_316)
);

CKINVDCx20_ASAP7_75t_R g317 ( 
.A(n_192),
.Y(n_317)
);

CKINVDCx5p33_ASAP7_75t_R g318 ( 
.A(n_249),
.Y(n_318)
);

INVxp67_ASAP7_75t_SL g319 ( 
.A(n_288),
.Y(n_319)
);

CKINVDCx20_ASAP7_75t_R g320 ( 
.A(n_200),
.Y(n_320)
);

CKINVDCx20_ASAP7_75t_R g321 ( 
.A(n_190),
.Y(n_321)
);

INVxp67_ASAP7_75t_SL g322 ( 
.A(n_176),
.Y(n_322)
);

CKINVDCx5p33_ASAP7_75t_R g323 ( 
.A(n_155),
.Y(n_323)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_250),
.Y(n_324)
);

INVxp67_ASAP7_75t_SL g325 ( 
.A(n_176),
.Y(n_325)
);

CKINVDCx5p33_ASAP7_75t_R g326 ( 
.A(n_158),
.Y(n_326)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_276),
.Y(n_327)
);

CKINVDCx5p33_ASAP7_75t_R g328 ( 
.A(n_161),
.Y(n_328)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_276),
.Y(n_329)
);

INVx2_ASAP7_75t_L g330 ( 
.A(n_164),
.Y(n_330)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_276),
.Y(n_331)
);

INVxp67_ASAP7_75t_L g332 ( 
.A(n_303),
.Y(n_332)
);

CKINVDCx5p33_ASAP7_75t_R g333 ( 
.A(n_162),
.Y(n_333)
);

HB1xp67_ASAP7_75t_L g334 ( 
.A(n_303),
.Y(n_334)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_223),
.Y(n_335)
);

CKINVDCx5p33_ASAP7_75t_R g336 ( 
.A(n_170),
.Y(n_336)
);

CKINVDCx20_ASAP7_75t_R g337 ( 
.A(n_211),
.Y(n_337)
);

INVx1_ASAP7_75t_L g338 ( 
.A(n_223),
.Y(n_338)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_231),
.Y(n_339)
);

CKINVDCx5p33_ASAP7_75t_R g340 ( 
.A(n_171),
.Y(n_340)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_231),
.Y(n_341)
);

INVx1_ASAP7_75t_L g342 ( 
.A(n_243),
.Y(n_342)
);

INVxp67_ASAP7_75t_L g343 ( 
.A(n_165),
.Y(n_343)
);

HB1xp67_ASAP7_75t_L g344 ( 
.A(n_301),
.Y(n_344)
);

INVx1_ASAP7_75t_L g345 ( 
.A(n_243),
.Y(n_345)
);

INVx1_ASAP7_75t_L g346 ( 
.A(n_290),
.Y(n_346)
);

INVx1_ASAP7_75t_L g347 ( 
.A(n_290),
.Y(n_347)
);

INVx1_ASAP7_75t_L g348 ( 
.A(n_160),
.Y(n_348)
);

INVx1_ASAP7_75t_L g349 ( 
.A(n_160),
.Y(n_349)
);

INVx1_ASAP7_75t_L g350 ( 
.A(n_166),
.Y(n_350)
);

CKINVDCx5p33_ASAP7_75t_R g351 ( 
.A(n_179),
.Y(n_351)
);

CKINVDCx20_ASAP7_75t_R g352 ( 
.A(n_180),
.Y(n_352)
);

CKINVDCx14_ASAP7_75t_R g353 ( 
.A(n_272),
.Y(n_353)
);

INVx1_ASAP7_75t_L g354 ( 
.A(n_166),
.Y(n_354)
);

INVx1_ASAP7_75t_L g355 ( 
.A(n_167),
.Y(n_355)
);

INVxp67_ASAP7_75t_SL g356 ( 
.A(n_272),
.Y(n_356)
);

CKINVDCx20_ASAP7_75t_R g357 ( 
.A(n_181),
.Y(n_357)
);

INVx1_ASAP7_75t_L g358 ( 
.A(n_167),
.Y(n_358)
);

INVx1_ASAP7_75t_L g359 ( 
.A(n_178),
.Y(n_359)
);

CKINVDCx20_ASAP7_75t_R g360 ( 
.A(n_183),
.Y(n_360)
);

INVx1_ASAP7_75t_L g361 ( 
.A(n_178),
.Y(n_361)
);

INVxp33_ASAP7_75t_L g362 ( 
.A(n_168),
.Y(n_362)
);

BUFx3_ASAP7_75t_L g363 ( 
.A(n_154),
.Y(n_363)
);

INVx1_ASAP7_75t_L g364 ( 
.A(n_184),
.Y(n_364)
);

CKINVDCx14_ASAP7_75t_R g365 ( 
.A(n_191),
.Y(n_365)
);

CKINVDCx5p33_ASAP7_75t_R g366 ( 
.A(n_186),
.Y(n_366)
);

INVx1_ASAP7_75t_L g367 ( 
.A(n_184),
.Y(n_367)
);

CKINVDCx20_ASAP7_75t_R g368 ( 
.A(n_189),
.Y(n_368)
);

CKINVDCx16_ASAP7_75t_R g369 ( 
.A(n_301),
.Y(n_369)
);

INVx1_ASAP7_75t_L g370 ( 
.A(n_205),
.Y(n_370)
);

INVxp67_ASAP7_75t_SL g371 ( 
.A(n_154),
.Y(n_371)
);

INVxp33_ASAP7_75t_L g372 ( 
.A(n_248),
.Y(n_372)
);

INVxp67_ASAP7_75t_SL g373 ( 
.A(n_282),
.Y(n_373)
);

CKINVDCx20_ASAP7_75t_R g374 ( 
.A(n_194),
.Y(n_374)
);

INVx1_ASAP7_75t_L g375 ( 
.A(n_205),
.Y(n_375)
);

CKINVDCx14_ASAP7_75t_R g376 ( 
.A(n_191),
.Y(n_376)
);

AND2x4_ASAP7_75t_L g377 ( 
.A(n_310),
.B(n_282),
.Y(n_377)
);

INVx1_ASAP7_75t_L g378 ( 
.A(n_310),
.Y(n_378)
);

NAND2xp5_ASAP7_75t_L g379 ( 
.A(n_371),
.B(n_232),
.Y(n_379)
);

INVx2_ASAP7_75t_L g380 ( 
.A(n_330),
.Y(n_380)
);

BUFx2_ASAP7_75t_L g381 ( 
.A(n_353),
.Y(n_381)
);

AOI22xp5_ASAP7_75t_L g382 ( 
.A1(n_369),
.A2(n_202),
.B1(n_230),
.B2(n_197),
.Y(n_382)
);

INVx1_ASAP7_75t_L g383 ( 
.A(n_313),
.Y(n_383)
);

AND2x2_ASAP7_75t_L g384 ( 
.A(n_373),
.B(n_282),
.Y(n_384)
);

HB1xp67_ASAP7_75t_L g385 ( 
.A(n_344),
.Y(n_385)
);

AND2x2_ASAP7_75t_L g386 ( 
.A(n_312),
.B(n_164),
.Y(n_386)
);

NAND2xp5_ASAP7_75t_L g387 ( 
.A(n_312),
.B(n_232),
.Y(n_387)
);

INVx1_ASAP7_75t_L g388 ( 
.A(n_313),
.Y(n_388)
);

INVx2_ASAP7_75t_L g389 ( 
.A(n_314),
.Y(n_389)
);

INVx3_ASAP7_75t_L g390 ( 
.A(n_330),
.Y(n_390)
);

BUFx6f_ASAP7_75t_L g391 ( 
.A(n_330),
.Y(n_391)
);

BUFx6f_ASAP7_75t_L g392 ( 
.A(n_314),
.Y(n_392)
);

INVx1_ASAP7_75t_L g393 ( 
.A(n_315),
.Y(n_393)
);

CKINVDCx16_ASAP7_75t_R g394 ( 
.A(n_369),
.Y(n_394)
);

INVx2_ASAP7_75t_L g395 ( 
.A(n_315),
.Y(n_395)
);

HB1xp67_ASAP7_75t_L g396 ( 
.A(n_334),
.Y(n_396)
);

HB1xp67_ASAP7_75t_L g397 ( 
.A(n_312),
.Y(n_397)
);

NOR2xp33_ASAP7_75t_L g398 ( 
.A(n_322),
.B(n_255),
.Y(n_398)
);

INVx2_ASAP7_75t_L g399 ( 
.A(n_316),
.Y(n_399)
);

INVx2_ASAP7_75t_L g400 ( 
.A(n_316),
.Y(n_400)
);

INVx2_ASAP7_75t_L g401 ( 
.A(n_324),
.Y(n_401)
);

INVx1_ASAP7_75t_L g402 ( 
.A(n_324),
.Y(n_402)
);

INVx1_ASAP7_75t_L g403 ( 
.A(n_348),
.Y(n_403)
);

OA21x2_ASAP7_75t_L g404 ( 
.A1(n_327),
.A2(n_225),
.B(n_216),
.Y(n_404)
);

BUFx2_ASAP7_75t_L g405 ( 
.A(n_363),
.Y(n_405)
);

NOR2xp33_ASAP7_75t_L g406 ( 
.A(n_325),
.B(n_268),
.Y(n_406)
);

BUFx6f_ASAP7_75t_L g407 ( 
.A(n_327),
.Y(n_407)
);

INVx1_ASAP7_75t_L g408 ( 
.A(n_348),
.Y(n_408)
);

INVx2_ASAP7_75t_L g409 ( 
.A(n_329),
.Y(n_409)
);

OR2x2_ASAP7_75t_L g410 ( 
.A(n_363),
.B(n_332),
.Y(n_410)
);

INVx1_ASAP7_75t_L g411 ( 
.A(n_349),
.Y(n_411)
);

NAND2xp5_ASAP7_75t_L g412 ( 
.A(n_363),
.B(n_306),
.Y(n_412)
);

BUFx6f_ASAP7_75t_L g413 ( 
.A(n_329),
.Y(n_413)
);

INVx1_ASAP7_75t_L g414 ( 
.A(n_349),
.Y(n_414)
);

NAND2xp5_ASAP7_75t_L g415 ( 
.A(n_350),
.B(n_198),
.Y(n_415)
);

INVx1_ASAP7_75t_L g416 ( 
.A(n_350),
.Y(n_416)
);

NOR2xp33_ASAP7_75t_R g417 ( 
.A(n_365),
.B(n_204),
.Y(n_417)
);

OAI22xp5_ASAP7_75t_L g418 ( 
.A1(n_343),
.A2(n_291),
.B1(n_274),
.B2(n_172),
.Y(n_418)
);

INVx1_ASAP7_75t_L g419 ( 
.A(n_354),
.Y(n_419)
);

BUFx8_ASAP7_75t_L g420 ( 
.A(n_376),
.Y(n_420)
);

INVx2_ASAP7_75t_L g421 ( 
.A(n_331),
.Y(n_421)
);

INVx1_ASAP7_75t_L g422 ( 
.A(n_354),
.Y(n_422)
);

AND2x2_ASAP7_75t_L g423 ( 
.A(n_331),
.B(n_164),
.Y(n_423)
);

AND2x4_ASAP7_75t_SL g424 ( 
.A(n_352),
.B(n_191),
.Y(n_424)
);

INVx2_ASAP7_75t_L g425 ( 
.A(n_335),
.Y(n_425)
);

INVx1_ASAP7_75t_L g426 ( 
.A(n_355),
.Y(n_426)
);

CKINVDCx5p33_ASAP7_75t_R g427 ( 
.A(n_323),
.Y(n_427)
);

INVx2_ASAP7_75t_L g428 ( 
.A(n_335),
.Y(n_428)
);

INVx2_ASAP7_75t_L g429 ( 
.A(n_338),
.Y(n_429)
);

INVx1_ASAP7_75t_L g430 ( 
.A(n_355),
.Y(n_430)
);

INVx1_ASAP7_75t_L g431 ( 
.A(n_358),
.Y(n_431)
);

NAND2xp5_ASAP7_75t_L g432 ( 
.A(n_358),
.B(n_359),
.Y(n_432)
);

INVxp67_ASAP7_75t_SL g433 ( 
.A(n_359),
.Y(n_433)
);

AND2x4_ASAP7_75t_L g434 ( 
.A(n_361),
.B(n_278),
.Y(n_434)
);

NAND2xp5_ASAP7_75t_L g435 ( 
.A(n_361),
.B(n_208),
.Y(n_435)
);

INVx2_ASAP7_75t_L g436 ( 
.A(n_338),
.Y(n_436)
);

BUFx6f_ASAP7_75t_L g437 ( 
.A(n_339),
.Y(n_437)
);

OAI21x1_ASAP7_75t_L g438 ( 
.A1(n_364),
.A2(n_278),
.B(n_195),
.Y(n_438)
);

AND2x4_ASAP7_75t_L g439 ( 
.A(n_364),
.B(n_195),
.Y(n_439)
);

AND2x2_ASAP7_75t_L g440 ( 
.A(n_356),
.B(n_339),
.Y(n_440)
);

INVx1_ASAP7_75t_L g441 ( 
.A(n_367),
.Y(n_441)
);

INVx2_ASAP7_75t_L g442 ( 
.A(n_389),
.Y(n_442)
);

INVx2_ASAP7_75t_L g443 ( 
.A(n_389),
.Y(n_443)
);

INVx2_ASAP7_75t_L g444 ( 
.A(n_389),
.Y(n_444)
);

INVx1_ASAP7_75t_L g445 ( 
.A(n_404),
.Y(n_445)
);

INVx1_ASAP7_75t_L g446 ( 
.A(n_404),
.Y(n_446)
);

INVx1_ASAP7_75t_L g447 ( 
.A(n_404),
.Y(n_447)
);

BUFx6f_ASAP7_75t_L g448 ( 
.A(n_404),
.Y(n_448)
);

AOI22xp33_ASAP7_75t_L g449 ( 
.A1(n_384),
.A2(n_319),
.B1(n_311),
.B2(n_267),
.Y(n_449)
);

INVx3_ASAP7_75t_L g450 ( 
.A(n_391),
.Y(n_450)
);

INVx1_ASAP7_75t_L g451 ( 
.A(n_404),
.Y(n_451)
);

NAND2xp5_ASAP7_75t_SL g452 ( 
.A(n_420),
.B(n_326),
.Y(n_452)
);

HB1xp67_ASAP7_75t_L g453 ( 
.A(n_397),
.Y(n_453)
);

INVx1_ASAP7_75t_SL g454 ( 
.A(n_381),
.Y(n_454)
);

INVx1_ASAP7_75t_L g455 ( 
.A(n_404),
.Y(n_455)
);

INVx1_ASAP7_75t_L g456 ( 
.A(n_378),
.Y(n_456)
);

INVx2_ASAP7_75t_L g457 ( 
.A(n_395),
.Y(n_457)
);

BUFx3_ASAP7_75t_L g458 ( 
.A(n_405),
.Y(n_458)
);

AOI22xp5_ASAP7_75t_L g459 ( 
.A1(n_398),
.A2(n_406),
.B1(n_360),
.B2(n_368),
.Y(n_459)
);

INVx3_ASAP7_75t_L g460 ( 
.A(n_391),
.Y(n_460)
);

INVx2_ASAP7_75t_L g461 ( 
.A(n_395),
.Y(n_461)
);

NOR2xp33_ASAP7_75t_L g462 ( 
.A(n_405),
.B(n_328),
.Y(n_462)
);

NAND2xp5_ASAP7_75t_L g463 ( 
.A(n_405),
.B(n_333),
.Y(n_463)
);

INVx2_ASAP7_75t_L g464 ( 
.A(n_395),
.Y(n_464)
);

INVx2_ASAP7_75t_L g465 ( 
.A(n_395),
.Y(n_465)
);

INVx2_ASAP7_75t_L g466 ( 
.A(n_399),
.Y(n_466)
);

AND2x2_ASAP7_75t_L g467 ( 
.A(n_384),
.B(n_341),
.Y(n_467)
);

NAND2xp33_ASAP7_75t_L g468 ( 
.A(n_397),
.B(n_195),
.Y(n_468)
);

INVx2_ASAP7_75t_L g469 ( 
.A(n_399),
.Y(n_469)
);

INVx1_ASAP7_75t_L g470 ( 
.A(n_378),
.Y(n_470)
);

AOI22xp5_ASAP7_75t_L g471 ( 
.A1(n_398),
.A2(n_357),
.B1(n_374),
.B2(n_366),
.Y(n_471)
);

INVx1_ASAP7_75t_L g472 ( 
.A(n_383),
.Y(n_472)
);

NOR2xp33_ASAP7_75t_L g473 ( 
.A(n_406),
.B(n_336),
.Y(n_473)
);

CKINVDCx5p33_ASAP7_75t_R g474 ( 
.A(n_417),
.Y(n_474)
);

INVx1_ASAP7_75t_L g475 ( 
.A(n_383),
.Y(n_475)
);

INVx4_ASAP7_75t_L g476 ( 
.A(n_392),
.Y(n_476)
);

INVx2_ASAP7_75t_L g477 ( 
.A(n_399),
.Y(n_477)
);

INVx1_ASAP7_75t_L g478 ( 
.A(n_388),
.Y(n_478)
);

NAND2xp5_ASAP7_75t_SL g479 ( 
.A(n_420),
.B(n_340),
.Y(n_479)
);

INVx2_ASAP7_75t_L g480 ( 
.A(n_399),
.Y(n_480)
);

NAND2xp5_ASAP7_75t_L g481 ( 
.A(n_412),
.B(n_351),
.Y(n_481)
);

INVx2_ASAP7_75t_SL g482 ( 
.A(n_410),
.Y(n_482)
);

INVx4_ASAP7_75t_L g483 ( 
.A(n_392),
.Y(n_483)
);

INVx1_ASAP7_75t_L g484 ( 
.A(n_388),
.Y(n_484)
);

INVx1_ASAP7_75t_L g485 ( 
.A(n_393),
.Y(n_485)
);

NOR2xp33_ASAP7_75t_L g486 ( 
.A(n_427),
.B(n_321),
.Y(n_486)
);

INVx2_ASAP7_75t_L g487 ( 
.A(n_400),
.Y(n_487)
);

INVx3_ASAP7_75t_L g488 ( 
.A(n_391),
.Y(n_488)
);

NAND2xp5_ASAP7_75t_L g489 ( 
.A(n_384),
.B(n_212),
.Y(n_489)
);

BUFx2_ASAP7_75t_L g490 ( 
.A(n_385),
.Y(n_490)
);

NOR2x1p5_ASAP7_75t_L g491 ( 
.A(n_433),
.B(n_309),
.Y(n_491)
);

INVx2_ASAP7_75t_L g492 ( 
.A(n_400),
.Y(n_492)
);

INVxp33_ASAP7_75t_SL g493 ( 
.A(n_417),
.Y(n_493)
);

NAND2xp5_ASAP7_75t_SL g494 ( 
.A(n_420),
.B(n_337),
.Y(n_494)
);

INVx1_ASAP7_75t_L g495 ( 
.A(n_393),
.Y(n_495)
);

INVx1_ASAP7_75t_L g496 ( 
.A(n_402),
.Y(n_496)
);

NAND2xp5_ASAP7_75t_SL g497 ( 
.A(n_420),
.B(n_318),
.Y(n_497)
);

INVx2_ASAP7_75t_L g498 ( 
.A(n_400),
.Y(n_498)
);

INVx1_ASAP7_75t_L g499 ( 
.A(n_402),
.Y(n_499)
);

OR2x6_ASAP7_75t_L g500 ( 
.A(n_410),
.B(n_267),
.Y(n_500)
);

NOR2xp33_ASAP7_75t_L g501 ( 
.A(n_410),
.B(n_362),
.Y(n_501)
);

NAND2xp5_ASAP7_75t_SL g502 ( 
.A(n_420),
.B(n_191),
.Y(n_502)
);

INVx1_ASAP7_75t_L g503 ( 
.A(n_403),
.Y(n_503)
);

INVx3_ASAP7_75t_L g504 ( 
.A(n_391),
.Y(n_504)
);

NAND2xp5_ASAP7_75t_SL g505 ( 
.A(n_381),
.B(n_193),
.Y(n_505)
);

INVx3_ASAP7_75t_L g506 ( 
.A(n_391),
.Y(n_506)
);

INVx2_ASAP7_75t_SL g507 ( 
.A(n_440),
.Y(n_507)
);

NAND2xp5_ASAP7_75t_L g508 ( 
.A(n_386),
.B(n_214),
.Y(n_508)
);

INVx1_ASAP7_75t_L g509 ( 
.A(n_403),
.Y(n_509)
);

INVx2_ASAP7_75t_L g510 ( 
.A(n_400),
.Y(n_510)
);

INVx2_ASAP7_75t_L g511 ( 
.A(n_401),
.Y(n_511)
);

INVx4_ASAP7_75t_L g512 ( 
.A(n_392),
.Y(n_512)
);

INVx2_ASAP7_75t_L g513 ( 
.A(n_401),
.Y(n_513)
);

INVx3_ASAP7_75t_L g514 ( 
.A(n_391),
.Y(n_514)
);

NAND2xp5_ASAP7_75t_L g515 ( 
.A(n_386),
.B(n_379),
.Y(n_515)
);

INVx1_ASAP7_75t_L g516 ( 
.A(n_408),
.Y(n_516)
);

NOR2x1p5_ASAP7_75t_L g517 ( 
.A(n_433),
.B(n_174),
.Y(n_517)
);

INVx1_ASAP7_75t_L g518 ( 
.A(n_408),
.Y(n_518)
);

INVx2_ASAP7_75t_L g519 ( 
.A(n_401),
.Y(n_519)
);

BUFx6f_ASAP7_75t_L g520 ( 
.A(n_438),
.Y(n_520)
);

INVx1_ASAP7_75t_L g521 ( 
.A(n_411),
.Y(n_521)
);

NOR2xp33_ASAP7_75t_L g522 ( 
.A(n_379),
.B(n_372),
.Y(n_522)
);

NOR2xp33_ASAP7_75t_L g523 ( 
.A(n_415),
.B(n_307),
.Y(n_523)
);

INVx1_ASAP7_75t_L g524 ( 
.A(n_411),
.Y(n_524)
);

INVx1_ASAP7_75t_L g525 ( 
.A(n_414),
.Y(n_525)
);

INVx2_ASAP7_75t_SL g526 ( 
.A(n_440),
.Y(n_526)
);

NAND2xp5_ASAP7_75t_SL g527 ( 
.A(n_381),
.B(n_193),
.Y(n_527)
);

CKINVDCx6p67_ASAP7_75t_R g528 ( 
.A(n_394),
.Y(n_528)
);

INVx2_ASAP7_75t_L g529 ( 
.A(n_401),
.Y(n_529)
);

INVx3_ASAP7_75t_L g530 ( 
.A(n_391),
.Y(n_530)
);

INVx2_ASAP7_75t_L g531 ( 
.A(n_380),
.Y(n_531)
);

INVx4_ASAP7_75t_L g532 ( 
.A(n_392),
.Y(n_532)
);

INVx2_ASAP7_75t_L g533 ( 
.A(n_380),
.Y(n_533)
);

INVx2_ASAP7_75t_L g534 ( 
.A(n_380),
.Y(n_534)
);

CKINVDCx5p33_ASAP7_75t_R g535 ( 
.A(n_394),
.Y(n_535)
);

NAND2xp5_ASAP7_75t_SL g536 ( 
.A(n_440),
.B(n_193),
.Y(n_536)
);

NAND2xp5_ASAP7_75t_L g537 ( 
.A(n_386),
.B(n_215),
.Y(n_537)
);

INVx2_ASAP7_75t_L g538 ( 
.A(n_380),
.Y(n_538)
);

INVx2_ASAP7_75t_L g539 ( 
.A(n_390),
.Y(n_539)
);

INVx1_ASAP7_75t_L g540 ( 
.A(n_414),
.Y(n_540)
);

NAND2xp5_ASAP7_75t_SL g541 ( 
.A(n_415),
.B(n_193),
.Y(n_541)
);

INVx1_ASAP7_75t_L g542 ( 
.A(n_416),
.Y(n_542)
);

INVx1_ASAP7_75t_L g543 ( 
.A(n_416),
.Y(n_543)
);

OR2x6_ASAP7_75t_L g544 ( 
.A(n_387),
.B(n_292),
.Y(n_544)
);

BUFx6f_ASAP7_75t_L g545 ( 
.A(n_438),
.Y(n_545)
);

OR2x6_ASAP7_75t_L g546 ( 
.A(n_387),
.B(n_292),
.Y(n_546)
);

NOR2xp33_ASAP7_75t_L g547 ( 
.A(n_435),
.B(n_385),
.Y(n_547)
);

BUFx6f_ASAP7_75t_SL g548 ( 
.A(n_377),
.Y(n_548)
);

INVx2_ASAP7_75t_L g549 ( 
.A(n_390),
.Y(n_549)
);

INVx3_ASAP7_75t_L g550 ( 
.A(n_391),
.Y(n_550)
);

INVx1_ASAP7_75t_L g551 ( 
.A(n_419),
.Y(n_551)
);

INVx2_ASAP7_75t_L g552 ( 
.A(n_390),
.Y(n_552)
);

NAND2xp5_ASAP7_75t_L g553 ( 
.A(n_377),
.B(n_218),
.Y(n_553)
);

INVx2_ASAP7_75t_L g554 ( 
.A(n_390),
.Y(n_554)
);

BUFx6f_ASAP7_75t_L g555 ( 
.A(n_438),
.Y(n_555)
);

INVx2_ASAP7_75t_SL g556 ( 
.A(n_396),
.Y(n_556)
);

BUFx3_ASAP7_75t_L g557 ( 
.A(n_377),
.Y(n_557)
);

NOR2xp33_ASAP7_75t_L g558 ( 
.A(n_435),
.B(n_396),
.Y(n_558)
);

NAND2xp5_ASAP7_75t_L g559 ( 
.A(n_377),
.B(n_222),
.Y(n_559)
);

NAND2xp5_ASAP7_75t_SL g560 ( 
.A(n_424),
.B(n_228),
.Y(n_560)
);

NAND2xp5_ASAP7_75t_L g561 ( 
.A(n_377),
.B(n_235),
.Y(n_561)
);

NAND3xp33_ASAP7_75t_SL g562 ( 
.A(n_382),
.B(n_210),
.C(n_182),
.Y(n_562)
);

INVx1_ASAP7_75t_L g563 ( 
.A(n_419),
.Y(n_563)
);

INVx1_ASAP7_75t_L g564 ( 
.A(n_422),
.Y(n_564)
);

INVx1_ASAP7_75t_L g565 ( 
.A(n_422),
.Y(n_565)
);

OR2x6_ASAP7_75t_L g566 ( 
.A(n_418),
.B(n_216),
.Y(n_566)
);

INVx1_ASAP7_75t_L g567 ( 
.A(n_426),
.Y(n_567)
);

INVx1_ASAP7_75t_L g568 ( 
.A(n_426),
.Y(n_568)
);

NAND2xp5_ASAP7_75t_L g569 ( 
.A(n_430),
.B(n_236),
.Y(n_569)
);

INVx1_ASAP7_75t_L g570 ( 
.A(n_430),
.Y(n_570)
);

BUFx6f_ASAP7_75t_SL g571 ( 
.A(n_434),
.Y(n_571)
);

NAND2xp5_ASAP7_75t_SL g572 ( 
.A(n_424),
.B(n_238),
.Y(n_572)
);

NAND2xp5_ASAP7_75t_L g573 ( 
.A(n_431),
.B(n_239),
.Y(n_573)
);

NAND2xp5_ASAP7_75t_L g574 ( 
.A(n_431),
.B(n_240),
.Y(n_574)
);

INVx1_ASAP7_75t_L g575 ( 
.A(n_441),
.Y(n_575)
);

INVx1_ASAP7_75t_L g576 ( 
.A(n_441),
.Y(n_576)
);

NAND3xp33_ASAP7_75t_L g577 ( 
.A(n_418),
.B(n_203),
.C(n_196),
.Y(n_577)
);

NOR2xp33_ASAP7_75t_L g578 ( 
.A(n_424),
.B(n_308),
.Y(n_578)
);

AND2x2_ASAP7_75t_L g579 ( 
.A(n_423),
.B(n_341),
.Y(n_579)
);

BUFx10_ASAP7_75t_L g580 ( 
.A(n_424),
.Y(n_580)
);

BUFx3_ASAP7_75t_L g581 ( 
.A(n_434),
.Y(n_581)
);

INVx3_ASAP7_75t_L g582 ( 
.A(n_392),
.Y(n_582)
);

NAND3xp33_ASAP7_75t_L g583 ( 
.A(n_382),
.B(n_254),
.C(n_226),
.Y(n_583)
);

INVx1_ASAP7_75t_L g584 ( 
.A(n_423),
.Y(n_584)
);

AND2x2_ASAP7_75t_L g585 ( 
.A(n_423),
.B(n_342),
.Y(n_585)
);

CKINVDCx20_ASAP7_75t_R g586 ( 
.A(n_432),
.Y(n_586)
);

AND3x2_ASAP7_75t_L g587 ( 
.A(n_439),
.B(n_157),
.C(n_156),
.Y(n_587)
);

NAND2xp5_ASAP7_75t_SL g588 ( 
.A(n_434),
.B(n_241),
.Y(n_588)
);

INVx8_ASAP7_75t_L g589 ( 
.A(n_500),
.Y(n_589)
);

NAND2xp5_ASAP7_75t_SL g590 ( 
.A(n_448),
.B(n_439),
.Y(n_590)
);

AND2x2_ASAP7_75t_L g591 ( 
.A(n_522),
.B(n_317),
.Y(n_591)
);

INVx2_ASAP7_75t_SL g592 ( 
.A(n_453),
.Y(n_592)
);

INVx2_ASAP7_75t_L g593 ( 
.A(n_448),
.Y(n_593)
);

INVx2_ASAP7_75t_L g594 ( 
.A(n_448),
.Y(n_594)
);

NAND2xp5_ASAP7_75t_SL g595 ( 
.A(n_448),
.B(n_439),
.Y(n_595)
);

NAND2xp5_ASAP7_75t_SL g596 ( 
.A(n_448),
.B(n_439),
.Y(n_596)
);

BUFx6f_ASAP7_75t_L g597 ( 
.A(n_557),
.Y(n_597)
);

AND2x6_ASAP7_75t_SL g598 ( 
.A(n_566),
.B(n_225),
.Y(n_598)
);

NAND2xp5_ASAP7_75t_L g599 ( 
.A(n_515),
.B(n_434),
.Y(n_599)
);

INVx3_ASAP7_75t_L g600 ( 
.A(n_557),
.Y(n_600)
);

NAND2xp5_ASAP7_75t_SL g601 ( 
.A(n_507),
.B(n_434),
.Y(n_601)
);

NAND2xp5_ASAP7_75t_L g602 ( 
.A(n_584),
.B(n_437),
.Y(n_602)
);

NAND2xp5_ASAP7_75t_L g603 ( 
.A(n_584),
.B(n_437),
.Y(n_603)
);

BUFx6f_ASAP7_75t_L g604 ( 
.A(n_581),
.Y(n_604)
);

NAND3xp33_ASAP7_75t_L g605 ( 
.A(n_558),
.B(n_219),
.C(n_217),
.Y(n_605)
);

NOR2xp33_ASAP7_75t_L g606 ( 
.A(n_547),
.B(n_247),
.Y(n_606)
);

NAND2xp5_ASAP7_75t_L g607 ( 
.A(n_473),
.B(n_437),
.Y(n_607)
);

NAND2xp5_ASAP7_75t_SL g608 ( 
.A(n_507),
.B(n_242),
.Y(n_608)
);

AND2x2_ASAP7_75t_L g609 ( 
.A(n_482),
.B(n_320),
.Y(n_609)
);

INVx2_ASAP7_75t_SL g610 ( 
.A(n_556),
.Y(n_610)
);

NAND2xp5_ASAP7_75t_L g611 ( 
.A(n_526),
.B(n_437),
.Y(n_611)
);

OAI22xp33_ASAP7_75t_L g612 ( 
.A1(n_526),
.A2(n_261),
.B1(n_280),
.B2(n_169),
.Y(n_612)
);

INVx2_ASAP7_75t_L g613 ( 
.A(n_445),
.Y(n_613)
);

NOR2xp33_ASAP7_75t_L g614 ( 
.A(n_482),
.B(n_220),
.Y(n_614)
);

NAND2xp33_ASAP7_75t_L g615 ( 
.A(n_481),
.B(n_244),
.Y(n_615)
);

AND2x2_ASAP7_75t_L g616 ( 
.A(n_501),
.B(n_432),
.Y(n_616)
);

O2A1O1Ixp33_ASAP7_75t_L g617 ( 
.A1(n_445),
.A2(n_447),
.B(n_451),
.C(n_446),
.Y(n_617)
);

BUFx12f_ASAP7_75t_L g618 ( 
.A(n_535),
.Y(n_618)
);

AOI22xp33_ASAP7_75t_L g619 ( 
.A1(n_446),
.A2(n_156),
.B1(n_157),
.B2(n_163),
.Y(n_619)
);

NAND2xp5_ASAP7_75t_SL g620 ( 
.A(n_520),
.B(n_246),
.Y(n_620)
);

NAND2xp33_ASAP7_75t_L g621 ( 
.A(n_520),
.B(n_251),
.Y(n_621)
);

NOR2xp33_ASAP7_75t_L g622 ( 
.A(n_463),
.B(n_224),
.Y(n_622)
);

NAND2xp5_ASAP7_75t_SL g623 ( 
.A(n_520),
.B(n_545),
.Y(n_623)
);

NOR2xp33_ASAP7_75t_L g624 ( 
.A(n_489),
.B(n_229),
.Y(n_624)
);

NOR3xp33_ASAP7_75t_L g625 ( 
.A(n_562),
.B(n_237),
.C(n_262),
.Y(n_625)
);

NAND2xp5_ASAP7_75t_L g626 ( 
.A(n_467),
.B(n_503),
.Y(n_626)
);

NAND2xp5_ASAP7_75t_L g627 ( 
.A(n_467),
.B(n_437),
.Y(n_627)
);

INVx1_ASAP7_75t_L g628 ( 
.A(n_579),
.Y(n_628)
);

OAI22xp5_ASAP7_75t_SL g629 ( 
.A1(n_459),
.A2(n_234),
.B1(n_258),
.B2(n_269),
.Y(n_629)
);

INVxp67_ASAP7_75t_L g630 ( 
.A(n_490),
.Y(n_630)
);

BUFx6f_ASAP7_75t_L g631 ( 
.A(n_581),
.Y(n_631)
);

INVx2_ASAP7_75t_L g632 ( 
.A(n_447),
.Y(n_632)
);

NAND2xp5_ASAP7_75t_SL g633 ( 
.A(n_520),
.B(n_253),
.Y(n_633)
);

NAND2xp5_ASAP7_75t_L g634 ( 
.A(n_503),
.B(n_437),
.Y(n_634)
);

INVx1_ASAP7_75t_L g635 ( 
.A(n_579),
.Y(n_635)
);

AOI22xp5_ASAP7_75t_L g636 ( 
.A1(n_523),
.A2(n_260),
.B1(n_264),
.B2(n_266),
.Y(n_636)
);

NAND2xp5_ASAP7_75t_L g637 ( 
.A(n_509),
.B(n_437),
.Y(n_637)
);

NAND2xp5_ASAP7_75t_L g638 ( 
.A(n_509),
.B(n_437),
.Y(n_638)
);

INVx1_ASAP7_75t_L g639 ( 
.A(n_585),
.Y(n_639)
);

NAND2xp5_ASAP7_75t_SL g640 ( 
.A(n_520),
.B(n_271),
.Y(n_640)
);

INVx1_ASAP7_75t_L g641 ( 
.A(n_585),
.Y(n_641)
);

INVx2_ASAP7_75t_L g642 ( 
.A(n_451),
.Y(n_642)
);

NAND2xp5_ASAP7_75t_SL g643 ( 
.A(n_462),
.B(n_273),
.Y(n_643)
);

NAND2xp5_ASAP7_75t_L g644 ( 
.A(n_516),
.B(n_163),
.Y(n_644)
);

INVx1_ASAP7_75t_L g645 ( 
.A(n_516),
.Y(n_645)
);

INVx3_ASAP7_75t_L g646 ( 
.A(n_545),
.Y(n_646)
);

NAND2xp5_ASAP7_75t_L g647 ( 
.A(n_518),
.B(n_169),
.Y(n_647)
);

NAND2xp5_ASAP7_75t_SL g648 ( 
.A(n_545),
.B(n_279),
.Y(n_648)
);

NOR2xp33_ASAP7_75t_L g649 ( 
.A(n_458),
.B(n_270),
.Y(n_649)
);

INVx2_ASAP7_75t_L g650 ( 
.A(n_455),
.Y(n_650)
);

AND2x2_ASAP7_75t_L g651 ( 
.A(n_556),
.B(n_367),
.Y(n_651)
);

AOI22xp33_ASAP7_75t_L g652 ( 
.A1(n_455),
.A2(n_206),
.B1(n_175),
.B2(n_177),
.Y(n_652)
);

INVx2_ASAP7_75t_L g653 ( 
.A(n_456),
.Y(n_653)
);

BUFx3_ASAP7_75t_L g654 ( 
.A(n_458),
.Y(n_654)
);

NAND2xp5_ASAP7_75t_L g655 ( 
.A(n_518),
.B(n_175),
.Y(n_655)
);

AND2x2_ASAP7_75t_L g656 ( 
.A(n_490),
.B(n_370),
.Y(n_656)
);

AND2x4_ASAP7_75t_L g657 ( 
.A(n_542),
.B(n_177),
.Y(n_657)
);

NOR2xp33_ASAP7_75t_L g658 ( 
.A(n_586),
.B(n_277),
.Y(n_658)
);

INVx2_ASAP7_75t_L g659 ( 
.A(n_456),
.Y(n_659)
);

INVx2_ASAP7_75t_L g660 ( 
.A(n_470),
.Y(n_660)
);

A2O1A1Ixp33_ASAP7_75t_L g661 ( 
.A1(n_543),
.A2(n_209),
.B(n_302),
.C(n_294),
.Y(n_661)
);

NOR2xp33_ASAP7_75t_L g662 ( 
.A(n_586),
.B(n_281),
.Y(n_662)
);

INVx1_ASAP7_75t_L g663 ( 
.A(n_521),
.Y(n_663)
);

AND2x2_ASAP7_75t_L g664 ( 
.A(n_454),
.B(n_370),
.Y(n_664)
);

NOR2xp33_ASAP7_75t_L g665 ( 
.A(n_536),
.B(n_283),
.Y(n_665)
);

NAND2xp5_ASAP7_75t_L g666 ( 
.A(n_521),
.B(n_185),
.Y(n_666)
);

AOI22xp33_ASAP7_75t_L g667 ( 
.A1(n_551),
.A2(n_201),
.B1(n_187),
.B2(n_188),
.Y(n_667)
);

AND2x2_ASAP7_75t_L g668 ( 
.A(n_471),
.B(n_375),
.Y(n_668)
);

INVx2_ASAP7_75t_L g669 ( 
.A(n_470),
.Y(n_669)
);

INVx2_ASAP7_75t_SL g670 ( 
.A(n_517),
.Y(n_670)
);

NAND2xp5_ASAP7_75t_SL g671 ( 
.A(n_545),
.B(n_289),
.Y(n_671)
);

OAI22x1_ASAP7_75t_L g672 ( 
.A1(n_577),
.A2(n_293),
.B1(n_295),
.B2(n_297),
.Y(n_672)
);

INVx1_ASAP7_75t_L g673 ( 
.A(n_524),
.Y(n_673)
);

INVx3_ASAP7_75t_L g674 ( 
.A(n_545),
.Y(n_674)
);

OR2x6_ASAP7_75t_L g675 ( 
.A(n_494),
.B(n_500),
.Y(n_675)
);

INVx2_ASAP7_75t_L g676 ( 
.A(n_472),
.Y(n_676)
);

NAND2xp5_ASAP7_75t_L g677 ( 
.A(n_524),
.B(n_185),
.Y(n_677)
);

OAI22xp5_ASAP7_75t_SL g678 ( 
.A1(n_566),
.A2(n_304),
.B1(n_286),
.B2(n_299),
.Y(n_678)
);

O2A1O1Ixp33_ASAP7_75t_L g679 ( 
.A1(n_468),
.A2(n_245),
.B(n_256),
.C(n_259),
.Y(n_679)
);

NAND2xp5_ASAP7_75t_SL g680 ( 
.A(n_555),
.B(n_296),
.Y(n_680)
);

INVx2_ASAP7_75t_L g681 ( 
.A(n_472),
.Y(n_681)
);

NAND2xp5_ASAP7_75t_L g682 ( 
.A(n_525),
.B(n_187),
.Y(n_682)
);

INVx2_ASAP7_75t_L g683 ( 
.A(n_475),
.Y(n_683)
);

INVx2_ASAP7_75t_L g684 ( 
.A(n_475),
.Y(n_684)
);

INVxp67_ASAP7_75t_L g685 ( 
.A(n_486),
.Y(n_685)
);

INVx2_ASAP7_75t_L g686 ( 
.A(n_478),
.Y(n_686)
);

INVx3_ASAP7_75t_L g687 ( 
.A(n_555),
.Y(n_687)
);

AOI22x1_ASAP7_75t_L g688 ( 
.A1(n_525),
.A2(n_188),
.B1(n_199),
.B2(n_201),
.Y(n_688)
);

INVx1_ASAP7_75t_L g689 ( 
.A(n_540),
.Y(n_689)
);

NOR2xp33_ASAP7_75t_L g690 ( 
.A(n_500),
.B(n_305),
.Y(n_690)
);

NAND2xp5_ASAP7_75t_L g691 ( 
.A(n_540),
.B(n_199),
.Y(n_691)
);

INVx1_ASAP7_75t_L g692 ( 
.A(n_563),
.Y(n_692)
);

O2A1O1Ixp33_ASAP7_75t_L g693 ( 
.A1(n_468),
.A2(n_285),
.B(n_245),
.C(n_256),
.Y(n_693)
);

INVx1_ASAP7_75t_L g694 ( 
.A(n_563),
.Y(n_694)
);

OR2x6_ASAP7_75t_L g695 ( 
.A(n_500),
.B(n_259),
.Y(n_695)
);

BUFx12f_ASAP7_75t_L g696 ( 
.A(n_535),
.Y(n_696)
);

INVx2_ASAP7_75t_L g697 ( 
.A(n_478),
.Y(n_697)
);

NAND2xp5_ASAP7_75t_L g698 ( 
.A(n_564),
.B(n_565),
.Y(n_698)
);

NAND2xp5_ASAP7_75t_SL g699 ( 
.A(n_555),
.B(n_298),
.Y(n_699)
);

NAND2xp5_ASAP7_75t_L g700 ( 
.A(n_564),
.B(n_206),
.Y(n_700)
);

BUFx6f_ASAP7_75t_L g701 ( 
.A(n_555),
.Y(n_701)
);

NAND2xp5_ASAP7_75t_L g702 ( 
.A(n_565),
.B(n_209),
.Y(n_702)
);

INVxp67_ASAP7_75t_L g703 ( 
.A(n_578),
.Y(n_703)
);

AOI22xp33_ASAP7_75t_L g704 ( 
.A1(n_567),
.A2(n_570),
.B1(n_568),
.B2(n_576),
.Y(n_704)
);

NAND2xp5_ASAP7_75t_SL g705 ( 
.A(n_555),
.B(n_213),
.Y(n_705)
);

OAI22xp33_ASAP7_75t_L g706 ( 
.A1(n_544),
.A2(n_302),
.B1(n_221),
.B2(n_227),
.Y(n_706)
);

NAND2xp5_ASAP7_75t_L g707 ( 
.A(n_567),
.B(n_213),
.Y(n_707)
);

NOR2xp33_ASAP7_75t_L g708 ( 
.A(n_541),
.B(n_221),
.Y(n_708)
);

NOR2xp33_ASAP7_75t_L g709 ( 
.A(n_569),
.B(n_227),
.Y(n_709)
);

NAND2xp5_ASAP7_75t_L g710 ( 
.A(n_568),
.B(n_233),
.Y(n_710)
);

INVx2_ASAP7_75t_SL g711 ( 
.A(n_491),
.Y(n_711)
);

AOI22xp5_ASAP7_75t_L g712 ( 
.A1(n_571),
.A2(n_233),
.B1(n_252),
.B2(n_257),
.Y(n_712)
);

NAND2xp5_ASAP7_75t_L g713 ( 
.A(n_570),
.B(n_252),
.Y(n_713)
);

INVx1_ASAP7_75t_L g714 ( 
.A(n_575),
.Y(n_714)
);

NAND2xp5_ASAP7_75t_L g715 ( 
.A(n_575),
.B(n_257),
.Y(n_715)
);

NAND2xp5_ASAP7_75t_L g716 ( 
.A(n_576),
.B(n_261),
.Y(n_716)
);

NAND2xp5_ASAP7_75t_L g717 ( 
.A(n_508),
.B(n_280),
.Y(n_717)
);

NOR2xp33_ASAP7_75t_L g718 ( 
.A(n_573),
.B(n_294),
.Y(n_718)
);

INVx2_ASAP7_75t_L g719 ( 
.A(n_484),
.Y(n_719)
);

AOI22xp5_ASAP7_75t_L g720 ( 
.A1(n_571),
.A2(n_436),
.B1(n_429),
.B2(n_428),
.Y(n_720)
);

INVx3_ASAP7_75t_L g721 ( 
.A(n_548),
.Y(n_721)
);

NAND2xp33_ASAP7_75t_SL g722 ( 
.A(n_502),
.B(n_263),
.Y(n_722)
);

NAND2xp33_ASAP7_75t_L g723 ( 
.A(n_553),
.B(n_392),
.Y(n_723)
);

INVx1_ASAP7_75t_L g724 ( 
.A(n_484),
.Y(n_724)
);

NAND2xp5_ASAP7_75t_L g725 ( 
.A(n_537),
.B(n_392),
.Y(n_725)
);

NAND2xp5_ASAP7_75t_L g726 ( 
.A(n_485),
.B(n_392),
.Y(n_726)
);

AOI22xp33_ASAP7_75t_L g727 ( 
.A1(n_548),
.A2(n_413),
.B1(n_407),
.B2(n_284),
.Y(n_727)
);

AND2x2_ASAP7_75t_L g728 ( 
.A(n_449),
.B(n_474),
.Y(n_728)
);

NAND2xp5_ASAP7_75t_L g729 ( 
.A(n_485),
.B(n_436),
.Y(n_729)
);

INVx1_ASAP7_75t_L g730 ( 
.A(n_495),
.Y(n_730)
);

A2O1A1Ixp33_ASAP7_75t_L g731 ( 
.A1(n_495),
.A2(n_499),
.B(n_496),
.C(n_561),
.Y(n_731)
);

AND2x2_ASAP7_75t_L g732 ( 
.A(n_474),
.B(n_375),
.Y(n_732)
);

NAND2xp5_ASAP7_75t_L g733 ( 
.A(n_496),
.B(n_436),
.Y(n_733)
);

NAND2xp5_ASAP7_75t_L g734 ( 
.A(n_499),
.B(n_436),
.Y(n_734)
);

NAND2xp5_ASAP7_75t_L g735 ( 
.A(n_574),
.B(n_429),
.Y(n_735)
);

NAND2xp5_ASAP7_75t_SL g736 ( 
.A(n_559),
.B(n_413),
.Y(n_736)
);

NAND2xp5_ASAP7_75t_SL g737 ( 
.A(n_493),
.B(n_413),
.Y(n_737)
);

AND2x2_ASAP7_75t_L g738 ( 
.A(n_544),
.B(n_346),
.Y(n_738)
);

OR2x2_ASAP7_75t_L g739 ( 
.A(n_544),
.B(n_263),
.Y(n_739)
);

INVx2_ASAP7_75t_L g740 ( 
.A(n_442),
.Y(n_740)
);

NAND2xp5_ASAP7_75t_SL g741 ( 
.A(n_450),
.B(n_413),
.Y(n_741)
);

INVx1_ASAP7_75t_L g742 ( 
.A(n_539),
.Y(n_742)
);

NOR2xp33_ASAP7_75t_L g743 ( 
.A(n_583),
.B(n_275),
.Y(n_743)
);

NAND2xp5_ASAP7_75t_L g744 ( 
.A(n_582),
.B(n_429),
.Y(n_744)
);

NAND2xp5_ASAP7_75t_SL g745 ( 
.A(n_450),
.B(n_413),
.Y(n_745)
);

AND2x2_ASAP7_75t_L g746 ( 
.A(n_544),
.B(n_347),
.Y(n_746)
);

BUFx6f_ASAP7_75t_L g747 ( 
.A(n_587),
.Y(n_747)
);

NAND2xp5_ASAP7_75t_L g748 ( 
.A(n_582),
.B(n_429),
.Y(n_748)
);

NAND2xp5_ASAP7_75t_L g749 ( 
.A(n_582),
.B(n_450),
.Y(n_749)
);

NAND2xp33_ASAP7_75t_L g750 ( 
.A(n_588),
.B(n_413),
.Y(n_750)
);

INVx1_ASAP7_75t_L g751 ( 
.A(n_539),
.Y(n_751)
);

O2A1O1Ixp33_ASAP7_75t_L g752 ( 
.A1(n_546),
.A2(n_275),
.B(n_284),
.C(n_285),
.Y(n_752)
);

INVxp33_ASAP7_75t_L g753 ( 
.A(n_505),
.Y(n_753)
);

INVx1_ASAP7_75t_L g754 ( 
.A(n_549),
.Y(n_754)
);

INVx2_ASAP7_75t_L g755 ( 
.A(n_442),
.Y(n_755)
);

INVx8_ASAP7_75t_L g756 ( 
.A(n_571),
.Y(n_756)
);

AND2x2_ASAP7_75t_L g757 ( 
.A(n_546),
.B(n_342),
.Y(n_757)
);

INVx2_ASAP7_75t_L g758 ( 
.A(n_443),
.Y(n_758)
);

NAND2xp5_ASAP7_75t_SL g759 ( 
.A(n_701),
.B(n_580),
.Y(n_759)
);

NOR2xp33_ASAP7_75t_SL g760 ( 
.A(n_618),
.B(n_528),
.Y(n_760)
);

NAND2xp5_ASAP7_75t_L g761 ( 
.A(n_616),
.B(n_546),
.Y(n_761)
);

INVx1_ASAP7_75t_L g762 ( 
.A(n_653),
.Y(n_762)
);

INVx2_ASAP7_75t_L g763 ( 
.A(n_653),
.Y(n_763)
);

NAND2xp5_ASAP7_75t_L g764 ( 
.A(n_606),
.B(n_546),
.Y(n_764)
);

BUFx6f_ASAP7_75t_L g765 ( 
.A(n_701),
.Y(n_765)
);

BUFx2_ASAP7_75t_L g766 ( 
.A(n_609),
.Y(n_766)
);

AOI22xp33_ASAP7_75t_L g767 ( 
.A1(n_606),
.A2(n_566),
.B1(n_287),
.B2(n_300),
.Y(n_767)
);

INVx2_ASAP7_75t_L g768 ( 
.A(n_659),
.Y(n_768)
);

INVx1_ASAP7_75t_L g769 ( 
.A(n_660),
.Y(n_769)
);

BUFx3_ASAP7_75t_L g770 ( 
.A(n_618),
.Y(n_770)
);

INVx1_ASAP7_75t_L g771 ( 
.A(n_660),
.Y(n_771)
);

INVx1_ASAP7_75t_L g772 ( 
.A(n_669),
.Y(n_772)
);

INVx1_ASAP7_75t_L g773 ( 
.A(n_669),
.Y(n_773)
);

INVx4_ASAP7_75t_L g774 ( 
.A(n_701),
.Y(n_774)
);

INVx5_ASAP7_75t_L g775 ( 
.A(n_701),
.Y(n_775)
);

BUFx12f_ASAP7_75t_L g776 ( 
.A(n_696),
.Y(n_776)
);

NAND2xp5_ASAP7_75t_SL g777 ( 
.A(n_610),
.B(n_580),
.Y(n_777)
);

AOI21xp5_ASAP7_75t_L g778 ( 
.A1(n_590),
.A2(n_488),
.B(n_460),
.Y(n_778)
);

BUFx8_ASAP7_75t_L g779 ( 
.A(n_696),
.Y(n_779)
);

AOI22xp33_ASAP7_75t_L g780 ( 
.A1(n_613),
.A2(n_566),
.B1(n_287),
.B2(n_300),
.Y(n_780)
);

INVx1_ASAP7_75t_L g781 ( 
.A(n_676),
.Y(n_781)
);

BUFx12f_ASAP7_75t_SL g782 ( 
.A(n_695),
.Y(n_782)
);

INVx2_ASAP7_75t_L g783 ( 
.A(n_676),
.Y(n_783)
);

AND2x6_ASAP7_75t_SL g784 ( 
.A(n_658),
.B(n_662),
.Y(n_784)
);

HB1xp67_ASAP7_75t_L g785 ( 
.A(n_630),
.Y(n_785)
);

NAND2xp5_ASAP7_75t_L g786 ( 
.A(n_709),
.B(n_460),
.Y(n_786)
);

AOI22xp5_ASAP7_75t_L g787 ( 
.A1(n_624),
.A2(n_548),
.B1(n_527),
.B2(n_452),
.Y(n_787)
);

INVx2_ASAP7_75t_SL g788 ( 
.A(n_664),
.Y(n_788)
);

AO22x1_ASAP7_75t_L g789 ( 
.A1(n_753),
.A2(n_580),
.B1(n_528),
.B2(n_345),
.Y(n_789)
);

INVx2_ASAP7_75t_L g790 ( 
.A(n_681),
.Y(n_790)
);

AOI22xp33_ASAP7_75t_L g791 ( 
.A1(n_613),
.A2(n_444),
.B1(n_443),
.B2(n_461),
.Y(n_791)
);

NAND2xp5_ASAP7_75t_L g792 ( 
.A(n_709),
.B(n_488),
.Y(n_792)
);

NAND2xp5_ASAP7_75t_L g793 ( 
.A(n_718),
.B(n_488),
.Y(n_793)
);

NAND2xp5_ASAP7_75t_L g794 ( 
.A(n_718),
.B(n_504),
.Y(n_794)
);

BUFx8_ASAP7_75t_L g795 ( 
.A(n_592),
.Y(n_795)
);

INVx2_ASAP7_75t_SL g796 ( 
.A(n_656),
.Y(n_796)
);

AOI22xp5_ASAP7_75t_L g797 ( 
.A1(n_624),
.A2(n_479),
.B1(n_572),
.B2(n_560),
.Y(n_797)
);

INVx2_ASAP7_75t_L g798 ( 
.A(n_681),
.Y(n_798)
);

HB1xp67_ASAP7_75t_L g799 ( 
.A(n_654),
.Y(n_799)
);

NAND2xp33_ASAP7_75t_L g800 ( 
.A(n_597),
.B(n_604),
.Y(n_800)
);

BUFx6f_ASAP7_75t_L g801 ( 
.A(n_597),
.Y(n_801)
);

NAND2xp5_ASAP7_75t_SL g802 ( 
.A(n_732),
.B(n_497),
.Y(n_802)
);

INVx1_ASAP7_75t_L g803 ( 
.A(n_683),
.Y(n_803)
);

AOI22xp5_ASAP7_75t_L g804 ( 
.A1(n_622),
.A2(n_514),
.B1(n_506),
.B2(n_550),
.Y(n_804)
);

INVx1_ASAP7_75t_L g805 ( 
.A(n_683),
.Y(n_805)
);

AOI22xp33_ASAP7_75t_L g806 ( 
.A1(n_632),
.A2(n_444),
.B1(n_487),
.B2(n_457),
.Y(n_806)
);

BUFx6f_ASAP7_75t_L g807 ( 
.A(n_597),
.Y(n_807)
);

NAND3xp33_ASAP7_75t_SL g808 ( 
.A(n_743),
.B(n_345),
.C(n_346),
.Y(n_808)
);

NAND2xp5_ASAP7_75t_SL g809 ( 
.A(n_604),
.B(n_504),
.Y(n_809)
);

NAND2xp5_ASAP7_75t_L g810 ( 
.A(n_626),
.B(n_645),
.Y(n_810)
);

AND2x6_ASAP7_75t_SL g811 ( 
.A(n_658),
.B(n_662),
.Y(n_811)
);

AOI22xp33_ASAP7_75t_L g812 ( 
.A1(n_632),
.A2(n_492),
.B1(n_457),
.B2(n_461),
.Y(n_812)
);

NAND2xp33_ASAP7_75t_L g813 ( 
.A(n_604),
.B(n_504),
.Y(n_813)
);

INVx1_ASAP7_75t_L g814 ( 
.A(n_684),
.Y(n_814)
);

CKINVDCx14_ASAP7_75t_R g815 ( 
.A(n_591),
.Y(n_815)
);

INVxp67_ASAP7_75t_L g816 ( 
.A(n_651),
.Y(n_816)
);

AND2x2_ASAP7_75t_L g817 ( 
.A(n_668),
.B(n_347),
.Y(n_817)
);

CKINVDCx5p33_ASAP7_75t_R g818 ( 
.A(n_685),
.Y(n_818)
);

AND2x2_ASAP7_75t_SL g819 ( 
.A(n_743),
.B(n_476),
.Y(n_819)
);

CKINVDCx5p33_ASAP7_75t_R g820 ( 
.A(n_703),
.Y(n_820)
);

NAND2xp5_ASAP7_75t_L g821 ( 
.A(n_663),
.B(n_506),
.Y(n_821)
);

NAND2xp5_ASAP7_75t_L g822 ( 
.A(n_673),
.B(n_689),
.Y(n_822)
);

INVx2_ASAP7_75t_L g823 ( 
.A(n_684),
.Y(n_823)
);

INVx2_ASAP7_75t_SL g824 ( 
.A(n_738),
.Y(n_824)
);

NAND2xp5_ASAP7_75t_SL g825 ( 
.A(n_604),
.B(n_506),
.Y(n_825)
);

NAND2xp5_ASAP7_75t_SL g826 ( 
.A(n_631),
.B(n_514),
.Y(n_826)
);

AND2x4_ASAP7_75t_L g827 ( 
.A(n_654),
.B(n_514),
.Y(n_827)
);

BUFx3_ASAP7_75t_L g828 ( 
.A(n_670),
.Y(n_828)
);

NAND3xp33_ASAP7_75t_SL g829 ( 
.A(n_665),
.B(n_428),
.C(n_425),
.Y(n_829)
);

INVx1_ASAP7_75t_L g830 ( 
.A(n_686),
.Y(n_830)
);

INVx1_ASAP7_75t_L g831 ( 
.A(n_686),
.Y(n_831)
);

BUFx3_ASAP7_75t_L g832 ( 
.A(n_711),
.Y(n_832)
);

AND2x2_ASAP7_75t_L g833 ( 
.A(n_728),
.B(n_425),
.Y(n_833)
);

NAND2xp5_ASAP7_75t_L g834 ( 
.A(n_692),
.B(n_530),
.Y(n_834)
);

NAND2xp5_ASAP7_75t_L g835 ( 
.A(n_694),
.B(n_530),
.Y(n_835)
);

INVx2_ASAP7_75t_L g836 ( 
.A(n_697),
.Y(n_836)
);

NOR2xp33_ASAP7_75t_SL g837 ( 
.A(n_756),
.B(n_549),
.Y(n_837)
);

NOR2xp33_ASAP7_75t_L g838 ( 
.A(n_622),
.B(n_476),
.Y(n_838)
);

NAND2xp5_ASAP7_75t_L g839 ( 
.A(n_714),
.B(n_530),
.Y(n_839)
);

INVx1_ASAP7_75t_L g840 ( 
.A(n_697),
.Y(n_840)
);

INVx1_ASAP7_75t_L g841 ( 
.A(n_719),
.Y(n_841)
);

NAND2xp5_ASAP7_75t_L g842 ( 
.A(n_724),
.B(n_550),
.Y(n_842)
);

INVx2_ASAP7_75t_SL g843 ( 
.A(n_746),
.Y(n_843)
);

NAND2x1p5_ASAP7_75t_L g844 ( 
.A(n_721),
.B(n_550),
.Y(n_844)
);

NAND2xp5_ASAP7_75t_L g845 ( 
.A(n_730),
.B(n_552),
.Y(n_845)
);

NAND2x1p5_ASAP7_75t_L g846 ( 
.A(n_721),
.B(n_476),
.Y(n_846)
);

NAND2xp5_ASAP7_75t_SL g847 ( 
.A(n_631),
.B(n_552),
.Y(n_847)
);

NAND2x1p5_ASAP7_75t_L g848 ( 
.A(n_600),
.B(n_483),
.Y(n_848)
);

CKINVDCx5p33_ASAP7_75t_R g849 ( 
.A(n_598),
.Y(n_849)
);

NAND2xp5_ASAP7_75t_L g850 ( 
.A(n_599),
.B(n_554),
.Y(n_850)
);

INVx1_ASAP7_75t_L g851 ( 
.A(n_719),
.Y(n_851)
);

NOR2x1p5_ASAP7_75t_L g852 ( 
.A(n_747),
.B(n_554),
.Y(n_852)
);

OR2x6_ASAP7_75t_L g853 ( 
.A(n_756),
.B(n_425),
.Y(n_853)
);

NAND2xp5_ASAP7_75t_SL g854 ( 
.A(n_631),
.B(n_483),
.Y(n_854)
);

AND2x4_ASAP7_75t_L g855 ( 
.A(n_628),
.B(n_512),
.Y(n_855)
);

BUFx6f_ASAP7_75t_L g856 ( 
.A(n_593),
.Y(n_856)
);

INVx5_ASAP7_75t_L g857 ( 
.A(n_646),
.Y(n_857)
);

AOI22xp33_ASAP7_75t_L g858 ( 
.A1(n_642),
.A2(n_487),
.B1(n_464),
.B2(n_465),
.Y(n_858)
);

AOI22xp5_ASAP7_75t_L g859 ( 
.A1(n_601),
.A2(n_512),
.B1(n_532),
.B2(n_465),
.Y(n_859)
);

INVx2_ASAP7_75t_L g860 ( 
.A(n_740),
.Y(n_860)
);

NAND2xp5_ASAP7_75t_L g861 ( 
.A(n_698),
.B(n_464),
.Y(n_861)
);

AND3x1_ASAP7_75t_L g862 ( 
.A(n_625),
.B(n_428),
.C(n_498),
.Y(n_862)
);

INVx1_ASAP7_75t_L g863 ( 
.A(n_635),
.Y(n_863)
);

HB1xp67_ASAP7_75t_SL g864 ( 
.A(n_690),
.Y(n_864)
);

INVx2_ASAP7_75t_L g865 ( 
.A(n_740),
.Y(n_865)
);

INVx2_ASAP7_75t_L g866 ( 
.A(n_755),
.Y(n_866)
);

AND2x6_ASAP7_75t_SL g867 ( 
.A(n_690),
.B(n_0),
.Y(n_867)
);

INVx4_ASAP7_75t_L g868 ( 
.A(n_756),
.Y(n_868)
);

BUFx6f_ASAP7_75t_L g869 ( 
.A(n_593),
.Y(n_869)
);

AND3x1_ASAP7_75t_L g870 ( 
.A(n_649),
.B(n_428),
.C(n_498),
.Y(n_870)
);

INVx1_ASAP7_75t_L g871 ( 
.A(n_639),
.Y(n_871)
);

BUFx6f_ASAP7_75t_L g872 ( 
.A(n_594),
.Y(n_872)
);

INVx3_ASAP7_75t_L g873 ( 
.A(n_600),
.Y(n_873)
);

NAND2xp5_ASAP7_75t_L g874 ( 
.A(n_704),
.B(n_492),
.Y(n_874)
);

NAND2xp5_ASAP7_75t_L g875 ( 
.A(n_601),
.B(n_510),
.Y(n_875)
);

NAND3xp33_ASAP7_75t_SL g876 ( 
.A(n_665),
.B(n_511),
.C(n_466),
.Y(n_876)
);

A2O1A1Ixp33_ASAP7_75t_L g877 ( 
.A1(n_708),
.A2(n_731),
.B(n_617),
.C(n_614),
.Y(n_877)
);

INVxp67_ASAP7_75t_L g878 ( 
.A(n_649),
.Y(n_878)
);

AOI22xp5_ASAP7_75t_L g879 ( 
.A1(n_641),
.A2(n_532),
.B1(n_466),
.B2(n_469),
.Y(n_879)
);

NAND2xp5_ASAP7_75t_SL g880 ( 
.A(n_708),
.B(n_532),
.Y(n_880)
);

CKINVDCx5p33_ASAP7_75t_R g881 ( 
.A(n_675),
.Y(n_881)
);

INVx2_ASAP7_75t_L g882 ( 
.A(n_755),
.Y(n_882)
);

A2O1A1Ixp33_ASAP7_75t_L g883 ( 
.A1(n_717),
.A2(n_510),
.B(n_469),
.C(n_477),
.Y(n_883)
);

AND2x2_ASAP7_75t_L g884 ( 
.A(n_757),
.B(n_513),
.Y(n_884)
);

AND2x4_ASAP7_75t_L g885 ( 
.A(n_695),
.B(n_70),
.Y(n_885)
);

INVx1_ASAP7_75t_L g886 ( 
.A(n_758),
.Y(n_886)
);

NAND2xp5_ASAP7_75t_SL g887 ( 
.A(n_594),
.B(n_511),
.Y(n_887)
);

NAND2xp5_ASAP7_75t_SL g888 ( 
.A(n_642),
.B(n_480),
.Y(n_888)
);

AND3x2_ASAP7_75t_SL g889 ( 
.A(n_678),
.B(n_0),
.C(n_2),
.Y(n_889)
);

INVx2_ASAP7_75t_L g890 ( 
.A(n_758),
.Y(n_890)
);

INVx1_ASAP7_75t_L g891 ( 
.A(n_742),
.Y(n_891)
);

INVx1_ASAP7_75t_L g892 ( 
.A(n_751),
.Y(n_892)
);

INVxp67_ASAP7_75t_L g893 ( 
.A(n_739),
.Y(n_893)
);

NOR2xp33_ASAP7_75t_R g894 ( 
.A(n_722),
.B(n_60),
.Y(n_894)
);

INVx1_ASAP7_75t_L g895 ( 
.A(n_754),
.Y(n_895)
);

NAND2xp5_ASAP7_75t_L g896 ( 
.A(n_650),
.B(n_480),
.Y(n_896)
);

NAND2xp5_ASAP7_75t_L g897 ( 
.A(n_650),
.B(n_513),
.Y(n_897)
);

AOI22xp33_ASAP7_75t_L g898 ( 
.A1(n_619),
.A2(n_477),
.B1(n_519),
.B2(n_529),
.Y(n_898)
);

INVx2_ASAP7_75t_L g899 ( 
.A(n_611),
.Y(n_899)
);

INVx2_ASAP7_75t_SL g900 ( 
.A(n_657),
.Y(n_900)
);

AOI22xp5_ASAP7_75t_L g901 ( 
.A1(n_620),
.A2(n_519),
.B1(n_529),
.B2(n_533),
.Y(n_901)
);

INVx2_ASAP7_75t_L g902 ( 
.A(n_726),
.Y(n_902)
);

INVx1_ASAP7_75t_L g903 ( 
.A(n_627),
.Y(n_903)
);

OR2x6_ASAP7_75t_L g904 ( 
.A(n_589),
.B(n_538),
.Y(n_904)
);

NAND2xp5_ASAP7_75t_SL g905 ( 
.A(n_607),
.B(n_538),
.Y(n_905)
);

AND2x6_ASAP7_75t_SL g906 ( 
.A(n_675),
.B(n_2),
.Y(n_906)
);

BUFx6f_ASAP7_75t_L g907 ( 
.A(n_646),
.Y(n_907)
);

AND3x1_ASAP7_75t_SL g908 ( 
.A(n_629),
.B(n_3),
.C(n_5),
.Y(n_908)
);

INVx1_ASAP7_75t_L g909 ( 
.A(n_729),
.Y(n_909)
);

AND2x4_ASAP7_75t_L g910 ( 
.A(n_695),
.B(n_657),
.Y(n_910)
);

INVx2_ASAP7_75t_L g911 ( 
.A(n_602),
.Y(n_911)
);

BUFx12f_ASAP7_75t_L g912 ( 
.A(n_747),
.Y(n_912)
);

AOI22xp5_ASAP7_75t_L g913 ( 
.A1(n_620),
.A2(n_534),
.B1(n_533),
.B2(n_531),
.Y(n_913)
);

NAND2xp5_ASAP7_75t_L g914 ( 
.A(n_652),
.B(n_534),
.Y(n_914)
);

INVx2_ASAP7_75t_L g915 ( 
.A(n_603),
.Y(n_915)
);

AOI21xp5_ASAP7_75t_L g916 ( 
.A1(n_590),
.A2(n_531),
.B(n_390),
.Y(n_916)
);

INVx1_ASAP7_75t_L g917 ( 
.A(n_733),
.Y(n_917)
);

NOR2xp33_ASAP7_75t_L g918 ( 
.A(n_608),
.B(n_3),
.Y(n_918)
);

INVx1_ASAP7_75t_L g919 ( 
.A(n_734),
.Y(n_919)
);

INVx2_ASAP7_75t_L g920 ( 
.A(n_749),
.Y(n_920)
);

INVx3_ASAP7_75t_L g921 ( 
.A(n_674),
.Y(n_921)
);

BUFx6f_ASAP7_75t_L g922 ( 
.A(n_674),
.Y(n_922)
);

BUFx4f_ASAP7_75t_L g923 ( 
.A(n_589),
.Y(n_923)
);

NAND2xp5_ASAP7_75t_L g924 ( 
.A(n_595),
.B(n_413),
.Y(n_924)
);

NOR2xp33_ASAP7_75t_L g925 ( 
.A(n_608),
.B(n_9),
.Y(n_925)
);

INVx2_ASAP7_75t_L g926 ( 
.A(n_596),
.Y(n_926)
);

INVx4_ASAP7_75t_L g927 ( 
.A(n_589),
.Y(n_927)
);

INVx4_ASAP7_75t_L g928 ( 
.A(n_687),
.Y(n_928)
);

INVx1_ASAP7_75t_L g929 ( 
.A(n_634),
.Y(n_929)
);

NAND2xp5_ASAP7_75t_L g930 ( 
.A(n_657),
.B(n_687),
.Y(n_930)
);

NAND2xp5_ASAP7_75t_L g931 ( 
.A(n_735),
.B(n_413),
.Y(n_931)
);

INVx1_ASAP7_75t_L g932 ( 
.A(n_637),
.Y(n_932)
);

NOR3xp33_ASAP7_75t_SL g933 ( 
.A(n_706),
.B(n_15),
.C(n_17),
.Y(n_933)
);

NAND2xp5_ASAP7_75t_L g934 ( 
.A(n_623),
.B(n_407),
.Y(n_934)
);

INVx2_ASAP7_75t_L g935 ( 
.A(n_744),
.Y(n_935)
);

NAND2xp5_ASAP7_75t_L g936 ( 
.A(n_623),
.B(n_407),
.Y(n_936)
);

INVx1_ASAP7_75t_L g937 ( 
.A(n_638),
.Y(n_937)
);

NOR2xp33_ASAP7_75t_R g938 ( 
.A(n_615),
.B(n_142),
.Y(n_938)
);

INVx2_ASAP7_75t_L g939 ( 
.A(n_748),
.Y(n_939)
);

BUFx4f_ASAP7_75t_SL g940 ( 
.A(n_747),
.Y(n_940)
);

OAI22xp5_ASAP7_75t_L g941 ( 
.A1(n_767),
.A2(n_705),
.B1(n_605),
.B2(n_675),
.Y(n_941)
);

INVx3_ASAP7_75t_SL g942 ( 
.A(n_820),
.Y(n_942)
);

AOI21xp5_ASAP7_75t_L g943 ( 
.A1(n_775),
.A2(n_621),
.B(n_725),
.Y(n_943)
);

CKINVDCx5p33_ASAP7_75t_R g944 ( 
.A(n_818),
.Y(n_944)
);

INVx1_ASAP7_75t_L g945 ( 
.A(n_762),
.Y(n_945)
);

HB1xp67_ASAP7_75t_L g946 ( 
.A(n_785),
.Y(n_946)
);

AND2x2_ASAP7_75t_L g947 ( 
.A(n_788),
.B(n_672),
.Y(n_947)
);

NAND3xp33_ASAP7_75t_L g948 ( 
.A(n_767),
.B(n_636),
.C(n_643),
.Y(n_948)
);

NAND2xp5_ASAP7_75t_L g949 ( 
.A(n_903),
.B(n_644),
.Y(n_949)
);

AOI21xp5_ASAP7_75t_L g950 ( 
.A1(n_775),
.A2(n_705),
.B(n_723),
.Y(n_950)
);

AOI21xp5_ASAP7_75t_L g951 ( 
.A1(n_850),
.A2(n_699),
.B(n_633),
.Y(n_951)
);

O2A1O1Ixp5_ASAP7_75t_SL g952 ( 
.A1(n_878),
.A2(n_671),
.B(n_633),
.C(n_680),
.Y(n_952)
);

A2O1A1Ixp33_ASAP7_75t_SL g953 ( 
.A1(n_838),
.A2(n_679),
.B(n_693),
.C(n_647),
.Y(n_953)
);

NAND2xp5_ASAP7_75t_L g954 ( 
.A(n_816),
.B(n_655),
.Y(n_954)
);

O2A1O1Ixp5_ASAP7_75t_L g955 ( 
.A1(n_838),
.A2(n_648),
.B(n_680),
.C(n_699),
.Y(n_955)
);

AOI21xp5_ASAP7_75t_L g956 ( 
.A1(n_800),
.A2(n_931),
.B(n_880),
.Y(n_956)
);

INVx1_ASAP7_75t_L g957 ( 
.A(n_769),
.Y(n_957)
);

INVx1_ASAP7_75t_SL g958 ( 
.A(n_785),
.Y(n_958)
);

O2A1O1Ixp33_ASAP7_75t_L g959 ( 
.A1(n_764),
.A2(n_612),
.B(n_752),
.C(n_702),
.Y(n_959)
);

INVx5_ASAP7_75t_L g960 ( 
.A(n_765),
.Y(n_960)
);

NAND2x1p5_ASAP7_75t_L g961 ( 
.A(n_774),
.B(n_737),
.Y(n_961)
);

OAI21x1_ASAP7_75t_L g962 ( 
.A1(n_778),
.A2(n_736),
.B(n_745),
.Y(n_962)
);

INVx2_ASAP7_75t_L g963 ( 
.A(n_763),
.Y(n_963)
);

NOR2xp33_ASAP7_75t_R g964 ( 
.A(n_815),
.B(n_750),
.Y(n_964)
);

NAND2xp5_ASAP7_75t_L g965 ( 
.A(n_816),
.B(n_691),
.Y(n_965)
);

AOI21xp5_ASAP7_75t_L g966 ( 
.A1(n_854),
.A2(n_671),
.B(n_648),
.Y(n_966)
);

AND2x2_ASAP7_75t_L g967 ( 
.A(n_796),
.B(n_712),
.Y(n_967)
);

AOI21xp5_ASAP7_75t_L g968 ( 
.A1(n_854),
.A2(n_640),
.B(n_736),
.Y(n_968)
);

INVx5_ASAP7_75t_L g969 ( 
.A(n_765),
.Y(n_969)
);

INVx2_ASAP7_75t_L g970 ( 
.A(n_768),
.Y(n_970)
);

INVx3_ASAP7_75t_L g971 ( 
.A(n_801),
.Y(n_971)
);

NAND2xp5_ASAP7_75t_SL g972 ( 
.A(n_797),
.B(n_727),
.Y(n_972)
);

INVx2_ASAP7_75t_L g973 ( 
.A(n_783),
.Y(n_973)
);

NOR2xp33_ASAP7_75t_L g974 ( 
.A(n_761),
.B(n_640),
.Y(n_974)
);

AOI22xp5_ASAP7_75t_L g975 ( 
.A1(n_824),
.A2(n_720),
.B1(n_666),
.B2(n_700),
.Y(n_975)
);

NOR2xp33_ASAP7_75t_L g976 ( 
.A(n_766),
.B(n_710),
.Y(n_976)
);

INVx2_ASAP7_75t_L g977 ( 
.A(n_790),
.Y(n_977)
);

O2A1O1Ixp33_ASAP7_75t_L g978 ( 
.A1(n_918),
.A2(n_707),
.B(n_677),
.C(n_716),
.Y(n_978)
);

INVx3_ASAP7_75t_L g979 ( 
.A(n_801),
.Y(n_979)
);

AOI21xp5_ASAP7_75t_L g980 ( 
.A1(n_848),
.A2(n_861),
.B(n_930),
.Y(n_980)
);

OAI22xp5_ASAP7_75t_L g981 ( 
.A1(n_780),
.A2(n_667),
.B1(n_715),
.B2(n_713),
.Y(n_981)
);

A2O1A1Ixp33_ASAP7_75t_L g982 ( 
.A1(n_918),
.A2(n_925),
.B(n_877),
.C(n_787),
.Y(n_982)
);

A2O1A1Ixp33_ASAP7_75t_L g983 ( 
.A1(n_925),
.A2(n_682),
.B(n_745),
.C(n_741),
.Y(n_983)
);

CKINVDCx5p33_ASAP7_75t_R g984 ( 
.A(n_776),
.Y(n_984)
);

INVx2_ASAP7_75t_L g985 ( 
.A(n_798),
.Y(n_985)
);

INVx1_ASAP7_75t_L g986 ( 
.A(n_771),
.Y(n_986)
);

BUFx6f_ASAP7_75t_L g987 ( 
.A(n_801),
.Y(n_987)
);

NAND2xp5_ASAP7_75t_L g988 ( 
.A(n_810),
.B(n_741),
.Y(n_988)
);

INVx2_ASAP7_75t_L g989 ( 
.A(n_823),
.Y(n_989)
);

HB1xp67_ASAP7_75t_L g990 ( 
.A(n_799),
.Y(n_990)
);

AOI33xp33_ASAP7_75t_L g991 ( 
.A1(n_863),
.A2(n_421),
.A3(n_409),
.B1(n_688),
.B2(n_661),
.B3(n_28),
.Y(n_991)
);

A2O1A1Ixp33_ASAP7_75t_L g992 ( 
.A1(n_900),
.A2(n_421),
.B(n_409),
.C(n_407),
.Y(n_992)
);

NAND2xp5_ASAP7_75t_L g993 ( 
.A(n_833),
.B(n_421),
.Y(n_993)
);

NOR2xp33_ASAP7_75t_L g994 ( 
.A(n_893),
.B(n_15),
.Y(n_994)
);

BUFx6f_ASAP7_75t_L g995 ( 
.A(n_801),
.Y(n_995)
);

AOI21x1_ASAP7_75t_L g996 ( 
.A1(n_905),
.A2(n_421),
.B(n_409),
.Y(n_996)
);

AND2x4_ASAP7_75t_L g997 ( 
.A(n_927),
.B(n_108),
.Y(n_997)
);

INVx1_ASAP7_75t_L g998 ( 
.A(n_772),
.Y(n_998)
);

O2A1O1Ixp33_ASAP7_75t_L g999 ( 
.A1(n_802),
.A2(n_409),
.B(n_25),
.C(n_26),
.Y(n_999)
);

CKINVDCx5p33_ASAP7_75t_R g1000 ( 
.A(n_779),
.Y(n_1000)
);

INVx1_ASAP7_75t_L g1001 ( 
.A(n_773),
.Y(n_1001)
);

NAND2xp5_ASAP7_75t_SL g1002 ( 
.A(n_910),
.B(n_843),
.Y(n_1002)
);

NAND2xp5_ASAP7_75t_L g1003 ( 
.A(n_817),
.B(n_407),
.Y(n_1003)
);

AOI22xp33_ASAP7_75t_L g1004 ( 
.A1(n_884),
.A2(n_407),
.B1(n_25),
.B2(n_29),
.Y(n_1004)
);

OAI22xp5_ASAP7_75t_L g1005 ( 
.A1(n_780),
.A2(n_407),
.B1(n_31),
.B2(n_33),
.Y(n_1005)
);

AOI21xp5_ASAP7_75t_L g1006 ( 
.A1(n_848),
.A2(n_407),
.B(n_140),
.Y(n_1006)
);

INVx1_ASAP7_75t_L g1007 ( 
.A(n_781),
.Y(n_1007)
);

AOI21xp5_ASAP7_75t_L g1008 ( 
.A1(n_813),
.A2(n_132),
.B(n_128),
.Y(n_1008)
);

NAND2xp5_ASAP7_75t_L g1009 ( 
.A(n_909),
.B(n_120),
.Y(n_1009)
);

HB1xp67_ASAP7_75t_L g1010 ( 
.A(n_799),
.Y(n_1010)
);

O2A1O1Ixp33_ASAP7_75t_L g1011 ( 
.A1(n_893),
.A2(n_23),
.B(n_34),
.C(n_35),
.Y(n_1011)
);

O2A1O1Ixp33_ASAP7_75t_L g1012 ( 
.A1(n_822),
.A2(n_35),
.B(n_36),
.C(n_37),
.Y(n_1012)
);

NAND2xp5_ASAP7_75t_L g1013 ( 
.A(n_917),
.B(n_119),
.Y(n_1013)
);

BUFx2_ASAP7_75t_SL g1014 ( 
.A(n_868),
.Y(n_1014)
);

A2O1A1Ixp33_ASAP7_75t_L g1015 ( 
.A1(n_926),
.A2(n_919),
.B(n_819),
.C(n_871),
.Y(n_1015)
);

HB1xp67_ASAP7_75t_L g1016 ( 
.A(n_910),
.Y(n_1016)
);

INVx4_ASAP7_75t_L g1017 ( 
.A(n_807),
.Y(n_1017)
);

INVx2_ASAP7_75t_L g1018 ( 
.A(n_836),
.Y(n_1018)
);

NAND2xp5_ASAP7_75t_SL g1019 ( 
.A(n_819),
.B(n_99),
.Y(n_1019)
);

INVx2_ASAP7_75t_L g1020 ( 
.A(n_860),
.Y(n_1020)
);

AND2x2_ASAP7_75t_L g1021 ( 
.A(n_885),
.B(n_832),
.Y(n_1021)
);

NAND2xp5_ASAP7_75t_SL g1022 ( 
.A(n_855),
.B(n_90),
.Y(n_1022)
);

NOR2xp33_ASAP7_75t_L g1023 ( 
.A(n_784),
.B(n_39),
.Y(n_1023)
);

NAND2xp5_ASAP7_75t_SL g1024 ( 
.A(n_855),
.B(n_89),
.Y(n_1024)
);

A2O1A1Ixp33_ASAP7_75t_L g1025 ( 
.A1(n_911),
.A2(n_40),
.B(n_42),
.C(n_43),
.Y(n_1025)
);

NOR2xp33_ASAP7_75t_L g1026 ( 
.A(n_811),
.B(n_42),
.Y(n_1026)
);

NOR3xp33_ASAP7_75t_SL g1027 ( 
.A(n_849),
.B(n_43),
.C(n_44),
.Y(n_1027)
);

AOI21xp5_ASAP7_75t_L g1028 ( 
.A1(n_786),
.A2(n_51),
.B(n_74),
.Y(n_1028)
);

INVx2_ASAP7_75t_L g1029 ( 
.A(n_865),
.Y(n_1029)
);

NAND2xp5_ASAP7_75t_SL g1030 ( 
.A(n_807),
.B(n_827),
.Y(n_1030)
);

AOI21xp5_ASAP7_75t_L g1031 ( 
.A1(n_792),
.A2(n_73),
.B(n_78),
.Y(n_1031)
);

INVx8_ASAP7_75t_L g1032 ( 
.A(n_904),
.Y(n_1032)
);

OAI22xp5_ASAP7_75t_L g1033 ( 
.A1(n_864),
.A2(n_45),
.B1(n_47),
.B2(n_48),
.Y(n_1033)
);

AOI21xp5_ASAP7_75t_L g1034 ( 
.A1(n_793),
.A2(n_47),
.B(n_50),
.Y(n_1034)
);

INVx2_ASAP7_75t_L g1035 ( 
.A(n_866),
.Y(n_1035)
);

NAND2xp5_ASAP7_75t_L g1036 ( 
.A(n_915),
.B(n_899),
.Y(n_1036)
);

AOI21xp5_ASAP7_75t_L g1037 ( 
.A1(n_794),
.A2(n_924),
.B(n_905),
.Y(n_1037)
);

AND2x4_ASAP7_75t_L g1038 ( 
.A(n_927),
.B(n_868),
.Y(n_1038)
);

NAND2xp5_ASAP7_75t_L g1039 ( 
.A(n_929),
.B(n_932),
.Y(n_1039)
);

BUFx2_ASAP7_75t_L g1040 ( 
.A(n_912),
.Y(n_1040)
);

OAI22x1_ASAP7_75t_L g1041 ( 
.A1(n_881),
.A2(n_889),
.B1(n_852),
.B2(n_885),
.Y(n_1041)
);

INVxp67_ASAP7_75t_L g1042 ( 
.A(n_795),
.Y(n_1042)
);

CKINVDCx20_ASAP7_75t_R g1043 ( 
.A(n_779),
.Y(n_1043)
);

NOR2xp33_ASAP7_75t_L g1044 ( 
.A(n_864),
.B(n_940),
.Y(n_1044)
);

AOI21xp5_ASAP7_75t_L g1045 ( 
.A1(n_914),
.A2(n_874),
.B(n_825),
.Y(n_1045)
);

AO21x1_ASAP7_75t_L g1046 ( 
.A1(n_759),
.A2(n_937),
.B(n_830),
.Y(n_1046)
);

INVx1_ASAP7_75t_L g1047 ( 
.A(n_803),
.Y(n_1047)
);

HB1xp67_ASAP7_75t_L g1048 ( 
.A(n_795),
.Y(n_1048)
);

AOI21x1_ASAP7_75t_L g1049 ( 
.A1(n_934),
.A2(n_936),
.B(n_825),
.Y(n_1049)
);

AOI21xp5_ASAP7_75t_L g1050 ( 
.A1(n_809),
.A2(n_897),
.B(n_896),
.Y(n_1050)
);

NOR2xp33_ASAP7_75t_L g1051 ( 
.A(n_940),
.B(n_828),
.Y(n_1051)
);

AND2x4_ASAP7_75t_L g1052 ( 
.A(n_904),
.B(n_827),
.Y(n_1052)
);

CKINVDCx5p33_ASAP7_75t_R g1053 ( 
.A(n_770),
.Y(n_1053)
);

INVxp67_ASAP7_75t_SL g1054 ( 
.A(n_765),
.Y(n_1054)
);

HB1xp67_ASAP7_75t_L g1055 ( 
.A(n_782),
.Y(n_1055)
);

A2O1A1Ixp33_ASAP7_75t_L g1056 ( 
.A1(n_805),
.A2(n_814),
.B(n_831),
.C(n_840),
.Y(n_1056)
);

CKINVDCx5p33_ASAP7_75t_R g1057 ( 
.A(n_923),
.Y(n_1057)
);

NAND2xp5_ASAP7_75t_L g1058 ( 
.A(n_902),
.B(n_935),
.Y(n_1058)
);

O2A1O1Ixp33_ASAP7_75t_L g1059 ( 
.A1(n_808),
.A2(n_933),
.B(n_777),
.C(n_891),
.Y(n_1059)
);

NOR2xp33_ASAP7_75t_L g1060 ( 
.A(n_789),
.B(n_856),
.Y(n_1060)
);

AOI21x1_ASAP7_75t_L g1061 ( 
.A1(n_809),
.A2(n_847),
.B(n_888),
.Y(n_1061)
);

OAI22xp5_ASAP7_75t_L g1062 ( 
.A1(n_841),
.A2(n_851),
.B1(n_933),
.B2(n_791),
.Y(n_1062)
);

NAND3xp33_ASAP7_75t_L g1063 ( 
.A(n_862),
.B(n_760),
.C(n_892),
.Y(n_1063)
);

OAI22xp5_ASAP7_75t_L g1064 ( 
.A1(n_791),
.A2(n_806),
.B1(n_858),
.B2(n_812),
.Y(n_1064)
);

AOI21xp5_ASAP7_75t_L g1065 ( 
.A1(n_875),
.A2(n_778),
.B(n_826),
.Y(n_1065)
);

OAI21x1_ASAP7_75t_L g1066 ( 
.A1(n_916),
.A2(n_887),
.B(n_888),
.Y(n_1066)
);

AOI21xp5_ASAP7_75t_L g1067 ( 
.A1(n_887),
.A2(n_857),
.B(n_920),
.Y(n_1067)
);

AOI21xp5_ASAP7_75t_L g1068 ( 
.A1(n_857),
.A2(n_939),
.B(n_774),
.Y(n_1068)
);

AOI21xp5_ASAP7_75t_L g1069 ( 
.A1(n_857),
.A2(n_928),
.B(n_834),
.Y(n_1069)
);

NAND2xp5_ASAP7_75t_L g1070 ( 
.A(n_856),
.B(n_869),
.Y(n_1070)
);

OAI21xp5_ASAP7_75t_L g1071 ( 
.A1(n_916),
.A2(n_883),
.B(n_829),
.Y(n_1071)
);

INVx5_ASAP7_75t_L g1072 ( 
.A(n_765),
.Y(n_1072)
);

AOI21xp5_ASAP7_75t_L g1073 ( 
.A1(n_857),
.A2(n_928),
.B(n_842),
.Y(n_1073)
);

AND2x4_ASAP7_75t_L g1074 ( 
.A(n_904),
.B(n_853),
.Y(n_1074)
);

A2O1A1Ixp33_ASAP7_75t_L g1075 ( 
.A1(n_895),
.A2(n_804),
.B(n_873),
.C(n_845),
.Y(n_1075)
);

O2A1O1Ixp33_ASAP7_75t_L g1076 ( 
.A1(n_808),
.A2(n_829),
.B(n_835),
.C(n_821),
.Y(n_1076)
);

NAND3xp33_ASAP7_75t_SL g1077 ( 
.A(n_938),
.B(n_894),
.C(n_837),
.Y(n_1077)
);

NAND2xp5_ASAP7_75t_L g1078 ( 
.A(n_856),
.B(n_869),
.Y(n_1078)
);

NAND2xp5_ASAP7_75t_L g1079 ( 
.A(n_1039),
.B(n_882),
.Y(n_1079)
);

OAI21x1_ASAP7_75t_SL g1080 ( 
.A1(n_1046),
.A2(n_839),
.B(n_879),
.Y(n_1080)
);

AO31x2_ASAP7_75t_L g1081 ( 
.A1(n_982),
.A2(n_886),
.A3(n_890),
.B(n_870),
.Y(n_1081)
);

NOR2xp67_ASAP7_75t_L g1082 ( 
.A(n_944),
.B(n_876),
.Y(n_1082)
);

AND2x4_ASAP7_75t_L g1083 ( 
.A(n_1038),
.B(n_853),
.Y(n_1083)
);

AO31x2_ASAP7_75t_L g1084 ( 
.A1(n_1015),
.A2(n_876),
.A3(n_901),
.B(n_913),
.Y(n_1084)
);

NAND2xp5_ASAP7_75t_L g1085 ( 
.A(n_976),
.B(n_872),
.Y(n_1085)
);

INVxp67_ASAP7_75t_SL g1086 ( 
.A(n_946),
.Y(n_1086)
);

NAND3xp33_ASAP7_75t_L g1087 ( 
.A(n_948),
.B(n_853),
.C(n_898),
.Y(n_1087)
);

A2O1A1Ixp33_ASAP7_75t_L g1088 ( 
.A1(n_974),
.A2(n_923),
.B(n_859),
.C(n_921),
.Y(n_1088)
);

OAI21x1_ASAP7_75t_L g1089 ( 
.A1(n_996),
.A2(n_844),
.B(n_806),
.Y(n_1089)
);

AOI21xp5_ASAP7_75t_L g1090 ( 
.A1(n_951),
.A2(n_846),
.B(n_921),
.Y(n_1090)
);

OAI21xp5_ASAP7_75t_L g1091 ( 
.A1(n_955),
.A2(n_898),
.B(n_812),
.Y(n_1091)
);

BUFx6f_ASAP7_75t_L g1092 ( 
.A(n_987),
.Y(n_1092)
);

NAND2x1p5_ASAP7_75t_L g1093 ( 
.A(n_960),
.B(n_856),
.Y(n_1093)
);

AOI21xp5_ASAP7_75t_L g1094 ( 
.A1(n_956),
.A2(n_846),
.B(n_869),
.Y(n_1094)
);

OAI21xp5_ASAP7_75t_L g1095 ( 
.A1(n_952),
.A2(n_858),
.B(n_844),
.Y(n_1095)
);

AOI21xp5_ASAP7_75t_L g1096 ( 
.A1(n_966),
.A2(n_869),
.B(n_872),
.Y(n_1096)
);

AND2x4_ASAP7_75t_L g1097 ( 
.A(n_1038),
.B(n_922),
.Y(n_1097)
);

AOI21xp5_ASAP7_75t_L g1098 ( 
.A1(n_1064),
.A2(n_907),
.B(n_922),
.Y(n_1098)
);

AOI21xp5_ASAP7_75t_L g1099 ( 
.A1(n_1064),
.A2(n_907),
.B(n_922),
.Y(n_1099)
);

INVx2_ASAP7_75t_SL g1100 ( 
.A(n_1040),
.Y(n_1100)
);

AOI21xp5_ASAP7_75t_L g1101 ( 
.A1(n_980),
.A2(n_907),
.B(n_922),
.Y(n_1101)
);

NAND2xp5_ASAP7_75t_L g1102 ( 
.A(n_1058),
.B(n_938),
.Y(n_1102)
);

NAND2xp5_ASAP7_75t_L g1103 ( 
.A(n_954),
.B(n_894),
.Y(n_1103)
);

OAI21x1_ASAP7_75t_L g1104 ( 
.A1(n_1066),
.A2(n_908),
.B(n_889),
.Y(n_1104)
);

OAI21xp5_ASAP7_75t_L g1105 ( 
.A1(n_1037),
.A2(n_908),
.B(n_906),
.Y(n_1105)
);

NAND2xp5_ASAP7_75t_L g1106 ( 
.A(n_965),
.B(n_867),
.Y(n_1106)
);

INVx2_ASAP7_75t_L g1107 ( 
.A(n_1020),
.Y(n_1107)
);

NAND2xp5_ASAP7_75t_L g1108 ( 
.A(n_1036),
.B(n_949),
.Y(n_1108)
);

OAI21xp5_ASAP7_75t_L g1109 ( 
.A1(n_1045),
.A2(n_968),
.B(n_1071),
.Y(n_1109)
);

INVx2_ASAP7_75t_L g1110 ( 
.A(n_1029),
.Y(n_1110)
);

AO31x2_ASAP7_75t_L g1111 ( 
.A1(n_992),
.A2(n_1075),
.A3(n_983),
.B(n_941),
.Y(n_1111)
);

AO31x2_ASAP7_75t_L g1112 ( 
.A1(n_941),
.A2(n_1062),
.A3(n_1056),
.B(n_943),
.Y(n_1112)
);

INVx1_ASAP7_75t_L g1113 ( 
.A(n_945),
.Y(n_1113)
);

OAI21xp5_ASAP7_75t_L g1114 ( 
.A1(n_1071),
.A2(n_1065),
.B(n_1050),
.Y(n_1114)
);

AOI21xp5_ASAP7_75t_L g1115 ( 
.A1(n_972),
.A2(n_950),
.B(n_949),
.Y(n_1115)
);

OAI21x1_ASAP7_75t_L g1116 ( 
.A1(n_962),
.A2(n_1049),
.B(n_1061),
.Y(n_1116)
);

AOI21xp5_ASAP7_75t_L g1117 ( 
.A1(n_978),
.A2(n_953),
.B(n_1003),
.Y(n_1117)
);

NAND3xp33_ASAP7_75t_L g1118 ( 
.A(n_1034),
.B(n_1059),
.C(n_1063),
.Y(n_1118)
);

INVxp67_ASAP7_75t_L g1119 ( 
.A(n_990),
.Y(n_1119)
);

AOI22xp5_ASAP7_75t_L g1120 ( 
.A1(n_1002),
.A2(n_1041),
.B1(n_947),
.B2(n_1019),
.Y(n_1120)
);

INVx1_ASAP7_75t_L g1121 ( 
.A(n_957),
.Y(n_1121)
);

NAND2xp5_ASAP7_75t_L g1122 ( 
.A(n_1036),
.B(n_988),
.Y(n_1122)
);

HB1xp67_ASAP7_75t_L g1123 ( 
.A(n_1010),
.Y(n_1123)
);

NAND2xp5_ASAP7_75t_L g1124 ( 
.A(n_967),
.B(n_993),
.Y(n_1124)
);

OAI21xp5_ASAP7_75t_L g1125 ( 
.A1(n_1076),
.A2(n_959),
.B(n_981),
.Y(n_1125)
);

OAI21x1_ASAP7_75t_L g1126 ( 
.A1(n_1067),
.A2(n_1073),
.B(n_1069),
.Y(n_1126)
);

OAI21xp5_ASAP7_75t_L g1127 ( 
.A1(n_981),
.A2(n_1013),
.B(n_1009),
.Y(n_1127)
);

AOI22xp5_ASAP7_75t_L g1128 ( 
.A1(n_1021),
.A2(n_1044),
.B1(n_1024),
.B2(n_1022),
.Y(n_1128)
);

OAI21x1_ASAP7_75t_L g1129 ( 
.A1(n_1068),
.A2(n_1006),
.B(n_961),
.Y(n_1129)
);

AOI21xp5_ASAP7_75t_L g1130 ( 
.A1(n_1009),
.A2(n_1013),
.B(n_1077),
.Y(n_1130)
);

AND2x2_ASAP7_75t_L g1131 ( 
.A(n_1016),
.B(n_942),
.Y(n_1131)
);

NOR2xp33_ASAP7_75t_L g1132 ( 
.A(n_1051),
.B(n_1057),
.Y(n_1132)
);

NAND2xp5_ASAP7_75t_L g1133 ( 
.A(n_1052),
.B(n_998),
.Y(n_1133)
);

AO31x2_ASAP7_75t_L g1134 ( 
.A1(n_1062),
.A2(n_1025),
.A3(n_1005),
.B(n_1060),
.Y(n_1134)
);

CKINVDCx5p33_ASAP7_75t_R g1135 ( 
.A(n_1000),
.Y(n_1135)
);

AOI21x1_ASAP7_75t_L g1136 ( 
.A1(n_1070),
.A2(n_1078),
.B(n_986),
.Y(n_1136)
);

AOI211x1_ASAP7_75t_L g1137 ( 
.A1(n_1033),
.A2(n_1005),
.B(n_1007),
.C(n_1047),
.Y(n_1137)
);

NAND2xp5_ASAP7_75t_L g1138 ( 
.A(n_1052),
.B(n_1001),
.Y(n_1138)
);

AOI221x1_ASAP7_75t_L g1139 ( 
.A1(n_1033),
.A2(n_1031),
.B1(n_1028),
.B2(n_1023),
.C(n_1026),
.Y(n_1139)
);

NAND2xp5_ASAP7_75t_L g1140 ( 
.A(n_963),
.B(n_973),
.Y(n_1140)
);

OAI21x1_ASAP7_75t_L g1141 ( 
.A1(n_961),
.A2(n_1078),
.B(n_1070),
.Y(n_1141)
);

NAND2xp5_ASAP7_75t_SL g1142 ( 
.A(n_964),
.B(n_1074),
.Y(n_1142)
);

AO21x2_ASAP7_75t_L g1143 ( 
.A1(n_975),
.A2(n_1008),
.B(n_1030),
.Y(n_1143)
);

INVx1_ASAP7_75t_SL g1144 ( 
.A(n_1053),
.Y(n_1144)
);

INVx1_ASAP7_75t_L g1145 ( 
.A(n_1035),
.Y(n_1145)
);

AND2x2_ASAP7_75t_L g1146 ( 
.A(n_994),
.B(n_1027),
.Y(n_1146)
);

INVx1_ASAP7_75t_L g1147 ( 
.A(n_970),
.Y(n_1147)
);

CKINVDCx11_ASAP7_75t_R g1148 ( 
.A(n_1043),
.Y(n_1148)
);

AND2x6_ASAP7_75t_L g1149 ( 
.A(n_997),
.B(n_1074),
.Y(n_1149)
);

NAND2xp5_ASAP7_75t_L g1150 ( 
.A(n_977),
.B(n_985),
.Y(n_1150)
);

A2O1A1Ixp33_ASAP7_75t_L g1151 ( 
.A1(n_999),
.A2(n_1011),
.B(n_1012),
.C(n_991),
.Y(n_1151)
);

NAND2xp5_ASAP7_75t_L g1152 ( 
.A(n_989),
.B(n_1018),
.Y(n_1152)
);

NAND2xp33_ASAP7_75t_L g1153 ( 
.A(n_1032),
.B(n_960),
.Y(n_1153)
);

INVx3_ASAP7_75t_L g1154 ( 
.A(n_960),
.Y(n_1154)
);

O2A1O1Ixp5_ASAP7_75t_SL g1155 ( 
.A1(n_971),
.A2(n_979),
.B(n_1042),
.C(n_1048),
.Y(n_1155)
);

AND2x2_ASAP7_75t_L g1156 ( 
.A(n_1055),
.B(n_997),
.Y(n_1156)
);

NAND2xp33_ASAP7_75t_L g1157 ( 
.A(n_1032),
.B(n_960),
.Y(n_1157)
);

NAND2xp5_ASAP7_75t_L g1158 ( 
.A(n_1004),
.B(n_1032),
.Y(n_1158)
);

NAND2xp5_ASAP7_75t_L g1159 ( 
.A(n_1054),
.B(n_971),
.Y(n_1159)
);

OR2x6_ASAP7_75t_L g1160 ( 
.A(n_1014),
.B(n_987),
.Y(n_1160)
);

NAND2xp5_ASAP7_75t_L g1161 ( 
.A(n_987),
.B(n_995),
.Y(n_1161)
);

OAI21xp5_ASAP7_75t_L g1162 ( 
.A1(n_1017),
.A2(n_969),
.B(n_1072),
.Y(n_1162)
);

INVx3_ASAP7_75t_L g1163 ( 
.A(n_969),
.Y(n_1163)
);

AOI21xp5_ASAP7_75t_L g1164 ( 
.A1(n_1072),
.A2(n_995),
.B(n_984),
.Y(n_1164)
);

NAND2xp5_ASAP7_75t_L g1165 ( 
.A(n_995),
.B(n_1039),
.Y(n_1165)
);

AND2x4_ASAP7_75t_L g1166 ( 
.A(n_1038),
.B(n_1052),
.Y(n_1166)
);

INVx4_ASAP7_75t_L g1167 ( 
.A(n_960),
.Y(n_1167)
);

CKINVDCx5p33_ASAP7_75t_R g1168 ( 
.A(n_944),
.Y(n_1168)
);

BUFx6f_ASAP7_75t_L g1169 ( 
.A(n_987),
.Y(n_1169)
);

BUFx2_ASAP7_75t_L g1170 ( 
.A(n_946),
.Y(n_1170)
);

AO31x2_ASAP7_75t_L g1171 ( 
.A1(n_1046),
.A2(n_982),
.A3(n_1015),
.B(n_951),
.Y(n_1171)
);

O2A1O1Ixp33_ASAP7_75t_L g1172 ( 
.A1(n_982),
.A2(n_606),
.B(n_878),
.C(n_685),
.Y(n_1172)
);

INVx2_ASAP7_75t_L g1173 ( 
.A(n_1020),
.Y(n_1173)
);

INVxp67_ASAP7_75t_SL g1174 ( 
.A(n_946),
.Y(n_1174)
);

NAND2xp5_ASAP7_75t_L g1175 ( 
.A(n_1039),
.B(n_616),
.Y(n_1175)
);

O2A1O1Ixp33_ASAP7_75t_SL g1176 ( 
.A1(n_982),
.A2(n_1015),
.B(n_972),
.C(n_877),
.Y(n_1176)
);

INVx1_ASAP7_75t_L g1177 ( 
.A(n_945),
.Y(n_1177)
);

INVx2_ASAP7_75t_L g1178 ( 
.A(n_1020),
.Y(n_1178)
);

NAND2xp5_ASAP7_75t_L g1179 ( 
.A(n_1039),
.B(n_616),
.Y(n_1179)
);

OAI21x1_ASAP7_75t_L g1180 ( 
.A1(n_996),
.A2(n_1066),
.B(n_1065),
.Y(n_1180)
);

INVx2_ASAP7_75t_SL g1181 ( 
.A(n_946),
.Y(n_1181)
);

OAI21x1_ASAP7_75t_L g1182 ( 
.A1(n_996),
.A2(n_1066),
.B(n_1065),
.Y(n_1182)
);

AOI21xp5_ASAP7_75t_L g1183 ( 
.A1(n_951),
.A2(n_701),
.B(n_775),
.Y(n_1183)
);

AOI21xp5_ASAP7_75t_L g1184 ( 
.A1(n_951),
.A2(n_701),
.B(n_775),
.Y(n_1184)
);

OAI21xp5_ASAP7_75t_L g1185 ( 
.A1(n_982),
.A2(n_955),
.B(n_951),
.Y(n_1185)
);

NAND2xp5_ASAP7_75t_L g1186 ( 
.A(n_1039),
.B(n_616),
.Y(n_1186)
);

OAI21x1_ASAP7_75t_L g1187 ( 
.A1(n_996),
.A2(n_1066),
.B(n_1065),
.Y(n_1187)
);

OAI22xp5_ASAP7_75t_L g1188 ( 
.A1(n_982),
.A2(n_767),
.B1(n_1064),
.B2(n_780),
.Y(n_1188)
);

BUFx6f_ASAP7_75t_L g1189 ( 
.A(n_987),
.Y(n_1189)
);

NOR2xp67_ASAP7_75t_L g1190 ( 
.A(n_944),
.B(n_788),
.Y(n_1190)
);

NAND2x1p5_ASAP7_75t_L g1191 ( 
.A(n_960),
.B(n_969),
.Y(n_1191)
);

OAI21x1_ASAP7_75t_L g1192 ( 
.A1(n_996),
.A2(n_1066),
.B(n_1065),
.Y(n_1192)
);

INVx3_ASAP7_75t_SL g1193 ( 
.A(n_944),
.Y(n_1193)
);

AND2x2_ASAP7_75t_L g1194 ( 
.A(n_976),
.B(n_788),
.Y(n_1194)
);

OAI21xp5_ASAP7_75t_L g1195 ( 
.A1(n_982),
.A2(n_955),
.B(n_951),
.Y(n_1195)
);

NAND2xp5_ASAP7_75t_L g1196 ( 
.A(n_1039),
.B(n_616),
.Y(n_1196)
);

CKINVDCx11_ASAP7_75t_R g1197 ( 
.A(n_1043),
.Y(n_1197)
);

INVx2_ASAP7_75t_L g1198 ( 
.A(n_1020),
.Y(n_1198)
);

NAND2xp5_ASAP7_75t_L g1199 ( 
.A(n_1039),
.B(n_616),
.Y(n_1199)
);

OAI21x1_ASAP7_75t_SL g1200 ( 
.A1(n_1046),
.A2(n_1059),
.B(n_1013),
.Y(n_1200)
);

AOI21xp5_ASAP7_75t_L g1201 ( 
.A1(n_951),
.A2(n_701),
.B(n_775),
.Y(n_1201)
);

NOR2xp33_ASAP7_75t_L g1202 ( 
.A(n_958),
.B(n_685),
.Y(n_1202)
);

OAI21x1_ASAP7_75t_L g1203 ( 
.A1(n_996),
.A2(n_1066),
.B(n_1065),
.Y(n_1203)
);

OAI21x1_ASAP7_75t_L g1204 ( 
.A1(n_996),
.A2(n_1066),
.B(n_1065),
.Y(n_1204)
);

AO31x2_ASAP7_75t_L g1205 ( 
.A1(n_1046),
.A2(n_982),
.A3(n_1015),
.B(n_951),
.Y(n_1205)
);

AOI21xp5_ASAP7_75t_L g1206 ( 
.A1(n_951),
.A2(n_701),
.B(n_775),
.Y(n_1206)
);

AOI21xp5_ASAP7_75t_L g1207 ( 
.A1(n_951),
.A2(n_701),
.B(n_775),
.Y(n_1207)
);

AOI221x1_ASAP7_75t_L g1208 ( 
.A1(n_982),
.A2(n_941),
.B1(n_1015),
.B2(n_951),
.C(n_966),
.Y(n_1208)
);

AOI21xp5_ASAP7_75t_L g1209 ( 
.A1(n_951),
.A2(n_701),
.B(n_775),
.Y(n_1209)
);

NAND2xp5_ASAP7_75t_L g1210 ( 
.A(n_1039),
.B(n_616),
.Y(n_1210)
);

A2O1A1Ixp33_ASAP7_75t_L g1211 ( 
.A1(n_982),
.A2(n_797),
.B(n_948),
.C(n_606),
.Y(n_1211)
);

INVx3_ASAP7_75t_L g1212 ( 
.A(n_1038),
.Y(n_1212)
);

OAI21x1_ASAP7_75t_L g1213 ( 
.A1(n_996),
.A2(n_1066),
.B(n_1065),
.Y(n_1213)
);

NAND2xp5_ASAP7_75t_L g1214 ( 
.A(n_1039),
.B(n_616),
.Y(n_1214)
);

OAI21x1_ASAP7_75t_L g1215 ( 
.A1(n_996),
.A2(n_1066),
.B(n_1065),
.Y(n_1215)
);

OAI21x1_ASAP7_75t_L g1216 ( 
.A1(n_996),
.A2(n_1066),
.B(n_1065),
.Y(n_1216)
);

AOI21xp5_ASAP7_75t_L g1217 ( 
.A1(n_951),
.A2(n_701),
.B(n_775),
.Y(n_1217)
);

OAI21xp5_ASAP7_75t_L g1218 ( 
.A1(n_1211),
.A2(n_1130),
.B(n_1127),
.Y(n_1218)
);

OAI21xp5_ASAP7_75t_L g1219 ( 
.A1(n_1127),
.A2(n_1172),
.B(n_1118),
.Y(n_1219)
);

HB1xp67_ASAP7_75t_L g1220 ( 
.A(n_1112),
.Y(n_1220)
);

OA21x2_ASAP7_75t_L g1221 ( 
.A1(n_1208),
.A2(n_1117),
.B(n_1185),
.Y(n_1221)
);

INVx2_ASAP7_75t_SL g1222 ( 
.A(n_1131),
.Y(n_1222)
);

OAI221xp5_ASAP7_75t_L g1223 ( 
.A1(n_1105),
.A2(n_1125),
.B1(n_1188),
.B2(n_1151),
.C(n_1118),
.Y(n_1223)
);

INVx1_ASAP7_75t_L g1224 ( 
.A(n_1113),
.Y(n_1224)
);

HB1xp67_ASAP7_75t_L g1225 ( 
.A(n_1112),
.Y(n_1225)
);

OAI21xp5_ASAP7_75t_L g1226 ( 
.A1(n_1115),
.A2(n_1125),
.B(n_1139),
.Y(n_1226)
);

BUFx12f_ASAP7_75t_L g1227 ( 
.A(n_1148),
.Y(n_1227)
);

AND2x2_ASAP7_75t_SL g1228 ( 
.A(n_1153),
.B(n_1157),
.Y(n_1228)
);

INVx1_ASAP7_75t_L g1229 ( 
.A(n_1121),
.Y(n_1229)
);

OAI21xp5_ASAP7_75t_L g1230 ( 
.A1(n_1103),
.A2(n_1188),
.B(n_1196),
.Y(n_1230)
);

NAND2xp5_ASAP7_75t_L g1231 ( 
.A(n_1175),
.B(n_1179),
.Y(n_1231)
);

AO21x2_ASAP7_75t_L g1232 ( 
.A1(n_1185),
.A2(n_1195),
.B(n_1200),
.Y(n_1232)
);

OR2x2_ASAP7_75t_L g1233 ( 
.A(n_1199),
.B(n_1210),
.Y(n_1233)
);

AO21x2_ASAP7_75t_L g1234 ( 
.A1(n_1195),
.A2(n_1114),
.B(n_1109),
.Y(n_1234)
);

OAI22xp5_ASAP7_75t_L g1235 ( 
.A1(n_1120),
.A2(n_1214),
.B1(n_1128),
.B2(n_1202),
.Y(n_1235)
);

AOI21xp33_ASAP7_75t_L g1236 ( 
.A1(n_1109),
.A2(n_1114),
.B(n_1175),
.Y(n_1236)
);

OAI21x1_ASAP7_75t_L g1237 ( 
.A1(n_1182),
.A2(n_1213),
.B(n_1204),
.Y(n_1237)
);

INVx2_ASAP7_75t_L g1238 ( 
.A(n_1107),
.Y(n_1238)
);

AO31x2_ASAP7_75t_L g1239 ( 
.A1(n_1098),
.A2(n_1099),
.A3(n_1209),
.B(n_1207),
.Y(n_1239)
);

O2A1O1Ixp33_ASAP7_75t_L g1240 ( 
.A1(n_1176),
.A2(n_1179),
.B(n_1186),
.C(n_1105),
.Y(n_1240)
);

OAI21xp5_ASAP7_75t_L g1241 ( 
.A1(n_1102),
.A2(n_1186),
.B(n_1087),
.Y(n_1241)
);

OA21x2_ASAP7_75t_L g1242 ( 
.A1(n_1095),
.A2(n_1187),
.B(n_1216),
.Y(n_1242)
);

OAI21x1_ASAP7_75t_L g1243 ( 
.A1(n_1192),
.A2(n_1215),
.B(n_1203),
.Y(n_1243)
);

BUFx3_ASAP7_75t_L g1244 ( 
.A(n_1170),
.Y(n_1244)
);

AO31x2_ASAP7_75t_L g1245 ( 
.A1(n_1183),
.A2(n_1217),
.A3(n_1206),
.B(n_1201),
.Y(n_1245)
);

OAI21x1_ASAP7_75t_L g1246 ( 
.A1(n_1096),
.A2(n_1094),
.B(n_1184),
.Y(n_1246)
);

INVx1_ASAP7_75t_L g1247 ( 
.A(n_1177),
.Y(n_1247)
);

NAND2xp5_ASAP7_75t_L g1248 ( 
.A(n_1122),
.B(n_1108),
.Y(n_1248)
);

INVx1_ASAP7_75t_L g1249 ( 
.A(n_1145),
.Y(n_1249)
);

INVx5_ASAP7_75t_L g1250 ( 
.A(n_1167),
.Y(n_1250)
);

BUFx6f_ASAP7_75t_L g1251 ( 
.A(n_1092),
.Y(n_1251)
);

INVx2_ASAP7_75t_L g1252 ( 
.A(n_1110),
.Y(n_1252)
);

OA21x2_ASAP7_75t_L g1253 ( 
.A1(n_1095),
.A2(n_1126),
.B(n_1091),
.Y(n_1253)
);

OAI21xp5_ASAP7_75t_L g1254 ( 
.A1(n_1087),
.A2(n_1088),
.B(n_1124),
.Y(n_1254)
);

AO21x2_ASAP7_75t_L g1255 ( 
.A1(n_1080),
.A2(n_1091),
.B(n_1136),
.Y(n_1255)
);

OAI21x1_ASAP7_75t_L g1256 ( 
.A1(n_1129),
.A2(n_1101),
.B(n_1089),
.Y(n_1256)
);

BUFx6f_ASAP7_75t_L g1257 ( 
.A(n_1092),
.Y(n_1257)
);

AO21x2_ASAP7_75t_L g1258 ( 
.A1(n_1143),
.A2(n_1141),
.B(n_1104),
.Y(n_1258)
);

INVx1_ASAP7_75t_L g1259 ( 
.A(n_1147),
.Y(n_1259)
);

BUFx2_ASAP7_75t_L g1260 ( 
.A(n_1086),
.Y(n_1260)
);

OAI21xp5_ASAP7_75t_L g1261 ( 
.A1(n_1082),
.A2(n_1155),
.B(n_1085),
.Y(n_1261)
);

INVx2_ASAP7_75t_SL g1262 ( 
.A(n_1168),
.Y(n_1262)
);

OAI22xp5_ASAP7_75t_L g1263 ( 
.A1(n_1158),
.A2(n_1106),
.B1(n_1194),
.B2(n_1174),
.Y(n_1263)
);

OAI22xp5_ASAP7_75t_L g1264 ( 
.A1(n_1190),
.A2(n_1119),
.B1(n_1146),
.B2(n_1181),
.Y(n_1264)
);

AND2x2_ASAP7_75t_L g1265 ( 
.A(n_1156),
.B(n_1166),
.Y(n_1265)
);

INVx1_ASAP7_75t_SL g1266 ( 
.A(n_1144),
.Y(n_1266)
);

INVx1_ASAP7_75t_L g1267 ( 
.A(n_1165),
.Y(n_1267)
);

BUFx2_ASAP7_75t_L g1268 ( 
.A(n_1123),
.Y(n_1268)
);

AOI22xp33_ASAP7_75t_L g1269 ( 
.A1(n_1149),
.A2(n_1143),
.B1(n_1079),
.B2(n_1173),
.Y(n_1269)
);

AOI22xp33_ASAP7_75t_SL g1270 ( 
.A1(n_1149),
.A2(n_1144),
.B1(n_1132),
.B2(n_1165),
.Y(n_1270)
);

A2O1A1Ixp33_ASAP7_75t_L g1271 ( 
.A1(n_1133),
.A2(n_1138),
.B(n_1198),
.C(n_1178),
.Y(n_1271)
);

OAI21x1_ASAP7_75t_L g1272 ( 
.A1(n_1162),
.A2(n_1093),
.B(n_1191),
.Y(n_1272)
);

INVx1_ASAP7_75t_L g1273 ( 
.A(n_1140),
.Y(n_1273)
);

OAI21x1_ASAP7_75t_L g1274 ( 
.A1(n_1154),
.A2(n_1163),
.B(n_1152),
.Y(n_1274)
);

O2A1O1Ixp33_ASAP7_75t_L g1275 ( 
.A1(n_1142),
.A2(n_1150),
.B(n_1100),
.C(n_1159),
.Y(n_1275)
);

HB1xp67_ASAP7_75t_L g1276 ( 
.A(n_1112),
.Y(n_1276)
);

AOI21xp33_ASAP7_75t_SL g1277 ( 
.A1(n_1193),
.A2(n_1135),
.B(n_1166),
.Y(n_1277)
);

BUFx2_ASAP7_75t_L g1278 ( 
.A(n_1161),
.Y(n_1278)
);

INVx1_ASAP7_75t_SL g1279 ( 
.A(n_1197),
.Y(n_1279)
);

NAND2x1p5_ASAP7_75t_L g1280 ( 
.A(n_1167),
.B(n_1212),
.Y(n_1280)
);

O2A1O1Ixp33_ASAP7_75t_SL g1281 ( 
.A1(n_1161),
.A2(n_1137),
.B(n_1212),
.C(n_1134),
.Y(n_1281)
);

NAND2xp5_ASAP7_75t_L g1282 ( 
.A(n_1134),
.B(n_1149),
.Y(n_1282)
);

OAI21xp5_ASAP7_75t_L g1283 ( 
.A1(n_1164),
.A2(n_1149),
.B(n_1083),
.Y(n_1283)
);

O2A1O1Ixp33_ASAP7_75t_SL g1284 ( 
.A1(n_1134),
.A2(n_1111),
.B(n_1081),
.C(n_1205),
.Y(n_1284)
);

CKINVDCx11_ASAP7_75t_R g1285 ( 
.A(n_1160),
.Y(n_1285)
);

CKINVDCx6p67_ASAP7_75t_R g1286 ( 
.A(n_1160),
.Y(n_1286)
);

OAI22x1_ASAP7_75t_L g1287 ( 
.A1(n_1083),
.A2(n_1097),
.B1(n_1111),
.B2(n_1171),
.Y(n_1287)
);

INVx1_ASAP7_75t_L g1288 ( 
.A(n_1081),
.Y(n_1288)
);

OAI222xp33_ASAP7_75t_L g1289 ( 
.A1(n_1160),
.A2(n_1111),
.B1(n_1097),
.B2(n_1205),
.C1(n_1171),
.C2(n_1084),
.Y(n_1289)
);

NAND2x1p5_ASAP7_75t_L g1290 ( 
.A(n_1092),
.B(n_1169),
.Y(n_1290)
);

OAI21x1_ASAP7_75t_L g1291 ( 
.A1(n_1084),
.A2(n_1171),
.B(n_1205),
.Y(n_1291)
);

INVx2_ASAP7_75t_SL g1292 ( 
.A(n_1169),
.Y(n_1292)
);

O2A1O1Ixp33_ASAP7_75t_SL g1293 ( 
.A1(n_1084),
.A2(n_1211),
.B(n_982),
.C(n_1188),
.Y(n_1293)
);

OAI21x1_ASAP7_75t_L g1294 ( 
.A1(n_1169),
.A2(n_1116),
.B(n_1090),
.Y(n_1294)
);

AOI221xp5_ASAP7_75t_L g1295 ( 
.A1(n_1189),
.A2(n_606),
.B1(n_1188),
.B2(n_767),
.C(n_1172),
.Y(n_1295)
);

INVx4_ASAP7_75t_L g1296 ( 
.A(n_1189),
.Y(n_1296)
);

AOI22xp33_ASAP7_75t_L g1297 ( 
.A1(n_1188),
.A2(n_606),
.B1(n_767),
.B2(n_918),
.Y(n_1297)
);

NOR3xp33_ASAP7_75t_SL g1298 ( 
.A(n_1211),
.B(n_1026),
.C(n_1023),
.Y(n_1298)
);

AOI21x1_ASAP7_75t_L g1299 ( 
.A1(n_1130),
.A2(n_966),
.B(n_1183),
.Y(n_1299)
);

OAI22xp5_ASAP7_75t_L g1300 ( 
.A1(n_1103),
.A2(n_606),
.B1(n_864),
.B2(n_982),
.Y(n_1300)
);

O2A1O1Ixp33_ASAP7_75t_L g1301 ( 
.A1(n_1211),
.A2(n_982),
.B(n_1172),
.C(n_606),
.Y(n_1301)
);

OA21x2_ASAP7_75t_L g1302 ( 
.A1(n_1208),
.A2(n_1117),
.B(n_1185),
.Y(n_1302)
);

NAND2xp5_ASAP7_75t_L g1303 ( 
.A(n_1175),
.B(n_1179),
.Y(n_1303)
);

OAI222xp33_ASAP7_75t_L g1304 ( 
.A1(n_1188),
.A2(n_1033),
.B1(n_1005),
.B2(n_767),
.C1(n_941),
.C2(n_972),
.Y(n_1304)
);

INVx2_ASAP7_75t_L g1305 ( 
.A(n_1107),
.Y(n_1305)
);

O2A1O1Ixp33_ASAP7_75t_L g1306 ( 
.A1(n_1211),
.A2(n_982),
.B(n_1172),
.C(n_606),
.Y(n_1306)
);

CKINVDCx20_ASAP7_75t_R g1307 ( 
.A(n_1148),
.Y(n_1307)
);

OAI21x1_ASAP7_75t_L g1308 ( 
.A1(n_1116),
.A2(n_1090),
.B(n_1180),
.Y(n_1308)
);

OAI22xp5_ASAP7_75t_L g1309 ( 
.A1(n_1103),
.A2(n_606),
.B1(n_864),
.B2(n_982),
.Y(n_1309)
);

AOI222xp33_ASAP7_75t_L g1310 ( 
.A1(n_1188),
.A2(n_606),
.B1(n_562),
.B2(n_418),
.C1(n_767),
.C2(n_678),
.Y(n_1310)
);

NOR2xp33_ASAP7_75t_L g1311 ( 
.A(n_1103),
.B(n_606),
.Y(n_1311)
);

INVx1_ASAP7_75t_L g1312 ( 
.A(n_1113),
.Y(n_1312)
);

INVx2_ASAP7_75t_L g1313 ( 
.A(n_1107),
.Y(n_1313)
);

AND2x4_ASAP7_75t_L g1314 ( 
.A(n_1166),
.B(n_1083),
.Y(n_1314)
);

AOI21xp5_ASAP7_75t_L g1315 ( 
.A1(n_1114),
.A2(n_1211),
.B(n_1109),
.Y(n_1315)
);

AO31x2_ASAP7_75t_L g1316 ( 
.A1(n_1208),
.A2(n_1211),
.A3(n_1046),
.B(n_982),
.Y(n_1316)
);

CKINVDCx5p33_ASAP7_75t_R g1317 ( 
.A(n_1168),
.Y(n_1317)
);

AOI22xp5_ASAP7_75t_L g1318 ( 
.A1(n_1082),
.A2(n_606),
.B1(n_591),
.B2(n_308),
.Y(n_1318)
);

AND2x2_ASAP7_75t_L g1319 ( 
.A(n_1194),
.B(n_732),
.Y(n_1319)
);

INVx2_ASAP7_75t_L g1320 ( 
.A(n_1107),
.Y(n_1320)
);

INVx1_ASAP7_75t_L g1321 ( 
.A(n_1113),
.Y(n_1321)
);

INVx1_ASAP7_75t_L g1322 ( 
.A(n_1113),
.Y(n_1322)
);

AO21x2_ASAP7_75t_L g1323 ( 
.A1(n_1185),
.A2(n_1195),
.B(n_1200),
.Y(n_1323)
);

OAI21x1_ASAP7_75t_L g1324 ( 
.A1(n_1116),
.A2(n_1090),
.B(n_1180),
.Y(n_1324)
);

AOI21xp5_ASAP7_75t_L g1325 ( 
.A1(n_1114),
.A2(n_1211),
.B(n_1109),
.Y(n_1325)
);

OAI21x1_ASAP7_75t_L g1326 ( 
.A1(n_1116),
.A2(n_1090),
.B(n_1180),
.Y(n_1326)
);

NOR2xp33_ASAP7_75t_L g1327 ( 
.A(n_1103),
.B(n_606),
.Y(n_1327)
);

INVx1_ASAP7_75t_SL g1328 ( 
.A(n_1170),
.Y(n_1328)
);

BUFx2_ASAP7_75t_R g1329 ( 
.A(n_1168),
.Y(n_1329)
);

INVx4_ASAP7_75t_L g1330 ( 
.A(n_1160),
.Y(n_1330)
);

AO31x2_ASAP7_75t_L g1331 ( 
.A1(n_1208),
.A2(n_1211),
.A3(n_1046),
.B(n_982),
.Y(n_1331)
);

AOI22xp5_ASAP7_75t_L g1332 ( 
.A1(n_1082),
.A2(n_606),
.B1(n_591),
.B2(n_308),
.Y(n_1332)
);

AOI22xp5_ASAP7_75t_L g1333 ( 
.A1(n_1082),
.A2(n_606),
.B1(n_591),
.B2(n_308),
.Y(n_1333)
);

INVx1_ASAP7_75t_L g1334 ( 
.A(n_1113),
.Y(n_1334)
);

AOI22xp33_ASAP7_75t_L g1335 ( 
.A1(n_1188),
.A2(n_606),
.B1(n_767),
.B2(n_918),
.Y(n_1335)
);

AO31x2_ASAP7_75t_L g1336 ( 
.A1(n_1208),
.A2(n_1211),
.A3(n_1046),
.B(n_982),
.Y(n_1336)
);

OAI21x1_ASAP7_75t_L g1337 ( 
.A1(n_1116),
.A2(n_1090),
.B(n_1180),
.Y(n_1337)
);

AO31x2_ASAP7_75t_L g1338 ( 
.A1(n_1208),
.A2(n_1211),
.A3(n_1046),
.B(n_982),
.Y(n_1338)
);

NOR2xp33_ASAP7_75t_L g1339 ( 
.A(n_1103),
.B(n_606),
.Y(n_1339)
);

OAI21xp5_ASAP7_75t_L g1340 ( 
.A1(n_1211),
.A2(n_473),
.B(n_982),
.Y(n_1340)
);

INVx2_ASAP7_75t_L g1341 ( 
.A(n_1288),
.Y(n_1341)
);

NAND2xp5_ASAP7_75t_L g1342 ( 
.A(n_1311),
.B(n_1327),
.Y(n_1342)
);

OR2x2_ASAP7_75t_SL g1343 ( 
.A(n_1233),
.B(n_1231),
.Y(n_1343)
);

CKINVDCx5p33_ASAP7_75t_R g1344 ( 
.A(n_1329),
.Y(n_1344)
);

AND2x2_ASAP7_75t_L g1345 ( 
.A(n_1298),
.B(n_1265),
.Y(n_1345)
);

INVxp67_ASAP7_75t_L g1346 ( 
.A(n_1260),
.Y(n_1346)
);

OAI22xp5_ASAP7_75t_L g1347 ( 
.A1(n_1297),
.A2(n_1335),
.B1(n_1318),
.B2(n_1333),
.Y(n_1347)
);

OAI22xp5_ASAP7_75t_L g1348 ( 
.A1(n_1297),
.A2(n_1335),
.B1(n_1332),
.B2(n_1298),
.Y(n_1348)
);

AOI21xp5_ASAP7_75t_SL g1349 ( 
.A1(n_1340),
.A2(n_1306),
.B(n_1301),
.Y(n_1349)
);

HB1xp67_ASAP7_75t_L g1350 ( 
.A(n_1220),
.Y(n_1350)
);

NAND2xp5_ASAP7_75t_L g1351 ( 
.A(n_1311),
.B(n_1327),
.Y(n_1351)
);

NAND2xp5_ASAP7_75t_L g1352 ( 
.A(n_1339),
.B(n_1248),
.Y(n_1352)
);

OAI22xp5_ASAP7_75t_L g1353 ( 
.A1(n_1223),
.A2(n_1339),
.B1(n_1235),
.B2(n_1263),
.Y(n_1353)
);

OAI22xp5_ASAP7_75t_SL g1354 ( 
.A1(n_1223),
.A2(n_1307),
.B1(n_1270),
.B2(n_1266),
.Y(n_1354)
);

AND2x2_ASAP7_75t_L g1355 ( 
.A(n_1278),
.B(n_1319),
.Y(n_1355)
);

AOI21xp5_ASAP7_75t_L g1356 ( 
.A1(n_1218),
.A2(n_1226),
.B(n_1325),
.Y(n_1356)
);

AND2x2_ASAP7_75t_L g1357 ( 
.A(n_1314),
.B(n_1267),
.Y(n_1357)
);

NAND2xp5_ASAP7_75t_L g1358 ( 
.A(n_1248),
.B(n_1231),
.Y(n_1358)
);

NAND2xp5_ASAP7_75t_L g1359 ( 
.A(n_1303),
.B(n_1273),
.Y(n_1359)
);

NAND2xp5_ASAP7_75t_L g1360 ( 
.A(n_1303),
.B(n_1230),
.Y(n_1360)
);

AOI21xp5_ASAP7_75t_SL g1361 ( 
.A1(n_1301),
.A2(n_1306),
.B(n_1295),
.Y(n_1361)
);

BUFx12f_ASAP7_75t_L g1362 ( 
.A(n_1227),
.Y(n_1362)
);

AOI21xp5_ASAP7_75t_L g1363 ( 
.A1(n_1315),
.A2(n_1325),
.B(n_1304),
.Y(n_1363)
);

AND2x4_ASAP7_75t_L g1364 ( 
.A(n_1283),
.B(n_1314),
.Y(n_1364)
);

AOI21x1_ASAP7_75t_SL g1365 ( 
.A1(n_1282),
.A2(n_1220),
.B(n_1276),
.Y(n_1365)
);

AND2x4_ASAP7_75t_SL g1366 ( 
.A(n_1330),
.B(n_1286),
.Y(n_1366)
);

OAI22xp5_ASAP7_75t_L g1367 ( 
.A1(n_1270),
.A2(n_1309),
.B1(n_1300),
.B2(n_1222),
.Y(n_1367)
);

AND2x4_ASAP7_75t_L g1368 ( 
.A(n_1229),
.B(n_1247),
.Y(n_1368)
);

AND2x2_ASAP7_75t_L g1369 ( 
.A(n_1238),
.B(n_1252),
.Y(n_1369)
);

AOI22xp5_ASAP7_75t_L g1370 ( 
.A1(n_1310),
.A2(n_1264),
.B1(n_1295),
.B2(n_1219),
.Y(n_1370)
);

AND2x2_ASAP7_75t_L g1371 ( 
.A(n_1305),
.B(n_1313),
.Y(n_1371)
);

AOI21xp5_ASAP7_75t_SL g1372 ( 
.A1(n_1240),
.A2(n_1275),
.B(n_1241),
.Y(n_1372)
);

OAI22xp5_ASAP7_75t_L g1373 ( 
.A1(n_1328),
.A2(n_1244),
.B1(n_1228),
.B2(n_1268),
.Y(n_1373)
);

AND2x2_ASAP7_75t_L g1374 ( 
.A(n_1320),
.B(n_1249),
.Y(n_1374)
);

OAI22xp5_ASAP7_75t_SL g1375 ( 
.A1(n_1279),
.A2(n_1262),
.B1(n_1317),
.B2(n_1228),
.Y(n_1375)
);

NAND2xp5_ASAP7_75t_L g1376 ( 
.A(n_1240),
.B(n_1275),
.Y(n_1376)
);

OA21x2_ASAP7_75t_L g1377 ( 
.A1(n_1291),
.A2(n_1246),
.B(n_1315),
.Y(n_1377)
);

AND2x2_ASAP7_75t_L g1378 ( 
.A(n_1259),
.B(n_1312),
.Y(n_1378)
);

NAND2x1_ASAP7_75t_L g1379 ( 
.A(n_1330),
.B(n_1254),
.Y(n_1379)
);

CKINVDCx5p33_ASAP7_75t_R g1380 ( 
.A(n_1329),
.Y(n_1380)
);

OAI22xp5_ASAP7_75t_L g1381 ( 
.A1(n_1282),
.A2(n_1269),
.B1(n_1271),
.B2(n_1321),
.Y(n_1381)
);

AOI21xp5_ASAP7_75t_L g1382 ( 
.A1(n_1304),
.A2(n_1234),
.B(n_1293),
.Y(n_1382)
);

AND2x2_ASAP7_75t_L g1383 ( 
.A(n_1322),
.B(n_1334),
.Y(n_1383)
);

AOI21xp5_ASAP7_75t_SL g1384 ( 
.A1(n_1271),
.A2(n_1261),
.B(n_1221),
.Y(n_1384)
);

OR2x2_ASAP7_75t_L g1385 ( 
.A(n_1234),
.B(n_1331),
.Y(n_1385)
);

AOI21xp5_ASAP7_75t_L g1386 ( 
.A1(n_1293),
.A2(n_1236),
.B(n_1302),
.Y(n_1386)
);

OAI22xp5_ASAP7_75t_SL g1387 ( 
.A1(n_1221),
.A2(n_1302),
.B1(n_1280),
.B2(n_1296),
.Y(n_1387)
);

AOI21x1_ASAP7_75t_SL g1388 ( 
.A1(n_1225),
.A2(n_1276),
.B(n_1289),
.Y(n_1388)
);

INVx1_ASAP7_75t_L g1389 ( 
.A(n_1287),
.Y(n_1389)
);

AOI21xp5_ASAP7_75t_L g1390 ( 
.A1(n_1236),
.A2(n_1232),
.B(n_1323),
.Y(n_1390)
);

AOI31xp33_ASAP7_75t_L g1391 ( 
.A1(n_1277),
.A2(n_1280),
.A3(n_1269),
.B(n_1281),
.Y(n_1391)
);

AND2x2_ASAP7_75t_L g1392 ( 
.A(n_1251),
.B(n_1257),
.Y(n_1392)
);

NAND2xp5_ASAP7_75t_L g1393 ( 
.A(n_1232),
.B(n_1323),
.Y(n_1393)
);

AO21x2_ASAP7_75t_L g1394 ( 
.A1(n_1299),
.A2(n_1324),
.B(n_1337),
.Y(n_1394)
);

OAI22xp5_ASAP7_75t_L g1395 ( 
.A1(n_1250),
.A2(n_1292),
.B1(n_1296),
.B2(n_1290),
.Y(n_1395)
);

AND2x2_ASAP7_75t_L g1396 ( 
.A(n_1257),
.B(n_1285),
.Y(n_1396)
);

OAI22xp5_ASAP7_75t_L g1397 ( 
.A1(n_1250),
.A2(n_1285),
.B1(n_1253),
.B2(n_1242),
.Y(n_1397)
);

O2A1O1Ixp33_ASAP7_75t_L g1398 ( 
.A1(n_1289),
.A2(n_1284),
.B(n_1255),
.C(n_1258),
.Y(n_1398)
);

O2A1O1Ixp5_ASAP7_75t_L g1399 ( 
.A1(n_1316),
.A2(n_1338),
.B(n_1336),
.C(n_1331),
.Y(n_1399)
);

BUFx6f_ASAP7_75t_L g1400 ( 
.A(n_1250),
.Y(n_1400)
);

NAND2xp5_ASAP7_75t_L g1401 ( 
.A(n_1316),
.B(n_1338),
.Y(n_1401)
);

O2A1O1Ixp5_ASAP7_75t_L g1402 ( 
.A1(n_1336),
.A2(n_1245),
.B(n_1239),
.C(n_1258),
.Y(n_1402)
);

AOI21x1_ASAP7_75t_SL g1403 ( 
.A1(n_1239),
.A2(n_1245),
.B(n_1294),
.Y(n_1403)
);

AND2x2_ASAP7_75t_L g1404 ( 
.A(n_1274),
.B(n_1272),
.Y(n_1404)
);

AOI21x1_ASAP7_75t_SL g1405 ( 
.A1(n_1239),
.A2(n_1245),
.B(n_1256),
.Y(n_1405)
);

AND2x4_ASAP7_75t_L g1406 ( 
.A(n_1245),
.B(n_1308),
.Y(n_1406)
);

OAI22xp5_ASAP7_75t_L g1407 ( 
.A1(n_1326),
.A2(n_1335),
.B1(n_1297),
.B2(n_864),
.Y(n_1407)
);

OAI22xp5_ASAP7_75t_L g1408 ( 
.A1(n_1237),
.A2(n_1335),
.B1(n_1297),
.B2(n_864),
.Y(n_1408)
);

AND2x4_ASAP7_75t_L g1409 ( 
.A(n_1243),
.B(n_1283),
.Y(n_1409)
);

AND2x2_ASAP7_75t_L g1410 ( 
.A(n_1298),
.B(n_1265),
.Y(n_1410)
);

OR2x2_ASAP7_75t_L g1411 ( 
.A(n_1263),
.B(n_1267),
.Y(n_1411)
);

OAI22xp5_ASAP7_75t_L g1412 ( 
.A1(n_1297),
.A2(n_1335),
.B1(n_864),
.B2(n_1332),
.Y(n_1412)
);

INVx1_ASAP7_75t_L g1413 ( 
.A(n_1224),
.Y(n_1413)
);

AND2x2_ASAP7_75t_L g1414 ( 
.A(n_1298),
.B(n_1265),
.Y(n_1414)
);

OA21x2_ASAP7_75t_L g1415 ( 
.A1(n_1226),
.A2(n_1208),
.B(n_1218),
.Y(n_1415)
);

BUFx3_ASAP7_75t_L g1416 ( 
.A(n_1244),
.Y(n_1416)
);

NAND2xp5_ASAP7_75t_L g1417 ( 
.A(n_1311),
.B(n_1327),
.Y(n_1417)
);

OAI22xp5_ASAP7_75t_L g1418 ( 
.A1(n_1297),
.A2(n_1335),
.B1(n_864),
.B2(n_1332),
.Y(n_1418)
);

O2A1O1Ixp33_ASAP7_75t_L g1419 ( 
.A1(n_1310),
.A2(n_1211),
.B(n_982),
.C(n_1340),
.Y(n_1419)
);

NAND2xp5_ASAP7_75t_L g1420 ( 
.A(n_1311),
.B(n_1327),
.Y(n_1420)
);

NOR2x1_ASAP7_75t_SL g1421 ( 
.A(n_1232),
.B(n_1323),
.Y(n_1421)
);

OA21x2_ASAP7_75t_L g1422 ( 
.A1(n_1226),
.A2(n_1208),
.B(n_1218),
.Y(n_1422)
);

INVx3_ASAP7_75t_SL g1423 ( 
.A(n_1317),
.Y(n_1423)
);

OR2x2_ASAP7_75t_L g1424 ( 
.A(n_1263),
.B(n_1267),
.Y(n_1424)
);

OAI22xp5_ASAP7_75t_L g1425 ( 
.A1(n_1297),
.A2(n_1335),
.B1(n_864),
.B2(n_1332),
.Y(n_1425)
);

AND2x2_ASAP7_75t_L g1426 ( 
.A(n_1298),
.B(n_1265),
.Y(n_1426)
);

INVx1_ASAP7_75t_L g1427 ( 
.A(n_1224),
.Y(n_1427)
);

AOI221xp5_ASAP7_75t_L g1428 ( 
.A1(n_1297),
.A2(n_606),
.B1(n_1335),
.B2(n_1223),
.C(n_1340),
.Y(n_1428)
);

BUFx2_ASAP7_75t_L g1429 ( 
.A(n_1244),
.Y(n_1429)
);

HB1xp67_ASAP7_75t_L g1430 ( 
.A(n_1350),
.Y(n_1430)
);

HB1xp67_ASAP7_75t_L g1431 ( 
.A(n_1350),
.Y(n_1431)
);

AOI22xp33_ASAP7_75t_L g1432 ( 
.A1(n_1347),
.A2(n_1348),
.B1(n_1428),
.B2(n_1418),
.Y(n_1432)
);

INVx2_ASAP7_75t_L g1433 ( 
.A(n_1341),
.Y(n_1433)
);

AO21x2_ASAP7_75t_L g1434 ( 
.A1(n_1356),
.A2(n_1363),
.B(n_1390),
.Y(n_1434)
);

AO21x2_ASAP7_75t_L g1435 ( 
.A1(n_1382),
.A2(n_1386),
.B(n_1421),
.Y(n_1435)
);

BUFx6f_ASAP7_75t_L g1436 ( 
.A(n_1409),
.Y(n_1436)
);

OAI21x1_ASAP7_75t_L g1437 ( 
.A1(n_1405),
.A2(n_1403),
.B(n_1402),
.Y(n_1437)
);

NAND2xp5_ASAP7_75t_L g1438 ( 
.A(n_1360),
.B(n_1358),
.Y(n_1438)
);

INVx1_ASAP7_75t_SL g1439 ( 
.A(n_1343),
.Y(n_1439)
);

INVx1_ASAP7_75t_L g1440 ( 
.A(n_1399),
.Y(n_1440)
);

INVx1_ASAP7_75t_L g1441 ( 
.A(n_1399),
.Y(n_1441)
);

OR2x2_ASAP7_75t_L g1442 ( 
.A(n_1385),
.B(n_1393),
.Y(n_1442)
);

INVx1_ASAP7_75t_L g1443 ( 
.A(n_1401),
.Y(n_1443)
);

AND2x2_ASAP7_75t_L g1444 ( 
.A(n_1415),
.B(n_1422),
.Y(n_1444)
);

BUFx4f_ASAP7_75t_L g1445 ( 
.A(n_1400),
.Y(n_1445)
);

HB1xp67_ASAP7_75t_SL g1446 ( 
.A(n_1344),
.Y(n_1446)
);

AOI22xp33_ASAP7_75t_L g1447 ( 
.A1(n_1412),
.A2(n_1425),
.B1(n_1353),
.B2(n_1370),
.Y(n_1447)
);

AND2x2_ASAP7_75t_L g1448 ( 
.A(n_1415),
.B(n_1422),
.Y(n_1448)
);

INVxp67_ASAP7_75t_SL g1449 ( 
.A(n_1376),
.Y(n_1449)
);

AND2x2_ASAP7_75t_L g1450 ( 
.A(n_1415),
.B(n_1422),
.Y(n_1450)
);

INVx2_ASAP7_75t_L g1451 ( 
.A(n_1377),
.Y(n_1451)
);

INVx2_ASAP7_75t_L g1452 ( 
.A(n_1377),
.Y(n_1452)
);

INVx2_ASAP7_75t_L g1453 ( 
.A(n_1377),
.Y(n_1453)
);

INVx1_ASAP7_75t_SL g1454 ( 
.A(n_1411),
.Y(n_1454)
);

AND2x4_ASAP7_75t_L g1455 ( 
.A(n_1409),
.B(n_1404),
.Y(n_1455)
);

AND2x2_ASAP7_75t_L g1456 ( 
.A(n_1389),
.B(n_1406),
.Y(n_1456)
);

OA21x2_ASAP7_75t_L g1457 ( 
.A1(n_1381),
.A2(n_1397),
.B(n_1407),
.Y(n_1457)
);

NAND2xp5_ASAP7_75t_L g1458 ( 
.A(n_1352),
.B(n_1359),
.Y(n_1458)
);

AND2x2_ASAP7_75t_L g1459 ( 
.A(n_1409),
.B(n_1368),
.Y(n_1459)
);

BUFx2_ASAP7_75t_L g1460 ( 
.A(n_1394),
.Y(n_1460)
);

HB1xp67_ASAP7_75t_L g1461 ( 
.A(n_1346),
.Y(n_1461)
);

AO21x2_ASAP7_75t_L g1462 ( 
.A1(n_1384),
.A2(n_1349),
.B(n_1398),
.Y(n_1462)
);

NAND2xp5_ASAP7_75t_L g1463 ( 
.A(n_1424),
.B(n_1342),
.Y(n_1463)
);

BUFx3_ASAP7_75t_L g1464 ( 
.A(n_1379),
.Y(n_1464)
);

AND2x2_ASAP7_75t_L g1465 ( 
.A(n_1368),
.B(n_1427),
.Y(n_1465)
);

AOI22xp33_ASAP7_75t_L g1466 ( 
.A1(n_1354),
.A2(n_1417),
.B1(n_1351),
.B2(n_1420),
.Y(n_1466)
);

INVx1_ASAP7_75t_SL g1467 ( 
.A(n_1368),
.Y(n_1467)
);

NAND2xp5_ASAP7_75t_L g1468 ( 
.A(n_1413),
.B(n_1346),
.Y(n_1468)
);

AND2x4_ASAP7_75t_L g1469 ( 
.A(n_1394),
.B(n_1364),
.Y(n_1469)
);

AO21x2_ASAP7_75t_L g1470 ( 
.A1(n_1361),
.A2(n_1372),
.B(n_1408),
.Y(n_1470)
);

INVxp67_ASAP7_75t_L g1471 ( 
.A(n_1378),
.Y(n_1471)
);

AOI22xp33_ASAP7_75t_L g1472 ( 
.A1(n_1432),
.A2(n_1367),
.B1(n_1345),
.B2(n_1414),
.Y(n_1472)
);

NAND2xp5_ASAP7_75t_L g1473 ( 
.A(n_1449),
.B(n_1454),
.Y(n_1473)
);

AND2x4_ASAP7_75t_L g1474 ( 
.A(n_1436),
.B(n_1364),
.Y(n_1474)
);

INVx1_ASAP7_75t_L g1475 ( 
.A(n_1433),
.Y(n_1475)
);

NAND2xp5_ASAP7_75t_L g1476 ( 
.A(n_1449),
.B(n_1383),
.Y(n_1476)
);

BUFx3_ASAP7_75t_L g1477 ( 
.A(n_1464),
.Y(n_1477)
);

OAI31xp33_ASAP7_75t_L g1478 ( 
.A1(n_1432),
.A2(n_1447),
.A3(n_1419),
.B(n_1466),
.Y(n_1478)
);

INVx2_ASAP7_75t_SL g1479 ( 
.A(n_1436),
.Y(n_1479)
);

NAND2xp5_ASAP7_75t_L g1480 ( 
.A(n_1454),
.B(n_1374),
.Y(n_1480)
);

HB1xp67_ASAP7_75t_L g1481 ( 
.A(n_1430),
.Y(n_1481)
);

NAND3xp33_ASAP7_75t_L g1482 ( 
.A(n_1466),
.B(n_1373),
.C(n_1426),
.Y(n_1482)
);

NAND2xp5_ASAP7_75t_L g1483 ( 
.A(n_1442),
.B(n_1355),
.Y(n_1483)
);

OR2x2_ASAP7_75t_L g1484 ( 
.A(n_1442),
.B(n_1387),
.Y(n_1484)
);

AND2x2_ASAP7_75t_L g1485 ( 
.A(n_1450),
.B(n_1410),
.Y(n_1485)
);

AND2x2_ASAP7_75t_L g1486 ( 
.A(n_1444),
.B(n_1448),
.Y(n_1486)
);

AND2x2_ASAP7_75t_L g1487 ( 
.A(n_1444),
.B(n_1357),
.Y(n_1487)
);

OR2x2_ASAP7_75t_L g1488 ( 
.A(n_1448),
.B(n_1391),
.Y(n_1488)
);

AND2x2_ASAP7_75t_L g1489 ( 
.A(n_1450),
.B(n_1392),
.Y(n_1489)
);

OA21x2_ASAP7_75t_L g1490 ( 
.A1(n_1437),
.A2(n_1365),
.B(n_1388),
.Y(n_1490)
);

INVxp67_ASAP7_75t_SL g1491 ( 
.A(n_1431),
.Y(n_1491)
);

AND2x2_ASAP7_75t_L g1492 ( 
.A(n_1450),
.B(n_1369),
.Y(n_1492)
);

OR2x2_ASAP7_75t_L g1493 ( 
.A(n_1440),
.B(n_1429),
.Y(n_1493)
);

NAND2xp5_ASAP7_75t_L g1494 ( 
.A(n_1463),
.B(n_1371),
.Y(n_1494)
);

BUFx2_ASAP7_75t_L g1495 ( 
.A(n_1477),
.Y(n_1495)
);

INVxp67_ASAP7_75t_L g1496 ( 
.A(n_1483),
.Y(n_1496)
);

OR2x6_ASAP7_75t_L g1497 ( 
.A(n_1479),
.B(n_1464),
.Y(n_1497)
);

AOI22xp33_ASAP7_75t_L g1498 ( 
.A1(n_1478),
.A2(n_1470),
.B1(n_1447),
.B2(n_1462),
.Y(n_1498)
);

NOR2x2_ASAP7_75t_L g1499 ( 
.A(n_1482),
.B(n_1446),
.Y(n_1499)
);

AOI22xp5_ASAP7_75t_L g1500 ( 
.A1(n_1472),
.A2(n_1470),
.B1(n_1462),
.B2(n_1439),
.Y(n_1500)
);

AND2x2_ASAP7_75t_L g1501 ( 
.A(n_1485),
.B(n_1459),
.Y(n_1501)
);

OAI31xp33_ASAP7_75t_L g1502 ( 
.A1(n_1478),
.A2(n_1439),
.A3(n_1464),
.B(n_1375),
.Y(n_1502)
);

BUFx2_ASAP7_75t_L g1503 ( 
.A(n_1477),
.Y(n_1503)
);

INVx1_ASAP7_75t_L g1504 ( 
.A(n_1475),
.Y(n_1504)
);

OAI33xp33_ASAP7_75t_L g1505 ( 
.A1(n_1473),
.A2(n_1463),
.A3(n_1468),
.B1(n_1438),
.B2(n_1458),
.B3(n_1443),
.Y(n_1505)
);

HB1xp67_ASAP7_75t_L g1506 ( 
.A(n_1481),
.Y(n_1506)
);

NAND3xp33_ASAP7_75t_L g1507 ( 
.A(n_1472),
.B(n_1457),
.C(n_1461),
.Y(n_1507)
);

INVx1_ASAP7_75t_L g1508 ( 
.A(n_1475),
.Y(n_1508)
);

AO21x1_ASAP7_75t_SL g1509 ( 
.A1(n_1488),
.A2(n_1484),
.B(n_1473),
.Y(n_1509)
);

NOR4xp25_ASAP7_75t_SL g1510 ( 
.A(n_1491),
.B(n_1344),
.C(n_1380),
.D(n_1460),
.Y(n_1510)
);

AND2x2_ASAP7_75t_L g1511 ( 
.A(n_1485),
.B(n_1459),
.Y(n_1511)
);

AOI221xp5_ASAP7_75t_L g1512 ( 
.A1(n_1482),
.A2(n_1438),
.B1(n_1458),
.B2(n_1461),
.C(n_1434),
.Y(n_1512)
);

AND2x2_ASAP7_75t_L g1513 ( 
.A(n_1485),
.B(n_1459),
.Y(n_1513)
);

NAND2xp33_ASAP7_75t_R g1514 ( 
.A(n_1476),
.B(n_1380),
.Y(n_1514)
);

OR2x2_ASAP7_75t_L g1515 ( 
.A(n_1493),
.B(n_1434),
.Y(n_1515)
);

NAND2xp33_ASAP7_75t_R g1516 ( 
.A(n_1476),
.B(n_1457),
.Y(n_1516)
);

AOI22xp33_ASAP7_75t_L g1517 ( 
.A1(n_1482),
.A2(n_1470),
.B1(n_1462),
.B2(n_1457),
.Y(n_1517)
);

AOI22xp33_ASAP7_75t_L g1518 ( 
.A1(n_1488),
.A2(n_1470),
.B1(n_1462),
.B2(n_1457),
.Y(n_1518)
);

AND2x2_ASAP7_75t_L g1519 ( 
.A(n_1485),
.B(n_1489),
.Y(n_1519)
);

HB1xp67_ASAP7_75t_L g1520 ( 
.A(n_1481),
.Y(n_1520)
);

AND2x2_ASAP7_75t_L g1521 ( 
.A(n_1489),
.B(n_1459),
.Y(n_1521)
);

AOI22xp33_ASAP7_75t_L g1522 ( 
.A1(n_1488),
.A2(n_1470),
.B1(n_1462),
.B2(n_1457),
.Y(n_1522)
);

NAND4xp25_ASAP7_75t_SL g1523 ( 
.A(n_1484),
.B(n_1396),
.C(n_1446),
.D(n_1467),
.Y(n_1523)
);

NAND2xp5_ASAP7_75t_L g1524 ( 
.A(n_1494),
.B(n_1465),
.Y(n_1524)
);

AOI221xp5_ASAP7_75t_L g1525 ( 
.A1(n_1483),
.A2(n_1434),
.B1(n_1468),
.B2(n_1471),
.C(n_1465),
.Y(n_1525)
);

OAI22xp5_ASAP7_75t_L g1526 ( 
.A1(n_1484),
.A2(n_1457),
.B1(n_1445),
.B2(n_1464),
.Y(n_1526)
);

OR2x6_ASAP7_75t_L g1527 ( 
.A(n_1479),
.B(n_1436),
.Y(n_1527)
);

INVx1_ASAP7_75t_L g1528 ( 
.A(n_1475),
.Y(n_1528)
);

AND2x2_ASAP7_75t_L g1529 ( 
.A(n_1489),
.B(n_1455),
.Y(n_1529)
);

OAI31xp33_ASAP7_75t_L g1530 ( 
.A1(n_1477),
.A2(n_1366),
.A3(n_1467),
.B(n_1493),
.Y(n_1530)
);

OA21x2_ASAP7_75t_L g1531 ( 
.A1(n_1512),
.A2(n_1525),
.B(n_1452),
.Y(n_1531)
);

HB1xp67_ASAP7_75t_L g1532 ( 
.A(n_1506),
.Y(n_1532)
);

INVx1_ASAP7_75t_L g1533 ( 
.A(n_1504),
.Y(n_1533)
);

INVx1_ASAP7_75t_SL g1534 ( 
.A(n_1499),
.Y(n_1534)
);

INVx1_ASAP7_75t_SL g1535 ( 
.A(n_1495),
.Y(n_1535)
);

OAI21xp5_ASAP7_75t_L g1536 ( 
.A1(n_1507),
.A2(n_1480),
.B(n_1494),
.Y(n_1536)
);

INVx1_ASAP7_75t_L g1537 ( 
.A(n_1504),
.Y(n_1537)
);

INVx1_ASAP7_75t_L g1538 ( 
.A(n_1508),
.Y(n_1538)
);

BUFx2_ASAP7_75t_L g1539 ( 
.A(n_1497),
.Y(n_1539)
);

INVx1_ASAP7_75t_L g1540 ( 
.A(n_1508),
.Y(n_1540)
);

INVx1_ASAP7_75t_L g1541 ( 
.A(n_1528),
.Y(n_1541)
);

AND2x4_ASAP7_75t_L g1542 ( 
.A(n_1497),
.B(n_1479),
.Y(n_1542)
);

AND4x1_ASAP7_75t_L g1543 ( 
.A(n_1502),
.B(n_1362),
.C(n_1441),
.D(n_1456),
.Y(n_1543)
);

OA21x2_ASAP7_75t_L g1544 ( 
.A1(n_1517),
.A2(n_1453),
.B(n_1451),
.Y(n_1544)
);

INVx1_ASAP7_75t_L g1545 ( 
.A(n_1520),
.Y(n_1545)
);

INVx1_ASAP7_75t_SL g1546 ( 
.A(n_1495),
.Y(n_1546)
);

AND2x2_ASAP7_75t_L g1547 ( 
.A(n_1519),
.B(n_1486),
.Y(n_1547)
);

NAND2xp5_ASAP7_75t_L g1548 ( 
.A(n_1496),
.B(n_1486),
.Y(n_1548)
);

AND2x2_ASAP7_75t_L g1549 ( 
.A(n_1519),
.B(n_1486),
.Y(n_1549)
);

AND2x2_ASAP7_75t_L g1550 ( 
.A(n_1509),
.B(n_1501),
.Y(n_1550)
);

NOR3xp33_ASAP7_75t_L g1551 ( 
.A(n_1507),
.B(n_1395),
.C(n_1416),
.Y(n_1551)
);

INVxp67_ASAP7_75t_L g1552 ( 
.A(n_1509),
.Y(n_1552)
);

NAND2xp5_ASAP7_75t_L g1553 ( 
.A(n_1524),
.B(n_1492),
.Y(n_1553)
);

INVxp67_ASAP7_75t_L g1554 ( 
.A(n_1516),
.Y(n_1554)
);

NAND2xp5_ASAP7_75t_L g1555 ( 
.A(n_1500),
.B(n_1492),
.Y(n_1555)
);

INVx1_ASAP7_75t_L g1556 ( 
.A(n_1533),
.Y(n_1556)
);

NAND2xp5_ASAP7_75t_L g1557 ( 
.A(n_1534),
.B(n_1500),
.Y(n_1557)
);

NAND2x1p5_ASAP7_75t_L g1558 ( 
.A(n_1550),
.B(n_1477),
.Y(n_1558)
);

AND2x2_ASAP7_75t_L g1559 ( 
.A(n_1550),
.B(n_1501),
.Y(n_1559)
);

AND2x2_ASAP7_75t_L g1560 ( 
.A(n_1550),
.B(n_1511),
.Y(n_1560)
);

AND2x2_ASAP7_75t_L g1561 ( 
.A(n_1552),
.B(n_1511),
.Y(n_1561)
);

AND2x2_ASAP7_75t_L g1562 ( 
.A(n_1552),
.B(n_1539),
.Y(n_1562)
);

NAND2x1p5_ASAP7_75t_L g1563 ( 
.A(n_1535),
.B(n_1503),
.Y(n_1563)
);

NAND2xp5_ASAP7_75t_L g1564 ( 
.A(n_1534),
.B(n_1513),
.Y(n_1564)
);

HB1xp67_ASAP7_75t_L g1565 ( 
.A(n_1532),
.Y(n_1565)
);

INVx1_ASAP7_75t_L g1566 ( 
.A(n_1533),
.Y(n_1566)
);

INVx1_ASAP7_75t_L g1567 ( 
.A(n_1537),
.Y(n_1567)
);

AND2x4_ASAP7_75t_L g1568 ( 
.A(n_1539),
.B(n_1497),
.Y(n_1568)
);

INVx1_ASAP7_75t_L g1569 ( 
.A(n_1537),
.Y(n_1569)
);

INVx1_ASAP7_75t_L g1570 ( 
.A(n_1538),
.Y(n_1570)
);

AND3x2_ASAP7_75t_L g1571 ( 
.A(n_1554),
.B(n_1503),
.C(n_1530),
.Y(n_1571)
);

AND2x2_ASAP7_75t_L g1572 ( 
.A(n_1539),
.B(n_1554),
.Y(n_1572)
);

AND2x4_ASAP7_75t_L g1573 ( 
.A(n_1542),
.B(n_1497),
.Y(n_1573)
);

NAND2xp5_ASAP7_75t_L g1574 ( 
.A(n_1536),
.B(n_1551),
.Y(n_1574)
);

INVx2_ASAP7_75t_L g1575 ( 
.A(n_1547),
.Y(n_1575)
);

NAND2xp5_ASAP7_75t_L g1576 ( 
.A(n_1536),
.B(n_1513),
.Y(n_1576)
);

NAND2xp5_ASAP7_75t_SL g1577 ( 
.A(n_1543),
.B(n_1530),
.Y(n_1577)
);

AOI21xp5_ASAP7_75t_L g1578 ( 
.A1(n_1531),
.A2(n_1498),
.B(n_1505),
.Y(n_1578)
);

OR2x2_ASAP7_75t_L g1579 ( 
.A(n_1555),
.B(n_1515),
.Y(n_1579)
);

NAND2xp5_ASAP7_75t_L g1580 ( 
.A(n_1551),
.B(n_1487),
.Y(n_1580)
);

INVx1_ASAP7_75t_L g1581 ( 
.A(n_1540),
.Y(n_1581)
);

AND2x2_ASAP7_75t_L g1582 ( 
.A(n_1547),
.B(n_1529),
.Y(n_1582)
);

INVxp33_ASAP7_75t_L g1583 ( 
.A(n_1548),
.Y(n_1583)
);

AND2x4_ASAP7_75t_L g1584 ( 
.A(n_1542),
.B(n_1497),
.Y(n_1584)
);

AND2x2_ASAP7_75t_L g1585 ( 
.A(n_1547),
.B(n_1529),
.Y(n_1585)
);

INVx4_ASAP7_75t_L g1586 ( 
.A(n_1532),
.Y(n_1586)
);

AOI21xp5_ASAP7_75t_L g1587 ( 
.A1(n_1531),
.A2(n_1523),
.B(n_1518),
.Y(n_1587)
);

CKINVDCx14_ASAP7_75t_R g1588 ( 
.A(n_1545),
.Y(n_1588)
);

INVx2_ASAP7_75t_L g1589 ( 
.A(n_1549),
.Y(n_1589)
);

AND2x2_ASAP7_75t_SL g1590 ( 
.A(n_1574),
.B(n_1543),
.Y(n_1590)
);

NAND2xp5_ASAP7_75t_L g1591 ( 
.A(n_1557),
.B(n_1545),
.Y(n_1591)
);

AND2x2_ASAP7_75t_L g1592 ( 
.A(n_1558),
.B(n_1535),
.Y(n_1592)
);

INVx2_ASAP7_75t_L g1593 ( 
.A(n_1563),
.Y(n_1593)
);

AND2x2_ASAP7_75t_L g1594 ( 
.A(n_1558),
.B(n_1559),
.Y(n_1594)
);

NAND2xp5_ASAP7_75t_L g1595 ( 
.A(n_1578),
.B(n_1546),
.Y(n_1595)
);

BUFx12f_ASAP7_75t_L g1596 ( 
.A(n_1586),
.Y(n_1596)
);

AND2x2_ASAP7_75t_L g1597 ( 
.A(n_1558),
.B(n_1546),
.Y(n_1597)
);

OR2x2_ASAP7_75t_L g1598 ( 
.A(n_1564),
.B(n_1565),
.Y(n_1598)
);

NOR2xp33_ASAP7_75t_L g1599 ( 
.A(n_1588),
.B(n_1362),
.Y(n_1599)
);

NAND3xp33_ASAP7_75t_SL g1600 ( 
.A(n_1587),
.B(n_1510),
.C(n_1522),
.Y(n_1600)
);

OAI22xp33_ASAP7_75t_L g1601 ( 
.A1(n_1577),
.A2(n_1514),
.B1(n_1531),
.B2(n_1526),
.Y(n_1601)
);

AOI21xp33_ASAP7_75t_SL g1602 ( 
.A1(n_1563),
.A2(n_1423),
.B(n_1531),
.Y(n_1602)
);

NAND2xp5_ASAP7_75t_L g1603 ( 
.A(n_1572),
.B(n_1548),
.Y(n_1603)
);

INVx1_ASAP7_75t_L g1604 ( 
.A(n_1556),
.Y(n_1604)
);

AOI21xp33_ASAP7_75t_L g1605 ( 
.A1(n_1562),
.A2(n_1531),
.B(n_1434),
.Y(n_1605)
);

NAND2xp5_ASAP7_75t_SL g1606 ( 
.A(n_1580),
.B(n_1542),
.Y(n_1606)
);

INVx1_ASAP7_75t_L g1607 ( 
.A(n_1556),
.Y(n_1607)
);

NAND2xp5_ASAP7_75t_L g1608 ( 
.A(n_1572),
.B(n_1553),
.Y(n_1608)
);

NAND2xp5_ASAP7_75t_L g1609 ( 
.A(n_1562),
.B(n_1553),
.Y(n_1609)
);

INVx1_ASAP7_75t_SL g1610 ( 
.A(n_1571),
.Y(n_1610)
);

BUFx3_ASAP7_75t_L g1611 ( 
.A(n_1563),
.Y(n_1611)
);

AND2x2_ASAP7_75t_L g1612 ( 
.A(n_1559),
.B(n_1542),
.Y(n_1612)
);

AOI22xp5_ASAP7_75t_L g1613 ( 
.A1(n_1576),
.A2(n_1435),
.B1(n_1544),
.B2(n_1490),
.Y(n_1613)
);

NAND2xp5_ASAP7_75t_L g1614 ( 
.A(n_1561),
.B(n_1521),
.Y(n_1614)
);

INVx1_ASAP7_75t_SL g1615 ( 
.A(n_1586),
.Y(n_1615)
);

AND2x4_ASAP7_75t_L g1616 ( 
.A(n_1560),
.B(n_1541),
.Y(n_1616)
);

AND2x2_ASAP7_75t_L g1617 ( 
.A(n_1560),
.B(n_1527),
.Y(n_1617)
);

INVx2_ASAP7_75t_L g1618 ( 
.A(n_1586),
.Y(n_1618)
);

AOI22xp33_ASAP7_75t_L g1619 ( 
.A1(n_1583),
.A2(n_1474),
.B1(n_1436),
.B2(n_1469),
.Y(n_1619)
);

INVx2_ASAP7_75t_L g1620 ( 
.A(n_1586),
.Y(n_1620)
);

AND2x2_ASAP7_75t_L g1621 ( 
.A(n_1561),
.B(n_1527),
.Y(n_1621)
);

NOR2xp33_ASAP7_75t_L g1622 ( 
.A(n_1579),
.B(n_1423),
.Y(n_1622)
);

INVx1_ASAP7_75t_L g1623 ( 
.A(n_1566),
.Y(n_1623)
);

NOR2xp33_ASAP7_75t_L g1624 ( 
.A(n_1599),
.B(n_1579),
.Y(n_1624)
);

NAND2xp5_ASAP7_75t_L g1625 ( 
.A(n_1590),
.B(n_1566),
.Y(n_1625)
);

NOR2xp33_ASAP7_75t_L g1626 ( 
.A(n_1590),
.B(n_1416),
.Y(n_1626)
);

AND2x2_ASAP7_75t_L g1627 ( 
.A(n_1594),
.B(n_1582),
.Y(n_1627)
);

INVx1_ASAP7_75t_L g1628 ( 
.A(n_1604),
.Y(n_1628)
);

OR2x2_ASAP7_75t_L g1629 ( 
.A(n_1598),
.B(n_1575),
.Y(n_1629)
);

AND2x2_ASAP7_75t_L g1630 ( 
.A(n_1594),
.B(n_1582),
.Y(n_1630)
);

AOI22xp33_ASAP7_75t_L g1631 ( 
.A1(n_1590),
.A2(n_1568),
.B1(n_1573),
.B2(n_1584),
.Y(n_1631)
);

INVx1_ASAP7_75t_SL g1632 ( 
.A(n_1610),
.Y(n_1632)
);

HB1xp67_ASAP7_75t_L g1633 ( 
.A(n_1615),
.Y(n_1633)
);

AND2x2_ASAP7_75t_L g1634 ( 
.A(n_1592),
.B(n_1585),
.Y(n_1634)
);

INVx1_ASAP7_75t_SL g1635 ( 
.A(n_1611),
.Y(n_1635)
);

AND2x2_ASAP7_75t_L g1636 ( 
.A(n_1592),
.B(n_1585),
.Y(n_1636)
);

INVx2_ASAP7_75t_L g1637 ( 
.A(n_1611),
.Y(n_1637)
);

AOI22xp33_ASAP7_75t_L g1638 ( 
.A1(n_1600),
.A2(n_1568),
.B1(n_1573),
.B2(n_1584),
.Y(n_1638)
);

INVxp67_ASAP7_75t_L g1639 ( 
.A(n_1622),
.Y(n_1639)
);

INVx2_ASAP7_75t_L g1640 ( 
.A(n_1611),
.Y(n_1640)
);

BUFx3_ASAP7_75t_L g1641 ( 
.A(n_1596),
.Y(n_1641)
);

OAI22xp5_ASAP7_75t_L g1642 ( 
.A1(n_1601),
.A2(n_1575),
.B1(n_1589),
.B2(n_1568),
.Y(n_1642)
);

INVx1_ASAP7_75t_L g1643 ( 
.A(n_1604),
.Y(n_1643)
);

INVx1_ASAP7_75t_SL g1644 ( 
.A(n_1615),
.Y(n_1644)
);

OR2x2_ASAP7_75t_L g1645 ( 
.A(n_1598),
.B(n_1589),
.Y(n_1645)
);

AND2x4_ASAP7_75t_L g1646 ( 
.A(n_1597),
.B(n_1568),
.Y(n_1646)
);

INVx1_ASAP7_75t_L g1647 ( 
.A(n_1623),
.Y(n_1647)
);

INVxp67_ASAP7_75t_L g1648 ( 
.A(n_1618),
.Y(n_1648)
);

INVx1_ASAP7_75t_L g1649 ( 
.A(n_1633),
.Y(n_1649)
);

NAND2xp5_ASAP7_75t_L g1650 ( 
.A(n_1632),
.B(n_1595),
.Y(n_1650)
);

AOI21xp5_ASAP7_75t_L g1651 ( 
.A1(n_1642),
.A2(n_1591),
.B(n_1602),
.Y(n_1651)
);

INVx1_ASAP7_75t_L g1652 ( 
.A(n_1628),
.Y(n_1652)
);

INVx1_ASAP7_75t_L g1653 ( 
.A(n_1628),
.Y(n_1653)
);

NAND2xp5_ASAP7_75t_SL g1654 ( 
.A(n_1632),
.B(n_1602),
.Y(n_1654)
);

NAND2xp5_ASAP7_75t_L g1655 ( 
.A(n_1635),
.B(n_1603),
.Y(n_1655)
);

AOI21xp5_ASAP7_75t_SL g1656 ( 
.A1(n_1626),
.A2(n_1620),
.B(n_1618),
.Y(n_1656)
);

NAND2xp5_ASAP7_75t_L g1657 ( 
.A(n_1635),
.B(n_1618),
.Y(n_1657)
);

OAI211xp5_ASAP7_75t_L g1658 ( 
.A1(n_1638),
.A2(n_1625),
.B(n_1642),
.C(n_1631),
.Y(n_1658)
);

OR2x6_ASAP7_75t_L g1659 ( 
.A(n_1641),
.B(n_1639),
.Y(n_1659)
);

AO221x1_ASAP7_75t_L g1660 ( 
.A1(n_1648),
.A2(n_1593),
.B1(n_1620),
.B2(n_1623),
.C(n_1607),
.Y(n_1660)
);

INVxp67_ASAP7_75t_L g1661 ( 
.A(n_1624),
.Y(n_1661)
);

NAND2xp5_ASAP7_75t_L g1662 ( 
.A(n_1644),
.B(n_1620),
.Y(n_1662)
);

AOI21xp33_ASAP7_75t_L g1663 ( 
.A1(n_1625),
.A2(n_1596),
.B(n_1593),
.Y(n_1663)
);

INVx1_ASAP7_75t_L g1664 ( 
.A(n_1643),
.Y(n_1664)
);

OR2x6_ASAP7_75t_L g1665 ( 
.A(n_1641),
.B(n_1596),
.Y(n_1665)
);

AOI22xp33_ASAP7_75t_SL g1666 ( 
.A1(n_1627),
.A2(n_1597),
.B1(n_1608),
.B2(n_1609),
.Y(n_1666)
);

NAND2xp5_ASAP7_75t_L g1667 ( 
.A(n_1644),
.B(n_1614),
.Y(n_1667)
);

AND2x2_ASAP7_75t_L g1668 ( 
.A(n_1659),
.B(n_1646),
.Y(n_1668)
);

OR2x2_ASAP7_75t_L g1669 ( 
.A(n_1650),
.B(n_1629),
.Y(n_1669)
);

NAND2xp5_ASAP7_75t_L g1670 ( 
.A(n_1649),
.B(n_1637),
.Y(n_1670)
);

INVx1_ASAP7_75t_L g1671 ( 
.A(n_1662),
.Y(n_1671)
);

NAND2xp5_ASAP7_75t_SL g1672 ( 
.A(n_1651),
.B(n_1637),
.Y(n_1672)
);

AND2x2_ASAP7_75t_L g1673 ( 
.A(n_1659),
.B(n_1646),
.Y(n_1673)
);

INVx2_ASAP7_75t_L g1674 ( 
.A(n_1660),
.Y(n_1674)
);

INVxp33_ASAP7_75t_L g1675 ( 
.A(n_1656),
.Y(n_1675)
);

AND2x2_ASAP7_75t_L g1676 ( 
.A(n_1666),
.B(n_1646),
.Y(n_1676)
);

AOI22xp33_ASAP7_75t_L g1677 ( 
.A1(n_1654),
.A2(n_1641),
.B1(n_1605),
.B2(n_1646),
.Y(n_1677)
);

INVx2_ASAP7_75t_L g1678 ( 
.A(n_1665),
.Y(n_1678)
);

INVx1_ASAP7_75t_L g1679 ( 
.A(n_1670),
.Y(n_1679)
);

AOI211xp5_ASAP7_75t_L g1680 ( 
.A1(n_1675),
.A2(n_1658),
.B(n_1663),
.C(n_1661),
.Y(n_1680)
);

OAI221xp5_ASAP7_75t_SL g1681 ( 
.A1(n_1677),
.A2(n_1665),
.B1(n_1667),
.B2(n_1655),
.C(n_1657),
.Y(n_1681)
);

OAI211xp5_ASAP7_75t_SL g1682 ( 
.A1(n_1672),
.A2(n_1637),
.B(n_1640),
.C(n_1648),
.Y(n_1682)
);

AOI21xp33_ASAP7_75t_L g1683 ( 
.A1(n_1675),
.A2(n_1640),
.B(n_1629),
.Y(n_1683)
);

NAND2xp33_ASAP7_75t_R g1684 ( 
.A(n_1668),
.B(n_1640),
.Y(n_1684)
);

A2O1A1Ixp33_ASAP7_75t_L g1685 ( 
.A1(n_1674),
.A2(n_1613),
.B(n_1664),
.C(n_1652),
.Y(n_1685)
);

OAI22xp5_ASAP7_75t_L g1686 ( 
.A1(n_1674),
.A2(n_1606),
.B1(n_1619),
.B2(n_1630),
.Y(n_1686)
);

NOR2xp33_ASAP7_75t_SL g1687 ( 
.A(n_1668),
.B(n_1673),
.Y(n_1687)
);

NAND2xp5_ASAP7_75t_SL g1688 ( 
.A(n_1669),
.B(n_1645),
.Y(n_1688)
);

NOR2xp33_ASAP7_75t_SL g1689 ( 
.A(n_1676),
.B(n_1678),
.Y(n_1689)
);

INVx1_ASAP7_75t_L g1690 ( 
.A(n_1688),
.Y(n_1690)
);

INVx1_ASAP7_75t_L g1691 ( 
.A(n_1679),
.Y(n_1691)
);

AOI221xp5_ASAP7_75t_L g1692 ( 
.A1(n_1681),
.A2(n_1672),
.B1(n_1671),
.B2(n_1678),
.C(n_1653),
.Y(n_1692)
);

AO22x1_ASAP7_75t_L g1693 ( 
.A1(n_1686),
.A2(n_1593),
.B1(n_1643),
.B2(n_1647),
.Y(n_1693)
);

OR2x2_ASAP7_75t_L g1694 ( 
.A(n_1685),
.B(n_1645),
.Y(n_1694)
);

NOR2x1_ASAP7_75t_L g1695 ( 
.A(n_1690),
.B(n_1682),
.Y(n_1695)
);

INVx1_ASAP7_75t_L g1696 ( 
.A(n_1694),
.Y(n_1696)
);

INVx1_ASAP7_75t_L g1697 ( 
.A(n_1691),
.Y(n_1697)
);

NAND2xp5_ASAP7_75t_L g1698 ( 
.A(n_1693),
.B(n_1689),
.Y(n_1698)
);

INVx3_ASAP7_75t_SL g1699 ( 
.A(n_1692),
.Y(n_1699)
);

AOI21xp5_ASAP7_75t_L g1700 ( 
.A1(n_1693),
.A2(n_1680),
.B(n_1687),
.Y(n_1700)
);

INVx2_ASAP7_75t_L g1701 ( 
.A(n_1698),
.Y(n_1701)
);

OAI211xp5_ASAP7_75t_L g1702 ( 
.A1(n_1695),
.A2(n_1683),
.B(n_1684),
.C(n_1647),
.Y(n_1702)
);

NAND2xp5_ASAP7_75t_L g1703 ( 
.A(n_1699),
.B(n_1607),
.Y(n_1703)
);

INVx1_ASAP7_75t_L g1704 ( 
.A(n_1696),
.Y(n_1704)
);

INVx1_ASAP7_75t_L g1705 ( 
.A(n_1697),
.Y(n_1705)
);

BUFx2_ASAP7_75t_L g1706 ( 
.A(n_1704),
.Y(n_1706)
);

AOI322xp5_ASAP7_75t_L g1707 ( 
.A1(n_1703),
.A2(n_1700),
.A3(n_1636),
.B1(n_1634),
.B2(n_1613),
.C1(n_1630),
.C2(n_1627),
.Y(n_1707)
);

CKINVDCx6p67_ASAP7_75t_R g1708 ( 
.A(n_1705),
.Y(n_1708)
);

BUFx2_ASAP7_75t_L g1709 ( 
.A(n_1706),
.Y(n_1709)
);

OAI221xp5_ASAP7_75t_SL g1710 ( 
.A1(n_1709),
.A2(n_1707),
.B1(n_1702),
.B2(n_1703),
.C(n_1701),
.Y(n_1710)
);

BUFx2_ASAP7_75t_L g1711 ( 
.A(n_1710),
.Y(n_1711)
);

OAI21xp5_ASAP7_75t_L g1712 ( 
.A1(n_1711),
.A2(n_1708),
.B(n_1636),
.Y(n_1712)
);

BUFx2_ASAP7_75t_L g1713 ( 
.A(n_1712),
.Y(n_1713)
);

INVx1_ASAP7_75t_L g1714 ( 
.A(n_1713),
.Y(n_1714)
);

OAI22x1_ASAP7_75t_L g1715 ( 
.A1(n_1713),
.A2(n_1634),
.B1(n_1616),
.B2(n_1612),
.Y(n_1715)
);

NOR2xp67_ASAP7_75t_L g1716 ( 
.A(n_1714),
.B(n_1616),
.Y(n_1716)
);

AOI21xp5_ASAP7_75t_L g1717 ( 
.A1(n_1715),
.A2(n_1616),
.B(n_1621),
.Y(n_1717)
);

INVx1_ASAP7_75t_L g1718 ( 
.A(n_1716),
.Y(n_1718)
);

NAND2x1_ASAP7_75t_L g1719 ( 
.A(n_1717),
.B(n_1616),
.Y(n_1719)
);

AOI322xp5_ASAP7_75t_L g1720 ( 
.A1(n_1719),
.A2(n_1718),
.A3(n_1621),
.B1(n_1612),
.B2(n_1617),
.C1(n_1584),
.C2(n_1573),
.Y(n_1720)
);

INVxp67_ASAP7_75t_L g1721 ( 
.A(n_1718),
.Y(n_1721)
);

AOI22xp5_ASAP7_75t_L g1722 ( 
.A1(n_1721),
.A2(n_1720),
.B1(n_1617),
.B2(n_1570),
.Y(n_1722)
);

AOI211xp5_ASAP7_75t_L g1723 ( 
.A1(n_1722),
.A2(n_1581),
.B(n_1567),
.C(n_1569),
.Y(n_1723)
);


endmodule