module fake_jpeg_25749_n_340 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_340);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_340;

wire n_253;
wire n_330;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVx4_ASAP7_75t_L g16 ( 
.A(n_1),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_14),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_9),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_1),
.Y(n_19)
);

BUFx24_ASAP7_75t_L g20 ( 
.A(n_12),
.Y(n_20)
);

NOR2xp33_ASAP7_75t_L g21 ( 
.A(n_5),
.B(n_15),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_8),
.Y(n_22)
);

INVx8_ASAP7_75t_L g23 ( 
.A(n_6),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_1),
.Y(n_24)
);

INVx8_ASAP7_75t_L g25 ( 
.A(n_4),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_11),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_2),
.Y(n_27)
);

INVx3_ASAP7_75t_L g28 ( 
.A(n_13),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_11),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_14),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_1),
.Y(n_31)
);

INVx8_ASAP7_75t_L g32 ( 
.A(n_10),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_9),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_10),
.Y(n_34)
);

BUFx5_ASAP7_75t_L g35 ( 
.A(n_12),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_20),
.Y(n_36)
);

CKINVDCx6p67_ASAP7_75t_R g60 ( 
.A(n_36),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_20),
.Y(n_37)
);

INVx2_ASAP7_75t_L g67 ( 
.A(n_37),
.Y(n_67)
);

INVx3_ASAP7_75t_L g38 ( 
.A(n_23),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_38),
.Y(n_50)
);

BUFx5_ASAP7_75t_L g39 ( 
.A(n_20),
.Y(n_39)
);

BUFx2_ASAP7_75t_L g73 ( 
.A(n_39),
.Y(n_73)
);

INVx5_ASAP7_75t_L g40 ( 
.A(n_23),
.Y(n_40)
);

INVx4_ASAP7_75t_L g56 ( 
.A(n_40),
.Y(n_56)
);

INVx6_ASAP7_75t_L g41 ( 
.A(n_30),
.Y(n_41)
);

INVx3_ASAP7_75t_L g53 ( 
.A(n_41),
.Y(n_53)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_17),
.Y(n_42)
);

NAND2xp5_ASAP7_75t_L g55 ( 
.A(n_42),
.B(n_19),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_20),
.Y(n_43)
);

INVx2_ASAP7_75t_L g51 ( 
.A(n_43),
.Y(n_51)
);

INVx4_ASAP7_75t_L g44 ( 
.A(n_30),
.Y(n_44)
);

INVx2_ASAP7_75t_L g54 ( 
.A(n_44),
.Y(n_54)
);

INVx4_ASAP7_75t_L g45 ( 
.A(n_30),
.Y(n_45)
);

INVx2_ASAP7_75t_L g72 ( 
.A(n_45),
.Y(n_72)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_20),
.Y(n_46)
);

INVx4_ASAP7_75t_L g68 ( 
.A(n_46),
.Y(n_68)
);

INVx2_ASAP7_75t_L g47 ( 
.A(n_16),
.Y(n_47)
);

BUFx3_ASAP7_75t_L g69 ( 
.A(n_47),
.Y(n_69)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_20),
.Y(n_48)
);

INVx3_ASAP7_75t_L g59 ( 
.A(n_48),
.Y(n_59)
);

AOI22xp33_ASAP7_75t_SL g49 ( 
.A1(n_16),
.A2(n_0),
.B1(n_2),
.B2(n_3),
.Y(n_49)
);

OAI22xp5_ASAP7_75t_L g65 ( 
.A1(n_49),
.A2(n_17),
.B1(n_19),
.B2(n_22),
.Y(n_65)
);

INVx5_ASAP7_75t_L g52 ( 
.A(n_39),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g79 ( 
.A(n_52),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_SL g84 ( 
.A(n_55),
.B(n_57),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_SL g57 ( 
.A(n_42),
.B(n_21),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_42),
.B(n_21),
.Y(n_58)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_58),
.Y(n_76)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_47),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_61),
.B(n_62),
.Y(n_101)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_47),
.Y(n_62)
);

OAI22xp33_ASAP7_75t_L g63 ( 
.A1(n_41),
.A2(n_16),
.B1(n_28),
.B2(n_32),
.Y(n_63)
);

OAI22xp5_ASAP7_75t_SL g107 ( 
.A1(n_63),
.A2(n_64),
.B1(n_45),
.B2(n_44),
.Y(n_107)
);

AOI22xp5_ASAP7_75t_L g64 ( 
.A1(n_41),
.A2(n_28),
.B1(n_16),
.B2(n_25),
.Y(n_64)
);

AOI22xp5_ASAP7_75t_L g80 ( 
.A1(n_65),
.A2(n_26),
.B1(n_29),
.B2(n_31),
.Y(n_80)
);

HB1xp67_ASAP7_75t_L g66 ( 
.A(n_38),
.Y(n_66)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_66),
.Y(n_77)
);

INVx3_ASAP7_75t_L g70 ( 
.A(n_36),
.Y(n_70)
);

INVx6_ASAP7_75t_L g112 ( 
.A(n_70),
.Y(n_112)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_44),
.Y(n_71)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_71),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_L g74 ( 
.A(n_49),
.B(n_27),
.Y(n_74)
);

AND2x2_ASAP7_75t_L g100 ( 
.A(n_74),
.B(n_34),
.Y(n_100)
);

INVx4_ASAP7_75t_SL g75 ( 
.A(n_39),
.Y(n_75)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_75),
.Y(n_98)
);

NOR2x1_ASAP7_75t_SL g78 ( 
.A(n_63),
.B(n_35),
.Y(n_78)
);

NAND2xp33_ASAP7_75t_SL g143 ( 
.A(n_78),
.B(n_35),
.Y(n_143)
);

OAI22xp5_ASAP7_75t_SL g116 ( 
.A1(n_80),
.A2(n_18),
.B1(n_33),
.B2(n_31),
.Y(n_116)
);

CKINVDCx20_ASAP7_75t_R g81 ( 
.A(n_73),
.Y(n_81)
);

OR2x2_ASAP7_75t_L g117 ( 
.A(n_81),
.B(n_37),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_L g82 ( 
.A(n_69),
.B(n_17),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_L g120 ( 
.A(n_82),
.B(n_95),
.Y(n_120)
);

INVx2_ASAP7_75t_L g83 ( 
.A(n_69),
.Y(n_83)
);

INVx2_ASAP7_75t_L g125 ( 
.A(n_83),
.Y(n_125)
);

INVx4_ASAP7_75t_L g85 ( 
.A(n_50),
.Y(n_85)
);

INVx2_ASAP7_75t_L g129 ( 
.A(n_85),
.Y(n_129)
);

AOI22xp33_ASAP7_75t_SL g86 ( 
.A1(n_52),
.A2(n_28),
.B1(n_25),
.B2(n_23),
.Y(n_86)
);

OAI22xp5_ASAP7_75t_L g141 ( 
.A1(n_86),
.A2(n_89),
.B1(n_99),
.B2(n_106),
.Y(n_141)
);

BUFx6f_ASAP7_75t_L g87 ( 
.A(n_59),
.Y(n_87)
);

BUFx6f_ASAP7_75t_L g146 ( 
.A(n_87),
.Y(n_146)
);

INVx2_ASAP7_75t_L g88 ( 
.A(n_54),
.Y(n_88)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_88),
.Y(n_118)
);

AOI22xp33_ASAP7_75t_SL g89 ( 
.A1(n_56),
.A2(n_25),
.B1(n_32),
.B2(n_23),
.Y(n_89)
);

INVx5_ASAP7_75t_L g90 ( 
.A(n_60),
.Y(n_90)
);

AOI22xp33_ASAP7_75t_SL g134 ( 
.A1(n_90),
.A2(n_96),
.B1(n_113),
.B2(n_48),
.Y(n_134)
);

INVx4_ASAP7_75t_L g91 ( 
.A(n_50),
.Y(n_91)
);

INVx3_ASAP7_75t_L g124 ( 
.A(n_91),
.Y(n_124)
);

INVx2_ASAP7_75t_L g92 ( 
.A(n_54),
.Y(n_92)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_92),
.Y(n_121)
);

INVx4_ASAP7_75t_L g94 ( 
.A(n_60),
.Y(n_94)
);

INVx3_ASAP7_75t_L g138 ( 
.A(n_94),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_L g95 ( 
.A(n_72),
.B(n_19),
.Y(n_95)
);

INVx5_ASAP7_75t_L g96 ( 
.A(n_60),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g97 ( 
.A(n_72),
.B(n_22),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_97),
.B(n_18),
.Y(n_127)
);

AOI22xp33_ASAP7_75t_SL g99 ( 
.A1(n_56),
.A2(n_32),
.B1(n_25),
.B2(n_22),
.Y(n_99)
);

OAI21xp5_ASAP7_75t_SL g131 ( 
.A1(n_100),
.A2(n_109),
.B(n_24),
.Y(n_131)
);

INVx3_ASAP7_75t_L g102 ( 
.A(n_60),
.Y(n_102)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_102),
.Y(n_128)
);

INVx3_ASAP7_75t_L g103 ( 
.A(n_73),
.Y(n_103)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_103),
.Y(n_130)
);

INVx2_ASAP7_75t_L g104 ( 
.A(n_51),
.Y(n_104)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_104),
.Y(n_136)
);

INVx2_ASAP7_75t_L g105 ( 
.A(n_51),
.Y(n_105)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_105),
.Y(n_139)
);

AOI22xp33_ASAP7_75t_SL g106 ( 
.A1(n_75),
.A2(n_32),
.B1(n_27),
.B2(n_41),
.Y(n_106)
);

AOI22xp5_ASAP7_75t_L g133 ( 
.A1(n_107),
.A2(n_115),
.B1(n_94),
.B2(n_102),
.Y(n_133)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_64),
.Y(n_108)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_108),
.Y(n_140)
);

AOI22xp5_ASAP7_75t_SL g109 ( 
.A1(n_53),
.A2(n_26),
.B1(n_18),
.B2(n_24),
.Y(n_109)
);

INVx2_ASAP7_75t_L g110 ( 
.A(n_67),
.Y(n_110)
);

BUFx5_ASAP7_75t_L g144 ( 
.A(n_110),
.Y(n_144)
);

AOI22xp33_ASAP7_75t_SL g111 ( 
.A1(n_53),
.A2(n_27),
.B1(n_40),
.B2(n_44),
.Y(n_111)
);

OAI22xp5_ASAP7_75t_L g145 ( 
.A1(n_111),
.A2(n_114),
.B1(n_48),
.B2(n_46),
.Y(n_145)
);

INVx2_ASAP7_75t_L g113 ( 
.A(n_68),
.Y(n_113)
);

AOI22xp33_ASAP7_75t_SL g114 ( 
.A1(n_68),
.A2(n_40),
.B1(n_45),
.B2(n_38),
.Y(n_114)
);

OAI22xp5_ASAP7_75t_SL g115 ( 
.A1(n_59),
.A2(n_45),
.B1(n_38),
.B2(n_40),
.Y(n_115)
);

AOI22xp5_ASAP7_75t_L g155 ( 
.A1(n_116),
.A2(n_119),
.B1(n_132),
.B2(n_123),
.Y(n_155)
);

CKINVDCx16_ASAP7_75t_R g158 ( 
.A(n_117),
.Y(n_158)
);

OAI22xp5_ASAP7_75t_SL g119 ( 
.A1(n_78),
.A2(n_80),
.B1(n_100),
.B2(n_107),
.Y(n_119)
);

NAND3xp33_ASAP7_75t_L g122 ( 
.A(n_84),
.B(n_15),
.C(n_2),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_SL g176 ( 
.A(n_122),
.B(n_0),
.Y(n_176)
);

AND2x2_ASAP7_75t_L g123 ( 
.A(n_95),
.B(n_36),
.Y(n_123)
);

OAI21xp5_ASAP7_75t_SL g150 ( 
.A1(n_123),
.A2(n_131),
.B(n_93),
.Y(n_150)
);

MAJIxp5_ASAP7_75t_L g126 ( 
.A(n_100),
.B(n_37),
.C(n_48),
.Y(n_126)
);

MAJIxp5_ASAP7_75t_L g160 ( 
.A(n_126),
.B(n_46),
.C(n_36),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_L g165 ( 
.A(n_127),
.B(n_137),
.Y(n_165)
);

OAI22xp5_ASAP7_75t_SL g132 ( 
.A1(n_97),
.A2(n_70),
.B1(n_24),
.B2(n_33),
.Y(n_132)
);

OAI22xp5_ASAP7_75t_L g154 ( 
.A1(n_133),
.A2(n_112),
.B1(n_85),
.B2(n_91),
.Y(n_154)
);

INVxp67_ASAP7_75t_L g164 ( 
.A(n_134),
.Y(n_164)
);

AOI22xp33_ASAP7_75t_SL g135 ( 
.A1(n_90),
.A2(n_96),
.B1(n_103),
.B2(n_76),
.Y(n_135)
);

INVxp67_ASAP7_75t_L g166 ( 
.A(n_135),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_L g137 ( 
.A(n_82),
.B(n_26),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_L g142 ( 
.A(n_109),
.B(n_29),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_L g169 ( 
.A(n_142),
.B(n_79),
.Y(n_169)
);

AND2x2_ASAP7_75t_L g163 ( 
.A(n_143),
.B(n_145),
.Y(n_163)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_117),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_SL g208 ( 
.A(n_147),
.B(n_161),
.Y(n_208)
);

INVx2_ASAP7_75t_L g148 ( 
.A(n_125),
.Y(n_148)
);

INVx2_ASAP7_75t_L g202 ( 
.A(n_148),
.Y(n_202)
);

XOR2xp5_ASAP7_75t_L g149 ( 
.A(n_120),
.B(n_101),
.Y(n_149)
);

XNOR2xp5_ASAP7_75t_SL g204 ( 
.A(n_149),
.B(n_168),
.Y(n_204)
);

XNOR2xp5_ASAP7_75t_L g183 ( 
.A(n_150),
.B(n_160),
.Y(n_183)
);

BUFx6f_ASAP7_75t_L g151 ( 
.A(n_124),
.Y(n_151)
);

NOR2xp33_ASAP7_75t_L g184 ( 
.A(n_151),
.B(n_159),
.Y(n_184)
);

OAI22xp5_ASAP7_75t_SL g152 ( 
.A1(n_133),
.A2(n_140),
.B1(n_120),
.B2(n_119),
.Y(n_152)
);

AOI22xp5_ASAP7_75t_L g188 ( 
.A1(n_152),
.A2(n_154),
.B1(n_156),
.B2(n_157),
.Y(n_188)
);

AOI21xp5_ASAP7_75t_L g153 ( 
.A1(n_131),
.A2(n_77),
.B(n_115),
.Y(n_153)
);

AOI21xp5_ASAP7_75t_L g209 ( 
.A1(n_153),
.A2(n_171),
.B(n_6),
.Y(n_209)
);

OAI22xp5_ASAP7_75t_L g182 ( 
.A1(n_155),
.A2(n_167),
.B1(n_138),
.B2(n_139),
.Y(n_182)
);

OAI22xp5_ASAP7_75t_L g156 ( 
.A1(n_140),
.A2(n_112),
.B1(n_110),
.B2(n_104),
.Y(n_156)
);

OAI22xp5_ASAP7_75t_SL g157 ( 
.A1(n_126),
.A2(n_105),
.B1(n_92),
.B2(n_88),
.Y(n_157)
);

BUFx5_ASAP7_75t_L g159 ( 
.A(n_124),
.Y(n_159)
);

CKINVDCx20_ASAP7_75t_R g161 ( 
.A(n_146),
.Y(n_161)
);

AOI22xp5_ASAP7_75t_L g162 ( 
.A1(n_123),
.A2(n_83),
.B1(n_113),
.B2(n_98),
.Y(n_162)
);

OAI22xp5_ASAP7_75t_SL g197 ( 
.A1(n_162),
.A2(n_172),
.B1(n_144),
.B2(n_43),
.Y(n_197)
);

AOI22xp33_ASAP7_75t_SL g167 ( 
.A1(n_141),
.A2(n_29),
.B1(n_31),
.B2(n_33),
.Y(n_167)
);

XNOR2xp5_ASAP7_75t_L g168 ( 
.A(n_137),
.B(n_35),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_L g186 ( 
.A(n_169),
.B(n_178),
.Y(n_186)
);

INVx2_ASAP7_75t_L g170 ( 
.A(n_125),
.Y(n_170)
);

BUFx6f_ASAP7_75t_L g185 ( 
.A(n_170),
.Y(n_185)
);

AND2x2_ASAP7_75t_L g171 ( 
.A(n_142),
.B(n_46),
.Y(n_171)
);

AOI22xp5_ASAP7_75t_L g172 ( 
.A1(n_116),
.A2(n_132),
.B1(n_127),
.B2(n_128),
.Y(n_172)
);

OAI22xp5_ASAP7_75t_SL g173 ( 
.A1(n_117),
.A2(n_87),
.B1(n_43),
.B2(n_37),
.Y(n_173)
);

AOI22xp5_ASAP7_75t_L g191 ( 
.A1(n_173),
.A2(n_138),
.B1(n_129),
.B2(n_118),
.Y(n_191)
);

A2O1A1Ixp33_ASAP7_75t_L g174 ( 
.A1(n_130),
.A2(n_15),
.B(n_34),
.C(n_30),
.Y(n_174)
);

A2O1A1Ixp33_ASAP7_75t_L g180 ( 
.A1(n_174),
.A2(n_128),
.B(n_34),
.C(n_121),
.Y(n_180)
);

XOR2xp5_ASAP7_75t_L g175 ( 
.A(n_130),
.B(n_79),
.Y(n_175)
);

MAJIxp5_ASAP7_75t_L g190 ( 
.A(n_175),
.B(n_121),
.C(n_118),
.Y(n_190)
);

NOR2xp33_ASAP7_75t_SL g192 ( 
.A(n_176),
.B(n_0),
.Y(n_192)
);

INVx3_ASAP7_75t_L g177 ( 
.A(n_146),
.Y(n_177)
);

NOR2xp33_ASAP7_75t_L g207 ( 
.A(n_177),
.B(n_159),
.Y(n_207)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_136),
.Y(n_178)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_136),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_L g187 ( 
.A(n_179),
.B(n_139),
.Y(n_187)
);

OAI21xp5_ASAP7_75t_SL g216 ( 
.A1(n_180),
.A2(n_181),
.B(n_209),
.Y(n_216)
);

AND2x2_ASAP7_75t_L g181 ( 
.A(n_169),
.B(n_43),
.Y(n_181)
);

AOI22xp5_ASAP7_75t_L g213 ( 
.A1(n_182),
.A2(n_197),
.B1(n_198),
.B2(n_205),
.Y(n_213)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_187),
.Y(n_220)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_175),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_L g221 ( 
.A(n_189),
.B(n_196),
.Y(n_221)
);

XOR2xp5_ASAP7_75t_L g217 ( 
.A(n_190),
.B(n_168),
.Y(n_217)
);

OAI22xp5_ASAP7_75t_L g240 ( 
.A1(n_191),
.A2(n_210),
.B1(n_212),
.B2(n_10),
.Y(n_240)
);

NAND2xp5_ASAP7_75t_SL g230 ( 
.A(n_192),
.B(n_193),
.Y(n_230)
);

AND2x6_ASAP7_75t_L g193 ( 
.A(n_163),
.B(n_152),
.Y(n_193)
);

MAJIxp5_ASAP7_75t_L g194 ( 
.A(n_149),
.B(n_129),
.C(n_146),
.Y(n_194)
);

MAJIxp5_ASAP7_75t_L g214 ( 
.A(n_194),
.B(n_201),
.C(n_157),
.Y(n_214)
);

NAND3xp33_ASAP7_75t_L g195 ( 
.A(n_165),
.B(n_0),
.C(n_2),
.Y(n_195)
);

INVxp67_ASAP7_75t_L g225 ( 
.A(n_195),
.Y(n_225)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_173),
.Y(n_196)
);

OAI22xp5_ASAP7_75t_SL g198 ( 
.A1(n_155),
.A2(n_144),
.B1(n_34),
.B2(n_5),
.Y(n_198)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_162),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_L g234 ( 
.A(n_199),
.B(n_211),
.Y(n_234)
);

AOI22xp5_ASAP7_75t_L g200 ( 
.A1(n_163),
.A2(n_3),
.B1(n_4),
.B2(n_5),
.Y(n_200)
);

OAI22xp5_ASAP7_75t_SL g223 ( 
.A1(n_200),
.A2(n_203),
.B1(n_211),
.B2(n_209),
.Y(n_223)
);

MAJIxp5_ASAP7_75t_L g201 ( 
.A(n_160),
.B(n_3),
.C(n_4),
.Y(n_201)
);

AOI22xp5_ASAP7_75t_L g203 ( 
.A1(n_163),
.A2(n_3),
.B1(n_4),
.B2(n_5),
.Y(n_203)
);

OAI22xp5_ASAP7_75t_SL g205 ( 
.A1(n_172),
.A2(n_6),
.B1(n_7),
.B2(n_8),
.Y(n_205)
);

OAI22xp5_ASAP7_75t_SL g206 ( 
.A1(n_153),
.A2(n_6),
.B1(n_7),
.B2(n_8),
.Y(n_206)
);

AOI22xp5_ASAP7_75t_L g227 ( 
.A1(n_206),
.A2(n_170),
.B1(n_148),
.B2(n_11),
.Y(n_227)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_207),
.Y(n_229)
);

OAI22xp5_ASAP7_75t_L g210 ( 
.A1(n_166),
.A2(n_164),
.B1(n_147),
.B2(n_158),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_L g211 ( 
.A(n_165),
.B(n_7),
.Y(n_211)
);

OAI22xp5_ASAP7_75t_L g212 ( 
.A1(n_166),
.A2(n_7),
.B1(n_8),
.B2(n_9),
.Y(n_212)
);

XNOR2xp5_ASAP7_75t_L g247 ( 
.A(n_214),
.B(n_183),
.Y(n_247)
);

CKINVDCx20_ASAP7_75t_R g215 ( 
.A(n_185),
.Y(n_215)
);

CKINVDCx20_ASAP7_75t_R g252 ( 
.A(n_215),
.Y(n_252)
);

MAJIxp5_ASAP7_75t_L g246 ( 
.A(n_217),
.B(n_218),
.C(n_222),
.Y(n_246)
);

MAJIxp5_ASAP7_75t_L g218 ( 
.A(n_204),
.B(n_150),
.C(n_171),
.Y(n_218)
);

INVx3_ASAP7_75t_L g219 ( 
.A(n_185),
.Y(n_219)
);

NOR2xp33_ASAP7_75t_L g242 ( 
.A(n_219),
.B(n_223),
.Y(n_242)
);

MAJIxp5_ASAP7_75t_L g222 ( 
.A(n_204),
.B(n_171),
.C(n_178),
.Y(n_222)
);

OAI22xp5_ASAP7_75t_SL g224 ( 
.A1(n_196),
.A2(n_164),
.B1(n_179),
.B2(n_177),
.Y(n_224)
);

AOI22xp5_ASAP7_75t_L g261 ( 
.A1(n_224),
.A2(n_240),
.B1(n_223),
.B2(n_219),
.Y(n_261)
);

OAI21xp5_ASAP7_75t_SL g226 ( 
.A1(n_189),
.A2(n_174),
.B(n_151),
.Y(n_226)
);

OAI21xp5_ASAP7_75t_SL g249 ( 
.A1(n_226),
.A2(n_227),
.B(n_232),
.Y(n_249)
);

INVxp67_ASAP7_75t_L g228 ( 
.A(n_184),
.Y(n_228)
);

NAND2xp5_ASAP7_75t_L g244 ( 
.A(n_228),
.B(n_235),
.Y(n_244)
);

CKINVDCx20_ASAP7_75t_R g231 ( 
.A(n_187),
.Y(n_231)
);

CKINVDCx20_ASAP7_75t_R g254 ( 
.A(n_231),
.Y(n_254)
);

OAI21xp5_ASAP7_75t_SL g232 ( 
.A1(n_186),
.A2(n_9),
.B(n_10),
.Y(n_232)
);

CKINVDCx20_ASAP7_75t_R g233 ( 
.A(n_208),
.Y(n_233)
);

NOR2xp33_ASAP7_75t_L g256 ( 
.A(n_233),
.B(n_237),
.Y(n_256)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_186),
.Y(n_235)
);

INVxp67_ASAP7_75t_L g236 ( 
.A(n_191),
.Y(n_236)
);

NAND2xp5_ASAP7_75t_L g250 ( 
.A(n_236),
.B(n_238),
.Y(n_250)
);

INVx2_ASAP7_75t_L g237 ( 
.A(n_202),
.Y(n_237)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_181),
.Y(n_238)
);

OA22x2_ASAP7_75t_L g239 ( 
.A1(n_180),
.A2(n_198),
.B1(n_199),
.B2(n_197),
.Y(n_239)
);

AND2x2_ASAP7_75t_L g263 ( 
.A(n_239),
.B(n_202),
.Y(n_263)
);

OAI21xp5_ASAP7_75t_L g241 ( 
.A1(n_230),
.A2(n_193),
.B(n_190),
.Y(n_241)
);

MAJIxp5_ASAP7_75t_SL g272 ( 
.A(n_241),
.B(n_243),
.C(n_245),
.Y(n_272)
);

AOI21xp5_ASAP7_75t_L g243 ( 
.A1(n_226),
.A2(n_216),
.B(n_221),
.Y(n_243)
);

OAI21xp5_ASAP7_75t_L g245 ( 
.A1(n_216),
.A2(n_221),
.B(n_238),
.Y(n_245)
);

MAJIxp5_ASAP7_75t_L g279 ( 
.A(n_247),
.B(n_248),
.C(n_11),
.Y(n_279)
);

MAJIxp5_ASAP7_75t_L g248 ( 
.A(n_217),
.B(n_194),
.C(n_183),
.Y(n_248)
);

HB1xp67_ASAP7_75t_L g251 ( 
.A(n_234),
.Y(n_251)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_251),
.Y(n_267)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_234),
.Y(n_253)
);

NOR2xp33_ASAP7_75t_L g271 ( 
.A(n_253),
.B(n_262),
.Y(n_271)
);

OAI21xp5_ASAP7_75t_L g255 ( 
.A1(n_236),
.A2(n_181),
.B(n_201),
.Y(n_255)
);

NAND2xp5_ASAP7_75t_SL g265 ( 
.A(n_255),
.B(n_214),
.Y(n_265)
);

XNOR2xp5_ASAP7_75t_L g257 ( 
.A(n_222),
.B(n_188),
.Y(n_257)
);

XOR2xp5_ASAP7_75t_L g273 ( 
.A(n_257),
.B(n_259),
.Y(n_273)
);

NOR2xp33_ASAP7_75t_L g258 ( 
.A(n_229),
.B(n_205),
.Y(n_258)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_258),
.Y(n_275)
);

XNOR2xp5_ASAP7_75t_L g259 ( 
.A(n_218),
.B(n_188),
.Y(n_259)
);

OAI22xp5_ASAP7_75t_SL g260 ( 
.A1(n_213),
.A2(n_200),
.B1(n_203),
.B2(n_206),
.Y(n_260)
);

AOI22xp5_ASAP7_75t_L g281 ( 
.A1(n_260),
.A2(n_14),
.B1(n_12),
.B2(n_13),
.Y(n_281)
);

OAI22xp5_ASAP7_75t_L g266 ( 
.A1(n_261),
.A2(n_213),
.B1(n_227),
.B2(n_220),
.Y(n_266)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_224),
.Y(n_262)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_263),
.Y(n_264)
);

XNOR2xp5_ASAP7_75t_L g291 ( 
.A(n_265),
.B(n_274),
.Y(n_291)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_266),
.Y(n_288)
);

OAI22xp5_ASAP7_75t_L g268 ( 
.A1(n_261),
.A2(n_225),
.B1(n_229),
.B2(n_235),
.Y(n_268)
);

CKINVDCx14_ASAP7_75t_R g298 ( 
.A(n_268),
.Y(n_298)
);

OAI22xp5_ASAP7_75t_L g269 ( 
.A1(n_242),
.A2(n_225),
.B1(n_220),
.B2(n_228),
.Y(n_269)
);

CKINVDCx16_ASAP7_75t_R g285 ( 
.A(n_269),
.Y(n_285)
);

OAI22xp5_ASAP7_75t_L g270 ( 
.A1(n_262),
.A2(n_239),
.B1(n_232),
.B2(n_215),
.Y(n_270)
);

OAI22xp5_ASAP7_75t_L g292 ( 
.A1(n_270),
.A2(n_281),
.B1(n_255),
.B2(n_252),
.Y(n_292)
);

XNOR2xp5_ASAP7_75t_SL g274 ( 
.A(n_241),
.B(n_239),
.Y(n_274)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_256),
.Y(n_276)
);

NOR2xp33_ASAP7_75t_L g289 ( 
.A(n_276),
.B(n_282),
.Y(n_289)
);

XNOR2xp5_ASAP7_75t_L g277 ( 
.A(n_259),
.B(n_239),
.Y(n_277)
);

XNOR2xp5_ASAP7_75t_L g296 ( 
.A(n_277),
.B(n_278),
.Y(n_296)
);

XNOR2xp5_ASAP7_75t_L g278 ( 
.A(n_257),
.B(n_237),
.Y(n_278)
);

MAJIxp5_ASAP7_75t_L g293 ( 
.A(n_279),
.B(n_280),
.C(n_246),
.Y(n_293)
);

XOR2xp5_ASAP7_75t_L g280 ( 
.A(n_246),
.B(n_248),
.Y(n_280)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_244),
.Y(n_282)
);

OAI21xp33_ASAP7_75t_L g283 ( 
.A1(n_243),
.A2(n_12),
.B(n_13),
.Y(n_283)
);

NAND2xp5_ASAP7_75t_SL g287 ( 
.A(n_283),
.B(n_249),
.Y(n_287)
);

AOI22xp5_ASAP7_75t_SL g284 ( 
.A1(n_275),
.A2(n_263),
.B1(n_260),
.B2(n_254),
.Y(n_284)
);

OAI21xp5_ASAP7_75t_SL g311 ( 
.A1(n_284),
.A2(n_286),
.B(n_295),
.Y(n_311)
);

AOI22xp5_ASAP7_75t_SL g286 ( 
.A1(n_272),
.A2(n_263),
.B1(n_254),
.B2(n_253),
.Y(n_286)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_287),
.Y(n_306)
);

CKINVDCx20_ASAP7_75t_R g290 ( 
.A(n_271),
.Y(n_290)
);

CKINVDCx20_ASAP7_75t_R g310 ( 
.A(n_290),
.Y(n_310)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_292),
.Y(n_312)
);

XNOR2xp5_ASAP7_75t_L g303 ( 
.A(n_293),
.B(n_278),
.Y(n_303)
);

MAJIxp5_ASAP7_75t_L g294 ( 
.A(n_279),
.B(n_273),
.C(n_280),
.Y(n_294)
);

NAND2xp5_ASAP7_75t_SL g302 ( 
.A(n_294),
.B(n_297),
.Y(n_302)
);

AND2x2_ASAP7_75t_L g295 ( 
.A(n_277),
.B(n_244),
.Y(n_295)
);

MAJIxp5_ASAP7_75t_L g297 ( 
.A(n_273),
.B(n_247),
.C(n_245),
.Y(n_297)
);

BUFx24_ASAP7_75t_SL g299 ( 
.A(n_272),
.Y(n_299)
);

NAND2xp5_ASAP7_75t_SL g305 ( 
.A(n_299),
.B(n_281),
.Y(n_305)
);

NOR2xp67_ASAP7_75t_L g300 ( 
.A(n_286),
.B(n_274),
.Y(n_300)
);

OAI22xp5_ASAP7_75t_L g318 ( 
.A1(n_300),
.A2(n_301),
.B1(n_308),
.B2(n_309),
.Y(n_318)
);

OAI22x1_ASAP7_75t_L g301 ( 
.A1(n_284),
.A2(n_249),
.B1(n_264),
.B2(n_283),
.Y(n_301)
);

XNOR2xp5_ASAP7_75t_L g317 ( 
.A(n_303),
.B(n_304),
.Y(n_317)
);

XNOR2xp5_ASAP7_75t_L g304 ( 
.A(n_296),
.B(n_250),
.Y(n_304)
);

NAND2xp5_ASAP7_75t_L g319 ( 
.A(n_305),
.B(n_307),
.Y(n_319)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_289),
.Y(n_307)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_295),
.Y(n_308)
);

OAI22xp5_ASAP7_75t_SL g309 ( 
.A1(n_285),
.A2(n_264),
.B1(n_282),
.B2(n_250),
.Y(n_309)
);

MAJIxp5_ASAP7_75t_L g313 ( 
.A(n_303),
.B(n_294),
.C(n_293),
.Y(n_313)
);

MAJIxp5_ASAP7_75t_L g324 ( 
.A(n_313),
.B(n_314),
.C(n_316),
.Y(n_324)
);

MAJIxp5_ASAP7_75t_L g314 ( 
.A(n_302),
.B(n_312),
.C(n_297),
.Y(n_314)
);

XOR2xp5_ASAP7_75t_L g315 ( 
.A(n_311),
.B(n_291),
.Y(n_315)
);

XOR2xp5_ASAP7_75t_L g327 ( 
.A(n_315),
.B(n_318),
.Y(n_327)
);

MAJIxp5_ASAP7_75t_L g316 ( 
.A(n_312),
.B(n_298),
.C(n_288),
.Y(n_316)
);

AOI21xp5_ASAP7_75t_L g320 ( 
.A1(n_311),
.A2(n_252),
.B(n_267),
.Y(n_320)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_320),
.Y(n_325)
);

INVx2_ASAP7_75t_L g321 ( 
.A(n_301),
.Y(n_321)
);

NOR2xp33_ASAP7_75t_L g323 ( 
.A(n_321),
.B(n_309),
.Y(n_323)
);

OAI21xp5_ASAP7_75t_SL g322 ( 
.A1(n_320),
.A2(n_310),
.B(n_306),
.Y(n_322)
);

NAND2xp5_ASAP7_75t_L g330 ( 
.A(n_322),
.B(n_326),
.Y(n_330)
);

INVxp33_ASAP7_75t_L g332 ( 
.A(n_323),
.Y(n_332)
);

NAND2xp5_ASAP7_75t_SL g326 ( 
.A(n_314),
.B(n_304),
.Y(n_326)
);

XOR2xp5_ASAP7_75t_L g329 ( 
.A(n_327),
.B(n_315),
.Y(n_329)
);

NOR2xp33_ASAP7_75t_L g328 ( 
.A(n_316),
.B(n_13),
.Y(n_328)
);

MAJIxp5_ASAP7_75t_L g331 ( 
.A(n_328),
.B(n_319),
.C(n_317),
.Y(n_331)
);

NOR2xp33_ASAP7_75t_L g333 ( 
.A(n_329),
.B(n_331),
.Y(n_333)
);

OAI21xp5_ASAP7_75t_L g334 ( 
.A1(n_330),
.A2(n_324),
.B(n_325),
.Y(n_334)
);

NAND2xp5_ASAP7_75t_L g335 ( 
.A(n_334),
.B(n_324),
.Y(n_335)
);

XOR2xp5_ASAP7_75t_L g336 ( 
.A(n_335),
.B(n_333),
.Y(n_336)
);

A2O1A1Ixp33_ASAP7_75t_L g337 ( 
.A1(n_336),
.A2(n_313),
.B(n_332),
.C(n_327),
.Y(n_337)
);

AOI21xp5_ASAP7_75t_L g338 ( 
.A1(n_337),
.A2(n_317),
.B(n_332),
.Y(n_338)
);

BUFx24_ASAP7_75t_SL g339 ( 
.A(n_338),
.Y(n_339)
);

NAND2xp5_ASAP7_75t_L g340 ( 
.A(n_339),
.B(n_14),
.Y(n_340)
);


endmodule