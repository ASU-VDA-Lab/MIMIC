module real_jpeg_25292_n_16 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_3, n_10, n_356, n_9, n_16);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_3;
input n_10;
input n_356;
input n_9;

output n_16;

wire n_37;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_300;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_199;
wire n_95;
wire n_238;
wire n_67;
wire n_350;
wire n_235;
wire n_107;
wire n_354;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_123;
wire n_50;
wire n_186;
wire n_137;
wire n_72;
wire n_171;
wire n_151;
wire n_272;
wire n_203;
wire n_198;
wire n_23;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_326;
wire n_339;
wire n_80;
wire n_30;
wire n_332;
wire n_149;
wire n_328;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_353;
wire n_230;
wire n_216;
wire n_128;
wire n_202;
wire n_127;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_348;
wire n_252;
wire n_310;
wire n_345;
wire n_78;
wire n_83;
wire n_288;
wire n_221;
wire n_104;
wire n_153;
wire n_337;
wire n_131;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_200;
wire n_335;
wire n_214;
wire n_113;
wire n_251;
wire n_139;
wire n_33;
wire n_175;
wire n_338;
wire n_156;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_77;
wire n_219;
wire n_122;
wire n_19;
wire n_262;
wire n_334;
wire n_17;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_195;
wire n_110;
wire n_289;
wire n_117;
wire n_193;
wire n_20;
wire n_278;
wire n_314;
wire n_103;
wire n_232;
wire n_212;
wire n_284;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_213;
wire n_25;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_341;
wire n_331;
wire n_49;
wire n_68;
wire n_146;
wire n_323;
wire n_286;
wire n_176;
wire n_166;
wire n_215;
wire n_312;
wire n_325;
wire n_316;
wire n_307;
wire n_161;
wire n_207;
wire n_237;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_140;
wire n_126;
wire n_342;
wire n_120;
wire n_155;
wire n_319;
wire n_93;
wire n_242;
wire n_142;
wire n_76;
wire n_79;
wire n_282;
wire n_147;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_18;
wire n_145;
wire n_266;
wire n_109;
wire n_148;
wire n_196;
wire n_298;
wire n_330;
wire n_333;
wire n_152;
wire n_270;
wire n_159;
wire n_347;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_336;
wire n_258;
wire n_150;
wire n_41;
wire n_74;
wire n_158;
wire n_204;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_75;
wire n_346;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_119;
wire n_283;
wire n_181;
wire n_256;
wire n_253;
wire n_273;
wire n_54;
wire n_168;
wire n_38;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_349;
wire n_292;
wire n_343;
wire n_64;
wire n_291;
wire n_236;
wire n_276;
wire n_287;
wire n_174;
wire n_255;
wire n_243;
wire n_299;
wire n_352;
wire n_56;
wire n_293;
wire n_275;
wire n_227;
wire n_229;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_45;
wire n_268;
wire n_42;
wire n_313;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_143;
wire n_351;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_303;
wire n_321;
wire n_100;
wire n_51;
wire n_205;
wire n_261;
wire n_86;
wire n_324;
wire n_70;
wire n_32;
wire n_228;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_133;
wire n_257;
wire n_344;
wire n_210;
wire n_206;
wire n_85;
wire n_96;
wire n_308;

AOI22xp33_ASAP7_75t_SL g44 ( 
.A1(n_0),
.A2(n_45),
.B1(n_46),
.B2(n_48),
.Y(n_44)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_0),
.Y(n_48)
);

AOI22xp5_ASAP7_75t_SL g108 ( 
.A1(n_0),
.A2(n_30),
.B1(n_31),
.B2(n_48),
.Y(n_108)
);

AOI22xp33_ASAP7_75t_SL g262 ( 
.A1(n_0),
.A2(n_48),
.B1(n_62),
.B2(n_65),
.Y(n_262)
);

AOI22xp33_ASAP7_75t_SL g302 ( 
.A1(n_0),
.A2(n_48),
.B1(n_77),
.B2(n_86),
.Y(n_302)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_1),
.Y(n_63)
);

OAI22xp33_ASAP7_75t_SL g61 ( 
.A1(n_2),
.A2(n_62),
.B1(n_64),
.B2(n_65),
.Y(n_61)
);

CKINVDCx16_ASAP7_75t_R g64 ( 
.A(n_2),
.Y(n_64)
);

OAI22xp33_ASAP7_75t_SL g98 ( 
.A1(n_2),
.A2(n_64),
.B1(n_76),
.B2(n_77),
.Y(n_98)
);

AOI22xp5_ASAP7_75t_SL g158 ( 
.A1(n_2),
.A2(n_45),
.B1(n_46),
.B2(n_64),
.Y(n_158)
);

AOI22xp33_ASAP7_75t_L g163 ( 
.A1(n_2),
.A2(n_30),
.B1(n_31),
.B2(n_64),
.Y(n_163)
);

INVx1_ASAP7_75t_SL g42 ( 
.A(n_3),
.Y(n_42)
);

BUFx12f_ASAP7_75t_L g31 ( 
.A(n_4),
.Y(n_31)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_5),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_5),
.B(n_88),
.Y(n_127)
);

MAJIxp5_ASAP7_75t_L g140 ( 
.A(n_5),
.B(n_31),
.C(n_43),
.Y(n_140)
);

OAI22xp5_ASAP7_75t_L g142 ( 
.A1(n_5),
.A2(n_45),
.B1(n_46),
.B2(n_78),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_L g155 ( 
.A(n_5),
.B(n_71),
.Y(n_155)
);

OAI22xp5_ASAP7_75t_L g173 ( 
.A1(n_5),
.A2(n_28),
.B1(n_170),
.B2(n_174),
.Y(n_173)
);

INVx8_ASAP7_75t_SL g82 ( 
.A(n_6),
.Y(n_82)
);

OAI22xp5_ASAP7_75t_L g35 ( 
.A1(n_7),
.A2(n_30),
.B1(n_31),
.B2(n_36),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_7),
.Y(n_36)
);

OAI22xp5_ASAP7_75t_L g229 ( 
.A1(n_7),
.A2(n_36),
.B1(n_45),
.B2(n_46),
.Y(n_229)
);

OAI22xp5_ASAP7_75t_L g277 ( 
.A1(n_7),
.A2(n_36),
.B1(n_62),
.B2(n_65),
.Y(n_277)
);

OAI22xp5_ASAP7_75t_L g322 ( 
.A1(n_7),
.A2(n_36),
.B1(n_259),
.B2(n_323),
.Y(n_322)
);

OAI22xp5_ASAP7_75t_SL g57 ( 
.A1(n_8),
.A2(n_45),
.B1(n_46),
.B2(n_58),
.Y(n_57)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_8),
.Y(n_58)
);

OAI22xp5_ASAP7_75t_L g103 ( 
.A1(n_8),
.A2(n_58),
.B1(n_62),
.B2(n_65),
.Y(n_103)
);

AOI22xp5_ASAP7_75t_L g152 ( 
.A1(n_8),
.A2(n_30),
.B1(n_31),
.B2(n_58),
.Y(n_152)
);

OAI22xp5_ASAP7_75t_SL g258 ( 
.A1(n_8),
.A2(n_58),
.B1(n_86),
.B2(n_259),
.Y(n_258)
);

BUFx12f_ASAP7_75t_L g68 ( 
.A(n_9),
.Y(n_68)
);

OAI22xp5_ASAP7_75t_L g38 ( 
.A1(n_10),
.A2(n_30),
.B1(n_31),
.B2(n_39),
.Y(n_38)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_10),
.Y(n_39)
);

AOI22xp33_ASAP7_75t_L g54 ( 
.A1(n_10),
.A2(n_39),
.B1(n_45),
.B2(n_46),
.Y(n_54)
);

AOI22xp33_ASAP7_75t_L g238 ( 
.A1(n_10),
.A2(n_39),
.B1(n_62),
.B2(n_65),
.Y(n_238)
);

OAI22xp5_ASAP7_75t_SL g288 ( 
.A1(n_10),
.A2(n_39),
.B1(n_76),
.B2(n_289),
.Y(n_288)
);

OAI22xp5_ASAP7_75t_L g72 ( 
.A1(n_11),
.A2(n_62),
.B1(n_65),
.B2(n_73),
.Y(n_72)
);

CKINVDCx20_ASAP7_75t_R g73 ( 
.A(n_11),
.Y(n_73)
);

AOI22xp5_ASAP7_75t_SL g148 ( 
.A1(n_11),
.A2(n_30),
.B1(n_31),
.B2(n_73),
.Y(n_148)
);

OAI22xp5_ASAP7_75t_L g195 ( 
.A1(n_11),
.A2(n_45),
.B1(n_46),
.B2(n_73),
.Y(n_195)
);

OAI22xp5_ASAP7_75t_L g235 ( 
.A1(n_11),
.A2(n_73),
.B1(n_85),
.B2(n_86),
.Y(n_235)
);

INVx13_ASAP7_75t_L g77 ( 
.A(n_12),
.Y(n_77)
);

NAND3xp33_ASAP7_75t_L g114 ( 
.A(n_12),
.B(n_65),
.C(n_83),
.Y(n_114)
);

AOI22xp33_ASAP7_75t_L g90 ( 
.A1(n_13),
.A2(n_85),
.B1(n_86),
.B2(n_91),
.Y(n_90)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_13),
.Y(n_91)
);

OAI22xp5_ASAP7_75t_L g130 ( 
.A1(n_13),
.A2(n_62),
.B1(n_65),
.B2(n_91),
.Y(n_130)
);

AOI22xp5_ASAP7_75t_L g145 ( 
.A1(n_13),
.A2(n_45),
.B1(n_46),
.B2(n_91),
.Y(n_145)
);

AOI22xp5_ASAP7_75t_L g170 ( 
.A1(n_13),
.A2(n_30),
.B1(n_31),
.B2(n_91),
.Y(n_170)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_14),
.Y(n_47)
);

INVx6_ASAP7_75t_L g33 ( 
.A(n_15),
.Y(n_33)
);

INVx6_ASAP7_75t_L g112 ( 
.A(n_15),
.Y(n_112)
);

INVx3_ASAP7_75t_L g174 ( 
.A(n_15),
.Y(n_174)
);

INVx2_ASAP7_75t_L g177 ( 
.A(n_15),
.Y(n_177)
);

MAJx2_ASAP7_75t_L g16 ( 
.A(n_17),
.B(n_349),
.C(n_354),
.Y(n_16)
);

OAI21xp5_ASAP7_75t_SL g17 ( 
.A1(n_18),
.A2(n_347),
.B(n_352),
.Y(n_17)
);

AOI21xp5_ASAP7_75t_L g18 ( 
.A1(n_19),
.A2(n_334),
.B(n_346),
.Y(n_18)
);

OAI321xp33_ASAP7_75t_L g19 ( 
.A1(n_20),
.A2(n_297),
.A3(n_327),
.B1(n_332),
.B2(n_333),
.C(n_356),
.Y(n_19)
);

AOI21xp5_ASAP7_75t_L g20 ( 
.A1(n_21),
.A2(n_270),
.B(n_296),
.Y(n_20)
);

OAI21xp5_ASAP7_75t_SL g21 ( 
.A1(n_22),
.A2(n_241),
.B(n_269),
.Y(n_21)
);

O2A1O1Ixp33_ASAP7_75t_SL g22 ( 
.A1(n_23),
.A2(n_132),
.B(n_220),
.C(n_240),
.Y(n_22)
);

AND2x2_ASAP7_75t_L g23 ( 
.A(n_24),
.B(n_116),
.Y(n_23)
);

NOR2xp33_ASAP7_75t_L g219 ( 
.A(n_24),
.B(n_116),
.Y(n_219)
);

XNOR2xp5_ASAP7_75t_L g24 ( 
.A(n_25),
.B(n_92),
.Y(n_24)
);

XNOR2xp5_ASAP7_75t_L g25 ( 
.A(n_26),
.B(n_55),
.Y(n_25)
);

MAJIxp5_ASAP7_75t_L g221 ( 
.A(n_26),
.B(n_55),
.C(n_92),
.Y(n_221)
);

XOR2xp5_ASAP7_75t_L g26 ( 
.A(n_27),
.B(n_40),
.Y(n_26)
);

NAND2xp5_ASAP7_75t_L g232 ( 
.A(n_27),
.B(n_40),
.Y(n_232)
);

OAI21xp5_ASAP7_75t_L g27 ( 
.A1(n_28),
.A2(n_34),
.B(n_37),
.Y(n_27)
);

OAI21xp5_ASAP7_75t_L g147 ( 
.A1(n_28),
.A2(n_148),
.B(n_149),
.Y(n_147)
);

OAI22xp5_ASAP7_75t_L g169 ( 
.A1(n_28),
.A2(n_163),
.B1(n_170),
.B2(n_171),
.Y(n_169)
);

OAI21xp5_ASAP7_75t_L g190 ( 
.A1(n_28),
.A2(n_37),
.B(n_152),
.Y(n_190)
);

AOI21xp5_ASAP7_75t_L g247 ( 
.A1(n_28),
.A2(n_152),
.B(n_174),
.Y(n_247)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_29),
.Y(n_28)
);

AOI22xp5_ASAP7_75t_L g106 ( 
.A1(n_29),
.A2(n_35),
.B1(n_107),
.B2(n_109),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_SL g125 ( 
.A(n_29),
.B(n_38),
.Y(n_125)
);

AOI22xp5_ASAP7_75t_L g161 ( 
.A1(n_29),
.A2(n_124),
.B1(n_162),
.B2(n_164),
.Y(n_161)
);

NOR2xp33_ASAP7_75t_L g29 ( 
.A(n_30),
.B(n_32),
.Y(n_29)
);

OA22x2_ASAP7_75t_L g41 ( 
.A1(n_30),
.A2(n_31),
.B1(n_42),
.B2(n_43),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g175 ( 
.A(n_30),
.B(n_176),
.Y(n_175)
);

INVx6_ASAP7_75t_L g30 ( 
.A(n_31),
.Y(n_30)
);

NAND2xp5_ASAP7_75t_SL g37 ( 
.A(n_32),
.B(n_38),
.Y(n_37)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_32),
.Y(n_171)
);

INVx2_ASAP7_75t_L g32 ( 
.A(n_33),
.Y(n_32)
);

INVx5_ASAP7_75t_L g124 ( 
.A(n_33),
.Y(n_124)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_35),
.Y(n_34)
);

OAI21xp5_ASAP7_75t_L g40 ( 
.A1(n_41),
.A2(n_44),
.B(n_49),
.Y(n_40)
);

NAND2xp5_ASAP7_75t_L g51 ( 
.A(n_41),
.B(n_52),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_41),
.B(n_54),
.Y(n_59)
);

CKINVDCx20_ASAP7_75t_R g143 ( 
.A(n_41),
.Y(n_143)
);

OAI22xp5_ASAP7_75t_SL g157 ( 
.A1(n_41),
.A2(n_51),
.B1(n_145),
.B2(n_158),
.Y(n_157)
);

NOR2xp33_ASAP7_75t_L g168 ( 
.A(n_41),
.B(n_78),
.Y(n_168)
);

AOI21xp5_ASAP7_75t_L g307 ( 
.A1(n_41),
.A2(n_51),
.B(n_308),
.Y(n_307)
);

INVx3_ASAP7_75t_SL g43 ( 
.A(n_42),
.Y(n_43)
);

OAI22xp33_ASAP7_75t_L g52 ( 
.A1(n_42),
.A2(n_43),
.B1(n_45),
.B2(n_46),
.Y(n_52)
);

CKINVDCx16_ASAP7_75t_R g228 ( 
.A(n_44),
.Y(n_228)
);

AOI22xp5_ASAP7_75t_L g70 ( 
.A1(n_45),
.A2(n_46),
.B1(n_68),
.B2(n_69),
.Y(n_70)
);

O2A1O1Ixp33_ASAP7_75t_L g185 ( 
.A1(n_45),
.A2(n_69),
.B(n_186),
.C(n_188),
.Y(n_185)
);

INVx3_ASAP7_75t_L g45 ( 
.A(n_46),
.Y(n_45)
);

NAND2xp5_ASAP7_75t_L g139 ( 
.A(n_46),
.B(n_140),
.Y(n_139)
);

NOR3xp33_ASAP7_75t_L g188 ( 
.A(n_46),
.B(n_65),
.C(n_68),
.Y(n_188)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_47),
.Y(n_46)
);

AND2x2_ASAP7_75t_L g278 ( 
.A(n_49),
.B(n_210),
.Y(n_278)
);

NAND2xp5_ASAP7_75t_SL g49 ( 
.A(n_50),
.B(n_53),
.Y(n_49)
);

AOI21xp5_ASAP7_75t_L g56 ( 
.A1(n_50),
.A2(n_57),
.B(n_59),
.Y(n_56)
);

AOI22xp5_ASAP7_75t_L g141 ( 
.A1(n_50),
.A2(n_142),
.B1(n_143),
.B2(n_144),
.Y(n_141)
);

AOI22xp5_ASAP7_75t_L g193 ( 
.A1(n_50),
.A2(n_143),
.B1(n_194),
.B2(n_195),
.Y(n_193)
);

AOI22xp5_ASAP7_75t_L g227 ( 
.A1(n_50),
.A2(n_143),
.B1(n_228),
.B2(n_229),
.Y(n_227)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_51),
.Y(n_50)
);

OAI21xp5_ASAP7_75t_SL g208 ( 
.A1(n_51),
.A2(n_209),
.B(n_210),
.Y(n_208)
);

OAI21xp5_ASAP7_75t_SL g248 ( 
.A1(n_51),
.A2(n_249),
.B(n_250),
.Y(n_248)
);

INVxp67_ASAP7_75t_L g53 ( 
.A(n_54),
.Y(n_53)
);

MAJIxp5_ASAP7_75t_L g55 ( 
.A(n_56),
.B(n_60),
.C(n_74),
.Y(n_55)
);

XOR2xp5_ASAP7_75t_L g118 ( 
.A(n_56),
.B(n_60),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_SL g210 ( 
.A(n_57),
.B(n_143),
.Y(n_210)
);

CKINVDCx16_ASAP7_75t_R g308 ( 
.A(n_57),
.Y(n_308)
);

INVxp67_ASAP7_75t_L g250 ( 
.A(n_59),
.Y(n_250)
);

AOI22xp5_ASAP7_75t_L g60 ( 
.A1(n_61),
.A2(n_66),
.B1(n_71),
.B2(n_72),
.Y(n_60)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_61),
.Y(n_131)
);

INVx5_ASAP7_75t_L g65 ( 
.A(n_62),
.Y(n_65)
);

OAI22xp5_ASAP7_75t_L g67 ( 
.A1(n_62),
.A2(n_65),
.B1(n_68),
.B2(n_69),
.Y(n_67)
);

AOI22xp5_ASAP7_75t_L g80 ( 
.A1(n_62),
.A2(n_65),
.B1(n_81),
.B2(n_83),
.Y(n_80)
);

A2O1A1Ixp33_ASAP7_75t_L g113 ( 
.A1(n_62),
.A2(n_75),
.B(n_81),
.C(n_114),
.Y(n_113)
);

HAxp5_ASAP7_75t_SL g187 ( 
.A(n_62),
.B(n_78),
.CON(n_187),
.SN(n_187)
);

BUFx12f_ASAP7_75t_L g62 ( 
.A(n_63),
.Y(n_62)
);

CKINVDCx20_ASAP7_75t_R g101 ( 
.A(n_66),
.Y(n_101)
);

AOI22xp5_ASAP7_75t_L g192 ( 
.A1(n_66),
.A2(n_71),
.B1(n_130),
.B2(n_187),
.Y(n_192)
);

AOI21xp5_ASAP7_75t_L g236 ( 
.A1(n_66),
.A2(n_103),
.B(n_237),
.Y(n_236)
);

NAND2xp5_ASAP7_75t_SL g263 ( 
.A(n_66),
.B(n_264),
.Y(n_263)
);

AOI22xp5_ASAP7_75t_L g275 ( 
.A1(n_66),
.A2(n_71),
.B1(n_276),
.B2(n_277),
.Y(n_275)
);

AOI21xp5_ASAP7_75t_L g310 ( 
.A1(n_66),
.A2(n_237),
.B(n_277),
.Y(n_310)
);

OAI21xp5_ASAP7_75t_SL g339 ( 
.A1(n_66),
.A2(n_71),
.B(n_103),
.Y(n_339)
);

AND2x2_ASAP7_75t_L g66 ( 
.A(n_67),
.B(n_70),
.Y(n_66)
);

INVx5_ASAP7_75t_L g69 ( 
.A(n_68),
.Y(n_69)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_70),
.Y(n_71)
);

OAI22xp5_ASAP7_75t_L g128 ( 
.A1(n_70),
.A2(n_101),
.B1(n_129),
.B2(n_131),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_L g237 ( 
.A(n_70),
.B(n_238),
.Y(n_237)
);

OAI21xp5_ASAP7_75t_L g261 ( 
.A1(n_70),
.A2(n_262),
.B(n_263),
.Y(n_261)
);

NAND2xp5_ASAP7_75t_SL g102 ( 
.A(n_71),
.B(n_103),
.Y(n_102)
);

CKINVDCx20_ASAP7_75t_R g100 ( 
.A(n_72),
.Y(n_100)
);

XOR2xp5_ASAP7_75t_L g117 ( 
.A(n_74),
.B(n_118),
.Y(n_117)
);

AOI22xp5_ASAP7_75t_L g74 ( 
.A1(n_75),
.A2(n_79),
.B1(n_88),
.B2(n_89),
.Y(n_74)
);

HAxp5_ASAP7_75t_SL g75 ( 
.A(n_76),
.B(n_78),
.CON(n_75),
.SN(n_75)
);

INVx11_ASAP7_75t_L g259 ( 
.A(n_76),
.Y(n_259)
);

INVx8_ASAP7_75t_L g76 ( 
.A(n_77),
.Y(n_76)
);

INVx11_ASAP7_75t_L g86 ( 
.A(n_77),
.Y(n_86)
);

INVx8_ASAP7_75t_L g87 ( 
.A(n_77),
.Y(n_87)
);

INVx6_ASAP7_75t_L g325 ( 
.A(n_77),
.Y(n_325)
);

NOR2xp33_ASAP7_75t_L g176 ( 
.A(n_78),
.B(n_177),
.Y(n_176)
);

CKINVDCx20_ASAP7_75t_R g96 ( 
.A(n_79),
.Y(n_96)
);

AOI22xp5_ASAP7_75t_L g234 ( 
.A1(n_79),
.A2(n_88),
.B1(n_98),
.B2(n_235),
.Y(n_234)
);

NAND2xp5_ASAP7_75t_L g303 ( 
.A(n_79),
.B(n_288),
.Y(n_303)
);

AOI22xp5_ASAP7_75t_L g320 ( 
.A1(n_79),
.A2(n_88),
.B1(n_321),
.B2(n_322),
.Y(n_320)
);

AOI21xp5_ASAP7_75t_L g340 ( 
.A1(n_79),
.A2(n_322),
.B(n_341),
.Y(n_340)
);

OAI21xp5_ASAP7_75t_SL g354 ( 
.A1(n_79),
.A2(n_88),
.B(n_258),
.Y(n_354)
);

AND2x2_ASAP7_75t_SL g79 ( 
.A(n_80),
.B(n_84),
.Y(n_79)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_80),
.Y(n_88)
);

OAI22xp5_ASAP7_75t_SL g95 ( 
.A1(n_80),
.A2(n_90),
.B1(n_96),
.B2(n_97),
.Y(n_95)
);

OAI21xp5_ASAP7_75t_L g301 ( 
.A1(n_80),
.A2(n_302),
.B(n_303),
.Y(n_301)
);

CKINVDCx5p33_ASAP7_75t_R g83 ( 
.A(n_81),
.Y(n_83)
);

OAI22xp33_ASAP7_75t_L g84 ( 
.A1(n_81),
.A2(n_83),
.B1(n_85),
.B2(n_87),
.Y(n_84)
);

INVx8_ASAP7_75t_L g81 ( 
.A(n_82),
.Y(n_81)
);

INVx8_ASAP7_75t_L g85 ( 
.A(n_86),
.Y(n_85)
);

INVx4_ASAP7_75t_L g289 ( 
.A(n_87),
.Y(n_289)
);

NAND2xp5_ASAP7_75t_SL g257 ( 
.A(n_88),
.B(n_258),
.Y(n_257)
);

NAND2xp5_ASAP7_75t_SL g287 ( 
.A(n_88),
.B(n_288),
.Y(n_287)
);

CKINVDCx14_ASAP7_75t_R g89 ( 
.A(n_90),
.Y(n_89)
);

OAI22xp5_ASAP7_75t_SL g92 ( 
.A1(n_93),
.A2(n_94),
.B1(n_104),
.B2(n_115),
.Y(n_92)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_94),
.Y(n_93)
);

XNOR2xp5_ASAP7_75t_SL g94 ( 
.A(n_95),
.B(n_99),
.Y(n_94)
);

MAJIxp5_ASAP7_75t_L g239 ( 
.A(n_95),
.B(n_99),
.C(n_115),
.Y(n_239)
);

OAI21xp5_ASAP7_75t_L g255 ( 
.A1(n_96),
.A2(n_256),
.B(n_257),
.Y(n_255)
);

OAI21xp5_ASAP7_75t_SL g285 ( 
.A1(n_96),
.A2(n_286),
.B(n_287),
.Y(n_285)
);

CKINVDCx14_ASAP7_75t_R g97 ( 
.A(n_98),
.Y(n_97)
);

OAI21xp5_ASAP7_75t_L g99 ( 
.A1(n_100),
.A2(n_101),
.B(n_102),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g319 ( 
.A(n_102),
.B(n_263),
.Y(n_319)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_104),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_L g104 ( 
.A(n_105),
.B(n_113),
.Y(n_104)
);

AOI22xp5_ASAP7_75t_L g119 ( 
.A1(n_105),
.A2(n_106),
.B1(n_113),
.B2(n_120),
.Y(n_119)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_106),
.Y(n_105)
);

CKINVDCx20_ASAP7_75t_R g107 ( 
.A(n_108),
.Y(n_107)
);

OAI21xp5_ASAP7_75t_L g122 ( 
.A1(n_108),
.A2(n_123),
.B(n_125),
.Y(n_122)
);

INVx3_ASAP7_75t_L g109 ( 
.A(n_110),
.Y(n_109)
);

INVx5_ASAP7_75t_L g110 ( 
.A(n_111),
.Y(n_110)
);

INVx8_ASAP7_75t_L g111 ( 
.A(n_112),
.Y(n_111)
);

INVx3_ASAP7_75t_SL g150 ( 
.A(n_112),
.Y(n_150)
);

CKINVDCx20_ASAP7_75t_R g120 ( 
.A(n_113),
.Y(n_120)
);

MAJIxp5_ASAP7_75t_L g116 ( 
.A(n_117),
.B(n_119),
.C(n_121),
.Y(n_116)
);

XNOR2xp5_ASAP7_75t_L g215 ( 
.A(n_117),
.B(n_216),
.Y(n_215)
);

XNOR2xp5_ASAP7_75t_L g216 ( 
.A(n_119),
.B(n_121),
.Y(n_216)
);

MAJIxp5_ASAP7_75t_L g121 ( 
.A(n_122),
.B(n_126),
.C(n_128),
.Y(n_121)
);

AOI22xp5_ASAP7_75t_L g203 ( 
.A1(n_122),
.A2(n_126),
.B1(n_127),
.B2(n_204),
.Y(n_203)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_122),
.Y(n_204)
);

INVx5_ASAP7_75t_L g123 ( 
.A(n_124),
.Y(n_123)
);

AND2x2_ASAP7_75t_L g226 ( 
.A(n_125),
.B(n_149),
.Y(n_226)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_127),
.Y(n_126)
);

XOR2xp5_ASAP7_75t_L g202 ( 
.A(n_128),
.B(n_203),
.Y(n_202)
);

CKINVDCx16_ASAP7_75t_R g129 ( 
.A(n_130),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_SL g132 ( 
.A(n_133),
.B(n_219),
.Y(n_132)
);

AOI21xp5_ASAP7_75t_L g133 ( 
.A1(n_134),
.A2(n_214),
.B(n_218),
.Y(n_133)
);

OAI21xp5_ASAP7_75t_SL g134 ( 
.A1(n_135),
.A2(n_198),
.B(n_213),
.Y(n_134)
);

AOI21xp5_ASAP7_75t_SL g135 ( 
.A1(n_136),
.A2(n_181),
.B(n_197),
.Y(n_135)
);

OAI21xp5_ASAP7_75t_SL g136 ( 
.A1(n_137),
.A2(n_159),
.B(n_180),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_L g137 ( 
.A(n_138),
.B(n_146),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_L g180 ( 
.A(n_138),
.B(n_146),
.Y(n_180)
);

NOR2xp33_ASAP7_75t_L g138 ( 
.A(n_139),
.B(n_141),
.Y(n_138)
);

XNOR2xp5_ASAP7_75t_L g165 ( 
.A(n_139),
.B(n_141),
.Y(n_165)
);

CKINVDCx14_ASAP7_75t_R g144 ( 
.A(n_145),
.Y(n_144)
);

XNOR2xp5_ASAP7_75t_L g146 ( 
.A(n_147),
.B(n_153),
.Y(n_146)
);

MAJIxp5_ASAP7_75t_L g196 ( 
.A(n_147),
.B(n_154),
.C(n_157),
.Y(n_196)
);

CKINVDCx14_ASAP7_75t_R g164 ( 
.A(n_148),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_L g149 ( 
.A(n_150),
.B(n_151),
.Y(n_149)
);

CKINVDCx16_ASAP7_75t_R g151 ( 
.A(n_152),
.Y(n_151)
);

AOI22xp5_ASAP7_75t_L g153 ( 
.A1(n_154),
.A2(n_155),
.B1(n_156),
.B2(n_157),
.Y(n_153)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_155),
.Y(n_154)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_157),
.Y(n_156)
);

CKINVDCx14_ASAP7_75t_R g194 ( 
.A(n_158),
.Y(n_194)
);

AOI21xp5_ASAP7_75t_L g159 ( 
.A1(n_160),
.A2(n_166),
.B(n_179),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_L g160 ( 
.A(n_161),
.B(n_165),
.Y(n_160)
);

NOR2xp33_ASAP7_75t_L g179 ( 
.A(n_161),
.B(n_165),
.Y(n_179)
);

CKINVDCx14_ASAP7_75t_R g162 ( 
.A(n_163),
.Y(n_162)
);

OAI21xp5_ASAP7_75t_SL g166 ( 
.A1(n_167),
.A2(n_172),
.B(n_178),
.Y(n_166)
);

NOR2xp33_ASAP7_75t_L g167 ( 
.A(n_168),
.B(n_169),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_L g178 ( 
.A(n_168),
.B(n_169),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_SL g172 ( 
.A(n_173),
.B(n_175),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_SL g181 ( 
.A(n_182),
.B(n_196),
.Y(n_181)
);

NOR2xp33_ASAP7_75t_L g197 ( 
.A(n_182),
.B(n_196),
.Y(n_197)
);

XNOR2xp5_ASAP7_75t_L g182 ( 
.A(n_183),
.B(n_191),
.Y(n_182)
);

MAJIxp5_ASAP7_75t_L g199 ( 
.A(n_183),
.B(n_192),
.C(n_193),
.Y(n_199)
);

AOI22xp5_ASAP7_75t_L g183 ( 
.A1(n_184),
.A2(n_185),
.B1(n_189),
.B2(n_190),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_L g207 ( 
.A(n_184),
.B(n_190),
.Y(n_207)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_185),
.Y(n_184)
);

CKINVDCx5p33_ASAP7_75t_R g186 ( 
.A(n_187),
.Y(n_186)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_190),
.Y(n_189)
);

XNOR2xp5_ASAP7_75t_L g191 ( 
.A(n_192),
.B(n_193),
.Y(n_191)
);

CKINVDCx14_ASAP7_75t_R g209 ( 
.A(n_195),
.Y(n_209)
);

NOR2xp33_ASAP7_75t_L g198 ( 
.A(n_199),
.B(n_200),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_L g213 ( 
.A(n_199),
.B(n_200),
.Y(n_213)
);

OAI22xp5_ASAP7_75t_SL g200 ( 
.A1(n_201),
.A2(n_202),
.B1(n_205),
.B2(n_206),
.Y(n_200)
);

MAJIxp5_ASAP7_75t_L g217 ( 
.A(n_201),
.B(n_208),
.C(n_211),
.Y(n_217)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_202),
.Y(n_201)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_206),
.Y(n_205)
);

OAI22xp5_ASAP7_75t_SL g206 ( 
.A1(n_207),
.A2(n_208),
.B1(n_211),
.B2(n_212),
.Y(n_206)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_207),
.Y(n_211)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_208),
.Y(n_212)
);

NAND2xp5_ASAP7_75t_SL g214 ( 
.A(n_215),
.B(n_217),
.Y(n_214)
);

NOR2xp33_ASAP7_75t_L g218 ( 
.A(n_215),
.B(n_217),
.Y(n_218)
);

NAND2xp5_ASAP7_75t_L g220 ( 
.A(n_221),
.B(n_222),
.Y(n_220)
);

NOR2xp33_ASAP7_75t_L g240 ( 
.A(n_221),
.B(n_222),
.Y(n_240)
);

XNOR2xp5_ASAP7_75t_L g222 ( 
.A(n_223),
.B(n_239),
.Y(n_222)
);

XNOR2xp5_ASAP7_75t_L g223 ( 
.A(n_224),
.B(n_231),
.Y(n_223)
);

MAJIxp5_ASAP7_75t_L g242 ( 
.A(n_224),
.B(n_231),
.C(n_239),
.Y(n_242)
);

AOI22xp5_ASAP7_75t_L g224 ( 
.A1(n_225),
.A2(n_226),
.B1(n_227),
.B2(n_230),
.Y(n_224)
);

NAND2xp5_ASAP7_75t_L g253 ( 
.A(n_225),
.B(n_230),
.Y(n_253)
);

CKINVDCx20_ASAP7_75t_R g225 ( 
.A(n_226),
.Y(n_225)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_227),
.Y(n_230)
);

CKINVDCx20_ASAP7_75t_R g249 ( 
.A(n_229),
.Y(n_249)
);

XOR2xp5_ASAP7_75t_L g231 ( 
.A(n_232),
.B(n_233),
.Y(n_231)
);

MAJIxp5_ASAP7_75t_L g268 ( 
.A(n_232),
.B(n_234),
.C(n_236),
.Y(n_268)
);

XOR2xp5_ASAP7_75t_L g233 ( 
.A(n_234),
.B(n_236),
.Y(n_233)
);

CKINVDCx20_ASAP7_75t_R g256 ( 
.A(n_235),
.Y(n_256)
);

INVxp67_ASAP7_75t_L g264 ( 
.A(n_238),
.Y(n_264)
);

NOR2xp33_ASAP7_75t_L g241 ( 
.A(n_242),
.B(n_243),
.Y(n_241)
);

NAND2xp5_ASAP7_75t_SL g269 ( 
.A(n_242),
.B(n_243),
.Y(n_269)
);

XNOR2xp5_ASAP7_75t_L g243 ( 
.A(n_244),
.B(n_268),
.Y(n_243)
);

AOI22xp5_ASAP7_75t_L g244 ( 
.A1(n_245),
.A2(n_252),
.B1(n_266),
.B2(n_267),
.Y(n_244)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_245),
.Y(n_266)
);

MAJIxp5_ASAP7_75t_L g271 ( 
.A(n_245),
.B(n_267),
.C(n_268),
.Y(n_271)
);

OAI22xp5_ASAP7_75t_L g245 ( 
.A1(n_246),
.A2(n_247),
.B1(n_248),
.B2(n_251),
.Y(n_245)
);

AOI22xp5_ASAP7_75t_L g283 ( 
.A1(n_246),
.A2(n_247),
.B1(n_284),
.B2(n_285),
.Y(n_283)
);

OAI21xp5_ASAP7_75t_L g312 ( 
.A1(n_246),
.A2(n_281),
.B(n_285),
.Y(n_312)
);

CKINVDCx20_ASAP7_75t_R g246 ( 
.A(n_247),
.Y(n_246)
);

NAND2xp5_ASAP7_75t_L g282 ( 
.A(n_247),
.B(n_248),
.Y(n_282)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_248),
.Y(n_251)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_252),
.Y(n_267)
);

XNOR2xp5_ASAP7_75t_SL g252 ( 
.A(n_253),
.B(n_254),
.Y(n_252)
);

MAJIxp5_ASAP7_75t_L g293 ( 
.A(n_253),
.B(n_260),
.C(n_265),
.Y(n_293)
);

AOI22xp5_ASAP7_75t_L g254 ( 
.A1(n_255),
.A2(n_260),
.B1(n_261),
.B2(n_265),
.Y(n_254)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_255),
.Y(n_265)
);

NAND2xp5_ASAP7_75t_SL g349 ( 
.A(n_257),
.B(n_303),
.Y(n_349)
);

CKINVDCx20_ASAP7_75t_R g286 ( 
.A(n_258),
.Y(n_286)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_261),
.Y(n_260)
);

CKINVDCx16_ASAP7_75t_R g276 ( 
.A(n_262),
.Y(n_276)
);

NAND2xp5_ASAP7_75t_L g270 ( 
.A(n_271),
.B(n_272),
.Y(n_270)
);

NOR2xp33_ASAP7_75t_SL g296 ( 
.A(n_271),
.B(n_272),
.Y(n_296)
);

AOI22xp5_ASAP7_75t_SL g272 ( 
.A1(n_273),
.A2(n_293),
.B1(n_294),
.B2(n_295),
.Y(n_272)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_273),
.Y(n_294)
);

AOI22xp5_ASAP7_75t_L g273 ( 
.A1(n_274),
.A2(n_280),
.B1(n_291),
.B2(n_292),
.Y(n_273)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_274),
.Y(n_291)
);

OAI21xp33_ASAP7_75t_L g274 ( 
.A1(n_275),
.A2(n_278),
.B(n_279),
.Y(n_274)
);

NAND2xp5_ASAP7_75t_SL g279 ( 
.A(n_275),
.B(n_278),
.Y(n_279)
);

CKINVDCx14_ASAP7_75t_R g311 ( 
.A(n_279),
.Y(n_311)
);

AOI22xp5_ASAP7_75t_L g330 ( 
.A1(n_279),
.A2(n_299),
.B1(n_311),
.B2(n_331),
.Y(n_330)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_280),
.Y(n_292)
);

MAJIxp5_ASAP7_75t_L g328 ( 
.A(n_280),
.B(n_291),
.C(n_295),
.Y(n_328)
);

AOI22xp5_ASAP7_75t_L g280 ( 
.A1(n_281),
.A2(n_282),
.B1(n_283),
.B2(n_290),
.Y(n_280)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_282),
.Y(n_281)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_283),
.Y(n_290)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_285),
.Y(n_284)
);

CKINVDCx20_ASAP7_75t_R g341 ( 
.A(n_287),
.Y(n_341)
);

CKINVDCx16_ASAP7_75t_R g295 ( 
.A(n_293),
.Y(n_295)
);

NOR2xp33_ASAP7_75t_L g297 ( 
.A(n_298),
.B(n_313),
.Y(n_297)
);

NAND2xp5_ASAP7_75t_L g333 ( 
.A(n_298),
.B(n_313),
.Y(n_333)
);

MAJIxp5_ASAP7_75t_L g298 ( 
.A(n_299),
.B(n_311),
.C(n_312),
.Y(n_298)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_299),
.Y(n_331)
);

AOI22xp5_ASAP7_75t_L g299 ( 
.A1(n_300),
.A2(n_301),
.B1(n_304),
.B2(n_305),
.Y(n_299)
);

AOI22xp5_ASAP7_75t_L g314 ( 
.A1(n_300),
.A2(n_301),
.B1(n_315),
.B2(n_316),
.Y(n_314)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_301),
.Y(n_300)
);

MAJIxp5_ASAP7_75t_L g326 ( 
.A(n_301),
.B(n_306),
.C(n_310),
.Y(n_326)
);

MAJIxp5_ASAP7_75t_L g335 ( 
.A(n_301),
.B(n_316),
.C(n_326),
.Y(n_335)
);

CKINVDCx20_ASAP7_75t_R g321 ( 
.A(n_302),
.Y(n_321)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_305),
.Y(n_304)
);

OAI22xp5_ASAP7_75t_SL g305 ( 
.A1(n_306),
.A2(n_307),
.B1(n_309),
.B2(n_310),
.Y(n_305)
);

AOI22xp5_ASAP7_75t_SL g317 ( 
.A1(n_306),
.A2(n_307),
.B1(n_318),
.B2(n_319),
.Y(n_317)
);

CKINVDCx16_ASAP7_75t_R g306 ( 
.A(n_307),
.Y(n_306)
);

MAJIxp5_ASAP7_75t_L g345 ( 
.A(n_307),
.B(n_318),
.C(n_320),
.Y(n_345)
);

CKINVDCx20_ASAP7_75t_R g309 ( 
.A(n_310),
.Y(n_309)
);

XOR2xp5_ASAP7_75t_L g329 ( 
.A(n_312),
.B(n_330),
.Y(n_329)
);

XNOR2xp5_ASAP7_75t_L g313 ( 
.A(n_314),
.B(n_326),
.Y(n_313)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_316),
.Y(n_315)
);

XOR2xp5_ASAP7_75t_L g316 ( 
.A(n_317),
.B(n_320),
.Y(n_316)
);

CKINVDCx20_ASAP7_75t_R g318 ( 
.A(n_319),
.Y(n_318)
);

INVx8_ASAP7_75t_L g323 ( 
.A(n_324),
.Y(n_323)
);

INVx8_ASAP7_75t_L g324 ( 
.A(n_325),
.Y(n_324)
);

NOR2xp33_ASAP7_75t_L g327 ( 
.A(n_328),
.B(n_329),
.Y(n_327)
);

NAND2xp5_ASAP7_75t_SL g332 ( 
.A(n_328),
.B(n_329),
.Y(n_332)
);

NAND2xp5_ASAP7_75t_SL g334 ( 
.A(n_335),
.B(n_336),
.Y(n_334)
);

NOR2xp33_ASAP7_75t_L g346 ( 
.A(n_335),
.B(n_336),
.Y(n_346)
);

AOI22xp5_ASAP7_75t_L g336 ( 
.A1(n_337),
.A2(n_338),
.B1(n_344),
.B2(n_345),
.Y(n_336)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_338),
.Y(n_337)
);

AOI22xp5_ASAP7_75t_L g338 ( 
.A1(n_339),
.A2(n_340),
.B1(n_342),
.B2(n_343),
.Y(n_338)
);

CKINVDCx20_ASAP7_75t_R g342 ( 
.A(n_339),
.Y(n_342)
);

CKINVDCx20_ASAP7_75t_R g343 ( 
.A(n_340),
.Y(n_343)
);

MAJIxp5_ASAP7_75t_L g351 ( 
.A(n_340),
.B(n_342),
.C(n_344),
.Y(n_351)
);

CKINVDCx20_ASAP7_75t_R g344 ( 
.A(n_345),
.Y(n_344)
);

INVxp67_ASAP7_75t_L g347 ( 
.A(n_348),
.Y(n_347)
);

NAND2xp5_ASAP7_75t_L g348 ( 
.A(n_349),
.B(n_350),
.Y(n_348)
);

CKINVDCx20_ASAP7_75t_R g353 ( 
.A(n_349),
.Y(n_353)
);

INVx1_ASAP7_75t_L g350 ( 
.A(n_351),
.Y(n_350)
);

NAND2xp5_ASAP7_75t_SL g352 ( 
.A(n_351),
.B(n_353),
.Y(n_352)
);


endmodule