module fake_jpeg_12522_n_132 (n_13, n_21, n_33, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_19, n_18, n_20, n_35, n_4, n_34, n_30, n_39, n_16, n_3, n_0, n_24, n_28, n_38, n_26, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_12, n_32, n_8, n_15, n_7, n_132);

input n_13;
input n_21;
input n_33;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_35;
input n_4;
input n_34;
input n_30;
input n_39;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_132;

wire n_117;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_73;
wire n_84;
wire n_59;
wire n_98;
wire n_65;
wire n_110;
wire n_42;
wire n_49;
wire n_76;
wire n_127;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_103;
wire n_50;
wire n_124;
wire n_57;
wire n_119;
wire n_69;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_106;
wire n_111;
wire n_44;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_67;
wire n_53;
wire n_54;
wire n_93;
wire n_91;
wire n_101;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_97;
wire n_62;
wire n_120;
wire n_43;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_96;

BUFx10_ASAP7_75t_L g40 ( 
.A(n_9),
.Y(n_40)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_20),
.Y(n_41)
);

BUFx3_ASAP7_75t_L g42 ( 
.A(n_6),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_32),
.Y(n_43)
);

INVx5_ASAP7_75t_L g44 ( 
.A(n_38),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_8),
.Y(n_45)
);

INVx5_ASAP7_75t_L g46 ( 
.A(n_35),
.Y(n_46)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_36),
.Y(n_47)
);

INVx4_ASAP7_75t_L g48 ( 
.A(n_37),
.Y(n_48)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_25),
.Y(n_49)
);

BUFx2_ASAP7_75t_L g50 ( 
.A(n_1),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g51 ( 
.A(n_4),
.B(n_16),
.Y(n_51)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_1),
.Y(n_52)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_11),
.Y(n_53)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_5),
.Y(n_54)
);

INVx2_ASAP7_75t_R g55 ( 
.A(n_21),
.Y(n_55)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_22),
.Y(n_56)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_52),
.Y(n_57)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_57),
.Y(n_80)
);

INVx4_ASAP7_75t_L g58 ( 
.A(n_42),
.Y(n_58)
);

INVx6_ASAP7_75t_L g78 ( 
.A(n_58),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_55),
.B(n_54),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_SL g76 ( 
.A(n_59),
.B(n_43),
.Y(n_76)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_48),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g79 ( 
.A(n_60),
.Y(n_79)
);

CKINVDCx20_ASAP7_75t_R g61 ( 
.A(n_51),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_61),
.B(n_64),
.Y(n_67)
);

INVx2_ASAP7_75t_L g62 ( 
.A(n_50),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_L g68 ( 
.A(n_62),
.B(n_40),
.Y(n_68)
);

BUFx12f_ASAP7_75t_L g63 ( 
.A(n_42),
.Y(n_63)
);

BUFx16f_ASAP7_75t_L g77 ( 
.A(n_63),
.Y(n_77)
);

INVx2_ASAP7_75t_SL g64 ( 
.A(n_40),
.Y(n_64)
);

BUFx3_ASAP7_75t_L g65 ( 
.A(n_50),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_65),
.B(n_46),
.Y(n_72)
);

INVx11_ASAP7_75t_L g66 ( 
.A(n_40),
.Y(n_66)
);

CKINVDCx20_ASAP7_75t_R g75 ( 
.A(n_66),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_L g91 ( 
.A(n_68),
.B(n_69),
.Y(n_91)
);

OR2x2_ASAP7_75t_SL g69 ( 
.A(n_58),
.B(n_55),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_L g70 ( 
.A(n_64),
.B(n_45),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_L g96 ( 
.A(n_70),
.B(n_73),
.Y(n_96)
);

OAI22xp33_ASAP7_75t_SL g71 ( 
.A1(n_65),
.A2(n_48),
.B1(n_56),
.B2(n_49),
.Y(n_71)
);

OAI22xp33_ASAP7_75t_SL g97 ( 
.A1(n_71),
.A2(n_2),
.B1(n_3),
.B2(n_4),
.Y(n_97)
);

INVxp67_ASAP7_75t_L g87 ( 
.A(n_72),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_L g73 ( 
.A(n_60),
.B(n_56),
.Y(n_73)
);

AOI22xp33_ASAP7_75t_SL g74 ( 
.A1(n_66),
.A2(n_46),
.B1(n_44),
.B2(n_53),
.Y(n_74)
);

AOI21xp5_ASAP7_75t_L g83 ( 
.A1(n_74),
.A2(n_63),
.B(n_47),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_76),
.B(n_41),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_81),
.B(n_82),
.Y(n_110)
);

O2A1O1Ixp33_ASAP7_75t_SL g82 ( 
.A1(n_71),
.A2(n_63),
.B(n_44),
.C(n_18),
.Y(n_82)
);

CKINVDCx16_ASAP7_75t_R g100 ( 
.A(n_83),
.Y(n_100)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_80),
.Y(n_84)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_84),
.Y(n_101)
);

OA22x2_ASAP7_75t_L g85 ( 
.A1(n_69),
.A2(n_15),
.B1(n_34),
.B2(n_33),
.Y(n_85)
);

OAI22xp5_ASAP7_75t_SL g98 ( 
.A1(n_85),
.A2(n_2),
.B1(n_3),
.B2(n_5),
.Y(n_98)
);

BUFx6f_ASAP7_75t_L g86 ( 
.A(n_79),
.Y(n_86)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_86),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_67),
.B(n_0),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_L g109 ( 
.A(n_88),
.B(n_90),
.Y(n_109)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_78),
.Y(n_89)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_89),
.Y(n_104)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_78),
.Y(n_90)
);

INVx2_ASAP7_75t_L g92 ( 
.A(n_79),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_SL g106 ( 
.A(n_92),
.B(n_93),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_75),
.B(n_0),
.Y(n_93)
);

OAI22xp5_ASAP7_75t_L g94 ( 
.A1(n_74),
.A2(n_14),
.B1(n_31),
.B2(n_30),
.Y(n_94)
);

AOI22xp5_ASAP7_75t_L g105 ( 
.A1(n_94),
.A2(n_97),
.B1(n_6),
.B2(n_7),
.Y(n_105)
);

INVx1_ASAP7_75t_SL g95 ( 
.A(n_77),
.Y(n_95)
);

CKINVDCx16_ASAP7_75t_R g108 ( 
.A(n_95),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_L g116 ( 
.A(n_98),
.B(n_111),
.Y(n_116)
);

OAI22xp5_ASAP7_75t_SL g99 ( 
.A1(n_91),
.A2(n_77),
.B1(n_7),
.B2(n_8),
.Y(n_99)
);

OAI22xp5_ASAP7_75t_L g115 ( 
.A1(n_99),
.A2(n_103),
.B1(n_105),
.B2(n_107),
.Y(n_115)
);

OAI22xp5_ASAP7_75t_SL g103 ( 
.A1(n_96),
.A2(n_87),
.B1(n_97),
.B2(n_82),
.Y(n_103)
);

OAI22xp5_ASAP7_75t_SL g107 ( 
.A1(n_87),
.A2(n_77),
.B1(n_10),
.B2(n_9),
.Y(n_107)
);

MAJIxp5_ASAP7_75t_L g111 ( 
.A(n_85),
.B(n_95),
.C(n_86),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_SL g112 ( 
.A(n_85),
.B(n_10),
.Y(n_112)
);

INVxp67_ASAP7_75t_L g113 ( 
.A(n_112),
.Y(n_113)
);

CKINVDCx20_ASAP7_75t_R g114 ( 
.A(n_109),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_SL g123 ( 
.A(n_114),
.B(n_117),
.Y(n_123)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_104),
.Y(n_117)
);

AO22x1_ASAP7_75t_L g118 ( 
.A1(n_100),
.A2(n_39),
.B1(n_13),
.B2(n_17),
.Y(n_118)
);

OAI21xp5_ASAP7_75t_L g121 ( 
.A1(n_118),
.A2(n_119),
.B(n_120),
.Y(n_121)
);

INVx3_ASAP7_75t_L g119 ( 
.A(n_101),
.Y(n_119)
);

AOI21xp5_ASAP7_75t_L g120 ( 
.A1(n_111),
.A2(n_110),
.B(n_106),
.Y(n_120)
);

AOI22xp5_ASAP7_75t_L g122 ( 
.A1(n_115),
.A2(n_99),
.B1(n_107),
.B2(n_98),
.Y(n_122)
);

OAI22xp5_ASAP7_75t_L g126 ( 
.A1(n_122),
.A2(n_105),
.B1(n_102),
.B2(n_108),
.Y(n_126)
);

OAI21xp5_ASAP7_75t_L g124 ( 
.A1(n_113),
.A2(n_116),
.B(n_118),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_SL g125 ( 
.A(n_124),
.B(n_113),
.Y(n_125)
);

BUFx4f_ASAP7_75t_SL g127 ( 
.A(n_125),
.Y(n_127)
);

NAND2x1p5_ASAP7_75t_L g128 ( 
.A(n_127),
.B(n_123),
.Y(n_128)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_128),
.Y(n_129)
);

AOI332xp33_ASAP7_75t_L g130 ( 
.A1(n_129),
.A2(n_121),
.A3(n_126),
.B1(n_23),
.B2(n_24),
.B3(n_26),
.C1(n_12),
.C2(n_28),
.Y(n_130)
);

MAJIxp5_ASAP7_75t_L g131 ( 
.A(n_130),
.B(n_19),
.C(n_27),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_L g132 ( 
.A(n_131),
.B(n_29),
.Y(n_132)
);


endmodule