module fake_jpeg_607_n_220 (n_13, n_21, n_33, n_1, n_45, n_10, n_23, n_27, n_6, n_22, n_47, n_51, n_14, n_40, n_19, n_18, n_20, n_35, n_48, n_52, n_46, n_41, n_4, n_34, n_30, n_39, n_42, n_16, n_49, n_3, n_0, n_24, n_28, n_38, n_26, n_44, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_43, n_50, n_12, n_32, n_8, n_15, n_7, n_220);

input n_13;
input n_21;
input n_33;
input n_1;
input n_45;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_47;
input n_51;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_48;
input n_52;
input n_46;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_42;
input n_16;
input n_49;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_44;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_43;
input n_50;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_220;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_64;
wire n_55;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_84;
wire n_59;
wire n_98;
wire n_178;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_127;
wire n_76;
wire n_154;
wire n_205;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_155;
wire n_207;
wire n_103;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_57;
wire n_171;
wire n_119;
wire n_69;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_143;
wire n_202;
wire n_122;
wire n_75;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_145;
wire n_108;
wire n_68;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_131;
wire n_56;
wire n_212;
wire n_211;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_216;
wire n_217;
wire n_184;
wire n_53;
wire n_91;
wire n_54;
wire n_93;
wire n_161;
wire n_209;
wire n_208;
wire n_138;
wire n_101;
wire n_210;
wire n_149;
wire n_157;
wire n_87;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

INVx4_ASAP7_75t_L g53 ( 
.A(n_14),
.Y(n_53)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_52),
.Y(n_54)
);

INVx6_ASAP7_75t_L g55 ( 
.A(n_16),
.Y(n_55)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_38),
.Y(n_56)
);

BUFx5_ASAP7_75t_L g57 ( 
.A(n_25),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_37),
.Y(n_58)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_0),
.Y(n_59)
);

INVx4_ASAP7_75t_L g60 ( 
.A(n_9),
.Y(n_60)
);

INVx6_ASAP7_75t_L g61 ( 
.A(n_22),
.Y(n_61)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_39),
.Y(n_62)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_17),
.Y(n_63)
);

CKINVDCx20_ASAP7_75t_R g64 ( 
.A(n_22),
.Y(n_64)
);

BUFx12_ASAP7_75t_L g65 ( 
.A(n_6),
.Y(n_65)
);

BUFx5_ASAP7_75t_L g66 ( 
.A(n_0),
.Y(n_66)
);

CKINVDCx20_ASAP7_75t_R g67 ( 
.A(n_34),
.Y(n_67)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_28),
.Y(n_68)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_2),
.Y(n_69)
);

BUFx10_ASAP7_75t_L g70 ( 
.A(n_11),
.Y(n_70)
);

CKINVDCx20_ASAP7_75t_R g71 ( 
.A(n_50),
.Y(n_71)
);

BUFx12f_ASAP7_75t_L g72 ( 
.A(n_48),
.Y(n_72)
);

CKINVDCx20_ASAP7_75t_R g73 ( 
.A(n_10),
.Y(n_73)
);

BUFx12f_ASAP7_75t_L g74 ( 
.A(n_46),
.Y(n_74)
);

CKINVDCx20_ASAP7_75t_R g75 ( 
.A(n_27),
.Y(n_75)
);

CKINVDCx20_ASAP7_75t_R g76 ( 
.A(n_26),
.Y(n_76)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_24),
.Y(n_77)
);

BUFx5_ASAP7_75t_L g78 ( 
.A(n_6),
.Y(n_78)
);

BUFx12f_ASAP7_75t_L g79 ( 
.A(n_65),
.Y(n_79)
);

INVx2_ASAP7_75t_SL g96 ( 
.A(n_79),
.Y(n_96)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_68),
.Y(n_80)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_80),
.Y(n_89)
);

INVx6_ASAP7_75t_L g81 ( 
.A(n_58),
.Y(n_81)
);

INVx2_ASAP7_75t_L g91 ( 
.A(n_81),
.Y(n_91)
);

BUFx5_ASAP7_75t_L g82 ( 
.A(n_56),
.Y(n_82)
);

BUFx5_ASAP7_75t_L g94 ( 
.A(n_82),
.Y(n_94)
);

INVx2_ASAP7_75t_L g83 ( 
.A(n_56),
.Y(n_83)
);

INVx2_ASAP7_75t_L g93 ( 
.A(n_83),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_64),
.B(n_1),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_84),
.B(n_54),
.Y(n_97)
);

INVx5_ASAP7_75t_L g85 ( 
.A(n_72),
.Y(n_85)
);

INVx3_ASAP7_75t_L g90 ( 
.A(n_85),
.Y(n_90)
);

INVx11_ASAP7_75t_L g86 ( 
.A(n_72),
.Y(n_86)
);

CKINVDCx6p67_ASAP7_75t_R g95 ( 
.A(n_86),
.Y(n_95)
);

BUFx12f_ASAP7_75t_L g87 ( 
.A(n_65),
.Y(n_87)
);

INVx2_ASAP7_75t_L g102 ( 
.A(n_87),
.Y(n_102)
);

INVx2_ASAP7_75t_L g88 ( 
.A(n_53),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_88),
.B(n_72),
.Y(n_103)
);

NOR2x1_ASAP7_75t_L g92 ( 
.A(n_88),
.B(n_63),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_92),
.B(n_97),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_80),
.B(n_69),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g118 ( 
.A(n_98),
.B(n_100),
.Y(n_118)
);

AOI22xp5_ASAP7_75t_L g99 ( 
.A1(n_83),
.A2(n_53),
.B1(n_60),
.B2(n_58),
.Y(n_99)
);

OAI22xp5_ASAP7_75t_SL g111 ( 
.A1(n_99),
.A2(n_55),
.B1(n_61),
.B2(n_60),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_79),
.B(n_59),
.Y(n_100)
);

CKINVDCx12_ASAP7_75t_R g101 ( 
.A(n_79),
.Y(n_101)
);

INVxp67_ASAP7_75t_L g104 ( 
.A(n_101),
.Y(n_104)
);

AND2x2_ASAP7_75t_L g123 ( 
.A(n_103),
.B(n_87),
.Y(n_123)
);

INVx3_ASAP7_75t_L g105 ( 
.A(n_90),
.Y(n_105)
);

INVx2_ASAP7_75t_L g130 ( 
.A(n_105),
.Y(n_130)
);

O2A1O1Ixp33_ASAP7_75t_L g106 ( 
.A1(n_92),
.A2(n_86),
.B(n_85),
.C(n_82),
.Y(n_106)
);

INVxp67_ASAP7_75t_L g139 ( 
.A(n_106),
.Y(n_139)
);

OAI22xp5_ASAP7_75t_L g107 ( 
.A1(n_99),
.A2(n_81),
.B1(n_55),
.B2(n_61),
.Y(n_107)
);

AOI22xp33_ASAP7_75t_L g141 ( 
.A1(n_107),
.A2(n_66),
.B1(n_57),
.B2(n_94),
.Y(n_141)
);

INVx4_ASAP7_75t_L g108 ( 
.A(n_90),
.Y(n_108)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_108),
.Y(n_126)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_89),
.Y(n_109)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_109),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_L g147 ( 
.A(n_111),
.B(n_117),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_SL g112 ( 
.A(n_93),
.B(n_77),
.Y(n_112)
);

NAND3xp33_ASAP7_75t_L g135 ( 
.A(n_112),
.B(n_122),
.C(n_123),
.Y(n_135)
);

OR2x4_ASAP7_75t_L g113 ( 
.A(n_95),
.B(n_70),
.Y(n_113)
);

OR2x2_ASAP7_75t_L g129 ( 
.A(n_113),
.B(n_70),
.Y(n_129)
);

INVx2_ASAP7_75t_L g114 ( 
.A(n_91),
.Y(n_114)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_114),
.Y(n_136)
);

AOI22xp33_ASAP7_75t_SL g115 ( 
.A1(n_96),
.A2(n_63),
.B1(n_59),
.B2(n_74),
.Y(n_115)
);

OAI22xp33_ASAP7_75t_SL g145 ( 
.A1(n_115),
.A2(n_5),
.B1(n_7),
.B2(n_8),
.Y(n_145)
);

INVx2_ASAP7_75t_L g116 ( 
.A(n_91),
.Y(n_116)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_116),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_93),
.B(n_62),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_L g119 ( 
.A(n_96),
.B(n_73),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_SL g138 ( 
.A(n_119),
.B(n_2),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_L g120 ( 
.A(n_102),
.B(n_62),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_120),
.B(n_75),
.Y(n_124)
);

OAI22xp5_ASAP7_75t_SL g121 ( 
.A1(n_102),
.A2(n_74),
.B1(n_77),
.B2(n_87),
.Y(n_121)
);

OAI22xp5_ASAP7_75t_SL g125 ( 
.A1(n_121),
.A2(n_79),
.B1(n_87),
.B2(n_95),
.Y(n_125)
);

CKINVDCx20_ASAP7_75t_R g122 ( 
.A(n_95),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_SL g153 ( 
.A(n_124),
.B(n_144),
.Y(n_153)
);

AOI22xp5_ASAP7_75t_L g159 ( 
.A1(n_125),
.A2(n_132),
.B1(n_142),
.B2(n_7),
.Y(n_159)
);

OA22x2_ASAP7_75t_SL g127 ( 
.A1(n_113),
.A2(n_95),
.B1(n_94),
.B2(n_70),
.Y(n_127)
);

OAI21xp33_ASAP7_75t_L g154 ( 
.A1(n_127),
.A2(n_40),
.B(n_47),
.Y(n_154)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_118),
.B(n_67),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_SL g161 ( 
.A(n_128),
.B(n_133),
.Y(n_161)
);

AND2x2_ASAP7_75t_L g163 ( 
.A(n_129),
.B(n_137),
.Y(n_163)
);

MAJIxp5_ASAP7_75t_L g131 ( 
.A(n_123),
.B(n_76),
.C(n_71),
.Y(n_131)
);

MAJIxp5_ASAP7_75t_L g167 ( 
.A(n_131),
.B(n_12),
.C(n_13),
.Y(n_167)
);

OAI22xp5_ASAP7_75t_SL g132 ( 
.A1(n_111),
.A2(n_74),
.B1(n_70),
.B2(n_78),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_L g133 ( 
.A(n_110),
.B(n_1),
.Y(n_133)
);

OAI32xp33_ASAP7_75t_L g137 ( 
.A1(n_106),
.A2(n_78),
.A3(n_66),
.B1(n_57),
.B2(n_65),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_SL g172 ( 
.A(n_138),
.B(n_140),
.Y(n_172)
);

NOR2xp33_ASAP7_75t_L g140 ( 
.A(n_104),
.B(n_3),
.Y(n_140)
);

OAI22xp5_ASAP7_75t_L g151 ( 
.A1(n_141),
.A2(n_108),
.B1(n_121),
.B2(n_116),
.Y(n_151)
);

OAI22xp5_ASAP7_75t_SL g142 ( 
.A1(n_123),
.A2(n_3),
.B1(n_4),
.B2(n_5),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_L g143 ( 
.A(n_114),
.B(n_51),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_L g157 ( 
.A(n_143),
.B(n_145),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_SL g144 ( 
.A(n_105),
.B(n_4),
.Y(n_144)
);

NOR2xp33_ASAP7_75t_L g148 ( 
.A(n_131),
.B(n_104),
.Y(n_148)
);

NOR2xp33_ASAP7_75t_L g177 ( 
.A(n_148),
.B(n_156),
.Y(n_177)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_136),
.Y(n_149)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_149),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_L g150 ( 
.A(n_147),
.B(n_143),
.Y(n_150)
);

A2O1A1O1Ixp25_ASAP7_75t_L g181 ( 
.A1(n_150),
.A2(n_127),
.B(n_32),
.C(n_33),
.D(n_45),
.Y(n_181)
);

AOI22xp5_ASAP7_75t_L g185 ( 
.A1(n_151),
.A2(n_159),
.B1(n_15),
.B2(n_16),
.Y(n_185)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_146),
.Y(n_152)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_152),
.Y(n_176)
);

OAI21xp5_ASAP7_75t_L g187 ( 
.A1(n_154),
.A2(n_173),
.B(n_17),
.Y(n_187)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_134),
.Y(n_155)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_155),
.Y(n_178)
);

CKINVDCx12_ASAP7_75t_R g156 ( 
.A(n_135),
.Y(n_156)
);

XNOR2xp5_ASAP7_75t_SL g158 ( 
.A(n_137),
.B(n_49),
.Y(n_158)
);

XNOR2xp5_ASAP7_75t_L g189 ( 
.A(n_158),
.B(n_165),
.Y(n_189)
);

AOI21xp5_ASAP7_75t_L g160 ( 
.A1(n_139),
.A2(n_8),
.B(n_9),
.Y(n_160)
);

OAI21xp5_ASAP7_75t_L g183 ( 
.A1(n_160),
.A2(n_14),
.B(n_15),
.Y(n_183)
);

NOR2xp33_ASAP7_75t_L g162 ( 
.A(n_142),
.B(n_10),
.Y(n_162)
);

NOR2xp33_ASAP7_75t_L g179 ( 
.A(n_162),
.B(n_164),
.Y(n_179)
);

NOR2xp33_ASAP7_75t_L g164 ( 
.A(n_126),
.B(n_11),
.Y(n_164)
);

XNOR2xp5_ASAP7_75t_SL g165 ( 
.A(n_129),
.B(n_29),
.Y(n_165)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_130),
.Y(n_166)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_166),
.Y(n_180)
);

NOR2xp33_ASAP7_75t_L g184 ( 
.A(n_167),
.B(n_168),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_SL g168 ( 
.A(n_130),
.B(n_12),
.Y(n_168)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_125),
.Y(n_169)
);

NOR2xp33_ASAP7_75t_L g186 ( 
.A(n_169),
.B(n_170),
.Y(n_186)
);

NOR2xp33_ASAP7_75t_L g170 ( 
.A(n_139),
.B(n_13),
.Y(n_170)
);

XNOR2xp5_ASAP7_75t_L g171 ( 
.A(n_132),
.B(n_31),
.Y(n_171)
);

MAJIxp5_ASAP7_75t_L g182 ( 
.A(n_171),
.B(n_44),
.C(n_43),
.Y(n_182)
);

INVx1_ASAP7_75t_SL g173 ( 
.A(n_127),
.Y(n_173)
);

INVx3_ASAP7_75t_SL g175 ( 
.A(n_163),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_L g192 ( 
.A(n_175),
.B(n_181),
.Y(n_192)
);

MAJIxp5_ASAP7_75t_L g197 ( 
.A(n_182),
.B(n_167),
.C(n_165),
.Y(n_197)
);

AOI21xp5_ASAP7_75t_L g199 ( 
.A1(n_183),
.A2(n_191),
.B(n_157),
.Y(n_199)
);

OAI22xp5_ASAP7_75t_L g194 ( 
.A1(n_185),
.A2(n_187),
.B1(n_190),
.B2(n_154),
.Y(n_194)
);

INVxp67_ASAP7_75t_L g188 ( 
.A(n_160),
.Y(n_188)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_188),
.Y(n_193)
);

AOI22xp5_ASAP7_75t_L g190 ( 
.A1(n_163),
.A2(n_18),
.B1(n_19),
.B2(n_20),
.Y(n_190)
);

A2O1A1O1Ixp25_ASAP7_75t_L g191 ( 
.A1(n_150),
.A2(n_30),
.B(n_41),
.C(n_36),
.D(n_35),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_L g207 ( 
.A(n_194),
.B(n_195),
.Y(n_207)
);

NOR2xp33_ASAP7_75t_L g195 ( 
.A(n_184),
.B(n_172),
.Y(n_195)
);

CKINVDCx20_ASAP7_75t_R g196 ( 
.A(n_178),
.Y(n_196)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_196),
.Y(n_205)
);

MAJIxp5_ASAP7_75t_L g203 ( 
.A(n_197),
.B(n_177),
.C(n_153),
.Y(n_203)
);

MAJIxp5_ASAP7_75t_L g198 ( 
.A(n_175),
.B(n_173),
.C(n_158),
.Y(n_198)
);

MAJIxp5_ASAP7_75t_L g202 ( 
.A(n_198),
.B(n_200),
.C(n_189),
.Y(n_202)
);

CKINVDCx16_ASAP7_75t_R g201 ( 
.A(n_199),
.Y(n_201)
);

MAJIxp5_ASAP7_75t_L g200 ( 
.A(n_189),
.B(n_171),
.C(n_159),
.Y(n_200)
);

XNOR2xp5_ASAP7_75t_L g209 ( 
.A(n_202),
.B(n_203),
.Y(n_209)
);

XNOR2x1_ASAP7_75t_L g204 ( 
.A(n_198),
.B(n_188),
.Y(n_204)
);

AOI21xp5_ASAP7_75t_L g211 ( 
.A1(n_204),
.A2(n_200),
.B(n_191),
.Y(n_211)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_193),
.Y(n_206)
);

AOI22xp5_ASAP7_75t_L g210 ( 
.A1(n_206),
.A2(n_176),
.B1(n_174),
.B2(n_186),
.Y(n_210)
);

OAI21xp5_ASAP7_75t_L g208 ( 
.A1(n_207),
.A2(n_192),
.B(n_181),
.Y(n_208)
);

MAJIxp5_ASAP7_75t_L g213 ( 
.A(n_208),
.B(n_211),
.C(n_202),
.Y(n_213)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_210),
.Y(n_212)
);

NOR2xp33_ASAP7_75t_SL g215 ( 
.A(n_213),
.B(n_182),
.Y(n_215)
);

AOI322xp5_ASAP7_75t_L g214 ( 
.A1(n_212),
.A2(n_201),
.A3(n_204),
.B1(n_205),
.B2(n_179),
.C1(n_209),
.C2(n_180),
.Y(n_214)
);

OAI21xp5_ASAP7_75t_L g216 ( 
.A1(n_214),
.A2(n_215),
.B(n_161),
.Y(n_216)
);

OR2x2_ASAP7_75t_L g217 ( 
.A(n_216),
.B(n_183),
.Y(n_217)
);

AOI322xp5_ASAP7_75t_L g218 ( 
.A1(n_217),
.A2(n_42),
.A3(n_19),
.B1(n_20),
.B2(n_21),
.C1(n_23),
.C2(n_18),
.Y(n_218)
);

NAND2xp5_ASAP7_75t_L g219 ( 
.A(n_218),
.B(n_21),
.Y(n_219)
);

NAND2x1_ASAP7_75t_L g220 ( 
.A(n_219),
.B(n_23),
.Y(n_220)
);


endmodule