module real_jpeg_18681_n_18 (n_17, n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_16, n_3, n_10, n_9, n_18);

input n_17;
input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_16;
input n_3;
input n_10;
input n_9;

output n_18;

wire n_384;
wire n_37;
wire n_430;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_460;
wire n_300;
wire n_415;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_518;
wire n_446;
wire n_199;
wire n_535;
wire n_95;
wire n_541;
wire n_441;
wire n_557;
wire n_238;
wire n_67;
wire n_350;
wire n_235;
wire n_107;
wire n_498;
wire n_369;
wire n_471;
wire n_376;
wire n_354;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_553;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_490;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_355;
wire n_123;
wire n_463;
wire n_425;
wire n_455;
wire n_462;
wire n_50;
wire n_409;
wire n_485;
wire n_186;
wire n_137;
wire n_491;
wire n_72;
wire n_440;
wire n_171;
wire n_151;
wire n_272;
wire n_461;
wire n_198;
wire n_203;
wire n_500;
wire n_23;
wire n_362;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_339;
wire n_326;
wire n_80;
wire n_30;
wire n_332;
wire n_149;
wire n_366;
wire n_328;
wire n_456;
wire n_259;
wire n_556;
wire n_57;
wire n_507;
wire n_157;
wire n_84;
wire n_560;
wire n_538;
wire n_527;
wire n_55;
wire n_499;
wire n_58;
wire n_52;
wire n_466;
wire n_353;
wire n_453;
wire n_551;
wire n_230;
wire n_417;
wire n_428;
wire n_128;
wire n_202;
wire n_216;
wire n_483;
wire n_367;
wire n_127;
wire n_365;
wire n_356;
wire n_464;
wire n_423;
wire n_36;
wire n_102;
wire n_81;
wire n_101;
wire n_422;
wire n_317;
wire n_506;
wire n_108;
wire n_550;
wire n_233;
wire n_73;
wire n_532;
wire n_348;
wire n_516;
wire n_473;
wire n_252;
wire n_363;
wire n_310;
wire n_345;
wire n_78;
wire n_83;
wire n_288;
wire n_525;
wire n_221;
wire n_393;
wire n_489;
wire n_104;
wire n_153;
wire n_443;
wire n_337;
wire n_544;
wire n_131;
wire n_439;
wire n_517;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_469;
wire n_378;
wire n_200;
wire n_432;
wire n_465;
wire n_335;
wire n_214;
wire n_113;
wire n_543;
wire n_251;
wire n_459;
wire n_139;
wire n_33;
wire n_175;
wire n_338;
wire n_488;
wire n_156;
wire n_387;
wire n_434;
wire n_66;
wire n_305;
wire n_505;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_390;
wire n_77;
wire n_399;
wire n_219;
wire n_372;
wire n_470;
wire n_122;
wire n_19;
wire n_262;
wire n_334;
wire n_383;
wire n_246;
wire n_523;
wire n_21;
wire n_476;
wire n_529;
wire n_69;
wire n_31;
wire n_426;
wire n_154;
wire n_495;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_371;
wire n_410;
wire n_421;
wire n_195;
wire n_110;
wire n_533;
wire n_289;
wire n_117;
wire n_193;
wire n_382;
wire n_411;
wire n_20;
wire n_278;
wire n_314;
wire n_103;
wire n_559;
wire n_232;
wire n_448;
wire n_212;
wire n_284;
wire n_402;
wire n_478;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_452;
wire n_213;
wire n_511;
wire n_524;
wire n_25;
wire n_480;
wire n_542;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_515;
wire n_89;
wire n_407;
wire n_419;
wire n_386;
wire n_521;
wire n_341;
wire n_331;
wire n_49;
wire n_514;
wire n_68;
wire n_497;
wire n_395;
wire n_146;
wire n_496;
wire n_323;
wire n_166;
wire n_176;
wire n_215;
wire n_286;
wire n_312;
wire n_325;
wire n_316;
wire n_307;
wire n_161;
wire n_207;
wire n_526;
wire n_431;
wire n_420;
wire n_357;
wire n_237;
wire n_445;
wire n_173;
wire n_115;
wire n_474;
wire n_184;
wire n_164;
wire n_380;
wire n_414;
wire n_140;
wire n_126;
wire n_342;
wire n_120;
wire n_155;
wire n_412;
wire n_405;
wire n_548;
wire n_319;
wire n_93;
wire n_487;
wire n_242;
wire n_493;
wire n_142;
wire n_522;
wire n_397;
wire n_76;
wire n_403;
wire n_79;
wire n_282;
wire n_147;
wire n_359;
wire n_265;
wire n_231;
wire n_44;
wire n_482;
wire n_208;
wire n_162;
wire n_449;
wire n_106;
wire n_172;
wire n_546;
wire n_285;
wire n_531;
wire n_112;
wire n_554;
wire n_508;
wire n_145;
wire n_266;
wire n_377;
wire n_109;
wire n_503;
wire n_391;
wire n_427;
wire n_401;
wire n_536;
wire n_148;
wire n_373;
wire n_558;
wire n_510;
wire n_396;
wire n_501;
wire n_392;
wire n_375;
wire n_196;
wire n_330;
wire n_298;
wire n_333;
wire n_450;
wire n_492;
wire n_152;
wire n_270;
wire n_159;
wire n_429;
wire n_347;
wire n_183;
wire n_248;
wire n_192;
wire n_537;
wire n_318;
wire n_90;
wire n_336;
wire n_258;
wire n_458;
wire n_150;
wire n_41;
wire n_74;
wire n_475;
wire n_404;
wire n_158;
wire n_204;
wire n_241;
wire n_504;
wire n_111;
wire n_479;
wire n_226;
wire n_125;
wire n_297;
wire n_413;
wire n_494;
wire n_539;
wire n_512;
wire n_75;
wire n_346;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_457;
wire n_119;
wire n_283;
wire n_181;
wire n_358;
wire n_534;
wire n_256;
wire n_520;
wire n_273;
wire n_253;
wire n_54;
wire n_168;
wire n_38;
wire n_442;
wire n_385;
wire n_201;
wire n_545;
wire n_484;
wire n_260;
wire n_247;
wire n_249;
wire n_349;
wire n_418;
wire n_502;
wire n_472;
wire n_292;
wire n_343;
wire n_486;
wire n_64;
wire n_291;
wire n_236;
wire n_370;
wire n_276;
wire n_374;
wire n_287;
wire n_388;
wire n_174;
wire n_400;
wire n_255;
wire n_243;
wire n_299;
wire n_352;
wire n_477;
wire n_56;
wire n_293;
wire n_275;
wire n_381;
wire n_227;
wire n_229;
wire n_454;
wire n_379;
wire n_141;
wire n_555;
wire n_65;
wire n_188;
wire n_444;
wire n_178;
wire n_360;
wire n_398;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_451;
wire n_45;
wire n_437;
wire n_268;
wire n_42;
wire n_313;
wire n_94;
wire n_547;
wire n_309;
wire n_294;
wire n_116;
wire n_416;
wire n_513;
wire n_143;
wire n_351;
wire n_467;
wire n_129;
wire n_135;
wire n_306;
wire n_540;
wire n_218;
wire n_528;
wire n_165;
wire n_406;
wire n_303;
wire n_321;
wire n_100;
wire n_368;
wire n_51;
wire n_509;
wire n_205;
wire n_519;
wire n_530;
wire n_361;
wire n_324;
wire n_86;
wire n_261;
wire n_549;
wire n_70;
wire n_435;
wire n_32;
wire n_228;
wire n_389;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_438;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_481;
wire n_191;
wire n_394;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_436;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_424;
wire n_133;
wire n_468;
wire n_257;
wire n_447;
wire n_344;
wire n_210;
wire n_206;
wire n_552;
wire n_408;
wire n_85;
wire n_96;
wire n_308;
wire n_433;
wire n_364;

NAND2xp5_ASAP7_75t_L g78 ( 
.A(n_0),
.B(n_79),
.Y(n_78)
);

OAI32xp33_ASAP7_75t_L g119 ( 
.A1(n_0),
.A2(n_39),
.A3(n_120),
.B1(n_121),
.B2(n_124),
.Y(n_119)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_0),
.Y(n_125)
);

AOI22xp33_ASAP7_75t_L g194 ( 
.A1(n_0),
.A2(n_125),
.B1(n_195),
.B2(n_201),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_L g266 ( 
.A(n_0),
.B(n_69),
.Y(n_266)
);

OAI22xp5_ASAP7_75t_SL g299 ( 
.A1(n_0),
.A2(n_92),
.B1(n_300),
.B2(n_306),
.Y(n_299)
);

OAI22xp5_ASAP7_75t_SL g70 ( 
.A1(n_1),
.A2(n_71),
.B1(n_72),
.B2(n_73),
.Y(n_70)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_1),
.Y(n_72)
);

OAI22xp5_ASAP7_75t_SL g186 ( 
.A1(n_1),
.A2(n_72),
.B1(n_126),
.B2(n_187),
.Y(n_186)
);

AOI22xp33_ASAP7_75t_SL g274 ( 
.A1(n_1),
.A2(n_72),
.B1(n_275),
.B2(n_277),
.Y(n_274)
);

AOI22xp5_ASAP7_75t_L g405 ( 
.A1(n_1),
.A2(n_72),
.B1(n_359),
.B2(n_406),
.Y(n_405)
);

AOI22xp5_ASAP7_75t_L g59 ( 
.A1(n_2),
.A2(n_60),
.B1(n_61),
.B2(n_68),
.Y(n_59)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_2),
.Y(n_68)
);

OAI22xp5_ASAP7_75t_SL g242 ( 
.A1(n_2),
.A2(n_68),
.B1(n_243),
.B2(n_244),
.Y(n_242)
);

AOI22xp5_ASAP7_75t_SL g300 ( 
.A1(n_2),
.A2(n_68),
.B1(n_301),
.B2(n_303),
.Y(n_300)
);

OAI22xp5_ASAP7_75t_L g365 ( 
.A1(n_2),
.A2(n_68),
.B1(n_366),
.B2(n_370),
.Y(n_365)
);

OAI22xp5_ASAP7_75t_SL g99 ( 
.A1(n_3),
.A2(n_100),
.B1(n_101),
.B2(n_102),
.Y(n_99)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_3),
.Y(n_101)
);

AOI22xp33_ASAP7_75t_L g382 ( 
.A1(n_3),
.A2(n_101),
.B1(n_383),
.B2(n_384),
.Y(n_382)
);

AOI22xp5_ASAP7_75t_SL g463 ( 
.A1(n_3),
.A2(n_101),
.B1(n_464),
.B2(n_469),
.Y(n_463)
);

AOI22xp5_ASAP7_75t_SL g556 ( 
.A1(n_3),
.A2(n_101),
.B1(n_370),
.B2(n_501),
.Y(n_556)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_4),
.Y(n_35)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_4),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_4),
.Y(n_52)
);

OAI22xp5_ASAP7_75t_SL g132 ( 
.A1(n_5),
.A2(n_133),
.B1(n_139),
.B2(n_140),
.Y(n_132)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_5),
.Y(n_139)
);

OAI22xp5_ASAP7_75t_L g172 ( 
.A1(n_5),
.A2(n_139),
.B1(n_173),
.B2(n_176),
.Y(n_172)
);

AOI22xp5_ASAP7_75t_L g397 ( 
.A1(n_5),
.A2(n_139),
.B1(n_398),
.B2(n_399),
.Y(n_397)
);

AOI22xp5_ASAP7_75t_L g497 ( 
.A1(n_5),
.A2(n_139),
.B1(n_498),
.B2(n_501),
.Y(n_497)
);

BUFx6f_ASAP7_75t_L g149 ( 
.A(n_6),
.Y(n_149)
);

BUFx5_ASAP7_75t_L g154 ( 
.A(n_6),
.Y(n_154)
);

BUFx6f_ASAP7_75t_L g160 ( 
.A(n_6),
.Y(n_160)
);

BUFx5_ASAP7_75t_L g231 ( 
.A(n_6),
.Y(n_231)
);

BUFx5_ASAP7_75t_L g94 ( 
.A(n_7),
.Y(n_94)
);

BUFx3_ASAP7_75t_L g109 ( 
.A(n_7),
.Y(n_109)
);

INVx2_ASAP7_75t_L g263 ( 
.A(n_7),
.Y(n_263)
);

BUFx5_ASAP7_75t_L g312 ( 
.A(n_7),
.Y(n_312)
);

OAI22xp33_ASAP7_75t_SL g110 ( 
.A1(n_8),
.A2(n_103),
.B1(n_111),
.B2(n_112),
.Y(n_110)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_8),
.Y(n_111)
);

AOI22xp33_ASAP7_75t_SL g422 ( 
.A1(n_8),
.A2(n_111),
.B1(n_423),
.B2(n_426),
.Y(n_422)
);

AOI22xp33_ASAP7_75t_SL g505 ( 
.A1(n_8),
.A2(n_62),
.B1(n_111),
.B2(n_506),
.Y(n_505)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_9),
.Y(n_49)
);

INVx3_ASAP7_75t_L g55 ( 
.A(n_9),
.Y(n_55)
);

BUFx3_ASAP7_75t_L g123 ( 
.A(n_9),
.Y(n_123)
);

BUFx6f_ASAP7_75t_L g162 ( 
.A(n_9),
.Y(n_162)
);

INVx2_ASAP7_75t_L g169 ( 
.A(n_9),
.Y(n_169)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_9),
.Y(n_190)
);

OAI22xp5_ASAP7_75t_L g164 ( 
.A1(n_10),
.A2(n_165),
.B1(n_166),
.B2(n_167),
.Y(n_164)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_10),
.Y(n_165)
);

AOI22xp5_ASAP7_75t_L g250 ( 
.A1(n_10),
.A2(n_165),
.B1(n_251),
.B2(n_254),
.Y(n_250)
);

OAI22xp5_ASAP7_75t_L g373 ( 
.A1(n_10),
.A2(n_165),
.B1(n_374),
.B2(n_375),
.Y(n_373)
);

AOI22xp5_ASAP7_75t_L g457 ( 
.A1(n_10),
.A2(n_165),
.B1(n_458),
.B2(n_459),
.Y(n_457)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_11),
.Y(n_83)
);

BUFx6f_ASAP7_75t_L g89 ( 
.A(n_11),
.Y(n_89)
);

BUFx6f_ASAP7_75t_L g353 ( 
.A(n_11),
.Y(n_353)
);

AOI22xp5_ASAP7_75t_L g431 ( 
.A1(n_12),
.A2(n_432),
.B1(n_435),
.B2(n_436),
.Y(n_431)
);

CKINVDCx20_ASAP7_75t_R g435 ( 
.A(n_12),
.Y(n_435)
);

AOI22xp33_ASAP7_75t_SL g510 ( 
.A1(n_12),
.A2(n_435),
.B1(n_511),
.B2(n_514),
.Y(n_510)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_13),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_13),
.Y(n_67)
);

AOI22xp5_ASAP7_75t_SL g330 ( 
.A1(n_14),
.A2(n_331),
.B1(n_332),
.B2(n_337),
.Y(n_330)
);

CKINVDCx20_ASAP7_75t_R g337 ( 
.A(n_14),
.Y(n_337)
);

AOI22xp33_ASAP7_75t_L g413 ( 
.A1(n_14),
.A2(n_337),
.B1(n_414),
.B2(n_416),
.Y(n_413)
);

AOI22xp5_ASAP7_75t_L g539 ( 
.A1(n_14),
.A2(n_337),
.B1(n_469),
.B2(n_540),
.Y(n_539)
);

BUFx12f_ASAP7_75t_L g98 ( 
.A(n_15),
.Y(n_98)
);

BUFx4f_ASAP7_75t_L g138 ( 
.A(n_15),
.Y(n_138)
);

INVx2_ASAP7_75t_L g143 ( 
.A(n_15),
.Y(n_143)
);

BUFx6f_ASAP7_75t_L g236 ( 
.A(n_15),
.Y(n_236)
);

AOI22xp33_ASAP7_75t_SL g444 ( 
.A1(n_16),
.A2(n_252),
.B1(n_445),
.B2(n_448),
.Y(n_444)
);

INVx1_ASAP7_75t_L g448 ( 
.A(n_16),
.Y(n_448)
);

OAI22xp5_ASAP7_75t_SL g546 ( 
.A1(n_16),
.A2(n_448),
.B1(n_547),
.B2(n_549),
.Y(n_546)
);

INVx2_ASAP7_75t_L g344 ( 
.A(n_17),
.Y(n_344)
);

BUFx5_ASAP7_75t_L g351 ( 
.A(n_17),
.Y(n_351)
);

BUFx3_ASAP7_75t_L g364 ( 
.A(n_17),
.Y(n_364)
);

BUFx8_ASAP7_75t_L g500 ( 
.A(n_17),
.Y(n_500)
);

XNOR2xp5_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_528),
.Y(n_18)
);

OAI21xp5_ASAP7_75t_SL g19 ( 
.A1(n_20),
.A2(n_486),
.B(n_526),
.Y(n_19)
);

AOI21xp5_ASAP7_75t_SL g20 ( 
.A1(n_21),
.A2(n_391),
.B(n_483),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_22),
.Y(n_21)
);

AOI21x1_ASAP7_75t_L g22 ( 
.A1(n_23),
.A2(n_324),
.B(n_390),
.Y(n_22)
);

OAI21x1_ASAP7_75t_L g23 ( 
.A1(n_24),
.A2(n_209),
.B(n_323),
.Y(n_23)
);

NOR2x1_ASAP7_75t_L g24 ( 
.A(n_25),
.B(n_182),
.Y(n_24)
);

NAND2xp5_ASAP7_75t_L g323 ( 
.A(n_25),
.B(n_182),
.Y(n_323)
);

OAI22xp5_ASAP7_75t_SL g25 ( 
.A1(n_26),
.A2(n_27),
.B1(n_116),
.B2(n_117),
.Y(n_25)
);

MAJIxp5_ASAP7_75t_L g389 ( 
.A(n_26),
.B(n_144),
.C(n_180),
.Y(n_389)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_27),
.Y(n_26)
);

XOR2x1_ASAP7_75t_L g27 ( 
.A(n_28),
.B(n_77),
.Y(n_27)
);

MAJIxp5_ASAP7_75t_L g354 ( 
.A(n_28),
.B(n_78),
.C(n_90),
.Y(n_354)
);

AOI22xp5_ASAP7_75t_SL g28 ( 
.A1(n_29),
.A2(n_58),
.B1(n_69),
.B2(n_70),
.Y(n_28)
);

AOI22xp5_ASAP7_75t_L g372 ( 
.A1(n_29),
.A2(n_69),
.B1(n_70),
.B2(n_373),
.Y(n_372)
);

AOI22xp5_ASAP7_75t_SL g536 ( 
.A1(n_29),
.A2(n_69),
.B1(n_537),
.B2(n_538),
.Y(n_536)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_30),
.Y(n_29)
);

OAI22xp5_ASAP7_75t_SL g193 ( 
.A1(n_30),
.A2(n_59),
.B1(n_194),
.B2(n_208),
.Y(n_193)
);

OAI22xp5_ASAP7_75t_L g395 ( 
.A1(n_30),
.A2(n_208),
.B1(n_396),
.B2(n_397),
.Y(n_395)
);

OAI22xp5_ASAP7_75t_L g462 ( 
.A1(n_30),
.A2(n_208),
.B1(n_397),
.B2(n_463),
.Y(n_462)
);

OAI22xp5_ASAP7_75t_L g504 ( 
.A1(n_30),
.A2(n_208),
.B1(n_463),
.B2(n_505),
.Y(n_504)
);

AO21x2_ASAP7_75t_SL g30 ( 
.A1(n_31),
.A2(n_39),
.B(n_47),
.Y(n_30)
);

NAND2xp5_ASAP7_75t_L g31 ( 
.A(n_32),
.B(n_36),
.Y(n_31)
);

INVx2_ASAP7_75t_L g32 ( 
.A(n_33),
.Y(n_32)
);

INVx3_ASAP7_75t_L g33 ( 
.A(n_34),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_35),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_35),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_36),
.Y(n_60)
);

INVx2_ASAP7_75t_L g36 ( 
.A(n_37),
.Y(n_36)
);

BUFx5_ASAP7_75t_L g37 ( 
.A(n_38),
.Y(n_37)
);

INVx2_ASAP7_75t_L g46 ( 
.A(n_38),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g200 ( 
.A(n_38),
.Y(n_200)
);

BUFx6f_ASAP7_75t_L g207 ( 
.A(n_38),
.Y(n_207)
);

BUFx6f_ASAP7_75t_L g471 ( 
.A(n_38),
.Y(n_471)
);

NAND2xp5_ASAP7_75t_L g39 ( 
.A(n_40),
.B(n_44),
.Y(n_39)
);

INVx4_ASAP7_75t_L g40 ( 
.A(n_41),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_42),
.Y(n_41)
);

INVx2_ASAP7_75t_L g42 ( 
.A(n_43),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g71 ( 
.A(n_44),
.Y(n_71)
);

INVx8_ASAP7_75t_L g44 ( 
.A(n_45),
.Y(n_44)
);

INVx4_ASAP7_75t_L g401 ( 
.A(n_45),
.Y(n_401)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_46),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g543 ( 
.A(n_46),
.Y(n_543)
);

BUFx2_ASAP7_75t_L g69 ( 
.A(n_47),
.Y(n_69)
);

OAI22xp5_ASAP7_75t_L g47 ( 
.A1(n_48),
.A2(n_50),
.B1(n_53),
.B2(n_56),
.Y(n_47)
);

INVx1_ASAP7_75t_L g383 ( 
.A(n_48),
.Y(n_383)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_49),
.Y(n_48)
);

INVx2_ASAP7_75t_L g129 ( 
.A(n_49),
.Y(n_129)
);

INVx6_ASAP7_75t_L g218 ( 
.A(n_49),
.Y(n_218)
);

INVx6_ASAP7_75t_L g50 ( 
.A(n_51),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_52),
.Y(n_51)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_54),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g179 ( 
.A(n_54),
.Y(n_179)
);

BUFx3_ASAP7_75t_L g415 ( 
.A(n_54),
.Y(n_415)
);

INVx2_ASAP7_75t_L g54 ( 
.A(n_55),
.Y(n_54)
);

INVx2_ASAP7_75t_L g157 ( 
.A(n_55),
.Y(n_157)
);

BUFx3_ASAP7_75t_L g175 ( 
.A(n_55),
.Y(n_175)
);

INVx1_ASAP7_75t_L g388 ( 
.A(n_55),
.Y(n_388)
);

BUFx3_ASAP7_75t_L g419 ( 
.A(n_55),
.Y(n_419)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_57),
.Y(n_56)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_59),
.Y(n_58)
);

INVx3_ASAP7_75t_SL g506 ( 
.A(n_60),
.Y(n_506)
);

INVx1_ASAP7_75t_SL g61 ( 
.A(n_62),
.Y(n_61)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_63),
.Y(n_62)
);

INVx2_ASAP7_75t_L g63 ( 
.A(n_64),
.Y(n_63)
);

INVx2_ASAP7_75t_L g64 ( 
.A(n_65),
.Y(n_64)
);

INVx2_ASAP7_75t_L g65 ( 
.A(n_66),
.Y(n_65)
);

INVx3_ASAP7_75t_L g66 ( 
.A(n_67),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g76 ( 
.A(n_67),
.Y(n_76)
);

BUFx6f_ASAP7_75t_L g85 ( 
.A(n_67),
.Y(n_85)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_67),
.Y(n_87)
);

INVx4_ASAP7_75t_L g468 ( 
.A(n_67),
.Y(n_468)
);

INVx2_ASAP7_75t_L g208 ( 
.A(n_69),
.Y(n_208)
);

INVx2_ASAP7_75t_L g120 ( 
.A(n_71),
.Y(n_120)
);

OAI22xp5_ASAP7_75t_L g338 ( 
.A1(n_71),
.A2(n_339),
.B1(n_345),
.B2(n_349),
.Y(n_338)
);

INVx1_ASAP7_75t_SL g73 ( 
.A(n_74),
.Y(n_73)
);

INVx6_ASAP7_75t_L g74 ( 
.A(n_75),
.Y(n_74)
);

INVx6_ASAP7_75t_L g75 ( 
.A(n_76),
.Y(n_75)
);

XOR2xp5_ASAP7_75t_SL g77 ( 
.A(n_78),
.B(n_90),
.Y(n_77)
);

AOI22xp5_ASAP7_75t_L g356 ( 
.A1(n_79),
.A2(n_357),
.B1(n_360),
.B2(n_365),
.Y(n_356)
);

AOI22xp5_ASAP7_75t_L g403 ( 
.A1(n_79),
.A2(n_360),
.B1(n_365),
.B2(n_404),
.Y(n_403)
);

INVx2_ASAP7_75t_L g461 ( 
.A(n_79),
.Y(n_461)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_80),
.Y(n_79)
);

OA21x2_ASAP7_75t_L g360 ( 
.A1(n_80),
.A2(n_350),
.B(n_361),
.Y(n_360)
);

AOI22xp5_ASAP7_75t_L g80 ( 
.A1(n_81),
.A2(n_84),
.B1(n_86),
.B2(n_88),
.Y(n_80)
);

INVx3_ASAP7_75t_L g81 ( 
.A(n_82),
.Y(n_81)
);

BUFx3_ASAP7_75t_L g82 ( 
.A(n_83),
.Y(n_82)
);

INVx2_ASAP7_75t_L g84 ( 
.A(n_85),
.Y(n_84)
);

INVx2_ASAP7_75t_SL g86 ( 
.A(n_87),
.Y(n_86)
);

INVx3_ASAP7_75t_L g88 ( 
.A(n_89),
.Y(n_88)
);

INVx2_ASAP7_75t_L g348 ( 
.A(n_89),
.Y(n_348)
);

INVx4_ASAP7_75t_L g362 ( 
.A(n_89),
.Y(n_362)
);

AOI22xp5_ASAP7_75t_L g90 ( 
.A1(n_91),
.A2(n_99),
.B1(n_104),
.B2(n_110),
.Y(n_90)
);

AOI22xp5_ASAP7_75t_L g131 ( 
.A1(n_91),
.A2(n_93),
.B1(n_99),
.B2(n_132),
.Y(n_131)
);

AOI22xp5_ASAP7_75t_L g272 ( 
.A1(n_91),
.A2(n_93),
.B1(n_273),
.B2(n_282),
.Y(n_272)
);

AOI22xp5_ASAP7_75t_L g429 ( 
.A1(n_91),
.A2(n_430),
.B1(n_440),
.B2(n_443),
.Y(n_429)
);

INVx1_ASAP7_75t_SL g91 ( 
.A(n_92),
.Y(n_91)
);

OAI22xp5_ASAP7_75t_L g249 ( 
.A1(n_92),
.A2(n_250),
.B1(n_258),
.B2(n_264),
.Y(n_249)
);

OAI22xp5_ASAP7_75t_SL g308 ( 
.A1(n_92),
.A2(n_274),
.B1(n_300),
.B2(n_309),
.Y(n_308)
);

OAI22xp5_ASAP7_75t_L g328 ( 
.A1(n_92),
.A2(n_306),
.B1(n_329),
.B2(n_330),
.Y(n_328)
);

OAI22xp5_ASAP7_75t_SL g452 ( 
.A1(n_92),
.A2(n_330),
.B1(n_431),
.B2(n_453),
.Y(n_452)
);

AOI21xp5_ASAP7_75t_L g519 ( 
.A1(n_92),
.A2(n_444),
.B(n_520),
.Y(n_519)
);

OR2x2_ASAP7_75t_L g92 ( 
.A(n_93),
.B(n_95),
.Y(n_92)
);

INVx6_ASAP7_75t_L g306 ( 
.A(n_93),
.Y(n_306)
);

BUFx12f_ASAP7_75t_L g93 ( 
.A(n_94),
.Y(n_93)
);

INVx2_ASAP7_75t_L g95 ( 
.A(n_96),
.Y(n_95)
);

HB1xp67_ASAP7_75t_L g103 ( 
.A(n_96),
.Y(n_103)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_97),
.Y(n_96)
);

INVx5_ASAP7_75t_L g97 ( 
.A(n_98),
.Y(n_97)
);

BUFx6f_ASAP7_75t_L g100 ( 
.A(n_98),
.Y(n_100)
);

INVx2_ASAP7_75t_L g115 ( 
.A(n_98),
.Y(n_115)
);

INVx4_ASAP7_75t_L g253 ( 
.A(n_98),
.Y(n_253)
);

INVx2_ASAP7_75t_L g281 ( 
.A(n_98),
.Y(n_281)
);

INVx2_ASAP7_75t_L g331 ( 
.A(n_98),
.Y(n_331)
);

INVx3_ASAP7_75t_L g434 ( 
.A(n_98),
.Y(n_434)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_103),
.Y(n_102)
);

BUFx2_ASAP7_75t_L g104 ( 
.A(n_105),
.Y(n_104)
);

INVx3_ASAP7_75t_L g105 ( 
.A(n_106),
.Y(n_105)
);

INVx5_ASAP7_75t_L g106 ( 
.A(n_107),
.Y(n_106)
);

INVx4_ASAP7_75t_L g107 ( 
.A(n_108),
.Y(n_107)
);

INVx3_ASAP7_75t_L g108 ( 
.A(n_109),
.Y(n_108)
);

BUFx3_ASAP7_75t_L g521 ( 
.A(n_109),
.Y(n_521)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_110),
.Y(n_329)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_113),
.Y(n_112)
);

HB1xp67_ASAP7_75t_L g113 ( 
.A(n_114),
.Y(n_113)
);

INVx2_ASAP7_75t_L g114 ( 
.A(n_115),
.Y(n_114)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_117),
.Y(n_116)
);

OAI22xp5_ASAP7_75t_SL g117 ( 
.A1(n_118),
.A2(n_144),
.B1(n_180),
.B2(n_181),
.Y(n_117)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_118),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_L g118 ( 
.A(n_119),
.B(n_130),
.Y(n_118)
);

AOI22xp5_ASAP7_75t_L g183 ( 
.A1(n_119),
.A2(n_130),
.B1(n_131),
.B2(n_184),
.Y(n_183)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_119),
.Y(n_184)
);

INVx3_ASAP7_75t_L g121 ( 
.A(n_122),
.Y(n_121)
);

INVx3_ASAP7_75t_L g122 ( 
.A(n_123),
.Y(n_122)
);

INVx2_ASAP7_75t_L g513 ( 
.A(n_123),
.Y(n_513)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_125),
.B(n_126),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_L g227 ( 
.A(n_125),
.B(n_228),
.Y(n_227)
);

OAI21xp33_ASAP7_75t_SL g239 ( 
.A1(n_125),
.A2(n_227),
.B(n_240),
.Y(n_239)
);

NOR2xp33_ASAP7_75t_SL g295 ( 
.A(n_125),
.B(n_296),
.Y(n_295)
);

NOR2xp33_ASAP7_75t_L g313 ( 
.A(n_125),
.B(n_170),
.Y(n_313)
);

NAND2xp5_ASAP7_75t_L g339 ( 
.A(n_125),
.B(n_340),
.Y(n_339)
);

OAI21xp33_ASAP7_75t_SL g357 ( 
.A1(n_125),
.A2(n_339),
.B(n_358),
.Y(n_357)
);

INVx4_ASAP7_75t_L g126 ( 
.A(n_127),
.Y(n_126)
);

BUFx6f_ASAP7_75t_L g127 ( 
.A(n_128),
.Y(n_127)
);

INVx5_ASAP7_75t_L g128 ( 
.A(n_129),
.Y(n_128)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_131),
.Y(n_130)
);

INVxp67_ASAP7_75t_L g264 ( 
.A(n_132),
.Y(n_264)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_134),
.Y(n_133)
);

HB1xp67_ASAP7_75t_L g134 ( 
.A(n_135),
.Y(n_134)
);

INVx2_ASAP7_75t_L g135 ( 
.A(n_136),
.Y(n_135)
);

HB1xp67_ASAP7_75t_L g276 ( 
.A(n_136),
.Y(n_276)
);

INVx2_ASAP7_75t_L g136 ( 
.A(n_137),
.Y(n_136)
);

INVx2_ASAP7_75t_L g137 ( 
.A(n_138),
.Y(n_137)
);

INVx3_ASAP7_75t_L g152 ( 
.A(n_138),
.Y(n_152)
);

INVx2_ASAP7_75t_L g257 ( 
.A(n_138),
.Y(n_257)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_141),
.Y(n_140)
);

INVx3_ASAP7_75t_L g141 ( 
.A(n_142),
.Y(n_141)
);

BUFx6f_ASAP7_75t_L g150 ( 
.A(n_142),
.Y(n_150)
);

BUFx6f_ASAP7_75t_L g142 ( 
.A(n_143),
.Y(n_142)
);

BUFx6f_ASAP7_75t_L g336 ( 
.A(n_143),
.Y(n_336)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_144),
.Y(n_181)
);

OAI22xp5_ASAP7_75t_SL g144 ( 
.A1(n_145),
.A2(n_163),
.B1(n_170),
.B2(n_171),
.Y(n_144)
);

OAI22xp5_ASAP7_75t_SL g451 ( 
.A1(n_145),
.A2(n_170),
.B1(n_382),
.B2(n_422),
.Y(n_451)
);

OAI22xp5_ASAP7_75t_SL g509 ( 
.A1(n_145),
.A2(n_170),
.B1(n_413),
.B2(n_510),
.Y(n_509)
);

INVx1_ASAP7_75t_SL g145 ( 
.A(n_146),
.Y(n_145)
);

AOI22xp5_ASAP7_75t_L g185 ( 
.A1(n_146),
.A2(n_164),
.B1(n_186),
.B2(n_191),
.Y(n_185)
);

AOI22xp5_ASAP7_75t_L g238 ( 
.A1(n_146),
.A2(n_191),
.B1(n_239),
.B2(n_242),
.Y(n_238)
);

AOI22xp5_ASAP7_75t_SL g268 ( 
.A1(n_146),
.A2(n_186),
.B1(n_191),
.B2(n_242),
.Y(n_268)
);

AOI22xp5_ASAP7_75t_L g380 ( 
.A1(n_146),
.A2(n_172),
.B1(n_191),
.B2(n_381),
.Y(n_380)
);

NAND2xp5_ASAP7_75t_SL g420 ( 
.A(n_146),
.B(n_421),
.Y(n_420)
);

AOI22xp5_ASAP7_75t_SL g544 ( 
.A1(n_146),
.A2(n_191),
.B1(n_545),
.B2(n_546),
.Y(n_544)
);

AND2x2_ASAP7_75t_SL g146 ( 
.A(n_147),
.B(n_155),
.Y(n_146)
);

BUFx3_ASAP7_75t_L g170 ( 
.A(n_147),
.Y(n_170)
);

AOI22xp5_ASAP7_75t_L g147 ( 
.A1(n_148),
.A2(n_150),
.B1(n_151),
.B2(n_153),
.Y(n_147)
);

OAI22xp33_ASAP7_75t_L g155 ( 
.A1(n_148),
.A2(n_156),
.B1(n_158),
.B2(n_161),
.Y(n_155)
);

BUFx3_ASAP7_75t_L g148 ( 
.A(n_149),
.Y(n_148)
);

INVx2_ASAP7_75t_L g220 ( 
.A(n_151),
.Y(n_220)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_152),
.Y(n_151)
);

INVx4_ASAP7_75t_L g153 ( 
.A(n_154),
.Y(n_153)
);

INVx2_ASAP7_75t_L g166 ( 
.A(n_156),
.Y(n_166)
);

INVx2_ASAP7_75t_L g548 ( 
.A(n_156),
.Y(n_548)
);

INVx5_ASAP7_75t_L g156 ( 
.A(n_157),
.Y(n_156)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_159),
.Y(n_158)
);

HB1xp67_ASAP7_75t_L g159 ( 
.A(n_160),
.Y(n_159)
);

INVx6_ASAP7_75t_L g226 ( 
.A(n_160),
.Y(n_226)
);

INVx2_ASAP7_75t_L g549 ( 
.A(n_161),
.Y(n_549)
);

BUFx12f_ASAP7_75t_L g161 ( 
.A(n_162),
.Y(n_161)
);

INVx4_ASAP7_75t_L g428 ( 
.A(n_162),
.Y(n_428)
);

INVxp67_ASAP7_75t_L g163 ( 
.A(n_164),
.Y(n_163)
);

BUFx6f_ASAP7_75t_L g167 ( 
.A(n_168),
.Y(n_167)
);

INVx6_ASAP7_75t_L g228 ( 
.A(n_168),
.Y(n_228)
);

BUFx6f_ASAP7_75t_L g168 ( 
.A(n_169),
.Y(n_168)
);

INVx2_ASAP7_75t_SL g191 ( 
.A(n_170),
.Y(n_191)
);

INVxp67_ASAP7_75t_L g171 ( 
.A(n_172),
.Y(n_171)
);

BUFx3_ASAP7_75t_L g173 ( 
.A(n_174),
.Y(n_173)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_175),
.Y(n_174)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_175),
.Y(n_241)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_175),
.Y(n_243)
);

INVx2_ASAP7_75t_L g176 ( 
.A(n_177),
.Y(n_176)
);

INVx3_ASAP7_75t_L g177 ( 
.A(n_178),
.Y(n_177)
);

INVx2_ASAP7_75t_L g178 ( 
.A(n_179),
.Y(n_178)
);

MAJIxp5_ASAP7_75t_L g182 ( 
.A(n_183),
.B(n_185),
.C(n_192),
.Y(n_182)
);

XOR2xp5_ASAP7_75t_L g319 ( 
.A(n_183),
.B(n_320),
.Y(n_319)
);

OAI22xp5_ASAP7_75t_SL g320 ( 
.A1(n_185),
.A2(n_192),
.B1(n_193),
.B2(n_321),
.Y(n_320)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_185),
.Y(n_321)
);

INVx3_ASAP7_75t_L g187 ( 
.A(n_188),
.Y(n_187)
);

INVx2_ASAP7_75t_L g188 ( 
.A(n_189),
.Y(n_188)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_190),
.Y(n_189)
);

INVx2_ASAP7_75t_L g517 ( 
.A(n_190),
.Y(n_517)
);

NAND2xp5_ASAP7_75t_SL g411 ( 
.A(n_191),
.B(n_412),
.Y(n_411)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_193),
.Y(n_192)
);

NOR2xp33_ASAP7_75t_L g345 ( 
.A(n_195),
.B(n_346),
.Y(n_345)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_196),
.Y(n_195)
);

INVx2_ASAP7_75t_L g196 ( 
.A(n_197),
.Y(n_196)
);

INVx1_ASAP7_75t_L g374 ( 
.A(n_197),
.Y(n_374)
);

INVx3_ASAP7_75t_L g197 ( 
.A(n_198),
.Y(n_197)
);

INVx2_ASAP7_75t_L g198 ( 
.A(n_199),
.Y(n_198)
);

INVx2_ASAP7_75t_L g199 ( 
.A(n_200),
.Y(n_199)
);

INVx1_ASAP7_75t_SL g201 ( 
.A(n_202),
.Y(n_201)
);

INVx2_ASAP7_75t_L g202 ( 
.A(n_203),
.Y(n_202)
);

BUFx6f_ASAP7_75t_L g203 ( 
.A(n_204),
.Y(n_203)
);

INVx2_ASAP7_75t_L g204 ( 
.A(n_205),
.Y(n_204)
);

INVx2_ASAP7_75t_L g205 ( 
.A(n_206),
.Y(n_205)
);

BUFx6f_ASAP7_75t_L g206 ( 
.A(n_207),
.Y(n_206)
);

INVx3_ASAP7_75t_L g379 ( 
.A(n_207),
.Y(n_379)
);

AOI21xp5_ASAP7_75t_L g209 ( 
.A1(n_210),
.A2(n_317),
.B(n_322),
.Y(n_209)
);

OAI21x1_ASAP7_75t_L g210 ( 
.A1(n_211),
.A2(n_270),
.B(n_316),
.Y(n_210)
);

AND2x2_ASAP7_75t_L g211 ( 
.A(n_212),
.B(n_248),
.Y(n_211)
);

OR2x2_ASAP7_75t_L g316 ( 
.A(n_212),
.B(n_248),
.Y(n_316)
);

NAND2xp5_ASAP7_75t_L g212 ( 
.A(n_213),
.B(n_237),
.Y(n_212)
);

HB1xp67_ASAP7_75t_L g213 ( 
.A(n_214),
.Y(n_213)
);

AOI22xp5_ASAP7_75t_L g283 ( 
.A1(n_214),
.A2(n_237),
.B1(n_238),
.B2(n_284),
.Y(n_283)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_214),
.Y(n_284)
);

OAI32xp33_ASAP7_75t_L g214 ( 
.A1(n_215),
.A2(n_219),
.A3(n_221),
.B1(n_227),
.B2(n_229),
.Y(n_214)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_216),
.Y(n_215)
);

HB1xp67_ASAP7_75t_L g216 ( 
.A(n_217),
.Y(n_216)
);

INVx2_ASAP7_75t_L g425 ( 
.A(n_217),
.Y(n_425)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_218),
.Y(n_217)
);

INVx2_ASAP7_75t_L g247 ( 
.A(n_218),
.Y(n_247)
);

INVx2_ASAP7_75t_L g219 ( 
.A(n_220),
.Y(n_219)
);

HB1xp67_ASAP7_75t_L g221 ( 
.A(n_222),
.Y(n_221)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_223),
.Y(n_222)
);

HB1xp67_ASAP7_75t_L g223 ( 
.A(n_224),
.Y(n_223)
);

INVx4_ASAP7_75t_L g224 ( 
.A(n_225),
.Y(n_224)
);

INVx3_ASAP7_75t_L g225 ( 
.A(n_226),
.Y(n_225)
);

NOR2xp33_ASAP7_75t_L g229 ( 
.A(n_230),
.B(n_232),
.Y(n_229)
);

INVx2_ASAP7_75t_SL g230 ( 
.A(n_231),
.Y(n_230)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_233),
.Y(n_232)
);

BUFx2_ASAP7_75t_L g233 ( 
.A(n_234),
.Y(n_233)
);

INVx5_ASAP7_75t_L g234 ( 
.A(n_235),
.Y(n_234)
);

INVx2_ASAP7_75t_L g235 ( 
.A(n_236),
.Y(n_235)
);

INVx3_ASAP7_75t_L g294 ( 
.A(n_236),
.Y(n_294)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_238),
.Y(n_237)
);

BUFx2_ASAP7_75t_L g240 ( 
.A(n_241),
.Y(n_240)
);

INVx3_ASAP7_75t_L g244 ( 
.A(n_245),
.Y(n_244)
);

INVx3_ASAP7_75t_L g245 ( 
.A(n_246),
.Y(n_245)
);

INVx2_ASAP7_75t_L g246 ( 
.A(n_247),
.Y(n_246)
);

XNOR2xp5_ASAP7_75t_L g248 ( 
.A(n_249),
.B(n_265),
.Y(n_248)
);

MAJIxp5_ASAP7_75t_L g318 ( 
.A(n_249),
.B(n_267),
.C(n_269),
.Y(n_318)
);

INVxp67_ASAP7_75t_L g282 ( 
.A(n_250),
.Y(n_282)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_252),
.Y(n_251)
);

INVx2_ASAP7_75t_L g252 ( 
.A(n_253),
.Y(n_252)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_255),
.Y(n_254)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_256),
.Y(n_255)
);

INVx2_ASAP7_75t_L g256 ( 
.A(n_257),
.Y(n_256)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_259),
.Y(n_258)
);

BUFx3_ASAP7_75t_L g259 ( 
.A(n_260),
.Y(n_259)
);

BUFx6f_ASAP7_75t_L g260 ( 
.A(n_261),
.Y(n_260)
);

INVx2_ASAP7_75t_L g453 ( 
.A(n_261),
.Y(n_453)
);

BUFx6f_ASAP7_75t_L g261 ( 
.A(n_262),
.Y(n_261)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_262),
.Y(n_298)
);

INVx2_ASAP7_75t_L g262 ( 
.A(n_263),
.Y(n_262)
);

INVx3_ASAP7_75t_L g442 ( 
.A(n_263),
.Y(n_442)
);

OAI22xp5_ASAP7_75t_L g265 ( 
.A1(n_266),
.A2(n_267),
.B1(n_268),
.B2(n_269),
.Y(n_265)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_266),
.Y(n_269)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_268),
.Y(n_267)
);

AOI21x1_ASAP7_75t_SL g270 ( 
.A1(n_271),
.A2(n_285),
.B(n_315),
.Y(n_270)
);

NAND2xp5_ASAP7_75t_L g271 ( 
.A(n_272),
.B(n_283),
.Y(n_271)
);

NOR2xp33_ASAP7_75t_L g315 ( 
.A(n_272),
.B(n_283),
.Y(n_315)
);

INVxp67_ASAP7_75t_L g273 ( 
.A(n_274),
.Y(n_273)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_276),
.Y(n_275)
);

BUFx3_ASAP7_75t_L g277 ( 
.A(n_278),
.Y(n_277)
);

INVx2_ASAP7_75t_L g278 ( 
.A(n_279),
.Y(n_278)
);

INVx2_ASAP7_75t_L g279 ( 
.A(n_280),
.Y(n_279)
);

INVx2_ASAP7_75t_L g280 ( 
.A(n_281),
.Y(n_280)
);

OAI21xp5_ASAP7_75t_L g285 ( 
.A1(n_286),
.A2(n_307),
.B(n_314),
.Y(n_285)
);

NAND2xp5_ASAP7_75t_L g286 ( 
.A(n_287),
.B(n_299),
.Y(n_286)
);

NOR2xp33_ASAP7_75t_L g287 ( 
.A(n_288),
.B(n_295),
.Y(n_287)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_289),
.Y(n_288)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_290),
.Y(n_289)
);

HB1xp67_ASAP7_75t_L g290 ( 
.A(n_291),
.Y(n_290)
);

INVx2_ASAP7_75t_L g291 ( 
.A(n_292),
.Y(n_291)
);

BUFx2_ASAP7_75t_L g302 ( 
.A(n_292),
.Y(n_302)
);

BUFx6f_ASAP7_75t_L g292 ( 
.A(n_293),
.Y(n_292)
);

INVx2_ASAP7_75t_L g293 ( 
.A(n_294),
.Y(n_293)
);

INVx2_ASAP7_75t_L g305 ( 
.A(n_294),
.Y(n_305)
);

INVx2_ASAP7_75t_L g439 ( 
.A(n_294),
.Y(n_439)
);

INVx2_ASAP7_75t_L g296 ( 
.A(n_297),
.Y(n_296)
);

INVx2_ASAP7_75t_L g297 ( 
.A(n_298),
.Y(n_297)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_302),
.Y(n_301)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_304),
.Y(n_303)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_305),
.Y(n_304)
);

NOR2xp33_ASAP7_75t_L g307 ( 
.A(n_308),
.B(n_313),
.Y(n_307)
);

NAND2xp5_ASAP7_75t_L g314 ( 
.A(n_308),
.B(n_313),
.Y(n_314)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_310),
.Y(n_309)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_311),
.Y(n_310)
);

INVx3_ASAP7_75t_L g311 ( 
.A(n_312),
.Y(n_311)
);

NAND2xp5_ASAP7_75t_L g317 ( 
.A(n_318),
.B(n_319),
.Y(n_317)
);

NOR2xp33_ASAP7_75t_L g322 ( 
.A(n_318),
.B(n_319),
.Y(n_322)
);

NAND2xp5_ASAP7_75t_SL g324 ( 
.A(n_325),
.B(n_389),
.Y(n_324)
);

NOR2xp33_ASAP7_75t_L g390 ( 
.A(n_325),
.B(n_389),
.Y(n_390)
);

XOR2xp5_ASAP7_75t_L g325 ( 
.A(n_326),
.B(n_355),
.Y(n_325)
);

XNOR2xp5_ASAP7_75t_L g326 ( 
.A(n_327),
.B(n_354),
.Y(n_326)
);

MAJIxp5_ASAP7_75t_L g479 ( 
.A(n_327),
.B(n_354),
.C(n_355),
.Y(n_479)
);

XOR2xp5_ASAP7_75t_L g327 ( 
.A(n_328),
.B(n_338),
.Y(n_327)
);

NAND2xp5_ASAP7_75t_L g402 ( 
.A(n_328),
.B(n_338),
.Y(n_402)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_333),
.Y(n_332)
);

HB1xp67_ASAP7_75t_L g333 ( 
.A(n_334),
.Y(n_333)
);

INVx3_ASAP7_75t_L g334 ( 
.A(n_335),
.Y(n_334)
);

INVx2_ASAP7_75t_L g335 ( 
.A(n_336),
.Y(n_335)
);

BUFx6f_ASAP7_75t_L g447 ( 
.A(n_336),
.Y(n_447)
);

INVx4_ASAP7_75t_L g340 ( 
.A(n_341),
.Y(n_340)
);

INVx6_ASAP7_75t_L g341 ( 
.A(n_342),
.Y(n_341)
);

INVx4_ASAP7_75t_L g359 ( 
.A(n_342),
.Y(n_359)
);

INVx5_ASAP7_75t_L g342 ( 
.A(n_343),
.Y(n_342)
);

INVx8_ASAP7_75t_L g460 ( 
.A(n_343),
.Y(n_460)
);

BUFx6f_ASAP7_75t_L g343 ( 
.A(n_344),
.Y(n_343)
);

BUFx6f_ASAP7_75t_L g369 ( 
.A(n_344),
.Y(n_369)
);

INVx1_ASAP7_75t_L g346 ( 
.A(n_347),
.Y(n_346)
);

INVx1_ASAP7_75t_L g347 ( 
.A(n_348),
.Y(n_347)
);

INVxp67_ASAP7_75t_L g349 ( 
.A(n_350),
.Y(n_349)
);

AND2x2_ASAP7_75t_L g350 ( 
.A(n_351),
.B(n_352),
.Y(n_350)
);

INVx2_ASAP7_75t_L g352 ( 
.A(n_353),
.Y(n_352)
);

XOR2xp5_ASAP7_75t_L g355 ( 
.A(n_356),
.B(n_371),
.Y(n_355)
);

MAJIxp5_ASAP7_75t_L g477 ( 
.A(n_356),
.B(n_372),
.C(n_380),
.Y(n_477)
);

INVx1_ASAP7_75t_L g358 ( 
.A(n_359),
.Y(n_358)
);

INVx3_ASAP7_75t_SL g456 ( 
.A(n_360),
.Y(n_456)
);

NOR2xp33_ASAP7_75t_L g361 ( 
.A(n_362),
.B(n_363),
.Y(n_361)
);

INVx5_ASAP7_75t_L g370 ( 
.A(n_363),
.Y(n_370)
);

BUFx6f_ASAP7_75t_L g363 ( 
.A(n_364),
.Y(n_363)
);

BUFx6f_ASAP7_75t_L g407 ( 
.A(n_364),
.Y(n_407)
);

BUFx12f_ASAP7_75t_L g503 ( 
.A(n_364),
.Y(n_503)
);

INVx2_ASAP7_75t_L g366 ( 
.A(n_367),
.Y(n_366)
);

INVx3_ASAP7_75t_L g367 ( 
.A(n_368),
.Y(n_367)
);

INVx6_ASAP7_75t_L g368 ( 
.A(n_369),
.Y(n_368)
);

XNOR2xp5_ASAP7_75t_L g371 ( 
.A(n_372),
.B(n_380),
.Y(n_371)
);

INVx1_ASAP7_75t_L g396 ( 
.A(n_373),
.Y(n_396)
);

INVx2_ASAP7_75t_L g375 ( 
.A(n_376),
.Y(n_375)
);

INVx2_ASAP7_75t_L g398 ( 
.A(n_376),
.Y(n_398)
);

INVx4_ASAP7_75t_L g376 ( 
.A(n_377),
.Y(n_376)
);

INVx2_ASAP7_75t_L g377 ( 
.A(n_378),
.Y(n_377)
);

INVx1_ASAP7_75t_L g378 ( 
.A(n_379),
.Y(n_378)
);

INVx1_ASAP7_75t_L g381 ( 
.A(n_382),
.Y(n_381)
);

INVx2_ASAP7_75t_L g384 ( 
.A(n_385),
.Y(n_384)
);

INVx2_ASAP7_75t_L g385 ( 
.A(n_386),
.Y(n_385)
);

INVx2_ASAP7_75t_L g386 ( 
.A(n_387),
.Y(n_386)
);

INVx2_ASAP7_75t_L g387 ( 
.A(n_388),
.Y(n_387)
);

AOI21x1_ASAP7_75t_L g391 ( 
.A1(n_392),
.A2(n_472),
.B(n_478),
.Y(n_391)
);

MAJIxp5_ASAP7_75t_L g484 ( 
.A(n_392),
.B(n_472),
.C(n_485),
.Y(n_484)
);

XNOR2x1_ASAP7_75t_L g392 ( 
.A(n_393),
.B(n_408),
.Y(n_392)
);

MAJIxp5_ASAP7_75t_L g525 ( 
.A(n_393),
.B(n_409),
.C(n_449),
.Y(n_525)
);

MAJIxp5_ASAP7_75t_L g393 ( 
.A(n_394),
.B(n_402),
.C(n_403),
.Y(n_393)
);

INVxp67_ASAP7_75t_L g394 ( 
.A(n_395),
.Y(n_394)
);

XNOR2xp5_ASAP7_75t_L g475 ( 
.A(n_395),
.B(n_403),
.Y(n_475)
);

INVx3_ASAP7_75t_L g399 ( 
.A(n_400),
.Y(n_399)
);

INVx2_ASAP7_75t_L g400 ( 
.A(n_401),
.Y(n_400)
);

XOR2x1_ASAP7_75t_SL g474 ( 
.A(n_402),
.B(n_475),
.Y(n_474)
);

INVx1_ASAP7_75t_L g404 ( 
.A(n_405),
.Y(n_404)
);

OAI22xp5_ASAP7_75t_L g455 ( 
.A1(n_405),
.A2(n_456),
.B1(n_457),
.B2(n_461),
.Y(n_455)
);

BUFx3_ASAP7_75t_L g406 ( 
.A(n_407),
.Y(n_406)
);

XOR2xp5_ASAP7_75t_L g408 ( 
.A(n_409),
.B(n_449),
.Y(n_408)
);

XNOR2xp5_ASAP7_75t_L g409 ( 
.A(n_410),
.B(n_429),
.Y(n_409)
);

NAND2xp5_ASAP7_75t_L g410 ( 
.A(n_411),
.B(n_420),
.Y(n_410)
);

AOI21xp5_ASAP7_75t_L g507 ( 
.A1(n_411),
.A2(n_420),
.B(n_429),
.Y(n_507)
);

INVx1_ASAP7_75t_L g412 ( 
.A(n_413),
.Y(n_412)
);

INVx1_ASAP7_75t_L g414 ( 
.A(n_415),
.Y(n_414)
);

INVx2_ASAP7_75t_L g416 ( 
.A(n_417),
.Y(n_416)
);

INVx2_ASAP7_75t_L g417 ( 
.A(n_418),
.Y(n_417)
);

INVx3_ASAP7_75t_L g418 ( 
.A(n_419),
.Y(n_418)
);

INVxp67_ASAP7_75t_L g421 ( 
.A(n_422),
.Y(n_421)
);

INVx2_ASAP7_75t_L g423 ( 
.A(n_424),
.Y(n_423)
);

INVx2_ASAP7_75t_L g424 ( 
.A(n_425),
.Y(n_424)
);

INVx1_ASAP7_75t_L g426 ( 
.A(n_427),
.Y(n_426)
);

HB1xp67_ASAP7_75t_L g427 ( 
.A(n_428),
.Y(n_427)
);

INVx1_ASAP7_75t_L g430 ( 
.A(n_431),
.Y(n_430)
);

INVx2_ASAP7_75t_L g432 ( 
.A(n_433),
.Y(n_432)
);

INVx4_ASAP7_75t_L g433 ( 
.A(n_434),
.Y(n_433)
);

BUFx6f_ASAP7_75t_L g436 ( 
.A(n_437),
.Y(n_436)
);

INVx3_ASAP7_75t_L g437 ( 
.A(n_438),
.Y(n_437)
);

INVx2_ASAP7_75t_L g438 ( 
.A(n_439),
.Y(n_438)
);

INVx6_ASAP7_75t_L g440 ( 
.A(n_441),
.Y(n_440)
);

INVx6_ASAP7_75t_L g441 ( 
.A(n_442),
.Y(n_441)
);

INVxp67_ASAP7_75t_L g443 ( 
.A(n_444),
.Y(n_443)
);

INVx1_ASAP7_75t_SL g445 ( 
.A(n_446),
.Y(n_445)
);

INVx3_ASAP7_75t_L g446 ( 
.A(n_447),
.Y(n_446)
);

XNOR2xp5_ASAP7_75t_L g449 ( 
.A(n_450),
.B(n_454),
.Y(n_449)
);

INVxp67_ASAP7_75t_L g490 ( 
.A(n_450),
.Y(n_490)
);

NAND2xp5_ASAP7_75t_SL g450 ( 
.A(n_451),
.B(n_452),
.Y(n_450)
);

XOR2x2_ASAP7_75t_SL g476 ( 
.A(n_451),
.B(n_452),
.Y(n_476)
);

XOR2xp5_ASAP7_75t_L g454 ( 
.A(n_455),
.B(n_462),
.Y(n_454)
);

HB1xp67_ASAP7_75t_L g491 ( 
.A(n_455),
.Y(n_491)
);

OAI22xp5_ASAP7_75t_L g496 ( 
.A1(n_456),
.A2(n_457),
.B1(n_461),
.B2(n_497),
.Y(n_496)
);

OAI22xp5_ASAP7_75t_SL g555 ( 
.A1(n_456),
.A2(n_461),
.B1(n_497),
.B2(n_556),
.Y(n_555)
);

INVx2_ASAP7_75t_L g458 ( 
.A(n_459),
.Y(n_458)
);

BUFx2_ASAP7_75t_L g459 ( 
.A(n_460),
.Y(n_459)
);

HB1xp67_ASAP7_75t_L g492 ( 
.A(n_462),
.Y(n_492)
);

INVx1_ASAP7_75t_L g464 ( 
.A(n_465),
.Y(n_464)
);

HB1xp67_ASAP7_75t_L g465 ( 
.A(n_466),
.Y(n_465)
);

HB1xp67_ASAP7_75t_L g466 ( 
.A(n_467),
.Y(n_466)
);

INVx6_ASAP7_75t_L g467 ( 
.A(n_468),
.Y(n_467)
);

INVx2_ASAP7_75t_L g469 ( 
.A(n_470),
.Y(n_469)
);

INVx2_ASAP7_75t_L g470 ( 
.A(n_471),
.Y(n_470)
);

MAJIxp5_ASAP7_75t_L g472 ( 
.A(n_473),
.B(n_476),
.C(n_477),
.Y(n_472)
);

AOI22xp5_ASAP7_75t_L g480 ( 
.A1(n_473),
.A2(n_474),
.B1(n_481),
.B2(n_482),
.Y(n_480)
);

INVx1_ASAP7_75t_L g473 ( 
.A(n_474),
.Y(n_473)
);

XNOR2xp5_ASAP7_75t_L g481 ( 
.A(n_476),
.B(n_477),
.Y(n_481)
);

AND2x2_ASAP7_75t_L g478 ( 
.A(n_479),
.B(n_480),
.Y(n_478)
);

OR2x2_ASAP7_75t_L g485 ( 
.A(n_479),
.B(n_480),
.Y(n_485)
);

INVx1_ASAP7_75t_L g482 ( 
.A(n_481),
.Y(n_482)
);

HB1xp67_ASAP7_75t_L g483 ( 
.A(n_484),
.Y(n_483)
);

INVxp67_ASAP7_75t_L g486 ( 
.A(n_487),
.Y(n_486)
);

NAND2xp5_ASAP7_75t_L g487 ( 
.A(n_488),
.B(n_525),
.Y(n_487)
);

NOR2xp33_ASAP7_75t_L g527 ( 
.A(n_488),
.B(n_525),
.Y(n_527)
);

XNOR2xp5_ASAP7_75t_L g488 ( 
.A(n_489),
.B(n_493),
.Y(n_488)
);

INVx1_ASAP7_75t_L g531 ( 
.A(n_489),
.Y(n_531)
);

MAJIxp5_ASAP7_75t_L g489 ( 
.A(n_490),
.B(n_491),
.C(n_492),
.Y(n_489)
);

AOI22xp5_ASAP7_75t_L g493 ( 
.A1(n_494),
.A2(n_508),
.B1(n_523),
.B2(n_524),
.Y(n_493)
);

INVx1_ASAP7_75t_L g524 ( 
.A(n_494),
.Y(n_524)
);

XNOR2xp5_ASAP7_75t_L g494 ( 
.A(n_495),
.B(n_507),
.Y(n_494)
);

XOR2xp5_ASAP7_75t_L g495 ( 
.A(n_496),
.B(n_504),
.Y(n_495)
);

MAJIxp5_ASAP7_75t_R g533 ( 
.A(n_496),
.B(n_504),
.C(n_507),
.Y(n_533)
);

BUFx2_ASAP7_75t_L g498 ( 
.A(n_499),
.Y(n_498)
);

INVx2_ASAP7_75t_L g499 ( 
.A(n_500),
.Y(n_499)
);

INVx2_ASAP7_75t_L g501 ( 
.A(n_502),
.Y(n_501)
);

INVx5_ASAP7_75t_L g502 ( 
.A(n_503),
.Y(n_502)
);

INVxp67_ASAP7_75t_L g537 ( 
.A(n_505),
.Y(n_537)
);

INVx1_ASAP7_75t_L g523 ( 
.A(n_508),
.Y(n_523)
);

MAJIxp5_ASAP7_75t_L g530 ( 
.A(n_508),
.B(n_524),
.C(n_531),
.Y(n_530)
);

OAI22xp5_ASAP7_75t_SL g508 ( 
.A1(n_509),
.A2(n_518),
.B1(n_519),
.B2(n_522),
.Y(n_508)
);

INVxp67_ASAP7_75t_L g522 ( 
.A(n_509),
.Y(n_522)
);

NAND2xp5_ASAP7_75t_L g557 ( 
.A(n_509),
.B(n_519),
.Y(n_557)
);

INVxp67_ASAP7_75t_L g545 ( 
.A(n_510),
.Y(n_545)
);

INVx1_ASAP7_75t_L g511 ( 
.A(n_512),
.Y(n_511)
);

INVx1_ASAP7_75t_L g512 ( 
.A(n_513),
.Y(n_512)
);

BUFx3_ASAP7_75t_L g514 ( 
.A(n_515),
.Y(n_514)
);

INVx3_ASAP7_75t_L g515 ( 
.A(n_516),
.Y(n_515)
);

INVx1_ASAP7_75t_L g516 ( 
.A(n_517),
.Y(n_516)
);

AOI22xp5_ASAP7_75t_L g553 ( 
.A1(n_518),
.A2(n_519),
.B1(n_554),
.B2(n_555),
.Y(n_553)
);

INVx1_ASAP7_75t_L g518 ( 
.A(n_519),
.Y(n_518)
);

INVx1_ASAP7_75t_L g520 ( 
.A(n_521),
.Y(n_520)
);

INVxp33_ASAP7_75t_L g526 ( 
.A(n_527),
.Y(n_526)
);

NOR2xp33_ASAP7_75t_L g528 ( 
.A(n_529),
.B(n_559),
.Y(n_528)
);

NOR2xp33_ASAP7_75t_L g529 ( 
.A(n_530),
.B(n_532),
.Y(n_529)
);

NAND2xp5_ASAP7_75t_SL g560 ( 
.A(n_530),
.B(n_532),
.Y(n_560)
);

XNOR2xp5_ASAP7_75t_L g532 ( 
.A(n_533),
.B(n_534),
.Y(n_532)
);

XNOR2xp5_ASAP7_75t_L g534 ( 
.A(n_535),
.B(n_551),
.Y(n_534)
);

OAI21xp5_ASAP7_75t_SL g535 ( 
.A1(n_536),
.A2(n_544),
.B(n_550),
.Y(n_535)
);

NAND2xp5_ASAP7_75t_L g550 ( 
.A(n_536),
.B(n_544),
.Y(n_550)
);

INVxp67_ASAP7_75t_L g538 ( 
.A(n_539),
.Y(n_538)
);

INVx4_ASAP7_75t_L g540 ( 
.A(n_541),
.Y(n_540)
);

INVx2_ASAP7_75t_L g541 ( 
.A(n_542),
.Y(n_541)
);

BUFx6f_ASAP7_75t_L g542 ( 
.A(n_543),
.Y(n_542)
);

BUFx2_ASAP7_75t_L g547 ( 
.A(n_548),
.Y(n_547)
);

OAI22xp5_ASAP7_75t_SL g551 ( 
.A1(n_552),
.A2(n_553),
.B1(n_557),
.B2(n_558),
.Y(n_551)
);

INVx1_ASAP7_75t_L g552 ( 
.A(n_553),
.Y(n_552)
);

INVx1_ASAP7_75t_L g554 ( 
.A(n_555),
.Y(n_554)
);

INVx1_ASAP7_75t_L g558 ( 
.A(n_557),
.Y(n_558)
);

INVxp33_ASAP7_75t_L g559 ( 
.A(n_560),
.Y(n_559)
);


endmodule