module real_aes_15977_n_344 (n_76, n_113, n_187, n_90, n_257, n_65, n_74, n_185, n_285, n_30, n_222, n_61, n_20, n_287, n_64, n_254, n_207, n_10, n_83, n_181, n_124, n_191, n_209, n_299, n_322, n_328, n_19, n_40, n_318, n_239, n_100, n_54, n_112, n_319, n_35, n_42, n_329, n_132, n_131, n_144, n_169, n_242, n_308, n_172, n_341, n_232, n_6, n_69, n_317, n_321, n_73, n_320, n_77, n_260, n_37, n_97, n_186, n_138, n_26, n_235, n_245, n_161, n_189, n_271, n_2, n_145, n_227, n_92, n_330, n_332, n_292, n_116, n_94, n_289, n_280, n_333, n_213, n_184, n_28, n_202, n_56, n_34, n_98, n_121, n_125, n_216, n_82, n_327, n_47, n_106, n_32, n_263, n_230, n_51, n_248, n_301, n_27, n_343, n_174, n_18, n_104, n_211, n_281, n_173, n_234, n_284, n_153, n_316, n_75, n_178, n_298, n_49, n_43, n_297, n_9, n_119, n_310, n_164, n_231, n_44, n_102, n_122, n_141, n_128, n_111, n_167, n_80, n_179, n_12, n_68, n_129, n_304, n_311, n_324, n_25, n_278, n_236, n_267, n_218, n_48, n_204, n_339, n_89, n_277, n_331, n_93, n_182, n_323, n_199, n_142, n_223, n_67, n_250, n_85, n_45, n_5, n_244, n_118, n_139, n_87, n_171, n_78, n_146, n_17, n_226, n_255, n_286, n_120, n_261, n_238, n_58, n_165, n_246, n_176, n_163, n_29, n_52, n_251, n_220, n_197, n_296, n_3, n_41, n_256, n_71, n_302, n_126, n_200, n_115, n_96, n_110, n_150, n_147, n_288, n_23, n_334, n_274, n_160, n_303, n_95, n_188, n_269, n_201, n_306, n_158, n_4, n_193, n_293, n_162, n_275, n_214, n_46, n_109, n_59, n_203, n_81, n_133, n_273, n_114, n_276, n_295, n_265, n_154, n_127, n_326, n_24, n_217, n_55, n_62, n_291, n_148, n_88, n_159, n_11, n_108, n_60, n_233, n_290, n_155, n_243, n_268, n_136, n_157, n_282, n_101, n_309, n_229, n_107, n_33, n_53, n_36, n_149, n_190, n_262, n_134, n_336, n_195, n_300, n_252, n_283, n_314, n_249, n_221, n_156, n_57, n_66, n_21, n_31, n_8, n_312, n_183, n_266, n_205, n_335, n_177, n_313, n_22, n_140, n_219, n_180, n_212, n_210, n_325, n_338, n_103, n_166, n_224, n_151, n_130, n_253, n_99, n_15, n_72, n_152, n_198, n_7, n_228, n_272, n_196, n_315, n_123, n_279, n_79, n_270, n_305, n_117, n_208, n_215, n_135, n_70, n_50, n_170, n_86, n_340, n_13, n_168, n_175, n_241, n_105, n_84, n_294, n_258, n_206, n_307, n_342, n_14, n_194, n_137, n_225, n_16, n_39, n_337, n_247, n_240, n_38, n_259, n_143, n_192, n_0, n_264, n_63, n_1, n_237, n_91, n_344);
input n_76;
input n_113;
input n_187;
input n_90;
input n_257;
input n_65;
input n_74;
input n_185;
input n_285;
input n_30;
input n_222;
input n_61;
input n_20;
input n_287;
input n_64;
input n_254;
input n_207;
input n_10;
input n_83;
input n_181;
input n_124;
input n_191;
input n_209;
input n_299;
input n_322;
input n_328;
input n_19;
input n_40;
input n_318;
input n_239;
input n_100;
input n_54;
input n_112;
input n_319;
input n_35;
input n_42;
input n_329;
input n_132;
input n_131;
input n_144;
input n_169;
input n_242;
input n_308;
input n_172;
input n_341;
input n_232;
input n_6;
input n_69;
input n_317;
input n_321;
input n_73;
input n_320;
input n_77;
input n_260;
input n_37;
input n_97;
input n_186;
input n_138;
input n_26;
input n_235;
input n_245;
input n_161;
input n_189;
input n_271;
input n_2;
input n_145;
input n_227;
input n_92;
input n_330;
input n_332;
input n_292;
input n_116;
input n_94;
input n_289;
input n_280;
input n_333;
input n_213;
input n_184;
input n_28;
input n_202;
input n_56;
input n_34;
input n_98;
input n_121;
input n_125;
input n_216;
input n_82;
input n_327;
input n_47;
input n_106;
input n_32;
input n_263;
input n_230;
input n_51;
input n_248;
input n_301;
input n_27;
input n_343;
input n_174;
input n_18;
input n_104;
input n_211;
input n_281;
input n_173;
input n_234;
input n_284;
input n_153;
input n_316;
input n_75;
input n_178;
input n_298;
input n_49;
input n_43;
input n_297;
input n_9;
input n_119;
input n_310;
input n_164;
input n_231;
input n_44;
input n_102;
input n_122;
input n_141;
input n_128;
input n_111;
input n_167;
input n_80;
input n_179;
input n_12;
input n_68;
input n_129;
input n_304;
input n_311;
input n_324;
input n_25;
input n_278;
input n_236;
input n_267;
input n_218;
input n_48;
input n_204;
input n_339;
input n_89;
input n_277;
input n_331;
input n_93;
input n_182;
input n_323;
input n_199;
input n_142;
input n_223;
input n_67;
input n_250;
input n_85;
input n_45;
input n_5;
input n_244;
input n_118;
input n_139;
input n_87;
input n_171;
input n_78;
input n_146;
input n_17;
input n_226;
input n_255;
input n_286;
input n_120;
input n_261;
input n_238;
input n_58;
input n_165;
input n_246;
input n_176;
input n_163;
input n_29;
input n_52;
input n_251;
input n_220;
input n_197;
input n_296;
input n_3;
input n_41;
input n_256;
input n_71;
input n_302;
input n_126;
input n_200;
input n_115;
input n_96;
input n_110;
input n_150;
input n_147;
input n_288;
input n_23;
input n_334;
input n_274;
input n_160;
input n_303;
input n_95;
input n_188;
input n_269;
input n_201;
input n_306;
input n_158;
input n_4;
input n_193;
input n_293;
input n_162;
input n_275;
input n_214;
input n_46;
input n_109;
input n_59;
input n_203;
input n_81;
input n_133;
input n_273;
input n_114;
input n_276;
input n_295;
input n_265;
input n_154;
input n_127;
input n_326;
input n_24;
input n_217;
input n_55;
input n_62;
input n_291;
input n_148;
input n_88;
input n_159;
input n_11;
input n_108;
input n_60;
input n_233;
input n_290;
input n_155;
input n_243;
input n_268;
input n_136;
input n_157;
input n_282;
input n_101;
input n_309;
input n_229;
input n_107;
input n_33;
input n_53;
input n_36;
input n_149;
input n_190;
input n_262;
input n_134;
input n_336;
input n_195;
input n_300;
input n_252;
input n_283;
input n_314;
input n_249;
input n_221;
input n_156;
input n_57;
input n_66;
input n_21;
input n_31;
input n_8;
input n_312;
input n_183;
input n_266;
input n_205;
input n_335;
input n_177;
input n_313;
input n_22;
input n_140;
input n_219;
input n_180;
input n_212;
input n_210;
input n_325;
input n_338;
input n_103;
input n_166;
input n_224;
input n_151;
input n_130;
input n_253;
input n_99;
input n_15;
input n_72;
input n_152;
input n_198;
input n_7;
input n_228;
input n_272;
input n_196;
input n_315;
input n_123;
input n_279;
input n_79;
input n_270;
input n_305;
input n_117;
input n_208;
input n_215;
input n_135;
input n_70;
input n_50;
input n_170;
input n_86;
input n_340;
input n_13;
input n_168;
input n_175;
input n_241;
input n_105;
input n_84;
input n_294;
input n_258;
input n_206;
input n_307;
input n_342;
input n_14;
input n_194;
input n_137;
input n_225;
input n_16;
input n_39;
input n_337;
input n_247;
input n_240;
input n_38;
input n_259;
input n_143;
input n_192;
input n_0;
input n_264;
input n_63;
input n_1;
input n_237;
input n_91;
output n_344;
wire n_476;
wire n_887;
wire n_599;
wire n_1279;
wire n_1314;
wire n_830;
wire n_1371;
wire n_624;
wire n_618;
wire n_1797;
wire n_933;
wire n_485;
wire n_822;
wire n_750;
wire n_1641;
wire n_503;
wire n_1781;
wire n_1762;
wire n_1591;
wire n_469;
wire n_1310;
wire n_1376;
wire n_592;
wire n_1621;
wire n_1729;
wire n_1737;
wire n_761;
wire n_421;
wire n_919;
wire n_1217;
wire n_1423;
wire n_571;
wire n_549;
wire n_1034;
wire n_1328;
wire n_1219;
wire n_952;
wire n_1166;
wire n_752;
wire n_448;
wire n_556;
wire n_593;
wire n_989;
wire n_431;
wire n_1044;
wire n_1730;
wire n_1744;
wire n_963;
wire n_551;
wire n_884;
wire n_814;
wire n_944;
wire n_1283;
wire n_983;
wire n_955;
wire n_975;
wire n_941;
wire n_1313;
wire n_1468;
wire n_1713;
wire n_870;
wire n_1248;
wire n_1602;
wire n_548;
wire n_572;
wire n_815;
wire n_1140;
wire n_1453;
wire n_1520;
wire n_786;
wire n_512;
wire n_395;
wire n_795;
wire n_1379;
wire n_400;
wire n_1597;
wire n_1415;
wire n_1160;
wire n_1287;
wire n_883;
wire n_478;
wire n_1575;
wire n_1687;
wire n_553;
wire n_1805;
wire n_1367;
wire n_744;
wire n_1325;
wire n_1225;
wire n_1441;
wire n_875;
wire n_951;
wire n_1199;
wire n_1382;
wire n_1543;
wire n_791;
wire n_976;
wire n_636;
wire n_906;
wire n_477;
wire n_1477;
wire n_595;
wire n_1282;
wire n_683;
wire n_840;
wire n_570;
wire n_675;
wire n_835;
wire n_732;
wire n_784;
wire n_962;
wire n_1599;
wire n_755;
wire n_409;
wire n_781;
wire n_576;
wire n_1688;
wire n_956;
wire n_1242;
wire n_1537;
wire n_874;
wire n_796;
wire n_1126;
wire n_383;
wire n_1607;
wire n_455;
wire n_1771;
wire n_1809;
wire n_682;
wire n_1745;
wire n_812;
wire n_817;
wire n_782;
wire n_760;
wire n_608;
wire n_534;
wire n_1454;
wire n_708;
wire n_1020;
wire n_885;
wire n_950;
wire n_381;
wire n_1196;
wire n_1013;
wire n_808;
wire n_1639;
wire n_1224;
wire n_1694;
wire n_688;
wire n_1042;
wire n_1588;
wire n_363;
wire n_1317;
wire n_417;
wire n_690;
wire n_1419;
wire n_499;
wire n_1142;
wire n_1731;
wire n_1589;
wire n_947;
wire n_970;
wire n_1677;
wire n_1149;
wire n_368;
wire n_527;
wire n_1676;
wire n_1342;
wire n_1440;
wire n_552;
wire n_1346;
wire n_1383;
wire n_1675;
wire n_590;
wire n_1293;
wire n_432;
wire n_1131;
wire n_1008;
wire n_1491;
wire n_805;
wire n_1600;
wire n_619;
wire n_1095;
wire n_1250;
wire n_1284;
wire n_360;
wire n_1583;
wire n_1465;
wire n_859;
wire n_1486;
wire n_1304;
wire n_685;
wire n_1080;
wire n_917;
wire n_1247;
wire n_501;
wire n_488;
wire n_1380;
wire n_1658;
wire n_954;
wire n_702;
wire n_1007;
wire n_351;
wire n_898;
wire n_562;
wire n_1022;
wire n_1502;
wire n_404;
wire n_1073;
wire n_728;
wire n_1301;
wire n_1632;
wire n_1201;
wire n_997;
wire n_1768;
wire n_1105;
wire n_1243;
wire n_1003;
wire n_346;
wire n_749;
wire n_914;
wire n_1286;
wire n_494;
wire n_1661;
wire n_927;
wire n_723;
wire n_1351;
wire n_972;
wire n_1813;
wire n_1628;
wire n_1587;
wire n_1570;
wire n_1209;
wire n_411;
wire n_498;
wire n_765;
wire n_1397;
wire n_1554;
wire n_648;
wire n_1487;
wire n_939;
wire n_1615;
wire n_1763;
wire n_928;
wire n_1384;
wire n_789;
wire n_1515;
wire n_738;
wire n_1387;
wire n_922;
wire n_1048;
wire n_1422;
wire n_787;
wire n_1214;
wire n_806;
wire n_715;
wire n_1714;
wire n_420;
wire n_1666;
wire n_1490;
wire n_1258;
wire n_873;
wire n_438;
wire n_1814;
wire n_446;
wire n_1281;
wire n_1559;
wire n_1495;
wire n_1510;
wire n_1727;
wire n_712;
wire n_422;
wire n_861;
wire n_1574;
wire n_479;
wire n_825;
wire n_541;
wire n_839;
wire n_811;
wire n_558;
wire n_1742;
wire n_724;
wire n_1648;
wire n_440;
wire n_1231;
wire n_1305;
wire n_1161;
wire n_686;
wire n_1299;
wire n_949;
wire n_586;
wire n_1508;
wire n_1421;
wire n_788;
wire n_441;
wire n_1045;
wire n_1339;
wire n_1793;
wire n_837;
wire n_1349;
wire n_1708;
wire n_1445;
wire n_1631;
wire n_829;
wire n_1030;
wire n_1348;
wire n_375;
wire n_1391;
wire n_597;
wire n_1036;
wire n_687;
wire n_1751;
wire n_1765;
wire n_652;
wire n_1538;
wire n_500;
wire n_804;
wire n_1173;
wire n_854;
wire n_1787;
wire n_424;
wire n_877;
wire n_802;
wire n_1488;
wire n_1572;
wire n_1514;
wire n_480;
wire n_1652;
wire n_684;
wire n_1178;
wire n_1531;
wire n_821;
wire n_1657;
wire n_1616;
wire n_1563;
wire n_1018;
wire n_980;
wire n_1233;
wire n_1106;
wire n_1205;
wire n_838;
wire n_1561;
wire n_635;
wire n_792;
wire n_1392;
wire n_1542;
wire n_665;
wire n_667;
wire n_991;
wire n_1712;
wire n_1556;
wire n_580;
wire n_1004;
wire n_1370;
wire n_1417;
wire n_1703;
wire n_1717;
wire n_1723;
wire n_979;
wire n_445;
wire n_596;
wire n_1740;
wire n_1197;
wire n_657;
wire n_1260;
wire n_355;
wire n_1606;
wire n_1760;
wire n_1129;
wire n_1285;
wire n_742;
wire n_1014;
wire n_1385;
wire n_1629;
wire n_1618;
wire n_461;
wire n_1770;
wire n_1047;
wire n_1016;
wire n_1545;
wire n_694;
wire n_1350;
wire n_894;
wire n_1750;
wire n_545;
wire n_1459;
wire n_1530;
wire n_401;
wire n_538;
wire n_1594;
wire n_537;
wire n_1767;
wire n_1651;
wire n_560;
wire n_1094;
wire n_1776;
wire n_1719;
wire n_1220;
wire n_696;
wire n_1147;
wire n_1425;
wire n_1613;
wire n_1504;
wire n_704;
wire n_453;
wire n_647;
wire n_1499;
wire n_948;
wire n_399;
wire n_700;
wire n_677;
wire n_1269;
wire n_378;
wire n_591;
wire n_1635;
wire n_1518;
wire n_1702;
wire n_1366;
wire n_678;
wire n_415;
wire n_1400;
wire n_564;
wire n_638;
wire n_1361;
wire n_510;
wire n_1358;
wire n_1577;
wire n_1642;
wire n_1406;
wire n_550;
wire n_966;
wire n_1568;
wire n_1368;
wire n_994;
wire n_1612;
wire n_384;
wire n_1479;
wire n_1128;
wire n_1098;
wire n_824;
wire n_1238;
wire n_1611;
wire n_992;
wire n_813;
wire n_981;
wire n_1338;
wire n_1182;
wire n_872;
wire n_1401;
wire n_1086;
wire n_1070;
wire n_1189;
wire n_1665;
wire n_535;
wire n_882;
wire n_1741;
wire n_1210;
wire n_1456;
wire n_746;
wire n_656;
wire n_1614;
wire n_1148;
wire n_748;
wire n_860;
wire n_1261;
wire n_1062;
wire n_1439;
wire n_651;
wire n_1585;
wire n_1500;
wire n_801;
wire n_1271;
wire n_1653;
wire n_529;
wire n_504;
wire n_973;
wire n_1364;
wire n_659;
wire n_634;
wire n_903;
wire n_1668;
wire n_565;
wire n_925;
wire n_1389;
wire n_1393;
wire n_457;
wire n_1121;
wire n_1059;
wire n_493;
wire n_1362;
wire n_610;
wire n_1035;
wire n_620;
wire n_722;
wire n_1174;
wire n_1193;
wire n_1553;
wire n_754;
wire n_508;
wire n_1141;
wire n_1769;
wire n_1812;
wire n_1112;
wire n_1485;
wire n_1408;
wire n_1680;
wire n_428;
wire n_783;
wire n_1107;
wire n_1564;
wire n_505;
wire n_600;
wire n_731;
wire n_964;
wire n_605;
wire n_1516;
wire n_1386;
wire n_406;
wire n_1493;
wire n_1579;
wire n_617;
wire n_602;
wire n_402;
wire n_733;
wire n_1404;
wire n_658;
wire n_676;
wire n_531;
wire n_1031;
wire n_1394;
wire n_807;
wire n_1011;
wire n_416;
wire n_1567;
wire n_895;
wire n_1569;
wire n_799;
wire n_490;
wire n_391;
wire n_695;
wire n_1181;
wire n_881;
wire n_1626;
wire n_645;
wire n_1145;
wire n_1529;
wire n_557;
wire n_1681;
wire n_1620;
wire n_777;
wire n_985;
wire n_1659;
wire n_910;
wire n_642;
wire n_613;
wire n_1773;
wire n_1125;
wire n_1347;
wire n_1655;
wire n_1766;
wire n_1522;
wire n_1163;
wire n_1278;
wire n_734;
wire n_1623;
wire n_735;
wire n_1179;
wire n_569;
wire n_1171;
wire n_785;
wire n_1203;
wire n_1716;
wire n_1232;
wire n_471;
wire n_853;
wire n_810;
wire n_1136;
wire n_699;
wire n_1187;
wire n_1000;
wire n_1580;
wire n_649;
wire n_358;
wire n_1234;
wire n_622;
wire n_1634;
wire n_1002;
wire n_1353;
wire n_1165;
wire n_1551;
wire n_1667;
wire n_1058;
wire n_1216;
wire n_662;
wire n_850;
wire n_354;
wire n_720;
wire n_1026;
wire n_1756;
wire n_1803;
wire n_492;
wire n_407;
wire n_419;
wire n_1023;
wire n_730;
wire n_1699;
wire n_1794;
wire n_1748;
wire n_643;
wire n_1403;
wire n_486;
wire n_779;
wire n_481;
wire n_691;
wire n_589;
wire n_365;
wire n_526;
wire n_1513;
wire n_1194;
wire n_389;
wire n_1609;
wire n_1462;
wire n_701;
wire n_809;
wire n_1532;
wire n_520;
wire n_679;
wire n_926;
wire n_1643;
wire n_942;
wire n_1374;
wire n_1120;
wire n_1497;
wire n_1784;
wire n_1548;
wire n_1526;
wire n_689;
wire n_1483;
wire n_946;
wire n_1409;
wire n_753;
wire n_1188;
wire n_623;
wire n_1032;
wire n_1474;
wire n_721;
wire n_1431;
wire n_1806;
wire n_1133;
wire n_1775;
wire n_1593;
wire n_739;
wire n_1322;
wire n_1525;
wire n_1732;
wire n_1162;
wire n_1463;
wire n_762;
wire n_1524;
wire n_1298;
wire n_442;
wire n_1633;
wire n_740;
wire n_1686;
wire n_1357;
wire n_639;
wire n_1186;
wire n_1365;
wire n_1807;
wire n_459;
wire n_1172;
wire n_998;
wire n_1689;
wire n_1625;
wire n_1395;
wire n_1276;
wire n_836;
wire n_1733;
wire n_1184;
wire n_583;
wire n_347;
wire n_414;
wire n_1336;
wire n_776;
wire n_1138;
wire n_890;
wire n_1306;
wire n_1413;
wire n_1783;
wire n_1759;
wire n_1266;
wire n_497;
wire n_911;
wire n_450;
wire n_1578;
wire n_1779;
wire n_473;
wire n_967;
wire n_1709;
wire n_474;
wire n_1159;
wire n_1315;
wire n_1055;
wire n_611;
wire n_380;
wire n_1576;
wire n_844;
wire n_968;
wire n_710;
wire n_1040;
wire n_1102;
wire n_661;
wire n_1185;
wire n_447;
wire n_1795;
wire n_403;
wire n_1039;
wire n_1119;
wire n_574;
wire n_1451;
wire n_1069;
wire n_842;
wire n_1788;
wire n_798;
wire n_1700;
wire n_668;
wire n_862;
wire n_869;
wire n_1811;
wire n_1066;
wire n_1377;
wire n_800;
wire n_1170;
wire n_778;
wire n_1175;
wire n_522;
wire n_1475;
wire n_943;
wire n_977;
wire n_357;
wire n_905;
wire n_386;
wire n_878;
wire n_1734;
wire n_1333;
wire n_577;
wire n_1610;
wire n_759;
wire n_1235;
wire n_900;
wire n_841;
wire n_1724;
wire n_1218;
wire n_736;
wire n_1706;
wire n_766;
wire n_1113;
wire n_852;
wire n_1268;
wire n_1695;
wire n_1089;
wire n_1122;
wire n_908;
wire n_1123;
wire n_923;
wire n_1302;
wire n_1289;
wire n_937;
wire n_1442;
wire n_773;
wire n_353;
wire n_1446;
wire n_1778;
wire n_865;
wire n_1644;
wire n_1736;
wire n_1707;
wire n_856;
wire n_594;
wire n_1146;
wire n_1685;
wire n_1810;
wire n_1435;
wire n_1800;
wire n_374;
wire n_932;
wire n_958;
wire n_1755;
wire n_775;
wire n_763;
wire n_1093;
wire n_427;
wire n_1540;
wire n_519;
wire n_1116;
wire n_709;
wire n_388;
wire n_1470;
wire n_816;
wire n_625;
wire n_953;
wire n_1565;
wire n_1373;
wire n_1558;
wire n_716;
wire n_1683;
wire n_356;
wire n_584;
wire n_896;
wire n_1722;
wire n_528;
wire n_1078;
wire n_495;
wire n_1072;
wire n_1638;
wire n_370;
wire n_1663;
wire n_352;
wire n_935;
wire n_1505;
wire n_467;
wire n_1213;
wire n_1053;
wire n_515;
wire n_1019;
wire n_680;
wire n_1180;
wire n_904;
wire n_920;
wire n_1117;
wire n_1168;
wire n_1598;
wire n_1309;
wire n_909;
wire n_996;
wire n_523;
wire n_439;
wire n_506;
wire n_606;
wire n_513;
wire n_1332;
wire n_1263;
wire n_1411;
wire n_1115;
wire n_725;
wire n_960;
wire n_671;
wire n_1084;
wire n_1726;
wire n_1656;
wire n_454;
wire n_1303;
wire n_1471;
wire n_443;
wire n_1029;
wire n_345;
wire n_1207;
wire n_1555;
wire n_664;
wire n_367;
wire n_1017;
wire n_581;
wire n_936;
wire n_1215;
wire n_582;
wire n_641;
wire n_1738;
wire n_940;
wire n_745;
wire n_1608;
wire n_1167;
wire n_1327;
wire n_609;
wire n_1743;
wire n_1752;
wire n_1792;
wire n_1006;
wire n_1259;
wire n_350;
wire n_561;
wire n_437;
wire n_1560;
wire n_405;
wire n_1223;
wire n_621;
wire n_1012;
wire n_1241;
wire n_1414;
wire n_1671;
wire n_502;
wire n_434;
wire n_769;
wire n_1212;
wire n_1455;
wire n_1054;
wire n_1669;
wire n_1308;
wire n_1050;
wire n_426;
wire n_1550;
wire n_1134;
wire n_1670;
wire n_1319;
wire n_1363;
wire n_616;
wire n_880;
wire n_1103;
wire n_1274;
wire n_832;
wire n_1321;
wire n_1429;
wire n_1660;
wire n_1060;
wire n_1154;
wire n_1786;
wire n_361;
wire n_632;
wire n_1344;
wire n_1450;
wire n_1603;
wire n_1720;
wire n_714;
wire n_1331;
wire n_1222;
wire n_1041;
wire n_1764;
wire n_1512;
wire n_957;
wire n_1255;
wire n_995;
wire n_1124;
wire n_1335;
wire n_1405;
wire n_912;
wire n_464;
wire n_1227;
wire n_1509;
wire n_945;
wire n_392;
wire n_563;
wire n_891;
wire n_568;
wire n_1586;
wire n_413;
wire n_1157;
wire n_902;
wire n_1749;
wire n_1158;
wire n_1079;
wire n_1330;
wire n_1033;
wire n_1464;
wire n_1028;
wire n_366;
wire n_727;
wire n_1083;
wire n_397;
wire n_1056;
wire n_1605;
wire n_1592;
wire n_1802;
wire n_663;
wire n_588;
wire n_1682;
wire n_1698;
wire n_1448;
wire n_707;
wire n_915;
wire n_1774;
wire n_1785;
wire n_1001;
wire n_1418;
wire n_711;
wire n_864;
wire n_1782;
wire n_1169;
wire n_377;
wire n_1139;
wire n_1482;
wire n_1798;
wire n_1038;
wire n_1085;
wire n_845;
wire n_1673;
wire n_1619;
wire n_1127;
wire n_1718;
wire n_484;
wire n_893;
wire n_1068;
wire n_747;
wire n_1672;
wire n_1753;
wire n_1244;
wire n_1581;
wire n_697;
wire n_978;
wire n_847;
wire n_1452;
wire n_826;
wire n_373;
wire n_628;
wire n_487;
wire n_831;
wire n_1772;
wire n_653;
wire n_1725;
wire n_692;
wire n_1433;
wire n_1051;
wire n_1696;
wire n_1355;
wire n_1494;
wire n_1517;
wire n_827;
wire n_472;
wire n_866;
wire n_452;
wire n_630;
wire n_820;
wire n_1208;
wire n_612;
wire n_1426;
wire n_858;
wire n_764;
wire n_741;
wire n_1090;
wire n_456;
wire n_359;
wire n_1469;
wire n_1164;
wire n_433;
wire n_627;
wire n_1693;
wire n_1791;
wire n_418;
wire n_771;
wire n_524;
wire n_1378;
wire n_1496;
wire n_705;
wire n_1191;
wire n_1206;
wire n_1270;
wire n_1566;
wire n_1399;
wire n_546;
wire n_1010;
wire n_1375;
wire n_1015;
wire n_1761;
wire n_863;
wire n_525;
wire n_1790;
wire n_1226;
wire n_1617;
wire n_644;
wire n_1150;
wire n_1341;
wire n_833;
wire n_1229;
wire n_1690;
wire n_1143;
wire n_929;
wire n_1190;
wire n_1728;
wire n_543;
wire n_1710;
wire n_585;
wire n_1457;
wire n_719;
wire n_1343;
wire n_465;
wire n_1604;
wire n_1156;
wire n_988;
wire n_1757;
wire n_1466;
wire n_921;
wire n_1396;
wire n_1799;
wire n_640;
wire n_1176;
wire n_1721;
wire n_1691;
wire n_1511;
wire n_1151;
wire n_1501;
wire n_1254;
wire n_1458;
wire n_646;
wire n_650;
wire n_1211;
wire n_743;
wire n_823;
wire n_393;
wire n_1804;
wire n_1480;
wire n_1101;
wire n_1251;
wire n_1076;
wire n_1434;
wire n_1461;
wire n_1449;
wire n_1715;
wire n_1407;
wire n_1104;
wire n_1061;
wire n_849;
wire n_554;
wire n_1153;
wire n_1337;
wire n_797;
wire n_1704;
wire n_1177;
wire n_758;
wire n_436;
wire n_390;
wire n_1096;
wire n_1316;
wire n_1590;
wire n_1420;
wire n_1552;
wire n_1544;
wire n_1571;
wire n_1092;
wire n_846;
wire n_631;
wire n_673;
wire n_1410;
wire n_1067;
wire n_518;
wire n_1292;
wire n_1192;
wire n_1478;
wire n_1507;
wire n_1240;
wire n_1789;
wire n_987;
wire n_1596;
wire n_362;
wire n_1065;
wire n_1064;
wire n_540;
wire n_1075;
wire n_718;
wire n_669;
wire n_1091;
wire n_423;
wire n_1221;
wire n_458;
wire n_1777;
wire n_444;
wire n_1200;
wire n_364;
wire n_555;
wire n_1295;
wire n_974;
wire n_1329;
wire n_857;
wire n_1424;
wire n_1674;
wire n_376;
wire n_491;
wire n_1294;
wire n_1110;
wire n_1137;
wire n_1533;
wire n_460;
wire n_1679;
wire n_1595;
wire n_1735;
wire n_666;
wire n_660;
wire n_1359;
wire n_886;
wire n_767;
wire n_889;
wire n_1398;
wire n_379;
wire n_1432;
wire n_1021;
wire n_1297;
wire n_1046;
wire n_1109;
wire n_961;
wire n_1447;
wire n_489;
wire n_1622;
wire n_1381;
wire n_1582;
wire n_1747;
wire n_573;
wire n_1099;
wire n_1654;
wire n_626;
wire n_539;
wire n_462;
wire n_615;
wire n_1118;
wire n_990;
wire n_1108;
wire n_670;
wire n_818;
wire n_918;
wire n_1272;
wire n_1541;
wire n_408;
wire n_1754;
wire n_372;
wire n_578;
wire n_892;
wire n_938;
wire n_774;
wire n_559;
wire n_1049;
wire n_466;
wire n_1277;
wire n_1584;
wire n_984;
wire n_726;
wire n_369;
wire n_517;
wire n_931;
wire n_780;
wire n_530;
wire n_834;
wire n_693;
wire n_496;
wire n_1360;
wire n_1082;
wire n_1257;
wire n_468;
wire n_532;
wire n_1025;
wire n_924;
wire n_1264;
wire n_1527;
wire n_1245;
wire n_1152;
wire n_1539;
wire n_1081;
wire n_547;
wire n_1324;
wire n_1198;
wire n_1678;
wire n_1307;
wire n_993;
wire n_819;
wire n_737;
wire n_1489;
wire n_1637;
wire n_1290;
wire n_1318;
wire n_1135;
wire n_1063;
wire n_828;
wire n_770;
wire n_867;
wire n_398;
wire n_1100;
wire n_1519;
wire n_425;
wire n_1650;
wire n_879;
wire n_1640;
wire n_449;
wire n_1340;
wire n_1562;
wire n_607;
wire n_629;
wire n_706;
wire n_901;
wire n_876;
wire n_1443;
wire n_655;
wire n_654;
wire n_1521;
wire n_672;
wire n_567;
wire n_916;
wire n_1354;
wire n_1780;
wire n_1547;
wire n_1334;
wire n_1291;
wire n_1437;
wire n_1473;
wire n_986;
wire n_451;
wire n_1037;
wire n_1267;
wire n_790;
wire n_1262;
wire n_410;
wire n_1684;
wire n_1444;
wire n_751;
wire n_999;
wire n_913;
wire n_1237;
wire n_1506;
wire n_1356;
wire n_1646;
wire n_768;
wire n_412;
wire n_542;
wire n_1256;
wire n_1427;
wire n_1077;
wire n_1111;
wire n_1503;
wire n_1249;
wire n_1416;
wire n_387;
wire n_1239;
wire n_1796;
wire n_1662;
wire n_969;
wire n_1535;
wire n_1009;
wire n_1202;
wire n_1498;
wire n_1801;
wire n_1549;
wire n_604;
wire n_848;
wire n_756;
wire n_713;
wire n_598;
wire n_430;
wire n_1252;
wire n_1647;
wire n_1132;
wire n_1649;
wire n_1275;
wire n_843;
wire n_579;
wire n_533;
wire n_1472;
wire n_385;
wire n_536;
wire n_470;
wire n_851;
wire n_1155;
wire n_934;
wire n_1636;
wire n_1027;
wire n_965;
wire n_1296;
wire n_382;
wire n_1484;
wire n_1043;
wire n_435;
wire n_511;
wire n_1808;
wire n_1492;
wire n_1467;
wire n_509;
wire n_1204;
wire n_930;
wire n_1265;
wire n_1057;
wire n_907;
wire n_1430;
wire n_1481;
wire n_1758;
wire n_1005;
wire n_1312;
wire n_1697;
wire n_899;
wire n_637;
wire n_544;
wire n_1476;
wire n_1087;
wire n_1536;
wire n_1746;
wire n_1711;
wire n_482;
wire n_633;
wire n_971;
wire n_1052;
wire n_1071;
wire n_1311;
wire n_1601;
wire n_1438;
wire n_1273;
wire n_959;
wire n_349;
wire n_1573;
wire n_1130;
wire n_794;
wire n_1228;
wire n_681;
wire n_982;
wire n_717;
wire n_1624;
wire n_1253;
wire n_1183;
wire n_516;
wire n_1460;
wire n_521;
wire n_1195;
wire n_575;
wire n_1300;
wire n_1372;
wire n_698;
wire n_371;
wire n_1345;
wire n_587;
wire n_1701;
wire n_1664;
wire n_1428;
wire n_1246;
wire n_1074;
wire n_674;
wire n_888;
wire n_1546;
wire n_1436;
wire n_793;
wire n_1390;
wire n_1815;
wire n_1412;
wire n_757;
wire n_1534;
wire n_803;
wire n_514;
wire n_507;
wire n_1557;
wire n_614;
wire n_772;
wire n_1114;
wire n_566;
wire n_871;
wire n_1739;
wire n_1088;
wire n_1230;
wire n_1326;
wire n_1402;
wire n_1388;
wire n_483;
wire n_1630;
wire n_394;
wire n_729;
wire n_1280;
wire n_1323;
wire n_1352;
wire n_703;
wire n_1369;
wire n_1097;
wire n_601;
wire n_463;
wire n_396;
wire n_1236;
wire n_1523;
wire n_348;
wire n_1528;
wire n_603;
wire n_1692;
wire n_1288;
wire n_868;
wire n_1705;
wire n_1024;
wire n_1144;
wire n_1627;
wire n_475;
wire n_897;
wire n_1320;
wire n_855;
wire n_1645;
wire n_429;
AOI22xp33_ASAP7_75t_L g1527 ( .A1(n_0), .A2(n_88), .B1(n_1494), .B2(n_1499), .Y(n_1527) );
INVx1_ASAP7_75t_L g1395 ( .A(n_1), .Y(n_1395) );
AO22x1_ASAP7_75t_L g1419 ( .A1(n_1), .A2(n_219), .B1(n_486), .B2(n_1341), .Y(n_1419) );
INVx1_ASAP7_75t_L g359 ( .A(n_2), .Y(n_359) );
AND2x2_ASAP7_75t_L g460 ( .A(n_2), .B(n_461), .Y(n_460) );
AND2x2_ASAP7_75t_L g492 ( .A(n_2), .B(n_243), .Y(n_492) );
NOR2xp33_ASAP7_75t_L g921 ( .A(n_2), .B(n_369), .Y(n_921) );
INVx1_ASAP7_75t_L g1404 ( .A(n_3), .Y(n_1404) );
AOI22xp33_ASAP7_75t_L g1418 ( .A1(n_3), .A2(n_117), .B1(n_491), .B2(n_654), .Y(n_1418) );
AOI22xp33_ASAP7_75t_SL g555 ( .A1(n_4), .A2(n_302), .B1(n_410), .B2(n_533), .Y(n_555) );
AOI221xp5_ASAP7_75t_L g582 ( .A1(n_4), .A2(n_5), .B1(n_583), .B2(n_585), .C(n_588), .Y(n_582) );
AOI22xp33_ASAP7_75t_SL g565 ( .A1(n_5), .A2(n_10), .B1(n_406), .B2(n_424), .Y(n_565) );
AOI22xp33_ASAP7_75t_SL g403 ( .A1(n_6), .A2(n_298), .B1(n_404), .B2(n_410), .Y(n_403) );
AOI221xp5_ASAP7_75t_L g471 ( .A1(n_6), .A2(n_252), .B1(n_472), .B2(n_476), .C(n_480), .Y(n_471) );
INVx1_ASAP7_75t_L g1106 ( .A(n_7), .Y(n_1106) );
XOR2x2_ASAP7_75t_L g1178 ( .A(n_8), .B(n_1179), .Y(n_1178) );
INVx1_ASAP7_75t_L g1295 ( .A(n_9), .Y(n_1295) );
OAI22xp5_ASAP7_75t_L g1311 ( .A1(n_9), .A2(n_330), .B1(n_519), .B2(n_704), .Y(n_1311) );
A2O1A1Ixp33_ASAP7_75t_L g600 ( .A1(n_10), .A2(n_601), .B(n_605), .C(n_611), .Y(n_600) );
OAI22xp5_ASAP7_75t_L g1173 ( .A1(n_11), .A2(n_207), .B1(n_438), .B2(n_689), .Y(n_1173) );
INVx1_ASAP7_75t_L g853 ( .A(n_12), .Y(n_853) );
AOI22xp33_ASAP7_75t_SL g1727 ( .A1(n_13), .A2(n_211), .B1(n_422), .B2(n_636), .Y(n_1727) );
INVxp67_ASAP7_75t_SL g1750 ( .A(n_13), .Y(n_1750) );
AOI221xp5_ASAP7_75t_L g865 ( .A1(n_14), .A2(n_292), .B1(n_736), .B2(n_866), .C(n_867), .Y(n_865) );
AOI22xp33_ASAP7_75t_SL g885 ( .A1(n_14), .A2(n_312), .B1(n_383), .B2(n_427), .Y(n_885) );
AOI22xp33_ASAP7_75t_L g643 ( .A1(n_15), .A2(n_277), .B1(n_640), .B2(n_644), .Y(n_643) );
AOI221xp5_ASAP7_75t_L g652 ( .A1(n_15), .A2(n_80), .B1(n_653), .B2(n_654), .C(n_655), .Y(n_652) );
AOI22xp33_ASAP7_75t_L g764 ( .A1(n_16), .A2(n_314), .B1(n_590), .B2(n_765), .Y(n_764) );
INVx1_ASAP7_75t_L g784 ( .A(n_16), .Y(n_784) );
CKINVDCx5p33_ASAP7_75t_R g1767 ( .A(n_17), .Y(n_1767) );
INVx2_ASAP7_75t_L g400 ( .A(n_18), .Y(n_400) );
INVx1_ASAP7_75t_L g805 ( .A(n_19), .Y(n_805) );
OAI222xp33_ASAP7_75t_L g835 ( .A1(n_19), .A2(n_165), .B1(n_666), .B2(n_687), .C1(n_836), .C2(n_841), .Y(n_835) );
INVx1_ASAP7_75t_L g1152 ( .A(n_20), .Y(n_1152) );
AOI22xp33_ASAP7_75t_L g642 ( .A1(n_21), .A2(n_215), .B1(n_427), .B2(n_638), .Y(n_642) );
AOI22xp33_ASAP7_75t_L g656 ( .A1(n_21), .A2(n_135), .B1(n_657), .B2(n_659), .Y(n_656) );
INVx1_ASAP7_75t_L g1480 ( .A(n_22), .Y(n_1480) );
AOI22xp33_ASAP7_75t_L g868 ( .A1(n_23), .A2(n_256), .B1(n_483), .B2(n_592), .Y(n_868) );
AOI22xp33_ASAP7_75t_L g887 ( .A1(n_23), .A2(n_253), .B1(n_645), .B2(n_888), .Y(n_887) );
AOI22xp5_ASAP7_75t_L g1708 ( .A1(n_24), .A2(n_1709), .B1(n_1710), .B2(n_1752), .Y(n_1708) );
CKINVDCx14_ASAP7_75t_R g1752 ( .A(n_24), .Y(n_1752) );
INVx1_ASAP7_75t_L g1150 ( .A(n_25), .Y(n_1150) );
AOI22xp33_ASAP7_75t_L g1164 ( .A1(n_25), .A2(n_63), .B1(n_1165), .B2(n_1166), .Y(n_1164) );
OAI22xp5_ASAP7_75t_L g1059 ( .A1(n_26), .A2(n_293), .B1(n_519), .B2(n_704), .Y(n_1059) );
CKINVDCx5p33_ASAP7_75t_R g692 ( .A(n_27), .Y(n_692) );
HB1xp67_ASAP7_75t_L g354 ( .A(n_28), .Y(n_354) );
AND2x2_ASAP7_75t_L g1495 ( .A(n_28), .B(n_352), .Y(n_1495) );
OAI22xp5_ASAP7_75t_SL g1454 ( .A1(n_29), .A2(n_278), .B1(n_1184), .B2(n_1196), .Y(n_1454) );
INVxp67_ASAP7_75t_SL g1483 ( .A(n_29), .Y(n_1483) );
AOI22xp33_ASAP7_75t_L g1051 ( .A1(n_30), .A2(n_209), .B1(n_427), .B2(n_1049), .Y(n_1051) );
AOI221xp5_ASAP7_75t_L g1078 ( .A1(n_30), .A2(n_305), .B1(n_507), .B2(n_1079), .C(n_1081), .Y(n_1078) );
CKINVDCx5p33_ASAP7_75t_R g1713 ( .A(n_31), .Y(n_1713) );
INVxp67_ASAP7_75t_L g377 ( .A(n_32), .Y(n_377) );
AOI22xp5_ASAP7_75t_L g874 ( .A1(n_33), .A2(n_312), .B1(n_483), .B2(n_765), .Y(n_874) );
AOI22xp5_ASAP7_75t_L g886 ( .A1(n_33), .A2(n_292), .B1(n_427), .B2(n_812), .Y(n_886) );
AOI22xp33_ASAP7_75t_L g1012 ( .A1(n_34), .A2(n_50), .B1(n_390), .B2(n_953), .Y(n_1012) );
INVx1_ASAP7_75t_L g1022 ( .A(n_34), .Y(n_1022) );
AOI22xp33_ASAP7_75t_L g1526 ( .A1(n_35), .A2(n_62), .B1(n_1502), .B2(n_1511), .Y(n_1526) );
INVx1_ASAP7_75t_L g1045 ( .A(n_36), .Y(n_1045) );
OAI221xp5_ASAP7_75t_L g1071 ( .A1(n_36), .A2(n_234), .B1(n_742), .B2(n_1072), .C(n_1073), .Y(n_1071) );
INVx1_ASAP7_75t_L g930 ( .A(n_37), .Y(n_930) );
INVx1_ASAP7_75t_L g832 ( .A(n_38), .Y(n_832) );
AOI22xp5_ASAP7_75t_L g896 ( .A1(n_39), .A2(n_46), .B1(n_897), .B2(n_898), .Y(n_896) );
AOI22xp33_ASAP7_75t_L g951 ( .A1(n_39), .A2(n_157), .B1(n_427), .B2(n_952), .Y(n_951) );
AOI22xp33_ASAP7_75t_L g556 ( .A1(n_40), .A2(n_91), .B1(n_389), .B2(n_557), .Y(n_556) );
AOI221xp5_ASAP7_75t_L g606 ( .A1(n_40), .A2(n_190), .B1(n_476), .B2(n_607), .C(n_608), .Y(n_606) );
AOI221xp5_ASAP7_75t_L g1001 ( .A1(n_41), .A2(n_333), .B1(n_412), .B2(n_1002), .C(n_1003), .Y(n_1001) );
AOI221xp5_ASAP7_75t_L g1020 ( .A1(n_41), .A2(n_113), .B1(n_736), .B2(n_761), .C(n_1021), .Y(n_1020) );
INVx1_ASAP7_75t_L g768 ( .A(n_42), .Y(n_768) );
AOI22xp33_ASAP7_75t_L g1725 ( .A1(n_43), .A2(n_273), .B1(n_426), .B2(n_1361), .Y(n_1725) );
INVx1_ASAP7_75t_L g1744 ( .A(n_43), .Y(n_1744) );
OAI21xp5_ASAP7_75t_L g878 ( .A1(n_44), .A2(n_703), .B(n_879), .Y(n_878) );
NAND5xp2_ASAP7_75t_L g1333 ( .A(n_45), .B(n_1334), .C(n_1357), .D(n_1367), .E(n_1372), .Y(n_1333) );
INVx1_ASAP7_75t_L g1380 ( .A(n_45), .Y(n_1380) );
AOI22xp33_ASAP7_75t_SL g942 ( .A1(n_46), .A2(n_168), .B1(n_943), .B2(n_944), .Y(n_942) );
INVx1_ASAP7_75t_L g767 ( .A(n_47), .Y(n_767) );
INVx1_ASAP7_75t_L g831 ( .A(n_48), .Y(n_831) );
AOI22xp33_ASAP7_75t_L g1300 ( .A1(n_49), .A2(n_179), .B1(n_485), .B2(n_499), .Y(n_1300) );
AOI22xp33_ASAP7_75t_SL g1319 ( .A1(n_49), .A2(n_307), .B1(n_645), .B2(n_1320), .Y(n_1319) );
INVx1_ASAP7_75t_L g1017 ( .A(n_50), .Y(n_1017) );
BUFx6f_ASAP7_75t_L g366 ( .A(n_51), .Y(n_366) );
XOR2x2_ASAP7_75t_L g1287 ( .A(n_52), .B(n_1288), .Y(n_1287) );
AOI22xp5_ASAP7_75t_L g1510 ( .A1(n_52), .A2(n_110), .B1(n_1502), .B2(n_1511), .Y(n_1510) );
AOI22xp5_ASAP7_75t_L g1518 ( .A1(n_53), .A2(n_247), .B1(n_1502), .B2(n_1511), .Y(n_1518) );
INVx1_ASAP7_75t_L g1721 ( .A(n_54), .Y(n_1721) );
INVx1_ASAP7_75t_L g629 ( .A(n_55), .Y(n_629) );
OAI222xp33_ASAP7_75t_L g665 ( .A1(n_55), .A2(n_342), .B1(n_666), .B2(n_667), .C1(n_678), .C2(n_686), .Y(n_665) );
CKINVDCx5p33_ASAP7_75t_R g664 ( .A(n_56), .Y(n_664) );
AOI221xp5_ASAP7_75t_L g1339 ( .A1(n_57), .A2(n_166), .B1(n_491), .B2(n_654), .C(n_867), .Y(n_1339) );
AOI22xp33_ASAP7_75t_L g1362 ( .A1(n_57), .A2(n_226), .B1(n_427), .B2(n_1218), .Y(n_1362) );
CKINVDCx5p33_ASAP7_75t_R g576 ( .A(n_58), .Y(n_576) );
AOI22xp33_ASAP7_75t_L g1340 ( .A1(n_59), .A2(n_226), .B1(n_765), .B2(n_1341), .Y(n_1340) );
AOI22xp33_ASAP7_75t_L g1360 ( .A1(n_59), .A2(n_166), .B1(n_427), .B2(n_1361), .Y(n_1360) );
INVx1_ASAP7_75t_L g1193 ( .A(n_60), .Y(n_1193) );
AOI22xp33_ASAP7_75t_L g425 ( .A1(n_61), .A2(n_154), .B1(n_382), .B2(n_426), .Y(n_425) );
AOI21xp33_ASAP7_75t_L g504 ( .A1(n_61), .A2(n_505), .B(n_507), .Y(n_504) );
AOI22xp5_ASAP7_75t_L g854 ( .A1(n_62), .A2(n_855), .B1(n_856), .B2(n_890), .Y(n_854) );
INVxp67_ASAP7_75t_SL g890 ( .A(n_62), .Y(n_890) );
INVx1_ASAP7_75t_L g1139 ( .A(n_63), .Y(n_1139) );
INVx1_ASAP7_75t_L g552 ( .A(n_64), .Y(n_552) );
AOI221xp5_ASAP7_75t_L g899 ( .A1(n_65), .A2(n_317), .B1(n_900), .B2(n_901), .C(n_903), .Y(n_899) );
AOI221xp5_ASAP7_75t_L g947 ( .A1(n_65), .A2(n_280), .B1(n_790), .B2(n_948), .C(n_950), .Y(n_947) );
AOI22xp33_ASAP7_75t_SL g1723 ( .A1(n_66), .A2(n_169), .B1(n_404), .B2(n_790), .Y(n_1723) );
INVxp67_ASAP7_75t_SL g1747 ( .A(n_66), .Y(n_1747) );
OAI211xp5_ASAP7_75t_SL g992 ( .A1(n_67), .A2(n_962), .B(n_969), .C(n_993), .Y(n_992) );
INVx1_ASAP7_75t_L g1027 ( .A(n_67), .Y(n_1027) );
CKINVDCx5p33_ASAP7_75t_R g1776 ( .A(n_68), .Y(n_1776) );
INVx1_ASAP7_75t_L g863 ( .A(n_69), .Y(n_863) );
OAI22xp5_ASAP7_75t_L g1226 ( .A1(n_70), .A2(n_241), .B1(n_1227), .B2(n_1231), .Y(n_1226) );
OAI22xp5_ASAP7_75t_L g1264 ( .A1(n_70), .A2(n_241), .B1(n_1265), .B2(n_1267), .Y(n_1264) );
CKINVDCx5p33_ASAP7_75t_R g436 ( .A(n_71), .Y(n_436) );
OAI21xp5_ASAP7_75t_SL g518 ( .A1(n_72), .A2(n_519), .B(n_531), .Y(n_518) );
CKINVDCx5p33_ASAP7_75t_R g1348 ( .A(n_73), .Y(n_1348) );
AOI22xp33_ASAP7_75t_L g1098 ( .A1(n_74), .A2(n_223), .B1(n_636), .B2(n_946), .Y(n_1098) );
AOI22xp33_ASAP7_75t_SL g1123 ( .A1(n_74), .A2(n_276), .B1(n_502), .B2(n_590), .Y(n_1123) );
INVxp67_ASAP7_75t_SL g935 ( .A(n_75), .Y(n_935) );
OAI22xp5_ASAP7_75t_L g954 ( .A1(n_75), .A2(n_327), .B1(n_955), .B2(n_958), .Y(n_954) );
AOI22xp33_ASAP7_75t_SL g1052 ( .A1(n_76), .A2(n_335), .B1(n_645), .B2(n_1053), .Y(n_1052) );
AOI221xp5_ASAP7_75t_L g1065 ( .A1(n_76), .A2(n_141), .B1(n_480), .B2(n_495), .C(n_1066), .Y(n_1065) );
AOI22xp33_ASAP7_75t_L g1533 ( .A1(n_77), .A2(n_235), .B1(n_1502), .B2(n_1511), .Y(n_1533) );
AOI22xp33_ASAP7_75t_SL g421 ( .A1(n_78), .A2(n_252), .B1(n_406), .B2(n_422), .Y(n_421) );
AOI22xp33_ASAP7_75t_L g498 ( .A1(n_78), .A2(n_298), .B1(n_499), .B2(n_502), .Y(n_498) );
INVx1_ASAP7_75t_L g864 ( .A(n_79), .Y(n_864) );
AOI22xp33_ASAP7_75t_L g637 ( .A1(n_80), .A2(n_124), .B1(n_638), .B2(n_640), .Y(n_637) );
AOI22xp5_ASAP7_75t_L g1493 ( .A1(n_81), .A2(n_242), .B1(n_1494), .B2(n_1499), .Y(n_1493) );
AOI22xp33_ASAP7_75t_SL g1097 ( .A1(n_82), .A2(n_214), .B1(n_944), .B2(n_1095), .Y(n_1097) );
INVx1_ASAP7_75t_L g1118 ( .A(n_82), .Y(n_1118) );
AOI22xp33_ASAP7_75t_SL g1457 ( .A1(n_83), .A2(n_156), .B1(n_486), .B2(n_829), .Y(n_1457) );
INVxp67_ASAP7_75t_SL g1476 ( .A(n_83), .Y(n_1476) );
AOI22xp5_ASAP7_75t_L g1501 ( .A1(n_84), .A2(n_101), .B1(n_1502), .B2(n_1504), .Y(n_1501) );
AO22x1_ASAP7_75t_L g1524 ( .A1(n_85), .A2(n_249), .B1(n_1494), .B2(n_1499), .Y(n_1524) );
AOI22xp33_ASAP7_75t_L g728 ( .A1(n_86), .A2(n_265), .B1(n_645), .B2(n_718), .Y(n_728) );
AOI221xp5_ASAP7_75t_L g735 ( .A1(n_86), .A2(n_262), .B1(n_584), .B2(n_588), .C(n_736), .Y(n_735) );
OAI21xp33_ASAP7_75t_L g688 ( .A1(n_87), .A2(n_689), .B(n_690), .Y(n_688) );
OAI22xp5_ASAP7_75t_L g1786 ( .A1(n_89), .A2(n_260), .B1(n_1787), .B2(n_1788), .Y(n_1786) );
OAI22xp5_ASAP7_75t_SL g1802 ( .A1(n_89), .A2(n_130), .B1(n_1233), .B2(n_1250), .Y(n_1802) );
INVx1_ASAP7_75t_L g716 ( .A(n_90), .Y(n_716) );
AOI22xp33_ASAP7_75t_L g737 ( .A1(n_90), .A2(n_284), .B1(n_499), .B2(n_592), .Y(n_737) );
AOI22xp33_ASAP7_75t_SL g589 ( .A1(n_91), .A2(n_131), .B1(n_590), .B2(n_591), .Y(n_589) );
CKINVDCx5p33_ASAP7_75t_R g1791 ( .A(n_92), .Y(n_1791) );
CKINVDCx5p33_ASAP7_75t_R g1766 ( .A(n_93), .Y(n_1766) );
INVx1_ASAP7_75t_L g1190 ( .A(n_94), .Y(n_1190) );
AOI22xp33_ASAP7_75t_SL g817 ( .A1(n_95), .A2(n_311), .B1(n_645), .B2(n_718), .Y(n_817) );
INVxp67_ASAP7_75t_SL g824 ( .A(n_95), .Y(n_824) );
INVx1_ASAP7_75t_L g1149 ( .A(n_96), .Y(n_1149) );
AOI221xp5_ASAP7_75t_L g1159 ( .A1(n_96), .A2(n_216), .B1(n_472), .B2(n_507), .C(n_653), .Y(n_1159) );
CKINVDCx5p33_ASAP7_75t_R g465 ( .A(n_97), .Y(n_465) );
XNOR2xp5_ASAP7_75t_L g755 ( .A(n_98), .B(n_756), .Y(n_755) );
OAI211xp5_ASAP7_75t_L g1344 ( .A1(n_99), .A2(n_1119), .B(n_1345), .C(n_1347), .Y(n_1344) );
INVx1_ASAP7_75t_L g1376 ( .A(n_99), .Y(n_1376) );
CKINVDCx5p33_ASAP7_75t_R g449 ( .A(n_100), .Y(n_449) );
OAI22xp5_ASAP7_75t_L g509 ( .A1(n_100), .A2(n_116), .B1(n_510), .B2(n_513), .Y(n_509) );
AOI22xp33_ASAP7_75t_L g1462 ( .A1(n_102), .A2(n_224), .B1(n_486), .B2(n_501), .Y(n_1462) );
AOI22xp33_ASAP7_75t_L g1473 ( .A1(n_102), .A2(n_248), .B1(n_406), .B2(n_946), .Y(n_1473) );
INVx1_ASAP7_75t_L g1205 ( .A(n_103), .Y(n_1205) );
CKINVDCx5p33_ASAP7_75t_R g1773 ( .A(n_104), .Y(n_1773) );
AOI21xp33_ASAP7_75t_L g774 ( .A1(n_105), .A2(n_736), .B(n_775), .Y(n_774) );
INVx1_ASAP7_75t_L g783 ( .A(n_105), .Y(n_783) );
INVx1_ASAP7_75t_L g701 ( .A(n_106), .Y(n_701) );
INVx1_ASAP7_75t_L g1447 ( .A(n_107), .Y(n_1447) );
INVx1_ASAP7_75t_L g352 ( .A(n_108), .Y(n_352) );
AOI221xp5_ASAP7_75t_L g760 ( .A1(n_109), .A2(n_246), .B1(n_588), .B2(n_761), .C(n_762), .Y(n_760) );
AOI22xp33_ASAP7_75t_L g785 ( .A1(n_109), .A2(n_172), .B1(n_411), .B2(n_645), .Y(n_785) );
AO221x2_ASAP7_75t_L g1611 ( .A1(n_111), .A2(n_319), .B1(n_1494), .B2(n_1499), .C(n_1612), .Y(n_1611) );
AOI22xp33_ASAP7_75t_L g1724 ( .A1(n_112), .A2(n_178), .B1(n_816), .B2(n_1361), .Y(n_1724) );
INVx1_ASAP7_75t_L g1745 ( .A(n_112), .Y(n_1745) );
INVx1_ASAP7_75t_L g1008 ( .A(n_113), .Y(n_1008) );
OAI22xp33_ASAP7_75t_L g1134 ( .A1(n_114), .A2(n_289), .B1(n_567), .B2(n_1135), .Y(n_1134) );
INVx1_ASAP7_75t_L g1169 ( .A(n_114), .Y(n_1169) );
OAI222xp33_ASAP7_75t_L g1409 ( .A1(n_115), .A2(n_316), .B1(n_965), .B2(n_967), .C1(n_1410), .C2(n_1412), .Y(n_1409) );
INVx1_ASAP7_75t_L g1422 ( .A(n_115), .Y(n_1422) );
CKINVDCx5p33_ASAP7_75t_R g445 ( .A(n_116), .Y(n_445) );
INVx1_ASAP7_75t_L g1400 ( .A(n_117), .Y(n_1400) );
OAI211xp5_ASAP7_75t_L g1449 ( .A1(n_118), .A2(n_837), .B(n_1450), .C(n_1451), .Y(n_1449) );
INVxp33_ASAP7_75t_SL g1466 ( .A(n_118), .Y(n_1466) );
CKINVDCx5p33_ASAP7_75t_R g724 ( .A(n_119), .Y(n_724) );
OAI22xp33_ASAP7_75t_L g972 ( .A1(n_120), .A2(n_164), .B1(n_973), .B2(n_976), .Y(n_972) );
INVxp67_ASAP7_75t_SL g979 ( .A(n_120), .Y(n_979) );
INVx1_ASAP7_75t_L g1141 ( .A(n_121), .Y(n_1141) );
AOI221xp5_ASAP7_75t_L g1162 ( .A1(n_121), .A2(n_271), .B1(n_607), .B2(n_653), .C(n_1163), .Y(n_1162) );
INVxp67_ASAP7_75t_SL g1303 ( .A(n_122), .Y(n_1303) );
AOI22xp33_ASAP7_75t_L g1321 ( .A1(n_122), .A2(n_250), .B1(n_813), .B2(n_1322), .Y(n_1321) );
INVx1_ASAP7_75t_L g872 ( .A(n_123), .Y(n_872) );
INVx1_ASAP7_75t_L g676 ( .A(n_124), .Y(n_676) );
INVx1_ASAP7_75t_L g711 ( .A(n_125), .Y(n_711) );
AOI21xp33_ASAP7_75t_L g747 ( .A1(n_125), .A2(n_507), .B(n_736), .Y(n_747) );
OAI22xp33_ASAP7_75t_SL g1797 ( .A1(n_126), .A2(n_130), .B1(n_1798), .B2(n_1799), .Y(n_1797) );
OAI22xp5_ASAP7_75t_L g1807 ( .A1(n_126), .A2(n_133), .B1(n_447), .B2(n_448), .Y(n_1807) );
OAI22xp5_ASAP7_75t_L g702 ( .A1(n_127), .A2(n_163), .B1(n_703), .B2(n_704), .Y(n_702) );
OAI211xp5_ASAP7_75t_L g733 ( .A1(n_127), .A2(n_650), .B(n_734), .C(n_738), .Y(n_733) );
INVx1_ASAP7_75t_L g1294 ( .A(n_128), .Y(n_1294) );
OAI22xp33_ASAP7_75t_L g1326 ( .A1(n_128), .A2(n_170), .B1(n_1055), .B2(n_1135), .Y(n_1326) );
INVx1_ASAP7_75t_L g1717 ( .A(n_129), .Y(n_1717) );
OAI222xp33_ASAP7_75t_L g1741 ( .A1(n_129), .A2(n_198), .B1(n_686), .B2(n_1742), .C1(n_1743), .C2(n_1746), .Y(n_1741) );
AOI22xp33_ASAP7_75t_L g560 ( .A1(n_131), .A2(n_190), .B1(n_389), .B2(n_561), .Y(n_560) );
INVxp67_ASAP7_75t_SL g1298 ( .A(n_132), .Y(n_1298) );
AOI22xp33_ASAP7_75t_SL g1323 ( .A1(n_132), .A2(n_189), .B1(n_1095), .B2(n_1324), .Y(n_1323) );
INVx1_ASAP7_75t_L g1792 ( .A(n_133), .Y(n_1792) );
AOI221xp5_ASAP7_75t_L g873 ( .A1(n_134), .A2(n_253), .B1(n_480), .B2(n_587), .C(n_761), .Y(n_873) );
AOI22xp33_ASAP7_75t_L g884 ( .A1(n_134), .A2(n_256), .B1(n_411), .B2(n_645), .Y(n_884) );
AOI22xp33_ASAP7_75t_SL g635 ( .A1(n_135), .A2(n_218), .B1(n_427), .B2(n_636), .Y(n_635) );
OAI22xp33_ASAP7_75t_L g991 ( .A1(n_136), .A2(n_341), .B1(n_973), .B2(n_976), .Y(n_991) );
INVxp33_ASAP7_75t_SL g1031 ( .A(n_136), .Y(n_1031) );
AO22x1_ASAP7_75t_L g1515 ( .A1(n_137), .A2(n_324), .B1(n_1494), .B2(n_1499), .Y(n_1515) );
INVx1_ASAP7_75t_L g1088 ( .A(n_138), .Y(n_1088) );
OAI221xp5_ASAP7_75t_L g1116 ( .A1(n_138), .A2(n_139), .B1(n_666), .B2(n_687), .C(n_1117), .Y(n_1116) );
INVx1_ASAP7_75t_L g1089 ( .A(n_139), .Y(n_1089) );
CKINVDCx5p33_ASAP7_75t_R g994 ( .A(n_140), .Y(n_994) );
AOI22xp33_ASAP7_75t_SL g1047 ( .A1(n_141), .A2(n_184), .B1(n_645), .B2(n_946), .Y(n_1047) );
INVx1_ASAP7_75t_L g998 ( .A(n_142), .Y(n_998) );
AOI221xp5_ASAP7_75t_L g1015 ( .A1(n_142), .A2(n_236), .B1(n_736), .B2(n_761), .C(n_1016), .Y(n_1015) );
CKINVDCx5p33_ASAP7_75t_R g1770 ( .A(n_143), .Y(n_1770) );
AOI221xp5_ASAP7_75t_L g914 ( .A1(n_144), .A2(n_157), .B1(n_898), .B2(n_915), .C(n_917), .Y(n_914) );
AOI221xp5_ASAP7_75t_L g945 ( .A1(n_144), .A2(n_317), .B1(n_645), .B2(n_820), .C(n_946), .Y(n_945) );
AOI22xp33_ASAP7_75t_L g1048 ( .A1(n_145), .A2(n_305), .B1(n_813), .B2(n_1049), .Y(n_1048) );
AOI22xp33_ASAP7_75t_L g1063 ( .A1(n_145), .A2(n_209), .B1(n_485), .B2(n_1064), .Y(n_1063) );
INVx1_ASAP7_75t_L g858 ( .A(n_146), .Y(n_858) );
INVx1_ASAP7_75t_L g1731 ( .A(n_147), .Y(n_1731) );
CKINVDCx5p33_ASAP7_75t_R g1058 ( .A(n_148), .Y(n_1058) );
OAI221xp5_ASAP7_75t_L g769 ( .A1(n_149), .A2(n_328), .B1(n_666), .B2(n_687), .C(n_770), .Y(n_769) );
OAI22xp33_ASAP7_75t_L g791 ( .A1(n_149), .A2(n_328), .B1(n_628), .B2(n_730), .Y(n_791) );
OAI22xp33_ASAP7_75t_L g1247 ( .A1(n_150), .A2(n_158), .B1(n_1248), .B2(n_1251), .Y(n_1247) );
OAI22xp33_ASAP7_75t_L g1259 ( .A1(n_150), .A2(n_158), .B1(n_1260), .B2(n_1261), .Y(n_1259) );
INVx1_ASAP7_75t_L g693 ( .A(n_151), .Y(n_693) );
AO22x1_ASAP7_75t_L g381 ( .A1(n_152), .A2(n_188), .B1(n_382), .B2(n_389), .Y(n_381) );
NAND2xp5_ASAP7_75t_L g494 ( .A(n_152), .B(n_495), .Y(n_494) );
INVx1_ASAP7_75t_L g1371 ( .A(n_153), .Y(n_1371) );
AOI22xp33_ASAP7_75t_SL g482 ( .A1(n_154), .A2(n_188), .B1(n_483), .B2(n_485), .Y(n_482) );
INVx1_ASAP7_75t_L g1238 ( .A(n_155), .Y(n_1238) );
INVx1_ASAP7_75t_L g1472 ( .A(n_156), .Y(n_1472) );
AO22x1_ASAP7_75t_L g1522 ( .A1(n_159), .A2(n_325), .B1(n_1502), .B2(n_1523), .Y(n_1522) );
CKINVDCx16_ASAP7_75t_R g1613 ( .A(n_160), .Y(n_1613) );
INVx1_ASAP7_75t_L g1199 ( .A(n_161), .Y(n_1199) );
CKINVDCx5p33_ASAP7_75t_R g1453 ( .A(n_162), .Y(n_1453) );
INVxp67_ASAP7_75t_SL g926 ( .A(n_164), .Y(n_926) );
INVx1_ASAP7_75t_L g803 ( .A(n_165), .Y(n_803) );
INVx1_ASAP7_75t_L g1397 ( .A(n_167), .Y(n_1397) );
AOI22xp33_ASAP7_75t_L g1430 ( .A1(n_167), .A2(n_254), .B1(n_765), .B2(n_1341), .Y(n_1430) );
INVx1_ASAP7_75t_L g918 ( .A(n_168), .Y(n_918) );
AOI221xp5_ASAP7_75t_L g1736 ( .A1(n_169), .A2(n_211), .B1(n_655), .B2(n_1737), .C(n_1738), .Y(n_1736) );
INVx1_ASAP7_75t_L g1292 ( .A(n_170), .Y(n_1292) );
CKINVDCx5p33_ASAP7_75t_R g1452 ( .A(n_171), .Y(n_1452) );
AOI22xp33_ASAP7_75t_SL g776 ( .A1(n_172), .A2(n_299), .B1(n_483), .B2(n_486), .Y(n_776) );
OAI211xp5_ASAP7_75t_L g758 ( .A1(n_173), .A2(n_650), .B(n_759), .C(n_766), .Y(n_758) );
OAI22xp5_ASAP7_75t_L g794 ( .A1(n_173), .A2(n_320), .B1(n_703), .B2(n_704), .Y(n_794) );
INVx1_ASAP7_75t_L g1460 ( .A(n_174), .Y(n_1460) );
AOI22xp33_ASAP7_75t_SL g1094 ( .A1(n_175), .A2(n_281), .B1(n_944), .B2(n_1095), .Y(n_1094) );
AOI22xp33_ASAP7_75t_L g1112 ( .A1(n_175), .A2(n_214), .B1(n_592), .B2(n_658), .Y(n_1112) );
OAI211xp5_ASAP7_75t_L g1335 ( .A1(n_176), .A2(n_1336), .B(n_1337), .C(n_1343), .Y(n_1335) );
NOR2xp33_ASAP7_75t_L g1356 ( .A(n_176), .B(n_438), .Y(n_1356) );
XNOR2x2_ASAP7_75t_L g1039 ( .A(n_177), .B(n_1040), .Y(n_1039) );
AOI22xp33_ASAP7_75t_L g1739 ( .A1(n_178), .A2(n_273), .B1(n_1064), .B2(n_1166), .Y(n_1739) );
AOI22xp33_ASAP7_75t_SL g1325 ( .A1(n_179), .A2(n_338), .B1(n_645), .B2(n_810), .Y(n_1325) );
INVx2_ASAP7_75t_L g1497 ( .A(n_180), .Y(n_1497) );
AND2x2_ASAP7_75t_L g1500 ( .A(n_180), .B(n_1498), .Y(n_1500) );
AND2x2_ASAP7_75t_L g1505 ( .A(n_180), .B(n_285), .Y(n_1505) );
AOI22xp33_ASAP7_75t_L g811 ( .A1(n_181), .A2(n_332), .B1(n_812), .B2(n_813), .Y(n_811) );
INVx1_ASAP7_75t_L g840 ( .A(n_181), .Y(n_840) );
INVx1_ASAP7_75t_L g740 ( .A(n_182), .Y(n_740) );
CKINVDCx5p33_ASAP7_75t_R g1772 ( .A(n_183), .Y(n_1772) );
INVxp67_ASAP7_75t_SL g1074 ( .A(n_184), .Y(n_1074) );
OAI22xp5_ASAP7_75t_L g577 ( .A1(n_185), .A2(n_275), .B1(n_438), .B2(n_519), .Y(n_577) );
OAI211xp5_ASAP7_75t_L g579 ( .A1(n_185), .A2(n_580), .B(n_581), .C(n_593), .Y(n_579) );
CKINVDCx5p33_ASAP7_75t_R g457 ( .A(n_186), .Y(n_457) );
OAI22xp33_ASAP7_75t_L g1054 ( .A1(n_187), .A2(n_255), .B1(n_573), .B2(n_1055), .Y(n_1054) );
INVx1_ASAP7_75t_L g1068 ( .A(n_187), .Y(n_1068) );
INVxp67_ASAP7_75t_SL g1304 ( .A(n_189), .Y(n_1304) );
INVx1_ASAP7_75t_L g1437 ( .A(n_191), .Y(n_1437) );
NOR2xp33_ASAP7_75t_L g1306 ( .A(n_192), .B(n_666), .Y(n_1306) );
INVx1_ASAP7_75t_L g1317 ( .A(n_192), .Y(n_1317) );
INVx1_ASAP7_75t_L g1730 ( .A(n_193), .Y(n_1730) );
AOI22xp33_ASAP7_75t_L g1338 ( .A1(n_194), .A2(n_270), .B1(n_501), .B2(n_765), .Y(n_1338) );
AOI22xp33_ASAP7_75t_SL g1363 ( .A1(n_194), .A2(n_283), .B1(n_645), .B2(n_888), .Y(n_1363) );
AOI22xp33_ASAP7_75t_SL g717 ( .A1(n_195), .A2(n_262), .B1(n_645), .B2(n_718), .Y(n_717) );
AOI22xp33_ASAP7_75t_SL g748 ( .A1(n_195), .A2(n_265), .B1(n_483), .B2(n_502), .Y(n_748) );
INVx1_ASAP7_75t_L g852 ( .A(n_196), .Y(n_852) );
INVx1_ASAP7_75t_L g1145 ( .A(n_197), .Y(n_1145) );
INVx1_ASAP7_75t_L g1718 ( .A(n_198), .Y(n_1718) );
INVx1_ASAP7_75t_L g632 ( .A(n_199), .Y(n_632) );
OAI211xp5_ASAP7_75t_L g649 ( .A1(n_199), .A2(n_650), .B(n_651), .C(n_661), .Y(n_649) );
OAI211xp5_ASAP7_75t_L g1234 ( .A1(n_200), .A2(n_1219), .B(n_1235), .C(n_1237), .Y(n_1234) );
INVx1_ASAP7_75t_L g1280 ( .A(n_200), .Y(n_1280) );
CKINVDCx5p33_ASAP7_75t_R g1399 ( .A(n_201), .Y(n_1399) );
CKINVDCx5p33_ASAP7_75t_R g771 ( .A(n_202), .Y(n_771) );
OAI22xp5_ASAP7_75t_L g1107 ( .A1(n_203), .A2(n_337), .B1(n_573), .B2(n_1055), .Y(n_1107) );
INVx1_ASAP7_75t_L g1114 ( .A(n_203), .Y(n_1114) );
CKINVDCx5p33_ASAP7_75t_R g1351 ( .A(n_204), .Y(n_1351) );
INVx2_ASAP7_75t_L g398 ( .A(n_205), .Y(n_398) );
INVx1_ASAP7_75t_L g420 ( .A(n_205), .Y(n_420) );
NAND2xp5_ASAP7_75t_L g530 ( .A(n_205), .B(n_400), .Y(n_530) );
CKINVDCx5p33_ASAP7_75t_R g662 ( .A(n_206), .Y(n_662) );
OAI211xp5_ASAP7_75t_L g1160 ( .A1(n_207), .A2(n_650), .B(n_1161), .C(n_1168), .Y(n_1160) );
INVx1_ASAP7_75t_L g1407 ( .A(n_208), .Y(n_1407) );
NAND2xp33_ASAP7_75t_SL g1431 ( .A(n_208), .B(n_491), .Y(n_1431) );
AOI22xp33_ASAP7_75t_L g815 ( .A1(n_210), .A2(n_301), .B1(n_723), .B2(n_816), .Y(n_815) );
INVx1_ASAP7_75t_L g838 ( .A(n_210), .Y(n_838) );
AOI22xp33_ASAP7_75t_SL g809 ( .A1(n_212), .A2(n_238), .B1(n_645), .B2(n_810), .Y(n_809) );
INVxp67_ASAP7_75t_SL g842 ( .A(n_212), .Y(n_842) );
INVx1_ASAP7_75t_L g1204 ( .A(n_213), .Y(n_1204) );
INVx1_ASAP7_75t_L g671 ( .A(n_215), .Y(n_671) );
INVx1_ASAP7_75t_L g1146 ( .A(n_216), .Y(n_1146) );
OAI22xp5_ASAP7_75t_L g1354 ( .A1(n_217), .A2(n_290), .B1(n_1345), .B2(n_1355), .Y(n_1354) );
INVx1_ASAP7_75t_L g1374 ( .A(n_217), .Y(n_1374) );
INVx1_ASAP7_75t_L g679 ( .A(n_218), .Y(n_679) );
AOI21xp5_ASAP7_75t_L g1408 ( .A1(n_219), .A2(n_820), .B(n_953), .Y(n_1408) );
INVx1_ASAP7_75t_L g1433 ( .A(n_220), .Y(n_1433) );
OAI21xp5_ASAP7_75t_L g846 ( .A1(n_221), .A2(n_703), .B(n_847), .Y(n_846) );
BUFx3_ASAP7_75t_L g388 ( .A(n_222), .Y(n_388) );
AOI221xp5_ASAP7_75t_L g1111 ( .A1(n_223), .A2(n_231), .B1(n_584), .B2(n_588), .C(n_736), .Y(n_1111) );
AOI22xp33_ASAP7_75t_L g1477 ( .A1(n_224), .A2(n_266), .B1(n_946), .B2(n_1478), .Y(n_1477) );
AOI22xp33_ASAP7_75t_L g1534 ( .A1(n_225), .A2(n_229), .B1(n_1494), .B2(n_1499), .Y(n_1534) );
CKINVDCx5p33_ASAP7_75t_R g995 ( .A(n_227), .Y(n_995) );
OAI22xp5_ASAP7_75t_L g1132 ( .A1(n_228), .A2(n_232), .B1(n_628), .B2(n_1133), .Y(n_1132) );
OAI221xp5_ASAP7_75t_L g1157 ( .A1(n_228), .A2(n_232), .B1(n_686), .B2(n_742), .C(n_1158), .Y(n_1157) );
INVx1_ASAP7_75t_L g1390 ( .A(n_230), .Y(n_1390) );
NOR2xp33_ASAP7_75t_L g1392 ( .A(n_230), .B(n_973), .Y(n_1392) );
AOI22xp33_ASAP7_75t_SL g1093 ( .A1(n_231), .A2(n_276), .B1(n_404), .B2(n_946), .Y(n_1093) );
AOI21xp33_ASAP7_75t_L g1461 ( .A1(n_233), .A2(n_736), .B(n_867), .Y(n_1461) );
INVx1_ASAP7_75t_L g1471 ( .A(n_233), .Y(n_1471) );
INVx1_ASAP7_75t_L g1044 ( .A(n_234), .Y(n_1044) );
INVx1_ASAP7_75t_L g1129 ( .A(n_235), .Y(n_1129) );
AOI21xp33_ASAP7_75t_L g1011 ( .A1(n_236), .A2(n_563), .B(n_950), .Y(n_1011) );
XOR2x2_ASAP7_75t_L g1442 ( .A(n_237), .B(n_1443), .Y(n_1442) );
AOI21xp33_ASAP7_75t_L g826 ( .A1(n_238), .A2(n_480), .B(n_827), .Y(n_826) );
NAND2xp5_ASAP7_75t_L g1083 ( .A(n_239), .B(n_1084), .Y(n_1083) );
AOI22xp5_ASAP7_75t_L g1101 ( .A1(n_239), .A2(n_1102), .B1(n_1103), .B2(n_1124), .Y(n_1101) );
INVx1_ASAP7_75t_L g1126 ( .A(n_239), .Y(n_1126) );
OAI22xp33_ASAP7_75t_L g566 ( .A1(n_240), .A2(n_259), .B1(n_567), .B2(n_573), .Y(n_566) );
INVx1_ASAP7_75t_L g594 ( .A(n_240), .Y(n_594) );
AOI22xp33_ASAP7_75t_L g1757 ( .A1(n_242), .A2(n_1758), .B1(n_1760), .B2(n_1811), .Y(n_1757) );
XOR2xp5_ASAP7_75t_L g1761 ( .A(n_242), .B(n_1762), .Y(n_1761) );
BUFx3_ASAP7_75t_L g369 ( .A(n_243), .Y(n_369) );
INVx1_ASAP7_75t_L g461 ( .A(n_243), .Y(n_461) );
CKINVDCx20_ASAP7_75t_R g1615 ( .A(n_244), .Y(n_1615) );
AOI22xp5_ASAP7_75t_L g1517 ( .A1(n_245), .A2(n_261), .B1(n_1494), .B2(n_1499), .Y(n_1517) );
AOI22xp33_ASAP7_75t_L g789 ( .A1(n_246), .A2(n_299), .B1(n_645), .B2(n_790), .Y(n_789) );
NAND2xp5_ASAP7_75t_SL g1456 ( .A(n_248), .B(n_736), .Y(n_1456) );
AOI21xp5_ASAP7_75t_L g1301 ( .A1(n_250), .A2(n_472), .B(n_867), .Y(n_1301) );
CKINVDCx5p33_ASAP7_75t_R g1000 ( .A(n_251), .Y(n_1000) );
INVx1_ASAP7_75t_L g1405 ( .A(n_254), .Y(n_1405) );
INVx1_ASAP7_75t_L g1069 ( .A(n_255), .Y(n_1069) );
CKINVDCx5p33_ASAP7_75t_R g1100 ( .A(n_257), .Y(n_1100) );
INVx1_ASAP7_75t_L g553 ( .A(n_258), .Y(n_553) );
INVx1_ASAP7_75t_L g597 ( .A(n_259), .Y(n_597) );
NOR2xp33_ASAP7_75t_L g1801 ( .A(n_260), .B(n_1229), .Y(n_1801) );
INVx1_ASAP7_75t_L g739 ( .A(n_263), .Y(n_739) );
CKINVDCx5p33_ASAP7_75t_R g1775 ( .A(n_264), .Y(n_1775) );
NAND2xp5_ASAP7_75t_SL g1458 ( .A(n_266), .B(n_1066), .Y(n_1458) );
AOI22xp5_ASAP7_75t_L g1509 ( .A1(n_267), .A2(n_331), .B1(n_1494), .B2(n_1499), .Y(n_1509) );
INVx1_ASAP7_75t_L g982 ( .A(n_268), .Y(n_982) );
AO22x1_ASAP7_75t_L g1514 ( .A1(n_268), .A2(n_274), .B1(n_1502), .B2(n_1511), .Y(n_1514) );
XNOR2x2_ASAP7_75t_L g547 ( .A(n_269), .B(n_548), .Y(n_547) );
AOI22xp33_ASAP7_75t_SL g1359 ( .A1(n_270), .A2(n_343), .B1(n_645), .B2(n_718), .Y(n_1359) );
INVx1_ASAP7_75t_L g1153 ( .A(n_271), .Y(n_1153) );
INVx1_ASAP7_75t_L g386 ( .A(n_272), .Y(n_386) );
INVx1_ASAP7_75t_L g394 ( .A(n_272), .Y(n_394) );
INVx1_ASAP7_75t_L g685 ( .A(n_277), .Y(n_685) );
OAI21xp33_ASAP7_75t_L g1464 ( .A1(n_278), .A2(n_1369), .B(n_1465), .Y(n_1464) );
INVx1_ASAP7_75t_L g807 ( .A(n_279), .Y(n_807) );
INVx1_ASAP7_75t_L g919 ( .A(n_280), .Y(n_919) );
AOI21xp33_ASAP7_75t_L g1120 ( .A1(n_281), .A2(n_507), .B(n_1121), .Y(n_1120) );
CKINVDCx5p33_ASAP7_75t_R g1389 ( .A(n_282), .Y(n_1389) );
AOI221xp5_ASAP7_75t_SL g1342 ( .A1(n_283), .A2(n_343), .B1(n_474), .B2(n_480), .C(n_491), .Y(n_1342) );
INVx1_ASAP7_75t_L g727 ( .A(n_284), .Y(n_727) );
INVx1_ASAP7_75t_L g1498 ( .A(n_285), .Y(n_1498) );
AND2x2_ASAP7_75t_L g1503 ( .A(n_285), .B(n_1497), .Y(n_1503) );
INVx1_ASAP7_75t_L g1243 ( .A(n_286), .Y(n_1243) );
OAI211xp5_ASAP7_75t_L g1273 ( .A1(n_286), .A2(n_1187), .B(n_1274), .C(n_1277), .Y(n_1273) );
OAI211xp5_ASAP7_75t_SL g1296 ( .A1(n_287), .A2(n_1072), .B(n_1297), .C(n_1302), .Y(n_1296) );
INVx1_ASAP7_75t_L g1315 ( .A(n_287), .Y(n_1315) );
INVx1_ASAP7_75t_L g877 ( .A(n_288), .Y(n_877) );
INVx1_ASAP7_75t_L g1170 ( .A(n_289), .Y(n_1170) );
INVx1_ASAP7_75t_L g1366 ( .A(n_290), .Y(n_1366) );
XNOR2xp5_ASAP7_75t_L g983 ( .A(n_291), .B(n_984), .Y(n_983) );
OAI211xp5_ASAP7_75t_L g1061 ( .A1(n_293), .A2(n_580), .B(n_1062), .C(n_1067), .Y(n_1061) );
INVx1_ASAP7_75t_L g1183 ( .A(n_294), .Y(n_1183) );
INVx1_ASAP7_75t_L g876 ( .A(n_295), .Y(n_876) );
INVxp67_ASAP7_75t_SL g1091 ( .A(n_296), .Y(n_1091) );
OAI211xp5_ASAP7_75t_L g1109 ( .A1(n_296), .A2(n_650), .B(n_1110), .C(n_1113), .Y(n_1109) );
CKINVDCx16_ASAP7_75t_R g1411 ( .A(n_297), .Y(n_1411) );
OAI211xp5_ASAP7_75t_SL g1789 ( .A1(n_300), .A2(n_902), .B(n_1790), .C(n_1794), .Y(n_1789) );
OAI211xp5_ASAP7_75t_SL g1803 ( .A1(n_300), .A2(n_1235), .B(n_1804), .C(n_1806), .Y(n_1803) );
AOI22xp5_ASAP7_75t_L g828 ( .A1(n_301), .A2(n_332), .B1(n_592), .B2(n_829), .Y(n_828) );
NAND2xp5_ASAP7_75t_L g609 ( .A(n_302), .B(n_610), .Y(n_609) );
OAI21xp33_ASAP7_75t_L g1728 ( .A1(n_303), .A2(n_519), .B(n_1729), .Y(n_1728) );
INVx1_ASAP7_75t_L g986 ( .A(n_304), .Y(n_986) );
INVx1_ASAP7_75t_L g1006 ( .A(n_306), .Y(n_1006) );
AOI221xp5_ASAP7_75t_L g1305 ( .A1(n_307), .A2(n_338), .B1(n_588), .B2(n_1079), .C(n_1081), .Y(n_1305) );
INVx1_ASAP7_75t_L g1198 ( .A(n_308), .Y(n_1198) );
INVx1_ASAP7_75t_L g1185 ( .A(n_309), .Y(n_1185) );
CKINVDCx5p33_ASAP7_75t_R g546 ( .A(n_310), .Y(n_546) );
INVxp67_ASAP7_75t_SL g844 ( .A(n_311), .Y(n_844) );
BUFx6f_ASAP7_75t_L g365 ( .A(n_313), .Y(n_365) );
INVx1_ASAP7_75t_L g788 ( .A(n_314), .Y(n_788) );
INVx1_ASAP7_75t_L g1310 ( .A(n_315), .Y(n_1310) );
NOR2xp33_ASAP7_75t_R g1424 ( .A(n_316), .B(n_1425), .Y(n_1424) );
INVx1_ASAP7_75t_L g1385 ( .A(n_318), .Y(n_1385) );
INVxp67_ASAP7_75t_SL g933 ( .A(n_321), .Y(n_933) );
OAI221xp5_ASAP7_75t_L g964 ( .A1(n_321), .A2(n_323), .B1(n_965), .B2(n_967), .C(n_969), .Y(n_964) );
INVx1_ASAP7_75t_L g793 ( .A(n_322), .Y(n_793) );
OAI221xp5_ASAP7_75t_L g905 ( .A1(n_323), .A2(n_327), .B1(n_906), .B2(n_911), .C(n_912), .Y(n_905) );
CKINVDCx5p33_ASAP7_75t_R g1769 ( .A(n_326), .Y(n_1769) );
INVx2_ASAP7_75t_L g402 ( .A(n_329), .Y(n_402) );
INVx1_ASAP7_75t_L g419 ( .A(n_329), .Y(n_419) );
INVx1_ASAP7_75t_L g443 ( .A(n_329), .Y(n_443) );
INVx1_ASAP7_75t_L g1018 ( .A(n_333), .Y(n_1018) );
CKINVDCx5p33_ASAP7_75t_R g1172 ( .A(n_334), .Y(n_1172) );
INVxp67_ASAP7_75t_SL g1077 ( .A(n_335), .Y(n_1077) );
OAI22xp33_ASAP7_75t_SL g729 ( .A1(n_336), .A2(n_340), .B1(n_628), .B2(n_730), .Y(n_729) );
OAI221xp5_ASAP7_75t_L g741 ( .A1(n_336), .A2(n_340), .B1(n_687), .B2(n_742), .C(n_743), .Y(n_741) );
INVx1_ASAP7_75t_L g1115 ( .A(n_337), .Y(n_1115) );
XNOR2xp5_ASAP7_75t_L g698 ( .A(n_339), .B(n_699), .Y(n_698) );
INVxp67_ASAP7_75t_SL g989 ( .A(n_341), .Y(n_989) );
INVx1_ASAP7_75t_L g626 ( .A(n_342), .Y(n_626) );
AOI21xp5_ASAP7_75t_L g344 ( .A1(n_345), .A2(n_370), .B(n_1485), .Y(n_344) );
INVx2_ASAP7_75t_SL g345 ( .A(n_346), .Y(n_345) );
INVx1_ASAP7_75t_L g346 ( .A(n_347), .Y(n_346) );
INVx3_ASAP7_75t_L g347 ( .A(n_348), .Y(n_347) );
OR2x2_ASAP7_75t_L g348 ( .A(n_349), .B(n_355), .Y(n_348) );
NOR2xp33_ASAP7_75t_L g1759 ( .A(n_349), .B(n_358), .Y(n_1759) );
INVx1_ASAP7_75t_L g349 ( .A(n_350), .Y(n_349) );
NOR2xp33_ASAP7_75t_L g350 ( .A(n_351), .B(n_353), .Y(n_350) );
NOR2xp33_ASAP7_75t_L g1756 ( .A(n_351), .B(n_354), .Y(n_1756) );
INVx1_ASAP7_75t_L g1812 ( .A(n_351), .Y(n_1812) );
HB1xp67_ASAP7_75t_L g351 ( .A(n_352), .Y(n_351) );
INVx1_ASAP7_75t_L g353 ( .A(n_354), .Y(n_353) );
NOR2xp33_ASAP7_75t_L g1815 ( .A(n_354), .B(n_1812), .Y(n_1815) );
INVx1_ASAP7_75t_L g355 ( .A(n_356), .Y(n_355) );
NAND2xp5_ASAP7_75t_L g356 ( .A(n_357), .B(n_360), .Y(n_356) );
INVx1_ASAP7_75t_L g357 ( .A(n_358), .Y(n_357) );
AND2x4_ASAP7_75t_L g1285 ( .A(n_358), .B(n_1286), .Y(n_1285) );
INVx1_ASAP7_75t_L g358 ( .A(n_359), .Y(n_358) );
AND2x4_ASAP7_75t_L g481 ( .A(n_359), .B(n_369), .Y(n_481) );
AND2x4_ASAP7_75t_L g508 ( .A(n_359), .B(n_368), .Y(n_508) );
INVx1_ASAP7_75t_L g1260 ( .A(n_360), .Y(n_1260) );
AND2x4_ASAP7_75t_SL g1758 ( .A(n_360), .B(n_1759), .Y(n_1758) );
INVx3_ASAP7_75t_L g360 ( .A(n_361), .Y(n_360) );
OR2x6_ASAP7_75t_L g361 ( .A(n_362), .B(n_367), .Y(n_361) );
INVxp67_ASAP7_75t_L g610 ( .A(n_362), .Y(n_610) );
OR2x6_ASAP7_75t_L g1266 ( .A(n_362), .B(n_1263), .Y(n_1266) );
OR2x2_ASAP7_75t_L g1798 ( .A(n_362), .B(n_1263), .Y(n_1798) );
INVx2_ASAP7_75t_L g362 ( .A(n_363), .Y(n_362) );
INVx3_ASAP7_75t_L g681 ( .A(n_363), .Y(n_681) );
BUFx4f_ASAP7_75t_L g1346 ( .A(n_363), .Y(n_1346) );
INVx3_ASAP7_75t_L g363 ( .A(n_364), .Y(n_363) );
OR2x2_ASAP7_75t_L g364 ( .A(n_365), .B(n_366), .Y(n_364) );
INVx2_ASAP7_75t_L g463 ( .A(n_365), .Y(n_463) );
AND2x2_ASAP7_75t_L g468 ( .A(n_365), .B(n_469), .Y(n_468) );
AND2x2_ASAP7_75t_L g479 ( .A(n_365), .B(n_366), .Y(n_479) );
INVx2_ASAP7_75t_L g488 ( .A(n_365), .Y(n_488) );
INVx1_ASAP7_75t_L g523 ( .A(n_365), .Y(n_523) );
NAND2x1_ASAP7_75t_L g670 ( .A(n_365), .B(n_366), .Y(n_670) );
INVx1_ASAP7_75t_L g464 ( .A(n_366), .Y(n_464) );
INVx2_ASAP7_75t_L g469 ( .A(n_366), .Y(n_469) );
AND2x2_ASAP7_75t_L g487 ( .A(n_366), .B(n_488), .Y(n_487) );
BUFx2_ASAP7_75t_L g516 ( .A(n_366), .Y(n_516) );
NAND2xp5_ASAP7_75t_L g604 ( .A(n_366), .B(n_488), .Y(n_604) );
OR2x2_ASAP7_75t_L g675 ( .A(n_366), .B(n_463), .Y(n_675) );
OR2x6_ASAP7_75t_L g1787 ( .A(n_367), .B(n_681), .Y(n_1787) );
INVxp67_ASAP7_75t_L g367 ( .A(n_368), .Y(n_367) );
INVx1_ASAP7_75t_L g1276 ( .A(n_368), .Y(n_1276) );
INVx2_ASAP7_75t_L g368 ( .A(n_369), .Y(n_368) );
BUFx2_ASAP7_75t_L g1272 ( .A(n_369), .Y(n_1272) );
AND2x4_ASAP7_75t_L g1283 ( .A(n_369), .B(n_522), .Y(n_1283) );
OAI22xp33_ASAP7_75t_L g370 ( .A1(n_371), .A2(n_372), .B1(n_1033), .B2(n_1484), .Y(n_370) );
INVx1_ASAP7_75t_L g371 ( .A(n_372), .Y(n_371) );
XNOR2xp5_ASAP7_75t_L g372 ( .A(n_373), .B(n_694), .Y(n_372) );
XNOR2xp5_ASAP7_75t_L g373 ( .A(n_374), .B(n_622), .Y(n_373) );
OAI22x1_ASAP7_75t_L g374 ( .A1(n_375), .A2(n_376), .B1(n_547), .B2(n_621), .Y(n_374) );
INVx2_ASAP7_75t_L g375 ( .A(n_376), .Y(n_375) );
XNOR2x1_ASAP7_75t_L g376 ( .A(n_377), .B(n_378), .Y(n_376) );
AND3x2_ASAP7_75t_L g378 ( .A(n_379), .B(n_454), .C(n_537), .Y(n_378) );
NOR2xp33_ASAP7_75t_SL g379 ( .A(n_380), .B(n_428), .Y(n_379) );
OAI21xp5_ASAP7_75t_SL g380 ( .A1(n_381), .A2(n_395), .B(n_413), .Y(n_380) );
HB1xp67_ASAP7_75t_L g382 ( .A(n_383), .Y(n_382) );
AND2x4_ASAP7_75t_L g536 ( .A(n_383), .B(n_535), .Y(n_536) );
INVx2_ASAP7_75t_SL g782 ( .A(n_383), .Y(n_782) );
INVx2_ASAP7_75t_SL g1148 ( .A(n_383), .Y(n_1148) );
BUFx8_ASAP7_75t_L g383 ( .A(n_384), .Y(n_383) );
INVx2_ASAP7_75t_L g559 ( .A(n_384), .Y(n_559) );
BUFx6f_ASAP7_75t_L g563 ( .A(n_384), .Y(n_563) );
BUFx6f_ASAP7_75t_L g723 ( .A(n_384), .Y(n_723) );
AND2x4_ASAP7_75t_L g384 ( .A(n_385), .B(n_387), .Y(n_384) );
INVxp67_ASAP7_75t_L g385 ( .A(n_386), .Y(n_385) );
INVx1_ASAP7_75t_L g409 ( .A(n_386), .Y(n_409) );
AND2x4_ASAP7_75t_L g407 ( .A(n_387), .B(n_408), .Y(n_407) );
INVx2_ASAP7_75t_L g387 ( .A(n_388), .Y(n_387) );
BUFx6f_ASAP7_75t_L g391 ( .A(n_388), .Y(n_391) );
AND2x4_ASAP7_75t_L g412 ( .A(n_388), .B(n_393), .Y(n_412) );
NAND2xp5_ASAP7_75t_L g543 ( .A(n_388), .B(n_394), .Y(n_543) );
OR2x2_ASAP7_75t_L g570 ( .A(n_388), .B(n_409), .Y(n_570) );
BUFx3_ASAP7_75t_L g389 ( .A(n_390), .Y(n_389) );
BUFx12f_ASAP7_75t_L g427 ( .A(n_390), .Y(n_427) );
INVx5_ASAP7_75t_L g814 ( .A(n_390), .Y(n_814) );
BUFx2_ASAP7_75t_L g944 ( .A(n_390), .Y(n_944) );
AND2x4_ASAP7_75t_L g977 ( .A(n_390), .B(n_975), .Y(n_977) );
BUFx3_ASAP7_75t_L g1324 ( .A(n_390), .Y(n_1324) );
AND2x4_ASAP7_75t_L g390 ( .A(n_391), .B(n_392), .Y(n_390) );
INVx2_ASAP7_75t_L g448 ( .A(n_391), .Y(n_448) );
NAND2x1p5_ASAP7_75t_L g526 ( .A(n_391), .B(n_527), .Y(n_526) );
BUFx2_ASAP7_75t_L g1242 ( .A(n_391), .Y(n_1242) );
INVx1_ASAP7_75t_L g453 ( .A(n_392), .Y(n_453) );
INVx1_ASAP7_75t_L g392 ( .A(n_393), .Y(n_392) );
INVx2_ASAP7_75t_L g393 ( .A(n_394), .Y(n_393) );
INVx1_ASAP7_75t_L g527 ( .A(n_394), .Y(n_527) );
NAND2xp5_ASAP7_75t_L g395 ( .A(n_396), .B(n_403), .Y(n_395) );
AOI33xp33_ASAP7_75t_L g554 ( .A1(n_396), .A2(n_555), .A3(n_556), .B1(n_560), .B2(n_564), .B3(n_565), .Y(n_554) );
AOI33xp33_ASAP7_75t_L g634 ( .A1(n_396), .A2(n_635), .A3(n_637), .B1(n_642), .B2(n_643), .B3(n_646), .Y(n_634) );
AOI33xp33_ASAP7_75t_L g1722 ( .A1(n_396), .A2(n_1723), .A3(n_1724), .B1(n_1725), .B2(n_1726), .B3(n_1727), .Y(n_1722) );
BUFx3_ASAP7_75t_L g396 ( .A(n_397), .Y(n_396) );
AOI33xp33_ASAP7_75t_L g808 ( .A1(n_397), .A2(n_809), .A3(n_811), .B1(n_815), .B2(n_817), .B3(n_818), .Y(n_808) );
AOI33xp33_ASAP7_75t_L g883 ( .A1(n_397), .A2(n_884), .A3(n_885), .B1(n_886), .B2(n_887), .B3(n_889), .Y(n_883) );
AOI33xp33_ASAP7_75t_L g1046 ( .A1(n_397), .A2(n_564), .A3(n_1047), .B1(n_1048), .B2(n_1051), .B3(n_1052), .Y(n_1046) );
AOI33xp33_ASAP7_75t_L g1092 ( .A1(n_397), .A2(n_646), .A3(n_1093), .B1(n_1094), .B2(n_1097), .B3(n_1098), .Y(n_1092) );
AOI33xp33_ASAP7_75t_L g1318 ( .A1(n_397), .A2(n_564), .A3(n_1319), .B1(n_1321), .B2(n_1323), .B3(n_1325), .Y(n_1318) );
AOI33xp33_ASAP7_75t_L g1358 ( .A1(n_397), .A2(n_1359), .A3(n_1360), .B1(n_1362), .B2(n_1363), .B3(n_1364), .Y(n_1358) );
AND3x4_ASAP7_75t_L g397 ( .A(n_398), .B(n_399), .C(n_401), .Y(n_397) );
INVx1_ASAP7_75t_L g434 ( .A(n_398), .Y(n_434) );
NAND2xp33_ASAP7_75t_SL g709 ( .A(n_398), .B(n_400), .Y(n_709) );
HB1xp67_ASAP7_75t_L g1255 ( .A(n_398), .Y(n_1255) );
AND2x2_ASAP7_75t_L g1401 ( .A(n_398), .B(n_399), .Y(n_1401) );
INVx3_ASAP7_75t_L g1241 ( .A(n_399), .Y(n_1241) );
AND2x2_ASAP7_75t_L g1808 ( .A(n_399), .B(n_453), .Y(n_1808) );
BUFx3_ASAP7_75t_L g399 ( .A(n_400), .Y(n_399) );
INVx3_ASAP7_75t_L g417 ( .A(n_400), .Y(n_417) );
INVx2_ASAP7_75t_SL g517 ( .A(n_401), .Y(n_517) );
INVx1_ASAP7_75t_L g620 ( .A(n_401), .Y(n_620) );
OAI31xp33_ASAP7_75t_SL g990 ( .A1(n_401), .A2(n_991), .A3(n_992), .B(n_996), .Y(n_990) );
OAI31xp33_ASAP7_75t_L g1391 ( .A1(n_401), .A2(n_1392), .A3(n_1393), .B(n_1409), .Y(n_1391) );
INVx2_ASAP7_75t_L g401 ( .A(n_402), .Y(n_401) );
BUFx2_ASAP7_75t_L g752 ( .A(n_402), .Y(n_752) );
NAND2xp5_ASAP7_75t_L g908 ( .A(n_402), .B(n_492), .Y(n_908) );
INVx2_ASAP7_75t_L g404 ( .A(n_405), .Y(n_404) );
INVx2_ASAP7_75t_SL g405 ( .A(n_406), .Y(n_405) );
BUFx3_ASAP7_75t_L g406 ( .A(n_407), .Y(n_406) );
NAND2x1p5_ASAP7_75t_L g439 ( .A(n_407), .B(n_433), .Y(n_439) );
INVx8_ASAP7_75t_L g534 ( .A(n_407), .Y(n_534) );
BUFx3_ASAP7_75t_L g953 ( .A(n_407), .Y(n_953) );
AND2x2_ASAP7_75t_L g956 ( .A(n_407), .B(n_957), .Y(n_956) );
HB1xp67_ASAP7_75t_L g1478 ( .A(n_407), .Y(n_1478) );
INVx1_ASAP7_75t_L g408 ( .A(n_409), .Y(n_408) );
BUFx2_ASAP7_75t_L g410 ( .A(n_411), .Y(n_410) );
AND2x4_ASAP7_75t_L g430 ( .A(n_411), .B(n_431), .Y(n_430) );
BUFx2_ASAP7_75t_L g411 ( .A(n_412), .Y(n_411) );
BUFx2_ASAP7_75t_L g424 ( .A(n_412), .Y(n_424) );
INVx2_ASAP7_75t_L g641 ( .A(n_412), .Y(n_641) );
BUFx2_ASAP7_75t_L g718 ( .A(n_412), .Y(n_718) );
BUFx3_ASAP7_75t_L g946 ( .A(n_412), .Y(n_946) );
AND2x2_ASAP7_75t_L g959 ( .A(n_412), .B(n_957), .Y(n_959) );
BUFx2_ASAP7_75t_L g1053 ( .A(n_412), .Y(n_1053) );
AND2x4_ASAP7_75t_L g1236 ( .A(n_412), .B(n_417), .Y(n_1236) );
BUFx2_ASAP7_75t_L g1320 ( .A(n_412), .Y(n_1320) );
NAND3xp33_ASAP7_75t_L g413 ( .A(n_414), .B(n_421), .C(n_425), .Y(n_413) );
INVx1_ASAP7_75t_L g1154 ( .A(n_414), .Y(n_1154) );
BUFx2_ASAP7_75t_L g414 ( .A(n_415), .Y(n_414) );
BUFx2_ASAP7_75t_L g564 ( .A(n_415), .Y(n_564) );
BUFx2_ASAP7_75t_L g646 ( .A(n_415), .Y(n_646) );
BUFx2_ASAP7_75t_L g1726 ( .A(n_415), .Y(n_1726) );
INVx3_ASAP7_75t_L g415 ( .A(n_416), .Y(n_415) );
INVx3_ASAP7_75t_L g720 ( .A(n_416), .Y(n_720) );
NAND3x1_ASAP7_75t_L g416 ( .A(n_417), .B(n_418), .C(n_420), .Y(n_416) );
AND2x4_ASAP7_75t_L g433 ( .A(n_417), .B(n_434), .Y(n_433) );
NAND2x1p5_ASAP7_75t_L g820 ( .A(n_417), .B(n_420), .Y(n_820) );
INVx1_ASAP7_75t_L g1230 ( .A(n_417), .Y(n_1230) );
OR2x6_ASAP7_75t_L g1233 ( .A(n_417), .B(n_715), .Y(n_1233) );
OR2x4_ASAP7_75t_L g1250 ( .A(n_417), .B(n_570), .Y(n_1250) );
INVx1_ASAP7_75t_L g418 ( .A(n_419), .Y(n_418) );
INVx1_ASAP7_75t_L g432 ( .A(n_419), .Y(n_432) );
NAND2xp5_ASAP7_75t_L g929 ( .A(n_419), .B(n_460), .Y(n_929) );
INVx1_ASAP7_75t_L g422 ( .A(n_423), .Y(n_422) );
INVx1_ASAP7_75t_L g423 ( .A(n_424), .Y(n_423) );
BUFx2_ASAP7_75t_L g426 ( .A(n_427), .Y(n_426) );
NAND3xp33_ASAP7_75t_L g428 ( .A(n_429), .B(n_435), .C(n_444), .Y(n_428) );
AND4x1_ASAP7_75t_L g801 ( .A(n_429), .B(n_802), .C(n_806), .D(n_808), .Y(n_801) );
INVx1_ASAP7_75t_L g1056 ( .A(n_429), .Y(n_1056) );
NAND4xp25_ASAP7_75t_SL g1086 ( .A(n_429), .B(n_1087), .C(n_1090), .D(n_1092), .Y(n_1086) );
NAND2xp5_ASAP7_75t_SL g1719 ( .A(n_429), .B(n_1720), .Y(n_1719) );
INVx3_ASAP7_75t_L g429 ( .A(n_430), .Y(n_429) );
HB1xp67_ASAP7_75t_L g574 ( .A(n_430), .Y(n_574) );
INVx3_ASAP7_75t_L g647 ( .A(n_430), .Y(n_647) );
NOR3xp33_ASAP7_75t_L g778 ( .A(n_430), .B(n_779), .C(n_791), .Y(n_778) );
AOI211xp5_ASAP7_75t_L g880 ( .A1(n_430), .A2(n_437), .B(n_872), .C(n_881), .Y(n_880) );
AOI221xp5_ASAP7_75t_L g1365 ( .A1(n_430), .A2(n_731), .B1(n_804), .B2(n_1348), .C(n_1366), .Y(n_1365) );
AND2x2_ASAP7_75t_L g446 ( .A(n_431), .B(n_447), .Y(n_446) );
AND2x4_ASAP7_75t_L g450 ( .A(n_431), .B(n_451), .Y(n_450) );
NAND2x1_ASAP7_75t_L g628 ( .A(n_431), .B(n_447), .Y(n_628) );
AND2x4_ASAP7_75t_SL g731 ( .A(n_431), .B(n_451), .Y(n_731) );
AND2x4_ASAP7_75t_SL g804 ( .A(n_431), .B(n_447), .Y(n_804) );
AND2x2_ASAP7_75t_L g1316 ( .A(n_431), .B(n_447), .Y(n_1316) );
AND2x4_ASAP7_75t_L g431 ( .A(n_432), .B(n_433), .Y(n_431) );
OR2x2_ASAP7_75t_L g544 ( .A(n_432), .B(n_545), .Y(n_544) );
INVx1_ASAP7_75t_L g924 ( .A(n_432), .Y(n_924) );
AND2x6_ASAP7_75t_L g966 ( .A(n_433), .B(n_447), .Y(n_966) );
AND2x2_ASAP7_75t_L g968 ( .A(n_433), .B(n_453), .Y(n_968) );
INVx1_ASAP7_75t_L g971 ( .A(n_433), .Y(n_971) );
NAND2xp5_ASAP7_75t_L g435 ( .A(n_436), .B(n_437), .Y(n_435) );
AOI221xp5_ASAP7_75t_SL g470 ( .A1(n_436), .A2(n_471), .B1(n_482), .B2(n_489), .C(n_490), .Y(n_470) );
INVx3_ASAP7_75t_L g437 ( .A(n_438), .Y(n_437) );
INVx5_ASAP7_75t_L g633 ( .A(n_438), .Y(n_633) );
OR2x6_ASAP7_75t_L g438 ( .A(n_439), .B(n_440), .Y(n_438) );
OR2x2_ASAP7_75t_L g704 ( .A(n_439), .B(n_440), .Y(n_704) );
INVx2_ASAP7_75t_L g963 ( .A(n_439), .Y(n_963) );
INVxp67_ASAP7_75t_L g440 ( .A(n_441), .Y(n_440) );
OR2x2_ASAP7_75t_L g520 ( .A(n_441), .B(n_521), .Y(n_520) );
OR2x2_ASAP7_75t_L g911 ( .A(n_441), .B(n_521), .Y(n_911) );
INVx1_ASAP7_75t_L g939 ( .A(n_441), .Y(n_939) );
INVx1_ASAP7_75t_L g1286 ( .A(n_441), .Y(n_1286) );
BUFx2_ASAP7_75t_L g441 ( .A(n_442), .Y(n_441) );
INVx2_ASAP7_75t_L g529 ( .A(n_442), .Y(n_529) );
INVx1_ASAP7_75t_L g442 ( .A(n_443), .Y(n_442) );
AOI22xp33_ASAP7_75t_L g444 ( .A1(n_445), .A2(n_446), .B1(n_449), .B2(n_450), .Y(n_444) );
AOI22xp33_ASAP7_75t_L g551 ( .A1(n_446), .A2(n_450), .B1(n_552), .B2(n_553), .Y(n_551) );
AO22x1_ASAP7_75t_L g1716 ( .A1(n_446), .A2(n_450), .B1(n_1717), .B2(n_1718), .Y(n_1716) );
INVx3_ASAP7_75t_L g447 ( .A(n_448), .Y(n_447) );
HB1xp67_ASAP7_75t_L g630 ( .A(n_450), .Y(n_630) );
AOI22xp33_ASAP7_75t_L g1043 ( .A1(n_450), .A2(n_627), .B1(n_1044), .B2(n_1045), .Y(n_1043) );
AOI22xp5_ASAP7_75t_L g1087 ( .A1(n_450), .A2(n_627), .B1(n_1088), .B2(n_1089), .Y(n_1087) );
AOI22xp33_ASAP7_75t_L g1314 ( .A1(n_450), .A2(n_1315), .B1(n_1316), .B2(n_1317), .Y(n_1314) );
AOI221x1_ASAP7_75t_L g1467 ( .A1(n_450), .A2(n_627), .B1(n_1447), .B2(n_1452), .C(n_1468), .Y(n_1467) );
INVx2_ASAP7_75t_L g451 ( .A(n_452), .Y(n_451) );
INVx1_ASAP7_75t_L g452 ( .A(n_453), .Y(n_452) );
AOI21xp5_ASAP7_75t_SL g454 ( .A1(n_455), .A2(n_517), .B(n_518), .Y(n_454) );
NAND3xp33_ASAP7_75t_L g455 ( .A(n_456), .B(n_470), .C(n_493), .Y(n_455) );
AOI22xp33_ASAP7_75t_L g456 ( .A1(n_457), .A2(n_458), .B1(n_465), .B2(n_466), .Y(n_456) );
AOI22xp33_ASAP7_75t_L g531 ( .A1(n_457), .A2(n_465), .B1(n_532), .B2(n_536), .Y(n_531) );
AOI22xp33_ASAP7_75t_L g738 ( .A1(n_458), .A2(n_466), .B1(n_739), .B2(n_740), .Y(n_738) );
AOI22xp5_ASAP7_75t_L g830 ( .A1(n_458), .A2(n_466), .B1(n_831), .B2(n_832), .Y(n_830) );
AOI22xp33_ASAP7_75t_L g875 ( .A1(n_458), .A2(n_466), .B1(n_876), .B2(n_877), .Y(n_875) );
AOI22xp33_ASAP7_75t_L g1113 ( .A1(n_458), .A2(n_466), .B1(n_1114), .B2(n_1115), .Y(n_1113) );
AOI22xp33_ASAP7_75t_L g1293 ( .A1(n_458), .A2(n_489), .B1(n_1294), .B2(n_1295), .Y(n_1293) );
BUFx6f_ASAP7_75t_L g458 ( .A(n_459), .Y(n_458) );
INVx1_ASAP7_75t_L g596 ( .A(n_459), .Y(n_596) );
AOI22xp33_ASAP7_75t_L g766 ( .A1(n_459), .A2(n_466), .B1(n_767), .B2(n_768), .Y(n_766) );
AND2x4_ASAP7_75t_L g938 ( .A(n_459), .B(n_939), .Y(n_938) );
AND2x2_ASAP7_75t_L g459 ( .A(n_460), .B(n_462), .Y(n_459) );
AND2x4_ASAP7_75t_L g466 ( .A(n_460), .B(n_467), .Y(n_466) );
AND2x4_ASAP7_75t_L g489 ( .A(n_460), .B(n_486), .Y(n_489) );
AND2x4_ASAP7_75t_SL g512 ( .A(n_460), .B(n_491), .Y(n_512) );
AND2x2_ASAP7_75t_L g870 ( .A(n_460), .B(n_871), .Y(n_870) );
AND2x2_ASAP7_75t_L g981 ( .A(n_460), .B(n_467), .Y(n_981) );
BUFx2_ASAP7_75t_L g1353 ( .A(n_460), .Y(n_1353) );
HB1xp67_ASAP7_75t_L g1263 ( .A(n_461), .Y(n_1263) );
INVx3_ASAP7_75t_L g484 ( .A(n_462), .Y(n_484) );
BUFx6f_ASAP7_75t_L g501 ( .A(n_462), .Y(n_501) );
NAND2xp5_ASAP7_75t_L g545 ( .A(n_462), .B(n_492), .Y(n_545) );
AND2x2_ASAP7_75t_L g462 ( .A(n_463), .B(n_464), .Y(n_462) );
HB1xp67_ASAP7_75t_L g1350 ( .A(n_463), .Y(n_1350) );
INVx1_ASAP7_75t_L g599 ( .A(n_466), .Y(n_599) );
HB1xp67_ASAP7_75t_L g663 ( .A(n_466), .Y(n_663) );
BUFx6f_ASAP7_75t_L g1070 ( .A(n_466), .Y(n_1070) );
AOI22xp33_ASAP7_75t_L g1734 ( .A1(n_466), .A2(n_595), .B1(n_1730), .B2(n_1731), .Y(n_1734) );
INVx2_ASAP7_75t_L g497 ( .A(n_467), .Y(n_497) );
INVx1_ASAP7_75t_L g763 ( .A(n_467), .Y(n_763) );
BUFx6f_ASAP7_75t_L g827 ( .A(n_467), .Y(n_827) );
BUFx6f_ASAP7_75t_L g467 ( .A(n_468), .Y(n_467) );
INVx2_ASAP7_75t_L g475 ( .A(n_468), .Y(n_475) );
BUFx3_ASAP7_75t_L g736 ( .A(n_468), .Y(n_736) );
AND2x4_ASAP7_75t_L g1262 ( .A(n_468), .B(n_1263), .Y(n_1262) );
INVx2_ASAP7_75t_L g472 ( .A(n_473), .Y(n_472) );
INVx2_ASAP7_75t_L g473 ( .A(n_474), .Y(n_473) );
HB1xp67_ASAP7_75t_L g607 ( .A(n_474), .Y(n_607) );
INVx1_ASAP7_75t_L g1080 ( .A(n_474), .Y(n_1080) );
INVx2_ASAP7_75t_L g474 ( .A(n_475), .Y(n_474) );
INVx2_ASAP7_75t_L g654 ( .A(n_475), .Y(n_654) );
INVx2_ASAP7_75t_L g476 ( .A(n_477), .Y(n_476) );
INVx1_ASAP7_75t_L g866 ( .A(n_477), .Y(n_866) );
INVx1_ASAP7_75t_L g1737 ( .A(n_477), .Y(n_1737) );
BUFx2_ASAP7_75t_L g477 ( .A(n_478), .Y(n_477) );
INVx1_ASAP7_75t_L g1796 ( .A(n_478), .Y(n_1796) );
INVx1_ASAP7_75t_L g478 ( .A(n_479), .Y(n_478) );
BUFx6f_ASAP7_75t_L g491 ( .A(n_479), .Y(n_491) );
INVx4_ASAP7_75t_L g480 ( .A(n_481), .Y(n_480) );
INVx4_ASAP7_75t_L g588 ( .A(n_481), .Y(n_588) );
INVx1_ASAP7_75t_SL g655 ( .A(n_481), .Y(n_655) );
AND2x2_ASAP7_75t_SL g904 ( .A(n_481), .B(n_529), .Y(n_904) );
AND2x4_ASAP7_75t_L g1023 ( .A(n_481), .B(n_1024), .Y(n_1023) );
NAND2xp5_ASAP7_75t_L g1202 ( .A(n_481), .B(n_1024), .Y(n_1202) );
NAND4xp25_ASAP7_75t_L g1455 ( .A(n_481), .B(n_1456), .C(n_1457), .D(n_1458), .Y(n_1455) );
INVx2_ASAP7_75t_SL g483 ( .A(n_484), .Y(n_483) );
INVx2_ASAP7_75t_L g590 ( .A(n_484), .Y(n_590) );
INVx1_ASAP7_75t_L g829 ( .A(n_484), .Y(n_829) );
INVx2_ASAP7_75t_L g1064 ( .A(n_484), .Y(n_1064) );
INVx1_ASAP7_75t_L g1165 ( .A(n_484), .Y(n_1165) );
INVx2_ASAP7_75t_L g1341 ( .A(n_484), .Y(n_1341) );
BUFx2_ASAP7_75t_L g485 ( .A(n_486), .Y(n_485) );
INVx1_ASAP7_75t_L g660 ( .A(n_486), .Y(n_660) );
BUFx6f_ASAP7_75t_L g486 ( .A(n_487), .Y(n_486) );
INVx2_ASAP7_75t_L g503 ( .A(n_487), .Y(n_503) );
BUFx3_ASAP7_75t_L g592 ( .A(n_487), .Y(n_592) );
BUFx3_ASAP7_75t_L g765 ( .A(n_487), .Y(n_765) );
INVx3_ASAP7_75t_L g580 ( .A(n_489), .Y(n_580) );
INVx2_ASAP7_75t_SL g650 ( .A(n_489), .Y(n_650) );
NAND2xp5_ASAP7_75t_L g833 ( .A(n_489), .B(n_807), .Y(n_833) );
NAND2xp5_ASAP7_75t_R g1740 ( .A(n_489), .B(n_1721), .Y(n_1740) );
AOI21xp5_ASAP7_75t_L g581 ( .A1(n_490), .A2(n_582), .B(n_589), .Y(n_581) );
AOI21xp5_ASAP7_75t_L g651 ( .A1(n_490), .A2(n_652), .B(n_656), .Y(n_651) );
AOI21xp5_ASAP7_75t_L g734 ( .A1(n_490), .A2(n_735), .B(n_737), .Y(n_734) );
AOI21xp5_ASAP7_75t_L g759 ( .A1(n_490), .A2(n_760), .B(n_764), .Y(n_759) );
INVx1_ASAP7_75t_L g834 ( .A(n_490), .Y(n_834) );
AOI221xp5_ASAP7_75t_L g869 ( .A1(n_490), .A2(n_870), .B1(n_872), .B2(n_873), .C(n_874), .Y(n_869) );
AOI21xp5_ASAP7_75t_L g1062 ( .A1(n_490), .A2(n_1063), .B(n_1065), .Y(n_1062) );
AOI21xp5_ASAP7_75t_L g1110 ( .A1(n_490), .A2(n_1111), .B(n_1112), .Y(n_1110) );
AOI21xp5_ASAP7_75t_L g1161 ( .A1(n_490), .A2(n_1162), .B(n_1164), .Y(n_1161) );
AOI21xp5_ASAP7_75t_L g1291 ( .A1(n_490), .A2(n_1070), .B(n_1292), .Y(n_1291) );
AOI21xp5_ASAP7_75t_L g1735 ( .A1(n_490), .A2(n_1736), .B(n_1739), .Y(n_1735) );
AND2x6_ASAP7_75t_L g490 ( .A(n_491), .B(n_492), .Y(n_490) );
INVx1_ASAP7_75t_L g506 ( .A(n_491), .Y(n_506) );
BUFx6f_ASAP7_75t_L g584 ( .A(n_491), .Y(n_584) );
BUFx3_ASAP7_75t_L g653 ( .A(n_491), .Y(n_653) );
BUFx3_ASAP7_75t_L g761 ( .A(n_491), .Y(n_761) );
BUFx3_ASAP7_75t_L g1066 ( .A(n_491), .Y(n_1066) );
BUFx3_ASAP7_75t_L g1081 ( .A(n_491), .Y(n_1081) );
AND2x2_ASAP7_75t_L g1275 ( .A(n_491), .B(n_1276), .Y(n_1275) );
AND2x2_ASAP7_75t_L g514 ( .A(n_492), .B(n_515), .Y(n_514) );
NAND2xp5_ASAP7_75t_L g521 ( .A(n_492), .B(n_522), .Y(n_521) );
INVx1_ASAP7_75t_L g614 ( .A(n_492), .Y(n_614) );
AOI31xp33_ASAP7_75t_L g493 ( .A1(n_494), .A2(n_498), .A3(n_504), .B(n_509), .Y(n_493) );
BUFx2_ASAP7_75t_L g495 ( .A(n_496), .Y(n_495) );
INVx2_ASAP7_75t_L g496 ( .A(n_497), .Y(n_496) );
INVx2_ASAP7_75t_L g587 ( .A(n_497), .Y(n_587) );
INVx2_ASAP7_75t_SL g499 ( .A(n_500), .Y(n_499) );
INVx3_ASAP7_75t_L g500 ( .A(n_501), .Y(n_500) );
BUFx6f_ASAP7_75t_L g658 ( .A(n_501), .Y(n_658) );
INVx1_ASAP7_75t_L g502 ( .A(n_503), .Y(n_502) );
INVx3_ASAP7_75t_L g871 ( .A(n_503), .Y(n_871) );
INVx1_ASAP7_75t_L g505 ( .A(n_506), .Y(n_505) );
INVx1_ASAP7_75t_L g677 ( .A(n_507), .Y(n_677) );
INVx2_ASAP7_75t_L g507 ( .A(n_508), .Y(n_507) );
INVx2_ASAP7_75t_L g608 ( .A(n_508), .Y(n_608) );
INVx1_ASAP7_75t_L g775 ( .A(n_508), .Y(n_775) );
INVx3_ASAP7_75t_L g867 ( .A(n_508), .Y(n_867) );
OAI221xp5_ASAP7_75t_L g1743 ( .A1(n_508), .A2(n_672), .B1(n_902), .B2(n_1744), .C(n_1745), .Y(n_1743) );
INVx1_ASAP7_75t_L g510 ( .A(n_511), .Y(n_510) );
AOI222xp33_ASAP7_75t_L g862 ( .A1(n_511), .A2(n_514), .B1(n_863), .B2(n_864), .C1(n_865), .C2(n_868), .Y(n_862) );
NAND2xp5_ASAP7_75t_L g1446 ( .A(n_511), .B(n_1447), .Y(n_1446) );
BUFx3_ASAP7_75t_L g511 ( .A(n_512), .Y(n_511) );
INVx2_ASAP7_75t_L g616 ( .A(n_512), .Y(n_616) );
INVx1_ASAP7_75t_L g513 ( .A(n_514), .Y(n_513) );
AOI22xp5_ASAP7_75t_L g1347 ( .A1(n_515), .A2(n_1348), .B1(n_1349), .B2(n_1351), .Y(n_1347) );
AOI22xp33_ASAP7_75t_L g1451 ( .A1(n_515), .A2(n_1349), .B1(n_1452), .B2(n_1453), .Y(n_1451) );
BUFx2_ASAP7_75t_L g515 ( .A(n_516), .Y(n_515) );
INVx1_ASAP7_75t_L g613 ( .A(n_516), .Y(n_613) );
INVx1_ASAP7_75t_L g910 ( .A(n_516), .Y(n_910) );
AND2x4_ASAP7_75t_L g1279 ( .A(n_516), .B(n_1272), .Y(n_1279) );
O2A1O1Ixp5_ASAP7_75t_L g648 ( .A1(n_517), .A2(n_649), .B(n_665), .C(n_688), .Y(n_648) );
OAI21xp5_ASAP7_75t_L g1060 ( .A1(n_517), .A2(n_1061), .B(n_1071), .Y(n_1060) );
HB1xp67_ASAP7_75t_L g689 ( .A(n_519), .Y(n_689) );
INVx2_ASAP7_75t_L g1105 ( .A(n_519), .Y(n_1105) );
AND2x4_ASAP7_75t_L g519 ( .A(n_520), .B(n_524), .Y(n_519) );
AND2x4_ASAP7_75t_L g703 ( .A(n_520), .B(n_524), .Y(n_703) );
INVx2_ASAP7_75t_SL g1029 ( .A(n_520), .Y(n_1029) );
INVx1_ASAP7_75t_L g522 ( .A(n_523), .Y(n_522) );
INVx2_ASAP7_75t_L g1373 ( .A(n_524), .Y(n_1373) );
OR2x2_ASAP7_75t_L g524 ( .A(n_525), .B(n_528), .Y(n_524) );
INVx3_ASAP7_75t_L g1010 ( .A(n_525), .Y(n_1010) );
BUFx6f_ASAP7_75t_L g1213 ( .A(n_525), .Y(n_1213) );
BUFx6f_ASAP7_75t_L g525 ( .A(n_526), .Y(n_525) );
BUFx2_ASAP7_75t_L g970 ( .A(n_526), .Y(n_970) );
BUFx3_ASAP7_75t_L g1220 ( .A(n_526), .Y(n_1220) );
BUFx2_ASAP7_75t_L g1246 ( .A(n_527), .Y(n_1246) );
INVx1_ASAP7_75t_L g535 ( .A(n_528), .Y(n_535) );
OR2x2_ASAP7_75t_L g540 ( .A(n_528), .B(n_541), .Y(n_540) );
INVx1_ASAP7_75t_L g572 ( .A(n_528), .Y(n_572) );
OR2x2_ASAP7_75t_L g528 ( .A(n_529), .B(n_530), .Y(n_528) );
OR2x2_ASAP7_75t_L g708 ( .A(n_529), .B(n_709), .Y(n_708) );
INVx1_ASAP7_75t_L g1025 ( .A(n_529), .Y(n_1025) );
HB1xp67_ASAP7_75t_L g1257 ( .A(n_529), .Y(n_1257) );
INVx1_ASAP7_75t_L g957 ( .A(n_530), .Y(n_957) );
INVx1_ASAP7_75t_L g975 ( .A(n_530), .Y(n_975) );
AOI22xp33_ASAP7_75t_L g690 ( .A1(n_532), .A2(n_536), .B1(n_662), .B2(n_664), .Y(n_690) );
AOI22xp33_ASAP7_75t_L g753 ( .A1(n_532), .A2(n_536), .B1(n_739), .B2(n_740), .Y(n_753) );
AOI22xp33_ASAP7_75t_L g795 ( .A1(n_532), .A2(n_536), .B1(n_767), .B2(n_768), .Y(n_795) );
AOI22xp33_ASAP7_75t_L g879 ( .A1(n_532), .A2(n_849), .B1(n_876), .B2(n_877), .Y(n_879) );
AOI22xp33_ASAP7_75t_L g1729 ( .A1(n_532), .A2(n_536), .B1(n_1730), .B2(n_1731), .Y(n_1729) );
AND2x4_ASAP7_75t_L g532 ( .A(n_533), .B(n_535), .Y(n_532) );
AND2x4_ASAP7_75t_L g848 ( .A(n_533), .B(n_535), .Y(n_848) );
AOI22xp5_ASAP7_75t_L g1410 ( .A1(n_533), .A2(n_888), .B1(n_1389), .B2(n_1411), .Y(n_1410) );
INVx2_ASAP7_75t_L g533 ( .A(n_534), .Y(n_533) );
INVx3_ASAP7_75t_L g636 ( .A(n_534), .Y(n_636) );
INVx8_ASAP7_75t_L g645 ( .A(n_534), .Y(n_645) );
CKINVDCx5p33_ASAP7_75t_R g1002 ( .A(n_534), .Y(n_1002) );
INVx2_ASAP7_75t_L g573 ( .A(n_536), .Y(n_573) );
INVx2_ASAP7_75t_L g1135 ( .A(n_536), .Y(n_1135) );
NAND2xp5_ASAP7_75t_L g537 ( .A(n_538), .B(n_546), .Y(n_537) );
AOI21xp5_ASAP7_75t_L g575 ( .A1(n_538), .A2(n_576), .B(n_577), .Y(n_575) );
NAND2xp5_ASAP7_75t_L g691 ( .A(n_538), .B(n_692), .Y(n_691) );
AOI21xp5_ASAP7_75t_L g700 ( .A1(n_538), .A2(n_701), .B(n_702), .Y(n_700) );
AOI21xp5_ASAP7_75t_L g792 ( .A1(n_538), .A2(n_793), .B(n_794), .Y(n_792) );
NAND2xp5_ASAP7_75t_L g851 ( .A(n_538), .B(n_852), .Y(n_851) );
NAND2xp5_ASAP7_75t_L g857 ( .A(n_538), .B(n_858), .Y(n_857) );
AOI21xp33_ASAP7_75t_SL g1057 ( .A1(n_538), .A2(n_1058), .B(n_1059), .Y(n_1057) );
NAND2xp33_ASAP7_75t_L g1099 ( .A(n_538), .B(n_1100), .Y(n_1099) );
AOI21xp33_ASAP7_75t_L g1171 ( .A1(n_538), .A2(n_1172), .B(n_1173), .Y(n_1171) );
AOI21xp33_ASAP7_75t_SL g1309 ( .A1(n_538), .A2(n_1310), .B(n_1311), .Y(n_1309) );
AOI211x1_ASAP7_75t_L g1712 ( .A1(n_538), .A2(n_1713), .B(n_1714), .C(n_1728), .Y(n_1712) );
INVx8_ASAP7_75t_L g538 ( .A(n_539), .Y(n_538) );
AND2x4_ASAP7_75t_L g539 ( .A(n_540), .B(n_544), .Y(n_539) );
INVx1_ASAP7_75t_L g1375 ( .A(n_540), .Y(n_1375) );
BUFx3_ASAP7_75t_L g999 ( .A(n_541), .Y(n_999) );
INVx1_ASAP7_75t_L g541 ( .A(n_542), .Y(n_541) );
BUFx6f_ASAP7_75t_L g726 ( .A(n_542), .Y(n_726) );
INVx1_ASAP7_75t_L g542 ( .A(n_543), .Y(n_542) );
BUFx2_ASAP7_75t_L g715 ( .A(n_543), .Y(n_715) );
NAND2xp5_ASAP7_75t_L g1438 ( .A(n_544), .B(n_1439), .Y(n_1438) );
INVx1_ASAP7_75t_L g925 ( .A(n_545), .Y(n_925) );
INVx1_ASAP7_75t_L g621 ( .A(n_547), .Y(n_621) );
NAND3xp33_ASAP7_75t_L g548 ( .A(n_549), .B(n_575), .C(n_578), .Y(n_548) );
NOR3xp33_ASAP7_75t_L g549 ( .A(n_550), .B(n_566), .C(n_574), .Y(n_549) );
NAND2xp5_ASAP7_75t_L g550 ( .A(n_551), .B(n_554), .Y(n_550) );
AOI22xp33_ASAP7_75t_L g611 ( .A1(n_552), .A2(n_553), .B1(n_612), .B2(n_615), .Y(n_611) );
INVx2_ASAP7_75t_L g557 ( .A(n_558), .Y(n_557) );
BUFx2_ASAP7_75t_L g558 ( .A(n_559), .Y(n_558) );
OAI221xp5_ASAP7_75t_L g710 ( .A1(n_559), .A2(n_711), .B1(n_712), .B2(n_716), .C(n_717), .Y(n_710) );
INVx3_ASAP7_75t_L g850 ( .A(n_559), .Y(n_850) );
INVx1_ASAP7_75t_L g943 ( .A(n_559), .Y(n_943) );
OR2x6_ASAP7_75t_SL g973 ( .A(n_559), .B(n_974), .Y(n_973) );
INVx8_ASAP7_75t_L g561 ( .A(n_562), .Y(n_561) );
BUFx3_ASAP7_75t_L g639 ( .A(n_562), .Y(n_639) );
OAI221xp5_ASAP7_75t_L g1475 ( .A1(n_562), .A2(n_999), .B1(n_1460), .B2(n_1476), .C(n_1477), .Y(n_1475) );
INVx5_ASAP7_75t_L g562 ( .A(n_563), .Y(n_562) );
INVx3_ASAP7_75t_L g949 ( .A(n_563), .Y(n_949) );
INVx2_ASAP7_75t_SL g1096 ( .A(n_563), .Y(n_1096) );
HB1xp67_ASAP7_75t_L g1322 ( .A(n_563), .Y(n_1322) );
INVx2_ASAP7_75t_SL g1403 ( .A(n_563), .Y(n_1403) );
NAND2xp5_ASAP7_75t_L g1481 ( .A(n_567), .B(n_937), .Y(n_1481) );
OR2x6_ASAP7_75t_L g567 ( .A(n_568), .B(n_571), .Y(n_567) );
OR2x2_ASAP7_75t_L g1055 ( .A(n_568), .B(n_571), .Y(n_1055) );
INVx2_ASAP7_75t_SL g1144 ( .A(n_568), .Y(n_1144) );
INVx2_ASAP7_75t_SL g568 ( .A(n_569), .Y(n_568) );
INVx2_ASAP7_75t_L g569 ( .A(n_570), .Y(n_569) );
BUFx4f_ASAP7_75t_L g1210 ( .A(n_570), .Y(n_1210) );
OR2x4_ASAP7_75t_L g1229 ( .A(n_570), .B(n_1230), .Y(n_1229) );
INVxp67_ASAP7_75t_L g571 ( .A(n_572), .Y(n_571) );
AND2x2_ASAP7_75t_L g849 ( .A(n_572), .B(n_850), .Y(n_849) );
NOR3xp33_ASAP7_75t_L g705 ( .A(n_574), .B(n_706), .C(n_729), .Y(n_705) );
OAI21xp5_ASAP7_75t_L g578 ( .A1(n_579), .A2(n_600), .B(n_617), .Y(n_578) );
BUFx2_ASAP7_75t_L g583 ( .A(n_584), .Y(n_583) );
INVx1_ASAP7_75t_L g585 ( .A(n_586), .Y(n_585) );
INVx1_ASAP7_75t_L g586 ( .A(n_587), .Y(n_586) );
HB1xp67_ASAP7_75t_SL g1163 ( .A(n_588), .Y(n_1163) );
BUFx3_ASAP7_75t_L g591 ( .A(n_592), .Y(n_591) );
INVx1_ASAP7_75t_SL g1167 ( .A(n_592), .Y(n_1167) );
AOI22xp33_ASAP7_75t_L g593 ( .A1(n_594), .A2(n_595), .B1(n_597), .B2(n_598), .Y(n_593) );
AOI22xp33_ASAP7_75t_L g661 ( .A1(n_595), .A2(n_662), .B1(n_663), .B2(n_664), .Y(n_661) );
AOI22xp5_ASAP7_75t_L g1067 ( .A1(n_595), .A2(n_1068), .B1(n_1069), .B2(n_1070), .Y(n_1067) );
AOI22xp33_ASAP7_75t_L g1168 ( .A1(n_595), .A2(n_663), .B1(n_1169), .B2(n_1170), .Y(n_1168) );
INVx2_ASAP7_75t_L g595 ( .A(n_596), .Y(n_595) );
INVx1_ASAP7_75t_L g598 ( .A(n_599), .Y(n_598) );
INVx5_ASAP7_75t_L g1751 ( .A(n_601), .Y(n_1751) );
BUFx6f_ASAP7_75t_L g601 ( .A(n_602), .Y(n_601) );
INVx2_ASAP7_75t_L g684 ( .A(n_602), .Y(n_684) );
INVx2_ASAP7_75t_L g845 ( .A(n_602), .Y(n_845) );
INVx2_ASAP7_75t_SL g1076 ( .A(n_602), .Y(n_1076) );
INVx4_ASAP7_75t_L g1196 ( .A(n_602), .Y(n_1196) );
INVx8_ASAP7_75t_L g602 ( .A(n_603), .Y(n_602) );
BUFx2_ASAP7_75t_L g916 ( .A(n_603), .Y(n_916) );
OR2x2_ASAP7_75t_L g1271 ( .A(n_603), .B(n_1272), .Y(n_1271) );
OR2x2_ASAP7_75t_L g1788 ( .A(n_603), .B(n_1276), .Y(n_1788) );
BUFx6f_ASAP7_75t_L g603 ( .A(n_604), .Y(n_603) );
NAND2xp5_ASAP7_75t_L g605 ( .A(n_606), .B(n_609), .Y(n_605) );
INVx1_ASAP7_75t_L g843 ( .A(n_610), .Y(n_843) );
INVx2_ASAP7_75t_L g687 ( .A(n_612), .Y(n_687) );
INVx2_ASAP7_75t_L g1072 ( .A(n_612), .Y(n_1072) );
NOR2x1_ASAP7_75t_L g612 ( .A(n_613), .B(n_614), .Y(n_612) );
INVx1_ASAP7_75t_L g1352 ( .A(n_614), .Y(n_1352) );
INVx2_ASAP7_75t_L g666 ( .A(n_615), .Y(n_666) );
INVx2_ASAP7_75t_L g742 ( .A(n_615), .Y(n_742) );
INVx1_ASAP7_75t_L g1742 ( .A(n_615), .Y(n_1742) );
INVx4_ASAP7_75t_L g615 ( .A(n_616), .Y(n_615) );
OAI21xp5_ASAP7_75t_L g1156 ( .A1(n_617), .A2(n_1157), .B(n_1160), .Y(n_1156) );
INVx2_ASAP7_75t_L g617 ( .A(n_618), .Y(n_617) );
INVx1_ASAP7_75t_L g618 ( .A(n_619), .Y(n_618) );
A2O1A1Ixp33_ASAP7_75t_L g940 ( .A1(n_619), .A2(n_941), .B(n_960), .C(n_978), .Y(n_940) );
INVx1_ASAP7_75t_L g1308 ( .A(n_619), .Y(n_1308) );
HB1xp67_ASAP7_75t_L g1463 ( .A(n_619), .Y(n_1463) );
BUFx2_ASAP7_75t_L g619 ( .A(n_620), .Y(n_619) );
BUFx2_ASAP7_75t_L g777 ( .A(n_620), .Y(n_777) );
AOI21x1_ASAP7_75t_L g1334 ( .A1(n_620), .A2(n_1335), .B(n_1356), .Y(n_1334) );
XOR2x2_ASAP7_75t_L g622 ( .A(n_623), .B(n_693), .Y(n_622) );
NAND3x1_ASAP7_75t_SL g623 ( .A(n_624), .B(n_648), .C(n_691), .Y(n_623) );
AND4x1_ASAP7_75t_L g624 ( .A(n_625), .B(n_631), .C(n_634), .D(n_647), .Y(n_624) );
AOI22xp33_ASAP7_75t_L g625 ( .A1(n_626), .A2(n_627), .B1(n_629), .B2(n_630), .Y(n_625) );
INVx2_ASAP7_75t_L g627 ( .A(n_628), .Y(n_627) );
INVx1_ASAP7_75t_L g1133 ( .A(n_630), .Y(n_1133) );
NAND2xp5_ASAP7_75t_L g631 ( .A(n_632), .B(n_633), .Y(n_631) );
NAND2xp5_ASAP7_75t_L g806 ( .A(n_633), .B(n_807), .Y(n_806) );
NAND2xp5_ASAP7_75t_L g1090 ( .A(n_633), .B(n_1091), .Y(n_1090) );
NAND2xp5_ASAP7_75t_L g1482 ( .A(n_633), .B(n_1483), .Y(n_1482) );
NAND2xp5_ASAP7_75t_L g1720 ( .A(n_633), .B(n_1721), .Y(n_1720) );
INVx1_ASAP7_75t_L g638 ( .A(n_639), .Y(n_638) );
OAI22xp5_ASAP7_75t_L g1142 ( .A1(n_639), .A2(n_1143), .B1(n_1145), .B2(n_1146), .Y(n_1142) );
INVx1_ASAP7_75t_L g640 ( .A(n_641), .Y(n_640) );
INVx2_ASAP7_75t_L g790 ( .A(n_641), .Y(n_790) );
INVx1_ASAP7_75t_L g810 ( .A(n_641), .Y(n_810) );
INVx2_ASAP7_75t_L g888 ( .A(n_641), .Y(n_888) );
BUFx2_ASAP7_75t_L g644 ( .A(n_645), .Y(n_644) );
INVx2_ASAP7_75t_SL g1155 ( .A(n_647), .Y(n_1155) );
AND5x1_ASAP7_75t_L g1443 ( .A(n_647), .B(n_1444), .C(n_1467), .D(n_1479), .E(n_1482), .Y(n_1443) );
HB1xp67_ASAP7_75t_L g657 ( .A(n_658), .Y(n_657) );
INVx1_ASAP7_75t_L g659 ( .A(n_660), .Y(n_659) );
OAI221xp5_ASAP7_75t_L g667 ( .A1(n_668), .A2(n_671), .B1(n_672), .B2(n_676), .C(n_677), .Y(n_667) );
BUFx2_ASAP7_75t_SL g668 ( .A(n_669), .Y(n_668) );
INVx2_ASAP7_75t_SL g773 ( .A(n_669), .Y(n_773) );
OR2x2_ASAP7_75t_L g932 ( .A(n_669), .B(n_929), .Y(n_932) );
OR2x2_ASAP7_75t_L g1425 ( .A(n_669), .B(n_929), .Y(n_1425) );
BUFx3_ASAP7_75t_L g669 ( .A(n_670), .Y(n_669) );
BUFx6f_ASAP7_75t_L g746 ( .A(n_670), .Y(n_746) );
INVx2_ASAP7_75t_L g672 ( .A(n_673), .Y(n_672) );
INVx4_ASAP7_75t_L g673 ( .A(n_674), .Y(n_673) );
BUFx2_ASAP7_75t_L g674 ( .A(n_675), .Y(n_674) );
BUFx3_ASAP7_75t_L g839 ( .A(n_675), .Y(n_839) );
BUFx2_ASAP7_75t_L g1184 ( .A(n_675), .Y(n_1184) );
INVx1_ASAP7_75t_L g1429 ( .A(n_675), .Y(n_1429) );
OAI221xp5_ASAP7_75t_L g836 ( .A1(n_677), .A2(n_837), .B1(n_838), .B2(n_839), .C(n_840), .Y(n_836) );
OAI22xp5_ASAP7_75t_L g678 ( .A1(n_679), .A2(n_680), .B1(n_682), .B2(n_685), .Y(n_678) );
INVx1_ASAP7_75t_L g898 ( .A(n_680), .Y(n_898) );
OAI221xp5_ASAP7_75t_L g1073 ( .A1(n_680), .A2(n_1074), .B1(n_1075), .B2(n_1077), .C(n_1078), .Y(n_1073) );
OAI221xp5_ASAP7_75t_SL g1158 ( .A1(n_680), .A2(n_682), .B1(n_1145), .B2(n_1152), .C(n_1159), .Y(n_1158) );
OAI221xp5_ASAP7_75t_L g1302 ( .A1(n_680), .A2(n_1075), .B1(n_1303), .B2(n_1304), .C(n_1305), .Y(n_1302) );
BUFx6f_ASAP7_75t_L g680 ( .A(n_681), .Y(n_680) );
OAI22xp5_ASAP7_75t_L g1016 ( .A1(n_681), .A2(n_845), .B1(n_1017), .B2(n_1018), .Y(n_1016) );
OAI22x1_ASAP7_75t_SL g1021 ( .A1(n_681), .A2(n_845), .B1(n_1000), .B2(n_1022), .Y(n_1021) );
INVx2_ASAP7_75t_SL g1192 ( .A(n_681), .Y(n_1192) );
BUFx3_ASAP7_75t_L g1781 ( .A(n_681), .Y(n_1781) );
BUFx2_ASAP7_75t_L g682 ( .A(n_683), .Y(n_682) );
INVx1_ASAP7_75t_L g897 ( .A(n_683), .Y(n_897) );
OAI22xp5_ASAP7_75t_L g1780 ( .A1(n_683), .A2(n_1766), .B1(n_1775), .B2(n_1781), .Y(n_1780) );
BUFx6f_ASAP7_75t_L g683 ( .A(n_684), .Y(n_683) );
BUFx2_ASAP7_75t_L g686 ( .A(n_687), .Y(n_686) );
HB1xp67_ASAP7_75t_L g694 ( .A(n_695), .Y(n_694) );
XNOR2x1_ASAP7_75t_L g695 ( .A(n_696), .B(n_797), .Y(n_695) );
INVx1_ASAP7_75t_L g696 ( .A(n_697), .Y(n_696) );
AO22x2_ASAP7_75t_L g697 ( .A1(n_698), .A2(n_754), .B1(n_755), .B2(n_796), .Y(n_697) );
INVx1_ASAP7_75t_L g796 ( .A(n_698), .Y(n_796) );
AND4x1_ASAP7_75t_L g699 ( .A(n_700), .B(n_705), .C(n_732), .D(n_753), .Y(n_699) );
NAND2xp5_ASAP7_75t_L g1434 ( .A(n_704), .B(n_1435), .Y(n_1434) );
OAI22xp5_ASAP7_75t_SL g706 ( .A1(n_707), .A2(n_710), .B1(n_719), .B2(n_721), .Y(n_706) );
BUFx3_ASAP7_75t_L g1207 ( .A(n_707), .Y(n_1207) );
OAI33xp33_ASAP7_75t_L g1764 ( .A1(n_707), .A2(n_1765), .A3(n_1768), .B1(n_1771), .B2(n_1774), .B3(n_1777), .Y(n_1764) );
BUFx4f_ASAP7_75t_L g707 ( .A(n_708), .Y(n_707) );
BUFx8_ASAP7_75t_L g780 ( .A(n_708), .Y(n_780) );
BUFx2_ASAP7_75t_L g1469 ( .A(n_708), .Y(n_1469) );
BUFx2_ASAP7_75t_L g950 ( .A(n_709), .Y(n_950) );
OAI221xp5_ASAP7_75t_L g781 ( .A1(n_712), .A2(n_782), .B1(n_783), .B2(n_784), .C(n_785), .Y(n_781) );
INVx3_ASAP7_75t_L g712 ( .A(n_713), .Y(n_712) );
BUFx2_ASAP7_75t_L g713 ( .A(n_714), .Y(n_713) );
INVx1_ASAP7_75t_L g714 ( .A(n_715), .Y(n_714) );
INVx2_ASAP7_75t_L g719 ( .A(n_720), .Y(n_719) );
CKINVDCx5p33_ASAP7_75t_R g786 ( .A(n_720), .Y(n_786) );
INVx2_ASAP7_75t_L g1474 ( .A(n_720), .Y(n_1474) );
OAI221xp5_ASAP7_75t_L g721 ( .A1(n_722), .A2(n_724), .B1(n_725), .B2(n_727), .C(n_728), .Y(n_721) );
INVx1_ASAP7_75t_L g812 ( .A(n_722), .Y(n_812) );
INVx2_ASAP7_75t_L g722 ( .A(n_723), .Y(n_722) );
INVx2_ASAP7_75t_L g1050 ( .A(n_723), .Y(n_1050) );
INVx2_ASAP7_75t_L g1215 ( .A(n_723), .Y(n_1215) );
BUFx6f_ASAP7_75t_L g1218 ( .A(n_723), .Y(n_1218) );
AND2x4_ASAP7_75t_L g1252 ( .A(n_723), .B(n_1230), .Y(n_1252) );
BUFx6f_ASAP7_75t_L g1361 ( .A(n_723), .Y(n_1361) );
OAI211xp5_ASAP7_75t_L g743 ( .A1(n_724), .A2(n_744), .B(n_747), .C(n_748), .Y(n_743) );
OAI221xp5_ASAP7_75t_L g787 ( .A1(n_725), .A2(n_771), .B1(n_782), .B2(n_788), .C(n_789), .Y(n_787) );
CKINVDCx8_ASAP7_75t_R g725 ( .A(n_726), .Y(n_725) );
INVx3_ASAP7_75t_L g1138 ( .A(n_726), .Y(n_1138) );
INVx3_ASAP7_75t_L g1224 ( .A(n_726), .Y(n_1224) );
INVx3_ASAP7_75t_L g1396 ( .A(n_726), .Y(n_1396) );
INVx1_ASAP7_75t_L g730 ( .A(n_731), .Y(n_730) );
AOI22xp5_ASAP7_75t_L g802 ( .A1(n_731), .A2(n_803), .B1(n_804), .B2(n_805), .Y(n_802) );
AOI22xp33_ASAP7_75t_L g882 ( .A1(n_731), .A2(n_804), .B1(n_863), .B2(n_864), .Y(n_882) );
OAI21xp5_ASAP7_75t_L g732 ( .A1(n_733), .A2(n_741), .B(n_749), .Y(n_732) );
INVx1_ASAP7_75t_L g1122 ( .A(n_736), .Y(n_1122) );
INVx1_ASAP7_75t_L g744 ( .A(n_745), .Y(n_744) );
INVx2_ASAP7_75t_L g837 ( .A(n_745), .Y(n_837) );
INVx2_ASAP7_75t_L g1119 ( .A(n_745), .Y(n_1119) );
INVx4_ASAP7_75t_L g745 ( .A(n_746), .Y(n_745) );
BUFx4f_ASAP7_75t_L g825 ( .A(n_746), .Y(n_825) );
BUFx4f_ASAP7_75t_L g902 ( .A(n_746), .Y(n_902) );
OR2x6_ASAP7_75t_L g912 ( .A(n_746), .B(n_913), .Y(n_912) );
BUFx6f_ASAP7_75t_L g1187 ( .A(n_746), .Y(n_1187) );
BUFx4f_ASAP7_75t_L g1299 ( .A(n_746), .Y(n_1299) );
BUFx4f_ASAP7_75t_L g1355 ( .A(n_746), .Y(n_1355) );
OAI21xp5_ASAP7_75t_L g1108 ( .A1(n_749), .A2(n_1109), .B(n_1116), .Y(n_1108) );
OAI21xp5_ASAP7_75t_L g1732 ( .A1(n_749), .A2(n_1733), .B(n_1741), .Y(n_1732) );
INVx2_ASAP7_75t_L g749 ( .A(n_750), .Y(n_749) );
INVx1_ASAP7_75t_L g860 ( .A(n_750), .Y(n_860) );
BUFx2_ASAP7_75t_L g750 ( .A(n_751), .Y(n_750) );
NAND2xp5_ASAP7_75t_L g1439 ( .A(n_751), .B(n_977), .Y(n_1439) );
INVx1_ASAP7_75t_L g751 ( .A(n_752), .Y(n_751) );
OR2x6_ASAP7_75t_L g819 ( .A(n_752), .B(n_820), .Y(n_819) );
AND2x4_ASAP7_75t_L g920 ( .A(n_752), .B(n_921), .Y(n_920) );
OR2x2_ASAP7_75t_L g1777 ( .A(n_752), .B(n_820), .Y(n_1777) );
INVx1_ASAP7_75t_L g754 ( .A(n_755), .Y(n_754) );
AND4x1_ASAP7_75t_L g756 ( .A(n_757), .B(n_778), .C(n_792), .D(n_795), .Y(n_756) );
OAI21xp5_ASAP7_75t_L g757 ( .A1(n_758), .A2(n_769), .B(n_777), .Y(n_757) );
INVx2_ASAP7_75t_SL g762 ( .A(n_763), .Y(n_762) );
OAI211xp5_ASAP7_75t_L g770 ( .A1(n_771), .A2(n_772), .B(n_774), .C(n_776), .Y(n_770) );
OAI211xp5_ASAP7_75t_L g1459 ( .A1(n_772), .A2(n_1460), .B(n_1461), .C(n_1462), .Y(n_1459) );
INVx5_ASAP7_75t_L g772 ( .A(n_773), .Y(n_772) );
O2A1O1Ixp5_ASAP7_75t_SL g821 ( .A1(n_777), .A2(n_822), .B(n_835), .C(n_846), .Y(n_821) );
OAI22xp5_ASAP7_75t_SL g779 ( .A1(n_780), .A2(n_781), .B1(n_786), .B2(n_787), .Y(n_779) );
OAI33xp33_ASAP7_75t_L g1136 ( .A1(n_780), .A2(n_1137), .A3(n_1142), .B1(n_1147), .B2(n_1151), .B3(n_1154), .Y(n_1136) );
XOR2xp5_ASAP7_75t_L g797 ( .A(n_798), .B(n_891), .Y(n_797) );
XNOR2xp5_ASAP7_75t_L g798 ( .A(n_799), .B(n_854), .Y(n_798) );
XOR2xp5_ASAP7_75t_L g799 ( .A(n_800), .B(n_853), .Y(n_799) );
NAND3xp33_ASAP7_75t_L g800 ( .A(n_801), .B(n_821), .C(n_851), .Y(n_800) );
INVx2_ASAP7_75t_R g813 ( .A(n_814), .Y(n_813) );
INVx2_ASAP7_75t_L g816 ( .A(n_814), .Y(n_816) );
INVx1_ASAP7_75t_L g818 ( .A(n_819), .Y(n_818) );
INVx1_ASAP7_75t_SL g889 ( .A(n_819), .Y(n_889) );
INVx1_ASAP7_75t_L g1364 ( .A(n_819), .Y(n_1364) );
INVx3_ASAP7_75t_L g1004 ( .A(n_820), .Y(n_1004) );
NAND4xp25_ASAP7_75t_L g822 ( .A(n_823), .B(n_830), .C(n_833), .D(n_834), .Y(n_822) );
OAI211xp5_ASAP7_75t_L g823 ( .A1(n_824), .A2(n_825), .B(n_826), .C(n_828), .Y(n_823) );
BUFx3_ASAP7_75t_L g1738 ( .A(n_827), .Y(n_1738) );
AOI22xp33_ASAP7_75t_L g847 ( .A1(n_831), .A2(n_832), .B1(n_848), .B2(n_849), .Y(n_847) );
OAI22xp5_ASAP7_75t_L g1783 ( .A1(n_837), .A2(n_839), .B1(n_1767), .B2(n_1776), .Y(n_1783) );
INVx2_ASAP7_75t_L g900 ( .A(n_839), .Y(n_900) );
OAI221xp5_ASAP7_75t_L g917 ( .A1(n_839), .A2(n_902), .B1(n_918), .B2(n_919), .C(n_920), .Y(n_917) );
OAI22xp5_ASAP7_75t_L g841 ( .A1(n_842), .A2(n_843), .B1(n_844), .B2(n_845), .Y(n_841) );
AOI222xp33_ASAP7_75t_L g1372 ( .A1(n_848), .A2(n_1351), .B1(n_1373), .B2(n_1374), .C1(n_1375), .C2(n_1376), .Y(n_1372) );
INVx2_ASAP7_75t_SL g1369 ( .A(n_849), .Y(n_1369) );
INVx1_ASAP7_75t_L g855 ( .A(n_856), .Y(n_855) );
NAND3xp33_ASAP7_75t_L g856 ( .A(n_857), .B(n_859), .C(n_880), .Y(n_856) );
AOI21xp5_ASAP7_75t_L g859 ( .A1(n_860), .A2(n_861), .B(n_878), .Y(n_859) );
NAND3xp33_ASAP7_75t_L g861 ( .A(n_862), .B(n_869), .C(n_875), .Y(n_861) );
INVx2_ASAP7_75t_L g1336 ( .A(n_870), .Y(n_1336) );
AND2x4_ASAP7_75t_L g927 ( .A(n_871), .B(n_928), .Y(n_927) );
NAND2xp5_ASAP7_75t_L g881 ( .A(n_882), .B(n_883), .Y(n_881) );
XNOR2x1_ASAP7_75t_L g891 ( .A(n_892), .B(n_983), .Y(n_891) );
XNOR2x1_ASAP7_75t_L g892 ( .A(n_893), .B(n_982), .Y(n_892) );
OR2x2_ASAP7_75t_L g893 ( .A(n_894), .B(n_940), .Y(n_893) );
NAND3xp33_ASAP7_75t_SL g894 ( .A(n_895), .B(n_922), .C(n_934), .Y(n_894) );
AOI211xp5_ASAP7_75t_SL g895 ( .A1(n_896), .A2(n_899), .B(n_905), .C(n_914), .Y(n_895) );
INVxp67_ASAP7_75t_SL g901 ( .A(n_902), .Y(n_901) );
OAI21xp5_ASAP7_75t_L g1426 ( .A1(n_903), .A2(n_912), .B(n_1427), .Y(n_1426) );
OAI33xp33_ASAP7_75t_L g1778 ( .A1(n_903), .A2(n_1779), .A3(n_1780), .B1(n_1782), .B2(n_1783), .B3(n_1784), .Y(n_1778) );
INVx2_ASAP7_75t_L g903 ( .A(n_904), .Y(n_903) );
INVx1_ASAP7_75t_L g1028 ( .A(n_906), .Y(n_1028) );
INVx2_ASAP7_75t_SL g1423 ( .A(n_906), .Y(n_1423) );
NAND2x2_ASAP7_75t_L g906 ( .A(n_907), .B(n_909), .Y(n_906) );
INVx1_ASAP7_75t_L g913 ( .A(n_907), .Y(n_913) );
INVx2_ASAP7_75t_L g907 ( .A(n_908), .Y(n_907) );
INVx2_ASAP7_75t_SL g909 ( .A(n_910), .Y(n_909) );
INVx1_ASAP7_75t_SL g1421 ( .A(n_911), .Y(n_1421) );
CKINVDCx5p33_ASAP7_75t_R g1032 ( .A(n_912), .Y(n_1032) );
INVx1_ASAP7_75t_L g915 ( .A(n_916), .Y(n_915) );
HB1xp67_ASAP7_75t_L g1019 ( .A(n_920), .Y(n_1019) );
INVx2_ASAP7_75t_L g1188 ( .A(n_920), .Y(n_1188) );
NAND2xp5_ASAP7_75t_L g1417 ( .A(n_920), .B(n_1418), .Y(n_1417) );
INVx2_ASAP7_75t_L g1779 ( .A(n_920), .Y(n_1779) );
AOI222xp33_ASAP7_75t_L g922 ( .A1(n_923), .A2(n_926), .B1(n_927), .B2(n_930), .C1(n_931), .C2(n_933), .Y(n_922) );
AOI21xp33_ASAP7_75t_SL g1030 ( .A1(n_923), .A2(n_1031), .B(n_1032), .Y(n_1030) );
AND2x4_ASAP7_75t_L g923 ( .A(n_924), .B(n_925), .Y(n_923) );
AOI222xp33_ASAP7_75t_L g1026 ( .A1(n_927), .A2(n_994), .B1(n_1006), .B2(n_1027), .C1(n_1028), .C2(n_1029), .Y(n_1026) );
INVx1_ASAP7_75t_L g1435 ( .A(n_927), .Y(n_1435) );
INVx1_ASAP7_75t_L g928 ( .A(n_929), .Y(n_928) );
AOI211xp5_ASAP7_75t_L g960 ( .A1(n_930), .A2(n_961), .B(n_964), .C(n_972), .Y(n_960) );
AOI222xp33_ASAP7_75t_L g1014 ( .A1(n_931), .A2(n_995), .B1(n_1015), .B2(n_1019), .C1(n_1020), .C2(n_1023), .Y(n_1014) );
INVx2_ASAP7_75t_L g931 ( .A(n_932), .Y(n_931) );
NAND2xp5_ASAP7_75t_L g934 ( .A(n_935), .B(n_936), .Y(n_934) );
INVx1_ASAP7_75t_L g936 ( .A(n_937), .Y(n_936) );
INVx3_ASAP7_75t_L g937 ( .A(n_938), .Y(n_937) );
HB1xp67_ASAP7_75t_L g985 ( .A(n_938), .Y(n_985) );
AOI22xp33_ASAP7_75t_L g1388 ( .A1(n_938), .A2(n_980), .B1(n_1389), .B2(n_1390), .Y(n_1388) );
AND2x4_ASAP7_75t_L g980 ( .A(n_939), .B(n_981), .Y(n_980) );
AOI221xp5_ASAP7_75t_L g941 ( .A1(n_942), .A2(n_945), .B1(n_947), .B2(n_951), .C(n_954), .Y(n_941) );
INVx2_ASAP7_75t_L g948 ( .A(n_949), .Y(n_948) );
OAI221xp5_ASAP7_75t_L g997 ( .A1(n_949), .A2(n_998), .B1(n_999), .B2(n_1000), .C(n_1001), .Y(n_997) );
OAI221xp5_ASAP7_75t_L g1398 ( .A1(n_949), .A2(n_970), .B1(n_1399), .B2(n_1400), .C(n_1401), .Y(n_1398) );
BUFx2_ASAP7_75t_L g952 ( .A(n_953), .Y(n_952) );
INVx2_ASAP7_75t_L g955 ( .A(n_956), .Y(n_955) );
AOI22xp5_ASAP7_75t_L g1005 ( .A1(n_956), .A2(n_959), .B1(n_986), .B2(n_1006), .Y(n_1005) );
INVx1_ASAP7_75t_L g958 ( .A(n_959), .Y(n_958) );
INVx1_ASAP7_75t_L g961 ( .A(n_962), .Y(n_961) );
INVx2_ASAP7_75t_L g962 ( .A(n_963), .Y(n_962) );
INVx4_ASAP7_75t_L g965 ( .A(n_966), .Y(n_965) );
AOI22xp33_ASAP7_75t_L g993 ( .A1(n_966), .A2(n_968), .B1(n_994), .B2(n_995), .Y(n_993) );
INVx2_ASAP7_75t_L g967 ( .A(n_968), .Y(n_967) );
OAI221xp5_ASAP7_75t_L g1393 ( .A1(n_969), .A2(n_1394), .B1(n_1398), .B2(n_1402), .C(n_1406), .Y(n_1393) );
OR2x6_ASAP7_75t_L g969 ( .A(n_970), .B(n_971), .Y(n_969) );
INVx2_ASAP7_75t_L g974 ( .A(n_975), .Y(n_974) );
HB1xp67_ASAP7_75t_L g1413 ( .A(n_975), .Y(n_1413) );
INVx3_ASAP7_75t_L g976 ( .A(n_977), .Y(n_976) );
NAND2xp5_ASAP7_75t_L g978 ( .A(n_979), .B(n_980), .Y(n_978) );
NAND2xp5_ASAP7_75t_L g988 ( .A(n_980), .B(n_989), .Y(n_988) );
INVx2_ASAP7_75t_L g1370 ( .A(n_980), .Y(n_1370) );
AOI211x1_ASAP7_75t_L g984 ( .A1(n_985), .A2(n_986), .B(n_987), .C(n_1013), .Y(n_984) );
NAND2xp5_ASAP7_75t_L g987 ( .A(n_988), .B(n_990), .Y(n_987) );
NAND3xp33_ASAP7_75t_L g996 ( .A(n_997), .B(n_1005), .C(n_1007), .Y(n_996) );
INVx3_ASAP7_75t_L g1003 ( .A(n_1004), .Y(n_1003) );
OAI211xp5_ASAP7_75t_L g1007 ( .A1(n_1008), .A2(n_1009), .B(n_1011), .C(n_1012), .Y(n_1007) );
OAI21xp5_ASAP7_75t_SL g1406 ( .A1(n_1009), .A2(n_1407), .B(n_1408), .Y(n_1406) );
OAI22xp5_ASAP7_75t_L g1765 ( .A1(n_1009), .A2(n_1210), .B1(n_1766), .B2(n_1767), .Y(n_1765) );
INVx3_ASAP7_75t_L g1009 ( .A(n_1010), .Y(n_1009) );
INVx2_ASAP7_75t_L g1140 ( .A(n_1010), .Y(n_1140) );
NAND3xp33_ASAP7_75t_L g1013 ( .A(n_1014), .B(n_1026), .C(n_1030), .Y(n_1013) );
INVx1_ASAP7_75t_L g1024 ( .A(n_1025), .Y(n_1024) );
INVxp67_ASAP7_75t_L g1484 ( .A(n_1033), .Y(n_1484) );
XNOR2xp5_ASAP7_75t_L g1033 ( .A(n_1034), .B(n_1175), .Y(n_1033) );
INVx2_ASAP7_75t_L g1034 ( .A(n_1035), .Y(n_1034) );
AO22x2_ASAP7_75t_L g1035 ( .A1(n_1036), .A2(n_1037), .B1(n_1128), .B2(n_1174), .Y(n_1035) );
INVx1_ASAP7_75t_L g1036 ( .A(n_1037), .Y(n_1036) );
OAI22xp5_ASAP7_75t_L g1037 ( .A1(n_1038), .A2(n_1039), .B1(n_1082), .B2(n_1127), .Y(n_1037) );
INVx2_ASAP7_75t_L g1038 ( .A(n_1039), .Y(n_1038) );
NAND3xp33_ASAP7_75t_L g1040 ( .A(n_1041), .B(n_1057), .C(n_1060), .Y(n_1040) );
NOR3xp33_ASAP7_75t_L g1041 ( .A(n_1042), .B(n_1054), .C(n_1056), .Y(n_1041) );
NAND2xp5_ASAP7_75t_L g1042 ( .A(n_1043), .B(n_1046), .Y(n_1042) );
INVx1_ASAP7_75t_L g1049 ( .A(n_1050), .Y(n_1049) );
OAI22xp5_ASAP7_75t_L g1768 ( .A1(n_1050), .A2(n_1396), .B1(n_1769), .B2(n_1770), .Y(n_1768) );
NOR3xp33_ASAP7_75t_L g1312 ( .A(n_1056), .B(n_1313), .C(n_1326), .Y(n_1312) );
HB1xp67_ASAP7_75t_L g1075 ( .A(n_1076), .Y(n_1075) );
INVx1_ASAP7_75t_L g1079 ( .A(n_1080), .Y(n_1079) );
INVx2_ASAP7_75t_L g1127 ( .A(n_1082), .Y(n_1127) );
NAND2x1p5_ASAP7_75t_L g1082 ( .A(n_1083), .B(n_1101), .Y(n_1082) );
NAND2xp5_ASAP7_75t_L g1084 ( .A(n_1085), .B(n_1099), .Y(n_1084) );
INVxp67_ASAP7_75t_L g1085 ( .A(n_1086), .Y(n_1085) );
NOR2xp33_ASAP7_75t_SL g1124 ( .A(n_1086), .B(n_1125), .Y(n_1124) );
INVx2_ASAP7_75t_L g1095 ( .A(n_1096), .Y(n_1095) );
NAND2xp5_ASAP7_75t_L g1125 ( .A(n_1099), .B(n_1126), .Y(n_1125) );
INVx1_ASAP7_75t_L g1102 ( .A(n_1103), .Y(n_1102) );
NAND2xp5_ASAP7_75t_L g1103 ( .A(n_1104), .B(n_1108), .Y(n_1103) );
AOI21xp5_ASAP7_75t_L g1104 ( .A1(n_1105), .A2(n_1106), .B(n_1107), .Y(n_1104) );
OAI211xp5_ASAP7_75t_L g1117 ( .A1(n_1118), .A2(n_1119), .B(n_1120), .C(n_1123), .Y(n_1117) );
INVx1_ASAP7_75t_L g1121 ( .A(n_1122), .Y(n_1121) );
INVx1_ASAP7_75t_L g1174 ( .A(n_1128), .Y(n_1174) );
XNOR2xp5_ASAP7_75t_SL g1128 ( .A(n_1129), .B(n_1130), .Y(n_1128) );
AND3x2_ASAP7_75t_L g1130 ( .A(n_1131), .B(n_1156), .C(n_1171), .Y(n_1130) );
NOR4xp25_ASAP7_75t_L g1131 ( .A(n_1132), .B(n_1134), .C(n_1136), .D(n_1155), .Y(n_1131) );
OAI22xp33_ASAP7_75t_L g1137 ( .A1(n_1138), .A2(n_1139), .B1(n_1140), .B2(n_1141), .Y(n_1137) );
OAI22xp5_ASAP7_75t_L g1147 ( .A1(n_1138), .A2(n_1148), .B1(n_1149), .B2(n_1150), .Y(n_1147) );
OAI22xp5_ASAP7_75t_L g1214 ( .A1(n_1138), .A2(n_1183), .B1(n_1198), .B2(n_1215), .Y(n_1214) );
OAI22xp5_ASAP7_75t_L g1402 ( .A1(n_1138), .A2(n_1403), .B1(n_1404), .B2(n_1405), .Y(n_1402) );
OAI22xp33_ASAP7_75t_L g1151 ( .A1(n_1140), .A2(n_1143), .B1(n_1152), .B2(n_1153), .Y(n_1151) );
INVx1_ASAP7_75t_L g1143 ( .A(n_1144), .Y(n_1143) );
OAI33xp33_ASAP7_75t_L g1206 ( .A1(n_1154), .A2(n_1207), .A3(n_1208), .B1(n_1214), .B2(n_1216), .B3(n_1221), .Y(n_1206) );
INVx1_ASAP7_75t_SL g1166 ( .A(n_1167), .Y(n_1166) );
XOR2xp5_ASAP7_75t_L g1175 ( .A(n_1176), .B(n_1328), .Y(n_1175) );
AOI22xp5_ASAP7_75t_L g1176 ( .A1(n_1177), .A2(n_1178), .B1(n_1287), .B2(n_1327), .Y(n_1176) );
INVx1_ASAP7_75t_L g1177 ( .A(n_1178), .Y(n_1177) );
NAND3xp33_ASAP7_75t_L g1179 ( .A(n_1180), .B(n_1225), .C(n_1258), .Y(n_1179) );
NOR2xp33_ASAP7_75t_L g1180 ( .A(n_1181), .B(n_1206), .Y(n_1180) );
OAI33xp33_ASAP7_75t_L g1181 ( .A1(n_1182), .A2(n_1188), .A3(n_1189), .B1(n_1197), .B2(n_1200), .B3(n_1203), .Y(n_1181) );
OAI22xp5_ASAP7_75t_L g1182 ( .A1(n_1183), .A2(n_1184), .B1(n_1185), .B2(n_1186), .Y(n_1182) );
OAI22xp5_ASAP7_75t_L g1203 ( .A1(n_1184), .A2(n_1194), .B1(n_1204), .B2(n_1205), .Y(n_1203) );
OAI22xp5_ASAP7_75t_L g1216 ( .A1(n_1185), .A2(n_1199), .B1(n_1217), .B2(n_1219), .Y(n_1216) );
HB1xp67_ASAP7_75t_L g1186 ( .A(n_1187), .Y(n_1186) );
OAI22xp33_ASAP7_75t_L g1197 ( .A1(n_1187), .A2(n_1191), .B1(n_1198), .B2(n_1199), .Y(n_1197) );
OAI22xp5_ASAP7_75t_L g1189 ( .A1(n_1190), .A2(n_1191), .B1(n_1193), .B2(n_1194), .Y(n_1189) );
OAI22xp33_ASAP7_75t_L g1208 ( .A1(n_1190), .A2(n_1204), .B1(n_1209), .B2(n_1211), .Y(n_1208) );
INVx2_ASAP7_75t_L g1191 ( .A(n_1192), .Y(n_1191) );
OAI22xp5_ASAP7_75t_L g1221 ( .A1(n_1193), .A2(n_1205), .B1(n_1222), .B2(n_1224), .Y(n_1221) );
INVx2_ASAP7_75t_L g1194 ( .A(n_1195), .Y(n_1194) );
INVx2_ASAP7_75t_L g1195 ( .A(n_1196), .Y(n_1195) );
OAI22xp5_ASAP7_75t_L g1784 ( .A1(n_1196), .A2(n_1770), .B1(n_1773), .B2(n_1781), .Y(n_1784) );
INVx2_ASAP7_75t_L g1200 ( .A(n_1201), .Y(n_1200) );
INVx1_ASAP7_75t_L g1201 ( .A(n_1202), .Y(n_1201) );
HB1xp67_ASAP7_75t_L g1209 ( .A(n_1210), .Y(n_1209) );
INVx1_ASAP7_75t_L g1223 ( .A(n_1210), .Y(n_1223) );
OAI22xp5_ASAP7_75t_L g1394 ( .A1(n_1210), .A2(n_1395), .B1(n_1396), .B2(n_1397), .Y(n_1394) );
OAI22xp5_ASAP7_75t_L g1774 ( .A1(n_1210), .A2(n_1220), .B1(n_1775), .B2(n_1776), .Y(n_1774) );
INVx2_ASAP7_75t_SL g1211 ( .A(n_1212), .Y(n_1211) );
INVx1_ASAP7_75t_L g1212 ( .A(n_1213), .Y(n_1212) );
INVx1_ASAP7_75t_L g1217 ( .A(n_1218), .Y(n_1217) );
BUFx6f_ASAP7_75t_L g1219 ( .A(n_1220), .Y(n_1219) );
INVx2_ASAP7_75t_L g1222 ( .A(n_1223), .Y(n_1222) );
OAI221xp5_ASAP7_75t_L g1470 ( .A1(n_1224), .A2(n_1403), .B1(n_1471), .B2(n_1472), .C(n_1473), .Y(n_1470) );
OAI22xp5_ASAP7_75t_L g1771 ( .A1(n_1224), .A2(n_1403), .B1(n_1772), .B2(n_1773), .Y(n_1771) );
OAI31xp33_ASAP7_75t_L g1225 ( .A1(n_1226), .A2(n_1234), .A3(n_1247), .B(n_1253), .Y(n_1225) );
INVx1_ASAP7_75t_L g1227 ( .A(n_1228), .Y(n_1227) );
INVx2_ASAP7_75t_SL g1228 ( .A(n_1229), .Y(n_1228) );
INVx2_ASAP7_75t_L g1231 ( .A(n_1232), .Y(n_1231) );
INVx2_ASAP7_75t_L g1232 ( .A(n_1233), .Y(n_1232) );
CKINVDCx8_ASAP7_75t_R g1235 ( .A(n_1236), .Y(n_1235) );
AOI22xp33_ASAP7_75t_L g1237 ( .A1(n_1238), .A2(n_1239), .B1(n_1243), .B2(n_1244), .Y(n_1237) );
AOI22xp33_ASAP7_75t_L g1277 ( .A1(n_1238), .A2(n_1278), .B1(n_1280), .B2(n_1281), .Y(n_1277) );
BUFx3_ASAP7_75t_L g1239 ( .A(n_1240), .Y(n_1239) );
AND2x2_ASAP7_75t_L g1240 ( .A(n_1241), .B(n_1242), .Y(n_1240) );
AND2x4_ASAP7_75t_L g1245 ( .A(n_1241), .B(n_1246), .Y(n_1245) );
AND2x2_ASAP7_75t_L g1805 ( .A(n_1241), .B(n_1246), .Y(n_1805) );
AND2x4_ASAP7_75t_L g1809 ( .A(n_1241), .B(n_1242), .Y(n_1809) );
BUFx6f_ASAP7_75t_L g1244 ( .A(n_1245), .Y(n_1244) );
INVx1_ASAP7_75t_L g1248 ( .A(n_1249), .Y(n_1248) );
INVx1_ASAP7_75t_L g1249 ( .A(n_1250), .Y(n_1249) );
INVx1_ASAP7_75t_L g1251 ( .A(n_1252), .Y(n_1251) );
AND2x2_ASAP7_75t_SL g1253 ( .A(n_1254), .B(n_1256), .Y(n_1253) );
AND2x2_ASAP7_75t_L g1810 ( .A(n_1254), .B(n_1256), .Y(n_1810) );
INVx1_ASAP7_75t_SL g1254 ( .A(n_1255), .Y(n_1254) );
INVx1_ASAP7_75t_L g1256 ( .A(n_1257), .Y(n_1256) );
OAI31xp33_ASAP7_75t_SL g1258 ( .A1(n_1259), .A2(n_1264), .A3(n_1273), .B(n_1284), .Y(n_1258) );
INVx3_ASAP7_75t_SL g1261 ( .A(n_1262), .Y(n_1261) );
INVx4_ASAP7_75t_L g1799 ( .A(n_1262), .Y(n_1799) );
HB1xp67_ASAP7_75t_L g1265 ( .A(n_1266), .Y(n_1265) );
INVx2_ASAP7_75t_L g1267 ( .A(n_1268), .Y(n_1267) );
INVx2_ASAP7_75t_L g1268 ( .A(n_1269), .Y(n_1268) );
INVx2_ASAP7_75t_L g1269 ( .A(n_1270), .Y(n_1269) );
INVx1_ASAP7_75t_L g1270 ( .A(n_1271), .Y(n_1270) );
INVx3_ASAP7_75t_L g1274 ( .A(n_1275), .Y(n_1274) );
AND2x2_ASAP7_75t_L g1795 ( .A(n_1276), .B(n_1796), .Y(n_1795) );
BUFx3_ASAP7_75t_L g1278 ( .A(n_1279), .Y(n_1278) );
AOI22xp5_ASAP7_75t_L g1790 ( .A1(n_1279), .A2(n_1791), .B1(n_1792), .B2(n_1793), .Y(n_1790) );
INVx2_ASAP7_75t_L g1281 ( .A(n_1282), .Y(n_1281) );
INVx2_ASAP7_75t_L g1282 ( .A(n_1283), .Y(n_1282) );
BUFx3_ASAP7_75t_L g1793 ( .A(n_1283), .Y(n_1793) );
BUFx3_ASAP7_75t_L g1284 ( .A(n_1285), .Y(n_1284) );
OAI31xp33_ASAP7_75t_L g1785 ( .A1(n_1285), .A2(n_1786), .A3(n_1789), .B(n_1797), .Y(n_1785) );
INVx1_ASAP7_75t_L g1327 ( .A(n_1287), .Y(n_1327) );
NAND3xp33_ASAP7_75t_L g1288 ( .A(n_1289), .B(n_1309), .C(n_1312), .Y(n_1288) );
OAI31xp33_ASAP7_75t_L g1289 ( .A1(n_1290), .A2(n_1296), .A3(n_1306), .B(n_1307), .Y(n_1289) );
NAND2xp5_ASAP7_75t_L g1290 ( .A(n_1291), .B(n_1293), .Y(n_1290) );
OAI211xp5_ASAP7_75t_L g1297 ( .A1(n_1298), .A2(n_1299), .B(n_1300), .C(n_1301), .Y(n_1297) );
INVx1_ASAP7_75t_L g1307 ( .A(n_1308), .Y(n_1307) );
NAND2xp5_ASAP7_75t_L g1313 ( .A(n_1314), .B(n_1318), .Y(n_1313) );
HB1xp67_ASAP7_75t_L g1328 ( .A(n_1329), .Y(n_1328) );
INVx1_ASAP7_75t_L g1329 ( .A(n_1330), .Y(n_1329) );
XNOR2xp5_ASAP7_75t_L g1330 ( .A(n_1331), .B(n_1442), .Y(n_1330) );
OAI22xp5_ASAP7_75t_L g1331 ( .A1(n_1332), .A2(n_1384), .B1(n_1440), .B2(n_1441), .Y(n_1331) );
INVx1_ASAP7_75t_L g1441 ( .A(n_1332), .Y(n_1441) );
NAND3xp33_ASAP7_75t_L g1332 ( .A(n_1333), .B(n_1377), .C(n_1381), .Y(n_1332) );
INVx1_ASAP7_75t_L g1378 ( .A(n_1334), .Y(n_1378) );
AOI22xp5_ASAP7_75t_L g1337 ( .A1(n_1338), .A2(n_1339), .B1(n_1340), .B2(n_1342), .Y(n_1337) );
AOI22xp5_ASAP7_75t_L g1343 ( .A1(n_1344), .A2(n_1352), .B1(n_1353), .B2(n_1354), .Y(n_1343) );
INVx3_ASAP7_75t_L g1345 ( .A(n_1346), .Y(n_1345) );
INVx4_ASAP7_75t_L g1450 ( .A(n_1346), .Y(n_1450) );
BUFx6f_ASAP7_75t_L g1749 ( .A(n_1346), .Y(n_1749) );
INVx1_ASAP7_75t_L g1349 ( .A(n_1350), .Y(n_1349) );
AOI22xp5_ASAP7_75t_L g1448 ( .A1(n_1352), .A2(n_1353), .B1(n_1449), .B2(n_1454), .Y(n_1448) );
OAI22xp5_ASAP7_75t_L g1782 ( .A1(n_1355), .A2(n_1428), .B1(n_1769), .B2(n_1772), .Y(n_1782) );
INVx1_ASAP7_75t_L g1379 ( .A(n_1357), .Y(n_1379) );
AND2x2_ASAP7_75t_L g1357 ( .A(n_1358), .B(n_1365), .Y(n_1357) );
INVx1_ASAP7_75t_L g1383 ( .A(n_1367), .Y(n_1383) );
NAND2xp5_ASAP7_75t_L g1367 ( .A(n_1368), .B(n_1371), .Y(n_1367) );
NAND2x1_ASAP7_75t_L g1368 ( .A(n_1369), .B(n_1370), .Y(n_1368) );
INVx1_ASAP7_75t_L g1382 ( .A(n_1372), .Y(n_1382) );
AOI22xp5_ASAP7_75t_L g1465 ( .A1(n_1373), .A2(n_1375), .B1(n_1453), .B2(n_1466), .Y(n_1465) );
OAI21xp5_ASAP7_75t_L g1377 ( .A1(n_1378), .A2(n_1379), .B(n_1380), .Y(n_1377) );
OAI21xp33_ASAP7_75t_L g1381 ( .A1(n_1380), .A2(n_1382), .B(n_1383), .Y(n_1381) );
INVx1_ASAP7_75t_L g1440 ( .A(n_1384), .Y(n_1440) );
XNOR2xp5_ASAP7_75t_L g1384 ( .A(n_1385), .B(n_1386), .Y(n_1384) );
NOR2x1_ASAP7_75t_L g1386 ( .A(n_1387), .B(n_1414), .Y(n_1386) );
NAND2xp5_ASAP7_75t_L g1387 ( .A(n_1388), .B(n_1391), .Y(n_1387) );
OAI211xp5_ASAP7_75t_L g1427 ( .A1(n_1399), .A2(n_1428), .B(n_1430), .C(n_1431), .Y(n_1427) );
AOI22xp5_ASAP7_75t_L g1420 ( .A1(n_1411), .A2(n_1421), .B1(n_1422), .B2(n_1423), .Y(n_1420) );
INVx1_ASAP7_75t_L g1412 ( .A(n_1413), .Y(n_1412) );
NAND3xp33_ASAP7_75t_L g1414 ( .A(n_1415), .B(n_1432), .C(n_1436), .Y(n_1414) );
NOR3xp33_ASAP7_75t_SL g1415 ( .A(n_1416), .B(n_1424), .C(n_1426), .Y(n_1415) );
OAI21xp5_ASAP7_75t_SL g1416 ( .A1(n_1417), .A2(n_1419), .B(n_1420), .Y(n_1416) );
INVx2_ASAP7_75t_L g1428 ( .A(n_1429), .Y(n_1428) );
NAND2xp5_ASAP7_75t_L g1432 ( .A(n_1433), .B(n_1434), .Y(n_1432) );
NAND2xp5_ASAP7_75t_L g1436 ( .A(n_1437), .B(n_1438), .Y(n_1436) );
AOI21xp5_ASAP7_75t_L g1444 ( .A1(n_1445), .A2(n_1463), .B(n_1464), .Y(n_1444) );
NAND4xp25_ASAP7_75t_L g1445 ( .A(n_1446), .B(n_1448), .C(n_1455), .D(n_1459), .Y(n_1445) );
OAI22xp5_ASAP7_75t_SL g1468 ( .A1(n_1469), .A2(n_1470), .B1(n_1474), .B2(n_1475), .Y(n_1468) );
NAND2xp5_ASAP7_75t_L g1479 ( .A(n_1480), .B(n_1481), .Y(n_1479) );
OAI221xp5_ASAP7_75t_L g1485 ( .A1(n_1486), .A2(n_1705), .B1(n_1708), .B2(n_1753), .C(n_1757), .Y(n_1485) );
AOI211xp5_ASAP7_75t_L g1486 ( .A1(n_1487), .A2(n_1610), .B(n_1617), .C(n_1683), .Y(n_1486) );
NAND5xp2_ASAP7_75t_L g1487 ( .A(n_1488), .B(n_1561), .C(n_1588), .D(n_1591), .E(n_1596), .Y(n_1487) );
AOI211xp5_ASAP7_75t_L g1488 ( .A1(n_1489), .A2(n_1519), .B(n_1528), .C(n_1556), .Y(n_1488) );
INVx1_ASAP7_75t_L g1489 ( .A(n_1490), .Y(n_1489) );
OR2x2_ASAP7_75t_L g1490 ( .A(n_1491), .B(n_1506), .Y(n_1490) );
OAI321xp33_ASAP7_75t_L g1528 ( .A1(n_1491), .A2(n_1529), .A3(n_1536), .B1(n_1541), .B2(n_1542), .C(n_1547), .Y(n_1528) );
AND2x2_ASAP7_75t_L g1549 ( .A(n_1491), .B(n_1507), .Y(n_1549) );
AND3x1_ASAP7_75t_L g1582 ( .A(n_1491), .B(n_1516), .C(n_1540), .Y(n_1582) );
AND2x2_ASAP7_75t_L g1587 ( .A(n_1491), .B(n_1574), .Y(n_1587) );
NAND2xp5_ASAP7_75t_L g1607 ( .A(n_1491), .B(n_1516), .Y(n_1607) );
OR2x2_ASAP7_75t_L g1634 ( .A(n_1491), .B(n_1635), .Y(n_1634) );
AND2x2_ASAP7_75t_L g1637 ( .A(n_1491), .B(n_1537), .Y(n_1637) );
NAND2xp5_ASAP7_75t_L g1676 ( .A(n_1491), .B(n_1540), .Y(n_1676) );
INVx2_ASAP7_75t_L g1491 ( .A(n_1492), .Y(n_1491) );
AND2x2_ASAP7_75t_L g1546 ( .A(n_1492), .B(n_1537), .Y(n_1546) );
BUFx2_ASAP7_75t_L g1552 ( .A(n_1492), .Y(n_1552) );
OR2x2_ASAP7_75t_L g1643 ( .A(n_1492), .B(n_1629), .Y(n_1643) );
AND2x2_ASAP7_75t_L g1655 ( .A(n_1492), .B(n_1574), .Y(n_1655) );
AND2x2_ASAP7_75t_L g1492 ( .A(n_1493), .B(n_1501), .Y(n_1492) );
AND2x4_ASAP7_75t_L g1494 ( .A(n_1495), .B(n_1496), .Y(n_1494) );
AND2x6_ASAP7_75t_L g1499 ( .A(n_1495), .B(n_1500), .Y(n_1499) );
AND2x6_ASAP7_75t_L g1502 ( .A(n_1495), .B(n_1503), .Y(n_1502) );
AND2x2_ASAP7_75t_L g1504 ( .A(n_1495), .B(n_1505), .Y(n_1504) );
AND2x2_ASAP7_75t_L g1511 ( .A(n_1495), .B(n_1505), .Y(n_1511) );
AND2x2_ASAP7_75t_L g1523 ( .A(n_1495), .B(n_1505), .Y(n_1523) );
NAND2xp5_ASAP7_75t_L g1707 ( .A(n_1495), .B(n_1496), .Y(n_1707) );
HB1xp67_ASAP7_75t_L g1813 ( .A(n_1496), .Y(n_1813) );
AND2x2_ASAP7_75t_L g1496 ( .A(n_1497), .B(n_1498), .Y(n_1496) );
INVx2_ASAP7_75t_L g1614 ( .A(n_1502), .Y(n_1614) );
NAND2xp5_ASAP7_75t_L g1506 ( .A(n_1507), .B(n_1512), .Y(n_1506) );
AND2x2_ASAP7_75t_L g1530 ( .A(n_1507), .B(n_1531), .Y(n_1530) );
NOR2xp33_ASAP7_75t_L g1564 ( .A(n_1507), .B(n_1565), .Y(n_1564) );
INVx1_ASAP7_75t_L g1599 ( .A(n_1507), .Y(n_1599) );
NAND2xp5_ASAP7_75t_L g1625 ( .A(n_1507), .B(n_1569), .Y(n_1625) );
NOR2xp33_ASAP7_75t_L g1659 ( .A(n_1507), .B(n_1660), .Y(n_1659) );
NAND2xp5_ASAP7_75t_L g1694 ( .A(n_1507), .B(n_1537), .Y(n_1694) );
INVx2_ASAP7_75t_L g1507 ( .A(n_1508), .Y(n_1507) );
INVx1_ASAP7_75t_L g1545 ( .A(n_1508), .Y(n_1545) );
AND2x2_ASAP7_75t_L g1551 ( .A(n_1508), .B(n_1552), .Y(n_1551) );
AND2x2_ASAP7_75t_L g1580 ( .A(n_1508), .B(n_1521), .Y(n_1580) );
NAND2xp5_ASAP7_75t_L g1629 ( .A(n_1508), .B(n_1512), .Y(n_1629) );
NOR2xp33_ASAP7_75t_L g1631 ( .A(n_1508), .B(n_1632), .Y(n_1631) );
AND2x2_ASAP7_75t_L g1675 ( .A(n_1508), .B(n_1532), .Y(n_1675) );
AND2x2_ASAP7_75t_L g1508 ( .A(n_1509), .B(n_1510), .Y(n_1508) );
INVxp67_ASAP7_75t_L g1616 ( .A(n_1511), .Y(n_1616) );
AND2x2_ASAP7_75t_L g1645 ( .A(n_1512), .B(n_1551), .Y(n_1645) );
AND2x2_ASAP7_75t_L g1512 ( .A(n_1513), .B(n_1516), .Y(n_1512) );
AND2x2_ASAP7_75t_L g1537 ( .A(n_1513), .B(n_1538), .Y(n_1537) );
INVx2_ASAP7_75t_L g1540 ( .A(n_1513), .Y(n_1540) );
NAND2xp5_ASAP7_75t_L g1565 ( .A(n_1513), .B(n_1552), .Y(n_1565) );
NAND3xp33_ASAP7_75t_L g1638 ( .A(n_1513), .B(n_1543), .C(n_1611), .Y(n_1638) );
OR2x2_ASAP7_75t_L g1513 ( .A(n_1514), .B(n_1515), .Y(n_1513) );
INVx1_ASAP7_75t_L g1538 ( .A(n_1516), .Y(n_1538) );
AND2x2_ASAP7_75t_L g1539 ( .A(n_1516), .B(n_1540), .Y(n_1539) );
AND2x2_ASAP7_75t_L g1624 ( .A(n_1516), .B(n_1552), .Y(n_1624) );
OR2x2_ASAP7_75t_L g1660 ( .A(n_1516), .B(n_1552), .Y(n_1660) );
AND2x2_ASAP7_75t_L g1516 ( .A(n_1517), .B(n_1518), .Y(n_1516) );
A2O1A1Ixp33_ASAP7_75t_L g1627 ( .A1(n_1519), .A2(n_1611), .B(n_1628), .C(n_1630), .Y(n_1627) );
INVx1_ASAP7_75t_L g1519 ( .A(n_1520), .Y(n_1519) );
OR2x2_ASAP7_75t_L g1520 ( .A(n_1521), .B(n_1525), .Y(n_1520) );
CKINVDCx6p67_ASAP7_75t_R g1554 ( .A(n_1521), .Y(n_1554) );
OR2x2_ASAP7_75t_L g1558 ( .A(n_1521), .B(n_1559), .Y(n_1558) );
NAND2xp5_ASAP7_75t_L g1601 ( .A(n_1521), .B(n_1569), .Y(n_1601) );
AND2x2_ASAP7_75t_L g1609 ( .A(n_1521), .B(n_1525), .Y(n_1609) );
NAND2xp5_ASAP7_75t_L g1691 ( .A(n_1521), .B(n_1611), .Y(n_1691) );
NAND2xp5_ASAP7_75t_L g1698 ( .A(n_1521), .B(n_1699), .Y(n_1698) );
OR2x6_ASAP7_75t_L g1521 ( .A(n_1522), .B(n_1524), .Y(n_1521) );
INVx1_ASAP7_75t_L g1535 ( .A(n_1525), .Y(n_1535) );
INVx3_ASAP7_75t_L g1541 ( .A(n_1525), .Y(n_1541) );
AND2x2_ASAP7_75t_L g1560 ( .A(n_1525), .B(n_1555), .Y(n_1560) );
OR2x2_ASAP7_75t_L g1563 ( .A(n_1525), .B(n_1532), .Y(n_1563) );
AND2x2_ASAP7_75t_L g1575 ( .A(n_1525), .B(n_1554), .Y(n_1575) );
AND2x2_ASAP7_75t_L g1578 ( .A(n_1525), .B(n_1532), .Y(n_1578) );
OR2x2_ASAP7_75t_L g1593 ( .A(n_1525), .B(n_1554), .Y(n_1593) );
OAI221xp5_ASAP7_75t_L g1652 ( .A1(n_1525), .A2(n_1653), .B1(n_1654), .B2(n_1656), .C(n_1657), .Y(n_1652) );
OAI32xp33_ASAP7_75t_L g1679 ( .A1(n_1525), .A2(n_1541), .A3(n_1543), .B1(n_1634), .B2(n_1680), .Y(n_1679) );
AND2x4_ASAP7_75t_L g1525 ( .A(n_1526), .B(n_1527), .Y(n_1525) );
OAI32xp33_ASAP7_75t_L g1696 ( .A1(n_1529), .A2(n_1543), .A3(n_1583), .B1(n_1697), .B2(n_1698), .Y(n_1696) );
INVx1_ASAP7_75t_L g1529 ( .A(n_1530), .Y(n_1529) );
INVx1_ASAP7_75t_L g1583 ( .A(n_1531), .Y(n_1583) );
AND2x2_ASAP7_75t_L g1640 ( .A(n_1531), .B(n_1554), .Y(n_1640) );
AND2x2_ASAP7_75t_L g1531 ( .A(n_1532), .B(n_1535), .Y(n_1531) );
INVx1_ASAP7_75t_L g1555 ( .A(n_1532), .Y(n_1555) );
AND2x2_ASAP7_75t_L g1532 ( .A(n_1533), .B(n_1534), .Y(n_1532) );
OR2x2_ASAP7_75t_L g1536 ( .A(n_1537), .B(n_1539), .Y(n_1536) );
AND2x2_ASAP7_75t_L g1550 ( .A(n_1537), .B(n_1551), .Y(n_1550) );
AND2x2_ASAP7_75t_L g1574 ( .A(n_1538), .B(n_1540), .Y(n_1574) );
O2A1O1Ixp33_ASAP7_75t_L g1647 ( .A1(n_1538), .A2(n_1648), .B(n_1649), .C(n_1650), .Y(n_1647) );
AND2x2_ASAP7_75t_L g1548 ( .A(n_1539), .B(n_1549), .Y(n_1548) );
INVx1_ASAP7_75t_L g1557 ( .A(n_1539), .Y(n_1557) );
AND2x2_ASAP7_75t_L g1595 ( .A(n_1539), .B(n_1552), .Y(n_1595) );
OAI322xp33_ASAP7_75t_L g1576 ( .A1(n_1540), .A2(n_1577), .A3(n_1579), .B1(n_1581), .B2(n_1583), .C1(n_1584), .C2(n_1586), .Y(n_1576) );
OR2x2_ASAP7_75t_L g1632 ( .A(n_1540), .B(n_1552), .Y(n_1632) );
AND2x2_ASAP7_75t_L g1681 ( .A(n_1540), .B(n_1552), .Y(n_1681) );
CKINVDCx14_ASAP7_75t_R g1672 ( .A(n_1541), .Y(n_1672) );
NAND2xp5_ASAP7_75t_L g1542 ( .A(n_1543), .B(n_1546), .Y(n_1542) );
NAND2xp5_ASAP7_75t_L g1669 ( .A(n_1543), .B(n_1637), .Y(n_1669) );
INVx1_ASAP7_75t_L g1543 ( .A(n_1544), .Y(n_1543) );
NAND2xp5_ASAP7_75t_L g1590 ( .A(n_1544), .B(n_1587), .Y(n_1590) );
NAND2xp5_ASAP7_75t_L g1648 ( .A(n_1544), .B(n_1585), .Y(n_1648) );
AND2x2_ASAP7_75t_L g1666 ( .A(n_1544), .B(n_1637), .Y(n_1666) );
INVx2_ASAP7_75t_L g1544 ( .A(n_1545), .Y(n_1544) );
AND2x2_ASAP7_75t_L g1594 ( .A(n_1545), .B(n_1595), .Y(n_1594) );
NAND2xp5_ASAP7_75t_L g1635 ( .A(n_1545), .B(n_1574), .Y(n_1635) );
AND2x2_ASAP7_75t_L g1685 ( .A(n_1545), .B(n_1585), .Y(n_1685) );
AND2x2_ASAP7_75t_L g1702 ( .A(n_1546), .B(n_1569), .Y(n_1702) );
OAI21xp5_ASAP7_75t_L g1547 ( .A1(n_1548), .A2(n_1550), .B(n_1553), .Y(n_1547) );
INVx1_ASAP7_75t_L g1626 ( .A(n_1548), .Y(n_1626) );
AND2x2_ASAP7_75t_L g1604 ( .A(n_1549), .B(n_1574), .Y(n_1604) );
INVx1_ASAP7_75t_L g1689 ( .A(n_1550), .Y(n_1689) );
INVx1_ASAP7_75t_L g1572 ( .A(n_1551), .Y(n_1572) );
INVx1_ASAP7_75t_L g1642 ( .A(n_1553), .Y(n_1642) );
NAND2xp5_ASAP7_75t_L g1654 ( .A(n_1553), .B(n_1655), .Y(n_1654) );
AND2x2_ASAP7_75t_L g1553 ( .A(n_1554), .B(n_1555), .Y(n_1553) );
NOR2xp33_ASAP7_75t_L g1562 ( .A(n_1554), .B(n_1563), .Y(n_1562) );
NAND2xp5_ASAP7_75t_L g1584 ( .A(n_1554), .B(n_1585), .Y(n_1584) );
NOR2xp33_ASAP7_75t_SL g1646 ( .A(n_1554), .B(n_1583), .Y(n_1646) );
NAND2xp5_ASAP7_75t_L g1650 ( .A(n_1554), .B(n_1611), .Y(n_1650) );
AND2x2_ASAP7_75t_L g1664 ( .A(n_1554), .B(n_1569), .Y(n_1664) );
INVx2_ASAP7_75t_L g1569 ( .A(n_1555), .Y(n_1569) );
NOR2xp33_ASAP7_75t_L g1556 ( .A(n_1557), .B(n_1558), .Y(n_1556) );
INVx1_ASAP7_75t_L g1695 ( .A(n_1558), .Y(n_1695) );
OAI22xp5_ASAP7_75t_L g1662 ( .A1(n_1559), .A2(n_1634), .B1(n_1663), .B2(n_1665), .Y(n_1662) );
OAI211xp5_ASAP7_75t_L g1670 ( .A1(n_1559), .A2(n_1636), .B(n_1671), .C(n_1677), .Y(n_1670) );
CKINVDCx6p67_ASAP7_75t_R g1559 ( .A(n_1560), .Y(n_1559) );
NAND2xp5_ASAP7_75t_L g1598 ( .A(n_1560), .B(n_1599), .Y(n_1598) );
AOI221xp5_ASAP7_75t_L g1561 ( .A1(n_1562), .A2(n_1564), .B1(n_1566), .B2(n_1575), .C(n_1576), .Y(n_1561) );
INVx2_ASAP7_75t_L g1585 ( .A(n_1563), .Y(n_1585) );
AND2x2_ASAP7_75t_L g1566 ( .A(n_1567), .B(n_1570), .Y(n_1566) );
AND2x2_ASAP7_75t_L g1658 ( .A(n_1567), .B(n_1659), .Y(n_1658) );
A2O1A1Ixp33_ASAP7_75t_L g1686 ( .A1(n_1567), .A2(n_1635), .B(n_1636), .C(n_1687), .Y(n_1686) );
INVx2_ASAP7_75t_L g1567 ( .A(n_1568), .Y(n_1567) );
NAND2xp5_ASAP7_75t_L g1588 ( .A(n_1568), .B(n_1589), .Y(n_1588) );
NAND2xp5_ASAP7_75t_L g1608 ( .A(n_1568), .B(n_1609), .Y(n_1608) );
NOR2xp33_ASAP7_75t_L g1688 ( .A(n_1568), .B(n_1689), .Y(n_1688) );
NAND2xp5_ASAP7_75t_L g1704 ( .A(n_1568), .B(n_1666), .Y(n_1704) );
INVx2_ASAP7_75t_L g1568 ( .A(n_1569), .Y(n_1568) );
OR2x2_ASAP7_75t_L g1653 ( .A(n_1569), .B(n_1571), .Y(n_1653) );
INVx1_ASAP7_75t_L g1570 ( .A(n_1571), .Y(n_1570) );
OR2x2_ASAP7_75t_L g1571 ( .A(n_1572), .B(n_1573), .Y(n_1571) );
INVx1_ASAP7_75t_L g1573 ( .A(n_1574), .Y(n_1573) );
INVx1_ASAP7_75t_L g1620 ( .A(n_1575), .Y(n_1620) );
AND2x2_ASAP7_75t_L g1630 ( .A(n_1575), .B(n_1631), .Y(n_1630) );
OAI22xp5_ASAP7_75t_L g1602 ( .A1(n_1577), .A2(n_1603), .B1(n_1605), .B2(n_1608), .Y(n_1602) );
NOR2xp33_ASAP7_75t_L g1678 ( .A(n_1577), .B(n_1581), .Y(n_1678) );
INVx2_ASAP7_75t_L g1577 ( .A(n_1578), .Y(n_1577) );
AOI22xp33_ASAP7_75t_L g1644 ( .A1(n_1578), .A2(n_1582), .B1(n_1645), .B2(n_1646), .Y(n_1644) );
CKINVDCx14_ASAP7_75t_R g1579 ( .A(n_1580), .Y(n_1579) );
INVx2_ASAP7_75t_L g1581 ( .A(n_1582), .Y(n_1581) );
INVx1_ASAP7_75t_L g1586 ( .A(n_1587), .Y(n_1586) );
O2A1O1Ixp33_ASAP7_75t_L g1692 ( .A1(n_1589), .A2(n_1693), .B(n_1695), .C(n_1696), .Y(n_1692) );
INVx1_ASAP7_75t_L g1589 ( .A(n_1590), .Y(n_1589) );
NAND2xp5_ASAP7_75t_L g1591 ( .A(n_1592), .B(n_1594), .Y(n_1591) );
INVx1_ASAP7_75t_L g1592 ( .A(n_1593), .Y(n_1592) );
O2A1O1Ixp33_ASAP7_75t_L g1596 ( .A1(n_1595), .A2(n_1597), .B(n_1600), .C(n_1602), .Y(n_1596) );
NOR2xp33_ASAP7_75t_L g1697 ( .A(n_1595), .B(n_1637), .Y(n_1697) );
INVx1_ASAP7_75t_L g1597 ( .A(n_1598), .Y(n_1597) );
NOR2xp33_ASAP7_75t_L g1606 ( .A(n_1599), .B(n_1607), .Y(n_1606) );
INVx1_ASAP7_75t_L g1600 ( .A(n_1601), .Y(n_1600) );
OAI221xp5_ASAP7_75t_L g1619 ( .A1(n_1601), .A2(n_1620), .B1(n_1621), .B2(n_1626), .C(n_1627), .Y(n_1619) );
INVx1_ASAP7_75t_L g1603 ( .A(n_1604), .Y(n_1603) );
INVx1_ASAP7_75t_L g1605 ( .A(n_1606), .Y(n_1605) );
OAI31xp33_ASAP7_75t_L g1700 ( .A1(n_1609), .A2(n_1701), .A3(n_1702), .B(n_1703), .Y(n_1700) );
INVx2_ASAP7_75t_SL g1610 ( .A(n_1611), .Y(n_1610) );
INVx2_ASAP7_75t_SL g1656 ( .A(n_1611), .Y(n_1656) );
OAI22xp5_ASAP7_75t_SL g1612 ( .A1(n_1613), .A2(n_1614), .B1(n_1615), .B2(n_1616), .Y(n_1612) );
NAND3xp33_ASAP7_75t_L g1617 ( .A(n_1618), .B(n_1651), .C(n_1667), .Y(n_1617) );
NOR4xp25_ASAP7_75t_L g1618 ( .A(n_1619), .B(n_1633), .C(n_1641), .D(n_1647), .Y(n_1618) );
INVx1_ASAP7_75t_L g1621 ( .A(n_1622), .Y(n_1621) );
OAI21xp5_ASAP7_75t_L g1657 ( .A1(n_1622), .A2(n_1658), .B(n_1661), .Y(n_1657) );
NOR2xp33_ASAP7_75t_L g1622 ( .A(n_1623), .B(n_1625), .Y(n_1622) );
A2O1A1Ixp33_ASAP7_75t_L g1684 ( .A1(n_1623), .A2(n_1685), .B(n_1686), .C(n_1690), .Y(n_1684) );
INVx1_ASAP7_75t_L g1623 ( .A(n_1624), .Y(n_1623) );
INVx1_ASAP7_75t_L g1628 ( .A(n_1629), .Y(n_1628) );
AOI31xp33_ASAP7_75t_L g1633 ( .A1(n_1634), .A2(n_1636), .A3(n_1638), .B(n_1639), .Y(n_1633) );
INVx1_ASAP7_75t_L g1701 ( .A(n_1634), .Y(n_1701) );
INVx1_ASAP7_75t_L g1636 ( .A(n_1637), .Y(n_1636) );
INVx1_ASAP7_75t_L g1639 ( .A(n_1640), .Y(n_1639) );
OAI21xp33_ASAP7_75t_L g1641 ( .A1(n_1642), .A2(n_1643), .B(n_1644), .Y(n_1641) );
INVx1_ASAP7_75t_L g1649 ( .A(n_1645), .Y(n_1649) );
INVx1_ASAP7_75t_L g1661 ( .A(n_1650), .Y(n_1661) );
NOR2xp33_ASAP7_75t_L g1651 ( .A(n_1652), .B(n_1662), .Y(n_1651) );
INVx3_ASAP7_75t_L g1682 ( .A(n_1656), .Y(n_1682) );
INVx1_ASAP7_75t_L g1663 ( .A(n_1664), .Y(n_1663) );
INVx1_ASAP7_75t_L g1665 ( .A(n_1666), .Y(n_1665) );
OAI31xp33_ASAP7_75t_L g1667 ( .A1(n_1668), .A2(n_1670), .A3(n_1679), .B(n_1682), .Y(n_1667) );
INVx1_ASAP7_75t_L g1668 ( .A(n_1669), .Y(n_1668) );
NAND2xp5_ASAP7_75t_L g1671 ( .A(n_1672), .B(n_1673), .Y(n_1671) );
NOR2xp33_ASAP7_75t_L g1673 ( .A(n_1674), .B(n_1676), .Y(n_1673) );
CKINVDCx14_ASAP7_75t_R g1674 ( .A(n_1675), .Y(n_1674) );
INVx1_ASAP7_75t_L g1699 ( .A(n_1676), .Y(n_1699) );
INVx1_ASAP7_75t_L g1677 ( .A(n_1678), .Y(n_1677) );
CKINVDCx14_ASAP7_75t_R g1680 ( .A(n_1681), .Y(n_1680) );
NAND3xp33_ASAP7_75t_L g1683 ( .A(n_1684), .B(n_1692), .C(n_1700), .Y(n_1683) );
INVxp67_ASAP7_75t_L g1687 ( .A(n_1688), .Y(n_1687) );
INVx1_ASAP7_75t_L g1690 ( .A(n_1691), .Y(n_1690) );
INVx1_ASAP7_75t_L g1693 ( .A(n_1694), .Y(n_1693) );
INVx1_ASAP7_75t_L g1703 ( .A(n_1704), .Y(n_1703) );
CKINVDCx20_ASAP7_75t_R g1705 ( .A(n_1706), .Y(n_1705) );
CKINVDCx5p33_ASAP7_75t_R g1706 ( .A(n_1707), .Y(n_1706) );
INVx1_ASAP7_75t_L g1709 ( .A(n_1710), .Y(n_1709) );
HB1xp67_ASAP7_75t_L g1710 ( .A(n_1711), .Y(n_1710) );
NAND2xp5_ASAP7_75t_SL g1711 ( .A(n_1712), .B(n_1732), .Y(n_1711) );
NAND2xp5_ASAP7_75t_L g1714 ( .A(n_1715), .B(n_1722), .Y(n_1714) );
NOR2xp33_ASAP7_75t_L g1715 ( .A(n_1716), .B(n_1719), .Y(n_1715) );
NAND3xp33_ASAP7_75t_SL g1733 ( .A(n_1734), .B(n_1735), .C(n_1740), .Y(n_1733) );
OAI22xp5_ASAP7_75t_L g1746 ( .A1(n_1747), .A2(n_1748), .B1(n_1750), .B2(n_1751), .Y(n_1746) );
INVx2_ASAP7_75t_L g1748 ( .A(n_1749), .Y(n_1748) );
CKINVDCx5p33_ASAP7_75t_R g1753 ( .A(n_1754), .Y(n_1753) );
BUFx2_ASAP7_75t_SL g1754 ( .A(n_1755), .Y(n_1754) );
BUFx3_ASAP7_75t_L g1755 ( .A(n_1756), .Y(n_1755) );
INVx1_ASAP7_75t_L g1760 ( .A(n_1761), .Y(n_1760) );
NAND3xp33_ASAP7_75t_L g1762 ( .A(n_1763), .B(n_1785), .C(n_1800), .Y(n_1762) );
NOR2xp33_ASAP7_75t_SL g1763 ( .A(n_1764), .B(n_1778), .Y(n_1763) );
AOI22xp5_ASAP7_75t_L g1806 ( .A1(n_1791), .A2(n_1807), .B1(n_1808), .B2(n_1809), .Y(n_1806) );
INVx2_ASAP7_75t_L g1794 ( .A(n_1795), .Y(n_1794) );
OAI31xp33_ASAP7_75t_SL g1800 ( .A1(n_1801), .A2(n_1802), .A3(n_1803), .B(n_1810), .Y(n_1800) );
INVxp67_ASAP7_75t_L g1804 ( .A(n_1805), .Y(n_1804) );
OAI21xp5_ASAP7_75t_L g1811 ( .A1(n_1812), .A2(n_1813), .B(n_1814), .Y(n_1811) );
INVx1_ASAP7_75t_L g1814 ( .A(n_1815), .Y(n_1814) );
endmodule