module fake_jpeg_26324_n_196 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_196);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_196;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_186;
wire n_44;
wire n_24;
wire n_143;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_177;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_128;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_183;
wire n_79;
wire n_170;
wire n_162;
wire n_132;
wire n_133;
wire n_67;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_161;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_189;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_140;
wire n_96;

BUFx16f_ASAP7_75t_L g16 ( 
.A(n_4),
.Y(n_16)
);

INVx2_ASAP7_75t_L g17 ( 
.A(n_8),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_7),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_9),
.Y(n_19)
);

INVx5_ASAP7_75t_L g20 ( 
.A(n_10),
.Y(n_20)
);

INVx11_ASAP7_75t_SL g21 ( 
.A(n_2),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_11),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_10),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_13),
.Y(n_24)
);

INVx2_ASAP7_75t_L g25 ( 
.A(n_14),
.Y(n_25)
);

BUFx12_ASAP7_75t_L g26 ( 
.A(n_8),
.Y(n_26)
);

INVx11_ASAP7_75t_L g27 ( 
.A(n_7),
.Y(n_27)
);

INVx3_ASAP7_75t_L g28 ( 
.A(n_6),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_3),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_6),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_15),
.Y(n_31)
);

BUFx6f_ASAP7_75t_SL g32 ( 
.A(n_0),
.Y(n_32)
);

INVx6_ASAP7_75t_L g33 ( 
.A(n_16),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_33),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_SL g34 ( 
.A(n_16),
.B(n_0),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_L g45 ( 
.A(n_34),
.B(n_37),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_32),
.Y(n_35)
);

INVx2_ASAP7_75t_L g50 ( 
.A(n_35),
.Y(n_50)
);

INVx5_ASAP7_75t_L g36 ( 
.A(n_16),
.Y(n_36)
);

INVx11_ASAP7_75t_L g55 ( 
.A(n_36),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_27),
.Y(n_37)
);

BUFx3_ASAP7_75t_L g38 ( 
.A(n_32),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_38),
.B(n_41),
.Y(n_56)
);

CKINVDCx9p33_ASAP7_75t_R g39 ( 
.A(n_21),
.Y(n_39)
);

BUFx8_ASAP7_75t_L g61 ( 
.A(n_39),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_SL g40 ( 
.A(n_30),
.B(n_0),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_SL g52 ( 
.A(n_40),
.B(n_18),
.Y(n_52)
);

INVx2_ASAP7_75t_SL g41 ( 
.A(n_21),
.Y(n_41)
);

INVx11_ASAP7_75t_L g42 ( 
.A(n_27),
.Y(n_42)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_42),
.Y(n_49)
);

INVx8_ASAP7_75t_L g43 ( 
.A(n_27),
.Y(n_43)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_43),
.Y(n_57)
);

OAI22xp5_ASAP7_75t_L g44 ( 
.A1(n_34),
.A2(n_28),
.B1(n_17),
.B2(n_25),
.Y(n_44)
);

AOI22xp5_ASAP7_75t_L g77 ( 
.A1(n_44),
.A2(n_51),
.B1(n_41),
.B2(n_42),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_L g46 ( 
.A(n_34),
.B(n_17),
.Y(n_46)
);

A2O1A1Ixp33_ASAP7_75t_L g74 ( 
.A1(n_46),
.A2(n_48),
.B(n_60),
.C(n_29),
.Y(n_74)
);

AOI22xp5_ASAP7_75t_L g47 ( 
.A1(n_42),
.A2(n_28),
.B1(n_25),
.B2(n_20),
.Y(n_47)
);

OAI22xp5_ASAP7_75t_SL g76 ( 
.A1(n_47),
.A2(n_41),
.B1(n_42),
.B2(n_43),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_L g48 ( 
.A(n_40),
.B(n_29),
.Y(n_48)
);

OAI22xp33_ASAP7_75t_SL g51 ( 
.A1(n_33),
.A2(n_28),
.B1(n_20),
.B2(n_30),
.Y(n_51)
);

OR2x2_ASAP7_75t_L g73 ( 
.A(n_52),
.B(n_59),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_40),
.B(n_31),
.Y(n_54)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_54),
.Y(n_80)
);

BUFx3_ASAP7_75t_L g58 ( 
.A(n_36),
.Y(n_58)
);

INVx2_ASAP7_75t_L g84 ( 
.A(n_58),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_SL g59 ( 
.A(n_36),
.B(n_31),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_SL g60 ( 
.A(n_43),
.B(n_18),
.Y(n_60)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_43),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_62),
.B(n_41),
.Y(n_63)
);

CKINVDCx16_ASAP7_75t_R g94 ( 
.A(n_63),
.Y(n_94)
);

CKINVDCx16_ASAP7_75t_R g64 ( 
.A(n_56),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_64),
.B(n_70),
.Y(n_88)
);

INVx2_ASAP7_75t_L g65 ( 
.A(n_50),
.Y(n_65)
);

INVx2_ASAP7_75t_L g95 ( 
.A(n_65),
.Y(n_95)
);

AOI22xp33_ASAP7_75t_SL g66 ( 
.A1(n_50),
.A2(n_20),
.B1(n_36),
.B2(n_33),
.Y(n_66)
);

BUFx10_ASAP7_75t_L g98 ( 
.A(n_66),
.Y(n_98)
);

INVx2_ASAP7_75t_L g67 ( 
.A(n_53),
.Y(n_67)
);

INVx2_ASAP7_75t_L g106 ( 
.A(n_67),
.Y(n_106)
);

AOI21xp33_ASAP7_75t_L g68 ( 
.A1(n_48),
.A2(n_19),
.B(n_24),
.Y(n_68)
);

MAJIxp5_ASAP7_75t_L g100 ( 
.A(n_68),
.B(n_26),
.C(n_35),
.Y(n_100)
);

AOI22xp5_ASAP7_75t_SL g69 ( 
.A1(n_44),
.A2(n_19),
.B1(n_22),
.B2(n_23),
.Y(n_69)
);

NOR2x1_ASAP7_75t_L g107 ( 
.A(n_69),
.B(n_77),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_59),
.B(n_22),
.Y(n_70)
);

INVxp67_ASAP7_75t_L g71 ( 
.A(n_56),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_SL g86 ( 
.A(n_71),
.B(n_78),
.Y(n_86)
);

OAI22xp5_ASAP7_75t_L g72 ( 
.A1(n_46),
.A2(n_23),
.B1(n_24),
.B2(n_33),
.Y(n_72)
);

AOI22xp5_ASAP7_75t_L g89 ( 
.A1(n_72),
.A2(n_76),
.B1(n_81),
.B2(n_45),
.Y(n_89)
);

XOR2xp5_ASAP7_75t_L g101 ( 
.A(n_74),
.B(n_38),
.Y(n_101)
);

INVx2_ASAP7_75t_L g75 ( 
.A(n_53),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_75),
.B(n_79),
.Y(n_91)
);

OR2x2_ASAP7_75t_L g78 ( 
.A(n_52),
.B(n_29),
.Y(n_78)
);

INVx3_ASAP7_75t_L g79 ( 
.A(n_53),
.Y(n_79)
);

AOI22xp5_ASAP7_75t_L g81 ( 
.A1(n_45),
.A2(n_41),
.B1(n_35),
.B2(n_38),
.Y(n_81)
);

INVx2_ASAP7_75t_L g82 ( 
.A(n_55),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_82),
.B(n_83),
.Y(n_97)
);

INVx2_ASAP7_75t_L g83 ( 
.A(n_55),
.Y(n_83)
);

BUFx12f_ASAP7_75t_SL g85 ( 
.A(n_61),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_85),
.B(n_58),
.Y(n_99)
);

CKINVDCx20_ASAP7_75t_R g87 ( 
.A(n_81),
.Y(n_87)
);

CKINVDCx20_ASAP7_75t_R g117 ( 
.A(n_87),
.Y(n_117)
);

AND2x2_ASAP7_75t_L g108 ( 
.A(n_89),
.B(n_101),
.Y(n_108)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_76),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_SL g123 ( 
.A(n_90),
.B(n_92),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_SL g92 ( 
.A(n_73),
.B(n_60),
.Y(n_92)
);

O2A1O1Ixp33_ASAP7_75t_L g93 ( 
.A1(n_71),
.A2(n_49),
.B(n_47),
.C(n_62),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_L g116 ( 
.A(n_93),
.B(n_96),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_L g96 ( 
.A(n_78),
.B(n_49),
.Y(n_96)
);

NOR3xp33_ASAP7_75t_L g126 ( 
.A(n_99),
.B(n_100),
.C(n_79),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_80),
.B(n_73),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_L g112 ( 
.A(n_102),
.B(n_103),
.Y(n_112)
);

INVx4_ASAP7_75t_L g103 ( 
.A(n_84),
.Y(n_103)
);

AOI22xp5_ASAP7_75t_L g104 ( 
.A1(n_74),
.A2(n_57),
.B1(n_35),
.B2(n_38),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_L g113 ( 
.A(n_104),
.B(n_105),
.Y(n_113)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_65),
.Y(n_105)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_91),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_SL g132 ( 
.A(n_109),
.B(n_114),
.Y(n_132)
);

NOR4xp25_ASAP7_75t_L g110 ( 
.A(n_86),
.B(n_69),
.C(n_85),
.D(n_26),
.Y(n_110)
);

MAJx2_ASAP7_75t_L g136 ( 
.A(n_110),
.B(n_100),
.C(n_94),
.Y(n_136)
);

XOR2xp5_ASAP7_75t_L g111 ( 
.A(n_101),
.B(n_77),
.Y(n_111)
);

XOR2xp5_ASAP7_75t_L g143 ( 
.A(n_111),
.B(n_98),
.Y(n_143)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_97),
.Y(n_114)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_93),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_L g141 ( 
.A(n_115),
.B(n_118),
.Y(n_141)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_104),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_L g119 ( 
.A(n_88),
.B(n_94),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_SL g144 ( 
.A(n_119),
.B(n_124),
.Y(n_144)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_96),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_L g135 ( 
.A(n_120),
.B(n_121),
.Y(n_135)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_105),
.Y(n_121)
);

CKINVDCx16_ASAP7_75t_R g122 ( 
.A(n_103),
.Y(n_122)
);

CKINVDCx16_ASAP7_75t_R g133 ( 
.A(n_122),
.Y(n_133)
);

CKINVDCx16_ASAP7_75t_R g124 ( 
.A(n_106),
.Y(n_124)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_95),
.Y(n_125)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_125),
.Y(n_128)
);

OAI21xp5_ASAP7_75t_SL g130 ( 
.A1(n_126),
.A2(n_123),
.B(n_108),
.Y(n_130)
);

CKINVDCx20_ASAP7_75t_R g127 ( 
.A(n_112),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_SL g151 ( 
.A(n_127),
.B(n_140),
.Y(n_151)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_113),
.Y(n_129)
);

OAI21xp5_ASAP7_75t_SL g155 ( 
.A1(n_129),
.A2(n_130),
.B(n_134),
.Y(n_155)
);

OAI22xp5_ASAP7_75t_L g131 ( 
.A1(n_118),
.A2(n_90),
.B1(n_87),
.B2(n_89),
.Y(n_131)
);

AOI22xp5_ASAP7_75t_L g147 ( 
.A1(n_131),
.A2(n_114),
.B1(n_109),
.B2(n_98),
.Y(n_147)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_121),
.Y(n_134)
);

XNOR2xp5_ASAP7_75t_L g156 ( 
.A(n_136),
.B(n_142),
.Y(n_156)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_116),
.Y(n_137)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_137),
.Y(n_148)
);

MAJIxp5_ASAP7_75t_L g138 ( 
.A(n_108),
.B(n_107),
.C(n_95),
.Y(n_138)
);

MAJIxp5_ASAP7_75t_L g145 ( 
.A(n_138),
.B(n_143),
.C(n_111),
.Y(n_145)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_116),
.Y(n_139)
);

AOI21xp5_ASAP7_75t_L g152 ( 
.A1(n_139),
.A2(n_1),
.B(n_2),
.Y(n_152)
);

CKINVDCx20_ASAP7_75t_R g140 ( 
.A(n_117),
.Y(n_140)
);

AOI22xp5_ASAP7_75t_SL g142 ( 
.A1(n_115),
.A2(n_98),
.B1(n_107),
.B2(n_67),
.Y(n_142)
);

MAJIxp5_ASAP7_75t_L g165 ( 
.A(n_145),
.B(n_146),
.C(n_129),
.Y(n_165)
);

MAJIxp5_ASAP7_75t_L g146 ( 
.A(n_143),
.B(n_108),
.C(n_120),
.Y(n_146)
);

OAI22xp5_ASAP7_75t_SL g168 ( 
.A1(n_147),
.A2(n_153),
.B1(n_142),
.B2(n_134),
.Y(n_168)
);

OAI322xp33_ASAP7_75t_L g149 ( 
.A1(n_136),
.A2(n_98),
.A3(n_26),
.B1(n_16),
.B2(n_125),
.C1(n_15),
.C2(n_14),
.Y(n_149)
);

AOI321xp33_ASAP7_75t_L g159 ( 
.A1(n_149),
.A2(n_157),
.A3(n_158),
.B1(n_155),
.B2(n_61),
.C(n_4),
.Y(n_159)
);

OAI21xp5_ASAP7_75t_L g150 ( 
.A1(n_141),
.A2(n_57),
.B(n_83),
.Y(n_150)
);

OAI21xp5_ASAP7_75t_L g162 ( 
.A1(n_150),
.A2(n_152),
.B(n_154),
.Y(n_162)
);

OAI22xp5_ASAP7_75t_SL g153 ( 
.A1(n_141),
.A2(n_75),
.B1(n_106),
.B2(n_82),
.Y(n_153)
);

AOI21xp5_ASAP7_75t_SL g154 ( 
.A1(n_137),
.A2(n_26),
.B(n_2),
.Y(n_154)
);

A2O1A1O1Ixp25_ASAP7_75t_L g157 ( 
.A1(n_138),
.A2(n_26),
.B(n_11),
.C(n_13),
.D(n_12),
.Y(n_157)
);

OAI21x1_ASAP7_75t_L g158 ( 
.A1(n_130),
.A2(n_12),
.B(n_9),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_SL g174 ( 
.A(n_159),
.B(n_163),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_L g160 ( 
.A(n_148),
.B(n_135),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_L g172 ( 
.A(n_160),
.B(n_161),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_L g161 ( 
.A(n_150),
.B(n_139),
.Y(n_161)
);

CKINVDCx20_ASAP7_75t_R g163 ( 
.A(n_151),
.Y(n_163)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_153),
.Y(n_164)
);

NOR2xp33_ASAP7_75t_L g176 ( 
.A(n_164),
.B(n_166),
.Y(n_176)
);

XOR2xp5_ASAP7_75t_L g171 ( 
.A(n_165),
.B(n_145),
.Y(n_171)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_147),
.Y(n_166)
);

NOR2xp33_ASAP7_75t_SL g167 ( 
.A(n_154),
.B(n_132),
.Y(n_167)
);

AOI21xp5_ASAP7_75t_L g170 ( 
.A1(n_167),
.A2(n_169),
.B(n_156),
.Y(n_170)
);

AOI22xp5_ASAP7_75t_SL g177 ( 
.A1(n_168),
.A2(n_35),
.B1(n_37),
.B2(n_4),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_SL g169 ( 
.A(n_146),
.B(n_144),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_L g179 ( 
.A(n_170),
.B(n_173),
.Y(n_179)
);

MAJIxp5_ASAP7_75t_L g180 ( 
.A(n_171),
.B(n_175),
.C(n_160),
.Y(n_180)
);

OAI22xp5_ASAP7_75t_SL g173 ( 
.A1(n_161),
.A2(n_156),
.B1(n_128),
.B2(n_157),
.Y(n_173)
);

MAJIxp5_ASAP7_75t_L g175 ( 
.A(n_165),
.B(n_128),
.C(n_133),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_SL g178 ( 
.A(n_177),
.B(n_162),
.Y(n_178)
);

AOI21xp5_ASAP7_75t_L g188 ( 
.A1(n_178),
.A2(n_182),
.B(n_183),
.Y(n_188)
);

AND2x2_ASAP7_75t_L g185 ( 
.A(n_180),
.B(n_171),
.Y(n_185)
);

NOR2xp33_ASAP7_75t_SL g181 ( 
.A(n_174),
.B(n_162),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_L g187 ( 
.A(n_181),
.B(n_176),
.Y(n_187)
);

OAI21xp5_ASAP7_75t_SL g182 ( 
.A1(n_172),
.A2(n_159),
.B(n_168),
.Y(n_182)
);

OAI21xp5_ASAP7_75t_L g183 ( 
.A1(n_175),
.A2(n_1),
.B(n_3),
.Y(n_183)
);

OAI21xp5_ASAP7_75t_SL g184 ( 
.A1(n_177),
.A2(n_1),
.B(n_3),
.Y(n_184)
);

AOI21xp5_ASAP7_75t_L g189 ( 
.A1(n_184),
.A2(n_5),
.B(n_6),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_SL g192 ( 
.A(n_185),
.B(n_186),
.Y(n_192)
);

NOR2xp33_ASAP7_75t_SL g186 ( 
.A(n_179),
.B(n_173),
.Y(n_186)
);

OAI321xp33_ASAP7_75t_L g190 ( 
.A1(n_187),
.A2(n_189),
.A3(n_178),
.B1(n_7),
.B2(n_5),
.C(n_61),
.Y(n_190)
);

OAI21xp5_ASAP7_75t_SL g193 ( 
.A1(n_190),
.A2(n_61),
.B(n_5),
.Y(n_193)
);

BUFx24_ASAP7_75t_SL g191 ( 
.A(n_188),
.Y(n_191)
);

MAJIxp5_ASAP7_75t_L g194 ( 
.A(n_191),
.B(n_37),
.C(n_192),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_L g195 ( 
.A(n_193),
.B(n_194),
.Y(n_195)
);

NOR2xp33_ASAP7_75t_L g196 ( 
.A(n_195),
.B(n_37),
.Y(n_196)
);


endmodule