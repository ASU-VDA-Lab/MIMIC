module fake_jpeg_16759_n_318 (n_13, n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_318);

input n_13;
input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_318;

wire n_253;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_15;
wire n_141;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_14;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

BUFx12_ASAP7_75t_L g14 ( 
.A(n_1),
.Y(n_14)
);

BUFx6f_ASAP7_75t_L g15 ( 
.A(n_12),
.Y(n_15)
);

INVx2_ASAP7_75t_L g16 ( 
.A(n_13),
.Y(n_16)
);

BUFx12f_ASAP7_75t_L g17 ( 
.A(n_7),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_4),
.Y(n_18)
);

INVx5_ASAP7_75t_L g19 ( 
.A(n_6),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_3),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_12),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_10),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_13),
.Y(n_23)
);

INVx3_ASAP7_75t_L g24 ( 
.A(n_10),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_3),
.Y(n_25)
);

INVx6_ASAP7_75t_L g26 ( 
.A(n_9),
.Y(n_26)
);

INVx11_ASAP7_75t_L g27 ( 
.A(n_12),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_3),
.Y(n_28)
);

BUFx3_ASAP7_75t_L g29 ( 
.A(n_11),
.Y(n_29)
);

INVx2_ASAP7_75t_L g30 ( 
.A(n_14),
.Y(n_30)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_30),
.Y(n_57)
);

INVx6_ASAP7_75t_L g31 ( 
.A(n_17),
.Y(n_31)
);

INVx8_ASAP7_75t_L g48 ( 
.A(n_31),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_25),
.Y(n_32)
);

INVx2_ASAP7_75t_L g44 ( 
.A(n_32),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_25),
.Y(n_33)
);

INVx2_ASAP7_75t_L g55 ( 
.A(n_33),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g34 ( 
.A(n_16),
.B(n_18),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_L g45 ( 
.A(n_34),
.B(n_35),
.Y(n_45)
);

INVx4_ASAP7_75t_L g35 ( 
.A(n_17),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_25),
.Y(n_36)
);

INVx3_ASAP7_75t_L g43 ( 
.A(n_36),
.Y(n_43)
);

BUFx12f_ASAP7_75t_L g37 ( 
.A(n_17),
.Y(n_37)
);

BUFx4f_ASAP7_75t_SL g46 ( 
.A(n_37),
.Y(n_46)
);

BUFx12f_ASAP7_75t_L g38 ( 
.A(n_17),
.Y(n_38)
);

INVx5_ASAP7_75t_L g40 ( 
.A(n_38),
.Y(n_40)
);

BUFx12f_ASAP7_75t_L g39 ( 
.A(n_17),
.Y(n_39)
);

INVx8_ASAP7_75t_L g49 ( 
.A(n_39),
.Y(n_49)
);

INVx6_ASAP7_75t_SL g41 ( 
.A(n_37),
.Y(n_41)
);

INVx4_ASAP7_75t_SL g72 ( 
.A(n_41),
.Y(n_72)
);

INVx11_ASAP7_75t_L g42 ( 
.A(n_32),
.Y(n_42)
);

BUFx24_ASAP7_75t_L g68 ( 
.A(n_42),
.Y(n_68)
);

AND2x2_ASAP7_75t_L g47 ( 
.A(n_37),
.B(n_0),
.Y(n_47)
);

AOI21xp5_ASAP7_75t_L g60 ( 
.A1(n_47),
.A2(n_51),
.B(n_19),
.Y(n_60)
);

INVx3_ASAP7_75t_L g50 ( 
.A(n_30),
.Y(n_50)
);

INVx3_ASAP7_75t_L g76 ( 
.A(n_50),
.Y(n_76)
);

AND2x2_ASAP7_75t_L g51 ( 
.A(n_37),
.B(n_0),
.Y(n_51)
);

INVx2_ASAP7_75t_SL g52 ( 
.A(n_37),
.Y(n_52)
);

INVx2_ASAP7_75t_L g62 ( 
.A(n_52),
.Y(n_62)
);

AOI22xp33_ASAP7_75t_SL g53 ( 
.A1(n_31),
.A2(n_26),
.B1(n_16),
.B2(n_27),
.Y(n_53)
);

AOI22xp33_ASAP7_75t_SL g67 ( 
.A1(n_53),
.A2(n_26),
.B1(n_27),
.B2(n_19),
.Y(n_67)
);

OAI22xp5_ASAP7_75t_L g54 ( 
.A1(n_34),
.A2(n_26),
.B1(n_16),
.B2(n_24),
.Y(n_54)
);

AOI22xp5_ASAP7_75t_L g73 ( 
.A1(n_54),
.A2(n_26),
.B1(n_24),
.B2(n_19),
.Y(n_73)
);

INVx2_ASAP7_75t_SL g56 ( 
.A(n_37),
.Y(n_56)
);

INVx2_ASAP7_75t_L g63 ( 
.A(n_56),
.Y(n_63)
);

INVx3_ASAP7_75t_L g58 ( 
.A(n_30),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_L g75 ( 
.A(n_58),
.B(n_17),
.Y(n_75)
);

BUFx12_ASAP7_75t_L g59 ( 
.A(n_38),
.Y(n_59)
);

INVx2_ASAP7_75t_L g77 ( 
.A(n_59),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_SL g101 ( 
.A(n_60),
.B(n_71),
.Y(n_101)
);

INVx1_ASAP7_75t_SL g61 ( 
.A(n_47),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_61),
.B(n_64),
.Y(n_93)
);

CKINVDCx16_ASAP7_75t_R g64 ( 
.A(n_57),
.Y(n_64)
);

INVx2_ASAP7_75t_L g65 ( 
.A(n_57),
.Y(n_65)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_65),
.Y(n_87)
);

INVx4_ASAP7_75t_L g66 ( 
.A(n_48),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_66),
.B(n_81),
.Y(n_95)
);

AOI22xp5_ASAP7_75t_SL g104 ( 
.A1(n_67),
.A2(n_69),
.B1(n_22),
.B2(n_21),
.Y(n_104)
);

AND2x2_ASAP7_75t_L g69 ( 
.A(n_54),
.B(n_0),
.Y(n_69)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_44),
.Y(n_70)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_70),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_SL g71 ( 
.A(n_45),
.B(n_21),
.Y(n_71)
);

OAI22xp5_ASAP7_75t_SL g102 ( 
.A1(n_73),
.A2(n_74),
.B1(n_78),
.B2(n_42),
.Y(n_102)
);

AOI22xp5_ASAP7_75t_L g74 ( 
.A1(n_47),
.A2(n_24),
.B1(n_31),
.B2(n_35),
.Y(n_74)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_75),
.Y(n_90)
);

OAI22xp5_ASAP7_75t_SL g78 ( 
.A1(n_45),
.A2(n_31),
.B1(n_27),
.B2(n_35),
.Y(n_78)
);

INVx2_ASAP7_75t_L g79 ( 
.A(n_44),
.Y(n_79)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_79),
.Y(n_105)
);

INVx2_ASAP7_75t_L g80 ( 
.A(n_55),
.Y(n_80)
);

INVx3_ASAP7_75t_L g86 ( 
.A(n_80),
.Y(n_86)
);

CKINVDCx16_ASAP7_75t_R g81 ( 
.A(n_47),
.Y(n_81)
);

BUFx12_ASAP7_75t_L g82 ( 
.A(n_46),
.Y(n_82)
);

INVxp67_ASAP7_75t_L g85 ( 
.A(n_82),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_SL g83 ( 
.A(n_69),
.B(n_51),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g115 ( 
.A(n_83),
.B(n_89),
.Y(n_115)
);

AOI22xp33_ASAP7_75t_SL g84 ( 
.A1(n_66),
.A2(n_40),
.B1(n_41),
.B2(n_49),
.Y(n_84)
);

AOI21xp5_ASAP7_75t_L g109 ( 
.A1(n_84),
.A2(n_68),
.B(n_40),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_61),
.B(n_51),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_SL g91 ( 
.A(n_69),
.B(n_51),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_SL g108 ( 
.A(n_91),
.B(n_92),
.Y(n_108)
);

FAx1_ASAP7_75t_SL g92 ( 
.A(n_74),
.B(n_50),
.CI(n_58),
.CON(n_92),
.SN(n_92)
);

NAND2xp5_ASAP7_75t_SL g94 ( 
.A(n_78),
.B(n_50),
.Y(n_94)
);

OAI21xp5_ASAP7_75t_L g126 ( 
.A1(n_94),
.A2(n_103),
.B(n_32),
.Y(n_126)
);

INVx8_ASAP7_75t_L g96 ( 
.A(n_76),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g122 ( 
.A(n_96),
.B(n_97),
.Y(n_122)
);

CKINVDCx16_ASAP7_75t_R g97 ( 
.A(n_60),
.Y(n_97)
);

A2O1A1Ixp33_ASAP7_75t_L g98 ( 
.A1(n_73),
.A2(n_20),
.B(n_18),
.C(n_21),
.Y(n_98)
);

OAI31xp33_ASAP7_75t_L g117 ( 
.A1(n_98),
.A2(n_22),
.A3(n_101),
.B(n_104),
.Y(n_117)
);

INVx3_ASAP7_75t_L g99 ( 
.A(n_76),
.Y(n_99)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_99),
.Y(n_107)
);

INVxp67_ASAP7_75t_L g100 ( 
.A(n_77),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g123 ( 
.A(n_100),
.B(n_106),
.Y(n_123)
);

AOI22xp5_ASAP7_75t_L g113 ( 
.A1(n_102),
.A2(n_43),
.B1(n_55),
.B2(n_79),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_SL g103 ( 
.A(n_65),
.B(n_48),
.Y(n_103)
);

AND2x2_ASAP7_75t_L g111 ( 
.A(n_104),
.B(n_22),
.Y(n_111)
);

CKINVDCx16_ASAP7_75t_R g106 ( 
.A(n_72),
.Y(n_106)
);

OAI21xp5_ASAP7_75t_L g140 ( 
.A1(n_109),
.A2(n_111),
.B(n_112),
.Y(n_140)
);

BUFx3_ASAP7_75t_L g110 ( 
.A(n_85),
.Y(n_110)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_110),
.Y(n_156)
);

AND2x2_ASAP7_75t_L g112 ( 
.A(n_89),
.B(n_0),
.Y(n_112)
);

OAI22xp5_ASAP7_75t_L g144 ( 
.A1(n_113),
.A2(n_114),
.B1(n_116),
.B2(n_121),
.Y(n_144)
);

OAI22xp5_ASAP7_75t_SL g114 ( 
.A1(n_97),
.A2(n_42),
.B1(n_43),
.B2(n_48),
.Y(n_114)
);

OAI22xp5_ASAP7_75t_L g116 ( 
.A1(n_94),
.A2(n_43),
.B1(n_80),
.B2(n_70),
.Y(n_116)
);

OAI21x1_ASAP7_75t_L g153 ( 
.A1(n_117),
.A2(n_98),
.B(n_84),
.Y(n_153)
);

OR2x2_ASAP7_75t_L g118 ( 
.A(n_92),
.B(n_63),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_L g133 ( 
.A(n_118),
.B(n_126),
.Y(n_133)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_103),
.Y(n_119)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_119),
.Y(n_132)
);

AOI21xp5_ASAP7_75t_L g120 ( 
.A1(n_95),
.A2(n_40),
.B(n_68),
.Y(n_120)
);

INVxp67_ASAP7_75t_L g146 ( 
.A(n_120),
.Y(n_146)
);

OAI22xp5_ASAP7_75t_L g121 ( 
.A1(n_90),
.A2(n_49),
.B1(n_72),
.B2(n_62),
.Y(n_121)
);

CKINVDCx20_ASAP7_75t_R g124 ( 
.A(n_88),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_SL g148 ( 
.A(n_124),
.B(n_87),
.Y(n_148)
);

BUFx2_ASAP7_75t_L g125 ( 
.A(n_99),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_L g141 ( 
.A(n_125),
.B(n_96),
.Y(n_141)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_86),
.Y(n_127)
);

INVx2_ASAP7_75t_L g135 ( 
.A(n_127),
.Y(n_135)
);

AOI22xp5_ASAP7_75t_L g128 ( 
.A1(n_95),
.A2(n_63),
.B1(n_62),
.B2(n_36),
.Y(n_128)
);

OAI22xp5_ASAP7_75t_L g150 ( 
.A1(n_128),
.A2(n_131),
.B1(n_96),
.B2(n_99),
.Y(n_150)
);

MAJIxp5_ASAP7_75t_L g129 ( 
.A(n_93),
.B(n_46),
.C(n_38),
.Y(n_129)
);

MAJIxp5_ASAP7_75t_L g142 ( 
.A(n_129),
.B(n_130),
.C(n_92),
.Y(n_142)
);

OAI21xp5_ASAP7_75t_L g130 ( 
.A1(n_83),
.A2(n_91),
.B(n_101),
.Y(n_130)
);

OAI22xp5_ASAP7_75t_SL g131 ( 
.A1(n_102),
.A2(n_36),
.B1(n_32),
.B2(n_33),
.Y(n_131)
);

BUFx3_ASAP7_75t_L g134 ( 
.A(n_110),
.Y(n_134)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_134),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_L g136 ( 
.A(n_118),
.B(n_90),
.Y(n_136)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_136),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_L g137 ( 
.A(n_118),
.B(n_93),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_L g171 ( 
.A(n_137),
.B(n_149),
.Y(n_171)
);

INVx3_ASAP7_75t_L g138 ( 
.A(n_125),
.Y(n_138)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_138),
.Y(n_182)
);

BUFx2_ASAP7_75t_L g139 ( 
.A(n_125),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_L g163 ( 
.A(n_139),
.B(n_151),
.Y(n_163)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_141),
.Y(n_185)
);

XNOR2xp5_ASAP7_75t_L g176 ( 
.A(n_142),
.B(n_143),
.Y(n_176)
);

MAJx2_ASAP7_75t_L g143 ( 
.A(n_130),
.B(n_108),
.C(n_115),
.Y(n_143)
);

NOR2xp33_ASAP7_75t_L g145 ( 
.A(n_121),
.B(n_107),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_SL g167 ( 
.A(n_145),
.B(n_148),
.Y(n_167)
);

BUFx12f_ASAP7_75t_SL g147 ( 
.A(n_117),
.Y(n_147)
);

AOI22xp5_ASAP7_75t_SL g159 ( 
.A1(n_147),
.A2(n_155),
.B1(n_111),
.B2(n_124),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_L g149 ( 
.A(n_108),
.B(n_92),
.Y(n_149)
);

AOI22xp5_ASAP7_75t_L g160 ( 
.A1(n_150),
.A2(n_116),
.B1(n_122),
.B2(n_119),
.Y(n_160)
);

INVx5_ASAP7_75t_L g151 ( 
.A(n_110),
.Y(n_151)
);

INVxp33_ASAP7_75t_L g152 ( 
.A(n_123),
.Y(n_152)
);

INVx1_ASAP7_75t_SL g170 ( 
.A(n_152),
.Y(n_170)
);

OAI21xp5_ASAP7_75t_L g161 ( 
.A1(n_153),
.A2(n_109),
.B(n_120),
.Y(n_161)
);

AND2x6_ASAP7_75t_L g154 ( 
.A(n_111),
.B(n_106),
.Y(n_154)
);

CKINVDCx20_ASAP7_75t_R g168 ( 
.A(n_154),
.Y(n_168)
);

INVx5_ASAP7_75t_L g155 ( 
.A(n_107),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_L g157 ( 
.A(n_123),
.B(n_86),
.Y(n_157)
);

CKINVDCx20_ASAP7_75t_R g183 ( 
.A(n_157),
.Y(n_183)
);

MAJIxp5_ASAP7_75t_L g158 ( 
.A(n_142),
.B(n_115),
.C(n_129),
.Y(n_158)
);

MAJIxp5_ASAP7_75t_L g190 ( 
.A(n_158),
.B(n_162),
.C(n_156),
.Y(n_190)
);

OAI21xp5_ASAP7_75t_L g201 ( 
.A1(n_159),
.A2(n_161),
.B(n_175),
.Y(n_201)
);

OAI22xp5_ASAP7_75t_L g208 ( 
.A1(n_160),
.A2(n_165),
.B1(n_180),
.B2(n_184),
.Y(n_208)
);

XOR2xp5_ASAP7_75t_L g162 ( 
.A(n_149),
.B(n_122),
.Y(n_162)
);

AND2x2_ASAP7_75t_L g164 ( 
.A(n_133),
.B(n_128),
.Y(n_164)
);

OAI21xp5_ASAP7_75t_SL g188 ( 
.A1(n_164),
.A2(n_169),
.B(n_178),
.Y(n_188)
);

AOI22xp5_ASAP7_75t_L g165 ( 
.A1(n_147),
.A2(n_112),
.B1(n_113),
.B2(n_131),
.Y(n_165)
);

AO21x2_ASAP7_75t_L g166 ( 
.A1(n_152),
.A2(n_114),
.B(n_126),
.Y(n_166)
);

AOI22xp5_ASAP7_75t_L g186 ( 
.A1(n_166),
.A2(n_155),
.B1(n_138),
.B2(n_135),
.Y(n_186)
);

AOI21xp5_ASAP7_75t_L g169 ( 
.A1(n_146),
.A2(n_112),
.B(n_127),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_L g173 ( 
.A(n_136),
.B(n_87),
.Y(n_173)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_173),
.Y(n_209)
);

NAND2xp5_ASAP7_75t_L g174 ( 
.A(n_132),
.B(n_98),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_L g199 ( 
.A(n_174),
.B(n_179),
.Y(n_199)
);

OAI21xp5_ASAP7_75t_L g175 ( 
.A1(n_133),
.A2(n_20),
.B(n_18),
.Y(n_175)
);

OAI21xp5_ASAP7_75t_L g177 ( 
.A1(n_140),
.A2(n_20),
.B(n_105),
.Y(n_177)
);

OAI21xp5_ASAP7_75t_L g203 ( 
.A1(n_177),
.A2(n_1),
.B(n_2),
.Y(n_203)
);

AOI21xp5_ASAP7_75t_L g178 ( 
.A1(n_146),
.A2(n_86),
.B(n_88),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_L g179 ( 
.A(n_132),
.B(n_105),
.Y(n_179)
);

AOI22xp5_ASAP7_75t_L g180 ( 
.A1(n_144),
.A2(n_49),
.B1(n_52),
.B2(n_56),
.Y(n_180)
);

OAI22xp5_ASAP7_75t_SL g184 ( 
.A1(n_137),
.A2(n_56),
.B1(n_52),
.B2(n_36),
.Y(n_184)
);

OAI22xp5_ASAP7_75t_SL g232 ( 
.A1(n_186),
.A2(n_187),
.B1(n_204),
.B2(n_175),
.Y(n_232)
);

AOI22xp5_ASAP7_75t_L g187 ( 
.A1(n_164),
.A2(n_154),
.B1(n_143),
.B2(n_140),
.Y(n_187)
);

XNOR2xp5_ASAP7_75t_SL g189 ( 
.A(n_176),
.B(n_158),
.Y(n_189)
);

XOR2xp5_ASAP7_75t_L g212 ( 
.A(n_189),
.B(n_207),
.Y(n_212)
);

MAJIxp5_ASAP7_75t_L g216 ( 
.A(n_190),
.B(n_191),
.C(n_194),
.Y(n_216)
);

XNOR2xp5_ASAP7_75t_L g191 ( 
.A(n_176),
.B(n_135),
.Y(n_191)
);

INVxp67_ASAP7_75t_L g192 ( 
.A(n_163),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_L g215 ( 
.A(n_192),
.B(n_196),
.Y(n_215)
);

NOR2xp33_ASAP7_75t_L g193 ( 
.A(n_181),
.B(n_134),
.Y(n_193)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_193),
.Y(n_219)
);

MAJIxp5_ASAP7_75t_L g194 ( 
.A(n_162),
.B(n_46),
.C(n_38),
.Y(n_194)
);

MAJIxp5_ASAP7_75t_L g195 ( 
.A(n_173),
.B(n_46),
.C(n_38),
.Y(n_195)
);

MAJIxp5_ASAP7_75t_L g217 ( 
.A(n_195),
.B(n_194),
.C(n_191),
.Y(n_217)
);

INVx5_ASAP7_75t_L g196 ( 
.A(n_166),
.Y(n_196)
);

NAND3xp33_ASAP7_75t_L g197 ( 
.A(n_168),
.B(n_151),
.C(n_13),
.Y(n_197)
);

NOR2xp33_ASAP7_75t_SL g221 ( 
.A(n_197),
.B(n_159),
.Y(n_221)
);

BUFx3_ASAP7_75t_L g198 ( 
.A(n_166),
.Y(n_198)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_198),
.Y(n_220)
);

CKINVDCx20_ASAP7_75t_R g200 ( 
.A(n_179),
.Y(n_200)
);

NAND2xp5_ASAP7_75t_SL g227 ( 
.A(n_200),
.B(n_203),
.Y(n_227)
);

NAND2xp5_ASAP7_75t_L g202 ( 
.A(n_183),
.B(n_11),
.Y(n_202)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_202),
.Y(n_225)
);

AOI22xp5_ASAP7_75t_L g204 ( 
.A1(n_164),
.A2(n_139),
.B1(n_56),
.B2(n_52),
.Y(n_204)
);

NAND2xp5_ASAP7_75t_L g205 ( 
.A(n_167),
.B(n_11),
.Y(n_205)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_205),
.Y(n_228)
);

AOI21xp33_ASAP7_75t_SL g206 ( 
.A1(n_166),
.A2(n_82),
.B(n_59),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_SL g233 ( 
.A(n_206),
.B(n_182),
.Y(n_233)
);

XOR2xp5_ASAP7_75t_L g207 ( 
.A(n_171),
.B(n_82),
.Y(n_207)
);

AOI21xp5_ASAP7_75t_L g210 ( 
.A1(n_161),
.A2(n_68),
.B(n_2),
.Y(n_210)
);

OAI22xp5_ASAP7_75t_L g213 ( 
.A1(n_210),
.A2(n_177),
.B1(n_174),
.B2(n_169),
.Y(n_213)
);

NAND2xp5_ASAP7_75t_L g211 ( 
.A(n_185),
.B(n_10),
.Y(n_211)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_211),
.Y(n_230)
);

AOI22xp5_ASAP7_75t_L g250 ( 
.A1(n_213),
.A2(n_9),
.B1(n_2),
.B2(n_3),
.Y(n_250)
);

XOR2xp5_ASAP7_75t_L g214 ( 
.A(n_189),
.B(n_171),
.Y(n_214)
);

XOR2xp5_ASAP7_75t_L g236 ( 
.A(n_214),
.B(n_224),
.Y(n_236)
);

MAJIxp5_ASAP7_75t_L g237 ( 
.A(n_217),
.B(n_226),
.C(n_231),
.Y(n_237)
);

AND2x2_ASAP7_75t_L g218 ( 
.A(n_186),
.B(n_204),
.Y(n_218)
);

INVx1_ASAP7_75t_SL g242 ( 
.A(n_218),
.Y(n_242)
);

NOR2xp33_ASAP7_75t_L g234 ( 
.A(n_221),
.B(n_201),
.Y(n_234)
);

AOI22xp5_ASAP7_75t_L g222 ( 
.A1(n_196),
.A2(n_166),
.B1(n_172),
.B2(n_170),
.Y(n_222)
);

OAI22xp5_ASAP7_75t_L g238 ( 
.A1(n_222),
.A2(n_229),
.B1(n_201),
.B2(n_210),
.Y(n_238)
);

NOR2xp33_ASAP7_75t_SL g223 ( 
.A(n_209),
.B(n_172),
.Y(n_223)
);

NAND2xp5_ASAP7_75t_L g240 ( 
.A(n_223),
.B(n_199),
.Y(n_240)
);

XOR2xp5_ASAP7_75t_L g224 ( 
.A(n_187),
.B(n_178),
.Y(n_224)
);

MAJIxp5_ASAP7_75t_L g226 ( 
.A(n_190),
.B(n_207),
.C(n_195),
.Y(n_226)
);

AOI22xp5_ASAP7_75t_L g229 ( 
.A1(n_208),
.A2(n_170),
.B1(n_160),
.B2(n_165),
.Y(n_229)
);

MAJIxp5_ASAP7_75t_L g231 ( 
.A(n_188),
.B(n_184),
.C(n_180),
.Y(n_231)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_232),
.Y(n_235)
);

OAI22xp5_ASAP7_75t_SL g245 ( 
.A1(n_233),
.A2(n_227),
.B1(n_231),
.B2(n_230),
.Y(n_245)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_234),
.Y(n_255)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_238),
.Y(n_259)
);

XNOR2xp5_ASAP7_75t_L g239 ( 
.A(n_216),
.B(n_188),
.Y(n_239)
);

MAJIxp5_ASAP7_75t_L g262 ( 
.A(n_239),
.B(n_248),
.C(n_252),
.Y(n_262)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_240),
.Y(n_260)
);

XOR2xp5_ASAP7_75t_L g241 ( 
.A(n_212),
.B(n_199),
.Y(n_241)
);

XOR2xp5_ASAP7_75t_L g254 ( 
.A(n_241),
.B(n_253),
.Y(n_254)
);

OAI21xp5_ASAP7_75t_L g243 ( 
.A1(n_226),
.A2(n_192),
.B(n_203),
.Y(n_243)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_243),
.Y(n_265)
);

XOR2xp5_ASAP7_75t_L g244 ( 
.A(n_212),
.B(n_198),
.Y(n_244)
);

XOR2xp5_ASAP7_75t_L g270 ( 
.A(n_244),
.B(n_39),
.Y(n_270)
);

NOR2xp33_ASAP7_75t_L g264 ( 
.A(n_245),
.B(n_232),
.Y(n_264)
);

NAND2xp5_ASAP7_75t_L g246 ( 
.A(n_219),
.B(n_228),
.Y(n_246)
);

CKINVDCx20_ASAP7_75t_R g258 ( 
.A(n_246),
.Y(n_258)
);

NAND2xp5_ASAP7_75t_L g247 ( 
.A(n_225),
.B(n_215),
.Y(n_247)
);

NOR2xp33_ASAP7_75t_SL g256 ( 
.A(n_247),
.B(n_222),
.Y(n_256)
);

XNOR2xp5_ASAP7_75t_L g248 ( 
.A(n_216),
.B(n_59),
.Y(n_248)
);

OAI22xp5_ASAP7_75t_L g249 ( 
.A1(n_229),
.A2(n_23),
.B1(n_15),
.B2(n_9),
.Y(n_249)
);

OAI22xp5_ASAP7_75t_L g269 ( 
.A1(n_249),
.A2(n_250),
.B1(n_15),
.B2(n_23),
.Y(n_269)
);

OAI21xp5_ASAP7_75t_L g251 ( 
.A1(n_218),
.A2(n_1),
.B(n_2),
.Y(n_251)
);

NAND2xp5_ASAP7_75t_L g263 ( 
.A(n_251),
.B(n_1),
.Y(n_263)
);

MAJIxp5_ASAP7_75t_L g252 ( 
.A(n_217),
.B(n_39),
.C(n_38),
.Y(n_252)
);

XNOR2x1_ASAP7_75t_L g253 ( 
.A(n_224),
.B(n_59),
.Y(n_253)
);

NAND2xp5_ASAP7_75t_SL g274 ( 
.A(n_256),
.B(n_264),
.Y(n_274)
);

XOR2xp5_ASAP7_75t_L g257 ( 
.A(n_236),
.B(n_244),
.Y(n_257)
);

XOR2xp5_ASAP7_75t_L g272 ( 
.A(n_257),
.B(n_270),
.Y(n_272)
);

XNOR2xp5_ASAP7_75t_L g261 ( 
.A(n_237),
.B(n_214),
.Y(n_261)
);

MAJIxp5_ASAP7_75t_L g278 ( 
.A(n_261),
.B(n_268),
.C(n_39),
.Y(n_278)
);

NOR2xp33_ASAP7_75t_L g271 ( 
.A(n_263),
.B(n_269),
.Y(n_271)
);

OAI22xp5_ASAP7_75t_SL g266 ( 
.A1(n_235),
.A2(n_220),
.B1(n_218),
.B2(n_33),
.Y(n_266)
);

NAND2xp5_ASAP7_75t_SL g279 ( 
.A(n_266),
.B(n_267),
.Y(n_279)
);

AO221x1_ASAP7_75t_L g267 ( 
.A1(n_253),
.A2(n_251),
.B1(n_242),
.B2(n_239),
.C(n_241),
.Y(n_267)
);

MAJIxp5_ASAP7_75t_L g268 ( 
.A(n_237),
.B(n_248),
.C(n_236),
.Y(n_268)
);

XNOR2xp5_ASAP7_75t_L g273 ( 
.A(n_261),
.B(n_252),
.Y(n_273)
);

MAJIxp5_ASAP7_75t_L g295 ( 
.A(n_273),
.B(n_275),
.C(n_278),
.Y(n_295)
);

XNOR2xp5_ASAP7_75t_L g275 ( 
.A(n_262),
.B(n_242),
.Y(n_275)
);

NOR2xp33_ASAP7_75t_L g276 ( 
.A(n_255),
.B(n_15),
.Y(n_276)
);

CKINVDCx20_ASAP7_75t_R g289 ( 
.A(n_276),
.Y(n_289)
);

XNOR2xp5_ASAP7_75t_L g277 ( 
.A(n_268),
.B(n_29),
.Y(n_277)
);

NAND2xp5_ASAP7_75t_SL g291 ( 
.A(n_277),
.B(n_280),
.Y(n_291)
);

XNOR2xp5_ASAP7_75t_L g280 ( 
.A(n_262),
.B(n_270),
.Y(n_280)
);

OAI21xp5_ASAP7_75t_L g281 ( 
.A1(n_265),
.A2(n_15),
.B(n_23),
.Y(n_281)
);

AOI21xp5_ASAP7_75t_L g286 ( 
.A1(n_281),
.A2(n_282),
.B(n_263),
.Y(n_286)
);

OAI21xp5_ASAP7_75t_L g282 ( 
.A1(n_258),
.A2(n_23),
.B(n_29),
.Y(n_282)
);

XNOR2xp5_ASAP7_75t_L g283 ( 
.A(n_257),
.B(n_29),
.Y(n_283)
);

XNOR2xp5_ASAP7_75t_L g287 ( 
.A(n_283),
.B(n_254),
.Y(n_287)
);

NOR2xp33_ASAP7_75t_L g284 ( 
.A(n_260),
.B(n_28),
.Y(n_284)
);

NAND2xp5_ASAP7_75t_L g288 ( 
.A(n_284),
.B(n_271),
.Y(n_288)
);

NOR2xp33_ASAP7_75t_SL g285 ( 
.A(n_259),
.B(n_4),
.Y(n_285)
);

NAND2xp5_ASAP7_75t_SL g293 ( 
.A(n_285),
.B(n_4),
.Y(n_293)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_286),
.Y(n_300)
);

NAND2xp5_ASAP7_75t_SL g302 ( 
.A(n_287),
.B(n_293),
.Y(n_302)
);

CKINVDCx20_ASAP7_75t_R g303 ( 
.A(n_288),
.Y(n_303)
);

OAI21xp5_ASAP7_75t_L g290 ( 
.A1(n_279),
.A2(n_266),
.B(n_254),
.Y(n_290)
);

AOI21xp5_ASAP7_75t_L g305 ( 
.A1(n_290),
.A2(n_272),
.B(n_6),
.Y(n_305)
);

AOI322xp5_ASAP7_75t_L g292 ( 
.A1(n_274),
.A2(n_33),
.A3(n_28),
.B1(n_25),
.B2(n_39),
.C1(n_8),
.C2(n_4),
.Y(n_292)
);

OAI21x1_ASAP7_75t_L g299 ( 
.A1(n_292),
.A2(n_296),
.B(n_5),
.Y(n_299)
);

NAND2xp5_ASAP7_75t_L g294 ( 
.A(n_275),
.B(n_39),
.Y(n_294)
);

NOR2xp33_ASAP7_75t_L g301 ( 
.A(n_294),
.B(n_297),
.Y(n_301)
);

AOI322xp5_ASAP7_75t_L g296 ( 
.A1(n_283),
.A2(n_28),
.A3(n_6),
.B1(n_7),
.B2(n_8),
.C1(n_5),
.C2(n_14),
.Y(n_296)
);

AOI22xp5_ASAP7_75t_L g297 ( 
.A1(n_278),
.A2(n_5),
.B1(n_6),
.B2(n_7),
.Y(n_297)
);

OAI21xp5_ASAP7_75t_L g298 ( 
.A1(n_295),
.A2(n_273),
.B(n_272),
.Y(n_298)
);

NAND2xp5_ASAP7_75t_L g311 ( 
.A(n_298),
.B(n_14),
.Y(n_311)
);

OAI21x1_ASAP7_75t_L g307 ( 
.A1(n_299),
.A2(n_28),
.B(n_8),
.Y(n_307)
);

O2A1O1Ixp33_ASAP7_75t_SL g304 ( 
.A1(n_291),
.A2(n_290),
.B(n_289),
.C(n_297),
.Y(n_304)
);

OAI21xp5_ASAP7_75t_L g310 ( 
.A1(n_304),
.A2(n_305),
.B(n_306),
.Y(n_310)
);

AOI21xp5_ASAP7_75t_L g306 ( 
.A1(n_287),
.A2(n_5),
.B(n_7),
.Y(n_306)
);

NAND2xp5_ASAP7_75t_L g313 ( 
.A(n_307),
.B(n_308),
.Y(n_313)
);

A2O1A1Ixp33_ASAP7_75t_L g308 ( 
.A1(n_300),
.A2(n_295),
.B(n_8),
.C(n_14),
.Y(n_308)
);

INVxp67_ASAP7_75t_L g309 ( 
.A(n_302),
.Y(n_309)
);

XOR2xp5_ASAP7_75t_L g314 ( 
.A(n_309),
.B(n_311),
.Y(n_314)
);

NAND2xp5_ASAP7_75t_L g312 ( 
.A(n_303),
.B(n_14),
.Y(n_312)
);

MAJIxp5_ASAP7_75t_L g315 ( 
.A(n_312),
.B(n_301),
.C(n_14),
.Y(n_315)
);

NAND2xp5_ASAP7_75t_L g316 ( 
.A(n_315),
.B(n_310),
.Y(n_316)
);

OAI21xp5_ASAP7_75t_L g317 ( 
.A1(n_316),
.A2(n_313),
.B(n_314),
.Y(n_317)
);

XOR2xp5_ASAP7_75t_L g318 ( 
.A(n_317),
.B(n_314),
.Y(n_318)
);


endmodule