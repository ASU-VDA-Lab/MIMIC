module fake_netlist_5_91_n_2496 (n_137, n_676, n_294, n_431, n_318, n_380, n_419, n_653, n_611, n_444, n_642, n_469, n_615, n_82, n_194, n_316, n_389, n_549, n_684, n_418, n_248, n_124, n_86, n_136, n_146, n_315, n_268, n_523, n_451, n_532, n_705, n_619, n_408, n_61, n_678, n_664, n_376, n_697, n_503, n_127, n_75, n_235, n_226, n_605, n_74, n_667, n_515, n_57, n_353, n_351, n_367, n_620, n_643, n_452, n_397, n_493, n_111, n_525, n_703, n_698, n_483, n_544, n_683, n_155, n_649, n_552, n_547, n_43, n_721, n_116, n_22, n_467, n_564, n_423, n_284, n_46, n_245, n_21, n_501, n_725, n_139, n_38, n_105, n_280, n_590, n_629, n_672, n_4, n_378, n_551, n_17, n_581, n_688, n_382, n_554, n_254, n_690, n_33, n_23, n_583, n_671, n_718, n_302, n_265, n_526, n_719, n_293, n_372, n_443, n_244, n_677, n_47, n_173, n_198, n_714, n_447, n_247, n_314, n_368, n_433, n_604, n_8, n_321, n_292, n_625, n_621, n_100, n_455, n_674, n_417, n_612, n_212, n_385, n_498, n_516, n_507, n_119, n_497, n_689, n_738, n_606, n_559, n_275, n_640, n_252, n_624, n_26, n_295, n_133, n_330, n_508, n_739, n_506, n_2, n_737, n_610, n_692, n_6, n_509, n_568, n_39, n_147, n_373, n_67, n_307, n_633, n_439, n_87, n_150, n_530, n_556, n_106, n_209, n_259, n_448, n_668, n_733, n_375, n_301, n_576, n_68, n_93, n_186, n_537, n_134, n_191, n_587, n_659, n_51, n_63, n_492, n_563, n_171, n_153, n_524, n_399, n_341, n_204, n_394, n_250, n_579, n_548, n_543, n_260, n_298, n_650, n_320, n_694, n_518, n_505, n_286, n_122, n_282, n_331, n_10, n_24, n_406, n_519, n_470, n_325, n_449, n_132, n_90, n_724, n_546, n_101, n_658, n_281, n_240, n_381, n_189, n_220, n_291, n_231, n_257, n_390, n_731, n_31, n_456, n_13, n_371, n_481, n_535, n_709, n_152, n_540, n_317, n_618, n_9, n_323, n_569, n_195, n_42, n_356, n_227, n_592, n_45, n_271, n_94, n_335, n_123, n_654, n_370, n_167, n_234, n_343, n_308, n_379, n_428, n_267, n_514, n_457, n_570, n_297, n_156, n_5, n_603, n_225, n_377, n_484, n_219, n_442, n_157, n_131, n_192, n_636, n_600, n_660, n_223, n_392, n_158, n_655, n_704, n_138, n_264, n_109, n_669, n_472, n_454, n_387, n_374, n_163, n_276, n_339, n_95, n_183, n_185, n_243, n_398, n_396, n_635, n_347, n_169, n_59, n_522, n_550, n_255, n_696, n_215, n_350, n_196, n_662, n_459, n_646, n_211, n_218, n_400, n_181, n_436, n_3, n_290, n_580, n_221, n_178, n_622, n_723, n_386, n_578, n_287, n_344, n_555, n_473, n_422, n_475, n_72, n_661, n_104, n_41, n_682, n_415, n_56, n_141, n_485, n_496, n_355, n_486, n_670, n_15, n_336, n_584, n_681, n_591, n_145, n_48, n_521, n_614, n_663, n_50, n_337, n_430, n_313, n_631, n_673, n_88, n_479, n_528, n_510, n_216, n_680, n_168, n_395, n_164, n_432, n_553, n_727, n_311, n_208, n_142, n_214, n_328, n_140, n_299, n_303, n_369, n_675, n_296, n_613, n_241, n_637, n_357, n_598, n_685, n_608, n_184, n_446, n_445, n_65, n_78, n_144, n_114, n_96, n_691, n_717, n_165, n_468, n_499, n_213, n_129, n_342, n_482, n_517, n_98, n_588, n_361, n_464, n_363, n_402, n_413, n_734, n_638, n_700, n_197, n_107, n_573, n_69, n_236, n_388, n_1, n_249, n_740, n_304, n_329, n_203, n_274, n_577, n_384, n_582, n_460, n_80, n_35, n_73, n_277, n_92, n_19, n_338, n_149, n_477, n_461, n_333, n_571, n_693, n_309, n_30, n_512, n_14, n_84, n_462, n_130, n_322, n_567, n_258, n_652, n_29, n_79, n_151, n_25, n_306, n_722, n_458, n_288, n_188, n_190, n_201, n_263, n_471, n_609, n_44, n_224, n_40, n_34, n_228, n_283, n_383, n_711, n_474, n_112, n_542, n_85, n_463, n_488, n_595, n_736, n_502, n_239, n_466, n_420, n_630, n_489, n_632, n_699, n_55, n_617, n_49, n_310, n_54, n_593, n_504, n_511, n_12, n_586, n_465, n_76, n_358, n_362, n_170, n_332, n_27, n_77, n_102, n_161, n_273, n_349, n_585, n_270, n_616, n_230, n_81, n_118, n_601, n_279, n_70, n_253, n_261, n_174, n_289, n_627, n_172, n_206, n_217, n_440, n_726, n_478, n_545, n_441, n_450, n_648, n_312, n_476, n_429, n_534, n_345, n_210, n_494, n_641, n_628, n_365, n_91, n_729, n_730, n_176, n_557, n_182, n_143, n_83, n_354, n_575, n_607, n_480, n_647, n_237, n_425, n_513, n_407, n_527, n_679, n_707, n_710, n_695, n_180, n_560, n_656, n_340, n_207, n_561, n_37, n_346, n_393, n_229, n_108, n_487, n_495, n_602, n_665, n_574, n_437, n_66, n_177, n_60, n_403, n_453, n_421, n_16, n_720, n_0, n_58, n_623, n_405, n_18, n_359, n_490, n_117, n_326, n_233, n_404, n_686, n_205, n_366, n_572, n_113, n_712, n_246, n_596, n_179, n_125, n_410, n_558, n_708, n_269, n_529, n_128, n_735, n_702, n_285, n_412, n_120, n_232, n_327, n_135, n_657, n_126, n_644, n_728, n_202, n_266, n_272, n_491, n_427, n_732, n_193, n_251, n_352, n_53, n_160, n_565, n_426, n_520, n_566, n_409, n_589, n_716, n_597, n_500, n_562, n_154, n_62, n_148, n_71, n_300, n_651, n_435, n_159, n_334, n_599, n_541, n_391, n_701, n_434, n_645, n_539, n_175, n_538, n_666, n_262, n_238, n_639, n_99, n_687, n_715, n_411, n_414, n_319, n_364, n_20, n_536, n_531, n_121, n_242, n_360, n_36, n_594, n_200, n_162, n_64, n_222, n_28, n_89, n_438, n_115, n_713, n_324, n_634, n_416, n_199, n_187, n_32, n_401, n_103, n_348, n_97, n_166, n_626, n_11, n_424, n_7, n_706, n_256, n_305, n_533, n_52, n_278, n_110, n_2496);

input n_137;
input n_676;
input n_294;
input n_431;
input n_318;
input n_380;
input n_419;
input n_653;
input n_611;
input n_444;
input n_642;
input n_469;
input n_615;
input n_82;
input n_194;
input n_316;
input n_389;
input n_549;
input n_684;
input n_418;
input n_248;
input n_124;
input n_86;
input n_136;
input n_146;
input n_315;
input n_268;
input n_523;
input n_451;
input n_532;
input n_705;
input n_619;
input n_408;
input n_61;
input n_678;
input n_664;
input n_376;
input n_697;
input n_503;
input n_127;
input n_75;
input n_235;
input n_226;
input n_605;
input n_74;
input n_667;
input n_515;
input n_57;
input n_353;
input n_351;
input n_367;
input n_620;
input n_643;
input n_452;
input n_397;
input n_493;
input n_111;
input n_525;
input n_703;
input n_698;
input n_483;
input n_544;
input n_683;
input n_155;
input n_649;
input n_552;
input n_547;
input n_43;
input n_721;
input n_116;
input n_22;
input n_467;
input n_564;
input n_423;
input n_284;
input n_46;
input n_245;
input n_21;
input n_501;
input n_725;
input n_139;
input n_38;
input n_105;
input n_280;
input n_590;
input n_629;
input n_672;
input n_4;
input n_378;
input n_551;
input n_17;
input n_581;
input n_688;
input n_382;
input n_554;
input n_254;
input n_690;
input n_33;
input n_23;
input n_583;
input n_671;
input n_718;
input n_302;
input n_265;
input n_526;
input n_719;
input n_293;
input n_372;
input n_443;
input n_244;
input n_677;
input n_47;
input n_173;
input n_198;
input n_714;
input n_447;
input n_247;
input n_314;
input n_368;
input n_433;
input n_604;
input n_8;
input n_321;
input n_292;
input n_625;
input n_621;
input n_100;
input n_455;
input n_674;
input n_417;
input n_612;
input n_212;
input n_385;
input n_498;
input n_516;
input n_507;
input n_119;
input n_497;
input n_689;
input n_738;
input n_606;
input n_559;
input n_275;
input n_640;
input n_252;
input n_624;
input n_26;
input n_295;
input n_133;
input n_330;
input n_508;
input n_739;
input n_506;
input n_2;
input n_737;
input n_610;
input n_692;
input n_6;
input n_509;
input n_568;
input n_39;
input n_147;
input n_373;
input n_67;
input n_307;
input n_633;
input n_439;
input n_87;
input n_150;
input n_530;
input n_556;
input n_106;
input n_209;
input n_259;
input n_448;
input n_668;
input n_733;
input n_375;
input n_301;
input n_576;
input n_68;
input n_93;
input n_186;
input n_537;
input n_134;
input n_191;
input n_587;
input n_659;
input n_51;
input n_63;
input n_492;
input n_563;
input n_171;
input n_153;
input n_524;
input n_399;
input n_341;
input n_204;
input n_394;
input n_250;
input n_579;
input n_548;
input n_543;
input n_260;
input n_298;
input n_650;
input n_320;
input n_694;
input n_518;
input n_505;
input n_286;
input n_122;
input n_282;
input n_331;
input n_10;
input n_24;
input n_406;
input n_519;
input n_470;
input n_325;
input n_449;
input n_132;
input n_90;
input n_724;
input n_546;
input n_101;
input n_658;
input n_281;
input n_240;
input n_381;
input n_189;
input n_220;
input n_291;
input n_231;
input n_257;
input n_390;
input n_731;
input n_31;
input n_456;
input n_13;
input n_371;
input n_481;
input n_535;
input n_709;
input n_152;
input n_540;
input n_317;
input n_618;
input n_9;
input n_323;
input n_569;
input n_195;
input n_42;
input n_356;
input n_227;
input n_592;
input n_45;
input n_271;
input n_94;
input n_335;
input n_123;
input n_654;
input n_370;
input n_167;
input n_234;
input n_343;
input n_308;
input n_379;
input n_428;
input n_267;
input n_514;
input n_457;
input n_570;
input n_297;
input n_156;
input n_5;
input n_603;
input n_225;
input n_377;
input n_484;
input n_219;
input n_442;
input n_157;
input n_131;
input n_192;
input n_636;
input n_600;
input n_660;
input n_223;
input n_392;
input n_158;
input n_655;
input n_704;
input n_138;
input n_264;
input n_109;
input n_669;
input n_472;
input n_454;
input n_387;
input n_374;
input n_163;
input n_276;
input n_339;
input n_95;
input n_183;
input n_185;
input n_243;
input n_398;
input n_396;
input n_635;
input n_347;
input n_169;
input n_59;
input n_522;
input n_550;
input n_255;
input n_696;
input n_215;
input n_350;
input n_196;
input n_662;
input n_459;
input n_646;
input n_211;
input n_218;
input n_400;
input n_181;
input n_436;
input n_3;
input n_290;
input n_580;
input n_221;
input n_178;
input n_622;
input n_723;
input n_386;
input n_578;
input n_287;
input n_344;
input n_555;
input n_473;
input n_422;
input n_475;
input n_72;
input n_661;
input n_104;
input n_41;
input n_682;
input n_415;
input n_56;
input n_141;
input n_485;
input n_496;
input n_355;
input n_486;
input n_670;
input n_15;
input n_336;
input n_584;
input n_681;
input n_591;
input n_145;
input n_48;
input n_521;
input n_614;
input n_663;
input n_50;
input n_337;
input n_430;
input n_313;
input n_631;
input n_673;
input n_88;
input n_479;
input n_528;
input n_510;
input n_216;
input n_680;
input n_168;
input n_395;
input n_164;
input n_432;
input n_553;
input n_727;
input n_311;
input n_208;
input n_142;
input n_214;
input n_328;
input n_140;
input n_299;
input n_303;
input n_369;
input n_675;
input n_296;
input n_613;
input n_241;
input n_637;
input n_357;
input n_598;
input n_685;
input n_608;
input n_184;
input n_446;
input n_445;
input n_65;
input n_78;
input n_144;
input n_114;
input n_96;
input n_691;
input n_717;
input n_165;
input n_468;
input n_499;
input n_213;
input n_129;
input n_342;
input n_482;
input n_517;
input n_98;
input n_588;
input n_361;
input n_464;
input n_363;
input n_402;
input n_413;
input n_734;
input n_638;
input n_700;
input n_197;
input n_107;
input n_573;
input n_69;
input n_236;
input n_388;
input n_1;
input n_249;
input n_740;
input n_304;
input n_329;
input n_203;
input n_274;
input n_577;
input n_384;
input n_582;
input n_460;
input n_80;
input n_35;
input n_73;
input n_277;
input n_92;
input n_19;
input n_338;
input n_149;
input n_477;
input n_461;
input n_333;
input n_571;
input n_693;
input n_309;
input n_30;
input n_512;
input n_14;
input n_84;
input n_462;
input n_130;
input n_322;
input n_567;
input n_258;
input n_652;
input n_29;
input n_79;
input n_151;
input n_25;
input n_306;
input n_722;
input n_458;
input n_288;
input n_188;
input n_190;
input n_201;
input n_263;
input n_471;
input n_609;
input n_44;
input n_224;
input n_40;
input n_34;
input n_228;
input n_283;
input n_383;
input n_711;
input n_474;
input n_112;
input n_542;
input n_85;
input n_463;
input n_488;
input n_595;
input n_736;
input n_502;
input n_239;
input n_466;
input n_420;
input n_630;
input n_489;
input n_632;
input n_699;
input n_55;
input n_617;
input n_49;
input n_310;
input n_54;
input n_593;
input n_504;
input n_511;
input n_12;
input n_586;
input n_465;
input n_76;
input n_358;
input n_362;
input n_170;
input n_332;
input n_27;
input n_77;
input n_102;
input n_161;
input n_273;
input n_349;
input n_585;
input n_270;
input n_616;
input n_230;
input n_81;
input n_118;
input n_601;
input n_279;
input n_70;
input n_253;
input n_261;
input n_174;
input n_289;
input n_627;
input n_172;
input n_206;
input n_217;
input n_440;
input n_726;
input n_478;
input n_545;
input n_441;
input n_450;
input n_648;
input n_312;
input n_476;
input n_429;
input n_534;
input n_345;
input n_210;
input n_494;
input n_641;
input n_628;
input n_365;
input n_91;
input n_729;
input n_730;
input n_176;
input n_557;
input n_182;
input n_143;
input n_83;
input n_354;
input n_575;
input n_607;
input n_480;
input n_647;
input n_237;
input n_425;
input n_513;
input n_407;
input n_527;
input n_679;
input n_707;
input n_710;
input n_695;
input n_180;
input n_560;
input n_656;
input n_340;
input n_207;
input n_561;
input n_37;
input n_346;
input n_393;
input n_229;
input n_108;
input n_487;
input n_495;
input n_602;
input n_665;
input n_574;
input n_437;
input n_66;
input n_177;
input n_60;
input n_403;
input n_453;
input n_421;
input n_16;
input n_720;
input n_0;
input n_58;
input n_623;
input n_405;
input n_18;
input n_359;
input n_490;
input n_117;
input n_326;
input n_233;
input n_404;
input n_686;
input n_205;
input n_366;
input n_572;
input n_113;
input n_712;
input n_246;
input n_596;
input n_179;
input n_125;
input n_410;
input n_558;
input n_708;
input n_269;
input n_529;
input n_128;
input n_735;
input n_702;
input n_285;
input n_412;
input n_120;
input n_232;
input n_327;
input n_135;
input n_657;
input n_126;
input n_644;
input n_728;
input n_202;
input n_266;
input n_272;
input n_491;
input n_427;
input n_732;
input n_193;
input n_251;
input n_352;
input n_53;
input n_160;
input n_565;
input n_426;
input n_520;
input n_566;
input n_409;
input n_589;
input n_716;
input n_597;
input n_500;
input n_562;
input n_154;
input n_62;
input n_148;
input n_71;
input n_300;
input n_651;
input n_435;
input n_159;
input n_334;
input n_599;
input n_541;
input n_391;
input n_701;
input n_434;
input n_645;
input n_539;
input n_175;
input n_538;
input n_666;
input n_262;
input n_238;
input n_639;
input n_99;
input n_687;
input n_715;
input n_411;
input n_414;
input n_319;
input n_364;
input n_20;
input n_536;
input n_531;
input n_121;
input n_242;
input n_360;
input n_36;
input n_594;
input n_200;
input n_162;
input n_64;
input n_222;
input n_28;
input n_89;
input n_438;
input n_115;
input n_713;
input n_324;
input n_634;
input n_416;
input n_199;
input n_187;
input n_32;
input n_401;
input n_103;
input n_348;
input n_97;
input n_166;
input n_626;
input n_11;
input n_424;
input n_7;
input n_706;
input n_256;
input n_305;
input n_533;
input n_52;
input n_278;
input n_110;

output n_2496;

wire n_924;
wire n_1263;
wire n_977;
wire n_1378;
wire n_2417;
wire n_2253;
wire n_1126;
wire n_1423;
wire n_1729;
wire n_1166;
wire n_2380;
wire n_1751;
wire n_1508;
wire n_785;
wire n_2200;
wire n_1161;
wire n_1859;
wire n_1677;
wire n_1150;
wire n_2327;
wire n_1780;
wire n_1488;
wire n_790;
wire n_1055;
wire n_2386;
wire n_1501;
wire n_2395;
wire n_880;
wire n_1007;
wire n_2369;
wire n_1528;
wire n_1370;
wire n_1292;
wire n_2347;
wire n_1198;
wire n_1360;
wire n_2388;
wire n_1099;
wire n_956;
wire n_1738;
wire n_2021;
wire n_2134;
wire n_2391;
wire n_1021;
wire n_1960;
wire n_2185;
wire n_2143;
wire n_2059;
wire n_1323;
wire n_1466;
wire n_1695;
wire n_2487;
wire n_1353;
wire n_800;
wire n_1347;
wire n_2495;
wire n_1535;
wire n_1789;
wire n_1666;
wire n_2389;
wire n_819;
wire n_1451;
wire n_1022;
wire n_2302;
wire n_915;
wire n_1545;
wire n_2374;
wire n_864;
wire n_859;
wire n_951;
wire n_1947;
wire n_1264;
wire n_2114;
wire n_2001;
wire n_1494;
wire n_854;
wire n_1462;
wire n_1799;
wire n_2069;
wire n_2396;
wire n_1580;
wire n_1939;
wire n_2486;
wire n_1806;
wire n_933;
wire n_2244;
wire n_2257;
wire n_1152;
wire n_1869;
wire n_1607;
wire n_1563;
wire n_2011;
wire n_2096;
wire n_877;
wire n_2105;
wire n_2024;
wire n_1696;
wire n_2483;
wire n_755;
wire n_1118;
wire n_1686;
wire n_947;
wire n_1285;
wire n_1860;
wire n_1359;
wire n_1728;
wire n_1107;
wire n_2076;
wire n_2031;
wire n_2482;
wire n_1230;
wire n_1896;
wire n_2165;
wire n_2147;
wire n_929;
wire n_1124;
wire n_1818;
wire n_2127;
wire n_902;
wire n_1576;
wire n_1104;
wire n_1294;
wire n_1705;
wire n_1257;
wire n_1182;
wire n_1698;
wire n_1261;
wire n_2329;
wire n_938;
wire n_1098;
wire n_2142;
wire n_1154;
wire n_2189;
wire n_1242;
wire n_1135;
wire n_2323;
wire n_2203;
wire n_1016;
wire n_1243;
wire n_2047;
wire n_1280;
wire n_1845;
wire n_2052;
wire n_2193;
wire n_2058;
wire n_2458;
wire n_2478;
wire n_1483;
wire n_1314;
wire n_1512;
wire n_1490;
wire n_1236;
wire n_1633;
wire n_2144;
wire n_1778;
wire n_2306;
wire n_920;
wire n_1289;
wire n_1517;
wire n_2091;
wire n_2466;
wire n_2085;
wire n_1669;
wire n_976;
wire n_1949;
wire n_1449;
wire n_1946;
wire n_1566;
wire n_2032;
wire n_2149;
wire n_1078;
wire n_1670;
wire n_775;
wire n_1484;
wire n_2071;
wire n_1374;
wire n_1328;
wire n_2141;
wire n_1948;
wire n_1984;
wire n_2099;
wire n_2408;
wire n_1877;
wire n_1831;
wire n_1598;
wire n_1723;
wire n_955;
wire n_1850;
wire n_1146;
wire n_882;
wire n_2384;
wire n_1036;
wire n_1097;
wire n_1749;
wire n_897;
wire n_798;
wire n_1428;
wire n_1394;
wire n_1414;
wire n_1216;
wire n_1040;
wire n_2202;
wire n_1872;
wire n_1852;
wire n_2159;
wire n_926;
wire n_2180;
wire n_2249;
wire n_2353;
wire n_1218;
wire n_1931;
wire n_2439;
wire n_2276;
wire n_1070;
wire n_777;
wire n_1547;
wire n_2089;
wire n_1030;
wire n_2470;
wire n_1755;
wire n_1071;
wire n_1165;
wire n_1267;
wire n_1561;
wire n_1801;
wire n_1391;
wire n_958;
wire n_1034;
wire n_1513;
wire n_1600;
wire n_845;
wire n_2235;
wire n_1862;
wire n_837;
wire n_1239;
wire n_2300;
wire n_1796;
wire n_1473;
wire n_1587;
wire n_901;
wire n_2432;
wire n_813;
wire n_1521;
wire n_1284;
wire n_1590;
wire n_2174;
wire n_1748;
wire n_1672;
wire n_888;
wire n_1880;
wire n_2337;
wire n_1167;
wire n_1626;
wire n_1384;
wire n_1556;
wire n_1863;
wire n_1064;
wire n_858;
wire n_2079;
wire n_2238;
wire n_923;
wire n_2118;
wire n_1151;
wire n_881;
wire n_1405;
wire n_2407;
wire n_1706;
wire n_1582;
wire n_1069;
wire n_1784;
wire n_1075;
wire n_1836;
wire n_1450;
wire n_1322;
wire n_2101;
wire n_1471;
wire n_1986;
wire n_2072;
wire n_1750;
wire n_1459;
wire n_889;
wire n_2358;
wire n_973;
wire n_1700;
wire n_1585;
wire n_1971;
wire n_1599;
wire n_2275;
wire n_1211;
wire n_1197;
wire n_1523;
wire n_1950;
wire n_907;
wire n_1447;
wire n_2251;
wire n_1377;
wire n_2370;
wire n_989;
wire n_1039;
wire n_2214;
wire n_2055;
wire n_1403;
wire n_2248;
wire n_2356;
wire n_892;
wire n_1000;
wire n_1202;
wire n_1278;
wire n_2062;
wire n_1002;
wire n_1463;
wire n_1581;
wire n_2100;
wire n_2258;
wire n_748;
wire n_1058;
wire n_1667;
wire n_838;
wire n_1053;
wire n_1224;
wire n_1926;
wire n_1248;
wire n_1331;
wire n_953;
wire n_1014;
wire n_1241;
wire n_2150;
wire n_2241;
wire n_2152;
wire n_963;
wire n_1052;
wire n_954;
wire n_1385;
wire n_793;
wire n_2140;
wire n_2385;
wire n_1819;
wire n_2330;
wire n_2139;
wire n_1527;
wire n_2042;
wire n_1882;
wire n_884;
wire n_944;
wire n_1754;
wire n_1623;
wire n_2175;
wire n_2324;
wire n_1854;
wire n_1565;
wire n_1809;
wire n_1856;
wire n_1072;
wire n_2218;
wire n_2267;
wire n_857;
wire n_832;
wire n_2305;
wire n_2450;
wire n_1319;
wire n_2379;
wire n_2154;
wire n_1825;
wire n_1951;
wire n_1883;
wire n_1906;
wire n_1712;
wire n_1387;
wire n_2262;
wire n_2462;
wire n_1532;
wire n_2322;
wire n_2271;
wire n_1027;
wire n_971;
wire n_1156;
wire n_794;
wire n_2331;
wire n_2293;
wire n_847;
wire n_1393;
wire n_2319;
wire n_1775;
wire n_2028;
wire n_1368;
wire n_1276;
wire n_822;
wire n_1412;
wire n_1709;
wire n_2108;
wire n_1162;
wire n_1538;
wire n_1838;
wire n_1199;
wire n_1847;
wire n_1779;
wire n_1884;
wire n_2434;
wire n_1038;
wire n_1369;
wire n_1841;
wire n_1660;
wire n_887;
wire n_1905;
wire n_2195;
wire n_809;
wire n_870;
wire n_931;
wire n_1711;
wire n_1662;
wire n_1891;
wire n_1481;
wire n_1942;
wire n_1978;
wire n_1544;
wire n_868;
wire n_2454;
wire n_914;
wire n_2120;
wire n_1629;
wire n_1293;
wire n_965;
wire n_1876;
wire n_1743;
wire n_935;
wire n_817;
wire n_1175;
wire n_1479;
wire n_1810;
wire n_2350;
wire n_1888;
wire n_2009;
wire n_759;
wire n_2222;
wire n_1892;
wire n_806;
wire n_1997;
wire n_1766;
wire n_1477;
wire n_1635;
wire n_1963;
wire n_2226;
wire n_1571;
wire n_1189;
wire n_2215;
wire n_1259;
wire n_1690;
wire n_746;
wire n_1649;
wire n_747;
wire n_2064;
wire n_784;
wire n_2449;
wire n_1733;
wire n_1244;
wire n_2413;
wire n_1194;
wire n_1925;
wire n_2297;
wire n_1815;
wire n_851;
wire n_1759;
wire n_843;
wire n_1788;
wire n_2177;
wire n_2491;
wire n_913;
wire n_1537;
wire n_865;
wire n_2227;
wire n_1222;
wire n_1679;
wire n_2190;
wire n_776;
wire n_1798;
wire n_2022;
wire n_1790;
wire n_1415;
wire n_1260;
wire n_1746;
wire n_1647;
wire n_2181;
wire n_2479;
wire n_1829;
wire n_1464;
wire n_1444;
wire n_1191;
wire n_2387;
wire n_1674;
wire n_1833;
wire n_1830;
wire n_2073;
wire n_1710;
wire n_1128;
wire n_1734;
wire n_744;
wire n_1308;
wire n_2178;
wire n_1767;
wire n_2336;
wire n_1680;
wire n_1233;
wire n_1615;
wire n_1529;
wire n_2005;
wire n_1916;
wire n_1333;
wire n_2469;
wire n_1121;
wire n_2007;
wire n_949;
wire n_1443;
wire n_1008;
wire n_946;
wire n_1539;
wire n_1001;
wire n_1503;
wire n_2054;
wire n_1468;
wire n_1559;
wire n_1765;
wire n_1866;
wire n_1624;
wire n_1510;
wire n_1380;
wire n_1744;
wire n_1617;
wire n_1010;
wire n_1994;
wire n_1231;
wire n_1279;
wire n_1406;
wire n_1195;
wire n_1839;
wire n_1837;
wire n_1760;
wire n_936;
wire n_1500;
wire n_1090;
wire n_757;
wire n_2342;
wire n_1832;
wire n_1851;
wire n_758;
wire n_999;
wire n_2046;
wire n_1933;
wire n_2290;
wire n_1656;
wire n_1158;
wire n_2045;
wire n_1509;
wire n_1874;
wire n_2040;
wire n_2060;
wire n_1987;
wire n_1145;
wire n_878;
wire n_1678;
wire n_1049;
wire n_1153;
wire n_2145;
wire n_741;
wire n_1639;
wire n_1306;
wire n_1068;
wire n_1871;
wire n_1964;
wire n_1163;
wire n_906;
wire n_2039;
wire n_1207;
wire n_919;
wire n_908;
wire n_2412;
wire n_2406;
wire n_1781;
wire n_2084;
wire n_2035;
wire n_2061;
wire n_2378;
wire n_1740;
wire n_2398;
wire n_1362;
wire n_1586;
wire n_959;
wire n_2459;
wire n_940;
wire n_1445;
wire n_1492;
wire n_2155;
wire n_1923;
wire n_1773;
wire n_1169;
wire n_1596;
wire n_1692;
wire n_1017;
wire n_2481;
wire n_2171;
wire n_978;
wire n_2116;
wire n_2314;
wire n_1434;
wire n_1054;
wire n_1474;
wire n_1665;
wire n_1269;
wire n_2420;
wire n_1095;
wire n_1828;
wire n_1614;
wire n_1079;
wire n_1045;
wire n_1208;
wire n_2093;
wire n_2038;
wire n_2320;
wire n_2339;
wire n_2473;
wire n_2137;
wire n_1431;
wire n_1593;
wire n_1033;
wire n_2299;
wire n_2087;
wire n_1640;
wire n_2162;
wire n_1732;
wire n_1009;
wire n_1148;
wire n_2051;
wire n_750;
wire n_742;
wire n_2029;
wire n_995;
wire n_2168;
wire n_1609;
wire n_1989;
wire n_2359;
wire n_1887;
wire n_1383;
wire n_1073;
wire n_2457;
wire n_2346;
wire n_2312;
wire n_962;
wire n_1215;
wire n_1171;
wire n_1578;
wire n_1920;
wire n_1065;
wire n_1592;
wire n_1336;
wire n_1721;
wire n_1959;
wire n_1758;
wire n_2338;
wire n_1574;
wire n_2399;
wire n_2048;
wire n_2355;
wire n_2133;
wire n_1921;
wire n_1309;
wire n_1878;
wire n_1426;
wire n_1043;
wire n_1800;
wire n_1548;
wire n_1421;
wire n_1286;
wire n_1177;
wire n_1355;
wire n_974;
wire n_1159;
wire n_957;
wire n_773;
wire n_2124;
wire n_743;
wire n_2081;
wire n_1119;
wire n_2156;
wire n_1240;
wire n_2261;
wire n_1820;
wire n_2418;
wire n_829;
wire n_1612;
wire n_2179;
wire n_1416;
wire n_2077;
wire n_1724;
wire n_2111;
wire n_1237;
wire n_1420;
wire n_1132;
wire n_1366;
wire n_1300;
wire n_1127;
wire n_2277;
wire n_761;
wire n_2477;
wire n_1785;
wire n_1568;
wire n_1006;
wire n_2110;
wire n_1270;
wire n_1664;
wire n_1486;
wire n_1332;
wire n_2231;
wire n_1390;
wire n_2017;
wire n_2474;
wire n_2090;
wire n_1870;
wire n_2367;
wire n_1591;
wire n_2033;
wire n_1682;
wire n_1980;
wire n_2390;
wire n_1249;
wire n_1111;
wire n_1365;
wire n_1927;
wire n_2132;
wire n_1349;
wire n_1093;
wire n_2400;
wire n_1031;
wire n_1041;
wire n_1265;
wire n_1909;
wire n_1562;
wire n_834;
wire n_765;
wire n_2255;
wire n_2424;
wire n_2272;
wire n_893;
wire n_1015;
wire n_1140;
wire n_891;
wire n_1651;
wire n_1965;
wire n_1902;
wire n_2151;
wire n_1941;
wire n_2106;
wire n_1913;
wire n_1823;
wire n_874;
wire n_2464;
wire n_1101;
wire n_1106;
wire n_1456;
wire n_2230;
wire n_2015;
wire n_2365;
wire n_1875;
wire n_1982;
wire n_1304;
wire n_1324;
wire n_987;
wire n_1846;
wire n_2066;
wire n_1885;
wire n_1455;
wire n_767;
wire n_993;
wire n_1903;
wire n_2490;
wire n_1407;
wire n_2452;
wire n_1551;
wire n_860;
wire n_1805;
wire n_2176;
wire n_2204;
wire n_1816;
wire n_948;
wire n_1217;
wire n_2220;
wire n_2455;
wire n_1849;
wire n_2410;
wire n_1131;
wire n_1084;
wire n_1961;
wire n_970;
wire n_1935;
wire n_911;
wire n_1430;
wire n_2467;
wire n_1094;
wire n_1354;
wire n_1534;
wire n_2288;
wire n_1351;
wire n_2240;
wire n_1044;
wire n_1205;
wire n_2436;
wire n_1209;
wire n_1552;
wire n_1435;
wire n_879;
wire n_2416;
wire n_2405;
wire n_2088;
wire n_824;
wire n_1645;
wire n_2461;
wire n_1327;
wire n_2243;
wire n_996;
wire n_921;
wire n_1684;
wire n_1717;
wire n_815;
wire n_1795;
wire n_2128;
wire n_1821;
wire n_1381;
wire n_1611;
wire n_1037;
wire n_2368;
wire n_1080;
wire n_2301;
wire n_1274;
wire n_1316;
wire n_1708;
wire n_2419;
wire n_1438;
wire n_1082;
wire n_1840;
wire n_1630;
wire n_2122;
wire n_1436;
wire n_1691;
wire n_952;
wire n_2092;
wire n_1229;
wire n_1437;
wire n_1023;
wire n_2075;
wire n_803;
wire n_1092;
wire n_1776;
wire n_2198;
wire n_2281;
wire n_2131;
wire n_2216;
wire n_1757;
wire n_890;
wire n_1897;
wire n_764;
wire n_1919;
wire n_1056;
wire n_1424;
wire n_960;
wire n_2308;
wire n_1893;
wire n_1290;
wire n_1123;
wire n_1467;
wire n_1047;
wire n_2053;
wire n_2163;
wire n_2328;
wire n_1958;
wire n_2254;
wire n_1252;
wire n_1382;
wire n_1029;
wire n_925;
wire n_1206;
wire n_1311;
wire n_2191;
wire n_1519;
wire n_950;
wire n_2428;
wire n_1553;
wire n_1811;
wire n_2443;
wire n_1346;
wire n_1299;
wire n_2158;
wire n_1808;
wire n_1060;
wire n_1141;
wire n_2266;
wire n_2465;
wire n_912;
wire n_968;
wire n_2440;
wire n_1386;
wire n_1699;
wire n_967;
wire n_1442;
wire n_1139;
wire n_2333;
wire n_885;
wire n_1432;
wire n_1357;
wire n_2125;
wire n_1632;
wire n_1057;
wire n_1051;
wire n_1085;
wire n_1066;
wire n_2402;
wire n_1157;
wire n_2403;
wire n_1050;
wire n_841;
wire n_802;
wire n_1954;
wire n_2265;
wire n_1608;
wire n_983;
wire n_1844;
wire n_1305;
wire n_873;
wire n_1826;
wire n_1112;
wire n_2304;
wire n_762;
wire n_1283;
wire n_1644;
wire n_2334;
wire n_1974;
wire n_2463;
wire n_2086;
wire n_2289;
wire n_1343;
wire n_2263;
wire n_1203;
wire n_1631;
wire n_2472;
wire n_821;
wire n_1763;
wire n_2341;
wire n_1966;
wire n_1768;
wire n_2294;
wire n_1179;
wire n_753;
wire n_2475;
wire n_1048;
wire n_1719;
wire n_1288;
wire n_2269;
wire n_2309;
wire n_2415;
wire n_1560;
wire n_1605;
wire n_2236;
wire n_1228;
wire n_2123;
wire n_972;
wire n_2037;
wire n_1953;
wire n_1938;
wire n_820;
wire n_1200;
wire n_1911;
wire n_2460;
wire n_1363;
wire n_1301;
wire n_1668;
wire n_1185;
wire n_991;
wire n_828;
wire n_1967;
wire n_779;
wire n_1143;
wire n_1579;
wire n_2233;
wire n_1329;
wire n_1312;
wire n_1439;
wire n_804;
wire n_1688;
wire n_945;
wire n_1504;
wire n_943;
wire n_992;
wire n_1932;
wire n_842;
wire n_984;
wire n_2082;
wire n_1992;
wire n_2429;
wire n_1643;
wire n_883;
wire n_1983;
wire n_1594;
wire n_1214;
wire n_1342;
wire n_1400;
wire n_900;
wire n_2362;
wire n_856;
wire n_1793;
wire n_1976;
wire n_2223;
wire n_918;
wire n_942;
wire n_2169;
wire n_1804;
wire n_1147;
wire n_1557;
wire n_1977;
wire n_2153;
wire n_2468;
wire n_1610;
wire n_1077;
wire n_1422;
wire n_2364;
wire n_896;
wire n_2310;
wire n_2287;
wire n_2291;
wire n_894;
wire n_1636;
wire n_2056;
wire n_1730;
wire n_831;
wire n_2280;
wire n_2192;
wire n_964;
wire n_1373;
wire n_1350;
wire n_1511;
wire n_1865;
wire n_1470;
wire n_1096;
wire n_2094;
wire n_1575;
wire n_1735;
wire n_1697;
wire n_833;
wire n_2318;
wire n_2393;
wire n_2020;
wire n_1646;
wire n_1307;
wire n_1881;
wire n_988;
wire n_2043;
wire n_1940;
wire n_814;
wire n_1549;
wire n_1934;
wire n_2311;
wire n_1201;
wire n_1114;
wire n_2025;
wire n_1616;
wire n_1446;
wire n_2285;
wire n_1458;
wire n_1176;
wire n_1472;
wire n_2298;
wire n_2471;
wire n_1807;
wire n_1149;
wire n_1671;
wire n_763;
wire n_1020;
wire n_1062;
wire n_2303;
wire n_1824;
wire n_1917;
wire n_2295;
wire n_1219;
wire n_1204;
wire n_2325;
wire n_2446;
wire n_1814;
wire n_1035;
wire n_783;
wire n_1848;
wire n_1928;
wire n_2126;
wire n_1188;
wire n_1722;
wire n_2441;
wire n_1802;
wire n_849;
wire n_1638;
wire n_1786;
wire n_2002;
wire n_2282;
wire n_2371;
wire n_830;
wire n_2098;
wire n_1296;
wire n_2352;
wire n_1413;
wire n_801;
wire n_2207;
wire n_2080;
wire n_2377;
wire n_2340;
wire n_2444;
wire n_2068;
wire n_875;
wire n_1110;
wire n_1655;
wire n_749;
wire n_1895;
wire n_1134;
wire n_1358;
wire n_939;
wire n_2361;
wire n_1088;
wire n_1173;
wire n_789;
wire n_1232;
wire n_1603;
wire n_866;
wire n_969;
wire n_1401;
wire n_2492;
wire n_1019;
wire n_1105;
wire n_1998;
wire n_1338;
wire n_2016;
wire n_1522;
wire n_1687;
wire n_1637;
wire n_2034;
wire n_1419;
wire n_1653;
wire n_2270;
wire n_1506;
wire n_836;
wire n_990;
wire n_1886;
wire n_1389;
wire n_1894;
wire n_975;
wire n_1908;
wire n_1256;
wire n_1702;
wire n_2259;
wire n_1465;
wire n_778;
wire n_1122;
wire n_770;
wire n_1375;
wire n_2494;
wire n_1102;
wire n_2392;
wire n_1843;
wire n_1499;
wire n_1187;
wire n_1441;
wire n_2435;
wire n_1392;
wire n_1597;
wire n_1929;
wire n_1164;
wire n_1659;
wire n_1834;
wire n_2097;
wire n_2313;
wire n_1174;
wire n_2431;
wire n_1371;
wire n_1303;
wire n_2206;
wire n_2063;
wire n_1572;
wire n_1968;
wire n_2252;
wire n_876;
wire n_1516;
wire n_1190;
wire n_1736;
wire n_1685;
wire n_2409;
wire n_917;
wire n_1714;
wire n_966;
wire n_1116;
wire n_2000;
wire n_1661;
wire n_1212;
wire n_2074;
wire n_1541;
wire n_982;
wire n_1573;
wire n_1453;
wire n_1731;
wire n_2217;
wire n_818;
wire n_2373;
wire n_1970;
wire n_861;
wire n_1713;
wire n_1183;
wire n_2307;
wire n_1658;
wire n_899;
wire n_1253;
wire n_1737;
wire n_2201;
wire n_2117;
wire n_1904;
wire n_1993;
wire n_774;
wire n_1628;
wire n_2493;
wire n_2205;
wire n_1335;
wire n_1514;
wire n_1777;
wire n_1957;
wire n_1059;
wire n_1345;
wire n_1133;
wire n_1771;
wire n_1912;
wire n_1899;
wire n_1410;
wire n_1005;
wire n_1003;
wire n_2067;
wire n_1168;
wire n_2219;
wire n_2437;
wire n_2148;
wire n_937;
wire n_2445;
wire n_1427;
wire n_1584;
wire n_1726;
wire n_1835;
wire n_1440;
wire n_2164;
wire n_1988;
wire n_2115;
wire n_1853;
wire n_1356;
wire n_1787;
wire n_910;
wire n_2232;
wire n_2212;
wire n_1657;
wire n_768;
wire n_1475;
wire n_1302;
wire n_1774;
wire n_1725;
wire n_1313;
wire n_1136;
wire n_1491;
wire n_754;
wire n_1496;
wire n_1125;
wire n_1812;
wire n_1915;
wire n_1109;
wire n_895;
wire n_1310;
wire n_2121;
wire n_1803;
wire n_1399;
wire n_1543;
wire n_1991;
wire n_1979;
wire n_791;
wire n_1533;
wire n_2224;
wire n_808;
wire n_2484;
wire n_797;
wire n_1025;
wire n_1930;
wire n_1955;
wire n_1067;
wire n_1720;
wire n_2401;
wire n_2003;
wire n_766;
wire n_1457;
wire n_2354;
wire n_2246;
wire n_2008;
wire n_1117;
wire n_799;
wire n_2264;
wire n_1742;
wire n_1480;
wire n_1482;
wire n_1213;
wire n_2489;
wire n_1266;
wire n_872;
wire n_2012;
wire n_1291;
wire n_1297;
wire n_1753;
wire n_2283;
wire n_1782;
wire n_2245;
wire n_1155;
wire n_1418;
wire n_1972;
wire n_1689;
wire n_1524;
wire n_1485;
wire n_1011;
wire n_1184;
wire n_2184;
wire n_985;
wire n_1855;
wire n_2425;
wire n_869;
wire n_810;
wire n_827;
wire n_1703;
wire n_1352;
wire n_2197;
wire n_2199;
wire n_1650;
wire n_1144;
wire n_1137;
wire n_1570;
wire n_1170;
wire n_2023;
wire n_2213;
wire n_2351;
wire n_2211;
wire n_2095;
wire n_2103;
wire n_2160;
wire n_2228;
wire n_1602;
wire n_855;
wire n_1178;
wire n_1461;
wire n_850;
wire n_2421;
wire n_2286;
wire n_1999;
wire n_2372;
wire n_2065;
wire n_2136;
wire n_2480;
wire n_1372;
wire n_1273;
wire n_1822;
wire n_2363;
wire n_2430;
wire n_916;
wire n_1081;
wire n_2332;
wire n_1235;
wire n_1115;
wire n_980;
wire n_2433;
wire n_1282;
wire n_1318;
wire n_1783;
wire n_780;
wire n_998;
wire n_2375;
wire n_1454;
wire n_1227;
wire n_1531;
wire n_840;
wire n_1334;
wire n_1907;
wire n_823;
wire n_2344;
wire n_1388;
wire n_1417;
wire n_1295;
wire n_2316;
wire n_1985;
wire n_1898;
wire n_2107;
wire n_1625;
wire n_2130;
wire n_2187;
wire n_2284;
wire n_898;
wire n_1762;
wire n_1013;
wire n_1452;
wire n_1120;
wire n_1791;
wire n_1890;
wire n_1747;
wire n_1683;
wire n_1817;
wire n_909;
wire n_1944;
wire n_1497;
wire n_1530;
wire n_997;
wire n_932;
wire n_2078;
wire n_1409;
wire n_788;
wire n_1326;
wire n_1268;
wire n_825;
wire n_1981;
wire n_2186;
wire n_1320;
wire n_1663;
wire n_1718;
wire n_986;
wire n_2315;
wire n_1317;
wire n_1518;
wire n_1715;
wire n_2102;
wire n_1281;
wire n_1952;
wire n_1192;
wire n_2221;
wire n_1024;
wire n_1063;
wire n_1889;
wire n_1792;
wire n_1564;
wire n_1868;
wire n_1613;
wire n_1489;
wire n_1922;
wire n_1376;
wire n_941;
wire n_2326;
wire n_981;
wire n_1569;
wire n_2188;
wire n_867;
wire n_2348;
wire n_2422;
wire n_2239;
wire n_792;
wire n_756;
wire n_1429;
wire n_1238;
wire n_2448;
wire n_812;
wire n_2104;
wire n_2057;
wire n_1772;
wire n_752;
wire n_905;
wire n_1476;
wire n_1108;
wire n_782;
wire n_1100;
wire n_1861;
wire n_2129;
wire n_1395;
wire n_862;
wire n_1425;
wire n_760;
wire n_1901;
wire n_1900;
wire n_1620;
wire n_1330;
wire n_1867;
wire n_1945;
wire n_1675;
wire n_1924;
wire n_1727;
wire n_1554;
wire n_1745;
wire n_769;
wire n_2006;
wire n_1995;
wire n_2411;
wire n_2138;
wire n_1046;
wire n_934;
wire n_1618;
wire n_2260;
wire n_826;
wire n_2343;
wire n_1813;
wire n_2447;
wire n_886;
wire n_2014;
wire n_1221;
wire n_2345;
wire n_1172;
wire n_1341;
wire n_1641;
wire n_1361;
wire n_2382;
wire n_1707;
wire n_853;
wire n_2317;
wire n_751;
wire n_2172;
wire n_1973;
wire n_1083;
wire n_786;
wire n_1142;
wire n_2376;
wire n_2488;
wire n_1129;
wire n_2476;
wire n_787;
wire n_1770;
wire n_2456;
wire n_961;
wire n_2250;
wire n_1756;
wire n_771;
wire n_1716;
wire n_1225;
wire n_1520;
wire n_2451;
wire n_1287;
wire n_1262;
wire n_930;
wire n_1873;
wire n_1411;
wire n_1962;
wire n_1577;
wire n_2423;
wire n_1087;
wire n_994;
wire n_1701;
wire n_2194;
wire n_848;
wire n_1550;
wire n_1498;
wire n_2167;
wire n_1223;
wire n_1272;
wire n_1567;
wire n_1247;
wire n_922;
wire n_816;
wire n_1648;
wire n_1536;
wire n_1857;
wire n_1344;
wire n_2041;
wire n_1246;
wire n_1339;
wire n_1478;
wire n_1797;
wire n_1769;
wire n_839;
wire n_1210;
wire n_1364;
wire n_2357;
wire n_2183;
wire n_2360;
wire n_2292;
wire n_1250;
wire n_2173;
wire n_1842;
wire n_871;
wire n_2442;
wire n_928;
wire n_1367;
wire n_1943;
wire n_1460;
wire n_772;
wire n_2018;
wire n_1555;
wire n_1589;
wire n_1086;
wire n_796;
wire n_1858;
wire n_1619;
wire n_2119;
wire n_1502;
wire n_2157;
wire n_1469;
wire n_1012;
wire n_1396;
wire n_1348;
wire n_2030;
wire n_903;
wire n_2453;
wire n_1525;
wire n_1752;
wire n_2397;
wire n_2208;
wire n_1404;
wire n_1794;
wire n_2182;
wire n_1315;
wire n_2234;
wire n_1061;
wire n_1910;
wire n_1298;
wire n_1652;
wire n_2209;
wire n_2050;
wire n_1193;
wire n_1676;
wire n_1255;
wire n_1113;
wire n_2321;
wire n_1226;
wire n_1277;
wire n_2146;
wire n_844;
wire n_852;
wire n_1487;
wire n_1864;
wire n_1028;
wire n_1601;
wire n_781;
wire n_1546;
wire n_1337;
wire n_1495;
wire n_979;
wire n_1515;
wire n_1627;
wire n_1245;
wire n_846;
wire n_2427;
wire n_2438;
wire n_1673;
wire n_1321;
wire n_1975;
wire n_2296;
wire n_2070;
wire n_1937;
wire n_2112;
wire n_1739;
wire n_2278;
wire n_2394;
wire n_1914;
wire n_2135;
wire n_2335;
wire n_745;
wire n_2381;
wire n_1654;
wire n_2349;
wire n_1103;
wire n_1379;
wire n_2196;
wire n_2170;
wire n_1076;
wire n_1091;
wire n_1408;
wire n_1761;
wire n_2036;
wire n_1325;
wire n_1595;
wire n_2161;
wire n_795;
wire n_2404;
wire n_2083;
wire n_1606;
wire n_1220;
wire n_1694;
wire n_1540;
wire n_2485;
wire n_1956;
wire n_1936;
wire n_1642;
wire n_2279;
wire n_2027;
wire n_1130;
wire n_2366;
wire n_1918;
wire n_1526;
wire n_863;
wire n_2210;
wire n_805;
wire n_1604;
wire n_1275;
wire n_1764;
wire n_2414;
wire n_1583;
wire n_2426;
wire n_1042;
wire n_1402;
wire n_2049;
wire n_2273;
wire n_1493;
wire n_1741;
wire n_2229;
wire n_1160;
wire n_1397;
wire n_1258;
wire n_1074;
wire n_2004;
wire n_1621;
wire n_2113;
wire n_1448;
wire n_2225;
wire n_1507;
wire n_1398;
wire n_2383;
wire n_1879;
wire n_1996;
wire n_1181;
wire n_1505;
wire n_1634;
wire n_1196;
wire n_2019;
wire n_1340;
wire n_2274;
wire n_811;
wire n_1558;
wire n_807;
wire n_2166;
wire n_835;
wire n_1433;
wire n_1704;
wire n_2256;
wire n_1254;
wire n_1026;
wire n_2026;
wire n_1969;
wire n_1234;
wire n_2109;
wire n_2044;
wire n_1138;
wire n_1089;
wire n_927;
wire n_2013;
wire n_1990;
wire n_1004;
wire n_1186;
wire n_1032;
wire n_1681;
wire n_2010;
wire n_1018;
wire n_2242;
wire n_2247;
wire n_1693;
wire n_904;
wire n_1588;
wire n_1622;
wire n_2237;
wire n_1180;
wire n_1827;
wire n_1271;
wire n_1542;
wire n_1251;
wire n_2268;

CKINVDCx20_ASAP7_75t_R g741 ( 
.A(n_96),
.Y(n_741)
);

INVx1_ASAP7_75t_L g742 ( 
.A(n_668),
.Y(n_742)
);

CKINVDCx5p33_ASAP7_75t_R g743 ( 
.A(n_698),
.Y(n_743)
);

CKINVDCx5p33_ASAP7_75t_R g744 ( 
.A(n_708),
.Y(n_744)
);

INVx2_ASAP7_75t_L g745 ( 
.A(n_678),
.Y(n_745)
);

CKINVDCx5p33_ASAP7_75t_R g746 ( 
.A(n_182),
.Y(n_746)
);

CKINVDCx16_ASAP7_75t_R g747 ( 
.A(n_178),
.Y(n_747)
);

CKINVDCx20_ASAP7_75t_R g748 ( 
.A(n_650),
.Y(n_748)
);

BUFx3_ASAP7_75t_L g749 ( 
.A(n_455),
.Y(n_749)
);

CKINVDCx20_ASAP7_75t_R g750 ( 
.A(n_732),
.Y(n_750)
);

CKINVDCx5p33_ASAP7_75t_R g751 ( 
.A(n_479),
.Y(n_751)
);

CKINVDCx5p33_ASAP7_75t_R g752 ( 
.A(n_737),
.Y(n_752)
);

CKINVDCx5p33_ASAP7_75t_R g753 ( 
.A(n_143),
.Y(n_753)
);

CKINVDCx5p33_ASAP7_75t_R g754 ( 
.A(n_679),
.Y(n_754)
);

INVx2_ASAP7_75t_L g755 ( 
.A(n_637),
.Y(n_755)
);

CKINVDCx20_ASAP7_75t_R g756 ( 
.A(n_666),
.Y(n_756)
);

CKINVDCx5p33_ASAP7_75t_R g757 ( 
.A(n_558),
.Y(n_757)
);

INVx2_ASAP7_75t_SL g758 ( 
.A(n_428),
.Y(n_758)
);

CKINVDCx16_ASAP7_75t_R g759 ( 
.A(n_630),
.Y(n_759)
);

INVx2_ASAP7_75t_SL g760 ( 
.A(n_348),
.Y(n_760)
);

CKINVDCx5p33_ASAP7_75t_R g761 ( 
.A(n_297),
.Y(n_761)
);

CKINVDCx5p33_ASAP7_75t_R g762 ( 
.A(n_211),
.Y(n_762)
);

CKINVDCx5p33_ASAP7_75t_R g763 ( 
.A(n_2),
.Y(n_763)
);

CKINVDCx5p33_ASAP7_75t_R g764 ( 
.A(n_285),
.Y(n_764)
);

INVx1_ASAP7_75t_L g765 ( 
.A(n_683),
.Y(n_765)
);

INVx1_ASAP7_75t_L g766 ( 
.A(n_722),
.Y(n_766)
);

BUFx10_ASAP7_75t_L g767 ( 
.A(n_665),
.Y(n_767)
);

CKINVDCx5p33_ASAP7_75t_R g768 ( 
.A(n_452),
.Y(n_768)
);

INVx1_ASAP7_75t_L g769 ( 
.A(n_523),
.Y(n_769)
);

CKINVDCx5p33_ASAP7_75t_R g770 ( 
.A(n_707),
.Y(n_770)
);

BUFx2_ASAP7_75t_L g771 ( 
.A(n_36),
.Y(n_771)
);

INVx2_ASAP7_75t_L g772 ( 
.A(n_723),
.Y(n_772)
);

CKINVDCx5p33_ASAP7_75t_R g773 ( 
.A(n_55),
.Y(n_773)
);

CKINVDCx5p33_ASAP7_75t_R g774 ( 
.A(n_727),
.Y(n_774)
);

CKINVDCx5p33_ASAP7_75t_R g775 ( 
.A(n_79),
.Y(n_775)
);

CKINVDCx5p33_ASAP7_75t_R g776 ( 
.A(n_439),
.Y(n_776)
);

INVxp67_ASAP7_75t_L g777 ( 
.A(n_697),
.Y(n_777)
);

CKINVDCx5p33_ASAP7_75t_R g778 ( 
.A(n_167),
.Y(n_778)
);

INVx1_ASAP7_75t_L g779 ( 
.A(n_734),
.Y(n_779)
);

CKINVDCx5p33_ASAP7_75t_R g780 ( 
.A(n_260),
.Y(n_780)
);

CKINVDCx5p33_ASAP7_75t_R g781 ( 
.A(n_475),
.Y(n_781)
);

BUFx3_ASAP7_75t_L g782 ( 
.A(n_638),
.Y(n_782)
);

CKINVDCx5p33_ASAP7_75t_R g783 ( 
.A(n_459),
.Y(n_783)
);

CKINVDCx5p33_ASAP7_75t_R g784 ( 
.A(n_581),
.Y(n_784)
);

INVx2_ASAP7_75t_L g785 ( 
.A(n_398),
.Y(n_785)
);

INVx2_ASAP7_75t_L g786 ( 
.A(n_664),
.Y(n_786)
);

INVx1_ASAP7_75t_L g787 ( 
.A(n_593),
.Y(n_787)
);

CKINVDCx5p33_ASAP7_75t_R g788 ( 
.A(n_661),
.Y(n_788)
);

CKINVDCx5p33_ASAP7_75t_R g789 ( 
.A(n_660),
.Y(n_789)
);

CKINVDCx5p33_ASAP7_75t_R g790 ( 
.A(n_16),
.Y(n_790)
);

BUFx2_ASAP7_75t_L g791 ( 
.A(n_440),
.Y(n_791)
);

CKINVDCx5p33_ASAP7_75t_R g792 ( 
.A(n_42),
.Y(n_792)
);

CKINVDCx5p33_ASAP7_75t_R g793 ( 
.A(n_385),
.Y(n_793)
);

BUFx2_ASAP7_75t_L g794 ( 
.A(n_235),
.Y(n_794)
);

INVx1_ASAP7_75t_SL g795 ( 
.A(n_531),
.Y(n_795)
);

CKINVDCx5p33_ASAP7_75t_R g796 ( 
.A(n_15),
.Y(n_796)
);

BUFx2_ASAP7_75t_L g797 ( 
.A(n_709),
.Y(n_797)
);

CKINVDCx5p33_ASAP7_75t_R g798 ( 
.A(n_27),
.Y(n_798)
);

INVx1_ASAP7_75t_L g799 ( 
.A(n_713),
.Y(n_799)
);

CKINVDCx5p33_ASAP7_75t_R g800 ( 
.A(n_113),
.Y(n_800)
);

INVx1_ASAP7_75t_L g801 ( 
.A(n_625),
.Y(n_801)
);

BUFx6f_ASAP7_75t_L g802 ( 
.A(n_718),
.Y(n_802)
);

CKINVDCx5p33_ASAP7_75t_R g803 ( 
.A(n_579),
.Y(n_803)
);

INVx1_ASAP7_75t_L g804 ( 
.A(n_545),
.Y(n_804)
);

INVx2_ASAP7_75t_L g805 ( 
.A(n_408),
.Y(n_805)
);

CKINVDCx5p33_ASAP7_75t_R g806 ( 
.A(n_674),
.Y(n_806)
);

CKINVDCx5p33_ASAP7_75t_R g807 ( 
.A(n_542),
.Y(n_807)
);

INVx1_ASAP7_75t_L g808 ( 
.A(n_544),
.Y(n_808)
);

INVx1_ASAP7_75t_L g809 ( 
.A(n_736),
.Y(n_809)
);

CKINVDCx16_ASAP7_75t_R g810 ( 
.A(n_367),
.Y(n_810)
);

CKINVDCx5p33_ASAP7_75t_R g811 ( 
.A(n_90),
.Y(n_811)
);

INVx1_ASAP7_75t_L g812 ( 
.A(n_460),
.Y(n_812)
);

CKINVDCx5p33_ASAP7_75t_R g813 ( 
.A(n_635),
.Y(n_813)
);

INVx1_ASAP7_75t_L g814 ( 
.A(n_96),
.Y(n_814)
);

CKINVDCx5p33_ASAP7_75t_R g815 ( 
.A(n_691),
.Y(n_815)
);

INVx1_ASAP7_75t_L g816 ( 
.A(n_506),
.Y(n_816)
);

INVx1_ASAP7_75t_L g817 ( 
.A(n_4),
.Y(n_817)
);

CKINVDCx5p33_ASAP7_75t_R g818 ( 
.A(n_261),
.Y(n_818)
);

CKINVDCx5p33_ASAP7_75t_R g819 ( 
.A(n_394),
.Y(n_819)
);

CKINVDCx5p33_ASAP7_75t_R g820 ( 
.A(n_569),
.Y(n_820)
);

CKINVDCx5p33_ASAP7_75t_R g821 ( 
.A(n_384),
.Y(n_821)
);

BUFx10_ASAP7_75t_L g822 ( 
.A(n_7),
.Y(n_822)
);

INVx1_ASAP7_75t_L g823 ( 
.A(n_183),
.Y(n_823)
);

CKINVDCx5p33_ASAP7_75t_R g824 ( 
.A(n_189),
.Y(n_824)
);

INVx1_ASAP7_75t_L g825 ( 
.A(n_67),
.Y(n_825)
);

CKINVDCx5p33_ASAP7_75t_R g826 ( 
.A(n_721),
.Y(n_826)
);

INVx1_ASAP7_75t_L g827 ( 
.A(n_655),
.Y(n_827)
);

INVx1_ASAP7_75t_L g828 ( 
.A(n_646),
.Y(n_828)
);

CKINVDCx5p33_ASAP7_75t_R g829 ( 
.A(n_288),
.Y(n_829)
);

CKINVDCx20_ASAP7_75t_R g830 ( 
.A(n_614),
.Y(n_830)
);

INVx1_ASAP7_75t_L g831 ( 
.A(n_671),
.Y(n_831)
);

CKINVDCx5p33_ASAP7_75t_R g832 ( 
.A(n_636),
.Y(n_832)
);

CKINVDCx20_ASAP7_75t_R g833 ( 
.A(n_454),
.Y(n_833)
);

CKINVDCx5p33_ASAP7_75t_R g834 ( 
.A(n_726),
.Y(n_834)
);

CKINVDCx5p33_ASAP7_75t_R g835 ( 
.A(n_156),
.Y(n_835)
);

CKINVDCx5p33_ASAP7_75t_R g836 ( 
.A(n_681),
.Y(n_836)
);

INVxp67_ASAP7_75t_L g837 ( 
.A(n_54),
.Y(n_837)
);

CKINVDCx5p33_ASAP7_75t_R g838 ( 
.A(n_693),
.Y(n_838)
);

INVx1_ASAP7_75t_L g839 ( 
.A(n_115),
.Y(n_839)
);

BUFx6f_ASAP7_75t_L g840 ( 
.A(n_474),
.Y(n_840)
);

CKINVDCx5p33_ASAP7_75t_R g841 ( 
.A(n_127),
.Y(n_841)
);

CKINVDCx5p33_ASAP7_75t_R g842 ( 
.A(n_323),
.Y(n_842)
);

CKINVDCx5p33_ASAP7_75t_R g843 ( 
.A(n_657),
.Y(n_843)
);

CKINVDCx5p33_ASAP7_75t_R g844 ( 
.A(n_316),
.Y(n_844)
);

INVx1_ASAP7_75t_L g845 ( 
.A(n_355),
.Y(n_845)
);

CKINVDCx5p33_ASAP7_75t_R g846 ( 
.A(n_31),
.Y(n_846)
);

CKINVDCx20_ASAP7_75t_R g847 ( 
.A(n_731),
.Y(n_847)
);

INVx1_ASAP7_75t_L g848 ( 
.A(n_382),
.Y(n_848)
);

CKINVDCx5p33_ASAP7_75t_R g849 ( 
.A(n_69),
.Y(n_849)
);

CKINVDCx5p33_ASAP7_75t_R g850 ( 
.A(n_392),
.Y(n_850)
);

CKINVDCx5p33_ASAP7_75t_R g851 ( 
.A(n_663),
.Y(n_851)
);

INVx1_ASAP7_75t_L g852 ( 
.A(n_642),
.Y(n_852)
);

CKINVDCx16_ASAP7_75t_R g853 ( 
.A(n_292),
.Y(n_853)
);

CKINVDCx5p33_ASAP7_75t_R g854 ( 
.A(n_714),
.Y(n_854)
);

INVx1_ASAP7_75t_L g855 ( 
.A(n_733),
.Y(n_855)
);

CKINVDCx5p33_ASAP7_75t_R g856 ( 
.A(n_574),
.Y(n_856)
);

INVx2_ASAP7_75t_L g857 ( 
.A(n_608),
.Y(n_857)
);

INVx1_ASAP7_75t_L g858 ( 
.A(n_602),
.Y(n_858)
);

CKINVDCx5p33_ASAP7_75t_R g859 ( 
.A(n_274),
.Y(n_859)
);

CKINVDCx5p33_ASAP7_75t_R g860 ( 
.A(n_705),
.Y(n_860)
);

CKINVDCx5p33_ASAP7_75t_R g861 ( 
.A(n_730),
.Y(n_861)
);

BUFx6f_ASAP7_75t_L g862 ( 
.A(n_41),
.Y(n_862)
);

CKINVDCx5p33_ASAP7_75t_R g863 ( 
.A(n_738),
.Y(n_863)
);

CKINVDCx5p33_ASAP7_75t_R g864 ( 
.A(n_552),
.Y(n_864)
);

CKINVDCx5p33_ASAP7_75t_R g865 ( 
.A(n_18),
.Y(n_865)
);

BUFx3_ASAP7_75t_L g866 ( 
.A(n_711),
.Y(n_866)
);

BUFx6f_ASAP7_75t_L g867 ( 
.A(n_411),
.Y(n_867)
);

CKINVDCx5p33_ASAP7_75t_R g868 ( 
.A(n_293),
.Y(n_868)
);

CKINVDCx5p33_ASAP7_75t_R g869 ( 
.A(n_712),
.Y(n_869)
);

INVx2_ASAP7_75t_L g870 ( 
.A(n_370),
.Y(n_870)
);

BUFx10_ASAP7_75t_L g871 ( 
.A(n_643),
.Y(n_871)
);

CKINVDCx5p33_ASAP7_75t_R g872 ( 
.A(n_652),
.Y(n_872)
);

INVx2_ASAP7_75t_L g873 ( 
.A(n_241),
.Y(n_873)
);

CKINVDCx5p33_ASAP7_75t_R g874 ( 
.A(n_667),
.Y(n_874)
);

CKINVDCx5p33_ASAP7_75t_R g875 ( 
.A(n_133),
.Y(n_875)
);

CKINVDCx5p33_ASAP7_75t_R g876 ( 
.A(n_3),
.Y(n_876)
);

INVx1_ASAP7_75t_L g877 ( 
.A(n_534),
.Y(n_877)
);

INVx1_ASAP7_75t_SL g878 ( 
.A(n_673),
.Y(n_878)
);

INVx2_ASAP7_75t_SL g879 ( 
.A(n_351),
.Y(n_879)
);

CKINVDCx5p33_ASAP7_75t_R g880 ( 
.A(n_729),
.Y(n_880)
);

INVxp67_ASAP7_75t_SL g881 ( 
.A(n_266),
.Y(n_881)
);

CKINVDCx20_ASAP7_75t_R g882 ( 
.A(n_567),
.Y(n_882)
);

INVx1_ASAP7_75t_L g883 ( 
.A(n_696),
.Y(n_883)
);

CKINVDCx5p33_ASAP7_75t_R g884 ( 
.A(n_530),
.Y(n_884)
);

BUFx2_ASAP7_75t_L g885 ( 
.A(n_447),
.Y(n_885)
);

CKINVDCx5p33_ASAP7_75t_R g886 ( 
.A(n_214),
.Y(n_886)
);

BUFx6f_ASAP7_75t_L g887 ( 
.A(n_155),
.Y(n_887)
);

CKINVDCx5p33_ASAP7_75t_R g888 ( 
.A(n_694),
.Y(n_888)
);

INVx1_ASAP7_75t_L g889 ( 
.A(n_689),
.Y(n_889)
);

INVx1_ASAP7_75t_L g890 ( 
.A(n_128),
.Y(n_890)
);

INVx1_ASAP7_75t_L g891 ( 
.A(n_670),
.Y(n_891)
);

BUFx6f_ASAP7_75t_L g892 ( 
.A(n_628),
.Y(n_892)
);

INVx2_ASAP7_75t_L g893 ( 
.A(n_114),
.Y(n_893)
);

CKINVDCx5p33_ASAP7_75t_R g894 ( 
.A(n_505),
.Y(n_894)
);

CKINVDCx5p33_ASAP7_75t_R g895 ( 
.A(n_326),
.Y(n_895)
);

CKINVDCx5p33_ASAP7_75t_R g896 ( 
.A(n_423),
.Y(n_896)
);

CKINVDCx5p33_ASAP7_75t_R g897 ( 
.A(n_605),
.Y(n_897)
);

INVx1_ASAP7_75t_L g898 ( 
.A(n_368),
.Y(n_898)
);

INVx1_ASAP7_75t_SL g899 ( 
.A(n_659),
.Y(n_899)
);

CKINVDCx20_ASAP7_75t_R g900 ( 
.A(n_662),
.Y(n_900)
);

CKINVDCx20_ASAP7_75t_R g901 ( 
.A(n_8),
.Y(n_901)
);

CKINVDCx20_ASAP7_75t_R g902 ( 
.A(n_379),
.Y(n_902)
);

CKINVDCx5p33_ASAP7_75t_R g903 ( 
.A(n_717),
.Y(n_903)
);

CKINVDCx5p33_ASAP7_75t_R g904 ( 
.A(n_59),
.Y(n_904)
);

CKINVDCx5p33_ASAP7_75t_R g905 ( 
.A(n_528),
.Y(n_905)
);

CKINVDCx5p33_ASAP7_75t_R g906 ( 
.A(n_383),
.Y(n_906)
);

CKINVDCx5p33_ASAP7_75t_R g907 ( 
.A(n_613),
.Y(n_907)
);

INVx1_ASAP7_75t_L g908 ( 
.A(n_572),
.Y(n_908)
);

INVx1_ASAP7_75t_L g909 ( 
.A(n_716),
.Y(n_909)
);

BUFx3_ASAP7_75t_L g910 ( 
.A(n_159),
.Y(n_910)
);

BUFx6f_ASAP7_75t_L g911 ( 
.A(n_617),
.Y(n_911)
);

CKINVDCx20_ASAP7_75t_R g912 ( 
.A(n_417),
.Y(n_912)
);

CKINVDCx5p33_ASAP7_75t_R g913 ( 
.A(n_704),
.Y(n_913)
);

CKINVDCx5p33_ASAP7_75t_R g914 ( 
.A(n_517),
.Y(n_914)
);

INVx1_ASAP7_75t_L g915 ( 
.A(n_216),
.Y(n_915)
);

INVx1_ASAP7_75t_L g916 ( 
.A(n_649),
.Y(n_916)
);

CKINVDCx5p33_ASAP7_75t_R g917 ( 
.A(n_735),
.Y(n_917)
);

INVx1_ASAP7_75t_L g918 ( 
.A(n_328),
.Y(n_918)
);

INVx1_ASAP7_75t_L g919 ( 
.A(n_60),
.Y(n_919)
);

CKINVDCx5p33_ASAP7_75t_R g920 ( 
.A(n_546),
.Y(n_920)
);

CKINVDCx5p33_ASAP7_75t_R g921 ( 
.A(n_177),
.Y(n_921)
);

INVx1_ASAP7_75t_L g922 ( 
.A(n_17),
.Y(n_922)
);

BUFx10_ASAP7_75t_L g923 ( 
.A(n_487),
.Y(n_923)
);

CKINVDCx5p33_ASAP7_75t_R g924 ( 
.A(n_641),
.Y(n_924)
);

INVx1_ASAP7_75t_L g925 ( 
.A(n_185),
.Y(n_925)
);

INVx1_ASAP7_75t_L g926 ( 
.A(n_174),
.Y(n_926)
);

INVx1_ASAP7_75t_L g927 ( 
.A(n_467),
.Y(n_927)
);

CKINVDCx5p33_ASAP7_75t_R g928 ( 
.A(n_241),
.Y(n_928)
);

CKINVDCx5p33_ASAP7_75t_R g929 ( 
.A(n_644),
.Y(n_929)
);

INVx1_ASAP7_75t_L g930 ( 
.A(n_684),
.Y(n_930)
);

CKINVDCx5p33_ASAP7_75t_R g931 ( 
.A(n_371),
.Y(n_931)
);

CKINVDCx20_ASAP7_75t_R g932 ( 
.A(n_267),
.Y(n_932)
);

INVx1_ASAP7_75t_L g933 ( 
.A(n_204),
.Y(n_933)
);

CKINVDCx5p33_ASAP7_75t_R g934 ( 
.A(n_688),
.Y(n_934)
);

CKINVDCx20_ASAP7_75t_R g935 ( 
.A(n_580),
.Y(n_935)
);

INVx1_ASAP7_75t_L g936 ( 
.A(n_543),
.Y(n_936)
);

BUFx10_ASAP7_75t_L g937 ( 
.A(n_724),
.Y(n_937)
);

INVx1_ASAP7_75t_L g938 ( 
.A(n_695),
.Y(n_938)
);

CKINVDCx5p33_ASAP7_75t_R g939 ( 
.A(n_529),
.Y(n_939)
);

INVx1_ASAP7_75t_L g940 ( 
.A(n_360),
.Y(n_940)
);

CKINVDCx5p33_ASAP7_75t_R g941 ( 
.A(n_703),
.Y(n_941)
);

CKINVDCx16_ASAP7_75t_R g942 ( 
.A(n_682),
.Y(n_942)
);

CKINVDCx5p33_ASAP7_75t_R g943 ( 
.A(n_143),
.Y(n_943)
);

CKINVDCx5p33_ASAP7_75t_R g944 ( 
.A(n_218),
.Y(n_944)
);

CKINVDCx5p33_ASAP7_75t_R g945 ( 
.A(n_706),
.Y(n_945)
);

INVx2_ASAP7_75t_SL g946 ( 
.A(n_653),
.Y(n_946)
);

CKINVDCx5p33_ASAP7_75t_R g947 ( 
.A(n_537),
.Y(n_947)
);

CKINVDCx5p33_ASAP7_75t_R g948 ( 
.A(n_248),
.Y(n_948)
);

INVx1_ASAP7_75t_L g949 ( 
.A(n_335),
.Y(n_949)
);

CKINVDCx5p33_ASAP7_75t_R g950 ( 
.A(n_318),
.Y(n_950)
);

CKINVDCx5p33_ASAP7_75t_R g951 ( 
.A(n_692),
.Y(n_951)
);

INVx2_ASAP7_75t_SL g952 ( 
.A(n_676),
.Y(n_952)
);

INVx1_ASAP7_75t_L g953 ( 
.A(n_550),
.Y(n_953)
);

CKINVDCx5p33_ASAP7_75t_R g954 ( 
.A(n_620),
.Y(n_954)
);

CKINVDCx5p33_ASAP7_75t_R g955 ( 
.A(n_425),
.Y(n_955)
);

CKINVDCx5p33_ASAP7_75t_R g956 ( 
.A(n_669),
.Y(n_956)
);

INVx1_ASAP7_75t_L g957 ( 
.A(n_316),
.Y(n_957)
);

INVx2_ASAP7_75t_L g958 ( 
.A(n_647),
.Y(n_958)
);

CKINVDCx20_ASAP7_75t_R g959 ( 
.A(n_395),
.Y(n_959)
);

INVx1_ASAP7_75t_L g960 ( 
.A(n_334),
.Y(n_960)
);

INVx1_ASAP7_75t_L g961 ( 
.A(n_677),
.Y(n_961)
);

INVx1_ASAP7_75t_L g962 ( 
.A(n_110),
.Y(n_962)
);

CKINVDCx5p33_ASAP7_75t_R g963 ( 
.A(n_720),
.Y(n_963)
);

BUFx6f_ASAP7_75t_L g964 ( 
.A(n_701),
.Y(n_964)
);

CKINVDCx20_ASAP7_75t_R g965 ( 
.A(n_640),
.Y(n_965)
);

CKINVDCx5p33_ASAP7_75t_R g966 ( 
.A(n_612),
.Y(n_966)
);

CKINVDCx5p33_ASAP7_75t_R g967 ( 
.A(n_107),
.Y(n_967)
);

BUFx10_ASAP7_75t_L g968 ( 
.A(n_632),
.Y(n_968)
);

CKINVDCx5p33_ASAP7_75t_R g969 ( 
.A(n_363),
.Y(n_969)
);

CKINVDCx5p33_ASAP7_75t_R g970 ( 
.A(n_686),
.Y(n_970)
);

CKINVDCx5p33_ASAP7_75t_R g971 ( 
.A(n_700),
.Y(n_971)
);

INVx2_ASAP7_75t_L g972 ( 
.A(n_1),
.Y(n_972)
);

INVx1_ASAP7_75t_SL g973 ( 
.A(n_685),
.Y(n_973)
);

CKINVDCx5p33_ASAP7_75t_R g974 ( 
.A(n_648),
.Y(n_974)
);

CKINVDCx5p33_ASAP7_75t_R g975 ( 
.A(n_257),
.Y(n_975)
);

BUFx2_ASAP7_75t_L g976 ( 
.A(n_189),
.Y(n_976)
);

BUFx3_ASAP7_75t_L g977 ( 
.A(n_47),
.Y(n_977)
);

CKINVDCx5p33_ASAP7_75t_R g978 ( 
.A(n_715),
.Y(n_978)
);

CKINVDCx5p33_ASAP7_75t_R g979 ( 
.A(n_699),
.Y(n_979)
);

INVx1_ASAP7_75t_L g980 ( 
.A(n_651),
.Y(n_980)
);

CKINVDCx5p33_ASAP7_75t_R g981 ( 
.A(n_388),
.Y(n_981)
);

INVx1_ASAP7_75t_L g982 ( 
.A(n_133),
.Y(n_982)
);

CKINVDCx20_ASAP7_75t_R g983 ( 
.A(n_339),
.Y(n_983)
);

CKINVDCx5p33_ASAP7_75t_R g984 ( 
.A(n_274),
.Y(n_984)
);

CKINVDCx20_ASAP7_75t_R g985 ( 
.A(n_86),
.Y(n_985)
);

CKINVDCx5p33_ASAP7_75t_R g986 ( 
.A(n_177),
.Y(n_986)
);

INVx2_ASAP7_75t_L g987 ( 
.A(n_373),
.Y(n_987)
);

CKINVDCx5p33_ASAP7_75t_R g988 ( 
.A(n_16),
.Y(n_988)
);

CKINVDCx5p33_ASAP7_75t_R g989 ( 
.A(n_675),
.Y(n_989)
);

CKINVDCx5p33_ASAP7_75t_R g990 ( 
.A(n_728),
.Y(n_990)
);

INVx1_ASAP7_75t_L g991 ( 
.A(n_312),
.Y(n_991)
);

CKINVDCx5p33_ASAP7_75t_R g992 ( 
.A(n_247),
.Y(n_992)
);

CKINVDCx5p33_ASAP7_75t_R g993 ( 
.A(n_208),
.Y(n_993)
);

CKINVDCx5p33_ASAP7_75t_R g994 ( 
.A(n_111),
.Y(n_994)
);

INVx1_ASAP7_75t_L g995 ( 
.A(n_654),
.Y(n_995)
);

CKINVDCx5p33_ASAP7_75t_R g996 ( 
.A(n_672),
.Y(n_996)
);

INVx1_ASAP7_75t_L g997 ( 
.A(n_58),
.Y(n_997)
);

INVx1_ASAP7_75t_SL g998 ( 
.A(n_719),
.Y(n_998)
);

INVx2_ASAP7_75t_SL g999 ( 
.A(n_658),
.Y(n_999)
);

CKINVDCx5p33_ASAP7_75t_R g1000 ( 
.A(n_211),
.Y(n_1000)
);

HB1xp67_ASAP7_75t_L g1001 ( 
.A(n_98),
.Y(n_1001)
);

CKINVDCx5p33_ASAP7_75t_R g1002 ( 
.A(n_215),
.Y(n_1002)
);

BUFx6f_ASAP7_75t_L g1003 ( 
.A(n_253),
.Y(n_1003)
);

INVx1_ASAP7_75t_L g1004 ( 
.A(n_645),
.Y(n_1004)
);

CKINVDCx5p33_ASAP7_75t_R g1005 ( 
.A(n_21),
.Y(n_1005)
);

INVxp67_ASAP7_75t_L g1006 ( 
.A(n_680),
.Y(n_1006)
);

INVx1_ASAP7_75t_L g1007 ( 
.A(n_639),
.Y(n_1007)
);

CKINVDCx5p33_ASAP7_75t_R g1008 ( 
.A(n_466),
.Y(n_1008)
);

INVx1_ASAP7_75t_L g1009 ( 
.A(n_633),
.Y(n_1009)
);

CKINVDCx5p33_ASAP7_75t_R g1010 ( 
.A(n_592),
.Y(n_1010)
);

INVx1_ASAP7_75t_L g1011 ( 
.A(n_442),
.Y(n_1011)
);

INVx1_ASAP7_75t_L g1012 ( 
.A(n_389),
.Y(n_1012)
);

CKINVDCx5p33_ASAP7_75t_R g1013 ( 
.A(n_687),
.Y(n_1013)
);

CKINVDCx5p33_ASAP7_75t_R g1014 ( 
.A(n_102),
.Y(n_1014)
);

CKINVDCx5p33_ASAP7_75t_R g1015 ( 
.A(n_284),
.Y(n_1015)
);

INVx1_ASAP7_75t_L g1016 ( 
.A(n_305),
.Y(n_1016)
);

INVx1_ASAP7_75t_L g1017 ( 
.A(n_623),
.Y(n_1017)
);

CKINVDCx5p33_ASAP7_75t_R g1018 ( 
.A(n_381),
.Y(n_1018)
);

INVx2_ASAP7_75t_L g1019 ( 
.A(n_516),
.Y(n_1019)
);

CKINVDCx5p33_ASAP7_75t_R g1020 ( 
.A(n_89),
.Y(n_1020)
);

CKINVDCx5p33_ASAP7_75t_R g1021 ( 
.A(n_710),
.Y(n_1021)
);

CKINVDCx5p33_ASAP7_75t_R g1022 ( 
.A(n_463),
.Y(n_1022)
);

INVx2_ASAP7_75t_L g1023 ( 
.A(n_702),
.Y(n_1023)
);

INVx1_ASAP7_75t_L g1024 ( 
.A(n_725),
.Y(n_1024)
);

CKINVDCx5p33_ASAP7_75t_R g1025 ( 
.A(n_634),
.Y(n_1025)
);

CKINVDCx5p33_ASAP7_75t_R g1026 ( 
.A(n_656),
.Y(n_1026)
);

BUFx3_ASAP7_75t_L g1027 ( 
.A(n_387),
.Y(n_1027)
);

INVx2_ASAP7_75t_SL g1028 ( 
.A(n_323),
.Y(n_1028)
);

CKINVDCx5p33_ASAP7_75t_R g1029 ( 
.A(n_165),
.Y(n_1029)
);

INVx1_ASAP7_75t_L g1030 ( 
.A(n_690),
.Y(n_1030)
);

INVx1_ASAP7_75t_L g1031 ( 
.A(n_862),
.Y(n_1031)
);

INVxp67_ASAP7_75t_L g1032 ( 
.A(n_771),
.Y(n_1032)
);

NOR2xp33_ASAP7_75t_L g1033 ( 
.A(n_791),
.B(n_1),
.Y(n_1033)
);

INVx1_ASAP7_75t_L g1034 ( 
.A(n_862),
.Y(n_1034)
);

CKINVDCx5p33_ASAP7_75t_R g1035 ( 
.A(n_743),
.Y(n_1035)
);

CKINVDCx5p33_ASAP7_75t_R g1036 ( 
.A(n_744),
.Y(n_1036)
);

INVx1_ASAP7_75t_L g1037 ( 
.A(n_862),
.Y(n_1037)
);

CKINVDCx5p33_ASAP7_75t_R g1038 ( 
.A(n_751),
.Y(n_1038)
);

CKINVDCx16_ASAP7_75t_R g1039 ( 
.A(n_747),
.Y(n_1039)
);

CKINVDCx5p33_ASAP7_75t_R g1040 ( 
.A(n_752),
.Y(n_1040)
);

CKINVDCx20_ASAP7_75t_R g1041 ( 
.A(n_748),
.Y(n_1041)
);

CKINVDCx20_ASAP7_75t_R g1042 ( 
.A(n_750),
.Y(n_1042)
);

CKINVDCx5p33_ASAP7_75t_R g1043 ( 
.A(n_754),
.Y(n_1043)
);

INVx1_ASAP7_75t_L g1044 ( 
.A(n_887),
.Y(n_1044)
);

CKINVDCx5p33_ASAP7_75t_R g1045 ( 
.A(n_757),
.Y(n_1045)
);

CKINVDCx5p33_ASAP7_75t_R g1046 ( 
.A(n_768),
.Y(n_1046)
);

INVx1_ASAP7_75t_L g1047 ( 
.A(n_887),
.Y(n_1047)
);

CKINVDCx5p33_ASAP7_75t_R g1048 ( 
.A(n_770),
.Y(n_1048)
);

INVx1_ASAP7_75t_L g1049 ( 
.A(n_887),
.Y(n_1049)
);

INVx1_ASAP7_75t_L g1050 ( 
.A(n_1003),
.Y(n_1050)
);

INVx1_ASAP7_75t_L g1051 ( 
.A(n_1003),
.Y(n_1051)
);

CKINVDCx5p33_ASAP7_75t_R g1052 ( 
.A(n_774),
.Y(n_1052)
);

OR2x2_ASAP7_75t_L g1053 ( 
.A(n_794),
.B(n_0),
.Y(n_1053)
);

INVxp67_ASAP7_75t_L g1054 ( 
.A(n_976),
.Y(n_1054)
);

NOR2xp33_ASAP7_75t_L g1055 ( 
.A(n_797),
.B(n_2),
.Y(n_1055)
);

INVxp67_ASAP7_75t_SL g1056 ( 
.A(n_885),
.Y(n_1056)
);

HB1xp67_ASAP7_75t_L g1057 ( 
.A(n_853),
.Y(n_1057)
);

INVx1_ASAP7_75t_L g1058 ( 
.A(n_1003),
.Y(n_1058)
);

INVx1_ASAP7_75t_L g1059 ( 
.A(n_910),
.Y(n_1059)
);

INVx3_ASAP7_75t_L g1060 ( 
.A(n_977),
.Y(n_1060)
);

INVx1_ASAP7_75t_L g1061 ( 
.A(n_1031),
.Y(n_1061)
);

INVx3_ASAP7_75t_L g1062 ( 
.A(n_1034),
.Y(n_1062)
);

NAND2xp5_ASAP7_75t_L g1063 ( 
.A(n_1035),
.B(n_758),
.Y(n_1063)
);

INVx1_ASAP7_75t_L g1064 ( 
.A(n_1037),
.Y(n_1064)
);

AND2x2_ASAP7_75t_L g1065 ( 
.A(n_1056),
.B(n_759),
.Y(n_1065)
);

AND2x2_ASAP7_75t_L g1066 ( 
.A(n_1036),
.B(n_810),
.Y(n_1066)
);

OA21x2_ASAP7_75t_L g1067 ( 
.A1(n_1044),
.A2(n_765),
.B(n_742),
.Y(n_1067)
);

INVx1_ASAP7_75t_L g1068 ( 
.A(n_1047),
.Y(n_1068)
);

BUFx6f_ASAP7_75t_L g1069 ( 
.A(n_1049),
.Y(n_1069)
);

INVx3_ASAP7_75t_L g1070 ( 
.A(n_1050),
.Y(n_1070)
);

INVx1_ASAP7_75t_L g1071 ( 
.A(n_1051),
.Y(n_1071)
);

CKINVDCx5p33_ASAP7_75t_R g1072 ( 
.A(n_1038),
.Y(n_1072)
);

INVx1_ASAP7_75t_L g1073 ( 
.A(n_1058),
.Y(n_1073)
);

AND2x4_ASAP7_75t_L g1074 ( 
.A(n_1032),
.B(n_749),
.Y(n_1074)
);

INVx2_ASAP7_75t_L g1075 ( 
.A(n_1060),
.Y(n_1075)
);

INVx1_ASAP7_75t_L g1076 ( 
.A(n_1059),
.Y(n_1076)
);

INVx4_ASAP7_75t_L g1077 ( 
.A(n_1040),
.Y(n_1077)
);

HB1xp67_ASAP7_75t_L g1078 ( 
.A(n_1057),
.Y(n_1078)
);

HB1xp67_ASAP7_75t_L g1079 ( 
.A(n_1039),
.Y(n_1079)
);

CKINVDCx5p33_ASAP7_75t_R g1080 ( 
.A(n_1043),
.Y(n_1080)
);

INVx1_ASAP7_75t_L g1081 ( 
.A(n_1060),
.Y(n_1081)
);

NAND2xp5_ASAP7_75t_SL g1082 ( 
.A(n_1033),
.B(n_942),
.Y(n_1082)
);

OAI21x1_ASAP7_75t_L g1083 ( 
.A1(n_1053),
.A2(n_755),
.B(n_745),
.Y(n_1083)
);

INVx1_ASAP7_75t_L g1084 ( 
.A(n_1045),
.Y(n_1084)
);

INVx2_ASAP7_75t_L g1085 ( 
.A(n_1046),
.Y(n_1085)
);

INVx1_ASAP7_75t_L g1086 ( 
.A(n_1048),
.Y(n_1086)
);

HB1xp67_ASAP7_75t_L g1087 ( 
.A(n_1052),
.Y(n_1087)
);

INVx2_ASAP7_75t_L g1088 ( 
.A(n_1054),
.Y(n_1088)
);

INVx3_ASAP7_75t_L g1089 ( 
.A(n_1055),
.Y(n_1089)
);

NAND2xp5_ASAP7_75t_L g1090 ( 
.A(n_1041),
.B(n_879),
.Y(n_1090)
);

INVx1_ASAP7_75t_L g1091 ( 
.A(n_1042),
.Y(n_1091)
);

INVx3_ASAP7_75t_L g1092 ( 
.A(n_1069),
.Y(n_1092)
);

NAND2xp33_ASAP7_75t_L g1093 ( 
.A(n_1089),
.B(n_802),
.Y(n_1093)
);

INVx2_ASAP7_75t_L g1094 ( 
.A(n_1069),
.Y(n_1094)
);

OAI22xp5_ASAP7_75t_L g1095 ( 
.A1(n_1089),
.A2(n_837),
.B1(n_881),
.B2(n_1001),
.Y(n_1095)
);

AND2x2_ASAP7_75t_L g1096 ( 
.A(n_1065),
.B(n_760),
.Y(n_1096)
);

INVx3_ASAP7_75t_L g1097 ( 
.A(n_1069),
.Y(n_1097)
);

AND2x2_ASAP7_75t_L g1098 ( 
.A(n_1075),
.B(n_1028),
.Y(n_1098)
);

AO21x2_ASAP7_75t_L g1099 ( 
.A1(n_1063),
.A2(n_1083),
.B(n_1084),
.Y(n_1099)
);

CKINVDCx5p33_ASAP7_75t_R g1100 ( 
.A(n_1072),
.Y(n_1100)
);

INVx1_ASAP7_75t_L g1101 ( 
.A(n_1076),
.Y(n_1101)
);

INVx1_ASAP7_75t_SL g1102 ( 
.A(n_1079),
.Y(n_1102)
);

INVxp33_ASAP7_75t_L g1103 ( 
.A(n_1078),
.Y(n_1103)
);

INVx2_ASAP7_75t_L g1104 ( 
.A(n_1061),
.Y(n_1104)
);

INVx2_ASAP7_75t_L g1105 ( 
.A(n_1064),
.Y(n_1105)
);

AND2x6_ASAP7_75t_L g1106 ( 
.A(n_1085),
.B(n_802),
.Y(n_1106)
);

INVx1_ASAP7_75t_L g1107 ( 
.A(n_1068),
.Y(n_1107)
);

AND2x6_ASAP7_75t_L g1108 ( 
.A(n_1086),
.B(n_802),
.Y(n_1108)
);

NAND2xp5_ASAP7_75t_SL g1109 ( 
.A(n_1066),
.B(n_767),
.Y(n_1109)
);

INVx1_ASAP7_75t_L g1110 ( 
.A(n_1071),
.Y(n_1110)
);

AOI22xp5_ASAP7_75t_L g1111 ( 
.A1(n_1082),
.A2(n_830),
.B1(n_833),
.B2(n_756),
.Y(n_1111)
);

INVx2_ASAP7_75t_L g1112 ( 
.A(n_1073),
.Y(n_1112)
);

BUFx6f_ASAP7_75t_L g1113 ( 
.A(n_1062),
.Y(n_1113)
);

INVx2_ASAP7_75t_L g1114 ( 
.A(n_1062),
.Y(n_1114)
);

NAND2xp5_ASAP7_75t_SL g1115 ( 
.A(n_1080),
.B(n_767),
.Y(n_1115)
);

INVx1_ASAP7_75t_L g1116 ( 
.A(n_1081),
.Y(n_1116)
);

INVx2_ASAP7_75t_L g1117 ( 
.A(n_1070),
.Y(n_1117)
);

INVx3_ASAP7_75t_L g1118 ( 
.A(n_1070),
.Y(n_1118)
);

INVx4_ASAP7_75t_L g1119 ( 
.A(n_1077),
.Y(n_1119)
);

INVx1_ASAP7_75t_L g1120 ( 
.A(n_1067),
.Y(n_1120)
);

INVx2_ASAP7_75t_L g1121 ( 
.A(n_1067),
.Y(n_1121)
);

AND2x2_ASAP7_75t_L g1122 ( 
.A(n_1074),
.B(n_814),
.Y(n_1122)
);

INVx3_ASAP7_75t_L g1123 ( 
.A(n_1074),
.Y(n_1123)
);

INVx1_ASAP7_75t_L g1124 ( 
.A(n_1088),
.Y(n_1124)
);

BUFx6f_ASAP7_75t_L g1125 ( 
.A(n_1090),
.Y(n_1125)
);

NAND2xp5_ASAP7_75t_L g1126 ( 
.A(n_1077),
.B(n_946),
.Y(n_1126)
);

AOI22xp33_ASAP7_75t_L g1127 ( 
.A1(n_1087),
.A2(n_893),
.B1(n_972),
.B2(n_873),
.Y(n_1127)
);

NOR2xp33_ASAP7_75t_L g1128 ( 
.A(n_1091),
.B(n_795),
.Y(n_1128)
);

INVx1_ASAP7_75t_L g1129 ( 
.A(n_1076),
.Y(n_1129)
);

OR2x6_ASAP7_75t_L g1130 ( 
.A(n_1079),
.B(n_817),
.Y(n_1130)
);

AND2x4_ASAP7_75t_L g1131 ( 
.A(n_1085),
.B(n_847),
.Y(n_1131)
);

INVx2_ASAP7_75t_L g1132 ( 
.A(n_1069),
.Y(n_1132)
);

INVx4_ASAP7_75t_L g1133 ( 
.A(n_1072),
.Y(n_1133)
);

BUFx2_ASAP7_75t_L g1134 ( 
.A(n_1079),
.Y(n_1134)
);

BUFx6f_ASAP7_75t_L g1135 ( 
.A(n_1069),
.Y(n_1135)
);

INVx1_ASAP7_75t_SL g1136 ( 
.A(n_1079),
.Y(n_1136)
);

OAI221xp5_ASAP7_75t_L g1137 ( 
.A1(n_1127),
.A2(n_839),
.B1(n_890),
.B2(n_825),
.C(n_823),
.Y(n_1137)
);

INVx1_ASAP7_75t_L g1138 ( 
.A(n_1107),
.Y(n_1138)
);

INVx1_ASAP7_75t_L g1139 ( 
.A(n_1110),
.Y(n_1139)
);

OAI221xp5_ASAP7_75t_L g1140 ( 
.A1(n_1095),
.A2(n_919),
.B1(n_922),
.B2(n_918),
.C(n_915),
.Y(n_1140)
);

NOR2xp67_ASAP7_75t_L g1141 ( 
.A(n_1133),
.B(n_777),
.Y(n_1141)
);

CKINVDCx5p33_ASAP7_75t_R g1142 ( 
.A(n_1100),
.Y(n_1142)
);

INVxp67_ASAP7_75t_L g1143 ( 
.A(n_1128),
.Y(n_1143)
);

INVx1_ASAP7_75t_L g1144 ( 
.A(n_1124),
.Y(n_1144)
);

BUFx8_ASAP7_75t_L g1145 ( 
.A(n_1134),
.Y(n_1145)
);

BUFx2_ASAP7_75t_L g1146 ( 
.A(n_1102),
.Y(n_1146)
);

AND2x2_ASAP7_75t_L g1147 ( 
.A(n_1096),
.B(n_822),
.Y(n_1147)
);

INVx1_ASAP7_75t_L g1148 ( 
.A(n_1101),
.Y(n_1148)
);

INVx1_ASAP7_75t_L g1149 ( 
.A(n_1129),
.Y(n_1149)
);

INVx1_ASAP7_75t_L g1150 ( 
.A(n_1116),
.Y(n_1150)
);

OR2x6_ASAP7_75t_L g1151 ( 
.A(n_1130),
.B(n_925),
.Y(n_1151)
);

INVx1_ASAP7_75t_L g1152 ( 
.A(n_1114),
.Y(n_1152)
);

INVx1_ASAP7_75t_L g1153 ( 
.A(n_1117),
.Y(n_1153)
);

INVx1_ASAP7_75t_L g1154 ( 
.A(n_1104),
.Y(n_1154)
);

OAI22xp33_ASAP7_75t_SL g1155 ( 
.A1(n_1109),
.A2(n_1006),
.B1(n_1030),
.B2(n_1024),
.Y(n_1155)
);

AND2x2_ASAP7_75t_L g1156 ( 
.A(n_1096),
.B(n_822),
.Y(n_1156)
);

AND3x1_ASAP7_75t_L g1157 ( 
.A(n_1111),
.B(n_933),
.C(n_926),
.Y(n_1157)
);

AND2x6_ASAP7_75t_L g1158 ( 
.A(n_1120),
.B(n_766),
.Y(n_1158)
);

INVx1_ASAP7_75t_L g1159 ( 
.A(n_1105),
.Y(n_1159)
);

AO22x2_ASAP7_75t_L g1160 ( 
.A1(n_1136),
.A2(n_997),
.B1(n_1016),
.B2(n_962),
.Y(n_1160)
);

INVx2_ASAP7_75t_L g1161 ( 
.A(n_1112),
.Y(n_1161)
);

INVx2_ASAP7_75t_SL g1162 ( 
.A(n_1125),
.Y(n_1162)
);

INVx1_ASAP7_75t_L g1163 ( 
.A(n_1118),
.Y(n_1163)
);

INVx1_ASAP7_75t_L g1164 ( 
.A(n_1098),
.Y(n_1164)
);

INVx1_ASAP7_75t_L g1165 ( 
.A(n_1098),
.Y(n_1165)
);

INVx1_ASAP7_75t_L g1166 ( 
.A(n_1123),
.Y(n_1166)
);

INVx1_ASAP7_75t_L g1167 ( 
.A(n_1113),
.Y(n_1167)
);

AND2x4_ASAP7_75t_L g1168 ( 
.A(n_1122),
.B(n_949),
.Y(n_1168)
);

INVx1_ASAP7_75t_L g1169 ( 
.A(n_1113),
.Y(n_1169)
);

NAND2x1p5_ASAP7_75t_L g1170 ( 
.A(n_1119),
.B(n_782),
.Y(n_1170)
);

AOI22xp5_ASAP7_75t_L g1171 ( 
.A1(n_1125),
.A2(n_882),
.B1(n_902),
.B2(n_900),
.Y(n_1171)
);

INVx1_ASAP7_75t_L g1172 ( 
.A(n_1122),
.Y(n_1172)
);

OAI221xp5_ASAP7_75t_L g1173 ( 
.A1(n_1126),
.A2(n_957),
.B1(n_991),
.B2(n_982),
.C(n_960),
.Y(n_1173)
);

NAND2x1p5_ASAP7_75t_L g1174 ( 
.A(n_1135),
.B(n_866),
.Y(n_1174)
);

AO22x2_ASAP7_75t_L g1175 ( 
.A1(n_1115),
.A2(n_973),
.B1(n_998),
.B2(n_878),
.Y(n_1175)
);

INVx2_ASAP7_75t_L g1176 ( 
.A(n_1135),
.Y(n_1176)
);

BUFx2_ASAP7_75t_L g1177 ( 
.A(n_1131),
.Y(n_1177)
);

BUFx6f_ASAP7_75t_SL g1178 ( 
.A(n_1130),
.Y(n_1178)
);

INVx1_ASAP7_75t_L g1179 ( 
.A(n_1094),
.Y(n_1179)
);

INVx2_ASAP7_75t_L g1180 ( 
.A(n_1132),
.Y(n_1180)
);

OAI221xp5_ASAP7_75t_L g1181 ( 
.A1(n_1093),
.A2(n_899),
.B1(n_848),
.B2(n_891),
.C(n_828),
.Y(n_1181)
);

INVx1_ASAP7_75t_L g1182 ( 
.A(n_1099),
.Y(n_1182)
);

INVx2_ASAP7_75t_SL g1183 ( 
.A(n_1092),
.Y(n_1183)
);

NAND2xp5_ASAP7_75t_L g1184 ( 
.A(n_1121),
.B(n_952),
.Y(n_1184)
);

BUFx3_ASAP7_75t_L g1185 ( 
.A(n_1097),
.Y(n_1185)
);

AO22x2_ASAP7_75t_L g1186 ( 
.A1(n_1103),
.A2(n_999),
.B1(n_769),
.B2(n_787),
.Y(n_1186)
);

AO22x2_ASAP7_75t_L g1187 ( 
.A1(n_1108),
.A2(n_799),
.B1(n_801),
.B2(n_779),
.Y(n_1187)
);

INVx1_ASAP7_75t_L g1188 ( 
.A(n_1106),
.Y(n_1188)
);

NAND2xp5_ASAP7_75t_L g1189 ( 
.A(n_1108),
.B(n_804),
.Y(n_1189)
);

NAND2xp5_ASAP7_75t_L g1190 ( 
.A(n_1108),
.B(n_808),
.Y(n_1190)
);

CKINVDCx20_ASAP7_75t_R g1191 ( 
.A(n_1106),
.Y(n_1191)
);

INVx1_ASAP7_75t_L g1192 ( 
.A(n_1106),
.Y(n_1192)
);

INVx1_ASAP7_75t_L g1193 ( 
.A(n_1107),
.Y(n_1193)
);

OAI22xp5_ASAP7_75t_L g1194 ( 
.A1(n_1111),
.A2(n_935),
.B1(n_959),
.B2(n_912),
.Y(n_1194)
);

AO22x2_ASAP7_75t_L g1195 ( 
.A1(n_1095),
.A2(n_812),
.B1(n_816),
.B2(n_809),
.Y(n_1195)
);

AO22x2_ASAP7_75t_L g1196 ( 
.A1(n_1095),
.A2(n_831),
.B1(n_845),
.B2(n_827),
.Y(n_1196)
);

INVx1_ASAP7_75t_L g1197 ( 
.A(n_1107),
.Y(n_1197)
);

AO22x2_ASAP7_75t_L g1198 ( 
.A1(n_1095),
.A2(n_855),
.B1(n_858),
.B2(n_852),
.Y(n_1198)
);

OAI22xp33_ASAP7_75t_L g1199 ( 
.A1(n_1111),
.A2(n_965),
.B1(n_940),
.B2(n_930),
.Y(n_1199)
);

CKINVDCx20_ASAP7_75t_R g1200 ( 
.A(n_1100),
.Y(n_1200)
);

OAI221xp5_ASAP7_75t_L g1201 ( 
.A1(n_1127),
.A2(n_1011),
.B1(n_889),
.B2(n_898),
.C(n_883),
.Y(n_1201)
);

INVx1_ASAP7_75t_L g1202 ( 
.A(n_1107),
.Y(n_1202)
);

INVx1_ASAP7_75t_L g1203 ( 
.A(n_1107),
.Y(n_1203)
);

NAND2xp5_ASAP7_75t_L g1204 ( 
.A(n_1096),
.B(n_877),
.Y(n_1204)
);

NAND2x1p5_ASAP7_75t_L g1205 ( 
.A(n_1133),
.B(n_1027),
.Y(n_1205)
);

INVx1_ASAP7_75t_L g1206 ( 
.A(n_1107),
.Y(n_1206)
);

INVx1_ASAP7_75t_L g1207 ( 
.A(n_1107),
.Y(n_1207)
);

CKINVDCx20_ASAP7_75t_R g1208 ( 
.A(n_1100),
.Y(n_1208)
);

NOR2xp33_ASAP7_75t_L g1209 ( 
.A(n_1125),
.B(n_746),
.Y(n_1209)
);

INVx1_ASAP7_75t_L g1210 ( 
.A(n_1107),
.Y(n_1210)
);

INVx1_ASAP7_75t_L g1211 ( 
.A(n_1107),
.Y(n_1211)
);

INVx1_ASAP7_75t_L g1212 ( 
.A(n_1107),
.Y(n_1212)
);

INVx1_ASAP7_75t_L g1213 ( 
.A(n_1107),
.Y(n_1213)
);

INVx1_ASAP7_75t_L g1214 ( 
.A(n_1107),
.Y(n_1214)
);

INVx1_ASAP7_75t_L g1215 ( 
.A(n_1107),
.Y(n_1215)
);

NAND2xp5_ASAP7_75t_L g1216 ( 
.A(n_1096),
.B(n_908),
.Y(n_1216)
);

AOI22xp33_ASAP7_75t_L g1217 ( 
.A1(n_1120),
.A2(n_785),
.B1(n_786),
.B2(n_772),
.Y(n_1217)
);

INVx1_ASAP7_75t_L g1218 ( 
.A(n_1107),
.Y(n_1218)
);

AO22x2_ASAP7_75t_L g1219 ( 
.A1(n_1095),
.A2(n_916),
.B1(n_927),
.B2(n_909),
.Y(n_1219)
);

INVx2_ASAP7_75t_L g1220 ( 
.A(n_1104),
.Y(n_1220)
);

AO22x2_ASAP7_75t_L g1221 ( 
.A1(n_1095),
.A2(n_938),
.B1(n_953),
.B2(n_936),
.Y(n_1221)
);

INVx1_ASAP7_75t_L g1222 ( 
.A(n_1107),
.Y(n_1222)
);

AND2x2_ASAP7_75t_L g1223 ( 
.A(n_1096),
.B(n_741),
.Y(n_1223)
);

INVxp67_ASAP7_75t_L g1224 ( 
.A(n_1128),
.Y(n_1224)
);

NOR2xp33_ASAP7_75t_L g1225 ( 
.A(n_1125),
.B(n_753),
.Y(n_1225)
);

AO22x2_ASAP7_75t_L g1226 ( 
.A1(n_1095),
.A2(n_980),
.B1(n_995),
.B2(n_961),
.Y(n_1226)
);

OR2x2_ASAP7_75t_SL g1227 ( 
.A(n_1125),
.B(n_901),
.Y(n_1227)
);

OA22x2_ASAP7_75t_L g1228 ( 
.A1(n_1095),
.A2(n_762),
.B1(n_763),
.B2(n_761),
.Y(n_1228)
);

NAND2x1p5_ASAP7_75t_L g1229 ( 
.A(n_1133),
.B(n_1004),
.Y(n_1229)
);

INVx1_ASAP7_75t_L g1230 ( 
.A(n_1107),
.Y(n_1230)
);

AND2x2_ASAP7_75t_L g1231 ( 
.A(n_1096),
.B(n_932),
.Y(n_1231)
);

INVx1_ASAP7_75t_L g1232 ( 
.A(n_1107),
.Y(n_1232)
);

NAND2xp5_ASAP7_75t_SL g1233 ( 
.A(n_1125),
.B(n_1018),
.Y(n_1233)
);

INVx1_ASAP7_75t_L g1234 ( 
.A(n_1107),
.Y(n_1234)
);

AO22x2_ASAP7_75t_L g1235 ( 
.A1(n_1095),
.A2(n_1009),
.B1(n_1012),
.B2(n_1007),
.Y(n_1235)
);

AO22x2_ASAP7_75t_L g1236 ( 
.A1(n_1095),
.A2(n_1017),
.B1(n_870),
.B2(n_805),
.Y(n_1236)
);

INVx2_ASAP7_75t_L g1237 ( 
.A(n_1104),
.Y(n_1237)
);

INVx2_ASAP7_75t_L g1238 ( 
.A(n_1104),
.Y(n_1238)
);

NAND2xp5_ASAP7_75t_SL g1239 ( 
.A(n_1143),
.B(n_776),
.Y(n_1239)
);

NAND2xp5_ASAP7_75t_SL g1240 ( 
.A(n_1224),
.B(n_781),
.Y(n_1240)
);

AND2x2_ASAP7_75t_L g1241 ( 
.A(n_1146),
.B(n_764),
.Y(n_1241)
);

NAND2xp5_ASAP7_75t_SL g1242 ( 
.A(n_1199),
.B(n_783),
.Y(n_1242)
);

NAND2xp5_ASAP7_75t_SL g1243 ( 
.A(n_1162),
.B(n_784),
.Y(n_1243)
);

NAND2xp5_ASAP7_75t_L g1244 ( 
.A(n_1138),
.B(n_857),
.Y(n_1244)
);

NAND2xp5_ASAP7_75t_SL g1245 ( 
.A(n_1171),
.B(n_1209),
.Y(n_1245)
);

NAND2xp5_ASAP7_75t_SL g1246 ( 
.A(n_1225),
.B(n_788),
.Y(n_1246)
);

NAND2xp5_ASAP7_75t_SL g1247 ( 
.A(n_1141),
.B(n_789),
.Y(n_1247)
);

AND2x4_ASAP7_75t_L g1248 ( 
.A(n_1185),
.B(n_958),
.Y(n_1248)
);

NAND2xp5_ASAP7_75t_L g1249 ( 
.A(n_1139),
.B(n_987),
.Y(n_1249)
);

NAND2xp33_ASAP7_75t_SL g1250 ( 
.A(n_1191),
.B(n_1142),
.Y(n_1250)
);

NAND2xp33_ASAP7_75t_SL g1251 ( 
.A(n_1177),
.B(n_983),
.Y(n_1251)
);

NAND2xp5_ASAP7_75t_L g1252 ( 
.A(n_1148),
.B(n_1149),
.Y(n_1252)
);

NAND2xp5_ASAP7_75t_SL g1253 ( 
.A(n_1193),
.B(n_793),
.Y(n_1253)
);

NAND2xp5_ASAP7_75t_SL g1254 ( 
.A(n_1197),
.B(n_803),
.Y(n_1254)
);

NAND2xp5_ASAP7_75t_SL g1255 ( 
.A(n_1202),
.B(n_806),
.Y(n_1255)
);

NAND2xp5_ASAP7_75t_SL g1256 ( 
.A(n_1203),
.B(n_1206),
.Y(n_1256)
);

NAND2xp5_ASAP7_75t_SL g1257 ( 
.A(n_1207),
.B(n_807),
.Y(n_1257)
);

NAND2xp5_ASAP7_75t_SL g1258 ( 
.A(n_1210),
.B(n_813),
.Y(n_1258)
);

NAND2xp5_ASAP7_75t_L g1259 ( 
.A(n_1211),
.B(n_1019),
.Y(n_1259)
);

NAND2xp5_ASAP7_75t_SL g1260 ( 
.A(n_1212),
.B(n_1213),
.Y(n_1260)
);

AND2x4_ASAP7_75t_L g1261 ( 
.A(n_1172),
.B(n_1023),
.Y(n_1261)
);

NAND2xp33_ASAP7_75t_SL g1262 ( 
.A(n_1200),
.B(n_985),
.Y(n_1262)
);

NAND2xp33_ASAP7_75t_SL g1263 ( 
.A(n_1208),
.B(n_815),
.Y(n_1263)
);

NAND2xp5_ASAP7_75t_SL g1264 ( 
.A(n_1214),
.B(n_819),
.Y(n_1264)
);

NAND2xp33_ASAP7_75t_SL g1265 ( 
.A(n_1147),
.B(n_820),
.Y(n_1265)
);

NAND2xp33_ASAP7_75t_SL g1266 ( 
.A(n_1156),
.B(n_821),
.Y(n_1266)
);

NAND2xp5_ASAP7_75t_SL g1267 ( 
.A(n_1215),
.B(n_826),
.Y(n_1267)
);

NAND2xp5_ASAP7_75t_SL g1268 ( 
.A(n_1218),
.B(n_832),
.Y(n_1268)
);

NAND2xp5_ASAP7_75t_SL g1269 ( 
.A(n_1222),
.B(n_834),
.Y(n_1269)
);

NAND2xp5_ASAP7_75t_SL g1270 ( 
.A(n_1230),
.B(n_1232),
.Y(n_1270)
);

NAND2xp5_ASAP7_75t_SL g1271 ( 
.A(n_1234),
.B(n_836),
.Y(n_1271)
);

NAND2xp5_ASAP7_75t_SL g1272 ( 
.A(n_1157),
.B(n_838),
.Y(n_1272)
);

NAND2xp5_ASAP7_75t_SL g1273 ( 
.A(n_1166),
.B(n_843),
.Y(n_1273)
);

NAND2xp33_ASAP7_75t_SL g1274 ( 
.A(n_1178),
.B(n_850),
.Y(n_1274)
);

NAND2xp33_ASAP7_75t_SL g1275 ( 
.A(n_1233),
.B(n_851),
.Y(n_1275)
);

NAND2xp5_ASAP7_75t_SL g1276 ( 
.A(n_1155),
.B(n_1194),
.Y(n_1276)
);

NAND2xp5_ASAP7_75t_SL g1277 ( 
.A(n_1150),
.B(n_854),
.Y(n_1277)
);

NAND2xp5_ASAP7_75t_L g1278 ( 
.A(n_1204),
.B(n_856),
.Y(n_1278)
);

NAND2xp33_ASAP7_75t_SL g1279 ( 
.A(n_1223),
.B(n_1231),
.Y(n_1279)
);

NAND2xp5_ASAP7_75t_SL g1280 ( 
.A(n_1164),
.B(n_860),
.Y(n_1280)
);

NAND2xp5_ASAP7_75t_SL g1281 ( 
.A(n_1165),
.B(n_861),
.Y(n_1281)
);

NAND2xp5_ASAP7_75t_SL g1282 ( 
.A(n_1216),
.B(n_863),
.Y(n_1282)
);

NAND2xp5_ASAP7_75t_SL g1283 ( 
.A(n_1161),
.B(n_1220),
.Y(n_1283)
);

NAND2xp5_ASAP7_75t_SL g1284 ( 
.A(n_1237),
.B(n_864),
.Y(n_1284)
);

NAND2xp5_ASAP7_75t_SL g1285 ( 
.A(n_1238),
.B(n_1163),
.Y(n_1285)
);

NAND2xp5_ASAP7_75t_SL g1286 ( 
.A(n_1144),
.B(n_869),
.Y(n_1286)
);

NAND2xp5_ASAP7_75t_SL g1287 ( 
.A(n_1154),
.B(n_872),
.Y(n_1287)
);

NAND2xp5_ASAP7_75t_L g1288 ( 
.A(n_1217),
.B(n_874),
.Y(n_1288)
);

NAND2xp33_ASAP7_75t_SL g1289 ( 
.A(n_1188),
.B(n_880),
.Y(n_1289)
);

NAND2xp5_ASAP7_75t_SL g1290 ( 
.A(n_1159),
.B(n_884),
.Y(n_1290)
);

NAND2xp5_ASAP7_75t_SL g1291 ( 
.A(n_1229),
.B(n_888),
.Y(n_1291)
);

NAND2xp5_ASAP7_75t_SL g1292 ( 
.A(n_1152),
.B(n_894),
.Y(n_1292)
);

NAND2xp5_ASAP7_75t_SL g1293 ( 
.A(n_1153),
.B(n_896),
.Y(n_1293)
);

NAND2xp5_ASAP7_75t_SL g1294 ( 
.A(n_1167),
.B(n_897),
.Y(n_1294)
);

NAND2xp5_ASAP7_75t_SL g1295 ( 
.A(n_1169),
.B(n_903),
.Y(n_1295)
);

NAND2xp33_ASAP7_75t_SL g1296 ( 
.A(n_1192),
.B(n_905),
.Y(n_1296)
);

NAND2xp33_ASAP7_75t_SL g1297 ( 
.A(n_1183),
.B(n_906),
.Y(n_1297)
);

NAND2xp5_ASAP7_75t_SL g1298 ( 
.A(n_1168),
.B(n_907),
.Y(n_1298)
);

AND2x2_ASAP7_75t_L g1299 ( 
.A(n_1186),
.B(n_773),
.Y(n_1299)
);

NAND2xp5_ASAP7_75t_SL g1300 ( 
.A(n_1205),
.B(n_913),
.Y(n_1300)
);

NAND2xp33_ASAP7_75t_SL g1301 ( 
.A(n_1176),
.B(n_914),
.Y(n_1301)
);

NAND2xp5_ASAP7_75t_SL g1302 ( 
.A(n_1179),
.B(n_917),
.Y(n_1302)
);

NAND2xp33_ASAP7_75t_SL g1303 ( 
.A(n_1189),
.B(n_920),
.Y(n_1303)
);

NAND2xp5_ASAP7_75t_L g1304 ( 
.A(n_1182),
.B(n_924),
.Y(n_1304)
);

NAND2xp5_ASAP7_75t_SL g1305 ( 
.A(n_1170),
.B(n_929),
.Y(n_1305)
);

NAND2xp5_ASAP7_75t_SL g1306 ( 
.A(n_1180),
.B(n_931),
.Y(n_1306)
);

AND2x2_ASAP7_75t_L g1307 ( 
.A(n_1160),
.B(n_775),
.Y(n_1307)
);

NAND2xp5_ASAP7_75t_SL g1308 ( 
.A(n_1228),
.B(n_934),
.Y(n_1308)
);

NAND2xp5_ASAP7_75t_SL g1309 ( 
.A(n_1190),
.B(n_939),
.Y(n_1309)
);

NOR2xp33_ASAP7_75t_L g1310 ( 
.A(n_1227),
.B(n_778),
.Y(n_1310)
);

NAND2xp5_ASAP7_75t_SL g1311 ( 
.A(n_1184),
.B(n_941),
.Y(n_1311)
);

NAND2xp33_ASAP7_75t_SL g1312 ( 
.A(n_1175),
.B(n_945),
.Y(n_1312)
);

NAND2xp5_ASAP7_75t_SL g1313 ( 
.A(n_1145),
.B(n_947),
.Y(n_1313)
);

NAND2xp5_ASAP7_75t_SL g1314 ( 
.A(n_1174),
.B(n_951),
.Y(n_1314)
);

NAND2xp5_ASAP7_75t_SL g1315 ( 
.A(n_1236),
.B(n_954),
.Y(n_1315)
);

NAND2xp5_ASAP7_75t_SL g1316 ( 
.A(n_1195),
.B(n_955),
.Y(n_1316)
);

NAND2xp5_ASAP7_75t_SL g1317 ( 
.A(n_1196),
.B(n_956),
.Y(n_1317)
);

NAND2xp5_ASAP7_75t_SL g1318 ( 
.A(n_1198),
.B(n_963),
.Y(n_1318)
);

NAND2xp5_ASAP7_75t_SL g1319 ( 
.A(n_1219),
.B(n_966),
.Y(n_1319)
);

NAND2xp5_ASAP7_75t_SL g1320 ( 
.A(n_1221),
.B(n_969),
.Y(n_1320)
);

NAND2xp5_ASAP7_75t_SL g1321 ( 
.A(n_1226),
.B(n_970),
.Y(n_1321)
);

NAND2xp5_ASAP7_75t_SL g1322 ( 
.A(n_1235),
.B(n_971),
.Y(n_1322)
);

NAND2xp33_ASAP7_75t_SL g1323 ( 
.A(n_1140),
.B(n_974),
.Y(n_1323)
);

NAND2xp5_ASAP7_75t_SL g1324 ( 
.A(n_1158),
.B(n_978),
.Y(n_1324)
);

NAND2xp33_ASAP7_75t_SL g1325 ( 
.A(n_1187),
.B(n_979),
.Y(n_1325)
);

NAND2xp5_ASAP7_75t_SL g1326 ( 
.A(n_1158),
.B(n_981),
.Y(n_1326)
);

NAND2xp5_ASAP7_75t_SL g1327 ( 
.A(n_1158),
.B(n_989),
.Y(n_1327)
);

NAND2xp33_ASAP7_75t_SL g1328 ( 
.A(n_1151),
.B(n_990),
.Y(n_1328)
);

NAND2xp5_ASAP7_75t_SL g1329 ( 
.A(n_1151),
.B(n_996),
.Y(n_1329)
);

NAND2xp5_ASAP7_75t_SL g1330 ( 
.A(n_1201),
.B(n_1008),
.Y(n_1330)
);

NAND2xp33_ASAP7_75t_SL g1331 ( 
.A(n_1181),
.B(n_1010),
.Y(n_1331)
);

NAND2xp5_ASAP7_75t_SL g1332 ( 
.A(n_1137),
.B(n_1013),
.Y(n_1332)
);

AND2x2_ASAP7_75t_L g1333 ( 
.A(n_1173),
.B(n_780),
.Y(n_1333)
);

NAND2xp5_ASAP7_75t_SL g1334 ( 
.A(n_1143),
.B(n_1021),
.Y(n_1334)
);

NAND2xp5_ASAP7_75t_SL g1335 ( 
.A(n_1143),
.B(n_1022),
.Y(n_1335)
);

AND2x4_ASAP7_75t_L g1336 ( 
.A(n_1162),
.B(n_350),
.Y(n_1336)
);

NAND2xp5_ASAP7_75t_SL g1337 ( 
.A(n_1143),
.B(n_1025),
.Y(n_1337)
);

NAND2xp5_ASAP7_75t_L g1338 ( 
.A(n_1143),
.B(n_1026),
.Y(n_1338)
);

NAND2xp5_ASAP7_75t_SL g1339 ( 
.A(n_1143),
.B(n_871),
.Y(n_1339)
);

NAND2xp5_ASAP7_75t_L g1340 ( 
.A(n_1143),
.B(n_840),
.Y(n_1340)
);

NAND2xp5_ASAP7_75t_SL g1341 ( 
.A(n_1143),
.B(n_871),
.Y(n_1341)
);

NAND2xp5_ASAP7_75t_SL g1342 ( 
.A(n_1143),
.B(n_923),
.Y(n_1342)
);

NAND2xp5_ASAP7_75t_SL g1343 ( 
.A(n_1143),
.B(n_923),
.Y(n_1343)
);

NAND2xp5_ASAP7_75t_SL g1344 ( 
.A(n_1143),
.B(n_937),
.Y(n_1344)
);

AND2x2_ASAP7_75t_L g1345 ( 
.A(n_1143),
.B(n_790),
.Y(n_1345)
);

NAND2xp5_ASAP7_75t_SL g1346 ( 
.A(n_1143),
.B(n_937),
.Y(n_1346)
);

NAND2xp5_ASAP7_75t_SL g1347 ( 
.A(n_1143),
.B(n_968),
.Y(n_1347)
);

NAND2xp5_ASAP7_75t_SL g1348 ( 
.A(n_1143),
.B(n_968),
.Y(n_1348)
);

NAND2xp5_ASAP7_75t_SL g1349 ( 
.A(n_1143),
.B(n_840),
.Y(n_1349)
);

NAND2xp5_ASAP7_75t_SL g1350 ( 
.A(n_1143),
.B(n_840),
.Y(n_1350)
);

NAND2xp5_ASAP7_75t_SL g1351 ( 
.A(n_1143),
.B(n_867),
.Y(n_1351)
);

NAND2xp5_ASAP7_75t_SL g1352 ( 
.A(n_1143),
.B(n_867),
.Y(n_1352)
);

NAND2xp33_ASAP7_75t_SL g1353 ( 
.A(n_1191),
.B(n_792),
.Y(n_1353)
);

NAND2xp5_ASAP7_75t_SL g1354 ( 
.A(n_1143),
.B(n_867),
.Y(n_1354)
);

NAND2xp5_ASAP7_75t_L g1355 ( 
.A(n_1143),
.B(n_892),
.Y(n_1355)
);

NAND2xp5_ASAP7_75t_SL g1356 ( 
.A(n_1143),
.B(n_892),
.Y(n_1356)
);

NAND2xp5_ASAP7_75t_SL g1357 ( 
.A(n_1143),
.B(n_892),
.Y(n_1357)
);

AND2x4_ASAP7_75t_L g1358 ( 
.A(n_1162),
.B(n_352),
.Y(n_1358)
);

NAND2xp5_ASAP7_75t_SL g1359 ( 
.A(n_1143),
.B(n_964),
.Y(n_1359)
);

NAND2xp5_ASAP7_75t_L g1360 ( 
.A(n_1143),
.B(n_911),
.Y(n_1360)
);

NAND2xp5_ASAP7_75t_SL g1361 ( 
.A(n_1143),
.B(n_964),
.Y(n_1361)
);

NAND2xp33_ASAP7_75t_SL g1362 ( 
.A(n_1191),
.B(n_796),
.Y(n_1362)
);

NAND2xp33_ASAP7_75t_SL g1363 ( 
.A(n_1191),
.B(n_798),
.Y(n_1363)
);

AND2x2_ASAP7_75t_L g1364 ( 
.A(n_1143),
.B(n_800),
.Y(n_1364)
);

NAND2xp5_ASAP7_75t_SL g1365 ( 
.A(n_1143),
.B(n_911),
.Y(n_1365)
);

NAND2xp5_ASAP7_75t_SL g1366 ( 
.A(n_1143),
.B(n_911),
.Y(n_1366)
);

NAND2xp33_ASAP7_75t_SL g1367 ( 
.A(n_1191),
.B(n_811),
.Y(n_1367)
);

NAND2xp5_ASAP7_75t_SL g1368 ( 
.A(n_1143),
.B(n_964),
.Y(n_1368)
);

NAND2xp5_ASAP7_75t_SL g1369 ( 
.A(n_1143),
.B(n_818),
.Y(n_1369)
);

AND2x2_ASAP7_75t_L g1370 ( 
.A(n_1143),
.B(n_824),
.Y(n_1370)
);

NAND2xp33_ASAP7_75t_SL g1371 ( 
.A(n_1191),
.B(n_829),
.Y(n_1371)
);

NAND2xp5_ASAP7_75t_SL g1372 ( 
.A(n_1143),
.B(n_835),
.Y(n_1372)
);

NAND2xp5_ASAP7_75t_SL g1373 ( 
.A(n_1143),
.B(n_841),
.Y(n_1373)
);

NAND2xp5_ASAP7_75t_SL g1374 ( 
.A(n_1143),
.B(n_842),
.Y(n_1374)
);

NAND2xp5_ASAP7_75t_SL g1375 ( 
.A(n_1143),
.B(n_844),
.Y(n_1375)
);

NAND2xp5_ASAP7_75t_L g1376 ( 
.A(n_1143),
.B(n_846),
.Y(n_1376)
);

NAND2xp5_ASAP7_75t_SL g1377 ( 
.A(n_1143),
.B(n_849),
.Y(n_1377)
);

NAND2xp5_ASAP7_75t_SL g1378 ( 
.A(n_1143),
.B(n_859),
.Y(n_1378)
);

AND2x4_ASAP7_75t_L g1379 ( 
.A(n_1162),
.B(n_353),
.Y(n_1379)
);

NAND2xp5_ASAP7_75t_SL g1380 ( 
.A(n_1143),
.B(n_865),
.Y(n_1380)
);

NAND2xp5_ASAP7_75t_SL g1381 ( 
.A(n_1143),
.B(n_868),
.Y(n_1381)
);

NAND2xp5_ASAP7_75t_L g1382 ( 
.A(n_1143),
.B(n_875),
.Y(n_1382)
);

NAND2xp5_ASAP7_75t_SL g1383 ( 
.A(n_1143),
.B(n_876),
.Y(n_1383)
);

AND2x2_ASAP7_75t_SL g1384 ( 
.A(n_1146),
.B(n_0),
.Y(n_1384)
);

NAND2xp5_ASAP7_75t_SL g1385 ( 
.A(n_1143),
.B(n_886),
.Y(n_1385)
);

NAND2xp33_ASAP7_75t_SL g1386 ( 
.A(n_1191),
.B(n_895),
.Y(n_1386)
);

NAND2xp5_ASAP7_75t_SL g1387 ( 
.A(n_1143),
.B(n_904),
.Y(n_1387)
);

NAND2xp5_ASAP7_75t_SL g1388 ( 
.A(n_1143),
.B(n_921),
.Y(n_1388)
);

NAND2xp5_ASAP7_75t_SL g1389 ( 
.A(n_1143),
.B(n_928),
.Y(n_1389)
);

AND2x2_ASAP7_75t_L g1390 ( 
.A(n_1143),
.B(n_943),
.Y(n_1390)
);

NAND2xp33_ASAP7_75t_SL g1391 ( 
.A(n_1191),
.B(n_944),
.Y(n_1391)
);

NAND2xp5_ASAP7_75t_L g1392 ( 
.A(n_1143),
.B(n_948),
.Y(n_1392)
);

NAND2xp5_ASAP7_75t_SL g1393 ( 
.A(n_1143),
.B(n_950),
.Y(n_1393)
);

NAND2xp5_ASAP7_75t_SL g1394 ( 
.A(n_1143),
.B(n_967),
.Y(n_1394)
);

A2O1A1Ixp33_ASAP7_75t_L g1395 ( 
.A1(n_1245),
.A2(n_984),
.B(n_986),
.C(n_975),
.Y(n_1395)
);

NOR2xp33_ASAP7_75t_L g1396 ( 
.A(n_1338),
.B(n_988),
.Y(n_1396)
);

AND2x6_ASAP7_75t_L g1397 ( 
.A(n_1336),
.B(n_354),
.Y(n_1397)
);

NAND2xp5_ASAP7_75t_L g1398 ( 
.A(n_1252),
.B(n_992),
.Y(n_1398)
);

AOI21xp5_ASAP7_75t_L g1399 ( 
.A1(n_1256),
.A2(n_357),
.B(n_356),
.Y(n_1399)
);

NAND2xp5_ASAP7_75t_L g1400 ( 
.A(n_1345),
.B(n_1364),
.Y(n_1400)
);

BUFx2_ASAP7_75t_L g1401 ( 
.A(n_1251),
.Y(n_1401)
);

AOI21xp5_ASAP7_75t_L g1402 ( 
.A1(n_1260),
.A2(n_359),
.B(n_358),
.Y(n_1402)
);

NAND2xp5_ASAP7_75t_L g1403 ( 
.A(n_1370),
.B(n_1390),
.Y(n_1403)
);

NAND3xp33_ASAP7_75t_L g1404 ( 
.A(n_1276),
.B(n_994),
.C(n_993),
.Y(n_1404)
);

CKINVDCx14_ASAP7_75t_R g1405 ( 
.A(n_1262),
.Y(n_1405)
);

AOI221x1_ASAP7_75t_L g1406 ( 
.A1(n_1312),
.A2(n_5),
.B1(n_3),
.B2(n_4),
.C(n_6),
.Y(n_1406)
);

NOR2xp33_ASAP7_75t_L g1407 ( 
.A(n_1376),
.B(n_1000),
.Y(n_1407)
);

AO31x2_ASAP7_75t_L g1408 ( 
.A1(n_1244),
.A2(n_362),
.A3(n_364),
.B(n_361),
.Y(n_1408)
);

NAND2xp5_ASAP7_75t_L g1409 ( 
.A(n_1340),
.B(n_1355),
.Y(n_1409)
);

AOI21xp5_ASAP7_75t_L g1410 ( 
.A1(n_1270),
.A2(n_366),
.B(n_365),
.Y(n_1410)
);

CKINVDCx5p33_ASAP7_75t_R g1411 ( 
.A(n_1250),
.Y(n_1411)
);

INVx3_ASAP7_75t_L g1412 ( 
.A(n_1248),
.Y(n_1412)
);

INVx2_ASAP7_75t_L g1413 ( 
.A(n_1283),
.Y(n_1413)
);

NAND2x1p5_ASAP7_75t_L g1414 ( 
.A(n_1336),
.B(n_369),
.Y(n_1414)
);

NAND2xp5_ASAP7_75t_L g1415 ( 
.A(n_1360),
.B(n_1002),
.Y(n_1415)
);

OR2x6_ASAP7_75t_L g1416 ( 
.A(n_1358),
.B(n_5),
.Y(n_1416)
);

NAND2xp5_ASAP7_75t_L g1417 ( 
.A(n_1382),
.B(n_1005),
.Y(n_1417)
);

OAI21x1_ASAP7_75t_L g1418 ( 
.A1(n_1249),
.A2(n_374),
.B(n_372),
.Y(n_1418)
);

AOI22xp33_ASAP7_75t_L g1419 ( 
.A1(n_1242),
.A2(n_1323),
.B1(n_1279),
.B2(n_1261),
.Y(n_1419)
);

OR2x2_ASAP7_75t_L g1420 ( 
.A(n_1392),
.B(n_1014),
.Y(n_1420)
);

AND2x4_ASAP7_75t_L g1421 ( 
.A(n_1248),
.B(n_375),
.Y(n_1421)
);

AOI21xp5_ASAP7_75t_L g1422 ( 
.A1(n_1311),
.A2(n_377),
.B(n_376),
.Y(n_1422)
);

AND3x2_ASAP7_75t_L g1423 ( 
.A(n_1310),
.B(n_6),
.C(n_7),
.Y(n_1423)
);

NAND2xp5_ASAP7_75t_SL g1424 ( 
.A(n_1358),
.B(n_1015),
.Y(n_1424)
);

AO31x2_ASAP7_75t_L g1425 ( 
.A1(n_1259),
.A2(n_1304),
.A3(n_1278),
.B(n_1288),
.Y(n_1425)
);

OAI21x1_ASAP7_75t_L g1426 ( 
.A1(n_1285),
.A2(n_380),
.B(n_378),
.Y(n_1426)
);

AND2x2_ASAP7_75t_L g1427 ( 
.A(n_1241),
.B(n_1020),
.Y(n_1427)
);

AOI21xp5_ASAP7_75t_L g1428 ( 
.A1(n_1280),
.A2(n_390),
.B(n_386),
.Y(n_1428)
);

INVx2_ASAP7_75t_L g1429 ( 
.A(n_1261),
.Y(n_1429)
);

BUFx3_ASAP7_75t_L g1430 ( 
.A(n_1379),
.Y(n_1430)
);

NOR2xp33_ASAP7_75t_L g1431 ( 
.A(n_1369),
.B(n_1029),
.Y(n_1431)
);

OA21x2_ASAP7_75t_L g1432 ( 
.A1(n_1306),
.A2(n_1302),
.B(n_1284),
.Y(n_1432)
);

AND2x4_ASAP7_75t_L g1433 ( 
.A(n_1379),
.B(n_1329),
.Y(n_1433)
);

BUFx2_ASAP7_75t_L g1434 ( 
.A(n_1353),
.Y(n_1434)
);

OA21x2_ASAP7_75t_L g1435 ( 
.A1(n_1292),
.A2(n_393),
.B(n_391),
.Y(n_1435)
);

OAI21xp5_ASAP7_75t_L g1436 ( 
.A1(n_1282),
.A2(n_397),
.B(n_396),
.Y(n_1436)
);

OAI21x1_ASAP7_75t_L g1437 ( 
.A1(n_1324),
.A2(n_400),
.B(n_399),
.Y(n_1437)
);

INVx2_ASAP7_75t_L g1438 ( 
.A(n_1273),
.Y(n_1438)
);

OAI21x1_ASAP7_75t_L g1439 ( 
.A1(n_1326),
.A2(n_402),
.B(n_401),
.Y(n_1439)
);

OAI21x1_ASAP7_75t_L g1440 ( 
.A1(n_1327),
.A2(n_1293),
.B(n_1309),
.Y(n_1440)
);

NAND2xp5_ASAP7_75t_L g1441 ( 
.A(n_1246),
.B(n_8),
.Y(n_1441)
);

AOI21xp5_ASAP7_75t_L g1442 ( 
.A1(n_1281),
.A2(n_404),
.B(n_403),
.Y(n_1442)
);

AND2x4_ASAP7_75t_L g1443 ( 
.A(n_1298),
.B(n_405),
.Y(n_1443)
);

INVx1_ASAP7_75t_L g1444 ( 
.A(n_1349),
.Y(n_1444)
);

O2A1O1Ixp5_ASAP7_75t_SL g1445 ( 
.A1(n_1316),
.A2(n_11),
.B(n_9),
.C(n_10),
.Y(n_1445)
);

INVx1_ASAP7_75t_SL g1446 ( 
.A(n_1384),
.Y(n_1446)
);

OR2x6_ASAP7_75t_L g1447 ( 
.A(n_1300),
.B(n_9),
.Y(n_1447)
);

OAI21x1_ASAP7_75t_L g1448 ( 
.A1(n_1287),
.A2(n_407),
.B(n_406),
.Y(n_1448)
);

NAND3x1_ASAP7_75t_L g1449 ( 
.A(n_1307),
.B(n_10),
.C(n_11),
.Y(n_1449)
);

INVx1_ASAP7_75t_SL g1450 ( 
.A(n_1263),
.Y(n_1450)
);

AOI21xp5_ASAP7_75t_L g1451 ( 
.A1(n_1253),
.A2(n_410),
.B(n_409),
.Y(n_1451)
);

AND2x2_ASAP7_75t_L g1452 ( 
.A(n_1333),
.B(n_12),
.Y(n_1452)
);

A2O1A1Ixp33_ASAP7_75t_L g1453 ( 
.A1(n_1265),
.A2(n_14),
.B(n_12),
.C(n_13),
.Y(n_1453)
);

OAI22xp5_ASAP7_75t_L g1454 ( 
.A1(n_1239),
.A2(n_413),
.B1(n_414),
.B2(n_412),
.Y(n_1454)
);

AOI21xp5_ASAP7_75t_L g1455 ( 
.A1(n_1254),
.A2(n_1257),
.B(n_1255),
.Y(n_1455)
);

NOR4xp25_ASAP7_75t_L g1456 ( 
.A(n_1317),
.B(n_15),
.C(n_13),
.D(n_14),
.Y(n_1456)
);

OAI21x1_ASAP7_75t_L g1457 ( 
.A1(n_1290),
.A2(n_1295),
.B(n_1294),
.Y(n_1457)
);

OAI21x1_ASAP7_75t_L g1458 ( 
.A1(n_1286),
.A2(n_416),
.B(n_415),
.Y(n_1458)
);

INVx1_ASAP7_75t_L g1459 ( 
.A(n_1350),
.Y(n_1459)
);

AOI21x1_ASAP7_75t_L g1460 ( 
.A1(n_1258),
.A2(n_419),
.B(n_418),
.Y(n_1460)
);

NAND2xp5_ASAP7_75t_SL g1461 ( 
.A(n_1266),
.B(n_420),
.Y(n_1461)
);

AOI21xp5_ASAP7_75t_L g1462 ( 
.A1(n_1264),
.A2(n_422),
.B(n_421),
.Y(n_1462)
);

CKINVDCx14_ASAP7_75t_R g1463 ( 
.A(n_1362),
.Y(n_1463)
);

NAND2x1p5_ASAP7_75t_L g1464 ( 
.A(n_1305),
.B(n_424),
.Y(n_1464)
);

OAI21x1_ASAP7_75t_L g1465 ( 
.A1(n_1267),
.A2(n_427),
.B(n_426),
.Y(n_1465)
);

OAI21x1_ASAP7_75t_SL g1466 ( 
.A1(n_1289),
.A2(n_430),
.B(n_429),
.Y(n_1466)
);

CKINVDCx5p33_ASAP7_75t_R g1467 ( 
.A(n_1363),
.Y(n_1467)
);

OAI21xp5_ASAP7_75t_SL g1468 ( 
.A1(n_1299),
.A2(n_17),
.B(n_18),
.Y(n_1468)
);

OAI21x1_ASAP7_75t_L g1469 ( 
.A1(n_1268),
.A2(n_1271),
.B(n_1269),
.Y(n_1469)
);

CKINVDCx20_ASAP7_75t_R g1470 ( 
.A(n_1367),
.Y(n_1470)
);

NAND2xp5_ASAP7_75t_L g1471 ( 
.A(n_1240),
.B(n_19),
.Y(n_1471)
);

OAI21xp5_ASAP7_75t_L g1472 ( 
.A1(n_1277),
.A2(n_432),
.B(n_431),
.Y(n_1472)
);

OAI22xp5_ASAP7_75t_L g1473 ( 
.A1(n_1334),
.A2(n_434),
.B1(n_435),
.B2(n_433),
.Y(n_1473)
);

NAND2xp5_ASAP7_75t_L g1474 ( 
.A(n_1335),
.B(n_19),
.Y(n_1474)
);

AND2x2_ASAP7_75t_L g1475 ( 
.A(n_1394),
.B(n_1372),
.Y(n_1475)
);

NAND2xp5_ASAP7_75t_L g1476 ( 
.A(n_1337),
.B(n_20),
.Y(n_1476)
);

AND2x2_ASAP7_75t_L g1477 ( 
.A(n_1373),
.B(n_20),
.Y(n_1477)
);

INVx1_ASAP7_75t_L g1478 ( 
.A(n_1351),
.Y(n_1478)
);

NAND2xp5_ASAP7_75t_SL g1479 ( 
.A(n_1318),
.B(n_436),
.Y(n_1479)
);

NAND2xp5_ASAP7_75t_L g1480 ( 
.A(n_1374),
.B(n_21),
.Y(n_1480)
);

O2A1O1Ixp5_ASAP7_75t_SL g1481 ( 
.A1(n_1319),
.A2(n_24),
.B(n_22),
.C(n_23),
.Y(n_1481)
);

NAND2xp5_ASAP7_75t_L g1482 ( 
.A(n_1375),
.B(n_22),
.Y(n_1482)
);

INVx1_ASAP7_75t_L g1483 ( 
.A(n_1352),
.Y(n_1483)
);

NAND2xp5_ASAP7_75t_L g1484 ( 
.A(n_1377),
.B(n_1387),
.Y(n_1484)
);

INVx1_ASAP7_75t_L g1485 ( 
.A(n_1354),
.Y(n_1485)
);

NOR2xp33_ASAP7_75t_L g1486 ( 
.A(n_1378),
.B(n_23),
.Y(n_1486)
);

OA21x2_ASAP7_75t_L g1487 ( 
.A1(n_1356),
.A2(n_438),
.B(n_437),
.Y(n_1487)
);

NOR2xp67_ASAP7_75t_L g1488 ( 
.A(n_1339),
.B(n_441),
.Y(n_1488)
);

AOI21xp5_ASAP7_75t_SL g1489 ( 
.A1(n_1291),
.A2(n_444),
.B(n_443),
.Y(n_1489)
);

OAI21x1_ASAP7_75t_L g1490 ( 
.A1(n_1315),
.A2(n_446),
.B(n_445),
.Y(n_1490)
);

AOI21xp5_ASAP7_75t_L g1491 ( 
.A1(n_1243),
.A2(n_449),
.B(n_448),
.Y(n_1491)
);

AOI221xp5_ASAP7_75t_L g1492 ( 
.A1(n_1371),
.A2(n_26),
.B1(n_24),
.B2(n_25),
.C(n_27),
.Y(n_1492)
);

AO21x2_ASAP7_75t_L g1493 ( 
.A1(n_1247),
.A2(n_451),
.B(n_450),
.Y(n_1493)
);

HB1xp67_ASAP7_75t_L g1494 ( 
.A(n_1308),
.Y(n_1494)
);

INVx1_ASAP7_75t_L g1495 ( 
.A(n_1357),
.Y(n_1495)
);

OAI21x1_ASAP7_75t_L g1496 ( 
.A1(n_1359),
.A2(n_456),
.B(n_453),
.Y(n_1496)
);

AOI21xp5_ASAP7_75t_L g1497 ( 
.A1(n_1330),
.A2(n_458),
.B(n_457),
.Y(n_1497)
);

AND2x6_ASAP7_75t_L g1498 ( 
.A(n_1320),
.B(n_461),
.Y(n_1498)
);

INVx2_ASAP7_75t_L g1499 ( 
.A(n_1361),
.Y(n_1499)
);

AOI21xp5_ASAP7_75t_L g1500 ( 
.A1(n_1303),
.A2(n_464),
.B(n_462),
.Y(n_1500)
);

A2O1A1Ixp33_ASAP7_75t_L g1501 ( 
.A1(n_1331),
.A2(n_1275),
.B(n_1322),
.C(n_1321),
.Y(n_1501)
);

NAND2xp5_ASAP7_75t_L g1502 ( 
.A(n_1380),
.B(n_25),
.Y(n_1502)
);

AOI21xp33_ASAP7_75t_L g1503 ( 
.A1(n_1381),
.A2(n_26),
.B(n_28),
.Y(n_1503)
);

OAI21x1_ASAP7_75t_L g1504 ( 
.A1(n_1365),
.A2(n_468),
.B(n_465),
.Y(n_1504)
);

AND2x2_ASAP7_75t_SL g1505 ( 
.A(n_1325),
.B(n_28),
.Y(n_1505)
);

NAND2xp5_ASAP7_75t_L g1506 ( 
.A(n_1383),
.B(n_29),
.Y(n_1506)
);

INVx5_ASAP7_75t_L g1507 ( 
.A(n_1274),
.Y(n_1507)
);

OAI21x1_ASAP7_75t_L g1508 ( 
.A1(n_1366),
.A2(n_470),
.B(n_469),
.Y(n_1508)
);

NAND2xp5_ASAP7_75t_L g1509 ( 
.A(n_1385),
.B(n_29),
.Y(n_1509)
);

NOR2xp33_ASAP7_75t_SL g1510 ( 
.A(n_1386),
.B(n_1391),
.Y(n_1510)
);

AOI221xp5_ASAP7_75t_L g1511 ( 
.A1(n_1341),
.A2(n_32),
.B1(n_30),
.B2(n_31),
.C(n_33),
.Y(n_1511)
);

NAND2xp5_ASAP7_75t_L g1512 ( 
.A(n_1388),
.B(n_30),
.Y(n_1512)
);

OAI21x1_ASAP7_75t_L g1513 ( 
.A1(n_1368),
.A2(n_472),
.B(n_471),
.Y(n_1513)
);

OAI21x1_ASAP7_75t_L g1514 ( 
.A1(n_1314),
.A2(n_476),
.B(n_473),
.Y(n_1514)
);

AO21x1_ASAP7_75t_L g1515 ( 
.A1(n_1409),
.A2(n_1272),
.B(n_1296),
.Y(n_1515)
);

OA21x2_ASAP7_75t_L g1516 ( 
.A1(n_1440),
.A2(n_1332),
.B(n_1389),
.Y(n_1516)
);

OAI21x1_ASAP7_75t_L g1517 ( 
.A1(n_1426),
.A2(n_1343),
.B(n_1342),
.Y(n_1517)
);

OAI21x1_ASAP7_75t_L g1518 ( 
.A1(n_1437),
.A2(n_1346),
.B(n_1344),
.Y(n_1518)
);

OAI21x1_ASAP7_75t_L g1519 ( 
.A1(n_1439),
.A2(n_1348),
.B(n_1347),
.Y(n_1519)
);

OAI221xp5_ASAP7_75t_L g1520 ( 
.A1(n_1400),
.A2(n_1393),
.B1(n_1328),
.B2(n_1313),
.C(n_1297),
.Y(n_1520)
);

INVx3_ASAP7_75t_L g1521 ( 
.A(n_1412),
.Y(n_1521)
);

AOI22xp5_ASAP7_75t_L g1522 ( 
.A1(n_1403),
.A2(n_1301),
.B1(n_34),
.B2(n_32),
.Y(n_1522)
);

INVx2_ASAP7_75t_SL g1523 ( 
.A(n_1430),
.Y(n_1523)
);

OAI21x1_ASAP7_75t_L g1524 ( 
.A1(n_1490),
.A2(n_478),
.B(n_477),
.Y(n_1524)
);

OAI221xp5_ASAP7_75t_L g1525 ( 
.A1(n_1431),
.A2(n_35),
.B1(n_33),
.B2(n_34),
.C(n_36),
.Y(n_1525)
);

A2O1A1Ixp33_ASAP7_75t_L g1526 ( 
.A1(n_1396),
.A2(n_38),
.B(n_35),
.C(n_37),
.Y(n_1526)
);

OAI21x1_ASAP7_75t_L g1527 ( 
.A1(n_1418),
.A2(n_1465),
.B(n_1458),
.Y(n_1527)
);

INVx1_ASAP7_75t_L g1528 ( 
.A(n_1413),
.Y(n_1528)
);

AOI21xp5_ASAP7_75t_L g1529 ( 
.A1(n_1455),
.A2(n_481),
.B(n_480),
.Y(n_1529)
);

AOI22x1_ASAP7_75t_L g1530 ( 
.A1(n_1499),
.A2(n_483),
.B1(n_484),
.B2(n_482),
.Y(n_1530)
);

OAI21x1_ASAP7_75t_L g1531 ( 
.A1(n_1448),
.A2(n_486),
.B(n_485),
.Y(n_1531)
);

OAI21x1_ASAP7_75t_L g1532 ( 
.A1(n_1514),
.A2(n_489),
.B(n_488),
.Y(n_1532)
);

AO31x2_ASAP7_75t_L g1533 ( 
.A1(n_1501),
.A2(n_491),
.A3(n_492),
.B(n_490),
.Y(n_1533)
);

NAND2xp5_ASAP7_75t_L g1534 ( 
.A(n_1407),
.B(n_37),
.Y(n_1534)
);

INVx1_ASAP7_75t_L g1535 ( 
.A(n_1429),
.Y(n_1535)
);

OAI21x1_ASAP7_75t_L g1536 ( 
.A1(n_1460),
.A2(n_494),
.B(n_493),
.Y(n_1536)
);

AND2x2_ASAP7_75t_L g1537 ( 
.A(n_1427),
.B(n_38),
.Y(n_1537)
);

INVx2_ASAP7_75t_L g1538 ( 
.A(n_1438),
.Y(n_1538)
);

INVx1_ASAP7_75t_L g1539 ( 
.A(n_1494),
.Y(n_1539)
);

INVx2_ASAP7_75t_L g1540 ( 
.A(n_1444),
.Y(n_1540)
);

INVx1_ASAP7_75t_L g1541 ( 
.A(n_1459),
.Y(n_1541)
);

NAND2x1_ASAP7_75t_L g1542 ( 
.A(n_1397),
.B(n_495),
.Y(n_1542)
);

AO31x2_ASAP7_75t_L g1543 ( 
.A1(n_1406),
.A2(n_497),
.A3(n_498),
.B(n_496),
.Y(n_1543)
);

A2O1A1Ixp33_ASAP7_75t_L g1544 ( 
.A1(n_1404),
.A2(n_41),
.B(n_39),
.C(n_40),
.Y(n_1544)
);

BUFx2_ASAP7_75t_L g1545 ( 
.A(n_1416),
.Y(n_1545)
);

INVx1_ASAP7_75t_L g1546 ( 
.A(n_1478),
.Y(n_1546)
);

OAI22xp5_ASAP7_75t_L g1547 ( 
.A1(n_1419),
.A2(n_1484),
.B1(n_1433),
.B2(n_1417),
.Y(n_1547)
);

CKINVDCx5p33_ASAP7_75t_R g1548 ( 
.A(n_1411),
.Y(n_1548)
);

INVx3_ASAP7_75t_L g1549 ( 
.A(n_1421),
.Y(n_1549)
);

A2O1A1Ixp33_ASAP7_75t_L g1550 ( 
.A1(n_1486),
.A2(n_42),
.B(n_39),
.C(n_40),
.Y(n_1550)
);

AO31x2_ASAP7_75t_L g1551 ( 
.A1(n_1453),
.A2(n_500),
.A3(n_501),
.B(n_499),
.Y(n_1551)
);

NAND2x1p5_ASAP7_75t_L g1552 ( 
.A(n_1507),
.B(n_511),
.Y(n_1552)
);

OAI21x1_ASAP7_75t_L g1553 ( 
.A1(n_1496),
.A2(n_503),
.B(n_502),
.Y(n_1553)
);

NAND2xp5_ASAP7_75t_L g1554 ( 
.A(n_1398),
.B(n_43),
.Y(n_1554)
);

INVx2_ASAP7_75t_L g1555 ( 
.A(n_1483),
.Y(n_1555)
);

NAND2x1p5_ASAP7_75t_L g1556 ( 
.A(n_1507),
.B(n_514),
.Y(n_1556)
);

HB1xp67_ASAP7_75t_L g1557 ( 
.A(n_1416),
.Y(n_1557)
);

OAI21x1_ASAP7_75t_L g1558 ( 
.A1(n_1504),
.A2(n_507),
.B(n_504),
.Y(n_1558)
);

INVx1_ASAP7_75t_L g1559 ( 
.A(n_1485),
.Y(n_1559)
);

OAI21x1_ASAP7_75t_L g1560 ( 
.A1(n_1508),
.A2(n_509),
.B(n_508),
.Y(n_1560)
);

OAI21xp5_ASAP7_75t_L g1561 ( 
.A1(n_1445),
.A2(n_512),
.B(n_510),
.Y(n_1561)
);

INVx1_ASAP7_75t_L g1562 ( 
.A(n_1495),
.Y(n_1562)
);

OAI22xp5_ASAP7_75t_L g1563 ( 
.A1(n_1415),
.A2(n_45),
.B1(n_43),
.B2(n_44),
.Y(n_1563)
);

NAND2xp5_ASAP7_75t_L g1564 ( 
.A(n_1452),
.B(n_1475),
.Y(n_1564)
);

INVx1_ASAP7_75t_L g1565 ( 
.A(n_1480),
.Y(n_1565)
);

AOI22xp33_ASAP7_75t_L g1566 ( 
.A1(n_1505),
.A2(n_46),
.B1(n_44),
.B2(n_45),
.Y(n_1566)
);

OA21x2_ASAP7_75t_L g1567 ( 
.A1(n_1469),
.A2(n_515),
.B(n_513),
.Y(n_1567)
);

OR2x2_ASAP7_75t_L g1568 ( 
.A(n_1446),
.B(n_1420),
.Y(n_1568)
);

OA21x2_ASAP7_75t_L g1569 ( 
.A1(n_1457),
.A2(n_519),
.B(n_518),
.Y(n_1569)
);

INVx2_ASAP7_75t_L g1570 ( 
.A(n_1425),
.Y(n_1570)
);

NAND2x1p5_ASAP7_75t_L g1571 ( 
.A(n_1450),
.B(n_522),
.Y(n_1571)
);

BUFx6f_ASAP7_75t_L g1572 ( 
.A(n_1434),
.Y(n_1572)
);

NAND2x1p5_ASAP7_75t_L g1573 ( 
.A(n_1461),
.B(n_524),
.Y(n_1573)
);

AOI22xp33_ASAP7_75t_L g1574 ( 
.A1(n_1401),
.A2(n_48),
.B1(n_46),
.B2(n_47),
.Y(n_1574)
);

CKINVDCx9p33_ASAP7_75t_R g1575 ( 
.A(n_1471),
.Y(n_1575)
);

CKINVDCx5p33_ASAP7_75t_R g1576 ( 
.A(n_1467),
.Y(n_1576)
);

OAI22xp33_ASAP7_75t_L g1577 ( 
.A1(n_1468),
.A2(n_50),
.B1(n_48),
.B2(n_49),
.Y(n_1577)
);

BUFx12f_ASAP7_75t_L g1578 ( 
.A(n_1447),
.Y(n_1578)
);

BUFx6f_ASAP7_75t_L g1579 ( 
.A(n_1443),
.Y(n_1579)
);

INVx2_ASAP7_75t_L g1580 ( 
.A(n_1425),
.Y(n_1580)
);

HB1xp67_ASAP7_75t_L g1581 ( 
.A(n_1414),
.Y(n_1581)
);

OAI21x1_ASAP7_75t_L g1582 ( 
.A1(n_1513),
.A2(n_521),
.B(n_520),
.Y(n_1582)
);

BUFx6f_ASAP7_75t_L g1583 ( 
.A(n_1447),
.Y(n_1583)
);

CKINVDCx6p67_ASAP7_75t_R g1584 ( 
.A(n_1470),
.Y(n_1584)
);

CKINVDCx8_ASAP7_75t_R g1585 ( 
.A(n_1498),
.Y(n_1585)
);

INVx1_ASAP7_75t_L g1586 ( 
.A(n_1482),
.Y(n_1586)
);

AO31x2_ASAP7_75t_L g1587 ( 
.A1(n_1497),
.A2(n_526),
.A3(n_527),
.B(n_525),
.Y(n_1587)
);

OAI22xp5_ASAP7_75t_L g1588 ( 
.A1(n_1424),
.A2(n_51),
.B1(n_49),
.B2(n_50),
.Y(n_1588)
);

NAND2xp5_ASAP7_75t_L g1589 ( 
.A(n_1477),
.B(n_51),
.Y(n_1589)
);

NAND2xp5_ASAP7_75t_L g1590 ( 
.A(n_1474),
.B(n_52),
.Y(n_1590)
);

OAI21x1_ASAP7_75t_SL g1591 ( 
.A1(n_1466),
.A2(n_533),
.B(n_532),
.Y(n_1591)
);

NAND2xp5_ASAP7_75t_L g1592 ( 
.A(n_1476),
.B(n_52),
.Y(n_1592)
);

NOR2xp33_ASAP7_75t_L g1593 ( 
.A(n_1405),
.B(n_53),
.Y(n_1593)
);

INVx1_ASAP7_75t_L g1594 ( 
.A(n_1502),
.Y(n_1594)
);

OA21x2_ASAP7_75t_L g1595 ( 
.A1(n_1436),
.A2(n_1472),
.B(n_1479),
.Y(n_1595)
);

INVx1_ASAP7_75t_L g1596 ( 
.A(n_1506),
.Y(n_1596)
);

NAND2x1p5_ASAP7_75t_L g1597 ( 
.A(n_1432),
.B(n_536),
.Y(n_1597)
);

AOI21x1_ASAP7_75t_L g1598 ( 
.A1(n_1441),
.A2(n_538),
.B(n_535),
.Y(n_1598)
);

OAI21xp5_ASAP7_75t_L g1599 ( 
.A1(n_1481),
.A2(n_540),
.B(n_539),
.Y(n_1599)
);

AO21x2_ASAP7_75t_L g1600 ( 
.A1(n_1500),
.A2(n_547),
.B(n_541),
.Y(n_1600)
);

OAI22xp33_ASAP7_75t_L g1601 ( 
.A1(n_1510),
.A2(n_1512),
.B1(n_1509),
.B2(n_1503),
.Y(n_1601)
);

AOI21xp5_ASAP7_75t_L g1602 ( 
.A1(n_1428),
.A2(n_549),
.B(n_548),
.Y(n_1602)
);

NOR2xp67_ASAP7_75t_L g1603 ( 
.A(n_1488),
.B(n_551),
.Y(n_1603)
);

OA21x2_ASAP7_75t_L g1604 ( 
.A1(n_1442),
.A2(n_554),
.B(n_553),
.Y(n_1604)
);

OAI21x1_ASAP7_75t_L g1605 ( 
.A1(n_1399),
.A2(n_556),
.B(n_555),
.Y(n_1605)
);

INVx1_ASAP7_75t_L g1606 ( 
.A(n_1397),
.Y(n_1606)
);

OAI21x1_ASAP7_75t_L g1607 ( 
.A1(n_1402),
.A2(n_559),
.B(n_557),
.Y(n_1607)
);

O2A1O1Ixp33_ASAP7_75t_L g1608 ( 
.A1(n_1395),
.A2(n_55),
.B(n_53),
.C(n_54),
.Y(n_1608)
);

NAND2x1_ASAP7_75t_L g1609 ( 
.A(n_1397),
.B(n_560),
.Y(n_1609)
);

INVx2_ASAP7_75t_L g1610 ( 
.A(n_1435),
.Y(n_1610)
);

AOI21xp5_ASAP7_75t_L g1611 ( 
.A1(n_1451),
.A2(n_562),
.B(n_561),
.Y(n_1611)
);

OAI22xp5_ASAP7_75t_L g1612 ( 
.A1(n_1449),
.A2(n_58),
.B1(n_56),
.B2(n_57),
.Y(n_1612)
);

INVx2_ASAP7_75t_L g1613 ( 
.A(n_1487),
.Y(n_1613)
);

BUFx6f_ASAP7_75t_L g1614 ( 
.A(n_1498),
.Y(n_1614)
);

OAI21x1_ASAP7_75t_L g1615 ( 
.A1(n_1410),
.A2(n_564),
.B(n_563),
.Y(n_1615)
);

NOR2x1_ASAP7_75t_SL g1616 ( 
.A(n_1493),
.B(n_1454),
.Y(n_1616)
);

NAND2xp5_ASAP7_75t_L g1617 ( 
.A(n_1498),
.B(n_56),
.Y(n_1617)
);

OAI21x1_ASAP7_75t_L g1618 ( 
.A1(n_1462),
.A2(n_566),
.B(n_565),
.Y(n_1618)
);

OR2x2_ASAP7_75t_L g1619 ( 
.A(n_1456),
.B(n_57),
.Y(n_1619)
);

NAND2xp5_ASAP7_75t_L g1620 ( 
.A(n_1511),
.B(n_1463),
.Y(n_1620)
);

INVx1_ASAP7_75t_L g1621 ( 
.A(n_1408),
.Y(n_1621)
);

OA21x2_ASAP7_75t_L g1622 ( 
.A1(n_1422),
.A2(n_570),
.B(n_568),
.Y(n_1622)
);

OAI21x1_ASAP7_75t_L g1623 ( 
.A1(n_1491),
.A2(n_573),
.B(n_571),
.Y(n_1623)
);

OAI21x1_ASAP7_75t_L g1624 ( 
.A1(n_1464),
.A2(n_576),
.B(n_575),
.Y(n_1624)
);

INVx1_ASAP7_75t_L g1625 ( 
.A(n_1408),
.Y(n_1625)
);

BUFx12f_ASAP7_75t_L g1626 ( 
.A(n_1423),
.Y(n_1626)
);

NOR2x1_ASAP7_75t_SL g1627 ( 
.A(n_1473),
.B(n_577),
.Y(n_1627)
);

OA21x2_ASAP7_75t_L g1628 ( 
.A1(n_1492),
.A2(n_582),
.B(n_578),
.Y(n_1628)
);

INVx1_ASAP7_75t_L g1629 ( 
.A(n_1489),
.Y(n_1629)
);

AND2x2_ASAP7_75t_L g1630 ( 
.A(n_1427),
.B(n_59),
.Y(n_1630)
);

OAI21x1_ASAP7_75t_L g1631 ( 
.A1(n_1426),
.A2(n_584),
.B(n_583),
.Y(n_1631)
);

BUFx2_ASAP7_75t_L g1632 ( 
.A(n_1416),
.Y(n_1632)
);

OAI21x1_ASAP7_75t_L g1633 ( 
.A1(n_1426),
.A2(n_586),
.B(n_585),
.Y(n_1633)
);

BUFx3_ASAP7_75t_L g1634 ( 
.A(n_1470),
.Y(n_1634)
);

INVx3_ASAP7_75t_L g1635 ( 
.A(n_1412),
.Y(n_1635)
);

NAND2xp5_ASAP7_75t_SL g1636 ( 
.A(n_1446),
.B(n_60),
.Y(n_1636)
);

INVx1_ASAP7_75t_L g1637 ( 
.A(n_1413),
.Y(n_1637)
);

INVx1_ASAP7_75t_L g1638 ( 
.A(n_1413),
.Y(n_1638)
);

NAND2xp5_ASAP7_75t_L g1639 ( 
.A(n_1400),
.B(n_61),
.Y(n_1639)
);

INVx1_ASAP7_75t_L g1640 ( 
.A(n_1413),
.Y(n_1640)
);

AOI21xp33_ASAP7_75t_L g1641 ( 
.A1(n_1407),
.A2(n_61),
.B(n_62),
.Y(n_1641)
);

AO31x2_ASAP7_75t_L g1642 ( 
.A1(n_1501),
.A2(n_588),
.A3(n_589),
.B(n_587),
.Y(n_1642)
);

AOI21xp5_ASAP7_75t_L g1643 ( 
.A1(n_1409),
.A2(n_591),
.B(n_590),
.Y(n_1643)
);

OAI21xp5_ASAP7_75t_L g1644 ( 
.A1(n_1534),
.A2(n_62),
.B(n_63),
.Y(n_1644)
);

AOI22xp33_ASAP7_75t_SL g1645 ( 
.A1(n_1578),
.A2(n_71),
.B1(n_79),
.B2(n_63),
.Y(n_1645)
);

OAI21x1_ASAP7_75t_L g1646 ( 
.A1(n_1527),
.A2(n_595),
.B(n_594),
.Y(n_1646)
);

BUFx3_ASAP7_75t_L g1647 ( 
.A(n_1572),
.Y(n_1647)
);

HB1xp67_ASAP7_75t_L g1648 ( 
.A(n_1539),
.Y(n_1648)
);

INVx2_ASAP7_75t_L g1649 ( 
.A(n_1540),
.Y(n_1649)
);

INVx1_ASAP7_75t_L g1650 ( 
.A(n_1528),
.Y(n_1650)
);

INVx1_ASAP7_75t_L g1651 ( 
.A(n_1637),
.Y(n_1651)
);

AOI21xp5_ASAP7_75t_L g1652 ( 
.A1(n_1595),
.A2(n_740),
.B(n_739),
.Y(n_1652)
);

BUFx10_ASAP7_75t_L g1653 ( 
.A(n_1576),
.Y(n_1653)
);

INVx2_ASAP7_75t_L g1654 ( 
.A(n_1555),
.Y(n_1654)
);

INVx1_ASAP7_75t_L g1655 ( 
.A(n_1638),
.Y(n_1655)
);

AOI22xp33_ASAP7_75t_L g1656 ( 
.A1(n_1601),
.A2(n_1577),
.B1(n_1641),
.B2(n_1547),
.Y(n_1656)
);

INVx1_ASAP7_75t_L g1657 ( 
.A(n_1640),
.Y(n_1657)
);

INVx1_ASAP7_75t_L g1658 ( 
.A(n_1541),
.Y(n_1658)
);

BUFx3_ASAP7_75t_L g1659 ( 
.A(n_1572),
.Y(n_1659)
);

AND2x2_ASAP7_75t_L g1660 ( 
.A(n_1537),
.B(n_64),
.Y(n_1660)
);

BUFx6f_ASAP7_75t_L g1661 ( 
.A(n_1579),
.Y(n_1661)
);

INVx2_ASAP7_75t_L g1662 ( 
.A(n_1538),
.Y(n_1662)
);

INVx4_ASAP7_75t_SL g1663 ( 
.A(n_1626),
.Y(n_1663)
);

BUFx2_ASAP7_75t_SL g1664 ( 
.A(n_1523),
.Y(n_1664)
);

INVx1_ASAP7_75t_L g1665 ( 
.A(n_1546),
.Y(n_1665)
);

INVx1_ASAP7_75t_L g1666 ( 
.A(n_1559),
.Y(n_1666)
);

AND2x4_ASAP7_75t_L g1667 ( 
.A(n_1549),
.B(n_596),
.Y(n_1667)
);

INVx1_ASAP7_75t_L g1668 ( 
.A(n_1562),
.Y(n_1668)
);

INVx2_ASAP7_75t_L g1669 ( 
.A(n_1535),
.Y(n_1669)
);

INVx2_ASAP7_75t_L g1670 ( 
.A(n_1565),
.Y(n_1670)
);

INVx2_ASAP7_75t_L g1671 ( 
.A(n_1586),
.Y(n_1671)
);

INVx1_ASAP7_75t_L g1672 ( 
.A(n_1594),
.Y(n_1672)
);

INVx1_ASAP7_75t_L g1673 ( 
.A(n_1596),
.Y(n_1673)
);

INVx2_ASAP7_75t_L g1674 ( 
.A(n_1521),
.Y(n_1674)
);

INVx1_ASAP7_75t_L g1675 ( 
.A(n_1639),
.Y(n_1675)
);

HB1xp67_ASAP7_75t_L g1676 ( 
.A(n_1568),
.Y(n_1676)
);

NOR2xp33_ASAP7_75t_SL g1677 ( 
.A(n_1548),
.B(n_597),
.Y(n_1677)
);

INVx2_ASAP7_75t_SL g1678 ( 
.A(n_1634),
.Y(n_1678)
);

BUFx6f_ASAP7_75t_L g1679 ( 
.A(n_1579),
.Y(n_1679)
);

BUFx8_ASAP7_75t_L g1680 ( 
.A(n_1545),
.Y(n_1680)
);

INVx1_ASAP7_75t_L g1681 ( 
.A(n_1590),
.Y(n_1681)
);

INVx3_ASAP7_75t_L g1682 ( 
.A(n_1635),
.Y(n_1682)
);

AO21x1_ASAP7_75t_L g1683 ( 
.A1(n_1608),
.A2(n_64),
.B(n_65),
.Y(n_1683)
);

NAND2xp5_ASAP7_75t_L g1684 ( 
.A(n_1564),
.B(n_1554),
.Y(n_1684)
);

INVx1_ASAP7_75t_L g1685 ( 
.A(n_1592),
.Y(n_1685)
);

BUFx2_ASAP7_75t_L g1686 ( 
.A(n_1557),
.Y(n_1686)
);

INVx1_ASAP7_75t_L g1687 ( 
.A(n_1619),
.Y(n_1687)
);

OR2x2_ASAP7_75t_L g1688 ( 
.A(n_1620),
.B(n_65),
.Y(n_1688)
);

NAND2x1p5_ASAP7_75t_L g1689 ( 
.A(n_1542),
.B(n_598),
.Y(n_1689)
);

HB1xp67_ASAP7_75t_L g1690 ( 
.A(n_1632),
.Y(n_1690)
);

HB1xp67_ASAP7_75t_L g1691 ( 
.A(n_1581),
.Y(n_1691)
);

BUFx2_ASAP7_75t_L g1692 ( 
.A(n_1575),
.Y(n_1692)
);

INVx1_ASAP7_75t_L g1693 ( 
.A(n_1606),
.Y(n_1693)
);

INVx1_ASAP7_75t_L g1694 ( 
.A(n_1589),
.Y(n_1694)
);

INVx1_ASAP7_75t_L g1695 ( 
.A(n_1533),
.Y(n_1695)
);

INVx1_ASAP7_75t_L g1696 ( 
.A(n_1533),
.Y(n_1696)
);

AOI21x1_ASAP7_75t_L g1697 ( 
.A1(n_1621),
.A2(n_600),
.B(n_599),
.Y(n_1697)
);

AND2x2_ASAP7_75t_L g1698 ( 
.A(n_1630),
.B(n_1566),
.Y(n_1698)
);

NAND3xp33_ASAP7_75t_L g1699 ( 
.A(n_1522),
.B(n_66),
.C(n_67),
.Y(n_1699)
);

INVx1_ASAP7_75t_L g1700 ( 
.A(n_1642),
.Y(n_1700)
);

HB1xp67_ASAP7_75t_L g1701 ( 
.A(n_1583),
.Y(n_1701)
);

OAI21x1_ASAP7_75t_L g1702 ( 
.A1(n_1631),
.A2(n_1633),
.B(n_1531),
.Y(n_1702)
);

INVx1_ASAP7_75t_L g1703 ( 
.A(n_1642),
.Y(n_1703)
);

INVx1_ASAP7_75t_L g1704 ( 
.A(n_1625),
.Y(n_1704)
);

INVx1_ASAP7_75t_SL g1705 ( 
.A(n_1584),
.Y(n_1705)
);

INVx2_ASAP7_75t_SL g1706 ( 
.A(n_1583),
.Y(n_1706)
);

INVx1_ASAP7_75t_L g1707 ( 
.A(n_1598),
.Y(n_1707)
);

INVx1_ASAP7_75t_L g1708 ( 
.A(n_1515),
.Y(n_1708)
);

INVx1_ASAP7_75t_L g1709 ( 
.A(n_1543),
.Y(n_1709)
);

INVx1_ASAP7_75t_L g1710 ( 
.A(n_1543),
.Y(n_1710)
);

INVx2_ASAP7_75t_L g1711 ( 
.A(n_1570),
.Y(n_1711)
);

INVx3_ASAP7_75t_L g1712 ( 
.A(n_1585),
.Y(n_1712)
);

INVx4_ASAP7_75t_SL g1713 ( 
.A(n_1614),
.Y(n_1713)
);

OAI22xp5_ASAP7_75t_L g1714 ( 
.A1(n_1520),
.A2(n_69),
.B1(n_66),
.B2(n_68),
.Y(n_1714)
);

INVx3_ASAP7_75t_SL g1715 ( 
.A(n_1614),
.Y(n_1715)
);

HB1xp67_ASAP7_75t_L g1716 ( 
.A(n_1636),
.Y(n_1716)
);

INVx1_ASAP7_75t_L g1717 ( 
.A(n_1580),
.Y(n_1717)
);

INVx1_ASAP7_75t_L g1718 ( 
.A(n_1516),
.Y(n_1718)
);

INVx2_ASAP7_75t_L g1719 ( 
.A(n_1597),
.Y(n_1719)
);

NAND2xp5_ASAP7_75t_L g1720 ( 
.A(n_1574),
.B(n_68),
.Y(n_1720)
);

INVx1_ASAP7_75t_L g1721 ( 
.A(n_1551),
.Y(n_1721)
);

BUFx6f_ASAP7_75t_L g1722 ( 
.A(n_1609),
.Y(n_1722)
);

NOR2xp33_ASAP7_75t_L g1723 ( 
.A(n_1593),
.B(n_601),
.Y(n_1723)
);

INVx1_ASAP7_75t_L g1724 ( 
.A(n_1551),
.Y(n_1724)
);

INVx1_ASAP7_75t_L g1725 ( 
.A(n_1544),
.Y(n_1725)
);

NOR2xp33_ASAP7_75t_R g1726 ( 
.A(n_1712),
.B(n_1617),
.Y(n_1726)
);

CKINVDCx16_ASAP7_75t_R g1727 ( 
.A(n_1653),
.Y(n_1727)
);

AND2x2_ASAP7_75t_L g1728 ( 
.A(n_1698),
.B(n_1550),
.Y(n_1728)
);

NAND2xp33_ASAP7_75t_R g1729 ( 
.A(n_1692),
.B(n_1628),
.Y(n_1729)
);

AND2x2_ASAP7_75t_L g1730 ( 
.A(n_1694),
.B(n_1526),
.Y(n_1730)
);

NAND2xp5_ASAP7_75t_L g1731 ( 
.A(n_1684),
.B(n_1563),
.Y(n_1731)
);

INVx1_ASAP7_75t_L g1732 ( 
.A(n_1658),
.Y(n_1732)
);

INVx1_ASAP7_75t_L g1733 ( 
.A(n_1665),
.Y(n_1733)
);

INVxp67_ASAP7_75t_L g1734 ( 
.A(n_1676),
.Y(n_1734)
);

NOR2xp33_ASAP7_75t_R g1735 ( 
.A(n_1715),
.B(n_1629),
.Y(n_1735)
);

NAND2xp33_ASAP7_75t_SL g1736 ( 
.A(n_1661),
.B(n_1612),
.Y(n_1736)
);

AND2x2_ASAP7_75t_L g1737 ( 
.A(n_1687),
.B(n_1571),
.Y(n_1737)
);

NOR2xp33_ASAP7_75t_R g1738 ( 
.A(n_1647),
.B(n_603),
.Y(n_1738)
);

XNOR2xp5_ASAP7_75t_L g1739 ( 
.A(n_1705),
.B(n_1588),
.Y(n_1739)
);

XNOR2xp5_ASAP7_75t_L g1740 ( 
.A(n_1678),
.B(n_1552),
.Y(n_1740)
);

NAND2xp5_ASAP7_75t_L g1741 ( 
.A(n_1675),
.B(n_1525),
.Y(n_1741)
);

AND2x4_ASAP7_75t_L g1742 ( 
.A(n_1659),
.B(n_1603),
.Y(n_1742)
);

NOR2xp33_ASAP7_75t_R g1743 ( 
.A(n_1661),
.B(n_604),
.Y(n_1743)
);

INVx2_ASAP7_75t_SL g1744 ( 
.A(n_1679),
.Y(n_1744)
);

NAND2xp5_ASAP7_75t_L g1745 ( 
.A(n_1681),
.B(n_1556),
.Y(n_1745)
);

NOR2xp33_ASAP7_75t_L g1746 ( 
.A(n_1723),
.B(n_1573),
.Y(n_1746)
);

NAND2xp5_ASAP7_75t_L g1747 ( 
.A(n_1685),
.B(n_1518),
.Y(n_1747)
);

INVx1_ASAP7_75t_L g1748 ( 
.A(n_1666),
.Y(n_1748)
);

AND2x2_ASAP7_75t_L g1749 ( 
.A(n_1660),
.B(n_1519),
.Y(n_1749)
);

OR2x6_ASAP7_75t_L g1750 ( 
.A(n_1664),
.B(n_1643),
.Y(n_1750)
);

INVxp67_ASAP7_75t_L g1751 ( 
.A(n_1648),
.Y(n_1751)
);

AND2x2_ASAP7_75t_L g1752 ( 
.A(n_1670),
.B(n_1671),
.Y(n_1752)
);

AND2x4_ASAP7_75t_L g1753 ( 
.A(n_1713),
.B(n_1624),
.Y(n_1753)
);

BUFx3_ASAP7_75t_L g1754 ( 
.A(n_1679),
.Y(n_1754)
);

AND2x4_ASAP7_75t_L g1755 ( 
.A(n_1713),
.B(n_1517),
.Y(n_1755)
);

CKINVDCx5p33_ASAP7_75t_R g1756 ( 
.A(n_1680),
.Y(n_1756)
);

CKINVDCx8_ASAP7_75t_R g1757 ( 
.A(n_1663),
.Y(n_1757)
);

AND2x2_ASAP7_75t_L g1758 ( 
.A(n_1649),
.B(n_1561),
.Y(n_1758)
);

NAND2xp5_ASAP7_75t_L g1759 ( 
.A(n_1672),
.B(n_1627),
.Y(n_1759)
);

AND2x4_ASAP7_75t_L g1760 ( 
.A(n_1706),
.B(n_1623),
.Y(n_1760)
);

NOR2xp33_ASAP7_75t_R g1761 ( 
.A(n_1677),
.B(n_606),
.Y(n_1761)
);

NAND2xp33_ASAP7_75t_R g1762 ( 
.A(n_1686),
.B(n_1567),
.Y(n_1762)
);

AND2x4_ASAP7_75t_L g1763 ( 
.A(n_1701),
.B(n_1618),
.Y(n_1763)
);

INVxp67_ASAP7_75t_SL g1764 ( 
.A(n_1673),
.Y(n_1764)
);

OR2x4_ASAP7_75t_L g1765 ( 
.A(n_1688),
.B(n_1591),
.Y(n_1765)
);

AND2x2_ASAP7_75t_L g1766 ( 
.A(n_1654),
.B(n_1599),
.Y(n_1766)
);

AND2x4_ASAP7_75t_L g1767 ( 
.A(n_1690),
.B(n_1667),
.Y(n_1767)
);

NAND2xp5_ASAP7_75t_L g1768 ( 
.A(n_1716),
.B(n_1529),
.Y(n_1768)
);

NAND2xp5_ASAP7_75t_L g1769 ( 
.A(n_1644),
.B(n_1587),
.Y(n_1769)
);

OR2x2_ASAP7_75t_L g1770 ( 
.A(n_1669),
.B(n_1587),
.Y(n_1770)
);

BUFx3_ASAP7_75t_L g1771 ( 
.A(n_1682),
.Y(n_1771)
);

NAND2xp5_ASAP7_75t_L g1772 ( 
.A(n_1662),
.B(n_1600),
.Y(n_1772)
);

OR2x6_ASAP7_75t_L g1773 ( 
.A(n_1722),
.B(n_1602),
.Y(n_1773)
);

AND2x2_ASAP7_75t_L g1774 ( 
.A(n_1650),
.B(n_1569),
.Y(n_1774)
);

INVx1_ASAP7_75t_L g1775 ( 
.A(n_1732),
.Y(n_1775)
);

OR2x2_ASAP7_75t_L g1776 ( 
.A(n_1734),
.B(n_1704),
.Y(n_1776)
);

BUFx2_ASAP7_75t_L g1777 ( 
.A(n_1735),
.Y(n_1777)
);

NAND2xp5_ASAP7_75t_L g1778 ( 
.A(n_1751),
.B(n_1668),
.Y(n_1778)
);

INVx2_ASAP7_75t_L g1779 ( 
.A(n_1752),
.Y(n_1779)
);

INVx1_ASAP7_75t_L g1780 ( 
.A(n_1764),
.Y(n_1780)
);

HB1xp67_ASAP7_75t_L g1781 ( 
.A(n_1770),
.Y(n_1781)
);

INVx1_ASAP7_75t_L g1782 ( 
.A(n_1733),
.Y(n_1782)
);

AOI22xp33_ASAP7_75t_SL g1783 ( 
.A1(n_1728),
.A2(n_1699),
.B1(n_1714),
.B2(n_1720),
.Y(n_1783)
);

INVxp67_ASAP7_75t_SL g1784 ( 
.A(n_1747),
.Y(n_1784)
);

INVxp67_ASAP7_75t_SL g1785 ( 
.A(n_1772),
.Y(n_1785)
);

AOI22xp33_ASAP7_75t_L g1786 ( 
.A1(n_1736),
.A2(n_1656),
.B1(n_1683),
.B2(n_1725),
.Y(n_1786)
);

NAND2xp5_ASAP7_75t_L g1787 ( 
.A(n_1748),
.B(n_1651),
.Y(n_1787)
);

AND2x4_ASAP7_75t_L g1788 ( 
.A(n_1749),
.B(n_1693),
.Y(n_1788)
);

NOR3xp33_ASAP7_75t_L g1789 ( 
.A(n_1746),
.B(n_1645),
.C(n_1708),
.Y(n_1789)
);

AND2x2_ASAP7_75t_L g1790 ( 
.A(n_1737),
.B(n_1691),
.Y(n_1790)
);

NAND2xp5_ASAP7_75t_SL g1791 ( 
.A(n_1726),
.B(n_1722),
.Y(n_1791)
);

INVx2_ASAP7_75t_L g1792 ( 
.A(n_1774),
.Y(n_1792)
);

AND2x2_ASAP7_75t_L g1793 ( 
.A(n_1767),
.B(n_1655),
.Y(n_1793)
);

INVxp33_ASAP7_75t_L g1794 ( 
.A(n_1740),
.Y(n_1794)
);

AND2x2_ASAP7_75t_L g1795 ( 
.A(n_1730),
.B(n_1657),
.Y(n_1795)
);

NAND2xp5_ASAP7_75t_L g1796 ( 
.A(n_1731),
.B(n_1717),
.Y(n_1796)
);

AND2x4_ASAP7_75t_L g1797 ( 
.A(n_1755),
.B(n_1711),
.Y(n_1797)
);

INVx1_ASAP7_75t_L g1798 ( 
.A(n_1759),
.Y(n_1798)
);

INVx1_ASAP7_75t_L g1799 ( 
.A(n_1758),
.Y(n_1799)
);

AND2x2_ASAP7_75t_L g1800 ( 
.A(n_1763),
.B(n_1674),
.Y(n_1800)
);

NAND2xp5_ASAP7_75t_L g1801 ( 
.A(n_1741),
.B(n_1707),
.Y(n_1801)
);

INVx3_ASAP7_75t_L g1802 ( 
.A(n_1760),
.Y(n_1802)
);

NAND2xp5_ASAP7_75t_L g1803 ( 
.A(n_1745),
.B(n_1709),
.Y(n_1803)
);

OAI21xp5_ASAP7_75t_SL g1804 ( 
.A1(n_1739),
.A2(n_1689),
.B(n_1611),
.Y(n_1804)
);

AND2x2_ASAP7_75t_L g1805 ( 
.A(n_1766),
.B(n_1721),
.Y(n_1805)
);

AND2x2_ASAP7_75t_L g1806 ( 
.A(n_1744),
.B(n_1754),
.Y(n_1806)
);

AOI22xp33_ASAP7_75t_SL g1807 ( 
.A1(n_1761),
.A2(n_1616),
.B1(n_1530),
.B2(n_1719),
.Y(n_1807)
);

INVx2_ASAP7_75t_L g1808 ( 
.A(n_1768),
.Y(n_1808)
);

INVx1_ASAP7_75t_L g1809 ( 
.A(n_1769),
.Y(n_1809)
);

INVx2_ASAP7_75t_L g1810 ( 
.A(n_1750),
.Y(n_1810)
);

INVx1_ASAP7_75t_L g1811 ( 
.A(n_1765),
.Y(n_1811)
);

NAND2xp5_ASAP7_75t_L g1812 ( 
.A(n_1742),
.B(n_1710),
.Y(n_1812)
);

AND2x2_ASAP7_75t_L g1813 ( 
.A(n_1771),
.B(n_1724),
.Y(n_1813)
);

INVxp67_ASAP7_75t_L g1814 ( 
.A(n_1729),
.Y(n_1814)
);

AND2x2_ASAP7_75t_L g1815 ( 
.A(n_1727),
.B(n_1695),
.Y(n_1815)
);

INVx1_ASAP7_75t_L g1816 ( 
.A(n_1750),
.Y(n_1816)
);

NAND2xp5_ASAP7_75t_L g1817 ( 
.A(n_1738),
.B(n_1696),
.Y(n_1817)
);

INVx1_ASAP7_75t_L g1818 ( 
.A(n_1753),
.Y(n_1818)
);

AOI22xp33_ASAP7_75t_L g1819 ( 
.A1(n_1743),
.A2(n_1703),
.B1(n_1700),
.B2(n_1604),
.Y(n_1819)
);

HB1xp67_ASAP7_75t_L g1820 ( 
.A(n_1762),
.Y(n_1820)
);

INVx1_ASAP7_75t_L g1821 ( 
.A(n_1773),
.Y(n_1821)
);

INVx1_ASAP7_75t_L g1822 ( 
.A(n_1773),
.Y(n_1822)
);

INVx1_ASAP7_75t_L g1823 ( 
.A(n_1757),
.Y(n_1823)
);

INVx1_ASAP7_75t_L g1824 ( 
.A(n_1756),
.Y(n_1824)
);

NAND2xp5_ASAP7_75t_L g1825 ( 
.A(n_1808),
.B(n_1718),
.Y(n_1825)
);

INVx1_ASAP7_75t_L g1826 ( 
.A(n_1775),
.Y(n_1826)
);

INVx1_ASAP7_75t_L g1827 ( 
.A(n_1775),
.Y(n_1827)
);

AND2x4_ASAP7_75t_L g1828 ( 
.A(n_1810),
.B(n_1663),
.Y(n_1828)
);

INVxp67_ASAP7_75t_L g1829 ( 
.A(n_1790),
.Y(n_1829)
);

AND2x2_ASAP7_75t_L g1830 ( 
.A(n_1815),
.B(n_1646),
.Y(n_1830)
);

INVx2_ASAP7_75t_L g1831 ( 
.A(n_1782),
.Y(n_1831)
);

NAND2xp5_ASAP7_75t_L g1832 ( 
.A(n_1798),
.B(n_1652),
.Y(n_1832)
);

INVx4_ASAP7_75t_L g1833 ( 
.A(n_1777),
.Y(n_1833)
);

INVx1_ASAP7_75t_L g1834 ( 
.A(n_1780),
.Y(n_1834)
);

AOI211xp5_ASAP7_75t_SL g1835 ( 
.A1(n_1814),
.A2(n_1610),
.B(n_1613),
.C(n_1697),
.Y(n_1835)
);

AND2x4_ASAP7_75t_L g1836 ( 
.A(n_1816),
.B(n_1702),
.Y(n_1836)
);

AND2x2_ASAP7_75t_L g1837 ( 
.A(n_1820),
.B(n_1524),
.Y(n_1837)
);

HB1xp67_ASAP7_75t_L g1838 ( 
.A(n_1781),
.Y(n_1838)
);

INVx1_ASAP7_75t_L g1839 ( 
.A(n_1776),
.Y(n_1839)
);

INVx1_ASAP7_75t_L g1840 ( 
.A(n_1787),
.Y(n_1840)
);

AND2x2_ASAP7_75t_L g1841 ( 
.A(n_1779),
.B(n_1532),
.Y(n_1841)
);

OAI31xp33_ASAP7_75t_L g1842 ( 
.A1(n_1804),
.A2(n_72),
.A3(n_70),
.B(n_71),
.Y(n_1842)
);

INVx1_ASAP7_75t_L g1843 ( 
.A(n_1778),
.Y(n_1843)
);

AOI22xp33_ASAP7_75t_L g1844 ( 
.A1(n_1789),
.A2(n_1622),
.B1(n_1605),
.B2(n_1615),
.Y(n_1844)
);

AOI211xp5_ASAP7_75t_L g1845 ( 
.A1(n_1811),
.A2(n_1607),
.B(n_1536),
.C(n_1558),
.Y(n_1845)
);

INVx3_ASAP7_75t_L g1846 ( 
.A(n_1806),
.Y(n_1846)
);

AND2x2_ASAP7_75t_L g1847 ( 
.A(n_1793),
.B(n_1553),
.Y(n_1847)
);

INVx2_ASAP7_75t_L g1848 ( 
.A(n_1788),
.Y(n_1848)
);

INVx1_ASAP7_75t_L g1849 ( 
.A(n_1809),
.Y(n_1849)
);

AND2x4_ASAP7_75t_SL g1850 ( 
.A(n_1800),
.B(n_1560),
.Y(n_1850)
);

INVx2_ASAP7_75t_L g1851 ( 
.A(n_1788),
.Y(n_1851)
);

AND2x2_ASAP7_75t_L g1852 ( 
.A(n_1799),
.B(n_1582),
.Y(n_1852)
);

AND2x2_ASAP7_75t_L g1853 ( 
.A(n_1802),
.B(n_70),
.Y(n_1853)
);

HB1xp67_ASAP7_75t_L g1854 ( 
.A(n_1792),
.Y(n_1854)
);

OR2x2_ASAP7_75t_L g1855 ( 
.A(n_1785),
.B(n_72),
.Y(n_1855)
);

INVx2_ASAP7_75t_L g1856 ( 
.A(n_1813),
.Y(n_1856)
);

INVx2_ASAP7_75t_L g1857 ( 
.A(n_1818),
.Y(n_1857)
);

AND2x2_ASAP7_75t_L g1858 ( 
.A(n_1795),
.B(n_73),
.Y(n_1858)
);

AND2x2_ASAP7_75t_L g1859 ( 
.A(n_1805),
.B(n_73),
.Y(n_1859)
);

AND2x2_ASAP7_75t_L g1860 ( 
.A(n_1821),
.B(n_74),
.Y(n_1860)
);

AND2x2_ASAP7_75t_L g1861 ( 
.A(n_1822),
.B(n_74),
.Y(n_1861)
);

OR2x2_ASAP7_75t_L g1862 ( 
.A(n_1784),
.B(n_75),
.Y(n_1862)
);

NOR2xp33_ASAP7_75t_L g1863 ( 
.A(n_1794),
.B(n_75),
.Y(n_1863)
);

INVx1_ASAP7_75t_L g1864 ( 
.A(n_1803),
.Y(n_1864)
);

BUFx3_ASAP7_75t_L g1865 ( 
.A(n_1823),
.Y(n_1865)
);

NAND4xp25_ASAP7_75t_L g1866 ( 
.A(n_1786),
.B(n_78),
.C(n_76),
.D(n_77),
.Y(n_1866)
);

NOR2x1_ASAP7_75t_SL g1867 ( 
.A(n_1791),
.B(n_77),
.Y(n_1867)
);

AND2x2_ASAP7_75t_L g1868 ( 
.A(n_1812),
.B(n_76),
.Y(n_1868)
);

INVx1_ASAP7_75t_L g1869 ( 
.A(n_1801),
.Y(n_1869)
);

HB1xp67_ASAP7_75t_L g1870 ( 
.A(n_1797),
.Y(n_1870)
);

NAND2xp5_ASAP7_75t_L g1871 ( 
.A(n_1796),
.B(n_78),
.Y(n_1871)
);

NAND2xp5_ASAP7_75t_L g1872 ( 
.A(n_1797),
.B(n_80),
.Y(n_1872)
);

OR2x2_ASAP7_75t_L g1873 ( 
.A(n_1817),
.B(n_80),
.Y(n_1873)
);

AND2x2_ASAP7_75t_L g1874 ( 
.A(n_1824),
.B(n_81),
.Y(n_1874)
);

OR2x2_ASAP7_75t_L g1875 ( 
.A(n_1819),
.B(n_81),
.Y(n_1875)
);

INVx1_ASAP7_75t_L g1876 ( 
.A(n_1807),
.Y(n_1876)
);

INVx1_ASAP7_75t_L g1877 ( 
.A(n_1783),
.Y(n_1877)
);

BUFx2_ASAP7_75t_L g1878 ( 
.A(n_1811),
.Y(n_1878)
);

NAND2xp5_ASAP7_75t_L g1879 ( 
.A(n_1808),
.B(n_82),
.Y(n_1879)
);

CKINVDCx20_ASAP7_75t_R g1880 ( 
.A(n_1777),
.Y(n_1880)
);

INVx1_ASAP7_75t_L g1881 ( 
.A(n_1775),
.Y(n_1881)
);

NAND2xp5_ASAP7_75t_L g1882 ( 
.A(n_1808),
.B(n_82),
.Y(n_1882)
);

INVx1_ASAP7_75t_L g1883 ( 
.A(n_1775),
.Y(n_1883)
);

NOR2xp33_ASAP7_75t_L g1884 ( 
.A(n_1794),
.B(n_83),
.Y(n_1884)
);

NOR2x1p5_ASAP7_75t_L g1885 ( 
.A(n_1811),
.B(n_83),
.Y(n_1885)
);

NAND2xp5_ASAP7_75t_L g1886 ( 
.A(n_1808),
.B(n_84),
.Y(n_1886)
);

AOI221xp5_ASAP7_75t_L g1887 ( 
.A1(n_1789),
.A2(n_86),
.B1(n_84),
.B2(n_85),
.C(n_87),
.Y(n_1887)
);

OR2x2_ASAP7_75t_L g1888 ( 
.A(n_1785),
.B(n_85),
.Y(n_1888)
);

AOI22xp33_ASAP7_75t_L g1889 ( 
.A1(n_1789),
.A2(n_89),
.B1(n_87),
.B2(n_88),
.Y(n_1889)
);

AND2x2_ASAP7_75t_L g1890 ( 
.A(n_1815),
.B(n_88),
.Y(n_1890)
);

INVx1_ASAP7_75t_L g1891 ( 
.A(n_1775),
.Y(n_1891)
);

NAND2xp5_ASAP7_75t_L g1892 ( 
.A(n_1808),
.B(n_90),
.Y(n_1892)
);

INVx2_ASAP7_75t_SL g1893 ( 
.A(n_1806),
.Y(n_1893)
);

OAI21xp5_ASAP7_75t_L g1894 ( 
.A1(n_1804),
.A2(n_91),
.B(n_92),
.Y(n_1894)
);

INVx1_ASAP7_75t_L g1895 ( 
.A(n_1775),
.Y(n_1895)
);

NOR2x1_ASAP7_75t_L g1896 ( 
.A(n_1833),
.B(n_91),
.Y(n_1896)
);

INVx2_ASAP7_75t_L g1897 ( 
.A(n_1849),
.Y(n_1897)
);

NAND2xp5_ASAP7_75t_L g1898 ( 
.A(n_1869),
.B(n_92),
.Y(n_1898)
);

AND2x2_ASAP7_75t_L g1899 ( 
.A(n_1848),
.B(n_93),
.Y(n_1899)
);

AND2x2_ASAP7_75t_L g1900 ( 
.A(n_1851),
.B(n_93),
.Y(n_1900)
);

NOR2x1p5_ASAP7_75t_L g1901 ( 
.A(n_1876),
.B(n_94),
.Y(n_1901)
);

OR2x2_ASAP7_75t_L g1902 ( 
.A(n_1838),
.B(n_94),
.Y(n_1902)
);

NOR2xp33_ASAP7_75t_L g1903 ( 
.A(n_1833),
.B(n_95),
.Y(n_1903)
);

AND2x2_ASAP7_75t_L g1904 ( 
.A(n_1856),
.B(n_95),
.Y(n_1904)
);

AND2x4_ASAP7_75t_L g1905 ( 
.A(n_1878),
.B(n_97),
.Y(n_1905)
);

OR2x2_ASAP7_75t_L g1906 ( 
.A(n_1839),
.B(n_97),
.Y(n_1906)
);

BUFx2_ASAP7_75t_L g1907 ( 
.A(n_1870),
.Y(n_1907)
);

BUFx2_ASAP7_75t_L g1908 ( 
.A(n_1846),
.Y(n_1908)
);

OR2x2_ASAP7_75t_L g1909 ( 
.A(n_1854),
.B(n_1829),
.Y(n_1909)
);

INVx1_ASAP7_75t_L g1910 ( 
.A(n_1826),
.Y(n_1910)
);

NAND2xp5_ASAP7_75t_L g1911 ( 
.A(n_1843),
.B(n_98),
.Y(n_1911)
);

INVx3_ASAP7_75t_L g1912 ( 
.A(n_1828),
.Y(n_1912)
);

INVxp67_ASAP7_75t_L g1913 ( 
.A(n_1873),
.Y(n_1913)
);

INVx1_ASAP7_75t_L g1914 ( 
.A(n_1827),
.Y(n_1914)
);

OR2x2_ASAP7_75t_L g1915 ( 
.A(n_1834),
.B(n_99),
.Y(n_1915)
);

INVx1_ASAP7_75t_L g1916 ( 
.A(n_1881),
.Y(n_1916)
);

INVx1_ASAP7_75t_L g1917 ( 
.A(n_1883),
.Y(n_1917)
);

AND2x2_ASAP7_75t_L g1918 ( 
.A(n_1893),
.B(n_99),
.Y(n_1918)
);

INVx1_ASAP7_75t_L g1919 ( 
.A(n_1891),
.Y(n_1919)
);

AND2x2_ASAP7_75t_L g1920 ( 
.A(n_1857),
.B(n_100),
.Y(n_1920)
);

AND2x2_ASAP7_75t_L g1921 ( 
.A(n_1840),
.B(n_100),
.Y(n_1921)
);

INVx1_ASAP7_75t_L g1922 ( 
.A(n_1895),
.Y(n_1922)
);

INVx2_ASAP7_75t_L g1923 ( 
.A(n_1831),
.Y(n_1923)
);

AND2x2_ASAP7_75t_L g1924 ( 
.A(n_1864),
.B(n_101),
.Y(n_1924)
);

INVx2_ASAP7_75t_SL g1925 ( 
.A(n_1865),
.Y(n_1925)
);

NAND2xp5_ASAP7_75t_L g1926 ( 
.A(n_1832),
.B(n_101),
.Y(n_1926)
);

NAND2xp5_ASAP7_75t_L g1927 ( 
.A(n_1825),
.B(n_102),
.Y(n_1927)
);

INVx2_ASAP7_75t_L g1928 ( 
.A(n_1836),
.Y(n_1928)
);

AND2x2_ASAP7_75t_L g1929 ( 
.A(n_1828),
.B(n_103),
.Y(n_1929)
);

NOR2x1_ASAP7_75t_SL g1930 ( 
.A(n_1830),
.B(n_103),
.Y(n_1930)
);

INVx1_ASAP7_75t_L g1931 ( 
.A(n_1836),
.Y(n_1931)
);

NAND2xp5_ASAP7_75t_L g1932 ( 
.A(n_1868),
.B(n_104),
.Y(n_1932)
);

NAND2xp5_ASAP7_75t_L g1933 ( 
.A(n_1877),
.B(n_104),
.Y(n_1933)
);

AND2x4_ASAP7_75t_L g1934 ( 
.A(n_1847),
.B(n_105),
.Y(n_1934)
);

INVx1_ASAP7_75t_SL g1935 ( 
.A(n_1880),
.Y(n_1935)
);

NAND2xp5_ASAP7_75t_L g1936 ( 
.A(n_1837),
.B(n_105),
.Y(n_1936)
);

INVx1_ASAP7_75t_L g1937 ( 
.A(n_1862),
.Y(n_1937)
);

INVx1_ASAP7_75t_SL g1938 ( 
.A(n_1874),
.Y(n_1938)
);

NAND2xp5_ASAP7_75t_L g1939 ( 
.A(n_1855),
.B(n_106),
.Y(n_1939)
);

INVx1_ASAP7_75t_L g1940 ( 
.A(n_1888),
.Y(n_1940)
);

INVx2_ASAP7_75t_L g1941 ( 
.A(n_1841),
.Y(n_1941)
);

NOR2x1_ASAP7_75t_L g1942 ( 
.A(n_1871),
.B(n_106),
.Y(n_1942)
);

AND2x2_ASAP7_75t_L g1943 ( 
.A(n_1890),
.B(n_107),
.Y(n_1943)
);

NAND2xp5_ASAP7_75t_L g1944 ( 
.A(n_1852),
.B(n_108),
.Y(n_1944)
);

AND2x2_ASAP7_75t_L g1945 ( 
.A(n_1859),
.B(n_108),
.Y(n_1945)
);

HB1xp67_ASAP7_75t_L g1946 ( 
.A(n_1872),
.Y(n_1946)
);

NAND2x1p5_ASAP7_75t_L g1947 ( 
.A(n_1853),
.B(n_607),
.Y(n_1947)
);

NAND2xp5_ASAP7_75t_L g1948 ( 
.A(n_1858),
.B(n_109),
.Y(n_1948)
);

NAND2xp5_ASAP7_75t_L g1949 ( 
.A(n_1879),
.B(n_109),
.Y(n_1949)
);

NAND2xp5_ASAP7_75t_L g1950 ( 
.A(n_1882),
.B(n_110),
.Y(n_1950)
);

OR2x2_ASAP7_75t_L g1951 ( 
.A(n_1886),
.B(n_111),
.Y(n_1951)
);

AND2x2_ASAP7_75t_L g1952 ( 
.A(n_1860),
.B(n_112),
.Y(n_1952)
);

AND2x2_ASAP7_75t_L g1953 ( 
.A(n_1861),
.B(n_112),
.Y(n_1953)
);

OR2x2_ASAP7_75t_L g1954 ( 
.A(n_1892),
.B(n_113),
.Y(n_1954)
);

NAND2xp5_ASAP7_75t_L g1955 ( 
.A(n_1875),
.B(n_114),
.Y(n_1955)
);

INVx1_ASAP7_75t_L g1956 ( 
.A(n_1850),
.Y(n_1956)
);

AND2x2_ASAP7_75t_L g1957 ( 
.A(n_1885),
.B(n_115),
.Y(n_1957)
);

INVx1_ASAP7_75t_L g1958 ( 
.A(n_1867),
.Y(n_1958)
);

AND2x2_ASAP7_75t_L g1959 ( 
.A(n_1863),
.B(n_116),
.Y(n_1959)
);

NOR2x1p5_ASAP7_75t_L g1960 ( 
.A(n_1866),
.B(n_116),
.Y(n_1960)
);

INVx2_ASAP7_75t_L g1961 ( 
.A(n_1884),
.Y(n_1961)
);

INVx1_ASAP7_75t_L g1962 ( 
.A(n_1845),
.Y(n_1962)
);

AND2x2_ASAP7_75t_L g1963 ( 
.A(n_1894),
.B(n_117),
.Y(n_1963)
);

AND2x2_ASAP7_75t_L g1964 ( 
.A(n_1835),
.B(n_117),
.Y(n_1964)
);

INVxp33_ASAP7_75t_L g1965 ( 
.A(n_1842),
.Y(n_1965)
);

AND2x2_ASAP7_75t_L g1966 ( 
.A(n_1844),
.B(n_118),
.Y(n_1966)
);

HB1xp67_ASAP7_75t_L g1967 ( 
.A(n_1887),
.Y(n_1967)
);

INVx1_ASAP7_75t_L g1968 ( 
.A(n_1889),
.Y(n_1968)
);

OR2x2_ASAP7_75t_L g1969 ( 
.A(n_1838),
.B(n_118),
.Y(n_1969)
);

AND2x2_ASAP7_75t_L g1970 ( 
.A(n_1848),
.B(n_119),
.Y(n_1970)
);

AND2x2_ASAP7_75t_L g1971 ( 
.A(n_1848),
.B(n_119),
.Y(n_1971)
);

NAND2xp5_ASAP7_75t_L g1972 ( 
.A(n_1869),
.B(n_120),
.Y(n_1972)
);

AND2x2_ASAP7_75t_L g1973 ( 
.A(n_1848),
.B(n_120),
.Y(n_1973)
);

AND2x2_ASAP7_75t_L g1974 ( 
.A(n_1848),
.B(n_121),
.Y(n_1974)
);

NAND2xp5_ASAP7_75t_L g1975 ( 
.A(n_1869),
.B(n_121),
.Y(n_1975)
);

INVx1_ASAP7_75t_L g1976 ( 
.A(n_1826),
.Y(n_1976)
);

INVx1_ASAP7_75t_L g1977 ( 
.A(n_1826),
.Y(n_1977)
);

NAND2xp5_ASAP7_75t_L g1978 ( 
.A(n_1869),
.B(n_122),
.Y(n_1978)
);

INVx1_ASAP7_75t_L g1979 ( 
.A(n_1826),
.Y(n_1979)
);

BUFx3_ASAP7_75t_L g1980 ( 
.A(n_1880),
.Y(n_1980)
);

AND2x2_ASAP7_75t_L g1981 ( 
.A(n_1848),
.B(n_122),
.Y(n_1981)
);

INVx1_ASAP7_75t_L g1982 ( 
.A(n_1826),
.Y(n_1982)
);

NAND2xp5_ASAP7_75t_SL g1983 ( 
.A(n_1833),
.B(n_123),
.Y(n_1983)
);

NAND2xp5_ASAP7_75t_L g1984 ( 
.A(n_1869),
.B(n_123),
.Y(n_1984)
);

NOR2xp33_ASAP7_75t_L g1985 ( 
.A(n_1833),
.B(n_124),
.Y(n_1985)
);

NAND2xp5_ASAP7_75t_L g1986 ( 
.A(n_1946),
.B(n_124),
.Y(n_1986)
);

OAI221xp5_ASAP7_75t_L g1987 ( 
.A1(n_1967),
.A2(n_127),
.B1(n_125),
.B2(n_126),
.C(n_128),
.Y(n_1987)
);

INVxp33_ASAP7_75t_SL g1988 ( 
.A(n_1935),
.Y(n_1988)
);

INVx3_ASAP7_75t_L g1989 ( 
.A(n_1912),
.Y(n_1989)
);

NAND2xp33_ASAP7_75t_SL g1990 ( 
.A(n_1901),
.B(n_1965),
.Y(n_1990)
);

NAND2xp5_ASAP7_75t_L g1991 ( 
.A(n_1962),
.B(n_126),
.Y(n_1991)
);

OR2x2_ASAP7_75t_L g1992 ( 
.A(n_1909),
.B(n_1907),
.Y(n_1992)
);

INVx1_ASAP7_75t_SL g1993 ( 
.A(n_1980),
.Y(n_1993)
);

NAND2xp5_ASAP7_75t_L g1994 ( 
.A(n_1937),
.B(n_129),
.Y(n_1994)
);

AOI22xp5_ASAP7_75t_L g1995 ( 
.A1(n_1960),
.A2(n_131),
.B1(n_129),
.B2(n_130),
.Y(n_1995)
);

NAND2xp5_ASAP7_75t_L g1996 ( 
.A(n_1940),
.B(n_130),
.Y(n_1996)
);

BUFx2_ASAP7_75t_L g1997 ( 
.A(n_1908),
.Y(n_1997)
);

INVx2_ASAP7_75t_L g1998 ( 
.A(n_1928),
.Y(n_1998)
);

INVx1_ASAP7_75t_SL g1999 ( 
.A(n_1925),
.Y(n_1999)
);

AND2x4_ASAP7_75t_L g2000 ( 
.A(n_1956),
.B(n_1934),
.Y(n_2000)
);

AO221x2_ASAP7_75t_L g2001 ( 
.A1(n_1961),
.A2(n_1958),
.B1(n_1955),
.B2(n_1933),
.C(n_1968),
.Y(n_2001)
);

NAND2xp5_ASAP7_75t_L g2002 ( 
.A(n_1913),
.B(n_131),
.Y(n_2002)
);

INVx4_ASAP7_75t_L g2003 ( 
.A(n_1905),
.Y(n_2003)
);

NAND2xp5_ASAP7_75t_L g2004 ( 
.A(n_1897),
.B(n_132),
.Y(n_2004)
);

OR2x2_ASAP7_75t_L g2005 ( 
.A(n_1941),
.B(n_132),
.Y(n_2005)
);

NAND2xp5_ASAP7_75t_L g2006 ( 
.A(n_1923),
.B(n_134),
.Y(n_2006)
);

NAND2xp5_ASAP7_75t_L g2007 ( 
.A(n_1936),
.B(n_134),
.Y(n_2007)
);

NOR2xp33_ASAP7_75t_L g2008 ( 
.A(n_1951),
.B(n_135),
.Y(n_2008)
);

AND2x2_ASAP7_75t_L g2009 ( 
.A(n_1931),
.B(n_135),
.Y(n_2009)
);

INVx1_ASAP7_75t_L g2010 ( 
.A(n_1910),
.Y(n_2010)
);

NAND2xp5_ASAP7_75t_L g2011 ( 
.A(n_1914),
.B(n_136),
.Y(n_2011)
);

NAND2xp5_ASAP7_75t_L g2012 ( 
.A(n_1916),
.B(n_136),
.Y(n_2012)
);

AO221x2_ASAP7_75t_L g2013 ( 
.A1(n_1939),
.A2(n_139),
.B1(n_137),
.B2(n_138),
.C(n_140),
.Y(n_2013)
);

BUFx12f_ASAP7_75t_L g2014 ( 
.A(n_1954),
.Y(n_2014)
);

OAI22xp33_ASAP7_75t_L g2015 ( 
.A1(n_1944),
.A2(n_139),
.B1(n_137),
.B2(n_138),
.Y(n_2015)
);

NAND2xp33_ASAP7_75t_R g2016 ( 
.A(n_1957),
.B(n_140),
.Y(n_2016)
);

INVx2_ASAP7_75t_L g2017 ( 
.A(n_1917),
.Y(n_2017)
);

NAND2xp5_ASAP7_75t_L g2018 ( 
.A(n_1919),
.B(n_141),
.Y(n_2018)
);

AOI22xp5_ASAP7_75t_L g2019 ( 
.A1(n_1963),
.A2(n_145),
.B1(n_142),
.B2(n_144),
.Y(n_2019)
);

INVx1_ASAP7_75t_SL g2020 ( 
.A(n_1938),
.Y(n_2020)
);

NAND2xp33_ASAP7_75t_SL g2021 ( 
.A(n_1983),
.B(n_142),
.Y(n_2021)
);

NAND2xp5_ASAP7_75t_L g2022 ( 
.A(n_1922),
.B(n_144),
.Y(n_2022)
);

NAND2xp5_ASAP7_75t_L g2023 ( 
.A(n_1976),
.B(n_145),
.Y(n_2023)
);

OR2x2_ASAP7_75t_L g2024 ( 
.A(n_1977),
.B(n_146),
.Y(n_2024)
);

NAND2xp33_ASAP7_75t_R g2025 ( 
.A(n_1905),
.B(n_146),
.Y(n_2025)
);

INVxp33_ASAP7_75t_SL g2026 ( 
.A(n_1896),
.Y(n_2026)
);

OAI22xp33_ASAP7_75t_L g2027 ( 
.A1(n_1926),
.A2(n_149),
.B1(n_147),
.B2(n_148),
.Y(n_2027)
);

NAND2xp5_ASAP7_75t_L g2028 ( 
.A(n_1979),
.B(n_147),
.Y(n_2028)
);

AO221x2_ASAP7_75t_L g2029 ( 
.A1(n_1932),
.A2(n_150),
.B1(n_148),
.B2(n_149),
.C(n_151),
.Y(n_2029)
);

OAI22xp33_ASAP7_75t_L g2030 ( 
.A1(n_1906),
.A2(n_152),
.B1(n_150),
.B2(n_151),
.Y(n_2030)
);

OAI22xp33_ASAP7_75t_L g2031 ( 
.A1(n_1902),
.A2(n_154),
.B1(n_152),
.B2(n_153),
.Y(n_2031)
);

NOR2x1_ASAP7_75t_L g2032 ( 
.A(n_1969),
.B(n_153),
.Y(n_2032)
);

NOR2x1_ASAP7_75t_L g2033 ( 
.A(n_1911),
.B(n_154),
.Y(n_2033)
);

INVxp67_ASAP7_75t_L g2034 ( 
.A(n_1942),
.Y(n_2034)
);

NOR2x1_ASAP7_75t_SL g2035 ( 
.A(n_1982),
.B(n_155),
.Y(n_2035)
);

NAND2xp5_ASAP7_75t_L g2036 ( 
.A(n_1927),
.B(n_156),
.Y(n_2036)
);

NAND2xp5_ASAP7_75t_L g2037 ( 
.A(n_1921),
.B(n_157),
.Y(n_2037)
);

OAI221xp5_ASAP7_75t_L g2038 ( 
.A1(n_1903),
.A2(n_159),
.B1(n_157),
.B2(n_158),
.C(n_160),
.Y(n_2038)
);

OAI22xp33_ASAP7_75t_L g2039 ( 
.A1(n_1966),
.A2(n_161),
.B1(n_158),
.B2(n_160),
.Y(n_2039)
);

AO221x2_ASAP7_75t_L g2040 ( 
.A1(n_1949),
.A2(n_163),
.B1(n_161),
.B2(n_162),
.C(n_164),
.Y(n_2040)
);

AO221x2_ASAP7_75t_L g2041 ( 
.A1(n_1950),
.A2(n_164),
.B1(n_162),
.B2(n_163),
.C(n_165),
.Y(n_2041)
);

NOR2xp33_ASAP7_75t_L g2042 ( 
.A(n_1898),
.B(n_166),
.Y(n_2042)
);

NAND2xp5_ASAP7_75t_L g2043 ( 
.A(n_1924),
.B(n_166),
.Y(n_2043)
);

INVxp67_ASAP7_75t_L g2044 ( 
.A(n_1930),
.Y(n_2044)
);

CKINVDCx5p33_ASAP7_75t_R g2045 ( 
.A(n_1929),
.Y(n_2045)
);

NAND2xp5_ASAP7_75t_L g2046 ( 
.A(n_1930),
.B(n_167),
.Y(n_2046)
);

NOR4xp25_ASAP7_75t_SL g2047 ( 
.A(n_1985),
.B(n_170),
.C(n_168),
.D(n_169),
.Y(n_2047)
);

INVx1_ASAP7_75t_SL g2048 ( 
.A(n_1918),
.Y(n_2048)
);

OAI221xp5_ASAP7_75t_L g2049 ( 
.A1(n_1964),
.A2(n_170),
.B1(n_168),
.B2(n_169),
.C(n_171),
.Y(n_2049)
);

INVx4_ASAP7_75t_L g2050 ( 
.A(n_1899),
.Y(n_2050)
);

INVxp67_ASAP7_75t_SL g2051 ( 
.A(n_1972),
.Y(n_2051)
);

OAI22xp5_ASAP7_75t_SL g2052 ( 
.A1(n_1948),
.A2(n_173),
.B1(n_171),
.B2(n_172),
.Y(n_2052)
);

NOR2xp33_ASAP7_75t_SL g2053 ( 
.A(n_1934),
.B(n_172),
.Y(n_2053)
);

NOR2xp33_ASAP7_75t_L g2054 ( 
.A(n_1975),
.B(n_173),
.Y(n_2054)
);

AOI22xp5_ASAP7_75t_L g2055 ( 
.A1(n_1959),
.A2(n_176),
.B1(n_174),
.B2(n_175),
.Y(n_2055)
);

NAND2xp5_ASAP7_75t_L g2056 ( 
.A(n_1920),
.B(n_175),
.Y(n_2056)
);

A2O1A1Ixp33_ASAP7_75t_L g2057 ( 
.A1(n_1915),
.A2(n_179),
.B(n_176),
.C(n_178),
.Y(n_2057)
);

CKINVDCx5p33_ASAP7_75t_R g2058 ( 
.A(n_1900),
.Y(n_2058)
);

AOI22xp5_ASAP7_75t_L g2059 ( 
.A1(n_1970),
.A2(n_181),
.B1(n_179),
.B2(n_180),
.Y(n_2059)
);

NOR2xp33_ASAP7_75t_R g2060 ( 
.A(n_1952),
.B(n_1953),
.Y(n_2060)
);

AO221x2_ASAP7_75t_L g2061 ( 
.A1(n_1978),
.A2(n_182),
.B1(n_180),
.B2(n_181),
.C(n_183),
.Y(n_2061)
);

NAND2xp5_ASAP7_75t_L g2062 ( 
.A(n_1984),
.B(n_184),
.Y(n_2062)
);

OAI22xp33_ASAP7_75t_L g2063 ( 
.A1(n_1947),
.A2(n_186),
.B1(n_184),
.B2(n_185),
.Y(n_2063)
);

AND2x2_ASAP7_75t_L g2064 ( 
.A(n_1971),
.B(n_186),
.Y(n_2064)
);

AO221x2_ASAP7_75t_L g2065 ( 
.A1(n_1943),
.A2(n_190),
.B1(n_187),
.B2(n_188),
.C(n_191),
.Y(n_2065)
);

NAND2xp5_ASAP7_75t_L g2066 ( 
.A(n_1904),
.B(n_1973),
.Y(n_2066)
);

INVxp67_ASAP7_75t_L g2067 ( 
.A(n_1974),
.Y(n_2067)
);

NAND2xp5_ASAP7_75t_L g2068 ( 
.A(n_1981),
.B(n_187),
.Y(n_2068)
);

NAND2xp5_ASAP7_75t_L g2069 ( 
.A(n_1945),
.B(n_188),
.Y(n_2069)
);

INVxp67_ASAP7_75t_L g2070 ( 
.A(n_1942),
.Y(n_2070)
);

CKINVDCx20_ASAP7_75t_R g2071 ( 
.A(n_1980),
.Y(n_2071)
);

INVx2_ASAP7_75t_SL g2072 ( 
.A(n_1925),
.Y(n_2072)
);

OR2x2_ASAP7_75t_L g2073 ( 
.A(n_1909),
.B(n_190),
.Y(n_2073)
);

OAI22xp33_ASAP7_75t_L g2074 ( 
.A1(n_1965),
.A2(n_193),
.B1(n_191),
.B2(n_192),
.Y(n_2074)
);

NOR4xp25_ASAP7_75t_SL g2075 ( 
.A(n_1962),
.B(n_194),
.C(n_192),
.D(n_193),
.Y(n_2075)
);

NOR2xp33_ASAP7_75t_L g2076 ( 
.A(n_1913),
.B(n_194),
.Y(n_2076)
);

INVx1_ASAP7_75t_L g2077 ( 
.A(n_1910),
.Y(n_2077)
);

NAND2xp5_ASAP7_75t_L g2078 ( 
.A(n_1946),
.B(n_195),
.Y(n_2078)
);

INVx2_ASAP7_75t_L g2079 ( 
.A(n_1928),
.Y(n_2079)
);

NAND2xp5_ASAP7_75t_L g2080 ( 
.A(n_1946),
.B(n_195),
.Y(n_2080)
);

INVx2_ASAP7_75t_SL g2081 ( 
.A(n_1925),
.Y(n_2081)
);

CKINVDCx5p33_ASAP7_75t_R g2082 ( 
.A(n_1980),
.Y(n_2082)
);

NOR4xp25_ASAP7_75t_SL g2083 ( 
.A(n_1962),
.B(n_198),
.C(n_196),
.D(n_197),
.Y(n_2083)
);

AOI22xp5_ASAP7_75t_L g2084 ( 
.A1(n_1965),
.A2(n_198),
.B1(n_196),
.B2(n_197),
.Y(n_2084)
);

OAI22xp33_ASAP7_75t_L g2085 ( 
.A1(n_1965),
.A2(n_201),
.B1(n_199),
.B2(n_200),
.Y(n_2085)
);

NAND2xp5_ASAP7_75t_L g2086 ( 
.A(n_1946),
.B(n_199),
.Y(n_2086)
);

OAI22xp33_ASAP7_75t_L g2087 ( 
.A1(n_1965),
.A2(n_202),
.B1(n_200),
.B2(n_201),
.Y(n_2087)
);

NOR2x1_ASAP7_75t_L g2088 ( 
.A(n_1896),
.B(n_202),
.Y(n_2088)
);

AOI22xp5_ASAP7_75t_L g2089 ( 
.A1(n_1965),
.A2(n_205),
.B1(n_203),
.B2(n_204),
.Y(n_2089)
);

AO221x2_ASAP7_75t_L g2090 ( 
.A1(n_1962),
.A2(n_206),
.B1(n_203),
.B2(n_205),
.C(n_207),
.Y(n_2090)
);

CKINVDCx20_ASAP7_75t_R g2091 ( 
.A(n_1980),
.Y(n_2091)
);

INVx1_ASAP7_75t_SL g2092 ( 
.A(n_1935),
.Y(n_2092)
);

INVx1_ASAP7_75t_L g2093 ( 
.A(n_2010),
.Y(n_2093)
);

NAND2xp33_ASAP7_75t_SL g2094 ( 
.A(n_2025),
.B(n_2016),
.Y(n_2094)
);

INVx1_ASAP7_75t_L g2095 ( 
.A(n_2077),
.Y(n_2095)
);

AND2x2_ASAP7_75t_L g2096 ( 
.A(n_1997),
.B(n_206),
.Y(n_2096)
);

AND2x4_ASAP7_75t_L g2097 ( 
.A(n_2044),
.B(n_207),
.Y(n_2097)
);

NOR2x1_ASAP7_75t_L g2098 ( 
.A(n_2088),
.B(n_208),
.Y(n_2098)
);

AOI22xp33_ASAP7_75t_L g2099 ( 
.A1(n_1990),
.A2(n_212),
.B1(n_209),
.B2(n_210),
.Y(n_2099)
);

INVx2_ASAP7_75t_L g2100 ( 
.A(n_1989),
.Y(n_2100)
);

NOR2xp33_ASAP7_75t_L g2101 ( 
.A(n_2026),
.B(n_209),
.Y(n_2101)
);

HB1xp67_ASAP7_75t_L g2102 ( 
.A(n_2017),
.Y(n_2102)
);

BUFx2_ASAP7_75t_L g2103 ( 
.A(n_2034),
.Y(n_2103)
);

NAND2xp5_ASAP7_75t_L g2104 ( 
.A(n_2001),
.B(n_212),
.Y(n_2104)
);

INVx2_ASAP7_75t_L g2105 ( 
.A(n_1992),
.Y(n_2105)
);

INVx2_ASAP7_75t_L g2106 ( 
.A(n_1998),
.Y(n_2106)
);

AOI22xp33_ASAP7_75t_L g2107 ( 
.A1(n_2001),
.A2(n_215),
.B1(n_213),
.B2(n_214),
.Y(n_2107)
);

AOI22xp5_ASAP7_75t_L g2108 ( 
.A1(n_2090),
.A2(n_2040),
.B1(n_2041),
.B2(n_2013),
.Y(n_2108)
);

HB1xp67_ASAP7_75t_L g2109 ( 
.A(n_2070),
.Y(n_2109)
);

INVx1_ASAP7_75t_SL g2110 ( 
.A(n_1999),
.Y(n_2110)
);

NOR2xp33_ASAP7_75t_L g2111 ( 
.A(n_1988),
.B(n_213),
.Y(n_2111)
);

AND2x4_ASAP7_75t_L g2112 ( 
.A(n_2003),
.B(n_216),
.Y(n_2112)
);

HB1xp67_ASAP7_75t_L g2113 ( 
.A(n_2020),
.Y(n_2113)
);

INVx1_ASAP7_75t_L g2114 ( 
.A(n_2006),
.Y(n_2114)
);

NAND2x1_ASAP7_75t_L g2115 ( 
.A(n_2072),
.B(n_217),
.Y(n_2115)
);

AND2x2_ASAP7_75t_L g2116 ( 
.A(n_2000),
.B(n_217),
.Y(n_2116)
);

INVx1_ASAP7_75t_L g2117 ( 
.A(n_2024),
.Y(n_2117)
);

INVx1_ASAP7_75t_L g2118 ( 
.A(n_2004),
.Y(n_2118)
);

INVx3_ASAP7_75t_L g2119 ( 
.A(n_2081),
.Y(n_2119)
);

OR2x2_ASAP7_75t_L g2120 ( 
.A(n_2073),
.B(n_218),
.Y(n_2120)
);

INVx1_ASAP7_75t_L g2121 ( 
.A(n_2005),
.Y(n_2121)
);

INVx1_ASAP7_75t_SL g2122 ( 
.A(n_2092),
.Y(n_2122)
);

AND2x2_ASAP7_75t_L g2123 ( 
.A(n_2048),
.B(n_219),
.Y(n_2123)
);

INVx1_ASAP7_75t_L g2124 ( 
.A(n_2011),
.Y(n_2124)
);

INVx1_ASAP7_75t_L g2125 ( 
.A(n_2012),
.Y(n_2125)
);

INVx1_ASAP7_75t_L g2126 ( 
.A(n_2018),
.Y(n_2126)
);

INVx1_ASAP7_75t_L g2127 ( 
.A(n_2022),
.Y(n_2127)
);

NAND2xp5_ASAP7_75t_L g2128 ( 
.A(n_2067),
.B(n_219),
.Y(n_2128)
);

INVx4_ASAP7_75t_L g2129 ( 
.A(n_2082),
.Y(n_2129)
);

OR2x2_ASAP7_75t_L g2130 ( 
.A(n_2079),
.B(n_220),
.Y(n_2130)
);

INVx1_ASAP7_75t_L g2131 ( 
.A(n_2023),
.Y(n_2131)
);

NAND2xp5_ASAP7_75t_L g2132 ( 
.A(n_2028),
.B(n_220),
.Y(n_2132)
);

BUFx3_ASAP7_75t_L g2133 ( 
.A(n_2071),
.Y(n_2133)
);

AOI21xp5_ASAP7_75t_L g2134 ( 
.A1(n_2021),
.A2(n_221),
.B(n_222),
.Y(n_2134)
);

INVx2_ASAP7_75t_L g2135 ( 
.A(n_2035),
.Y(n_2135)
);

INVx1_ASAP7_75t_L g2136 ( 
.A(n_1986),
.Y(n_2136)
);

AND2x2_ASAP7_75t_L g2137 ( 
.A(n_2009),
.B(n_221),
.Y(n_2137)
);

NAND2xp5_ASAP7_75t_SL g2138 ( 
.A(n_1993),
.B(n_222),
.Y(n_2138)
);

INVx1_ASAP7_75t_SL g2139 ( 
.A(n_2091),
.Y(n_2139)
);

OR2x2_ASAP7_75t_L g2140 ( 
.A(n_1994),
.B(n_1996),
.Y(n_2140)
);

INVxp67_ASAP7_75t_SL g2141 ( 
.A(n_2032),
.Y(n_2141)
);

INVx2_ASAP7_75t_L g2142 ( 
.A(n_2050),
.Y(n_2142)
);

AOI22xp33_ASAP7_75t_L g2143 ( 
.A1(n_2090),
.A2(n_225),
.B1(n_223),
.B2(n_224),
.Y(n_2143)
);

OR2x2_ASAP7_75t_L g2144 ( 
.A(n_2078),
.B(n_2080),
.Y(n_2144)
);

INVx1_ASAP7_75t_SL g2145 ( 
.A(n_2060),
.Y(n_2145)
);

NAND2xp5_ASAP7_75t_L g2146 ( 
.A(n_2086),
.B(n_223),
.Y(n_2146)
);

OR2x2_ASAP7_75t_L g2147 ( 
.A(n_2066),
.B(n_224),
.Y(n_2147)
);

CKINVDCx16_ASAP7_75t_R g2148 ( 
.A(n_2053),
.Y(n_2148)
);

NAND2xp5_ASAP7_75t_L g2149 ( 
.A(n_2076),
.B(n_225),
.Y(n_2149)
);

AND2x2_ASAP7_75t_L g2150 ( 
.A(n_2014),
.B(n_226),
.Y(n_2150)
);

AOI22xp33_ASAP7_75t_L g2151 ( 
.A1(n_2040),
.A2(n_228),
.B1(n_226),
.B2(n_227),
.Y(n_2151)
);

INVx1_ASAP7_75t_L g2152 ( 
.A(n_2002),
.Y(n_2152)
);

NAND3xp33_ASAP7_75t_L g2153 ( 
.A(n_2084),
.B(n_227),
.C(n_228),
.Y(n_2153)
);

INVx2_ASAP7_75t_L g2154 ( 
.A(n_2046),
.Y(n_2154)
);

NAND2xp5_ASAP7_75t_L g2155 ( 
.A(n_2033),
.B(n_229),
.Y(n_2155)
);

INVx1_ASAP7_75t_L g2156 ( 
.A(n_1991),
.Y(n_2156)
);

HB1xp67_ASAP7_75t_L g2157 ( 
.A(n_2058),
.Y(n_2157)
);

INVx1_ASAP7_75t_SL g2158 ( 
.A(n_2045),
.Y(n_2158)
);

INVxp67_ASAP7_75t_L g2159 ( 
.A(n_2008),
.Y(n_2159)
);

INVx1_ASAP7_75t_L g2160 ( 
.A(n_2036),
.Y(n_2160)
);

AND2x2_ASAP7_75t_L g2161 ( 
.A(n_2064),
.B(n_229),
.Y(n_2161)
);

OR2x2_ASAP7_75t_L g2162 ( 
.A(n_2007),
.B(n_230),
.Y(n_2162)
);

INVxp67_ASAP7_75t_L g2163 ( 
.A(n_2042),
.Y(n_2163)
);

INVx1_ASAP7_75t_SL g2164 ( 
.A(n_2037),
.Y(n_2164)
);

INVx1_ASAP7_75t_L g2165 ( 
.A(n_2062),
.Y(n_2165)
);

INVx1_ASAP7_75t_SL g2166 ( 
.A(n_2043),
.Y(n_2166)
);

INVx2_ASAP7_75t_SL g2167 ( 
.A(n_2065),
.Y(n_2167)
);

AND2x4_ASAP7_75t_L g2168 ( 
.A(n_2056),
.B(n_230),
.Y(n_2168)
);

HB1xp67_ASAP7_75t_L g2169 ( 
.A(n_2061),
.Y(n_2169)
);

INVx1_ASAP7_75t_SL g2170 ( 
.A(n_2068),
.Y(n_2170)
);

AND2x2_ASAP7_75t_L g2171 ( 
.A(n_2069),
.B(n_231),
.Y(n_2171)
);

INVx2_ASAP7_75t_SL g2172 ( 
.A(n_2065),
.Y(n_2172)
);

NAND2xp5_ASAP7_75t_L g2173 ( 
.A(n_2054),
.B(n_231),
.Y(n_2173)
);

INVx2_ASAP7_75t_L g2174 ( 
.A(n_2013),
.Y(n_2174)
);

AND2x2_ASAP7_75t_L g2175 ( 
.A(n_2029),
.B(n_232),
.Y(n_2175)
);

AND2x2_ASAP7_75t_L g2176 ( 
.A(n_2029),
.B(n_232),
.Y(n_2176)
);

NAND3xp33_ASAP7_75t_SL g2177 ( 
.A(n_2089),
.B(n_233),
.C(n_234),
.Y(n_2177)
);

BUFx2_ASAP7_75t_L g2178 ( 
.A(n_2019),
.Y(n_2178)
);

INVx1_ASAP7_75t_L g2179 ( 
.A(n_2061),
.Y(n_2179)
);

OAI22xp5_ASAP7_75t_L g2180 ( 
.A1(n_2049),
.A2(n_235),
.B1(n_233),
.B2(n_234),
.Y(n_2180)
);

AND2x2_ASAP7_75t_L g2181 ( 
.A(n_2041),
.B(n_236),
.Y(n_2181)
);

AND2x2_ASAP7_75t_L g2182 ( 
.A(n_2059),
.B(n_236),
.Y(n_2182)
);

AOI22xp33_ASAP7_75t_L g2183 ( 
.A1(n_1987),
.A2(n_239),
.B1(n_237),
.B2(n_238),
.Y(n_2183)
);

NAND2xp5_ASAP7_75t_L g2184 ( 
.A(n_2027),
.B(n_237),
.Y(n_2184)
);

INVx2_ASAP7_75t_L g2185 ( 
.A(n_2052),
.Y(n_2185)
);

INVx1_ASAP7_75t_L g2186 ( 
.A(n_2030),
.Y(n_2186)
);

INVx1_ASAP7_75t_L g2187 ( 
.A(n_2031),
.Y(n_2187)
);

AO21x2_ASAP7_75t_L g2188 ( 
.A1(n_2074),
.A2(n_238),
.B(n_239),
.Y(n_2188)
);

AND2x2_ASAP7_75t_L g2189 ( 
.A(n_2055),
.B(n_240),
.Y(n_2189)
);

INVx1_ASAP7_75t_SL g2190 ( 
.A(n_1995),
.Y(n_2190)
);

INVx1_ASAP7_75t_SL g2191 ( 
.A(n_2063),
.Y(n_2191)
);

INVx1_ASAP7_75t_L g2192 ( 
.A(n_2015),
.Y(n_2192)
);

OAI22xp5_ASAP7_75t_L g2193 ( 
.A1(n_2038),
.A2(n_2057),
.B1(n_2083),
.B2(n_2075),
.Y(n_2193)
);

INVx2_ASAP7_75t_L g2194 ( 
.A(n_2047),
.Y(n_2194)
);

AOI22xp5_ASAP7_75t_L g2195 ( 
.A1(n_2085),
.A2(n_243),
.B1(n_240),
.B2(n_242),
.Y(n_2195)
);

AND2x2_ASAP7_75t_L g2196 ( 
.A(n_2039),
.B(n_242),
.Y(n_2196)
);

NOR2xp33_ASAP7_75t_L g2197 ( 
.A(n_2087),
.B(n_243),
.Y(n_2197)
);

AND2x2_ASAP7_75t_L g2198 ( 
.A(n_1997),
.B(n_244),
.Y(n_2198)
);

OR2x2_ASAP7_75t_L g2199 ( 
.A(n_1992),
.B(n_244),
.Y(n_2199)
);

INVx1_ASAP7_75t_L g2200 ( 
.A(n_2010),
.Y(n_2200)
);

INVx1_ASAP7_75t_L g2201 ( 
.A(n_2010),
.Y(n_2201)
);

AND2x2_ASAP7_75t_L g2202 ( 
.A(n_1997),
.B(n_245),
.Y(n_2202)
);

AND2x4_ASAP7_75t_L g2203 ( 
.A(n_2003),
.B(n_245),
.Y(n_2203)
);

NOR2xp33_ASAP7_75t_L g2204 ( 
.A(n_2026),
.B(n_246),
.Y(n_2204)
);

INVx1_ASAP7_75t_L g2205 ( 
.A(n_2010),
.Y(n_2205)
);

INVx1_ASAP7_75t_L g2206 ( 
.A(n_2010),
.Y(n_2206)
);

INVx1_ASAP7_75t_L g2207 ( 
.A(n_2010),
.Y(n_2207)
);

AND3x1_ASAP7_75t_L g2208 ( 
.A(n_2053),
.B(n_246),
.C(n_247),
.Y(n_2208)
);

INVx2_ASAP7_75t_L g2209 ( 
.A(n_1997),
.Y(n_2209)
);

AND3x2_ASAP7_75t_L g2210 ( 
.A(n_2034),
.B(n_248),
.C(n_249),
.Y(n_2210)
);

INVx3_ASAP7_75t_L g2211 ( 
.A(n_2003),
.Y(n_2211)
);

AND2x2_ASAP7_75t_L g2212 ( 
.A(n_1997),
.B(n_250),
.Y(n_2212)
);

AOI22xp33_ASAP7_75t_SL g2213 ( 
.A1(n_2026),
.A2(n_252),
.B1(n_250),
.B2(n_251),
.Y(n_2213)
);

NOR2xp33_ASAP7_75t_L g2214 ( 
.A(n_2026),
.B(n_252),
.Y(n_2214)
);

AND2x2_ASAP7_75t_L g2215 ( 
.A(n_1997),
.B(n_253),
.Y(n_2215)
);

INVx1_ASAP7_75t_L g2216 ( 
.A(n_2010),
.Y(n_2216)
);

NAND2xp5_ASAP7_75t_L g2217 ( 
.A(n_2051),
.B(n_254),
.Y(n_2217)
);

INVx1_ASAP7_75t_L g2218 ( 
.A(n_2010),
.Y(n_2218)
);

NAND2xp5_ASAP7_75t_L g2219 ( 
.A(n_2051),
.B(n_254),
.Y(n_2219)
);

INVx1_ASAP7_75t_L g2220 ( 
.A(n_2010),
.Y(n_2220)
);

INVx1_ASAP7_75t_L g2221 ( 
.A(n_2010),
.Y(n_2221)
);

AND2x4_ASAP7_75t_L g2222 ( 
.A(n_2044),
.B(n_255),
.Y(n_2222)
);

INVx3_ASAP7_75t_L g2223 ( 
.A(n_2003),
.Y(n_2223)
);

AND2x2_ASAP7_75t_L g2224 ( 
.A(n_1997),
.B(n_255),
.Y(n_2224)
);

AND2x2_ASAP7_75t_L g2225 ( 
.A(n_1997),
.B(n_256),
.Y(n_2225)
);

HB1xp67_ASAP7_75t_L g2226 ( 
.A(n_1997),
.Y(n_2226)
);

AND2x4_ASAP7_75t_L g2227 ( 
.A(n_2044),
.B(n_256),
.Y(n_2227)
);

INVx1_ASAP7_75t_SL g2228 ( 
.A(n_2026),
.Y(n_2228)
);

INVx1_ASAP7_75t_L g2229 ( 
.A(n_2010),
.Y(n_2229)
);

INVx1_ASAP7_75t_L g2230 ( 
.A(n_2010),
.Y(n_2230)
);

HB1xp67_ASAP7_75t_L g2231 ( 
.A(n_1997),
.Y(n_2231)
);

INVx2_ASAP7_75t_SL g2232 ( 
.A(n_1997),
.Y(n_2232)
);

OR2x2_ASAP7_75t_L g2233 ( 
.A(n_1992),
.B(n_257),
.Y(n_2233)
);

INVx2_ASAP7_75t_L g2234 ( 
.A(n_1997),
.Y(n_2234)
);

NOR2xp33_ASAP7_75t_L g2235 ( 
.A(n_2026),
.B(n_258),
.Y(n_2235)
);

OR2x2_ASAP7_75t_L g2236 ( 
.A(n_1992),
.B(n_258),
.Y(n_2236)
);

INVx2_ASAP7_75t_SL g2237 ( 
.A(n_1997),
.Y(n_2237)
);

NAND2xp5_ASAP7_75t_L g2238 ( 
.A(n_2051),
.B(n_259),
.Y(n_2238)
);

OAI22xp5_ASAP7_75t_L g2239 ( 
.A1(n_2026),
.A2(n_261),
.B1(n_259),
.B2(n_260),
.Y(n_2239)
);

AND2x2_ASAP7_75t_L g2240 ( 
.A(n_1997),
.B(n_262),
.Y(n_2240)
);

INVx1_ASAP7_75t_SL g2241 ( 
.A(n_2026),
.Y(n_2241)
);

AOI221xp5_ASAP7_75t_L g2242 ( 
.A1(n_2074),
.A2(n_264),
.B1(n_262),
.B2(n_263),
.C(n_265),
.Y(n_2242)
);

AND2x2_ASAP7_75t_L g2243 ( 
.A(n_1997),
.B(n_263),
.Y(n_2243)
);

INVxp67_ASAP7_75t_SL g2244 ( 
.A(n_2034),
.Y(n_2244)
);

AOI22xp33_ASAP7_75t_L g2245 ( 
.A1(n_1990),
.A2(n_266),
.B1(n_264),
.B2(n_265),
.Y(n_2245)
);

OAI22xp33_ASAP7_75t_L g2246 ( 
.A1(n_2108),
.A2(n_269),
.B1(n_267),
.B2(n_268),
.Y(n_2246)
);

INVx1_ASAP7_75t_L g2247 ( 
.A(n_2093),
.Y(n_2247)
);

NAND2xp5_ASAP7_75t_L g2248 ( 
.A(n_2141),
.B(n_2244),
.Y(n_2248)
);

OAI22xp33_ASAP7_75t_L g2249 ( 
.A1(n_2169),
.A2(n_270),
.B1(n_268),
.B2(n_269),
.Y(n_2249)
);

OAI22xp5_ASAP7_75t_L g2250 ( 
.A1(n_2107),
.A2(n_272),
.B1(n_270),
.B2(n_271),
.Y(n_2250)
);

NAND2xp5_ASAP7_75t_L g2251 ( 
.A(n_2109),
.B(n_271),
.Y(n_2251)
);

AOI21xp5_ASAP7_75t_L g2252 ( 
.A1(n_2094),
.A2(n_272),
.B(n_273),
.Y(n_2252)
);

O2A1O1Ixp33_ASAP7_75t_SL g2253 ( 
.A1(n_2167),
.A2(n_276),
.B(n_273),
.C(n_275),
.Y(n_2253)
);

NAND4xp25_ASAP7_75t_L g2254 ( 
.A(n_2151),
.B(n_277),
.C(n_275),
.D(n_276),
.Y(n_2254)
);

INVx1_ASAP7_75t_SL g2255 ( 
.A(n_2228),
.Y(n_2255)
);

CKINVDCx14_ASAP7_75t_R g2256 ( 
.A(n_2175),
.Y(n_2256)
);

OAI21xp5_ASAP7_75t_L g2257 ( 
.A1(n_2098),
.A2(n_277),
.B(n_278),
.Y(n_2257)
);

OAI31xp33_ASAP7_75t_L g2258 ( 
.A1(n_2193),
.A2(n_280),
.A3(n_278),
.B(n_279),
.Y(n_2258)
);

INVx1_ASAP7_75t_L g2259 ( 
.A(n_2095),
.Y(n_2259)
);

OAI21xp5_ASAP7_75t_L g2260 ( 
.A1(n_2104),
.A2(n_279),
.B(n_280),
.Y(n_2260)
);

A2O1A1Ixp33_ASAP7_75t_L g2261 ( 
.A1(n_2172),
.A2(n_283),
.B(n_281),
.C(n_282),
.Y(n_2261)
);

NAND2x1p5_ASAP7_75t_L g2262 ( 
.A(n_2122),
.B(n_281),
.Y(n_2262)
);

OAI21xp33_ASAP7_75t_L g2263 ( 
.A1(n_2143),
.A2(n_282),
.B(n_283),
.Y(n_2263)
);

NAND2xp5_ASAP7_75t_L g2264 ( 
.A(n_2103),
.B(n_284),
.Y(n_2264)
);

NOR2xp33_ASAP7_75t_L g2265 ( 
.A(n_2241),
.B(n_285),
.Y(n_2265)
);

INVx1_ASAP7_75t_L g2266 ( 
.A(n_2200),
.Y(n_2266)
);

AOI221xp5_ASAP7_75t_L g2267 ( 
.A1(n_2178),
.A2(n_288),
.B1(n_286),
.B2(n_287),
.C(n_289),
.Y(n_2267)
);

OR4x1_ASAP7_75t_L g2268 ( 
.A(n_2232),
.B(n_289),
.C(n_286),
.D(n_287),
.Y(n_2268)
);

INVx1_ASAP7_75t_L g2269 ( 
.A(n_2201),
.Y(n_2269)
);

INVx1_ASAP7_75t_L g2270 ( 
.A(n_2205),
.Y(n_2270)
);

AOI21xp33_ASAP7_75t_L g2271 ( 
.A1(n_2184),
.A2(n_2145),
.B(n_2190),
.Y(n_2271)
);

INVx1_ASAP7_75t_L g2272 ( 
.A(n_2206),
.Y(n_2272)
);

OR2x2_ASAP7_75t_L g2273 ( 
.A(n_2105),
.B(n_290),
.Y(n_2273)
);

NAND2xp5_ASAP7_75t_L g2274 ( 
.A(n_2113),
.B(n_290),
.Y(n_2274)
);

O2A1O1Ixp33_ASAP7_75t_L g2275 ( 
.A1(n_2179),
.A2(n_293),
.B(n_291),
.C(n_292),
.Y(n_2275)
);

INVx2_ASAP7_75t_L g2276 ( 
.A(n_2211),
.Y(n_2276)
);

OAI21xp5_ASAP7_75t_L g2277 ( 
.A1(n_2153),
.A2(n_291),
.B(n_294),
.Y(n_2277)
);

NAND2xp5_ASAP7_75t_SL g2278 ( 
.A(n_2148),
.B(n_294),
.Y(n_2278)
);

INVx1_ASAP7_75t_L g2279 ( 
.A(n_2207),
.Y(n_2279)
);

AND2x2_ASAP7_75t_L g2280 ( 
.A(n_2223),
.B(n_295),
.Y(n_2280)
);

INVx1_ASAP7_75t_L g2281 ( 
.A(n_2216),
.Y(n_2281)
);

OAI21xp5_ASAP7_75t_L g2282 ( 
.A1(n_2134),
.A2(n_295),
.B(n_296),
.Y(n_2282)
);

OAI22xp33_ASAP7_75t_L g2283 ( 
.A1(n_2174),
.A2(n_298),
.B1(n_296),
.B2(n_297),
.Y(n_2283)
);

AOI21xp33_ASAP7_75t_L g2284 ( 
.A1(n_2192),
.A2(n_298),
.B(n_299),
.Y(n_2284)
);

OAI22xp33_ASAP7_75t_L g2285 ( 
.A1(n_2237),
.A2(n_301),
.B1(n_299),
.B2(n_300),
.Y(n_2285)
);

AO22x1_ASAP7_75t_L g2286 ( 
.A1(n_2135),
.A2(n_302),
.B1(n_300),
.B2(n_301),
.Y(n_2286)
);

NAND2x1_ASAP7_75t_SL g2287 ( 
.A(n_2226),
.B(n_302),
.Y(n_2287)
);

INVx1_ASAP7_75t_L g2288 ( 
.A(n_2218),
.Y(n_2288)
);

OAI322xp33_ASAP7_75t_L g2289 ( 
.A1(n_2197),
.A2(n_303),
.A3(n_304),
.B1(n_305),
.B2(n_306),
.C1(n_307),
.C2(n_308),
.Y(n_2289)
);

AOI321xp33_ASAP7_75t_L g2290 ( 
.A1(n_2208),
.A2(n_306),
.A3(n_308),
.B1(n_303),
.B2(n_304),
.C(n_307),
.Y(n_2290)
);

INVx2_ASAP7_75t_L g2291 ( 
.A(n_2119),
.Y(n_2291)
);

NAND2xp5_ASAP7_75t_L g2292 ( 
.A(n_2154),
.B(n_309),
.Y(n_2292)
);

AOI22xp5_ASAP7_75t_L g2293 ( 
.A1(n_2177),
.A2(n_311),
.B1(n_309),
.B2(n_310),
.Y(n_2293)
);

INVx1_ASAP7_75t_L g2294 ( 
.A(n_2220),
.Y(n_2294)
);

AOI222xp33_ASAP7_75t_L g2295 ( 
.A1(n_2181),
.A2(n_312),
.B1(n_314),
.B2(n_310),
.C1(n_311),
.C2(n_313),
.Y(n_2295)
);

INVxp67_ASAP7_75t_L g2296 ( 
.A(n_2231),
.Y(n_2296)
);

INVx1_ASAP7_75t_L g2297 ( 
.A(n_2221),
.Y(n_2297)
);

OA21x2_ASAP7_75t_L g2298 ( 
.A1(n_2209),
.A2(n_313),
.B(n_314),
.Y(n_2298)
);

AOI222xp33_ASAP7_75t_L g2299 ( 
.A1(n_2176),
.A2(n_318),
.B1(n_320),
.B2(n_315),
.C1(n_317),
.C2(n_319),
.Y(n_2299)
);

INVx1_ASAP7_75t_L g2300 ( 
.A(n_2229),
.Y(n_2300)
);

NOR2xp33_ASAP7_75t_L g2301 ( 
.A(n_2170),
.B(n_2164),
.Y(n_2301)
);

AOI22xp33_ASAP7_75t_L g2302 ( 
.A1(n_2186),
.A2(n_2185),
.B1(n_2187),
.B2(n_2191),
.Y(n_2302)
);

NAND2xp5_ASAP7_75t_L g2303 ( 
.A(n_2156),
.B(n_2166),
.Y(n_2303)
);

INVxp67_ASAP7_75t_SL g2304 ( 
.A(n_2157),
.Y(n_2304)
);

AOI211xp5_ASAP7_75t_SL g2305 ( 
.A1(n_2180),
.A2(n_2242),
.B(n_2239),
.C(n_2195),
.Y(n_2305)
);

OAI21xp5_ASAP7_75t_L g2306 ( 
.A1(n_2099),
.A2(n_315),
.B(n_317),
.Y(n_2306)
);

NAND2xp5_ASAP7_75t_L g2307 ( 
.A(n_2117),
.B(n_319),
.Y(n_2307)
);

O2A1O1Ixp5_ASAP7_75t_SL g2308 ( 
.A1(n_2138),
.A2(n_2159),
.B(n_2163),
.C(n_2155),
.Y(n_2308)
);

INVx1_ASAP7_75t_L g2309 ( 
.A(n_2230),
.Y(n_2309)
);

NAND2xp5_ASAP7_75t_L g2310 ( 
.A(n_2160),
.B(n_320),
.Y(n_2310)
);

AOI21xp33_ASAP7_75t_L g2311 ( 
.A1(n_2188),
.A2(n_2194),
.B(n_2144),
.Y(n_2311)
);

OAI21xp33_ASAP7_75t_L g2312 ( 
.A1(n_2183),
.A2(n_321),
.B(n_322),
.Y(n_2312)
);

AOI221xp5_ASAP7_75t_L g2313 ( 
.A1(n_2101),
.A2(n_325),
.B1(n_322),
.B2(n_324),
.C(n_326),
.Y(n_2313)
);

NAND2xp5_ASAP7_75t_L g2314 ( 
.A(n_2165),
.B(n_2121),
.Y(n_2314)
);

OR2x2_ASAP7_75t_L g2315 ( 
.A(n_2234),
.B(n_324),
.Y(n_2315)
);

OAI21xp33_ASAP7_75t_L g2316 ( 
.A1(n_2245),
.A2(n_325),
.B(n_327),
.Y(n_2316)
);

AOI221xp5_ASAP7_75t_L g2317 ( 
.A1(n_2204),
.A2(n_330),
.B1(n_328),
.B2(n_329),
.C(n_331),
.Y(n_2317)
);

INVxp67_ASAP7_75t_L g2318 ( 
.A(n_2097),
.Y(n_2318)
);

AOI22xp5_ASAP7_75t_L g2319 ( 
.A1(n_2110),
.A2(n_331),
.B1(n_329),
.B2(n_330),
.Y(n_2319)
);

INVx1_ASAP7_75t_L g2320 ( 
.A(n_2102),
.Y(n_2320)
);

O2A1O1Ixp33_ASAP7_75t_SL g2321 ( 
.A1(n_2115),
.A2(n_334),
.B(n_332),
.C(n_333),
.Y(n_2321)
);

INVx1_ASAP7_75t_L g2322 ( 
.A(n_2114),
.Y(n_2322)
);

NAND2xp5_ASAP7_75t_L g2323 ( 
.A(n_2136),
.B(n_332),
.Y(n_2323)
);

INVx1_ASAP7_75t_L g2324 ( 
.A(n_2118),
.Y(n_2324)
);

INVx1_ASAP7_75t_L g2325 ( 
.A(n_2124),
.Y(n_2325)
);

NAND2xp5_ASAP7_75t_L g2326 ( 
.A(n_2152),
.B(n_335),
.Y(n_2326)
);

INVx2_ASAP7_75t_L g2327 ( 
.A(n_2142),
.Y(n_2327)
);

INVx1_ASAP7_75t_L g2328 ( 
.A(n_2125),
.Y(n_2328)
);

AO21x1_ASAP7_75t_L g2329 ( 
.A1(n_2214),
.A2(n_336),
.B(n_337),
.Y(n_2329)
);

NOR2xp33_ASAP7_75t_L g2330 ( 
.A(n_2129),
.B(n_2140),
.Y(n_2330)
);

NOR2xp33_ASAP7_75t_L g2331 ( 
.A(n_2158),
.B(n_336),
.Y(n_2331)
);

NOR2xp33_ASAP7_75t_SL g2332 ( 
.A(n_2139),
.B(n_337),
.Y(n_2332)
);

NAND2x1_ASAP7_75t_L g2333 ( 
.A(n_2100),
.B(n_338),
.Y(n_2333)
);

INVx1_ASAP7_75t_L g2334 ( 
.A(n_2126),
.Y(n_2334)
);

NAND2xp5_ASAP7_75t_L g2335 ( 
.A(n_2127),
.B(n_338),
.Y(n_2335)
);

INVx1_ASAP7_75t_L g2336 ( 
.A(n_2131),
.Y(n_2336)
);

NAND2xp5_ASAP7_75t_L g2337 ( 
.A(n_2097),
.B(n_339),
.Y(n_2337)
);

AOI22xp5_ASAP7_75t_L g2338 ( 
.A1(n_2196),
.A2(n_342),
.B1(n_340),
.B2(n_341),
.Y(n_2338)
);

AOI211xp5_ASAP7_75t_L g2339 ( 
.A1(n_2235),
.A2(n_342),
.B(n_340),
.C(n_341),
.Y(n_2339)
);

INVx2_ASAP7_75t_L g2340 ( 
.A(n_2106),
.Y(n_2340)
);

INVx1_ASAP7_75t_L g2341 ( 
.A(n_2130),
.Y(n_2341)
);

NAND2xp5_ASAP7_75t_L g2342 ( 
.A(n_2222),
.B(n_343),
.Y(n_2342)
);

AOI211x1_ASAP7_75t_L g2343 ( 
.A1(n_2189),
.A2(n_345),
.B(n_343),
.C(n_344),
.Y(n_2343)
);

INVxp67_ASAP7_75t_L g2344 ( 
.A(n_2222),
.Y(n_2344)
);

INVxp33_ASAP7_75t_L g2345 ( 
.A(n_2111),
.Y(n_2345)
);

OR2x2_ASAP7_75t_L g2346 ( 
.A(n_2199),
.B(n_344),
.Y(n_2346)
);

NAND2xp5_ASAP7_75t_L g2347 ( 
.A(n_2227),
.B(n_345),
.Y(n_2347)
);

INVxp67_ASAP7_75t_SL g2348 ( 
.A(n_2227),
.Y(n_2348)
);

A2O1A1Ixp33_ASAP7_75t_L g2349 ( 
.A1(n_2182),
.A2(n_348),
.B(n_346),
.C(n_347),
.Y(n_2349)
);

NAND3xp33_ASAP7_75t_L g2350 ( 
.A(n_2213),
.B(n_346),
.C(n_347),
.Y(n_2350)
);

NAND2xp33_ASAP7_75t_SL g2351 ( 
.A(n_2096),
.B(n_349),
.Y(n_2351)
);

NAND2xp5_ASAP7_75t_SL g2352 ( 
.A(n_2133),
.B(n_349),
.Y(n_2352)
);

AND2x2_ASAP7_75t_L g2353 ( 
.A(n_2198),
.B(n_2202),
.Y(n_2353)
);

NAND3xp33_ASAP7_75t_L g2354 ( 
.A(n_2210),
.B(n_609),
.C(n_610),
.Y(n_2354)
);

INVx1_ASAP7_75t_L g2355 ( 
.A(n_2217),
.Y(n_2355)
);

AND2x2_ASAP7_75t_L g2356 ( 
.A(n_2255),
.B(n_2116),
.Y(n_2356)
);

OR2x2_ASAP7_75t_L g2357 ( 
.A(n_2248),
.B(n_2233),
.Y(n_2357)
);

INVx1_ASAP7_75t_L g2358 ( 
.A(n_2341),
.Y(n_2358)
);

INVx1_ASAP7_75t_L g2359 ( 
.A(n_2247),
.Y(n_2359)
);

NAND2xp5_ASAP7_75t_L g2360 ( 
.A(n_2348),
.B(n_2212),
.Y(n_2360)
);

NAND2xp5_ASAP7_75t_L g2361 ( 
.A(n_2256),
.B(n_2215),
.Y(n_2361)
);

INVx1_ASAP7_75t_L g2362 ( 
.A(n_2259),
.Y(n_2362)
);

NAND2xp5_ASAP7_75t_L g2363 ( 
.A(n_2304),
.B(n_2224),
.Y(n_2363)
);

NAND2xp5_ASAP7_75t_L g2364 ( 
.A(n_2318),
.B(n_2225),
.Y(n_2364)
);

AND2x2_ASAP7_75t_L g2365 ( 
.A(n_2344),
.B(n_2123),
.Y(n_2365)
);

AOI221xp5_ASAP7_75t_L g2366 ( 
.A1(n_2311),
.A2(n_2238),
.B1(n_2219),
.B2(n_2173),
.C(n_2149),
.Y(n_2366)
);

NOR2x1_ASAP7_75t_SL g2367 ( 
.A(n_2291),
.B(n_2240),
.Y(n_2367)
);

AND2x2_ASAP7_75t_L g2368 ( 
.A(n_2276),
.B(n_2150),
.Y(n_2368)
);

NAND2xp5_ASAP7_75t_L g2369 ( 
.A(n_2302),
.B(n_2243),
.Y(n_2369)
);

INVx1_ASAP7_75t_L g2370 ( 
.A(n_2266),
.Y(n_2370)
);

NAND2xp5_ASAP7_75t_L g2371 ( 
.A(n_2296),
.B(n_2236),
.Y(n_2371)
);

AND2x2_ASAP7_75t_L g2372 ( 
.A(n_2353),
.B(n_2171),
.Y(n_2372)
);

INVx1_ASAP7_75t_L g2373 ( 
.A(n_2269),
.Y(n_2373)
);

INVx2_ASAP7_75t_L g2374 ( 
.A(n_2315),
.Y(n_2374)
);

NAND2xp5_ASAP7_75t_SL g2375 ( 
.A(n_2330),
.B(n_2290),
.Y(n_2375)
);

INVx1_ASAP7_75t_L g2376 ( 
.A(n_2270),
.Y(n_2376)
);

AND2x2_ASAP7_75t_L g2377 ( 
.A(n_2327),
.B(n_2112),
.Y(n_2377)
);

NAND2xp5_ASAP7_75t_L g2378 ( 
.A(n_2308),
.B(n_2168),
.Y(n_2378)
);

AOI22xp5_ASAP7_75t_L g2379 ( 
.A1(n_2350),
.A2(n_2203),
.B1(n_2146),
.B2(n_2132),
.Y(n_2379)
);

HB1xp67_ASAP7_75t_L g2380 ( 
.A(n_2298),
.Y(n_2380)
);

INVx1_ASAP7_75t_L g2381 ( 
.A(n_2272),
.Y(n_2381)
);

INVx1_ASAP7_75t_L g2382 ( 
.A(n_2279),
.Y(n_2382)
);

NOR2xp33_ASAP7_75t_L g2383 ( 
.A(n_2345),
.B(n_2147),
.Y(n_2383)
);

NAND2xp5_ASAP7_75t_L g2384 ( 
.A(n_2258),
.B(n_2137),
.Y(n_2384)
);

NAND2xp5_ASAP7_75t_L g2385 ( 
.A(n_2301),
.B(n_2128),
.Y(n_2385)
);

NAND2xp5_ASAP7_75t_L g2386 ( 
.A(n_2305),
.B(n_2161),
.Y(n_2386)
);

NAND2xp33_ASAP7_75t_SL g2387 ( 
.A(n_2287),
.B(n_2120),
.Y(n_2387)
);

NAND2xp5_ASAP7_75t_L g2388 ( 
.A(n_2252),
.B(n_2162),
.Y(n_2388)
);

NAND2xp5_ASAP7_75t_L g2389 ( 
.A(n_2286),
.B(n_2355),
.Y(n_2389)
);

INVx1_ASAP7_75t_L g2390 ( 
.A(n_2281),
.Y(n_2390)
);

INVx1_ASAP7_75t_L g2391 ( 
.A(n_2288),
.Y(n_2391)
);

NAND2xp5_ASAP7_75t_SL g2392 ( 
.A(n_2271),
.B(n_611),
.Y(n_2392)
);

INVxp67_ASAP7_75t_L g2393 ( 
.A(n_2351),
.Y(n_2393)
);

NAND2xp5_ASAP7_75t_L g2394 ( 
.A(n_2329),
.B(n_615),
.Y(n_2394)
);

BUFx2_ASAP7_75t_L g2395 ( 
.A(n_2298),
.Y(n_2395)
);

INVx1_ASAP7_75t_L g2396 ( 
.A(n_2294),
.Y(n_2396)
);

NAND2xp5_ASAP7_75t_L g2397 ( 
.A(n_2260),
.B(n_616),
.Y(n_2397)
);

NAND2xp5_ASAP7_75t_L g2398 ( 
.A(n_2320),
.B(n_618),
.Y(n_2398)
);

BUFx2_ASAP7_75t_L g2399 ( 
.A(n_2262),
.Y(n_2399)
);

INVx1_ASAP7_75t_L g2400 ( 
.A(n_2297),
.Y(n_2400)
);

NAND2xp5_ASAP7_75t_L g2401 ( 
.A(n_2325),
.B(n_619),
.Y(n_2401)
);

INVx1_ASAP7_75t_L g2402 ( 
.A(n_2300),
.Y(n_2402)
);

INVx1_ASAP7_75t_L g2403 ( 
.A(n_2309),
.Y(n_2403)
);

OR2x2_ASAP7_75t_L g2404 ( 
.A(n_2303),
.B(n_621),
.Y(n_2404)
);

NAND2xp5_ASAP7_75t_L g2405 ( 
.A(n_2328),
.B(n_622),
.Y(n_2405)
);

NAND2xp5_ASAP7_75t_L g2406 ( 
.A(n_2334),
.B(n_624),
.Y(n_2406)
);

AOI221xp5_ASAP7_75t_L g2407 ( 
.A1(n_2246),
.A2(n_2249),
.B1(n_2275),
.B2(n_2268),
.C(n_2289),
.Y(n_2407)
);

AOI22xp33_ASAP7_75t_L g2408 ( 
.A1(n_2263),
.A2(n_629),
.B1(n_626),
.B2(n_627),
.Y(n_2408)
);

NAND2xp5_ASAP7_75t_L g2409 ( 
.A(n_2336),
.B(n_631),
.Y(n_2409)
);

INVx1_ASAP7_75t_SL g2410 ( 
.A(n_2278),
.Y(n_2410)
);

CKINVDCx5p33_ASAP7_75t_R g2411 ( 
.A(n_2399),
.Y(n_2411)
);

INVx2_ASAP7_75t_L g2412 ( 
.A(n_2368),
.Y(n_2412)
);

INVx1_ASAP7_75t_L g2413 ( 
.A(n_2380),
.Y(n_2413)
);

INVx1_ASAP7_75t_L g2414 ( 
.A(n_2395),
.Y(n_2414)
);

AND2x2_ASAP7_75t_L g2415 ( 
.A(n_2356),
.B(n_2340),
.Y(n_2415)
);

INVxp67_ASAP7_75t_L g2416 ( 
.A(n_2387),
.Y(n_2416)
);

HB1xp67_ASAP7_75t_L g2417 ( 
.A(n_2393),
.Y(n_2417)
);

INVx1_ASAP7_75t_L g2418 ( 
.A(n_2365),
.Y(n_2418)
);

INVx1_ASAP7_75t_L g2419 ( 
.A(n_2374),
.Y(n_2419)
);

NAND2xp5_ASAP7_75t_SL g2420 ( 
.A(n_2407),
.B(n_2257),
.Y(n_2420)
);

INVx1_ASAP7_75t_L g2421 ( 
.A(n_2359),
.Y(n_2421)
);

INVx1_ASAP7_75t_SL g2422 ( 
.A(n_2410),
.Y(n_2422)
);

NAND2xp5_ASAP7_75t_L g2423 ( 
.A(n_2372),
.B(n_2322),
.Y(n_2423)
);

INVx1_ASAP7_75t_L g2424 ( 
.A(n_2362),
.Y(n_2424)
);

INVx1_ASAP7_75t_L g2425 ( 
.A(n_2370),
.Y(n_2425)
);

NOR2xp33_ASAP7_75t_L g2426 ( 
.A(n_2375),
.B(n_2335),
.Y(n_2426)
);

INVx1_ASAP7_75t_L g2427 ( 
.A(n_2373),
.Y(n_2427)
);

INVx1_ASAP7_75t_L g2428 ( 
.A(n_2376),
.Y(n_2428)
);

INVx1_ASAP7_75t_L g2429 ( 
.A(n_2381),
.Y(n_2429)
);

INVx1_ASAP7_75t_L g2430 ( 
.A(n_2382),
.Y(n_2430)
);

INVx1_ASAP7_75t_L g2431 ( 
.A(n_2390),
.Y(n_2431)
);

INVx1_ASAP7_75t_L g2432 ( 
.A(n_2391),
.Y(n_2432)
);

INVx1_ASAP7_75t_L g2433 ( 
.A(n_2396),
.Y(n_2433)
);

HB1xp67_ASAP7_75t_L g2434 ( 
.A(n_2363),
.Y(n_2434)
);

INVx1_ASAP7_75t_L g2435 ( 
.A(n_2400),
.Y(n_2435)
);

INVx2_ASAP7_75t_L g2436 ( 
.A(n_2367),
.Y(n_2436)
);

INVxp67_ASAP7_75t_L g2437 ( 
.A(n_2361),
.Y(n_2437)
);

INVx1_ASAP7_75t_L g2438 ( 
.A(n_2402),
.Y(n_2438)
);

INVx2_ASAP7_75t_L g2439 ( 
.A(n_2377),
.Y(n_2439)
);

NOR2xp33_ASAP7_75t_L g2440 ( 
.A(n_2384),
.B(n_2310),
.Y(n_2440)
);

INVx1_ASAP7_75t_L g2441 ( 
.A(n_2403),
.Y(n_2441)
);

INVx1_ASAP7_75t_L g2442 ( 
.A(n_2358),
.Y(n_2442)
);

OA211x2_ASAP7_75t_L g2443 ( 
.A1(n_2416),
.A2(n_2378),
.B(n_2332),
.C(n_2333),
.Y(n_2443)
);

OAI21xp33_ASAP7_75t_L g2444 ( 
.A1(n_2420),
.A2(n_2386),
.B(n_2389),
.Y(n_2444)
);

NOR2xp33_ASAP7_75t_L g2445 ( 
.A(n_2411),
.B(n_2422),
.Y(n_2445)
);

NOR3xp33_ASAP7_75t_L g2446 ( 
.A(n_2426),
.B(n_2383),
.C(n_2366),
.Y(n_2446)
);

AOI211xp5_ASAP7_75t_L g2447 ( 
.A1(n_2440),
.A2(n_2267),
.B(n_2277),
.C(n_2284),
.Y(n_2447)
);

NAND3xp33_ASAP7_75t_SL g2448 ( 
.A(n_2422),
.B(n_2339),
.C(n_2299),
.Y(n_2448)
);

OAI21xp33_ASAP7_75t_L g2449 ( 
.A1(n_2417),
.A2(n_2371),
.B(n_2360),
.Y(n_2449)
);

NOR2xp67_ASAP7_75t_L g2450 ( 
.A(n_2436),
.B(n_2364),
.Y(n_2450)
);

INVxp67_ASAP7_75t_SL g2451 ( 
.A(n_2414),
.Y(n_2451)
);

O2A1O1Ixp33_ASAP7_75t_L g2452 ( 
.A1(n_2413),
.A2(n_2394),
.B(n_2261),
.C(n_2253),
.Y(n_2452)
);

AOI211xp5_ASAP7_75t_L g2453 ( 
.A1(n_2437),
.A2(n_2283),
.B(n_2317),
.C(n_2313),
.Y(n_2453)
);

NAND3xp33_ASAP7_75t_L g2454 ( 
.A(n_2434),
.B(n_2295),
.C(n_2354),
.Y(n_2454)
);

NAND2xp5_ASAP7_75t_L g2455 ( 
.A(n_2415),
.B(n_2369),
.Y(n_2455)
);

NOR2x1_ASAP7_75t_L g2456 ( 
.A(n_2418),
.B(n_2388),
.Y(n_2456)
);

AND4x1_ASAP7_75t_L g2457 ( 
.A(n_2419),
.B(n_2349),
.C(n_2293),
.D(n_2265),
.Y(n_2457)
);

NOR3x1_ASAP7_75t_L g2458 ( 
.A(n_2423),
.B(n_2385),
.C(n_2357),
.Y(n_2458)
);

NAND3x1_ASAP7_75t_L g2459 ( 
.A(n_2442),
.B(n_2264),
.C(n_2251),
.Y(n_2459)
);

NAND4xp75_ASAP7_75t_L g2460 ( 
.A(n_2421),
.B(n_2343),
.C(n_2282),
.D(n_2424),
.Y(n_2460)
);

OAI221xp5_ASAP7_75t_L g2461 ( 
.A1(n_2444),
.A2(n_2412),
.B1(n_2439),
.B2(n_2338),
.C(n_2319),
.Y(n_2461)
);

OAI221xp5_ASAP7_75t_SL g2462 ( 
.A1(n_2452),
.A2(n_2312),
.B1(n_2316),
.B2(n_2379),
.C(n_2254),
.Y(n_2462)
);

BUFx2_ASAP7_75t_L g2463 ( 
.A(n_2451),
.Y(n_2463)
);

OAI221xp5_ASAP7_75t_L g2464 ( 
.A1(n_2454),
.A2(n_2306),
.B1(n_2379),
.B2(n_2392),
.C(n_2352),
.Y(n_2464)
);

NAND5xp2_ASAP7_75t_L g2465 ( 
.A(n_2446),
.B(n_2425),
.C(n_2429),
.D(n_2428),
.E(n_2427),
.Y(n_2465)
);

AOI221xp5_ASAP7_75t_L g2466 ( 
.A1(n_2448),
.A2(n_2431),
.B1(n_2433),
.B2(n_2432),
.C(n_2430),
.Y(n_2466)
);

INVx1_ASAP7_75t_SL g2467 ( 
.A(n_2456),
.Y(n_2467)
);

OAI211xp5_ASAP7_75t_L g2468 ( 
.A1(n_2453),
.A2(n_2321),
.B(n_2438),
.C(n_2435),
.Y(n_2468)
);

INVx1_ASAP7_75t_SL g2469 ( 
.A(n_2459),
.Y(n_2469)
);

OR2x2_ASAP7_75t_L g2470 ( 
.A(n_2463),
.B(n_2455),
.Y(n_2470)
);

NOR2xp33_ASAP7_75t_L g2471 ( 
.A(n_2462),
.B(n_2445),
.Y(n_2471)
);

XNOR2xp5_ASAP7_75t_L g2472 ( 
.A(n_2464),
.B(n_2457),
.Y(n_2472)
);

NOR2xp67_ASAP7_75t_L g2473 ( 
.A(n_2468),
.B(n_2450),
.Y(n_2473)
);

NAND2xp5_ASAP7_75t_L g2474 ( 
.A(n_2469),
.B(n_2447),
.Y(n_2474)
);

NOR3xp33_ASAP7_75t_SL g2475 ( 
.A(n_2465),
.B(n_2449),
.C(n_2460),
.Y(n_2475)
);

NOR2x1_ASAP7_75t_L g2476 ( 
.A(n_2467),
.B(n_2274),
.Y(n_2476)
);

INVx1_ASAP7_75t_L g2477 ( 
.A(n_2461),
.Y(n_2477)
);

NAND3xp33_ASAP7_75t_L g2478 ( 
.A(n_2475),
.B(n_2466),
.C(n_2441),
.Y(n_2478)
);

NAND2xp5_ASAP7_75t_SL g2479 ( 
.A(n_2473),
.B(n_2324),
.Y(n_2479)
);

NOR2xp33_ASAP7_75t_R g2480 ( 
.A(n_2470),
.B(n_2331),
.Y(n_2480)
);

NAND3xp33_ASAP7_75t_L g2481 ( 
.A(n_2472),
.B(n_2397),
.C(n_2401),
.Y(n_2481)
);

NAND2xp5_ASAP7_75t_SL g2482 ( 
.A(n_2476),
.B(n_2285),
.Y(n_2482)
);

NOR2xp33_ASAP7_75t_L g2483 ( 
.A(n_2482),
.B(n_2474),
.Y(n_2483)
);

NAND2xp5_ASAP7_75t_L g2484 ( 
.A(n_2480),
.B(n_2471),
.Y(n_2484)
);

INVxp67_ASAP7_75t_L g2485 ( 
.A(n_2483),
.Y(n_2485)
);

NAND5xp2_ASAP7_75t_L g2486 ( 
.A(n_2485),
.B(n_2477),
.C(n_2484),
.D(n_2478),
.E(n_2479),
.Y(n_2486)
);

AOI22xp33_ASAP7_75t_L g2487 ( 
.A1(n_2486),
.A2(n_2443),
.B1(n_2481),
.B2(n_2250),
.Y(n_2487)
);

AOI22xp33_ASAP7_75t_L g2488 ( 
.A1(n_2486),
.A2(n_2458),
.B1(n_2273),
.B2(n_2280),
.Y(n_2488)
);

AO22x2_ASAP7_75t_L g2489 ( 
.A1(n_2487),
.A2(n_2326),
.B1(n_2323),
.B2(n_2337),
.Y(n_2489)
);

NAND2xp5_ASAP7_75t_L g2490 ( 
.A(n_2488),
.B(n_2314),
.Y(n_2490)
);

AOI21xp5_ASAP7_75t_L g2491 ( 
.A1(n_2490),
.A2(n_2307),
.B(n_2292),
.Y(n_2491)
);

OAI22xp5_ASAP7_75t_L g2492 ( 
.A1(n_2489),
.A2(n_2346),
.B1(n_2347),
.B2(n_2342),
.Y(n_2492)
);

INVx1_ASAP7_75t_L g2493 ( 
.A(n_2492),
.Y(n_2493)
);

INVx1_ASAP7_75t_L g2494 ( 
.A(n_2491),
.Y(n_2494)
);

OAI221xp5_ASAP7_75t_R g2495 ( 
.A1(n_2493),
.A2(n_2408),
.B1(n_2404),
.B2(n_2398),
.C(n_2406),
.Y(n_2495)
);

AOI211xp5_ASAP7_75t_L g2496 ( 
.A1(n_2495),
.A2(n_2494),
.B(n_2409),
.C(n_2405),
.Y(n_2496)
);


endmodule