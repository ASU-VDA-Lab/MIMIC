module fake_jpeg_27028_n_76 (n_13, n_21, n_1, n_10, n_6, n_22, n_14, n_19, n_18, n_20, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_76);

input n_13;
input n_21;
input n_1;
input n_10;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_76;

wire n_57;
wire n_53;
wire n_33;
wire n_54;
wire n_61;
wire n_45;
wire n_23;
wire n_69;
wire n_27;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_40;
wire n_73;
wire n_71;
wire n_35;
wire n_48;
wire n_68;
wire n_52;
wire n_59;
wire n_46;
wire n_58;
wire n_41;
wire n_60;
wire n_65;
wire n_63;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_49;
wire n_72;
wire n_24;
wire n_28;
wire n_44;
wire n_26;
wire n_38;
wire n_36;
wire n_74;
wire n_62;
wire n_25;
wire n_31;
wire n_56;
wire n_67;
wire n_75;
wire n_29;
wire n_37;
wire n_50;
wire n_43;
wire n_32;
wire n_70;
wire n_66;

INVx1_ASAP7_75t_L g23 ( 
.A(n_15),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_11),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_3),
.Y(n_25)
);

INVx4_ASAP7_75t_L g26 ( 
.A(n_21),
.Y(n_26)
);

INVx13_ASAP7_75t_L g27 ( 
.A(n_9),
.Y(n_27)
);

INVx2_ASAP7_75t_L g28 ( 
.A(n_3),
.Y(n_28)
);

CKINVDCx9p33_ASAP7_75t_R g29 ( 
.A(n_18),
.Y(n_29)
);

OR2x2_ASAP7_75t_SL g30 ( 
.A(n_22),
.B(n_0),
.Y(n_30)
);

INVx5_ASAP7_75t_L g31 ( 
.A(n_0),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_4),
.Y(n_32)
);

INVx2_ASAP7_75t_L g33 ( 
.A(n_14),
.Y(n_33)
);

BUFx3_ASAP7_75t_L g34 ( 
.A(n_6),
.Y(n_34)
);

NAND2xp5_ASAP7_75t_L g35 ( 
.A(n_17),
.B(n_19),
.Y(n_35)
);

INVx3_ASAP7_75t_L g36 ( 
.A(n_10),
.Y(n_36)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_16),
.Y(n_37)
);

INVx4_ASAP7_75t_L g38 ( 
.A(n_4),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_20),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_1),
.Y(n_40)
);

INVx11_ASAP7_75t_L g41 ( 
.A(n_7),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_8),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_5),
.Y(n_43)
);

INVx8_ASAP7_75t_L g44 ( 
.A(n_2),
.Y(n_44)
);

INVx6_ASAP7_75t_L g45 ( 
.A(n_39),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_45),
.B(n_46),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_L g46 ( 
.A(n_35),
.B(n_1),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g47 ( 
.A(n_30),
.B(n_2),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_47),
.B(n_48),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_SL g48 ( 
.A(n_25),
.B(n_12),
.Y(n_48)
);

INVxp67_ASAP7_75t_L g49 ( 
.A(n_29),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_L g59 ( 
.A(n_49),
.B(n_50),
.Y(n_59)
);

BUFx2_ASAP7_75t_L g50 ( 
.A(n_27),
.Y(n_50)
);

OAI22xp5_ASAP7_75t_SL g51 ( 
.A1(n_36),
.A2(n_33),
.B1(n_26),
.B2(n_28),
.Y(n_51)
);

OAI22xp5_ASAP7_75t_SL g60 ( 
.A1(n_51),
.A2(n_57),
.B1(n_58),
.B2(n_31),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_SL g52 ( 
.A(n_32),
.B(n_13),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_L g62 ( 
.A(n_52),
.B(n_53),
.Y(n_62)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_24),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_SL g54 ( 
.A(n_40),
.B(n_27),
.Y(n_54)
);

MAJIxp5_ASAP7_75t_L g65 ( 
.A(n_54),
.B(n_55),
.C(n_56),
.Y(n_65)
);

INVx1_ASAP7_75t_SL g55 ( 
.A(n_34),
.Y(n_55)
);

INVx11_ASAP7_75t_L g56 ( 
.A(n_39),
.Y(n_56)
);

INVx8_ASAP7_75t_L g57 ( 
.A(n_41),
.Y(n_57)
);

INVx13_ASAP7_75t_L g58 ( 
.A(n_42),
.Y(n_58)
);

AOI22xp5_ASAP7_75t_L g67 ( 
.A1(n_60),
.A2(n_61),
.B1(n_44),
.B2(n_49),
.Y(n_67)
);

OAI22xp5_ASAP7_75t_SL g61 ( 
.A1(n_45),
.A2(n_23),
.B1(n_37),
.B2(n_38),
.Y(n_61)
);

OAI22xp5_ASAP7_75t_SL g66 ( 
.A1(n_64),
.A2(n_58),
.B1(n_65),
.B2(n_44),
.Y(n_66)
);

XNOR2xp5_ASAP7_75t_SL g70 ( 
.A(n_66),
.B(n_68),
.Y(n_70)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_67),
.Y(n_71)
);

XOR2xp5_ASAP7_75t_L g68 ( 
.A(n_64),
.B(n_42),
.Y(n_68)
);

XNOR2xp5_ASAP7_75t_SL g69 ( 
.A(n_63),
.B(n_43),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_L g72 ( 
.A(n_71),
.B(n_62),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_72),
.B(n_73),
.Y(n_74)
);

A2O1A1Ixp33_ASAP7_75t_SL g73 ( 
.A1(n_70),
.A2(n_69),
.B(n_43),
.C(n_50),
.Y(n_73)
);

OAI21xp5_ASAP7_75t_SL g75 ( 
.A1(n_74),
.A2(n_69),
.B(n_59),
.Y(n_75)
);

XOR2xp5_ASAP7_75t_L g76 ( 
.A(n_75),
.B(n_57),
.Y(n_76)
);


endmodule