module fake_jpeg_25868_n_380 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_380);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_380;

wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_340;
wire n_377;
wire n_291;
wire n_236;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_370;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_137;
wire n_74;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_368;
wire n_298;
wire n_106;
wire n_327;
wire n_122;
wire n_75;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_39;
wire n_371;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_367;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_360;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_378;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_379;
wire n_114;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_356;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_375;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVx2_ASAP7_75t_L g17 ( 
.A(n_4),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_16),
.Y(n_18)
);

INVx2_ASAP7_75t_L g19 ( 
.A(n_0),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_1),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_14),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_5),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_11),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_4),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_5),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_8),
.Y(n_26)
);

INVx2_ASAP7_75t_L g27 ( 
.A(n_8),
.Y(n_27)
);

CKINVDCx16_ASAP7_75t_R g28 ( 
.A(n_6),
.Y(n_28)
);

INVx8_ASAP7_75t_L g29 ( 
.A(n_8),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_8),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_6),
.Y(n_31)
);

NOR2xp33_ASAP7_75t_L g32 ( 
.A(n_3),
.B(n_2),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_5),
.Y(n_33)
);

INVx2_ASAP7_75t_L g34 ( 
.A(n_2),
.Y(n_34)
);

BUFx12f_ASAP7_75t_L g35 ( 
.A(n_12),
.Y(n_35)
);

BUFx3_ASAP7_75t_L g36 ( 
.A(n_5),
.Y(n_36)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_14),
.Y(n_37)
);

INVx2_ASAP7_75t_L g38 ( 
.A(n_1),
.Y(n_38)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_1),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_15),
.Y(n_40)
);

INVx2_ASAP7_75t_L g41 ( 
.A(n_17),
.Y(n_41)
);

INVx2_ASAP7_75t_L g79 ( 
.A(n_41),
.Y(n_79)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_35),
.Y(n_42)
);

INVx6_ASAP7_75t_L g78 ( 
.A(n_42),
.Y(n_78)
);

INVx2_ASAP7_75t_L g43 ( 
.A(n_17),
.Y(n_43)
);

INVx2_ASAP7_75t_L g106 ( 
.A(n_43),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g44 ( 
.A(n_32),
.B(n_16),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_SL g108 ( 
.A(n_44),
.B(n_57),
.Y(n_108)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_35),
.Y(n_45)
);

INVx6_ASAP7_75t_L g80 ( 
.A(n_45),
.Y(n_80)
);

INVx6_ASAP7_75t_L g46 ( 
.A(n_22),
.Y(n_46)
);

INVx3_ASAP7_75t_L g72 ( 
.A(n_46),
.Y(n_72)
);

AOI22xp5_ASAP7_75t_L g47 ( 
.A1(n_19),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_47)
);

OAI22xp5_ASAP7_75t_SL g82 ( 
.A1(n_47),
.A2(n_20),
.B1(n_33),
.B2(n_31),
.Y(n_82)
);

BUFx12f_ASAP7_75t_L g48 ( 
.A(n_35),
.Y(n_48)
);

BUFx12f_ASAP7_75t_L g86 ( 
.A(n_48),
.Y(n_86)
);

INVx3_ASAP7_75t_L g49 ( 
.A(n_40),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g97 ( 
.A(n_49),
.Y(n_97)
);

BUFx3_ASAP7_75t_L g50 ( 
.A(n_35),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_50),
.B(n_59),
.Y(n_89)
);

BUFx12f_ASAP7_75t_L g51 ( 
.A(n_35),
.Y(n_51)
);

BUFx12f_ASAP7_75t_L g105 ( 
.A(n_51),
.Y(n_105)
);

BUFx5_ASAP7_75t_L g52 ( 
.A(n_22),
.Y(n_52)
);

BUFx3_ASAP7_75t_L g102 ( 
.A(n_52),
.Y(n_102)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_19),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g109 ( 
.A(n_53),
.Y(n_109)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_32),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_L g88 ( 
.A(n_54),
.B(n_56),
.Y(n_88)
);

INVx3_ASAP7_75t_L g55 ( 
.A(n_40),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g112 ( 
.A(n_55),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_L g56 ( 
.A(n_27),
.B(n_0),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g57 ( 
.A(n_18),
.B(n_16),
.Y(n_57)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_29),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_L g96 ( 
.A(n_58),
.B(n_70),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_SL g59 ( 
.A(n_18),
.B(n_21),
.Y(n_59)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_27),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g113 ( 
.A(n_60),
.Y(n_113)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_34),
.Y(n_61)
);

INVx4_ASAP7_75t_L g71 ( 
.A(n_61),
.Y(n_71)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_34),
.Y(n_62)
);

INVx4_ASAP7_75t_L g73 ( 
.A(n_62),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_21),
.B(n_15),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_63),
.B(n_69),
.Y(n_99)
);

INVx6_ASAP7_75t_SL g64 ( 
.A(n_36),
.Y(n_64)
);

CKINVDCx16_ASAP7_75t_R g111 ( 
.A(n_64),
.Y(n_111)
);

INVx8_ASAP7_75t_L g65 ( 
.A(n_29),
.Y(n_65)
);

INVx5_ASAP7_75t_L g94 ( 
.A(n_65),
.Y(n_94)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_38),
.Y(n_66)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_66),
.Y(n_74)
);

INVx2_ASAP7_75t_L g67 ( 
.A(n_38),
.Y(n_67)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_67),
.Y(n_84)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_29),
.Y(n_68)
);

INVx4_ASAP7_75t_L g75 ( 
.A(n_68),
.Y(n_75)
);

INVx3_ASAP7_75t_L g69 ( 
.A(n_40),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_37),
.B(n_15),
.Y(n_70)
);

INVx3_ASAP7_75t_L g76 ( 
.A(n_42),
.Y(n_76)
);

INVx6_ASAP7_75t_L g138 ( 
.A(n_76),
.Y(n_138)
);

INVx2_ASAP7_75t_SL g77 ( 
.A(n_45),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g142 ( 
.A(n_77),
.B(n_81),
.Y(n_142)
);

A2O1A1Ixp33_ASAP7_75t_L g81 ( 
.A1(n_56),
.A2(n_37),
.B(n_28),
.C(n_25),
.Y(n_81)
);

AOI22xp5_ASAP7_75t_L g128 ( 
.A1(n_82),
.A2(n_90),
.B1(n_93),
.B2(n_0),
.Y(n_128)
);

AOI22xp33_ASAP7_75t_SL g83 ( 
.A1(n_46),
.A2(n_25),
.B1(n_24),
.B2(n_39),
.Y(n_83)
);

AOI22xp33_ASAP7_75t_SL g117 ( 
.A1(n_83),
.A2(n_91),
.B1(n_69),
.B2(n_58),
.Y(n_117)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_65),
.Y(n_85)
);

INVxp33_ASAP7_75t_L g132 ( 
.A(n_85),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_L g87 ( 
.A(n_54),
.B(n_39),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_L g123 ( 
.A(n_87),
.B(n_98),
.Y(n_123)
);

OAI22xp5_ASAP7_75t_SL g90 ( 
.A1(n_47),
.A2(n_26),
.B1(n_33),
.B2(n_31),
.Y(n_90)
);

AOI22xp33_ASAP7_75t_SL g91 ( 
.A1(n_49),
.A2(n_24),
.B1(n_23),
.B2(n_20),
.Y(n_91)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_41),
.Y(n_92)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_92),
.Y(n_114)
);

OAI22xp5_ASAP7_75t_L g93 ( 
.A1(n_55),
.A2(n_23),
.B1(n_30),
.B2(n_26),
.Y(n_93)
);

AND2x2_ASAP7_75t_SL g95 ( 
.A(n_53),
.B(n_22),
.Y(n_95)
);

AND2x2_ASAP7_75t_L g133 ( 
.A(n_95),
.B(n_100),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_L g98 ( 
.A(n_43),
.B(n_30),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g100 ( 
.A(n_60),
.B(n_28),
.Y(n_100)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_66),
.Y(n_101)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_101),
.Y(n_129)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_67),
.Y(n_103)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_103),
.Y(n_146)
);

INVx4_ASAP7_75t_L g104 ( 
.A(n_48),
.Y(n_104)
);

INVx2_ASAP7_75t_L g131 ( 
.A(n_104),
.Y(n_131)
);

INVx11_ASAP7_75t_L g107 ( 
.A(n_48),
.Y(n_107)
);

INVx5_ASAP7_75t_L g116 ( 
.A(n_107),
.Y(n_116)
);

CKINVDCx20_ASAP7_75t_R g110 ( 
.A(n_61),
.Y(n_110)
);

CKINVDCx20_ASAP7_75t_R g126 ( 
.A(n_110),
.Y(n_126)
);

HB1xp67_ASAP7_75t_L g115 ( 
.A(n_98),
.Y(n_115)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_115),
.Y(n_168)
);

AOI22xp5_ASAP7_75t_SL g165 ( 
.A1(n_117),
.A2(n_140),
.B1(n_141),
.B2(n_151),
.Y(n_165)
);

INVx4_ASAP7_75t_L g118 ( 
.A(n_107),
.Y(n_118)
);

BUFx6f_ASAP7_75t_L g160 ( 
.A(n_118),
.Y(n_160)
);

AOI22xp33_ASAP7_75t_L g119 ( 
.A1(n_71),
.A2(n_62),
.B1(n_22),
.B2(n_68),
.Y(n_119)
);

AOI22xp5_ASAP7_75t_L g178 ( 
.A1(n_119),
.A2(n_120),
.B1(n_122),
.B2(n_125),
.Y(n_178)
);

OAI22xp5_ASAP7_75t_SL g120 ( 
.A1(n_88),
.A2(n_71),
.B1(n_73),
.B2(n_72),
.Y(n_120)
);

AOI22xp33_ASAP7_75t_SL g121 ( 
.A1(n_94),
.A2(n_14),
.B1(n_13),
.B2(n_36),
.Y(n_121)
);

AOI22xp33_ASAP7_75t_SL g179 ( 
.A1(n_121),
.A2(n_124),
.B1(n_130),
.B2(n_134),
.Y(n_179)
);

OAI22xp33_ASAP7_75t_SL g122 ( 
.A1(n_82),
.A2(n_52),
.B1(n_36),
.B2(n_64),
.Y(n_122)
);

AOI22xp33_ASAP7_75t_SL g124 ( 
.A1(n_94),
.A2(n_13),
.B1(n_2),
.B2(n_3),
.Y(n_124)
);

OAI22xp5_ASAP7_75t_L g125 ( 
.A1(n_95),
.A2(n_50),
.B1(n_51),
.B2(n_13),
.Y(n_125)
);

INVxp67_ASAP7_75t_L g127 ( 
.A(n_91),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_L g159 ( 
.A(n_127),
.B(n_136),
.Y(n_159)
);

OR2x2_ASAP7_75t_L g157 ( 
.A(n_128),
.B(n_108),
.Y(n_157)
);

AOI22xp33_ASAP7_75t_SL g130 ( 
.A1(n_75),
.A2(n_3),
.B1(n_4),
.B2(n_6),
.Y(n_130)
);

INVx5_ASAP7_75t_L g134 ( 
.A(n_86),
.Y(n_134)
);

OAI22xp5_ASAP7_75t_L g135 ( 
.A1(n_95),
.A2(n_51),
.B1(n_4),
.B2(n_6),
.Y(n_135)
);

OAI22xp5_ASAP7_75t_SL g156 ( 
.A1(n_135),
.A2(n_143),
.B1(n_145),
.B2(n_148),
.Y(n_156)
);

INVx3_ASAP7_75t_L g136 ( 
.A(n_113),
.Y(n_136)
);

INVx2_ASAP7_75t_L g137 ( 
.A(n_79),
.Y(n_137)
);

INVx2_ASAP7_75t_L g158 ( 
.A(n_137),
.Y(n_158)
);

AND2x4_ASAP7_75t_SL g139 ( 
.A(n_81),
.B(n_3),
.Y(n_139)
);

AND2x2_ASAP7_75t_L g172 ( 
.A(n_139),
.B(n_86),
.Y(n_172)
);

OAI22xp5_ASAP7_75t_SL g140 ( 
.A1(n_73),
.A2(n_7),
.B1(n_9),
.B2(n_10),
.Y(n_140)
);

AOI22xp33_ASAP7_75t_SL g141 ( 
.A1(n_75),
.A2(n_12),
.B1(n_9),
.B2(n_10),
.Y(n_141)
);

AOI22xp5_ASAP7_75t_L g143 ( 
.A1(n_90),
.A2(n_7),
.B1(n_9),
.B2(n_10),
.Y(n_143)
);

INVx2_ASAP7_75t_L g144 ( 
.A(n_79),
.Y(n_144)
);

INVx2_ASAP7_75t_L g162 ( 
.A(n_144),
.Y(n_162)
);

AOI22xp33_ASAP7_75t_L g145 ( 
.A1(n_72),
.A2(n_7),
.B1(n_9),
.B2(n_10),
.Y(n_145)
);

INVx2_ASAP7_75t_L g147 ( 
.A(n_106),
.Y(n_147)
);

INVx2_ASAP7_75t_L g174 ( 
.A(n_147),
.Y(n_174)
);

O2A1O1Ixp33_ASAP7_75t_L g148 ( 
.A1(n_106),
.A2(n_84),
.B(n_74),
.C(n_83),
.Y(n_148)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_87),
.Y(n_149)
);

NOR2xp33_ASAP7_75t_L g161 ( 
.A(n_149),
.B(n_152),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_L g150 ( 
.A(n_99),
.B(n_7),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_L g170 ( 
.A(n_150),
.B(n_111),
.Y(n_170)
);

AOI22xp33_ASAP7_75t_SL g151 ( 
.A1(n_104),
.A2(n_78),
.B1(n_80),
.B2(n_76),
.Y(n_151)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_96),
.Y(n_152)
);

AOI22xp33_ASAP7_75t_L g153 ( 
.A1(n_78),
.A2(n_11),
.B1(n_12),
.B2(n_80),
.Y(n_153)
);

OAI22xp5_ASAP7_75t_SL g188 ( 
.A1(n_153),
.A2(n_154),
.B1(n_155),
.B2(n_102),
.Y(n_188)
);

AOI22xp33_ASAP7_75t_L g154 ( 
.A1(n_77),
.A2(n_11),
.B1(n_12),
.B2(n_109),
.Y(n_154)
);

AOI22xp33_ASAP7_75t_SL g155 ( 
.A1(n_102),
.A2(n_11),
.B1(n_89),
.B2(n_97),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_SL g208 ( 
.A(n_157),
.B(n_170),
.Y(n_208)
);

CKINVDCx20_ASAP7_75t_R g163 ( 
.A(n_126),
.Y(n_163)
);

NOR2xp33_ASAP7_75t_L g198 ( 
.A(n_163),
.B(n_167),
.Y(n_198)
);

NOR2xp33_ASAP7_75t_L g164 ( 
.A(n_149),
.B(n_113),
.Y(n_164)
);

NOR2xp33_ASAP7_75t_SL g205 ( 
.A(n_164),
.B(n_166),
.Y(n_205)
);

NOR2xp33_ASAP7_75t_L g166 ( 
.A(n_152),
.B(n_97),
.Y(n_166)
);

CKINVDCx20_ASAP7_75t_R g167 ( 
.A(n_126),
.Y(n_167)
);

NOR2xp33_ASAP7_75t_L g169 ( 
.A(n_123),
.B(n_112),
.Y(n_169)
);

NOR2xp33_ASAP7_75t_L g203 ( 
.A(n_169),
.B(n_171),
.Y(n_203)
);

NOR2xp33_ASAP7_75t_L g171 ( 
.A(n_123),
.B(n_112),
.Y(n_171)
);

OAI21xp5_ASAP7_75t_SL g207 ( 
.A1(n_172),
.A2(n_173),
.B(n_175),
.Y(n_207)
);

AND2x2_ASAP7_75t_L g173 ( 
.A(n_142),
.B(n_135),
.Y(n_173)
);

AND2x2_ASAP7_75t_L g175 ( 
.A(n_142),
.B(n_109),
.Y(n_175)
);

CKINVDCx20_ASAP7_75t_R g176 ( 
.A(n_120),
.Y(n_176)
);

CKINVDCx20_ASAP7_75t_R g224 ( 
.A(n_176),
.Y(n_224)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_148),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_SL g215 ( 
.A(n_177),
.B(n_180),
.Y(n_215)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_148),
.Y(n_180)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_115),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_SL g220 ( 
.A(n_181),
.B(n_182),
.Y(n_220)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_137),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_L g183 ( 
.A(n_133),
.B(n_86),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_L g195 ( 
.A(n_183),
.B(n_184),
.Y(n_195)
);

NOR2xp33_ASAP7_75t_L g184 ( 
.A(n_150),
.B(n_105),
.Y(n_184)
);

INVx13_ASAP7_75t_L g185 ( 
.A(n_134),
.Y(n_185)
);

INVx13_ASAP7_75t_L g196 ( 
.A(n_185),
.Y(n_196)
);

NAND2xp5_ASAP7_75t_SL g186 ( 
.A(n_133),
.B(n_105),
.Y(n_186)
);

CKINVDCx16_ASAP7_75t_R g217 ( 
.A(n_186),
.Y(n_217)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_144),
.Y(n_187)
);

NOR2xp33_ASAP7_75t_L g201 ( 
.A(n_187),
.B(n_190),
.Y(n_201)
);

AOI22xp33_ASAP7_75t_L g218 ( 
.A1(n_188),
.A2(n_134),
.B1(n_116),
.B2(n_118),
.Y(n_218)
);

INVx2_ASAP7_75t_L g189 ( 
.A(n_147),
.Y(n_189)
);

BUFx24_ASAP7_75t_L g226 ( 
.A(n_189),
.Y(n_226)
);

INVx2_ASAP7_75t_L g190 ( 
.A(n_131),
.Y(n_190)
);

NOR2xp33_ASAP7_75t_SL g191 ( 
.A(n_139),
.B(n_105),
.Y(n_191)
);

NOR2xp33_ASAP7_75t_L g212 ( 
.A(n_191),
.B(n_132),
.Y(n_212)
);

NAND2xp5_ASAP7_75t_SL g192 ( 
.A(n_133),
.B(n_128),
.Y(n_192)
);

OAI21xp5_ASAP7_75t_SL g211 ( 
.A1(n_192),
.A2(n_129),
.B(n_146),
.Y(n_211)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_166),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_SL g229 ( 
.A(n_193),
.B(n_204),
.Y(n_229)
);

MAJIxp5_ASAP7_75t_SL g194 ( 
.A(n_178),
.B(n_143),
.C(n_125),
.Y(n_194)
);

OAI21xp5_ASAP7_75t_SL g248 ( 
.A1(n_194),
.A2(n_210),
.B(n_211),
.Y(n_248)
);

AOI22xp5_ASAP7_75t_L g197 ( 
.A1(n_177),
.A2(n_139),
.B1(n_140),
.B2(n_136),
.Y(n_197)
);

OAI22xp5_ASAP7_75t_SL g242 ( 
.A1(n_197),
.A2(n_200),
.B1(n_202),
.B2(n_206),
.Y(n_242)
);

INVxp67_ASAP7_75t_L g199 ( 
.A(n_159),
.Y(n_199)
);

NOR2xp33_ASAP7_75t_L g245 ( 
.A(n_199),
.B(n_216),
.Y(n_245)
);

AOI22xp5_ASAP7_75t_L g200 ( 
.A1(n_180),
.A2(n_139),
.B1(n_138),
.B2(n_114),
.Y(n_200)
);

AO22x2_ASAP7_75t_L g202 ( 
.A1(n_156),
.A2(n_153),
.B1(n_138),
.B2(n_114),
.Y(n_202)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_164),
.Y(n_204)
);

OA22x2_ASAP7_75t_L g206 ( 
.A1(n_176),
.A2(n_138),
.B1(n_116),
.B2(n_118),
.Y(n_206)
);

AOI22xp5_ASAP7_75t_L g209 ( 
.A1(n_156),
.A2(n_173),
.B1(n_192),
.B2(n_175),
.Y(n_209)
);

OAI22xp5_ASAP7_75t_SL g257 ( 
.A1(n_209),
.A2(n_218),
.B1(n_219),
.B2(n_221),
.Y(n_257)
);

NAND2x1p5_ASAP7_75t_L g210 ( 
.A(n_175),
.B(n_173),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_SL g243 ( 
.A(n_212),
.B(n_214),
.Y(n_243)
);

AO22x1_ASAP7_75t_SL g213 ( 
.A1(n_178),
.A2(n_129),
.B1(n_146),
.B2(n_116),
.Y(n_213)
);

NAND2xp5_ASAP7_75t_L g231 ( 
.A(n_213),
.B(n_222),
.Y(n_231)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_169),
.Y(n_214)
);

NOR2xp33_ASAP7_75t_L g216 ( 
.A(n_163),
.B(n_131),
.Y(n_216)
);

AOI22xp5_ASAP7_75t_L g219 ( 
.A1(n_173),
.A2(n_175),
.B1(n_188),
.B2(n_171),
.Y(n_219)
);

OAI22xp5_ASAP7_75t_L g221 ( 
.A1(n_165),
.A2(n_181),
.B1(n_168),
.B2(n_159),
.Y(n_221)
);

OR2x2_ASAP7_75t_L g222 ( 
.A(n_191),
.B(n_172),
.Y(n_222)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_167),
.Y(n_223)
);

NAND2xp5_ASAP7_75t_SL g250 ( 
.A(n_223),
.B(n_228),
.Y(n_250)
);

BUFx24_ASAP7_75t_SL g225 ( 
.A(n_161),
.Y(n_225)
);

CKINVDCx20_ASAP7_75t_R g235 ( 
.A(n_225),
.Y(n_235)
);

NOR2xp33_ASAP7_75t_L g227 ( 
.A(n_157),
.B(n_161),
.Y(n_227)
);

NOR2xp33_ASAP7_75t_L g253 ( 
.A(n_227),
.B(n_203),
.Y(n_253)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_182),
.Y(n_228)
);

NAND2xp33_ASAP7_75t_R g230 ( 
.A(n_210),
.B(n_172),
.Y(n_230)
);

OAI21xp5_ASAP7_75t_SL g283 ( 
.A1(n_230),
.A2(n_237),
.B(n_252),
.Y(n_283)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_201),
.Y(n_232)
);

NAND2xp5_ASAP7_75t_L g273 ( 
.A(n_232),
.B(n_233),
.Y(n_273)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_198),
.Y(n_233)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_198),
.Y(n_234)
);

NAND2xp5_ASAP7_75t_L g276 ( 
.A(n_234),
.B(n_247),
.Y(n_276)
);

CKINVDCx16_ASAP7_75t_R g236 ( 
.A(n_220),
.Y(n_236)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_236),
.Y(n_261)
);

INVx1_ASAP7_75t_SL g237 ( 
.A(n_206),
.Y(n_237)
);

MAJIxp5_ASAP7_75t_L g238 ( 
.A(n_207),
.B(n_183),
.C(n_186),
.Y(n_238)
);

MAJIxp5_ASAP7_75t_L g274 ( 
.A(n_238),
.B(n_222),
.C(n_195),
.Y(n_274)
);

NAND3xp33_ASAP7_75t_L g239 ( 
.A(n_210),
.B(n_170),
.C(n_157),
.Y(n_239)
);

AOI21xp33_ASAP7_75t_L g262 ( 
.A1(n_239),
.A2(n_258),
.B(n_259),
.Y(n_262)
);

OAI32xp33_ASAP7_75t_L g240 ( 
.A1(n_208),
.A2(n_168),
.A3(n_172),
.B1(n_184),
.B2(n_165),
.Y(n_240)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_240),
.Y(n_266)
);

CKINVDCx20_ASAP7_75t_R g241 ( 
.A(n_220),
.Y(n_241)
);

CKINVDCx20_ASAP7_75t_R g271 ( 
.A(n_241),
.Y(n_271)
);

INVx13_ASAP7_75t_L g244 ( 
.A(n_196),
.Y(n_244)
);

INVx2_ASAP7_75t_L g263 ( 
.A(n_244),
.Y(n_263)
);

CKINVDCx20_ASAP7_75t_R g246 ( 
.A(n_205),
.Y(n_246)
);

CKINVDCx20_ASAP7_75t_R g279 ( 
.A(n_246),
.Y(n_279)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_206),
.Y(n_247)
);

XOR2xp5_ASAP7_75t_L g249 ( 
.A(n_207),
.B(n_209),
.Y(n_249)
);

XOR2xp5_ASAP7_75t_L g264 ( 
.A(n_249),
.B(n_255),
.Y(n_264)
);

CKINVDCx20_ASAP7_75t_R g251 ( 
.A(n_205),
.Y(n_251)
);

NOR2xp33_ASAP7_75t_SL g265 ( 
.A(n_251),
.B(n_253),
.Y(n_265)
);

AOI21xp5_ASAP7_75t_L g252 ( 
.A1(n_215),
.A2(n_179),
.B(n_187),
.Y(n_252)
);

NAND2xp5_ASAP7_75t_SL g254 ( 
.A(n_223),
.B(n_158),
.Y(n_254)
);

OAI32xp33_ASAP7_75t_L g268 ( 
.A1(n_254),
.A2(n_214),
.A3(n_224),
.B1(n_202),
.B2(n_208),
.Y(n_268)
);

XOR2xp5_ASAP7_75t_L g255 ( 
.A(n_195),
.B(n_158),
.Y(n_255)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_206),
.Y(n_256)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_256),
.Y(n_272)
);

NOR2xp33_ASAP7_75t_L g258 ( 
.A(n_204),
.B(n_190),
.Y(n_258)
);

NOR2xp33_ASAP7_75t_L g259 ( 
.A(n_193),
.B(n_162),
.Y(n_259)
);

CKINVDCx16_ASAP7_75t_R g260 ( 
.A(n_203),
.Y(n_260)
);

OAI22xp5_ASAP7_75t_L g277 ( 
.A1(n_260),
.A2(n_224),
.B1(n_217),
.B2(n_202),
.Y(n_277)
);

AOI22xp5_ASAP7_75t_L g267 ( 
.A1(n_242),
.A2(n_202),
.B1(n_221),
.B2(n_215),
.Y(n_267)
);

OAI22xp5_ASAP7_75t_SL g288 ( 
.A1(n_267),
.A2(n_278),
.B1(n_231),
.B2(n_272),
.Y(n_288)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_268),
.Y(n_289)
);

XNOR2xp5_ASAP7_75t_L g269 ( 
.A(n_240),
.B(n_211),
.Y(n_269)
);

XOR2xp5_ASAP7_75t_L g293 ( 
.A(n_269),
.B(n_284),
.Y(n_293)
);

A2O1A1O1Ixp25_ASAP7_75t_L g270 ( 
.A1(n_230),
.A2(n_222),
.B(n_219),
.C(n_202),
.D(n_200),
.Y(n_270)
);

NAND3xp33_ASAP7_75t_L g305 ( 
.A(n_270),
.B(n_281),
.C(n_262),
.Y(n_305)
);

MAJIxp5_ASAP7_75t_L g299 ( 
.A(n_274),
.B(n_275),
.C(n_255),
.Y(n_299)
);

MAJIxp5_ASAP7_75t_L g275 ( 
.A(n_249),
.B(n_217),
.C(n_213),
.Y(n_275)
);

NAND2xp5_ASAP7_75t_L g294 ( 
.A(n_277),
.B(n_237),
.Y(n_294)
);

AOI22xp5_ASAP7_75t_L g278 ( 
.A1(n_242),
.A2(n_194),
.B1(n_213),
.B2(n_197),
.Y(n_278)
);

OAI22xp5_ASAP7_75t_L g280 ( 
.A1(n_237),
.A2(n_213),
.B1(n_206),
.B2(n_228),
.Y(n_280)
);

AOI22xp5_ASAP7_75t_L g306 ( 
.A1(n_280),
.A2(n_282),
.B1(n_250),
.B2(n_254),
.Y(n_306)
);

OA21x2_ASAP7_75t_SL g281 ( 
.A1(n_252),
.A2(n_162),
.B(n_174),
.Y(n_281)
);

OAI22xp5_ASAP7_75t_SL g282 ( 
.A1(n_247),
.A2(n_174),
.B1(n_189),
.B2(n_196),
.Y(n_282)
);

XNOR2xp5_ASAP7_75t_L g284 ( 
.A(n_248),
.B(n_185),
.Y(n_284)
);

AOI21xp5_ASAP7_75t_L g285 ( 
.A1(n_248),
.A2(n_196),
.B(n_185),
.Y(n_285)
);

OAI21xp5_ASAP7_75t_L g287 ( 
.A1(n_285),
.A2(n_256),
.B(n_231),
.Y(n_287)
);

INVx1_ASAP7_75t_SL g286 ( 
.A(n_273),
.Y(n_286)
);

NAND2xp5_ASAP7_75t_L g321 ( 
.A(n_286),
.B(n_290),
.Y(n_321)
);

OAI22xp5_ASAP7_75t_SL g312 ( 
.A1(n_287),
.A2(n_288),
.B1(n_294),
.B2(n_304),
.Y(n_312)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_276),
.Y(n_290)
);

NOR2xp33_ASAP7_75t_SL g291 ( 
.A(n_279),
.B(n_246),
.Y(n_291)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_291),
.Y(n_317)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_276),
.Y(n_292)
);

NOR2xp33_ASAP7_75t_L g314 ( 
.A(n_292),
.B(n_295),
.Y(n_314)
);

CKINVDCx20_ASAP7_75t_R g295 ( 
.A(n_279),
.Y(n_295)
);

XNOR2x2_ASAP7_75t_SL g296 ( 
.A(n_275),
.B(n_238),
.Y(n_296)
);

OAI322xp33_ASAP7_75t_L g313 ( 
.A1(n_296),
.A2(n_266),
.A3(n_270),
.B1(n_269),
.B2(n_284),
.C1(n_281),
.C2(n_285),
.Y(n_313)
);

CKINVDCx20_ASAP7_75t_R g297 ( 
.A(n_273),
.Y(n_297)
);

NOR2xp33_ASAP7_75t_L g324 ( 
.A(n_297),
.B(n_258),
.Y(n_324)
);

AND2x2_ASAP7_75t_L g298 ( 
.A(n_271),
.B(n_253),
.Y(n_298)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_298),
.Y(n_315)
);

MAJIxp5_ASAP7_75t_L g309 ( 
.A(n_299),
.B(n_300),
.C(n_301),
.Y(n_309)
);

MAJIxp5_ASAP7_75t_L g300 ( 
.A(n_264),
.B(n_257),
.C(n_233),
.Y(n_300)
);

MAJIxp5_ASAP7_75t_L g301 ( 
.A(n_264),
.B(n_257),
.C(n_234),
.Y(n_301)
);

MAJIxp5_ASAP7_75t_L g302 ( 
.A(n_274),
.B(n_260),
.C(n_241),
.Y(n_302)
);

MAJIxp5_ASAP7_75t_L g316 ( 
.A(n_302),
.B(n_283),
.C(n_261),
.Y(n_316)
);

NAND2xp5_ASAP7_75t_SL g303 ( 
.A(n_265),
.B(n_251),
.Y(n_303)
);

NAND2xp5_ASAP7_75t_SL g308 ( 
.A(n_303),
.B(n_305),
.Y(n_308)
);

OAI22xp5_ASAP7_75t_SL g304 ( 
.A1(n_278),
.A2(n_250),
.B1(n_229),
.B2(n_236),
.Y(n_304)
);

OAI22xp5_ASAP7_75t_L g311 ( 
.A1(n_306),
.A2(n_267),
.B1(n_266),
.B2(n_272),
.Y(n_311)
);

NAND2xp5_ASAP7_75t_L g307 ( 
.A(n_271),
.B(n_229),
.Y(n_307)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_307),
.Y(n_319)
);

INVxp67_ASAP7_75t_L g310 ( 
.A(n_298),
.Y(n_310)
);

NAND2xp5_ASAP7_75t_L g335 ( 
.A(n_310),
.B(n_323),
.Y(n_335)
);

AOI22xp5_ASAP7_75t_L g334 ( 
.A1(n_311),
.A2(n_289),
.B1(n_290),
.B2(n_292),
.Y(n_334)
);

XNOR2xp5_ASAP7_75t_L g327 ( 
.A(n_313),
.B(n_293),
.Y(n_327)
);

MAJIxp5_ASAP7_75t_L g330 ( 
.A(n_316),
.B(n_318),
.C(n_320),
.Y(n_330)
);

MAJIxp5_ASAP7_75t_L g318 ( 
.A(n_299),
.B(n_283),
.C(n_261),
.Y(n_318)
);

MAJIxp5_ASAP7_75t_L g320 ( 
.A(n_300),
.B(n_232),
.C(n_245),
.Y(n_320)
);

MAJIxp5_ASAP7_75t_L g322 ( 
.A(n_301),
.B(n_245),
.C(n_265),
.Y(n_322)
);

MAJIxp5_ASAP7_75t_L g338 ( 
.A(n_322),
.B(n_325),
.C(n_307),
.Y(n_338)
);

INVx1_ASAP7_75t_SL g323 ( 
.A(n_298),
.Y(n_323)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_324),
.Y(n_337)
);

MAJIxp5_ASAP7_75t_L g325 ( 
.A(n_302),
.B(n_243),
.C(n_259),
.Y(n_325)
);

NOR2xp33_ASAP7_75t_L g326 ( 
.A(n_291),
.B(n_263),
.Y(n_326)
);

NAND2xp5_ASAP7_75t_SL g328 ( 
.A(n_326),
.B(n_295),
.Y(n_328)
);

NAND2xp5_ASAP7_75t_SL g344 ( 
.A(n_327),
.B(n_331),
.Y(n_344)
);

INVx1_ASAP7_75t_L g351 ( 
.A(n_328),
.Y(n_351)
);

AOI22xp5_ASAP7_75t_SL g329 ( 
.A1(n_312),
.A2(n_288),
.B1(n_304),
.B2(n_289),
.Y(n_329)
);

AOI22xp5_ASAP7_75t_SL g345 ( 
.A1(n_329),
.A2(n_333),
.B1(n_315),
.B2(n_287),
.Y(n_345)
);

XNOR2xp5_ASAP7_75t_L g331 ( 
.A(n_309),
.B(n_293),
.Y(n_331)
);

BUFx24_ASAP7_75t_SL g332 ( 
.A(n_308),
.Y(n_332)
);

NAND2xp5_ASAP7_75t_L g349 ( 
.A(n_332),
.B(n_338),
.Y(n_349)
);

AND2x4_ASAP7_75t_L g333 ( 
.A(n_323),
.B(n_286),
.Y(n_333)
);

NOR2xp33_ASAP7_75t_L g346 ( 
.A(n_334),
.B(n_336),
.Y(n_346)
);

AOI22xp5_ASAP7_75t_L g336 ( 
.A1(n_312),
.A2(n_297),
.B1(n_282),
.B2(n_243),
.Y(n_336)
);

AOI22xp5_ASAP7_75t_L g339 ( 
.A1(n_310),
.A2(n_306),
.B1(n_296),
.B2(n_294),
.Y(n_339)
);

INVxp67_ASAP7_75t_L g343 ( 
.A(n_339),
.Y(n_343)
);

NOR2xp33_ASAP7_75t_L g340 ( 
.A(n_317),
.B(n_263),
.Y(n_340)
);

CKINVDCx20_ASAP7_75t_R g352 ( 
.A(n_340),
.Y(n_352)
);

NOR2xp33_ASAP7_75t_L g341 ( 
.A(n_325),
.B(n_226),
.Y(n_341)
);

OAI21xp5_ASAP7_75t_SL g350 ( 
.A1(n_341),
.A2(n_321),
.B(n_318),
.Y(n_350)
);

AOI22xp5_ASAP7_75t_L g342 ( 
.A1(n_333),
.A2(n_315),
.B1(n_319),
.B2(n_314),
.Y(n_342)
);

NAND2xp5_ASAP7_75t_L g358 ( 
.A(n_342),
.B(n_345),
.Y(n_358)
);

XOR2xp5_ASAP7_75t_L g347 ( 
.A(n_330),
.B(n_309),
.Y(n_347)
);

XOR2xp5_ASAP7_75t_L g354 ( 
.A(n_347),
.B(n_333),
.Y(n_354)
);

MAJIxp5_ASAP7_75t_L g348 ( 
.A(n_338),
.B(n_320),
.C(n_322),
.Y(n_348)
);

NAND2xp5_ASAP7_75t_L g361 ( 
.A(n_348),
.B(n_353),
.Y(n_361)
);

AOI21xp5_ASAP7_75t_L g356 ( 
.A1(n_350),
.A2(n_337),
.B(n_335),
.Y(n_356)
);

MAJIxp5_ASAP7_75t_L g353 ( 
.A(n_330),
.B(n_316),
.C(n_321),
.Y(n_353)
);

XNOR2xp5_ASAP7_75t_L g366 ( 
.A(n_354),
.B(n_355),
.Y(n_366)
);

MAJx2_ASAP7_75t_L g355 ( 
.A(n_353),
.B(n_348),
.C(n_343),
.Y(n_355)
);

INVx1_ASAP7_75t_L g370 ( 
.A(n_356),
.Y(n_370)
);

BUFx4f_ASAP7_75t_SL g357 ( 
.A(n_352),
.Y(n_357)
);

CKINVDCx20_ASAP7_75t_R g367 ( 
.A(n_357),
.Y(n_367)
);

MAJIxp5_ASAP7_75t_L g359 ( 
.A(n_347),
.B(n_329),
.C(n_235),
.Y(n_359)
);

NAND2xp5_ASAP7_75t_L g364 ( 
.A(n_359),
.B(n_362),
.Y(n_364)
);

AOI21xp5_ASAP7_75t_L g360 ( 
.A1(n_343),
.A2(n_268),
.B(n_244),
.Y(n_360)
);

OAI21xp5_ASAP7_75t_L g365 ( 
.A1(n_360),
.A2(n_363),
.B(n_346),
.Y(n_365)
);

NOR2xp33_ASAP7_75t_SL g362 ( 
.A(n_351),
.B(n_235),
.Y(n_362)
);

NOR2xp33_ASAP7_75t_SL g363 ( 
.A(n_349),
.B(n_226),
.Y(n_363)
);

AOI21xp5_ASAP7_75t_L g372 ( 
.A1(n_365),
.A2(n_368),
.B(n_160),
.Y(n_372)
);

A2O1A1Ixp33_ASAP7_75t_SL g368 ( 
.A1(n_358),
.A2(n_345),
.B(n_342),
.C(n_244),
.Y(n_368)
);

MAJIxp5_ASAP7_75t_L g369 ( 
.A(n_355),
.B(n_344),
.C(n_160),
.Y(n_369)
);

AND2x2_ASAP7_75t_L g374 ( 
.A(n_369),
.B(n_226),
.Y(n_374)
);

AOI31xp67_ASAP7_75t_L g371 ( 
.A1(n_364),
.A2(n_357),
.A3(n_361),
.B(n_354),
.Y(n_371)
);

AOI21xp5_ASAP7_75t_L g376 ( 
.A1(n_371),
.A2(n_374),
.B(n_367),
.Y(n_376)
);

NOR2xp33_ASAP7_75t_L g375 ( 
.A(n_372),
.B(n_373),
.Y(n_375)
);

XNOR2xp5_ASAP7_75t_L g373 ( 
.A(n_369),
.B(n_160),
.Y(n_373)
);

NOR2xp33_ASAP7_75t_SL g377 ( 
.A(n_376),
.B(n_366),
.Y(n_377)
);

AOI21xp5_ASAP7_75t_L g378 ( 
.A1(n_377),
.A2(n_370),
.B(n_375),
.Y(n_378)
);

OAI21xp5_ASAP7_75t_L g379 ( 
.A1(n_378),
.A2(n_368),
.B(n_226),
.Y(n_379)
);

XNOR2xp5_ASAP7_75t_L g380 ( 
.A(n_379),
.B(n_368),
.Y(n_380)
);


endmodule