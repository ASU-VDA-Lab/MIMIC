module real_jpeg_12513_n_18 (n_17, n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_16, n_3, n_10, n_9, n_18);

input n_17;
input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_16;
input n_3;
input n_10;
input n_9;

output n_18;

wire n_37;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_300;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_199;
wire n_95;
wire n_238;
wire n_67;
wire n_235;
wire n_107;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_123;
wire n_50;
wire n_186;
wire n_137;
wire n_72;
wire n_171;
wire n_151;
wire n_272;
wire n_198;
wire n_203;
wire n_23;
wire n_71;
wire n_61;
wire n_99;
wire n_80;
wire n_30;
wire n_149;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_230;
wire n_128;
wire n_202;
wire n_216;
wire n_127;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_252;
wire n_310;
wire n_83;
wire n_78;
wire n_288;
wire n_221;
wire n_104;
wire n_153;
wire n_131;
wire n_87;
wire n_40;
wire n_98;
wire n_200;
wire n_214;
wire n_113;
wire n_251;
wire n_139;
wire n_33;
wire n_175;
wire n_156;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_77;
wire n_219;
wire n_122;
wire n_19;
wire n_262;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_20;
wire n_314;
wire n_278;
wire n_103;
wire n_232;
wire n_212;
wire n_284;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_213;
wire n_25;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_49;
wire n_68;
wire n_146;
wire n_286;
wire n_166;
wire n_176;
wire n_215;
wire n_312;
wire n_316;
wire n_307;
wire n_161;
wire n_207;
wire n_237;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_140;
wire n_126;
wire n_120;
wire n_155;
wire n_319;
wire n_93;
wire n_242;
wire n_142;
wire n_76;
wire n_79;
wire n_282;
wire n_147;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_145;
wire n_266;
wire n_109;
wire n_148;
wire n_196;
wire n_298;
wire n_152;
wire n_270;
wire n_159;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_258;
wire n_150;
wire n_41;
wire n_74;
wire n_158;
wire n_204;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_75;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_119;
wire n_283;
wire n_181;
wire n_256;
wire n_253;
wire n_273;
wire n_54;
wire n_168;
wire n_38;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_292;
wire n_64;
wire n_291;
wire n_236;
wire n_276;
wire n_287;
wire n_174;
wire n_255;
wire n_299;
wire n_243;
wire n_56;
wire n_293;
wire n_275;
wire n_227;
wire n_229;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_45;
wire n_268;
wire n_42;
wire n_313;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_143;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_303;
wire n_321;
wire n_100;
wire n_51;
wire n_205;
wire n_261;
wire n_86;
wire n_70;
wire n_32;
wire n_228;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_133;
wire n_257;
wire n_210;
wire n_206;
wire n_85;
wire n_96;
wire n_308;

BUFx12f_ASAP7_75t_L g98 ( 
.A(n_0),
.Y(n_98)
);

BUFx16f_ASAP7_75t_L g47 ( 
.A(n_1),
.Y(n_47)
);

BUFx12_ASAP7_75t_L g60 ( 
.A(n_2),
.Y(n_60)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_3),
.Y(n_190)
);

AOI21xp33_ASAP7_75t_L g208 ( 
.A1(n_3),
.A2(n_59),
.B(n_209),
.Y(n_208)
);

NAND2xp5_ASAP7_75t_L g224 ( 
.A(n_3),
.B(n_81),
.Y(n_224)
);

OAI22xp33_ASAP7_75t_L g260 ( 
.A1(n_3),
.A2(n_34),
.B1(n_35),
.B2(n_190),
.Y(n_260)
);

O2A1O1Ixp33_ASAP7_75t_L g262 ( 
.A1(n_3),
.A2(n_35),
.B(n_47),
.C(n_263),
.Y(n_262)
);

NAND2xp5_ASAP7_75t_SL g266 ( 
.A(n_3),
.B(n_72),
.Y(n_266)
);

NAND2xp5_ASAP7_75t_L g284 ( 
.A(n_3),
.B(n_98),
.Y(n_284)
);

NAND2xp5_ASAP7_75t_L g287 ( 
.A(n_3),
.B(n_41),
.Y(n_287)
);

A2O1A1Ixp33_ASAP7_75t_L g296 ( 
.A1(n_3),
.A2(n_27),
.B(n_29),
.C(n_297),
.Y(n_296)
);

AOI22xp33_ASAP7_75t_L g197 ( 
.A1(n_4),
.A2(n_59),
.B1(n_60),
.B2(n_198),
.Y(n_197)
);

CKINVDCx20_ASAP7_75t_R g198 ( 
.A(n_4),
.Y(n_198)
);

AOI22xp33_ASAP7_75t_SL g222 ( 
.A1(n_4),
.A2(n_29),
.B1(n_30),
.B2(n_198),
.Y(n_222)
);

OAI22xp5_ASAP7_75t_L g261 ( 
.A1(n_4),
.A2(n_34),
.B1(n_35),
.B2(n_198),
.Y(n_261)
);

OAI22xp33_ASAP7_75t_SL g282 ( 
.A1(n_4),
.A2(n_43),
.B1(n_48),
.B2(n_198),
.Y(n_282)
);

BUFx16f_ASAP7_75t_L g34 ( 
.A(n_5),
.Y(n_34)
);

AOI22xp33_ASAP7_75t_SL g170 ( 
.A1(n_6),
.A2(n_59),
.B1(n_60),
.B2(n_171),
.Y(n_170)
);

CKINVDCx20_ASAP7_75t_R g171 ( 
.A(n_6),
.Y(n_171)
);

AOI22xp33_ASAP7_75t_SL g212 ( 
.A1(n_6),
.A2(n_29),
.B1(n_30),
.B2(n_171),
.Y(n_212)
);

OAI22xp5_ASAP7_75t_L g268 ( 
.A1(n_6),
.A2(n_34),
.B1(n_35),
.B2(n_171),
.Y(n_268)
);

OAI22xp33_ASAP7_75t_SL g275 ( 
.A1(n_6),
.A2(n_43),
.B1(n_48),
.B2(n_171),
.Y(n_275)
);

BUFx12f_ASAP7_75t_L g30 ( 
.A(n_7),
.Y(n_30)
);

AOI22xp33_ASAP7_75t_L g36 ( 
.A1(n_8),
.A2(n_29),
.B1(n_30),
.B2(n_37),
.Y(n_36)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_8),
.Y(n_37)
);

OAI22xp5_ASAP7_75t_L g80 ( 
.A1(n_8),
.A2(n_37),
.B1(n_59),
.B2(n_60),
.Y(n_80)
);

OAI22xp5_ASAP7_75t_L g103 ( 
.A1(n_8),
.A2(n_34),
.B1(n_35),
.B2(n_37),
.Y(n_103)
);

AOI22xp33_ASAP7_75t_L g134 ( 
.A1(n_8),
.A2(n_37),
.B1(n_43),
.B2(n_48),
.Y(n_134)
);

BUFx12_ASAP7_75t_L g31 ( 
.A(n_9),
.Y(n_31)
);

AOI22xp33_ASAP7_75t_SL g66 ( 
.A1(n_10),
.A2(n_59),
.B1(n_60),
.B2(n_67),
.Y(n_66)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_10),
.Y(n_67)
);

AOI22xp33_ASAP7_75t_SL g140 ( 
.A1(n_10),
.A2(n_29),
.B1(n_30),
.B2(n_67),
.Y(n_140)
);

OAI22xp5_ASAP7_75t_L g165 ( 
.A1(n_10),
.A2(n_34),
.B1(n_35),
.B2(n_67),
.Y(n_165)
);

OAI22xp5_ASAP7_75t_L g226 ( 
.A1(n_10),
.A2(n_43),
.B1(n_48),
.B2(n_67),
.Y(n_226)
);

AOI22xp33_ASAP7_75t_SL g38 ( 
.A1(n_11),
.A2(n_29),
.B1(n_30),
.B2(n_39),
.Y(n_38)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_11),
.Y(n_39)
);

OAI22xp5_ASAP7_75t_SL g51 ( 
.A1(n_11),
.A2(n_34),
.B1(n_35),
.B2(n_39),
.Y(n_51)
);

OAI22xp5_ASAP7_75t_L g99 ( 
.A1(n_11),
.A2(n_39),
.B1(n_43),
.B2(n_48),
.Y(n_99)
);

BUFx8_ASAP7_75t_L g57 ( 
.A(n_12),
.Y(n_57)
);

AOI22xp33_ASAP7_75t_SL g105 ( 
.A1(n_13),
.A2(n_59),
.B1(n_60),
.B2(n_106),
.Y(n_105)
);

CKINVDCx20_ASAP7_75t_R g106 ( 
.A(n_13),
.Y(n_106)
);

AOI22xp33_ASAP7_75t_SL g168 ( 
.A1(n_13),
.A2(n_29),
.B1(n_30),
.B2(n_106),
.Y(n_168)
);

OAI22xp5_ASAP7_75t_L g214 ( 
.A1(n_13),
.A2(n_34),
.B1(n_35),
.B2(n_106),
.Y(n_214)
);

OAI22xp5_ASAP7_75t_SL g249 ( 
.A1(n_13),
.A2(n_43),
.B1(n_48),
.B2(n_106),
.Y(n_249)
);

AOI22xp33_ASAP7_75t_SL g142 ( 
.A1(n_14),
.A2(n_59),
.B1(n_60),
.B2(n_143),
.Y(n_142)
);

CKINVDCx20_ASAP7_75t_R g143 ( 
.A(n_14),
.Y(n_143)
);

AOI22xp33_ASAP7_75t_SL g193 ( 
.A1(n_14),
.A2(n_29),
.B1(n_30),
.B2(n_143),
.Y(n_193)
);

AOI22xp33_ASAP7_75t_SL g241 ( 
.A1(n_14),
.A2(n_34),
.B1(n_35),
.B2(n_143),
.Y(n_241)
);

OAI22xp5_ASAP7_75t_SL g270 ( 
.A1(n_14),
.A2(n_43),
.B1(n_48),
.B2(n_143),
.Y(n_270)
);

AOI22xp33_ASAP7_75t_SL g63 ( 
.A1(n_15),
.A2(n_59),
.B1(n_60),
.B2(n_64),
.Y(n_63)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_15),
.Y(n_64)
);

OAI22xp5_ASAP7_75t_L g70 ( 
.A1(n_15),
.A2(n_29),
.B1(n_30),
.B2(n_64),
.Y(n_70)
);

OAI22xp5_ASAP7_75t_L g102 ( 
.A1(n_15),
.A2(n_34),
.B1(n_35),
.B2(n_64),
.Y(n_102)
);

OAI22xp5_ASAP7_75t_L g162 ( 
.A1(n_15),
.A2(n_43),
.B1(n_48),
.B2(n_64),
.Y(n_162)
);

INVx11_ASAP7_75t_L g45 ( 
.A(n_16),
.Y(n_45)
);

AOI22xp33_ASAP7_75t_SL g61 ( 
.A1(n_17),
.A2(n_59),
.B1(n_60),
.B2(n_62),
.Y(n_61)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_17),
.Y(n_62)
);

AOI22xp33_ASAP7_75t_SL g111 ( 
.A1(n_17),
.A2(n_29),
.B1(n_30),
.B2(n_62),
.Y(n_111)
);

AOI22xp33_ASAP7_75t_L g138 ( 
.A1(n_17),
.A2(n_34),
.B1(n_35),
.B2(n_62),
.Y(n_138)
);

OAI22xp5_ASAP7_75t_L g186 ( 
.A1(n_17),
.A2(n_43),
.B1(n_48),
.B2(n_62),
.Y(n_186)
);

XOR2xp5_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_87),
.Y(n_18)
);

NAND2xp5_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_85),
.Y(n_19)
);

NAND2xp5_ASAP7_75t_SL g20 ( 
.A(n_21),
.B(n_73),
.Y(n_20)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_21),
.B(n_73),
.Y(n_86)
);

MAJIxp5_ASAP7_75t_L g21 ( 
.A(n_22),
.B(n_65),
.C(n_68),
.Y(n_21)
);

AOI22xp5_ASAP7_75t_SL g147 ( 
.A1(n_22),
.A2(n_65),
.B1(n_114),
.B2(n_148),
.Y(n_147)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_22),
.Y(n_148)
);

XNOR2xp5_ASAP7_75t_L g22 ( 
.A(n_23),
.B(n_53),
.Y(n_22)
);

AOI22xp5_ASAP7_75t_L g23 ( 
.A1(n_24),
.A2(n_25),
.B1(n_40),
.B2(n_52),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_25),
.Y(n_24)
);

MAJIxp5_ASAP7_75t_L g84 ( 
.A(n_25),
.B(n_40),
.C(n_53),
.Y(n_84)
);

OAI22xp5_ASAP7_75t_SL g25 ( 
.A1(n_26),
.A2(n_33),
.B1(n_36),
.B2(n_38),
.Y(n_25)
);

OAI22xp5_ASAP7_75t_SL g139 ( 
.A1(n_26),
.A2(n_33),
.B1(n_111),
.B2(n_140),
.Y(n_139)
);

OAI22xp5_ASAP7_75t_SL g167 ( 
.A1(n_26),
.A2(n_33),
.B1(n_140),
.B2(n_168),
.Y(n_167)
);

OAI22xp5_ASAP7_75t_SL g211 ( 
.A1(n_26),
.A2(n_33),
.B1(n_193),
.B2(n_212),
.Y(n_211)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_27),
.Y(n_26)
);

AOI22xp5_ASAP7_75t_SL g69 ( 
.A1(n_27),
.A2(n_70),
.B1(n_71),
.B2(n_72),
.Y(n_69)
);

OAI21xp5_ASAP7_75t_SL g75 ( 
.A1(n_27),
.A2(n_72),
.B(n_76),
.Y(n_75)
);

AOI22xp5_ASAP7_75t_L g109 ( 
.A1(n_27),
.A2(n_70),
.B1(n_72),
.B2(n_110),
.Y(n_109)
);

AOI22xp5_ASAP7_75t_L g191 ( 
.A1(n_27),
.A2(n_72),
.B1(n_192),
.B2(n_194),
.Y(n_191)
);

AOI22xp5_ASAP7_75t_L g220 ( 
.A1(n_27),
.A2(n_72),
.B1(n_221),
.B2(n_223),
.Y(n_220)
);

AND2x2_ASAP7_75t_L g27 ( 
.A(n_28),
.B(n_33),
.Y(n_27)
);

OAI22xp5_ASAP7_75t_SL g28 ( 
.A1(n_29),
.A2(n_30),
.B1(n_31),
.B2(n_32),
.Y(n_28)
);

OA22x2_ASAP7_75t_L g55 ( 
.A1(n_29),
.A2(n_30),
.B1(n_56),
.B2(n_57),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g188 ( 
.A(n_29),
.B(n_56),
.Y(n_188)
);

OAI32xp33_ASAP7_75t_L g245 ( 
.A1(n_29),
.A2(n_31),
.A3(n_34),
.B1(n_246),
.B2(n_247),
.Y(n_245)
);

INVx5_ASAP7_75t_L g29 ( 
.A(n_30),
.Y(n_29)
);

OAI32xp33_ASAP7_75t_L g187 ( 
.A1(n_30),
.A2(n_57),
.A3(n_59),
.B1(n_188),
.B2(n_189),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_SL g246 ( 
.A(n_30),
.B(n_190),
.Y(n_246)
);

INVx8_ASAP7_75t_L g32 ( 
.A(n_31),
.Y(n_32)
);

OA22x2_ASAP7_75t_L g33 ( 
.A1(n_31),
.A2(n_32),
.B1(n_34),
.B2(n_35),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_L g247 ( 
.A(n_32),
.B(n_35),
.Y(n_247)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_33),
.Y(n_72)
);

OAI21xp5_ASAP7_75t_L g295 ( 
.A1(n_33),
.A2(n_222),
.B(n_296),
.Y(n_295)
);

INVx5_ASAP7_75t_L g35 ( 
.A(n_34),
.Y(n_35)
);

OAI22xp5_ASAP7_75t_L g50 ( 
.A1(n_34),
.A2(n_35),
.B1(n_46),
.B2(n_47),
.Y(n_50)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_36),
.Y(n_71)
);

CKINVDCx16_ASAP7_75t_R g76 ( 
.A(n_38),
.Y(n_76)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_40),
.Y(n_52)
);

MAJIxp5_ASAP7_75t_L g68 ( 
.A(n_40),
.B(n_65),
.C(n_69),
.Y(n_68)
);

OAI22xp5_ASAP7_75t_SL g116 ( 
.A1(n_40),
.A2(n_52),
.B1(n_69),
.B2(n_117),
.Y(n_116)
);

OAI21xp5_ASAP7_75t_L g40 ( 
.A1(n_41),
.A2(n_49),
.B(n_51),
.Y(n_40)
);

AOI22xp5_ASAP7_75t_L g101 ( 
.A1(n_41),
.A2(n_49),
.B1(n_102),
.B2(n_103),
.Y(n_101)
);

AOI22xp5_ASAP7_75t_L g112 ( 
.A1(n_41),
.A2(n_49),
.B1(n_51),
.B2(n_103),
.Y(n_112)
);

AOI22xp5_ASAP7_75t_L g136 ( 
.A1(n_41),
.A2(n_49),
.B1(n_102),
.B2(n_137),
.Y(n_136)
);

AOI22xp5_ASAP7_75t_L g213 ( 
.A1(n_41),
.A2(n_49),
.B1(n_165),
.B2(n_214),
.Y(n_213)
);

AOI22xp5_ASAP7_75t_L g239 ( 
.A1(n_41),
.A2(n_49),
.B1(n_214),
.B2(n_240),
.Y(n_239)
);

AOI22xp5_ASAP7_75t_L g259 ( 
.A1(n_41),
.A2(n_49),
.B1(n_260),
.B2(n_261),
.Y(n_259)
);

AOI22xp5_ASAP7_75t_L g267 ( 
.A1(n_41),
.A2(n_49),
.B1(n_261),
.B2(n_268),
.Y(n_267)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_42),
.Y(n_41)
);

AND2x2_ASAP7_75t_L g49 ( 
.A(n_42),
.B(n_50),
.Y(n_49)
);

OAI22xp5_ASAP7_75t_L g163 ( 
.A1(n_42),
.A2(n_138),
.B1(n_164),
.B2(n_166),
.Y(n_163)
);

OAI22xp5_ASAP7_75t_SL g298 ( 
.A1(n_42),
.A2(n_166),
.B1(n_241),
.B2(n_299),
.Y(n_298)
);

OA22x2_ASAP7_75t_L g42 ( 
.A1(n_43),
.A2(n_46),
.B1(n_47),
.B2(n_48),
.Y(n_42)
);

INVx6_ASAP7_75t_L g48 ( 
.A(n_43),
.Y(n_48)
);

AND2x2_ASAP7_75t_L g96 ( 
.A(n_43),
.B(n_97),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_SL g283 ( 
.A(n_43),
.B(n_284),
.Y(n_283)
);

BUFx12f_ASAP7_75t_L g43 ( 
.A(n_44),
.Y(n_43)
);

INVx8_ASAP7_75t_L g44 ( 
.A(n_45),
.Y(n_44)
);

OAI21xp33_ASAP7_75t_L g263 ( 
.A1(n_46),
.A2(n_48),
.B(n_190),
.Y(n_263)
);

INVx6_ASAP7_75t_L g46 ( 
.A(n_47),
.Y(n_46)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_49),
.Y(n_166)
);

OAI22xp5_ASAP7_75t_SL g53 ( 
.A1(n_54),
.A2(n_55),
.B1(n_61),
.B2(n_63),
.Y(n_53)
);

OAI22xp5_ASAP7_75t_L g65 ( 
.A1(n_54),
.A2(n_55),
.B1(n_61),
.B2(n_66),
.Y(n_65)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_54),
.Y(n_79)
);

OAI22xp5_ASAP7_75t_SL g104 ( 
.A1(n_54),
.A2(n_55),
.B1(n_66),
.B2(n_105),
.Y(n_104)
);

OAI22xp5_ASAP7_75t_SL g141 ( 
.A1(n_54),
.A2(n_55),
.B1(n_105),
.B2(n_142),
.Y(n_141)
);

OAI22xp5_ASAP7_75t_SL g169 ( 
.A1(n_54),
.A2(n_55),
.B1(n_142),
.B2(n_170),
.Y(n_169)
);

OAI22xp5_ASAP7_75t_SL g207 ( 
.A1(n_54),
.A2(n_55),
.B1(n_197),
.B2(n_208),
.Y(n_207)
);

NAND2xp5_ASAP7_75t_SL g54 ( 
.A(n_55),
.B(n_58),
.Y(n_54)
);

CKINVDCx14_ASAP7_75t_R g81 ( 
.A(n_55),
.Y(n_81)
);

OAI22xp5_ASAP7_75t_SL g58 ( 
.A1(n_56),
.A2(n_57),
.B1(n_59),
.B2(n_60),
.Y(n_58)
);

INVx11_ASAP7_75t_L g56 ( 
.A(n_57),
.Y(n_56)
);

INVx4_ASAP7_75t_L g59 ( 
.A(n_60),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_SL g189 ( 
.A(n_60),
.B(n_190),
.Y(n_189)
);

CKINVDCx20_ASAP7_75t_R g78 ( 
.A(n_63),
.Y(n_78)
);

AOI22xp5_ASAP7_75t_L g113 ( 
.A1(n_65),
.A2(n_114),
.B1(n_115),
.B2(n_116),
.Y(n_113)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_65),
.Y(n_114)
);

XNOR2xp5_ASAP7_75t_L g146 ( 
.A(n_68),
.B(n_147),
.Y(n_146)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_69),
.Y(n_117)
);

XNOR2xp5_ASAP7_75t_L g73 ( 
.A(n_74),
.B(n_84),
.Y(n_73)
);

AOI22xp5_ASAP7_75t_L g74 ( 
.A1(n_75),
.A2(n_77),
.B1(n_82),
.B2(n_83),
.Y(n_74)
);

CKINVDCx20_ASAP7_75t_R g82 ( 
.A(n_75),
.Y(n_82)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_77),
.Y(n_83)
);

AOI22xp5_ASAP7_75t_L g77 ( 
.A1(n_78),
.A2(n_79),
.B1(n_80),
.B2(n_81),
.Y(n_77)
);

AOI22xp5_ASAP7_75t_L g195 ( 
.A1(n_79),
.A2(n_81),
.B1(n_196),
.B2(n_199),
.Y(n_195)
);

INVxp67_ASAP7_75t_L g85 ( 
.A(n_86),
.Y(n_85)
);

AO21x1_ASAP7_75t_L g87 ( 
.A1(n_88),
.A2(n_149),
.B(n_319),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_89),
.B(n_144),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_SL g89 ( 
.A(n_90),
.B(n_120),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g320 ( 
.A(n_90),
.B(n_120),
.Y(n_320)
);

XOR2xp5_ASAP7_75t_L g90 ( 
.A(n_91),
.B(n_107),
.Y(n_90)
);

MAJIxp5_ASAP7_75t_L g145 ( 
.A(n_91),
.B(n_113),
.C(n_118),
.Y(n_145)
);

OAI21xp5_ASAP7_75t_L g91 ( 
.A1(n_92),
.A2(n_95),
.B(n_104),
.Y(n_91)
);

OAI22xp5_ASAP7_75t_L g122 ( 
.A1(n_92),
.A2(n_93),
.B1(n_123),
.B2(n_124),
.Y(n_122)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_93),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_L g93 ( 
.A(n_94),
.B(n_100),
.Y(n_93)
);

AOI22xp5_ASAP7_75t_L g124 ( 
.A1(n_94),
.A2(n_95),
.B1(n_104),
.B2(n_125),
.Y(n_124)
);

AOI22xp5_ASAP7_75t_L g155 ( 
.A1(n_94),
.A2(n_95),
.B1(n_100),
.B2(n_101),
.Y(n_155)
);

CKINVDCx16_ASAP7_75t_R g94 ( 
.A(n_95),
.Y(n_94)
);

OAI21xp5_ASAP7_75t_SL g95 ( 
.A1(n_96),
.A2(n_98),
.B(n_99),
.Y(n_95)
);

AOI22xp5_ASAP7_75t_L g132 ( 
.A1(n_96),
.A2(n_98),
.B1(n_99),
.B2(n_133),
.Y(n_132)
);

CKINVDCx16_ASAP7_75t_R g160 ( 
.A(n_96),
.Y(n_160)
);

AOI22xp5_ASAP7_75t_L g185 ( 
.A1(n_96),
.A2(n_98),
.B1(n_162),
.B2(n_186),
.Y(n_185)
);

AOI22xp5_ASAP7_75t_L g225 ( 
.A1(n_96),
.A2(n_98),
.B1(n_186),
.B2(n_226),
.Y(n_225)
);

AOI22xp5_ASAP7_75t_L g248 ( 
.A1(n_96),
.A2(n_98),
.B1(n_226),
.B2(n_249),
.Y(n_248)
);

AOI22xp5_ASAP7_75t_SL g269 ( 
.A1(n_96),
.A2(n_98),
.B1(n_249),
.B2(n_270),
.Y(n_269)
);

AOI22xp5_ASAP7_75t_SL g281 ( 
.A1(n_96),
.A2(n_98),
.B1(n_190),
.B2(n_282),
.Y(n_281)
);

AOI22xp33_ASAP7_75t_L g286 ( 
.A1(n_96),
.A2(n_98),
.B1(n_275),
.B2(n_282),
.Y(n_286)
);

OAI22xp5_ASAP7_75t_L g159 ( 
.A1(n_97),
.A2(n_134),
.B1(n_160),
.B2(n_161),
.Y(n_159)
);

OAI22xp5_ASAP7_75t_SL g273 ( 
.A1(n_97),
.A2(n_160),
.B1(n_274),
.B2(n_276),
.Y(n_273)
);

INVx4_ASAP7_75t_L g97 ( 
.A(n_98),
.Y(n_97)
);

CKINVDCx20_ASAP7_75t_R g100 ( 
.A(n_101),
.Y(n_100)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_104),
.Y(n_125)
);

AOI22xp5_ASAP7_75t_L g107 ( 
.A1(n_108),
.A2(n_113),
.B1(n_118),
.B2(n_119),
.Y(n_107)
);

CKINVDCx20_ASAP7_75t_R g118 ( 
.A(n_108),
.Y(n_118)
);

OAI21xp33_ASAP7_75t_L g127 ( 
.A1(n_108),
.A2(n_109),
.B(n_112),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_L g108 ( 
.A(n_109),
.B(n_112),
.Y(n_108)
);

INVxp67_ASAP7_75t_L g110 ( 
.A(n_111),
.Y(n_110)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_113),
.Y(n_119)
);

CKINVDCx16_ASAP7_75t_R g115 ( 
.A(n_116),
.Y(n_115)
);

MAJIxp5_ASAP7_75t_L g120 ( 
.A(n_121),
.B(n_126),
.C(n_128),
.Y(n_120)
);

AOI22xp5_ASAP7_75t_L g173 ( 
.A1(n_121),
.A2(n_122),
.B1(n_126),
.B2(n_127),
.Y(n_173)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_122),
.Y(n_121)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_124),
.Y(n_123)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_127),
.Y(n_126)
);

XOR2xp5_ASAP7_75t_L g172 ( 
.A(n_128),
.B(n_173),
.Y(n_172)
);

MAJIxp5_ASAP7_75t_L g128 ( 
.A(n_129),
.B(n_139),
.C(n_141),
.Y(n_128)
);

AOI22xp5_ASAP7_75t_L g152 ( 
.A1(n_129),
.A2(n_130),
.B1(n_153),
.B2(n_154),
.Y(n_152)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_130),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_L g130 ( 
.A(n_131),
.B(n_135),
.Y(n_130)
);

OAI22xp5_ASAP7_75t_SL g181 ( 
.A1(n_131),
.A2(n_132),
.B1(n_135),
.B2(n_136),
.Y(n_181)
);

CKINVDCx20_ASAP7_75t_R g131 ( 
.A(n_132),
.Y(n_131)
);

INVxp67_ASAP7_75t_L g133 ( 
.A(n_134),
.Y(n_133)
);

CKINVDCx14_ASAP7_75t_R g135 ( 
.A(n_136),
.Y(n_135)
);

INVxp67_ASAP7_75t_L g137 ( 
.A(n_138),
.Y(n_137)
);

XOR2xp5_ASAP7_75t_L g154 ( 
.A(n_139),
.B(n_141),
.Y(n_154)
);

OAI21xp5_ASAP7_75t_L g319 ( 
.A1(n_144),
.A2(n_320),
.B(n_321),
.Y(n_319)
);

NOR2xp33_ASAP7_75t_L g144 ( 
.A(n_145),
.B(n_146),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_L g321 ( 
.A(n_145),
.B(n_146),
.Y(n_321)
);

OAI21x1_ASAP7_75t_SL g149 ( 
.A1(n_150),
.A2(n_174),
.B(n_318),
.Y(n_149)
);

NOR2xp33_ASAP7_75t_L g150 ( 
.A(n_151),
.B(n_172),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_L g318 ( 
.A(n_151),
.B(n_172),
.Y(n_318)
);

MAJIxp5_ASAP7_75t_L g151 ( 
.A(n_152),
.B(n_155),
.C(n_156),
.Y(n_151)
);

XNOR2xp5_ASAP7_75t_L g201 ( 
.A(n_152),
.B(n_155),
.Y(n_201)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_154),
.Y(n_153)
);

XNOR2xp5_ASAP7_75t_L g200 ( 
.A(n_156),
.B(n_201),
.Y(n_200)
);

MAJIxp5_ASAP7_75t_L g156 ( 
.A(n_157),
.B(n_167),
.C(n_169),
.Y(n_156)
);

AOI22xp5_ASAP7_75t_L g178 ( 
.A1(n_157),
.A2(n_158),
.B1(n_179),
.B2(n_180),
.Y(n_178)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_158),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_L g158 ( 
.A(n_159),
.B(n_163),
.Y(n_158)
);

XNOR2xp5_ASAP7_75t_L g230 ( 
.A(n_159),
.B(n_163),
.Y(n_230)
);

CKINVDCx16_ASAP7_75t_R g161 ( 
.A(n_162),
.Y(n_161)
);

CKINVDCx16_ASAP7_75t_R g164 ( 
.A(n_165),
.Y(n_164)
);

XOR2xp5_ASAP7_75t_L g180 ( 
.A(n_167),
.B(n_169),
.Y(n_180)
);

INVxp67_ASAP7_75t_L g194 ( 
.A(n_168),
.Y(n_194)
);

INVxp67_ASAP7_75t_L g199 ( 
.A(n_170),
.Y(n_199)
);

AOI21xp5_ASAP7_75t_SL g174 ( 
.A1(n_175),
.A2(n_202),
.B(n_317),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_L g175 ( 
.A(n_176),
.B(n_200),
.Y(n_175)
);

NOR2xp33_ASAP7_75t_L g317 ( 
.A(n_176),
.B(n_200),
.Y(n_317)
);

MAJIxp5_ASAP7_75t_L g176 ( 
.A(n_177),
.B(n_181),
.C(n_182),
.Y(n_176)
);

AOI22xp5_ASAP7_75t_L g314 ( 
.A1(n_177),
.A2(n_178),
.B1(n_181),
.B2(n_315),
.Y(n_314)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_178),
.Y(n_177)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_180),
.Y(n_179)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_181),
.Y(n_315)
);

XNOR2xp5_ASAP7_75t_L g313 ( 
.A(n_182),
.B(n_314),
.Y(n_313)
);

MAJIxp5_ASAP7_75t_L g182 ( 
.A(n_183),
.B(n_191),
.C(n_195),
.Y(n_182)
);

XOR2xp5_ASAP7_75t_L g231 ( 
.A(n_183),
.B(n_232),
.Y(n_231)
);

NAND2xp5_ASAP7_75t_SL g183 ( 
.A(n_184),
.B(n_187),
.Y(n_183)
);

OAI22xp5_ASAP7_75t_SL g217 ( 
.A1(n_184),
.A2(n_185),
.B1(n_187),
.B2(n_218),
.Y(n_217)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_185),
.Y(n_184)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_187),
.Y(n_218)
);

INVxp67_ASAP7_75t_L g209 ( 
.A(n_189),
.Y(n_209)
);

XOR2xp5_ASAP7_75t_L g232 ( 
.A(n_191),
.B(n_195),
.Y(n_232)
);

INVxp67_ASAP7_75t_L g192 ( 
.A(n_193),
.Y(n_192)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_197),
.Y(n_196)
);

A2O1A1Ixp33_ASAP7_75t_SL g202 ( 
.A1(n_203),
.A2(n_233),
.B(n_311),
.C(n_316),
.Y(n_202)
);

OR2x2_ASAP7_75t_L g203 ( 
.A(n_204),
.B(n_227),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_L g310 ( 
.A(n_204),
.B(n_227),
.Y(n_310)
);

MAJIxp5_ASAP7_75t_L g204 ( 
.A(n_205),
.B(n_217),
.C(n_219),
.Y(n_204)
);

OAI22xp5_ASAP7_75t_SL g250 ( 
.A1(n_205),
.A2(n_206),
.B1(n_251),
.B2(n_252),
.Y(n_250)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_206),
.Y(n_205)
);

XOR2xp5_ASAP7_75t_L g206 ( 
.A(n_207),
.B(n_210),
.Y(n_206)
);

MAJIxp5_ASAP7_75t_L g229 ( 
.A(n_207),
.B(n_211),
.C(n_216),
.Y(n_229)
);

AOI22xp5_ASAP7_75t_L g210 ( 
.A1(n_211),
.A2(n_213),
.B1(n_215),
.B2(n_216),
.Y(n_210)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_211),
.Y(n_215)
);

INVxp67_ASAP7_75t_L g223 ( 
.A(n_212),
.Y(n_223)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_213),
.Y(n_216)
);

XNOR2xp5_ASAP7_75t_SL g251 ( 
.A(n_217),
.B(n_219),
.Y(n_251)
);

MAJIxp5_ASAP7_75t_L g219 ( 
.A(n_220),
.B(n_224),
.C(n_225),
.Y(n_219)
);

XNOR2xp5_ASAP7_75t_SL g237 ( 
.A(n_220),
.B(n_238),
.Y(n_237)
);

INVxp67_ASAP7_75t_L g221 ( 
.A(n_222),
.Y(n_221)
);

XNOR2xp5_ASAP7_75t_L g238 ( 
.A(n_224),
.B(n_225),
.Y(n_238)
);

XNOR2xp5_ASAP7_75t_L g227 ( 
.A(n_228),
.B(n_231),
.Y(n_227)
);

XNOR2xp5_ASAP7_75t_L g228 ( 
.A(n_229),
.B(n_230),
.Y(n_228)
);

MAJIxp5_ASAP7_75t_L g312 ( 
.A(n_229),
.B(n_230),
.C(n_231),
.Y(n_312)
);

NAND2xp5_ASAP7_75t_SL g233 ( 
.A(n_234),
.B(n_310),
.Y(n_233)
);

OAI21xp5_ASAP7_75t_L g234 ( 
.A1(n_235),
.A2(n_253),
.B(n_309),
.Y(n_234)
);

NOR2xp33_ASAP7_75t_L g235 ( 
.A(n_236),
.B(n_250),
.Y(n_235)
);

NAND2xp5_ASAP7_75t_SL g309 ( 
.A(n_236),
.B(n_250),
.Y(n_309)
);

MAJIxp5_ASAP7_75t_L g236 ( 
.A(n_237),
.B(n_239),
.C(n_242),
.Y(n_236)
);

XOR2xp5_ASAP7_75t_L g305 ( 
.A(n_237),
.B(n_306),
.Y(n_305)
);

OAI22xp5_ASAP7_75t_L g306 ( 
.A1(n_239),
.A2(n_242),
.B1(n_243),
.B2(n_307),
.Y(n_306)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_239),
.Y(n_307)
);

INVxp67_ASAP7_75t_L g240 ( 
.A(n_241),
.Y(n_240)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_243),
.Y(n_242)
);

NOR2xp33_ASAP7_75t_L g243 ( 
.A(n_244),
.B(n_248),
.Y(n_243)
);

OAI22xp5_ASAP7_75t_SL g300 ( 
.A1(n_244),
.A2(n_245),
.B1(n_248),
.B2(n_301),
.Y(n_300)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_245),
.Y(n_244)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_246),
.Y(n_297)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_248),
.Y(n_301)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_251),
.Y(n_252)
);

AOI21xp5_ASAP7_75t_L g253 ( 
.A1(n_254),
.A2(n_303),
.B(n_308),
.Y(n_253)
);

OAI21xp5_ASAP7_75t_SL g254 ( 
.A1(n_255),
.A2(n_291),
.B(n_302),
.Y(n_254)
);

AOI21xp5_ASAP7_75t_L g255 ( 
.A1(n_256),
.A2(n_271),
.B(n_290),
.Y(n_255)
);

NAND2xp5_ASAP7_75t_L g256 ( 
.A(n_257),
.B(n_264),
.Y(n_256)
);

NOR2xp33_ASAP7_75t_SL g290 ( 
.A(n_257),
.B(n_264),
.Y(n_290)
);

NAND2xp5_ASAP7_75t_SL g257 ( 
.A(n_258),
.B(n_262),
.Y(n_257)
);

OAI22xp5_ASAP7_75t_SL g277 ( 
.A1(n_258),
.A2(n_259),
.B1(n_262),
.B2(n_278),
.Y(n_277)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_259),
.Y(n_258)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_262),
.Y(n_278)
);

XNOR2xp5_ASAP7_75t_L g264 ( 
.A(n_265),
.B(n_269),
.Y(n_264)
);

XNOR2xp5_ASAP7_75t_L g265 ( 
.A(n_266),
.B(n_267),
.Y(n_265)
);

MAJIxp5_ASAP7_75t_L g292 ( 
.A(n_266),
.B(n_267),
.C(n_269),
.Y(n_292)
);

INVxp67_ASAP7_75t_L g299 ( 
.A(n_268),
.Y(n_299)
);

CKINVDCx14_ASAP7_75t_R g276 ( 
.A(n_270),
.Y(n_276)
);

OAI21xp5_ASAP7_75t_SL g271 ( 
.A1(n_272),
.A2(n_279),
.B(n_289),
.Y(n_271)
);

NOR2xp33_ASAP7_75t_L g272 ( 
.A(n_273),
.B(n_277),
.Y(n_272)
);

NAND2xp5_ASAP7_75t_SL g289 ( 
.A(n_273),
.B(n_277),
.Y(n_289)
);

INVxp67_ASAP7_75t_L g274 ( 
.A(n_275),
.Y(n_274)
);

AOI21xp5_ASAP7_75t_L g279 ( 
.A1(n_280),
.A2(n_285),
.B(n_288),
.Y(n_279)
);

NOR2xp33_ASAP7_75t_SL g280 ( 
.A(n_281),
.B(n_283),
.Y(n_280)
);

NAND2xp5_ASAP7_75t_L g285 ( 
.A(n_286),
.B(n_287),
.Y(n_285)
);

NOR2xp33_ASAP7_75t_SL g288 ( 
.A(n_286),
.B(n_287),
.Y(n_288)
);

NOR2xp33_ASAP7_75t_L g291 ( 
.A(n_292),
.B(n_293),
.Y(n_291)
);

NAND2xp5_ASAP7_75t_SL g302 ( 
.A(n_292),
.B(n_293),
.Y(n_302)
);

XNOR2xp5_ASAP7_75t_L g293 ( 
.A(n_294),
.B(n_300),
.Y(n_293)
);

XNOR2xp5_ASAP7_75t_L g294 ( 
.A(n_295),
.B(n_298),
.Y(n_294)
);

MAJIxp5_ASAP7_75t_L g304 ( 
.A(n_295),
.B(n_298),
.C(n_300),
.Y(n_304)
);

NAND2xp5_ASAP7_75t_L g303 ( 
.A(n_304),
.B(n_305),
.Y(n_303)
);

NOR2xp33_ASAP7_75t_SL g308 ( 
.A(n_304),
.B(n_305),
.Y(n_308)
);

NOR2xp33_ASAP7_75t_L g311 ( 
.A(n_312),
.B(n_313),
.Y(n_311)
);

NAND2xp5_ASAP7_75t_L g316 ( 
.A(n_312),
.B(n_313),
.Y(n_316)
);


endmodule