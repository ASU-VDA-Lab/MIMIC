module fake_jpeg_30360_n_519 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_519);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_519;

wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_252;
wire n_19;
wire n_182;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_17;
wire n_431;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_513;
wire n_283;
wire n_107;
wire n_490;
wire n_517;
wire n_415;
wire n_479;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_48;
wire n_465;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_256;
wire n_221;
wire n_454;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_508;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_474;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_511;
wire n_305;
wire n_161;
wire n_441;
wire n_342;
wire n_101;
wire n_226;
wire n_509;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_510;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_296;
wire n_384;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_491;
wire n_24;
wire n_467;
wire n_269;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_473;
wire n_45;
wire n_476;
wire n_337;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_481;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_333;
wire n_518;
wire n_378;
wire n_132;
wire n_133;
wire n_419;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_199;
wire n_260;
wire n_413;
wire n_275;
wire n_494;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_492;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_515;
wire n_347;
wire n_424;
wire n_55;
wire n_358;
wire n_312;
wire n_47;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_472;
wire n_279;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_484;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_469;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_482;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_512;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_516;
wire n_183;
wire n_409;
wire n_249;
wire n_412;
wire n_217;
wire n_471;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_402;
wire n_504;
wire n_438;
wire n_475;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_514;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

INVx1_ASAP7_75t_L g17 ( 
.A(n_8),
.Y(n_17)
);

BUFx5_ASAP7_75t_L g18 ( 
.A(n_16),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_16),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_8),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_4),
.Y(n_21)
);

BUFx5_ASAP7_75t_L g22 ( 
.A(n_14),
.Y(n_22)
);

BUFx10_ASAP7_75t_L g23 ( 
.A(n_11),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_9),
.Y(n_24)
);

BUFx12_ASAP7_75t_L g25 ( 
.A(n_10),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_1),
.Y(n_26)
);

INVx6_ASAP7_75t_L g27 ( 
.A(n_16),
.Y(n_27)
);

INVx3_ASAP7_75t_L g28 ( 
.A(n_5),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_10),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_9),
.Y(n_30)
);

INVxp67_ASAP7_75t_L g31 ( 
.A(n_7),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_8),
.Y(n_32)
);

CKINVDCx14_ASAP7_75t_R g33 ( 
.A(n_7),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_6),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_3),
.Y(n_35)
);

BUFx16f_ASAP7_75t_L g36 ( 
.A(n_6),
.Y(n_36)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_2),
.Y(n_37)
);

INVx2_ASAP7_75t_L g38 ( 
.A(n_10),
.Y(n_38)
);

BUFx6f_ASAP7_75t_SL g39 ( 
.A(n_14),
.Y(n_39)
);

INVx5_ASAP7_75t_L g40 ( 
.A(n_10),
.Y(n_40)
);

BUFx8_ASAP7_75t_L g41 ( 
.A(n_14),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_7),
.Y(n_42)
);

BUFx5_ASAP7_75t_L g43 ( 
.A(n_13),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_9),
.Y(n_44)
);

BUFx4f_ASAP7_75t_SL g45 ( 
.A(n_1),
.Y(n_45)
);

BUFx12f_ASAP7_75t_L g46 ( 
.A(n_7),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_2),
.Y(n_47)
);

BUFx12f_ASAP7_75t_L g48 ( 
.A(n_13),
.Y(n_48)
);

BUFx12f_ASAP7_75t_L g49 ( 
.A(n_13),
.Y(n_49)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_9),
.Y(n_50)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_4),
.Y(n_51)
);

BUFx16f_ASAP7_75t_L g52 ( 
.A(n_13),
.Y(n_52)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_23),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g130 ( 
.A(n_53),
.B(n_76),
.Y(n_130)
);

INVx11_ASAP7_75t_L g54 ( 
.A(n_36),
.Y(n_54)
);

INVx6_ASAP7_75t_L g122 ( 
.A(n_54),
.Y(n_122)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_38),
.Y(n_55)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_55),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_31),
.B(n_6),
.Y(n_56)
);

AND2x2_ASAP7_75t_L g107 ( 
.A(n_56),
.B(n_60),
.Y(n_107)
);

BUFx4f_ASAP7_75t_L g57 ( 
.A(n_39),
.Y(n_57)
);

BUFx2_ASAP7_75t_L g109 ( 
.A(n_57),
.Y(n_109)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_29),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g113 ( 
.A(n_58),
.Y(n_113)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_29),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g115 ( 
.A(n_59),
.Y(n_115)
);

AND2x2_ASAP7_75t_SL g60 ( 
.A(n_38),
.B(n_6),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_29),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g131 ( 
.A(n_61),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g62 ( 
.A(n_20),
.B(n_8),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_L g120 ( 
.A(n_62),
.B(n_69),
.Y(n_120)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_44),
.Y(n_63)
);

BUFx6f_ASAP7_75t_L g137 ( 
.A(n_63),
.Y(n_137)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_44),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g147 ( 
.A(n_64),
.Y(n_147)
);

INVx2_ASAP7_75t_L g65 ( 
.A(n_28),
.Y(n_65)
);

INVx2_ASAP7_75t_L g118 ( 
.A(n_65),
.Y(n_118)
);

INVx8_ASAP7_75t_L g66 ( 
.A(n_22),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g152 ( 
.A(n_66),
.Y(n_152)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_44),
.Y(n_67)
);

INVx6_ASAP7_75t_L g139 ( 
.A(n_67),
.Y(n_139)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_27),
.Y(n_68)
);

INVx6_ASAP7_75t_L g150 ( 
.A(n_68),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_L g69 ( 
.A(n_20),
.B(n_16),
.Y(n_69)
);

INVx3_ASAP7_75t_L g70 ( 
.A(n_46),
.Y(n_70)
);

INVx3_ASAP7_75t_L g106 ( 
.A(n_70),
.Y(n_106)
);

BUFx3_ASAP7_75t_L g71 ( 
.A(n_22),
.Y(n_71)
);

BUFx3_ASAP7_75t_L g144 ( 
.A(n_71),
.Y(n_144)
);

INVx3_ASAP7_75t_L g72 ( 
.A(n_22),
.Y(n_72)
);

INVx3_ASAP7_75t_L g108 ( 
.A(n_72),
.Y(n_108)
);

INVx3_ASAP7_75t_L g73 ( 
.A(n_46),
.Y(n_73)
);

INVx3_ASAP7_75t_L g110 ( 
.A(n_73),
.Y(n_110)
);

BUFx5_ASAP7_75t_L g74 ( 
.A(n_46),
.Y(n_74)
);

BUFx2_ASAP7_75t_L g158 ( 
.A(n_74),
.Y(n_158)
);

INVx2_ASAP7_75t_L g75 ( 
.A(n_28),
.Y(n_75)
);

INVx2_ASAP7_75t_L g123 ( 
.A(n_75),
.Y(n_123)
);

OR2x2_ASAP7_75t_L g76 ( 
.A(n_34),
.B(n_15),
.Y(n_76)
);

BUFx12f_ASAP7_75t_L g77 ( 
.A(n_36),
.Y(n_77)
);

INVx3_ASAP7_75t_L g111 ( 
.A(n_77),
.Y(n_111)
);

BUFx5_ASAP7_75t_L g78 ( 
.A(n_46),
.Y(n_78)
);

INVx4_ASAP7_75t_L g112 ( 
.A(n_78),
.Y(n_112)
);

BUFx6f_ASAP7_75t_L g79 ( 
.A(n_27),
.Y(n_79)
);

INVx6_ASAP7_75t_L g159 ( 
.A(n_79),
.Y(n_159)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_17),
.Y(n_80)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_80),
.Y(n_151)
);

INVx2_ASAP7_75t_L g81 ( 
.A(n_28),
.Y(n_81)
);

INVx2_ASAP7_75t_L g125 ( 
.A(n_81),
.Y(n_125)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_17),
.Y(n_82)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_82),
.Y(n_162)
);

BUFx6f_ASAP7_75t_L g83 ( 
.A(n_27),
.Y(n_83)
);

INVx3_ASAP7_75t_L g114 ( 
.A(n_83),
.Y(n_114)
);

INVx6_ASAP7_75t_L g84 ( 
.A(n_26),
.Y(n_84)
);

INVx2_ASAP7_75t_L g135 ( 
.A(n_84),
.Y(n_135)
);

BUFx6f_ASAP7_75t_L g85 ( 
.A(n_26),
.Y(n_85)
);

INVx3_ASAP7_75t_L g128 ( 
.A(n_85),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_SL g86 ( 
.A(n_34),
.B(n_15),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_L g146 ( 
.A(n_86),
.B(n_101),
.Y(n_146)
);

BUFx5_ASAP7_75t_L g87 ( 
.A(n_46),
.Y(n_87)
);

INVx4_ASAP7_75t_L g149 ( 
.A(n_87),
.Y(n_149)
);

INVx4_ASAP7_75t_L g88 ( 
.A(n_40),
.Y(n_88)
);

INVx3_ASAP7_75t_L g142 ( 
.A(n_88),
.Y(n_142)
);

BUFx6f_ASAP7_75t_L g89 ( 
.A(n_26),
.Y(n_89)
);

INVx4_ASAP7_75t_L g157 ( 
.A(n_89),
.Y(n_157)
);

BUFx6f_ASAP7_75t_L g90 ( 
.A(n_47),
.Y(n_90)
);

INVx2_ASAP7_75t_L g153 ( 
.A(n_90),
.Y(n_153)
);

INVx4_ASAP7_75t_L g91 ( 
.A(n_40),
.Y(n_91)
);

INVx3_ASAP7_75t_L g124 ( 
.A(n_91),
.Y(n_124)
);

BUFx6f_ASAP7_75t_L g92 ( 
.A(n_47),
.Y(n_92)
);

INVx2_ASAP7_75t_L g155 ( 
.A(n_92),
.Y(n_155)
);

BUFx6f_ASAP7_75t_L g93 ( 
.A(n_47),
.Y(n_93)
);

INVx2_ASAP7_75t_L g160 ( 
.A(n_93),
.Y(n_160)
);

INVx2_ASAP7_75t_L g94 ( 
.A(n_40),
.Y(n_94)
);

NAND2xp33_ASAP7_75t_SL g165 ( 
.A(n_94),
.B(n_97),
.Y(n_165)
);

BUFx6f_ASAP7_75t_L g95 ( 
.A(n_39),
.Y(n_95)
);

BUFx12f_ASAP7_75t_L g117 ( 
.A(n_95),
.Y(n_117)
);

INVx6_ASAP7_75t_L g96 ( 
.A(n_18),
.Y(n_96)
);

INVx3_ASAP7_75t_L g136 ( 
.A(n_96),
.Y(n_136)
);

INVx2_ASAP7_75t_L g97 ( 
.A(n_19),
.Y(n_97)
);

INVx2_ASAP7_75t_L g98 ( 
.A(n_19),
.Y(n_98)
);

INVx3_ASAP7_75t_L g166 ( 
.A(n_98),
.Y(n_166)
);

INVx2_ASAP7_75t_SL g99 ( 
.A(n_36),
.Y(n_99)
);

BUFx4f_ASAP7_75t_SL g129 ( 
.A(n_99),
.Y(n_129)
);

BUFx3_ASAP7_75t_L g100 ( 
.A(n_18),
.Y(n_100)
);

CKINVDCx20_ASAP7_75t_R g116 ( 
.A(n_100),
.Y(n_116)
);

BUFx6f_ASAP7_75t_L g101 ( 
.A(n_36),
.Y(n_101)
);

INVx8_ASAP7_75t_L g102 ( 
.A(n_43),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_L g133 ( 
.A(n_102),
.B(n_104),
.Y(n_133)
);

BUFx3_ASAP7_75t_L g103 ( 
.A(n_43),
.Y(n_103)
);

CKINVDCx20_ASAP7_75t_R g132 ( 
.A(n_103),
.Y(n_132)
);

BUFx5_ASAP7_75t_L g104 ( 
.A(n_48),
.Y(n_104)
);

BUFx6f_ASAP7_75t_L g105 ( 
.A(n_52),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_L g163 ( 
.A(n_105),
.B(n_41),
.Y(n_163)
);

AOI22xp33_ASAP7_75t_SL g119 ( 
.A1(n_100),
.A2(n_33),
.B1(n_48),
.B2(n_49),
.Y(n_119)
);

OAI22xp5_ASAP7_75t_L g179 ( 
.A1(n_119),
.A2(n_121),
.B1(n_126),
.B2(n_134),
.Y(n_179)
);

AOI22xp33_ASAP7_75t_SL g121 ( 
.A1(n_103),
.A2(n_33),
.B1(n_96),
.B2(n_102),
.Y(n_121)
);

AOI22xp33_ASAP7_75t_SL g126 ( 
.A1(n_57),
.A2(n_48),
.B1(n_49),
.B2(n_52),
.Y(n_126)
);

AOI22xp33_ASAP7_75t_L g134 ( 
.A1(n_84),
.A2(n_58),
.B1(n_63),
.B2(n_61),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_L g138 ( 
.A(n_76),
.B(n_42),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_SL g169 ( 
.A(n_138),
.B(n_141),
.Y(n_169)
);

AOI22xp5_ASAP7_75t_L g140 ( 
.A1(n_60),
.A2(n_59),
.B1(n_67),
.B2(n_64),
.Y(n_140)
);

OAI22xp5_ASAP7_75t_L g217 ( 
.A1(n_140),
.A2(n_143),
.B1(n_148),
.B2(n_156),
.Y(n_217)
);

NOR2xp33_ASAP7_75t_SL g141 ( 
.A(n_77),
.B(n_42),
.Y(n_141)
);

AOI22xp33_ASAP7_75t_L g143 ( 
.A1(n_85),
.A2(n_48),
.B1(n_49),
.B2(n_21),
.Y(n_143)
);

NOR2xp33_ASAP7_75t_L g145 ( 
.A(n_77),
.B(n_35),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_SL g182 ( 
.A(n_145),
.B(n_154),
.Y(n_182)
);

AOI22xp5_ASAP7_75t_L g148 ( 
.A1(n_68),
.A2(n_24),
.B1(n_30),
.B2(n_50),
.Y(n_148)
);

NOR2xp33_ASAP7_75t_L g154 ( 
.A(n_99),
.B(n_35),
.Y(n_154)
);

AOI22xp33_ASAP7_75t_SL g156 ( 
.A1(n_71),
.A2(n_49),
.B1(n_48),
.B2(n_52),
.Y(n_156)
);

AOI22xp5_ASAP7_75t_SL g161 ( 
.A1(n_88),
.A2(n_21),
.B1(n_32),
.B2(n_50),
.Y(n_161)
);

AND2x2_ASAP7_75t_L g212 ( 
.A(n_161),
.B(n_163),
.Y(n_212)
);

AOI22xp33_ASAP7_75t_SL g164 ( 
.A1(n_95),
.A2(n_49),
.B1(n_52),
.B2(n_24),
.Y(n_164)
);

AOI22xp33_ASAP7_75t_SL g178 ( 
.A1(n_164),
.A2(n_66),
.B1(n_158),
.B2(n_112),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_L g167 ( 
.A(n_120),
.B(n_107),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_L g236 ( 
.A(n_167),
.B(n_172),
.Y(n_236)
);

HB1xp67_ASAP7_75t_L g168 ( 
.A(n_124),
.Y(n_168)
);

INVx2_ASAP7_75t_L g221 ( 
.A(n_168),
.Y(n_221)
);

NOR2xp33_ASAP7_75t_L g170 ( 
.A(n_130),
.B(n_30),
.Y(n_170)
);

NOR2xp33_ASAP7_75t_L g224 ( 
.A(n_170),
.B(n_175),
.Y(n_224)
);

INVx2_ASAP7_75t_L g171 ( 
.A(n_106),
.Y(n_171)
);

INVx2_ASAP7_75t_L g229 ( 
.A(n_171),
.Y(n_229)
);

NAND2xp5_ASAP7_75t_L g172 ( 
.A(n_107),
.B(n_146),
.Y(n_172)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_151),
.Y(n_173)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_173),
.Y(n_220)
);

BUFx2_ASAP7_75t_SL g174 ( 
.A(n_129),
.Y(n_174)
);

INVxp67_ASAP7_75t_L g234 ( 
.A(n_174),
.Y(n_234)
);

CKINVDCx20_ASAP7_75t_R g175 ( 
.A(n_109),
.Y(n_175)
);

INVx5_ASAP7_75t_L g176 ( 
.A(n_122),
.Y(n_176)
);

INVx4_ASAP7_75t_L g225 ( 
.A(n_176),
.Y(n_225)
);

INVx2_ASAP7_75t_L g177 ( 
.A(n_110),
.Y(n_177)
);

INVx2_ASAP7_75t_L g235 ( 
.A(n_177),
.Y(n_235)
);

AOI22xp33_ASAP7_75t_SL g226 ( 
.A1(n_178),
.A2(n_191),
.B1(n_204),
.B2(n_206),
.Y(n_226)
);

INVx2_ASAP7_75t_L g180 ( 
.A(n_135),
.Y(n_180)
);

INVx2_ASAP7_75t_L g239 ( 
.A(n_180),
.Y(n_239)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_162),
.Y(n_181)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_181),
.Y(n_240)
);

NAND2xp5_ASAP7_75t_SL g183 ( 
.A(n_127),
.B(n_32),
.Y(n_183)
);

NOR2xp33_ASAP7_75t_L g245 ( 
.A(n_183),
.B(n_201),
.Y(n_245)
);

INVx11_ASAP7_75t_L g184 ( 
.A(n_152),
.Y(n_184)
);

INVx6_ASAP7_75t_L g251 ( 
.A(n_184),
.Y(n_251)
);

INVx3_ASAP7_75t_L g185 ( 
.A(n_122),
.Y(n_185)
);

INVx4_ASAP7_75t_L g228 ( 
.A(n_185),
.Y(n_228)
);

INVx3_ASAP7_75t_L g186 ( 
.A(n_117),
.Y(n_186)
);

INVx3_ASAP7_75t_L g222 ( 
.A(n_186),
.Y(n_222)
);

INVx2_ASAP7_75t_L g187 ( 
.A(n_153),
.Y(n_187)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_187),
.Y(n_223)
);

AOI22xp33_ASAP7_75t_L g188 ( 
.A1(n_139),
.A2(n_93),
.B1(n_92),
.B2(n_90),
.Y(n_188)
);

OAI22xp5_ASAP7_75t_SL g238 ( 
.A1(n_188),
.A2(n_196),
.B1(n_121),
.B2(n_119),
.Y(n_238)
);

INVx3_ASAP7_75t_L g189 ( 
.A(n_117),
.Y(n_189)
);

INVx3_ASAP7_75t_L g254 ( 
.A(n_189),
.Y(n_254)
);

NAND2xp5_ASAP7_75t_L g190 ( 
.A(n_166),
.B(n_37),
.Y(n_190)
);

NAND2xp5_ASAP7_75t_L g246 ( 
.A(n_190),
.B(n_203),
.Y(n_246)
);

AOI22xp33_ASAP7_75t_SL g191 ( 
.A1(n_166),
.A2(n_91),
.B1(n_70),
.B2(n_73),
.Y(n_191)
);

INVx4_ASAP7_75t_L g192 ( 
.A(n_124),
.Y(n_192)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_192),
.Y(n_243)
);

INVx2_ASAP7_75t_L g193 ( 
.A(n_155),
.Y(n_193)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_193),
.Y(n_249)
);

INVx2_ASAP7_75t_L g194 ( 
.A(n_160),
.Y(n_194)
);

BUFx3_ASAP7_75t_L g230 ( 
.A(n_194),
.Y(n_230)
);

BUFx2_ASAP7_75t_L g195 ( 
.A(n_136),
.Y(n_195)
);

CKINVDCx20_ASAP7_75t_R g231 ( 
.A(n_195),
.Y(n_231)
);

AOI22xp33_ASAP7_75t_L g196 ( 
.A1(n_139),
.A2(n_89),
.B1(n_83),
.B2(n_79),
.Y(n_196)
);

INVx2_ASAP7_75t_L g197 ( 
.A(n_118),
.Y(n_197)
);

BUFx3_ASAP7_75t_L g250 ( 
.A(n_197),
.Y(n_250)
);

OR2x2_ASAP7_75t_SL g198 ( 
.A(n_165),
.B(n_143),
.Y(n_198)
);

OR2x2_ASAP7_75t_L g242 ( 
.A(n_198),
.B(n_205),
.Y(n_242)
);

INVx2_ASAP7_75t_L g199 ( 
.A(n_123),
.Y(n_199)
);

BUFx6f_ASAP7_75t_L g241 ( 
.A(n_199),
.Y(n_241)
);

BUFx2_ASAP7_75t_L g200 ( 
.A(n_136),
.Y(n_200)
);

CKINVDCx16_ASAP7_75t_R g218 ( 
.A(n_200),
.Y(n_218)
);

CKINVDCx16_ASAP7_75t_R g201 ( 
.A(n_133),
.Y(n_201)
);

INVx2_ASAP7_75t_L g202 ( 
.A(n_125),
.Y(n_202)
);

CKINVDCx16_ASAP7_75t_R g227 ( 
.A(n_202),
.Y(n_227)
);

NAND2xp5_ASAP7_75t_L g203 ( 
.A(n_129),
.B(n_51),
.Y(n_203)
);

INVx6_ASAP7_75t_L g204 ( 
.A(n_113),
.Y(n_204)
);

NOR2xp33_ASAP7_75t_L g205 ( 
.A(n_116),
.B(n_54),
.Y(n_205)
);

INVx4_ASAP7_75t_L g206 ( 
.A(n_152),
.Y(n_206)
);

AOI22xp33_ASAP7_75t_SL g207 ( 
.A1(n_157),
.A2(n_51),
.B1(n_37),
.B2(n_105),
.Y(n_207)
);

AOI22xp33_ASAP7_75t_SL g232 ( 
.A1(n_207),
.A2(n_208),
.B1(n_209),
.B2(n_210),
.Y(n_232)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_108),
.Y(n_208)
);

INVx2_ASAP7_75t_L g209 ( 
.A(n_157),
.Y(n_209)
);

INVx2_ASAP7_75t_L g210 ( 
.A(n_128),
.Y(n_210)
);

NOR2xp33_ASAP7_75t_L g211 ( 
.A(n_132),
.B(n_25),
.Y(n_211)
);

NAND2xp5_ASAP7_75t_L g248 ( 
.A(n_211),
.B(n_213),
.Y(n_248)
);

INVx4_ASAP7_75t_L g213 ( 
.A(n_142),
.Y(n_213)
);

INVx5_ASAP7_75t_L g214 ( 
.A(n_111),
.Y(n_214)
);

OAI22xp33_ASAP7_75t_SL g256 ( 
.A1(n_214),
.A2(n_158),
.B1(n_149),
.B2(n_109),
.Y(n_256)
);

AND2x2_ASAP7_75t_L g215 ( 
.A(n_112),
.B(n_41),
.Y(n_215)
);

XNOR2xp5_ASAP7_75t_L g244 ( 
.A(n_215),
.B(n_216),
.Y(n_244)
);

NOR2xp33_ASAP7_75t_L g216 ( 
.A(n_129),
.B(n_25),
.Y(n_216)
);

AOI22xp5_ASAP7_75t_L g219 ( 
.A1(n_217),
.A2(n_159),
.B1(n_150),
.B2(n_114),
.Y(n_219)
);

AND2x2_ASAP7_75t_L g284 ( 
.A(n_219),
.B(n_237),
.Y(n_284)
);

MAJIxp5_ASAP7_75t_L g233 ( 
.A(n_212),
.B(n_144),
.C(n_149),
.Y(n_233)
);

XNOR2xp5_ASAP7_75t_L g283 ( 
.A(n_233),
.B(n_247),
.Y(n_283)
);

AOI22xp5_ASAP7_75t_L g237 ( 
.A1(n_212),
.A2(n_159),
.B1(n_150),
.B2(n_134),
.Y(n_237)
);

AOI22xp5_ASAP7_75t_L g265 ( 
.A1(n_238),
.A2(n_252),
.B1(n_253),
.B2(n_256),
.Y(n_265)
);

XNOR2xp5_ASAP7_75t_L g247 ( 
.A(n_212),
.B(n_156),
.Y(n_247)
);

AOI22xp5_ASAP7_75t_L g252 ( 
.A1(n_179),
.A2(n_115),
.B1(n_113),
.B2(n_131),
.Y(n_252)
);

AOI22xp5_ASAP7_75t_L g253 ( 
.A1(n_198),
.A2(n_115),
.B1(n_131),
.B2(n_137),
.Y(n_253)
);

MAJIxp5_ASAP7_75t_L g255 ( 
.A(n_190),
.B(n_203),
.C(n_182),
.Y(n_255)
);

XNOR2xp5_ASAP7_75t_SL g267 ( 
.A(n_255),
.B(n_215),
.Y(n_267)
);

NAND2xp5_ASAP7_75t_L g257 ( 
.A(n_246),
.B(n_199),
.Y(n_257)
);

NAND2xp5_ASAP7_75t_L g317 ( 
.A(n_257),
.B(n_270),
.Y(n_317)
);

CKINVDCx20_ASAP7_75t_R g258 ( 
.A(n_250),
.Y(n_258)
);

NOR2xp33_ASAP7_75t_L g300 ( 
.A(n_258),
.B(n_260),
.Y(n_300)
);

OAI21xp5_ASAP7_75t_L g259 ( 
.A1(n_242),
.A2(n_215),
.B(n_169),
.Y(n_259)
);

OAI21xp5_ASAP7_75t_L g295 ( 
.A1(n_259),
.A2(n_280),
.B(n_41),
.Y(n_295)
);

CKINVDCx20_ASAP7_75t_R g260 ( 
.A(n_250),
.Y(n_260)
);

NOR2xp33_ASAP7_75t_L g261 ( 
.A(n_245),
.B(n_213),
.Y(n_261)
);

NAND2xp5_ASAP7_75t_SL g307 ( 
.A(n_261),
.B(n_268),
.Y(n_307)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_223),
.Y(n_262)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_262),
.Y(n_291)
);

BUFx2_ASAP7_75t_L g263 ( 
.A(n_251),
.Y(n_263)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_263),
.Y(n_292)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_223),
.Y(n_264)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_264),
.Y(n_294)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_249),
.Y(n_266)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_266),
.Y(n_298)
);

XOR2xp5_ASAP7_75t_L g318 ( 
.A(n_267),
.B(n_221),
.Y(n_318)
);

CKINVDCx20_ASAP7_75t_R g268 ( 
.A(n_230),
.Y(n_268)
);

INVx3_ASAP7_75t_L g269 ( 
.A(n_228),
.Y(n_269)
);

BUFx3_ASAP7_75t_L g301 ( 
.A(n_269),
.Y(n_301)
);

NAND2xp5_ASAP7_75t_L g270 ( 
.A(n_246),
.B(n_197),
.Y(n_270)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_249),
.Y(n_271)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_271),
.Y(n_299)
);

BUFx6f_ASAP7_75t_L g272 ( 
.A(n_251),
.Y(n_272)
);

BUFx3_ASAP7_75t_L g305 ( 
.A(n_272),
.Y(n_305)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_239),
.Y(n_273)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_273),
.Y(n_306)
);

NOR2xp33_ASAP7_75t_L g274 ( 
.A(n_224),
.B(n_214),
.Y(n_274)
);

NAND2xp5_ASAP7_75t_SL g314 ( 
.A(n_274),
.B(n_275),
.Y(n_314)
);

NOR2xp33_ASAP7_75t_SL g275 ( 
.A(n_236),
.B(n_255),
.Y(n_275)
);

AOI22xp5_ASAP7_75t_L g276 ( 
.A1(n_247),
.A2(n_202),
.B1(n_137),
.B2(n_147),
.Y(n_276)
);

OAI22xp5_ASAP7_75t_SL g302 ( 
.A1(n_276),
.A2(n_226),
.B1(n_232),
.B2(n_231),
.Y(n_302)
);

INVxp33_ASAP7_75t_L g277 ( 
.A(n_218),
.Y(n_277)
);

CKINVDCx16_ASAP7_75t_R g296 ( 
.A(n_277),
.Y(n_296)
);

AOI21x1_ASAP7_75t_L g278 ( 
.A1(n_248),
.A2(n_126),
.B(n_164),
.Y(n_278)
);

OAI21xp5_ASAP7_75t_SL g313 ( 
.A1(n_278),
.A2(n_290),
.B(n_234),
.Y(n_313)
);

INVx4_ASAP7_75t_L g279 ( 
.A(n_222),
.Y(n_279)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_279),
.Y(n_309)
);

OAI21xp5_ASAP7_75t_L g280 ( 
.A1(n_242),
.A2(n_45),
.B(n_41),
.Y(n_280)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_239),
.Y(n_281)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_281),
.Y(n_311)
);

INVx2_ASAP7_75t_L g282 ( 
.A(n_241),
.Y(n_282)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_282),
.Y(n_312)
);

NAND2xp5_ASAP7_75t_L g285 ( 
.A(n_236),
.B(n_180),
.Y(n_285)
);

NAND2xp5_ASAP7_75t_SL g316 ( 
.A(n_285),
.B(n_287),
.Y(n_316)
);

MAJx2_ASAP7_75t_L g286 ( 
.A(n_233),
.B(n_171),
.C(n_177),
.Y(n_286)
);

MAJIxp5_ASAP7_75t_L g303 ( 
.A(n_286),
.B(n_244),
.C(n_243),
.Y(n_303)
);

NAND2xp5_ASAP7_75t_L g287 ( 
.A(n_248),
.B(n_193),
.Y(n_287)
);

OR2x6_ASAP7_75t_L g288 ( 
.A(n_253),
.B(n_206),
.Y(n_288)
);

AND2x2_ASAP7_75t_L g297 ( 
.A(n_288),
.B(n_238),
.Y(n_297)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_243),
.Y(n_289)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_289),
.Y(n_320)
);

OAI21xp33_ASAP7_75t_L g290 ( 
.A1(n_244),
.A2(n_192),
.B(n_195),
.Y(n_290)
);

OAI22xp5_ASAP7_75t_L g293 ( 
.A1(n_265),
.A2(n_219),
.B1(n_252),
.B2(n_237),
.Y(n_293)
);

AOI22xp5_ASAP7_75t_L g324 ( 
.A1(n_293),
.A2(n_302),
.B1(n_322),
.B2(n_288),
.Y(n_324)
);

OAI21xp5_ASAP7_75t_L g345 ( 
.A1(n_295),
.A2(n_315),
.B(n_296),
.Y(n_345)
);

OAI21xp5_ASAP7_75t_SL g323 ( 
.A1(n_297),
.A2(n_319),
.B(n_278),
.Y(n_323)
);

XNOR2xp5_ASAP7_75t_L g331 ( 
.A(n_303),
.B(n_313),
.Y(n_331)
);

AOI22xp5_ASAP7_75t_L g304 ( 
.A1(n_284),
.A2(n_220),
.B1(n_240),
.B2(n_147),
.Y(n_304)
);

OAI22xp5_ASAP7_75t_SL g335 ( 
.A1(n_304),
.A2(n_308),
.B1(n_310),
.B2(n_273),
.Y(n_335)
);

AOI22xp5_ASAP7_75t_L g308 ( 
.A1(n_284),
.A2(n_204),
.B1(n_227),
.B2(n_228),
.Y(n_308)
);

AOI22xp5_ASAP7_75t_L g310 ( 
.A1(n_284),
.A2(n_210),
.B1(n_187),
.B2(n_194),
.Y(n_310)
);

OAI21xp5_ASAP7_75t_L g315 ( 
.A1(n_280),
.A2(n_234),
.B(n_221),
.Y(n_315)
);

MAJIxp5_ASAP7_75t_L g332 ( 
.A(n_318),
.B(n_321),
.C(n_267),
.Y(n_332)
);

XOR2x2_ASAP7_75t_L g319 ( 
.A(n_283),
.B(n_235),
.Y(n_319)
);

MAJIxp5_ASAP7_75t_L g321 ( 
.A(n_283),
.B(n_229),
.C(n_235),
.Y(n_321)
);

OAI22xp5_ASAP7_75t_SL g322 ( 
.A1(n_265),
.A2(n_184),
.B1(n_200),
.B2(n_209),
.Y(n_322)
);

AOI21xp5_ASAP7_75t_L g359 ( 
.A1(n_323),
.A2(n_327),
.B(n_343),
.Y(n_359)
);

OAI22xp5_ASAP7_75t_L g372 ( 
.A1(n_324),
.A2(n_342),
.B1(n_347),
.B2(n_310),
.Y(n_372)
);

OAI32xp33_ASAP7_75t_L g325 ( 
.A1(n_317),
.A2(n_288),
.A3(n_257),
.B1(n_270),
.B2(n_285),
.Y(n_325)
);

INVx1_ASAP7_75t_L g361 ( 
.A(n_325),
.Y(n_361)
);

NOR2xp33_ASAP7_75t_L g326 ( 
.A(n_300),
.B(n_287),
.Y(n_326)
);

CKINVDCx20_ASAP7_75t_R g354 ( 
.A(n_326),
.Y(n_354)
);

OAI21xp5_ASAP7_75t_SL g327 ( 
.A1(n_297),
.A2(n_288),
.B(n_286),
.Y(n_327)
);

OAI22xp5_ASAP7_75t_L g328 ( 
.A1(n_297),
.A2(n_288),
.B1(n_276),
.B2(n_259),
.Y(n_328)
);

AOI22xp5_ASAP7_75t_L g357 ( 
.A1(n_328),
.A2(n_335),
.B1(n_336),
.B2(n_351),
.Y(n_357)
);

CKINVDCx20_ASAP7_75t_R g329 ( 
.A(n_307),
.Y(n_329)
);

CKINVDCx20_ASAP7_75t_R g381 ( 
.A(n_329),
.Y(n_381)
);

NOR2xp33_ASAP7_75t_L g330 ( 
.A(n_296),
.B(n_277),
.Y(n_330)
);

CKINVDCx20_ASAP7_75t_R g355 ( 
.A(n_330),
.Y(n_355)
);

MAJIxp5_ASAP7_75t_L g363 ( 
.A(n_332),
.B(n_340),
.C(n_294),
.Y(n_363)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_320),
.Y(n_333)
);

INVx1_ASAP7_75t_L g364 ( 
.A(n_333),
.Y(n_364)
);

AOI21xp5_ASAP7_75t_SL g334 ( 
.A1(n_295),
.A2(n_289),
.B(n_266),
.Y(n_334)
);

OAI21xp5_ASAP7_75t_L g379 ( 
.A1(n_334),
.A2(n_345),
.B(n_346),
.Y(n_379)
);

OAI22xp5_ASAP7_75t_SL g336 ( 
.A1(n_293),
.A2(n_316),
.B1(n_317),
.B2(n_314),
.Y(n_336)
);

XNOR2x2_ASAP7_75t_SL g337 ( 
.A(n_319),
.B(n_264),
.Y(n_337)
);

NAND2xp5_ASAP7_75t_L g366 ( 
.A(n_337),
.B(n_350),
.Y(n_366)
);

NAND2xp5_ASAP7_75t_L g338 ( 
.A(n_316),
.B(n_262),
.Y(n_338)
);

INVx1_ASAP7_75t_L g368 ( 
.A(n_338),
.Y(n_368)
);

CKINVDCx20_ASAP7_75t_R g339 ( 
.A(n_307),
.Y(n_339)
);

CKINVDCx20_ASAP7_75t_R g378 ( 
.A(n_339),
.Y(n_378)
);

MAJIxp5_ASAP7_75t_L g340 ( 
.A(n_319),
.B(n_271),
.C(n_281),
.Y(n_340)
);

CKINVDCx20_ASAP7_75t_R g341 ( 
.A(n_301),
.Y(n_341)
);

NOR2xp33_ASAP7_75t_L g362 ( 
.A(n_341),
.B(n_349),
.Y(n_362)
);

AOI22xp5_ASAP7_75t_L g342 ( 
.A1(n_302),
.A2(n_260),
.B1(n_263),
.B2(n_279),
.Y(n_342)
);

AOI22xp5_ASAP7_75t_SL g343 ( 
.A1(n_322),
.A2(n_269),
.B1(n_282),
.B2(n_225),
.Y(n_343)
);

INVx1_ASAP7_75t_L g344 ( 
.A(n_320),
.Y(n_344)
);

INVx1_ASAP7_75t_L g380 ( 
.A(n_344),
.Y(n_380)
);

AOI22xp5_ASAP7_75t_SL g346 ( 
.A1(n_313),
.A2(n_315),
.B1(n_291),
.B2(n_299),
.Y(n_346)
);

AOI22xp5_ASAP7_75t_L g347 ( 
.A1(n_314),
.A2(n_272),
.B1(n_225),
.B2(n_241),
.Y(n_347)
);

INVx1_ASAP7_75t_L g348 ( 
.A(n_291),
.Y(n_348)
);

INVx1_ASAP7_75t_SL g370 ( 
.A(n_348),
.Y(n_370)
);

CKINVDCx20_ASAP7_75t_R g349 ( 
.A(n_301),
.Y(n_349)
);

NAND2xp5_ASAP7_75t_L g350 ( 
.A(n_321),
.B(n_229),
.Y(n_350)
);

OAI22xp5_ASAP7_75t_SL g351 ( 
.A1(n_304),
.A2(n_185),
.B1(n_230),
.B2(n_176),
.Y(n_351)
);

INVx1_ASAP7_75t_L g352 ( 
.A(n_294),
.Y(n_352)
);

INVx2_ASAP7_75t_L g382 ( 
.A(n_352),
.Y(n_382)
);

NOR2x1p5_ASAP7_75t_SL g353 ( 
.A(n_318),
.B(n_45),
.Y(n_353)
);

AOI22xp5_ASAP7_75t_L g365 ( 
.A1(n_353),
.A2(n_298),
.B1(n_309),
.B2(n_311),
.Y(n_365)
);

XOR2x2_ASAP7_75t_L g356 ( 
.A(n_353),
.B(n_303),
.Y(n_356)
);

XNOR2xp5_ASAP7_75t_L g392 ( 
.A(n_356),
.B(n_358),
.Y(n_392)
);

XOR2x2_ASAP7_75t_L g358 ( 
.A(n_353),
.B(n_308),
.Y(n_358)
);

NAND3xp33_ASAP7_75t_L g360 ( 
.A(n_329),
.B(n_299),
.C(n_298),
.Y(n_360)
);

NOR2xp33_ASAP7_75t_L g390 ( 
.A(n_360),
.B(n_371),
.Y(n_390)
);

MAJIxp5_ASAP7_75t_L g385 ( 
.A(n_363),
.B(n_367),
.C(n_373),
.Y(n_385)
);

OAI22xp5_ASAP7_75t_SL g389 ( 
.A1(n_365),
.A2(n_369),
.B1(n_370),
.B2(n_357),
.Y(n_389)
);

MAJIxp5_ASAP7_75t_L g367 ( 
.A(n_332),
.B(n_311),
.C(n_306),
.Y(n_367)
);

AOI22xp5_ASAP7_75t_L g369 ( 
.A1(n_328),
.A2(n_292),
.B1(n_306),
.B2(n_309),
.Y(n_369)
);

HB1xp67_ASAP7_75t_L g371 ( 
.A(n_333),
.Y(n_371)
);

AOI22xp5_ASAP7_75t_L g397 ( 
.A1(n_372),
.A2(n_335),
.B1(n_351),
.B2(n_342),
.Y(n_397)
);

MAJIxp5_ASAP7_75t_L g373 ( 
.A(n_331),
.B(n_292),
.C(n_312),
.Y(n_373)
);

MAJIxp5_ASAP7_75t_L g374 ( 
.A(n_331),
.B(n_312),
.C(n_254),
.Y(n_374)
);

MAJIxp5_ASAP7_75t_L g387 ( 
.A(n_374),
.B(n_377),
.C(n_327),
.Y(n_387)
);

XOR2xp5_ASAP7_75t_L g375 ( 
.A(n_340),
.B(n_254),
.Y(n_375)
);

XOR2xp5_ASAP7_75t_L g388 ( 
.A(n_375),
.B(n_383),
.Y(n_388)
);

NOR2xp33_ASAP7_75t_L g376 ( 
.A(n_339),
.B(n_336),
.Y(n_376)
);

CKINVDCx14_ASAP7_75t_R g410 ( 
.A(n_376),
.Y(n_410)
);

MAJIxp5_ASAP7_75t_L g377 ( 
.A(n_350),
.B(n_222),
.C(n_305),
.Y(n_377)
);

XNOR2xp5_ASAP7_75t_L g383 ( 
.A(n_323),
.B(n_144),
.Y(n_383)
);

NAND2xp5_ASAP7_75t_SL g384 ( 
.A(n_326),
.B(n_189),
.Y(n_384)
);

CKINVDCx16_ASAP7_75t_R g396 ( 
.A(n_384),
.Y(n_396)
);

OAI21xp5_ASAP7_75t_SL g386 ( 
.A1(n_359),
.A2(n_334),
.B(n_346),
.Y(n_386)
);

NOR2xp33_ASAP7_75t_L g423 ( 
.A(n_386),
.B(n_359),
.Y(n_423)
);

XNOR2x1_ASAP7_75t_L g413 ( 
.A(n_387),
.B(n_374),
.Y(n_413)
);

AOI22xp5_ASAP7_75t_SL g428 ( 
.A1(n_389),
.A2(n_394),
.B1(n_403),
.B2(n_404),
.Y(n_428)
);

INVx1_ASAP7_75t_L g391 ( 
.A(n_364),
.Y(n_391)
);

INVx1_ASAP7_75t_L g414 ( 
.A(n_391),
.Y(n_414)
);

XOR2xp5_ASAP7_75t_L g393 ( 
.A(n_375),
.B(n_345),
.Y(n_393)
);

XOR2xp5_ASAP7_75t_L g417 ( 
.A(n_393),
.B(n_405),
.Y(n_417)
);

OAI22xp5_ASAP7_75t_SL g394 ( 
.A1(n_357),
.A2(n_361),
.B1(n_324),
.B2(n_369),
.Y(n_394)
);

NAND2xp5_ASAP7_75t_L g395 ( 
.A(n_381),
.B(n_338),
.Y(n_395)
);

INVx1_ASAP7_75t_L g418 ( 
.A(n_395),
.Y(n_418)
);

OAI22xp5_ASAP7_75t_SL g432 ( 
.A1(n_397),
.A2(n_399),
.B1(n_408),
.B2(n_365),
.Y(n_432)
);

NAND2xp5_ASAP7_75t_L g398 ( 
.A(n_381),
.B(n_344),
.Y(n_398)
);

INVx1_ASAP7_75t_L g421 ( 
.A(n_398),
.Y(n_421)
);

AOI22xp5_ASAP7_75t_L g399 ( 
.A1(n_361),
.A2(n_325),
.B1(n_337),
.B2(n_348),
.Y(n_399)
);

MAJIxp5_ASAP7_75t_L g400 ( 
.A(n_363),
.B(n_337),
.C(n_347),
.Y(n_400)
);

MAJIxp5_ASAP7_75t_L g426 ( 
.A(n_400),
.B(n_356),
.C(n_358),
.Y(n_426)
);

INVx1_ASAP7_75t_L g401 ( 
.A(n_364),
.Y(n_401)
);

INVx1_ASAP7_75t_L g434 ( 
.A(n_401),
.Y(n_434)
);

INVx1_ASAP7_75t_L g402 ( 
.A(n_380),
.Y(n_402)
);

INVx1_ASAP7_75t_L g435 ( 
.A(n_402),
.Y(n_435)
);

OAI22xp5_ASAP7_75t_SL g403 ( 
.A1(n_368),
.A2(n_343),
.B1(n_352),
.B2(n_330),
.Y(n_403)
);

OAI22xp5_ASAP7_75t_L g404 ( 
.A1(n_378),
.A2(n_349),
.B1(n_341),
.B2(n_305),
.Y(n_404)
);

XOR2xp5_ASAP7_75t_L g405 ( 
.A(n_373),
.B(n_101),
.Y(n_405)
);

NAND2xp5_ASAP7_75t_SL g406 ( 
.A(n_354),
.B(n_186),
.Y(n_406)
);

NAND2xp5_ASAP7_75t_L g415 ( 
.A(n_406),
.B(n_407),
.Y(n_415)
);

NAND2xp5_ASAP7_75t_SL g407 ( 
.A(n_354),
.B(n_12),
.Y(n_407)
);

AOI22xp5_ASAP7_75t_SL g408 ( 
.A1(n_355),
.A2(n_23),
.B1(n_117),
.B2(n_45),
.Y(n_408)
);

INVx1_ASAP7_75t_L g409 ( 
.A(n_380),
.Y(n_409)
);

CKINVDCx16_ASAP7_75t_R g420 ( 
.A(n_409),
.Y(n_420)
);

CKINVDCx20_ASAP7_75t_R g411 ( 
.A(n_362),
.Y(n_411)
);

NAND2xp5_ASAP7_75t_L g416 ( 
.A(n_411),
.B(n_412),
.Y(n_416)
);

NAND2xp5_ASAP7_75t_L g412 ( 
.A(n_368),
.B(n_0),
.Y(n_412)
);

XOR2xp5_ASAP7_75t_L g440 ( 
.A(n_413),
.B(n_425),
.Y(n_440)
);

XNOR2xp5_ASAP7_75t_L g419 ( 
.A(n_405),
.B(n_385),
.Y(n_419)
);

XNOR2xp5_ASAP7_75t_L g442 ( 
.A(n_419),
.B(n_422),
.Y(n_442)
);

XNOR2xp5_ASAP7_75t_L g422 ( 
.A(n_385),
.B(n_387),
.Y(n_422)
);

AOI21xp5_ASAP7_75t_L g446 ( 
.A1(n_423),
.A2(n_401),
.B(n_408),
.Y(n_446)
);

OAI21xp5_ASAP7_75t_L g424 ( 
.A1(n_399),
.A2(n_379),
.B(n_366),
.Y(n_424)
);

OAI21xp5_ASAP7_75t_L g449 ( 
.A1(n_424),
.A2(n_382),
.B(n_45),
.Y(n_449)
);

XOR2xp5_ASAP7_75t_L g425 ( 
.A(n_388),
.B(n_367),
.Y(n_425)
);

XOR2xp5_ASAP7_75t_L g445 ( 
.A(n_426),
.B(n_430),
.Y(n_445)
);

XNOR2xp5_ASAP7_75t_L g427 ( 
.A(n_388),
.B(n_379),
.Y(n_427)
);

NOR2xp33_ASAP7_75t_L g436 ( 
.A(n_427),
.B(n_410),
.Y(n_436)
);

MAJIxp5_ASAP7_75t_L g429 ( 
.A(n_400),
.B(n_377),
.C(n_366),
.Y(n_429)
);

MAJIxp5_ASAP7_75t_L g441 ( 
.A(n_429),
.B(n_398),
.C(n_395),
.Y(n_441)
);

XOR2xp5_ASAP7_75t_L g430 ( 
.A(n_392),
.B(n_383),
.Y(n_430)
);

XOR2xp5_ASAP7_75t_L g431 ( 
.A(n_392),
.B(n_393),
.Y(n_431)
);

XOR2xp5_ASAP7_75t_L g447 ( 
.A(n_431),
.B(n_433),
.Y(n_447)
);

AOI22xp5_ASAP7_75t_SL g439 ( 
.A1(n_432),
.A2(n_394),
.B1(n_403),
.B2(n_389),
.Y(n_439)
);

XNOR2xp5_ASAP7_75t_SL g433 ( 
.A(n_386),
.B(n_370),
.Y(n_433)
);

XNOR2xp5_ASAP7_75t_L g463 ( 
.A(n_436),
.B(n_448),
.Y(n_463)
);

OAI22xp5_ASAP7_75t_L g437 ( 
.A1(n_428),
.A2(n_390),
.B1(n_397),
.B2(n_396),
.Y(n_437)
);

INVx1_ASAP7_75t_L g459 ( 
.A(n_437),
.Y(n_459)
);

NAND2xp5_ASAP7_75t_L g438 ( 
.A(n_415),
.B(n_411),
.Y(n_438)
);

NAND2xp5_ASAP7_75t_L g456 ( 
.A(n_438),
.B(n_443),
.Y(n_456)
);

OAI22xp5_ASAP7_75t_SL g471 ( 
.A1(n_439),
.A2(n_454),
.B1(n_12),
.B2(n_1),
.Y(n_471)
);

NAND2xp5_ASAP7_75t_SL g457 ( 
.A(n_441),
.B(n_446),
.Y(n_457)
);

OAI22xp5_ASAP7_75t_L g443 ( 
.A1(n_428),
.A2(n_409),
.B1(n_391),
.B2(n_402),
.Y(n_443)
);

NOR2xp33_ASAP7_75t_L g444 ( 
.A(n_416),
.B(n_404),
.Y(n_444)
);

NAND2xp5_ASAP7_75t_L g460 ( 
.A(n_444),
.B(n_450),
.Y(n_460)
);

XOR2xp5_ASAP7_75t_L g448 ( 
.A(n_417),
.B(n_412),
.Y(n_448)
);

XNOR2xp5_ASAP7_75t_L g464 ( 
.A(n_449),
.B(n_433),
.Y(n_464)
);

BUFx24_ASAP7_75t_SL g450 ( 
.A(n_422),
.Y(n_450)
);

OAI21xp5_ASAP7_75t_SL g451 ( 
.A1(n_426),
.A2(n_382),
.B(n_11),
.Y(n_451)
);

NAND2xp5_ASAP7_75t_SL g458 ( 
.A(n_451),
.B(n_420),
.Y(n_458)
);

OAI22xp5_ASAP7_75t_SL g452 ( 
.A1(n_424),
.A2(n_11),
.B1(n_15),
.B2(n_14),
.Y(n_452)
);

NAND2xp5_ASAP7_75t_L g467 ( 
.A(n_452),
.B(n_453),
.Y(n_467)
);

OAI22xp5_ASAP7_75t_SL g453 ( 
.A1(n_418),
.A2(n_15),
.B1(n_12),
.B2(n_11),
.Y(n_453)
);

AOI22xp5_ASAP7_75t_L g454 ( 
.A1(n_432),
.A2(n_12),
.B1(n_1),
.B2(n_2),
.Y(n_454)
);

NOR2xp33_ASAP7_75t_L g455 ( 
.A(n_441),
.B(n_429),
.Y(n_455)
);

NAND2xp5_ASAP7_75t_L g472 ( 
.A(n_455),
.B(n_458),
.Y(n_472)
);

NAND2xp5_ASAP7_75t_SL g461 ( 
.A(n_442),
.B(n_419),
.Y(n_461)
);

NAND2xp5_ASAP7_75t_L g473 ( 
.A(n_461),
.B(n_464),
.Y(n_473)
);

MAJIxp5_ASAP7_75t_L g462 ( 
.A(n_442),
.B(n_413),
.C(n_425),
.Y(n_462)
);

MAJIxp5_ASAP7_75t_L g474 ( 
.A(n_462),
.B(n_466),
.C(n_470),
.Y(n_474)
);

OAI21xp5_ASAP7_75t_L g465 ( 
.A1(n_439),
.A2(n_421),
.B(n_434),
.Y(n_465)
);

XNOR2xp5_ASAP7_75t_SL g484 ( 
.A(n_465),
.B(n_0),
.Y(n_484)
);

MAJIxp5_ASAP7_75t_L g466 ( 
.A(n_440),
.B(n_417),
.C(n_431),
.Y(n_466)
);

AND2x2_ASAP7_75t_L g468 ( 
.A(n_449),
.B(n_427),
.Y(n_468)
);

AND2x2_ASAP7_75t_L g476 ( 
.A(n_468),
.B(n_447),
.Y(n_476)
);

NAND2xp5_ASAP7_75t_SL g469 ( 
.A(n_445),
.B(n_435),
.Y(n_469)
);

NAND2xp5_ASAP7_75t_L g481 ( 
.A(n_469),
.B(n_463),
.Y(n_481)
);

MAJIxp5_ASAP7_75t_L g470 ( 
.A(n_440),
.B(n_430),
.C(n_414),
.Y(n_470)
);

XOR2xp5_ASAP7_75t_L g475 ( 
.A(n_471),
.B(n_452),
.Y(n_475)
);

AOI22xp5_ASAP7_75t_L g487 ( 
.A1(n_475),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_487)
);

NAND2xp5_ASAP7_75t_L g494 ( 
.A(n_476),
.B(n_482),
.Y(n_494)
);

MAJIxp5_ASAP7_75t_L g477 ( 
.A(n_462),
.B(n_445),
.C(n_448),
.Y(n_477)
);

NAND2xp5_ASAP7_75t_SL g492 ( 
.A(n_477),
.B(n_478),
.Y(n_492)
);

XNOR2xp5_ASAP7_75t_L g478 ( 
.A(n_470),
.B(n_463),
.Y(n_478)
);

AOI21xp33_ASAP7_75t_L g479 ( 
.A1(n_457),
.A2(n_446),
.B(n_447),
.Y(n_479)
);

INVx1_ASAP7_75t_L g489 ( 
.A(n_479),
.Y(n_489)
);

OAI21xp5_ASAP7_75t_SL g480 ( 
.A1(n_460),
.A2(n_453),
.B(n_454),
.Y(n_480)
);

INVx1_ASAP7_75t_L g498 ( 
.A(n_480),
.Y(n_498)
);

NOR2xp33_ASAP7_75t_L g488 ( 
.A(n_481),
.B(n_484),
.Y(n_488)
);

OAI21xp5_ASAP7_75t_L g482 ( 
.A1(n_456),
.A2(n_459),
.B(n_468),
.Y(n_482)
);

OAI211xp5_ASAP7_75t_L g483 ( 
.A1(n_467),
.A2(n_465),
.B(n_464),
.C(n_471),
.Y(n_483)
);

NOR2xp33_ASAP7_75t_SL g495 ( 
.A(n_483),
.B(n_3),
.Y(n_495)
);

NAND2xp5_ASAP7_75t_L g485 ( 
.A(n_466),
.B(n_23),
.Y(n_485)
);

NOR2xp33_ASAP7_75t_L g496 ( 
.A(n_485),
.B(n_486),
.Y(n_496)
);

NOR2xp33_ASAP7_75t_L g486 ( 
.A(n_455),
.B(n_25),
.Y(n_486)
);

NOR2xp33_ASAP7_75t_L g501 ( 
.A(n_487),
.B(n_484),
.Y(n_501)
);

OAI21xp5_ASAP7_75t_SL g490 ( 
.A1(n_472),
.A2(n_0),
.B(n_2),
.Y(n_490)
);

AOI21xp5_ASAP7_75t_L g500 ( 
.A1(n_490),
.A2(n_3),
.B(n_4),
.Y(n_500)
);

AOI22xp5_ASAP7_75t_L g491 ( 
.A1(n_475),
.A2(n_0),
.B1(n_3),
.B2(n_4),
.Y(n_491)
);

NAND2xp5_ASAP7_75t_L g504 ( 
.A(n_491),
.B(n_493),
.Y(n_504)
);

OAI22xp5_ASAP7_75t_SL g493 ( 
.A1(n_473),
.A2(n_23),
.B1(n_4),
.B2(n_5),
.Y(n_493)
);

NAND2xp5_ASAP7_75t_L g505 ( 
.A(n_495),
.B(n_497),
.Y(n_505)
);

NOR2xp33_ASAP7_75t_L g497 ( 
.A(n_474),
.B(n_477),
.Y(n_497)
);

OAI21xp5_ASAP7_75t_SL g499 ( 
.A1(n_489),
.A2(n_474),
.B(n_476),
.Y(n_499)
);

NAND2xp5_ASAP7_75t_SL g508 ( 
.A(n_499),
.B(n_500),
.Y(n_508)
);

INVxp67_ASAP7_75t_L g507 ( 
.A(n_501),
.Y(n_507)
);

NOR2xp33_ASAP7_75t_L g502 ( 
.A(n_492),
.B(n_25),
.Y(n_502)
);

NOR2xp33_ASAP7_75t_SL g510 ( 
.A(n_502),
.B(n_496),
.Y(n_510)
);

NOR2xp33_ASAP7_75t_L g503 ( 
.A(n_494),
.B(n_3),
.Y(n_503)
);

OAI21xp5_ASAP7_75t_L g509 ( 
.A1(n_503),
.A2(n_506),
.B(n_488),
.Y(n_509)
);

AOI21xp5_ASAP7_75t_SL g506 ( 
.A1(n_494),
.A2(n_23),
.B(n_5),
.Y(n_506)
);

INVx1_ASAP7_75t_L g512 ( 
.A(n_509),
.Y(n_512)
);

INVx1_ASAP7_75t_L g513 ( 
.A(n_510),
.Y(n_513)
);

A2O1A1O1Ixp25_ASAP7_75t_SL g511 ( 
.A1(n_503),
.A2(n_498),
.B(n_487),
.C(n_491),
.D(n_490),
.Y(n_511)
);

MAJx2_ASAP7_75t_L g514 ( 
.A(n_511),
.B(n_504),
.C(n_505),
.Y(n_514)
);

XOR2xp5_ASAP7_75t_L g516 ( 
.A(n_514),
.B(n_493),
.Y(n_516)
);

AOI21xp5_ASAP7_75t_L g515 ( 
.A1(n_512),
.A2(n_508),
.B(n_507),
.Y(n_515)
);

AOI21xp5_ASAP7_75t_SL g517 ( 
.A1(n_515),
.A2(n_516),
.B(n_513),
.Y(n_517)
);

INVx1_ASAP7_75t_L g518 ( 
.A(n_517),
.Y(n_518)
);

XOR2xp5_ASAP7_75t_L g519 ( 
.A(n_518),
.B(n_5),
.Y(n_519)
);


endmodule