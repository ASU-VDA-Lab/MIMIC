module fake_jpeg_28635_n_168 (n_13, n_21, n_33, n_1, n_45, n_10, n_23, n_27, n_6, n_22, n_47, n_14, n_40, n_19, n_18, n_20, n_35, n_48, n_46, n_41, n_4, n_34, n_30, n_39, n_42, n_16, n_49, n_3, n_0, n_24, n_28, n_38, n_26, n_44, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_43, n_50, n_12, n_32, n_8, n_15, n_7, n_168);

input n_13;
input n_21;
input n_33;
input n_1;
input n_45;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_47;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_48;
input n_46;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_42;
input n_16;
input n_49;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_44;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_43;
input n_50;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_168;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_51;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_84;
wire n_59;
wire n_98;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_76;
wire n_127;
wire n_154;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_155;
wire n_103;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_57;
wire n_119;
wire n_69;
wire n_83;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_106;
wire n_111;
wire n_143;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_139;
wire n_78;
wire n_165;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_162;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_91;
wire n_54;
wire n_93;
wire n_161;
wire n_138;
wire n_101;
wire n_149;
wire n_157;
wire n_87;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_153;
wire n_135;
wire n_62;
wire n_167;
wire n_120;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_40),
.Y(n_51)
);

INVx2_ASAP7_75t_L g52 ( 
.A(n_45),
.Y(n_52)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_15),
.Y(n_53)
);

BUFx3_ASAP7_75t_L g54 ( 
.A(n_11),
.Y(n_54)
);

CKINVDCx20_ASAP7_75t_R g55 ( 
.A(n_19),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_SL g56 ( 
.A(n_46),
.B(n_38),
.Y(n_56)
);

BUFx3_ASAP7_75t_L g57 ( 
.A(n_18),
.Y(n_57)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_35),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_13),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_SL g60 ( 
.A(n_5),
.B(n_29),
.Y(n_60)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_8),
.Y(n_61)
);

CKINVDCx20_ASAP7_75t_R g62 ( 
.A(n_10),
.Y(n_62)
);

CKINVDCx20_ASAP7_75t_R g63 ( 
.A(n_28),
.Y(n_63)
);

CKINVDCx20_ASAP7_75t_R g64 ( 
.A(n_23),
.Y(n_64)
);

BUFx4f_ASAP7_75t_L g65 ( 
.A(n_2),
.Y(n_65)
);

INVx3_ASAP7_75t_L g66 ( 
.A(n_48),
.Y(n_66)
);

BUFx10_ASAP7_75t_L g67 ( 
.A(n_49),
.Y(n_67)
);

INVx5_ASAP7_75t_L g68 ( 
.A(n_2),
.Y(n_68)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_17),
.Y(n_69)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_39),
.Y(n_70)
);

BUFx16f_ASAP7_75t_L g71 ( 
.A(n_31),
.Y(n_71)
);

BUFx10_ASAP7_75t_L g72 ( 
.A(n_8),
.Y(n_72)
);

CKINVDCx20_ASAP7_75t_R g73 ( 
.A(n_25),
.Y(n_73)
);

CKINVDCx20_ASAP7_75t_R g74 ( 
.A(n_11),
.Y(n_74)
);

INVx11_ASAP7_75t_L g75 ( 
.A(n_71),
.Y(n_75)
);

INVx5_ASAP7_75t_L g84 ( 
.A(n_75),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g76 ( 
.A(n_56),
.B(n_61),
.Y(n_76)
);

XOR2xp5_ASAP7_75t_L g92 ( 
.A(n_76),
.B(n_56),
.Y(n_92)
);

BUFx5_ASAP7_75t_L g77 ( 
.A(n_71),
.Y(n_77)
);

INVx3_ASAP7_75t_SL g94 ( 
.A(n_77),
.Y(n_94)
);

BUFx12f_ASAP7_75t_L g78 ( 
.A(n_68),
.Y(n_78)
);

INVx3_ASAP7_75t_L g88 ( 
.A(n_78),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_62),
.B(n_0),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_79),
.B(n_81),
.Y(n_85)
);

BUFx6f_ASAP7_75t_L g80 ( 
.A(n_51),
.Y(n_80)
);

INVx11_ASAP7_75t_L g98 ( 
.A(n_80),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_74),
.B(n_0),
.Y(n_81)
);

INVx3_ASAP7_75t_L g82 ( 
.A(n_54),
.Y(n_82)
);

INVx3_ASAP7_75t_L g91 ( 
.A(n_82),
.Y(n_91)
);

CKINVDCx16_ASAP7_75t_R g83 ( 
.A(n_65),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_83),
.B(n_73),
.Y(n_86)
);

AND2x2_ASAP7_75t_L g105 ( 
.A(n_86),
.B(n_69),
.Y(n_105)
);

INVx5_ASAP7_75t_L g87 ( 
.A(n_77),
.Y(n_87)
);

BUFx3_ASAP7_75t_L g104 ( 
.A(n_87),
.Y(n_104)
);

AOI22xp5_ASAP7_75t_L g89 ( 
.A1(n_80),
.A2(n_65),
.B1(n_51),
.B2(n_59),
.Y(n_89)
);

OAI22xp5_ASAP7_75t_L g108 ( 
.A1(n_89),
.A2(n_59),
.B1(n_67),
.B2(n_72),
.Y(n_108)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_82),
.Y(n_90)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_90),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_L g112 ( 
.A(n_92),
.B(n_3),
.Y(n_112)
);

AOI21xp33_ASAP7_75t_L g93 ( 
.A1(n_76),
.A2(n_60),
.B(n_70),
.Y(n_93)
);

OAI32xp33_ASAP7_75t_L g106 ( 
.A1(n_93),
.A2(n_63),
.A3(n_67),
.B1(n_72),
.B2(n_54),
.Y(n_106)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_75),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_95),
.B(n_55),
.Y(n_101)
);

O2A1O1Ixp33_ASAP7_75t_L g96 ( 
.A1(n_78),
.A2(n_52),
.B(n_64),
.C(n_53),
.Y(n_96)
);

OA22x2_ASAP7_75t_L g116 ( 
.A1(n_96),
.A2(n_94),
.B1(n_87),
.B2(n_6),
.Y(n_116)
);

INVx4_ASAP7_75t_L g97 ( 
.A(n_78),
.Y(n_97)
);

INVx3_ASAP7_75t_L g110 ( 
.A(n_97),
.Y(n_110)
);

AOI22xp5_ASAP7_75t_SL g99 ( 
.A1(n_96),
.A2(n_72),
.B1(n_66),
.B2(n_67),
.Y(n_99)
);

OR2x2_ASAP7_75t_L g128 ( 
.A(n_99),
.B(n_116),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_SL g100 ( 
.A(n_85),
.B(n_58),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_L g133 ( 
.A(n_100),
.B(n_109),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_L g123 ( 
.A(n_101),
.B(n_105),
.Y(n_123)
);

CKINVDCx20_ASAP7_75t_R g102 ( 
.A(n_84),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_SL g121 ( 
.A(n_102),
.B(n_115),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_SL g126 ( 
.A(n_106),
.B(n_107),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_91),
.B(n_57),
.Y(n_107)
);

AOI22xp5_ASAP7_75t_L g122 ( 
.A1(n_108),
.A2(n_113),
.B1(n_27),
.B2(n_43),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_88),
.B(n_1),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_97),
.B(n_1),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_L g137 ( 
.A(n_111),
.B(n_114),
.Y(n_137)
);

XNOR2xp5_ASAP7_75t_SL g138 ( 
.A(n_112),
.B(n_21),
.Y(n_138)
);

OAI22xp5_ASAP7_75t_L g113 ( 
.A1(n_98),
.A2(n_26),
.B1(n_47),
.B2(n_44),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_L g114 ( 
.A(n_84),
.B(n_3),
.Y(n_114)
);

CKINVDCx20_ASAP7_75t_R g115 ( 
.A(n_98),
.Y(n_115)
);

AO21x1_ASAP7_75t_L g124 ( 
.A1(n_116),
.A2(n_117),
.B(n_119),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_L g117 ( 
.A(n_94),
.B(n_4),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_SL g118 ( 
.A(n_85),
.B(n_4),
.Y(n_118)
);

OAI21xp5_ASAP7_75t_L g129 ( 
.A1(n_118),
.A2(n_7),
.B(n_9),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_L g119 ( 
.A(n_92),
.B(n_5),
.Y(n_119)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_103),
.Y(n_120)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_120),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_L g145 ( 
.A(n_122),
.B(n_129),
.Y(n_145)
);

XOR2xp5_ASAP7_75t_L g125 ( 
.A(n_99),
.B(n_24),
.Y(n_125)
);

MAJIxp5_ASAP7_75t_L g140 ( 
.A(n_125),
.B(n_136),
.C(n_22),
.Y(n_140)
);

AOI22xp5_ASAP7_75t_SL g127 ( 
.A1(n_116),
.A2(n_6),
.B1(n_7),
.B2(n_9),
.Y(n_127)
);

XNOR2xp5_ASAP7_75t_L g148 ( 
.A(n_127),
.B(n_135),
.Y(n_148)
);

OAI21xp5_ASAP7_75t_SL g143 ( 
.A1(n_128),
.A2(n_30),
.B(n_33),
.Y(n_143)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_110),
.Y(n_130)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_130),
.Y(n_149)
);

INVxp67_ASAP7_75t_L g131 ( 
.A(n_104),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_L g142 ( 
.A(n_131),
.B(n_132),
.Y(n_142)
);

INVx1_ASAP7_75t_SL g132 ( 
.A(n_104),
.Y(n_132)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_106),
.Y(n_134)
);

CKINVDCx20_ASAP7_75t_R g144 ( 
.A(n_134),
.Y(n_144)
);

OAI22xp5_ASAP7_75t_SL g135 ( 
.A1(n_99),
.A2(n_10),
.B1(n_12),
.B2(n_14),
.Y(n_135)
);

MAJIxp5_ASAP7_75t_L g136 ( 
.A(n_112),
.B(n_16),
.C(n_20),
.Y(n_136)
);

FAx1_ASAP7_75t_SL g141 ( 
.A(n_138),
.B(n_50),
.CI(n_32),
.CON(n_141),
.SN(n_141)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_103),
.Y(n_139)
);

XNOR2xp5_ASAP7_75t_L g150 ( 
.A(n_139),
.B(n_36),
.Y(n_150)
);

XNOR2xp5_ASAP7_75t_L g154 ( 
.A(n_140),
.B(n_141),
.Y(n_154)
);

AOI22xp5_ASAP7_75t_SL g152 ( 
.A1(n_143),
.A2(n_132),
.B1(n_131),
.B2(n_125),
.Y(n_152)
);

XOR2xp5_ASAP7_75t_L g147 ( 
.A(n_138),
.B(n_34),
.Y(n_147)
);

MAJIxp5_ASAP7_75t_L g157 ( 
.A(n_147),
.B(n_150),
.C(n_151),
.Y(n_157)
);

MAJIxp5_ASAP7_75t_L g151 ( 
.A(n_126),
.B(n_42),
.C(n_37),
.Y(n_151)
);

XNOR2xp5_ASAP7_75t_L g161 ( 
.A(n_152),
.B(n_137),
.Y(n_161)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_146),
.Y(n_153)
);

OAI21xp33_ASAP7_75t_L g159 ( 
.A1(n_153),
.A2(n_155),
.B(n_156),
.Y(n_159)
);

CKINVDCx20_ASAP7_75t_R g155 ( 
.A(n_142),
.Y(n_155)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_149),
.Y(n_156)
);

A2O1A1O1Ixp25_ASAP7_75t_L g158 ( 
.A1(n_144),
.A2(n_124),
.B(n_145),
.C(n_128),
.D(n_121),
.Y(n_158)
);

A2O1A1Ixp33_ASAP7_75t_SL g160 ( 
.A1(n_158),
.A2(n_124),
.B(n_148),
.C(n_141),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_L g162 ( 
.A(n_160),
.B(n_154),
.Y(n_162)
);

AOI21xp5_ASAP7_75t_L g163 ( 
.A1(n_161),
.A2(n_157),
.B(n_123),
.Y(n_163)
);

MAJIxp5_ASAP7_75t_L g164 ( 
.A(n_162),
.B(n_163),
.C(n_133),
.Y(n_164)
);

OAI21xp5_ASAP7_75t_L g165 ( 
.A1(n_164),
.A2(n_142),
.B(n_159),
.Y(n_165)
);

HB1xp67_ASAP7_75t_L g166 ( 
.A(n_165),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_SL g167 ( 
.A(n_166),
.B(n_41),
.Y(n_167)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_167),
.Y(n_168)
);


endmodule