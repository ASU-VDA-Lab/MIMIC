module fake_jpeg_4976_n_20 (n_0, n_2, n_1, n_20);

input n_0;
input n_2;
input n_1;

output n_20;

wire n_13;
wire n_10;
wire n_6;
wire n_14;
wire n_19;
wire n_18;
wire n_4;
wire n_16;
wire n_3;
wire n_9;
wire n_5;
wire n_11;
wire n_17;
wire n_12;
wire n_8;
wire n_15;
wire n_7;

BUFx4f_ASAP7_75t_L g3 ( 
.A(n_2),
.Y(n_3)
);

INVx3_ASAP7_75t_L g4 ( 
.A(n_2),
.Y(n_4)
);

NOR2xp33_ASAP7_75t_SL g5 ( 
.A(n_1),
.B(n_0),
.Y(n_5)
);

CKINVDCx20_ASAP7_75t_R g6 ( 
.A(n_0),
.Y(n_6)
);

INVx1_ASAP7_75t_L g7 ( 
.A(n_5),
.Y(n_7)
);

INVx1_ASAP7_75t_L g11 ( 
.A(n_7),
.Y(n_11)
);

NAND2xp5_ASAP7_75t_L g8 ( 
.A(n_6),
.B(n_0),
.Y(n_8)
);

CKINVDCx20_ASAP7_75t_R g10 ( 
.A(n_8),
.Y(n_10)
);

NAND2xp5_ASAP7_75t_L g9 ( 
.A(n_6),
.B(n_1),
.Y(n_9)
);

NAND2xp5_ASAP7_75t_L g12 ( 
.A(n_10),
.B(n_8),
.Y(n_12)
);

NAND2xp5_ASAP7_75t_SL g15 ( 
.A(n_12),
.B(n_13),
.Y(n_15)
);

XNOR2xp5_ASAP7_75t_L g13 ( 
.A(n_10),
.B(n_9),
.Y(n_13)
);

XOR2x1_ASAP7_75t_SL g14 ( 
.A(n_13),
.B(n_3),
.Y(n_14)
);

NOR3xp33_ASAP7_75t_SL g16 ( 
.A(n_14),
.B(n_3),
.C(n_15),
.Y(n_16)
);

OAI21xp5_ASAP7_75t_L g18 ( 
.A1(n_16),
.A2(n_17),
.B(n_11),
.Y(n_18)
);

HB1xp67_ASAP7_75t_L g17 ( 
.A(n_14),
.Y(n_17)
);

AOI22xp5_ASAP7_75t_SL g19 ( 
.A1(n_18),
.A2(n_11),
.B1(n_4),
.B2(n_3),
.Y(n_19)
);

OAI21xp5_ASAP7_75t_L g20 ( 
.A1(n_19),
.A2(n_4),
.B(n_1),
.Y(n_20)
);


endmodule