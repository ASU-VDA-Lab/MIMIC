module fake_jpeg_24295_n_258 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_258);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_258;

wire n_159;
wire n_117;
wire n_253;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_251;
wire n_252;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_223;
wire n_187;
wire n_21;
wire n_57;
wire n_234;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_44;
wire n_24;
wire n_143;
wire n_202;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_217;
wire n_216;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_7),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_0),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_11),
.Y(n_18)
);

BUFx16f_ASAP7_75t_L g19 ( 
.A(n_1),
.Y(n_19)
);

INVx2_ASAP7_75t_L g20 ( 
.A(n_4),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_12),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_1),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_1),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_11),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_12),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_3),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_6),
.Y(n_27)
);

INVx11_ASAP7_75t_SL g28 ( 
.A(n_7),
.Y(n_28)
);

BUFx8_ASAP7_75t_L g29 ( 
.A(n_9),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_15),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_7),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_1),
.Y(n_32)
);

INVx4_ASAP7_75t_L g33 ( 
.A(n_29),
.Y(n_33)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_33),
.Y(n_44)
);

AND2x2_ASAP7_75t_SL g34 ( 
.A(n_20),
.B(n_0),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_34),
.B(n_35),
.Y(n_48)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_16),
.Y(n_35)
);

BUFx12f_ASAP7_75t_L g36 ( 
.A(n_29),
.Y(n_36)
);

BUFx3_ASAP7_75t_L g42 ( 
.A(n_36),
.Y(n_42)
);

INVx2_ASAP7_75t_L g37 ( 
.A(n_19),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g49 ( 
.A(n_37),
.B(n_29),
.Y(n_49)
);

BUFx12f_ASAP7_75t_L g38 ( 
.A(n_29),
.Y(n_38)
);

INVx4_ASAP7_75t_L g53 ( 
.A(n_38),
.Y(n_53)
);

BUFx3_ASAP7_75t_L g39 ( 
.A(n_29),
.Y(n_39)
);

INVx3_ASAP7_75t_L g54 ( 
.A(n_39),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_23),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_40),
.Y(n_50)
);

AOI22xp5_ASAP7_75t_L g41 ( 
.A1(n_34),
.A2(n_20),
.B1(n_22),
.B2(n_26),
.Y(n_41)
);

OAI22xp5_ASAP7_75t_L g74 ( 
.A1(n_41),
.A2(n_34),
.B1(n_32),
.B2(n_26),
.Y(n_74)
);

INVx2_ASAP7_75t_L g43 ( 
.A(n_39),
.Y(n_43)
);

INVx6_ASAP7_75t_L g76 ( 
.A(n_43),
.Y(n_76)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_33),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_45),
.B(n_47),
.Y(n_65)
);

INVx3_ASAP7_75t_L g46 ( 
.A(n_39),
.Y(n_46)
);

BUFx2_ASAP7_75t_SL g57 ( 
.A(n_46),
.Y(n_57)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_33),
.Y(n_47)
);

CKINVDCx16_ASAP7_75t_R g64 ( 
.A(n_49),
.Y(n_64)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_33),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_L g56 ( 
.A(n_51),
.B(n_34),
.Y(n_56)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_35),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_SL g60 ( 
.A(n_52),
.B(n_35),
.Y(n_60)
);

AOI22xp33_ASAP7_75t_SL g55 ( 
.A1(n_36),
.A2(n_28),
.B1(n_20),
.B2(n_18),
.Y(n_55)
);

AOI22xp33_ASAP7_75t_SL g69 ( 
.A1(n_55),
.A2(n_36),
.B1(n_38),
.B2(n_28),
.Y(n_69)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_56),
.Y(n_91)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_41),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_SL g98 ( 
.A(n_58),
.B(n_60),
.Y(n_98)
);

AOI22xp33_ASAP7_75t_L g59 ( 
.A1(n_48),
.A2(n_25),
.B1(n_27),
.B2(n_30),
.Y(n_59)
);

OAI22xp5_ASAP7_75t_L g93 ( 
.A1(n_59),
.A2(n_69),
.B1(n_72),
.B2(n_82),
.Y(n_93)
);

AND2x2_ASAP7_75t_L g61 ( 
.A(n_48),
.B(n_34),
.Y(n_61)
);

OR2x4_ASAP7_75t_L g105 ( 
.A(n_61),
.B(n_40),
.Y(n_105)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_49),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_62),
.B(n_63),
.Y(n_90)
);

CKINVDCx20_ASAP7_75t_R g63 ( 
.A(n_52),
.Y(n_63)
);

INVx8_ASAP7_75t_L g66 ( 
.A(n_50),
.Y(n_66)
);

INVx2_ASAP7_75t_L g86 ( 
.A(n_66),
.Y(n_86)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_53),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_67),
.B(n_68),
.Y(n_104)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_53),
.Y(n_68)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_53),
.Y(n_70)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_70),
.Y(n_95)
);

OAI21xp5_ASAP7_75t_L g71 ( 
.A1(n_44),
.A2(n_34),
.B(n_38),
.Y(n_71)
);

CKINVDCx14_ASAP7_75t_R g87 ( 
.A(n_71),
.Y(n_87)
);

AOI22xp33_ASAP7_75t_SL g72 ( 
.A1(n_54),
.A2(n_24),
.B1(n_18),
.B2(n_21),
.Y(n_72)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_42),
.Y(n_73)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_73),
.Y(n_97)
);

AOI22xp5_ASAP7_75t_L g96 ( 
.A1(n_74),
.A2(n_77),
.B1(n_83),
.B2(n_84),
.Y(n_96)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_42),
.Y(n_75)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_75),
.Y(n_108)
);

AO22x2_ASAP7_75t_L g77 ( 
.A1(n_42),
.A2(n_36),
.B1(n_38),
.B2(n_34),
.Y(n_77)
);

BUFx5_ASAP7_75t_L g78 ( 
.A(n_46),
.Y(n_78)
);

BUFx12_ASAP7_75t_L g107 ( 
.A(n_78),
.Y(n_107)
);

CKINVDCx20_ASAP7_75t_R g79 ( 
.A(n_54),
.Y(n_79)
);

NOR3xp33_ASAP7_75t_L g100 ( 
.A(n_79),
.B(n_36),
.C(n_38),
.Y(n_100)
);

INVx4_ASAP7_75t_L g80 ( 
.A(n_54),
.Y(n_80)
);

BUFx6f_ASAP7_75t_L g103 ( 
.A(n_80),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_SL g81 ( 
.A(n_44),
.B(n_25),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g92 ( 
.A(n_81),
.B(n_85),
.Y(n_92)
);

AOI22xp5_ASAP7_75t_L g82 ( 
.A1(n_51),
.A2(n_37),
.B1(n_47),
.B2(n_45),
.Y(n_82)
);

AOI22xp5_ASAP7_75t_L g83 ( 
.A1(n_43),
.A2(n_37),
.B1(n_39),
.B2(n_40),
.Y(n_83)
);

AOI22xp5_ASAP7_75t_L g84 ( 
.A1(n_50),
.A2(n_37),
.B1(n_40),
.B2(n_38),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g85 ( 
.A(n_50),
.B(n_23),
.Y(n_85)
);

CKINVDCx16_ASAP7_75t_R g88 ( 
.A(n_65),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_88),
.B(n_94),
.Y(n_111)
);

AND2x6_ASAP7_75t_L g89 ( 
.A(n_77),
.B(n_38),
.Y(n_89)
);

A2O1A1O1Ixp25_ASAP7_75t_L g132 ( 
.A1(n_89),
.A2(n_83),
.B(n_84),
.C(n_85),
.D(n_76),
.Y(n_132)
);

INVx3_ASAP7_75t_L g94 ( 
.A(n_78),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_61),
.B(n_40),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g113 ( 
.A(n_99),
.B(n_106),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_L g116 ( 
.A(n_100),
.B(n_29),
.Y(n_116)
);

AOI22xp33_ASAP7_75t_L g101 ( 
.A1(n_58),
.A2(n_36),
.B1(n_21),
.B2(n_18),
.Y(n_101)
);

OAI22xp5_ASAP7_75t_SL g124 ( 
.A1(n_101),
.A2(n_110),
.B1(n_24),
.B2(n_31),
.Y(n_124)
);

OR2x2_ASAP7_75t_L g102 ( 
.A(n_63),
.B(n_36),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_SL g122 ( 
.A(n_102),
.B(n_81),
.Y(n_122)
);

OAI21xp5_ASAP7_75t_SL g117 ( 
.A1(n_105),
.A2(n_77),
.B(n_71),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_L g106 ( 
.A(n_61),
.B(n_19),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_L g109 ( 
.A(n_56),
.B(n_19),
.Y(n_109)
);

XOR2xp5_ASAP7_75t_L g121 ( 
.A(n_109),
.B(n_82),
.Y(n_121)
);

AOI22xp5_ASAP7_75t_L g110 ( 
.A1(n_74),
.A2(n_24),
.B1(n_31),
.B2(n_21),
.Y(n_110)
);

CKINVDCx16_ASAP7_75t_R g112 ( 
.A(n_104),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_L g157 ( 
.A(n_112),
.B(n_126),
.Y(n_157)
);

OAI21xp5_ASAP7_75t_L g114 ( 
.A1(n_87),
.A2(n_105),
.B(n_98),
.Y(n_114)
);

MAJIxp5_ASAP7_75t_SL g145 ( 
.A(n_114),
.B(n_128),
.C(n_132),
.Y(n_145)
);

OA21x2_ASAP7_75t_L g115 ( 
.A1(n_102),
.A2(n_77),
.B(n_96),
.Y(n_115)
);

OAI21xp5_ASAP7_75t_SL g140 ( 
.A1(n_115),
.A2(n_116),
.B(n_117),
.Y(n_140)
);

AOI22xp5_ASAP7_75t_L g118 ( 
.A1(n_93),
.A2(n_77),
.B1(n_64),
.B2(n_62),
.Y(n_118)
);

OAI22xp5_ASAP7_75t_L g155 ( 
.A1(n_118),
.A2(n_86),
.B1(n_66),
.B2(n_68),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_L g119 ( 
.A(n_94),
.B(n_79),
.Y(n_119)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_119),
.Y(n_138)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_90),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_L g160 ( 
.A(n_120),
.B(n_125),
.Y(n_160)
);

XNOR2xp5_ASAP7_75t_L g148 ( 
.A(n_121),
.B(n_23),
.Y(n_148)
);

OAI21xp5_ASAP7_75t_SL g144 ( 
.A1(n_122),
.A2(n_133),
.B(n_134),
.Y(n_144)
);

XOR2xp5_ASAP7_75t_L g123 ( 
.A(n_99),
.B(n_64),
.Y(n_123)
);

MAJIxp5_ASAP7_75t_L g137 ( 
.A(n_123),
.B(n_130),
.C(n_136),
.Y(n_137)
);

OAI22xp33_ASAP7_75t_SL g142 ( 
.A1(n_124),
.A2(n_135),
.B1(n_80),
.B2(n_76),
.Y(n_142)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_92),
.Y(n_125)
);

CKINVDCx16_ASAP7_75t_R g126 ( 
.A(n_103),
.Y(n_126)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_92),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_L g162 ( 
.A(n_127),
.B(n_129),
.Y(n_162)
);

NOR2xp67_ASAP7_75t_SL g128 ( 
.A(n_89),
.B(n_57),
.Y(n_128)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_110),
.Y(n_129)
);

MAJIxp5_ASAP7_75t_L g130 ( 
.A(n_106),
.B(n_91),
.C(n_109),
.Y(n_130)
);

CKINVDCx20_ASAP7_75t_R g131 ( 
.A(n_103),
.Y(n_131)
);

CKINVDCx20_ASAP7_75t_R g139 ( 
.A(n_131),
.Y(n_139)
);

AND2x2_ASAP7_75t_L g133 ( 
.A(n_96),
.B(n_0),
.Y(n_133)
);

CKINVDCx20_ASAP7_75t_R g134 ( 
.A(n_103),
.Y(n_134)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_95),
.Y(n_135)
);

MAJIxp5_ASAP7_75t_L g136 ( 
.A(n_91),
.B(n_67),
.C(n_70),
.Y(n_136)
);

OAI22xp5_ASAP7_75t_SL g141 ( 
.A1(n_128),
.A2(n_93),
.B1(n_86),
.B2(n_76),
.Y(n_141)
);

AOI22xp5_ASAP7_75t_L g164 ( 
.A1(n_141),
.A2(n_155),
.B1(n_124),
.B2(n_129),
.Y(n_164)
);

AOI22xp33_ASAP7_75t_L g165 ( 
.A1(n_142),
.A2(n_66),
.B1(n_131),
.B2(n_134),
.Y(n_165)
);

CKINVDCx16_ASAP7_75t_R g143 ( 
.A(n_111),
.Y(n_143)
);

NOR2xp33_ASAP7_75t_L g174 ( 
.A(n_143),
.B(n_146),
.Y(n_174)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_136),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_L g147 ( 
.A(n_125),
.B(n_60),
.Y(n_147)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_147),
.Y(n_168)
);

XNOR2xp5_ASAP7_75t_SL g184 ( 
.A(n_148),
.B(n_150),
.Y(n_184)
);

XNOR2xp5_ASAP7_75t_L g149 ( 
.A(n_123),
.B(n_95),
.Y(n_149)
);

MAJIxp5_ASAP7_75t_L g170 ( 
.A(n_149),
.B(n_151),
.C(n_154),
.Y(n_170)
);

XNOR2xp5_ASAP7_75t_SL g150 ( 
.A(n_118),
.B(n_19),
.Y(n_150)
);

XNOR2xp5_ASAP7_75t_L g151 ( 
.A(n_114),
.B(n_108),
.Y(n_151)
);

FAx1_ASAP7_75t_SL g152 ( 
.A(n_130),
.B(n_97),
.CI(n_108),
.CON(n_152),
.SN(n_152)
);

NOR2xp33_ASAP7_75t_L g176 ( 
.A(n_152),
.B(n_153),
.Y(n_176)
);

BUFx5_ASAP7_75t_L g153 ( 
.A(n_126),
.Y(n_153)
);

XNOR2xp5_ASAP7_75t_L g154 ( 
.A(n_113),
.B(n_97),
.Y(n_154)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_135),
.Y(n_156)
);

NOR2xp33_ASAP7_75t_L g183 ( 
.A(n_156),
.B(n_163),
.Y(n_183)
);

XOR2xp5_ASAP7_75t_L g158 ( 
.A(n_117),
.B(n_19),
.Y(n_158)
);

MAJIxp5_ASAP7_75t_L g177 ( 
.A(n_158),
.B(n_159),
.C(n_161),
.Y(n_177)
);

XOR2xp5_ASAP7_75t_L g159 ( 
.A(n_113),
.B(n_23),
.Y(n_159)
);

MAJIxp5_ASAP7_75t_L g161 ( 
.A(n_121),
.B(n_75),
.C(n_73),
.Y(n_161)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_122),
.Y(n_163)
);

OAI22xp5_ASAP7_75t_SL g187 ( 
.A1(n_164),
.A2(n_165),
.B1(n_166),
.B2(n_167),
.Y(n_187)
);

AOI22xp5_ASAP7_75t_L g166 ( 
.A1(n_141),
.A2(n_115),
.B1(n_132),
.B2(n_133),
.Y(n_166)
);

OAI22xp5_ASAP7_75t_SL g167 ( 
.A1(n_145),
.A2(n_115),
.B1(n_127),
.B2(n_133),
.Y(n_167)
);

O2A1O1Ixp33_ASAP7_75t_L g169 ( 
.A1(n_162),
.A2(n_115),
.B(n_17),
.C(n_112),
.Y(n_169)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_169),
.Y(n_191)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_160),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_L g198 ( 
.A(n_171),
.B(n_173),
.Y(n_198)
);

AND2x2_ASAP7_75t_L g172 ( 
.A(n_151),
.B(n_0),
.Y(n_172)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_172),
.Y(n_196)
);

AOI22xp5_ASAP7_75t_L g173 ( 
.A1(n_145),
.A2(n_161),
.B1(n_140),
.B2(n_150),
.Y(n_173)
);

BUFx12_ASAP7_75t_L g175 ( 
.A(n_153),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_SL g200 ( 
.A(n_175),
.B(n_178),
.Y(n_200)
);

OAI22xp5_ASAP7_75t_SL g178 ( 
.A1(n_140),
.A2(n_120),
.B1(n_32),
.B2(n_22),
.Y(n_178)
);

MAJIxp5_ASAP7_75t_L g179 ( 
.A(n_137),
.B(n_107),
.C(n_32),
.Y(n_179)
);

MAJIxp5_ASAP7_75t_L g192 ( 
.A(n_179),
.B(n_138),
.C(n_139),
.Y(n_192)
);

AOI22xp5_ASAP7_75t_L g180 ( 
.A1(n_137),
.A2(n_27),
.B1(n_25),
.B2(n_26),
.Y(n_180)
);

AOI22xp5_ASAP7_75t_SL g201 ( 
.A1(n_180),
.A2(n_185),
.B1(n_17),
.B2(n_10),
.Y(n_201)
);

OAI32xp33_ASAP7_75t_L g181 ( 
.A1(n_158),
.A2(n_31),
.A3(n_22),
.B1(n_4),
.B2(n_2),
.Y(n_181)
);

XOR2xp5_ASAP7_75t_L g189 ( 
.A(n_181),
.B(n_144),
.Y(n_189)
);

OAI21xp5_ASAP7_75t_L g182 ( 
.A1(n_147),
.A2(n_27),
.B(n_17),
.Y(n_182)
);

AOI21xp5_ASAP7_75t_SL g190 ( 
.A1(n_182),
.A2(n_186),
.B(n_144),
.Y(n_190)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_157),
.Y(n_185)
);

NOR2xp33_ASAP7_75t_SL g186 ( 
.A(n_159),
.B(n_16),
.Y(n_186)
);

XNOR2xp5_ASAP7_75t_L g188 ( 
.A(n_184),
.B(n_177),
.Y(n_188)
);

XOR2xp5_ASAP7_75t_L g211 ( 
.A(n_188),
.B(n_195),
.Y(n_211)
);

NAND2xp5_ASAP7_75t_SL g215 ( 
.A(n_189),
.B(n_172),
.Y(n_215)
);

NOR2xp33_ASAP7_75t_SL g210 ( 
.A(n_190),
.B(n_202),
.Y(n_210)
);

MAJIxp5_ASAP7_75t_L g212 ( 
.A(n_192),
.B(n_193),
.C(n_194),
.Y(n_212)
);

MAJIxp5_ASAP7_75t_L g193 ( 
.A(n_177),
.B(n_149),
.C(n_148),
.Y(n_193)
);

MAJIxp5_ASAP7_75t_L g194 ( 
.A(n_179),
.B(n_152),
.C(n_154),
.Y(n_194)
);

MAJIxp5_ASAP7_75t_L g195 ( 
.A(n_170),
.B(n_152),
.C(n_107),
.Y(n_195)
);

XNOR2xp5_ASAP7_75t_SL g197 ( 
.A(n_173),
.B(n_11),
.Y(n_197)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_197),
.Y(n_207)
);

MAJIxp5_ASAP7_75t_L g199 ( 
.A(n_170),
.B(n_107),
.C(n_30),
.Y(n_199)
);

NOR2xp33_ASAP7_75t_L g204 ( 
.A(n_199),
.B(n_201),
.Y(n_204)
);

MAJIxp5_ASAP7_75t_L g202 ( 
.A(n_184),
.B(n_107),
.C(n_9),
.Y(n_202)
);

XOR2xp5_ASAP7_75t_L g203 ( 
.A(n_167),
.B(n_9),
.Y(n_203)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_203),
.Y(n_216)
);

AOI21xp5_ASAP7_75t_SL g205 ( 
.A1(n_190),
.A2(n_176),
.B(n_168),
.Y(n_205)
);

AOI21xp5_ASAP7_75t_L g224 ( 
.A1(n_205),
.A2(n_213),
.B(n_210),
.Y(n_224)
);

OAI22xp5_ASAP7_75t_L g206 ( 
.A1(n_198),
.A2(n_164),
.B1(n_166),
.B2(n_171),
.Y(n_206)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_206),
.Y(n_228)
);

HB1xp67_ASAP7_75t_L g208 ( 
.A(n_192),
.Y(n_208)
);

HB1xp67_ASAP7_75t_L g225 ( 
.A(n_208),
.Y(n_225)
);

AOI21x1_ASAP7_75t_L g209 ( 
.A1(n_189),
.A2(n_169),
.B(n_168),
.Y(n_209)
);

OAI22x1_ASAP7_75t_L g220 ( 
.A1(n_209),
.A2(n_217),
.B1(n_200),
.B2(n_203),
.Y(n_220)
);

INVxp67_ASAP7_75t_L g213 ( 
.A(n_187),
.Y(n_213)
);

OAI22xp5_ASAP7_75t_L g214 ( 
.A1(n_191),
.A2(n_174),
.B1(n_185),
.B2(n_183),
.Y(n_214)
);

NAND2xp5_ASAP7_75t_SL g222 ( 
.A(n_214),
.B(n_175),
.Y(n_222)
);

MAJIxp5_ASAP7_75t_L g221 ( 
.A(n_215),
.B(n_195),
.C(n_182),
.Y(n_221)
);

AOI22xp5_ASAP7_75t_L g217 ( 
.A1(n_196),
.A2(n_178),
.B1(n_186),
.B2(n_181),
.Y(n_217)
);

NAND3xp33_ASAP7_75t_L g218 ( 
.A(n_197),
.B(n_172),
.C(n_180),
.Y(n_218)
);

NOR2xp33_ASAP7_75t_L g223 ( 
.A(n_218),
.B(n_175),
.Y(n_223)
);

XNOR2xp5_ASAP7_75t_L g219 ( 
.A(n_212),
.B(n_193),
.Y(n_219)
);

XNOR2xp5_ASAP7_75t_L g236 ( 
.A(n_219),
.B(n_221),
.Y(n_236)
);

A2O1A1O1Ixp25_ASAP7_75t_L g237 ( 
.A1(n_220),
.A2(n_223),
.B(n_216),
.C(n_211),
.D(n_10),
.Y(n_237)
);

NAND2xp5_ASAP7_75t_L g233 ( 
.A(n_222),
.B(n_204),
.Y(n_233)
);

CKINVDCx20_ASAP7_75t_R g231 ( 
.A(n_224),
.Y(n_231)
);

NOR2xp33_ASAP7_75t_L g226 ( 
.A(n_205),
.B(n_8),
.Y(n_226)
);

NAND2xp5_ASAP7_75t_SL g235 ( 
.A(n_226),
.B(n_10),
.Y(n_235)
);

NAND2xp5_ASAP7_75t_L g227 ( 
.A(n_217),
.B(n_8),
.Y(n_227)
);

NAND2xp5_ASAP7_75t_L g238 ( 
.A(n_227),
.B(n_8),
.Y(n_238)
);

MAJIxp5_ASAP7_75t_L g229 ( 
.A(n_212),
.B(n_2),
.C(n_3),
.Y(n_229)
);

MAJIxp5_ASAP7_75t_L g232 ( 
.A(n_229),
.B(n_216),
.C(n_207),
.Y(n_232)
);

NOR2xp33_ASAP7_75t_L g230 ( 
.A(n_228),
.B(n_213),
.Y(n_230)
);

CKINVDCx20_ASAP7_75t_R g239 ( 
.A(n_230),
.Y(n_239)
);

AOI21xp5_ASAP7_75t_L g245 ( 
.A1(n_232),
.A2(n_237),
.B(n_6),
.Y(n_245)
);

NAND2xp5_ASAP7_75t_L g241 ( 
.A(n_233),
.B(n_235),
.Y(n_241)
);

AND2x2_ASAP7_75t_L g234 ( 
.A(n_220),
.B(n_209),
.Y(n_234)
);

NAND3xp33_ASAP7_75t_SL g243 ( 
.A(n_234),
.B(n_225),
.C(n_12),
.Y(n_243)
);

NOR2xp33_ASAP7_75t_L g240 ( 
.A(n_238),
.B(n_231),
.Y(n_240)
);

CKINVDCx20_ASAP7_75t_R g246 ( 
.A(n_240),
.Y(n_246)
);

AOI22xp5_ASAP7_75t_L g242 ( 
.A1(n_234),
.A2(n_225),
.B1(n_229),
.B2(n_211),
.Y(n_242)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_242),
.Y(n_247)
);

AND2x2_ASAP7_75t_L g249 ( 
.A(n_243),
.B(n_13),
.Y(n_249)
);

NOR2xp33_ASAP7_75t_L g244 ( 
.A(n_236),
.B(n_6),
.Y(n_244)
);

MAJIxp5_ASAP7_75t_L g248 ( 
.A(n_244),
.B(n_245),
.C(n_241),
.Y(n_248)
);

AOI21xp5_ASAP7_75t_L g251 ( 
.A1(n_248),
.A2(n_250),
.B(n_243),
.Y(n_251)
);

AOI322xp5_ASAP7_75t_L g253 ( 
.A1(n_249),
.A2(n_5),
.A3(n_13),
.B1(n_14),
.B2(n_15),
.C1(n_3),
.C2(n_4),
.Y(n_253)
);

MAJIxp5_ASAP7_75t_L g250 ( 
.A(n_239),
.B(n_232),
.C(n_237),
.Y(n_250)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_251),
.Y(n_254)
);

AOI322xp5_ASAP7_75t_L g252 ( 
.A1(n_246),
.A2(n_5),
.A3(n_13),
.B1(n_14),
.B2(n_15),
.C1(n_3),
.C2(n_4),
.Y(n_252)
);

AOI22xp33_ASAP7_75t_SL g255 ( 
.A1(n_252),
.A2(n_253),
.B1(n_247),
.B2(n_5),
.Y(n_255)
);

MAJIxp5_ASAP7_75t_L g256 ( 
.A(n_255),
.B(n_14),
.C(n_2),
.Y(n_256)
);

XNOR2xp5_ASAP7_75t_L g257 ( 
.A(n_256),
.B(n_2),
.Y(n_257)
);

XNOR2xp5_ASAP7_75t_L g258 ( 
.A(n_257),
.B(n_254),
.Y(n_258)
);


endmodule