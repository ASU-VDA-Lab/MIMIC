module fake_jpeg_21581_n_77 (n_3, n_2, n_1, n_0, n_4, n_6, n_5, n_7, n_77);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_6;
input n_5;
input n_7;

output n_77;

wire n_10;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_59;
wire n_65;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_28;
wire n_38;
wire n_26;
wire n_74;
wire n_31;
wire n_29;
wire n_50;
wire n_15;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_69;
wire n_27;
wire n_40;
wire n_71;
wire n_30;
wire n_24;
wire n_44;
wire n_17;
wire n_25;
wire n_75;
wire n_37;
wire n_70;
wire n_66;
wire n_61;
wire n_45;
wire n_18;
wire n_20;
wire n_68;
wire n_52;
wire n_58;
wire n_41;
wire n_60;
wire n_63;
wire n_34;
wire n_39;
wire n_72;
wire n_11;
wire n_56;
wire n_12;
wire n_8;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_22;
wire n_35;
wire n_48;
wire n_46;
wire n_9;
wire n_36;
wire n_62;
wire n_43;
wire n_32;

INVx1_ASAP7_75t_L g8 ( 
.A(n_6),
.Y(n_8)
);

INVx1_ASAP7_75t_L g9 ( 
.A(n_1),
.Y(n_9)
);

CKINVDCx20_ASAP7_75t_R g10 ( 
.A(n_6),
.Y(n_10)
);

CKINVDCx20_ASAP7_75t_R g11 ( 
.A(n_4),
.Y(n_11)
);

BUFx12f_ASAP7_75t_L g12 ( 
.A(n_5),
.Y(n_12)
);

INVx6_ASAP7_75t_SL g13 ( 
.A(n_5),
.Y(n_13)
);

CKINVDCx20_ASAP7_75t_R g14 ( 
.A(n_2),
.Y(n_14)
);

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_2),
.Y(n_15)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_4),
.Y(n_16)
);

BUFx12f_ASAP7_75t_L g17 ( 
.A(n_12),
.Y(n_17)
);

BUFx3_ASAP7_75t_L g24 ( 
.A(n_17),
.Y(n_24)
);

INVx4_ASAP7_75t_L g18 ( 
.A(n_12),
.Y(n_18)
);

INVx3_ASAP7_75t_L g22 ( 
.A(n_18),
.Y(n_22)
);

BUFx2_ASAP7_75t_L g19 ( 
.A(n_12),
.Y(n_19)
);

NOR2xp33_ASAP7_75t_L g23 ( 
.A(n_19),
.B(n_13),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_12),
.Y(n_20)
);

INVx3_ASAP7_75t_L g26 ( 
.A(n_20),
.Y(n_26)
);

NAND2xp5_ASAP7_75t_L g21 ( 
.A(n_12),
.B(n_0),
.Y(n_21)
);

NAND2xp5_ASAP7_75t_L g25 ( 
.A(n_21),
.B(n_15),
.Y(n_25)
);

AO21x1_ASAP7_75t_L g29 ( 
.A1(n_23),
.A2(n_13),
.B(n_19),
.Y(n_29)
);

XOR2xp5_ASAP7_75t_L g33 ( 
.A(n_25),
.B(n_27),
.Y(n_33)
);

MAJIxp5_ASAP7_75t_L g27 ( 
.A(n_21),
.B(n_9),
.C(n_15),
.Y(n_27)
);

INVx13_ASAP7_75t_L g28 ( 
.A(n_24),
.Y(n_28)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_28),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g38 ( 
.A(n_29),
.B(n_32),
.Y(n_38)
);

OAI22xp5_ASAP7_75t_SL g30 ( 
.A1(n_25),
.A2(n_18),
.B1(n_14),
.B2(n_9),
.Y(n_30)
);

OAI22xp5_ASAP7_75t_L g40 ( 
.A1(n_30),
.A2(n_35),
.B1(n_26),
.B2(n_10),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_24),
.Y(n_31)
);

INVx4_ASAP7_75t_L g45 ( 
.A(n_31),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g32 ( 
.A(n_27),
.B(n_11),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_22),
.Y(n_34)
);

AOI22xp33_ASAP7_75t_SL g43 ( 
.A1(n_34),
.A2(n_36),
.B1(n_17),
.B2(n_20),
.Y(n_43)
);

OAI22xp5_ASAP7_75t_SL g35 ( 
.A1(n_26),
.A2(n_18),
.B1(n_14),
.B2(n_19),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_22),
.Y(n_36)
);

INVxp67_ASAP7_75t_L g37 ( 
.A(n_35),
.Y(n_37)
);

NAND2xp5_ASAP7_75t_SL g50 ( 
.A(n_37),
.B(n_39),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_L g39 ( 
.A(n_33),
.B(n_19),
.Y(n_39)
);

AND2x2_ASAP7_75t_L g49 ( 
.A(n_40),
.B(n_16),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_L g41 ( 
.A(n_33),
.B(n_17),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_41),
.B(n_42),
.Y(n_52)
);

INVx3_ASAP7_75t_L g42 ( 
.A(n_28),
.Y(n_42)
);

CKINVDCx16_ASAP7_75t_R g54 ( 
.A(n_43),
.Y(n_54)
);

AOI21xp5_ASAP7_75t_SL g46 ( 
.A1(n_30),
.A2(n_8),
.B(n_16),
.Y(n_46)
);

OAI21xp5_ASAP7_75t_L g51 ( 
.A1(n_46),
.A2(n_10),
.B(n_11),
.Y(n_51)
);

INVxp33_ASAP7_75t_L g47 ( 
.A(n_45),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g57 ( 
.A(n_47),
.B(n_45),
.Y(n_57)
);

INVxp67_ASAP7_75t_L g48 ( 
.A(n_38),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_L g56 ( 
.A(n_48),
.B(n_51),
.Y(n_56)
);

AOI22xp5_ASAP7_75t_L g59 ( 
.A1(n_49),
.A2(n_44),
.B1(n_42),
.B2(n_7),
.Y(n_59)
);

NOR3xp33_ASAP7_75t_L g53 ( 
.A(n_46),
.B(n_29),
.C(n_37),
.Y(n_53)
);

NOR3xp33_ASAP7_75t_L g60 ( 
.A(n_53),
.B(n_39),
.C(n_17),
.Y(n_60)
);

MAJIxp5_ASAP7_75t_L g55 ( 
.A(n_41),
.B(n_17),
.C(n_20),
.Y(n_55)
);

MAJIxp5_ASAP7_75t_L g61 ( 
.A(n_55),
.B(n_20),
.C(n_31),
.Y(n_61)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_57),
.Y(n_64)
);

AND2x2_ASAP7_75t_L g58 ( 
.A(n_52),
.B(n_8),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_L g65 ( 
.A(n_58),
.B(n_59),
.Y(n_65)
);

INVx11_ASAP7_75t_L g62 ( 
.A(n_60),
.Y(n_62)
);

MAJIxp5_ASAP7_75t_L g63 ( 
.A(n_61),
.B(n_54),
.C(n_50),
.Y(n_63)
);

AOI22xp5_ASAP7_75t_SL g66 ( 
.A1(n_63),
.A2(n_49),
.B1(n_56),
.B2(n_57),
.Y(n_66)
);

MAJIxp5_ASAP7_75t_L g71 ( 
.A(n_66),
.B(n_67),
.C(n_65),
.Y(n_71)
);

OA21x2_ASAP7_75t_SL g67 ( 
.A1(n_62),
.A2(n_7),
.B(n_47),
.Y(n_67)
);

AOI22xp5_ASAP7_75t_L g68 ( 
.A1(n_65),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_68)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_68),
.Y(n_70)
);

INVxp33_ASAP7_75t_L g69 ( 
.A(n_66),
.Y(n_69)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_69),
.Y(n_72)
);

AOI21xp5_ASAP7_75t_L g73 ( 
.A1(n_71),
.A2(n_64),
.B(n_62),
.Y(n_73)
);

AOI322xp5_ASAP7_75t_L g74 ( 
.A1(n_73),
.A2(n_70),
.A3(n_64),
.B1(n_63),
.B2(n_62),
.C1(n_3),
.C2(n_1),
.Y(n_74)
);

CKINVDCx20_ASAP7_75t_R g75 ( 
.A(n_74),
.Y(n_75)
);

AOI22xp33_ASAP7_75t_L g76 ( 
.A1(n_75),
.A2(n_72),
.B1(n_0),
.B2(n_3),
.Y(n_76)
);

XOR2xp5_ASAP7_75t_L g77 ( 
.A(n_76),
.B(n_3),
.Y(n_77)
);


endmodule