module real_jpeg_13826_n_17 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_335, n_7, n_16, n_3, n_10, n_9, n_17);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_335;
input n_7;
input n_16;
input n_3;
input n_10;
input n_9;

output n_17;

wire n_37;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_300;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_199;
wire n_95;
wire n_238;
wire n_67;
wire n_235;
wire n_107;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_123;
wire n_50;
wire n_186;
wire n_137;
wire n_72;
wire n_171;
wire n_151;
wire n_272;
wire n_203;
wire n_198;
wire n_23;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_326;
wire n_80;
wire n_30;
wire n_328;
wire n_149;
wire n_332;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_230;
wire n_128;
wire n_202;
wire n_216;
wire n_127;
wire n_36;
wire n_102;
wire n_81;
wire n_101;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_252;
wire n_310;
wire n_78;
wire n_83;
wire n_288;
wire n_221;
wire n_104;
wire n_153;
wire n_131;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_200;
wire n_214;
wire n_113;
wire n_251;
wire n_139;
wire n_33;
wire n_175;
wire n_156;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_77;
wire n_219;
wire n_122;
wire n_19;
wire n_262;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_20;
wire n_314;
wire n_278;
wire n_103;
wire n_232;
wire n_212;
wire n_284;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_213;
wire n_25;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_331;
wire n_49;
wire n_68;
wire n_146;
wire n_323;
wire n_215;
wire n_176;
wire n_166;
wire n_286;
wire n_312;
wire n_325;
wire n_316;
wire n_307;
wire n_161;
wire n_207;
wire n_237;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_140;
wire n_126;
wire n_120;
wire n_155;
wire n_319;
wire n_93;
wire n_242;
wire n_142;
wire n_76;
wire n_79;
wire n_282;
wire n_147;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_18;
wire n_145;
wire n_266;
wire n_109;
wire n_148;
wire n_196;
wire n_330;
wire n_298;
wire n_333;
wire n_152;
wire n_270;
wire n_159;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_258;
wire n_150;
wire n_41;
wire n_74;
wire n_158;
wire n_204;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_75;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_119;
wire n_283;
wire n_181;
wire n_256;
wire n_253;
wire n_273;
wire n_54;
wire n_168;
wire n_38;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_292;
wire n_64;
wire n_291;
wire n_236;
wire n_276;
wire n_287;
wire n_174;
wire n_255;
wire n_243;
wire n_299;
wire n_56;
wire n_293;
wire n_275;
wire n_227;
wire n_229;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_45;
wire n_313;
wire n_42;
wire n_268;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_143;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_303;
wire n_321;
wire n_100;
wire n_51;
wire n_205;
wire n_261;
wire n_86;
wire n_324;
wire n_70;
wire n_32;
wire n_228;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_133;
wire n_257;
wire n_210;
wire n_206;
wire n_85;
wire n_96;
wire n_308;

BUFx2_ASAP7_75t_L g54 ( 
.A(n_0),
.Y(n_54)
);

BUFx12_ASAP7_75t_L g30 ( 
.A(n_1),
.Y(n_30)
);

OAI22xp5_ASAP7_75t_SL g31 ( 
.A1(n_2),
.A2(n_29),
.B1(n_30),
.B2(n_32),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_2),
.Y(n_32)
);

AOI22xp33_ASAP7_75t_SL g56 ( 
.A1(n_2),
.A2(n_32),
.B1(n_51),
.B2(n_52),
.Y(n_56)
);

AOI22xp33_ASAP7_75t_SL g93 ( 
.A1(n_2),
.A2(n_32),
.B1(n_61),
.B2(n_62),
.Y(n_93)
);

AOI22xp33_ASAP7_75t_SL g143 ( 
.A1(n_2),
.A2(n_23),
.B1(n_24),
.B2(n_32),
.Y(n_143)
);

BUFx16f_ASAP7_75t_L g65 ( 
.A(n_3),
.Y(n_65)
);

AOI22xp5_ASAP7_75t_SL g169 ( 
.A1(n_4),
.A2(n_61),
.B1(n_62),
.B2(n_170),
.Y(n_169)
);

CKINVDCx20_ASAP7_75t_R g170 ( 
.A(n_4),
.Y(n_170)
);

AOI22xp33_ASAP7_75t_L g180 ( 
.A1(n_4),
.A2(n_51),
.B1(n_52),
.B2(n_170),
.Y(n_180)
);

AOI22xp33_ASAP7_75t_SL g221 ( 
.A1(n_4),
.A2(n_23),
.B1(n_24),
.B2(n_170),
.Y(n_221)
);

AOI22xp33_ASAP7_75t_SL g272 ( 
.A1(n_4),
.A2(n_29),
.B1(n_30),
.B2(n_170),
.Y(n_272)
);

BUFx12f_ASAP7_75t_L g61 ( 
.A(n_5),
.Y(n_61)
);

OAI22xp5_ASAP7_75t_L g59 ( 
.A1(n_6),
.A2(n_60),
.B1(n_61),
.B2(n_62),
.Y(n_59)
);

CKINVDCx20_ASAP7_75t_R g60 ( 
.A(n_6),
.Y(n_60)
);

AOI22xp33_ASAP7_75t_SL g90 ( 
.A1(n_6),
.A2(n_23),
.B1(n_24),
.B2(n_60),
.Y(n_90)
);

AOI22xp33_ASAP7_75t_SL g139 ( 
.A1(n_6),
.A2(n_29),
.B1(n_30),
.B2(n_60),
.Y(n_139)
);

OAI22xp33_ASAP7_75t_SL g262 ( 
.A1(n_6),
.A2(n_51),
.B1(n_52),
.B2(n_60),
.Y(n_262)
);

BUFx12f_ASAP7_75t_L g24 ( 
.A(n_7),
.Y(n_24)
);

INVx4_ASAP7_75t_L g84 ( 
.A(n_8),
.Y(n_84)
);

OAI22xp5_ASAP7_75t_L g35 ( 
.A1(n_9),
.A2(n_29),
.B1(n_30),
.B2(n_36),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_9),
.Y(n_36)
);

AOI22xp33_ASAP7_75t_SL g69 ( 
.A1(n_9),
.A2(n_36),
.B1(n_61),
.B2(n_62),
.Y(n_69)
);

AOI22xp5_ASAP7_75t_L g99 ( 
.A1(n_9),
.A2(n_23),
.B1(n_24),
.B2(n_36),
.Y(n_99)
);

OAI22xp5_ASAP7_75t_L g120 ( 
.A1(n_9),
.A2(n_36),
.B1(n_51),
.B2(n_52),
.Y(n_120)
);

AOI22xp5_ASAP7_75t_SL g87 ( 
.A1(n_10),
.A2(n_23),
.B1(n_24),
.B2(n_88),
.Y(n_87)
);

CKINVDCx14_ASAP7_75t_R g88 ( 
.A(n_10),
.Y(n_88)
);

AOI22xp33_ASAP7_75t_SL g106 ( 
.A1(n_10),
.A2(n_29),
.B1(n_30),
.B2(n_88),
.Y(n_106)
);

OAI22xp5_ASAP7_75t_L g125 ( 
.A1(n_10),
.A2(n_61),
.B1(n_62),
.B2(n_88),
.Y(n_125)
);

AOI22xp5_ASAP7_75t_SL g228 ( 
.A1(n_10),
.A2(n_51),
.B1(n_52),
.B2(n_88),
.Y(n_228)
);

AOI22xp5_ASAP7_75t_L g22 ( 
.A1(n_11),
.A2(n_23),
.B1(n_24),
.B2(n_25),
.Y(n_22)
);

INVx4_ASAP7_75t_L g25 ( 
.A(n_11),
.Y(n_25)
);

OAI22xp5_ASAP7_75t_SL g28 ( 
.A1(n_11),
.A2(n_25),
.B1(n_29),
.B2(n_30),
.Y(n_28)
);

NAND2xp33_ASAP7_75t_SL g258 ( 
.A(n_11),
.B(n_24),
.Y(n_258)
);

AOI22xp33_ASAP7_75t_L g157 ( 
.A1(n_12),
.A2(n_61),
.B1(n_62),
.B2(n_158),
.Y(n_157)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_12),
.Y(n_158)
);

MAJIxp5_ASAP7_75t_L g162 ( 
.A(n_12),
.B(n_52),
.C(n_65),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_L g166 ( 
.A(n_12),
.B(n_86),
.Y(n_166)
);

OAI21xp33_ASAP7_75t_L g190 ( 
.A1(n_12),
.A2(n_121),
.B(n_174),
.Y(n_190)
);

O2A1O1Ixp33_ASAP7_75t_L g200 ( 
.A1(n_12),
.A2(n_23),
.B(n_85),
.C(n_201),
.Y(n_200)
);

AOI22xp33_ASAP7_75t_L g206 ( 
.A1(n_12),
.A2(n_23),
.B1(n_24),
.B2(n_158),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_L g225 ( 
.A(n_12),
.B(n_21),
.Y(n_225)
);

NOR2xp33_ASAP7_75t_L g245 ( 
.A(n_12),
.B(n_29),
.Y(n_245)
);

AOI22xp33_ASAP7_75t_SL g72 ( 
.A1(n_13),
.A2(n_29),
.B1(n_30),
.B2(n_73),
.Y(n_72)
);

CKINVDCx20_ASAP7_75t_R g73 ( 
.A(n_13),
.Y(n_73)
);

AOI22xp33_ASAP7_75t_SL g127 ( 
.A1(n_13),
.A2(n_23),
.B1(n_24),
.B2(n_73),
.Y(n_127)
);

AOI22xp33_ASAP7_75t_SL g203 ( 
.A1(n_13),
.A2(n_51),
.B1(n_52),
.B2(n_73),
.Y(n_203)
);

OAI22xp5_ASAP7_75t_L g251 ( 
.A1(n_13),
.A2(n_61),
.B1(n_62),
.B2(n_73),
.Y(n_251)
);

AOI22xp33_ASAP7_75t_L g76 ( 
.A1(n_14),
.A2(n_29),
.B1(n_30),
.B2(n_77),
.Y(n_76)
);

CKINVDCx20_ASAP7_75t_R g77 ( 
.A(n_14),
.Y(n_77)
);

OAI22xp5_ASAP7_75t_SL g160 ( 
.A1(n_14),
.A2(n_61),
.B1(n_62),
.B2(n_77),
.Y(n_160)
);

OAI22xp5_ASAP7_75t_SL g175 ( 
.A1(n_14),
.A2(n_51),
.B1(n_52),
.B2(n_77),
.Y(n_175)
);

OAI22xp33_ASAP7_75t_SL g208 ( 
.A1(n_14),
.A2(n_23),
.B1(n_24),
.B2(n_77),
.Y(n_208)
);

AOI22xp33_ASAP7_75t_SL g129 ( 
.A1(n_15),
.A2(n_29),
.B1(n_30),
.B2(n_130),
.Y(n_129)
);

CKINVDCx20_ASAP7_75t_R g130 ( 
.A(n_15),
.Y(n_130)
);

AOI22xp5_ASAP7_75t_SL g173 ( 
.A1(n_15),
.A2(n_51),
.B1(n_52),
.B2(n_130),
.Y(n_173)
);

OAI22xp5_ASAP7_75t_L g211 ( 
.A1(n_15),
.A2(n_61),
.B1(n_62),
.B2(n_130),
.Y(n_211)
);

AOI22xp33_ASAP7_75t_SL g248 ( 
.A1(n_15),
.A2(n_23),
.B1(n_24),
.B2(n_130),
.Y(n_248)
);

INVx11_ASAP7_75t_L g53 ( 
.A(n_16),
.Y(n_53)
);

XOR2xp5_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_39),
.Y(n_17)
);

NAND2xp5_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_37),
.Y(n_18)
);

NAND2xp5_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_33),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_20),
.Y(n_38)
);

OAI21xp5_ASAP7_75t_SL g20 ( 
.A1(n_21),
.A2(n_26),
.B(n_31),
.Y(n_20)
);

AOI22xp5_ASAP7_75t_L g34 ( 
.A1(n_21),
.A2(n_26),
.B1(n_31),
.B2(n_35),
.Y(n_34)
);

AOI22xp5_ASAP7_75t_L g322 ( 
.A1(n_21),
.A2(n_26),
.B1(n_35),
.B2(n_323),
.Y(n_322)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_22),
.Y(n_21)
);

NAND2xp5_ASAP7_75t_SL g27 ( 
.A(n_22),
.B(n_28),
.Y(n_27)
);

OAI21xp5_ASAP7_75t_L g71 ( 
.A1(n_22),
.A2(n_72),
.B(n_74),
.Y(n_71)
);

OAI22xp5_ASAP7_75t_L g105 ( 
.A1(n_22),
.A2(n_27),
.B1(n_72),
.B2(n_106),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g132 ( 
.A(n_22),
.B(n_76),
.Y(n_132)
);

OAI22xp5_ASAP7_75t_SL g138 ( 
.A1(n_22),
.A2(n_27),
.B1(n_106),
.B2(n_139),
.Y(n_138)
);

OAI21xp5_ASAP7_75t_L g271 ( 
.A1(n_22),
.A2(n_74),
.B(n_272),
.Y(n_271)
);

OAI22xp5_ASAP7_75t_SL g285 ( 
.A1(n_22),
.A2(n_27),
.B1(n_129),
.B2(n_272),
.Y(n_285)
);

AOI22xp33_ASAP7_75t_L g83 ( 
.A1(n_23),
.A2(n_24),
.B1(n_84),
.B2(n_85),
.Y(n_83)
);

AOI32xp33_ASAP7_75t_L g257 ( 
.A1(n_23),
.A2(n_25),
.A3(n_30),
.B1(n_245),
.B2(n_258),
.Y(n_257)
);

INVx8_ASAP7_75t_L g23 ( 
.A(n_24),
.Y(n_23)
);

NAND2xp5_ASAP7_75t_SL g74 ( 
.A(n_26),
.B(n_75),
.Y(n_74)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_27),
.Y(n_26)
);

OAI21xp5_ASAP7_75t_L g128 ( 
.A1(n_27),
.A2(n_129),
.B(n_131),
.Y(n_128)
);

O2A1O1Ixp33_ASAP7_75t_L g243 ( 
.A1(n_27),
.A2(n_30),
.B(n_158),
.C(n_244),
.Y(n_243)
);

INVx4_ASAP7_75t_L g29 ( 
.A(n_30),
.Y(n_29)
);

NOR2xp33_ASAP7_75t_L g332 ( 
.A(n_33),
.B(n_333),
.Y(n_332)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_34),
.Y(n_33)
);

NAND2xp5_ASAP7_75t_L g37 ( 
.A(n_34),
.B(n_38),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g329 ( 
.A(n_34),
.B(n_330),
.Y(n_329)
);

OAI21xp5_ASAP7_75t_L g39 ( 
.A1(n_40),
.A2(n_329),
.B(n_331),
.Y(n_39)
);

AOI21xp5_ASAP7_75t_L g40 ( 
.A1(n_41),
.A2(n_317),
.B(n_328),
.Y(n_40)
);

AO21x1_ASAP7_75t_L g41 ( 
.A1(n_42),
.A2(n_146),
.B(n_314),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g42 ( 
.A(n_43),
.B(n_133),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g43 ( 
.A(n_44),
.B(n_108),
.Y(n_43)
);

NAND2xp5_ASAP7_75t_L g315 ( 
.A(n_44),
.B(n_108),
.Y(n_315)
);

XOR2xp5_ASAP7_75t_L g44 ( 
.A(n_45),
.B(n_78),
.Y(n_44)
);

MAJIxp5_ASAP7_75t_L g145 ( 
.A(n_45),
.B(n_79),
.C(n_94),
.Y(n_145)
);

OAI21xp5_ASAP7_75t_L g45 ( 
.A1(n_46),
.A2(n_49),
.B(n_71),
.Y(n_45)
);

OAI22xp5_ASAP7_75t_SL g110 ( 
.A1(n_46),
.A2(n_47),
.B1(n_111),
.B2(n_112),
.Y(n_110)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_47),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_L g47 ( 
.A(n_48),
.B(n_57),
.Y(n_47)
);

AOI22xp5_ASAP7_75t_L g112 ( 
.A1(n_48),
.A2(n_49),
.B1(n_71),
.B2(n_113),
.Y(n_112)
);

AOI22xp5_ASAP7_75t_L g301 ( 
.A1(n_48),
.A2(n_49),
.B1(n_57),
.B2(n_58),
.Y(n_301)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_49),
.Y(n_48)
);

OAI21xp5_ASAP7_75t_SL g49 ( 
.A1(n_50),
.A2(n_54),
.B(n_55),
.Y(n_49)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_50),
.Y(n_121)
);

AOI22xp5_ASAP7_75t_SL g178 ( 
.A1(n_50),
.A2(n_54),
.B1(n_179),
.B2(n_181),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_L g188 ( 
.A(n_50),
.B(n_175),
.Y(n_188)
);

AOI22xp5_ASAP7_75t_L g276 ( 
.A1(n_50),
.A2(n_54),
.B1(n_120),
.B2(n_262),
.Y(n_276)
);

NOR2xp33_ASAP7_75t_SL g50 ( 
.A(n_51),
.B(n_54),
.Y(n_50)
);

OA22x2_ASAP7_75t_L g67 ( 
.A1(n_51),
.A2(n_52),
.B1(n_65),
.B2(n_66),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_SL g191 ( 
.A(n_51),
.B(n_192),
.Y(n_191)
);

INVx5_ASAP7_75t_L g51 ( 
.A(n_52),
.Y(n_51)
);

INVx8_ASAP7_75t_L g52 ( 
.A(n_53),
.Y(n_52)
);

CKINVDCx20_ASAP7_75t_R g122 ( 
.A(n_54),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_SL g174 ( 
.A(n_54),
.B(n_175),
.Y(n_174)
);

INVxp67_ASAP7_75t_L g55 ( 
.A(n_56),
.Y(n_55)
);

OAI22xp5_ASAP7_75t_SL g118 ( 
.A1(n_56),
.A2(n_119),
.B1(n_121),
.B2(n_122),
.Y(n_118)
);

CKINVDCx20_ASAP7_75t_R g57 ( 
.A(n_58),
.Y(n_57)
);

AOI22xp5_ASAP7_75t_L g58 ( 
.A1(n_59),
.A2(n_63),
.B1(n_68),
.B2(n_70),
.Y(n_58)
);

AOI22xp5_ASAP7_75t_L g124 ( 
.A1(n_59),
.A2(n_63),
.B1(n_70),
.B2(n_125),
.Y(n_124)
);

INVx6_ASAP7_75t_L g62 ( 
.A(n_61),
.Y(n_62)
);

OAI22xp33_ASAP7_75t_L g64 ( 
.A1(n_61),
.A2(n_62),
.B1(n_65),
.B2(n_66),
.Y(n_64)
);

AO22x1_ASAP7_75t_SL g86 ( 
.A1(n_61),
.A2(n_62),
.B1(n_84),
.B2(n_85),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_SL g161 ( 
.A(n_61),
.B(n_162),
.Y(n_161)
);

OAI21xp33_ASAP7_75t_L g201 ( 
.A1(n_62),
.A2(n_84),
.B(n_158),
.Y(n_201)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_63),
.Y(n_92)
);

OAI21xp5_ASAP7_75t_L g101 ( 
.A1(n_63),
.A2(n_70),
.B(n_102),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_SL g171 ( 
.A(n_63),
.B(n_160),
.Y(n_171)
);

AOI22xp5_ASAP7_75t_L g209 ( 
.A1(n_63),
.A2(n_70),
.B1(n_210),
.B2(n_211),
.Y(n_209)
);

AOI22xp5_ASAP7_75t_L g277 ( 
.A1(n_63),
.A2(n_70),
.B1(n_125),
.B2(n_251),
.Y(n_277)
);

AND2x2_ASAP7_75t_L g63 ( 
.A(n_64),
.B(n_67),
.Y(n_63)
);

INVx6_ASAP7_75t_L g66 ( 
.A(n_65),
.Y(n_66)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_67),
.Y(n_70)
);

OAI22xp5_ASAP7_75t_SL g91 ( 
.A1(n_67),
.A2(n_69),
.B1(n_92),
.B2(n_93),
.Y(n_91)
);

OAI21xp5_ASAP7_75t_L g168 ( 
.A1(n_67),
.A2(n_169),
.B(n_171),
.Y(n_168)
);

NOR2xp33_ASAP7_75t_SL g186 ( 
.A(n_67),
.B(n_158),
.Y(n_186)
);

OAI21xp5_ASAP7_75t_L g249 ( 
.A1(n_67),
.A2(n_171),
.B(n_250),
.Y(n_249)
);

INVxp67_ASAP7_75t_L g68 ( 
.A(n_69),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_L g159 ( 
.A(n_70),
.B(n_160),
.Y(n_159)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_71),
.Y(n_113)
);

INVxp67_ASAP7_75t_L g75 ( 
.A(n_76),
.Y(n_75)
);

XNOR2xp5_ASAP7_75t_L g78 ( 
.A(n_79),
.B(n_94),
.Y(n_78)
);

AOI21xp5_ASAP7_75t_L g114 ( 
.A1(n_79),
.A2(n_80),
.B(n_91),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_80),
.B(n_91),
.Y(n_79)
);

OAI22xp5_ASAP7_75t_SL g80 ( 
.A1(n_81),
.A2(n_87),
.B1(n_89),
.B2(n_90),
.Y(n_80)
);

OAI22xp5_ASAP7_75t_SL g126 ( 
.A1(n_81),
.A2(n_87),
.B1(n_89),
.B2(n_127),
.Y(n_126)
);

OAI22xp5_ASAP7_75t_SL g142 ( 
.A1(n_81),
.A2(n_89),
.B1(n_99),
.B2(n_143),
.Y(n_142)
);

OAI21xp5_ASAP7_75t_SL g205 ( 
.A1(n_81),
.A2(n_206),
.B(n_207),
.Y(n_205)
);

OAI22xp5_ASAP7_75t_SL g247 ( 
.A1(n_81),
.A2(n_89),
.B1(n_221),
.B2(n_248),
.Y(n_247)
);

OAI21xp5_ASAP7_75t_L g270 ( 
.A1(n_81),
.A2(n_207),
.B(n_248),
.Y(n_270)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_82),
.Y(n_81)
);

AOI22xp5_ASAP7_75t_L g96 ( 
.A1(n_82),
.A2(n_86),
.B1(n_97),
.B2(n_98),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g222 ( 
.A(n_82),
.B(n_208),
.Y(n_222)
);

OAI21xp5_ASAP7_75t_SL g320 ( 
.A1(n_82),
.A2(n_86),
.B(n_321),
.Y(n_320)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_83),
.B(n_86),
.Y(n_82)
);

INVx8_ASAP7_75t_L g85 ( 
.A(n_84),
.Y(n_85)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_86),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g207 ( 
.A(n_86),
.B(n_208),
.Y(n_207)
);

OAI21xp5_ASAP7_75t_SL g220 ( 
.A1(n_89),
.A2(n_221),
.B(n_222),
.Y(n_220)
);

OAI21xp5_ASAP7_75t_SL g286 ( 
.A1(n_89),
.A2(n_127),
.B(n_222),
.Y(n_286)
);

INVxp67_ASAP7_75t_L g97 ( 
.A(n_90),
.Y(n_97)
);

OAI21xp33_ASAP7_75t_SL g156 ( 
.A1(n_92),
.A2(n_157),
.B(n_159),
.Y(n_156)
);

OAI21xp5_ASAP7_75t_SL g232 ( 
.A1(n_92),
.A2(n_159),
.B(n_233),
.Y(n_232)
);

INVxp67_ASAP7_75t_L g102 ( 
.A(n_93),
.Y(n_102)
);

AOI22xp5_ASAP7_75t_L g94 ( 
.A1(n_95),
.A2(n_104),
.B1(n_105),
.B2(n_107),
.Y(n_94)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_95),
.Y(n_107)
);

AOI22xp5_ASAP7_75t_L g95 ( 
.A1(n_96),
.A2(n_100),
.B1(n_101),
.B2(n_103),
.Y(n_95)
);

CKINVDCx16_ASAP7_75t_R g103 ( 
.A(n_96),
.Y(n_103)
);

MAJIxp5_ASAP7_75t_SL g144 ( 
.A(n_96),
.B(n_101),
.C(n_105),
.Y(n_144)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_99),
.Y(n_98)
);

AOI22xp5_ASAP7_75t_L g140 ( 
.A1(n_100),
.A2(n_101),
.B1(n_141),
.B2(n_142),
.Y(n_140)
);

CKINVDCx16_ASAP7_75t_R g100 ( 
.A(n_101),
.Y(n_100)
);

MAJIxp5_ASAP7_75t_L g326 ( 
.A(n_101),
.B(n_138),
.C(n_142),
.Y(n_326)
);

AOI22xp5_ASAP7_75t_L g135 ( 
.A1(n_104),
.A2(n_105),
.B1(n_136),
.B2(n_137),
.Y(n_135)
);

CKINVDCx20_ASAP7_75t_R g104 ( 
.A(n_105),
.Y(n_104)
);

MAJIxp5_ASAP7_75t_L g327 ( 
.A(n_105),
.B(n_137),
.C(n_144),
.Y(n_327)
);

MAJIxp5_ASAP7_75t_L g108 ( 
.A(n_109),
.B(n_114),
.C(n_115),
.Y(n_108)
);

AOI22xp5_ASAP7_75t_L g311 ( 
.A1(n_109),
.A2(n_110),
.B1(n_114),
.B2(n_312),
.Y(n_311)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_110),
.Y(n_109)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_112),
.Y(n_111)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_114),
.Y(n_312)
);

XOR2xp5_ASAP7_75t_L g310 ( 
.A(n_115),
.B(n_311),
.Y(n_310)
);

MAJIxp5_ASAP7_75t_L g115 ( 
.A(n_116),
.B(n_126),
.C(n_128),
.Y(n_115)
);

OAI22xp5_ASAP7_75t_SL g303 ( 
.A1(n_116),
.A2(n_117),
.B1(n_304),
.B2(n_305),
.Y(n_303)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_117),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_L g117 ( 
.A(n_118),
.B(n_123),
.Y(n_117)
);

OAI22xp5_ASAP7_75t_SL g281 ( 
.A1(n_118),
.A2(n_123),
.B1(n_124),
.B2(n_282),
.Y(n_281)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_118),
.Y(n_282)
);

CKINVDCx16_ASAP7_75t_R g119 ( 
.A(n_120),
.Y(n_119)
);

OAI21xp5_ASAP7_75t_L g172 ( 
.A1(n_121),
.A2(n_173),
.B(n_174),
.Y(n_172)
);

OAI22xp5_ASAP7_75t_SL g227 ( 
.A1(n_121),
.A2(n_122),
.B1(n_203),
.B2(n_228),
.Y(n_227)
);

OAI22xp5_ASAP7_75t_SL g260 ( 
.A1(n_121),
.A2(n_122),
.B1(n_228),
.B2(n_261),
.Y(n_260)
);

OAI21xp5_ASAP7_75t_SL g187 ( 
.A1(n_122),
.A2(n_180),
.B(n_188),
.Y(n_187)
);

NOR2xp33_ASAP7_75t_L g192 ( 
.A(n_122),
.B(n_158),
.Y(n_192)
);

OAI21xp5_ASAP7_75t_L g202 ( 
.A1(n_122),
.A2(n_188),
.B(n_203),
.Y(n_202)
);

CKINVDCx16_ASAP7_75t_R g123 ( 
.A(n_124),
.Y(n_123)
);

XNOR2xp5_ASAP7_75t_SL g305 ( 
.A(n_126),
.B(n_128),
.Y(n_305)
);

INVxp67_ASAP7_75t_L g131 ( 
.A(n_132),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_SL g242 ( 
.A(n_132),
.B(n_243),
.Y(n_242)
);

OAI21xp33_ASAP7_75t_L g314 ( 
.A1(n_133),
.A2(n_315),
.B(n_316),
.Y(n_314)
);

NOR2xp33_ASAP7_75t_SL g133 ( 
.A(n_134),
.B(n_145),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_L g316 ( 
.A(n_134),
.B(n_145),
.Y(n_316)
);

XNOR2xp5_ASAP7_75t_L g134 ( 
.A(n_135),
.B(n_144),
.Y(n_134)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_137),
.Y(n_136)
);

XNOR2xp5_ASAP7_75t_L g137 ( 
.A(n_138),
.B(n_140),
.Y(n_137)
);

CKINVDCx20_ASAP7_75t_R g323 ( 
.A(n_139),
.Y(n_323)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_142),
.Y(n_141)
);

CKINVDCx16_ASAP7_75t_R g321 ( 
.A(n_143),
.Y(n_321)
);

OAI21xp5_ASAP7_75t_SL g146 ( 
.A1(n_147),
.A2(n_308),
.B(n_313),
.Y(n_146)
);

AOI21xp5_ASAP7_75t_SL g147 ( 
.A1(n_148),
.A2(n_296),
.B(n_307),
.Y(n_147)
);

OAI321xp33_ASAP7_75t_L g148 ( 
.A1(n_149),
.A2(n_264),
.A3(n_289),
.B1(n_294),
.B2(n_295),
.C(n_335),
.Y(n_148)
);

AOI21xp5_ASAP7_75t_SL g149 ( 
.A1(n_150),
.A2(n_237),
.B(n_263),
.Y(n_149)
);

OAI21xp5_ASAP7_75t_L g150 ( 
.A1(n_151),
.A2(n_215),
.B(n_236),
.Y(n_150)
);

AOI21xp5_ASAP7_75t_L g151 ( 
.A1(n_152),
.A2(n_196),
.B(n_214),
.Y(n_151)
);

OAI21xp5_ASAP7_75t_SL g152 ( 
.A1(n_153),
.A2(n_176),
.B(n_195),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_L g153 ( 
.A(n_154),
.B(n_163),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_SL g195 ( 
.A(n_154),
.B(n_163),
.Y(n_195)
);

NOR2xp33_ASAP7_75t_SL g154 ( 
.A(n_155),
.B(n_161),
.Y(n_154)
);

AOI22xp5_ASAP7_75t_SL g182 ( 
.A1(n_155),
.A2(n_156),
.B1(n_161),
.B2(n_183),
.Y(n_182)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_156),
.Y(n_155)
);

CKINVDCx16_ASAP7_75t_R g183 ( 
.A(n_161),
.Y(n_183)
);

XNOR2xp5_ASAP7_75t_L g163 ( 
.A(n_164),
.B(n_172),
.Y(n_163)
);

AOI22xp5_ASAP7_75t_L g164 ( 
.A1(n_165),
.A2(n_166),
.B1(n_167),
.B2(n_168),
.Y(n_164)
);

MAJIxp5_ASAP7_75t_L g197 ( 
.A(n_165),
.B(n_168),
.C(n_172),
.Y(n_197)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_166),
.Y(n_165)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_168),
.Y(n_167)
);

INVxp67_ASAP7_75t_L g210 ( 
.A(n_169),
.Y(n_210)
);

CKINVDCx14_ASAP7_75t_R g181 ( 
.A(n_173),
.Y(n_181)
);

AOI21xp5_ASAP7_75t_L g176 ( 
.A1(n_177),
.A2(n_184),
.B(n_194),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_L g177 ( 
.A(n_178),
.B(n_182),
.Y(n_177)
);

NOR2xp33_ASAP7_75t_SL g194 ( 
.A(n_178),
.B(n_182),
.Y(n_194)
);

INVxp67_ASAP7_75t_L g179 ( 
.A(n_180),
.Y(n_179)
);

OAI21xp5_ASAP7_75t_SL g184 ( 
.A1(n_185),
.A2(n_189),
.B(n_193),
.Y(n_184)
);

NOR2xp33_ASAP7_75t_L g185 ( 
.A(n_186),
.B(n_187),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_SL g193 ( 
.A(n_186),
.B(n_187),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_SL g189 ( 
.A(n_190),
.B(n_191),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_L g196 ( 
.A(n_197),
.B(n_198),
.Y(n_196)
);

NOR2xp33_ASAP7_75t_SL g214 ( 
.A(n_197),
.B(n_198),
.Y(n_214)
);

XNOR2xp5_ASAP7_75t_L g198 ( 
.A(n_199),
.B(n_204),
.Y(n_198)
);

MAJIxp5_ASAP7_75t_L g216 ( 
.A(n_199),
.B(n_209),
.C(n_213),
.Y(n_216)
);

XNOR2xp5_ASAP7_75t_SL g199 ( 
.A(n_200),
.B(n_202),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_L g231 ( 
.A(n_200),
.B(n_202),
.Y(n_231)
);

AOI22xp5_ASAP7_75t_L g204 ( 
.A1(n_205),
.A2(n_209),
.B1(n_212),
.B2(n_213),
.Y(n_204)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_205),
.Y(n_213)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_209),
.Y(n_212)
);

CKINVDCx16_ASAP7_75t_R g233 ( 
.A(n_211),
.Y(n_233)
);

NOR2xp33_ASAP7_75t_L g215 ( 
.A(n_216),
.B(n_217),
.Y(n_215)
);

NAND2xp5_ASAP7_75t_SL g236 ( 
.A(n_216),
.B(n_217),
.Y(n_236)
);

OAI22xp5_ASAP7_75t_SL g217 ( 
.A1(n_218),
.A2(n_219),
.B1(n_229),
.B2(n_230),
.Y(n_217)
);

MAJIxp5_ASAP7_75t_L g238 ( 
.A(n_218),
.B(n_232),
.C(n_234),
.Y(n_238)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_219),
.Y(n_218)
);

XOR2xp5_ASAP7_75t_L g219 ( 
.A(n_220),
.B(n_223),
.Y(n_219)
);

MAJIxp5_ASAP7_75t_L g254 ( 
.A(n_220),
.B(n_224),
.C(n_227),
.Y(n_254)
);

AOI22xp5_ASAP7_75t_L g223 ( 
.A1(n_224),
.A2(n_225),
.B1(n_226),
.B2(n_227),
.Y(n_223)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_225),
.Y(n_224)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_227),
.Y(n_226)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_230),
.Y(n_229)
);

OAI22xp5_ASAP7_75t_SL g230 ( 
.A1(n_231),
.A2(n_232),
.B1(n_234),
.B2(n_235),
.Y(n_230)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_231),
.Y(n_234)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_232),
.Y(n_235)
);

NAND2xp5_ASAP7_75t_L g237 ( 
.A(n_238),
.B(n_239),
.Y(n_237)
);

NOR2xp33_ASAP7_75t_L g263 ( 
.A(n_238),
.B(n_239),
.Y(n_263)
);

XNOR2xp5_ASAP7_75t_L g239 ( 
.A(n_240),
.B(n_253),
.Y(n_239)
);

MAJIxp5_ASAP7_75t_L g290 ( 
.A(n_240),
.B(n_254),
.C(n_255),
.Y(n_290)
);

AOI22xp5_ASAP7_75t_L g240 ( 
.A1(n_241),
.A2(n_242),
.B1(n_246),
.B2(n_252),
.Y(n_240)
);

MAJIxp5_ASAP7_75t_L g278 ( 
.A(n_241),
.B(n_247),
.C(n_249),
.Y(n_278)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_242),
.Y(n_241)
);

INVxp67_ASAP7_75t_L g244 ( 
.A(n_245),
.Y(n_244)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_246),
.Y(n_252)
);

XNOR2xp5_ASAP7_75t_SL g246 ( 
.A(n_247),
.B(n_249),
.Y(n_246)
);

CKINVDCx20_ASAP7_75t_R g250 ( 
.A(n_251),
.Y(n_250)
);

XNOR2xp5_ASAP7_75t_L g253 ( 
.A(n_254),
.B(n_255),
.Y(n_253)
);

AOI22xp5_ASAP7_75t_L g255 ( 
.A1(n_256),
.A2(n_257),
.B1(n_259),
.B2(n_260),
.Y(n_255)
);

NAND2xp5_ASAP7_75t_L g274 ( 
.A(n_256),
.B(n_260),
.Y(n_274)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_257),
.Y(n_256)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_260),
.Y(n_259)
);

INVxp67_ASAP7_75t_L g261 ( 
.A(n_262),
.Y(n_261)
);

NOR2xp33_ASAP7_75t_L g264 ( 
.A(n_265),
.B(n_279),
.Y(n_264)
);

NAND2xp5_ASAP7_75t_L g295 ( 
.A(n_265),
.B(n_279),
.Y(n_295)
);

MAJIxp5_ASAP7_75t_L g265 ( 
.A(n_266),
.B(n_275),
.C(n_278),
.Y(n_265)
);

OAI22xp5_ASAP7_75t_SL g291 ( 
.A1(n_266),
.A2(n_267),
.B1(n_292),
.B2(n_293),
.Y(n_291)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_267),
.Y(n_266)
);

XOR2xp5_ASAP7_75t_L g267 ( 
.A(n_268),
.B(n_274),
.Y(n_267)
);

AOI22xp5_ASAP7_75t_L g268 ( 
.A1(n_269),
.A2(n_270),
.B1(n_271),
.B2(n_273),
.Y(n_268)
);

MAJIxp5_ASAP7_75t_L g288 ( 
.A(n_269),
.B(n_273),
.C(n_274),
.Y(n_288)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_270),
.Y(n_269)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_271),
.Y(n_273)
);

XNOR2xp5_ASAP7_75t_SL g293 ( 
.A(n_275),
.B(n_278),
.Y(n_293)
);

XNOR2xp5_ASAP7_75t_L g275 ( 
.A(n_276),
.B(n_277),
.Y(n_275)
);

NOR2xp33_ASAP7_75t_L g287 ( 
.A(n_276),
.B(n_277),
.Y(n_287)
);

XNOR2xp5_ASAP7_75t_L g279 ( 
.A(n_280),
.B(n_288),
.Y(n_279)
);

XNOR2xp5_ASAP7_75t_L g280 ( 
.A(n_281),
.B(n_283),
.Y(n_280)
);

MAJIxp5_ASAP7_75t_L g306 ( 
.A(n_281),
.B(n_283),
.C(n_288),
.Y(n_306)
);

XNOR2xp5_ASAP7_75t_SL g283 ( 
.A(n_284),
.B(n_287),
.Y(n_283)
);

XNOR2xp5_ASAP7_75t_L g284 ( 
.A(n_285),
.B(n_286),
.Y(n_284)
);

MAJIxp5_ASAP7_75t_L g298 ( 
.A(n_285),
.B(n_286),
.C(n_287),
.Y(n_298)
);

NOR2xp33_ASAP7_75t_L g289 ( 
.A(n_290),
.B(n_291),
.Y(n_289)
);

NAND2xp5_ASAP7_75t_SL g294 ( 
.A(n_290),
.B(n_291),
.Y(n_294)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_293),
.Y(n_292)
);

NAND2xp5_ASAP7_75t_SL g296 ( 
.A(n_297),
.B(n_306),
.Y(n_296)
);

NOR2xp33_ASAP7_75t_L g307 ( 
.A(n_297),
.B(n_306),
.Y(n_307)
);

XNOR2xp5_ASAP7_75t_L g297 ( 
.A(n_298),
.B(n_299),
.Y(n_297)
);

MAJIxp5_ASAP7_75t_L g309 ( 
.A(n_298),
.B(n_301),
.C(n_302),
.Y(n_309)
);

AOI22xp5_ASAP7_75t_L g299 ( 
.A1(n_300),
.A2(n_301),
.B1(n_302),
.B2(n_303),
.Y(n_299)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_301),
.Y(n_300)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_303),
.Y(n_302)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_305),
.Y(n_304)
);

NOR2xp33_ASAP7_75t_L g308 ( 
.A(n_309),
.B(n_310),
.Y(n_308)
);

NAND2xp5_ASAP7_75t_L g313 ( 
.A(n_309),
.B(n_310),
.Y(n_313)
);

NAND2xp5_ASAP7_75t_L g317 ( 
.A(n_318),
.B(n_327),
.Y(n_317)
);

NOR2xp33_ASAP7_75t_L g328 ( 
.A(n_318),
.B(n_327),
.Y(n_328)
);

XNOR2xp5_ASAP7_75t_L g318 ( 
.A(n_319),
.B(n_326),
.Y(n_318)
);

AOI22xp5_ASAP7_75t_L g319 ( 
.A1(n_320),
.A2(n_322),
.B1(n_324),
.B2(n_325),
.Y(n_319)
);

CKINVDCx20_ASAP7_75t_R g324 ( 
.A(n_320),
.Y(n_324)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_322),
.Y(n_325)
);

MAJIxp5_ASAP7_75t_L g330 ( 
.A(n_322),
.B(n_324),
.C(n_326),
.Y(n_330)
);

CKINVDCx16_ASAP7_75t_R g333 ( 
.A(n_330),
.Y(n_333)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_332),
.Y(n_331)
);


endmodule