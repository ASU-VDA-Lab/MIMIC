module real_jpeg_16201_n_18 (n_17, n_8, n_0, n_2, n_10, n_9, n_12, n_584, n_6, n_11, n_14, n_7, n_3, n_5, n_4, n_1, n_16, n_15, n_13, n_18);

input n_17;
input n_8;
input n_0;
input n_2;
input n_10;
input n_9;
input n_12;
input n_584;
input n_6;
input n_11;
input n_14;
input n_7;
input n_3;
input n_5;
input n_4;
input n_1;
input n_16;
input n_15;
input n_13;

output n_18;

wire n_384;
wire n_37;
wire n_430;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_460;
wire n_300;
wire n_415;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_518;
wire n_446;
wire n_199;
wire n_535;
wire n_95;
wire n_541;
wire n_441;
wire n_557;
wire n_238;
wire n_67;
wire n_350;
wire n_235;
wire n_107;
wire n_369;
wire n_498;
wire n_471;
wire n_376;
wire n_354;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_553;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_574;
wire n_490;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_355;
wire n_123;
wire n_463;
wire n_425;
wire n_455;
wire n_462;
wire n_50;
wire n_409;
wire n_485;
wire n_186;
wire n_137;
wire n_491;
wire n_72;
wire n_440;
wire n_171;
wire n_151;
wire n_272;
wire n_461;
wire n_198;
wire n_203;
wire n_500;
wire n_562;
wire n_23;
wire n_362;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_339;
wire n_326;
wire n_80;
wire n_30;
wire n_328;
wire n_149;
wire n_366;
wire n_332;
wire n_578;
wire n_456;
wire n_259;
wire n_556;
wire n_57;
wire n_507;
wire n_157;
wire n_84;
wire n_560;
wire n_538;
wire n_527;
wire n_55;
wire n_499;
wire n_58;
wire n_52;
wire n_565;
wire n_466;
wire n_353;
wire n_453;
wire n_551;
wire n_230;
wire n_417;
wire n_428;
wire n_128;
wire n_202;
wire n_216;
wire n_483;
wire n_367;
wire n_127;
wire n_356;
wire n_365;
wire n_423;
wire n_464;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_422;
wire n_317;
wire n_506;
wire n_108;
wire n_550;
wire n_233;
wire n_73;
wire n_532;
wire n_516;
wire n_348;
wire n_473;
wire n_252;
wire n_363;
wire n_310;
wire n_345;
wire n_525;
wire n_78;
wire n_83;
wire n_288;
wire n_221;
wire n_393;
wire n_489;
wire n_104;
wire n_153;
wire n_443;
wire n_337;
wire n_544;
wire n_131;
wire n_439;
wire n_517;
wire n_322;
wire n_87;
wire n_40;
wire n_561;
wire n_98;
wire n_469;
wire n_378;
wire n_200;
wire n_432;
wire n_465;
wire n_569;
wire n_335;
wire n_214;
wire n_113;
wire n_566;
wire n_543;
wire n_251;
wire n_459;
wire n_576;
wire n_139;
wire n_33;
wire n_338;
wire n_175;
wire n_488;
wire n_156;
wire n_387;
wire n_434;
wire n_66;
wire n_577;
wire n_305;
wire n_505;
wire n_62;
wire n_254;
wire n_250;
wire n_564;
wire n_304;
wire n_390;
wire n_77;
wire n_399;
wire n_470;
wire n_219;
wire n_372;
wire n_122;
wire n_19;
wire n_262;
wire n_334;
wire n_383;
wire n_246;
wire n_523;
wire n_21;
wire n_476;
wire n_529;
wire n_69;
wire n_31;
wire n_426;
wire n_154;
wire n_495;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_371;
wire n_410;
wire n_421;
wire n_110;
wire n_195;
wire n_533;
wire n_289;
wire n_117;
wire n_193;
wire n_382;
wire n_411;
wire n_20;
wire n_278;
wire n_314;
wire n_103;
wire n_559;
wire n_232;
wire n_582;
wire n_448;
wire n_212;
wire n_284;
wire n_579;
wire n_402;
wire n_478;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_452;
wire n_213;
wire n_511;
wire n_524;
wire n_25;
wire n_542;
wire n_480;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_515;
wire n_89;
wire n_407;
wire n_419;
wire n_386;
wire n_521;
wire n_341;
wire n_331;
wire n_49;
wire n_514;
wire n_68;
wire n_497;
wire n_395;
wire n_146;
wire n_496;
wire n_323;
wire n_215;
wire n_176;
wire n_166;
wire n_286;
wire n_312;
wire n_325;
wire n_307;
wire n_316;
wire n_161;
wire n_207;
wire n_526;
wire n_431;
wire n_420;
wire n_357;
wire n_237;
wire n_445;
wire n_173;
wire n_115;
wire n_474;
wire n_184;
wire n_164;
wire n_380;
wire n_414;
wire n_140;
wire n_126;
wire n_342;
wire n_120;
wire n_155;
wire n_572;
wire n_405;
wire n_412;
wire n_548;
wire n_319;
wire n_93;
wire n_487;
wire n_242;
wire n_493;
wire n_142;
wire n_522;
wire n_397;
wire n_76;
wire n_403;
wire n_79;
wire n_282;
wire n_147;
wire n_359;
wire n_265;
wire n_231;
wire n_44;
wire n_482;
wire n_208;
wire n_162;
wire n_449;
wire n_106;
wire n_172;
wire n_531;
wire n_285;
wire n_546;
wire n_112;
wire n_554;
wire n_508;
wire n_145;
wire n_266;
wire n_377;
wire n_109;
wire n_503;
wire n_391;
wire n_427;
wire n_401;
wire n_536;
wire n_148;
wire n_373;
wire n_563;
wire n_558;
wire n_510;
wire n_396;
wire n_501;
wire n_392;
wire n_575;
wire n_375;
wire n_196;
wire n_298;
wire n_330;
wire n_333;
wire n_450;
wire n_492;
wire n_152;
wire n_270;
wire n_159;
wire n_429;
wire n_347;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_537;
wire n_90;
wire n_336;
wire n_258;
wire n_458;
wire n_150;
wire n_41;
wire n_74;
wire n_475;
wire n_404;
wire n_158;
wire n_204;
wire n_241;
wire n_504;
wire n_111;
wire n_479;
wire n_226;
wire n_125;
wire n_297;
wire n_413;
wire n_494;
wire n_539;
wire n_512;
wire n_75;
wire n_581;
wire n_346;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_457;
wire n_119;
wire n_283;
wire n_181;
wire n_358;
wire n_534;
wire n_256;
wire n_520;
wire n_273;
wire n_253;
wire n_54;
wire n_168;
wire n_38;
wire n_442;
wire n_385;
wire n_201;
wire n_545;
wire n_484;
wire n_260;
wire n_247;
wire n_249;
wire n_349;
wire n_418;
wire n_502;
wire n_472;
wire n_292;
wire n_343;
wire n_486;
wire n_64;
wire n_291;
wire n_236;
wire n_370;
wire n_276;
wire n_374;
wire n_287;
wire n_388;
wire n_174;
wire n_400;
wire n_255;
wire n_299;
wire n_243;
wire n_352;
wire n_477;
wire n_56;
wire n_293;
wire n_275;
wire n_381;
wire n_227;
wire n_229;
wire n_454;
wire n_571;
wire n_573;
wire n_379;
wire n_141;
wire n_555;
wire n_65;
wire n_188;
wire n_178;
wire n_444;
wire n_360;
wire n_398;
wire n_189;
wire n_170;
wire n_570;
wire n_28;
wire n_245;
wire n_451;
wire n_45;
wire n_437;
wire n_268;
wire n_42;
wire n_313;
wire n_94;
wire n_547;
wire n_309;
wire n_294;
wire n_116;
wire n_416;
wire n_513;
wire n_143;
wire n_351;
wire n_467;
wire n_129;
wire n_135;
wire n_306;
wire n_540;
wire n_218;
wire n_528;
wire n_165;
wire n_406;
wire n_303;
wire n_321;
wire n_100;
wire n_368;
wire n_567;
wire n_51;
wire n_509;
wire n_205;
wire n_519;
wire n_530;
wire n_361;
wire n_324;
wire n_86;
wire n_261;
wire n_549;
wire n_70;
wire n_568;
wire n_435;
wire n_32;
wire n_228;
wire n_389;
wire n_580;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_438;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_481;
wire n_191;
wire n_394;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_436;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_424;
wire n_468;
wire n_133;
wire n_257;
wire n_447;
wire n_344;
wire n_210;
wire n_206;
wire n_552;
wire n_408;
wire n_85;
wire n_96;
wire n_308;
wire n_433;
wire n_364;

INVx1_ASAP7_75t_L g165 ( 
.A(n_0),
.Y(n_165)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_0),
.Y(n_174)
);

BUFx6f_ASAP7_75t_L g181 ( 
.A(n_0),
.Y(n_181)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_1),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_1),
.Y(n_37)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_1),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_1),
.Y(n_50)
);

INVx1_ASAP7_75t_L g415 ( 
.A(n_1),
.Y(n_415)
);

AOI22xp5_ASAP7_75t_L g244 ( 
.A1(n_2),
.A2(n_245),
.B1(n_248),
.B2(n_249),
.Y(n_244)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_2),
.Y(n_248)
);

OAI22xp5_ASAP7_75t_SL g350 ( 
.A1(n_2),
.A2(n_248),
.B1(n_351),
.B2(n_353),
.Y(n_350)
);

OAI22xp5_ASAP7_75t_SL g459 ( 
.A1(n_2),
.A2(n_248),
.B1(n_460),
.B2(n_463),
.Y(n_459)
);

AOI22xp33_ASAP7_75t_SL g469 ( 
.A1(n_2),
.A2(n_248),
.B1(n_266),
.B2(n_470),
.Y(n_469)
);

AOI22xp33_ASAP7_75t_L g97 ( 
.A1(n_3),
.A2(n_98),
.B1(n_103),
.B2(n_109),
.Y(n_97)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_3),
.Y(n_109)
);

OAI22xp5_ASAP7_75t_SL g217 ( 
.A1(n_3),
.A2(n_56),
.B1(n_109),
.B2(n_218),
.Y(n_217)
);

AOI22xp33_ASAP7_75t_SL g52 ( 
.A1(n_4),
.A2(n_53),
.B1(n_56),
.B2(n_60),
.Y(n_52)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_4),
.Y(n_60)
);

AOI22xp33_ASAP7_75t_SL g189 ( 
.A1(n_4),
.A2(n_60),
.B1(n_190),
.B2(n_191),
.Y(n_189)
);

OAI22xp33_ASAP7_75t_SL g323 ( 
.A1(n_4),
.A2(n_60),
.B1(n_91),
.B2(n_324),
.Y(n_323)
);

AOI22xp33_ASAP7_75t_SL g570 ( 
.A1(n_4),
.A2(n_60),
.B1(n_571),
.B2(n_572),
.Y(n_570)
);

INVx2_ASAP7_75t_L g80 ( 
.A(n_5),
.Y(n_80)
);

BUFx3_ASAP7_75t_L g334 ( 
.A(n_5),
.Y(n_334)
);

BUFx5_ASAP7_75t_L g394 ( 
.A(n_5),
.Y(n_394)
);

BUFx5_ASAP7_75t_L g486 ( 
.A(n_5),
.Y(n_486)
);

INVxp67_ASAP7_75t_L g310 ( 
.A(n_6),
.Y(n_310)
);

NAND2xp5_ASAP7_75t_L g395 ( 
.A(n_6),
.B(n_150),
.Y(n_395)
);

NAND2xp5_ASAP7_75t_L g456 ( 
.A(n_6),
.B(n_188),
.Y(n_456)
);

OAI22xp5_ASAP7_75t_SL g487 ( 
.A1(n_6),
.A2(n_77),
.B1(n_482),
.B2(n_488),
.Y(n_487)
);

OAI32xp33_ASAP7_75t_L g510 ( 
.A1(n_6),
.A2(n_170),
.A3(n_511),
.B1(n_513),
.B2(n_516),
.Y(n_510)
);

AOI22xp33_ASAP7_75t_SL g524 ( 
.A1(n_6),
.A2(n_310),
.B1(n_525),
.B2(n_526),
.Y(n_524)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_7),
.Y(n_33)
);

INVx2_ASAP7_75t_L g55 ( 
.A(n_7),
.Y(n_55)
);

BUFx3_ASAP7_75t_L g59 ( 
.A(n_7),
.Y(n_59)
);

INVx3_ASAP7_75t_L g74 ( 
.A(n_7),
.Y(n_74)
);

BUFx6f_ASAP7_75t_L g183 ( 
.A(n_7),
.Y(n_183)
);

BUFx3_ASAP7_75t_L g214 ( 
.A(n_7),
.Y(n_214)
);

BUFx5_ASAP7_75t_L g430 ( 
.A(n_7),
.Y(n_430)
);

AOI22xp33_ASAP7_75t_L g85 ( 
.A1(n_8),
.A2(n_86),
.B1(n_90),
.B2(n_91),
.Y(n_85)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_8),
.Y(n_90)
);

AOI22xp33_ASAP7_75t_SL g209 ( 
.A1(n_8),
.A2(n_90),
.B1(n_210),
.B2(n_215),
.Y(n_209)
);

AOI22xp5_ASAP7_75t_L g575 ( 
.A1(n_8),
.A2(n_90),
.B1(n_201),
.B2(n_576),
.Y(n_575)
);

AOI22xp5_ASAP7_75t_SL g152 ( 
.A1(n_9),
.A2(n_153),
.B1(n_155),
.B2(n_159),
.Y(n_152)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_9),
.Y(n_159)
);

AOI22xp5_ASAP7_75t_SL g227 ( 
.A1(n_9),
.A2(n_143),
.B1(n_159),
.B2(n_228),
.Y(n_227)
);

AOI22xp33_ASAP7_75t_L g256 ( 
.A1(n_9),
.A2(n_159),
.B1(n_257),
.B2(n_259),
.Y(n_256)
);

OAI22xp5_ASAP7_75t_SL g383 ( 
.A1(n_9),
.A2(n_159),
.B1(n_384),
.B2(n_388),
.Y(n_383)
);

OAI22xp5_ASAP7_75t_L g336 ( 
.A1(n_10),
.A2(n_139),
.B1(n_143),
.B2(n_337),
.Y(n_336)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_10),
.Y(n_337)
);

AOI22xp5_ASAP7_75t_L g375 ( 
.A1(n_10),
.A2(n_337),
.B1(n_376),
.B2(n_380),
.Y(n_375)
);

OAI22xp5_ASAP7_75t_SL g426 ( 
.A1(n_10),
.A2(n_337),
.B1(n_427),
.B2(n_431),
.Y(n_426)
);

AOI22xp5_ASAP7_75t_SL g488 ( 
.A1(n_10),
.A2(n_337),
.B1(n_489),
.B2(n_495),
.Y(n_488)
);

INVx6_ASAP7_75t_L g116 ( 
.A(n_11),
.Y(n_116)
);

BUFx6f_ASAP7_75t_L g122 ( 
.A(n_11),
.Y(n_122)
);

BUFx6f_ASAP7_75t_L g126 ( 
.A(n_11),
.Y(n_126)
);

BUFx6f_ASAP7_75t_L g130 ( 
.A(n_12),
.Y(n_130)
);

BUFx6f_ASAP7_75t_L g158 ( 
.A(n_12),
.Y(n_158)
);

AOI22xp5_ASAP7_75t_L g133 ( 
.A1(n_13),
.A2(n_134),
.B1(n_138),
.B2(n_139),
.Y(n_133)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_13),
.Y(n_138)
);

OAI22xp5_ASAP7_75t_L g298 ( 
.A1(n_13),
.A2(n_138),
.B1(n_299),
.B2(n_304),
.Y(n_298)
);

AOI22xp5_ASAP7_75t_L g435 ( 
.A1(n_13),
.A2(n_138),
.B1(n_436),
.B2(n_440),
.Y(n_435)
);

OAI22xp5_ASAP7_75t_L g530 ( 
.A1(n_13),
.A2(n_53),
.B1(n_138),
.B2(n_531),
.Y(n_530)
);

BUFx12f_ASAP7_75t_L g44 ( 
.A(n_14),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_14),
.Y(n_47)
);

BUFx4f_ASAP7_75t_L g89 ( 
.A(n_14),
.Y(n_89)
);

INVx2_ASAP7_75t_L g108 ( 
.A(n_14),
.Y(n_108)
);

AOI22xp33_ASAP7_75t_L g65 ( 
.A1(n_15),
.A2(n_66),
.B1(n_69),
.B2(n_70),
.Y(n_65)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_15),
.Y(n_69)
);

AOI22xp5_ASAP7_75t_L g200 ( 
.A1(n_15),
.A2(n_69),
.B1(n_201),
.B2(n_205),
.Y(n_200)
);

AOI22xp5_ASAP7_75t_SL g262 ( 
.A1(n_15),
.A2(n_69),
.B1(n_263),
.B2(n_267),
.Y(n_262)
);

AOI22xp5_ASAP7_75t_L g142 ( 
.A1(n_16),
.A2(n_143),
.B1(n_145),
.B2(n_146),
.Y(n_142)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_16),
.Y(n_145)
);

AOI22xp5_ASAP7_75t_L g276 ( 
.A1(n_16),
.A2(n_145),
.B1(n_277),
.B2(n_282),
.Y(n_276)
);

OAI22xp5_ASAP7_75t_L g359 ( 
.A1(n_16),
.A2(n_145),
.B1(n_360),
.B2(n_361),
.Y(n_359)
);

OAI22xp5_ASAP7_75t_SL g448 ( 
.A1(n_16),
.A2(n_145),
.B1(n_449),
.B2(n_451),
.Y(n_448)
);

BUFx3_ASAP7_75t_L g118 ( 
.A(n_17),
.Y(n_118)
);

INVx2_ASAP7_75t_L g137 ( 
.A(n_17),
.Y(n_137)
);

BUFx8_ASAP7_75t_L g141 ( 
.A(n_17),
.Y(n_141)
);

BUFx5_ASAP7_75t_L g229 ( 
.A(n_17),
.Y(n_229)
);

XOR2xp5_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_559),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_20),
.Y(n_19)
);

INVxp67_ASAP7_75t_SL g20 ( 
.A(n_21),
.Y(n_20)
);

OAI21xp5_ASAP7_75t_L g21 ( 
.A1(n_22),
.A2(n_399),
.B(n_554),
.Y(n_21)
);

NAND3xp33_ASAP7_75t_L g22 ( 
.A(n_23),
.B(n_285),
.C(n_339),
.Y(n_22)
);

A2O1A1O1Ixp25_ASAP7_75t_L g554 ( 
.A1(n_23),
.A2(n_285),
.B(n_555),
.C(n_557),
.D(n_558),
.Y(n_554)
);

NAND2xp5_ASAP7_75t_SL g23 ( 
.A(n_24),
.B(n_235),
.Y(n_23)
);

NOR2xp33_ASAP7_75t_L g558 ( 
.A(n_24),
.B(n_235),
.Y(n_558)
);

XNOR2xp5_ASAP7_75t_L g24 ( 
.A(n_25),
.B(n_194),
.Y(n_24)
);

MAJIxp5_ASAP7_75t_L g561 ( 
.A(n_25),
.B(n_562),
.C(n_563),
.Y(n_561)
);

MAJIxp5_ASAP7_75t_L g25 ( 
.A(n_26),
.B(n_110),
.C(n_151),
.Y(n_25)
);

XNOR2xp5_ASAP7_75t_L g237 ( 
.A(n_26),
.B(n_238),
.Y(n_237)
);

AOI21xp5_ASAP7_75t_L g26 ( 
.A1(n_27),
.A2(n_61),
.B(n_75),
.Y(n_26)
);

NAND2xp5_ASAP7_75t_L g293 ( 
.A(n_27),
.B(n_61),
.Y(n_293)
);

NAND2xp5_ASAP7_75t_SL g27 ( 
.A(n_28),
.B(n_51),
.Y(n_27)
);

AOI22xp5_ASAP7_75t_SL g207 ( 
.A1(n_28),
.A2(n_62),
.B1(n_208),
.B2(n_217),
.Y(n_207)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_28),
.Y(n_233)
);

AOI22xp5_ASAP7_75t_L g358 ( 
.A1(n_28),
.A2(n_62),
.B1(n_359),
.B2(n_366),
.Y(n_358)
);

AOI22xp5_ASAP7_75t_L g421 ( 
.A1(n_28),
.A2(n_62),
.B1(n_422),
.B2(n_426),
.Y(n_421)
);

AOI22xp5_ASAP7_75t_SL g458 ( 
.A1(n_28),
.A2(n_62),
.B1(n_426),
.B2(n_459),
.Y(n_458)
);

AOI22xp5_ASAP7_75t_L g529 ( 
.A1(n_28),
.A2(n_62),
.B1(n_459),
.B2(n_530),
.Y(n_529)
);

OA21x2_ASAP7_75t_L g578 ( 
.A1(n_28),
.A2(n_62),
.B(n_217),
.Y(n_578)
);

AND2x2_ASAP7_75t_L g28 ( 
.A(n_29),
.B(n_39),
.Y(n_28)
);

OAI22xp33_ASAP7_75t_L g29 ( 
.A1(n_30),
.A2(n_34),
.B1(n_36),
.B2(n_38),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_31),
.Y(n_30)
);

INVx2_ASAP7_75t_L g31 ( 
.A(n_32),
.Y(n_31)
);

INVx2_ASAP7_75t_L g38 ( 
.A(n_32),
.Y(n_38)
);

INVx1_ASAP7_75t_L g409 ( 
.A(n_32),
.Y(n_409)
);

INVx6_ASAP7_75t_L g32 ( 
.A(n_33),
.Y(n_32)
);

INVx2_ASAP7_75t_L g178 ( 
.A(n_33),
.Y(n_178)
);

BUFx6f_ASAP7_75t_L g462 ( 
.A(n_33),
.Y(n_462)
);

BUFx3_ASAP7_75t_L g34 ( 
.A(n_35),
.Y(n_34)
);

INVx6_ASAP7_75t_L g36 ( 
.A(n_37),
.Y(n_36)
);

BUFx3_ASAP7_75t_L g63 ( 
.A(n_39),
.Y(n_63)
);

AOI22xp5_ASAP7_75t_L g39 ( 
.A1(n_40),
.A2(n_43),
.B1(n_45),
.B2(n_48),
.Y(n_39)
);

INVx4_ASAP7_75t_L g40 ( 
.A(n_41),
.Y(n_40)
);

BUFx3_ASAP7_75t_L g41 ( 
.A(n_42),
.Y(n_41)
);

INVx4_ASAP7_75t_L g43 ( 
.A(n_44),
.Y(n_43)
);

INVx5_ASAP7_75t_L g387 ( 
.A(n_44),
.Y(n_387)
);

BUFx6f_ASAP7_75t_L g419 ( 
.A(n_44),
.Y(n_419)
);

INVx2_ASAP7_75t_L g494 ( 
.A(n_44),
.Y(n_494)
);

INVx2_ASAP7_75t_L g45 ( 
.A(n_46),
.Y(n_45)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_47),
.Y(n_46)
);

INVx2_ASAP7_75t_L g83 ( 
.A(n_47),
.Y(n_83)
);

INVx3_ASAP7_75t_L g102 ( 
.A(n_47),
.Y(n_102)
);

INVx3_ASAP7_75t_L g48 ( 
.A(n_49),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_50),
.Y(n_49)
);

INVxp67_ASAP7_75t_L g51 ( 
.A(n_52),
.Y(n_51)
);

OAI22xp5_ASAP7_75t_SL g255 ( 
.A1(n_52),
.A2(n_63),
.B1(n_233),
.B2(n_256),
.Y(n_255)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_54),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_55),
.Y(n_54)
);

INVx2_ASAP7_75t_L g68 ( 
.A(n_55),
.Y(n_68)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_57),
.Y(n_56)
);

BUFx2_ASAP7_75t_L g57 ( 
.A(n_58),
.Y(n_57)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_59),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_SL g61 ( 
.A(n_62),
.B(n_64),
.Y(n_61)
);

INVx2_ASAP7_75t_SL g62 ( 
.A(n_63),
.Y(n_62)
);

OAI22xp5_ASAP7_75t_SL g232 ( 
.A1(n_63),
.A2(n_65),
.B1(n_209),
.B2(n_233),
.Y(n_232)
);

NOR2xp33_ASAP7_75t_L g502 ( 
.A(n_63),
.B(n_310),
.Y(n_502)
);

OAI22xp5_ASAP7_75t_SL g541 ( 
.A1(n_63),
.A2(n_233),
.B1(n_542),
.B2(n_543),
.Y(n_541)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_65),
.Y(n_64)
);

INVx4_ASAP7_75t_L g66 ( 
.A(n_67),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_68),
.Y(n_67)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_71),
.Y(n_70)
);

INVx2_ASAP7_75t_L g71 ( 
.A(n_72),
.Y(n_71)
);

INVx3_ASAP7_75t_L g72 ( 
.A(n_73),
.Y(n_72)
);

BUFx3_ASAP7_75t_L g73 ( 
.A(n_74),
.Y(n_73)
);

INVx2_ASAP7_75t_L g260 ( 
.A(n_74),
.Y(n_260)
);

INVx2_ASAP7_75t_L g365 ( 
.A(n_74),
.Y(n_365)
);

BUFx3_ASAP7_75t_L g425 ( 
.A(n_74),
.Y(n_425)
);

XNOR2xp5_ASAP7_75t_L g292 ( 
.A(n_75),
.B(n_293),
.Y(n_292)
);

AOI22xp5_ASAP7_75t_L g75 ( 
.A1(n_76),
.A2(n_84),
.B1(n_94),
.B2(n_96),
.Y(n_75)
);

AOI22x1_ASAP7_75t_SL g382 ( 
.A1(n_76),
.A2(n_323),
.B1(n_383),
.B2(n_392),
.Y(n_382)
);

AOI22xp5_ASAP7_75t_L g467 ( 
.A1(n_76),
.A2(n_468),
.B1(n_471),
.B2(n_473),
.Y(n_467)
);

AOI22xp5_ASAP7_75t_L g518 ( 
.A1(n_76),
.A2(n_273),
.B1(n_383),
.B2(n_448),
.Y(n_518)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_77),
.Y(n_76)
);

AO21x2_ASAP7_75t_L g224 ( 
.A1(n_77),
.A2(n_97),
.B(n_225),
.Y(n_224)
);

OAI22xp5_ASAP7_75t_SL g261 ( 
.A1(n_77),
.A2(n_85),
.B1(n_262),
.B2(n_272),
.Y(n_261)
);

OAI22xp5_ASAP7_75t_L g321 ( 
.A1(n_77),
.A2(n_262),
.B1(n_322),
.B2(n_328),
.Y(n_321)
);

OAI22xp5_ASAP7_75t_L g434 ( 
.A1(n_77),
.A2(n_435),
.B1(n_443),
.B2(n_447),
.Y(n_434)
);

OAI22xp5_ASAP7_75t_SL g499 ( 
.A1(n_77),
.A2(n_469),
.B1(n_488),
.B2(n_500),
.Y(n_499)
);

OR2x2_ASAP7_75t_L g77 ( 
.A(n_78),
.B(n_81),
.Y(n_77)
);

BUFx6f_ASAP7_75t_L g95 ( 
.A(n_78),
.Y(n_95)
);

BUFx6f_ASAP7_75t_L g78 ( 
.A(n_79),
.Y(n_78)
);

INVx1_ASAP7_75t_L g446 ( 
.A(n_79),
.Y(n_446)
);

INVx2_ASAP7_75t_L g79 ( 
.A(n_80),
.Y(n_79)
);

INVx3_ASAP7_75t_L g274 ( 
.A(n_80),
.Y(n_274)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_82),
.Y(n_81)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_83),
.Y(n_82)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_85),
.Y(n_84)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_87),
.Y(n_86)
);

INVx2_ASAP7_75t_L g87 ( 
.A(n_88),
.Y(n_87)
);

BUFx6f_ASAP7_75t_L g411 ( 
.A(n_88),
.Y(n_411)
);

INVx2_ASAP7_75t_L g88 ( 
.A(n_89),
.Y(n_88)
);

INVx2_ASAP7_75t_L g93 ( 
.A(n_89),
.Y(n_93)
);

INVx2_ASAP7_75t_L g439 ( 
.A(n_89),
.Y(n_439)
);

HB1xp67_ASAP7_75t_L g91 ( 
.A(n_92),
.Y(n_91)
);

INVx2_ASAP7_75t_L g92 ( 
.A(n_93),
.Y(n_92)
);

BUFx3_ASAP7_75t_L g94 ( 
.A(n_95),
.Y(n_94)
);

INVx2_ASAP7_75t_L g225 ( 
.A(n_95),
.Y(n_225)
);

INVxp67_ASAP7_75t_L g96 ( 
.A(n_97),
.Y(n_96)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_99),
.Y(n_98)
);

INVx3_ASAP7_75t_L g99 ( 
.A(n_100),
.Y(n_99)
);

INVx2_ASAP7_75t_L g100 ( 
.A(n_101),
.Y(n_100)
);

INVx2_ASAP7_75t_L g101 ( 
.A(n_102),
.Y(n_101)
);

INVx2_ASAP7_75t_L g391 ( 
.A(n_102),
.Y(n_391)
);

INVx2_ASAP7_75t_L g454 ( 
.A(n_102),
.Y(n_454)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_104),
.Y(n_103)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_105),
.Y(n_104)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_106),
.Y(n_105)
);

BUFx6f_ASAP7_75t_L g106 ( 
.A(n_107),
.Y(n_106)
);

INVx2_ASAP7_75t_L g266 ( 
.A(n_107),
.Y(n_266)
);

INVx3_ASAP7_75t_L g271 ( 
.A(n_107),
.Y(n_271)
);

BUFx6f_ASAP7_75t_L g107 ( 
.A(n_108),
.Y(n_107)
);

BUFx6f_ASAP7_75t_L g327 ( 
.A(n_108),
.Y(n_327)
);

XOR2xp5_ASAP7_75t_L g238 ( 
.A(n_110),
.B(n_151),
.Y(n_238)
);

OAI22x1_ASAP7_75t_SL g110 ( 
.A1(n_111),
.A2(n_133),
.B1(n_142),
.B2(n_149),
.Y(n_110)
);

OAI22x1_ASAP7_75t_L g226 ( 
.A1(n_111),
.A2(n_142),
.B1(n_149),
.B2(n_227),
.Y(n_226)
);

OAI22xp5_ASAP7_75t_L g243 ( 
.A1(n_111),
.A2(n_133),
.B1(n_149),
.B2(n_244),
.Y(n_243)
);

OAI22xp5_ASAP7_75t_SL g569 ( 
.A1(n_111),
.A2(n_149),
.B1(n_227),
.B2(n_570),
.Y(n_569)
);

INVx2_ASAP7_75t_L g111 ( 
.A(n_112),
.Y(n_111)
);

AOI22xp5_ASAP7_75t_L g335 ( 
.A1(n_112),
.A2(n_150),
.B1(n_336),
.B2(n_338),
.Y(n_335)
);

AOI22xp5_ASAP7_75t_L g355 ( 
.A1(n_112),
.A2(n_150),
.B1(n_336),
.B2(n_356),
.Y(n_355)
);

OA21x2_ASAP7_75t_L g112 ( 
.A1(n_113),
.A2(n_119),
.B(n_123),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_L g113 ( 
.A(n_114),
.B(n_117),
.Y(n_113)
);

AOI22xp5_ASAP7_75t_SL g123 ( 
.A1(n_114),
.A2(n_124),
.B1(n_127),
.B2(n_131),
.Y(n_123)
);

INVx6_ASAP7_75t_L g114 ( 
.A(n_115),
.Y(n_114)
);

INVx4_ASAP7_75t_L g115 ( 
.A(n_116),
.Y(n_115)
);

BUFx6f_ASAP7_75t_L g316 ( 
.A(n_116),
.Y(n_316)
);

BUFx3_ASAP7_75t_L g357 ( 
.A(n_117),
.Y(n_357)
);

BUFx6f_ASAP7_75t_L g117 ( 
.A(n_118),
.Y(n_117)
);

BUFx6f_ASAP7_75t_L g120 ( 
.A(n_118),
.Y(n_120)
);

BUFx6f_ASAP7_75t_L g144 ( 
.A(n_118),
.Y(n_144)
);

INVxp67_ASAP7_75t_L g320 ( 
.A(n_119),
.Y(n_320)
);

AND2x2_ASAP7_75t_L g119 ( 
.A(n_120),
.B(n_121),
.Y(n_119)
);

INVx2_ASAP7_75t_L g121 ( 
.A(n_122),
.Y(n_121)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_123),
.Y(n_150)
);

INVx2_ASAP7_75t_L g124 ( 
.A(n_125),
.Y(n_124)
);

INVx2_ASAP7_75t_L g125 ( 
.A(n_126),
.Y(n_125)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_128),
.Y(n_127)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_129),
.Y(n_128)
);

INVx2_ASAP7_75t_SL g306 ( 
.A(n_129),
.Y(n_306)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_130),
.Y(n_129)
);

INVx4_ASAP7_75t_L g132 ( 
.A(n_130),
.Y(n_132)
);

BUFx6f_ASAP7_75t_L g154 ( 
.A(n_130),
.Y(n_154)
);

INVx4_ASAP7_75t_L g284 ( 
.A(n_131),
.Y(n_284)
);

INVx6_ASAP7_75t_L g131 ( 
.A(n_132),
.Y(n_131)
);

INVx4_ASAP7_75t_L g134 ( 
.A(n_135),
.Y(n_134)
);

INVx5_ASAP7_75t_L g135 ( 
.A(n_136),
.Y(n_135)
);

INVx8_ASAP7_75t_L g148 ( 
.A(n_136),
.Y(n_148)
);

INVx4_ASAP7_75t_L g312 ( 
.A(n_136),
.Y(n_312)
);

BUFx6f_ASAP7_75t_L g136 ( 
.A(n_137),
.Y(n_136)
);

BUFx6f_ASAP7_75t_L g247 ( 
.A(n_137),
.Y(n_247)
);

INVx2_ASAP7_75t_L g139 ( 
.A(n_140),
.Y(n_139)
);

INVx3_ASAP7_75t_L g140 ( 
.A(n_141),
.Y(n_140)
);

INVx5_ASAP7_75t_L g143 ( 
.A(n_144),
.Y(n_143)
);

INVx2_ASAP7_75t_L g571 ( 
.A(n_146),
.Y(n_571)
);

INVx3_ASAP7_75t_L g146 ( 
.A(n_147),
.Y(n_146)
);

INVx6_ASAP7_75t_L g147 ( 
.A(n_148),
.Y(n_147)
);

BUFx2_ASAP7_75t_L g572 ( 
.A(n_148),
.Y(n_572)
);

INVx2_ASAP7_75t_L g149 ( 
.A(n_150),
.Y(n_149)
);

OAI22xp5_ASAP7_75t_L g151 ( 
.A1(n_152),
.A2(n_160),
.B1(n_187),
.B2(n_189),
.Y(n_151)
);

OAI22xp5_ASAP7_75t_L g275 ( 
.A1(n_152),
.A2(n_160),
.B1(n_187),
.B2(n_276),
.Y(n_275)
);

INVx6_ASAP7_75t_L g354 ( 
.A(n_153),
.Y(n_354)
);

INVx6_ASAP7_75t_L g153 ( 
.A(n_154),
.Y(n_153)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_155),
.Y(n_190)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_156),
.Y(n_155)
);

INVx2_ASAP7_75t_L g204 ( 
.A(n_156),
.Y(n_204)
);

INVx2_ASAP7_75t_L g156 ( 
.A(n_157),
.Y(n_156)
);

BUFx3_ASAP7_75t_L g381 ( 
.A(n_157),
.Y(n_381)
);

BUFx6f_ASAP7_75t_L g157 ( 
.A(n_158),
.Y(n_157)
);

INVx2_ASAP7_75t_L g169 ( 
.A(n_158),
.Y(n_169)
);

BUFx6f_ASAP7_75t_L g281 ( 
.A(n_158),
.Y(n_281)
);

BUFx5_ASAP7_75t_L g303 ( 
.A(n_158),
.Y(n_303)
);

BUFx6f_ASAP7_75t_L g379 ( 
.A(n_158),
.Y(n_379)
);

INVx2_ASAP7_75t_L g197 ( 
.A(n_160),
.Y(n_197)
);

OAI22xp5_ASAP7_75t_L g296 ( 
.A1(n_160),
.A2(n_187),
.B1(n_276),
.B2(n_297),
.Y(n_296)
);

OAI22xp5_ASAP7_75t_SL g523 ( 
.A1(n_160),
.A2(n_187),
.B1(n_375),
.B2(n_524),
.Y(n_523)
);

OAI22xp5_ASAP7_75t_L g574 ( 
.A1(n_160),
.A2(n_187),
.B1(n_200),
.B2(n_575),
.Y(n_574)
);

AO21x2_ASAP7_75t_SL g160 ( 
.A1(n_161),
.A2(n_170),
.B(n_176),
.Y(n_160)
);

NAND2xp33_ASAP7_75t_SL g161 ( 
.A(n_162),
.B(n_166),
.Y(n_161)
);

BUFx2_ASAP7_75t_L g162 ( 
.A(n_163),
.Y(n_162)
);

INVx3_ASAP7_75t_L g163 ( 
.A(n_164),
.Y(n_163)
);

BUFx6f_ASAP7_75t_L g164 ( 
.A(n_165),
.Y(n_164)
);

INVx2_ASAP7_75t_L g166 ( 
.A(n_167),
.Y(n_166)
);

INVx2_ASAP7_75t_L g167 ( 
.A(n_168),
.Y(n_167)
);

INVx4_ASAP7_75t_L g175 ( 
.A(n_168),
.Y(n_175)
);

INVx1_ASAP7_75t_L g515 ( 
.A(n_168),
.Y(n_515)
);

BUFx6f_ASAP7_75t_L g527 ( 
.A(n_168),
.Y(n_527)
);

BUFx6f_ASAP7_75t_L g168 ( 
.A(n_169),
.Y(n_168)
);

BUFx6f_ASAP7_75t_L g193 ( 
.A(n_169),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_L g170 ( 
.A(n_171),
.B(n_175),
.Y(n_170)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_172),
.Y(n_171)
);

INVx2_ASAP7_75t_L g172 ( 
.A(n_173),
.Y(n_172)
);

BUFx3_ASAP7_75t_L g173 ( 
.A(n_174),
.Y(n_173)
);

BUFx3_ASAP7_75t_L g188 ( 
.A(n_176),
.Y(n_188)
);

OAI22xp5_ASAP7_75t_L g176 ( 
.A1(n_177),
.A2(n_179),
.B1(n_182),
.B2(n_184),
.Y(n_176)
);

BUFx6f_ASAP7_75t_L g360 ( 
.A(n_177),
.Y(n_360)
);

INVx5_ASAP7_75t_L g177 ( 
.A(n_178),
.Y(n_177)
);

INVx6_ASAP7_75t_L g179 ( 
.A(n_180),
.Y(n_179)
);

BUFx6f_ASAP7_75t_L g180 ( 
.A(n_181),
.Y(n_180)
);

BUFx6f_ASAP7_75t_L g186 ( 
.A(n_181),
.Y(n_186)
);

INVx3_ASAP7_75t_L g216 ( 
.A(n_182),
.Y(n_216)
);

INVx2_ASAP7_75t_L g219 ( 
.A(n_182),
.Y(n_219)
);

INVx4_ASAP7_75t_L g182 ( 
.A(n_183),
.Y(n_182)
);

BUFx12f_ASAP7_75t_L g258 ( 
.A(n_183),
.Y(n_258)
);

INVx3_ASAP7_75t_L g184 ( 
.A(n_185),
.Y(n_184)
);

INVx3_ASAP7_75t_L g185 ( 
.A(n_186),
.Y(n_185)
);

INVx2_ASAP7_75t_L g187 ( 
.A(n_188),
.Y(n_187)
);

AOI22xp5_ASAP7_75t_SL g196 ( 
.A1(n_188),
.A2(n_197),
.B1(n_198),
.B2(n_199),
.Y(n_196)
);

AOI22xp5_ASAP7_75t_L g349 ( 
.A1(n_188),
.A2(n_197),
.B1(n_298),
.B2(n_350),
.Y(n_349)
);

AOI22xp5_ASAP7_75t_SL g373 ( 
.A1(n_188),
.A2(n_197),
.B1(n_350),
.B2(n_374),
.Y(n_373)
);

INVxp67_ASAP7_75t_L g198 ( 
.A(n_189),
.Y(n_198)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_191),
.Y(n_317)
);

BUFx2_ASAP7_75t_L g191 ( 
.A(n_192),
.Y(n_191)
);

INVx2_ASAP7_75t_L g206 ( 
.A(n_192),
.Y(n_206)
);

INVx4_ASAP7_75t_L g192 ( 
.A(n_193),
.Y(n_192)
);

XNOR2xp5_ASAP7_75t_L g194 ( 
.A(n_195),
.B(n_221),
.Y(n_194)
);

INVx1_ASAP7_75t_L g563 ( 
.A(n_195),
.Y(n_563)
);

OAI21xp5_ASAP7_75t_SL g195 ( 
.A1(n_196),
.A2(n_207),
.B(n_220),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_L g220 ( 
.A(n_196),
.B(n_207),
.Y(n_220)
);

INVxp67_ASAP7_75t_L g199 ( 
.A(n_200),
.Y(n_199)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_202),
.Y(n_201)
);

INVx2_ASAP7_75t_L g202 ( 
.A(n_203),
.Y(n_202)
);

INVx3_ASAP7_75t_L g203 ( 
.A(n_204),
.Y(n_203)
);

INVx1_ASAP7_75t_L g525 ( 
.A(n_205),
.Y(n_525)
);

INVx3_ASAP7_75t_L g205 ( 
.A(n_206),
.Y(n_205)
);

INVxp67_ASAP7_75t_L g208 ( 
.A(n_209),
.Y(n_208)
);

INVx2_ASAP7_75t_L g210 ( 
.A(n_211),
.Y(n_210)
);

HB1xp67_ASAP7_75t_L g211 ( 
.A(n_212),
.Y(n_211)
);

INVx2_ASAP7_75t_L g212 ( 
.A(n_213),
.Y(n_212)
);

INVx2_ASAP7_75t_L g512 ( 
.A(n_213),
.Y(n_512)
);

INVx3_ASAP7_75t_L g213 ( 
.A(n_214),
.Y(n_213)
);

HB1xp67_ASAP7_75t_L g215 ( 
.A(n_216),
.Y(n_215)
);

INVx2_ASAP7_75t_L g218 ( 
.A(n_219),
.Y(n_218)
);

AOI22xp5_ASAP7_75t_L g566 ( 
.A1(n_220),
.A2(n_567),
.B1(n_580),
.B2(n_581),
.Y(n_566)
);

INVx1_ASAP7_75t_L g580 ( 
.A(n_220),
.Y(n_580)
);

INVxp67_ASAP7_75t_L g562 ( 
.A(n_221),
.Y(n_562)
);

OAI22xp5_ASAP7_75t_SL g221 ( 
.A1(n_222),
.A2(n_223),
.B1(n_230),
.B2(n_234),
.Y(n_221)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_223),
.Y(n_222)
);

XNOR2xp5_ASAP7_75t_SL g223 ( 
.A(n_224),
.B(n_226),
.Y(n_223)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_224),
.Y(n_231)
);

OAI22xp5_ASAP7_75t_SL g239 ( 
.A1(n_224),
.A2(n_231),
.B1(n_232),
.B2(n_240),
.Y(n_239)
);

AOI22xp5_ASAP7_75t_SL g565 ( 
.A1(n_224),
.A2(n_226),
.B1(n_234),
.B2(n_584),
.Y(n_565)
);

BUFx6f_ASAP7_75t_L g228 ( 
.A(n_229),
.Y(n_228)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_230),
.Y(n_234)
);

NAND2xp5_ASAP7_75t_L g230 ( 
.A(n_231),
.B(n_232),
.Y(n_230)
);

INVxp67_ASAP7_75t_L g240 ( 
.A(n_232),
.Y(n_240)
);

MAJIxp5_ASAP7_75t_L g235 ( 
.A(n_236),
.B(n_239),
.C(n_241),
.Y(n_235)
);

AOI22xp5_ASAP7_75t_L g287 ( 
.A1(n_236),
.A2(n_237),
.B1(n_239),
.B2(n_288),
.Y(n_287)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_237),
.Y(n_236)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_239),
.Y(n_288)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_242),
.Y(n_241)
);

XNOR2xp5_ASAP7_75t_L g286 ( 
.A(n_242),
.B(n_287),
.Y(n_286)
);

MAJIxp5_ASAP7_75t_L g242 ( 
.A(n_243),
.B(n_253),
.C(n_275),
.Y(n_242)
);

XOR2xp5_ASAP7_75t_L g291 ( 
.A(n_243),
.B(n_275),
.Y(n_291)
);

INVx1_ASAP7_75t_L g338 ( 
.A(n_244),
.Y(n_338)
);

INVx3_ASAP7_75t_L g245 ( 
.A(n_246),
.Y(n_245)
);

INVx4_ASAP7_75t_L g246 ( 
.A(n_247),
.Y(n_246)
);

INVx6_ASAP7_75t_L g252 ( 
.A(n_247),
.Y(n_252)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_250),
.Y(n_249)
);

INVx3_ASAP7_75t_L g250 ( 
.A(n_251),
.Y(n_250)
);

BUFx6f_ASAP7_75t_L g251 ( 
.A(n_252),
.Y(n_251)
);

INVxp67_ASAP7_75t_L g253 ( 
.A(n_254),
.Y(n_253)
);

XNOR2xp5_ASAP7_75t_L g290 ( 
.A(n_254),
.B(n_291),
.Y(n_290)
);

NAND2xp5_ASAP7_75t_SL g254 ( 
.A(n_255),
.B(n_261),
.Y(n_254)
);

XOR2xp5_ASAP7_75t_L g346 ( 
.A(n_255),
.B(n_261),
.Y(n_346)
);

INVx1_ASAP7_75t_L g366 ( 
.A(n_256),
.Y(n_366)
);

INVx2_ASAP7_75t_L g257 ( 
.A(n_258),
.Y(n_257)
);

INVx1_ASAP7_75t_SL g463 ( 
.A(n_258),
.Y(n_463)
);

INVx1_ASAP7_75t_L g517 ( 
.A(n_259),
.Y(n_517)
);

HB1xp67_ASAP7_75t_L g259 ( 
.A(n_260),
.Y(n_259)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_264),
.Y(n_263)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_265),
.Y(n_264)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_266),
.Y(n_265)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_268),
.Y(n_267)
);

INVx1_ASAP7_75t_SL g268 ( 
.A(n_269),
.Y(n_268)
);

INVx2_ASAP7_75t_L g269 ( 
.A(n_270),
.Y(n_269)
);

INVx2_ASAP7_75t_SL g270 ( 
.A(n_271),
.Y(n_270)
);

INVx1_ASAP7_75t_L g470 ( 
.A(n_271),
.Y(n_470)
);

INVx2_ASAP7_75t_L g272 ( 
.A(n_273),
.Y(n_272)
);

BUFx6f_ASAP7_75t_L g273 ( 
.A(n_274),
.Y(n_273)
);

INVx6_ASAP7_75t_L g472 ( 
.A(n_274),
.Y(n_472)
);

BUFx2_ASAP7_75t_L g277 ( 
.A(n_278),
.Y(n_277)
);

INVx2_ASAP7_75t_L g278 ( 
.A(n_279),
.Y(n_278)
);

INVx2_ASAP7_75t_L g279 ( 
.A(n_280),
.Y(n_279)
);

INVx4_ASAP7_75t_L g280 ( 
.A(n_281),
.Y(n_280)
);

BUFx6f_ASAP7_75t_L g352 ( 
.A(n_281),
.Y(n_352)
);

INVx2_ASAP7_75t_L g577 ( 
.A(n_281),
.Y(n_577)
);

HB1xp67_ASAP7_75t_L g282 ( 
.A(n_283),
.Y(n_282)
);

INVx2_ASAP7_75t_L g319 ( 
.A(n_283),
.Y(n_319)
);

INVx5_ASAP7_75t_L g283 ( 
.A(n_284),
.Y(n_283)
);

NAND2xp5_ASAP7_75t_SL g285 ( 
.A(n_286),
.B(n_289),
.Y(n_285)
);

NOR2xp33_ASAP7_75t_L g557 ( 
.A(n_286),
.B(n_289),
.Y(n_557)
);

MAJIxp5_ASAP7_75t_L g289 ( 
.A(n_290),
.B(n_292),
.C(n_294),
.Y(n_289)
);

XOR2xp5_ASAP7_75t_L g341 ( 
.A(n_290),
.B(n_292),
.Y(n_341)
);

XNOR2xp5_ASAP7_75t_L g340 ( 
.A(n_294),
.B(n_341),
.Y(n_340)
);

MAJIxp5_ASAP7_75t_L g294 ( 
.A(n_295),
.B(n_307),
.C(n_335),
.Y(n_294)
);

INVxp67_ASAP7_75t_L g295 ( 
.A(n_296),
.Y(n_295)
);

XNOR2xp5_ASAP7_75t_L g345 ( 
.A(n_296),
.B(n_335),
.Y(n_345)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_298),
.Y(n_297)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_300),
.Y(n_299)
);

INVx3_ASAP7_75t_L g300 ( 
.A(n_301),
.Y(n_300)
);

INVx2_ASAP7_75t_L g301 ( 
.A(n_302),
.Y(n_301)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_303),
.Y(n_302)
);

INVx1_ASAP7_75t_SL g304 ( 
.A(n_305),
.Y(n_304)
);

BUFx3_ASAP7_75t_L g305 ( 
.A(n_306),
.Y(n_305)
);

XOR2xp5_ASAP7_75t_L g344 ( 
.A(n_307),
.B(n_345),
.Y(n_344)
);

NAND2xp5_ASAP7_75t_L g307 ( 
.A(n_308),
.B(n_321),
.Y(n_307)
);

XOR2xp5_ASAP7_75t_L g371 ( 
.A(n_308),
.B(n_321),
.Y(n_371)
);

OAI22xp5_ASAP7_75t_L g308 ( 
.A1(n_309),
.A2(n_313),
.B1(n_318),
.B2(n_320),
.Y(n_308)
);

OAI21xp33_ASAP7_75t_SL g356 ( 
.A1(n_309),
.A2(n_310),
.B(n_357),
.Y(n_356)
);

NAND2xp5_ASAP7_75t_L g309 ( 
.A(n_310),
.B(n_311),
.Y(n_309)
);

NAND2xp5_ASAP7_75t_L g416 ( 
.A(n_310),
.B(n_360),
.Y(n_416)
);

OAI21xp33_ASAP7_75t_SL g422 ( 
.A1(n_310),
.A2(n_416),
.B(n_423),
.Y(n_422)
);

NOR2xp33_ASAP7_75t_SL g481 ( 
.A(n_310),
.B(n_482),
.Y(n_481)
);

NOR2xp33_ASAP7_75t_L g516 ( 
.A(n_310),
.B(n_517),
.Y(n_516)
);

BUFx6f_ASAP7_75t_L g311 ( 
.A(n_312),
.Y(n_311)
);

NOR2xp33_ASAP7_75t_L g313 ( 
.A(n_314),
.B(n_317),
.Y(n_313)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_315),
.Y(n_314)
);

INVx2_ASAP7_75t_L g315 ( 
.A(n_316),
.Y(n_315)
);

INVx2_ASAP7_75t_L g318 ( 
.A(n_319),
.Y(n_318)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_323),
.Y(n_322)
);

INVx2_ASAP7_75t_L g324 ( 
.A(n_325),
.Y(n_324)
);

BUFx6f_ASAP7_75t_L g325 ( 
.A(n_326),
.Y(n_325)
);

INVx4_ASAP7_75t_L g326 ( 
.A(n_327),
.Y(n_326)
);

BUFx6f_ASAP7_75t_L g497 ( 
.A(n_327),
.Y(n_497)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_329),
.Y(n_328)
);

BUFx2_ASAP7_75t_L g329 ( 
.A(n_330),
.Y(n_329)
);

INVx3_ASAP7_75t_L g330 ( 
.A(n_331),
.Y(n_330)
);

INVx5_ASAP7_75t_L g331 ( 
.A(n_332),
.Y(n_331)
);

INVx4_ASAP7_75t_L g332 ( 
.A(n_333),
.Y(n_332)
);

INVx3_ASAP7_75t_L g333 ( 
.A(n_334),
.Y(n_333)
);

BUFx3_ASAP7_75t_L g501 ( 
.A(n_334),
.Y(n_501)
);

AOI21xp5_ASAP7_75t_L g339 ( 
.A1(n_340),
.A2(n_342),
.B(n_367),
.Y(n_339)
);

MAJIxp5_ASAP7_75t_L g555 ( 
.A(n_340),
.B(n_342),
.C(n_556),
.Y(n_555)
);

MAJIxp5_ASAP7_75t_L g342 ( 
.A(n_343),
.B(n_346),
.C(n_347),
.Y(n_342)
);

AOI22xp5_ASAP7_75t_L g396 ( 
.A1(n_343),
.A2(n_344),
.B1(n_397),
.B2(n_398),
.Y(n_396)
);

INVx1_ASAP7_75t_L g343 ( 
.A(n_344),
.Y(n_343)
);

XNOR2xp5_ASAP7_75t_L g397 ( 
.A(n_346),
.B(n_348),
.Y(n_397)
);

HB1xp67_ASAP7_75t_L g347 ( 
.A(n_348),
.Y(n_347)
);

MAJIxp5_ASAP7_75t_L g348 ( 
.A(n_349),
.B(n_355),
.C(n_358),
.Y(n_348)
);

XNOR2xp5_ASAP7_75t_L g370 ( 
.A(n_349),
.B(n_358),
.Y(n_370)
);

BUFx3_ASAP7_75t_L g351 ( 
.A(n_352),
.Y(n_351)
);

INVx1_ASAP7_75t_SL g353 ( 
.A(n_354),
.Y(n_353)
);

XOR2xp5_ASAP7_75t_L g369 ( 
.A(n_355),
.B(n_370),
.Y(n_369)
);

INVxp67_ASAP7_75t_L g543 ( 
.A(n_359),
.Y(n_543)
);

INVx2_ASAP7_75t_L g361 ( 
.A(n_362),
.Y(n_361)
);

INVx3_ASAP7_75t_L g362 ( 
.A(n_363),
.Y(n_362)
);

INVx2_ASAP7_75t_L g363 ( 
.A(n_364),
.Y(n_363)
);

BUFx6f_ASAP7_75t_L g364 ( 
.A(n_365),
.Y(n_364)
);

AND2x2_ASAP7_75t_L g367 ( 
.A(n_368),
.B(n_396),
.Y(n_367)
);

OR2x2_ASAP7_75t_L g556 ( 
.A(n_368),
.B(n_396),
.Y(n_556)
);

MAJIxp5_ASAP7_75t_L g368 ( 
.A(n_369),
.B(n_371),
.C(n_372),
.Y(n_368)
);

XOR2xp5_ASAP7_75t_L g549 ( 
.A(n_369),
.B(n_550),
.Y(n_549)
);

XNOR2xp5_ASAP7_75t_L g550 ( 
.A(n_371),
.B(n_551),
.Y(n_550)
);

MAJIxp5_ASAP7_75t_L g372 ( 
.A(n_373),
.B(n_382),
.C(n_395),
.Y(n_372)
);

XOR2xp5_ASAP7_75t_SL g536 ( 
.A(n_373),
.B(n_537),
.Y(n_536)
);

MAJIxp5_ASAP7_75t_L g551 ( 
.A(n_373),
.B(n_382),
.C(n_395),
.Y(n_551)
);

INVx1_ASAP7_75t_L g374 ( 
.A(n_375),
.Y(n_374)
);

INVx1_ASAP7_75t_L g376 ( 
.A(n_377),
.Y(n_376)
);

BUFx2_ASAP7_75t_L g377 ( 
.A(n_378),
.Y(n_377)
);

BUFx6f_ASAP7_75t_L g378 ( 
.A(n_379),
.Y(n_378)
);

BUFx6f_ASAP7_75t_L g380 ( 
.A(n_381),
.Y(n_380)
);

XOR2xp5_ASAP7_75t_SL g537 ( 
.A(n_382),
.B(n_395),
.Y(n_537)
);

INVx1_ASAP7_75t_L g384 ( 
.A(n_385),
.Y(n_384)
);

INVx1_ASAP7_75t_L g385 ( 
.A(n_386),
.Y(n_385)
);

INVx1_ASAP7_75t_L g386 ( 
.A(n_387),
.Y(n_386)
);

INVx3_ASAP7_75t_L g442 ( 
.A(n_387),
.Y(n_442)
);

INVx1_ASAP7_75t_L g388 ( 
.A(n_389),
.Y(n_388)
);

INVx1_ASAP7_75t_L g389 ( 
.A(n_390),
.Y(n_389)
);

INVx1_ASAP7_75t_L g390 ( 
.A(n_391),
.Y(n_390)
);

INVx1_ASAP7_75t_L g392 ( 
.A(n_393),
.Y(n_392)
);

INVx3_ASAP7_75t_L g393 ( 
.A(n_394),
.Y(n_393)
);

INVx1_ASAP7_75t_L g398 ( 
.A(n_397),
.Y(n_398)
);

AOI21x1_ASAP7_75t_L g399 ( 
.A1(n_400),
.A2(n_548),
.B(n_553),
.Y(n_399)
);

OAI21x1_ASAP7_75t_L g400 ( 
.A1(n_401),
.A2(n_533),
.B(n_547),
.Y(n_400)
);

AOI21x1_ASAP7_75t_L g401 ( 
.A1(n_402),
.A2(n_506),
.B(n_532),
.Y(n_401)
);

OAI21x1_ASAP7_75t_L g402 ( 
.A1(n_403),
.A2(n_465),
.B(n_505),
.Y(n_402)
);

AND2x2_ASAP7_75t_L g403 ( 
.A(n_404),
.B(n_433),
.Y(n_403)
);

OR2x2_ASAP7_75t_L g505 ( 
.A(n_404),
.B(n_433),
.Y(n_505)
);

NAND2xp5_ASAP7_75t_L g404 ( 
.A(n_405),
.B(n_420),
.Y(n_404)
);

AOI22xp5_ASAP7_75t_L g474 ( 
.A1(n_405),
.A2(n_420),
.B1(n_421),
.B2(n_475),
.Y(n_474)
);

INVx1_ASAP7_75t_L g475 ( 
.A(n_405),
.Y(n_475)
);

OAI32xp33_ASAP7_75t_L g405 ( 
.A1(n_406),
.A2(n_410),
.A3(n_412),
.B1(n_416),
.B2(n_417),
.Y(n_405)
);

INVx2_ASAP7_75t_L g406 ( 
.A(n_407),
.Y(n_406)
);

INVx2_ASAP7_75t_L g407 ( 
.A(n_408),
.Y(n_407)
);

INVx2_ASAP7_75t_L g408 ( 
.A(n_409),
.Y(n_408)
);

INVx3_ASAP7_75t_L g410 ( 
.A(n_411),
.Y(n_410)
);

INVx1_ASAP7_75t_L g412 ( 
.A(n_413),
.Y(n_412)
);

NOR2xp33_ASAP7_75t_L g417 ( 
.A(n_413),
.B(n_418),
.Y(n_417)
);

INVx1_ASAP7_75t_L g413 ( 
.A(n_414),
.Y(n_413)
);

INVx2_ASAP7_75t_L g414 ( 
.A(n_415),
.Y(n_414)
);

INVx2_ASAP7_75t_L g418 ( 
.A(n_419),
.Y(n_418)
);

INVx1_ASAP7_75t_L g420 ( 
.A(n_421),
.Y(n_420)
);

BUFx2_ASAP7_75t_L g423 ( 
.A(n_424),
.Y(n_423)
);

INVx1_ASAP7_75t_L g424 ( 
.A(n_425),
.Y(n_424)
);

INVx1_ASAP7_75t_L g531 ( 
.A(n_425),
.Y(n_531)
);

INVx2_ASAP7_75t_L g427 ( 
.A(n_428),
.Y(n_427)
);

INVx4_ASAP7_75t_L g428 ( 
.A(n_429),
.Y(n_428)
);

BUFx6f_ASAP7_75t_L g429 ( 
.A(n_430),
.Y(n_429)
);

INVx1_ASAP7_75t_L g432 ( 
.A(n_430),
.Y(n_432)
);

BUFx2_ASAP7_75t_L g431 ( 
.A(n_432),
.Y(n_431)
);

XNOR2xp5_ASAP7_75t_L g433 ( 
.A(n_434),
.B(n_455),
.Y(n_433)
);

MAJIxp5_ASAP7_75t_L g507 ( 
.A(n_434),
.B(n_457),
.C(n_464),
.Y(n_507)
);

INVxp67_ASAP7_75t_L g473 ( 
.A(n_435),
.Y(n_473)
);

BUFx2_ASAP7_75t_L g436 ( 
.A(n_437),
.Y(n_436)
);

INVx1_ASAP7_75t_L g437 ( 
.A(n_438),
.Y(n_437)
);

INVx2_ASAP7_75t_L g438 ( 
.A(n_439),
.Y(n_438)
);

INVx1_ASAP7_75t_L g440 ( 
.A(n_441),
.Y(n_440)
);

INVx2_ASAP7_75t_L g441 ( 
.A(n_442),
.Y(n_441)
);

INVx1_ASAP7_75t_L g450 ( 
.A(n_442),
.Y(n_450)
);

INVx1_ASAP7_75t_L g443 ( 
.A(n_444),
.Y(n_443)
);

BUFx2_ASAP7_75t_L g444 ( 
.A(n_445),
.Y(n_444)
);

INVx2_ASAP7_75t_L g445 ( 
.A(n_446),
.Y(n_445)
);

INVxp67_ASAP7_75t_L g447 ( 
.A(n_448),
.Y(n_447)
);

INVx2_ASAP7_75t_L g449 ( 
.A(n_450),
.Y(n_449)
);

INVx1_ASAP7_75t_L g480 ( 
.A(n_451),
.Y(n_480)
);

HB1xp67_ASAP7_75t_L g451 ( 
.A(n_452),
.Y(n_451)
);

INVx2_ASAP7_75t_L g452 ( 
.A(n_453),
.Y(n_452)
);

BUFx6f_ASAP7_75t_L g453 ( 
.A(n_454),
.Y(n_453)
);

OAI22xp5_ASAP7_75t_L g455 ( 
.A1(n_456),
.A2(n_457),
.B1(n_458),
.B2(n_464),
.Y(n_455)
);

INVx1_ASAP7_75t_L g464 ( 
.A(n_456),
.Y(n_464)
);

INVx1_ASAP7_75t_L g457 ( 
.A(n_458),
.Y(n_457)
);

INVx1_ASAP7_75t_L g460 ( 
.A(n_461),
.Y(n_460)
);

INVx4_ASAP7_75t_L g461 ( 
.A(n_462),
.Y(n_461)
);

AOI21xp5_ASAP7_75t_L g465 ( 
.A1(n_466),
.A2(n_476),
.B(n_504),
.Y(n_465)
);

NAND2xp5_ASAP7_75t_L g466 ( 
.A(n_467),
.B(n_474),
.Y(n_466)
);

NOR2xp33_ASAP7_75t_L g504 ( 
.A(n_467),
.B(n_474),
.Y(n_504)
);

INVxp67_ASAP7_75t_L g468 ( 
.A(n_469),
.Y(n_468)
);

INVx6_ASAP7_75t_L g471 ( 
.A(n_472),
.Y(n_471)
);

OAI21xp5_ASAP7_75t_L g476 ( 
.A1(n_477),
.A2(n_498),
.B(n_503),
.Y(n_476)
);

NAND2xp5_ASAP7_75t_L g477 ( 
.A(n_478),
.B(n_487),
.Y(n_477)
);

NOR2xp33_ASAP7_75t_L g478 ( 
.A(n_479),
.B(n_481),
.Y(n_478)
);

INVx1_ASAP7_75t_L g479 ( 
.A(n_480),
.Y(n_479)
);

INVx1_ASAP7_75t_L g482 ( 
.A(n_483),
.Y(n_482)
);

INVx4_ASAP7_75t_L g483 ( 
.A(n_484),
.Y(n_483)
);

INVx6_ASAP7_75t_L g484 ( 
.A(n_485),
.Y(n_484)
);

BUFx12f_ASAP7_75t_L g485 ( 
.A(n_486),
.Y(n_485)
);

INVx2_ASAP7_75t_L g489 ( 
.A(n_490),
.Y(n_489)
);

BUFx3_ASAP7_75t_L g490 ( 
.A(n_491),
.Y(n_490)
);

INVx2_ASAP7_75t_L g491 ( 
.A(n_492),
.Y(n_491)
);

INVx2_ASAP7_75t_L g492 ( 
.A(n_493),
.Y(n_492)
);

INVx2_ASAP7_75t_L g493 ( 
.A(n_494),
.Y(n_493)
);

INVx1_ASAP7_75t_L g495 ( 
.A(n_496),
.Y(n_495)
);

BUFx3_ASAP7_75t_L g496 ( 
.A(n_497),
.Y(n_496)
);

NOR2xp33_ASAP7_75t_L g498 ( 
.A(n_499),
.B(n_502),
.Y(n_498)
);

NAND2xp5_ASAP7_75t_L g503 ( 
.A(n_499),
.B(n_502),
.Y(n_503)
);

INVx1_ASAP7_75t_L g500 ( 
.A(n_501),
.Y(n_500)
);

NAND2xp5_ASAP7_75t_L g506 ( 
.A(n_507),
.B(n_508),
.Y(n_506)
);

NOR2xp33_ASAP7_75t_L g532 ( 
.A(n_507),
.B(n_508),
.Y(n_532)
);

XOR2xp5_ASAP7_75t_L g508 ( 
.A(n_509),
.B(n_521),
.Y(n_508)
);

MAJIxp5_ASAP7_75t_L g546 ( 
.A(n_509),
.B(n_522),
.C(n_529),
.Y(n_546)
);

AOI22xp5_ASAP7_75t_L g509 ( 
.A1(n_510),
.A2(n_518),
.B1(n_519),
.B2(n_520),
.Y(n_509)
);

INVx1_ASAP7_75t_L g519 ( 
.A(n_510),
.Y(n_519)
);

NAND2xp5_ASAP7_75t_L g540 ( 
.A(n_510),
.B(n_520),
.Y(n_540)
);

BUFx3_ASAP7_75t_L g511 ( 
.A(n_512),
.Y(n_511)
);

INVx8_ASAP7_75t_L g513 ( 
.A(n_514),
.Y(n_513)
);

BUFx6f_ASAP7_75t_L g514 ( 
.A(n_515),
.Y(n_514)
);

INVx1_ASAP7_75t_L g520 ( 
.A(n_518),
.Y(n_520)
);

OAI22xp5_ASAP7_75t_SL g521 ( 
.A1(n_522),
.A2(n_523),
.B1(n_528),
.B2(n_529),
.Y(n_521)
);

INVx1_ASAP7_75t_L g522 ( 
.A(n_523),
.Y(n_522)
);

INVx3_ASAP7_75t_L g526 ( 
.A(n_527),
.Y(n_526)
);

INVx1_ASAP7_75t_L g528 ( 
.A(n_529),
.Y(n_528)
);

INVxp67_ASAP7_75t_L g542 ( 
.A(n_530),
.Y(n_542)
);

NOR2xp67_ASAP7_75t_SL g533 ( 
.A(n_534),
.B(n_546),
.Y(n_533)
);

NAND2xp5_ASAP7_75t_L g547 ( 
.A(n_534),
.B(n_546),
.Y(n_547)
);

OAI22xp5_ASAP7_75t_SL g534 ( 
.A1(n_535),
.A2(n_536),
.B1(n_538),
.B2(n_539),
.Y(n_534)
);

MAJIxp5_ASAP7_75t_L g552 ( 
.A(n_535),
.B(n_541),
.C(n_544),
.Y(n_552)
);

INVx1_ASAP7_75t_L g535 ( 
.A(n_536),
.Y(n_535)
);

INVx1_ASAP7_75t_L g538 ( 
.A(n_539),
.Y(n_538)
);

OAI22xp5_ASAP7_75t_SL g539 ( 
.A1(n_540),
.A2(n_541),
.B1(n_544),
.B2(n_545),
.Y(n_539)
);

INVx1_ASAP7_75t_L g544 ( 
.A(n_540),
.Y(n_544)
);

INVx1_ASAP7_75t_L g545 ( 
.A(n_541),
.Y(n_545)
);

NAND2xp5_ASAP7_75t_SL g548 ( 
.A(n_549),
.B(n_552),
.Y(n_548)
);

NOR2xp33_ASAP7_75t_L g553 ( 
.A(n_549),
.B(n_552),
.Y(n_553)
);

NAND2xp5_ASAP7_75t_L g559 ( 
.A(n_560),
.B(n_582),
.Y(n_559)
);

OR2x2_ASAP7_75t_L g560 ( 
.A(n_561),
.B(n_564),
.Y(n_560)
);

NAND2xp5_ASAP7_75t_L g582 ( 
.A(n_561),
.B(n_564),
.Y(n_582)
);

XOR2xp5_ASAP7_75t_L g564 ( 
.A(n_565),
.B(n_566),
.Y(n_564)
);

INVx1_ASAP7_75t_L g581 ( 
.A(n_567),
.Y(n_581)
);

AOI22xp5_ASAP7_75t_L g567 ( 
.A1(n_568),
.A2(n_569),
.B1(n_573),
.B2(n_579),
.Y(n_567)
);

INVx1_ASAP7_75t_L g568 ( 
.A(n_569),
.Y(n_568)
);

INVx1_ASAP7_75t_L g579 ( 
.A(n_573),
.Y(n_579)
);

XNOR2xp5_ASAP7_75t_L g573 ( 
.A(n_574),
.B(n_578),
.Y(n_573)
);

INVx1_ASAP7_75t_L g576 ( 
.A(n_577),
.Y(n_576)
);


endmodule