module fake_jpeg_10179_n_225 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_225);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_225;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_223;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_24;
wire n_44;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_212;
wire n_131;
wire n_56;
wire n_211;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_216;
wire n_217;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

BUFx3_ASAP7_75t_L g15 ( 
.A(n_9),
.Y(n_15)
);

BUFx6f_ASAP7_75t_L g16 ( 
.A(n_2),
.Y(n_16)
);

INVx2_ASAP7_75t_L g17 ( 
.A(n_5),
.Y(n_17)
);

BUFx12f_ASAP7_75t_L g18 ( 
.A(n_8),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_5),
.Y(n_19)
);

INVx13_ASAP7_75t_L g20 ( 
.A(n_2),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_2),
.Y(n_21)
);

BUFx5_ASAP7_75t_L g22 ( 
.A(n_5),
.Y(n_22)
);

INVx8_ASAP7_75t_L g23 ( 
.A(n_3),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_7),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_1),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_7),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_3),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_14),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_0),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_7),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_18),
.Y(n_31)
);

INVx6_ASAP7_75t_L g42 ( 
.A(n_31),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g32 ( 
.A(n_20),
.B(n_0),
.Y(n_32)
);

NOR2xp33_ASAP7_75t_SL g61 ( 
.A(n_32),
.B(n_35),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_18),
.Y(n_33)
);

INVx6_ASAP7_75t_L g45 ( 
.A(n_33),
.Y(n_45)
);

INVx4_ASAP7_75t_L g34 ( 
.A(n_18),
.Y(n_34)
);

INVx11_ASAP7_75t_L g43 ( 
.A(n_34),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g35 ( 
.A(n_20),
.B(n_0),
.Y(n_35)
);

BUFx3_ASAP7_75t_L g36 ( 
.A(n_22),
.Y(n_36)
);

INVx3_ASAP7_75t_L g44 ( 
.A(n_36),
.Y(n_44)
);

INVx3_ASAP7_75t_L g37 ( 
.A(n_16),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g51 ( 
.A(n_37),
.B(n_38),
.Y(n_51)
);

INVx4_ASAP7_75t_L g38 ( 
.A(n_18),
.Y(n_38)
);

INVx3_ASAP7_75t_L g39 ( 
.A(n_16),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_39),
.B(n_41),
.Y(n_54)
);

BUFx3_ASAP7_75t_L g40 ( 
.A(n_22),
.Y(n_40)
);

CKINVDCx6p67_ASAP7_75t_R g55 ( 
.A(n_40),
.Y(n_55)
);

INVx3_ASAP7_75t_L g41 ( 
.A(n_16),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_32),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_SL g67 ( 
.A(n_46),
.B(n_52),
.Y(n_67)
);

AOI22xp33_ASAP7_75t_SL g47 ( 
.A1(n_37),
.A2(n_17),
.B1(n_23),
.B2(n_20),
.Y(n_47)
);

AOI22xp33_ASAP7_75t_SL g79 ( 
.A1(n_47),
.A2(n_58),
.B1(n_28),
.B2(n_24),
.Y(n_79)
);

AOI22xp33_ASAP7_75t_L g48 ( 
.A1(n_41),
.A2(n_17),
.B1(n_23),
.B2(n_30),
.Y(n_48)
);

OAI22xp5_ASAP7_75t_L g77 ( 
.A1(n_48),
.A2(n_29),
.B1(n_27),
.B2(n_28),
.Y(n_77)
);

AO22x2_ASAP7_75t_L g49 ( 
.A1(n_39),
.A2(n_22),
.B1(n_26),
.B2(n_25),
.Y(n_49)
);

AOI22xp5_ASAP7_75t_L g83 ( 
.A1(n_49),
.A2(n_19),
.B1(n_26),
.B2(n_16),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g50 ( 
.A(n_35),
.B(n_18),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_L g71 ( 
.A(n_50),
.B(n_53),
.Y(n_71)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_31),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_L g53 ( 
.A(n_31),
.B(n_25),
.Y(n_53)
);

AND2x2_ASAP7_75t_L g56 ( 
.A(n_36),
.B(n_21),
.Y(n_56)
);

OAI21xp33_ASAP7_75t_L g65 ( 
.A1(n_56),
.A2(n_59),
.B(n_46),
.Y(n_65)
);

OR2x2_ASAP7_75t_L g57 ( 
.A(n_34),
.B(n_30),
.Y(n_57)
);

NAND2xp33_ASAP7_75t_L g63 ( 
.A(n_57),
.B(n_15),
.Y(n_63)
);

AOI22xp33_ASAP7_75t_SL g58 ( 
.A1(n_38),
.A2(n_23),
.B1(n_21),
.B2(n_27),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_33),
.B(n_29),
.Y(n_59)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_33),
.Y(n_60)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_60),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_L g62 ( 
.A(n_40),
.B(n_25),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_L g72 ( 
.A(n_62),
.B(n_25),
.Y(n_72)
);

AND2x2_ASAP7_75t_L g105 ( 
.A(n_63),
.B(n_65),
.Y(n_105)
);

INVx4_ASAP7_75t_L g64 ( 
.A(n_43),
.Y(n_64)
);

INVx4_ASAP7_75t_L g91 ( 
.A(n_64),
.Y(n_91)
);

CKINVDCx20_ASAP7_75t_R g66 ( 
.A(n_42),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_66),
.B(n_68),
.Y(n_89)
);

INVx2_ASAP7_75t_L g68 ( 
.A(n_43),
.Y(n_68)
);

INVx8_ASAP7_75t_L g69 ( 
.A(n_55),
.Y(n_69)
);

AOI22xp33_ASAP7_75t_SL g102 ( 
.A1(n_69),
.A2(n_44),
.B1(n_45),
.B2(n_55),
.Y(n_102)
);

CKINVDCx20_ASAP7_75t_R g70 ( 
.A(n_42),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_70),
.B(n_74),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_L g92 ( 
.A(n_72),
.B(n_75),
.Y(n_92)
);

CKINVDCx20_ASAP7_75t_R g74 ( 
.A(n_42),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_L g75 ( 
.A(n_57),
.B(n_56),
.Y(n_75)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_54),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_76),
.B(n_78),
.Y(n_97)
);

AOI22xp33_ASAP7_75t_L g103 ( 
.A1(n_77),
.A2(n_45),
.B1(n_44),
.B2(n_55),
.Y(n_103)
);

INVx2_ASAP7_75t_L g78 ( 
.A(n_43),
.Y(n_78)
);

OAI22xp5_ASAP7_75t_L g100 ( 
.A1(n_79),
.A2(n_80),
.B1(n_50),
.B2(n_59),
.Y(n_100)
);

OAI22xp5_ASAP7_75t_L g80 ( 
.A1(n_49),
.A2(n_24),
.B1(n_19),
.B2(n_26),
.Y(n_80)
);

INVx5_ASAP7_75t_L g81 ( 
.A(n_55),
.Y(n_81)
);

INVx2_ASAP7_75t_L g96 ( 
.A(n_81),
.Y(n_96)
);

INVx2_ASAP7_75t_SL g82 ( 
.A(n_49),
.Y(n_82)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_82),
.Y(n_84)
);

OAI22xp5_ASAP7_75t_SL g86 ( 
.A1(n_83),
.A2(n_49),
.B1(n_53),
.B2(n_62),
.Y(n_86)
);

AOI22xp5_ASAP7_75t_L g85 ( 
.A1(n_82),
.A2(n_49),
.B1(n_54),
.B2(n_51),
.Y(n_85)
);

AOI22xp5_ASAP7_75t_L g107 ( 
.A1(n_85),
.A2(n_86),
.B1(n_90),
.B2(n_104),
.Y(n_107)
);

INVxp67_ASAP7_75t_L g87 ( 
.A(n_67),
.Y(n_87)
);

INVxp67_ASAP7_75t_L g118 ( 
.A(n_87),
.Y(n_118)
);

HB1xp67_ASAP7_75t_L g88 ( 
.A(n_68),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_88),
.B(n_95),
.Y(n_108)
);

OAI22xp5_ASAP7_75t_L g90 ( 
.A1(n_82),
.A2(n_49),
.B1(n_45),
.B2(n_60),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_L g93 ( 
.A(n_71),
.B(n_57),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_L g109 ( 
.A(n_93),
.B(n_98),
.Y(n_109)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_67),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g98 ( 
.A(n_71),
.B(n_56),
.Y(n_98)
);

CKINVDCx20_ASAP7_75t_R g99 ( 
.A(n_77),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g126 ( 
.A(n_99),
.B(n_69),
.Y(n_126)
);

AOI22xp5_ASAP7_75t_SL g123 ( 
.A1(n_100),
.A2(n_103),
.B1(n_104),
.B2(n_99),
.Y(n_123)
);

MAJIxp5_ASAP7_75t_L g101 ( 
.A(n_72),
.B(n_51),
.C(n_52),
.Y(n_101)
);

AND2x2_ASAP7_75t_L g112 ( 
.A(n_101),
.B(n_73),
.Y(n_112)
);

AOI21xp5_ASAP7_75t_L g113 ( 
.A1(n_102),
.A2(n_81),
.B(n_74),
.Y(n_113)
);

AO22x2_ASAP7_75t_L g104 ( 
.A1(n_63),
.A2(n_55),
.B1(n_26),
.B2(n_15),
.Y(n_104)
);

O2A1O1Ixp33_ASAP7_75t_L g106 ( 
.A1(n_84),
.A2(n_80),
.B(n_83),
.C(n_76),
.Y(n_106)
);

AOI22xp5_ASAP7_75t_L g134 ( 
.A1(n_106),
.A2(n_123),
.B1(n_126),
.B2(n_96),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_L g110 ( 
.A(n_92),
.B(n_75),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_L g138 ( 
.A(n_110),
.B(n_114),
.Y(n_138)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_94),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_SL g133 ( 
.A(n_111),
.B(n_112),
.Y(n_133)
);

INVxp67_ASAP7_75t_L g129 ( 
.A(n_113),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_L g114 ( 
.A(n_92),
.B(n_61),
.Y(n_114)
);

XNOR2x2_ASAP7_75t_L g115 ( 
.A(n_104),
.B(n_61),
.Y(n_115)
);

XOR2xp5_ASAP7_75t_L g130 ( 
.A(n_115),
.B(n_104),
.Y(n_130)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_89),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_SL g135 ( 
.A(n_116),
.B(n_117),
.Y(n_135)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_97),
.Y(n_117)
);

CKINVDCx20_ASAP7_75t_R g119 ( 
.A(n_93),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_L g132 ( 
.A(n_119),
.B(n_122),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_L g120 ( 
.A(n_87),
.B(n_70),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_L g140 ( 
.A(n_120),
.B(n_121),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_SL g121 ( 
.A(n_95),
.B(n_66),
.Y(n_121)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_90),
.Y(n_122)
);

CKINVDCx16_ASAP7_75t_R g124 ( 
.A(n_104),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_L g139 ( 
.A(n_124),
.B(n_84),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_L g125 ( 
.A(n_101),
.B(n_73),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_L g142 ( 
.A(n_125),
.B(n_105),
.Y(n_142)
);

MAJIxp5_ASAP7_75t_L g127 ( 
.A(n_125),
.B(n_98),
.C(n_86),
.Y(n_127)
);

MAJIxp5_ASAP7_75t_L g151 ( 
.A(n_127),
.B(n_137),
.C(n_145),
.Y(n_151)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_108),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_L g149 ( 
.A(n_128),
.B(n_131),
.Y(n_149)
);

XNOR2xp5_ASAP7_75t_SL g155 ( 
.A(n_130),
.B(n_107),
.Y(n_155)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_108),
.Y(n_131)
);

OAI22xp5_ASAP7_75t_SL g150 ( 
.A1(n_134),
.A2(n_146),
.B1(n_126),
.B2(n_124),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_SL g136 ( 
.A(n_111),
.B(n_105),
.Y(n_136)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_136),
.Y(n_147)
);

XOR2xp5_ASAP7_75t_L g137 ( 
.A(n_109),
.B(n_105),
.Y(n_137)
);

AOI22xp5_ASAP7_75t_L g162 ( 
.A1(n_139),
.A2(n_106),
.B1(n_115),
.B2(n_118),
.Y(n_162)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_120),
.Y(n_141)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_141),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_L g154 ( 
.A(n_142),
.B(n_110),
.Y(n_154)
);

NOR2xp33_ASAP7_75t_L g143 ( 
.A(n_116),
.B(n_96),
.Y(n_143)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_143),
.Y(n_152)
);

AND2x2_ASAP7_75t_L g144 ( 
.A(n_115),
.B(n_85),
.Y(n_144)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_144),
.Y(n_153)
);

MAJIxp5_ASAP7_75t_L g145 ( 
.A(n_109),
.B(n_69),
.C(n_91),
.Y(n_145)
);

AOI22xp5_ASAP7_75t_L g146 ( 
.A1(n_122),
.A2(n_78),
.B1(n_64),
.B2(n_91),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_L g175 ( 
.A(n_150),
.B(n_164),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_L g179 ( 
.A(n_154),
.B(n_156),
.Y(n_179)
);

XNOR2xp5_ASAP7_75t_L g170 ( 
.A(n_155),
.B(n_130),
.Y(n_170)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_140),
.Y(n_156)
);

MAJIxp5_ASAP7_75t_L g157 ( 
.A(n_127),
.B(n_119),
.C(n_112),
.Y(n_157)
);

MAJIxp5_ASAP7_75t_L g169 ( 
.A(n_157),
.B(n_159),
.C(n_137),
.Y(n_169)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_135),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_SL g167 ( 
.A(n_158),
.B(n_161),
.Y(n_167)
);

MAJIxp5_ASAP7_75t_L g159 ( 
.A(n_142),
.B(n_112),
.C(n_107),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_L g160 ( 
.A(n_140),
.B(n_114),
.Y(n_160)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_160),
.Y(n_165)
);

INVxp67_ASAP7_75t_L g161 ( 
.A(n_146),
.Y(n_161)
);

OAI21xp5_ASAP7_75t_L g172 ( 
.A1(n_162),
.A2(n_153),
.B(n_129),
.Y(n_172)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_132),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_SL g176 ( 
.A(n_163),
.B(n_145),
.Y(n_176)
);

OAI321xp33_ASAP7_75t_L g164 ( 
.A1(n_138),
.A2(n_123),
.A3(n_106),
.B1(n_113),
.B2(n_121),
.C(n_117),
.Y(n_164)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_149),
.Y(n_166)
);

NOR2xp33_ASAP7_75t_L g187 ( 
.A(n_166),
.B(n_168),
.Y(n_187)
);

HB1xp67_ASAP7_75t_L g168 ( 
.A(n_161),
.Y(n_168)
);

MAJIxp5_ASAP7_75t_L g189 ( 
.A(n_169),
.B(n_177),
.C(n_151),
.Y(n_189)
);

XOR2xp5_ASAP7_75t_L g182 ( 
.A(n_170),
.B(n_155),
.Y(n_182)
);

CKINVDCx16_ASAP7_75t_R g171 ( 
.A(n_150),
.Y(n_171)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_171),
.Y(n_186)
);

OAI21xp5_ASAP7_75t_SL g181 ( 
.A1(n_172),
.A2(n_174),
.B(n_162),
.Y(n_181)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_160),
.Y(n_173)
);

NOR2xp33_ASAP7_75t_L g188 ( 
.A(n_173),
.B(n_178),
.Y(n_188)
);

AOI22xp5_ASAP7_75t_SL g174 ( 
.A1(n_153),
.A2(n_129),
.B1(n_134),
.B2(n_144),
.Y(n_174)
);

NOR2xp33_ASAP7_75t_SL g183 ( 
.A(n_176),
.B(n_147),
.Y(n_183)
);

XNOR2xp5_ASAP7_75t_L g177 ( 
.A(n_151),
.B(n_133),
.Y(n_177)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_152),
.Y(n_178)
);

AOI21xp5_ASAP7_75t_SL g180 ( 
.A1(n_172),
.A2(n_144),
.B(n_156),
.Y(n_180)
);

OAI31xp33_ASAP7_75t_L g194 ( 
.A1(n_180),
.A2(n_179),
.A3(n_165),
.B(n_170),
.Y(n_194)
);

XNOR2xp5_ASAP7_75t_SL g199 ( 
.A(n_181),
.B(n_1),
.Y(n_199)
);

XOR2xp5_ASAP7_75t_L g197 ( 
.A(n_182),
.B(n_169),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_L g201 ( 
.A(n_183),
.B(n_184),
.Y(n_201)
);

NOR2xp33_ASAP7_75t_SL g184 ( 
.A(n_175),
.B(n_138),
.Y(n_184)
);

AOI21xp5_ASAP7_75t_L g185 ( 
.A1(n_174),
.A2(n_159),
.B(n_148),
.Y(n_185)
);

NOR2xp33_ASAP7_75t_L g195 ( 
.A(n_185),
.B(n_191),
.Y(n_195)
);

XOR2xp5_ASAP7_75t_L g198 ( 
.A(n_189),
.B(n_182),
.Y(n_198)
);

AOI22xp5_ASAP7_75t_L g190 ( 
.A1(n_167),
.A2(n_157),
.B1(n_154),
.B2(n_64),
.Y(n_190)
);

CKINVDCx16_ASAP7_75t_R g193 ( 
.A(n_190),
.Y(n_193)
);

AOI21xp5_ASAP7_75t_L g191 ( 
.A1(n_179),
.A2(n_15),
.B(n_3),
.Y(n_191)
);

XNOR2xp5_ASAP7_75t_L g192 ( 
.A(n_189),
.B(n_177),
.Y(n_192)
);

XNOR2xp5_ASAP7_75t_L g205 ( 
.A(n_192),
.B(n_196),
.Y(n_205)
);

OAI21xp33_ASAP7_75t_SL g207 ( 
.A1(n_194),
.A2(n_199),
.B(n_200),
.Y(n_207)
);

NOR2xp33_ASAP7_75t_L g196 ( 
.A(n_191),
.B(n_187),
.Y(n_196)
);

XOR2xp5_ASAP7_75t_L g206 ( 
.A(n_197),
.B(n_198),
.Y(n_206)
);

XOR2xp5_ASAP7_75t_L g200 ( 
.A(n_181),
.B(n_1),
.Y(n_200)
);

OAI21xp5_ASAP7_75t_SL g202 ( 
.A1(n_193),
.A2(n_185),
.B(n_180),
.Y(n_202)
);

AOI21xp5_ASAP7_75t_SL g212 ( 
.A1(n_202),
.A2(n_207),
.B(n_206),
.Y(n_212)
);

AOI22xp5_ASAP7_75t_L g203 ( 
.A1(n_195),
.A2(n_186),
.B1(n_188),
.B2(n_190),
.Y(n_203)
);

OAI22xp5_ASAP7_75t_SL g209 ( 
.A1(n_203),
.A2(n_200),
.B1(n_197),
.B2(n_8),
.Y(n_209)
);

AOI31xp67_ASAP7_75t_SL g204 ( 
.A1(n_201),
.A2(n_4),
.A3(n_6),
.B(n_8),
.Y(n_204)
);

OAI21x1_ASAP7_75t_L g210 ( 
.A1(n_204),
.A2(n_208),
.B(n_4),
.Y(n_210)
);

AOI21x1_ASAP7_75t_L g208 ( 
.A1(n_199),
.A2(n_4),
.B(n_6),
.Y(n_208)
);

NOR2xp33_ASAP7_75t_L g215 ( 
.A(n_209),
.B(n_210),
.Y(n_215)
);

NAND2xp5_ASAP7_75t_L g211 ( 
.A(n_205),
.B(n_6),
.Y(n_211)
);

NOR2xp33_ASAP7_75t_L g217 ( 
.A(n_211),
.B(n_212),
.Y(n_217)
);

AND2x2_ASAP7_75t_L g213 ( 
.A(n_206),
.B(n_207),
.Y(n_213)
);

MAJx2_ASAP7_75t_L g216 ( 
.A(n_213),
.B(n_9),
.C(n_10),
.Y(n_216)
);

OAI21xp5_ASAP7_75t_L g214 ( 
.A1(n_203),
.A2(n_9),
.B(n_10),
.Y(n_214)
);

MAJIxp5_ASAP7_75t_L g218 ( 
.A(n_214),
.B(n_10),
.C(n_11),
.Y(n_218)
);

AOI31xp33_ASAP7_75t_L g221 ( 
.A1(n_216),
.A2(n_12),
.A3(n_13),
.B(n_14),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_L g220 ( 
.A(n_218),
.B(n_11),
.Y(n_220)
);

XNOR2xp5_ASAP7_75t_L g219 ( 
.A(n_217),
.B(n_11),
.Y(n_219)
);

NAND2xp5_ASAP7_75t_SL g223 ( 
.A(n_219),
.B(n_220),
.Y(n_223)
);

OAI21xp5_ASAP7_75t_L g222 ( 
.A1(n_221),
.A2(n_215),
.B(n_13),
.Y(n_222)
);

AOI22xp5_ASAP7_75t_L g224 ( 
.A1(n_222),
.A2(n_12),
.B1(n_13),
.B2(n_14),
.Y(n_224)
);

XNOR2xp5_ASAP7_75t_L g225 ( 
.A(n_224),
.B(n_223),
.Y(n_225)
);


endmodule