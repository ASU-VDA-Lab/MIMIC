module fake_jpeg_12300_n_183 (n_13, n_21, n_33, n_1, n_45, n_10, n_23, n_27, n_6, n_22, n_47, n_14, n_40, n_19, n_18, n_20, n_35, n_48, n_46, n_41, n_4, n_34, n_30, n_39, n_42, n_16, n_49, n_3, n_0, n_24, n_28, n_38, n_26, n_44, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_43, n_50, n_12, n_32, n_8, n_15, n_7, n_183);

input n_13;
input n_21;
input n_33;
input n_1;
input n_45;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_47;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_48;
input n_46;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_42;
input n_16;
input n_49;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_44;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_43;
input n_50;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_183;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_64;
wire n_55;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_84;
wire n_59;
wire n_98;
wire n_178;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_76;
wire n_154;
wire n_127;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_155;
wire n_103;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_175;
wire n_57;
wire n_171;
wire n_119;
wire n_69;
wire n_83;
wire n_179;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_168;
wire n_106;
wire n_111;
wire n_143;
wire n_122;
wire n_75;
wire n_102;
wire n_121;
wire n_99;
wire n_130;
wire n_70;
wire n_177;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_128;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_91;
wire n_54;
wire n_93;
wire n_161;
wire n_138;
wire n_101;
wire n_149;
wire n_157;
wire n_87;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_176;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_62;
wire n_167;
wire n_174;
wire n_120;
wire n_100;
wire n_118;
wire n_82;
wire n_140;
wire n_96;

INVx1_ASAP7_75t_L g51 ( 
.A(n_50),
.Y(n_51)
);

INVx3_ASAP7_75t_L g52 ( 
.A(n_45),
.Y(n_52)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_5),
.Y(n_53)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_30),
.Y(n_54)
);

INVx4_ASAP7_75t_L g55 ( 
.A(n_18),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_17),
.Y(n_56)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_4),
.Y(n_57)
);

INVx13_ASAP7_75t_L g58 ( 
.A(n_0),
.Y(n_58)
);

BUFx12f_ASAP7_75t_L g59 ( 
.A(n_32),
.Y(n_59)
);

CKINVDCx20_ASAP7_75t_R g60 ( 
.A(n_9),
.Y(n_60)
);

BUFx5_ASAP7_75t_L g61 ( 
.A(n_16),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_34),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_8),
.Y(n_63)
);

CKINVDCx20_ASAP7_75t_R g64 ( 
.A(n_20),
.Y(n_64)
);

BUFx12f_ASAP7_75t_L g65 ( 
.A(n_29),
.Y(n_65)
);

CKINVDCx20_ASAP7_75t_R g66 ( 
.A(n_47),
.Y(n_66)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_27),
.Y(n_67)
);

BUFx16f_ASAP7_75t_L g68 ( 
.A(n_49),
.Y(n_68)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_19),
.Y(n_69)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_35),
.Y(n_70)
);

BUFx16f_ASAP7_75t_L g71 ( 
.A(n_5),
.Y(n_71)
);

CKINVDCx20_ASAP7_75t_R g72 ( 
.A(n_37),
.Y(n_72)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_4),
.Y(n_73)
);

BUFx6f_ASAP7_75t_L g74 ( 
.A(n_41),
.Y(n_74)
);

CKINVDCx20_ASAP7_75t_R g75 ( 
.A(n_13),
.Y(n_75)
);

CKINVDCx20_ASAP7_75t_R g76 ( 
.A(n_42),
.Y(n_76)
);

BUFx2_ASAP7_75t_L g77 ( 
.A(n_7),
.Y(n_77)
);

BUFx2_ASAP7_75t_L g78 ( 
.A(n_28),
.Y(n_78)
);

INVx2_ASAP7_75t_L g79 ( 
.A(n_77),
.Y(n_79)
);

INVx2_ASAP7_75t_L g89 ( 
.A(n_79),
.Y(n_89)
);

BUFx6f_ASAP7_75t_L g80 ( 
.A(n_56),
.Y(n_80)
);

BUFx6f_ASAP7_75t_L g91 ( 
.A(n_80),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_53),
.B(n_0),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_SL g97 ( 
.A(n_81),
.B(n_72),
.Y(n_97)
);

BUFx6f_ASAP7_75t_L g82 ( 
.A(n_56),
.Y(n_82)
);

BUFx3_ASAP7_75t_L g99 ( 
.A(n_82),
.Y(n_99)
);

BUFx6f_ASAP7_75t_L g83 ( 
.A(n_62),
.Y(n_83)
);

BUFx12f_ASAP7_75t_L g92 ( 
.A(n_83),
.Y(n_92)
);

OAI22xp5_ASAP7_75t_SL g84 ( 
.A1(n_63),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_84)
);

AOI22xp33_ASAP7_75t_SL g96 ( 
.A1(n_84),
.A2(n_59),
.B1(n_65),
.B2(n_78),
.Y(n_96)
);

INVx2_ASAP7_75t_L g85 ( 
.A(n_77),
.Y(n_85)
);

INVx2_ASAP7_75t_L g100 ( 
.A(n_85),
.Y(n_100)
);

INVx6_ASAP7_75t_L g86 ( 
.A(n_62),
.Y(n_86)
);

INVx4_ASAP7_75t_L g103 ( 
.A(n_86),
.Y(n_103)
);

CKINVDCx20_ASAP7_75t_R g87 ( 
.A(n_64),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_87),
.B(n_66),
.Y(n_95)
);

BUFx6f_ASAP7_75t_L g88 ( 
.A(n_74),
.Y(n_88)
);

INVx5_ASAP7_75t_L g93 ( 
.A(n_88),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_L g90 ( 
.A(n_86),
.B(n_60),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_L g119 ( 
.A(n_90),
.B(n_94),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_L g94 ( 
.A(n_80),
.B(n_73),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g112 ( 
.A(n_95),
.B(n_96),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_L g122 ( 
.A(n_97),
.B(n_98),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_SL g98 ( 
.A(n_82),
.B(n_57),
.Y(n_98)
);

INVx5_ASAP7_75t_SL g101 ( 
.A(n_83),
.Y(n_101)
);

INVx4_ASAP7_75t_SL g107 ( 
.A(n_101),
.Y(n_107)
);

FAx1_ASAP7_75t_SL g102 ( 
.A(n_88),
.B(n_58),
.CI(n_2),
.CON(n_102),
.SN(n_102)
);

OR2x2_ASAP7_75t_L g115 ( 
.A(n_102),
.B(n_61),
.Y(n_115)
);

INVx13_ASAP7_75t_L g104 ( 
.A(n_101),
.Y(n_104)
);

NOR3xp33_ASAP7_75t_L g129 ( 
.A(n_104),
.B(n_109),
.C(n_111),
.Y(n_129)
);

OAI22xp33_ASAP7_75t_SL g105 ( 
.A1(n_96),
.A2(n_78),
.B1(n_63),
.B2(n_74),
.Y(n_105)
);

OAI22xp5_ASAP7_75t_SL g131 ( 
.A1(n_105),
.A2(n_108),
.B1(n_120),
.B2(n_65),
.Y(n_131)
);

INVx2_ASAP7_75t_L g106 ( 
.A(n_89),
.Y(n_106)
);

INVx3_ASAP7_75t_L g127 ( 
.A(n_106),
.Y(n_127)
);

AOI22xp5_ASAP7_75t_L g108 ( 
.A1(n_102),
.A2(n_55),
.B1(n_52),
.B2(n_54),
.Y(n_108)
);

AOI22xp5_ASAP7_75t_SL g109 ( 
.A1(n_100),
.A2(n_59),
.B1(n_65),
.B2(n_58),
.Y(n_109)
);

INVx8_ASAP7_75t_L g110 ( 
.A(n_91),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_SL g128 ( 
.A(n_110),
.B(n_115),
.Y(n_128)
);

AND2x6_ASAP7_75t_L g111 ( 
.A(n_103),
.B(n_38),
.Y(n_111)
);

MAJIxp5_ASAP7_75t_L g113 ( 
.A(n_91),
.B(n_69),
.C(n_67),
.Y(n_113)
);

MAJIxp5_ASAP7_75t_L g136 ( 
.A(n_113),
.B(n_71),
.C(n_68),
.Y(n_136)
);

INVxp67_ASAP7_75t_L g114 ( 
.A(n_92),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_L g133 ( 
.A(n_114),
.B(n_116),
.Y(n_133)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_103),
.Y(n_116)
);

INVx8_ASAP7_75t_L g117 ( 
.A(n_92),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_SL g132 ( 
.A(n_117),
.B(n_68),
.Y(n_132)
);

CKINVDCx20_ASAP7_75t_R g118 ( 
.A(n_93),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_L g135 ( 
.A(n_118),
.B(n_121),
.Y(n_135)
);

AOI22xp5_ASAP7_75t_L g120 ( 
.A1(n_99),
.A2(n_70),
.B1(n_51),
.B2(n_76),
.Y(n_120)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_92),
.Y(n_121)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_99),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_L g137 ( 
.A(n_123),
.B(n_124),
.Y(n_137)
);

INVxp67_ASAP7_75t_L g124 ( 
.A(n_98),
.Y(n_124)
);

INVx13_ASAP7_75t_L g125 ( 
.A(n_101),
.Y(n_125)
);

CKINVDCx20_ASAP7_75t_R g134 ( 
.A(n_125),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_SL g126 ( 
.A(n_122),
.B(n_75),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_L g156 ( 
.A(n_126),
.B(n_136),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_L g130 ( 
.A(n_119),
.B(n_59),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_L g159 ( 
.A(n_130),
.B(n_131),
.Y(n_159)
);

CKINVDCx14_ASAP7_75t_R g157 ( 
.A(n_132),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_L g138 ( 
.A(n_115),
.B(n_25),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_L g160 ( 
.A(n_138),
.B(n_140),
.Y(n_160)
);

NOR2xp33_ASAP7_75t_SL g139 ( 
.A(n_112),
.B(n_1),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_L g164 ( 
.A(n_139),
.B(n_141),
.Y(n_164)
);

NOR2xp33_ASAP7_75t_L g140 ( 
.A(n_117),
.B(n_71),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_L g141 ( 
.A(n_110),
.B(n_3),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_L g142 ( 
.A(n_111),
.B(n_6),
.Y(n_142)
);

XOR2xp5_ASAP7_75t_L g155 ( 
.A(n_142),
.B(n_145),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_SL g143 ( 
.A(n_107),
.B(n_6),
.Y(n_143)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_143),
.Y(n_149)
);

NOR2xp33_ASAP7_75t_SL g144 ( 
.A(n_107),
.B(n_7),
.Y(n_144)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_144),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_L g145 ( 
.A(n_104),
.B(n_8),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_L g146 ( 
.A(n_105),
.B(n_48),
.Y(n_146)
);

XNOR2xp5_ASAP7_75t_SL g153 ( 
.A(n_146),
.B(n_10),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_L g147 ( 
.A(n_125),
.B(n_9),
.Y(n_147)
);

OAI21xp5_ASAP7_75t_SL g151 ( 
.A1(n_147),
.A2(n_148),
.B(n_31),
.Y(n_151)
);

NOR2xp33_ASAP7_75t_L g148 ( 
.A(n_122),
.B(n_10),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_L g171 ( 
.A(n_151),
.B(n_152),
.Y(n_171)
);

OAI22x1_ASAP7_75t_L g152 ( 
.A1(n_128),
.A2(n_33),
.B1(n_46),
.B2(n_44),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_L g167 ( 
.A(n_153),
.B(n_161),
.Y(n_167)
);

OAI21xp5_ASAP7_75t_SL g154 ( 
.A1(n_138),
.A2(n_11),
.B(n_12),
.Y(n_154)
);

OAI21xp5_ASAP7_75t_L g168 ( 
.A1(n_154),
.A2(n_158),
.B(n_162),
.Y(n_168)
);

AOI21xp5_ASAP7_75t_L g158 ( 
.A1(n_135),
.A2(n_11),
.B(n_12),
.Y(n_158)
);

XNOR2xp5_ASAP7_75t_SL g161 ( 
.A(n_130),
.B(n_14),
.Y(n_161)
);

INVx2_ASAP7_75t_L g162 ( 
.A(n_127),
.Y(n_162)
);

OAI22xp5_ASAP7_75t_SL g163 ( 
.A1(n_146),
.A2(n_15),
.B1(n_21),
.B2(n_22),
.Y(n_163)
);

OAI22xp5_ASAP7_75t_L g166 ( 
.A1(n_163),
.A2(n_136),
.B1(n_134),
.B2(n_133),
.Y(n_166)
);

NOR3xp33_ASAP7_75t_SL g165 ( 
.A(n_160),
.B(n_129),
.C(n_137),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_SL g175 ( 
.A(n_165),
.B(n_166),
.Y(n_175)
);

OAI21xp5_ASAP7_75t_L g169 ( 
.A1(n_159),
.A2(n_131),
.B(n_127),
.Y(n_169)
);

AOI21xp5_ASAP7_75t_SL g174 ( 
.A1(n_169),
.A2(n_155),
.B(n_152),
.Y(n_174)
);

OAI22xp5_ASAP7_75t_L g170 ( 
.A1(n_153),
.A2(n_23),
.B1(n_24),
.B2(n_26),
.Y(n_170)
);

OAI22xp5_ASAP7_75t_SL g173 ( 
.A1(n_170),
.A2(n_164),
.B1(n_150),
.B2(n_149),
.Y(n_173)
);

MAJIxp5_ASAP7_75t_L g172 ( 
.A(n_167),
.B(n_161),
.C(n_156),
.Y(n_172)
);

MAJIxp5_ASAP7_75t_L g177 ( 
.A(n_172),
.B(n_168),
.C(n_167),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_SL g176 ( 
.A(n_173),
.B(n_174),
.Y(n_176)
);

MAJIxp5_ASAP7_75t_L g178 ( 
.A(n_177),
.B(n_175),
.C(n_171),
.Y(n_178)
);

OAI21xp5_ASAP7_75t_L g179 ( 
.A1(n_178),
.A2(n_176),
.B(n_157),
.Y(n_179)
);

XNOR2xp5_ASAP7_75t_L g180 ( 
.A(n_179),
.B(n_157),
.Y(n_180)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_180),
.Y(n_181)
);

O2A1O1Ixp33_ASAP7_75t_L g182 ( 
.A1(n_181),
.A2(n_36),
.B(n_39),
.C(n_40),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_L g183 ( 
.A(n_182),
.B(n_43),
.Y(n_183)
);


endmodule