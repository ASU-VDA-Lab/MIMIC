module real_aes_7347_n_100 (n_17, n_28, n_76, n_56, n_34, n_98, n_90, n_82, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_83, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_91, n_43, n_96, n_54, n_35, n_42, n_99, n_15, n_9, n_23, n_72, n_95, n_44, n_7, n_4, n_80, n_6, n_12, n_68, n_79, n_69, n_46, n_59, n_25, n_73, n_77, n_81, n_48, n_37, n_97, n_70, n_50, n_89, n_26, n_86, n_93, n_13, n_24, n_2, n_55, n_62, n_84, n_67, n_92, n_33, n_88, n_14, n_11, n_85, n_16, n_94, n_39, n_5, n_45, n_60, n_38, n_87, n_0, n_78, n_63, n_1, n_53, n_36, n_100);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_98;
input n_90;
input n_82;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_83;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_91;
input n_43;
input n_96;
input n_54;
input n_35;
input n_42;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_95;
input n_44;
input n_7;
input n_4;
input n_80;
input n_6;
input n_12;
input n_68;
input n_79;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_81;
input n_48;
input n_37;
input n_97;
input n_70;
input n_50;
input n_89;
input n_26;
input n_86;
input n_93;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_84;
input n_67;
input n_92;
input n_33;
input n_88;
input n_14;
input n_11;
input n_85;
input n_16;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_87;
input n_0;
input n_78;
input n_63;
input n_1;
input n_53;
input n_36;
output n_100;
wire n_480;
wire n_113;
wire n_476;
wire n_599;
wire n_187;
wire n_436;
wire n_684;
wire n_257;
wire n_390;
wire n_185;
wire n_285;
wire n_624;
wire n_618;
wire n_522;
wire n_485;
wire n_222;
wire n_750;
wire n_631;
wire n_287;
wire n_357;
wire n_503;
wire n_635;
wire n_386;
wire n_673;
wire n_518;
wire n_254;
wire n_207;
wire n_665;
wire n_667;
wire n_580;
wire n_577;
wire n_469;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_718;
wire n_318;
wire n_355;
wire n_239;
wire n_669;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_742;
wire n_112;
wire n_364;
wire n_319;
wire n_555;
wire n_421;
wire n_329;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_169;
wire n_242;
wire n_376;
wire n_549;
wire n_571;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_448;
wire n_556;
wire n_341;
wire n_545;
wire n_593;
wire n_232;
wire n_460;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_537;
wire n_551;
wire n_320;
wire n_666;
wire n_560;
wire n_260;
wire n_660;
wire n_594;
wire n_186;
wire n_138;
wire n_696;
wire n_704;
wire n_453;
wire n_374;
wire n_379;
wire n_647;
wire n_235;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_161;
wire n_189;
wire n_271;
wire n_489;
wire n_548;
wire n_427;
wire n_678;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_519;
wire n_564;
wire n_638;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_512;
wire n_395;
wire n_332;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_116;
wire n_625;
wire n_462;
wire n_289;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_716;
wire n_213;
wire n_356;
wire n_478;
wire n_584;
wire n_408;
wire n_553;
wire n_184;
wire n_372;
wire n_528;
wire n_578;
wire n_202;
wire n_495;
wire n_370;
wire n_384;
wire n_744;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_467;
wire n_327;
wire n_106;
wire n_559;
wire n_466;
wire n_636;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_726;
wire n_517;
wire n_683;
wire n_174;
wire n_570;
wire n_675;
wire n_530;
wire n_104;
wire n_535;
wire n_732;
wire n_211;
wire n_281;
wire n_496;
wire n_693;
wire n_173;
wire n_468;
wire n_234;
wire n_746;
wire n_284;
wire n_153;
wire n_532;
wire n_316;
wire n_656;
wire n_178;
wire n_409;
wire n_748;
wire n_298;
wire n_523;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_297;
wire n_383;
wire n_529;
wire n_455;
wire n_119;
wire n_504;
wire n_310;
wire n_725;
wire n_164;
wire n_671;
wire n_231;
wire n_102;
wire n_547;
wire n_659;
wire n_634;
wire n_682;
wire n_454;
wire n_122;
wire n_443;
wire n_565;
wire n_608;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_267;
wire n_218;
wire n_737;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_722;
wire n_745;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_331;
wire n_449;
wire n_182;
wire n_363;
wire n_417;
wire n_607;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_561;
wire n_142;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_655;
wire n_654;
wire n_505;
wire n_434;
wire n_502;
wire n_527;
wire n_600;
wire n_731;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_602;
wire n_552;
wire n_402;
wire n_617;
wire n_733;
wire n_171;
wire n_676;
wire n_658;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_432;
wire n_146;
wire n_226;
wire n_255;
wire n_286;
wire n_416;
wire n_410;
wire n_120;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_695;
wire n_685;
wire n_165;
wire n_361;
wire n_632;
wire n_246;
wire n_176;
wire n_412;
wire n_163;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_501;
wire n_488;
wire n_251;
wire n_642;
wire n_613;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_702;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_734;
wire n_110;
wire n_392;
wire n_562;
wire n_150;
wire n_147;
wire n_404;
wire n_288;
wire n_713;
wire n_598;
wire n_735;
wire n_728;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_569;
wire n_563;
wire n_188;
wire n_269;
wire n_430;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_193;
wire n_397;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_649;
wire n_663;
wire n_749;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_707;
wire n_622;
wire n_470;
wire n_133;
wire n_494;
wire n_711;
wire n_377;
wire n_273;
wire n_723;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_265;
wire n_354;
wire n_720;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_730;
wire n_643;
wire n_747;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_148;
wire n_498;
wire n_481;
wire n_691;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_487;
wire n_233;
wire n_290;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_155;
wire n_243;
wire n_692;
wire n_544;
wire n_268;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_101;
wire n_738;
wire n_701;
wire n_309;
wire n_344;
wire n_107;
wire n_229;
wire n_482;
wire n_520;
wire n_633;
wire n_679;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_262;
wire n_630;
wire n_689;
wire n_715;
wire n_134;
wire n_349;
wire n_336;
wire n_420;
wire n_612;
wire n_195;
wire n_438;
wire n_300;
wire n_252;
wire n_283;
wire n_314;
wire n_741;
wire n_249;
wire n_623;
wire n_446;
wire n_721;
wire n_221;
wire n_681;
wire n_156;
wire n_359;
wire n_456;
wire n_717;
wire n_312;
wire n_266;
wire n_183;
wire n_712;
wire n_205;
wire n_433;
wire n_335;
wire n_177;
wire n_516;
wire n_313;
wire n_627;
wire n_739;
wire n_140;
wire n_521;
wire n_418;
wire n_422;
wire n_219;
wire n_524;
wire n_705;
wire n_180;
wire n_212;
wire n_210;
wire n_575;
wire n_325;
wire n_338;
wire n_479;
wire n_442;
wire n_740;
wire n_371;
wire n_698;
wire n_103;
wire n_166;
wire n_541;
wire n_224;
wire n_151;
wire n_546;
wire n_639;
wire n_587;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_724;
wire n_440;
wire n_525;
wire n_674;
wire n_644;
wire n_152;
wire n_198;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_414;
wire n_123;
wire n_279;
wire n_686;
wire n_543;
wire n_497;
wire n_514;
wire n_270;
wire n_507;
wire n_614;
wire n_305;
wire n_586;
wire n_450;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_473;
wire n_465;
wire n_719;
wire n_566;
wire n_474;
wire n_170;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_168;
wire n_241;
wire n_175;
wire n_687;
wire n_729;
wire n_646;
wire n_650;
wire n_710;
wire n_743;
wire n_105;
wire n_294;
wire n_393;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_500;
wire n_307;
wire n_601;
wire n_661;
wire n_463;
wire n_396;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_143;
wire n_192;
wire n_475;
wire n_554;
wire n_264;
wire n_237;
wire n_668;
A2O1A1Ixp33_ASAP7_75t_SL g243 ( .A1(n_0), .A2(n_244), .B(n_245), .C(n_248), .Y(n_243) );
NAND2xp5_ASAP7_75t_L g249 ( .A(n_1), .B(n_232), .Y(n_249) );
INVx1_ASAP7_75t_L g439 ( .A(n_2), .Y(n_439) );
NAND2xp5_ASAP7_75t_SL g159 ( .A(n_3), .B(n_160), .Y(n_159) );
A2O1A1Ixp33_ASAP7_75t_L g531 ( .A1(n_4), .A2(n_121), .B(n_124), .C(n_532), .Y(n_531) );
AOI21xp5_ASAP7_75t_L g555 ( .A1(n_5), .A2(n_116), .B(n_556), .Y(n_555) );
AOI21xp5_ASAP7_75t_L g225 ( .A1(n_6), .A2(n_116), .B(n_226), .Y(n_225) );
NAND2xp5_ASAP7_75t_L g562 ( .A(n_7), .B(n_232), .Y(n_562) );
AO21x2_ASAP7_75t_L g187 ( .A1(n_8), .A2(n_151), .B(n_188), .Y(n_187) );
AND2x6_ASAP7_75t_L g121 ( .A(n_9), .B(n_122), .Y(n_121) );
A2O1A1Ixp33_ASAP7_75t_L g204 ( .A1(n_10), .A2(n_121), .B(n_124), .C(n_205), .Y(n_204) );
INVx1_ASAP7_75t_L g500 ( .A(n_11), .Y(n_500) );
NOR2xp33_ASAP7_75t_L g440 ( .A(n_12), .B(n_40), .Y(n_440) );
NAND2xp5_ASAP7_75t_SL g534 ( .A(n_13), .B(n_208), .Y(n_534) );
INVx1_ASAP7_75t_L g142 ( .A(n_14), .Y(n_142) );
NAND2xp5_ASAP7_75t_SL g194 ( .A(n_15), .B(n_160), .Y(n_194) );
A2O1A1Ixp33_ASAP7_75t_L g517 ( .A1(n_16), .A2(n_161), .B(n_518), .C(n_520), .Y(n_517) );
NAND2xp5_ASAP7_75t_L g521 ( .A(n_17), .B(n_232), .Y(n_521) );
NAND2xp5_ASAP7_75t_L g491 ( .A(n_18), .B(n_136), .Y(n_491) );
A2O1A1Ixp33_ASAP7_75t_L g123 ( .A1(n_19), .A2(n_124), .B(n_127), .C(n_135), .Y(n_123) );
A2O1A1Ixp33_ASAP7_75t_L g507 ( .A1(n_20), .A2(n_196), .B(n_247), .C(n_508), .Y(n_507) );
NAND2xp5_ASAP7_75t_SL g551 ( .A(n_21), .B(n_208), .Y(n_551) );
AOI222xp33_ASAP7_75t_L g100 ( .A1(n_22), .A2(n_101), .B1(n_443), .B2(n_450), .C1(n_743), .C2(n_748), .Y(n_100) );
AOI22xp5_ASAP7_75t_L g102 ( .A1(n_22), .A2(n_103), .B1(n_104), .B2(n_432), .Y(n_102) );
CKINVDCx20_ASAP7_75t_R g432 ( .A(n_22), .Y(n_432) );
NAND2xp5_ASAP7_75t_SL g473 ( .A(n_23), .B(n_208), .Y(n_473) );
CKINVDCx16_ASAP7_75t_R g547 ( .A(n_24), .Y(n_547) );
INVx1_ASAP7_75t_L g472 ( .A(n_25), .Y(n_472) );
A2O1A1Ixp33_ASAP7_75t_L g190 ( .A1(n_26), .A2(n_124), .B(n_135), .C(n_191), .Y(n_190) );
BUFx6f_ASAP7_75t_L g120 ( .A(n_27), .Y(n_120) );
CKINVDCx20_ASAP7_75t_R g530 ( .A(n_28), .Y(n_530) );
INVx1_ASAP7_75t_L g488 ( .A(n_29), .Y(n_488) );
NAND2xp5_ASAP7_75t_SL g441 ( .A(n_30), .B(n_442), .Y(n_441) );
AOI21xp5_ASAP7_75t_L g240 ( .A1(n_31), .A2(n_116), .B(n_241), .Y(n_240) );
INVx2_ASAP7_75t_L g119 ( .A(n_32), .Y(n_119) );
A2O1A1Ixp33_ASAP7_75t_L g172 ( .A1(n_33), .A2(n_164), .B(n_173), .C(n_175), .Y(n_172) );
CKINVDCx20_ASAP7_75t_R g537 ( .A(n_34), .Y(n_537) );
A2O1A1Ixp33_ASAP7_75t_L g558 ( .A1(n_35), .A2(n_247), .B(n_559), .C(n_561), .Y(n_558) );
INVxp67_ASAP7_75t_L g489 ( .A(n_36), .Y(n_489) );
NAND2xp5_ASAP7_75t_L g192 ( .A(n_37), .B(n_193), .Y(n_192) );
A2O1A1Ixp33_ASAP7_75t_L g470 ( .A1(n_38), .A2(n_124), .B(n_135), .C(n_471), .Y(n_470) );
CKINVDCx14_ASAP7_75t_R g557 ( .A(n_39), .Y(n_557) );
A2O1A1Ixp33_ASAP7_75t_L g497 ( .A1(n_41), .A2(n_248), .B(n_498), .C(n_499), .Y(n_497) );
NAND2xp5_ASAP7_75t_L g114 ( .A(n_42), .B(n_115), .Y(n_114) );
CKINVDCx20_ASAP7_75t_R g210 ( .A(n_43), .Y(n_210) );
NAND2xp5_ASAP7_75t_L g219 ( .A(n_44), .B(n_160), .Y(n_219) );
NAND2xp5_ASAP7_75t_L g189 ( .A(n_45), .B(n_116), .Y(n_189) );
CKINVDCx20_ASAP7_75t_R g475 ( .A(n_46), .Y(n_475) );
CKINVDCx20_ASAP7_75t_R g485 ( .A(n_47), .Y(n_485) );
A2O1A1Ixp33_ASAP7_75t_L g216 ( .A1(n_48), .A2(n_164), .B(n_173), .C(n_217), .Y(n_216) );
INVx1_ASAP7_75t_L g246 ( .A(n_49), .Y(n_246) );
OAI22xp5_ASAP7_75t_L g104 ( .A1(n_50), .A2(n_105), .B1(n_106), .B2(n_431), .Y(n_104) );
CKINVDCx16_ASAP7_75t_R g105 ( .A(n_50), .Y(n_105) );
INVx1_ASAP7_75t_L g218 ( .A(n_51), .Y(n_218) );
INVx1_ASAP7_75t_L g506 ( .A(n_52), .Y(n_506) );
NAND2xp5_ASAP7_75t_L g215 ( .A(n_53), .B(n_116), .Y(n_215) );
CKINVDCx20_ASAP7_75t_R g144 ( .A(n_54), .Y(n_144) );
CKINVDCx14_ASAP7_75t_R g496 ( .A(n_55), .Y(n_496) );
INVx1_ASAP7_75t_L g122 ( .A(n_56), .Y(n_122) );
NAND2xp5_ASAP7_75t_L g166 ( .A(n_57), .B(n_116), .Y(n_166) );
NAND2xp5_ASAP7_75t_L g231 ( .A(n_58), .B(n_232), .Y(n_231) );
A2O1A1Ixp33_ASAP7_75t_L g228 ( .A1(n_59), .A2(n_134), .B(n_157), .C(n_229), .Y(n_228) );
INVx1_ASAP7_75t_L g141 ( .A(n_60), .Y(n_141) );
OAI22xp5_ASAP7_75t_L g452 ( .A1(n_61), .A2(n_99), .B1(n_453), .B2(n_454), .Y(n_452) );
CKINVDCx20_ASAP7_75t_R g454 ( .A(n_61), .Y(n_454) );
INVx1_ASAP7_75t_SL g560 ( .A(n_62), .Y(n_560) );
CKINVDCx20_ASAP7_75t_R g446 ( .A(n_63), .Y(n_446) );
NAND2xp5_ASAP7_75t_SL g177 ( .A(n_64), .B(n_160), .Y(n_177) );
NAND2xp5_ASAP7_75t_L g510 ( .A(n_65), .B(n_232), .Y(n_510) );
NAND2xp5_ASAP7_75t_L g206 ( .A(n_66), .B(n_161), .Y(n_206) );
INVx1_ASAP7_75t_L g550 ( .A(n_67), .Y(n_550) );
CKINVDCx16_ASAP7_75t_R g242 ( .A(n_68), .Y(n_242) );
NAND2xp5_ASAP7_75t_L g128 ( .A(n_69), .B(n_129), .Y(n_128) );
A2O1A1Ixp33_ASAP7_75t_L g154 ( .A1(n_70), .A2(n_124), .B(n_155), .C(n_164), .Y(n_154) );
CKINVDCx16_ASAP7_75t_R g227 ( .A(n_71), .Y(n_227) );
INVx1_ASAP7_75t_L g449 ( .A(n_72), .Y(n_449) );
AOI21xp5_ASAP7_75t_L g494 ( .A1(n_73), .A2(n_116), .B(n_495), .Y(n_494) );
CKINVDCx20_ASAP7_75t_R g553 ( .A(n_74), .Y(n_553) );
AOI21xp5_ASAP7_75t_L g514 ( .A1(n_75), .A2(n_116), .B(n_515), .Y(n_514) );
AOI222xp33_ASAP7_75t_SL g451 ( .A1(n_76), .A2(n_452), .B1(n_455), .B2(n_735), .C1(n_736), .C2(n_740), .Y(n_451) );
AOI21xp5_ASAP7_75t_L g483 ( .A1(n_77), .A2(n_115), .B(n_484), .Y(n_483) );
CKINVDCx16_ASAP7_75t_R g469 ( .A(n_78), .Y(n_469) );
INVx1_ASAP7_75t_L g516 ( .A(n_79), .Y(n_516) );
NAND2xp5_ASAP7_75t_SL g131 ( .A(n_80), .B(n_132), .Y(n_131) );
CKINVDCx20_ASAP7_75t_R g181 ( .A(n_81), .Y(n_181) );
AOI21xp5_ASAP7_75t_L g504 ( .A1(n_82), .A2(n_116), .B(n_505), .Y(n_504) );
INVx1_ASAP7_75t_L g519 ( .A(n_83), .Y(n_519) );
INVx2_ASAP7_75t_L g139 ( .A(n_84), .Y(n_139) );
INVx1_ASAP7_75t_L g533 ( .A(n_85), .Y(n_533) );
CKINVDCx20_ASAP7_75t_R g168 ( .A(n_86), .Y(n_168) );
NAND2xp5_ASAP7_75t_SL g207 ( .A(n_87), .B(n_208), .Y(n_207) );
OR2x2_ASAP7_75t_L g436 ( .A(n_88), .B(n_437), .Y(n_436) );
OR2x2_ASAP7_75t_L g458 ( .A(n_88), .B(n_438), .Y(n_458) );
INVx2_ASAP7_75t_L g460 ( .A(n_88), .Y(n_460) );
A2O1A1Ixp33_ASAP7_75t_L g548 ( .A1(n_89), .A2(n_124), .B(n_164), .C(n_549), .Y(n_548) );
NAND2xp5_ASAP7_75t_L g171 ( .A(n_90), .B(n_116), .Y(n_171) );
INVx1_ASAP7_75t_L g176 ( .A(n_91), .Y(n_176) );
INVxp67_ASAP7_75t_L g230 ( .A(n_92), .Y(n_230) );
NAND2xp5_ASAP7_75t_L g501 ( .A(n_93), .B(n_151), .Y(n_501) );
INVx1_ASAP7_75t_L g156 ( .A(n_94), .Y(n_156) );
INVx1_ASAP7_75t_L g202 ( .A(n_95), .Y(n_202) );
NAND2xp5_ASAP7_75t_L g448 ( .A(n_96), .B(n_449), .Y(n_448) );
INVx2_ASAP7_75t_L g509 ( .A(n_97), .Y(n_509) );
AND2x2_ASAP7_75t_L g220 ( .A(n_98), .B(n_138), .Y(n_220) );
CKINVDCx20_ASAP7_75t_R g453 ( .A(n_99), .Y(n_453) );
OAI21xp5_ASAP7_75t_SL g101 ( .A1(n_102), .A2(n_433), .B(n_441), .Y(n_101) );
INVxp67_ASAP7_75t_L g103 ( .A(n_104), .Y(n_103) );
OAI22xp5_ASAP7_75t_SL g736 ( .A1(n_106), .A2(n_462), .B1(n_737), .B2(n_738), .Y(n_736) );
INVx1_ASAP7_75t_L g106 ( .A(n_107), .Y(n_106) );
BUFx2_ASAP7_75t_L g431 ( .A(n_107), .Y(n_431) );
AND3x1_ASAP7_75t_L g107 ( .A(n_108), .B(n_335), .C(n_392), .Y(n_107) );
NOR3xp33_ASAP7_75t_L g108 ( .A(n_109), .B(n_280), .C(n_316), .Y(n_108) );
OAI211xp5_ASAP7_75t_L g109 ( .A1(n_110), .A2(n_182), .B(n_234), .C(n_267), .Y(n_109) );
NAND2xp5_ASAP7_75t_L g110 ( .A(n_111), .B(n_146), .Y(n_110) );
HB1xp67_ASAP7_75t_L g111 ( .A(n_112), .Y(n_111) );
AND2x4_ASAP7_75t_L g237 ( .A(n_112), .B(n_238), .Y(n_237) );
INVx5_ASAP7_75t_L g266 ( .A(n_112), .Y(n_266) );
AND2x2_ASAP7_75t_L g339 ( .A(n_112), .B(n_255), .Y(n_339) );
AND2x2_ASAP7_75t_L g377 ( .A(n_112), .B(n_283), .Y(n_377) );
AND2x2_ASAP7_75t_L g397 ( .A(n_112), .B(n_239), .Y(n_397) );
OR2x6_ASAP7_75t_L g112 ( .A(n_113), .B(n_143), .Y(n_112) );
AOI21xp5_ASAP7_75t_SL g113 ( .A1(n_114), .A2(n_123), .B(n_136), .Y(n_113) );
BUFx2_ASAP7_75t_L g115 ( .A(n_116), .Y(n_115) );
AND2x4_ASAP7_75t_L g116 ( .A(n_117), .B(n_121), .Y(n_116) );
NAND2x1p5_ASAP7_75t_L g203 ( .A(n_117), .B(n_121), .Y(n_203) );
AND2x2_ASAP7_75t_L g117 ( .A(n_118), .B(n_120), .Y(n_117) );
INVx1_ASAP7_75t_L g134 ( .A(n_118), .Y(n_134) );
INVx1_ASAP7_75t_L g118 ( .A(n_119), .Y(n_118) );
INVx2_ASAP7_75t_L g125 ( .A(n_119), .Y(n_125) );
INVx1_ASAP7_75t_L g197 ( .A(n_119), .Y(n_197) );
INVx1_ASAP7_75t_L g126 ( .A(n_120), .Y(n_126) );
BUFx6f_ASAP7_75t_L g130 ( .A(n_120), .Y(n_130) );
INVx3_ASAP7_75t_L g161 ( .A(n_120), .Y(n_161) );
INVx1_ASAP7_75t_L g193 ( .A(n_120), .Y(n_193) );
BUFx6f_ASAP7_75t_L g208 ( .A(n_120), .Y(n_208) );
BUFx3_ASAP7_75t_L g135 ( .A(n_121), .Y(n_135) );
INVx4_ASAP7_75t_SL g165 ( .A(n_121), .Y(n_165) );
INVx5_ASAP7_75t_L g174 ( .A(n_124), .Y(n_174) );
AND2x6_ASAP7_75t_L g124 ( .A(n_125), .B(n_126), .Y(n_124) );
BUFx6f_ASAP7_75t_L g163 ( .A(n_125), .Y(n_163) );
BUFx3_ASAP7_75t_L g179 ( .A(n_125), .Y(n_179) );
AOI21xp5_ASAP7_75t_L g127 ( .A1(n_128), .A2(n_131), .B(n_133), .Y(n_127) );
INVx2_ASAP7_75t_L g132 ( .A(n_129), .Y(n_132) );
INVx2_ASAP7_75t_L g129 ( .A(n_130), .Y(n_129) );
INVx4_ASAP7_75t_L g158 ( .A(n_130), .Y(n_158) );
O2A1O1Ixp33_ASAP7_75t_L g175 ( .A1(n_132), .A2(n_176), .B(n_177), .C(n_178), .Y(n_175) );
O2A1O1Ixp33_ASAP7_75t_L g217 ( .A1(n_132), .A2(n_178), .B(n_218), .C(n_219), .Y(n_217) );
O2A1O1Ixp5_ASAP7_75t_L g532 ( .A1(n_132), .A2(n_533), .B(n_534), .C(n_535), .Y(n_532) );
O2A1O1Ixp33_ASAP7_75t_L g549 ( .A1(n_132), .A2(n_535), .B(n_550), .C(n_551), .Y(n_549) );
O2A1O1Ixp33_ASAP7_75t_L g471 ( .A1(n_133), .A2(n_160), .B(n_472), .C(n_473), .Y(n_471) );
INVx2_ASAP7_75t_L g133 ( .A(n_134), .Y(n_133) );
NAND2xp5_ASAP7_75t_SL g486 ( .A(n_134), .B(n_487), .Y(n_486) );
INVx1_ASAP7_75t_L g136 ( .A(n_137), .Y(n_136) );
NOR2xp33_ASAP7_75t_L g552 ( .A(n_137), .B(n_553), .Y(n_552) );
INVx2_ASAP7_75t_L g137 ( .A(n_138), .Y(n_137) );
INVx1_ASAP7_75t_L g145 ( .A(n_138), .Y(n_145) );
AOI21xp5_ASAP7_75t_L g170 ( .A1(n_138), .A2(n_171), .B(n_172), .Y(n_170) );
AOI21xp5_ASAP7_75t_L g214 ( .A1(n_138), .A2(n_215), .B(n_216), .Y(n_214) );
O2A1O1Ixp33_ASAP7_75t_L g468 ( .A1(n_138), .A2(n_203), .B(n_469), .C(n_470), .Y(n_468) );
OA21x2_ASAP7_75t_L g493 ( .A1(n_138), .A2(n_494), .B(n_501), .Y(n_493) );
AND2x2_ASAP7_75t_SL g138 ( .A(n_139), .B(n_140), .Y(n_138) );
AND2x2_ASAP7_75t_L g152 ( .A(n_139), .B(n_140), .Y(n_152) );
NAND2xp5_ASAP7_75t_L g140 ( .A(n_141), .B(n_142), .Y(n_140) );
NOR2xp33_ASAP7_75t_L g143 ( .A(n_144), .B(n_145), .Y(n_143) );
AO21x2_ASAP7_75t_L g528 ( .A1(n_145), .A2(n_529), .B(n_536), .Y(n_528) );
NAND2xp5_ASAP7_75t_L g269 ( .A(n_146), .B(n_270), .Y(n_269) );
AND2x2_ASAP7_75t_L g146 ( .A(n_147), .B(n_169), .Y(n_146) );
HB1xp67_ASAP7_75t_L g278 ( .A(n_147), .Y(n_278) );
AND2x2_ASAP7_75t_L g292 ( .A(n_147), .B(n_238), .Y(n_292) );
INVx1_ASAP7_75t_L g315 ( .A(n_147), .Y(n_315) );
NAND2xp5_ASAP7_75t_L g354 ( .A(n_147), .B(n_266), .Y(n_354) );
OR2x2_ASAP7_75t_L g391 ( .A(n_147), .B(n_236), .Y(n_391) );
INVx2_ASAP7_75t_L g147 ( .A(n_148), .Y(n_147) );
HB1xp67_ASAP7_75t_L g327 ( .A(n_148), .Y(n_327) );
AND2x2_ASAP7_75t_L g334 ( .A(n_148), .B(n_239), .Y(n_334) );
INVx2_ASAP7_75t_L g148 ( .A(n_149), .Y(n_148) );
AND2x2_ASAP7_75t_L g255 ( .A(n_149), .B(n_239), .Y(n_255) );
BUFx2_ASAP7_75t_L g283 ( .A(n_149), .Y(n_283) );
AO21x2_ASAP7_75t_L g149 ( .A1(n_150), .A2(n_153), .B(n_167), .Y(n_149) );
NOR2xp33_ASAP7_75t_L g167 ( .A(n_150), .B(n_168), .Y(n_167) );
NOR2xp33_ASAP7_75t_L g180 ( .A(n_150), .B(n_181), .Y(n_180) );
AO21x2_ASAP7_75t_L g200 ( .A1(n_150), .A2(n_201), .B(n_209), .Y(n_200) );
INVx3_ASAP7_75t_L g232 ( .A(n_150), .Y(n_232) );
NOR2xp33_ASAP7_75t_L g474 ( .A(n_150), .B(n_475), .Y(n_474) );
NOR2xp33_ASAP7_75t_L g536 ( .A(n_150), .B(n_537), .Y(n_536) );
AO21x2_ASAP7_75t_L g545 ( .A1(n_150), .A2(n_546), .B(n_552), .Y(n_545) );
INVx4_ASAP7_75t_L g150 ( .A(n_151), .Y(n_150) );
AOI21xp5_ASAP7_75t_L g188 ( .A1(n_151), .A2(n_189), .B(n_190), .Y(n_188) );
HB1xp67_ASAP7_75t_L g224 ( .A(n_151), .Y(n_224) );
BUFx6f_ASAP7_75t_L g151 ( .A(n_152), .Y(n_151) );
INVx1_ASAP7_75t_L g211 ( .A(n_152), .Y(n_211) );
NAND2xp5_ASAP7_75t_L g153 ( .A(n_154), .B(n_166), .Y(n_153) );
O2A1O1Ixp33_ASAP7_75t_L g155 ( .A1(n_156), .A2(n_157), .B(n_159), .C(n_162), .Y(n_155) );
INVx1_ASAP7_75t_L g157 ( .A(n_158), .Y(n_157) );
OAI22xp33_ASAP7_75t_L g487 ( .A1(n_158), .A2(n_160), .B1(n_488), .B2(n_489), .Y(n_487) );
NOR2xp33_ASAP7_75t_L g508 ( .A(n_158), .B(n_509), .Y(n_508) );
NOR2xp33_ASAP7_75t_L g518 ( .A(n_158), .B(n_519), .Y(n_518) );
NOR2xp33_ASAP7_75t_L g229 ( .A(n_160), .B(n_230), .Y(n_229) );
INVx2_ASAP7_75t_L g244 ( .A(n_160), .Y(n_244) );
INVx5_ASAP7_75t_L g160 ( .A(n_161), .Y(n_160) );
NOR2xp33_ASAP7_75t_L g499 ( .A(n_161), .B(n_500), .Y(n_499) );
HB1xp67_ASAP7_75t_L g162 ( .A(n_163), .Y(n_162) );
INVx3_ASAP7_75t_L g561 ( .A(n_163), .Y(n_561) );
INVx1_ASAP7_75t_L g164 ( .A(n_165), .Y(n_164) );
O2A1O1Ixp33_ASAP7_75t_L g226 ( .A1(n_165), .A2(n_174), .B(n_227), .C(n_228), .Y(n_226) );
O2A1O1Ixp33_ASAP7_75t_SL g241 ( .A1(n_165), .A2(n_174), .B(n_242), .C(n_243), .Y(n_241) );
O2A1O1Ixp33_ASAP7_75t_SL g484 ( .A1(n_165), .A2(n_174), .B(n_485), .C(n_486), .Y(n_484) );
O2A1O1Ixp33_ASAP7_75t_SL g495 ( .A1(n_165), .A2(n_174), .B(n_496), .C(n_497), .Y(n_495) );
O2A1O1Ixp33_ASAP7_75t_SL g505 ( .A1(n_165), .A2(n_174), .B(n_506), .C(n_507), .Y(n_505) );
O2A1O1Ixp33_ASAP7_75t_SL g515 ( .A1(n_165), .A2(n_174), .B(n_516), .C(n_517), .Y(n_515) );
O2A1O1Ixp33_ASAP7_75t_L g556 ( .A1(n_165), .A2(n_174), .B(n_557), .C(n_558), .Y(n_556) );
INVx5_ASAP7_75t_L g236 ( .A(n_169), .Y(n_236) );
BUFx2_ASAP7_75t_L g259 ( .A(n_169), .Y(n_259) );
AND2x2_ASAP7_75t_L g416 ( .A(n_169), .B(n_270), .Y(n_416) );
OR2x6_ASAP7_75t_L g169 ( .A(n_170), .B(n_180), .Y(n_169) );
INVx2_ASAP7_75t_L g173 ( .A(n_174), .Y(n_173) );
HB1xp67_ASAP7_75t_L g178 ( .A(n_179), .Y(n_178) );
INVx2_ASAP7_75t_L g248 ( .A(n_179), .Y(n_248) );
INVx1_ASAP7_75t_L g520 ( .A(n_179), .Y(n_520) );
INVx1_ASAP7_75t_L g182 ( .A(n_183), .Y(n_182) );
NAND2xp33_ASAP7_75t_L g183 ( .A(n_184), .B(n_221), .Y(n_183) );
OAI221xp5_ASAP7_75t_L g316 ( .A1(n_184), .A2(n_317), .B1(n_324), .B2(n_325), .C(n_328), .Y(n_316) );
OR2x2_ASAP7_75t_L g184 ( .A(n_185), .B(n_198), .Y(n_184) );
AND2x2_ASAP7_75t_L g222 ( .A(n_185), .B(n_223), .Y(n_222) );
NAND2xp5_ASAP7_75t_L g310 ( .A(n_185), .B(n_311), .Y(n_310) );
INVx1_ASAP7_75t_SL g185 ( .A(n_186), .Y(n_185) );
AND2x2_ASAP7_75t_L g251 ( .A(n_186), .B(n_199), .Y(n_251) );
NAND2xp5_ASAP7_75t_SL g261 ( .A(n_186), .B(n_200), .Y(n_261) );
OR2x2_ASAP7_75t_L g272 ( .A(n_186), .B(n_223), .Y(n_272) );
AND2x2_ASAP7_75t_L g275 ( .A(n_186), .B(n_263), .Y(n_275) );
AND2x2_ASAP7_75t_L g291 ( .A(n_186), .B(n_212), .Y(n_291) );
OR2x2_ASAP7_75t_L g307 ( .A(n_186), .B(n_200), .Y(n_307) );
NAND2xp5_ASAP7_75t_L g369 ( .A(n_186), .B(n_223), .Y(n_369) );
INVx2_ASAP7_75t_L g186 ( .A(n_187), .Y(n_186) );
NAND2xp5_ASAP7_75t_L g361 ( .A(n_187), .B(n_212), .Y(n_361) );
AND2x2_ASAP7_75t_L g364 ( .A(n_187), .B(n_200), .Y(n_364) );
AOI21xp5_ASAP7_75t_L g191 ( .A1(n_192), .A2(n_194), .B(n_195), .Y(n_191) );
AOI21xp5_ASAP7_75t_L g205 ( .A1(n_195), .A2(n_206), .B(n_207), .Y(n_205) );
INVx2_ASAP7_75t_L g195 ( .A(n_196), .Y(n_195) );
INVx3_ASAP7_75t_L g196 ( .A(n_197), .Y(n_196) );
OR2x2_ASAP7_75t_L g285 ( .A(n_198), .B(n_272), .Y(n_285) );
INVx2_ASAP7_75t_L g311 ( .A(n_198), .Y(n_311) );
OR2x2_ASAP7_75t_L g198 ( .A(n_199), .B(n_212), .Y(n_198) );
AND2x2_ASAP7_75t_L g233 ( .A(n_199), .B(n_213), .Y(n_233) );
NAND2xp5_ASAP7_75t_L g290 ( .A(n_199), .B(n_223), .Y(n_290) );
OR2x2_ASAP7_75t_L g301 ( .A(n_199), .B(n_213), .Y(n_301) );
NAND2xp5_ASAP7_75t_L g360 ( .A(n_199), .B(n_263), .Y(n_360) );
OAI221xp5_ASAP7_75t_L g393 ( .A1(n_199), .A2(n_394), .B1(n_396), .B2(n_398), .C(n_401), .Y(n_393) );
INVx5_ASAP7_75t_SL g199 ( .A(n_200), .Y(n_199) );
NAND2xp5_ASAP7_75t_L g332 ( .A(n_200), .B(n_223), .Y(n_332) );
OAI21xp5_ASAP7_75t_L g201 ( .A1(n_202), .A2(n_203), .B(n_204), .Y(n_201) );
OAI21xp5_ASAP7_75t_L g529 ( .A1(n_203), .A2(n_530), .B(n_531), .Y(n_529) );
OAI21xp5_ASAP7_75t_L g546 ( .A1(n_203), .A2(n_547), .B(n_548), .Y(n_546) );
INVx4_ASAP7_75t_L g247 ( .A(n_208), .Y(n_247) );
INVx2_ASAP7_75t_L g498 ( .A(n_208), .Y(n_498) );
NOR2xp33_ASAP7_75t_L g209 ( .A(n_210), .B(n_211), .Y(n_209) );
INVx2_ASAP7_75t_L g481 ( .A(n_211), .Y(n_481) );
NAND2xp5_ASAP7_75t_L g262 ( .A(n_212), .B(n_263), .Y(n_262) );
NOR2xp33_ASAP7_75t_L g273 ( .A(n_212), .B(n_274), .Y(n_273) );
AND2x2_ASAP7_75t_L g279 ( .A(n_212), .B(n_251), .Y(n_279) );
OR2x2_ASAP7_75t_L g323 ( .A(n_212), .B(n_223), .Y(n_323) );
NAND2xp5_ASAP7_75t_L g342 ( .A(n_212), .B(n_275), .Y(n_342) );
NAND2xp5_ASAP7_75t_L g367 ( .A(n_212), .B(n_368), .Y(n_367) );
AND2x2_ASAP7_75t_L g388 ( .A(n_212), .B(n_389), .Y(n_388) );
INVx5_ASAP7_75t_SL g212 ( .A(n_213), .Y(n_212) );
AND2x2_ASAP7_75t_SL g252 ( .A(n_213), .B(n_222), .Y(n_252) );
O2A1O1Ixp33_ASAP7_75t_SL g256 ( .A1(n_213), .A2(n_257), .B(n_260), .C(n_264), .Y(n_256) );
OR2x2_ASAP7_75t_L g294 ( .A(n_213), .B(n_290), .Y(n_294) );
OR2x2_ASAP7_75t_L g330 ( .A(n_213), .B(n_272), .Y(n_330) );
OAI311xp33_ASAP7_75t_L g336 ( .A1(n_213), .A2(n_275), .A3(n_337), .B1(n_340), .C1(n_347), .Y(n_336) );
AND2x2_ASAP7_75t_L g387 ( .A(n_213), .B(n_223), .Y(n_387) );
AND2x2_ASAP7_75t_L g395 ( .A(n_213), .B(n_250), .Y(n_395) );
HB1xp67_ASAP7_75t_L g413 ( .A(n_213), .Y(n_413) );
AND2x2_ASAP7_75t_L g430 ( .A(n_213), .B(n_251), .Y(n_430) );
OR2x6_ASAP7_75t_L g213 ( .A(n_214), .B(n_220), .Y(n_213) );
NAND2xp5_ASAP7_75t_L g221 ( .A(n_222), .B(n_233), .Y(n_221) );
AND2x2_ASAP7_75t_L g258 ( .A(n_222), .B(n_259), .Y(n_258) );
INVx2_ASAP7_75t_L g414 ( .A(n_222), .Y(n_414) );
AND2x2_ASAP7_75t_L g250 ( .A(n_223), .B(n_251), .Y(n_250) );
INVx3_ASAP7_75t_L g263 ( .A(n_223), .Y(n_263) );
HB1xp67_ASAP7_75t_L g306 ( .A(n_223), .Y(n_306) );
INVxp67_ASAP7_75t_L g345 ( .A(n_223), .Y(n_345) );
OA21x2_ASAP7_75t_L g223 ( .A1(n_224), .A2(n_225), .B(n_231), .Y(n_223) );
OA21x2_ASAP7_75t_L g503 ( .A1(n_224), .A2(n_504), .B(n_510), .Y(n_503) );
OA21x2_ASAP7_75t_L g513 ( .A1(n_224), .A2(n_514), .B(n_521), .Y(n_513) );
OA21x2_ASAP7_75t_L g554 ( .A1(n_224), .A2(n_555), .B(n_562), .Y(n_554) );
OA21x2_ASAP7_75t_L g239 ( .A1(n_232), .A2(n_240), .B(n_249), .Y(n_239) );
AND2x2_ASAP7_75t_L g423 ( .A(n_233), .B(n_271), .Y(n_423) );
AOI221xp5_ASAP7_75t_L g234 ( .A1(n_235), .A2(n_250), .B1(n_252), .B2(n_253), .C(n_256), .Y(n_234) );
AND2x2_ASAP7_75t_L g235 ( .A(n_236), .B(n_237), .Y(n_235) );
NAND2xp5_ASAP7_75t_L g254 ( .A(n_236), .B(n_255), .Y(n_254) );
AND2x2_ASAP7_75t_L g276 ( .A(n_236), .B(n_266), .Y(n_276) );
AND2x2_ASAP7_75t_L g284 ( .A(n_236), .B(n_238), .Y(n_284) );
OR2x2_ASAP7_75t_L g296 ( .A(n_236), .B(n_297), .Y(n_296) );
AND2x2_ASAP7_75t_L g314 ( .A(n_236), .B(n_315), .Y(n_314) );
AND2x2_ASAP7_75t_L g338 ( .A(n_236), .B(n_339), .Y(n_338) );
HB1xp67_ASAP7_75t_L g358 ( .A(n_236), .Y(n_358) );
AND2x2_ASAP7_75t_L g410 ( .A(n_236), .B(n_334), .Y(n_410) );
OAI31xp33_ASAP7_75t_L g418 ( .A1(n_236), .A2(n_287), .A3(n_386), .B(n_419), .Y(n_418) );
NAND2xp5_ASAP7_75t_L g313 ( .A(n_237), .B(n_314), .Y(n_313) );
INVx1_ASAP7_75t_SL g382 ( .A(n_237), .Y(n_382) );
NOR2xp33_ASAP7_75t_L g390 ( .A(n_237), .B(n_391), .Y(n_390) );
AND2x4_ASAP7_75t_L g270 ( .A(n_238), .B(n_266), .Y(n_270) );
INVx1_ASAP7_75t_L g357 ( .A(n_238), .Y(n_357) );
INVx2_ASAP7_75t_L g238 ( .A(n_239), .Y(n_238) );
AND2x2_ASAP7_75t_L g407 ( .A(n_239), .B(n_266), .Y(n_407) );
NOR2xp33_ASAP7_75t_L g245 ( .A(n_246), .B(n_247), .Y(n_245) );
NOR2xp33_ASAP7_75t_L g559 ( .A(n_247), .B(n_560), .Y(n_559) );
INVx2_ASAP7_75t_L g535 ( .A(n_248), .Y(n_535) );
INVx1_ASAP7_75t_SL g417 ( .A(n_250), .Y(n_417) );
NAND2xp5_ASAP7_75t_L g321 ( .A(n_251), .B(n_322), .Y(n_321) );
AOI22xp5_ASAP7_75t_L g401 ( .A1(n_252), .A2(n_364), .B1(n_402), .B2(n_405), .Y(n_401) );
INVx1_ASAP7_75t_L g253 ( .A(n_254), .Y(n_253) );
AND2x2_ASAP7_75t_L g265 ( .A(n_255), .B(n_266), .Y(n_265) );
INVx1_ASAP7_75t_L g324 ( .A(n_255), .Y(n_324) );
NAND2xp5_ASAP7_75t_L g429 ( .A(n_255), .B(n_276), .Y(n_429) );
INVx1_ASAP7_75t_SL g257 ( .A(n_258), .Y(n_257) );
AND2x2_ASAP7_75t_L g399 ( .A(n_258), .B(n_400), .Y(n_399) );
AOI21xp5_ASAP7_75t_L g317 ( .A1(n_259), .A2(n_318), .B(n_320), .Y(n_317) );
OR2x2_ASAP7_75t_L g325 ( .A(n_259), .B(n_326), .Y(n_325) );
AND2x2_ASAP7_75t_L g346 ( .A(n_259), .B(n_334), .Y(n_346) );
NAND2xp5_ASAP7_75t_L g385 ( .A(n_259), .B(n_357), .Y(n_385) );
NAND2xp5_ASAP7_75t_L g396 ( .A(n_259), .B(n_397), .Y(n_396) );
OAI221xp5_ASAP7_75t_SL g373 ( .A1(n_260), .A2(n_374), .B1(n_379), .B2(n_382), .C(n_383), .Y(n_373) );
OR2x2_ASAP7_75t_L g260 ( .A(n_261), .B(n_262), .Y(n_260) );
OR2x2_ASAP7_75t_L g350 ( .A(n_261), .B(n_323), .Y(n_350) );
INVx1_ASAP7_75t_L g389 ( .A(n_261), .Y(n_389) );
INVx2_ASAP7_75t_L g365 ( .A(n_262), .Y(n_365) );
INVx1_ASAP7_75t_L g299 ( .A(n_263), .Y(n_299) );
INVx1_ASAP7_75t_SL g264 ( .A(n_265), .Y(n_264) );
INVx2_ASAP7_75t_L g304 ( .A(n_266), .Y(n_304) );
NAND2xp5_ASAP7_75t_L g326 ( .A(n_266), .B(n_327), .Y(n_326) );
AND2x2_ASAP7_75t_L g333 ( .A(n_266), .B(n_334), .Y(n_333) );
OR2x2_ASAP7_75t_L g421 ( .A(n_266), .B(n_391), .Y(n_421) );
AOI222xp33_ASAP7_75t_L g267 ( .A1(n_268), .A2(n_271), .B1(n_273), .B2(n_276), .C1(n_277), .C2(n_279), .Y(n_267) );
INVxp67_ASAP7_75t_L g268 ( .A(n_269), .Y(n_268) );
AND2x2_ASAP7_75t_L g277 ( .A(n_270), .B(n_278), .Y(n_277) );
AOI22xp33_ASAP7_75t_L g347 ( .A1(n_270), .A2(n_320), .B1(n_348), .B2(n_349), .Y(n_347) );
NAND2xp5_ASAP7_75t_L g403 ( .A(n_270), .B(n_404), .Y(n_403) );
INVx1_ASAP7_75t_SL g271 ( .A(n_272), .Y(n_271) );
INVx1_ASAP7_75t_SL g274 ( .A(n_275), .Y(n_274) );
OAI21xp33_ASAP7_75t_SL g308 ( .A1(n_279), .A2(n_309), .B(n_312), .Y(n_308) );
OAI211xp5_ASAP7_75t_SL g280 ( .A1(n_281), .A2(n_285), .B(n_286), .C(n_308), .Y(n_280) );
INVxp67_ASAP7_75t_L g281 ( .A(n_282), .Y(n_281) );
AND2x2_ASAP7_75t_L g282 ( .A(n_283), .B(n_284), .Y(n_282) );
AOI221xp5_ASAP7_75t_L g286 ( .A1(n_284), .A2(n_287), .B1(n_292), .B2(n_293), .C(n_295), .Y(n_286) );
NAND2xp5_ASAP7_75t_L g371 ( .A(n_284), .B(n_372), .Y(n_371) );
INVxp67_ASAP7_75t_L g378 ( .A(n_284), .Y(n_378) );
INVx1_ASAP7_75t_L g287 ( .A(n_288), .Y(n_287) );
NAND2xp5_ASAP7_75t_L g288 ( .A(n_289), .B(n_291), .Y(n_288) );
AND2x2_ASAP7_75t_L g380 ( .A(n_289), .B(n_381), .Y(n_380) );
INVx1_ASAP7_75t_SL g289 ( .A(n_290), .Y(n_289) );
INVx1_ASAP7_75t_L g297 ( .A(n_292), .Y(n_297) );
AND2x2_ASAP7_75t_L g303 ( .A(n_292), .B(n_304), .Y(n_303) );
INVx1_ASAP7_75t_L g293 ( .A(n_294), .Y(n_293) );
OAI22xp5_ASAP7_75t_L g295 ( .A1(n_296), .A2(n_298), .B1(n_302), .B2(n_305), .Y(n_295) );
NAND2xp5_ASAP7_75t_L g298 ( .A(n_299), .B(n_300), .Y(n_298) );
NAND2xp5_ASAP7_75t_L g319 ( .A(n_299), .B(n_311), .Y(n_319) );
NAND2xp5_ASAP7_75t_L g344 ( .A(n_300), .B(n_345), .Y(n_344) );
INVx1_ASAP7_75t_SL g300 ( .A(n_301), .Y(n_300) );
INVx1_ASAP7_75t_L g302 ( .A(n_303), .Y(n_302) );
INVx1_ASAP7_75t_L g400 ( .A(n_304), .Y(n_400) );
AND2x2_ASAP7_75t_L g419 ( .A(n_304), .B(n_334), .Y(n_419) );
OR2x2_ASAP7_75t_L g305 ( .A(n_306), .B(n_307), .Y(n_305) );
INVx1_ASAP7_75t_L g309 ( .A(n_310), .Y(n_309) );
NAND2xp5_ASAP7_75t_L g427 ( .A(n_311), .B(n_368), .Y(n_427) );
INVx1_ASAP7_75t_L g312 ( .A(n_313), .Y(n_312) );
NOR2xp33_ASAP7_75t_L g425 ( .A(n_314), .B(n_382), .Y(n_425) );
INVx1_ASAP7_75t_L g318 ( .A(n_319), .Y(n_318) );
INVx1_ASAP7_75t_L g320 ( .A(n_321), .Y(n_320) );
INVx1_ASAP7_75t_L g322 ( .A(n_323), .Y(n_322) );
INVx1_ASAP7_75t_L g348 ( .A(n_326), .Y(n_348) );
BUFx2_ASAP7_75t_L g372 ( .A(n_327), .Y(n_372) );
OAI21xp5_ASAP7_75t_SL g328 ( .A1(n_329), .A2(n_331), .B(n_333), .Y(n_328) );
INVx1_ASAP7_75t_L g329 ( .A(n_330), .Y(n_329) );
INVx1_ASAP7_75t_L g331 ( .A(n_332), .Y(n_331) );
NOR3xp33_ASAP7_75t_L g335 ( .A(n_336), .B(n_351), .C(n_373), .Y(n_335) );
INVx1_ASAP7_75t_L g337 ( .A(n_338), .Y(n_337) );
OAI21xp5_ASAP7_75t_L g340 ( .A1(n_341), .A2(n_343), .B(n_346), .Y(n_340) );
INVx1_ASAP7_75t_L g341 ( .A(n_342), .Y(n_341) );
INVx1_ASAP7_75t_L g343 ( .A(n_344), .Y(n_343) );
INVx1_ASAP7_75t_SL g349 ( .A(n_350), .Y(n_349) );
A2O1A1Ixp33_ASAP7_75t_SL g351 ( .A1(n_352), .A2(n_355), .B(n_359), .C(n_362), .Y(n_351) );
NAND2xp5_ASAP7_75t_SL g384 ( .A(n_352), .B(n_385), .Y(n_384) );
INVx1_ASAP7_75t_L g352 ( .A(n_353), .Y(n_352) );
INVx1_ASAP7_75t_L g353 ( .A(n_354), .Y(n_353) );
INVx1_ASAP7_75t_L g355 ( .A(n_356), .Y(n_355) );
NOR2xp67_ASAP7_75t_SL g356 ( .A(n_357), .B(n_358), .Y(n_356) );
OR2x2_ASAP7_75t_L g359 ( .A(n_360), .B(n_361), .Y(n_359) );
INVx1_ASAP7_75t_SL g381 ( .A(n_361), .Y(n_381) );
OAI21xp5_ASAP7_75t_L g362 ( .A1(n_363), .A2(n_366), .B(n_370), .Y(n_362) );
AND2x4_ASAP7_75t_L g363 ( .A(n_364), .B(n_365), .Y(n_363) );
AND2x2_ASAP7_75t_L g386 ( .A(n_364), .B(n_387), .Y(n_386) );
INVx1_ASAP7_75t_L g366 ( .A(n_367), .Y(n_366) );
INVx1_ASAP7_75t_SL g368 ( .A(n_369), .Y(n_368) );
INVx1_ASAP7_75t_L g370 ( .A(n_371), .Y(n_370) );
INVx1_ASAP7_75t_L g374 ( .A(n_375), .Y(n_374) );
NOR2xp33_ASAP7_75t_L g375 ( .A(n_376), .B(n_378), .Y(n_375) );
INVx2_ASAP7_75t_L g376 ( .A(n_377), .Y(n_376) );
INVx1_ASAP7_75t_L g379 ( .A(n_380), .Y(n_379) );
AOI22xp33_ASAP7_75t_L g383 ( .A1(n_384), .A2(n_386), .B1(n_388), .B2(n_390), .Y(n_383) );
INVx2_ASAP7_75t_SL g404 ( .A(n_391), .Y(n_404) );
NOR3xp33_ASAP7_75t_L g392 ( .A(n_393), .B(n_408), .C(n_420), .Y(n_392) );
INVx1_ASAP7_75t_L g394 ( .A(n_395), .Y(n_394) );
INVxp67_ASAP7_75t_L g398 ( .A(n_399), .Y(n_398) );
INVxp67_ASAP7_75t_L g402 ( .A(n_403), .Y(n_402) );
NAND2xp5_ASAP7_75t_L g406 ( .A(n_404), .B(n_407), .Y(n_406) );
INVx1_ASAP7_75t_L g405 ( .A(n_406), .Y(n_405) );
OAI221xp5_ASAP7_75t_L g408 ( .A1(n_409), .A2(n_411), .B1(n_415), .B2(n_417), .C(n_418), .Y(n_408) );
A2O1A1Ixp33_ASAP7_75t_L g420 ( .A1(n_409), .A2(n_421), .B(n_422), .C(n_424), .Y(n_420) );
INVx1_ASAP7_75t_SL g409 ( .A(n_410), .Y(n_409) );
INVxp67_ASAP7_75t_L g411 ( .A(n_412), .Y(n_411) );
NOR2xp33_ASAP7_75t_L g412 ( .A(n_413), .B(n_414), .Y(n_412) );
INVx1_ASAP7_75t_L g415 ( .A(n_416), .Y(n_415) );
INVx1_ASAP7_75t_L g422 ( .A(n_423), .Y(n_422) );
AOI22xp5_ASAP7_75t_L g424 ( .A1(n_425), .A2(n_426), .B1(n_428), .B2(n_430), .Y(n_424) );
INVx1_ASAP7_75t_L g426 ( .A(n_427), .Y(n_426) );
INVx1_ASAP7_75t_L g428 ( .A(n_429), .Y(n_428) );
OAI22xp5_ASAP7_75t_L g455 ( .A1(n_431), .A2(n_456), .B1(n_459), .B2(n_461), .Y(n_455) );
INVx1_ASAP7_75t_L g433 ( .A(n_434), .Y(n_433) );
INVx1_ASAP7_75t_SL g434 ( .A(n_435), .Y(n_434) );
INVx1_ASAP7_75t_SL g435 ( .A(n_436), .Y(n_435) );
INVx2_ASAP7_75t_L g442 ( .A(n_436), .Y(n_442) );
INVx1_ASAP7_75t_SL g747 ( .A(n_436), .Y(n_747) );
BUFx2_ASAP7_75t_L g750 ( .A(n_436), .Y(n_750) );
NOR2x2_ASAP7_75t_L g742 ( .A(n_437), .B(n_460), .Y(n_742) );
INVx2_ASAP7_75t_L g437 ( .A(n_438), .Y(n_437) );
OR2x2_ASAP7_75t_L g459 ( .A(n_438), .B(n_460), .Y(n_459) );
AND2x2_ASAP7_75t_L g438 ( .A(n_439), .B(n_440), .Y(n_438) );
AND2x2_ASAP7_75t_L g443 ( .A(n_444), .B(n_447), .Y(n_443) );
INVx1_ASAP7_75t_L g444 ( .A(n_445), .Y(n_444) );
INVx1_ASAP7_75t_L g445 ( .A(n_446), .Y(n_445) );
NOR2xp33_ASAP7_75t_SL g745 ( .A(n_446), .B(n_448), .Y(n_745) );
OA21x2_ASAP7_75t_L g749 ( .A1(n_446), .A2(n_447), .B(n_750), .Y(n_749) );
INVx1_ASAP7_75t_SL g447 ( .A(n_448), .Y(n_447) );
INVxp67_ASAP7_75t_L g450 ( .A(n_451), .Y(n_450) );
INVx1_ASAP7_75t_L g735 ( .A(n_452), .Y(n_735) );
INVx2_ASAP7_75t_L g456 ( .A(n_457), .Y(n_456) );
INVx2_ASAP7_75t_L g737 ( .A(n_457), .Y(n_737) );
INVx1_ASAP7_75t_L g457 ( .A(n_458), .Y(n_457) );
INVx1_ASAP7_75t_L g739 ( .A(n_459), .Y(n_739) );
INVx1_ASAP7_75t_SL g461 ( .A(n_462), .Y(n_461) );
OR5x1_ASAP7_75t_L g462 ( .A(n_463), .B(n_629), .C(n_693), .D(n_709), .E(n_724), .Y(n_462) );
NAND4xp25_ASAP7_75t_L g463 ( .A(n_464), .B(n_563), .C(n_590), .D(n_613), .Y(n_463) );
AOI21xp5_ASAP7_75t_L g464 ( .A1(n_465), .A2(n_511), .B(n_522), .Y(n_464) );
NOR2xp33_ASAP7_75t_L g465 ( .A(n_466), .B(n_476), .Y(n_465) );
HB1xp67_ASAP7_75t_L g466 ( .A(n_467), .Y(n_466) );
INVx3_ASAP7_75t_SL g542 ( .A(n_467), .Y(n_542) );
AND2x4_ASAP7_75t_L g576 ( .A(n_467), .B(n_565), .Y(n_576) );
OR2x2_ASAP7_75t_L g586 ( .A(n_467), .B(n_544), .Y(n_586) );
OR2x2_ASAP7_75t_L g632 ( .A(n_467), .B(n_479), .Y(n_632) );
AND2x2_ASAP7_75t_L g646 ( .A(n_467), .B(n_543), .Y(n_646) );
AND2x2_ASAP7_75t_L g689 ( .A(n_467), .B(n_579), .Y(n_689) );
AND2x2_ASAP7_75t_L g696 ( .A(n_467), .B(n_554), .Y(n_696) );
AND2x2_ASAP7_75t_L g715 ( .A(n_467), .B(n_605), .Y(n_715) );
AND2x2_ASAP7_75t_L g733 ( .A(n_467), .B(n_575), .Y(n_733) );
OR2x6_ASAP7_75t_L g467 ( .A(n_468), .B(n_474), .Y(n_467) );
INVx1_ASAP7_75t_L g698 ( .A(n_476), .Y(n_698) );
NAND2xp5_ASAP7_75t_L g476 ( .A(n_477), .B(n_492), .Y(n_476) );
AND2x2_ASAP7_75t_L g608 ( .A(n_477), .B(n_543), .Y(n_608) );
NAND2xp5_ASAP7_75t_L g627 ( .A(n_477), .B(n_628), .Y(n_627) );
AOI32xp33_ASAP7_75t_L g641 ( .A1(n_477), .A2(n_642), .A3(n_645), .B1(n_647), .B2(n_651), .Y(n_641) );
AND2x2_ASAP7_75t_L g711 ( .A(n_477), .B(n_605), .Y(n_711) );
INVx2_ASAP7_75t_L g477 ( .A(n_478), .Y(n_477) );
INVx1_ASAP7_75t_SL g478 ( .A(n_479), .Y(n_478) );
AND2x2_ASAP7_75t_L g575 ( .A(n_479), .B(n_544), .Y(n_575) );
NAND2xp5_ASAP7_75t_L g584 ( .A(n_479), .B(n_585), .Y(n_584) );
AND2x2_ASAP7_75t_L g617 ( .A(n_479), .B(n_564), .Y(n_617) );
NAND2xp5_ASAP7_75t_L g695 ( .A(n_479), .B(n_696), .Y(n_695) );
AO21x2_ASAP7_75t_L g479 ( .A1(n_480), .A2(n_482), .B(n_490), .Y(n_479) );
INVx1_ASAP7_75t_L g580 ( .A(n_480), .Y(n_580) );
INVx1_ASAP7_75t_L g480 ( .A(n_481), .Y(n_480) );
INVx1_ASAP7_75t_L g482 ( .A(n_483), .Y(n_482) );
OA21x2_ASAP7_75t_L g579 ( .A1(n_483), .A2(n_491), .B(n_580), .Y(n_579) );
INVx1_ASAP7_75t_L g490 ( .A(n_491), .Y(n_490) );
AND2x2_ASAP7_75t_L g582 ( .A(n_492), .B(n_526), .Y(n_582) );
AND2x2_ASAP7_75t_L g658 ( .A(n_492), .B(n_659), .Y(n_658) );
INVx1_ASAP7_75t_SL g730 ( .A(n_492), .Y(n_730) );
AND2x2_ASAP7_75t_L g492 ( .A(n_493), .B(n_502), .Y(n_492) );
OR2x2_ASAP7_75t_L g525 ( .A(n_493), .B(n_503), .Y(n_525) );
AND2x2_ASAP7_75t_L g539 ( .A(n_493), .B(n_540), .Y(n_539) );
NOR2xp33_ASAP7_75t_L g567 ( .A(n_493), .B(n_568), .Y(n_567) );
INVx2_ASAP7_75t_L g589 ( .A(n_493), .Y(n_589) );
AND2x2_ASAP7_75t_L g616 ( .A(n_493), .B(n_503), .Y(n_616) );
BUFx3_ASAP7_75t_L g619 ( .A(n_493), .Y(n_619) );
NAND2xp5_ASAP7_75t_L g626 ( .A(n_493), .B(n_594), .Y(n_626) );
NAND2xp5_ASAP7_75t_L g712 ( .A(n_493), .B(n_713), .Y(n_712) );
INVx2_ASAP7_75t_L g570 ( .A(n_502), .Y(n_570) );
AND2x2_ASAP7_75t_L g588 ( .A(n_502), .B(n_568), .Y(n_588) );
INVx2_ASAP7_75t_L g502 ( .A(n_503), .Y(n_502) );
AND2x2_ASAP7_75t_L g599 ( .A(n_503), .B(n_513), .Y(n_599) );
HB1xp67_ASAP7_75t_L g612 ( .A(n_503), .Y(n_612) );
INVx1_ASAP7_75t_L g511 ( .A(n_512), .Y(n_511) );
NAND2xp5_ASAP7_75t_L g669 ( .A(n_512), .B(n_619), .Y(n_669) );
HB1xp67_ASAP7_75t_L g512 ( .A(n_513), .Y(n_512) );
INVx1_ASAP7_75t_SL g540 ( .A(n_513), .Y(n_540) );
NAND3xp33_ASAP7_75t_L g587 ( .A(n_513), .B(n_588), .C(n_589), .Y(n_587) );
OR2x2_ASAP7_75t_L g595 ( .A(n_513), .B(n_568), .Y(n_595) );
AND2x2_ASAP7_75t_L g615 ( .A(n_513), .B(n_568), .Y(n_615) );
AND2x2_ASAP7_75t_L g659 ( .A(n_513), .B(n_528), .Y(n_659) );
AOI21xp5_ASAP7_75t_L g522 ( .A1(n_523), .A2(n_538), .B(n_541), .Y(n_522) );
NAND2xp5_ASAP7_75t_SL g523 ( .A(n_524), .B(n_526), .Y(n_523) );
AND2x2_ASAP7_75t_L g734 ( .A(n_524), .B(n_659), .Y(n_734) );
INVx1_ASAP7_75t_L g524 ( .A(n_525), .Y(n_524) );
OAI22xp5_ASAP7_75t_L g673 ( .A1(n_525), .A2(n_632), .B1(n_674), .B2(n_676), .Y(n_673) );
OR2x2_ASAP7_75t_L g680 ( .A(n_525), .B(n_595), .Y(n_680) );
OR2x2_ASAP7_75t_L g704 ( .A(n_525), .B(n_705), .Y(n_704) );
NOR2xp33_ASAP7_75t_L g717 ( .A(n_525), .B(n_624), .Y(n_717) );
AND2x2_ASAP7_75t_L g610 ( .A(n_526), .B(n_611), .Y(n_610) );
AOI21xp5_ASAP7_75t_L g697 ( .A1(n_526), .A2(n_683), .B(n_698), .Y(n_697) );
AOI32xp33_ASAP7_75t_L g718 ( .A1(n_526), .A2(n_608), .A3(n_719), .B1(n_721), .B2(n_722), .Y(n_718) );
OR2x2_ASAP7_75t_L g729 ( .A(n_526), .B(n_730), .Y(n_729) );
CKINVDCx16_ASAP7_75t_R g526 ( .A(n_527), .Y(n_526) );
OR2x2_ASAP7_75t_L g597 ( .A(n_527), .B(n_598), .Y(n_597) );
NAND2xp5_ASAP7_75t_L g676 ( .A(n_527), .B(n_611), .Y(n_676) );
BUFx3_ASAP7_75t_L g527 ( .A(n_528), .Y(n_527) );
INVx4_ASAP7_75t_L g568 ( .A(n_528), .Y(n_568) );
AND2x2_ASAP7_75t_L g634 ( .A(n_528), .B(n_599), .Y(n_634) );
AND3x2_ASAP7_75t_L g643 ( .A(n_528), .B(n_539), .C(n_644), .Y(n_643) );
INVx1_ASAP7_75t_L g538 ( .A(n_539), .Y(n_538) );
AND2x2_ASAP7_75t_L g569 ( .A(n_540), .B(n_570), .Y(n_569) );
HB1xp67_ASAP7_75t_L g624 ( .A(n_540), .Y(n_624) );
NAND2xp5_ASAP7_75t_L g705 ( .A(n_540), .B(n_568), .Y(n_705) );
NAND2xp5_ASAP7_75t_L g541 ( .A(n_542), .B(n_543), .Y(n_541) );
AND2x2_ASAP7_75t_L g564 ( .A(n_542), .B(n_565), .Y(n_564) );
AND2x2_ASAP7_75t_L g604 ( .A(n_542), .B(n_605), .Y(n_604) );
AND2x2_ASAP7_75t_L g622 ( .A(n_542), .B(n_554), .Y(n_622) );
AND2x2_ASAP7_75t_L g640 ( .A(n_542), .B(n_544), .Y(n_640) );
OR2x2_ASAP7_75t_L g654 ( .A(n_542), .B(n_655), .Y(n_654) );
AND2x2_ASAP7_75t_L g700 ( .A(n_542), .B(n_628), .Y(n_700) );
NAND2xp5_ASAP7_75t_L g578 ( .A(n_543), .B(n_579), .Y(n_578) );
AND2x2_ASAP7_75t_L g543 ( .A(n_544), .B(n_554), .Y(n_543) );
AND2x2_ASAP7_75t_L g601 ( .A(n_544), .B(n_579), .Y(n_601) );
OR2x2_ASAP7_75t_L g655 ( .A(n_544), .B(n_579), .Y(n_655) );
AND2x2_ASAP7_75t_L g708 ( .A(n_544), .B(n_565), .Y(n_708) );
INVx2_ASAP7_75t_SL g544 ( .A(n_545), .Y(n_544) );
BUFx2_ASAP7_75t_L g606 ( .A(n_545), .Y(n_606) );
AND2x2_ASAP7_75t_L g628 ( .A(n_545), .B(n_554), .Y(n_628) );
INVx2_ASAP7_75t_L g565 ( .A(n_554), .Y(n_565) );
INVx1_ASAP7_75t_L g585 ( .A(n_554), .Y(n_585) );
AOI211xp5_ASAP7_75t_L g563 ( .A1(n_564), .A2(n_566), .B(n_571), .C(n_583), .Y(n_563) );
NAND2xp5_ASAP7_75t_L g674 ( .A(n_564), .B(n_675), .Y(n_674) );
INVx1_ASAP7_75t_L g727 ( .A(n_564), .Y(n_727) );
AND2x2_ASAP7_75t_L g605 ( .A(n_565), .B(n_606), .Y(n_605) );
AND2x2_ASAP7_75t_L g566 ( .A(n_567), .B(n_569), .Y(n_566) );
NAND2xp5_ASAP7_75t_L g577 ( .A(n_568), .B(n_569), .Y(n_577) );
INVx1_ASAP7_75t_L g662 ( .A(n_568), .Y(n_662) );
NAND2xp5_ASAP7_75t_L g686 ( .A(n_568), .B(n_589), .Y(n_686) );
AND2x2_ASAP7_75t_L g702 ( .A(n_568), .B(n_616), .Y(n_702) );
NAND2xp5_ASAP7_75t_SL g684 ( .A(n_569), .B(n_685), .Y(n_684) );
INVx2_ASAP7_75t_L g593 ( .A(n_570), .Y(n_593) );
OAI22xp5_ASAP7_75t_L g571 ( .A1(n_572), .A2(n_577), .B1(n_578), .B2(n_581), .Y(n_571) );
INVx1_ASAP7_75t_L g572 ( .A(n_573), .Y(n_572) );
NOR2xp33_ASAP7_75t_L g573 ( .A(n_574), .B(n_576), .Y(n_573) );
NOR2xp33_ASAP7_75t_L g726 ( .A(n_574), .B(n_727), .Y(n_726) );
INVx1_ASAP7_75t_L g574 ( .A(n_575), .Y(n_574) );
NAND2xp5_ASAP7_75t_L g621 ( .A(n_575), .B(n_622), .Y(n_621) );
AND2x2_ASAP7_75t_L g600 ( .A(n_576), .B(n_601), .Y(n_600) );
AOI221xp5_ASAP7_75t_SL g665 ( .A1(n_576), .A2(n_618), .B1(n_666), .B2(n_671), .C(n_673), .Y(n_665) );
NAND2xp5_ASAP7_75t_L g672 ( .A(n_576), .B(n_639), .Y(n_672) );
INVx1_ASAP7_75t_L g732 ( .A(n_578), .Y(n_732) );
BUFx3_ASAP7_75t_L g639 ( .A(n_579), .Y(n_639) );
INVx1_ASAP7_75t_L g581 ( .A(n_582), .Y(n_581) );
AOI21xp33_ASAP7_75t_SL g583 ( .A1(n_584), .A2(n_586), .B(n_587), .Y(n_583) );
INVx1_ASAP7_75t_L g648 ( .A(n_585), .Y(n_648) );
NAND2xp5_ASAP7_75t_L g692 ( .A(n_585), .B(n_639), .Y(n_692) );
INVx1_ASAP7_75t_L g649 ( .A(n_586), .Y(n_649) );
NAND2xp5_ASAP7_75t_SL g650 ( .A(n_586), .B(n_639), .Y(n_650) );
INVxp67_ASAP7_75t_L g670 ( .A(n_588), .Y(n_670) );
AND2x2_ASAP7_75t_L g611 ( .A(n_589), .B(n_612), .Y(n_611) );
O2A1O1Ixp33_ASAP7_75t_L g590 ( .A1(n_591), .A2(n_596), .B(n_600), .C(n_602), .Y(n_590) );
INVx1_ASAP7_75t_L g591 ( .A(n_592), .Y(n_591) );
NAND2xp5_ASAP7_75t_L g592 ( .A(n_593), .B(n_594), .Y(n_592) );
INVx1_ASAP7_75t_SL g625 ( .A(n_593), .Y(n_625) );
NAND2xp5_ASAP7_75t_L g636 ( .A(n_594), .B(n_625), .Y(n_636) );
NAND2xp5_ASAP7_75t_L g667 ( .A(n_594), .B(n_616), .Y(n_667) );
INVx2_ASAP7_75t_SL g594 ( .A(n_595), .Y(n_594) );
INVx1_ASAP7_75t_L g596 ( .A(n_597), .Y(n_596) );
OAI22xp5_ASAP7_75t_L g602 ( .A1(n_597), .A2(n_603), .B1(n_607), .B2(n_609), .Y(n_602) );
INVx1_ASAP7_75t_SL g598 ( .A(n_599), .Y(n_598) );
AND2x2_ASAP7_75t_L g618 ( .A(n_599), .B(n_619), .Y(n_618) );
AND2x2_ASAP7_75t_L g663 ( .A(n_599), .B(n_664), .Y(n_663) );
OAI21xp33_ASAP7_75t_L g666 ( .A1(n_601), .A2(n_667), .B(n_668), .Y(n_666) );
INVx1_ASAP7_75t_SL g603 ( .A(n_604), .Y(n_603) );
AOI221xp5_ASAP7_75t_L g613 ( .A1(n_605), .A2(n_614), .B1(n_617), .B2(n_618), .C(n_620), .Y(n_613) );
NAND2xp5_ASAP7_75t_L g682 ( .A(n_605), .B(n_639), .Y(n_682) );
NAND2xp5_ASAP7_75t_L g688 ( .A(n_605), .B(n_689), .Y(n_688) );
INVx1_ASAP7_75t_L g607 ( .A(n_608), .Y(n_607) );
INVx1_ASAP7_75t_L g609 ( .A(n_610), .Y(n_609) );
INVx1_ASAP7_75t_L g721 ( .A(n_611), .Y(n_721) );
INVxp67_ASAP7_75t_L g644 ( .A(n_612), .Y(n_644) );
INVx1_ASAP7_75t_L g651 ( .A(n_614), .Y(n_651) );
AND2x2_ASAP7_75t_L g614 ( .A(n_615), .B(n_616), .Y(n_614) );
AND2x2_ASAP7_75t_L g690 ( .A(n_615), .B(n_619), .Y(n_690) );
INVx1_ASAP7_75t_L g664 ( .A(n_619), .Y(n_664) );
NAND2xp5_ASAP7_75t_SL g694 ( .A(n_619), .B(n_634), .Y(n_694) );
OAI32xp33_ASAP7_75t_L g620 ( .A1(n_621), .A2(n_623), .A3(n_625), .B1(n_626), .B2(n_627), .Y(n_620) );
INVx1_ASAP7_75t_L g623 ( .A(n_624), .Y(n_623) );
INVx2_ASAP7_75t_SL g633 ( .A(n_628), .Y(n_633) );
NAND2xp5_ASAP7_75t_L g677 ( .A(n_628), .B(n_660), .Y(n_677) );
NAND2xp5_ASAP7_75t_L g720 ( .A(n_628), .B(n_689), .Y(n_720) );
NAND2x1p5_ASAP7_75t_L g728 ( .A(n_628), .B(n_639), .Y(n_728) );
NAND5xp2_ASAP7_75t_L g629 ( .A(n_630), .B(n_652), .C(n_665), .D(n_677), .E(n_678), .Y(n_629) );
AOI221xp5_ASAP7_75t_L g630 ( .A1(n_631), .A2(n_634), .B1(n_635), .B2(n_637), .C(n_641), .Y(n_630) );
NOR2xp33_ASAP7_75t_L g631 ( .A(n_632), .B(n_633), .Y(n_631) );
INVx1_ASAP7_75t_L g635 ( .A(n_636), .Y(n_635) );
NAND2xp33_ASAP7_75t_SL g656 ( .A(n_636), .B(n_657), .Y(n_656) );
INVx1_ASAP7_75t_L g637 ( .A(n_638), .Y(n_637) );
NAND2xp5_ASAP7_75t_L g638 ( .A(n_639), .B(n_640), .Y(n_638) );
NAND2xp5_ASAP7_75t_L g707 ( .A(n_639), .B(n_708), .Y(n_707) );
AOI22xp33_ASAP7_75t_L g652 ( .A1(n_640), .A2(n_653), .B1(n_656), .B2(n_660), .Y(n_652) );
INVx2_ASAP7_75t_SL g642 ( .A(n_643), .Y(n_642) );
OAI211xp5_ASAP7_75t_SL g647 ( .A1(n_643), .A2(n_648), .B(n_649), .C(n_650), .Y(n_647) );
INVx1_ASAP7_75t_L g645 ( .A(n_646), .Y(n_645) );
INVx1_ASAP7_75t_L g653 ( .A(n_654), .Y(n_653) );
INVx1_ASAP7_75t_SL g675 ( .A(n_655), .Y(n_675) );
INVx1_ASAP7_75t_SL g657 ( .A(n_658), .Y(n_657) );
INVx1_ASAP7_75t_SL g660 ( .A(n_661), .Y(n_660) );
NAND2xp5_ASAP7_75t_L g661 ( .A(n_662), .B(n_663), .Y(n_661) );
NAND2xp5_ASAP7_75t_L g723 ( .A(n_664), .B(n_713), .Y(n_723) );
OR2x2_ASAP7_75t_L g668 ( .A(n_669), .B(n_670), .Y(n_668) );
INVx1_ASAP7_75t_L g671 ( .A(n_672), .Y(n_671) );
AOI222xp33_ASAP7_75t_L g678 ( .A1(n_679), .A2(n_681), .B1(n_683), .B2(n_687), .C1(n_690), .C2(n_691), .Y(n_678) );
INVx1_ASAP7_75t_L g679 ( .A(n_680), .Y(n_679) );
INVx1_ASAP7_75t_L g681 ( .A(n_682), .Y(n_681) );
INVx1_ASAP7_75t_L g683 ( .A(n_684), .Y(n_683) );
INVx1_ASAP7_75t_L g685 ( .A(n_686), .Y(n_685) );
INVx1_ASAP7_75t_L g687 ( .A(n_688), .Y(n_687) );
INVx1_ASAP7_75t_L g691 ( .A(n_692), .Y(n_691) );
OAI221xp5_ASAP7_75t_L g693 ( .A1(n_694), .A2(n_695), .B1(n_697), .B2(n_699), .C(n_701), .Y(n_693) );
INVx1_ASAP7_75t_SL g699 ( .A(n_700), .Y(n_699) );
OAI21xp33_ASAP7_75t_L g701 ( .A1(n_702), .A2(n_703), .B(n_706), .Y(n_701) );
INVx2_ASAP7_75t_L g703 ( .A(n_704), .Y(n_703) );
INVx1_ASAP7_75t_L g713 ( .A(n_705), .Y(n_713) );
INVx1_ASAP7_75t_L g706 ( .A(n_707), .Y(n_706) );
OAI221xp5_ASAP7_75t_L g709 ( .A1(n_710), .A2(n_712), .B1(n_714), .B2(n_716), .C(n_718), .Y(n_709) );
INVx1_ASAP7_75t_L g710 ( .A(n_711), .Y(n_710) );
INVx1_ASAP7_75t_SL g714 ( .A(n_715), .Y(n_714) );
INVxp67_ASAP7_75t_L g716 ( .A(n_717), .Y(n_716) );
INVx1_ASAP7_75t_L g719 ( .A(n_720), .Y(n_719) );
INVx1_ASAP7_75t_L g722 ( .A(n_723), .Y(n_722) );
A2O1A1Ixp33_ASAP7_75t_L g724 ( .A1(n_725), .A2(n_728), .B(n_729), .C(n_731), .Y(n_724) );
INVxp67_ASAP7_75t_L g725 ( .A(n_726), .Y(n_725) );
OAI21xp33_ASAP7_75t_L g731 ( .A1(n_732), .A2(n_733), .B(n_734), .Y(n_731) );
INVx2_ASAP7_75t_L g738 ( .A(n_739), .Y(n_738) );
INVx1_ASAP7_75t_SL g740 ( .A(n_741), .Y(n_740) );
INVx3_ASAP7_75t_SL g741 ( .A(n_742), .Y(n_741) );
INVx1_ASAP7_75t_SL g743 ( .A(n_744), .Y(n_743) );
NAND2xp33_ASAP7_75t_L g744 ( .A(n_745), .B(n_746), .Y(n_744) );
INVx1_ASAP7_75t_SL g746 ( .A(n_747), .Y(n_746) );
INVx1_ASAP7_75t_SL g748 ( .A(n_749), .Y(n_748) );
endmodule