module fake_netlist_1_3684_n_11 (n_1, n_2, n_0, n_11);
input n_1;
input n_2;
input n_0;
output n_11;
wire n_6;
wire n_4;
wire n_3;
wire n_9;
wire n_5;
wire n_7;
wire n_8;
BUFx6f_ASAP7_75t_L g3 ( .A(n_2), .Y(n_3) );
INVx1_ASAP7_75t_SL g4 ( .A(n_0), .Y(n_4) );
INVx2_ASAP7_75t_L g5 ( .A(n_3), .Y(n_5) );
OR2x2_ASAP7_75t_L g6 ( .A(n_4), .B(n_0), .Y(n_6) );
AOI33xp33_ASAP7_75t_L g7 ( .A1(n_5), .A2(n_0), .A3(n_1), .B1(n_2), .B2(n_3), .B3(n_6), .Y(n_7) );
INVx1_ASAP7_75t_L g8 ( .A(n_7), .Y(n_8) );
AOI22xp5_ASAP7_75t_L g9 ( .A1(n_8), .A2(n_1), .B1(n_3), .B2(n_6), .Y(n_9) );
HB1xp67_ASAP7_75t_L g10 ( .A(n_9), .Y(n_10) );
UNKNOWN g11 ( );
endmodule