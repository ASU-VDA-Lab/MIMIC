module fake_netlist_5_251_n_2457 (n_137, n_210, n_168, n_164, n_191, n_91, n_208, n_82, n_122, n_194, n_142, n_176, n_10, n_214, n_140, n_24, n_124, n_86, n_136, n_146, n_182, n_143, n_83, n_132, n_61, n_237, n_90, n_127, n_75, n_101, n_180, n_184, n_226, n_235, n_65, n_78, n_74, n_144, n_207, n_114, n_57, n_96, n_37, n_189, n_220, n_165, n_111, n_229, n_108, n_231, n_213, n_129, n_31, n_13, n_66, n_98, n_177, n_60, n_155, n_152, n_197, n_16, n_43, n_107, n_0, n_58, n_9, n_69, n_236, n_18, n_116, n_195, n_42, n_22, n_227, n_1, n_45, n_117, n_46, n_233, n_21, n_94, n_203, n_205, n_113, n_38, n_123, n_139, n_105, n_80, n_4, n_179, n_125, n_35, n_167, n_128, n_73, n_234, n_17, n_92, n_19, n_149, n_120, n_232, n_135, n_30, n_156, n_5, n_33, n_126, n_14, n_225, n_84, n_23, n_202, n_130, n_219, n_157, n_29, n_79, n_193, n_131, n_151, n_47, n_173, n_192, n_25, n_53, n_160, n_198, n_223, n_188, n_190, n_8, n_201, n_158, n_44, n_224, n_40, n_34, n_100, n_62, n_138, n_148, n_71, n_154, n_228, n_109, n_112, n_212, n_85, n_159, n_163, n_95, n_119, n_183, n_185, n_175, n_169, n_59, n_26, n_133, n_238, n_215, n_55, n_196, n_99, n_2, n_211, n_218, n_181, n_3, n_49, n_20, n_6, n_39, n_54, n_147, n_178, n_221, n_12, n_67, n_121, n_36, n_76, n_200, n_87, n_150, n_162, n_27, n_170, n_64, n_77, n_102, n_106, n_161, n_209, n_222, n_230, n_81, n_118, n_28, n_89, n_70, n_115, n_68, n_93, n_72, n_174, n_186, n_199, n_134, n_187, n_32, n_41, n_104, n_172, n_103, n_56, n_51, n_63, n_97, n_141, n_166, n_11, n_206, n_217, n_171, n_153, n_7, n_15, n_145, n_48, n_204, n_50, n_52, n_88, n_110, n_216, n_2457);

input n_137;
input n_210;
input n_168;
input n_164;
input n_191;
input n_91;
input n_208;
input n_82;
input n_122;
input n_194;
input n_142;
input n_176;
input n_10;
input n_214;
input n_140;
input n_24;
input n_124;
input n_86;
input n_136;
input n_146;
input n_182;
input n_143;
input n_83;
input n_132;
input n_61;
input n_237;
input n_90;
input n_127;
input n_75;
input n_101;
input n_180;
input n_184;
input n_226;
input n_235;
input n_65;
input n_78;
input n_74;
input n_144;
input n_207;
input n_114;
input n_57;
input n_96;
input n_37;
input n_189;
input n_220;
input n_165;
input n_111;
input n_229;
input n_108;
input n_231;
input n_213;
input n_129;
input n_31;
input n_13;
input n_66;
input n_98;
input n_177;
input n_60;
input n_155;
input n_152;
input n_197;
input n_16;
input n_43;
input n_107;
input n_0;
input n_58;
input n_9;
input n_69;
input n_236;
input n_18;
input n_116;
input n_195;
input n_42;
input n_22;
input n_227;
input n_1;
input n_45;
input n_117;
input n_46;
input n_233;
input n_21;
input n_94;
input n_203;
input n_205;
input n_113;
input n_38;
input n_123;
input n_139;
input n_105;
input n_80;
input n_4;
input n_179;
input n_125;
input n_35;
input n_167;
input n_128;
input n_73;
input n_234;
input n_17;
input n_92;
input n_19;
input n_149;
input n_120;
input n_232;
input n_135;
input n_30;
input n_156;
input n_5;
input n_33;
input n_126;
input n_14;
input n_225;
input n_84;
input n_23;
input n_202;
input n_130;
input n_219;
input n_157;
input n_29;
input n_79;
input n_193;
input n_131;
input n_151;
input n_47;
input n_173;
input n_192;
input n_25;
input n_53;
input n_160;
input n_198;
input n_223;
input n_188;
input n_190;
input n_8;
input n_201;
input n_158;
input n_44;
input n_224;
input n_40;
input n_34;
input n_100;
input n_62;
input n_138;
input n_148;
input n_71;
input n_154;
input n_228;
input n_109;
input n_112;
input n_212;
input n_85;
input n_159;
input n_163;
input n_95;
input n_119;
input n_183;
input n_185;
input n_175;
input n_169;
input n_59;
input n_26;
input n_133;
input n_238;
input n_215;
input n_55;
input n_196;
input n_99;
input n_2;
input n_211;
input n_218;
input n_181;
input n_3;
input n_49;
input n_20;
input n_6;
input n_39;
input n_54;
input n_147;
input n_178;
input n_221;
input n_12;
input n_67;
input n_121;
input n_36;
input n_76;
input n_200;
input n_87;
input n_150;
input n_162;
input n_27;
input n_170;
input n_64;
input n_77;
input n_102;
input n_106;
input n_161;
input n_209;
input n_222;
input n_230;
input n_81;
input n_118;
input n_28;
input n_89;
input n_70;
input n_115;
input n_68;
input n_93;
input n_72;
input n_174;
input n_186;
input n_199;
input n_134;
input n_187;
input n_32;
input n_41;
input n_104;
input n_172;
input n_103;
input n_56;
input n_51;
input n_63;
input n_97;
input n_141;
input n_166;
input n_11;
input n_206;
input n_217;
input n_171;
input n_153;
input n_7;
input n_15;
input n_145;
input n_48;
input n_204;
input n_50;
input n_52;
input n_88;
input n_110;
input n_216;

output n_2457;

wire n_924;
wire n_1263;
wire n_977;
wire n_1378;
wire n_2253;
wire n_2417;
wire n_611;
wire n_1126;
wire n_1423;
wire n_1729;
wire n_1166;
wire n_2380;
wire n_1751;
wire n_469;
wire n_1508;
wire n_785;
wire n_549;
wire n_2200;
wire n_532;
wire n_1161;
wire n_1859;
wire n_1677;
wire n_1150;
wire n_2327;
wire n_1780;
wire n_1488;
wire n_667;
wire n_790;
wire n_1055;
wire n_2386;
wire n_1501;
wire n_2395;
wire n_880;
wire n_544;
wire n_1007;
wire n_2369;
wire n_552;
wire n_1528;
wire n_1370;
wire n_1292;
wire n_2347;
wire n_1198;
wire n_1360;
wire n_2388;
wire n_1099;
wire n_956;
wire n_564;
wire n_423;
wire n_1738;
wire n_2021;
wire n_2134;
wire n_2391;
wire n_1021;
wire n_1960;
wire n_2185;
wire n_551;
wire n_2143;
wire n_2059;
wire n_1323;
wire n_1466;
wire n_688;
wire n_1695;
wire n_1353;
wire n_800;
wire n_1347;
wire n_1535;
wire n_1789;
wire n_1666;
wire n_2389;
wire n_671;
wire n_819;
wire n_1451;
wire n_1022;
wire n_2302;
wire n_915;
wire n_1545;
wire n_2374;
wire n_864;
wire n_859;
wire n_951;
wire n_1947;
wire n_1264;
wire n_2114;
wire n_447;
wire n_247;
wire n_2001;
wire n_1494;
wire n_292;
wire n_625;
wire n_854;
wire n_1462;
wire n_1799;
wire n_2069;
wire n_2396;
wire n_1580;
wire n_674;
wire n_417;
wire n_1939;
wire n_1806;
wire n_516;
wire n_933;
wire n_2244;
wire n_2257;
wire n_1152;
wire n_497;
wire n_1869;
wire n_1607;
wire n_1563;
wire n_606;
wire n_275;
wire n_2011;
wire n_2096;
wire n_877;
wire n_2105;
wire n_2024;
wire n_1696;
wire n_1118;
wire n_755;
wire n_1686;
wire n_947;
wire n_1285;
wire n_373;
wire n_307;
wire n_1860;
wire n_1359;
wire n_530;
wire n_1107;
wire n_1728;
wire n_556;
wire n_2031;
wire n_2076;
wire n_1230;
wire n_668;
wire n_375;
wire n_301;
wire n_1896;
wire n_2165;
wire n_2147;
wire n_929;
wire n_1124;
wire n_1818;
wire n_2127;
wire n_902;
wire n_1576;
wire n_1104;
wire n_1294;
wire n_659;
wire n_1705;
wire n_1257;
wire n_1182;
wire n_579;
wire n_1698;
wire n_1261;
wire n_2329;
wire n_938;
wire n_1098;
wire n_2142;
wire n_320;
wire n_1154;
wire n_2189;
wire n_1242;
wire n_1135;
wire n_406;
wire n_519;
wire n_2323;
wire n_2203;
wire n_1016;
wire n_1243;
wire n_546;
wire n_2047;
wire n_1280;
wire n_1845;
wire n_281;
wire n_240;
wire n_2052;
wire n_2193;
wire n_2058;
wire n_291;
wire n_257;
wire n_731;
wire n_371;
wire n_1483;
wire n_1314;
wire n_1512;
wire n_709;
wire n_1490;
wire n_317;
wire n_1236;
wire n_1633;
wire n_569;
wire n_2144;
wire n_1778;
wire n_2306;
wire n_920;
wire n_1289;
wire n_1517;
wire n_2091;
wire n_335;
wire n_2085;
wire n_1669;
wire n_370;
wire n_976;
wire n_1949;
wire n_343;
wire n_1449;
wire n_308;
wire n_1946;
wire n_1566;
wire n_2032;
wire n_297;
wire n_2149;
wire n_1078;
wire n_1670;
wire n_775;
wire n_600;
wire n_1484;
wire n_2071;
wire n_1374;
wire n_1328;
wire n_2141;
wire n_1948;
wire n_1984;
wire n_2099;
wire n_2408;
wire n_264;
wire n_1877;
wire n_1831;
wire n_1598;
wire n_1723;
wire n_955;
wire n_1850;
wire n_339;
wire n_1146;
wire n_882;
wire n_243;
wire n_2384;
wire n_1036;
wire n_1097;
wire n_1749;
wire n_347;
wire n_550;
wire n_696;
wire n_897;
wire n_798;
wire n_350;
wire n_646;
wire n_1428;
wire n_436;
wire n_1394;
wire n_1414;
wire n_1216;
wire n_580;
wire n_290;
wire n_1040;
wire n_2202;
wire n_1872;
wire n_1852;
wire n_2159;
wire n_578;
wire n_926;
wire n_2180;
wire n_2249;
wire n_344;
wire n_2353;
wire n_1218;
wire n_1931;
wire n_2439;
wire n_2276;
wire n_422;
wire n_475;
wire n_1070;
wire n_777;
wire n_1547;
wire n_2089;
wire n_1030;
wire n_1755;
wire n_415;
wire n_1071;
wire n_485;
wire n_1165;
wire n_1267;
wire n_1561;
wire n_496;
wire n_1801;
wire n_1391;
wire n_958;
wire n_1034;
wire n_670;
wire n_1513;
wire n_1600;
wire n_521;
wire n_663;
wire n_845;
wire n_2235;
wire n_1862;
wire n_673;
wire n_837;
wire n_1239;
wire n_528;
wire n_2300;
wire n_1796;
wire n_680;
wire n_1473;
wire n_1587;
wire n_395;
wire n_901;
wire n_553;
wire n_2432;
wire n_813;
wire n_1521;
wire n_1284;
wire n_1590;
wire n_2174;
wire n_1748;
wire n_1672;
wire n_675;
wire n_888;
wire n_1880;
wire n_2337;
wire n_1167;
wire n_1626;
wire n_637;
wire n_1384;
wire n_1556;
wire n_446;
wire n_1863;
wire n_1064;
wire n_858;
wire n_2079;
wire n_2238;
wire n_923;
wire n_2118;
wire n_691;
wire n_1151;
wire n_881;
wire n_1405;
wire n_2407;
wire n_1706;
wire n_468;
wire n_342;
wire n_464;
wire n_363;
wire n_1582;
wire n_1069;
wire n_1784;
wire n_1075;
wire n_1836;
wire n_1450;
wire n_1322;
wire n_2101;
wire n_1471;
wire n_1986;
wire n_2072;
wire n_1750;
wire n_1459;
wire n_460;
wire n_889;
wire n_2358;
wire n_973;
wire n_1700;
wire n_477;
wire n_571;
wire n_1585;
wire n_461;
wire n_1971;
wire n_1599;
wire n_2275;
wire n_1211;
wire n_1197;
wire n_1523;
wire n_1950;
wire n_907;
wire n_1447;
wire n_2251;
wire n_1377;
wire n_2370;
wire n_989;
wire n_1039;
wire n_2214;
wire n_2055;
wire n_283;
wire n_1403;
wire n_2248;
wire n_2356;
wire n_488;
wire n_736;
wire n_892;
wire n_1000;
wire n_1202;
wire n_1278;
wire n_2062;
wire n_1002;
wire n_1581;
wire n_1463;
wire n_2100;
wire n_310;
wire n_593;
wire n_2258;
wire n_748;
wire n_586;
wire n_1058;
wire n_1667;
wire n_838;
wire n_332;
wire n_1053;
wire n_1224;
wire n_349;
wire n_1926;
wire n_1248;
wire n_1331;
wire n_953;
wire n_279;
wire n_1014;
wire n_1241;
wire n_2150;
wire n_2241;
wire n_2152;
wire n_289;
wire n_963;
wire n_1052;
wire n_954;
wire n_627;
wire n_1385;
wire n_440;
wire n_793;
wire n_478;
wire n_2140;
wire n_2385;
wire n_1819;
wire n_2330;
wire n_2139;
wire n_476;
wire n_1527;
wire n_2042;
wire n_534;
wire n_1882;
wire n_884;
wire n_345;
wire n_944;
wire n_1754;
wire n_1623;
wire n_2175;
wire n_2324;
wire n_1854;
wire n_1565;
wire n_1809;
wire n_1856;
wire n_647;
wire n_407;
wire n_1072;
wire n_2218;
wire n_2267;
wire n_857;
wire n_832;
wire n_2305;
wire n_2450;
wire n_1319;
wire n_561;
wire n_2379;
wire n_2154;
wire n_1825;
wire n_1951;
wire n_1906;
wire n_1883;
wire n_1712;
wire n_1387;
wire n_2262;
wire n_1532;
wire n_2322;
wire n_2271;
wire n_1027;
wire n_971;
wire n_1156;
wire n_326;
wire n_794;
wire n_404;
wire n_2331;
wire n_2293;
wire n_686;
wire n_847;
wire n_1393;
wire n_2319;
wire n_596;
wire n_1775;
wire n_2028;
wire n_1368;
wire n_558;
wire n_702;
wire n_1276;
wire n_822;
wire n_1412;
wire n_1709;
wire n_2108;
wire n_728;
wire n_266;
wire n_1162;
wire n_272;
wire n_1538;
wire n_1838;
wire n_1199;
wire n_1847;
wire n_1779;
wire n_352;
wire n_1884;
wire n_2434;
wire n_1038;
wire n_520;
wire n_1369;
wire n_409;
wire n_1841;
wire n_1660;
wire n_887;
wire n_1905;
wire n_2195;
wire n_300;
wire n_809;
wire n_931;
wire n_870;
wire n_599;
wire n_1711;
wire n_1662;
wire n_1891;
wire n_1481;
wire n_1942;
wire n_434;
wire n_1978;
wire n_1544;
wire n_868;
wire n_2454;
wire n_639;
wire n_914;
wire n_2120;
wire n_411;
wire n_414;
wire n_1629;
wire n_1293;
wire n_965;
wire n_1876;
wire n_1743;
wire n_935;
wire n_817;
wire n_1175;
wire n_360;
wire n_1479;
wire n_1810;
wire n_2350;
wire n_1888;
wire n_2009;
wire n_759;
wire n_2222;
wire n_1892;
wire n_806;
wire n_1997;
wire n_1766;
wire n_1477;
wire n_324;
wire n_1635;
wire n_1963;
wire n_2226;
wire n_1571;
wire n_1189;
wire n_2215;
wire n_1259;
wire n_1690;
wire n_706;
wire n_746;
wire n_1649;
wire n_747;
wire n_2064;
wire n_784;
wire n_2449;
wire n_1733;
wire n_1244;
wire n_2413;
wire n_431;
wire n_1194;
wire n_1925;
wire n_2297;
wire n_1815;
wire n_615;
wire n_851;
wire n_1759;
wire n_843;
wire n_1788;
wire n_2177;
wire n_523;
wire n_913;
wire n_1537;
wire n_705;
wire n_865;
wire n_2227;
wire n_678;
wire n_697;
wire n_1222;
wire n_1679;
wire n_2190;
wire n_776;
wire n_1798;
wire n_2022;
wire n_1790;
wire n_1415;
wire n_367;
wire n_452;
wire n_525;
wire n_1260;
wire n_1746;
wire n_1647;
wire n_2181;
wire n_1829;
wire n_1464;
wire n_649;
wire n_547;
wire n_1444;
wire n_1191;
wire n_2387;
wire n_1674;
wire n_1833;
wire n_1830;
wire n_2073;
wire n_1710;
wire n_284;
wire n_1128;
wire n_1734;
wire n_744;
wire n_590;
wire n_629;
wire n_1308;
wire n_2178;
wire n_1767;
wire n_2336;
wire n_254;
wire n_1680;
wire n_1233;
wire n_1615;
wire n_1529;
wire n_2005;
wire n_526;
wire n_1916;
wire n_293;
wire n_372;
wire n_677;
wire n_244;
wire n_1333;
wire n_1121;
wire n_368;
wire n_604;
wire n_314;
wire n_433;
wire n_2007;
wire n_949;
wire n_1443;
wire n_1008;
wire n_946;
wire n_1539;
wire n_1001;
wire n_1503;
wire n_2054;
wire n_498;
wire n_1468;
wire n_1559;
wire n_1765;
wire n_1866;
wire n_689;
wire n_738;
wire n_1624;
wire n_640;
wire n_1510;
wire n_252;
wire n_624;
wire n_1380;
wire n_1744;
wire n_1617;
wire n_295;
wire n_1010;
wire n_1994;
wire n_1231;
wire n_739;
wire n_1279;
wire n_1406;
wire n_1195;
wire n_1839;
wire n_1837;
wire n_610;
wire n_1760;
wire n_936;
wire n_568;
wire n_1500;
wire n_1090;
wire n_757;
wire n_2342;
wire n_633;
wire n_439;
wire n_1832;
wire n_259;
wire n_448;
wire n_1851;
wire n_999;
wire n_758;
wire n_2046;
wire n_1933;
wire n_2290;
wire n_1656;
wire n_1158;
wire n_2045;
wire n_1509;
wire n_1874;
wire n_2040;
wire n_563;
wire n_2060;
wire n_1987;
wire n_1145;
wire n_878;
wire n_524;
wire n_394;
wire n_1678;
wire n_1049;
wire n_1153;
wire n_2145;
wire n_741;
wire n_1639;
wire n_1306;
wire n_1068;
wire n_1871;
wire n_1964;
wire n_331;
wire n_906;
wire n_1163;
wire n_2039;
wire n_1207;
wire n_919;
wire n_908;
wire n_2412;
wire n_2406;
wire n_724;
wire n_1781;
wire n_2084;
wire n_2035;
wire n_658;
wire n_2061;
wire n_2378;
wire n_1740;
wire n_2398;
wire n_1362;
wire n_1586;
wire n_456;
wire n_959;
wire n_535;
wire n_940;
wire n_1445;
wire n_1492;
wire n_2155;
wire n_1923;
wire n_1773;
wire n_592;
wire n_1169;
wire n_1692;
wire n_1596;
wire n_1017;
wire n_2171;
wire n_978;
wire n_2116;
wire n_2314;
wire n_1434;
wire n_1054;
wire n_1474;
wire n_1665;
wire n_1269;
wire n_2420;
wire n_1095;
wire n_1828;
wire n_1614;
wire n_267;
wire n_514;
wire n_1079;
wire n_457;
wire n_1045;
wire n_1208;
wire n_2093;
wire n_2038;
wire n_2320;
wire n_2339;
wire n_2137;
wire n_603;
wire n_1431;
wire n_484;
wire n_1593;
wire n_1033;
wire n_442;
wire n_2299;
wire n_636;
wire n_660;
wire n_2087;
wire n_1640;
wire n_2162;
wire n_1732;
wire n_1009;
wire n_1148;
wire n_2051;
wire n_750;
wire n_742;
wire n_2029;
wire n_995;
wire n_454;
wire n_2168;
wire n_1609;
wire n_374;
wire n_1989;
wire n_2359;
wire n_396;
wire n_1887;
wire n_1383;
wire n_1073;
wire n_255;
wire n_2346;
wire n_662;
wire n_459;
wire n_2312;
wire n_962;
wire n_1215;
wire n_1171;
wire n_1578;
wire n_723;
wire n_1920;
wire n_1065;
wire n_1592;
wire n_1336;
wire n_1721;
wire n_1959;
wire n_1758;
wire n_2338;
wire n_1574;
wire n_2399;
wire n_473;
wire n_2048;
wire n_2355;
wire n_2133;
wire n_1921;
wire n_1309;
wire n_1878;
wire n_1426;
wire n_1043;
wire n_355;
wire n_486;
wire n_1800;
wire n_1548;
wire n_614;
wire n_337;
wire n_1421;
wire n_1286;
wire n_1177;
wire n_1355;
wire n_974;
wire n_727;
wire n_1159;
wire n_957;
wire n_773;
wire n_2124;
wire n_743;
wire n_2081;
wire n_299;
wire n_303;
wire n_296;
wire n_613;
wire n_1119;
wire n_2156;
wire n_1240;
wire n_2261;
wire n_1820;
wire n_2418;
wire n_829;
wire n_1612;
wire n_2179;
wire n_1416;
wire n_2077;
wire n_1724;
wire n_2111;
wire n_361;
wire n_1237;
wire n_700;
wire n_573;
wire n_1420;
wire n_1132;
wire n_388;
wire n_1366;
wire n_1300;
wire n_1127;
wire n_2277;
wire n_761;
wire n_1785;
wire n_1568;
wire n_1006;
wire n_2110;
wire n_329;
wire n_274;
wire n_1270;
wire n_1664;
wire n_1486;
wire n_582;
wire n_1332;
wire n_2231;
wire n_1390;
wire n_2017;
wire n_2090;
wire n_1870;
wire n_309;
wire n_512;
wire n_2367;
wire n_1591;
wire n_2033;
wire n_322;
wire n_1682;
wire n_1980;
wire n_2390;
wire n_1249;
wire n_652;
wire n_1111;
wire n_1365;
wire n_1927;
wire n_2132;
wire n_1349;
wire n_1093;
wire n_288;
wire n_2400;
wire n_1031;
wire n_263;
wire n_609;
wire n_1041;
wire n_1265;
wire n_1909;
wire n_1562;
wire n_383;
wire n_834;
wire n_765;
wire n_2255;
wire n_2424;
wire n_2272;
wire n_893;
wire n_1015;
wire n_1140;
wire n_891;
wire n_1651;
wire n_1965;
wire n_239;
wire n_630;
wire n_1902;
wire n_2151;
wire n_1941;
wire n_2106;
wire n_1913;
wire n_504;
wire n_1823;
wire n_511;
wire n_874;
wire n_358;
wire n_1101;
wire n_1106;
wire n_1456;
wire n_2230;
wire n_2015;
wire n_2365;
wire n_1875;
wire n_1982;
wire n_1304;
wire n_1324;
wire n_987;
wire n_1846;
wire n_261;
wire n_2066;
wire n_1885;
wire n_1455;
wire n_767;
wire n_993;
wire n_1903;
wire n_1407;
wire n_2452;
wire n_1551;
wire n_545;
wire n_441;
wire n_860;
wire n_450;
wire n_1805;
wire n_2176;
wire n_2204;
wire n_1816;
wire n_429;
wire n_948;
wire n_1217;
wire n_2220;
wire n_2455;
wire n_628;
wire n_365;
wire n_1849;
wire n_2410;
wire n_729;
wire n_1131;
wire n_1084;
wire n_1961;
wire n_970;
wire n_1935;
wire n_911;
wire n_1430;
wire n_513;
wire n_1094;
wire n_1354;
wire n_560;
wire n_1534;
wire n_340;
wire n_2288;
wire n_1351;
wire n_2240;
wire n_1044;
wire n_1205;
wire n_2436;
wire n_346;
wire n_1209;
wire n_1552;
wire n_495;
wire n_602;
wire n_574;
wire n_1435;
wire n_879;
wire n_2416;
wire n_2405;
wire n_623;
wire n_2088;
wire n_405;
wire n_824;
wire n_359;
wire n_1645;
wire n_490;
wire n_1327;
wire n_2243;
wire n_996;
wire n_921;
wire n_1684;
wire n_1717;
wire n_572;
wire n_366;
wire n_815;
wire n_1795;
wire n_2128;
wire n_1821;
wire n_327;
wire n_1381;
wire n_1611;
wire n_1037;
wire n_2368;
wire n_1080;
wire n_2301;
wire n_1274;
wire n_1316;
wire n_1708;
wire n_2419;
wire n_426;
wire n_1438;
wire n_1082;
wire n_1840;
wire n_589;
wire n_716;
wire n_1630;
wire n_2122;
wire n_562;
wire n_1436;
wire n_1691;
wire n_952;
wire n_2092;
wire n_1229;
wire n_391;
wire n_701;
wire n_1437;
wire n_1023;
wire n_2075;
wire n_645;
wire n_539;
wire n_803;
wire n_1092;
wire n_1776;
wire n_2198;
wire n_2281;
wire n_2131;
wire n_2216;
wire n_531;
wire n_1757;
wire n_890;
wire n_1897;
wire n_764;
wire n_1919;
wire n_1056;
wire n_1424;
wire n_960;
wire n_2308;
wire n_1893;
wire n_1290;
wire n_1123;
wire n_1467;
wire n_1047;
wire n_2053;
wire n_2163;
wire n_634;
wire n_2328;
wire n_1958;
wire n_2254;
wire n_1252;
wire n_348;
wire n_1382;
wire n_1029;
wire n_925;
wire n_1206;
wire n_424;
wire n_1311;
wire n_2191;
wire n_1519;
wire n_256;
wire n_950;
wire n_2428;
wire n_1553;
wire n_1811;
wire n_2443;
wire n_380;
wire n_419;
wire n_1346;
wire n_444;
wire n_1299;
wire n_2158;
wire n_1808;
wire n_1060;
wire n_1141;
wire n_316;
wire n_2266;
wire n_389;
wire n_418;
wire n_248;
wire n_912;
wire n_315;
wire n_968;
wire n_451;
wire n_619;
wire n_408;
wire n_2440;
wire n_1386;
wire n_1699;
wire n_376;
wire n_967;
wire n_1442;
wire n_1139;
wire n_515;
wire n_2333;
wire n_351;
wire n_885;
wire n_397;
wire n_1432;
wire n_1357;
wire n_483;
wire n_2125;
wire n_683;
wire n_1632;
wire n_1057;
wire n_1051;
wire n_1085;
wire n_1066;
wire n_721;
wire n_2402;
wire n_1157;
wire n_2403;
wire n_841;
wire n_1050;
wire n_802;
wire n_1954;
wire n_2265;
wire n_1608;
wire n_983;
wire n_1844;
wire n_280;
wire n_1305;
wire n_873;
wire n_1826;
wire n_378;
wire n_1112;
wire n_2304;
wire n_762;
wire n_1283;
wire n_1644;
wire n_2334;
wire n_690;
wire n_1974;
wire n_583;
wire n_2086;
wire n_2289;
wire n_302;
wire n_1343;
wire n_2263;
wire n_1203;
wire n_1631;
wire n_821;
wire n_1763;
wire n_2341;
wire n_1966;
wire n_1768;
wire n_321;
wire n_2294;
wire n_1179;
wire n_621;
wire n_753;
wire n_455;
wire n_1048;
wire n_1719;
wire n_1288;
wire n_385;
wire n_507;
wire n_2269;
wire n_2309;
wire n_2415;
wire n_1560;
wire n_1605;
wire n_2236;
wire n_330;
wire n_1228;
wire n_2123;
wire n_972;
wire n_692;
wire n_2037;
wire n_1953;
wire n_1938;
wire n_820;
wire n_1200;
wire n_1911;
wire n_1363;
wire n_1301;
wire n_1668;
wire n_1185;
wire n_991;
wire n_828;
wire n_1967;
wire n_779;
wire n_576;
wire n_1143;
wire n_1579;
wire n_2233;
wire n_1329;
wire n_1312;
wire n_1439;
wire n_804;
wire n_537;
wire n_1688;
wire n_945;
wire n_492;
wire n_1504;
wire n_943;
wire n_341;
wire n_250;
wire n_992;
wire n_1932;
wire n_543;
wire n_260;
wire n_842;
wire n_650;
wire n_984;
wire n_694;
wire n_2082;
wire n_286;
wire n_1992;
wire n_2429;
wire n_1643;
wire n_883;
wire n_1983;
wire n_470;
wire n_325;
wire n_449;
wire n_1594;
wire n_1214;
wire n_1342;
wire n_1400;
wire n_900;
wire n_2362;
wire n_856;
wire n_1793;
wire n_1976;
wire n_2223;
wire n_918;
wire n_942;
wire n_2169;
wire n_1804;
wire n_1147;
wire n_1557;
wire n_1977;
wire n_2153;
wire n_1610;
wire n_1077;
wire n_1422;
wire n_2364;
wire n_540;
wire n_618;
wire n_896;
wire n_2310;
wire n_323;
wire n_2287;
wire n_356;
wire n_2291;
wire n_894;
wire n_1636;
wire n_2056;
wire n_1730;
wire n_831;
wire n_2280;
wire n_2192;
wire n_964;
wire n_1373;
wire n_1350;
wire n_1511;
wire n_1865;
wire n_1470;
wire n_1096;
wire n_2094;
wire n_1575;
wire n_1697;
wire n_1735;
wire n_833;
wire n_2318;
wire n_2393;
wire n_2020;
wire n_1646;
wire n_1307;
wire n_1881;
wire n_988;
wire n_2043;
wire n_1940;
wire n_814;
wire n_1549;
wire n_1934;
wire n_2311;
wire n_1201;
wire n_1114;
wire n_655;
wire n_2025;
wire n_1616;
wire n_1446;
wire n_2285;
wire n_669;
wire n_472;
wire n_1458;
wire n_1176;
wire n_1472;
wire n_2298;
wire n_1807;
wire n_387;
wire n_1149;
wire n_398;
wire n_1671;
wire n_635;
wire n_763;
wire n_1020;
wire n_1062;
wire n_2303;
wire n_1824;
wire n_1917;
wire n_2295;
wire n_1219;
wire n_1204;
wire n_2325;
wire n_2446;
wire n_1814;
wire n_1035;
wire n_287;
wire n_555;
wire n_783;
wire n_1928;
wire n_1848;
wire n_2126;
wire n_1188;
wire n_1722;
wire n_661;
wire n_2441;
wire n_1802;
wire n_849;
wire n_584;
wire n_681;
wire n_336;
wire n_1638;
wire n_1786;
wire n_430;
wire n_2002;
wire n_2282;
wire n_510;
wire n_2371;
wire n_311;
wire n_830;
wire n_2098;
wire n_1296;
wire n_2352;
wire n_1413;
wire n_801;
wire n_2207;
wire n_2080;
wire n_2377;
wire n_2340;
wire n_2444;
wire n_2068;
wire n_241;
wire n_875;
wire n_357;
wire n_1110;
wire n_1655;
wire n_445;
wire n_749;
wire n_1895;
wire n_1134;
wire n_1358;
wire n_717;
wire n_939;
wire n_482;
wire n_2361;
wire n_1088;
wire n_588;
wire n_1173;
wire n_789;
wire n_1232;
wire n_1603;
wire n_734;
wire n_638;
wire n_866;
wire n_969;
wire n_1401;
wire n_1019;
wire n_1105;
wire n_249;
wire n_1998;
wire n_304;
wire n_1338;
wire n_577;
wire n_2016;
wire n_1522;
wire n_1687;
wire n_1637;
wire n_2034;
wire n_1419;
wire n_338;
wire n_1653;
wire n_693;
wire n_2270;
wire n_1506;
wire n_990;
wire n_836;
wire n_1886;
wire n_1389;
wire n_1894;
wire n_975;
wire n_1908;
wire n_1256;
wire n_1702;
wire n_2259;
wire n_567;
wire n_1465;
wire n_778;
wire n_1122;
wire n_306;
wire n_458;
wire n_770;
wire n_1375;
wire n_1102;
wire n_2392;
wire n_1843;
wire n_711;
wire n_1499;
wire n_1187;
wire n_1441;
wire n_2435;
wire n_1392;
wire n_1597;
wire n_1929;
wire n_1164;
wire n_1659;
wire n_1834;
wire n_2097;
wire n_2313;
wire n_489;
wire n_1174;
wire n_2431;
wire n_1371;
wire n_617;
wire n_1303;
wire n_2206;
wire n_2063;
wire n_1572;
wire n_1968;
wire n_2252;
wire n_876;
wire n_1516;
wire n_1190;
wire n_1736;
wire n_1685;
wire n_2409;
wire n_601;
wire n_917;
wire n_1714;
wire n_966;
wire n_253;
wire n_1116;
wire n_2000;
wire n_1661;
wire n_1212;
wire n_2074;
wire n_1541;
wire n_726;
wire n_982;
wire n_1573;
wire n_1453;
wire n_1731;
wire n_2217;
wire n_818;
wire n_2373;
wire n_1970;
wire n_861;
wire n_1713;
wire n_1183;
wire n_2307;
wire n_1658;
wire n_899;
wire n_1253;
wire n_1737;
wire n_2201;
wire n_2117;
wire n_1904;
wire n_1993;
wire n_774;
wire n_1628;
wire n_2205;
wire n_1335;
wire n_1514;
wire n_1777;
wire n_1957;
wire n_1059;
wire n_1345;
wire n_1133;
wire n_1771;
wire n_1912;
wire n_1899;
wire n_557;
wire n_1410;
wire n_1005;
wire n_607;
wire n_1003;
wire n_679;
wire n_710;
wire n_2067;
wire n_527;
wire n_707;
wire n_1168;
wire n_2219;
wire n_2437;
wire n_2148;
wire n_937;
wire n_2445;
wire n_1427;
wire n_393;
wire n_487;
wire n_1726;
wire n_665;
wire n_1584;
wire n_1835;
wire n_1440;
wire n_2164;
wire n_421;
wire n_1988;
wire n_2115;
wire n_1853;
wire n_1356;
wire n_1787;
wire n_910;
wire n_2232;
wire n_2212;
wire n_1657;
wire n_768;
wire n_1475;
wire n_1302;
wire n_1774;
wire n_1725;
wire n_1136;
wire n_1313;
wire n_1491;
wire n_754;
wire n_1496;
wire n_1125;
wire n_410;
wire n_708;
wire n_529;
wire n_1812;
wire n_735;
wire n_1915;
wire n_1109;
wire n_895;
wire n_1310;
wire n_2121;
wire n_1803;
wire n_427;
wire n_1399;
wire n_1543;
wire n_1991;
wire n_1979;
wire n_791;
wire n_732;
wire n_1533;
wire n_2224;
wire n_808;
wire n_797;
wire n_1025;
wire n_1930;
wire n_1955;
wire n_500;
wire n_1067;
wire n_1720;
wire n_2401;
wire n_435;
wire n_2003;
wire n_766;
wire n_1457;
wire n_541;
wire n_538;
wire n_2354;
wire n_2246;
wire n_2008;
wire n_1117;
wire n_799;
wire n_2264;
wire n_687;
wire n_715;
wire n_1742;
wire n_1480;
wire n_1482;
wire n_1213;
wire n_1266;
wire n_536;
wire n_872;
wire n_2012;
wire n_594;
wire n_1291;
wire n_1297;
wire n_1753;
wire n_2283;
wire n_1782;
wire n_2245;
wire n_1155;
wire n_1418;
wire n_1972;
wire n_1524;
wire n_1689;
wire n_1485;
wire n_1011;
wire n_1184;
wire n_2184;
wire n_985;
wire n_1855;
wire n_2425;
wire n_869;
wire n_810;
wire n_416;
wire n_827;
wire n_401;
wire n_1703;
wire n_1352;
wire n_626;
wire n_2197;
wire n_2199;
wire n_1650;
wire n_1144;
wire n_1137;
wire n_1570;
wire n_1170;
wire n_305;
wire n_2023;
wire n_2213;
wire n_2351;
wire n_2211;
wire n_2095;
wire n_676;
wire n_294;
wire n_318;
wire n_2103;
wire n_653;
wire n_2160;
wire n_642;
wire n_2228;
wire n_1602;
wire n_855;
wire n_1178;
wire n_1461;
wire n_850;
wire n_684;
wire n_268;
wire n_2421;
wire n_2286;
wire n_664;
wire n_1999;
wire n_503;
wire n_2372;
wire n_2065;
wire n_2136;
wire n_1372;
wire n_605;
wire n_1273;
wire n_1822;
wire n_353;
wire n_620;
wire n_643;
wire n_2363;
wire n_2430;
wire n_916;
wire n_1081;
wire n_493;
wire n_2332;
wire n_1235;
wire n_703;
wire n_698;
wire n_980;
wire n_1115;
wire n_2433;
wire n_1282;
wire n_1318;
wire n_1783;
wire n_780;
wire n_998;
wire n_2375;
wire n_1454;
wire n_467;
wire n_1227;
wire n_1531;
wire n_840;
wire n_1334;
wire n_1907;
wire n_501;
wire n_823;
wire n_245;
wire n_725;
wire n_2344;
wire n_1388;
wire n_1417;
wire n_1295;
wire n_2316;
wire n_672;
wire n_1985;
wire n_1898;
wire n_2107;
wire n_581;
wire n_382;
wire n_554;
wire n_1625;
wire n_2130;
wire n_2187;
wire n_2284;
wire n_898;
wire n_1762;
wire n_1013;
wire n_1452;
wire n_718;
wire n_265;
wire n_1120;
wire n_719;
wire n_443;
wire n_1791;
wire n_1890;
wire n_1747;
wire n_714;
wire n_1683;
wire n_1944;
wire n_909;
wire n_1817;
wire n_1497;
wire n_1530;
wire n_997;
wire n_932;
wire n_612;
wire n_2078;
wire n_1409;
wire n_788;
wire n_1326;
wire n_1268;
wire n_559;
wire n_825;
wire n_1981;
wire n_508;
wire n_2186;
wire n_506;
wire n_1320;
wire n_1663;
wire n_737;
wire n_1718;
wire n_986;
wire n_2315;
wire n_509;
wire n_1317;
wire n_1518;
wire n_1715;
wire n_2102;
wire n_1281;
wire n_1952;
wire n_1192;
wire n_2221;
wire n_1024;
wire n_1063;
wire n_1889;
wire n_1792;
wire n_1564;
wire n_1868;
wire n_1613;
wire n_733;
wire n_1489;
wire n_1922;
wire n_1376;
wire n_941;
wire n_2326;
wire n_981;
wire n_1569;
wire n_2188;
wire n_867;
wire n_2348;
wire n_2422;
wire n_2239;
wire n_587;
wire n_792;
wire n_756;
wire n_1429;
wire n_399;
wire n_1238;
wire n_2448;
wire n_548;
wire n_812;
wire n_298;
wire n_2104;
wire n_518;
wire n_505;
wire n_2057;
wire n_1772;
wire n_282;
wire n_752;
wire n_905;
wire n_1476;
wire n_1108;
wire n_782;
wire n_1100;
wire n_1861;
wire n_2129;
wire n_1395;
wire n_862;
wire n_1425;
wire n_760;
wire n_1901;
wire n_1900;
wire n_1620;
wire n_381;
wire n_390;
wire n_1330;
wire n_1867;
wire n_1945;
wire n_481;
wire n_1675;
wire n_1924;
wire n_1727;
wire n_1554;
wire n_1745;
wire n_769;
wire n_2006;
wire n_1995;
wire n_2411;
wire n_2138;
wire n_1046;
wire n_271;
wire n_934;
wire n_1618;
wire n_2260;
wire n_826;
wire n_2343;
wire n_1813;
wire n_2447;
wire n_886;
wire n_2014;
wire n_1221;
wire n_2345;
wire n_654;
wire n_1172;
wire n_379;
wire n_428;
wire n_1341;
wire n_570;
wire n_1641;
wire n_1361;
wire n_2382;
wire n_1707;
wire n_853;
wire n_377;
wire n_2317;
wire n_751;
wire n_2172;
wire n_1973;
wire n_786;
wire n_1083;
wire n_1142;
wire n_2376;
wire n_1129;
wire n_392;
wire n_704;
wire n_787;
wire n_1770;
wire n_2456;
wire n_961;
wire n_2250;
wire n_1756;
wire n_771;
wire n_276;
wire n_1716;
wire n_1225;
wire n_1520;
wire n_2451;
wire n_522;
wire n_1287;
wire n_1262;
wire n_400;
wire n_930;
wire n_1873;
wire n_1411;
wire n_622;
wire n_1962;
wire n_1577;
wire n_2423;
wire n_1087;
wire n_386;
wire n_994;
wire n_1701;
wire n_2194;
wire n_848;
wire n_1550;
wire n_1498;
wire n_2167;
wire n_1223;
wire n_1272;
wire n_682;
wire n_1567;
wire n_1247;
wire n_922;
wire n_816;
wire n_1648;
wire n_591;
wire n_1536;
wire n_1857;
wire n_1344;
wire n_2041;
wire n_313;
wire n_631;
wire n_479;
wire n_1246;
wire n_1339;
wire n_1478;
wire n_1797;
wire n_432;
wire n_1769;
wire n_839;
wire n_1210;
wire n_1364;
wire n_2357;
wire n_2183;
wire n_2360;
wire n_328;
wire n_2292;
wire n_1250;
wire n_2173;
wire n_369;
wire n_1842;
wire n_871;
wire n_2442;
wire n_598;
wire n_685;
wire n_608;
wire n_928;
wire n_1367;
wire n_1943;
wire n_1460;
wire n_772;
wire n_2018;
wire n_1555;
wire n_499;
wire n_1589;
wire n_517;
wire n_402;
wire n_413;
wire n_1086;
wire n_796;
wire n_1858;
wire n_1619;
wire n_2119;
wire n_1502;
wire n_2157;
wire n_1469;
wire n_1012;
wire n_1396;
wire n_1348;
wire n_2030;
wire n_903;
wire n_2453;
wire n_1525;
wire n_1752;
wire n_2397;
wire n_740;
wire n_384;
wire n_2208;
wire n_1404;
wire n_1794;
wire n_2182;
wire n_1315;
wire n_2234;
wire n_277;
wire n_1061;
wire n_1910;
wire n_333;
wire n_1298;
wire n_1652;
wire n_2209;
wire n_462;
wire n_2050;
wire n_1193;
wire n_1676;
wire n_1255;
wire n_258;
wire n_1113;
wire n_2321;
wire n_1226;
wire n_722;
wire n_1277;
wire n_2146;
wire n_844;
wire n_471;
wire n_852;
wire n_1487;
wire n_1864;
wire n_1028;
wire n_1601;
wire n_781;
wire n_474;
wire n_542;
wire n_463;
wire n_1546;
wire n_595;
wire n_502;
wire n_466;
wire n_1337;
wire n_420;
wire n_1495;
wire n_632;
wire n_699;
wire n_979;
wire n_1515;
wire n_1627;
wire n_1245;
wire n_846;
wire n_2427;
wire n_2438;
wire n_1673;
wire n_465;
wire n_362;
wire n_1321;
wire n_1975;
wire n_2296;
wire n_2070;
wire n_273;
wire n_1937;
wire n_585;
wire n_2112;
wire n_1739;
wire n_270;
wire n_616;
wire n_2278;
wire n_2394;
wire n_1914;
wire n_2135;
wire n_2335;
wire n_745;
wire n_2381;
wire n_1654;
wire n_2349;
wire n_1103;
wire n_648;
wire n_1379;
wire n_312;
wire n_2196;
wire n_2170;
wire n_1076;
wire n_1091;
wire n_1408;
wire n_494;
wire n_1761;
wire n_641;
wire n_730;
wire n_2036;
wire n_1325;
wire n_1595;
wire n_2161;
wire n_354;
wire n_575;
wire n_480;
wire n_425;
wire n_795;
wire n_2404;
wire n_2083;
wire n_695;
wire n_656;
wire n_1606;
wire n_1220;
wire n_1694;
wire n_1540;
wire n_1936;
wire n_1956;
wire n_437;
wire n_1642;
wire n_2279;
wire n_2027;
wire n_453;
wire n_403;
wire n_1130;
wire n_720;
wire n_2366;
wire n_1918;
wire n_1526;
wire n_863;
wire n_2210;
wire n_805;
wire n_1604;
wire n_1275;
wire n_1764;
wire n_712;
wire n_2414;
wire n_246;
wire n_1583;
wire n_2426;
wire n_1042;
wire n_1402;
wire n_269;
wire n_2049;
wire n_2273;
wire n_285;
wire n_412;
wire n_1493;
wire n_657;
wire n_644;
wire n_1741;
wire n_2229;
wire n_1160;
wire n_1397;
wire n_491;
wire n_1258;
wire n_1074;
wire n_2004;
wire n_1621;
wire n_2113;
wire n_251;
wire n_566;
wire n_565;
wire n_1448;
wire n_2225;
wire n_1507;
wire n_1398;
wire n_2383;
wire n_1879;
wire n_597;
wire n_1996;
wire n_1181;
wire n_1505;
wire n_1634;
wire n_1196;
wire n_2019;
wire n_651;
wire n_1340;
wire n_2274;
wire n_334;
wire n_811;
wire n_1558;
wire n_807;
wire n_2166;
wire n_835;
wire n_666;
wire n_262;
wire n_1433;
wire n_1704;
wire n_2256;
wire n_1254;
wire n_1026;
wire n_2026;
wire n_1969;
wire n_1234;
wire n_2109;
wire n_319;
wire n_364;
wire n_1138;
wire n_927;
wire n_1089;
wire n_2044;
wire n_1990;
wire n_2013;
wire n_1004;
wire n_1186;
wire n_242;
wire n_1032;
wire n_1681;
wire n_2010;
wire n_1018;
wire n_2242;
wire n_2247;
wire n_1693;
wire n_438;
wire n_713;
wire n_904;
wire n_1588;
wire n_1622;
wire n_2237;
wire n_1180;
wire n_1827;
wire n_1271;
wire n_533;
wire n_1542;
wire n_1251;
wire n_278;
wire n_2268;

CKINVDCx5p33_ASAP7_75t_R g239 ( 
.A(n_30),
.Y(n_239)
);

INVx2_ASAP7_75t_L g240 ( 
.A(n_148),
.Y(n_240)
);

CKINVDCx5p33_ASAP7_75t_R g241 ( 
.A(n_101),
.Y(n_241)
);

CKINVDCx5p33_ASAP7_75t_R g242 ( 
.A(n_76),
.Y(n_242)
);

INVxp67_ASAP7_75t_L g243 ( 
.A(n_214),
.Y(n_243)
);

CKINVDCx5p33_ASAP7_75t_R g244 ( 
.A(n_77),
.Y(n_244)
);

CKINVDCx5p33_ASAP7_75t_R g245 ( 
.A(n_176),
.Y(n_245)
);

CKINVDCx5p33_ASAP7_75t_R g246 ( 
.A(n_13),
.Y(n_246)
);

CKINVDCx5p33_ASAP7_75t_R g247 ( 
.A(n_86),
.Y(n_247)
);

CKINVDCx5p33_ASAP7_75t_R g248 ( 
.A(n_61),
.Y(n_248)
);

CKINVDCx5p33_ASAP7_75t_R g249 ( 
.A(n_67),
.Y(n_249)
);

CKINVDCx5p33_ASAP7_75t_R g250 ( 
.A(n_44),
.Y(n_250)
);

CKINVDCx20_ASAP7_75t_R g251 ( 
.A(n_233),
.Y(n_251)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_189),
.Y(n_252)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_81),
.Y(n_253)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_89),
.Y(n_254)
);

CKINVDCx5p33_ASAP7_75t_R g255 ( 
.A(n_75),
.Y(n_255)
);

INVx2_ASAP7_75t_L g256 ( 
.A(n_48),
.Y(n_256)
);

CKINVDCx5p33_ASAP7_75t_R g257 ( 
.A(n_74),
.Y(n_257)
);

INVx2_ASAP7_75t_L g258 ( 
.A(n_49),
.Y(n_258)
);

INVx1_ASAP7_75t_SL g259 ( 
.A(n_200),
.Y(n_259)
);

CKINVDCx5p33_ASAP7_75t_R g260 ( 
.A(n_167),
.Y(n_260)
);

CKINVDCx20_ASAP7_75t_R g261 ( 
.A(n_74),
.Y(n_261)
);

CKINVDCx5p33_ASAP7_75t_R g262 ( 
.A(n_57),
.Y(n_262)
);

CKINVDCx20_ASAP7_75t_R g263 ( 
.A(n_115),
.Y(n_263)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_88),
.Y(n_264)
);

BUFx3_ASAP7_75t_L g265 ( 
.A(n_199),
.Y(n_265)
);

BUFx3_ASAP7_75t_L g266 ( 
.A(n_99),
.Y(n_266)
);

CKINVDCx5p33_ASAP7_75t_R g267 ( 
.A(n_222),
.Y(n_267)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_92),
.Y(n_268)
);

INVx2_ASAP7_75t_SL g269 ( 
.A(n_146),
.Y(n_269)
);

CKINVDCx5p33_ASAP7_75t_R g270 ( 
.A(n_114),
.Y(n_270)
);

CKINVDCx5p33_ASAP7_75t_R g271 ( 
.A(n_82),
.Y(n_271)
);

CKINVDCx5p33_ASAP7_75t_R g272 ( 
.A(n_100),
.Y(n_272)
);

CKINVDCx5p33_ASAP7_75t_R g273 ( 
.A(n_72),
.Y(n_273)
);

CKINVDCx5p33_ASAP7_75t_R g274 ( 
.A(n_226),
.Y(n_274)
);

CKINVDCx5p33_ASAP7_75t_R g275 ( 
.A(n_73),
.Y(n_275)
);

CKINVDCx5p33_ASAP7_75t_R g276 ( 
.A(n_195),
.Y(n_276)
);

INVx2_ASAP7_75t_L g277 ( 
.A(n_180),
.Y(n_277)
);

CKINVDCx5p33_ASAP7_75t_R g278 ( 
.A(n_112),
.Y(n_278)
);

CKINVDCx5p33_ASAP7_75t_R g279 ( 
.A(n_53),
.Y(n_279)
);

INVx2_ASAP7_75t_L g280 ( 
.A(n_215),
.Y(n_280)
);

CKINVDCx5p33_ASAP7_75t_R g281 ( 
.A(n_196),
.Y(n_281)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_117),
.Y(n_282)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_143),
.Y(n_283)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_190),
.Y(n_284)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_11),
.Y(n_285)
);

CKINVDCx5p33_ASAP7_75t_R g286 ( 
.A(n_219),
.Y(n_286)
);

CKINVDCx5p33_ASAP7_75t_R g287 ( 
.A(n_47),
.Y(n_287)
);

CKINVDCx5p33_ASAP7_75t_R g288 ( 
.A(n_90),
.Y(n_288)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_70),
.Y(n_289)
);

INVx2_ASAP7_75t_L g290 ( 
.A(n_238),
.Y(n_290)
);

CKINVDCx5p33_ASAP7_75t_R g291 ( 
.A(n_72),
.Y(n_291)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_92),
.Y(n_292)
);

BUFx3_ASAP7_75t_L g293 ( 
.A(n_28),
.Y(n_293)
);

CKINVDCx5p33_ASAP7_75t_R g294 ( 
.A(n_79),
.Y(n_294)
);

CKINVDCx5p33_ASAP7_75t_R g295 ( 
.A(n_1),
.Y(n_295)
);

CKINVDCx20_ASAP7_75t_R g296 ( 
.A(n_40),
.Y(n_296)
);

CKINVDCx5p33_ASAP7_75t_R g297 ( 
.A(n_217),
.Y(n_297)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_168),
.Y(n_298)
);

CKINVDCx5p33_ASAP7_75t_R g299 ( 
.A(n_152),
.Y(n_299)
);

CKINVDCx5p33_ASAP7_75t_R g300 ( 
.A(n_194),
.Y(n_300)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_67),
.Y(n_301)
);

CKINVDCx5p33_ASAP7_75t_R g302 ( 
.A(n_166),
.Y(n_302)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_187),
.Y(n_303)
);

CKINVDCx5p33_ASAP7_75t_R g304 ( 
.A(n_51),
.Y(n_304)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_232),
.Y(n_305)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_93),
.Y(n_306)
);

CKINVDCx5p33_ASAP7_75t_R g307 ( 
.A(n_132),
.Y(n_307)
);

BUFx3_ASAP7_75t_L g308 ( 
.A(n_55),
.Y(n_308)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_31),
.Y(n_309)
);

CKINVDCx5p33_ASAP7_75t_R g310 ( 
.A(n_95),
.Y(n_310)
);

BUFx5_ASAP7_75t_L g311 ( 
.A(n_141),
.Y(n_311)
);

CKINVDCx5p33_ASAP7_75t_R g312 ( 
.A(n_0),
.Y(n_312)
);

INVx2_ASAP7_75t_L g313 ( 
.A(n_118),
.Y(n_313)
);

CKINVDCx5p33_ASAP7_75t_R g314 ( 
.A(n_42),
.Y(n_314)
);

CKINVDCx5p33_ASAP7_75t_R g315 ( 
.A(n_125),
.Y(n_315)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_174),
.Y(n_316)
);

CKINVDCx16_ASAP7_75t_R g317 ( 
.A(n_98),
.Y(n_317)
);

BUFx10_ASAP7_75t_L g318 ( 
.A(n_10),
.Y(n_318)
);

CKINVDCx5p33_ASAP7_75t_R g319 ( 
.A(n_133),
.Y(n_319)
);

CKINVDCx20_ASAP7_75t_R g320 ( 
.A(n_164),
.Y(n_320)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_136),
.Y(n_321)
);

CKINVDCx5p33_ASAP7_75t_R g322 ( 
.A(n_227),
.Y(n_322)
);

CKINVDCx5p33_ASAP7_75t_R g323 ( 
.A(n_49),
.Y(n_323)
);

BUFx2_ASAP7_75t_SL g324 ( 
.A(n_121),
.Y(n_324)
);

CKINVDCx5p33_ASAP7_75t_R g325 ( 
.A(n_25),
.Y(n_325)
);

CKINVDCx5p33_ASAP7_75t_R g326 ( 
.A(n_38),
.Y(n_326)
);

CKINVDCx5p33_ASAP7_75t_R g327 ( 
.A(n_140),
.Y(n_327)
);

CKINVDCx5p33_ASAP7_75t_R g328 ( 
.A(n_235),
.Y(n_328)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_216),
.Y(n_329)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_208),
.Y(n_330)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_188),
.Y(n_331)
);

CKINVDCx5p33_ASAP7_75t_R g332 ( 
.A(n_151),
.Y(n_332)
);

HB1xp67_ASAP7_75t_L g333 ( 
.A(n_32),
.Y(n_333)
);

BUFx2_ASAP7_75t_L g334 ( 
.A(n_129),
.Y(n_334)
);

CKINVDCx20_ASAP7_75t_R g335 ( 
.A(n_137),
.Y(n_335)
);

CKINVDCx5p33_ASAP7_75t_R g336 ( 
.A(n_69),
.Y(n_336)
);

CKINVDCx5p33_ASAP7_75t_R g337 ( 
.A(n_27),
.Y(n_337)
);

INVx2_ASAP7_75t_L g338 ( 
.A(n_183),
.Y(n_338)
);

CKINVDCx5p33_ASAP7_75t_R g339 ( 
.A(n_76),
.Y(n_339)
);

BUFx2_ASAP7_75t_L g340 ( 
.A(n_32),
.Y(n_340)
);

CKINVDCx5p33_ASAP7_75t_R g341 ( 
.A(n_191),
.Y(n_341)
);

CKINVDCx16_ASAP7_75t_R g342 ( 
.A(n_77),
.Y(n_342)
);

CKINVDCx5p33_ASAP7_75t_R g343 ( 
.A(n_16),
.Y(n_343)
);

INVx1_ASAP7_75t_L g344 ( 
.A(n_25),
.Y(n_344)
);

CKINVDCx5p33_ASAP7_75t_R g345 ( 
.A(n_171),
.Y(n_345)
);

INVx1_ASAP7_75t_L g346 ( 
.A(n_98),
.Y(n_346)
);

CKINVDCx5p33_ASAP7_75t_R g347 ( 
.A(n_48),
.Y(n_347)
);

CKINVDCx5p33_ASAP7_75t_R g348 ( 
.A(n_73),
.Y(n_348)
);

CKINVDCx5p33_ASAP7_75t_R g349 ( 
.A(n_229),
.Y(n_349)
);

CKINVDCx5p33_ASAP7_75t_R g350 ( 
.A(n_101),
.Y(n_350)
);

CKINVDCx5p33_ASAP7_75t_R g351 ( 
.A(n_102),
.Y(n_351)
);

CKINVDCx5p33_ASAP7_75t_R g352 ( 
.A(n_55),
.Y(n_352)
);

INVx1_ASAP7_75t_L g353 ( 
.A(n_126),
.Y(n_353)
);

CKINVDCx5p33_ASAP7_75t_R g354 ( 
.A(n_159),
.Y(n_354)
);

CKINVDCx5p33_ASAP7_75t_R g355 ( 
.A(n_175),
.Y(n_355)
);

INVx1_ASAP7_75t_L g356 ( 
.A(n_213),
.Y(n_356)
);

CKINVDCx5p33_ASAP7_75t_R g357 ( 
.A(n_17),
.Y(n_357)
);

BUFx10_ASAP7_75t_L g358 ( 
.A(n_157),
.Y(n_358)
);

INVx1_ASAP7_75t_L g359 ( 
.A(n_155),
.Y(n_359)
);

INVx1_ASAP7_75t_SL g360 ( 
.A(n_186),
.Y(n_360)
);

INVx1_ASAP7_75t_L g361 ( 
.A(n_6),
.Y(n_361)
);

CKINVDCx5p33_ASAP7_75t_R g362 ( 
.A(n_54),
.Y(n_362)
);

CKINVDCx20_ASAP7_75t_R g363 ( 
.A(n_30),
.Y(n_363)
);

INVx1_ASAP7_75t_L g364 ( 
.A(n_205),
.Y(n_364)
);

INVx1_ASAP7_75t_L g365 ( 
.A(n_149),
.Y(n_365)
);

CKINVDCx5p33_ASAP7_75t_R g366 ( 
.A(n_43),
.Y(n_366)
);

INVx1_ASAP7_75t_L g367 ( 
.A(n_211),
.Y(n_367)
);

CKINVDCx5p33_ASAP7_75t_R g368 ( 
.A(n_116),
.Y(n_368)
);

BUFx6f_ASAP7_75t_L g369 ( 
.A(n_64),
.Y(n_369)
);

CKINVDCx5p33_ASAP7_75t_R g370 ( 
.A(n_165),
.Y(n_370)
);

CKINVDCx5p33_ASAP7_75t_R g371 ( 
.A(n_94),
.Y(n_371)
);

CKINVDCx20_ASAP7_75t_R g372 ( 
.A(n_87),
.Y(n_372)
);

CKINVDCx5p33_ASAP7_75t_R g373 ( 
.A(n_120),
.Y(n_373)
);

CKINVDCx5p33_ASAP7_75t_R g374 ( 
.A(n_69),
.Y(n_374)
);

HB1xp67_ASAP7_75t_L g375 ( 
.A(n_78),
.Y(n_375)
);

CKINVDCx5p33_ASAP7_75t_R g376 ( 
.A(n_81),
.Y(n_376)
);

CKINVDCx5p33_ASAP7_75t_R g377 ( 
.A(n_225),
.Y(n_377)
);

INVx1_ASAP7_75t_L g378 ( 
.A(n_24),
.Y(n_378)
);

INVx1_ASAP7_75t_SL g379 ( 
.A(n_202),
.Y(n_379)
);

CKINVDCx5p33_ASAP7_75t_R g380 ( 
.A(n_10),
.Y(n_380)
);

INVx1_ASAP7_75t_L g381 ( 
.A(n_193),
.Y(n_381)
);

CKINVDCx5p33_ASAP7_75t_R g382 ( 
.A(n_109),
.Y(n_382)
);

CKINVDCx20_ASAP7_75t_R g383 ( 
.A(n_124),
.Y(n_383)
);

CKINVDCx5p33_ASAP7_75t_R g384 ( 
.A(n_197),
.Y(n_384)
);

CKINVDCx20_ASAP7_75t_R g385 ( 
.A(n_20),
.Y(n_385)
);

CKINVDCx5p33_ASAP7_75t_R g386 ( 
.A(n_128),
.Y(n_386)
);

BUFx6f_ASAP7_75t_L g387 ( 
.A(n_103),
.Y(n_387)
);

BUFx5_ASAP7_75t_L g388 ( 
.A(n_105),
.Y(n_388)
);

CKINVDCx5p33_ASAP7_75t_R g389 ( 
.A(n_8),
.Y(n_389)
);

CKINVDCx5p33_ASAP7_75t_R g390 ( 
.A(n_56),
.Y(n_390)
);

CKINVDCx5p33_ASAP7_75t_R g391 ( 
.A(n_236),
.Y(n_391)
);

CKINVDCx5p33_ASAP7_75t_R g392 ( 
.A(n_161),
.Y(n_392)
);

INVx2_ASAP7_75t_L g393 ( 
.A(n_147),
.Y(n_393)
);

CKINVDCx5p33_ASAP7_75t_R g394 ( 
.A(n_153),
.Y(n_394)
);

CKINVDCx5p33_ASAP7_75t_R g395 ( 
.A(n_11),
.Y(n_395)
);

INVx2_ASAP7_75t_L g396 ( 
.A(n_29),
.Y(n_396)
);

CKINVDCx5p33_ASAP7_75t_R g397 ( 
.A(n_119),
.Y(n_397)
);

CKINVDCx5p33_ASAP7_75t_R g398 ( 
.A(n_1),
.Y(n_398)
);

CKINVDCx5p33_ASAP7_75t_R g399 ( 
.A(n_95),
.Y(n_399)
);

INVx1_ASAP7_75t_L g400 ( 
.A(n_18),
.Y(n_400)
);

INVx1_ASAP7_75t_SL g401 ( 
.A(n_104),
.Y(n_401)
);

INVx1_ASAP7_75t_L g402 ( 
.A(n_163),
.Y(n_402)
);

INVx1_ASAP7_75t_L g403 ( 
.A(n_234),
.Y(n_403)
);

CKINVDCx5p33_ASAP7_75t_R g404 ( 
.A(n_31),
.Y(n_404)
);

CKINVDCx5p33_ASAP7_75t_R g405 ( 
.A(n_5),
.Y(n_405)
);

INVx2_ASAP7_75t_SL g406 ( 
.A(n_220),
.Y(n_406)
);

BUFx3_ASAP7_75t_L g407 ( 
.A(n_0),
.Y(n_407)
);

CKINVDCx5p33_ASAP7_75t_R g408 ( 
.A(n_71),
.Y(n_408)
);

INVx1_ASAP7_75t_L g409 ( 
.A(n_109),
.Y(n_409)
);

CKINVDCx5p33_ASAP7_75t_R g410 ( 
.A(n_169),
.Y(n_410)
);

CKINVDCx5p33_ASAP7_75t_R g411 ( 
.A(n_113),
.Y(n_411)
);

INVx1_ASAP7_75t_SL g412 ( 
.A(n_7),
.Y(n_412)
);

CKINVDCx5p33_ASAP7_75t_R g413 ( 
.A(n_54),
.Y(n_413)
);

INVx1_ASAP7_75t_L g414 ( 
.A(n_24),
.Y(n_414)
);

BUFx3_ASAP7_75t_L g415 ( 
.A(n_89),
.Y(n_415)
);

CKINVDCx5p33_ASAP7_75t_R g416 ( 
.A(n_23),
.Y(n_416)
);

CKINVDCx5p33_ASAP7_75t_R g417 ( 
.A(n_192),
.Y(n_417)
);

CKINVDCx20_ASAP7_75t_R g418 ( 
.A(n_78),
.Y(n_418)
);

CKINVDCx20_ASAP7_75t_R g419 ( 
.A(n_97),
.Y(n_419)
);

CKINVDCx5p33_ASAP7_75t_R g420 ( 
.A(n_41),
.Y(n_420)
);

CKINVDCx5p33_ASAP7_75t_R g421 ( 
.A(n_130),
.Y(n_421)
);

CKINVDCx5p33_ASAP7_75t_R g422 ( 
.A(n_123),
.Y(n_422)
);

CKINVDCx5p33_ASAP7_75t_R g423 ( 
.A(n_100),
.Y(n_423)
);

CKINVDCx5p33_ASAP7_75t_R g424 ( 
.A(n_6),
.Y(n_424)
);

INVx1_ASAP7_75t_L g425 ( 
.A(n_170),
.Y(n_425)
);

CKINVDCx5p33_ASAP7_75t_R g426 ( 
.A(n_37),
.Y(n_426)
);

INVx1_ASAP7_75t_L g427 ( 
.A(n_20),
.Y(n_427)
);

INVx1_ASAP7_75t_L g428 ( 
.A(n_162),
.Y(n_428)
);

INVx1_ASAP7_75t_L g429 ( 
.A(n_33),
.Y(n_429)
);

CKINVDCx5p33_ASAP7_75t_R g430 ( 
.A(n_90),
.Y(n_430)
);

INVx1_ASAP7_75t_L g431 ( 
.A(n_22),
.Y(n_431)
);

INVx1_ASAP7_75t_L g432 ( 
.A(n_13),
.Y(n_432)
);

INVx1_ASAP7_75t_L g433 ( 
.A(n_83),
.Y(n_433)
);

INVx1_ASAP7_75t_L g434 ( 
.A(n_68),
.Y(n_434)
);

CKINVDCx5p33_ASAP7_75t_R g435 ( 
.A(n_33),
.Y(n_435)
);

INVx1_ASAP7_75t_L g436 ( 
.A(n_182),
.Y(n_436)
);

HB1xp67_ASAP7_75t_L g437 ( 
.A(n_75),
.Y(n_437)
);

CKINVDCx5p33_ASAP7_75t_R g438 ( 
.A(n_223),
.Y(n_438)
);

INVx3_ASAP7_75t_L g439 ( 
.A(n_91),
.Y(n_439)
);

CKINVDCx5p33_ASAP7_75t_R g440 ( 
.A(n_178),
.Y(n_440)
);

CKINVDCx5p33_ASAP7_75t_R g441 ( 
.A(n_207),
.Y(n_441)
);

INVx2_ASAP7_75t_L g442 ( 
.A(n_36),
.Y(n_442)
);

CKINVDCx5p33_ASAP7_75t_R g443 ( 
.A(n_184),
.Y(n_443)
);

BUFx2_ASAP7_75t_SL g444 ( 
.A(n_41),
.Y(n_444)
);

CKINVDCx5p33_ASAP7_75t_R g445 ( 
.A(n_35),
.Y(n_445)
);

CKINVDCx5p33_ASAP7_75t_R g446 ( 
.A(n_210),
.Y(n_446)
);

CKINVDCx5p33_ASAP7_75t_R g447 ( 
.A(n_26),
.Y(n_447)
);

INVx1_ASAP7_75t_L g448 ( 
.A(n_7),
.Y(n_448)
);

CKINVDCx5p33_ASAP7_75t_R g449 ( 
.A(n_83),
.Y(n_449)
);

INVx2_ASAP7_75t_L g450 ( 
.A(n_91),
.Y(n_450)
);

CKINVDCx5p33_ASAP7_75t_R g451 ( 
.A(n_28),
.Y(n_451)
);

INVx3_ASAP7_75t_L g452 ( 
.A(n_16),
.Y(n_452)
);

CKINVDCx5p33_ASAP7_75t_R g453 ( 
.A(n_56),
.Y(n_453)
);

INVx1_ASAP7_75t_L g454 ( 
.A(n_110),
.Y(n_454)
);

BUFx3_ASAP7_75t_L g455 ( 
.A(n_70),
.Y(n_455)
);

CKINVDCx5p33_ASAP7_75t_R g456 ( 
.A(n_9),
.Y(n_456)
);

CKINVDCx5p33_ASAP7_75t_R g457 ( 
.A(n_37),
.Y(n_457)
);

INVx2_ASAP7_75t_L g458 ( 
.A(n_179),
.Y(n_458)
);

INVx1_ASAP7_75t_L g459 ( 
.A(n_110),
.Y(n_459)
);

INVx1_ASAP7_75t_L g460 ( 
.A(n_135),
.Y(n_460)
);

CKINVDCx5p33_ASAP7_75t_R g461 ( 
.A(n_106),
.Y(n_461)
);

CKINVDCx20_ASAP7_75t_R g462 ( 
.A(n_209),
.Y(n_462)
);

CKINVDCx5p33_ASAP7_75t_R g463 ( 
.A(n_38),
.Y(n_463)
);

CKINVDCx20_ASAP7_75t_R g464 ( 
.A(n_17),
.Y(n_464)
);

CKINVDCx5p33_ASAP7_75t_R g465 ( 
.A(n_111),
.Y(n_465)
);

INVx1_ASAP7_75t_L g466 ( 
.A(n_53),
.Y(n_466)
);

INVx1_ASAP7_75t_SL g467 ( 
.A(n_14),
.Y(n_467)
);

INVx1_ASAP7_75t_L g468 ( 
.A(n_122),
.Y(n_468)
);

CKINVDCx5p33_ASAP7_75t_R g469 ( 
.A(n_80),
.Y(n_469)
);

INVx1_ASAP7_75t_L g470 ( 
.A(n_154),
.Y(n_470)
);

INVx1_ASAP7_75t_L g471 ( 
.A(n_388),
.Y(n_471)
);

CKINVDCx20_ASAP7_75t_R g472 ( 
.A(n_251),
.Y(n_472)
);

INVx1_ASAP7_75t_L g473 ( 
.A(n_388),
.Y(n_473)
);

INVx1_ASAP7_75t_L g474 ( 
.A(n_388),
.Y(n_474)
);

CKINVDCx16_ASAP7_75t_R g475 ( 
.A(n_317),
.Y(n_475)
);

CKINVDCx5p33_ASAP7_75t_R g476 ( 
.A(n_245),
.Y(n_476)
);

INVx1_ASAP7_75t_L g477 ( 
.A(n_388),
.Y(n_477)
);

INVx1_ASAP7_75t_L g478 ( 
.A(n_388),
.Y(n_478)
);

BUFx2_ASAP7_75t_L g479 ( 
.A(n_340),
.Y(n_479)
);

CKINVDCx5p33_ASAP7_75t_R g480 ( 
.A(n_260),
.Y(n_480)
);

CKINVDCx20_ASAP7_75t_R g481 ( 
.A(n_263),
.Y(n_481)
);

INVxp67_ASAP7_75t_SL g482 ( 
.A(n_334),
.Y(n_482)
);

CKINVDCx5p33_ASAP7_75t_R g483 ( 
.A(n_267),
.Y(n_483)
);

NOR2xp33_ASAP7_75t_L g484 ( 
.A(n_334),
.B(n_2),
.Y(n_484)
);

INVxp67_ASAP7_75t_SL g485 ( 
.A(n_439),
.Y(n_485)
);

NOR2xp67_ASAP7_75t_L g486 ( 
.A(n_439),
.B(n_2),
.Y(n_486)
);

CKINVDCx5p33_ASAP7_75t_R g487 ( 
.A(n_270),
.Y(n_487)
);

INVx1_ASAP7_75t_L g488 ( 
.A(n_388),
.Y(n_488)
);

CKINVDCx20_ASAP7_75t_R g489 ( 
.A(n_320),
.Y(n_489)
);

INVx1_ASAP7_75t_L g490 ( 
.A(n_388),
.Y(n_490)
);

INVx1_ASAP7_75t_L g491 ( 
.A(n_388),
.Y(n_491)
);

INVx1_ASAP7_75t_L g492 ( 
.A(n_388),
.Y(n_492)
);

NOR2xp67_ASAP7_75t_L g493 ( 
.A(n_439),
.B(n_3),
.Y(n_493)
);

CKINVDCx20_ASAP7_75t_R g494 ( 
.A(n_462),
.Y(n_494)
);

INVx1_ASAP7_75t_L g495 ( 
.A(n_388),
.Y(n_495)
);

CKINVDCx20_ASAP7_75t_R g496 ( 
.A(n_335),
.Y(n_496)
);

INVx1_ASAP7_75t_L g497 ( 
.A(n_369),
.Y(n_497)
);

INVx1_ASAP7_75t_L g498 ( 
.A(n_369),
.Y(n_498)
);

INVx1_ASAP7_75t_L g499 ( 
.A(n_369),
.Y(n_499)
);

INVx1_ASAP7_75t_L g500 ( 
.A(n_369),
.Y(n_500)
);

INVx1_ASAP7_75t_L g501 ( 
.A(n_369),
.Y(n_501)
);

INVx1_ASAP7_75t_L g502 ( 
.A(n_369),
.Y(n_502)
);

INVx1_ASAP7_75t_L g503 ( 
.A(n_387),
.Y(n_503)
);

CKINVDCx20_ASAP7_75t_R g504 ( 
.A(n_335),
.Y(n_504)
);

INVx1_ASAP7_75t_L g505 ( 
.A(n_387),
.Y(n_505)
);

INVx1_ASAP7_75t_L g506 ( 
.A(n_387),
.Y(n_506)
);

INVx1_ASAP7_75t_L g507 ( 
.A(n_387),
.Y(n_507)
);

CKINVDCx5p33_ASAP7_75t_R g508 ( 
.A(n_274),
.Y(n_508)
);

INVx1_ASAP7_75t_L g509 ( 
.A(n_387),
.Y(n_509)
);

CKINVDCx5p33_ASAP7_75t_R g510 ( 
.A(n_276),
.Y(n_510)
);

CKINVDCx5p33_ASAP7_75t_R g511 ( 
.A(n_278),
.Y(n_511)
);

NOR2xp67_ASAP7_75t_L g512 ( 
.A(n_439),
.B(n_3),
.Y(n_512)
);

CKINVDCx5p33_ASAP7_75t_R g513 ( 
.A(n_281),
.Y(n_513)
);

CKINVDCx16_ASAP7_75t_R g514 ( 
.A(n_317),
.Y(n_514)
);

CKINVDCx20_ASAP7_75t_R g515 ( 
.A(n_383),
.Y(n_515)
);

OR2x2_ASAP7_75t_L g516 ( 
.A(n_253),
.B(n_4),
.Y(n_516)
);

INVxp33_ASAP7_75t_SL g517 ( 
.A(n_333),
.Y(n_517)
);

INVx1_ASAP7_75t_L g518 ( 
.A(n_387),
.Y(n_518)
);

INVxp67_ASAP7_75t_L g519 ( 
.A(n_333),
.Y(n_519)
);

CKINVDCx5p33_ASAP7_75t_R g520 ( 
.A(n_286),
.Y(n_520)
);

CKINVDCx5p33_ASAP7_75t_R g521 ( 
.A(n_297),
.Y(n_521)
);

CKINVDCx5p33_ASAP7_75t_R g522 ( 
.A(n_299),
.Y(n_522)
);

INVx1_ASAP7_75t_L g523 ( 
.A(n_452),
.Y(n_523)
);

INVx1_ASAP7_75t_L g524 ( 
.A(n_252),
.Y(n_524)
);

CKINVDCx20_ASAP7_75t_R g525 ( 
.A(n_383),
.Y(n_525)
);

CKINVDCx5p33_ASAP7_75t_R g526 ( 
.A(n_300),
.Y(n_526)
);

INVx1_ASAP7_75t_L g527 ( 
.A(n_452),
.Y(n_527)
);

INVx1_ASAP7_75t_L g528 ( 
.A(n_452),
.Y(n_528)
);

BUFx2_ASAP7_75t_L g529 ( 
.A(n_340),
.Y(n_529)
);

INVx1_ASAP7_75t_L g530 ( 
.A(n_452),
.Y(n_530)
);

NOR2xp33_ASAP7_75t_L g531 ( 
.A(n_243),
.B(n_4),
.Y(n_531)
);

CKINVDCx5p33_ASAP7_75t_R g532 ( 
.A(n_302),
.Y(n_532)
);

INVx1_ASAP7_75t_L g533 ( 
.A(n_256),
.Y(n_533)
);

CKINVDCx20_ASAP7_75t_R g534 ( 
.A(n_307),
.Y(n_534)
);

CKINVDCx20_ASAP7_75t_R g535 ( 
.A(n_315),
.Y(n_535)
);

CKINVDCx5p33_ASAP7_75t_R g536 ( 
.A(n_319),
.Y(n_536)
);

CKINVDCx20_ASAP7_75t_R g537 ( 
.A(n_322),
.Y(n_537)
);

CKINVDCx5p33_ASAP7_75t_R g538 ( 
.A(n_327),
.Y(n_538)
);

INVx1_ASAP7_75t_L g539 ( 
.A(n_256),
.Y(n_539)
);

CKINVDCx5p33_ASAP7_75t_R g540 ( 
.A(n_328),
.Y(n_540)
);

INVx1_ASAP7_75t_L g541 ( 
.A(n_256),
.Y(n_541)
);

INVx1_ASAP7_75t_L g542 ( 
.A(n_258),
.Y(n_542)
);

INVx1_ASAP7_75t_L g543 ( 
.A(n_258),
.Y(n_543)
);

NOR2xp33_ASAP7_75t_L g544 ( 
.A(n_243),
.B(n_5),
.Y(n_544)
);

CKINVDCx5p33_ASAP7_75t_R g545 ( 
.A(n_332),
.Y(n_545)
);

NOR2xp33_ASAP7_75t_L g546 ( 
.A(n_269),
.B(n_8),
.Y(n_546)
);

CKINVDCx5p33_ASAP7_75t_R g547 ( 
.A(n_341),
.Y(n_547)
);

NOR2xp33_ASAP7_75t_L g548 ( 
.A(n_269),
.B(n_9),
.Y(n_548)
);

INVxp67_ASAP7_75t_SL g549 ( 
.A(n_265),
.Y(n_549)
);

INVx1_ASAP7_75t_L g550 ( 
.A(n_258),
.Y(n_550)
);

CKINVDCx5p33_ASAP7_75t_R g551 ( 
.A(n_345),
.Y(n_551)
);

CKINVDCx5p33_ASAP7_75t_R g552 ( 
.A(n_349),
.Y(n_552)
);

INVx1_ASAP7_75t_L g553 ( 
.A(n_396),
.Y(n_553)
);

CKINVDCx5p33_ASAP7_75t_R g554 ( 
.A(n_354),
.Y(n_554)
);

CKINVDCx5p33_ASAP7_75t_R g555 ( 
.A(n_355),
.Y(n_555)
);

INVxp67_ASAP7_75t_L g556 ( 
.A(n_375),
.Y(n_556)
);

INVx1_ASAP7_75t_L g557 ( 
.A(n_396),
.Y(n_557)
);

CKINVDCx16_ASAP7_75t_R g558 ( 
.A(n_342),
.Y(n_558)
);

CKINVDCx5p33_ASAP7_75t_R g559 ( 
.A(n_368),
.Y(n_559)
);

CKINVDCx20_ASAP7_75t_R g560 ( 
.A(n_370),
.Y(n_560)
);

INVx1_ASAP7_75t_L g561 ( 
.A(n_396),
.Y(n_561)
);

INVx1_ASAP7_75t_L g562 ( 
.A(n_442),
.Y(n_562)
);

INVx1_ASAP7_75t_L g563 ( 
.A(n_442),
.Y(n_563)
);

CKINVDCx20_ASAP7_75t_R g564 ( 
.A(n_373),
.Y(n_564)
);

CKINVDCx5p33_ASAP7_75t_R g565 ( 
.A(n_377),
.Y(n_565)
);

INVx1_ASAP7_75t_L g566 ( 
.A(n_442),
.Y(n_566)
);

CKINVDCx5p33_ASAP7_75t_R g567 ( 
.A(n_384),
.Y(n_567)
);

INVx1_ASAP7_75t_L g568 ( 
.A(n_450),
.Y(n_568)
);

BUFx3_ASAP7_75t_L g569 ( 
.A(n_265),
.Y(n_569)
);

INVx1_ASAP7_75t_L g570 ( 
.A(n_450),
.Y(n_570)
);

INVx1_ASAP7_75t_L g571 ( 
.A(n_450),
.Y(n_571)
);

CKINVDCx5p33_ASAP7_75t_R g572 ( 
.A(n_386),
.Y(n_572)
);

INVx1_ASAP7_75t_L g573 ( 
.A(n_266),
.Y(n_573)
);

INVx1_ASAP7_75t_L g574 ( 
.A(n_266),
.Y(n_574)
);

INVx1_ASAP7_75t_L g575 ( 
.A(n_266),
.Y(n_575)
);

CKINVDCx5p33_ASAP7_75t_R g576 ( 
.A(n_391),
.Y(n_576)
);

INVx1_ASAP7_75t_L g577 ( 
.A(n_293),
.Y(n_577)
);

INVx1_ASAP7_75t_L g578 ( 
.A(n_293),
.Y(n_578)
);

CKINVDCx5p33_ASAP7_75t_R g579 ( 
.A(n_392),
.Y(n_579)
);

CKINVDCx5p33_ASAP7_75t_R g580 ( 
.A(n_394),
.Y(n_580)
);

INVx1_ASAP7_75t_L g581 ( 
.A(n_293),
.Y(n_581)
);

INVxp67_ASAP7_75t_SL g582 ( 
.A(n_265),
.Y(n_582)
);

INVx1_ASAP7_75t_L g583 ( 
.A(n_252),
.Y(n_583)
);

INVx1_ASAP7_75t_L g584 ( 
.A(n_308),
.Y(n_584)
);

CKINVDCx20_ASAP7_75t_R g585 ( 
.A(n_397),
.Y(n_585)
);

INVxp33_ASAP7_75t_SL g586 ( 
.A(n_375),
.Y(n_586)
);

CKINVDCx20_ASAP7_75t_R g587 ( 
.A(n_410),
.Y(n_587)
);

NAND2xp5_ASAP7_75t_L g588 ( 
.A(n_269),
.B(n_406),
.Y(n_588)
);

NOR2xp67_ASAP7_75t_L g589 ( 
.A(n_437),
.B(n_12),
.Y(n_589)
);

AND2x2_ASAP7_75t_L g590 ( 
.A(n_437),
.B(n_12),
.Y(n_590)
);

INVx2_ASAP7_75t_L g591 ( 
.A(n_240),
.Y(n_591)
);

INVx1_ASAP7_75t_L g592 ( 
.A(n_308),
.Y(n_592)
);

CKINVDCx5p33_ASAP7_75t_R g593 ( 
.A(n_411),
.Y(n_593)
);

CKINVDCx5p33_ASAP7_75t_R g594 ( 
.A(n_417),
.Y(n_594)
);

CKINVDCx16_ASAP7_75t_R g595 ( 
.A(n_342),
.Y(n_595)
);

CKINVDCx5p33_ASAP7_75t_R g596 ( 
.A(n_421),
.Y(n_596)
);

INVxp67_ASAP7_75t_L g597 ( 
.A(n_444),
.Y(n_597)
);

INVx1_ASAP7_75t_L g598 ( 
.A(n_308),
.Y(n_598)
);

CKINVDCx20_ASAP7_75t_R g599 ( 
.A(n_422),
.Y(n_599)
);

INVxp33_ASAP7_75t_L g600 ( 
.A(n_253),
.Y(n_600)
);

INVx1_ASAP7_75t_L g601 ( 
.A(n_407),
.Y(n_601)
);

CKINVDCx5p33_ASAP7_75t_R g602 ( 
.A(n_476),
.Y(n_602)
);

INVx3_ASAP7_75t_L g603 ( 
.A(n_471),
.Y(n_603)
);

INVx1_ASAP7_75t_L g604 ( 
.A(n_497),
.Y(n_604)
);

CKINVDCx5p33_ASAP7_75t_R g605 ( 
.A(n_480),
.Y(n_605)
);

BUFx6f_ASAP7_75t_L g606 ( 
.A(n_591),
.Y(n_606)
);

CKINVDCx5p33_ASAP7_75t_R g607 ( 
.A(n_483),
.Y(n_607)
);

CKINVDCx5p33_ASAP7_75t_R g608 ( 
.A(n_487),
.Y(n_608)
);

INVx2_ASAP7_75t_L g609 ( 
.A(n_497),
.Y(n_609)
);

NAND2xp5_ASAP7_75t_L g610 ( 
.A(n_485),
.B(n_406),
.Y(n_610)
);

INVx1_ASAP7_75t_L g611 ( 
.A(n_498),
.Y(n_611)
);

INVx1_ASAP7_75t_L g612 ( 
.A(n_498),
.Y(n_612)
);

CKINVDCx20_ASAP7_75t_R g613 ( 
.A(n_472),
.Y(n_613)
);

AND2x4_ASAP7_75t_L g614 ( 
.A(n_486),
.B(n_406),
.Y(n_614)
);

CKINVDCx5p33_ASAP7_75t_R g615 ( 
.A(n_508),
.Y(n_615)
);

CKINVDCx5p33_ASAP7_75t_R g616 ( 
.A(n_510),
.Y(n_616)
);

BUFx6f_ASAP7_75t_L g617 ( 
.A(n_591),
.Y(n_617)
);

INVx2_ASAP7_75t_L g618 ( 
.A(n_499),
.Y(n_618)
);

INVx1_ASAP7_75t_L g619 ( 
.A(n_499),
.Y(n_619)
);

CKINVDCx16_ASAP7_75t_R g620 ( 
.A(n_475),
.Y(n_620)
);

INVx1_ASAP7_75t_L g621 ( 
.A(n_500),
.Y(n_621)
);

CKINVDCx5p33_ASAP7_75t_R g622 ( 
.A(n_511),
.Y(n_622)
);

INVx1_ASAP7_75t_L g623 ( 
.A(n_500),
.Y(n_623)
);

AND2x4_ASAP7_75t_L g624 ( 
.A(n_493),
.B(n_240),
.Y(n_624)
);

INVx1_ASAP7_75t_L g625 ( 
.A(n_501),
.Y(n_625)
);

BUFx2_ASAP7_75t_L g626 ( 
.A(n_514),
.Y(n_626)
);

INVx1_ASAP7_75t_L g627 ( 
.A(n_501),
.Y(n_627)
);

NOR2xp33_ASAP7_75t_R g628 ( 
.A(n_534),
.B(n_438),
.Y(n_628)
);

INVx1_ASAP7_75t_L g629 ( 
.A(n_502),
.Y(n_629)
);

BUFx6f_ASAP7_75t_L g630 ( 
.A(n_502),
.Y(n_630)
);

CKINVDCx5p33_ASAP7_75t_R g631 ( 
.A(n_513),
.Y(n_631)
);

INVx1_ASAP7_75t_L g632 ( 
.A(n_503),
.Y(n_632)
);

AND2x2_ASAP7_75t_L g633 ( 
.A(n_549),
.B(n_407),
.Y(n_633)
);

CKINVDCx5p33_ASAP7_75t_R g634 ( 
.A(n_520),
.Y(n_634)
);

CKINVDCx20_ASAP7_75t_R g635 ( 
.A(n_481),
.Y(n_635)
);

AND2x2_ASAP7_75t_L g636 ( 
.A(n_582),
.B(n_407),
.Y(n_636)
);

BUFx6f_ASAP7_75t_L g637 ( 
.A(n_503),
.Y(n_637)
);

CKINVDCx5p33_ASAP7_75t_R g638 ( 
.A(n_521),
.Y(n_638)
);

INVxp67_ASAP7_75t_L g639 ( 
.A(n_479),
.Y(n_639)
);

INVx1_ASAP7_75t_L g640 ( 
.A(n_505),
.Y(n_640)
);

AND2x2_ASAP7_75t_L g641 ( 
.A(n_573),
.B(n_574),
.Y(n_641)
);

NOR2xp67_ASAP7_75t_L g642 ( 
.A(n_471),
.B(n_240),
.Y(n_642)
);

INVx1_ASAP7_75t_L g643 ( 
.A(n_505),
.Y(n_643)
);

INVx2_ASAP7_75t_L g644 ( 
.A(n_506),
.Y(n_644)
);

CKINVDCx5p33_ASAP7_75t_R g645 ( 
.A(n_522),
.Y(n_645)
);

BUFx6f_ASAP7_75t_L g646 ( 
.A(n_506),
.Y(n_646)
);

CKINVDCx5p33_ASAP7_75t_R g647 ( 
.A(n_526),
.Y(n_647)
);

INVx1_ASAP7_75t_L g648 ( 
.A(n_507),
.Y(n_648)
);

CKINVDCx5p33_ASAP7_75t_R g649 ( 
.A(n_532),
.Y(n_649)
);

INVx1_ASAP7_75t_L g650 ( 
.A(n_507),
.Y(n_650)
);

CKINVDCx5p33_ASAP7_75t_R g651 ( 
.A(n_536),
.Y(n_651)
);

INVx2_ASAP7_75t_SL g652 ( 
.A(n_569),
.Y(n_652)
);

INVx1_ASAP7_75t_L g653 ( 
.A(n_509),
.Y(n_653)
);

INVx1_ASAP7_75t_L g654 ( 
.A(n_509),
.Y(n_654)
);

CKINVDCx5p33_ASAP7_75t_R g655 ( 
.A(n_538),
.Y(n_655)
);

INVx1_ASAP7_75t_L g656 ( 
.A(n_518),
.Y(n_656)
);

AND2x2_ASAP7_75t_L g657 ( 
.A(n_573),
.B(n_415),
.Y(n_657)
);

CKINVDCx5p33_ASAP7_75t_R g658 ( 
.A(n_540),
.Y(n_658)
);

INVxp67_ASAP7_75t_L g659 ( 
.A(n_479),
.Y(n_659)
);

INVx1_ASAP7_75t_L g660 ( 
.A(n_518),
.Y(n_660)
);

CKINVDCx5p33_ASAP7_75t_R g661 ( 
.A(n_545),
.Y(n_661)
);

CKINVDCx20_ASAP7_75t_R g662 ( 
.A(n_489),
.Y(n_662)
);

INVx1_ASAP7_75t_L g663 ( 
.A(n_523),
.Y(n_663)
);

INVx1_ASAP7_75t_L g664 ( 
.A(n_523),
.Y(n_664)
);

INVx1_ASAP7_75t_L g665 ( 
.A(n_527),
.Y(n_665)
);

INVx2_ASAP7_75t_L g666 ( 
.A(n_473),
.Y(n_666)
);

CKINVDCx20_ASAP7_75t_R g667 ( 
.A(n_494),
.Y(n_667)
);

CKINVDCx5p33_ASAP7_75t_R g668 ( 
.A(n_547),
.Y(n_668)
);

CKINVDCx5p33_ASAP7_75t_R g669 ( 
.A(n_551),
.Y(n_669)
);

INVx2_ASAP7_75t_L g670 ( 
.A(n_473),
.Y(n_670)
);

INVx3_ASAP7_75t_L g671 ( 
.A(n_474),
.Y(n_671)
);

INVx1_ASAP7_75t_L g672 ( 
.A(n_527),
.Y(n_672)
);

INVx2_ASAP7_75t_L g673 ( 
.A(n_474),
.Y(n_673)
);

CKINVDCx20_ASAP7_75t_R g674 ( 
.A(n_496),
.Y(n_674)
);

CKINVDCx5p33_ASAP7_75t_R g675 ( 
.A(n_552),
.Y(n_675)
);

INVxp67_ASAP7_75t_SL g676 ( 
.A(n_588),
.Y(n_676)
);

INVx1_ASAP7_75t_L g677 ( 
.A(n_528),
.Y(n_677)
);

CKINVDCx5p33_ASAP7_75t_R g678 ( 
.A(n_554),
.Y(n_678)
);

INVx2_ASAP7_75t_L g679 ( 
.A(n_477),
.Y(n_679)
);

INVx2_ASAP7_75t_L g680 ( 
.A(n_477),
.Y(n_680)
);

AOI22xp5_ASAP7_75t_L g681 ( 
.A1(n_517),
.A2(n_372),
.B1(n_261),
.B2(n_363),
.Y(n_681)
);

INVxp67_ASAP7_75t_L g682 ( 
.A(n_529),
.Y(n_682)
);

AND2x6_ASAP7_75t_L g683 ( 
.A(n_590),
.B(n_277),
.Y(n_683)
);

HB1xp67_ASAP7_75t_L g684 ( 
.A(n_569),
.Y(n_684)
);

INVx2_ASAP7_75t_L g685 ( 
.A(n_478),
.Y(n_685)
);

AND2x2_ASAP7_75t_L g686 ( 
.A(n_574),
.B(n_415),
.Y(n_686)
);

INVx1_ASAP7_75t_L g687 ( 
.A(n_528),
.Y(n_687)
);

INVx1_ASAP7_75t_L g688 ( 
.A(n_530),
.Y(n_688)
);

CKINVDCx5p33_ASAP7_75t_R g689 ( 
.A(n_555),
.Y(n_689)
);

CKINVDCx20_ASAP7_75t_R g690 ( 
.A(n_504),
.Y(n_690)
);

NOR2xp33_ASAP7_75t_R g691 ( 
.A(n_535),
.B(n_537),
.Y(n_691)
);

INVx1_ASAP7_75t_L g692 ( 
.A(n_530),
.Y(n_692)
);

HB1xp67_ASAP7_75t_L g693 ( 
.A(n_529),
.Y(n_693)
);

INVx2_ASAP7_75t_L g694 ( 
.A(n_478),
.Y(n_694)
);

CKINVDCx5p33_ASAP7_75t_R g695 ( 
.A(n_559),
.Y(n_695)
);

AND2x2_ASAP7_75t_L g696 ( 
.A(n_575),
.B(n_415),
.Y(n_696)
);

INVx1_ASAP7_75t_L g697 ( 
.A(n_488),
.Y(n_697)
);

CKINVDCx5p33_ASAP7_75t_R g698 ( 
.A(n_565),
.Y(n_698)
);

INVx2_ASAP7_75t_L g699 ( 
.A(n_488),
.Y(n_699)
);

INVx1_ASAP7_75t_L g700 ( 
.A(n_490),
.Y(n_700)
);

NAND2xp5_ASAP7_75t_L g701 ( 
.A(n_676),
.B(n_567),
.Y(n_701)
);

INVx1_ASAP7_75t_SL g702 ( 
.A(n_691),
.Y(n_702)
);

INVx2_ASAP7_75t_L g703 ( 
.A(n_606),
.Y(n_703)
);

NAND2xp5_ASAP7_75t_L g704 ( 
.A(n_676),
.B(n_572),
.Y(n_704)
);

INVx3_ASAP7_75t_L g705 ( 
.A(n_606),
.Y(n_705)
);

AOI22xp33_ASAP7_75t_L g706 ( 
.A1(n_683),
.A2(n_590),
.B1(n_586),
.B2(n_482),
.Y(n_706)
);

BUFx3_ASAP7_75t_L g707 ( 
.A(n_652),
.Y(n_707)
);

INVx4_ASAP7_75t_L g708 ( 
.A(n_606),
.Y(n_708)
);

INVx1_ASAP7_75t_L g709 ( 
.A(n_697),
.Y(n_709)
);

INVx4_ASAP7_75t_L g710 ( 
.A(n_606),
.Y(n_710)
);

HB1xp67_ASAP7_75t_L g711 ( 
.A(n_684),
.Y(n_711)
);

INVx2_ASAP7_75t_L g712 ( 
.A(n_606),
.Y(n_712)
);

INVx1_ASAP7_75t_L g713 ( 
.A(n_697),
.Y(n_713)
);

INVx4_ASAP7_75t_L g714 ( 
.A(n_606),
.Y(n_714)
);

AND2x2_ASAP7_75t_L g715 ( 
.A(n_641),
.B(n_575),
.Y(n_715)
);

INVx2_ASAP7_75t_L g716 ( 
.A(n_617),
.Y(n_716)
);

INVx1_ASAP7_75t_L g717 ( 
.A(n_700),
.Y(n_717)
);

AOI22xp5_ASAP7_75t_L g718 ( 
.A1(n_639),
.A2(n_484),
.B1(n_589),
.B2(n_372),
.Y(n_718)
);

AO21x2_ASAP7_75t_L g719 ( 
.A1(n_642),
.A2(n_283),
.B(n_282),
.Y(n_719)
);

AND2x4_ASAP7_75t_L g720 ( 
.A(n_652),
.B(n_512),
.Y(n_720)
);

AND2x4_ASAP7_75t_L g721 ( 
.A(n_652),
.B(n_282),
.Y(n_721)
);

INVx2_ASAP7_75t_L g722 ( 
.A(n_617),
.Y(n_722)
);

NAND2x1p5_ASAP7_75t_L g723 ( 
.A(n_624),
.B(n_259),
.Y(n_723)
);

NAND2xp5_ASAP7_75t_SL g724 ( 
.A(n_602),
.B(n_576),
.Y(n_724)
);

INVx1_ASAP7_75t_L g725 ( 
.A(n_700),
.Y(n_725)
);

INVx3_ASAP7_75t_L g726 ( 
.A(n_617),
.Y(n_726)
);

AND2x4_ASAP7_75t_L g727 ( 
.A(n_624),
.B(n_283),
.Y(n_727)
);

BUFx6f_ASAP7_75t_L g728 ( 
.A(n_617),
.Y(n_728)
);

INVx2_ASAP7_75t_L g729 ( 
.A(n_617),
.Y(n_729)
);

INVx1_ASAP7_75t_L g730 ( 
.A(n_666),
.Y(n_730)
);

INVx1_ASAP7_75t_L g731 ( 
.A(n_666),
.Y(n_731)
);

BUFx6f_ASAP7_75t_L g732 ( 
.A(n_617),
.Y(n_732)
);

NAND2x1p5_ASAP7_75t_L g733 ( 
.A(n_624),
.B(n_259),
.Y(n_733)
);

NAND2xp5_ASAP7_75t_SL g734 ( 
.A(n_605),
.B(n_579),
.Y(n_734)
);

NAND2xp5_ASAP7_75t_L g735 ( 
.A(n_614),
.B(n_580),
.Y(n_735)
);

CKINVDCx5p33_ASAP7_75t_R g736 ( 
.A(n_607),
.Y(n_736)
);

NOR2xp33_ASAP7_75t_L g737 ( 
.A(n_684),
.B(n_593),
.Y(n_737)
);

INVx4_ASAP7_75t_L g738 ( 
.A(n_630),
.Y(n_738)
);

NAND2xp5_ASAP7_75t_L g739 ( 
.A(n_614),
.B(n_594),
.Y(n_739)
);

OR2x2_ASAP7_75t_L g740 ( 
.A(n_693),
.B(n_558),
.Y(n_740)
);

BUFx3_ASAP7_75t_L g741 ( 
.A(n_683),
.Y(n_741)
);

INVx1_ASAP7_75t_L g742 ( 
.A(n_666),
.Y(n_742)
);

NAND2xp5_ASAP7_75t_L g743 ( 
.A(n_614),
.B(n_683),
.Y(n_743)
);

BUFx6f_ASAP7_75t_L g744 ( 
.A(n_630),
.Y(n_744)
);

NAND2xp5_ASAP7_75t_L g745 ( 
.A(n_614),
.B(n_596),
.Y(n_745)
);

INVx2_ASAP7_75t_L g746 ( 
.A(n_609),
.Y(n_746)
);

NAND2xp5_ASAP7_75t_L g747 ( 
.A(n_683),
.B(n_546),
.Y(n_747)
);

INVx1_ASAP7_75t_L g748 ( 
.A(n_670),
.Y(n_748)
);

AOI22xp5_ASAP7_75t_L g749 ( 
.A1(n_639),
.A2(n_261),
.B1(n_544),
.B2(n_531),
.Y(n_749)
);

CKINVDCx16_ASAP7_75t_R g750 ( 
.A(n_620),
.Y(n_750)
);

INVx1_ASAP7_75t_L g751 ( 
.A(n_670),
.Y(n_751)
);

BUFx6f_ASAP7_75t_L g752 ( 
.A(n_630),
.Y(n_752)
);

NAND2xp5_ASAP7_75t_SL g753 ( 
.A(n_608),
.B(n_595),
.Y(n_753)
);

INVx4_ASAP7_75t_L g754 ( 
.A(n_630),
.Y(n_754)
);

INVx2_ASAP7_75t_L g755 ( 
.A(n_609),
.Y(n_755)
);

NOR2xp33_ASAP7_75t_L g756 ( 
.A(n_615),
.B(n_560),
.Y(n_756)
);

INVx2_ASAP7_75t_L g757 ( 
.A(n_609),
.Y(n_757)
);

INVx2_ASAP7_75t_L g758 ( 
.A(n_618),
.Y(n_758)
);

BUFx2_ASAP7_75t_L g759 ( 
.A(n_626),
.Y(n_759)
);

OR2x2_ASAP7_75t_L g760 ( 
.A(n_693),
.B(n_597),
.Y(n_760)
);

INVx8_ASAP7_75t_L g761 ( 
.A(n_683),
.Y(n_761)
);

AND2x4_ASAP7_75t_L g762 ( 
.A(n_624),
.B(n_284),
.Y(n_762)
);

INVx1_ASAP7_75t_L g763 ( 
.A(n_670),
.Y(n_763)
);

AND2x2_ASAP7_75t_L g764 ( 
.A(n_641),
.B(n_577),
.Y(n_764)
);

INVx1_ASAP7_75t_L g765 ( 
.A(n_673),
.Y(n_765)
);

INVx1_ASAP7_75t_L g766 ( 
.A(n_673),
.Y(n_766)
);

AND2x4_ASAP7_75t_L g767 ( 
.A(n_641),
.B(n_284),
.Y(n_767)
);

INVx1_ASAP7_75t_L g768 ( 
.A(n_673),
.Y(n_768)
);

INVx2_ASAP7_75t_L g769 ( 
.A(n_618),
.Y(n_769)
);

BUFx6f_ASAP7_75t_L g770 ( 
.A(n_630),
.Y(n_770)
);

INVx3_ASAP7_75t_L g771 ( 
.A(n_630),
.Y(n_771)
);

NAND2xp5_ASAP7_75t_L g772 ( 
.A(n_683),
.B(n_633),
.Y(n_772)
);

INVxp67_ASAP7_75t_SL g773 ( 
.A(n_603),
.Y(n_773)
);

INVx1_ASAP7_75t_L g774 ( 
.A(n_679),
.Y(n_774)
);

INVx1_ASAP7_75t_L g775 ( 
.A(n_679),
.Y(n_775)
);

OR2x6_ASAP7_75t_L g776 ( 
.A(n_633),
.B(n_324),
.Y(n_776)
);

INVx2_ASAP7_75t_L g777 ( 
.A(n_618),
.Y(n_777)
);

NAND2xp5_ASAP7_75t_L g778 ( 
.A(n_683),
.B(n_548),
.Y(n_778)
);

BUFx2_ASAP7_75t_L g779 ( 
.A(n_626),
.Y(n_779)
);

INVx2_ASAP7_75t_L g780 ( 
.A(n_644),
.Y(n_780)
);

INVx1_ASAP7_75t_L g781 ( 
.A(n_679),
.Y(n_781)
);

AOI22xp33_ASAP7_75t_L g782 ( 
.A1(n_683),
.A2(n_633),
.B1(n_636),
.B2(n_610),
.Y(n_782)
);

INVx4_ASAP7_75t_L g783 ( 
.A(n_637),
.Y(n_783)
);

NAND2xp5_ASAP7_75t_L g784 ( 
.A(n_636),
.B(n_524),
.Y(n_784)
);

NAND2xp5_ASAP7_75t_L g785 ( 
.A(n_636),
.B(n_610),
.Y(n_785)
);

NAND2xp5_ASAP7_75t_SL g786 ( 
.A(n_616),
.B(n_564),
.Y(n_786)
);

BUFx6f_ASAP7_75t_L g787 ( 
.A(n_637),
.Y(n_787)
);

BUFx3_ASAP7_75t_L g788 ( 
.A(n_603),
.Y(n_788)
);

INVx3_ASAP7_75t_L g789 ( 
.A(n_637),
.Y(n_789)
);

INVx3_ASAP7_75t_L g790 ( 
.A(n_637),
.Y(n_790)
);

NAND2xp5_ASAP7_75t_L g791 ( 
.A(n_603),
.B(n_583),
.Y(n_791)
);

AOI22xp33_ASAP7_75t_L g792 ( 
.A1(n_657),
.A2(n_556),
.B1(n_519),
.B2(n_516),
.Y(n_792)
);

BUFx3_ASAP7_75t_L g793 ( 
.A(n_603),
.Y(n_793)
);

INVx3_ASAP7_75t_L g794 ( 
.A(n_637),
.Y(n_794)
);

NOR2xp33_ASAP7_75t_L g795 ( 
.A(n_622),
.B(n_585),
.Y(n_795)
);

NOR2xp33_ASAP7_75t_L g796 ( 
.A(n_631),
.B(n_587),
.Y(n_796)
);

BUFx6f_ASAP7_75t_L g797 ( 
.A(n_637),
.Y(n_797)
);

AND2x2_ASAP7_75t_L g798 ( 
.A(n_657),
.B(n_601),
.Y(n_798)
);

INVx3_ASAP7_75t_L g799 ( 
.A(n_646),
.Y(n_799)
);

AND2x2_ASAP7_75t_L g800 ( 
.A(n_657),
.B(n_601),
.Y(n_800)
);

BUFx4f_ASAP7_75t_L g801 ( 
.A(n_646),
.Y(n_801)
);

CKINVDCx5p33_ASAP7_75t_R g802 ( 
.A(n_634),
.Y(n_802)
);

INVx3_ASAP7_75t_L g803 ( 
.A(n_646),
.Y(n_803)
);

NAND2xp5_ASAP7_75t_SL g804 ( 
.A(n_638),
.B(n_599),
.Y(n_804)
);

INVx3_ASAP7_75t_L g805 ( 
.A(n_646),
.Y(n_805)
);

NOR2xp33_ASAP7_75t_L g806 ( 
.A(n_645),
.B(n_600),
.Y(n_806)
);

NAND2xp5_ASAP7_75t_L g807 ( 
.A(n_671),
.B(n_490),
.Y(n_807)
);

BUFx10_ASAP7_75t_L g808 ( 
.A(n_647),
.Y(n_808)
);

NAND2xp5_ASAP7_75t_L g809 ( 
.A(n_671),
.B(n_491),
.Y(n_809)
);

AND2x2_ASAP7_75t_L g810 ( 
.A(n_686),
.B(n_598),
.Y(n_810)
);

INVx1_ASAP7_75t_L g811 ( 
.A(n_680),
.Y(n_811)
);

AND2x2_ASAP7_75t_L g812 ( 
.A(n_686),
.B(n_598),
.Y(n_812)
);

AOI22xp33_ASAP7_75t_L g813 ( 
.A1(n_686),
.A2(n_516),
.B1(n_455),
.B2(n_264),
.Y(n_813)
);

AND2x4_ASAP7_75t_L g814 ( 
.A(n_696),
.B(n_298),
.Y(n_814)
);

BUFx3_ASAP7_75t_L g815 ( 
.A(n_671),
.Y(n_815)
);

INVx1_ASAP7_75t_L g816 ( 
.A(n_680),
.Y(n_816)
);

INVx2_ASAP7_75t_L g817 ( 
.A(n_644),
.Y(n_817)
);

INVx2_ASAP7_75t_L g818 ( 
.A(n_644),
.Y(n_818)
);

BUFx6f_ASAP7_75t_L g819 ( 
.A(n_646),
.Y(n_819)
);

INVx1_ASAP7_75t_L g820 ( 
.A(n_680),
.Y(n_820)
);

NAND2xp33_ASAP7_75t_L g821 ( 
.A(n_649),
.B(n_440),
.Y(n_821)
);

OR2x2_ASAP7_75t_L g822 ( 
.A(n_659),
.B(n_577),
.Y(n_822)
);

INVx1_ASAP7_75t_L g823 ( 
.A(n_685),
.Y(n_823)
);

BUFx6f_ASAP7_75t_L g824 ( 
.A(n_646),
.Y(n_824)
);

INVx1_ASAP7_75t_L g825 ( 
.A(n_685),
.Y(n_825)
);

AND2x4_ASAP7_75t_L g826 ( 
.A(n_696),
.B(n_298),
.Y(n_826)
);

CKINVDCx5p33_ASAP7_75t_R g827 ( 
.A(n_651),
.Y(n_827)
);

BUFx3_ASAP7_75t_L g828 ( 
.A(n_671),
.Y(n_828)
);

INVx2_ASAP7_75t_L g829 ( 
.A(n_685),
.Y(n_829)
);

BUFx6f_ASAP7_75t_L g830 ( 
.A(n_694),
.Y(n_830)
);

INVxp67_ASAP7_75t_L g831 ( 
.A(n_696),
.Y(n_831)
);

AND2x6_ASAP7_75t_L g832 ( 
.A(n_694),
.B(n_277),
.Y(n_832)
);

NOR3xp33_ASAP7_75t_L g833 ( 
.A(n_659),
.B(n_412),
.C(n_401),
.Y(n_833)
);

AND2x4_ASAP7_75t_L g834 ( 
.A(n_663),
.B(n_303),
.Y(n_834)
);

INVx2_ASAP7_75t_L g835 ( 
.A(n_694),
.Y(n_835)
);

NAND2xp5_ASAP7_75t_L g836 ( 
.A(n_699),
.B(n_491),
.Y(n_836)
);

INVx1_ASAP7_75t_L g837 ( 
.A(n_699),
.Y(n_837)
);

INVx2_ASAP7_75t_L g838 ( 
.A(n_699),
.Y(n_838)
);

INVx1_ASAP7_75t_SL g839 ( 
.A(n_674),
.Y(n_839)
);

AOI22xp33_ASAP7_75t_L g840 ( 
.A1(n_663),
.A2(n_455),
.B1(n_264),
.B2(n_268),
.Y(n_840)
);

INVxp67_ASAP7_75t_L g841 ( 
.A(n_682),
.Y(n_841)
);

INVx1_ASAP7_75t_L g842 ( 
.A(n_604),
.Y(n_842)
);

NOR2xp33_ASAP7_75t_L g843 ( 
.A(n_655),
.B(n_578),
.Y(n_843)
);

INVx4_ASAP7_75t_L g844 ( 
.A(n_604),
.Y(n_844)
);

AND2x2_ASAP7_75t_L g845 ( 
.A(n_664),
.B(n_578),
.Y(n_845)
);

AND2x2_ASAP7_75t_SL g846 ( 
.A(n_620),
.B(n_277),
.Y(n_846)
);

NAND2xp5_ASAP7_75t_L g847 ( 
.A(n_611),
.B(n_492),
.Y(n_847)
);

INVx3_ASAP7_75t_L g848 ( 
.A(n_611),
.Y(n_848)
);

BUFx2_ASAP7_75t_L g849 ( 
.A(n_682),
.Y(n_849)
);

CKINVDCx5p33_ASAP7_75t_R g850 ( 
.A(n_658),
.Y(n_850)
);

AND2x6_ASAP7_75t_L g851 ( 
.A(n_664),
.B(n_280),
.Y(n_851)
);

AND2x4_ASAP7_75t_L g852 ( 
.A(n_665),
.B(n_672),
.Y(n_852)
);

INVx2_ASAP7_75t_L g853 ( 
.A(n_612),
.Y(n_853)
);

NAND2xp5_ASAP7_75t_SL g854 ( 
.A(n_661),
.B(n_358),
.Y(n_854)
);

OR2x2_ASAP7_75t_L g855 ( 
.A(n_681),
.B(n_581),
.Y(n_855)
);

NOR2xp33_ASAP7_75t_L g856 ( 
.A(n_668),
.B(n_581),
.Y(n_856)
);

AND2x4_ASAP7_75t_L g857 ( 
.A(n_665),
.B(n_303),
.Y(n_857)
);

INVx1_ASAP7_75t_L g858 ( 
.A(n_612),
.Y(n_858)
);

INVx1_ASAP7_75t_L g859 ( 
.A(n_619),
.Y(n_859)
);

INVx4_ASAP7_75t_L g860 ( 
.A(n_619),
.Y(n_860)
);

NAND2xp5_ASAP7_75t_SL g861 ( 
.A(n_698),
.B(n_358),
.Y(n_861)
);

CKINVDCx5p33_ASAP7_75t_R g862 ( 
.A(n_669),
.Y(n_862)
);

NAND2xp5_ASAP7_75t_L g863 ( 
.A(n_621),
.B(n_492),
.Y(n_863)
);

INVx1_ASAP7_75t_L g864 ( 
.A(n_621),
.Y(n_864)
);

AOI22xp5_ASAP7_75t_L g865 ( 
.A1(n_782),
.A2(n_681),
.B1(n_385),
.B2(n_418),
.Y(n_865)
);

OAI221xp5_ASAP7_75t_L g866 ( 
.A1(n_706),
.A2(n_285),
.B1(n_289),
.B2(n_268),
.C(n_254),
.Y(n_866)
);

OR2x6_ASAP7_75t_L g867 ( 
.A(n_776),
.B(n_324),
.Y(n_867)
);

INVx5_ASAP7_75t_L g868 ( 
.A(n_761),
.Y(n_868)
);

AND2x2_ASAP7_75t_L g869 ( 
.A(n_798),
.B(n_672),
.Y(n_869)
);

AOI22xp5_ASAP7_75t_L g870 ( 
.A1(n_846),
.A2(n_678),
.B1(n_689),
.B2(n_675),
.Y(n_870)
);

NOR2xp33_ASAP7_75t_L g871 ( 
.A(n_806),
.B(n_695),
.Y(n_871)
);

NAND2xp5_ASAP7_75t_L g872 ( 
.A(n_785),
.B(n_677),
.Y(n_872)
);

BUFx6f_ASAP7_75t_L g873 ( 
.A(n_741),
.Y(n_873)
);

INVx2_ASAP7_75t_L g874 ( 
.A(n_853),
.Y(n_874)
);

BUFx6f_ASAP7_75t_L g875 ( 
.A(n_741),
.Y(n_875)
);

NOR2xp33_ASAP7_75t_SL g876 ( 
.A(n_702),
.B(n_613),
.Y(n_876)
);

OAI22xp5_ASAP7_75t_L g877 ( 
.A1(n_723),
.A2(n_379),
.B1(n_360),
.B2(n_290),
.Y(n_877)
);

AND2x2_ASAP7_75t_L g878 ( 
.A(n_798),
.B(n_677),
.Y(n_878)
);

INVx2_ASAP7_75t_L g879 ( 
.A(n_853),
.Y(n_879)
);

NAND2x1p5_ASAP7_75t_L g880 ( 
.A(n_741),
.B(n_305),
.Y(n_880)
);

AO221x1_ASAP7_75t_L g881 ( 
.A1(n_831),
.A2(n_321),
.B1(n_329),
.B2(n_316),
.C(n_305),
.Y(n_881)
);

OAI21xp5_ASAP7_75t_L g882 ( 
.A1(n_772),
.A2(n_642),
.B(n_495),
.Y(n_882)
);

NAND2xp5_ASAP7_75t_L g883 ( 
.A(n_707),
.B(n_687),
.Y(n_883)
);

AOI21xp5_ASAP7_75t_L g884 ( 
.A1(n_743),
.A2(n_773),
.B(n_784),
.Y(n_884)
);

INVx2_ASAP7_75t_L g885 ( 
.A(n_709),
.Y(n_885)
);

NAND2xp5_ASAP7_75t_L g886 ( 
.A(n_707),
.B(n_687),
.Y(n_886)
);

NAND2xp5_ASAP7_75t_L g887 ( 
.A(n_707),
.B(n_688),
.Y(n_887)
);

INVx3_ASAP7_75t_L g888 ( 
.A(n_788),
.Y(n_888)
);

NAND2xp5_ASAP7_75t_SL g889 ( 
.A(n_701),
.B(n_628),
.Y(n_889)
);

INVx2_ASAP7_75t_L g890 ( 
.A(n_709),
.Y(n_890)
);

NAND2xp5_ASAP7_75t_L g891 ( 
.A(n_720),
.B(n_688),
.Y(n_891)
);

INVx1_ASAP7_75t_L g892 ( 
.A(n_713),
.Y(n_892)
);

NAND2xp5_ASAP7_75t_L g893 ( 
.A(n_720),
.B(n_692),
.Y(n_893)
);

AND2x2_ASAP7_75t_L g894 ( 
.A(n_800),
.B(n_692),
.Y(n_894)
);

NAND2xp5_ASAP7_75t_SL g895 ( 
.A(n_704),
.B(n_360),
.Y(n_895)
);

NAND2xp5_ASAP7_75t_L g896 ( 
.A(n_720),
.B(n_623),
.Y(n_896)
);

INVx2_ASAP7_75t_L g897 ( 
.A(n_713),
.Y(n_897)
);

INVx2_ASAP7_75t_L g898 ( 
.A(n_717),
.Y(n_898)
);

NAND2xp5_ASAP7_75t_L g899 ( 
.A(n_720),
.B(n_623),
.Y(n_899)
);

OAI22xp5_ASAP7_75t_L g900 ( 
.A1(n_723),
.A2(n_733),
.B1(n_776),
.B2(n_747),
.Y(n_900)
);

INVx1_ASAP7_75t_L g901 ( 
.A(n_717),
.Y(n_901)
);

NAND2xp5_ASAP7_75t_L g902 ( 
.A(n_725),
.B(n_625),
.Y(n_902)
);

AND2x4_ASAP7_75t_L g903 ( 
.A(n_800),
.B(n_316),
.Y(n_903)
);

NAND2xp5_ASAP7_75t_L g904 ( 
.A(n_725),
.B(n_625),
.Y(n_904)
);

BUFx8_ASAP7_75t_L g905 ( 
.A(n_759),
.Y(n_905)
);

NAND2xp5_ASAP7_75t_L g906 ( 
.A(n_852),
.B(n_627),
.Y(n_906)
);

INVx2_ASAP7_75t_SL g907 ( 
.A(n_810),
.Y(n_907)
);

NAND2xp5_ASAP7_75t_L g908 ( 
.A(n_852),
.B(n_627),
.Y(n_908)
);

A2O1A1Ixp33_ASAP7_75t_L g909 ( 
.A1(n_778),
.A2(n_280),
.B(n_313),
.C(n_290),
.Y(n_909)
);

NAND2xp5_ASAP7_75t_SL g910 ( 
.A(n_846),
.B(n_379),
.Y(n_910)
);

OAI22xp33_ASAP7_75t_L g911 ( 
.A1(n_749),
.A2(n_329),
.B1(n_330),
.B2(n_321),
.Y(n_911)
);

INVx1_ASAP7_75t_L g912 ( 
.A(n_852),
.Y(n_912)
);

NAND2xp5_ASAP7_75t_L g913 ( 
.A(n_852),
.B(n_629),
.Y(n_913)
);

NAND2xp5_ASAP7_75t_L g914 ( 
.A(n_723),
.B(n_629),
.Y(n_914)
);

AOI22xp5_ASAP7_75t_L g915 ( 
.A1(n_846),
.A2(n_525),
.B1(n_515),
.B2(n_443),
.Y(n_915)
);

NOR2xp33_ASAP7_75t_SL g916 ( 
.A(n_736),
.B(n_635),
.Y(n_916)
);

NAND2xp5_ASAP7_75t_L g917 ( 
.A(n_733),
.B(n_632),
.Y(n_917)
);

AND2x2_ASAP7_75t_L g918 ( 
.A(n_810),
.B(n_584),
.Y(n_918)
);

OR2x6_ASAP7_75t_L g919 ( 
.A(n_776),
.B(n_444),
.Y(n_919)
);

OR2x2_ASAP7_75t_L g920 ( 
.A(n_760),
.B(n_401),
.Y(n_920)
);

NOR2xp33_ASAP7_75t_L g921 ( 
.A(n_843),
.B(n_662),
.Y(n_921)
);

INVx2_ASAP7_75t_L g922 ( 
.A(n_842),
.Y(n_922)
);

AND2x2_ASAP7_75t_L g923 ( 
.A(n_812),
.B(n_584),
.Y(n_923)
);

INVx4_ASAP7_75t_L g924 ( 
.A(n_761),
.Y(n_924)
);

INVx3_ASAP7_75t_L g925 ( 
.A(n_788),
.Y(n_925)
);

NAND2xp5_ASAP7_75t_SL g926 ( 
.A(n_733),
.B(n_441),
.Y(n_926)
);

NOR2xp33_ASAP7_75t_L g927 ( 
.A(n_856),
.B(n_667),
.Y(n_927)
);

NAND2xp5_ASAP7_75t_SL g928 ( 
.A(n_735),
.B(n_446),
.Y(n_928)
);

NAND2xp5_ASAP7_75t_L g929 ( 
.A(n_715),
.B(n_632),
.Y(n_929)
);

NOR2xp33_ASAP7_75t_L g930 ( 
.A(n_841),
.B(n_690),
.Y(n_930)
);

NOR2xp33_ASAP7_75t_SL g931 ( 
.A(n_802),
.B(n_296),
.Y(n_931)
);

NAND2xp5_ASAP7_75t_L g932 ( 
.A(n_715),
.B(n_640),
.Y(n_932)
);

NOR2xp33_ASAP7_75t_L g933 ( 
.A(n_737),
.B(n_739),
.Y(n_933)
);

AOI22xp5_ASAP7_75t_L g934 ( 
.A1(n_776),
.A2(n_465),
.B1(n_331),
.B2(n_353),
.Y(n_934)
);

AOI22xp5_ASAP7_75t_L g935 ( 
.A1(n_776),
.A2(n_331),
.B1(n_353),
.B2(n_330),
.Y(n_935)
);

NOR2xp33_ASAP7_75t_L g936 ( 
.A(n_745),
.B(n_412),
.Y(n_936)
);

NAND2xp5_ASAP7_75t_L g937 ( 
.A(n_764),
.B(n_844),
.Y(n_937)
);

AND2x6_ASAP7_75t_SL g938 ( 
.A(n_756),
.B(n_254),
.Y(n_938)
);

AOI22xp33_ASAP7_75t_L g939 ( 
.A1(n_814),
.A2(n_826),
.B1(n_767),
.B2(n_727),
.Y(n_939)
);

NAND2xp5_ASAP7_75t_L g940 ( 
.A(n_764),
.B(n_640),
.Y(n_940)
);

HB1xp67_ASAP7_75t_L g941 ( 
.A(n_759),
.Y(n_941)
);

NOR2x1p5_ASAP7_75t_L g942 ( 
.A(n_740),
.B(n_455),
.Y(n_942)
);

NAND2xp5_ASAP7_75t_SL g943 ( 
.A(n_822),
.B(n_358),
.Y(n_943)
);

CKINVDCx5p33_ASAP7_75t_R g944 ( 
.A(n_827),
.Y(n_944)
);

NAND2xp5_ASAP7_75t_L g945 ( 
.A(n_844),
.B(n_643),
.Y(n_945)
);

NAND2xp33_ASAP7_75t_L g946 ( 
.A(n_761),
.B(n_311),
.Y(n_946)
);

INVx2_ASAP7_75t_L g947 ( 
.A(n_842),
.Y(n_947)
);

INVx2_ASAP7_75t_L g948 ( 
.A(n_858),
.Y(n_948)
);

AOI22xp33_ASAP7_75t_L g949 ( 
.A1(n_814),
.A2(n_290),
.B1(n_313),
.B2(n_280),
.Y(n_949)
);

INVx2_ASAP7_75t_L g950 ( 
.A(n_858),
.Y(n_950)
);

NAND2xp5_ASAP7_75t_SL g951 ( 
.A(n_822),
.B(n_358),
.Y(n_951)
);

INVx1_ASAP7_75t_L g952 ( 
.A(n_859),
.Y(n_952)
);

NAND2xp5_ASAP7_75t_L g953 ( 
.A(n_844),
.B(n_643),
.Y(n_953)
);

NAND2xp5_ASAP7_75t_L g954 ( 
.A(n_844),
.B(n_648),
.Y(n_954)
);

NAND2xp5_ASAP7_75t_SL g955 ( 
.A(n_760),
.B(n_356),
.Y(n_955)
);

INVx2_ASAP7_75t_SL g956 ( 
.A(n_812),
.Y(n_956)
);

BUFx8_ASAP7_75t_L g957 ( 
.A(n_779),
.Y(n_957)
);

AND2x4_ASAP7_75t_L g958 ( 
.A(n_814),
.B(n_356),
.Y(n_958)
);

INVxp67_ASAP7_75t_L g959 ( 
.A(n_849),
.Y(n_959)
);

INVxp67_ASAP7_75t_L g960 ( 
.A(n_849),
.Y(n_960)
);

INVx1_ASAP7_75t_L g961 ( 
.A(n_859),
.Y(n_961)
);

NAND2xp5_ASAP7_75t_L g962 ( 
.A(n_860),
.B(n_648),
.Y(n_962)
);

INVx2_ASAP7_75t_L g963 ( 
.A(n_864),
.Y(n_963)
);

NAND2xp5_ASAP7_75t_L g964 ( 
.A(n_860),
.B(n_650),
.Y(n_964)
);

NAND3xp33_ASAP7_75t_L g965 ( 
.A(n_749),
.B(n_241),
.C(n_239),
.Y(n_965)
);

INVx1_ASAP7_75t_L g966 ( 
.A(n_864),
.Y(n_966)
);

CKINVDCx5p33_ASAP7_75t_R g967 ( 
.A(n_850),
.Y(n_967)
);

INVx2_ASAP7_75t_L g968 ( 
.A(n_829),
.Y(n_968)
);

NAND2xp5_ASAP7_75t_L g969 ( 
.A(n_860),
.B(n_650),
.Y(n_969)
);

OAI22xp5_ASAP7_75t_L g970 ( 
.A1(n_718),
.A2(n_338),
.B1(n_393),
.B2(n_313),
.Y(n_970)
);

AOI22xp33_ASAP7_75t_L g971 ( 
.A1(n_814),
.A2(n_338),
.B1(n_458),
.B2(n_393),
.Y(n_971)
);

NAND2xp5_ASAP7_75t_L g972 ( 
.A(n_860),
.B(n_653),
.Y(n_972)
);

OR2x2_ASAP7_75t_L g973 ( 
.A(n_740),
.B(n_467),
.Y(n_973)
);

AOI22xp33_ASAP7_75t_L g974 ( 
.A1(n_826),
.A2(n_338),
.B1(n_458),
.B2(n_393),
.Y(n_974)
);

NAND2xp5_ASAP7_75t_L g975 ( 
.A(n_721),
.B(n_653),
.Y(n_975)
);

INVx1_ASAP7_75t_L g976 ( 
.A(n_848),
.Y(n_976)
);

A2O1A1Ixp33_ASAP7_75t_L g977 ( 
.A1(n_767),
.A2(n_458),
.B(n_495),
.C(n_364),
.Y(n_977)
);

NOR2xp33_ASAP7_75t_L g978 ( 
.A(n_711),
.B(n_467),
.Y(n_978)
);

INVxp67_ASAP7_75t_SL g979 ( 
.A(n_830),
.Y(n_979)
);

NAND2xp5_ASAP7_75t_L g980 ( 
.A(n_721),
.B(n_654),
.Y(n_980)
);

AOI22xp33_ASAP7_75t_L g981 ( 
.A1(n_826),
.A2(n_359),
.B1(n_365),
.B2(n_364),
.Y(n_981)
);

NOR2xp33_ASAP7_75t_L g982 ( 
.A(n_724),
.B(n_734),
.Y(n_982)
);

AOI22xp33_ASAP7_75t_L g983 ( 
.A1(n_826),
.A2(n_359),
.B1(n_367),
.B2(n_365),
.Y(n_983)
);

NAND2xp5_ASAP7_75t_SL g984 ( 
.A(n_718),
.B(n_367),
.Y(n_984)
);

A2O1A1Ixp33_ASAP7_75t_L g985 ( 
.A1(n_767),
.A2(n_402),
.B(n_403),
.C(n_381),
.Y(n_985)
);

AOI22xp33_ASAP7_75t_L g986 ( 
.A1(n_767),
.A2(n_762),
.B1(n_727),
.B2(n_834),
.Y(n_986)
);

NAND2xp5_ASAP7_75t_L g987 ( 
.A(n_721),
.B(n_654),
.Y(n_987)
);

NAND2xp5_ASAP7_75t_SL g988 ( 
.A(n_808),
.B(n_381),
.Y(n_988)
);

AND2x2_ASAP7_75t_L g989 ( 
.A(n_845),
.B(n_592),
.Y(n_989)
);

INVx1_ASAP7_75t_L g990 ( 
.A(n_848),
.Y(n_990)
);

NAND2xp5_ASAP7_75t_SL g991 ( 
.A(n_808),
.B(n_402),
.Y(n_991)
);

INVx1_ASAP7_75t_L g992 ( 
.A(n_848),
.Y(n_992)
);

NAND2xp5_ASAP7_75t_L g993 ( 
.A(n_721),
.B(n_656),
.Y(n_993)
);

OAI22xp5_ASAP7_75t_L g994 ( 
.A1(n_727),
.A2(n_425),
.B1(n_428),
.B2(n_403),
.Y(n_994)
);

NAND2xp5_ASAP7_75t_L g995 ( 
.A(n_727),
.B(n_656),
.Y(n_995)
);

NAND2xp5_ASAP7_75t_SL g996 ( 
.A(n_808),
.B(n_425),
.Y(n_996)
);

INVx2_ASAP7_75t_SL g997 ( 
.A(n_762),
.Y(n_997)
);

INVx2_ASAP7_75t_SL g998 ( 
.A(n_762),
.Y(n_998)
);

BUFx6f_ASAP7_75t_L g999 ( 
.A(n_788),
.Y(n_999)
);

AOI22xp33_ASAP7_75t_L g1000 ( 
.A1(n_762),
.A2(n_428),
.B1(n_460),
.B2(n_436),
.Y(n_1000)
);

NOR2xp67_ASAP7_75t_SL g1001 ( 
.A(n_793),
.B(n_436),
.Y(n_1001)
);

AOI22xp33_ASAP7_75t_L g1002 ( 
.A1(n_834),
.A2(n_460),
.B1(n_470),
.B2(n_468),
.Y(n_1002)
);

INVx1_ASAP7_75t_L g1003 ( 
.A(n_848),
.Y(n_1003)
);

NAND2xp5_ASAP7_75t_SL g1004 ( 
.A(n_808),
.B(n_792),
.Y(n_1004)
);

NAND2xp5_ASAP7_75t_SL g1005 ( 
.A(n_854),
.B(n_468),
.Y(n_1005)
);

INVx2_ASAP7_75t_L g1006 ( 
.A(n_829),
.Y(n_1006)
);

NAND2xp5_ASAP7_75t_L g1007 ( 
.A(n_793),
.B(n_660),
.Y(n_1007)
);

O2A1O1Ixp33_ASAP7_75t_L g1008 ( 
.A1(n_855),
.A2(n_592),
.B(n_289),
.C(n_292),
.Y(n_1008)
);

INVx1_ASAP7_75t_L g1009 ( 
.A(n_730),
.Y(n_1009)
);

NAND2xp5_ASAP7_75t_L g1010 ( 
.A(n_793),
.B(n_660),
.Y(n_1010)
);

INVx2_ASAP7_75t_L g1011 ( 
.A(n_835),
.Y(n_1011)
);

NAND2xp5_ASAP7_75t_SL g1012 ( 
.A(n_861),
.B(n_813),
.Y(n_1012)
);

INVx2_ASAP7_75t_L g1013 ( 
.A(n_835),
.Y(n_1013)
);

NAND2xp5_ASAP7_75t_L g1014 ( 
.A(n_815),
.B(n_470),
.Y(n_1014)
);

O2A1O1Ixp5_ASAP7_75t_L g1015 ( 
.A1(n_791),
.A2(n_539),
.B(n_541),
.C(n_533),
.Y(n_1015)
);

AOI22xp33_ASAP7_75t_L g1016 ( 
.A1(n_834),
.A2(n_311),
.B1(n_292),
.B2(n_301),
.Y(n_1016)
);

BUFx6f_ASAP7_75t_L g1017 ( 
.A(n_815),
.Y(n_1017)
);

BUFx3_ASAP7_75t_L g1018 ( 
.A(n_779),
.Y(n_1018)
);

NAND2xp5_ASAP7_75t_SL g1019 ( 
.A(n_862),
.B(n_242),
.Y(n_1019)
);

AOI22xp33_ASAP7_75t_L g1020 ( 
.A1(n_834),
.A2(n_311),
.B1(n_301),
.B2(n_306),
.Y(n_1020)
);

AOI22xp5_ASAP7_75t_L g1021 ( 
.A1(n_821),
.A2(n_419),
.B1(n_464),
.B2(n_311),
.Y(n_1021)
);

INVx2_ASAP7_75t_L g1022 ( 
.A(n_838),
.Y(n_1022)
);

INVx1_ASAP7_75t_L g1023 ( 
.A(n_730),
.Y(n_1023)
);

AOI22xp5_ASAP7_75t_L g1024 ( 
.A1(n_857),
.A2(n_246),
.B1(n_247),
.B2(n_244),
.Y(n_1024)
);

INVx1_ASAP7_75t_L g1025 ( 
.A(n_731),
.Y(n_1025)
);

NAND2xp5_ASAP7_75t_SL g1026 ( 
.A(n_855),
.B(n_248),
.Y(n_1026)
);

INVx2_ASAP7_75t_L g1027 ( 
.A(n_838),
.Y(n_1027)
);

NAND2xp5_ASAP7_75t_SL g1028 ( 
.A(n_750),
.B(n_249),
.Y(n_1028)
);

INVx2_ASAP7_75t_L g1029 ( 
.A(n_746),
.Y(n_1029)
);

NAND2xp5_ASAP7_75t_SL g1030 ( 
.A(n_750),
.B(n_250),
.Y(n_1030)
);

NAND2xp5_ASAP7_75t_L g1031 ( 
.A(n_815),
.B(n_311),
.Y(n_1031)
);

NAND2xp5_ASAP7_75t_L g1032 ( 
.A(n_828),
.B(n_311),
.Y(n_1032)
);

NAND2xp5_ASAP7_75t_SL g1033 ( 
.A(n_857),
.B(n_845),
.Y(n_1033)
);

A2O1A1Ixp33_ASAP7_75t_SL g1034 ( 
.A1(n_705),
.A2(n_448),
.B(n_306),
.C(n_309),
.Y(n_1034)
);

CKINVDCx5p33_ASAP7_75t_R g1035 ( 
.A(n_795),
.Y(n_1035)
);

O2A1O1Ixp5_ASAP7_75t_L g1036 ( 
.A1(n_807),
.A2(n_571),
.B(n_570),
.C(n_568),
.Y(n_1036)
);

INVx2_ASAP7_75t_L g1037 ( 
.A(n_746),
.Y(n_1037)
);

INVx1_ASAP7_75t_L g1038 ( 
.A(n_731),
.Y(n_1038)
);

NAND2xp5_ASAP7_75t_L g1039 ( 
.A(n_828),
.B(n_311),
.Y(n_1039)
);

INVx4_ASAP7_75t_L g1040 ( 
.A(n_873),
.Y(n_1040)
);

CKINVDCx5p33_ASAP7_75t_R g1041 ( 
.A(n_944),
.Y(n_1041)
);

NAND2xp5_ASAP7_75t_L g1042 ( 
.A(n_933),
.B(n_828),
.Y(n_1042)
);

INVx2_ASAP7_75t_L g1043 ( 
.A(n_885),
.Y(n_1043)
);

INVx2_ASAP7_75t_L g1044 ( 
.A(n_885),
.Y(n_1044)
);

INVx3_ASAP7_75t_L g1045 ( 
.A(n_873),
.Y(n_1045)
);

NOR2x1_ASAP7_75t_L g1046 ( 
.A(n_889),
.B(n_786),
.Y(n_1046)
);

NOR2xp33_ASAP7_75t_L g1047 ( 
.A(n_871),
.B(n_796),
.Y(n_1047)
);

NAND2xp5_ASAP7_75t_L g1048 ( 
.A(n_872),
.B(n_857),
.Y(n_1048)
);

NOR2xp33_ASAP7_75t_R g1049 ( 
.A(n_944),
.B(n_839),
.Y(n_1049)
);

NAND2xp5_ASAP7_75t_L g1050 ( 
.A(n_907),
.B(n_857),
.Y(n_1050)
);

AOI22xp33_ASAP7_75t_L g1051 ( 
.A1(n_866),
.A2(n_851),
.B1(n_833),
.B2(n_761),
.Y(n_1051)
);

NAND2xp5_ASAP7_75t_SL g1052 ( 
.A(n_873),
.B(n_761),
.Y(n_1052)
);

INVx5_ASAP7_75t_L g1053 ( 
.A(n_868),
.Y(n_1053)
);

AND2x2_ASAP7_75t_L g1054 ( 
.A(n_907),
.B(n_956),
.Y(n_1054)
);

BUFx2_ASAP7_75t_L g1055 ( 
.A(n_1018),
.Y(n_1055)
);

BUFx6f_ASAP7_75t_L g1056 ( 
.A(n_873),
.Y(n_1056)
);

INVx2_ASAP7_75t_L g1057 ( 
.A(n_890),
.Y(n_1057)
);

INVx3_ASAP7_75t_L g1058 ( 
.A(n_873),
.Y(n_1058)
);

CKINVDCx14_ASAP7_75t_R g1059 ( 
.A(n_967),
.Y(n_1059)
);

CKINVDCx6p67_ASAP7_75t_R g1060 ( 
.A(n_1018),
.Y(n_1060)
);

OR2x6_ASAP7_75t_L g1061 ( 
.A(n_919),
.B(n_804),
.Y(n_1061)
);

AOI22xp5_ASAP7_75t_L g1062 ( 
.A1(n_900),
.A2(n_753),
.B1(n_851),
.B2(n_809),
.Y(n_1062)
);

BUFx12f_ASAP7_75t_L g1063 ( 
.A(n_905),
.Y(n_1063)
);

AND2x2_ASAP7_75t_L g1064 ( 
.A(n_956),
.B(n_719),
.Y(n_1064)
);

AOI21xp5_ASAP7_75t_L g1065 ( 
.A1(n_868),
.A2(n_801),
.B(n_710),
.Y(n_1065)
);

AND2x2_ASAP7_75t_L g1066 ( 
.A(n_918),
.B(n_719),
.Y(n_1066)
);

BUFx6f_ASAP7_75t_L g1067 ( 
.A(n_875),
.Y(n_1067)
);

INVx1_ASAP7_75t_L g1068 ( 
.A(n_912),
.Y(n_1068)
);

NOR2xp33_ASAP7_75t_L g1069 ( 
.A(n_959),
.B(n_830),
.Y(n_1069)
);

INVx1_ASAP7_75t_L g1070 ( 
.A(n_912),
.Y(n_1070)
);

AND2x2_ASAP7_75t_L g1071 ( 
.A(n_918),
.B(n_719),
.Y(n_1071)
);

OR2x6_ASAP7_75t_L g1072 ( 
.A(n_919),
.B(n_847),
.Y(n_1072)
);

OR2x2_ASAP7_75t_L g1073 ( 
.A(n_920),
.B(n_840),
.Y(n_1073)
);

AND2x2_ASAP7_75t_L g1074 ( 
.A(n_923),
.B(n_742),
.Y(n_1074)
);

AND2x4_ASAP7_75t_SL g1075 ( 
.A(n_941),
.B(n_318),
.Y(n_1075)
);

AND2x2_ASAP7_75t_L g1076 ( 
.A(n_923),
.B(n_742),
.Y(n_1076)
);

NOR2xp33_ASAP7_75t_L g1077 ( 
.A(n_960),
.B(n_830),
.Y(n_1077)
);

AND3x1_ASAP7_75t_SL g1078 ( 
.A(n_942),
.B(n_309),
.C(n_285),
.Y(n_1078)
);

NOR2xp67_ASAP7_75t_L g1079 ( 
.A(n_967),
.B(n_863),
.Y(n_1079)
);

OAI221xp5_ASAP7_75t_L g1080 ( 
.A1(n_984),
.A2(n_459),
.B1(n_427),
.B2(n_414),
.C(n_409),
.Y(n_1080)
);

BUFx12f_ASAP7_75t_L g1081 ( 
.A(n_905),
.Y(n_1081)
);

BUFx3_ASAP7_75t_L g1082 ( 
.A(n_905),
.Y(n_1082)
);

BUFx3_ASAP7_75t_L g1083 ( 
.A(n_957),
.Y(n_1083)
);

INVx1_ASAP7_75t_L g1084 ( 
.A(n_976),
.Y(n_1084)
);

NOR2xp33_ASAP7_75t_R g1085 ( 
.A(n_1035),
.B(n_771),
.Y(n_1085)
);

NAND2xp5_ASAP7_75t_L g1086 ( 
.A(n_892),
.B(n_748),
.Y(n_1086)
);

INVx1_ASAP7_75t_L g1087 ( 
.A(n_976),
.Y(n_1087)
);

NAND2xp33_ASAP7_75t_SL g1088 ( 
.A(n_875),
.B(n_344),
.Y(n_1088)
);

INVx3_ASAP7_75t_L g1089 ( 
.A(n_875),
.Y(n_1089)
);

INVx4_ASAP7_75t_L g1090 ( 
.A(n_875),
.Y(n_1090)
);

INVx2_ASAP7_75t_SL g1091 ( 
.A(n_869),
.Y(n_1091)
);

INVx3_ASAP7_75t_L g1092 ( 
.A(n_875),
.Y(n_1092)
);

HB1xp67_ASAP7_75t_L g1093 ( 
.A(n_942),
.Y(n_1093)
);

HB1xp67_ASAP7_75t_L g1094 ( 
.A(n_973),
.Y(n_1094)
);

INVx3_ASAP7_75t_L g1095 ( 
.A(n_888),
.Y(n_1095)
);

INVx3_ASAP7_75t_L g1096 ( 
.A(n_888),
.Y(n_1096)
);

INVx1_ASAP7_75t_L g1097 ( 
.A(n_990),
.Y(n_1097)
);

NAND2xp5_ASAP7_75t_L g1098 ( 
.A(n_892),
.B(n_748),
.Y(n_1098)
);

INVx1_ASAP7_75t_L g1099 ( 
.A(n_990),
.Y(n_1099)
);

INVxp33_ASAP7_75t_L g1100 ( 
.A(n_978),
.Y(n_1100)
);

NAND2xp5_ASAP7_75t_L g1101 ( 
.A(n_901),
.B(n_751),
.Y(n_1101)
);

OR2x6_ASAP7_75t_L g1102 ( 
.A(n_919),
.B(n_830),
.Y(n_1102)
);

INVx1_ASAP7_75t_L g1103 ( 
.A(n_992),
.Y(n_1103)
);

AND2x2_ASAP7_75t_SL g1104 ( 
.A(n_982),
.B(n_344),
.Y(n_1104)
);

BUFx6f_ASAP7_75t_L g1105 ( 
.A(n_999),
.Y(n_1105)
);

INVx1_ASAP7_75t_L g1106 ( 
.A(n_992),
.Y(n_1106)
);

INVx2_ASAP7_75t_L g1107 ( 
.A(n_890),
.Y(n_1107)
);

NAND2xp5_ASAP7_75t_L g1108 ( 
.A(n_901),
.B(n_751),
.Y(n_1108)
);

INVx1_ASAP7_75t_L g1109 ( 
.A(n_1003),
.Y(n_1109)
);

NOR3xp33_ASAP7_75t_SL g1110 ( 
.A(n_911),
.B(n_257),
.C(n_255),
.Y(n_1110)
);

AND2x4_ASAP7_75t_L g1111 ( 
.A(n_997),
.B(n_703),
.Y(n_1111)
);

OR2x6_ASAP7_75t_L g1112 ( 
.A(n_919),
.B(n_830),
.Y(n_1112)
);

BUFx8_ASAP7_75t_L g1113 ( 
.A(n_973),
.Y(n_1113)
);

HB1xp67_ASAP7_75t_L g1114 ( 
.A(n_920),
.Y(n_1114)
);

INVx1_ASAP7_75t_L g1115 ( 
.A(n_1003),
.Y(n_1115)
);

AND2x4_ASAP7_75t_L g1116 ( 
.A(n_997),
.B(n_703),
.Y(n_1116)
);

NAND2xp5_ASAP7_75t_L g1117 ( 
.A(n_952),
.B(n_763),
.Y(n_1117)
);

INVxp67_ASAP7_75t_L g1118 ( 
.A(n_936),
.Y(n_1118)
);

NAND2xp5_ASAP7_75t_SL g1119 ( 
.A(n_868),
.B(n_830),
.Y(n_1119)
);

NOR2xp33_ASAP7_75t_L g1120 ( 
.A(n_921),
.B(n_262),
.Y(n_1120)
);

INVx1_ASAP7_75t_L g1121 ( 
.A(n_897),
.Y(n_1121)
);

OR2x4_ASAP7_75t_L g1122 ( 
.A(n_930),
.B(n_927),
.Y(n_1122)
);

AND3x1_ASAP7_75t_SL g1123 ( 
.A(n_938),
.B(n_361),
.C(n_346),
.Y(n_1123)
);

INVx2_ASAP7_75t_L g1124 ( 
.A(n_897),
.Y(n_1124)
);

INVx1_ASAP7_75t_L g1125 ( 
.A(n_898),
.Y(n_1125)
);

INVx1_ASAP7_75t_L g1126 ( 
.A(n_898),
.Y(n_1126)
);

INVx1_ASAP7_75t_SL g1127 ( 
.A(n_876),
.Y(n_1127)
);

AO22x1_ASAP7_75t_L g1128 ( 
.A1(n_970),
.A2(n_272),
.B1(n_273),
.B2(n_271),
.Y(n_1128)
);

INVx2_ASAP7_75t_L g1129 ( 
.A(n_922),
.Y(n_1129)
);

INVxp67_ASAP7_75t_L g1130 ( 
.A(n_955),
.Y(n_1130)
);

INVx1_ASAP7_75t_L g1131 ( 
.A(n_922),
.Y(n_1131)
);

HB1xp67_ASAP7_75t_L g1132 ( 
.A(n_989),
.Y(n_1132)
);

BUFx6f_ASAP7_75t_L g1133 ( 
.A(n_999),
.Y(n_1133)
);

HB1xp67_ASAP7_75t_L g1134 ( 
.A(n_989),
.Y(n_1134)
);

BUFx8_ASAP7_75t_L g1135 ( 
.A(n_958),
.Y(n_1135)
);

BUFx6f_ASAP7_75t_L g1136 ( 
.A(n_999),
.Y(n_1136)
);

HB1xp67_ASAP7_75t_L g1137 ( 
.A(n_869),
.Y(n_1137)
);

BUFx8_ASAP7_75t_L g1138 ( 
.A(n_958),
.Y(n_1138)
);

AND2x4_ASAP7_75t_SL g1139 ( 
.A(n_867),
.B(n_939),
.Y(n_1139)
);

INVx1_ASAP7_75t_L g1140 ( 
.A(n_947),
.Y(n_1140)
);

NAND2xp5_ASAP7_75t_L g1141 ( 
.A(n_952),
.B(n_763),
.Y(n_1141)
);

CKINVDCx6p67_ASAP7_75t_R g1142 ( 
.A(n_1004),
.Y(n_1142)
);

INVx1_ASAP7_75t_L g1143 ( 
.A(n_947),
.Y(n_1143)
);

AND2x2_ASAP7_75t_L g1144 ( 
.A(n_878),
.B(n_894),
.Y(n_1144)
);

NAND2xp5_ASAP7_75t_L g1145 ( 
.A(n_961),
.B(n_765),
.Y(n_1145)
);

INVx2_ASAP7_75t_L g1146 ( 
.A(n_948),
.Y(n_1146)
);

INVx3_ASAP7_75t_L g1147 ( 
.A(n_888),
.Y(n_1147)
);

NAND2xp5_ASAP7_75t_L g1148 ( 
.A(n_961),
.B(n_765),
.Y(n_1148)
);

INVx1_ASAP7_75t_L g1149 ( 
.A(n_948),
.Y(n_1149)
);

INVx2_ASAP7_75t_SL g1150 ( 
.A(n_878),
.Y(n_1150)
);

AOI22xp5_ASAP7_75t_SL g1151 ( 
.A1(n_1035),
.A2(n_279),
.B1(n_287),
.B2(n_275),
.Y(n_1151)
);

AND2x4_ASAP7_75t_L g1152 ( 
.A(n_998),
.B(n_712),
.Y(n_1152)
);

AND2x2_ASAP7_75t_L g1153 ( 
.A(n_894),
.B(n_766),
.Y(n_1153)
);

INVx3_ASAP7_75t_L g1154 ( 
.A(n_925),
.Y(n_1154)
);

INVx1_ASAP7_75t_L g1155 ( 
.A(n_950),
.Y(n_1155)
);

NOR2xp33_ASAP7_75t_R g1156 ( 
.A(n_916),
.B(n_931),
.Y(n_1156)
);

INVx2_ASAP7_75t_L g1157 ( 
.A(n_950),
.Y(n_1157)
);

INVx6_ASAP7_75t_L g1158 ( 
.A(n_999),
.Y(n_1158)
);

INVx1_ASAP7_75t_L g1159 ( 
.A(n_963),
.Y(n_1159)
);

OR2x2_ASAP7_75t_L g1160 ( 
.A(n_865),
.B(n_288),
.Y(n_1160)
);

INVx2_ASAP7_75t_L g1161 ( 
.A(n_963),
.Y(n_1161)
);

BUFx8_ASAP7_75t_L g1162 ( 
.A(n_958),
.Y(n_1162)
);

OAI22xp5_ASAP7_75t_L g1163 ( 
.A1(n_986),
.A2(n_768),
.B1(n_774),
.B2(n_766),
.Y(n_1163)
);

INVx1_ASAP7_75t_L g1164 ( 
.A(n_1009),
.Y(n_1164)
);

BUFx6f_ASAP7_75t_L g1165 ( 
.A(n_999),
.Y(n_1165)
);

AND2x6_ASAP7_75t_L g1166 ( 
.A(n_966),
.B(n_925),
.Y(n_1166)
);

INVx2_ASAP7_75t_L g1167 ( 
.A(n_874),
.Y(n_1167)
);

INVx1_ASAP7_75t_L g1168 ( 
.A(n_1009),
.Y(n_1168)
);

BUFx3_ASAP7_75t_L g1169 ( 
.A(n_957),
.Y(n_1169)
);

OR2x2_ASAP7_75t_L g1170 ( 
.A(n_865),
.B(n_291),
.Y(n_1170)
);

INVx3_ASAP7_75t_L g1171 ( 
.A(n_925),
.Y(n_1171)
);

INVx1_ASAP7_75t_L g1172 ( 
.A(n_1023),
.Y(n_1172)
);

INVx1_ASAP7_75t_L g1173 ( 
.A(n_1023),
.Y(n_1173)
);

INVx2_ASAP7_75t_L g1174 ( 
.A(n_874),
.Y(n_1174)
);

BUFx4f_ASAP7_75t_L g1175 ( 
.A(n_867),
.Y(n_1175)
);

AND2x4_ASAP7_75t_L g1176 ( 
.A(n_998),
.B(n_712),
.Y(n_1176)
);

AND2x4_ASAP7_75t_L g1177 ( 
.A(n_903),
.B(n_716),
.Y(n_1177)
);

INVx1_ASAP7_75t_SL g1178 ( 
.A(n_1028),
.Y(n_1178)
);

NAND2xp5_ASAP7_75t_L g1179 ( 
.A(n_966),
.B(n_768),
.Y(n_1179)
);

HB1xp67_ASAP7_75t_L g1180 ( 
.A(n_903),
.Y(n_1180)
);

NOR2xp33_ASAP7_75t_L g1181 ( 
.A(n_895),
.B(n_910),
.Y(n_1181)
);

CKINVDCx5p33_ASAP7_75t_R g1182 ( 
.A(n_957),
.Y(n_1182)
);

NAND2xp5_ASAP7_75t_L g1183 ( 
.A(n_937),
.B(n_774),
.Y(n_1183)
);

INVx3_ASAP7_75t_SL g1184 ( 
.A(n_1030),
.Y(n_1184)
);

NAND2xp5_ASAP7_75t_L g1185 ( 
.A(n_891),
.B(n_775),
.Y(n_1185)
);

NAND2xp5_ASAP7_75t_L g1186 ( 
.A(n_893),
.B(n_775),
.Y(n_1186)
);

INVx1_ASAP7_75t_L g1187 ( 
.A(n_1025),
.Y(n_1187)
);

NOR2xp33_ASAP7_75t_L g1188 ( 
.A(n_1012),
.B(n_294),
.Y(n_1188)
);

INVx2_ASAP7_75t_L g1189 ( 
.A(n_879),
.Y(n_1189)
);

INVx1_ASAP7_75t_L g1190 ( 
.A(n_1038),
.Y(n_1190)
);

INVx1_ASAP7_75t_L g1191 ( 
.A(n_1038),
.Y(n_1191)
);

BUFx12f_ASAP7_75t_L g1192 ( 
.A(n_867),
.Y(n_1192)
);

INVx1_ASAP7_75t_L g1193 ( 
.A(n_879),
.Y(n_1193)
);

INVx2_ASAP7_75t_L g1194 ( 
.A(n_968),
.Y(n_1194)
);

HB1xp67_ASAP7_75t_L g1195 ( 
.A(n_903),
.Y(n_1195)
);

NOR3xp33_ASAP7_75t_SL g1196 ( 
.A(n_965),
.B(n_304),
.C(n_295),
.Y(n_1196)
);

NAND2xp5_ASAP7_75t_L g1197 ( 
.A(n_929),
.B(n_781),
.Y(n_1197)
);

NOR3xp33_ASAP7_75t_SL g1198 ( 
.A(n_1026),
.B(n_312),
.C(n_310),
.Y(n_1198)
);

INVxp67_ASAP7_75t_SL g1199 ( 
.A(n_1017),
.Y(n_1199)
);

NAND2xp5_ASAP7_75t_SL g1200 ( 
.A(n_868),
.B(n_924),
.Y(n_1200)
);

AND2x2_ASAP7_75t_SL g1201 ( 
.A(n_934),
.B(n_346),
.Y(n_1201)
);

BUFx3_ASAP7_75t_L g1202 ( 
.A(n_1017),
.Y(n_1202)
);

BUFx3_ASAP7_75t_L g1203 ( 
.A(n_1017),
.Y(n_1203)
);

AND3x1_ASAP7_75t_L g1204 ( 
.A(n_915),
.B(n_378),
.C(n_361),
.Y(n_1204)
);

NOR3xp33_ASAP7_75t_SL g1205 ( 
.A(n_943),
.B(n_323),
.C(n_314),
.Y(n_1205)
);

NAND2xp5_ASAP7_75t_L g1206 ( 
.A(n_932),
.B(n_781),
.Y(n_1206)
);

HB1xp67_ASAP7_75t_L g1207 ( 
.A(n_940),
.Y(n_1207)
);

INVx2_ASAP7_75t_L g1208 ( 
.A(n_968),
.Y(n_1208)
);

NAND2xp5_ASAP7_75t_L g1209 ( 
.A(n_884),
.B(n_811),
.Y(n_1209)
);

CKINVDCx5p33_ASAP7_75t_R g1210 ( 
.A(n_870),
.Y(n_1210)
);

NAND2xp5_ASAP7_75t_SL g1211 ( 
.A(n_868),
.B(n_716),
.Y(n_1211)
);

INVx2_ASAP7_75t_L g1212 ( 
.A(n_1006),
.Y(n_1212)
);

BUFx4f_ASAP7_75t_L g1213 ( 
.A(n_867),
.Y(n_1213)
);

INVx1_ASAP7_75t_L g1214 ( 
.A(n_906),
.Y(n_1214)
);

INVx1_ASAP7_75t_L g1215 ( 
.A(n_908),
.Y(n_1215)
);

INVx2_ASAP7_75t_L g1216 ( 
.A(n_1006),
.Y(n_1216)
);

CKINVDCx5p33_ASAP7_75t_R g1217 ( 
.A(n_1021),
.Y(n_1217)
);

AOI22xp5_ASAP7_75t_L g1218 ( 
.A1(n_1033),
.A2(n_851),
.B1(n_816),
.B2(n_820),
.Y(n_1218)
);

INVx1_ASAP7_75t_SL g1219 ( 
.A(n_1019),
.Y(n_1219)
);

NAND2xp5_ASAP7_75t_SL g1220 ( 
.A(n_924),
.B(n_722),
.Y(n_1220)
);

OR2x6_ASAP7_75t_L g1221 ( 
.A(n_880),
.B(n_738),
.Y(n_1221)
);

INVx1_ASAP7_75t_L g1222 ( 
.A(n_913),
.Y(n_1222)
);

AOI22xp33_ASAP7_75t_L g1223 ( 
.A1(n_877),
.A2(n_851),
.B1(n_816),
.B2(n_820),
.Y(n_1223)
);

NOR2xp33_ASAP7_75t_L g1224 ( 
.A(n_951),
.B(n_325),
.Y(n_1224)
);

NAND2xp5_ASAP7_75t_L g1225 ( 
.A(n_883),
.B(n_811),
.Y(n_1225)
);

NOR2xp33_ASAP7_75t_L g1226 ( 
.A(n_988),
.B(n_326),
.Y(n_1226)
);

INVx5_ASAP7_75t_L g1227 ( 
.A(n_924),
.Y(n_1227)
);

AOI22xp5_ASAP7_75t_L g1228 ( 
.A1(n_914),
.A2(n_851),
.B1(n_825),
.B2(n_837),
.Y(n_1228)
);

INVx2_ASAP7_75t_L g1229 ( 
.A(n_1011),
.Y(n_1229)
);

BUFx6f_ASAP7_75t_L g1230 ( 
.A(n_1017),
.Y(n_1230)
);

NAND2xp5_ASAP7_75t_L g1231 ( 
.A(n_886),
.B(n_823),
.Y(n_1231)
);

AND2x4_ASAP7_75t_L g1232 ( 
.A(n_1017),
.B(n_722),
.Y(n_1232)
);

BUFx6f_ASAP7_75t_L g1233 ( 
.A(n_880),
.Y(n_1233)
);

INVx2_ASAP7_75t_SL g1234 ( 
.A(n_1055),
.Y(n_1234)
);

OAI21xp5_ASAP7_75t_L g1235 ( 
.A1(n_1066),
.A2(n_1071),
.B(n_1064),
.Y(n_1235)
);

INVx1_ASAP7_75t_L g1236 ( 
.A(n_1164),
.Y(n_1236)
);

OAI21x1_ASAP7_75t_L g1237 ( 
.A1(n_1065),
.A2(n_1032),
.B(n_1031),
.Y(n_1237)
);

NAND2xp5_ASAP7_75t_SL g1238 ( 
.A(n_1227),
.B(n_917),
.Y(n_1238)
);

BUFx2_ASAP7_75t_SL g1239 ( 
.A(n_1055),
.Y(n_1239)
);

AND2x4_ASAP7_75t_L g1240 ( 
.A(n_1144),
.B(n_991),
.Y(n_1240)
);

NAND2xp5_ASAP7_75t_L g1241 ( 
.A(n_1207),
.B(n_887),
.Y(n_1241)
);

NAND2xp5_ASAP7_75t_L g1242 ( 
.A(n_1047),
.B(n_1024),
.Y(n_1242)
);

NAND2xp5_ASAP7_75t_L g1243 ( 
.A(n_1144),
.B(n_1024),
.Y(n_1243)
);

INVx1_ASAP7_75t_L g1244 ( 
.A(n_1168),
.Y(n_1244)
);

NAND3xp33_ASAP7_75t_SL g1245 ( 
.A(n_1120),
.B(n_1005),
.C(n_996),
.Y(n_1245)
);

OAI21xp33_ASAP7_75t_L g1246 ( 
.A1(n_1100),
.A2(n_935),
.B(n_1008),
.Y(n_1246)
);

NAND2xp5_ASAP7_75t_L g1247 ( 
.A(n_1118),
.B(n_896),
.Y(n_1247)
);

INVx1_ASAP7_75t_L g1248 ( 
.A(n_1172),
.Y(n_1248)
);

AOI21xp5_ASAP7_75t_L g1249 ( 
.A1(n_1227),
.A2(n_1053),
.B(n_1200),
.Y(n_1249)
);

OAI21xp5_ASAP7_75t_L g1250 ( 
.A1(n_1066),
.A2(n_882),
.B(n_995),
.Y(n_1250)
);

OAI21xp5_ASAP7_75t_L g1251 ( 
.A1(n_1071),
.A2(n_899),
.B(n_975),
.Y(n_1251)
);

O2A1O1Ixp5_ASAP7_75t_L g1252 ( 
.A1(n_1188),
.A2(n_926),
.B(n_1042),
.C(n_1181),
.Y(n_1252)
);

CKINVDCx5p33_ASAP7_75t_R g1253 ( 
.A(n_1041),
.Y(n_1253)
);

NOR4xp25_ASAP7_75t_L g1254 ( 
.A(n_1080),
.B(n_1160),
.C(n_1170),
.D(n_1224),
.Y(n_1254)
);

INVx2_ASAP7_75t_L g1255 ( 
.A(n_1043),
.Y(n_1255)
);

BUFx6f_ASAP7_75t_L g1256 ( 
.A(n_1056),
.Y(n_1256)
);

NAND2xp5_ASAP7_75t_L g1257 ( 
.A(n_1091),
.B(n_1150),
.Y(n_1257)
);

NAND2xp5_ASAP7_75t_L g1258 ( 
.A(n_1091),
.B(n_902),
.Y(n_1258)
);

NAND2xp5_ASAP7_75t_L g1259 ( 
.A(n_1150),
.B(n_904),
.Y(n_1259)
);

AOI21xp5_ASAP7_75t_L g1260 ( 
.A1(n_1227),
.A2(n_979),
.B(n_801),
.Y(n_1260)
);

INVx3_ASAP7_75t_L g1261 ( 
.A(n_1040),
.Y(n_1261)
);

NAND2xp5_ASAP7_75t_L g1262 ( 
.A(n_1132),
.B(n_981),
.Y(n_1262)
);

NAND2xp5_ASAP7_75t_L g1263 ( 
.A(n_1134),
.B(n_983),
.Y(n_1263)
);

AND2x2_ASAP7_75t_L g1264 ( 
.A(n_1100),
.B(n_928),
.Y(n_1264)
);

OAI21x1_ASAP7_75t_L g1265 ( 
.A1(n_1209),
.A2(n_1039),
.B(n_1010),
.Y(n_1265)
);

OAI21x1_ASAP7_75t_L g1266 ( 
.A1(n_1052),
.A2(n_1007),
.B(n_880),
.Y(n_1266)
);

BUFx2_ASAP7_75t_L g1267 ( 
.A(n_1113),
.Y(n_1267)
);

NAND2xp5_ASAP7_75t_L g1268 ( 
.A(n_1054),
.B(n_980),
.Y(n_1268)
);

OAI21xp33_ASAP7_75t_L g1269 ( 
.A1(n_1104),
.A2(n_1002),
.B(n_1000),
.Y(n_1269)
);

A2O1A1Ixp33_ASAP7_75t_L g1270 ( 
.A1(n_1104),
.A2(n_949),
.B(n_974),
.C(n_971),
.Y(n_1270)
);

OAI21x1_ASAP7_75t_L g1271 ( 
.A1(n_1052),
.A2(n_1014),
.B(n_953),
.Y(n_1271)
);

AND2x4_ASAP7_75t_L g1272 ( 
.A(n_1180),
.B(n_1011),
.Y(n_1272)
);

NAND2xp5_ASAP7_75t_L g1273 ( 
.A(n_1054),
.B(n_987),
.Y(n_1273)
);

NOR2xp33_ASAP7_75t_L g1274 ( 
.A(n_1217),
.B(n_945),
.Y(n_1274)
);

AOI22xp5_ASAP7_75t_L g1275 ( 
.A1(n_1217),
.A2(n_946),
.B1(n_994),
.B2(n_993),
.Y(n_1275)
);

OAI21xp5_ASAP7_75t_L g1276 ( 
.A1(n_1064),
.A2(n_962),
.B(n_954),
.Y(n_1276)
);

BUFx2_ASAP7_75t_L g1277 ( 
.A(n_1113),
.Y(n_1277)
);

INVxp67_ASAP7_75t_L g1278 ( 
.A(n_1114),
.Y(n_1278)
);

NAND2xp5_ASAP7_75t_L g1279 ( 
.A(n_1214),
.B(n_964),
.Y(n_1279)
);

OR2x2_ASAP7_75t_L g1280 ( 
.A(n_1094),
.B(n_1013),
.Y(n_1280)
);

OAI21xp5_ASAP7_75t_L g1281 ( 
.A1(n_1048),
.A2(n_972),
.B(n_969),
.Y(n_1281)
);

BUFx6f_ASAP7_75t_L g1282 ( 
.A(n_1056),
.Y(n_1282)
);

CKINVDCx8_ASAP7_75t_R g1283 ( 
.A(n_1041),
.Y(n_1283)
);

BUFx3_ASAP7_75t_L g1284 ( 
.A(n_1060),
.Y(n_1284)
);

OAI21x1_ASAP7_75t_SL g1285 ( 
.A1(n_1040),
.A2(n_1020),
.B(n_1016),
.Y(n_1285)
);

NAND2xp5_ASAP7_75t_L g1286 ( 
.A(n_1215),
.B(n_1037),
.Y(n_1286)
);

CKINVDCx11_ASAP7_75t_R g1287 ( 
.A(n_1063),
.Y(n_1287)
);

OAI22xp5_ASAP7_75t_L g1288 ( 
.A1(n_1222),
.A2(n_1013),
.B1(n_1027),
.B2(n_1022),
.Y(n_1288)
);

NAND2xp5_ASAP7_75t_L g1289 ( 
.A(n_1153),
.B(n_1022),
.Y(n_1289)
);

AOI22xp5_ASAP7_75t_L g1290 ( 
.A1(n_1142),
.A2(n_946),
.B1(n_851),
.B2(n_1027),
.Y(n_1290)
);

NAND2xp5_ASAP7_75t_L g1291 ( 
.A(n_1153),
.B(n_1037),
.Y(n_1291)
);

NAND2xp5_ASAP7_75t_L g1292 ( 
.A(n_1137),
.B(n_1029),
.Y(n_1292)
);

OAI21xp5_ASAP7_75t_L g1293 ( 
.A1(n_1050),
.A2(n_1029),
.B(n_909),
.Y(n_1293)
);

BUFx6f_ASAP7_75t_L g1294 ( 
.A(n_1056),
.Y(n_1294)
);

NAND2xp5_ASAP7_75t_L g1295 ( 
.A(n_1074),
.B(n_823),
.Y(n_1295)
);

NAND2xp5_ASAP7_75t_L g1296 ( 
.A(n_1074),
.B(n_825),
.Y(n_1296)
);

NAND2xp5_ASAP7_75t_L g1297 ( 
.A(n_1076),
.B(n_837),
.Y(n_1297)
);

INVx1_ASAP7_75t_SL g1298 ( 
.A(n_1049),
.Y(n_1298)
);

OAI21x1_ASAP7_75t_L g1299 ( 
.A1(n_1200),
.A2(n_1036),
.B(n_1015),
.Y(n_1299)
);

INVx2_ASAP7_75t_L g1300 ( 
.A(n_1043),
.Y(n_1300)
);

AOI21xp5_ASAP7_75t_L g1301 ( 
.A1(n_1227),
.A2(n_801),
.B(n_710),
.Y(n_1301)
);

NAND2xp5_ASAP7_75t_L g1302 ( 
.A(n_1076),
.B(n_985),
.Y(n_1302)
);

OAI21x1_ASAP7_75t_L g1303 ( 
.A1(n_1220),
.A2(n_729),
.B(n_726),
.Y(n_1303)
);

INVxp67_ASAP7_75t_L g1304 ( 
.A(n_1093),
.Y(n_1304)
);

INVx1_ASAP7_75t_L g1305 ( 
.A(n_1173),
.Y(n_1305)
);

INVx3_ASAP7_75t_L g1306 ( 
.A(n_1040),
.Y(n_1306)
);

BUFx8_ASAP7_75t_SL g1307 ( 
.A(n_1063),
.Y(n_1307)
);

INVx4_ASAP7_75t_L g1308 ( 
.A(n_1056),
.Y(n_1308)
);

INVxp67_ASAP7_75t_SL g1309 ( 
.A(n_1056),
.Y(n_1309)
);

NAND2xp5_ASAP7_75t_L g1310 ( 
.A(n_1195),
.B(n_881),
.Y(n_1310)
);

OAI22xp5_ASAP7_75t_L g1311 ( 
.A1(n_1139),
.A2(n_977),
.B1(n_726),
.B2(n_705),
.Y(n_1311)
);

OAI21x1_ASAP7_75t_L g1312 ( 
.A1(n_1220),
.A2(n_729),
.B(n_726),
.Y(n_1312)
);

AND2x4_ASAP7_75t_L g1313 ( 
.A(n_1202),
.B(n_771),
.Y(n_1313)
);

AOI21xp5_ASAP7_75t_L g1314 ( 
.A1(n_1227),
.A2(n_710),
.B(n_708),
.Y(n_1314)
);

NAND2xp5_ASAP7_75t_L g1315 ( 
.A(n_1069),
.B(n_1077),
.Y(n_1315)
);

NOR2x1_ASAP7_75t_SL g1316 ( 
.A(n_1067),
.B(n_770),
.Y(n_1316)
);

OAI21x1_ASAP7_75t_L g1317 ( 
.A1(n_1119),
.A2(n_726),
.B(n_705),
.Y(n_1317)
);

INVx1_ASAP7_75t_L g1318 ( 
.A(n_1187),
.Y(n_1318)
);

INVx1_ASAP7_75t_L g1319 ( 
.A(n_1190),
.Y(n_1319)
);

AOI21xp5_ASAP7_75t_L g1320 ( 
.A1(n_1053),
.A2(n_1183),
.B(n_1221),
.Y(n_1320)
);

NOR2xp67_ASAP7_75t_L g1321 ( 
.A(n_1130),
.B(n_127),
.Y(n_1321)
);

NAND2xp5_ASAP7_75t_L g1322 ( 
.A(n_1197),
.B(n_881),
.Y(n_1322)
);

NAND2xp5_ASAP7_75t_L g1323 ( 
.A(n_1206),
.B(n_836),
.Y(n_1323)
);

NAND2xp5_ASAP7_75t_L g1324 ( 
.A(n_1191),
.B(n_1068),
.Y(n_1324)
);

A2O1A1Ixp33_ASAP7_75t_L g1325 ( 
.A1(n_1139),
.A2(n_400),
.B(n_409),
.C(n_378),
.Y(n_1325)
);

NOR2x1_ASAP7_75t_L g1326 ( 
.A(n_1046),
.B(n_705),
.Y(n_1326)
);

NAND2xp5_ASAP7_75t_L g1327 ( 
.A(n_1070),
.B(n_755),
.Y(n_1327)
);

AOI21x1_ASAP7_75t_L g1328 ( 
.A1(n_1086),
.A2(n_1001),
.B(n_757),
.Y(n_1328)
);

OAI22xp5_ASAP7_75t_L g1329 ( 
.A1(n_1142),
.A2(n_789),
.B1(n_790),
.B2(n_771),
.Y(n_1329)
);

INVx2_ASAP7_75t_L g1330 ( 
.A(n_1044),
.Y(n_1330)
);

INVx2_ASAP7_75t_L g1331 ( 
.A(n_1044),
.Y(n_1331)
);

OAI21x1_ASAP7_75t_L g1332 ( 
.A1(n_1119),
.A2(n_789),
.B(n_771),
.Y(n_1332)
);

OAI21xp5_ASAP7_75t_L g1333 ( 
.A1(n_1062),
.A2(n_757),
.B(n_755),
.Y(n_1333)
);

INVx3_ASAP7_75t_L g1334 ( 
.A(n_1090),
.Y(n_1334)
);

INVx3_ASAP7_75t_L g1335 ( 
.A(n_1090),
.Y(n_1335)
);

AOI21x1_ASAP7_75t_SL g1336 ( 
.A1(n_1185),
.A2(n_1001),
.B(n_1034),
.Y(n_1336)
);

AOI21xp5_ASAP7_75t_L g1337 ( 
.A1(n_1053),
.A2(n_710),
.B(n_708),
.Y(n_1337)
);

AOI221x1_ASAP7_75t_L g1338 ( 
.A1(n_1088),
.A2(n_427),
.B1(n_400),
.B2(n_429),
.C(n_431),
.Y(n_1338)
);

BUFx6f_ASAP7_75t_L g1339 ( 
.A(n_1067),
.Y(n_1339)
);

A2O1A1Ixp33_ASAP7_75t_L g1340 ( 
.A1(n_1201),
.A2(n_414),
.B(n_429),
.C(n_431),
.Y(n_1340)
);

AND3x4_ASAP7_75t_L g1341 ( 
.A(n_1198),
.B(n_318),
.C(n_336),
.Y(n_1341)
);

OAI21xp5_ASAP7_75t_L g1342 ( 
.A1(n_1228),
.A2(n_769),
.B(n_758),
.Y(n_1342)
);

OAI21xp5_ASAP7_75t_L g1343 ( 
.A1(n_1186),
.A2(n_1218),
.B(n_1225),
.Y(n_1343)
);

INVx1_ASAP7_75t_L g1344 ( 
.A(n_1057),
.Y(n_1344)
);

OAI22x1_ASAP7_75t_L g1345 ( 
.A1(n_1210),
.A2(n_339),
.B1(n_337),
.B2(n_343),
.Y(n_1345)
);

INVx1_ASAP7_75t_L g1346 ( 
.A(n_1057),
.Y(n_1346)
);

A2O1A1Ixp33_ASAP7_75t_L g1347 ( 
.A1(n_1201),
.A2(n_459),
.B(n_432),
.C(n_433),
.Y(n_1347)
);

AND2x2_ASAP7_75t_L g1348 ( 
.A(n_1127),
.B(n_1073),
.Y(n_1348)
);

AOI21x1_ASAP7_75t_L g1349 ( 
.A1(n_1098),
.A2(n_769),
.B(n_758),
.Y(n_1349)
);

AOI21xp5_ASAP7_75t_L g1350 ( 
.A1(n_1053),
.A2(n_1221),
.B(n_1090),
.Y(n_1350)
);

NAND2xp5_ASAP7_75t_SL g1351 ( 
.A(n_1067),
.B(n_1156),
.Y(n_1351)
);

AOI21xp5_ASAP7_75t_L g1352 ( 
.A1(n_1053),
.A2(n_714),
.B(n_708),
.Y(n_1352)
);

BUFx2_ASAP7_75t_SL g1353 ( 
.A(n_1082),
.Y(n_1353)
);

INVx4_ASAP7_75t_L g1354 ( 
.A(n_1067),
.Y(n_1354)
);

AOI21xp5_ASAP7_75t_L g1355 ( 
.A1(n_1221),
.A2(n_714),
.B(n_708),
.Y(n_1355)
);

OAI21xp5_ASAP7_75t_L g1356 ( 
.A1(n_1231),
.A2(n_780),
.B(n_777),
.Y(n_1356)
);

NOR2xp67_ASAP7_75t_L g1357 ( 
.A(n_1081),
.B(n_131),
.Y(n_1357)
);

INVxp67_ASAP7_75t_SL g1358 ( 
.A(n_1136),
.Y(n_1358)
);

AOI21xp5_ASAP7_75t_L g1359 ( 
.A1(n_1221),
.A2(n_714),
.B(n_738),
.Y(n_1359)
);

OAI21x1_ASAP7_75t_L g1360 ( 
.A1(n_1211),
.A2(n_790),
.B(n_789),
.Y(n_1360)
);

BUFx3_ASAP7_75t_L g1361 ( 
.A(n_1060),
.Y(n_1361)
);

A2O1A1Ixp33_ASAP7_75t_L g1362 ( 
.A1(n_1226),
.A2(n_432),
.B(n_433),
.C(n_434),
.Y(n_1362)
);

BUFx3_ASAP7_75t_L g1363 ( 
.A(n_1135),
.Y(n_1363)
);

NOR2xp33_ASAP7_75t_L g1364 ( 
.A(n_1122),
.B(n_347),
.Y(n_1364)
);

INVx1_ASAP7_75t_L g1365 ( 
.A(n_1107),
.Y(n_1365)
);

INVx3_ASAP7_75t_L g1366 ( 
.A(n_1095),
.Y(n_1366)
);

NAND2xp5_ASAP7_75t_L g1367 ( 
.A(n_1107),
.B(n_780),
.Y(n_1367)
);

NAND2xp5_ASAP7_75t_L g1368 ( 
.A(n_1124),
.B(n_817),
.Y(n_1368)
);

NAND2xp5_ASAP7_75t_SL g1369 ( 
.A(n_1233),
.B(n_789),
.Y(n_1369)
);

OAI21xp5_ASAP7_75t_L g1370 ( 
.A1(n_1163),
.A2(n_818),
.B(n_817),
.Y(n_1370)
);

NOR2xp33_ASAP7_75t_L g1371 ( 
.A(n_1122),
.B(n_348),
.Y(n_1371)
);

OAI21x1_ASAP7_75t_L g1372 ( 
.A1(n_1211),
.A2(n_794),
.B(n_790),
.Y(n_1372)
);

AOI21xp5_ASAP7_75t_L g1373 ( 
.A1(n_1199),
.A2(n_1096),
.B(n_1095),
.Y(n_1373)
);

NAND3xp33_ASAP7_75t_L g1374 ( 
.A(n_1110),
.B(n_1151),
.C(n_1196),
.Y(n_1374)
);

INVx1_ASAP7_75t_L g1375 ( 
.A(n_1124),
.Y(n_1375)
);

OAI21x1_ASAP7_75t_L g1376 ( 
.A1(n_1101),
.A2(n_794),
.B(n_790),
.Y(n_1376)
);

NAND2xp5_ASAP7_75t_L g1377 ( 
.A(n_1129),
.B(n_818),
.Y(n_1377)
);

OAI21x1_ASAP7_75t_L g1378 ( 
.A1(n_1108),
.A2(n_799),
.B(n_794),
.Y(n_1378)
);

INVx1_ASAP7_75t_L g1379 ( 
.A(n_1129),
.Y(n_1379)
);

NAND2xp5_ASAP7_75t_L g1380 ( 
.A(n_1146),
.B(n_794),
.Y(n_1380)
);

NAND2xp5_ASAP7_75t_L g1381 ( 
.A(n_1146),
.B(n_799),
.Y(n_1381)
);

BUFx2_ASAP7_75t_L g1382 ( 
.A(n_1113),
.Y(n_1382)
);

AO21x2_ASAP7_75t_L g1383 ( 
.A1(n_1117),
.A2(n_539),
.B(n_533),
.Y(n_1383)
);

INVxp67_ASAP7_75t_L g1384 ( 
.A(n_1178),
.Y(n_1384)
);

NOR2xp33_ASAP7_75t_L g1385 ( 
.A(n_1160),
.B(n_350),
.Y(n_1385)
);

NAND2xp5_ASAP7_75t_L g1386 ( 
.A(n_1157),
.B(n_799),
.Y(n_1386)
);

NAND2xp33_ASAP7_75t_SL g1387 ( 
.A(n_1233),
.B(n_770),
.Y(n_1387)
);

OAI21x1_ASAP7_75t_L g1388 ( 
.A1(n_1141),
.A2(n_803),
.B(n_799),
.Y(n_1388)
);

INVx2_ASAP7_75t_SL g1389 ( 
.A(n_1075),
.Y(n_1389)
);

INVx1_ASAP7_75t_L g1390 ( 
.A(n_1157),
.Y(n_1390)
);

OAI21x1_ASAP7_75t_L g1391 ( 
.A1(n_1145),
.A2(n_805),
.B(n_803),
.Y(n_1391)
);

NAND2xp5_ASAP7_75t_SL g1392 ( 
.A(n_1233),
.B(n_803),
.Y(n_1392)
);

NAND2xp5_ASAP7_75t_L g1393 ( 
.A(n_1161),
.B(n_803),
.Y(n_1393)
);

OAI21x1_ASAP7_75t_L g1394 ( 
.A1(n_1148),
.A2(n_805),
.B(n_542),
.Y(n_1394)
);

NOR2xp67_ASAP7_75t_L g1395 ( 
.A(n_1081),
.B(n_134),
.Y(n_1395)
);

NAND2x1_ASAP7_75t_L g1396 ( 
.A(n_1166),
.B(n_714),
.Y(n_1396)
);

AOI21xp5_ASAP7_75t_L g1397 ( 
.A1(n_1095),
.A2(n_754),
.B(n_738),
.Y(n_1397)
);

AND2x4_ASAP7_75t_L g1398 ( 
.A(n_1202),
.B(n_805),
.Y(n_1398)
);

INVx4_ASAP7_75t_L g1399 ( 
.A(n_1136),
.Y(n_1399)
);

INVx3_ASAP7_75t_L g1400 ( 
.A(n_1096),
.Y(n_1400)
);

AO32x2_ASAP7_75t_L g1401 ( 
.A1(n_1078),
.A2(n_783),
.A3(n_754),
.B1(n_738),
.B2(n_832),
.Y(n_1401)
);

A2O1A1Ixp33_ASAP7_75t_L g1402 ( 
.A1(n_1242),
.A2(n_1175),
.B(n_1213),
.C(n_1205),
.Y(n_1402)
);

AOI22xp33_ASAP7_75t_L g1403 ( 
.A1(n_1385),
.A2(n_1210),
.B1(n_1170),
.B2(n_1061),
.Y(n_1403)
);

NAND2xp5_ASAP7_75t_L g1404 ( 
.A(n_1274),
.B(n_1079),
.Y(n_1404)
);

AOI22xp33_ASAP7_75t_L g1405 ( 
.A1(n_1385),
.A2(n_1061),
.B1(n_1192),
.B2(n_1219),
.Y(n_1405)
);

INVx1_ASAP7_75t_L g1406 ( 
.A(n_1255),
.Y(n_1406)
);

AOI22xp33_ASAP7_75t_L g1407 ( 
.A1(n_1348),
.A2(n_1061),
.B1(n_1192),
.B2(n_1175),
.Y(n_1407)
);

INVx3_ASAP7_75t_L g1408 ( 
.A(n_1261),
.Y(n_1408)
);

OAI21x1_ASAP7_75t_L g1409 ( 
.A1(n_1376),
.A2(n_1179),
.B(n_1161),
.Y(n_1409)
);

OAI21xp5_ASAP7_75t_L g1410 ( 
.A1(n_1252),
.A2(n_1250),
.B(n_1251),
.Y(n_1410)
);

INVx2_ASAP7_75t_L g1411 ( 
.A(n_1300),
.Y(n_1411)
);

O2A1O1Ixp33_ASAP7_75t_L g1412 ( 
.A1(n_1340),
.A2(n_1184),
.B(n_1061),
.C(n_1059),
.Y(n_1412)
);

AND2x2_ASAP7_75t_L g1413 ( 
.A(n_1235),
.B(n_1121),
.Y(n_1413)
);

AOI222xp33_ASAP7_75t_L g1414 ( 
.A1(n_1269),
.A2(n_1128),
.B1(n_318),
.B2(n_448),
.C1(n_454),
.C2(n_466),
.Y(n_1414)
);

AND2x4_ASAP7_75t_L g1415 ( 
.A(n_1240),
.B(n_1203),
.Y(n_1415)
);

AO32x2_ASAP7_75t_L g1416 ( 
.A1(n_1311),
.A2(n_1204),
.A3(n_1088),
.B1(n_1175),
.B2(n_1213),
.Y(n_1416)
);

NOR2x1_ASAP7_75t_SL g1417 ( 
.A(n_1238),
.B(n_1233),
.Y(n_1417)
);

INVx1_ASAP7_75t_L g1418 ( 
.A(n_1300),
.Y(n_1418)
);

AO21x1_ASAP7_75t_L g1419 ( 
.A1(n_1322),
.A2(n_1126),
.B(n_1125),
.Y(n_1419)
);

AOI22xp33_ASAP7_75t_L g1420 ( 
.A1(n_1245),
.A2(n_1213),
.B1(n_1138),
.B2(n_1162),
.Y(n_1420)
);

OAI21xp5_ASAP7_75t_L g1421 ( 
.A1(n_1343),
.A2(n_1223),
.B(n_1051),
.Y(n_1421)
);

INVx2_ASAP7_75t_L g1422 ( 
.A(n_1330),
.Y(n_1422)
);

INVx1_ASAP7_75t_L g1423 ( 
.A(n_1330),
.Y(n_1423)
);

OA21x2_ASAP7_75t_L g1424 ( 
.A1(n_1394),
.A2(n_1140),
.B(n_1131),
.Y(n_1424)
);

AOI22x1_ASAP7_75t_L g1425 ( 
.A1(n_1281),
.A2(n_1143),
.B1(n_1155),
.B2(n_1149),
.Y(n_1425)
);

INVx2_ASAP7_75t_L g1426 ( 
.A(n_1331),
.Y(n_1426)
);

AO21x2_ASAP7_75t_L g1427 ( 
.A1(n_1376),
.A2(n_1159),
.B(n_1087),
.Y(n_1427)
);

NAND2xp5_ASAP7_75t_L g1428 ( 
.A(n_1274),
.B(n_1085),
.Y(n_1428)
);

AOI21xp5_ASAP7_75t_L g1429 ( 
.A1(n_1315),
.A2(n_1233),
.B(n_1112),
.Y(n_1429)
);

OAI21x1_ASAP7_75t_L g1430 ( 
.A1(n_1378),
.A2(n_1391),
.B(n_1388),
.Y(n_1430)
);

NAND2xp5_ASAP7_75t_L g1431 ( 
.A(n_1241),
.B(n_1247),
.Y(n_1431)
);

HB1xp67_ASAP7_75t_L g1432 ( 
.A(n_1278),
.Y(n_1432)
);

OAI21x1_ASAP7_75t_SL g1433 ( 
.A1(n_1350),
.A2(n_1097),
.B(n_1084),
.Y(n_1433)
);

AND2x2_ASAP7_75t_L g1434 ( 
.A(n_1240),
.B(n_1177),
.Y(n_1434)
);

AOI22xp33_ASAP7_75t_L g1435 ( 
.A1(n_1374),
.A2(n_1138),
.B1(n_1162),
.B2(n_1135),
.Y(n_1435)
);

OAI21x1_ASAP7_75t_L g1436 ( 
.A1(n_1378),
.A2(n_1147),
.B(n_1096),
.Y(n_1436)
);

AND2x2_ASAP7_75t_L g1437 ( 
.A(n_1240),
.B(n_1177),
.Y(n_1437)
);

O2A1O1Ixp33_ASAP7_75t_SL g1438 ( 
.A1(n_1270),
.A2(n_1103),
.B(n_1106),
.C(n_1099),
.Y(n_1438)
);

OAI21x1_ASAP7_75t_L g1439 ( 
.A1(n_1388),
.A2(n_1154),
.B(n_1147),
.Y(n_1439)
);

INVx1_ASAP7_75t_L g1440 ( 
.A(n_1331),
.Y(n_1440)
);

OAI21x1_ASAP7_75t_L g1441 ( 
.A1(n_1391),
.A2(n_1394),
.B(n_1332),
.Y(n_1441)
);

OAI221xp5_ASAP7_75t_L g1442 ( 
.A1(n_1254),
.A2(n_1184),
.B1(n_1082),
.B2(n_1083),
.C(n_1169),
.Y(n_1442)
);

AOI22xp33_ASAP7_75t_L g1443 ( 
.A1(n_1246),
.A2(n_1138),
.B1(n_1162),
.B2(n_1135),
.Y(n_1443)
);

OAI21x1_ASAP7_75t_L g1444 ( 
.A1(n_1332),
.A2(n_1154),
.B(n_1147),
.Y(n_1444)
);

OR2x6_ASAP7_75t_L g1445 ( 
.A(n_1351),
.B(n_1102),
.Y(n_1445)
);

OAI21x1_ASAP7_75t_L g1446 ( 
.A1(n_1237),
.A2(n_1171),
.B(n_1154),
.Y(n_1446)
);

OAI22xp33_ASAP7_75t_L g1447 ( 
.A1(n_1243),
.A2(n_1182),
.B1(n_1169),
.B2(n_1083),
.Y(n_1447)
);

AND2x2_ASAP7_75t_L g1448 ( 
.A(n_1268),
.B(n_1177),
.Y(n_1448)
);

OAI21x1_ASAP7_75t_L g1449 ( 
.A1(n_1237),
.A2(n_1171),
.B(n_1167),
.Y(n_1449)
);

AOI22xp33_ASAP7_75t_L g1450 ( 
.A1(n_1364),
.A2(n_1371),
.B1(n_1264),
.B2(n_1345),
.Y(n_1450)
);

AOI21xp5_ASAP7_75t_L g1451 ( 
.A1(n_1320),
.A2(n_1112),
.B(n_1102),
.Y(n_1451)
);

OAI21x1_ASAP7_75t_L g1452 ( 
.A1(n_1317),
.A2(n_1171),
.B(n_1167),
.Y(n_1452)
);

INVx1_ASAP7_75t_L g1453 ( 
.A(n_1344),
.Y(n_1453)
);

INVx2_ASAP7_75t_SL g1454 ( 
.A(n_1339),
.Y(n_1454)
);

INVx2_ASAP7_75t_L g1455 ( 
.A(n_1346),
.Y(n_1455)
);

INVx1_ASAP7_75t_L g1456 ( 
.A(n_1365),
.Y(n_1456)
);

BUFx6f_ASAP7_75t_L g1457 ( 
.A(n_1256),
.Y(n_1457)
);

INVx1_ASAP7_75t_L g1458 ( 
.A(n_1375),
.Y(n_1458)
);

INVx1_ASAP7_75t_L g1459 ( 
.A(n_1379),
.Y(n_1459)
);

NAND2xp5_ASAP7_75t_L g1460 ( 
.A(n_1273),
.B(n_1174),
.Y(n_1460)
);

OAI21x1_ASAP7_75t_L g1461 ( 
.A1(n_1317),
.A2(n_1189),
.B(n_1174),
.Y(n_1461)
);

INVx2_ASAP7_75t_L g1462 ( 
.A(n_1390),
.Y(n_1462)
);

OAI21x1_ASAP7_75t_L g1463 ( 
.A1(n_1349),
.A2(n_1189),
.B(n_1194),
.Y(n_1463)
);

NAND2xp5_ASAP7_75t_L g1464 ( 
.A(n_1279),
.B(n_1193),
.Y(n_1464)
);

NAND2x1p5_ASAP7_75t_L g1465 ( 
.A(n_1261),
.B(n_1045),
.Y(n_1465)
);

AOI31xp67_ASAP7_75t_L g1466 ( 
.A1(n_1238),
.A2(n_1208),
.A3(n_1194),
.B(n_1229),
.Y(n_1466)
);

NOR2xp33_ASAP7_75t_L g1467 ( 
.A(n_1298),
.B(n_1059),
.Y(n_1467)
);

NOR2x1_ASAP7_75t_R g1468 ( 
.A(n_1253),
.B(n_1182),
.Y(n_1468)
);

INVx4_ASAP7_75t_L g1469 ( 
.A(n_1339),
.Y(n_1469)
);

OAI21x1_ASAP7_75t_L g1470 ( 
.A1(n_1360),
.A2(n_1372),
.B(n_1266),
.Y(n_1470)
);

OAI21x1_ASAP7_75t_L g1471 ( 
.A1(n_1360),
.A2(n_1372),
.B(n_1266),
.Y(n_1471)
);

AO21x2_ASAP7_75t_L g1472 ( 
.A1(n_1333),
.A2(n_1115),
.B(n_1109),
.Y(n_1472)
);

OAI21x1_ASAP7_75t_L g1473 ( 
.A1(n_1303),
.A2(n_1212),
.B(n_1208),
.Y(n_1473)
);

INVx3_ASAP7_75t_L g1474 ( 
.A(n_1261),
.Y(n_1474)
);

AO31x2_ASAP7_75t_L g1475 ( 
.A1(n_1338),
.A2(n_1212),
.A3(n_1216),
.B(n_1229),
.Y(n_1475)
);

NAND2xp5_ASAP7_75t_L g1476 ( 
.A(n_1258),
.B(n_1111),
.Y(n_1476)
);

OAI21x1_ASAP7_75t_L g1477 ( 
.A1(n_1303),
.A2(n_1216),
.B(n_1058),
.Y(n_1477)
);

HB1xp67_ASAP7_75t_L g1478 ( 
.A(n_1234),
.Y(n_1478)
);

BUFx2_ASAP7_75t_SL g1479 ( 
.A(n_1283),
.Y(n_1479)
);

INVx1_ASAP7_75t_L g1480 ( 
.A(n_1289),
.Y(n_1480)
);

NAND2xp5_ASAP7_75t_L g1481 ( 
.A(n_1259),
.B(n_1111),
.Y(n_1481)
);

BUFx6f_ASAP7_75t_L g1482 ( 
.A(n_1256),
.Y(n_1482)
);

INVx3_ASAP7_75t_L g1483 ( 
.A(n_1306),
.Y(n_1483)
);

OAI21x1_ASAP7_75t_L g1484 ( 
.A1(n_1312),
.A2(n_1058),
.B(n_1045),
.Y(n_1484)
);

OAI21x1_ASAP7_75t_L g1485 ( 
.A1(n_1312),
.A2(n_1058),
.B(n_1045),
.Y(n_1485)
);

INVx1_ASAP7_75t_L g1486 ( 
.A(n_1291),
.Y(n_1486)
);

AOI21xp5_ASAP7_75t_L g1487 ( 
.A1(n_1323),
.A2(n_1112),
.B(n_1102),
.Y(n_1487)
);

INVx3_ASAP7_75t_L g1488 ( 
.A(n_1306),
.Y(n_1488)
);

NAND2x1p5_ASAP7_75t_L g1489 ( 
.A(n_1306),
.B(n_1334),
.Y(n_1489)
);

HB1xp67_ASAP7_75t_L g1490 ( 
.A(n_1384),
.Y(n_1490)
);

AND2x2_ASAP7_75t_L g1491 ( 
.A(n_1272),
.B(n_1111),
.Y(n_1491)
);

INVx2_ASAP7_75t_L g1492 ( 
.A(n_1236),
.Y(n_1492)
);

OAI21xp5_ASAP7_75t_L g1493 ( 
.A1(n_1270),
.A2(n_1276),
.B(n_1275),
.Y(n_1493)
);

OR2x6_ASAP7_75t_L g1494 ( 
.A(n_1351),
.B(n_1102),
.Y(n_1494)
);

AND2x4_ASAP7_75t_L g1495 ( 
.A(n_1272),
.B(n_1203),
.Y(n_1495)
);

OAI21x1_ASAP7_75t_L g1496 ( 
.A1(n_1271),
.A2(n_1092),
.B(n_1089),
.Y(n_1496)
);

INVx4_ASAP7_75t_L g1497 ( 
.A(n_1339),
.Y(n_1497)
);

INVx1_ASAP7_75t_L g1498 ( 
.A(n_1286),
.Y(n_1498)
);

AOI22xp33_ASAP7_75t_SL g1499 ( 
.A1(n_1267),
.A2(n_1075),
.B1(n_1166),
.B2(n_1112),
.Y(n_1499)
);

AOI221xp5_ASAP7_75t_L g1500 ( 
.A1(n_1362),
.A2(n_413),
.B1(n_351),
.B2(n_416),
.C(n_352),
.Y(n_1500)
);

INVx1_ASAP7_75t_SL g1501 ( 
.A(n_1253),
.Y(n_1501)
);

AOI21xp33_ASAP7_75t_SL g1502 ( 
.A1(n_1341),
.A2(n_362),
.B(n_357),
.Y(n_1502)
);

AOI21xp33_ASAP7_75t_L g1503 ( 
.A1(n_1364),
.A2(n_1371),
.B(n_1263),
.Y(n_1503)
);

AND2x4_ASAP7_75t_L g1504 ( 
.A(n_1272),
.B(n_1313),
.Y(n_1504)
);

INVx1_ASAP7_75t_L g1505 ( 
.A(n_1367),
.Y(n_1505)
);

OAI21x1_ASAP7_75t_L g1506 ( 
.A1(n_1271),
.A2(n_1092),
.B(n_1089),
.Y(n_1506)
);

INVx1_ASAP7_75t_L g1507 ( 
.A(n_1368),
.Y(n_1507)
);

BUFx12f_ASAP7_75t_L g1508 ( 
.A(n_1287),
.Y(n_1508)
);

NAND2xp5_ASAP7_75t_L g1509 ( 
.A(n_1292),
.B(n_1116),
.Y(n_1509)
);

OA21x2_ASAP7_75t_L g1510 ( 
.A1(n_1265),
.A2(n_542),
.B(n_541),
.Y(n_1510)
);

OAI21x1_ASAP7_75t_L g1511 ( 
.A1(n_1328),
.A2(n_1092),
.B(n_1089),
.Y(n_1511)
);

INVx1_ASAP7_75t_L g1512 ( 
.A(n_1377),
.Y(n_1512)
);

INVx1_ASAP7_75t_L g1513 ( 
.A(n_1324),
.Y(n_1513)
);

OA21x2_ASAP7_75t_L g1514 ( 
.A1(n_1265),
.A2(n_1293),
.B(n_1370),
.Y(n_1514)
);

OAI21x1_ASAP7_75t_L g1515 ( 
.A1(n_1299),
.A2(n_805),
.B(n_550),
.Y(n_1515)
);

NAND3x1_ASAP7_75t_L g1516 ( 
.A(n_1310),
.B(n_466),
.C(n_1123),
.Y(n_1516)
);

AO32x2_ASAP7_75t_L g1517 ( 
.A1(n_1288),
.A2(n_1072),
.A3(n_754),
.B1(n_783),
.B2(n_1166),
.Y(n_1517)
);

AND2x4_ASAP7_75t_L g1518 ( 
.A(n_1313),
.B(n_1232),
.Y(n_1518)
);

INVx2_ASAP7_75t_L g1519 ( 
.A(n_1244),
.Y(n_1519)
);

OR2x2_ASAP7_75t_L g1520 ( 
.A(n_1302),
.B(n_1072),
.Y(n_1520)
);

BUFx3_ASAP7_75t_L g1521 ( 
.A(n_1284),
.Y(n_1521)
);

AOI22xp33_ASAP7_75t_L g1522 ( 
.A1(n_1341),
.A2(n_1262),
.B1(n_1321),
.B2(n_1305),
.Y(n_1522)
);

HB1xp67_ASAP7_75t_L g1523 ( 
.A(n_1280),
.Y(n_1523)
);

AOI21xp5_ASAP7_75t_L g1524 ( 
.A1(n_1387),
.A2(n_1232),
.B(n_1230),
.Y(n_1524)
);

OAI21xp5_ASAP7_75t_L g1525 ( 
.A1(n_1290),
.A2(n_1152),
.B(n_1116),
.Y(n_1525)
);

OAI21x1_ASAP7_75t_L g1526 ( 
.A1(n_1299),
.A2(n_550),
.B(n_543),
.Y(n_1526)
);

INVx1_ASAP7_75t_L g1527 ( 
.A(n_1248),
.Y(n_1527)
);

INVx1_ASAP7_75t_L g1528 ( 
.A(n_1318),
.Y(n_1528)
);

OAI21xp5_ASAP7_75t_L g1529 ( 
.A1(n_1295),
.A2(n_1176),
.B(n_1152),
.Y(n_1529)
);

OAI21x1_ASAP7_75t_L g1530 ( 
.A1(n_1249),
.A2(n_553),
.B(n_543),
.Y(n_1530)
);

INVxp67_ASAP7_75t_L g1531 ( 
.A(n_1239),
.Y(n_1531)
);

AND2x4_ASAP7_75t_L g1532 ( 
.A(n_1313),
.B(n_1232),
.Y(n_1532)
);

HB1xp67_ASAP7_75t_L g1533 ( 
.A(n_1304),
.Y(n_1533)
);

AOI22xp33_ASAP7_75t_L g1534 ( 
.A1(n_1319),
.A2(n_1176),
.B1(n_1166),
.B2(n_1158),
.Y(n_1534)
);

OAI21x1_ASAP7_75t_L g1535 ( 
.A1(n_1355),
.A2(n_557),
.B(n_553),
.Y(n_1535)
);

BUFx2_ASAP7_75t_SL g1536 ( 
.A(n_1256),
.Y(n_1536)
);

HB1xp67_ASAP7_75t_L g1537 ( 
.A(n_1257),
.Y(n_1537)
);

OAI21x1_ASAP7_75t_L g1538 ( 
.A1(n_1359),
.A2(n_561),
.B(n_557),
.Y(n_1538)
);

O2A1O1Ixp33_ASAP7_75t_L g1539 ( 
.A1(n_1347),
.A2(n_571),
.B(n_570),
.C(n_568),
.Y(n_1539)
);

OAI21x1_ASAP7_75t_L g1540 ( 
.A1(n_1260),
.A2(n_562),
.B(n_561),
.Y(n_1540)
);

AO21x1_ASAP7_75t_L g1541 ( 
.A1(n_1387),
.A2(n_563),
.B(n_562),
.Y(n_1541)
);

AND2x4_ASAP7_75t_L g1542 ( 
.A(n_1398),
.B(n_1363),
.Y(n_1542)
);

AOI21xp5_ASAP7_75t_L g1543 ( 
.A1(n_1301),
.A2(n_1314),
.B(n_1373),
.Y(n_1543)
);

AOI21x1_ASAP7_75t_L g1544 ( 
.A1(n_1369),
.A2(n_566),
.B(n_563),
.Y(n_1544)
);

INVx2_ASAP7_75t_L g1545 ( 
.A(n_1366),
.Y(n_1545)
);

OAI21x1_ASAP7_75t_L g1546 ( 
.A1(n_1342),
.A2(n_566),
.B(n_1166),
.Y(n_1546)
);

AOI21xp5_ASAP7_75t_L g1547 ( 
.A1(n_1356),
.A2(n_1230),
.B(n_1136),
.Y(n_1547)
);

AOI21x1_ASAP7_75t_L g1548 ( 
.A1(n_1369),
.A2(n_1166),
.B(n_1136),
.Y(n_1548)
);

INVx2_ASAP7_75t_L g1549 ( 
.A(n_1366),
.Y(n_1549)
);

OAI21x1_ASAP7_75t_L g1550 ( 
.A1(n_1397),
.A2(n_1352),
.B(n_1337),
.Y(n_1550)
);

O2A1O1Ixp33_ASAP7_75t_L g1551 ( 
.A1(n_1347),
.A2(n_318),
.B(n_374),
.C(n_371),
.Y(n_1551)
);

INVx2_ASAP7_75t_L g1552 ( 
.A(n_1366),
.Y(n_1552)
);

OAI21x1_ASAP7_75t_L g1553 ( 
.A1(n_1336),
.A2(n_1230),
.B(n_1136),
.Y(n_1553)
);

OR2x2_ASAP7_75t_L g1554 ( 
.A(n_1296),
.B(n_1230),
.Y(n_1554)
);

NAND2xp5_ASAP7_75t_L g1555 ( 
.A(n_1297),
.B(n_1105),
.Y(n_1555)
);

OAI211xp5_ASAP7_75t_L g1556 ( 
.A1(n_1362),
.A2(n_426),
.B(n_376),
.C(n_380),
.Y(n_1556)
);

NAND2xp5_ASAP7_75t_L g1557 ( 
.A(n_1325),
.B(n_1105),
.Y(n_1557)
);

BUFx3_ASAP7_75t_L g1558 ( 
.A(n_1284),
.Y(n_1558)
);

AO31x2_ASAP7_75t_L g1559 ( 
.A1(n_1329),
.A2(n_754),
.A3(n_783),
.B(n_832),
.Y(n_1559)
);

BUFx2_ASAP7_75t_L g1560 ( 
.A(n_1309),
.Y(n_1560)
);

OR2x2_ASAP7_75t_L g1561 ( 
.A(n_1327),
.B(n_1105),
.Y(n_1561)
);

AOI22xp33_ASAP7_75t_L g1562 ( 
.A1(n_1285),
.A2(n_1158),
.B1(n_851),
.B2(n_1133),
.Y(n_1562)
);

HB1xp67_ASAP7_75t_L g1563 ( 
.A(n_1361),
.Y(n_1563)
);

OAI21x1_ASAP7_75t_L g1564 ( 
.A1(n_1396),
.A2(n_1158),
.B(n_1165),
.Y(n_1564)
);

OAI21x1_ASAP7_75t_L g1565 ( 
.A1(n_1392),
.A2(n_1158),
.B(n_1165),
.Y(n_1565)
);

OAI22xp5_ASAP7_75t_L g1566 ( 
.A1(n_1358),
.A2(n_1165),
.B1(n_1133),
.B2(n_1105),
.Y(n_1566)
);

OAI21xp5_ASAP7_75t_L g1567 ( 
.A1(n_1326),
.A2(n_832),
.B(n_783),
.Y(n_1567)
);

NAND2x1p5_ASAP7_75t_L g1568 ( 
.A(n_1334),
.B(n_1133),
.Y(n_1568)
);

CKINVDCx5p33_ASAP7_75t_R g1569 ( 
.A(n_1307),
.Y(n_1569)
);

OA21x2_ASAP7_75t_L g1570 ( 
.A1(n_1380),
.A2(n_1386),
.B(n_1381),
.Y(n_1570)
);

OAI21x1_ASAP7_75t_L g1571 ( 
.A1(n_1392),
.A2(n_1393),
.B(n_1400),
.Y(n_1571)
);

INVx2_ASAP7_75t_SL g1572 ( 
.A(n_1339),
.Y(n_1572)
);

INVx1_ASAP7_75t_L g1573 ( 
.A(n_1400),
.Y(n_1573)
);

OAI21x1_ASAP7_75t_L g1574 ( 
.A1(n_1400),
.A2(n_1165),
.B(n_1133),
.Y(n_1574)
);

AND2x4_ASAP7_75t_L g1575 ( 
.A(n_1398),
.B(n_138),
.Y(n_1575)
);

OAI21xp5_ASAP7_75t_L g1576 ( 
.A1(n_1398),
.A2(n_832),
.B(n_447),
.Y(n_1576)
);

NAND2x1_ASAP7_75t_L g1577 ( 
.A(n_1334),
.B(n_728),
.Y(n_1577)
);

OAI21x1_ASAP7_75t_L g1578 ( 
.A1(n_1335),
.A2(n_1401),
.B(n_1316),
.Y(n_1578)
);

AOI21xp5_ASAP7_75t_L g1579 ( 
.A1(n_1335),
.A2(n_728),
.B(n_732),
.Y(n_1579)
);

INVx2_ASAP7_75t_L g1580 ( 
.A(n_1383),
.Y(n_1580)
);

HB1xp67_ASAP7_75t_L g1581 ( 
.A(n_1361),
.Y(n_1581)
);

OAI21x1_ASAP7_75t_L g1582 ( 
.A1(n_1401),
.A2(n_832),
.B(n_728),
.Y(n_1582)
);

OAI21x1_ASAP7_75t_L g1583 ( 
.A1(n_1401),
.A2(n_832),
.B(n_728),
.Y(n_1583)
);

BUFx2_ASAP7_75t_L g1584 ( 
.A(n_1490),
.Y(n_1584)
);

OR2x2_ASAP7_75t_L g1585 ( 
.A(n_1523),
.B(n_1277),
.Y(n_1585)
);

AOI221x1_ASAP7_75t_L g1586 ( 
.A1(n_1503),
.A2(n_1399),
.B1(n_1308),
.B2(n_1256),
.C(n_1294),
.Y(n_1586)
);

CKINVDCx6p67_ASAP7_75t_R g1587 ( 
.A(n_1508),
.Y(n_1587)
);

O2A1O1Ixp33_ASAP7_75t_L g1588 ( 
.A1(n_1404),
.A2(n_1389),
.B(n_1382),
.C(n_1395),
.Y(n_1588)
);

CKINVDCx5p33_ASAP7_75t_R g1589 ( 
.A(n_1479),
.Y(n_1589)
);

INVx6_ASAP7_75t_L g1590 ( 
.A(n_1504),
.Y(n_1590)
);

AOI22xp33_ASAP7_75t_L g1591 ( 
.A1(n_1403),
.A2(n_1363),
.B1(n_1353),
.B2(n_1357),
.Y(n_1591)
);

AOI22xp5_ASAP7_75t_L g1592 ( 
.A1(n_1428),
.A2(n_1287),
.B1(n_404),
.B2(n_405),
.Y(n_1592)
);

AOI22xp5_ASAP7_75t_L g1593 ( 
.A1(n_1405),
.A2(n_461),
.B1(n_430),
.B2(n_435),
.Y(n_1593)
);

AND2x4_ASAP7_75t_L g1594 ( 
.A(n_1504),
.B(n_1354),
.Y(n_1594)
);

AND2x2_ASAP7_75t_L g1595 ( 
.A(n_1480),
.B(n_1401),
.Y(n_1595)
);

OAI22xp5_ASAP7_75t_L g1596 ( 
.A1(n_1522),
.A2(n_1399),
.B1(n_1308),
.B2(n_1354),
.Y(n_1596)
);

INVx3_ASAP7_75t_L g1597 ( 
.A(n_1408),
.Y(n_1597)
);

INVx1_ASAP7_75t_L g1598 ( 
.A(n_1492),
.Y(n_1598)
);

AOI22xp33_ASAP7_75t_L g1599 ( 
.A1(n_1493),
.A2(n_1383),
.B1(n_311),
.B2(n_457),
.Y(n_1599)
);

INVx1_ASAP7_75t_L g1600 ( 
.A(n_1492),
.Y(n_1600)
);

NAND2xp5_ASAP7_75t_L g1601 ( 
.A(n_1431),
.B(n_1354),
.Y(n_1601)
);

NOR2xp33_ASAP7_75t_L g1602 ( 
.A(n_1501),
.B(n_1307),
.Y(n_1602)
);

A2O1A1Ixp33_ASAP7_75t_L g1603 ( 
.A1(n_1421),
.A2(n_366),
.B(n_382),
.C(n_389),
.Y(n_1603)
);

AOI211xp5_ASAP7_75t_L g1604 ( 
.A1(n_1502),
.A2(n_1412),
.B(n_1500),
.C(n_1551),
.Y(n_1604)
);

INVx1_ASAP7_75t_L g1605 ( 
.A(n_1519),
.Y(n_1605)
);

AOI22xp33_ASAP7_75t_L g1606 ( 
.A1(n_1414),
.A2(n_1450),
.B1(n_1437),
.B2(n_1434),
.Y(n_1606)
);

INVx1_ASAP7_75t_L g1607 ( 
.A(n_1519),
.Y(n_1607)
);

HB1xp67_ASAP7_75t_L g1608 ( 
.A(n_1432),
.Y(n_1608)
);

OAI22xp5_ASAP7_75t_L g1609 ( 
.A1(n_1513),
.A2(n_1294),
.B1(n_1282),
.B2(n_456),
.Y(n_1609)
);

INVxp67_ASAP7_75t_SL g1610 ( 
.A(n_1560),
.Y(n_1610)
);

INVx2_ASAP7_75t_SL g1611 ( 
.A(n_1521),
.Y(n_1611)
);

INVx3_ASAP7_75t_L g1612 ( 
.A(n_1408),
.Y(n_1612)
);

OR2x2_ASAP7_75t_L g1613 ( 
.A(n_1537),
.B(n_1282),
.Y(n_1613)
);

AOI21x1_ASAP7_75t_L g1614 ( 
.A1(n_1451),
.A2(n_1294),
.B(n_1282),
.Y(n_1614)
);

OAI22xp33_ASAP7_75t_L g1615 ( 
.A1(n_1442),
.A2(n_453),
.B1(n_395),
.B2(n_398),
.Y(n_1615)
);

INVx1_ASAP7_75t_L g1616 ( 
.A(n_1527),
.Y(n_1616)
);

NAND2xp5_ASAP7_75t_L g1617 ( 
.A(n_1513),
.B(n_390),
.Y(n_1617)
);

OAI22xp5_ASAP7_75t_L g1618 ( 
.A1(n_1407),
.A2(n_1282),
.B1(n_469),
.B2(n_463),
.Y(n_1618)
);

NOR2xp33_ASAP7_75t_L g1619 ( 
.A(n_1467),
.B(n_399),
.Y(n_1619)
);

AOI22xp33_ASAP7_75t_L g1620 ( 
.A1(n_1434),
.A2(n_311),
.B1(n_408),
.B2(n_420),
.Y(n_1620)
);

INVx3_ASAP7_75t_L g1621 ( 
.A(n_1408),
.Y(n_1621)
);

INVx2_ASAP7_75t_L g1622 ( 
.A(n_1411),
.Y(n_1622)
);

HB1xp67_ASAP7_75t_L g1623 ( 
.A(n_1533),
.Y(n_1623)
);

AND2x4_ASAP7_75t_L g1624 ( 
.A(n_1504),
.B(n_139),
.Y(n_1624)
);

NAND2xp5_ASAP7_75t_L g1625 ( 
.A(n_1498),
.B(n_423),
.Y(n_1625)
);

NAND2xp33_ASAP7_75t_R g1626 ( 
.A(n_1445),
.B(n_142),
.Y(n_1626)
);

INVx4_ASAP7_75t_SL g1627 ( 
.A(n_1445),
.Y(n_1627)
);

AND2x4_ASAP7_75t_L g1628 ( 
.A(n_1518),
.B(n_144),
.Y(n_1628)
);

INVx1_ASAP7_75t_L g1629 ( 
.A(n_1527),
.Y(n_1629)
);

OAI22xp5_ASAP7_75t_L g1630 ( 
.A1(n_1420),
.A2(n_424),
.B1(n_445),
.B2(n_449),
.Y(n_1630)
);

BUFx2_ASAP7_75t_L g1631 ( 
.A(n_1478),
.Y(n_1631)
);

INVx2_ASAP7_75t_L g1632 ( 
.A(n_1411),
.Y(n_1632)
);

INVx2_ASAP7_75t_L g1633 ( 
.A(n_1422),
.Y(n_1633)
);

OR2x2_ASAP7_75t_L g1634 ( 
.A(n_1520),
.B(n_451),
.Y(n_1634)
);

OAI22xp33_ASAP7_75t_L g1635 ( 
.A1(n_1445),
.A2(n_744),
.B1(n_752),
.B2(n_787),
.Y(n_1635)
);

NAND2xp5_ASAP7_75t_L g1636 ( 
.A(n_1498),
.B(n_832),
.Y(n_1636)
);

INVx1_ASAP7_75t_L g1637 ( 
.A(n_1528),
.Y(n_1637)
);

CKINVDCx5p33_ASAP7_75t_R g1638 ( 
.A(n_1479),
.Y(n_1638)
);

BUFx2_ASAP7_75t_L g1639 ( 
.A(n_1531),
.Y(n_1639)
);

INVx2_ASAP7_75t_L g1640 ( 
.A(n_1422),
.Y(n_1640)
);

AOI221x1_ASAP7_75t_L g1641 ( 
.A1(n_1410),
.A2(n_728),
.B1(n_732),
.B2(n_797),
.C(n_824),
.Y(n_1641)
);

INVx3_ASAP7_75t_L g1642 ( 
.A(n_1474),
.Y(n_1642)
);

AOI22xp33_ASAP7_75t_SL g1643 ( 
.A1(n_1556),
.A2(n_311),
.B1(n_15),
.B2(n_18),
.Y(n_1643)
);

CKINVDCx5p33_ASAP7_75t_R g1644 ( 
.A(n_1569),
.Y(n_1644)
);

NAND2xp5_ASAP7_75t_L g1645 ( 
.A(n_1480),
.B(n_14),
.Y(n_1645)
);

AO21x2_ASAP7_75t_L g1646 ( 
.A1(n_1419),
.A2(n_728),
.B(n_732),
.Y(n_1646)
);

AND2x2_ASAP7_75t_L g1647 ( 
.A(n_1486),
.B(n_145),
.Y(n_1647)
);

NAND2xp33_ASAP7_75t_R g1648 ( 
.A(n_1445),
.B(n_1494),
.Y(n_1648)
);

OA21x2_ASAP7_75t_L g1649 ( 
.A1(n_1449),
.A2(n_732),
.B(n_819),
.Y(n_1649)
);

INVx1_ASAP7_75t_SL g1650 ( 
.A(n_1521),
.Y(n_1650)
);

OR2x2_ASAP7_75t_L g1651 ( 
.A(n_1520),
.B(n_732),
.Y(n_1651)
);

INVx1_ASAP7_75t_SL g1652 ( 
.A(n_1558),
.Y(n_1652)
);

INVx3_ASAP7_75t_L g1653 ( 
.A(n_1474),
.Y(n_1653)
);

NAND2xp5_ASAP7_75t_L g1654 ( 
.A(n_1486),
.B(n_15),
.Y(n_1654)
);

INVx1_ASAP7_75t_L g1655 ( 
.A(n_1453),
.Y(n_1655)
);

CKINVDCx8_ASAP7_75t_R g1656 ( 
.A(n_1569),
.Y(n_1656)
);

BUFx2_ASAP7_75t_L g1657 ( 
.A(n_1542),
.Y(n_1657)
);

AOI22xp33_ASAP7_75t_SL g1658 ( 
.A1(n_1508),
.A2(n_19),
.B1(n_21),
.B2(n_22),
.Y(n_1658)
);

AND2x2_ASAP7_75t_L g1659 ( 
.A(n_1437),
.B(n_150),
.Y(n_1659)
);

INVx1_ASAP7_75t_L g1660 ( 
.A(n_1453),
.Y(n_1660)
);

OR2x6_ASAP7_75t_L g1661 ( 
.A(n_1494),
.B(n_732),
.Y(n_1661)
);

HB1xp67_ASAP7_75t_L g1662 ( 
.A(n_1560),
.Y(n_1662)
);

BUFx3_ASAP7_75t_L g1663 ( 
.A(n_1558),
.Y(n_1663)
);

AO21x1_ASAP7_75t_L g1664 ( 
.A1(n_1487),
.A2(n_19),
.B(n_21),
.Y(n_1664)
);

INVx2_ASAP7_75t_L g1665 ( 
.A(n_1426),
.Y(n_1665)
);

AOI22xp33_ASAP7_75t_L g1666 ( 
.A1(n_1443),
.A2(n_1448),
.B1(n_1415),
.B2(n_1494),
.Y(n_1666)
);

HB1xp67_ASAP7_75t_L g1667 ( 
.A(n_1491),
.Y(n_1667)
);

INVx1_ASAP7_75t_L g1668 ( 
.A(n_1456),
.Y(n_1668)
);

AND2x2_ASAP7_75t_L g1669 ( 
.A(n_1413),
.B(n_156),
.Y(n_1669)
);

OAI22xp5_ASAP7_75t_L g1670 ( 
.A1(n_1402),
.A2(n_787),
.B1(n_752),
.B2(n_744),
.Y(n_1670)
);

AND2x2_ASAP7_75t_L g1671 ( 
.A(n_1413),
.B(n_158),
.Y(n_1671)
);

INVx2_ASAP7_75t_L g1672 ( 
.A(n_1426),
.Y(n_1672)
);

AND2x2_ASAP7_75t_L g1673 ( 
.A(n_1448),
.B(n_160),
.Y(n_1673)
);

OAI221xp5_ASAP7_75t_L g1674 ( 
.A1(n_1502),
.A2(n_824),
.B1(n_819),
.B2(n_797),
.C(n_770),
.Y(n_1674)
);

BUFx2_ASAP7_75t_L g1675 ( 
.A(n_1542),
.Y(n_1675)
);

AOI221xp5_ASAP7_75t_L g1676 ( 
.A1(n_1447),
.A2(n_23),
.B1(n_26),
.B2(n_27),
.C(n_29),
.Y(n_1676)
);

HB1xp67_ASAP7_75t_L g1677 ( 
.A(n_1491),
.Y(n_1677)
);

NAND2x1p5_ASAP7_75t_L g1678 ( 
.A(n_1474),
.B(n_744),
.Y(n_1678)
);

CKINVDCx5p33_ASAP7_75t_R g1679 ( 
.A(n_1563),
.Y(n_1679)
);

BUFx2_ASAP7_75t_L g1680 ( 
.A(n_1542),
.Y(n_1680)
);

HB1xp67_ASAP7_75t_L g1681 ( 
.A(n_1495),
.Y(n_1681)
);

AOI22xp33_ASAP7_75t_L g1682 ( 
.A1(n_1494),
.A2(n_824),
.B1(n_819),
.B2(n_797),
.Y(n_1682)
);

AND2x2_ASAP7_75t_L g1683 ( 
.A(n_1455),
.B(n_172),
.Y(n_1683)
);

BUFx2_ASAP7_75t_L g1684 ( 
.A(n_1581),
.Y(n_1684)
);

AND2x2_ASAP7_75t_L g1685 ( 
.A(n_1455),
.B(n_173),
.Y(n_1685)
);

INVx4_ASAP7_75t_L g1686 ( 
.A(n_1495),
.Y(n_1686)
);

OR2x6_ASAP7_75t_L g1687 ( 
.A(n_1429),
.B(n_744),
.Y(n_1687)
);

INVx1_ASAP7_75t_L g1688 ( 
.A(n_1456),
.Y(n_1688)
);

NAND2xp5_ASAP7_75t_L g1689 ( 
.A(n_1464),
.B(n_34),
.Y(n_1689)
);

NAND2xp5_ASAP7_75t_L g1690 ( 
.A(n_1476),
.B(n_34),
.Y(n_1690)
);

AOI21xp5_ASAP7_75t_L g1691 ( 
.A1(n_1543),
.A2(n_787),
.B(n_752),
.Y(n_1691)
);

CKINVDCx5p33_ASAP7_75t_R g1692 ( 
.A(n_1435),
.Y(n_1692)
);

INVx1_ASAP7_75t_L g1693 ( 
.A(n_1458),
.Y(n_1693)
);

AND2x2_ASAP7_75t_L g1694 ( 
.A(n_1462),
.B(n_177),
.Y(n_1694)
);

INVx2_ASAP7_75t_L g1695 ( 
.A(n_1406),
.Y(n_1695)
);

INVx1_ASAP7_75t_L g1696 ( 
.A(n_1458),
.Y(n_1696)
);

NAND2xp33_ASAP7_75t_R g1697 ( 
.A(n_1495),
.B(n_181),
.Y(n_1697)
);

AOI22xp33_ASAP7_75t_L g1698 ( 
.A1(n_1518),
.A2(n_770),
.B1(n_787),
.B2(n_752),
.Y(n_1698)
);

AO31x2_ASAP7_75t_L g1699 ( 
.A1(n_1419),
.A2(n_35),
.A3(n_36),
.B(n_39),
.Y(n_1699)
);

INVx1_ASAP7_75t_L g1700 ( 
.A(n_1459),
.Y(n_1700)
);

AOI22xp33_ASAP7_75t_L g1701 ( 
.A1(n_1518),
.A2(n_770),
.B1(n_744),
.B2(n_42),
.Y(n_1701)
);

BUFx2_ASAP7_75t_L g1702 ( 
.A(n_1532),
.Y(n_1702)
);

INVx1_ASAP7_75t_L g1703 ( 
.A(n_1459),
.Y(n_1703)
);

OAI221xp5_ASAP7_75t_L g1704 ( 
.A1(n_1499),
.A2(n_39),
.B1(n_40),
.B2(n_43),
.C(n_44),
.Y(n_1704)
);

AOI22xp33_ASAP7_75t_SL g1705 ( 
.A1(n_1417),
.A2(n_45),
.B1(n_46),
.B2(n_47),
.Y(n_1705)
);

INVx4_ASAP7_75t_L g1706 ( 
.A(n_1457),
.Y(n_1706)
);

AOI22xp33_ASAP7_75t_L g1707 ( 
.A1(n_1518),
.A2(n_45),
.B1(n_46),
.B2(n_50),
.Y(n_1707)
);

AOI22xp33_ASAP7_75t_SL g1708 ( 
.A1(n_1417),
.A2(n_1575),
.B1(n_1576),
.B2(n_1557),
.Y(n_1708)
);

AND2x2_ASAP7_75t_L g1709 ( 
.A(n_1462),
.B(n_237),
.Y(n_1709)
);

AND2x2_ASAP7_75t_L g1710 ( 
.A(n_1406),
.B(n_231),
.Y(n_1710)
);

AOI22xp33_ASAP7_75t_L g1711 ( 
.A1(n_1575),
.A2(n_50),
.B1(n_51),
.B2(n_52),
.Y(n_1711)
);

NOR2xp33_ASAP7_75t_L g1712 ( 
.A(n_1532),
.B(n_230),
.Y(n_1712)
);

INVx4_ASAP7_75t_L g1713 ( 
.A(n_1457),
.Y(n_1713)
);

NAND2x1p5_ASAP7_75t_L g1714 ( 
.A(n_1483),
.B(n_1488),
.Y(n_1714)
);

AOI21xp5_ASAP7_75t_L g1715 ( 
.A1(n_1514),
.A2(n_228),
.B(n_224),
.Y(n_1715)
);

OR2x2_ASAP7_75t_L g1716 ( 
.A(n_1481),
.B(n_52),
.Y(n_1716)
);

CKINVDCx20_ASAP7_75t_R g1717 ( 
.A(n_1468),
.Y(n_1717)
);

AOI22xp33_ASAP7_75t_L g1718 ( 
.A1(n_1575),
.A2(n_57),
.B1(n_58),
.B2(n_59),
.Y(n_1718)
);

INVx1_ASAP7_75t_L g1719 ( 
.A(n_1418),
.Y(n_1719)
);

OAI21x1_ASAP7_75t_L g1720 ( 
.A1(n_1430),
.A2(n_221),
.B(n_218),
.Y(n_1720)
);

NAND2xp5_ASAP7_75t_L g1721 ( 
.A(n_1509),
.B(n_58),
.Y(n_1721)
);

CKINVDCx5p33_ASAP7_75t_R g1722 ( 
.A(n_1468),
.Y(n_1722)
);

NOR2xp33_ASAP7_75t_L g1723 ( 
.A(n_1532),
.B(n_212),
.Y(n_1723)
);

AO21x1_ASAP7_75t_L g1724 ( 
.A1(n_1547),
.A2(n_59),
.B(n_60),
.Y(n_1724)
);

INVx1_ASAP7_75t_L g1725 ( 
.A(n_1418),
.Y(n_1725)
);

AOI221xp5_ASAP7_75t_L g1726 ( 
.A1(n_1438),
.A2(n_60),
.B1(n_61),
.B2(n_62),
.C(n_63),
.Y(n_1726)
);

AND2x2_ASAP7_75t_L g1727 ( 
.A(n_1423),
.B(n_206),
.Y(n_1727)
);

AOI22xp33_ASAP7_75t_L g1728 ( 
.A1(n_1525),
.A2(n_62),
.B1(n_63),
.B2(n_64),
.Y(n_1728)
);

INVx3_ASAP7_75t_L g1729 ( 
.A(n_1483),
.Y(n_1729)
);

OAI22xp5_ASAP7_75t_L g1730 ( 
.A1(n_1534),
.A2(n_65),
.B1(n_66),
.B2(n_68),
.Y(n_1730)
);

CKINVDCx11_ASAP7_75t_R g1731 ( 
.A(n_1457),
.Y(n_1731)
);

OR2x2_ASAP7_75t_L g1732 ( 
.A(n_1460),
.B(n_65),
.Y(n_1732)
);

A2O1A1Ixp33_ASAP7_75t_L g1733 ( 
.A1(n_1529),
.A2(n_66),
.B(n_71),
.C(n_79),
.Y(n_1733)
);

BUFx2_ASAP7_75t_L g1734 ( 
.A(n_1454),
.Y(n_1734)
);

CKINVDCx6p67_ASAP7_75t_R g1735 ( 
.A(n_1536),
.Y(n_1735)
);

HB1xp67_ASAP7_75t_L g1736 ( 
.A(n_1554),
.Y(n_1736)
);

INVx8_ASAP7_75t_L g1737 ( 
.A(n_1457),
.Y(n_1737)
);

INVx3_ASAP7_75t_L g1738 ( 
.A(n_1483),
.Y(n_1738)
);

NAND2xp5_ASAP7_75t_L g1739 ( 
.A(n_1505),
.B(n_84),
.Y(n_1739)
);

INVx1_ASAP7_75t_L g1740 ( 
.A(n_1423),
.Y(n_1740)
);

INVx1_ASAP7_75t_L g1741 ( 
.A(n_1440),
.Y(n_1741)
);

AOI22xp33_ASAP7_75t_L g1742 ( 
.A1(n_1433),
.A2(n_85),
.B1(n_86),
.B2(n_87),
.Y(n_1742)
);

AOI22xp33_ASAP7_75t_L g1743 ( 
.A1(n_1425),
.A2(n_88),
.B1(n_93),
.B2(n_94),
.Y(n_1743)
);

AOI21xp33_ASAP7_75t_L g1744 ( 
.A1(n_1425),
.A2(n_96),
.B(n_97),
.Y(n_1744)
);

AND2x2_ASAP7_75t_L g1745 ( 
.A(n_1440),
.B(n_204),
.Y(n_1745)
);

INVx1_ASAP7_75t_L g1746 ( 
.A(n_1573),
.Y(n_1746)
);

A2O1A1Ixp33_ASAP7_75t_L g1747 ( 
.A1(n_1524),
.A2(n_96),
.B(n_99),
.C(n_102),
.Y(n_1747)
);

AOI22xp33_ASAP7_75t_L g1748 ( 
.A1(n_1505),
.A2(n_103),
.B1(n_104),
.B2(n_105),
.Y(n_1748)
);

INVx6_ASAP7_75t_L g1749 ( 
.A(n_1469),
.Y(n_1749)
);

INVx2_ASAP7_75t_L g1750 ( 
.A(n_1466),
.Y(n_1750)
);

OR2x6_ASAP7_75t_SL g1751 ( 
.A(n_1561),
.B(n_106),
.Y(n_1751)
);

NAND2x1_ASAP7_75t_L g1752 ( 
.A(n_1488),
.B(n_185),
.Y(n_1752)
);

HB1xp67_ASAP7_75t_L g1753 ( 
.A(n_1454),
.Y(n_1753)
);

OR2x2_ASAP7_75t_L g1754 ( 
.A(n_1555),
.B(n_107),
.Y(n_1754)
);

AND2x2_ASAP7_75t_L g1755 ( 
.A(n_1545),
.B(n_203),
.Y(n_1755)
);

AND2x2_ASAP7_75t_L g1756 ( 
.A(n_1545),
.B(n_198),
.Y(n_1756)
);

INVx1_ASAP7_75t_L g1757 ( 
.A(n_1573),
.Y(n_1757)
);

INVx4_ASAP7_75t_L g1758 ( 
.A(n_1482),
.Y(n_1758)
);

AOI22xp33_ASAP7_75t_L g1759 ( 
.A1(n_1507),
.A2(n_107),
.B1(n_108),
.B2(n_201),
.Y(n_1759)
);

OAI21xp5_ASAP7_75t_L g1760 ( 
.A1(n_1516),
.A2(n_108),
.B(n_1546),
.Y(n_1760)
);

AOI21xp5_ASAP7_75t_L g1761 ( 
.A1(n_1514),
.A2(n_1550),
.B(n_1472),
.Y(n_1761)
);

NAND2xp33_ASAP7_75t_SL g1762 ( 
.A(n_1482),
.B(n_1488),
.Y(n_1762)
);

INVx4_ASAP7_75t_L g1763 ( 
.A(n_1482),
.Y(n_1763)
);

AOI22xp33_ASAP7_75t_L g1764 ( 
.A1(n_1507),
.A2(n_1512),
.B1(n_1549),
.B2(n_1552),
.Y(n_1764)
);

NAND2xp5_ASAP7_75t_L g1765 ( 
.A(n_1512),
.B(n_1516),
.Y(n_1765)
);

AOI22xp33_ASAP7_75t_SL g1766 ( 
.A1(n_1416),
.A2(n_1536),
.B1(n_1514),
.B2(n_1489),
.Y(n_1766)
);

NAND2xp33_ASAP7_75t_R g1767 ( 
.A(n_1514),
.B(n_1570),
.Y(n_1767)
);

AOI21xp5_ASAP7_75t_L g1768 ( 
.A1(n_1550),
.A2(n_1472),
.B(n_1579),
.Y(n_1768)
);

AOI22xp33_ASAP7_75t_L g1769 ( 
.A1(n_1552),
.A2(n_1561),
.B1(n_1472),
.B2(n_1562),
.Y(n_1769)
);

AOI222xp33_ASAP7_75t_L g1770 ( 
.A1(n_1416),
.A2(n_1566),
.B1(n_1580),
.B2(n_1567),
.C1(n_1546),
.C2(n_1572),
.Y(n_1770)
);

O2A1O1Ixp33_ASAP7_75t_SL g1771 ( 
.A1(n_1577),
.A2(n_1572),
.B(n_1580),
.C(n_1416),
.Y(n_1771)
);

NAND2xp5_ASAP7_75t_L g1772 ( 
.A(n_1469),
.B(n_1497),
.Y(n_1772)
);

CKINVDCx5p33_ASAP7_75t_R g1773 ( 
.A(n_1482),
.Y(n_1773)
);

BUFx6f_ASAP7_75t_L g1774 ( 
.A(n_1482),
.Y(n_1774)
);

INVx6_ASAP7_75t_L g1775 ( 
.A(n_1469),
.Y(n_1775)
);

AOI22xp33_ASAP7_75t_SL g1776 ( 
.A1(n_1416),
.A2(n_1489),
.B1(n_1578),
.B2(n_1582),
.Y(n_1776)
);

NAND2xp5_ASAP7_75t_L g1777 ( 
.A(n_1497),
.B(n_1489),
.Y(n_1777)
);

AOI22xp33_ASAP7_75t_L g1778 ( 
.A1(n_1676),
.A2(n_1541),
.B1(n_1570),
.B2(n_1424),
.Y(n_1778)
);

CKINVDCx5p33_ASAP7_75t_R g1779 ( 
.A(n_1644),
.Y(n_1779)
);

AOI22xp5_ASAP7_75t_L g1780 ( 
.A1(n_1692),
.A2(n_1541),
.B1(n_1497),
.B2(n_1465),
.Y(n_1780)
);

AND2x4_ASAP7_75t_L g1781 ( 
.A(n_1686),
.B(n_1565),
.Y(n_1781)
);

OAI211xp5_ASAP7_75t_L g1782 ( 
.A1(n_1658),
.A2(n_1539),
.B(n_1416),
.C(n_1510),
.Y(n_1782)
);

OR2x2_ASAP7_75t_L g1783 ( 
.A(n_1736),
.B(n_1475),
.Y(n_1783)
);

OAI211xp5_ASAP7_75t_L g1784 ( 
.A1(n_1733),
.A2(n_1510),
.B(n_1530),
.C(n_1544),
.Y(n_1784)
);

INVx1_ASAP7_75t_L g1785 ( 
.A(n_1616),
.Y(n_1785)
);

AOI22xp33_ASAP7_75t_L g1786 ( 
.A1(n_1726),
.A2(n_1570),
.B1(n_1424),
.B2(n_1427),
.Y(n_1786)
);

NAND2xp5_ASAP7_75t_L g1787 ( 
.A(n_1601),
.B(n_1475),
.Y(n_1787)
);

OAI22xp5_ASAP7_75t_L g1788 ( 
.A1(n_1692),
.A2(n_1568),
.B1(n_1465),
.B2(n_1548),
.Y(n_1788)
);

OA21x2_ASAP7_75t_L g1789 ( 
.A1(n_1641),
.A2(n_1430),
.B(n_1441),
.Y(n_1789)
);

OAI22xp5_ASAP7_75t_L g1790 ( 
.A1(n_1606),
.A2(n_1568),
.B1(n_1548),
.B2(n_1570),
.Y(n_1790)
);

OAI221xp5_ASAP7_75t_L g1791 ( 
.A1(n_1604),
.A2(n_1510),
.B1(n_1424),
.B2(n_1544),
.C(n_1517),
.Y(n_1791)
);

AOI22xp33_ASAP7_75t_L g1792 ( 
.A1(n_1728),
.A2(n_1424),
.B1(n_1427),
.B2(n_1583),
.Y(n_1792)
);

OAI22xp33_ASAP7_75t_L g1793 ( 
.A1(n_1697),
.A2(n_1510),
.B1(n_1517),
.B2(n_1583),
.Y(n_1793)
);

AOI21xp33_ASAP7_75t_L g1794 ( 
.A1(n_1615),
.A2(n_1538),
.B(n_1535),
.Y(n_1794)
);

AOI22xp33_ASAP7_75t_L g1795 ( 
.A1(n_1704),
.A2(n_1582),
.B1(n_1540),
.B2(n_1409),
.Y(n_1795)
);

A2O1A1Ixp33_ASAP7_75t_L g1796 ( 
.A1(n_1603),
.A2(n_1578),
.B(n_1571),
.C(n_1553),
.Y(n_1796)
);

AND2x2_ASAP7_75t_L g1797 ( 
.A(n_1667),
.B(n_1677),
.Y(n_1797)
);

BUFx6f_ASAP7_75t_L g1798 ( 
.A(n_1731),
.Y(n_1798)
);

INVx1_ASAP7_75t_L g1799 ( 
.A(n_1629),
.Y(n_1799)
);

AOI22xp33_ASAP7_75t_SL g1800 ( 
.A1(n_1697),
.A2(n_1517),
.B1(n_1553),
.B2(n_1574),
.Y(n_1800)
);

AOI22xp33_ASAP7_75t_L g1801 ( 
.A1(n_1707),
.A2(n_1409),
.B1(n_1571),
.B2(n_1538),
.Y(n_1801)
);

INVx6_ASAP7_75t_L g1802 ( 
.A(n_1686),
.Y(n_1802)
);

BUFx10_ASAP7_75t_L g1803 ( 
.A(n_1644),
.Y(n_1803)
);

OAI221xp5_ASAP7_75t_L g1804 ( 
.A1(n_1603),
.A2(n_1517),
.B1(n_1559),
.B2(n_1530),
.C(n_1475),
.Y(n_1804)
);

HB1xp67_ASAP7_75t_L g1805 ( 
.A(n_1662),
.Y(n_1805)
);

NAND2xp5_ASAP7_75t_L g1806 ( 
.A(n_1608),
.B(n_1475),
.Y(n_1806)
);

HB1xp67_ASAP7_75t_L g1807 ( 
.A(n_1610),
.Y(n_1807)
);

AND2x2_ASAP7_75t_L g1808 ( 
.A(n_1681),
.B(n_1475),
.Y(n_1808)
);

INVxp67_ASAP7_75t_L g1809 ( 
.A(n_1623),
.Y(n_1809)
);

INVx2_ASAP7_75t_L g1810 ( 
.A(n_1600),
.Y(n_1810)
);

INVx3_ASAP7_75t_L g1811 ( 
.A(n_1749),
.Y(n_1811)
);

NAND2xp5_ASAP7_75t_L g1812 ( 
.A(n_1721),
.B(n_1565),
.Y(n_1812)
);

INVx2_ASAP7_75t_SL g1813 ( 
.A(n_1663),
.Y(n_1813)
);

AOI222xp33_ASAP7_75t_L g1814 ( 
.A1(n_1711),
.A2(n_1463),
.B1(n_1473),
.B2(n_1461),
.C1(n_1446),
.C2(n_1511),
.Y(n_1814)
);

AOI22xp33_ASAP7_75t_L g1815 ( 
.A1(n_1643),
.A2(n_1496),
.B1(n_1506),
.B2(n_1511),
.Y(n_1815)
);

OAI22xp5_ASAP7_75t_L g1816 ( 
.A1(n_1679),
.A2(n_1559),
.B1(n_1574),
.B2(n_1564),
.Y(n_1816)
);

OAI22xp33_ASAP7_75t_L g1817 ( 
.A1(n_1751),
.A2(n_1559),
.B1(n_1463),
.B2(n_1473),
.Y(n_1817)
);

AOI22xp33_ASAP7_75t_L g1818 ( 
.A1(n_1705),
.A2(n_1506),
.B1(n_1496),
.B2(n_1446),
.Y(n_1818)
);

OAI21xp33_ASAP7_75t_L g1819 ( 
.A1(n_1733),
.A2(n_1747),
.B(n_1718),
.Y(n_1819)
);

OAI21xp5_ASAP7_75t_SL g1820 ( 
.A1(n_1592),
.A2(n_1559),
.B(n_1564),
.Y(n_1820)
);

OAI22xp5_ASAP7_75t_L g1821 ( 
.A1(n_1679),
.A2(n_1559),
.B1(n_1444),
.B2(n_1485),
.Y(n_1821)
);

AND2x2_ASAP7_75t_L g1822 ( 
.A(n_1702),
.B(n_1444),
.Y(n_1822)
);

AOI31xp67_ASAP7_75t_L g1823 ( 
.A1(n_1750),
.A2(n_1515),
.A3(n_1449),
.B(n_1526),
.Y(n_1823)
);

AOI21xp5_ASAP7_75t_L g1824 ( 
.A1(n_1687),
.A2(n_1470),
.B(n_1471),
.Y(n_1824)
);

AOI221xp5_ASAP7_75t_L g1825 ( 
.A1(n_1744),
.A2(n_1461),
.B1(n_1439),
.B2(n_1436),
.C(n_1477),
.Y(n_1825)
);

AOI22xp33_ASAP7_75t_L g1826 ( 
.A1(n_1666),
.A2(n_1436),
.B1(n_1439),
.B2(n_1484),
.Y(n_1826)
);

AOI22xp33_ASAP7_75t_L g1827 ( 
.A1(n_1619),
.A2(n_1484),
.B1(n_1485),
.B2(n_1470),
.Y(n_1827)
);

INVx1_ASAP7_75t_L g1828 ( 
.A(n_1637),
.Y(n_1828)
);

AOI221xp5_ASAP7_75t_L g1829 ( 
.A1(n_1747),
.A2(n_1452),
.B1(n_1630),
.B2(n_1743),
.C(n_1748),
.Y(n_1829)
);

BUFx2_ASAP7_75t_L g1830 ( 
.A(n_1663),
.Y(n_1830)
);

OAI221xp5_ASAP7_75t_L g1831 ( 
.A1(n_1593),
.A2(n_1634),
.B1(n_1620),
.B2(n_1742),
.C(n_1617),
.Y(n_1831)
);

OAI211xp5_ASAP7_75t_L g1832 ( 
.A1(n_1759),
.A2(n_1760),
.B(n_1689),
.C(n_1701),
.Y(n_1832)
);

AND2x4_ASAP7_75t_L g1833 ( 
.A(n_1657),
.B(n_1675),
.Y(n_1833)
);

CKINVDCx5p33_ASAP7_75t_R g1834 ( 
.A(n_1656),
.Y(n_1834)
);

INVx3_ASAP7_75t_SL g1835 ( 
.A(n_1589),
.Y(n_1835)
);

AOI22xp33_ASAP7_75t_SL g1836 ( 
.A1(n_1730),
.A2(n_1751),
.B1(n_1669),
.B2(n_1671),
.Y(n_1836)
);

AOI221xp5_ASAP7_75t_L g1837 ( 
.A1(n_1664),
.A2(n_1724),
.B1(n_1625),
.B2(n_1765),
.C(n_1654),
.Y(n_1837)
);

INVx1_ASAP7_75t_L g1838 ( 
.A(n_1655),
.Y(n_1838)
);

AOI211xp5_ASAP7_75t_L g1839 ( 
.A1(n_1588),
.A2(n_1724),
.B(n_1618),
.C(n_1690),
.Y(n_1839)
);

AOI22xp33_ASAP7_75t_L g1840 ( 
.A1(n_1716),
.A2(n_1645),
.B1(n_1732),
.B2(n_1739),
.Y(n_1840)
);

AO221x2_ASAP7_75t_L g1841 ( 
.A1(n_1635),
.A2(n_1670),
.B1(n_1626),
.B2(n_1699),
.C(n_1771),
.Y(n_1841)
);

AOI22xp33_ASAP7_75t_SL g1842 ( 
.A1(n_1669),
.A2(n_1671),
.B1(n_1626),
.B2(n_1647),
.Y(n_1842)
);

OR2x6_ASAP7_75t_L g1843 ( 
.A(n_1661),
.B(n_1687),
.Y(n_1843)
);

NAND2xp5_ASAP7_75t_L g1844 ( 
.A(n_1584),
.B(n_1754),
.Y(n_1844)
);

AND2x2_ASAP7_75t_L g1845 ( 
.A(n_1680),
.B(n_1673),
.Y(n_1845)
);

OR2x6_ASAP7_75t_L g1846 ( 
.A(n_1661),
.B(n_1687),
.Y(n_1846)
);

INVxp67_ASAP7_75t_SL g1847 ( 
.A(n_1750),
.Y(n_1847)
);

AOI222xp33_ASAP7_75t_L g1848 ( 
.A1(n_1631),
.A2(n_1639),
.B1(n_1599),
.B2(n_1684),
.C1(n_1624),
.C2(n_1628),
.Y(n_1848)
);

INVx1_ASAP7_75t_L g1849 ( 
.A(n_1660),
.Y(n_1849)
);

AOI22xp33_ASAP7_75t_SL g1850 ( 
.A1(n_1647),
.A2(n_1628),
.B1(n_1624),
.B2(n_1673),
.Y(n_1850)
);

INVx2_ASAP7_75t_L g1851 ( 
.A(n_1605),
.Y(n_1851)
);

AOI222xp33_ASAP7_75t_L g1852 ( 
.A1(n_1624),
.A2(n_1628),
.B1(n_1602),
.B2(n_1627),
.C1(n_1712),
.C2(n_1723),
.Y(n_1852)
);

CKINVDCx11_ASAP7_75t_R g1853 ( 
.A(n_1656),
.Y(n_1853)
);

AOI221xp5_ASAP7_75t_L g1854 ( 
.A1(n_1771),
.A2(n_1609),
.B1(n_1715),
.B2(n_1769),
.C(n_1764),
.Y(n_1854)
);

AOI22xp33_ASAP7_75t_SL g1855 ( 
.A1(n_1661),
.A2(n_1638),
.B1(n_1589),
.B2(n_1717),
.Y(n_1855)
);

AOI22xp33_ASAP7_75t_L g1856 ( 
.A1(n_1708),
.A2(n_1659),
.B1(n_1590),
.B2(n_1585),
.Y(n_1856)
);

AND2x2_ASAP7_75t_L g1857 ( 
.A(n_1659),
.B(n_1613),
.Y(n_1857)
);

NOR2xp33_ASAP7_75t_SL g1858 ( 
.A(n_1638),
.B(n_1722),
.Y(n_1858)
);

OAI22xp33_ASAP7_75t_L g1859 ( 
.A1(n_1648),
.A2(n_1587),
.B1(n_1586),
.B2(n_1652),
.Y(n_1859)
);

AOI22xp33_ASAP7_75t_SL g1860 ( 
.A1(n_1717),
.A2(n_1674),
.B1(n_1685),
.B2(n_1709),
.Y(n_1860)
);

AOI22xp33_ASAP7_75t_L g1861 ( 
.A1(n_1590),
.A2(n_1594),
.B1(n_1694),
.B2(n_1683),
.Y(n_1861)
);

NAND3xp33_ASAP7_75t_L g1862 ( 
.A(n_1683),
.B(n_1727),
.C(n_1745),
.Y(n_1862)
);

INVx2_ASAP7_75t_L g1863 ( 
.A(n_1607),
.Y(n_1863)
);

A2O1A1Ixp33_ASAP7_75t_L g1864 ( 
.A1(n_1762),
.A2(n_1611),
.B(n_1682),
.C(n_1720),
.Y(n_1864)
);

AOI22xp5_ASAP7_75t_L g1865 ( 
.A1(n_1722),
.A2(n_1648),
.B1(n_1650),
.B2(n_1596),
.Y(n_1865)
);

OAI211xp5_ASAP7_75t_SL g1866 ( 
.A1(n_1770),
.A2(n_1651),
.B(n_1761),
.C(n_1636),
.Y(n_1866)
);

AOI221xp5_ASAP7_75t_L g1867 ( 
.A1(n_1668),
.A2(n_1696),
.B1(n_1703),
.B2(n_1688),
.C(n_1700),
.Y(n_1867)
);

OAI211xp5_ASAP7_75t_L g1868 ( 
.A1(n_1766),
.A2(n_1693),
.B(n_1727),
.C(n_1710),
.Y(n_1868)
);

HB1xp67_ASAP7_75t_L g1869 ( 
.A(n_1614),
.Y(n_1869)
);

BUFx6f_ASAP7_75t_L g1870 ( 
.A(n_1731),
.Y(n_1870)
);

NAND3xp33_ASAP7_75t_L g1871 ( 
.A(n_1710),
.B(n_1745),
.C(n_1755),
.Y(n_1871)
);

OR2x2_ASAP7_75t_L g1872 ( 
.A(n_1651),
.B(n_1695),
.Y(n_1872)
);

AOI22xp5_ASAP7_75t_L g1873 ( 
.A1(n_1611),
.A2(n_1627),
.B1(n_1752),
.B2(n_1762),
.Y(n_1873)
);

AO21x2_ASAP7_75t_L g1874 ( 
.A1(n_1646),
.A2(n_1746),
.B(n_1757),
.Y(n_1874)
);

AOI22xp5_ASAP7_75t_L g1875 ( 
.A1(n_1627),
.A2(n_1755),
.B1(n_1756),
.B2(n_1773),
.Y(n_1875)
);

OAI211xp5_ASAP7_75t_L g1876 ( 
.A1(n_1719),
.A2(n_1725),
.B(n_1740),
.C(n_1741),
.Y(n_1876)
);

BUFx2_ASAP7_75t_L g1877 ( 
.A(n_1773),
.Y(n_1877)
);

OAI22xp5_ASAP7_75t_L g1878 ( 
.A1(n_1735),
.A2(n_1698),
.B1(n_1777),
.B2(n_1772),
.Y(n_1878)
);

AOI21xp5_ASAP7_75t_L g1879 ( 
.A1(n_1649),
.A2(n_1646),
.B(n_1776),
.Y(n_1879)
);

AOI21x1_ASAP7_75t_L g1880 ( 
.A1(n_1753),
.A2(n_1734),
.B(n_1665),
.Y(n_1880)
);

OAI22xp5_ASAP7_75t_L g1881 ( 
.A1(n_1735),
.A2(n_1775),
.B1(n_1749),
.B2(n_1714),
.Y(n_1881)
);

OAI22xp5_ASAP7_75t_SL g1882 ( 
.A1(n_1749),
.A2(n_1775),
.B1(n_1763),
.B2(n_1758),
.Y(n_1882)
);

AOI221xp5_ASAP7_75t_L g1883 ( 
.A1(n_1595),
.A2(n_1672),
.B1(n_1640),
.B2(n_1633),
.C(n_1622),
.Y(n_1883)
);

AOI22xp33_ASAP7_75t_SL g1884 ( 
.A1(n_1595),
.A2(n_1646),
.B1(n_1775),
.B2(n_1737),
.Y(n_1884)
);

OAI221xp5_ASAP7_75t_L g1885 ( 
.A1(n_1597),
.A2(n_1612),
.B1(n_1621),
.B2(n_1729),
.C(n_1738),
.Y(n_1885)
);

OR2x2_ASAP7_75t_L g1886 ( 
.A(n_1632),
.B(n_1640),
.Y(n_1886)
);

AOI221xp5_ASAP7_75t_SL g1887 ( 
.A1(n_1774),
.A2(n_1642),
.B1(n_1653),
.B2(n_1738),
.C(n_1729),
.Y(n_1887)
);

AOI22xp33_ASAP7_75t_L g1888 ( 
.A1(n_1653),
.A2(n_1763),
.B1(n_1706),
.B2(n_1713),
.Y(n_1888)
);

OAI21x1_ASAP7_75t_L g1889 ( 
.A1(n_1678),
.A2(n_1767),
.B(n_1706),
.Y(n_1889)
);

AOI22xp33_ASAP7_75t_L g1890 ( 
.A1(n_1706),
.A2(n_1758),
.B1(n_1763),
.B2(n_1713),
.Y(n_1890)
);

AOI22xp5_ASAP7_75t_L g1891 ( 
.A1(n_1758),
.A2(n_1774),
.B1(n_1737),
.B2(n_1767),
.Y(n_1891)
);

OAI22xp33_ASAP7_75t_L g1892 ( 
.A1(n_1737),
.A2(n_1774),
.B1(n_1678),
.B2(n_1699),
.Y(n_1892)
);

HB1xp67_ASAP7_75t_L g1893 ( 
.A(n_1699),
.Y(n_1893)
);

AND2x4_ASAP7_75t_L g1894 ( 
.A(n_1699),
.B(n_1737),
.Y(n_1894)
);

INVx4_ASAP7_75t_L g1895 ( 
.A(n_1735),
.Y(n_1895)
);

BUFx6f_ASAP7_75t_L g1896 ( 
.A(n_1731),
.Y(n_1896)
);

OAI22xp5_ASAP7_75t_L g1897 ( 
.A1(n_1591),
.A2(n_1047),
.B1(n_1403),
.B2(n_1242),
.Y(n_1897)
);

OAI211xp5_ASAP7_75t_L g1898 ( 
.A1(n_1676),
.A2(n_1047),
.B(n_749),
.C(n_718),
.Y(n_1898)
);

OAI22xp5_ASAP7_75t_L g1899 ( 
.A1(n_1591),
.A2(n_1047),
.B1(n_1403),
.B2(n_1242),
.Y(n_1899)
);

BUFx6f_ASAP7_75t_L g1900 ( 
.A(n_1731),
.Y(n_1900)
);

AOI22xp33_ASAP7_75t_L g1901 ( 
.A1(n_1676),
.A2(n_1104),
.B1(n_1242),
.B2(n_1047),
.Y(n_1901)
);

AOI221xp5_ASAP7_75t_L g1902 ( 
.A1(n_1676),
.A2(n_1047),
.B1(n_1254),
.B2(n_911),
.C(n_1120),
.Y(n_1902)
);

AOI22xp33_ASAP7_75t_L g1903 ( 
.A1(n_1676),
.A2(n_1047),
.B1(n_1120),
.B2(n_1403),
.Y(n_1903)
);

OAI22xp33_ASAP7_75t_L g1904 ( 
.A1(n_1697),
.A2(n_1242),
.B1(n_1751),
.B2(n_1626),
.Y(n_1904)
);

NAND2xp5_ASAP7_75t_L g1905 ( 
.A(n_1601),
.B(n_1047),
.Y(n_1905)
);

OAI21x1_ASAP7_75t_L g1906 ( 
.A1(n_1691),
.A2(n_1550),
.B(n_1543),
.Y(n_1906)
);

AOI221xp5_ASAP7_75t_L g1907 ( 
.A1(n_1676),
.A2(n_1047),
.B1(n_1254),
.B2(n_911),
.C(n_1120),
.Y(n_1907)
);

AND2x2_ASAP7_75t_L g1908 ( 
.A(n_1667),
.B(n_1677),
.Y(n_1908)
);

AOI22xp5_ASAP7_75t_L g1909 ( 
.A1(n_1692),
.A2(n_1047),
.B1(n_1035),
.B2(n_1120),
.Y(n_1909)
);

OAI22xp5_ASAP7_75t_L g1910 ( 
.A1(n_1591),
.A2(n_1047),
.B1(n_1403),
.B2(n_1242),
.Y(n_1910)
);

INVx1_ASAP7_75t_L g1911 ( 
.A(n_1616),
.Y(n_1911)
);

BUFx2_ASAP7_75t_L g1912 ( 
.A(n_1679),
.Y(n_1912)
);

OAI21x1_ASAP7_75t_L g1913 ( 
.A1(n_1691),
.A2(n_1550),
.B(n_1543),
.Y(n_1913)
);

AND2x4_ASAP7_75t_L g1914 ( 
.A(n_1686),
.B(n_1657),
.Y(n_1914)
);

AOI21xp5_ASAP7_75t_L g1915 ( 
.A1(n_1768),
.A2(n_1421),
.B(n_1047),
.Y(n_1915)
);

AND2x2_ASAP7_75t_L g1916 ( 
.A(n_1667),
.B(n_1677),
.Y(n_1916)
);

OAI22xp5_ASAP7_75t_SL g1917 ( 
.A1(n_1658),
.A2(n_1047),
.B1(n_1035),
.B2(n_1403),
.Y(n_1917)
);

CKINVDCx20_ASAP7_75t_R g1918 ( 
.A(n_1717),
.Y(n_1918)
);

BUFx3_ASAP7_75t_L g1919 ( 
.A(n_1663),
.Y(n_1919)
);

AOI221xp5_ASAP7_75t_L g1920 ( 
.A1(n_1676),
.A2(n_1047),
.B1(n_1254),
.B2(n_911),
.C(n_1120),
.Y(n_1920)
);

INVx1_ASAP7_75t_SL g1921 ( 
.A(n_1584),
.Y(n_1921)
);

OAI221xp5_ASAP7_75t_L g1922 ( 
.A1(n_1604),
.A2(n_1047),
.B1(n_1403),
.B2(n_1120),
.C(n_1385),
.Y(n_1922)
);

AOI221xp5_ASAP7_75t_L g1923 ( 
.A1(n_1676),
.A2(n_1047),
.B1(n_1254),
.B2(n_911),
.C(n_1120),
.Y(n_1923)
);

AOI22xp33_ASAP7_75t_L g1924 ( 
.A1(n_1676),
.A2(n_1047),
.B1(n_1120),
.B2(n_1403),
.Y(n_1924)
);

INVx2_ASAP7_75t_L g1925 ( 
.A(n_1598),
.Y(n_1925)
);

AOI221xp5_ASAP7_75t_L g1926 ( 
.A1(n_1676),
.A2(n_1047),
.B1(n_1254),
.B2(n_911),
.C(n_1120),
.Y(n_1926)
);

AOI221xp5_ASAP7_75t_L g1927 ( 
.A1(n_1676),
.A2(n_1047),
.B1(n_1254),
.B2(n_911),
.C(n_1120),
.Y(n_1927)
);

AOI22xp33_ASAP7_75t_SL g1928 ( 
.A1(n_1704),
.A2(n_1104),
.B1(n_1047),
.B2(n_504),
.Y(n_1928)
);

OR2x2_ASAP7_75t_L g1929 ( 
.A(n_1736),
.B(n_1634),
.Y(n_1929)
);

BUFx2_ASAP7_75t_L g1930 ( 
.A(n_1679),
.Y(n_1930)
);

OAI22xp5_ASAP7_75t_SL g1931 ( 
.A1(n_1658),
.A2(n_1047),
.B1(n_1035),
.B2(n_1403),
.Y(n_1931)
);

INVx1_ASAP7_75t_L g1932 ( 
.A(n_1616),
.Y(n_1932)
);

AOI221xp5_ASAP7_75t_L g1933 ( 
.A1(n_1676),
.A2(n_1047),
.B1(n_1254),
.B2(n_911),
.C(n_1120),
.Y(n_1933)
);

OAI211xp5_ASAP7_75t_L g1934 ( 
.A1(n_1676),
.A2(n_1047),
.B(n_749),
.C(n_718),
.Y(n_1934)
);

AND2x2_ASAP7_75t_L g1935 ( 
.A(n_1667),
.B(n_1677),
.Y(n_1935)
);

AOI221xp5_ASAP7_75t_L g1936 ( 
.A1(n_1676),
.A2(n_1047),
.B1(n_1254),
.B2(n_911),
.C(n_1120),
.Y(n_1936)
);

INVx2_ASAP7_75t_L g1937 ( 
.A(n_1598),
.Y(n_1937)
);

AND2x2_ASAP7_75t_L g1938 ( 
.A(n_1667),
.B(n_1677),
.Y(n_1938)
);

AOI22xp33_ASAP7_75t_L g1939 ( 
.A1(n_1676),
.A2(n_1104),
.B1(n_1242),
.B2(n_1047),
.Y(n_1939)
);

INVx1_ASAP7_75t_SL g1940 ( 
.A(n_1584),
.Y(n_1940)
);

OAI21xp5_ASAP7_75t_L g1941 ( 
.A1(n_1603),
.A2(n_1047),
.B(n_1120),
.Y(n_1941)
);

OAI211xp5_ASAP7_75t_L g1942 ( 
.A1(n_1676),
.A2(n_1047),
.B(n_749),
.C(n_718),
.Y(n_1942)
);

NAND2xp5_ASAP7_75t_L g1943 ( 
.A(n_1601),
.B(n_1047),
.Y(n_1943)
);

OAI22xp33_ASAP7_75t_L g1944 ( 
.A1(n_1697),
.A2(n_1242),
.B1(n_1751),
.B2(n_1626),
.Y(n_1944)
);

AND2x4_ASAP7_75t_L g1945 ( 
.A(n_1686),
.B(n_1657),
.Y(n_1945)
);

NOR2xp33_ASAP7_75t_L g1946 ( 
.A(n_1909),
.B(n_1922),
.Y(n_1946)
);

NAND2xp5_ASAP7_75t_L g1947 ( 
.A(n_1807),
.B(n_1806),
.Y(n_1947)
);

AND2x2_ASAP7_75t_L g1948 ( 
.A(n_1884),
.B(n_1800),
.Y(n_1948)
);

AND2x2_ASAP7_75t_L g1949 ( 
.A(n_1884),
.B(n_1800),
.Y(n_1949)
);

OR2x2_ASAP7_75t_L g1950 ( 
.A(n_1783),
.B(n_1787),
.Y(n_1950)
);

INVx1_ASAP7_75t_L g1951 ( 
.A(n_1785),
.Y(n_1951)
);

AND2x2_ASAP7_75t_L g1952 ( 
.A(n_1808),
.B(n_1799),
.Y(n_1952)
);

INVx1_ASAP7_75t_L g1953 ( 
.A(n_1828),
.Y(n_1953)
);

INVx2_ASAP7_75t_L g1954 ( 
.A(n_1874),
.Y(n_1954)
);

INVx3_ASAP7_75t_L g1955 ( 
.A(n_1781),
.Y(n_1955)
);

INVx2_ASAP7_75t_L g1956 ( 
.A(n_1874),
.Y(n_1956)
);

OAI22xp5_ASAP7_75t_L g1957 ( 
.A1(n_1928),
.A2(n_1901),
.B1(n_1939),
.B2(n_1924),
.Y(n_1957)
);

INVx4_ASAP7_75t_SL g1958 ( 
.A(n_1843),
.Y(n_1958)
);

AOI22xp33_ASAP7_75t_L g1959 ( 
.A1(n_1928),
.A2(n_1941),
.B1(n_1819),
.B2(n_1944),
.Y(n_1959)
);

OR2x2_ASAP7_75t_L g1960 ( 
.A(n_1893),
.B(n_1807),
.Y(n_1960)
);

NAND2xp5_ASAP7_75t_L g1961 ( 
.A(n_1805),
.B(n_1905),
.Y(n_1961)
);

AND2x4_ASAP7_75t_L g1962 ( 
.A(n_1822),
.B(n_1894),
.Y(n_1962)
);

NAND2xp5_ASAP7_75t_L g1963 ( 
.A(n_1805),
.B(n_1943),
.Y(n_1963)
);

OAI22xp5_ASAP7_75t_L g1964 ( 
.A1(n_1901),
.A2(n_1939),
.B1(n_1903),
.B2(n_1944),
.Y(n_1964)
);

INVx2_ASAP7_75t_L g1965 ( 
.A(n_1838),
.Y(n_1965)
);

AND2x4_ASAP7_75t_L g1966 ( 
.A(n_1894),
.B(n_1889),
.Y(n_1966)
);

HB1xp67_ASAP7_75t_L g1967 ( 
.A(n_1869),
.Y(n_1967)
);

INVx2_ASAP7_75t_L g1968 ( 
.A(n_1849),
.Y(n_1968)
);

INVx2_ASAP7_75t_L g1969 ( 
.A(n_1911),
.Y(n_1969)
);

NOR2x1_ASAP7_75t_SL g1970 ( 
.A(n_1843),
.B(n_1846),
.Y(n_1970)
);

CKINVDCx5p33_ASAP7_75t_R g1971 ( 
.A(n_1853),
.Y(n_1971)
);

AND2x2_ASAP7_75t_L g1972 ( 
.A(n_1932),
.B(n_1857),
.Y(n_1972)
);

BUFx2_ASAP7_75t_L g1973 ( 
.A(n_1869),
.Y(n_1973)
);

INVx4_ASAP7_75t_L g1974 ( 
.A(n_1798),
.Y(n_1974)
);

NOR2xp33_ASAP7_75t_L g1975 ( 
.A(n_1921),
.B(n_1940),
.Y(n_1975)
);

OR2x2_ASAP7_75t_L g1976 ( 
.A(n_1872),
.B(n_1929),
.Y(n_1976)
);

AOI31xp33_ASAP7_75t_L g1977 ( 
.A1(n_1904),
.A2(n_1836),
.A3(n_1842),
.B(n_1839),
.Y(n_1977)
);

OR2x2_ASAP7_75t_L g1978 ( 
.A(n_1812),
.B(n_1821),
.Y(n_1978)
);

OR2x2_ASAP7_75t_L g1979 ( 
.A(n_1844),
.B(n_1809),
.Y(n_1979)
);

AOI22xp33_ASAP7_75t_L g1980 ( 
.A1(n_1904),
.A2(n_1902),
.B1(n_1936),
.B2(n_1933),
.Y(n_1980)
);

AND2x2_ASAP7_75t_L g1981 ( 
.A(n_1847),
.B(n_1879),
.Y(n_1981)
);

HB1xp67_ASAP7_75t_L g1982 ( 
.A(n_1880),
.Y(n_1982)
);

INVx1_ASAP7_75t_L g1983 ( 
.A(n_1810),
.Y(n_1983)
);

AOI221xp5_ASAP7_75t_L g1984 ( 
.A1(n_1898),
.A2(n_1942),
.B1(n_1934),
.B2(n_1920),
.C(n_1907),
.Y(n_1984)
);

INVx5_ASAP7_75t_L g1985 ( 
.A(n_1846),
.Y(n_1985)
);

INVxp67_ASAP7_75t_L g1986 ( 
.A(n_1876),
.Y(n_1986)
);

INVx2_ASAP7_75t_L g1987 ( 
.A(n_1823),
.Y(n_1987)
);

INVx1_ASAP7_75t_L g1988 ( 
.A(n_1851),
.Y(n_1988)
);

AND2x2_ASAP7_75t_L g1989 ( 
.A(n_1841),
.B(n_1789),
.Y(n_1989)
);

OR2x2_ASAP7_75t_L g1990 ( 
.A(n_1809),
.B(n_1797),
.Y(n_1990)
);

AND2x2_ASAP7_75t_L g1991 ( 
.A(n_1841),
.B(n_1789),
.Y(n_1991)
);

AND2x2_ASAP7_75t_L g1992 ( 
.A(n_1826),
.B(n_1796),
.Y(n_1992)
);

AOI22xp33_ASAP7_75t_L g1993 ( 
.A1(n_1923),
.A2(n_1927),
.B1(n_1926),
.B2(n_1917),
.Y(n_1993)
);

INVx1_ASAP7_75t_L g1994 ( 
.A(n_1863),
.Y(n_1994)
);

INVx1_ASAP7_75t_L g1995 ( 
.A(n_1925),
.Y(n_1995)
);

INVx2_ASAP7_75t_L g1996 ( 
.A(n_1937),
.Y(n_1996)
);

AND2x2_ASAP7_75t_L g1997 ( 
.A(n_1915),
.B(n_1824),
.Y(n_1997)
);

NAND2xp5_ASAP7_75t_L g1998 ( 
.A(n_1837),
.B(n_1867),
.Y(n_1998)
);

INVx2_ASAP7_75t_L g1999 ( 
.A(n_1886),
.Y(n_1999)
);

AND2x2_ASAP7_75t_L g2000 ( 
.A(n_1827),
.B(n_1818),
.Y(n_2000)
);

INVx2_ASAP7_75t_L g2001 ( 
.A(n_1906),
.Y(n_2001)
);

INVx1_ASAP7_75t_L g2002 ( 
.A(n_1817),
.Y(n_2002)
);

INVx1_ASAP7_75t_L g2003 ( 
.A(n_1817),
.Y(n_2003)
);

AND2x2_ASAP7_75t_L g2004 ( 
.A(n_1814),
.B(n_1816),
.Y(n_2004)
);

BUFx2_ASAP7_75t_L g2005 ( 
.A(n_1830),
.Y(n_2005)
);

AND2x2_ASAP7_75t_L g2006 ( 
.A(n_1790),
.B(n_1815),
.Y(n_2006)
);

BUFx3_ASAP7_75t_L g2007 ( 
.A(n_1798),
.Y(n_2007)
);

HB1xp67_ASAP7_75t_L g2008 ( 
.A(n_1887),
.Y(n_2008)
);

NOR2x1_ASAP7_75t_SL g2009 ( 
.A(n_1868),
.B(n_1881),
.Y(n_2009)
);

INVx2_ASAP7_75t_L g2010 ( 
.A(n_1913),
.Y(n_2010)
);

AND2x2_ASAP7_75t_L g2011 ( 
.A(n_1792),
.B(n_1825),
.Y(n_2011)
);

OR2x2_ASAP7_75t_L g2012 ( 
.A(n_1908),
.B(n_1916),
.Y(n_2012)
);

OR2x2_ASAP7_75t_L g2013 ( 
.A(n_1935),
.B(n_1938),
.Y(n_2013)
);

INVx2_ASAP7_75t_L g2014 ( 
.A(n_1791),
.Y(n_2014)
);

OR2x2_ASAP7_75t_L g2015 ( 
.A(n_1840),
.B(n_1804),
.Y(n_2015)
);

INVx4_ASAP7_75t_L g2016 ( 
.A(n_1798),
.Y(n_2016)
);

OAI21xp5_ASAP7_75t_L g2017 ( 
.A1(n_1897),
.A2(n_1910),
.B(n_1899),
.Y(n_2017)
);

INVx2_ASAP7_75t_L g2018 ( 
.A(n_1885),
.Y(n_2018)
);

INVx1_ASAP7_75t_L g2019 ( 
.A(n_1892),
.Y(n_2019)
);

AND2x2_ASAP7_75t_L g2020 ( 
.A(n_1842),
.B(n_1845),
.Y(n_2020)
);

INVx1_ASAP7_75t_L g2021 ( 
.A(n_1892),
.Y(n_2021)
);

INVx1_ASAP7_75t_L g2022 ( 
.A(n_1883),
.Y(n_2022)
);

NAND2xp5_ASAP7_75t_L g2023 ( 
.A(n_1840),
.B(n_1859),
.Y(n_2023)
);

CKINVDCx5p33_ASAP7_75t_R g2024 ( 
.A(n_1779),
.Y(n_2024)
);

OAI21x1_ASAP7_75t_L g2025 ( 
.A1(n_1795),
.A2(n_1801),
.B(n_1788),
.Y(n_2025)
);

INVx2_ASAP7_75t_L g2026 ( 
.A(n_1891),
.Y(n_2026)
);

INVx1_ASAP7_75t_L g2027 ( 
.A(n_1793),
.Y(n_2027)
);

INVx1_ASAP7_75t_L g2028 ( 
.A(n_1793),
.Y(n_2028)
);

AO21x2_ASAP7_75t_L g2029 ( 
.A1(n_1784),
.A2(n_1859),
.B(n_1794),
.Y(n_2029)
);

INVx1_ASAP7_75t_L g2030 ( 
.A(n_1866),
.Y(n_2030)
);

INVx1_ASAP7_75t_L g2031 ( 
.A(n_1866),
.Y(n_2031)
);

BUFx2_ASAP7_75t_L g2032 ( 
.A(n_1877),
.Y(n_2032)
);

AND2x2_ASAP7_75t_L g2033 ( 
.A(n_1801),
.B(n_1795),
.Y(n_2033)
);

OAI22xp33_ASAP7_75t_SL g2034 ( 
.A1(n_1831),
.A2(n_1865),
.B1(n_1780),
.B2(n_1858),
.Y(n_2034)
);

AND2x2_ASAP7_75t_L g2035 ( 
.A(n_1786),
.B(n_1820),
.Y(n_2035)
);

AND2x2_ASAP7_75t_L g2036 ( 
.A(n_1786),
.B(n_1850),
.Y(n_2036)
);

OR2x2_ASAP7_75t_L g2037 ( 
.A(n_1862),
.B(n_1871),
.Y(n_2037)
);

INVx1_ASAP7_75t_L g2038 ( 
.A(n_1864),
.Y(n_2038)
);

INVxp67_ASAP7_75t_SL g2039 ( 
.A(n_1888),
.Y(n_2039)
);

INVx1_ASAP7_75t_L g2040 ( 
.A(n_1873),
.Y(n_2040)
);

AND2x2_ASAP7_75t_L g2041 ( 
.A(n_1850),
.B(n_1860),
.Y(n_2041)
);

INVx1_ASAP7_75t_L g2042 ( 
.A(n_1888),
.Y(n_2042)
);

HB1xp67_ASAP7_75t_L g2043 ( 
.A(n_1833),
.Y(n_2043)
);

NAND2xp5_ASAP7_75t_L g2044 ( 
.A(n_1860),
.B(n_1878),
.Y(n_2044)
);

AND2x2_ASAP7_75t_SL g2045 ( 
.A(n_1798),
.B(n_1900),
.Y(n_2045)
);

NAND2xp5_ASAP7_75t_L g2046 ( 
.A(n_1854),
.B(n_1836),
.Y(n_2046)
);

AND2x2_ASAP7_75t_L g2047 ( 
.A(n_1856),
.B(n_1875),
.Y(n_2047)
);

AND2x2_ASAP7_75t_L g2048 ( 
.A(n_1782),
.B(n_1861),
.Y(n_2048)
);

AND2x2_ASAP7_75t_L g2049 ( 
.A(n_1813),
.B(n_1833),
.Y(n_2049)
);

INVx1_ASAP7_75t_L g2050 ( 
.A(n_1951),
.Y(n_2050)
);

AOI22xp33_ASAP7_75t_SL g2051 ( 
.A1(n_1957),
.A2(n_1964),
.B1(n_2017),
.B2(n_1946),
.Y(n_2051)
);

NOR2x1_ASAP7_75t_SL g2052 ( 
.A(n_2037),
.B(n_1900),
.Y(n_2052)
);

NOR3xp33_ASAP7_75t_L g2053 ( 
.A(n_1984),
.B(n_1832),
.C(n_1931),
.Y(n_2053)
);

INVx1_ASAP7_75t_SL g2054 ( 
.A(n_1976),
.Y(n_2054)
);

INVx1_ASAP7_75t_L g2055 ( 
.A(n_1953),
.Y(n_2055)
);

NAND2xp33_ASAP7_75t_R g2056 ( 
.A(n_1971),
.B(n_2024),
.Y(n_2056)
);

NAND2xp33_ASAP7_75t_L g2057 ( 
.A(n_1959),
.B(n_1900),
.Y(n_2057)
);

NAND3xp33_ASAP7_75t_L g2058 ( 
.A(n_1984),
.B(n_1829),
.C(n_1848),
.Y(n_2058)
);

AOI222xp33_ASAP7_75t_L g2059 ( 
.A1(n_1957),
.A2(n_1778),
.B1(n_1930),
.B2(n_1912),
.C1(n_1918),
.C2(n_1835),
.Y(n_2059)
);

AO21x2_ASAP7_75t_L g2060 ( 
.A1(n_1987),
.A2(n_1945),
.B(n_1914),
.Y(n_2060)
);

OAI31xp33_ASAP7_75t_L g2061 ( 
.A1(n_2034),
.A2(n_1919),
.A3(n_1882),
.B(n_1811),
.Y(n_2061)
);

INVx2_ASAP7_75t_L g2062 ( 
.A(n_1965),
.Y(n_2062)
);

AND2x2_ASAP7_75t_L g2063 ( 
.A(n_1948),
.B(n_1900),
.Y(n_2063)
);

INVx1_ASAP7_75t_L g2064 ( 
.A(n_1965),
.Y(n_2064)
);

AOI221xp5_ASAP7_75t_L g2065 ( 
.A1(n_1977),
.A2(n_1855),
.B1(n_1895),
.B2(n_1811),
.C(n_1834),
.Y(n_2065)
);

OAI22xp5_ASAP7_75t_L g2066 ( 
.A1(n_1993),
.A2(n_1855),
.B1(n_1835),
.B2(n_1896),
.Y(n_2066)
);

CKINVDCx5p33_ASAP7_75t_R g2067 ( 
.A(n_2032),
.Y(n_2067)
);

AND2x2_ASAP7_75t_L g2068 ( 
.A(n_1948),
.B(n_1870),
.Y(n_2068)
);

AOI22xp33_ASAP7_75t_L g2069 ( 
.A1(n_2017),
.A2(n_1852),
.B1(n_1870),
.B2(n_1896),
.Y(n_2069)
);

INVx2_ASAP7_75t_L g2070 ( 
.A(n_1965),
.Y(n_2070)
);

INVx1_ASAP7_75t_L g2071 ( 
.A(n_1968),
.Y(n_2071)
);

NOR2x1_ASAP7_75t_L g2072 ( 
.A(n_1961),
.B(n_1895),
.Y(n_2072)
);

OA21x2_ASAP7_75t_L g2073 ( 
.A1(n_1954),
.A2(n_1890),
.B(n_1802),
.Y(n_2073)
);

OR2x2_ASAP7_75t_L g2074 ( 
.A(n_2027),
.B(n_1870),
.Y(n_2074)
);

NAND2xp33_ASAP7_75t_SL g2075 ( 
.A(n_1998),
.B(n_1870),
.Y(n_2075)
);

OR2x2_ASAP7_75t_L g2076 ( 
.A(n_2027),
.B(n_1896),
.Y(n_2076)
);

INVx1_ASAP7_75t_L g2077 ( 
.A(n_1968),
.Y(n_2077)
);

AOI22xp33_ASAP7_75t_L g2078 ( 
.A1(n_1964),
.A2(n_1896),
.B1(n_1803),
.B2(n_1890),
.Y(n_2078)
);

NAND2xp5_ASAP7_75t_L g2079 ( 
.A(n_1961),
.B(n_1803),
.Y(n_2079)
);

AND2x4_ASAP7_75t_SL g2080 ( 
.A(n_1974),
.B(n_2016),
.Y(n_2080)
);

AOI22xp33_ASAP7_75t_L g2081 ( 
.A1(n_1980),
.A2(n_2034),
.B1(n_2046),
.B2(n_2015),
.Y(n_2081)
);

INVx1_ASAP7_75t_L g2082 ( 
.A(n_1969),
.Y(n_2082)
);

INVxp67_ASAP7_75t_L g2083 ( 
.A(n_1976),
.Y(n_2083)
);

AND2x4_ASAP7_75t_L g2084 ( 
.A(n_1958),
.B(n_1966),
.Y(n_2084)
);

OAI22xp33_ASAP7_75t_L g2085 ( 
.A1(n_1977),
.A2(n_2046),
.B1(n_2044),
.B2(n_1998),
.Y(n_2085)
);

NAND2xp5_ASAP7_75t_L g2086 ( 
.A(n_1963),
.B(n_1979),
.Y(n_2086)
);

OAI221xp5_ASAP7_75t_SL g2087 ( 
.A1(n_2015),
.A2(n_2023),
.B1(n_2044),
.B2(n_2030),
.C(n_2031),
.Y(n_2087)
);

INVx1_ASAP7_75t_L g2088 ( 
.A(n_1969),
.Y(n_2088)
);

INVx2_ASAP7_75t_SL g2089 ( 
.A(n_2005),
.Y(n_2089)
);

INVx4_ASAP7_75t_L g2090 ( 
.A(n_1974),
.Y(n_2090)
);

AND2x2_ASAP7_75t_L g2091 ( 
.A(n_1948),
.B(n_1949),
.Y(n_2091)
);

AND2x2_ASAP7_75t_L g2092 ( 
.A(n_1949),
.B(n_1952),
.Y(n_2092)
);

AO21x2_ASAP7_75t_L g2093 ( 
.A1(n_1954),
.A2(n_1956),
.B(n_2001),
.Y(n_2093)
);

CKINVDCx14_ASAP7_75t_R g2094 ( 
.A(n_2007),
.Y(n_2094)
);

OAI22xp5_ASAP7_75t_L g2095 ( 
.A1(n_1986),
.A2(n_2023),
.B1(n_2031),
.B2(n_2030),
.Y(n_2095)
);

INVx1_ASAP7_75t_L g2096 ( 
.A(n_1983),
.Y(n_2096)
);

AOI31xp33_ASAP7_75t_L g2097 ( 
.A1(n_2037),
.A2(n_1986),
.A3(n_2041),
.B(n_2040),
.Y(n_2097)
);

INVx1_ASAP7_75t_SL g2098 ( 
.A(n_2049),
.Y(n_2098)
);

AND2x4_ASAP7_75t_L g2099 ( 
.A(n_1958),
.B(n_1966),
.Y(n_2099)
);

OAI221xp5_ASAP7_75t_L g2100 ( 
.A1(n_2038),
.A2(n_2014),
.B1(n_2040),
.B2(n_1963),
.C(n_2018),
.Y(n_2100)
);

INVx2_ASAP7_75t_SL g2101 ( 
.A(n_2005),
.Y(n_2101)
);

INVx1_ASAP7_75t_L g2102 ( 
.A(n_1983),
.Y(n_2102)
);

OAI22xp33_ASAP7_75t_L g2103 ( 
.A1(n_2038),
.A2(n_2014),
.B1(n_2041),
.B2(n_1985),
.Y(n_2103)
);

OAI211xp5_ASAP7_75t_L g2104 ( 
.A1(n_2014),
.A2(n_2035),
.B(n_2011),
.C(n_2004),
.Y(n_2104)
);

INVx2_ASAP7_75t_L g2105 ( 
.A(n_1996),
.Y(n_2105)
);

AO21x2_ASAP7_75t_L g2106 ( 
.A1(n_1954),
.A2(n_1956),
.B(n_2010),
.Y(n_2106)
);

INVx1_ASAP7_75t_L g2107 ( 
.A(n_1988),
.Y(n_2107)
);

INVx1_ASAP7_75t_L g2108 ( 
.A(n_1988),
.Y(n_2108)
);

OAI22xp5_ASAP7_75t_L g2109 ( 
.A1(n_2041),
.A2(n_2045),
.B1(n_2032),
.B2(n_2035),
.Y(n_2109)
);

AOI22xp33_ASAP7_75t_L g2110 ( 
.A1(n_2047),
.A2(n_2035),
.B1(n_2036),
.B2(n_2048),
.Y(n_2110)
);

INVx1_ASAP7_75t_L g2111 ( 
.A(n_1994),
.Y(n_2111)
);

BUFx2_ASAP7_75t_L g2112 ( 
.A(n_1955),
.Y(n_2112)
);

NAND3xp33_ASAP7_75t_L g2113 ( 
.A(n_1997),
.B(n_2011),
.C(n_2018),
.Y(n_2113)
);

OAI211xp5_ASAP7_75t_L g2114 ( 
.A1(n_2011),
.A2(n_2004),
.B(n_1992),
.C(n_2036),
.Y(n_2114)
);

OR2x2_ASAP7_75t_L g2115 ( 
.A(n_2028),
.B(n_1950),
.Y(n_2115)
);

NOR2x1_ASAP7_75t_L g2116 ( 
.A(n_2007),
.B(n_1974),
.Y(n_2116)
);

HB1xp67_ASAP7_75t_L g2117 ( 
.A(n_2008),
.Y(n_2117)
);

INVx1_ASAP7_75t_L g2118 ( 
.A(n_1994),
.Y(n_2118)
);

AO21x1_ASAP7_75t_SL g2119 ( 
.A1(n_2019),
.A2(n_2021),
.B(n_2028),
.Y(n_2119)
);

INVx2_ASAP7_75t_L g2120 ( 
.A(n_1996),
.Y(n_2120)
);

OAI221xp5_ASAP7_75t_L g2121 ( 
.A1(n_2018),
.A2(n_1979),
.B1(n_2039),
.B2(n_1992),
.C(n_1975),
.Y(n_2121)
);

NAND2xp5_ASAP7_75t_L g2122 ( 
.A(n_1972),
.B(n_1999),
.Y(n_2122)
);

INVx1_ASAP7_75t_L g2123 ( 
.A(n_1995),
.Y(n_2123)
);

NOR4xp25_ASAP7_75t_SL g2124 ( 
.A(n_1973),
.B(n_2039),
.C(n_2019),
.D(n_2021),
.Y(n_2124)
);

OR2x2_ASAP7_75t_L g2125 ( 
.A(n_1950),
.B(n_1947),
.Y(n_2125)
);

OR2x2_ASAP7_75t_L g2126 ( 
.A(n_1947),
.B(n_2002),
.Y(n_2126)
);

BUFx3_ASAP7_75t_L g2127 ( 
.A(n_2080),
.Y(n_2127)
);

INVx1_ASAP7_75t_L g2128 ( 
.A(n_2062),
.Y(n_2128)
);

AND2x2_ASAP7_75t_L g2129 ( 
.A(n_2092),
.B(n_1949),
.Y(n_2129)
);

BUFx2_ASAP7_75t_L g2130 ( 
.A(n_2084),
.Y(n_2130)
);

INVx2_ASAP7_75t_L g2131 ( 
.A(n_2093),
.Y(n_2131)
);

INVx2_ASAP7_75t_L g2132 ( 
.A(n_2093),
.Y(n_2132)
);

AND2x4_ASAP7_75t_L g2133 ( 
.A(n_2084),
.B(n_1966),
.Y(n_2133)
);

INVx1_ASAP7_75t_L g2134 ( 
.A(n_2062),
.Y(n_2134)
);

AND2x2_ASAP7_75t_L g2135 ( 
.A(n_2092),
.B(n_1989),
.Y(n_2135)
);

AND2x4_ASAP7_75t_L g2136 ( 
.A(n_2084),
.B(n_1966),
.Y(n_2136)
);

INVx2_ASAP7_75t_L g2137 ( 
.A(n_2093),
.Y(n_2137)
);

INVxp67_ASAP7_75t_SL g2138 ( 
.A(n_2117),
.Y(n_2138)
);

INVxp67_ASAP7_75t_L g2139 ( 
.A(n_2086),
.Y(n_2139)
);

INVx1_ASAP7_75t_L g2140 ( 
.A(n_2070),
.Y(n_2140)
);

AND2x2_ASAP7_75t_L g2141 ( 
.A(n_2091),
.B(n_1989),
.Y(n_2141)
);

BUFx2_ASAP7_75t_L g2142 ( 
.A(n_2099),
.Y(n_2142)
);

NAND2xp5_ASAP7_75t_L g2143 ( 
.A(n_2125),
.B(n_1967),
.Y(n_2143)
);

INVx1_ASAP7_75t_L g2144 ( 
.A(n_2070),
.Y(n_2144)
);

OR2x2_ASAP7_75t_L g2145 ( 
.A(n_2115),
.B(n_2002),
.Y(n_2145)
);

AND2x4_ASAP7_75t_L g2146 ( 
.A(n_2099),
.B(n_1970),
.Y(n_2146)
);

HB1xp67_ASAP7_75t_L g2147 ( 
.A(n_2089),
.Y(n_2147)
);

NAND2xp33_ASAP7_75t_L g2148 ( 
.A(n_2053),
.B(n_2008),
.Y(n_2148)
);

AND2x2_ASAP7_75t_L g2149 ( 
.A(n_2091),
.B(n_1989),
.Y(n_2149)
);

OR2x2_ASAP7_75t_L g2150 ( 
.A(n_2115),
.B(n_2003),
.Y(n_2150)
);

OR2x2_ASAP7_75t_L g2151 ( 
.A(n_2125),
.B(n_2003),
.Y(n_2151)
);

BUFx2_ASAP7_75t_L g2152 ( 
.A(n_2099),
.Y(n_2152)
);

INVx3_ASAP7_75t_L g2153 ( 
.A(n_2060),
.Y(n_2153)
);

INVx1_ASAP7_75t_L g2154 ( 
.A(n_2064),
.Y(n_2154)
);

INVx2_ASAP7_75t_L g2155 ( 
.A(n_2106),
.Y(n_2155)
);

AND2x4_ASAP7_75t_L g2156 ( 
.A(n_2060),
.B(n_1970),
.Y(n_2156)
);

AND2x2_ASAP7_75t_L g2157 ( 
.A(n_2054),
.B(n_1991),
.Y(n_2157)
);

NAND2xp5_ASAP7_75t_L g2158 ( 
.A(n_2126),
.B(n_1967),
.Y(n_2158)
);

INVx1_ASAP7_75t_L g2159 ( 
.A(n_2071),
.Y(n_2159)
);

INVx5_ASAP7_75t_L g2160 ( 
.A(n_2090),
.Y(n_2160)
);

OR2x2_ASAP7_75t_L g2161 ( 
.A(n_2126),
.B(n_2083),
.Y(n_2161)
);

AND2x2_ASAP7_75t_SL g2162 ( 
.A(n_2057),
.B(n_1992),
.Y(n_2162)
);

INVx1_ASAP7_75t_L g2163 ( 
.A(n_2077),
.Y(n_2163)
);

NAND2xp5_ASAP7_75t_L g2164 ( 
.A(n_2113),
.B(n_1973),
.Y(n_2164)
);

NAND2xp5_ASAP7_75t_L g2165 ( 
.A(n_2096),
.B(n_1982),
.Y(n_2165)
);

NAND2xp5_ASAP7_75t_L g2166 ( 
.A(n_2102),
.B(n_1982),
.Y(n_2166)
);

AND2x2_ASAP7_75t_L g2167 ( 
.A(n_2063),
.B(n_1991),
.Y(n_2167)
);

AND2x2_ASAP7_75t_L g2168 ( 
.A(n_2063),
.B(n_1991),
.Y(n_2168)
);

AND2x2_ASAP7_75t_L g2169 ( 
.A(n_2068),
.B(n_2098),
.Y(n_2169)
);

AND2x2_ASAP7_75t_L g2170 ( 
.A(n_2068),
.B(n_2112),
.Y(n_2170)
);

OR2x2_ASAP7_75t_L g2171 ( 
.A(n_2122),
.B(n_1978),
.Y(n_2171)
);

AND2x2_ASAP7_75t_L g2172 ( 
.A(n_2112),
.B(n_1962),
.Y(n_2172)
);

OR2x2_ASAP7_75t_L g2173 ( 
.A(n_2089),
.B(n_1978),
.Y(n_2173)
);

NAND2xp5_ASAP7_75t_L g2174 ( 
.A(n_2107),
.B(n_1952),
.Y(n_2174)
);

INVx1_ASAP7_75t_L g2175 ( 
.A(n_2082),
.Y(n_2175)
);

INVx1_ASAP7_75t_L g2176 ( 
.A(n_2088),
.Y(n_2176)
);

AND2x2_ASAP7_75t_L g2177 ( 
.A(n_2101),
.B(n_1962),
.Y(n_2177)
);

OR2x2_ASAP7_75t_L g2178 ( 
.A(n_2101),
.B(n_1960),
.Y(n_2178)
);

NAND2xp5_ASAP7_75t_L g2179 ( 
.A(n_2108),
.B(n_1981),
.Y(n_2179)
);

OR2x2_ASAP7_75t_SL g2180 ( 
.A(n_2058),
.B(n_1990),
.Y(n_2180)
);

NAND2xp5_ASAP7_75t_SL g2181 ( 
.A(n_2051),
.B(n_2045),
.Y(n_2181)
);

INVx2_ASAP7_75t_L g2182 ( 
.A(n_2106),
.Y(n_2182)
);

INVx1_ASAP7_75t_L g2183 ( 
.A(n_2105),
.Y(n_2183)
);

INVx3_ASAP7_75t_L g2184 ( 
.A(n_2060),
.Y(n_2184)
);

AND2x4_ASAP7_75t_L g2185 ( 
.A(n_2116),
.B(n_1958),
.Y(n_2185)
);

INVx1_ASAP7_75t_L g2186 ( 
.A(n_2120),
.Y(n_2186)
);

INVx1_ASAP7_75t_L g2187 ( 
.A(n_2050),
.Y(n_2187)
);

NAND2x1_ASAP7_75t_L g2188 ( 
.A(n_2072),
.B(n_2073),
.Y(n_2188)
);

NAND2xp5_ASAP7_75t_L g2189 ( 
.A(n_2139),
.B(n_2110),
.Y(n_2189)
);

AOI221xp5_ASAP7_75t_L g2190 ( 
.A1(n_2148),
.A2(n_2085),
.B1(n_2097),
.B2(n_2095),
.C(n_2087),
.Y(n_2190)
);

OR2x2_ASAP7_75t_L g2191 ( 
.A(n_2164),
.B(n_1990),
.Y(n_2191)
);

NOR2x1p5_ASAP7_75t_L g2192 ( 
.A(n_2146),
.B(n_2007),
.Y(n_2192)
);

NAND2xp5_ASAP7_75t_L g2193 ( 
.A(n_2129),
.B(n_2164),
.Y(n_2193)
);

INVx1_ASAP7_75t_L g2194 ( 
.A(n_2187),
.Y(n_2194)
);

INVx1_ASAP7_75t_L g2195 ( 
.A(n_2187),
.Y(n_2195)
);

INVx1_ASAP7_75t_L g2196 ( 
.A(n_2154),
.Y(n_2196)
);

NAND2xp5_ASAP7_75t_SL g2197 ( 
.A(n_2162),
.B(n_2114),
.Y(n_2197)
);

INVx1_ASAP7_75t_L g2198 ( 
.A(n_2154),
.Y(n_2198)
);

AND2x2_ASAP7_75t_L g2199 ( 
.A(n_2130),
.B(n_2094),
.Y(n_2199)
);

INVx1_ASAP7_75t_L g2200 ( 
.A(n_2159),
.Y(n_2200)
);

INVx1_ASAP7_75t_L g2201 ( 
.A(n_2159),
.Y(n_2201)
);

INVx1_ASAP7_75t_L g2202 ( 
.A(n_2163),
.Y(n_2202)
);

AND2x2_ASAP7_75t_L g2203 ( 
.A(n_2130),
.B(n_2094),
.Y(n_2203)
);

AND2x2_ASAP7_75t_L g2204 ( 
.A(n_2142),
.B(n_2119),
.Y(n_2204)
);

INVx2_ASAP7_75t_L g2205 ( 
.A(n_2131),
.Y(n_2205)
);

INVx1_ASAP7_75t_L g2206 ( 
.A(n_2163),
.Y(n_2206)
);

OR2x2_ASAP7_75t_L g2207 ( 
.A(n_2151),
.B(n_2012),
.Y(n_2207)
);

HB1xp67_ASAP7_75t_L g2208 ( 
.A(n_2145),
.Y(n_2208)
);

NAND2xp5_ASAP7_75t_L g2209 ( 
.A(n_2129),
.B(n_2079),
.Y(n_2209)
);

INVx4_ASAP7_75t_L g2210 ( 
.A(n_2160),
.Y(n_2210)
);

OR2x2_ASAP7_75t_L g2211 ( 
.A(n_2151),
.B(n_2012),
.Y(n_2211)
);

OR2x2_ASAP7_75t_L g2212 ( 
.A(n_2143),
.B(n_2013),
.Y(n_2212)
);

INVx1_ASAP7_75t_L g2213 ( 
.A(n_2175),
.Y(n_2213)
);

NAND2xp5_ASAP7_75t_L g2214 ( 
.A(n_2171),
.B(n_2013),
.Y(n_2214)
);

AND2x2_ASAP7_75t_L g2215 ( 
.A(n_2142),
.B(n_2119),
.Y(n_2215)
);

INVx1_ASAP7_75t_L g2216 ( 
.A(n_2175),
.Y(n_2216)
);

OR2x2_ASAP7_75t_L g2217 ( 
.A(n_2143),
.B(n_2074),
.Y(n_2217)
);

NOR2x1_ASAP7_75t_L g2218 ( 
.A(n_2188),
.B(n_2104),
.Y(n_2218)
);

INVx1_ASAP7_75t_L g2219 ( 
.A(n_2176),
.Y(n_2219)
);

AND2x2_ASAP7_75t_L g2220 ( 
.A(n_2152),
.B(n_2135),
.Y(n_2220)
);

OR2x2_ASAP7_75t_L g2221 ( 
.A(n_2145),
.B(n_2074),
.Y(n_2221)
);

INVx1_ASAP7_75t_L g2222 ( 
.A(n_2176),
.Y(n_2222)
);

OR2x2_ASAP7_75t_L g2223 ( 
.A(n_2150),
.B(n_2076),
.Y(n_2223)
);

NAND2xp5_ASAP7_75t_L g2224 ( 
.A(n_2171),
.B(n_1972),
.Y(n_2224)
);

INVx1_ASAP7_75t_L g2225 ( 
.A(n_2165),
.Y(n_2225)
);

INVx1_ASAP7_75t_L g2226 ( 
.A(n_2165),
.Y(n_2226)
);

INVx2_ASAP7_75t_L g2227 ( 
.A(n_2131),
.Y(n_2227)
);

INVxp67_ASAP7_75t_L g2228 ( 
.A(n_2138),
.Y(n_2228)
);

OAI31xp33_ASAP7_75t_L g2229 ( 
.A1(n_2181),
.A2(n_2061),
.A3(n_2121),
.B(n_2066),
.Y(n_2229)
);

AND2x4_ASAP7_75t_L g2230 ( 
.A(n_2146),
.B(n_2052),
.Y(n_2230)
);

NAND2xp5_ASAP7_75t_L g2231 ( 
.A(n_2141),
.B(n_2111),
.Y(n_2231)
);

NAND2xp5_ASAP7_75t_L g2232 ( 
.A(n_2141),
.B(n_2118),
.Y(n_2232)
);

INVx1_ASAP7_75t_L g2233 ( 
.A(n_2166),
.Y(n_2233)
);

INVx1_ASAP7_75t_L g2234 ( 
.A(n_2166),
.Y(n_2234)
);

NOR2xp33_ASAP7_75t_L g2235 ( 
.A(n_2180),
.B(n_2100),
.Y(n_2235)
);

OAI21xp33_ASAP7_75t_L g2236 ( 
.A1(n_2162),
.A2(n_2081),
.B(n_2059),
.Y(n_2236)
);

INVx1_ASAP7_75t_L g2237 ( 
.A(n_2161),
.Y(n_2237)
);

INVx1_ASAP7_75t_L g2238 ( 
.A(n_2161),
.Y(n_2238)
);

INVx1_ASAP7_75t_L g2239 ( 
.A(n_2150),
.Y(n_2239)
);

NAND2xp5_ASAP7_75t_L g2240 ( 
.A(n_2149),
.B(n_2123),
.Y(n_2240)
);

INVx1_ASAP7_75t_L g2241 ( 
.A(n_2174),
.Y(n_2241)
);

INVx2_ASAP7_75t_L g2242 ( 
.A(n_2205),
.Y(n_2242)
);

NOR2x1_ASAP7_75t_L g2243 ( 
.A(n_2218),
.B(n_2188),
.Y(n_2243)
);

INVx1_ASAP7_75t_L g2244 ( 
.A(n_2206),
.Y(n_2244)
);

OR2x2_ASAP7_75t_L g2245 ( 
.A(n_2193),
.B(n_2179),
.Y(n_2245)
);

INVx1_ASAP7_75t_L g2246 ( 
.A(n_2206),
.Y(n_2246)
);

AOI221xp5_ASAP7_75t_L g2247 ( 
.A1(n_2235),
.A2(n_2190),
.B1(n_2236),
.B2(n_2197),
.C(n_2229),
.Y(n_2247)
);

OAI21xp33_ASAP7_75t_SL g2248 ( 
.A1(n_2235),
.A2(n_2197),
.B(n_2192),
.Y(n_2248)
);

AND2x2_ASAP7_75t_L g2249 ( 
.A(n_2230),
.B(n_2152),
.Y(n_2249)
);

INVx1_ASAP7_75t_L g2250 ( 
.A(n_2194),
.Y(n_2250)
);

NAND3xp33_ASAP7_75t_L g2251 ( 
.A(n_2189),
.B(n_2057),
.C(n_2065),
.Y(n_2251)
);

INVx1_ASAP7_75t_L g2252 ( 
.A(n_2195),
.Y(n_2252)
);

OR2x2_ASAP7_75t_L g2253 ( 
.A(n_2217),
.B(n_2179),
.Y(n_2253)
);

INVx1_ASAP7_75t_SL g2254 ( 
.A(n_2199),
.Y(n_2254)
);

NOR2xp33_ASAP7_75t_L g2255 ( 
.A(n_2209),
.B(n_2180),
.Y(n_2255)
);

NAND2xp5_ASAP7_75t_SL g2256 ( 
.A(n_2230),
.B(n_2162),
.Y(n_2256)
);

NAND2xp5_ASAP7_75t_SL g2257 ( 
.A(n_2230),
.B(n_2185),
.Y(n_2257)
);

AND2x2_ASAP7_75t_L g2258 ( 
.A(n_2204),
.B(n_2133),
.Y(n_2258)
);

AND2x2_ASAP7_75t_L g2259 ( 
.A(n_2204),
.B(n_2133),
.Y(n_2259)
);

INVx2_ASAP7_75t_L g2260 ( 
.A(n_2205),
.Y(n_2260)
);

NAND2xp5_ASAP7_75t_L g2261 ( 
.A(n_2228),
.B(n_2149),
.Y(n_2261)
);

NAND2xp5_ASAP7_75t_L g2262 ( 
.A(n_2241),
.B(n_2157),
.Y(n_2262)
);

NAND2xp5_ASAP7_75t_L g2263 ( 
.A(n_2214),
.B(n_2157),
.Y(n_2263)
);

NAND2xp5_ASAP7_75t_L g2264 ( 
.A(n_2237),
.B(n_2167),
.Y(n_2264)
);

INVxp67_ASAP7_75t_L g2265 ( 
.A(n_2191),
.Y(n_2265)
);

NAND2xp5_ASAP7_75t_L g2266 ( 
.A(n_2238),
.B(n_2167),
.Y(n_2266)
);

AOI21xp5_ASAP7_75t_L g2267 ( 
.A1(n_2226),
.A2(n_2075),
.B(n_2052),
.Y(n_2267)
);

NAND2xp5_ASAP7_75t_L g2268 ( 
.A(n_2212),
.B(n_2168),
.Y(n_2268)
);

INVx1_ASAP7_75t_L g2269 ( 
.A(n_2196),
.Y(n_2269)
);

AND2x4_ASAP7_75t_SL g2270 ( 
.A(n_2199),
.B(n_2185),
.Y(n_2270)
);

OR2x2_ASAP7_75t_L g2271 ( 
.A(n_2217),
.B(n_2158),
.Y(n_2271)
);

INVx2_ASAP7_75t_SL g2272 ( 
.A(n_2203),
.Y(n_2272)
);

INVx1_ASAP7_75t_L g2273 ( 
.A(n_2198),
.Y(n_2273)
);

AND2x2_ASAP7_75t_L g2274 ( 
.A(n_2215),
.B(n_2133),
.Y(n_2274)
);

AND2x2_ASAP7_75t_L g2275 ( 
.A(n_2215),
.B(n_2220),
.Y(n_2275)
);

AOI21xp33_ASAP7_75t_L g2276 ( 
.A1(n_2233),
.A2(n_2103),
.B(n_2109),
.Y(n_2276)
);

NAND2xp5_ASAP7_75t_L g2277 ( 
.A(n_2212),
.B(n_2168),
.Y(n_2277)
);

OR2x2_ASAP7_75t_L g2278 ( 
.A(n_2221),
.B(n_2158),
.Y(n_2278)
);

INVx1_ASAP7_75t_L g2279 ( 
.A(n_2200),
.Y(n_2279)
);

NOR3xp33_ASAP7_75t_SL g2280 ( 
.A(n_2234),
.B(n_2056),
.C(n_2075),
.Y(n_2280)
);

AND2x2_ASAP7_75t_L g2281 ( 
.A(n_2220),
.B(n_2133),
.Y(n_2281)
);

AND2x2_ASAP7_75t_L g2282 ( 
.A(n_2203),
.B(n_2136),
.Y(n_2282)
);

INVx2_ASAP7_75t_SL g2283 ( 
.A(n_2210),
.Y(n_2283)
);

AND2x2_ASAP7_75t_L g2284 ( 
.A(n_2208),
.B(n_2136),
.Y(n_2284)
);

AND2x2_ASAP7_75t_L g2285 ( 
.A(n_2239),
.B(n_2136),
.Y(n_2285)
);

INVx1_ASAP7_75t_L g2286 ( 
.A(n_2201),
.Y(n_2286)
);

AOI22xp33_ASAP7_75t_L g2287 ( 
.A1(n_2191),
.A2(n_2036),
.B1(n_2006),
.B2(n_2004),
.Y(n_2287)
);

INVx1_ASAP7_75t_L g2288 ( 
.A(n_2202),
.Y(n_2288)
);

AND2x2_ASAP7_75t_L g2289 ( 
.A(n_2221),
.B(n_2136),
.Y(n_2289)
);

AND2x2_ASAP7_75t_L g2290 ( 
.A(n_2223),
.B(n_2146),
.Y(n_2290)
);

INVx6_ASAP7_75t_L g2291 ( 
.A(n_2210),
.Y(n_2291)
);

OR2x2_ASAP7_75t_L g2292 ( 
.A(n_2223),
.B(n_2173),
.Y(n_2292)
);

A2O1A1Ixp33_ASAP7_75t_L g2293 ( 
.A1(n_2247),
.A2(n_2069),
.B(n_2078),
.C(n_2047),
.Y(n_2293)
);

AND2x2_ASAP7_75t_L g2294 ( 
.A(n_2275),
.B(n_2146),
.Y(n_2294)
);

AOI221xp5_ASAP7_75t_L g2295 ( 
.A1(n_2248),
.A2(n_2225),
.B1(n_1997),
.B2(n_2213),
.C(n_2219),
.Y(n_2295)
);

AOI22xp33_ASAP7_75t_L g2296 ( 
.A1(n_2255),
.A2(n_2006),
.B1(n_2000),
.B2(n_1997),
.Y(n_2296)
);

NOR2xp33_ASAP7_75t_L g2297 ( 
.A(n_2251),
.B(n_2224),
.Y(n_2297)
);

AOI21xp5_ASAP7_75t_L g2298 ( 
.A1(n_2243),
.A2(n_2009),
.B(n_2225),
.Y(n_2298)
);

NAND2xp5_ASAP7_75t_L g2299 ( 
.A(n_2287),
.B(n_2207),
.Y(n_2299)
);

AND2x4_ASAP7_75t_L g2300 ( 
.A(n_2270),
.B(n_2210),
.Y(n_2300)
);

AND2x2_ASAP7_75t_L g2301 ( 
.A(n_2275),
.B(n_2135),
.Y(n_2301)
);

INVxp67_ASAP7_75t_L g2302 ( 
.A(n_2272),
.Y(n_2302)
);

INVx1_ASAP7_75t_L g2303 ( 
.A(n_2244),
.Y(n_2303)
);

NAND2xp5_ASAP7_75t_L g2304 ( 
.A(n_2254),
.B(n_2207),
.Y(n_2304)
);

O2A1O1Ixp33_ASAP7_75t_L g2305 ( 
.A1(n_2280),
.A2(n_2076),
.B(n_2029),
.C(n_2048),
.Y(n_2305)
);

OAI21xp5_ASAP7_75t_L g2306 ( 
.A1(n_2267),
.A2(n_2156),
.B(n_2025),
.Y(n_2306)
);

NAND2xp5_ASAP7_75t_SL g2307 ( 
.A(n_2272),
.B(n_2045),
.Y(n_2307)
);

OAI22xp5_ASAP7_75t_L g2308 ( 
.A1(n_2270),
.A2(n_2256),
.B1(n_2257),
.B2(n_2265),
.Y(n_2308)
);

INVx1_ASAP7_75t_L g2309 ( 
.A(n_2244),
.Y(n_2309)
);

INVx1_ASAP7_75t_L g2310 ( 
.A(n_2246),
.Y(n_2310)
);

NAND2xp5_ASAP7_75t_L g2311 ( 
.A(n_2285),
.B(n_2211),
.Y(n_2311)
);

AND2x4_ASAP7_75t_L g2312 ( 
.A(n_2282),
.B(n_2156),
.Y(n_2312)
);

OR2x2_ASAP7_75t_L g2313 ( 
.A(n_2271),
.B(n_2211),
.Y(n_2313)
);

AND2x2_ASAP7_75t_L g2314 ( 
.A(n_2282),
.B(n_2170),
.Y(n_2314)
);

AND2x2_ASAP7_75t_L g2315 ( 
.A(n_2258),
.B(n_2170),
.Y(n_2315)
);

NAND2xp5_ASAP7_75t_L g2316 ( 
.A(n_2285),
.B(n_2231),
.Y(n_2316)
);

NAND2xp5_ASAP7_75t_L g2317 ( 
.A(n_2276),
.B(n_2240),
.Y(n_2317)
);

INVx1_ASAP7_75t_L g2318 ( 
.A(n_2246),
.Y(n_2318)
);

INVx1_ASAP7_75t_L g2319 ( 
.A(n_2250),
.Y(n_2319)
);

AOI21xp5_ASAP7_75t_L g2320 ( 
.A1(n_2283),
.A2(n_2009),
.B(n_2124),
.Y(n_2320)
);

AND2x2_ASAP7_75t_L g2321 ( 
.A(n_2258),
.B(n_2156),
.Y(n_2321)
);

INVxp67_ASAP7_75t_L g2322 ( 
.A(n_2283),
.Y(n_2322)
);

INVx1_ASAP7_75t_L g2323 ( 
.A(n_2250),
.Y(n_2323)
);

OAI21xp33_ASAP7_75t_SL g2324 ( 
.A1(n_2281),
.A2(n_2169),
.B(n_2232),
.Y(n_2324)
);

INVx1_ASAP7_75t_L g2325 ( 
.A(n_2252),
.Y(n_2325)
);

INVx1_ASAP7_75t_L g2326 ( 
.A(n_2252),
.Y(n_2326)
);

OAI221xp5_ASAP7_75t_L g2327 ( 
.A1(n_2291),
.A2(n_2271),
.B1(n_2261),
.B2(n_2253),
.C(n_2249),
.Y(n_2327)
);

INVx1_ASAP7_75t_L g2328 ( 
.A(n_2269),
.Y(n_2328)
);

OAI21xp5_ASAP7_75t_SL g2329 ( 
.A1(n_2249),
.A2(n_2006),
.B(n_2048),
.Y(n_2329)
);

NAND2xp5_ASAP7_75t_L g2330 ( 
.A(n_2284),
.B(n_2289),
.Y(n_2330)
);

O2A1O1Ixp33_ASAP7_75t_L g2331 ( 
.A1(n_2269),
.A2(n_2029),
.B(n_2022),
.C(n_2033),
.Y(n_2331)
);

AND2x2_ASAP7_75t_L g2332 ( 
.A(n_2259),
.B(n_2156),
.Y(n_2332)
);

INVx2_ASAP7_75t_L g2333 ( 
.A(n_2289),
.Y(n_2333)
);

INVx1_ASAP7_75t_L g2334 ( 
.A(n_2303),
.Y(n_2334)
);

NOR2xp33_ASAP7_75t_L g2335 ( 
.A(n_2297),
.B(n_2291),
.Y(n_2335)
);

AND2x2_ASAP7_75t_L g2336 ( 
.A(n_2300),
.B(n_2259),
.Y(n_2336)
);

OAI22xp5_ASAP7_75t_L g2337 ( 
.A1(n_2296),
.A2(n_2291),
.B1(n_2274),
.B2(n_2277),
.Y(n_2337)
);

AOI22xp5_ASAP7_75t_L g2338 ( 
.A1(n_2308),
.A2(n_2291),
.B1(n_2284),
.B2(n_2274),
.Y(n_2338)
);

OAI221xp5_ASAP7_75t_L g2339 ( 
.A1(n_2295),
.A2(n_2278),
.B1(n_2253),
.B2(n_2288),
.C(n_2286),
.Y(n_2339)
);

O2A1O1Ixp5_ASAP7_75t_L g2340 ( 
.A1(n_2298),
.A2(n_2286),
.B(n_2288),
.C(n_2273),
.Y(n_2340)
);

INVx1_ASAP7_75t_L g2341 ( 
.A(n_2303),
.Y(n_2341)
);

INVx1_ASAP7_75t_L g2342 ( 
.A(n_2318),
.Y(n_2342)
);

INVx2_ASAP7_75t_SL g2343 ( 
.A(n_2300),
.Y(n_2343)
);

AOI32xp33_ASAP7_75t_L g2344 ( 
.A1(n_2327),
.A2(n_2290),
.A3(n_2281),
.B1(n_2279),
.B2(n_2273),
.Y(n_2344)
);

INVx2_ASAP7_75t_SL g2345 ( 
.A(n_2300),
.Y(n_2345)
);

OAI21xp33_ASAP7_75t_SL g2346 ( 
.A1(n_2307),
.A2(n_2290),
.B(n_2268),
.Y(n_2346)
);

NOR2x1_ASAP7_75t_L g2347 ( 
.A(n_2307),
.B(n_2279),
.Y(n_2347)
);

AND2x2_ASAP7_75t_L g2348 ( 
.A(n_2314),
.B(n_2292),
.Y(n_2348)
);

OAI21xp5_ASAP7_75t_L g2349 ( 
.A1(n_2305),
.A2(n_2331),
.B(n_2293),
.Y(n_2349)
);

INVx1_ASAP7_75t_L g2350 ( 
.A(n_2318),
.Y(n_2350)
);

INVxp67_ASAP7_75t_L g2351 ( 
.A(n_2322),
.Y(n_2351)
);

AND2x4_ASAP7_75t_SL g2352 ( 
.A(n_2312),
.B(n_2185),
.Y(n_2352)
);

AND2x2_ASAP7_75t_L g2353 ( 
.A(n_2314),
.B(n_2292),
.Y(n_2353)
);

INVxp33_ASAP7_75t_L g2354 ( 
.A(n_2320),
.Y(n_2354)
);

AOI22xp5_ASAP7_75t_L g2355 ( 
.A1(n_2302),
.A2(n_2185),
.B1(n_2262),
.B2(n_2266),
.Y(n_2355)
);

INVx1_ASAP7_75t_SL g2356 ( 
.A(n_2304),
.Y(n_2356)
);

OAI21xp5_ASAP7_75t_SL g2357 ( 
.A1(n_2293),
.A2(n_2000),
.B(n_2033),
.Y(n_2357)
);

NAND4xp25_ASAP7_75t_L g2358 ( 
.A(n_2317),
.B(n_2245),
.C(n_2278),
.D(n_2264),
.Y(n_2358)
);

NAND2xp5_ASAP7_75t_L g2359 ( 
.A(n_2329),
.B(n_2245),
.Y(n_2359)
);

NOR2xp33_ASAP7_75t_L g2360 ( 
.A(n_2299),
.B(n_2263),
.Y(n_2360)
);

NAND2xp5_ASAP7_75t_L g2361 ( 
.A(n_2333),
.B(n_2301),
.Y(n_2361)
);

INVx1_ASAP7_75t_SL g2362 ( 
.A(n_2330),
.Y(n_2362)
);

INVx1_ASAP7_75t_L g2363 ( 
.A(n_2325),
.Y(n_2363)
);

INVx1_ASAP7_75t_L g2364 ( 
.A(n_2325),
.Y(n_2364)
);

INVx1_ASAP7_75t_L g2365 ( 
.A(n_2334),
.Y(n_2365)
);

INVx1_ASAP7_75t_L g2366 ( 
.A(n_2341),
.Y(n_2366)
);

INVx1_ASAP7_75t_L g2367 ( 
.A(n_2342),
.Y(n_2367)
);

NOR2x1_ASAP7_75t_L g2368 ( 
.A(n_2347),
.B(n_2319),
.Y(n_2368)
);

CKINVDCx5p33_ASAP7_75t_R g2369 ( 
.A(n_2351),
.Y(n_2369)
);

INVx2_ASAP7_75t_SL g2370 ( 
.A(n_2352),
.Y(n_2370)
);

AOI211x1_ASAP7_75t_L g2371 ( 
.A1(n_2349),
.A2(n_2306),
.B(n_2294),
.C(n_2316),
.Y(n_2371)
);

NAND2xp5_ASAP7_75t_SL g2372 ( 
.A(n_2335),
.B(n_2313),
.Y(n_2372)
);

AND2x2_ASAP7_75t_L g2373 ( 
.A(n_2336),
.B(n_2294),
.Y(n_2373)
);

CKINVDCx20_ASAP7_75t_R g2374 ( 
.A(n_2335),
.Y(n_2374)
);

AND2x2_ASAP7_75t_L g2375 ( 
.A(n_2343),
.B(n_2315),
.Y(n_2375)
);

NAND2xp5_ASAP7_75t_L g2376 ( 
.A(n_2351),
.B(n_2333),
.Y(n_2376)
);

INVxp67_ASAP7_75t_L g2377 ( 
.A(n_2345),
.Y(n_2377)
);

INVx1_ASAP7_75t_L g2378 ( 
.A(n_2350),
.Y(n_2378)
);

INVxp67_ASAP7_75t_L g2379 ( 
.A(n_2338),
.Y(n_2379)
);

INVx1_ASAP7_75t_SL g2380 ( 
.A(n_2356),
.Y(n_2380)
);

INVx1_ASAP7_75t_L g2381 ( 
.A(n_2363),
.Y(n_2381)
);

NAND2xp5_ASAP7_75t_L g2382 ( 
.A(n_2362),
.B(n_2315),
.Y(n_2382)
);

INVx1_ASAP7_75t_SL g2383 ( 
.A(n_2352),
.Y(n_2383)
);

INVx1_ASAP7_75t_L g2384 ( 
.A(n_2364),
.Y(n_2384)
);

OR2x2_ASAP7_75t_L g2385 ( 
.A(n_2358),
.B(n_2313),
.Y(n_2385)
);

INVx2_ASAP7_75t_L g2386 ( 
.A(n_2348),
.Y(n_2386)
);

INVx1_ASAP7_75t_L g2387 ( 
.A(n_2361),
.Y(n_2387)
);

INVx2_ASAP7_75t_SL g2388 ( 
.A(n_2353),
.Y(n_2388)
);

NAND2xp5_ASAP7_75t_L g2389 ( 
.A(n_2360),
.B(n_2301),
.Y(n_2389)
);

INVx1_ASAP7_75t_L g2390 ( 
.A(n_2376),
.Y(n_2390)
);

HB1xp67_ASAP7_75t_L g2391 ( 
.A(n_2368),
.Y(n_2391)
);

NAND4xp25_ASAP7_75t_L g2392 ( 
.A(n_2380),
.B(n_2344),
.C(n_2357),
.D(n_2340),
.Y(n_2392)
);

NAND2xp5_ASAP7_75t_L g2393 ( 
.A(n_2369),
.B(n_2360),
.Y(n_2393)
);

A2O1A1Ixp33_ASAP7_75t_L g2394 ( 
.A1(n_2379),
.A2(n_2340),
.B(n_2354),
.C(n_2346),
.Y(n_2394)
);

INVxp67_ASAP7_75t_SL g2395 ( 
.A(n_2374),
.Y(n_2395)
);

XOR2x2_ASAP7_75t_L g2396 ( 
.A(n_2372),
.B(n_2337),
.Y(n_2396)
);

OR2x2_ASAP7_75t_L g2397 ( 
.A(n_2385),
.B(n_2359),
.Y(n_2397)
);

NOR2xp67_ASAP7_75t_L g2398 ( 
.A(n_2388),
.B(n_2355),
.Y(n_2398)
);

NAND3xp33_ASAP7_75t_L g2399 ( 
.A(n_2369),
.B(n_2354),
.C(n_2339),
.Y(n_2399)
);

AOI21xp33_ASAP7_75t_L g2400 ( 
.A1(n_2374),
.A2(n_2328),
.B(n_2326),
.Y(n_2400)
);

AND3x2_ASAP7_75t_L g2401 ( 
.A(n_2377),
.B(n_2323),
.C(n_2309),
.Y(n_2401)
);

INVx1_ASAP7_75t_L g2402 ( 
.A(n_2386),
.Y(n_2402)
);

NAND3xp33_ASAP7_75t_SL g2403 ( 
.A(n_2383),
.B(n_2067),
.C(n_2311),
.Y(n_2403)
);

NAND3xp33_ASAP7_75t_L g2404 ( 
.A(n_2371),
.B(n_2310),
.C(n_2324),
.Y(n_2404)
);

AND4x1_ASAP7_75t_L g2405 ( 
.A(n_2399),
.B(n_2387),
.C(n_2375),
.D(n_2382),
.Y(n_2405)
);

AOI211xp5_ASAP7_75t_L g2406 ( 
.A1(n_2394),
.A2(n_2385),
.B(n_2370),
.C(n_2388),
.Y(n_2406)
);

NOR3x1_ASAP7_75t_L g2407 ( 
.A(n_2395),
.B(n_2370),
.C(n_2389),
.Y(n_2407)
);

AOI21xp33_ASAP7_75t_SL g2408 ( 
.A1(n_2391),
.A2(n_2386),
.B(n_2375),
.Y(n_2408)
);

NOR3xp33_ASAP7_75t_L g2409 ( 
.A(n_2393),
.B(n_2384),
.C(n_2381),
.Y(n_2409)
);

OAI211xp5_ASAP7_75t_SL g2410 ( 
.A1(n_2397),
.A2(n_2366),
.B(n_2367),
.C(n_2365),
.Y(n_2410)
);

AOI21xp5_ASAP7_75t_L g2411 ( 
.A1(n_2392),
.A2(n_2378),
.B(n_2365),
.Y(n_2411)
);

AOI221xp5_ASAP7_75t_L g2412 ( 
.A1(n_2400),
.A2(n_2378),
.B1(n_2373),
.B2(n_2312),
.C(n_2321),
.Y(n_2412)
);

NOR3xp33_ASAP7_75t_SL g2413 ( 
.A(n_2403),
.B(n_2067),
.C(n_2373),
.Y(n_2413)
);

AOI221xp5_ASAP7_75t_L g2414 ( 
.A1(n_2400),
.A2(n_2404),
.B1(n_2390),
.B2(n_2402),
.C(n_2396),
.Y(n_2414)
);

AOI211xp5_ASAP7_75t_L g2415 ( 
.A1(n_2398),
.A2(n_2312),
.B(n_2321),
.C(n_2332),
.Y(n_2415)
);

AO221x1_ASAP7_75t_L g2416 ( 
.A1(n_2401),
.A2(n_2184),
.B1(n_2153),
.B2(n_2242),
.C(n_2260),
.Y(n_2416)
);

OAI21xp5_ASAP7_75t_L g2417 ( 
.A1(n_2394),
.A2(n_2332),
.B(n_2260),
.Y(n_2417)
);

NAND2xp33_ASAP7_75t_R g2418 ( 
.A(n_2413),
.B(n_2169),
.Y(n_2418)
);

INVx1_ASAP7_75t_L g2419 ( 
.A(n_2407),
.Y(n_2419)
);

INVx1_ASAP7_75t_L g2420 ( 
.A(n_2408),
.Y(n_2420)
);

OAI22xp5_ASAP7_75t_L g2421 ( 
.A1(n_2406),
.A2(n_2173),
.B1(n_2127),
.B2(n_2242),
.Y(n_2421)
);

AOI221xp5_ASAP7_75t_L g2422 ( 
.A1(n_2414),
.A2(n_2227),
.B1(n_2216),
.B2(n_2222),
.C(n_2153),
.Y(n_2422)
);

AOI221xp5_ASAP7_75t_L g2423 ( 
.A1(n_2411),
.A2(n_2227),
.B1(n_2184),
.B2(n_2153),
.C(n_2022),
.Y(n_2423)
);

AO22x2_ASAP7_75t_L g2424 ( 
.A1(n_2409),
.A2(n_2417),
.B1(n_2405),
.B2(n_2410),
.Y(n_2424)
);

XNOR2xp5_ASAP7_75t_L g2425 ( 
.A(n_2424),
.B(n_2419),
.Y(n_2425)
);

OAI221xp5_ASAP7_75t_L g2426 ( 
.A1(n_2422),
.A2(n_2412),
.B1(n_2415),
.B2(n_2416),
.C(n_2016),
.Y(n_2426)
);

XNOR2x1_ASAP7_75t_L g2427 ( 
.A(n_2420),
.B(n_2020),
.Y(n_2427)
);

NOR2xp67_ASAP7_75t_SL g2428 ( 
.A(n_2418),
.B(n_1974),
.Y(n_2428)
);

AOI311xp33_ASAP7_75t_L g2429 ( 
.A1(n_2421),
.A2(n_2134),
.A3(n_2128),
.B(n_2140),
.C(n_2144),
.Y(n_2429)
);

XNOR2xp5_ASAP7_75t_L g2430 ( 
.A(n_2423),
.B(n_2049),
.Y(n_2430)
);

NOR4xp75_ASAP7_75t_SL g2431 ( 
.A(n_2421),
.B(n_2174),
.C(n_2160),
.D(n_2016),
.Y(n_2431)
);

NAND4xp75_ASAP7_75t_L g2432 ( 
.A(n_2420),
.B(n_2172),
.C(n_2177),
.D(n_2020),
.Y(n_2432)
);

AOI221xp5_ASAP7_75t_L g2433 ( 
.A1(n_2425),
.A2(n_2184),
.B1(n_2153),
.B2(n_2147),
.C(n_2131),
.Y(n_2433)
);

AOI22xp5_ASAP7_75t_L g2434 ( 
.A1(n_2428),
.A2(n_2016),
.B1(n_2127),
.B2(n_2160),
.Y(n_2434)
);

NAND3xp33_ASAP7_75t_SL g2435 ( 
.A(n_2426),
.B(n_2178),
.C(n_2090),
.Y(n_2435)
);

AND2x2_ASAP7_75t_L g2436 ( 
.A(n_2427),
.B(n_2432),
.Y(n_2436)
);

NOR3xp33_ASAP7_75t_SL g2437 ( 
.A(n_2430),
.B(n_2042),
.C(n_2055),
.Y(n_2437)
);

XOR2xp5_ASAP7_75t_L g2438 ( 
.A(n_2431),
.B(n_2043),
.Y(n_2438)
);

AOI22xp5_ASAP7_75t_L g2439 ( 
.A1(n_2429),
.A2(n_2127),
.B1(n_2160),
.B2(n_2184),
.Y(n_2439)
);

AND2x2_ASAP7_75t_L g2440 ( 
.A(n_2436),
.B(n_2437),
.Y(n_2440)
);

XOR2xp5_ASAP7_75t_L g2441 ( 
.A(n_2435),
.B(n_2429),
.Y(n_2441)
);

CKINVDCx20_ASAP7_75t_R g2442 ( 
.A(n_2438),
.Y(n_2442)
);

HB1xp67_ASAP7_75t_L g2443 ( 
.A(n_2434),
.Y(n_2443)
);

AOI22xp5_ASAP7_75t_L g2444 ( 
.A1(n_2442),
.A2(n_2433),
.B1(n_2439),
.B2(n_2160),
.Y(n_2444)
);

AOI22xp5_ASAP7_75t_L g2445 ( 
.A1(n_2440),
.A2(n_2441),
.B1(n_2443),
.B2(n_2160),
.Y(n_2445)
);

OAI21xp5_ASAP7_75t_L g2446 ( 
.A1(n_2445),
.A2(n_2444),
.B(n_2182),
.Y(n_2446)
);

INVx1_ASAP7_75t_L g2447 ( 
.A(n_2445),
.Y(n_2447)
);

HB1xp67_ASAP7_75t_L g2448 ( 
.A(n_2447),
.Y(n_2448)
);

INVx1_ASAP7_75t_L g2449 ( 
.A(n_2446),
.Y(n_2449)
);

INVxp33_ASAP7_75t_SL g2450 ( 
.A(n_2447),
.Y(n_2450)
);

OAI21xp5_ASAP7_75t_L g2451 ( 
.A1(n_2448),
.A2(n_2132),
.B(n_2137),
.Y(n_2451)
);

AOI222xp33_ASAP7_75t_SL g2452 ( 
.A1(n_2450),
.A2(n_2137),
.B1(n_2182),
.B2(n_2155),
.C1(n_2132),
.C2(n_2026),
.Y(n_2452)
);

NAND2x1p5_ASAP7_75t_L g2453 ( 
.A(n_2452),
.B(n_2449),
.Y(n_2453)
);

INVx1_ASAP7_75t_SL g2454 ( 
.A(n_2451),
.Y(n_2454)
);

OAI221xp5_ASAP7_75t_R g2455 ( 
.A1(n_2453),
.A2(n_2132),
.B1(n_2155),
.B2(n_2182),
.C(n_2137),
.Y(n_2455)
);

AOI221xp5_ASAP7_75t_L g2456 ( 
.A1(n_2455),
.A2(n_2454),
.B1(n_2155),
.B2(n_2186),
.C(n_2183),
.Y(n_2456)
);

AOI211xp5_ASAP7_75t_L g2457 ( 
.A1(n_2456),
.A2(n_2178),
.B(n_2186),
.C(n_2183),
.Y(n_2457)
);


endmodule