module fake_jpeg_20676_n_323 (n_3, n_2, n_1, n_0, n_10, n_4, n_8, n_9, n_6, n_5, n_7, n_323);

input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_323;

wire n_253;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_15;
wire n_141;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_13;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_11;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_14;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_317;
wire n_18;
wire n_145;
wire n_20;
wire n_303;
wire n_259;
wire n_90;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_12;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVx1_ASAP7_75t_L g11 ( 
.A(n_6),
.Y(n_11)
);

INVx11_ASAP7_75t_L g12 ( 
.A(n_9),
.Y(n_12)
);

CKINVDCx20_ASAP7_75t_R g13 ( 
.A(n_5),
.Y(n_13)
);

CKINVDCx20_ASAP7_75t_R g14 ( 
.A(n_5),
.Y(n_14)
);

INVx1_ASAP7_75t_L g15 ( 
.A(n_8),
.Y(n_15)
);

INVx4_ASAP7_75t_L g16 ( 
.A(n_5),
.Y(n_16)
);

BUFx6f_ASAP7_75t_L g17 ( 
.A(n_7),
.Y(n_17)
);

BUFx5_ASAP7_75t_L g18 ( 
.A(n_3),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_3),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_5),
.Y(n_20)
);

INVx2_ASAP7_75t_L g21 ( 
.A(n_9),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_8),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_7),
.Y(n_23)
);

INVx2_ASAP7_75t_L g24 ( 
.A(n_18),
.Y(n_24)
);

INVx4_ASAP7_75t_L g45 ( 
.A(n_24),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_17),
.Y(n_25)
);

INVx3_ASAP7_75t_SL g44 ( 
.A(n_25),
.Y(n_44)
);

INVx8_ASAP7_75t_L g26 ( 
.A(n_17),
.Y(n_26)
);

NOR2xp33_ASAP7_75t_L g39 ( 
.A(n_26),
.B(n_27),
.Y(n_39)
);

INVx2_ASAP7_75t_SL g27 ( 
.A(n_17),
.Y(n_27)
);

BUFx12f_ASAP7_75t_L g28 ( 
.A(n_17),
.Y(n_28)
);

BUFx3_ASAP7_75t_L g37 ( 
.A(n_28),
.Y(n_37)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_11),
.Y(n_29)
);

NOR2xp33_ASAP7_75t_L g41 ( 
.A(n_29),
.B(n_32),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_17),
.Y(n_30)
);

INVx2_ASAP7_75t_L g38 ( 
.A(n_30),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_21),
.Y(n_31)
);

INVx2_ASAP7_75t_L g46 ( 
.A(n_31),
.Y(n_46)
);

CKINVDCx14_ASAP7_75t_R g32 ( 
.A(n_22),
.Y(n_32)
);

INVx8_ASAP7_75t_L g33 ( 
.A(n_12),
.Y(n_33)
);

BUFx3_ASAP7_75t_L g40 ( 
.A(n_33),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_21),
.Y(n_34)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_34),
.Y(n_43)
);

INVx6_ASAP7_75t_L g35 ( 
.A(n_12),
.Y(n_35)
);

HB1xp67_ASAP7_75t_L g36 ( 
.A(n_35),
.Y(n_36)
);

CKINVDCx14_ASAP7_75t_R g42 ( 
.A(n_32),
.Y(n_42)
);

NAND2xp5_ASAP7_75t_L g49 ( 
.A(n_42),
.B(n_24),
.Y(n_49)
);

OAI21xp5_ASAP7_75t_SL g47 ( 
.A1(n_41),
.A2(n_29),
.B(n_19),
.Y(n_47)
);

INVxp67_ASAP7_75t_L g72 ( 
.A(n_47),
.Y(n_72)
);

INVx2_ASAP7_75t_L g48 ( 
.A(n_40),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g78 ( 
.A(n_48),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_49),
.B(n_56),
.Y(n_69)
);

OAI22xp5_ASAP7_75t_L g50 ( 
.A1(n_41),
.A2(n_26),
.B1(n_27),
.B2(n_21),
.Y(n_50)
);

AOI22xp5_ASAP7_75t_L g67 ( 
.A1(n_50),
.A2(n_51),
.B1(n_61),
.B2(n_44),
.Y(n_67)
);

OAI22xp5_ASAP7_75t_SL g51 ( 
.A1(n_46),
.A2(n_27),
.B1(n_26),
.B2(n_24),
.Y(n_51)
);

AOI22xp33_ASAP7_75t_SL g52 ( 
.A1(n_44),
.A2(n_21),
.B1(n_12),
.B2(n_16),
.Y(n_52)
);

AOI22xp33_ASAP7_75t_SL g70 ( 
.A1(n_52),
.A2(n_44),
.B1(n_35),
.B2(n_33),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_L g53 ( 
.A(n_42),
.B(n_34),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_L g68 ( 
.A(n_53),
.B(n_44),
.Y(n_68)
);

INVx2_ASAP7_75t_L g54 ( 
.A(n_40),
.Y(n_54)
);

INVx4_ASAP7_75t_L g79 ( 
.A(n_54),
.Y(n_79)
);

BUFx3_ASAP7_75t_L g55 ( 
.A(n_37),
.Y(n_55)
);

BUFx12f_ASAP7_75t_L g73 ( 
.A(n_55),
.Y(n_73)
);

INVx3_ASAP7_75t_L g56 ( 
.A(n_45),
.Y(n_56)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_40),
.Y(n_57)
);

INVx3_ASAP7_75t_L g63 ( 
.A(n_57),
.Y(n_63)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_38),
.Y(n_58)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_58),
.Y(n_74)
);

INVx2_ASAP7_75t_L g59 ( 
.A(n_37),
.Y(n_59)
);

INVx3_ASAP7_75t_L g66 ( 
.A(n_59),
.Y(n_66)
);

INVx11_ASAP7_75t_L g60 ( 
.A(n_36),
.Y(n_60)
);

INVx13_ASAP7_75t_L g65 ( 
.A(n_60),
.Y(n_65)
);

OAI22xp5_ASAP7_75t_L g61 ( 
.A1(n_46),
.A2(n_26),
.B1(n_27),
.B2(n_16),
.Y(n_61)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_39),
.Y(n_62)
);

INVx1_ASAP7_75t_SL g71 ( 
.A(n_62),
.Y(n_71)
);

AND2x2_ASAP7_75t_L g64 ( 
.A(n_62),
.B(n_39),
.Y(n_64)
);

INVx1_ASAP7_75t_SL g90 ( 
.A(n_64),
.Y(n_90)
);

AND2x2_ASAP7_75t_L g93 ( 
.A(n_67),
.B(n_77),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_L g87 ( 
.A(n_68),
.B(n_51),
.Y(n_87)
);

INVxp67_ASAP7_75t_L g86 ( 
.A(n_70),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_47),
.B(n_49),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_SL g88 ( 
.A(n_75),
.B(n_76),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_53),
.B(n_22),
.Y(n_76)
);

OR2x2_ASAP7_75t_SL g77 ( 
.A(n_50),
.B(n_18),
.Y(n_77)
);

CKINVDCx20_ASAP7_75t_R g80 ( 
.A(n_51),
.Y(n_80)
);

OR2x2_ASAP7_75t_L g96 ( 
.A(n_80),
.B(n_61),
.Y(n_96)
);

AOI21xp5_ASAP7_75t_SL g81 ( 
.A1(n_75),
.A2(n_15),
.B(n_11),
.Y(n_81)
);

OAI21xp5_ASAP7_75t_SL g127 ( 
.A1(n_81),
.A2(n_82),
.B(n_89),
.Y(n_127)
);

OA22x2_ASAP7_75t_L g82 ( 
.A1(n_77),
.A2(n_43),
.B1(n_45),
.B2(n_46),
.Y(n_82)
);

OAI22xp5_ASAP7_75t_SL g83 ( 
.A1(n_80),
.A2(n_52),
.B1(n_43),
.B2(n_38),
.Y(n_83)
);

AOI22xp5_ASAP7_75t_L g109 ( 
.A1(n_83),
.A2(n_94),
.B1(n_99),
.B2(n_74),
.Y(n_109)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_65),
.Y(n_84)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_84),
.Y(n_111)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_65),
.Y(n_85)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_85),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_L g116 ( 
.A(n_87),
.B(n_95),
.Y(n_116)
);

OA22x2_ASAP7_75t_L g89 ( 
.A1(n_71),
.A2(n_45),
.B1(n_38),
.B2(n_56),
.Y(n_89)
);

HB1xp67_ASAP7_75t_L g91 ( 
.A(n_66),
.Y(n_91)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_91),
.Y(n_126)
);

INVx3_ASAP7_75t_L g92 ( 
.A(n_73),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g112 ( 
.A(n_92),
.B(n_73),
.Y(n_112)
);

OAI22xp5_ASAP7_75t_L g94 ( 
.A1(n_67),
.A2(n_56),
.B1(n_48),
.B2(n_54),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_L g95 ( 
.A(n_76),
.B(n_68),
.Y(n_95)
);

AND2x2_ASAP7_75t_L g108 ( 
.A(n_96),
.B(n_34),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_L g97 ( 
.A(n_69),
.B(n_58),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g124 ( 
.A(n_97),
.B(n_74),
.Y(n_124)
);

BUFx8_ASAP7_75t_L g98 ( 
.A(n_73),
.Y(n_98)
);

INVxp67_ASAP7_75t_SL g129 ( 
.A(n_98),
.Y(n_129)
);

OAI22xp5_ASAP7_75t_SL g99 ( 
.A1(n_72),
.A2(n_48),
.B1(n_54),
.B2(n_57),
.Y(n_99)
);

MAJIxp5_ASAP7_75t_L g100 ( 
.A(n_64),
.B(n_34),
.C(n_31),
.Y(n_100)
);

MAJIxp5_ASAP7_75t_L g114 ( 
.A(n_100),
.B(n_25),
.C(n_30),
.Y(n_114)
);

INVx1_ASAP7_75t_SL g101 ( 
.A(n_89),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_L g134 ( 
.A(n_101),
.B(n_103),
.Y(n_134)
);

AOI22xp33_ASAP7_75t_L g102 ( 
.A1(n_96),
.A2(n_71),
.B1(n_69),
.B2(n_64),
.Y(n_102)
);

OAI22xp33_ASAP7_75t_SL g157 ( 
.A1(n_102),
.A2(n_16),
.B1(n_58),
.B2(n_33),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_SL g103 ( 
.A(n_95),
.B(n_31),
.Y(n_103)
);

OAI21xp5_ASAP7_75t_L g104 ( 
.A1(n_93),
.A2(n_22),
.B(n_11),
.Y(n_104)
);

OAI21xp5_ASAP7_75t_L g145 ( 
.A1(n_104),
.A2(n_115),
.B(n_11),
.Y(n_145)
);

INVxp67_ASAP7_75t_L g105 ( 
.A(n_99),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_L g137 ( 
.A(n_105),
.B(n_106),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_SL g106 ( 
.A(n_88),
.B(n_97),
.Y(n_106)
);

CKINVDCx20_ASAP7_75t_R g107 ( 
.A(n_84),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_L g130 ( 
.A(n_107),
.B(n_110),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_L g155 ( 
.A(n_108),
.B(n_113),
.Y(n_155)
);

OAI22xp5_ASAP7_75t_L g143 ( 
.A1(n_109),
.A2(n_123),
.B1(n_59),
.B2(n_60),
.Y(n_143)
);

CKINVDCx20_ASAP7_75t_R g110 ( 
.A(n_85),
.Y(n_110)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_112),
.Y(n_139)
);

CKINVDCx14_ASAP7_75t_R g113 ( 
.A(n_81),
.Y(n_113)
);

XNOR2xp5_ASAP7_75t_L g148 ( 
.A(n_114),
.B(n_30),
.Y(n_148)
);

XNOR2x1_ASAP7_75t_SL g115 ( 
.A(n_93),
.B(n_65),
.Y(n_115)
);

OAI22xp33_ASAP7_75t_SL g117 ( 
.A1(n_86),
.A2(n_96),
.B1(n_90),
.B2(n_83),
.Y(n_117)
);

AOI22xp5_ASAP7_75t_L g144 ( 
.A1(n_117),
.A2(n_60),
.B1(n_16),
.B2(n_35),
.Y(n_144)
);

CKINVDCx20_ASAP7_75t_R g118 ( 
.A(n_89),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_L g138 ( 
.A(n_118),
.B(n_128),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_L g119 ( 
.A(n_88),
.B(n_66),
.Y(n_119)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_119),
.Y(n_156)
);

INVxp67_ASAP7_75t_L g120 ( 
.A(n_82),
.Y(n_120)
);

INVxp67_ASAP7_75t_L g154 ( 
.A(n_120),
.Y(n_154)
);

OR2x2_ASAP7_75t_L g121 ( 
.A(n_90),
.B(n_79),
.Y(n_121)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_121),
.Y(n_141)
);

AOI22xp33_ASAP7_75t_SL g123 ( 
.A1(n_86),
.A2(n_79),
.B1(n_57),
.B2(n_59),
.Y(n_123)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_124),
.Y(n_164)
);

NOR2xp33_ASAP7_75t_L g125 ( 
.A(n_89),
.B(n_63),
.Y(n_125)
);

CKINVDCx16_ASAP7_75t_R g162 ( 
.A(n_125),
.Y(n_162)
);

INVxp67_ASAP7_75t_L g128 ( 
.A(n_82),
.Y(n_128)
);

AOI21xp5_ASAP7_75t_L g131 ( 
.A1(n_115),
.A2(n_93),
.B(n_94),
.Y(n_131)
);

OAI21xp5_ASAP7_75t_SL g180 ( 
.A1(n_131),
.A2(n_136),
.B(n_147),
.Y(n_180)
);

CKINVDCx20_ASAP7_75t_R g132 ( 
.A(n_112),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_SL g170 ( 
.A(n_132),
.B(n_150),
.Y(n_170)
);

AOI22xp5_ASAP7_75t_SL g133 ( 
.A1(n_115),
.A2(n_100),
.B1(n_82),
.B2(n_92),
.Y(n_133)
);

OAI21xp5_ASAP7_75t_L g166 ( 
.A1(n_133),
.A2(n_163),
.B(n_165),
.Y(n_166)
);

MAJIxp5_ASAP7_75t_L g135 ( 
.A(n_116),
.B(n_87),
.C(n_63),
.Y(n_135)
);

XOR2xp5_ASAP7_75t_L g191 ( 
.A(n_135),
.B(n_140),
.Y(n_191)
);

AOI21xp5_ASAP7_75t_SL g136 ( 
.A1(n_127),
.A2(n_23),
.B(n_15),
.Y(n_136)
);

MAJIxp5_ASAP7_75t_L g140 ( 
.A(n_116),
.B(n_79),
.C(n_78),
.Y(n_140)
);

XOR2xp5_ASAP7_75t_L g142 ( 
.A(n_106),
.B(n_36),
.Y(n_142)
);

XOR2xp5_ASAP7_75t_L g195 ( 
.A(n_142),
.B(n_148),
.Y(n_195)
);

AOI22xp5_ASAP7_75t_L g179 ( 
.A1(n_143),
.A2(n_157),
.B1(n_160),
.B2(n_107),
.Y(n_179)
);

OAI22xp5_ASAP7_75t_L g175 ( 
.A1(n_144),
.A2(n_146),
.B1(n_161),
.B2(n_125),
.Y(n_175)
);

AO21x1_ASAP7_75t_L g187 ( 
.A1(n_145),
.A2(n_111),
.B(n_18),
.Y(n_187)
);

AOI22xp5_ASAP7_75t_L g146 ( 
.A1(n_117),
.A2(n_16),
.B1(n_35),
.B2(n_33),
.Y(n_146)
);

AOI21xp5_ASAP7_75t_L g147 ( 
.A1(n_127),
.A2(n_98),
.B(n_73),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_L g149 ( 
.A(n_119),
.B(n_78),
.Y(n_149)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_149),
.Y(n_185)
);

NOR2xp33_ASAP7_75t_L g150 ( 
.A(n_102),
.B(n_78),
.Y(n_150)
);

MAJIxp5_ASAP7_75t_L g151 ( 
.A(n_114),
.B(n_31),
.C(n_58),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_SL g194 ( 
.A(n_151),
.B(n_152),
.Y(n_194)
);

CKINVDCx20_ASAP7_75t_R g152 ( 
.A(n_126),
.Y(n_152)
);

INVx2_ASAP7_75t_L g153 ( 
.A(n_129),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_L g188 ( 
.A(n_153),
.B(n_159),
.Y(n_188)
);

NOR2xp33_ASAP7_75t_SL g158 ( 
.A(n_103),
.B(n_13),
.Y(n_158)
);

NOR2xp33_ASAP7_75t_SL g173 ( 
.A(n_158),
.B(n_13),
.Y(n_173)
);

INVx2_ASAP7_75t_L g159 ( 
.A(n_129),
.Y(n_159)
);

OAI22xp5_ASAP7_75t_SL g160 ( 
.A1(n_101),
.A2(n_19),
.B1(n_15),
.B2(n_23),
.Y(n_160)
);

AOI22xp5_ASAP7_75t_L g161 ( 
.A1(n_118),
.A2(n_12),
.B1(n_30),
.B2(n_25),
.Y(n_161)
);

OAI21xp5_ASAP7_75t_L g163 ( 
.A1(n_113),
.A2(n_98),
.B(n_23),
.Y(n_163)
);

AOI21xp5_ASAP7_75t_L g165 ( 
.A1(n_121),
.A2(n_98),
.B(n_10),
.Y(n_165)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_130),
.Y(n_167)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_167),
.Y(n_205)
);

AOI22xp5_ASAP7_75t_SL g168 ( 
.A1(n_162),
.A2(n_104),
.B1(n_101),
.B2(n_108),
.Y(n_168)
);

INVxp67_ASAP7_75t_L g211 ( 
.A(n_168),
.Y(n_211)
);

CKINVDCx20_ASAP7_75t_R g169 ( 
.A(n_156),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_SL g220 ( 
.A(n_169),
.B(n_184),
.Y(n_220)
);

NAND3xp33_ASAP7_75t_L g171 ( 
.A(n_137),
.B(n_139),
.C(n_155),
.Y(n_171)
);

NOR2xp33_ASAP7_75t_SL g216 ( 
.A(n_171),
.B(n_173),
.Y(n_216)
);

XNOR2xp5_ASAP7_75t_SL g172 ( 
.A(n_142),
.B(n_124),
.Y(n_172)
);

XNOR2xp5_ASAP7_75t_SL g213 ( 
.A(n_172),
.B(n_186),
.Y(n_213)
);

CKINVDCx20_ASAP7_75t_R g174 ( 
.A(n_139),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_SL g209 ( 
.A(n_174),
.B(n_182),
.Y(n_209)
);

CKINVDCx14_ASAP7_75t_R g210 ( 
.A(n_175),
.Y(n_210)
);

AOI22x1_ASAP7_75t_L g176 ( 
.A1(n_131),
.A2(n_108),
.B1(n_109),
.B2(n_121),
.Y(n_176)
);

OA22x2_ASAP7_75t_L g196 ( 
.A1(n_176),
.A2(n_141),
.B1(n_144),
.B2(n_146),
.Y(n_196)
);

INVxp67_ASAP7_75t_L g177 ( 
.A(n_147),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_L g215 ( 
.A(n_177),
.B(n_55),
.Y(n_215)
);

OAI21xp5_ASAP7_75t_L g178 ( 
.A1(n_133),
.A2(n_108),
.B(n_110),
.Y(n_178)
);

AOI21xp5_ASAP7_75t_L g204 ( 
.A1(n_178),
.A2(n_163),
.B(n_136),
.Y(n_204)
);

OAI22xp5_ASAP7_75t_L g208 ( 
.A1(n_179),
.A2(n_160),
.B1(n_19),
.B2(n_25),
.Y(n_208)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_164),
.Y(n_181)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_181),
.Y(n_214)
);

NOR2xp33_ASAP7_75t_SL g182 ( 
.A(n_137),
.B(n_126),
.Y(n_182)
);

AOI22xp5_ASAP7_75t_L g183 ( 
.A1(n_138),
.A2(n_122),
.B1(n_111),
.B2(n_12),
.Y(n_183)
);

OAI22xp5_ASAP7_75t_SL g202 ( 
.A1(n_183),
.A2(n_189),
.B1(n_154),
.B2(n_151),
.Y(n_202)
);

CKINVDCx20_ASAP7_75t_R g184 ( 
.A(n_164),
.Y(n_184)
);

XNOR2x1_ASAP7_75t_L g186 ( 
.A(n_135),
.B(n_122),
.Y(n_186)
);

NOR2xp33_ASAP7_75t_L g197 ( 
.A(n_187),
.B(n_165),
.Y(n_197)
);

AOI22xp5_ASAP7_75t_L g189 ( 
.A1(n_134),
.A2(n_154),
.B1(n_141),
.B2(n_148),
.Y(n_189)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_134),
.Y(n_190)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_190),
.Y(n_201)
);

OR2x2_ASAP7_75t_L g192 ( 
.A(n_155),
.B(n_13),
.Y(n_192)
);

CKINVDCx20_ASAP7_75t_R g199 ( 
.A(n_192),
.Y(n_199)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_140),
.Y(n_193)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_193),
.Y(n_203)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_196),
.Y(n_243)
);

NOR2xp33_ASAP7_75t_L g225 ( 
.A(n_197),
.B(n_187),
.Y(n_225)
);

XNOR2xp5_ASAP7_75t_L g198 ( 
.A(n_191),
.B(n_145),
.Y(n_198)
);

XNOR2xp5_ASAP7_75t_L g240 ( 
.A(n_198),
.B(n_204),
.Y(n_240)
);

INVx2_ASAP7_75t_L g200 ( 
.A(n_186),
.Y(n_200)
);

AOI22xp33_ASAP7_75t_L g230 ( 
.A1(n_200),
.A2(n_176),
.B1(n_180),
.B2(n_177),
.Y(n_230)
);

AOI22xp5_ASAP7_75t_L g224 ( 
.A1(n_202),
.A2(n_207),
.B1(n_208),
.B2(n_172),
.Y(n_224)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_188),
.Y(n_206)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_206),
.Y(n_226)
);

OAI22xp5_ASAP7_75t_SL g207 ( 
.A1(n_190),
.A2(n_161),
.B1(n_159),
.B2(n_153),
.Y(n_207)
);

AND2x2_ASAP7_75t_SL g212 ( 
.A(n_181),
.B(n_55),
.Y(n_212)
);

AOI21xp5_ASAP7_75t_L g241 ( 
.A1(n_212),
.A2(n_0),
.B(n_1),
.Y(n_241)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_215),
.Y(n_227)
);

NAND2xp5_ASAP7_75t_SL g217 ( 
.A(n_167),
.B(n_15),
.Y(n_217)
);

CKINVDCx20_ASAP7_75t_R g232 ( 
.A(n_217),
.Y(n_232)
);

AOI22xp5_ASAP7_75t_SL g218 ( 
.A1(n_178),
.A2(n_23),
.B1(n_19),
.B2(n_13),
.Y(n_218)
);

XOR2xp5_ASAP7_75t_L g234 ( 
.A(n_218),
.B(n_183),
.Y(n_234)
);

MAJIxp5_ASAP7_75t_L g219 ( 
.A(n_191),
.B(n_28),
.C(n_37),
.Y(n_219)
);

MAJIxp5_ASAP7_75t_L g221 ( 
.A(n_219),
.B(n_195),
.C(n_193),
.Y(n_221)
);

XNOR2xp5_ASAP7_75t_L g252 ( 
.A(n_221),
.B(n_234),
.Y(n_252)
);

OAI22xp5_ASAP7_75t_L g222 ( 
.A1(n_216),
.A2(n_179),
.B1(n_170),
.B2(n_166),
.Y(n_222)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_222),
.Y(n_247)
);

OAI22xp5_ASAP7_75t_L g223 ( 
.A1(n_210),
.A2(n_166),
.B1(n_185),
.B2(n_192),
.Y(n_223)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_223),
.Y(n_249)
);

OAI22xp5_ASAP7_75t_SL g244 ( 
.A1(n_224),
.A2(n_233),
.B1(n_239),
.B2(n_211),
.Y(n_244)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_225),
.Y(n_250)
);

MAJIxp5_ASAP7_75t_L g228 ( 
.A(n_219),
.B(n_195),
.C(n_194),
.Y(n_228)
);

MAJIxp5_ASAP7_75t_L g258 ( 
.A(n_228),
.B(n_229),
.C(n_235),
.Y(n_258)
);

MAJIxp5_ASAP7_75t_L g229 ( 
.A(n_198),
.B(n_189),
.C(n_180),
.Y(n_229)
);

XOR2xp5_ASAP7_75t_L g245 ( 
.A(n_230),
.B(n_215),
.Y(n_245)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_209),
.Y(n_231)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_231),
.Y(n_260)
);

AOI22xp5_ASAP7_75t_L g233 ( 
.A1(n_202),
.A2(n_176),
.B1(n_168),
.B2(n_188),
.Y(n_233)
);

MAJIxp5_ASAP7_75t_L g235 ( 
.A(n_203),
.B(n_28),
.C(n_20),
.Y(n_235)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_220),
.Y(n_236)
);

CKINVDCx20_ASAP7_75t_R g256 ( 
.A(n_236),
.Y(n_256)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_212),
.Y(n_237)
);

NAND2xp5_ASAP7_75t_SL g257 ( 
.A(n_237),
.B(n_238),
.Y(n_257)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_212),
.Y(n_238)
);

AOI22xp5_ASAP7_75t_L g239 ( 
.A1(n_211),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_239)
);

OAI21xp5_ASAP7_75t_L g261 ( 
.A1(n_241),
.A2(n_14),
.B(n_20),
.Y(n_261)
);

MAJIxp5_ASAP7_75t_L g242 ( 
.A(n_203),
.B(n_28),
.C(n_20),
.Y(n_242)
);

MAJIxp5_ASAP7_75t_L g259 ( 
.A(n_242),
.B(n_218),
.C(n_214),
.Y(n_259)
);

NOR2xp33_ASAP7_75t_L g272 ( 
.A(n_244),
.B(n_259),
.Y(n_272)
);

XOR2xp5_ASAP7_75t_L g273 ( 
.A(n_245),
.B(n_246),
.Y(n_273)
);

MAJx2_ASAP7_75t_L g246 ( 
.A(n_240),
.B(n_204),
.C(n_213),
.Y(n_246)
);

AOI22xp5_ASAP7_75t_L g248 ( 
.A1(n_243),
.A2(n_206),
.B1(n_207),
.B2(n_201),
.Y(n_248)
);

OAI22xp5_ASAP7_75t_SL g266 ( 
.A1(n_248),
.A2(n_253),
.B1(n_245),
.B2(n_259),
.Y(n_266)
);

NOR2xp33_ASAP7_75t_SL g251 ( 
.A(n_232),
.B(n_205),
.Y(n_251)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_251),
.Y(n_264)
);

INVxp67_ASAP7_75t_L g253 ( 
.A(n_235),
.Y(n_253)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_253),
.Y(n_268)
);

OAI22xp5_ASAP7_75t_SL g254 ( 
.A1(n_224),
.A2(n_199),
.B1(n_200),
.B2(n_201),
.Y(n_254)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_254),
.Y(n_270)
);

OAI22xp5_ASAP7_75t_L g255 ( 
.A1(n_243),
.A2(n_233),
.B1(n_229),
.B2(n_227),
.Y(n_255)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_255),
.Y(n_276)
);

OAI22xp5_ASAP7_75t_SL g265 ( 
.A1(n_261),
.A2(n_241),
.B1(n_239),
.B2(n_226),
.Y(n_265)
);

XOR2xp5_ASAP7_75t_L g262 ( 
.A(n_240),
.B(n_213),
.Y(n_262)
);

XOR2xp5_ASAP7_75t_L g277 ( 
.A(n_262),
.B(n_196),
.Y(n_277)
);

MAJIxp5_ASAP7_75t_L g263 ( 
.A(n_258),
.B(n_221),
.C(n_228),
.Y(n_263)
);

MAJIxp5_ASAP7_75t_L g280 ( 
.A(n_263),
.B(n_269),
.C(n_271),
.Y(n_280)
);

NOR2xp33_ASAP7_75t_L g290 ( 
.A(n_265),
.B(n_6),
.Y(n_290)
);

AOI22xp5_ASAP7_75t_L g283 ( 
.A1(n_266),
.A2(n_7),
.B1(n_10),
.B2(n_9),
.Y(n_283)
);

HB1xp67_ASAP7_75t_L g267 ( 
.A(n_258),
.Y(n_267)
);

XOR2xp5_ASAP7_75t_L g278 ( 
.A(n_267),
.B(n_274),
.Y(n_278)
);

MAJIxp5_ASAP7_75t_L g269 ( 
.A(n_252),
.B(n_247),
.C(n_249),
.Y(n_269)
);

MAJIxp5_ASAP7_75t_L g271 ( 
.A(n_252),
.B(n_234),
.C(n_242),
.Y(n_271)
);

HB1xp67_ASAP7_75t_L g274 ( 
.A(n_261),
.Y(n_274)
);

NOR2xp33_ASAP7_75t_L g275 ( 
.A(n_256),
.B(n_196),
.Y(n_275)
);

NOR2xp33_ASAP7_75t_SL g284 ( 
.A(n_275),
.B(n_7),
.Y(n_284)
);

XOR2xp5_ASAP7_75t_L g287 ( 
.A(n_277),
.B(n_273),
.Y(n_287)
);

OAI22xp5_ASAP7_75t_L g279 ( 
.A1(n_276),
.A2(n_250),
.B1(n_260),
.B2(n_257),
.Y(n_279)
);

NAND2xp5_ASAP7_75t_SL g302 ( 
.A(n_279),
.B(n_283),
.Y(n_302)
);

AOI22xp33_ASAP7_75t_L g281 ( 
.A1(n_270),
.A2(n_248),
.B1(n_196),
.B2(n_246),
.Y(n_281)
);

NOR2xp33_ASAP7_75t_L g296 ( 
.A(n_281),
.B(n_284),
.Y(n_296)
);

XNOR2x1_ASAP7_75t_L g282 ( 
.A(n_273),
.B(n_262),
.Y(n_282)
);

MAJx2_ASAP7_75t_L g295 ( 
.A(n_282),
.B(n_10),
.C(n_9),
.Y(n_295)
);

MAJIxp5_ASAP7_75t_L g285 ( 
.A(n_263),
.B(n_28),
.C(n_18),
.Y(n_285)
);

MAJIxp5_ASAP7_75t_L g292 ( 
.A(n_285),
.B(n_14),
.C(n_1),
.Y(n_292)
);

AOI21xp5_ASAP7_75t_SL g286 ( 
.A1(n_268),
.A2(n_272),
.B(n_264),
.Y(n_286)
);

OAI21xp5_ASAP7_75t_L g291 ( 
.A1(n_286),
.A2(n_289),
.B(n_20),
.Y(n_291)
);

XNOR2xp5_ASAP7_75t_L g294 ( 
.A(n_287),
.B(n_288),
.Y(n_294)
);

XNOR2xp5_ASAP7_75t_L g288 ( 
.A(n_271),
.B(n_28),
.Y(n_288)
);

MAJx2_ASAP7_75t_L g289 ( 
.A(n_266),
.B(n_269),
.C(n_277),
.Y(n_289)
);

INVxp67_ASAP7_75t_L g297 ( 
.A(n_290),
.Y(n_297)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_291),
.Y(n_304)
);

NAND2xp5_ASAP7_75t_SL g310 ( 
.A(n_292),
.B(n_295),
.Y(n_310)
);

MAJIxp5_ASAP7_75t_L g293 ( 
.A(n_280),
.B(n_14),
.C(n_10),
.Y(n_293)
);

NAND2xp5_ASAP7_75t_L g307 ( 
.A(n_293),
.B(n_298),
.Y(n_307)
);

INVxp67_ASAP7_75t_L g298 ( 
.A(n_286),
.Y(n_298)
);

AOI21xp5_ASAP7_75t_L g299 ( 
.A1(n_282),
.A2(n_8),
.B(n_6),
.Y(n_299)
);

NAND2xp5_ASAP7_75t_L g308 ( 
.A(n_299),
.B(n_300),
.Y(n_308)
);

MAJIxp5_ASAP7_75t_L g300 ( 
.A(n_278),
.B(n_14),
.C(n_8),
.Y(n_300)
);

AOI321xp33_ASAP7_75t_L g301 ( 
.A1(n_289),
.A2(n_6),
.A3(n_1),
.B1(n_2),
.B2(n_3),
.C(n_4),
.Y(n_301)
);

NOR2xp33_ASAP7_75t_SL g305 ( 
.A(n_301),
.B(n_296),
.Y(n_305)
);

MAJIxp5_ASAP7_75t_L g303 ( 
.A(n_294),
.B(n_302),
.C(n_296),
.Y(n_303)
);

HB1xp67_ASAP7_75t_L g315 ( 
.A(n_303),
.Y(n_315)
);

OAI21xp5_ASAP7_75t_L g312 ( 
.A1(n_305),
.A2(n_311),
.B(n_0),
.Y(n_312)
);

AOI22xp5_ASAP7_75t_L g306 ( 
.A1(n_297),
.A2(n_281),
.B1(n_1),
.B2(n_2),
.Y(n_306)
);

AOI21xp5_ASAP7_75t_L g314 ( 
.A1(n_306),
.A2(n_309),
.B(n_310),
.Y(n_314)
);

NOR2xp33_ASAP7_75t_L g309 ( 
.A(n_295),
.B(n_0),
.Y(n_309)
);

AOI21xp5_ASAP7_75t_SL g311 ( 
.A1(n_291),
.A2(n_0),
.B(n_2),
.Y(n_311)
);

AOI21xp5_ASAP7_75t_L g316 ( 
.A1(n_312),
.A2(n_313),
.B(n_310),
.Y(n_316)
);

OAI21xp5_ASAP7_75t_SL g313 ( 
.A1(n_307),
.A2(n_2),
.B(n_3),
.Y(n_313)
);

INVxp67_ASAP7_75t_L g317 ( 
.A(n_314),
.Y(n_317)
);

INVxp33_ASAP7_75t_L g318 ( 
.A(n_316),
.Y(n_318)
);

AO21x1_ASAP7_75t_L g319 ( 
.A1(n_318),
.A2(n_317),
.B(n_315),
.Y(n_319)
);

AOI21x1_ASAP7_75t_SL g320 ( 
.A1(n_319),
.A2(n_304),
.B(n_308),
.Y(n_320)
);

AOI21xp5_ASAP7_75t_L g321 ( 
.A1(n_320),
.A2(n_3),
.B(n_4),
.Y(n_321)
);

AO21x1_ASAP7_75t_L g322 ( 
.A1(n_321),
.A2(n_4),
.B(n_5),
.Y(n_322)
);

NOR2xp33_ASAP7_75t_L g323 ( 
.A(n_322),
.B(n_4),
.Y(n_323)
);


endmodule