module fake_jpeg_1974_n_108 (n_13, n_21, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_19, n_18, n_20, n_4, n_16, n_3, n_0, n_24, n_28, n_26, n_9, n_5, n_11, n_17, n_25, n_2, n_12, n_8, n_15, n_7, n_108);

input n_13;
input n_21;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_4;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_26;
input n_9;
input n_5;
input n_11;
input n_17;
input n_25;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_108;

wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_73;
wire n_84;
wire n_59;
wire n_98;
wire n_65;
wire n_42;
wire n_49;
wire n_76;
wire n_38;
wire n_88;
wire n_74;
wire n_31;
wire n_29;
wire n_103;
wire n_50;
wire n_57;
wire n_69;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_30;
wire n_106;
wire n_44;
wire n_75;
wire n_37;
wire n_102;
wire n_99;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_56;
wire n_79;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_101;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_95;
wire n_97;
wire n_36;
wire n_62;
wire n_43;
wire n_32;
wire n_100;
wire n_82;
wire n_96;

INVx2_ASAP7_75t_L g29 ( 
.A(n_25),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_23),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_21),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_10),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_11),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_20),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_2),
.Y(n_35)
);

INVx8_ASAP7_75t_L g36 ( 
.A(n_1),
.Y(n_36)
);

BUFx5_ASAP7_75t_L g37 ( 
.A(n_16),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_17),
.Y(n_38)
);

BUFx3_ASAP7_75t_L g39 ( 
.A(n_7),
.Y(n_39)
);

INVx4_ASAP7_75t_L g40 ( 
.A(n_37),
.Y(n_40)
);

INVx4_ASAP7_75t_L g50 ( 
.A(n_40),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_29),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_41),
.Y(n_52)
);

BUFx12f_ASAP7_75t_L g42 ( 
.A(n_36),
.Y(n_42)
);

INVx11_ASAP7_75t_L g51 ( 
.A(n_42),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g43 ( 
.A(n_35),
.B(n_0),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g49 ( 
.A(n_43),
.B(n_45),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_L g44 ( 
.A(n_29),
.B(n_39),
.Y(n_44)
);

NAND2xp5_ASAP7_75t_L g48 ( 
.A(n_44),
.B(n_19),
.Y(n_48)
);

INVx3_ASAP7_75t_L g45 ( 
.A(n_39),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_SL g46 ( 
.A(n_32),
.B(n_0),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_46),
.B(n_32),
.Y(n_53)
);

INVx6_ASAP7_75t_L g47 ( 
.A(n_41),
.Y(n_47)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_47),
.Y(n_58)
);

AND2x2_ASAP7_75t_L g60 ( 
.A(n_48),
.B(n_33),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_L g61 ( 
.A(n_53),
.B(n_54),
.Y(n_61)
);

INVx6_ASAP7_75t_L g54 ( 
.A(n_42),
.Y(n_54)
);

CKINVDCx20_ASAP7_75t_R g55 ( 
.A(n_46),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_55),
.B(n_49),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_SL g66 ( 
.A(n_56),
.B(n_57),
.Y(n_66)
);

FAx1_ASAP7_75t_SL g57 ( 
.A(n_48),
.B(n_44),
.CI(n_45),
.CON(n_57),
.SN(n_57)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_55),
.B(n_34),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_SL g70 ( 
.A(n_59),
.B(n_60),
.Y(n_70)
);

AOI22xp5_ASAP7_75t_L g62 ( 
.A1(n_52),
.A2(n_30),
.B1(n_34),
.B2(n_40),
.Y(n_62)
);

OAI22xp5_ASAP7_75t_L g75 ( 
.A1(n_62),
.A2(n_63),
.B1(n_51),
.B2(n_54),
.Y(n_75)
);

AOI22xp5_ASAP7_75t_L g63 ( 
.A1(n_52),
.A2(n_30),
.B1(n_36),
.B2(n_33),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_50),
.B(n_38),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_64),
.B(n_65),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_50),
.B(n_31),
.Y(n_65)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_58),
.Y(n_67)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_67),
.Y(n_88)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_62),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_L g83 ( 
.A(n_68),
.B(n_69),
.Y(n_83)
);

BUFx3_ASAP7_75t_L g69 ( 
.A(n_63),
.Y(n_69)
);

AOI22xp5_ASAP7_75t_L g72 ( 
.A1(n_57),
.A2(n_47),
.B1(n_42),
.B2(n_51),
.Y(n_72)
);

OAI22xp5_ASAP7_75t_SL g86 ( 
.A1(n_72),
.A2(n_76),
.B1(n_15),
.B2(n_27),
.Y(n_86)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_61),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_L g85 ( 
.A(n_73),
.B(n_5),
.Y(n_85)
);

AND2x2_ASAP7_75t_L g74 ( 
.A(n_60),
.B(n_42),
.Y(n_74)
);

INVxp67_ASAP7_75t_L g81 ( 
.A(n_74),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g87 ( 
.A(n_75),
.B(n_5),
.Y(n_87)
);

AOI22xp5_ASAP7_75t_L g76 ( 
.A1(n_57),
.A2(n_37),
.B1(n_2),
.B2(n_3),
.Y(n_76)
);

AOI22xp5_ASAP7_75t_L g77 ( 
.A1(n_72),
.A2(n_60),
.B1(n_13),
.B2(n_14),
.Y(n_77)
);

OAI22xp5_ASAP7_75t_L g93 ( 
.A1(n_77),
.A2(n_78),
.B1(n_87),
.B2(n_6),
.Y(n_93)
);

AOI22xp5_ASAP7_75t_L g78 ( 
.A1(n_68),
.A2(n_69),
.B1(n_66),
.B2(n_76),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_70),
.B(n_1),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_L g91 ( 
.A(n_79),
.B(n_82),
.Y(n_91)
);

OAI21xp5_ASAP7_75t_L g80 ( 
.A1(n_74),
.A2(n_3),
.B(n_4),
.Y(n_80)
);

XNOR2xp5_ASAP7_75t_L g89 ( 
.A(n_80),
.B(n_6),
.Y(n_89)
);

CKINVDCx20_ASAP7_75t_R g82 ( 
.A(n_71),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_73),
.B(n_4),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g92 ( 
.A(n_84),
.B(n_85),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_SL g97 ( 
.A(n_86),
.B(n_7),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g100 ( 
.A(n_89),
.B(n_90),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_L g90 ( 
.A(n_83),
.B(n_18),
.Y(n_90)
);

AO221x1_ASAP7_75t_L g98 ( 
.A1(n_93),
.A2(n_94),
.B1(n_95),
.B2(n_96),
.C(n_97),
.Y(n_98)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_88),
.Y(n_94)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_81),
.Y(n_95)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_81),
.Y(n_96)
);

OAI22xp5_ASAP7_75t_SL g99 ( 
.A1(n_90),
.A2(n_78),
.B1(n_77),
.B2(n_80),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_99),
.B(n_91),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_SL g102 ( 
.A(n_101),
.B(n_99),
.Y(n_102)
);

MAJIxp5_ASAP7_75t_L g103 ( 
.A(n_102),
.B(n_100),
.C(n_92),
.Y(n_103)
);

XNOR2xp5_ASAP7_75t_L g104 ( 
.A(n_103),
.B(n_89),
.Y(n_104)
);

AOI21xp33_ASAP7_75t_L g105 ( 
.A1(n_104),
.A2(n_98),
.B(n_9),
.Y(n_105)
);

MAJIxp5_ASAP7_75t_L g106 ( 
.A(n_105),
.B(n_12),
.C(n_22),
.Y(n_106)
);

AOI31xp33_ASAP7_75t_L g107 ( 
.A1(n_106),
.A2(n_24),
.A3(n_26),
.B(n_28),
.Y(n_107)
);

XNOR2xp5_ASAP7_75t_L g108 ( 
.A(n_107),
.B(n_8),
.Y(n_108)
);


endmodule