module fake_jpeg_16536_n_49 (n_13, n_21, n_1, n_10, n_6, n_14, n_19, n_18, n_20, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_49);

input n_13;
input n_21;
input n_1;
input n_10;
input n_6;
input n_14;
input n_19;
input n_18;
input n_20;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_49;

wire n_33;
wire n_45;
wire n_23;
wire n_27;
wire n_47;
wire n_22;
wire n_40;
wire n_35;
wire n_48;
wire n_46;
wire n_41;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_24;
wire n_28;
wire n_38;
wire n_44;
wire n_26;
wire n_36;
wire n_31;
wire n_25;
wire n_29;
wire n_37;
wire n_43;
wire n_32;

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_17),
.Y(n_22)
);

BUFx3_ASAP7_75t_L g23 ( 
.A(n_6),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_1),
.Y(n_24)
);

BUFx12f_ASAP7_75t_L g25 ( 
.A(n_4),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_18),
.Y(n_26)
);

INVx2_ASAP7_75t_L g27 ( 
.A(n_9),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_7),
.Y(n_28)
);

OAI22xp5_ASAP7_75t_L g29 ( 
.A1(n_27),
.A2(n_11),
.B1(n_20),
.B2(n_19),
.Y(n_29)
);

AOI22xp5_ASAP7_75t_L g38 ( 
.A1(n_29),
.A2(n_14),
.B1(n_16),
.B2(n_15),
.Y(n_38)
);

NAND2xp5_ASAP7_75t_L g30 ( 
.A(n_24),
.B(n_0),
.Y(n_30)
);

NAND2xp5_ASAP7_75t_L g39 ( 
.A(n_30),
.B(n_31),
.Y(n_39)
);

NAND2xp5_ASAP7_75t_L g31 ( 
.A(n_24),
.B(n_0),
.Y(n_31)
);

MAJIxp5_ASAP7_75t_L g32 ( 
.A(n_28),
.B(n_21),
.C(n_10),
.Y(n_32)
);

NOR2xp33_ASAP7_75t_SL g35 ( 
.A(n_32),
.B(n_33),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_SL g33 ( 
.A(n_23),
.B(n_1),
.Y(n_33)
);

INVx2_ASAP7_75t_SL g34 ( 
.A(n_25),
.Y(n_34)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_34),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g37 ( 
.A(n_32),
.B(n_2),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g42 ( 
.A(n_37),
.B(n_3),
.Y(n_42)
);

OAI22xp5_ASAP7_75t_SL g40 ( 
.A1(n_38),
.A2(n_2),
.B1(n_3),
.B2(n_4),
.Y(n_40)
);

AOI22xp5_ASAP7_75t_L g43 ( 
.A1(n_40),
.A2(n_41),
.B1(n_42),
.B2(n_5),
.Y(n_43)
);

INVxp67_ASAP7_75t_L g41 ( 
.A(n_36),
.Y(n_41)
);

OAI22xp5_ASAP7_75t_SL g44 ( 
.A1(n_43),
.A2(n_39),
.B1(n_38),
.B2(n_41),
.Y(n_44)
);

XNOR2xp5_ASAP7_75t_L g45 ( 
.A(n_44),
.B(n_35),
.Y(n_45)
);

OAI21xp5_ASAP7_75t_SL g46 ( 
.A1(n_45),
.A2(n_25),
.B(n_5),
.Y(n_46)
);

OAI22xp5_ASAP7_75t_SL g47 ( 
.A1(n_46),
.A2(n_34),
.B1(n_12),
.B2(n_13),
.Y(n_47)
);

AO21x1_ASAP7_75t_L g48 ( 
.A1(n_47),
.A2(n_8),
.B(n_28),
.Y(n_48)
);

AOI21xp5_ASAP7_75t_L g49 ( 
.A1(n_48),
.A2(n_22),
.B(n_26),
.Y(n_49)
);


endmodule