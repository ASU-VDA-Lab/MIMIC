module real_jpeg_15992_n_14 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_2, n_13, n_6, n_7, n_3, n_10, n_9, n_14);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_2;
input n_13;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_14;

wire n_384;
wire n_37;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_300;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_199;
wire n_95;
wire n_238;
wire n_67;
wire n_350;
wire n_235;
wire n_107;
wire n_369;
wire n_376;
wire n_354;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_355;
wire n_123;
wire n_50;
wire n_186;
wire n_137;
wire n_72;
wire n_171;
wire n_151;
wire n_272;
wire n_203;
wire n_198;
wire n_23;
wire n_362;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_326;
wire n_339;
wire n_80;
wire n_30;
wire n_328;
wire n_149;
wire n_332;
wire n_366;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_353;
wire n_230;
wire n_128;
wire n_202;
wire n_216;
wire n_367;
wire n_127;
wire n_365;
wire n_356;
wire n_36;
wire n_102;
wire n_81;
wire n_101;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_348;
wire n_252;
wire n_363;
wire n_310;
wire n_345;
wire n_78;
wire n_83;
wire n_288;
wire n_221;
wire n_393;
wire n_104;
wire n_153;
wire n_337;
wire n_131;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_378;
wire n_200;
wire n_335;
wire n_214;
wire n_113;
wire n_251;
wire n_139;
wire n_33;
wire n_175;
wire n_338;
wire n_156;
wire n_387;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_390;
wire n_77;
wire n_219;
wire n_372;
wire n_122;
wire n_19;
wire n_262;
wire n_334;
wire n_17;
wire n_383;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_371;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_382;
wire n_20;
wire n_278;
wire n_314;
wire n_103;
wire n_232;
wire n_212;
wire n_284;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_213;
wire n_25;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_386;
wire n_341;
wire n_331;
wire n_49;
wire n_68;
wire n_395;
wire n_146;
wire n_286;
wire n_323;
wire n_176;
wire n_166;
wire n_215;
wire n_312;
wire n_325;
wire n_316;
wire n_307;
wire n_161;
wire n_207;
wire n_357;
wire n_237;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_380;
wire n_140;
wire n_126;
wire n_342;
wire n_120;
wire n_155;
wire n_319;
wire n_93;
wire n_242;
wire n_142;
wire n_76;
wire n_79;
wire n_282;
wire n_147;
wire n_359;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_18;
wire n_145;
wire n_266;
wire n_377;
wire n_109;
wire n_391;
wire n_148;
wire n_373;
wire n_396;
wire n_392;
wire n_375;
wire n_196;
wire n_298;
wire n_330;
wire n_333;
wire n_152;
wire n_270;
wire n_159;
wire n_347;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_336;
wire n_258;
wire n_150;
wire n_41;
wire n_74;
wire n_204;
wire n_158;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_75;
wire n_346;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_119;
wire n_283;
wire n_181;
wire n_358;
wire n_256;
wire n_253;
wire n_273;
wire n_16;
wire n_54;
wire n_168;
wire n_38;
wire n_385;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_349;
wire n_343;
wire n_292;
wire n_64;
wire n_291;
wire n_236;
wire n_370;
wire n_276;
wire n_374;
wire n_287;
wire n_388;
wire n_174;
wire n_255;
wire n_243;
wire n_299;
wire n_352;
wire n_56;
wire n_293;
wire n_275;
wire n_381;
wire n_227;
wire n_229;
wire n_379;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_360;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_45;
wire n_268;
wire n_42;
wire n_313;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_143;
wire n_351;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_303;
wire n_321;
wire n_100;
wire n_368;
wire n_51;
wire n_205;
wire n_361;
wire n_261;
wire n_86;
wire n_324;
wire n_70;
wire n_32;
wire n_228;
wire n_389;
wire n_15;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_394;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_169;
wire n_88;
wire n_167;
wire n_295;
wire n_133;
wire n_257;
wire n_344;
wire n_210;
wire n_206;
wire n_85;
wire n_96;
wire n_308;
wire n_364;

AOI21xp5_ASAP7_75t_L g14 ( 
.A1(n_0),
.A2(n_15),
.B(n_395),
.Y(n_14)
);

NOR2xp33_ASAP7_75t_L g395 ( 
.A(n_0),
.B(n_396),
.Y(n_395)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_1),
.Y(n_27)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_1),
.Y(n_59)
);

NAND2x1_ASAP7_75t_L g23 ( 
.A(n_2),
.B(n_24),
.Y(n_23)
);

AND2x2_ASAP7_75t_L g54 ( 
.A(n_2),
.B(n_55),
.Y(n_54)
);

AND2x2_ASAP7_75t_L g57 ( 
.A(n_2),
.B(n_58),
.Y(n_57)
);

AND2x2_ASAP7_75t_L g67 ( 
.A(n_2),
.B(n_68),
.Y(n_67)
);

AND2x2_ASAP7_75t_L g78 ( 
.A(n_2),
.B(n_79),
.Y(n_78)
);

NAND2x1_ASAP7_75t_SL g83 ( 
.A(n_2),
.B(n_84),
.Y(n_83)
);

AND2x2_ASAP7_75t_L g118 ( 
.A(n_2),
.B(n_119),
.Y(n_118)
);

AND2x4_ASAP7_75t_L g120 ( 
.A(n_2),
.B(n_121),
.Y(n_120)
);

BUFx6f_ASAP7_75t_L g70 ( 
.A(n_3),
.Y(n_70)
);

BUFx5_ASAP7_75t_L g119 ( 
.A(n_4),
.Y(n_119)
);

BUFx3_ASAP7_75t_L g194 ( 
.A(n_4),
.Y(n_194)
);

INVx2_ASAP7_75t_L g208 ( 
.A(n_4),
.Y(n_208)
);

CKINVDCx20_ASAP7_75t_R g396 ( 
.A(n_5),
.Y(n_396)
);

AND2x2_ASAP7_75t_L g25 ( 
.A(n_6),
.B(n_26),
.Y(n_25)
);

INVx2_ASAP7_75t_SL g38 ( 
.A(n_6),
.Y(n_38)
);

NAND2xp5_ASAP7_75t_SL g48 ( 
.A(n_6),
.B(n_49),
.Y(n_48)
);

AND2x2_ASAP7_75t_L g63 ( 
.A(n_6),
.B(n_64),
.Y(n_63)
);

AND2x2_ASAP7_75t_L g85 ( 
.A(n_6),
.B(n_86),
.Y(n_85)
);

AND2x2_ASAP7_75t_L g153 ( 
.A(n_6),
.B(n_79),
.Y(n_153)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_7),
.Y(n_55)
);

INVx3_ASAP7_75t_L g87 ( 
.A(n_7),
.Y(n_87)
);

BUFx6f_ASAP7_75t_L g106 ( 
.A(n_7),
.Y(n_106)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_7),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_L g29 ( 
.A(n_8),
.B(n_30),
.Y(n_29)
);

NAND2xp5_ASAP7_75t_L g34 ( 
.A(n_8),
.B(n_35),
.Y(n_34)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_8),
.B(n_90),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g103 ( 
.A(n_8),
.B(n_104),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_8),
.B(n_128),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_L g196 ( 
.A(n_8),
.B(n_197),
.Y(n_196)
);

NAND2xp5_ASAP7_75t_SL g203 ( 
.A(n_8),
.B(n_204),
.Y(n_203)
);

AND2x2_ASAP7_75t_L g216 ( 
.A(n_8),
.B(n_217),
.Y(n_216)
);

AND2x2_ASAP7_75t_SL g154 ( 
.A(n_9),
.B(n_155),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_SL g157 ( 
.A(n_9),
.B(n_158),
.Y(n_157)
);

AND2x2_ASAP7_75t_SL g163 ( 
.A(n_9),
.B(n_164),
.Y(n_163)
);

AND2x2_ASAP7_75t_L g169 ( 
.A(n_9),
.B(n_170),
.Y(n_169)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_9),
.Y(n_178)
);

AND2x2_ASAP7_75t_SL g189 ( 
.A(n_9),
.B(n_190),
.Y(n_189)
);

AND2x2_ASAP7_75t_L g297 ( 
.A(n_9),
.B(n_298),
.Y(n_297)
);

NAND2xp5_ASAP7_75t_L g307 ( 
.A(n_9),
.B(n_308),
.Y(n_307)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_10),
.Y(n_36)
);

INVx6_ASAP7_75t_L g65 ( 
.A(n_10),
.Y(n_65)
);

BUFx6f_ASAP7_75t_L g84 ( 
.A(n_10),
.Y(n_84)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_11),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_11),
.Y(n_43)
);

BUFx12f_ASAP7_75t_L g79 ( 
.A(n_12),
.Y(n_79)
);

BUFx4f_ASAP7_75t_L g199 ( 
.A(n_12),
.Y(n_199)
);

BUFx8_ASAP7_75t_L g24 ( 
.A(n_13),
.Y(n_24)
);

INVx2_ASAP7_75t_L g51 ( 
.A(n_13),
.Y(n_51)
);

BUFx5_ASAP7_75t_L g190 ( 
.A(n_13),
.Y(n_190)
);

XOR2xp5_ASAP7_75t_L g15 ( 
.A(n_16),
.B(n_142),
.Y(n_15)
);

NOR2xp33_ASAP7_75t_L g16 ( 
.A(n_17),
.B(n_141),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_18),
.Y(n_17)
);

NAND2xp5_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_122),
.Y(n_18)
);

NOR2xp33_ASAP7_75t_L g141 ( 
.A(n_19),
.B(n_122),
.Y(n_141)
);

MAJIxp5_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_73),
.C(n_91),
.Y(n_19)
);

XOR2xp5_ASAP7_75t_L g390 ( 
.A(n_20),
.B(n_73),
.Y(n_390)
);

AOI22xp5_ASAP7_75t_L g20 ( 
.A1(n_21),
.A2(n_45),
.B1(n_46),
.B2(n_72),
.Y(n_20)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_21),
.Y(n_72)
);

XNOR2xp5_ASAP7_75t_L g21 ( 
.A(n_22),
.B(n_32),
.Y(n_21)
);

MAJIxp5_ASAP7_75t_L g139 ( 
.A(n_22),
.B(n_34),
.C(n_37),
.Y(n_139)
);

MAJIxp5_ASAP7_75t_L g22 ( 
.A(n_23),
.B(n_25),
.C(n_28),
.Y(n_22)
);

AOI22xp5_ASAP7_75t_L g111 ( 
.A1(n_23),
.A2(n_112),
.B1(n_113),
.B2(n_115),
.Y(n_111)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_23),
.Y(n_115)
);

MAJIxp5_ASAP7_75t_L g116 ( 
.A(n_23),
.B(n_117),
.C(n_120),
.Y(n_116)
);

MAJx2_ASAP7_75t_L g174 ( 
.A(n_23),
.B(n_54),
.C(n_67),
.Y(n_174)
);

OAI22xp5_ASAP7_75t_SL g241 ( 
.A1(n_23),
.A2(n_75),
.B1(n_76),
.B2(n_115),
.Y(n_241)
);

OAI22xp5_ASAP7_75t_L g279 ( 
.A1(n_23),
.A2(n_115),
.B1(n_120),
.B2(n_138),
.Y(n_279)
);

MAJIxp5_ASAP7_75t_L g99 ( 
.A(n_25),
.B(n_100),
.C(n_102),
.Y(n_99)
);

OAI22xp5_ASAP7_75t_SL g113 ( 
.A1(n_25),
.A2(n_28),
.B1(n_29),
.B2(n_114),
.Y(n_113)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_25),
.Y(n_114)
);

O2A1O1Ixp5_ASAP7_75t_L g162 ( 
.A1(n_25),
.A2(n_67),
.B(n_163),
.C(n_168),
.Y(n_162)
);

AO22x1_ASAP7_75t_L g267 ( 
.A1(n_25),
.A2(n_102),
.B1(n_103),
.B2(n_114),
.Y(n_267)
);

OAI22xp5_ASAP7_75t_SL g347 ( 
.A1(n_25),
.A2(n_66),
.B1(n_67),
.B2(n_114),
.Y(n_347)
);

BUFx2_ASAP7_75t_L g158 ( 
.A(n_26),
.Y(n_158)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_27),
.Y(n_26)
);

BUFx5_ASAP7_75t_L g90 ( 
.A(n_27),
.Y(n_90)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_29),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_31),
.Y(n_30)
);

OAI22xp5_ASAP7_75t_SL g32 ( 
.A1(n_33),
.A2(n_34),
.B1(n_37),
.B2(n_44),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_34),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_36),
.Y(n_35)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_37),
.Y(n_44)
);

MAJIxp5_ASAP7_75t_L g77 ( 
.A(n_37),
.B(n_66),
.C(n_78),
.Y(n_77)
);

AOI22xp5_ASAP7_75t_L g95 ( 
.A1(n_37),
.A2(n_44),
.B1(n_96),
.B2(n_97),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g202 ( 
.A(n_37),
.B(n_203),
.Y(n_202)
);

OAI21xp5_ASAP7_75t_L g244 ( 
.A1(n_37),
.A2(n_202),
.B(n_203),
.Y(n_244)
);

OR2x2_ASAP7_75t_L g37 ( 
.A(n_38),
.B(n_39),
.Y(n_37)
);

OR2x4_ASAP7_75t_SL g101 ( 
.A(n_38),
.B(n_69),
.Y(n_101)
);

OR2x2_ASAP7_75t_L g192 ( 
.A(n_38),
.B(n_193),
.Y(n_192)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_40),
.Y(n_39)
);

INVx2_ASAP7_75t_L g40 ( 
.A(n_41),
.Y(n_40)
);

INVx3_ASAP7_75t_L g41 ( 
.A(n_42),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_43),
.Y(n_42)
);

BUFx5_ASAP7_75t_L g121 ( 
.A(n_43),
.Y(n_121)
);

BUFx6f_ASAP7_75t_L g180 ( 
.A(n_43),
.Y(n_180)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_46),
.Y(n_45)
);

XOR2xp5_ASAP7_75t_L g46 ( 
.A(n_47),
.B(n_60),
.Y(n_46)
);

MAJIxp5_ASAP7_75t_L g140 ( 
.A(n_47),
.B(n_60),
.C(n_72),
.Y(n_140)
);

XNOR2xp5_ASAP7_75t_L g47 ( 
.A(n_48),
.B(n_52),
.Y(n_47)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_48),
.Y(n_132)
);

XNOR2xp5_ASAP7_75t_L g227 ( 
.A(n_48),
.B(n_228),
.Y(n_227)
);

OAI21xp5_ASAP7_75t_SL g265 ( 
.A1(n_48),
.A2(n_118),
.B(n_153),
.Y(n_265)
);

INVx5_ASAP7_75t_L g49 ( 
.A(n_50),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_51),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g129 ( 
.A(n_51),
.Y(n_129)
);

OAI22xp5_ASAP7_75t_L g52 ( 
.A1(n_53),
.A2(n_54),
.B1(n_56),
.B2(n_57),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_L g61 ( 
.A(n_53),
.B(n_62),
.Y(n_61)
);

OAI22xp5_ASAP7_75t_SL g182 ( 
.A1(n_53),
.A2(n_54),
.B1(n_136),
.B2(n_137),
.Y(n_182)
);

OAI22xp5_ASAP7_75t_SL g334 ( 
.A1(n_53),
.A2(n_54),
.B1(n_169),
.B2(n_311),
.Y(n_334)
);

INVx1_ASAP7_75t_SL g53 ( 
.A(n_54),
.Y(n_53)
);

AND2x2_ASAP7_75t_L g71 ( 
.A(n_54),
.B(n_63),
.Y(n_71)
);

XNOR2xp5_ASAP7_75t_L g75 ( 
.A(n_54),
.B(n_66),
.Y(n_75)
);

MAJIxp5_ASAP7_75t_L g131 ( 
.A(n_54),
.B(n_56),
.C(n_132),
.Y(n_131)
);

AND2x2_ASAP7_75t_L g168 ( 
.A(n_54),
.B(n_169),
.Y(n_168)
);

O2A1O1Ixp33_ASAP7_75t_SL g321 ( 
.A1(n_54),
.A2(n_168),
.B(n_169),
.C(n_322),
.Y(n_321)
);

OAI22xp5_ASAP7_75t_SL g232 ( 
.A1(n_56),
.A2(n_57),
.B1(n_154),
.B2(n_156),
.Y(n_232)
);

AOI22xp5_ASAP7_75t_L g293 ( 
.A1(n_56),
.A2(n_57),
.B1(n_100),
.B2(n_101),
.Y(n_293)
);

MAJIxp5_ASAP7_75t_L g318 ( 
.A(n_56),
.B(n_101),
.C(n_294),
.Y(n_318)
);

INVx2_ASAP7_75t_SL g56 ( 
.A(n_57),
.Y(n_56)
);

XNOR2xp5_ASAP7_75t_L g136 ( 
.A(n_57),
.B(n_62),
.Y(n_136)
);

AO21x1_ASAP7_75t_L g225 ( 
.A1(n_57),
.A2(n_61),
.B(n_71),
.Y(n_225)
);

MAJIxp5_ASAP7_75t_L g253 ( 
.A(n_57),
.B(n_85),
.C(n_154),
.Y(n_253)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_59),
.Y(n_58)
);

AOI21xp5_ASAP7_75t_L g60 ( 
.A1(n_61),
.A2(n_66),
.B(n_71),
.Y(n_60)
);

OAI22xp5_ASAP7_75t_SL g74 ( 
.A1(n_62),
.A2(n_63),
.B1(n_75),
.B2(n_76),
.Y(n_74)
);

INVx1_ASAP7_75t_SL g62 ( 
.A(n_63),
.Y(n_62)
);

INVx4_ASAP7_75t_L g64 ( 
.A(n_65),
.Y(n_64)
);

INVx3_ASAP7_75t_SL g155 ( 
.A(n_65),
.Y(n_155)
);

OAI22xp5_ASAP7_75t_SL g97 ( 
.A1(n_66),
.A2(n_67),
.B1(n_78),
.B2(n_98),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_SL g329 ( 
.A(n_66),
.B(n_330),
.Y(n_329)
);

NOR2xp33_ASAP7_75t_L g331 ( 
.A(n_66),
.B(n_330),
.Y(n_331)
);

INVx2_ASAP7_75t_SL g66 ( 
.A(n_67),
.Y(n_66)
);

INVx3_ASAP7_75t_L g68 ( 
.A(n_69),
.Y(n_68)
);

INVx2_ASAP7_75t_L g217 ( 
.A(n_69),
.Y(n_217)
);

INVx6_ASAP7_75t_L g69 ( 
.A(n_70),
.Y(n_69)
);

BUFx6f_ASAP7_75t_L g172 ( 
.A(n_70),
.Y(n_172)
);

MAJIxp5_ASAP7_75t_L g73 ( 
.A(n_74),
.B(n_77),
.C(n_80),
.Y(n_73)
);

XOR2xp5_ASAP7_75t_L g384 ( 
.A(n_74),
.B(n_385),
.Y(n_384)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_75),
.Y(n_76)
);

OAI22xp5_ASAP7_75t_SL g385 ( 
.A1(n_77),
.A2(n_80),
.B1(n_81),
.B2(n_386),
.Y(n_385)
);

INVx1_ASAP7_75t_L g386 ( 
.A(n_77),
.Y(n_386)
);

INVx2_ASAP7_75t_SL g98 ( 
.A(n_78),
.Y(n_98)
);

NAND2x1_ASAP7_75t_L g243 ( 
.A(n_78),
.B(n_118),
.Y(n_243)
);

OAI21xp5_ASAP7_75t_L g269 ( 
.A1(n_78),
.A2(n_118),
.B(n_243),
.Y(n_269)
);

OAI22xp5_ASAP7_75t_SL g353 ( 
.A1(n_78),
.A2(n_98),
.B1(n_192),
.B2(n_200),
.Y(n_353)
);

INVx3_ASAP7_75t_L g299 ( 
.A(n_79),
.Y(n_299)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_81),
.Y(n_80)
);

MAJIxp5_ASAP7_75t_L g81 ( 
.A(n_82),
.B(n_85),
.C(n_88),
.Y(n_81)
);

AOI22xp5_ASAP7_75t_L g107 ( 
.A1(n_82),
.A2(n_83),
.B1(n_108),
.B2(n_109),
.Y(n_107)
);

OAI22xp5_ASAP7_75t_SL g268 ( 
.A1(n_82),
.A2(n_83),
.B1(n_269),
.B2(n_270),
.Y(n_268)
);

OAI22xp5_ASAP7_75t_SL g343 ( 
.A1(n_82),
.A2(n_83),
.B1(n_176),
.B2(n_177),
.Y(n_343)
);

INVx1_ASAP7_75t_SL g82 ( 
.A(n_83),
.Y(n_82)
);

MAJIxp5_ASAP7_75t_L g117 ( 
.A(n_83),
.B(n_98),
.C(n_118),
.Y(n_117)
);

MAJIxp5_ASAP7_75t_L g242 ( 
.A(n_83),
.B(n_177),
.C(n_243),
.Y(n_242)
);

OAI22xp5_ASAP7_75t_SL g109 ( 
.A1(n_85),
.A2(n_88),
.B1(n_89),
.B2(n_110),
.Y(n_109)
);

INVx1_ASAP7_75t_SL g110 ( 
.A(n_85),
.Y(n_110)
);

AOI22xp5_ASAP7_75t_L g314 ( 
.A1(n_85),
.A2(n_110),
.B1(n_315),
.B2(n_316),
.Y(n_314)
);

MAJIxp5_ASAP7_75t_L g351 ( 
.A(n_85),
.B(n_120),
.C(n_210),
.Y(n_351)
);

INVx2_ASAP7_75t_L g86 ( 
.A(n_87),
.Y(n_86)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_89),
.Y(n_88)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_92),
.Y(n_91)
);

XNOR2xp5_ASAP7_75t_L g389 ( 
.A(n_92),
.B(n_390),
.Y(n_389)
);

MAJIxp5_ASAP7_75t_L g92 ( 
.A(n_93),
.B(n_111),
.C(n_116),
.Y(n_92)
);

INVxp33_ASAP7_75t_L g93 ( 
.A(n_94),
.Y(n_93)
);

XNOR2xp5_ASAP7_75t_L g382 ( 
.A(n_94),
.B(n_383),
.Y(n_382)
);

MAJIxp5_ASAP7_75t_L g94 ( 
.A(n_95),
.B(n_99),
.C(n_107),
.Y(n_94)
);

XNOR2xp5_ASAP7_75t_L g274 ( 
.A(n_95),
.B(n_275),
.Y(n_274)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_97),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g306 ( 
.A(n_98),
.B(n_307),
.Y(n_306)
);

XOR2xp5_ASAP7_75t_L g275 ( 
.A(n_99),
.B(n_107),
.Y(n_275)
);

OAI22xp5_ASAP7_75t_SL g175 ( 
.A1(n_100),
.A2(n_101),
.B1(n_176),
.B2(n_177),
.Y(n_175)
);

MAJIxp5_ASAP7_75t_L g212 ( 
.A(n_100),
.B(n_174),
.C(n_176),
.Y(n_212)
);

CKINVDCx14_ASAP7_75t_R g100 ( 
.A(n_101),
.Y(n_100)
);

XNOR2xp5_ASAP7_75t_L g266 ( 
.A(n_101),
.B(n_267),
.Y(n_266)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_103),
.Y(n_102)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_105),
.Y(n_104)
);

INVx6_ASAP7_75t_L g105 ( 
.A(n_106),
.Y(n_105)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_109),
.Y(n_108)
);

XNOR2xp5_ASAP7_75t_L g231 ( 
.A(n_110),
.B(n_232),
.Y(n_231)
);

XNOR2xp5_ASAP7_75t_L g383 ( 
.A(n_111),
.B(n_116),
.Y(n_383)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_113),
.Y(n_112)
);

XNOR2xp5_ASAP7_75t_L g278 ( 
.A(n_117),
.B(n_279),
.Y(n_278)
);

NAND2xp5_ASAP7_75t_SL g160 ( 
.A(n_118),
.B(n_153),
.Y(n_160)
);

OAI22xp5_ASAP7_75t_SL g228 ( 
.A1(n_118),
.A2(n_152),
.B1(n_153),
.B2(n_229),
.Y(n_228)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_118),
.Y(n_229)
);

OAI22xp5_ASAP7_75t_SL g301 ( 
.A1(n_118),
.A2(n_229),
.B1(n_297),
.B2(n_302),
.Y(n_301)
);

OAI22xp5_ASAP7_75t_SL g135 ( 
.A1(n_120),
.A2(n_136),
.B1(n_137),
.B2(n_138),
.Y(n_135)
);

INVx2_ASAP7_75t_SL g138 ( 
.A(n_120),
.Y(n_138)
);

AOI22x1_ASAP7_75t_SL g215 ( 
.A1(n_120),
.A2(n_138),
.B1(n_216),
.B2(n_218),
.Y(n_215)
);

MAJIxp5_ASAP7_75t_L g250 ( 
.A(n_120),
.B(n_214),
.C(n_216),
.Y(n_250)
);

XNOR2xp5_ASAP7_75t_L g255 ( 
.A(n_120),
.B(n_188),
.Y(n_255)
);

XNOR2xp5_ASAP7_75t_L g316 ( 
.A(n_120),
.B(n_157),
.Y(n_316)
);

XOR2xp5_ASAP7_75t_L g122 ( 
.A(n_123),
.B(n_140),
.Y(n_122)
);

XOR2xp5_ASAP7_75t_L g123 ( 
.A(n_124),
.B(n_139),
.Y(n_123)
);

OAI22xp5_ASAP7_75t_SL g124 ( 
.A1(n_125),
.A2(n_126),
.B1(n_134),
.B2(n_135),
.Y(n_124)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_126),
.Y(n_125)
);

AOI22xp5_ASAP7_75t_L g126 ( 
.A1(n_127),
.A2(n_130),
.B1(n_131),
.B2(n_133),
.Y(n_126)
);

CKINVDCx16_ASAP7_75t_R g133 ( 
.A(n_127),
.Y(n_133)
);

INVx4_ASAP7_75t_L g128 ( 
.A(n_129),
.Y(n_128)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_131),
.Y(n_130)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_135),
.Y(n_134)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_136),
.Y(n_137)
);

MAJIxp5_ASAP7_75t_L g280 ( 
.A(n_138),
.B(n_188),
.C(n_252),
.Y(n_280)
);

OAI21xp5_ASAP7_75t_SL g142 ( 
.A1(n_143),
.A2(n_387),
.B(n_392),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_L g143 ( 
.A(n_144),
.B(n_376),
.Y(n_143)
);

OAI321xp33_ASAP7_75t_L g144 ( 
.A1(n_145),
.A2(n_245),
.A3(n_286),
.B1(n_369),
.B2(n_370),
.C(n_375),
.Y(n_144)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_146),
.Y(n_145)
);

AOI31xp33_ASAP7_75t_L g370 ( 
.A1(n_146),
.A2(n_282),
.A3(n_371),
.B(n_374),
.Y(n_370)
);

OR2x2_ASAP7_75t_L g146 ( 
.A(n_147),
.B(n_233),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_L g372 ( 
.A(n_147),
.B(n_233),
.Y(n_372)
);

XOR2xp5_ASAP7_75t_L g147 ( 
.A(n_148),
.B(n_183),
.Y(n_147)
);

MAJIxp5_ASAP7_75t_L g285 ( 
.A(n_148),
.B(n_184),
.C(n_222),
.Y(n_285)
);

MAJIxp5_ASAP7_75t_L g148 ( 
.A(n_149),
.B(n_173),
.C(n_181),
.Y(n_148)
);

XOR2xp5_ASAP7_75t_L g234 ( 
.A(n_149),
.B(n_235),
.Y(n_234)
);

MAJIxp5_ASAP7_75t_L g149 ( 
.A(n_150),
.B(n_159),
.C(n_161),
.Y(n_149)
);

XNOR2xp5_ASAP7_75t_L g360 ( 
.A(n_150),
.B(n_361),
.Y(n_360)
);

XNOR2xp5_ASAP7_75t_SL g150 ( 
.A(n_151),
.B(n_157),
.Y(n_150)
);

OAI22xp5_ASAP7_75t_SL g151 ( 
.A1(n_152),
.A2(n_153),
.B1(n_154),
.B2(n_156),
.Y(n_151)
);

OAI22xp5_ASAP7_75t_SL g322 ( 
.A1(n_152),
.A2(n_153),
.B1(n_307),
.B2(n_323),
.Y(n_322)
);

INVx1_ASAP7_75t_SL g152 ( 
.A(n_153),
.Y(n_152)
);

MAJIxp5_ASAP7_75t_L g209 ( 
.A(n_153),
.B(n_154),
.C(n_210),
.Y(n_209)
);

CKINVDCx16_ASAP7_75t_R g156 ( 
.A(n_154),
.Y(n_156)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_157),
.Y(n_210)
);

XNOR2xp5_ASAP7_75t_L g361 ( 
.A(n_159),
.B(n_162),
.Y(n_361)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_160),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_SL g264 ( 
.A(n_160),
.B(n_265),
.Y(n_264)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_162),
.Y(n_161)
);

AOI22xp5_ASAP7_75t_L g292 ( 
.A1(n_163),
.A2(n_293),
.B1(n_294),
.B2(n_295),
.Y(n_292)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_163),
.Y(n_294)
);

OAI22xp5_ASAP7_75t_L g346 ( 
.A1(n_163),
.A2(n_294),
.B1(n_347),
.B2(n_348),
.Y(n_346)
);

INVx3_ASAP7_75t_L g164 ( 
.A(n_165),
.Y(n_164)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_166),
.Y(n_165)
);

INVx2_ASAP7_75t_L g166 ( 
.A(n_167),
.Y(n_166)
);

OAI22xp5_ASAP7_75t_L g310 ( 
.A1(n_169),
.A2(n_269),
.B1(n_270),
.B2(n_311),
.Y(n_310)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_169),
.Y(n_311)
);

OAI21xp5_ASAP7_75t_SL g344 ( 
.A1(n_169),
.A2(n_270),
.B(n_306),
.Y(n_344)
);

INVx2_ASAP7_75t_L g170 ( 
.A(n_171),
.Y(n_170)
);

INVx3_ASAP7_75t_L g171 ( 
.A(n_172),
.Y(n_171)
);

OAI22xp5_ASAP7_75t_L g235 ( 
.A1(n_173),
.A2(n_181),
.B1(n_182),
.B2(n_236),
.Y(n_235)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_173),
.Y(n_236)
);

XNOR2xp5_ASAP7_75t_L g173 ( 
.A(n_174),
.B(n_175),
.Y(n_173)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_177),
.Y(n_176)
);

OR2x2_ASAP7_75t_L g177 ( 
.A(n_178),
.B(n_179),
.Y(n_177)
);

INVx2_ASAP7_75t_L g179 ( 
.A(n_180),
.Y(n_179)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_182),
.Y(n_181)
);

OAI22xp5_ASAP7_75t_SL g183 ( 
.A1(n_184),
.A2(n_185),
.B1(n_221),
.B2(n_222),
.Y(n_183)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_185),
.Y(n_184)
);

XNOR2xp5_ASAP7_75t_L g185 ( 
.A(n_186),
.B(n_211),
.Y(n_185)
);

INVxp67_ASAP7_75t_L g260 ( 
.A(n_186),
.Y(n_260)
);

MAJIxp5_ASAP7_75t_L g186 ( 
.A(n_187),
.B(n_201),
.C(n_209),
.Y(n_186)
);

XOR2xp5_ASAP7_75t_L g237 ( 
.A(n_187),
.B(n_238),
.Y(n_237)
);

XNOR2xp5_ASAP7_75t_L g187 ( 
.A(n_188),
.B(n_191),
.Y(n_187)
);

INVx1_ASAP7_75t_SL g188 ( 
.A(n_189),
.Y(n_188)
);

MAJIxp5_ASAP7_75t_L g214 ( 
.A(n_189),
.B(n_192),
.C(n_196),
.Y(n_214)
);

OAI22xp5_ASAP7_75t_SL g191 ( 
.A1(n_192),
.A2(n_195),
.B1(n_196),
.B2(n_200),
.Y(n_191)
);

INVx1_ASAP7_75t_SL g200 ( 
.A(n_192),
.Y(n_200)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_194),
.Y(n_193)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_196),
.Y(n_195)
);

INVx2_ASAP7_75t_L g197 ( 
.A(n_198),
.Y(n_197)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_199),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_L g296 ( 
.A(n_200),
.B(n_297),
.Y(n_296)
);

OAI21xp5_ASAP7_75t_SL g330 ( 
.A1(n_200),
.A2(n_296),
.B(n_297),
.Y(n_330)
);

OAI22xp5_ASAP7_75t_SL g238 ( 
.A1(n_201),
.A2(n_202),
.B1(n_209),
.B2(n_239),
.Y(n_238)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_202),
.Y(n_201)
);

BUFx2_ASAP7_75t_L g204 ( 
.A(n_205),
.Y(n_204)
);

INVx2_ASAP7_75t_L g205 ( 
.A(n_206),
.Y(n_205)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_207),
.Y(n_206)
);

INVx2_ASAP7_75t_L g207 ( 
.A(n_208),
.Y(n_207)
);

INVx3_ASAP7_75t_L g309 ( 
.A(n_208),
.Y(n_309)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_209),
.Y(n_239)
);

OAI22xp5_ASAP7_75t_L g211 ( 
.A1(n_212),
.A2(n_213),
.B1(n_219),
.B2(n_220),
.Y(n_211)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_212),
.Y(n_220)
);

MAJIxp5_ASAP7_75t_L g259 ( 
.A(n_212),
.B(n_260),
.C(n_261),
.Y(n_259)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_213),
.Y(n_219)
);

XNOR2xp5_ASAP7_75t_L g213 ( 
.A(n_214),
.B(n_215),
.Y(n_213)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_216),
.Y(n_218)
);

HB1xp67_ASAP7_75t_L g261 ( 
.A(n_219),
.Y(n_261)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_222),
.Y(n_221)
);

XNOR2x1_ASAP7_75t_L g222 ( 
.A(n_223),
.B(n_230),
.Y(n_222)
);

OAI22xp5_ASAP7_75t_SL g223 ( 
.A1(n_224),
.A2(n_225),
.B1(n_226),
.B2(n_227),
.Y(n_223)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_225),
.Y(n_224)
);

MAJIxp5_ASAP7_75t_L g258 ( 
.A(n_225),
.B(n_226),
.C(n_231),
.Y(n_258)
);

INVx1_ASAP7_75t_SL g226 ( 
.A(n_227),
.Y(n_226)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_231),
.Y(n_230)
);

MAJIxp5_ASAP7_75t_L g233 ( 
.A(n_234),
.B(n_237),
.C(n_240),
.Y(n_233)
);

XNOR2xp5_ASAP7_75t_L g367 ( 
.A(n_234),
.B(n_368),
.Y(n_367)
);

XOR2xp5_ASAP7_75t_L g368 ( 
.A(n_237),
.B(n_240),
.Y(n_368)
);

MAJIxp5_ASAP7_75t_L g240 ( 
.A(n_241),
.B(n_242),
.C(n_244),
.Y(n_240)
);

XOR2xp5_ASAP7_75t_L g363 ( 
.A(n_241),
.B(n_244),
.Y(n_363)
);

XNOR2xp5_ASAP7_75t_SL g362 ( 
.A(n_242),
.B(n_363),
.Y(n_362)
);

XOR2xp5_ASAP7_75t_L g342 ( 
.A(n_243),
.B(n_343),
.Y(n_342)
);

NAND2xp5_ASAP7_75t_SL g245 ( 
.A(n_246),
.B(n_282),
.Y(n_245)
);

INVx1_ASAP7_75t_L g369 ( 
.A(n_246),
.Y(n_369)
);

NAND2xp5_ASAP7_75t_L g246 ( 
.A(n_247),
.B(n_271),
.Y(n_246)
);

OR2x2_ASAP7_75t_L g375 ( 
.A(n_247),
.B(n_271),
.Y(n_375)
);

MAJIxp5_ASAP7_75t_L g247 ( 
.A(n_248),
.B(n_259),
.C(n_262),
.Y(n_247)
);

XOR2xp5_ASAP7_75t_L g284 ( 
.A(n_248),
.B(n_262),
.Y(n_284)
);

XNOR2xp5_ASAP7_75t_L g248 ( 
.A(n_249),
.B(n_258),
.Y(n_248)
);

OAI22xp5_ASAP7_75t_L g249 ( 
.A1(n_250),
.A2(n_251),
.B1(n_256),
.B2(n_257),
.Y(n_249)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_250),
.Y(n_256)
);

MAJIxp5_ASAP7_75t_L g272 ( 
.A(n_250),
.B(n_257),
.C(n_258),
.Y(n_272)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_251),
.Y(n_257)
);

OAI22xp5_ASAP7_75t_SL g251 ( 
.A1(n_252),
.A2(n_253),
.B1(n_254),
.B2(n_255),
.Y(n_251)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_253),
.Y(n_252)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_255),
.Y(n_254)
);

XNOR2xp5_ASAP7_75t_L g283 ( 
.A(n_259),
.B(n_284),
.Y(n_283)
);

XOR2x1_ASAP7_75t_L g262 ( 
.A(n_263),
.B(n_268),
.Y(n_262)
);

XOR2xp5_ASAP7_75t_L g263 ( 
.A(n_264),
.B(n_266),
.Y(n_263)
);

MAJIxp5_ASAP7_75t_L g281 ( 
.A(n_264),
.B(n_266),
.C(n_268),
.Y(n_281)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_269),
.Y(n_270)
);

XNOR2xp5_ASAP7_75t_L g271 ( 
.A(n_272),
.B(n_273),
.Y(n_271)
);

MAJIxp5_ASAP7_75t_R g378 ( 
.A(n_272),
.B(n_274),
.C(n_276),
.Y(n_378)
);

XOR2xp5_ASAP7_75t_L g273 ( 
.A(n_274),
.B(n_276),
.Y(n_273)
);

XNOR2xp5_ASAP7_75t_L g276 ( 
.A(n_277),
.B(n_281),
.Y(n_276)
);

XOR2xp5_ASAP7_75t_L g277 ( 
.A(n_278),
.B(n_280),
.Y(n_277)
);

MAJIxp5_ASAP7_75t_L g380 ( 
.A(n_278),
.B(n_280),
.C(n_281),
.Y(n_380)
);

NAND2xp5_ASAP7_75t_SL g282 ( 
.A(n_283),
.B(n_285),
.Y(n_282)
);

NOR2x1_ASAP7_75t_L g374 ( 
.A(n_283),
.B(n_285),
.Y(n_374)
);

NAND2xp5_ASAP7_75t_L g286 ( 
.A(n_287),
.B(n_365),
.Y(n_286)
);

OAI21xp5_ASAP7_75t_SL g287 ( 
.A1(n_288),
.A2(n_355),
.B(n_364),
.Y(n_287)
);

AOI21xp5_ASAP7_75t_L g288 ( 
.A1(n_289),
.A2(n_338),
.B(n_354),
.Y(n_288)
);

OAI21xp5_ASAP7_75t_SL g289 ( 
.A1(n_290),
.A2(n_319),
.B(n_337),
.Y(n_289)
);

NOR2xp33_ASAP7_75t_L g290 ( 
.A(n_291),
.B(n_303),
.Y(n_290)
);

NAND2xp5_ASAP7_75t_L g337 ( 
.A(n_291),
.B(n_303),
.Y(n_337)
);

MAJIxp5_ASAP7_75t_L g291 ( 
.A(n_292),
.B(n_296),
.C(n_300),
.Y(n_291)
);

XOR2xp5_ASAP7_75t_L g324 ( 
.A(n_292),
.B(n_325),
.Y(n_324)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_293),
.Y(n_295)
);

OAI22xp5_ASAP7_75t_SL g325 ( 
.A1(n_296),
.A2(n_300),
.B1(n_301),
.B2(n_326),
.Y(n_325)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_296),
.Y(n_326)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_297),
.Y(n_302)
);

INVx4_ASAP7_75t_L g298 ( 
.A(n_299),
.Y(n_298)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_301),
.Y(n_300)
);

XOR2xp5_ASAP7_75t_L g303 ( 
.A(n_304),
.B(n_312),
.Y(n_303)
);

MAJIxp5_ASAP7_75t_L g339 ( 
.A(n_304),
.B(n_313),
.C(n_318),
.Y(n_339)
);

XNOR2xp5_ASAP7_75t_L g304 ( 
.A(n_305),
.B(n_310),
.Y(n_304)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_306),
.Y(n_305)
);

AOI21xp5_ASAP7_75t_L g328 ( 
.A1(n_306),
.A2(n_329),
.B(n_331),
.Y(n_328)
);

INVxp67_ASAP7_75t_L g323 ( 
.A(n_307),
.Y(n_323)
);

BUFx3_ASAP7_75t_L g308 ( 
.A(n_309),
.Y(n_308)
);

OAI22xp5_ASAP7_75t_SL g312 ( 
.A1(n_313),
.A2(n_314),
.B1(n_317),
.B2(n_318),
.Y(n_312)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_314),
.Y(n_313)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_316),
.Y(n_315)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_318),
.Y(n_317)
);

AOI21xp5_ASAP7_75t_L g319 ( 
.A1(n_320),
.A2(n_327),
.B(n_336),
.Y(n_319)
);

NAND2xp5_ASAP7_75t_L g320 ( 
.A(n_321),
.B(n_324),
.Y(n_320)
);

NOR2xp33_ASAP7_75t_L g336 ( 
.A(n_321),
.B(n_324),
.Y(n_336)
);

XOR2xp5_ASAP7_75t_L g333 ( 
.A(n_322),
.B(n_334),
.Y(n_333)
);

NOR2xp33_ASAP7_75t_L g332 ( 
.A(n_326),
.B(n_333),
.Y(n_332)
);

NAND2xp5_ASAP7_75t_L g335 ( 
.A(n_326),
.B(n_333),
.Y(n_335)
);

OAI21xp5_ASAP7_75t_L g327 ( 
.A1(n_328),
.A2(n_332),
.B(n_335),
.Y(n_327)
);

NAND2xp5_ASAP7_75t_L g338 ( 
.A(n_339),
.B(n_340),
.Y(n_338)
);

NOR2xp33_ASAP7_75t_L g354 ( 
.A(n_339),
.B(n_340),
.Y(n_354)
);

XOR2x2_ASAP7_75t_L g340 ( 
.A(n_341),
.B(n_345),
.Y(n_340)
);

XOR2xp5_ASAP7_75t_L g341 ( 
.A(n_342),
.B(n_344),
.Y(n_341)
);

MAJIxp5_ASAP7_75t_L g356 ( 
.A(n_342),
.B(n_344),
.C(n_345),
.Y(n_356)
);

XNOR2xp5_ASAP7_75t_SL g345 ( 
.A(n_346),
.B(n_349),
.Y(n_345)
);

MAJIxp5_ASAP7_75t_L g359 ( 
.A(n_346),
.B(n_350),
.C(n_353),
.Y(n_359)
);

INVx1_ASAP7_75t_L g348 ( 
.A(n_347),
.Y(n_348)
);

OAI22xp5_ASAP7_75t_SL g349 ( 
.A1(n_350),
.A2(n_351),
.B1(n_352),
.B2(n_353),
.Y(n_349)
);

INVx1_ASAP7_75t_L g350 ( 
.A(n_351),
.Y(n_350)
);

INVx1_ASAP7_75t_L g352 ( 
.A(n_353),
.Y(n_352)
);

NOR2xp67_ASAP7_75t_SL g355 ( 
.A(n_356),
.B(n_357),
.Y(n_355)
);

NAND2xp5_ASAP7_75t_L g364 ( 
.A(n_356),
.B(n_357),
.Y(n_364)
);

XNOR2xp5_ASAP7_75t_L g357 ( 
.A(n_358),
.B(n_362),
.Y(n_357)
);

XOR2xp5_ASAP7_75t_L g358 ( 
.A(n_359),
.B(n_360),
.Y(n_358)
);

MAJIxp5_ASAP7_75t_L g366 ( 
.A(n_359),
.B(n_360),
.C(n_362),
.Y(n_366)
);

OR2x2_ASAP7_75t_L g365 ( 
.A(n_366),
.B(n_367),
.Y(n_365)
);

NAND2xp5_ASAP7_75t_L g373 ( 
.A(n_366),
.B(n_367),
.Y(n_373)
);

NAND2xp5_ASAP7_75t_SL g371 ( 
.A(n_372),
.B(n_373),
.Y(n_371)
);

CKINVDCx12_ASAP7_75t_R g376 ( 
.A(n_377),
.Y(n_376)
);

AND2x2_ASAP7_75t_L g377 ( 
.A(n_378),
.B(n_379),
.Y(n_377)
);

NOR2xp33_ASAP7_75t_L g393 ( 
.A(n_378),
.B(n_379),
.Y(n_393)
);

XNOR2xp5_ASAP7_75t_L g379 ( 
.A(n_380),
.B(n_381),
.Y(n_379)
);

MAJIxp5_ASAP7_75t_L g391 ( 
.A(n_380),
.B(n_382),
.C(n_384),
.Y(n_391)
);

XOR2xp5_ASAP7_75t_L g381 ( 
.A(n_382),
.B(n_384),
.Y(n_381)
);

INVx1_ASAP7_75t_L g387 ( 
.A(n_388),
.Y(n_387)
);

AOI21xp5_ASAP7_75t_SL g392 ( 
.A1(n_388),
.A2(n_393),
.B(n_394),
.Y(n_392)
);

NAND2xp5_ASAP7_75t_SL g388 ( 
.A(n_389),
.B(n_391),
.Y(n_388)
);

NOR2xp33_ASAP7_75t_L g394 ( 
.A(n_389),
.B(n_391),
.Y(n_394)
);


endmodule