module real_aes_16505_n_101 (n_17, n_28, n_76, n_56, n_34, n_98, n_90, n_82, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_83, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_91, n_100, n_43, n_96, n_54, n_35, n_42, n_99, n_15, n_9, n_23, n_72, n_95, n_44, n_7, n_4, n_80, n_6, n_12, n_68, n_79, n_69, n_46, n_59, n_25, n_73, n_77, n_81, n_48, n_37, n_97, n_70, n_50, n_89, n_26, n_86, n_93, n_13, n_24, n_2, n_55, n_62, n_84, n_67, n_92, n_33, n_88, n_14, n_11, n_85, n_16, n_94, n_39, n_5, n_45, n_60, n_38, n_87, n_0, n_78, n_63, n_1, n_53, n_36, n_101);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_98;
input n_90;
input n_82;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_83;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_91;
input n_100;
input n_43;
input n_96;
input n_54;
input n_35;
input n_42;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_95;
input n_44;
input n_7;
input n_4;
input n_80;
input n_6;
input n_12;
input n_68;
input n_79;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_81;
input n_48;
input n_37;
input n_97;
input n_70;
input n_50;
input n_89;
input n_26;
input n_86;
input n_93;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_84;
input n_67;
input n_92;
input n_33;
input n_88;
input n_14;
input n_11;
input n_85;
input n_16;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_87;
input n_0;
input n_78;
input n_63;
input n_1;
input n_53;
input n_36;
output n_101;
wire n_480;
wire n_113;
wire n_476;
wire n_758;
wire n_599;
wire n_187;
wire n_436;
wire n_684;
wire n_257;
wire n_390;
wire n_821;
wire n_830;
wire n_185;
wire n_285;
wire n_624;
wire n_618;
wire n_778;
wire n_800;
wire n_522;
wire n_838;
wire n_485;
wire n_822;
wire n_846;
wire n_222;
wire n_750;
wire n_631;
wire n_287;
wire n_357;
wire n_503;
wire n_635;
wire n_386;
wire n_673;
wire n_792;
wire n_518;
wire n_254;
wire n_207;
wire n_665;
wire n_667;
wire n_577;
wire n_580;
wire n_469;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_759;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_718;
wire n_318;
wire n_841;
wire n_355;
wire n_239;
wire n_669;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_761;
wire n_742;
wire n_112;
wire n_319;
wire n_364;
wire n_555;
wire n_421;
wire n_329;
wire n_766;
wire n_852;
wire n_132;
wire n_857;
wire n_131;
wire n_144;
wire n_461;
wire n_169;
wire n_242;
wire n_376;
wire n_549;
wire n_571;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_752;
wire n_448;
wire n_545;
wire n_556;
wire n_341;
wire n_593;
wire n_232;
wire n_460;
wire n_773;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_865;
wire n_537;
wire n_320;
wire n_666;
wire n_551;
wire n_560;
wire n_260;
wire n_660;
wire n_814;
wire n_594;
wire n_856;
wire n_186;
wire n_767;
wire n_138;
wire n_696;
wire n_704;
wire n_379;
wire n_374;
wire n_453;
wire n_647;
wire n_235;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_775;
wire n_161;
wire n_763;
wire n_189;
wire n_870;
wire n_271;
wire n_489;
wire n_548;
wire n_427;
wire n_678;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_564;
wire n_519;
wire n_815;
wire n_638;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_786;
wire n_512;
wire n_395;
wire n_332;
wire n_795;
wire n_816;
wire n_292;
wire n_539;
wire n_400;
wire n_626;
wire n_116;
wire n_625;
wire n_289;
wire n_462;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_818;
wire n_716;
wire n_213;
wire n_356;
wire n_478;
wire n_584;
wire n_408;
wire n_553;
wire n_184;
wire n_578;
wire n_372;
wire n_528;
wire n_202;
wire n_495;
wire n_370;
wire n_384;
wire n_744;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_824;
wire n_467;
wire n_327;
wire n_774;
wire n_813;
wire n_106;
wire n_791;
wire n_466;
wire n_559;
wire n_636;
wire n_872;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_726;
wire n_517;
wire n_683;
wire n_780;
wire n_174;
wire n_840;
wire n_570;
wire n_675;
wire n_530;
wire n_835;
wire n_104;
wire n_535;
wire n_732;
wire n_834;
wire n_784;
wire n_211;
wire n_281;
wire n_496;
wire n_693;
wire n_173;
wire n_468;
wire n_234;
wire n_755;
wire n_284;
wire n_153;
wire n_532;
wire n_316;
wire n_656;
wire n_746;
wire n_178;
wire n_409;
wire n_748;
wire n_781;
wire n_860;
wire n_298;
wire n_523;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_796;
wire n_297;
wire n_801;
wire n_383;
wire n_529;
wire n_119;
wire n_310;
wire n_455;
wire n_504;
wire n_725;
wire n_164;
wire n_671;
wire n_231;
wire n_102;
wire n_547;
wire n_659;
wire n_634;
wire n_682;
wire n_454;
wire n_122;
wire n_812;
wire n_817;
wire n_443;
wire n_565;
wire n_782;
wire n_760;
wire n_608;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_819;
wire n_267;
wire n_218;
wire n_737;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_828;
wire n_808;
wire n_770;
wire n_722;
wire n_745;
wire n_867;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_331;
wire n_182;
wire n_417;
wire n_363;
wire n_449;
wire n_607;
wire n_754;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_142;
wire n_561;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_783;
wire n_655;
wire n_654;
wire n_502;
wire n_434;
wire n_505;
wire n_527;
wire n_769;
wire n_600;
wire n_731;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_617;
wire n_552;
wire n_402;
wire n_602;
wire n_733;
wire n_171;
wire n_658;
wire n_676;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_146;
wire n_432;
wire n_807;
wire n_226;
wire n_255;
wire n_286;
wire n_416;
wire n_790;
wire n_832;
wire n_410;
wire n_120;
wire n_799;
wire n_805;
wire n_751;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_859;
wire n_695;
wire n_685;
wire n_165;
wire n_361;
wire n_632;
wire n_246;
wire n_176;
wire n_768;
wire n_412;
wire n_163;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_777;
wire n_488;
wire n_501;
wire n_251;
wire n_642;
wire n_613;
wire n_869;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_702;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_734;
wire n_110;
wire n_848;
wire n_392;
wire n_562;
wire n_150;
wire n_147;
wire n_288;
wire n_404;
wire n_598;
wire n_713;
wire n_735;
wire n_728;
wire n_756;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_569;
wire n_563;
wire n_785;
wire n_188;
wire n_269;
wire n_430;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_853;
wire n_810;
wire n_843;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_193;
wire n_397;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_649;
wire n_663;
wire n_749;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_707;
wire n_622;
wire n_470;
wire n_851;
wire n_133;
wire n_494;
wire n_711;
wire n_864;
wire n_377;
wire n_273;
wire n_723;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_845;
wire n_850;
wire n_265;
wire n_354;
wire n_720;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_730;
wire n_643;
wire n_747;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_847;
wire n_779;
wire n_148;
wire n_498;
wire n_481;
wire n_691;
wire n_765;
wire n_826;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_233;
wire n_487;
wire n_831;
wire n_290;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_155;
wire n_243;
wire n_692;
wire n_544;
wire n_268;
wire n_789;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_738;
wire n_701;
wire n_309;
wire n_344;
wire n_107;
wire n_229;
wire n_827;
wire n_809;
wire n_482;
wire n_520;
wire n_633;
wire n_679;
wire n_149;
wire n_472;
wire n_866;
wire n_452;
wire n_190;
wire n_787;
wire n_262;
wire n_630;
wire n_806;
wire n_689;
wire n_820;
wire n_715;
wire n_134;
wire n_349;
wire n_420;
wire n_336;
wire n_612;
wire n_858;
wire n_873;
wire n_195;
wire n_438;
wire n_764;
wire n_794;
wire n_300;
wire n_252;
wire n_283;
wire n_314;
wire n_741;
wire n_753;
wire n_249;
wire n_623;
wire n_446;
wire n_721;
wire n_221;
wire n_681;
wire n_156;
wire n_359;
wire n_456;
wire n_717;
wire n_312;
wire n_183;
wire n_266;
wire n_712;
wire n_205;
wire n_433;
wire n_335;
wire n_177;
wire n_516;
wire n_313;
wire n_627;
wire n_739;
wire n_140;
wire n_521;
wire n_418;
wire n_422;
wire n_771;
wire n_219;
wire n_524;
wire n_861;
wire n_705;
wire n_180;
wire n_212;
wire n_575;
wire n_210;
wire n_325;
wire n_762;
wire n_338;
wire n_479;
wire n_442;
wire n_825;
wire n_740;
wire n_371;
wire n_698;
wire n_103;
wire n_166;
wire n_541;
wire n_224;
wire n_839;
wire n_546;
wire n_151;
wire n_587;
wire n_639;
wire n_811;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_863;
wire n_724;
wire n_440;
wire n_525;
wire n_674;
wire n_644;
wire n_152;
wire n_198;
wire n_836;
wire n_793;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_833;
wire n_414;
wire n_757;
wire n_123;
wire n_279;
wire n_686;
wire n_776;
wire n_803;
wire n_543;
wire n_497;
wire n_514;
wire n_507;
wire n_270;
wire n_614;
wire n_305;
wire n_586;
wire n_772;
wire n_450;
wire n_788;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_465;
wire n_473;
wire n_719;
wire n_566;
wire n_837;
wire n_871;
wire n_474;
wire n_829;
wire n_170;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_168;
wire n_175;
wire n_241;
wire n_729;
wire n_687;
wire n_844;
wire n_646;
wire n_650;
wire n_710;
wire n_105;
wire n_743;
wire n_823;
wire n_294;
wire n_393;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_307;
wire n_500;
wire n_601;
wire n_661;
wire n_463;
wire n_396;
wire n_804;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_854;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_802;
wire n_868;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_842;
wire n_259;
wire n_143;
wire n_849;
wire n_192;
wire n_554;
wire n_475;
wire n_855;
wire n_264;
wire n_798;
wire n_237;
wire n_668;
wire n_797;
wire n_862;
AND2x4_ASAP7_75t_L g864 ( .A(n_0), .B(n_865), .Y(n_864) );
AOI22xp5_ASAP7_75t_L g248 ( .A1(n_1), .A2(n_5), .B1(n_249), .B2(n_250), .Y(n_248) );
INVx1_ASAP7_75t_L g872 ( .A(n_2), .Y(n_872) );
AOI22xp33_ASAP7_75t_L g545 ( .A1(n_3), .A2(n_45), .B1(n_120), .B2(n_149), .Y(n_545) );
AOI22xp33_ASAP7_75t_L g235 ( .A1(n_4), .A2(n_26), .B1(n_149), .B2(n_230), .Y(n_235) );
AOI22xp5_ASAP7_75t_L g592 ( .A1(n_6), .A2(n_17), .B1(n_510), .B2(n_593), .Y(n_592) );
AOI22xp5_ASAP7_75t_L g105 ( .A1(n_7), .A2(n_32), .B1(n_106), .B2(n_107), .Y(n_105) );
INVx1_ASAP7_75t_L g107 ( .A(n_7), .Y(n_107) );
AOI22xp33_ASAP7_75t_L g185 ( .A1(n_8), .A2(n_62), .B1(n_157), .B2(n_186), .Y(n_185) );
AOI22xp5_ASAP7_75t_L g119 ( .A1(n_9), .A2(n_18), .B1(n_120), .B2(n_122), .Y(n_119) );
INVx1_ASAP7_75t_L g865 ( .A(n_10), .Y(n_865) );
CKINVDCx5p33_ASAP7_75t_R g229 ( .A(n_11), .Y(n_229) );
CKINVDCx5p33_ASAP7_75t_R g563 ( .A(n_12), .Y(n_563) );
AOI22xp5_ASAP7_75t_L g530 ( .A1(n_13), .A2(n_20), .B1(n_531), .B2(n_532), .Y(n_530) );
OR2x2_ASAP7_75t_L g832 ( .A(n_14), .B(n_41), .Y(n_832) );
BUFx2_ASAP7_75t_L g870 ( .A(n_14), .Y(n_870) );
BUFx6f_ASAP7_75t_L g121 ( .A(n_15), .Y(n_121) );
CKINVDCx5p33_ASAP7_75t_R g595 ( .A(n_16), .Y(n_595) );
AOI21xp5_ASAP7_75t_L g847 ( .A1(n_19), .A2(n_848), .B(n_855), .Y(n_847) );
AOI22xp5_ASAP7_75t_L g509 ( .A1(n_21), .A2(n_99), .B1(n_250), .B2(n_510), .Y(n_509) );
AOI22xp33_ASAP7_75t_L g591 ( .A1(n_22), .A2(n_40), .B1(n_192), .B2(n_567), .Y(n_591) );
NAND2xp5_ASAP7_75t_SL g564 ( .A(n_23), .B(n_191), .Y(n_564) );
OAI21x1_ASAP7_75t_L g132 ( .A1(n_24), .A2(n_59), .B(n_133), .Y(n_132) );
CKINVDCx5p33_ASAP7_75t_R g239 ( .A(n_25), .Y(n_239) );
CKINVDCx5p33_ASAP7_75t_R g515 ( .A(n_27), .Y(n_515) );
NAND2xp5_ASAP7_75t_L g205 ( .A(n_28), .B(n_125), .Y(n_205) );
INVx4_ASAP7_75t_R g173 ( .A(n_29), .Y(n_173) );
AOI22xp33_ASAP7_75t_L g546 ( .A1(n_30), .A2(n_49), .B1(n_127), .B2(n_247), .Y(n_546) );
AOI22xp33_ASAP7_75t_L g520 ( .A1(n_31), .A2(n_55), .B1(n_127), .B2(n_510), .Y(n_520) );
INVx1_ASAP7_75t_L g106 ( .A(n_32), .Y(n_106) );
CKINVDCx5p33_ASAP7_75t_R g579 ( .A(n_33), .Y(n_579) );
NAND2xp5_ASAP7_75t_L g566 ( .A(n_34), .B(n_567), .Y(n_566) );
CKINVDCx5p33_ASAP7_75t_R g556 ( .A(n_35), .Y(n_556) );
NAND2xp5_ASAP7_75t_SL g212 ( .A(n_36), .B(n_149), .Y(n_212) );
INVx1_ASAP7_75t_L g254 ( .A(n_37), .Y(n_254) );
A2O1A1Ixp33_ASAP7_75t_SL g227 ( .A1(n_38), .A2(n_120), .B(n_124), .C(n_228), .Y(n_227) );
AOI22xp33_ASAP7_75t_L g236 ( .A1(n_39), .A2(n_56), .B1(n_120), .B2(n_127), .Y(n_236) );
HB1xp67_ASAP7_75t_L g868 ( .A(n_41), .Y(n_868) );
AOI22xp5_ASAP7_75t_L g575 ( .A1(n_42), .A2(n_87), .B1(n_120), .B2(n_576), .Y(n_575) );
CKINVDCx5p33_ASAP7_75t_R g225 ( .A(n_43), .Y(n_225) );
AOI22xp33_ASAP7_75t_L g533 ( .A1(n_44), .A2(n_48), .B1(n_120), .B2(n_122), .Y(n_533) );
OAI22xp5_ASAP7_75t_L g837 ( .A1(n_46), .A2(n_69), .B1(n_838), .B2(n_839), .Y(n_837) );
CKINVDCx5p33_ASAP7_75t_R g839 ( .A(n_46), .Y(n_839) );
AOI22xp33_ASAP7_75t_L g511 ( .A1(n_47), .A2(n_60), .B1(n_510), .B2(n_512), .Y(n_511) );
INVx1_ASAP7_75t_L g209 ( .A(n_50), .Y(n_209) );
NAND2xp5_ASAP7_75t_L g211 ( .A(n_51), .B(n_120), .Y(n_211) );
CKINVDCx5p33_ASAP7_75t_R g147 ( .A(n_52), .Y(n_147) );
INVx2_ASAP7_75t_L g827 ( .A(n_53), .Y(n_827) );
BUFx3_ASAP7_75t_L g830 ( .A(n_54), .Y(n_830) );
INVx1_ASAP7_75t_L g846 ( .A(n_54), .Y(n_846) );
CKINVDCx5p33_ASAP7_75t_R g175 ( .A(n_57), .Y(n_175) );
AOI22xp33_ASAP7_75t_L g126 ( .A1(n_58), .A2(n_88), .B1(n_120), .B2(n_127), .Y(n_126) );
CKINVDCx20_ASAP7_75t_R g857 ( .A(n_61), .Y(n_857) );
AOI22xp33_ASAP7_75t_L g519 ( .A1(n_63), .A2(n_76), .B1(n_247), .B2(n_512), .Y(n_519) );
CKINVDCx5p33_ASAP7_75t_R g138 ( .A(n_64), .Y(n_138) );
AOI22xp33_ASAP7_75t_L g554 ( .A1(n_65), .A2(n_79), .B1(n_120), .B2(n_122), .Y(n_554) );
AOI22xp5_ASAP7_75t_L g553 ( .A1(n_66), .A2(n_97), .B1(n_510), .B2(n_532), .Y(n_553) );
INVx1_ASAP7_75t_L g133 ( .A(n_67), .Y(n_133) );
AND2x4_ASAP7_75t_L g135 ( .A(n_68), .B(n_136), .Y(n_135) );
INVx1_ASAP7_75t_L g838 ( .A(n_69), .Y(n_838) );
AOI22xp33_ASAP7_75t_L g246 ( .A1(n_70), .A2(n_90), .B1(n_127), .B2(n_247), .Y(n_246) );
AO22x1_ASAP7_75t_L g189 ( .A1(n_71), .A2(n_77), .B1(n_190), .B2(n_192), .Y(n_189) );
INVx1_ASAP7_75t_L g136 ( .A(n_72), .Y(n_136) );
AND2x2_ASAP7_75t_L g231 ( .A(n_73), .B(n_143), .Y(n_231) );
NAND2xp5_ASAP7_75t_L g156 ( .A(n_74), .B(n_157), .Y(n_156) );
CKINVDCx5p33_ASAP7_75t_R g222 ( .A(n_75), .Y(n_222) );
NAND2xp5_ASAP7_75t_L g148 ( .A(n_78), .B(n_149), .Y(n_148) );
INVx2_ASAP7_75t_L g125 ( .A(n_80), .Y(n_125) );
CKINVDCx5p33_ASAP7_75t_R g170 ( .A(n_81), .Y(n_170) );
NAND2xp5_ASAP7_75t_L g202 ( .A(n_82), .B(n_143), .Y(n_202) );
AOI22xp33_ASAP7_75t_L g577 ( .A1(n_83), .A2(n_98), .B1(n_127), .B2(n_157), .Y(n_577) );
CKINVDCx5p33_ASAP7_75t_R g522 ( .A(n_84), .Y(n_522) );
NAND2xp5_ASAP7_75t_L g187 ( .A(n_85), .B(n_131), .Y(n_187) );
CKINVDCx5p33_ASAP7_75t_R g548 ( .A(n_86), .Y(n_548) );
NAND2xp5_ASAP7_75t_SL g570 ( .A(n_89), .B(n_143), .Y(n_570) );
CKINVDCx5p33_ASAP7_75t_R g536 ( .A(n_91), .Y(n_536) );
NAND2xp5_ASAP7_75t_SL g142 ( .A(n_92), .B(n_143), .Y(n_142) );
INVx1_ASAP7_75t_L g497 ( .A(n_93), .Y(n_497) );
NOR2xp33_ASAP7_75t_L g844 ( .A(n_93), .B(n_845), .Y(n_844) );
NAND2xp33_ASAP7_75t_L g568 ( .A(n_94), .B(n_191), .Y(n_568) );
A2O1A1Ixp33_ASAP7_75t_L g167 ( .A1(n_95), .A2(n_129), .B(n_157), .C(n_168), .Y(n_167) );
AND2x2_ASAP7_75t_L g177 ( .A(n_96), .B(n_178), .Y(n_177) );
NAND2xp33_ASAP7_75t_L g154 ( .A(n_100), .B(n_155), .Y(n_154) );
AOI21xp33_ASAP7_75t_L g101 ( .A1(n_102), .A2(n_858), .B(n_871), .Y(n_101) );
AO21x2_ASAP7_75t_L g102 ( .A1(n_103), .A2(n_823), .B(n_833), .Y(n_102) );
OAI22xp5_ASAP7_75t_L g103 ( .A1(n_104), .A2(n_105), .B1(n_108), .B2(n_822), .Y(n_103) );
INVx1_ASAP7_75t_L g104 ( .A(n_105), .Y(n_104) );
INVx2_ASAP7_75t_L g822 ( .A(n_108), .Y(n_822) );
OAI22x1_ASAP7_75t_L g108 ( .A1(n_109), .A2(n_494), .B1(n_498), .B2(n_819), .Y(n_108) );
AND2x2_ASAP7_75t_L g109 ( .A(n_110), .B(n_403), .Y(n_109) );
NOR3xp33_ASAP7_75t_L g110 ( .A(n_111), .B(n_319), .C(n_350), .Y(n_110) );
NAND2xp5_ASAP7_75t_L g111 ( .A(n_112), .B(n_285), .Y(n_111) );
AOI211x1_ASAP7_75t_SL g112 ( .A1(n_113), .A2(n_197), .B(n_240), .C(n_271), .Y(n_112) );
INVx1_ASAP7_75t_L g113 ( .A(n_114), .Y(n_113) );
NAND2xp5_ASAP7_75t_L g114 ( .A(n_115), .B(n_161), .Y(n_114) );
AND2x2_ASAP7_75t_L g426 ( .A(n_115), .B(n_301), .Y(n_426) );
AND2x2_ASAP7_75t_L g115 ( .A(n_116), .B(n_140), .Y(n_115) );
INVx1_ASAP7_75t_L g311 ( .A(n_116), .Y(n_311) );
OR2x2_ASAP7_75t_L g432 ( .A(n_116), .B(n_283), .Y(n_432) );
INVx2_ASAP7_75t_L g116 ( .A(n_117), .Y(n_116) );
AND2x2_ASAP7_75t_L g268 ( .A(n_117), .B(n_141), .Y(n_268) );
NAND2xp5_ASAP7_75t_L g282 ( .A(n_117), .B(n_283), .Y(n_282) );
INVx2_ASAP7_75t_L g300 ( .A(n_117), .Y(n_300) );
OR2x2_ASAP7_75t_L g331 ( .A(n_117), .B(n_162), .Y(n_331) );
AND2x2_ASAP7_75t_L g345 ( .A(n_117), .B(n_162), .Y(n_345) );
AND2x2_ASAP7_75t_L g382 ( .A(n_117), .B(n_338), .Y(n_382) );
AO31x2_ASAP7_75t_L g117 ( .A1(n_118), .A2(n_130), .A3(n_134), .B(n_137), .Y(n_117) );
OAI22x1_ASAP7_75t_L g118 ( .A1(n_119), .A2(n_123), .B1(n_126), .B2(n_128), .Y(n_118) );
INVx4_ASAP7_75t_L g122 ( .A(n_120), .Y(n_122) );
INVx1_ASAP7_75t_L g512 ( .A(n_120), .Y(n_512) );
INVx1_ASAP7_75t_L g532 ( .A(n_120), .Y(n_532) );
INVx3_ASAP7_75t_L g120 ( .A(n_121), .Y(n_120) );
BUFx6f_ASAP7_75t_L g127 ( .A(n_121), .Y(n_127) );
BUFx6f_ASAP7_75t_L g149 ( .A(n_121), .Y(n_149) );
BUFx6f_ASAP7_75t_L g155 ( .A(n_121), .Y(n_155) );
INVx1_ASAP7_75t_L g157 ( .A(n_121), .Y(n_157) );
INVx1_ASAP7_75t_L g169 ( .A(n_121), .Y(n_169) );
INVx1_ASAP7_75t_L g174 ( .A(n_121), .Y(n_174) );
BUFx6f_ASAP7_75t_L g191 ( .A(n_121), .Y(n_191) );
INVx1_ASAP7_75t_L g193 ( .A(n_121), .Y(n_193) );
INVx1_ASAP7_75t_L g224 ( .A(n_121), .Y(n_224) );
INVx2_ASAP7_75t_L g230 ( .A(n_121), .Y(n_230) );
O2A1O1Ixp33_ASAP7_75t_L g146 ( .A1(n_122), .A2(n_147), .B(n_148), .C(n_150), .Y(n_146) );
O2A1O1Ixp5_ASAP7_75t_L g562 ( .A1(n_122), .A2(n_124), .B(n_563), .C(n_564), .Y(n_562) );
OAI22xp5_ASAP7_75t_L g234 ( .A1(n_123), .A2(n_183), .B1(n_235), .B2(n_236), .Y(n_234) );
OAI22xp5_ASAP7_75t_L g245 ( .A1(n_123), .A2(n_128), .B1(n_246), .B2(n_248), .Y(n_245) );
OAI22xp5_ASAP7_75t_L g508 ( .A1(n_123), .A2(n_509), .B1(n_511), .B2(n_513), .Y(n_508) );
OAI22xp5_ASAP7_75t_L g518 ( .A1(n_123), .A2(n_513), .B1(n_519), .B2(n_520), .Y(n_518) );
OAI22xp5_ASAP7_75t_L g529 ( .A1(n_123), .A2(n_530), .B1(n_533), .B2(n_534), .Y(n_529) );
OAI22xp5_ASAP7_75t_L g544 ( .A1(n_123), .A2(n_513), .B1(n_545), .B2(n_546), .Y(n_544) );
OAI22xp5_ASAP7_75t_L g552 ( .A1(n_123), .A2(n_534), .B1(n_553), .B2(n_554), .Y(n_552) );
AOI21xp5_ASAP7_75t_L g565 ( .A1(n_123), .A2(n_566), .B(n_568), .Y(n_565) );
OAI22xp5_ASAP7_75t_L g574 ( .A1(n_123), .A2(n_128), .B1(n_575), .B2(n_577), .Y(n_574) );
OAI22xp5_ASAP7_75t_L g590 ( .A1(n_123), .A2(n_513), .B1(n_591), .B2(n_592), .Y(n_590) );
INVx6_ASAP7_75t_L g123 ( .A(n_124), .Y(n_123) );
AOI21xp5_ASAP7_75t_L g153 ( .A1(n_124), .A2(n_154), .B(n_156), .Y(n_153) );
NAND2xp5_ASAP7_75t_L g188 ( .A(n_124), .B(n_189), .Y(n_188) );
A2O1A1Ixp33_ASAP7_75t_L g284 ( .A1(n_124), .A2(n_182), .B(n_189), .C(n_195), .Y(n_284) );
BUFx8_ASAP7_75t_L g124 ( .A(n_125), .Y(n_124) );
INVx1_ASAP7_75t_L g129 ( .A(n_125), .Y(n_129) );
INVx2_ASAP7_75t_L g152 ( .A(n_125), .Y(n_152) );
INVx1_ASAP7_75t_L g208 ( .A(n_125), .Y(n_208) );
NAND2xp5_ASAP7_75t_L g206 ( .A(n_127), .B(n_207), .Y(n_206) );
INVx2_ASAP7_75t_L g249 ( .A(n_127), .Y(n_249) );
NAND2xp5_ASAP7_75t_SL g171 ( .A(n_128), .B(n_172), .Y(n_171) );
INVx1_ASAP7_75t_L g128 ( .A(n_129), .Y(n_128) );
INVx1_ASAP7_75t_SL g534 ( .A(n_129), .Y(n_534) );
NOR2xp33_ASAP7_75t_L g514 ( .A(n_130), .B(n_515), .Y(n_514) );
NOR2xp33_ASAP7_75t_L g521 ( .A(n_130), .B(n_522), .Y(n_521) );
INVx2_ASAP7_75t_L g130 ( .A(n_131), .Y(n_130) );
INVx2_ASAP7_75t_L g139 ( .A(n_131), .Y(n_139) );
INVx2_ASAP7_75t_L g165 ( .A(n_131), .Y(n_165) );
OAI21xp33_ASAP7_75t_L g195 ( .A1(n_131), .A2(n_187), .B(n_196), .Y(n_195) );
INVx2_ASAP7_75t_L g131 ( .A(n_132), .Y(n_131) );
BUFx6f_ASAP7_75t_L g144 ( .A(n_132), .Y(n_144) );
INVx2_ASAP7_75t_L g176 ( .A(n_134), .Y(n_176) );
AO31x2_ASAP7_75t_L g528 ( .A1(n_134), .A2(n_218), .A3(n_529), .B(n_535), .Y(n_528) );
AO31x2_ASAP7_75t_L g543 ( .A1(n_134), .A2(n_237), .A3(n_544), .B(n_547), .Y(n_543) );
AO31x2_ASAP7_75t_L g589 ( .A1(n_134), .A2(n_573), .A3(n_590), .B(n_594), .Y(n_589) );
BUFx10_ASAP7_75t_L g134 ( .A(n_135), .Y(n_134) );
BUFx10_ASAP7_75t_L g160 ( .A(n_135), .Y(n_160) );
INVx1_ASAP7_75t_L g196 ( .A(n_135), .Y(n_196) );
INVx1_ASAP7_75t_L g252 ( .A(n_135), .Y(n_252) );
NOR2xp33_ASAP7_75t_L g137 ( .A(n_138), .B(n_139), .Y(n_137) );
INVx2_ASAP7_75t_L g178 ( .A(n_139), .Y(n_178) );
BUFx2_ASAP7_75t_L g218 ( .A(n_139), .Y(n_218) );
NOR2xp33_ASAP7_75t_L g238 ( .A(n_139), .B(n_239), .Y(n_238) );
NOR2xp33_ASAP7_75t_L g253 ( .A(n_139), .B(n_254), .Y(n_253) );
BUFx2_ASAP7_75t_L g262 ( .A(n_140), .Y(n_262) );
AND2x2_ASAP7_75t_L g313 ( .A(n_140), .B(n_179), .Y(n_313) );
AND2x2_ASAP7_75t_L g456 ( .A(n_140), .B(n_162), .Y(n_456) );
INVx2_ASAP7_75t_L g140 ( .A(n_141), .Y(n_140) );
BUFx3_ASAP7_75t_L g280 ( .A(n_141), .Y(n_280) );
AND2x2_ASAP7_75t_L g299 ( .A(n_141), .B(n_300), .Y(n_299) );
INVx1_ASAP7_75t_L g336 ( .A(n_141), .Y(n_336) );
AND2x2_ASAP7_75t_L g360 ( .A(n_141), .B(n_162), .Y(n_360) );
NAND2x1p5_ASAP7_75t_L g141 ( .A(n_142), .B(n_145), .Y(n_141) );
NOR2x1_ASAP7_75t_L g158 ( .A(n_143), .B(n_159), .Y(n_158) );
INVx2_ASAP7_75t_L g237 ( .A(n_143), .Y(n_237) );
INVx4_ASAP7_75t_L g143 ( .A(n_144), .Y(n_143) );
AND2x2_ASAP7_75t_L g213 ( .A(n_144), .B(n_160), .Y(n_213) );
NOR2xp33_ASAP7_75t_L g547 ( .A(n_144), .B(n_548), .Y(n_547) );
NOR2xp33_ASAP7_75t_L g555 ( .A(n_144), .B(n_556), .Y(n_555) );
INVx2_ASAP7_75t_SL g560 ( .A(n_144), .Y(n_560) );
BUFx3_ASAP7_75t_L g573 ( .A(n_144), .Y(n_573) );
NOR2xp33_ASAP7_75t_L g594 ( .A(n_144), .B(n_595), .Y(n_594) );
OAI21x1_ASAP7_75t_L g145 ( .A1(n_146), .A2(n_153), .B(n_158), .Y(n_145) );
NOR2xp33_ASAP7_75t_L g221 ( .A(n_149), .B(n_222), .Y(n_221) );
INVx2_ASAP7_75t_SL g150 ( .A(n_151), .Y(n_150) );
INVx2_ASAP7_75t_L g151 ( .A(n_152), .Y(n_151) );
BUFx3_ASAP7_75t_L g184 ( .A(n_152), .Y(n_184) );
OAI22xp33_ASAP7_75t_L g172 ( .A1(n_155), .A2(n_173), .B1(n_174), .B2(n_175), .Y(n_172) );
INVx2_ASAP7_75t_L g247 ( .A(n_155), .Y(n_247) );
INVx1_ASAP7_75t_L g567 ( .A(n_155), .Y(n_567) );
INVx1_ASAP7_75t_L g159 ( .A(n_160), .Y(n_159) );
AO31x2_ASAP7_75t_L g233 ( .A1(n_160), .A2(n_234), .A3(n_237), .B(n_238), .Y(n_233) );
HB1xp67_ASAP7_75t_L g260 ( .A(n_161), .Y(n_260) );
AND2x2_ASAP7_75t_L g321 ( .A(n_161), .B(n_310), .Y(n_321) );
INVx2_ASAP7_75t_L g453 ( .A(n_161), .Y(n_453) );
AND2x2_ASAP7_75t_L g161 ( .A(n_162), .B(n_179), .Y(n_161) );
INVx1_ASAP7_75t_L g258 ( .A(n_162), .Y(n_258) );
AND2x4_ASAP7_75t_L g270 ( .A(n_162), .B(n_180), .Y(n_270) );
INVx2_ASAP7_75t_L g338 ( .A(n_162), .Y(n_338) );
AO21x2_ASAP7_75t_L g162 ( .A1(n_163), .A2(n_166), .B(n_177), .Y(n_162) );
AO31x2_ASAP7_75t_L g506 ( .A1(n_163), .A2(n_507), .A3(n_508), .B(n_514), .Y(n_506) );
AO31x2_ASAP7_75t_L g517 ( .A1(n_163), .A2(n_251), .A3(n_518), .B(n_521), .Y(n_517) );
INVx2_ASAP7_75t_L g163 ( .A(n_164), .Y(n_163) );
INVx2_ASAP7_75t_L g164 ( .A(n_165), .Y(n_164) );
NOR2xp33_ASAP7_75t_SL g535 ( .A(n_165), .B(n_536), .Y(n_535) );
NOR2xp33_ASAP7_75t_L g578 ( .A(n_165), .B(n_579), .Y(n_578) );
AOI21xp5_ASAP7_75t_L g166 ( .A1(n_167), .A2(n_171), .B(n_176), .Y(n_166) );
NOR2xp33_ASAP7_75t_L g168 ( .A(n_169), .B(n_170), .Y(n_168) );
INVx2_ASAP7_75t_L g186 ( .A(n_169), .Y(n_186) );
INVx1_ASAP7_75t_L g593 ( .A(n_174), .Y(n_593) );
INVx1_ASAP7_75t_L g507 ( .A(n_176), .Y(n_507) );
AND2x2_ASAP7_75t_L g337 ( .A(n_179), .B(n_338), .Y(n_337) );
INVx1_ASAP7_75t_L g344 ( .A(n_179), .Y(n_344) );
INVx2_ASAP7_75t_L g179 ( .A(n_180), .Y(n_179) );
AND2x2_ASAP7_75t_L g422 ( .A(n_180), .B(n_338), .Y(n_422) );
AOI21x1_ASAP7_75t_L g180 ( .A1(n_181), .A2(n_188), .B(n_194), .Y(n_180) );
INVx1_ASAP7_75t_L g181 ( .A(n_182), .Y(n_181) );
OAI21x1_ASAP7_75t_L g182 ( .A1(n_183), .A2(n_185), .B(n_187), .Y(n_182) );
AOI21xp5_ASAP7_75t_L g210 ( .A1(n_183), .A2(n_211), .B(n_212), .Y(n_210) );
INVx2_ASAP7_75t_L g183 ( .A(n_184), .Y(n_183) );
INVx2_ASAP7_75t_L g513 ( .A(n_184), .Y(n_513) );
INVx1_ASAP7_75t_L g531 ( .A(n_186), .Y(n_531) );
INVxp67_ASAP7_75t_SL g190 ( .A(n_191), .Y(n_190) );
INVx3_ASAP7_75t_L g510 ( .A(n_191), .Y(n_510) );
OAI21xp33_ASAP7_75t_SL g204 ( .A1(n_192), .A2(n_205), .B(n_206), .Y(n_204) );
INVx1_ASAP7_75t_L g192 ( .A(n_193), .Y(n_192) );
INVx1_ASAP7_75t_L g194 ( .A(n_195), .Y(n_194) );
AOI21xp5_ASAP7_75t_L g219 ( .A1(n_196), .A2(n_220), .B(n_227), .Y(n_219) );
INVx1_ASAP7_75t_L g197 ( .A(n_198), .Y(n_197) );
NAND2xp5_ASAP7_75t_L g198 ( .A(n_199), .B(n_214), .Y(n_198) );
OR2x2_ASAP7_75t_L g327 ( .A(n_199), .B(n_215), .Y(n_327) );
AND2x2_ASAP7_75t_L g465 ( .A(n_199), .B(n_409), .Y(n_465) );
INVx2_ASAP7_75t_L g199 ( .A(n_200), .Y(n_199) );
AND2x4_ASAP7_75t_L g242 ( .A(n_200), .B(n_243), .Y(n_242) );
OR2x2_ASAP7_75t_L g347 ( .A(n_200), .B(n_348), .Y(n_347) );
NAND2xp5_ASAP7_75t_L g389 ( .A(n_200), .B(n_289), .Y(n_389) );
NAND2xp5_ASAP7_75t_L g402 ( .A(n_200), .B(n_265), .Y(n_402) );
INVx3_ASAP7_75t_L g200 ( .A(n_201), .Y(n_200) );
INVx1_ASAP7_75t_L g259 ( .A(n_201), .Y(n_259) );
AND2x2_ASAP7_75t_L g275 ( .A(n_201), .B(n_276), .Y(n_275) );
NAND2x1p5_ASAP7_75t_SL g288 ( .A(n_201), .B(n_289), .Y(n_288) );
OR2x2_ASAP7_75t_L g296 ( .A(n_201), .B(n_297), .Y(n_296) );
NAND2xp5_ASAP7_75t_L g367 ( .A(n_201), .B(n_265), .Y(n_367) );
AND2x2_ASAP7_75t_L g415 ( .A(n_201), .B(n_244), .Y(n_415) );
NAND2xp5_ASAP7_75t_L g458 ( .A(n_201), .B(n_243), .Y(n_458) );
BUFx2_ASAP7_75t_L g477 ( .A(n_201), .Y(n_477) );
AND2x4_ASAP7_75t_L g201 ( .A(n_202), .B(n_203), .Y(n_201) );
OAI21xp5_ASAP7_75t_L g203 ( .A1(n_204), .A2(n_210), .B(n_213), .Y(n_203) );
NOR2xp33_ASAP7_75t_L g207 ( .A(n_208), .B(n_209), .Y(n_207) );
BUFx4f_ASAP7_75t_L g226 ( .A(n_208), .Y(n_226) );
INVx1_ASAP7_75t_L g214 ( .A(n_215), .Y(n_214) );
OR2x2_ASAP7_75t_L g261 ( .A(n_215), .B(n_262), .Y(n_261) );
INVx2_ASAP7_75t_L g374 ( .A(n_215), .Y(n_374) );
OR2x2_ASAP7_75t_L g215 ( .A(n_216), .B(n_232), .Y(n_215) );
NOR2xp33_ASAP7_75t_L g277 ( .A(n_216), .B(n_244), .Y(n_277) );
INVx2_ASAP7_75t_L g289 ( .A(n_216), .Y(n_289) );
AND2x2_ASAP7_75t_L g325 ( .A(n_216), .B(n_233), .Y(n_325) );
INVx2_ASAP7_75t_L g216 ( .A(n_217), .Y(n_216) );
INVx1_ASAP7_75t_L g265 ( .A(n_217), .Y(n_265) );
AOI21x1_ASAP7_75t_L g217 ( .A1(n_218), .A2(n_219), .B(n_231), .Y(n_217) );
AO31x2_ASAP7_75t_L g244 ( .A1(n_218), .A2(n_245), .A3(n_251), .B(n_253), .Y(n_244) );
AO31x2_ASAP7_75t_L g551 ( .A1(n_218), .A2(n_507), .A3(n_552), .B(n_555), .Y(n_551) );
OAI21xp5_ASAP7_75t_L g220 ( .A1(n_221), .A2(n_223), .B(n_226), .Y(n_220) );
NOR2xp33_ASAP7_75t_L g223 ( .A(n_224), .B(n_225), .Y(n_223) );
INVx2_ASAP7_75t_L g250 ( .A(n_224), .Y(n_250) );
NOR2xp33_ASAP7_75t_L g228 ( .A(n_229), .B(n_230), .Y(n_228) );
INVx2_ASAP7_75t_SL g576 ( .A(n_230), .Y(n_576) );
INVx1_ASAP7_75t_L g349 ( .A(n_232), .Y(n_349) );
NAND2xp5_ASAP7_75t_L g366 ( .A(n_232), .B(n_244), .Y(n_366) );
INVx2_ASAP7_75t_SL g232 ( .A(n_233), .Y(n_232) );
BUFx2_ASAP7_75t_L g276 ( .A(n_233), .Y(n_276) );
OR2x2_ASAP7_75t_L g308 ( .A(n_233), .B(n_244), .Y(n_308) );
NAND2xp5_ASAP7_75t_L g386 ( .A(n_233), .B(n_244), .Y(n_386) );
OAI22xp5_ASAP7_75t_L g240 ( .A1(n_241), .A2(n_261), .B1(n_263), .B2(n_267), .Y(n_240) );
AOI22xp5_ASAP7_75t_L g241 ( .A1(n_242), .A2(n_255), .B1(n_259), .B2(n_260), .Y(n_241) );
INVx2_ASAP7_75t_L g266 ( .A(n_242), .Y(n_266) );
NAND2xp5_ASAP7_75t_L g339 ( .A(n_242), .B(n_325), .Y(n_339) );
AND2x2_ASAP7_75t_L g373 ( .A(n_242), .B(n_374), .Y(n_373) );
INVx1_ASAP7_75t_L g243 ( .A(n_244), .Y(n_243) );
INVx1_ASAP7_75t_L g291 ( .A(n_244), .Y(n_291) );
INVx1_ASAP7_75t_L g297 ( .A(n_244), .Y(n_297) );
AO31x2_ASAP7_75t_L g572 ( .A1(n_251), .A2(n_573), .A3(n_574), .B(n_578), .Y(n_572) );
INVx2_ASAP7_75t_SL g251 ( .A(n_252), .Y(n_251) );
INVx2_ASAP7_75t_SL g569 ( .A(n_252), .Y(n_569) );
INVx1_ASAP7_75t_L g255 ( .A(n_256), .Y(n_255) );
INVx1_ASAP7_75t_L g256 ( .A(n_257), .Y(n_256) );
OR2x2_ASAP7_75t_L g431 ( .A(n_257), .B(n_432), .Y(n_431) );
INVx1_ASAP7_75t_L g257 ( .A(n_258), .Y(n_257) );
INVx1_ASAP7_75t_L g312 ( .A(n_258), .Y(n_312) );
AND3x1_ASAP7_75t_L g416 ( .A(n_258), .B(n_279), .C(n_417), .Y(n_416) );
INVx1_ASAP7_75t_L g372 ( .A(n_259), .Y(n_372) );
AND2x4_ASAP7_75t_L g408 ( .A(n_259), .B(n_409), .Y(n_408) );
INVx1_ASAP7_75t_L g446 ( .A(n_262), .Y(n_446) );
INVx1_ASAP7_75t_L g450 ( .A(n_263), .Y(n_450) );
OR2x2_ASAP7_75t_L g263 ( .A(n_264), .B(n_266), .Y(n_263) );
OR2x2_ASAP7_75t_L g423 ( .A(n_264), .B(n_424), .Y(n_423) );
INVxp67_ASAP7_75t_SL g471 ( .A(n_264), .Y(n_471) );
INVxp67_ASAP7_75t_L g264 ( .A(n_265), .Y(n_264) );
OR2x2_ASAP7_75t_L g371 ( .A(n_265), .B(n_349), .Y(n_371) );
AND2x2_ASAP7_75t_L g413 ( .A(n_265), .B(n_280), .Y(n_413) );
HB1xp67_ASAP7_75t_L g417 ( .A(n_265), .Y(n_417) );
NAND2xp5_ASAP7_75t_SL g267 ( .A(n_268), .B(n_269), .Y(n_267) );
O2A1O1Ixp33_ASAP7_75t_L g332 ( .A1(n_268), .A2(n_269), .B(n_333), .C(n_339), .Y(n_332) );
NAND2x1_ASAP7_75t_L g376 ( .A(n_268), .B(n_377), .Y(n_376) );
NOR2xp33_ASAP7_75t_L g472 ( .A(n_268), .B(n_426), .Y(n_472) );
INVx3_ASAP7_75t_L g269 ( .A(n_270), .Y(n_269) );
NAND2xp5_ASAP7_75t_L g318 ( .A(n_270), .B(n_299), .Y(n_318) );
INVx1_ASAP7_75t_L g271 ( .A(n_272), .Y(n_271) );
NAND2xp5_ASAP7_75t_SL g272 ( .A(n_273), .B(n_278), .Y(n_272) );
INVx2_ASAP7_75t_L g273 ( .A(n_274), .Y(n_273) );
NAND2xp5_ASAP7_75t_L g274 ( .A(n_275), .B(n_277), .Y(n_274) );
INVx2_ASAP7_75t_L g294 ( .A(n_276), .Y(n_294) );
HB1xp67_ASAP7_75t_L g355 ( .A(n_277), .Y(n_355) );
NOR2xp33_ASAP7_75t_L g419 ( .A(n_278), .B(n_420), .Y(n_419) );
AND2x2_ASAP7_75t_L g278 ( .A(n_279), .B(n_281), .Y(n_278) );
AND2x2_ASAP7_75t_L g328 ( .A(n_279), .B(n_329), .Y(n_328) );
NAND2xp5_ASAP7_75t_L g392 ( .A(n_279), .B(n_345), .Y(n_392) );
NAND2x1p5_ASAP7_75t_L g398 ( .A(n_279), .B(n_399), .Y(n_398) );
NAND2xp5_ASAP7_75t_L g493 ( .A(n_279), .B(n_337), .Y(n_493) );
INVx3_ASAP7_75t_L g279 ( .A(n_280), .Y(n_279) );
BUFx2_ASAP7_75t_L g476 ( .A(n_280), .Y(n_476) );
INVx1_ASAP7_75t_L g281 ( .A(n_282), .Y(n_281) );
INVx2_ASAP7_75t_L g302 ( .A(n_283), .Y(n_302) );
INVx1_ASAP7_75t_L g283 ( .A(n_284), .Y(n_283) );
AOI21xp5_ASAP7_75t_L g285 ( .A1(n_286), .A2(n_298), .B(n_303), .Y(n_285) );
NAND2xp5_ASAP7_75t_L g286 ( .A(n_287), .B(n_292), .Y(n_286) );
OR2x2_ASAP7_75t_L g287 ( .A(n_288), .B(n_290), .Y(n_287) );
OAI33xp33_ASAP7_75t_L g352 ( .A1(n_288), .A2(n_293), .A3(n_353), .B1(n_354), .B2(n_356), .B3(n_357), .Y(n_352) );
OR2x2_ASAP7_75t_L g484 ( .A(n_288), .B(n_308), .Y(n_484) );
INVx2_ASAP7_75t_L g486 ( .A(n_288), .Y(n_486) );
INVx1_ASAP7_75t_L g307 ( .A(n_289), .Y(n_307) );
OR2x2_ASAP7_75t_L g348 ( .A(n_289), .B(n_349), .Y(n_348) );
INVx1_ASAP7_75t_L g290 ( .A(n_291), .Y(n_290) );
NAND2xp5_ASAP7_75t_L g292 ( .A(n_293), .B(n_295), .Y(n_292) );
INVx1_ASAP7_75t_L g356 ( .A(n_293), .Y(n_356) );
NOR3xp33_ASAP7_75t_L g474 ( .A(n_293), .B(n_475), .C(n_477), .Y(n_474) );
INVx2_ASAP7_75t_L g293 ( .A(n_294), .Y(n_293) );
NOR2xp33_ASAP7_75t_L g433 ( .A(n_294), .B(n_434), .Y(n_433) );
NOR2xp33_ASAP7_75t_L g462 ( .A(n_294), .B(n_458), .Y(n_462) );
AND2x4_ASAP7_75t_L g491 ( .A(n_294), .B(n_492), .Y(n_491) );
INVxp67_ASAP7_75t_SL g295 ( .A(n_296), .Y(n_295) );
INVx1_ASAP7_75t_L g317 ( .A(n_296), .Y(n_317) );
OR2x2_ASAP7_75t_L g323 ( .A(n_296), .B(n_324), .Y(n_323) );
OR2x2_ASAP7_75t_L g436 ( .A(n_296), .B(n_371), .Y(n_436) );
INVx1_ASAP7_75t_L g492 ( .A(n_296), .Y(n_492) );
AND2x4_ASAP7_75t_SL g298 ( .A(n_299), .B(n_301), .Y(n_298) );
INVx1_ASAP7_75t_L g315 ( .A(n_299), .Y(n_315) );
INVx1_ASAP7_75t_L g358 ( .A(n_300), .Y(n_358) );
AND2x2_ASAP7_75t_L g399 ( .A(n_300), .B(n_302), .Y(n_399) );
INVx1_ASAP7_75t_L g439 ( .A(n_301), .Y(n_439) );
INVx2_ASAP7_75t_L g301 ( .A(n_302), .Y(n_301) );
OR2x2_ASAP7_75t_L g330 ( .A(n_302), .B(n_331), .Y(n_330) );
OAI22xp33_ASAP7_75t_L g303 ( .A1(n_304), .A2(n_309), .B1(n_316), .B2(n_318), .Y(n_303) );
INVx2_ASAP7_75t_L g304 ( .A(n_305), .Y(n_304) );
INVx2_ASAP7_75t_L g305 ( .A(n_306), .Y(n_305) );
OR2x2_ASAP7_75t_L g306 ( .A(n_307), .B(n_308), .Y(n_306) );
INVx2_ASAP7_75t_L g395 ( .A(n_308), .Y(n_395) );
INVx2_ASAP7_75t_L g409 ( .A(n_308), .Y(n_409) );
AOI211xp5_ASAP7_75t_L g309 ( .A1(n_310), .A2(n_312), .B(n_313), .C(n_314), .Y(n_309) );
INVx1_ASAP7_75t_L g353 ( .A(n_310), .Y(n_353) );
INVx1_ASAP7_75t_L g310 ( .A(n_311), .Y(n_310) );
NAND2xp5_ASAP7_75t_L g438 ( .A(n_311), .B(n_336), .Y(n_438) );
OR2x2_ASAP7_75t_L g454 ( .A(n_311), .B(n_455), .Y(n_454) );
INVx1_ASAP7_75t_L g467 ( .A(n_311), .Y(n_467) );
NAND2xp5_ASAP7_75t_L g442 ( .A(n_313), .B(n_381), .Y(n_442) );
INVx1_ASAP7_75t_L g314 ( .A(n_315), .Y(n_314) );
INVx1_ASAP7_75t_L g316 ( .A(n_317), .Y(n_316) );
NAND2xp5_ASAP7_75t_SL g319 ( .A(n_320), .B(n_340), .Y(n_319) );
AOI221xp5_ASAP7_75t_L g320 ( .A1(n_321), .A2(n_322), .B1(n_326), .B2(n_328), .C(n_332), .Y(n_320) );
INVx2_ASAP7_75t_L g322 ( .A(n_323), .Y(n_322) );
OAI32xp33_ASAP7_75t_L g489 ( .A1(n_323), .A2(n_420), .A3(n_438), .B1(n_490), .B2(n_493), .Y(n_489) );
INVx1_ASAP7_75t_L g324 ( .A(n_325), .Y(n_324) );
INVx1_ASAP7_75t_L g459 ( .A(n_325), .Y(n_459) );
INVx2_ASAP7_75t_L g326 ( .A(n_327), .Y(n_326) );
OAI21xp5_ASAP7_75t_L g340 ( .A1(n_328), .A2(n_341), .B(n_346), .Y(n_340) );
NAND2x1_ASAP7_75t_L g488 ( .A(n_329), .B(n_476), .Y(n_488) );
INVx2_ASAP7_75t_L g329 ( .A(n_330), .Y(n_329) );
INVx2_ASAP7_75t_L g363 ( .A(n_331), .Y(n_363) );
INVx1_ASAP7_75t_L g333 ( .A(n_334), .Y(n_333) );
AND2x2_ASAP7_75t_L g334 ( .A(n_335), .B(n_337), .Y(n_334) );
AND2x2_ASAP7_75t_L g482 ( .A(n_335), .B(n_363), .Y(n_482) );
INVx2_ASAP7_75t_L g335 ( .A(n_336), .Y(n_335) );
INVx1_ASAP7_75t_L g430 ( .A(n_336), .Y(n_430) );
INVx2_ASAP7_75t_L g383 ( .A(n_337), .Y(n_383) );
INVx2_ASAP7_75t_SL g341 ( .A(n_342), .Y(n_341) );
NAND2xp5_ASAP7_75t_L g342 ( .A(n_343), .B(n_345), .Y(n_342) );
AND2x2_ASAP7_75t_L g359 ( .A(n_343), .B(n_360), .Y(n_359) );
INVx1_ASAP7_75t_L g343 ( .A(n_344), .Y(n_343) );
INVx2_ASAP7_75t_L g378 ( .A(n_344), .Y(n_378) );
INVx1_ASAP7_75t_L g346 ( .A(n_347), .Y(n_346) );
NAND4xp25_ASAP7_75t_L g350 ( .A(n_351), .B(n_368), .C(n_379), .D(n_390), .Y(n_350) );
AOI22xp5_ASAP7_75t_L g351 ( .A1(n_352), .A2(n_359), .B1(n_361), .B2(n_364), .Y(n_351) );
OAI22xp5_ASAP7_75t_L g480 ( .A1(n_353), .A2(n_481), .B1(n_483), .B2(n_484), .Y(n_480) );
INVx1_ASAP7_75t_L g354 ( .A(n_355), .Y(n_354) );
INVx1_ASAP7_75t_L g357 ( .A(n_358), .Y(n_357) );
AND2x2_ASAP7_75t_L g463 ( .A(n_358), .B(n_422), .Y(n_463) );
AND2x2_ASAP7_75t_L g466 ( .A(n_360), .B(n_467), .Y(n_466) );
AOI22xp5_ASAP7_75t_L g379 ( .A1(n_361), .A2(n_380), .B1(n_384), .B2(n_387), .Y(n_379) );
INVx1_ASAP7_75t_L g361 ( .A(n_362), .Y(n_361) );
INVx1_ASAP7_75t_L g362 ( .A(n_363), .Y(n_362) );
INVx2_ASAP7_75t_L g364 ( .A(n_365), .Y(n_364) );
OR2x2_ASAP7_75t_L g365 ( .A(n_366), .B(n_367), .Y(n_365) );
OR2x2_ASAP7_75t_L g401 ( .A(n_366), .B(n_402), .Y(n_401) );
OR2x2_ASAP7_75t_L g385 ( .A(n_367), .B(n_386), .Y(n_385) );
INVx1_ASAP7_75t_L g396 ( .A(n_367), .Y(n_396) );
OAI21xp5_ASAP7_75t_L g368 ( .A1(n_369), .A2(n_373), .B(n_375), .Y(n_368) );
O2A1O1Ixp33_ASAP7_75t_L g473 ( .A1(n_369), .A2(n_474), .B(n_478), .C(n_480), .Y(n_473) );
AND2x2_ASAP7_75t_L g369 ( .A(n_370), .B(n_372), .Y(n_369) );
INVxp67_ASAP7_75t_L g370 ( .A(n_371), .Y(n_370) );
INVx1_ASAP7_75t_L g448 ( .A(n_371), .Y(n_448) );
AND2x4_ASAP7_75t_L g441 ( .A(n_374), .B(n_415), .Y(n_441) );
INVx2_ASAP7_75t_SL g375 ( .A(n_376), .Y(n_375) );
INVx1_ASAP7_75t_L g377 ( .A(n_378), .Y(n_377) );
NAND2xp5_ASAP7_75t_L g380 ( .A(n_381), .B(n_383), .Y(n_380) );
OAI21xp33_ASAP7_75t_L g406 ( .A1(n_381), .A2(n_407), .B(n_410), .Y(n_406) );
INVx2_ASAP7_75t_L g381 ( .A(n_382), .Y(n_381) );
AND2x2_ASAP7_75t_L g412 ( .A(n_382), .B(n_413), .Y(n_412) );
NAND2xp5_ASAP7_75t_L g445 ( .A(n_382), .B(n_446), .Y(n_445) );
INVx2_ASAP7_75t_L g384 ( .A(n_385), .Y(n_384) );
OR2x2_ASAP7_75t_L g388 ( .A(n_386), .B(n_389), .Y(n_388) );
INVx1_ASAP7_75t_L g387 ( .A(n_388), .Y(n_387) );
OAI22xp5_ASAP7_75t_L g418 ( .A1(n_388), .A2(n_419), .B1(n_423), .B2(n_425), .Y(n_418) );
AOI22xp33_ASAP7_75t_L g390 ( .A1(n_391), .A2(n_393), .B1(n_397), .B2(n_400), .Y(n_390) );
INVx1_ASAP7_75t_L g391 ( .A(n_392), .Y(n_391) );
INVx1_ASAP7_75t_L g393 ( .A(n_394), .Y(n_393) );
NAND2xp5_ASAP7_75t_L g394 ( .A(n_395), .B(n_396), .Y(n_394) );
HB1xp67_ASAP7_75t_L g411 ( .A(n_395), .Y(n_411) );
INVx1_ASAP7_75t_L g397 ( .A(n_398), .Y(n_397) );
INVx1_ASAP7_75t_L g400 ( .A(n_401), .Y(n_400) );
NOR2xp33_ASAP7_75t_L g403 ( .A(n_404), .B(n_468), .Y(n_403) );
NAND4xp25_ASAP7_75t_L g404 ( .A(n_405), .B(n_427), .C(n_443), .D(n_460), .Y(n_404) );
NOR2xp33_ASAP7_75t_L g405 ( .A(n_406), .B(n_418), .Y(n_405) );
INVx2_ASAP7_75t_L g407 ( .A(n_408), .Y(n_407) );
AND2x2_ASAP7_75t_L g470 ( .A(n_408), .B(n_471), .Y(n_470) );
AOI22xp5_ASAP7_75t_L g410 ( .A1(n_411), .A2(n_412), .B1(n_414), .B2(n_416), .Y(n_410) );
INVxp67_ASAP7_75t_L g434 ( .A(n_414), .Y(n_434) );
BUFx2_ASAP7_75t_SL g414 ( .A(n_415), .Y(n_414) );
INVx1_ASAP7_75t_L g424 ( .A(n_415), .Y(n_424) );
AND2x2_ASAP7_75t_L g447 ( .A(n_415), .B(n_448), .Y(n_447) );
INVx3_ASAP7_75t_L g420 ( .A(n_421), .Y(n_420) );
INVx2_ASAP7_75t_L g421 ( .A(n_422), .Y(n_421) );
INVx1_ASAP7_75t_L g425 ( .A(n_426), .Y(n_425) );
AOI21xp5_ASAP7_75t_L g427 ( .A1(n_428), .A2(n_433), .B(n_435), .Y(n_427) );
NOR2x1_ASAP7_75t_L g428 ( .A(n_429), .B(n_431), .Y(n_428) );
INVx1_ASAP7_75t_L g429 ( .A(n_430), .Y(n_429) );
OR2x6_ASAP7_75t_L g452 ( .A(n_430), .B(n_453), .Y(n_452) );
INVx3_ASAP7_75t_L g449 ( .A(n_431), .Y(n_449) );
OAI32xp33_ASAP7_75t_L g435 ( .A1(n_436), .A2(n_437), .A3(n_439), .B1(n_440), .B2(n_442), .Y(n_435) );
INVx2_ASAP7_75t_L g437 ( .A(n_438), .Y(n_437) );
INVx1_ASAP7_75t_L g440 ( .A(n_441), .Y(n_440) );
AOI221xp5_ASAP7_75t_L g443 ( .A1(n_444), .A2(n_447), .B1(n_449), .B2(n_450), .C(n_451), .Y(n_443) );
INVx1_ASAP7_75t_L g444 ( .A(n_445), .Y(n_444) );
AOI21xp5_ASAP7_75t_L g451 ( .A1(n_452), .A2(n_454), .B(n_457), .Y(n_451) );
INVx2_ASAP7_75t_SL g455 ( .A(n_456), .Y(n_455) );
OR2x2_ASAP7_75t_L g457 ( .A(n_458), .B(n_459), .Y(n_457) );
NOR2x1_ASAP7_75t_L g460 ( .A(n_461), .B(n_464), .Y(n_460) );
AND2x2_ASAP7_75t_L g461 ( .A(n_462), .B(n_463), .Y(n_461) );
INVx1_ASAP7_75t_L g483 ( .A(n_462), .Y(n_483) );
INVx1_ASAP7_75t_L g479 ( .A(n_463), .Y(n_479) );
AND2x2_ASAP7_75t_L g464 ( .A(n_465), .B(n_466), .Y(n_464) );
OAI211xp5_ASAP7_75t_SL g468 ( .A1(n_469), .A2(n_472), .B(n_473), .C(n_485), .Y(n_468) );
INVx1_ASAP7_75t_L g469 ( .A(n_470), .Y(n_469) );
INVx1_ASAP7_75t_L g475 ( .A(n_476), .Y(n_475) );
INVxp67_ASAP7_75t_L g478 ( .A(n_479), .Y(n_478) );
INVx1_ASAP7_75t_SL g481 ( .A(n_482), .Y(n_481) );
AOI21xp33_ASAP7_75t_L g485 ( .A1(n_486), .A2(n_487), .B(n_489), .Y(n_485) );
INVx2_ASAP7_75t_L g487 ( .A(n_488), .Y(n_487) );
INVx2_ASAP7_75t_L g490 ( .A(n_491), .Y(n_490) );
CKINVDCx5p33_ASAP7_75t_R g494 ( .A(n_495), .Y(n_494) );
BUFx8_ASAP7_75t_SL g495 ( .A(n_496), .Y(n_495) );
AND2x2_ASAP7_75t_L g853 ( .A(n_496), .B(n_854), .Y(n_853) );
INVx2_ASAP7_75t_L g496 ( .A(n_497), .Y(n_496) );
BUFx2_ASAP7_75t_L g821 ( .A(n_497), .Y(n_821) );
XNOR2x1_ASAP7_75t_L g836 ( .A(n_498), .B(n_837), .Y(n_836) );
AND3x4_ASAP7_75t_L g498 ( .A(n_499), .B(n_681), .C(n_735), .Y(n_498) );
NOR2x1_ASAP7_75t_L g499 ( .A(n_500), .B(n_641), .Y(n_499) );
NAND3xp33_ASAP7_75t_L g500 ( .A(n_501), .B(n_580), .C(n_623), .Y(n_500) );
OAI21xp33_ASAP7_75t_L g501 ( .A1(n_502), .A2(n_523), .B(n_538), .Y(n_501) );
INVx1_ASAP7_75t_L g502 ( .A(n_503), .Y(n_502) );
HB1xp67_ASAP7_75t_L g503 ( .A(n_504), .Y(n_503) );
OR2x2_ASAP7_75t_L g673 ( .A(n_504), .B(n_584), .Y(n_673) );
INVx2_ASAP7_75t_L g699 ( .A(n_504), .Y(n_699) );
OR2x2_ASAP7_75t_L g504 ( .A(n_505), .B(n_516), .Y(n_504) );
INVx1_ASAP7_75t_L g598 ( .A(n_505), .Y(n_598) );
INVx2_ASAP7_75t_L g713 ( .A(n_505), .Y(n_713) );
INVx2_ASAP7_75t_L g505 ( .A(n_506), .Y(n_505) );
INVx2_ASAP7_75t_L g526 ( .A(n_506), .Y(n_526) );
AND2x4_ASAP7_75t_L g656 ( .A(n_506), .B(n_618), .Y(n_656) );
INVx1_ASAP7_75t_L g709 ( .A(n_516), .Y(n_709) );
INVx2_ASAP7_75t_L g516 ( .A(n_517), .Y(n_516) );
INVx1_ASAP7_75t_L g537 ( .A(n_517), .Y(n_537) );
AND2x4_ASAP7_75t_L g587 ( .A(n_517), .B(n_588), .Y(n_587) );
HB1xp67_ASAP7_75t_L g615 ( .A(n_517), .Y(n_615) );
INVx2_ASAP7_75t_L g618 ( .A(n_517), .Y(n_618) );
OR2x2_ASAP7_75t_L g632 ( .A(n_517), .B(n_589), .Y(n_632) );
AND2x2_ASAP7_75t_L g734 ( .A(n_517), .B(n_528), .Y(n_734) );
INVx1_ASAP7_75t_L g523 ( .A(n_524), .Y(n_523) );
NAND2xp5_ASAP7_75t_SL g789 ( .A(n_524), .B(n_790), .Y(n_789) );
OR2x2_ASAP7_75t_L g524 ( .A(n_525), .B(n_527), .Y(n_524) );
OR2x2_ASAP7_75t_L g616 ( .A(n_525), .B(n_617), .Y(n_616) );
NAND2xp5_ASAP7_75t_SL g680 ( .A(n_525), .B(n_635), .Y(n_680) );
AND2x2_ASAP7_75t_L g745 ( .A(n_525), .B(n_721), .Y(n_745) );
INVx4_ASAP7_75t_L g779 ( .A(n_525), .Y(n_779) );
INVx3_ASAP7_75t_L g525 ( .A(n_526), .Y(n_525) );
AND2x2_ASAP7_75t_L g614 ( .A(n_526), .B(n_615), .Y(n_614) );
AND2x2_ASAP7_75t_L g652 ( .A(n_526), .B(n_586), .Y(n_652) );
AND2x2_ASAP7_75t_L g762 ( .A(n_526), .B(n_589), .Y(n_762) );
AND2x2_ASAP7_75t_L g796 ( .A(n_526), .B(n_618), .Y(n_796) );
NAND2xp5_ASAP7_75t_L g527 ( .A(n_528), .B(n_537), .Y(n_527) );
INVx4_ASAP7_75t_SL g586 ( .A(n_528), .Y(n_586) );
NAND2xp5_ASAP7_75t_L g611 ( .A(n_528), .B(n_612), .Y(n_611) );
AND2x2_ASAP7_75t_L g697 ( .A(n_528), .B(n_589), .Y(n_697) );
BUFx2_ASAP7_75t_L g715 ( .A(n_528), .Y(n_715) );
AOI222xp33_ASAP7_75t_L g623 ( .A1(n_537), .A2(n_624), .B1(n_629), .B2(n_630), .C1(n_633), .C2(n_637), .Y(n_623) );
INVx1_ASAP7_75t_L g754 ( .A(n_537), .Y(n_754) );
AND2x2_ASAP7_75t_L g538 ( .A(n_539), .B(n_549), .Y(n_538) );
AND2x2_ASAP7_75t_L g791 ( .A(n_539), .B(n_603), .Y(n_791) );
INVx1_ASAP7_75t_L g539 ( .A(n_540), .Y(n_539) );
AND2x2_ASAP7_75t_L g812 ( .A(n_540), .B(n_813), .Y(n_812) );
INVx1_ASAP7_75t_L g540 ( .A(n_541), .Y(n_540) );
AND2x4_ASAP7_75t_L g621 ( .A(n_541), .B(n_622), .Y(n_621) );
NAND2xp5_ASAP7_75t_L g760 ( .A(n_541), .B(n_604), .Y(n_760) );
INVx2_ASAP7_75t_L g541 ( .A(n_542), .Y(n_541) );
NAND2xp5_ASAP7_75t_L g650 ( .A(n_542), .B(n_608), .Y(n_650) );
AND2x2_ASAP7_75t_L g678 ( .A(n_542), .B(n_558), .Y(n_678) );
INVx2_ASAP7_75t_L g542 ( .A(n_543), .Y(n_542) );
AND2x2_ASAP7_75t_L g607 ( .A(n_543), .B(n_608), .Y(n_607) );
OR2x2_ASAP7_75t_L g640 ( .A(n_543), .B(n_572), .Y(n_640) );
INVx1_ASAP7_75t_L g668 ( .A(n_543), .Y(n_668) );
HB1xp67_ASAP7_75t_L g774 ( .A(n_543), .Y(n_774) );
AOI222xp33_ASAP7_75t_L g723 ( .A1(n_549), .A2(n_666), .B1(n_724), .B2(n_725), .C1(n_727), .C2(n_729), .Y(n_723) );
AND2x4_ASAP7_75t_L g549 ( .A(n_550), .B(n_557), .Y(n_549) );
INVx1_ASAP7_75t_L g658 ( .A(n_550), .Y(n_658) );
BUFx2_ASAP7_75t_L g550 ( .A(n_551), .Y(n_550) );
INVx3_ASAP7_75t_L g604 ( .A(n_551), .Y(n_604) );
AND2x2_ASAP7_75t_L g609 ( .A(n_551), .B(n_572), .Y(n_609) );
AND2x2_ASAP7_75t_L g669 ( .A(n_551), .B(n_571), .Y(n_669) );
AND2x2_ASAP7_75t_L g657 ( .A(n_557), .B(n_658), .Y(n_657) );
AND2x4_ASAP7_75t_L g752 ( .A(n_557), .B(n_668), .Y(n_752) );
NAND2xp5_ASAP7_75t_L g758 ( .A(n_557), .B(n_759), .Y(n_758) );
AND3x1_ASAP7_75t_L g817 ( .A(n_557), .B(n_587), .C(n_818), .Y(n_817) );
AND2x4_ASAP7_75t_L g557 ( .A(n_558), .B(n_571), .Y(n_557) );
AND2x2_ASAP7_75t_L g638 ( .A(n_558), .B(n_604), .Y(n_638) );
NAND2xp5_ASAP7_75t_L g787 ( .A(n_558), .B(n_740), .Y(n_787) );
INVx2_ASAP7_75t_L g558 ( .A(n_559), .Y(n_558) );
BUFx2_ASAP7_75t_L g601 ( .A(n_559), .Y(n_601) );
OAI21x1_ASAP7_75t_L g559 ( .A1(n_560), .A2(n_561), .B(n_570), .Y(n_559) );
OAI21x1_ASAP7_75t_L g608 ( .A1(n_560), .A2(n_561), .B(n_570), .Y(n_608) );
OAI21x1_ASAP7_75t_L g561 ( .A1(n_562), .A2(n_565), .B(n_569), .Y(n_561) );
INVx2_ASAP7_75t_L g571 ( .A(n_572), .Y(n_571) );
AND2x4_ASAP7_75t_L g603 ( .A(n_572), .B(n_604), .Y(n_603) );
OR2x2_ASAP7_75t_L g636 ( .A(n_572), .B(n_622), .Y(n_636) );
INVx1_ASAP7_75t_L g646 ( .A(n_572), .Y(n_646) );
BUFx2_ASAP7_75t_L g740 ( .A(n_572), .Y(n_740) );
AOI21xp5_ASAP7_75t_L g580 ( .A1(n_581), .A2(n_599), .B(n_605), .Y(n_580) );
INVx1_ASAP7_75t_L g581 ( .A(n_582), .Y(n_581) );
NAND2x1_ASAP7_75t_L g582 ( .A(n_583), .B(n_596), .Y(n_582) );
AOI221xp5_ASAP7_75t_SL g663 ( .A1(n_583), .A2(n_664), .B1(n_670), .B2(n_674), .C(n_679), .Y(n_663) );
AND2x4_ASAP7_75t_L g583 ( .A(n_584), .B(n_587), .Y(n_583) );
INVx2_ASAP7_75t_L g584 ( .A(n_585), .Y(n_584) );
NAND2xp5_ASAP7_75t_L g784 ( .A(n_585), .B(n_598), .Y(n_784) );
INVx2_ASAP7_75t_L g585 ( .A(n_586), .Y(n_585) );
NAND2xp5_ASAP7_75t_L g617 ( .A(n_586), .B(n_618), .Y(n_617) );
AND2x4_ASAP7_75t_L g626 ( .A(n_586), .B(n_627), .Y(n_626) );
INVx1_ASAP7_75t_L g662 ( .A(n_586), .Y(n_662) );
INVx1_ASAP7_75t_L g672 ( .A(n_586), .Y(n_672) );
AND2x2_ASAP7_75t_L g691 ( .A(n_586), .B(n_692), .Y(n_691) );
OR2x2_ASAP7_75t_L g703 ( .A(n_586), .B(n_704), .Y(n_703) );
NAND2xp5_ASAP7_75t_L g816 ( .A(n_586), .B(n_709), .Y(n_816) );
INVx2_ASAP7_75t_L g651 ( .A(n_587), .Y(n_651) );
AND2x2_ASAP7_75t_L g661 ( .A(n_587), .B(n_662), .Y(n_661) );
NAND2xp5_ASAP7_75t_L g671 ( .A(n_587), .B(n_672), .Y(n_671) );
NAND2xp5_ASAP7_75t_L g804 ( .A(n_587), .B(n_805), .Y(n_804) );
INVx2_ASAP7_75t_L g588 ( .A(n_589), .Y(n_588) );
INVx1_ASAP7_75t_L g612 ( .A(n_589), .Y(n_612) );
HB1xp67_ASAP7_75t_L g655 ( .A(n_589), .Y(n_655) );
INVx1_ASAP7_75t_L g692 ( .A(n_589), .Y(n_692) );
NAND2xp5_ASAP7_75t_L g708 ( .A(n_589), .B(n_709), .Y(n_708) );
INVx1_ASAP7_75t_L g596 ( .A(n_597), .Y(n_596) );
OR2x2_ASAP7_75t_L g631 ( .A(n_597), .B(n_632), .Y(n_631) );
NAND2xp5_ASAP7_75t_L g733 ( .A(n_597), .B(n_734), .Y(n_733) );
INVx1_ASAP7_75t_L g597 ( .A(n_598), .Y(n_597) );
HB1xp67_ASAP7_75t_L g690 ( .A(n_598), .Y(n_690) );
NOR2xp33_ASAP7_75t_R g599 ( .A(n_600), .B(n_602), .Y(n_599) );
INVx1_ASAP7_75t_L g600 ( .A(n_601), .Y(n_600) );
NOR3xp33_ASAP7_75t_L g679 ( .A(n_601), .B(n_671), .C(n_680), .Y(n_679) );
AND2x2_ASAP7_75t_L g702 ( .A(n_601), .B(n_609), .Y(n_702) );
AND2x2_ASAP7_75t_L g731 ( .A(n_601), .B(n_701), .Y(n_731) );
OR2x2_ASAP7_75t_L g798 ( .A(n_601), .B(n_799), .Y(n_798) );
INVx1_ASAP7_75t_L g602 ( .A(n_603), .Y(n_602) );
AND2x4_ASAP7_75t_L g724 ( .A(n_603), .B(n_607), .Y(n_724) );
INVx2_ASAP7_75t_SL g808 ( .A(n_603), .Y(n_808) );
INVx2_ASAP7_75t_L g635 ( .A(n_604), .Y(n_635) );
NAND2xp5_ASAP7_75t_L g648 ( .A(n_604), .B(n_649), .Y(n_648) );
INVx3_ASAP7_75t_L g677 ( .A(n_604), .Y(n_677) );
HB1xp67_ASAP7_75t_L g750 ( .A(n_604), .Y(n_750) );
OAI32xp33_ASAP7_75t_L g605 ( .A1(n_606), .A2(n_610), .A3(n_613), .B1(n_616), .B2(n_619), .Y(n_605) );
NAND2xp5_ASAP7_75t_L g606 ( .A(n_607), .B(n_609), .Y(n_606) );
AND2x2_ASAP7_75t_L g629 ( .A(n_607), .B(n_609), .Y(n_629) );
AND2x2_ASAP7_75t_L g687 ( .A(n_607), .B(n_669), .Y(n_687) );
NAND2xp5_ASAP7_75t_L g695 ( .A(n_607), .B(n_669), .Y(n_695) );
INVx1_ASAP7_75t_L g622 ( .A(n_608), .Y(n_622) );
AND2x4_ASAP7_75t_SL g620 ( .A(n_609), .B(n_621), .Y(n_620) );
INVx1_ASAP7_75t_SL g764 ( .A(n_609), .Y(n_764) );
INVx2_ASAP7_75t_L g799 ( .A(n_609), .Y(n_799) );
AND2x2_ASAP7_75t_L g811 ( .A(n_609), .B(n_678), .Y(n_811) );
NOR3xp33_ASAP7_75t_L g741 ( .A(n_610), .B(n_732), .C(n_742), .Y(n_741) );
INVx1_ASAP7_75t_L g610 ( .A(n_611), .Y(n_610) );
INVx1_ASAP7_75t_L g627 ( .A(n_612), .Y(n_627) );
AOI321xp33_ASAP7_75t_L g810 ( .A1(n_613), .A2(n_672), .A3(n_811), .B1(n_812), .B2(n_814), .C(n_817), .Y(n_810) );
INVx2_ASAP7_75t_L g613 ( .A(n_614), .Y(n_613) );
INVx1_ASAP7_75t_L g628 ( .A(n_615), .Y(n_628) );
OAI22xp5_ASAP7_75t_L g814 ( .A1(n_617), .A2(n_636), .B1(n_815), .B2(n_816), .Y(n_814) );
INVx3_ASAP7_75t_L g619 ( .A(n_620), .Y(n_619) );
AND2x2_ASAP7_75t_L g717 ( .A(n_621), .B(n_676), .Y(n_717) );
INVx1_ASAP7_75t_L g624 ( .A(n_625), .Y(n_624) );
NAND2xp5_ASAP7_75t_SL g625 ( .A(n_626), .B(n_628), .Y(n_625) );
INVx1_ASAP7_75t_L g751 ( .A(n_626), .Y(n_751) );
NAND2x1_ASAP7_75t_L g778 ( .A(n_626), .B(n_779), .Y(n_778) );
NAND2xp5_ASAP7_75t_L g795 ( .A(n_626), .B(n_796), .Y(n_795) );
AND2x2_ASAP7_75t_L g776 ( .A(n_628), .B(n_762), .Y(n_776) );
INVx2_ASAP7_75t_L g630 ( .A(n_631), .Y(n_630) );
INVx2_ASAP7_75t_L g716 ( .A(n_632), .Y(n_716) );
OR2x2_ASAP7_75t_L g783 ( .A(n_632), .B(n_784), .Y(n_783) );
INVx1_ASAP7_75t_L g633 ( .A(n_634), .Y(n_633) );
OR2x2_ASAP7_75t_L g634 ( .A(n_635), .B(n_636), .Y(n_634) );
NOR2xp33_ASAP7_75t_L g660 ( .A(n_635), .B(n_636), .Y(n_660) );
NOR2x1p5_ASAP7_75t_L g701 ( .A(n_635), .B(n_640), .Y(n_701) );
INVx1_ASAP7_75t_L g771 ( .A(n_635), .Y(n_771) );
NOR2x1_ASAP7_75t_L g772 ( .A(n_636), .B(n_773), .Y(n_772) );
AND2x2_ASAP7_75t_L g637 ( .A(n_638), .B(n_639), .Y(n_637) );
INVxp67_ASAP7_75t_SL g815 ( .A(n_638), .Y(n_815) );
INVx1_ASAP7_75t_L g639 ( .A(n_640), .Y(n_639) );
NAND3xp33_ASAP7_75t_L g641 ( .A(n_642), .B(n_653), .C(n_663), .Y(n_641) );
NAND3xp33_ASAP7_75t_L g642 ( .A(n_643), .B(n_651), .C(n_652), .Y(n_642) );
AND2x4_ASAP7_75t_L g643 ( .A(n_644), .B(n_647), .Y(n_643) );
INVx1_ASAP7_75t_L g644 ( .A(n_645), .Y(n_644) );
BUFx2_ASAP7_75t_L g645 ( .A(n_646), .Y(n_645) );
INVx1_ASAP7_75t_L g793 ( .A(n_647), .Y(n_793) );
INVx1_ASAP7_75t_L g647 ( .A(n_648), .Y(n_647) );
INVxp67_ASAP7_75t_SL g649 ( .A(n_650), .Y(n_649) );
INVx1_ASAP7_75t_L g685 ( .A(n_650), .Y(n_685) );
INVx1_ASAP7_75t_L g721 ( .A(n_650), .Y(n_721) );
NAND2xp33_ASAP7_75t_L g725 ( .A(n_651), .B(n_726), .Y(n_725) );
INVx1_ASAP7_75t_L g729 ( .A(n_651), .Y(n_729) );
INVx1_ASAP7_75t_L g755 ( .A(n_652), .Y(n_755) );
AOI21xp5_ASAP7_75t_L g653 ( .A1(n_654), .A2(n_657), .B(n_659), .Y(n_653) );
AND2x4_ASAP7_75t_L g654 ( .A(n_655), .B(n_656), .Y(n_654) );
INVx3_ASAP7_75t_L g704 ( .A(n_656), .Y(n_704) );
AND2x2_ASAP7_75t_L g659 ( .A(n_660), .B(n_661), .Y(n_659) );
INVxp67_ASAP7_75t_L g664 ( .A(n_665), .Y(n_664) );
INVx1_ASAP7_75t_L g665 ( .A(n_666), .Y(n_665) );
AND2x2_ASAP7_75t_L g666 ( .A(n_667), .B(n_669), .Y(n_666) );
INVx2_ASAP7_75t_L g667 ( .A(n_668), .Y(n_667) );
AND2x2_ASAP7_75t_L g781 ( .A(n_668), .B(n_771), .Y(n_781) );
AND2x2_ASAP7_75t_L g684 ( .A(n_669), .B(n_685), .Y(n_684) );
INVx1_ASAP7_75t_L g749 ( .A(n_669), .Y(n_749) );
NAND2xp5_ASAP7_75t_L g670 ( .A(n_671), .B(n_673), .Y(n_670) );
OR2x2_ASAP7_75t_L g707 ( .A(n_672), .B(n_708), .Y(n_707) );
INVx2_ASAP7_75t_L g686 ( .A(n_673), .Y(n_686) );
INVx1_ASAP7_75t_L g674 ( .A(n_675), .Y(n_674) );
NAND2xp5_ASAP7_75t_L g675 ( .A(n_676), .B(n_678), .Y(n_675) );
INVx2_ASAP7_75t_L g676 ( .A(n_677), .Y(n_676) );
AND2x4_ASAP7_75t_L g720 ( .A(n_677), .B(n_721), .Y(n_720) );
INVx1_ASAP7_75t_L g809 ( .A(n_678), .Y(n_809) );
NOR2xp67_ASAP7_75t_L g681 ( .A(n_682), .B(n_718), .Y(n_681) );
NAND3xp33_ASAP7_75t_SL g682 ( .A(n_683), .B(n_693), .C(n_705), .Y(n_682) );
AOI22xp33_ASAP7_75t_L g683 ( .A1(n_684), .A2(n_686), .B1(n_687), .B2(n_688), .Y(n_683) );
INVx1_ASAP7_75t_L g688 ( .A(n_689), .Y(n_688) );
NAND2xp5_ASAP7_75t_L g689 ( .A(n_690), .B(n_691), .Y(n_689) );
INVx1_ASAP7_75t_L g726 ( .A(n_691), .Y(n_726) );
AND2x2_ASAP7_75t_L g801 ( .A(n_691), .B(n_712), .Y(n_801) );
INVx1_ASAP7_75t_L g748 ( .A(n_692), .Y(n_748) );
INVx1_ASAP7_75t_L g693 ( .A(n_694), .Y(n_693) );
OAI32xp33_ASAP7_75t_L g694 ( .A1(n_695), .A2(n_696), .A3(n_698), .B1(n_700), .B2(n_703), .Y(n_694) );
INVx1_ASAP7_75t_L g696 ( .A(n_697), .Y(n_696) );
INVx2_ASAP7_75t_L g728 ( .A(n_697), .Y(n_728) );
NAND2x1_ASAP7_75t_L g766 ( .A(n_697), .B(n_767), .Y(n_766) );
HB1xp67_ASAP7_75t_L g698 ( .A(n_699), .Y(n_698) );
AND2x2_ASAP7_75t_L g727 ( .A(n_699), .B(n_728), .Y(n_727) );
NOR2x1_ASAP7_75t_L g700 ( .A(n_701), .B(n_702), .Y(n_700) );
OAI211xp5_ASAP7_75t_SL g753 ( .A1(n_704), .A2(n_747), .B(n_754), .C(n_755), .Y(n_753) );
INVx2_ASAP7_75t_L g767 ( .A(n_704), .Y(n_767) );
OAI21xp5_ASAP7_75t_L g705 ( .A1(n_706), .A2(n_710), .B(n_717), .Y(n_705) );
INVx1_ASAP7_75t_L g706 ( .A(n_707), .Y(n_706) );
INVx1_ASAP7_75t_L g710 ( .A(n_711), .Y(n_710) );
HB1xp67_ASAP7_75t_L g722 ( .A(n_711), .Y(n_722) );
NAND2x1_ASAP7_75t_L g711 ( .A(n_712), .B(n_714), .Y(n_711) );
INVx2_ASAP7_75t_L g805 ( .A(n_712), .Y(n_805) );
INVx3_ASAP7_75t_L g712 ( .A(n_713), .Y(n_712) );
AND2x2_ASAP7_75t_L g813 ( .A(n_713), .B(n_748), .Y(n_813) );
AND2x2_ASAP7_75t_L g818 ( .A(n_713), .B(n_774), .Y(n_818) );
AND2x4_ASAP7_75t_L g714 ( .A(n_715), .B(n_716), .Y(n_714) );
INVx1_ASAP7_75t_L g743 ( .A(n_716), .Y(n_743) );
OAI211xp5_ASAP7_75t_L g718 ( .A1(n_719), .A2(n_722), .B(n_723), .C(n_730), .Y(n_718) );
INVxp67_ASAP7_75t_SL g719 ( .A(n_720), .Y(n_719) );
NAND2x1p5_ASAP7_75t_L g737 ( .A(n_720), .B(n_738), .Y(n_737) );
NAND2xp5_ASAP7_75t_L g730 ( .A(n_731), .B(n_732), .Y(n_730) );
INVx2_ASAP7_75t_SL g732 ( .A(n_733), .Y(n_732) );
NOR3xp33_ASAP7_75t_L g735 ( .A(n_736), .B(n_768), .C(n_797), .Y(n_735) );
OAI211xp5_ASAP7_75t_L g736 ( .A1(n_737), .A2(n_741), .B(n_744), .C(n_756), .Y(n_736) );
INVx1_ASAP7_75t_L g738 ( .A(n_739), .Y(n_738) );
INVx1_ASAP7_75t_L g739 ( .A(n_740), .Y(n_739) );
AOI22xp5_ASAP7_75t_L g780 ( .A1(n_742), .A2(n_781), .B1(n_782), .B2(n_785), .Y(n_780) );
INVx1_ASAP7_75t_L g742 ( .A(n_743), .Y(n_742) );
AOI22xp5_ASAP7_75t_L g744 ( .A1(n_745), .A2(n_746), .B1(n_752), .B2(n_753), .Y(n_744) );
OAI22xp33_ASAP7_75t_L g746 ( .A1(n_747), .A2(n_749), .B1(n_750), .B2(n_751), .Y(n_746) );
NAND2xp5_ASAP7_75t_L g790 ( .A(n_747), .B(n_779), .Y(n_790) );
INVx1_ASAP7_75t_L g747 ( .A(n_748), .Y(n_747) );
AND2x2_ASAP7_75t_L g761 ( .A(n_754), .B(n_762), .Y(n_761) );
AOI22xp5_ASAP7_75t_L g756 ( .A1(n_757), .A2(n_761), .B1(n_763), .B2(n_765), .Y(n_756) );
INVx1_ASAP7_75t_L g757 ( .A(n_758), .Y(n_757) );
INVx1_ASAP7_75t_L g759 ( .A(n_760), .Y(n_759) );
OR2x2_ASAP7_75t_L g786 ( .A(n_760), .B(n_787), .Y(n_786) );
INVx2_ASAP7_75t_L g763 ( .A(n_764), .Y(n_763) );
INVx1_ASAP7_75t_L g765 ( .A(n_766), .Y(n_765) );
OAI211xp5_ASAP7_75t_SL g768 ( .A1(n_769), .A2(n_775), .B(n_780), .C(n_788), .Y(n_768) );
INVx2_ASAP7_75t_L g769 ( .A(n_770), .Y(n_769) );
AND2x2_ASAP7_75t_L g770 ( .A(n_771), .B(n_772), .Y(n_770) );
INVx1_ASAP7_75t_L g773 ( .A(n_774), .Y(n_773) );
NOR2xp33_ASAP7_75t_L g775 ( .A(n_776), .B(n_777), .Y(n_775) );
INVx2_ASAP7_75t_L g777 ( .A(n_778), .Y(n_777) );
INVx1_ASAP7_75t_L g782 ( .A(n_783), .Y(n_782) );
INVx2_ASAP7_75t_SL g785 ( .A(n_786), .Y(n_785) );
AOI22xp5_ASAP7_75t_L g788 ( .A1(n_789), .A2(n_791), .B1(n_792), .B2(n_794), .Y(n_788) );
INVx1_ASAP7_75t_L g792 ( .A(n_793), .Y(n_792) );
INVx1_ASAP7_75t_L g794 ( .A(n_795), .Y(n_794) );
OAI211xp5_ASAP7_75t_SL g797 ( .A1(n_798), .A2(n_800), .B(n_802), .C(n_810), .Y(n_797) );
INVxp67_ASAP7_75t_L g800 ( .A(n_801), .Y(n_800) );
NAND2xp5_ASAP7_75t_L g802 ( .A(n_803), .B(n_806), .Y(n_802) );
INVx1_ASAP7_75t_L g803 ( .A(n_804), .Y(n_803) );
INVx1_ASAP7_75t_L g806 ( .A(n_807), .Y(n_806) );
OR2x2_ASAP7_75t_L g807 ( .A(n_808), .B(n_809), .Y(n_807) );
INVx4_ASAP7_75t_L g819 ( .A(n_820), .Y(n_819) );
BUFx6f_ASAP7_75t_L g820 ( .A(n_821), .Y(n_820) );
NOR3xp33_ASAP7_75t_L g862 ( .A(n_821), .B(n_863), .C(n_866), .Y(n_862) );
INVx1_ASAP7_75t_L g823 ( .A(n_824), .Y(n_823) );
INVx4_ASAP7_75t_L g824 ( .A(n_825), .Y(n_824) );
AND2x6_ASAP7_75t_SL g825 ( .A(n_826), .B(n_828), .Y(n_825) );
BUFx3_ASAP7_75t_L g834 ( .A(n_826), .Y(n_834) );
INVx1_ASAP7_75t_L g826 ( .A(n_827), .Y(n_826) );
NOR2xp33_ASAP7_75t_L g851 ( .A(n_827), .B(n_852), .Y(n_851) );
NAND2xp5_ASAP7_75t_L g828 ( .A(n_829), .B(n_831), .Y(n_828) );
INVx1_ASAP7_75t_L g829 ( .A(n_830), .Y(n_829) );
NOR2x1_ASAP7_75t_L g854 ( .A(n_830), .B(n_832), .Y(n_854) );
AND2x6_ASAP7_75t_SL g843 ( .A(n_831), .B(n_844), .Y(n_843) );
INVx1_ASAP7_75t_L g831 ( .A(n_832), .Y(n_831) );
OAI21xp5_ASAP7_75t_L g833 ( .A1(n_834), .A2(n_835), .B(n_847), .Y(n_833) );
NAND2xp5_ASAP7_75t_L g835 ( .A(n_836), .B(n_840), .Y(n_835) );
INVx3_ASAP7_75t_L g840 ( .A(n_841), .Y(n_840) );
INVx3_ASAP7_75t_L g841 ( .A(n_842), .Y(n_841) );
CKINVDCx8_ASAP7_75t_R g842 ( .A(n_843), .Y(n_842) );
CKINVDCx5p33_ASAP7_75t_R g856 ( .A(n_843), .Y(n_856) );
INVx1_ASAP7_75t_L g845 ( .A(n_846), .Y(n_845) );
HB1xp67_ASAP7_75t_L g866 ( .A(n_846), .Y(n_866) );
INVx3_ASAP7_75t_L g848 ( .A(n_849), .Y(n_848) );
INVx6_ASAP7_75t_L g849 ( .A(n_850), .Y(n_849) );
BUFx10_ASAP7_75t_L g850 ( .A(n_851), .Y(n_850) );
INVx1_ASAP7_75t_L g852 ( .A(n_853), .Y(n_852) );
NOR2xp33_ASAP7_75t_L g855 ( .A(n_856), .B(n_857), .Y(n_855) );
CKINVDCx6p67_ASAP7_75t_R g858 ( .A(n_859), .Y(n_858) );
BUFx12f_ASAP7_75t_L g859 ( .A(n_860), .Y(n_859) );
INVx4_ASAP7_75t_L g873 ( .A(n_860), .Y(n_873) );
BUFx6f_ASAP7_75t_L g860 ( .A(n_861), .Y(n_860) );
NAND2xp5_ASAP7_75t_SL g861 ( .A(n_862), .B(n_867), .Y(n_861) );
INVx2_ASAP7_75t_SL g863 ( .A(n_864), .Y(n_863) );
NOR2x1p5_ASAP7_75t_L g867 ( .A(n_868), .B(n_869), .Y(n_867) );
INVx1_ASAP7_75t_L g869 ( .A(n_870), .Y(n_869) );
NOR2xp33_ASAP7_75t_L g871 ( .A(n_872), .B(n_873), .Y(n_871) );
endmodule