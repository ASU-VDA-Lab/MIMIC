module real_aes_8453_n_99 (n_17, n_28, n_76, n_56, n_34, n_98, n_90, n_82, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_714, n_18, n_21, n_31, n_8, n_10, n_83, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_91, n_43, n_96, n_54, n_35, n_42, n_15, n_9, n_23, n_72, n_95, n_44, n_7, n_4, n_80, n_6, n_12, n_68, n_79, n_69, n_46, n_59, n_25, n_73, n_77, n_81, n_48, n_37, n_97, n_70, n_50, n_89, n_26, n_86, n_93, n_13, n_24, n_2, n_55, n_62, n_84, n_67, n_92, n_33, n_88, n_14, n_11, n_85, n_16, n_94, n_39, n_5, n_45, n_60, n_38, n_87, n_0, n_78, n_63, n_1, n_53, n_36, n_99);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_98;
input n_90;
input n_82;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_714;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_83;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_91;
input n_43;
input n_96;
input n_54;
input n_35;
input n_42;
input n_15;
input n_9;
input n_23;
input n_72;
input n_95;
input n_44;
input n_7;
input n_4;
input n_80;
input n_6;
input n_12;
input n_68;
input n_79;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_81;
input n_48;
input n_37;
input n_97;
input n_70;
input n_50;
input n_89;
input n_26;
input n_86;
input n_93;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_84;
input n_67;
input n_92;
input n_33;
input n_88;
input n_14;
input n_11;
input n_85;
input n_16;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_87;
input n_0;
input n_78;
input n_63;
input n_1;
input n_53;
input n_36;
output n_99;
wire n_480;
wire n_113;
wire n_476;
wire n_599;
wire n_187;
wire n_436;
wire n_684;
wire n_257;
wire n_390;
wire n_185;
wire n_285;
wire n_624;
wire n_618;
wire n_522;
wire n_485;
wire n_222;
wire n_631;
wire n_287;
wire n_357;
wire n_503;
wire n_635;
wire n_386;
wire n_673;
wire n_518;
wire n_254;
wire n_207;
wire n_665;
wire n_667;
wire n_580;
wire n_577;
wire n_469;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_318;
wire n_355;
wire n_239;
wire n_669;
wire n_100;
wire n_423;
wire n_458;
wire n_444;
wire n_112;
wire n_319;
wire n_364;
wire n_421;
wire n_555;
wire n_329;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_242;
wire n_169;
wire n_376;
wire n_549;
wire n_571;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_448;
wire n_545;
wire n_341;
wire n_556;
wire n_593;
wire n_232;
wire n_460;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_551;
wire n_320;
wire n_537;
wire n_666;
wire n_560;
wire n_260;
wire n_660;
wire n_594;
wire n_186;
wire n_138;
wire n_696;
wire n_704;
wire n_379;
wire n_374;
wire n_453;
wire n_647;
wire n_235;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_161;
wire n_189;
wire n_271;
wire n_489;
wire n_427;
wire n_548;
wire n_678;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_564;
wire n_519;
wire n_638;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_512;
wire n_395;
wire n_332;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_116;
wire n_625;
wire n_289;
wire n_462;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_213;
wire n_356;
wire n_478;
wire n_584;
wire n_408;
wire n_553;
wire n_184;
wire n_372;
wire n_528;
wire n_578;
wire n_202;
wire n_495;
wire n_370;
wire n_384;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_467;
wire n_327;
wire n_106;
wire n_466;
wire n_559;
wire n_636;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_517;
wire n_683;
wire n_174;
wire n_570;
wire n_675;
wire n_530;
wire n_104;
wire n_535;
wire n_211;
wire n_281;
wire n_496;
wire n_693;
wire n_173;
wire n_468;
wire n_234;
wire n_284;
wire n_153;
wire n_316;
wire n_532;
wire n_656;
wire n_178;
wire n_409;
wire n_298;
wire n_523;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_297;
wire n_383;
wire n_529;
wire n_455;
wire n_119;
wire n_310;
wire n_504;
wire n_164;
wire n_671;
wire n_231;
wire n_102;
wire n_547;
wire n_659;
wire n_634;
wire n_682;
wire n_454;
wire n_122;
wire n_443;
wire n_565;
wire n_608;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_267;
wire n_218;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_331;
wire n_182;
wire n_363;
wire n_417;
wire n_449;
wire n_607;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_142;
wire n_561;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_655;
wire n_654;
wire n_505;
wire n_434;
wire n_502;
wire n_527;
wire n_600;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_602;
wire n_402;
wire n_552;
wire n_617;
wire n_171;
wire n_676;
wire n_658;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_146;
wire n_432;
wire n_226;
wire n_255;
wire n_286;
wire n_416;
wire n_410;
wire n_120;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_695;
wire n_685;
wire n_165;
wire n_361;
wire n_632;
wire n_246;
wire n_176;
wire n_412;
wire n_163;
wire n_542;
wire n_645;
wire n_557;
wire n_501;
wire n_488;
wire n_251;
wire n_642;
wire n_613;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_702;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_110;
wire n_392;
wire n_562;
wire n_150;
wire n_147;
wire n_288;
wire n_404;
wire n_598;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_569;
wire n_563;
wire n_188;
wire n_430;
wire n_269;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_193;
wire n_397;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_649;
wire n_663;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_707;
wire n_622;
wire n_470;
wire n_133;
wire n_494;
wire n_711;
wire n_377;
wire n_273;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_265;
wire n_354;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_643;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_148;
wire n_498;
wire n_481;
wire n_691;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_233;
wire n_487;
wire n_290;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_155;
wire n_243;
wire n_692;
wire n_544;
wire n_268;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_101;
wire n_701;
wire n_309;
wire n_344;
wire n_107;
wire n_229;
wire n_482;
wire n_520;
wire n_633;
wire n_679;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_262;
wire n_630;
wire n_689;
wire n_134;
wire n_349;
wire n_336;
wire n_420;
wire n_612;
wire n_195;
wire n_438;
wire n_300;
wire n_252;
wire n_314;
wire n_283;
wire n_249;
wire n_623;
wire n_446;
wire n_221;
wire n_681;
wire n_156;
wire n_456;
wire n_359;
wire n_312;
wire n_183;
wire n_266;
wire n_712;
wire n_205;
wire n_433;
wire n_335;
wire n_177;
wire n_516;
wire n_313;
wire n_627;
wire n_521;
wire n_140;
wire n_418;
wire n_422;
wire n_524;
wire n_219;
wire n_705;
wire n_180;
wire n_212;
wire n_210;
wire n_575;
wire n_325;
wire n_338;
wire n_479;
wire n_442;
wire n_698;
wire n_371;
wire n_103;
wire n_166;
wire n_541;
wire n_224;
wire n_151;
wire n_546;
wire n_639;
wire n_587;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_440;
wire n_525;
wire n_644;
wire n_674;
wire n_152;
wire n_198;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_414;
wire n_123;
wire n_279;
wire n_686;
wire n_543;
wire n_497;
wire n_514;
wire n_507;
wire n_270;
wire n_614;
wire n_305;
wire n_586;
wire n_450;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_473;
wire n_465;
wire n_566;
wire n_474;
wire n_170;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_168;
wire n_175;
wire n_241;
wire n_687;
wire n_646;
wire n_710;
wire n_650;
wire n_105;
wire n_294;
wire n_393;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_500;
wire n_307;
wire n_601;
wire n_661;
wire n_463;
wire n_396;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_194;
wire n_137;
wire n_424;
wire n_225;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_143;
wire n_192;
wire n_475;
wire n_554;
wire n_264;
wire n_237;
wire n_668;
A2O1A1Ixp33_ASAP7_75t_SL g443 ( .A1(n_0), .A2(n_181), .B(n_444), .C(n_447), .Y(n_443) );
NAND2xp5_ASAP7_75t_L g448 ( .A(n_1), .B(n_438), .Y(n_448) );
INVx1_ASAP7_75t_L g678 ( .A(n_2), .Y(n_678) );
INVx1_ASAP7_75t_L g216 ( .A(n_3), .Y(n_216) );
NAND2xp5_ASAP7_75t_SL g428 ( .A(n_4), .B(n_133), .Y(n_428) );
AOI21xp5_ASAP7_75t_L g520 ( .A1(n_5), .A2(n_433), .B(n_521), .Y(n_520) );
AO21x2_ASAP7_75t_L g482 ( .A1(n_6), .A2(n_156), .B(n_483), .Y(n_482) );
AOI22xp33_ASAP7_75t_L g180 ( .A1(n_7), .A2(n_36), .B1(n_126), .B2(n_150), .Y(n_180) );
NAND2xp5_ASAP7_75t_L g228 ( .A(n_8), .B(n_156), .Y(n_228) );
AND2x6_ASAP7_75t_L g141 ( .A(n_9), .B(n_142), .Y(n_141) );
A2O1A1Ixp33_ASAP7_75t_L g496 ( .A1(n_10), .A2(n_141), .B(n_424), .C(n_497), .Y(n_496) );
NOR2xp33_ASAP7_75t_L g679 ( .A(n_11), .B(n_37), .Y(n_679) );
INVx1_ASAP7_75t_L g122 ( .A(n_12), .Y(n_122) );
NAND2xp5_ASAP7_75t_L g164 ( .A(n_13), .B(n_131), .Y(n_164) );
INVx1_ASAP7_75t_L g208 ( .A(n_14), .Y(n_208) );
NAND2xp5_ASAP7_75t_SL g488 ( .A(n_15), .B(n_133), .Y(n_488) );
NAND2xp5_ASAP7_75t_L g195 ( .A(n_16), .B(n_157), .Y(n_195) );
AO32x2_ASAP7_75t_L g178 ( .A1(n_17), .A2(n_155), .A3(n_156), .B1(n_179), .B2(n_183), .Y(n_178) );
NAND2xp5_ASAP7_75t_SL g168 ( .A(n_18), .B(n_126), .Y(n_168) );
NAND2xp5_ASAP7_75t_L g218 ( .A(n_19), .B(n_157), .Y(n_218) );
AOI22xp33_ASAP7_75t_L g182 ( .A1(n_20), .A2(n_52), .B1(n_126), .B2(n_150), .Y(n_182) );
AOI22xp33_ASAP7_75t_SL g153 ( .A1(n_21), .A2(n_78), .B1(n_126), .B2(n_131), .Y(n_153) );
NAND2xp5_ASAP7_75t_SL g137 ( .A(n_22), .B(n_126), .Y(n_137) );
A2O1A1Ixp33_ASAP7_75t_L g470 ( .A1(n_23), .A2(n_155), .B(n_424), .C(n_471), .Y(n_470) );
A2O1A1Ixp33_ASAP7_75t_L g485 ( .A1(n_24), .A2(n_155), .B(n_424), .C(n_486), .Y(n_485) );
BUFx6f_ASAP7_75t_L g135 ( .A(n_25), .Y(n_135) );
NAND2xp5_ASAP7_75t_L g237 ( .A(n_26), .B(n_118), .Y(n_237) );
OAI22xp5_ASAP7_75t_L g102 ( .A1(n_27), .A2(n_103), .B1(n_104), .B2(n_105), .Y(n_102) );
CKINVDCx20_ASAP7_75t_R g103 ( .A(n_27), .Y(n_103) );
AOI21xp5_ASAP7_75t_L g439 ( .A1(n_28), .A2(n_433), .B(n_440), .Y(n_439) );
NAND2xp5_ASAP7_75t_L g143 ( .A(n_29), .B(n_118), .Y(n_143) );
INVx2_ASAP7_75t_L g128 ( .A(n_30), .Y(n_128) );
A2O1A1Ixp33_ASAP7_75t_L g455 ( .A1(n_31), .A2(n_430), .B(n_456), .C(n_457), .Y(n_455) );
NAND2xp5_ASAP7_75t_SL g232 ( .A(n_32), .B(n_126), .Y(n_232) );
NAND2xp5_ASAP7_75t_L g171 ( .A(n_33), .B(n_118), .Y(n_171) );
AOI222xp33_ASAP7_75t_L g99 ( .A1(n_34), .A2(n_100), .B1(n_683), .B2(n_692), .C1(n_704), .C2(n_710), .Y(n_99) );
OAI22xp5_ASAP7_75t_SL g697 ( .A1(n_34), .A2(n_41), .B1(n_414), .B2(n_698), .Y(n_697) );
CKINVDCx20_ASAP7_75t_R g698 ( .A(n_34), .Y(n_698) );
NAND2xp5_ASAP7_75t_L g487 ( .A(n_35), .B(n_166), .Y(n_487) );
NAND2xp5_ASAP7_75t_L g468 ( .A(n_38), .B(n_469), .Y(n_468) );
CKINVDCx20_ASAP7_75t_R g501 ( .A(n_39), .Y(n_501) );
NAND2xp5_ASAP7_75t_L g509 ( .A(n_40), .B(n_133), .Y(n_509) );
OAI22xp5_ASAP7_75t_SL g108 ( .A1(n_41), .A2(n_109), .B1(n_414), .B2(n_415), .Y(n_108) );
INVx1_ASAP7_75t_L g414 ( .A(n_41), .Y(n_414) );
NAND2xp5_ASAP7_75t_L g484 ( .A(n_42), .B(n_433), .Y(n_484) );
A2O1A1Ixp33_ASAP7_75t_L g506 ( .A1(n_43), .A2(n_430), .B(n_456), .C(n_507), .Y(n_506) );
NAND2xp5_ASAP7_75t_SL g223 ( .A(n_44), .B(n_126), .Y(n_223) );
INVx1_ASAP7_75t_L g445 ( .A(n_45), .Y(n_445) );
AOI22xp33_ASAP7_75t_L g149 ( .A1(n_46), .A2(n_86), .B1(n_150), .B2(n_151), .Y(n_149) );
INVx1_ASAP7_75t_L g508 ( .A(n_47), .Y(n_508) );
NAND2xp5_ASAP7_75t_SL g226 ( .A(n_48), .B(n_126), .Y(n_226) );
NAND2xp5_ASAP7_75t_L g210 ( .A(n_49), .B(n_126), .Y(n_210) );
NAND2xp5_ASAP7_75t_L g505 ( .A(n_50), .B(n_433), .Y(n_505) );
NAND2xp5_ASAP7_75t_L g227 ( .A(n_51), .B(n_214), .Y(n_227) );
AOI22xp33_ASAP7_75t_SL g199 ( .A1(n_53), .A2(n_57), .B1(n_126), .B2(n_131), .Y(n_199) );
CKINVDCx20_ASAP7_75t_R g476 ( .A(n_54), .Y(n_476) );
NAND2xp5_ASAP7_75t_SL g163 ( .A(n_55), .B(n_126), .Y(n_163) );
NAND2xp5_ASAP7_75t_SL g236 ( .A(n_56), .B(n_126), .Y(n_236) );
INVx1_ASAP7_75t_L g142 ( .A(n_58), .Y(n_142) );
NAND2xp5_ASAP7_75t_L g432 ( .A(n_59), .B(n_433), .Y(n_432) );
NAND2xp5_ASAP7_75t_L g526 ( .A(n_60), .B(n_438), .Y(n_526) );
A2O1A1Ixp33_ASAP7_75t_L g523 ( .A1(n_61), .A2(n_211), .B(n_214), .C(n_524), .Y(n_523) );
NAND2xp5_ASAP7_75t_L g217 ( .A(n_62), .B(n_126), .Y(n_217) );
INVx1_ASAP7_75t_L g121 ( .A(n_63), .Y(n_121) );
CKINVDCx20_ASAP7_75t_R g688 ( .A(n_64), .Y(n_688) );
NAND2xp5_ASAP7_75t_SL g461 ( .A(n_65), .B(n_133), .Y(n_461) );
AO32x2_ASAP7_75t_L g147 ( .A1(n_66), .A2(n_148), .A3(n_154), .B1(n_155), .B2(n_156), .Y(n_147) );
NAND2xp5_ASAP7_75t_L g498 ( .A(n_67), .B(n_134), .Y(n_498) );
INVx1_ASAP7_75t_L g235 ( .A(n_68), .Y(n_235) );
INVx1_ASAP7_75t_L g129 ( .A(n_69), .Y(n_129) );
CKINVDCx16_ASAP7_75t_R g441 ( .A(n_70), .Y(n_441) );
NAND2xp5_ASAP7_75t_L g472 ( .A(n_71), .B(n_460), .Y(n_472) );
A2O1A1Ixp33_ASAP7_75t_L g423 ( .A1(n_72), .A2(n_424), .B(n_426), .C(n_430), .Y(n_423) );
NAND2xp5_ASAP7_75t_SL g130 ( .A(n_73), .B(n_131), .Y(n_130) );
CKINVDCx16_ASAP7_75t_R g522 ( .A(n_74), .Y(n_522) );
INVx1_ASAP7_75t_L g687 ( .A(n_75), .Y(n_687) );
NAND2xp5_ASAP7_75t_SL g473 ( .A(n_76), .B(n_459), .Y(n_473) );
AOI22xp5_ASAP7_75t_SL g101 ( .A1(n_77), .A2(n_102), .B1(n_676), .B2(n_680), .Y(n_101) );
NAND2xp5_ASAP7_75t_L g169 ( .A(n_79), .B(n_150), .Y(n_169) );
CKINVDCx20_ASAP7_75t_R g464 ( .A(n_80), .Y(n_464) );
NAND2xp5_ASAP7_75t_SL g138 ( .A(n_81), .B(n_131), .Y(n_138) );
INVx2_ASAP7_75t_L g119 ( .A(n_82), .Y(n_119) );
CKINVDCx20_ASAP7_75t_R g436 ( .A(n_83), .Y(n_436) );
NAND2xp5_ASAP7_75t_SL g499 ( .A(n_84), .B(n_152), .Y(n_499) );
NAND2xp5_ASAP7_75t_L g224 ( .A(n_85), .B(n_131), .Y(n_224) );
INVx2_ASAP7_75t_L g107 ( .A(n_87), .Y(n_107) );
OR2x2_ASAP7_75t_L g691 ( .A(n_87), .B(n_676), .Y(n_691) );
AOI22xp33_ASAP7_75t_L g198 ( .A1(n_88), .A2(n_98), .B1(n_131), .B2(n_132), .Y(n_198) );
NAND2xp5_ASAP7_75t_L g454 ( .A(n_89), .B(n_433), .Y(n_454) );
INVx1_ASAP7_75t_L g458 ( .A(n_90), .Y(n_458) );
CKINVDCx20_ASAP7_75t_R g701 ( .A(n_91), .Y(n_701) );
INVxp67_ASAP7_75t_L g525 ( .A(n_92), .Y(n_525) );
NAND2xp5_ASAP7_75t_L g233 ( .A(n_93), .B(n_131), .Y(n_233) );
INVx1_ASAP7_75t_L g427 ( .A(n_94), .Y(n_427) );
INVx1_ASAP7_75t_L g494 ( .A(n_95), .Y(n_494) );
NAND2xp5_ASAP7_75t_L g686 ( .A(n_96), .B(n_687), .Y(n_686) );
AND2x2_ASAP7_75t_L g510 ( .A(n_97), .B(n_118), .Y(n_510) );
INVxp67_ASAP7_75t_L g100 ( .A(n_101), .Y(n_100) );
INVx1_ASAP7_75t_L g104 ( .A(n_105), .Y(n_104) );
INVx1_ASAP7_75t_L g105 ( .A(n_106), .Y(n_105) );
AO22x2_ASAP7_75t_SL g106 ( .A1(n_107), .A2(n_108), .B1(n_416), .B2(n_675), .Y(n_106) );
INVx1_ASAP7_75t_L g675 ( .A(n_107), .Y(n_675) );
NOR2x2_ASAP7_75t_L g682 ( .A(n_107), .B(n_676), .Y(n_682) );
INVx1_ASAP7_75t_L g415 ( .A(n_109), .Y(n_415) );
OAI22xp5_ASAP7_75t_SL g695 ( .A1(n_109), .A2(n_415), .B1(n_696), .B2(n_697), .Y(n_695) );
OR2x2_ASAP7_75t_L g109 ( .A(n_110), .B(n_335), .Y(n_109) );
NAND3xp33_ASAP7_75t_L g110 ( .A(n_111), .B(n_284), .C(n_326), .Y(n_110) );
AOI211xp5_ASAP7_75t_L g111 ( .A1(n_112), .A2(n_189), .B(n_238), .C(n_260), .Y(n_111) );
OAI211xp5_ASAP7_75t_SL g112 ( .A1(n_113), .A2(n_144), .B(n_172), .C(n_184), .Y(n_112) );
INVxp67_ASAP7_75t_L g113 ( .A(n_114), .Y(n_113) );
NAND2xp5_ASAP7_75t_L g241 ( .A(n_114), .B(n_242), .Y(n_241) );
AND2x2_ASAP7_75t_L g347 ( .A(n_114), .B(n_264), .Y(n_347) );
BUFx2_ASAP7_75t_L g114 ( .A(n_115), .Y(n_114) );
AND2x2_ASAP7_75t_L g249 ( .A(n_115), .B(n_175), .Y(n_249) );
NAND2xp5_ASAP7_75t_L g366 ( .A(n_115), .B(n_160), .Y(n_366) );
INVx1_ASAP7_75t_L g384 ( .A(n_115), .Y(n_384) );
AND2x2_ASAP7_75t_L g393 ( .A(n_115), .B(n_281), .Y(n_393) );
INVx2_ASAP7_75t_L g115 ( .A(n_116), .Y(n_115) );
OR2x2_ASAP7_75t_L g276 ( .A(n_116), .B(n_160), .Y(n_276) );
AND2x2_ASAP7_75t_L g334 ( .A(n_116), .B(n_281), .Y(n_334) );
INVx1_ASAP7_75t_L g378 ( .A(n_116), .Y(n_378) );
INVx2_ASAP7_75t_L g116 ( .A(n_117), .Y(n_116) );
OR2x2_ASAP7_75t_L g255 ( .A(n_117), .B(n_256), .Y(n_255) );
INVx2_ASAP7_75t_L g263 ( .A(n_117), .Y(n_263) );
HB1xp67_ASAP7_75t_L g303 ( .A(n_117), .Y(n_303) );
OA21x2_ASAP7_75t_L g117 ( .A1(n_118), .A2(n_123), .B(n_143), .Y(n_117) );
INVx2_ASAP7_75t_L g154 ( .A(n_118), .Y(n_154) );
OA21x2_ASAP7_75t_L g160 ( .A1(n_118), .A2(n_161), .B(n_171), .Y(n_160) );
AOI21xp5_ASAP7_75t_L g453 ( .A1(n_118), .A2(n_454), .B(n_455), .Y(n_453) );
INVx1_ASAP7_75t_L g477 ( .A(n_118), .Y(n_477) );
AOI21xp5_ASAP7_75t_L g504 ( .A1(n_118), .A2(n_505), .B(n_506), .Y(n_504) );
AND2x2_ASAP7_75t_SL g118 ( .A(n_119), .B(n_120), .Y(n_118) );
AND2x2_ASAP7_75t_L g157 ( .A(n_119), .B(n_120), .Y(n_157) );
NAND2xp5_ASAP7_75t_L g120 ( .A(n_121), .B(n_122), .Y(n_120) );
OAI21xp5_ASAP7_75t_L g123 ( .A1(n_124), .A2(n_136), .B(n_141), .Y(n_123) );
O2A1O1Ixp5_ASAP7_75t_SL g124 ( .A1(n_125), .A2(n_129), .B(n_130), .C(n_133), .Y(n_124) );
INVx3_ASAP7_75t_L g125 ( .A(n_126), .Y(n_125) );
HB1xp67_ASAP7_75t_L g429 ( .A(n_126), .Y(n_429) );
BUFx6f_ASAP7_75t_L g126 ( .A(n_127), .Y(n_126) );
INVx1_ASAP7_75t_L g150 ( .A(n_127), .Y(n_150) );
BUFx3_ASAP7_75t_L g151 ( .A(n_127), .Y(n_151) );
AND2x6_ASAP7_75t_L g424 ( .A(n_127), .B(n_425), .Y(n_424) );
INVx2_ASAP7_75t_L g127 ( .A(n_128), .Y(n_127) );
INVx1_ASAP7_75t_L g132 ( .A(n_128), .Y(n_132) );
INVx1_ASAP7_75t_L g215 ( .A(n_128), .Y(n_215) );
INVx2_ASAP7_75t_L g209 ( .A(n_131), .Y(n_209) );
INVx3_ASAP7_75t_L g131 ( .A(n_132), .Y(n_131) );
INVx2_ASAP7_75t_L g181 ( .A(n_133), .Y(n_181) );
AOI21xp5_ASAP7_75t_L g222 ( .A1(n_133), .A2(n_223), .B(n_224), .Y(n_222) );
AOI21xp5_ASAP7_75t_L g231 ( .A1(n_133), .A2(n_232), .B(n_233), .Y(n_231) );
NOR2xp33_ASAP7_75t_L g524 ( .A(n_133), .B(n_525), .Y(n_524) );
INVx5_ASAP7_75t_L g133 ( .A(n_134), .Y(n_133) );
OAI22xp5_ASAP7_75t_SL g148 ( .A1(n_134), .A2(n_149), .B1(n_152), .B2(n_153), .Y(n_148) );
INVx3_ASAP7_75t_L g134 ( .A(n_135), .Y(n_134) );
BUFx6f_ASAP7_75t_L g140 ( .A(n_135), .Y(n_140) );
BUFx6f_ASAP7_75t_L g152 ( .A(n_135), .Y(n_152) );
INVx1_ASAP7_75t_L g166 ( .A(n_135), .Y(n_166) );
INVx1_ASAP7_75t_L g425 ( .A(n_135), .Y(n_425) );
AND2x2_ASAP7_75t_L g434 ( .A(n_135), .B(n_215), .Y(n_434) );
AOI21xp5_ASAP7_75t_L g136 ( .A1(n_137), .A2(n_138), .B(n_139), .Y(n_136) );
INVx1_ASAP7_75t_L g211 ( .A(n_139), .Y(n_211) );
INVx4_ASAP7_75t_L g139 ( .A(n_140), .Y(n_139) );
INVx2_ASAP7_75t_L g460 ( .A(n_140), .Y(n_460) );
BUFx3_ASAP7_75t_L g155 ( .A(n_141), .Y(n_155) );
OAI21xp5_ASAP7_75t_L g161 ( .A1(n_141), .A2(n_162), .B(n_167), .Y(n_161) );
OAI21xp5_ASAP7_75t_L g206 ( .A1(n_141), .A2(n_207), .B(n_212), .Y(n_206) );
OAI21xp5_ASAP7_75t_L g221 ( .A1(n_141), .A2(n_222), .B(n_225), .Y(n_221) );
INVx4_ASAP7_75t_SL g431 ( .A(n_141), .Y(n_431) );
AND2x4_ASAP7_75t_L g433 ( .A(n_141), .B(n_434), .Y(n_433) );
NAND2x1p5_ASAP7_75t_L g495 ( .A(n_141), .B(n_434), .Y(n_495) );
INVxp67_ASAP7_75t_L g144 ( .A(n_145), .Y(n_144) );
NAND2xp5_ASAP7_75t_L g145 ( .A(n_146), .B(n_158), .Y(n_145) );
AND2x2_ASAP7_75t_L g242 ( .A(n_146), .B(n_243), .Y(n_242) );
INVx2_ASAP7_75t_L g275 ( .A(n_146), .Y(n_275) );
OR2x2_ASAP7_75t_L g401 ( .A(n_146), .B(n_402), .Y(n_401) );
NOR2xp33_ASAP7_75t_L g405 ( .A(n_146), .B(n_160), .Y(n_405) );
BUFx6f_ASAP7_75t_L g146 ( .A(n_147), .Y(n_146) );
INVx1_ASAP7_75t_L g175 ( .A(n_147), .Y(n_175) );
INVx1_ASAP7_75t_L g187 ( .A(n_147), .Y(n_187) );
AND2x2_ASAP7_75t_L g264 ( .A(n_147), .B(n_177), .Y(n_264) );
AND2x2_ASAP7_75t_L g304 ( .A(n_147), .B(n_178), .Y(n_304) );
INVx2_ASAP7_75t_L g447 ( .A(n_151), .Y(n_447) );
HB1xp67_ASAP7_75t_L g462 ( .A(n_151), .Y(n_462) );
INVx2_ASAP7_75t_L g170 ( .A(n_152), .Y(n_170) );
OAI22xp5_ASAP7_75t_L g179 ( .A1(n_152), .A2(n_180), .B1(n_181), .B2(n_182), .Y(n_179) );
OAI22xp5_ASAP7_75t_L g197 ( .A1(n_152), .A2(n_181), .B1(n_198), .B2(n_199), .Y(n_197) );
INVx4_ASAP7_75t_L g446 ( .A(n_152), .Y(n_446) );
INVx1_ASAP7_75t_L g474 ( .A(n_154), .Y(n_474) );
NAND3xp33_ASAP7_75t_L g196 ( .A(n_155), .B(n_197), .C(n_200), .Y(n_196) );
OAI21xp5_ASAP7_75t_L g230 ( .A1(n_155), .A2(n_231), .B(n_234), .Y(n_230) );
INVx4_ASAP7_75t_L g200 ( .A(n_156), .Y(n_200) );
OA21x2_ASAP7_75t_L g220 ( .A1(n_156), .A2(n_221), .B(n_228), .Y(n_220) );
AOI21xp5_ASAP7_75t_L g483 ( .A1(n_156), .A2(n_484), .B(n_485), .Y(n_483) );
HB1xp67_ASAP7_75t_L g519 ( .A(n_156), .Y(n_519) );
BUFx6f_ASAP7_75t_L g156 ( .A(n_157), .Y(n_156) );
INVx1_ASAP7_75t_L g183 ( .A(n_157), .Y(n_183) );
INVxp67_ASAP7_75t_L g346 ( .A(n_158), .Y(n_346) );
AND2x4_ASAP7_75t_L g371 ( .A(n_158), .B(n_264), .Y(n_371) );
BUFx3_ASAP7_75t_L g158 ( .A(n_159), .Y(n_158) );
AND2x2_ASAP7_75t_SL g262 ( .A(n_159), .B(n_263), .Y(n_262) );
INVx1_ASAP7_75t_L g159 ( .A(n_160), .Y(n_159) );
AND2x2_ASAP7_75t_L g176 ( .A(n_160), .B(n_177), .Y(n_176) );
AND2x2_ASAP7_75t_L g250 ( .A(n_160), .B(n_178), .Y(n_250) );
INVx1_ASAP7_75t_L g256 ( .A(n_160), .Y(n_256) );
INVx2_ASAP7_75t_L g282 ( .A(n_160), .Y(n_282) );
AND2x2_ASAP7_75t_L g298 ( .A(n_160), .B(n_299), .Y(n_298) );
AOI21xp5_ASAP7_75t_L g162 ( .A1(n_163), .A2(n_164), .B(n_165), .Y(n_162) );
INVx1_ASAP7_75t_L g165 ( .A(n_166), .Y(n_165) );
AOI21xp5_ASAP7_75t_L g167 ( .A1(n_168), .A2(n_169), .B(n_170), .Y(n_167) );
O2A1O1Ixp5_ASAP7_75t_L g234 ( .A1(n_170), .A2(n_213), .B(n_235), .C(n_236), .Y(n_234) );
INVx1_ASAP7_75t_L g172 ( .A(n_173), .Y(n_172) );
NAND2xp5_ASAP7_75t_L g286 ( .A(n_173), .B(n_287), .Y(n_286) );
AND2x2_ASAP7_75t_L g173 ( .A(n_174), .B(n_176), .Y(n_173) );
INVx1_ASAP7_75t_L g174 ( .A(n_175), .Y(n_174) );
BUFx2_ASAP7_75t_L g253 ( .A(n_175), .Y(n_253) );
AND2x2_ASAP7_75t_L g361 ( .A(n_175), .B(n_177), .Y(n_361) );
AND2x2_ASAP7_75t_L g278 ( .A(n_176), .B(n_263), .Y(n_278) );
AND2x2_ASAP7_75t_L g377 ( .A(n_176), .B(n_378), .Y(n_377) );
NOR2xp67_ASAP7_75t_L g299 ( .A(n_177), .B(n_300), .Y(n_299) );
OR2x2_ASAP7_75t_L g402 ( .A(n_177), .B(n_263), .Y(n_402) );
INVx2_ASAP7_75t_L g177 ( .A(n_178), .Y(n_177) );
BUFx2_ASAP7_75t_L g188 ( .A(n_178), .Y(n_188) );
AND2x2_ASAP7_75t_L g281 ( .A(n_178), .B(n_282), .Y(n_281) );
O2A1O1Ixp33_ASAP7_75t_L g212 ( .A1(n_181), .A2(n_213), .B(n_216), .C(n_217), .Y(n_212) );
AOI21xp5_ASAP7_75t_L g225 ( .A1(n_181), .A2(n_226), .B(n_227), .Y(n_225) );
INVx2_ASAP7_75t_L g205 ( .A(n_183), .Y(n_205) );
NOR2xp33_ASAP7_75t_L g500 ( .A(n_183), .B(n_501), .Y(n_500) );
INVx1_ASAP7_75t_L g184 ( .A(n_185), .Y(n_184) );
AND2x2_ASAP7_75t_L g185 ( .A(n_186), .B(n_188), .Y(n_185) );
AND2x2_ASAP7_75t_L g327 ( .A(n_186), .B(n_262), .Y(n_327) );
HB1xp67_ASAP7_75t_L g186 ( .A(n_187), .Y(n_186) );
NAND2xp5_ASAP7_75t_L g312 ( .A(n_187), .B(n_263), .Y(n_312) );
INVx2_ASAP7_75t_L g311 ( .A(n_188), .Y(n_311) );
OAI222xp33_ASAP7_75t_L g315 ( .A1(n_188), .A2(n_255), .B1(n_316), .B2(n_318), .C1(n_319), .C2(n_322), .Y(n_315) );
INVx1_ASAP7_75t_L g189 ( .A(n_190), .Y(n_189) );
NAND2xp5_ASAP7_75t_L g190 ( .A(n_191), .B(n_201), .Y(n_190) );
INVx1_ASAP7_75t_L g191 ( .A(n_192), .Y(n_191) );
INVx1_ASAP7_75t_L g192 ( .A(n_193), .Y(n_192) );
INVx2_ASAP7_75t_L g240 ( .A(n_193), .Y(n_240) );
OR2x2_ASAP7_75t_L g351 ( .A(n_193), .B(n_352), .Y(n_351) );
INVx2_ASAP7_75t_L g193 ( .A(n_194), .Y(n_193) );
INVx3_ASAP7_75t_L g273 ( .A(n_194), .Y(n_273) );
NOR2x1_ASAP7_75t_L g324 ( .A(n_194), .B(n_325), .Y(n_324) );
AND2x2_ASAP7_75t_L g330 ( .A(n_194), .B(n_244), .Y(n_330) );
AND2x4_ASAP7_75t_L g194 ( .A(n_195), .B(n_196), .Y(n_194) );
INVx1_ASAP7_75t_L g291 ( .A(n_195), .Y(n_291) );
AO21x1_ASAP7_75t_L g290 ( .A1(n_197), .A2(n_200), .B(n_291), .Y(n_290) );
AO21x2_ASAP7_75t_L g421 ( .A1(n_200), .A2(n_422), .B(n_435), .Y(n_421) );
NOR2xp33_ASAP7_75t_L g435 ( .A(n_200), .B(n_436), .Y(n_435) );
INVx3_ASAP7_75t_L g438 ( .A(n_200), .Y(n_438) );
NOR2xp33_ASAP7_75t_L g463 ( .A(n_200), .B(n_464), .Y(n_463) );
AO21x2_ASAP7_75t_L g492 ( .A1(n_200), .A2(n_493), .B(n_500), .Y(n_492) );
AOI22xp5_ASAP7_75t_L g332 ( .A1(n_201), .A2(n_294), .B1(n_333), .B2(n_334), .Y(n_332) );
AND2x2_ASAP7_75t_L g201 ( .A(n_202), .B(n_219), .Y(n_201) );
INVx3_ASAP7_75t_L g266 ( .A(n_202), .Y(n_266) );
OR2x2_ASAP7_75t_L g399 ( .A(n_202), .B(n_275), .Y(n_399) );
INVx2_ASAP7_75t_L g202 ( .A(n_203), .Y(n_202) );
AND2x2_ASAP7_75t_L g272 ( .A(n_203), .B(n_273), .Y(n_272) );
AND2x2_ASAP7_75t_L g288 ( .A(n_203), .B(n_289), .Y(n_288) );
AND2x2_ASAP7_75t_L g296 ( .A(n_203), .B(n_244), .Y(n_296) );
NAND2xp5_ASAP7_75t_L g352 ( .A(n_203), .B(n_220), .Y(n_352) );
INVx2_ASAP7_75t_L g203 ( .A(n_204), .Y(n_203) );
AND2x2_ASAP7_75t_L g243 ( .A(n_204), .B(n_244), .Y(n_243) );
AND2x2_ASAP7_75t_L g247 ( .A(n_204), .B(n_220), .Y(n_247) );
AND2x2_ASAP7_75t_L g323 ( .A(n_204), .B(n_270), .Y(n_323) );
NAND2xp5_ASAP7_75t_L g363 ( .A(n_204), .B(n_229), .Y(n_363) );
OA21x2_ASAP7_75t_L g204 ( .A1(n_205), .A2(n_206), .B(n_218), .Y(n_204) );
OA21x2_ASAP7_75t_L g229 ( .A1(n_205), .A2(n_230), .B(n_237), .Y(n_229) );
O2A1O1Ixp33_ASAP7_75t_L g207 ( .A1(n_208), .A2(n_209), .B(n_210), .C(n_211), .Y(n_207) );
AOI21xp5_ASAP7_75t_L g486 ( .A1(n_209), .A2(n_487), .B(n_488), .Y(n_486) );
AOI21xp5_ASAP7_75t_L g497 ( .A1(n_209), .A2(n_498), .B(n_499), .Y(n_497) );
O2A1O1Ixp33_ASAP7_75t_L g426 ( .A1(n_211), .A2(n_427), .B(n_428), .C(n_429), .Y(n_426) );
AOI21xp5_ASAP7_75t_L g471 ( .A1(n_213), .A2(n_472), .B(n_473), .Y(n_471) );
INVx2_ASAP7_75t_L g213 ( .A(n_214), .Y(n_213) );
INVx1_ASAP7_75t_L g214 ( .A(n_215), .Y(n_214) );
NAND2xp5_ASAP7_75t_L g265 ( .A(n_219), .B(n_266), .Y(n_265) );
AND2x2_ASAP7_75t_L g279 ( .A(n_219), .B(n_240), .Y(n_279) );
AND2x2_ASAP7_75t_L g283 ( .A(n_219), .B(n_273), .Y(n_283) );
AND2x2_ASAP7_75t_L g219 ( .A(n_220), .B(n_229), .Y(n_219) );
INVx3_ASAP7_75t_L g244 ( .A(n_220), .Y(n_244) );
AND2x2_ASAP7_75t_L g269 ( .A(n_220), .B(n_270), .Y(n_269) );
AND2x2_ASAP7_75t_L g404 ( .A(n_220), .B(n_387), .Y(n_404) );
HB1xp67_ASAP7_75t_L g258 ( .A(n_229), .Y(n_258) );
INVx2_ASAP7_75t_L g270 ( .A(n_229), .Y(n_270) );
AND2x2_ASAP7_75t_L g314 ( .A(n_229), .B(n_290), .Y(n_314) );
INVx1_ASAP7_75t_L g357 ( .A(n_229), .Y(n_357) );
OR2x2_ASAP7_75t_L g388 ( .A(n_229), .B(n_290), .Y(n_388) );
AND2x2_ASAP7_75t_L g408 ( .A(n_229), .B(n_244), .Y(n_408) );
OAI21xp5_ASAP7_75t_L g238 ( .A1(n_239), .A2(n_241), .B(n_245), .Y(n_238) );
INVx1_ASAP7_75t_L g239 ( .A(n_240), .Y(n_239) );
AND2x2_ASAP7_75t_L g246 ( .A(n_240), .B(n_247), .Y(n_246) );
NAND2xp5_ASAP7_75t_L g373 ( .A(n_240), .B(n_374), .Y(n_373) );
INVx1_ASAP7_75t_L g365 ( .A(n_242), .Y(n_365) );
INVx2_ASAP7_75t_SL g259 ( .A(n_243), .Y(n_259) );
AND2x2_ASAP7_75t_L g379 ( .A(n_243), .B(n_273), .Y(n_379) );
INVx2_ASAP7_75t_L g325 ( .A(n_244), .Y(n_325) );
NAND2xp5_ASAP7_75t_L g356 ( .A(n_244), .B(n_357), .Y(n_356) );
AOI22xp5_ASAP7_75t_L g245 ( .A1(n_246), .A2(n_248), .B1(n_251), .B2(n_257), .Y(n_245) );
NAND2xp5_ASAP7_75t_L g391 ( .A(n_247), .B(n_392), .Y(n_391) );
INVx1_ASAP7_75t_SL g413 ( .A(n_247), .Y(n_413) );
AND2x2_ASAP7_75t_L g248 ( .A(n_249), .B(n_250), .Y(n_248) );
INVx1_ASAP7_75t_L g338 ( .A(n_249), .Y(n_338) );
NAND2xp5_ASAP7_75t_L g350 ( .A(n_249), .B(n_281), .Y(n_350) );
NOR2xp33_ASAP7_75t_L g337 ( .A(n_250), .B(n_338), .Y(n_337) );
AND2x2_ASAP7_75t_L g354 ( .A(n_250), .B(n_303), .Y(n_354) );
INVx2_ASAP7_75t_L g410 ( .A(n_250), .Y(n_410) );
INVx1_ASAP7_75t_L g251 ( .A(n_252), .Y(n_251) );
NAND2xp5_ASAP7_75t_L g252 ( .A(n_253), .B(n_254), .Y(n_252) );
AND2x2_ASAP7_75t_L g280 ( .A(n_253), .B(n_281), .Y(n_280) );
NAND2xp5_ASAP7_75t_L g331 ( .A(n_253), .B(n_298), .Y(n_331) );
INVx2_ASAP7_75t_L g254 ( .A(n_255), .Y(n_254) );
NOR2xp33_ASAP7_75t_L g333 ( .A(n_255), .B(n_275), .Y(n_333) );
NOR2xp33_ASAP7_75t_L g257 ( .A(n_258), .B(n_259), .Y(n_257) );
INVx1_ASAP7_75t_L g392 ( .A(n_258), .Y(n_392) );
O2A1O1Ixp33_ASAP7_75t_SL g342 ( .A1(n_259), .A2(n_343), .B(n_345), .C(n_348), .Y(n_342) );
OR2x2_ASAP7_75t_L g369 ( .A(n_259), .B(n_273), .Y(n_369) );
OAI221xp5_ASAP7_75t_SL g260 ( .A1(n_261), .A2(n_265), .B1(n_267), .B2(n_274), .C(n_277), .Y(n_260) );
NAND2xp5_ASAP7_75t_SL g261 ( .A(n_262), .B(n_264), .Y(n_261) );
NAND2xp5_ASAP7_75t_L g318 ( .A(n_262), .B(n_311), .Y(n_318) );
AND2x2_ASAP7_75t_L g360 ( .A(n_262), .B(n_361), .Y(n_360) );
INVx2_ASAP7_75t_L g396 ( .A(n_262), .Y(n_396) );
HB1xp67_ASAP7_75t_L g287 ( .A(n_263), .Y(n_287) );
INVx1_ASAP7_75t_L g300 ( .A(n_263), .Y(n_300) );
NOR2xp67_ASAP7_75t_L g320 ( .A(n_266), .B(n_321), .Y(n_320) );
INVxp67_ASAP7_75t_L g374 ( .A(n_266), .Y(n_374) );
NAND2xp5_ASAP7_75t_SL g390 ( .A(n_266), .B(n_314), .Y(n_390) );
INVx2_ASAP7_75t_L g376 ( .A(n_267), .Y(n_376) );
OR2x2_ASAP7_75t_L g267 ( .A(n_268), .B(n_271), .Y(n_267) );
INVx1_ASAP7_75t_L g268 ( .A(n_269), .Y(n_268) );
AND2x2_ASAP7_75t_L g317 ( .A(n_269), .B(n_288), .Y(n_317) );
O2A1O1Ixp33_ASAP7_75t_L g326 ( .A1(n_269), .A2(n_285), .B(n_327), .C(n_328), .Y(n_326) );
AND2x2_ASAP7_75t_L g295 ( .A(n_270), .B(n_290), .Y(n_295) );
INVx1_ASAP7_75t_L g271 ( .A(n_272), .Y(n_271) );
NOR2xp33_ASAP7_75t_L g372 ( .A(n_274), .B(n_373), .Y(n_372) );
OR2x2_ASAP7_75t_L g274 ( .A(n_275), .B(n_276), .Y(n_274) );
OR2x2_ASAP7_75t_L g343 ( .A(n_275), .B(n_344), .Y(n_343) );
AOI22xp5_ASAP7_75t_L g277 ( .A1(n_278), .A2(n_279), .B1(n_280), .B2(n_283), .Y(n_277) );
INVx1_ASAP7_75t_L g397 ( .A(n_279), .Y(n_397) );
INVx1_ASAP7_75t_L g344 ( .A(n_281), .Y(n_344) );
INVx1_ASAP7_75t_L g395 ( .A(n_283), .Y(n_395) );
AOI211xp5_ASAP7_75t_SL g284 ( .A1(n_285), .A2(n_288), .B(n_292), .C(n_315), .Y(n_284) );
INVx1_ASAP7_75t_L g285 ( .A(n_286), .Y(n_285) );
OR2x2_ASAP7_75t_L g307 ( .A(n_287), .B(n_308), .Y(n_307) );
INVx1_ASAP7_75t_L g358 ( .A(n_288), .Y(n_358) );
AND2x2_ASAP7_75t_L g407 ( .A(n_288), .B(n_408), .Y(n_407) );
INVx1_ASAP7_75t_L g289 ( .A(n_290), .Y(n_289) );
OAI21xp33_ASAP7_75t_L g292 ( .A1(n_293), .A2(n_297), .B(n_305), .Y(n_292) );
INVx1_ASAP7_75t_SL g293 ( .A(n_294), .Y(n_293) );
AND2x2_ASAP7_75t_L g294 ( .A(n_295), .B(n_296), .Y(n_294) );
INVx2_ASAP7_75t_L g321 ( .A(n_295), .Y(n_321) );
NAND2xp5_ASAP7_75t_L g340 ( .A(n_295), .B(n_341), .Y(n_340) );
AND2x2_ASAP7_75t_L g313 ( .A(n_296), .B(n_314), .Y(n_313) );
INVx2_ASAP7_75t_L g389 ( .A(n_296), .Y(n_389) );
OAI32xp33_ASAP7_75t_L g400 ( .A1(n_296), .A2(n_348), .A3(n_355), .B1(n_396), .B2(n_401), .Y(n_400) );
NOR2xp33_ASAP7_75t_SL g297 ( .A(n_298), .B(n_301), .Y(n_297) );
INVx1_ASAP7_75t_SL g368 ( .A(n_298), .Y(n_368) );
AND2x2_ASAP7_75t_L g301 ( .A(n_302), .B(n_304), .Y(n_301) );
INVx1_ASAP7_75t_L g302 ( .A(n_303), .Y(n_302) );
INVx1_ASAP7_75t_SL g308 ( .A(n_304), .Y(n_308) );
OAI21xp33_ASAP7_75t_L g305 ( .A1(n_306), .A2(n_309), .B(n_313), .Y(n_305) );
INVx1_ASAP7_75t_L g306 ( .A(n_307), .Y(n_306) );
OAI22xp33_ASAP7_75t_L g380 ( .A1(n_307), .A2(n_355), .B1(n_381), .B2(n_383), .Y(n_380) );
INVx1_ASAP7_75t_L g309 ( .A(n_310), .Y(n_309) );
OR2x2_ASAP7_75t_L g310 ( .A(n_311), .B(n_312), .Y(n_310) );
NAND2xp5_ASAP7_75t_L g383 ( .A(n_311), .B(n_384), .Y(n_383) );
INVx1_ASAP7_75t_L g348 ( .A(n_314), .Y(n_348) );
INVx1_ASAP7_75t_L g316 ( .A(n_317), .Y(n_316) );
INVx1_ASAP7_75t_L g319 ( .A(n_320), .Y(n_319) );
NAND2x1p5_ASAP7_75t_L g322 ( .A(n_323), .B(n_324), .Y(n_322) );
INVx1_ASAP7_75t_L g341 ( .A(n_325), .Y(n_341) );
OAI21xp5_ASAP7_75t_L g328 ( .A1(n_329), .A2(n_331), .B(n_332), .Y(n_328) );
INVx1_ASAP7_75t_L g329 ( .A(n_330), .Y(n_329) );
AOI221xp5_ASAP7_75t_L g375 ( .A1(n_334), .A2(n_376), .B1(n_377), .B2(n_379), .C(n_380), .Y(n_375) );
NAND5xp2_ASAP7_75t_L g335 ( .A(n_336), .B(n_359), .C(n_375), .D(n_385), .E(n_403), .Y(n_335) );
AOI211xp5_ASAP7_75t_SL g336 ( .A1(n_337), .A2(n_339), .B(n_342), .C(n_349), .Y(n_336) );
INVx1_ASAP7_75t_L g339 ( .A(n_340), .Y(n_339) );
INVx1_ASAP7_75t_L g406 ( .A(n_343), .Y(n_406) );
NAND2xp5_ASAP7_75t_L g345 ( .A(n_346), .B(n_347), .Y(n_345) );
OAI22xp33_ASAP7_75t_L g349 ( .A1(n_350), .A2(n_351), .B1(n_353), .B2(n_355), .Y(n_349) );
INVx1_ASAP7_75t_SL g382 ( .A(n_352), .Y(n_382) );
INVx1_ASAP7_75t_L g353 ( .A(n_354), .Y(n_353) );
OAI322xp33_ASAP7_75t_L g364 ( .A1(n_355), .A2(n_365), .A3(n_366), .B1(n_367), .B2(n_368), .C1(n_369), .C2(n_370), .Y(n_364) );
OR2x2_ASAP7_75t_L g355 ( .A(n_356), .B(n_358), .Y(n_355) );
INVx1_ASAP7_75t_L g367 ( .A(n_357), .Y(n_367) );
NAND2xp5_ASAP7_75t_L g381 ( .A(n_357), .B(n_382), .Y(n_381) );
AOI211xp5_ASAP7_75t_SL g359 ( .A1(n_360), .A2(n_362), .B(n_364), .C(n_372), .Y(n_359) );
INVx1_ASAP7_75t_L g362 ( .A(n_363), .Y(n_362) );
OAI22xp33_ASAP7_75t_L g394 ( .A1(n_368), .A2(n_395), .B1(n_396), .B2(n_397), .Y(n_394) );
INVx1_ASAP7_75t_SL g370 ( .A(n_371), .Y(n_370) );
INVx1_ASAP7_75t_L g411 ( .A(n_378), .Y(n_411) );
AOI221xp5_ASAP7_75t_L g385 ( .A1(n_386), .A2(n_393), .B1(n_394), .B2(n_398), .C(n_400), .Y(n_385) );
OAI211xp5_ASAP7_75t_SL g386 ( .A1(n_387), .A2(n_389), .B(n_390), .C(n_391), .Y(n_386) );
INVx1_ASAP7_75t_SL g387 ( .A(n_388), .Y(n_387) );
OR2x2_ASAP7_75t_L g412 ( .A(n_388), .B(n_413), .Y(n_412) );
INVx1_ASAP7_75t_L g398 ( .A(n_399), .Y(n_398) );
AOI221xp5_ASAP7_75t_L g403 ( .A1(n_404), .A2(n_405), .B1(n_406), .B2(n_407), .C(n_409), .Y(n_403) );
AOI21xp33_ASAP7_75t_SL g409 ( .A1(n_410), .A2(n_411), .B(n_412), .Y(n_409) );
NAND2x1p5_ASAP7_75t_L g416 ( .A(n_417), .B(n_618), .Y(n_416) );
AND4x1_ASAP7_75t_L g417 ( .A(n_418), .B(n_558), .C(n_573), .D(n_598), .Y(n_417) );
NOR2xp33_ASAP7_75t_SL g418 ( .A(n_419), .B(n_531), .Y(n_418) );
OAI21xp33_ASAP7_75t_L g419 ( .A1(n_420), .A2(n_449), .B(n_511), .Y(n_419) );
AND2x2_ASAP7_75t_L g561 ( .A(n_420), .B(n_466), .Y(n_561) );
AND2x2_ASAP7_75t_L g574 ( .A(n_420), .B(n_465), .Y(n_574) );
NAND2xp5_ASAP7_75t_L g624 ( .A(n_420), .B(n_450), .Y(n_624) );
INVx1_ASAP7_75t_L g628 ( .A(n_420), .Y(n_628) );
AND2x2_ASAP7_75t_L g420 ( .A(n_421), .B(n_437), .Y(n_420) );
INVx2_ASAP7_75t_L g545 ( .A(n_421), .Y(n_545) );
BUFx2_ASAP7_75t_L g572 ( .A(n_421), .Y(n_572) );
NAND2xp5_ASAP7_75t_L g422 ( .A(n_423), .B(n_432), .Y(n_422) );
INVx5_ASAP7_75t_L g442 ( .A(n_424), .Y(n_442) );
INVx1_ASAP7_75t_L g430 ( .A(n_431), .Y(n_430) );
O2A1O1Ixp33_ASAP7_75t_SL g440 ( .A1(n_431), .A2(n_441), .B(n_442), .C(n_443), .Y(n_440) );
O2A1O1Ixp33_ASAP7_75t_L g521 ( .A1(n_431), .A2(n_442), .B(n_522), .C(n_523), .Y(n_521) );
BUFx2_ASAP7_75t_L g469 ( .A(n_433), .Y(n_469) );
AND2x2_ASAP7_75t_L g512 ( .A(n_437), .B(n_466), .Y(n_512) );
INVx2_ASAP7_75t_L g528 ( .A(n_437), .Y(n_528) );
AND2x2_ASAP7_75t_L g537 ( .A(n_437), .B(n_465), .Y(n_537) );
AND2x2_ASAP7_75t_L g616 ( .A(n_437), .B(n_545), .Y(n_616) );
OA21x2_ASAP7_75t_L g437 ( .A1(n_438), .A2(n_439), .B(n_448), .Y(n_437) );
INVx2_ASAP7_75t_L g456 ( .A(n_442), .Y(n_456) );
NOR2xp33_ASAP7_75t_L g444 ( .A(n_445), .B(n_446), .Y(n_444) );
NAND2xp5_ASAP7_75t_L g449 ( .A(n_450), .B(n_478), .Y(n_449) );
NAND2xp5_ASAP7_75t_L g581 ( .A(n_450), .B(n_543), .Y(n_581) );
INVx1_ASAP7_75t_L g669 ( .A(n_450), .Y(n_669) );
AND2x2_ASAP7_75t_L g450 ( .A(n_451), .B(n_465), .Y(n_450) );
AND2x2_ASAP7_75t_L g527 ( .A(n_451), .B(n_528), .Y(n_527) );
OR2x2_ASAP7_75t_L g541 ( .A(n_451), .B(n_542), .Y(n_541) );
HB1xp67_ASAP7_75t_L g570 ( .A(n_451), .Y(n_570) );
OR2x2_ASAP7_75t_L g602 ( .A(n_451), .B(n_544), .Y(n_602) );
AND2x2_ASAP7_75t_L g610 ( .A(n_451), .B(n_611), .Y(n_610) );
AND2x2_ASAP7_75t_L g643 ( .A(n_451), .B(n_612), .Y(n_643) );
NAND2xp5_ASAP7_75t_L g660 ( .A(n_451), .B(n_512), .Y(n_660) );
NAND2xp5_ASAP7_75t_L g668 ( .A(n_451), .B(n_572), .Y(n_668) );
AND2x2_ASAP7_75t_L g674 ( .A(n_451), .B(n_561), .Y(n_674) );
INVx5_ASAP7_75t_L g451 ( .A(n_452), .Y(n_451) );
BUFx2_ASAP7_75t_L g534 ( .A(n_452), .Y(n_534) );
AND2x2_ASAP7_75t_L g564 ( .A(n_452), .B(n_544), .Y(n_564) );
AND2x2_ASAP7_75t_L g597 ( .A(n_452), .B(n_557), .Y(n_597) );
AND2x2_ASAP7_75t_L g617 ( .A(n_452), .B(n_466), .Y(n_617) );
AND2x2_ASAP7_75t_L g651 ( .A(n_452), .B(n_517), .Y(n_651) );
OR2x6_ASAP7_75t_L g452 ( .A(n_453), .B(n_463), .Y(n_452) );
O2A1O1Ixp33_ASAP7_75t_L g457 ( .A1(n_458), .A2(n_459), .B(n_461), .C(n_462), .Y(n_457) );
O2A1O1Ixp33_ASAP7_75t_L g507 ( .A1(n_459), .A2(n_462), .B(n_508), .C(n_509), .Y(n_507) );
INVx2_ASAP7_75t_L g459 ( .A(n_460), .Y(n_459) );
AND2x4_ASAP7_75t_L g557 ( .A(n_465), .B(n_528), .Y(n_557) );
AND2x2_ASAP7_75t_L g568 ( .A(n_465), .B(n_564), .Y(n_568) );
NAND2xp5_ASAP7_75t_L g607 ( .A(n_465), .B(n_544), .Y(n_607) );
INVx2_ASAP7_75t_L g622 ( .A(n_465), .Y(n_622) );
NOR2xp33_ASAP7_75t_L g645 ( .A(n_465), .B(n_556), .Y(n_645) );
AND2x2_ASAP7_75t_L g664 ( .A(n_465), .B(n_616), .Y(n_664) );
INVx5_ASAP7_75t_L g465 ( .A(n_466), .Y(n_465) );
HB1xp67_ASAP7_75t_L g563 ( .A(n_466), .Y(n_563) );
AND2x2_ASAP7_75t_L g571 ( .A(n_466), .B(n_572), .Y(n_571) );
AND2x4_ASAP7_75t_L g612 ( .A(n_466), .B(n_528), .Y(n_612) );
OR2x6_ASAP7_75t_L g466 ( .A(n_467), .B(n_475), .Y(n_466) );
AOI21xp5_ASAP7_75t_SL g467 ( .A1(n_468), .A2(n_470), .B(n_474), .Y(n_467) );
NOR2xp33_ASAP7_75t_L g475 ( .A(n_476), .B(n_477), .Y(n_475) );
INVx1_ASAP7_75t_L g478 ( .A(n_479), .Y(n_478) );
NAND2xp5_ASAP7_75t_L g479 ( .A(n_480), .B(n_489), .Y(n_479) );
AND2x2_ASAP7_75t_L g535 ( .A(n_480), .B(n_518), .Y(n_535) );
INVx1_ASAP7_75t_SL g480 ( .A(n_481), .Y(n_480) );
NAND2xp5_ASAP7_75t_SL g515 ( .A(n_481), .B(n_492), .Y(n_515) );
OR2x2_ASAP7_75t_L g548 ( .A(n_481), .B(n_518), .Y(n_548) );
NAND2xp5_ASAP7_75t_L g553 ( .A(n_481), .B(n_518), .Y(n_553) );
AND2x2_ASAP7_75t_L g580 ( .A(n_481), .B(n_517), .Y(n_580) );
AND2x2_ASAP7_75t_L g632 ( .A(n_481), .B(n_491), .Y(n_632) );
INVx2_ASAP7_75t_L g481 ( .A(n_482), .Y(n_481) );
NAND2xp5_ASAP7_75t_L g540 ( .A(n_482), .B(n_502), .Y(n_540) );
AND2x2_ASAP7_75t_L g576 ( .A(n_482), .B(n_492), .Y(n_576) );
NAND2xp5_ASAP7_75t_L g639 ( .A(n_489), .B(n_640), .Y(n_639) );
INVx2_ASAP7_75t_L g489 ( .A(n_490), .Y(n_489) );
OR2x2_ASAP7_75t_L g566 ( .A(n_490), .B(n_548), .Y(n_566) );
OR2x2_ASAP7_75t_L g490 ( .A(n_491), .B(n_502), .Y(n_490) );
OAI322xp33_ASAP7_75t_L g531 ( .A1(n_491), .A2(n_532), .A3(n_536), .B1(n_538), .B2(n_541), .C1(n_546), .C2(n_554), .Y(n_531) );
NAND2xp5_ASAP7_75t_L g539 ( .A(n_491), .B(n_517), .Y(n_539) );
OR2x2_ASAP7_75t_L g549 ( .A(n_491), .B(n_503), .Y(n_549) );
AND2x2_ASAP7_75t_L g551 ( .A(n_491), .B(n_503), .Y(n_551) );
NOR2xp33_ASAP7_75t_L g552 ( .A(n_491), .B(n_553), .Y(n_552) );
NAND2xp5_ASAP7_75t_L g613 ( .A(n_491), .B(n_518), .Y(n_613) );
NOR2xp33_ASAP7_75t_L g646 ( .A(n_491), .B(n_647), .Y(n_646) );
INVx5_ASAP7_75t_SL g491 ( .A(n_492), .Y(n_491) );
NAND2xp5_ASAP7_75t_L g661 ( .A(n_492), .B(n_535), .Y(n_661) );
OAI21xp5_ASAP7_75t_L g493 ( .A1(n_494), .A2(n_495), .B(n_496), .Y(n_493) );
NAND2xp5_ASAP7_75t_L g516 ( .A(n_502), .B(n_517), .Y(n_516) );
AND2x2_ASAP7_75t_L g529 ( .A(n_502), .B(n_530), .Y(n_529) );
NAND2xp5_ASAP7_75t_L g579 ( .A(n_502), .B(n_580), .Y(n_579) );
OR2x2_ASAP7_75t_L g591 ( .A(n_502), .B(n_518), .Y(n_591) );
AOI211xp5_ASAP7_75t_SL g619 ( .A1(n_502), .A2(n_620), .B(n_623), .C(n_635), .Y(n_619) );
NAND2xp5_ASAP7_75t_L g625 ( .A(n_502), .B(n_626), .Y(n_625) );
AND2x2_ASAP7_75t_L g657 ( .A(n_502), .B(n_632), .Y(n_657) );
INVx5_ASAP7_75t_SL g502 ( .A(n_503), .Y(n_502) );
AND2x2_ASAP7_75t_L g585 ( .A(n_503), .B(n_518), .Y(n_585) );
HB1xp67_ASAP7_75t_L g594 ( .A(n_503), .Y(n_594) );
AND2x2_ASAP7_75t_L g634 ( .A(n_503), .B(n_632), .Y(n_634) );
AND2x2_ASAP7_75t_SL g665 ( .A(n_503), .B(n_535), .Y(n_665) );
AND2x2_ASAP7_75t_L g672 ( .A(n_503), .B(n_631), .Y(n_672) );
OR2x6_ASAP7_75t_L g503 ( .A(n_504), .B(n_510), .Y(n_503) );
AOI22xp33_ASAP7_75t_L g511 ( .A1(n_512), .A2(n_513), .B1(n_527), .B2(n_529), .Y(n_511) );
NAND2xp5_ASAP7_75t_L g582 ( .A(n_512), .B(n_534), .Y(n_582) );
INVx2_ASAP7_75t_L g513 ( .A(n_514), .Y(n_513) );
OR2x2_ASAP7_75t_L g514 ( .A(n_515), .B(n_516), .Y(n_514) );
INVx1_ASAP7_75t_L g530 ( .A(n_515), .Y(n_530) );
OR2x2_ASAP7_75t_L g590 ( .A(n_515), .B(n_591), .Y(n_590) );
OAI221xp5_ASAP7_75t_SL g638 ( .A1(n_515), .A2(n_639), .B1(n_641), .B2(n_642), .C(n_644), .Y(n_638) );
INVx2_ASAP7_75t_L g577 ( .A(n_516), .Y(n_577) );
AND2x2_ASAP7_75t_L g550 ( .A(n_517), .B(n_551), .Y(n_550) );
INVx1_ASAP7_75t_L g640 ( .A(n_517), .Y(n_640) );
NAND2xp5_ASAP7_75t_L g653 ( .A(n_517), .B(n_632), .Y(n_653) );
INVx3_ASAP7_75t_L g517 ( .A(n_518), .Y(n_517) );
INVxp67_ASAP7_75t_L g595 ( .A(n_518), .Y(n_595) );
AND2x2_ASAP7_75t_L g631 ( .A(n_518), .B(n_632), .Y(n_631) );
OA21x2_ASAP7_75t_L g518 ( .A1(n_519), .A2(n_520), .B(n_526), .Y(n_518) );
AND2x2_ASAP7_75t_L g633 ( .A(n_527), .B(n_572), .Y(n_633) );
AND2x2_ASAP7_75t_L g543 ( .A(n_528), .B(n_544), .Y(n_543) );
NAND2xp5_ASAP7_75t_L g600 ( .A(n_528), .B(n_601), .Y(n_600) );
NOR2xp33_ASAP7_75t_SL g614 ( .A(n_530), .B(n_577), .Y(n_614) );
INVx1_ASAP7_75t_SL g532 ( .A(n_533), .Y(n_532) );
AND2x2_ASAP7_75t_L g620 ( .A(n_533), .B(n_621), .Y(n_620) );
AND2x2_ASAP7_75t_L g533 ( .A(n_534), .B(n_535), .Y(n_533) );
OR2x2_ASAP7_75t_L g606 ( .A(n_534), .B(n_607), .Y(n_606) );
AND2x2_ASAP7_75t_L g671 ( .A(n_534), .B(n_616), .Y(n_671) );
INVx2_ASAP7_75t_L g604 ( .A(n_535), .Y(n_604) );
NAND4xp25_ASAP7_75t_SL g667 ( .A(n_536), .B(n_668), .C(n_669), .D(n_670), .Y(n_667) );
INVx1_ASAP7_75t_L g536 ( .A(n_537), .Y(n_536) );
NAND2xp5_ASAP7_75t_L g636 ( .A(n_537), .B(n_601), .Y(n_636) );
OR2x2_ASAP7_75t_L g538 ( .A(n_539), .B(n_540), .Y(n_538) );
INVx1_ASAP7_75t_SL g673 ( .A(n_540), .Y(n_673) );
O2A1O1Ixp33_ASAP7_75t_SL g635 ( .A1(n_541), .A2(n_604), .B(n_608), .C(n_636), .Y(n_635) );
INVx1_ASAP7_75t_L g542 ( .A(n_543), .Y(n_542) );
AND2x2_ASAP7_75t_L g630 ( .A(n_543), .B(n_622), .Y(n_630) );
HB1xp67_ASAP7_75t_L g556 ( .A(n_544), .Y(n_556) );
INVx1_ASAP7_75t_L g611 ( .A(n_544), .Y(n_611) );
INVx2_ASAP7_75t_L g544 ( .A(n_545), .Y(n_544) );
HB1xp67_ASAP7_75t_L g588 ( .A(n_545), .Y(n_588) );
AOI211xp5_ASAP7_75t_L g546 ( .A1(n_547), .A2(n_549), .B(n_550), .C(n_552), .Y(n_546) );
AND2x2_ASAP7_75t_L g567 ( .A(n_547), .B(n_551), .Y(n_567) );
OAI322xp33_ASAP7_75t_SL g605 ( .A1(n_547), .A2(n_606), .A3(n_608), .B1(n_609), .B2(n_613), .C1(n_614), .C2(n_615), .Y(n_605) );
INVx1_ASAP7_75t_SL g547 ( .A(n_548), .Y(n_547) );
OR2x2_ASAP7_75t_L g627 ( .A(n_549), .B(n_553), .Y(n_627) );
INVx1_ASAP7_75t_L g608 ( .A(n_551), .Y(n_608) );
INVx1_ASAP7_75t_SL g626 ( .A(n_553), .Y(n_626) );
INVx2_ASAP7_75t_L g554 ( .A(n_555), .Y(n_554) );
AND2x2_ASAP7_75t_L g555 ( .A(n_556), .B(n_557), .Y(n_555) );
AOI222xp33_ASAP7_75t_L g558 ( .A1(n_559), .A2(n_565), .B1(n_567), .B2(n_568), .C1(n_569), .C2(n_714), .Y(n_558) );
NAND2xp5_ASAP7_75t_SL g559 ( .A(n_560), .B(n_562), .Y(n_559) );
OAI322xp33_ASAP7_75t_L g648 ( .A1(n_560), .A2(n_622), .A3(n_627), .B1(n_649), .B2(n_650), .C1(n_652), .C2(n_653), .Y(n_648) );
INVx1_ASAP7_75t_L g560 ( .A(n_561), .Y(n_560) );
AOI221xp5_ASAP7_75t_L g598 ( .A1(n_561), .A2(n_575), .B1(n_599), .B2(n_603), .C(n_605), .Y(n_598) );
NAND2xp5_ASAP7_75t_L g562 ( .A(n_563), .B(n_564), .Y(n_562) );
INVx1_ASAP7_75t_SL g565 ( .A(n_566), .Y(n_565) );
OAI222xp33_ASAP7_75t_L g578 ( .A1(n_566), .A2(n_579), .B1(n_581), .B2(n_582), .C1(n_583), .C2(n_586), .Y(n_578) );
AOI22xp5_ASAP7_75t_L g644 ( .A1(n_568), .A2(n_575), .B1(n_645), .B2(n_646), .Y(n_644) );
AND2x2_ASAP7_75t_L g569 ( .A(n_570), .B(n_571), .Y(n_569) );
AOI211xp5_ASAP7_75t_L g573 ( .A1(n_574), .A2(n_575), .B(n_578), .C(n_589), .Y(n_573) );
O2A1O1Ixp33_ASAP7_75t_L g654 ( .A1(n_575), .A2(n_612), .B(n_655), .C(n_658), .Y(n_654) );
AND2x4_ASAP7_75t_L g575 ( .A(n_576), .B(n_577), .Y(n_575) );
AND2x2_ASAP7_75t_L g584 ( .A(n_576), .B(n_585), .Y(n_584) );
INVx1_ASAP7_75t_SL g647 ( .A(n_580), .Y(n_647) );
INVx1_ASAP7_75t_L g583 ( .A(n_584), .Y(n_583) );
INVx1_ASAP7_75t_L g586 ( .A(n_587), .Y(n_586) );
NAND2xp5_ASAP7_75t_L g641 ( .A(n_587), .B(n_612), .Y(n_641) );
BUFx2_ASAP7_75t_L g587 ( .A(n_588), .Y(n_587) );
AOI21xp33_ASAP7_75t_L g589 ( .A1(n_590), .A2(n_592), .B(n_596), .Y(n_589) );
OAI221xp5_ASAP7_75t_SL g658 ( .A1(n_590), .A2(n_659), .B1(n_660), .B2(n_661), .C(n_662), .Y(n_658) );
INVxp33_ASAP7_75t_L g592 ( .A(n_593), .Y(n_592) );
NOR2xp33_ASAP7_75t_L g593 ( .A(n_594), .B(n_595), .Y(n_593) );
NOR2xp33_ASAP7_75t_L g603 ( .A(n_594), .B(n_604), .Y(n_603) );
INVx1_ASAP7_75t_L g596 ( .A(n_597), .Y(n_596) );
INVx1_ASAP7_75t_L g599 ( .A(n_600), .Y(n_599) );
NAND2xp5_ASAP7_75t_L g652 ( .A(n_601), .B(n_612), .Y(n_652) );
INVx2_ASAP7_75t_SL g601 ( .A(n_602), .Y(n_601) );
NAND2xp5_ASAP7_75t_L g609 ( .A(n_610), .B(n_612), .Y(n_609) );
NAND2xp5_ASAP7_75t_L g615 ( .A(n_616), .B(n_617), .Y(n_615) );
AND2x2_ASAP7_75t_L g663 ( .A(n_616), .B(n_622), .Y(n_663) );
AND4x1_ASAP7_75t_L g618 ( .A(n_619), .B(n_637), .C(n_654), .D(n_666), .Y(n_618) );
INVx1_ASAP7_75t_L g621 ( .A(n_622), .Y(n_621) );
OAI221xp5_ASAP7_75t_SL g623 ( .A1(n_624), .A2(n_625), .B1(n_627), .B2(n_628), .C(n_629), .Y(n_623) );
AOI22xp5_ASAP7_75t_L g629 ( .A1(n_630), .A2(n_631), .B1(n_633), .B2(n_634), .Y(n_629) );
INVx1_ASAP7_75t_L g659 ( .A(n_630), .Y(n_659) );
INVx1_ASAP7_75t_SL g649 ( .A(n_634), .Y(n_649) );
NOR2xp33_ASAP7_75t_SL g637 ( .A(n_638), .B(n_648), .Y(n_637) );
INVx1_ASAP7_75t_L g642 ( .A(n_643), .Y(n_642) );
NOR2xp33_ASAP7_75t_L g655 ( .A(n_650), .B(n_656), .Y(n_655) );
INVx1_ASAP7_75t_L g650 ( .A(n_651), .Y(n_650) );
INVx1_ASAP7_75t_L g656 ( .A(n_657), .Y(n_656) );
AOI22xp33_ASAP7_75t_L g662 ( .A1(n_657), .A2(n_663), .B1(n_664), .B2(n_665), .Y(n_662) );
AOI22xp5_ASAP7_75t_L g666 ( .A1(n_667), .A2(n_672), .B1(n_673), .B2(n_674), .Y(n_666) );
INVx1_ASAP7_75t_L g670 ( .A(n_671), .Y(n_670) );
INVx2_ASAP7_75t_L g676 ( .A(n_677), .Y(n_676) );
AND2x2_ASAP7_75t_L g677 ( .A(n_678), .B(n_679), .Y(n_677) );
INVx1_ASAP7_75t_SL g680 ( .A(n_681), .Y(n_680) );
INVx3_ASAP7_75t_SL g681 ( .A(n_682), .Y(n_681) );
INVx1_ASAP7_75t_L g683 ( .A(n_684), .Y(n_683) );
NAND2xp33_ASAP7_75t_L g684 ( .A(n_685), .B(n_689), .Y(n_684) );
NOR2xp33_ASAP7_75t_SL g685 ( .A(n_686), .B(n_688), .Y(n_685) );
INVx1_ASAP7_75t_SL g709 ( .A(n_686), .Y(n_709) );
INVx1_ASAP7_75t_L g708 ( .A(n_688), .Y(n_708) );
OA21x2_ASAP7_75t_L g711 ( .A1(n_688), .A2(n_709), .B(n_712), .Y(n_711) );
INVx1_ASAP7_75t_SL g689 ( .A(n_690), .Y(n_689) );
INVx1_ASAP7_75t_SL g690 ( .A(n_691), .Y(n_690) );
HB1xp67_ASAP7_75t_L g699 ( .A(n_691), .Y(n_699) );
INVx2_ASAP7_75t_L g703 ( .A(n_691), .Y(n_703) );
BUFx2_ASAP7_75t_L g712 ( .A(n_691), .Y(n_712) );
INVxp67_ASAP7_75t_L g692 ( .A(n_693), .Y(n_692) );
AOI21xp5_ASAP7_75t_L g693 ( .A1(n_694), .A2(n_699), .B(n_700), .Y(n_693) );
HB1xp67_ASAP7_75t_L g694 ( .A(n_695), .Y(n_694) );
INVx1_ASAP7_75t_L g696 ( .A(n_697), .Y(n_696) );
NOR2xp33_ASAP7_75t_L g700 ( .A(n_701), .B(n_702), .Y(n_700) );
INVx1_ASAP7_75t_L g702 ( .A(n_703), .Y(n_702) );
INVx1_ASAP7_75t_SL g704 ( .A(n_705), .Y(n_704) );
CKINVDCx6p67_ASAP7_75t_R g705 ( .A(n_706), .Y(n_705) );
AND2x2_ASAP7_75t_L g706 ( .A(n_707), .B(n_709), .Y(n_706) );
INVx1_ASAP7_75t_L g707 ( .A(n_708), .Y(n_707) );
INVx2_ASAP7_75t_SL g710 ( .A(n_711), .Y(n_710) );
endmodule