module fake_jpeg_28851_n_39 (n_11, n_3, n_2, n_1, n_0, n_10, n_4, n_8, n_9, n_6, n_5, n_7, n_39);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_39;

wire n_13;
wire n_21;
wire n_33;
wire n_23;
wire n_27;
wire n_22;
wire n_14;
wire n_19;
wire n_18;
wire n_20;
wire n_35;
wire n_34;
wire n_30;
wire n_16;
wire n_24;
wire n_28;
wire n_38;
wire n_26;
wire n_36;
wire n_25;
wire n_31;
wire n_17;
wire n_29;
wire n_37;
wire n_12;
wire n_32;
wire n_15;

NAND2xp5_ASAP7_75t_L g12 ( 
.A(n_10),
.B(n_0),
.Y(n_12)
);

INVx2_ASAP7_75t_L g13 ( 
.A(n_4),
.Y(n_13)
);

BUFx3_ASAP7_75t_L g14 ( 
.A(n_0),
.Y(n_14)
);

BUFx6f_ASAP7_75t_L g15 ( 
.A(n_1),
.Y(n_15)
);

NOR2xp33_ASAP7_75t_L g16 ( 
.A(n_2),
.B(n_9),
.Y(n_16)
);

INVx11_ASAP7_75t_L g17 ( 
.A(n_8),
.Y(n_17)
);

NAND2xp5_ASAP7_75t_L g18 ( 
.A(n_5),
.B(n_1),
.Y(n_18)
);

INVx6_ASAP7_75t_L g19 ( 
.A(n_3),
.Y(n_19)
);

INVx2_ASAP7_75t_L g20 ( 
.A(n_7),
.Y(n_20)
);

INVx2_ASAP7_75t_SL g21 ( 
.A(n_3),
.Y(n_21)
);

CKINVDCx14_ASAP7_75t_R g22 ( 
.A(n_2),
.Y(n_22)
);

INVx6_ASAP7_75t_L g23 ( 
.A(n_11),
.Y(n_23)
);

INVx11_ASAP7_75t_L g24 ( 
.A(n_6),
.Y(n_24)
);

INVx4_ASAP7_75t_L g25 ( 
.A(n_14),
.Y(n_25)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_25),
.Y(n_32)
);

INVx13_ASAP7_75t_L g26 ( 
.A(n_21),
.Y(n_26)
);

OAI21xp5_ASAP7_75t_L g34 ( 
.A1(n_26),
.A2(n_27),
.B(n_28),
.Y(n_34)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_15),
.Y(n_27)
);

NOR2xp33_ASAP7_75t_SL g28 ( 
.A(n_16),
.B(n_12),
.Y(n_28)
);

INVx8_ASAP7_75t_L g29 ( 
.A(n_15),
.Y(n_29)
);

AOI21xp5_ASAP7_75t_L g33 ( 
.A1(n_29),
.A2(n_30),
.B(n_31),
.Y(n_33)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_19),
.Y(n_30)
);

AND2x6_ASAP7_75t_L g31 ( 
.A(n_18),
.B(n_22),
.Y(n_31)
);

NAND2xp5_ASAP7_75t_L g35 ( 
.A(n_34),
.B(n_16),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_SL g37 ( 
.A(n_35),
.B(n_36),
.Y(n_37)
);

OAI22xp5_ASAP7_75t_L g36 ( 
.A1(n_33),
.A2(n_31),
.B1(n_13),
.B2(n_20),
.Y(n_36)
);

AOI322xp5_ASAP7_75t_L g38 ( 
.A1(n_37),
.A2(n_23),
.A3(n_26),
.B1(n_32),
.B2(n_22),
.C1(n_21),
.C2(n_29),
.Y(n_38)
);

MAJIxp5_ASAP7_75t_L g39 ( 
.A(n_38),
.B(n_17),
.C(n_24),
.Y(n_39)
);


endmodule