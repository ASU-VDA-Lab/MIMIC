module fake_ariane_2888_n_2270 (n_295, n_356, n_170, n_190, n_160, n_64, n_180, n_119, n_124, n_386, n_307, n_332, n_294, n_197, n_176, n_34, n_172, n_347, n_183, n_373, n_299, n_12, n_133, n_66, n_205, n_341, n_71, n_109, n_245, n_96, n_319, n_49, n_20, n_283, n_50, n_187, n_367, n_345, n_374, n_318, n_103, n_244, n_226, n_220, n_261, n_36, n_370, n_189, n_72, n_286, n_57, n_387, n_117, n_139, n_85, n_130, n_349, n_391, n_346, n_214, n_348, n_2, n_32, n_379, n_138, n_162, n_264, n_137, n_122, n_198, n_232, n_52, n_385, n_73, n_327, n_77, n_372, n_377, n_15, n_23, n_87, n_279, n_207, n_363, n_354, n_41, n_140, n_151, n_28, n_146, n_230, n_270, n_194, n_154, n_338, n_142, n_285, n_186, n_202, n_145, n_193, n_59, n_336, n_315, n_311, n_239, n_35, n_272, n_54, n_8, n_339, n_167, n_90, n_38, n_47, n_153, n_18, n_269, n_75, n_158, n_69, n_259, n_95, n_143, n_152, n_120, n_169, n_106, n_173, n_242, n_309, n_320, n_115, n_331, n_267, n_335, n_350, n_291, n_344, n_381, n_62, n_210, n_200, n_166, n_253, n_218, n_79, n_3, n_271, n_247, n_91, n_240, n_369, n_128, n_224, n_44, n_82, n_31, n_222, n_256, n_326, n_227, n_48, n_188, n_323, n_330, n_11, n_129, n_126, n_282, n_328, n_368, n_277, n_248, n_301, n_293, n_228, n_325, n_276, n_93, n_108, n_303, n_168, n_81, n_1, n_206, n_352, n_238, n_365, n_136, n_334, n_192, n_300, n_14, n_163, n_88, n_141, n_390, n_104, n_314, n_16, n_273, n_305, n_312, n_233, n_56, n_60, n_388, n_333, n_392, n_376, n_221, n_321, n_86, n_361, n_89, n_149, n_383, n_237, n_175, n_74, n_19, n_40, n_181, n_53, n_260, n_362, n_310, n_236, n_281, n_24, n_7, n_209, n_262, n_17, n_225, n_235, n_297, n_290, n_46, n_84, n_371, n_199, n_107, n_217, n_178, n_42, n_308, n_201, n_70, n_343, n_10, n_287, n_302, n_380, n_6, n_94, n_284, n_4, n_249, n_37, n_58, n_65, n_123, n_212, n_355, n_278, n_255, n_257, n_148, n_135, n_171, n_384, n_61, n_102, n_182, n_316, n_196, n_125, n_43, n_13, n_27, n_254, n_219, n_55, n_231, n_366, n_234, n_280, n_215, n_252, n_161, n_298, n_68, n_78, n_63, n_99, n_216, n_5, n_223, n_25, n_83, n_389, n_288, n_179, n_195, n_213, n_110, n_304, n_67, n_306, n_313, n_92, n_203, n_378, n_150, n_98, n_375, n_113, n_114, n_33, n_324, n_337, n_111, n_21, n_274, n_296, n_265, n_208, n_156, n_292, n_174, n_275, n_100, n_132, n_147, n_204, n_51, n_76, n_342, n_26, n_246, n_0, n_159, n_358, n_105, n_30, n_131, n_263, n_360, n_229, n_394, n_250, n_165, n_144, n_317, n_101, n_243, n_134, n_329, n_185, n_340, n_289, n_9, n_112, n_45, n_268, n_266, n_164, n_157, n_184, n_177, n_364, n_258, n_118, n_121, n_353, n_22, n_241, n_29, n_357, n_191, n_382, n_80, n_211, n_97, n_322, n_251, n_116, n_351, n_39, n_393, n_359, n_155, n_127, n_2270);

input n_295;
input n_356;
input n_170;
input n_190;
input n_160;
input n_64;
input n_180;
input n_119;
input n_124;
input n_386;
input n_307;
input n_332;
input n_294;
input n_197;
input n_176;
input n_34;
input n_172;
input n_347;
input n_183;
input n_373;
input n_299;
input n_12;
input n_133;
input n_66;
input n_205;
input n_341;
input n_71;
input n_109;
input n_245;
input n_96;
input n_319;
input n_49;
input n_20;
input n_283;
input n_50;
input n_187;
input n_367;
input n_345;
input n_374;
input n_318;
input n_103;
input n_244;
input n_226;
input n_220;
input n_261;
input n_36;
input n_370;
input n_189;
input n_72;
input n_286;
input n_57;
input n_387;
input n_117;
input n_139;
input n_85;
input n_130;
input n_349;
input n_391;
input n_346;
input n_214;
input n_348;
input n_2;
input n_32;
input n_379;
input n_138;
input n_162;
input n_264;
input n_137;
input n_122;
input n_198;
input n_232;
input n_52;
input n_385;
input n_73;
input n_327;
input n_77;
input n_372;
input n_377;
input n_15;
input n_23;
input n_87;
input n_279;
input n_207;
input n_363;
input n_354;
input n_41;
input n_140;
input n_151;
input n_28;
input n_146;
input n_230;
input n_270;
input n_194;
input n_154;
input n_338;
input n_142;
input n_285;
input n_186;
input n_202;
input n_145;
input n_193;
input n_59;
input n_336;
input n_315;
input n_311;
input n_239;
input n_35;
input n_272;
input n_54;
input n_8;
input n_339;
input n_167;
input n_90;
input n_38;
input n_47;
input n_153;
input n_18;
input n_269;
input n_75;
input n_158;
input n_69;
input n_259;
input n_95;
input n_143;
input n_152;
input n_120;
input n_169;
input n_106;
input n_173;
input n_242;
input n_309;
input n_320;
input n_115;
input n_331;
input n_267;
input n_335;
input n_350;
input n_291;
input n_344;
input n_381;
input n_62;
input n_210;
input n_200;
input n_166;
input n_253;
input n_218;
input n_79;
input n_3;
input n_271;
input n_247;
input n_91;
input n_240;
input n_369;
input n_128;
input n_224;
input n_44;
input n_82;
input n_31;
input n_222;
input n_256;
input n_326;
input n_227;
input n_48;
input n_188;
input n_323;
input n_330;
input n_11;
input n_129;
input n_126;
input n_282;
input n_328;
input n_368;
input n_277;
input n_248;
input n_301;
input n_293;
input n_228;
input n_325;
input n_276;
input n_93;
input n_108;
input n_303;
input n_168;
input n_81;
input n_1;
input n_206;
input n_352;
input n_238;
input n_365;
input n_136;
input n_334;
input n_192;
input n_300;
input n_14;
input n_163;
input n_88;
input n_141;
input n_390;
input n_104;
input n_314;
input n_16;
input n_273;
input n_305;
input n_312;
input n_233;
input n_56;
input n_60;
input n_388;
input n_333;
input n_392;
input n_376;
input n_221;
input n_321;
input n_86;
input n_361;
input n_89;
input n_149;
input n_383;
input n_237;
input n_175;
input n_74;
input n_19;
input n_40;
input n_181;
input n_53;
input n_260;
input n_362;
input n_310;
input n_236;
input n_281;
input n_24;
input n_7;
input n_209;
input n_262;
input n_17;
input n_225;
input n_235;
input n_297;
input n_290;
input n_46;
input n_84;
input n_371;
input n_199;
input n_107;
input n_217;
input n_178;
input n_42;
input n_308;
input n_201;
input n_70;
input n_343;
input n_10;
input n_287;
input n_302;
input n_380;
input n_6;
input n_94;
input n_284;
input n_4;
input n_249;
input n_37;
input n_58;
input n_65;
input n_123;
input n_212;
input n_355;
input n_278;
input n_255;
input n_257;
input n_148;
input n_135;
input n_171;
input n_384;
input n_61;
input n_102;
input n_182;
input n_316;
input n_196;
input n_125;
input n_43;
input n_13;
input n_27;
input n_254;
input n_219;
input n_55;
input n_231;
input n_366;
input n_234;
input n_280;
input n_215;
input n_252;
input n_161;
input n_298;
input n_68;
input n_78;
input n_63;
input n_99;
input n_216;
input n_5;
input n_223;
input n_25;
input n_83;
input n_389;
input n_288;
input n_179;
input n_195;
input n_213;
input n_110;
input n_304;
input n_67;
input n_306;
input n_313;
input n_92;
input n_203;
input n_378;
input n_150;
input n_98;
input n_375;
input n_113;
input n_114;
input n_33;
input n_324;
input n_337;
input n_111;
input n_21;
input n_274;
input n_296;
input n_265;
input n_208;
input n_156;
input n_292;
input n_174;
input n_275;
input n_100;
input n_132;
input n_147;
input n_204;
input n_51;
input n_76;
input n_342;
input n_26;
input n_246;
input n_0;
input n_159;
input n_358;
input n_105;
input n_30;
input n_131;
input n_263;
input n_360;
input n_229;
input n_394;
input n_250;
input n_165;
input n_144;
input n_317;
input n_101;
input n_243;
input n_134;
input n_329;
input n_185;
input n_340;
input n_289;
input n_9;
input n_112;
input n_45;
input n_268;
input n_266;
input n_164;
input n_157;
input n_184;
input n_177;
input n_364;
input n_258;
input n_118;
input n_121;
input n_353;
input n_22;
input n_241;
input n_29;
input n_357;
input n_191;
input n_382;
input n_80;
input n_211;
input n_97;
input n_322;
input n_251;
input n_116;
input n_351;
input n_39;
input n_393;
input n_359;
input n_155;
input n_127;

output n_2270;

wire n_913;
wire n_1681;
wire n_2163;
wire n_1507;
wire n_1486;
wire n_1938;
wire n_589;
wire n_1174;
wire n_1469;
wire n_691;
wire n_1353;
wire n_1355;
wire n_2131;
wire n_423;
wire n_1383;
wire n_2182;
wire n_603;
wire n_2135;
wire n_1250;
wire n_2030;
wire n_1169;
wire n_789;
wire n_850;
wire n_1916;
wire n_610;
wire n_1713;
wire n_1436;
wire n_690;
wire n_416;
wire n_1109;
wire n_1430;
wire n_525;
wire n_2002;
wire n_1463;
wire n_2243;
wire n_1238;
wire n_2011;
wire n_1515;
wire n_817;
wire n_1837;
wire n_924;
wire n_781;
wire n_2013;
wire n_1566;
wire n_717;
wire n_2006;
wire n_952;
wire n_864;
wire n_1096;
wire n_1379;
wire n_1706;
wire n_2207;
wire n_524;
wire n_1214;
wire n_634;
wire n_1839;
wire n_1246;
wire n_1138;
wire n_2042;
wire n_2123;
wire n_1853;
wire n_764;
wire n_1503;
wire n_2238;
wire n_462;
wire n_1196;
wire n_1181;
wire n_1999;
wire n_410;
wire n_1187;
wire n_1131;
wire n_1225;
wire n_737;
wire n_1298;
wire n_1745;
wire n_1366;
wire n_2084;
wire n_568;
wire n_1088;
wire n_1424;
wire n_766;
wire n_1835;
wire n_1457;
wire n_1682;
wire n_1836;
wire n_520;
wire n_870;
wire n_1453;
wire n_945;
wire n_958;
wire n_2248;
wire n_813;
wire n_419;
wire n_1985;
wire n_995;
wire n_1909;
wire n_2156;
wire n_1184;
wire n_1961;
wire n_1535;
wire n_500;
wire n_754;
wire n_665;
wire n_903;
wire n_871;
wire n_1073;
wire n_402;
wire n_1979;
wire n_1277;
wire n_2107;
wire n_1746;
wire n_829;
wire n_1761;
wire n_1062;
wire n_738;
wire n_1690;
wire n_2221;
wire n_672;
wire n_740;
wire n_1283;
wire n_1974;
wire n_1736;
wire n_1018;
wire n_2200;
wire n_953;
wire n_1364;
wire n_1888;
wire n_1224;
wire n_2109;
wire n_1425;
wire n_625;
wire n_557;
wire n_1107;
wire n_1688;
wire n_989;
wire n_645;
wire n_1944;
wire n_559;
wire n_2233;
wire n_495;
wire n_1988;
wire n_795;
wire n_721;
wire n_1084;
wire n_1718;
wire n_1276;
wire n_1936;
wire n_2149;
wire n_1428;
wire n_1284;
wire n_1241;
wire n_821;
wire n_561;
wire n_770;
wire n_1514;
wire n_1528;
wire n_507;
wire n_486;
wire n_901;
wire n_569;
wire n_2078;
wire n_1145;
wire n_971;
wire n_2201;
wire n_787;
wire n_1650;
wire n_1519;
wire n_1195;
wire n_2049;
wire n_1522;
wire n_518;
wire n_1207;
wire n_786;
wire n_1404;
wire n_868;
wire n_2232;
wire n_1847;
wire n_1542;
wire n_1314;
wire n_1512;
wire n_2227;
wire n_1539;
wire n_884;
wire n_1851;
wire n_2162;
wire n_1415;
wire n_1034;
wire n_1652;
wire n_2192;
wire n_1676;
wire n_1085;
wire n_1636;
wire n_432;
wire n_823;
wire n_1900;
wire n_620;
wire n_1074;
wire n_859;
wire n_1765;
wire n_1889;
wire n_587;
wire n_1977;
wire n_693;
wire n_863;
wire n_1254;
wire n_929;
wire n_899;
wire n_1703;
wire n_611;
wire n_1295;
wire n_2060;
wire n_1850;
wire n_2004;
wire n_1013;
wire n_1495;
wire n_1637;
wire n_661;
wire n_2098;
wire n_1751;
wire n_533;
wire n_1917;
wire n_1924;
wire n_438;
wire n_1560;
wire n_1654;
wire n_1548;
wire n_1811;
wire n_2045;
wire n_440;
wire n_1396;
wire n_1230;
wire n_612;
wire n_1840;
wire n_512;
wire n_1597;
wire n_1771;
wire n_1544;
wire n_579;
wire n_844;
wire n_1012;
wire n_1267;
wire n_2061;
wire n_2094;
wire n_1354;
wire n_1790;
wire n_1213;
wire n_2043;
wire n_780;
wire n_1918;
wire n_1021;
wire n_1443;
wire n_491;
wire n_1465;
wire n_1949;
wire n_1595;
wire n_1142;
wire n_1140;
wire n_705;
wire n_570;
wire n_942;
wire n_1437;
wire n_2077;
wire n_1378;
wire n_461;
wire n_1121;
wire n_1416;
wire n_490;
wire n_1461;
wire n_1391;
wire n_1947;
wire n_1599;
wire n_1876;
wire n_1006;
wire n_1830;
wire n_575;
wire n_546;
wire n_503;
wire n_1112;
wire n_700;
wire n_1159;
wire n_772;
wire n_1216;
wire n_1245;
wire n_1669;
wire n_1675;
wire n_676;
wire n_2038;
wire n_2263;
wire n_2116;
wire n_2145;
wire n_1838;
wire n_1594;
wire n_680;
wire n_1935;
wire n_1716;
wire n_1872;
wire n_1585;
wire n_1432;
wire n_2245;
wire n_1108;
wire n_851;
wire n_444;
wire n_1590;
wire n_1351;
wire n_2216;
wire n_1274;
wire n_652;
wire n_1819;
wire n_475;
wire n_947;
wire n_2134;
wire n_1260;
wire n_930;
wire n_1179;
wire n_468;
wire n_1442;
wire n_696;
wire n_482;
wire n_798;
wire n_1833;
wire n_577;
wire n_407;
wire n_1691;
wire n_916;
wire n_1386;
wire n_912;
wire n_1884;
wire n_460;
wire n_1555;
wire n_1842;
wire n_762;
wire n_1253;
wire n_1468;
wire n_1661;
wire n_555;
wire n_804;
wire n_1656;
wire n_1382;
wire n_992;
wire n_966;
wire n_955;
wire n_1182;
wire n_794;
wire n_2166;
wire n_1692;
wire n_1562;
wire n_514;
wire n_418;
wire n_2185;
wire n_1376;
wire n_513;
wire n_1292;
wire n_1972;
wire n_2015;
wire n_1178;
wire n_1435;
wire n_1750;
wire n_1026;
wire n_1506;
wire n_1610;
wire n_2202;
wire n_2072;
wire n_436;
wire n_2087;
wire n_669;
wire n_1491;
wire n_931;
wire n_619;
wire n_437;
wire n_1083;
wire n_967;
wire n_2161;
wire n_1418;
wire n_746;
wire n_1357;
wire n_1079;
wire n_1787;
wire n_1389;
wire n_2155;
wire n_615;
wire n_1139;
wire n_517;
wire n_1312;
wire n_1717;
wire n_1812;
wire n_824;
wire n_428;
wire n_2172;
wire n_892;
wire n_1880;
wire n_959;
wire n_2257;
wire n_1399;
wire n_1101;
wire n_1567;
wire n_1343;
wire n_563;
wire n_2219;
wire n_1855;
wire n_2100;
wire n_1623;
wire n_990;
wire n_1903;
wire n_867;
wire n_2147;
wire n_1226;
wire n_2224;
wire n_944;
wire n_749;
wire n_1932;
wire n_1780;
wire n_1970;
wire n_1920;
wire n_2083;
wire n_815;
wire n_542;
wire n_2167;
wire n_1340;
wire n_470;
wire n_1240;
wire n_1087;
wire n_632;
wire n_477;
wire n_650;
wire n_425;
wire n_1433;
wire n_1911;
wire n_1825;
wire n_1908;
wire n_1155;
wire n_1071;
wire n_976;
wire n_712;
wire n_909;
wire n_1392;
wire n_767;
wire n_1832;
wire n_1841;
wire n_1680;
wire n_2066;
wire n_964;
wire n_1627;
wire n_2220;
wire n_489;
wire n_974;
wire n_506;
wire n_1731;
wire n_799;
wire n_1147;
wire n_397;
wire n_471;
wire n_1914;
wire n_965;
wire n_2253;
wire n_934;
wire n_2213;
wire n_1447;
wire n_1220;
wire n_2019;
wire n_698;
wire n_2130;
wire n_1674;
wire n_2021;
wire n_2025;
wire n_2160;
wire n_1992;
wire n_1209;
wire n_1020;
wire n_1563;
wire n_646;
wire n_2142;
wire n_1633;
wire n_404;
wire n_1913;
wire n_2069;
wire n_1058;
wire n_1042;
wire n_1234;
wire n_479;
wire n_1578;
wire n_2261;
wire n_1455;
wire n_836;
wire n_2223;
wire n_1279;
wire n_2144;
wire n_564;
wire n_1029;
wire n_1247;
wire n_760;
wire n_522;
wire n_1568;
wire n_1483;
wire n_1363;
wire n_1111;
wire n_1689;
wire n_970;
wire n_713;
wire n_1255;
wire n_1646;
wire n_598;
wire n_2262;
wire n_1237;
wire n_927;
wire n_1095;
wire n_1728;
wire n_706;
wire n_2120;
wire n_1401;
wire n_1419;
wire n_1531;
wire n_776;
wire n_424;
wire n_2041;
wire n_2113;
wire n_1933;
wire n_1651;
wire n_1387;
wire n_466;
wire n_1263;
wire n_1817;
wire n_2168;
wire n_552;
wire n_670;
wire n_1826;
wire n_441;
wire n_1951;
wire n_1032;
wire n_1217;
wire n_1496;
wire n_637;
wire n_1592;
wire n_1259;
wire n_1177;
wire n_1231;
wire n_2132;
wire n_980;
wire n_1618;
wire n_1869;
wire n_1743;
wire n_905;
wire n_720;
wire n_926;
wire n_1943;
wire n_1802;
wire n_2178;
wire n_2112;
wire n_1163;
wire n_1795;
wire n_1384;
wire n_2237;
wire n_2146;
wire n_1868;
wire n_1501;
wire n_2241;
wire n_1173;
wire n_1068;
wire n_1198;
wire n_1570;
wire n_2099;
wire n_487;
wire n_1518;
wire n_1456;
wire n_1879;
wire n_1886;
wire n_1648;
wire n_2187;
wire n_1413;
wire n_2129;
wire n_855;
wire n_808;
wire n_1365;
wire n_553;
wire n_2059;
wire n_1439;
wire n_814;
wire n_578;
wire n_2074;
wire n_1665;
wire n_1287;
wire n_405;
wire n_1611;
wire n_2122;
wire n_1414;
wire n_1134;
wire n_2067;
wire n_1484;
wire n_1901;
wire n_647;
wire n_2055;
wire n_2027;
wire n_1423;
wire n_2117;
wire n_481;
wire n_600;
wire n_1053;
wire n_1609;
wire n_1939;
wire n_2242;
wire n_1906;
wire n_529;
wire n_1899;
wire n_2195;
wire n_502;
wire n_2194;
wire n_1467;
wire n_1828;
wire n_2159;
wire n_1798;
wire n_1304;
wire n_1608;
wire n_1744;
wire n_2267;
wire n_1105;
wire n_547;
wire n_439;
wire n_604;
wire n_677;
wire n_478;
wire n_703;
wire n_1349;
wire n_1709;
wire n_1061;
wire n_2102;
wire n_681;
wire n_874;
wire n_2023;
wire n_1278;
wire n_707;
wire n_983;
wire n_699;
wire n_727;
wire n_590;
wire n_1726;
wire n_2075;
wire n_1945;
wire n_1015;
wire n_545;
wire n_1377;
wire n_1162;
wire n_536;
wire n_1614;
wire n_2031;
wire n_2118;
wire n_1740;
wire n_1602;
wire n_688;
wire n_636;
wire n_427;
wire n_1098;
wire n_1490;
wire n_442;
wire n_777;
wire n_1553;
wire n_1080;
wire n_920;
wire n_1760;
wire n_1086;
wire n_1092;
wire n_2225;
wire n_986;
wire n_1104;
wire n_1963;
wire n_729;
wire n_887;
wire n_2057;
wire n_2218;
wire n_1122;
wire n_1205;
wire n_1408;
wire n_1693;
wire n_2125;
wire n_1132;
wire n_1156;
wire n_501;
wire n_2184;
wire n_1823;
wire n_1120;
wire n_1202;
wire n_627;
wire n_2254;
wire n_1188;
wire n_1498;
wire n_1371;
wire n_2033;
wire n_1402;
wire n_957;
wire n_1242;
wire n_1607;
wire n_1489;
wire n_1218;
wire n_2217;
wire n_2226;
wire n_1586;
wire n_861;
wire n_1543;
wire n_1431;
wire n_877;
wire n_1119;
wire n_1863;
wire n_1763;
wire n_1666;
wire n_1500;
wire n_616;
wire n_2214;
wire n_1055;
wire n_1395;
wire n_1346;
wire n_2256;
wire n_1189;
wire n_1089;
wire n_1859;
wire n_1502;
wire n_1523;
wire n_2190;
wire n_1478;
wire n_1883;
wire n_1969;
wire n_735;
wire n_1005;
wire n_527;
wire n_1294;
wire n_1667;
wire n_845;
wire n_888;
wire n_1649;
wire n_1677;
wire n_1927;
wire n_1297;
wire n_551;
wire n_417;
wire n_1708;
wire n_1222;
wire n_1844;
wire n_582;
wire n_1957;
wire n_1953;
wire n_755;
wire n_1097;
wire n_1219;
wire n_1711;
wire n_1919;
wire n_710;
wire n_534;
wire n_1791;
wire n_2124;
wire n_1894;
wire n_1460;
wire n_1239;
wire n_2266;
wire n_560;
wire n_890;
wire n_842;
wire n_1898;
wire n_451;
wire n_745;
wire n_1741;
wire n_1572;
wire n_1907;
wire n_1793;
wire n_742;
wire n_1081;
wire n_1373;
wire n_1975;
wire n_1388;
wire n_1266;
wire n_1540;
wire n_1719;
wire n_2119;
wire n_769;
wire n_1797;
wire n_1753;
wire n_1990;
wire n_1372;
wire n_476;
wire n_832;
wire n_535;
wire n_744;
wire n_1895;
wire n_982;
wire n_1800;
wire n_915;
wire n_1075;
wire n_2008;
wire n_454;
wire n_1331;
wire n_1890;
wire n_1529;
wire n_1227;
wire n_2127;
wire n_655;
wire n_1734;
wire n_1860;
wire n_403;
wire n_1007;
wire n_1580;
wire n_1319;
wire n_657;
wire n_837;
wire n_812;
wire n_2211;
wire n_606;
wire n_951;
wire n_862;
wire n_1700;
wire n_659;
wire n_1332;
wire n_509;
wire n_1854;
wire n_666;
wire n_1747;
wire n_2071;
wire n_430;
wire n_1206;
wire n_1729;
wire n_722;
wire n_1508;
wire n_2082;
wire n_1532;
wire n_1171;
wire n_1030;
wire n_785;
wire n_1309;
wire n_999;
wire n_1766;
wire n_1338;
wire n_1342;
wire n_456;
wire n_1867;
wire n_852;
wire n_1394;
wire n_704;
wire n_1060;
wire n_1044;
wire n_1714;
wire n_521;
wire n_2140;
wire n_873;
wire n_1301;
wire n_1748;
wire n_2157;
wire n_1966;
wire n_1243;
wire n_2171;
wire n_1400;
wire n_2035;
wire n_1466;
wire n_1527;
wire n_1513;
wire n_1783;
wire n_608;
wire n_1538;
wire n_2128;
wire n_1037;
wire n_1329;
wire n_1993;
wire n_1545;
wire n_1257;
wire n_1480;
wire n_1954;
wire n_1668;
wire n_1878;
wire n_1605;
wire n_1078;
wire n_1897;
wire n_2137;
wire n_1161;
wire n_811;
wire n_624;
wire n_791;
wire n_876;
wire n_1191;
wire n_618;
wire n_736;
wire n_1025;
wire n_1215;
wire n_1449;
wire n_2265;
wire n_687;
wire n_797;
wire n_2026;
wire n_1786;
wire n_480;
wire n_1327;
wire n_1475;
wire n_642;
wire n_1804;
wire n_2106;
wire n_408;
wire n_1406;
wire n_595;
wire n_1405;
wire n_602;
wire n_1757;
wire n_592;
wire n_1499;
wire n_854;
wire n_1318;
wire n_2091;
wire n_1632;
wire n_1769;
wire n_474;
wire n_1929;
wire n_1950;
wire n_2264;
wire n_805;
wire n_2032;
wire n_2090;
wire n_1658;
wire n_2249;
wire n_1072;
wire n_695;
wire n_1526;
wire n_1305;
wire n_730;
wire n_1596;
wire n_1281;
wire n_516;
wire n_1997;
wire n_1137;
wire n_1873;
wire n_1258;
wire n_640;
wire n_1733;
wire n_463;
wire n_1476;
wire n_1524;
wire n_1856;
wire n_2016;
wire n_943;
wire n_1118;
wire n_678;
wire n_651;
wire n_1874;
wire n_1293;
wire n_961;
wire n_469;
wire n_1046;
wire n_1807;
wire n_1123;
wire n_726;
wire n_1657;
wire n_878;
wire n_1784;
wire n_771;
wire n_1321;
wire n_752;
wire n_1488;
wire n_985;
wire n_421;
wire n_1330;
wire n_906;
wire n_1180;
wire n_1697;
wire n_806;
wire n_1984;
wire n_1350;
wire n_1556;
wire n_649;
wire n_1561;
wire n_1352;
wire n_1824;
wire n_643;
wire n_1492;
wire n_1441;
wire n_1822;
wire n_682;
wire n_1616;
wire n_819;
wire n_1971;
wire n_1429;
wire n_1324;
wire n_586;
wire n_2064;
wire n_1778;
wire n_1776;
wire n_686;
wire n_605;
wire n_1154;
wire n_584;
wire n_1557;
wire n_1759;
wire n_1829;
wire n_1130;
wire n_1450;
wire n_756;
wire n_2022;
wire n_1016;
wire n_1149;
wire n_1505;
wire n_979;
wire n_1642;
wire n_1815;
wire n_897;
wire n_949;
wire n_1493;
wire n_515;
wire n_807;
wire n_891;
wire n_885;
wire n_1659;
wire n_1864;
wire n_1887;
wire n_1208;
wire n_1987;
wire n_396;
wire n_802;
wire n_1151;
wire n_554;
wire n_960;
wire n_1256;
wire n_714;
wire n_2170;
wire n_790;
wire n_2244;
wire n_2143;
wire n_725;
wire n_1577;
wire n_1448;
wire n_2198;
wire n_1009;
wire n_1133;
wire n_883;
wire n_473;
wire n_1852;
wire n_801;
wire n_1286;
wire n_818;
wire n_1685;
wire n_779;
wire n_594;
wire n_2222;
wire n_1995;
wire n_1877;
wire n_1397;
wire n_1052;
wire n_1333;
wire n_1306;
wire n_1849;
wire n_2076;
wire n_2133;
wire n_2203;
wire n_833;
wire n_1426;
wire n_2250;
wire n_2247;
wire n_2230;
wire n_879;
wire n_1117;
wire n_422;
wire n_1269;
wire n_1303;
wire n_1547;
wire n_1438;
wire n_1541;
wire n_597;
wire n_2001;
wire n_1047;
wire n_1472;
wire n_1593;
wire n_1050;
wire n_566;
wire n_2158;
wire n_1288;
wire n_1201;
wire n_858;
wire n_1185;
wire n_2173;
wire n_1035;
wire n_1143;
wire n_2070;
wire n_2136;
wire n_426;
wire n_433;
wire n_398;
wire n_1090;
wire n_1367;
wire n_2044;
wire n_928;
wire n_1153;
wire n_465;
wire n_825;
wire n_1103;
wire n_732;
wire n_1565;
wire n_1192;
wire n_894;
wire n_1380;
wire n_1624;
wire n_1801;
wire n_420;
wire n_1291;
wire n_562;
wire n_2020;
wire n_748;
wire n_510;
wire n_1045;
wire n_1160;
wire n_1882;
wire n_1976;
wire n_1023;
wire n_1881;
wire n_988;
wire n_914;
wire n_689;
wire n_400;
wire n_1116;
wire n_1958;
wire n_467;
wire n_1511;
wire n_2177;
wire n_1422;
wire n_1965;
wire n_644;
wire n_1197;
wire n_497;
wire n_1165;
wire n_1641;
wire n_538;
wire n_1517;
wire n_2036;
wire n_576;
wire n_843;
wire n_511;
wire n_455;
wire n_429;
wire n_588;
wire n_638;
wire n_2003;
wire n_2210;
wire n_1307;
wire n_1128;
wire n_2053;
wire n_1671;
wire n_1417;
wire n_1048;
wire n_775;
wire n_667;
wire n_1049;
wire n_869;
wire n_846;
wire n_1398;
wire n_1921;
wire n_1356;
wire n_1341;
wire n_2234;
wire n_1504;
wire n_1955;
wire n_2110;
wire n_1773;
wire n_1440;
wire n_1603;
wire n_1370;
wire n_728;
wire n_413;
wire n_715;
wire n_889;
wire n_1066;
wire n_1549;
wire n_935;
wire n_685;
wire n_911;
wire n_623;
wire n_1712;
wire n_1403;
wire n_1065;
wire n_453;
wire n_1534;
wire n_1948;
wire n_810;
wire n_1290;
wire n_1959;
wire n_617;
wire n_543;
wire n_1362;
wire n_1559;
wire n_2121;
wire n_601;
wire n_683;
wire n_565;
wire n_628;
wire n_1300;
wire n_1960;
wire n_2068;
wire n_743;
wire n_1194;
wire n_1647;
wire n_1546;
wire n_1420;
wire n_907;
wire n_1454;
wire n_660;
wire n_464;
wire n_962;
wire n_941;
wire n_1210;
wire n_847;
wire n_747;
wire n_1622;
wire n_1135;
wire n_918;
wire n_1968;
wire n_1885;
wire n_639;
wire n_452;
wire n_673;
wire n_2196;
wire n_1038;
wire n_1978;
wire n_414;
wire n_571;
wire n_1521;
wire n_1694;
wire n_1940;
wire n_593;
wire n_1695;
wire n_1164;
wire n_609;
wire n_1193;
wire n_1345;
wire n_613;
wire n_1022;
wire n_1336;
wire n_1033;
wire n_1774;
wire n_409;
wire n_519;
wire n_1166;
wire n_1056;
wire n_2007;
wire n_526;
wire n_1994;
wire n_1767;
wire n_1040;
wire n_674;
wire n_1158;
wire n_1973;
wire n_1444;
wire n_1803;
wire n_820;
wire n_1749;
wire n_872;
wire n_1653;
wire n_1157;
wire n_1584;
wire n_848;
wire n_1664;
wire n_629;
wire n_1739;
wire n_1814;
wire n_532;
wire n_2154;
wire n_2236;
wire n_1789;
wire n_763;
wire n_1986;
wire n_2174;
wire n_540;
wire n_692;
wire n_2054;
wire n_1857;
wire n_984;
wire n_1687;
wire n_2073;
wire n_2150;
wire n_1552;
wire n_750;
wire n_834;
wire n_1612;
wire n_800;
wire n_2046;
wire n_1816;
wire n_1910;
wire n_1756;
wire n_1606;
wire n_2189;
wire n_395;
wire n_621;
wire n_1587;
wire n_2093;
wire n_2018;
wire n_1772;
wire n_1014;
wire n_724;
wire n_2204;
wire n_1427;
wire n_1481;
wire n_2040;
wire n_493;
wire n_1311;
wire n_2199;
wire n_1956;
wire n_1589;
wire n_2151;
wire n_1100;
wire n_585;
wire n_875;
wire n_1617;
wire n_827;
wire n_2231;
wire n_697;
wire n_622;
wire n_1626;
wire n_1962;
wire n_1335;
wire n_1715;
wire n_880;
wire n_793;
wire n_2114;
wire n_1175;
wire n_751;
wire n_1027;
wire n_1070;
wire n_1621;
wire n_739;
wire n_1485;
wire n_1028;
wire n_1221;
wire n_530;
wire n_1785;
wire n_792;
wire n_1262;
wire n_1942;
wire n_2180;
wire n_580;
wire n_1579;
wire n_494;
wire n_2181;
wire n_434;
wire n_2014;
wire n_975;
wire n_923;
wire n_1645;
wire n_1124;
wire n_1381;
wire n_1494;
wire n_932;
wire n_1893;
wire n_1183;
wire n_1326;
wire n_1805;
wire n_981;
wire n_2141;
wire n_1758;
wire n_1110;
wire n_1407;
wire n_1204;
wire n_1554;
wire n_994;
wire n_1360;
wire n_973;
wire n_972;
wire n_2251;
wire n_856;
wire n_1248;
wire n_1176;
wire n_1564;
wire n_2010;
wire n_1054;
wire n_508;
wire n_1679;
wire n_2126;
wire n_1952;
wire n_1858;
wire n_1678;
wire n_1482;
wire n_1361;
wire n_1601;
wire n_1057;
wire n_1834;
wire n_978;
wire n_1011;
wire n_1520;
wire n_1509;
wire n_828;
wire n_1411;
wire n_1359;
wire n_558;
wire n_1721;
wire n_653;
wire n_1445;
wire n_1317;
wire n_2050;
wire n_2197;
wire n_783;
wire n_556;
wire n_1127;
wire n_1536;
wire n_1471;
wire n_1008;
wire n_581;
wire n_1024;
wire n_830;
wire n_1980;
wire n_987;
wire n_936;
wire n_1620;
wire n_1385;
wire n_1525;
wire n_1998;
wire n_2165;
wire n_541;
wire n_499;
wire n_1775;
wire n_788;
wire n_908;
wire n_1036;
wire n_2169;
wire n_1270;
wire n_1167;
wire n_1272;
wire n_549;
wire n_591;
wire n_969;
wire n_2028;
wire n_919;
wire n_1663;
wire n_2092;
wire n_2175;
wire n_1625;
wire n_2086;
wire n_1926;
wire n_1458;
wire n_679;
wire n_1630;
wire n_663;
wire n_1720;
wire n_443;
wire n_2176;
wire n_1412;
wire n_1738;
wire n_1550;
wire n_528;
wire n_1358;
wire n_1200;
wire n_406;
wire n_826;
wire n_1922;
wire n_1735;
wire n_1788;
wire n_940;
wire n_1537;
wire n_2138;
wire n_2065;
wire n_1077;
wire n_607;
wire n_956;
wire n_445;
wire n_1930;
wire n_765;
wire n_1809;
wire n_1843;
wire n_1904;
wire n_2000;
wire n_1268;
wire n_917;
wire n_1271;
wire n_2096;
wire n_2186;
wire n_1530;
wire n_2215;
wire n_631;
wire n_399;
wire n_1170;
wire n_2258;
wire n_1261;
wire n_702;
wire n_898;
wire n_857;
wire n_968;
wire n_1067;
wire n_1235;
wire n_1323;
wire n_1462;
wire n_1937;
wire n_2012;
wire n_1064;
wire n_633;
wire n_900;
wire n_1446;
wire n_1282;
wire n_1701;
wire n_1093;
wire n_1551;
wire n_2039;
wire n_1755;
wire n_1285;
wire n_733;
wire n_761;
wire n_2212;
wire n_731;
wire n_1813;
wire n_2268;
wire n_1452;
wire n_1573;
wire n_668;
wire n_758;
wire n_2252;
wire n_2111;
wire n_1996;
wire n_1106;
wire n_2009;
wire n_648;
wire n_784;
wire n_816;
wire n_1322;
wire n_1473;
wire n_835;
wire n_446;
wire n_1076;
wire n_2024;
wire n_1348;
wire n_753;
wire n_1770;
wire n_1003;
wire n_701;
wire n_1125;
wire n_2103;
wire n_1710;
wire n_1865;
wire n_1344;
wire n_1390;
wire n_401;
wire n_485;
wire n_1792;
wire n_504;
wire n_2062;
wire n_483;
wire n_435;
wire n_1141;
wire n_1629;
wire n_1640;
wire n_822;
wire n_1094;
wire n_840;
wire n_1459;
wire n_2153;
wire n_1510;
wire n_2139;
wire n_1099;
wire n_839;
wire n_1754;
wire n_759;
wire n_567;
wire n_1727;
wire n_2235;
wire n_1991;
wire n_1575;
wire n_1848;
wire n_1892;
wire n_1172;
wire n_614;
wire n_1212;
wire n_831;
wire n_778;
wire n_1619;
wire n_2260;
wire n_550;
wire n_1660;
wire n_1315;
wire n_1902;
wire n_997;
wire n_635;
wire n_2206;
wire n_694;
wire n_1643;
wire n_1320;
wire n_1113;
wire n_1152;
wire n_2034;
wire n_1845;
wire n_1934;
wire n_2101;
wire n_921;
wire n_1615;
wire n_1236;
wire n_2104;
wire n_1265;
wire n_1576;
wire n_2105;
wire n_1470;
wire n_1533;
wire n_1806;
wire n_671;
wire n_1684;
wire n_1148;
wire n_1588;
wire n_1409;
wire n_1673;
wire n_1334;
wire n_654;
wire n_2088;
wire n_1275;
wire n_488;
wire n_904;
wire n_505;
wire n_2005;
wire n_2048;
wire n_1696;
wire n_498;
wire n_1875;
wire n_1059;
wire n_684;
wire n_2108;
wire n_1039;
wire n_2246;
wire n_539;
wire n_1150;
wire n_977;
wire n_449;
wire n_1628;
wire n_1289;
wire n_1831;
wire n_2191;
wire n_1497;
wire n_1866;
wire n_2056;
wire n_459;
wire n_1136;
wire n_1782;
wire n_458;
wire n_1600;
wire n_1190;
wire n_1144;
wire n_838;
wire n_1558;
wire n_1941;
wire n_1316;
wire n_950;
wire n_1017;
wire n_711;
wire n_734;
wire n_1915;
wire n_723;
wire n_1393;
wire n_2240;
wire n_658;
wire n_630;
wire n_1369;
wire n_1781;
wire n_709;
wire n_809;
wire n_2085;
wire n_1686;
wire n_1964;
wire n_881;
wire n_1019;
wire n_1477;
wire n_1777;
wire n_2188;
wire n_1982;
wire n_2097;
wire n_662;
wire n_641;
wire n_910;
wire n_741;
wire n_1410;
wire n_939;
wire n_1114;
wire n_1325;
wire n_1742;
wire n_708;
wire n_1223;
wire n_1768;
wire n_2193;
wire n_572;
wire n_1199;
wire n_865;
wire n_1273;
wire n_1983;
wire n_1041;
wire n_2115;
wire n_993;
wire n_1862;
wire n_948;
wire n_2017;
wire n_922;
wire n_1004;
wire n_1810;
wire n_448;
wire n_1347;
wire n_860;
wire n_1043;
wire n_450;
wire n_1923;
wire n_1764;
wire n_896;
wire n_1737;
wire n_1479;
wire n_1613;
wire n_902;
wire n_1031;
wire n_1723;
wire n_1638;
wire n_853;
wire n_716;
wire n_1571;
wire n_1698;
wire n_1337;
wire n_774;
wire n_1946;
wire n_2148;
wire n_933;
wire n_1779;
wire n_596;
wire n_954;
wire n_2051;
wire n_1168;
wire n_1821;
wire n_1310;
wire n_656;
wire n_492;
wire n_574;
wire n_1591;
wire n_664;
wire n_1229;
wire n_1683;
wire n_1896;
wire n_2164;
wire n_1732;
wire n_415;
wire n_1967;
wire n_2179;
wire n_1280;
wire n_544;
wire n_1516;
wire n_1186;
wire n_1705;
wire n_599;
wire n_768;
wire n_1091;
wire n_2052;
wire n_1063;
wire n_537;
wire n_991;
wire n_2205;
wire n_2183;
wire n_1724;
wire n_1670;
wire n_1707;
wire n_1799;
wire n_2080;
wire n_2058;
wire n_1126;
wire n_2029;
wire n_1846;
wire n_1912;
wire n_938;
wire n_1891;
wire n_1328;
wire n_895;
wire n_1639;
wire n_583;
wire n_2209;
wire n_1302;
wire n_1000;
wire n_626;
wire n_1581;
wire n_1928;
wire n_946;
wire n_757;
wire n_2047;
wire n_1655;
wire n_1818;
wire n_1146;
wire n_1634;
wire n_1203;
wire n_998;
wire n_1699;
wire n_1598;
wire n_2269;
wire n_472;
wire n_937;
wire n_1474;
wire n_2081;
wire n_1583;
wire n_1604;
wire n_1631;
wire n_1702;
wire n_1794;
wire n_1375;
wire n_1232;
wire n_996;
wire n_1211;
wire n_1368;
wire n_963;
wire n_1264;
wire n_1082;
wire n_1725;
wire n_496;
wire n_1827;
wire n_866;
wire n_925;
wire n_1752;
wire n_1313;
wire n_1001;
wire n_1722;
wire n_1115;
wire n_2229;
wire n_1339;
wire n_1002;
wire n_1644;
wire n_1051;
wire n_719;
wire n_1102;
wire n_2255;
wire n_1252;
wire n_1129;
wire n_2239;
wire n_1464;
wire n_1296;
wire n_773;
wire n_1010;
wire n_882;
wire n_1249;
wire n_803;
wire n_1871;
wire n_718;
wire n_1434;
wire n_1905;
wire n_1569;
wire n_548;
wire n_523;
wire n_1662;
wire n_457;
wire n_1299;
wire n_1870;
wire n_2063;
wire n_1925;
wire n_782;
wire n_431;
wire n_1861;
wire n_2079;
wire n_1228;
wire n_2152;
wire n_1931;
wire n_1244;
wire n_1796;
wire n_411;
wire n_484;
wire n_2259;
wire n_849;
wire n_2095;
wire n_1820;
wire n_412;
wire n_1251;
wire n_1989;
wire n_447;
wire n_1421;
wire n_2208;
wire n_1762;
wire n_1233;
wire n_1808;
wire n_1574;
wire n_1672;
wire n_2228;
wire n_1635;
wire n_1704;
wire n_893;
wire n_1582;
wire n_841;
wire n_886;
wire n_1981;
wire n_1069;
wire n_2037;
wire n_1308;
wire n_573;
wire n_796;
wire n_531;
wire n_1730;
wire n_1374;
wire n_1451;
wire n_2089;
wire n_1487;
wire n_675;

INVx1_ASAP7_75t_L g395 ( 
.A(n_99),
.Y(n_395)
);

CKINVDCx5p33_ASAP7_75t_R g396 ( 
.A(n_190),
.Y(n_396)
);

CKINVDCx5p33_ASAP7_75t_R g397 ( 
.A(n_374),
.Y(n_397)
);

INVx2_ASAP7_75t_L g398 ( 
.A(n_298),
.Y(n_398)
);

CKINVDCx5p33_ASAP7_75t_R g399 ( 
.A(n_321),
.Y(n_399)
);

CKINVDCx5p33_ASAP7_75t_R g400 ( 
.A(n_175),
.Y(n_400)
);

CKINVDCx5p33_ASAP7_75t_R g401 ( 
.A(n_253),
.Y(n_401)
);

BUFx3_ASAP7_75t_L g402 ( 
.A(n_362),
.Y(n_402)
);

CKINVDCx5p33_ASAP7_75t_R g403 ( 
.A(n_375),
.Y(n_403)
);

CKINVDCx5p33_ASAP7_75t_R g404 ( 
.A(n_360),
.Y(n_404)
);

CKINVDCx5p33_ASAP7_75t_R g405 ( 
.A(n_25),
.Y(n_405)
);

INVx1_ASAP7_75t_L g406 ( 
.A(n_226),
.Y(n_406)
);

INVx1_ASAP7_75t_L g407 ( 
.A(n_389),
.Y(n_407)
);

CKINVDCx5p33_ASAP7_75t_R g408 ( 
.A(n_306),
.Y(n_408)
);

CKINVDCx5p33_ASAP7_75t_R g409 ( 
.A(n_90),
.Y(n_409)
);

INVx1_ASAP7_75t_L g410 ( 
.A(n_130),
.Y(n_410)
);

INVx1_ASAP7_75t_L g411 ( 
.A(n_127),
.Y(n_411)
);

CKINVDCx5p33_ASAP7_75t_R g412 ( 
.A(n_166),
.Y(n_412)
);

INVx1_ASAP7_75t_L g413 ( 
.A(n_243),
.Y(n_413)
);

INVx1_ASAP7_75t_L g414 ( 
.A(n_3),
.Y(n_414)
);

CKINVDCx5p33_ASAP7_75t_R g415 ( 
.A(n_133),
.Y(n_415)
);

CKINVDCx5p33_ASAP7_75t_R g416 ( 
.A(n_393),
.Y(n_416)
);

INVx1_ASAP7_75t_L g417 ( 
.A(n_31),
.Y(n_417)
);

CKINVDCx16_ASAP7_75t_R g418 ( 
.A(n_223),
.Y(n_418)
);

CKINVDCx5p33_ASAP7_75t_R g419 ( 
.A(n_136),
.Y(n_419)
);

CKINVDCx5p33_ASAP7_75t_R g420 ( 
.A(n_195),
.Y(n_420)
);

CKINVDCx5p33_ASAP7_75t_R g421 ( 
.A(n_247),
.Y(n_421)
);

CKINVDCx20_ASAP7_75t_R g422 ( 
.A(n_96),
.Y(n_422)
);

CKINVDCx5p33_ASAP7_75t_R g423 ( 
.A(n_23),
.Y(n_423)
);

INVx1_ASAP7_75t_L g424 ( 
.A(n_134),
.Y(n_424)
);

CKINVDCx5p33_ASAP7_75t_R g425 ( 
.A(n_338),
.Y(n_425)
);

INVx2_ASAP7_75t_L g426 ( 
.A(n_54),
.Y(n_426)
);

CKINVDCx20_ASAP7_75t_R g427 ( 
.A(n_354),
.Y(n_427)
);

CKINVDCx5p33_ASAP7_75t_R g428 ( 
.A(n_267),
.Y(n_428)
);

CKINVDCx20_ASAP7_75t_R g429 ( 
.A(n_380),
.Y(n_429)
);

INVx1_ASAP7_75t_L g430 ( 
.A(n_99),
.Y(n_430)
);

CKINVDCx5p33_ASAP7_75t_R g431 ( 
.A(n_266),
.Y(n_431)
);

INVx1_ASAP7_75t_L g432 ( 
.A(n_4),
.Y(n_432)
);

CKINVDCx5p33_ASAP7_75t_R g433 ( 
.A(n_16),
.Y(n_433)
);

INVx1_ASAP7_75t_L g434 ( 
.A(n_104),
.Y(n_434)
);

INVx1_ASAP7_75t_L g435 ( 
.A(n_43),
.Y(n_435)
);

CKINVDCx5p33_ASAP7_75t_R g436 ( 
.A(n_216),
.Y(n_436)
);

CKINVDCx20_ASAP7_75t_R g437 ( 
.A(n_361),
.Y(n_437)
);

CKINVDCx5p33_ASAP7_75t_R g438 ( 
.A(n_157),
.Y(n_438)
);

BUFx5_ASAP7_75t_L g439 ( 
.A(n_5),
.Y(n_439)
);

BUFx3_ASAP7_75t_L g440 ( 
.A(n_1),
.Y(n_440)
);

CKINVDCx5p33_ASAP7_75t_R g441 ( 
.A(n_94),
.Y(n_441)
);

CKINVDCx5p33_ASAP7_75t_R g442 ( 
.A(n_275),
.Y(n_442)
);

BUFx10_ASAP7_75t_L g443 ( 
.A(n_67),
.Y(n_443)
);

CKINVDCx5p33_ASAP7_75t_R g444 ( 
.A(n_232),
.Y(n_444)
);

CKINVDCx5p33_ASAP7_75t_R g445 ( 
.A(n_348),
.Y(n_445)
);

INVx1_ASAP7_75t_L g446 ( 
.A(n_141),
.Y(n_446)
);

INVx1_ASAP7_75t_L g447 ( 
.A(n_251),
.Y(n_447)
);

INVx1_ASAP7_75t_L g448 ( 
.A(n_259),
.Y(n_448)
);

CKINVDCx5p33_ASAP7_75t_R g449 ( 
.A(n_392),
.Y(n_449)
);

INVxp67_ASAP7_75t_L g450 ( 
.A(n_215),
.Y(n_450)
);

INVx1_ASAP7_75t_L g451 ( 
.A(n_278),
.Y(n_451)
);

INVx2_ASAP7_75t_L g452 ( 
.A(n_387),
.Y(n_452)
);

CKINVDCx5p33_ASAP7_75t_R g453 ( 
.A(n_364),
.Y(n_453)
);

INVx1_ASAP7_75t_L g454 ( 
.A(n_274),
.Y(n_454)
);

CKINVDCx5p33_ASAP7_75t_R g455 ( 
.A(n_337),
.Y(n_455)
);

INVx1_ASAP7_75t_L g456 ( 
.A(n_207),
.Y(n_456)
);

CKINVDCx5p33_ASAP7_75t_R g457 ( 
.A(n_17),
.Y(n_457)
);

CKINVDCx5p33_ASAP7_75t_R g458 ( 
.A(n_2),
.Y(n_458)
);

INVx2_ASAP7_75t_L g459 ( 
.A(n_208),
.Y(n_459)
);

CKINVDCx5p33_ASAP7_75t_R g460 ( 
.A(n_119),
.Y(n_460)
);

CKINVDCx5p33_ASAP7_75t_R g461 ( 
.A(n_386),
.Y(n_461)
);

INVx2_ASAP7_75t_L g462 ( 
.A(n_183),
.Y(n_462)
);

INVx1_ASAP7_75t_L g463 ( 
.A(n_107),
.Y(n_463)
);

INVx1_ASAP7_75t_L g464 ( 
.A(n_98),
.Y(n_464)
);

CKINVDCx16_ASAP7_75t_R g465 ( 
.A(n_326),
.Y(n_465)
);

INVx1_ASAP7_75t_SL g466 ( 
.A(n_367),
.Y(n_466)
);

CKINVDCx5p33_ASAP7_75t_R g467 ( 
.A(n_296),
.Y(n_467)
);

CKINVDCx5p33_ASAP7_75t_R g468 ( 
.A(n_24),
.Y(n_468)
);

CKINVDCx5p33_ASAP7_75t_R g469 ( 
.A(n_104),
.Y(n_469)
);

CKINVDCx5p33_ASAP7_75t_R g470 ( 
.A(n_369),
.Y(n_470)
);

INVx1_ASAP7_75t_L g471 ( 
.A(n_276),
.Y(n_471)
);

INVx1_ASAP7_75t_L g472 ( 
.A(n_382),
.Y(n_472)
);

CKINVDCx5p33_ASAP7_75t_R g473 ( 
.A(n_39),
.Y(n_473)
);

CKINVDCx5p33_ASAP7_75t_R g474 ( 
.A(n_333),
.Y(n_474)
);

INVx1_ASAP7_75t_L g475 ( 
.A(n_27),
.Y(n_475)
);

CKINVDCx5p33_ASAP7_75t_R g476 ( 
.A(n_315),
.Y(n_476)
);

CKINVDCx5p33_ASAP7_75t_R g477 ( 
.A(n_301),
.Y(n_477)
);

CKINVDCx5p33_ASAP7_75t_R g478 ( 
.A(n_344),
.Y(n_478)
);

INVx1_ASAP7_75t_L g479 ( 
.A(n_73),
.Y(n_479)
);

CKINVDCx5p33_ASAP7_75t_R g480 ( 
.A(n_288),
.Y(n_480)
);

INVx1_ASAP7_75t_L g481 ( 
.A(n_0),
.Y(n_481)
);

INVx1_ASAP7_75t_L g482 ( 
.A(n_295),
.Y(n_482)
);

CKINVDCx20_ASAP7_75t_R g483 ( 
.A(n_62),
.Y(n_483)
);

CKINVDCx5p33_ASAP7_75t_R g484 ( 
.A(n_149),
.Y(n_484)
);

CKINVDCx5p33_ASAP7_75t_R g485 ( 
.A(n_192),
.Y(n_485)
);

INVx1_ASAP7_75t_L g486 ( 
.A(n_336),
.Y(n_486)
);

CKINVDCx5p33_ASAP7_75t_R g487 ( 
.A(n_311),
.Y(n_487)
);

BUFx2_ASAP7_75t_L g488 ( 
.A(n_52),
.Y(n_488)
);

INVx1_ASAP7_75t_L g489 ( 
.A(n_307),
.Y(n_489)
);

CKINVDCx5p33_ASAP7_75t_R g490 ( 
.A(n_231),
.Y(n_490)
);

CKINVDCx5p33_ASAP7_75t_R g491 ( 
.A(n_261),
.Y(n_491)
);

INVx1_ASAP7_75t_L g492 ( 
.A(n_319),
.Y(n_492)
);

CKINVDCx5p33_ASAP7_75t_R g493 ( 
.A(n_75),
.Y(n_493)
);

CKINVDCx5p33_ASAP7_75t_R g494 ( 
.A(n_302),
.Y(n_494)
);

INVx1_ASAP7_75t_L g495 ( 
.A(n_217),
.Y(n_495)
);

BUFx6f_ASAP7_75t_L g496 ( 
.A(n_293),
.Y(n_496)
);

CKINVDCx5p33_ASAP7_75t_R g497 ( 
.A(n_233),
.Y(n_497)
);

CKINVDCx5p33_ASAP7_75t_R g498 ( 
.A(n_76),
.Y(n_498)
);

CKINVDCx5p33_ASAP7_75t_R g499 ( 
.A(n_38),
.Y(n_499)
);

BUFx3_ASAP7_75t_L g500 ( 
.A(n_18),
.Y(n_500)
);

BUFx3_ASAP7_75t_L g501 ( 
.A(n_67),
.Y(n_501)
);

INVx1_ASAP7_75t_L g502 ( 
.A(n_280),
.Y(n_502)
);

CKINVDCx5p33_ASAP7_75t_R g503 ( 
.A(n_55),
.Y(n_503)
);

CKINVDCx5p33_ASAP7_75t_R g504 ( 
.A(n_327),
.Y(n_504)
);

INVx1_ASAP7_75t_L g505 ( 
.A(n_352),
.Y(n_505)
);

HB1xp67_ASAP7_75t_L g506 ( 
.A(n_167),
.Y(n_506)
);

CKINVDCx5p33_ASAP7_75t_R g507 ( 
.A(n_40),
.Y(n_507)
);

INVx1_ASAP7_75t_L g508 ( 
.A(n_10),
.Y(n_508)
);

CKINVDCx5p33_ASAP7_75t_R g509 ( 
.A(n_26),
.Y(n_509)
);

CKINVDCx5p33_ASAP7_75t_R g510 ( 
.A(n_299),
.Y(n_510)
);

INVx2_ASAP7_75t_L g511 ( 
.A(n_41),
.Y(n_511)
);

BUFx10_ASAP7_75t_L g512 ( 
.A(n_347),
.Y(n_512)
);

CKINVDCx12_ASAP7_75t_R g513 ( 
.A(n_196),
.Y(n_513)
);

INVx1_ASAP7_75t_L g514 ( 
.A(n_200),
.Y(n_514)
);

INVx1_ASAP7_75t_L g515 ( 
.A(n_66),
.Y(n_515)
);

CKINVDCx5p33_ASAP7_75t_R g516 ( 
.A(n_51),
.Y(n_516)
);

CKINVDCx5p33_ASAP7_75t_R g517 ( 
.A(n_123),
.Y(n_517)
);

CKINVDCx5p33_ASAP7_75t_R g518 ( 
.A(n_160),
.Y(n_518)
);

INVx1_ASAP7_75t_L g519 ( 
.A(n_291),
.Y(n_519)
);

CKINVDCx20_ASAP7_75t_R g520 ( 
.A(n_105),
.Y(n_520)
);

CKINVDCx5p33_ASAP7_75t_R g521 ( 
.A(n_241),
.Y(n_521)
);

CKINVDCx5p33_ASAP7_75t_R g522 ( 
.A(n_235),
.Y(n_522)
);

INVx1_ASAP7_75t_L g523 ( 
.A(n_179),
.Y(n_523)
);

CKINVDCx5p33_ASAP7_75t_R g524 ( 
.A(n_110),
.Y(n_524)
);

CKINVDCx5p33_ASAP7_75t_R g525 ( 
.A(n_228),
.Y(n_525)
);

INVx1_ASAP7_75t_L g526 ( 
.A(n_282),
.Y(n_526)
);

INVx1_ASAP7_75t_L g527 ( 
.A(n_109),
.Y(n_527)
);

INVx1_ASAP7_75t_L g528 ( 
.A(n_309),
.Y(n_528)
);

CKINVDCx5p33_ASAP7_75t_R g529 ( 
.A(n_92),
.Y(n_529)
);

CKINVDCx20_ASAP7_75t_R g530 ( 
.A(n_209),
.Y(n_530)
);

CKINVDCx5p33_ASAP7_75t_R g531 ( 
.A(n_388),
.Y(n_531)
);

CKINVDCx5p33_ASAP7_75t_R g532 ( 
.A(n_10),
.Y(n_532)
);

CKINVDCx5p33_ASAP7_75t_R g533 ( 
.A(n_151),
.Y(n_533)
);

INVx1_ASAP7_75t_L g534 ( 
.A(n_28),
.Y(n_534)
);

INVx1_ASAP7_75t_L g535 ( 
.A(n_94),
.Y(n_535)
);

CKINVDCx5p33_ASAP7_75t_R g536 ( 
.A(n_6),
.Y(n_536)
);

CKINVDCx5p33_ASAP7_75t_R g537 ( 
.A(n_281),
.Y(n_537)
);

INVx2_ASAP7_75t_SL g538 ( 
.A(n_61),
.Y(n_538)
);

INVx1_ASAP7_75t_L g539 ( 
.A(n_5),
.Y(n_539)
);

CKINVDCx5p33_ASAP7_75t_R g540 ( 
.A(n_365),
.Y(n_540)
);

CKINVDCx5p33_ASAP7_75t_R g541 ( 
.A(n_40),
.Y(n_541)
);

CKINVDCx16_ASAP7_75t_R g542 ( 
.A(n_73),
.Y(n_542)
);

CKINVDCx5p33_ASAP7_75t_R g543 ( 
.A(n_144),
.Y(n_543)
);

CKINVDCx20_ASAP7_75t_R g544 ( 
.A(n_25),
.Y(n_544)
);

CKINVDCx5p33_ASAP7_75t_R g545 ( 
.A(n_371),
.Y(n_545)
);

CKINVDCx5p33_ASAP7_75t_R g546 ( 
.A(n_89),
.Y(n_546)
);

INVx1_ASAP7_75t_L g547 ( 
.A(n_258),
.Y(n_547)
);

INVx2_ASAP7_75t_L g548 ( 
.A(n_57),
.Y(n_548)
);

CKINVDCx5p33_ASAP7_75t_R g549 ( 
.A(n_169),
.Y(n_549)
);

CKINVDCx5p33_ASAP7_75t_R g550 ( 
.A(n_4),
.Y(n_550)
);

BUFx10_ASAP7_75t_L g551 ( 
.A(n_264),
.Y(n_551)
);

CKINVDCx5p33_ASAP7_75t_R g552 ( 
.A(n_373),
.Y(n_552)
);

CKINVDCx5p33_ASAP7_75t_R g553 ( 
.A(n_23),
.Y(n_553)
);

CKINVDCx5p33_ASAP7_75t_R g554 ( 
.A(n_36),
.Y(n_554)
);

CKINVDCx5p33_ASAP7_75t_R g555 ( 
.A(n_370),
.Y(n_555)
);

CKINVDCx5p33_ASAP7_75t_R g556 ( 
.A(n_14),
.Y(n_556)
);

CKINVDCx5p33_ASAP7_75t_R g557 ( 
.A(n_21),
.Y(n_557)
);

CKINVDCx5p33_ASAP7_75t_R g558 ( 
.A(n_56),
.Y(n_558)
);

CKINVDCx5p33_ASAP7_75t_R g559 ( 
.A(n_42),
.Y(n_559)
);

CKINVDCx5p33_ASAP7_75t_R g560 ( 
.A(n_378),
.Y(n_560)
);

BUFx6f_ASAP7_75t_L g561 ( 
.A(n_294),
.Y(n_561)
);

CKINVDCx5p33_ASAP7_75t_R g562 ( 
.A(n_285),
.Y(n_562)
);

CKINVDCx5p33_ASAP7_75t_R g563 ( 
.A(n_260),
.Y(n_563)
);

CKINVDCx20_ASAP7_75t_R g564 ( 
.A(n_245),
.Y(n_564)
);

CKINVDCx5p33_ASAP7_75t_R g565 ( 
.A(n_156),
.Y(n_565)
);

INVx1_ASAP7_75t_L g566 ( 
.A(n_84),
.Y(n_566)
);

INVx1_ASAP7_75t_L g567 ( 
.A(n_172),
.Y(n_567)
);

CKINVDCx5p33_ASAP7_75t_R g568 ( 
.A(n_24),
.Y(n_568)
);

CKINVDCx16_ASAP7_75t_R g569 ( 
.A(n_363),
.Y(n_569)
);

CKINVDCx5p33_ASAP7_75t_R g570 ( 
.A(n_116),
.Y(n_570)
);

CKINVDCx20_ASAP7_75t_R g571 ( 
.A(n_246),
.Y(n_571)
);

CKINVDCx5p33_ASAP7_75t_R g572 ( 
.A(n_72),
.Y(n_572)
);

CKINVDCx5p33_ASAP7_75t_R g573 ( 
.A(n_31),
.Y(n_573)
);

CKINVDCx5p33_ASAP7_75t_R g574 ( 
.A(n_342),
.Y(n_574)
);

INVx1_ASAP7_75t_SL g575 ( 
.A(n_0),
.Y(n_575)
);

BUFx10_ASAP7_75t_L g576 ( 
.A(n_390),
.Y(n_576)
);

CKINVDCx5p33_ASAP7_75t_R g577 ( 
.A(n_237),
.Y(n_577)
);

CKINVDCx5p33_ASAP7_75t_R g578 ( 
.A(n_332),
.Y(n_578)
);

INVx1_ASAP7_75t_L g579 ( 
.A(n_77),
.Y(n_579)
);

INVx1_ASAP7_75t_L g580 ( 
.A(n_16),
.Y(n_580)
);

INVx1_ASAP7_75t_L g581 ( 
.A(n_366),
.Y(n_581)
);

INVx1_ASAP7_75t_L g582 ( 
.A(n_153),
.Y(n_582)
);

CKINVDCx5p33_ASAP7_75t_R g583 ( 
.A(n_322),
.Y(n_583)
);

INVx1_ASAP7_75t_L g584 ( 
.A(n_11),
.Y(n_584)
);

INVx1_ASAP7_75t_L g585 ( 
.A(n_152),
.Y(n_585)
);

CKINVDCx5p33_ASAP7_75t_R g586 ( 
.A(n_229),
.Y(n_586)
);

CKINVDCx5p33_ASAP7_75t_R g587 ( 
.A(n_95),
.Y(n_587)
);

INVx1_ASAP7_75t_L g588 ( 
.A(n_287),
.Y(n_588)
);

INVx1_ASAP7_75t_SL g589 ( 
.A(n_185),
.Y(n_589)
);

INVxp67_ASAP7_75t_L g590 ( 
.A(n_201),
.Y(n_590)
);

CKINVDCx5p33_ASAP7_75t_R g591 ( 
.A(n_34),
.Y(n_591)
);

CKINVDCx5p33_ASAP7_75t_R g592 ( 
.A(n_262),
.Y(n_592)
);

CKINVDCx5p33_ASAP7_75t_R g593 ( 
.A(n_191),
.Y(n_593)
);

CKINVDCx5p33_ASAP7_75t_R g594 ( 
.A(n_202),
.Y(n_594)
);

INVx1_ASAP7_75t_L g595 ( 
.A(n_203),
.Y(n_595)
);

INVx3_ASAP7_75t_L g596 ( 
.A(n_350),
.Y(n_596)
);

CKINVDCx5p33_ASAP7_75t_R g597 ( 
.A(n_227),
.Y(n_597)
);

CKINVDCx5p33_ASAP7_75t_R g598 ( 
.A(n_383),
.Y(n_598)
);

CKINVDCx5p33_ASAP7_75t_R g599 ( 
.A(n_106),
.Y(n_599)
);

INVx1_ASAP7_75t_L g600 ( 
.A(n_178),
.Y(n_600)
);

CKINVDCx5p33_ASAP7_75t_R g601 ( 
.A(n_45),
.Y(n_601)
);

CKINVDCx5p33_ASAP7_75t_R g602 ( 
.A(n_30),
.Y(n_602)
);

INVx1_ASAP7_75t_L g603 ( 
.A(n_238),
.Y(n_603)
);

CKINVDCx5p33_ASAP7_75t_R g604 ( 
.A(n_125),
.Y(n_604)
);

CKINVDCx5p33_ASAP7_75t_R g605 ( 
.A(n_341),
.Y(n_605)
);

INVx1_ASAP7_75t_L g606 ( 
.A(n_372),
.Y(n_606)
);

CKINVDCx5p33_ASAP7_75t_R g607 ( 
.A(n_340),
.Y(n_607)
);

CKINVDCx5p33_ASAP7_75t_R g608 ( 
.A(n_45),
.Y(n_608)
);

CKINVDCx5p33_ASAP7_75t_R g609 ( 
.A(n_112),
.Y(n_609)
);

INVx1_ASAP7_75t_L g610 ( 
.A(n_305),
.Y(n_610)
);

INVx1_ASAP7_75t_L g611 ( 
.A(n_221),
.Y(n_611)
);

BUFx3_ASAP7_75t_L g612 ( 
.A(n_43),
.Y(n_612)
);

INVxp67_ASAP7_75t_L g613 ( 
.A(n_358),
.Y(n_613)
);

BUFx6f_ASAP7_75t_L g614 ( 
.A(n_165),
.Y(n_614)
);

CKINVDCx5p33_ASAP7_75t_R g615 ( 
.A(n_310),
.Y(n_615)
);

INVx1_ASAP7_75t_L g616 ( 
.A(n_317),
.Y(n_616)
);

BUFx2_ASAP7_75t_L g617 ( 
.A(n_64),
.Y(n_617)
);

CKINVDCx5p33_ASAP7_75t_R g618 ( 
.A(n_129),
.Y(n_618)
);

INVx2_ASAP7_75t_L g619 ( 
.A(n_58),
.Y(n_619)
);

BUFx3_ASAP7_75t_L g620 ( 
.A(n_182),
.Y(n_620)
);

CKINVDCx20_ASAP7_75t_R g621 ( 
.A(n_19),
.Y(n_621)
);

BUFx2_ASAP7_75t_SL g622 ( 
.A(n_312),
.Y(n_622)
);

INVx1_ASAP7_75t_SL g623 ( 
.A(n_313),
.Y(n_623)
);

INVx1_ASAP7_75t_L g624 ( 
.A(n_81),
.Y(n_624)
);

CKINVDCx5p33_ASAP7_75t_R g625 ( 
.A(n_145),
.Y(n_625)
);

INVx1_ASAP7_75t_L g626 ( 
.A(n_35),
.Y(n_626)
);

INVx1_ASAP7_75t_L g627 ( 
.A(n_64),
.Y(n_627)
);

CKINVDCx5p33_ASAP7_75t_R g628 ( 
.A(n_297),
.Y(n_628)
);

CKINVDCx14_ASAP7_75t_R g629 ( 
.A(n_9),
.Y(n_629)
);

CKINVDCx5p33_ASAP7_75t_R g630 ( 
.A(n_168),
.Y(n_630)
);

CKINVDCx5p33_ASAP7_75t_R g631 ( 
.A(n_118),
.Y(n_631)
);

INVx1_ASAP7_75t_L g632 ( 
.A(n_102),
.Y(n_632)
);

CKINVDCx20_ASAP7_75t_R g633 ( 
.A(n_19),
.Y(n_633)
);

INVx1_ASAP7_75t_L g634 ( 
.A(n_131),
.Y(n_634)
);

CKINVDCx5p33_ASAP7_75t_R g635 ( 
.A(n_65),
.Y(n_635)
);

INVx1_ASAP7_75t_L g636 ( 
.A(n_356),
.Y(n_636)
);

INVx1_ASAP7_75t_L g637 ( 
.A(n_66),
.Y(n_637)
);

CKINVDCx5p33_ASAP7_75t_R g638 ( 
.A(n_65),
.Y(n_638)
);

CKINVDCx5p33_ASAP7_75t_R g639 ( 
.A(n_339),
.Y(n_639)
);

CKINVDCx5p33_ASAP7_75t_R g640 ( 
.A(n_38),
.Y(n_640)
);

CKINVDCx5p33_ASAP7_75t_R g641 ( 
.A(n_206),
.Y(n_641)
);

BUFx10_ASAP7_75t_L g642 ( 
.A(n_263),
.Y(n_642)
);

INVx1_ASAP7_75t_L g643 ( 
.A(n_53),
.Y(n_643)
);

CKINVDCx5p33_ASAP7_75t_R g644 ( 
.A(n_355),
.Y(n_644)
);

INVx1_ASAP7_75t_L g645 ( 
.A(n_74),
.Y(n_645)
);

INVx1_ASAP7_75t_L g646 ( 
.A(n_349),
.Y(n_646)
);

INVx1_ASAP7_75t_L g647 ( 
.A(n_391),
.Y(n_647)
);

INVx1_ASAP7_75t_L g648 ( 
.A(n_111),
.Y(n_648)
);

INVx2_ASAP7_75t_L g649 ( 
.A(n_345),
.Y(n_649)
);

CKINVDCx14_ASAP7_75t_R g650 ( 
.A(n_239),
.Y(n_650)
);

CKINVDCx20_ASAP7_75t_R g651 ( 
.A(n_385),
.Y(n_651)
);

CKINVDCx20_ASAP7_75t_R g652 ( 
.A(n_189),
.Y(n_652)
);

CKINVDCx5p33_ASAP7_75t_R g653 ( 
.A(n_324),
.Y(n_653)
);

CKINVDCx5p33_ASAP7_75t_R g654 ( 
.A(n_230),
.Y(n_654)
);

CKINVDCx5p33_ASAP7_75t_R g655 ( 
.A(n_81),
.Y(n_655)
);

INVx1_ASAP7_75t_L g656 ( 
.A(n_84),
.Y(n_656)
);

BUFx10_ASAP7_75t_L g657 ( 
.A(n_249),
.Y(n_657)
);

CKINVDCx5p33_ASAP7_75t_R g658 ( 
.A(n_384),
.Y(n_658)
);

INVx1_ASAP7_75t_L g659 ( 
.A(n_173),
.Y(n_659)
);

BUFx2_ASAP7_75t_L g660 ( 
.A(n_316),
.Y(n_660)
);

CKINVDCx5p33_ASAP7_75t_R g661 ( 
.A(n_91),
.Y(n_661)
);

CKINVDCx5p33_ASAP7_75t_R g662 ( 
.A(n_334),
.Y(n_662)
);

INVx1_ASAP7_75t_L g663 ( 
.A(n_70),
.Y(n_663)
);

CKINVDCx5p33_ASAP7_75t_R g664 ( 
.A(n_158),
.Y(n_664)
);

CKINVDCx5p33_ASAP7_75t_R g665 ( 
.A(n_368),
.Y(n_665)
);

BUFx6f_ASAP7_75t_L g666 ( 
.A(n_273),
.Y(n_666)
);

INVx1_ASAP7_75t_L g667 ( 
.A(n_1),
.Y(n_667)
);

INVx1_ASAP7_75t_L g668 ( 
.A(n_318),
.Y(n_668)
);

CKINVDCx14_ASAP7_75t_R g669 ( 
.A(n_284),
.Y(n_669)
);

CKINVDCx5p33_ASAP7_75t_R g670 ( 
.A(n_213),
.Y(n_670)
);

CKINVDCx5p33_ASAP7_75t_R g671 ( 
.A(n_346),
.Y(n_671)
);

CKINVDCx5p33_ASAP7_75t_R g672 ( 
.A(n_46),
.Y(n_672)
);

CKINVDCx5p33_ASAP7_75t_R g673 ( 
.A(n_381),
.Y(n_673)
);

CKINVDCx5p33_ASAP7_75t_R g674 ( 
.A(n_325),
.Y(n_674)
);

CKINVDCx5p33_ASAP7_75t_R g675 ( 
.A(n_335),
.Y(n_675)
);

INVx3_ASAP7_75t_L g676 ( 
.A(n_269),
.Y(n_676)
);

CKINVDCx5p33_ASAP7_75t_R g677 ( 
.A(n_320),
.Y(n_677)
);

CKINVDCx5p33_ASAP7_75t_R g678 ( 
.A(n_137),
.Y(n_678)
);

INVx1_ASAP7_75t_L g679 ( 
.A(n_351),
.Y(n_679)
);

CKINVDCx5p33_ASAP7_75t_R g680 ( 
.A(n_331),
.Y(n_680)
);

CKINVDCx5p33_ASAP7_75t_R g681 ( 
.A(n_343),
.Y(n_681)
);

INVx1_ASAP7_75t_L g682 ( 
.A(n_50),
.Y(n_682)
);

CKINVDCx5p33_ASAP7_75t_R g683 ( 
.A(n_193),
.Y(n_683)
);

CKINVDCx5p33_ASAP7_75t_R g684 ( 
.A(n_150),
.Y(n_684)
);

CKINVDCx5p33_ASAP7_75t_R g685 ( 
.A(n_323),
.Y(n_685)
);

CKINVDCx5p33_ASAP7_75t_R g686 ( 
.A(n_376),
.Y(n_686)
);

CKINVDCx20_ASAP7_75t_R g687 ( 
.A(n_244),
.Y(n_687)
);

CKINVDCx5p33_ASAP7_75t_R g688 ( 
.A(n_330),
.Y(n_688)
);

INVx1_ASAP7_75t_L g689 ( 
.A(n_194),
.Y(n_689)
);

CKINVDCx5p33_ASAP7_75t_R g690 ( 
.A(n_359),
.Y(n_690)
);

CKINVDCx20_ASAP7_75t_R g691 ( 
.A(n_74),
.Y(n_691)
);

BUFx6f_ASAP7_75t_L g692 ( 
.A(n_46),
.Y(n_692)
);

CKINVDCx5p33_ASAP7_75t_R g693 ( 
.A(n_314),
.Y(n_693)
);

CKINVDCx5p33_ASAP7_75t_R g694 ( 
.A(n_42),
.Y(n_694)
);

CKINVDCx5p33_ASAP7_75t_R g695 ( 
.A(n_80),
.Y(n_695)
);

CKINVDCx5p33_ASAP7_75t_R g696 ( 
.A(n_163),
.Y(n_696)
);

CKINVDCx5p33_ASAP7_75t_R g697 ( 
.A(n_256),
.Y(n_697)
);

CKINVDCx20_ASAP7_75t_R g698 ( 
.A(n_98),
.Y(n_698)
);

INVx2_ASAP7_75t_L g699 ( 
.A(n_394),
.Y(n_699)
);

CKINVDCx5p33_ASAP7_75t_R g700 ( 
.A(n_3),
.Y(n_700)
);

CKINVDCx5p33_ASAP7_75t_R g701 ( 
.A(n_357),
.Y(n_701)
);

CKINVDCx5p33_ASAP7_75t_R g702 ( 
.A(n_180),
.Y(n_702)
);

HB1xp67_ASAP7_75t_L g703 ( 
.A(n_188),
.Y(n_703)
);

CKINVDCx5p33_ASAP7_75t_R g704 ( 
.A(n_135),
.Y(n_704)
);

INVx1_ASAP7_75t_L g705 ( 
.A(n_184),
.Y(n_705)
);

CKINVDCx5p33_ASAP7_75t_R g706 ( 
.A(n_270),
.Y(n_706)
);

CKINVDCx5p33_ASAP7_75t_R g707 ( 
.A(n_155),
.Y(n_707)
);

BUFx3_ASAP7_75t_L g708 ( 
.A(n_39),
.Y(n_708)
);

BUFx10_ASAP7_75t_L g709 ( 
.A(n_77),
.Y(n_709)
);

CKINVDCx5p33_ASAP7_75t_R g710 ( 
.A(n_252),
.Y(n_710)
);

INVx1_ASAP7_75t_L g711 ( 
.A(n_283),
.Y(n_711)
);

CKINVDCx5p33_ASAP7_75t_R g712 ( 
.A(n_128),
.Y(n_712)
);

CKINVDCx5p33_ASAP7_75t_R g713 ( 
.A(n_52),
.Y(n_713)
);

INVx1_ASAP7_75t_SL g714 ( 
.A(n_55),
.Y(n_714)
);

CKINVDCx5p33_ASAP7_75t_R g715 ( 
.A(n_51),
.Y(n_715)
);

CKINVDCx5p33_ASAP7_75t_R g716 ( 
.A(n_17),
.Y(n_716)
);

CKINVDCx16_ASAP7_75t_R g717 ( 
.A(n_308),
.Y(n_717)
);

INVx2_ASAP7_75t_L g718 ( 
.A(n_377),
.Y(n_718)
);

CKINVDCx5p33_ASAP7_75t_R g719 ( 
.A(n_102),
.Y(n_719)
);

INVx1_ASAP7_75t_L g720 ( 
.A(n_328),
.Y(n_720)
);

INVx1_ASAP7_75t_L g721 ( 
.A(n_289),
.Y(n_721)
);

INVx1_ASAP7_75t_L g722 ( 
.A(n_329),
.Y(n_722)
);

INVx1_ASAP7_75t_L g723 ( 
.A(n_57),
.Y(n_723)
);

CKINVDCx5p33_ASAP7_75t_R g724 ( 
.A(n_250),
.Y(n_724)
);

CKINVDCx5p33_ASAP7_75t_R g725 ( 
.A(n_304),
.Y(n_725)
);

CKINVDCx5p33_ASAP7_75t_R g726 ( 
.A(n_353),
.Y(n_726)
);

INVx2_ASAP7_75t_SL g727 ( 
.A(n_379),
.Y(n_727)
);

INVx1_ASAP7_75t_L g728 ( 
.A(n_138),
.Y(n_728)
);

CKINVDCx5p33_ASAP7_75t_R g729 ( 
.A(n_56),
.Y(n_729)
);

CKINVDCx5p33_ASAP7_75t_R g730 ( 
.A(n_199),
.Y(n_730)
);

CKINVDCx5p33_ASAP7_75t_R g731 ( 
.A(n_255),
.Y(n_731)
);

INVx1_ASAP7_75t_L g732 ( 
.A(n_440),
.Y(n_732)
);

CKINVDCx5p33_ASAP7_75t_R g733 ( 
.A(n_542),
.Y(n_733)
);

INVx1_ASAP7_75t_L g734 ( 
.A(n_440),
.Y(n_734)
);

INVx1_ASAP7_75t_L g735 ( 
.A(n_500),
.Y(n_735)
);

CKINVDCx5p33_ASAP7_75t_R g736 ( 
.A(n_429),
.Y(n_736)
);

INVx1_ASAP7_75t_L g737 ( 
.A(n_500),
.Y(n_737)
);

INVx1_ASAP7_75t_L g738 ( 
.A(n_501),
.Y(n_738)
);

INVx1_ASAP7_75t_L g739 ( 
.A(n_501),
.Y(n_739)
);

INVx1_ASAP7_75t_L g740 ( 
.A(n_612),
.Y(n_740)
);

INVx1_ASAP7_75t_L g741 ( 
.A(n_612),
.Y(n_741)
);

INVx1_ASAP7_75t_L g742 ( 
.A(n_708),
.Y(n_742)
);

CKINVDCx16_ASAP7_75t_R g743 ( 
.A(n_629),
.Y(n_743)
);

INVx1_ASAP7_75t_L g744 ( 
.A(n_708),
.Y(n_744)
);

INVx1_ASAP7_75t_L g745 ( 
.A(n_439),
.Y(n_745)
);

INVxp67_ASAP7_75t_SL g746 ( 
.A(n_426),
.Y(n_746)
);

INVx1_ASAP7_75t_L g747 ( 
.A(n_439),
.Y(n_747)
);

INVx1_ASAP7_75t_L g748 ( 
.A(n_439),
.Y(n_748)
);

INVxp67_ASAP7_75t_SL g749 ( 
.A(n_426),
.Y(n_749)
);

INVxp33_ASAP7_75t_SL g750 ( 
.A(n_488),
.Y(n_750)
);

INVxp67_ASAP7_75t_SL g751 ( 
.A(n_511),
.Y(n_751)
);

INVx1_ASAP7_75t_L g752 ( 
.A(n_439),
.Y(n_752)
);

INVx1_ASAP7_75t_L g753 ( 
.A(n_439),
.Y(n_753)
);

INVx1_ASAP7_75t_L g754 ( 
.A(n_439),
.Y(n_754)
);

CKINVDCx20_ASAP7_75t_R g755 ( 
.A(n_629),
.Y(n_755)
);

INVx1_ASAP7_75t_L g756 ( 
.A(n_439),
.Y(n_756)
);

INVx1_ASAP7_75t_L g757 ( 
.A(n_395),
.Y(n_757)
);

INVx1_ASAP7_75t_L g758 ( 
.A(n_414),
.Y(n_758)
);

INVxp67_ASAP7_75t_L g759 ( 
.A(n_617),
.Y(n_759)
);

BUFx5_ASAP7_75t_L g760 ( 
.A(n_406),
.Y(n_760)
);

BUFx3_ASAP7_75t_L g761 ( 
.A(n_660),
.Y(n_761)
);

INVx1_ASAP7_75t_L g762 ( 
.A(n_417),
.Y(n_762)
);

INVx1_ASAP7_75t_L g763 ( 
.A(n_430),
.Y(n_763)
);

CKINVDCx16_ASAP7_75t_R g764 ( 
.A(n_418),
.Y(n_764)
);

INVx1_ASAP7_75t_L g765 ( 
.A(n_432),
.Y(n_765)
);

INVx2_ASAP7_75t_L g766 ( 
.A(n_692),
.Y(n_766)
);

INVx1_ASAP7_75t_L g767 ( 
.A(n_434),
.Y(n_767)
);

INVxp67_ASAP7_75t_L g768 ( 
.A(n_511),
.Y(n_768)
);

CKINVDCx20_ASAP7_75t_R g769 ( 
.A(n_427),
.Y(n_769)
);

INVx1_ASAP7_75t_L g770 ( 
.A(n_435),
.Y(n_770)
);

INVxp67_ASAP7_75t_L g771 ( 
.A(n_548),
.Y(n_771)
);

INVx1_ASAP7_75t_L g772 ( 
.A(n_464),
.Y(n_772)
);

INVx1_ASAP7_75t_L g773 ( 
.A(n_475),
.Y(n_773)
);

CKINVDCx16_ASAP7_75t_R g774 ( 
.A(n_465),
.Y(n_774)
);

INVx1_ASAP7_75t_L g775 ( 
.A(n_479),
.Y(n_775)
);

INVx2_ASAP7_75t_L g776 ( 
.A(n_692),
.Y(n_776)
);

INVxp33_ASAP7_75t_L g777 ( 
.A(n_548),
.Y(n_777)
);

INVxp67_ASAP7_75t_SL g778 ( 
.A(n_619),
.Y(n_778)
);

INVxp33_ASAP7_75t_L g779 ( 
.A(n_481),
.Y(n_779)
);

INVx1_ASAP7_75t_L g780 ( 
.A(n_508),
.Y(n_780)
);

INVxp33_ASAP7_75t_L g781 ( 
.A(n_515),
.Y(n_781)
);

INVx1_ASAP7_75t_L g782 ( 
.A(n_534),
.Y(n_782)
);

INVx1_ASAP7_75t_L g783 ( 
.A(n_535),
.Y(n_783)
);

INVx1_ASAP7_75t_L g784 ( 
.A(n_539),
.Y(n_784)
);

CKINVDCx5p33_ASAP7_75t_R g785 ( 
.A(n_437),
.Y(n_785)
);

INVx1_ASAP7_75t_L g786 ( 
.A(n_566),
.Y(n_786)
);

INVxp67_ASAP7_75t_SL g787 ( 
.A(n_619),
.Y(n_787)
);

INVx2_ASAP7_75t_L g788 ( 
.A(n_692),
.Y(n_788)
);

INVx2_ASAP7_75t_L g789 ( 
.A(n_692),
.Y(n_789)
);

INVx3_ASAP7_75t_L g790 ( 
.A(n_443),
.Y(n_790)
);

CKINVDCx20_ASAP7_75t_R g791 ( 
.A(n_427),
.Y(n_791)
);

INVxp67_ASAP7_75t_SL g792 ( 
.A(n_579),
.Y(n_792)
);

INVx2_ASAP7_75t_L g793 ( 
.A(n_402),
.Y(n_793)
);

INVx1_ASAP7_75t_L g794 ( 
.A(n_580),
.Y(n_794)
);

INVxp33_ASAP7_75t_SL g795 ( 
.A(n_405),
.Y(n_795)
);

INVx1_ASAP7_75t_L g796 ( 
.A(n_584),
.Y(n_796)
);

INVx1_ASAP7_75t_L g797 ( 
.A(n_624),
.Y(n_797)
);

INVxp67_ASAP7_75t_SL g798 ( 
.A(n_626),
.Y(n_798)
);

INVxp33_ASAP7_75t_L g799 ( 
.A(n_627),
.Y(n_799)
);

BUFx3_ASAP7_75t_L g800 ( 
.A(n_512),
.Y(n_800)
);

INVx1_ASAP7_75t_L g801 ( 
.A(n_632),
.Y(n_801)
);

CKINVDCx14_ASAP7_75t_R g802 ( 
.A(n_650),
.Y(n_802)
);

INVx1_ASAP7_75t_L g803 ( 
.A(n_637),
.Y(n_803)
);

INVx2_ASAP7_75t_L g804 ( 
.A(n_402),
.Y(n_804)
);

INVxp33_ASAP7_75t_SL g805 ( 
.A(n_409),
.Y(n_805)
);

INVx1_ASAP7_75t_L g806 ( 
.A(n_643),
.Y(n_806)
);

INVx1_ASAP7_75t_L g807 ( 
.A(n_645),
.Y(n_807)
);

INVx2_ASAP7_75t_L g808 ( 
.A(n_620),
.Y(n_808)
);

INVx2_ASAP7_75t_L g809 ( 
.A(n_620),
.Y(n_809)
);

INVx1_ASAP7_75t_L g810 ( 
.A(n_656),
.Y(n_810)
);

CKINVDCx5p33_ASAP7_75t_R g811 ( 
.A(n_520),
.Y(n_811)
);

INVx1_ASAP7_75t_L g812 ( 
.A(n_663),
.Y(n_812)
);

CKINVDCx16_ASAP7_75t_R g813 ( 
.A(n_569),
.Y(n_813)
);

INVx1_ASAP7_75t_L g814 ( 
.A(n_667),
.Y(n_814)
);

INVx1_ASAP7_75t_L g815 ( 
.A(n_682),
.Y(n_815)
);

INVx1_ASAP7_75t_L g816 ( 
.A(n_723),
.Y(n_816)
);

INVx1_ASAP7_75t_L g817 ( 
.A(n_506),
.Y(n_817)
);

CKINVDCx5p33_ASAP7_75t_R g818 ( 
.A(n_530),
.Y(n_818)
);

INVx1_ASAP7_75t_L g819 ( 
.A(n_703),
.Y(n_819)
);

INVx1_ASAP7_75t_L g820 ( 
.A(n_538),
.Y(n_820)
);

INVx1_ASAP7_75t_L g821 ( 
.A(n_512),
.Y(n_821)
);

CKINVDCx5p33_ASAP7_75t_R g822 ( 
.A(n_423),
.Y(n_822)
);

INVx1_ASAP7_75t_L g823 ( 
.A(n_512),
.Y(n_823)
);

INVx1_ASAP7_75t_L g824 ( 
.A(n_551),
.Y(n_824)
);

INVx1_ASAP7_75t_L g825 ( 
.A(n_551),
.Y(n_825)
);

INVx1_ASAP7_75t_L g826 ( 
.A(n_551),
.Y(n_826)
);

CKINVDCx5p33_ASAP7_75t_R g827 ( 
.A(n_433),
.Y(n_827)
);

CKINVDCx20_ASAP7_75t_R g828 ( 
.A(n_564),
.Y(n_828)
);

INVxp67_ASAP7_75t_SL g829 ( 
.A(n_596),
.Y(n_829)
);

INVx1_ASAP7_75t_L g830 ( 
.A(n_576),
.Y(n_830)
);

CKINVDCx20_ASAP7_75t_R g831 ( 
.A(n_564),
.Y(n_831)
);

INVx2_ASAP7_75t_SL g832 ( 
.A(n_443),
.Y(n_832)
);

INVx1_ASAP7_75t_L g833 ( 
.A(n_576),
.Y(n_833)
);

INVx1_ASAP7_75t_L g834 ( 
.A(n_576),
.Y(n_834)
);

INVx1_ASAP7_75t_L g835 ( 
.A(n_642),
.Y(n_835)
);

INVxp67_ASAP7_75t_L g836 ( 
.A(n_443),
.Y(n_836)
);

INVx1_ASAP7_75t_L g837 ( 
.A(n_642),
.Y(n_837)
);

XNOR2xp5_ASAP7_75t_L g838 ( 
.A(n_422),
.B(n_2),
.Y(n_838)
);

INVxp67_ASAP7_75t_L g839 ( 
.A(n_709),
.Y(n_839)
);

CKINVDCx5p33_ASAP7_75t_R g840 ( 
.A(n_441),
.Y(n_840)
);

INVx1_ASAP7_75t_L g841 ( 
.A(n_642),
.Y(n_841)
);

NOR2xp67_ASAP7_75t_L g842 ( 
.A(n_596),
.B(n_6),
.Y(n_842)
);

INVx1_ASAP7_75t_L g843 ( 
.A(n_657),
.Y(n_843)
);

INVx1_ASAP7_75t_L g844 ( 
.A(n_657),
.Y(n_844)
);

INVx1_ASAP7_75t_L g845 ( 
.A(n_657),
.Y(n_845)
);

INVx1_ASAP7_75t_L g846 ( 
.A(n_709),
.Y(n_846)
);

INVx1_ASAP7_75t_L g847 ( 
.A(n_709),
.Y(n_847)
);

INVx1_ASAP7_75t_L g848 ( 
.A(n_407),
.Y(n_848)
);

INVx1_ASAP7_75t_L g849 ( 
.A(n_410),
.Y(n_849)
);

INVxp67_ASAP7_75t_SL g850 ( 
.A(n_596),
.Y(n_850)
);

BUFx10_ASAP7_75t_L g851 ( 
.A(n_457),
.Y(n_851)
);

CKINVDCx20_ASAP7_75t_R g852 ( 
.A(n_571),
.Y(n_852)
);

INVxp67_ASAP7_75t_SL g853 ( 
.A(n_676),
.Y(n_853)
);

CKINVDCx5p33_ASAP7_75t_R g854 ( 
.A(n_458),
.Y(n_854)
);

INVx1_ASAP7_75t_L g855 ( 
.A(n_411),
.Y(n_855)
);

INVx1_ASAP7_75t_L g856 ( 
.A(n_413),
.Y(n_856)
);

CKINVDCx20_ASAP7_75t_R g857 ( 
.A(n_571),
.Y(n_857)
);

INVxp33_ASAP7_75t_L g858 ( 
.A(n_398),
.Y(n_858)
);

INVx1_ASAP7_75t_L g859 ( 
.A(n_424),
.Y(n_859)
);

CKINVDCx5p33_ASAP7_75t_R g860 ( 
.A(n_468),
.Y(n_860)
);

BUFx6f_ASAP7_75t_L g861 ( 
.A(n_496),
.Y(n_861)
);

CKINVDCx5p33_ASAP7_75t_R g862 ( 
.A(n_469),
.Y(n_862)
);

INVx1_ASAP7_75t_L g863 ( 
.A(n_446),
.Y(n_863)
);

INVx1_ASAP7_75t_L g864 ( 
.A(n_447),
.Y(n_864)
);

INVx1_ASAP7_75t_L g865 ( 
.A(n_448),
.Y(n_865)
);

INVx1_ASAP7_75t_L g866 ( 
.A(n_451),
.Y(n_866)
);

INVxp33_ASAP7_75t_L g867 ( 
.A(n_398),
.Y(n_867)
);

BUFx3_ASAP7_75t_L g868 ( 
.A(n_454),
.Y(n_868)
);

INVx1_ASAP7_75t_L g869 ( 
.A(n_456),
.Y(n_869)
);

CKINVDCx20_ASAP7_75t_R g870 ( 
.A(n_651),
.Y(n_870)
);

INVx2_ASAP7_75t_L g871 ( 
.A(n_463),
.Y(n_871)
);

INVx1_ASAP7_75t_L g872 ( 
.A(n_471),
.Y(n_872)
);

INVx2_ASAP7_75t_L g873 ( 
.A(n_472),
.Y(n_873)
);

INVx1_ASAP7_75t_L g874 ( 
.A(n_482),
.Y(n_874)
);

CKINVDCx5p33_ASAP7_75t_R g875 ( 
.A(n_473),
.Y(n_875)
);

INVx1_ASAP7_75t_L g876 ( 
.A(n_486),
.Y(n_876)
);

INVx1_ASAP7_75t_L g877 ( 
.A(n_489),
.Y(n_877)
);

CKINVDCx5p33_ASAP7_75t_R g878 ( 
.A(n_493),
.Y(n_878)
);

INVx1_ASAP7_75t_L g879 ( 
.A(n_492),
.Y(n_879)
);

INVxp33_ASAP7_75t_SL g880 ( 
.A(n_498),
.Y(n_880)
);

INVxp67_ASAP7_75t_SL g881 ( 
.A(n_676),
.Y(n_881)
);

INVx1_ASAP7_75t_L g882 ( 
.A(n_495),
.Y(n_882)
);

INVxp33_ASAP7_75t_L g883 ( 
.A(n_452),
.Y(n_883)
);

INVx1_ASAP7_75t_L g884 ( 
.A(n_502),
.Y(n_884)
);

CKINVDCx20_ASAP7_75t_R g885 ( 
.A(n_651),
.Y(n_885)
);

HB1xp67_ASAP7_75t_L g886 ( 
.A(n_499),
.Y(n_886)
);

INVx2_ASAP7_75t_L g887 ( 
.A(n_505),
.Y(n_887)
);

INVx1_ASAP7_75t_L g888 ( 
.A(n_514),
.Y(n_888)
);

INVx2_ASAP7_75t_L g889 ( 
.A(n_519),
.Y(n_889)
);

NOR2xp67_ASAP7_75t_L g890 ( 
.A(n_676),
.B(n_7),
.Y(n_890)
);

INVx1_ASAP7_75t_L g891 ( 
.A(n_523),
.Y(n_891)
);

INVxp67_ASAP7_75t_SL g892 ( 
.A(n_452),
.Y(n_892)
);

BUFx3_ASAP7_75t_L g893 ( 
.A(n_526),
.Y(n_893)
);

INVx1_ASAP7_75t_L g894 ( 
.A(n_527),
.Y(n_894)
);

INVxp33_ASAP7_75t_L g895 ( 
.A(n_459),
.Y(n_895)
);

BUFx6f_ASAP7_75t_L g896 ( 
.A(n_496),
.Y(n_896)
);

INVx1_ASAP7_75t_L g897 ( 
.A(n_528),
.Y(n_897)
);

INVx3_ASAP7_75t_L g898 ( 
.A(n_503),
.Y(n_898)
);

CKINVDCx5p33_ASAP7_75t_R g899 ( 
.A(n_507),
.Y(n_899)
);

CKINVDCx5p33_ASAP7_75t_R g900 ( 
.A(n_509),
.Y(n_900)
);

INVx1_ASAP7_75t_L g901 ( 
.A(n_547),
.Y(n_901)
);

INVx1_ASAP7_75t_L g902 ( 
.A(n_567),
.Y(n_902)
);

INVx1_ASAP7_75t_L g903 ( 
.A(n_581),
.Y(n_903)
);

INVx1_ASAP7_75t_L g904 ( 
.A(n_582),
.Y(n_904)
);

INVxp33_ASAP7_75t_SL g905 ( 
.A(n_516),
.Y(n_905)
);

INVxp33_ASAP7_75t_L g906 ( 
.A(n_459),
.Y(n_906)
);

INVx2_ASAP7_75t_L g907 ( 
.A(n_585),
.Y(n_907)
);

INVxp67_ASAP7_75t_SL g908 ( 
.A(n_462),
.Y(n_908)
);

INVx1_ASAP7_75t_L g909 ( 
.A(n_588),
.Y(n_909)
);

INVx1_ASAP7_75t_L g910 ( 
.A(n_595),
.Y(n_910)
);

INVxp33_ASAP7_75t_SL g911 ( 
.A(n_529),
.Y(n_911)
);

INVx1_ASAP7_75t_L g912 ( 
.A(n_600),
.Y(n_912)
);

INVx1_ASAP7_75t_L g913 ( 
.A(n_603),
.Y(n_913)
);

INVx1_ASAP7_75t_L g914 ( 
.A(n_606),
.Y(n_914)
);

BUFx6f_ASAP7_75t_L g915 ( 
.A(n_496),
.Y(n_915)
);

INVx1_ASAP7_75t_L g916 ( 
.A(n_610),
.Y(n_916)
);

INVx1_ASAP7_75t_L g917 ( 
.A(n_611),
.Y(n_917)
);

INVx1_ASAP7_75t_L g918 ( 
.A(n_616),
.Y(n_918)
);

INVxp67_ASAP7_75t_SL g919 ( 
.A(n_462),
.Y(n_919)
);

INVx1_ASAP7_75t_L g920 ( 
.A(n_634),
.Y(n_920)
);

INVx1_ASAP7_75t_L g921 ( 
.A(n_636),
.Y(n_921)
);

INVxp67_ASAP7_75t_SL g922 ( 
.A(n_649),
.Y(n_922)
);

INVx1_ASAP7_75t_SL g923 ( 
.A(n_483),
.Y(n_923)
);

INVxp33_ASAP7_75t_L g924 ( 
.A(n_649),
.Y(n_924)
);

INVx1_ASAP7_75t_L g925 ( 
.A(n_646),
.Y(n_925)
);

INVx1_ASAP7_75t_L g926 ( 
.A(n_647),
.Y(n_926)
);

INVxp67_ASAP7_75t_SL g927 ( 
.A(n_699),
.Y(n_927)
);

CKINVDCx20_ASAP7_75t_R g928 ( 
.A(n_652),
.Y(n_928)
);

INVxp33_ASAP7_75t_L g929 ( 
.A(n_699),
.Y(n_929)
);

INVx1_ASAP7_75t_L g930 ( 
.A(n_648),
.Y(n_930)
);

INVx1_ASAP7_75t_L g931 ( 
.A(n_659),
.Y(n_931)
);

INVx1_ASAP7_75t_L g932 ( 
.A(n_668),
.Y(n_932)
);

CKINVDCx20_ASAP7_75t_R g933 ( 
.A(n_652),
.Y(n_933)
);

INVxp67_ASAP7_75t_SL g934 ( 
.A(n_718),
.Y(n_934)
);

INVx1_ASAP7_75t_L g935 ( 
.A(n_679),
.Y(n_935)
);

INVx1_ASAP7_75t_L g936 ( 
.A(n_689),
.Y(n_936)
);

INVx2_ASAP7_75t_L g937 ( 
.A(n_705),
.Y(n_937)
);

INVx1_ASAP7_75t_L g938 ( 
.A(n_711),
.Y(n_938)
);

INVx1_ASAP7_75t_L g939 ( 
.A(n_720),
.Y(n_939)
);

INVx2_ASAP7_75t_L g940 ( 
.A(n_721),
.Y(n_940)
);

INVx1_ASAP7_75t_L g941 ( 
.A(n_722),
.Y(n_941)
);

INVx1_ASAP7_75t_L g942 ( 
.A(n_728),
.Y(n_942)
);

BUFx3_ASAP7_75t_L g943 ( 
.A(n_396),
.Y(n_943)
);

INVx2_ASAP7_75t_L g944 ( 
.A(n_718),
.Y(n_944)
);

INVx1_ASAP7_75t_L g945 ( 
.A(n_513),
.Y(n_945)
);

INVx1_ASAP7_75t_L g946 ( 
.A(n_532),
.Y(n_946)
);

INVx1_ASAP7_75t_L g947 ( 
.A(n_536),
.Y(n_947)
);

INVx1_ASAP7_75t_L g948 ( 
.A(n_541),
.Y(n_948)
);

INVx2_ASAP7_75t_L g949 ( 
.A(n_727),
.Y(n_949)
);

INVx1_ASAP7_75t_L g950 ( 
.A(n_546),
.Y(n_950)
);

INVx2_ASAP7_75t_L g951 ( 
.A(n_496),
.Y(n_951)
);

INVx1_ASAP7_75t_L g952 ( 
.A(n_550),
.Y(n_952)
);

INVx1_ASAP7_75t_L g953 ( 
.A(n_553),
.Y(n_953)
);

INVxp67_ASAP7_75t_SL g954 ( 
.A(n_450),
.Y(n_954)
);

INVx1_ASAP7_75t_L g955 ( 
.A(n_554),
.Y(n_955)
);

BUFx6f_ASAP7_75t_L g956 ( 
.A(n_561),
.Y(n_956)
);

INVxp67_ASAP7_75t_SL g957 ( 
.A(n_590),
.Y(n_957)
);

INVx1_ASAP7_75t_L g958 ( 
.A(n_556),
.Y(n_958)
);

INVxp33_ASAP7_75t_SL g959 ( 
.A(n_557),
.Y(n_959)
);

INVx1_ASAP7_75t_L g960 ( 
.A(n_558),
.Y(n_960)
);

INVx1_ASAP7_75t_L g961 ( 
.A(n_559),
.Y(n_961)
);

INVx1_ASAP7_75t_L g962 ( 
.A(n_568),
.Y(n_962)
);

CKINVDCx20_ASAP7_75t_R g963 ( 
.A(n_687),
.Y(n_963)
);

INVx1_ASAP7_75t_L g964 ( 
.A(n_572),
.Y(n_964)
);

INVx1_ASAP7_75t_L g965 ( 
.A(n_573),
.Y(n_965)
);

INVx1_ASAP7_75t_L g966 ( 
.A(n_587),
.Y(n_966)
);

INVx1_ASAP7_75t_L g967 ( 
.A(n_591),
.Y(n_967)
);

INVx1_ASAP7_75t_L g968 ( 
.A(n_601),
.Y(n_968)
);

CKINVDCx20_ASAP7_75t_R g969 ( 
.A(n_687),
.Y(n_969)
);

INVx1_ASAP7_75t_L g970 ( 
.A(n_602),
.Y(n_970)
);

INVxp67_ASAP7_75t_L g971 ( 
.A(n_608),
.Y(n_971)
);

CKINVDCx20_ASAP7_75t_R g972 ( 
.A(n_422),
.Y(n_972)
);

INVx1_ASAP7_75t_L g973 ( 
.A(n_635),
.Y(n_973)
);

INVx1_ASAP7_75t_L g974 ( 
.A(n_638),
.Y(n_974)
);

INVx1_ASAP7_75t_L g975 ( 
.A(n_640),
.Y(n_975)
);

INVx1_ASAP7_75t_L g976 ( 
.A(n_655),
.Y(n_976)
);

INVxp67_ASAP7_75t_L g977 ( 
.A(n_661),
.Y(n_977)
);

INVx2_ASAP7_75t_L g978 ( 
.A(n_561),
.Y(n_978)
);

INVxp33_ASAP7_75t_L g979 ( 
.A(n_544),
.Y(n_979)
);

INVx2_ASAP7_75t_L g980 ( 
.A(n_561),
.Y(n_980)
);

INVx1_ASAP7_75t_L g981 ( 
.A(n_672),
.Y(n_981)
);

CKINVDCx20_ASAP7_75t_R g982 ( 
.A(n_544),
.Y(n_982)
);

INVx1_ASAP7_75t_L g983 ( 
.A(n_694),
.Y(n_983)
);

INVxp67_ASAP7_75t_SL g984 ( 
.A(n_613),
.Y(n_984)
);

INVx1_ASAP7_75t_L g985 ( 
.A(n_695),
.Y(n_985)
);

INVx1_ASAP7_75t_L g986 ( 
.A(n_700),
.Y(n_986)
);

INVxp67_ASAP7_75t_L g987 ( 
.A(n_713),
.Y(n_987)
);

INVx1_ASAP7_75t_L g988 ( 
.A(n_715),
.Y(n_988)
);

CKINVDCx20_ASAP7_75t_R g989 ( 
.A(n_621),
.Y(n_989)
);

INVx1_ASAP7_75t_L g990 ( 
.A(n_716),
.Y(n_990)
);

INVx1_ASAP7_75t_L g991 ( 
.A(n_719),
.Y(n_991)
);

CKINVDCx5p33_ASAP7_75t_R g992 ( 
.A(n_729),
.Y(n_992)
);

INVx1_ASAP7_75t_L g993 ( 
.A(n_622),
.Y(n_993)
);

INVx2_ASAP7_75t_L g994 ( 
.A(n_561),
.Y(n_994)
);

INVx1_ASAP7_75t_L g995 ( 
.A(n_575),
.Y(n_995)
);

INVx1_ASAP7_75t_L g996 ( 
.A(n_714),
.Y(n_996)
);

INVx1_ASAP7_75t_L g997 ( 
.A(n_397),
.Y(n_997)
);

INVx1_ASAP7_75t_L g998 ( 
.A(n_399),
.Y(n_998)
);

INVx1_ASAP7_75t_L g999 ( 
.A(n_400),
.Y(n_999)
);

CKINVDCx16_ASAP7_75t_R g1000 ( 
.A(n_717),
.Y(n_1000)
);

INVx1_ASAP7_75t_L g1001 ( 
.A(n_401),
.Y(n_1001)
);

INVx1_ASAP7_75t_L g1002 ( 
.A(n_403),
.Y(n_1002)
);

CKINVDCx20_ASAP7_75t_R g1003 ( 
.A(n_621),
.Y(n_1003)
);

INVx1_ASAP7_75t_L g1004 ( 
.A(n_404),
.Y(n_1004)
);

CKINVDCx5p33_ASAP7_75t_R g1005 ( 
.A(n_408),
.Y(n_1005)
);

INVx1_ASAP7_75t_L g1006 ( 
.A(n_412),
.Y(n_1006)
);

INVxp33_ASAP7_75t_L g1007 ( 
.A(n_633),
.Y(n_1007)
);

INVxp33_ASAP7_75t_SL g1008 ( 
.A(n_415),
.Y(n_1008)
);

BUFx3_ASAP7_75t_L g1009 ( 
.A(n_943),
.Y(n_1009)
);

NAND2xp5_ASAP7_75t_L g1010 ( 
.A(n_829),
.B(n_650),
.Y(n_1010)
);

AND2x4_ASAP7_75t_L g1011 ( 
.A(n_790),
.B(n_466),
.Y(n_1011)
);

INVx1_ASAP7_75t_L g1012 ( 
.A(n_745),
.Y(n_1012)
);

INVx5_ASAP7_75t_L g1013 ( 
.A(n_861),
.Y(n_1013)
);

BUFx3_ASAP7_75t_L g1014 ( 
.A(n_793),
.Y(n_1014)
);

NAND2xp5_ASAP7_75t_L g1015 ( 
.A(n_829),
.B(n_669),
.Y(n_1015)
);

INVx1_ASAP7_75t_L g1016 ( 
.A(n_747),
.Y(n_1016)
);

BUFx6f_ASAP7_75t_L g1017 ( 
.A(n_861),
.Y(n_1017)
);

BUFx8_ASAP7_75t_SL g1018 ( 
.A(n_972),
.Y(n_1018)
);

INVx2_ASAP7_75t_L g1019 ( 
.A(n_951),
.Y(n_1019)
);

INVx2_ASAP7_75t_SL g1020 ( 
.A(n_800),
.Y(n_1020)
);

INVx1_ASAP7_75t_L g1021 ( 
.A(n_748),
.Y(n_1021)
);

BUFx3_ASAP7_75t_L g1022 ( 
.A(n_804),
.Y(n_1022)
);

NAND2xp5_ASAP7_75t_L g1023 ( 
.A(n_850),
.B(n_669),
.Y(n_1023)
);

BUFx6f_ASAP7_75t_L g1024 ( 
.A(n_861),
.Y(n_1024)
);

AND2x4_ASAP7_75t_L g1025 ( 
.A(n_790),
.B(n_589),
.Y(n_1025)
);

INVx1_ASAP7_75t_L g1026 ( 
.A(n_752),
.Y(n_1026)
);

INVx2_ASAP7_75t_L g1027 ( 
.A(n_978),
.Y(n_1027)
);

BUFx8_ASAP7_75t_SL g1028 ( 
.A(n_982),
.Y(n_1028)
);

BUFx2_ASAP7_75t_L g1029 ( 
.A(n_733),
.Y(n_1029)
);

BUFx6f_ASAP7_75t_L g1030 ( 
.A(n_861),
.Y(n_1030)
);

BUFx6f_ASAP7_75t_L g1031 ( 
.A(n_896),
.Y(n_1031)
);

BUFx8_ASAP7_75t_L g1032 ( 
.A(n_945),
.Y(n_1032)
);

BUFx2_ASAP7_75t_L g1033 ( 
.A(n_822),
.Y(n_1033)
);

INVx5_ASAP7_75t_L g1034 ( 
.A(n_896),
.Y(n_1034)
);

NOR2xp33_ASAP7_75t_R g1035 ( 
.A(n_802),
.B(n_416),
.Y(n_1035)
);

INVx6_ASAP7_75t_L g1036 ( 
.A(n_851),
.Y(n_1036)
);

AOI22xp5_ASAP7_75t_L g1037 ( 
.A1(n_750),
.A2(n_633),
.B1(n_698),
.B2(n_691),
.Y(n_1037)
);

BUFx6f_ASAP7_75t_L g1038 ( 
.A(n_896),
.Y(n_1038)
);

INVx2_ASAP7_75t_L g1039 ( 
.A(n_980),
.Y(n_1039)
);

BUFx6f_ASAP7_75t_L g1040 ( 
.A(n_896),
.Y(n_1040)
);

INVx3_ASAP7_75t_L g1041 ( 
.A(n_808),
.Y(n_1041)
);

INVx1_ASAP7_75t_L g1042 ( 
.A(n_753),
.Y(n_1042)
);

BUFx6f_ASAP7_75t_L g1043 ( 
.A(n_915),
.Y(n_1043)
);

INVx2_ASAP7_75t_L g1044 ( 
.A(n_994),
.Y(n_1044)
);

AND2x4_ASAP7_75t_L g1045 ( 
.A(n_761),
.B(n_623),
.Y(n_1045)
);

INVx1_ASAP7_75t_L g1046 ( 
.A(n_754),
.Y(n_1046)
);

HB1xp67_ASAP7_75t_L g1047 ( 
.A(n_827),
.Y(n_1047)
);

NOR2xp33_ASAP7_75t_L g1048 ( 
.A(n_997),
.B(n_998),
.Y(n_1048)
);

AND2x4_ASAP7_75t_L g1049 ( 
.A(n_821),
.B(n_691),
.Y(n_1049)
);

NOR2x1_ASAP7_75t_L g1050 ( 
.A(n_993),
.B(n_614),
.Y(n_1050)
);

BUFx6f_ASAP7_75t_L g1051 ( 
.A(n_915),
.Y(n_1051)
);

INVx1_ASAP7_75t_L g1052 ( 
.A(n_756),
.Y(n_1052)
);

INVx3_ASAP7_75t_L g1053 ( 
.A(n_809),
.Y(n_1053)
);

BUFx8_ASAP7_75t_L g1054 ( 
.A(n_995),
.Y(n_1054)
);

INVx2_ASAP7_75t_L g1055 ( 
.A(n_766),
.Y(n_1055)
);

INVx2_ASAP7_75t_L g1056 ( 
.A(n_776),
.Y(n_1056)
);

OA21x2_ASAP7_75t_L g1057 ( 
.A1(n_944),
.A2(n_420),
.B(n_419),
.Y(n_1057)
);

CKINVDCx5p33_ASAP7_75t_R g1058 ( 
.A(n_736),
.Y(n_1058)
);

BUFx8_ASAP7_75t_SL g1059 ( 
.A(n_989),
.Y(n_1059)
);

BUFx6f_ASAP7_75t_L g1060 ( 
.A(n_915),
.Y(n_1060)
);

INVx5_ASAP7_75t_L g1061 ( 
.A(n_915),
.Y(n_1061)
);

INVx1_ASAP7_75t_L g1062 ( 
.A(n_757),
.Y(n_1062)
);

BUFx3_ASAP7_75t_L g1063 ( 
.A(n_1005),
.Y(n_1063)
);

INVx1_ASAP7_75t_L g1064 ( 
.A(n_788),
.Y(n_1064)
);

INVx1_ASAP7_75t_L g1065 ( 
.A(n_758),
.Y(n_1065)
);

INVx3_ASAP7_75t_L g1066 ( 
.A(n_789),
.Y(n_1066)
);

BUFx6f_ASAP7_75t_L g1067 ( 
.A(n_956),
.Y(n_1067)
);

BUFx3_ASAP7_75t_L g1068 ( 
.A(n_732),
.Y(n_1068)
);

BUFx6f_ASAP7_75t_L g1069 ( 
.A(n_956),
.Y(n_1069)
);

BUFx6f_ASAP7_75t_L g1070 ( 
.A(n_956),
.Y(n_1070)
);

INVx1_ASAP7_75t_L g1071 ( 
.A(n_762),
.Y(n_1071)
);

BUFx3_ASAP7_75t_L g1072 ( 
.A(n_734),
.Y(n_1072)
);

BUFx12f_ASAP7_75t_L g1073 ( 
.A(n_785),
.Y(n_1073)
);

INVx5_ASAP7_75t_L g1074 ( 
.A(n_956),
.Y(n_1074)
);

HB1xp67_ASAP7_75t_L g1075 ( 
.A(n_840),
.Y(n_1075)
);

INVx1_ASAP7_75t_L g1076 ( 
.A(n_850),
.Y(n_1076)
);

INVx5_ASAP7_75t_L g1077 ( 
.A(n_898),
.Y(n_1077)
);

BUFx6f_ASAP7_75t_L g1078 ( 
.A(n_871),
.Y(n_1078)
);

AOI22xp5_ASAP7_75t_L g1079 ( 
.A1(n_759),
.A2(n_698),
.B1(n_425),
.B2(n_428),
.Y(n_1079)
);

INVx5_ASAP7_75t_L g1080 ( 
.A(n_898),
.Y(n_1080)
);

OAI21x1_ASAP7_75t_L g1081 ( 
.A1(n_853),
.A2(n_666),
.B(n_614),
.Y(n_1081)
);

BUFx6f_ASAP7_75t_L g1082 ( 
.A(n_873),
.Y(n_1082)
);

INVx2_ASAP7_75t_L g1083 ( 
.A(n_760),
.Y(n_1083)
);

CKINVDCx5p33_ASAP7_75t_R g1084 ( 
.A(n_811),
.Y(n_1084)
);

INVx3_ASAP7_75t_L g1085 ( 
.A(n_887),
.Y(n_1085)
);

INVx2_ASAP7_75t_L g1086 ( 
.A(n_760),
.Y(n_1086)
);

BUFx6f_ASAP7_75t_L g1087 ( 
.A(n_889),
.Y(n_1087)
);

AND2x6_ASAP7_75t_L g1088 ( 
.A(n_848),
.B(n_614),
.Y(n_1088)
);

INVx2_ASAP7_75t_L g1089 ( 
.A(n_760),
.Y(n_1089)
);

INVx2_ASAP7_75t_L g1090 ( 
.A(n_760),
.Y(n_1090)
);

BUFx6f_ASAP7_75t_L g1091 ( 
.A(n_907),
.Y(n_1091)
);

INVx2_ASAP7_75t_L g1092 ( 
.A(n_760),
.Y(n_1092)
);

INVx3_ASAP7_75t_L g1093 ( 
.A(n_937),
.Y(n_1093)
);

INVx2_ASAP7_75t_L g1094 ( 
.A(n_760),
.Y(n_1094)
);

NAND2xp5_ASAP7_75t_SL g1095 ( 
.A(n_743),
.B(n_421),
.Y(n_1095)
);

AOI22xp5_ASAP7_75t_L g1096 ( 
.A1(n_759),
.A2(n_436),
.B1(n_438),
.B2(n_431),
.Y(n_1096)
);

NOR2xp33_ASAP7_75t_L g1097 ( 
.A(n_999),
.B(n_442),
.Y(n_1097)
);

INVx2_ASAP7_75t_L g1098 ( 
.A(n_735),
.Y(n_1098)
);

CKINVDCx20_ASAP7_75t_R g1099 ( 
.A(n_769),
.Y(n_1099)
);

NAND2xp5_ASAP7_75t_L g1100 ( 
.A(n_853),
.B(n_444),
.Y(n_1100)
);

HB1xp67_ASAP7_75t_L g1101 ( 
.A(n_854),
.Y(n_1101)
);

BUFx3_ASAP7_75t_L g1102 ( 
.A(n_737),
.Y(n_1102)
);

CKINVDCx20_ASAP7_75t_R g1103 ( 
.A(n_791),
.Y(n_1103)
);

INVx2_ASAP7_75t_L g1104 ( 
.A(n_738),
.Y(n_1104)
);

AND2x2_ASAP7_75t_L g1105 ( 
.A(n_867),
.B(n_445),
.Y(n_1105)
);

OAI22xp5_ASAP7_75t_SL g1106 ( 
.A1(n_838),
.A2(n_453),
.B1(n_455),
.B2(n_449),
.Y(n_1106)
);

BUFx6f_ASAP7_75t_L g1107 ( 
.A(n_940),
.Y(n_1107)
);

AND2x4_ASAP7_75t_L g1108 ( 
.A(n_823),
.B(n_614),
.Y(n_1108)
);

BUFx2_ASAP7_75t_L g1109 ( 
.A(n_860),
.Y(n_1109)
);

BUFx3_ASAP7_75t_L g1110 ( 
.A(n_739),
.Y(n_1110)
);

CKINVDCx6p67_ASAP7_75t_R g1111 ( 
.A(n_764),
.Y(n_1111)
);

INVx2_ASAP7_75t_L g1112 ( 
.A(n_740),
.Y(n_1112)
);

HB1xp67_ASAP7_75t_L g1113 ( 
.A(n_862),
.Y(n_1113)
);

AND2x6_ASAP7_75t_L g1114 ( 
.A(n_849),
.B(n_666),
.Y(n_1114)
);

CKINVDCx14_ASAP7_75t_R g1115 ( 
.A(n_802),
.Y(n_1115)
);

INVx2_ASAP7_75t_L g1116 ( 
.A(n_741),
.Y(n_1116)
);

INVx1_ASAP7_75t_L g1117 ( 
.A(n_763),
.Y(n_1117)
);

INVx1_ASAP7_75t_L g1118 ( 
.A(n_881),
.Y(n_1118)
);

INVx1_ASAP7_75t_L g1119 ( 
.A(n_765),
.Y(n_1119)
);

CKINVDCx20_ASAP7_75t_R g1120 ( 
.A(n_828),
.Y(n_1120)
);

BUFx6f_ASAP7_75t_L g1121 ( 
.A(n_868),
.Y(n_1121)
);

INVx3_ASAP7_75t_L g1122 ( 
.A(n_893),
.Y(n_1122)
);

BUFx6f_ASAP7_75t_L g1123 ( 
.A(n_767),
.Y(n_1123)
);

INVx4_ASAP7_75t_L g1124 ( 
.A(n_875),
.Y(n_1124)
);

OAI21x1_ASAP7_75t_L g1125 ( 
.A1(n_881),
.A2(n_666),
.B(n_461),
.Y(n_1125)
);

AND2x4_ASAP7_75t_L g1126 ( 
.A(n_824),
.B(n_666),
.Y(n_1126)
);

CKINVDCx20_ASAP7_75t_R g1127 ( 
.A(n_831),
.Y(n_1127)
);

NAND2xp5_ASAP7_75t_L g1128 ( 
.A(n_1001),
.B(n_460),
.Y(n_1128)
);

BUFx6f_ASAP7_75t_L g1129 ( 
.A(n_770),
.Y(n_1129)
);

INVx1_ASAP7_75t_L g1130 ( 
.A(n_855),
.Y(n_1130)
);

CKINVDCx11_ASAP7_75t_R g1131 ( 
.A(n_1003),
.Y(n_1131)
);

INVx1_ASAP7_75t_L g1132 ( 
.A(n_856),
.Y(n_1132)
);

INVx4_ASAP7_75t_L g1133 ( 
.A(n_878),
.Y(n_1133)
);

AND2x4_ASAP7_75t_L g1134 ( 
.A(n_825),
.B(n_467),
.Y(n_1134)
);

AND2x4_ASAP7_75t_L g1135 ( 
.A(n_826),
.B(n_470),
.Y(n_1135)
);

NAND2xp5_ASAP7_75t_L g1136 ( 
.A(n_1002),
.B(n_474),
.Y(n_1136)
);

BUFx6f_ASAP7_75t_L g1137 ( 
.A(n_772),
.Y(n_1137)
);

INVx1_ASAP7_75t_L g1138 ( 
.A(n_859),
.Y(n_1138)
);

INVx5_ASAP7_75t_L g1139 ( 
.A(n_851),
.Y(n_1139)
);

INVx2_ASAP7_75t_L g1140 ( 
.A(n_742),
.Y(n_1140)
);

INVx3_ASAP7_75t_L g1141 ( 
.A(n_949),
.Y(n_1141)
);

INVx1_ASAP7_75t_L g1142 ( 
.A(n_863),
.Y(n_1142)
);

BUFx8_ASAP7_75t_SL g1143 ( 
.A(n_852),
.Y(n_1143)
);

BUFx6f_ASAP7_75t_L g1144 ( 
.A(n_773),
.Y(n_1144)
);

AND2x2_ASAP7_75t_L g1145 ( 
.A(n_895),
.B(n_476),
.Y(n_1145)
);

INVx5_ASAP7_75t_L g1146 ( 
.A(n_832),
.Y(n_1146)
);

AND2x2_ASAP7_75t_L g1147 ( 
.A(n_924),
.B(n_477),
.Y(n_1147)
);

INVx2_ASAP7_75t_L g1148 ( 
.A(n_744),
.Y(n_1148)
);

BUFx8_ASAP7_75t_L g1149 ( 
.A(n_996),
.Y(n_1149)
);

AND2x2_ASAP7_75t_L g1150 ( 
.A(n_777),
.B(n_478),
.Y(n_1150)
);

INVx3_ASAP7_75t_L g1151 ( 
.A(n_864),
.Y(n_1151)
);

INVx3_ASAP7_75t_L g1152 ( 
.A(n_865),
.Y(n_1152)
);

AND2x2_ASAP7_75t_L g1153 ( 
.A(n_777),
.B(n_480),
.Y(n_1153)
);

INVx1_ASAP7_75t_L g1154 ( 
.A(n_775),
.Y(n_1154)
);

NAND2xp5_ASAP7_75t_L g1155 ( 
.A(n_1004),
.B(n_484),
.Y(n_1155)
);

AND2x2_ASAP7_75t_L g1156 ( 
.A(n_858),
.B(n_485),
.Y(n_1156)
);

INVx5_ASAP7_75t_L g1157 ( 
.A(n_774),
.Y(n_1157)
);

AND2x4_ASAP7_75t_L g1158 ( 
.A(n_830),
.B(n_487),
.Y(n_1158)
);

INVx2_ASAP7_75t_L g1159 ( 
.A(n_780),
.Y(n_1159)
);

BUFx12f_ASAP7_75t_L g1160 ( 
.A(n_818),
.Y(n_1160)
);

CKINVDCx5p33_ASAP7_75t_R g1161 ( 
.A(n_857),
.Y(n_1161)
);

INVx1_ASAP7_75t_L g1162 ( 
.A(n_782),
.Y(n_1162)
);

BUFx6f_ASAP7_75t_L g1163 ( 
.A(n_783),
.Y(n_1163)
);

INVx6_ASAP7_75t_L g1164 ( 
.A(n_813),
.Y(n_1164)
);

NAND2xp5_ASAP7_75t_L g1165 ( 
.A(n_1006),
.B(n_954),
.Y(n_1165)
);

NAND2xp5_ASAP7_75t_L g1166 ( 
.A(n_954),
.B(n_490),
.Y(n_1166)
);

AND2x2_ASAP7_75t_L g1167 ( 
.A(n_858),
.B(n_883),
.Y(n_1167)
);

NAND2xp5_ASAP7_75t_L g1168 ( 
.A(n_957),
.B(n_491),
.Y(n_1168)
);

AOI22xp5_ASAP7_75t_L g1169 ( 
.A1(n_836),
.A2(n_497),
.B1(n_504),
.B2(n_494),
.Y(n_1169)
);

CKINVDCx5p33_ASAP7_75t_R g1170 ( 
.A(n_870),
.Y(n_1170)
);

HB1xp67_ASAP7_75t_L g1171 ( 
.A(n_899),
.Y(n_1171)
);

HB1xp67_ASAP7_75t_L g1172 ( 
.A(n_900),
.Y(n_1172)
);

BUFx12f_ASAP7_75t_L g1173 ( 
.A(n_992),
.Y(n_1173)
);

INVx5_ASAP7_75t_L g1174 ( 
.A(n_1000),
.Y(n_1174)
);

INVx1_ASAP7_75t_L g1175 ( 
.A(n_784),
.Y(n_1175)
);

INVx2_ASAP7_75t_L g1176 ( 
.A(n_786),
.Y(n_1176)
);

CKINVDCx5p33_ASAP7_75t_R g1177 ( 
.A(n_885),
.Y(n_1177)
);

BUFx6f_ASAP7_75t_L g1178 ( 
.A(n_794),
.Y(n_1178)
);

INVx1_ASAP7_75t_L g1179 ( 
.A(n_866),
.Y(n_1179)
);

BUFx8_ASAP7_75t_SL g1180 ( 
.A(n_928),
.Y(n_1180)
);

INVx1_ASAP7_75t_L g1181 ( 
.A(n_869),
.Y(n_1181)
);

INVx1_ASAP7_75t_L g1182 ( 
.A(n_872),
.Y(n_1182)
);

INVx1_ASAP7_75t_L g1183 ( 
.A(n_874),
.Y(n_1183)
);

AND2x2_ASAP7_75t_L g1184 ( 
.A(n_883),
.B(n_510),
.Y(n_1184)
);

AOI22x1_ASAP7_75t_SL g1185 ( 
.A1(n_933),
.A2(n_963),
.B1(n_969),
.B2(n_755),
.Y(n_1185)
);

INVx3_ASAP7_75t_L g1186 ( 
.A(n_876),
.Y(n_1186)
);

BUFx3_ASAP7_75t_L g1187 ( 
.A(n_1008),
.Y(n_1187)
);

AND2x4_ASAP7_75t_L g1188 ( 
.A(n_833),
.B(n_517),
.Y(n_1188)
);

CKINVDCx16_ASAP7_75t_R g1189 ( 
.A(n_923),
.Y(n_1189)
);

BUFx8_ASAP7_75t_L g1190 ( 
.A(n_846),
.Y(n_1190)
);

INVx5_ASAP7_75t_L g1191 ( 
.A(n_906),
.Y(n_1191)
);

INVx2_ASAP7_75t_L g1192 ( 
.A(n_796),
.Y(n_1192)
);

AND2x4_ASAP7_75t_L g1193 ( 
.A(n_834),
.B(n_518),
.Y(n_1193)
);

AND2x4_ASAP7_75t_L g1194 ( 
.A(n_1191),
.B(n_1122),
.Y(n_1194)
);

INVx1_ASAP7_75t_L g1195 ( 
.A(n_1014),
.Y(n_1195)
);

NAND2xp5_ASAP7_75t_L g1196 ( 
.A(n_1012),
.B(n_906),
.Y(n_1196)
);

NAND2xp5_ASAP7_75t_SL g1197 ( 
.A(n_1124),
.B(n_795),
.Y(n_1197)
);

AND2x2_ASAP7_75t_L g1198 ( 
.A(n_1167),
.B(n_836),
.Y(n_1198)
);

INVx2_ASAP7_75t_L g1199 ( 
.A(n_1041),
.Y(n_1199)
);

NAND2xp5_ASAP7_75t_SL g1200 ( 
.A(n_1124),
.B(n_805),
.Y(n_1200)
);

AND2x2_ASAP7_75t_L g1201 ( 
.A(n_1191),
.B(n_839),
.Y(n_1201)
);

INVx4_ASAP7_75t_L g1202 ( 
.A(n_1139),
.Y(n_1202)
);

BUFx6f_ASAP7_75t_L g1203 ( 
.A(n_1078),
.Y(n_1203)
);

INVx6_ASAP7_75t_L g1204 ( 
.A(n_1157),
.Y(n_1204)
);

INVx2_ASAP7_75t_L g1205 ( 
.A(n_1041),
.Y(n_1205)
);

HB1xp67_ASAP7_75t_L g1206 ( 
.A(n_1058),
.Y(n_1206)
);

INVx1_ASAP7_75t_L g1207 ( 
.A(n_1022),
.Y(n_1207)
);

INVxp67_ASAP7_75t_L g1208 ( 
.A(n_1029),
.Y(n_1208)
);

AND2x4_ASAP7_75t_L g1209 ( 
.A(n_1191),
.B(n_835),
.Y(n_1209)
);

AND2x4_ASAP7_75t_L g1210 ( 
.A(n_1122),
.B(n_837),
.Y(n_1210)
);

INVx2_ASAP7_75t_L g1211 ( 
.A(n_1053),
.Y(n_1211)
);

NAND2xp5_ASAP7_75t_L g1212 ( 
.A(n_1012),
.B(n_929),
.Y(n_1212)
);

INVx2_ASAP7_75t_L g1213 ( 
.A(n_1053),
.Y(n_1213)
);

INVx1_ASAP7_75t_L g1214 ( 
.A(n_1098),
.Y(n_1214)
);

INVx1_ASAP7_75t_L g1215 ( 
.A(n_1104),
.Y(n_1215)
);

INVx3_ASAP7_75t_L g1216 ( 
.A(n_1078),
.Y(n_1216)
);

NAND2xp5_ASAP7_75t_L g1217 ( 
.A(n_1016),
.B(n_929),
.Y(n_1217)
);

INVx2_ASAP7_75t_L g1218 ( 
.A(n_1078),
.Y(n_1218)
);

CKINVDCx5p33_ASAP7_75t_R g1219 ( 
.A(n_1084),
.Y(n_1219)
);

AND2x2_ASAP7_75t_SL g1220 ( 
.A(n_1033),
.B(n_886),
.Y(n_1220)
);

INVx2_ASAP7_75t_L g1221 ( 
.A(n_1082),
.Y(n_1221)
);

NAND2xp5_ASAP7_75t_L g1222 ( 
.A(n_1016),
.B(n_892),
.Y(n_1222)
);

INVx1_ASAP7_75t_L g1223 ( 
.A(n_1112),
.Y(n_1223)
);

INVx1_ASAP7_75t_L g1224 ( 
.A(n_1116),
.Y(n_1224)
);

BUFx6f_ASAP7_75t_L g1225 ( 
.A(n_1082),
.Y(n_1225)
);

INVx2_ASAP7_75t_L g1226 ( 
.A(n_1082),
.Y(n_1226)
);

BUFx6f_ASAP7_75t_L g1227 ( 
.A(n_1087),
.Y(n_1227)
);

INVx3_ASAP7_75t_L g1228 ( 
.A(n_1087),
.Y(n_1228)
);

AND2x4_ASAP7_75t_L g1229 ( 
.A(n_1011),
.B(n_1025),
.Y(n_1229)
);

AND2x2_ASAP7_75t_L g1230 ( 
.A(n_1045),
.B(n_839),
.Y(n_1230)
);

OA21x2_ASAP7_75t_L g1231 ( 
.A1(n_1081),
.A2(n_1125),
.B(n_1086),
.Y(n_1231)
);

INVx2_ASAP7_75t_L g1232 ( 
.A(n_1087),
.Y(n_1232)
);

AND2x2_ASAP7_75t_SL g1233 ( 
.A(n_1109),
.B(n_886),
.Y(n_1233)
);

AND2x2_ASAP7_75t_L g1234 ( 
.A(n_1045),
.B(n_971),
.Y(n_1234)
);

INVx1_ASAP7_75t_L g1235 ( 
.A(n_1140),
.Y(n_1235)
);

BUFx6f_ASAP7_75t_L g1236 ( 
.A(n_1091),
.Y(n_1236)
);

INVx1_ASAP7_75t_L g1237 ( 
.A(n_1148),
.Y(n_1237)
);

INVx2_ASAP7_75t_L g1238 ( 
.A(n_1091),
.Y(n_1238)
);

INVx1_ASAP7_75t_L g1239 ( 
.A(n_1159),
.Y(n_1239)
);

BUFx6f_ASAP7_75t_L g1240 ( 
.A(n_1091),
.Y(n_1240)
);

NAND2xp5_ASAP7_75t_L g1241 ( 
.A(n_1021),
.B(n_892),
.Y(n_1241)
);

INVx1_ASAP7_75t_L g1242 ( 
.A(n_1176),
.Y(n_1242)
);

INVx1_ASAP7_75t_L g1243 ( 
.A(n_1192),
.Y(n_1243)
);

BUFx6f_ASAP7_75t_L g1244 ( 
.A(n_1107),
.Y(n_1244)
);

BUFx6f_ASAP7_75t_L g1245 ( 
.A(n_1107),
.Y(n_1245)
);

INVx1_ASAP7_75t_L g1246 ( 
.A(n_1130),
.Y(n_1246)
);

INVx3_ASAP7_75t_L g1247 ( 
.A(n_1107),
.Y(n_1247)
);

INVx1_ASAP7_75t_L g1248 ( 
.A(n_1130),
.Y(n_1248)
);

INVx2_ASAP7_75t_L g1249 ( 
.A(n_1019),
.Y(n_1249)
);

BUFx2_ASAP7_75t_L g1250 ( 
.A(n_1173),
.Y(n_1250)
);

BUFx2_ASAP7_75t_L g1251 ( 
.A(n_1164),
.Y(n_1251)
);

INVx2_ASAP7_75t_L g1252 ( 
.A(n_1027),
.Y(n_1252)
);

AND2x2_ASAP7_75t_L g1253 ( 
.A(n_1105),
.B(n_971),
.Y(n_1253)
);

INVx1_ASAP7_75t_L g1254 ( 
.A(n_1132),
.Y(n_1254)
);

NAND2xp5_ASAP7_75t_L g1255 ( 
.A(n_1021),
.B(n_1052),
.Y(n_1255)
);

BUFx6f_ASAP7_75t_L g1256 ( 
.A(n_1017),
.Y(n_1256)
);

OAI22xp5_ASAP7_75t_SL g1257 ( 
.A1(n_1037),
.A2(n_1007),
.B1(n_979),
.B2(n_1099),
.Y(n_1257)
);

HB1xp67_ASAP7_75t_L g1258 ( 
.A(n_1145),
.Y(n_1258)
);

NOR2x1_ASAP7_75t_L g1259 ( 
.A(n_1010),
.B(n_877),
.Y(n_1259)
);

INVx2_ASAP7_75t_L g1260 ( 
.A(n_1039),
.Y(n_1260)
);

INVx1_ASAP7_75t_L g1261 ( 
.A(n_1132),
.Y(n_1261)
);

NAND2xp5_ASAP7_75t_L g1262 ( 
.A(n_1052),
.B(n_908),
.Y(n_1262)
);

HB1xp67_ASAP7_75t_L g1263 ( 
.A(n_1147),
.Y(n_1263)
);

AND2x4_ASAP7_75t_L g1264 ( 
.A(n_1011),
.B(n_1025),
.Y(n_1264)
);

INVx2_ASAP7_75t_L g1265 ( 
.A(n_1044),
.Y(n_1265)
);

CKINVDCx11_ASAP7_75t_R g1266 ( 
.A(n_1131),
.Y(n_1266)
);

INVx2_ASAP7_75t_L g1267 ( 
.A(n_1055),
.Y(n_1267)
);

NOR2xp33_ASAP7_75t_L g1268 ( 
.A(n_1128),
.B(n_880),
.Y(n_1268)
);

INVx2_ASAP7_75t_L g1269 ( 
.A(n_1056),
.Y(n_1269)
);

AND2x4_ASAP7_75t_L g1270 ( 
.A(n_1108),
.B(n_841),
.Y(n_1270)
);

NAND2xp5_ASAP7_75t_L g1271 ( 
.A(n_1026),
.B(n_1042),
.Y(n_1271)
);

AND2x2_ASAP7_75t_L g1272 ( 
.A(n_1150),
.B(n_977),
.Y(n_1272)
);

AND2x2_ASAP7_75t_L g1273 ( 
.A(n_1153),
.B(n_977),
.Y(n_1273)
);

INVx1_ASAP7_75t_L g1274 ( 
.A(n_1138),
.Y(n_1274)
);

BUFx8_ASAP7_75t_L g1275 ( 
.A(n_1073),
.Y(n_1275)
);

AND2x2_ASAP7_75t_L g1276 ( 
.A(n_1036),
.B(n_987),
.Y(n_1276)
);

BUFx8_ASAP7_75t_L g1277 ( 
.A(n_1160),
.Y(n_1277)
);

NOR2xp33_ASAP7_75t_L g1278 ( 
.A(n_1136),
.B(n_905),
.Y(n_1278)
);

INVx5_ASAP7_75t_L g1279 ( 
.A(n_1088),
.Y(n_1279)
);

AND2x4_ASAP7_75t_L g1280 ( 
.A(n_1108),
.B(n_843),
.Y(n_1280)
);

NAND2xp5_ASAP7_75t_SL g1281 ( 
.A(n_1133),
.B(n_911),
.Y(n_1281)
);

INVx2_ASAP7_75t_L g1282 ( 
.A(n_1066),
.Y(n_1282)
);

AND2x2_ASAP7_75t_L g1283 ( 
.A(n_1036),
.B(n_1115),
.Y(n_1283)
);

BUFx3_ASAP7_75t_L g1284 ( 
.A(n_1121),
.Y(n_1284)
);

NAND2xp5_ASAP7_75t_SL g1285 ( 
.A(n_1133),
.B(n_959),
.Y(n_1285)
);

INVx1_ASAP7_75t_L g1286 ( 
.A(n_1138),
.Y(n_1286)
);

NAND2xp5_ASAP7_75t_L g1287 ( 
.A(n_1046),
.B(n_1076),
.Y(n_1287)
);

INVx1_ASAP7_75t_L g1288 ( 
.A(n_1142),
.Y(n_1288)
);

INVxp67_ASAP7_75t_L g1289 ( 
.A(n_1156),
.Y(n_1289)
);

INVx2_ASAP7_75t_L g1290 ( 
.A(n_1066),
.Y(n_1290)
);

INVx1_ASAP7_75t_L g1291 ( 
.A(n_1142),
.Y(n_1291)
);

AND2x4_ASAP7_75t_L g1292 ( 
.A(n_1126),
.B(n_844),
.Y(n_1292)
);

INVx1_ASAP7_75t_L g1293 ( 
.A(n_1179),
.Y(n_1293)
);

XNOR2xp5_ASAP7_75t_L g1294 ( 
.A(n_1103),
.B(n_845),
.Y(n_1294)
);

OA21x2_ASAP7_75t_L g1295 ( 
.A1(n_1083),
.A2(n_882),
.B(n_879),
.Y(n_1295)
);

NAND2xp33_ASAP7_75t_SL g1296 ( 
.A(n_1035),
.B(n_799),
.Y(n_1296)
);

CKINVDCx8_ASAP7_75t_R g1297 ( 
.A(n_1189),
.Y(n_1297)
);

INVx3_ASAP7_75t_L g1298 ( 
.A(n_1151),
.Y(n_1298)
);

INVx1_ASAP7_75t_L g1299 ( 
.A(n_1179),
.Y(n_1299)
);

AND2x2_ASAP7_75t_L g1300 ( 
.A(n_1184),
.B(n_1020),
.Y(n_1300)
);

NAND2xp5_ASAP7_75t_L g1301 ( 
.A(n_1076),
.B(n_908),
.Y(n_1301)
);

INVx1_ASAP7_75t_L g1302 ( 
.A(n_1181),
.Y(n_1302)
);

HB1xp67_ASAP7_75t_L g1303 ( 
.A(n_1164),
.Y(n_1303)
);

INVx3_ASAP7_75t_L g1304 ( 
.A(n_1151),
.Y(n_1304)
);

NAND2xp5_ASAP7_75t_L g1305 ( 
.A(n_1118),
.B(n_919),
.Y(n_1305)
);

NAND2xp5_ASAP7_75t_L g1306 ( 
.A(n_1118),
.B(n_919),
.Y(n_1306)
);

AND2x2_ASAP7_75t_L g1307 ( 
.A(n_1187),
.B(n_987),
.Y(n_1307)
);

INVx1_ASAP7_75t_L g1308 ( 
.A(n_1181),
.Y(n_1308)
);

INVx1_ASAP7_75t_L g1309 ( 
.A(n_1182),
.Y(n_1309)
);

INVx1_ASAP7_75t_L g1310 ( 
.A(n_1182),
.Y(n_1310)
);

NAND2xp5_ASAP7_75t_L g1311 ( 
.A(n_1089),
.B(n_1090),
.Y(n_1311)
);

NAND2xp5_ASAP7_75t_SL g1312 ( 
.A(n_1139),
.B(n_946),
.Y(n_1312)
);

INVx1_ASAP7_75t_L g1313 ( 
.A(n_1183),
.Y(n_1313)
);

INVx2_ASAP7_75t_L g1314 ( 
.A(n_1085),
.Y(n_1314)
);

NAND2xp5_ASAP7_75t_L g1315 ( 
.A(n_1092),
.B(n_922),
.Y(n_1315)
);

INVx1_ASAP7_75t_L g1316 ( 
.A(n_1183),
.Y(n_1316)
);

BUFx6f_ASAP7_75t_L g1317 ( 
.A(n_1024),
.Y(n_1317)
);

AND2x4_ASAP7_75t_L g1318 ( 
.A(n_1126),
.B(n_847),
.Y(n_1318)
);

INVx1_ASAP7_75t_L g1319 ( 
.A(n_1062),
.Y(n_1319)
);

AND2x2_ASAP7_75t_L g1320 ( 
.A(n_1157),
.B(n_957),
.Y(n_1320)
);

INVx1_ASAP7_75t_L g1321 ( 
.A(n_1065),
.Y(n_1321)
);

BUFx2_ASAP7_75t_L g1322 ( 
.A(n_1018),
.Y(n_1322)
);

INVx1_ASAP7_75t_L g1323 ( 
.A(n_1071),
.Y(n_1323)
);

OA21x2_ASAP7_75t_L g1324 ( 
.A1(n_1094),
.A2(n_888),
.B(n_884),
.Y(n_1324)
);

BUFx2_ASAP7_75t_L g1325 ( 
.A(n_1028),
.Y(n_1325)
);

BUFx6f_ASAP7_75t_L g1326 ( 
.A(n_1024),
.Y(n_1326)
);

CKINVDCx5p33_ASAP7_75t_R g1327 ( 
.A(n_1059),
.Y(n_1327)
);

OAI22xp5_ASAP7_75t_SL g1328 ( 
.A1(n_1120),
.A2(n_819),
.B1(n_817),
.B2(n_781),
.Y(n_1328)
);

INVx1_ASAP7_75t_L g1329 ( 
.A(n_1117),
.Y(n_1329)
);

INVx1_ASAP7_75t_L g1330 ( 
.A(n_1119),
.Y(n_1330)
);

CKINVDCx8_ASAP7_75t_R g1331 ( 
.A(n_1161),
.Y(n_1331)
);

INVx1_ASAP7_75t_L g1332 ( 
.A(n_1154),
.Y(n_1332)
);

INVx1_ASAP7_75t_L g1333 ( 
.A(n_1162),
.Y(n_1333)
);

AND2x2_ASAP7_75t_L g1334 ( 
.A(n_1157),
.B(n_984),
.Y(n_1334)
);

NOR2xp33_ASAP7_75t_L g1335 ( 
.A(n_1155),
.B(n_1100),
.Y(n_1335)
);

INVx1_ASAP7_75t_L g1336 ( 
.A(n_1175),
.Y(n_1336)
);

BUFx6f_ASAP7_75t_L g1337 ( 
.A(n_1030),
.Y(n_1337)
);

INVx1_ASAP7_75t_L g1338 ( 
.A(n_1123),
.Y(n_1338)
);

NAND2xp5_ASAP7_75t_L g1339 ( 
.A(n_1015),
.B(n_922),
.Y(n_1339)
);

BUFx6f_ASAP7_75t_L g1340 ( 
.A(n_1030),
.Y(n_1340)
);

AND2x2_ASAP7_75t_L g1341 ( 
.A(n_1174),
.B(n_984),
.Y(n_1341)
);

CKINVDCx5p33_ASAP7_75t_R g1342 ( 
.A(n_1143),
.Y(n_1342)
);

NAND2xp33_ASAP7_75t_L g1343 ( 
.A(n_1139),
.B(n_947),
.Y(n_1343)
);

INVxp67_ASAP7_75t_L g1344 ( 
.A(n_1023),
.Y(n_1344)
);

CKINVDCx5p33_ASAP7_75t_R g1345 ( 
.A(n_1180),
.Y(n_1345)
);

INVx2_ASAP7_75t_L g1346 ( 
.A(n_1085),
.Y(n_1346)
);

AND2x2_ASAP7_75t_L g1347 ( 
.A(n_1174),
.B(n_779),
.Y(n_1347)
);

INVx2_ASAP7_75t_L g1348 ( 
.A(n_1093),
.Y(n_1348)
);

INVxp67_ASAP7_75t_L g1349 ( 
.A(n_1166),
.Y(n_1349)
);

BUFx8_ASAP7_75t_L g1350 ( 
.A(n_1063),
.Y(n_1350)
);

OAI22xp33_ASAP7_75t_L g1351 ( 
.A1(n_1339),
.A2(n_1079),
.B1(n_799),
.B2(n_1165),
.Y(n_1351)
);

INVx1_ASAP7_75t_L g1352 ( 
.A(n_1246),
.Y(n_1352)
);

INVx2_ASAP7_75t_L g1353 ( 
.A(n_1199),
.Y(n_1353)
);

INVx2_ASAP7_75t_L g1354 ( 
.A(n_1205),
.Y(n_1354)
);

INVxp67_ASAP7_75t_SL g1355 ( 
.A(n_1229),
.Y(n_1355)
);

NAND2xp5_ASAP7_75t_SL g1356 ( 
.A(n_1272),
.B(n_1047),
.Y(n_1356)
);

INVx2_ASAP7_75t_SL g1357 ( 
.A(n_1229),
.Y(n_1357)
);

INVx1_ASAP7_75t_L g1358 ( 
.A(n_1248),
.Y(n_1358)
);

INVx2_ASAP7_75t_SL g1359 ( 
.A(n_1264),
.Y(n_1359)
);

INVx1_ASAP7_75t_SL g1360 ( 
.A(n_1264),
.Y(n_1360)
);

INVx2_ASAP7_75t_L g1361 ( 
.A(n_1211),
.Y(n_1361)
);

INVx2_ASAP7_75t_L g1362 ( 
.A(n_1213),
.Y(n_1362)
);

INVx1_ASAP7_75t_L g1363 ( 
.A(n_1254),
.Y(n_1363)
);

AND2x6_ASAP7_75t_L g1364 ( 
.A(n_1283),
.B(n_1193),
.Y(n_1364)
);

INVx3_ASAP7_75t_L g1365 ( 
.A(n_1203),
.Y(n_1365)
);

INVx1_ASAP7_75t_L g1366 ( 
.A(n_1261),
.Y(n_1366)
);

INVx1_ASAP7_75t_L g1367 ( 
.A(n_1274),
.Y(n_1367)
);

NAND2xp5_ASAP7_75t_SL g1368 ( 
.A(n_1273),
.B(n_1075),
.Y(n_1368)
);

BUFx2_ASAP7_75t_L g1369 ( 
.A(n_1251),
.Y(n_1369)
);

INVx2_ASAP7_75t_L g1370 ( 
.A(n_1314),
.Y(n_1370)
);

NAND2xp5_ASAP7_75t_SL g1371 ( 
.A(n_1320),
.B(n_1101),
.Y(n_1371)
);

INVx2_ASAP7_75t_L g1372 ( 
.A(n_1346),
.Y(n_1372)
);

INVx1_ASAP7_75t_L g1373 ( 
.A(n_1286),
.Y(n_1373)
);

CKINVDCx5p33_ASAP7_75t_R g1374 ( 
.A(n_1219),
.Y(n_1374)
);

INVx2_ASAP7_75t_L g1375 ( 
.A(n_1348),
.Y(n_1375)
);

INVx1_ASAP7_75t_L g1376 ( 
.A(n_1288),
.Y(n_1376)
);

NOR3xp33_ASAP7_75t_L g1377 ( 
.A(n_1198),
.B(n_1106),
.C(n_1168),
.Y(n_1377)
);

INVx2_ASAP7_75t_L g1378 ( 
.A(n_1282),
.Y(n_1378)
);

INVx4_ASAP7_75t_L g1379 ( 
.A(n_1204),
.Y(n_1379)
);

INVx2_ASAP7_75t_L g1380 ( 
.A(n_1290),
.Y(n_1380)
);

INVx2_ASAP7_75t_L g1381 ( 
.A(n_1249),
.Y(n_1381)
);

BUFx6f_ASAP7_75t_L g1382 ( 
.A(n_1203),
.Y(n_1382)
);

AND2x2_ASAP7_75t_L g1383 ( 
.A(n_1230),
.B(n_1113),
.Y(n_1383)
);

NOR2x1p5_ASAP7_75t_L g1384 ( 
.A(n_1327),
.B(n_1111),
.Y(n_1384)
);

INVx1_ASAP7_75t_L g1385 ( 
.A(n_1291),
.Y(n_1385)
);

NAND2xp5_ASAP7_75t_L g1386 ( 
.A(n_1335),
.B(n_1048),
.Y(n_1386)
);

INVx3_ASAP7_75t_L g1387 ( 
.A(n_1203),
.Y(n_1387)
);

AND2x6_ASAP7_75t_L g1388 ( 
.A(n_1234),
.B(n_1259),
.Y(n_1388)
);

NAND3xp33_ASAP7_75t_L g1389 ( 
.A(n_1344),
.B(n_1097),
.C(n_1152),
.Y(n_1389)
);

INVx1_ASAP7_75t_L g1390 ( 
.A(n_1293),
.Y(n_1390)
);

INVx2_ASAP7_75t_L g1391 ( 
.A(n_1252),
.Y(n_1391)
);

CKINVDCx5p33_ASAP7_75t_R g1392 ( 
.A(n_1342),
.Y(n_1392)
);

INVx3_ASAP7_75t_L g1393 ( 
.A(n_1225),
.Y(n_1393)
);

NAND2xp5_ASAP7_75t_L g1394 ( 
.A(n_1344),
.B(n_1152),
.Y(n_1394)
);

OAI22xp5_ASAP7_75t_L g1395 ( 
.A1(n_1289),
.A2(n_890),
.B1(n_842),
.B2(n_1096),
.Y(n_1395)
);

INVx2_ASAP7_75t_L g1396 ( 
.A(n_1260),
.Y(n_1396)
);

INVx1_ASAP7_75t_L g1397 ( 
.A(n_1299),
.Y(n_1397)
);

INVx2_ASAP7_75t_L g1398 ( 
.A(n_1265),
.Y(n_1398)
);

INVxp67_ASAP7_75t_L g1399 ( 
.A(n_1307),
.Y(n_1399)
);

INVx2_ASAP7_75t_L g1400 ( 
.A(n_1267),
.Y(n_1400)
);

INVx2_ASAP7_75t_SL g1401 ( 
.A(n_1276),
.Y(n_1401)
);

INVx4_ASAP7_75t_L g1402 ( 
.A(n_1204),
.Y(n_1402)
);

NOR2xp33_ASAP7_75t_L g1403 ( 
.A(n_1349),
.B(n_1171),
.Y(n_1403)
);

INVx2_ASAP7_75t_L g1404 ( 
.A(n_1269),
.Y(n_1404)
);

NAND2xp5_ASAP7_75t_L g1405 ( 
.A(n_1339),
.B(n_1186),
.Y(n_1405)
);

NOR2xp33_ASAP7_75t_L g1406 ( 
.A(n_1349),
.B(n_1172),
.Y(n_1406)
);

INVxp67_ASAP7_75t_SL g1407 ( 
.A(n_1301),
.Y(n_1407)
);

INVx2_ASAP7_75t_L g1408 ( 
.A(n_1214),
.Y(n_1408)
);

INVx1_ASAP7_75t_L g1409 ( 
.A(n_1302),
.Y(n_1409)
);

NAND2xp33_ASAP7_75t_SL g1410 ( 
.A(n_1253),
.B(n_1206),
.Y(n_1410)
);

INVx1_ASAP7_75t_L g1411 ( 
.A(n_1308),
.Y(n_1411)
);

AND3x2_ASAP7_75t_L g1412 ( 
.A(n_1250),
.B(n_1049),
.C(n_771),
.Y(n_1412)
);

BUFx2_ASAP7_75t_L g1413 ( 
.A(n_1208),
.Y(n_1413)
);

BUFx3_ASAP7_75t_L g1414 ( 
.A(n_1350),
.Y(n_1414)
);

INVx2_ASAP7_75t_L g1415 ( 
.A(n_1215),
.Y(n_1415)
);

INVx3_ASAP7_75t_L g1416 ( 
.A(n_1225),
.Y(n_1416)
);

INVx2_ASAP7_75t_L g1417 ( 
.A(n_1223),
.Y(n_1417)
);

AND2x6_ASAP7_75t_L g1418 ( 
.A(n_1259),
.B(n_1193),
.Y(n_1418)
);

INVx1_ASAP7_75t_L g1419 ( 
.A(n_1309),
.Y(n_1419)
);

BUFx2_ASAP7_75t_L g1420 ( 
.A(n_1303),
.Y(n_1420)
);

INVx2_ASAP7_75t_L g1421 ( 
.A(n_1224),
.Y(n_1421)
);

NAND2xp5_ASAP7_75t_SL g1422 ( 
.A(n_1334),
.B(n_1134),
.Y(n_1422)
);

NAND2xp5_ASAP7_75t_L g1423 ( 
.A(n_1287),
.B(n_1186),
.Y(n_1423)
);

INVx2_ASAP7_75t_L g1424 ( 
.A(n_1235),
.Y(n_1424)
);

INVx2_ASAP7_75t_L g1425 ( 
.A(n_1237),
.Y(n_1425)
);

NAND2xp5_ASAP7_75t_L g1426 ( 
.A(n_1287),
.B(n_1134),
.Y(n_1426)
);

NAND2xp5_ASAP7_75t_L g1427 ( 
.A(n_1255),
.B(n_1135),
.Y(n_1427)
);

AOI22x1_ASAP7_75t_L g1428 ( 
.A1(n_1310),
.A2(n_1158),
.B1(n_1188),
.B2(n_1135),
.Y(n_1428)
);

INVx2_ASAP7_75t_SL g1429 ( 
.A(n_1347),
.Y(n_1429)
);

NAND3xp33_ASAP7_75t_L g1430 ( 
.A(n_1289),
.B(n_1080),
.C(n_1077),
.Y(n_1430)
);

INVx1_ASAP7_75t_L g1431 ( 
.A(n_1313),
.Y(n_1431)
);

BUFx3_ASAP7_75t_L g1432 ( 
.A(n_1350),
.Y(n_1432)
);

NAND2xp5_ASAP7_75t_SL g1433 ( 
.A(n_1341),
.B(n_1158),
.Y(n_1433)
);

INVx3_ASAP7_75t_L g1434 ( 
.A(n_1225),
.Y(n_1434)
);

OAI22xp33_ASAP7_75t_L g1435 ( 
.A1(n_1258),
.A2(n_1169),
.B1(n_1174),
.B2(n_1146),
.Y(n_1435)
);

AOI22xp33_ASAP7_75t_SL g1436 ( 
.A1(n_1220),
.A2(n_1049),
.B1(n_1185),
.B2(n_934),
.Y(n_1436)
);

AND2x4_ASAP7_75t_L g1437 ( 
.A(n_1194),
.B(n_1009),
.Y(n_1437)
);

BUFx3_ASAP7_75t_L g1438 ( 
.A(n_1297),
.Y(n_1438)
);

INVx1_ASAP7_75t_L g1439 ( 
.A(n_1316),
.Y(n_1439)
);

NOR2x1p5_ASAP7_75t_L g1440 ( 
.A(n_1345),
.B(n_1188),
.Y(n_1440)
);

INVx3_ASAP7_75t_L g1441 ( 
.A(n_1227),
.Y(n_1441)
);

INVx6_ASAP7_75t_L g1442 ( 
.A(n_1275),
.Y(n_1442)
);

AOI22xp33_ASAP7_75t_L g1443 ( 
.A1(n_1328),
.A2(n_1057),
.B1(n_934),
.B2(n_927),
.Y(n_1443)
);

NAND2xp5_ASAP7_75t_L g1444 ( 
.A(n_1255),
.B(n_1057),
.Y(n_1444)
);

INVx2_ASAP7_75t_SL g1445 ( 
.A(n_1300),
.Y(n_1445)
);

BUFx3_ASAP7_75t_L g1446 ( 
.A(n_1331),
.Y(n_1446)
);

INVx4_ASAP7_75t_L g1447 ( 
.A(n_1194),
.Y(n_1447)
);

INVx1_ASAP7_75t_L g1448 ( 
.A(n_1319),
.Y(n_1448)
);

INVx1_ASAP7_75t_L g1449 ( 
.A(n_1321),
.Y(n_1449)
);

INVx2_ASAP7_75t_L g1450 ( 
.A(n_1239),
.Y(n_1450)
);

INVx8_ASAP7_75t_L g1451 ( 
.A(n_1210),
.Y(n_1451)
);

AOI22xp33_ASAP7_75t_L g1452 ( 
.A1(n_1328),
.A2(n_927),
.B1(n_1129),
.B2(n_1123),
.Y(n_1452)
);

OR2x2_ASAP7_75t_L g1453 ( 
.A(n_1257),
.B(n_1170),
.Y(n_1453)
);

INVx1_ASAP7_75t_L g1454 ( 
.A(n_1323),
.Y(n_1454)
);

AND2x2_ASAP7_75t_L g1455 ( 
.A(n_1233),
.B(n_1121),
.Y(n_1455)
);

INVx2_ASAP7_75t_L g1456 ( 
.A(n_1242),
.Y(n_1456)
);

NOR3xp33_ASAP7_75t_L g1457 ( 
.A(n_1296),
.B(n_1095),
.C(n_950),
.Y(n_1457)
);

NAND2xp5_ASAP7_75t_SL g1458 ( 
.A(n_1268),
.B(n_1077),
.Y(n_1458)
);

INVx2_ASAP7_75t_L g1459 ( 
.A(n_1243),
.Y(n_1459)
);

NAND3xp33_ASAP7_75t_L g1460 ( 
.A(n_1271),
.B(n_1080),
.C(n_1077),
.Y(n_1460)
);

BUFx6f_ASAP7_75t_L g1461 ( 
.A(n_1227),
.Y(n_1461)
);

NOR2xp33_ASAP7_75t_L g1462 ( 
.A(n_1278),
.B(n_1146),
.Y(n_1462)
);

INVx1_ASAP7_75t_L g1463 ( 
.A(n_1329),
.Y(n_1463)
);

NAND2xp5_ASAP7_75t_L g1464 ( 
.A(n_1196),
.B(n_1080),
.Y(n_1464)
);

INVx1_ASAP7_75t_L g1465 ( 
.A(n_1330),
.Y(n_1465)
);

INVx2_ASAP7_75t_L g1466 ( 
.A(n_1295),
.Y(n_1466)
);

BUFx6f_ASAP7_75t_L g1467 ( 
.A(n_1227),
.Y(n_1467)
);

INVx2_ASAP7_75t_L g1468 ( 
.A(n_1295),
.Y(n_1468)
);

AOI22xp5_ASAP7_75t_L g1469 ( 
.A1(n_1196),
.A2(n_798),
.B1(n_792),
.B2(n_1050),
.Y(n_1469)
);

CKINVDCx20_ASAP7_75t_R g1470 ( 
.A(n_1266),
.Y(n_1470)
);

NAND2xp5_ASAP7_75t_L g1471 ( 
.A(n_1212),
.B(n_1123),
.Y(n_1471)
);

AND2x2_ASAP7_75t_L g1472 ( 
.A(n_1263),
.B(n_1121),
.Y(n_1472)
);

CKINVDCx20_ASAP7_75t_R g1473 ( 
.A(n_1322),
.Y(n_1473)
);

INVx1_ASAP7_75t_L g1474 ( 
.A(n_1332),
.Y(n_1474)
);

NAND2xp5_ASAP7_75t_SL g1475 ( 
.A(n_1201),
.B(n_1146),
.Y(n_1475)
);

BUFx6f_ASAP7_75t_L g1476 ( 
.A(n_1236),
.Y(n_1476)
);

NOR2xp33_ASAP7_75t_L g1477 ( 
.A(n_1197),
.B(n_1177),
.Y(n_1477)
);

INVx5_ASAP7_75t_L g1478 ( 
.A(n_1202),
.Y(n_1478)
);

INVx2_ASAP7_75t_L g1479 ( 
.A(n_1324),
.Y(n_1479)
);

INVx1_ASAP7_75t_L g1480 ( 
.A(n_1333),
.Y(n_1480)
);

NAND2xp5_ASAP7_75t_SL g1481 ( 
.A(n_1212),
.B(n_1129),
.Y(n_1481)
);

INVx1_ASAP7_75t_L g1482 ( 
.A(n_1336),
.Y(n_1482)
);

INVx1_ASAP7_75t_L g1483 ( 
.A(n_1271),
.Y(n_1483)
);

OAI22xp33_ASAP7_75t_L g1484 ( 
.A1(n_1217),
.A2(n_1137),
.B1(n_1144),
.B2(n_1129),
.Y(n_1484)
);

NAND2xp5_ASAP7_75t_L g1485 ( 
.A(n_1217),
.B(n_1137),
.Y(n_1485)
);

BUFx6f_ASAP7_75t_L g1486 ( 
.A(n_1236),
.Y(n_1486)
);

AND2x4_ASAP7_75t_L g1487 ( 
.A(n_1355),
.B(n_1284),
.Y(n_1487)
);

INVx1_ASAP7_75t_L g1488 ( 
.A(n_1448),
.Y(n_1488)
);

AND2x2_ASAP7_75t_L g1489 ( 
.A(n_1383),
.B(n_1386),
.Y(n_1489)
);

NAND2xp5_ASAP7_75t_L g1490 ( 
.A(n_1386),
.B(n_1301),
.Y(n_1490)
);

AND2x4_ASAP7_75t_L g1491 ( 
.A(n_1355),
.B(n_1202),
.Y(n_1491)
);

INVx4_ASAP7_75t_L g1492 ( 
.A(n_1374),
.Y(n_1492)
);

AOI22xp33_ASAP7_75t_SL g1493 ( 
.A1(n_1453),
.A2(n_1257),
.B1(n_1185),
.B2(n_1127),
.Y(n_1493)
);

INVx1_ASAP7_75t_L g1494 ( 
.A(n_1449),
.Y(n_1494)
);

INVx1_ASAP7_75t_SL g1495 ( 
.A(n_1369),
.Y(n_1495)
);

INVx1_ASAP7_75t_L g1496 ( 
.A(n_1454),
.Y(n_1496)
);

INVx2_ASAP7_75t_SL g1497 ( 
.A(n_1420),
.Y(n_1497)
);

NOR2xp33_ASAP7_75t_L g1498 ( 
.A(n_1403),
.B(n_1200),
.Y(n_1498)
);

AOI22xp5_ASAP7_75t_L g1499 ( 
.A1(n_1351),
.A2(n_1210),
.B1(n_1209),
.B2(n_1343),
.Y(n_1499)
);

AND2x4_ASAP7_75t_L g1500 ( 
.A(n_1437),
.B(n_1298),
.Y(n_1500)
);

INVx1_ASAP7_75t_L g1501 ( 
.A(n_1463),
.Y(n_1501)
);

INVx1_ASAP7_75t_L g1502 ( 
.A(n_1465),
.Y(n_1502)
);

OR2x2_ASAP7_75t_L g1503 ( 
.A(n_1399),
.B(n_1294),
.Y(n_1503)
);

INVx1_ASAP7_75t_L g1504 ( 
.A(n_1474),
.Y(n_1504)
);

AND2x4_ASAP7_75t_L g1505 ( 
.A(n_1437),
.B(n_1298),
.Y(n_1505)
);

AND2x2_ASAP7_75t_L g1506 ( 
.A(n_1399),
.B(n_1318),
.Y(n_1506)
);

INVx2_ASAP7_75t_L g1507 ( 
.A(n_1381),
.Y(n_1507)
);

BUFx2_ASAP7_75t_L g1508 ( 
.A(n_1413),
.Y(n_1508)
);

INVx1_ASAP7_75t_SL g1509 ( 
.A(n_1455),
.Y(n_1509)
);

AND2x4_ASAP7_75t_L g1510 ( 
.A(n_1447),
.B(n_1304),
.Y(n_1510)
);

INVx2_ASAP7_75t_L g1511 ( 
.A(n_1391),
.Y(n_1511)
);

AND2x2_ASAP7_75t_L g1512 ( 
.A(n_1360),
.B(n_1318),
.Y(n_1512)
);

BUFx6f_ASAP7_75t_L g1513 ( 
.A(n_1382),
.Y(n_1513)
);

INVx4_ASAP7_75t_L g1514 ( 
.A(n_1451),
.Y(n_1514)
);

OAI221xp5_ASAP7_75t_L g1515 ( 
.A1(n_1406),
.A2(n_798),
.B1(n_792),
.B2(n_1285),
.C(n_1281),
.Y(n_1515)
);

INVx2_ASAP7_75t_SL g1516 ( 
.A(n_1451),
.Y(n_1516)
);

AND2x2_ASAP7_75t_L g1517 ( 
.A(n_1360),
.B(n_1270),
.Y(n_1517)
);

NAND2xp5_ASAP7_75t_SL g1518 ( 
.A(n_1426),
.B(n_1304),
.Y(n_1518)
);

BUFx6f_ASAP7_75t_L g1519 ( 
.A(n_1382),
.Y(n_1519)
);

NOR2xp33_ASAP7_75t_L g1520 ( 
.A(n_1401),
.B(n_1305),
.Y(n_1520)
);

AND2x2_ASAP7_75t_L g1521 ( 
.A(n_1357),
.B(n_1359),
.Y(n_1521)
);

INVx2_ASAP7_75t_L g1522 ( 
.A(n_1396),
.Y(n_1522)
);

INVx2_ASAP7_75t_L g1523 ( 
.A(n_1398),
.Y(n_1523)
);

OAI22xp5_ASAP7_75t_L g1524 ( 
.A1(n_1483),
.A2(n_1426),
.B1(n_1427),
.B2(n_1423),
.Y(n_1524)
);

NAND2xp5_ASAP7_75t_SL g1525 ( 
.A(n_1427),
.B(n_1209),
.Y(n_1525)
);

AND2x4_ASAP7_75t_L g1526 ( 
.A(n_1447),
.B(n_1379),
.Y(n_1526)
);

NAND2xp5_ASAP7_75t_SL g1527 ( 
.A(n_1394),
.B(n_1305),
.Y(n_1527)
);

AND2x4_ASAP7_75t_L g1528 ( 
.A(n_1379),
.B(n_1195),
.Y(n_1528)
);

NOR2x1p5_ASAP7_75t_L g1529 ( 
.A(n_1392),
.B(n_1275),
.Y(n_1529)
);

CKINVDCx8_ASAP7_75t_R g1530 ( 
.A(n_1364),
.Y(n_1530)
);

BUFx6f_ASAP7_75t_L g1531 ( 
.A(n_1382),
.Y(n_1531)
);

OR2x2_ASAP7_75t_L g1532 ( 
.A(n_1356),
.B(n_1325),
.Y(n_1532)
);

BUFx6f_ASAP7_75t_L g1533 ( 
.A(n_1461),
.Y(n_1533)
);

INVx1_ASAP7_75t_L g1534 ( 
.A(n_1480),
.Y(n_1534)
);

INVx1_ASAP7_75t_L g1535 ( 
.A(n_1482),
.Y(n_1535)
);

AND2x6_ASAP7_75t_L g1536 ( 
.A(n_1414),
.B(n_1270),
.Y(n_1536)
);

INVx1_ASAP7_75t_L g1537 ( 
.A(n_1352),
.Y(n_1537)
);

OAI22xp33_ASAP7_75t_SL g1538 ( 
.A1(n_1395),
.A2(n_771),
.B1(n_768),
.B2(n_1280),
.Y(n_1538)
);

INVx4_ASAP7_75t_L g1539 ( 
.A(n_1451),
.Y(n_1539)
);

INVxp33_ASAP7_75t_L g1540 ( 
.A(n_1477),
.Y(n_1540)
);

AND2x6_ASAP7_75t_L g1541 ( 
.A(n_1432),
.B(n_1280),
.Y(n_1541)
);

NAND2xp5_ASAP7_75t_L g1542 ( 
.A(n_1407),
.B(n_1306),
.Y(n_1542)
);

INVx4_ASAP7_75t_L g1543 ( 
.A(n_1402),
.Y(n_1543)
);

HB1xp67_ASAP7_75t_L g1544 ( 
.A(n_1472),
.Y(n_1544)
);

NAND2xp5_ASAP7_75t_L g1545 ( 
.A(n_1407),
.B(n_1306),
.Y(n_1545)
);

BUFx6f_ASAP7_75t_L g1546 ( 
.A(n_1461),
.Y(n_1546)
);

INVx3_ASAP7_75t_L g1547 ( 
.A(n_1442),
.Y(n_1547)
);

BUFx3_ASAP7_75t_L g1548 ( 
.A(n_1446),
.Y(n_1548)
);

AND2x4_ASAP7_75t_L g1549 ( 
.A(n_1402),
.B(n_1207),
.Y(n_1549)
);

NAND2xp5_ASAP7_75t_L g1550 ( 
.A(n_1394),
.B(n_1222),
.Y(n_1550)
);

INVx1_ASAP7_75t_L g1551 ( 
.A(n_1358),
.Y(n_1551)
);

AND2x6_ASAP7_75t_L g1552 ( 
.A(n_1438),
.B(n_1466),
.Y(n_1552)
);

BUFx6f_ASAP7_75t_L g1553 ( 
.A(n_1461),
.Y(n_1553)
);

BUFx6f_ASAP7_75t_L g1554 ( 
.A(n_1467),
.Y(n_1554)
);

INVx1_ASAP7_75t_L g1555 ( 
.A(n_1363),
.Y(n_1555)
);

NAND2xp5_ASAP7_75t_L g1556 ( 
.A(n_1423),
.B(n_1222),
.Y(n_1556)
);

NAND2xp5_ASAP7_75t_SL g1557 ( 
.A(n_1377),
.B(n_1241),
.Y(n_1557)
);

BUFx4f_ASAP7_75t_L g1558 ( 
.A(n_1442),
.Y(n_1558)
);

INVx6_ASAP7_75t_L g1559 ( 
.A(n_1440),
.Y(n_1559)
);

BUFx2_ASAP7_75t_L g1560 ( 
.A(n_1473),
.Y(n_1560)
);

INVx1_ASAP7_75t_L g1561 ( 
.A(n_1366),
.Y(n_1561)
);

HB1xp67_ASAP7_75t_L g1562 ( 
.A(n_1445),
.Y(n_1562)
);

INVx4_ASAP7_75t_L g1563 ( 
.A(n_1478),
.Y(n_1563)
);

INVx1_ASAP7_75t_SL g1564 ( 
.A(n_1410),
.Y(n_1564)
);

AND2x2_ASAP7_75t_L g1565 ( 
.A(n_1368),
.B(n_1292),
.Y(n_1565)
);

INVx4_ASAP7_75t_L g1566 ( 
.A(n_1364),
.Y(n_1566)
);

AND2x4_ASAP7_75t_L g1567 ( 
.A(n_1429),
.B(n_1292),
.Y(n_1567)
);

INVx1_ASAP7_75t_L g1568 ( 
.A(n_1367),
.Y(n_1568)
);

INVx2_ASAP7_75t_L g1569 ( 
.A(n_1400),
.Y(n_1569)
);

INVx2_ASAP7_75t_L g1570 ( 
.A(n_1404),
.Y(n_1570)
);

NAND2xp5_ASAP7_75t_L g1571 ( 
.A(n_1405),
.B(n_1471),
.Y(n_1571)
);

INVx1_ASAP7_75t_L g1572 ( 
.A(n_1373),
.Y(n_1572)
);

INVx4_ASAP7_75t_L g1573 ( 
.A(n_1478),
.Y(n_1573)
);

INVxp67_ASAP7_75t_SL g1574 ( 
.A(n_1467),
.Y(n_1574)
);

AND2x4_ASAP7_75t_L g1575 ( 
.A(n_1364),
.B(n_1216),
.Y(n_1575)
);

BUFx6f_ASAP7_75t_L g1576 ( 
.A(n_1467),
.Y(n_1576)
);

INVx4_ASAP7_75t_L g1577 ( 
.A(n_1478),
.Y(n_1577)
);

INVx2_ASAP7_75t_L g1578 ( 
.A(n_1353),
.Y(n_1578)
);

INVx2_ASAP7_75t_L g1579 ( 
.A(n_1354),
.Y(n_1579)
);

INVx1_ASAP7_75t_L g1580 ( 
.A(n_1376),
.Y(n_1580)
);

INVx2_ASAP7_75t_L g1581 ( 
.A(n_1361),
.Y(n_1581)
);

AOI21x1_ASAP7_75t_L g1582 ( 
.A1(n_1444),
.A2(n_1231),
.B(n_1311),
.Y(n_1582)
);

BUFx6f_ASAP7_75t_L g1583 ( 
.A(n_1476),
.Y(n_1583)
);

NAND2xp5_ASAP7_75t_L g1584 ( 
.A(n_1489),
.B(n_1351),
.Y(n_1584)
);

OR2x6_ASAP7_75t_L g1585 ( 
.A(n_1548),
.B(n_1384),
.Y(n_1585)
);

INVx2_ASAP7_75t_L g1586 ( 
.A(n_1507),
.Y(n_1586)
);

INVx1_ASAP7_75t_L g1587 ( 
.A(n_1488),
.Y(n_1587)
);

INVx1_ASAP7_75t_L g1588 ( 
.A(n_1494),
.Y(n_1588)
);

INVx2_ASAP7_75t_L g1589 ( 
.A(n_1511),
.Y(n_1589)
);

INVx1_ASAP7_75t_L g1590 ( 
.A(n_1496),
.Y(n_1590)
);

INVx2_ASAP7_75t_L g1591 ( 
.A(n_1522),
.Y(n_1591)
);

NAND2xp5_ASAP7_75t_L g1592 ( 
.A(n_1490),
.B(n_1388),
.Y(n_1592)
);

NAND2xp5_ASAP7_75t_L g1593 ( 
.A(n_1520),
.B(n_1388),
.Y(n_1593)
);

NAND2xp5_ASAP7_75t_L g1594 ( 
.A(n_1498),
.B(n_1388),
.Y(n_1594)
);

NAND2xp5_ASAP7_75t_SL g1595 ( 
.A(n_1540),
.B(n_1435),
.Y(n_1595)
);

BUFx6f_ASAP7_75t_L g1596 ( 
.A(n_1514),
.Y(n_1596)
);

NOR2xp33_ASAP7_75t_L g1597 ( 
.A(n_1508),
.B(n_1462),
.Y(n_1597)
);

NOR2xp33_ASAP7_75t_L g1598 ( 
.A(n_1508),
.B(n_1371),
.Y(n_1598)
);

INVxp67_ASAP7_75t_SL g1599 ( 
.A(n_1487),
.Y(n_1599)
);

INVx2_ASAP7_75t_SL g1600 ( 
.A(n_1558),
.Y(n_1600)
);

NAND2xp5_ASAP7_75t_L g1601 ( 
.A(n_1524),
.B(n_1388),
.Y(n_1601)
);

AOI22xp5_ASAP7_75t_L g1602 ( 
.A1(n_1557),
.A2(n_1377),
.B1(n_1433),
.B2(n_1422),
.Y(n_1602)
);

HB1xp67_ASAP7_75t_L g1603 ( 
.A(n_1495),
.Y(n_1603)
);

NAND2xp5_ASAP7_75t_L g1604 ( 
.A(n_1550),
.B(n_1405),
.Y(n_1604)
);

INVx2_ASAP7_75t_L g1605 ( 
.A(n_1523),
.Y(n_1605)
);

NAND2xp5_ASAP7_75t_SL g1606 ( 
.A(n_1491),
.B(n_1436),
.Y(n_1606)
);

INVx1_ASAP7_75t_L g1607 ( 
.A(n_1501),
.Y(n_1607)
);

NOR2xp33_ASAP7_75t_L g1608 ( 
.A(n_1503),
.B(n_1389),
.Y(n_1608)
);

INVx2_ASAP7_75t_SL g1609 ( 
.A(n_1559),
.Y(n_1609)
);

INVx1_ASAP7_75t_L g1610 ( 
.A(n_1502),
.Y(n_1610)
);

OR2x6_ASAP7_75t_L g1611 ( 
.A(n_1566),
.B(n_1471),
.Y(n_1611)
);

INVx1_ASAP7_75t_L g1612 ( 
.A(n_1504),
.Y(n_1612)
);

OAI21xp5_ASAP7_75t_L g1613 ( 
.A1(n_1571),
.A2(n_1444),
.B(n_1311),
.Y(n_1613)
);

NAND2xp5_ASAP7_75t_SL g1614 ( 
.A(n_1491),
.B(n_1436),
.Y(n_1614)
);

NAND2xp5_ASAP7_75t_SL g1615 ( 
.A(n_1487),
.B(n_1389),
.Y(n_1615)
);

OR2x2_ASAP7_75t_L g1616 ( 
.A(n_1509),
.B(n_1452),
.Y(n_1616)
);

INVx3_ASAP7_75t_L g1617 ( 
.A(n_1530),
.Y(n_1617)
);

NAND2xp5_ASAP7_75t_SL g1618 ( 
.A(n_1526),
.B(n_1428),
.Y(n_1618)
);

NAND2xp5_ASAP7_75t_L g1619 ( 
.A(n_1556),
.B(n_1469),
.Y(n_1619)
);

INVx1_ASAP7_75t_L g1620 ( 
.A(n_1534),
.Y(n_1620)
);

INVx2_ASAP7_75t_SL g1621 ( 
.A(n_1559),
.Y(n_1621)
);

NOR2xp33_ASAP7_75t_L g1622 ( 
.A(n_1564),
.B(n_1412),
.Y(n_1622)
);

HB1xp67_ASAP7_75t_L g1623 ( 
.A(n_1497),
.Y(n_1623)
);

AOI22xp5_ASAP7_75t_L g1624 ( 
.A1(n_1506),
.A2(n_1499),
.B1(n_1525),
.B2(n_1418),
.Y(n_1624)
);

NAND2xp5_ASAP7_75t_L g1625 ( 
.A(n_1542),
.B(n_1469),
.Y(n_1625)
);

OAI21xp33_ASAP7_75t_L g1626 ( 
.A1(n_1515),
.A2(n_952),
.B(n_948),
.Y(n_1626)
);

AOI22xp33_ASAP7_75t_L g1627 ( 
.A1(n_1493),
.A2(n_1418),
.B1(n_1395),
.B2(n_1364),
.Y(n_1627)
);

INVxp33_ASAP7_75t_L g1628 ( 
.A(n_1560),
.Y(n_1628)
);

OR2x2_ASAP7_75t_L g1629 ( 
.A(n_1560),
.B(n_1443),
.Y(n_1629)
);

BUFx3_ASAP7_75t_L g1630 ( 
.A(n_1547),
.Y(n_1630)
);

NAND2xp5_ASAP7_75t_L g1631 ( 
.A(n_1545),
.B(n_1485),
.Y(n_1631)
);

NAND2xp5_ASAP7_75t_L g1632 ( 
.A(n_1512),
.B(n_1485),
.Y(n_1632)
);

INVx5_ASAP7_75t_L g1633 ( 
.A(n_1536),
.Y(n_1633)
);

INVx5_ASAP7_75t_L g1634 ( 
.A(n_1536),
.Y(n_1634)
);

NAND2xp5_ASAP7_75t_L g1635 ( 
.A(n_1517),
.B(n_1418),
.Y(n_1635)
);

INVx1_ASAP7_75t_L g1636 ( 
.A(n_1535),
.Y(n_1636)
);

AOI22xp5_ASAP7_75t_L g1637 ( 
.A1(n_1565),
.A2(n_1418),
.B1(n_1457),
.B2(n_1484),
.Y(n_1637)
);

NOR2x1p5_ASAP7_75t_L g1638 ( 
.A(n_1492),
.B(n_1430),
.Y(n_1638)
);

OAI21xp5_ASAP7_75t_L g1639 ( 
.A1(n_1518),
.A2(n_1464),
.B(n_1481),
.Y(n_1639)
);

AND2x2_ASAP7_75t_L g1640 ( 
.A(n_1544),
.B(n_1567),
.Y(n_1640)
);

INVxp67_ASAP7_75t_L g1641 ( 
.A(n_1562),
.Y(n_1641)
);

NAND2xp5_ASAP7_75t_L g1642 ( 
.A(n_1527),
.B(n_1385),
.Y(n_1642)
);

INVx2_ASAP7_75t_SL g1643 ( 
.A(n_1536),
.Y(n_1643)
);

INVx1_ASAP7_75t_L g1644 ( 
.A(n_1537),
.Y(n_1644)
);

INVx2_ASAP7_75t_L g1645 ( 
.A(n_1586),
.Y(n_1645)
);

NAND2xp5_ASAP7_75t_L g1646 ( 
.A(n_1619),
.B(n_1551),
.Y(n_1646)
);

INVx1_ASAP7_75t_L g1647 ( 
.A(n_1587),
.Y(n_1647)
);

BUFx4f_ASAP7_75t_L g1648 ( 
.A(n_1600),
.Y(n_1648)
);

NOR2xp33_ASAP7_75t_L g1649 ( 
.A(n_1594),
.B(n_1608),
.Y(n_1649)
);

NOR2xp33_ASAP7_75t_L g1650 ( 
.A(n_1593),
.B(n_1538),
.Y(n_1650)
);

INVx2_ASAP7_75t_L g1651 ( 
.A(n_1589),
.Y(n_1651)
);

INVx1_ASAP7_75t_L g1652 ( 
.A(n_1588),
.Y(n_1652)
);

AND2x4_ASAP7_75t_L g1653 ( 
.A(n_1633),
.B(n_1514),
.Y(n_1653)
);

INVx4_ASAP7_75t_L g1654 ( 
.A(n_1633),
.Y(n_1654)
);

INVx5_ASAP7_75t_L g1655 ( 
.A(n_1633),
.Y(n_1655)
);

NAND2xp5_ASAP7_75t_SL g1656 ( 
.A(n_1601),
.B(n_1513),
.Y(n_1656)
);

NAND2xp5_ASAP7_75t_L g1657 ( 
.A(n_1604),
.B(n_1555),
.Y(n_1657)
);

O2A1O1Ixp33_ASAP7_75t_L g1658 ( 
.A1(n_1584),
.A2(n_1464),
.B(n_1457),
.C(n_1458),
.Y(n_1658)
);

INVx3_ASAP7_75t_L g1659 ( 
.A(n_1634),
.Y(n_1659)
);

INVx4_ASAP7_75t_L g1660 ( 
.A(n_1634),
.Y(n_1660)
);

NOR2x1p5_ASAP7_75t_L g1661 ( 
.A(n_1617),
.B(n_1532),
.Y(n_1661)
);

INVx3_ASAP7_75t_L g1662 ( 
.A(n_1634),
.Y(n_1662)
);

INVx2_ASAP7_75t_L g1663 ( 
.A(n_1591),
.Y(n_1663)
);

OR2x2_ASAP7_75t_SL g1664 ( 
.A(n_1629),
.B(n_1529),
.Y(n_1664)
);

INVx1_ASAP7_75t_L g1665 ( 
.A(n_1590),
.Y(n_1665)
);

BUFx3_ASAP7_75t_L g1666 ( 
.A(n_1630),
.Y(n_1666)
);

INVx1_ASAP7_75t_L g1667 ( 
.A(n_1607),
.Y(n_1667)
);

AND2x6_ASAP7_75t_L g1668 ( 
.A(n_1624),
.B(n_1468),
.Y(n_1668)
);

NAND2xp5_ASAP7_75t_L g1669 ( 
.A(n_1625),
.B(n_1561),
.Y(n_1669)
);

INVx1_ASAP7_75t_L g1670 ( 
.A(n_1610),
.Y(n_1670)
);

AND2x4_ASAP7_75t_L g1671 ( 
.A(n_1617),
.B(n_1539),
.Y(n_1671)
);

OR2x2_ASAP7_75t_L g1672 ( 
.A(n_1603),
.B(n_1568),
.Y(n_1672)
);

BUFx6f_ASAP7_75t_L g1673 ( 
.A(n_1596),
.Y(n_1673)
);

INVx4_ASAP7_75t_L g1674 ( 
.A(n_1596),
.Y(n_1674)
);

INVx1_ASAP7_75t_L g1675 ( 
.A(n_1612),
.Y(n_1675)
);

INVx2_ASAP7_75t_L g1676 ( 
.A(n_1605),
.Y(n_1676)
);

INVx1_ASAP7_75t_L g1677 ( 
.A(n_1620),
.Y(n_1677)
);

INVx2_ASAP7_75t_SL g1678 ( 
.A(n_1609),
.Y(n_1678)
);

OR2x2_ASAP7_75t_SL g1679 ( 
.A(n_1623),
.B(n_1470),
.Y(n_1679)
);

BUFx4f_ASAP7_75t_L g1680 ( 
.A(n_1585),
.Y(n_1680)
);

NAND2xp5_ASAP7_75t_L g1681 ( 
.A(n_1631),
.B(n_1572),
.Y(n_1681)
);

INVx3_ASAP7_75t_L g1682 ( 
.A(n_1596),
.Y(n_1682)
);

AOI22xp5_ASAP7_75t_L g1683 ( 
.A1(n_1597),
.A2(n_1541),
.B1(n_1567),
.B2(n_1500),
.Y(n_1683)
);

CKINVDCx5p33_ASAP7_75t_R g1684 ( 
.A(n_1585),
.Y(n_1684)
);

INVx1_ASAP7_75t_SL g1685 ( 
.A(n_1640),
.Y(n_1685)
);

AND2x2_ASAP7_75t_L g1686 ( 
.A(n_1685),
.B(n_1598),
.Y(n_1686)
);

CKINVDCx5p33_ASAP7_75t_R g1687 ( 
.A(n_1666),
.Y(n_1687)
);

INVx1_ASAP7_75t_L g1688 ( 
.A(n_1647),
.Y(n_1688)
);

AOI221xp5_ASAP7_75t_L g1689 ( 
.A1(n_1649),
.A2(n_1626),
.B1(n_1595),
.B2(n_1627),
.C(n_1602),
.Y(n_1689)
);

NAND2xp5_ASAP7_75t_L g1690 ( 
.A(n_1649),
.B(n_1599),
.Y(n_1690)
);

A2O1A1Ixp33_ASAP7_75t_L g1691 ( 
.A1(n_1650),
.A2(n_1602),
.B(n_1626),
.C(n_1637),
.Y(n_1691)
);

INVx4_ASAP7_75t_L g1692 ( 
.A(n_1648),
.Y(n_1692)
);

NAND3xp33_ASAP7_75t_L g1693 ( 
.A(n_1650),
.B(n_1637),
.C(n_1615),
.Y(n_1693)
);

NOR2xp33_ASAP7_75t_R g1694 ( 
.A(n_1684),
.B(n_1277),
.Y(n_1694)
);

NOR2xp33_ASAP7_75t_L g1695 ( 
.A(n_1678),
.B(n_1628),
.Y(n_1695)
);

NAND2xp5_ASAP7_75t_SL g1696 ( 
.A(n_1655),
.B(n_1592),
.Y(n_1696)
);

NAND2xp5_ASAP7_75t_L g1697 ( 
.A(n_1657),
.B(n_1636),
.Y(n_1697)
);

AOI22xp33_ASAP7_75t_L g1698 ( 
.A1(n_1668),
.A2(n_1614),
.B1(n_1606),
.B2(n_1616),
.Y(n_1698)
);

AOI21xp5_ASAP7_75t_L g1699 ( 
.A1(n_1657),
.A2(n_1613),
.B(n_1618),
.Y(n_1699)
);

NAND2xp5_ASAP7_75t_L g1700 ( 
.A(n_1669),
.B(n_1644),
.Y(n_1700)
);

NOR2xp33_ASAP7_75t_L g1701 ( 
.A(n_1648),
.B(n_1641),
.Y(n_1701)
);

O2A1O1Ixp33_ASAP7_75t_L g1702 ( 
.A1(n_1658),
.A2(n_1312),
.B(n_1397),
.C(n_1390),
.Y(n_1702)
);

NAND2xp5_ASAP7_75t_L g1703 ( 
.A(n_1669),
.B(n_1632),
.Y(n_1703)
);

BUFx3_ASAP7_75t_L g1704 ( 
.A(n_1680),
.Y(n_1704)
);

NOR2xp67_ASAP7_75t_SL g1705 ( 
.A(n_1655),
.B(n_1539),
.Y(n_1705)
);

AOI22xp5_ASAP7_75t_L g1706 ( 
.A1(n_1683),
.A2(n_1624),
.B1(n_1622),
.B2(n_1541),
.Y(n_1706)
);

O2A1O1Ixp5_ASAP7_75t_L g1707 ( 
.A1(n_1656),
.A2(n_1639),
.B(n_1613),
.C(n_1642),
.Y(n_1707)
);

NOR2xp33_ASAP7_75t_L g1708 ( 
.A(n_1685),
.B(n_1621),
.Y(n_1708)
);

NAND2xp5_ASAP7_75t_L g1709 ( 
.A(n_1646),
.B(n_1580),
.Y(n_1709)
);

OR2x6_ASAP7_75t_L g1710 ( 
.A(n_1661),
.B(n_1585),
.Y(n_1710)
);

NAND2xp5_ASAP7_75t_SL g1711 ( 
.A(n_1655),
.B(n_1635),
.Y(n_1711)
);

BUFx2_ASAP7_75t_L g1712 ( 
.A(n_1673),
.Y(n_1712)
);

INVx2_ASAP7_75t_SL g1713 ( 
.A(n_1680),
.Y(n_1713)
);

INVx3_ASAP7_75t_L g1714 ( 
.A(n_1654),
.Y(n_1714)
);

OAI21xp33_ASAP7_75t_SL g1715 ( 
.A1(n_1681),
.A2(n_1638),
.B(n_1611),
.Y(n_1715)
);

NOR2xp33_ASAP7_75t_L g1716 ( 
.A(n_1679),
.B(n_1500),
.Y(n_1716)
);

AOI21xp5_ASAP7_75t_L g1717 ( 
.A1(n_1681),
.A2(n_1611),
.B(n_1574),
.Y(n_1717)
);

INVx1_ASAP7_75t_L g1718 ( 
.A(n_1652),
.Y(n_1718)
);

NAND2xp5_ASAP7_75t_L g1719 ( 
.A(n_1646),
.B(n_1505),
.Y(n_1719)
);

AOI21xp5_ASAP7_75t_L g1720 ( 
.A1(n_1656),
.A2(n_1611),
.B(n_1460),
.Y(n_1720)
);

NAND2xp5_ASAP7_75t_L g1721 ( 
.A(n_1672),
.B(n_1505),
.Y(n_1721)
);

AND2x4_ASAP7_75t_L g1722 ( 
.A(n_1653),
.B(n_1643),
.Y(n_1722)
);

NAND2x1p5_ASAP7_75t_L g1723 ( 
.A(n_1655),
.B(n_1653),
.Y(n_1723)
);

O2A1O1Ixp33_ASAP7_75t_L g1724 ( 
.A1(n_1658),
.A2(n_1411),
.B(n_1419),
.C(n_1409),
.Y(n_1724)
);

AOI22xp5_ASAP7_75t_L g1725 ( 
.A1(n_1671),
.A2(n_1541),
.B1(n_1190),
.B2(n_1510),
.Y(n_1725)
);

O2A1O1Ixp5_ASAP7_75t_L g1726 ( 
.A1(n_1674),
.A2(n_1387),
.B(n_1393),
.C(n_1365),
.Y(n_1726)
);

AND2x6_ASAP7_75t_L g1727 ( 
.A(n_1659),
.B(n_1575),
.Y(n_1727)
);

NAND2xp33_ASAP7_75t_L g1728 ( 
.A(n_1691),
.B(n_1673),
.Y(n_1728)
);

AOI222xp33_ASAP7_75t_L g1729 ( 
.A1(n_1689),
.A2(n_768),
.B1(n_749),
.B2(n_778),
.C1(n_751),
.C2(n_746),
.Y(n_1729)
);

NAND2xp5_ASAP7_75t_L g1730 ( 
.A(n_1690),
.B(n_1665),
.Y(n_1730)
);

BUFx6f_ASAP7_75t_L g1731 ( 
.A(n_1704),
.Y(n_1731)
);

NOR2xp67_ASAP7_75t_L g1732 ( 
.A(n_1692),
.B(n_1674),
.Y(n_1732)
);

BUFx3_ASAP7_75t_L g1733 ( 
.A(n_1687),
.Y(n_1733)
);

HB1xp67_ASAP7_75t_L g1734 ( 
.A(n_1688),
.Y(n_1734)
);

AND2x4_ASAP7_75t_L g1735 ( 
.A(n_1710),
.B(n_1673),
.Y(n_1735)
);

AOI22xp33_ASAP7_75t_L g1736 ( 
.A1(n_1693),
.A2(n_1668),
.B1(n_1149),
.B2(n_1054),
.Y(n_1736)
);

INVx1_ASAP7_75t_L g1737 ( 
.A(n_1718),
.Y(n_1737)
);

BUFx2_ASAP7_75t_L g1738 ( 
.A(n_1712),
.Y(n_1738)
);

HAxp5_ASAP7_75t_L g1739 ( 
.A(n_1695),
.B(n_7),
.CON(n_1739),
.SN(n_1739)
);

AO31x2_ASAP7_75t_L g1740 ( 
.A1(n_1720),
.A2(n_1479),
.A3(n_1670),
.B(n_1667),
.Y(n_1740)
);

AOI22xp5_ASAP7_75t_L g1741 ( 
.A1(n_1706),
.A2(n_1575),
.B1(n_1671),
.B2(n_1668),
.Y(n_1741)
);

INVx5_ASAP7_75t_L g1742 ( 
.A(n_1710),
.Y(n_1742)
);

INVx4_ASAP7_75t_L g1743 ( 
.A(n_1692),
.Y(n_1743)
);

INVx1_ASAP7_75t_L g1744 ( 
.A(n_1700),
.Y(n_1744)
);

CKINVDCx20_ASAP7_75t_R g1745 ( 
.A(n_1694),
.Y(n_1745)
);

CKINVDCx8_ASAP7_75t_R g1746 ( 
.A(n_1701),
.Y(n_1746)
);

BUFx6f_ASAP7_75t_L g1747 ( 
.A(n_1713),
.Y(n_1747)
);

AND2x2_ASAP7_75t_L g1748 ( 
.A(n_1686),
.B(n_1675),
.Y(n_1748)
);

INVx3_ASAP7_75t_L g1749 ( 
.A(n_1714),
.Y(n_1749)
);

BUFx2_ASAP7_75t_SL g1750 ( 
.A(n_1722),
.Y(n_1750)
);

AO21x1_ASAP7_75t_L g1751 ( 
.A1(n_1709),
.A2(n_1677),
.B(n_894),
.Y(n_1751)
);

NAND2xp5_ASAP7_75t_L g1752 ( 
.A(n_1703),
.B(n_1668),
.Y(n_1752)
);

NAND2xp5_ASAP7_75t_L g1753 ( 
.A(n_1697),
.B(n_1699),
.Y(n_1753)
);

INVx1_ASAP7_75t_L g1754 ( 
.A(n_1719),
.Y(n_1754)
);

INVx2_ASAP7_75t_L g1755 ( 
.A(n_1721),
.Y(n_1755)
);

INVx2_ASAP7_75t_L g1756 ( 
.A(n_1707),
.Y(n_1756)
);

BUFx6f_ASAP7_75t_L g1757 ( 
.A(n_1722),
.Y(n_1757)
);

AOI22xp33_ASAP7_75t_L g1758 ( 
.A1(n_1698),
.A2(n_1668),
.B1(n_1149),
.B2(n_1054),
.Y(n_1758)
);

NAND2xp5_ASAP7_75t_L g1759 ( 
.A(n_1715),
.B(n_1673),
.Y(n_1759)
);

INVx1_ASAP7_75t_L g1760 ( 
.A(n_1708),
.Y(n_1760)
);

BUFx2_ASAP7_75t_L g1761 ( 
.A(n_1714),
.Y(n_1761)
);

A2O1A1Ixp33_ASAP7_75t_L g1762 ( 
.A1(n_1725),
.A2(n_1430),
.B(n_1460),
.C(n_897),
.Y(n_1762)
);

BUFx3_ASAP7_75t_L g1763 ( 
.A(n_1727),
.Y(n_1763)
);

INVx1_ASAP7_75t_L g1764 ( 
.A(n_1696),
.Y(n_1764)
);

BUFx2_ASAP7_75t_L g1765 ( 
.A(n_1723),
.Y(n_1765)
);

NOR2xp33_ASAP7_75t_L g1766 ( 
.A(n_1716),
.B(n_1664),
.Y(n_1766)
);

INVx2_ASAP7_75t_L g1767 ( 
.A(n_1711),
.Y(n_1767)
);

NAND2xp5_ASAP7_75t_L g1768 ( 
.A(n_1717),
.B(n_1724),
.Y(n_1768)
);

O2A1O1Ixp33_ASAP7_75t_L g1769 ( 
.A1(n_1702),
.A2(n_1439),
.B(n_1431),
.C(n_1726),
.Y(n_1769)
);

INVx1_ASAP7_75t_L g1770 ( 
.A(n_1727),
.Y(n_1770)
);

A2O1A1Ixp33_ASAP7_75t_L g1771 ( 
.A1(n_1736),
.A2(n_901),
.B(n_902),
.C(n_891),
.Y(n_1771)
);

NOR2xp67_ASAP7_75t_L g1772 ( 
.A(n_1753),
.B(n_1682),
.Y(n_1772)
);

AOI21xp5_ASAP7_75t_L g1773 ( 
.A1(n_1768),
.A2(n_1662),
.B(n_1659),
.Y(n_1773)
);

AO31x2_ASAP7_75t_L g1774 ( 
.A1(n_1751),
.A2(n_1651),
.A3(n_1663),
.B(n_1645),
.Y(n_1774)
);

O2A1O1Ixp33_ASAP7_75t_SL g1775 ( 
.A1(n_1745),
.A2(n_1734),
.B(n_1730),
.C(n_1753),
.Y(n_1775)
);

AND2x2_ASAP7_75t_L g1776 ( 
.A(n_1748),
.B(n_1682),
.Y(n_1776)
);

AOI21xp5_ASAP7_75t_L g1777 ( 
.A1(n_1768),
.A2(n_1728),
.B(n_1769),
.Y(n_1777)
);

CKINVDCx20_ASAP7_75t_R g1778 ( 
.A(n_1733),
.Y(n_1778)
);

NAND2xp5_ASAP7_75t_L g1779 ( 
.A(n_1730),
.B(n_903),
.Y(n_1779)
);

AND2x6_ASAP7_75t_L g1780 ( 
.A(n_1763),
.B(n_1741),
.Y(n_1780)
);

NAND2xp5_ASAP7_75t_L g1781 ( 
.A(n_1744),
.B(n_904),
.Y(n_1781)
);

NAND2xp5_ASAP7_75t_L g1782 ( 
.A(n_1734),
.B(n_909),
.Y(n_1782)
);

OAI22xp5_ASAP7_75t_L g1783 ( 
.A1(n_1758),
.A2(n_1662),
.B1(n_1654),
.B2(n_1660),
.Y(n_1783)
);

INVx1_ASAP7_75t_L g1784 ( 
.A(n_1737),
.Y(n_1784)
);

NAND2x1_ASAP7_75t_L g1785 ( 
.A(n_1761),
.B(n_1705),
.Y(n_1785)
);

INVx1_ASAP7_75t_L g1786 ( 
.A(n_1755),
.Y(n_1786)
);

INVx1_ASAP7_75t_L g1787 ( 
.A(n_1754),
.Y(n_1787)
);

O2A1O1Ixp33_ASAP7_75t_L g1788 ( 
.A1(n_1739),
.A2(n_749),
.B(n_751),
.C(n_746),
.Y(n_1788)
);

INVx1_ASAP7_75t_L g1789 ( 
.A(n_1764),
.Y(n_1789)
);

CKINVDCx5p33_ASAP7_75t_R g1790 ( 
.A(n_1746),
.Y(n_1790)
);

BUFx3_ASAP7_75t_L g1791 ( 
.A(n_1731),
.Y(n_1791)
);

OAI221xp5_ASAP7_75t_L g1792 ( 
.A1(n_1766),
.A2(n_820),
.B1(n_787),
.B2(n_778),
.C(n_801),
.Y(n_1792)
);

AOI22xp33_ASAP7_75t_L g1793 ( 
.A1(n_1752),
.A2(n_1552),
.B1(n_1676),
.B2(n_1415),
.Y(n_1793)
);

AOI21xp5_ASAP7_75t_L g1794 ( 
.A1(n_1769),
.A2(n_1756),
.B(n_1759),
.Y(n_1794)
);

INVx2_ASAP7_75t_SL g1795 ( 
.A(n_1731),
.Y(n_1795)
);

NAND3xp33_ASAP7_75t_SL g1796 ( 
.A(n_1729),
.B(n_803),
.C(n_797),
.Y(n_1796)
);

AOI221x1_ASAP7_75t_L g1797 ( 
.A1(n_1760),
.A2(n_1064),
.B1(n_913),
.B2(n_914),
.C(n_912),
.Y(n_1797)
);

BUFx6f_ASAP7_75t_L g1798 ( 
.A(n_1731),
.Y(n_1798)
);

AOI22xp5_ASAP7_75t_L g1799 ( 
.A1(n_1729),
.A2(n_1752),
.B1(n_1750),
.B2(n_1770),
.Y(n_1799)
);

OAI21xp5_ASAP7_75t_L g1800 ( 
.A1(n_1762),
.A2(n_916),
.B(n_910),
.Y(n_1800)
);

INVx2_ASAP7_75t_L g1801 ( 
.A(n_1767),
.Y(n_1801)
);

O2A1O1Ixp33_ASAP7_75t_L g1802 ( 
.A1(n_1759),
.A2(n_787),
.B(n_918),
.C(n_917),
.Y(n_1802)
);

HB1xp67_ASAP7_75t_L g1803 ( 
.A(n_1738),
.Y(n_1803)
);

NOR2xp33_ASAP7_75t_L g1804 ( 
.A(n_1747),
.B(n_8),
.Y(n_1804)
);

INVx1_ASAP7_75t_L g1805 ( 
.A(n_1740),
.Y(n_1805)
);

INVx1_ASAP7_75t_L g1806 ( 
.A(n_1740),
.Y(n_1806)
);

OAI21xp5_ASAP7_75t_L g1807 ( 
.A1(n_1732),
.A2(n_921),
.B(n_920),
.Y(n_1807)
);

AOI21xp5_ASAP7_75t_L g1808 ( 
.A1(n_1749),
.A2(n_1660),
.B(n_1526),
.Y(n_1808)
);

AOI22xp33_ASAP7_75t_L g1809 ( 
.A1(n_1742),
.A2(n_1552),
.B1(n_1417),
.B2(n_1421),
.Y(n_1809)
);

A2O1A1Ixp33_ASAP7_75t_L g1810 ( 
.A1(n_1742),
.A2(n_926),
.B(n_930),
.C(n_925),
.Y(n_1810)
);

OAI21xp5_ASAP7_75t_SL g1811 ( 
.A1(n_1735),
.A2(n_1412),
.B(n_807),
.Y(n_1811)
);

AOI21xp5_ASAP7_75t_L g1812 ( 
.A1(n_1749),
.A2(n_1516),
.B(n_1563),
.Y(n_1812)
);

NAND2xp5_ASAP7_75t_L g1813 ( 
.A(n_1747),
.B(n_931),
.Y(n_1813)
);

A2O1A1Ixp33_ASAP7_75t_L g1814 ( 
.A1(n_1742),
.A2(n_1735),
.B(n_935),
.C(n_936),
.Y(n_1814)
);

OAI21xp5_ASAP7_75t_L g1815 ( 
.A1(n_1743),
.A2(n_938),
.B(n_932),
.Y(n_1815)
);

INVx1_ASAP7_75t_L g1816 ( 
.A(n_1740),
.Y(n_1816)
);

AO32x2_ASAP7_75t_L g1817 ( 
.A1(n_1743),
.A2(n_1563),
.A3(n_1577),
.B1(n_1573),
.B2(n_1543),
.Y(n_1817)
);

INVx2_ASAP7_75t_SL g1818 ( 
.A(n_1747),
.Y(n_1818)
);

OAI221xp5_ASAP7_75t_SL g1819 ( 
.A1(n_1765),
.A2(n_812),
.B1(n_814),
.B2(n_810),
.C(n_806),
.Y(n_1819)
);

AO32x2_ASAP7_75t_L g1820 ( 
.A1(n_1742),
.A2(n_1577),
.A3(n_1573),
.B1(n_1543),
.B2(n_1582),
.Y(n_1820)
);

INVx1_ASAP7_75t_L g1821 ( 
.A(n_1757),
.Y(n_1821)
);

O2A1O1Ixp33_ASAP7_75t_L g1822 ( 
.A1(n_1757),
.A2(n_941),
.B(n_942),
.C(n_939),
.Y(n_1822)
);

AOI21xp5_ASAP7_75t_L g1823 ( 
.A1(n_1757),
.A2(n_1510),
.B(n_1513),
.Y(n_1823)
);

AOI21xp5_ASAP7_75t_L g1824 ( 
.A1(n_1768),
.A2(n_1519),
.B(n_1513),
.Y(n_1824)
);

AOI22xp5_ASAP7_75t_L g1825 ( 
.A1(n_1728),
.A2(n_1727),
.B1(n_1552),
.B2(n_1190),
.Y(n_1825)
);

BUFx2_ASAP7_75t_L g1826 ( 
.A(n_1738),
.Y(n_1826)
);

INVx1_ASAP7_75t_L g1827 ( 
.A(n_1734),
.Y(n_1827)
);

AOI22xp5_ASAP7_75t_L g1828 ( 
.A1(n_1728),
.A2(n_1727),
.B1(n_1528),
.B2(n_1549),
.Y(n_1828)
);

NAND2x1p5_ASAP7_75t_L g1829 ( 
.A(n_1742),
.B(n_1519),
.Y(n_1829)
);

AOI22xp33_ASAP7_75t_L g1830 ( 
.A1(n_1758),
.A2(n_1408),
.B1(n_1425),
.B2(n_1424),
.Y(n_1830)
);

NOR2xp33_ASAP7_75t_L g1831 ( 
.A(n_1746),
.B(n_8),
.Y(n_1831)
);

AOI22xp33_ASAP7_75t_L g1832 ( 
.A1(n_1830),
.A2(n_1456),
.B1(n_1459),
.B2(n_1450),
.Y(n_1832)
);

OA21x2_ASAP7_75t_L g1833 ( 
.A1(n_1794),
.A2(n_1064),
.B(n_816),
.Y(n_1833)
);

INVx1_ASAP7_75t_L g1834 ( 
.A(n_1827),
.Y(n_1834)
);

OR2x2_ASAP7_75t_L g1835 ( 
.A(n_1803),
.B(n_815),
.Y(n_1835)
);

AND2x2_ASAP7_75t_L g1836 ( 
.A(n_1826),
.B(n_1776),
.Y(n_1836)
);

INVx1_ASAP7_75t_SL g1837 ( 
.A(n_1790),
.Y(n_1837)
);

NAND2xp5_ASAP7_75t_L g1838 ( 
.A(n_1789),
.B(n_1141),
.Y(n_1838)
);

AND2x4_ASAP7_75t_L g1839 ( 
.A(n_1772),
.B(n_1093),
.Y(n_1839)
);

INVx2_ASAP7_75t_SL g1840 ( 
.A(n_1791),
.Y(n_1840)
);

BUFx6f_ASAP7_75t_L g1841 ( 
.A(n_1798),
.Y(n_1841)
);

NAND2xp5_ASAP7_75t_L g1842 ( 
.A(n_1787),
.B(n_1141),
.Y(n_1842)
);

OR2x2_ASAP7_75t_L g1843 ( 
.A(n_1784),
.B(n_1137),
.Y(n_1843)
);

AOI22xp5_ASAP7_75t_L g1844 ( 
.A1(n_1780),
.A2(n_1338),
.B1(n_1032),
.B2(n_1528),
.Y(n_1844)
);

INVx1_ASAP7_75t_L g1845 ( 
.A(n_1801),
.Y(n_1845)
);

AOI22xp33_ASAP7_75t_SL g1846 ( 
.A1(n_1780),
.A2(n_1277),
.B1(n_1032),
.B2(n_1521),
.Y(n_1846)
);

AND2x6_ASAP7_75t_L g1847 ( 
.A(n_1828),
.B(n_1583),
.Y(n_1847)
);

CKINVDCx5p33_ASAP7_75t_R g1848 ( 
.A(n_1778),
.Y(n_1848)
);

NOR2xp67_ASAP7_75t_SL g1849 ( 
.A(n_1777),
.B(n_1583),
.Y(n_1849)
);

AOI22xp33_ASAP7_75t_L g1850 ( 
.A1(n_1780),
.A2(n_1799),
.B1(n_1793),
.B2(n_1786),
.Y(n_1850)
);

INVx2_ASAP7_75t_SL g1851 ( 
.A(n_1798),
.Y(n_1851)
);

AOI22xp33_ASAP7_75t_L g1852 ( 
.A1(n_1831),
.A2(n_1579),
.B1(n_1581),
.B2(n_1578),
.Y(n_1852)
);

AND2x6_ASAP7_75t_L g1853 ( 
.A(n_1825),
.B(n_1519),
.Y(n_1853)
);

INVx2_ASAP7_75t_L g1854 ( 
.A(n_1821),
.Y(n_1854)
);

INVx2_ASAP7_75t_L g1855 ( 
.A(n_1805),
.Y(n_1855)
);

OAI22xp33_ASAP7_75t_L g1856 ( 
.A1(n_1797),
.A2(n_1533),
.B1(n_1546),
.B2(n_1531),
.Y(n_1856)
);

CKINVDCx8_ASAP7_75t_R g1857 ( 
.A(n_1804),
.Y(n_1857)
);

AOI22xp5_ASAP7_75t_L g1858 ( 
.A1(n_1811),
.A2(n_1549),
.B1(n_1218),
.B2(n_1226),
.Y(n_1858)
);

AO31x2_ASAP7_75t_L g1859 ( 
.A1(n_1806),
.A2(n_1232),
.A3(n_1238),
.B(n_1221),
.Y(n_1859)
);

AOI22xp33_ASAP7_75t_SL g1860 ( 
.A1(n_1779),
.A2(n_1570),
.B1(n_1569),
.B2(n_1370),
.Y(n_1860)
);

INVx4_ASAP7_75t_L g1861 ( 
.A(n_1795),
.Y(n_1861)
);

AOI22xp5_ASAP7_75t_L g1862 ( 
.A1(n_1783),
.A2(n_1387),
.B1(n_1393),
.B2(n_1365),
.Y(n_1862)
);

INVxp67_ASAP7_75t_L g1863 ( 
.A(n_1782),
.Y(n_1863)
);

AOI22xp33_ASAP7_75t_L g1864 ( 
.A1(n_1796),
.A2(n_1240),
.B1(n_1244),
.B2(n_1236),
.Y(n_1864)
);

CKINVDCx20_ASAP7_75t_R g1865 ( 
.A(n_1818),
.Y(n_1865)
);

AOI22xp33_ASAP7_75t_L g1866 ( 
.A1(n_1809),
.A2(n_1244),
.B1(n_1245),
.B2(n_1240),
.Y(n_1866)
);

INVx3_ASAP7_75t_L g1867 ( 
.A(n_1785),
.Y(n_1867)
);

AOI22xp33_ASAP7_75t_L g1868 ( 
.A1(n_1816),
.A2(n_1244),
.B1(n_1245),
.B2(n_1240),
.Y(n_1868)
);

AND2x4_ASAP7_75t_L g1869 ( 
.A(n_1824),
.B(n_1531),
.Y(n_1869)
);

BUFx3_ASAP7_75t_L g1870 ( 
.A(n_1813),
.Y(n_1870)
);

INVx2_ASAP7_75t_L g1871 ( 
.A(n_1774),
.Y(n_1871)
);

CKINVDCx11_ASAP7_75t_R g1872 ( 
.A(n_1819),
.Y(n_1872)
);

OAI22xp5_ASAP7_75t_L g1873 ( 
.A1(n_1814),
.A2(n_1533),
.B1(n_1546),
.B2(n_1531),
.Y(n_1873)
);

AOI22xp5_ASAP7_75t_L g1874 ( 
.A1(n_1775),
.A2(n_1434),
.B1(n_1441),
.B2(n_1416),
.Y(n_1874)
);

INVx3_ASAP7_75t_L g1875 ( 
.A(n_1829),
.Y(n_1875)
);

AND2x2_ASAP7_75t_L g1876 ( 
.A(n_1773),
.B(n_9),
.Y(n_1876)
);

NOR2xp33_ASAP7_75t_L g1877 ( 
.A(n_1781),
.B(n_11),
.Y(n_1877)
);

INVx1_ASAP7_75t_L g1878 ( 
.A(n_1834),
.Y(n_1878)
);

AOI21x1_ASAP7_75t_L g1879 ( 
.A1(n_1849),
.A2(n_1808),
.B(n_1812),
.Y(n_1879)
);

INVx1_ASAP7_75t_L g1880 ( 
.A(n_1838),
.Y(n_1880)
);

INVx2_ASAP7_75t_L g1881 ( 
.A(n_1855),
.Y(n_1881)
);

INVx3_ASAP7_75t_L g1882 ( 
.A(n_1867),
.Y(n_1882)
);

INVx2_ASAP7_75t_L g1883 ( 
.A(n_1843),
.Y(n_1883)
);

AO31x2_ASAP7_75t_L g1884 ( 
.A1(n_1871),
.A2(n_1845),
.A3(n_1854),
.B(n_1842),
.Y(n_1884)
);

OA21x2_ASAP7_75t_L g1885 ( 
.A1(n_1850),
.A2(n_1807),
.B(n_1815),
.Y(n_1885)
);

INVx2_ASAP7_75t_L g1886 ( 
.A(n_1870),
.Y(n_1886)
);

AND2x2_ASAP7_75t_L g1887 ( 
.A(n_1836),
.B(n_1820),
.Y(n_1887)
);

AOI22xp5_ASAP7_75t_L g1888 ( 
.A1(n_1872),
.A2(n_1810),
.B1(n_1792),
.B2(n_1771),
.Y(n_1888)
);

AND2x4_ASAP7_75t_L g1889 ( 
.A(n_1840),
.B(n_1774),
.Y(n_1889)
);

HB1xp67_ASAP7_75t_L g1890 ( 
.A(n_1863),
.Y(n_1890)
);

OAI22xp5_ASAP7_75t_L g1891 ( 
.A1(n_1876),
.A2(n_1823),
.B1(n_1802),
.B2(n_1800),
.Y(n_1891)
);

INVx1_ASAP7_75t_L g1892 ( 
.A(n_1835),
.Y(n_1892)
);

INVx1_ASAP7_75t_L g1893 ( 
.A(n_1859),
.Y(n_1893)
);

INVx4_ASAP7_75t_SL g1894 ( 
.A(n_1853),
.Y(n_1894)
);

INVx2_ASAP7_75t_L g1895 ( 
.A(n_1859),
.Y(n_1895)
);

OAI21xp5_ASAP7_75t_L g1896 ( 
.A1(n_1877),
.A2(n_1788),
.B(n_1822),
.Y(n_1896)
);

INVx2_ASAP7_75t_L g1897 ( 
.A(n_1859),
.Y(n_1897)
);

O2A1O1Ixp5_ASAP7_75t_L g1898 ( 
.A1(n_1849),
.A2(n_955),
.B(n_958),
.C(n_953),
.Y(n_1898)
);

INVx1_ASAP7_75t_L g1899 ( 
.A(n_1861),
.Y(n_1899)
);

INVx1_ASAP7_75t_L g1900 ( 
.A(n_1869),
.Y(n_1900)
);

NAND2x1p5_ASAP7_75t_L g1901 ( 
.A(n_1833),
.B(n_1820),
.Y(n_1901)
);

HB1xp67_ASAP7_75t_L g1902 ( 
.A(n_1851),
.Y(n_1902)
);

AND2x4_ASAP7_75t_L g1903 ( 
.A(n_1869),
.B(n_12),
.Y(n_1903)
);

AND2x2_ASAP7_75t_L g1904 ( 
.A(n_1865),
.B(n_1820),
.Y(n_1904)
);

INVx2_ASAP7_75t_L g1905 ( 
.A(n_1833),
.Y(n_1905)
);

NOR2xp33_ASAP7_75t_L g1906 ( 
.A(n_1848),
.B(n_1837),
.Y(n_1906)
);

OAI211xp5_ASAP7_75t_L g1907 ( 
.A1(n_1896),
.A2(n_1857),
.B(n_1846),
.C(n_1844),
.Y(n_1907)
);

OAI22xp5_ASAP7_75t_L g1908 ( 
.A1(n_1904),
.A2(n_1874),
.B1(n_1862),
.B2(n_1841),
.Y(n_1908)
);

OAI22xp5_ASAP7_75t_L g1909 ( 
.A1(n_1904),
.A2(n_1841),
.B1(n_1875),
.B2(n_1839),
.Y(n_1909)
);

INVx2_ASAP7_75t_L g1910 ( 
.A(n_1884),
.Y(n_1910)
);

AOI22xp33_ASAP7_75t_L g1911 ( 
.A1(n_1885),
.A2(n_1853),
.B1(n_1847),
.B2(n_1839),
.Y(n_1911)
);

BUFx12f_ASAP7_75t_L g1912 ( 
.A(n_1903),
.Y(n_1912)
);

OAI22xp5_ASAP7_75t_L g1913 ( 
.A1(n_1903),
.A2(n_1841),
.B1(n_1856),
.B2(n_1852),
.Y(n_1913)
);

OAI22xp33_ASAP7_75t_L g1914 ( 
.A1(n_1885),
.A2(n_1873),
.B1(n_1858),
.B2(n_1847),
.Y(n_1914)
);

AOI22xp33_ASAP7_75t_L g1915 ( 
.A1(n_1885),
.A2(n_1853),
.B1(n_1847),
.B2(n_1860),
.Y(n_1915)
);

AND2x6_ASAP7_75t_SL g1916 ( 
.A(n_1906),
.B(n_960),
.Y(n_1916)
);

AOI221x1_ASAP7_75t_SL g1917 ( 
.A1(n_1892),
.A2(n_1880),
.B1(n_1878),
.B2(n_1900),
.C(n_1899),
.Y(n_1917)
);

NAND2xp5_ASAP7_75t_L g1918 ( 
.A(n_1890),
.B(n_1868),
.Y(n_1918)
);

AOI21xp5_ASAP7_75t_L g1919 ( 
.A1(n_1891),
.A2(n_1866),
.B(n_1864),
.Y(n_1919)
);

AOI21xp33_ASAP7_75t_L g1920 ( 
.A1(n_1883),
.A2(n_1832),
.B(n_12),
.Y(n_1920)
);

OAI22xp5_ASAP7_75t_L g1921 ( 
.A1(n_1903),
.A2(n_1546),
.B1(n_1553),
.B2(n_1533),
.Y(n_1921)
);

OAI21x1_ASAP7_75t_L g1922 ( 
.A1(n_1882),
.A2(n_1582),
.B(n_1434),
.Y(n_1922)
);

OAI22xp5_ASAP7_75t_L g1923 ( 
.A1(n_1892),
.A2(n_1554),
.B1(n_1576),
.B2(n_1553),
.Y(n_1923)
);

OR2x2_ASAP7_75t_L g1924 ( 
.A(n_1883),
.B(n_13),
.Y(n_1924)
);

INVx2_ASAP7_75t_L g1925 ( 
.A(n_1884),
.Y(n_1925)
);

INVx1_ASAP7_75t_L g1926 ( 
.A(n_1884),
.Y(n_1926)
);

BUFx6f_ASAP7_75t_SL g1927 ( 
.A(n_1889),
.Y(n_1927)
);

OR2x2_ASAP7_75t_L g1928 ( 
.A(n_1887),
.B(n_1902),
.Y(n_1928)
);

BUFx6f_ASAP7_75t_L g1929 ( 
.A(n_1879),
.Y(n_1929)
);

AOI22xp33_ASAP7_75t_L g1930 ( 
.A1(n_1888),
.A2(n_1245),
.B1(n_1228),
.B2(n_1216),
.Y(n_1930)
);

AOI21xp33_ASAP7_75t_SL g1931 ( 
.A1(n_1882),
.A2(n_13),
.B(n_14),
.Y(n_1931)
);

AOI22xp33_ASAP7_75t_L g1932 ( 
.A1(n_1886),
.A2(n_1247),
.B1(n_1228),
.B2(n_1324),
.Y(n_1932)
);

HB1xp67_ASAP7_75t_L g1933 ( 
.A(n_1928),
.Y(n_1933)
);

NAND2xp5_ASAP7_75t_L g1934 ( 
.A(n_1917),
.B(n_1887),
.Y(n_1934)
);

INVx2_ASAP7_75t_L g1935 ( 
.A(n_1910),
.Y(n_1935)
);

AND2x2_ASAP7_75t_L g1936 ( 
.A(n_1929),
.B(n_1882),
.Y(n_1936)
);

AND2x2_ASAP7_75t_L g1937 ( 
.A(n_1929),
.B(n_1894),
.Y(n_1937)
);

AO31x2_ASAP7_75t_L g1938 ( 
.A1(n_1925),
.A2(n_1895),
.A3(n_1897),
.B(n_1905),
.Y(n_1938)
);

OR2x2_ASAP7_75t_L g1939 ( 
.A(n_1918),
.B(n_1884),
.Y(n_1939)
);

HB1xp67_ASAP7_75t_L g1940 ( 
.A(n_1929),
.Y(n_1940)
);

HB1xp67_ASAP7_75t_L g1941 ( 
.A(n_1909),
.Y(n_1941)
);

AOI22xp33_ASAP7_75t_L g1942 ( 
.A1(n_1914),
.A2(n_1905),
.B1(n_1901),
.B2(n_1886),
.Y(n_1942)
);

INVx1_ASAP7_75t_L g1943 ( 
.A(n_1924),
.Y(n_1943)
);

BUFx2_ASAP7_75t_L g1944 ( 
.A(n_1912),
.Y(n_1944)
);

INVx1_ASAP7_75t_L g1945 ( 
.A(n_1926),
.Y(n_1945)
);

NAND2xp5_ASAP7_75t_L g1946 ( 
.A(n_1908),
.B(n_1884),
.Y(n_1946)
);

BUFx2_ASAP7_75t_L g1947 ( 
.A(n_1922),
.Y(n_1947)
);

HB1xp67_ASAP7_75t_L g1948 ( 
.A(n_1913),
.Y(n_1948)
);

NAND2xp5_ASAP7_75t_L g1949 ( 
.A(n_1931),
.B(n_1889),
.Y(n_1949)
);

BUFx6f_ASAP7_75t_L g1950 ( 
.A(n_1916),
.Y(n_1950)
);

AND2x4_ASAP7_75t_L g1951 ( 
.A(n_1911),
.B(n_1894),
.Y(n_1951)
);

AND2x2_ASAP7_75t_L g1952 ( 
.A(n_1915),
.B(n_1894),
.Y(n_1952)
);

NAND2xp5_ASAP7_75t_L g1953 ( 
.A(n_1931),
.B(n_1889),
.Y(n_1953)
);

INVx2_ASAP7_75t_L g1954 ( 
.A(n_1927),
.Y(n_1954)
);

AND2x2_ASAP7_75t_L g1955 ( 
.A(n_1923),
.B(n_1894),
.Y(n_1955)
);

INVx1_ASAP7_75t_L g1956 ( 
.A(n_1927),
.Y(n_1956)
);

AND2x2_ASAP7_75t_L g1957 ( 
.A(n_1921),
.B(n_1879),
.Y(n_1957)
);

INVx1_ASAP7_75t_L g1958 ( 
.A(n_1919),
.Y(n_1958)
);

BUFx6f_ASAP7_75t_L g1959 ( 
.A(n_1907),
.Y(n_1959)
);

OR2x2_ASAP7_75t_SL g1960 ( 
.A(n_1920),
.B(n_1881),
.Y(n_1960)
);

INVx1_ASAP7_75t_L g1961 ( 
.A(n_1930),
.Y(n_1961)
);

AND2x2_ASAP7_75t_L g1962 ( 
.A(n_1932),
.B(n_1901),
.Y(n_1962)
);

INVx1_ASAP7_75t_L g1963 ( 
.A(n_1924),
.Y(n_1963)
);

NAND2xp5_ASAP7_75t_L g1964 ( 
.A(n_1917),
.B(n_1901),
.Y(n_1964)
);

INVx1_ASAP7_75t_L g1965 ( 
.A(n_1943),
.Y(n_1965)
);

OAI22xp5_ASAP7_75t_L g1966 ( 
.A1(n_1934),
.A2(n_1881),
.B1(n_1893),
.B2(n_1895),
.Y(n_1966)
);

AND2x2_ASAP7_75t_L g1967 ( 
.A(n_1944),
.B(n_1898),
.Y(n_1967)
);

AND2x4_ASAP7_75t_L g1968 ( 
.A(n_1944),
.B(n_1893),
.Y(n_1968)
);

INVx2_ASAP7_75t_L g1969 ( 
.A(n_1940),
.Y(n_1969)
);

AND2x2_ASAP7_75t_L g1970 ( 
.A(n_1933),
.B(n_1817),
.Y(n_1970)
);

AOI22xp5_ASAP7_75t_L g1971 ( 
.A1(n_1959),
.A2(n_1958),
.B1(n_1950),
.B2(n_1948),
.Y(n_1971)
);

OAI22xp5_ASAP7_75t_L g1972 ( 
.A1(n_1964),
.A2(n_1897),
.B1(n_962),
.B2(n_964),
.Y(n_1972)
);

AO31x2_ASAP7_75t_L g1973 ( 
.A1(n_1954),
.A2(n_965),
.A3(n_966),
.B(n_961),
.Y(n_1973)
);

INVxp67_ASAP7_75t_L g1974 ( 
.A(n_1950),
.Y(n_1974)
);

AND2x2_ASAP7_75t_L g1975 ( 
.A(n_1937),
.B(n_1817),
.Y(n_1975)
);

INVxp67_ASAP7_75t_SL g1976 ( 
.A(n_1959),
.Y(n_1976)
);

INVx2_ASAP7_75t_L g1977 ( 
.A(n_1963),
.Y(n_1977)
);

OR2x2_ASAP7_75t_L g1978 ( 
.A(n_1949),
.B(n_15),
.Y(n_1978)
);

INVx2_ASAP7_75t_L g1979 ( 
.A(n_1936),
.Y(n_1979)
);

NAND3xp33_ASAP7_75t_SL g1980 ( 
.A(n_1942),
.B(n_968),
.C(n_967),
.Y(n_1980)
);

AOI222xp33_ASAP7_75t_L g1981 ( 
.A1(n_1959),
.A2(n_976),
.B1(n_981),
.B2(n_983),
.C1(n_985),
.C2(n_986),
.Y(n_1981)
);

OAI21xp5_ASAP7_75t_L g1982 ( 
.A1(n_1953),
.A2(n_973),
.B(n_970),
.Y(n_1982)
);

AO221x2_ASAP7_75t_L g1983 ( 
.A1(n_1956),
.A2(n_988),
.B1(n_990),
.B2(n_975),
.C(n_974),
.Y(n_1983)
);

OR2x2_ASAP7_75t_L g1984 ( 
.A(n_1941),
.B(n_1954),
.Y(n_1984)
);

INVx1_ASAP7_75t_SL g1985 ( 
.A(n_1950),
.Y(n_1985)
);

AOI22xp33_ASAP7_75t_L g1986 ( 
.A1(n_1959),
.A2(n_1962),
.B1(n_1950),
.B2(n_1952),
.Y(n_1986)
);

OR2x2_ASAP7_75t_L g1987 ( 
.A(n_1984),
.B(n_1960),
.Y(n_1987)
);

AND2x2_ASAP7_75t_L g1988 ( 
.A(n_1967),
.B(n_1937),
.Y(n_1988)
);

AND2x2_ASAP7_75t_L g1989 ( 
.A(n_1979),
.B(n_1936),
.Y(n_1989)
);

AND2x4_ASAP7_75t_SL g1990 ( 
.A(n_1969),
.B(n_1951),
.Y(n_1990)
);

OR2x2_ASAP7_75t_L g1991 ( 
.A(n_1965),
.B(n_1960),
.Y(n_1991)
);

INVx1_ASAP7_75t_L g1992 ( 
.A(n_1977),
.Y(n_1992)
);

HB1xp67_ASAP7_75t_L g1993 ( 
.A(n_1972),
.Y(n_1993)
);

AND2x4_ASAP7_75t_L g1994 ( 
.A(n_1976),
.B(n_1985),
.Y(n_1994)
);

INVx1_ASAP7_75t_L g1995 ( 
.A(n_1973),
.Y(n_1995)
);

AND2x2_ASAP7_75t_L g1996 ( 
.A(n_1968),
.B(n_1952),
.Y(n_1996)
);

NAND2xp5_ASAP7_75t_SL g1997 ( 
.A(n_1971),
.B(n_1951),
.Y(n_1997)
);

OR2x2_ASAP7_75t_L g1998 ( 
.A(n_1978),
.B(n_1961),
.Y(n_1998)
);

AND2x2_ASAP7_75t_L g1999 ( 
.A(n_1968),
.B(n_1951),
.Y(n_1999)
);

AND2x4_ASAP7_75t_SL g2000 ( 
.A(n_1971),
.B(n_1955),
.Y(n_2000)
);

AND2x4_ASAP7_75t_L g2001 ( 
.A(n_1985),
.B(n_1955),
.Y(n_2001)
);

NOR2xp33_ASAP7_75t_L g2002 ( 
.A(n_1994),
.B(n_1974),
.Y(n_2002)
);

OR2x2_ASAP7_75t_L g2003 ( 
.A(n_1987),
.B(n_1966),
.Y(n_2003)
);

INVx1_ASAP7_75t_L g2004 ( 
.A(n_1992),
.Y(n_2004)
);

NAND2xp5_ASAP7_75t_L g2005 ( 
.A(n_1994),
.B(n_1983),
.Y(n_2005)
);

OAI221xp5_ASAP7_75t_SL g2006 ( 
.A1(n_1991),
.A2(n_1986),
.B1(n_1981),
.B2(n_1946),
.C(n_1939),
.Y(n_2006)
);

HB1xp67_ASAP7_75t_L g2007 ( 
.A(n_1988),
.Y(n_2007)
);

OAI33xp33_ASAP7_75t_L g2008 ( 
.A1(n_1997),
.A2(n_1939),
.A3(n_1945),
.B1(n_1935),
.B2(n_1981),
.B3(n_1983),
.Y(n_2008)
);

NAND2xp5_ASAP7_75t_L g2009 ( 
.A(n_1993),
.B(n_1973),
.Y(n_2009)
);

AOI22xp33_ASAP7_75t_L g2010 ( 
.A1(n_1993),
.A2(n_1962),
.B1(n_1975),
.B2(n_1957),
.Y(n_2010)
);

OR2x2_ASAP7_75t_L g2011 ( 
.A(n_2007),
.B(n_2001),
.Y(n_2011)
);

AND2x2_ASAP7_75t_L g2012 ( 
.A(n_2002),
.B(n_1989),
.Y(n_2012)
);

AND2x2_ASAP7_75t_L g2013 ( 
.A(n_2005),
.B(n_2001),
.Y(n_2013)
);

INVx2_ASAP7_75t_L g2014 ( 
.A(n_2009),
.Y(n_2014)
);

INVx1_ASAP7_75t_L g2015 ( 
.A(n_2004),
.Y(n_2015)
);

INVx1_ASAP7_75t_L g2016 ( 
.A(n_2003),
.Y(n_2016)
);

NAND2xp5_ASAP7_75t_L g2017 ( 
.A(n_2010),
.B(n_2000),
.Y(n_2017)
);

NOR2xp33_ASAP7_75t_L g2018 ( 
.A(n_2011),
.B(n_1997),
.Y(n_2018)
);

NAND2xp5_ASAP7_75t_L g2019 ( 
.A(n_2016),
.B(n_1973),
.Y(n_2019)
);

AOI31xp33_ASAP7_75t_L g2020 ( 
.A1(n_2016),
.A2(n_2017),
.A3(n_2012),
.B(n_2013),
.Y(n_2020)
);

NAND5xp2_ASAP7_75t_L g2021 ( 
.A(n_2015),
.B(n_2006),
.C(n_1996),
.D(n_1999),
.E(n_2000),
.Y(n_2021)
);

OAI21xp5_ASAP7_75t_L g2022 ( 
.A1(n_2014),
.A2(n_1957),
.B(n_1998),
.Y(n_2022)
);

INVx1_ASAP7_75t_L g2023 ( 
.A(n_2019),
.Y(n_2023)
);

INVx2_ASAP7_75t_L g2024 ( 
.A(n_2018),
.Y(n_2024)
);

AND2x2_ASAP7_75t_L g2025 ( 
.A(n_2022),
.B(n_1990),
.Y(n_2025)
);

AOI211xp5_ASAP7_75t_L g2026 ( 
.A1(n_2024),
.A2(n_2021),
.B(n_2008),
.C(n_1995),
.Y(n_2026)
);

NAND3xp33_ASAP7_75t_L g2027 ( 
.A(n_2024),
.B(n_2020),
.C(n_1982),
.Y(n_2027)
);

OAI22xp5_ASAP7_75t_L g2028 ( 
.A1(n_2027),
.A2(n_2025),
.B1(n_2023),
.B2(n_1970),
.Y(n_2028)
);

INVx1_ASAP7_75t_L g2029 ( 
.A(n_2026),
.Y(n_2029)
);

AOI222xp33_ASAP7_75t_L g2030 ( 
.A1(n_2027),
.A2(n_1980),
.B1(n_1935),
.B2(n_1947),
.C1(n_991),
.C2(n_1938),
.Y(n_2030)
);

INVx2_ASAP7_75t_L g2031 ( 
.A(n_2029),
.Y(n_2031)
);

HB1xp67_ASAP7_75t_L g2032 ( 
.A(n_2028),
.Y(n_2032)
);

INVx1_ASAP7_75t_L g2033 ( 
.A(n_2032),
.Y(n_2033)
);

INVx1_ASAP7_75t_L g2034 ( 
.A(n_2031),
.Y(n_2034)
);

INVx1_ASAP7_75t_L g2035 ( 
.A(n_2032),
.Y(n_2035)
);

NAND3xp33_ASAP7_75t_SL g2036 ( 
.A(n_2033),
.B(n_2030),
.C(n_1947),
.Y(n_2036)
);

NOR3x1_ASAP7_75t_L g2037 ( 
.A(n_2035),
.B(n_15),
.C(n_18),
.Y(n_2037)
);

OAI21xp5_ASAP7_75t_SL g2038 ( 
.A1(n_2034),
.A2(n_1163),
.B(n_1144),
.Y(n_2038)
);

BUFx12f_ASAP7_75t_L g2039 ( 
.A(n_2034),
.Y(n_2039)
);

NAND2xp5_ASAP7_75t_SL g2040 ( 
.A(n_2039),
.B(n_1144),
.Y(n_2040)
);

NOR3xp33_ASAP7_75t_L g2041 ( 
.A(n_2036),
.B(n_1475),
.C(n_1072),
.Y(n_2041)
);

INVx1_ASAP7_75t_L g2042 ( 
.A(n_2037),
.Y(n_2042)
);

NOR2x1_ASAP7_75t_L g2043 ( 
.A(n_2038),
.B(n_1068),
.Y(n_2043)
);

OAI21xp5_ASAP7_75t_L g2044 ( 
.A1(n_2042),
.A2(n_1110),
.B(n_1102),
.Y(n_2044)
);

OAI22xp5_ASAP7_75t_L g2045 ( 
.A1(n_2041),
.A2(n_1178),
.B1(n_1163),
.B2(n_1362),
.Y(n_2045)
);

NOR3xp33_ASAP7_75t_L g2046 ( 
.A(n_2040),
.B(n_1247),
.C(n_1241),
.Y(n_2046)
);

NAND4xp25_ASAP7_75t_L g2047 ( 
.A(n_2043),
.B(n_22),
.C(n_20),
.D(n_21),
.Y(n_2047)
);

INVx1_ASAP7_75t_L g2048 ( 
.A(n_2042),
.Y(n_2048)
);

OA33x2_ASAP7_75t_L g2049 ( 
.A1(n_2042),
.A2(n_20),
.A3(n_22),
.B1(n_26),
.B2(n_27),
.B3(n_28),
.Y(n_2049)
);

AND2x2_ASAP7_75t_L g2050 ( 
.A(n_2042),
.B(n_1938),
.Y(n_2050)
);

AOI221xp5_ASAP7_75t_L g2051 ( 
.A1(n_2042),
.A2(n_1178),
.B1(n_1163),
.B2(n_1375),
.C(n_1372),
.Y(n_2051)
);

INVx2_ASAP7_75t_L g2052 ( 
.A(n_2042),
.Y(n_2052)
);

O2A1O1Ixp33_ASAP7_75t_SL g2053 ( 
.A1(n_2042),
.A2(n_32),
.B(n_29),
.C(n_30),
.Y(n_2053)
);

INVxp67_ASAP7_75t_L g2054 ( 
.A(n_2042),
.Y(n_2054)
);

OAI22xp5_ASAP7_75t_L g2055 ( 
.A1(n_2042),
.A2(n_1178),
.B1(n_1380),
.B2(n_1378),
.Y(n_2055)
);

INVx1_ASAP7_75t_L g2056 ( 
.A(n_2042),
.Y(n_2056)
);

INVxp33_ASAP7_75t_SL g2057 ( 
.A(n_2052),
.Y(n_2057)
);

NAND2xp5_ASAP7_75t_L g2058 ( 
.A(n_2054),
.B(n_1938),
.Y(n_2058)
);

NAND2x1p5_ASAP7_75t_L g2059 ( 
.A(n_2048),
.B(n_1416),
.Y(n_2059)
);

NOR2x1_ASAP7_75t_L g2060 ( 
.A(n_2056),
.B(n_29),
.Y(n_2060)
);

NOR2xp67_ASAP7_75t_L g2061 ( 
.A(n_2047),
.B(n_32),
.Y(n_2061)
);

NOR2xp33_ASAP7_75t_L g2062 ( 
.A(n_2053),
.B(n_33),
.Y(n_2062)
);

NOR2x1_ASAP7_75t_L g2063 ( 
.A(n_2044),
.B(n_33),
.Y(n_2063)
);

NOR2xp33_ASAP7_75t_L g2064 ( 
.A(n_2050),
.B(n_34),
.Y(n_2064)
);

NOR2x1_ASAP7_75t_L g2065 ( 
.A(n_2055),
.B(n_35),
.Y(n_2065)
);

NOR3xp33_ASAP7_75t_L g2066 ( 
.A(n_2051),
.B(n_2045),
.C(n_2046),
.Y(n_2066)
);

INVxp33_ASAP7_75t_L g2067 ( 
.A(n_2049),
.Y(n_2067)
);

AOI211xp5_ASAP7_75t_L g2068 ( 
.A1(n_2054),
.A2(n_41),
.B(n_36),
.C(n_37),
.Y(n_2068)
);

NAND2xp5_ASAP7_75t_SL g2069 ( 
.A(n_2052),
.B(n_521),
.Y(n_2069)
);

NOR2x1_ASAP7_75t_L g2070 ( 
.A(n_2052),
.B(n_37),
.Y(n_2070)
);

INVx1_ASAP7_75t_L g2071 ( 
.A(n_2053),
.Y(n_2071)
);

NOR3xp33_ASAP7_75t_L g2072 ( 
.A(n_2054),
.B(n_1262),
.C(n_524),
.Y(n_2072)
);

NOR3xp33_ASAP7_75t_L g2073 ( 
.A(n_2054),
.B(n_1262),
.C(n_525),
.Y(n_2073)
);

XNOR2x1_ASAP7_75t_L g2074 ( 
.A(n_2052),
.B(n_44),
.Y(n_2074)
);

NOR2xp33_ASAP7_75t_L g2075 ( 
.A(n_2054),
.B(n_44),
.Y(n_2075)
);

NOR2x1_ASAP7_75t_L g2076 ( 
.A(n_2052),
.B(n_47),
.Y(n_2076)
);

AND2x2_ASAP7_75t_L g2077 ( 
.A(n_2052),
.B(n_1938),
.Y(n_2077)
);

NAND5xp2_ASAP7_75t_L g2078 ( 
.A(n_2048),
.B(n_49),
.C(n_47),
.D(n_48),
.E(n_50),
.Y(n_2078)
);

NAND4xp25_ASAP7_75t_L g2079 ( 
.A(n_2054),
.B(n_53),
.C(n_48),
.D(n_49),
.Y(n_2079)
);

NAND3xp33_ASAP7_75t_SL g2080 ( 
.A(n_2052),
.B(n_531),
.C(n_522),
.Y(n_2080)
);

NOR4xp25_ASAP7_75t_L g2081 ( 
.A(n_2054),
.B(n_59),
.C(n_54),
.D(n_58),
.Y(n_2081)
);

AND5x1_ASAP7_75t_L g2082 ( 
.A(n_2051),
.B(n_61),
.C(n_59),
.D(n_60),
.E(n_62),
.Y(n_2082)
);

NOR3xp33_ASAP7_75t_L g2083 ( 
.A(n_2054),
.B(n_537),
.C(n_533),
.Y(n_2083)
);

NAND4xp75_ASAP7_75t_L g2084 ( 
.A(n_2048),
.B(n_68),
.C(n_60),
.D(n_63),
.Y(n_2084)
);

NAND3xp33_ASAP7_75t_SL g2085 ( 
.A(n_2052),
.B(n_543),
.C(n_540),
.Y(n_2085)
);

AND2x2_ASAP7_75t_L g2086 ( 
.A(n_2052),
.B(n_63),
.Y(n_2086)
);

NOR3xp33_ASAP7_75t_L g2087 ( 
.A(n_2054),
.B(n_549),
.C(n_545),
.Y(n_2087)
);

NOR4xp25_ASAP7_75t_L g2088 ( 
.A(n_2054),
.B(n_70),
.C(n_68),
.D(n_69),
.Y(n_2088)
);

INVx1_ASAP7_75t_L g2089 ( 
.A(n_2053),
.Y(n_2089)
);

NAND3xp33_ASAP7_75t_L g2090 ( 
.A(n_2054),
.B(n_555),
.C(n_552),
.Y(n_2090)
);

NOR2xp33_ASAP7_75t_L g2091 ( 
.A(n_2054),
.B(n_69),
.Y(n_2091)
);

NAND2xp5_ASAP7_75t_L g2092 ( 
.A(n_2054),
.B(n_71),
.Y(n_2092)
);

AOI211x1_ASAP7_75t_L g2093 ( 
.A1(n_2056),
.A2(n_75),
.B(n_71),
.C(n_72),
.Y(n_2093)
);

AND2x2_ASAP7_75t_L g2094 ( 
.A(n_2067),
.B(n_76),
.Y(n_2094)
);

NAND4xp75_ASAP7_75t_L g2095 ( 
.A(n_2060),
.B(n_80),
.C(n_78),
.D(n_79),
.Y(n_2095)
);

INVxp67_ASAP7_75t_L g2096 ( 
.A(n_2070),
.Y(n_2096)
);

AOI21xp33_ASAP7_75t_SL g2097 ( 
.A1(n_2057),
.A2(n_78),
.B(n_79),
.Y(n_2097)
);

OAI21xp5_ASAP7_75t_L g2098 ( 
.A1(n_2076),
.A2(n_562),
.B(n_560),
.Y(n_2098)
);

OAI22x1_ASAP7_75t_L g2099 ( 
.A1(n_2071),
.A2(n_85),
.B1(n_82),
.B2(n_83),
.Y(n_2099)
);

INVxp67_ASAP7_75t_L g2100 ( 
.A(n_2062),
.Y(n_2100)
);

AOI211xp5_ASAP7_75t_L g2101 ( 
.A1(n_2081),
.A2(n_85),
.B(n_82),
.C(n_83),
.Y(n_2101)
);

NOR2x1_ASAP7_75t_L g2102 ( 
.A(n_2092),
.B(n_86),
.Y(n_2102)
);

OAI211xp5_ASAP7_75t_L g2103 ( 
.A1(n_2089),
.A2(n_88),
.B(n_86),
.C(n_87),
.Y(n_2103)
);

NAND3x1_ASAP7_75t_L g2104 ( 
.A(n_2083),
.B(n_2087),
.C(n_2075),
.Y(n_2104)
);

OAI211xp5_ASAP7_75t_L g2105 ( 
.A1(n_2088),
.A2(n_89),
.B(n_87),
.C(n_88),
.Y(n_2105)
);

AOI22xp33_ASAP7_75t_L g2106 ( 
.A1(n_2061),
.A2(n_565),
.B1(n_570),
.B2(n_563),
.Y(n_2106)
);

AOI21xp5_ASAP7_75t_L g2107 ( 
.A1(n_2069),
.A2(n_577),
.B(n_574),
.Y(n_2107)
);

OAI211xp5_ASAP7_75t_SL g2108 ( 
.A1(n_2058),
.A2(n_92),
.B(n_90),
.C(n_91),
.Y(n_2108)
);

OAI211xp5_ASAP7_75t_L g2109 ( 
.A1(n_2093),
.A2(n_96),
.B(n_93),
.C(n_95),
.Y(n_2109)
);

OAI221xp5_ASAP7_75t_SL g2110 ( 
.A1(n_2082),
.A2(n_93),
.B1(n_97),
.B2(n_100),
.C(n_101),
.Y(n_2110)
);

O2A1O1Ixp33_ASAP7_75t_L g2111 ( 
.A1(n_2080),
.A2(n_101),
.B(n_97),
.C(n_100),
.Y(n_2111)
);

AOI21xp5_ASAP7_75t_L g2112 ( 
.A1(n_2085),
.A2(n_583),
.B(n_578),
.Y(n_2112)
);

INVx1_ASAP7_75t_L g2113 ( 
.A(n_2086),
.Y(n_2113)
);

NAND2xp5_ASAP7_75t_SL g2114 ( 
.A(n_2068),
.B(n_586),
.Y(n_2114)
);

AND2x4_ASAP7_75t_L g2115 ( 
.A(n_2063),
.B(n_103),
.Y(n_2115)
);

INVx2_ASAP7_75t_L g2116 ( 
.A(n_2074),
.Y(n_2116)
);

OAI21xp33_ASAP7_75t_L g2117 ( 
.A1(n_2078),
.A2(n_593),
.B(n_592),
.Y(n_2117)
);

OAI211xp5_ASAP7_75t_SL g2118 ( 
.A1(n_2064),
.A2(n_103),
.B(n_1441),
.C(n_1315),
.Y(n_2118)
);

OAI21xp33_ASAP7_75t_SL g2119 ( 
.A1(n_2077),
.A2(n_2091),
.B(n_2065),
.Y(n_2119)
);

OAI211xp5_ASAP7_75t_L g2120 ( 
.A1(n_2072),
.A2(n_597),
.B(n_598),
.C(n_594),
.Y(n_2120)
);

NAND2x1p5_ASAP7_75t_L g2121 ( 
.A(n_2084),
.B(n_1476),
.Y(n_2121)
);

NOR3xp33_ASAP7_75t_L g2122 ( 
.A(n_2090),
.B(n_604),
.C(n_599),
.Y(n_2122)
);

A2O1A1Ixp33_ASAP7_75t_L g2123 ( 
.A1(n_2073),
.A2(n_607),
.B(n_609),
.C(n_605),
.Y(n_2123)
);

NAND2xp5_ASAP7_75t_L g2124 ( 
.A(n_2059),
.B(n_2079),
.Y(n_2124)
);

NAND2xp5_ASAP7_75t_L g2125 ( 
.A(n_2066),
.B(n_615),
.Y(n_2125)
);

INVx2_ASAP7_75t_L g2126 ( 
.A(n_2070),
.Y(n_2126)
);

INVx1_ASAP7_75t_L g2127 ( 
.A(n_2060),
.Y(n_2127)
);

OA22x2_ASAP7_75t_L g2128 ( 
.A1(n_2071),
.A2(n_625),
.B1(n_628),
.B2(n_618),
.Y(n_2128)
);

OAI221xp5_ASAP7_75t_L g2129 ( 
.A1(n_2071),
.A2(n_724),
.B1(n_631),
.B2(n_639),
.C(n_641),
.Y(n_2129)
);

INVx1_ASAP7_75t_SL g2130 ( 
.A(n_2086),
.Y(n_2130)
);

INVx1_ASAP7_75t_L g2131 ( 
.A(n_2060),
.Y(n_2131)
);

NOR5xp2_ASAP7_75t_L g2132 ( 
.A(n_2090),
.B(n_731),
.C(n_730),
.D(n_726),
.E(n_725),
.Y(n_2132)
);

HB1xp67_ASAP7_75t_L g2133 ( 
.A(n_2060),
.Y(n_2133)
);

NAND3xp33_ASAP7_75t_L g2134 ( 
.A(n_2060),
.B(n_644),
.C(n_630),
.Y(n_2134)
);

AOI21xp5_ASAP7_75t_L g2135 ( 
.A1(n_2057),
.A2(n_654),
.B(n_653),
.Y(n_2135)
);

BUFx2_ASAP7_75t_L g2136 ( 
.A(n_2060),
.Y(n_2136)
);

AND3x4_ASAP7_75t_L g2137 ( 
.A(n_2061),
.B(n_1817),
.C(n_108),
.Y(n_2137)
);

NAND4xp25_ASAP7_75t_L g2138 ( 
.A(n_2057),
.B(n_1315),
.C(n_712),
.D(n_710),
.Y(n_2138)
);

OAI211xp5_ASAP7_75t_SL g2139 ( 
.A1(n_2071),
.A2(n_707),
.B(n_706),
.C(n_704),
.Y(n_2139)
);

NOR3xp33_ASAP7_75t_SL g2140 ( 
.A(n_2080),
.B(n_662),
.C(n_658),
.Y(n_2140)
);

INVx1_ASAP7_75t_L g2141 ( 
.A(n_2136),
.Y(n_2141)
);

NOR3xp33_ASAP7_75t_L g2142 ( 
.A(n_2130),
.B(n_2113),
.C(n_2116),
.Y(n_2142)
);

NAND2x1p5_ASAP7_75t_L g2143 ( 
.A(n_2094),
.B(n_1476),
.Y(n_2143)
);

INVx1_ASAP7_75t_L g2144 ( 
.A(n_2133),
.Y(n_2144)
);

NOR2xp67_ASAP7_75t_L g2145 ( 
.A(n_2103),
.B(n_113),
.Y(n_2145)
);

NAND2xp5_ASAP7_75t_SL g2146 ( 
.A(n_2097),
.B(n_664),
.Y(n_2146)
);

NOR2xp33_ASAP7_75t_L g2147 ( 
.A(n_2096),
.B(n_665),
.Y(n_2147)
);

INVx1_ASAP7_75t_SL g2148 ( 
.A(n_2115),
.Y(n_2148)
);

AND3x2_ASAP7_75t_L g2149 ( 
.A(n_2100),
.B(n_671),
.C(n_670),
.Y(n_2149)
);

NAND3xp33_ASAP7_75t_L g2150 ( 
.A(n_2127),
.B(n_674),
.C(n_673),
.Y(n_2150)
);

INVx2_ASAP7_75t_L g2151 ( 
.A(n_2115),
.Y(n_2151)
);

AND2x2_ASAP7_75t_L g2152 ( 
.A(n_2131),
.B(n_675),
.Y(n_2152)
);

NOR3xp33_ASAP7_75t_SL g2153 ( 
.A(n_2119),
.B(n_678),
.C(n_677),
.Y(n_2153)
);

NAND5xp2_ASAP7_75t_L g2154 ( 
.A(n_2101),
.B(n_114),
.C(n_115),
.D(n_117),
.E(n_120),
.Y(n_2154)
);

AOI22xp33_ASAP7_75t_R g2155 ( 
.A1(n_2126),
.A2(n_2108),
.B1(n_2110),
.B2(n_2102),
.Y(n_2155)
);

NAND2xp5_ASAP7_75t_L g2156 ( 
.A(n_2117),
.B(n_680),
.Y(n_2156)
);

INVx1_ASAP7_75t_L g2157 ( 
.A(n_2137),
.Y(n_2157)
);

NAND2xp5_ASAP7_75t_L g2158 ( 
.A(n_2106),
.B(n_681),
.Y(n_2158)
);

NOR3xp33_ASAP7_75t_L g2159 ( 
.A(n_2138),
.B(n_684),
.C(n_683),
.Y(n_2159)
);

INVxp67_ASAP7_75t_L g2160 ( 
.A(n_2095),
.Y(n_2160)
);

AOI21xp33_ASAP7_75t_SL g2161 ( 
.A1(n_2099),
.A2(n_686),
.B(n_685),
.Y(n_2161)
);

NOR3xp33_ASAP7_75t_L g2162 ( 
.A(n_2139),
.B(n_690),
.C(n_688),
.Y(n_2162)
);

OR2x2_ASAP7_75t_L g2163 ( 
.A(n_2105),
.B(n_121),
.Y(n_2163)
);

NAND4xp75_ASAP7_75t_L g2164 ( 
.A(n_2098),
.B(n_1231),
.C(n_702),
.D(n_701),
.Y(n_2164)
);

AOI211x1_ASAP7_75t_SL g2165 ( 
.A1(n_2134),
.A2(n_1070),
.B(n_1030),
.C(n_1031),
.Y(n_2165)
);

NOR3xp33_ASAP7_75t_L g2166 ( 
.A(n_2125),
.B(n_696),
.C(n_693),
.Y(n_2166)
);

INVx1_ASAP7_75t_L g2167 ( 
.A(n_2128),
.Y(n_2167)
);

NAND4xp75_ASAP7_75t_L g2168 ( 
.A(n_2135),
.B(n_697),
.C(n_124),
.D(n_126),
.Y(n_2168)
);

NOR4xp75_ASAP7_75t_SL g2169 ( 
.A(n_2104),
.B(n_122),
.C(n_132),
.D(n_139),
.Y(n_2169)
);

INVx1_ASAP7_75t_L g2170 ( 
.A(n_2121),
.Y(n_2170)
);

OR2x2_ASAP7_75t_L g2171 ( 
.A(n_2109),
.B(n_140),
.Y(n_2171)
);

INVx1_ASAP7_75t_L g2172 ( 
.A(n_2124),
.Y(n_2172)
);

AOI21xp5_ASAP7_75t_L g2173 ( 
.A1(n_2112),
.A2(n_1038),
.B(n_1031),
.Y(n_2173)
);

NOR2xp33_ASAP7_75t_R g2174 ( 
.A(n_2132),
.B(n_142),
.Y(n_2174)
);

INVxp67_ASAP7_75t_SL g2175 ( 
.A(n_2107),
.Y(n_2175)
);

NAND5xp2_ASAP7_75t_L g2176 ( 
.A(n_2140),
.B(n_143),
.C(n_146),
.D(n_147),
.E(n_148),
.Y(n_2176)
);

INVx2_ASAP7_75t_L g2177 ( 
.A(n_2114),
.Y(n_2177)
);

NOR3xp33_ASAP7_75t_L g2178 ( 
.A(n_2141),
.B(n_2144),
.C(n_2142),
.Y(n_2178)
);

AND4x1_ASAP7_75t_L g2179 ( 
.A(n_2153),
.B(n_2123),
.C(n_2111),
.D(n_2122),
.Y(n_2179)
);

OA22x2_ASAP7_75t_L g2180 ( 
.A1(n_2149),
.A2(n_2120),
.B1(n_2118),
.B2(n_2129),
.Y(n_2180)
);

XOR2xp5_ASAP7_75t_L g2181 ( 
.A(n_2155),
.B(n_154),
.Y(n_2181)
);

HB1xp67_ASAP7_75t_L g2182 ( 
.A(n_2151),
.Y(n_2182)
);

NOR2x1p5_ASAP7_75t_L g2183 ( 
.A(n_2157),
.B(n_2171),
.Y(n_2183)
);

AO22x2_ASAP7_75t_L g2184 ( 
.A1(n_2148),
.A2(n_159),
.B1(n_161),
.B2(n_162),
.Y(n_2184)
);

BUFx2_ASAP7_75t_L g2185 ( 
.A(n_2174),
.Y(n_2185)
);

AND4x1_ASAP7_75t_L g2186 ( 
.A(n_2172),
.B(n_2159),
.C(n_2170),
.D(n_2147),
.Y(n_2186)
);

NOR4xp75_ASAP7_75t_L g2187 ( 
.A(n_2146),
.B(n_164),
.C(n_170),
.D(n_171),
.Y(n_2187)
);

NOR2xp33_ASAP7_75t_L g2188 ( 
.A(n_2176),
.B(n_174),
.Y(n_2188)
);

INVx1_ASAP7_75t_L g2189 ( 
.A(n_2163),
.Y(n_2189)
);

AOI221x1_ASAP7_75t_L g2190 ( 
.A1(n_2150),
.A2(n_1031),
.B1(n_1038),
.B2(n_1040),
.C(n_1043),
.Y(n_2190)
);

OAI22xp5_ASAP7_75t_L g2191 ( 
.A1(n_2167),
.A2(n_2175),
.B1(n_2160),
.B2(n_2164),
.Y(n_2191)
);

AOI21xp5_ASAP7_75t_L g2192 ( 
.A1(n_2156),
.A2(n_1013),
.B(n_1034),
.Y(n_2192)
);

INVx1_ASAP7_75t_L g2193 ( 
.A(n_2145),
.Y(n_2193)
);

OAI221xp5_ASAP7_75t_L g2194 ( 
.A1(n_2162),
.A2(n_1486),
.B1(n_1583),
.B2(n_1554),
.C(n_1553),
.Y(n_2194)
);

AOI31xp33_ASAP7_75t_L g2195 ( 
.A1(n_2152),
.A2(n_176),
.A3(n_177),
.B(n_181),
.Y(n_2195)
);

OA22x2_ASAP7_75t_L g2196 ( 
.A1(n_2177),
.A2(n_186),
.B1(n_187),
.B2(n_197),
.Y(n_2196)
);

NAND4xp25_ASAP7_75t_L g2197 ( 
.A(n_2154),
.B(n_198),
.C(n_204),
.D(n_205),
.Y(n_2197)
);

AOI211x1_ASAP7_75t_L g2198 ( 
.A1(n_2173),
.A2(n_210),
.B(n_211),
.C(n_212),
.Y(n_2198)
);

NOR2xp33_ASAP7_75t_L g2199 ( 
.A(n_2143),
.B(n_214),
.Y(n_2199)
);

AOI221x1_ASAP7_75t_L g2200 ( 
.A1(n_2166),
.A2(n_1038),
.B1(n_1040),
.B2(n_1043),
.C(n_1051),
.Y(n_2200)
);

AOI22xp5_ASAP7_75t_SL g2201 ( 
.A1(n_2158),
.A2(n_1088),
.B1(n_1114),
.B2(n_1576),
.Y(n_2201)
);

OAI22xp5_ASAP7_75t_L g2202 ( 
.A1(n_2161),
.A2(n_1576),
.B1(n_1554),
.B2(n_1486),
.Y(n_2202)
);

INVx1_ASAP7_75t_L g2203 ( 
.A(n_2165),
.Y(n_2203)
);

XNOR2xp5_ASAP7_75t_L g2204 ( 
.A(n_2168),
.B(n_218),
.Y(n_2204)
);

INVx2_ASAP7_75t_L g2205 ( 
.A(n_2169),
.Y(n_2205)
);

AOI22xp33_ASAP7_75t_L g2206 ( 
.A1(n_2141),
.A2(n_1088),
.B1(n_1114),
.B2(n_1043),
.Y(n_2206)
);

AOI221xp5_ASAP7_75t_L g2207 ( 
.A1(n_2141),
.A2(n_1040),
.B1(n_1067),
.B2(n_1069),
.C(n_1070),
.Y(n_2207)
);

HB1xp67_ASAP7_75t_L g2208 ( 
.A(n_2151),
.Y(n_2208)
);

NOR2x1p5_ASAP7_75t_L g2209 ( 
.A(n_2141),
.B(n_1051),
.Y(n_2209)
);

A2O1A1Ixp33_ASAP7_75t_L g2210 ( 
.A1(n_2144),
.A2(n_1486),
.B(n_1051),
.C(n_1060),
.Y(n_2210)
);

NAND2xp5_ASAP7_75t_L g2211 ( 
.A(n_2178),
.B(n_1088),
.Y(n_2211)
);

INVx2_ASAP7_75t_L g2212 ( 
.A(n_2205),
.Y(n_2212)
);

AOI21xp33_ASAP7_75t_L g2213 ( 
.A1(n_2182),
.A2(n_219),
.B(n_220),
.Y(n_2213)
);

NAND4xp75_ASAP7_75t_L g2214 ( 
.A(n_2193),
.B(n_222),
.C(n_224),
.D(n_225),
.Y(n_2214)
);

AOI211xp5_ASAP7_75t_L g2215 ( 
.A1(n_2208),
.A2(n_1060),
.B(n_1067),
.C(n_1069),
.Y(n_2215)
);

O2A1O1Ixp33_ASAP7_75t_L g2216 ( 
.A1(n_2185),
.A2(n_234),
.B(n_236),
.C(n_240),
.Y(n_2216)
);

XOR2x1_ASAP7_75t_L g2217 ( 
.A(n_2183),
.B(n_242),
.Y(n_2217)
);

NAND2xp5_ASAP7_75t_L g2218 ( 
.A(n_2189),
.B(n_1114),
.Y(n_2218)
);

BUFx2_ASAP7_75t_L g2219 ( 
.A(n_2181),
.Y(n_2219)
);

INVx2_ASAP7_75t_L g2220 ( 
.A(n_2184),
.Y(n_2220)
);

NAND2xp5_ASAP7_75t_L g2221 ( 
.A(n_2188),
.B(n_1114),
.Y(n_2221)
);

OR3x2_ASAP7_75t_L g2222 ( 
.A(n_2197),
.B(n_248),
.C(n_254),
.Y(n_2222)
);

INVx2_ASAP7_75t_L g2223 ( 
.A(n_2184),
.Y(n_2223)
);

INVx2_ASAP7_75t_SL g2224 ( 
.A(n_2196),
.Y(n_2224)
);

AOI21x1_ASAP7_75t_L g2225 ( 
.A1(n_2191),
.A2(n_257),
.B(n_265),
.Y(n_2225)
);

AO22x2_ASAP7_75t_L g2226 ( 
.A1(n_2203),
.A2(n_2200),
.B1(n_2198),
.B2(n_2192),
.Y(n_2226)
);

OAI22xp5_ASAP7_75t_SL g2227 ( 
.A1(n_2204),
.A2(n_1279),
.B1(n_1067),
.B2(n_1069),
.Y(n_2227)
);

BUFx2_ASAP7_75t_L g2228 ( 
.A(n_2180),
.Y(n_2228)
);

INVx1_ASAP7_75t_L g2229 ( 
.A(n_2199),
.Y(n_2229)
);

CKINVDCx20_ASAP7_75t_R g2230 ( 
.A(n_2186),
.Y(n_2230)
);

NAND2xp5_ASAP7_75t_L g2231 ( 
.A(n_2179),
.B(n_268),
.Y(n_2231)
);

INVxp67_ASAP7_75t_SL g2232 ( 
.A(n_2209),
.Y(n_2232)
);

NAND2xp5_ASAP7_75t_L g2233 ( 
.A(n_2195),
.B(n_271),
.Y(n_2233)
);

AND2x2_ASAP7_75t_L g2234 ( 
.A(n_2202),
.B(n_272),
.Y(n_2234)
);

NAND3xp33_ASAP7_75t_L g2235 ( 
.A(n_2228),
.B(n_2207),
.C(n_2201),
.Y(n_2235)
);

OAI221xp5_ASAP7_75t_L g2236 ( 
.A1(n_2224),
.A2(n_2194),
.B1(n_2210),
.B2(n_2206),
.C(n_2187),
.Y(n_2236)
);

NOR2xp67_ASAP7_75t_L g2237 ( 
.A(n_2220),
.B(n_2190),
.Y(n_2237)
);

INVx1_ASAP7_75t_L g2238 ( 
.A(n_2217),
.Y(n_2238)
);

INVx2_ASAP7_75t_L g2239 ( 
.A(n_2230),
.Y(n_2239)
);

OAI22xp5_ASAP7_75t_L g2240 ( 
.A1(n_2212),
.A2(n_1060),
.B1(n_1070),
.B2(n_1013),
.Y(n_2240)
);

NAND3xp33_ASAP7_75t_SL g2241 ( 
.A(n_2219),
.B(n_277),
.C(n_279),
.Y(n_2241)
);

INVx1_ASAP7_75t_L g2242 ( 
.A(n_2223),
.Y(n_2242)
);

INVx2_ASAP7_75t_L g2243 ( 
.A(n_2222),
.Y(n_2243)
);

OAI22x1_ASAP7_75t_L g2244 ( 
.A1(n_2225),
.A2(n_1279),
.B1(n_1074),
.B2(n_1061),
.Y(n_2244)
);

XOR2xp5_ASAP7_75t_L g2245 ( 
.A(n_2229),
.B(n_286),
.Y(n_2245)
);

NOR3xp33_ASAP7_75t_L g2246 ( 
.A(n_2231),
.B(n_290),
.C(n_292),
.Y(n_2246)
);

NOR3xp33_ASAP7_75t_L g2247 ( 
.A(n_2211),
.B(n_300),
.C(n_303),
.Y(n_2247)
);

INVx2_ASAP7_75t_L g2248 ( 
.A(n_2239),
.Y(n_2248)
);

OAI22xp5_ASAP7_75t_SL g2249 ( 
.A1(n_2238),
.A2(n_2232),
.B1(n_2221),
.B2(n_2227),
.Y(n_2249)
);

XNOR2xp5_ASAP7_75t_L g2250 ( 
.A(n_2242),
.B(n_2226),
.Y(n_2250)
);

INVx1_ASAP7_75t_L g2251 ( 
.A(n_2243),
.Y(n_2251)
);

XNOR2xp5_ASAP7_75t_L g2252 ( 
.A(n_2245),
.B(n_2226),
.Y(n_2252)
);

NAND4xp75_ASAP7_75t_L g2253 ( 
.A(n_2237),
.B(n_2233),
.C(n_2218),
.D(n_2234),
.Y(n_2253)
);

INVx2_ASAP7_75t_L g2254 ( 
.A(n_2244),
.Y(n_2254)
);

INVx1_ASAP7_75t_L g2255 ( 
.A(n_2246),
.Y(n_2255)
);

AND4x2_ASAP7_75t_L g2256 ( 
.A(n_2250),
.B(n_2235),
.C(n_2236),
.D(n_2247),
.Y(n_2256)
);

XNOR2x1_ASAP7_75t_L g2257 ( 
.A(n_2248),
.B(n_2252),
.Y(n_2257)
);

INVx1_ASAP7_75t_SL g2258 ( 
.A(n_2251),
.Y(n_2258)
);

OAI222xp33_ASAP7_75t_L g2259 ( 
.A1(n_2255),
.A2(n_2216),
.B1(n_2240),
.B2(n_2241),
.C1(n_2215),
.C2(n_2213),
.Y(n_2259)
);

HB1xp67_ASAP7_75t_L g2260 ( 
.A(n_2257),
.Y(n_2260)
);

NAND2xp5_ASAP7_75t_L g2261 ( 
.A(n_2258),
.B(n_2253),
.Y(n_2261)
);

INVx1_ASAP7_75t_L g2262 ( 
.A(n_2260),
.Y(n_2262)
);

OAI22xp5_ASAP7_75t_L g2263 ( 
.A1(n_2261),
.A2(n_2254),
.B1(n_2249),
.B2(n_2256),
.Y(n_2263)
);

OAI22xp5_ASAP7_75t_L g2264 ( 
.A1(n_2262),
.A2(n_2259),
.B1(n_2214),
.B2(n_1279),
.Y(n_2264)
);

AOI222xp33_ASAP7_75t_L g2265 ( 
.A1(n_2264),
.A2(n_2263),
.B1(n_1340),
.B2(n_1337),
.C1(n_1326),
.C2(n_1317),
.Y(n_2265)
);

AOI22xp33_ASAP7_75t_L g2266 ( 
.A1(n_2265),
.A2(n_1340),
.B1(n_1337),
.B2(n_1326),
.Y(n_2266)
);

INVxp67_ASAP7_75t_L g2267 ( 
.A(n_2266),
.Y(n_2267)
);

OR2x6_ASAP7_75t_L g2268 ( 
.A(n_2267),
.B(n_1256),
.Y(n_2268)
);

AOI21xp5_ASAP7_75t_L g2269 ( 
.A1(n_2268),
.A2(n_1013),
.B(n_1034),
.Y(n_2269)
);

AOI211xp5_ASAP7_75t_L g2270 ( 
.A1(n_2269),
.A2(n_1340),
.B(n_1337),
.C(n_1326),
.Y(n_2270)
);


endmodule