module real_jpeg_25981_n_16 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_3, n_10, n_9, n_16);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_16;

wire n_37;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_300;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_199;
wire n_95;
wire n_238;
wire n_67;
wire n_235;
wire n_107;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_123;
wire n_50;
wire n_186;
wire n_137;
wire n_72;
wire n_171;
wire n_151;
wire n_272;
wire n_198;
wire n_203;
wire n_23;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_326;
wire n_80;
wire n_30;
wire n_332;
wire n_149;
wire n_328;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_230;
wire n_216;
wire n_128;
wire n_202;
wire n_127;
wire n_36;
wire n_102;
wire n_81;
wire n_101;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_252;
wire n_310;
wire n_83;
wire n_78;
wire n_288;
wire n_221;
wire n_104;
wire n_153;
wire n_337;
wire n_131;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_200;
wire n_335;
wire n_214;
wire n_113;
wire n_251;
wire n_139;
wire n_33;
wire n_175;
wire n_156;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_77;
wire n_219;
wire n_122;
wire n_19;
wire n_262;
wire n_334;
wire n_17;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_20;
wire n_278;
wire n_314;
wire n_103;
wire n_232;
wire n_212;
wire n_284;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_213;
wire n_25;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_331;
wire n_49;
wire n_68;
wire n_146;
wire n_286;
wire n_215;
wire n_166;
wire n_176;
wire n_323;
wire n_312;
wire n_325;
wire n_307;
wire n_316;
wire n_161;
wire n_207;
wire n_237;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_140;
wire n_126;
wire n_120;
wire n_155;
wire n_319;
wire n_93;
wire n_242;
wire n_142;
wire n_76;
wire n_79;
wire n_282;
wire n_147;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_18;
wire n_145;
wire n_266;
wire n_109;
wire n_148;
wire n_196;
wire n_298;
wire n_330;
wire n_333;
wire n_152;
wire n_270;
wire n_159;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_336;
wire n_258;
wire n_150;
wire n_41;
wire n_74;
wire n_204;
wire n_158;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_75;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_119;
wire n_283;
wire n_181;
wire n_256;
wire n_253;
wire n_273;
wire n_54;
wire n_168;
wire n_38;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_292;
wire n_64;
wire n_291;
wire n_236;
wire n_276;
wire n_287;
wire n_174;
wire n_255;
wire n_243;
wire n_299;
wire n_56;
wire n_293;
wire n_275;
wire n_227;
wire n_229;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_45;
wire n_268;
wire n_42;
wire n_313;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_143;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_303;
wire n_321;
wire n_100;
wire n_51;
wire n_205;
wire n_261;
wire n_86;
wire n_324;
wire n_70;
wire n_32;
wire n_228;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_169;
wire n_88;
wire n_167;
wire n_295;
wire n_133;
wire n_257;
wire n_210;
wire n_206;
wire n_85;
wire n_96;
wire n_308;

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_0),
.Y(n_29)
);

AOI22xp33_ASAP7_75t_L g168 ( 
.A1(n_1),
.A2(n_58),
.B1(n_59),
.B2(n_169),
.Y(n_168)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_1),
.Y(n_169)
);

AOI21xp5_ASAP7_75t_L g174 ( 
.A1(n_1),
.A2(n_61),
.B(n_66),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_L g178 ( 
.A(n_1),
.B(n_91),
.Y(n_178)
);

OAI22xp5_ASAP7_75t_SL g203 ( 
.A1(n_1),
.A2(n_111),
.B1(n_199),
.B2(n_204),
.Y(n_203)
);

AOI21xp5_ASAP7_75t_L g215 ( 
.A1(n_1),
.A2(n_26),
.B(n_216),
.Y(n_215)
);

NAND2xp5_ASAP7_75t_L g244 ( 
.A(n_1),
.B(n_51),
.Y(n_244)
);

OAI22xp5_ASAP7_75t_L g171 ( 
.A1(n_2),
.A2(n_58),
.B1(n_59),
.B2(n_172),
.Y(n_171)
);

CKINVDCx14_ASAP7_75t_R g172 ( 
.A(n_2),
.Y(n_172)
);

AOI22xp33_ASAP7_75t_L g199 ( 
.A1(n_2),
.A2(n_65),
.B1(n_66),
.B2(n_172),
.Y(n_199)
);

AOI22xp33_ASAP7_75t_L g219 ( 
.A1(n_2),
.A2(n_26),
.B1(n_27),
.B2(n_172),
.Y(n_219)
);

OAI22xp5_ASAP7_75t_SL g282 ( 
.A1(n_2),
.A2(n_37),
.B1(n_38),
.B2(n_172),
.Y(n_282)
);

BUFx12f_ASAP7_75t_L g62 ( 
.A(n_3),
.Y(n_62)
);

OAI22xp5_ASAP7_75t_L g180 ( 
.A1(n_4),
.A2(n_58),
.B1(n_59),
.B2(n_181),
.Y(n_180)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_4),
.Y(n_181)
);

AOI22xp33_ASAP7_75t_L g189 ( 
.A1(n_4),
.A2(n_65),
.B1(n_66),
.B2(n_181),
.Y(n_189)
);

OAI22xp5_ASAP7_75t_L g241 ( 
.A1(n_4),
.A2(n_26),
.B1(n_27),
.B2(n_181),
.Y(n_241)
);

AOI22xp33_ASAP7_75t_SL g294 ( 
.A1(n_4),
.A2(n_37),
.B1(n_46),
.B2(n_181),
.Y(n_294)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_5),
.Y(n_67)
);

INVx8_ASAP7_75t_SL g25 ( 
.A(n_6),
.Y(n_25)
);

OAI22xp5_ASAP7_75t_L g69 ( 
.A1(n_7),
.A2(n_58),
.B1(n_59),
.B2(n_70),
.Y(n_69)
);

CKINVDCx20_ASAP7_75t_R g70 ( 
.A(n_7),
.Y(n_70)
);

AOI22xp5_ASAP7_75t_L g78 ( 
.A1(n_7),
.A2(n_26),
.B1(n_27),
.B2(n_70),
.Y(n_78)
);

OAI22xp5_ASAP7_75t_L g117 ( 
.A1(n_7),
.A2(n_65),
.B1(n_66),
.B2(n_70),
.Y(n_117)
);

OAI22xp5_ASAP7_75t_SL g126 ( 
.A1(n_7),
.A2(n_31),
.B1(n_42),
.B2(n_70),
.Y(n_126)
);

OAI22xp5_ASAP7_75t_SL g36 ( 
.A1(n_8),
.A2(n_37),
.B1(n_40),
.B2(n_41),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_8),
.Y(n_40)
);

OAI22xp5_ASAP7_75t_SL g82 ( 
.A1(n_8),
.A2(n_26),
.B1(n_27),
.B2(n_40),
.Y(n_82)
);

AOI22xp5_ASAP7_75t_L g103 ( 
.A1(n_8),
.A2(n_40),
.B1(n_58),
.B2(n_59),
.Y(n_103)
);

OAI22xp5_ASAP7_75t_SL g144 ( 
.A1(n_8),
.A2(n_40),
.B1(n_65),
.B2(n_66),
.Y(n_144)
);

OAI22xp5_ASAP7_75t_L g52 ( 
.A1(n_9),
.A2(n_38),
.B1(n_42),
.B2(n_53),
.Y(n_52)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_9),
.Y(n_53)
);

OAI22xp5_ASAP7_75t_L g88 ( 
.A1(n_9),
.A2(n_26),
.B1(n_27),
.B2(n_53),
.Y(n_88)
);

AOI22xp5_ASAP7_75t_L g120 ( 
.A1(n_9),
.A2(n_53),
.B1(n_58),
.B2(n_59),
.Y(n_120)
);

OAI22xp5_ASAP7_75t_L g269 ( 
.A1(n_9),
.A2(n_53),
.B1(n_65),
.B2(n_66),
.Y(n_269)
);

BUFx12f_ASAP7_75t_L g76 ( 
.A(n_10),
.Y(n_76)
);

INVx13_ASAP7_75t_L g33 ( 
.A(n_11),
.Y(n_33)
);

NAND2xp5_ASAP7_75t_L g262 ( 
.A(n_11),
.B(n_169),
.Y(n_262)
);

BUFx12f_ASAP7_75t_L g60 ( 
.A(n_12),
.Y(n_60)
);

AOI22xp33_ASAP7_75t_SL g30 ( 
.A1(n_13),
.A2(n_31),
.B1(n_32),
.B2(n_34),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_13),
.Y(n_34)
);

AOI22xp33_ASAP7_75t_SL g106 ( 
.A1(n_13),
.A2(n_26),
.B1(n_27),
.B2(n_34),
.Y(n_106)
);

AOI22xp5_ASAP7_75t_SL g149 ( 
.A1(n_13),
.A2(n_34),
.B1(n_58),
.B2(n_59),
.Y(n_149)
);

AOI22xp33_ASAP7_75t_L g247 ( 
.A1(n_13),
.A2(n_34),
.B1(n_65),
.B2(n_66),
.Y(n_247)
);

AOI22xp5_ASAP7_75t_SL g151 ( 
.A1(n_14),
.A2(n_33),
.B1(n_37),
.B2(n_152),
.Y(n_151)
);

CKINVDCx20_ASAP7_75t_R g152 ( 
.A(n_14),
.Y(n_152)
);

AOI22xp5_ASAP7_75t_L g184 ( 
.A1(n_14),
.A2(n_65),
.B1(n_66),
.B2(n_152),
.Y(n_184)
);

OAI22xp5_ASAP7_75t_L g221 ( 
.A1(n_14),
.A2(n_58),
.B1(n_59),
.B2(n_152),
.Y(n_221)
);

OAI22xp5_ASAP7_75t_L g278 ( 
.A1(n_14),
.A2(n_26),
.B1(n_27),
.B2(n_152),
.Y(n_278)
);

INVx6_ASAP7_75t_L g114 ( 
.A(n_15),
.Y(n_114)
);

INVx2_ASAP7_75t_L g147 ( 
.A(n_15),
.Y(n_147)
);

INVx6_ASAP7_75t_L g192 ( 
.A(n_15),
.Y(n_192)
);

XOR2xp5_ASAP7_75t_L g16 ( 
.A(n_17),
.B(n_130),
.Y(n_16)
);

NAND2xp5_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_128),
.Y(n_17)
);

NAND2xp5_ASAP7_75t_SL g18 ( 
.A(n_19),
.B(n_92),
.Y(n_18)
);

NOR2xp33_ASAP7_75t_L g129 ( 
.A(n_19),
.B(n_92),
.Y(n_129)
);

XNOR2xp5_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_86),
.Y(n_19)
);

AOI22xp5_ASAP7_75t_L g20 ( 
.A1(n_21),
.A2(n_48),
.B1(n_84),
.B2(n_85),
.Y(n_20)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_21),
.Y(n_84)
);

MAJIxp5_ASAP7_75t_L g86 ( 
.A(n_21),
.B(n_55),
.C(n_87),
.Y(n_86)
);

AOI22xp5_ASAP7_75t_L g93 ( 
.A1(n_21),
.A2(n_84),
.B1(n_94),
.B2(n_96),
.Y(n_93)
);

OAI21xp5_ASAP7_75t_L g21 ( 
.A1(n_22),
.A2(n_30),
.B(n_35),
.Y(n_21)
);

NAND2xp5_ASAP7_75t_SL g44 ( 
.A(n_22),
.B(n_45),
.Y(n_44)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_22),
.Y(n_51)
);

OAI22xp5_ASAP7_75t_SL g305 ( 
.A1(n_22),
.A2(n_44),
.B1(n_151),
.B2(n_294),
.Y(n_305)
);

AOI22xp5_ASAP7_75t_L g22 ( 
.A1(n_23),
.A2(n_24),
.B1(n_26),
.B2(n_27),
.Y(n_22)
);

OAI22xp33_ASAP7_75t_L g45 ( 
.A1(n_23),
.A2(n_24),
.B1(n_46),
.B2(n_47),
.Y(n_45)
);

OAI32xp33_ASAP7_75t_L g261 ( 
.A1(n_23),
.A2(n_27),
.A3(n_31),
.B1(n_262),
.B2(n_263),
.Y(n_261)
);

INVx4_ASAP7_75t_L g23 ( 
.A(n_24),
.Y(n_23)
);

NOR2xp33_ASAP7_75t_L g263 ( 
.A(n_24),
.B(n_26),
.Y(n_263)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_25),
.Y(n_24)
);

OAI22xp5_ASAP7_75t_L g81 ( 
.A1(n_26),
.A2(n_27),
.B1(n_76),
.B2(n_77),
.Y(n_81)
);

OAI32xp33_ASAP7_75t_L g225 ( 
.A1(n_26),
.A2(n_59),
.A3(n_76),
.B1(n_217),
.B2(n_226),
.Y(n_225)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_27),
.Y(n_26)
);

NAND2xp5_ASAP7_75t_L g217 ( 
.A(n_27),
.B(n_169),
.Y(n_217)
);

BUFx12f_ASAP7_75t_L g27 ( 
.A(n_28),
.Y(n_27)
);

BUFx12f_ASAP7_75t_L g28 ( 
.A(n_29),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_30),
.Y(n_50)
);

INVx8_ASAP7_75t_L g31 ( 
.A(n_32),
.Y(n_31)
);

INVx11_ASAP7_75t_L g32 ( 
.A(n_33),
.Y(n_32)
);

INVx6_ASAP7_75t_L g39 ( 
.A(n_33),
.Y(n_39)
);

INVx8_ASAP7_75t_L g42 ( 
.A(n_33),
.Y(n_42)
);

INVx8_ASAP7_75t_L g47 ( 
.A(n_33),
.Y(n_47)
);

NAND2xp5_ASAP7_75t_L g35 ( 
.A(n_36),
.B(n_43),
.Y(n_35)
);

NAND2xp5_ASAP7_75t_SL g127 ( 
.A(n_36),
.B(n_51),
.Y(n_127)
);

OAI21xp33_ASAP7_75t_L g281 ( 
.A1(n_37),
.A2(n_169),
.B(n_262),
.Y(n_281)
);

INVx8_ASAP7_75t_L g37 ( 
.A(n_38),
.Y(n_37)
);

INVx8_ASAP7_75t_L g38 ( 
.A(n_39),
.Y(n_38)
);

INVx11_ASAP7_75t_L g41 ( 
.A(n_42),
.Y(n_41)
);

AOI22xp5_ASAP7_75t_L g49 ( 
.A1(n_43),
.A2(n_50),
.B1(n_51),
.B2(n_52),
.Y(n_49)
);

AOI22xp5_ASAP7_75t_SL g280 ( 
.A1(n_43),
.A2(n_51),
.B1(n_281),
.B2(n_282),
.Y(n_280)
);

AOI22xp5_ASAP7_75t_L g292 ( 
.A1(n_43),
.A2(n_51),
.B1(n_282),
.B2(n_293),
.Y(n_292)
);

CKINVDCx16_ASAP7_75t_R g43 ( 
.A(n_44),
.Y(n_43)
);

OAI21xp5_ASAP7_75t_SL g124 ( 
.A1(n_44),
.A2(n_125),
.B(n_127),
.Y(n_124)
);

OAI21xp5_ASAP7_75t_SL g150 ( 
.A1(n_44),
.A2(n_151),
.B(n_153),
.Y(n_150)
);

INVx4_ASAP7_75t_L g46 ( 
.A(n_47),
.Y(n_46)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_48),
.Y(n_85)
);

XNOR2xp5_ASAP7_75t_SL g48 ( 
.A(n_49),
.B(n_54),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_SL g153 ( 
.A(n_51),
.B(n_126),
.Y(n_153)
);

AOI22xp5_ASAP7_75t_L g54 ( 
.A1(n_55),
.A2(n_71),
.B1(n_72),
.B2(n_83),
.Y(n_54)
);

CKINVDCx16_ASAP7_75t_R g83 ( 
.A(n_55),
.Y(n_83)
);

AOI22xp5_ASAP7_75t_L g94 ( 
.A1(n_55),
.A2(n_83),
.B1(n_87),
.B2(n_95),
.Y(n_94)
);

OAI21xp5_ASAP7_75t_SL g55 ( 
.A1(n_56),
.A2(n_68),
.B(n_69),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_L g101 ( 
.A(n_56),
.B(n_102),
.Y(n_101)
);

CKINVDCx20_ASAP7_75t_R g119 ( 
.A(n_56),
.Y(n_119)
);

AOI22xp5_ASAP7_75t_L g179 ( 
.A1(n_56),
.A2(n_68),
.B1(n_171),
.B2(n_180),
.Y(n_179)
);

AOI22xp5_ASAP7_75t_L g220 ( 
.A1(n_56),
.A2(n_68),
.B1(n_180),
.B2(n_221),
.Y(n_220)
);

AOI21xp5_ASAP7_75t_L g279 ( 
.A1(n_56),
.A2(n_69),
.B(n_122),
.Y(n_279)
);

AND2x2_ASAP7_75t_L g56 ( 
.A(n_57),
.B(n_64),
.Y(n_56)
);

OAI22xp33_ASAP7_75t_L g57 ( 
.A1(n_58),
.A2(n_59),
.B1(n_61),
.B2(n_63),
.Y(n_57)
);

AOI22xp5_ASAP7_75t_L g75 ( 
.A1(n_58),
.A2(n_59),
.B1(n_76),
.B2(n_77),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_SL g226 ( 
.A(n_58),
.B(n_77),
.Y(n_226)
);

INVx8_ASAP7_75t_L g58 ( 
.A(n_59),
.Y(n_58)
);

A2O1A1Ixp33_ASAP7_75t_SL g173 ( 
.A1(n_59),
.A2(n_63),
.B(n_169),
.C(n_174),
.Y(n_173)
);

BUFx12f_ASAP7_75t_L g59 ( 
.A(n_60),
.Y(n_59)
);

INVx13_ASAP7_75t_L g63 ( 
.A(n_61),
.Y(n_63)
);

AOI22xp5_ASAP7_75t_L g64 ( 
.A1(n_61),
.A2(n_63),
.B1(n_65),
.B2(n_66),
.Y(n_64)
);

BUFx24_ASAP7_75t_L g61 ( 
.A(n_62),
.Y(n_61)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_64),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g122 ( 
.A(n_64),
.B(n_103),
.Y(n_122)
);

OAI22xp5_ASAP7_75t_L g148 ( 
.A1(n_64),
.A2(n_119),
.B1(n_120),
.B2(n_149),
.Y(n_148)
);

OAI22xp5_ASAP7_75t_L g167 ( 
.A1(n_64),
.A2(n_119),
.B1(n_168),
.B2(n_170),
.Y(n_167)
);

NOR2xp33_ASAP7_75t_SL g197 ( 
.A(n_64),
.B(n_169),
.Y(n_197)
);

OAI21xp5_ASAP7_75t_L g299 ( 
.A1(n_64),
.A2(n_101),
.B(n_149),
.Y(n_299)
);

NOR2xp33_ASAP7_75t_L g112 ( 
.A(n_65),
.B(n_113),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_SL g205 ( 
.A(n_65),
.B(n_206),
.Y(n_205)
);

INVx5_ASAP7_75t_L g65 ( 
.A(n_66),
.Y(n_65)
);

BUFx12f_ASAP7_75t_L g66 ( 
.A(n_67),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_SL g100 ( 
.A(n_68),
.B(n_69),
.Y(n_100)
);

CKINVDCx20_ASAP7_75t_R g71 ( 
.A(n_72),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_L g72 ( 
.A(n_73),
.B(n_79),
.Y(n_72)
);

INVxp67_ASAP7_75t_L g73 ( 
.A(n_74),
.Y(n_73)
);

AOI21xp5_ASAP7_75t_L g291 ( 
.A1(n_74),
.A2(n_80),
.B(n_278),
.Y(n_291)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_75),
.B(n_78),
.Y(n_74)
);

AND2x2_ASAP7_75t_L g80 ( 
.A(n_75),
.B(n_81),
.Y(n_80)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_75),
.Y(n_91)
);

OAI21xp5_ASAP7_75t_L g154 ( 
.A1(n_75),
.A2(n_79),
.B(n_106),
.Y(n_154)
);

OAI22xp5_ASAP7_75t_L g214 ( 
.A1(n_75),
.A2(n_215),
.B1(n_218),
.B2(n_219),
.Y(n_214)
);

INVx5_ASAP7_75t_L g77 ( 
.A(n_76),
.Y(n_77)
);

OAI21xp5_ASAP7_75t_SL g306 ( 
.A1(n_78),
.A2(n_90),
.B(n_218),
.Y(n_306)
);

NAND2xp5_ASAP7_75t_SL g79 ( 
.A(n_80),
.B(n_82),
.Y(n_79)
);

AOI21xp5_ASAP7_75t_L g87 ( 
.A1(n_80),
.A2(n_88),
.B(n_89),
.Y(n_87)
);

AOI22xp5_ASAP7_75t_L g104 ( 
.A1(n_80),
.A2(n_88),
.B1(n_91),
.B2(n_105),
.Y(n_104)
);

CKINVDCx20_ASAP7_75t_R g218 ( 
.A(n_80),
.Y(n_218)
);

AOI22xp5_ASAP7_75t_L g239 ( 
.A1(n_80),
.A2(n_91),
.B1(n_240),
.B2(n_241),
.Y(n_239)
);

AOI22xp5_ASAP7_75t_L g277 ( 
.A1(n_80),
.A2(n_91),
.B1(n_241),
.B2(n_278),
.Y(n_277)
);

NAND2xp5_ASAP7_75t_L g90 ( 
.A(n_82),
.B(n_91),
.Y(n_90)
);

CKINVDCx20_ASAP7_75t_R g95 ( 
.A(n_87),
.Y(n_95)
);

INVxp67_ASAP7_75t_L g89 ( 
.A(n_90),
.Y(n_89)
);

MAJIxp5_ASAP7_75t_L g92 ( 
.A(n_93),
.B(n_97),
.C(n_107),
.Y(n_92)
);

AOI22xp5_ASAP7_75t_L g156 ( 
.A1(n_93),
.A2(n_97),
.B1(n_98),
.B2(n_157),
.Y(n_156)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_93),
.Y(n_157)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_94),
.Y(n_96)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_98),
.Y(n_97)
);

OAI21xp5_ASAP7_75t_L g138 ( 
.A1(n_98),
.A2(n_99),
.B(n_104),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_SL g98 ( 
.A(n_99),
.B(n_104),
.Y(n_98)
);

AND2x2_ASAP7_75t_L g99 ( 
.A(n_100),
.B(n_101),
.Y(n_99)
);

OAI21xp5_ASAP7_75t_SL g251 ( 
.A1(n_100),
.A2(n_119),
.B(n_252),
.Y(n_251)
);

CKINVDCx20_ASAP7_75t_R g102 ( 
.A(n_103),
.Y(n_102)
);

CKINVDCx14_ASAP7_75t_R g105 ( 
.A(n_106),
.Y(n_105)
);

XOR2xp5_ASAP7_75t_L g155 ( 
.A(n_107),
.B(n_156),
.Y(n_155)
);

OAI21xp5_ASAP7_75t_L g107 ( 
.A1(n_108),
.A2(n_123),
.B(n_124),
.Y(n_107)
);

AOI22xp5_ASAP7_75t_L g133 ( 
.A1(n_108),
.A2(n_109),
.B1(n_134),
.B2(n_136),
.Y(n_133)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_109),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_L g109 ( 
.A(n_110),
.B(n_118),
.Y(n_109)
);

CKINVDCx16_ASAP7_75t_R g123 ( 
.A(n_110),
.Y(n_123)
);

AOI22xp5_ASAP7_75t_L g134 ( 
.A1(n_110),
.A2(n_123),
.B1(n_124),
.B2(n_135),
.Y(n_134)
);

AOI22xp5_ASAP7_75t_L g321 ( 
.A1(n_110),
.A2(n_118),
.B1(n_123),
.B2(n_322),
.Y(n_321)
);

AOI21xp5_ASAP7_75t_L g110 ( 
.A1(n_111),
.A2(n_115),
.B(n_116),
.Y(n_110)
);

OAI21xp5_ASAP7_75t_L g183 ( 
.A1(n_111),
.A2(n_145),
.B(n_184),
.Y(n_183)
);

OAI22xp5_ASAP7_75t_SL g198 ( 
.A1(n_111),
.A2(n_189),
.B1(n_199),
.B2(n_200),
.Y(n_198)
);

OAI21xp5_ASAP7_75t_L g227 ( 
.A1(n_111),
.A2(n_116),
.B(n_228),
.Y(n_227)
);

OAI21xp5_ASAP7_75t_L g297 ( 
.A1(n_111),
.A2(n_228),
.B(n_298),
.Y(n_297)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_112),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_SL g143 ( 
.A(n_112),
.B(n_144),
.Y(n_143)
);

AOI22xp5_ASAP7_75t_SL g187 ( 
.A1(n_112),
.A2(n_188),
.B1(n_190),
.B2(n_191),
.Y(n_187)
);

AOI22xp5_ASAP7_75t_L g264 ( 
.A1(n_112),
.A2(n_265),
.B1(n_266),
.B2(n_269),
.Y(n_264)
);

INVx2_ASAP7_75t_L g115 ( 
.A(n_113),
.Y(n_115)
);

INVx5_ASAP7_75t_L g113 ( 
.A(n_114),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_L g206 ( 
.A(n_114),
.B(n_169),
.Y(n_206)
);

INVx8_ASAP7_75t_L g268 ( 
.A(n_114),
.Y(n_268)
);

OAI21xp5_ASAP7_75t_L g246 ( 
.A1(n_115),
.A2(n_143),
.B(n_247),
.Y(n_246)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_117),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_SL g145 ( 
.A(n_117),
.B(n_146),
.Y(n_145)
);

INVxp67_ASAP7_75t_L g322 ( 
.A(n_118),
.Y(n_322)
);

OAI21xp5_ASAP7_75t_SL g118 ( 
.A1(n_119),
.A2(n_120),
.B(n_121),
.Y(n_118)
);

INVxp67_ASAP7_75t_L g121 ( 
.A(n_122),
.Y(n_121)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_124),
.Y(n_135)
);

CKINVDCx16_ASAP7_75t_R g125 ( 
.A(n_126),
.Y(n_125)
);

INVxp67_ASAP7_75t_L g128 ( 
.A(n_129),
.Y(n_128)
);

OAI21xp5_ASAP7_75t_L g130 ( 
.A1(n_131),
.A2(n_158),
.B(n_337),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_L g131 ( 
.A(n_132),
.B(n_155),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_SL g337 ( 
.A(n_132),
.B(n_155),
.Y(n_337)
);

MAJIxp5_ASAP7_75t_L g132 ( 
.A(n_133),
.B(n_137),
.C(n_139),
.Y(n_132)
);

AOI22xp5_ASAP7_75t_L g325 ( 
.A1(n_133),
.A2(n_137),
.B1(n_138),
.B2(n_326),
.Y(n_325)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_133),
.Y(n_326)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_134),
.Y(n_136)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_138),
.Y(n_137)
);

XOR2xp5_ASAP7_75t_L g324 ( 
.A(n_139),
.B(n_325),
.Y(n_324)
);

MAJIxp5_ASAP7_75t_L g139 ( 
.A(n_140),
.B(n_150),
.C(n_154),
.Y(n_139)
);

AOI22xp5_ASAP7_75t_L g318 ( 
.A1(n_140),
.A2(n_141),
.B1(n_319),
.B2(n_320),
.Y(n_318)
);

CKINVDCx14_ASAP7_75t_R g140 ( 
.A(n_141),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_L g141 ( 
.A(n_142),
.B(n_148),
.Y(n_141)
);

XOR2xp5_ASAP7_75t_L g308 ( 
.A(n_142),
.B(n_148),
.Y(n_308)
);

NAND2xp5_ASAP7_75t_L g142 ( 
.A(n_143),
.B(n_145),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_L g228 ( 
.A(n_144),
.B(n_229),
.Y(n_228)
);

INVx2_ASAP7_75t_L g146 ( 
.A(n_147),
.Y(n_146)
);

BUFx2_ASAP7_75t_L g230 ( 
.A(n_147),
.Y(n_230)
);

XNOR2xp5_ASAP7_75t_SL g319 ( 
.A(n_150),
.B(n_154),
.Y(n_319)
);

AOI311xp33_ASAP7_75t_L g158 ( 
.A1(n_159),
.A2(n_315),
.A3(n_327),
.B(n_331),
.C(n_332),
.Y(n_158)
);

NOR3xp33_ASAP7_75t_L g159 ( 
.A(n_160),
.B(n_284),
.C(n_310),
.Y(n_159)
);

AOI21xp5_ASAP7_75t_L g160 ( 
.A1(n_161),
.A2(n_256),
.B(n_283),
.Y(n_160)
);

OAI21xp5_ASAP7_75t_SL g161 ( 
.A1(n_162),
.A2(n_234),
.B(n_255),
.Y(n_161)
);

AOI21xp5_ASAP7_75t_L g162 ( 
.A1(n_163),
.A2(n_210),
.B(n_233),
.Y(n_162)
);

OAI21xp5_ASAP7_75t_SL g163 ( 
.A1(n_164),
.A2(n_185),
.B(n_209),
.Y(n_163)
);

NOR2xp33_ASAP7_75t_L g164 ( 
.A(n_165),
.B(n_175),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_SL g209 ( 
.A(n_165),
.B(n_175),
.Y(n_209)
);

NOR2xp33_ASAP7_75t_SL g165 ( 
.A(n_166),
.B(n_173),
.Y(n_165)
);

AOI22xp5_ASAP7_75t_SL g193 ( 
.A1(n_166),
.A2(n_167),
.B1(n_173),
.B2(n_194),
.Y(n_193)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_167),
.Y(n_166)
);

CKINVDCx16_ASAP7_75t_R g170 ( 
.A(n_171),
.Y(n_170)
);

CKINVDCx20_ASAP7_75t_R g194 ( 
.A(n_173),
.Y(n_194)
);

XNOR2xp5_ASAP7_75t_L g175 ( 
.A(n_176),
.B(n_183),
.Y(n_175)
);

AOI22xp5_ASAP7_75t_L g176 ( 
.A1(n_177),
.A2(n_178),
.B1(n_179),
.B2(n_182),
.Y(n_176)
);

MAJIxp5_ASAP7_75t_L g211 ( 
.A(n_177),
.B(n_182),
.C(n_183),
.Y(n_211)
);

CKINVDCx14_ASAP7_75t_R g177 ( 
.A(n_178),
.Y(n_177)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_179),
.Y(n_182)
);

CKINVDCx20_ASAP7_75t_R g190 ( 
.A(n_184),
.Y(n_190)
);

AOI21xp5_ASAP7_75t_L g185 ( 
.A1(n_186),
.A2(n_195),
.B(n_208),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_L g186 ( 
.A(n_187),
.B(n_193),
.Y(n_186)
);

NOR2xp33_ASAP7_75t_SL g208 ( 
.A(n_187),
.B(n_193),
.Y(n_208)
);

CKINVDCx16_ASAP7_75t_R g188 ( 
.A(n_189),
.Y(n_188)
);

INVx5_ASAP7_75t_L g204 ( 
.A(n_191),
.Y(n_204)
);

INVx5_ASAP7_75t_L g191 ( 
.A(n_192),
.Y(n_191)
);

INVx2_ASAP7_75t_L g201 ( 
.A(n_192),
.Y(n_201)
);

OAI21xp5_ASAP7_75t_SL g195 ( 
.A1(n_196),
.A2(n_202),
.B(n_207),
.Y(n_195)
);

NOR2xp33_ASAP7_75t_L g196 ( 
.A(n_197),
.B(n_198),
.Y(n_196)
);

NAND2xp5_ASAP7_75t_SL g207 ( 
.A(n_197),
.B(n_198),
.Y(n_207)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_201),
.Y(n_200)
);

NAND2xp5_ASAP7_75t_SL g202 ( 
.A(n_203),
.B(n_205),
.Y(n_202)
);

NAND2xp5_ASAP7_75t_L g210 ( 
.A(n_211),
.B(n_212),
.Y(n_210)
);

NOR2xp33_ASAP7_75t_SL g233 ( 
.A(n_211),
.B(n_212),
.Y(n_233)
);

AOI22xp5_ASAP7_75t_SL g212 ( 
.A1(n_213),
.A2(n_224),
.B1(n_231),
.B2(n_232),
.Y(n_212)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_213),
.Y(n_232)
);

AOI22xp5_ASAP7_75t_L g213 ( 
.A1(n_214),
.A2(n_220),
.B1(n_222),
.B2(n_223),
.Y(n_213)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_214),
.Y(n_223)
);

CKINVDCx20_ASAP7_75t_R g216 ( 
.A(n_217),
.Y(n_216)
);

CKINVDCx14_ASAP7_75t_R g240 ( 
.A(n_219),
.Y(n_240)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_220),
.Y(n_222)
);

MAJIxp5_ASAP7_75t_L g235 ( 
.A(n_220),
.B(n_223),
.C(n_231),
.Y(n_235)
);

CKINVDCx20_ASAP7_75t_R g252 ( 
.A(n_221),
.Y(n_252)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_224),
.Y(n_231)
);

XOR2xp5_ASAP7_75t_L g224 ( 
.A(n_225),
.B(n_227),
.Y(n_224)
);

NAND2xp5_ASAP7_75t_L g250 ( 
.A(n_225),
.B(n_227),
.Y(n_250)
);

CKINVDCx20_ASAP7_75t_R g229 ( 
.A(n_230),
.Y(n_229)
);

NOR2xp33_ASAP7_75t_L g234 ( 
.A(n_235),
.B(n_236),
.Y(n_234)
);

NAND2xp5_ASAP7_75t_SL g255 ( 
.A(n_235),
.B(n_236),
.Y(n_255)
);

OAI22xp5_ASAP7_75t_SL g236 ( 
.A1(n_237),
.A2(n_238),
.B1(n_248),
.B2(n_249),
.Y(n_236)
);

MAJIxp5_ASAP7_75t_L g257 ( 
.A(n_237),
.B(n_251),
.C(n_253),
.Y(n_257)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_238),
.Y(n_237)
);

XNOR2xp5_ASAP7_75t_SL g238 ( 
.A(n_239),
.B(n_242),
.Y(n_238)
);

MAJIxp5_ASAP7_75t_L g272 ( 
.A(n_239),
.B(n_244),
.C(n_245),
.Y(n_272)
);

AOI22xp5_ASAP7_75t_L g242 ( 
.A1(n_243),
.A2(n_244),
.B1(n_245),
.B2(n_246),
.Y(n_242)
);

CKINVDCx16_ASAP7_75t_R g243 ( 
.A(n_244),
.Y(n_243)
);

CKINVDCx16_ASAP7_75t_R g245 ( 
.A(n_246),
.Y(n_245)
);

INVxp67_ASAP7_75t_L g265 ( 
.A(n_247),
.Y(n_265)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_249),
.Y(n_248)
);

OAI22xp5_ASAP7_75t_SL g249 ( 
.A1(n_250),
.A2(n_251),
.B1(n_253),
.B2(n_254),
.Y(n_249)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_250),
.Y(n_253)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_251),
.Y(n_254)
);

NAND2xp5_ASAP7_75t_L g256 ( 
.A(n_257),
.B(n_258),
.Y(n_256)
);

NOR2xp33_ASAP7_75t_SL g283 ( 
.A(n_257),
.B(n_258),
.Y(n_283)
);

XOR2xp5_ASAP7_75t_L g258 ( 
.A(n_259),
.B(n_275),
.Y(n_258)
);

OAI22xp5_ASAP7_75t_L g259 ( 
.A1(n_260),
.A2(n_272),
.B1(n_273),
.B2(n_274),
.Y(n_259)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_260),
.Y(n_273)
);

MAJIxp5_ASAP7_75t_L g311 ( 
.A(n_260),
.B(n_274),
.C(n_275),
.Y(n_311)
);

AOI22xp5_ASAP7_75t_L g260 ( 
.A1(n_261),
.A2(n_264),
.B1(n_270),
.B2(n_271),
.Y(n_260)
);

CKINVDCx14_ASAP7_75t_R g271 ( 
.A(n_261),
.Y(n_271)
);

NAND2xp5_ASAP7_75t_L g289 ( 
.A(n_261),
.B(n_270),
.Y(n_289)
);

CKINVDCx20_ASAP7_75t_R g270 ( 
.A(n_264),
.Y(n_270)
);

INVx3_ASAP7_75t_L g266 ( 
.A(n_267),
.Y(n_266)
);

INVx5_ASAP7_75t_L g267 ( 
.A(n_268),
.Y(n_267)
);

INVxp67_ASAP7_75t_L g298 ( 
.A(n_269),
.Y(n_298)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_272),
.Y(n_274)
);

XOR2xp5_ASAP7_75t_L g275 ( 
.A(n_276),
.B(n_280),
.Y(n_275)
);

XOR2xp5_ASAP7_75t_L g276 ( 
.A(n_277),
.B(n_279),
.Y(n_276)
);

MAJIxp5_ASAP7_75t_L g295 ( 
.A(n_277),
.B(n_279),
.C(n_280),
.Y(n_295)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_285),
.Y(n_284)
);

AOI21xp33_ASAP7_75t_L g333 ( 
.A1(n_285),
.A2(n_334),
.B(n_335),
.Y(n_333)
);

NAND2xp5_ASAP7_75t_L g285 ( 
.A(n_286),
.B(n_300),
.Y(n_285)
);

NOR2xp33_ASAP7_75t_SL g335 ( 
.A(n_286),
.B(n_300),
.Y(n_335)
);

MAJIxp5_ASAP7_75t_L g286 ( 
.A(n_287),
.B(n_295),
.C(n_296),
.Y(n_286)
);

OAI22xp5_ASAP7_75t_L g312 ( 
.A1(n_287),
.A2(n_288),
.B1(n_313),
.B2(n_314),
.Y(n_312)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_288),
.Y(n_287)
);

XOR2xp5_ASAP7_75t_L g288 ( 
.A(n_289),
.B(n_290),
.Y(n_288)
);

MAJIxp5_ASAP7_75t_L g309 ( 
.A(n_289),
.B(n_291),
.C(n_292),
.Y(n_309)
);

XOR2xp5_ASAP7_75t_L g290 ( 
.A(n_291),
.B(n_292),
.Y(n_290)
);

INVxp67_ASAP7_75t_L g293 ( 
.A(n_294),
.Y(n_293)
);

XNOR2xp5_ASAP7_75t_SL g314 ( 
.A(n_295),
.B(n_296),
.Y(n_314)
);

XOR2xp5_ASAP7_75t_L g296 ( 
.A(n_297),
.B(n_299),
.Y(n_296)
);

NAND2xp5_ASAP7_75t_L g302 ( 
.A(n_297),
.B(n_299),
.Y(n_302)
);

CKINVDCx5p33_ASAP7_75t_R g329 ( 
.A(n_300),
.Y(n_329)
);

FAx1_ASAP7_75t_SL g300 ( 
.A(n_301),
.B(n_308),
.CI(n_309),
.CON(n_300),
.SN(n_300)
);

OAI22xp5_ASAP7_75t_L g301 ( 
.A1(n_302),
.A2(n_303),
.B1(n_304),
.B2(n_307),
.Y(n_301)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_302),
.Y(n_307)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_304),
.Y(n_303)
);

XNOR2xp5_ASAP7_75t_SL g304 ( 
.A(n_305),
.B(n_306),
.Y(n_304)
);

MAJIxp5_ASAP7_75t_L g323 ( 
.A(n_305),
.B(n_306),
.C(n_307),
.Y(n_323)
);

NOR2xp33_ASAP7_75t_L g310 ( 
.A(n_311),
.B(n_312),
.Y(n_310)
);

AND2x2_ASAP7_75t_L g334 ( 
.A(n_311),
.B(n_312),
.Y(n_334)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_314),
.Y(n_313)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_316),
.Y(n_315)
);

O2A1O1Ixp33_ASAP7_75t_SL g332 ( 
.A1(n_316),
.A2(n_328),
.B(n_333),
.C(n_336),
.Y(n_332)
);

NOR2xp33_ASAP7_75t_L g316 ( 
.A(n_317),
.B(n_324),
.Y(n_316)
);

AND2x2_ASAP7_75t_L g331 ( 
.A(n_317),
.B(n_324),
.Y(n_331)
);

MAJIxp5_ASAP7_75t_L g317 ( 
.A(n_318),
.B(n_321),
.C(n_323),
.Y(n_317)
);

FAx1_ASAP7_75t_L g330 ( 
.A(n_318),
.B(n_321),
.CI(n_323),
.CON(n_330),
.SN(n_330)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_319),
.Y(n_320)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_328),
.Y(n_327)
);

NOR2xp33_ASAP7_75t_L g328 ( 
.A(n_329),
.B(n_330),
.Y(n_328)
);

NAND2xp5_ASAP7_75t_SL g336 ( 
.A(n_329),
.B(n_330),
.Y(n_336)
);

BUFx24_ASAP7_75t_SL g338 ( 
.A(n_330),
.Y(n_338)
);


endmodule