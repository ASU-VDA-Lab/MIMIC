module real_jpeg_8443_n_18 (n_17, n_8, n_0, n_2, n_10, n_9, n_12, n_6, n_11, n_14, n_7, n_3, n_5, n_4, n_299, n_1, n_16, n_15, n_13, n_18);

input n_17;
input n_8;
input n_0;
input n_2;
input n_10;
input n_9;
input n_12;
input n_6;
input n_11;
input n_14;
input n_7;
input n_3;
input n_5;
input n_4;
input n_299;
input n_1;
input n_16;
input n_15;
input n_13;

output n_18;

wire n_108;
wire n_54;
wire n_37;
wire n_233;
wire n_168;
wire n_73;
wire n_35;
wire n_38;
wire n_29;
wire n_91;
wire n_49;
wire n_114;
wire n_201;
wire n_252;
wire n_68;
wire n_260;
wire n_247;
wire n_146;
wire n_83;
wire n_78;
wire n_249;
wire n_166;
wire n_176;
wire n_221;
wire n_215;
wire n_292;
wire n_288;
wire n_286;
wire n_104;
wire n_153;
wire n_194;
wire n_161;
wire n_207;
wire n_280;
wire n_64;
wire n_177;
wire n_291;
wire n_236;
wire n_131;
wire n_47;
wire n_271;
wire n_281;
wire n_163;
wire n_276;
wire n_22;
wire n_287;
wire n_174;
wire n_237;
wire n_87;
wire n_197;
wire n_40;
wire n_173;
wire n_105;
wire n_255;
wire n_115;
wire n_243;
wire n_98;
wire n_27;
wire n_56;
wire n_184;
wire n_48;
wire n_164;
wire n_200;
wire n_293;
wire n_275;
wire n_140;
wire n_227;
wire n_126;
wire n_229;
wire n_214;
wire n_120;
wire n_155;
wire n_113;
wire n_199;
wire n_251;
wire n_93;
wire n_95;
wire n_141;
wire n_242;
wire n_65;
wire n_33;
wire n_139;
wire n_188;
wire n_142;
wire n_175;
wire n_178;
wire n_76;
wire n_67;
wire n_79;
wire n_238;
wire n_235;
wire n_107;
wire n_156;
wire n_282;
wire n_147;
wire n_265;
wire n_189;
wire n_170;
wire n_66;
wire n_231;
wire n_136;
wire n_28;
wire n_44;
wire n_267;
wire n_208;
wire n_62;
wire n_162;
wire n_290;
wire n_239;
wire n_245;
wire n_254;
wire n_250;
wire n_121;
wire n_234;
wire n_106;
wire n_160;
wire n_172;
wire n_211;
wire n_45;
wire n_285;
wire n_112;
wire n_42;
wire n_268;
wire n_145;
wire n_266;
wire n_77;
wire n_109;
wire n_39;
wire n_219;
wire n_122;
wire n_94;
wire n_26;
wire n_19;
wire n_148;
wire n_222;
wire n_262;
wire n_118;
wire n_220;
wire n_294;
wire n_123;
wire n_116;
wire n_246;
wire n_21;
wire n_50;
wire n_143;
wire n_196;
wire n_69;
wire n_186;
wire n_31;
wire n_137;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_218;
wire n_165;
wire n_296;
wire n_134;
wire n_270;
wire n_223;
wire n_72;
wire n_159;
wire n_171;
wire n_151;
wire n_183;
wire n_248;
wire n_272;
wire n_203;
wire n_192;
wire n_100;
wire n_198;
wire n_23;
wire n_51;
wire n_71;
wire n_90;
wire n_61;
wire n_195;
wire n_110;
wire n_205;
wire n_258;
wire n_289;
wire n_117;
wire n_99;
wire n_193;
wire n_261;
wire n_86;
wire n_70;
wire n_41;
wire n_74;
wire n_80;
wire n_32;
wire n_20;
wire n_150;
wire n_228;
wire n_30;
wire n_158;
wire n_204;
wire n_149;
wire n_144;
wire n_130;
wire n_278;
wire n_241;
wire n_103;
wire n_225;
wire n_259;
wire n_232;
wire n_57;
wire n_43;
wire n_157;
wire n_84;
wire n_212;
wire n_82;
wire n_111;
wire n_132;
wire n_284;
wire n_277;
wire n_226;
wire n_185;
wire n_125;
wire n_240;
wire n_55;
wire n_209;
wire n_180;
wire n_58;
wire n_52;
wire n_191;
wire n_63;
wire n_124;
wire n_24;
wire n_92;
wire n_264;
wire n_75;
wire n_97;
wire n_187;
wire n_34;
wire n_190;
wire n_230;
wire n_60;
wire n_263;
wire n_46;
wire n_88;
wire n_279;
wire n_59;
wire n_169;
wire n_167;
wire n_244;
wire n_295;
wire n_179;
wire n_128;
wire n_202;
wire n_133;
wire n_213;
wire n_216;
wire n_138;
wire n_25;
wire n_257;
wire n_217;
wire n_53;
wire n_206;
wire n_127;
wire n_210;
wire n_224;
wire n_119;
wire n_36;
wire n_81;
wire n_102;
wire n_85;
wire n_283;
wire n_181;
wire n_101;
wire n_256;
wire n_274;
wire n_182;
wire n_273;
wire n_96;
wire n_269;
wire n_253;
wire n_89;

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_0),
.Y(n_32)
);

AOI22xp33_ASAP7_75t_SL g50 ( 
.A1(n_1),
.A2(n_31),
.B1(n_32),
.B2(n_51),
.Y(n_50)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_1),
.Y(n_51)
);

AOI22xp33_ASAP7_75t_SL g67 ( 
.A1(n_1),
.A2(n_45),
.B1(n_46),
.B2(n_51),
.Y(n_67)
);

AOI22xp33_ASAP7_75t_SL g109 ( 
.A1(n_1),
.A2(n_51),
.B1(n_57),
.B2(n_58),
.Y(n_109)
);

INVx2_ASAP7_75t_SL g28 ( 
.A(n_2),
.Y(n_28)
);

AOI22xp5_ASAP7_75t_SL g30 ( 
.A1(n_2),
.A2(n_28),
.B1(n_31),
.B2(n_32),
.Y(n_30)
);

AOI21xp33_ASAP7_75t_L g214 ( 
.A1(n_2),
.A2(n_11),
.B(n_32),
.Y(n_214)
);

AOI22xp33_ASAP7_75t_SL g33 ( 
.A1(n_3),
.A2(n_27),
.B1(n_34),
.B2(n_35),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_3),
.Y(n_35)
);

AOI22xp33_ASAP7_75t_SL g118 ( 
.A1(n_3),
.A2(n_31),
.B1(n_32),
.B2(n_35),
.Y(n_118)
);

OAI22xp5_ASAP7_75t_SL g183 ( 
.A1(n_3),
.A2(n_35),
.B1(n_57),
.B2(n_58),
.Y(n_183)
);

OAI22xp5_ASAP7_75t_SL g228 ( 
.A1(n_3),
.A2(n_35),
.B1(n_45),
.B2(n_46),
.Y(n_228)
);

BUFx10_ASAP7_75t_L g74 ( 
.A(n_4),
.Y(n_74)
);

BUFx12f_ASAP7_75t_L g58 ( 
.A(n_5),
.Y(n_58)
);

A2O1A1Ixp33_ASAP7_75t_SL g54 ( 
.A1(n_6),
.A2(n_45),
.B(n_55),
.C(n_56),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_6),
.B(n_45),
.Y(n_55)
);

AOI22xp5_ASAP7_75t_SL g56 ( 
.A1(n_6),
.A2(n_57),
.B1(n_58),
.B2(n_59),
.Y(n_56)
);

INVx3_ASAP7_75t_L g59 ( 
.A(n_6),
.Y(n_59)
);

BUFx6f_ASAP7_75t_SL g42 ( 
.A(n_7),
.Y(n_42)
);

BUFx3_ASAP7_75t_L g46 ( 
.A(n_8),
.Y(n_46)
);

AOI22xp5_ASAP7_75t_SL g60 ( 
.A1(n_9),
.A2(n_45),
.B1(n_46),
.B2(n_61),
.Y(n_60)
);

CKINVDCx20_ASAP7_75t_R g61 ( 
.A(n_9),
.Y(n_61)
);

AOI22xp33_ASAP7_75t_L g76 ( 
.A1(n_9),
.A2(n_57),
.B1(n_58),
.B2(n_61),
.Y(n_76)
);

AOI22xp33_ASAP7_75t_SL g92 ( 
.A1(n_9),
.A2(n_31),
.B1(n_32),
.B2(n_61),
.Y(n_92)
);

AOI22xp33_ASAP7_75t_SL g36 ( 
.A1(n_10),
.A2(n_27),
.B1(n_34),
.B2(n_37),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_10),
.Y(n_37)
);

AOI22xp33_ASAP7_75t_SL g65 ( 
.A1(n_10),
.A2(n_31),
.B1(n_32),
.B2(n_37),
.Y(n_65)
);

AOI22xp33_ASAP7_75t_SL g111 ( 
.A1(n_10),
.A2(n_37),
.B1(n_45),
.B2(n_46),
.Y(n_111)
);

OAI22xp5_ASAP7_75t_L g197 ( 
.A1(n_10),
.A2(n_37),
.B1(n_57),
.B2(n_58),
.Y(n_197)
);

AOI21xp5_ASAP7_75t_L g137 ( 
.A1(n_11),
.A2(n_45),
.B(n_138),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_L g138 ( 
.A(n_11),
.B(n_45),
.Y(n_138)
);

CKINVDCx20_ASAP7_75t_R g151 ( 
.A(n_11),
.Y(n_151)
);

OAI22xp5_ASAP7_75t_L g153 ( 
.A1(n_11),
.A2(n_72),
.B1(n_75),
.B2(n_149),
.Y(n_153)
);

AOI21xp5_ASAP7_75t_L g173 ( 
.A1(n_11),
.A2(n_31),
.B(n_174),
.Y(n_173)
);

NOR2xp33_ASAP7_75t_L g174 ( 
.A(n_11),
.B(n_31),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_L g194 ( 
.A(n_11),
.B(n_195),
.Y(n_194)
);

OAI22xp33_ASAP7_75t_SL g235 ( 
.A1(n_11),
.A2(n_27),
.B1(n_34),
.B2(n_151),
.Y(n_235)
);

AOI22xp33_ASAP7_75t_SL g139 ( 
.A1(n_12),
.A2(n_45),
.B1(n_46),
.B2(n_140),
.Y(n_139)
);

CKINVDCx20_ASAP7_75t_R g140 ( 
.A(n_12),
.Y(n_140)
);

AOI22xp33_ASAP7_75t_SL g149 ( 
.A1(n_12),
.A2(n_57),
.B1(n_58),
.B2(n_140),
.Y(n_149)
);

AOI22xp5_ASAP7_75t_L g175 ( 
.A1(n_12),
.A2(n_31),
.B1(n_32),
.B2(n_140),
.Y(n_175)
);

OAI22xp5_ASAP7_75t_SL g236 ( 
.A1(n_12),
.A2(n_27),
.B1(n_34),
.B2(n_140),
.Y(n_236)
);

BUFx2_ASAP7_75t_L g27 ( 
.A(n_13),
.Y(n_27)
);

AOI22xp33_ASAP7_75t_SL g48 ( 
.A1(n_14),
.A2(n_31),
.B1(n_32),
.B2(n_49),
.Y(n_48)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_14),
.Y(n_49)
);

AOI22xp33_ASAP7_75t_L g78 ( 
.A1(n_14),
.A2(n_45),
.B1(n_46),
.B2(n_49),
.Y(n_78)
);

AOI22xp33_ASAP7_75t_SL g88 ( 
.A1(n_14),
.A2(n_27),
.B1(n_34),
.B2(n_49),
.Y(n_88)
);

AOI22xp33_ASAP7_75t_SL g218 ( 
.A1(n_14),
.A2(n_49),
.B1(n_57),
.B2(n_58),
.Y(n_218)
);

AOI22xp33_ASAP7_75t_SL g114 ( 
.A1(n_15),
.A2(n_27),
.B1(n_34),
.B2(n_115),
.Y(n_114)
);

CKINVDCx20_ASAP7_75t_R g115 ( 
.A(n_15),
.Y(n_115)
);

AOI22xp33_ASAP7_75t_SL g133 ( 
.A1(n_15),
.A2(n_57),
.B1(n_58),
.B2(n_115),
.Y(n_133)
);

AOI22xp33_ASAP7_75t_L g171 ( 
.A1(n_15),
.A2(n_45),
.B1(n_46),
.B2(n_115),
.Y(n_171)
);

AOI22xp33_ASAP7_75t_SL g232 ( 
.A1(n_15),
.A2(n_31),
.B1(n_32),
.B2(n_115),
.Y(n_232)
);

AOI22xp33_ASAP7_75t_SL g81 ( 
.A1(n_16),
.A2(n_27),
.B1(n_34),
.B2(n_82),
.Y(n_81)
);

CKINVDCx20_ASAP7_75t_R g82 ( 
.A(n_16),
.Y(n_82)
);

AOI22xp33_ASAP7_75t_SL g166 ( 
.A1(n_16),
.A2(n_57),
.B1(n_58),
.B2(n_82),
.Y(n_166)
);

AOI22xp33_ASAP7_75t_SL g203 ( 
.A1(n_16),
.A2(n_45),
.B1(n_46),
.B2(n_82),
.Y(n_203)
);

AOI22xp33_ASAP7_75t_SL g244 ( 
.A1(n_16),
.A2(n_31),
.B1(n_32),
.B2(n_82),
.Y(n_244)
);

AOI22xp33_ASAP7_75t_SL g130 ( 
.A1(n_17),
.A2(n_57),
.B1(n_58),
.B2(n_131),
.Y(n_130)
);

CKINVDCx20_ASAP7_75t_R g131 ( 
.A(n_17),
.Y(n_131)
);

AOI22xp33_ASAP7_75t_SL g164 ( 
.A1(n_17),
.A2(n_45),
.B1(n_46),
.B2(n_131),
.Y(n_164)
);

AOI22xp33_ASAP7_75t_SL g191 ( 
.A1(n_17),
.A2(n_31),
.B1(n_32),
.B2(n_131),
.Y(n_191)
);

AOI22xp33_ASAP7_75t_SL g248 ( 
.A1(n_17),
.A2(n_27),
.B1(n_34),
.B2(n_131),
.Y(n_248)
);

XOR2xp5_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_97),
.Y(n_18)
);

NAND2xp5_ASAP7_75t_SL g19 ( 
.A(n_20),
.B(n_96),
.Y(n_19)
);

INVxp67_ASAP7_75t_L g20 ( 
.A(n_21),
.Y(n_20)
);

NOR2xp33_ASAP7_75t_L g21 ( 
.A(n_22),
.B(n_83),
.Y(n_21)
);

NAND2xp5_ASAP7_75t_L g96 ( 
.A(n_22),
.B(n_83),
.Y(n_96)
);

MAJIxp5_ASAP7_75t_L g22 ( 
.A(n_23),
.B(n_63),
.C(n_68),
.Y(n_22)
);

FAx1_ASAP7_75t_SL g119 ( 
.A(n_23),
.B(n_63),
.CI(n_68),
.CON(n_119),
.SN(n_119)
);

AOI22xp5_ASAP7_75t_L g23 ( 
.A1(n_24),
.A2(n_25),
.B1(n_38),
.B2(n_39),
.Y(n_23)
);

OAI22xp5_ASAP7_75t_SL g84 ( 
.A1(n_24),
.A2(n_25),
.B1(n_85),
.B2(n_86),
.Y(n_84)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_25),
.Y(n_24)
);

MAJIxp5_ASAP7_75t_L g95 ( 
.A(n_25),
.B(n_52),
.C(n_62),
.Y(n_95)
);

OAI22xp5_ASAP7_75t_SL g25 ( 
.A1(n_26),
.A2(n_30),
.B1(n_33),
.B2(n_36),
.Y(n_25)
);

OAI22xp5_ASAP7_75t_SL g80 ( 
.A1(n_26),
.A2(n_30),
.B1(n_33),
.B2(n_81),
.Y(n_80)
);

OAI22xp5_ASAP7_75t_SL g87 ( 
.A1(n_26),
.A2(n_30),
.B1(n_36),
.B2(n_88),
.Y(n_87)
);

OAI22xp5_ASAP7_75t_SL g113 ( 
.A1(n_26),
.A2(n_30),
.B1(n_81),
.B2(n_114),
.Y(n_113)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_26),
.Y(n_234)
);

OAI22xp5_ASAP7_75t_SL g246 ( 
.A1(n_26),
.A2(n_30),
.B1(n_247),
.B2(n_248),
.Y(n_246)
);

OAI22xp5_ASAP7_75t_SL g265 ( 
.A1(n_26),
.A2(n_30),
.B1(n_114),
.B2(n_248),
.Y(n_265)
);

A2O1A1Ixp33_ASAP7_75t_L g26 ( 
.A1(n_27),
.A2(n_28),
.B(n_29),
.C(n_30),
.Y(n_26)
);

NOR2xp33_ASAP7_75t_L g29 ( 
.A(n_27),
.B(n_28),
.Y(n_29)
);

INVx3_ASAP7_75t_L g34 ( 
.A(n_27),
.Y(n_34)
);

A2O1A1Ixp33_ASAP7_75t_L g213 ( 
.A1(n_27),
.A2(n_28),
.B(n_151),
.C(n_214),
.Y(n_213)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_30),
.Y(n_195)
);

A2O1A1Ixp33_ASAP7_75t_L g41 ( 
.A1(n_31),
.A2(n_42),
.B(n_43),
.C(n_44),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g43 ( 
.A(n_31),
.B(n_42),
.Y(n_43)
);

INVx11_ASAP7_75t_L g31 ( 
.A(n_32),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_39),
.Y(n_38)
);

OAI22xp5_ASAP7_75t_L g39 ( 
.A1(n_40),
.A2(n_52),
.B1(n_53),
.B2(n_62),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g62 ( 
.A(n_40),
.Y(n_62)
);

OAI22xp5_ASAP7_75t_SL g40 ( 
.A1(n_41),
.A2(n_44),
.B1(n_48),
.B2(n_50),
.Y(n_40)
);

OAI22xp5_ASAP7_75t_SL g64 ( 
.A1(n_41),
.A2(n_44),
.B1(n_48),
.B2(n_65),
.Y(n_64)
);

OAI22xp5_ASAP7_75t_SL g91 ( 
.A1(n_41),
.A2(n_44),
.B1(n_50),
.B2(n_92),
.Y(n_91)
);

OAI22xp5_ASAP7_75t_SL g117 ( 
.A1(n_41),
.A2(n_44),
.B1(n_65),
.B2(n_118),
.Y(n_117)
);

OAI22xp5_ASAP7_75t_L g172 ( 
.A1(n_41),
.A2(n_44),
.B1(n_173),
.B2(n_175),
.Y(n_172)
);

OAI22xp5_ASAP7_75t_SL g190 ( 
.A1(n_41),
.A2(n_44),
.B1(n_175),
.B2(n_191),
.Y(n_190)
);

OAI22xp5_ASAP7_75t_L g231 ( 
.A1(n_41),
.A2(n_44),
.B1(n_191),
.B2(n_232),
.Y(n_231)
);

OAI22xp5_ASAP7_75t_SL g243 ( 
.A1(n_41),
.A2(n_44),
.B1(n_232),
.B2(n_244),
.Y(n_243)
);

OAI22xp5_ASAP7_75t_SL g263 ( 
.A1(n_41),
.A2(n_44),
.B1(n_118),
.B2(n_244),
.Y(n_263)
);

AOI22xp5_ASAP7_75t_SL g44 ( 
.A1(n_42),
.A2(n_45),
.B1(n_46),
.B2(n_47),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_42),
.Y(n_47)
);

INVxp67_ASAP7_75t_L g180 ( 
.A(n_43),
.Y(n_180)
);

NOR2xp33_ASAP7_75t_L g162 ( 
.A(n_44),
.B(n_151),
.Y(n_162)
);

NOR2xp33_ASAP7_75t_SL g179 ( 
.A(n_45),
.B(n_47),
.Y(n_179)
);

INVx4_ASAP7_75t_L g45 ( 
.A(n_46),
.Y(n_45)
);

OAI22xp5_ASAP7_75t_L g177 ( 
.A1(n_46),
.A2(n_178),
.B1(n_179),
.B2(n_180),
.Y(n_177)
);

OAI22xp5_ASAP7_75t_L g90 ( 
.A1(n_52),
.A2(n_53),
.B1(n_91),
.B2(n_93),
.Y(n_90)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_53),
.Y(n_52)
);

AOI21xp5_ASAP7_75t_SL g53 ( 
.A1(n_54),
.A2(n_56),
.B(n_60),
.Y(n_53)
);

OAI22xp5_ASAP7_75t_SL g66 ( 
.A1(n_54),
.A2(n_56),
.B1(n_60),
.B2(n_67),
.Y(n_66)
);

OAI22xp5_ASAP7_75t_SL g77 ( 
.A1(n_54),
.A2(n_56),
.B1(n_67),
.B2(n_78),
.Y(n_77)
);

OAI22xp5_ASAP7_75t_L g110 ( 
.A1(n_54),
.A2(n_56),
.B1(n_78),
.B2(n_111),
.Y(n_110)
);

OAI22xp5_ASAP7_75t_L g136 ( 
.A1(n_54),
.A2(n_56),
.B1(n_137),
.B2(n_139),
.Y(n_136)
);

OAI22xp5_ASAP7_75t_SL g163 ( 
.A1(n_54),
.A2(n_56),
.B1(n_139),
.B2(n_164),
.Y(n_163)
);

OAI22xp5_ASAP7_75t_L g170 ( 
.A1(n_54),
.A2(n_56),
.B1(n_164),
.B2(n_171),
.Y(n_170)
);

OAI22xp5_ASAP7_75t_SL g202 ( 
.A1(n_54),
.A2(n_56),
.B1(n_171),
.B2(n_203),
.Y(n_202)
);

INVxp67_ASAP7_75t_L g227 ( 
.A(n_54),
.Y(n_227)
);

OAI22xp5_ASAP7_75t_L g253 ( 
.A1(n_54),
.A2(n_56),
.B1(n_111),
.B2(n_254),
.Y(n_253)
);

INVxp67_ASAP7_75t_L g144 ( 
.A(n_55),
.Y(n_144)
);

NOR2xp33_ASAP7_75t_SL g150 ( 
.A(n_56),
.B(n_151),
.Y(n_150)
);

CKINVDCx20_ASAP7_75t_R g229 ( 
.A(n_56),
.Y(n_229)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_57),
.B(n_74),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_SL g142 ( 
.A(n_57),
.B(n_59),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_SL g154 ( 
.A(n_57),
.B(n_155),
.Y(n_154)
);

CKINVDCx20_ASAP7_75t_R g57 ( 
.A(n_58),
.Y(n_57)
);

OAI22xp5_ASAP7_75t_L g141 ( 
.A1(n_58),
.A2(n_142),
.B1(n_143),
.B2(n_144),
.Y(n_141)
);

AOI21xp5_ASAP7_75t_L g104 ( 
.A1(n_63),
.A2(n_64),
.B(n_66),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_64),
.B(n_66),
.Y(n_63)
);

OAI21xp5_ASAP7_75t_L g68 ( 
.A1(n_69),
.A2(n_79),
.B(n_80),
.Y(n_68)
);

AOI22xp5_ASAP7_75t_L g100 ( 
.A1(n_69),
.A2(n_70),
.B1(n_101),
.B2(n_102),
.Y(n_100)
);

CKINVDCx20_ASAP7_75t_R g69 ( 
.A(n_70),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_L g70 ( 
.A(n_71),
.B(n_77),
.Y(n_70)
);

CKINVDCx20_ASAP7_75t_R g79 ( 
.A(n_71),
.Y(n_79)
);

OAI22xp5_ASAP7_75t_L g102 ( 
.A1(n_71),
.A2(n_79),
.B1(n_80),
.B2(n_103),
.Y(n_102)
);

OAI22xp5_ASAP7_75t_L g278 ( 
.A1(n_71),
.A2(n_77),
.B1(n_79),
.B2(n_279),
.Y(n_278)
);

AOI21xp5_ASAP7_75t_L g71 ( 
.A1(n_72),
.A2(n_75),
.B(n_76),
.Y(n_71)
);

OAI22xp5_ASAP7_75t_L g108 ( 
.A1(n_72),
.A2(n_75),
.B1(n_76),
.B2(n_109),
.Y(n_108)
);

OAI22xp5_ASAP7_75t_SL g148 ( 
.A1(n_72),
.A2(n_75),
.B1(n_130),
.B2(n_149),
.Y(n_148)
);

OAI22xp5_ASAP7_75t_L g165 ( 
.A1(n_72),
.A2(n_75),
.B1(n_133),
.B2(n_166),
.Y(n_165)
);

OAI22xp5_ASAP7_75t_L g181 ( 
.A1(n_72),
.A2(n_75),
.B1(n_166),
.B2(n_182),
.Y(n_181)
);

OAI22xp5_ASAP7_75t_SL g216 ( 
.A1(n_72),
.A2(n_75),
.B1(n_217),
.B2(n_218),
.Y(n_216)
);

OAI22xp5_ASAP7_75t_L g252 ( 
.A1(n_72),
.A2(n_75),
.B1(n_109),
.B2(n_218),
.Y(n_252)
);

CKINVDCx16_ASAP7_75t_R g72 ( 
.A(n_73),
.Y(n_72)
);

AOI22xp5_ASAP7_75t_SL g128 ( 
.A1(n_73),
.A2(n_74),
.B1(n_129),
.B2(n_132),
.Y(n_128)
);

AOI22xp5_ASAP7_75t_L g196 ( 
.A1(n_73),
.A2(n_74),
.B1(n_183),
.B2(n_197),
.Y(n_196)
);

CKINVDCx16_ASAP7_75t_R g75 ( 
.A(n_74),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g155 ( 
.A(n_75),
.B(n_151),
.Y(n_155)
);

CKINVDCx20_ASAP7_75t_R g279 ( 
.A(n_77),
.Y(n_279)
);

CKINVDCx20_ASAP7_75t_R g103 ( 
.A(n_80),
.Y(n_103)
);

XOR2xp5_ASAP7_75t_L g83 ( 
.A(n_84),
.B(n_95),
.Y(n_83)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_86),
.Y(n_85)
);

AOI22xp5_ASAP7_75t_L g86 ( 
.A1(n_87),
.A2(n_89),
.B1(n_90),
.B2(n_94),
.Y(n_86)
);

CKINVDCx20_ASAP7_75t_R g94 ( 
.A(n_87),
.Y(n_94)
);

CKINVDCx20_ASAP7_75t_R g89 ( 
.A(n_90),
.Y(n_89)
);

CKINVDCx20_ASAP7_75t_R g93 ( 
.A(n_91),
.Y(n_93)
);

OAI21xp5_ASAP7_75t_L g97 ( 
.A1(n_98),
.A2(n_120),
.B(n_296),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_99),
.B(n_119),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_SL g296 ( 
.A(n_99),
.B(n_119),
.Y(n_296)
);

MAJIxp5_ASAP7_75t_L g99 ( 
.A(n_100),
.B(n_104),
.C(n_105),
.Y(n_99)
);

XOR2xp5_ASAP7_75t_L g283 ( 
.A(n_100),
.B(n_104),
.Y(n_283)
);

CKINVDCx20_ASAP7_75t_R g101 ( 
.A(n_102),
.Y(n_101)
);

AOI22xp5_ASAP7_75t_SL g281 ( 
.A1(n_105),
.A2(n_106),
.B1(n_282),
.B2(n_283),
.Y(n_281)
);

CKINVDCx20_ASAP7_75t_R g105 ( 
.A(n_106),
.Y(n_105)
);

MAJIxp5_ASAP7_75t_L g106 ( 
.A(n_107),
.B(n_112),
.C(n_116),
.Y(n_106)
);

XOR2xp5_ASAP7_75t_L g276 ( 
.A(n_107),
.B(n_277),
.Y(n_276)
);

NAND2xp5_ASAP7_75t_L g107 ( 
.A(n_108),
.B(n_110),
.Y(n_107)
);

XNOR2xp5_ASAP7_75t_L g259 ( 
.A(n_108),
.B(n_110),
.Y(n_259)
);

OAI22xp5_ASAP7_75t_SL g277 ( 
.A1(n_112),
.A2(n_113),
.B1(n_116),
.B2(n_117),
.Y(n_277)
);

CKINVDCx20_ASAP7_75t_R g112 ( 
.A(n_113),
.Y(n_112)
);

CKINVDCx20_ASAP7_75t_R g116 ( 
.A(n_117),
.Y(n_116)
);

BUFx24_ASAP7_75t_SL g298 ( 
.A(n_119),
.Y(n_298)
);

AOI321xp33_ASAP7_75t_L g120 ( 
.A1(n_121),
.A2(n_273),
.A3(n_284),
.B1(n_290),
.B2(n_295),
.C(n_299),
.Y(n_120)
);

NOR3xp33_ASAP7_75t_L g121 ( 
.A(n_122),
.B(n_238),
.C(n_269),
.Y(n_121)
);

AOI21xp5_ASAP7_75t_L g122 ( 
.A1(n_123),
.A2(n_207),
.B(n_237),
.Y(n_122)
);

OAI21xp5_ASAP7_75t_SL g123 ( 
.A1(n_124),
.A2(n_185),
.B(n_206),
.Y(n_123)
);

AOI21xp5_ASAP7_75t_L g124 ( 
.A1(n_125),
.A2(n_168),
.B(n_184),
.Y(n_124)
);

OAI21xp5_ASAP7_75t_SL g125 ( 
.A1(n_126),
.A2(n_158),
.B(n_167),
.Y(n_125)
);

AOI21xp5_ASAP7_75t_L g126 ( 
.A1(n_127),
.A2(n_146),
.B(n_157),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_128),
.B(n_134),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_SL g157 ( 
.A(n_128),
.B(n_134),
.Y(n_157)
);

CKINVDCx20_ASAP7_75t_R g129 ( 
.A(n_130),
.Y(n_129)
);

CKINVDCx20_ASAP7_75t_R g132 ( 
.A(n_133),
.Y(n_132)
);

AOI22xp5_ASAP7_75t_SL g134 ( 
.A1(n_135),
.A2(n_136),
.B1(n_141),
.B2(n_145),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_SL g159 ( 
.A(n_135),
.B(n_145),
.Y(n_159)
);

CKINVDCx20_ASAP7_75t_R g135 ( 
.A(n_136),
.Y(n_135)
);

CKINVDCx20_ASAP7_75t_R g143 ( 
.A(n_138),
.Y(n_143)
);

CKINVDCx20_ASAP7_75t_R g145 ( 
.A(n_141),
.Y(n_145)
);

OAI21xp5_ASAP7_75t_SL g146 ( 
.A1(n_147),
.A2(n_152),
.B(n_156),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_L g147 ( 
.A(n_148),
.B(n_150),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_L g156 ( 
.A(n_148),
.B(n_150),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_SL g152 ( 
.A(n_153),
.B(n_154),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_L g158 ( 
.A(n_159),
.B(n_160),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_SL g167 ( 
.A(n_159),
.B(n_160),
.Y(n_167)
);

CKINVDCx5p33_ASAP7_75t_R g160 ( 
.A(n_161),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_L g168 ( 
.A(n_161),
.B(n_169),
.Y(n_168)
);

NOR2xp33_ASAP7_75t_SL g184 ( 
.A(n_161),
.B(n_169),
.Y(n_184)
);

FAx1_ASAP7_75t_SL g161 ( 
.A(n_162),
.B(n_163),
.CI(n_165),
.CON(n_161),
.SN(n_161)
);

CKINVDCx5p33_ASAP7_75t_R g186 ( 
.A(n_169),
.Y(n_186)
);

FAx1_ASAP7_75t_SL g169 ( 
.A(n_170),
.B(n_172),
.CI(n_176),
.CON(n_169),
.SN(n_169)
);

CKINVDCx16_ASAP7_75t_R g178 ( 
.A(n_174),
.Y(n_178)
);

XOR2xp5_ASAP7_75t_L g176 ( 
.A(n_177),
.B(n_181),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_L g201 ( 
.A(n_177),
.B(n_181),
.Y(n_201)
);

CKINVDCx20_ASAP7_75t_R g182 ( 
.A(n_183),
.Y(n_182)
);

NOR2xp33_ASAP7_75t_L g185 ( 
.A(n_186),
.B(n_187),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_SL g206 ( 
.A(n_186),
.B(n_187),
.Y(n_206)
);

OAI22xp5_ASAP7_75t_SL g187 ( 
.A1(n_188),
.A2(n_189),
.B1(n_199),
.B2(n_200),
.Y(n_187)
);

MAJIxp5_ASAP7_75t_L g208 ( 
.A(n_188),
.B(n_202),
.C(n_204),
.Y(n_208)
);

CKINVDCx16_ASAP7_75t_R g188 ( 
.A(n_189),
.Y(n_188)
);

AOI22xp5_ASAP7_75t_L g189 ( 
.A1(n_190),
.A2(n_192),
.B1(n_193),
.B2(n_198),
.Y(n_189)
);

CKINVDCx20_ASAP7_75t_R g198 ( 
.A(n_190),
.Y(n_198)
);

CKINVDCx20_ASAP7_75t_R g192 ( 
.A(n_193),
.Y(n_192)
);

XOR2xp5_ASAP7_75t_L g193 ( 
.A(n_194),
.B(n_196),
.Y(n_193)
);

MAJIxp5_ASAP7_75t_L g219 ( 
.A(n_194),
.B(n_196),
.C(n_198),
.Y(n_219)
);

AOI22xp5_ASAP7_75t_SL g233 ( 
.A1(n_195),
.A2(n_234),
.B1(n_235),
.B2(n_236),
.Y(n_233)
);

CKINVDCx20_ASAP7_75t_R g217 ( 
.A(n_197),
.Y(n_217)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_200),
.Y(n_199)
);

OAI22xp5_ASAP7_75t_SL g200 ( 
.A1(n_201),
.A2(n_202),
.B1(n_204),
.B2(n_205),
.Y(n_200)
);

CKINVDCx20_ASAP7_75t_R g204 ( 
.A(n_201),
.Y(n_204)
);

CKINVDCx20_ASAP7_75t_R g205 ( 
.A(n_202),
.Y(n_205)
);

CKINVDCx20_ASAP7_75t_R g226 ( 
.A(n_203),
.Y(n_226)
);

NAND2xp5_ASAP7_75t_L g207 ( 
.A(n_208),
.B(n_209),
.Y(n_207)
);

NOR2xp33_ASAP7_75t_SL g237 ( 
.A(n_208),
.B(n_209),
.Y(n_237)
);

XOR2xp5_ASAP7_75t_L g209 ( 
.A(n_210),
.B(n_222),
.Y(n_209)
);

OAI22xp5_ASAP7_75t_L g210 ( 
.A1(n_211),
.A2(n_219),
.B1(n_220),
.B2(n_221),
.Y(n_210)
);

CKINVDCx20_ASAP7_75t_R g220 ( 
.A(n_211),
.Y(n_220)
);

MAJIxp5_ASAP7_75t_L g270 ( 
.A(n_211),
.B(n_221),
.C(n_222),
.Y(n_270)
);

AOI22xp5_ASAP7_75t_L g211 ( 
.A1(n_212),
.A2(n_213),
.B1(n_215),
.B2(n_216),
.Y(n_211)
);

NAND2xp5_ASAP7_75t_L g250 ( 
.A(n_212),
.B(n_216),
.Y(n_250)
);

CKINVDCx20_ASAP7_75t_R g212 ( 
.A(n_213),
.Y(n_212)
);

CKINVDCx20_ASAP7_75t_R g215 ( 
.A(n_216),
.Y(n_215)
);

CKINVDCx20_ASAP7_75t_R g221 ( 
.A(n_219),
.Y(n_221)
);

XOR2xp5_ASAP7_75t_L g222 ( 
.A(n_223),
.B(n_233),
.Y(n_222)
);

OAI22xp5_ASAP7_75t_L g223 ( 
.A1(n_224),
.A2(n_225),
.B1(n_230),
.B2(n_231),
.Y(n_223)
);

CKINVDCx20_ASAP7_75t_R g224 ( 
.A(n_225),
.Y(n_224)
);

MAJIxp5_ASAP7_75t_L g255 ( 
.A(n_225),
.B(n_230),
.C(n_233),
.Y(n_255)
);

AOI22xp5_ASAP7_75t_L g225 ( 
.A1(n_226),
.A2(n_227),
.B1(n_228),
.B2(n_229),
.Y(n_225)
);

CKINVDCx20_ASAP7_75t_R g254 ( 
.A(n_228),
.Y(n_254)
);

CKINVDCx20_ASAP7_75t_R g230 ( 
.A(n_231),
.Y(n_230)
);

CKINVDCx20_ASAP7_75t_R g247 ( 
.A(n_236),
.Y(n_247)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_239),
.Y(n_238)
);

AOI21xp33_ASAP7_75t_L g291 ( 
.A1(n_239),
.A2(n_292),
.B(n_293),
.Y(n_291)
);

NAND2xp5_ASAP7_75t_L g239 ( 
.A(n_240),
.B(n_256),
.Y(n_239)
);

NOR2xp33_ASAP7_75t_SL g293 ( 
.A(n_240),
.B(n_256),
.Y(n_293)
);

MAJIxp5_ASAP7_75t_L g240 ( 
.A(n_241),
.B(n_251),
.C(n_255),
.Y(n_240)
);

XNOR2xp5_ASAP7_75t_L g271 ( 
.A(n_241),
.B(n_272),
.Y(n_271)
);

XNOR2xp5_ASAP7_75t_SL g241 ( 
.A(n_242),
.B(n_250),
.Y(n_241)
);

OAI22xp5_ASAP7_75t_SL g242 ( 
.A1(n_243),
.A2(n_245),
.B1(n_246),
.B2(n_249),
.Y(n_242)
);

CKINVDCx20_ASAP7_75t_R g249 ( 
.A(n_243),
.Y(n_249)
);

MAJIxp5_ASAP7_75t_SL g267 ( 
.A(n_245),
.B(n_249),
.C(n_250),
.Y(n_267)
);

CKINVDCx20_ASAP7_75t_R g245 ( 
.A(n_246),
.Y(n_245)
);

XNOR2xp5_ASAP7_75t_L g272 ( 
.A(n_251),
.B(n_255),
.Y(n_272)
);

XOR2xp5_ASAP7_75t_L g251 ( 
.A(n_252),
.B(n_253),
.Y(n_251)
);

NAND2xp5_ASAP7_75t_L g261 ( 
.A(n_252),
.B(n_253),
.Y(n_261)
);

AOI22xp5_ASAP7_75t_SL g256 ( 
.A1(n_257),
.A2(n_258),
.B1(n_267),
.B2(n_268),
.Y(n_256)
);

CKINVDCx16_ASAP7_75t_R g257 ( 
.A(n_258),
.Y(n_257)
);

XOR2xp5_ASAP7_75t_L g258 ( 
.A(n_259),
.B(n_260),
.Y(n_258)
);

MAJIxp5_ASAP7_75t_L g286 ( 
.A(n_259),
.B(n_260),
.C(n_268),
.Y(n_286)
);

XOR2xp5_ASAP7_75t_L g260 ( 
.A(n_261),
.B(n_262),
.Y(n_260)
);

MAJIxp5_ASAP7_75t_L g280 ( 
.A(n_261),
.B(n_264),
.C(n_266),
.Y(n_280)
);

OAI22xp5_ASAP7_75t_SL g262 ( 
.A1(n_263),
.A2(n_264),
.B1(n_265),
.B2(n_266),
.Y(n_262)
);

CKINVDCx20_ASAP7_75t_R g266 ( 
.A(n_263),
.Y(n_266)
);

CKINVDCx20_ASAP7_75t_R g264 ( 
.A(n_265),
.Y(n_264)
);

CKINVDCx20_ASAP7_75t_R g268 ( 
.A(n_267),
.Y(n_268)
);

NOR2xp33_ASAP7_75t_L g269 ( 
.A(n_270),
.B(n_271),
.Y(n_269)
);

AND2x2_ASAP7_75t_L g292 ( 
.A(n_270),
.B(n_271),
.Y(n_292)
);

NAND2xp5_ASAP7_75t_L g273 ( 
.A(n_274),
.B(n_281),
.Y(n_273)
);

NOR2xp33_ASAP7_75t_SL g295 ( 
.A(n_274),
.B(n_281),
.Y(n_295)
);

MAJIxp5_ASAP7_75t_L g274 ( 
.A(n_275),
.B(n_278),
.C(n_280),
.Y(n_274)
);

AOI22xp5_ASAP7_75t_L g288 ( 
.A1(n_275),
.A2(n_276),
.B1(n_278),
.B2(n_289),
.Y(n_288)
);

CKINVDCx20_ASAP7_75t_R g275 ( 
.A(n_276),
.Y(n_275)
);

CKINVDCx20_ASAP7_75t_R g289 ( 
.A(n_278),
.Y(n_289)
);

XNOR2xp5_ASAP7_75t_L g287 ( 
.A(n_280),
.B(n_288),
.Y(n_287)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_283),
.Y(n_282)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_285),
.Y(n_284)
);

OAI21xp5_ASAP7_75t_L g290 ( 
.A1(n_285),
.A2(n_291),
.B(n_294),
.Y(n_290)
);

NOR2xp33_ASAP7_75t_L g285 ( 
.A(n_286),
.B(n_287),
.Y(n_285)
);

NAND2xp5_ASAP7_75t_SL g294 ( 
.A(n_286),
.B(n_287),
.Y(n_294)
);


endmodule