module fake_netlist_1_591_n_27 (n_1, n_2, n_6, n_4, n_3, n_9, n_5, n_7, n_10, n_8, n_0, n_27);
input n_1;
input n_2;
input n_6;
input n_4;
input n_3;
input n_9;
input n_5;
input n_7;
input n_10;
input n_8;
input n_0;
output n_27;
wire n_20;
wire n_23;
wire n_22;
wire n_11;
wire n_25;
wire n_16;
wire n_26;
wire n_13;
wire n_18;
wire n_12;
wire n_17;
wire n_14;
wire n_15;
wire n_24;
wire n_19;
wire n_21;
CKINVDCx5p33_ASAP7_75t_R g11 ( .A(n_6), .Y(n_11) );
HB1xp67_ASAP7_75t_L g12 ( .A(n_10), .Y(n_12) );
BUFx2_ASAP7_75t_L g13 ( .A(n_8), .Y(n_13) );
BUFx2_ASAP7_75t_L g14 ( .A(n_2), .Y(n_14) );
BUFx3_ASAP7_75t_L g15 ( .A(n_7), .Y(n_15) );
OR2x6_ASAP7_75t_L g16 ( .A(n_14), .B(n_0), .Y(n_16) );
INVx2_ASAP7_75t_L g17 ( .A(n_15), .Y(n_17) );
AO221x2_ASAP7_75t_L g18 ( .A1(n_16), .A2(n_0), .B1(n_1), .B2(n_2), .C(n_3), .Y(n_18) );
AND2x2_ASAP7_75t_L g19 ( .A(n_18), .B(n_16), .Y(n_19) );
INVx2_ASAP7_75t_L g20 ( .A(n_19), .Y(n_20) );
OR2x2_ASAP7_75t_L g21 ( .A(n_20), .B(n_19), .Y(n_21) );
OAI22xp33_ASAP7_75t_SL g22 ( .A1(n_21), .A2(n_11), .B1(n_13), .B2(n_12), .Y(n_22) );
OAI32xp33_ASAP7_75t_L g23 ( .A1(n_21), .A2(n_15), .A3(n_11), .B1(n_17), .B2(n_5), .Y(n_23) );
NOR2xp33_ASAP7_75t_SL g24 ( .A(n_22), .B(n_1), .Y(n_24) );
BUFx4f_ASAP7_75t_SL g25 ( .A(n_24), .Y(n_25) );
AOI221xp5_ASAP7_75t_L g26 ( .A1(n_25), .A2(n_23), .B1(n_4), .B2(n_5), .C(n_3), .Y(n_26) );
NAND3xp33_ASAP7_75t_L g27 ( .A(n_26), .B(n_4), .C(n_9), .Y(n_27) );
endmodule