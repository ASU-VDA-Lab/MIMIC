module real_jpeg_30580_n_12 (n_5, n_4, n_8, n_0, n_1, n_11, n_2, n_6, n_7, n_3, n_10, n_9, n_12);

input n_5;
input n_4;
input n_8;
input n_0;
input n_1;
input n_11;
input n_2;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_12;

wire n_384;
wire n_37;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_300;
wire n_415;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_271;
wire n_47;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_13;
wire n_199;
wire n_95;
wire n_238;
wire n_67;
wire n_350;
wire n_235;
wire n_107;
wire n_369;
wire n_376;
wire n_354;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_355;
wire n_123;
wire n_50;
wire n_409;
wire n_186;
wire n_137;
wire n_72;
wire n_171;
wire n_151;
wire n_272;
wire n_198;
wire n_203;
wire n_23;
wire n_362;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_326;
wire n_339;
wire n_80;
wire n_30;
wire n_332;
wire n_149;
wire n_366;
wire n_328;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_353;
wire n_230;
wire n_417;
wire n_216;
wire n_128;
wire n_202;
wire n_367;
wire n_127;
wire n_356;
wire n_365;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_348;
wire n_252;
wire n_363;
wire n_310;
wire n_345;
wire n_78;
wire n_83;
wire n_288;
wire n_221;
wire n_393;
wire n_104;
wire n_153;
wire n_337;
wire n_131;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_378;
wire n_200;
wire n_335;
wire n_214;
wire n_113;
wire n_251;
wire n_139;
wire n_33;
wire n_338;
wire n_175;
wire n_156;
wire n_387;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_390;
wire n_77;
wire n_399;
wire n_372;
wire n_219;
wire n_122;
wire n_19;
wire n_262;
wire n_334;
wire n_17;
wire n_383;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_371;
wire n_410;
wire n_421;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_382;
wire n_411;
wire n_20;
wire n_278;
wire n_314;
wire n_103;
wire n_232;
wire n_212;
wire n_284;
wire n_402;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_213;
wire n_25;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_407;
wire n_419;
wire n_386;
wire n_341;
wire n_331;
wire n_49;
wire n_68;
wire n_395;
wire n_146;
wire n_286;
wire n_166;
wire n_176;
wire n_215;
wire n_323;
wire n_312;
wire n_325;
wire n_316;
wire n_307;
wire n_161;
wire n_207;
wire n_420;
wire n_357;
wire n_237;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_380;
wire n_414;
wire n_140;
wire n_126;
wire n_342;
wire n_120;
wire n_155;
wire n_412;
wire n_405;
wire n_319;
wire n_93;
wire n_242;
wire n_142;
wire n_397;
wire n_76;
wire n_403;
wire n_79;
wire n_282;
wire n_147;
wire n_359;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_18;
wire n_145;
wire n_266;
wire n_377;
wire n_109;
wire n_391;
wire n_401;
wire n_148;
wire n_373;
wire n_396;
wire n_392;
wire n_196;
wire n_375;
wire n_298;
wire n_330;
wire n_333;
wire n_152;
wire n_270;
wire n_159;
wire n_347;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_336;
wire n_258;
wire n_150;
wire n_41;
wire n_74;
wire n_404;
wire n_204;
wire n_158;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_413;
wire n_75;
wire n_346;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_119;
wire n_283;
wire n_181;
wire n_358;
wire n_256;
wire n_253;
wire n_273;
wire n_16;
wire n_54;
wire n_168;
wire n_38;
wire n_385;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_349;
wire n_418;
wire n_292;
wire n_343;
wire n_64;
wire n_291;
wire n_236;
wire n_370;
wire n_276;
wire n_374;
wire n_287;
wire n_388;
wire n_174;
wire n_400;
wire n_255;
wire n_243;
wire n_299;
wire n_352;
wire n_56;
wire n_293;
wire n_275;
wire n_381;
wire n_227;
wire n_229;
wire n_379;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_360;
wire n_398;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_45;
wire n_268;
wire n_42;
wire n_313;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_416;
wire n_143;
wire n_351;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_406;
wire n_303;
wire n_321;
wire n_100;
wire n_368;
wire n_51;
wire n_14;
wire n_205;
wire n_361;
wire n_261;
wire n_86;
wire n_324;
wire n_70;
wire n_32;
wire n_228;
wire n_389;
wire n_144;
wire n_15;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_394;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_133;
wire n_257;
wire n_344;
wire n_210;
wire n_206;
wire n_408;
wire n_85;
wire n_96;
wire n_308;
wire n_364;

BUFx12f_ASAP7_75t_L g131 ( 
.A(n_0),
.Y(n_131)
);

BUFx6f_ASAP7_75t_L g166 ( 
.A(n_0),
.Y(n_166)
);

BUFx3_ASAP7_75t_L g206 ( 
.A(n_0),
.Y(n_206)
);

HB1xp67_ASAP7_75t_L g259 ( 
.A(n_0),
.Y(n_259)
);

BUFx3_ASAP7_75t_L g296 ( 
.A(n_1),
.Y(n_296)
);

BUFx6f_ASAP7_75t_L g315 ( 
.A(n_1),
.Y(n_315)
);

BUFx6f_ASAP7_75t_L g82 ( 
.A(n_2),
.Y(n_82)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_2),
.Y(n_86)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_3),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_3),
.Y(n_35)
);

INVx4_ASAP7_75t_L g136 ( 
.A(n_3),
.Y(n_136)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_3),
.Y(n_242)
);

BUFx6f_ASAP7_75t_L g72 ( 
.A(n_4),
.Y(n_72)
);

BUFx6f_ASAP7_75t_L g98 ( 
.A(n_4),
.Y(n_98)
);

INVx2_ASAP7_75t_L g104 ( 
.A(n_4),
.Y(n_104)
);

BUFx6f_ASAP7_75t_L g305 ( 
.A(n_4),
.Y(n_305)
);

INVx2_ASAP7_75t_L g42 ( 
.A(n_5),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_5),
.Y(n_46)
);

BUFx3_ASAP7_75t_L g88 ( 
.A(n_5),
.Y(n_88)
);

BUFx6f_ASAP7_75t_L g151 ( 
.A(n_5),
.Y(n_151)
);

BUFx6f_ASAP7_75t_L g177 ( 
.A(n_6),
.Y(n_177)
);

OAI22xp5_ASAP7_75t_SL g61 ( 
.A1(n_7),
.A2(n_62),
.B1(n_63),
.B2(n_64),
.Y(n_61)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_7),
.Y(n_63)
);

OAI22xp5_ASAP7_75t_L g167 ( 
.A1(n_7),
.A2(n_63),
.B1(n_168),
.B2(n_170),
.Y(n_167)
);

AO22x2_ASAP7_75t_L g186 ( 
.A1(n_7),
.A2(n_63),
.B1(n_187),
.B2(n_189),
.Y(n_186)
);

OAI22xp5_ASAP7_75t_SL g350 ( 
.A1(n_7),
.A2(n_63),
.B1(n_351),
.B2(n_352),
.Y(n_350)
);

INVx2_ASAP7_75t_L g27 ( 
.A(n_8),
.Y(n_27)
);

INVx4_ASAP7_75t_L g33 ( 
.A(n_8),
.Y(n_33)
);

AOI22x1_ASAP7_75t_SL g91 ( 
.A1(n_9),
.A2(n_92),
.B1(n_94),
.B2(n_95),
.Y(n_91)
);

INVx2_ASAP7_75t_SL g94 ( 
.A(n_9),
.Y(n_94)
);

NAND2xp33_ASAP7_75t_SL g125 ( 
.A(n_9),
.B(n_126),
.Y(n_125)
);

AO22x1_ASAP7_75t_SL g138 ( 
.A1(n_9),
.A2(n_94),
.B1(n_139),
.B2(n_141),
.Y(n_138)
);

OAI22xp5_ASAP7_75t_SL g148 ( 
.A1(n_9),
.A2(n_94),
.B1(n_149),
.B2(n_152),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_SL g201 ( 
.A(n_9),
.B(n_75),
.Y(n_201)
);

OAI32xp33_ASAP7_75t_L g224 ( 
.A1(n_9),
.A2(n_225),
.A3(n_226),
.B1(n_230),
.B2(n_237),
.Y(n_224)
);

OAI22xp33_ASAP7_75t_L g36 ( 
.A1(n_10),
.A2(n_37),
.B1(n_38),
.B2(n_43),
.Y(n_36)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_10),
.Y(n_37)
);

OAI22xp33_ASAP7_75t_L g69 ( 
.A1(n_10),
.A2(n_37),
.B1(n_70),
.B2(n_73),
.Y(n_69)
);

OAI22xp33_ASAP7_75t_SL g208 ( 
.A1(n_10),
.A2(n_37),
.B1(n_209),
.B2(n_213),
.Y(n_208)
);

OAI22xp5_ASAP7_75t_SL g310 ( 
.A1(n_10),
.A2(n_37),
.B1(n_311),
.B2(n_316),
.Y(n_310)
);

AOI22xp5_ASAP7_75t_L g280 ( 
.A1(n_11),
.A2(n_225),
.B1(n_281),
.B2(n_282),
.Y(n_280)
);

INVx2_ASAP7_75t_SL g282 ( 
.A(n_11),
.Y(n_282)
);

OAI22xp5_ASAP7_75t_SL g361 ( 
.A1(n_11),
.A2(n_282),
.B1(n_362),
.B2(n_366),
.Y(n_361)
);

XNOR2xp5_ASAP7_75t_L g12 ( 
.A(n_13),
.B(n_394),
.Y(n_12)
);

INVx1_ASAP7_75t_L g13 ( 
.A(n_14),
.Y(n_13)
);

AOI21x1_ASAP7_75t_L g14 ( 
.A1(n_15),
.A2(n_338),
.B(n_389),
.Y(n_14)
);

BUFx2_ASAP7_75t_L g15 ( 
.A(n_16),
.Y(n_15)
);

AO21x1_ASAP7_75t_L g16 ( 
.A1(n_17),
.A2(n_272),
.B(n_337),
.Y(n_16)
);

OAI21x1_ASAP7_75t_SL g17 ( 
.A1(n_18),
.A2(n_194),
.B(n_271),
.Y(n_17)
);

NOR2x1_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_144),
.Y(n_18)
);

NAND2xp5_ASAP7_75t_L g271 ( 
.A(n_19),
.B(n_144),
.Y(n_271)
);

MAJIxp5_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_66),
.C(n_114),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_21),
.Y(n_20)
);

XOR2xp5_ASAP7_75t_L g216 ( 
.A(n_21),
.B(n_67),
.Y(n_216)
);

NAND2xp5_ASAP7_75t_L g21 ( 
.A(n_22),
.B(n_47),
.Y(n_21)
);

NAND2xp5_ASAP7_75t_L g244 ( 
.A(n_22),
.B(n_245),
.Y(n_244)
);

NAND2xp5_ASAP7_75t_L g22 ( 
.A(n_23),
.B(n_36),
.Y(n_22)
);

NAND2xp5_ASAP7_75t_L g147 ( 
.A(n_23),
.B(n_148),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_SL g199 ( 
.A(n_23),
.B(n_61),
.Y(n_199)
);

OA21x2_ASAP7_75t_L g335 ( 
.A1(n_23),
.A2(n_48),
.B(n_148),
.Y(n_335)
);

NAND2xp5_ASAP7_75t_L g360 ( 
.A(n_23),
.B(n_361),
.Y(n_360)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_24),
.Y(n_23)
);

AND2x2_ASAP7_75t_L g48 ( 
.A(n_24),
.B(n_49),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_R g250 ( 
.A(n_24),
.B(n_94),
.Y(n_250)
);

OA22x2_ASAP7_75t_L g24 ( 
.A1(n_25),
.A2(n_28),
.B1(n_31),
.B2(n_34),
.Y(n_24)
);

BUFx3_ASAP7_75t_L g25 ( 
.A(n_26),
.Y(n_25)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_26),
.Y(n_60)
);

INVx4_ASAP7_75t_L g236 ( 
.A(n_26),
.Y(n_236)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_27),
.Y(n_26)
);

INVx2_ASAP7_75t_L g28 ( 
.A(n_29),
.Y(n_28)
);

BUFx2_ASAP7_75t_L g255 ( 
.A(n_29),
.Y(n_255)
);

INVx6_ASAP7_75t_L g29 ( 
.A(n_30),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g140 ( 
.A(n_30),
.Y(n_140)
);

INVx2_ASAP7_75t_L g31 ( 
.A(n_32),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_33),
.Y(n_32)
);

INVx2_ASAP7_75t_L g54 ( 
.A(n_33),
.Y(n_54)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_35),
.Y(n_34)
);

INVx2_ASAP7_75t_L g142 ( 
.A(n_35),
.Y(n_142)
);

BUFx6f_ASAP7_75t_L g169 ( 
.A(n_35),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_L g155 ( 
.A(n_36),
.B(n_48),
.Y(n_155)
);

INVx2_ASAP7_75t_L g38 ( 
.A(n_39),
.Y(n_38)
);

INVx2_ASAP7_75t_L g39 ( 
.A(n_40),
.Y(n_39)
);

INVx2_ASAP7_75t_L g40 ( 
.A(n_41),
.Y(n_40)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_41),
.Y(n_62)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_41),
.Y(n_65)
);

BUFx5_ASAP7_75t_L g41 ( 
.A(n_42),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_42),
.Y(n_58)
);

BUFx3_ASAP7_75t_L g229 ( 
.A(n_42),
.Y(n_229)
);

INVx2_ASAP7_75t_L g43 ( 
.A(n_44),
.Y(n_43)
);

INVx2_ASAP7_75t_L g44 ( 
.A(n_45),
.Y(n_44)
);

INVx2_ASAP7_75t_L g45 ( 
.A(n_46),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_46),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g78 ( 
.A(n_46),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_L g359 ( 
.A(n_47),
.B(n_360),
.Y(n_359)
);

AOI22xp5_ASAP7_75t_L g413 ( 
.A1(n_47),
.A2(n_204),
.B1(n_265),
.B2(n_360),
.Y(n_413)
);

NAND2xp5_ASAP7_75t_L g47 ( 
.A(n_48),
.B(n_61),
.Y(n_47)
);

NAND2xp5_ASAP7_75t_L g245 ( 
.A(n_48),
.B(n_148),
.Y(n_245)
);

INVxp67_ASAP7_75t_L g409 ( 
.A(n_48),
.Y(n_409)
);

OAI22xp33_ASAP7_75t_L g49 ( 
.A1(n_50),
.A2(n_52),
.B1(n_55),
.B2(n_59),
.Y(n_49)
);

INVx4_ASAP7_75t_L g50 ( 
.A(n_51),
.Y(n_50)
);

INVx1_ASAP7_75t_SL g52 ( 
.A(n_53),
.Y(n_52)
);

INVx2_ASAP7_75t_SL g53 ( 
.A(n_54),
.Y(n_53)
);

INVx2_ASAP7_75t_L g55 ( 
.A(n_56),
.Y(n_55)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_57),
.Y(n_56)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_58),
.Y(n_57)
);

INVxp67_ASAP7_75t_SL g59 ( 
.A(n_60),
.Y(n_59)
);

INVx3_ASAP7_75t_L g123 ( 
.A(n_64),
.Y(n_123)
);

INVx2_ASAP7_75t_L g64 ( 
.A(n_65),
.Y(n_64)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_67),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_L g67 ( 
.A(n_68),
.B(n_89),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_L g332 ( 
.A(n_68),
.B(n_333),
.Y(n_332)
);

NAND2xp33_ASAP7_75t_SL g68 ( 
.A(n_69),
.B(n_75),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_L g192 ( 
.A(n_69),
.B(n_193),
.Y(n_192)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_71),
.Y(n_70)
);

INVx2_ASAP7_75t_L g74 ( 
.A(n_71),
.Y(n_74)
);

INVx2_ASAP7_75t_L g93 ( 
.A(n_71),
.Y(n_93)
);

INVx3_ASAP7_75t_L g188 ( 
.A(n_71),
.Y(n_188)
);

INVx8_ASAP7_75t_L g71 ( 
.A(n_72),
.Y(n_71)
);

INVx3_ASAP7_75t_L g110 ( 
.A(n_72),
.Y(n_110)
);

INVx2_ASAP7_75t_L g73 ( 
.A(n_74),
.Y(n_73)
);

AND2x4_ASAP7_75t_L g185 ( 
.A(n_75),
.B(n_186),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_L g345 ( 
.A(n_75),
.B(n_346),
.Y(n_345)
);

INVx1_ASAP7_75t_L g372 ( 
.A(n_75),
.Y(n_372)
);

INVx2_ASAP7_75t_L g75 ( 
.A(n_76),
.Y(n_75)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_77),
.Y(n_76)
);

AO21x2_ASAP7_75t_L g99 ( 
.A1(n_77),
.A2(n_100),
.B(n_108),
.Y(n_99)
);

OAI22xp5_ASAP7_75t_L g77 ( 
.A1(n_78),
.A2(n_79),
.B1(n_83),
.B2(n_87),
.Y(n_77)
);

INVx2_ASAP7_75t_L g79 ( 
.A(n_80),
.Y(n_79)
);

INVx2_ASAP7_75t_L g80 ( 
.A(n_81),
.Y(n_80)
);

INVx3_ASAP7_75t_L g81 ( 
.A(n_82),
.Y(n_81)
);

BUFx6f_ASAP7_75t_L g107 ( 
.A(n_82),
.Y(n_107)
);

INVx2_ASAP7_75t_L g83 ( 
.A(n_84),
.Y(n_83)
);

INVx2_ASAP7_75t_L g84 ( 
.A(n_85),
.Y(n_84)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_86),
.Y(n_85)
);

BUFx6f_ASAP7_75t_L g113 ( 
.A(n_86),
.Y(n_113)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_88),
.Y(n_87)
);

BUFx6f_ASAP7_75t_L g128 ( 
.A(n_88),
.Y(n_128)
);

INVx2_ASAP7_75t_L g365 ( 
.A(n_88),
.Y(n_365)
);

INVxp67_ASAP7_75t_L g89 ( 
.A(n_90),
.Y(n_89)
);

NOR2x1_ASAP7_75t_L g415 ( 
.A(n_90),
.B(n_185),
.Y(n_415)
);

NOR2x1_ASAP7_75t_L g90 ( 
.A(n_91),
.B(n_99),
.Y(n_90)
);

INVx1_ASAP7_75t_L g346 ( 
.A(n_91),
.Y(n_346)
);

AOI21x1_ASAP7_75t_L g371 ( 
.A1(n_91),
.A2(n_99),
.B(n_372),
.Y(n_371)
);

INVxp67_ASAP7_75t_SL g92 ( 
.A(n_93),
.Y(n_92)
);

AOI32xp33_ASAP7_75t_L g117 ( 
.A1(n_94),
.A2(n_118),
.A3(n_122),
.B1(n_124),
.B2(n_125),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_SL g173 ( 
.A(n_94),
.B(n_174),
.Y(n_173)
);

NOR2xp33_ASAP7_75t_L g237 ( 
.A(n_94),
.B(n_238),
.Y(n_237)
);

NOR2xp33_ASAP7_75t_L g256 ( 
.A(n_94),
.B(n_257),
.Y(n_256)
);

NAND2xp5_ASAP7_75t_L g292 ( 
.A(n_94),
.B(n_293),
.Y(n_292)
);

OAI21xp5_ASAP7_75t_SL g319 ( 
.A1(n_94),
.A2(n_292),
.B(n_320),
.Y(n_319)
);

INVx2_ASAP7_75t_L g95 ( 
.A(n_96),
.Y(n_95)
);

INVx3_ASAP7_75t_L g96 ( 
.A(n_97),
.Y(n_96)
);

BUFx6f_ASAP7_75t_L g97 ( 
.A(n_98),
.Y(n_97)
);

BUFx6f_ASAP7_75t_L g121 ( 
.A(n_98),
.Y(n_121)
);

BUFx6f_ASAP7_75t_L g179 ( 
.A(n_98),
.Y(n_179)
);

BUFx6f_ASAP7_75t_L g191 ( 
.A(n_98),
.Y(n_191)
);

INVx2_ASAP7_75t_L g193 ( 
.A(n_99),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_L g100 ( 
.A(n_101),
.B(n_105),
.Y(n_100)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_102),
.Y(n_101)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_103),
.Y(n_102)
);

BUFx6f_ASAP7_75t_L g103 ( 
.A(n_104),
.Y(n_103)
);

BUFx6f_ASAP7_75t_L g178 ( 
.A(n_104),
.Y(n_178)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_106),
.Y(n_105)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_107),
.Y(n_106)
);

INVxp33_ASAP7_75t_L g124 ( 
.A(n_108),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_L g108 ( 
.A(n_109),
.B(n_111),
.Y(n_108)
);

INVx3_ASAP7_75t_SL g109 ( 
.A(n_110),
.Y(n_109)
);

INVx4_ASAP7_75t_L g111 ( 
.A(n_112),
.Y(n_111)
);

INVx5_ASAP7_75t_L g112 ( 
.A(n_113),
.Y(n_112)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_115),
.Y(n_114)
);

XNOR2xp5_ASAP7_75t_L g215 ( 
.A(n_115),
.B(n_216),
.Y(n_215)
);

OAI22xp33_ASAP7_75t_L g115 ( 
.A1(n_116),
.A2(n_117),
.B1(n_129),
.B2(n_143),
.Y(n_115)
);

INVxp67_ASAP7_75t_L g116 ( 
.A(n_117),
.Y(n_116)
);

NOR2x1_ASAP7_75t_SL g156 ( 
.A(n_117),
.B(n_129),
.Y(n_156)
);

INVx3_ASAP7_75t_L g118 ( 
.A(n_119),
.Y(n_118)
);

BUFx3_ASAP7_75t_L g119 ( 
.A(n_120),
.Y(n_119)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_121),
.Y(n_120)
);

INVx4_ASAP7_75t_L g122 ( 
.A(n_123),
.Y(n_122)
);

INVx4_ASAP7_75t_L g126 ( 
.A(n_127),
.Y(n_126)
);

INVx4_ASAP7_75t_L g127 ( 
.A(n_128),
.Y(n_127)
);

BUFx6f_ASAP7_75t_L g367 ( 
.A(n_128),
.Y(n_367)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_129),
.Y(n_143)
);

OAI22xp5_ASAP7_75t_L g405 ( 
.A1(n_129),
.A2(n_143),
.B1(n_406),
.B2(n_410),
.Y(n_405)
);

AO21x2_ASAP7_75t_L g129 ( 
.A1(n_130),
.A2(n_132),
.B(n_137),
.Y(n_129)
);

AND2x2_ASAP7_75t_L g133 ( 
.A(n_130),
.B(n_134),
.Y(n_133)
);

INVx4_ASAP7_75t_SL g130 ( 
.A(n_131),
.Y(n_130)
);

OAI21xp33_ASAP7_75t_L g260 ( 
.A1(n_132),
.A2(n_137),
.B(n_261),
.Y(n_260)
);

OAI21xp5_ASAP7_75t_L g377 ( 
.A1(n_132),
.A2(n_162),
.B(n_280),
.Y(n_377)
);

INVx2_ASAP7_75t_L g132 ( 
.A(n_133),
.Y(n_132)
);

AOI21xp5_ASAP7_75t_L g160 ( 
.A1(n_133),
.A2(n_138),
.B(n_161),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_SL g207 ( 
.A(n_133),
.B(n_208),
.Y(n_207)
);

NAND2xp5_ASAP7_75t_SL g265 ( 
.A(n_133),
.B(n_167),
.Y(n_265)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_134),
.Y(n_281)
);

BUFx6f_ASAP7_75t_L g134 ( 
.A(n_135),
.Y(n_134)
);

INVx2_ASAP7_75t_L g135 ( 
.A(n_136),
.Y(n_135)
);

BUFx6f_ASAP7_75t_L g171 ( 
.A(n_136),
.Y(n_171)
);

BUFx6f_ASAP7_75t_L g212 ( 
.A(n_136),
.Y(n_212)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_138),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_L g204 ( 
.A(n_138),
.B(n_205),
.Y(n_204)
);

INVx2_ASAP7_75t_L g139 ( 
.A(n_140),
.Y(n_139)
);

INVx4_ASAP7_75t_L g141 ( 
.A(n_142),
.Y(n_141)
);

XOR2xp5_ASAP7_75t_L g144 ( 
.A(n_145),
.B(n_157),
.Y(n_144)
);

XOR2xp5_ASAP7_75t_L g145 ( 
.A(n_146),
.B(n_156),
.Y(n_145)
);

MAJIxp5_ASAP7_75t_L g273 ( 
.A(n_146),
.B(n_156),
.C(n_157),
.Y(n_273)
);

NAND2xp5_ASAP7_75t_L g146 ( 
.A(n_147),
.B(n_155),
.Y(n_146)
);

BUFx6f_ASAP7_75t_L g149 ( 
.A(n_150),
.Y(n_149)
);

INVx5_ASAP7_75t_L g233 ( 
.A(n_150),
.Y(n_233)
);

BUFx6f_ASAP7_75t_L g150 ( 
.A(n_151),
.Y(n_150)
);

INVx2_ASAP7_75t_L g154 ( 
.A(n_151),
.Y(n_154)
);

INVx2_ASAP7_75t_SL g152 ( 
.A(n_153),
.Y(n_152)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_154),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_L g198 ( 
.A(n_155),
.B(n_199),
.Y(n_198)
);

XOR2x2_ASAP7_75t_L g157 ( 
.A(n_158),
.B(n_182),
.Y(n_157)
);

OAI22xp5_ASAP7_75t_SL g158 ( 
.A1(n_159),
.A2(n_160),
.B1(n_172),
.B2(n_173),
.Y(n_158)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_160),
.Y(n_159)
);

MAJx2_ASAP7_75t_L g306 ( 
.A(n_160),
.B(n_172),
.C(n_183),
.Y(n_306)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_162),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_L g249 ( 
.A(n_162),
.B(n_207),
.Y(n_249)
);

NAND2xp5_ASAP7_75t_L g162 ( 
.A(n_163),
.B(n_167),
.Y(n_162)
);

BUFx6f_ASAP7_75t_L g163 ( 
.A(n_164),
.Y(n_163)
);

INVx3_ASAP7_75t_L g164 ( 
.A(n_165),
.Y(n_164)
);

INVx2_ASAP7_75t_L g165 ( 
.A(n_166),
.Y(n_165)
);

BUFx3_ASAP7_75t_L g279 ( 
.A(n_166),
.Y(n_279)
);

INVx2_ASAP7_75t_L g168 ( 
.A(n_169),
.Y(n_168)
);

BUFx2_ASAP7_75t_SL g214 ( 
.A(n_169),
.Y(n_214)
);

INVx6_ASAP7_75t_L g170 ( 
.A(n_171),
.Y(n_170)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_173),
.Y(n_172)
);

INVx1_ASAP7_75t_L g353 ( 
.A(n_174),
.Y(n_353)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_175),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_SL g309 ( 
.A(n_175),
.B(n_310),
.Y(n_309)
);

NOR2x1p5_ASAP7_75t_L g323 ( 
.A(n_175),
.B(n_324),
.Y(n_323)
);

AO22x2_ASAP7_75t_L g175 ( 
.A1(n_176),
.A2(n_178),
.B1(n_179),
.B2(n_180),
.Y(n_175)
);

BUFx2_ASAP7_75t_L g301 ( 
.A(n_176),
.Y(n_301)
);

BUFx6f_ASAP7_75t_L g176 ( 
.A(n_177),
.Y(n_176)
);

BUFx6f_ASAP7_75t_L g181 ( 
.A(n_177),
.Y(n_181)
);

BUFx6f_ASAP7_75t_L g288 ( 
.A(n_177),
.Y(n_288)
);

INVx2_ASAP7_75t_L g330 ( 
.A(n_177),
.Y(n_330)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_178),
.Y(n_290)
);

INVx2_ASAP7_75t_L g180 ( 
.A(n_181),
.Y(n_180)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_183),
.Y(n_182)
);

AND2x2_ASAP7_75t_L g183 ( 
.A(n_184),
.B(n_192),
.Y(n_183)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_185),
.Y(n_184)
);

NAND2x1_ASAP7_75t_L g333 ( 
.A(n_186),
.B(n_193),
.Y(n_333)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_188),
.Y(n_187)
);

INVx3_ASAP7_75t_L g189 ( 
.A(n_190),
.Y(n_189)
);

INVx2_ASAP7_75t_L g190 ( 
.A(n_191),
.Y(n_190)
);

NAND2xp5_ASAP7_75t_L g344 ( 
.A(n_192),
.B(n_345),
.Y(n_344)
);

AOI21x1_ASAP7_75t_L g194 ( 
.A1(n_195),
.A2(n_217),
.B(n_270),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_L g195 ( 
.A(n_196),
.B(n_215),
.Y(n_195)
);

NOR2xp67_ASAP7_75t_SL g270 ( 
.A(n_196),
.B(n_215),
.Y(n_270)
);

MAJIxp5_ASAP7_75t_L g196 ( 
.A(n_197),
.B(n_200),
.C(n_202),
.Y(n_196)
);

HB1xp67_ASAP7_75t_L g197 ( 
.A(n_198),
.Y(n_197)
);

OAI22xp5_ASAP7_75t_L g220 ( 
.A1(n_198),
.A2(n_200),
.B1(n_201),
.B2(n_221),
.Y(n_220)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_198),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_L g376 ( 
.A(n_199),
.B(n_245),
.Y(n_376)
);

OAI21xp5_ASAP7_75t_L g407 ( 
.A1(n_199),
.A2(n_408),
.B(n_409),
.Y(n_407)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_201),
.Y(n_200)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_203),
.Y(n_202)
);

XNOR2xp5_ASAP7_75t_L g219 ( 
.A(n_203),
.B(n_220),
.Y(n_219)
);

AND2x2_ASAP7_75t_L g203 ( 
.A(n_204),
.B(n_207),
.Y(n_203)
);

AND2x2_ASAP7_75t_L g368 ( 
.A(n_204),
.B(n_265),
.Y(n_368)
);

BUFx6f_ASAP7_75t_L g205 ( 
.A(n_206),
.Y(n_205)
);

NAND2xp5_ASAP7_75t_L g261 ( 
.A(n_208),
.B(n_258),
.Y(n_261)
);

INVx4_ASAP7_75t_L g209 ( 
.A(n_210),
.Y(n_209)
);

INVx2_ASAP7_75t_L g210 ( 
.A(n_211),
.Y(n_210)
);

INVx2_ASAP7_75t_L g211 ( 
.A(n_212),
.Y(n_211)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_212),
.Y(n_225)
);

INVx2_ASAP7_75t_L g213 ( 
.A(n_214),
.Y(n_213)
);

OAI21xp5_ASAP7_75t_L g217 ( 
.A1(n_218),
.A2(n_246),
.B(n_269),
.Y(n_217)
);

NOR2xp67_ASAP7_75t_L g218 ( 
.A(n_219),
.B(n_222),
.Y(n_218)
);

NAND2xp5_ASAP7_75t_L g269 ( 
.A(n_219),
.B(n_222),
.Y(n_269)
);

NOR2xp33_ASAP7_75t_L g222 ( 
.A(n_223),
.B(n_243),
.Y(n_222)
);

NAND2xp33_ASAP7_75t_SL g266 ( 
.A(n_223),
.B(n_244),
.Y(n_266)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_224),
.Y(n_223)
);

NAND2xp5_ASAP7_75t_L g267 ( 
.A(n_224),
.B(n_243),
.Y(n_267)
);

INVx3_ASAP7_75t_L g226 ( 
.A(n_227),
.Y(n_226)
);

INVx4_ASAP7_75t_L g227 ( 
.A(n_228),
.Y(n_227)
);

BUFx3_ASAP7_75t_L g228 ( 
.A(n_229),
.Y(n_228)
);

NAND2xp5_ASAP7_75t_L g230 ( 
.A(n_231),
.B(n_234),
.Y(n_230)
);

INVx2_ASAP7_75t_L g231 ( 
.A(n_232),
.Y(n_231)
);

BUFx6f_ASAP7_75t_L g232 ( 
.A(n_233),
.Y(n_232)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_235),
.Y(n_234)
);

HB1xp67_ASAP7_75t_L g235 ( 
.A(n_236),
.Y(n_235)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_239),
.Y(n_238)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_240),
.Y(n_239)
);

INVx2_ASAP7_75t_L g240 ( 
.A(n_241),
.Y(n_240)
);

INVx2_ASAP7_75t_L g241 ( 
.A(n_242),
.Y(n_241)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_244),
.Y(n_243)
);

AOI21x1_ASAP7_75t_SL g246 ( 
.A1(n_247),
.A2(n_263),
.B(n_268),
.Y(n_246)
);

OAI21xp5_ASAP7_75t_L g247 ( 
.A1(n_248),
.A2(n_251),
.B(n_262),
.Y(n_247)
);

NOR2xp33_ASAP7_75t_SL g248 ( 
.A(n_249),
.B(n_250),
.Y(n_248)
);

NAND2xp5_ASAP7_75t_L g262 ( 
.A(n_249),
.B(n_250),
.Y(n_262)
);

NAND2xp5_ASAP7_75t_L g251 ( 
.A(n_252),
.B(n_260),
.Y(n_251)
);

NOR2xp33_ASAP7_75t_L g252 ( 
.A(n_253),
.B(n_256),
.Y(n_252)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_254),
.Y(n_253)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_255),
.Y(n_254)
);

INVx2_ASAP7_75t_L g257 ( 
.A(n_258),
.Y(n_257)
);

BUFx4f_ASAP7_75t_L g258 ( 
.A(n_259),
.Y(n_258)
);

AND2x2_ASAP7_75t_L g264 ( 
.A(n_261),
.B(n_265),
.Y(n_264)
);

NAND3xp33_ASAP7_75t_SL g263 ( 
.A(n_264),
.B(n_266),
.C(n_267),
.Y(n_263)
);

AOI21xp5_ASAP7_75t_L g268 ( 
.A1(n_264),
.A2(n_266),
.B(n_267),
.Y(n_268)
);

OAI21xp5_ASAP7_75t_L g277 ( 
.A1(n_265),
.A2(n_278),
.B(n_280),
.Y(n_277)
);

NAND2xp5_ASAP7_75t_L g272 ( 
.A(n_273),
.B(n_274),
.Y(n_272)
);

NOR2xp67_ASAP7_75t_L g337 ( 
.A(n_273),
.B(n_274),
.Y(n_337)
);

XOR2xp5_ASAP7_75t_L g274 ( 
.A(n_275),
.B(n_307),
.Y(n_274)
);

XOR2xp5_ASAP7_75t_L g275 ( 
.A(n_276),
.B(n_306),
.Y(n_275)
);

MAJIxp5_ASAP7_75t_L g386 ( 
.A(n_276),
.B(n_306),
.C(n_307),
.Y(n_386)
);

XNOR2xp5_ASAP7_75t_L g276 ( 
.A(n_277),
.B(n_283),
.Y(n_276)
);

OAI21xp5_ASAP7_75t_L g354 ( 
.A1(n_277),
.A2(n_355),
.B(n_356),
.Y(n_354)
);

INVx3_ASAP7_75t_L g278 ( 
.A(n_279),
.Y(n_278)
);

NAND2xp5_ASAP7_75t_L g283 ( 
.A(n_284),
.B(n_297),
.Y(n_283)
);

INVx1_ASAP7_75t_L g356 ( 
.A(n_284),
.Y(n_356)
);

OAI21xp5_ASAP7_75t_L g284 ( 
.A1(n_285),
.A2(n_289),
.B(n_291),
.Y(n_284)
);

INVx1_ASAP7_75t_SL g285 ( 
.A(n_286),
.Y(n_285)
);

INVx2_ASAP7_75t_L g286 ( 
.A(n_287),
.Y(n_286)
);

INVx2_ASAP7_75t_L g287 ( 
.A(n_288),
.Y(n_287)
);

INVx2_ASAP7_75t_L g326 ( 
.A(n_288),
.Y(n_326)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_290),
.Y(n_289)
);

INVxp67_ASAP7_75t_L g291 ( 
.A(n_292),
.Y(n_291)
);

INVx3_ASAP7_75t_L g352 ( 
.A(n_293),
.Y(n_352)
);

INVx2_ASAP7_75t_L g293 ( 
.A(n_294),
.Y(n_293)
);

BUFx6f_ASAP7_75t_L g299 ( 
.A(n_294),
.Y(n_299)
);

INVx2_ASAP7_75t_L g325 ( 
.A(n_294),
.Y(n_325)
);

INVx6_ASAP7_75t_L g294 ( 
.A(n_295),
.Y(n_294)
);

BUFx6f_ASAP7_75t_L g295 ( 
.A(n_296),
.Y(n_295)
);

BUFx6f_ASAP7_75t_L g328 ( 
.A(n_296),
.Y(n_328)
);

INVx1_ASAP7_75t_L g355 ( 
.A(n_297),
.Y(n_355)
);

NAND3xp33_ASAP7_75t_L g297 ( 
.A(n_298),
.B(n_300),
.C(n_302),
.Y(n_297)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_299),
.Y(n_298)
);

INVx2_ASAP7_75t_L g300 ( 
.A(n_301),
.Y(n_300)
);

INVx3_ASAP7_75t_SL g302 ( 
.A(n_303),
.Y(n_302)
);

INVx4_ASAP7_75t_L g303 ( 
.A(n_304),
.Y(n_303)
);

INVx8_ASAP7_75t_L g304 ( 
.A(n_305),
.Y(n_304)
);

XNOR2xp5_ASAP7_75t_L g307 ( 
.A(n_308),
.B(n_331),
.Y(n_307)
);

MAJx2_ASAP7_75t_L g382 ( 
.A(n_308),
.B(n_332),
.C(n_335),
.Y(n_382)
);

NAND2xp5_ASAP7_75t_L g308 ( 
.A(n_309),
.B(n_318),
.Y(n_308)
);

NAND2xp5_ASAP7_75t_L g373 ( 
.A(n_309),
.B(n_374),
.Y(n_373)
);

NAND2xp5_ASAP7_75t_L g348 ( 
.A(n_310),
.B(n_323),
.Y(n_348)
);

INVx2_ASAP7_75t_L g311 ( 
.A(n_312),
.Y(n_311)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_313),
.Y(n_312)
);

INVx3_ASAP7_75t_L g313 ( 
.A(n_314),
.Y(n_313)
);

INVx6_ASAP7_75t_L g314 ( 
.A(n_315),
.Y(n_314)
);

BUFx6f_ASAP7_75t_L g317 ( 
.A(n_315),
.Y(n_317)
);

BUFx3_ASAP7_75t_L g322 ( 
.A(n_315),
.Y(n_322)
);

INVx2_ASAP7_75t_L g316 ( 
.A(n_317),
.Y(n_316)
);

BUFx6f_ASAP7_75t_L g351 ( 
.A(n_317),
.Y(n_351)
);

NAND2xp5_ASAP7_75t_L g318 ( 
.A(n_319),
.B(n_323),
.Y(n_318)
);

NAND2xp5_ASAP7_75t_L g417 ( 
.A(n_319),
.B(n_353),
.Y(n_417)
);

INVx4_ASAP7_75t_L g320 ( 
.A(n_321),
.Y(n_320)
);

INVx2_ASAP7_75t_L g321 ( 
.A(n_322),
.Y(n_321)
);

NAND2xp5_ASAP7_75t_L g374 ( 
.A(n_323),
.B(n_350),
.Y(n_374)
);

AOI22xp5_ASAP7_75t_L g324 ( 
.A1(n_325),
.A2(n_326),
.B1(n_327),
.B2(n_329),
.Y(n_324)
);

INVx2_ASAP7_75t_L g327 ( 
.A(n_328),
.Y(n_327)
);

INVx4_ASAP7_75t_L g329 ( 
.A(n_330),
.Y(n_329)
);

OAI22xp33_ASAP7_75t_SL g331 ( 
.A1(n_332),
.A2(n_334),
.B1(n_335),
.B2(n_336),
.Y(n_331)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_332),
.Y(n_336)
);

INVx2_ASAP7_75t_SL g334 ( 
.A(n_335),
.Y(n_334)
);

INVxp67_ASAP7_75t_L g338 ( 
.A(n_339),
.Y(n_338)
);

NAND2xp5_ASAP7_75t_L g339 ( 
.A(n_340),
.B(n_385),
.Y(n_339)
);

NAND2xp5_ASAP7_75t_L g391 ( 
.A(n_340),
.B(n_392),
.Y(n_391)
);

NAND2x1_ASAP7_75t_L g340 ( 
.A(n_341),
.B(n_378),
.Y(n_340)
);

OR2x2_ASAP7_75t_L g393 ( 
.A(n_341),
.B(n_378),
.Y(n_393)
);

XNOR2xp5_ASAP7_75t_L g341 ( 
.A(n_342),
.B(n_357),
.Y(n_341)
);

MAJIxp5_ASAP7_75t_L g396 ( 
.A(n_342),
.B(n_358),
.C(n_397),
.Y(n_396)
);

MAJIxp5_ASAP7_75t_L g342 ( 
.A(n_343),
.B(n_347),
.C(n_354),
.Y(n_342)
);

OAI22xp5_ASAP7_75t_L g380 ( 
.A1(n_343),
.A2(n_344),
.B1(n_347),
.B2(n_381),
.Y(n_380)
);

INVx1_ASAP7_75t_L g343 ( 
.A(n_344),
.Y(n_343)
);

INVx1_ASAP7_75t_L g381 ( 
.A(n_347),
.Y(n_381)
);

AND2x2_ASAP7_75t_L g347 ( 
.A(n_348),
.B(n_349),
.Y(n_347)
);

NAND2xp5_ASAP7_75t_L g416 ( 
.A(n_348),
.B(n_417),
.Y(n_416)
);

AND2x2_ASAP7_75t_L g419 ( 
.A(n_348),
.B(n_417),
.Y(n_419)
);

NAND2xp5_ASAP7_75t_L g349 ( 
.A(n_350),
.B(n_353),
.Y(n_349)
);

XNOR2xp5_ASAP7_75t_L g379 ( 
.A(n_354),
.B(n_380),
.Y(n_379)
);

XOR2xp5_ASAP7_75t_L g357 ( 
.A(n_358),
.B(n_369),
.Y(n_357)
);

XNOR2x2_ASAP7_75t_L g358 ( 
.A(n_359),
.B(n_368),
.Y(n_358)
);

INVx1_ASAP7_75t_L g408 ( 
.A(n_361),
.Y(n_408)
);

INVx1_ASAP7_75t_L g362 ( 
.A(n_363),
.Y(n_362)
);

INVx2_ASAP7_75t_L g363 ( 
.A(n_364),
.Y(n_363)
);

INVx3_ASAP7_75t_SL g364 ( 
.A(n_365),
.Y(n_364)
);

INVx3_ASAP7_75t_L g366 ( 
.A(n_367),
.Y(n_366)
);

HB1xp67_ASAP7_75t_L g397 ( 
.A(n_369),
.Y(n_397)
);

XNOR2xp5_ASAP7_75t_L g369 ( 
.A(n_370),
.B(n_375),
.Y(n_369)
);

XOR2xp5_ASAP7_75t_L g370 ( 
.A(n_371),
.B(n_373),
.Y(n_370)
);

HB1xp67_ASAP7_75t_L g403 ( 
.A(n_371),
.Y(n_403)
);

HB1xp67_ASAP7_75t_L g402 ( 
.A(n_373),
.Y(n_402)
);

HB1xp67_ASAP7_75t_L g401 ( 
.A(n_375),
.Y(n_401)
);

NAND2xp5_ASAP7_75t_L g375 ( 
.A(n_376),
.B(n_377),
.Y(n_375)
);

INVx1_ASAP7_75t_L g384 ( 
.A(n_376),
.Y(n_384)
);

XNOR2x1_ASAP7_75t_L g383 ( 
.A(n_377),
.B(n_384),
.Y(n_383)
);

MAJIxp5_ASAP7_75t_L g378 ( 
.A(n_379),
.B(n_382),
.C(n_383),
.Y(n_378)
);

XOR2xp5_ASAP7_75t_L g387 ( 
.A(n_379),
.B(n_388),
.Y(n_387)
);

XOR2xp5_ASAP7_75t_L g388 ( 
.A(n_382),
.B(n_383),
.Y(n_388)
);

OR2x2_ASAP7_75t_L g385 ( 
.A(n_386),
.B(n_387),
.Y(n_385)
);

AND2x2_ASAP7_75t_L g392 ( 
.A(n_386),
.B(n_387),
.Y(n_392)
);

NAND2xp5_ASAP7_75t_SL g389 ( 
.A(n_390),
.B(n_393),
.Y(n_389)
);

HB1xp67_ASAP7_75t_L g390 ( 
.A(n_391),
.Y(n_390)
);

NOR2xp33_ASAP7_75t_L g394 ( 
.A(n_395),
.B(n_420),
.Y(n_394)
);

AND2x2_ASAP7_75t_L g395 ( 
.A(n_396),
.B(n_398),
.Y(n_395)
);

OR2x2_ASAP7_75t_L g421 ( 
.A(n_396),
.B(n_398),
.Y(n_421)
);

XNOR2xp5_ASAP7_75t_L g398 ( 
.A(n_399),
.B(n_404),
.Y(n_398)
);

MAJIxp5_ASAP7_75t_L g399 ( 
.A(n_400),
.B(n_402),
.C(n_403),
.Y(n_399)
);

INVxp67_ASAP7_75t_SL g400 ( 
.A(n_401),
.Y(n_400)
);

XOR2xp5_ASAP7_75t_L g404 ( 
.A(n_405),
.B(n_411),
.Y(n_404)
);

INVx1_ASAP7_75t_L g410 ( 
.A(n_406),
.Y(n_410)
);

INVx1_ASAP7_75t_L g406 ( 
.A(n_407),
.Y(n_406)
);

XNOR2x1_ASAP7_75t_L g411 ( 
.A(n_412),
.B(n_414),
.Y(n_411)
);

INVx1_ASAP7_75t_L g412 ( 
.A(n_413),
.Y(n_412)
);

AOI22x1_ASAP7_75t_L g414 ( 
.A1(n_415),
.A2(n_416),
.B1(n_418),
.B2(n_419),
.Y(n_414)
);

INVx2_ASAP7_75t_L g418 ( 
.A(n_415),
.Y(n_418)
);

INVx2_ASAP7_75t_L g420 ( 
.A(n_421),
.Y(n_420)
);


endmodule