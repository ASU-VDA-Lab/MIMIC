module fake_jpeg_29311_n_179 (n_13, n_21, n_33, n_1, n_45, n_10, n_23, n_27, n_6, n_22, n_47, n_14, n_40, n_19, n_18, n_20, n_35, n_48, n_46, n_41, n_4, n_34, n_30, n_39, n_42, n_16, n_49, n_3, n_0, n_24, n_28, n_38, n_26, n_44, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_43, n_50, n_12, n_32, n_8, n_15, n_7, n_179);

input n_13;
input n_21;
input n_33;
input n_1;
input n_45;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_47;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_48;
input n_46;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_42;
input n_16;
input n_49;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_44;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_43;
input n_50;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_179;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_51;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_84;
wire n_59;
wire n_98;
wire n_178;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_76;
wire n_154;
wire n_127;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_155;
wire n_103;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_175;
wire n_57;
wire n_171;
wire n_119;
wire n_69;
wire n_83;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_168;
wire n_106;
wire n_111;
wire n_143;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_177;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_54;
wire n_91;
wire n_93;
wire n_161;
wire n_138;
wire n_101;
wire n_149;
wire n_157;
wire n_87;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_176;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_62;
wire n_167;
wire n_174;
wire n_120;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_20),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_31),
.Y(n_52)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_34),
.Y(n_53)
);

INVx13_ASAP7_75t_L g54 ( 
.A(n_29),
.Y(n_54)
);

CKINVDCx20_ASAP7_75t_R g55 ( 
.A(n_9),
.Y(n_55)
);

INVx11_ASAP7_75t_L g56 ( 
.A(n_15),
.Y(n_56)
);

CKINVDCx20_ASAP7_75t_R g57 ( 
.A(n_11),
.Y(n_57)
);

INVx11_ASAP7_75t_L g58 ( 
.A(n_18),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_25),
.Y(n_59)
);

INVx3_ASAP7_75t_L g60 ( 
.A(n_11),
.Y(n_60)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_42),
.Y(n_61)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_37),
.Y(n_62)
);

CKINVDCx20_ASAP7_75t_R g63 ( 
.A(n_49),
.Y(n_63)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_46),
.Y(n_64)
);

CKINVDCx20_ASAP7_75t_R g65 ( 
.A(n_41),
.Y(n_65)
);

CKINVDCx20_ASAP7_75t_R g66 ( 
.A(n_30),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_16),
.Y(n_67)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_3),
.Y(n_68)
);

CKINVDCx20_ASAP7_75t_R g69 ( 
.A(n_33),
.Y(n_69)
);

BUFx12_ASAP7_75t_L g70 ( 
.A(n_6),
.Y(n_70)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_35),
.Y(n_71)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_44),
.Y(n_72)
);

CKINVDCx20_ASAP7_75t_R g73 ( 
.A(n_26),
.Y(n_73)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_45),
.Y(n_74)
);

INVx11_ASAP7_75t_L g75 ( 
.A(n_9),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_SL g76 ( 
.A(n_55),
.B(n_0),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_L g91 ( 
.A(n_76),
.B(n_1),
.Y(n_91)
);

INVx3_ASAP7_75t_L g77 ( 
.A(n_54),
.Y(n_77)
);

INVx4_ASAP7_75t_L g89 ( 
.A(n_77),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_57),
.B(n_0),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_78),
.B(n_79),
.Y(n_86)
);

CKINVDCx20_ASAP7_75t_R g79 ( 
.A(n_51),
.Y(n_79)
);

INVx8_ASAP7_75t_L g80 ( 
.A(n_52),
.Y(n_80)
);

INVx4_ASAP7_75t_L g90 ( 
.A(n_80),
.Y(n_90)
);

INVx2_ASAP7_75t_L g81 ( 
.A(n_60),
.Y(n_81)
);

INVx2_ASAP7_75t_L g97 ( 
.A(n_81),
.Y(n_97)
);

CKINVDCx20_ASAP7_75t_R g82 ( 
.A(n_53),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_82),
.B(n_66),
.Y(n_96)
);

INVx4_ASAP7_75t_L g83 ( 
.A(n_60),
.Y(n_83)
);

INVx4_ASAP7_75t_L g99 ( 
.A(n_83),
.Y(n_99)
);

BUFx12f_ASAP7_75t_L g84 ( 
.A(n_54),
.Y(n_84)
);

INVx1_ASAP7_75t_SL g85 ( 
.A(n_84),
.Y(n_85)
);

CKINVDCx20_ASAP7_75t_R g87 ( 
.A(n_79),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_SL g108 ( 
.A(n_87),
.B(n_82),
.Y(n_108)
);

CKINVDCx12_ASAP7_75t_R g88 ( 
.A(n_84),
.Y(n_88)
);

INVxp67_ASAP7_75t_L g116 ( 
.A(n_88),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_SL g100 ( 
.A(n_91),
.B(n_68),
.Y(n_100)
);

AOI22xp33_ASAP7_75t_SL g92 ( 
.A1(n_83),
.A2(n_52),
.B1(n_59),
.B2(n_67),
.Y(n_92)
);

OAI22xp5_ASAP7_75t_L g117 ( 
.A1(n_92),
.A2(n_74),
.B1(n_62),
.B2(n_71),
.Y(n_117)
);

AOI21xp5_ASAP7_75t_L g93 ( 
.A1(n_81),
.A2(n_39),
.B(n_40),
.Y(n_93)
);

OAI21xp33_ASAP7_75t_L g111 ( 
.A1(n_93),
.A2(n_99),
.B(n_89),
.Y(n_111)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_77),
.Y(n_94)
);

INVx1_ASAP7_75t_SL g109 ( 
.A(n_94),
.Y(n_109)
);

OR2x2_ASAP7_75t_L g95 ( 
.A(n_84),
.B(n_68),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_95),
.B(n_96),
.Y(n_101)
);

HB1xp67_ASAP7_75t_L g98 ( 
.A(n_80),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g105 ( 
.A(n_98),
.B(n_69),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_SL g120 ( 
.A(n_100),
.B(n_103),
.Y(n_120)
);

AOI22xp33_ASAP7_75t_L g102 ( 
.A1(n_97),
.A2(n_67),
.B1(n_59),
.B2(n_75),
.Y(n_102)
);

OAI22xp5_ASAP7_75t_SL g132 ( 
.A1(n_102),
.A2(n_114),
.B1(n_115),
.B2(n_70),
.Y(n_132)
);

CKINVDCx20_ASAP7_75t_R g103 ( 
.A(n_95),
.Y(n_103)
);

INVx6_ASAP7_75t_L g104 ( 
.A(n_90),
.Y(n_104)
);

INVx3_ASAP7_75t_L g127 ( 
.A(n_104),
.Y(n_127)
);

AND2x2_ASAP7_75t_L g124 ( 
.A(n_105),
.B(n_111),
.Y(n_124)
);

INVx3_ASAP7_75t_L g106 ( 
.A(n_90),
.Y(n_106)
);

BUFx3_ASAP7_75t_L g136 ( 
.A(n_106),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_L g107 ( 
.A(n_86),
.B(n_93),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_L g121 ( 
.A(n_107),
.B(n_113),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_L g126 ( 
.A(n_108),
.B(n_112),
.Y(n_126)
);

INVx3_ASAP7_75t_L g110 ( 
.A(n_99),
.Y(n_110)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_110),
.Y(n_122)
);

AOI32xp33_ASAP7_75t_L g112 ( 
.A1(n_92),
.A2(n_61),
.A3(n_74),
.B1(n_64),
.B2(n_72),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_L g113 ( 
.A(n_89),
.B(n_61),
.Y(n_113)
);

OAI22xp33_ASAP7_75t_L g114 ( 
.A1(n_85),
.A2(n_75),
.B1(n_56),
.B2(n_58),
.Y(n_114)
);

AOI22xp33_ASAP7_75t_L g115 ( 
.A1(n_85),
.A2(n_56),
.B1(n_58),
.B2(n_72),
.Y(n_115)
);

AOI21xp5_ASAP7_75t_L g131 ( 
.A1(n_117),
.A2(n_1),
.B(n_2),
.Y(n_131)
);

A2O1A1O1Ixp25_ASAP7_75t_L g118 ( 
.A1(n_86),
.A2(n_62),
.B(n_71),
.C(n_64),
.D(n_38),
.Y(n_118)
);

AND2x2_ASAP7_75t_L g128 ( 
.A(n_118),
.B(n_22),
.Y(n_128)
);

BUFx12f_ASAP7_75t_L g119 ( 
.A(n_88),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_L g137 ( 
.A(n_119),
.B(n_4),
.Y(n_137)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_109),
.Y(n_123)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_123),
.Y(n_146)
);

OAI22xp33_ASAP7_75t_SL g125 ( 
.A1(n_111),
.A2(n_70),
.B1(n_73),
.B2(n_65),
.Y(n_125)
);

OAI22xp5_ASAP7_75t_L g149 ( 
.A1(n_125),
.A2(n_129),
.B1(n_131),
.B2(n_134),
.Y(n_149)
);

NOR2xp33_ASAP7_75t_L g142 ( 
.A(n_128),
.B(n_130),
.Y(n_142)
);

OAI22x1_ASAP7_75t_L g129 ( 
.A1(n_102),
.A2(n_70),
.B1(n_63),
.B2(n_21),
.Y(n_129)
);

CKINVDCx20_ASAP7_75t_R g130 ( 
.A(n_101),
.Y(n_130)
);

OR2x2_ASAP7_75t_L g147 ( 
.A(n_132),
.B(n_10),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_SL g133 ( 
.A(n_116),
.B(n_2),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_L g141 ( 
.A(n_133),
.B(n_138),
.Y(n_141)
);

OAI22xp33_ASAP7_75t_SL g134 ( 
.A1(n_115),
.A2(n_23),
.B1(n_50),
.B2(n_48),
.Y(n_134)
);

AOI22xp33_ASAP7_75t_L g135 ( 
.A1(n_119),
.A2(n_3),
.B1(n_4),
.B2(n_5),
.Y(n_135)
);

OAI22xp5_ASAP7_75t_SL g155 ( 
.A1(n_135),
.A2(n_14),
.B1(n_17),
.B2(n_19),
.Y(n_155)
);

INVxp67_ASAP7_75t_L g143 ( 
.A(n_137),
.Y(n_143)
);

NOR2xp33_ASAP7_75t_L g138 ( 
.A(n_119),
.B(n_5),
.Y(n_138)
);

MAJx2_ASAP7_75t_L g139 ( 
.A(n_107),
.B(n_24),
.C(n_47),
.Y(n_139)
);

XOR2xp5_ASAP7_75t_L g144 ( 
.A(n_139),
.B(n_7),
.Y(n_144)
);

NOR2xp33_ASAP7_75t_L g140 ( 
.A(n_108),
.B(n_6),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_L g145 ( 
.A(n_140),
.B(n_8),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_SL g165 ( 
.A(n_144),
.B(n_145),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_L g163 ( 
.A(n_147),
.B(n_154),
.Y(n_163)
);

AND2x6_ASAP7_75t_L g148 ( 
.A(n_125),
.B(n_27),
.Y(n_148)
);

NOR2xp33_ASAP7_75t_L g162 ( 
.A(n_148),
.B(n_150),
.Y(n_162)
);

NOR4xp25_ASAP7_75t_SL g150 ( 
.A(n_126),
.B(n_28),
.C(n_43),
.D(n_36),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_L g151 ( 
.A(n_121),
.B(n_10),
.Y(n_151)
);

NOR2xp33_ASAP7_75t_L g164 ( 
.A(n_151),
.B(n_153),
.Y(n_164)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_122),
.Y(n_152)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_152),
.Y(n_160)
);

OAI21xp5_ASAP7_75t_SL g153 ( 
.A1(n_124),
.A2(n_12),
.B(n_13),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_L g154 ( 
.A(n_120),
.B(n_14),
.Y(n_154)
);

AOI22xp5_ASAP7_75t_L g158 ( 
.A1(n_155),
.A2(n_157),
.B1(n_134),
.B2(n_129),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_L g156 ( 
.A(n_124),
.B(n_32),
.Y(n_156)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_156),
.Y(n_161)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_136),
.Y(n_157)
);

OAI22xp5_ASAP7_75t_SL g167 ( 
.A1(n_158),
.A2(n_159),
.B1(n_147),
.B2(n_143),
.Y(n_167)
);

AOI22xp5_ASAP7_75t_L g159 ( 
.A1(n_149),
.A2(n_127),
.B1(n_135),
.B2(n_136),
.Y(n_159)
);

NOR2xp67_ASAP7_75t_SL g166 ( 
.A(n_163),
.B(n_153),
.Y(n_166)
);

XNOR2xp5_ASAP7_75t_L g170 ( 
.A(n_166),
.B(n_168),
.Y(n_170)
);

AOI22xp5_ASAP7_75t_L g171 ( 
.A1(n_167),
.A2(n_169),
.B1(n_146),
.B2(n_143),
.Y(n_171)
);

XNOR2x2_ASAP7_75t_SL g168 ( 
.A(n_163),
.B(n_141),
.Y(n_168)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_160),
.Y(n_169)
);

AOI22xp5_ASAP7_75t_SL g172 ( 
.A1(n_171),
.A2(n_155),
.B1(n_159),
.B2(n_161),
.Y(n_172)
);

XOR2xp5_ASAP7_75t_L g173 ( 
.A(n_172),
.B(n_158),
.Y(n_173)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_173),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_L g175 ( 
.A(n_174),
.B(n_162),
.Y(n_175)
);

NOR2xp33_ASAP7_75t_L g176 ( 
.A(n_175),
.B(n_170),
.Y(n_176)
);

AO221x1_ASAP7_75t_L g177 ( 
.A1(n_176),
.A2(n_168),
.B1(n_164),
.B2(n_142),
.C(n_165),
.Y(n_177)
);

XNOR2xp5_ASAP7_75t_L g178 ( 
.A(n_177),
.B(n_144),
.Y(n_178)
);

XNOR2xp5_ASAP7_75t_L g179 ( 
.A(n_178),
.B(n_139),
.Y(n_179)
);


endmodule