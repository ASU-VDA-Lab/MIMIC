module fake_jpeg_4777_n_140 (n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_140);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_140;

wire n_117;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_29;
wire n_103;
wire n_50;
wire n_15;
wire n_124;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_30;
wire n_106;
wire n_111;
wire n_24;
wire n_44;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_78;
wire n_20;
wire n_18;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_97;
wire n_135;
wire n_36;
wire n_62;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_96;

BUFx6f_ASAP7_75t_L g13 ( 
.A(n_6),
.Y(n_13)
);

BUFx6f_ASAP7_75t_L g14 ( 
.A(n_11),
.Y(n_14)
);

INVx1_ASAP7_75t_SL g15 ( 
.A(n_11),
.Y(n_15)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_6),
.Y(n_16)
);

BUFx12f_ASAP7_75t_L g17 ( 
.A(n_3),
.Y(n_17)
);

INVx11_ASAP7_75t_L g18 ( 
.A(n_8),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_9),
.Y(n_19)
);

INVx6_ASAP7_75t_SL g20 ( 
.A(n_0),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_5),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_10),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_0),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_7),
.Y(n_24)
);

CKINVDCx14_ASAP7_75t_R g25 ( 
.A(n_9),
.Y(n_25)
);

CKINVDCx5p33_ASAP7_75t_R g26 ( 
.A(n_3),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_0),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_20),
.Y(n_28)
);

INVx6_ASAP7_75t_L g43 ( 
.A(n_28),
.Y(n_43)
);

NAND2xp5_ASAP7_75t_SL g29 ( 
.A(n_23),
.B(n_26),
.Y(n_29)
);

AOI22xp5_ASAP7_75t_SL g38 ( 
.A1(n_29),
.A2(n_30),
.B1(n_25),
.B2(n_16),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_L g30 ( 
.A(n_26),
.B(n_1),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_20),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_31),
.Y(n_47)
);

INVx4_ASAP7_75t_L g32 ( 
.A(n_18),
.Y(n_32)
);

INVx5_ASAP7_75t_L g46 ( 
.A(n_32),
.Y(n_46)
);

INVx8_ASAP7_75t_L g33 ( 
.A(n_13),
.Y(n_33)
);

INVx4_ASAP7_75t_L g37 ( 
.A(n_33),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_13),
.Y(n_34)
);

INVx2_ASAP7_75t_L g45 ( 
.A(n_34),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_13),
.Y(n_35)
);

BUFx8_ASAP7_75t_L g44 ( 
.A(n_35),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_14),
.Y(n_36)
);

BUFx12f_ASAP7_75t_L g42 ( 
.A(n_36),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_38),
.B(n_24),
.Y(n_53)
);

AOI22xp33_ASAP7_75t_L g39 ( 
.A1(n_33),
.A2(n_21),
.B1(n_18),
.B2(n_27),
.Y(n_39)
);

AOI22xp33_ASAP7_75t_SL g49 ( 
.A1(n_39),
.A2(n_40),
.B1(n_25),
.B2(n_16),
.Y(n_49)
);

OAI22xp5_ASAP7_75t_L g40 ( 
.A1(n_33),
.A2(n_21),
.B1(n_27),
.B2(n_18),
.Y(n_40)
);

CKINVDCx5p33_ASAP7_75t_R g41 ( 
.A(n_29),
.Y(n_41)
);

NAND2xp5_ASAP7_75t_SL g50 ( 
.A(n_41),
.B(n_30),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_L g48 ( 
.A(n_38),
.B(n_23),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_L g68 ( 
.A(n_48),
.B(n_59),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_49),
.B(n_54),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_SL g84 ( 
.A(n_50),
.B(n_51),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g51 ( 
.A(n_41),
.B(n_24),
.Y(n_51)
);

BUFx12f_ASAP7_75t_L g52 ( 
.A(n_46),
.Y(n_52)
);

CKINVDCx20_ASAP7_75t_R g81 ( 
.A(n_52),
.Y(n_81)
);

A2O1A1O1Ixp25_ASAP7_75t_L g82 ( 
.A1(n_53),
.A2(n_14),
.B(n_19),
.C(n_4),
.D(n_5),
.Y(n_82)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_46),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_43),
.B(n_31),
.Y(n_55)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_55),
.Y(n_71)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_44),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_56),
.B(n_60),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g57 ( 
.A(n_43),
.B(n_31),
.Y(n_57)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_57),
.Y(n_73)
);

OAI21xp5_ASAP7_75t_L g58 ( 
.A1(n_37),
.A2(n_15),
.B(n_28),
.Y(n_58)
);

AOI21xp5_ASAP7_75t_L g74 ( 
.A1(n_58),
.A2(n_17),
.B(n_14),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_L g59 ( 
.A(n_44),
.B(n_22),
.Y(n_59)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_45),
.Y(n_60)
);

INVx3_ASAP7_75t_L g61 ( 
.A(n_44),
.Y(n_61)
);

INVx5_ASAP7_75t_L g76 ( 
.A(n_61),
.Y(n_76)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_45),
.Y(n_62)
);

INVx4_ASAP7_75t_L g77 ( 
.A(n_62),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_L g63 ( 
.A(n_42),
.B(n_17),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_L g69 ( 
.A(n_63),
.B(n_64),
.Y(n_69)
);

AND2x2_ASAP7_75t_L g64 ( 
.A(n_47),
.B(n_15),
.Y(n_64)
);

MAJIxp5_ASAP7_75t_L g65 ( 
.A(n_37),
.B(n_22),
.C(n_32),
.Y(n_65)
);

MAJIxp5_ASAP7_75t_L g70 ( 
.A(n_65),
.B(n_17),
.C(n_31),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_L g66 ( 
.A(n_42),
.B(n_17),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_L g80 ( 
.A(n_66),
.B(n_42),
.Y(n_80)
);

INVx3_ASAP7_75t_L g67 ( 
.A(n_47),
.Y(n_67)
);

AO22x1_ASAP7_75t_L g72 ( 
.A1(n_67),
.A2(n_35),
.B1(n_36),
.B2(n_34),
.Y(n_72)
);

XNOR2xp5_ASAP7_75t_L g92 ( 
.A(n_70),
.B(n_52),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_72),
.B(n_1),
.Y(n_98)
);

OAI22xp5_ASAP7_75t_L g91 ( 
.A1(n_74),
.A2(n_19),
.B1(n_61),
.B2(n_34),
.Y(n_91)
);

XOR2xp5_ASAP7_75t_L g78 ( 
.A(n_48),
.B(n_32),
.Y(n_78)
);

MAJIxp5_ASAP7_75t_L g87 ( 
.A(n_78),
.B(n_66),
.C(n_64),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_L g94 ( 
.A(n_80),
.B(n_83),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_SL g89 ( 
.A(n_82),
.B(n_64),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g83 ( 
.A(n_63),
.B(n_42),
.Y(n_83)
);

OAI22xp5_ASAP7_75t_SL g85 ( 
.A1(n_75),
.A2(n_65),
.B1(n_58),
.B2(n_67),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_85),
.B(n_93),
.Y(n_104)
);

CKINVDCx20_ASAP7_75t_R g86 ( 
.A(n_79),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_SL g103 ( 
.A(n_86),
.B(n_88),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_L g101 ( 
.A(n_87),
.B(n_94),
.Y(n_101)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_80),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_SL g107 ( 
.A(n_89),
.B(n_90),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_SL g90 ( 
.A(n_68),
.B(n_56),
.Y(n_90)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_91),
.Y(n_99)
);

AND2x2_ASAP7_75t_L g108 ( 
.A(n_92),
.B(n_72),
.Y(n_108)
);

OAI22xp5_ASAP7_75t_SL g93 ( 
.A1(n_69),
.A2(n_36),
.B1(n_35),
.B2(n_19),
.Y(n_93)
);

OAI21xp33_ASAP7_75t_L g95 ( 
.A1(n_69),
.A2(n_1),
.B(n_2),
.Y(n_95)
);

OAI21xp5_ASAP7_75t_SL g102 ( 
.A1(n_95),
.A2(n_74),
.B(n_84),
.Y(n_102)
);

AOI22xp5_ASAP7_75t_L g96 ( 
.A1(n_78),
.A2(n_36),
.B1(n_35),
.B2(n_52),
.Y(n_96)
);

OAI22xp5_ASAP7_75t_SL g100 ( 
.A1(n_96),
.A2(n_70),
.B1(n_68),
.B2(n_71),
.Y(n_100)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_83),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g106 ( 
.A(n_97),
.B(n_98),
.Y(n_106)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_100),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g113 ( 
.A(n_101),
.B(n_105),
.Y(n_113)
);

AOI21xp5_ASAP7_75t_L g115 ( 
.A1(n_102),
.A2(n_87),
.B(n_95),
.Y(n_115)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_94),
.Y(n_105)
);

XNOR2x1_ASAP7_75t_L g117 ( 
.A(n_108),
.B(n_72),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_93),
.B(n_81),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_SL g116 ( 
.A(n_109),
.B(n_82),
.Y(n_116)
);

INVxp67_ASAP7_75t_L g110 ( 
.A(n_104),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_SL g118 ( 
.A(n_110),
.B(n_116),
.Y(n_118)
);

INVx2_ASAP7_75t_L g111 ( 
.A(n_103),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_L g119 ( 
.A(n_111),
.B(n_73),
.Y(n_119)
);

OAI22xp5_ASAP7_75t_L g112 ( 
.A1(n_99),
.A2(n_85),
.B1(n_96),
.B2(n_92),
.Y(n_112)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_112),
.Y(n_120)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_115),
.Y(n_123)
);

AOI32xp33_ASAP7_75t_L g122 ( 
.A1(n_117),
.A2(n_108),
.A3(n_106),
.B1(n_102),
.B2(n_100),
.Y(n_122)
);

AOI21xp5_ASAP7_75t_L g125 ( 
.A1(n_119),
.A2(n_121),
.B(n_110),
.Y(n_125)
);

INVxp67_ASAP7_75t_L g121 ( 
.A(n_117),
.Y(n_121)
);

AOI22xp5_ASAP7_75t_SL g124 ( 
.A1(n_122),
.A2(n_121),
.B1(n_123),
.B2(n_120),
.Y(n_124)
);

OAI21xp5_ASAP7_75t_L g132 ( 
.A1(n_124),
.A2(n_125),
.B(n_76),
.Y(n_132)
);

XNOR2xp5_ASAP7_75t_L g126 ( 
.A(n_118),
.B(n_101),
.Y(n_126)
);

BUFx24_ASAP7_75t_SL g129 ( 
.A(n_126),
.Y(n_129)
);

OAI22xp33_ASAP7_75t_L g127 ( 
.A1(n_121),
.A2(n_113),
.B1(n_108),
.B2(n_114),
.Y(n_127)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_127),
.Y(n_131)
);

AOI22xp5_ASAP7_75t_L g128 ( 
.A1(n_120),
.A2(n_107),
.B1(n_76),
.B2(n_2),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_L g130 ( 
.A(n_128),
.B(n_10),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_SL g134 ( 
.A(n_130),
.B(n_132),
.Y(n_134)
);

AOI21x1_ASAP7_75t_L g133 ( 
.A1(n_131),
.A2(n_127),
.B(n_2),
.Y(n_133)
);

OAI22xp5_ASAP7_75t_SL g137 ( 
.A1(n_133),
.A2(n_12),
.B1(n_77),
.B2(n_134),
.Y(n_137)
);

AOI21xp33_ASAP7_75t_L g135 ( 
.A1(n_129),
.A2(n_4),
.B(n_7),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_L g136 ( 
.A(n_135),
.B(n_8),
.Y(n_136)
);

INVxp67_ASAP7_75t_L g138 ( 
.A(n_136),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_L g139 ( 
.A(n_138),
.B(n_137),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_SL g140 ( 
.A(n_139),
.B(n_137),
.Y(n_140)
);


endmodule