module real_jpeg_16800_n_8 (n_5, n_4, n_0, n_1, n_2, n_6, n_7, n_3, n_8);

input n_5;
input n_4;
input n_0;
input n_1;
input n_2;
input n_6;
input n_7;
input n_3;

output n_8;

wire n_17;
wire n_43;
wire n_37;
wire n_21;
wire n_33;
wire n_35;
wire n_38;
wire n_29;
wire n_10;
wire n_31;
wire n_9;
wire n_12;
wire n_24;
wire n_34;
wire n_44;
wire n_28;
wire n_46;
wire n_23;
wire n_11;
wire n_14;
wire n_45;
wire n_25;
wire n_42;
wire n_22;
wire n_18;
wire n_40;
wire n_39;
wire n_36;
wire n_41;
wire n_26;
wire n_32;
wire n_20;
wire n_19;
wire n_27;
wire n_30;
wire n_16;
wire n_15;
wire n_13;

AOI22xp5_ASAP7_75t_SL g39 ( 
.A1(n_0),
.A2(n_40),
.B1(n_44),
.B2(n_46),
.Y(n_39)
);

INVx5_ASAP7_75t_L g31 ( 
.A(n_1),
.Y(n_31)
);

INVx2_ASAP7_75t_SL g38 ( 
.A(n_1),
.Y(n_38)
);

CKINVDCx6p67_ASAP7_75t_R g45 ( 
.A(n_1),
.Y(n_45)
);

INVx1_ASAP7_75t_L g11 ( 
.A(n_2),
.Y(n_11)
);

NAND2xp5_ASAP7_75t_L g17 ( 
.A(n_2),
.B(n_18),
.Y(n_17)
);

NAND2xp5_ASAP7_75t_L g10 ( 
.A(n_3),
.B(n_11),
.Y(n_10)
);

INVx2_ASAP7_75t_L g18 ( 
.A(n_3),
.Y(n_18)
);

OAI322xp33_ASAP7_75t_L g40 ( 
.A1(n_3),
.A2(n_11),
.A3(n_13),
.B1(n_14),
.B2(n_20),
.C1(n_41),
.C2(n_42),
.Y(n_40)
);

NAND2xp5_ASAP7_75t_SL g41 ( 
.A(n_3),
.B(n_25),
.Y(n_41)
);

AND2x2_ASAP7_75t_SL g43 ( 
.A(n_3),
.B(n_5),
.Y(n_43)
);

INVx2_ASAP7_75t_R g30 ( 
.A(n_4),
.Y(n_30)
);

OR2x4_ASAP7_75t_L g36 ( 
.A(n_4),
.B(n_14),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g22 ( 
.A(n_5),
.B(n_7),
.Y(n_22)
);

INVx2_ASAP7_75t_R g25 ( 
.A(n_5),
.Y(n_25)
);

AOI22xp33_ASAP7_75t_SL g32 ( 
.A1(n_5),
.A2(n_18),
.B1(n_25),
.B2(n_33),
.Y(n_32)
);

AOI221xp5_ASAP7_75t_L g12 ( 
.A1(n_6),
.A2(n_13),
.B1(n_14),
.B2(n_15),
.C(n_16),
.Y(n_12)
);

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_6),
.Y(n_15)
);

INVx2_ASAP7_75t_L g14 ( 
.A(n_7),
.Y(n_14)
);

OAI221xp5_ASAP7_75t_L g8 ( 
.A1(n_9),
.A2(n_31),
.B1(n_32),
.B2(n_34),
.C(n_39),
.Y(n_8)
);

AOI32xp33_ASAP7_75t_SL g9 ( 
.A1(n_10),
.A2(n_12),
.A3(n_19),
.B1(n_26),
.B2(n_29),
.Y(n_9)
);

OAI21xp33_ASAP7_75t_L g26 ( 
.A1(n_10),
.A2(n_25),
.B(n_27),
.Y(n_26)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_10),
.Y(n_33)
);

INVx2_ASAP7_75t_R g13 ( 
.A(n_14),
.Y(n_13)
);

NOR2xp33_ASAP7_75t_R g24 ( 
.A(n_14),
.B(n_25),
.Y(n_24)
);

AND2x4_ASAP7_75t_L g29 ( 
.A(n_14),
.B(n_30),
.Y(n_29)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_17),
.Y(n_16)
);

AND2x2_ASAP7_75t_SL g28 ( 
.A(n_18),
.B(n_25),
.Y(n_28)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_20),
.Y(n_19)
);

NAND2xp5_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_23),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_22),
.Y(n_21)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_24),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_28),
.Y(n_27)
);

NOR2xp33_ASAP7_75t_L g44 ( 
.A(n_30),
.B(n_45),
.Y(n_44)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_35),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_SL g35 ( 
.A(n_36),
.B(n_37),
.Y(n_35)
);

BUFx12f_ASAP7_75t_SL g37 ( 
.A(n_38),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_38),
.Y(n_46)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_43),
.Y(n_42)
);


endmodule