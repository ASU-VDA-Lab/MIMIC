module fake_jpeg_11673_n_82 (n_13, n_21, n_1, n_10, n_6, n_22, n_14, n_19, n_18, n_20, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_82);

input n_13;
input n_21;
input n_1;
input n_10;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_82;

wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_73;
wire n_59;
wire n_65;
wire n_42;
wire n_49;
wire n_76;
wire n_28;
wire n_38;
wire n_26;
wire n_74;
wire n_31;
wire n_29;
wire n_50;
wire n_57;
wire n_23;
wire n_69;
wire n_27;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_30;
wire n_24;
wire n_44;
wire n_25;
wire n_75;
wire n_37;
wire n_70;
wire n_66;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_68;
wire n_52;
wire n_58;
wire n_41;
wire n_60;
wire n_63;
wire n_34;
wire n_39;
wire n_72;
wire n_56;
wire n_79;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_35;
wire n_48;
wire n_46;
wire n_36;
wire n_62;
wire n_43;
wire n_32;

CKINVDCx16_ASAP7_75t_R g23 ( 
.A(n_2),
.Y(n_23)
);

NOR2xp33_ASAP7_75t_L g24 ( 
.A(n_9),
.B(n_10),
.Y(n_24)
);

BUFx8_ASAP7_75t_L g25 ( 
.A(n_22),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_2),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_6),
.Y(n_27)
);

CKINVDCx14_ASAP7_75t_R g28 ( 
.A(n_17),
.Y(n_28)
);

BUFx3_ASAP7_75t_L g29 ( 
.A(n_3),
.Y(n_29)
);

INVx4_ASAP7_75t_L g30 ( 
.A(n_29),
.Y(n_30)
);

INVx4_ASAP7_75t_L g40 ( 
.A(n_30),
.Y(n_40)
);

INVx5_ASAP7_75t_L g31 ( 
.A(n_29),
.Y(n_31)
);

INVx5_ASAP7_75t_L g44 ( 
.A(n_31),
.Y(n_44)
);

BUFx12f_ASAP7_75t_L g32 ( 
.A(n_25),
.Y(n_32)
);

BUFx4f_ASAP7_75t_SL g43 ( 
.A(n_32),
.Y(n_43)
);

BUFx12f_ASAP7_75t_L g33 ( 
.A(n_25),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_33),
.Y(n_39)
);

INVx2_ASAP7_75t_L g34 ( 
.A(n_26),
.Y(n_34)
);

INVx2_ASAP7_75t_L g38 ( 
.A(n_34),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_L g35 ( 
.A(n_27),
.B(n_0),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g37 ( 
.A(n_35),
.B(n_28),
.Y(n_37)
);

CKINVDCx14_ASAP7_75t_R g36 ( 
.A(n_25),
.Y(n_36)
);

OR2x2_ASAP7_75t_L g41 ( 
.A(n_36),
.B(n_23),
.Y(n_41)
);

NAND2xp5_ASAP7_75t_SL g51 ( 
.A(n_37),
.B(n_42),
.Y(n_51)
);

AND2x2_ASAP7_75t_L g50 ( 
.A(n_41),
.B(n_7),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g42 ( 
.A(n_36),
.B(n_28),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g45 ( 
.A(n_41),
.B(n_24),
.Y(n_45)
);

NAND2xp5_ASAP7_75t_L g60 ( 
.A(n_45),
.B(n_49),
.Y(n_60)
);

INVx2_ASAP7_75t_L g46 ( 
.A(n_38),
.Y(n_46)
);

HB1xp67_ASAP7_75t_L g55 ( 
.A(n_46),
.Y(n_55)
);

AOI22xp33_ASAP7_75t_SL g47 ( 
.A1(n_40),
.A2(n_1),
.B1(n_4),
.B2(n_5),
.Y(n_47)
);

XOR2xp5_ASAP7_75t_L g63 ( 
.A(n_47),
.B(n_21),
.Y(n_63)
);

MAJIxp5_ASAP7_75t_R g48 ( 
.A(n_43),
.B(n_5),
.C(n_6),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_48),
.B(n_52),
.Y(n_62)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_43),
.Y(n_49)
);

AND2x2_ASAP7_75t_L g58 ( 
.A(n_50),
.B(n_53),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_L g52 ( 
.A(n_44),
.B(n_8),
.Y(n_52)
);

OAI21xp33_ASAP7_75t_SL g53 ( 
.A1(n_39),
.A2(n_11),
.B(n_12),
.Y(n_53)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_53),
.Y(n_54)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_54),
.Y(n_71)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_51),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_L g66 ( 
.A(n_56),
.B(n_57),
.Y(n_66)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_50),
.Y(n_57)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_46),
.Y(n_59)
);

INVx2_ASAP7_75t_L g69 ( 
.A(n_59),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_51),
.B(n_13),
.Y(n_61)
);

CKINVDCx16_ASAP7_75t_R g68 ( 
.A(n_61),
.Y(n_68)
);

MAJIxp5_ASAP7_75t_L g65 ( 
.A(n_63),
.B(n_64),
.C(n_15),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_51),
.B(n_14),
.Y(n_64)
);

MAJIxp5_ASAP7_75t_L g74 ( 
.A(n_65),
.B(n_67),
.C(n_58),
.Y(n_74)
);

MAJIxp5_ASAP7_75t_L g67 ( 
.A(n_60),
.B(n_16),
.C(n_18),
.Y(n_67)
);

OAI21xp33_ASAP7_75t_L g70 ( 
.A1(n_58),
.A2(n_19),
.B(n_20),
.Y(n_70)
);

CKINVDCx20_ASAP7_75t_R g72 ( 
.A(n_70),
.Y(n_72)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_69),
.Y(n_73)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_73),
.Y(n_77)
);

NOR3xp33_ASAP7_75t_SL g76 ( 
.A(n_74),
.B(n_75),
.C(n_70),
.Y(n_76)
);

CKINVDCx20_ASAP7_75t_R g75 ( 
.A(n_66),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_76),
.B(n_72),
.Y(n_78)
);

MAJIxp5_ASAP7_75t_L g79 ( 
.A(n_78),
.B(n_62),
.C(n_64),
.Y(n_79)
);

MAJIxp5_ASAP7_75t_L g80 ( 
.A(n_79),
.B(n_68),
.C(n_62),
.Y(n_80)
);

MAJIxp5_ASAP7_75t_L g81 ( 
.A(n_80),
.B(n_71),
.C(n_77),
.Y(n_81)
);

XOR2xp5_ASAP7_75t_L g82 ( 
.A(n_81),
.B(n_55),
.Y(n_82)
);


endmodule