module fake_jpeg_28823_n_532 (n_13, n_1, n_10, n_6, n_14, n_18, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_532);

input n_13;
input n_1;
input n_10;
input n_6;
input n_14;
input n_18;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_532;

wire n_529;
wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_525;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_519;
wire n_276;
wire n_143;
wire n_431;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_513;
wire n_283;
wire n_107;
wire n_490;
wire n_517;
wire n_415;
wire n_479;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_48;
wire n_465;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_221;
wire n_256;
wire n_454;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_508;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_393;
wire n_349;
wire n_234;
wire n_530;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_474;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_511;
wire n_305;
wire n_161;
wire n_441;
wire n_342;
wire n_101;
wire n_226;
wire n_509;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_510;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_531;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_523;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_296;
wire n_384;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_491;
wire n_24;
wire n_526;
wire n_467;
wire n_269;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_473;
wire n_45;
wire n_520;
wire n_476;
wire n_337;
wire n_317;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_344;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_481;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_522;
wire n_333;
wire n_518;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_302;
wire n_216;
wire n_528;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_199;
wire n_260;
wire n_413;
wire n_275;
wire n_494;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_492;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_515;
wire n_347;
wire n_521;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_472;
wire n_279;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_484;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_469;
wire n_111;
wire n_197;
wire n_396;
wire n_375;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_527;
wire n_482;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_512;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_516;
wire n_183;
wire n_409;
wire n_249;
wire n_412;
wire n_217;
wire n_471;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_524;
wire n_402;
wire n_504;
wire n_438;
wire n_475;
wire n_247;
wire n_157;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_514;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

INVx2_ASAP7_75t_L g19 ( 
.A(n_10),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_16),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_6),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_13),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_11),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_6),
.Y(n_24)
);

BUFx5_ASAP7_75t_L g25 ( 
.A(n_13),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_4),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_6),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_17),
.Y(n_28)
);

INVx2_ASAP7_75t_L g29 ( 
.A(n_8),
.Y(n_29)
);

NOR2xp33_ASAP7_75t_L g30 ( 
.A(n_17),
.B(n_1),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_16),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_10),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_1),
.Y(n_33)
);

BUFx5_ASAP7_75t_L g34 ( 
.A(n_1),
.Y(n_34)
);

INVx11_ASAP7_75t_L g35 ( 
.A(n_10),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_8),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_10),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_11),
.Y(n_38)
);

INVx13_ASAP7_75t_L g39 ( 
.A(n_16),
.Y(n_39)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_15),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_13),
.Y(n_41)
);

BUFx12_ASAP7_75t_L g42 ( 
.A(n_14),
.Y(n_42)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_17),
.Y(n_43)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_5),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_4),
.Y(n_45)
);

BUFx2_ASAP7_75t_L g46 ( 
.A(n_6),
.Y(n_46)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_7),
.Y(n_47)
);

INVx6_ASAP7_75t_SL g48 ( 
.A(n_14),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_14),
.Y(n_49)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_18),
.Y(n_50)
);

INVx8_ASAP7_75t_L g51 ( 
.A(n_34),
.Y(n_51)
);

INVx8_ASAP7_75t_L g120 ( 
.A(n_51),
.Y(n_120)
);

INVx8_ASAP7_75t_L g52 ( 
.A(n_34),
.Y(n_52)
);

INVx8_ASAP7_75t_L g160 ( 
.A(n_52),
.Y(n_160)
);

INVx2_ASAP7_75t_L g53 ( 
.A(n_19),
.Y(n_53)
);

INVx2_ASAP7_75t_L g102 ( 
.A(n_53),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_30),
.B(n_18),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_54),
.B(n_69),
.Y(n_111)
);

INVx2_ASAP7_75t_L g55 ( 
.A(n_19),
.Y(n_55)
);

INVx2_ASAP7_75t_L g113 ( 
.A(n_55),
.Y(n_113)
);

INVx3_ASAP7_75t_L g56 ( 
.A(n_25),
.Y(n_56)
);

INVx3_ASAP7_75t_L g103 ( 
.A(n_56),
.Y(n_103)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_19),
.Y(n_57)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_57),
.Y(n_110)
);

INVx8_ASAP7_75t_L g58 ( 
.A(n_34),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g112 ( 
.A(n_58),
.Y(n_112)
);

INVx2_ASAP7_75t_L g59 ( 
.A(n_29),
.Y(n_59)
);

INVx2_ASAP7_75t_L g136 ( 
.A(n_59),
.Y(n_136)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_21),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g130 ( 
.A(n_60),
.Y(n_130)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_29),
.Y(n_61)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_61),
.Y(n_122)
);

INVx4_ASAP7_75t_L g62 ( 
.A(n_29),
.Y(n_62)
);

INVx4_ASAP7_75t_L g124 ( 
.A(n_62),
.Y(n_124)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_21),
.Y(n_63)
);

BUFx6f_ASAP7_75t_L g131 ( 
.A(n_63),
.Y(n_131)
);

INVx4_ASAP7_75t_L g64 ( 
.A(n_25),
.Y(n_64)
);

INVx4_ASAP7_75t_L g134 ( 
.A(n_64),
.Y(n_134)
);

INVx8_ASAP7_75t_L g65 ( 
.A(n_25),
.Y(n_65)
);

INVx5_ASAP7_75t_L g104 ( 
.A(n_65),
.Y(n_104)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_21),
.Y(n_66)
);

INVx6_ASAP7_75t_L g135 ( 
.A(n_66),
.Y(n_135)
);

INVx2_ASAP7_75t_L g67 ( 
.A(n_46),
.Y(n_67)
);

INVx2_ASAP7_75t_L g147 ( 
.A(n_67),
.Y(n_147)
);

INVx11_ASAP7_75t_L g68 ( 
.A(n_21),
.Y(n_68)
);

INVx6_ASAP7_75t_L g143 ( 
.A(n_68),
.Y(n_143)
);

CKINVDCx20_ASAP7_75t_R g69 ( 
.A(n_46),
.Y(n_69)
);

BUFx6f_ASAP7_75t_L g70 ( 
.A(n_38),
.Y(n_70)
);

INVx6_ASAP7_75t_L g144 ( 
.A(n_70),
.Y(n_144)
);

INVx3_ASAP7_75t_L g71 ( 
.A(n_39),
.Y(n_71)
);

INVx3_ASAP7_75t_L g107 ( 
.A(n_71),
.Y(n_107)
);

INVx2_ASAP7_75t_L g72 ( 
.A(n_46),
.Y(n_72)
);

INVx2_ASAP7_75t_L g151 ( 
.A(n_72),
.Y(n_151)
);

BUFx6f_ASAP7_75t_L g73 ( 
.A(n_38),
.Y(n_73)
);

INVx6_ASAP7_75t_L g145 ( 
.A(n_73),
.Y(n_145)
);

BUFx6f_ASAP7_75t_L g74 ( 
.A(n_38),
.Y(n_74)
);

INVx6_ASAP7_75t_L g127 ( 
.A(n_74),
.Y(n_127)
);

CKINVDCx20_ASAP7_75t_R g75 ( 
.A(n_46),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g126 ( 
.A(n_75),
.B(n_76),
.Y(n_126)
);

CKINVDCx20_ASAP7_75t_R g76 ( 
.A(n_30),
.Y(n_76)
);

INVx4_ASAP7_75t_L g77 ( 
.A(n_38),
.Y(n_77)
);

INVx3_ASAP7_75t_L g108 ( 
.A(n_77),
.Y(n_108)
);

INVx4_ASAP7_75t_L g78 ( 
.A(n_20),
.Y(n_78)
);

INVx3_ASAP7_75t_L g115 ( 
.A(n_78),
.Y(n_115)
);

BUFx6f_ASAP7_75t_L g79 ( 
.A(n_20),
.Y(n_79)
);

INVx3_ASAP7_75t_SL g114 ( 
.A(n_79),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_SL g80 ( 
.A(n_28),
.B(n_18),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g132 ( 
.A(n_80),
.B(n_87),
.Y(n_132)
);

INVx3_ASAP7_75t_L g81 ( 
.A(n_39),
.Y(n_81)
);

INVx3_ASAP7_75t_L g154 ( 
.A(n_81),
.Y(n_154)
);

BUFx3_ASAP7_75t_L g82 ( 
.A(n_35),
.Y(n_82)
);

INVx5_ASAP7_75t_L g118 ( 
.A(n_82),
.Y(n_118)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_22),
.Y(n_83)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_83),
.Y(n_125)
);

BUFx2_ASAP7_75t_L g84 ( 
.A(n_20),
.Y(n_84)
);

INVx3_ASAP7_75t_L g159 ( 
.A(n_84),
.Y(n_159)
);

BUFx6f_ASAP7_75t_L g85 ( 
.A(n_20),
.Y(n_85)
);

BUFx2_ASAP7_75t_L g129 ( 
.A(n_85),
.Y(n_129)
);

INVx2_ASAP7_75t_L g86 ( 
.A(n_41),
.Y(n_86)
);

INVx2_ASAP7_75t_L g162 ( 
.A(n_86),
.Y(n_162)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_28),
.B(n_15),
.Y(n_87)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_22),
.Y(n_88)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_88),
.Y(n_128)
);

BUFx6f_ASAP7_75t_L g89 ( 
.A(n_41),
.Y(n_89)
);

INVx5_ASAP7_75t_L g119 ( 
.A(n_89),
.Y(n_119)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_22),
.Y(n_90)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_90),
.Y(n_133)
);

INVx8_ASAP7_75t_L g91 ( 
.A(n_41),
.Y(n_91)
);

INVx5_ASAP7_75t_L g149 ( 
.A(n_91),
.Y(n_149)
);

INVx6_ASAP7_75t_L g92 ( 
.A(n_41),
.Y(n_92)
);

INVx5_ASAP7_75t_L g156 ( 
.A(n_92),
.Y(n_156)
);

INVx2_ASAP7_75t_L g93 ( 
.A(n_49),
.Y(n_93)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_93),
.Y(n_137)
);

BUFx10_ASAP7_75t_L g94 ( 
.A(n_48),
.Y(n_94)
);

INVx2_ASAP7_75t_SL g152 ( 
.A(n_94),
.Y(n_152)
);

BUFx6f_ASAP7_75t_L g95 ( 
.A(n_49),
.Y(n_95)
);

INVx5_ASAP7_75t_L g158 ( 
.A(n_95),
.Y(n_158)
);

CKINVDCx16_ASAP7_75t_R g96 ( 
.A(n_48),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g148 ( 
.A(n_96),
.B(n_97),
.Y(n_148)
);

CKINVDCx16_ASAP7_75t_R g97 ( 
.A(n_48),
.Y(n_97)
);

AOI22xp33_ASAP7_75t_SL g98 ( 
.A1(n_49),
.A2(n_32),
.B1(n_44),
.B2(n_37),
.Y(n_98)
);

OAI22xp5_ASAP7_75t_L g116 ( 
.A1(n_98),
.A2(n_32),
.B1(n_37),
.B2(n_44),
.Y(n_116)
);

INVx3_ASAP7_75t_L g99 ( 
.A(n_39),
.Y(n_99)
);

BUFx3_ASAP7_75t_L g117 ( 
.A(n_99),
.Y(n_117)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_31),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_SL g106 ( 
.A(n_100),
.B(n_28),
.Y(n_106)
);

BUFx12_ASAP7_75t_L g101 ( 
.A(n_39),
.Y(n_101)
);

INVx4_ASAP7_75t_SL g105 ( 
.A(n_101),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g168 ( 
.A(n_106),
.B(n_109),
.Y(n_168)
);

CKINVDCx20_ASAP7_75t_R g109 ( 
.A(n_94),
.Y(n_109)
);

AOI22xp5_ASAP7_75t_L g186 ( 
.A1(n_116),
.A2(n_146),
.B1(n_23),
.B2(n_33),
.Y(n_186)
);

AOI22xp33_ASAP7_75t_L g121 ( 
.A1(n_92),
.A2(n_49),
.B1(n_36),
.B2(n_47),
.Y(n_121)
);

OAI22xp5_ASAP7_75t_SL g167 ( 
.A1(n_121),
.A2(n_140),
.B1(n_37),
.B2(n_32),
.Y(n_167)
);

NOR2xp33_ASAP7_75t_SL g123 ( 
.A(n_64),
.B(n_26),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_L g172 ( 
.A(n_123),
.B(n_138),
.Y(n_172)
);

CKINVDCx20_ASAP7_75t_R g138 ( 
.A(n_94),
.Y(n_138)
);

BUFx12f_ASAP7_75t_L g139 ( 
.A(n_101),
.Y(n_139)
);

INVx3_ASAP7_75t_L g195 ( 
.A(n_139),
.Y(n_195)
);

AOI22xp33_ASAP7_75t_L g140 ( 
.A1(n_79),
.A2(n_36),
.B1(n_47),
.B2(n_24),
.Y(n_140)
);

BUFx3_ASAP7_75t_L g141 ( 
.A(n_51),
.Y(n_141)
);

BUFx3_ASAP7_75t_L g198 ( 
.A(n_141),
.Y(n_198)
);

AOI22xp33_ASAP7_75t_SL g142 ( 
.A1(n_84),
.A2(n_50),
.B1(n_31),
.B2(n_43),
.Y(n_142)
);

AOI22xp33_ASAP7_75t_SL g179 ( 
.A1(n_142),
.A2(n_47),
.B1(n_24),
.B2(n_33),
.Y(n_179)
);

OAI22xp5_ASAP7_75t_L g146 ( 
.A1(n_98),
.A2(n_26),
.B1(n_45),
.B2(n_27),
.Y(n_146)
);

BUFx12f_ASAP7_75t_L g150 ( 
.A(n_101),
.Y(n_150)
);

INVx13_ASAP7_75t_L g200 ( 
.A(n_150),
.Y(n_200)
);

BUFx12f_ASAP7_75t_L g153 ( 
.A(n_85),
.Y(n_153)
);

INVx1_ASAP7_75t_SL g213 ( 
.A(n_153),
.Y(n_213)
);

CKINVDCx20_ASAP7_75t_R g155 ( 
.A(n_82),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_L g178 ( 
.A(n_155),
.B(n_71),
.Y(n_178)
);

INVx6_ASAP7_75t_SL g157 ( 
.A(n_89),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_SL g176 ( 
.A(n_157),
.B(n_164),
.Y(n_176)
);

BUFx12f_ASAP7_75t_L g161 ( 
.A(n_95),
.Y(n_161)
);

INVxp67_ASAP7_75t_L g169 ( 
.A(n_161),
.Y(n_169)
);

HAxp5_ASAP7_75t_SL g163 ( 
.A(n_62),
.B(n_44),
.CON(n_163),
.SN(n_163)
);

OR2x4_ASAP7_75t_L g201 ( 
.A(n_163),
.B(n_33),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_SL g164 ( 
.A(n_99),
.B(n_27),
.Y(n_164)
);

NOR2xp33_ASAP7_75t_SL g165 ( 
.A(n_132),
.B(n_45),
.Y(n_165)
);

NOR2xp33_ASAP7_75t_SL g253 ( 
.A(n_165),
.B(n_187),
.Y(n_253)
);

INVx2_ASAP7_75t_L g166 ( 
.A(n_162),
.Y(n_166)
);

INVx2_ASAP7_75t_L g228 ( 
.A(n_166),
.Y(n_228)
);

AOI22xp5_ASAP7_75t_L g233 ( 
.A1(n_167),
.A2(n_206),
.B1(n_135),
.B2(n_144),
.Y(n_233)
);

INVx8_ASAP7_75t_L g170 ( 
.A(n_112),
.Y(n_170)
);

INVx11_ASAP7_75t_L g254 ( 
.A(n_170),
.Y(n_254)
);

NAND2xp5_ASAP7_75t_L g171 ( 
.A(n_125),
.B(n_36),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_L g238 ( 
.A(n_171),
.B(n_173),
.Y(n_238)
);

NAND2xp5_ASAP7_75t_L g173 ( 
.A(n_128),
.B(n_133),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_L g174 ( 
.A(n_111),
.B(n_24),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_L g243 ( 
.A(n_174),
.B(n_184),
.Y(n_243)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_110),
.Y(n_175)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_175),
.Y(n_236)
);

OR2x2_ASAP7_75t_L g177 ( 
.A(n_132),
.B(n_40),
.Y(n_177)
);

CKINVDCx14_ASAP7_75t_R g249 ( 
.A(n_177),
.Y(n_249)
);

NOR2xp33_ASAP7_75t_L g226 ( 
.A(n_178),
.B(n_189),
.Y(n_226)
);

OAI22xp5_ASAP7_75t_L g235 ( 
.A1(n_179),
.A2(n_119),
.B1(n_158),
.B2(n_104),
.Y(n_235)
);

AOI22xp33_ASAP7_75t_SL g180 ( 
.A1(n_163),
.A2(n_50),
.B1(n_43),
.B2(n_40),
.Y(n_180)
);

AOI22xp33_ASAP7_75t_SL g227 ( 
.A1(n_180),
.A2(n_225),
.B1(n_114),
.B2(n_201),
.Y(n_227)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_122),
.Y(n_181)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_181),
.Y(n_251)
);

INVx2_ASAP7_75t_L g182 ( 
.A(n_102),
.Y(n_182)
);

INVx2_ASAP7_75t_L g229 ( 
.A(n_182),
.Y(n_229)
);

BUFx6f_ASAP7_75t_L g183 ( 
.A(n_130),
.Y(n_183)
);

INVx3_ASAP7_75t_SL g275 ( 
.A(n_183),
.Y(n_275)
);

NAND2xp5_ASAP7_75t_L g184 ( 
.A(n_111),
.B(n_23),
.Y(n_184)
);

AOI21xp33_ASAP7_75t_L g185 ( 
.A1(n_126),
.A2(n_40),
.B(n_50),
.Y(n_185)
);

NOR3xp33_ASAP7_75t_L g250 ( 
.A(n_185),
.B(n_161),
.C(n_153),
.Y(n_250)
);

OA22x2_ASAP7_75t_L g259 ( 
.A1(n_186),
.A2(n_222),
.B1(n_224),
.B2(n_0),
.Y(n_259)
);

NAND2xp5_ASAP7_75t_SL g187 ( 
.A(n_126),
.B(n_43),
.Y(n_187)
);

HB1xp67_ASAP7_75t_L g188 ( 
.A(n_108),
.Y(n_188)
);

INVx2_ASAP7_75t_L g240 ( 
.A(n_188),
.Y(n_240)
);

CKINVDCx20_ASAP7_75t_R g189 ( 
.A(n_117),
.Y(n_189)
);

INVx2_ASAP7_75t_L g190 ( 
.A(n_113),
.Y(n_190)
);

INVx2_ASAP7_75t_L g245 ( 
.A(n_190),
.Y(n_245)
);

AND2x4_ASAP7_75t_L g191 ( 
.A(n_142),
.B(n_77),
.Y(n_191)
);

AND2x2_ASAP7_75t_L g248 ( 
.A(n_191),
.B(n_201),
.Y(n_248)
);

NAND2xp5_ASAP7_75t_SL g192 ( 
.A(n_148),
.B(n_31),
.Y(n_192)
);

NOR2xp33_ASAP7_75t_L g230 ( 
.A(n_192),
.B(n_194),
.Y(n_230)
);

NAND2xp5_ASAP7_75t_L g193 ( 
.A(n_136),
.B(n_23),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_L g247 ( 
.A(n_193),
.B(n_203),
.Y(n_247)
);

CKINVDCx12_ASAP7_75t_R g194 ( 
.A(n_105),
.Y(n_194)
);

MAJIxp5_ASAP7_75t_L g196 ( 
.A(n_137),
.B(n_78),
.C(n_52),
.Y(n_196)
);

MAJIxp5_ASAP7_75t_L g244 ( 
.A(n_196),
.B(n_120),
.C(n_160),
.Y(n_244)
);

BUFx12_ASAP7_75t_L g197 ( 
.A(n_118),
.Y(n_197)
);

NOR2xp33_ASAP7_75t_L g232 ( 
.A(n_197),
.B(n_204),
.Y(n_232)
);

INVx2_ASAP7_75t_L g199 ( 
.A(n_147),
.Y(n_199)
);

INVx2_ASAP7_75t_L g262 ( 
.A(n_199),
.Y(n_262)
);

INVx11_ASAP7_75t_L g202 ( 
.A(n_112),
.Y(n_202)
);

INVx6_ASAP7_75t_L g234 ( 
.A(n_202),
.Y(n_234)
);

NAND2xp5_ASAP7_75t_L g203 ( 
.A(n_151),
.B(n_74),
.Y(n_203)
);

OR2x2_ASAP7_75t_L g204 ( 
.A(n_148),
.B(n_42),
.Y(n_204)
);

NAND2xp5_ASAP7_75t_L g205 ( 
.A(n_124),
.B(n_145),
.Y(n_205)
);

NAND2xp5_ASAP7_75t_L g267 ( 
.A(n_205),
.B(n_11),
.Y(n_267)
);

OAI22xp5_ASAP7_75t_L g206 ( 
.A1(n_127),
.A2(n_66),
.B1(n_73),
.B2(n_70),
.Y(n_206)
);

CKINVDCx16_ASAP7_75t_R g207 ( 
.A(n_105),
.Y(n_207)
);

NOR2xp33_ASAP7_75t_L g252 ( 
.A(n_207),
.B(n_210),
.Y(n_252)
);

BUFx6f_ASAP7_75t_L g208 ( 
.A(n_130),
.Y(n_208)
);

BUFx2_ASAP7_75t_L g231 ( 
.A(n_208),
.Y(n_231)
);

INVx2_ASAP7_75t_L g209 ( 
.A(n_115),
.Y(n_209)
);

INVx2_ASAP7_75t_L g270 ( 
.A(n_209),
.Y(n_270)
);

CKINVDCx16_ASAP7_75t_R g210 ( 
.A(n_152),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_SL g211 ( 
.A(n_103),
.B(n_12),
.Y(n_211)
);

NOR2xp33_ASAP7_75t_L g258 ( 
.A(n_211),
.B(n_212),
.Y(n_258)
);

NAND2xp5_ASAP7_75t_SL g212 ( 
.A(n_152),
.B(n_12),
.Y(n_212)
);

NOR2xp33_ASAP7_75t_L g214 ( 
.A(n_154),
.B(n_42),
.Y(n_214)
);

NOR2xp33_ASAP7_75t_L g264 ( 
.A(n_214),
.B(n_216),
.Y(n_264)
);

BUFx6f_ASAP7_75t_L g215 ( 
.A(n_131),
.Y(n_215)
);

INVx3_ASAP7_75t_L g237 ( 
.A(n_215),
.Y(n_237)
);

CKINVDCx16_ASAP7_75t_R g216 ( 
.A(n_139),
.Y(n_216)
);

INVx11_ASAP7_75t_L g217 ( 
.A(n_120),
.Y(n_217)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_217),
.Y(n_271)
);

BUFx6f_ASAP7_75t_L g218 ( 
.A(n_131),
.Y(n_218)
);

INVx3_ASAP7_75t_L g239 ( 
.A(n_218),
.Y(n_239)
);

OR2x2_ASAP7_75t_L g219 ( 
.A(n_140),
.B(n_42),
.Y(n_219)
);

NOR2xp33_ASAP7_75t_L g265 ( 
.A(n_219),
.B(n_220),
.Y(n_265)
);

NAND2xp5_ASAP7_75t_SL g220 ( 
.A(n_107),
.B(n_12),
.Y(n_220)
);

NOR2xp33_ASAP7_75t_L g221 ( 
.A(n_134),
.B(n_150),
.Y(n_221)
);

NOR2xp33_ASAP7_75t_L g268 ( 
.A(n_221),
.B(n_0),
.Y(n_268)
);

AOI22xp5_ASAP7_75t_SL g222 ( 
.A1(n_114),
.A2(n_65),
.B1(n_58),
.B2(n_91),
.Y(n_222)
);

AOI22xp33_ASAP7_75t_L g223 ( 
.A1(n_129),
.A2(n_68),
.B1(n_63),
.B2(n_60),
.Y(n_223)
);

OAI22xp5_ASAP7_75t_SL g261 ( 
.A1(n_223),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_261)
);

AO22x1_ASAP7_75t_SL g224 ( 
.A1(n_121),
.A2(n_42),
.B1(n_35),
.B2(n_2),
.Y(n_224)
);

AOI22xp33_ASAP7_75t_SL g225 ( 
.A1(n_129),
.A2(n_42),
.B1(n_35),
.B2(n_15),
.Y(n_225)
);

INVxp67_ASAP7_75t_L g316 ( 
.A(n_227),
.Y(n_316)
);

OA22x2_ASAP7_75t_L g293 ( 
.A1(n_233),
.A2(n_259),
.B1(n_222),
.B2(n_190),
.Y(n_293)
);

AOI22xp5_ASAP7_75t_L g313 ( 
.A1(n_235),
.A2(n_261),
.B1(n_169),
.B2(n_218),
.Y(n_313)
);

AOI22xp33_ASAP7_75t_L g241 ( 
.A1(n_167),
.A2(n_156),
.B1(n_143),
.B2(n_135),
.Y(n_241)
);

OAI22xp5_ASAP7_75t_SL g277 ( 
.A1(n_241),
.A2(n_256),
.B1(n_263),
.B2(n_272),
.Y(n_277)
);

INVx1_ASAP7_75t_SL g242 ( 
.A(n_175),
.Y(n_242)
);

INVx13_ASAP7_75t_L g288 ( 
.A(n_242),
.Y(n_288)
);

XOR2xp5_ASAP7_75t_L g302 ( 
.A(n_244),
.B(n_217),
.Y(n_302)
);

AOI22xp33_ASAP7_75t_SL g246 ( 
.A1(n_191),
.A2(n_160),
.B1(n_159),
.B2(n_149),
.Y(n_246)
);

AOI22xp33_ASAP7_75t_SL g280 ( 
.A1(n_246),
.A2(n_213),
.B1(n_170),
.B2(n_198),
.Y(n_280)
);

NAND2xp5_ASAP7_75t_SL g292 ( 
.A(n_250),
.B(n_257),
.Y(n_292)
);

NOR2x1_ASAP7_75t_SL g255 ( 
.A(n_204),
.B(n_42),
.Y(n_255)
);

A2O1A1Ixp33_ASAP7_75t_L g321 ( 
.A1(n_255),
.A2(n_200),
.B(n_197),
.C(n_202),
.Y(n_321)
);

AOI22xp33_ASAP7_75t_L g256 ( 
.A1(n_186),
.A2(n_143),
.B1(n_145),
.B2(n_144),
.Y(n_256)
);

CKINVDCx20_ASAP7_75t_R g257 ( 
.A(n_173),
.Y(n_257)
);

HB1xp67_ASAP7_75t_L g260 ( 
.A(n_209),
.Y(n_260)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_260),
.Y(n_278)
);

AOI22xp5_ASAP7_75t_L g263 ( 
.A1(n_191),
.A2(n_219),
.B1(n_224),
.B2(n_206),
.Y(n_263)
);

AOI22xp5_ASAP7_75t_SL g266 ( 
.A1(n_191),
.A2(n_0),
.B1(n_2),
.B2(n_3),
.Y(n_266)
);

OAI21xp5_ASAP7_75t_L g307 ( 
.A1(n_266),
.A2(n_213),
.B(n_169),
.Y(n_307)
);

NAND2xp5_ASAP7_75t_L g295 ( 
.A(n_267),
.B(n_276),
.Y(n_295)
);

NOR2xp33_ASAP7_75t_L g279 ( 
.A(n_268),
.B(n_269),
.Y(n_279)
);

NOR2xp33_ASAP7_75t_L g269 ( 
.A(n_168),
.B(n_172),
.Y(n_269)
);

AOI22xp5_ASAP7_75t_L g272 ( 
.A1(n_224),
.A2(n_2),
.B1(n_3),
.B2(n_4),
.Y(n_272)
);

INVx1_ASAP7_75t_SL g273 ( 
.A(n_181),
.Y(n_273)
);

INVx13_ASAP7_75t_L g301 ( 
.A(n_273),
.Y(n_301)
);

AOI22xp5_ASAP7_75t_L g274 ( 
.A1(n_176),
.A2(n_11),
.B1(n_4),
.B2(n_5),
.Y(n_274)
);

OAI22xp5_ASAP7_75t_L g284 ( 
.A1(n_274),
.A2(n_184),
.B1(n_174),
.B2(n_177),
.Y(n_284)
);

NAND2xp5_ASAP7_75t_L g276 ( 
.A(n_171),
.B(n_193),
.Y(n_276)
);

INVxp67_ASAP7_75t_L g326 ( 
.A(n_280),
.Y(n_326)
);

CKINVDCx20_ASAP7_75t_R g281 ( 
.A(n_226),
.Y(n_281)
);

NAND2xp5_ASAP7_75t_SL g328 ( 
.A(n_281),
.B(n_286),
.Y(n_328)
);

OAI21xp5_ASAP7_75t_SL g282 ( 
.A1(n_248),
.A2(n_196),
.B(n_205),
.Y(n_282)
);

OAI21xp5_ASAP7_75t_SL g340 ( 
.A1(n_282),
.A2(n_321),
.B(n_238),
.Y(n_340)
);

INVx2_ASAP7_75t_L g283 ( 
.A(n_270),
.Y(n_283)
);

INVx2_ASAP7_75t_L g323 ( 
.A(n_283),
.Y(n_323)
);

AOI22xp5_ASAP7_75t_L g333 ( 
.A1(n_284),
.A2(n_265),
.B1(n_232),
.B2(n_248),
.Y(n_333)
);

BUFx4f_ASAP7_75t_SL g285 ( 
.A(n_275),
.Y(n_285)
);

INVxp67_ASAP7_75t_L g362 ( 
.A(n_285),
.Y(n_362)
);

CKINVDCx16_ASAP7_75t_R g286 ( 
.A(n_252),
.Y(n_286)
);

NOR2xp33_ASAP7_75t_L g287 ( 
.A(n_253),
.B(n_165),
.Y(n_287)
);

NOR2xp33_ASAP7_75t_SL g352 ( 
.A(n_287),
.B(n_291),
.Y(n_352)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_236),
.Y(n_289)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_289),
.Y(n_332)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_236),
.Y(n_290)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_290),
.Y(n_337)
);

NOR2xp33_ASAP7_75t_L g291 ( 
.A(n_253),
.B(n_189),
.Y(n_291)
);

AND2x2_ASAP7_75t_L g330 ( 
.A(n_293),
.B(n_307),
.Y(n_330)
);

BUFx3_ASAP7_75t_L g294 ( 
.A(n_254),
.Y(n_294)
);

INVx2_ASAP7_75t_L g324 ( 
.A(n_294),
.Y(n_324)
);

NOR2xp33_ASAP7_75t_L g296 ( 
.A(n_230),
.B(n_210),
.Y(n_296)
);

NOR2xp33_ASAP7_75t_L g325 ( 
.A(n_296),
.B(n_297),
.Y(n_325)
);

NOR2xp33_ASAP7_75t_L g297 ( 
.A(n_257),
.B(n_207),
.Y(n_297)
);

INVx2_ASAP7_75t_L g298 ( 
.A(n_270),
.Y(n_298)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_298),
.Y(n_336)
);

INVx2_ASAP7_75t_L g299 ( 
.A(n_228),
.Y(n_299)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_299),
.Y(n_341)
);

NOR2xp33_ASAP7_75t_SL g300 ( 
.A(n_249),
.B(n_203),
.Y(n_300)
);

NAND3xp33_ASAP7_75t_L g342 ( 
.A(n_300),
.B(n_305),
.C(n_317),
.Y(n_342)
);

XNOR2xp5_ASAP7_75t_SL g351 ( 
.A(n_302),
.B(n_320),
.Y(n_351)
);

INVx3_ASAP7_75t_L g303 ( 
.A(n_234),
.Y(n_303)
);

INVx1_ASAP7_75t_L g345 ( 
.A(n_303),
.Y(n_345)
);

NOR2xp33_ASAP7_75t_L g304 ( 
.A(n_243),
.B(n_216),
.Y(n_304)
);

NOR2xp33_ASAP7_75t_L g349 ( 
.A(n_304),
.B(n_311),
.Y(n_349)
);

NOR2xp33_ASAP7_75t_SL g305 ( 
.A(n_243),
.B(n_182),
.Y(n_305)
);

NAND2xp5_ASAP7_75t_L g306 ( 
.A(n_276),
.B(n_199),
.Y(n_306)
);

NAND2xp5_ASAP7_75t_L g329 ( 
.A(n_306),
.B(n_315),
.Y(n_329)
);

AOI22xp33_ASAP7_75t_SL g308 ( 
.A1(n_255),
.A2(n_235),
.B1(n_259),
.B2(n_198),
.Y(n_308)
);

AOI22xp33_ASAP7_75t_SL g359 ( 
.A1(n_308),
.A2(n_312),
.B1(n_314),
.B2(n_231),
.Y(n_359)
);

CKINVDCx10_ASAP7_75t_R g309 ( 
.A(n_275),
.Y(n_309)
);

CKINVDCx16_ASAP7_75t_R g331 ( 
.A(n_309),
.Y(n_331)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_251),
.Y(n_310)
);

INVx1_ASAP7_75t_L g358 ( 
.A(n_310),
.Y(n_358)
);

INVx3_ASAP7_75t_L g311 ( 
.A(n_234),
.Y(n_311)
);

INVx3_ASAP7_75t_L g312 ( 
.A(n_237),
.Y(n_312)
);

OAI22xp5_ASAP7_75t_L g348 ( 
.A1(n_313),
.A2(n_275),
.B1(n_208),
.B2(n_239),
.Y(n_348)
);

INVx13_ASAP7_75t_L g314 ( 
.A(n_237),
.Y(n_314)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_251),
.Y(n_315)
);

NOR2xp33_ASAP7_75t_L g317 ( 
.A(n_264),
.B(n_195),
.Y(n_317)
);

NAND2xp5_ASAP7_75t_L g318 ( 
.A(n_247),
.B(n_166),
.Y(n_318)
);

NAND2xp5_ASAP7_75t_L g338 ( 
.A(n_318),
.B(n_320),
.Y(n_338)
);

AOI22xp5_ASAP7_75t_L g319 ( 
.A1(n_248),
.A2(n_215),
.B1(n_208),
.B2(n_183),
.Y(n_319)
);

OAI22xp5_ASAP7_75t_SL g327 ( 
.A1(n_319),
.A2(n_233),
.B1(n_263),
.B2(n_244),
.Y(n_327)
);

NAND2xp5_ASAP7_75t_L g320 ( 
.A(n_247),
.B(n_215),
.Y(n_320)
);

NAND2xp5_ASAP7_75t_L g322 ( 
.A(n_238),
.B(n_183),
.Y(n_322)
);

NAND2xp5_ASAP7_75t_L g339 ( 
.A(n_322),
.B(n_267),
.Y(n_339)
);

AOI22xp5_ASAP7_75t_L g378 ( 
.A1(n_327),
.A2(n_347),
.B1(n_348),
.B2(n_354),
.Y(n_378)
);

NAND2xp5_ASAP7_75t_SL g392 ( 
.A(n_333),
.B(n_356),
.Y(n_392)
);

MAJIxp5_ASAP7_75t_L g334 ( 
.A(n_302),
.B(n_282),
.C(n_295),
.Y(n_334)
);

MAJIxp5_ASAP7_75t_L g370 ( 
.A(n_334),
.B(n_344),
.C(n_351),
.Y(n_370)
);

MAJIxp5_ASAP7_75t_SL g335 ( 
.A(n_292),
.B(n_266),
.C(n_259),
.Y(n_335)
);

AOI21xp33_ASAP7_75t_L g393 ( 
.A1(n_335),
.A2(n_342),
.B(n_356),
.Y(n_393)
);

NAND2xp5_ASAP7_75t_L g368 ( 
.A(n_339),
.B(n_355),
.Y(n_368)
);

XNOR2xp5_ASAP7_75t_SL g387 ( 
.A(n_340),
.B(n_343),
.Y(n_387)
);

XOR2x1_ASAP7_75t_L g343 ( 
.A(n_300),
.B(n_259),
.Y(n_343)
);

MAJx2_ASAP7_75t_L g344 ( 
.A(n_295),
.B(n_258),
.C(n_273),
.Y(n_344)
);

OAI32xp33_ASAP7_75t_L g346 ( 
.A1(n_306),
.A2(n_272),
.A3(n_274),
.B1(n_271),
.B2(n_261),
.Y(n_346)
);

INVx1_ASAP7_75t_L g372 ( 
.A(n_346),
.Y(n_372)
);

OAI22xp5_ASAP7_75t_SL g347 ( 
.A1(n_316),
.A2(n_242),
.B1(n_271),
.B2(n_218),
.Y(n_347)
);

AOI22xp5_ASAP7_75t_L g350 ( 
.A1(n_277),
.A2(n_240),
.B1(n_239),
.B2(n_262),
.Y(n_350)
);

OAI22xp5_ASAP7_75t_SL g367 ( 
.A1(n_350),
.A2(n_353),
.B1(n_361),
.B2(n_313),
.Y(n_367)
);

AOI22xp5_ASAP7_75t_L g353 ( 
.A1(n_277),
.A2(n_240),
.B1(n_228),
.B2(n_245),
.Y(n_353)
);

OAI22xp5_ASAP7_75t_SL g354 ( 
.A1(n_316),
.A2(n_231),
.B1(n_254),
.B2(n_262),
.Y(n_354)
);

NAND2xp5_ASAP7_75t_L g355 ( 
.A(n_322),
.B(n_245),
.Y(n_355)
);

OAI21xp5_ASAP7_75t_SL g356 ( 
.A1(n_321),
.A2(n_229),
.B(n_195),
.Y(n_356)
);

NAND2xp5_ASAP7_75t_L g357 ( 
.A(n_318),
.B(n_229),
.Y(n_357)
);

NAND2xp5_ASAP7_75t_L g377 ( 
.A(n_357),
.B(n_360),
.Y(n_377)
);

AOI22xp33_ASAP7_75t_SL g363 ( 
.A1(n_359),
.A2(n_309),
.B1(n_294),
.B2(n_312),
.Y(n_363)
);

NAND2xp5_ASAP7_75t_L g360 ( 
.A(n_305),
.B(n_231),
.Y(n_360)
);

AOI22xp5_ASAP7_75t_L g361 ( 
.A1(n_293),
.A2(n_197),
.B1(n_5),
.B2(n_7),
.Y(n_361)
);

OAI22xp5_ASAP7_75t_L g399 ( 
.A1(n_363),
.A2(n_393),
.B1(n_326),
.B2(n_362),
.Y(n_399)
);

AND2x2_ASAP7_75t_L g364 ( 
.A(n_330),
.B(n_293),
.Y(n_364)
);

AO21x1_ASAP7_75t_L g407 ( 
.A1(n_364),
.A2(n_382),
.B(n_391),
.Y(n_407)
);

NOR2xp33_ASAP7_75t_L g365 ( 
.A(n_352),
.B(n_281),
.Y(n_365)
);

INVx1_ASAP7_75t_L g401 ( 
.A(n_365),
.Y(n_401)
);

CKINVDCx16_ASAP7_75t_R g366 ( 
.A(n_328),
.Y(n_366)
);

NOR2xp33_ASAP7_75t_L g400 ( 
.A(n_366),
.B(n_369),
.Y(n_400)
);

AOI22xp5_ASAP7_75t_L g398 ( 
.A1(n_367),
.A2(n_381),
.B1(n_327),
.B2(n_347),
.Y(n_398)
);

INVxp67_ASAP7_75t_SL g369 ( 
.A(n_360),
.Y(n_369)
);

OAI21xp33_ASAP7_75t_L g371 ( 
.A1(n_335),
.A2(n_286),
.B(n_279),
.Y(n_371)
);

AOI22xp5_ASAP7_75t_SL g418 ( 
.A1(n_371),
.A2(n_324),
.B1(n_336),
.B2(n_341),
.Y(n_418)
);

NOR2x1_ASAP7_75t_L g373 ( 
.A(n_333),
.B(n_319),
.Y(n_373)
);

NAND2xp5_ASAP7_75t_L g423 ( 
.A(n_373),
.B(n_396),
.Y(n_423)
);

CKINVDCx16_ASAP7_75t_R g374 ( 
.A(n_332),
.Y(n_374)
);

NOR2xp33_ASAP7_75t_L g402 ( 
.A(n_374),
.B(n_389),
.Y(n_402)
);

HB1xp67_ASAP7_75t_L g375 ( 
.A(n_324),
.Y(n_375)
);

INVx1_ASAP7_75t_L g415 ( 
.A(n_375),
.Y(n_415)
);

INVx1_ASAP7_75t_L g376 ( 
.A(n_355),
.Y(n_376)
);

INVx1_ASAP7_75t_L g417 ( 
.A(n_376),
.Y(n_417)
);

CKINVDCx20_ASAP7_75t_R g379 ( 
.A(n_357),
.Y(n_379)
);

CKINVDCx20_ASAP7_75t_R g421 ( 
.A(n_379),
.Y(n_421)
);

INVx2_ASAP7_75t_L g380 ( 
.A(n_323),
.Y(n_380)
);

INVx2_ASAP7_75t_L g425 ( 
.A(n_380),
.Y(n_425)
);

OAI22xp5_ASAP7_75t_SL g381 ( 
.A1(n_361),
.A2(n_293),
.B1(n_307),
.B2(n_315),
.Y(n_381)
);

AND2x2_ASAP7_75t_L g382 ( 
.A(n_330),
.B(n_289),
.Y(n_382)
);

MAJIxp5_ASAP7_75t_L g383 ( 
.A(n_334),
.B(n_278),
.C(n_284),
.Y(n_383)
);

MAJIxp5_ASAP7_75t_L g403 ( 
.A(n_383),
.B(n_388),
.C(n_370),
.Y(n_403)
);

NAND2xp5_ASAP7_75t_L g384 ( 
.A(n_339),
.B(n_290),
.Y(n_384)
);

INVx1_ASAP7_75t_L g397 ( 
.A(n_384),
.Y(n_397)
);

OAI32xp33_ASAP7_75t_L g385 ( 
.A1(n_343),
.A2(n_310),
.A3(n_278),
.B1(n_283),
.B2(n_298),
.Y(n_385)
);

INVx1_ASAP7_75t_L g411 ( 
.A(n_385),
.Y(n_411)
);

NAND2xp5_ASAP7_75t_L g386 ( 
.A(n_338),
.B(n_329),
.Y(n_386)
);

INVx1_ASAP7_75t_L g424 ( 
.A(n_386),
.Y(n_424)
);

MAJIxp5_ASAP7_75t_L g388 ( 
.A(n_351),
.B(n_311),
.C(n_303),
.Y(n_388)
);

CKINVDCx16_ASAP7_75t_R g389 ( 
.A(n_337),
.Y(n_389)
);

NAND3xp33_ASAP7_75t_L g390 ( 
.A(n_325),
.B(n_288),
.C(n_301),
.Y(n_390)
);

NOR2xp33_ASAP7_75t_L g405 ( 
.A(n_390),
.B(n_394),
.Y(n_405)
);

OAI21xp5_ASAP7_75t_L g391 ( 
.A1(n_330),
.A2(n_285),
.B(n_301),
.Y(n_391)
);

NOR2xp33_ASAP7_75t_L g394 ( 
.A(n_349),
.B(n_299),
.Y(n_394)
);

INVx1_ASAP7_75t_L g395 ( 
.A(n_358),
.Y(n_395)
);

INVx2_ASAP7_75t_L g426 ( 
.A(n_395),
.Y(n_426)
);

CKINVDCx20_ASAP7_75t_R g396 ( 
.A(n_329),
.Y(n_396)
);

OAI22xp5_ASAP7_75t_SL g432 ( 
.A1(n_398),
.A2(n_409),
.B1(n_413),
.B2(n_376),
.Y(n_432)
);

AOI22xp33_ASAP7_75t_L g445 ( 
.A1(n_399),
.A2(n_367),
.B1(n_373),
.B2(n_395),
.Y(n_445)
);

MAJIxp5_ASAP7_75t_L g442 ( 
.A(n_403),
.B(n_420),
.C(n_389),
.Y(n_442)
);

FAx1_ASAP7_75t_SL g404 ( 
.A(n_387),
.B(n_338),
.CI(n_340),
.CON(n_404),
.SN(n_404)
);

NAND2xp5_ASAP7_75t_L g431 ( 
.A(n_404),
.B(n_364),
.Y(n_431)
);

XNOR2xp5_ASAP7_75t_SL g406 ( 
.A(n_370),
.B(n_344),
.Y(n_406)
);

XNOR2xp5_ASAP7_75t_SL g437 ( 
.A(n_406),
.B(n_408),
.Y(n_437)
);

XNOR2xp5_ASAP7_75t_SL g408 ( 
.A(n_387),
.B(n_383),
.Y(n_408)
);

AOI22xp5_ASAP7_75t_L g409 ( 
.A1(n_372),
.A2(n_326),
.B1(n_346),
.B2(n_354),
.Y(n_409)
);

NOR2xp33_ASAP7_75t_SL g410 ( 
.A(n_396),
.B(n_331),
.Y(n_410)
);

CKINVDCx14_ASAP7_75t_R g444 ( 
.A(n_410),
.Y(n_444)
);

INVx3_ASAP7_75t_L g412 ( 
.A(n_380),
.Y(n_412)
);

INVx2_ASAP7_75t_L g439 ( 
.A(n_412),
.Y(n_439)
);

AOI22xp5_ASAP7_75t_L g413 ( 
.A1(n_372),
.A2(n_350),
.B1(n_353),
.B2(n_362),
.Y(n_413)
);

XOR2xp5_ASAP7_75t_L g414 ( 
.A(n_388),
.B(n_345),
.Y(n_414)
);

XOR2xp5_ASAP7_75t_L g436 ( 
.A(n_414),
.B(n_381),
.Y(n_436)
);

XNOR2xp5_ASAP7_75t_SL g416 ( 
.A(n_392),
.B(n_288),
.Y(n_416)
);

XNOR2xp5_ASAP7_75t_SL g443 ( 
.A(n_416),
.B(n_377),
.Y(n_443)
);

OAI22xp5_ASAP7_75t_L g430 ( 
.A1(n_418),
.A2(n_391),
.B1(n_378),
.B2(n_382),
.Y(n_430)
);

OAI22xp5_ASAP7_75t_L g419 ( 
.A1(n_378),
.A2(n_336),
.B1(n_323),
.B2(n_285),
.Y(n_419)
);

INVx1_ASAP7_75t_L g427 ( 
.A(n_419),
.Y(n_427)
);

MAJIxp5_ASAP7_75t_L g420 ( 
.A(n_384),
.B(n_314),
.C(n_197),
.Y(n_420)
);

INVxp67_ASAP7_75t_SL g422 ( 
.A(n_377),
.Y(n_422)
);

NOR2xp33_ASAP7_75t_L g440 ( 
.A(n_422),
.B(n_400),
.Y(n_440)
);

INVx1_ASAP7_75t_L g428 ( 
.A(n_401),
.Y(n_428)
);

INVx1_ASAP7_75t_L g456 ( 
.A(n_428),
.Y(n_456)
);

OAI21xp5_ASAP7_75t_L g429 ( 
.A1(n_423),
.A2(n_364),
.B(n_382),
.Y(n_429)
);

NAND2xp5_ASAP7_75t_L g454 ( 
.A(n_429),
.B(n_407),
.Y(n_454)
);

AOI22xp5_ASAP7_75t_L g470 ( 
.A1(n_430),
.A2(n_432),
.B1(n_446),
.B2(n_450),
.Y(n_470)
);

NAND2xp5_ASAP7_75t_SL g462 ( 
.A(n_431),
.B(n_447),
.Y(n_462)
);

NAND2xp5_ASAP7_75t_L g433 ( 
.A(n_421),
.B(n_379),
.Y(n_433)
);

INVx1_ASAP7_75t_L g464 ( 
.A(n_433),
.Y(n_464)
);

OAI22xp5_ASAP7_75t_L g434 ( 
.A1(n_411),
.A2(n_398),
.B1(n_405),
.B2(n_409),
.Y(n_434)
);

INVx1_ASAP7_75t_L g467 ( 
.A(n_434),
.Y(n_467)
);

XOR2x2_ASAP7_75t_SL g435 ( 
.A(n_404),
.B(n_385),
.Y(n_435)
);

XNOR2xp5_ASAP7_75t_L g459 ( 
.A(n_435),
.B(n_448),
.Y(n_459)
);

XOR2xp5_ASAP7_75t_L g458 ( 
.A(n_436),
.B(n_441),
.Y(n_458)
);

XNOR2x2_ASAP7_75t_SL g438 ( 
.A(n_423),
.B(n_386),
.Y(n_438)
);

OAI22xp5_ASAP7_75t_L g453 ( 
.A1(n_438),
.A2(n_445),
.B1(n_418),
.B2(n_417),
.Y(n_453)
);

INVx1_ASAP7_75t_L g469 ( 
.A(n_440),
.Y(n_469)
);

XOR2xp5_ASAP7_75t_L g441 ( 
.A(n_403),
.B(n_368),
.Y(n_441)
);

MAJIxp5_ASAP7_75t_L g455 ( 
.A(n_442),
.B(n_408),
.C(n_406),
.Y(n_455)
);

XOR2xp5_ASAP7_75t_L g465 ( 
.A(n_443),
.B(n_407),
.Y(n_465)
);

OAI22xp5_ASAP7_75t_SL g446 ( 
.A1(n_411),
.A2(n_413),
.B1(n_397),
.B2(n_424),
.Y(n_446)
);

NOR2xp33_ASAP7_75t_SL g447 ( 
.A(n_402),
.B(n_368),
.Y(n_447)
);

XNOR2xp5_ASAP7_75t_L g448 ( 
.A(n_414),
.B(n_200),
.Y(n_448)
);

INVx1_ASAP7_75t_L g449 ( 
.A(n_426),
.Y(n_449)
);

INVx1_ASAP7_75t_L g471 ( 
.A(n_449),
.Y(n_471)
);

OAI22xp5_ASAP7_75t_SL g450 ( 
.A1(n_397),
.A2(n_285),
.B1(n_5),
.B2(n_7),
.Y(n_450)
);

NAND2xp5_ASAP7_75t_L g451 ( 
.A(n_424),
.B(n_3),
.Y(n_451)
);

INVx1_ASAP7_75t_L g472 ( 
.A(n_451),
.Y(n_472)
);

NOR2xp33_ASAP7_75t_L g452 ( 
.A(n_420),
.B(n_3),
.Y(n_452)
);

CKINVDCx16_ASAP7_75t_R g457 ( 
.A(n_452),
.Y(n_457)
);

XNOR2xp5_ASAP7_75t_SL g477 ( 
.A(n_453),
.B(n_454),
.Y(n_477)
);

MAJIxp5_ASAP7_75t_L g475 ( 
.A(n_455),
.B(n_463),
.C(n_466),
.Y(n_475)
);

NAND2xp5_ASAP7_75t_L g460 ( 
.A(n_433),
.B(n_426),
.Y(n_460)
);

INVx1_ASAP7_75t_L g482 ( 
.A(n_460),
.Y(n_482)
);

XNOR2xp5_ASAP7_75t_L g461 ( 
.A(n_436),
.B(n_416),
.Y(n_461)
);

XNOR2xp5_ASAP7_75t_L g485 ( 
.A(n_461),
.B(n_465),
.Y(n_485)
);

MAJIxp5_ASAP7_75t_L g463 ( 
.A(n_441),
.B(n_404),
.C(n_415),
.Y(n_463)
);

MAJIxp5_ASAP7_75t_L g466 ( 
.A(n_442),
.B(n_425),
.C(n_412),
.Y(n_466)
);

HB1xp67_ASAP7_75t_L g468 ( 
.A(n_439),
.Y(n_468)
);

INVx1_ASAP7_75t_L g483 ( 
.A(n_468),
.Y(n_483)
);

INVx1_ASAP7_75t_L g473 ( 
.A(n_451),
.Y(n_473)
);

INVx1_ASAP7_75t_L g487 ( 
.A(n_473),
.Y(n_487)
);

CKINVDCx20_ASAP7_75t_R g474 ( 
.A(n_460),
.Y(n_474)
);

NAND2xp5_ASAP7_75t_SL g503 ( 
.A(n_474),
.B(n_480),
.Y(n_503)
);

NOR3xp33_ASAP7_75t_SL g476 ( 
.A(n_462),
.B(n_435),
.C(n_444),
.Y(n_476)
);

CKINVDCx20_ASAP7_75t_R g500 ( 
.A(n_476),
.Y(n_500)
);

AOI22xp5_ASAP7_75t_L g478 ( 
.A1(n_467),
.A2(n_432),
.B1(n_427),
.B2(n_446),
.Y(n_478)
);

INVx1_ASAP7_75t_L g497 ( 
.A(n_478),
.Y(n_497)
);

NAND2xp5_ASAP7_75t_L g479 ( 
.A(n_464),
.B(n_450),
.Y(n_479)
);

CKINVDCx14_ASAP7_75t_R g499 ( 
.A(n_479),
.Y(n_499)
);

OAI22xp5_ASAP7_75t_SL g480 ( 
.A1(n_470),
.A2(n_454),
.B1(n_429),
.B2(n_431),
.Y(n_480)
);

AOI21xp5_ASAP7_75t_L g481 ( 
.A1(n_470),
.A2(n_438),
.B(n_448),
.Y(n_481)
);

OAI21xp5_ASAP7_75t_SL g492 ( 
.A1(n_481),
.A2(n_463),
.B(n_465),
.Y(n_492)
);

INVx1_ASAP7_75t_L g484 ( 
.A(n_456),
.Y(n_484)
);

AOI22xp33_ASAP7_75t_SL g496 ( 
.A1(n_484),
.A2(n_482),
.B1(n_487),
.B2(n_483),
.Y(n_496)
);

NAND2xp5_ASAP7_75t_L g486 ( 
.A(n_473),
.B(n_425),
.Y(n_486)
);

NOR2xp33_ASAP7_75t_L g495 ( 
.A(n_486),
.B(n_488),
.Y(n_495)
);

NAND2xp5_ASAP7_75t_SL g488 ( 
.A(n_469),
.B(n_439),
.Y(n_488)
);

MAJIxp5_ASAP7_75t_L g489 ( 
.A(n_466),
.B(n_437),
.C(n_443),
.Y(n_489)
);

MAJIxp5_ASAP7_75t_L g498 ( 
.A(n_489),
.B(n_458),
.C(n_455),
.Y(n_498)
);

NOR2xp33_ASAP7_75t_SL g490 ( 
.A(n_457),
.B(n_437),
.Y(n_490)
);

NOR2xp33_ASAP7_75t_L g501 ( 
.A(n_490),
.B(n_459),
.Y(n_501)
);

XOR2xp5_ASAP7_75t_L g491 ( 
.A(n_485),
.B(n_458),
.Y(n_491)
);

MAJIxp5_ASAP7_75t_L g505 ( 
.A(n_491),
.B(n_498),
.C(n_502),
.Y(n_505)
);

INVx1_ASAP7_75t_L g507 ( 
.A(n_492),
.Y(n_507)
);

OAI21xp5_ASAP7_75t_L g493 ( 
.A1(n_481),
.A2(n_472),
.B(n_471),
.Y(n_493)
);

AND2x2_ASAP7_75t_L g512 ( 
.A(n_493),
.B(n_475),
.Y(n_512)
);

BUFx24_ASAP7_75t_SL g494 ( 
.A(n_478),
.Y(n_494)
);

NOR2xp33_ASAP7_75t_SL g514 ( 
.A(n_494),
.B(n_504),
.Y(n_514)
);

INVx1_ASAP7_75t_L g508 ( 
.A(n_496),
.Y(n_508)
);

INVx1_ASAP7_75t_L g510 ( 
.A(n_501),
.Y(n_510)
);

XOR2xp5_ASAP7_75t_L g502 ( 
.A(n_485),
.B(n_461),
.Y(n_502)
);

NOR2xp33_ASAP7_75t_L g504 ( 
.A(n_480),
.B(n_459),
.Y(n_504)
);

AOI22xp5_ASAP7_75t_L g506 ( 
.A1(n_503),
.A2(n_476),
.B1(n_477),
.B2(n_479),
.Y(n_506)
);

INVxp67_ASAP7_75t_L g517 ( 
.A(n_506),
.Y(n_517)
);

AOI22xp5_ASAP7_75t_L g509 ( 
.A1(n_499),
.A2(n_477),
.B1(n_484),
.B2(n_486),
.Y(n_509)
);

XOR2xp5_ASAP7_75t_L g515 ( 
.A(n_509),
.B(n_512),
.Y(n_515)
);

FAx1_ASAP7_75t_SL g511 ( 
.A(n_493),
.B(n_500),
.CI(n_489),
.CON(n_511),
.SN(n_511)
);

NOR2xp67_ASAP7_75t_L g519 ( 
.A(n_511),
.B(n_498),
.Y(n_519)
);

MAJIxp5_ASAP7_75t_L g513 ( 
.A(n_491),
.B(n_475),
.C(n_8),
.Y(n_513)
);

OAI21xp5_ASAP7_75t_L g520 ( 
.A1(n_513),
.A2(n_495),
.B(n_497),
.Y(n_520)
);

NAND2x1_ASAP7_75t_L g516 ( 
.A(n_511),
.B(n_492),
.Y(n_516)
);

NAND2xp5_ASAP7_75t_SL g524 ( 
.A(n_516),
.B(n_512),
.Y(n_524)
);

INVxp33_ASAP7_75t_L g518 ( 
.A(n_514),
.Y(n_518)
);

NAND2xp5_ASAP7_75t_L g523 ( 
.A(n_518),
.B(n_520),
.Y(n_523)
);

OAI21xp5_ASAP7_75t_SL g521 ( 
.A1(n_519),
.A2(n_507),
.B(n_505),
.Y(n_521)
);

INVx1_ASAP7_75t_L g526 ( 
.A(n_521),
.Y(n_526)
);

XOR2xp5_ASAP7_75t_L g522 ( 
.A(n_515),
.B(n_505),
.Y(n_522)
);

AND2x2_ASAP7_75t_L g525 ( 
.A(n_522),
.B(n_524),
.Y(n_525)
);

A2O1A1O1Ixp25_ASAP7_75t_SL g527 ( 
.A1(n_526),
.A2(n_517),
.B(n_516),
.C(n_497),
.D(n_508),
.Y(n_527)
);

O2A1O1Ixp33_ASAP7_75t_SL g528 ( 
.A1(n_527),
.A2(n_523),
.B(n_509),
.C(n_506),
.Y(n_528)
);

AOI322xp5_ASAP7_75t_L g529 ( 
.A1(n_528),
.A2(n_510),
.A3(n_525),
.B1(n_513),
.B2(n_502),
.C1(n_7),
.C2(n_9),
.Y(n_529)
);

AND2x2_ASAP7_75t_L g530 ( 
.A(n_529),
.B(n_8),
.Y(n_530)
);

OAI21xp5_ASAP7_75t_L g531 ( 
.A1(n_530),
.A2(n_9),
.B(n_523),
.Y(n_531)
);

XOR2xp5_ASAP7_75t_L g532 ( 
.A(n_531),
.B(n_9),
.Y(n_532)
);


endmodule