module fake_jpeg_29282_n_553 (n_13, n_1, n_10, n_6, n_14, n_18, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_553);

input n_13;
input n_1;
input n_10;
input n_6;
input n_14;
input n_18;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_553;

wire n_529;
wire n_390;
wire n_552;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_525;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_519;
wire n_276;
wire n_143;
wire n_431;
wire n_102;
wire n_549;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_172;
wire n_547;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_513;
wire n_283;
wire n_107;
wire n_490;
wire n_517;
wire n_415;
wire n_479;
wire n_543;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_542;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_48;
wire n_465;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_221;
wire n_256;
wire n_454;
wire n_540;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_508;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_544;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_530;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_298;
wire n_106;
wire n_545;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_474;
wire n_539;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_511;
wire n_305;
wire n_161;
wire n_441;
wire n_342;
wire n_101;
wire n_226;
wire n_509;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_510;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_536;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_537;
wire n_110;
wire n_531;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_352;
wire n_350;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_523;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_533;
wire n_296;
wire n_384;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_491;
wire n_24;
wire n_526;
wire n_467;
wire n_269;
wire n_546;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_473;
wire n_45;
wire n_520;
wire n_476;
wire n_337;
wire n_317;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_481;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_522;
wire n_333;
wire n_518;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_302;
wire n_216;
wire n_528;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_199;
wire n_260;
wire n_550;
wire n_413;
wire n_275;
wire n_494;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_551;
wire n_36;
wire n_62;
wire n_492;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_515;
wire n_347;
wire n_521;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_538;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_534;
wire n_472;
wire n_279;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_484;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_469;
wire n_111;
wire n_197;
wire n_396;
wire n_375;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_527;
wire n_482;
wire n_58;
wire n_41;
wire n_266;
wire n_548;
wire n_72;
wire n_512;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_516;
wire n_183;
wire n_409;
wire n_532;
wire n_249;
wire n_412;
wire n_217;
wire n_471;
wire n_541;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_535;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_524;
wire n_402;
wire n_504;
wire n_438;
wire n_475;
wire n_247;
wire n_157;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_514;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_3),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_14),
.Y(n_20)
);

BUFx8_ASAP7_75t_L g21 ( 
.A(n_9),
.Y(n_21)
);

BUFx3_ASAP7_75t_L g22 ( 
.A(n_9),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_1),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_14),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_5),
.Y(n_25)
);

INVx11_ASAP7_75t_L g26 ( 
.A(n_9),
.Y(n_26)
);

BUFx3_ASAP7_75t_L g27 ( 
.A(n_15),
.Y(n_27)
);

BUFx4f_ASAP7_75t_SL g28 ( 
.A(n_3),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_8),
.Y(n_29)
);

INVx2_ASAP7_75t_L g30 ( 
.A(n_1),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_15),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_2),
.Y(n_32)
);

BUFx12f_ASAP7_75t_L g33 ( 
.A(n_15),
.Y(n_33)
);

BUFx3_ASAP7_75t_L g34 ( 
.A(n_17),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_8),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_16),
.Y(n_36)
);

BUFx16f_ASAP7_75t_L g37 ( 
.A(n_1),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_14),
.Y(n_38)
);

INVx4_ASAP7_75t_L g39 ( 
.A(n_1),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_16),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_18),
.Y(n_41)
);

INVx11_ASAP7_75t_L g42 ( 
.A(n_8),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_3),
.Y(n_43)
);

INVx13_ASAP7_75t_L g44 ( 
.A(n_11),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_2),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_18),
.Y(n_46)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_4),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_4),
.Y(n_48)
);

INVx8_ASAP7_75t_L g49 ( 
.A(n_17),
.Y(n_49)
);

BUFx5_ASAP7_75t_L g50 ( 
.A(n_3),
.Y(n_50)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_0),
.Y(n_51)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_31),
.Y(n_52)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_52),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_20),
.B(n_18),
.Y(n_53)
);

AND2x2_ASAP7_75t_L g129 ( 
.A(n_53),
.B(n_79),
.Y(n_129)
);

BUFx12f_ASAP7_75t_L g54 ( 
.A(n_44),
.Y(n_54)
);

BUFx8_ASAP7_75t_L g133 ( 
.A(n_54),
.Y(n_133)
);

INVx3_ASAP7_75t_L g55 ( 
.A(n_33),
.Y(n_55)
);

INVx3_ASAP7_75t_L g118 ( 
.A(n_55),
.Y(n_118)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_48),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g116 ( 
.A(n_56),
.Y(n_116)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_48),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g123 ( 
.A(n_57),
.Y(n_123)
);

INVx8_ASAP7_75t_L g58 ( 
.A(n_21),
.Y(n_58)
);

INVx8_ASAP7_75t_L g131 ( 
.A(n_58),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_SL g59 ( 
.A(n_20),
.B(n_10),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_L g107 ( 
.A(n_59),
.B(n_63),
.Y(n_107)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_48),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g135 ( 
.A(n_60),
.Y(n_135)
);

BUFx5_ASAP7_75t_L g61 ( 
.A(n_33),
.Y(n_61)
);

INVx5_ASAP7_75t_L g146 ( 
.A(n_61),
.Y(n_146)
);

INVx8_ASAP7_75t_L g62 ( 
.A(n_21),
.Y(n_62)
);

INVx8_ASAP7_75t_L g150 ( 
.A(n_62),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_L g63 ( 
.A(n_24),
.B(n_10),
.Y(n_63)
);

INVx11_ASAP7_75t_L g64 ( 
.A(n_37),
.Y(n_64)
);

INVx6_ASAP7_75t_L g105 ( 
.A(n_64),
.Y(n_105)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_31),
.Y(n_65)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_65),
.Y(n_125)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_30),
.Y(n_66)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_66),
.Y(n_156)
);

INVx4_ASAP7_75t_L g67 ( 
.A(n_39),
.Y(n_67)
);

INVx4_ASAP7_75t_L g155 ( 
.A(n_67),
.Y(n_155)
);

INVx8_ASAP7_75t_L g68 ( 
.A(n_21),
.Y(n_68)
);

BUFx6f_ASAP7_75t_L g142 ( 
.A(n_68),
.Y(n_142)
);

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_48),
.Y(n_69)
);

INVx6_ASAP7_75t_L g114 ( 
.A(n_69),
.Y(n_114)
);

INVx8_ASAP7_75t_L g70 ( 
.A(n_21),
.Y(n_70)
);

INVx5_ASAP7_75t_L g168 ( 
.A(n_70),
.Y(n_168)
);

CKINVDCx16_ASAP7_75t_R g71 ( 
.A(n_37),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_71),
.B(n_72),
.Y(n_109)
);

CKINVDCx20_ASAP7_75t_R g72 ( 
.A(n_22),
.Y(n_72)
);

INVx8_ASAP7_75t_L g73 ( 
.A(n_21),
.Y(n_73)
);

INVx6_ASAP7_75t_L g122 ( 
.A(n_73),
.Y(n_122)
);

INVx2_ASAP7_75t_L g74 ( 
.A(n_30),
.Y(n_74)
);

INVx2_ASAP7_75t_L g115 ( 
.A(n_74),
.Y(n_115)
);

BUFx12f_ASAP7_75t_L g75 ( 
.A(n_44),
.Y(n_75)
);

INVx3_ASAP7_75t_L g130 ( 
.A(n_75),
.Y(n_130)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_30),
.Y(n_76)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_76),
.Y(n_157)
);

BUFx3_ASAP7_75t_L g77 ( 
.A(n_50),
.Y(n_77)
);

BUFx3_ASAP7_75t_L g153 ( 
.A(n_77),
.Y(n_153)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_35),
.Y(n_78)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_78),
.Y(n_163)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_24),
.B(n_10),
.Y(n_79)
);

INVx2_ASAP7_75t_L g80 ( 
.A(n_39),
.Y(n_80)
);

INVx2_ASAP7_75t_L g120 ( 
.A(n_80),
.Y(n_120)
);

BUFx6f_ASAP7_75t_L g81 ( 
.A(n_29),
.Y(n_81)
);

INVx6_ASAP7_75t_L g128 ( 
.A(n_81),
.Y(n_128)
);

INVx1_ASAP7_75t_SL g82 ( 
.A(n_37),
.Y(n_82)
);

AND2x2_ASAP7_75t_L g136 ( 
.A(n_82),
.B(n_91),
.Y(n_136)
);

BUFx12f_ASAP7_75t_L g83 ( 
.A(n_44),
.Y(n_83)
);

INVx3_ASAP7_75t_L g148 ( 
.A(n_83),
.Y(n_148)
);

INVx2_ASAP7_75t_L g84 ( 
.A(n_39),
.Y(n_84)
);

INVx2_ASAP7_75t_L g126 ( 
.A(n_84),
.Y(n_126)
);

BUFx3_ASAP7_75t_L g85 ( 
.A(n_50),
.Y(n_85)
);

INVx4_ASAP7_75t_L g159 ( 
.A(n_85),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_SL g86 ( 
.A(n_38),
.B(n_7),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_L g132 ( 
.A(n_86),
.B(n_46),
.Y(n_132)
);

BUFx6f_ASAP7_75t_L g87 ( 
.A(n_29),
.Y(n_87)
);

INVx6_ASAP7_75t_L g145 ( 
.A(n_87),
.Y(n_145)
);

CKINVDCx20_ASAP7_75t_R g88 ( 
.A(n_22),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g119 ( 
.A(n_88),
.B(n_93),
.Y(n_119)
);

BUFx8_ASAP7_75t_L g89 ( 
.A(n_33),
.Y(n_89)
);

BUFx2_ASAP7_75t_L g108 ( 
.A(n_89),
.Y(n_108)
);

BUFx5_ASAP7_75t_L g90 ( 
.A(n_33),
.Y(n_90)
);

INVx5_ASAP7_75t_SL g117 ( 
.A(n_90),
.Y(n_117)
);

INVx3_ASAP7_75t_SL g91 ( 
.A(n_50),
.Y(n_91)
);

BUFx6f_ASAP7_75t_L g92 ( 
.A(n_29),
.Y(n_92)
);

INVx2_ASAP7_75t_L g134 ( 
.A(n_92),
.Y(n_134)
);

CKINVDCx20_ASAP7_75t_R g93 ( 
.A(n_22),
.Y(n_93)
);

INVx2_ASAP7_75t_R g94 ( 
.A(n_37),
.Y(n_94)
);

OR2x2_ASAP7_75t_L g151 ( 
.A(n_94),
.B(n_23),
.Y(n_151)
);

NOR2xp33_ASAP7_75t_SL g95 ( 
.A(n_38),
.B(n_7),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g121 ( 
.A(n_95),
.B(n_98),
.Y(n_121)
);

BUFx8_ASAP7_75t_L g96 ( 
.A(n_33),
.Y(n_96)
);

BUFx12f_ASAP7_75t_L g124 ( 
.A(n_96),
.Y(n_124)
);

INVx4_ASAP7_75t_L g97 ( 
.A(n_37),
.Y(n_97)
);

HB1xp67_ASAP7_75t_L g110 ( 
.A(n_97),
.Y(n_110)
);

INVxp67_ASAP7_75t_L g98 ( 
.A(n_35),
.Y(n_98)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_35),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g137 ( 
.A(n_99),
.B(n_102),
.Y(n_137)
);

INVx3_ASAP7_75t_L g100 ( 
.A(n_27),
.Y(n_100)
);

INVx2_ASAP7_75t_L g141 ( 
.A(n_100),
.Y(n_141)
);

BUFx3_ASAP7_75t_L g101 ( 
.A(n_26),
.Y(n_101)
);

INVx2_ASAP7_75t_L g144 ( 
.A(n_101),
.Y(n_144)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_41),
.B(n_17),
.Y(n_102)
);

INVx8_ASAP7_75t_L g103 ( 
.A(n_29),
.Y(n_103)
);

INVx2_ASAP7_75t_L g147 ( 
.A(n_103),
.Y(n_147)
);

BUFx6f_ASAP7_75t_L g104 ( 
.A(n_40),
.Y(n_104)
);

INVx2_ASAP7_75t_L g158 ( 
.A(n_104),
.Y(n_158)
);

OAI22xp5_ASAP7_75t_L g106 ( 
.A1(n_81),
.A2(n_40),
.B1(n_46),
.B2(n_41),
.Y(n_106)
);

AOI22xp5_ASAP7_75t_L g183 ( 
.A1(n_106),
.A2(n_36),
.B1(n_45),
.B2(n_43),
.Y(n_183)
);

AOI22xp33_ASAP7_75t_SL g111 ( 
.A1(n_94),
.A2(n_49),
.B1(n_27),
.B2(n_34),
.Y(n_111)
);

AOI22xp33_ASAP7_75t_SL g175 ( 
.A1(n_111),
.A2(n_112),
.B1(n_73),
.B2(n_68),
.Y(n_175)
);

AOI22xp33_ASAP7_75t_SL g112 ( 
.A1(n_58),
.A2(n_49),
.B1(n_27),
.B2(n_34),
.Y(n_112)
);

CKINVDCx20_ASAP7_75t_R g127 ( 
.A(n_101),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_L g179 ( 
.A(n_127),
.B(n_138),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_L g174 ( 
.A(n_132),
.B(n_143),
.Y(n_174)
);

NOR2xp33_ASAP7_75t_SL g138 ( 
.A(n_98),
.B(n_25),
.Y(n_138)
);

NOR2xp67_ASAP7_75t_L g139 ( 
.A(n_54),
.B(n_25),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_L g187 ( 
.A(n_139),
.B(n_154),
.Y(n_187)
);

AOI22xp5_ASAP7_75t_L g140 ( 
.A1(n_87),
.A2(n_40),
.B1(n_36),
.B2(n_34),
.Y(n_140)
);

OAI22xp5_ASAP7_75t_SL g211 ( 
.A1(n_140),
.A2(n_42),
.B1(n_26),
.B2(n_64),
.Y(n_211)
);

NOR2xp33_ASAP7_75t_L g143 ( 
.A(n_54),
.B(n_43),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_L g149 ( 
.A(n_75),
.B(n_23),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_L g210 ( 
.A(n_149),
.B(n_152),
.Y(n_210)
);

INVxp67_ASAP7_75t_L g177 ( 
.A(n_151),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_L g152 ( 
.A(n_75),
.B(n_51),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_L g154 ( 
.A(n_83),
.B(n_51),
.Y(n_154)
);

INVx2_ASAP7_75t_L g160 ( 
.A(n_55),
.Y(n_160)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_160),
.Y(n_170)
);

AND2x2_ASAP7_75t_SL g161 ( 
.A(n_67),
.B(n_40),
.Y(n_161)
);

MAJIxp5_ASAP7_75t_L g220 ( 
.A(n_161),
.B(n_28),
.C(n_42),
.Y(n_220)
);

NOR2xp33_ASAP7_75t_L g162 ( 
.A(n_83),
.B(n_19),
.Y(n_162)
);

NOR2xp33_ASAP7_75t_L g189 ( 
.A(n_162),
.B(n_167),
.Y(n_189)
);

BUFx12f_ASAP7_75t_L g164 ( 
.A(n_56),
.Y(n_164)
);

INVx3_ASAP7_75t_L g180 ( 
.A(n_164),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_L g165 ( 
.A(n_82),
.B(n_19),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_SL g171 ( 
.A(n_165),
.B(n_45),
.Y(n_171)
);

AOI21xp33_ASAP7_75t_L g166 ( 
.A1(n_91),
.A2(n_36),
.B(n_32),
.Y(n_166)
);

AOI21xp33_ASAP7_75t_L g217 ( 
.A1(n_166),
.A2(n_96),
.B(n_89),
.Y(n_217)
);

OR2x2_ASAP7_75t_L g167 ( 
.A(n_89),
.B(n_47),
.Y(n_167)
);

AND2x2_ASAP7_75t_SL g169 ( 
.A(n_115),
.B(n_97),
.Y(n_169)
);

FAx1_ASAP7_75t_SL g231 ( 
.A(n_169),
.B(n_136),
.CI(n_124),
.CON(n_231),
.SN(n_231)
);

NAND3xp33_ASAP7_75t_L g242 ( 
.A(n_171),
.B(n_16),
.C(n_13),
.Y(n_242)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_163),
.Y(n_172)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_172),
.Y(n_232)
);

BUFx6f_ASAP7_75t_L g173 ( 
.A(n_116),
.Y(n_173)
);

BUFx6f_ASAP7_75t_L g235 ( 
.A(n_173),
.Y(n_235)
);

AO21x1_ASAP7_75t_L g241 ( 
.A1(n_175),
.A2(n_188),
.B(n_193),
.Y(n_241)
);

INVx5_ASAP7_75t_L g176 ( 
.A(n_168),
.Y(n_176)
);

INVx5_ASAP7_75t_L g270 ( 
.A(n_176),
.Y(n_270)
);

INVx4_ASAP7_75t_L g178 ( 
.A(n_144),
.Y(n_178)
);

INVx1_ASAP7_75t_SL g258 ( 
.A(n_178),
.Y(n_258)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_113),
.Y(n_181)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_181),
.Y(n_236)
);

CKINVDCx12_ASAP7_75t_R g182 ( 
.A(n_133),
.Y(n_182)
);

CKINVDCx16_ASAP7_75t_R g248 ( 
.A(n_182),
.Y(n_248)
);

OAI22xp5_ASAP7_75t_L g254 ( 
.A1(n_183),
.A2(n_194),
.B1(n_201),
.B2(n_203),
.Y(n_254)
);

BUFx10_ASAP7_75t_L g184 ( 
.A(n_133),
.Y(n_184)
);

CKINVDCx20_ASAP7_75t_R g252 ( 
.A(n_184),
.Y(n_252)
);

INVx6_ASAP7_75t_L g185 ( 
.A(n_116),
.Y(n_185)
);

BUFx6f_ASAP7_75t_L g262 ( 
.A(n_185),
.Y(n_262)
);

BUFx6f_ASAP7_75t_L g186 ( 
.A(n_123),
.Y(n_186)
);

BUFx2_ASAP7_75t_L g246 ( 
.A(n_186),
.Y(n_246)
);

AOI22xp33_ASAP7_75t_SL g188 ( 
.A1(n_117),
.A2(n_49),
.B1(n_100),
.B2(n_62),
.Y(n_188)
);

NOR2xp33_ASAP7_75t_L g190 ( 
.A(n_121),
.B(n_137),
.Y(n_190)
);

NOR2xp33_ASAP7_75t_SL g255 ( 
.A(n_190),
.B(n_192),
.Y(n_255)
);

NAND2xp5_ASAP7_75t_SL g191 ( 
.A(n_107),
.B(n_47),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_L g233 ( 
.A(n_191),
.B(n_216),
.Y(n_233)
);

NOR2xp33_ASAP7_75t_L g192 ( 
.A(n_129),
.B(n_96),
.Y(n_192)
);

AOI22xp33_ASAP7_75t_SL g193 ( 
.A1(n_117),
.A2(n_70),
.B1(n_103),
.B2(n_85),
.Y(n_193)
);

AOI22xp33_ASAP7_75t_SL g194 ( 
.A1(n_156),
.A2(n_77),
.B1(n_32),
.B2(n_90),
.Y(n_194)
);

INVx2_ASAP7_75t_L g195 ( 
.A(n_110),
.Y(n_195)
);

INVx2_ASAP7_75t_L g234 ( 
.A(n_195),
.Y(n_234)
);

INVx2_ASAP7_75t_L g196 ( 
.A(n_110),
.Y(n_196)
);

INVx2_ASAP7_75t_L g244 ( 
.A(n_196),
.Y(n_244)
);

INVx11_ASAP7_75t_L g197 ( 
.A(n_142),
.Y(n_197)
);

BUFx3_ASAP7_75t_L g274 ( 
.A(n_197),
.Y(n_274)
);

INVx3_ASAP7_75t_L g198 ( 
.A(n_105),
.Y(n_198)
);

INVx1_ASAP7_75t_SL g271 ( 
.A(n_198),
.Y(n_271)
);

BUFx12_ASAP7_75t_L g199 ( 
.A(n_146),
.Y(n_199)
);

NOR2xp33_ASAP7_75t_L g239 ( 
.A(n_199),
.B(n_221),
.Y(n_239)
);

BUFx3_ASAP7_75t_L g200 ( 
.A(n_153),
.Y(n_200)
);

INVx4_ASAP7_75t_L g249 ( 
.A(n_200),
.Y(n_249)
);

AOI22xp33_ASAP7_75t_SL g201 ( 
.A1(n_157),
.A2(n_32),
.B1(n_92),
.B2(n_104),
.Y(n_201)
);

CKINVDCx20_ASAP7_75t_R g202 ( 
.A(n_119),
.Y(n_202)
);

NAND2xp5_ASAP7_75t_SL g240 ( 
.A(n_202),
.B(n_204),
.Y(n_240)
);

AOI22xp33_ASAP7_75t_SL g203 ( 
.A1(n_111),
.A2(n_57),
.B1(n_69),
.B2(n_60),
.Y(n_203)
);

CKINVDCx20_ASAP7_75t_R g204 ( 
.A(n_109),
.Y(n_204)
);

INVx2_ASAP7_75t_L g205 ( 
.A(n_118),
.Y(n_205)
);

INVx2_ASAP7_75t_L g277 ( 
.A(n_205),
.Y(n_277)
);

BUFx12f_ASAP7_75t_L g206 ( 
.A(n_142),
.Y(n_206)
);

INVx3_ASAP7_75t_L g237 ( 
.A(n_206),
.Y(n_237)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_125),
.Y(n_207)
);

CKINVDCx16_ASAP7_75t_R g268 ( 
.A(n_207),
.Y(n_268)
);

INVx13_ASAP7_75t_L g208 ( 
.A(n_130),
.Y(n_208)
);

INVx3_ASAP7_75t_L g257 ( 
.A(n_208),
.Y(n_257)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_120),
.Y(n_209)
);

CKINVDCx16_ASAP7_75t_R g283 ( 
.A(n_209),
.Y(n_283)
);

AOI22xp5_ASAP7_75t_L g245 ( 
.A1(n_211),
.A2(n_145),
.B1(n_128),
.B2(n_114),
.Y(n_245)
);

BUFx3_ASAP7_75t_L g212 ( 
.A(n_153),
.Y(n_212)
);

INVx4_ASAP7_75t_L g263 ( 
.A(n_212),
.Y(n_263)
);

INVx2_ASAP7_75t_L g213 ( 
.A(n_134),
.Y(n_213)
);

INVx4_ASAP7_75t_L g280 ( 
.A(n_213),
.Y(n_280)
);

BUFx2_ASAP7_75t_L g214 ( 
.A(n_131),
.Y(n_214)
);

INVx3_ASAP7_75t_L g261 ( 
.A(n_214),
.Y(n_261)
);

INVx5_ASAP7_75t_L g215 ( 
.A(n_105),
.Y(n_215)
);

INVx3_ASAP7_75t_L g265 ( 
.A(n_215),
.Y(n_265)
);

NAND2xp5_ASAP7_75t_SL g216 ( 
.A(n_129),
.B(n_12),
.Y(n_216)
);

AND2x2_ASAP7_75t_L g250 ( 
.A(n_217),
.B(n_220),
.Y(n_250)
);

NAND2xp5_ASAP7_75t_L g218 ( 
.A(n_151),
.B(n_28),
.Y(n_218)
);

NAND2xp5_ASAP7_75t_L g279 ( 
.A(n_218),
.B(n_177),
.Y(n_279)
);

AOI22xp33_ASAP7_75t_SL g219 ( 
.A1(n_112),
.A2(n_28),
.B1(n_42),
.B2(n_26),
.Y(n_219)
);

AOI22xp33_ASAP7_75t_SL g243 ( 
.A1(n_219),
.A2(n_227),
.B1(n_108),
.B2(n_164),
.Y(n_243)
);

CKINVDCx20_ASAP7_75t_R g221 ( 
.A(n_167),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_SL g222 ( 
.A(n_136),
.B(n_7),
.Y(n_222)
);

NAND2xp5_ASAP7_75t_L g251 ( 
.A(n_222),
.B(n_13),
.Y(n_251)
);

INVx2_ASAP7_75t_L g223 ( 
.A(n_158),
.Y(n_223)
);

CKINVDCx20_ASAP7_75t_R g264 ( 
.A(n_223),
.Y(n_264)
);

BUFx6f_ASAP7_75t_L g224 ( 
.A(n_123),
.Y(n_224)
);

INVxp33_ASAP7_75t_L g259 ( 
.A(n_224),
.Y(n_259)
);

OAI21xp33_ASAP7_75t_L g225 ( 
.A1(n_161),
.A2(n_28),
.B(n_2),
.Y(n_225)
);

AOI21xp5_ASAP7_75t_SL g267 ( 
.A1(n_225),
.A2(n_147),
.B(n_108),
.Y(n_267)
);

INVx5_ASAP7_75t_L g226 ( 
.A(n_148),
.Y(n_226)
);

NOR2xp33_ASAP7_75t_L g247 ( 
.A(n_226),
.B(n_228),
.Y(n_247)
);

AOI22xp33_ASAP7_75t_SL g227 ( 
.A1(n_159),
.A2(n_28),
.B1(n_11),
.B2(n_12),
.Y(n_227)
);

INVx3_ASAP7_75t_L g228 ( 
.A(n_164),
.Y(n_228)
);

CKINVDCx12_ASAP7_75t_R g229 ( 
.A(n_124),
.Y(n_229)
);

NOR2xp33_ASAP7_75t_L g253 ( 
.A(n_229),
.B(n_230),
.Y(n_253)
);

CKINVDCx12_ASAP7_75t_R g230 ( 
.A(n_124),
.Y(n_230)
);

AND2x2_ASAP7_75t_L g320 ( 
.A(n_231),
.B(n_279),
.Y(n_320)
);

OAI22xp5_ASAP7_75t_SL g238 ( 
.A1(n_183),
.A2(n_128),
.B1(n_145),
.B2(n_114),
.Y(n_238)
);

OAI22xp5_ASAP7_75t_L g329 ( 
.A1(n_238),
.A2(n_245),
.B1(n_185),
.B2(n_224),
.Y(n_329)
);

NOR2xp33_ASAP7_75t_L g287 ( 
.A(n_242),
.B(n_273),
.Y(n_287)
);

INVxp67_ASAP7_75t_L g285 ( 
.A(n_243),
.Y(n_285)
);

NAND2xp5_ASAP7_75t_SL g286 ( 
.A(n_251),
.B(n_256),
.Y(n_286)
);

NAND2xp5_ASAP7_75t_L g256 ( 
.A(n_210),
.B(n_126),
.Y(n_256)
);

NOR2xp33_ASAP7_75t_L g260 ( 
.A(n_179),
.B(n_141),
.Y(n_260)
);

NAND2xp5_ASAP7_75t_SL g321 ( 
.A(n_260),
.B(n_272),
.Y(n_321)
);

XNOR2xp5_ASAP7_75t_L g266 ( 
.A(n_218),
.B(n_155),
.Y(n_266)
);

MAJIxp5_ASAP7_75t_L g331 ( 
.A(n_266),
.B(n_269),
.C(n_282),
.Y(n_331)
);

OAI21xp5_ASAP7_75t_SL g302 ( 
.A1(n_267),
.A2(n_178),
.B(n_196),
.Y(n_302)
);

MAJIxp5_ASAP7_75t_L g269 ( 
.A(n_220),
.B(n_159),
.C(n_122),
.Y(n_269)
);

NOR2xp33_ASAP7_75t_L g272 ( 
.A(n_189),
.B(n_150),
.Y(n_272)
);

CKINVDCx20_ASAP7_75t_R g273 ( 
.A(n_184),
.Y(n_273)
);

NOR2xp33_ASAP7_75t_L g275 ( 
.A(n_187),
.B(n_150),
.Y(n_275)
);

NOR2xp33_ASAP7_75t_L g290 ( 
.A(n_275),
.B(n_278),
.Y(n_290)
);

AOI22xp33_ASAP7_75t_SL g276 ( 
.A1(n_214),
.A2(n_131),
.B1(n_122),
.B2(n_135),
.Y(n_276)
);

INVxp67_ASAP7_75t_L g313 ( 
.A(n_276),
.Y(n_313)
);

NOR2xp33_ASAP7_75t_SL g278 ( 
.A(n_174),
.B(n_13),
.Y(n_278)
);

NOR2xp33_ASAP7_75t_L g281 ( 
.A(n_177),
.B(n_12),
.Y(n_281)
);

NOR2xp33_ASAP7_75t_L g291 ( 
.A(n_281),
.B(n_199),
.Y(n_291)
);

MAJIxp5_ASAP7_75t_L g282 ( 
.A(n_169),
.B(n_135),
.C(n_11),
.Y(n_282)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_234),
.Y(n_284)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_284),
.Y(n_334)
);

INVx13_ASAP7_75t_L g288 ( 
.A(n_257),
.Y(n_288)
);

INVx13_ASAP7_75t_L g355 ( 
.A(n_288),
.Y(n_355)
);

NAND2xp5_ASAP7_75t_L g289 ( 
.A(n_266),
.B(n_279),
.Y(n_289)
);

NAND2xp5_ASAP7_75t_L g343 ( 
.A(n_289),
.B(n_293),
.Y(n_343)
);

CKINVDCx14_ASAP7_75t_R g337 ( 
.A(n_291),
.Y(n_337)
);

NOR2xp33_ASAP7_75t_L g292 ( 
.A(n_239),
.B(n_208),
.Y(n_292)
);

NAND2xp5_ASAP7_75t_SL g340 ( 
.A(n_292),
.B(n_298),
.Y(n_340)
);

OAI22xp5_ASAP7_75t_SL g293 ( 
.A1(n_245),
.A2(n_211),
.B1(n_225),
.B2(n_213),
.Y(n_293)
);

INVx3_ASAP7_75t_L g294 ( 
.A(n_235),
.Y(n_294)
);

BUFx2_ASAP7_75t_L g372 ( 
.A(n_294),
.Y(n_372)
);

INVx2_ASAP7_75t_L g295 ( 
.A(n_277),
.Y(n_295)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_295),
.Y(n_339)
);

NAND2xp5_ASAP7_75t_L g296 ( 
.A(n_250),
.B(n_169),
.Y(n_296)
);

NAND2xp5_ASAP7_75t_L g344 ( 
.A(n_296),
.B(n_299),
.Y(n_344)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_234),
.Y(n_297)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_297),
.Y(n_336)
);

NOR2xp33_ASAP7_75t_L g298 ( 
.A(n_268),
.B(n_226),
.Y(n_298)
);

NAND2xp5_ASAP7_75t_L g299 ( 
.A(n_250),
.B(n_195),
.Y(n_299)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_244),
.Y(n_300)
);

INVx1_ASAP7_75t_L g356 ( 
.A(n_300),
.Y(n_356)
);

NOR2xp33_ASAP7_75t_L g301 ( 
.A(n_240),
.B(n_205),
.Y(n_301)
);

NAND2xp5_ASAP7_75t_SL g354 ( 
.A(n_301),
.B(n_303),
.Y(n_354)
);

AOI21xp5_ASAP7_75t_L g347 ( 
.A1(n_302),
.A2(n_318),
.B(n_327),
.Y(n_347)
);

OR2x2_ASAP7_75t_L g303 ( 
.A(n_231),
.B(n_170),
.Y(n_303)
);

INVx5_ASAP7_75t_L g304 ( 
.A(n_270),
.Y(n_304)
);

INVx1_ASAP7_75t_L g350 ( 
.A(n_304),
.Y(n_350)
);

NOR2xp33_ASAP7_75t_L g305 ( 
.A(n_255),
.B(n_199),
.Y(n_305)
);

NOR2xp33_ASAP7_75t_L g338 ( 
.A(n_305),
.B(n_307),
.Y(n_338)
);

INVx6_ASAP7_75t_L g306 ( 
.A(n_235),
.Y(n_306)
);

INVx1_ASAP7_75t_L g363 ( 
.A(n_306),
.Y(n_363)
);

NOR2xp33_ASAP7_75t_L g307 ( 
.A(n_232),
.B(n_176),
.Y(n_307)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_244),
.Y(n_308)
);

INVx1_ASAP7_75t_L g357 ( 
.A(n_308),
.Y(n_357)
);

BUFx6f_ASAP7_75t_L g309 ( 
.A(n_262),
.Y(n_309)
);

INVx1_ASAP7_75t_L g370 ( 
.A(n_309),
.Y(n_370)
);

INVx2_ASAP7_75t_L g310 ( 
.A(n_277),
.Y(n_310)
);

INVx1_ASAP7_75t_L g361 ( 
.A(n_310),
.Y(n_361)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_236),
.Y(n_311)
);

INVx1_ASAP7_75t_L g362 ( 
.A(n_311),
.Y(n_362)
);

INVx3_ASAP7_75t_L g312 ( 
.A(n_274),
.Y(n_312)
);

INVxp67_ASAP7_75t_L g341 ( 
.A(n_312),
.Y(n_341)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_280),
.Y(n_314)
);

INVx1_ASAP7_75t_L g364 ( 
.A(n_314),
.Y(n_364)
);

INVx13_ASAP7_75t_L g315 ( 
.A(n_257),
.Y(n_315)
);

INVxp67_ASAP7_75t_L g342 ( 
.A(n_315),
.Y(n_342)
);

AND2x6_ASAP7_75t_L g316 ( 
.A(n_250),
.B(n_200),
.Y(n_316)
);

OAI21xp5_ASAP7_75t_SL g352 ( 
.A1(n_316),
.A2(n_263),
.B(n_249),
.Y(n_352)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_280),
.Y(n_317)
);

INVx1_ASAP7_75t_L g365 ( 
.A(n_317),
.Y(n_365)
);

OAI21xp5_ASAP7_75t_SL g318 ( 
.A1(n_267),
.A2(n_223),
.B(n_198),
.Y(n_318)
);

NOR2xp33_ASAP7_75t_L g319 ( 
.A(n_233),
.B(n_206),
.Y(n_319)
);

INVxp67_ASAP7_75t_L g358 ( 
.A(n_319),
.Y(n_358)
);

CKINVDCx20_ASAP7_75t_R g322 ( 
.A(n_247),
.Y(n_322)
);

CKINVDCx20_ASAP7_75t_R g335 ( 
.A(n_322),
.Y(n_335)
);

INVxp67_ASAP7_75t_L g323 ( 
.A(n_253),
.Y(n_323)
);

NAND2xp5_ASAP7_75t_L g348 ( 
.A(n_323),
.B(n_328),
.Y(n_348)
);

INVx3_ASAP7_75t_L g324 ( 
.A(n_274),
.Y(n_324)
);

INVx1_ASAP7_75t_L g367 ( 
.A(n_324),
.Y(n_367)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_271),
.Y(n_325)
);

AND2x2_ASAP7_75t_L g333 ( 
.A(n_325),
.B(n_326),
.Y(n_333)
);

INVx3_ASAP7_75t_L g326 ( 
.A(n_262),
.Y(n_326)
);

AOI21xp5_ASAP7_75t_L g327 ( 
.A1(n_241),
.A2(n_212),
.B(n_228),
.Y(n_327)
);

CKINVDCx5p33_ASAP7_75t_R g328 ( 
.A(n_231),
.Y(n_328)
);

AND2x2_ASAP7_75t_L g349 ( 
.A(n_329),
.B(n_330),
.Y(n_349)
);

AND2x2_ASAP7_75t_L g330 ( 
.A(n_269),
.B(n_180),
.Y(n_330)
);

OAI22xp5_ASAP7_75t_SL g332 ( 
.A1(n_299),
.A2(n_254),
.B1(n_241),
.B2(n_238),
.Y(n_332)
);

AOI22xp5_ASAP7_75t_L g390 ( 
.A1(n_332),
.A2(n_353),
.B1(n_293),
.B2(n_325),
.Y(n_390)
);

XOR2xp5_ASAP7_75t_L g345 ( 
.A(n_331),
.B(n_282),
.Y(n_345)
);

MAJIxp5_ASAP7_75t_L g379 ( 
.A(n_345),
.B(n_368),
.C(n_369),
.Y(n_379)
);

XNOR2xp5_ASAP7_75t_L g346 ( 
.A(n_289),
.B(n_283),
.Y(n_346)
);

XNOR2xp5_ASAP7_75t_SL g392 ( 
.A(n_346),
.B(n_366),
.Y(n_392)
);

NAND2xp5_ASAP7_75t_L g351 ( 
.A(n_320),
.B(n_331),
.Y(n_351)
);

NAND2xp5_ASAP7_75t_L g380 ( 
.A(n_351),
.B(n_359),
.Y(n_380)
);

INVxp67_ASAP7_75t_L g375 ( 
.A(n_352),
.Y(n_375)
);

OAI22xp5_ASAP7_75t_SL g353 ( 
.A1(n_285),
.A2(n_264),
.B1(n_186),
.B2(n_173),
.Y(n_353)
);

NAND2xp5_ASAP7_75t_L g359 ( 
.A(n_320),
.B(n_252),
.Y(n_359)
);

OA21x2_ASAP7_75t_L g360 ( 
.A1(n_327),
.A2(n_258),
.B(n_271),
.Y(n_360)
);

NAND2xp5_ASAP7_75t_L g383 ( 
.A(n_360),
.B(n_371),
.Y(n_383)
);

XNOR2xp5_ASAP7_75t_L g366 ( 
.A(n_320),
.B(n_248),
.Y(n_366)
);

MAJIxp5_ASAP7_75t_L g368 ( 
.A(n_330),
.B(n_258),
.C(n_263),
.Y(n_368)
);

MAJIxp5_ASAP7_75t_L g369 ( 
.A(n_330),
.B(n_249),
.C(n_265),
.Y(n_369)
);

NAND2xp5_ASAP7_75t_L g371 ( 
.A(n_303),
.B(n_261),
.Y(n_371)
);

CKINVDCx20_ASAP7_75t_R g373 ( 
.A(n_321),
.Y(n_373)
);

NOR2xp33_ASAP7_75t_L g388 ( 
.A(n_373),
.B(n_323),
.Y(n_388)
);

OAI22xp5_ASAP7_75t_L g374 ( 
.A1(n_347),
.A2(n_285),
.B1(n_313),
.B2(n_316),
.Y(n_374)
);

NAND2xp5_ASAP7_75t_L g410 ( 
.A(n_374),
.B(n_376),
.Y(n_410)
);

INVx1_ASAP7_75t_SL g376 ( 
.A(n_333),
.Y(n_376)
);

NOR2xp33_ASAP7_75t_SL g377 ( 
.A(n_348),
.B(n_290),
.Y(n_377)
);

NOR2xp33_ASAP7_75t_SL g421 ( 
.A(n_377),
.B(n_388),
.Y(n_421)
);

INVx1_ASAP7_75t_L g378 ( 
.A(n_362),
.Y(n_378)
);

INVx1_ASAP7_75t_L g413 ( 
.A(n_378),
.Y(n_413)
);

MAJIxp5_ASAP7_75t_L g381 ( 
.A(n_351),
.B(n_296),
.C(n_302),
.Y(n_381)
);

MAJIxp5_ASAP7_75t_L g437 ( 
.A(n_381),
.B(n_300),
.C(n_297),
.Y(n_437)
);

OAI21xp5_ASAP7_75t_SL g382 ( 
.A1(n_347),
.A2(n_328),
.B(n_313),
.Y(n_382)
);

NAND2xp5_ASAP7_75t_SL g434 ( 
.A(n_382),
.B(n_389),
.Y(n_434)
);

NAND2xp5_ASAP7_75t_L g384 ( 
.A(n_348),
.B(n_286),
.Y(n_384)
);

INVx1_ASAP7_75t_L g418 ( 
.A(n_384),
.Y(n_418)
);

OAI22xp5_ASAP7_75t_L g385 ( 
.A1(n_349),
.A2(n_343),
.B1(n_332),
.B2(n_359),
.Y(n_385)
);

NAND2xp5_ASAP7_75t_L g431 ( 
.A(n_385),
.B(n_386),
.Y(n_431)
);

INVx1_ASAP7_75t_SL g386 ( 
.A(n_333),
.Y(n_386)
);

INVx1_ASAP7_75t_L g387 ( 
.A(n_365),
.Y(n_387)
);

INVx1_ASAP7_75t_L g424 ( 
.A(n_387),
.Y(n_424)
);

NOR2xp33_ASAP7_75t_L g389 ( 
.A(n_335),
.B(n_287),
.Y(n_389)
);

OAI22xp5_ASAP7_75t_SL g412 ( 
.A1(n_390),
.A2(n_401),
.B1(n_408),
.B2(n_360),
.Y(n_412)
);

AOI21xp5_ASAP7_75t_L g391 ( 
.A1(n_352),
.A2(n_318),
.B(n_304),
.Y(n_391)
);

OAI21xp5_ASAP7_75t_L g441 ( 
.A1(n_391),
.A2(n_406),
.B(n_383),
.Y(n_441)
);

CKINVDCx12_ASAP7_75t_R g393 ( 
.A(n_342),
.Y(n_393)
);

INVxp67_ASAP7_75t_L g415 ( 
.A(n_393),
.Y(n_415)
);

NOR2xp33_ASAP7_75t_L g394 ( 
.A(n_338),
.B(n_311),
.Y(n_394)
);

CKINVDCx16_ASAP7_75t_R g427 ( 
.A(n_394),
.Y(n_427)
);

INVx1_ASAP7_75t_L g395 ( 
.A(n_334),
.Y(n_395)
);

INVx1_ASAP7_75t_L g435 ( 
.A(n_395),
.Y(n_435)
);

NOR2xp33_ASAP7_75t_L g396 ( 
.A(n_337),
.B(n_358),
.Y(n_396)
);

NOR2xp33_ASAP7_75t_L g411 ( 
.A(n_396),
.B(n_398),
.Y(n_411)
);

INVx1_ASAP7_75t_L g397 ( 
.A(n_336),
.Y(n_397)
);

INVx1_ASAP7_75t_L g440 ( 
.A(n_397),
.Y(n_440)
);

NOR2xp33_ASAP7_75t_L g398 ( 
.A(n_358),
.B(n_315),
.Y(n_398)
);

NOR2xp33_ASAP7_75t_L g399 ( 
.A(n_340),
.B(n_288),
.Y(n_399)
);

NOR2xp33_ASAP7_75t_L g426 ( 
.A(n_399),
.B(n_404),
.Y(n_426)
);

INVx13_ASAP7_75t_L g400 ( 
.A(n_355),
.Y(n_400)
);

INVxp67_ASAP7_75t_L g419 ( 
.A(n_400),
.Y(n_419)
);

AOI22xp5_ASAP7_75t_L g401 ( 
.A1(n_349),
.A2(n_326),
.B1(n_306),
.B2(n_294),
.Y(n_401)
);

INVx1_ASAP7_75t_L g402 ( 
.A(n_356),
.Y(n_402)
);

NAND2xp5_ASAP7_75t_L g432 ( 
.A(n_402),
.B(n_403),
.Y(n_432)
);

INVx1_ASAP7_75t_L g403 ( 
.A(n_357),
.Y(n_403)
);

NAND2xp5_ASAP7_75t_L g404 ( 
.A(n_371),
.B(n_308),
.Y(n_404)
);

NAND2xp5_ASAP7_75t_L g405 ( 
.A(n_343),
.B(n_284),
.Y(n_405)
);

NOR2xp33_ASAP7_75t_L g428 ( 
.A(n_405),
.B(n_407),
.Y(n_428)
);

OR2x2_ASAP7_75t_L g406 ( 
.A(n_349),
.B(n_261),
.Y(n_406)
);

OAI22x1_ASAP7_75t_R g414 ( 
.A1(n_406),
.A2(n_333),
.B1(n_353),
.B2(n_341),
.Y(n_414)
);

NOR2xp33_ASAP7_75t_L g407 ( 
.A(n_354),
.B(n_346),
.Y(n_407)
);

OAI22xp5_ASAP7_75t_SL g408 ( 
.A1(n_344),
.A2(n_369),
.B1(n_368),
.B2(n_360),
.Y(n_408)
);

OAI22xp5_ASAP7_75t_L g409 ( 
.A1(n_344),
.A2(n_309),
.B1(n_246),
.B2(n_324),
.Y(n_409)
);

OAI22xp5_ASAP7_75t_L g425 ( 
.A1(n_409),
.A2(n_372),
.B1(n_339),
.B2(n_361),
.Y(n_425)
);

AOI22xp5_ASAP7_75t_SL g461 ( 
.A1(n_412),
.A2(n_416),
.B1(n_420),
.B2(n_425),
.Y(n_461)
);

INVxp67_ASAP7_75t_L g454 ( 
.A(n_414),
.Y(n_454)
);

OAI22xp5_ASAP7_75t_SL g416 ( 
.A1(n_390),
.A2(n_363),
.B1(n_370),
.B2(n_350),
.Y(n_416)
);

OAI22xp5_ASAP7_75t_L g417 ( 
.A1(n_377),
.A2(n_363),
.B1(n_350),
.B2(n_341),
.Y(n_417)
);

INVx1_ASAP7_75t_L g442 ( 
.A(n_417),
.Y(n_442)
);

OAI22xp5_ASAP7_75t_SL g420 ( 
.A1(n_375),
.A2(n_370),
.B1(n_345),
.B2(n_366),
.Y(n_420)
);

XNOR2xp5_ASAP7_75t_L g422 ( 
.A(n_392),
.B(n_364),
.Y(n_422)
);

XNOR2xp5_ASAP7_75t_L g459 ( 
.A(n_422),
.B(n_392),
.Y(n_459)
);

OAI22xp33_ASAP7_75t_SL g423 ( 
.A1(n_375),
.A2(n_372),
.B1(n_367),
.B2(n_342),
.Y(n_423)
);

INVx1_ASAP7_75t_L g443 ( 
.A(n_423),
.Y(n_443)
);

NOR2xp33_ASAP7_75t_SL g429 ( 
.A(n_384),
.B(n_339),
.Y(n_429)
);

NAND2xp5_ASAP7_75t_SL g456 ( 
.A(n_429),
.B(n_404),
.Y(n_456)
);

NOR3xp33_ASAP7_75t_SL g430 ( 
.A(n_382),
.B(n_355),
.C(n_184),
.Y(n_430)
);

NOR2xp33_ASAP7_75t_SL g458 ( 
.A(n_430),
.B(n_393),
.Y(n_458)
);

NOR2xp33_ASAP7_75t_L g433 ( 
.A(n_380),
.B(n_312),
.Y(n_433)
);

INVx1_ASAP7_75t_L g445 ( 
.A(n_433),
.Y(n_445)
);

NOR2xp33_ASAP7_75t_L g436 ( 
.A(n_380),
.B(n_317),
.Y(n_436)
);

INVx1_ASAP7_75t_L g448 ( 
.A(n_436),
.Y(n_448)
);

MAJIxp5_ASAP7_75t_L g453 ( 
.A(n_437),
.B(n_379),
.C(n_381),
.Y(n_453)
);

NOR2xp33_ASAP7_75t_L g438 ( 
.A(n_385),
.B(n_310),
.Y(n_438)
);

INVx1_ASAP7_75t_L g450 ( 
.A(n_438),
.Y(n_450)
);

NOR2xp33_ASAP7_75t_L g439 ( 
.A(n_408),
.B(n_295),
.Y(n_439)
);

INVx1_ASAP7_75t_L g467 ( 
.A(n_439),
.Y(n_467)
);

OAI21xp5_ASAP7_75t_L g457 ( 
.A1(n_441),
.A2(n_406),
.B(n_414),
.Y(n_457)
);

NOR2xp33_ASAP7_75t_L g444 ( 
.A(n_421),
.B(n_378),
.Y(n_444)
);

INVx1_ASAP7_75t_L g474 ( 
.A(n_444),
.Y(n_474)
);

INVx2_ASAP7_75t_L g446 ( 
.A(n_413),
.Y(n_446)
);

INVx1_ASAP7_75t_L g477 ( 
.A(n_446),
.Y(n_477)
);

NOR2xp33_ASAP7_75t_L g447 ( 
.A(n_421),
.B(n_383),
.Y(n_447)
);

INVx1_ASAP7_75t_L g478 ( 
.A(n_447),
.Y(n_478)
);

INVxp33_ASAP7_75t_SL g449 ( 
.A(n_414),
.Y(n_449)
);

INVx1_ASAP7_75t_L g485 ( 
.A(n_449),
.Y(n_485)
);

XOR2xp5_ASAP7_75t_L g451 ( 
.A(n_422),
.B(n_379),
.Y(n_451)
);

XOR2xp5_ASAP7_75t_L g489 ( 
.A(n_451),
.B(n_457),
.Y(n_489)
);

INVx2_ASAP7_75t_L g452 ( 
.A(n_413),
.Y(n_452)
);

NOR2xp33_ASAP7_75t_L g483 ( 
.A(n_452),
.B(n_455),
.Y(n_483)
);

MAJIxp5_ASAP7_75t_L g469 ( 
.A(n_453),
.B(n_465),
.C(n_466),
.Y(n_469)
);

OAI21xp5_ASAP7_75t_SL g455 ( 
.A1(n_410),
.A2(n_391),
.B(n_374),
.Y(n_455)
);

OAI22xp5_ASAP7_75t_L g476 ( 
.A1(n_456),
.A2(n_458),
.B1(n_426),
.B2(n_411),
.Y(n_476)
);

XNOR2xp5_ASAP7_75t_SL g475 ( 
.A(n_459),
.B(n_462),
.Y(n_475)
);

HB1xp67_ASAP7_75t_L g460 ( 
.A(n_425),
.Y(n_460)
);

NOR2xp33_ASAP7_75t_L g484 ( 
.A(n_460),
.B(n_464),
.Y(n_484)
);

XOR2xp5_ASAP7_75t_L g462 ( 
.A(n_420),
.B(n_405),
.Y(n_462)
);

AOI22xp5_ASAP7_75t_SL g463 ( 
.A1(n_412),
.A2(n_376),
.B1(n_386),
.B2(n_409),
.Y(n_463)
);

OAI22xp5_ASAP7_75t_SL g472 ( 
.A1(n_463),
.A2(n_441),
.B1(n_431),
.B2(n_415),
.Y(n_472)
);

NOR2xp33_ASAP7_75t_L g464 ( 
.A(n_427),
.B(n_387),
.Y(n_464)
);

XNOR2xp5_ASAP7_75t_L g465 ( 
.A(n_437),
.B(n_401),
.Y(n_465)
);

MAJIxp5_ASAP7_75t_L g466 ( 
.A(n_410),
.B(n_403),
.C(n_402),
.Y(n_466)
);

INVx1_ASAP7_75t_L g468 ( 
.A(n_432),
.Y(n_468)
);

AOI22xp33_ASAP7_75t_SL g480 ( 
.A1(n_468),
.A2(n_440),
.B1(n_435),
.B2(n_424),
.Y(n_480)
);

AOI22xp5_ASAP7_75t_L g470 ( 
.A1(n_442),
.A2(n_414),
.B1(n_416),
.B2(n_418),
.Y(n_470)
);

OAI22xp5_ASAP7_75t_L g502 ( 
.A1(n_470),
.A2(n_486),
.B1(n_487),
.B2(n_446),
.Y(n_502)
);

AOI22xp5_ASAP7_75t_SL g471 ( 
.A1(n_443),
.A2(n_418),
.B1(n_430),
.B2(n_415),
.Y(n_471)
);

XOR2xp5_ASAP7_75t_L g494 ( 
.A(n_471),
.B(n_463),
.Y(n_494)
);

AOI22xp5_ASAP7_75t_SL g500 ( 
.A1(n_472),
.A2(n_488),
.B1(n_454),
.B2(n_485),
.Y(n_500)
);

MAJIxp5_ASAP7_75t_L g473 ( 
.A(n_453),
.B(n_431),
.C(n_434),
.Y(n_473)
);

MAJIxp5_ASAP7_75t_L g495 ( 
.A(n_473),
.B(n_490),
.C(n_465),
.Y(n_495)
);

INVx1_ASAP7_75t_L g493 ( 
.A(n_476),
.Y(n_493)
);

OAI22xp5_ASAP7_75t_SL g479 ( 
.A1(n_461),
.A2(n_428),
.B1(n_429),
.B2(n_432),
.Y(n_479)
);

NAND2xp5_ASAP7_75t_L g491 ( 
.A(n_479),
.B(n_482),
.Y(n_491)
);

INVx1_ASAP7_75t_L g508 ( 
.A(n_480),
.Y(n_508)
);

OAI22xp5_ASAP7_75t_L g481 ( 
.A1(n_467),
.A2(n_440),
.B1(n_435),
.B2(n_424),
.Y(n_481)
);

INVx1_ASAP7_75t_L g497 ( 
.A(n_481),
.Y(n_497)
);

FAx1_ASAP7_75t_SL g482 ( 
.A(n_457),
.B(n_397),
.CI(n_395),
.CON(n_482),
.SN(n_482)
);

AOI22xp5_ASAP7_75t_L g486 ( 
.A1(n_450),
.A2(n_419),
.B1(n_246),
.B2(n_400),
.Y(n_486)
);

AOI22xp5_ASAP7_75t_L g487 ( 
.A1(n_454),
.A2(n_419),
.B1(n_400),
.B2(n_270),
.Y(n_487)
);

XOR2x2_ASAP7_75t_SL g488 ( 
.A(n_455),
.B(n_184),
.Y(n_488)
);

MAJIxp5_ASAP7_75t_L g490 ( 
.A(n_451),
.B(n_265),
.C(n_237),
.Y(n_490)
);

NOR2xp33_ASAP7_75t_L g492 ( 
.A(n_473),
.B(n_448),
.Y(n_492)
);

NAND2xp5_ASAP7_75t_L g509 ( 
.A(n_492),
.B(n_496),
.Y(n_509)
);

XNOR2xp5_ASAP7_75t_L g521 ( 
.A(n_494),
.B(n_495),
.Y(n_521)
);

NOR2xp33_ASAP7_75t_SL g496 ( 
.A(n_474),
.B(n_445),
.Y(n_496)
);

XNOR2xp5_ASAP7_75t_L g498 ( 
.A(n_469),
.B(n_461),
.Y(n_498)
);

MAJIxp5_ASAP7_75t_L g511 ( 
.A(n_498),
.B(n_504),
.C(n_505),
.Y(n_511)
);

NOR2xp33_ASAP7_75t_L g499 ( 
.A(n_478),
.B(n_466),
.Y(n_499)
);

INVx1_ASAP7_75t_L g522 ( 
.A(n_499),
.Y(n_522)
);

OR2x2_ASAP7_75t_L g518 ( 
.A(n_500),
.B(n_494),
.Y(n_518)
);

AOI21xp5_ASAP7_75t_L g501 ( 
.A1(n_483),
.A2(n_462),
.B(n_452),
.Y(n_501)
);

AOI21xp5_ASAP7_75t_L g517 ( 
.A1(n_501),
.A2(n_486),
.B(n_487),
.Y(n_517)
);

AOI22xp5_ASAP7_75t_SL g512 ( 
.A1(n_502),
.A2(n_472),
.B1(n_477),
.B2(n_482),
.Y(n_512)
);

NOR2xp33_ASAP7_75t_L g503 ( 
.A(n_479),
.B(n_259),
.Y(n_503)
);

INVx1_ASAP7_75t_L g523 ( 
.A(n_503),
.Y(n_523)
);

XOR2xp5_ASAP7_75t_L g504 ( 
.A(n_489),
.B(n_459),
.Y(n_504)
);

MAJIxp5_ASAP7_75t_L g505 ( 
.A(n_469),
.B(n_237),
.C(n_180),
.Y(n_505)
);

NOR2xp33_ASAP7_75t_L g506 ( 
.A(n_484),
.B(n_259),
.Y(n_506)
);

NOR2xp33_ASAP7_75t_SL g514 ( 
.A(n_506),
.B(n_507),
.Y(n_514)
);

BUFx24_ASAP7_75t_SL g507 ( 
.A(n_471),
.Y(n_507)
);

OAI21xp5_ASAP7_75t_SL g510 ( 
.A1(n_493),
.A2(n_488),
.B(n_490),
.Y(n_510)
);

AOI21xp5_ASAP7_75t_L g528 ( 
.A1(n_510),
.A2(n_513),
.B(n_515),
.Y(n_528)
);

OAI22xp5_ASAP7_75t_L g525 ( 
.A1(n_512),
.A2(n_491),
.B1(n_504),
.B2(n_215),
.Y(n_525)
);

MAJIxp5_ASAP7_75t_L g513 ( 
.A(n_495),
.B(n_489),
.C(n_475),
.Y(n_513)
);

MAJIxp5_ASAP7_75t_L g515 ( 
.A(n_498),
.B(n_475),
.C(n_470),
.Y(n_515)
);

INVx11_ASAP7_75t_L g516 ( 
.A(n_500),
.Y(n_516)
);

OR2x2_ASAP7_75t_L g532 ( 
.A(n_516),
.B(n_6),
.Y(n_532)
);

NAND2xp5_ASAP7_75t_SL g526 ( 
.A(n_517),
.B(n_518),
.Y(n_526)
);

HB1xp67_ASAP7_75t_L g519 ( 
.A(n_501),
.Y(n_519)
);

NAND2xp5_ASAP7_75t_L g527 ( 
.A(n_519),
.B(n_520),
.Y(n_527)
);

NOR2xp33_ASAP7_75t_SL g520 ( 
.A(n_505),
.B(n_482),
.Y(n_520)
);

MAJIxp5_ASAP7_75t_L g524 ( 
.A(n_511),
.B(n_508),
.C(n_497),
.Y(n_524)
);

NAND2xp5_ASAP7_75t_L g536 ( 
.A(n_524),
.B(n_530),
.Y(n_536)
);

INVxp67_ASAP7_75t_L g538 ( 
.A(n_525),
.Y(n_538)
);

AOI21xp5_ASAP7_75t_L g529 ( 
.A1(n_521),
.A2(n_491),
.B(n_206),
.Y(n_529)
);

OAI21xp5_ASAP7_75t_L g535 ( 
.A1(n_529),
.A2(n_531),
.B(n_534),
.Y(n_535)
);

NAND2xp5_ASAP7_75t_L g530 ( 
.A(n_509),
.B(n_0),
.Y(n_530)
);

AND2x2_ASAP7_75t_L g531 ( 
.A(n_521),
.B(n_197),
.Y(n_531)
);

NOR2xp33_ASAP7_75t_L g540 ( 
.A(n_532),
.B(n_533),
.Y(n_540)
);

NOR2xp33_ASAP7_75t_L g533 ( 
.A(n_514),
.B(n_0),
.Y(n_533)
);

OAI21xp5_ASAP7_75t_L g534 ( 
.A1(n_511),
.A2(n_0),
.B(n_2),
.Y(n_534)
);

MAJIxp5_ASAP7_75t_L g537 ( 
.A(n_528),
.B(n_522),
.C(n_513),
.Y(n_537)
);

NAND2xp5_ASAP7_75t_L g544 ( 
.A(n_537),
.B(n_541),
.Y(n_544)
);

AOI211xp5_ASAP7_75t_L g539 ( 
.A1(n_526),
.A2(n_523),
.B(n_516),
.C(n_512),
.Y(n_539)
);

CKINVDCx20_ASAP7_75t_R g542 ( 
.A(n_539),
.Y(n_542)
);

NOR2xp33_ASAP7_75t_L g541 ( 
.A(n_527),
.B(n_518),
.Y(n_541)
);

MAJIxp5_ASAP7_75t_L g543 ( 
.A(n_536),
.B(n_538),
.C(n_526),
.Y(n_543)
);

NOR2xp33_ASAP7_75t_L g546 ( 
.A(n_543),
.B(n_545),
.Y(n_546)
);

AOI21xp5_ASAP7_75t_L g545 ( 
.A1(n_538),
.A2(n_525),
.B(n_515),
.Y(n_545)
);

NOR2xp33_ASAP7_75t_L g547 ( 
.A(n_544),
.B(n_540),
.Y(n_547)
);

NOR2xp33_ASAP7_75t_L g548 ( 
.A(n_547),
.B(n_542),
.Y(n_548)
);

MAJIxp5_ASAP7_75t_L g549 ( 
.A(n_548),
.B(n_546),
.C(n_535),
.Y(n_549)
);

OAI21x1_ASAP7_75t_L g550 ( 
.A1(n_549),
.A2(n_517),
.B(n_5),
.Y(n_550)
);

OAI22xp5_ASAP7_75t_L g551 ( 
.A1(n_550),
.A2(n_6),
.B1(n_4),
.B2(n_5),
.Y(n_551)
);

AOI21xp5_ASAP7_75t_L g552 ( 
.A1(n_551),
.A2(n_4),
.B(n_5),
.Y(n_552)
);

AOI21xp5_ASAP7_75t_L g553 ( 
.A1(n_552),
.A2(n_6),
.B(n_551),
.Y(n_553)
);


endmodule