module real_jpeg_2606_n_17 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_16, n_3, n_10, n_9, n_17);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_16;
input n_3;
input n_10;
input n_9;

output n_17;

wire n_108;
wire n_54;
wire n_37;
wire n_168;
wire n_73;
wire n_38;
wire n_35;
wire n_29;
wire n_91;
wire n_49;
wire n_114;
wire n_201;
wire n_68;
wire n_146;
wire n_83;
wire n_78;
wire n_166;
wire n_176;
wire n_221;
wire n_215;
wire n_104;
wire n_153;
wire n_194;
wire n_161;
wire n_207;
wire n_64;
wire n_177;
wire n_47;
wire n_131;
wire n_163;
wire n_22;
wire n_174;
wire n_87;
wire n_197;
wire n_40;
wire n_105;
wire n_173;
wire n_115;
wire n_98;
wire n_27;
wire n_56;
wire n_184;
wire n_48;
wire n_164;
wire n_200;
wire n_140;
wire n_227;
wire n_126;
wire n_229;
wire n_214;
wire n_113;
wire n_120;
wire n_155;
wire n_199;
wire n_93;
wire n_95;
wire n_141;
wire n_65;
wire n_33;
wire n_139;
wire n_188;
wire n_142;
wire n_175;
wire n_76;
wire n_178;
wire n_67;
wire n_79;
wire n_107;
wire n_156;
wire n_147;
wire n_189;
wire n_170;
wire n_66;
wire n_231;
wire n_136;
wire n_28;
wire n_44;
wire n_208;
wire n_62;
wire n_162;
wire n_121;
wire n_106;
wire n_172;
wire n_160;
wire n_211;
wire n_45;
wire n_112;
wire n_42;
wire n_18;
wire n_145;
wire n_77;
wire n_109;
wire n_39;
wire n_219;
wire n_122;
wire n_94;
wire n_26;
wire n_19;
wire n_148;
wire n_222;
wire n_118;
wire n_220;
wire n_123;
wire n_116;
wire n_21;
wire n_50;
wire n_143;
wire n_196;
wire n_69;
wire n_186;
wire n_31;
wire n_137;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_218;
wire n_165;
wire n_134;
wire n_223;
wire n_72;
wire n_159;
wire n_171;
wire n_151;
wire n_183;
wire n_192;
wire n_203;
wire n_100;
wire n_198;
wire n_23;
wire n_51;
wire n_71;
wire n_90;
wire n_61;
wire n_110;
wire n_205;
wire n_195;
wire n_117;
wire n_99;
wire n_193;
wire n_86;
wire n_70;
wire n_41;
wire n_74;
wire n_80;
wire n_32;
wire n_20;
wire n_150;
wire n_228;
wire n_30;
wire n_158;
wire n_204;
wire n_149;
wire n_144;
wire n_130;
wire n_103;
wire n_225;
wire n_57;
wire n_43;
wire n_157;
wire n_84;
wire n_212;
wire n_82;
wire n_111;
wire n_132;
wire n_226;
wire n_125;
wire n_185;
wire n_55;
wire n_209;
wire n_180;
wire n_58;
wire n_52;
wire n_191;
wire n_63;
wire n_124;
wire n_24;
wire n_92;
wire n_75;
wire n_97;
wire n_187;
wire n_34;
wire n_190;
wire n_230;
wire n_60;
wire n_46;
wire n_169;
wire n_88;
wire n_59;
wire n_167;
wire n_128;
wire n_202;
wire n_179;
wire n_216;
wire n_213;
wire n_133;
wire n_138;
wire n_25;
wire n_217;
wire n_210;
wire n_127;
wire n_53;
wire n_206;
wire n_224;
wire n_119;
wire n_36;
wire n_81;
wire n_102;
wire n_85;
wire n_181;
wire n_101;
wire n_182;
wire n_96;
wire n_89;

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_0),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g33 ( 
.A(n_1),
.B(n_34),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g103 ( 
.A(n_1),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_L g150 ( 
.A(n_1),
.B(n_115),
.Y(n_150)
);

O2A1O1Ixp33_ASAP7_75t_L g166 ( 
.A1(n_1),
.A2(n_6),
.B(n_24),
.C(n_167),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_L g181 ( 
.A(n_1),
.B(n_55),
.Y(n_181)
);

AOI22xp5_ASAP7_75t_SL g190 ( 
.A1(n_1),
.A2(n_24),
.B1(n_25),
.B2(n_103),
.Y(n_190)
);

MAJIxp5_ASAP7_75t_L g199 ( 
.A(n_1),
.B(n_41),
.C(n_82),
.Y(n_199)
);

AOI22xp33_ASAP7_75t_L g201 ( 
.A1(n_1),
.A2(n_56),
.B1(n_57),
.B2(n_103),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_L g210 ( 
.A(n_1),
.B(n_46),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_L g215 ( 
.A(n_1),
.B(n_86),
.Y(n_215)
);

BUFx12f_ASAP7_75t_L g46 ( 
.A(n_2),
.Y(n_46)
);

OAI22xp5_ASAP7_75t_SL g48 ( 
.A1(n_3),
.A2(n_40),
.B1(n_41),
.B2(n_49),
.Y(n_48)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_3),
.Y(n_49)
);

OAI22xp5_ASAP7_75t_L g129 ( 
.A1(n_3),
.A2(n_49),
.B1(n_56),
.B2(n_57),
.Y(n_129)
);

OAI22xp5_ASAP7_75t_L g78 ( 
.A1(n_4),
.A2(n_56),
.B1(n_57),
.B2(n_79),
.Y(n_78)
);

CKINVDCx20_ASAP7_75t_R g79 ( 
.A(n_4),
.Y(n_79)
);

AOI22xp5_ASAP7_75t_SL g118 ( 
.A1(n_4),
.A2(n_24),
.B1(n_25),
.B2(n_79),
.Y(n_118)
);

AOI22xp33_ASAP7_75t_SL g152 ( 
.A1(n_4),
.A2(n_40),
.B1(n_41),
.B2(n_79),
.Y(n_152)
);

OAI22xp33_ASAP7_75t_SL g89 ( 
.A1(n_5),
.A2(n_40),
.B1(n_41),
.B2(n_90),
.Y(n_89)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_5),
.Y(n_90)
);

O2A1O1Ixp33_ASAP7_75t_L g53 ( 
.A1(n_6),
.A2(n_24),
.B(n_54),
.C(n_55),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_SL g54 ( 
.A(n_6),
.B(n_24),
.Y(n_54)
);

AO22x2_ASAP7_75t_L g55 ( 
.A1(n_6),
.A2(n_56),
.B1(n_57),
.B2(n_59),
.Y(n_55)
);

INVx5_ASAP7_75t_L g59 ( 
.A(n_6),
.Y(n_59)
);

OAI22xp5_ASAP7_75t_SL g61 ( 
.A1(n_7),
.A2(n_24),
.B1(n_25),
.B2(n_62),
.Y(n_61)
);

CKINVDCx20_ASAP7_75t_R g62 ( 
.A(n_7),
.Y(n_62)
);

OAI22xp5_ASAP7_75t_L g114 ( 
.A1(n_7),
.A2(n_30),
.B1(n_34),
.B2(n_62),
.Y(n_114)
);

AOI22xp5_ASAP7_75t_SL g162 ( 
.A1(n_7),
.A2(n_56),
.B1(n_57),
.B2(n_62),
.Y(n_162)
);

AOI22xp5_ASAP7_75t_SL g184 ( 
.A1(n_7),
.A2(n_40),
.B1(n_41),
.B2(n_62),
.Y(n_184)
);

INVx4_ASAP7_75t_L g32 ( 
.A(n_8),
.Y(n_32)
);

OAI22xp33_ASAP7_75t_SL g64 ( 
.A1(n_9),
.A2(n_24),
.B1(n_25),
.B2(n_65),
.Y(n_64)
);

CKINVDCx20_ASAP7_75t_R g65 ( 
.A(n_9),
.Y(n_65)
);

AOI22xp33_ASAP7_75t_L g73 ( 
.A1(n_9),
.A2(n_30),
.B1(n_34),
.B2(n_65),
.Y(n_73)
);

OAI22xp5_ASAP7_75t_SL g97 ( 
.A1(n_9),
.A2(n_56),
.B1(n_57),
.B2(n_65),
.Y(n_97)
);

AOI22xp33_ASAP7_75t_L g171 ( 
.A1(n_9),
.A2(n_40),
.B1(n_41),
.B2(n_65),
.Y(n_171)
);

AOI22xp33_ASAP7_75t_SL g126 ( 
.A1(n_10),
.A2(n_40),
.B1(n_41),
.B2(n_127),
.Y(n_126)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_10),
.Y(n_127)
);

BUFx10_ASAP7_75t_L g82 ( 
.A(n_11),
.Y(n_82)
);

INVx2_ASAP7_75t_L g27 ( 
.A(n_12),
.Y(n_27)
);

OAI22xp5_ASAP7_75t_L g68 ( 
.A1(n_13),
.A2(n_30),
.B1(n_34),
.B2(n_69),
.Y(n_68)
);

CKINVDCx20_ASAP7_75t_R g69 ( 
.A(n_13),
.Y(n_69)
);

OAI22xp33_ASAP7_75t_SL g99 ( 
.A1(n_13),
.A2(n_24),
.B1(n_25),
.B2(n_69),
.Y(n_99)
);

AOI22xp5_ASAP7_75t_SL g180 ( 
.A1(n_13),
.A2(n_56),
.B1(n_57),
.B2(n_69),
.Y(n_180)
);

OAI22xp5_ASAP7_75t_L g214 ( 
.A1(n_13),
.A2(n_40),
.B1(n_41),
.B2(n_69),
.Y(n_214)
);

AOI22xp33_ASAP7_75t_SL g39 ( 
.A1(n_14),
.A2(n_40),
.B1(n_41),
.B2(n_43),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_14),
.Y(n_43)
);

OAI22xp5_ASAP7_75t_L g85 ( 
.A1(n_14),
.A2(n_43),
.B1(n_56),
.B2(n_57),
.Y(n_85)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_15),
.Y(n_29)
);

BUFx12f_ASAP7_75t_L g58 ( 
.A(n_16),
.Y(n_58)
);

XOR2xp5_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_134),
.Y(n_17)
);

NAND2xp5_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_132),
.Y(n_18)
);

NAND2xp5_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_106),
.Y(n_19)
);

NOR2xp33_ASAP7_75t_SL g133 ( 
.A(n_20),
.B(n_106),
.Y(n_133)
);

MAJIxp5_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_76),
.C(n_91),
.Y(n_20)
);

XOR2xp5_ASAP7_75t_L g137 ( 
.A(n_21),
.B(n_138),
.Y(n_137)
);

XOR2xp5_ASAP7_75t_L g21 ( 
.A(n_22),
.B(n_50),
.Y(n_21)
);

MAJIxp5_ASAP7_75t_L g107 ( 
.A(n_22),
.B(n_51),
.C(n_66),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_L g22 ( 
.A(n_23),
.B(n_37),
.Y(n_22)
);

AOI22xp5_ASAP7_75t_L g144 ( 
.A1(n_23),
.A2(n_37),
.B1(n_38),
.B2(n_145),
.Y(n_144)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_23),
.Y(n_145)
);

AOI32xp33_ASAP7_75t_L g23 ( 
.A1(n_24),
.A2(n_28),
.A3(n_30),
.B1(n_33),
.B2(n_35),
.Y(n_23)
);

OA22x2_ASAP7_75t_L g70 ( 
.A1(n_24),
.A2(n_25),
.B1(n_28),
.B2(n_36),
.Y(n_70)
);

INVx4_ASAP7_75t_L g24 ( 
.A(n_25),
.Y(n_24)
);

NAND2xp33_ASAP7_75t_SL g35 ( 
.A(n_25),
.B(n_36),
.Y(n_35)
);

INVx11_ASAP7_75t_L g25 ( 
.A(n_26),
.Y(n_25)
);

BUFx12f_ASAP7_75t_L g26 ( 
.A(n_27),
.Y(n_26)
);

INVx3_ASAP7_75t_SL g36 ( 
.A(n_28),
.Y(n_36)
);

OAI22xp5_ASAP7_75t_SL g75 ( 
.A1(n_28),
.A2(n_30),
.B1(n_34),
.B2(n_36),
.Y(n_75)
);

INVx8_ASAP7_75t_L g28 ( 
.A(n_29),
.Y(n_28)
);

INVx2_ASAP7_75t_L g34 ( 
.A(n_30),
.Y(n_34)
);

O2A1O1Ixp33_ASAP7_75t_L g102 ( 
.A1(n_30),
.A2(n_103),
.B(n_104),
.C(n_105),
.Y(n_102)
);

BUFx4f_ASAP7_75t_L g30 ( 
.A(n_31),
.Y(n_30)
);

INVx4_ASAP7_75t_L g31 ( 
.A(n_32),
.Y(n_31)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_33),
.Y(n_104)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_38),
.Y(n_37)
);

OAI22xp5_ASAP7_75t_SL g38 ( 
.A1(n_39),
.A2(n_44),
.B1(n_45),
.B2(n_47),
.Y(n_38)
);

OAI22xp5_ASAP7_75t_SL g151 ( 
.A1(n_39),
.A2(n_44),
.B1(n_45),
.B2(n_152),
.Y(n_151)
);

OA22x2_ASAP7_75t_L g84 ( 
.A1(n_40),
.A2(n_41),
.B1(n_82),
.B2(n_83),
.Y(n_84)
);

INVx2_ASAP7_75t_SL g40 ( 
.A(n_41),
.Y(n_40)
);

NAND2xp5_ASAP7_75t_L g44 ( 
.A(n_41),
.B(n_45),
.Y(n_44)
);

NAND2xp5_ASAP7_75t_L g209 ( 
.A(n_41),
.B(n_210),
.Y(n_209)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_42),
.Y(n_41)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_44),
.Y(n_88)
);

OAI22xp5_ASAP7_75t_SL g124 ( 
.A1(n_44),
.A2(n_45),
.B1(n_125),
.B2(n_126),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_L g170 ( 
.A(n_44),
.B(n_171),
.Y(n_170)
);

OAI21xp5_ASAP7_75t_L g183 ( 
.A1(n_44),
.A2(n_184),
.B(n_185),
.Y(n_183)
);

OAI22xp5_ASAP7_75t_SL g218 ( 
.A1(n_44),
.A2(n_45),
.B1(n_184),
.B2(n_219),
.Y(n_218)
);

OAI21xp5_ASAP7_75t_L g168 ( 
.A1(n_45),
.A2(n_152),
.B(n_169),
.Y(n_168)
);

NOR2xp33_ASAP7_75t_L g186 ( 
.A(n_45),
.B(n_171),
.Y(n_186)
);

INVx4_ASAP7_75t_L g45 ( 
.A(n_46),
.Y(n_45)
);

AOI22xp5_ASAP7_75t_L g87 ( 
.A1(n_46),
.A2(n_48),
.B1(n_88),
.B2(n_89),
.Y(n_87)
);

AOI21xp5_ASAP7_75t_L g213 ( 
.A1(n_46),
.A2(n_170),
.B(n_214),
.Y(n_213)
);

CKINVDCx14_ASAP7_75t_R g47 ( 
.A(n_48),
.Y(n_47)
);

XNOR2xp5_ASAP7_75t_L g50 ( 
.A(n_51),
.B(n_66),
.Y(n_50)
);

OAI21xp5_ASAP7_75t_SL g51 ( 
.A1(n_52),
.A2(n_60),
.B(n_63),
.Y(n_51)
);

OAI21xp5_ASAP7_75t_SL g189 ( 
.A1(n_52),
.A2(n_63),
.B(n_190),
.Y(n_189)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_53),
.Y(n_52)
);

AOI22xp5_ASAP7_75t_L g98 ( 
.A1(n_53),
.A2(n_55),
.B1(n_61),
.B2(n_99),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g120 ( 
.A(n_53),
.B(n_64),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_L g63 ( 
.A(n_55),
.B(n_64),
.Y(n_63)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_55),
.Y(n_119)
);

OAI22xp33_ASAP7_75t_L g81 ( 
.A1(n_56),
.A2(n_57),
.B1(n_82),
.B2(n_83),
.Y(n_81)
);

OAI21xp33_ASAP7_75t_L g167 ( 
.A1(n_56),
.A2(n_59),
.B(n_103),
.Y(n_167)
);

INVx4_ASAP7_75t_L g56 ( 
.A(n_57),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_L g198 ( 
.A(n_57),
.B(n_199),
.Y(n_198)
);

BUFx12f_ASAP7_75t_L g57 ( 
.A(n_58),
.Y(n_57)
);

INVxp67_ASAP7_75t_L g60 ( 
.A(n_61),
.Y(n_60)
);

OAI21xp5_ASAP7_75t_L g66 ( 
.A1(n_67),
.A2(n_70),
.B(n_71),
.Y(n_66)
);

INVxp67_ASAP7_75t_L g67 ( 
.A(n_68),
.Y(n_67)
);

AOI22xp5_ASAP7_75t_L g113 ( 
.A1(n_68),
.A2(n_74),
.B1(n_114),
.B2(n_115),
.Y(n_113)
);

AND2x2_ASAP7_75t_SL g74 ( 
.A(n_70),
.B(n_75),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_70),
.B(n_73),
.Y(n_101)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_70),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_L g71 ( 
.A(n_72),
.B(n_74),
.Y(n_71)
);

INVxp67_ASAP7_75t_L g72 ( 
.A(n_73),
.Y(n_72)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_74),
.Y(n_105)
);

AOI22xp5_ASAP7_75t_SL g138 ( 
.A1(n_76),
.A2(n_91),
.B1(n_92),
.B2(n_139),
.Y(n_138)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_76),
.Y(n_139)
);

XNOR2xp5_ASAP7_75t_L g76 ( 
.A(n_77),
.B(n_87),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_SL g110 ( 
.A(n_77),
.B(n_87),
.Y(n_110)
);

AOI22xp5_ASAP7_75t_L g77 ( 
.A1(n_78),
.A2(n_80),
.B1(n_85),
.B2(n_86),
.Y(n_77)
);

CKINVDCx14_ASAP7_75t_R g95 ( 
.A(n_78),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_SL g96 ( 
.A(n_80),
.B(n_97),
.Y(n_96)
);

AOI22xp5_ASAP7_75t_L g128 ( 
.A1(n_80),
.A2(n_85),
.B1(n_86),
.B2(n_129),
.Y(n_128)
);

AOI21xp5_ASAP7_75t_L g160 ( 
.A1(n_80),
.A2(n_161),
.B(n_163),
.Y(n_160)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_80),
.Y(n_192)
);

AND2x2_ASAP7_75t_L g80 ( 
.A(n_81),
.B(n_84),
.Y(n_80)
);

INVx13_ASAP7_75t_L g83 ( 
.A(n_82),
.Y(n_83)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_84),
.Y(n_86)
);

OAI21xp5_ASAP7_75t_SL g94 ( 
.A1(n_84),
.A2(n_95),
.B(n_96),
.Y(n_94)
);

OAI21xp5_ASAP7_75t_L g179 ( 
.A1(n_84),
.A2(n_96),
.B(n_180),
.Y(n_179)
);

OAI22xp5_ASAP7_75t_SL g191 ( 
.A1(n_84),
.A2(n_162),
.B1(n_180),
.B2(n_192),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_L g164 ( 
.A(n_86),
.B(n_97),
.Y(n_164)
);

AOI21xp5_ASAP7_75t_L g211 ( 
.A1(n_88),
.A2(n_103),
.B(n_186),
.Y(n_211)
);

INVxp67_ASAP7_75t_L g125 ( 
.A(n_89),
.Y(n_125)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_92),
.Y(n_91)
);

MAJIxp5_ASAP7_75t_L g92 ( 
.A(n_93),
.B(n_98),
.C(n_100),
.Y(n_92)
);

AOI22xp5_ASAP7_75t_L g142 ( 
.A1(n_93),
.A2(n_94),
.B1(n_98),
.B2(n_143),
.Y(n_142)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_94),
.Y(n_93)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_98),
.Y(n_143)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_99),
.Y(n_148)
);

XNOR2xp5_ASAP7_75t_SL g141 ( 
.A(n_100),
.B(n_142),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_SL g100 ( 
.A(n_101),
.B(n_102),
.Y(n_100)
);

XOR2xp5_ASAP7_75t_L g106 ( 
.A(n_107),
.B(n_108),
.Y(n_106)
);

XNOR2xp5_ASAP7_75t_L g108 ( 
.A(n_109),
.B(n_123),
.Y(n_108)
);

AOI22xp5_ASAP7_75t_L g109 ( 
.A1(n_110),
.A2(n_111),
.B1(n_121),
.B2(n_122),
.Y(n_109)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_110),
.Y(n_121)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_111),
.Y(n_122)
);

AOI22xp5_ASAP7_75t_L g111 ( 
.A1(n_112),
.A2(n_113),
.B1(n_116),
.B2(n_117),
.Y(n_111)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_113),
.Y(n_112)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_117),
.Y(n_116)
);

OAI21xp5_ASAP7_75t_L g117 ( 
.A1(n_118),
.A2(n_119),
.B(n_120),
.Y(n_117)
);

OAI21xp5_ASAP7_75t_SL g147 ( 
.A1(n_119),
.A2(n_120),
.B(n_148),
.Y(n_147)
);

AOI22xp5_ASAP7_75t_L g123 ( 
.A1(n_124),
.A2(n_128),
.B1(n_130),
.B2(n_131),
.Y(n_123)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_124),
.Y(n_130)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_128),
.Y(n_131)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_133),
.Y(n_132)
);

OAI21xp5_ASAP7_75t_L g134 ( 
.A1(n_135),
.A2(n_153),
.B(n_231),
.Y(n_134)
);

INVxp67_ASAP7_75t_L g135 ( 
.A(n_136),
.Y(n_135)
);

OR2x2_ASAP7_75t_L g136 ( 
.A(n_137),
.B(n_140),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_L g231 ( 
.A(n_137),
.B(n_140),
.Y(n_231)
);

MAJIxp5_ASAP7_75t_L g140 ( 
.A(n_141),
.B(n_144),
.C(n_146),
.Y(n_140)
);

XOR2xp5_ASAP7_75t_L g172 ( 
.A(n_141),
.B(n_173),
.Y(n_172)
);

XNOR2xp5_ASAP7_75t_L g173 ( 
.A(n_144),
.B(n_146),
.Y(n_173)
);

MAJIxp5_ASAP7_75t_L g146 ( 
.A(n_147),
.B(n_149),
.C(n_151),
.Y(n_146)
);

XOR2xp5_ASAP7_75t_L g157 ( 
.A(n_147),
.B(n_158),
.Y(n_157)
);

AOI22xp5_ASAP7_75t_L g158 ( 
.A1(n_149),
.A2(n_150),
.B1(n_151),
.B2(n_159),
.Y(n_158)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_150),
.Y(n_149)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_151),
.Y(n_159)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_154),
.Y(n_153)
);

OAI21xp5_ASAP7_75t_L g154 ( 
.A1(n_155),
.A2(n_174),
.B(n_230),
.Y(n_154)
);

NOR2xp33_ASAP7_75t_L g155 ( 
.A(n_156),
.B(n_172),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_L g230 ( 
.A(n_156),
.B(n_172),
.Y(n_230)
);

MAJIxp5_ASAP7_75t_L g156 ( 
.A(n_157),
.B(n_160),
.C(n_165),
.Y(n_156)
);

XNOR2xp5_ASAP7_75t_L g226 ( 
.A(n_157),
.B(n_227),
.Y(n_226)
);

XNOR2xp5_ASAP7_75t_L g227 ( 
.A(n_160),
.B(n_165),
.Y(n_227)
);

INVxp67_ASAP7_75t_L g161 ( 
.A(n_162),
.Y(n_161)
);

INVxp67_ASAP7_75t_L g163 ( 
.A(n_164),
.Y(n_163)
);

OAI21xp5_ASAP7_75t_SL g200 ( 
.A1(n_164),
.A2(n_192),
.B(n_201),
.Y(n_200)
);

NAND2xp5_ASAP7_75t_L g165 ( 
.A(n_166),
.B(n_168),
.Y(n_165)
);

XOR2xp5_ASAP7_75t_L g193 ( 
.A(n_166),
.B(n_168),
.Y(n_193)
);

INVxp67_ASAP7_75t_L g169 ( 
.A(n_170),
.Y(n_169)
);

AOI21xp5_ASAP7_75t_SL g174 ( 
.A1(n_175),
.A2(n_225),
.B(n_229),
.Y(n_174)
);

OAI21xp5_ASAP7_75t_L g175 ( 
.A1(n_176),
.A2(n_194),
.B(n_224),
.Y(n_175)
);

NOR2xp33_ASAP7_75t_L g176 ( 
.A(n_177),
.B(n_187),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_L g224 ( 
.A(n_177),
.B(n_187),
.Y(n_224)
);

MAJIxp5_ASAP7_75t_L g177 ( 
.A(n_178),
.B(n_181),
.C(n_182),
.Y(n_177)
);

AOI22xp5_ASAP7_75t_L g203 ( 
.A1(n_178),
.A2(n_179),
.B1(n_181),
.B2(n_204),
.Y(n_203)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_179),
.Y(n_178)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_181),
.Y(n_204)
);

AOI22xp5_ASAP7_75t_L g202 ( 
.A1(n_182),
.A2(n_183),
.B1(n_203),
.B2(n_205),
.Y(n_202)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_183),
.Y(n_182)
);

INVxp67_ASAP7_75t_L g185 ( 
.A(n_186),
.Y(n_185)
);

XNOR2xp5_ASAP7_75t_L g187 ( 
.A(n_188),
.B(n_193),
.Y(n_187)
);

XNOR2xp5_ASAP7_75t_L g188 ( 
.A(n_189),
.B(n_191),
.Y(n_188)
);

MAJIxp5_ASAP7_75t_L g228 ( 
.A(n_189),
.B(n_191),
.C(n_193),
.Y(n_228)
);

AOI21xp5_ASAP7_75t_L g194 ( 
.A1(n_195),
.A2(n_206),
.B(n_223),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_L g195 ( 
.A(n_196),
.B(n_202),
.Y(n_195)
);

NOR2xp33_ASAP7_75t_L g223 ( 
.A(n_196),
.B(n_202),
.Y(n_223)
);

NAND2xp5_ASAP7_75t_L g196 ( 
.A(n_197),
.B(n_200),
.Y(n_196)
);

OAI22xp5_ASAP7_75t_SL g220 ( 
.A1(n_197),
.A2(n_198),
.B1(n_200),
.B2(n_221),
.Y(n_220)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_198),
.Y(n_197)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_200),
.Y(n_221)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_203),
.Y(n_205)
);

OAI21xp5_ASAP7_75t_L g206 ( 
.A1(n_207),
.A2(n_217),
.B(n_222),
.Y(n_206)
);

AOI21xp5_ASAP7_75t_L g207 ( 
.A1(n_208),
.A2(n_212),
.B(n_216),
.Y(n_207)
);

NOR2xp33_ASAP7_75t_L g208 ( 
.A(n_209),
.B(n_211),
.Y(n_208)
);

NAND2xp5_ASAP7_75t_SL g212 ( 
.A(n_213),
.B(n_215),
.Y(n_212)
);

NOR2xp33_ASAP7_75t_L g216 ( 
.A(n_213),
.B(n_215),
.Y(n_216)
);

INVxp67_ASAP7_75t_L g219 ( 
.A(n_214),
.Y(n_219)
);

NOR2xp33_ASAP7_75t_L g217 ( 
.A(n_218),
.B(n_220),
.Y(n_217)
);

NAND2xp5_ASAP7_75t_L g222 ( 
.A(n_218),
.B(n_220),
.Y(n_222)
);

NAND2xp5_ASAP7_75t_SL g225 ( 
.A(n_226),
.B(n_228),
.Y(n_225)
);

NOR2xp33_ASAP7_75t_L g229 ( 
.A(n_226),
.B(n_228),
.Y(n_229)
);


endmodule