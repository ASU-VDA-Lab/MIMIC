module fake_jpeg_15861_n_344 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_344);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_344;

wire n_253;
wire n_330;
wire n_158;
wire n_73;
wire n_152;
wire n_252;
wire n_19;
wire n_182;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_340;
wire n_291;
wire n_236;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_260;
wire n_199;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_247;
wire n_157;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_8),
.Y(n_16)
);

INVx8_ASAP7_75t_SL g17 ( 
.A(n_13),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_9),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_6),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_8),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_3),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_10),
.Y(n_22)
);

INVx6_ASAP7_75t_L g23 ( 
.A(n_9),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_5),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_10),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_1),
.Y(n_26)
);

INVx3_ASAP7_75t_L g27 ( 
.A(n_13),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_3),
.Y(n_28)
);

INVx2_ASAP7_75t_L g29 ( 
.A(n_6),
.Y(n_29)
);

BUFx8_ASAP7_75t_L g30 ( 
.A(n_8),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_2),
.Y(n_31)
);

INVx2_ASAP7_75t_L g32 ( 
.A(n_5),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_7),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_3),
.Y(n_34)
);

INVx1_ASAP7_75t_SL g35 ( 
.A(n_6),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_21),
.Y(n_36)
);

INVx3_ASAP7_75t_SL g62 ( 
.A(n_36),
.Y(n_62)
);

OR2x2_ASAP7_75t_L g37 ( 
.A(n_16),
.B(n_0),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_SL g67 ( 
.A(n_37),
.B(n_47),
.Y(n_67)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_29),
.Y(n_38)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_38),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_L g39 ( 
.A(n_29),
.B(n_0),
.Y(n_39)
);

AND2x2_ASAP7_75t_L g53 ( 
.A(n_39),
.B(n_44),
.Y(n_53)
);

BUFx24_ASAP7_75t_L g40 ( 
.A(n_30),
.Y(n_40)
);

INVx3_ASAP7_75t_SL g75 ( 
.A(n_40),
.Y(n_75)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_21),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_41),
.Y(n_59)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_18),
.Y(n_42)
);

NAND2xp5_ASAP7_75t_SL g74 ( 
.A(n_42),
.B(n_45),
.Y(n_74)
);

BUFx3_ASAP7_75t_L g43 ( 
.A(n_21),
.Y(n_43)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_43),
.Y(n_73)
);

AND2x2_ASAP7_75t_SL g44 ( 
.A(n_26),
.B(n_0),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_18),
.Y(n_45)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_29),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_L g54 ( 
.A(n_46),
.B(n_32),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g47 ( 
.A(n_35),
.B(n_15),
.Y(n_47)
);

CKINVDCx16_ASAP7_75t_R g48 ( 
.A(n_26),
.Y(n_48)
);

BUFx2_ASAP7_75t_L g77 ( 
.A(n_48),
.Y(n_77)
);

BUFx12_ASAP7_75t_L g49 ( 
.A(n_30),
.Y(n_49)
);

BUFx12f_ASAP7_75t_L g52 ( 
.A(n_49),
.Y(n_52)
);

INVx6_ASAP7_75t_L g50 ( 
.A(n_36),
.Y(n_50)
);

INVx2_ASAP7_75t_L g78 ( 
.A(n_50),
.Y(n_78)
);

AOI22xp33_ASAP7_75t_SL g51 ( 
.A1(n_38),
.A2(n_23),
.B1(n_27),
.B2(n_35),
.Y(n_51)
);

AOI22xp33_ASAP7_75t_SL g95 ( 
.A1(n_51),
.A2(n_64),
.B1(n_66),
.B2(n_71),
.Y(n_95)
);

AND2x2_ASAP7_75t_L g94 ( 
.A(n_54),
.B(n_63),
.Y(n_94)
);

BUFx10_ASAP7_75t_L g55 ( 
.A(n_40),
.Y(n_55)
);

HB1xp67_ASAP7_75t_L g104 ( 
.A(n_55),
.Y(n_104)
);

INVx5_ASAP7_75t_L g56 ( 
.A(n_43),
.Y(n_56)
);

INVx3_ASAP7_75t_L g87 ( 
.A(n_56),
.Y(n_87)
);

OAI22xp5_ASAP7_75t_L g57 ( 
.A1(n_39),
.A2(n_23),
.B1(n_32),
.B2(n_27),
.Y(n_57)
);

AOI22xp5_ASAP7_75t_L g114 ( 
.A1(n_57),
.A2(n_25),
.B1(n_1),
.B2(n_2),
.Y(n_114)
);

INVx6_ASAP7_75t_L g58 ( 
.A(n_36),
.Y(n_58)
);

INVx2_ASAP7_75t_L g85 ( 
.A(n_58),
.Y(n_85)
);

AOI22xp33_ASAP7_75t_L g60 ( 
.A1(n_48),
.A2(n_23),
.B1(n_27),
.B2(n_32),
.Y(n_60)
);

OAI22xp5_ASAP7_75t_SL g91 ( 
.A1(n_60),
.A2(n_69),
.B1(n_45),
.B2(n_42),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_L g63 ( 
.A(n_44),
.B(n_34),
.Y(n_63)
);

AOI22xp33_ASAP7_75t_SL g64 ( 
.A1(n_38),
.A2(n_23),
.B1(n_35),
.B2(n_18),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_36),
.Y(n_65)
);

CKINVDCx20_ASAP7_75t_R g81 ( 
.A(n_65),
.Y(n_81)
);

AOI22xp33_ASAP7_75t_SL g66 ( 
.A1(n_46),
.A2(n_22),
.B1(n_16),
.B2(n_31),
.Y(n_66)
);

INVx3_ASAP7_75t_L g68 ( 
.A(n_41),
.Y(n_68)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_68),
.Y(n_83)
);

AOI22xp33_ASAP7_75t_L g69 ( 
.A1(n_46),
.A2(n_22),
.B1(n_16),
.B2(n_31),
.Y(n_69)
);

INVx3_ASAP7_75t_L g70 ( 
.A(n_41),
.Y(n_70)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_70),
.Y(n_86)
);

AOI22xp33_ASAP7_75t_SL g71 ( 
.A1(n_42),
.A2(n_22),
.B1(n_19),
.B2(n_31),
.Y(n_71)
);

INVx4_ASAP7_75t_L g72 ( 
.A(n_41),
.Y(n_72)
);

INVx2_ASAP7_75t_L g89 ( 
.A(n_72),
.Y(n_89)
);

BUFx6f_ASAP7_75t_L g76 ( 
.A(n_43),
.Y(n_76)
);

CKINVDCx20_ASAP7_75t_R g84 ( 
.A(n_76),
.Y(n_84)
);

CKINVDCx20_ASAP7_75t_R g79 ( 
.A(n_61),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g122 ( 
.A(n_79),
.B(n_106),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_L g80 ( 
.A(n_53),
.B(n_44),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_L g121 ( 
.A(n_80),
.B(n_88),
.Y(n_121)
);

INVx2_ASAP7_75t_SL g82 ( 
.A(n_55),
.Y(n_82)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_82),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_L g88 ( 
.A(n_53),
.B(n_44),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_SL g90 ( 
.A(n_67),
.B(n_37),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_SL g135 ( 
.A(n_90),
.B(n_105),
.Y(n_135)
);

AOI22xp33_ASAP7_75t_L g116 ( 
.A1(n_91),
.A2(n_98),
.B1(n_68),
.B2(n_75),
.Y(n_116)
);

OAI22xp5_ASAP7_75t_SL g92 ( 
.A1(n_54),
.A2(n_39),
.B1(n_34),
.B2(n_26),
.Y(n_92)
);

OAI22xp5_ASAP7_75t_L g120 ( 
.A1(n_92),
.A2(n_96),
.B1(n_101),
.B2(n_114),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_L g93 ( 
.A(n_53),
.B(n_44),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_L g126 ( 
.A(n_93),
.B(n_97),
.Y(n_126)
);

OAI22xp5_ASAP7_75t_SL g96 ( 
.A1(n_57),
.A2(n_34),
.B1(n_24),
.B2(n_28),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g97 ( 
.A(n_63),
.B(n_37),
.Y(n_97)
);

AOI22xp33_ASAP7_75t_L g98 ( 
.A1(n_50),
.A2(n_45),
.B1(n_24),
.B2(n_19),
.Y(n_98)
);

OAI22xp33_ASAP7_75t_SL g99 ( 
.A1(n_58),
.A2(n_24),
.B1(n_19),
.B2(n_20),
.Y(n_99)
);

OAI22xp33_ASAP7_75t_SL g136 ( 
.A1(n_99),
.A2(n_102),
.B1(n_25),
.B2(n_30),
.Y(n_136)
);

OR2x2_ASAP7_75t_SL g100 ( 
.A(n_67),
.B(n_47),
.Y(n_100)
);

OAI21xp33_ASAP7_75t_L g117 ( 
.A1(n_100),
.A2(n_97),
.B(n_93),
.Y(n_117)
);

OAI22xp5_ASAP7_75t_SL g101 ( 
.A1(n_61),
.A2(n_28),
.B1(n_20),
.B2(n_43),
.Y(n_101)
);

OAI22xp33_ASAP7_75t_SL g102 ( 
.A1(n_62),
.A2(n_20),
.B1(n_28),
.B2(n_25),
.Y(n_102)
);

INVx2_ASAP7_75t_L g103 ( 
.A(n_73),
.Y(n_103)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_103),
.Y(n_134)
);

A2O1A1Ixp33_ASAP7_75t_L g105 ( 
.A1(n_74),
.A2(n_37),
.B(n_17),
.C(n_30),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_SL g106 ( 
.A(n_73),
.B(n_11),
.Y(n_106)
);

INVx2_ASAP7_75t_L g107 ( 
.A(n_76),
.Y(n_107)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_107),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_SL g108 ( 
.A(n_52),
.B(n_11),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_L g141 ( 
.A(n_108),
.B(n_77),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_L g109 ( 
.A(n_62),
.B(n_21),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_109),
.B(n_110),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_L g110 ( 
.A(n_62),
.B(n_33),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_L g111 ( 
.A(n_72),
.B(n_70),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_L g128 ( 
.A(n_111),
.B(n_59),
.Y(n_128)
);

INVx2_ASAP7_75t_L g112 ( 
.A(n_56),
.Y(n_112)
);

INVx3_ASAP7_75t_L g137 ( 
.A(n_112),
.Y(n_137)
);

MAJIxp5_ASAP7_75t_L g113 ( 
.A(n_52),
.B(n_40),
.C(n_30),
.Y(n_113)
);

MAJIxp5_ASAP7_75t_L g115 ( 
.A(n_113),
.B(n_40),
.C(n_75),
.Y(n_115)
);

AND2x2_ASAP7_75t_L g159 ( 
.A(n_115),
.B(n_128),
.Y(n_159)
);

AO21x1_ASAP7_75t_SL g175 ( 
.A1(n_116),
.A2(n_117),
.B(n_136),
.Y(n_175)
);

INVx8_ASAP7_75t_L g118 ( 
.A(n_87),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_L g154 ( 
.A(n_118),
.B(n_123),
.Y(n_154)
);

AOI21xp5_ASAP7_75t_L g119 ( 
.A1(n_95),
.A2(n_40),
.B(n_52),
.Y(n_119)
);

OAI21xp5_ASAP7_75t_L g180 ( 
.A1(n_119),
.A2(n_139),
.B(n_145),
.Y(n_180)
);

INVxp67_ASAP7_75t_L g123 ( 
.A(n_112),
.Y(n_123)
);

OAI22xp5_ASAP7_75t_L g124 ( 
.A1(n_114),
.A2(n_65),
.B1(n_59),
.B2(n_75),
.Y(n_124)
);

AOI22xp5_ASAP7_75t_L g148 ( 
.A1(n_124),
.A2(n_78),
.B1(n_85),
.B2(n_81),
.Y(n_148)
);

CKINVDCx20_ASAP7_75t_R g125 ( 
.A(n_111),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_L g170 ( 
.A(n_125),
.B(n_131),
.Y(n_170)
);

BUFx6f_ASAP7_75t_L g129 ( 
.A(n_87),
.Y(n_129)
);

INVx2_ASAP7_75t_L g160 ( 
.A(n_129),
.Y(n_160)
);

AOI22xp5_ASAP7_75t_SL g130 ( 
.A1(n_100),
.A2(n_17),
.B1(n_25),
.B2(n_33),
.Y(n_130)
);

INVxp67_ASAP7_75t_L g174 ( 
.A(n_130),
.Y(n_174)
);

INVx1_ASAP7_75t_SL g131 ( 
.A(n_82),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_SL g133 ( 
.A(n_92),
.B(n_52),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_L g171 ( 
.A(n_133),
.B(n_33),
.Y(n_171)
);

INVxp67_ASAP7_75t_L g138 ( 
.A(n_89),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_L g178 ( 
.A(n_138),
.B(n_141),
.Y(n_178)
);

OAI21xp5_ASAP7_75t_L g139 ( 
.A1(n_80),
.A2(n_77),
.B(n_30),
.Y(n_139)
);

INVxp67_ASAP7_75t_L g142 ( 
.A(n_89),
.Y(n_142)
);

CKINVDCx16_ASAP7_75t_R g153 ( 
.A(n_142),
.Y(n_153)
);

AOI22xp5_ASAP7_75t_L g143 ( 
.A1(n_94),
.A2(n_10),
.B1(n_9),
.B2(n_15),
.Y(n_143)
);

OAI22xp5_ASAP7_75t_L g152 ( 
.A1(n_143),
.A2(n_78),
.B1(n_85),
.B2(n_105),
.Y(n_152)
);

INVx4_ASAP7_75t_L g144 ( 
.A(n_83),
.Y(n_144)
);

CKINVDCx16_ASAP7_75t_R g179 ( 
.A(n_144),
.Y(n_179)
);

AND2x2_ASAP7_75t_L g145 ( 
.A(n_88),
.B(n_0),
.Y(n_145)
);

CKINVDCx20_ASAP7_75t_R g146 ( 
.A(n_134),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_SL g186 ( 
.A(n_146),
.B(n_152),
.Y(n_186)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_134),
.Y(n_147)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_147),
.Y(n_182)
);

OAI22xp5_ASAP7_75t_SL g194 ( 
.A1(n_148),
.A2(n_151),
.B1(n_161),
.B2(n_144),
.Y(n_194)
);

MAJIxp5_ASAP7_75t_L g149 ( 
.A(n_121),
.B(n_113),
.C(n_94),
.Y(n_149)
);

MAJIxp5_ASAP7_75t_L g198 ( 
.A(n_149),
.B(n_157),
.C(n_163),
.Y(n_198)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_128),
.Y(n_150)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_150),
.Y(n_197)
);

OAI22xp5_ASAP7_75t_SL g151 ( 
.A1(n_125),
.A2(n_110),
.B1(n_109),
.B2(n_91),
.Y(n_151)
);

CKINVDCx20_ASAP7_75t_R g155 ( 
.A(n_140),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_SL g205 ( 
.A(n_155),
.B(n_132),
.Y(n_205)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_137),
.Y(n_156)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_156),
.Y(n_199)
);

MAJx2_ASAP7_75t_L g157 ( 
.A(n_121),
.B(n_94),
.C(n_96),
.Y(n_157)
);

AOI21xp5_ASAP7_75t_L g158 ( 
.A1(n_139),
.A2(n_83),
.B(n_86),
.Y(n_158)
);

OAI21xp5_ASAP7_75t_SL g191 ( 
.A1(n_158),
.A2(n_162),
.B(n_171),
.Y(n_191)
);

AOI22xp5_ASAP7_75t_L g161 ( 
.A1(n_120),
.A2(n_86),
.B1(n_81),
.B2(n_103),
.Y(n_161)
);

A2O1A1O1Ixp25_ASAP7_75t_L g162 ( 
.A1(n_145),
.A2(n_101),
.B(n_40),
.C(n_49),
.D(n_55),
.Y(n_162)
);

MAJIxp5_ASAP7_75t_L g163 ( 
.A(n_126),
.B(n_55),
.C(n_84),
.Y(n_163)
);

MAJIxp5_ASAP7_75t_L g164 ( 
.A(n_126),
.B(n_84),
.C(n_82),
.Y(n_164)
);

MAJIxp5_ASAP7_75t_L g206 ( 
.A(n_164),
.B(n_169),
.C(n_172),
.Y(n_206)
);

OAI22xp5_ASAP7_75t_L g165 ( 
.A1(n_133),
.A2(n_107),
.B1(n_33),
.B2(n_11),
.Y(n_165)
);

OAI22xp33_ASAP7_75t_SL g204 ( 
.A1(n_165),
.A2(n_131),
.B1(n_13),
.B2(n_15),
.Y(n_204)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_137),
.Y(n_166)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_166),
.Y(n_208)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_132),
.Y(n_167)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_167),
.Y(n_184)
);

INVx2_ASAP7_75t_L g168 ( 
.A(n_129),
.Y(n_168)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_168),
.Y(n_187)
);

XOR2xp5_ASAP7_75t_L g169 ( 
.A(n_145),
.B(n_49),
.Y(n_169)
);

XNOR2xp5_ASAP7_75t_L g172 ( 
.A(n_115),
.B(n_104),
.Y(n_172)
);

AND2x2_ASAP7_75t_L g173 ( 
.A(n_127),
.B(n_1),
.Y(n_173)
);

AOI22xp5_ASAP7_75t_SL g193 ( 
.A1(n_173),
.A2(n_118),
.B1(n_144),
.B2(n_131),
.Y(n_193)
);

AOI22xp5_ASAP7_75t_SL g176 ( 
.A1(n_119),
.A2(n_130),
.B1(n_120),
.B2(n_135),
.Y(n_176)
);

INVxp67_ASAP7_75t_L g200 ( 
.A(n_176),
.Y(n_200)
);

NAND2xp5_ASAP7_75t_L g177 ( 
.A(n_127),
.B(n_1),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_L g188 ( 
.A(n_177),
.B(n_143),
.Y(n_188)
);

CKINVDCx20_ASAP7_75t_R g181 ( 
.A(n_156),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_SL g229 ( 
.A(n_181),
.B(n_189),
.Y(n_229)
);

XNOR2xp5_ASAP7_75t_L g183 ( 
.A(n_172),
.B(n_141),
.Y(n_183)
);

MAJIxp5_ASAP7_75t_L g221 ( 
.A(n_183),
.B(n_195),
.C(n_201),
.Y(n_221)
);

INVx1_ASAP7_75t_SL g185 ( 
.A(n_176),
.Y(n_185)
);

NOR2xp33_ASAP7_75t_L g236 ( 
.A(n_185),
.B(n_194),
.Y(n_236)
);

NAND2xp5_ASAP7_75t_L g219 ( 
.A(n_188),
.B(n_212),
.Y(n_219)
);

NOR2xp33_ASAP7_75t_L g189 ( 
.A(n_154),
.B(n_118),
.Y(n_189)
);

CKINVDCx20_ASAP7_75t_R g190 ( 
.A(n_166),
.Y(n_190)
);

NAND2xp5_ASAP7_75t_SL g232 ( 
.A(n_190),
.B(n_192),
.Y(n_232)
);

CKINVDCx14_ASAP7_75t_R g192 ( 
.A(n_178),
.Y(n_192)
);

NOR2xp33_ASAP7_75t_SL g216 ( 
.A(n_193),
.B(n_202),
.Y(n_216)
);

XNOR2xp5_ASAP7_75t_L g195 ( 
.A(n_149),
.B(n_122),
.Y(n_195)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_160),
.Y(n_196)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_196),
.Y(n_223)
);

XNOR2xp5_ASAP7_75t_L g201 ( 
.A(n_180),
.B(n_122),
.Y(n_201)
);

NOR2xp33_ASAP7_75t_SL g202 ( 
.A(n_177),
.B(n_135),
.Y(n_202)
);

NAND2xp5_ASAP7_75t_L g203 ( 
.A(n_150),
.B(n_124),
.Y(n_203)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_203),
.Y(n_230)
);

OAI22xp5_ASAP7_75t_L g237 ( 
.A1(n_204),
.A2(n_12),
.B1(n_14),
.B2(n_6),
.Y(n_237)
);

CKINVDCx20_ASAP7_75t_R g222 ( 
.A(n_205),
.Y(n_222)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_160),
.Y(n_207)
);

NOR2xp33_ASAP7_75t_L g239 ( 
.A(n_207),
.B(n_214),
.Y(n_239)
);

OAI22xp5_ASAP7_75t_SL g209 ( 
.A1(n_161),
.A2(n_140),
.B1(n_129),
.B2(n_49),
.Y(n_209)
);

OAI22xp5_ASAP7_75t_L g218 ( 
.A1(n_209),
.A2(n_148),
.B1(n_179),
.B2(n_170),
.Y(n_218)
);

MAJIxp5_ASAP7_75t_L g210 ( 
.A(n_164),
.B(n_49),
.C(n_14),
.Y(n_210)
);

MAJIxp5_ASAP7_75t_L g235 ( 
.A(n_210),
.B(n_211),
.C(n_168),
.Y(n_235)
);

XOR2xp5_ASAP7_75t_L g211 ( 
.A(n_159),
.B(n_49),
.Y(n_211)
);

NAND2xp5_ASAP7_75t_L g212 ( 
.A(n_173),
.B(n_2),
.Y(n_212)
);

OAI211xp5_ASAP7_75t_SL g213 ( 
.A1(n_157),
.A2(n_2),
.B(n_3),
.C(n_4),
.Y(n_213)
);

OAI21x1_ASAP7_75t_L g215 ( 
.A1(n_213),
.A2(n_162),
.B(n_175),
.Y(n_215)
);

BUFx24_ASAP7_75t_SL g214 ( 
.A(n_173),
.Y(n_214)
);

NAND2xp5_ASAP7_75t_L g248 ( 
.A(n_215),
.B(n_226),
.Y(n_248)
);

AOI21xp5_ASAP7_75t_L g217 ( 
.A1(n_185),
.A2(n_180),
.B(n_174),
.Y(n_217)
);

AOI21xp5_ASAP7_75t_L g261 ( 
.A1(n_217),
.A2(n_233),
.B(n_238),
.Y(n_261)
);

AOI22xp5_ASAP7_75t_L g244 ( 
.A1(n_218),
.A2(n_242),
.B1(n_213),
.B2(n_186),
.Y(n_244)
);

OAI22xp5_ASAP7_75t_SL g220 ( 
.A1(n_200),
.A2(n_174),
.B1(n_158),
.B2(n_171),
.Y(n_220)
);

OAI22xp5_ASAP7_75t_SL g255 ( 
.A1(n_220),
.A2(n_225),
.B1(n_226),
.B2(n_215),
.Y(n_255)
);

FAx1_ASAP7_75t_SL g224 ( 
.A(n_198),
.B(n_169),
.CI(n_163),
.CON(n_224),
.SN(n_224)
);

XNOR2xp5_ASAP7_75t_L g258 ( 
.A(n_224),
.B(n_227),
.Y(n_258)
);

AOI22xp5_ASAP7_75t_L g225 ( 
.A1(n_200),
.A2(n_159),
.B1(n_175),
.B2(n_151),
.Y(n_225)
);

INVx1_ASAP7_75t_SL g226 ( 
.A(n_193),
.Y(n_226)
);

NAND2xp5_ASAP7_75t_L g227 ( 
.A(n_197),
.B(n_195),
.Y(n_227)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_227),
.Y(n_256)
);

INVxp67_ASAP7_75t_L g228 ( 
.A(n_209),
.Y(n_228)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_228),
.Y(n_257)
);

XOR2xp5_ASAP7_75t_L g231 ( 
.A(n_198),
.B(n_159),
.Y(n_231)
);

MAJIxp5_ASAP7_75t_L g247 ( 
.A(n_231),
.B(n_235),
.C(n_241),
.Y(n_247)
);

AND2x2_ASAP7_75t_L g233 ( 
.A(n_211),
.B(n_201),
.Y(n_233)
);

NAND2xp5_ASAP7_75t_L g234 ( 
.A(n_197),
.B(n_153),
.Y(n_234)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_234),
.Y(n_259)
);

CKINVDCx16_ASAP7_75t_R g253 ( 
.A(n_237),
.Y(n_253)
);

OAI21xp5_ASAP7_75t_SL g238 ( 
.A1(n_191),
.A2(n_4),
.B(n_5),
.Y(n_238)
);

NOR2xp33_ASAP7_75t_SL g240 ( 
.A(n_188),
.B(n_12),
.Y(n_240)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_240),
.Y(n_245)
);

MAJIxp5_ASAP7_75t_L g241 ( 
.A(n_206),
.B(n_12),
.C(n_14),
.Y(n_241)
);

OAI22xp5_ASAP7_75t_L g242 ( 
.A1(n_203),
.A2(n_4),
.B1(n_5),
.B2(n_7),
.Y(n_242)
);

XNOR2xp5_ASAP7_75t_SL g243 ( 
.A(n_221),
.B(n_183),
.Y(n_243)
);

XOR2xp5_ASAP7_75t_L g279 ( 
.A(n_243),
.B(n_249),
.Y(n_279)
);

OAI22xp5_ASAP7_75t_L g277 ( 
.A1(n_244),
.A2(n_216),
.B1(n_240),
.B2(n_212),
.Y(n_277)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_223),
.Y(n_246)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_246),
.Y(n_271)
);

XNOR2xp5_ASAP7_75t_SL g249 ( 
.A(n_221),
.B(n_206),
.Y(n_249)
);

CKINVDCx20_ASAP7_75t_R g250 ( 
.A(n_232),
.Y(n_250)
);

NAND2xp5_ASAP7_75t_SL g283 ( 
.A(n_250),
.B(n_266),
.Y(n_283)
);

XOR2xp5_ASAP7_75t_L g251 ( 
.A(n_231),
.B(n_191),
.Y(n_251)
);

MAJIxp5_ASAP7_75t_L g278 ( 
.A(n_251),
.B(n_254),
.C(n_258),
.Y(n_278)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_223),
.Y(n_252)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_252),
.Y(n_272)
);

MAJIxp5_ASAP7_75t_L g254 ( 
.A(n_224),
.B(n_210),
.C(n_194),
.Y(n_254)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_255),
.Y(n_286)
);

NOR2xp67_ASAP7_75t_SL g260 ( 
.A(n_222),
.B(n_184),
.Y(n_260)
);

OAI21xp5_ASAP7_75t_SL g270 ( 
.A1(n_260),
.A2(n_262),
.B(n_217),
.Y(n_270)
);

AOI21xp5_ASAP7_75t_L g262 ( 
.A1(n_236),
.A2(n_208),
.B(n_199),
.Y(n_262)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_234),
.Y(n_263)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_263),
.Y(n_276)
);

MAJIxp5_ASAP7_75t_L g264 ( 
.A(n_224),
.B(n_208),
.C(n_199),
.Y(n_264)
);

NOR2xp33_ASAP7_75t_L g280 ( 
.A(n_264),
.B(n_216),
.Y(n_280)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_229),
.Y(n_265)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_265),
.Y(n_282)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_230),
.Y(n_266)
);

OAI22xp5_ASAP7_75t_L g267 ( 
.A1(n_257),
.A2(n_230),
.B1(n_228),
.B2(n_259),
.Y(n_267)
);

AOI22xp5_ASAP7_75t_L g287 ( 
.A1(n_267),
.A2(n_277),
.B1(n_248),
.B2(n_233),
.Y(n_287)
);

NAND2xp5_ASAP7_75t_L g268 ( 
.A(n_259),
.B(n_222),
.Y(n_268)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_268),
.Y(n_293)
);

INVxp67_ASAP7_75t_L g269 ( 
.A(n_262),
.Y(n_269)
);

NAND2xp5_ASAP7_75t_L g298 ( 
.A(n_269),
.B(n_275),
.Y(n_298)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_270),
.Y(n_288)
);

NAND2xp5_ASAP7_75t_L g273 ( 
.A(n_256),
.B(n_219),
.Y(n_273)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_273),
.Y(n_302)
);

OAI22xp5_ASAP7_75t_SL g274 ( 
.A1(n_257),
.A2(n_225),
.B1(n_219),
.B2(n_235),
.Y(n_274)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_274),
.Y(n_295)
);

NAND2xp5_ASAP7_75t_L g275 ( 
.A(n_256),
.B(n_242),
.Y(n_275)
);

MAJIxp5_ASAP7_75t_L g292 ( 
.A(n_280),
.B(n_254),
.C(n_258),
.Y(n_292)
);

OAI21xp5_ASAP7_75t_L g281 ( 
.A1(n_248),
.A2(n_233),
.B(n_220),
.Y(n_281)
);

AO21x1_ASAP7_75t_L g291 ( 
.A1(n_281),
.A2(n_261),
.B(n_255),
.Y(n_291)
);

OAI22xp5_ASAP7_75t_L g284 ( 
.A1(n_253),
.A2(n_218),
.B1(n_241),
.B2(n_238),
.Y(n_284)
);

INVxp67_ASAP7_75t_L g294 ( 
.A(n_284),
.Y(n_294)
);

NOR2xp33_ASAP7_75t_L g285 ( 
.A(n_245),
.B(n_182),
.Y(n_285)
);

NOR2xp33_ASAP7_75t_L g290 ( 
.A(n_285),
.B(n_244),
.Y(n_290)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_287),
.Y(n_308)
);

NOR2xp67_ASAP7_75t_SL g289 ( 
.A(n_283),
.B(n_264),
.Y(n_289)
);

AOI21xp5_ASAP7_75t_L g312 ( 
.A1(n_289),
.A2(n_301),
.B(n_270),
.Y(n_312)
);

NOR2xp33_ASAP7_75t_SL g307 ( 
.A(n_290),
.B(n_292),
.Y(n_307)
);

XOR2xp5_ASAP7_75t_L g316 ( 
.A(n_291),
.B(n_275),
.Y(n_316)
);

XNOR2x1_ASAP7_75t_L g296 ( 
.A(n_281),
.B(n_261),
.Y(n_296)
);

XNOR2xp5_ASAP7_75t_SL g315 ( 
.A(n_296),
.B(n_274),
.Y(n_315)
);

INVx1_ASAP7_75t_SL g297 ( 
.A(n_269),
.Y(n_297)
);

NAND2xp5_ASAP7_75t_L g313 ( 
.A(n_297),
.B(n_299),
.Y(n_313)
);

NOR2xp33_ASAP7_75t_L g299 ( 
.A(n_282),
.B(n_187),
.Y(n_299)
);

INVx13_ASAP7_75t_L g300 ( 
.A(n_271),
.Y(n_300)
);

AOI22xp5_ASAP7_75t_L g306 ( 
.A1(n_300),
.A2(n_272),
.B1(n_267),
.B2(n_276),
.Y(n_306)
);

NAND2xp5_ASAP7_75t_L g301 ( 
.A(n_273),
.B(n_251),
.Y(n_301)
);

MAJIxp5_ASAP7_75t_L g303 ( 
.A(n_295),
.B(n_247),
.C(n_249),
.Y(n_303)
);

MAJIxp5_ASAP7_75t_L g321 ( 
.A(n_303),
.B(n_304),
.C(n_309),
.Y(n_321)
);

MAJIxp5_ASAP7_75t_L g304 ( 
.A(n_293),
.B(n_247),
.C(n_279),
.Y(n_304)
);

OAI21xp5_ASAP7_75t_SL g305 ( 
.A1(n_294),
.A2(n_282),
.B(n_271),
.Y(n_305)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_305),
.Y(n_320)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_306),
.Y(n_325)
);

MAJIxp5_ASAP7_75t_L g309 ( 
.A(n_293),
.B(n_279),
.C(n_278),
.Y(n_309)
);

MAJIxp5_ASAP7_75t_L g310 ( 
.A(n_301),
.B(n_292),
.C(n_278),
.Y(n_310)
);

NAND2xp5_ASAP7_75t_L g318 ( 
.A(n_310),
.B(n_311),
.Y(n_318)
);

NOR2xp33_ASAP7_75t_SL g311 ( 
.A(n_287),
.B(n_239),
.Y(n_311)
);

XOR2xp5_ASAP7_75t_L g324 ( 
.A(n_312),
.B(n_315),
.Y(n_324)
);

OAI21xp5_ASAP7_75t_L g314 ( 
.A1(n_294),
.A2(n_286),
.B(n_268),
.Y(n_314)
);

XNOR2xp5_ASAP7_75t_L g322 ( 
.A(n_314),
.B(n_298),
.Y(n_322)
);

XOR2xp5_ASAP7_75t_L g326 ( 
.A(n_316),
.B(n_291),
.Y(n_326)
);

AOI21xp5_ASAP7_75t_SL g317 ( 
.A1(n_308),
.A2(n_296),
.B(n_288),
.Y(n_317)
);

NAND2xp5_ASAP7_75t_L g327 ( 
.A(n_317),
.B(n_322),
.Y(n_327)
);

OAI22xp5_ASAP7_75t_SL g319 ( 
.A1(n_316),
.A2(n_286),
.B1(n_298),
.B2(n_276),
.Y(n_319)
);

MAJIxp5_ASAP7_75t_L g329 ( 
.A(n_319),
.B(n_326),
.C(n_315),
.Y(n_329)
);

NOR2xp33_ASAP7_75t_L g323 ( 
.A(n_307),
.B(n_297),
.Y(n_323)
);

NAND2xp5_ASAP7_75t_L g328 ( 
.A(n_323),
.B(n_313),
.Y(n_328)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_328),
.Y(n_335)
);

INVxp67_ASAP7_75t_L g334 ( 
.A(n_329),
.Y(n_334)
);

NAND2xp5_ASAP7_75t_L g330 ( 
.A(n_320),
.B(n_272),
.Y(n_330)
);

NAND2xp5_ASAP7_75t_L g336 ( 
.A(n_330),
.B(n_331),
.Y(n_336)
);

INVxp33_ASAP7_75t_L g331 ( 
.A(n_317),
.Y(n_331)
);

A2O1A1Ixp33_ASAP7_75t_L g332 ( 
.A1(n_318),
.A2(n_302),
.B(n_325),
.C(n_324),
.Y(n_332)
);

NAND2xp5_ASAP7_75t_L g337 ( 
.A(n_332),
.B(n_333),
.Y(n_337)
);

OAI21xp5_ASAP7_75t_SL g333 ( 
.A1(n_326),
.A2(n_302),
.B(n_309),
.Y(n_333)
);

AOI211x1_ASAP7_75t_L g338 ( 
.A1(n_337),
.A2(n_331),
.B(n_324),
.C(n_327),
.Y(n_338)
);

AOI21xp5_ASAP7_75t_L g340 ( 
.A1(n_338),
.A2(n_339),
.B(n_334),
.Y(n_340)
);

AND2x2_ASAP7_75t_L g339 ( 
.A(n_336),
.B(n_321),
.Y(n_339)
);

AOI321xp33_ASAP7_75t_L g341 ( 
.A1(n_340),
.A2(n_335),
.A3(n_321),
.B1(n_310),
.B2(n_304),
.C(n_303),
.Y(n_341)
);

MAJIxp5_ASAP7_75t_L g342 ( 
.A(n_341),
.B(n_243),
.C(n_300),
.Y(n_342)
);

AOI22xp5_ASAP7_75t_L g343 ( 
.A1(n_342),
.A2(n_4),
.B1(n_7),
.B2(n_8),
.Y(n_343)
);

XOR2xp5_ASAP7_75t_L g344 ( 
.A(n_343),
.B(n_7),
.Y(n_344)
);


endmodule