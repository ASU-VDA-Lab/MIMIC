module fake_ariane_1270_n_2532 (n_295, n_356, n_170, n_190, n_160, n_64, n_180, n_119, n_124, n_386, n_307, n_516, n_332, n_294, n_197, n_463, n_176, n_34, n_404, n_172, n_347, n_423, n_183, n_469, n_479, n_373, n_299, n_499, n_12, n_133, n_66, n_205, n_341, n_71, n_109, n_245, n_421, n_96, n_522, n_319, n_49, n_20, n_416, n_283, n_50, n_187, n_525, n_367, n_345, n_374, n_318, n_103, n_244, n_226, n_220, n_261, n_36, n_370, n_189, n_72, n_286, n_443, n_57, n_424, n_528, n_387, n_406, n_117, n_139, n_524, n_85, n_130, n_349, n_391, n_466, n_346, n_214, n_348, n_2, n_462, n_32, n_410, n_379, n_445, n_515, n_138, n_162, n_264, n_137, n_122, n_198, n_232, n_52, n_441, n_385, n_73, n_327, n_77, n_372, n_377, n_15, n_396, n_23, n_399, n_520, n_87, n_279, n_207, n_363, n_354, n_41, n_140, n_419, n_151, n_28, n_146, n_230, n_270, n_194, n_154, n_338, n_142, n_285, n_473, n_186, n_202, n_145, n_193, n_500, n_59, n_336, n_315, n_311, n_239, n_402, n_35, n_272, n_54, n_8, n_339, n_487, n_167, n_90, n_38, n_422, n_47, n_153, n_18, n_269, n_75, n_158, n_69, n_259, n_95, n_446, n_143, n_152, n_405, n_120, n_169, n_106, n_173, n_242, n_309, n_320, n_115, n_331, n_401, n_485, n_267, n_495, n_504, n_483, n_335, n_435, n_350, n_291, n_344, n_381, n_426, n_433, n_481, n_398, n_62, n_210, n_200, n_529, n_502, n_166, n_253, n_218, n_79, n_3, n_271, n_465, n_486, n_507, n_247, n_91, n_240, n_369, n_128, n_224, n_44, n_82, n_31, n_420, n_518, n_439, n_222, n_478, n_510, n_256, n_326, n_227, n_48, n_188, n_323, n_330, n_400, n_11, n_129, n_126, n_282, n_328, n_368, n_277, n_248, n_301, n_467, n_432, n_536, n_293, n_228, n_325, n_276, n_93, n_427, n_108, n_497, n_303, n_442, n_168, n_81, n_1, n_206, n_352, n_511, n_238, n_365, n_429, n_455, n_136, n_334, n_192, n_488, n_300, n_533, n_505, n_14, n_163, n_88, n_141, n_390, n_498, n_104, n_501, n_438, n_314, n_16, n_440, n_273, n_305, n_312, n_233, n_56, n_60, n_388, n_333, n_449, n_413, n_392, n_376, n_512, n_459, n_221, n_321, n_86, n_361, n_458, n_89, n_149, n_383, n_237, n_175, n_453, n_74, n_491, n_19, n_40, n_181, n_53, n_260, n_362, n_310, n_236, n_281, n_24, n_7, n_461, n_209, n_262, n_490, n_17, n_225, n_235, n_464, n_297, n_503, n_290, n_527, n_46, n_84, n_371, n_199, n_107, n_217, n_452, n_178, n_42, n_308, n_417, n_201, n_70, n_343, n_10, n_414, n_287, n_302, n_380, n_6, n_94, n_284, n_4, n_448, n_249, n_534, n_37, n_58, n_65, n_123, n_212, n_355, n_444, n_278, n_255, n_450, n_257, n_148, n_451, n_475, n_135, n_409, n_171, n_519, n_384, n_468, n_61, n_526, n_102, n_182, n_482, n_316, n_196, n_125, n_43, n_407, n_13, n_27, n_254, n_476, n_460, n_219, n_55, n_535, n_231, n_366, n_234, n_492, n_280, n_215, n_252, n_161, n_454, n_298, n_532, n_68, n_415, n_78, n_63, n_99, n_216, n_5, n_514, n_418, n_223, n_403, n_25, n_83, n_389, n_513, n_288, n_179, n_395, n_195, n_213, n_110, n_304, n_67, n_509, n_306, n_313, n_92, n_430, n_493, n_203, n_378, n_436, n_150, n_98, n_375, n_113, n_114, n_33, n_324, n_337, n_437, n_111, n_21, n_274, n_472, n_296, n_265, n_208, n_456, n_156, n_292, n_174, n_275, n_100, n_132, n_147, n_204, n_521, n_51, n_496, n_76, n_342, n_26, n_246, n_517, n_530, n_0, n_428, n_159, n_358, n_105, n_30, n_494, n_131, n_263, n_434, n_360, n_229, n_394, n_250, n_165, n_144, n_317, n_101, n_243, n_134, n_329, n_185, n_340, n_289, n_9, n_112, n_45, n_523, n_268, n_266, n_470, n_457, n_164, n_157, n_184, n_177, n_477, n_364, n_258, n_425, n_431, n_508, n_118, n_121, n_411, n_484, n_353, n_22, n_241, n_29, n_357, n_412, n_447, n_191, n_382, n_489, n_80, n_480, n_211, n_97, n_408, n_322, n_251, n_506, n_116, n_397, n_471, n_351, n_39, n_393, n_474, n_359, n_155, n_127, n_531, n_2532);

input n_295;
input n_356;
input n_170;
input n_190;
input n_160;
input n_64;
input n_180;
input n_119;
input n_124;
input n_386;
input n_307;
input n_516;
input n_332;
input n_294;
input n_197;
input n_463;
input n_176;
input n_34;
input n_404;
input n_172;
input n_347;
input n_423;
input n_183;
input n_469;
input n_479;
input n_373;
input n_299;
input n_499;
input n_12;
input n_133;
input n_66;
input n_205;
input n_341;
input n_71;
input n_109;
input n_245;
input n_421;
input n_96;
input n_522;
input n_319;
input n_49;
input n_20;
input n_416;
input n_283;
input n_50;
input n_187;
input n_525;
input n_367;
input n_345;
input n_374;
input n_318;
input n_103;
input n_244;
input n_226;
input n_220;
input n_261;
input n_36;
input n_370;
input n_189;
input n_72;
input n_286;
input n_443;
input n_57;
input n_424;
input n_528;
input n_387;
input n_406;
input n_117;
input n_139;
input n_524;
input n_85;
input n_130;
input n_349;
input n_391;
input n_466;
input n_346;
input n_214;
input n_348;
input n_2;
input n_462;
input n_32;
input n_410;
input n_379;
input n_445;
input n_515;
input n_138;
input n_162;
input n_264;
input n_137;
input n_122;
input n_198;
input n_232;
input n_52;
input n_441;
input n_385;
input n_73;
input n_327;
input n_77;
input n_372;
input n_377;
input n_15;
input n_396;
input n_23;
input n_399;
input n_520;
input n_87;
input n_279;
input n_207;
input n_363;
input n_354;
input n_41;
input n_140;
input n_419;
input n_151;
input n_28;
input n_146;
input n_230;
input n_270;
input n_194;
input n_154;
input n_338;
input n_142;
input n_285;
input n_473;
input n_186;
input n_202;
input n_145;
input n_193;
input n_500;
input n_59;
input n_336;
input n_315;
input n_311;
input n_239;
input n_402;
input n_35;
input n_272;
input n_54;
input n_8;
input n_339;
input n_487;
input n_167;
input n_90;
input n_38;
input n_422;
input n_47;
input n_153;
input n_18;
input n_269;
input n_75;
input n_158;
input n_69;
input n_259;
input n_95;
input n_446;
input n_143;
input n_152;
input n_405;
input n_120;
input n_169;
input n_106;
input n_173;
input n_242;
input n_309;
input n_320;
input n_115;
input n_331;
input n_401;
input n_485;
input n_267;
input n_495;
input n_504;
input n_483;
input n_335;
input n_435;
input n_350;
input n_291;
input n_344;
input n_381;
input n_426;
input n_433;
input n_481;
input n_398;
input n_62;
input n_210;
input n_200;
input n_529;
input n_502;
input n_166;
input n_253;
input n_218;
input n_79;
input n_3;
input n_271;
input n_465;
input n_486;
input n_507;
input n_247;
input n_91;
input n_240;
input n_369;
input n_128;
input n_224;
input n_44;
input n_82;
input n_31;
input n_420;
input n_518;
input n_439;
input n_222;
input n_478;
input n_510;
input n_256;
input n_326;
input n_227;
input n_48;
input n_188;
input n_323;
input n_330;
input n_400;
input n_11;
input n_129;
input n_126;
input n_282;
input n_328;
input n_368;
input n_277;
input n_248;
input n_301;
input n_467;
input n_432;
input n_536;
input n_293;
input n_228;
input n_325;
input n_276;
input n_93;
input n_427;
input n_108;
input n_497;
input n_303;
input n_442;
input n_168;
input n_81;
input n_1;
input n_206;
input n_352;
input n_511;
input n_238;
input n_365;
input n_429;
input n_455;
input n_136;
input n_334;
input n_192;
input n_488;
input n_300;
input n_533;
input n_505;
input n_14;
input n_163;
input n_88;
input n_141;
input n_390;
input n_498;
input n_104;
input n_501;
input n_438;
input n_314;
input n_16;
input n_440;
input n_273;
input n_305;
input n_312;
input n_233;
input n_56;
input n_60;
input n_388;
input n_333;
input n_449;
input n_413;
input n_392;
input n_376;
input n_512;
input n_459;
input n_221;
input n_321;
input n_86;
input n_361;
input n_458;
input n_89;
input n_149;
input n_383;
input n_237;
input n_175;
input n_453;
input n_74;
input n_491;
input n_19;
input n_40;
input n_181;
input n_53;
input n_260;
input n_362;
input n_310;
input n_236;
input n_281;
input n_24;
input n_7;
input n_461;
input n_209;
input n_262;
input n_490;
input n_17;
input n_225;
input n_235;
input n_464;
input n_297;
input n_503;
input n_290;
input n_527;
input n_46;
input n_84;
input n_371;
input n_199;
input n_107;
input n_217;
input n_452;
input n_178;
input n_42;
input n_308;
input n_417;
input n_201;
input n_70;
input n_343;
input n_10;
input n_414;
input n_287;
input n_302;
input n_380;
input n_6;
input n_94;
input n_284;
input n_4;
input n_448;
input n_249;
input n_534;
input n_37;
input n_58;
input n_65;
input n_123;
input n_212;
input n_355;
input n_444;
input n_278;
input n_255;
input n_450;
input n_257;
input n_148;
input n_451;
input n_475;
input n_135;
input n_409;
input n_171;
input n_519;
input n_384;
input n_468;
input n_61;
input n_526;
input n_102;
input n_182;
input n_482;
input n_316;
input n_196;
input n_125;
input n_43;
input n_407;
input n_13;
input n_27;
input n_254;
input n_476;
input n_460;
input n_219;
input n_55;
input n_535;
input n_231;
input n_366;
input n_234;
input n_492;
input n_280;
input n_215;
input n_252;
input n_161;
input n_454;
input n_298;
input n_532;
input n_68;
input n_415;
input n_78;
input n_63;
input n_99;
input n_216;
input n_5;
input n_514;
input n_418;
input n_223;
input n_403;
input n_25;
input n_83;
input n_389;
input n_513;
input n_288;
input n_179;
input n_395;
input n_195;
input n_213;
input n_110;
input n_304;
input n_67;
input n_509;
input n_306;
input n_313;
input n_92;
input n_430;
input n_493;
input n_203;
input n_378;
input n_436;
input n_150;
input n_98;
input n_375;
input n_113;
input n_114;
input n_33;
input n_324;
input n_337;
input n_437;
input n_111;
input n_21;
input n_274;
input n_472;
input n_296;
input n_265;
input n_208;
input n_456;
input n_156;
input n_292;
input n_174;
input n_275;
input n_100;
input n_132;
input n_147;
input n_204;
input n_521;
input n_51;
input n_496;
input n_76;
input n_342;
input n_26;
input n_246;
input n_517;
input n_530;
input n_0;
input n_428;
input n_159;
input n_358;
input n_105;
input n_30;
input n_494;
input n_131;
input n_263;
input n_434;
input n_360;
input n_229;
input n_394;
input n_250;
input n_165;
input n_144;
input n_317;
input n_101;
input n_243;
input n_134;
input n_329;
input n_185;
input n_340;
input n_289;
input n_9;
input n_112;
input n_45;
input n_523;
input n_268;
input n_266;
input n_470;
input n_457;
input n_164;
input n_157;
input n_184;
input n_177;
input n_477;
input n_364;
input n_258;
input n_425;
input n_431;
input n_508;
input n_118;
input n_121;
input n_411;
input n_484;
input n_353;
input n_22;
input n_241;
input n_29;
input n_357;
input n_412;
input n_447;
input n_191;
input n_382;
input n_489;
input n_80;
input n_480;
input n_211;
input n_97;
input n_408;
input n_322;
input n_251;
input n_506;
input n_116;
input n_397;
input n_471;
input n_351;
input n_39;
input n_393;
input n_474;
input n_359;
input n_155;
input n_127;
input n_531;

output n_2532;

wire n_913;
wire n_1681;
wire n_2163;
wire n_1486;
wire n_1507;
wire n_1938;
wire n_589;
wire n_2484;
wire n_1174;
wire n_2346;
wire n_1469;
wire n_691;
wire n_1353;
wire n_1355;
wire n_2131;
wire n_2500;
wire n_2509;
wire n_1383;
wire n_2182;
wire n_603;
wire n_2135;
wire n_2334;
wire n_1250;
wire n_2030;
wire n_1169;
wire n_789;
wire n_850;
wire n_1916;
wire n_610;
wire n_1713;
wire n_1436;
wire n_2407;
wire n_690;
wire n_1109;
wire n_1430;
wire n_2002;
wire n_1463;
wire n_2243;
wire n_1238;
wire n_2011;
wire n_1515;
wire n_817;
wire n_1837;
wire n_924;
wire n_781;
wire n_2013;
wire n_1566;
wire n_717;
wire n_2006;
wire n_952;
wire n_864;
wire n_2446;
wire n_1096;
wire n_1379;
wire n_2436;
wire n_2376;
wire n_2367;
wire n_1706;
wire n_2207;
wire n_2461;
wire n_634;
wire n_1214;
wire n_1839;
wire n_1246;
wire n_1138;
wire n_2042;
wire n_2123;
wire n_1853;
wire n_764;
wire n_1503;
wire n_2238;
wire n_2529;
wire n_2374;
wire n_1196;
wire n_1181;
wire n_1999;
wire n_2380;
wire n_1187;
wire n_1131;
wire n_1225;
wire n_737;
wire n_1298;
wire n_1745;
wire n_1366;
wire n_2084;
wire n_568;
wire n_2278;
wire n_1088;
wire n_1424;
wire n_766;
wire n_1835;
wire n_1457;
wire n_2482;
wire n_1682;
wire n_1836;
wire n_870;
wire n_1453;
wire n_958;
wire n_945;
wire n_2248;
wire n_813;
wire n_1985;
wire n_2288;
wire n_995;
wire n_1909;
wire n_2156;
wire n_1184;
wire n_1961;
wire n_1535;
wire n_665;
wire n_754;
wire n_903;
wire n_871;
wire n_2323;
wire n_1073;
wire n_1979;
wire n_1277;
wire n_2107;
wire n_1746;
wire n_1761;
wire n_829;
wire n_1062;
wire n_738;
wire n_1690;
wire n_2221;
wire n_672;
wire n_740;
wire n_1283;
wire n_2317;
wire n_1974;
wire n_1736;
wire n_1018;
wire n_2342;
wire n_2200;
wire n_2442;
wire n_953;
wire n_1364;
wire n_2390;
wire n_1888;
wire n_1224;
wire n_2109;
wire n_1425;
wire n_625;
wire n_557;
wire n_2322;
wire n_1107;
wire n_1688;
wire n_989;
wire n_645;
wire n_1944;
wire n_559;
wire n_2233;
wire n_2370;
wire n_1988;
wire n_795;
wire n_721;
wire n_1084;
wire n_1718;
wire n_1276;
wire n_1936;
wire n_2149;
wire n_2277;
wire n_1428;
wire n_1284;
wire n_1241;
wire n_821;
wire n_561;
wire n_770;
wire n_1514;
wire n_1528;
wire n_901;
wire n_569;
wire n_2078;
wire n_1145;
wire n_971;
wire n_2359;
wire n_2201;
wire n_787;
wire n_1650;
wire n_1519;
wire n_1195;
wire n_2049;
wire n_1522;
wire n_1207;
wire n_786;
wire n_1404;
wire n_868;
wire n_2232;
wire n_1847;
wire n_2458;
wire n_1542;
wire n_1314;
wire n_1512;
wire n_2227;
wire n_2301;
wire n_1539;
wire n_884;
wire n_1851;
wire n_2162;
wire n_1415;
wire n_1034;
wire n_1652;
wire n_2192;
wire n_1676;
wire n_1085;
wire n_1636;
wire n_823;
wire n_1900;
wire n_620;
wire n_1074;
wire n_859;
wire n_1765;
wire n_1889;
wire n_587;
wire n_1977;
wire n_693;
wire n_863;
wire n_1254;
wire n_929;
wire n_2433;
wire n_1703;
wire n_899;
wire n_2332;
wire n_2391;
wire n_611;
wire n_1295;
wire n_2060;
wire n_1850;
wire n_2004;
wire n_1013;
wire n_1495;
wire n_1637;
wire n_2427;
wire n_661;
wire n_2098;
wire n_1751;
wire n_1917;
wire n_2456;
wire n_1924;
wire n_1560;
wire n_1654;
wire n_2341;
wire n_1548;
wire n_1811;
wire n_2045;
wire n_1396;
wire n_1230;
wire n_612;
wire n_1840;
wire n_1597;
wire n_1771;
wire n_1544;
wire n_579;
wire n_844;
wire n_1012;
wire n_1267;
wire n_2061;
wire n_2094;
wire n_2512;
wire n_1354;
wire n_1790;
wire n_1213;
wire n_2382;
wire n_2043;
wire n_780;
wire n_2349;
wire n_1918;
wire n_1021;
wire n_1443;
wire n_1465;
wire n_1949;
wire n_1595;
wire n_1142;
wire n_1140;
wire n_705;
wire n_570;
wire n_942;
wire n_1437;
wire n_2077;
wire n_1378;
wire n_1121;
wire n_1416;
wire n_1461;
wire n_1391;
wire n_1947;
wire n_1599;
wire n_1876;
wire n_1006;
wire n_1830;
wire n_575;
wire n_546;
wire n_2527;
wire n_1112;
wire n_1159;
wire n_700;
wire n_772;
wire n_1216;
wire n_1245;
wire n_1669;
wire n_1675;
wire n_2466;
wire n_676;
wire n_2038;
wire n_2263;
wire n_2116;
wire n_2271;
wire n_2145;
wire n_2326;
wire n_1838;
wire n_1594;
wire n_680;
wire n_1935;
wire n_1716;
wire n_1872;
wire n_1585;
wire n_2281;
wire n_1432;
wire n_2245;
wire n_1108;
wire n_851;
wire n_1590;
wire n_1351;
wire n_2216;
wire n_1274;
wire n_2426;
wire n_652;
wire n_1819;
wire n_947;
wire n_2134;
wire n_930;
wire n_1260;
wire n_1179;
wire n_696;
wire n_1442;
wire n_798;
wire n_577;
wire n_1833;
wire n_1691;
wire n_916;
wire n_1386;
wire n_912;
wire n_1884;
wire n_1555;
wire n_1842;
wire n_2499;
wire n_762;
wire n_1253;
wire n_1468;
wire n_1661;
wire n_555;
wire n_804;
wire n_1656;
wire n_1382;
wire n_992;
wire n_966;
wire n_955;
wire n_1182;
wire n_794;
wire n_2166;
wire n_1692;
wire n_1562;
wire n_2185;
wire n_2398;
wire n_1376;
wire n_1292;
wire n_1178;
wire n_2015;
wire n_1972;
wire n_1435;
wire n_1750;
wire n_1026;
wire n_1506;
wire n_1610;
wire n_2202;
wire n_2072;
wire n_2415;
wire n_2087;
wire n_931;
wire n_669;
wire n_1491;
wire n_619;
wire n_967;
wire n_1083;
wire n_2161;
wire n_1418;
wire n_746;
wire n_1357;
wire n_1079;
wire n_1787;
wire n_2462;
wire n_1389;
wire n_2155;
wire n_615;
wire n_1139;
wire n_2439;
wire n_1312;
wire n_1717;
wire n_1812;
wire n_824;
wire n_2172;
wire n_892;
wire n_1880;
wire n_959;
wire n_2365;
wire n_2257;
wire n_1399;
wire n_1101;
wire n_1567;
wire n_1343;
wire n_563;
wire n_2219;
wire n_1855;
wire n_2100;
wire n_2333;
wire n_990;
wire n_1623;
wire n_1903;
wire n_867;
wire n_2147;
wire n_2435;
wire n_1226;
wire n_2224;
wire n_944;
wire n_749;
wire n_1932;
wire n_1780;
wire n_1970;
wire n_1920;
wire n_2083;
wire n_815;
wire n_542;
wire n_2167;
wire n_2293;
wire n_1340;
wire n_1240;
wire n_1087;
wire n_2400;
wire n_632;
wire n_650;
wire n_2388;
wire n_2273;
wire n_1433;
wire n_1911;
wire n_1908;
wire n_1825;
wire n_1155;
wire n_1071;
wire n_976;
wire n_712;
wire n_909;
wire n_1392;
wire n_767;
wire n_1832;
wire n_1841;
wire n_1680;
wire n_2066;
wire n_2302;
wire n_964;
wire n_1627;
wire n_2220;
wire n_2294;
wire n_2274;
wire n_974;
wire n_1731;
wire n_799;
wire n_1147;
wire n_2378;
wire n_2467;
wire n_965;
wire n_1914;
wire n_2253;
wire n_934;
wire n_2213;
wire n_1447;
wire n_2363;
wire n_1220;
wire n_2019;
wire n_698;
wire n_2130;
wire n_1674;
wire n_2021;
wire n_2025;
wire n_2160;
wire n_1992;
wire n_1209;
wire n_1020;
wire n_1563;
wire n_646;
wire n_2507;
wire n_2142;
wire n_1633;
wire n_1913;
wire n_2069;
wire n_2495;
wire n_1058;
wire n_2328;
wire n_2434;
wire n_1042;
wire n_1234;
wire n_2311;
wire n_1578;
wire n_2261;
wire n_1455;
wire n_2287;
wire n_836;
wire n_2223;
wire n_1279;
wire n_2473;
wire n_2144;
wire n_2511;
wire n_564;
wire n_1029;
wire n_1247;
wire n_760;
wire n_2438;
wire n_1568;
wire n_1483;
wire n_1363;
wire n_1111;
wire n_970;
wire n_1689;
wire n_713;
wire n_1255;
wire n_1646;
wire n_598;
wire n_2262;
wire n_1237;
wire n_927;
wire n_1095;
wire n_1728;
wire n_2335;
wire n_706;
wire n_2120;
wire n_1401;
wire n_1419;
wire n_1531;
wire n_776;
wire n_2041;
wire n_2113;
wire n_1933;
wire n_1651;
wire n_1387;
wire n_1263;
wire n_1817;
wire n_2404;
wire n_2168;
wire n_552;
wire n_2312;
wire n_670;
wire n_1826;
wire n_2483;
wire n_1951;
wire n_2490;
wire n_1032;
wire n_1217;
wire n_1496;
wire n_637;
wire n_1592;
wire n_1259;
wire n_1177;
wire n_1231;
wire n_2132;
wire n_980;
wire n_1618;
wire n_1869;
wire n_1743;
wire n_905;
wire n_720;
wire n_926;
wire n_1943;
wire n_2296;
wire n_1802;
wire n_2178;
wire n_2112;
wire n_1163;
wire n_1795;
wire n_1384;
wire n_2237;
wire n_2146;
wire n_1868;
wire n_1501;
wire n_2241;
wire n_2373;
wire n_1173;
wire n_2350;
wire n_1068;
wire n_1198;
wire n_2531;
wire n_1570;
wire n_2099;
wire n_1518;
wire n_1456;
wire n_1879;
wire n_1886;
wire n_1648;
wire n_2187;
wire n_1413;
wire n_2481;
wire n_2129;
wire n_855;
wire n_2327;
wire n_808;
wire n_1365;
wire n_2476;
wire n_553;
wire n_2059;
wire n_2437;
wire n_1439;
wire n_814;
wire n_578;
wire n_2074;
wire n_1665;
wire n_1287;
wire n_1611;
wire n_2122;
wire n_2399;
wire n_1414;
wire n_1134;
wire n_2067;
wire n_1484;
wire n_1901;
wire n_647;
wire n_2055;
wire n_2027;
wire n_1423;
wire n_2117;
wire n_600;
wire n_1609;
wire n_1053;
wire n_1939;
wire n_2308;
wire n_2242;
wire n_1906;
wire n_1899;
wire n_2195;
wire n_2194;
wire n_1467;
wire n_1828;
wire n_2159;
wire n_1798;
wire n_1304;
wire n_1608;
wire n_1744;
wire n_2267;
wire n_1105;
wire n_547;
wire n_604;
wire n_677;
wire n_703;
wire n_1349;
wire n_1709;
wire n_1061;
wire n_2102;
wire n_681;
wire n_874;
wire n_2286;
wire n_2023;
wire n_1278;
wire n_707;
wire n_983;
wire n_590;
wire n_699;
wire n_727;
wire n_1726;
wire n_2075;
wire n_2523;
wire n_1945;
wire n_1015;
wire n_545;
wire n_2418;
wire n_1377;
wire n_1162;
wire n_1614;
wire n_2031;
wire n_2496;
wire n_2118;
wire n_1740;
wire n_1602;
wire n_688;
wire n_636;
wire n_1098;
wire n_1490;
wire n_2338;
wire n_777;
wire n_1553;
wire n_1080;
wire n_920;
wire n_1760;
wire n_1086;
wire n_1092;
wire n_2225;
wire n_986;
wire n_1104;
wire n_1963;
wire n_729;
wire n_887;
wire n_2057;
wire n_2218;
wire n_1122;
wire n_1205;
wire n_1408;
wire n_1693;
wire n_2125;
wire n_1132;
wire n_1156;
wire n_2184;
wire n_1823;
wire n_1120;
wire n_1202;
wire n_627;
wire n_2254;
wire n_1188;
wire n_1498;
wire n_1371;
wire n_2033;
wire n_957;
wire n_1402;
wire n_1242;
wire n_1607;
wire n_1489;
wire n_1218;
wire n_2217;
wire n_2226;
wire n_1586;
wire n_861;
wire n_1543;
wire n_1431;
wire n_877;
wire n_1119;
wire n_1863;
wire n_1763;
wire n_1666;
wire n_1500;
wire n_616;
wire n_2214;
wire n_1055;
wire n_1395;
wire n_1346;
wire n_2256;
wire n_1189;
wire n_1089;
wire n_1859;
wire n_1502;
wire n_1523;
wire n_2190;
wire n_1478;
wire n_1883;
wire n_2516;
wire n_1969;
wire n_735;
wire n_1005;
wire n_2379;
wire n_1294;
wire n_1667;
wire n_845;
wire n_888;
wire n_2300;
wire n_1649;
wire n_2452;
wire n_1677;
wire n_2470;
wire n_1927;
wire n_1297;
wire n_551;
wire n_1708;
wire n_1222;
wire n_2284;
wire n_1844;
wire n_2283;
wire n_582;
wire n_2526;
wire n_1957;
wire n_1953;
wire n_755;
wire n_1097;
wire n_1219;
wire n_1711;
wire n_710;
wire n_1919;
wire n_1791;
wire n_2508;
wire n_2124;
wire n_1894;
wire n_1460;
wire n_1239;
wire n_2266;
wire n_2449;
wire n_560;
wire n_890;
wire n_842;
wire n_1898;
wire n_745;
wire n_1741;
wire n_1572;
wire n_1907;
wire n_1793;
wire n_742;
wire n_1373;
wire n_1081;
wire n_1975;
wire n_1388;
wire n_1266;
wire n_1540;
wire n_1719;
wire n_2119;
wire n_769;
wire n_1797;
wire n_2366;
wire n_2493;
wire n_1753;
wire n_1990;
wire n_1372;
wire n_832;
wire n_744;
wire n_1895;
wire n_2474;
wire n_982;
wire n_1800;
wire n_915;
wire n_1075;
wire n_2008;
wire n_1331;
wire n_1890;
wire n_1529;
wire n_1227;
wire n_2127;
wire n_655;
wire n_1734;
wire n_1860;
wire n_2460;
wire n_1007;
wire n_1580;
wire n_1319;
wire n_657;
wire n_837;
wire n_812;
wire n_2448;
wire n_2211;
wire n_2292;
wire n_2480;
wire n_606;
wire n_951;
wire n_862;
wire n_1700;
wire n_659;
wire n_1332;
wire n_2306;
wire n_1854;
wire n_666;
wire n_1747;
wire n_2071;
wire n_2424;
wire n_1206;
wire n_1729;
wire n_722;
wire n_1508;
wire n_2414;
wire n_2082;
wire n_1532;
wire n_1171;
wire n_1030;
wire n_785;
wire n_2389;
wire n_1309;
wire n_999;
wire n_2280;
wire n_1766;
wire n_1338;
wire n_1342;
wire n_1867;
wire n_852;
wire n_1394;
wire n_704;
wire n_1060;
wire n_1044;
wire n_1714;
wire n_2140;
wire n_873;
wire n_1301;
wire n_1748;
wire n_2157;
wire n_1966;
wire n_1243;
wire n_2171;
wire n_2468;
wire n_1400;
wire n_2035;
wire n_1466;
wire n_1527;
wire n_1513;
wire n_1783;
wire n_608;
wire n_2494;
wire n_1538;
wire n_2457;
wire n_2128;
wire n_1037;
wire n_1329;
wire n_1993;
wire n_1545;
wire n_1257;
wire n_1480;
wire n_1954;
wire n_1668;
wire n_1878;
wire n_1605;
wire n_1078;
wire n_2486;
wire n_1897;
wire n_2520;
wire n_2137;
wire n_1161;
wire n_2489;
wire n_811;
wire n_624;
wire n_791;
wire n_876;
wire n_1191;
wire n_618;
wire n_2492;
wire n_736;
wire n_1025;
wire n_1215;
wire n_1449;
wire n_2337;
wire n_2265;
wire n_687;
wire n_797;
wire n_2026;
wire n_1786;
wire n_1327;
wire n_1475;
wire n_642;
wire n_1804;
wire n_2106;
wire n_1406;
wire n_595;
wire n_1405;
wire n_602;
wire n_2272;
wire n_1757;
wire n_592;
wire n_1499;
wire n_854;
wire n_1318;
wire n_2091;
wire n_1769;
wire n_1632;
wire n_1929;
wire n_1950;
wire n_2264;
wire n_805;
wire n_2032;
wire n_2090;
wire n_1658;
wire n_2249;
wire n_1072;
wire n_695;
wire n_1526;
wire n_1305;
wire n_730;
wire n_1596;
wire n_2348;
wire n_1281;
wire n_2364;
wire n_1997;
wire n_1137;
wire n_1873;
wire n_1258;
wire n_640;
wire n_1733;
wire n_1476;
wire n_1524;
wire n_1856;
wire n_2016;
wire n_943;
wire n_1118;
wire n_678;
wire n_651;
wire n_1874;
wire n_1293;
wire n_961;
wire n_1046;
wire n_1807;
wire n_1123;
wire n_726;
wire n_1657;
wire n_878;
wire n_1784;
wire n_771;
wire n_1321;
wire n_752;
wire n_2307;
wire n_1488;
wire n_985;
wire n_1330;
wire n_906;
wire n_1180;
wire n_1697;
wire n_2295;
wire n_806;
wire n_1984;
wire n_1350;
wire n_1556;
wire n_649;
wire n_1561;
wire n_2412;
wire n_1352;
wire n_2405;
wire n_1824;
wire n_643;
wire n_1492;
wire n_2383;
wire n_1441;
wire n_1822;
wire n_682;
wire n_1616;
wire n_2416;
wire n_819;
wire n_2386;
wire n_1971;
wire n_586;
wire n_1324;
wire n_1429;
wire n_2064;
wire n_2353;
wire n_2528;
wire n_1778;
wire n_1776;
wire n_686;
wire n_605;
wire n_1154;
wire n_584;
wire n_1557;
wire n_1759;
wire n_1829;
wire n_2325;
wire n_1130;
wire n_1450;
wire n_756;
wire n_2022;
wire n_1016;
wire n_2298;
wire n_1149;
wire n_1505;
wire n_2408;
wire n_2320;
wire n_979;
wire n_2329;
wire n_1642;
wire n_2417;
wire n_2525;
wire n_1815;
wire n_897;
wire n_949;
wire n_2454;
wire n_1493;
wire n_807;
wire n_891;
wire n_885;
wire n_1659;
wire n_2354;
wire n_1864;
wire n_1887;
wire n_1208;
wire n_1987;
wire n_2368;
wire n_802;
wire n_1151;
wire n_554;
wire n_960;
wire n_2352;
wire n_2502;
wire n_1256;
wire n_714;
wire n_2170;
wire n_790;
wire n_2244;
wire n_2143;
wire n_2393;
wire n_725;
wire n_2377;
wire n_1577;
wire n_1448;
wire n_2198;
wire n_1009;
wire n_1133;
wire n_883;
wire n_1852;
wire n_801;
wire n_1286;
wire n_818;
wire n_1685;
wire n_779;
wire n_2410;
wire n_2314;
wire n_2477;
wire n_2279;
wire n_594;
wire n_2222;
wire n_1995;
wire n_1877;
wire n_1397;
wire n_1052;
wire n_1333;
wire n_1306;
wire n_1849;
wire n_2076;
wire n_2133;
wire n_2203;
wire n_833;
wire n_1426;
wire n_2250;
wire n_2497;
wire n_2247;
wire n_2230;
wire n_879;
wire n_1117;
wire n_1269;
wire n_1303;
wire n_1547;
wire n_1438;
wire n_1541;
wire n_597;
wire n_2001;
wire n_1047;
wire n_2506;
wire n_1472;
wire n_2413;
wire n_1593;
wire n_1050;
wire n_566;
wire n_2158;
wire n_2285;
wire n_1288;
wire n_1201;
wire n_858;
wire n_1185;
wire n_2475;
wire n_2173;
wire n_1035;
wire n_1143;
wire n_2070;
wire n_2136;
wire n_1090;
wire n_2403;
wire n_1367;
wire n_2044;
wire n_928;
wire n_1153;
wire n_1103;
wire n_825;
wire n_732;
wire n_1565;
wire n_1192;
wire n_894;
wire n_1380;
wire n_1624;
wire n_1801;
wire n_1291;
wire n_562;
wire n_2020;
wire n_748;
wire n_2310;
wire n_1045;
wire n_1160;
wire n_1882;
wire n_1976;
wire n_1023;
wire n_1881;
wire n_988;
wire n_914;
wire n_689;
wire n_1116;
wire n_1958;
wire n_1511;
wire n_2177;
wire n_1422;
wire n_1965;
wire n_644;
wire n_1197;
wire n_1165;
wire n_1641;
wire n_538;
wire n_1517;
wire n_2036;
wire n_576;
wire n_843;
wire n_588;
wire n_638;
wire n_2003;
wire n_2210;
wire n_1307;
wire n_1128;
wire n_2053;
wire n_1671;
wire n_1417;
wire n_1048;
wire n_2343;
wire n_775;
wire n_667;
wire n_2419;
wire n_1049;
wire n_2330;
wire n_869;
wire n_846;
wire n_1398;
wire n_1921;
wire n_2450;
wire n_2411;
wire n_1356;
wire n_1341;
wire n_2234;
wire n_2309;
wire n_1504;
wire n_1955;
wire n_2110;
wire n_2431;
wire n_1773;
wire n_1440;
wire n_1370;
wire n_1603;
wire n_728;
wire n_2401;
wire n_715;
wire n_889;
wire n_1066;
wire n_1549;
wire n_2331;
wire n_935;
wire n_2478;
wire n_685;
wire n_911;
wire n_623;
wire n_1712;
wire n_1403;
wire n_1065;
wire n_1534;
wire n_1948;
wire n_810;
wire n_1290;
wire n_1959;
wire n_617;
wire n_2396;
wire n_543;
wire n_1362;
wire n_1559;
wire n_2121;
wire n_601;
wire n_683;
wire n_565;
wire n_628;
wire n_1300;
wire n_1960;
wire n_2068;
wire n_743;
wire n_1194;
wire n_1647;
wire n_1546;
wire n_1420;
wire n_907;
wire n_1454;
wire n_660;
wire n_2459;
wire n_962;
wire n_941;
wire n_1210;
wire n_847;
wire n_747;
wire n_1622;
wire n_1135;
wire n_918;
wire n_1968;
wire n_1885;
wire n_639;
wire n_673;
wire n_2196;
wire n_1038;
wire n_2371;
wire n_1978;
wire n_571;
wire n_1521;
wire n_1694;
wire n_1940;
wire n_593;
wire n_1695;
wire n_1164;
wire n_2313;
wire n_609;
wire n_1193;
wire n_1345;
wire n_613;
wire n_1022;
wire n_1336;
wire n_1033;
wire n_1774;
wire n_1166;
wire n_1056;
wire n_2007;
wire n_1994;
wire n_1767;
wire n_1040;
wire n_674;
wire n_1158;
wire n_1973;
wire n_1444;
wire n_1803;
wire n_820;
wire n_1749;
wire n_872;
wire n_1653;
wire n_2303;
wire n_1157;
wire n_1584;
wire n_848;
wire n_1664;
wire n_629;
wire n_1739;
wire n_1814;
wire n_2154;
wire n_2441;
wire n_2236;
wire n_1789;
wire n_763;
wire n_1986;
wire n_2174;
wire n_540;
wire n_692;
wire n_2054;
wire n_1857;
wire n_2315;
wire n_984;
wire n_1687;
wire n_2073;
wire n_2150;
wire n_1552;
wire n_750;
wire n_834;
wire n_1612;
wire n_2498;
wire n_800;
wire n_2046;
wire n_1816;
wire n_1910;
wire n_1756;
wire n_1606;
wire n_2189;
wire n_621;
wire n_1587;
wire n_2093;
wire n_2340;
wire n_2018;
wire n_1772;
wire n_2444;
wire n_1014;
wire n_724;
wire n_2204;
wire n_1427;
wire n_1481;
wire n_2040;
wire n_1311;
wire n_2199;
wire n_1956;
wire n_1589;
wire n_2151;
wire n_1100;
wire n_585;
wire n_875;
wire n_1617;
wire n_2455;
wire n_827;
wire n_2231;
wire n_697;
wire n_622;
wire n_1626;
wire n_1962;
wire n_1335;
wire n_1715;
wire n_2305;
wire n_880;
wire n_793;
wire n_2114;
wire n_1175;
wire n_2289;
wire n_2530;
wire n_2299;
wire n_751;
wire n_1027;
wire n_1070;
wire n_2406;
wire n_1621;
wire n_739;
wire n_1485;
wire n_1028;
wire n_1221;
wire n_1785;
wire n_792;
wire n_1262;
wire n_1942;
wire n_2180;
wire n_580;
wire n_1579;
wire n_2181;
wire n_2014;
wire n_975;
wire n_923;
wire n_1645;
wire n_1124;
wire n_1381;
wire n_1494;
wire n_932;
wire n_1893;
wire n_1183;
wire n_1326;
wire n_2276;
wire n_1805;
wire n_2282;
wire n_981;
wire n_2141;
wire n_1110;
wire n_1758;
wire n_2503;
wire n_2270;
wire n_2443;
wire n_1407;
wire n_2465;
wire n_1204;
wire n_1554;
wire n_994;
wire n_2428;
wire n_1360;
wire n_973;
wire n_972;
wire n_2251;
wire n_856;
wire n_1248;
wire n_1176;
wire n_1564;
wire n_2010;
wire n_1054;
wire n_1679;
wire n_2126;
wire n_1952;
wire n_2425;
wire n_2394;
wire n_1858;
wire n_1678;
wire n_1482;
wire n_1361;
wire n_2356;
wire n_1601;
wire n_1057;
wire n_2487;
wire n_1834;
wire n_1011;
wire n_978;
wire n_1520;
wire n_2488;
wire n_1509;
wire n_828;
wire n_1411;
wire n_1359;
wire n_558;
wire n_1721;
wire n_653;
wire n_1445;
wire n_1317;
wire n_2050;
wire n_2197;
wire n_783;
wire n_556;
wire n_1127;
wire n_1536;
wire n_1471;
wire n_2385;
wire n_2387;
wire n_1008;
wire n_581;
wire n_1024;
wire n_830;
wire n_2291;
wire n_1980;
wire n_2518;
wire n_987;
wire n_936;
wire n_2510;
wire n_1620;
wire n_2501;
wire n_1385;
wire n_1525;
wire n_1998;
wire n_2165;
wire n_541;
wire n_1775;
wire n_788;
wire n_908;
wire n_1036;
wire n_2169;
wire n_1270;
wire n_1167;
wire n_1272;
wire n_549;
wire n_591;
wire n_969;
wire n_2028;
wire n_919;
wire n_1663;
wire n_2092;
wire n_2175;
wire n_1625;
wire n_2086;
wire n_1926;
wire n_2402;
wire n_1458;
wire n_679;
wire n_1630;
wire n_663;
wire n_1720;
wire n_2409;
wire n_2176;
wire n_1412;
wire n_1738;
wire n_1550;
wire n_1358;
wire n_1200;
wire n_826;
wire n_2453;
wire n_2344;
wire n_1922;
wire n_1735;
wire n_1788;
wire n_940;
wire n_2392;
wire n_1537;
wire n_2138;
wire n_2065;
wire n_2321;
wire n_1077;
wire n_607;
wire n_956;
wire n_1930;
wire n_765;
wire n_1809;
wire n_1904;
wire n_1843;
wire n_2000;
wire n_1268;
wire n_2395;
wire n_917;
wire n_1271;
wire n_2096;
wire n_2440;
wire n_2186;
wire n_1530;
wire n_2215;
wire n_631;
wire n_1170;
wire n_2258;
wire n_1261;
wire n_2471;
wire n_702;
wire n_857;
wire n_898;
wire n_968;
wire n_1067;
wire n_1235;
wire n_1323;
wire n_2375;
wire n_1462;
wire n_1937;
wire n_2012;
wire n_1064;
wire n_633;
wire n_900;
wire n_1446;
wire n_1282;
wire n_1701;
wire n_1093;
wire n_1551;
wire n_2039;
wire n_1755;
wire n_1285;
wire n_733;
wire n_761;
wire n_2212;
wire n_731;
wire n_1813;
wire n_2268;
wire n_1452;
wire n_1573;
wire n_668;
wire n_758;
wire n_2252;
wire n_2111;
wire n_2420;
wire n_1996;
wire n_1106;
wire n_2009;
wire n_648;
wire n_784;
wire n_816;
wire n_1322;
wire n_1473;
wire n_835;
wire n_1076;
wire n_2024;
wire n_1348;
wire n_753;
wire n_2445;
wire n_1770;
wire n_701;
wire n_1003;
wire n_2469;
wire n_1125;
wire n_2103;
wire n_2358;
wire n_1710;
wire n_1865;
wire n_2522;
wire n_2463;
wire n_1344;
wire n_2355;
wire n_1390;
wire n_1792;
wire n_2062;
wire n_1141;
wire n_1629;
wire n_1640;
wire n_822;
wire n_1094;
wire n_840;
wire n_1459;
wire n_2153;
wire n_2324;
wire n_1510;
wire n_2505;
wire n_2139;
wire n_1099;
wire n_839;
wire n_1754;
wire n_759;
wire n_567;
wire n_2397;
wire n_2521;
wire n_1727;
wire n_2235;
wire n_1991;
wire n_1575;
wire n_1848;
wire n_1892;
wire n_1172;
wire n_614;
wire n_1212;
wire n_831;
wire n_778;
wire n_1619;
wire n_2351;
wire n_2260;
wire n_550;
wire n_1315;
wire n_1660;
wire n_1902;
wire n_997;
wire n_635;
wire n_2206;
wire n_694;
wire n_1643;
wire n_1320;
wire n_1113;
wire n_2347;
wire n_1152;
wire n_2447;
wire n_2034;
wire n_1845;
wire n_1934;
wire n_2101;
wire n_921;
wire n_2362;
wire n_1615;
wire n_1236;
wire n_2104;
wire n_1265;
wire n_1576;
wire n_2105;
wire n_1470;
wire n_671;
wire n_1533;
wire n_1806;
wire n_2372;
wire n_1409;
wire n_1148;
wire n_1588;
wire n_1684;
wire n_1673;
wire n_2422;
wire n_1334;
wire n_654;
wire n_2290;
wire n_2088;
wire n_1275;
wire n_904;
wire n_2005;
wire n_2048;
wire n_1696;
wire n_1875;
wire n_1059;
wire n_684;
wire n_2429;
wire n_2108;
wire n_1039;
wire n_2246;
wire n_539;
wire n_1150;
wire n_977;
wire n_2339;
wire n_1628;
wire n_1289;
wire n_1831;
wire n_2191;
wire n_1497;
wire n_1866;
wire n_2472;
wire n_2056;
wire n_1136;
wire n_2515;
wire n_1782;
wire n_1190;
wire n_1600;
wire n_1144;
wire n_838;
wire n_1558;
wire n_1941;
wire n_1316;
wire n_2519;
wire n_950;
wire n_1017;
wire n_711;
wire n_734;
wire n_1915;
wire n_2360;
wire n_723;
wire n_1393;
wire n_2240;
wire n_658;
wire n_630;
wire n_1369;
wire n_1781;
wire n_709;
wire n_809;
wire n_2085;
wire n_2432;
wire n_1686;
wire n_1964;
wire n_881;
wire n_1019;
wire n_1477;
wire n_1777;
wire n_2188;
wire n_1982;
wire n_2097;
wire n_662;
wire n_641;
wire n_2430;
wire n_2504;
wire n_910;
wire n_741;
wire n_939;
wire n_1410;
wire n_2297;
wire n_1114;
wire n_1325;
wire n_1742;
wire n_708;
wire n_1223;
wire n_1768;
wire n_2513;
wire n_2193;
wire n_2369;
wire n_572;
wire n_1199;
wire n_865;
wire n_1273;
wire n_1983;
wire n_1041;
wire n_2451;
wire n_2115;
wire n_993;
wire n_1862;
wire n_948;
wire n_2017;
wire n_922;
wire n_1004;
wire n_1810;
wire n_1347;
wire n_860;
wire n_1043;
wire n_1923;
wire n_1764;
wire n_896;
wire n_1737;
wire n_1479;
wire n_1613;
wire n_902;
wire n_1031;
wire n_1723;
wire n_1638;
wire n_853;
wire n_716;
wire n_1571;
wire n_1698;
wire n_1337;
wire n_774;
wire n_1946;
wire n_2148;
wire n_933;
wire n_1779;
wire n_596;
wire n_954;
wire n_2051;
wire n_1168;
wire n_1821;
wire n_1310;
wire n_656;
wire n_574;
wire n_664;
wire n_1591;
wire n_1229;
wire n_1683;
wire n_1896;
wire n_2164;
wire n_1732;
wire n_2381;
wire n_1967;
wire n_2384;
wire n_2179;
wire n_1280;
wire n_544;
wire n_1516;
wire n_1186;
wire n_1705;
wire n_599;
wire n_768;
wire n_1091;
wire n_2052;
wire n_2485;
wire n_537;
wire n_1063;
wire n_991;
wire n_2183;
wire n_2205;
wire n_2275;
wire n_1724;
wire n_1670;
wire n_1707;
wire n_1799;
wire n_2080;
wire n_2058;
wire n_1126;
wire n_2357;
wire n_2029;
wire n_1846;
wire n_1912;
wire n_938;
wire n_1891;
wire n_1328;
wire n_895;
wire n_1639;
wire n_583;
wire n_2209;
wire n_2421;
wire n_1302;
wire n_1000;
wire n_626;
wire n_1581;
wire n_1928;
wire n_946;
wire n_757;
wire n_2047;
wire n_1655;
wire n_1818;
wire n_1146;
wire n_1634;
wire n_1203;
wire n_998;
wire n_1699;
wire n_1598;
wire n_2269;
wire n_2081;
wire n_937;
wire n_1474;
wire n_2524;
wire n_1583;
wire n_1604;
wire n_1631;
wire n_1702;
wire n_1794;
wire n_1375;
wire n_1232;
wire n_996;
wire n_1211;
wire n_1368;
wire n_963;
wire n_1264;
wire n_1082;
wire n_1725;
wire n_2318;
wire n_1827;
wire n_866;
wire n_925;
wire n_1752;
wire n_1313;
wire n_1001;
wire n_1722;
wire n_2361;
wire n_1115;
wire n_2229;
wire n_1339;
wire n_1002;
wire n_1644;
wire n_1051;
wire n_719;
wire n_1102;
wire n_2255;
wire n_1129;
wire n_1252;
wire n_2239;
wire n_1464;
wire n_1296;
wire n_773;
wire n_2316;
wire n_2464;
wire n_1010;
wire n_882;
wire n_2304;
wire n_1249;
wire n_803;
wire n_1871;
wire n_2514;
wire n_718;
wire n_1434;
wire n_1905;
wire n_1569;
wire n_548;
wire n_2336;
wire n_1662;
wire n_1299;
wire n_1870;
wire n_2063;
wire n_1925;
wire n_782;
wire n_2491;
wire n_1861;
wire n_2079;
wire n_1228;
wire n_2319;
wire n_2152;
wire n_2517;
wire n_1931;
wire n_1244;
wire n_1796;
wire n_2259;
wire n_849;
wire n_2095;
wire n_1820;
wire n_1251;
wire n_1989;
wire n_1421;
wire n_2208;
wire n_2423;
wire n_1762;
wire n_1233;
wire n_1808;
wire n_1574;
wire n_1672;
wire n_2228;
wire n_1635;
wire n_1704;
wire n_893;
wire n_1582;
wire n_841;
wire n_2479;
wire n_886;
wire n_1069;
wire n_1981;
wire n_2037;
wire n_1308;
wire n_796;
wire n_573;
wire n_2345;
wire n_1730;
wire n_1374;
wire n_1451;
wire n_2089;
wire n_1487;
wire n_675;

CKINVDCx5p33_ASAP7_75t_R g537 ( 
.A(n_106),
.Y(n_537)
);

CKINVDCx5p33_ASAP7_75t_R g538 ( 
.A(n_241),
.Y(n_538)
);

CKINVDCx5p33_ASAP7_75t_R g539 ( 
.A(n_262),
.Y(n_539)
);

CKINVDCx5p33_ASAP7_75t_R g540 ( 
.A(n_450),
.Y(n_540)
);

CKINVDCx20_ASAP7_75t_R g541 ( 
.A(n_484),
.Y(n_541)
);

CKINVDCx5p33_ASAP7_75t_R g542 ( 
.A(n_519),
.Y(n_542)
);

INVx2_ASAP7_75t_L g543 ( 
.A(n_22),
.Y(n_543)
);

CKINVDCx5p33_ASAP7_75t_R g544 ( 
.A(n_356),
.Y(n_544)
);

CKINVDCx5p33_ASAP7_75t_R g545 ( 
.A(n_402),
.Y(n_545)
);

CKINVDCx5p33_ASAP7_75t_R g546 ( 
.A(n_490),
.Y(n_546)
);

INVx1_ASAP7_75t_L g547 ( 
.A(n_204),
.Y(n_547)
);

INVx1_ASAP7_75t_L g548 ( 
.A(n_181),
.Y(n_548)
);

CKINVDCx5p33_ASAP7_75t_R g549 ( 
.A(n_414),
.Y(n_549)
);

BUFx10_ASAP7_75t_L g550 ( 
.A(n_121),
.Y(n_550)
);

INVx1_ASAP7_75t_L g551 ( 
.A(n_99),
.Y(n_551)
);

CKINVDCx5p33_ASAP7_75t_R g552 ( 
.A(n_524),
.Y(n_552)
);

BUFx3_ASAP7_75t_L g553 ( 
.A(n_497),
.Y(n_553)
);

CKINVDCx5p33_ASAP7_75t_R g554 ( 
.A(n_494),
.Y(n_554)
);

INVx1_ASAP7_75t_L g555 ( 
.A(n_417),
.Y(n_555)
);

INVx1_ASAP7_75t_L g556 ( 
.A(n_91),
.Y(n_556)
);

INVx1_ASAP7_75t_L g557 ( 
.A(n_521),
.Y(n_557)
);

INVxp67_ASAP7_75t_L g558 ( 
.A(n_527),
.Y(n_558)
);

CKINVDCx5p33_ASAP7_75t_R g559 ( 
.A(n_266),
.Y(n_559)
);

CKINVDCx5p33_ASAP7_75t_R g560 ( 
.A(n_21),
.Y(n_560)
);

BUFx6f_ASAP7_75t_L g561 ( 
.A(n_510),
.Y(n_561)
);

INVx1_ASAP7_75t_L g562 ( 
.A(n_508),
.Y(n_562)
);

CKINVDCx5p33_ASAP7_75t_R g563 ( 
.A(n_514),
.Y(n_563)
);

CKINVDCx5p33_ASAP7_75t_R g564 ( 
.A(n_350),
.Y(n_564)
);

CKINVDCx16_ASAP7_75t_R g565 ( 
.A(n_433),
.Y(n_565)
);

CKINVDCx5p33_ASAP7_75t_R g566 ( 
.A(n_200),
.Y(n_566)
);

INVx1_ASAP7_75t_L g567 ( 
.A(n_137),
.Y(n_567)
);

INVx2_ASAP7_75t_L g568 ( 
.A(n_24),
.Y(n_568)
);

CKINVDCx5p33_ASAP7_75t_R g569 ( 
.A(n_75),
.Y(n_569)
);

CKINVDCx5p33_ASAP7_75t_R g570 ( 
.A(n_163),
.Y(n_570)
);

INVx1_ASAP7_75t_L g571 ( 
.A(n_218),
.Y(n_571)
);

INVx2_ASAP7_75t_L g572 ( 
.A(n_307),
.Y(n_572)
);

CKINVDCx5p33_ASAP7_75t_R g573 ( 
.A(n_486),
.Y(n_573)
);

CKINVDCx5p33_ASAP7_75t_R g574 ( 
.A(n_506),
.Y(n_574)
);

INVx1_ASAP7_75t_L g575 ( 
.A(n_438),
.Y(n_575)
);

CKINVDCx5p33_ASAP7_75t_R g576 ( 
.A(n_43),
.Y(n_576)
);

INVx1_ASAP7_75t_L g577 ( 
.A(n_134),
.Y(n_577)
);

CKINVDCx14_ASAP7_75t_R g578 ( 
.A(n_254),
.Y(n_578)
);

INVxp67_ASAP7_75t_SL g579 ( 
.A(n_53),
.Y(n_579)
);

CKINVDCx5p33_ASAP7_75t_R g580 ( 
.A(n_535),
.Y(n_580)
);

CKINVDCx5p33_ASAP7_75t_R g581 ( 
.A(n_395),
.Y(n_581)
);

CKINVDCx5p33_ASAP7_75t_R g582 ( 
.A(n_485),
.Y(n_582)
);

CKINVDCx20_ASAP7_75t_R g583 ( 
.A(n_220),
.Y(n_583)
);

CKINVDCx5p33_ASAP7_75t_R g584 ( 
.A(n_134),
.Y(n_584)
);

INVx1_ASAP7_75t_L g585 ( 
.A(n_456),
.Y(n_585)
);

CKINVDCx5p33_ASAP7_75t_R g586 ( 
.A(n_489),
.Y(n_586)
);

CKINVDCx5p33_ASAP7_75t_R g587 ( 
.A(n_169),
.Y(n_587)
);

CKINVDCx5p33_ASAP7_75t_R g588 ( 
.A(n_79),
.Y(n_588)
);

CKINVDCx5p33_ASAP7_75t_R g589 ( 
.A(n_58),
.Y(n_589)
);

INVx1_ASAP7_75t_L g590 ( 
.A(n_493),
.Y(n_590)
);

INVx1_ASAP7_75t_L g591 ( 
.A(n_491),
.Y(n_591)
);

CKINVDCx5p33_ASAP7_75t_R g592 ( 
.A(n_386),
.Y(n_592)
);

INVx1_ASAP7_75t_L g593 ( 
.A(n_502),
.Y(n_593)
);

BUFx8_ASAP7_75t_SL g594 ( 
.A(n_348),
.Y(n_594)
);

CKINVDCx5p33_ASAP7_75t_R g595 ( 
.A(n_220),
.Y(n_595)
);

INVx1_ASAP7_75t_L g596 ( 
.A(n_32),
.Y(n_596)
);

CKINVDCx5p33_ASAP7_75t_R g597 ( 
.A(n_511),
.Y(n_597)
);

BUFx10_ASAP7_75t_L g598 ( 
.A(n_530),
.Y(n_598)
);

CKINVDCx5p33_ASAP7_75t_R g599 ( 
.A(n_503),
.Y(n_599)
);

INVx1_ASAP7_75t_L g600 ( 
.A(n_487),
.Y(n_600)
);

BUFx6f_ASAP7_75t_L g601 ( 
.A(n_515),
.Y(n_601)
);

CKINVDCx5p33_ASAP7_75t_R g602 ( 
.A(n_516),
.Y(n_602)
);

INVx1_ASAP7_75t_L g603 ( 
.A(n_179),
.Y(n_603)
);

INVx1_ASAP7_75t_L g604 ( 
.A(n_498),
.Y(n_604)
);

CKINVDCx5p33_ASAP7_75t_R g605 ( 
.A(n_193),
.Y(n_605)
);

INVx1_ASAP7_75t_L g606 ( 
.A(n_407),
.Y(n_606)
);

INVx1_ASAP7_75t_L g607 ( 
.A(n_212),
.Y(n_607)
);

INVx2_ASAP7_75t_L g608 ( 
.A(n_449),
.Y(n_608)
);

CKINVDCx20_ASAP7_75t_R g609 ( 
.A(n_281),
.Y(n_609)
);

INVx1_ASAP7_75t_SL g610 ( 
.A(n_5),
.Y(n_610)
);

CKINVDCx5p33_ASAP7_75t_R g611 ( 
.A(n_49),
.Y(n_611)
);

CKINVDCx5p33_ASAP7_75t_R g612 ( 
.A(n_403),
.Y(n_612)
);

CKINVDCx5p33_ASAP7_75t_R g613 ( 
.A(n_146),
.Y(n_613)
);

CKINVDCx5p33_ASAP7_75t_R g614 ( 
.A(n_492),
.Y(n_614)
);

CKINVDCx5p33_ASAP7_75t_R g615 ( 
.A(n_522),
.Y(n_615)
);

CKINVDCx5p33_ASAP7_75t_R g616 ( 
.A(n_337),
.Y(n_616)
);

INVx1_ASAP7_75t_L g617 ( 
.A(n_353),
.Y(n_617)
);

CKINVDCx5p33_ASAP7_75t_R g618 ( 
.A(n_426),
.Y(n_618)
);

CKINVDCx5p33_ASAP7_75t_R g619 ( 
.A(n_251),
.Y(n_619)
);

CKINVDCx5p33_ASAP7_75t_R g620 ( 
.A(n_174),
.Y(n_620)
);

HB1xp67_ASAP7_75t_L g621 ( 
.A(n_488),
.Y(n_621)
);

INVx1_ASAP7_75t_L g622 ( 
.A(n_400),
.Y(n_622)
);

INVx1_ASAP7_75t_L g623 ( 
.A(n_461),
.Y(n_623)
);

CKINVDCx5p33_ASAP7_75t_R g624 ( 
.A(n_513),
.Y(n_624)
);

INVx1_ASAP7_75t_L g625 ( 
.A(n_120),
.Y(n_625)
);

CKINVDCx5p33_ASAP7_75t_R g626 ( 
.A(n_283),
.Y(n_626)
);

INVx1_ASAP7_75t_SL g627 ( 
.A(n_218),
.Y(n_627)
);

INVx2_ASAP7_75t_L g628 ( 
.A(n_219),
.Y(n_628)
);

INVx1_ASAP7_75t_L g629 ( 
.A(n_183),
.Y(n_629)
);

CKINVDCx5p33_ASAP7_75t_R g630 ( 
.A(n_451),
.Y(n_630)
);

CKINVDCx5p33_ASAP7_75t_R g631 ( 
.A(n_293),
.Y(n_631)
);

CKINVDCx5p33_ASAP7_75t_R g632 ( 
.A(n_428),
.Y(n_632)
);

CKINVDCx5p33_ASAP7_75t_R g633 ( 
.A(n_533),
.Y(n_633)
);

CKINVDCx5p33_ASAP7_75t_R g634 ( 
.A(n_57),
.Y(n_634)
);

INVx1_ASAP7_75t_L g635 ( 
.A(n_164),
.Y(n_635)
);

CKINVDCx5p33_ASAP7_75t_R g636 ( 
.A(n_4),
.Y(n_636)
);

CKINVDCx5p33_ASAP7_75t_R g637 ( 
.A(n_499),
.Y(n_637)
);

CKINVDCx20_ASAP7_75t_R g638 ( 
.A(n_318),
.Y(n_638)
);

BUFx8_ASAP7_75t_SL g639 ( 
.A(n_140),
.Y(n_639)
);

CKINVDCx5p33_ASAP7_75t_R g640 ( 
.A(n_64),
.Y(n_640)
);

CKINVDCx5p33_ASAP7_75t_R g641 ( 
.A(n_277),
.Y(n_641)
);

INVx1_ASAP7_75t_L g642 ( 
.A(n_313),
.Y(n_642)
);

INVx2_ASAP7_75t_L g643 ( 
.A(n_453),
.Y(n_643)
);

BUFx2_ASAP7_75t_R g644 ( 
.A(n_250),
.Y(n_644)
);

INVx1_ASAP7_75t_L g645 ( 
.A(n_430),
.Y(n_645)
);

CKINVDCx20_ASAP7_75t_R g646 ( 
.A(n_302),
.Y(n_646)
);

INVx1_ASAP7_75t_L g647 ( 
.A(n_207),
.Y(n_647)
);

INVx1_ASAP7_75t_L g648 ( 
.A(n_22),
.Y(n_648)
);

INVx1_ASAP7_75t_L g649 ( 
.A(n_8),
.Y(n_649)
);

INVx1_ASAP7_75t_L g650 ( 
.A(n_339),
.Y(n_650)
);

BUFx6f_ASAP7_75t_L g651 ( 
.A(n_365),
.Y(n_651)
);

CKINVDCx20_ASAP7_75t_R g652 ( 
.A(n_131),
.Y(n_652)
);

CKINVDCx5p33_ASAP7_75t_R g653 ( 
.A(n_387),
.Y(n_653)
);

CKINVDCx20_ASAP7_75t_R g654 ( 
.A(n_370),
.Y(n_654)
);

CKINVDCx5p33_ASAP7_75t_R g655 ( 
.A(n_518),
.Y(n_655)
);

BUFx2_ASAP7_75t_L g656 ( 
.A(n_14),
.Y(n_656)
);

CKINVDCx5p33_ASAP7_75t_R g657 ( 
.A(n_483),
.Y(n_657)
);

BUFx2_ASAP7_75t_L g658 ( 
.A(n_377),
.Y(n_658)
);

CKINVDCx5p33_ASAP7_75t_R g659 ( 
.A(n_7),
.Y(n_659)
);

INVx1_ASAP7_75t_L g660 ( 
.A(n_419),
.Y(n_660)
);

CKINVDCx14_ASAP7_75t_R g661 ( 
.A(n_211),
.Y(n_661)
);

CKINVDCx5p33_ASAP7_75t_R g662 ( 
.A(n_23),
.Y(n_662)
);

INVx1_ASAP7_75t_L g663 ( 
.A(n_394),
.Y(n_663)
);

CKINVDCx5p33_ASAP7_75t_R g664 ( 
.A(n_82),
.Y(n_664)
);

INVx1_ASAP7_75t_L g665 ( 
.A(n_409),
.Y(n_665)
);

INVx1_ASAP7_75t_L g666 ( 
.A(n_289),
.Y(n_666)
);

INVx1_ASAP7_75t_L g667 ( 
.A(n_175),
.Y(n_667)
);

CKINVDCx5p33_ASAP7_75t_R g668 ( 
.A(n_100),
.Y(n_668)
);

CKINVDCx5p33_ASAP7_75t_R g669 ( 
.A(n_139),
.Y(n_669)
);

CKINVDCx5p33_ASAP7_75t_R g670 ( 
.A(n_3),
.Y(n_670)
);

CKINVDCx20_ASAP7_75t_R g671 ( 
.A(n_505),
.Y(n_671)
);

INVx1_ASAP7_75t_L g672 ( 
.A(n_142),
.Y(n_672)
);

INVx1_ASAP7_75t_L g673 ( 
.A(n_5),
.Y(n_673)
);

CKINVDCx5p33_ASAP7_75t_R g674 ( 
.A(n_8),
.Y(n_674)
);

INVx1_ASAP7_75t_L g675 ( 
.A(n_235),
.Y(n_675)
);

CKINVDCx5p33_ASAP7_75t_R g676 ( 
.A(n_334),
.Y(n_676)
);

INVx1_ASAP7_75t_L g677 ( 
.A(n_473),
.Y(n_677)
);

CKINVDCx5p33_ASAP7_75t_R g678 ( 
.A(n_517),
.Y(n_678)
);

INVx1_ASAP7_75t_L g679 ( 
.A(n_101),
.Y(n_679)
);

INVx2_ASAP7_75t_L g680 ( 
.A(n_20),
.Y(n_680)
);

CKINVDCx5p33_ASAP7_75t_R g681 ( 
.A(n_341),
.Y(n_681)
);

BUFx10_ASAP7_75t_L g682 ( 
.A(n_531),
.Y(n_682)
);

CKINVDCx5p33_ASAP7_75t_R g683 ( 
.A(n_159),
.Y(n_683)
);

CKINVDCx5p33_ASAP7_75t_R g684 ( 
.A(n_297),
.Y(n_684)
);

INVx1_ASAP7_75t_L g685 ( 
.A(n_520),
.Y(n_685)
);

CKINVDCx5p33_ASAP7_75t_R g686 ( 
.A(n_131),
.Y(n_686)
);

INVx1_ASAP7_75t_L g687 ( 
.A(n_35),
.Y(n_687)
);

CKINVDCx5p33_ASAP7_75t_R g688 ( 
.A(n_374),
.Y(n_688)
);

INVx1_ASAP7_75t_L g689 ( 
.A(n_267),
.Y(n_689)
);

CKINVDCx5p33_ASAP7_75t_R g690 ( 
.A(n_238),
.Y(n_690)
);

BUFx2_ASAP7_75t_L g691 ( 
.A(n_232),
.Y(n_691)
);

CKINVDCx5p33_ASAP7_75t_R g692 ( 
.A(n_393),
.Y(n_692)
);

CKINVDCx5p33_ASAP7_75t_R g693 ( 
.A(n_279),
.Y(n_693)
);

CKINVDCx20_ASAP7_75t_R g694 ( 
.A(n_148),
.Y(n_694)
);

INVx1_ASAP7_75t_L g695 ( 
.A(n_270),
.Y(n_695)
);

CKINVDCx5p33_ASAP7_75t_R g696 ( 
.A(n_183),
.Y(n_696)
);

INVx1_ASAP7_75t_L g697 ( 
.A(n_340),
.Y(n_697)
);

CKINVDCx5p33_ASAP7_75t_R g698 ( 
.A(n_269),
.Y(n_698)
);

INVx1_ASAP7_75t_L g699 ( 
.A(n_421),
.Y(n_699)
);

INVx1_ASAP7_75t_L g700 ( 
.A(n_306),
.Y(n_700)
);

INVx1_ASAP7_75t_L g701 ( 
.A(n_225),
.Y(n_701)
);

INVx1_ASAP7_75t_L g702 ( 
.A(n_507),
.Y(n_702)
);

CKINVDCx5p33_ASAP7_75t_R g703 ( 
.A(n_106),
.Y(n_703)
);

CKINVDCx5p33_ASAP7_75t_R g704 ( 
.A(n_107),
.Y(n_704)
);

INVx1_ASAP7_75t_L g705 ( 
.A(n_178),
.Y(n_705)
);

CKINVDCx5p33_ASAP7_75t_R g706 ( 
.A(n_193),
.Y(n_706)
);

INVx2_ASAP7_75t_L g707 ( 
.A(n_75),
.Y(n_707)
);

CKINVDCx5p33_ASAP7_75t_R g708 ( 
.A(n_185),
.Y(n_708)
);

BUFx6f_ASAP7_75t_L g709 ( 
.A(n_0),
.Y(n_709)
);

INVx2_ASAP7_75t_L g710 ( 
.A(n_496),
.Y(n_710)
);

CKINVDCx5p33_ASAP7_75t_R g711 ( 
.A(n_63),
.Y(n_711)
);

CKINVDCx5p33_ASAP7_75t_R g712 ( 
.A(n_87),
.Y(n_712)
);

INVx1_ASAP7_75t_L g713 ( 
.A(n_276),
.Y(n_713)
);

CKINVDCx5p33_ASAP7_75t_R g714 ( 
.A(n_452),
.Y(n_714)
);

CKINVDCx5p33_ASAP7_75t_R g715 ( 
.A(n_432),
.Y(n_715)
);

CKINVDCx5p33_ASAP7_75t_R g716 ( 
.A(n_431),
.Y(n_716)
);

CKINVDCx20_ASAP7_75t_R g717 ( 
.A(n_125),
.Y(n_717)
);

CKINVDCx5p33_ASAP7_75t_R g718 ( 
.A(n_398),
.Y(n_718)
);

INVx2_ASAP7_75t_SL g719 ( 
.A(n_230),
.Y(n_719)
);

INVx1_ASAP7_75t_SL g720 ( 
.A(n_424),
.Y(n_720)
);

BUFx3_ASAP7_75t_L g721 ( 
.A(n_308),
.Y(n_721)
);

INVx2_ASAP7_75t_L g722 ( 
.A(n_207),
.Y(n_722)
);

INVx1_ASAP7_75t_L g723 ( 
.A(n_240),
.Y(n_723)
);

BUFx6f_ASAP7_75t_L g724 ( 
.A(n_444),
.Y(n_724)
);

CKINVDCx5p33_ASAP7_75t_R g725 ( 
.A(n_102),
.Y(n_725)
);

INVx1_ASAP7_75t_L g726 ( 
.A(n_310),
.Y(n_726)
);

INVx1_ASAP7_75t_L g727 ( 
.A(n_525),
.Y(n_727)
);

CKINVDCx5p33_ASAP7_75t_R g728 ( 
.A(n_80),
.Y(n_728)
);

INVx1_ASAP7_75t_L g729 ( 
.A(n_279),
.Y(n_729)
);

CKINVDCx5p33_ASAP7_75t_R g730 ( 
.A(n_495),
.Y(n_730)
);

INVx1_ASAP7_75t_L g731 ( 
.A(n_6),
.Y(n_731)
);

CKINVDCx5p33_ASAP7_75t_R g732 ( 
.A(n_126),
.Y(n_732)
);

INVx1_ASAP7_75t_L g733 ( 
.A(n_509),
.Y(n_733)
);

INVx1_ASAP7_75t_L g734 ( 
.A(n_504),
.Y(n_734)
);

CKINVDCx5p33_ASAP7_75t_R g735 ( 
.A(n_181),
.Y(n_735)
);

INVx2_ASAP7_75t_L g736 ( 
.A(n_221),
.Y(n_736)
);

BUFx5_ASAP7_75t_L g737 ( 
.A(n_39),
.Y(n_737)
);

INVx1_ASAP7_75t_SL g738 ( 
.A(n_465),
.Y(n_738)
);

CKINVDCx5p33_ASAP7_75t_R g739 ( 
.A(n_165),
.Y(n_739)
);

CKINVDCx5p33_ASAP7_75t_R g740 ( 
.A(n_122),
.Y(n_740)
);

INVx1_ASAP7_75t_SL g741 ( 
.A(n_298),
.Y(n_741)
);

CKINVDCx5p33_ASAP7_75t_R g742 ( 
.A(n_99),
.Y(n_742)
);

CKINVDCx5p33_ASAP7_75t_R g743 ( 
.A(n_252),
.Y(n_743)
);

INVx1_ASAP7_75t_L g744 ( 
.A(n_89),
.Y(n_744)
);

CKINVDCx5p33_ASAP7_75t_R g745 ( 
.A(n_174),
.Y(n_745)
);

CKINVDCx5p33_ASAP7_75t_R g746 ( 
.A(n_512),
.Y(n_746)
);

CKINVDCx5p33_ASAP7_75t_R g747 ( 
.A(n_501),
.Y(n_747)
);

INVx1_ASAP7_75t_L g748 ( 
.A(n_454),
.Y(n_748)
);

CKINVDCx5p33_ASAP7_75t_R g749 ( 
.A(n_40),
.Y(n_749)
);

CKINVDCx5p33_ASAP7_75t_R g750 ( 
.A(n_154),
.Y(n_750)
);

CKINVDCx5p33_ASAP7_75t_R g751 ( 
.A(n_371),
.Y(n_751)
);

CKINVDCx5p33_ASAP7_75t_R g752 ( 
.A(n_269),
.Y(n_752)
);

CKINVDCx5p33_ASAP7_75t_R g753 ( 
.A(n_94),
.Y(n_753)
);

CKINVDCx5p33_ASAP7_75t_R g754 ( 
.A(n_355),
.Y(n_754)
);

CKINVDCx5p33_ASAP7_75t_R g755 ( 
.A(n_500),
.Y(n_755)
);

CKINVDCx5p33_ASAP7_75t_R g756 ( 
.A(n_85),
.Y(n_756)
);

CKINVDCx20_ASAP7_75t_R g757 ( 
.A(n_467),
.Y(n_757)
);

BUFx3_ASAP7_75t_L g758 ( 
.A(n_529),
.Y(n_758)
);

CKINVDCx5p33_ASAP7_75t_R g759 ( 
.A(n_242),
.Y(n_759)
);

INVx1_ASAP7_75t_L g760 ( 
.A(n_329),
.Y(n_760)
);

CKINVDCx5p33_ASAP7_75t_R g761 ( 
.A(n_523),
.Y(n_761)
);

INVx1_ASAP7_75t_L g762 ( 
.A(n_165),
.Y(n_762)
);

INVx1_ASAP7_75t_SL g763 ( 
.A(n_469),
.Y(n_763)
);

HB1xp67_ASAP7_75t_L g764 ( 
.A(n_243),
.Y(n_764)
);

INVx1_ASAP7_75t_L g765 ( 
.A(n_20),
.Y(n_765)
);

INVx1_ASAP7_75t_L g766 ( 
.A(n_149),
.Y(n_766)
);

INVx1_ASAP7_75t_L g767 ( 
.A(n_180),
.Y(n_767)
);

CKINVDCx5p33_ASAP7_75t_R g768 ( 
.A(n_578),
.Y(n_768)
);

INVx1_ASAP7_75t_L g769 ( 
.A(n_737),
.Y(n_769)
);

INVx1_ASAP7_75t_L g770 ( 
.A(n_737),
.Y(n_770)
);

INVxp33_ASAP7_75t_L g771 ( 
.A(n_764),
.Y(n_771)
);

CKINVDCx20_ASAP7_75t_R g772 ( 
.A(n_609),
.Y(n_772)
);

INVx1_ASAP7_75t_L g773 ( 
.A(n_737),
.Y(n_773)
);

INVx1_ASAP7_75t_L g774 ( 
.A(n_737),
.Y(n_774)
);

INVx1_ASAP7_75t_L g775 ( 
.A(n_737),
.Y(n_775)
);

INVx1_ASAP7_75t_L g776 ( 
.A(n_737),
.Y(n_776)
);

INVx1_ASAP7_75t_L g777 ( 
.A(n_737),
.Y(n_777)
);

INVx2_ASAP7_75t_L g778 ( 
.A(n_709),
.Y(n_778)
);

INVx1_ASAP7_75t_L g779 ( 
.A(n_547),
.Y(n_779)
);

INVx1_ASAP7_75t_L g780 ( 
.A(n_548),
.Y(n_780)
);

INVx1_ASAP7_75t_L g781 ( 
.A(n_551),
.Y(n_781)
);

INVx1_ASAP7_75t_SL g782 ( 
.A(n_639),
.Y(n_782)
);

INVx1_ASAP7_75t_L g783 ( 
.A(n_556),
.Y(n_783)
);

INVx1_ASAP7_75t_L g784 ( 
.A(n_567),
.Y(n_784)
);

CKINVDCx14_ASAP7_75t_R g785 ( 
.A(n_578),
.Y(n_785)
);

INVx1_ASAP7_75t_L g786 ( 
.A(n_571),
.Y(n_786)
);

INVx1_ASAP7_75t_L g787 ( 
.A(n_577),
.Y(n_787)
);

INVxp33_ASAP7_75t_SL g788 ( 
.A(n_621),
.Y(n_788)
);

INVx1_ASAP7_75t_L g789 ( 
.A(n_596),
.Y(n_789)
);

INVx1_ASAP7_75t_L g790 ( 
.A(n_603),
.Y(n_790)
);

CKINVDCx5p33_ASAP7_75t_R g791 ( 
.A(n_661),
.Y(n_791)
);

INVxp33_ASAP7_75t_SL g792 ( 
.A(n_656),
.Y(n_792)
);

INVx1_ASAP7_75t_L g793 ( 
.A(n_607),
.Y(n_793)
);

INVxp67_ASAP7_75t_SL g794 ( 
.A(n_709),
.Y(n_794)
);

INVx1_ASAP7_75t_L g795 ( 
.A(n_625),
.Y(n_795)
);

INVx1_ASAP7_75t_L g796 ( 
.A(n_629),
.Y(n_796)
);

INVx1_ASAP7_75t_L g797 ( 
.A(n_635),
.Y(n_797)
);

INVx1_ASAP7_75t_L g798 ( 
.A(n_647),
.Y(n_798)
);

INVx1_ASAP7_75t_L g799 ( 
.A(n_648),
.Y(n_799)
);

INVxp67_ASAP7_75t_SL g800 ( 
.A(n_709),
.Y(n_800)
);

CKINVDCx5p33_ASAP7_75t_R g801 ( 
.A(n_661),
.Y(n_801)
);

CKINVDCx5p33_ASAP7_75t_R g802 ( 
.A(n_639),
.Y(n_802)
);

INVxp33_ASAP7_75t_SL g803 ( 
.A(n_691),
.Y(n_803)
);

INVx1_ASAP7_75t_L g804 ( 
.A(n_649),
.Y(n_804)
);

INVx1_ASAP7_75t_L g805 ( 
.A(n_666),
.Y(n_805)
);

INVx1_ASAP7_75t_L g806 ( 
.A(n_667),
.Y(n_806)
);

INVx1_ASAP7_75t_L g807 ( 
.A(n_672),
.Y(n_807)
);

INVx1_ASAP7_75t_L g808 ( 
.A(n_673),
.Y(n_808)
);

CKINVDCx5p33_ASAP7_75t_R g809 ( 
.A(n_565),
.Y(n_809)
);

INVx1_ASAP7_75t_L g810 ( 
.A(n_675),
.Y(n_810)
);

HB1xp67_ASAP7_75t_L g811 ( 
.A(n_537),
.Y(n_811)
);

INVx1_ASAP7_75t_L g812 ( 
.A(n_679),
.Y(n_812)
);

CKINVDCx5p33_ASAP7_75t_R g813 ( 
.A(n_594),
.Y(n_813)
);

CKINVDCx20_ASAP7_75t_R g814 ( 
.A(n_609),
.Y(n_814)
);

INVx1_ASAP7_75t_L g815 ( 
.A(n_687),
.Y(n_815)
);

INVx1_ASAP7_75t_L g816 ( 
.A(n_689),
.Y(n_816)
);

INVx1_ASAP7_75t_L g817 ( 
.A(n_695),
.Y(n_817)
);

INVx1_ASAP7_75t_L g818 ( 
.A(n_701),
.Y(n_818)
);

INVxp67_ASAP7_75t_L g819 ( 
.A(n_719),
.Y(n_819)
);

CKINVDCx5p33_ASAP7_75t_R g820 ( 
.A(n_594),
.Y(n_820)
);

INVx1_ASAP7_75t_L g821 ( 
.A(n_705),
.Y(n_821)
);

INVxp67_ASAP7_75t_SL g822 ( 
.A(n_709),
.Y(n_822)
);

CKINVDCx16_ASAP7_75t_R g823 ( 
.A(n_550),
.Y(n_823)
);

INVxp67_ASAP7_75t_SL g824 ( 
.A(n_543),
.Y(n_824)
);

INVx1_ASAP7_75t_L g825 ( 
.A(n_713),
.Y(n_825)
);

INVx1_ASAP7_75t_L g826 ( 
.A(n_723),
.Y(n_826)
);

INVx1_ASAP7_75t_L g827 ( 
.A(n_729),
.Y(n_827)
);

INVx1_ASAP7_75t_L g828 ( 
.A(n_731),
.Y(n_828)
);

INVx1_ASAP7_75t_L g829 ( 
.A(n_744),
.Y(n_829)
);

CKINVDCx5p33_ASAP7_75t_R g830 ( 
.A(n_658),
.Y(n_830)
);

INVx1_ASAP7_75t_L g831 ( 
.A(n_762),
.Y(n_831)
);

INVx1_ASAP7_75t_L g832 ( 
.A(n_765),
.Y(n_832)
);

INVx1_ASAP7_75t_L g833 ( 
.A(n_766),
.Y(n_833)
);

INVx1_ASAP7_75t_L g834 ( 
.A(n_767),
.Y(n_834)
);

INVx1_ASAP7_75t_L g835 ( 
.A(n_543),
.Y(n_835)
);

INVx1_ASAP7_75t_L g836 ( 
.A(n_568),
.Y(n_836)
);

INVx2_ASAP7_75t_SL g837 ( 
.A(n_550),
.Y(n_837)
);

CKINVDCx16_ASAP7_75t_R g838 ( 
.A(n_550),
.Y(n_838)
);

INVx1_ASAP7_75t_L g839 ( 
.A(n_568),
.Y(n_839)
);

CKINVDCx5p33_ASAP7_75t_R g840 ( 
.A(n_541),
.Y(n_840)
);

INVx1_ASAP7_75t_L g841 ( 
.A(n_628),
.Y(n_841)
);

INVx1_ASAP7_75t_SL g842 ( 
.A(n_644),
.Y(n_842)
);

INVxp67_ASAP7_75t_SL g843 ( 
.A(n_628),
.Y(n_843)
);

INVx1_ASAP7_75t_L g844 ( 
.A(n_680),
.Y(n_844)
);

INVx1_ASAP7_75t_L g845 ( 
.A(n_680),
.Y(n_845)
);

INVx1_ASAP7_75t_L g846 ( 
.A(n_707),
.Y(n_846)
);

INVx1_ASAP7_75t_L g847 ( 
.A(n_707),
.Y(n_847)
);

INVx1_ASAP7_75t_L g848 ( 
.A(n_722),
.Y(n_848)
);

INVx1_ASAP7_75t_L g849 ( 
.A(n_722),
.Y(n_849)
);

INVx1_ASAP7_75t_L g850 ( 
.A(n_736),
.Y(n_850)
);

BUFx2_ASAP7_75t_L g851 ( 
.A(n_736),
.Y(n_851)
);

INVx1_ASAP7_75t_L g852 ( 
.A(n_598),
.Y(n_852)
);

INVx1_ASAP7_75t_L g853 ( 
.A(n_598),
.Y(n_853)
);

INVx1_ASAP7_75t_L g854 ( 
.A(n_598),
.Y(n_854)
);

INVxp67_ASAP7_75t_SL g855 ( 
.A(n_553),
.Y(n_855)
);

INVxp33_ASAP7_75t_L g856 ( 
.A(n_572),
.Y(n_856)
);

CKINVDCx20_ASAP7_75t_R g857 ( 
.A(n_652),
.Y(n_857)
);

INVxp33_ASAP7_75t_SL g858 ( 
.A(n_538),
.Y(n_858)
);

INVx1_ASAP7_75t_L g859 ( 
.A(n_682),
.Y(n_859)
);

INVx1_ASAP7_75t_L g860 ( 
.A(n_682),
.Y(n_860)
);

INVx2_ASAP7_75t_L g861 ( 
.A(n_553),
.Y(n_861)
);

INVx1_ASAP7_75t_L g862 ( 
.A(n_682),
.Y(n_862)
);

CKINVDCx5p33_ASAP7_75t_R g863 ( 
.A(n_541),
.Y(n_863)
);

INVxp67_ASAP7_75t_SL g864 ( 
.A(n_721),
.Y(n_864)
);

INVx1_ASAP7_75t_L g865 ( 
.A(n_579),
.Y(n_865)
);

INVx1_ASAP7_75t_L g866 ( 
.A(n_555),
.Y(n_866)
);

INVx1_ASAP7_75t_L g867 ( 
.A(n_557),
.Y(n_867)
);

INVx1_ASAP7_75t_L g868 ( 
.A(n_562),
.Y(n_868)
);

BUFx6f_ASAP7_75t_L g869 ( 
.A(n_778),
.Y(n_869)
);

INVx1_ASAP7_75t_L g870 ( 
.A(n_769),
.Y(n_870)
);

INVx2_ASAP7_75t_L g871 ( 
.A(n_778),
.Y(n_871)
);

BUFx6f_ASAP7_75t_L g872 ( 
.A(n_770),
.Y(n_872)
);

INVx2_ASAP7_75t_L g873 ( 
.A(n_773),
.Y(n_873)
);

BUFx6f_ASAP7_75t_L g874 ( 
.A(n_774),
.Y(n_874)
);

INVx1_ASAP7_75t_L g875 ( 
.A(n_775),
.Y(n_875)
);

INVx2_ASAP7_75t_L g876 ( 
.A(n_776),
.Y(n_876)
);

AND2x2_ASAP7_75t_L g877 ( 
.A(n_785),
.B(n_721),
.Y(n_877)
);

INVx2_ASAP7_75t_L g878 ( 
.A(n_777),
.Y(n_878)
);

INVxp67_ASAP7_75t_L g879 ( 
.A(n_811),
.Y(n_879)
);

OA21x2_ASAP7_75t_L g880 ( 
.A1(n_866),
.A2(n_585),
.B(n_575),
.Y(n_880)
);

BUFx6f_ASAP7_75t_L g881 ( 
.A(n_861),
.Y(n_881)
);

AOI22x1_ASAP7_75t_SL g882 ( 
.A1(n_772),
.A2(n_652),
.B1(n_717),
.B2(n_694),
.Y(n_882)
);

OAI21x1_ASAP7_75t_L g883 ( 
.A1(n_867),
.A2(n_591),
.B(n_590),
.Y(n_883)
);

INVx3_ASAP7_75t_L g884 ( 
.A(n_861),
.Y(n_884)
);

NOR2xp33_ASAP7_75t_L g885 ( 
.A(n_788),
.B(n_558),
.Y(n_885)
);

AND2x4_ASAP7_75t_SL g886 ( 
.A(n_852),
.B(n_638),
.Y(n_886)
);

INVx1_ASAP7_75t_L g887 ( 
.A(n_794),
.Y(n_887)
);

INVx4_ASAP7_75t_L g888 ( 
.A(n_868),
.Y(n_888)
);

AND2x4_ASAP7_75t_L g889 ( 
.A(n_855),
.B(n_864),
.Y(n_889)
);

AND2x4_ASAP7_75t_L g890 ( 
.A(n_800),
.B(n_758),
.Y(n_890)
);

BUFx6f_ASAP7_75t_L g891 ( 
.A(n_835),
.Y(n_891)
);

BUFx2_ASAP7_75t_L g892 ( 
.A(n_813),
.Y(n_892)
);

INVx4_ASAP7_75t_L g893 ( 
.A(n_768),
.Y(n_893)
);

INVx2_ASAP7_75t_L g894 ( 
.A(n_836),
.Y(n_894)
);

INVx2_ASAP7_75t_SL g895 ( 
.A(n_768),
.Y(n_895)
);

INVx1_ASAP7_75t_L g896 ( 
.A(n_822),
.Y(n_896)
);

INVx2_ASAP7_75t_L g897 ( 
.A(n_839),
.Y(n_897)
);

INVx1_ASAP7_75t_L g898 ( 
.A(n_841),
.Y(n_898)
);

AND2x4_ASAP7_75t_L g899 ( 
.A(n_853),
.B(n_758),
.Y(n_899)
);

AND2x4_ASAP7_75t_L g900 ( 
.A(n_854),
.B(n_572),
.Y(n_900)
);

NOR2xp33_ASAP7_75t_L g901 ( 
.A(n_788),
.B(n_600),
.Y(n_901)
);

HB1xp67_ASAP7_75t_L g902 ( 
.A(n_782),
.Y(n_902)
);

OAI22x1_ASAP7_75t_R g903 ( 
.A1(n_772),
.A2(n_694),
.B1(n_717),
.B2(n_583),
.Y(n_903)
);

AND2x2_ASAP7_75t_L g904 ( 
.A(n_785),
.B(n_856),
.Y(n_904)
);

INVx3_ASAP7_75t_L g905 ( 
.A(n_844),
.Y(n_905)
);

AND2x4_ASAP7_75t_L g906 ( 
.A(n_859),
.B(n_860),
.Y(n_906)
);

INVx2_ASAP7_75t_L g907 ( 
.A(n_845),
.Y(n_907)
);

INVx2_ASAP7_75t_L g908 ( 
.A(n_846),
.Y(n_908)
);

NOR2xp33_ASAP7_75t_L g909 ( 
.A(n_862),
.B(n_593),
.Y(n_909)
);

BUFx3_ASAP7_75t_L g910 ( 
.A(n_779),
.Y(n_910)
);

INVx3_ASAP7_75t_L g911 ( 
.A(n_847),
.Y(n_911)
);

BUFx6f_ASAP7_75t_L g912 ( 
.A(n_848),
.Y(n_912)
);

BUFx12f_ASAP7_75t_L g913 ( 
.A(n_813),
.Y(n_913)
);

BUFx6f_ASAP7_75t_L g914 ( 
.A(n_849),
.Y(n_914)
);

INVx2_ASAP7_75t_L g915 ( 
.A(n_850),
.Y(n_915)
);

NAND2xp5_ASAP7_75t_L g916 ( 
.A(n_856),
.B(n_604),
.Y(n_916)
);

HB1xp67_ASAP7_75t_L g917 ( 
.A(n_802),
.Y(n_917)
);

HB1xp67_ASAP7_75t_L g918 ( 
.A(n_802),
.Y(n_918)
);

AND2x4_ASAP7_75t_L g919 ( 
.A(n_824),
.B(n_608),
.Y(n_919)
);

INVx4_ASAP7_75t_L g920 ( 
.A(n_791),
.Y(n_920)
);

INVx2_ASAP7_75t_L g921 ( 
.A(n_780),
.Y(n_921)
);

INVx2_ASAP7_75t_L g922 ( 
.A(n_781),
.Y(n_922)
);

OAI22x1_ASAP7_75t_SL g923 ( 
.A1(n_814),
.A2(n_610),
.B1(n_627),
.B2(n_749),
.Y(n_923)
);

INVx2_ASAP7_75t_L g924 ( 
.A(n_783),
.Y(n_924)
);

INVx2_ASAP7_75t_L g925 ( 
.A(n_784),
.Y(n_925)
);

NOR2xp33_ASAP7_75t_L g926 ( 
.A(n_791),
.B(n_606),
.Y(n_926)
);

INVx1_ASAP7_75t_L g927 ( 
.A(n_786),
.Y(n_927)
);

INVx1_ASAP7_75t_L g928 ( 
.A(n_787),
.Y(n_928)
);

INVx5_ASAP7_75t_L g929 ( 
.A(n_851),
.Y(n_929)
);

BUFx6f_ASAP7_75t_L g930 ( 
.A(n_789),
.Y(n_930)
);

INVx1_ASAP7_75t_L g931 ( 
.A(n_790),
.Y(n_931)
);

HB1xp67_ASAP7_75t_L g932 ( 
.A(n_820),
.Y(n_932)
);

AND2x4_ASAP7_75t_L g933 ( 
.A(n_843),
.B(n_608),
.Y(n_933)
);

INVx1_ASAP7_75t_L g934 ( 
.A(n_921),
.Y(n_934)
);

BUFx6f_ASAP7_75t_L g935 ( 
.A(n_881),
.Y(n_935)
);

BUFx6f_ASAP7_75t_L g936 ( 
.A(n_881),
.Y(n_936)
);

BUFx3_ASAP7_75t_L g937 ( 
.A(n_887),
.Y(n_937)
);

CKINVDCx5p33_ASAP7_75t_R g938 ( 
.A(n_913),
.Y(n_938)
);

INVx1_ASAP7_75t_L g939 ( 
.A(n_921),
.Y(n_939)
);

INVx2_ASAP7_75t_L g940 ( 
.A(n_873),
.Y(n_940)
);

CKINVDCx5p33_ASAP7_75t_R g941 ( 
.A(n_913),
.Y(n_941)
);

CKINVDCx20_ASAP7_75t_R g942 ( 
.A(n_903),
.Y(n_942)
);

CKINVDCx5p33_ASAP7_75t_R g943 ( 
.A(n_892),
.Y(n_943)
);

BUFx6f_ASAP7_75t_L g944 ( 
.A(n_881),
.Y(n_944)
);

INVx3_ASAP7_75t_L g945 ( 
.A(n_881),
.Y(n_945)
);

NAND2xp5_ASAP7_75t_L g946 ( 
.A(n_889),
.B(n_801),
.Y(n_946)
);

NAND2xp5_ASAP7_75t_L g947 ( 
.A(n_889),
.B(n_801),
.Y(n_947)
);

INVx1_ASAP7_75t_L g948 ( 
.A(n_922),
.Y(n_948)
);

INVx3_ASAP7_75t_L g949 ( 
.A(n_881),
.Y(n_949)
);

INVx1_ASAP7_75t_L g950 ( 
.A(n_922),
.Y(n_950)
);

AND2x6_ASAP7_75t_L g951 ( 
.A(n_904),
.B(n_643),
.Y(n_951)
);

INVx1_ASAP7_75t_L g952 ( 
.A(n_924),
.Y(n_952)
);

INVx2_ASAP7_75t_L g953 ( 
.A(n_873),
.Y(n_953)
);

INVx1_ASAP7_75t_L g954 ( 
.A(n_924),
.Y(n_954)
);

NOR2xp33_ASAP7_75t_L g955 ( 
.A(n_887),
.B(n_858),
.Y(n_955)
);

BUFx6f_ASAP7_75t_L g956 ( 
.A(n_881),
.Y(n_956)
);

AND2x2_ASAP7_75t_L g957 ( 
.A(n_904),
.B(n_823),
.Y(n_957)
);

NAND2xp5_ASAP7_75t_L g958 ( 
.A(n_889),
.B(n_830),
.Y(n_958)
);

HB1xp67_ASAP7_75t_L g959 ( 
.A(n_902),
.Y(n_959)
);

BUFx6f_ASAP7_75t_L g960 ( 
.A(n_891),
.Y(n_960)
);

INVx2_ASAP7_75t_L g961 ( 
.A(n_876),
.Y(n_961)
);

INVx1_ASAP7_75t_L g962 ( 
.A(n_925),
.Y(n_962)
);

BUFx2_ASAP7_75t_L g963 ( 
.A(n_879),
.Y(n_963)
);

AND2x4_ASAP7_75t_L g964 ( 
.A(n_889),
.B(n_837),
.Y(n_964)
);

INVx1_ASAP7_75t_L g965 ( 
.A(n_925),
.Y(n_965)
);

BUFx6f_ASAP7_75t_L g966 ( 
.A(n_891),
.Y(n_966)
);

INVx1_ASAP7_75t_L g967 ( 
.A(n_896),
.Y(n_967)
);

INVx1_ASAP7_75t_L g968 ( 
.A(n_896),
.Y(n_968)
);

XOR2xp5_ASAP7_75t_L g969 ( 
.A(n_932),
.B(n_840),
.Y(n_969)
);

CKINVDCx5p33_ASAP7_75t_R g970 ( 
.A(n_892),
.Y(n_970)
);

NAND2xp5_ASAP7_75t_L g971 ( 
.A(n_929),
.B(n_830),
.Y(n_971)
);

INVx2_ASAP7_75t_L g972 ( 
.A(n_876),
.Y(n_972)
);

INVx2_ASAP7_75t_L g973 ( 
.A(n_878),
.Y(n_973)
);

INVx2_ASAP7_75t_L g974 ( 
.A(n_878),
.Y(n_974)
);

CKINVDCx5p33_ASAP7_75t_R g975 ( 
.A(n_917),
.Y(n_975)
);

INVx1_ASAP7_75t_L g976 ( 
.A(n_927),
.Y(n_976)
);

INVx1_ASAP7_75t_L g977 ( 
.A(n_927),
.Y(n_977)
);

CKINVDCx5p33_ASAP7_75t_R g978 ( 
.A(n_918),
.Y(n_978)
);

BUFx6f_ASAP7_75t_L g979 ( 
.A(n_891),
.Y(n_979)
);

CKINVDCx5p33_ASAP7_75t_R g980 ( 
.A(n_882),
.Y(n_980)
);

OA21x2_ASAP7_75t_L g981 ( 
.A1(n_883),
.A2(n_710),
.B(n_643),
.Y(n_981)
);

INVx2_ASAP7_75t_L g982 ( 
.A(n_872),
.Y(n_982)
);

INVx2_ASAP7_75t_L g983 ( 
.A(n_872),
.Y(n_983)
);

NAND2xp5_ASAP7_75t_L g984 ( 
.A(n_929),
.B(n_837),
.Y(n_984)
);

CKINVDCx20_ASAP7_75t_R g985 ( 
.A(n_903),
.Y(n_985)
);

INVx1_ASAP7_75t_L g986 ( 
.A(n_928),
.Y(n_986)
);

INVx1_ASAP7_75t_L g987 ( 
.A(n_928),
.Y(n_987)
);

INVx1_ASAP7_75t_L g988 ( 
.A(n_931),
.Y(n_988)
);

INVx1_ASAP7_75t_L g989 ( 
.A(n_931),
.Y(n_989)
);

CKINVDCx5p33_ASAP7_75t_R g990 ( 
.A(n_895),
.Y(n_990)
);

INVx2_ASAP7_75t_L g991 ( 
.A(n_872),
.Y(n_991)
);

CKINVDCx5p33_ASAP7_75t_R g992 ( 
.A(n_895),
.Y(n_992)
);

NAND2xp5_ASAP7_75t_SL g993 ( 
.A(n_893),
.B(n_809),
.Y(n_993)
);

BUFx3_ASAP7_75t_L g994 ( 
.A(n_872),
.Y(n_994)
);

CKINVDCx20_ASAP7_75t_R g995 ( 
.A(n_882),
.Y(n_995)
);

CKINVDCx20_ASAP7_75t_R g996 ( 
.A(n_886),
.Y(n_996)
);

INVx1_ASAP7_75t_L g997 ( 
.A(n_870),
.Y(n_997)
);

NAND2xp33_ASAP7_75t_R g998 ( 
.A(n_885),
.B(n_840),
.Y(n_998)
);

AND2x4_ASAP7_75t_L g999 ( 
.A(n_929),
.B(n_865),
.Y(n_999)
);

INVx1_ASAP7_75t_L g1000 ( 
.A(n_870),
.Y(n_1000)
);

CKINVDCx5p33_ASAP7_75t_R g1001 ( 
.A(n_893),
.Y(n_1001)
);

INVx2_ASAP7_75t_L g1002 ( 
.A(n_872),
.Y(n_1002)
);

AND2x2_ASAP7_75t_L g1003 ( 
.A(n_929),
.B(n_838),
.Y(n_1003)
);

INVx1_ASAP7_75t_L g1004 ( 
.A(n_875),
.Y(n_1004)
);

HB1xp67_ASAP7_75t_L g1005 ( 
.A(n_886),
.Y(n_1005)
);

AND2x2_ASAP7_75t_L g1006 ( 
.A(n_929),
.B(n_771),
.Y(n_1006)
);

INVxp67_ASAP7_75t_SL g1007 ( 
.A(n_884),
.Y(n_1007)
);

INVx2_ASAP7_75t_L g1008 ( 
.A(n_872),
.Y(n_1008)
);

HB1xp67_ASAP7_75t_L g1009 ( 
.A(n_886),
.Y(n_1009)
);

CKINVDCx5p33_ASAP7_75t_R g1010 ( 
.A(n_910),
.Y(n_1010)
);

INVx1_ASAP7_75t_L g1011 ( 
.A(n_875),
.Y(n_1011)
);

INVx1_ASAP7_75t_L g1012 ( 
.A(n_930),
.Y(n_1012)
);

HB1xp67_ASAP7_75t_L g1013 ( 
.A(n_929),
.Y(n_1013)
);

INVx1_ASAP7_75t_L g1014 ( 
.A(n_930),
.Y(n_1014)
);

CKINVDCx20_ASAP7_75t_R g1015 ( 
.A(n_877),
.Y(n_1015)
);

CKINVDCx5p33_ASAP7_75t_R g1016 ( 
.A(n_910),
.Y(n_1016)
);

INVx1_ASAP7_75t_L g1017 ( 
.A(n_930),
.Y(n_1017)
);

CKINVDCx5p33_ASAP7_75t_R g1018 ( 
.A(n_910),
.Y(n_1018)
);

INVxp67_ASAP7_75t_L g1019 ( 
.A(n_901),
.Y(n_1019)
);

NAND2xp5_ASAP7_75t_L g1020 ( 
.A(n_890),
.B(n_809),
.Y(n_1020)
);

AND2x2_ASAP7_75t_L g1021 ( 
.A(n_877),
.B(n_771),
.Y(n_1021)
);

AND2x4_ASAP7_75t_L g1022 ( 
.A(n_900),
.B(n_851),
.Y(n_1022)
);

INVx1_ASAP7_75t_L g1023 ( 
.A(n_930),
.Y(n_1023)
);

INVx2_ASAP7_75t_L g1024 ( 
.A(n_940),
.Y(n_1024)
);

AO22x2_ASAP7_75t_L g1025 ( 
.A1(n_942),
.A2(n_842),
.B1(n_857),
.B2(n_814),
.Y(n_1025)
);

INVx6_ASAP7_75t_L g1026 ( 
.A(n_1022),
.Y(n_1026)
);

NAND2xp5_ASAP7_75t_L g1027 ( 
.A(n_1019),
.B(n_893),
.Y(n_1027)
);

NAND2xp5_ASAP7_75t_SL g1028 ( 
.A(n_1010),
.B(n_893),
.Y(n_1028)
);

INVx2_ASAP7_75t_L g1029 ( 
.A(n_940),
.Y(n_1029)
);

INVx1_ASAP7_75t_L g1030 ( 
.A(n_953),
.Y(n_1030)
);

NAND2xp5_ASAP7_75t_SL g1031 ( 
.A(n_1016),
.B(n_920),
.Y(n_1031)
);

INVx1_ASAP7_75t_L g1032 ( 
.A(n_953),
.Y(n_1032)
);

INVx2_ASAP7_75t_L g1033 ( 
.A(n_961),
.Y(n_1033)
);

INVx4_ASAP7_75t_L g1034 ( 
.A(n_990),
.Y(n_1034)
);

AOI22xp33_ASAP7_75t_L g1035 ( 
.A1(n_951),
.A2(n_803),
.B1(n_792),
.B2(n_919),
.Y(n_1035)
);

INVx3_ASAP7_75t_L g1036 ( 
.A(n_937),
.Y(n_1036)
);

INVx1_ASAP7_75t_SL g1037 ( 
.A(n_963),
.Y(n_1037)
);

BUFx6f_ASAP7_75t_L g1038 ( 
.A(n_994),
.Y(n_1038)
);

OR2x6_ASAP7_75t_L g1039 ( 
.A(n_959),
.B(n_1005),
.Y(n_1039)
);

BUFx2_ASAP7_75t_L g1040 ( 
.A(n_943),
.Y(n_1040)
);

AOI22xp5_ASAP7_75t_L g1041 ( 
.A1(n_955),
.A2(n_926),
.B1(n_906),
.B2(n_920),
.Y(n_1041)
);

INVx4_ASAP7_75t_SL g1042 ( 
.A(n_951),
.Y(n_1042)
);

INVx3_ASAP7_75t_L g1043 ( 
.A(n_937),
.Y(n_1043)
);

XNOR2xp5_ASAP7_75t_L g1044 ( 
.A(n_969),
.B(n_863),
.Y(n_1044)
);

INVx6_ASAP7_75t_L g1045 ( 
.A(n_1022),
.Y(n_1045)
);

INVx2_ASAP7_75t_L g1046 ( 
.A(n_961),
.Y(n_1046)
);

INVx2_ASAP7_75t_L g1047 ( 
.A(n_972),
.Y(n_1047)
);

INVx2_ASAP7_75t_L g1048 ( 
.A(n_972),
.Y(n_1048)
);

CKINVDCx5p33_ASAP7_75t_R g1049 ( 
.A(n_938),
.Y(n_1049)
);

AND2x2_ASAP7_75t_SL g1050 ( 
.A(n_957),
.B(n_1009),
.Y(n_1050)
);

NOR2xp33_ASAP7_75t_L g1051 ( 
.A(n_992),
.B(n_858),
.Y(n_1051)
);

INVx3_ASAP7_75t_L g1052 ( 
.A(n_973),
.Y(n_1052)
);

AND2x6_ASAP7_75t_L g1053 ( 
.A(n_964),
.B(n_906),
.Y(n_1053)
);

AOI22xp5_ASAP7_75t_L g1054 ( 
.A1(n_955),
.A2(n_906),
.B1(n_920),
.B2(n_654),
.Y(n_1054)
);

INVx2_ASAP7_75t_L g1055 ( 
.A(n_973),
.Y(n_1055)
);

INVx2_ASAP7_75t_L g1056 ( 
.A(n_974),
.Y(n_1056)
);

INVx2_ASAP7_75t_L g1057 ( 
.A(n_974),
.Y(n_1057)
);

INVxp33_ASAP7_75t_L g1058 ( 
.A(n_1021),
.Y(n_1058)
);

INVxp67_ASAP7_75t_SL g1059 ( 
.A(n_994),
.Y(n_1059)
);

INVx1_ASAP7_75t_L g1060 ( 
.A(n_997),
.Y(n_1060)
);

INVx1_ASAP7_75t_L g1061 ( 
.A(n_1000),
.Y(n_1061)
);

INVx1_ASAP7_75t_L g1062 ( 
.A(n_1004),
.Y(n_1062)
);

NAND2xp5_ASAP7_75t_L g1063 ( 
.A(n_964),
.B(n_920),
.Y(n_1063)
);

NOR2xp33_ASAP7_75t_L g1064 ( 
.A(n_958),
.B(n_863),
.Y(n_1064)
);

BUFx6f_ASAP7_75t_L g1065 ( 
.A(n_960),
.Y(n_1065)
);

INVx1_ASAP7_75t_L g1066 ( 
.A(n_1011),
.Y(n_1066)
);

NAND2xp5_ASAP7_75t_L g1067 ( 
.A(n_964),
.B(n_919),
.Y(n_1067)
);

INVx2_ASAP7_75t_L g1068 ( 
.A(n_934),
.Y(n_1068)
);

INVx4_ASAP7_75t_L g1069 ( 
.A(n_1018),
.Y(n_1069)
);

NAND2xp33_ASAP7_75t_L g1070 ( 
.A(n_1001),
.B(n_874),
.Y(n_1070)
);

OR2x6_ASAP7_75t_L g1071 ( 
.A(n_1022),
.B(n_906),
.Y(n_1071)
);

NAND2xp33_ASAP7_75t_L g1072 ( 
.A(n_1001),
.B(n_874),
.Y(n_1072)
);

INVx2_ASAP7_75t_SL g1073 ( 
.A(n_1015),
.Y(n_1073)
);

BUFx10_ASAP7_75t_L g1074 ( 
.A(n_941),
.Y(n_1074)
);

INVx3_ASAP7_75t_L g1075 ( 
.A(n_960),
.Y(n_1075)
);

INVx2_ASAP7_75t_L g1076 ( 
.A(n_939),
.Y(n_1076)
);

BUFx10_ASAP7_75t_L g1077 ( 
.A(n_970),
.Y(n_1077)
);

INVx1_ASAP7_75t_L g1078 ( 
.A(n_967),
.Y(n_1078)
);

NAND2xp5_ASAP7_75t_SL g1079 ( 
.A(n_971),
.B(n_899),
.Y(n_1079)
);

INVx1_ASAP7_75t_L g1080 ( 
.A(n_968),
.Y(n_1080)
);

BUFx3_ASAP7_75t_L g1081 ( 
.A(n_975),
.Y(n_1081)
);

AOI22xp33_ASAP7_75t_L g1082 ( 
.A1(n_951),
.A2(n_803),
.B1(n_792),
.B2(n_919),
.Y(n_1082)
);

INVx1_ASAP7_75t_L g1083 ( 
.A(n_948),
.Y(n_1083)
);

OAI22xp5_ASAP7_75t_L g1084 ( 
.A1(n_976),
.A2(n_888),
.B1(n_654),
.B2(n_671),
.Y(n_1084)
);

INVx2_ASAP7_75t_L g1085 ( 
.A(n_950),
.Y(n_1085)
);

NAND2xp5_ASAP7_75t_SL g1086 ( 
.A(n_946),
.B(n_947),
.Y(n_1086)
);

NOR2xp33_ASAP7_75t_L g1087 ( 
.A(n_1020),
.B(n_820),
.Y(n_1087)
);

NAND2xp5_ASAP7_75t_SL g1088 ( 
.A(n_1003),
.B(n_899),
.Y(n_1088)
);

INVx2_ASAP7_75t_L g1089 ( 
.A(n_952),
.Y(n_1089)
);

INVx1_ASAP7_75t_L g1090 ( 
.A(n_954),
.Y(n_1090)
);

NAND2xp5_ASAP7_75t_SL g1091 ( 
.A(n_993),
.B(n_1006),
.Y(n_1091)
);

INVx2_ASAP7_75t_L g1092 ( 
.A(n_962),
.Y(n_1092)
);

BUFx3_ASAP7_75t_L g1093 ( 
.A(n_978),
.Y(n_1093)
);

INVx2_ASAP7_75t_L g1094 ( 
.A(n_965),
.Y(n_1094)
);

NAND2xp5_ASAP7_75t_L g1095 ( 
.A(n_999),
.B(n_919),
.Y(n_1095)
);

AND2x6_ASAP7_75t_L g1096 ( 
.A(n_999),
.B(n_900),
.Y(n_1096)
);

BUFx6f_ASAP7_75t_L g1097 ( 
.A(n_960),
.Y(n_1097)
);

INVx4_ASAP7_75t_L g1098 ( 
.A(n_951),
.Y(n_1098)
);

XNOR2xp5_ASAP7_75t_L g1099 ( 
.A(n_942),
.B(n_985),
.Y(n_1099)
);

INVx5_ASAP7_75t_L g1100 ( 
.A(n_951),
.Y(n_1100)
);

AND2x4_ASAP7_75t_SL g1101 ( 
.A(n_1015),
.B(n_996),
.Y(n_1101)
);

BUFx6f_ASAP7_75t_SL g1102 ( 
.A(n_999),
.Y(n_1102)
);

NOR2xp33_ASAP7_75t_L g1103 ( 
.A(n_993),
.B(n_888),
.Y(n_1103)
);

INVx4_ASAP7_75t_L g1104 ( 
.A(n_960),
.Y(n_1104)
);

INVx2_ASAP7_75t_L g1105 ( 
.A(n_982),
.Y(n_1105)
);

O2A1O1Ixp33_ASAP7_75t_L g1106 ( 
.A1(n_977),
.A2(n_909),
.B(n_911),
.C(n_905),
.Y(n_1106)
);

INVx2_ASAP7_75t_L g1107 ( 
.A(n_982),
.Y(n_1107)
);

INVx2_ASAP7_75t_L g1108 ( 
.A(n_983),
.Y(n_1108)
);

NOR2xp33_ASAP7_75t_L g1109 ( 
.A(n_986),
.B(n_888),
.Y(n_1109)
);

NAND2xp5_ASAP7_75t_L g1110 ( 
.A(n_987),
.B(n_933),
.Y(n_1110)
);

BUFx6f_ASAP7_75t_L g1111 ( 
.A(n_966),
.Y(n_1111)
);

INVx1_ASAP7_75t_L g1112 ( 
.A(n_988),
.Y(n_1112)
);

NOR2xp33_ASAP7_75t_L g1113 ( 
.A(n_989),
.B(n_888),
.Y(n_1113)
);

INVx1_ASAP7_75t_L g1114 ( 
.A(n_1023),
.Y(n_1114)
);

INVx5_ASAP7_75t_L g1115 ( 
.A(n_966),
.Y(n_1115)
);

INVx1_ASAP7_75t_L g1116 ( 
.A(n_1012),
.Y(n_1116)
);

INVx2_ASAP7_75t_L g1117 ( 
.A(n_983),
.Y(n_1117)
);

INVx2_ASAP7_75t_L g1118 ( 
.A(n_991),
.Y(n_1118)
);

INVx5_ASAP7_75t_L g1119 ( 
.A(n_966),
.Y(n_1119)
);

INVx2_ASAP7_75t_L g1120 ( 
.A(n_991),
.Y(n_1120)
);

BUFx10_ASAP7_75t_L g1121 ( 
.A(n_966),
.Y(n_1121)
);

NAND2xp5_ASAP7_75t_SL g1122 ( 
.A(n_984),
.B(n_899),
.Y(n_1122)
);

INVx4_ASAP7_75t_SL g1123 ( 
.A(n_979),
.Y(n_1123)
);

OR2x6_ASAP7_75t_L g1124 ( 
.A(n_996),
.B(n_900),
.Y(n_1124)
);

INVx1_ASAP7_75t_L g1125 ( 
.A(n_1014),
.Y(n_1125)
);

NAND2xp5_ASAP7_75t_SL g1126 ( 
.A(n_979),
.B(n_899),
.Y(n_1126)
);

INVx1_ASAP7_75t_L g1127 ( 
.A(n_1017),
.Y(n_1127)
);

INVx4_ASAP7_75t_L g1128 ( 
.A(n_979),
.Y(n_1128)
);

INVx1_ASAP7_75t_L g1129 ( 
.A(n_1007),
.Y(n_1129)
);

INVx1_ASAP7_75t_SL g1130 ( 
.A(n_985),
.Y(n_1130)
);

INVx2_ASAP7_75t_L g1131 ( 
.A(n_1002),
.Y(n_1131)
);

NOR2xp33_ASAP7_75t_L g1132 ( 
.A(n_1013),
.B(n_916),
.Y(n_1132)
);

INVx3_ASAP7_75t_L g1133 ( 
.A(n_979),
.Y(n_1133)
);

OAI22xp5_ASAP7_75t_L g1134 ( 
.A1(n_1002),
.A2(n_671),
.B1(n_757),
.B2(n_638),
.Y(n_1134)
);

INVx1_ASAP7_75t_L g1135 ( 
.A(n_1008),
.Y(n_1135)
);

INVx2_ASAP7_75t_L g1136 ( 
.A(n_1008),
.Y(n_1136)
);

OR2x6_ASAP7_75t_L g1137 ( 
.A(n_998),
.B(n_900),
.Y(n_1137)
);

INVx1_ASAP7_75t_L g1138 ( 
.A(n_945),
.Y(n_1138)
);

CKINVDCx20_ASAP7_75t_R g1139 ( 
.A(n_995),
.Y(n_1139)
);

INVx2_ASAP7_75t_L g1140 ( 
.A(n_945),
.Y(n_1140)
);

AOI22xp33_ASAP7_75t_L g1141 ( 
.A1(n_949),
.A2(n_933),
.B1(n_880),
.B2(n_930),
.Y(n_1141)
);

INVx2_ASAP7_75t_L g1142 ( 
.A(n_949),
.Y(n_1142)
);

INVxp67_ASAP7_75t_SL g1143 ( 
.A(n_935),
.Y(n_1143)
);

BUFx3_ASAP7_75t_L g1144 ( 
.A(n_995),
.Y(n_1144)
);

INVx2_ASAP7_75t_SL g1145 ( 
.A(n_981),
.Y(n_1145)
);

NOR2xp33_ASAP7_75t_L g1146 ( 
.A(n_935),
.B(n_933),
.Y(n_1146)
);

INVx6_ASAP7_75t_L g1147 ( 
.A(n_935),
.Y(n_1147)
);

INVx1_ASAP7_75t_L g1148 ( 
.A(n_935),
.Y(n_1148)
);

INVx1_ASAP7_75t_L g1149 ( 
.A(n_936),
.Y(n_1149)
);

INVx1_ASAP7_75t_L g1150 ( 
.A(n_936),
.Y(n_1150)
);

INVx2_ASAP7_75t_L g1151 ( 
.A(n_936),
.Y(n_1151)
);

INVx1_ASAP7_75t_L g1152 ( 
.A(n_936),
.Y(n_1152)
);

OAI22xp5_ASAP7_75t_L g1153 ( 
.A1(n_998),
.A2(n_757),
.B1(n_646),
.B2(n_559),
.Y(n_1153)
);

INVx2_ASAP7_75t_SL g1154 ( 
.A(n_981),
.Y(n_1154)
);

BUFx6f_ASAP7_75t_L g1155 ( 
.A(n_944),
.Y(n_1155)
);

INVx2_ASAP7_75t_L g1156 ( 
.A(n_944),
.Y(n_1156)
);

BUFx4f_ASAP7_75t_L g1157 ( 
.A(n_944),
.Y(n_1157)
);

NAND3xp33_ASAP7_75t_L g1158 ( 
.A(n_944),
.B(n_930),
.C(n_874),
.Y(n_1158)
);

NOR2xp33_ASAP7_75t_L g1159 ( 
.A(n_956),
.B(n_933),
.Y(n_1159)
);

NAND2xp5_ASAP7_75t_SL g1160 ( 
.A(n_956),
.B(n_890),
.Y(n_1160)
);

BUFx4f_ASAP7_75t_L g1161 ( 
.A(n_956),
.Y(n_1161)
);

INVx3_ASAP7_75t_L g1162 ( 
.A(n_956),
.Y(n_1162)
);

INVx2_ASAP7_75t_L g1163 ( 
.A(n_1052),
.Y(n_1163)
);

INVx2_ASAP7_75t_SL g1164 ( 
.A(n_1037),
.Y(n_1164)
);

INVx2_ASAP7_75t_SL g1165 ( 
.A(n_1081),
.Y(n_1165)
);

NAND2xp33_ASAP7_75t_L g1166 ( 
.A(n_1053),
.B(n_874),
.Y(n_1166)
);

INVx4_ASAP7_75t_L g1167 ( 
.A(n_1026),
.Y(n_1167)
);

NAND2xp5_ASAP7_75t_SL g1168 ( 
.A(n_1069),
.B(n_890),
.Y(n_1168)
);

BUFx10_ASAP7_75t_L g1169 ( 
.A(n_1051),
.Y(n_1169)
);

BUFx10_ASAP7_75t_L g1170 ( 
.A(n_1049),
.Y(n_1170)
);

INVx1_ASAP7_75t_L g1171 ( 
.A(n_1030),
.Y(n_1171)
);

AND2x4_ASAP7_75t_L g1172 ( 
.A(n_1071),
.B(n_898),
.Y(n_1172)
);

BUFx6f_ASAP7_75t_L g1173 ( 
.A(n_1038),
.Y(n_1173)
);

BUFx3_ASAP7_75t_L g1174 ( 
.A(n_1093),
.Y(n_1174)
);

INVx1_ASAP7_75t_L g1175 ( 
.A(n_1078),
.Y(n_1175)
);

AND2x4_ASAP7_75t_L g1176 ( 
.A(n_1071),
.B(n_898),
.Y(n_1176)
);

INVx2_ASAP7_75t_L g1177 ( 
.A(n_1052),
.Y(n_1177)
);

BUFx6f_ASAP7_75t_L g1178 ( 
.A(n_1038),
.Y(n_1178)
);

INVx1_ASAP7_75t_L g1179 ( 
.A(n_1080),
.Y(n_1179)
);

AND2x4_ASAP7_75t_L g1180 ( 
.A(n_1042),
.B(n_890),
.Y(n_1180)
);

NAND2x1_ASAP7_75t_L g1181 ( 
.A(n_1098),
.B(n_981),
.Y(n_1181)
);

INVx2_ASAP7_75t_L g1182 ( 
.A(n_1030),
.Y(n_1182)
);

AND2x4_ASAP7_75t_L g1183 ( 
.A(n_1042),
.B(n_905),
.Y(n_1183)
);

AND2x6_ASAP7_75t_L g1184 ( 
.A(n_1036),
.B(n_710),
.Y(n_1184)
);

NAND2xp5_ASAP7_75t_SL g1185 ( 
.A(n_1069),
.B(n_874),
.Y(n_1185)
);

AND2x6_ASAP7_75t_L g1186 ( 
.A(n_1036),
.B(n_884),
.Y(n_1186)
);

AND2x4_ASAP7_75t_L g1187 ( 
.A(n_1137),
.B(n_905),
.Y(n_1187)
);

INVx1_ASAP7_75t_L g1188 ( 
.A(n_1060),
.Y(n_1188)
);

INVx2_ASAP7_75t_L g1189 ( 
.A(n_1032),
.Y(n_1189)
);

INVx1_ASAP7_75t_L g1190 ( 
.A(n_1060),
.Y(n_1190)
);

INVx2_ASAP7_75t_L g1191 ( 
.A(n_1032),
.Y(n_1191)
);

NAND2xp5_ASAP7_75t_L g1192 ( 
.A(n_1027),
.B(n_884),
.Y(n_1192)
);

INVx3_ASAP7_75t_L g1193 ( 
.A(n_1121),
.Y(n_1193)
);

INVx4_ASAP7_75t_L g1194 ( 
.A(n_1026),
.Y(n_1194)
);

INVx1_ASAP7_75t_L g1195 ( 
.A(n_1061),
.Y(n_1195)
);

NAND2x1p5_ASAP7_75t_L g1196 ( 
.A(n_1043),
.B(n_884),
.Y(n_1196)
);

INVx1_ASAP7_75t_L g1197 ( 
.A(n_1061),
.Y(n_1197)
);

INVx1_ASAP7_75t_L g1198 ( 
.A(n_1062),
.Y(n_1198)
);

INVx1_ASAP7_75t_L g1199 ( 
.A(n_1062),
.Y(n_1199)
);

AND2x4_ASAP7_75t_L g1200 ( 
.A(n_1137),
.B(n_1039),
.Y(n_1200)
);

NAND2xp5_ASAP7_75t_SL g1201 ( 
.A(n_1041),
.B(n_874),
.Y(n_1201)
);

INVx3_ASAP7_75t_L g1202 ( 
.A(n_1121),
.Y(n_1202)
);

INVx2_ASAP7_75t_L g1203 ( 
.A(n_1135),
.Y(n_1203)
);

INVx1_ASAP7_75t_L g1204 ( 
.A(n_1066),
.Y(n_1204)
);

INVx1_ASAP7_75t_L g1205 ( 
.A(n_1066),
.Y(n_1205)
);

INVx4_ASAP7_75t_L g1206 ( 
.A(n_1045),
.Y(n_1206)
);

BUFx3_ASAP7_75t_L g1207 ( 
.A(n_1040),
.Y(n_1207)
);

INVx3_ASAP7_75t_L g1208 ( 
.A(n_1038),
.Y(n_1208)
);

INVx1_ASAP7_75t_L g1209 ( 
.A(n_1112),
.Y(n_1209)
);

NAND2x1p5_ASAP7_75t_L g1210 ( 
.A(n_1043),
.B(n_905),
.Y(n_1210)
);

INVx1_ASAP7_75t_L g1211 ( 
.A(n_1112),
.Y(n_1211)
);

CKINVDCx5p33_ASAP7_75t_R g1212 ( 
.A(n_1074),
.Y(n_1212)
);

INVx2_ASAP7_75t_L g1213 ( 
.A(n_1135),
.Y(n_1213)
);

INVx1_ASAP7_75t_L g1214 ( 
.A(n_1083),
.Y(n_1214)
);

OAI221xp5_ASAP7_75t_L g1215 ( 
.A1(n_1054),
.A2(n_819),
.B1(n_566),
.B2(n_569),
.C(n_560),
.Y(n_1215)
);

NAND2x1p5_ASAP7_75t_L g1216 ( 
.A(n_1100),
.B(n_911),
.Y(n_1216)
);

CKINVDCx5p33_ASAP7_75t_R g1217 ( 
.A(n_1074),
.Y(n_1217)
);

INVx1_ASAP7_75t_L g1218 ( 
.A(n_1083),
.Y(n_1218)
);

NOR2xp33_ASAP7_75t_L g1219 ( 
.A(n_1153),
.B(n_857),
.Y(n_1219)
);

INVx1_ASAP7_75t_L g1220 ( 
.A(n_1090),
.Y(n_1220)
);

INVx2_ASAP7_75t_SL g1221 ( 
.A(n_1101),
.Y(n_1221)
);

INVx1_ASAP7_75t_L g1222 ( 
.A(n_1090),
.Y(n_1222)
);

INVx2_ASAP7_75t_L g1223 ( 
.A(n_1024),
.Y(n_1223)
);

INVxp67_ASAP7_75t_L g1224 ( 
.A(n_1073),
.Y(n_1224)
);

INVx1_ASAP7_75t_L g1225 ( 
.A(n_1029),
.Y(n_1225)
);

CKINVDCx5p33_ASAP7_75t_R g1226 ( 
.A(n_1077),
.Y(n_1226)
);

INVx2_ASAP7_75t_SL g1227 ( 
.A(n_1077),
.Y(n_1227)
);

INVx1_ASAP7_75t_L g1228 ( 
.A(n_1068),
.Y(n_1228)
);

INVx1_ASAP7_75t_L g1229 ( 
.A(n_1076),
.Y(n_1229)
);

BUFx6f_ASAP7_75t_L g1230 ( 
.A(n_1065),
.Y(n_1230)
);

CKINVDCx5p33_ASAP7_75t_R g1231 ( 
.A(n_1044),
.Y(n_1231)
);

INVxp67_ASAP7_75t_L g1232 ( 
.A(n_1134),
.Y(n_1232)
);

NAND2xp5_ASAP7_75t_SL g1233 ( 
.A(n_1034),
.B(n_911),
.Y(n_1233)
);

INVxp67_ASAP7_75t_L g1234 ( 
.A(n_1064),
.Y(n_1234)
);

INVx1_ASAP7_75t_L g1235 ( 
.A(n_1085),
.Y(n_1235)
);

INVx1_ASAP7_75t_SL g1236 ( 
.A(n_1039),
.Y(n_1236)
);

NAND2x1p5_ASAP7_75t_L g1237 ( 
.A(n_1100),
.B(n_911),
.Y(n_1237)
);

NAND3xp33_ASAP7_75t_L g1238 ( 
.A(n_1084),
.B(n_605),
.C(n_588),
.Y(n_1238)
);

INVx1_ASAP7_75t_L g1239 ( 
.A(n_1089),
.Y(n_1239)
);

BUFx2_ASAP7_75t_L g1240 ( 
.A(n_1045),
.Y(n_1240)
);

NOR3xp33_ASAP7_75t_L g1241 ( 
.A(n_1034),
.B(n_570),
.C(n_539),
.Y(n_1241)
);

INVx2_ASAP7_75t_L g1242 ( 
.A(n_1033),
.Y(n_1242)
);

AND2x6_ASAP7_75t_L g1243 ( 
.A(n_1150),
.B(n_617),
.Y(n_1243)
);

INVx1_ASAP7_75t_L g1244 ( 
.A(n_1092),
.Y(n_1244)
);

INVx1_ASAP7_75t_L g1245 ( 
.A(n_1094),
.Y(n_1245)
);

HB1xp67_ASAP7_75t_L g1246 ( 
.A(n_1124),
.Y(n_1246)
);

NAND2xp5_ASAP7_75t_L g1247 ( 
.A(n_1132),
.B(n_891),
.Y(n_1247)
);

INVxp67_ASAP7_75t_L g1248 ( 
.A(n_1124),
.Y(n_1248)
);

INVx2_ASAP7_75t_L g1249 ( 
.A(n_1046),
.Y(n_1249)
);

HB1xp67_ASAP7_75t_L g1250 ( 
.A(n_1102),
.Y(n_1250)
);

INVxp67_ASAP7_75t_L g1251 ( 
.A(n_1053),
.Y(n_1251)
);

INVx3_ASAP7_75t_L g1252 ( 
.A(n_1157),
.Y(n_1252)
);

INVx1_ASAP7_75t_L g1253 ( 
.A(n_1114),
.Y(n_1253)
);

AND2x2_ASAP7_75t_L g1254 ( 
.A(n_1058),
.B(n_894),
.Y(n_1254)
);

OR2x2_ASAP7_75t_L g1255 ( 
.A(n_1130),
.B(n_1087),
.Y(n_1255)
);

NAND2x1p5_ASAP7_75t_L g1256 ( 
.A(n_1100),
.B(n_894),
.Y(n_1256)
);

NAND2xp5_ASAP7_75t_L g1257 ( 
.A(n_1067),
.B(n_891),
.Y(n_1257)
);

OR2x6_ASAP7_75t_L g1258 ( 
.A(n_1144),
.B(n_897),
.Y(n_1258)
);

NAND2x1p5_ASAP7_75t_L g1259 ( 
.A(n_1050),
.B(n_897),
.Y(n_1259)
);

INVx2_ASAP7_75t_SL g1260 ( 
.A(n_1053),
.Y(n_1260)
);

INVx2_ASAP7_75t_L g1261 ( 
.A(n_1047),
.Y(n_1261)
);

CKINVDCx5p33_ASAP7_75t_R g1262 ( 
.A(n_1099),
.Y(n_1262)
);

INVx1_ASAP7_75t_L g1263 ( 
.A(n_1114),
.Y(n_1263)
);

INVx1_ASAP7_75t_L g1264 ( 
.A(n_1116),
.Y(n_1264)
);

AND2x4_ASAP7_75t_L g1265 ( 
.A(n_1053),
.B(n_907),
.Y(n_1265)
);

NAND2xp5_ASAP7_75t_L g1266 ( 
.A(n_1086),
.B(n_891),
.Y(n_1266)
);

BUFx2_ASAP7_75t_L g1267 ( 
.A(n_1096),
.Y(n_1267)
);

AO22x2_ASAP7_75t_L g1268 ( 
.A1(n_1025),
.A2(n_923),
.B1(n_1091),
.B2(n_1088),
.Y(n_1268)
);

INVx1_ASAP7_75t_L g1269 ( 
.A(n_1116),
.Y(n_1269)
);

INVx1_ASAP7_75t_L g1270 ( 
.A(n_1125),
.Y(n_1270)
);

BUFx2_ASAP7_75t_L g1271 ( 
.A(n_1096),
.Y(n_1271)
);

BUFx6f_ASAP7_75t_L g1272 ( 
.A(n_1065),
.Y(n_1272)
);

INVxp67_ASAP7_75t_L g1273 ( 
.A(n_1102),
.Y(n_1273)
);

INVx1_ASAP7_75t_L g1274 ( 
.A(n_1125),
.Y(n_1274)
);

INVx2_ASAP7_75t_L g1275 ( 
.A(n_1048),
.Y(n_1275)
);

INVxp67_ASAP7_75t_L g1276 ( 
.A(n_1095),
.Y(n_1276)
);

BUFx3_ASAP7_75t_L g1277 ( 
.A(n_1139),
.Y(n_1277)
);

NAND2xp5_ASAP7_75t_SL g1278 ( 
.A(n_1063),
.B(n_912),
.Y(n_1278)
);

INVx2_ASAP7_75t_L g1279 ( 
.A(n_1055),
.Y(n_1279)
);

INVx1_ASAP7_75t_L g1280 ( 
.A(n_1056),
.Y(n_1280)
);

AND2x4_ASAP7_75t_L g1281 ( 
.A(n_1098),
.B(n_907),
.Y(n_1281)
);

BUFx6f_ASAP7_75t_L g1282 ( 
.A(n_1065),
.Y(n_1282)
);

INVx2_ASAP7_75t_L g1283 ( 
.A(n_1057),
.Y(n_1283)
);

AND2x4_ASAP7_75t_L g1284 ( 
.A(n_1123),
.B(n_908),
.Y(n_1284)
);

INVx1_ASAP7_75t_L g1285 ( 
.A(n_1127),
.Y(n_1285)
);

NAND2xp5_ASAP7_75t_L g1286 ( 
.A(n_1129),
.B(n_1110),
.Y(n_1286)
);

INVx2_ASAP7_75t_L g1287 ( 
.A(n_1127),
.Y(n_1287)
);

INVx1_ASAP7_75t_SL g1288 ( 
.A(n_1025),
.Y(n_1288)
);

NAND2xp5_ASAP7_75t_SL g1289 ( 
.A(n_1035),
.B(n_912),
.Y(n_1289)
);

AND2x4_ASAP7_75t_L g1290 ( 
.A(n_1123),
.B(n_908),
.Y(n_1290)
);

AND2x4_ASAP7_75t_L g1291 ( 
.A(n_1096),
.B(n_915),
.Y(n_1291)
);

NAND2xp5_ASAP7_75t_L g1292 ( 
.A(n_1129),
.B(n_912),
.Y(n_1292)
);

HB1xp67_ASAP7_75t_L g1293 ( 
.A(n_1096),
.Y(n_1293)
);

INVx1_ASAP7_75t_SL g1294 ( 
.A(n_1126),
.Y(n_1294)
);

INVx1_ASAP7_75t_L g1295 ( 
.A(n_1138),
.Y(n_1295)
);

INVx5_ASAP7_75t_L g1296 ( 
.A(n_1097),
.Y(n_1296)
);

NOR2xp33_ASAP7_75t_L g1297 ( 
.A(n_1082),
.B(n_1079),
.Y(n_1297)
);

NOR2xp33_ASAP7_75t_L g1298 ( 
.A(n_1103),
.B(n_923),
.Y(n_1298)
);

INVx2_ASAP7_75t_L g1299 ( 
.A(n_1105),
.Y(n_1299)
);

INVx2_ASAP7_75t_L g1300 ( 
.A(n_1107),
.Y(n_1300)
);

INVx1_ASAP7_75t_L g1301 ( 
.A(n_1138),
.Y(n_1301)
);

NAND2x1p5_ASAP7_75t_L g1302 ( 
.A(n_1115),
.B(n_915),
.Y(n_1302)
);

BUFx3_ASAP7_75t_L g1303 ( 
.A(n_1147),
.Y(n_1303)
);

A2O1A1Ixp33_ASAP7_75t_L g1304 ( 
.A1(n_1106),
.A2(n_883),
.B(n_622),
.C(n_642),
.Y(n_1304)
);

BUFx6f_ASAP7_75t_L g1305 ( 
.A(n_1097),
.Y(n_1305)
);

OR2x2_ASAP7_75t_L g1306 ( 
.A(n_1160),
.B(n_980),
.Y(n_1306)
);

AND2x4_ASAP7_75t_L g1307 ( 
.A(n_1115),
.B(n_793),
.Y(n_1307)
);

HB1xp67_ASAP7_75t_L g1308 ( 
.A(n_1146),
.Y(n_1308)
);

INVx2_ASAP7_75t_L g1309 ( 
.A(n_1108),
.Y(n_1309)
);

INVx4_ASAP7_75t_SL g1310 ( 
.A(n_1147),
.Y(n_1310)
);

INVx2_ASAP7_75t_L g1311 ( 
.A(n_1117),
.Y(n_1311)
);

BUFx3_ASAP7_75t_L g1312 ( 
.A(n_1157),
.Y(n_1312)
);

OAI22xp33_ASAP7_75t_L g1313 ( 
.A1(n_1109),
.A2(n_584),
.B1(n_587),
.B2(n_576),
.Y(n_1313)
);

INVx2_ASAP7_75t_L g1314 ( 
.A(n_1118),
.Y(n_1314)
);

INVx2_ASAP7_75t_L g1315 ( 
.A(n_1120),
.Y(n_1315)
);

NAND2xp5_ASAP7_75t_L g1316 ( 
.A(n_1159),
.B(n_912),
.Y(n_1316)
);

AND2x2_ASAP7_75t_L g1317 ( 
.A(n_1113),
.B(n_795),
.Y(n_1317)
);

INVx1_ASAP7_75t_L g1318 ( 
.A(n_1131),
.Y(n_1318)
);

CKINVDCx5p33_ASAP7_75t_R g1319 ( 
.A(n_1097),
.Y(n_1319)
);

INVx2_ASAP7_75t_L g1320 ( 
.A(n_1136),
.Y(n_1320)
);

INVx2_ASAP7_75t_L g1321 ( 
.A(n_1140),
.Y(n_1321)
);

INVx1_ASAP7_75t_L g1322 ( 
.A(n_1142),
.Y(n_1322)
);

INVxp67_ASAP7_75t_L g1323 ( 
.A(n_1122),
.Y(n_1323)
);

AND2x2_ASAP7_75t_L g1324 ( 
.A(n_1141),
.B(n_796),
.Y(n_1324)
);

INVx1_ASAP7_75t_L g1325 ( 
.A(n_1150),
.Y(n_1325)
);

INVx1_ASAP7_75t_L g1326 ( 
.A(n_1152),
.Y(n_1326)
);

NAND2xp5_ASAP7_75t_L g1327 ( 
.A(n_1028),
.B(n_912),
.Y(n_1327)
);

INVx1_ASAP7_75t_L g1328 ( 
.A(n_1152),
.Y(n_1328)
);

AND2x6_ASAP7_75t_L g1329 ( 
.A(n_1075),
.B(n_623),
.Y(n_1329)
);

INVx1_ASAP7_75t_L g1330 ( 
.A(n_1148),
.Y(n_1330)
);

AND2x4_ASAP7_75t_L g1331 ( 
.A(n_1115),
.B(n_1119),
.Y(n_1331)
);

AND2x2_ASAP7_75t_L g1332 ( 
.A(n_1031),
.B(n_797),
.Y(n_1332)
);

NOR2xp33_ASAP7_75t_L g1333 ( 
.A(n_1149),
.B(n_980),
.Y(n_1333)
);

INVx1_ASAP7_75t_L g1334 ( 
.A(n_1151),
.Y(n_1334)
);

NOR2xp33_ASAP7_75t_L g1335 ( 
.A(n_1075),
.B(n_589),
.Y(n_1335)
);

OR2x2_ASAP7_75t_SL g1336 ( 
.A(n_1158),
.B(n_798),
.Y(n_1336)
);

INVx1_ASAP7_75t_L g1337 ( 
.A(n_1156),
.Y(n_1337)
);

AND2x4_ASAP7_75t_L g1338 ( 
.A(n_1119),
.B(n_799),
.Y(n_1338)
);

INVx1_ASAP7_75t_L g1339 ( 
.A(n_1133),
.Y(n_1339)
);

INVx2_ASAP7_75t_L g1340 ( 
.A(n_1162),
.Y(n_1340)
);

INVx1_ASAP7_75t_L g1341 ( 
.A(n_1133),
.Y(n_1341)
);

NOR2xp33_ASAP7_75t_L g1342 ( 
.A(n_1059),
.B(n_595),
.Y(n_1342)
);

INVx1_ASAP7_75t_L g1343 ( 
.A(n_1162),
.Y(n_1343)
);

AND2x4_ASAP7_75t_L g1344 ( 
.A(n_1119),
.B(n_1104),
.Y(n_1344)
);

NOR2xp33_ASAP7_75t_L g1345 ( 
.A(n_1104),
.B(n_611),
.Y(n_1345)
);

BUFx2_ASAP7_75t_L g1346 ( 
.A(n_1111),
.Y(n_1346)
);

NAND2xp5_ASAP7_75t_SL g1347 ( 
.A(n_1161),
.B(n_912),
.Y(n_1347)
);

INVx1_ASAP7_75t_L g1348 ( 
.A(n_1111),
.Y(n_1348)
);

OAI22xp5_ASAP7_75t_SL g1349 ( 
.A1(n_1128),
.A2(n_619),
.B1(n_620),
.B2(n_613),
.Y(n_1349)
);

OR2x2_ASAP7_75t_L g1350 ( 
.A(n_1111),
.B(n_804),
.Y(n_1350)
);

AOI22xp33_ASAP7_75t_L g1351 ( 
.A1(n_1128),
.A2(n_880),
.B1(n_914),
.B2(n_634),
.Y(n_1351)
);

INVx1_ASAP7_75t_L g1352 ( 
.A(n_1155),
.Y(n_1352)
);

CKINVDCx5p33_ASAP7_75t_R g1353 ( 
.A(n_1161),
.Y(n_1353)
);

INVx1_ASAP7_75t_L g1354 ( 
.A(n_1155),
.Y(n_1354)
);

NAND3xp33_ASAP7_75t_L g1355 ( 
.A(n_1070),
.B(n_728),
.C(n_690),
.Y(n_1355)
);

INVx2_ASAP7_75t_L g1356 ( 
.A(n_1155),
.Y(n_1356)
);

INVx1_ASAP7_75t_L g1357 ( 
.A(n_1145),
.Y(n_1357)
);

AO22x2_ASAP7_75t_L g1358 ( 
.A1(n_1154),
.A2(n_806),
.B1(n_807),
.B2(n_805),
.Y(n_1358)
);

INVx2_ASAP7_75t_L g1359 ( 
.A(n_1143),
.Y(n_1359)
);

INVx2_ASAP7_75t_L g1360 ( 
.A(n_1072),
.Y(n_1360)
);

INVx2_ASAP7_75t_L g1361 ( 
.A(n_1052),
.Y(n_1361)
);

HB1xp67_ASAP7_75t_L g1362 ( 
.A(n_1037),
.Y(n_1362)
);

BUFx3_ASAP7_75t_L g1363 ( 
.A(n_1081),
.Y(n_1363)
);

INVx2_ASAP7_75t_L g1364 ( 
.A(n_1052),
.Y(n_1364)
);

AND2x6_ASAP7_75t_L g1365 ( 
.A(n_1042),
.B(n_645),
.Y(n_1365)
);

NOR2xp33_ASAP7_75t_L g1366 ( 
.A(n_1234),
.B(n_626),
.Y(n_1366)
);

NAND2xp5_ASAP7_75t_L g1367 ( 
.A(n_1317),
.B(n_914),
.Y(n_1367)
);

AOI22xp5_ASAP7_75t_L g1368 ( 
.A1(n_1219),
.A2(n_640),
.B1(n_641),
.B2(n_636),
.Y(n_1368)
);

INVx2_ASAP7_75t_L g1369 ( 
.A(n_1182),
.Y(n_1369)
);

CKINVDCx5p33_ASAP7_75t_R g1370 ( 
.A(n_1212),
.Y(n_1370)
);

INVx1_ASAP7_75t_L g1371 ( 
.A(n_1188),
.Y(n_1371)
);

INVx2_ASAP7_75t_L g1372 ( 
.A(n_1189),
.Y(n_1372)
);

NAND2xp5_ASAP7_75t_L g1373 ( 
.A(n_1232),
.B(n_914),
.Y(n_1373)
);

AOI22xp33_ASAP7_75t_L g1374 ( 
.A1(n_1298),
.A2(n_914),
.B1(n_880),
.B2(n_659),
.Y(n_1374)
);

NAND2xp33_ASAP7_75t_SL g1375 ( 
.A(n_1353),
.B(n_662),
.Y(n_1375)
);

NAND2xp5_ASAP7_75t_L g1376 ( 
.A(n_1286),
.B(n_880),
.Y(n_1376)
);

NOR3x1_ASAP7_75t_L g1377 ( 
.A(n_1227),
.B(n_1215),
.C(n_1165),
.Y(n_1377)
);

INVx5_ASAP7_75t_L g1378 ( 
.A(n_1365),
.Y(n_1378)
);

NAND2xp5_ASAP7_75t_L g1379 ( 
.A(n_1190),
.B(n_914),
.Y(n_1379)
);

HB1xp67_ASAP7_75t_L g1380 ( 
.A(n_1362),
.Y(n_1380)
);

NAND2xp5_ASAP7_75t_L g1381 ( 
.A(n_1195),
.B(n_914),
.Y(n_1381)
);

AOI21xp5_ASAP7_75t_L g1382 ( 
.A1(n_1166),
.A2(n_738),
.B(n_720),
.Y(n_1382)
);

NAND2xp5_ASAP7_75t_L g1383 ( 
.A(n_1308),
.B(n_808),
.Y(n_1383)
);

NAND2xp5_ASAP7_75t_L g1384 ( 
.A(n_1276),
.B(n_810),
.Y(n_1384)
);

NAND2xp5_ASAP7_75t_L g1385 ( 
.A(n_1197),
.B(n_812),
.Y(n_1385)
);

NAND2xp5_ASAP7_75t_L g1386 ( 
.A(n_1198),
.B(n_815),
.Y(n_1386)
);

A2O1A1Ixp33_ASAP7_75t_L g1387 ( 
.A1(n_1297),
.A2(n_660),
.B(n_663),
.C(n_650),
.Y(n_1387)
);

AND3x1_ASAP7_75t_L g1388 ( 
.A(n_1241),
.B(n_817),
.C(n_816),
.Y(n_1388)
);

INVx1_ASAP7_75t_L g1389 ( 
.A(n_1199),
.Y(n_1389)
);

NOR2xp33_ASAP7_75t_L g1390 ( 
.A(n_1255),
.B(n_1169),
.Y(n_1390)
);

NAND2xp5_ASAP7_75t_L g1391 ( 
.A(n_1204),
.B(n_818),
.Y(n_1391)
);

NAND2xp5_ASAP7_75t_SL g1392 ( 
.A(n_1169),
.B(n_664),
.Y(n_1392)
);

NAND2xp5_ASAP7_75t_L g1393 ( 
.A(n_1205),
.B(n_821),
.Y(n_1393)
);

NAND2xp5_ASAP7_75t_SL g1394 ( 
.A(n_1164),
.B(n_668),
.Y(n_1394)
);

INVx3_ASAP7_75t_L g1395 ( 
.A(n_1331),
.Y(n_1395)
);

AND2x6_ASAP7_75t_SL g1396 ( 
.A(n_1258),
.B(n_825),
.Y(n_1396)
);

NAND2xp5_ASAP7_75t_L g1397 ( 
.A(n_1209),
.B(n_826),
.Y(n_1397)
);

NAND2xp5_ASAP7_75t_L g1398 ( 
.A(n_1211),
.B(n_827),
.Y(n_1398)
);

NAND2xp5_ASAP7_75t_L g1399 ( 
.A(n_1254),
.B(n_828),
.Y(n_1399)
);

AOI22xp33_ASAP7_75t_L g1400 ( 
.A1(n_1268),
.A2(n_1238),
.B1(n_1306),
.B2(n_1246),
.Y(n_1400)
);

INVx1_ASAP7_75t_L g1401 ( 
.A(n_1175),
.Y(n_1401)
);

NAND2xp5_ASAP7_75t_L g1402 ( 
.A(n_1172),
.B(n_829),
.Y(n_1402)
);

INVx2_ASAP7_75t_L g1403 ( 
.A(n_1191),
.Y(n_1403)
);

INVx1_ASAP7_75t_L g1404 ( 
.A(n_1179),
.Y(n_1404)
);

NAND2xp5_ASAP7_75t_L g1405 ( 
.A(n_1172),
.B(n_831),
.Y(n_1405)
);

INVx2_ASAP7_75t_SL g1406 ( 
.A(n_1174),
.Y(n_1406)
);

INVx2_ASAP7_75t_L g1407 ( 
.A(n_1203),
.Y(n_1407)
);

AOI22xp5_ASAP7_75t_L g1408 ( 
.A1(n_1176),
.A2(n_669),
.B1(n_674),
.B2(n_670),
.Y(n_1408)
);

INVx1_ASAP7_75t_L g1409 ( 
.A(n_1214),
.Y(n_1409)
);

BUFx6f_ASAP7_75t_L g1410 ( 
.A(n_1331),
.Y(n_1410)
);

NAND2xp5_ASAP7_75t_L g1411 ( 
.A(n_1176),
.B(n_832),
.Y(n_1411)
);

INVx1_ASAP7_75t_L g1412 ( 
.A(n_1218),
.Y(n_1412)
);

NAND2xp5_ASAP7_75t_L g1413 ( 
.A(n_1220),
.B(n_833),
.Y(n_1413)
);

HB1xp67_ASAP7_75t_L g1414 ( 
.A(n_1207),
.Y(n_1414)
);

INVx5_ASAP7_75t_L g1415 ( 
.A(n_1365),
.Y(n_1415)
);

NAND2xp5_ASAP7_75t_SL g1416 ( 
.A(n_1167),
.B(n_683),
.Y(n_1416)
);

AOI22xp33_ASAP7_75t_SL g1417 ( 
.A1(n_1268),
.A2(n_693),
.B1(n_696),
.B2(n_686),
.Y(n_1417)
);

AND2x2_ASAP7_75t_L g1418 ( 
.A(n_1200),
.B(n_834),
.Y(n_1418)
);

AOI22xp33_ASAP7_75t_L g1419 ( 
.A1(n_1333),
.A2(n_1228),
.B1(n_1235),
.B2(n_1229),
.Y(n_1419)
);

AOI22xp5_ASAP7_75t_L g1420 ( 
.A1(n_1251),
.A2(n_703),
.B1(n_704),
.B2(n_698),
.Y(n_1420)
);

NAND2xp5_ASAP7_75t_L g1421 ( 
.A(n_1222),
.B(n_706),
.Y(n_1421)
);

NAND2xp5_ASAP7_75t_L g1422 ( 
.A(n_1342),
.B(n_708),
.Y(n_1422)
);

NOR2xp33_ASAP7_75t_L g1423 ( 
.A(n_1167),
.B(n_711),
.Y(n_1423)
);

AND3x1_ASAP7_75t_L g1424 ( 
.A(n_1221),
.B(n_677),
.C(n_665),
.Y(n_1424)
);

NAND2xp5_ASAP7_75t_L g1425 ( 
.A(n_1324),
.B(n_750),
.Y(n_1425)
);

AOI22xp33_ASAP7_75t_L g1426 ( 
.A1(n_1239),
.A2(n_725),
.B1(n_732),
.B2(n_712),
.Y(n_1426)
);

INVx2_ASAP7_75t_L g1427 ( 
.A(n_1213),
.Y(n_1427)
);

INVx2_ASAP7_75t_SL g1428 ( 
.A(n_1363),
.Y(n_1428)
);

NAND2xp5_ASAP7_75t_L g1429 ( 
.A(n_1187),
.B(n_753),
.Y(n_1429)
);

NAND2xp5_ASAP7_75t_SL g1430 ( 
.A(n_1194),
.B(n_735),
.Y(n_1430)
);

NAND2xp5_ASAP7_75t_L g1431 ( 
.A(n_1187),
.B(n_1194),
.Y(n_1431)
);

INVx2_ASAP7_75t_SL g1432 ( 
.A(n_1170),
.Y(n_1432)
);

NAND2xp5_ASAP7_75t_L g1433 ( 
.A(n_1206),
.B(n_756),
.Y(n_1433)
);

AOI221xp5_ASAP7_75t_SL g1434 ( 
.A1(n_1285),
.A2(n_699),
.B1(n_700),
.B2(n_697),
.C(n_685),
.Y(n_1434)
);

INVx2_ASAP7_75t_L g1435 ( 
.A(n_1171),
.Y(n_1435)
);

INVx1_ASAP7_75t_L g1436 ( 
.A(n_1253),
.Y(n_1436)
);

NAND2xp5_ASAP7_75t_L g1437 ( 
.A(n_1285),
.B(n_702),
.Y(n_1437)
);

NAND2xp5_ASAP7_75t_L g1438 ( 
.A(n_1206),
.B(n_739),
.Y(n_1438)
);

AOI22xp5_ASAP7_75t_L g1439 ( 
.A1(n_1224),
.A2(n_742),
.B1(n_743),
.B2(n_740),
.Y(n_1439)
);

INVx2_ASAP7_75t_L g1440 ( 
.A(n_1171),
.Y(n_1440)
);

NAND2xp33_ASAP7_75t_L g1441 ( 
.A(n_1186),
.B(n_745),
.Y(n_1441)
);

NAND2x1_ASAP7_75t_L g1442 ( 
.A(n_1252),
.B(n_869),
.Y(n_1442)
);

INVx1_ASAP7_75t_L g1443 ( 
.A(n_1263),
.Y(n_1443)
);

NAND2xp5_ASAP7_75t_L g1444 ( 
.A(n_1259),
.B(n_752),
.Y(n_1444)
);

NOR2xp33_ASAP7_75t_L g1445 ( 
.A(n_1231),
.B(n_759),
.Y(n_1445)
);

AOI22xp5_ASAP7_75t_L g1446 ( 
.A1(n_1260),
.A2(n_727),
.B1(n_733),
.B2(n_726),
.Y(n_1446)
);

INVx1_ASAP7_75t_L g1447 ( 
.A(n_1264),
.Y(n_1447)
);

NAND3xp33_ASAP7_75t_L g1448 ( 
.A(n_1345),
.B(n_748),
.C(n_734),
.Y(n_1448)
);

NAND2xp5_ASAP7_75t_SL g1449 ( 
.A(n_1319),
.B(n_755),
.Y(n_1449)
);

INVx1_ASAP7_75t_L g1450 ( 
.A(n_1269),
.Y(n_1450)
);

NAND2xp5_ASAP7_75t_SL g1451 ( 
.A(n_1312),
.B(n_761),
.Y(n_1451)
);

AOI22xp33_ASAP7_75t_L g1452 ( 
.A1(n_1244),
.A2(n_741),
.B1(n_763),
.B2(n_760),
.Y(n_1452)
);

INVx2_ASAP7_75t_L g1453 ( 
.A(n_1287),
.Y(n_1453)
);

INVx1_ASAP7_75t_L g1454 ( 
.A(n_1270),
.Y(n_1454)
);

BUFx6f_ASAP7_75t_L g1455 ( 
.A(n_1296),
.Y(n_1455)
);

NAND2xp5_ASAP7_75t_SL g1456 ( 
.A(n_1267),
.B(n_540),
.Y(n_1456)
);

INVx2_ASAP7_75t_L g1457 ( 
.A(n_1295),
.Y(n_1457)
);

A2O1A1Ixp33_ASAP7_75t_L g1458 ( 
.A1(n_1323),
.A2(n_871),
.B(n_869),
.C(n_582),
.Y(n_1458)
);

NAND2xp5_ASAP7_75t_SL g1459 ( 
.A(n_1271),
.B(n_684),
.Y(n_1459)
);

NAND2xp5_ASAP7_75t_L g1460 ( 
.A(n_1274),
.B(n_871),
.Y(n_1460)
);

OAI21xp5_ASAP7_75t_L g1461 ( 
.A1(n_1304),
.A2(n_544),
.B(n_542),
.Y(n_1461)
);

BUFx3_ASAP7_75t_L g1462 ( 
.A(n_1170),
.Y(n_1462)
);

INVx2_ASAP7_75t_L g1463 ( 
.A(n_1301),
.Y(n_1463)
);

NAND2xp5_ASAP7_75t_L g1464 ( 
.A(n_1225),
.B(n_869),
.Y(n_1464)
);

NOR2xp33_ASAP7_75t_L g1465 ( 
.A(n_1248),
.B(n_545),
.Y(n_1465)
);

INVx2_ASAP7_75t_L g1466 ( 
.A(n_1245),
.Y(n_1466)
);

INVx2_ASAP7_75t_L g1467 ( 
.A(n_1223),
.Y(n_1467)
);

NAND2xp5_ASAP7_75t_SL g1468 ( 
.A(n_1252),
.B(n_715),
.Y(n_1468)
);

INVxp67_ASAP7_75t_L g1469 ( 
.A(n_1240),
.Y(n_1469)
);

O2A1O1Ixp33_ASAP7_75t_L g1470 ( 
.A1(n_1313),
.A2(n_2),
.B(n_0),
.C(n_1),
.Y(n_1470)
);

HB1xp67_ASAP7_75t_L g1471 ( 
.A(n_1200),
.Y(n_1471)
);

INVx1_ASAP7_75t_L g1472 ( 
.A(n_1225),
.Y(n_1472)
);

NAND2xp33_ASAP7_75t_L g1473 ( 
.A(n_1186),
.B(n_546),
.Y(n_1473)
);

AND2x2_ASAP7_75t_L g1474 ( 
.A(n_1236),
.B(n_869),
.Y(n_1474)
);

INVx1_ASAP7_75t_L g1475 ( 
.A(n_1280),
.Y(n_1475)
);

OAI22x1_ASAP7_75t_L g1476 ( 
.A1(n_1288),
.A2(n_552),
.B1(n_554),
.B2(n_549),
.Y(n_1476)
);

AOI22xp33_ASAP7_75t_SL g1477 ( 
.A1(n_1349),
.A2(n_601),
.B1(n_651),
.B2(n_561),
.Y(n_1477)
);

NAND2xp5_ASAP7_75t_L g1478 ( 
.A(n_1307),
.B(n_1),
.Y(n_1478)
);

INVx1_ASAP7_75t_L g1479 ( 
.A(n_1280),
.Y(n_1479)
);

NOR2xp33_ASAP7_75t_L g1480 ( 
.A(n_1262),
.B(n_1226),
.Y(n_1480)
);

NAND2xp5_ASAP7_75t_L g1481 ( 
.A(n_1307),
.B(n_2),
.Y(n_1481)
);

INVx1_ASAP7_75t_L g1482 ( 
.A(n_1350),
.Y(n_1482)
);

NAND2xp5_ASAP7_75t_L g1483 ( 
.A(n_1338),
.B(n_3),
.Y(n_1483)
);

NOR2xp33_ASAP7_75t_L g1484 ( 
.A(n_1294),
.B(n_563),
.Y(n_1484)
);

NAND2xp5_ASAP7_75t_L g1485 ( 
.A(n_1338),
.B(n_4),
.Y(n_1485)
);

INVx3_ASAP7_75t_L g1486 ( 
.A(n_1344),
.Y(n_1486)
);

NAND3xp33_ASAP7_75t_SL g1487 ( 
.A(n_1217),
.B(n_573),
.C(n_564),
.Y(n_1487)
);

NAND2xp5_ASAP7_75t_L g1488 ( 
.A(n_1291),
.B(n_6),
.Y(n_1488)
);

NAND2xp5_ASAP7_75t_L g1489 ( 
.A(n_1291),
.B(n_7),
.Y(n_1489)
);

AND2x4_ASAP7_75t_L g1490 ( 
.A(n_1310),
.B(n_869),
.Y(n_1490)
);

NAND2xp5_ASAP7_75t_SL g1491 ( 
.A(n_1265),
.B(n_1180),
.Y(n_1491)
);

INVx2_ASAP7_75t_SL g1492 ( 
.A(n_1250),
.Y(n_1492)
);

NAND2xp5_ASAP7_75t_L g1493 ( 
.A(n_1332),
.B(n_9),
.Y(n_1493)
);

INVx2_ASAP7_75t_L g1494 ( 
.A(n_1242),
.Y(n_1494)
);

NAND2xp5_ASAP7_75t_L g1495 ( 
.A(n_1265),
.B(n_1293),
.Y(n_1495)
);

NAND2xp5_ASAP7_75t_L g1496 ( 
.A(n_1335),
.B(n_9),
.Y(n_1496)
);

INVx3_ASAP7_75t_L g1497 ( 
.A(n_1344),
.Y(n_1497)
);

NAND2xp5_ASAP7_75t_L g1498 ( 
.A(n_1180),
.B(n_10),
.Y(n_1498)
);

NAND2xp5_ASAP7_75t_L g1499 ( 
.A(n_1193),
.B(n_10),
.Y(n_1499)
);

AOI22xp5_ASAP7_75t_L g1500 ( 
.A1(n_1168),
.A2(n_574),
.B1(n_581),
.B2(n_580),
.Y(n_1500)
);

NOR2xp33_ASAP7_75t_L g1501 ( 
.A(n_1273),
.B(n_1303),
.Y(n_1501)
);

NAND2xp5_ASAP7_75t_SL g1502 ( 
.A(n_1296),
.B(n_586),
.Y(n_1502)
);

AND2x4_ASAP7_75t_L g1503 ( 
.A(n_1310),
.B(n_869),
.Y(n_1503)
);

INVx1_ASAP7_75t_L g1504 ( 
.A(n_1249),
.Y(n_1504)
);

INVx2_ASAP7_75t_L g1505 ( 
.A(n_1261),
.Y(n_1505)
);

AOI22xp33_ASAP7_75t_L g1506 ( 
.A1(n_1275),
.A2(n_601),
.B1(n_651),
.B2(n_561),
.Y(n_1506)
);

A2O1A1Ixp33_ASAP7_75t_L g1507 ( 
.A1(n_1247),
.A2(n_592),
.B(n_599),
.C(n_597),
.Y(n_1507)
);

AND2x4_ASAP7_75t_L g1508 ( 
.A(n_1183),
.B(n_11),
.Y(n_1508)
);

NAND2xp5_ASAP7_75t_L g1509 ( 
.A(n_1193),
.B(n_11),
.Y(n_1509)
);

INVx1_ASAP7_75t_L g1510 ( 
.A(n_1279),
.Y(n_1510)
);

INVx1_ASAP7_75t_L g1511 ( 
.A(n_1283),
.Y(n_1511)
);

NOR2xp33_ASAP7_75t_L g1512 ( 
.A(n_1258),
.B(n_602),
.Y(n_1512)
);

AOI22xp5_ASAP7_75t_L g1513 ( 
.A1(n_1329),
.A2(n_614),
.B1(n_615),
.B2(n_612),
.Y(n_1513)
);

CKINVDCx5p33_ASAP7_75t_R g1514 ( 
.A(n_1277),
.Y(n_1514)
);

AND2x4_ASAP7_75t_L g1515 ( 
.A(n_1183),
.B(n_1284),
.Y(n_1515)
);

HB1xp67_ASAP7_75t_L g1516 ( 
.A(n_1346),
.Y(n_1516)
);

INVx1_ASAP7_75t_L g1517 ( 
.A(n_1318),
.Y(n_1517)
);

AOI22xp33_ASAP7_75t_L g1518 ( 
.A1(n_1299),
.A2(n_601),
.B1(n_651),
.B2(n_561),
.Y(n_1518)
);

BUFx3_ASAP7_75t_L g1519 ( 
.A(n_1173),
.Y(n_1519)
);

INVx3_ASAP7_75t_L g1520 ( 
.A(n_1230),
.Y(n_1520)
);

INVx2_ASAP7_75t_L g1521 ( 
.A(n_1300),
.Y(n_1521)
);

AND2x2_ASAP7_75t_L g1522 ( 
.A(n_1358),
.B(n_12),
.Y(n_1522)
);

CKINVDCx20_ASAP7_75t_R g1523 ( 
.A(n_1296),
.Y(n_1523)
);

INVx2_ASAP7_75t_SL g1524 ( 
.A(n_1173),
.Y(n_1524)
);

INVx1_ASAP7_75t_L g1525 ( 
.A(n_1309),
.Y(n_1525)
);

INVx1_ASAP7_75t_L g1526 ( 
.A(n_1311),
.Y(n_1526)
);

INVx1_ASAP7_75t_L g1527 ( 
.A(n_1314),
.Y(n_1527)
);

BUFx4f_ASAP7_75t_L g1528 ( 
.A(n_1365),
.Y(n_1528)
);

INVx1_ASAP7_75t_L g1529 ( 
.A(n_1315),
.Y(n_1529)
);

AOI22xp33_ASAP7_75t_L g1530 ( 
.A1(n_1320),
.A2(n_601),
.B1(n_651),
.B2(n_561),
.Y(n_1530)
);

AOI22xp5_ASAP7_75t_SL g1531 ( 
.A1(n_1243),
.A2(n_754),
.B1(n_618),
.B2(n_624),
.Y(n_1531)
);

AND2x2_ASAP7_75t_L g1532 ( 
.A(n_1358),
.B(n_12),
.Y(n_1532)
);

AOI21xp5_ASAP7_75t_L g1533 ( 
.A1(n_1201),
.A2(n_630),
.B(n_616),
.Y(n_1533)
);

INVx1_ASAP7_75t_L g1534 ( 
.A(n_1325),
.Y(n_1534)
);

AND2x2_ASAP7_75t_L g1535 ( 
.A(n_1284),
.B(n_13),
.Y(n_1535)
);

NAND2xp5_ASAP7_75t_L g1536 ( 
.A(n_1202),
.B(n_13),
.Y(n_1536)
);

NAND2xp5_ASAP7_75t_L g1537 ( 
.A(n_1202),
.B(n_14),
.Y(n_1537)
);

NAND3xp33_ASAP7_75t_SL g1538 ( 
.A(n_1233),
.B(n_1185),
.C(n_1355),
.Y(n_1538)
);

INVx1_ASAP7_75t_L g1539 ( 
.A(n_1326),
.Y(n_1539)
);

INVx2_ASAP7_75t_SL g1540 ( 
.A(n_1173),
.Y(n_1540)
);

INVx1_ASAP7_75t_L g1541 ( 
.A(n_1328),
.Y(n_1541)
);

INVx2_ASAP7_75t_L g1542 ( 
.A(n_1321),
.Y(n_1542)
);

O2A1O1Ixp5_ASAP7_75t_L g1543 ( 
.A1(n_1181),
.A2(n_17),
.B(n_15),
.C(n_16),
.Y(n_1543)
);

HB1xp67_ASAP7_75t_L g1544 ( 
.A(n_1178),
.Y(n_1544)
);

NAND2xp5_ASAP7_75t_L g1545 ( 
.A(n_1243),
.B(n_15),
.Y(n_1545)
);

HB1xp67_ASAP7_75t_L g1546 ( 
.A(n_1178),
.Y(n_1546)
);

AND2x6_ASAP7_75t_SL g1547 ( 
.A(n_1290),
.B(n_16),
.Y(n_1547)
);

INVx1_ASAP7_75t_L g1548 ( 
.A(n_1330),
.Y(n_1548)
);

NAND2xp5_ASAP7_75t_L g1549 ( 
.A(n_1243),
.B(n_17),
.Y(n_1549)
);

INVx1_ASAP7_75t_L g1550 ( 
.A(n_1322),
.Y(n_1550)
);

NAND2xp5_ASAP7_75t_L g1551 ( 
.A(n_1243),
.B(n_18),
.Y(n_1551)
);

NAND2xp5_ASAP7_75t_SL g1552 ( 
.A(n_1178),
.B(n_631),
.Y(n_1552)
);

NAND2xp5_ASAP7_75t_SL g1553 ( 
.A(n_1281),
.B(n_751),
.Y(n_1553)
);

INVx2_ASAP7_75t_L g1554 ( 
.A(n_1163),
.Y(n_1554)
);

AO22x1_ASAP7_75t_L g1555 ( 
.A1(n_1365),
.A2(n_633),
.B1(n_637),
.B2(n_632),
.Y(n_1555)
);

NAND2xp5_ASAP7_75t_L g1556 ( 
.A(n_1281),
.B(n_18),
.Y(n_1556)
);

INVx1_ASAP7_75t_L g1557 ( 
.A(n_1334),
.Y(n_1557)
);

INVx1_ASAP7_75t_L g1558 ( 
.A(n_1337),
.Y(n_1558)
);

NAND2xp5_ASAP7_75t_SL g1559 ( 
.A(n_1230),
.B(n_1272),
.Y(n_1559)
);

INVx1_ASAP7_75t_L g1560 ( 
.A(n_1177),
.Y(n_1560)
);

NAND2xp5_ASAP7_75t_L g1561 ( 
.A(n_1361),
.B(n_19),
.Y(n_1561)
);

INVx2_ASAP7_75t_L g1562 ( 
.A(n_1364),
.Y(n_1562)
);

INVx2_ASAP7_75t_L g1563 ( 
.A(n_1340),
.Y(n_1563)
);

INVx1_ASAP7_75t_L g1564 ( 
.A(n_1292),
.Y(n_1564)
);

OAI22xp33_ASAP7_75t_L g1565 ( 
.A1(n_1360),
.A2(n_655),
.B1(n_657),
.B2(n_653),
.Y(n_1565)
);

O2A1O1Ixp33_ASAP7_75t_L g1566 ( 
.A1(n_1192),
.A2(n_23),
.B(n_19),
.C(n_21),
.Y(n_1566)
);

INVx1_ASAP7_75t_L g1567 ( 
.A(n_1266),
.Y(n_1567)
);

BUFx6f_ASAP7_75t_L g1568 ( 
.A(n_1230),
.Y(n_1568)
);

NAND2x1p5_ASAP7_75t_L g1569 ( 
.A(n_1208),
.B(n_724),
.Y(n_1569)
);

BUFx12f_ASAP7_75t_L g1570 ( 
.A(n_1272),
.Y(n_1570)
);

NAND2xp5_ASAP7_75t_L g1571 ( 
.A(n_1329),
.B(n_24),
.Y(n_1571)
);

NAND2xp5_ASAP7_75t_L g1572 ( 
.A(n_1329),
.B(n_25),
.Y(n_1572)
);

BUFx3_ASAP7_75t_L g1573 ( 
.A(n_1208),
.Y(n_1573)
);

BUFx6f_ASAP7_75t_L g1574 ( 
.A(n_1272),
.Y(n_1574)
);

NAND2xp5_ASAP7_75t_L g1575 ( 
.A(n_1329),
.B(n_1186),
.Y(n_1575)
);

INVx1_ASAP7_75t_L g1576 ( 
.A(n_1339),
.Y(n_1576)
);

INVx5_ASAP7_75t_L g1577 ( 
.A(n_1455),
.Y(n_1577)
);

NOR2x1_ASAP7_75t_L g1578 ( 
.A(n_1523),
.B(n_1354),
.Y(n_1578)
);

INVx1_ASAP7_75t_L g1579 ( 
.A(n_1401),
.Y(n_1579)
);

INVx1_ASAP7_75t_L g1580 ( 
.A(n_1404),
.Y(n_1580)
);

INVx1_ASAP7_75t_L g1581 ( 
.A(n_1371),
.Y(n_1581)
);

BUFx6f_ASAP7_75t_L g1582 ( 
.A(n_1455),
.Y(n_1582)
);

NAND3xp33_ASAP7_75t_SL g1583 ( 
.A(n_1368),
.B(n_678),
.C(n_676),
.Y(n_1583)
);

INVx1_ASAP7_75t_L g1584 ( 
.A(n_1389),
.Y(n_1584)
);

AND2x4_ASAP7_75t_L g1585 ( 
.A(n_1515),
.B(n_1290),
.Y(n_1585)
);

INVx2_ASAP7_75t_L g1586 ( 
.A(n_1466),
.Y(n_1586)
);

AND2x2_ASAP7_75t_L g1587 ( 
.A(n_1418),
.B(n_1390),
.Y(n_1587)
);

NAND2xp5_ASAP7_75t_SL g1588 ( 
.A(n_1531),
.B(n_1282),
.Y(n_1588)
);

NAND2xp5_ASAP7_75t_L g1589 ( 
.A(n_1482),
.B(n_1354),
.Y(n_1589)
);

NAND2xp5_ASAP7_75t_SL g1590 ( 
.A(n_1531),
.B(n_1282),
.Y(n_1590)
);

HB1xp67_ASAP7_75t_L g1591 ( 
.A(n_1380),
.Y(n_1591)
);

INVx2_ASAP7_75t_L g1592 ( 
.A(n_1453),
.Y(n_1592)
);

OR2x4_ASAP7_75t_L g1593 ( 
.A(n_1480),
.B(n_1341),
.Y(n_1593)
);

INVxp67_ASAP7_75t_L g1594 ( 
.A(n_1414),
.Y(n_1594)
);

INVx1_ASAP7_75t_L g1595 ( 
.A(n_1409),
.Y(n_1595)
);

AOI22xp33_ASAP7_75t_L g1596 ( 
.A1(n_1417),
.A2(n_1289),
.B1(n_1184),
.B2(n_1359),
.Y(n_1596)
);

INVx1_ASAP7_75t_L g1597 ( 
.A(n_1412),
.Y(n_1597)
);

NOR3xp33_ASAP7_75t_SL g1598 ( 
.A(n_1370),
.B(n_1343),
.C(n_1327),
.Y(n_1598)
);

INVx3_ASAP7_75t_L g1599 ( 
.A(n_1455),
.Y(n_1599)
);

NOR2xp33_ASAP7_75t_R g1600 ( 
.A(n_1514),
.B(n_1282),
.Y(n_1600)
);

NOR2xp33_ASAP7_75t_L g1601 ( 
.A(n_1445),
.B(n_1356),
.Y(n_1601)
);

INVx2_ASAP7_75t_L g1602 ( 
.A(n_1369),
.Y(n_1602)
);

INVx2_ASAP7_75t_L g1603 ( 
.A(n_1372),
.Y(n_1603)
);

NAND2xp5_ASAP7_75t_SL g1604 ( 
.A(n_1388),
.B(n_1305),
.Y(n_1604)
);

NOR2xp33_ASAP7_75t_L g1605 ( 
.A(n_1469),
.B(n_1348),
.Y(n_1605)
);

BUFx2_ASAP7_75t_L g1606 ( 
.A(n_1570),
.Y(n_1606)
);

INVx1_ASAP7_75t_L g1607 ( 
.A(n_1436),
.Y(n_1607)
);

INVx3_ASAP7_75t_L g1608 ( 
.A(n_1568),
.Y(n_1608)
);

NAND2xp5_ASAP7_75t_L g1609 ( 
.A(n_1399),
.B(n_1184),
.Y(n_1609)
);

INVx1_ASAP7_75t_L g1610 ( 
.A(n_1443),
.Y(n_1610)
);

INVx2_ASAP7_75t_L g1611 ( 
.A(n_1403),
.Y(n_1611)
);

INVx1_ASAP7_75t_L g1612 ( 
.A(n_1447),
.Y(n_1612)
);

AOI21xp5_ASAP7_75t_L g1613 ( 
.A1(n_1473),
.A2(n_1181),
.B(n_1357),
.Y(n_1613)
);

AND2x4_ASAP7_75t_L g1614 ( 
.A(n_1515),
.B(n_1305),
.Y(n_1614)
);

BUFx4f_ASAP7_75t_L g1615 ( 
.A(n_1406),
.Y(n_1615)
);

NAND2x1p5_ASAP7_75t_L g1616 ( 
.A(n_1410),
.B(n_1305),
.Y(n_1616)
);

NAND2xp5_ASAP7_75t_L g1617 ( 
.A(n_1383),
.B(n_1184),
.Y(n_1617)
);

NAND2xp5_ASAP7_75t_L g1618 ( 
.A(n_1402),
.B(n_1184),
.Y(n_1618)
);

NAND2xp5_ASAP7_75t_L g1619 ( 
.A(n_1405),
.B(n_1352),
.Y(n_1619)
);

AND2x2_ASAP7_75t_L g1620 ( 
.A(n_1471),
.B(n_1196),
.Y(n_1620)
);

OR2x6_ASAP7_75t_L g1621 ( 
.A(n_1428),
.B(n_1302),
.Y(n_1621)
);

INVx1_ASAP7_75t_L g1622 ( 
.A(n_1450),
.Y(n_1622)
);

AND2x2_ASAP7_75t_L g1623 ( 
.A(n_1508),
.B(n_1210),
.Y(n_1623)
);

BUFx6f_ASAP7_75t_L g1624 ( 
.A(n_1410),
.Y(n_1624)
);

INVx1_ASAP7_75t_L g1625 ( 
.A(n_1454),
.Y(n_1625)
);

HB1xp67_ASAP7_75t_L g1626 ( 
.A(n_1516),
.Y(n_1626)
);

INVxp67_ASAP7_75t_L g1627 ( 
.A(n_1501),
.Y(n_1627)
);

AND2x4_ASAP7_75t_L g1628 ( 
.A(n_1395),
.B(n_1186),
.Y(n_1628)
);

OR2x2_ASAP7_75t_L g1629 ( 
.A(n_1411),
.B(n_1336),
.Y(n_1629)
);

INVx1_ASAP7_75t_SL g1630 ( 
.A(n_1396),
.Y(n_1630)
);

NOR3xp33_ASAP7_75t_SL g1631 ( 
.A(n_1487),
.B(n_1392),
.C(n_1366),
.Y(n_1631)
);

AND2x4_ASAP7_75t_L g1632 ( 
.A(n_1395),
.B(n_1347),
.Y(n_1632)
);

CKINVDCx5p33_ASAP7_75t_R g1633 ( 
.A(n_1462),
.Y(n_1633)
);

AND2x2_ASAP7_75t_L g1634 ( 
.A(n_1508),
.B(n_25),
.Y(n_1634)
);

NOR2xp67_ASAP7_75t_L g1635 ( 
.A(n_1432),
.B(n_1257),
.Y(n_1635)
);

BUFx2_ASAP7_75t_SL g1636 ( 
.A(n_1410),
.Y(n_1636)
);

BUFx6f_ASAP7_75t_L g1637 ( 
.A(n_1568),
.Y(n_1637)
);

INVx3_ASAP7_75t_L g1638 ( 
.A(n_1519),
.Y(n_1638)
);

BUFx2_ASAP7_75t_L g1639 ( 
.A(n_1396),
.Y(n_1639)
);

INVx1_ASAP7_75t_L g1640 ( 
.A(n_1457),
.Y(n_1640)
);

AND2x4_ASAP7_75t_L g1641 ( 
.A(n_1491),
.B(n_1357),
.Y(n_1641)
);

AOI21xp5_ASAP7_75t_L g1642 ( 
.A1(n_1367),
.A2(n_1316),
.B(n_1278),
.Y(n_1642)
);

AND2x4_ASAP7_75t_L g1643 ( 
.A(n_1486),
.B(n_1351),
.Y(n_1643)
);

NOR2xp33_ASAP7_75t_R g1644 ( 
.A(n_1375),
.B(n_681),
.Y(n_1644)
);

INVx2_ASAP7_75t_L g1645 ( 
.A(n_1407),
.Y(n_1645)
);

CKINVDCx5p33_ASAP7_75t_R g1646 ( 
.A(n_1547),
.Y(n_1646)
);

INVx1_ASAP7_75t_L g1647 ( 
.A(n_1463),
.Y(n_1647)
);

INVx4_ASAP7_75t_L g1648 ( 
.A(n_1568),
.Y(n_1648)
);

AND2x4_ASAP7_75t_L g1649 ( 
.A(n_1486),
.B(n_1256),
.Y(n_1649)
);

NAND2xp5_ASAP7_75t_L g1650 ( 
.A(n_1384),
.B(n_1237),
.Y(n_1650)
);

O2A1O1Ixp5_ASAP7_75t_L g1651 ( 
.A1(n_1496),
.A2(n_1216),
.B(n_28),
.C(n_26),
.Y(n_1651)
);

HB1xp67_ASAP7_75t_L g1652 ( 
.A(n_1556),
.Y(n_1652)
);

INVx3_ASAP7_75t_L g1653 ( 
.A(n_1573),
.Y(n_1653)
);

BUFx3_ASAP7_75t_L g1654 ( 
.A(n_1492),
.Y(n_1654)
);

CKINVDCx5p33_ASAP7_75t_R g1655 ( 
.A(n_1547),
.Y(n_1655)
);

AOI22xp33_ASAP7_75t_L g1656 ( 
.A1(n_1448),
.A2(n_724),
.B1(n_692),
.B2(n_714),
.Y(n_1656)
);

INVx4_ASAP7_75t_L g1657 ( 
.A(n_1574),
.Y(n_1657)
);

AND2x6_ASAP7_75t_L g1658 ( 
.A(n_1522),
.B(n_724),
.Y(n_1658)
);

BUFx3_ASAP7_75t_L g1659 ( 
.A(n_1574),
.Y(n_1659)
);

AND2x4_ASAP7_75t_L g1660 ( 
.A(n_1497),
.B(n_290),
.Y(n_1660)
);

AND2x2_ASAP7_75t_L g1661 ( 
.A(n_1535),
.B(n_26),
.Y(n_1661)
);

NOR3xp33_ASAP7_75t_SL g1662 ( 
.A(n_1416),
.B(n_747),
.C(n_716),
.Y(n_1662)
);

INVx1_ASAP7_75t_L g1663 ( 
.A(n_1548),
.Y(n_1663)
);

NAND2x1p5_ASAP7_75t_L g1664 ( 
.A(n_1497),
.B(n_724),
.Y(n_1664)
);

OR2x2_ASAP7_75t_L g1665 ( 
.A(n_1425),
.B(n_27),
.Y(n_1665)
);

BUFx2_ASAP7_75t_L g1666 ( 
.A(n_1544),
.Y(n_1666)
);

INVx1_ASAP7_75t_L g1667 ( 
.A(n_1534),
.Y(n_1667)
);

NAND2xp5_ASAP7_75t_L g1668 ( 
.A(n_1484),
.B(n_27),
.Y(n_1668)
);

NAND2xp5_ASAP7_75t_SL g1669 ( 
.A(n_1388),
.B(n_746),
.Y(n_1669)
);

INVx1_ASAP7_75t_L g1670 ( 
.A(n_1539),
.Y(n_1670)
);

AOI22xp5_ASAP7_75t_L g1671 ( 
.A1(n_1448),
.A2(n_718),
.B1(n_730),
.B2(n_688),
.Y(n_1671)
);

NAND2xp5_ASAP7_75t_L g1672 ( 
.A(n_1422),
.B(n_28),
.Y(n_1672)
);

AND2x4_ASAP7_75t_L g1673 ( 
.A(n_1431),
.B(n_291),
.Y(n_1673)
);

NOR3xp33_ASAP7_75t_SL g1674 ( 
.A(n_1430),
.B(n_29),
.C(n_30),
.Y(n_1674)
);

AOI22xp5_ASAP7_75t_L g1675 ( 
.A1(n_1423),
.A2(n_31),
.B1(n_29),
.B2(n_30),
.Y(n_1675)
);

NAND2xp5_ASAP7_75t_L g1676 ( 
.A(n_1435),
.B(n_31),
.Y(n_1676)
);

INVx1_ASAP7_75t_L g1677 ( 
.A(n_1541),
.Y(n_1677)
);

NAND2xp5_ASAP7_75t_SL g1678 ( 
.A(n_1378),
.B(n_1415),
.Y(n_1678)
);

INVx2_ASAP7_75t_L g1679 ( 
.A(n_1427),
.Y(n_1679)
);

NOR2xp33_ASAP7_75t_R g1680 ( 
.A(n_1528),
.B(n_292),
.Y(n_1680)
);

INVx1_ASAP7_75t_L g1681 ( 
.A(n_1517),
.Y(n_1681)
);

INVx3_ASAP7_75t_L g1682 ( 
.A(n_1574),
.Y(n_1682)
);

CKINVDCx11_ASAP7_75t_R g1683 ( 
.A(n_1554),
.Y(n_1683)
);

NOR2x2_ASAP7_75t_L g1684 ( 
.A(n_1440),
.B(n_32),
.Y(n_1684)
);

CKINVDCx5p33_ASAP7_75t_R g1685 ( 
.A(n_1546),
.Y(n_1685)
);

NOR2xp33_ASAP7_75t_R g1686 ( 
.A(n_1528),
.B(n_294),
.Y(n_1686)
);

INVx2_ASAP7_75t_L g1687 ( 
.A(n_1467),
.Y(n_1687)
);

INVx2_ASAP7_75t_L g1688 ( 
.A(n_1494),
.Y(n_1688)
);

INVx1_ASAP7_75t_L g1689 ( 
.A(n_1472),
.Y(n_1689)
);

BUFx3_ASAP7_75t_L g1690 ( 
.A(n_1524),
.Y(n_1690)
);

INVxp67_ASAP7_75t_L g1691 ( 
.A(n_1512),
.Y(n_1691)
);

INVx1_ASAP7_75t_L g1692 ( 
.A(n_1475),
.Y(n_1692)
);

NAND2xp5_ASAP7_75t_SL g1693 ( 
.A(n_1378),
.B(n_33),
.Y(n_1693)
);

INVx2_ASAP7_75t_L g1694 ( 
.A(n_1505),
.Y(n_1694)
);

NAND2xp33_ASAP7_75t_L g1695 ( 
.A(n_1378),
.B(n_33),
.Y(n_1695)
);

INVx4_ASAP7_75t_L g1696 ( 
.A(n_1415),
.Y(n_1696)
);

NOR3xp33_ASAP7_75t_SL g1697 ( 
.A(n_1499),
.B(n_34),
.C(n_35),
.Y(n_1697)
);

INVx5_ASAP7_75t_L g1698 ( 
.A(n_1415),
.Y(n_1698)
);

INVx1_ASAP7_75t_L g1699 ( 
.A(n_1479),
.Y(n_1699)
);

INVx1_ASAP7_75t_L g1700 ( 
.A(n_1550),
.Y(n_1700)
);

CKINVDCx5p33_ASAP7_75t_R g1701 ( 
.A(n_1540),
.Y(n_1701)
);

INVx1_ASAP7_75t_L g1702 ( 
.A(n_1557),
.Y(n_1702)
);

INVx3_ASAP7_75t_SL g1703 ( 
.A(n_1394),
.Y(n_1703)
);

CKINVDCx14_ASAP7_75t_R g1704 ( 
.A(n_1465),
.Y(n_1704)
);

INVx2_ASAP7_75t_L g1705 ( 
.A(n_1521),
.Y(n_1705)
);

AND2x4_ASAP7_75t_L g1706 ( 
.A(n_1495),
.B(n_536),
.Y(n_1706)
);

BUFx3_ASAP7_75t_L g1707 ( 
.A(n_1520),
.Y(n_1707)
);

NAND2xp5_ASAP7_75t_L g1708 ( 
.A(n_1385),
.B(n_34),
.Y(n_1708)
);

INVx4_ASAP7_75t_L g1709 ( 
.A(n_1520),
.Y(n_1709)
);

AND2x4_ASAP7_75t_L g1710 ( 
.A(n_1490),
.B(n_534),
.Y(n_1710)
);

AOI22xp33_ASAP7_75t_L g1711 ( 
.A1(n_1532),
.A2(n_38),
.B1(n_36),
.B2(n_37),
.Y(n_1711)
);

CKINVDCx5p33_ASAP7_75t_R g1712 ( 
.A(n_1449),
.Y(n_1712)
);

NAND2xp5_ASAP7_75t_SL g1713 ( 
.A(n_1424),
.B(n_36),
.Y(n_1713)
);

INVx3_ASAP7_75t_L g1714 ( 
.A(n_1490),
.Y(n_1714)
);

INVx2_ASAP7_75t_SL g1715 ( 
.A(n_1474),
.Y(n_1715)
);

NAND2xp5_ASAP7_75t_SL g1716 ( 
.A(n_1424),
.B(n_37),
.Y(n_1716)
);

BUFx12f_ASAP7_75t_L g1717 ( 
.A(n_1503),
.Y(n_1717)
);

NAND2xp5_ASAP7_75t_L g1718 ( 
.A(n_1386),
.B(n_38),
.Y(n_1718)
);

INVx1_ASAP7_75t_L g1719 ( 
.A(n_1558),
.Y(n_1719)
);

BUFx2_ASAP7_75t_L g1720 ( 
.A(n_1478),
.Y(n_1720)
);

CKINVDCx5p33_ASAP7_75t_R g1721 ( 
.A(n_1476),
.Y(n_1721)
);

NAND2xp5_ASAP7_75t_L g1722 ( 
.A(n_1391),
.B(n_39),
.Y(n_1722)
);

NOR2xp33_ASAP7_75t_L g1723 ( 
.A(n_1433),
.B(n_40),
.Y(n_1723)
);

INVx1_ASAP7_75t_L g1724 ( 
.A(n_1504),
.Y(n_1724)
);

BUFx6f_ASAP7_75t_L g1725 ( 
.A(n_1503),
.Y(n_1725)
);

BUFx6f_ASAP7_75t_L g1726 ( 
.A(n_1559),
.Y(n_1726)
);

NAND2xp5_ASAP7_75t_L g1727 ( 
.A(n_1393),
.B(n_41),
.Y(n_1727)
);

INVx2_ASAP7_75t_L g1728 ( 
.A(n_1510),
.Y(n_1728)
);

CKINVDCx5p33_ASAP7_75t_R g1729 ( 
.A(n_1451),
.Y(n_1729)
);

NAND2xp5_ASAP7_75t_L g1730 ( 
.A(n_1397),
.B(n_41),
.Y(n_1730)
);

HB1xp67_ASAP7_75t_L g1731 ( 
.A(n_1488),
.Y(n_1731)
);

BUFx2_ASAP7_75t_L g1732 ( 
.A(n_1481),
.Y(n_1732)
);

BUFx6f_ASAP7_75t_L g1733 ( 
.A(n_1569),
.Y(n_1733)
);

BUFx2_ASAP7_75t_L g1734 ( 
.A(n_1483),
.Y(n_1734)
);

INVx5_ASAP7_75t_L g1735 ( 
.A(n_1563),
.Y(n_1735)
);

BUFx2_ASAP7_75t_L g1736 ( 
.A(n_1485),
.Y(n_1736)
);

BUFx3_ASAP7_75t_L g1737 ( 
.A(n_1542),
.Y(n_1737)
);

AND2x4_ASAP7_75t_L g1738 ( 
.A(n_1562),
.B(n_295),
.Y(n_1738)
);

BUFx6f_ASAP7_75t_L g1739 ( 
.A(n_1569),
.Y(n_1739)
);

INVx2_ASAP7_75t_L g1740 ( 
.A(n_1511),
.Y(n_1740)
);

INVx1_ASAP7_75t_L g1741 ( 
.A(n_1525),
.Y(n_1741)
);

HB1xp67_ASAP7_75t_L g1742 ( 
.A(n_1489),
.Y(n_1742)
);

INVx1_ASAP7_75t_L g1743 ( 
.A(n_1526),
.Y(n_1743)
);

NAND2xp5_ASAP7_75t_L g1744 ( 
.A(n_1398),
.B(n_42),
.Y(n_1744)
);

AND2x2_ASAP7_75t_L g1745 ( 
.A(n_1408),
.B(n_42),
.Y(n_1745)
);

INVx1_ASAP7_75t_L g1746 ( 
.A(n_1527),
.Y(n_1746)
);

CKINVDCx8_ASAP7_75t_R g1747 ( 
.A(n_1377),
.Y(n_1747)
);

NAND2xp5_ASAP7_75t_L g1748 ( 
.A(n_1413),
.B(n_43),
.Y(n_1748)
);

BUFx2_ASAP7_75t_L g1749 ( 
.A(n_1498),
.Y(n_1749)
);

NAND2xp5_ASAP7_75t_SL g1750 ( 
.A(n_1575),
.B(n_44),
.Y(n_1750)
);

NOR2xp33_ASAP7_75t_L g1751 ( 
.A(n_1438),
.B(n_44),
.Y(n_1751)
);

HB1xp67_ASAP7_75t_L g1752 ( 
.A(n_1560),
.Y(n_1752)
);

INVx1_ASAP7_75t_L g1753 ( 
.A(n_1529),
.Y(n_1753)
);

INVx2_ASAP7_75t_L g1754 ( 
.A(n_1576),
.Y(n_1754)
);

BUFx3_ASAP7_75t_L g1755 ( 
.A(n_1429),
.Y(n_1755)
);

INVx5_ASAP7_75t_L g1756 ( 
.A(n_1441),
.Y(n_1756)
);

AOI21xp33_ASAP7_75t_L g1757 ( 
.A1(n_1461),
.A2(n_45),
.B(n_46),
.Y(n_1757)
);

NAND2x1p5_ASAP7_75t_L g1758 ( 
.A(n_1502),
.B(n_296),
.Y(n_1758)
);

INVx2_ASAP7_75t_L g1759 ( 
.A(n_1561),
.Y(n_1759)
);

INVx1_ASAP7_75t_L g1760 ( 
.A(n_1561),
.Y(n_1760)
);

A2O1A1Ixp33_ASAP7_75t_L g1761 ( 
.A1(n_1387),
.A2(n_47),
.B(n_45),
.C(n_46),
.Y(n_1761)
);

AND2x4_ASAP7_75t_L g1762 ( 
.A(n_1419),
.B(n_532),
.Y(n_1762)
);

BUFx6f_ASAP7_75t_L g1763 ( 
.A(n_1442),
.Y(n_1763)
);

NAND2xp5_ASAP7_75t_L g1764 ( 
.A(n_1493),
.B(n_47),
.Y(n_1764)
);

INVx5_ASAP7_75t_L g1765 ( 
.A(n_1555),
.Y(n_1765)
);

NAND2xp5_ASAP7_75t_L g1766 ( 
.A(n_1437),
.B(n_48),
.Y(n_1766)
);

AND2x4_ASAP7_75t_L g1767 ( 
.A(n_1553),
.B(n_528),
.Y(n_1767)
);

NAND2xp5_ASAP7_75t_L g1768 ( 
.A(n_1437),
.B(n_48),
.Y(n_1768)
);

INVx2_ASAP7_75t_SL g1769 ( 
.A(n_1509),
.Y(n_1769)
);

INVx1_ASAP7_75t_L g1770 ( 
.A(n_1460),
.Y(n_1770)
);

NAND2xp5_ASAP7_75t_SL g1771 ( 
.A(n_1477),
.B(n_1545),
.Y(n_1771)
);

NAND2xp5_ASAP7_75t_L g1772 ( 
.A(n_1400),
.B(n_49),
.Y(n_1772)
);

NOR2xp33_ASAP7_75t_L g1773 ( 
.A(n_1444),
.B(n_50),
.Y(n_1773)
);

OAI21x1_ASAP7_75t_L g1774 ( 
.A1(n_1613),
.A2(n_1464),
.B(n_1376),
.Y(n_1774)
);

NAND2xp5_ASAP7_75t_L g1775 ( 
.A(n_1587),
.B(n_1536),
.Y(n_1775)
);

OA22x2_ASAP7_75t_L g1776 ( 
.A1(n_1630),
.A2(n_1446),
.B1(n_1420),
.B2(n_1513),
.Y(n_1776)
);

INVx2_ASAP7_75t_SL g1777 ( 
.A(n_1615),
.Y(n_1777)
);

AOI21x1_ASAP7_75t_L g1778 ( 
.A1(n_1771),
.A2(n_1376),
.B(n_1373),
.Y(n_1778)
);

AND3x4_ASAP7_75t_L g1779 ( 
.A(n_1631),
.B(n_1439),
.C(n_1426),
.Y(n_1779)
);

AOI21xp5_ASAP7_75t_L g1780 ( 
.A1(n_1695),
.A2(n_1564),
.B(n_1461),
.Y(n_1780)
);

OAI21x1_ASAP7_75t_L g1781 ( 
.A1(n_1642),
.A2(n_1464),
.B(n_1381),
.Y(n_1781)
);

INVx4_ASAP7_75t_L g1782 ( 
.A(n_1633),
.Y(n_1782)
);

AND2x2_ASAP7_75t_L g1783 ( 
.A(n_1634),
.B(n_1421),
.Y(n_1783)
);

AOI21x1_ASAP7_75t_L g1784 ( 
.A1(n_1588),
.A2(n_1381),
.B(n_1379),
.Y(n_1784)
);

BUFx3_ASAP7_75t_L g1785 ( 
.A(n_1683),
.Y(n_1785)
);

OAI21x1_ASAP7_75t_L g1786 ( 
.A1(n_1770),
.A2(n_1379),
.B(n_1567),
.Y(n_1786)
);

NAND2xp5_ASAP7_75t_SL g1787 ( 
.A(n_1765),
.B(n_1549),
.Y(n_1787)
);

AND2x4_ASAP7_75t_L g1788 ( 
.A(n_1585),
.B(n_1551),
.Y(n_1788)
);

OAI21x1_ASAP7_75t_L g1789 ( 
.A1(n_1759),
.A2(n_1460),
.B(n_1543),
.Y(n_1789)
);

AO31x2_ASAP7_75t_L g1790 ( 
.A1(n_1760),
.A2(n_1458),
.A3(n_1692),
.B(n_1689),
.Y(n_1790)
);

A2O1A1Ixp33_ASAP7_75t_L g1791 ( 
.A1(n_1762),
.A2(n_1470),
.B(n_1382),
.C(n_1566),
.Y(n_1791)
);

NAND2xp5_ASAP7_75t_L g1792 ( 
.A(n_1591),
.B(n_1537),
.Y(n_1792)
);

AOI21xp5_ASAP7_75t_SL g1793 ( 
.A1(n_1762),
.A2(n_1572),
.B(n_1571),
.Y(n_1793)
);

OAI21xp5_ASAP7_75t_L g1794 ( 
.A1(n_1757),
.A2(n_1434),
.B(n_1507),
.Y(n_1794)
);

OR2x2_ASAP7_75t_L g1795 ( 
.A(n_1626),
.B(n_1374),
.Y(n_1795)
);

NOR2xp33_ASAP7_75t_L g1796 ( 
.A(n_1627),
.B(n_1552),
.Y(n_1796)
);

NAND2xp5_ASAP7_75t_L g1797 ( 
.A(n_1601),
.B(n_1434),
.Y(n_1797)
);

AOI21x1_ASAP7_75t_L g1798 ( 
.A1(n_1590),
.A2(n_1533),
.B(n_1468),
.Y(n_1798)
);

NAND2xp5_ASAP7_75t_L g1799 ( 
.A(n_1720),
.B(n_1452),
.Y(n_1799)
);

A2O1A1Ixp33_ASAP7_75t_L g1800 ( 
.A1(n_1773),
.A2(n_1500),
.B(n_1459),
.C(n_1456),
.Y(n_1800)
);

OAI21xp5_ASAP7_75t_L g1801 ( 
.A1(n_1668),
.A2(n_1565),
.B(n_1538),
.Y(n_1801)
);

INVx2_ASAP7_75t_SL g1802 ( 
.A(n_1600),
.Y(n_1802)
);

OAI21xp5_ASAP7_75t_L g1803 ( 
.A1(n_1672),
.A2(n_1518),
.B(n_1506),
.Y(n_1803)
);

INVx1_ASAP7_75t_L g1804 ( 
.A(n_1699),
.Y(n_1804)
);

O2A1O1Ixp5_ASAP7_75t_L g1805 ( 
.A1(n_1604),
.A2(n_1530),
.B(n_52),
.C(n_50),
.Y(n_1805)
);

AOI21xp5_ASAP7_75t_L g1806 ( 
.A1(n_1756),
.A2(n_1768),
.B(n_1766),
.Y(n_1806)
);

NOR2xp33_ASAP7_75t_L g1807 ( 
.A(n_1704),
.B(n_51),
.Y(n_1807)
);

NAND2xp5_ASAP7_75t_L g1808 ( 
.A(n_1732),
.B(n_51),
.Y(n_1808)
);

AND2x4_ASAP7_75t_L g1809 ( 
.A(n_1585),
.B(n_52),
.Y(n_1809)
);

INVx1_ASAP7_75t_L g1810 ( 
.A(n_1581),
.Y(n_1810)
);

OAI21xp5_ASAP7_75t_L g1811 ( 
.A1(n_1761),
.A2(n_53),
.B(n_54),
.Y(n_1811)
);

OAI21x1_ASAP7_75t_L g1812 ( 
.A1(n_1651),
.A2(n_300),
.B(n_299),
.Y(n_1812)
);

A2O1A1Ixp33_ASAP7_75t_L g1813 ( 
.A1(n_1723),
.A2(n_56),
.B(n_54),
.C(n_55),
.Y(n_1813)
);

INVx1_ASAP7_75t_SL g1814 ( 
.A(n_1685),
.Y(n_1814)
);

NAND2x1p5_ASAP7_75t_L g1815 ( 
.A(n_1698),
.B(n_301),
.Y(n_1815)
);

NOR2x1_ASAP7_75t_L g1816 ( 
.A(n_1635),
.B(n_55),
.Y(n_1816)
);

NAND2xp5_ASAP7_75t_L g1817 ( 
.A(n_1734),
.B(n_56),
.Y(n_1817)
);

NAND2xp5_ASAP7_75t_L g1818 ( 
.A(n_1736),
.B(n_57),
.Y(n_1818)
);

OAI21xp5_ASAP7_75t_L g1819 ( 
.A1(n_1751),
.A2(n_1764),
.B(n_1675),
.Y(n_1819)
);

A2O1A1Ixp33_ASAP7_75t_L g1820 ( 
.A1(n_1767),
.A2(n_60),
.B(n_58),
.C(n_59),
.Y(n_1820)
);

BUFx2_ASAP7_75t_L g1821 ( 
.A(n_1593),
.Y(n_1821)
);

OAI21xp5_ASAP7_75t_L g1822 ( 
.A1(n_1583),
.A2(n_59),
.B(n_60),
.Y(n_1822)
);

A2O1A1Ixp33_ASAP7_75t_L g1823 ( 
.A1(n_1767),
.A2(n_63),
.B(n_61),
.C(n_62),
.Y(n_1823)
);

AOI21xp5_ASAP7_75t_L g1824 ( 
.A1(n_1756),
.A2(n_61),
.B(n_62),
.Y(n_1824)
);

NAND2xp5_ASAP7_75t_L g1825 ( 
.A(n_1749),
.B(n_64),
.Y(n_1825)
);

OAI21x1_ASAP7_75t_SL g1826 ( 
.A1(n_1769),
.A2(n_65),
.B(n_66),
.Y(n_1826)
);

NAND2xp5_ASAP7_75t_L g1827 ( 
.A(n_1652),
.B(n_65),
.Y(n_1827)
);

OAI21x1_ASAP7_75t_SL g1828 ( 
.A1(n_1676),
.A2(n_66),
.B(n_67),
.Y(n_1828)
);

INVx4_ASAP7_75t_L g1829 ( 
.A(n_1577),
.Y(n_1829)
);

BUFx12f_ASAP7_75t_L g1830 ( 
.A(n_1606),
.Y(n_1830)
);

OAI21xp33_ASAP7_75t_L g1831 ( 
.A1(n_1697),
.A2(n_1711),
.B(n_1674),
.Y(n_1831)
);

AND2x2_ASAP7_75t_L g1832 ( 
.A(n_1661),
.B(n_67),
.Y(n_1832)
);

NAND2xp5_ASAP7_75t_L g1833 ( 
.A(n_1589),
.B(n_68),
.Y(n_1833)
);

INVx5_ASAP7_75t_L g1834 ( 
.A(n_1698),
.Y(n_1834)
);

OAI21x1_ASAP7_75t_L g1835 ( 
.A1(n_1678),
.A2(n_304),
.B(n_303),
.Y(n_1835)
);

AOI21x1_ASAP7_75t_L g1836 ( 
.A1(n_1731),
.A2(n_309),
.B(n_305),
.Y(n_1836)
);

O2A1O1Ixp5_ASAP7_75t_L g1837 ( 
.A1(n_1750),
.A2(n_70),
.B(n_68),
.C(n_69),
.Y(n_1837)
);

OA21x2_ASAP7_75t_L g1838 ( 
.A1(n_1609),
.A2(n_312),
.B(n_311),
.Y(n_1838)
);

AOI21xp5_ASAP7_75t_L g1839 ( 
.A1(n_1756),
.A2(n_69),
.B(n_70),
.Y(n_1839)
);

AOI21xp5_ASAP7_75t_L g1840 ( 
.A1(n_1617),
.A2(n_71),
.B(n_72),
.Y(n_1840)
);

OAI21x1_ASAP7_75t_L g1841 ( 
.A1(n_1664),
.A2(n_1595),
.B(n_1584),
.Y(n_1841)
);

AOI21xp5_ASAP7_75t_L g1842 ( 
.A1(n_1698),
.A2(n_71),
.B(n_72),
.Y(n_1842)
);

AOI21xp5_ASAP7_75t_L g1843 ( 
.A1(n_1650),
.A2(n_73),
.B(n_74),
.Y(n_1843)
);

INVx1_ASAP7_75t_L g1844 ( 
.A(n_1597),
.Y(n_1844)
);

A2O1A1Ixp33_ASAP7_75t_L g1845 ( 
.A1(n_1665),
.A2(n_76),
.B(n_73),
.C(n_74),
.Y(n_1845)
);

AOI21xp5_ASAP7_75t_L g1846 ( 
.A1(n_1618),
.A2(n_76),
.B(n_77),
.Y(n_1846)
);

OAI21x1_ASAP7_75t_L g1847 ( 
.A1(n_1607),
.A2(n_315),
.B(n_314),
.Y(n_1847)
);

OAI21x1_ASAP7_75t_L g1848 ( 
.A1(n_1610),
.A2(n_317),
.B(n_316),
.Y(n_1848)
);

INVx2_ASAP7_75t_L g1849 ( 
.A(n_1586),
.Y(n_1849)
);

INVx1_ASAP7_75t_SL g1850 ( 
.A(n_1703),
.Y(n_1850)
);

AOI21xp33_ASAP7_75t_L g1851 ( 
.A1(n_1629),
.A2(n_77),
.B(n_78),
.Y(n_1851)
);

AOI21xp5_ASAP7_75t_L g1852 ( 
.A1(n_1628),
.A2(n_78),
.B(n_79),
.Y(n_1852)
);

AND2x4_ASAP7_75t_L g1853 ( 
.A(n_1614),
.B(n_80),
.Y(n_1853)
);

NAND2xp5_ASAP7_75t_L g1854 ( 
.A(n_1640),
.B(n_81),
.Y(n_1854)
);

NOR2xp33_ASAP7_75t_L g1855 ( 
.A(n_1691),
.B(n_81),
.Y(n_1855)
);

OAI21x1_ASAP7_75t_L g1856 ( 
.A1(n_1612),
.A2(n_320),
.B(n_319),
.Y(n_1856)
);

OAI22xp5_ASAP7_75t_L g1857 ( 
.A1(n_1708),
.A2(n_84),
.B1(n_82),
.B2(n_83),
.Y(n_1857)
);

BUFx2_ASAP7_75t_L g1858 ( 
.A(n_1666),
.Y(n_1858)
);

A2O1A1Ixp33_ASAP7_75t_L g1859 ( 
.A1(n_1718),
.A2(n_85),
.B(n_83),
.C(n_84),
.Y(n_1859)
);

AOI21xp5_ASAP7_75t_L g1860 ( 
.A1(n_1628),
.A2(n_86),
.B(n_87),
.Y(n_1860)
);

OAI21x1_ASAP7_75t_L g1861 ( 
.A1(n_1622),
.A2(n_322),
.B(n_321),
.Y(n_1861)
);

AND2x2_ASAP7_75t_L g1862 ( 
.A(n_1745),
.B(n_86),
.Y(n_1862)
);

OAI21xp5_ASAP7_75t_L g1863 ( 
.A1(n_1656),
.A2(n_88),
.B(n_89),
.Y(n_1863)
);

AOI21xp5_ASAP7_75t_L g1864 ( 
.A1(n_1710),
.A2(n_88),
.B(n_90),
.Y(n_1864)
);

INVx2_ASAP7_75t_L g1865 ( 
.A(n_1592),
.Y(n_1865)
);

AOI21xp33_ASAP7_75t_L g1866 ( 
.A1(n_1596),
.A2(n_90),
.B(n_91),
.Y(n_1866)
);

OAI21xp5_ASAP7_75t_L g1867 ( 
.A1(n_1671),
.A2(n_92),
.B(n_93),
.Y(n_1867)
);

AOI21xp5_ASAP7_75t_L g1868 ( 
.A1(n_1710),
.A2(n_92),
.B(n_93),
.Y(n_1868)
);

OAI22xp5_ASAP7_75t_L g1869 ( 
.A1(n_1722),
.A2(n_96),
.B1(n_94),
.B2(n_95),
.Y(n_1869)
);

OAI21x1_ASAP7_75t_L g1870 ( 
.A1(n_1625),
.A2(n_324),
.B(n_323),
.Y(n_1870)
);

OAI21x1_ASAP7_75t_L g1871 ( 
.A1(n_1667),
.A2(n_326),
.B(n_325),
.Y(n_1871)
);

NOR3xp33_ASAP7_75t_L g1872 ( 
.A(n_1713),
.B(n_1716),
.C(n_1772),
.Y(n_1872)
);

NAND2xp5_ASAP7_75t_L g1873 ( 
.A(n_1647),
.B(n_95),
.Y(n_1873)
);

AOI21xp5_ASAP7_75t_L g1874 ( 
.A1(n_1660),
.A2(n_96),
.B(n_97),
.Y(n_1874)
);

NAND2xp5_ASAP7_75t_L g1875 ( 
.A(n_1755),
.B(n_1742),
.Y(n_1875)
);

A2O1A1Ixp33_ASAP7_75t_L g1876 ( 
.A1(n_1727),
.A2(n_100),
.B(n_97),
.C(n_98),
.Y(n_1876)
);

AND2x2_ASAP7_75t_L g1877 ( 
.A(n_1623),
.B(n_98),
.Y(n_1877)
);

AOI21xp5_ASAP7_75t_L g1878 ( 
.A1(n_1660),
.A2(n_101),
.B(n_102),
.Y(n_1878)
);

AOI21xp5_ASAP7_75t_L g1879 ( 
.A1(n_1738),
.A2(n_103),
.B(n_104),
.Y(n_1879)
);

AOI21xp5_ASAP7_75t_L g1880 ( 
.A1(n_1738),
.A2(n_1744),
.B(n_1730),
.Y(n_1880)
);

NAND2xp5_ASAP7_75t_L g1881 ( 
.A(n_1594),
.B(n_103),
.Y(n_1881)
);

NAND2xp5_ASAP7_75t_L g1882 ( 
.A(n_1579),
.B(n_104),
.Y(n_1882)
);

OAI21x1_ASAP7_75t_L g1883 ( 
.A1(n_1670),
.A2(n_1677),
.B(n_1681),
.Y(n_1883)
);

OAI21x1_ASAP7_75t_L g1884 ( 
.A1(n_1700),
.A2(n_328),
.B(n_327),
.Y(n_1884)
);

AOI21xp5_ASAP7_75t_L g1885 ( 
.A1(n_1748),
.A2(n_1693),
.B(n_1641),
.Y(n_1885)
);

NAND2xp5_ASAP7_75t_SL g1886 ( 
.A(n_1765),
.B(n_105),
.Y(n_1886)
);

O2A1O1Ixp5_ASAP7_75t_L g1887 ( 
.A1(n_1669),
.A2(n_108),
.B(n_105),
.C(n_107),
.Y(n_1887)
);

A2O1A1Ixp33_ASAP7_75t_L g1888 ( 
.A1(n_1765),
.A2(n_110),
.B(n_108),
.C(n_109),
.Y(n_1888)
);

BUFx3_ASAP7_75t_L g1889 ( 
.A(n_1654),
.Y(n_1889)
);

NAND2xp5_ASAP7_75t_L g1890 ( 
.A(n_1580),
.B(n_109),
.Y(n_1890)
);

OAI21x1_ASAP7_75t_L g1891 ( 
.A1(n_1702),
.A2(n_331),
.B(n_330),
.Y(n_1891)
);

NOR2xp33_ASAP7_75t_L g1892 ( 
.A(n_1747),
.B(n_110),
.Y(n_1892)
);

CKINVDCx20_ASAP7_75t_R g1893 ( 
.A(n_1701),
.Y(n_1893)
);

A2O1A1Ixp33_ASAP7_75t_L g1894 ( 
.A1(n_1662),
.A2(n_113),
.B(n_111),
.C(n_112),
.Y(n_1894)
);

BUFx3_ASAP7_75t_L g1895 ( 
.A(n_1653),
.Y(n_1895)
);

INVx1_ASAP7_75t_L g1896 ( 
.A(n_1719),
.Y(n_1896)
);

AO31x2_ASAP7_75t_L g1897 ( 
.A1(n_1724),
.A2(n_333),
.A3(n_335),
.B(n_332),
.Y(n_1897)
);

OAI21x1_ASAP7_75t_L g1898 ( 
.A1(n_1754),
.A2(n_1758),
.B(n_1663),
.Y(n_1898)
);

INVx3_ASAP7_75t_L g1899 ( 
.A(n_1696),
.Y(n_1899)
);

NAND2xp5_ASAP7_75t_L g1900 ( 
.A(n_1752),
.B(n_111),
.Y(n_1900)
);

OAI22xp5_ASAP7_75t_L g1901 ( 
.A1(n_1598),
.A2(n_114),
.B1(n_112),
.B2(n_113),
.Y(n_1901)
);

OAI21xp5_ASAP7_75t_L g1902 ( 
.A1(n_1605),
.A2(n_114),
.B(n_115),
.Y(n_1902)
);

NAND2x1p5_ASAP7_75t_L g1903 ( 
.A(n_1577),
.B(n_336),
.Y(n_1903)
);

INVx2_ASAP7_75t_L g1904 ( 
.A(n_1602),
.Y(n_1904)
);

AOI221x1_ASAP7_75t_L g1905 ( 
.A1(n_1706),
.A2(n_117),
.B1(n_115),
.B2(n_116),
.C(n_118),
.Y(n_1905)
);

NAND2xp5_ASAP7_75t_L g1906 ( 
.A(n_1619),
.B(n_116),
.Y(n_1906)
);

INVx2_ASAP7_75t_L g1907 ( 
.A(n_1603),
.Y(n_1907)
);

AOI21xp5_ASAP7_75t_L g1908 ( 
.A1(n_1641),
.A2(n_117),
.B(n_118),
.Y(n_1908)
);

BUFx3_ASAP7_75t_L g1909 ( 
.A(n_1638),
.Y(n_1909)
);

NAND2x1p5_ASAP7_75t_L g1910 ( 
.A(n_1577),
.B(n_338),
.Y(n_1910)
);

AOI21x1_ASAP7_75t_L g1911 ( 
.A1(n_1578),
.A2(n_343),
.B(n_342),
.Y(n_1911)
);

AO31x2_ASAP7_75t_L g1912 ( 
.A1(n_1741),
.A2(n_345),
.A3(n_346),
.B(n_344),
.Y(n_1912)
);

INVx4_ASAP7_75t_L g1913 ( 
.A(n_1637),
.Y(n_1913)
);

NAND2xp5_ASAP7_75t_L g1914 ( 
.A(n_1614),
.B(n_119),
.Y(n_1914)
);

AND2x2_ASAP7_75t_L g1915 ( 
.A(n_1639),
.B(n_119),
.Y(n_1915)
);

NAND2xp5_ASAP7_75t_L g1916 ( 
.A(n_1620),
.B(n_120),
.Y(n_1916)
);

AOI21xp5_ASAP7_75t_L g1917 ( 
.A1(n_1763),
.A2(n_121),
.B(n_122),
.Y(n_1917)
);

A2O1A1Ixp33_ASAP7_75t_L g1918 ( 
.A1(n_1673),
.A2(n_125),
.B(n_123),
.C(n_124),
.Y(n_1918)
);

OAI21x1_ASAP7_75t_L g1919 ( 
.A1(n_1714),
.A2(n_349),
.B(n_347),
.Y(n_1919)
);

OAI21xp5_ASAP7_75t_L g1920 ( 
.A1(n_1658),
.A2(n_123),
.B(n_124),
.Y(n_1920)
);

AOI21xp5_ASAP7_75t_L g1921 ( 
.A1(n_1763),
.A2(n_126),
.B(n_127),
.Y(n_1921)
);

AND2x4_ASAP7_75t_L g1922 ( 
.A(n_1735),
.B(n_127),
.Y(n_1922)
);

OAI21xp5_ASAP7_75t_L g1923 ( 
.A1(n_1658),
.A2(n_128),
.B(n_129),
.Y(n_1923)
);

AND2x2_ASAP7_75t_L g1924 ( 
.A(n_1646),
.B(n_128),
.Y(n_1924)
);

BUFx6f_ASAP7_75t_L g1925 ( 
.A(n_1725),
.Y(n_1925)
);

AO31x2_ASAP7_75t_L g1926 ( 
.A1(n_1743),
.A2(n_352),
.A3(n_354),
.B(n_351),
.Y(n_1926)
);

NOR2xp33_ASAP7_75t_L g1927 ( 
.A(n_1712),
.B(n_129),
.Y(n_1927)
);

AND2x2_ASAP7_75t_L g1928 ( 
.A(n_1655),
.B(n_130),
.Y(n_1928)
);

AOI21xp5_ASAP7_75t_L g1929 ( 
.A1(n_1763),
.A2(n_130),
.B(n_132),
.Y(n_1929)
);

AOI22xp5_ASAP7_75t_SL g1930 ( 
.A1(n_1658),
.A2(n_135),
.B1(n_132),
.B2(n_133),
.Y(n_1930)
);

OR2x6_ASAP7_75t_L g1931 ( 
.A(n_1717),
.B(n_357),
.Y(n_1931)
);

HB1xp67_ASAP7_75t_L g1932 ( 
.A(n_1637),
.Y(n_1932)
);

AND2x4_ASAP7_75t_L g1933 ( 
.A(n_1735),
.B(n_133),
.Y(n_1933)
);

AO21x1_ASAP7_75t_L g1934 ( 
.A1(n_1673),
.A2(n_135),
.B(n_136),
.Y(n_1934)
);

AOI21xp5_ASAP7_75t_L g1935 ( 
.A1(n_1706),
.A2(n_136),
.B(n_137),
.Y(n_1935)
);

OAI21xp5_ASAP7_75t_L g1936 ( 
.A1(n_1658),
.A2(n_138),
.B(n_139),
.Y(n_1936)
);

AOI21x1_ASAP7_75t_L g1937 ( 
.A1(n_1643),
.A2(n_359),
.B(n_358),
.Y(n_1937)
);

BUFx3_ASAP7_75t_L g1938 ( 
.A(n_1690),
.Y(n_1938)
);

A2O1A1Ixp33_ASAP7_75t_L g1939 ( 
.A1(n_1643),
.A2(n_141),
.B(n_138),
.C(n_140),
.Y(n_1939)
);

OAI21xp5_ASAP7_75t_L g1940 ( 
.A1(n_1632),
.A2(n_1715),
.B(n_1729),
.Y(n_1940)
);

AOI21xp5_ASAP7_75t_SL g1941 ( 
.A1(n_1696),
.A2(n_141),
.B(n_142),
.Y(n_1941)
);

CKINVDCx5p33_ASAP7_75t_R g1942 ( 
.A(n_1721),
.Y(n_1942)
);

NAND2xp5_ASAP7_75t_L g1943 ( 
.A(n_1746),
.B(n_1753),
.Y(n_1943)
);

OR2x6_ASAP7_75t_L g1944 ( 
.A(n_1931),
.B(n_1636),
.Y(n_1944)
);

AOI21xp5_ASAP7_75t_L g1945 ( 
.A1(n_1780),
.A2(n_1739),
.B(n_1733),
.Y(n_1945)
);

OR2x6_ASAP7_75t_L g1946 ( 
.A(n_1931),
.B(n_1621),
.Y(n_1946)
);

NAND2xp5_ASAP7_75t_L g1947 ( 
.A(n_1858),
.B(n_1728),
.Y(n_1947)
);

AOI22xp5_ASAP7_75t_L g1948 ( 
.A1(n_1779),
.A2(n_1632),
.B1(n_1649),
.B2(n_1621),
.Y(n_1948)
);

AOI21xp5_ASAP7_75t_L g1949 ( 
.A1(n_1793),
.A2(n_1739),
.B(n_1733),
.Y(n_1949)
);

AOI22xp5_ASAP7_75t_L g1950 ( 
.A1(n_1831),
.A2(n_1649),
.B1(n_1714),
.B2(n_1725),
.Y(n_1950)
);

INVx8_ASAP7_75t_L g1951 ( 
.A(n_1830),
.Y(n_1951)
);

INVx2_ASAP7_75t_SL g1952 ( 
.A(n_1938),
.Y(n_1952)
);

AND2x4_ASAP7_75t_L g1953 ( 
.A(n_1810),
.B(n_1735),
.Y(n_1953)
);

NAND2xp5_ASAP7_75t_L g1954 ( 
.A(n_1792),
.B(n_1740),
.Y(n_1954)
);

CKINVDCx5p33_ASAP7_75t_R g1955 ( 
.A(n_1893),
.Y(n_1955)
);

NAND2xp5_ASAP7_75t_L g1956 ( 
.A(n_1810),
.B(n_1582),
.Y(n_1956)
);

OR2x2_ASAP7_75t_L g1957 ( 
.A(n_1844),
.B(n_1611),
.Y(n_1957)
);

NAND2x1p5_ASAP7_75t_L g1958 ( 
.A(n_1834),
.B(n_1582),
.Y(n_1958)
);

HB1xp67_ASAP7_75t_L g1959 ( 
.A(n_1790),
.Y(n_1959)
);

CKINVDCx20_ASAP7_75t_R g1960 ( 
.A(n_1785),
.Y(n_1960)
);

AND2x4_ASAP7_75t_L g1961 ( 
.A(n_1844),
.B(n_1582),
.Y(n_1961)
);

INVx2_ASAP7_75t_L g1962 ( 
.A(n_1849),
.Y(n_1962)
);

INVx1_ASAP7_75t_L g1963 ( 
.A(n_1896),
.Y(n_1963)
);

O2A1O1Ixp33_ASAP7_75t_L g1964 ( 
.A1(n_1819),
.A2(n_1707),
.B(n_1599),
.C(n_1682),
.Y(n_1964)
);

NAND2xp5_ASAP7_75t_L g1965 ( 
.A(n_1896),
.B(n_1804),
.Y(n_1965)
);

INVx2_ASAP7_75t_L g1966 ( 
.A(n_1865),
.Y(n_1966)
);

OR2x6_ASAP7_75t_L g1967 ( 
.A(n_1802),
.B(n_1624),
.Y(n_1967)
);

INVx1_ASAP7_75t_L g1968 ( 
.A(n_1804),
.Y(n_1968)
);

NAND2xp5_ASAP7_75t_L g1969 ( 
.A(n_1797),
.B(n_1599),
.Y(n_1969)
);

INVxp67_ASAP7_75t_SL g1970 ( 
.A(n_1875),
.Y(n_1970)
);

INVx1_ASAP7_75t_L g1971 ( 
.A(n_1883),
.Y(n_1971)
);

INVx2_ASAP7_75t_SL g1972 ( 
.A(n_1889),
.Y(n_1972)
);

AOI22xp33_ASAP7_75t_L g1973 ( 
.A1(n_1776),
.A2(n_1737),
.B1(n_1645),
.B2(n_1679),
.Y(n_1973)
);

INVx1_ASAP7_75t_L g1974 ( 
.A(n_1943),
.Y(n_1974)
);

INVx1_ASAP7_75t_L g1975 ( 
.A(n_1790),
.Y(n_1975)
);

BUFx3_ASAP7_75t_L g1976 ( 
.A(n_1895),
.Y(n_1976)
);

AND2x2_ASAP7_75t_L g1977 ( 
.A(n_1877),
.B(n_1783),
.Y(n_1977)
);

BUFx6f_ASAP7_75t_L g1978 ( 
.A(n_1909),
.Y(n_1978)
);

NAND2xp5_ASAP7_75t_L g1979 ( 
.A(n_1775),
.B(n_1659),
.Y(n_1979)
);

INVx2_ASAP7_75t_SL g1980 ( 
.A(n_1782),
.Y(n_1980)
);

BUFx2_ASAP7_75t_L g1981 ( 
.A(n_1821),
.Y(n_1981)
);

INVx1_ASAP7_75t_L g1982 ( 
.A(n_1790),
.Y(n_1982)
);

INVx4_ASAP7_75t_L g1983 ( 
.A(n_1782),
.Y(n_1983)
);

BUFx2_ASAP7_75t_SL g1984 ( 
.A(n_1834),
.Y(n_1984)
);

AOI22xp5_ASAP7_75t_L g1985 ( 
.A1(n_1872),
.A2(n_1725),
.B1(n_1624),
.B2(n_1726),
.Y(n_1985)
);

BUFx3_ASAP7_75t_L g1986 ( 
.A(n_1777),
.Y(n_1986)
);

INVx1_ASAP7_75t_L g1987 ( 
.A(n_1904),
.Y(n_1987)
);

NAND2xp5_ASAP7_75t_L g1988 ( 
.A(n_1880),
.B(n_1833),
.Y(n_1988)
);

NAND2xp5_ASAP7_75t_L g1989 ( 
.A(n_1862),
.B(n_1906),
.Y(n_1989)
);

INVx3_ASAP7_75t_SL g1990 ( 
.A(n_1814),
.Y(n_1990)
);

OR2x6_ASAP7_75t_L g1991 ( 
.A(n_1940),
.B(n_1624),
.Y(n_1991)
);

AND2x4_ASAP7_75t_L g1992 ( 
.A(n_1788),
.B(n_1648),
.Y(n_1992)
);

INVx2_ASAP7_75t_L g1993 ( 
.A(n_1907),
.Y(n_1993)
);

NOR2x1p5_ASAP7_75t_L g1994 ( 
.A(n_1829),
.B(n_1942),
.Y(n_1994)
);

INVx3_ASAP7_75t_L g1995 ( 
.A(n_1925),
.Y(n_1995)
);

INVx1_ASAP7_75t_L g1996 ( 
.A(n_1786),
.Y(n_1996)
);

BUFx2_ASAP7_75t_L g1997 ( 
.A(n_1932),
.Y(n_1997)
);

BUFx6f_ASAP7_75t_L g1998 ( 
.A(n_1925),
.Y(n_1998)
);

INVx1_ASAP7_75t_L g1999 ( 
.A(n_1882),
.Y(n_1999)
);

AOI21xp5_ASAP7_75t_L g2000 ( 
.A1(n_1791),
.A2(n_1739),
.B(n_1733),
.Y(n_2000)
);

AOI21xp5_ASAP7_75t_L g2001 ( 
.A1(n_1794),
.A2(n_1709),
.B(n_1682),
.Y(n_2001)
);

HB1xp67_ASAP7_75t_L g2002 ( 
.A(n_1898),
.Y(n_2002)
);

AOI22xp5_ASAP7_75t_L g2003 ( 
.A1(n_1902),
.A2(n_1726),
.B1(n_1608),
.B2(n_1709),
.Y(n_2003)
);

INVx5_ASAP7_75t_L g2004 ( 
.A(n_1834),
.Y(n_2004)
);

INVx1_ASAP7_75t_L g2005 ( 
.A(n_1890),
.Y(n_2005)
);

BUFx3_ASAP7_75t_L g2006 ( 
.A(n_1850),
.Y(n_2006)
);

NAND2xp5_ASAP7_75t_L g2007 ( 
.A(n_1806),
.B(n_1608),
.Y(n_2007)
);

INVx5_ASAP7_75t_L g2008 ( 
.A(n_1829),
.Y(n_2008)
);

NOR2xp33_ASAP7_75t_L g2009 ( 
.A(n_1807),
.B(n_1648),
.Y(n_2009)
);

AOI221xp5_ASAP7_75t_L g2010 ( 
.A1(n_1851),
.A2(n_1644),
.B1(n_1684),
.B2(n_1726),
.C(n_1686),
.Y(n_2010)
);

BUFx2_ASAP7_75t_R g2011 ( 
.A(n_1799),
.Y(n_2011)
);

AOI22xp33_ASAP7_75t_L g2012 ( 
.A1(n_1811),
.A2(n_1934),
.B1(n_1867),
.B2(n_1866),
.Y(n_2012)
);

AOI22xp5_ASAP7_75t_L g2013 ( 
.A1(n_1927),
.A2(n_1616),
.B1(n_1657),
.B2(n_1637),
.Y(n_2013)
);

INVx3_ASAP7_75t_L g2014 ( 
.A(n_1925),
.Y(n_2014)
);

BUFx12f_ASAP7_75t_L g2015 ( 
.A(n_1922),
.Y(n_2015)
);

AND2x2_ASAP7_75t_L g2016 ( 
.A(n_1832),
.B(n_1657),
.Y(n_2016)
);

NAND2xp5_ASAP7_75t_SL g2017 ( 
.A(n_1801),
.B(n_1680),
.Y(n_2017)
);

OR2x6_ASAP7_75t_L g2018 ( 
.A(n_1922),
.B(n_1705),
.Y(n_2018)
);

AOI221xp5_ASAP7_75t_L g2019 ( 
.A1(n_1813),
.A2(n_1694),
.B1(n_1688),
.B2(n_1687),
.C(n_145),
.Y(n_2019)
);

NAND2xp5_ASAP7_75t_L g2020 ( 
.A(n_1900),
.B(n_143),
.Y(n_2020)
);

BUFx2_ASAP7_75t_L g2021 ( 
.A(n_1899),
.Y(n_2021)
);

OR2x6_ASAP7_75t_L g2022 ( 
.A(n_1933),
.B(n_360),
.Y(n_2022)
);

INVx3_ASAP7_75t_L g2023 ( 
.A(n_1913),
.Y(n_2023)
);

BUFx6f_ASAP7_75t_L g2024 ( 
.A(n_1853),
.Y(n_2024)
);

A2O1A1Ixp33_ASAP7_75t_L g2025 ( 
.A1(n_1800),
.A2(n_145),
.B(n_143),
.C(n_144),
.Y(n_2025)
);

NOR2xp67_ASAP7_75t_L g2026 ( 
.A(n_1796),
.B(n_144),
.Y(n_2026)
);

INVx1_ASAP7_75t_L g2027 ( 
.A(n_1854),
.Y(n_2027)
);

INVx1_ASAP7_75t_L g2028 ( 
.A(n_1873),
.Y(n_2028)
);

NAND2x1_ASAP7_75t_L g2029 ( 
.A(n_1899),
.B(n_361),
.Y(n_2029)
);

AND2x4_ASAP7_75t_L g2030 ( 
.A(n_1788),
.B(n_362),
.Y(n_2030)
);

INVx2_ASAP7_75t_SL g2031 ( 
.A(n_1933),
.Y(n_2031)
);

AND2x4_ASAP7_75t_L g2032 ( 
.A(n_1913),
.B(n_363),
.Y(n_2032)
);

AOI22xp33_ASAP7_75t_L g2033 ( 
.A1(n_1920),
.A2(n_148),
.B1(n_146),
.B2(n_147),
.Y(n_2033)
);

NOR2xp67_ASAP7_75t_L g2034 ( 
.A(n_1827),
.B(n_147),
.Y(n_2034)
);

INVx2_ASAP7_75t_SL g2035 ( 
.A(n_1809),
.Y(n_2035)
);

AND2x2_ASAP7_75t_L g2036 ( 
.A(n_1809),
.B(n_149),
.Y(n_2036)
);

INVx3_ASAP7_75t_L g2037 ( 
.A(n_1853),
.Y(n_2037)
);

CKINVDCx5p33_ASAP7_75t_R g2038 ( 
.A(n_1924),
.Y(n_2038)
);

BUFx10_ASAP7_75t_L g2039 ( 
.A(n_1855),
.Y(n_2039)
);

BUFx6f_ASAP7_75t_L g2040 ( 
.A(n_1914),
.Y(n_2040)
);

INVx3_ASAP7_75t_L g2041 ( 
.A(n_1903),
.Y(n_2041)
);

INVx2_ASAP7_75t_L g2042 ( 
.A(n_1841),
.Y(n_2042)
);

BUFx3_ASAP7_75t_L g2043 ( 
.A(n_1916),
.Y(n_2043)
);

BUFx2_ASAP7_75t_L g2044 ( 
.A(n_1774),
.Y(n_2044)
);

NAND2x1p5_ASAP7_75t_L g2045 ( 
.A(n_1816),
.B(n_364),
.Y(n_2045)
);

HB1xp67_ASAP7_75t_L g2046 ( 
.A(n_1778),
.Y(n_2046)
);

BUFx4f_ASAP7_75t_L g2047 ( 
.A(n_1910),
.Y(n_2047)
);

NAND2xp5_ASAP7_75t_SL g2048 ( 
.A(n_1885),
.B(n_366),
.Y(n_2048)
);

INVx2_ASAP7_75t_L g2049 ( 
.A(n_1789),
.Y(n_2049)
);

BUFx3_ASAP7_75t_L g2050 ( 
.A(n_1808),
.Y(n_2050)
);

INVx1_ASAP7_75t_L g2051 ( 
.A(n_1784),
.Y(n_2051)
);

BUFx2_ASAP7_75t_L g2052 ( 
.A(n_1781),
.Y(n_2052)
);

BUFx6f_ASAP7_75t_L g2053 ( 
.A(n_1787),
.Y(n_2053)
);

INVx1_ASAP7_75t_L g2054 ( 
.A(n_1965),
.Y(n_2054)
);

INVxp33_ASAP7_75t_L g2055 ( 
.A(n_2009),
.Y(n_2055)
);

INVx1_ASAP7_75t_L g2056 ( 
.A(n_1963),
.Y(n_2056)
);

INVx2_ASAP7_75t_L g2057 ( 
.A(n_1968),
.Y(n_2057)
);

BUFx2_ASAP7_75t_L g2058 ( 
.A(n_1981),
.Y(n_2058)
);

NOR2xp67_ASAP7_75t_L g2059 ( 
.A(n_1983),
.B(n_1988),
.Y(n_2059)
);

CKINVDCx11_ASAP7_75t_R g2060 ( 
.A(n_1960),
.Y(n_2060)
);

OAI21x1_ASAP7_75t_L g2061 ( 
.A1(n_1945),
.A2(n_1937),
.B(n_1836),
.Y(n_2061)
);

OA21x2_ASAP7_75t_L g2062 ( 
.A1(n_1975),
.A2(n_1936),
.B(n_1923),
.Y(n_2062)
);

INVx1_ASAP7_75t_L g2063 ( 
.A(n_1957),
.Y(n_2063)
);

NAND2x1p5_ASAP7_75t_L g2064 ( 
.A(n_2004),
.B(n_1930),
.Y(n_2064)
);

AOI21x1_ASAP7_75t_L g2065 ( 
.A1(n_2046),
.A2(n_1911),
.B(n_1798),
.Y(n_2065)
);

OAI21x1_ASAP7_75t_SL g2066 ( 
.A1(n_1964),
.A2(n_1828),
.B(n_1822),
.Y(n_2066)
);

INVx1_ASAP7_75t_L g2067 ( 
.A(n_1974),
.Y(n_2067)
);

BUFx2_ASAP7_75t_L g2068 ( 
.A(n_1981),
.Y(n_2068)
);

OAI21x1_ASAP7_75t_L g2069 ( 
.A1(n_2000),
.A2(n_2001),
.B(n_1949),
.Y(n_2069)
);

INVx3_ASAP7_75t_L g2070 ( 
.A(n_1961),
.Y(n_2070)
);

OAI21x1_ASAP7_75t_L g2071 ( 
.A1(n_2051),
.A2(n_1812),
.B(n_1847),
.Y(n_2071)
);

AOI221xp5_ASAP7_75t_L g2072 ( 
.A1(n_2025),
.A2(n_1869),
.B1(n_1857),
.B2(n_1845),
.C(n_1859),
.Y(n_2072)
);

OAI21x1_ASAP7_75t_L g2073 ( 
.A1(n_2049),
.A2(n_1856),
.B(n_1848),
.Y(n_2073)
);

AO21x2_ASAP7_75t_L g2074 ( 
.A1(n_1982),
.A2(n_1840),
.B(n_1826),
.Y(n_2074)
);

INVx2_ASAP7_75t_L g2075 ( 
.A(n_1962),
.Y(n_2075)
);

NOR2xp33_ASAP7_75t_L g2076 ( 
.A(n_1969),
.B(n_1817),
.Y(n_2076)
);

BUFx6f_ASAP7_75t_L g2077 ( 
.A(n_2047),
.Y(n_2077)
);

INVxp67_ASAP7_75t_L g2078 ( 
.A(n_1997),
.Y(n_2078)
);

AOI21xp5_ASAP7_75t_L g2079 ( 
.A1(n_2048),
.A2(n_1935),
.B(n_1879),
.Y(n_2079)
);

INVx4_ASAP7_75t_L g2080 ( 
.A(n_2008),
.Y(n_2080)
);

INVx2_ASAP7_75t_L g2081 ( 
.A(n_1966),
.Y(n_2081)
);

CKINVDCx11_ASAP7_75t_R g2082 ( 
.A(n_1990),
.Y(n_2082)
);

NOR2xp67_ASAP7_75t_L g2083 ( 
.A(n_1980),
.B(n_1818),
.Y(n_2083)
);

INVx1_ASAP7_75t_L g2084 ( 
.A(n_1970),
.Y(n_2084)
);

OA21x2_ASAP7_75t_L g2085 ( 
.A1(n_2052),
.A2(n_2044),
.B(n_1996),
.Y(n_2085)
);

INVx2_ASAP7_75t_L g2086 ( 
.A(n_1993),
.Y(n_2086)
);

O2A1O1Ixp33_ASAP7_75t_L g2087 ( 
.A1(n_2017),
.A2(n_1820),
.B(n_1823),
.C(n_1894),
.Y(n_2087)
);

OAI21x1_ASAP7_75t_L g2088 ( 
.A1(n_2007),
.A2(n_1870),
.B(n_1861),
.Y(n_2088)
);

OA21x2_ASAP7_75t_L g2089 ( 
.A1(n_2052),
.A2(n_1905),
.B(n_1884),
.Y(n_2089)
);

OR2x2_ASAP7_75t_L g2090 ( 
.A(n_1947),
.B(n_1997),
.Y(n_2090)
);

OAI21x1_ASAP7_75t_L g2091 ( 
.A1(n_2042),
.A2(n_1891),
.B(n_1871),
.Y(n_2091)
);

OAI21x1_ASAP7_75t_L g2092 ( 
.A1(n_2029),
.A2(n_1919),
.B(n_1838),
.Y(n_2092)
);

OAI222xp33_ASAP7_75t_L g2093 ( 
.A1(n_2012),
.A2(n_1795),
.B1(n_1901),
.B2(n_1908),
.C1(n_1868),
.C2(n_1864),
.Y(n_2093)
);

NAND2x1p5_ASAP7_75t_L g2094 ( 
.A(n_2004),
.B(n_1838),
.Y(n_2094)
);

INVx2_ASAP7_75t_L g2095 ( 
.A(n_1987),
.Y(n_2095)
);

INVx1_ASAP7_75t_L g2096 ( 
.A(n_1954),
.Y(n_2096)
);

INVx1_ASAP7_75t_L g2097 ( 
.A(n_1956),
.Y(n_2097)
);

OR2x6_ASAP7_75t_L g2098 ( 
.A(n_1984),
.B(n_1815),
.Y(n_2098)
);

OAI21xp5_ASAP7_75t_L g2099 ( 
.A1(n_2034),
.A2(n_1888),
.B(n_1876),
.Y(n_2099)
);

AND2x2_ASAP7_75t_L g2100 ( 
.A(n_1977),
.B(n_1915),
.Y(n_2100)
);

OAI21x1_ASAP7_75t_L g2101 ( 
.A1(n_2029),
.A2(n_1835),
.B(n_1824),
.Y(n_2101)
);

AO21x2_ASAP7_75t_L g2102 ( 
.A1(n_1959),
.A2(n_1846),
.B(n_1939),
.Y(n_2102)
);

OA21x2_ASAP7_75t_L g2103 ( 
.A1(n_2044),
.A2(n_1839),
.B(n_1887),
.Y(n_2103)
);

OAI21xp5_ASAP7_75t_L g2104 ( 
.A1(n_2033),
.A2(n_1918),
.B(n_1843),
.Y(n_2104)
);

INVx1_ASAP7_75t_L g2105 ( 
.A(n_1971),
.Y(n_2105)
);

AOI21xp5_ASAP7_75t_L g2106 ( 
.A1(n_2002),
.A2(n_1863),
.B(n_1874),
.Y(n_2106)
);

NOR3xp33_ASAP7_75t_SL g2107 ( 
.A(n_1955),
.B(n_1892),
.C(n_1917),
.Y(n_2107)
);

OA21x2_ASAP7_75t_L g2108 ( 
.A1(n_2021),
.A2(n_1837),
.B(n_1842),
.Y(n_2108)
);

OAI21x1_ASAP7_75t_L g2109 ( 
.A1(n_1958),
.A2(n_1878),
.B(n_1805),
.Y(n_2109)
);

INVx2_ASAP7_75t_L g2110 ( 
.A(n_1961),
.Y(n_2110)
);

OAI22xp33_ASAP7_75t_L g2111 ( 
.A1(n_2022),
.A2(n_1825),
.B1(n_1886),
.B2(n_1860),
.Y(n_2111)
);

A2O1A1Ixp33_ASAP7_75t_L g2112 ( 
.A1(n_2019),
.A2(n_1852),
.B(n_1929),
.C(n_1921),
.Y(n_2112)
);

CKINVDCx6p67_ASAP7_75t_R g2113 ( 
.A(n_1951),
.Y(n_2113)
);

OAI21x1_ASAP7_75t_L g2114 ( 
.A1(n_2023),
.A2(n_1803),
.B(n_1941),
.Y(n_2114)
);

OAI21x1_ASAP7_75t_L g2115 ( 
.A1(n_1995),
.A2(n_2014),
.B(n_2045),
.Y(n_2115)
);

INVx3_ASAP7_75t_L g2116 ( 
.A(n_2080),
.Y(n_2116)
);

AOI22xp33_ASAP7_75t_L g2117 ( 
.A1(n_2072),
.A2(n_2010),
.B1(n_1989),
.B2(n_2026),
.Y(n_2117)
);

AOI221xp5_ASAP7_75t_L g2118 ( 
.A1(n_2099),
.A2(n_2020),
.B1(n_2028),
.B2(n_2027),
.C(n_1999),
.Y(n_2118)
);

AND2x2_ASAP7_75t_L g2119 ( 
.A(n_2058),
.B(n_2016),
.Y(n_2119)
);

AOI22xp33_ASAP7_75t_L g2120 ( 
.A1(n_2104),
.A2(n_2043),
.B1(n_2050),
.B2(n_2005),
.Y(n_2120)
);

INVx4_ASAP7_75t_SL g2121 ( 
.A(n_2098),
.Y(n_2121)
);

OR2x6_ASAP7_75t_L g2122 ( 
.A(n_2064),
.B(n_1984),
.Y(n_2122)
);

OR2x2_ASAP7_75t_L g2123 ( 
.A(n_2090),
.B(n_1979),
.Y(n_2123)
);

AND2x2_ASAP7_75t_L g2124 ( 
.A(n_2068),
.B(n_2006),
.Y(n_2124)
);

NOR2xp33_ASAP7_75t_L g2125 ( 
.A(n_2055),
.B(n_2039),
.Y(n_2125)
);

AOI22xp33_ASAP7_75t_L g2126 ( 
.A1(n_2062),
.A2(n_1928),
.B1(n_2022),
.B2(n_1946),
.Y(n_2126)
);

AND2x2_ASAP7_75t_L g2127 ( 
.A(n_2055),
.B(n_1976),
.Y(n_2127)
);

OAI22xp5_ASAP7_75t_L g2128 ( 
.A1(n_2111),
.A2(n_2087),
.B1(n_2107),
.B2(n_2112),
.Y(n_2128)
);

AND2x2_ASAP7_75t_L g2129 ( 
.A(n_2078),
.B(n_2021),
.Y(n_2129)
);

AO221x2_ASAP7_75t_L g2130 ( 
.A1(n_2111),
.A2(n_1881),
.B1(n_2011),
.B2(n_1994),
.C(n_152),
.Y(n_2130)
);

AOI21xp5_ASAP7_75t_L g2131 ( 
.A1(n_2106),
.A2(n_1944),
.B(n_2004),
.Y(n_2131)
);

OR2x6_ASAP7_75t_L g2132 ( 
.A(n_2064),
.B(n_1944),
.Y(n_2132)
);

INVx1_ASAP7_75t_L g2133 ( 
.A(n_2057),
.Y(n_2133)
);

OR2x6_ASAP7_75t_L g2134 ( 
.A(n_2098),
.B(n_2069),
.Y(n_2134)
);

HB1xp67_ASAP7_75t_L g2135 ( 
.A(n_2078),
.Y(n_2135)
);

AND2x4_ASAP7_75t_L g2136 ( 
.A(n_2070),
.B(n_1953),
.Y(n_2136)
);

CKINVDCx5p33_ASAP7_75t_R g2137 ( 
.A(n_2060),
.Y(n_2137)
);

NAND2xp5_ASAP7_75t_L g2138 ( 
.A(n_2084),
.B(n_1953),
.Y(n_2138)
);

INVx2_ASAP7_75t_L g2139 ( 
.A(n_2105),
.Y(n_2139)
);

AND2x2_ASAP7_75t_L g2140 ( 
.A(n_2100),
.B(n_1952),
.Y(n_2140)
);

NAND2xp33_ASAP7_75t_L g2141 ( 
.A(n_2077),
.B(n_1978),
.Y(n_2141)
);

BUFx3_ASAP7_75t_L g2142 ( 
.A(n_2082),
.Y(n_2142)
);

AOI22xp33_ASAP7_75t_L g2143 ( 
.A1(n_2062),
.A2(n_1946),
.B1(n_2040),
.B2(n_2036),
.Y(n_2143)
);

INVx1_ASAP7_75t_L g2144 ( 
.A(n_2057),
.Y(n_2144)
);

INVx1_ASAP7_75t_L g2145 ( 
.A(n_2056),
.Y(n_2145)
);

AOI21xp33_ASAP7_75t_L g2146 ( 
.A1(n_2066),
.A2(n_2053),
.B(n_1991),
.Y(n_2146)
);

NOR2x1p5_ASAP7_75t_L g2147 ( 
.A(n_2113),
.B(n_2015),
.Y(n_2147)
);

OAI22xp33_ASAP7_75t_L g2148 ( 
.A1(n_2098),
.A2(n_2037),
.B1(n_2035),
.B2(n_2003),
.Y(n_2148)
);

INVx2_ASAP7_75t_L g2149 ( 
.A(n_2075),
.Y(n_2149)
);

AOI222xp33_ASAP7_75t_L g2150 ( 
.A1(n_2093),
.A2(n_1973),
.B1(n_2040),
.B2(n_2030),
.C1(n_2024),
.C2(n_2031),
.Y(n_2150)
);

BUFx3_ASAP7_75t_L g2151 ( 
.A(n_2082),
.Y(n_2151)
);

INVx4_ASAP7_75t_L g2152 ( 
.A(n_2077),
.Y(n_2152)
);

AND2x2_ASAP7_75t_L g2153 ( 
.A(n_2070),
.B(n_1972),
.Y(n_2153)
);

AND2x2_ASAP7_75t_L g2154 ( 
.A(n_2119),
.B(n_2059),
.Y(n_2154)
);

INVx1_ASAP7_75t_L g2155 ( 
.A(n_2139),
.Y(n_2155)
);

INVx1_ASAP7_75t_SL g2156 ( 
.A(n_2137),
.Y(n_2156)
);

INVx2_ASAP7_75t_L g2157 ( 
.A(n_2139),
.Y(n_2157)
);

AND2x4_ASAP7_75t_L g2158 ( 
.A(n_2134),
.B(n_2110),
.Y(n_2158)
);

INVx1_ASAP7_75t_L g2159 ( 
.A(n_2133),
.Y(n_2159)
);

INVx1_ASAP7_75t_L g2160 ( 
.A(n_2144),
.Y(n_2160)
);

INVx1_ASAP7_75t_L g2161 ( 
.A(n_2145),
.Y(n_2161)
);

INVx2_ASAP7_75t_L g2162 ( 
.A(n_2149),
.Y(n_2162)
);

INVx1_ASAP7_75t_L g2163 ( 
.A(n_2135),
.Y(n_2163)
);

INVx1_ASAP7_75t_L g2164 ( 
.A(n_2129),
.Y(n_2164)
);

INVx2_ASAP7_75t_L g2165 ( 
.A(n_2149),
.Y(n_2165)
);

INVx1_ASAP7_75t_L g2166 ( 
.A(n_2123),
.Y(n_2166)
);

INVx1_ASAP7_75t_L g2167 ( 
.A(n_2138),
.Y(n_2167)
);

NAND2xp5_ASAP7_75t_L g2168 ( 
.A(n_2124),
.B(n_2076),
.Y(n_2168)
);

NAND2xp5_ASAP7_75t_SL g2169 ( 
.A(n_2121),
.B(n_2083),
.Y(n_2169)
);

INVx2_ASAP7_75t_L g2170 ( 
.A(n_2134),
.Y(n_2170)
);

HB1xp67_ASAP7_75t_L g2171 ( 
.A(n_2134),
.Y(n_2171)
);

INVx2_ASAP7_75t_L g2172 ( 
.A(n_2122),
.Y(n_2172)
);

INVx2_ASAP7_75t_L g2173 ( 
.A(n_2122),
.Y(n_2173)
);

OR2x6_ASAP7_75t_L g2174 ( 
.A(n_2132),
.B(n_2094),
.Y(n_2174)
);

OR2x2_ASAP7_75t_L g2175 ( 
.A(n_2136),
.B(n_2097),
.Y(n_2175)
);

INVx2_ASAP7_75t_L g2176 ( 
.A(n_2122),
.Y(n_2176)
);

AND2x4_ASAP7_75t_L g2177 ( 
.A(n_2172),
.B(n_2121),
.Y(n_2177)
);

OAI22xp5_ASAP7_75t_L g2178 ( 
.A1(n_2168),
.A2(n_2128),
.B1(n_2126),
.B2(n_2120),
.Y(n_2178)
);

INVx2_ASAP7_75t_SL g2179 ( 
.A(n_2156),
.Y(n_2179)
);

INVx1_ASAP7_75t_SL g2180 ( 
.A(n_2154),
.Y(n_2180)
);

OAI22xp5_ASAP7_75t_L g2181 ( 
.A1(n_2167),
.A2(n_2126),
.B1(n_2120),
.B2(n_2132),
.Y(n_2181)
);

OAI211xp5_ASAP7_75t_L g2182 ( 
.A1(n_2163),
.A2(n_2117),
.B(n_2107),
.C(n_2118),
.Y(n_2182)
);

OAI22xp33_ASAP7_75t_L g2183 ( 
.A1(n_2174),
.A2(n_2132),
.B1(n_2148),
.B2(n_2131),
.Y(n_2183)
);

OAI221xp5_ASAP7_75t_L g2184 ( 
.A1(n_2171),
.A2(n_2117),
.B1(n_2143),
.B2(n_2150),
.C(n_2112),
.Y(n_2184)
);

OAI22xp5_ASAP7_75t_L g2185 ( 
.A1(n_2164),
.A2(n_2125),
.B1(n_2143),
.B2(n_2148),
.Y(n_2185)
);

AND2x2_ASAP7_75t_L g2186 ( 
.A(n_2172),
.B(n_2127),
.Y(n_2186)
);

NAND3xp33_ASAP7_75t_L g2187 ( 
.A(n_2171),
.B(n_2130),
.C(n_2076),
.Y(n_2187)
);

OR2x2_ASAP7_75t_L g2188 ( 
.A(n_2180),
.B(n_2166),
.Y(n_2188)
);

INVx1_ASAP7_75t_SL g2189 ( 
.A(n_2179),
.Y(n_2189)
);

NAND2xp5_ASAP7_75t_L g2190 ( 
.A(n_2182),
.B(n_2161),
.Y(n_2190)
);

NOR2xp67_ASAP7_75t_L g2191 ( 
.A(n_2187),
.B(n_2137),
.Y(n_2191)
);

OR2x2_ASAP7_75t_L g2192 ( 
.A(n_2178),
.B(n_2175),
.Y(n_2192)
);

NAND2xp5_ASAP7_75t_L g2193 ( 
.A(n_2186),
.B(n_2159),
.Y(n_2193)
);

INVxp67_ASAP7_75t_L g2194 ( 
.A(n_2191),
.Y(n_2194)
);

NAND2xp5_ASAP7_75t_L g2195 ( 
.A(n_2190),
.B(n_2189),
.Y(n_2195)
);

AO21x2_ASAP7_75t_L g2196 ( 
.A1(n_2192),
.A2(n_2183),
.B(n_2184),
.Y(n_2196)
);

AOI31xp33_ASAP7_75t_L g2197 ( 
.A1(n_2188),
.A2(n_2125),
.A3(n_2038),
.B(n_2169),
.Y(n_2197)
);

OAI31xp33_ASAP7_75t_L g2198 ( 
.A1(n_2193),
.A2(n_2181),
.A3(n_2130),
.B(n_2093),
.Y(n_2198)
);

NAND2xp5_ASAP7_75t_L g2199 ( 
.A(n_2190),
.B(n_2185),
.Y(n_2199)
);

OR2x2_ASAP7_75t_L g2200 ( 
.A(n_2190),
.B(n_2173),
.Y(n_2200)
);

AND2x2_ASAP7_75t_L g2201 ( 
.A(n_2189),
.B(n_2142),
.Y(n_2201)
);

AO21x2_ASAP7_75t_L g2202 ( 
.A1(n_2190),
.A2(n_2146),
.B(n_2169),
.Y(n_2202)
);

XOR2x2_ASAP7_75t_L g2203 ( 
.A(n_2199),
.B(n_2142),
.Y(n_2203)
);

AND2x2_ASAP7_75t_L g2204 ( 
.A(n_2201),
.B(n_2151),
.Y(n_2204)
);

NAND3xp33_ASAP7_75t_L g2205 ( 
.A(n_2198),
.B(n_2130),
.C(n_2079),
.Y(n_2205)
);

AOI22xp33_ASAP7_75t_L g2206 ( 
.A1(n_2198),
.A2(n_2196),
.B1(n_2195),
.B2(n_2200),
.Y(n_2206)
);

OR2x2_ASAP7_75t_L g2207 ( 
.A(n_2194),
.B(n_2151),
.Y(n_2207)
);

AND2x2_ASAP7_75t_L g2208 ( 
.A(n_2196),
.B(n_2060),
.Y(n_2208)
);

AOI22xp33_ASAP7_75t_L g2209 ( 
.A1(n_2202),
.A2(n_2170),
.B1(n_2102),
.B2(n_2174),
.Y(n_2209)
);

NOR3xp33_ASAP7_75t_L g2210 ( 
.A(n_2197),
.B(n_2152),
.C(n_2141),
.Y(n_2210)
);

AND2x2_ASAP7_75t_L g2211 ( 
.A(n_2202),
.B(n_2147),
.Y(n_2211)
);

NAND2xp5_ASAP7_75t_SL g2212 ( 
.A(n_2197),
.B(n_2173),
.Y(n_2212)
);

AND2x2_ASAP7_75t_L g2213 ( 
.A(n_2201),
.B(n_2140),
.Y(n_2213)
);

INVx1_ASAP7_75t_L g2214 ( 
.A(n_2205),
.Y(n_2214)
);

OAI31xp33_ASAP7_75t_L g2215 ( 
.A1(n_2206),
.A2(n_2170),
.A3(n_2177),
.B(n_2176),
.Y(n_2215)
);

OR2x2_ASAP7_75t_L g2216 ( 
.A(n_2208),
.B(n_2176),
.Y(n_2216)
);

OR2x2_ASAP7_75t_L g2217 ( 
.A(n_2207),
.B(n_2160),
.Y(n_2217)
);

OAI221xp5_ASAP7_75t_L g2218 ( 
.A1(n_2206),
.A2(n_2209),
.B1(n_2211),
.B2(n_2203),
.C(n_2212),
.Y(n_2218)
);

NAND3xp33_ASAP7_75t_L g2219 ( 
.A(n_2204),
.B(n_2141),
.C(n_2152),
.Y(n_2219)
);

BUFx3_ASAP7_75t_L g2220 ( 
.A(n_2213),
.Y(n_2220)
);

AND2x2_ASAP7_75t_L g2221 ( 
.A(n_2210),
.B(n_1978),
.Y(n_2221)
);

OR2x2_ASAP7_75t_L g2222 ( 
.A(n_2210),
.B(n_2155),
.Y(n_2222)
);

AND2x2_ASAP7_75t_L g2223 ( 
.A(n_2220),
.B(n_1986),
.Y(n_2223)
);

INVx1_ASAP7_75t_L g2224 ( 
.A(n_2217),
.Y(n_2224)
);

AND2x2_ASAP7_75t_L g2225 ( 
.A(n_2221),
.B(n_2214),
.Y(n_2225)
);

NAND2xp5_ASAP7_75t_L g2226 ( 
.A(n_2214),
.B(n_2157),
.Y(n_2226)
);

AND2x2_ASAP7_75t_L g2227 ( 
.A(n_2223),
.B(n_2219),
.Y(n_2227)
);

OR2x2_ASAP7_75t_L g2228 ( 
.A(n_2224),
.B(n_2216),
.Y(n_2228)
);

INVx2_ASAP7_75t_L g2229 ( 
.A(n_2225),
.Y(n_2229)
);

INVx4_ASAP7_75t_L g2230 ( 
.A(n_2226),
.Y(n_2230)
);

OR2x6_ASAP7_75t_L g2231 ( 
.A(n_2229),
.B(n_1951),
.Y(n_2231)
);

A2O1A1Ixp33_ASAP7_75t_L g2232 ( 
.A1(n_2228),
.A2(n_2218),
.B(n_2215),
.C(n_2226),
.Y(n_2232)
);

INVx1_ASAP7_75t_L g2233 ( 
.A(n_2230),
.Y(n_2233)
);

BUFx3_ASAP7_75t_L g2234 ( 
.A(n_2227),
.Y(n_2234)
);

NAND2xp5_ASAP7_75t_L g2235 ( 
.A(n_2230),
.B(n_2222),
.Y(n_2235)
);

AND2x2_ASAP7_75t_L g2236 ( 
.A(n_2229),
.B(n_2152),
.Y(n_2236)
);

NAND2xp5_ASAP7_75t_L g2237 ( 
.A(n_2234),
.B(n_2233),
.Y(n_2237)
);

AOI22xp5_ASAP7_75t_L g2238 ( 
.A1(n_2231),
.A2(n_2077),
.B1(n_2177),
.B2(n_2174),
.Y(n_2238)
);

INVx1_ASAP7_75t_L g2239 ( 
.A(n_2235),
.Y(n_2239)
);

INVx1_ASAP7_75t_SL g2240 ( 
.A(n_2231),
.Y(n_2240)
);

INVx1_ASAP7_75t_L g2241 ( 
.A(n_2236),
.Y(n_2241)
);

INVx1_ASAP7_75t_L g2242 ( 
.A(n_2232),
.Y(n_2242)
);

NAND3xp33_ASAP7_75t_L g2243 ( 
.A(n_2234),
.B(n_2032),
.C(n_2077),
.Y(n_2243)
);

INVxp67_ASAP7_75t_L g2244 ( 
.A(n_2234),
.Y(n_2244)
);

NAND2xp5_ASAP7_75t_L g2245 ( 
.A(n_2234),
.B(n_2157),
.Y(n_2245)
);

A2O1A1Ixp33_ASAP7_75t_L g2246 ( 
.A1(n_2232),
.A2(n_2114),
.B(n_2115),
.C(n_1948),
.Y(n_2246)
);

XNOR2x2_ASAP7_75t_L g2247 ( 
.A(n_2240),
.B(n_2013),
.Y(n_2247)
);

INVx1_ASAP7_75t_L g2248 ( 
.A(n_2244),
.Y(n_2248)
);

OAI22xp5_ASAP7_75t_L g2249 ( 
.A1(n_2239),
.A2(n_2174),
.B1(n_2041),
.B2(n_2116),
.Y(n_2249)
);

AOI21xp33_ASAP7_75t_L g2250 ( 
.A1(n_2242),
.A2(n_2067),
.B(n_2030),
.Y(n_2250)
);

AND2x2_ASAP7_75t_L g2251 ( 
.A(n_2241),
.B(n_2153),
.Y(n_2251)
);

XOR2xp5_ASAP7_75t_L g2252 ( 
.A(n_2243),
.B(n_2024),
.Y(n_2252)
);

AOI22xp33_ASAP7_75t_SL g2253 ( 
.A1(n_2245),
.A2(n_2089),
.B1(n_2102),
.B2(n_2103),
.Y(n_2253)
);

NAND2xp5_ASAP7_75t_L g2254 ( 
.A(n_2237),
.B(n_2054),
.Y(n_2254)
);

NOR2x1_ASAP7_75t_L g2255 ( 
.A(n_2246),
.B(n_2032),
.Y(n_2255)
);

NAND2xp5_ASAP7_75t_L g2256 ( 
.A(n_2238),
.B(n_2085),
.Y(n_2256)
);

INVx1_ASAP7_75t_L g2257 ( 
.A(n_2244),
.Y(n_2257)
);

NOR2xp33_ASAP7_75t_L g2258 ( 
.A(n_2244),
.B(n_1967),
.Y(n_2258)
);

INVx1_ASAP7_75t_L g2259 ( 
.A(n_2244),
.Y(n_2259)
);

NAND2xp5_ASAP7_75t_L g2260 ( 
.A(n_2251),
.B(n_150),
.Y(n_2260)
);

AOI21xp33_ASAP7_75t_L g2261 ( 
.A1(n_2248),
.A2(n_150),
.B(n_151),
.Y(n_2261)
);

BUFx2_ASAP7_75t_L g2262 ( 
.A(n_2257),
.Y(n_2262)
);

NAND2xp5_ASAP7_75t_L g2263 ( 
.A(n_2259),
.B(n_151),
.Y(n_2263)
);

AND2x2_ASAP7_75t_L g2264 ( 
.A(n_2258),
.B(n_2116),
.Y(n_2264)
);

INVx1_ASAP7_75t_L g2265 ( 
.A(n_2254),
.Y(n_2265)
);

INVx1_ASAP7_75t_L g2266 ( 
.A(n_2247),
.Y(n_2266)
);

INVx1_ASAP7_75t_L g2267 ( 
.A(n_2252),
.Y(n_2267)
);

XOR2x2_ASAP7_75t_L g2268 ( 
.A(n_2255),
.B(n_1950),
.Y(n_2268)
);

XNOR2x1_ASAP7_75t_L g2269 ( 
.A(n_2249),
.B(n_2256),
.Y(n_2269)
);

INVx1_ASAP7_75t_L g2270 ( 
.A(n_2250),
.Y(n_2270)
);

NOR2xp33_ASAP7_75t_L g2271 ( 
.A(n_2253),
.B(n_152),
.Y(n_2271)
);

INVx1_ASAP7_75t_L g2272 ( 
.A(n_2248),
.Y(n_2272)
);

NAND2xp5_ASAP7_75t_L g2273 ( 
.A(n_2251),
.B(n_153),
.Y(n_2273)
);

INVx1_ASAP7_75t_L g2274 ( 
.A(n_2248),
.Y(n_2274)
);

NOR2xp33_ASAP7_75t_L g2275 ( 
.A(n_2262),
.B(n_153),
.Y(n_2275)
);

AO22x2_ASAP7_75t_L g2276 ( 
.A1(n_2266),
.A2(n_2121),
.B1(n_156),
.B2(n_154),
.Y(n_2276)
);

AOI22xp5_ASAP7_75t_L g2277 ( 
.A1(n_2272),
.A2(n_2103),
.B1(n_2089),
.B2(n_1967),
.Y(n_2277)
);

OA21x2_ASAP7_75t_L g2278 ( 
.A1(n_2260),
.A2(n_2115),
.B(n_2114),
.Y(n_2278)
);

OR2x2_ASAP7_75t_L g2279 ( 
.A(n_2273),
.B(n_155),
.Y(n_2279)
);

NAND2x1_ASAP7_75t_SL g2280 ( 
.A(n_2274),
.B(n_155),
.Y(n_2280)
);

AOI21xp5_ASAP7_75t_L g2281 ( 
.A1(n_2263),
.A2(n_156),
.B(n_157),
.Y(n_2281)
);

INVx1_ASAP7_75t_L g2282 ( 
.A(n_2265),
.Y(n_2282)
);

NOR3xp33_ASAP7_75t_L g2283 ( 
.A(n_2261),
.B(n_2065),
.C(n_157),
.Y(n_2283)
);

NAND2xp5_ASAP7_75t_L g2284 ( 
.A(n_2261),
.B(n_158),
.Y(n_2284)
);

AOI211x1_ASAP7_75t_L g2285 ( 
.A1(n_2264),
.A2(n_160),
.B(n_158),
.C(n_159),
.Y(n_2285)
);

INVx1_ASAP7_75t_L g2286 ( 
.A(n_2271),
.Y(n_2286)
);

AOI22x1_ASAP7_75t_SL g2287 ( 
.A1(n_2267),
.A2(n_162),
.B1(n_160),
.B2(n_161),
.Y(n_2287)
);

AOI22xp5_ASAP7_75t_L g2288 ( 
.A1(n_2269),
.A2(n_2103),
.B1(n_2089),
.B2(n_2108),
.Y(n_2288)
);

AND2x4_ASAP7_75t_L g2289 ( 
.A(n_2282),
.B(n_2270),
.Y(n_2289)
);

OAI21xp5_ASAP7_75t_SL g2290 ( 
.A1(n_2275),
.A2(n_2268),
.B(n_161),
.Y(n_2290)
);

AOI22xp5_ASAP7_75t_L g2291 ( 
.A1(n_2283),
.A2(n_2108),
.B1(n_2074),
.B2(n_2018),
.Y(n_2291)
);

NAND4xp25_ASAP7_75t_L g2292 ( 
.A(n_2285),
.B(n_164),
.C(n_162),
.D(n_163),
.Y(n_2292)
);

NAND5xp2_ASAP7_75t_L g2293 ( 
.A(n_2286),
.B(n_2094),
.C(n_168),
.D(n_166),
.E(n_167),
.Y(n_2293)
);

NAND2x1_ASAP7_75t_L g2294 ( 
.A(n_2276),
.B(n_2108),
.Y(n_2294)
);

A2O1A1Ixp33_ASAP7_75t_L g2295 ( 
.A1(n_2280),
.A2(n_2281),
.B(n_2284),
.C(n_2279),
.Y(n_2295)
);

NOR2x1_ASAP7_75t_L g2296 ( 
.A(n_2287),
.B(n_166),
.Y(n_2296)
);

INVx1_ASAP7_75t_L g2297 ( 
.A(n_2276),
.Y(n_2297)
);

AOI22xp5_ASAP7_75t_L g2298 ( 
.A1(n_2288),
.A2(n_2074),
.B1(n_2018),
.B2(n_2158),
.Y(n_2298)
);

XNOR2xp5_ASAP7_75t_L g2299 ( 
.A(n_2278),
.B(n_167),
.Y(n_2299)
);

AOI221x1_ASAP7_75t_L g2300 ( 
.A1(n_2277),
.A2(n_170),
.B1(n_168),
.B2(n_169),
.C(n_171),
.Y(n_2300)
);

XOR2xp5_ASAP7_75t_L g2301 ( 
.A(n_2287),
.B(n_170),
.Y(n_2301)
);

INVx1_ASAP7_75t_L g2302 ( 
.A(n_2276),
.Y(n_2302)
);

NAND3xp33_ASAP7_75t_L g2303 ( 
.A(n_2275),
.B(n_171),
.C(n_172),
.Y(n_2303)
);

NOR3xp33_ASAP7_75t_L g2304 ( 
.A(n_2275),
.B(n_172),
.C(n_173),
.Y(n_2304)
);

INVx1_ASAP7_75t_L g2305 ( 
.A(n_2276),
.Y(n_2305)
);

OAI22xp5_ASAP7_75t_L g2306 ( 
.A1(n_2282),
.A2(n_1985),
.B1(n_1991),
.B2(n_2080),
.Y(n_2306)
);

INVx2_ASAP7_75t_SL g2307 ( 
.A(n_2280),
.Y(n_2307)
);

XOR2xp5_ASAP7_75t_L g2308 ( 
.A(n_2287),
.B(n_173),
.Y(n_2308)
);

OAI21xp33_ASAP7_75t_L g2309 ( 
.A1(n_2275),
.A2(n_2109),
.B(n_2101),
.Y(n_2309)
);

NAND2xp5_ASAP7_75t_L g2310 ( 
.A(n_2280),
.B(n_175),
.Y(n_2310)
);

INVx1_ASAP7_75t_L g2311 ( 
.A(n_2296),
.Y(n_2311)
);

INVx1_ASAP7_75t_L g2312 ( 
.A(n_2301),
.Y(n_2312)
);

INVx1_ASAP7_75t_L g2313 ( 
.A(n_2308),
.Y(n_2313)
);

AOI22xp5_ASAP7_75t_L g2314 ( 
.A1(n_2289),
.A2(n_2158),
.B1(n_2085),
.B2(n_2096),
.Y(n_2314)
);

NOR4xp25_ASAP7_75t_L g2315 ( 
.A(n_2307),
.B(n_178),
.C(n_176),
.D(n_177),
.Y(n_2315)
);

OAI22xp5_ASAP7_75t_L g2316 ( 
.A1(n_2289),
.A2(n_2085),
.B1(n_2008),
.B2(n_2162),
.Y(n_2316)
);

NAND2xp5_ASAP7_75t_L g2317 ( 
.A(n_2295),
.B(n_176),
.Y(n_2317)
);

INVx1_ASAP7_75t_L g2318 ( 
.A(n_2310),
.Y(n_2318)
);

OA22x2_ASAP7_75t_L g2319 ( 
.A1(n_2290),
.A2(n_2136),
.B1(n_2158),
.B2(n_2092),
.Y(n_2319)
);

INVx1_ASAP7_75t_L g2320 ( 
.A(n_2297),
.Y(n_2320)
);

INVx1_ASAP7_75t_L g2321 ( 
.A(n_2302),
.Y(n_2321)
);

NOR2xp33_ASAP7_75t_L g2322 ( 
.A(n_2293),
.B(n_177),
.Y(n_2322)
);

AOI22xp5_ASAP7_75t_L g2323 ( 
.A1(n_2305),
.A2(n_2162),
.B1(n_2165),
.B2(n_2136),
.Y(n_2323)
);

OA22x2_ASAP7_75t_L g2324 ( 
.A1(n_2300),
.A2(n_182),
.B1(n_179),
.B2(n_180),
.Y(n_2324)
);

AOI22xp5_ASAP7_75t_L g2325 ( 
.A1(n_2292),
.A2(n_2165),
.B1(n_1998),
.B2(n_2053),
.Y(n_2325)
);

NAND2xp5_ASAP7_75t_L g2326 ( 
.A(n_2304),
.B(n_182),
.Y(n_2326)
);

AOI22xp5_ASAP7_75t_L g2327 ( 
.A1(n_2291),
.A2(n_1998),
.B1(n_2061),
.B2(n_2062),
.Y(n_2327)
);

AOI22xp5_ASAP7_75t_L g2328 ( 
.A1(n_2294),
.A2(n_2088),
.B1(n_1992),
.B2(n_2071),
.Y(n_2328)
);

AOI31xp33_ASAP7_75t_L g2329 ( 
.A1(n_2303),
.A2(n_186),
.A3(n_184),
.B(n_185),
.Y(n_2329)
);

NAND2xp5_ASAP7_75t_L g2330 ( 
.A(n_2299),
.B(n_184),
.Y(n_2330)
);

INVx1_ASAP7_75t_L g2331 ( 
.A(n_2306),
.Y(n_2331)
);

HB1xp67_ASAP7_75t_L g2332 ( 
.A(n_2298),
.Y(n_2332)
);

AOI22xp5_ASAP7_75t_L g2333 ( 
.A1(n_2309),
.A2(n_1992),
.B1(n_2008),
.B2(n_2063),
.Y(n_2333)
);

INVx1_ASAP7_75t_L g2334 ( 
.A(n_2296),
.Y(n_2334)
);

AOI22xp5_ASAP7_75t_L g2335 ( 
.A1(n_2289),
.A2(n_2095),
.B1(n_2073),
.B2(n_2091),
.Y(n_2335)
);

NAND2xp5_ASAP7_75t_SL g2336 ( 
.A(n_2289),
.B(n_186),
.Y(n_2336)
);

AOI31xp33_ASAP7_75t_L g2337 ( 
.A1(n_2307),
.A2(n_189),
.A3(n_187),
.B(n_188),
.Y(n_2337)
);

INVx2_ASAP7_75t_L g2338 ( 
.A(n_2296),
.Y(n_2338)
);

AOI22xp5_ASAP7_75t_L g2339 ( 
.A1(n_2289),
.A2(n_2095),
.B1(n_2073),
.B2(n_2110),
.Y(n_2339)
);

INVxp67_ASAP7_75t_SL g2340 ( 
.A(n_2296),
.Y(n_2340)
);

INVx3_ASAP7_75t_L g2341 ( 
.A(n_2289),
.Y(n_2341)
);

INVx1_ASAP7_75t_L g2342 ( 
.A(n_2296),
.Y(n_2342)
);

NAND2xp5_ASAP7_75t_L g2343 ( 
.A(n_2307),
.B(n_187),
.Y(n_2343)
);

AOI22xp5_ASAP7_75t_L g2344 ( 
.A1(n_2289),
.A2(n_2081),
.B1(n_2086),
.B2(n_2075),
.Y(n_2344)
);

AOI221xp5_ASAP7_75t_L g2345 ( 
.A1(n_2307),
.A2(n_188),
.B1(n_189),
.B2(n_190),
.C(n_191),
.Y(n_2345)
);

HB1xp67_ASAP7_75t_L g2346 ( 
.A(n_2341),
.Y(n_2346)
);

O2A1O1Ixp33_ASAP7_75t_L g2347 ( 
.A1(n_2340),
.A2(n_192),
.B(n_190),
.C(n_191),
.Y(n_2347)
);

NAND4xp25_ASAP7_75t_L g2348 ( 
.A(n_2322),
.B(n_195),
.C(n_192),
.D(n_194),
.Y(n_2348)
);

OAI322xp33_ASAP7_75t_L g2349 ( 
.A1(n_2311),
.A2(n_194),
.A3(n_195),
.B1(n_196),
.B2(n_197),
.C1(n_198),
.C2(n_199),
.Y(n_2349)
);

INVx1_ASAP7_75t_SL g2350 ( 
.A(n_2334),
.Y(n_2350)
);

AOI221xp5_ASAP7_75t_L g2351 ( 
.A1(n_2342),
.A2(n_2313),
.B1(n_2312),
.B2(n_2338),
.C(n_2321),
.Y(n_2351)
);

INVx1_ASAP7_75t_L g2352 ( 
.A(n_2324),
.Y(n_2352)
);

INVx1_ASAP7_75t_L g2353 ( 
.A(n_2337),
.Y(n_2353)
);

OAI211xp5_ASAP7_75t_SL g2354 ( 
.A1(n_2320),
.A2(n_198),
.B(n_196),
.C(n_197),
.Y(n_2354)
);

INVx1_ASAP7_75t_L g2355 ( 
.A(n_2336),
.Y(n_2355)
);

NAND2xp5_ASAP7_75t_L g2356 ( 
.A(n_2315),
.B(n_199),
.Y(n_2356)
);

NOR2xp33_ASAP7_75t_R g2357 ( 
.A(n_2343),
.B(n_200),
.Y(n_2357)
);

AOI22xp33_ASAP7_75t_SL g2358 ( 
.A1(n_2318),
.A2(n_203),
.B1(n_201),
.B2(n_202),
.Y(n_2358)
);

INVx1_ASAP7_75t_SL g2359 ( 
.A(n_2330),
.Y(n_2359)
);

NAND2xp5_ASAP7_75t_SL g2360 ( 
.A(n_2345),
.B(n_201),
.Y(n_2360)
);

NAND4xp25_ASAP7_75t_L g2361 ( 
.A(n_2317),
.B(n_204),
.C(n_202),
.D(n_203),
.Y(n_2361)
);

AOI22xp5_ASAP7_75t_L g2362 ( 
.A1(n_2327),
.A2(n_2086),
.B1(n_2081),
.B2(n_208),
.Y(n_2362)
);

NOR2xp67_ASAP7_75t_L g2363 ( 
.A(n_2326),
.B(n_205),
.Y(n_2363)
);

OAI221xp5_ASAP7_75t_L g2364 ( 
.A1(n_2328),
.A2(n_2329),
.B1(n_2332),
.B2(n_2333),
.C(n_2331),
.Y(n_2364)
);

INVx2_ASAP7_75t_L g2365 ( 
.A(n_2319),
.Y(n_2365)
);

AOI221xp5_ASAP7_75t_L g2366 ( 
.A1(n_2316),
.A2(n_205),
.B1(n_206),
.B2(n_208),
.C(n_209),
.Y(n_2366)
);

NAND4xp75_ASAP7_75t_L g2367 ( 
.A(n_2323),
.B(n_2314),
.C(n_2325),
.D(n_2335),
.Y(n_2367)
);

INVx1_ASAP7_75t_L g2368 ( 
.A(n_2344),
.Y(n_2368)
);

NAND2xp5_ASAP7_75t_L g2369 ( 
.A(n_2339),
.B(n_206),
.Y(n_2369)
);

INVx1_ASAP7_75t_SL g2370 ( 
.A(n_2341),
.Y(n_2370)
);

OAI322xp33_ASAP7_75t_L g2371 ( 
.A1(n_2311),
.A2(n_209),
.A3(n_210),
.B1(n_211),
.B2(n_212),
.C1(n_213),
.C2(n_214),
.Y(n_2371)
);

INVx2_ASAP7_75t_L g2372 ( 
.A(n_2341),
.Y(n_2372)
);

OAI221xp5_ASAP7_75t_SL g2373 ( 
.A1(n_2341),
.A2(n_210),
.B1(n_213),
.B2(n_214),
.C(n_215),
.Y(n_2373)
);

NOR2x1p5_ASAP7_75t_L g2374 ( 
.A(n_2341),
.B(n_215),
.Y(n_2374)
);

NOR2x1_ASAP7_75t_L g2375 ( 
.A(n_2372),
.B(n_216),
.Y(n_2375)
);

AND2x2_ASAP7_75t_L g2376 ( 
.A(n_2346),
.B(n_216),
.Y(n_2376)
);

INVx1_ASAP7_75t_L g2377 ( 
.A(n_2374),
.Y(n_2377)
);

INVx1_ASAP7_75t_L g2378 ( 
.A(n_2356),
.Y(n_2378)
);

AND2x2_ASAP7_75t_SL g2379 ( 
.A(n_2352),
.B(n_217),
.Y(n_2379)
);

OR2x2_ASAP7_75t_L g2380 ( 
.A(n_2370),
.B(n_217),
.Y(n_2380)
);

NAND4xp75_ASAP7_75t_L g2381 ( 
.A(n_2351),
.B(n_222),
.C(n_219),
.D(n_221),
.Y(n_2381)
);

AOI22xp5_ASAP7_75t_SL g2382 ( 
.A1(n_2350),
.A2(n_224),
.B1(n_222),
.B2(n_223),
.Y(n_2382)
);

INVx1_ASAP7_75t_L g2383 ( 
.A(n_2363),
.Y(n_2383)
);

XNOR2xp5_ASAP7_75t_L g2384 ( 
.A(n_2348),
.B(n_223),
.Y(n_2384)
);

AOI22xp33_ASAP7_75t_SL g2385 ( 
.A1(n_2365),
.A2(n_226),
.B1(n_224),
.B2(n_225),
.Y(n_2385)
);

INVx1_ASAP7_75t_L g2386 ( 
.A(n_2353),
.Y(n_2386)
);

NAND2xp5_ASAP7_75t_L g2387 ( 
.A(n_2359),
.B(n_226),
.Y(n_2387)
);

INVx1_ASAP7_75t_L g2388 ( 
.A(n_2355),
.Y(n_2388)
);

AND2x4_ASAP7_75t_L g2389 ( 
.A(n_2360),
.B(n_227),
.Y(n_2389)
);

HB1xp67_ASAP7_75t_L g2390 ( 
.A(n_2357),
.Y(n_2390)
);

AOI22xp5_ASAP7_75t_L g2391 ( 
.A1(n_2364),
.A2(n_229),
.B1(n_227),
.B2(n_228),
.Y(n_2391)
);

NOR2x1_ASAP7_75t_L g2392 ( 
.A(n_2349),
.B(n_228),
.Y(n_2392)
);

NAND3xp33_ASAP7_75t_SL g2393 ( 
.A(n_2347),
.B(n_2358),
.C(n_2366),
.Y(n_2393)
);

INVx1_ASAP7_75t_L g2394 ( 
.A(n_2354),
.Y(n_2394)
);

OR2x2_ASAP7_75t_L g2395 ( 
.A(n_2361),
.B(n_229),
.Y(n_2395)
);

NAND4xp75_ASAP7_75t_L g2396 ( 
.A(n_2368),
.B(n_2369),
.C(n_2362),
.D(n_2373),
.Y(n_2396)
);

XNOR2xp5_ASAP7_75t_L g2397 ( 
.A(n_2367),
.B(n_230),
.Y(n_2397)
);

AND3x4_ASAP7_75t_L g2398 ( 
.A(n_2371),
.B(n_231),
.C(n_232),
.Y(n_2398)
);

INVx2_ASAP7_75t_L g2399 ( 
.A(n_2374),
.Y(n_2399)
);

O2A1O1Ixp33_ASAP7_75t_L g2400 ( 
.A1(n_2346),
.A2(n_234),
.B(n_231),
.C(n_233),
.Y(n_2400)
);

INVx1_ASAP7_75t_L g2401 ( 
.A(n_2346),
.Y(n_2401)
);

AOI22xp5_ASAP7_75t_L g2402 ( 
.A1(n_2350),
.A2(n_235),
.B1(n_233),
.B2(n_234),
.Y(n_2402)
);

INVx1_ASAP7_75t_L g2403 ( 
.A(n_2346),
.Y(n_2403)
);

NOR2x1_ASAP7_75t_L g2404 ( 
.A(n_2372),
.B(n_236),
.Y(n_2404)
);

INVx2_ASAP7_75t_L g2405 ( 
.A(n_2374),
.Y(n_2405)
);

INVxp67_ASAP7_75t_L g2406 ( 
.A(n_2346),
.Y(n_2406)
);

XNOR2xp5_ASAP7_75t_L g2407 ( 
.A(n_2346),
.B(n_236),
.Y(n_2407)
);

NOR2x1_ASAP7_75t_L g2408 ( 
.A(n_2372),
.B(n_237),
.Y(n_2408)
);

INVx1_ASAP7_75t_L g2409 ( 
.A(n_2346),
.Y(n_2409)
);

AOI22xp5_ASAP7_75t_L g2410 ( 
.A1(n_2350),
.A2(n_239),
.B1(n_237),
.B2(n_238),
.Y(n_2410)
);

INVx1_ASAP7_75t_L g2411 ( 
.A(n_2346),
.Y(n_2411)
);

AOI221xp5_ASAP7_75t_SL g2412 ( 
.A1(n_2406),
.A2(n_239),
.B1(n_240),
.B2(n_241),
.C(n_242),
.Y(n_2412)
);

OAI322xp33_ASAP7_75t_L g2413 ( 
.A1(n_2401),
.A2(n_243),
.A3(n_244),
.B1(n_245),
.B2(n_246),
.C1(n_247),
.C2(n_248),
.Y(n_2413)
);

NOR5xp2_ASAP7_75t_L g2414 ( 
.A(n_2403),
.B(n_244),
.C(n_245),
.D(n_246),
.E(n_247),
.Y(n_2414)
);

OAI211xp5_ASAP7_75t_L g2415 ( 
.A1(n_2409),
.A2(n_248),
.B(n_249),
.C(n_250),
.Y(n_2415)
);

NAND2xp5_ASAP7_75t_SL g2416 ( 
.A(n_2411),
.B(n_249),
.Y(n_2416)
);

OAI22xp33_ASAP7_75t_SL g2417 ( 
.A1(n_2378),
.A2(n_251),
.B1(n_252),
.B2(n_253),
.Y(n_2417)
);

OAI221xp5_ASAP7_75t_L g2418 ( 
.A1(n_2385),
.A2(n_253),
.B1(n_254),
.B2(n_255),
.C(n_256),
.Y(n_2418)
);

NAND4xp75_ASAP7_75t_L g2419 ( 
.A(n_2379),
.B(n_255),
.C(n_256),
.D(n_257),
.Y(n_2419)
);

NAND3xp33_ASAP7_75t_SL g2420 ( 
.A(n_2377),
.B(n_257),
.C(n_258),
.Y(n_2420)
);

AOI22x1_ASAP7_75t_SL g2421 ( 
.A1(n_2386),
.A2(n_258),
.B1(n_259),
.B2(n_260),
.Y(n_2421)
);

NOR4xp25_ASAP7_75t_L g2422 ( 
.A(n_2388),
.B(n_2405),
.C(n_2399),
.D(n_2383),
.Y(n_2422)
);

AOI211xp5_ASAP7_75t_L g2423 ( 
.A1(n_2400),
.A2(n_259),
.B(n_260),
.C(n_261),
.Y(n_2423)
);

INVx2_ASAP7_75t_L g2424 ( 
.A(n_2375),
.Y(n_2424)
);

AOI221xp5_ASAP7_75t_L g2425 ( 
.A1(n_2393),
.A2(n_261),
.B1(n_262),
.B2(n_263),
.C(n_264),
.Y(n_2425)
);

AOI22xp33_ASAP7_75t_SL g2426 ( 
.A1(n_2390),
.A2(n_263),
.B1(n_264),
.B2(n_265),
.Y(n_2426)
);

OAI22xp5_ASAP7_75t_L g2427 ( 
.A1(n_2402),
.A2(n_265),
.B1(n_266),
.B2(n_267),
.Y(n_2427)
);

INVx1_ASAP7_75t_L g2428 ( 
.A(n_2404),
.Y(n_2428)
);

OR3x1_ASAP7_75t_L g2429 ( 
.A(n_2394),
.B(n_268),
.C(n_270),
.Y(n_2429)
);

AOI221xp5_ASAP7_75t_L g2430 ( 
.A1(n_2389),
.A2(n_268),
.B1(n_271),
.B2(n_272),
.C(n_273),
.Y(n_2430)
);

O2A1O1Ixp33_ASAP7_75t_L g2431 ( 
.A1(n_2387),
.A2(n_271),
.B(n_272),
.C(n_273),
.Y(n_2431)
);

OAI321xp33_ASAP7_75t_L g2432 ( 
.A1(n_2391),
.A2(n_274),
.A3(n_275),
.B1(n_276),
.B2(n_277),
.C(n_278),
.Y(n_2432)
);

OAI21xp5_ASAP7_75t_SL g2433 ( 
.A1(n_2397),
.A2(n_274),
.B(n_275),
.Y(n_2433)
);

CKINVDCx20_ASAP7_75t_R g2434 ( 
.A(n_2384),
.Y(n_2434)
);

AOI21xp5_ASAP7_75t_L g2435 ( 
.A1(n_2407),
.A2(n_278),
.B(n_280),
.Y(n_2435)
);

AOI221x1_ASAP7_75t_L g2436 ( 
.A1(n_2389),
.A2(n_280),
.B1(n_281),
.B2(n_282),
.C(n_283),
.Y(n_2436)
);

AOI22xp5_ASAP7_75t_L g2437 ( 
.A1(n_2398),
.A2(n_282),
.B1(n_284),
.B2(n_285),
.Y(n_2437)
);

AOI221xp5_ASAP7_75t_L g2438 ( 
.A1(n_2395),
.A2(n_284),
.B1(n_285),
.B2(n_286),
.C(n_287),
.Y(n_2438)
);

NOR3xp33_ASAP7_75t_L g2439 ( 
.A(n_2408),
.B(n_2380),
.C(n_2376),
.Y(n_2439)
);

AO22x2_ASAP7_75t_L g2440 ( 
.A1(n_2381),
.A2(n_286),
.B1(n_287),
.B2(n_288),
.Y(n_2440)
);

OAI21xp33_ASAP7_75t_L g2441 ( 
.A1(n_2392),
.A2(n_288),
.B(n_289),
.Y(n_2441)
);

OAI211xp5_ASAP7_75t_L g2442 ( 
.A1(n_2410),
.A2(n_367),
.B(n_368),
.C(n_369),
.Y(n_2442)
);

AOI221xp5_ASAP7_75t_L g2443 ( 
.A1(n_2382),
.A2(n_1926),
.B1(n_1912),
.B2(n_1897),
.C(n_376),
.Y(n_2443)
);

NAND3x1_ASAP7_75t_L g2444 ( 
.A(n_2439),
.B(n_2396),
.C(n_372),
.Y(n_2444)
);

OR2x6_ASAP7_75t_L g2445 ( 
.A(n_2424),
.B(n_373),
.Y(n_2445)
);

XNOR2x1_ASAP7_75t_L g2446 ( 
.A(n_2419),
.B(n_375),
.Y(n_2446)
);

INVx1_ASAP7_75t_L g2447 ( 
.A(n_2429),
.Y(n_2447)
);

INVx2_ASAP7_75t_L g2448 ( 
.A(n_2428),
.Y(n_2448)
);

NAND2xp5_ASAP7_75t_L g2449 ( 
.A(n_2422),
.B(n_1897),
.Y(n_2449)
);

NAND2xp5_ASAP7_75t_L g2450 ( 
.A(n_2433),
.B(n_1897),
.Y(n_2450)
);

XOR2xp5_ASAP7_75t_L g2451 ( 
.A(n_2434),
.B(n_378),
.Y(n_2451)
);

INVx1_ASAP7_75t_L g2452 ( 
.A(n_2421),
.Y(n_2452)
);

XNOR2xp5_ASAP7_75t_L g2453 ( 
.A(n_2437),
.B(n_379),
.Y(n_2453)
);

OR2x2_ASAP7_75t_L g2454 ( 
.A(n_2420),
.B(n_1912),
.Y(n_2454)
);

INVx1_ASAP7_75t_L g2455 ( 
.A(n_2440),
.Y(n_2455)
);

NAND4xp75_ASAP7_75t_L g2456 ( 
.A(n_2436),
.B(n_380),
.C(n_381),
.D(n_382),
.Y(n_2456)
);

OAI22xp5_ASAP7_75t_SL g2457 ( 
.A1(n_2426),
.A2(n_1926),
.B1(n_1912),
.B2(n_385),
.Y(n_2457)
);

BUFx2_ASAP7_75t_L g2458 ( 
.A(n_2440),
.Y(n_2458)
);

OR2x2_ASAP7_75t_L g2459 ( 
.A(n_2416),
.B(n_1926),
.Y(n_2459)
);

XNOR2x1_ASAP7_75t_L g2460 ( 
.A(n_2427),
.B(n_383),
.Y(n_2460)
);

INVx1_ASAP7_75t_L g2461 ( 
.A(n_2417),
.Y(n_2461)
);

AND2x4_ASAP7_75t_L g2462 ( 
.A(n_2435),
.B(n_384),
.Y(n_2462)
);

HB1xp67_ASAP7_75t_L g2463 ( 
.A(n_2412),
.Y(n_2463)
);

INVx2_ASAP7_75t_L g2464 ( 
.A(n_2418),
.Y(n_2464)
);

OA22x2_ASAP7_75t_L g2465 ( 
.A1(n_2441),
.A2(n_388),
.B1(n_389),
.B2(n_390),
.Y(n_2465)
);

AOI22xp5_ASAP7_75t_L g2466 ( 
.A1(n_2415),
.A2(n_391),
.B1(n_392),
.B2(n_396),
.Y(n_2466)
);

NAND2xp5_ASAP7_75t_L g2467 ( 
.A(n_2423),
.B(n_526),
.Y(n_2467)
);

INVx2_ASAP7_75t_L g2468 ( 
.A(n_2414),
.Y(n_2468)
);

NOR2xp67_ASAP7_75t_SL g2469 ( 
.A(n_2442),
.B(n_397),
.Y(n_2469)
);

AOI22xp33_ASAP7_75t_L g2470 ( 
.A1(n_2438),
.A2(n_399),
.B1(n_401),
.B2(n_404),
.Y(n_2470)
);

NAND3xp33_ASAP7_75t_L g2471 ( 
.A(n_2425),
.B(n_405),
.C(n_406),
.Y(n_2471)
);

AND2x2_ASAP7_75t_SL g2472 ( 
.A(n_2430),
.B(n_408),
.Y(n_2472)
);

NAND4xp25_ASAP7_75t_L g2473 ( 
.A(n_2431),
.B(n_410),
.C(n_411),
.D(n_412),
.Y(n_2473)
);

CKINVDCx5p33_ASAP7_75t_R g2474 ( 
.A(n_2432),
.Y(n_2474)
);

INVx1_ASAP7_75t_L g2475 ( 
.A(n_2413),
.Y(n_2475)
);

AOI22xp5_ASAP7_75t_L g2476 ( 
.A1(n_2448),
.A2(n_2443),
.B1(n_415),
.B2(n_416),
.Y(n_2476)
);

CKINVDCx5p33_ASAP7_75t_R g2477 ( 
.A(n_2458),
.Y(n_2477)
);

OA21x2_ASAP7_75t_L g2478 ( 
.A1(n_2452),
.A2(n_413),
.B(n_418),
.Y(n_2478)
);

NOR2xp33_ASAP7_75t_L g2479 ( 
.A(n_2455),
.B(n_420),
.Y(n_2479)
);

BUFx4f_ASAP7_75t_SL g2480 ( 
.A(n_2447),
.Y(n_2480)
);

INVx1_ASAP7_75t_L g2481 ( 
.A(n_2444),
.Y(n_2481)
);

AOI22xp33_ASAP7_75t_L g2482 ( 
.A1(n_2468),
.A2(n_422),
.B1(n_423),
.B2(n_425),
.Y(n_2482)
);

NAND3x2_ASAP7_75t_L g2483 ( 
.A(n_2475),
.B(n_2461),
.C(n_2462),
.Y(n_2483)
);

INVx3_ASAP7_75t_SL g2484 ( 
.A(n_2474),
.Y(n_2484)
);

CKINVDCx5p33_ASAP7_75t_R g2485 ( 
.A(n_2463),
.Y(n_2485)
);

AND2x4_ASAP7_75t_L g2486 ( 
.A(n_2464),
.B(n_427),
.Y(n_2486)
);

CKINVDCx5p33_ASAP7_75t_R g2487 ( 
.A(n_2453),
.Y(n_2487)
);

CKINVDCx12_ASAP7_75t_R g2488 ( 
.A(n_2445),
.Y(n_2488)
);

OR2x6_ASAP7_75t_L g2489 ( 
.A(n_2467),
.B(n_429),
.Y(n_2489)
);

NAND2xp5_ASAP7_75t_SL g2490 ( 
.A(n_2466),
.B(n_434),
.Y(n_2490)
);

OAI221xp5_ASAP7_75t_L g2491 ( 
.A1(n_2449),
.A2(n_435),
.B1(n_436),
.B2(n_437),
.C(n_439),
.Y(n_2491)
);

INVx1_ASAP7_75t_L g2492 ( 
.A(n_2446),
.Y(n_2492)
);

AOI22xp5_ASAP7_75t_L g2493 ( 
.A1(n_2477),
.A2(n_2472),
.B1(n_2469),
.B2(n_2460),
.Y(n_2493)
);

INVx1_ASAP7_75t_L g2494 ( 
.A(n_2488),
.Y(n_2494)
);

AOI21xp33_ASAP7_75t_L g2495 ( 
.A1(n_2485),
.A2(n_2451),
.B(n_2445),
.Y(n_2495)
);

HB1xp67_ASAP7_75t_L g2496 ( 
.A(n_2480),
.Y(n_2496)
);

INVx1_ASAP7_75t_SL g2497 ( 
.A(n_2484),
.Y(n_2497)
);

INVx1_ASAP7_75t_L g2498 ( 
.A(n_2481),
.Y(n_2498)
);

AND2x2_ASAP7_75t_L g2499 ( 
.A(n_2489),
.B(n_2465),
.Y(n_2499)
);

NAND4xp75_ASAP7_75t_L g2500 ( 
.A(n_2492),
.B(n_2450),
.C(n_2456),
.D(n_2473),
.Y(n_2500)
);

OAI21xp5_ASAP7_75t_L g2501 ( 
.A1(n_2483),
.A2(n_2471),
.B(n_2491),
.Y(n_2501)
);

INVx1_ASAP7_75t_L g2502 ( 
.A(n_2489),
.Y(n_2502)
);

NAND2xp5_ASAP7_75t_L g2503 ( 
.A(n_2487),
.B(n_2470),
.Y(n_2503)
);

INVx3_ASAP7_75t_L g2504 ( 
.A(n_2486),
.Y(n_2504)
);

INVxp67_ASAP7_75t_L g2505 ( 
.A(n_2479),
.Y(n_2505)
);

INVx1_ASAP7_75t_L g2506 ( 
.A(n_2478),
.Y(n_2506)
);

AND2x2_ASAP7_75t_L g2507 ( 
.A(n_2476),
.B(n_2454),
.Y(n_2507)
);

AOI22xp33_ASAP7_75t_L g2508 ( 
.A1(n_2497),
.A2(n_2490),
.B1(n_2459),
.B2(n_2457),
.Y(n_2508)
);

INVx2_ASAP7_75t_L g2509 ( 
.A(n_2506),
.Y(n_2509)
);

AOI22xp5_ASAP7_75t_L g2510 ( 
.A1(n_2496),
.A2(n_2482),
.B1(n_441),
.B2(n_442),
.Y(n_2510)
);

INVx1_ASAP7_75t_L g2511 ( 
.A(n_2504),
.Y(n_2511)
);

INVx1_ASAP7_75t_L g2512 ( 
.A(n_2502),
.Y(n_2512)
);

OAI321xp33_ASAP7_75t_L g2513 ( 
.A1(n_2494),
.A2(n_440),
.A3(n_443),
.B1(n_445),
.B2(n_446),
.C(n_447),
.Y(n_2513)
);

XOR2xp5_ASAP7_75t_L g2514 ( 
.A(n_2493),
.B(n_448),
.Y(n_2514)
);

INVx1_ASAP7_75t_L g2515 ( 
.A(n_2499),
.Y(n_2515)
);

AOI22xp33_ASAP7_75t_L g2516 ( 
.A1(n_2509),
.A2(n_2495),
.B1(n_2498),
.B2(n_2505),
.Y(n_2516)
);

AOI221xp5_ASAP7_75t_L g2517 ( 
.A1(n_2511),
.A2(n_2501),
.B1(n_2507),
.B2(n_2503),
.C(n_2500),
.Y(n_2517)
);

OAI22xp33_ASAP7_75t_L g2518 ( 
.A1(n_2515),
.A2(n_455),
.B1(n_457),
.B2(n_458),
.Y(n_2518)
);

INVx1_ASAP7_75t_L g2519 ( 
.A(n_2516),
.Y(n_2519)
);

CKINVDCx20_ASAP7_75t_R g2520 ( 
.A(n_2517),
.Y(n_2520)
);

INVx1_ASAP7_75t_L g2521 ( 
.A(n_2518),
.Y(n_2521)
);

OAI222xp33_ASAP7_75t_L g2522 ( 
.A1(n_2519),
.A2(n_2512),
.B1(n_2508),
.B2(n_2514),
.C1(n_2510),
.C2(n_2513),
.Y(n_2522)
);

OAI222xp33_ASAP7_75t_L g2523 ( 
.A1(n_2520),
.A2(n_459),
.B1(n_460),
.B2(n_462),
.C1(n_463),
.C2(n_464),
.Y(n_2523)
);

AOI222xp33_ASAP7_75t_SL g2524 ( 
.A1(n_2521),
.A2(n_466),
.B1(n_468),
.B2(n_470),
.C1(n_471),
.C2(n_472),
.Y(n_2524)
);

AOI21xp5_ASAP7_75t_L g2525 ( 
.A1(n_2519),
.A2(n_474),
.B(n_475),
.Y(n_2525)
);

INVxp67_ASAP7_75t_SL g2526 ( 
.A(n_2522),
.Y(n_2526)
);

INVx1_ASAP7_75t_L g2527 ( 
.A(n_2525),
.Y(n_2527)
);

NAND2xp5_ASAP7_75t_L g2528 ( 
.A(n_2526),
.B(n_2524),
.Y(n_2528)
);

OAI22xp5_ASAP7_75t_SL g2529 ( 
.A1(n_2528),
.A2(n_2527),
.B1(n_2523),
.B2(n_478),
.Y(n_2529)
);

NAND2xp5_ASAP7_75t_L g2530 ( 
.A(n_2529),
.B(n_476),
.Y(n_2530)
);

AOI21xp5_ASAP7_75t_L g2531 ( 
.A1(n_2530),
.A2(n_477),
.B(n_479),
.Y(n_2531)
);

AOI211xp5_ASAP7_75t_L g2532 ( 
.A1(n_2531),
.A2(n_480),
.B(n_481),
.C(n_482),
.Y(n_2532)
);


endmodule