module fake_ariane_2657_n_1019 (n_83, n_8, n_56, n_60, n_170, n_190, n_160, n_64, n_179, n_180, n_119, n_124, n_167, n_90, n_195, n_38, n_213, n_47, n_110, n_153, n_18, n_197, n_86, n_75, n_89, n_67, n_176, n_149, n_34, n_158, n_172, n_69, n_95, n_175, n_92, n_143, n_183, n_203, n_150, n_98, n_74, n_113, n_114, n_33, n_19, n_40, n_181, n_152, n_120, n_169, n_106, n_12, n_53, n_173, n_111, n_21, n_115, n_133, n_66, n_205, n_71, n_24, n_7, n_109, n_208, n_96, n_156, n_209, n_49, n_20, n_174, n_100, n_17, n_50, n_187, n_132, n_62, n_210, n_147, n_204, n_200, n_51, n_166, n_76, n_218, n_103, n_79, n_26, n_3, n_46, n_220, n_0, n_84, n_36, n_199, n_91, n_159, n_107, n_189, n_72, n_105, n_128, n_217, n_44, n_30, n_82, n_178, n_31, n_42, n_57, n_131, n_201, n_70, n_10, n_117, n_139, n_165, n_85, n_130, n_144, n_6, n_214, n_48, n_94, n_101, n_4, n_134, n_188, n_185, n_2, n_32, n_37, n_58, n_65, n_123, n_212, n_9, n_138, n_112, n_45, n_162, n_11, n_129, n_126, n_137, n_122, n_198, n_148, n_164, n_52, n_157, n_184, n_177, n_135, n_73, n_77, n_171, n_15, n_118, n_93, n_121, n_23, n_61, n_108, n_102, n_182, n_196, n_125, n_22, n_168, n_43, n_1, n_81, n_87, n_206, n_13, n_27, n_207, n_29, n_41, n_219, n_140, n_55, n_191, n_151, n_136, n_192, n_28, n_80, n_146, n_211, n_194, n_97, n_154, n_215, n_142, n_161, n_14, n_163, n_88, n_186, n_141, n_68, n_116, n_104, n_202, n_145, n_78, n_193, n_39, n_59, n_63, n_99, n_216, n_16, n_5, n_155, n_127, n_35, n_54, n_25, n_1019);

input n_83;
input n_8;
input n_56;
input n_60;
input n_170;
input n_190;
input n_160;
input n_64;
input n_179;
input n_180;
input n_119;
input n_124;
input n_167;
input n_90;
input n_195;
input n_38;
input n_213;
input n_47;
input n_110;
input n_153;
input n_18;
input n_197;
input n_86;
input n_75;
input n_89;
input n_67;
input n_176;
input n_149;
input n_34;
input n_158;
input n_172;
input n_69;
input n_95;
input n_175;
input n_92;
input n_143;
input n_183;
input n_203;
input n_150;
input n_98;
input n_74;
input n_113;
input n_114;
input n_33;
input n_19;
input n_40;
input n_181;
input n_152;
input n_120;
input n_169;
input n_106;
input n_12;
input n_53;
input n_173;
input n_111;
input n_21;
input n_115;
input n_133;
input n_66;
input n_205;
input n_71;
input n_24;
input n_7;
input n_109;
input n_208;
input n_96;
input n_156;
input n_209;
input n_49;
input n_20;
input n_174;
input n_100;
input n_17;
input n_50;
input n_187;
input n_132;
input n_62;
input n_210;
input n_147;
input n_204;
input n_200;
input n_51;
input n_166;
input n_76;
input n_218;
input n_103;
input n_79;
input n_26;
input n_3;
input n_46;
input n_220;
input n_0;
input n_84;
input n_36;
input n_199;
input n_91;
input n_159;
input n_107;
input n_189;
input n_72;
input n_105;
input n_128;
input n_217;
input n_44;
input n_30;
input n_82;
input n_178;
input n_31;
input n_42;
input n_57;
input n_131;
input n_201;
input n_70;
input n_10;
input n_117;
input n_139;
input n_165;
input n_85;
input n_130;
input n_144;
input n_6;
input n_214;
input n_48;
input n_94;
input n_101;
input n_4;
input n_134;
input n_188;
input n_185;
input n_2;
input n_32;
input n_37;
input n_58;
input n_65;
input n_123;
input n_212;
input n_9;
input n_138;
input n_112;
input n_45;
input n_162;
input n_11;
input n_129;
input n_126;
input n_137;
input n_122;
input n_198;
input n_148;
input n_164;
input n_52;
input n_157;
input n_184;
input n_177;
input n_135;
input n_73;
input n_77;
input n_171;
input n_15;
input n_118;
input n_93;
input n_121;
input n_23;
input n_61;
input n_108;
input n_102;
input n_182;
input n_196;
input n_125;
input n_22;
input n_168;
input n_43;
input n_1;
input n_81;
input n_87;
input n_206;
input n_13;
input n_27;
input n_207;
input n_29;
input n_41;
input n_219;
input n_140;
input n_55;
input n_191;
input n_151;
input n_136;
input n_192;
input n_28;
input n_80;
input n_146;
input n_211;
input n_194;
input n_97;
input n_154;
input n_215;
input n_142;
input n_161;
input n_14;
input n_163;
input n_88;
input n_186;
input n_141;
input n_68;
input n_116;
input n_104;
input n_202;
input n_145;
input n_78;
input n_193;
input n_39;
input n_59;
input n_63;
input n_99;
input n_216;
input n_16;
input n_5;
input n_155;
input n_127;
input n_35;
input n_54;
input n_25;

output n_1019;

wire n_295;
wire n_356;
wire n_556;
wire n_698;
wire n_695;
wire n_913;
wire n_730;
wire n_386;
wire n_307;
wire n_516;
wire n_589;
wire n_332;
wire n_1008;
wire n_581;
wire n_294;
wire n_646;
wire n_640;
wire n_463;
wire n_830;
wire n_691;
wire n_404;
wire n_943;
wire n_678;
wire n_651;
wire n_987;
wire n_936;
wire n_347;
wire n_423;
wire n_961;
wire n_469;
wire n_479;
wire n_726;
wire n_603;
wire n_878;
wire n_373;
wire n_299;
wire n_836;
wire n_541;
wire n_499;
wire n_789;
wire n_788;
wire n_850;
wire n_908;
wire n_771;
wire n_564;
wire n_610;
wire n_752;
wire n_341;
wire n_985;
wire n_245;
wire n_421;
wire n_549;
wire n_522;
wire n_319;
wire n_591;
wire n_760;
wire n_690;
wire n_906;
wire n_416;
wire n_969;
wire n_283;
wire n_919;
wire n_525;
wire n_806;
wire n_367;
wire n_970;
wire n_713;
wire n_649;
wire n_598;
wire n_345;
wire n_374;
wire n_318;
wire n_817;
wire n_244;
wire n_643;
wire n_679;
wire n_226;
wire n_924;
wire n_927;
wire n_781;
wire n_261;
wire n_682;
wire n_663;
wire n_370;
wire n_706;
wire n_819;
wire n_717;
wire n_443;
wire n_286;
wire n_586;
wire n_864;
wire n_952;
wire n_686;
wire n_605;
wire n_776;
wire n_424;
wire n_584;
wire n_528;
wire n_387;
wire n_406;
wire n_826;
wire n_524;
wire n_349;
wire n_391;
wire n_634;
wire n_466;
wire n_756;
wire n_940;
wire n_346;
wire n_1016;
wire n_764;
wire n_979;
wire n_348;
wire n_552;
wire n_462;
wire n_607;
wire n_670;
wire n_897;
wire n_949;
wire n_956;
wire n_410;
wire n_445;
wire n_379;
wire n_515;
wire n_807;
wire n_765;
wire n_264;
wire n_891;
wire n_737;
wire n_885;
wire n_232;
wire n_441;
wire n_568;
wire n_385;
wire n_637;
wire n_917;
wire n_327;
wire n_766;
wire n_372;
wire n_377;
wire n_396;
wire n_802;
wire n_631;
wire n_399;
wire n_554;
wire n_960;
wire n_520;
wire n_980;
wire n_870;
wire n_714;
wire n_279;
wire n_945;
wire n_702;
wire n_958;
wire n_905;
wire n_790;
wire n_898;
wire n_857;
wire n_363;
wire n_720;
wire n_968;
wire n_354;
wire n_813;
wire n_926;
wire n_725;
wire n_419;
wire n_1009;
wire n_230;
wire n_270;
wire n_633;
wire n_900;
wire n_883;
wire n_338;
wire n_995;
wire n_285;
wire n_473;
wire n_801;
wire n_733;
wire n_761;
wire n_818;
wire n_500;
wire n_665;
wire n_336;
wire n_754;
wire n_731;
wire n_903;
wire n_871;
wire n_315;
wire n_779;
wire n_594;
wire n_311;
wire n_239;
wire n_402;
wire n_272;
wire n_829;
wire n_668;
wire n_339;
wire n_738;
wire n_758;
wire n_833;
wire n_672;
wire n_487;
wire n_740;
wire n_879;
wire n_422;
wire n_648;
wire n_784;
wire n_269;
wire n_597;
wire n_816;
wire n_1018;
wire n_855;
wire n_259;
wire n_835;
wire n_953;
wire n_808;
wire n_446;
wire n_553;
wire n_753;
wire n_566;
wire n_814;
wire n_578;
wire n_701;
wire n_1003;
wire n_625;
wire n_405;
wire n_557;
wire n_858;
wire n_242;
wire n_645;
wire n_989;
wire n_320;
wire n_331;
wire n_309;
wire n_559;
wire n_401;
wire n_485;
wire n_267;
wire n_495;
wire n_504;
wire n_647;
wire n_483;
wire n_335;
wire n_435;
wire n_350;
wire n_291;
wire n_822;
wire n_344;
wire n_381;
wire n_840;
wire n_426;
wire n_481;
wire n_433;
wire n_600;
wire n_721;
wire n_795;
wire n_398;
wire n_529;
wire n_502;
wire n_253;
wire n_561;
wire n_821;
wire n_770;
wire n_839;
wire n_928;
wire n_271;
wire n_465;
wire n_486;
wire n_507;
wire n_901;
wire n_759;
wire n_247;
wire n_569;
wire n_567;
wire n_825;
wire n_732;
wire n_971;
wire n_240;
wire n_369;
wire n_224;
wire n_787;
wire n_894;
wire n_547;
wire n_420;
wire n_562;
wire n_518;
wire n_439;
wire n_604;
wire n_614;
wire n_677;
wire n_222;
wire n_478;
wire n_703;
wire n_748;
wire n_786;
wire n_510;
wire n_831;
wire n_256;
wire n_868;
wire n_326;
wire n_681;
wire n_778;
wire n_227;
wire n_874;
wire n_323;
wire n_550;
wire n_988;
wire n_635;
wire n_707;
wire n_997;
wire n_330;
wire n_914;
wire n_400;
wire n_689;
wire n_694;
wire n_884;
wire n_983;
wire n_282;
wire n_328;
wire n_368;
wire n_590;
wire n_699;
wire n_727;
wire n_301;
wire n_248;
wire n_277;
wire n_467;
wire n_432;
wire n_545;
wire n_1015;
wire n_536;
wire n_644;
wire n_293;
wire n_823;
wire n_921;
wire n_620;
wire n_228;
wire n_325;
wire n_276;
wire n_688;
wire n_859;
wire n_636;
wire n_427;
wire n_587;
wire n_497;
wire n_693;
wire n_863;
wire n_303;
wire n_671;
wire n_442;
wire n_777;
wire n_929;
wire n_352;
wire n_538;
wire n_920;
wire n_899;
wire n_576;
wire n_843;
wire n_511;
wire n_611;
wire n_238;
wire n_365;
wire n_429;
wire n_455;
wire n_654;
wire n_588;
wire n_1013;
wire n_986;
wire n_638;
wire n_334;
wire n_729;
wire n_887;
wire n_661;
wire n_488;
wire n_775;
wire n_667;
wire n_300;
wire n_533;
wire n_904;
wire n_505;
wire n_869;
wire n_846;
wire n_390;
wire n_498;
wire n_501;
wire n_438;
wire n_314;
wire n_684;
wire n_440;
wire n_627;
wire n_273;
wire n_305;
wire n_539;
wire n_312;
wire n_233;
wire n_728;
wire n_388;
wire n_333;
wire n_449;
wire n_612;
wire n_413;
wire n_392;
wire n_376;
wire n_957;
wire n_977;
wire n_512;
wire n_715;
wire n_889;
wire n_935;
wire n_579;
wire n_844;
wire n_1012;
wire n_459;
wire n_685;
wire n_221;
wire n_321;
wire n_911;
wire n_361;
wire n_458;
wire n_383;
wire n_623;
wire n_838;
wire n_237;
wire n_861;
wire n_780;
wire n_950;
wire n_1017;
wire n_711;
wire n_877;
wire n_453;
wire n_734;
wire n_491;
wire n_810;
wire n_723;
wire n_616;
wire n_617;
wire n_658;
wire n_630;
wire n_705;
wire n_570;
wire n_362;
wire n_260;
wire n_543;
wire n_942;
wire n_310;
wire n_709;
wire n_236;
wire n_601;
wire n_683;
wire n_565;
wire n_281;
wire n_628;
wire n_809;
wire n_461;
wire n_490;
wire n_262;
wire n_743;
wire n_225;
wire n_907;
wire n_235;
wire n_1006;
wire n_881;
wire n_660;
wire n_464;
wire n_735;
wire n_575;
wire n_546;
wire n_297;
wire n_962;
wire n_662;
wire n_641;
wire n_1005;
wire n_503;
wire n_941;
wire n_700;
wire n_910;
wire n_290;
wire n_527;
wire n_741;
wire n_747;
wire n_772;
wire n_847;
wire n_939;
wire n_371;
wire n_845;
wire n_888;
wire n_918;
wire n_639;
wire n_452;
wire n_673;
wire n_676;
wire n_551;
wire n_308;
wire n_708;
wire n_417;
wire n_572;
wire n_343;
wire n_865;
wire n_414;
wire n_571;
wire n_680;
wire n_287;
wire n_302;
wire n_993;
wire n_380;
wire n_948;
wire n_582;
wire n_284;
wire n_922;
wire n_1004;
wire n_448;
wire n_593;
wire n_755;
wire n_710;
wire n_860;
wire n_249;
wire n_534;
wire n_355;
wire n_444;
wire n_609;
wire n_278;
wire n_851;
wire n_255;
wire n_560;
wire n_450;
wire n_890;
wire n_257;
wire n_842;
wire n_652;
wire n_451;
wire n_613;
wire n_745;
wire n_475;
wire n_896;
wire n_409;
wire n_947;
wire n_930;
wire n_519;
wire n_902;
wire n_384;
wire n_468;
wire n_853;
wire n_526;
wire n_716;
wire n_742;
wire n_696;
wire n_674;
wire n_482;
wire n_316;
wire n_798;
wire n_769;
wire n_820;
wire n_577;
wire n_407;
wire n_774;
wire n_872;
wire n_933;
wire n_916;
wire n_254;
wire n_596;
wire n_954;
wire n_912;
wire n_476;
wire n_460;
wire n_832;
wire n_535;
wire n_231;
wire n_366;
wire n_744;
wire n_762;
wire n_656;
wire n_555;
wire n_234;
wire n_492;
wire n_574;
wire n_848;
wire n_804;
wire n_280;
wire n_982;
wire n_915;
wire n_252;
wire n_629;
wire n_664;
wire n_454;
wire n_966;
wire n_992;
wire n_298;
wire n_955;
wire n_532;
wire n_415;
wire n_794;
wire n_763;
wire n_655;
wire n_544;
wire n_540;
wire n_692;
wire n_599;
wire n_768;
wire n_514;
wire n_418;
wire n_984;
wire n_537;
wire n_223;
wire n_403;
wire n_750;
wire n_834;
wire n_991;
wire n_389;
wire n_1007;
wire n_800;
wire n_657;
wire n_513;
wire n_837;
wire n_288;
wire n_812;
wire n_395;
wire n_621;
wire n_606;
wire n_951;
wire n_938;
wire n_895;
wire n_304;
wire n_862;
wire n_659;
wire n_583;
wire n_509;
wire n_1014;
wire n_724;
wire n_306;
wire n_666;
wire n_1000;
wire n_313;
wire n_430;
wire n_626;
wire n_493;
wire n_722;
wire n_378;
wire n_436;
wire n_946;
wire n_757;
wire n_375;
wire n_324;
wire n_585;
wire n_875;
wire n_669;
wire n_785;
wire n_827;
wire n_931;
wire n_619;
wire n_337;
wire n_437;
wire n_274;
wire n_622;
wire n_697;
wire n_967;
wire n_998;
wire n_999;
wire n_472;
wire n_937;
wire n_296;
wire n_265;
wire n_746;
wire n_456;
wire n_292;
wire n_880;
wire n_793;
wire n_852;
wire n_275;
wire n_704;
wire n_751;
wire n_615;
wire n_996;
wire n_521;
wire n_963;
wire n_873;
wire n_496;
wire n_739;
wire n_342;
wire n_866;
wire n_246;
wire n_517;
wire n_925;
wire n_530;
wire n_792;
wire n_1001;
wire n_824;
wire n_428;
wire n_1002;
wire n_358;
wire n_580;
wire n_892;
wire n_608;
wire n_959;
wire n_494;
wire n_719;
wire n_263;
wire n_434;
wire n_360;
wire n_975;
wire n_563;
wire n_229;
wire n_394;
wire n_923;
wire n_250;
wire n_932;
wire n_773;
wire n_981;
wire n_1010;
wire n_882;
wire n_990;
wire n_317;
wire n_867;
wire n_243;
wire n_803;
wire n_329;
wire n_718;
wire n_340;
wire n_944;
wire n_749;
wire n_994;
wire n_289;
wire n_548;
wire n_542;
wire n_815;
wire n_973;
wire n_523;
wire n_268;
wire n_972;
wire n_266;
wire n_470;
wire n_457;
wire n_632;
wire n_477;
wire n_364;
wire n_258;
wire n_650;
wire n_782;
wire n_856;
wire n_425;
wire n_431;
wire n_811;
wire n_508;
wire n_624;
wire n_791;
wire n_876;
wire n_618;
wire n_411;
wire n_484;
wire n_712;
wire n_849;
wire n_909;
wire n_976;
wire n_353;
wire n_736;
wire n_767;
wire n_241;
wire n_357;
wire n_412;
wire n_687;
wire n_447;
wire n_964;
wire n_382;
wire n_797;
wire n_489;
wire n_480;
wire n_978;
wire n_642;
wire n_1011;
wire n_408;
wire n_828;
wire n_595;
wire n_322;
wire n_251;
wire n_974;
wire n_506;
wire n_893;
wire n_602;
wire n_799;
wire n_558;
wire n_592;
wire n_397;
wire n_841;
wire n_854;
wire n_471;
wire n_351;
wire n_886;
wire n_965;
wire n_393;
wire n_474;
wire n_653;
wire n_359;
wire n_573;
wire n_796;
wire n_805;
wire n_531;
wire n_934;
wire n_783;
wire n_675;

INVx1_ASAP7_75t_L g221 ( 
.A(n_77),
.Y(n_221)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_200),
.Y(n_222)
);

HB1xp67_ASAP7_75t_L g223 ( 
.A(n_44),
.Y(n_223)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_101),
.Y(n_224)
);

CKINVDCx16_ASAP7_75t_R g225 ( 
.A(n_4),
.Y(n_225)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_79),
.Y(n_226)
);

CKINVDCx5p33_ASAP7_75t_R g227 ( 
.A(n_43),
.Y(n_227)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_31),
.Y(n_228)
);

CKINVDCx5p33_ASAP7_75t_R g229 ( 
.A(n_11),
.Y(n_229)
);

CKINVDCx5p33_ASAP7_75t_R g230 ( 
.A(n_164),
.Y(n_230)
);

CKINVDCx5p33_ASAP7_75t_R g231 ( 
.A(n_155),
.Y(n_231)
);

CKINVDCx5p33_ASAP7_75t_R g232 ( 
.A(n_207),
.Y(n_232)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_41),
.Y(n_233)
);

CKINVDCx5p33_ASAP7_75t_R g234 ( 
.A(n_16),
.Y(n_234)
);

CKINVDCx5p33_ASAP7_75t_R g235 ( 
.A(n_191),
.Y(n_235)
);

CKINVDCx5p33_ASAP7_75t_R g236 ( 
.A(n_13),
.Y(n_236)
);

CKINVDCx5p33_ASAP7_75t_R g237 ( 
.A(n_42),
.Y(n_237)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_56),
.Y(n_238)
);

INVx2_ASAP7_75t_L g239 ( 
.A(n_209),
.Y(n_239)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_63),
.Y(n_240)
);

CKINVDCx5p33_ASAP7_75t_R g241 ( 
.A(n_51),
.Y(n_241)
);

INVx2_ASAP7_75t_L g242 ( 
.A(n_9),
.Y(n_242)
);

BUFx3_ASAP7_75t_L g243 ( 
.A(n_71),
.Y(n_243)
);

BUFx2_ASAP7_75t_SL g244 ( 
.A(n_75),
.Y(n_244)
);

CKINVDCx5p33_ASAP7_75t_R g245 ( 
.A(n_98),
.Y(n_245)
);

CKINVDCx5p33_ASAP7_75t_R g246 ( 
.A(n_34),
.Y(n_246)
);

CKINVDCx5p33_ASAP7_75t_R g247 ( 
.A(n_66),
.Y(n_247)
);

CKINVDCx5p33_ASAP7_75t_R g248 ( 
.A(n_192),
.Y(n_248)
);

INVx2_ASAP7_75t_SL g249 ( 
.A(n_181),
.Y(n_249)
);

CKINVDCx20_ASAP7_75t_R g250 ( 
.A(n_24),
.Y(n_250)
);

CKINVDCx5p33_ASAP7_75t_R g251 ( 
.A(n_21),
.Y(n_251)
);

INVx2_ASAP7_75t_L g252 ( 
.A(n_172),
.Y(n_252)
);

CKINVDCx5p33_ASAP7_75t_R g253 ( 
.A(n_1),
.Y(n_253)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_78),
.Y(n_254)
);

INVx2_ASAP7_75t_SL g255 ( 
.A(n_60),
.Y(n_255)
);

CKINVDCx5p33_ASAP7_75t_R g256 ( 
.A(n_97),
.Y(n_256)
);

CKINVDCx5p33_ASAP7_75t_R g257 ( 
.A(n_133),
.Y(n_257)
);

INVx1_ASAP7_75t_SL g258 ( 
.A(n_95),
.Y(n_258)
);

INVx2_ASAP7_75t_L g259 ( 
.A(n_109),
.Y(n_259)
);

CKINVDCx5p33_ASAP7_75t_R g260 ( 
.A(n_139),
.Y(n_260)
);

CKINVDCx5p33_ASAP7_75t_R g261 ( 
.A(n_183),
.Y(n_261)
);

CKINVDCx5p33_ASAP7_75t_R g262 ( 
.A(n_130),
.Y(n_262)
);

CKINVDCx5p33_ASAP7_75t_R g263 ( 
.A(n_159),
.Y(n_263)
);

CKINVDCx5p33_ASAP7_75t_R g264 ( 
.A(n_173),
.Y(n_264)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_152),
.Y(n_265)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_49),
.Y(n_266)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_55),
.Y(n_267)
);

CKINVDCx5p33_ASAP7_75t_R g268 ( 
.A(n_212),
.Y(n_268)
);

CKINVDCx20_ASAP7_75t_R g269 ( 
.A(n_3),
.Y(n_269)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_89),
.Y(n_270)
);

CKINVDCx5p33_ASAP7_75t_R g271 ( 
.A(n_113),
.Y(n_271)
);

CKINVDCx5p33_ASAP7_75t_R g272 ( 
.A(n_33),
.Y(n_272)
);

CKINVDCx20_ASAP7_75t_R g273 ( 
.A(n_84),
.Y(n_273)
);

INVx2_ASAP7_75t_L g274 ( 
.A(n_197),
.Y(n_274)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_119),
.Y(n_275)
);

CKINVDCx5p33_ASAP7_75t_R g276 ( 
.A(n_120),
.Y(n_276)
);

CKINVDCx5p33_ASAP7_75t_R g277 ( 
.A(n_153),
.Y(n_277)
);

CKINVDCx5p33_ASAP7_75t_R g278 ( 
.A(n_132),
.Y(n_278)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_22),
.Y(n_279)
);

INVx2_ASAP7_75t_L g280 ( 
.A(n_81),
.Y(n_280)
);

BUFx5_ASAP7_75t_L g281 ( 
.A(n_187),
.Y(n_281)
);

BUFx10_ASAP7_75t_L g282 ( 
.A(n_111),
.Y(n_282)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_13),
.Y(n_283)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_21),
.Y(n_284)
);

CKINVDCx5p33_ASAP7_75t_R g285 ( 
.A(n_147),
.Y(n_285)
);

CKINVDCx5p33_ASAP7_75t_R g286 ( 
.A(n_126),
.Y(n_286)
);

CKINVDCx5p33_ASAP7_75t_R g287 ( 
.A(n_166),
.Y(n_287)
);

CKINVDCx5p33_ASAP7_75t_R g288 ( 
.A(n_12),
.Y(n_288)
);

CKINVDCx5p33_ASAP7_75t_R g289 ( 
.A(n_178),
.Y(n_289)
);

CKINVDCx20_ASAP7_75t_R g290 ( 
.A(n_215),
.Y(n_290)
);

CKINVDCx5p33_ASAP7_75t_R g291 ( 
.A(n_108),
.Y(n_291)
);

CKINVDCx5p33_ASAP7_75t_R g292 ( 
.A(n_28),
.Y(n_292)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_0),
.Y(n_293)
);

CKINVDCx5p33_ASAP7_75t_R g294 ( 
.A(n_72),
.Y(n_294)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_202),
.Y(n_295)
);

INVxp67_ASAP7_75t_SL g296 ( 
.A(n_134),
.Y(n_296)
);

CKINVDCx5p33_ASAP7_75t_R g297 ( 
.A(n_127),
.Y(n_297)
);

CKINVDCx5p33_ASAP7_75t_R g298 ( 
.A(n_190),
.Y(n_298)
);

CKINVDCx5p33_ASAP7_75t_R g299 ( 
.A(n_195),
.Y(n_299)
);

CKINVDCx5p33_ASAP7_75t_R g300 ( 
.A(n_35),
.Y(n_300)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_91),
.Y(n_301)
);

INVx1_ASAP7_75t_SL g302 ( 
.A(n_216),
.Y(n_302)
);

BUFx10_ASAP7_75t_L g303 ( 
.A(n_169),
.Y(n_303)
);

CKINVDCx5p33_ASAP7_75t_R g304 ( 
.A(n_143),
.Y(n_304)
);

CKINVDCx5p33_ASAP7_75t_R g305 ( 
.A(n_138),
.Y(n_305)
);

INVx2_ASAP7_75t_SL g306 ( 
.A(n_18),
.Y(n_306)
);

CKINVDCx5p33_ASAP7_75t_R g307 ( 
.A(n_196),
.Y(n_307)
);

CKINVDCx5p33_ASAP7_75t_R g308 ( 
.A(n_104),
.Y(n_308)
);

CKINVDCx5p33_ASAP7_75t_R g309 ( 
.A(n_194),
.Y(n_309)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_76),
.Y(n_310)
);

CKINVDCx5p33_ASAP7_75t_R g311 ( 
.A(n_3),
.Y(n_311)
);

CKINVDCx5p33_ASAP7_75t_R g312 ( 
.A(n_213),
.Y(n_312)
);

CKINVDCx5p33_ASAP7_75t_R g313 ( 
.A(n_4),
.Y(n_313)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_174),
.Y(n_314)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_228),
.Y(n_315)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_279),
.Y(n_316)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_283),
.Y(n_317)
);

CKINVDCx16_ASAP7_75t_R g318 ( 
.A(n_225),
.Y(n_318)
);

CKINVDCx5p33_ASAP7_75t_R g319 ( 
.A(n_229),
.Y(n_319)
);

CKINVDCx20_ASAP7_75t_R g320 ( 
.A(n_250),
.Y(n_320)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_284),
.Y(n_321)
);

CKINVDCx5p33_ASAP7_75t_R g322 ( 
.A(n_234),
.Y(n_322)
);

NOR2xp33_ASAP7_75t_L g323 ( 
.A(n_223),
.B(n_0),
.Y(n_323)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_293),
.Y(n_324)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_242),
.Y(n_325)
);

CKINVDCx20_ASAP7_75t_R g326 ( 
.A(n_250),
.Y(n_326)
);

INVxp33_ASAP7_75t_SL g327 ( 
.A(n_236),
.Y(n_327)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_242),
.Y(n_328)
);

CKINVDCx5p33_ASAP7_75t_R g329 ( 
.A(n_251),
.Y(n_329)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_306),
.Y(n_330)
);

CKINVDCx5p33_ASAP7_75t_R g331 ( 
.A(n_253),
.Y(n_331)
);

CKINVDCx20_ASAP7_75t_R g332 ( 
.A(n_273),
.Y(n_332)
);

INVxp33_ASAP7_75t_SL g333 ( 
.A(n_272),
.Y(n_333)
);

BUFx6f_ASAP7_75t_L g334 ( 
.A(n_243),
.Y(n_334)
);

CKINVDCx20_ASAP7_75t_R g335 ( 
.A(n_273),
.Y(n_335)
);

NOR2xp67_ASAP7_75t_L g336 ( 
.A(n_288),
.B(n_1),
.Y(n_336)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_282),
.Y(n_337)
);

CKINVDCx5p33_ASAP7_75t_R g338 ( 
.A(n_292),
.Y(n_338)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_282),
.Y(n_339)
);

NOR2xp33_ASAP7_75t_L g340 ( 
.A(n_314),
.B(n_2),
.Y(n_340)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_282),
.Y(n_341)
);

BUFx2_ASAP7_75t_L g342 ( 
.A(n_311),
.Y(n_342)
);

NOR2xp33_ASAP7_75t_L g343 ( 
.A(n_221),
.B(n_2),
.Y(n_343)
);

INVx2_ASAP7_75t_L g344 ( 
.A(n_243),
.Y(n_344)
);

CKINVDCx20_ASAP7_75t_R g345 ( 
.A(n_269),
.Y(n_345)
);

INVx1_ASAP7_75t_L g346 ( 
.A(n_303),
.Y(n_346)
);

CKINVDCx5p33_ASAP7_75t_R g347 ( 
.A(n_313),
.Y(n_347)
);

CKINVDCx20_ASAP7_75t_R g348 ( 
.A(n_269),
.Y(n_348)
);

INVxp67_ASAP7_75t_L g349 ( 
.A(n_303),
.Y(n_349)
);

INVxp67_ASAP7_75t_SL g350 ( 
.A(n_239),
.Y(n_350)
);

CKINVDCx5p33_ASAP7_75t_R g351 ( 
.A(n_227),
.Y(n_351)
);

CKINVDCx16_ASAP7_75t_R g352 ( 
.A(n_290),
.Y(n_352)
);

CKINVDCx5p33_ASAP7_75t_R g353 ( 
.A(n_230),
.Y(n_353)
);

INVx2_ASAP7_75t_L g354 ( 
.A(n_222),
.Y(n_354)
);

INVxp33_ASAP7_75t_SL g355 ( 
.A(n_244),
.Y(n_355)
);

INVx1_ASAP7_75t_L g356 ( 
.A(n_303),
.Y(n_356)
);

INVx2_ASAP7_75t_L g357 ( 
.A(n_224),
.Y(n_357)
);

INVxp33_ASAP7_75t_L g358 ( 
.A(n_239),
.Y(n_358)
);

CKINVDCx5p33_ASAP7_75t_R g359 ( 
.A(n_231),
.Y(n_359)
);

INVx1_ASAP7_75t_L g360 ( 
.A(n_226),
.Y(n_360)
);

CKINVDCx5p33_ASAP7_75t_R g361 ( 
.A(n_232),
.Y(n_361)
);

INVx1_ASAP7_75t_L g362 ( 
.A(n_233),
.Y(n_362)
);

CKINVDCx14_ASAP7_75t_R g363 ( 
.A(n_290),
.Y(n_363)
);

CKINVDCx20_ASAP7_75t_R g364 ( 
.A(n_235),
.Y(n_364)
);

CKINVDCx20_ASAP7_75t_R g365 ( 
.A(n_237),
.Y(n_365)
);

CKINVDCx5p33_ASAP7_75t_R g366 ( 
.A(n_241),
.Y(n_366)
);

INVx1_ASAP7_75t_L g367 ( 
.A(n_238),
.Y(n_367)
);

INVx1_ASAP7_75t_L g368 ( 
.A(n_240),
.Y(n_368)
);

INVx2_ASAP7_75t_L g369 ( 
.A(n_254),
.Y(n_369)
);

INVx1_ASAP7_75t_L g370 ( 
.A(n_265),
.Y(n_370)
);

NAND2xp5_ASAP7_75t_L g371 ( 
.A(n_266),
.B(n_5),
.Y(n_371)
);

NAND2xp5_ASAP7_75t_L g372 ( 
.A(n_337),
.B(n_339),
.Y(n_372)
);

HB1xp67_ASAP7_75t_L g373 ( 
.A(n_318),
.Y(n_373)
);

INVx1_ASAP7_75t_L g374 ( 
.A(n_354),
.Y(n_374)
);

INVx1_ASAP7_75t_L g375 ( 
.A(n_354),
.Y(n_375)
);

INVx2_ASAP7_75t_L g376 ( 
.A(n_357),
.Y(n_376)
);

INVx1_ASAP7_75t_L g377 ( 
.A(n_357),
.Y(n_377)
);

INVx3_ASAP7_75t_L g378 ( 
.A(n_369),
.Y(n_378)
);

INVx3_ASAP7_75t_L g379 ( 
.A(n_369),
.Y(n_379)
);

NAND2xp5_ASAP7_75t_L g380 ( 
.A(n_341),
.B(n_267),
.Y(n_380)
);

INVx2_ASAP7_75t_L g381 ( 
.A(n_344),
.Y(n_381)
);

INVx3_ASAP7_75t_L g382 ( 
.A(n_334),
.Y(n_382)
);

INVx2_ASAP7_75t_L g383 ( 
.A(n_344),
.Y(n_383)
);

INVx1_ASAP7_75t_L g384 ( 
.A(n_360),
.Y(n_384)
);

NAND3xp33_ASAP7_75t_L g385 ( 
.A(n_323),
.B(n_259),
.C(n_252),
.Y(n_385)
);

INVx1_ASAP7_75t_L g386 ( 
.A(n_362),
.Y(n_386)
);

INVx1_ASAP7_75t_L g387 ( 
.A(n_367),
.Y(n_387)
);

NAND2xp5_ASAP7_75t_SL g388 ( 
.A(n_351),
.B(n_252),
.Y(n_388)
);

INVx1_ASAP7_75t_L g389 ( 
.A(n_368),
.Y(n_389)
);

BUFx6f_ASAP7_75t_L g390 ( 
.A(n_334),
.Y(n_390)
);

CKINVDCx6p67_ASAP7_75t_R g391 ( 
.A(n_364),
.Y(n_391)
);

INVx1_ASAP7_75t_L g392 ( 
.A(n_370),
.Y(n_392)
);

BUFx6f_ASAP7_75t_L g393 ( 
.A(n_334),
.Y(n_393)
);

INVx2_ASAP7_75t_L g394 ( 
.A(n_334),
.Y(n_394)
);

NAND2xp5_ASAP7_75t_L g395 ( 
.A(n_346),
.B(n_270),
.Y(n_395)
);

INVx1_ASAP7_75t_L g396 ( 
.A(n_325),
.Y(n_396)
);

INVx1_ASAP7_75t_L g397 ( 
.A(n_328),
.Y(n_397)
);

INVx2_ASAP7_75t_L g398 ( 
.A(n_315),
.Y(n_398)
);

XOR2xp5_ASAP7_75t_L g399 ( 
.A(n_320),
.B(n_5),
.Y(n_399)
);

INVx1_ASAP7_75t_L g400 ( 
.A(n_350),
.Y(n_400)
);

INVx2_ASAP7_75t_L g401 ( 
.A(n_316),
.Y(n_401)
);

INVx2_ASAP7_75t_L g402 ( 
.A(n_317),
.Y(n_402)
);

INVx2_ASAP7_75t_L g403 ( 
.A(n_321),
.Y(n_403)
);

NAND3xp33_ASAP7_75t_L g404 ( 
.A(n_319),
.B(n_274),
.C(n_259),
.Y(n_404)
);

NAND2xp5_ASAP7_75t_SL g405 ( 
.A(n_353),
.B(n_274),
.Y(n_405)
);

INVx1_ASAP7_75t_L g406 ( 
.A(n_371),
.Y(n_406)
);

INVx1_ASAP7_75t_L g407 ( 
.A(n_324),
.Y(n_407)
);

INVx1_ASAP7_75t_L g408 ( 
.A(n_340),
.Y(n_408)
);

INVx3_ASAP7_75t_L g409 ( 
.A(n_330),
.Y(n_409)
);

INVx2_ASAP7_75t_L g410 ( 
.A(n_343),
.Y(n_410)
);

INVx1_ASAP7_75t_L g411 ( 
.A(n_358),
.Y(n_411)
);

NOR2xp33_ASAP7_75t_L g412 ( 
.A(n_355),
.B(n_275),
.Y(n_412)
);

INVx1_ASAP7_75t_L g413 ( 
.A(n_358),
.Y(n_413)
);

INVx1_ASAP7_75t_L g414 ( 
.A(n_356),
.Y(n_414)
);

NAND2xp33_ASAP7_75t_SL g415 ( 
.A(n_364),
.B(n_249),
.Y(n_415)
);

OAI22xp5_ASAP7_75t_L g416 ( 
.A1(n_349),
.A2(n_296),
.B1(n_310),
.B2(n_295),
.Y(n_416)
);

NOR2xp33_ASAP7_75t_L g417 ( 
.A(n_366),
.B(n_301),
.Y(n_417)
);

INVx2_ASAP7_75t_L g418 ( 
.A(n_359),
.Y(n_418)
);

BUFx6f_ASAP7_75t_L g419 ( 
.A(n_361),
.Y(n_419)
);

INVx2_ASAP7_75t_L g420 ( 
.A(n_342),
.Y(n_420)
);

INVx3_ASAP7_75t_L g421 ( 
.A(n_322),
.Y(n_421)
);

NAND2xp5_ASAP7_75t_L g422 ( 
.A(n_329),
.B(n_255),
.Y(n_422)
);

INVx1_ASAP7_75t_L g423 ( 
.A(n_336),
.Y(n_423)
);

INVx1_ASAP7_75t_L g424 ( 
.A(n_331),
.Y(n_424)
);

BUFx6f_ASAP7_75t_L g425 ( 
.A(n_338),
.Y(n_425)
);

NOR2xp33_ASAP7_75t_L g426 ( 
.A(n_327),
.B(n_258),
.Y(n_426)
);

NAND2xp5_ASAP7_75t_L g427 ( 
.A(n_347),
.B(n_280),
.Y(n_427)
);

INVx2_ASAP7_75t_L g428 ( 
.A(n_365),
.Y(n_428)
);

INVx2_ASAP7_75t_L g429 ( 
.A(n_365),
.Y(n_429)
);

CKINVDCx5p33_ASAP7_75t_R g430 ( 
.A(n_391),
.Y(n_430)
);

OR2x6_ASAP7_75t_L g431 ( 
.A(n_373),
.B(n_363),
.Y(n_431)
);

AND2x2_ASAP7_75t_L g432 ( 
.A(n_411),
.B(n_363),
.Y(n_432)
);

NOR2xp33_ASAP7_75t_L g433 ( 
.A(n_411),
.B(n_333),
.Y(n_433)
);

NAND2x1p5_ASAP7_75t_L g434 ( 
.A(n_419),
.B(n_425),
.Y(n_434)
);

OR2x2_ASAP7_75t_L g435 ( 
.A(n_420),
.B(n_352),
.Y(n_435)
);

INVx1_ASAP7_75t_L g436 ( 
.A(n_398),
.Y(n_436)
);

OR2x2_ASAP7_75t_L g437 ( 
.A(n_420),
.B(n_332),
.Y(n_437)
);

OR2x2_ASAP7_75t_L g438 ( 
.A(n_413),
.B(n_335),
.Y(n_438)
);

NOR2xp33_ASAP7_75t_SL g439 ( 
.A(n_426),
.B(n_302),
.Y(n_439)
);

BUFx6f_ASAP7_75t_L g440 ( 
.A(n_390),
.Y(n_440)
);

OR2x2_ASAP7_75t_L g441 ( 
.A(n_413),
.B(n_428),
.Y(n_441)
);

INVx1_ASAP7_75t_L g442 ( 
.A(n_398),
.Y(n_442)
);

INVx2_ASAP7_75t_L g443 ( 
.A(n_382),
.Y(n_443)
);

BUFx6f_ASAP7_75t_L g444 ( 
.A(n_390),
.Y(n_444)
);

BUFx4f_ASAP7_75t_L g445 ( 
.A(n_425),
.Y(n_445)
);

INVx1_ASAP7_75t_L g446 ( 
.A(n_401),
.Y(n_446)
);

INVx1_ASAP7_75t_L g447 ( 
.A(n_401),
.Y(n_447)
);

NOR2xp33_ASAP7_75t_L g448 ( 
.A(n_414),
.B(n_280),
.Y(n_448)
);

OR2x2_ASAP7_75t_L g449 ( 
.A(n_428),
.B(n_320),
.Y(n_449)
);

INVx1_ASAP7_75t_L g450 ( 
.A(n_402),
.Y(n_450)
);

INVx1_ASAP7_75t_L g451 ( 
.A(n_402),
.Y(n_451)
);

INVx1_ASAP7_75t_L g452 ( 
.A(n_403),
.Y(n_452)
);

NAND2xp5_ASAP7_75t_SL g453 ( 
.A(n_419),
.B(n_245),
.Y(n_453)
);

INVx2_ASAP7_75t_L g454 ( 
.A(n_382),
.Y(n_454)
);

AND2x2_ASAP7_75t_L g455 ( 
.A(n_421),
.B(n_326),
.Y(n_455)
);

NAND2xp5_ASAP7_75t_L g456 ( 
.A(n_406),
.B(n_281),
.Y(n_456)
);

INVx1_ASAP7_75t_SL g457 ( 
.A(n_429),
.Y(n_457)
);

INVx2_ASAP7_75t_L g458 ( 
.A(n_382),
.Y(n_458)
);

BUFx3_ASAP7_75t_L g459 ( 
.A(n_425),
.Y(n_459)
);

INVx3_ASAP7_75t_L g460 ( 
.A(n_390),
.Y(n_460)
);

AND2x2_ASAP7_75t_SL g461 ( 
.A(n_425),
.B(n_6),
.Y(n_461)
);

INVx2_ASAP7_75t_L g462 ( 
.A(n_394),
.Y(n_462)
);

HB1xp67_ASAP7_75t_L g463 ( 
.A(n_429),
.Y(n_463)
);

AND2x4_ASAP7_75t_L g464 ( 
.A(n_414),
.B(n_6),
.Y(n_464)
);

INVx1_ASAP7_75t_L g465 ( 
.A(n_403),
.Y(n_465)
);

NAND2xp5_ASAP7_75t_L g466 ( 
.A(n_406),
.B(n_281),
.Y(n_466)
);

NAND2xp5_ASAP7_75t_L g467 ( 
.A(n_410),
.B(n_281),
.Y(n_467)
);

OAI22xp5_ASAP7_75t_SL g468 ( 
.A1(n_399),
.A2(n_348),
.B1(n_345),
.B2(n_326),
.Y(n_468)
);

NAND3xp33_ASAP7_75t_L g469 ( 
.A(n_412),
.B(n_247),
.C(n_246),
.Y(n_469)
);

NAND2xp5_ASAP7_75t_L g470 ( 
.A(n_410),
.B(n_281),
.Y(n_470)
);

NOR2xp33_ASAP7_75t_L g471 ( 
.A(n_372),
.B(n_248),
.Y(n_471)
);

BUFx6f_ASAP7_75t_L g472 ( 
.A(n_390),
.Y(n_472)
);

AND2x4_ASAP7_75t_L g473 ( 
.A(n_400),
.B(n_7),
.Y(n_473)
);

INVx1_ASAP7_75t_L g474 ( 
.A(n_384),
.Y(n_474)
);

AND2x4_ASAP7_75t_L g475 ( 
.A(n_400),
.B(n_7),
.Y(n_475)
);

INVx2_ASAP7_75t_L g476 ( 
.A(n_394),
.Y(n_476)
);

INVx1_ASAP7_75t_L g477 ( 
.A(n_384),
.Y(n_477)
);

BUFx10_ASAP7_75t_L g478 ( 
.A(n_419),
.Y(n_478)
);

BUFx6f_ASAP7_75t_L g479 ( 
.A(n_390),
.Y(n_479)
);

BUFx3_ASAP7_75t_L g480 ( 
.A(n_425),
.Y(n_480)
);

INVx1_ASAP7_75t_L g481 ( 
.A(n_386),
.Y(n_481)
);

NAND2xp5_ASAP7_75t_SL g482 ( 
.A(n_419),
.B(n_256),
.Y(n_482)
);

AND2x2_ASAP7_75t_L g483 ( 
.A(n_421),
.B(n_348),
.Y(n_483)
);

INVx3_ASAP7_75t_L g484 ( 
.A(n_393),
.Y(n_484)
);

INVx1_ASAP7_75t_L g485 ( 
.A(n_386),
.Y(n_485)
);

AOI22xp33_ASAP7_75t_L g486 ( 
.A1(n_408),
.A2(n_281),
.B1(n_312),
.B2(n_309),
.Y(n_486)
);

NAND2xp5_ASAP7_75t_L g487 ( 
.A(n_408),
.B(n_381),
.Y(n_487)
);

AND2x4_ASAP7_75t_L g488 ( 
.A(n_418),
.B(n_8),
.Y(n_488)
);

AOI22xp33_ASAP7_75t_L g489 ( 
.A1(n_385),
.A2(n_281),
.B1(n_308),
.B2(n_307),
.Y(n_489)
);

INVx2_ASAP7_75t_L g490 ( 
.A(n_381),
.Y(n_490)
);

AND2x2_ASAP7_75t_L g491 ( 
.A(n_421),
.B(n_424),
.Y(n_491)
);

AND2x2_ASAP7_75t_L g492 ( 
.A(n_424),
.B(n_345),
.Y(n_492)
);

NAND2xp5_ASAP7_75t_L g493 ( 
.A(n_383),
.B(n_376),
.Y(n_493)
);

NAND2xp5_ASAP7_75t_SL g494 ( 
.A(n_419),
.B(n_257),
.Y(n_494)
);

INVx1_ASAP7_75t_L g495 ( 
.A(n_387),
.Y(n_495)
);

INVx2_ASAP7_75t_L g496 ( 
.A(n_383),
.Y(n_496)
);

CKINVDCx5p33_ASAP7_75t_R g497 ( 
.A(n_391),
.Y(n_497)
);

INVx4_ASAP7_75t_SL g498 ( 
.A(n_393),
.Y(n_498)
);

INVx3_ASAP7_75t_L g499 ( 
.A(n_393),
.Y(n_499)
);

INVx1_ASAP7_75t_L g500 ( 
.A(n_387),
.Y(n_500)
);

INVx1_ASAP7_75t_L g501 ( 
.A(n_389),
.Y(n_501)
);

NOR2xp33_ASAP7_75t_L g502 ( 
.A(n_427),
.B(n_260),
.Y(n_502)
);

AND2x6_ASAP7_75t_L g503 ( 
.A(n_418),
.B(n_281),
.Y(n_503)
);

INVx4_ASAP7_75t_L g504 ( 
.A(n_393),
.Y(n_504)
);

INVx1_ASAP7_75t_L g505 ( 
.A(n_389),
.Y(n_505)
);

INVx1_ASAP7_75t_L g506 ( 
.A(n_392),
.Y(n_506)
);

AO22x2_ASAP7_75t_L g507 ( 
.A1(n_449),
.A2(n_399),
.B1(n_416),
.B2(n_404),
.Y(n_507)
);

AO22x2_ASAP7_75t_L g508 ( 
.A1(n_437),
.A2(n_423),
.B1(n_388),
.B2(n_405),
.Y(n_508)
);

NAND2xp5_ASAP7_75t_L g509 ( 
.A(n_502),
.B(n_417),
.Y(n_509)
);

INVx2_ASAP7_75t_L g510 ( 
.A(n_490),
.Y(n_510)
);

INVx2_ASAP7_75t_L g511 ( 
.A(n_496),
.Y(n_511)
);

AND2x4_ASAP7_75t_L g512 ( 
.A(n_491),
.B(n_457),
.Y(n_512)
);

AND2x6_ASAP7_75t_L g513 ( 
.A(n_488),
.B(n_423),
.Y(n_513)
);

NAND2xp5_ASAP7_75t_SL g514 ( 
.A(n_439),
.B(n_422),
.Y(n_514)
);

INVx2_ASAP7_75t_L g515 ( 
.A(n_462),
.Y(n_515)
);

OAI221xp5_ASAP7_75t_L g516 ( 
.A1(n_439),
.A2(n_380),
.B1(n_395),
.B2(n_407),
.C(n_392),
.Y(n_516)
);

INVx2_ASAP7_75t_L g517 ( 
.A(n_476),
.Y(n_517)
);

INVx2_ASAP7_75t_L g518 ( 
.A(n_443),
.Y(n_518)
);

OAI22xp5_ASAP7_75t_SL g519 ( 
.A1(n_468),
.A2(n_415),
.B1(n_409),
.B2(n_397),
.Y(n_519)
);

NAND2xp5_ASAP7_75t_SL g520 ( 
.A(n_445),
.B(n_409),
.Y(n_520)
);

AO22x2_ASAP7_75t_L g521 ( 
.A1(n_457),
.A2(n_397),
.B1(n_396),
.B2(n_374),
.Y(n_521)
);

INVx1_ASAP7_75t_L g522 ( 
.A(n_474),
.Y(n_522)
);

OAI221xp5_ASAP7_75t_L g523 ( 
.A1(n_486),
.A2(n_409),
.B1(n_396),
.B2(n_374),
.C(n_377),
.Y(n_523)
);

INVx1_ASAP7_75t_L g524 ( 
.A(n_477),
.Y(n_524)
);

INVx1_ASAP7_75t_L g525 ( 
.A(n_481),
.Y(n_525)
);

INVx1_ASAP7_75t_L g526 ( 
.A(n_485),
.Y(n_526)
);

INVx2_ASAP7_75t_L g527 ( 
.A(n_454),
.Y(n_527)
);

INVx2_ASAP7_75t_L g528 ( 
.A(n_458),
.Y(n_528)
);

INVx1_ASAP7_75t_L g529 ( 
.A(n_495),
.Y(n_529)
);

BUFx8_ASAP7_75t_L g530 ( 
.A(n_455),
.Y(n_530)
);

INVx1_ASAP7_75t_L g531 ( 
.A(n_500),
.Y(n_531)
);

AND2x2_ASAP7_75t_L g532 ( 
.A(n_432),
.B(n_378),
.Y(n_532)
);

BUFx6f_ASAP7_75t_SL g533 ( 
.A(n_431),
.Y(n_533)
);

NAND2xp5_ASAP7_75t_L g534 ( 
.A(n_502),
.B(n_378),
.Y(n_534)
);

INVx1_ASAP7_75t_L g535 ( 
.A(n_501),
.Y(n_535)
);

NAND2xp5_ASAP7_75t_L g536 ( 
.A(n_471),
.B(n_378),
.Y(n_536)
);

AO22x2_ASAP7_75t_L g537 ( 
.A1(n_492),
.A2(n_375),
.B1(n_377),
.B2(n_376),
.Y(n_537)
);

OAI221xp5_ASAP7_75t_L g538 ( 
.A1(n_486),
.A2(n_375),
.B1(n_379),
.B2(n_393),
.C(n_305),
.Y(n_538)
);

INVx1_ASAP7_75t_L g539 ( 
.A(n_505),
.Y(n_539)
);

AO22x2_ASAP7_75t_L g540 ( 
.A1(n_438),
.A2(n_379),
.B1(n_9),
.B2(n_10),
.Y(n_540)
);

INVx1_ASAP7_75t_L g541 ( 
.A(n_506),
.Y(n_541)
);

AND2x2_ASAP7_75t_L g542 ( 
.A(n_433),
.B(n_379),
.Y(n_542)
);

INVx1_ASAP7_75t_L g543 ( 
.A(n_436),
.Y(n_543)
);

INVx1_ASAP7_75t_L g544 ( 
.A(n_442),
.Y(n_544)
);

NAND2xp5_ASAP7_75t_L g545 ( 
.A(n_471),
.B(n_261),
.Y(n_545)
);

NAND2xp5_ASAP7_75t_L g546 ( 
.A(n_433),
.B(n_262),
.Y(n_546)
);

AND2x4_ASAP7_75t_L g547 ( 
.A(n_473),
.B(n_8),
.Y(n_547)
);

INVx1_ASAP7_75t_L g548 ( 
.A(n_446),
.Y(n_548)
);

INVx1_ASAP7_75t_L g549 ( 
.A(n_447),
.Y(n_549)
);

INVx2_ASAP7_75t_L g550 ( 
.A(n_450),
.Y(n_550)
);

INVx1_ASAP7_75t_L g551 ( 
.A(n_451),
.Y(n_551)
);

INVx1_ASAP7_75t_L g552 ( 
.A(n_452),
.Y(n_552)
);

INVxp67_ASAP7_75t_L g553 ( 
.A(n_435),
.Y(n_553)
);

INVx1_ASAP7_75t_L g554 ( 
.A(n_465),
.Y(n_554)
);

AND2x2_ASAP7_75t_L g555 ( 
.A(n_463),
.B(n_10),
.Y(n_555)
);

AO22x2_ASAP7_75t_L g556 ( 
.A1(n_483),
.A2(n_11),
.B1(n_12),
.B2(n_14),
.Y(n_556)
);

INVxp67_ASAP7_75t_L g557 ( 
.A(n_463),
.Y(n_557)
);

INVx1_ASAP7_75t_L g558 ( 
.A(n_493),
.Y(n_558)
);

AND2x4_ASAP7_75t_L g559 ( 
.A(n_473),
.B(n_14),
.Y(n_559)
);

AO22x2_ASAP7_75t_L g560 ( 
.A1(n_488),
.A2(n_15),
.B1(n_16),
.B2(n_17),
.Y(n_560)
);

AO22x2_ASAP7_75t_L g561 ( 
.A1(n_441),
.A2(n_15),
.B1(n_17),
.B2(n_18),
.Y(n_561)
);

NAND2x1p5_ASAP7_75t_L g562 ( 
.A(n_459),
.B(n_480),
.Y(n_562)
);

BUFx8_ASAP7_75t_L g563 ( 
.A(n_464),
.Y(n_563)
);

AOI22xp5_ASAP7_75t_L g564 ( 
.A1(n_461),
.A2(n_494),
.B1(n_453),
.B2(n_475),
.Y(n_564)
);

AND2x4_ASAP7_75t_L g565 ( 
.A(n_475),
.B(n_19),
.Y(n_565)
);

INVxp67_ASAP7_75t_L g566 ( 
.A(n_431),
.Y(n_566)
);

INVx1_ASAP7_75t_L g567 ( 
.A(n_493),
.Y(n_567)
);

AO22x2_ASAP7_75t_L g568 ( 
.A1(n_464),
.A2(n_19),
.B1(n_20),
.B2(n_22),
.Y(n_568)
);

AO22x2_ASAP7_75t_L g569 ( 
.A1(n_461),
.A2(n_20),
.B1(n_23),
.B2(n_24),
.Y(n_569)
);

NAND2x1p5_ASAP7_75t_L g570 ( 
.A(n_445),
.B(n_23),
.Y(n_570)
);

INVx1_ASAP7_75t_L g571 ( 
.A(n_487),
.Y(n_571)
);

NAND2x1p5_ASAP7_75t_L g572 ( 
.A(n_453),
.B(n_25),
.Y(n_572)
);

HB1xp67_ASAP7_75t_L g573 ( 
.A(n_431),
.Y(n_573)
);

INVx1_ASAP7_75t_L g574 ( 
.A(n_487),
.Y(n_574)
);

NOR2xp33_ASAP7_75t_L g575 ( 
.A(n_494),
.B(n_263),
.Y(n_575)
);

OAI221xp5_ASAP7_75t_L g576 ( 
.A1(n_489),
.A2(n_304),
.B1(n_300),
.B2(n_299),
.C(n_298),
.Y(n_576)
);

AOI22xp5_ASAP7_75t_L g577 ( 
.A1(n_489),
.A2(n_297),
.B1(n_294),
.B2(n_291),
.Y(n_577)
);

INVx1_ASAP7_75t_L g578 ( 
.A(n_456),
.Y(n_578)
);

BUFx6f_ASAP7_75t_SL g579 ( 
.A(n_478),
.Y(n_579)
);

INVx1_ASAP7_75t_L g580 ( 
.A(n_456),
.Y(n_580)
);

AO22x2_ASAP7_75t_L g581 ( 
.A1(n_469),
.A2(n_466),
.B1(n_482),
.B2(n_497),
.Y(n_581)
);

INVxp67_ASAP7_75t_L g582 ( 
.A(n_448),
.Y(n_582)
);

INVx1_ASAP7_75t_L g583 ( 
.A(n_466),
.Y(n_583)
);

NAND2xp5_ASAP7_75t_L g584 ( 
.A(n_448),
.B(n_264),
.Y(n_584)
);

INVx1_ASAP7_75t_L g585 ( 
.A(n_467),
.Y(n_585)
);

OAI22xp5_ASAP7_75t_L g586 ( 
.A1(n_434),
.A2(n_278),
.B1(n_287),
.B2(n_286),
.Y(n_586)
);

INVx2_ASAP7_75t_L g587 ( 
.A(n_460),
.Y(n_587)
);

INVx1_ASAP7_75t_L g588 ( 
.A(n_467),
.Y(n_588)
);

NAND2xp5_ASAP7_75t_L g589 ( 
.A(n_434),
.B(n_268),
.Y(n_589)
);

INVx1_ASAP7_75t_L g590 ( 
.A(n_470),
.Y(n_590)
);

INVxp67_ASAP7_75t_L g591 ( 
.A(n_430),
.Y(n_591)
);

NAND2xp5_ASAP7_75t_L g592 ( 
.A(n_509),
.B(n_478),
.Y(n_592)
);

NAND2xp33_ASAP7_75t_SL g593 ( 
.A(n_579),
.B(n_470),
.Y(n_593)
);

NAND2xp5_ASAP7_75t_SL g594 ( 
.A(n_512),
.B(n_504),
.Y(n_594)
);

NAND2xp5_ASAP7_75t_SL g595 ( 
.A(n_512),
.B(n_504),
.Y(n_595)
);

NAND2xp5_ASAP7_75t_SL g596 ( 
.A(n_564),
.B(n_547),
.Y(n_596)
);

NAND2xp5_ASAP7_75t_SL g597 ( 
.A(n_547),
.B(n_440),
.Y(n_597)
);

NAND2xp5_ASAP7_75t_L g598 ( 
.A(n_582),
.B(n_503),
.Y(n_598)
);

NAND2xp5_ASAP7_75t_SL g599 ( 
.A(n_559),
.B(n_565),
.Y(n_599)
);

NAND2xp5_ASAP7_75t_SL g600 ( 
.A(n_559),
.B(n_440),
.Y(n_600)
);

NAND2xp5_ASAP7_75t_SL g601 ( 
.A(n_565),
.B(n_571),
.Y(n_601)
);

NAND2xp5_ASAP7_75t_SL g602 ( 
.A(n_574),
.B(n_440),
.Y(n_602)
);

NAND2xp5_ASAP7_75t_SL g603 ( 
.A(n_542),
.B(n_444),
.Y(n_603)
);

NAND2xp5_ASAP7_75t_SL g604 ( 
.A(n_563),
.B(n_444),
.Y(n_604)
);

NAND2xp33_ASAP7_75t_SL g605 ( 
.A(n_546),
.B(n_460),
.Y(n_605)
);

NAND2xp5_ASAP7_75t_SL g606 ( 
.A(n_563),
.B(n_444),
.Y(n_606)
);

NAND2xp5_ASAP7_75t_SL g607 ( 
.A(n_557),
.B(n_472),
.Y(n_607)
);

NAND2xp5_ASAP7_75t_L g608 ( 
.A(n_513),
.B(n_503),
.Y(n_608)
);

NAND2xp5_ASAP7_75t_SL g609 ( 
.A(n_514),
.B(n_472),
.Y(n_609)
);

NAND2xp5_ASAP7_75t_L g610 ( 
.A(n_513),
.B(n_503),
.Y(n_610)
);

NAND2xp5_ASAP7_75t_L g611 ( 
.A(n_513),
.B(n_503),
.Y(n_611)
);

NAND2xp5_ASAP7_75t_SL g612 ( 
.A(n_519),
.B(n_472),
.Y(n_612)
);

NAND2xp5_ASAP7_75t_SL g613 ( 
.A(n_545),
.B(n_479),
.Y(n_613)
);

NAND2xp33_ASAP7_75t_SL g614 ( 
.A(n_555),
.B(n_484),
.Y(n_614)
);

NAND2xp5_ASAP7_75t_SL g615 ( 
.A(n_575),
.B(n_479),
.Y(n_615)
);

NAND2xp5_ASAP7_75t_SL g616 ( 
.A(n_536),
.B(n_479),
.Y(n_616)
);

NAND2xp5_ASAP7_75t_SL g617 ( 
.A(n_534),
.B(n_484),
.Y(n_617)
);

NAND2xp5_ASAP7_75t_SL g618 ( 
.A(n_532),
.B(n_499),
.Y(n_618)
);

NAND2xp33_ASAP7_75t_SL g619 ( 
.A(n_522),
.B(n_499),
.Y(n_619)
);

NAND2xp5_ASAP7_75t_SL g620 ( 
.A(n_584),
.B(n_498),
.Y(n_620)
);

NAND2xp33_ASAP7_75t_SL g621 ( 
.A(n_524),
.B(n_271),
.Y(n_621)
);

NAND2xp33_ASAP7_75t_SL g622 ( 
.A(n_525),
.B(n_276),
.Y(n_622)
);

NAND2xp5_ASAP7_75t_L g623 ( 
.A(n_567),
.B(n_503),
.Y(n_623)
);

NAND2xp5_ASAP7_75t_SL g624 ( 
.A(n_553),
.B(n_498),
.Y(n_624)
);

NAND2xp5_ASAP7_75t_SL g625 ( 
.A(n_558),
.B(n_498),
.Y(n_625)
);

NAND2xp5_ASAP7_75t_SL g626 ( 
.A(n_558),
.B(n_277),
.Y(n_626)
);

NAND2xp5_ASAP7_75t_SL g627 ( 
.A(n_526),
.B(n_285),
.Y(n_627)
);

NAND2xp5_ASAP7_75t_L g628 ( 
.A(n_578),
.B(n_289),
.Y(n_628)
);

NAND2xp5_ASAP7_75t_SL g629 ( 
.A(n_529),
.B(n_25),
.Y(n_629)
);

NAND2xp5_ASAP7_75t_L g630 ( 
.A(n_580),
.B(n_26),
.Y(n_630)
);

NAND2xp5_ASAP7_75t_SL g631 ( 
.A(n_531),
.B(n_26),
.Y(n_631)
);

NAND2xp5_ASAP7_75t_L g632 ( 
.A(n_583),
.B(n_27),
.Y(n_632)
);

NAND2xp5_ASAP7_75t_SL g633 ( 
.A(n_535),
.B(n_27),
.Y(n_633)
);

NAND2xp5_ASAP7_75t_SL g634 ( 
.A(n_539),
.B(n_28),
.Y(n_634)
);

NAND2xp33_ASAP7_75t_SL g635 ( 
.A(n_541),
.B(n_29),
.Y(n_635)
);

NAND2xp5_ASAP7_75t_SL g636 ( 
.A(n_591),
.B(n_29),
.Y(n_636)
);

NAND2xp5_ASAP7_75t_SL g637 ( 
.A(n_589),
.B(n_30),
.Y(n_637)
);

AND2x4_ASAP7_75t_L g638 ( 
.A(n_566),
.B(n_30),
.Y(n_638)
);

AND2x2_ASAP7_75t_L g639 ( 
.A(n_507),
.B(n_31),
.Y(n_639)
);

NAND2xp5_ASAP7_75t_SL g640 ( 
.A(n_572),
.B(n_32),
.Y(n_640)
);

NAND2xp5_ASAP7_75t_SL g641 ( 
.A(n_586),
.B(n_32),
.Y(n_641)
);

NAND2xp5_ASAP7_75t_SL g642 ( 
.A(n_577),
.B(n_33),
.Y(n_642)
);

NAND2xp33_ASAP7_75t_SL g643 ( 
.A(n_533),
.B(n_520),
.Y(n_643)
);

NOR2xp33_ASAP7_75t_SL g644 ( 
.A(n_530),
.B(n_36),
.Y(n_644)
);

NAND2xp5_ASAP7_75t_SL g645 ( 
.A(n_570),
.B(n_37),
.Y(n_645)
);

NAND2xp5_ASAP7_75t_L g646 ( 
.A(n_585),
.B(n_588),
.Y(n_646)
);

NAND2xp5_ASAP7_75t_SL g647 ( 
.A(n_562),
.B(n_38),
.Y(n_647)
);

NAND2xp5_ASAP7_75t_SL g648 ( 
.A(n_590),
.B(n_530),
.Y(n_648)
);

NAND2xp33_ASAP7_75t_SL g649 ( 
.A(n_573),
.B(n_39),
.Y(n_649)
);

NAND2xp5_ASAP7_75t_SL g650 ( 
.A(n_543),
.B(n_40),
.Y(n_650)
);

NAND2xp33_ASAP7_75t_SL g651 ( 
.A(n_544),
.B(n_45),
.Y(n_651)
);

NAND2xp5_ASAP7_75t_SL g652 ( 
.A(n_548),
.B(n_46),
.Y(n_652)
);

NAND2xp33_ASAP7_75t_SL g653 ( 
.A(n_549),
.B(n_47),
.Y(n_653)
);

NAND2xp5_ASAP7_75t_SL g654 ( 
.A(n_551),
.B(n_48),
.Y(n_654)
);

NAND2xp33_ASAP7_75t_SL g655 ( 
.A(n_552),
.B(n_554),
.Y(n_655)
);

NAND2xp33_ASAP7_75t_SL g656 ( 
.A(n_587),
.B(n_550),
.Y(n_656)
);

AND2x4_ASAP7_75t_L g657 ( 
.A(n_518),
.B(n_50),
.Y(n_657)
);

NAND2xp5_ASAP7_75t_SL g658 ( 
.A(n_527),
.B(n_52),
.Y(n_658)
);

A2O1A1Ixp33_ASAP7_75t_L g659 ( 
.A1(n_655),
.A2(n_592),
.B(n_646),
.C(n_596),
.Y(n_659)
);

NAND2xp5_ASAP7_75t_L g660 ( 
.A(n_601),
.B(n_537),
.Y(n_660)
);

AOI221xp5_ASAP7_75t_SL g661 ( 
.A1(n_641),
.A2(n_523),
.B1(n_516),
.B2(n_538),
.C(n_576),
.Y(n_661)
);

OAI21x1_ASAP7_75t_L g662 ( 
.A1(n_616),
.A2(n_528),
.B(n_515),
.Y(n_662)
);

NAND2xp5_ASAP7_75t_L g663 ( 
.A(n_599),
.B(n_537),
.Y(n_663)
);

NAND2xp5_ASAP7_75t_SL g664 ( 
.A(n_598),
.B(n_510),
.Y(n_664)
);

A2O1A1Ixp33_ASAP7_75t_L g665 ( 
.A1(n_642),
.A2(n_511),
.B(n_517),
.C(n_569),
.Y(n_665)
);

AO21x1_ASAP7_75t_L g666 ( 
.A1(n_651),
.A2(n_569),
.B(n_521),
.Y(n_666)
);

INVx3_ASAP7_75t_L g667 ( 
.A(n_657),
.Y(n_667)
);

OAI21xp5_ASAP7_75t_L g668 ( 
.A1(n_630),
.A2(n_581),
.B(n_521),
.Y(n_668)
);

INVx1_ASAP7_75t_L g669 ( 
.A(n_632),
.Y(n_669)
);

NAND3xp33_ASAP7_75t_SL g670 ( 
.A(n_635),
.B(n_644),
.C(n_636),
.Y(n_670)
);

OAI21xp5_ASAP7_75t_L g671 ( 
.A1(n_623),
.A2(n_581),
.B(n_508),
.Y(n_671)
);

NAND2xp5_ASAP7_75t_L g672 ( 
.A(n_638),
.B(n_508),
.Y(n_672)
);

AO31x2_ASAP7_75t_L g673 ( 
.A1(n_628),
.A2(n_540),
.A3(n_560),
.B(n_556),
.Y(n_673)
);

AO31x2_ASAP7_75t_L g674 ( 
.A1(n_608),
.A2(n_540),
.A3(n_560),
.B(n_556),
.Y(n_674)
);

NAND2xp5_ASAP7_75t_L g675 ( 
.A(n_638),
.B(n_507),
.Y(n_675)
);

AOI21x1_ASAP7_75t_SL g676 ( 
.A1(n_610),
.A2(n_568),
.B(n_561),
.Y(n_676)
);

CKINVDCx5p33_ASAP7_75t_R g677 ( 
.A(n_648),
.Y(n_677)
);

NOR2xp33_ASAP7_75t_L g678 ( 
.A(n_597),
.B(n_53),
.Y(n_678)
);

AND2x2_ASAP7_75t_L g679 ( 
.A(n_639),
.B(n_568),
.Y(n_679)
);

OAI21xp5_ASAP7_75t_L g680 ( 
.A1(n_618),
.A2(n_561),
.B(n_57),
.Y(n_680)
);

OAI21x1_ASAP7_75t_L g681 ( 
.A1(n_620),
.A2(n_54),
.B(n_58),
.Y(n_681)
);

OAI21xp5_ASAP7_75t_L g682 ( 
.A1(n_617),
.A2(n_603),
.B(n_637),
.Y(n_682)
);

INVx1_ASAP7_75t_L g683 ( 
.A(n_638),
.Y(n_683)
);

AOI21x1_ASAP7_75t_SL g684 ( 
.A1(n_611),
.A2(n_59),
.B(n_61),
.Y(n_684)
);

AO31x2_ASAP7_75t_L g685 ( 
.A1(n_605),
.A2(n_62),
.A3(n_64),
.B(n_65),
.Y(n_685)
);

NAND2xp5_ASAP7_75t_L g686 ( 
.A(n_600),
.B(n_67),
.Y(n_686)
);

O2A1O1Ixp33_ASAP7_75t_L g687 ( 
.A1(n_629),
.A2(n_68),
.B(n_69),
.C(n_70),
.Y(n_687)
);

AO21x1_ASAP7_75t_L g688 ( 
.A1(n_653),
.A2(n_73),
.B(n_74),
.Y(n_688)
);

OAI21xp5_ASAP7_75t_L g689 ( 
.A1(n_650),
.A2(n_80),
.B(n_82),
.Y(n_689)
);

AOI21xp5_ASAP7_75t_L g690 ( 
.A1(n_613),
.A2(n_619),
.B(n_614),
.Y(n_690)
);

NAND2xp5_ASAP7_75t_L g691 ( 
.A(n_612),
.B(n_83),
.Y(n_691)
);

HB1xp67_ASAP7_75t_L g692 ( 
.A(n_657),
.Y(n_692)
);

AOI21x1_ASAP7_75t_L g693 ( 
.A1(n_615),
.A2(n_85),
.B(n_86),
.Y(n_693)
);

NAND3xp33_ASAP7_75t_L g694 ( 
.A(n_640),
.B(n_87),
.C(n_88),
.Y(n_694)
);

INVx2_ASAP7_75t_L g695 ( 
.A(n_657),
.Y(n_695)
);

AOI21x1_ASAP7_75t_L g696 ( 
.A1(n_609),
.A2(n_90),
.B(n_92),
.Y(n_696)
);

AND2x2_ASAP7_75t_L g697 ( 
.A(n_604),
.B(n_93),
.Y(n_697)
);

OAI21x1_ASAP7_75t_L g698 ( 
.A1(n_625),
.A2(n_94),
.B(n_96),
.Y(n_698)
);

NAND2xp5_ASAP7_75t_L g699 ( 
.A(n_594),
.B(n_99),
.Y(n_699)
);

INVx1_ASAP7_75t_L g700 ( 
.A(n_631),
.Y(n_700)
);

OAI21xp33_ASAP7_75t_L g701 ( 
.A1(n_633),
.A2(n_100),
.B(n_102),
.Y(n_701)
);

OA21x2_ASAP7_75t_L g702 ( 
.A1(n_652),
.A2(n_654),
.B(n_602),
.Y(n_702)
);

OAI21x1_ASAP7_75t_L g703 ( 
.A1(n_658),
.A2(n_103),
.B(n_105),
.Y(n_703)
);

AO31x2_ASAP7_75t_L g704 ( 
.A1(n_656),
.A2(n_106),
.A3(n_107),
.B(n_110),
.Y(n_704)
);

OAI21x1_ASAP7_75t_L g705 ( 
.A1(n_647),
.A2(n_112),
.B(n_114),
.Y(n_705)
);

AOI221x1_ASAP7_75t_L g706 ( 
.A1(n_649),
.A2(n_115),
.B1(n_116),
.B2(n_117),
.C(n_118),
.Y(n_706)
);

AOI21xp5_ASAP7_75t_L g707 ( 
.A1(n_626),
.A2(n_607),
.B(n_627),
.Y(n_707)
);

NAND2xp5_ASAP7_75t_L g708 ( 
.A(n_595),
.B(n_121),
.Y(n_708)
);

NAND2x1_ASAP7_75t_L g709 ( 
.A(n_593),
.B(n_122),
.Y(n_709)
);

INVx1_ASAP7_75t_L g710 ( 
.A(n_634),
.Y(n_710)
);

INVx1_ASAP7_75t_L g711 ( 
.A(n_624),
.Y(n_711)
);

INVx1_ASAP7_75t_L g712 ( 
.A(n_606),
.Y(n_712)
);

INVx5_ASAP7_75t_L g713 ( 
.A(n_643),
.Y(n_713)
);

INVx1_ASAP7_75t_L g714 ( 
.A(n_683),
.Y(n_714)
);

BUFx2_ASAP7_75t_L g715 ( 
.A(n_677),
.Y(n_715)
);

CKINVDCx6p67_ASAP7_75t_R g716 ( 
.A(n_713),
.Y(n_716)
);

OAI21x1_ASAP7_75t_L g717 ( 
.A1(n_684),
.A2(n_645),
.B(n_622),
.Y(n_717)
);

BUFx2_ASAP7_75t_L g718 ( 
.A(n_712),
.Y(n_718)
);

INVx1_ASAP7_75t_L g719 ( 
.A(n_700),
.Y(n_719)
);

NAND2xp5_ASAP7_75t_L g720 ( 
.A(n_669),
.B(n_621),
.Y(n_720)
);

INVx1_ASAP7_75t_L g721 ( 
.A(n_710),
.Y(n_721)
);

AND2x4_ASAP7_75t_L g722 ( 
.A(n_713),
.B(n_123),
.Y(n_722)
);

NAND2xp5_ASAP7_75t_L g723 ( 
.A(n_679),
.B(n_713),
.Y(n_723)
);

AO21x2_ASAP7_75t_L g724 ( 
.A1(n_671),
.A2(n_124),
.B(n_125),
.Y(n_724)
);

OAI21x1_ASAP7_75t_L g725 ( 
.A1(n_690),
.A2(n_128),
.B(n_129),
.Y(n_725)
);

AOI22xp33_ASAP7_75t_L g726 ( 
.A1(n_666),
.A2(n_131),
.B1(n_135),
.B2(n_136),
.Y(n_726)
);

NAND2xp5_ASAP7_75t_L g727 ( 
.A(n_673),
.B(n_220),
.Y(n_727)
);

INVx6_ASAP7_75t_SL g728 ( 
.A(n_670),
.Y(n_728)
);

OAI21x1_ASAP7_75t_L g729 ( 
.A1(n_681),
.A2(n_137),
.B(n_140),
.Y(n_729)
);

NOR2xp67_ASAP7_75t_L g730 ( 
.A(n_707),
.B(n_141),
.Y(n_730)
);

AOI21xp5_ASAP7_75t_L g731 ( 
.A1(n_659),
.A2(n_667),
.B(n_689),
.Y(n_731)
);

INVx2_ASAP7_75t_L g732 ( 
.A(n_662),
.Y(n_732)
);

BUFx2_ASAP7_75t_L g733 ( 
.A(n_674),
.Y(n_733)
);

BUFx2_ASAP7_75t_L g734 ( 
.A(n_674),
.Y(n_734)
);

AND2x4_ASAP7_75t_L g735 ( 
.A(n_667),
.B(n_142),
.Y(n_735)
);

AOI21x1_ASAP7_75t_L g736 ( 
.A1(n_668),
.A2(n_144),
.B(n_145),
.Y(n_736)
);

CKINVDCx9p33_ASAP7_75t_R g737 ( 
.A(n_678),
.Y(n_737)
);

OR2x2_ASAP7_75t_L g738 ( 
.A(n_675),
.B(n_146),
.Y(n_738)
);

INVx4_ASAP7_75t_L g739 ( 
.A(n_692),
.Y(n_739)
);

NAND2xp5_ASAP7_75t_L g740 ( 
.A(n_673),
.B(n_219),
.Y(n_740)
);

INVx2_ASAP7_75t_L g741 ( 
.A(n_695),
.Y(n_741)
);

BUFx2_ASAP7_75t_L g742 ( 
.A(n_674),
.Y(n_742)
);

AOI21xp5_ASAP7_75t_SL g743 ( 
.A1(n_665),
.A2(n_148),
.B(n_149),
.Y(n_743)
);

OA21x2_ASAP7_75t_L g744 ( 
.A1(n_706),
.A2(n_150),
.B(n_151),
.Y(n_744)
);

OA21x2_ASAP7_75t_L g745 ( 
.A1(n_661),
.A2(n_154),
.B(n_156),
.Y(n_745)
);

CKINVDCx9p33_ASAP7_75t_R g746 ( 
.A(n_691),
.Y(n_746)
);

NOR3xp33_ASAP7_75t_L g747 ( 
.A(n_680),
.B(n_157),
.C(n_158),
.Y(n_747)
);

OR2x2_ASAP7_75t_L g748 ( 
.A(n_672),
.B(n_160),
.Y(n_748)
);

INVx1_ASAP7_75t_L g749 ( 
.A(n_711),
.Y(n_749)
);

OAI21x1_ASAP7_75t_L g750 ( 
.A1(n_693),
.A2(n_161),
.B(n_162),
.Y(n_750)
);

INVx2_ASAP7_75t_L g751 ( 
.A(n_698),
.Y(n_751)
);

AND2x4_ASAP7_75t_L g752 ( 
.A(n_663),
.B(n_163),
.Y(n_752)
);

OA21x2_ASAP7_75t_L g753 ( 
.A1(n_661),
.A2(n_165),
.B(n_167),
.Y(n_753)
);

INVx1_ASAP7_75t_L g754 ( 
.A(n_660),
.Y(n_754)
);

AOI21x1_ASAP7_75t_L g755 ( 
.A1(n_664),
.A2(n_168),
.B(n_170),
.Y(n_755)
);

NAND2xp5_ASAP7_75t_L g756 ( 
.A(n_673),
.B(n_171),
.Y(n_756)
);

OAI21x1_ASAP7_75t_L g757 ( 
.A1(n_696),
.A2(n_175),
.B(n_176),
.Y(n_757)
);

AOI21xp5_ASAP7_75t_L g758 ( 
.A1(n_689),
.A2(n_177),
.B(n_179),
.Y(n_758)
);

OAI21x1_ASAP7_75t_L g759 ( 
.A1(n_703),
.A2(n_180),
.B(n_182),
.Y(n_759)
);

INVxp67_ASAP7_75t_L g760 ( 
.A(n_697),
.Y(n_760)
);

BUFx3_ASAP7_75t_L g761 ( 
.A(n_709),
.Y(n_761)
);

NOR2xp67_ASAP7_75t_L g762 ( 
.A(n_686),
.B(n_184),
.Y(n_762)
);

INVxp67_ASAP7_75t_L g763 ( 
.A(n_682),
.Y(n_763)
);

INVx1_ASAP7_75t_L g764 ( 
.A(n_682),
.Y(n_764)
);

AOI22xp33_ASAP7_75t_L g765 ( 
.A1(n_701),
.A2(n_185),
.B1(n_186),
.B2(n_188),
.Y(n_765)
);

INVx4_ASAP7_75t_L g766 ( 
.A(n_716),
.Y(n_766)
);

AND2x2_ASAP7_75t_L g767 ( 
.A(n_764),
.B(n_704),
.Y(n_767)
);

INVx2_ASAP7_75t_L g768 ( 
.A(n_741),
.Y(n_768)
);

INVx1_ASAP7_75t_L g769 ( 
.A(n_733),
.Y(n_769)
);

NAND2xp5_ASAP7_75t_L g770 ( 
.A(n_763),
.B(n_701),
.Y(n_770)
);

O2A1O1Ixp33_ASAP7_75t_SL g771 ( 
.A1(n_720),
.A2(n_694),
.B(n_687),
.C(n_699),
.Y(n_771)
);

BUFx12f_ASAP7_75t_L g772 ( 
.A(n_715),
.Y(n_772)
);

INVx1_ASAP7_75t_L g773 ( 
.A(n_734),
.Y(n_773)
);

CKINVDCx6p67_ASAP7_75t_R g774 ( 
.A(n_746),
.Y(n_774)
);

OR2x2_ASAP7_75t_L g775 ( 
.A(n_742),
.B(n_704),
.Y(n_775)
);

INVx1_ASAP7_75t_L g776 ( 
.A(n_754),
.Y(n_776)
);

INVx1_ASAP7_75t_L g777 ( 
.A(n_714),
.Y(n_777)
);

OR2x2_ASAP7_75t_L g778 ( 
.A(n_723),
.B(n_704),
.Y(n_778)
);

INVx1_ASAP7_75t_L g779 ( 
.A(n_732),
.Y(n_779)
);

AOI22xp33_ASAP7_75t_L g780 ( 
.A1(n_747),
.A2(n_694),
.B1(n_688),
.B2(n_702),
.Y(n_780)
);

INVx2_ASAP7_75t_L g781 ( 
.A(n_749),
.Y(n_781)
);

INVx2_ASAP7_75t_L g782 ( 
.A(n_719),
.Y(n_782)
);

AOI22xp33_ASAP7_75t_L g783 ( 
.A1(n_752),
.A2(n_702),
.B1(n_676),
.B2(n_708),
.Y(n_783)
);

AND2x4_ASAP7_75t_L g784 ( 
.A(n_752),
.B(n_685),
.Y(n_784)
);

AND2x2_ASAP7_75t_L g785 ( 
.A(n_721),
.B(n_718),
.Y(n_785)
);

INVx1_ASAP7_75t_L g786 ( 
.A(n_727),
.Y(n_786)
);

INVx1_ASAP7_75t_L g787 ( 
.A(n_740),
.Y(n_787)
);

INVx1_ASAP7_75t_L g788 ( 
.A(n_756),
.Y(n_788)
);

INVx2_ASAP7_75t_L g789 ( 
.A(n_751),
.Y(n_789)
);

NAND2xp5_ASAP7_75t_L g790 ( 
.A(n_760),
.B(n_685),
.Y(n_790)
);

BUFx12f_ASAP7_75t_L g791 ( 
.A(n_722),
.Y(n_791)
);

NAND2xp5_ASAP7_75t_L g792 ( 
.A(n_716),
.B(n_685),
.Y(n_792)
);

INVx1_ASAP7_75t_L g793 ( 
.A(n_724),
.Y(n_793)
);

OAI21x1_ASAP7_75t_L g794 ( 
.A1(n_725),
.A2(n_705),
.B(n_193),
.Y(n_794)
);

INVx2_ASAP7_75t_L g795 ( 
.A(n_751),
.Y(n_795)
);

OAI21x1_ASAP7_75t_L g796 ( 
.A1(n_725),
.A2(n_731),
.B(n_750),
.Y(n_796)
);

INVx1_ASAP7_75t_L g797 ( 
.A(n_724),
.Y(n_797)
);

HB1xp67_ASAP7_75t_L g798 ( 
.A(n_739),
.Y(n_798)
);

INVx1_ASAP7_75t_L g799 ( 
.A(n_736),
.Y(n_799)
);

INVx1_ASAP7_75t_L g800 ( 
.A(n_745),
.Y(n_800)
);

AO21x1_ASAP7_75t_SL g801 ( 
.A1(n_765),
.A2(n_189),
.B(n_198),
.Y(n_801)
);

HB1xp67_ASAP7_75t_L g802 ( 
.A(n_739),
.Y(n_802)
);

BUFx2_ASAP7_75t_L g803 ( 
.A(n_739),
.Y(n_803)
);

INVx2_ASAP7_75t_L g804 ( 
.A(n_745),
.Y(n_804)
);

INVx1_ASAP7_75t_L g805 ( 
.A(n_745),
.Y(n_805)
);

NAND2xp5_ASAP7_75t_L g806 ( 
.A(n_752),
.B(n_199),
.Y(n_806)
);

INVx1_ASAP7_75t_L g807 ( 
.A(n_753),
.Y(n_807)
);

INVx1_ASAP7_75t_L g808 ( 
.A(n_753),
.Y(n_808)
);

INVx2_ASAP7_75t_L g809 ( 
.A(n_753),
.Y(n_809)
);

INVx1_ASAP7_75t_L g810 ( 
.A(n_730),
.Y(n_810)
);

INVx2_ASAP7_75t_L g811 ( 
.A(n_744),
.Y(n_811)
);

AND2x2_ASAP7_75t_L g812 ( 
.A(n_735),
.B(n_201),
.Y(n_812)
);

INVx2_ASAP7_75t_L g813 ( 
.A(n_744),
.Y(n_813)
);

HB1xp67_ASAP7_75t_L g814 ( 
.A(n_735),
.Y(n_814)
);

INVx1_ASAP7_75t_L g815 ( 
.A(n_744),
.Y(n_815)
);

OAI22xp5_ASAP7_75t_L g816 ( 
.A1(n_728),
.A2(n_203),
.B1(n_204),
.B2(n_205),
.Y(n_816)
);

INVx2_ASAP7_75t_L g817 ( 
.A(n_757),
.Y(n_817)
);

INVx1_ASAP7_75t_L g818 ( 
.A(n_755),
.Y(n_818)
);

AND2x2_ASAP7_75t_L g819 ( 
.A(n_735),
.B(n_206),
.Y(n_819)
);

INVx6_ASAP7_75t_L g820 ( 
.A(n_722),
.Y(n_820)
);

INVx1_ASAP7_75t_L g821 ( 
.A(n_748),
.Y(n_821)
);

INVxp67_ASAP7_75t_L g822 ( 
.A(n_785),
.Y(n_822)
);

XNOR2xp5_ASAP7_75t_L g823 ( 
.A(n_785),
.B(n_722),
.Y(n_823)
);

NAND2xp5_ASAP7_75t_L g824 ( 
.A(n_781),
.B(n_738),
.Y(n_824)
);

CKINVDCx20_ASAP7_75t_R g825 ( 
.A(n_772),
.Y(n_825)
);

OR2x6_ASAP7_75t_L g826 ( 
.A(n_791),
.B(n_743),
.Y(n_826)
);

NAND2xp33_ASAP7_75t_R g827 ( 
.A(n_812),
.B(n_728),
.Y(n_827)
);

BUFx3_ASAP7_75t_L g828 ( 
.A(n_772),
.Y(n_828)
);

CKINVDCx20_ASAP7_75t_R g829 ( 
.A(n_774),
.Y(n_829)
);

AND2x4_ASAP7_75t_L g830 ( 
.A(n_803),
.B(n_781),
.Y(n_830)
);

HB1xp67_ASAP7_75t_L g831 ( 
.A(n_798),
.Y(n_831)
);

AND2x2_ASAP7_75t_L g832 ( 
.A(n_814),
.B(n_726),
.Y(n_832)
);

AND2x4_ASAP7_75t_L g833 ( 
.A(n_803),
.B(n_761),
.Y(n_833)
);

INVx1_ASAP7_75t_L g834 ( 
.A(n_782),
.Y(n_834)
);

XOR2x2_ASAP7_75t_SL g835 ( 
.A(n_784),
.B(n_728),
.Y(n_835)
);

INVx1_ASAP7_75t_L g836 ( 
.A(n_782),
.Y(n_836)
);

CKINVDCx5p33_ASAP7_75t_R g837 ( 
.A(n_774),
.Y(n_837)
);

AND2x4_ASAP7_75t_L g838 ( 
.A(n_802),
.B(n_761),
.Y(n_838)
);

NAND2xp5_ASAP7_75t_L g839 ( 
.A(n_777),
.B(n_821),
.Y(n_839)
);

OR2x2_ASAP7_75t_L g840 ( 
.A(n_777),
.B(n_726),
.Y(n_840)
);

CKINVDCx5p33_ASAP7_75t_R g841 ( 
.A(n_791),
.Y(n_841)
);

OR2x2_ASAP7_75t_L g842 ( 
.A(n_776),
.B(n_743),
.Y(n_842)
);

INVxp67_ASAP7_75t_L g843 ( 
.A(n_776),
.Y(n_843)
);

NOR2xp33_ASAP7_75t_R g844 ( 
.A(n_820),
.B(n_737),
.Y(n_844)
);

NAND2xp5_ASAP7_75t_L g845 ( 
.A(n_821),
.B(n_770),
.Y(n_845)
);

OR2x6_ASAP7_75t_L g846 ( 
.A(n_820),
.B(n_758),
.Y(n_846)
);

NAND2xp33_ASAP7_75t_R g847 ( 
.A(n_812),
.B(n_819),
.Y(n_847)
);

OR2x6_ASAP7_75t_L g848 ( 
.A(n_820),
.B(n_762),
.Y(n_848)
);

AND2x4_ASAP7_75t_L g849 ( 
.A(n_766),
.B(n_765),
.Y(n_849)
);

AND2x4_ASAP7_75t_L g850 ( 
.A(n_766),
.B(n_717),
.Y(n_850)
);

AND2x2_ASAP7_75t_L g851 ( 
.A(n_819),
.B(n_717),
.Y(n_851)
);

NAND2xp33_ASAP7_75t_R g852 ( 
.A(n_784),
.B(n_737),
.Y(n_852)
);

NAND2xp33_ASAP7_75t_R g853 ( 
.A(n_784),
.B(n_746),
.Y(n_853)
);

NAND2xp33_ASAP7_75t_R g854 ( 
.A(n_784),
.B(n_759),
.Y(n_854)
);

CKINVDCx5p33_ASAP7_75t_R g855 ( 
.A(n_766),
.Y(n_855)
);

XOR2xp5_ASAP7_75t_L g856 ( 
.A(n_778),
.B(n_208),
.Y(n_856)
);

XOR2x2_ASAP7_75t_SL g857 ( 
.A(n_806),
.B(n_210),
.Y(n_857)
);

INVxp67_ASAP7_75t_L g858 ( 
.A(n_790),
.Y(n_858)
);

AND2x2_ASAP7_75t_L g859 ( 
.A(n_820),
.B(n_759),
.Y(n_859)
);

INVx1_ASAP7_75t_L g860 ( 
.A(n_768),
.Y(n_860)
);

BUFx10_ASAP7_75t_L g861 ( 
.A(n_810),
.Y(n_861)
);

NAND2xp5_ASAP7_75t_SL g862 ( 
.A(n_766),
.B(n_757),
.Y(n_862)
);

NOR2xp33_ASAP7_75t_R g863 ( 
.A(n_792),
.B(n_810),
.Y(n_863)
);

NAND2xp5_ASAP7_75t_L g864 ( 
.A(n_786),
.B(n_750),
.Y(n_864)
);

NAND2xp33_ASAP7_75t_SL g865 ( 
.A(n_816),
.B(n_729),
.Y(n_865)
);

OR2x6_ASAP7_75t_L g866 ( 
.A(n_778),
.B(n_773),
.Y(n_866)
);

NAND2xp5_ASAP7_75t_L g867 ( 
.A(n_845),
.B(n_767),
.Y(n_867)
);

INVx1_ASAP7_75t_L g868 ( 
.A(n_834),
.Y(n_868)
);

AND2x4_ASAP7_75t_L g869 ( 
.A(n_830),
.B(n_767),
.Y(n_869)
);

AND2x4_ASAP7_75t_L g870 ( 
.A(n_830),
.B(n_789),
.Y(n_870)
);

NAND2xp5_ASAP7_75t_L g871 ( 
.A(n_843),
.B(n_786),
.Y(n_871)
);

BUFx2_ASAP7_75t_L g872 ( 
.A(n_831),
.Y(n_872)
);

AND2x2_ASAP7_75t_L g873 ( 
.A(n_822),
.B(n_815),
.Y(n_873)
);

INVx2_ASAP7_75t_L g874 ( 
.A(n_860),
.Y(n_874)
);

AND2x2_ASAP7_75t_L g875 ( 
.A(n_866),
.B(n_815),
.Y(n_875)
);

NAND2xp5_ASAP7_75t_L g876 ( 
.A(n_858),
.B(n_788),
.Y(n_876)
);

AND2x2_ASAP7_75t_L g877 ( 
.A(n_866),
.B(n_851),
.Y(n_877)
);

INVx2_ASAP7_75t_L g878 ( 
.A(n_836),
.Y(n_878)
);

AND2x4_ASAP7_75t_L g879 ( 
.A(n_850),
.B(n_789),
.Y(n_879)
);

BUFx2_ASAP7_75t_L g880 ( 
.A(n_833),
.Y(n_880)
);

INVx2_ASAP7_75t_L g881 ( 
.A(n_864),
.Y(n_881)
);

INVx2_ASAP7_75t_L g882 ( 
.A(n_839),
.Y(n_882)
);

AOI22xp33_ASAP7_75t_L g883 ( 
.A1(n_856),
.A2(n_832),
.B1(n_840),
.B2(n_801),
.Y(n_883)
);

NAND2xp5_ASAP7_75t_L g884 ( 
.A(n_824),
.B(n_788),
.Y(n_884)
);

AND2x2_ASAP7_75t_L g885 ( 
.A(n_859),
.B(n_813),
.Y(n_885)
);

INVx1_ASAP7_75t_L g886 ( 
.A(n_842),
.Y(n_886)
);

HB1xp67_ASAP7_75t_L g887 ( 
.A(n_863),
.Y(n_887)
);

INVx1_ASAP7_75t_L g888 ( 
.A(n_850),
.Y(n_888)
);

INVx1_ASAP7_75t_L g889 ( 
.A(n_861),
.Y(n_889)
);

BUFx2_ASAP7_75t_L g890 ( 
.A(n_833),
.Y(n_890)
);

NAND2xp5_ASAP7_75t_L g891 ( 
.A(n_838),
.B(n_787),
.Y(n_891)
);

AOI22xp33_ASAP7_75t_L g892 ( 
.A1(n_849),
.A2(n_801),
.B1(n_787),
.B2(n_783),
.Y(n_892)
);

HB1xp67_ASAP7_75t_L g893 ( 
.A(n_838),
.Y(n_893)
);

OR2x2_ASAP7_75t_L g894 ( 
.A(n_823),
.B(n_773),
.Y(n_894)
);

CKINVDCx11_ASAP7_75t_R g895 ( 
.A(n_825),
.Y(n_895)
);

INVx1_ASAP7_75t_L g896 ( 
.A(n_849),
.Y(n_896)
);

AND2x2_ASAP7_75t_L g897 ( 
.A(n_846),
.B(n_813),
.Y(n_897)
);

NAND2xp5_ASAP7_75t_L g898 ( 
.A(n_855),
.B(n_769),
.Y(n_898)
);

AND2x2_ASAP7_75t_L g899 ( 
.A(n_846),
.B(n_811),
.Y(n_899)
);

AND2x2_ASAP7_75t_L g900 ( 
.A(n_877),
.B(n_811),
.Y(n_900)
);

AND2x2_ASAP7_75t_L g901 ( 
.A(n_877),
.B(n_795),
.Y(n_901)
);

OR2x2_ASAP7_75t_L g902 ( 
.A(n_872),
.B(n_775),
.Y(n_902)
);

INVx3_ASAP7_75t_L g903 ( 
.A(n_888),
.Y(n_903)
);

AOI31xp33_ASAP7_75t_L g904 ( 
.A1(n_887),
.A2(n_847),
.A3(n_837),
.B(n_827),
.Y(n_904)
);

AND2x2_ASAP7_75t_L g905 ( 
.A(n_880),
.B(n_795),
.Y(n_905)
);

INVx1_ASAP7_75t_L g906 ( 
.A(n_868),
.Y(n_906)
);

INVx1_ASAP7_75t_L g907 ( 
.A(n_868),
.Y(n_907)
);

AND2x2_ASAP7_75t_L g908 ( 
.A(n_880),
.B(n_890),
.Y(n_908)
);

AND2x4_ASAP7_75t_L g909 ( 
.A(n_888),
.B(n_826),
.Y(n_909)
);

INVx2_ASAP7_75t_L g910 ( 
.A(n_878),
.Y(n_910)
);

INVx2_ASAP7_75t_L g911 ( 
.A(n_878),
.Y(n_911)
);

OR2x2_ASAP7_75t_L g912 ( 
.A(n_872),
.B(n_867),
.Y(n_912)
);

NOR2xp33_ASAP7_75t_L g913 ( 
.A(n_895),
.B(n_828),
.Y(n_913)
);

HB1xp67_ASAP7_75t_L g914 ( 
.A(n_873),
.Y(n_914)
);

NOR3xp33_ASAP7_75t_L g915 ( 
.A(n_889),
.B(n_865),
.C(n_862),
.Y(n_915)
);

NOR2x1_ASAP7_75t_L g916 ( 
.A(n_871),
.B(n_829),
.Y(n_916)
);

AOI22xp33_ASAP7_75t_L g917 ( 
.A1(n_883),
.A2(n_793),
.B1(n_797),
.B2(n_775),
.Y(n_917)
);

NAND2xp5_ASAP7_75t_L g918 ( 
.A(n_882),
.B(n_769),
.Y(n_918)
);

INVx1_ASAP7_75t_L g919 ( 
.A(n_878),
.Y(n_919)
);

AND2x2_ASAP7_75t_L g920 ( 
.A(n_908),
.B(n_890),
.Y(n_920)
);

AND2x2_ASAP7_75t_L g921 ( 
.A(n_908),
.B(n_893),
.Y(n_921)
);

NOR2xp33_ASAP7_75t_L g922 ( 
.A(n_913),
.B(n_889),
.Y(n_922)
);

INVxp67_ASAP7_75t_SL g923 ( 
.A(n_903),
.Y(n_923)
);

NAND2xp5_ASAP7_75t_L g924 ( 
.A(n_912),
.B(n_882),
.Y(n_924)
);

INVx1_ASAP7_75t_L g925 ( 
.A(n_906),
.Y(n_925)
);

INVx1_ASAP7_75t_L g926 ( 
.A(n_906),
.Y(n_926)
);

NAND2xp5_ASAP7_75t_L g927 ( 
.A(n_912),
.B(n_882),
.Y(n_927)
);

OR2x2_ASAP7_75t_L g928 ( 
.A(n_902),
.B(n_873),
.Y(n_928)
);

INVx1_ASAP7_75t_L g929 ( 
.A(n_907),
.Y(n_929)
);

INVx3_ASAP7_75t_L g930 ( 
.A(n_903),
.Y(n_930)
);

OR2x2_ASAP7_75t_L g931 ( 
.A(n_902),
.B(n_886),
.Y(n_931)
);

AND2x2_ASAP7_75t_L g932 ( 
.A(n_914),
.B(n_916),
.Y(n_932)
);

INVx2_ASAP7_75t_SL g933 ( 
.A(n_903),
.Y(n_933)
);

NAND2xp67_ASAP7_75t_L g934 ( 
.A(n_904),
.B(n_876),
.Y(n_934)
);

OAI22xp33_ASAP7_75t_L g935 ( 
.A1(n_928),
.A2(n_853),
.B1(n_852),
.B2(n_896),
.Y(n_935)
);

NOR2xp33_ASAP7_75t_L g936 ( 
.A(n_922),
.B(n_916),
.Y(n_936)
);

NAND2xp33_ASAP7_75t_SL g937 ( 
.A(n_932),
.B(n_844),
.Y(n_937)
);

NOR2xp33_ASAP7_75t_L g938 ( 
.A(n_934),
.B(n_841),
.Y(n_938)
);

NAND2xp33_ASAP7_75t_SL g939 ( 
.A(n_932),
.B(n_898),
.Y(n_939)
);

NOR4xp25_ASAP7_75t_SL g940 ( 
.A(n_923),
.B(n_854),
.C(n_907),
.D(n_919),
.Y(n_940)
);

NOR2xp33_ASAP7_75t_R g941 ( 
.A(n_921),
.B(n_891),
.Y(n_941)
);

NOR4xp25_ASAP7_75t_SL g942 ( 
.A(n_925),
.B(n_919),
.C(n_886),
.D(n_896),
.Y(n_942)
);

NOR2xp33_ASAP7_75t_L g943 ( 
.A(n_936),
.B(n_926),
.Y(n_943)
);

INVx2_ASAP7_75t_L g944 ( 
.A(n_938),
.Y(n_944)
);

INVx2_ASAP7_75t_L g945 ( 
.A(n_942),
.Y(n_945)
);

AND2x2_ASAP7_75t_L g946 ( 
.A(n_941),
.B(n_921),
.Y(n_946)
);

NAND2xp5_ASAP7_75t_L g947 ( 
.A(n_939),
.B(n_929),
.Y(n_947)
);

INVx1_ASAP7_75t_L g948 ( 
.A(n_935),
.Y(n_948)
);

INVx1_ASAP7_75t_SL g949 ( 
.A(n_937),
.Y(n_949)
);

INVx1_ASAP7_75t_L g950 ( 
.A(n_940),
.Y(n_950)
);

OAI211xp5_ASAP7_75t_L g951 ( 
.A1(n_949),
.A2(n_915),
.B(n_930),
.C(n_933),
.Y(n_951)
);

AOI21xp5_ASAP7_75t_L g952 ( 
.A1(n_943),
.A2(n_933),
.B(n_927),
.Y(n_952)
);

NAND2xp5_ASAP7_75t_L g953 ( 
.A(n_943),
.B(n_924),
.Y(n_953)
);

NAND2xp5_ASAP7_75t_L g954 ( 
.A(n_947),
.B(n_928),
.Y(n_954)
);

INVxp67_ASAP7_75t_SL g955 ( 
.A(n_950),
.Y(n_955)
);

OAI21xp33_ASAP7_75t_L g956 ( 
.A1(n_955),
.A2(n_947),
.B(n_945),
.Y(n_956)
);

NAND2xp5_ASAP7_75t_SL g957 ( 
.A(n_951),
.B(n_944),
.Y(n_957)
);

AND2x4_ASAP7_75t_L g958 ( 
.A(n_954),
.B(n_946),
.Y(n_958)
);

AND2x2_ASAP7_75t_L g959 ( 
.A(n_952),
.B(n_920),
.Y(n_959)
);

INVx1_ASAP7_75t_L g960 ( 
.A(n_958),
.Y(n_960)
);

INVx2_ASAP7_75t_L g961 ( 
.A(n_958),
.Y(n_961)
);

INVx1_ASAP7_75t_L g962 ( 
.A(n_956),
.Y(n_962)
);

NOR2xp33_ASAP7_75t_L g963 ( 
.A(n_957),
.B(n_953),
.Y(n_963)
);

BUFx2_ASAP7_75t_L g964 ( 
.A(n_959),
.Y(n_964)
);

NAND4xp25_ASAP7_75t_L g965 ( 
.A(n_962),
.B(n_948),
.C(n_920),
.D(n_930),
.Y(n_965)
);

AND2x2_ASAP7_75t_L g966 ( 
.A(n_964),
.B(n_930),
.Y(n_966)
);

NAND4xp75_ASAP7_75t_L g967 ( 
.A(n_963),
.B(n_857),
.C(n_876),
.D(n_891),
.Y(n_967)
);

NAND2xp5_ASAP7_75t_L g968 ( 
.A(n_963),
.B(n_931),
.Y(n_968)
);

AOI32xp33_ASAP7_75t_L g969 ( 
.A1(n_960),
.A2(n_892),
.A3(n_917),
.B1(n_780),
.B2(n_909),
.Y(n_969)
);

INVx2_ASAP7_75t_SL g970 ( 
.A(n_961),
.Y(n_970)
);

NAND3xp33_ASAP7_75t_L g971 ( 
.A(n_962),
.B(n_771),
.C(n_931),
.Y(n_971)
);

NAND4xp75_ASAP7_75t_L g972 ( 
.A(n_962),
.B(n_875),
.C(n_884),
.D(n_899),
.Y(n_972)
);

AOI21xp5_ASAP7_75t_L g973 ( 
.A1(n_968),
.A2(n_826),
.B(n_918),
.Y(n_973)
);

NAND4xp75_ASAP7_75t_L g974 ( 
.A(n_970),
.B(n_875),
.C(n_905),
.D(n_897),
.Y(n_974)
);

BUFx2_ASAP7_75t_L g975 ( 
.A(n_966),
.Y(n_975)
);

BUFx2_ASAP7_75t_L g976 ( 
.A(n_965),
.Y(n_976)
);

AOI222xp33_ASAP7_75t_L g977 ( 
.A1(n_971),
.A2(n_797),
.B1(n_793),
.B2(n_799),
.C1(n_805),
.C2(n_808),
.Y(n_977)
);

AOI222xp33_ASAP7_75t_L g978 ( 
.A1(n_967),
.A2(n_799),
.B1(n_800),
.B2(n_808),
.C1(n_807),
.C2(n_805),
.Y(n_978)
);

AOI221xp5_ASAP7_75t_L g979 ( 
.A1(n_969),
.A2(n_818),
.B1(n_807),
.B2(n_800),
.C(n_881),
.Y(n_979)
);

AOI221xp5_ASAP7_75t_SL g980 ( 
.A1(n_972),
.A2(n_881),
.B1(n_897),
.B2(n_899),
.C(n_900),
.Y(n_980)
);

INVx1_ASAP7_75t_L g981 ( 
.A(n_975),
.Y(n_981)
);

INVx1_ASAP7_75t_SL g982 ( 
.A(n_976),
.Y(n_982)
);

AOI22xp5_ASAP7_75t_L g983 ( 
.A1(n_979),
.A2(n_848),
.B1(n_909),
.B2(n_900),
.Y(n_983)
);

NOR2xp67_ASAP7_75t_L g984 ( 
.A(n_973),
.B(n_894),
.Y(n_984)
);

XNOR2x1_ASAP7_75t_L g985 ( 
.A(n_974),
.B(n_848),
.Y(n_985)
);

INVx1_ASAP7_75t_L g986 ( 
.A(n_977),
.Y(n_986)
);

XNOR2xp5_ASAP7_75t_L g987 ( 
.A(n_980),
.B(n_909),
.Y(n_987)
);

CKINVDCx11_ASAP7_75t_R g988 ( 
.A(n_978),
.Y(n_988)
);

NAND3xp33_ASAP7_75t_L g989 ( 
.A(n_981),
.B(n_988),
.C(n_986),
.Y(n_989)
);

NOR2xp33_ASAP7_75t_R g990 ( 
.A(n_982),
.B(n_211),
.Y(n_990)
);

NOR2xp33_ASAP7_75t_R g991 ( 
.A(n_987),
.B(n_214),
.Y(n_991)
);

NAND2xp5_ASAP7_75t_SL g992 ( 
.A(n_984),
.B(n_909),
.Y(n_992)
);

NOR2xp33_ASAP7_75t_R g993 ( 
.A(n_985),
.B(n_217),
.Y(n_993)
);

NAND2xp5_ASAP7_75t_SL g994 ( 
.A(n_983),
.B(n_881),
.Y(n_994)
);

NAND2xp5_ASAP7_75t_L g995 ( 
.A(n_981),
.B(n_905),
.Y(n_995)
);

NAND5xp2_ASAP7_75t_L g996 ( 
.A(n_995),
.B(n_818),
.C(n_835),
.D(n_885),
.E(n_901),
.Y(n_996)
);

AOI22xp5_ASAP7_75t_L g997 ( 
.A1(n_989),
.A2(n_894),
.B1(n_885),
.B2(n_901),
.Y(n_997)
);

XNOR2xp5_ASAP7_75t_L g998 ( 
.A(n_992),
.B(n_218),
.Y(n_998)
);

OAI22x1_ASAP7_75t_L g999 ( 
.A1(n_990),
.A2(n_911),
.B1(n_910),
.B2(n_879),
.Y(n_999)
);

INVx2_ASAP7_75t_L g1000 ( 
.A(n_994),
.Y(n_1000)
);

INVx1_ASAP7_75t_L g1001 ( 
.A(n_991),
.Y(n_1001)
);

INVx1_ASAP7_75t_L g1002 ( 
.A(n_1000),
.Y(n_1002)
);

OR4x2_ASAP7_75t_L g1003 ( 
.A(n_996),
.B(n_998),
.C(n_993),
.D(n_1001),
.Y(n_1003)
);

AOI22x1_ASAP7_75t_L g1004 ( 
.A1(n_999),
.A2(n_809),
.B1(n_804),
.B2(n_911),
.Y(n_1004)
);

INVx1_ASAP7_75t_L g1005 ( 
.A(n_997),
.Y(n_1005)
);

AND2x4_ASAP7_75t_L g1006 ( 
.A(n_1000),
.B(n_879),
.Y(n_1006)
);

CKINVDCx20_ASAP7_75t_R g1007 ( 
.A(n_1002),
.Y(n_1007)
);

OAI22x1_ASAP7_75t_L g1008 ( 
.A1(n_1005),
.A2(n_910),
.B1(n_879),
.B2(n_869),
.Y(n_1008)
);

OAI22xp5_ASAP7_75t_L g1009 ( 
.A1(n_1006),
.A2(n_1004),
.B1(n_1003),
.B2(n_809),
.Y(n_1009)
);

AOI31xp33_ASAP7_75t_L g1010 ( 
.A1(n_1007),
.A2(n_804),
.A3(n_879),
.B(n_869),
.Y(n_1010)
);

AOI31xp33_ASAP7_75t_L g1011 ( 
.A1(n_1009),
.A2(n_869),
.A3(n_817),
.B(n_870),
.Y(n_1011)
);

XOR2xp5_ASAP7_75t_L g1012 ( 
.A(n_1011),
.B(n_1008),
.Y(n_1012)
);

NOR3xp33_ASAP7_75t_L g1013 ( 
.A(n_1010),
.B(n_729),
.C(n_794),
.Y(n_1013)
);

OR2x2_ASAP7_75t_L g1014 ( 
.A(n_1012),
.B(n_796),
.Y(n_1014)
);

INVxp67_ASAP7_75t_L g1015 ( 
.A(n_1013),
.Y(n_1015)
);

NAND2xp5_ASAP7_75t_L g1016 ( 
.A(n_1015),
.B(n_794),
.Y(n_1016)
);

INVx1_ASAP7_75t_L g1017 ( 
.A(n_1014),
.Y(n_1017)
);

OAI221xp5_ASAP7_75t_R g1018 ( 
.A1(n_1017),
.A2(n_1016),
.B1(n_796),
.B2(n_869),
.C(n_817),
.Y(n_1018)
);

AOI211xp5_ASAP7_75t_L g1019 ( 
.A1(n_1018),
.A2(n_874),
.B(n_779),
.C(n_870),
.Y(n_1019)
);


endmodule