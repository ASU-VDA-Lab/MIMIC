module fake_jpeg_31866_n_72 (n_3, n_2, n_1, n_0, n_4, n_6, n_5, n_7, n_72);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_6;
input n_5;
input n_7;

output n_72;

wire n_13;
wire n_21;
wire n_57;
wire n_53;
wire n_33;
wire n_54;
wire n_61;
wire n_45;
wire n_10;
wire n_23;
wire n_69;
wire n_27;
wire n_55;
wire n_64;
wire n_22;
wire n_47;
wire n_51;
wire n_14;
wire n_40;
wire n_19;
wire n_18;
wire n_20;
wire n_59;
wire n_35;
wire n_48;
wire n_68;
wire n_52;
wire n_71;
wire n_46;
wire n_58;
wire n_41;
wire n_60;
wire n_63;
wire n_65;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_16;
wire n_49;
wire n_24;
wire n_28;
wire n_38;
wire n_26;
wire n_44;
wire n_9;
wire n_36;
wire n_11;
wire n_62;
wire n_17;
wire n_31;
wire n_25;
wire n_56;
wire n_67;
wire n_29;
wire n_37;
wire n_43;
wire n_50;
wire n_12;
wire n_32;
wire n_8;
wire n_70;
wire n_15;
wire n_66;

BUFx5_ASAP7_75t_L g8 ( 
.A(n_6),
.Y(n_8)
);

BUFx10_ASAP7_75t_L g9 ( 
.A(n_2),
.Y(n_9)
);

INVx1_ASAP7_75t_L g10 ( 
.A(n_0),
.Y(n_10)
);

INVx1_ASAP7_75t_L g11 ( 
.A(n_3),
.Y(n_11)
);

INVx11_ASAP7_75t_L g12 ( 
.A(n_4),
.Y(n_12)
);

INVx1_ASAP7_75t_L g13 ( 
.A(n_0),
.Y(n_13)
);

BUFx6f_ASAP7_75t_L g14 ( 
.A(n_1),
.Y(n_14)
);

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_4),
.Y(n_15)
);

BUFx6f_ASAP7_75t_L g16 ( 
.A(n_14),
.Y(n_16)
);

INVx11_ASAP7_75t_L g26 ( 
.A(n_16),
.Y(n_26)
);

INVx8_ASAP7_75t_L g17 ( 
.A(n_14),
.Y(n_17)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_17),
.Y(n_25)
);

INVx8_ASAP7_75t_L g18 ( 
.A(n_14),
.Y(n_18)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_18),
.Y(n_27)
);

CKINVDCx16_ASAP7_75t_R g19 ( 
.A(n_10),
.Y(n_19)
);

CKINVDCx14_ASAP7_75t_R g23 ( 
.A(n_19),
.Y(n_23)
);

NOR2xp33_ASAP7_75t_L g20 ( 
.A(n_15),
.B(n_0),
.Y(n_20)
);

NAND2xp5_ASAP7_75t_L g24 ( 
.A(n_20),
.B(n_21),
.Y(n_24)
);

INVx2_ASAP7_75t_L g21 ( 
.A(n_14),
.Y(n_21)
);

AOI22xp33_ASAP7_75t_L g22 ( 
.A1(n_21),
.A2(n_16),
.B1(n_19),
.B2(n_18),
.Y(n_22)
);

AOI22xp5_ASAP7_75t_L g32 ( 
.A1(n_22),
.A2(n_28),
.B1(n_17),
.B2(n_11),
.Y(n_32)
);

AOI22xp33_ASAP7_75t_L g28 ( 
.A1(n_16),
.A2(n_10),
.B1(n_12),
.B2(n_13),
.Y(n_28)
);

OAI22xp33_ASAP7_75t_SL g29 ( 
.A1(n_24),
.A2(n_18),
.B1(n_17),
.B2(n_16),
.Y(n_29)
);

OAI22xp5_ASAP7_75t_L g37 ( 
.A1(n_29),
.A2(n_32),
.B1(n_26),
.B2(n_27),
.Y(n_37)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_22),
.Y(n_30)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_30),
.Y(n_41)
);

AOI22xp5_ASAP7_75t_SL g31 ( 
.A1(n_23),
.A2(n_13),
.B1(n_11),
.B2(n_10),
.Y(n_31)
);

OAI21xp5_ASAP7_75t_SL g38 ( 
.A1(n_31),
.A2(n_11),
.B(n_25),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_SL g33 ( 
.A(n_24),
.B(n_20),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_L g36 ( 
.A(n_33),
.B(n_35),
.Y(n_36)
);

NAND2xp5_ASAP7_75t_L g34 ( 
.A(n_23),
.B(n_9),
.Y(n_34)
);

NAND2xp5_ASAP7_75t_L g40 ( 
.A(n_34),
.B(n_9),
.Y(n_40)
);

OR2x2_ASAP7_75t_L g35 ( 
.A(n_28),
.B(n_15),
.Y(n_35)
);

OAI22xp5_ASAP7_75t_L g43 ( 
.A1(n_37),
.A2(n_32),
.B1(n_30),
.B2(n_34),
.Y(n_43)
);

OAI21xp5_ASAP7_75t_L g47 ( 
.A1(n_38),
.A2(n_12),
.B(n_25),
.Y(n_47)
);

AND2x6_ASAP7_75t_L g39 ( 
.A(n_35),
.B(n_31),
.Y(n_39)
);

XNOR2xp5_ASAP7_75t_L g48 ( 
.A(n_39),
.B(n_40),
.Y(n_48)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_41),
.Y(n_42)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_42),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_L g50 ( 
.A(n_43),
.B(n_44),
.Y(n_50)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_38),
.Y(n_44)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_36),
.Y(n_45)
);

INVxp67_ASAP7_75t_L g49 ( 
.A(n_45),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_39),
.Y(n_46)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_46),
.Y(n_52)
);

MAJIxp5_ASAP7_75t_L g54 ( 
.A(n_47),
.B(n_9),
.C(n_8),
.Y(n_54)
);

MAJx2_ASAP7_75t_L g51 ( 
.A(n_48),
.B(n_27),
.C(n_8),
.Y(n_51)
);

MAJIxp5_ASAP7_75t_L g59 ( 
.A(n_51),
.B(n_9),
.C(n_1),
.Y(n_59)
);

OAI22xp5_ASAP7_75t_L g57 ( 
.A1(n_54),
.A2(n_8),
.B1(n_42),
.B2(n_12),
.Y(n_57)
);

AO21x1_ASAP7_75t_L g55 ( 
.A1(n_50),
.A2(n_47),
.B(n_48),
.Y(n_55)
);

AOI21x1_ASAP7_75t_L g63 ( 
.A1(n_55),
.A2(n_58),
.B(n_3),
.Y(n_63)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_53),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_L g62 ( 
.A(n_56),
.B(n_55),
.Y(n_62)
);

MAJIxp5_ASAP7_75t_L g60 ( 
.A(n_57),
.B(n_59),
.C(n_52),
.Y(n_60)
);

A2O1A1O1Ixp25_ASAP7_75t_L g58 ( 
.A1(n_51),
.A2(n_9),
.B(n_1),
.C(n_2),
.D(n_5),
.Y(n_58)
);

INVxp67_ASAP7_75t_L g65 ( 
.A(n_60),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_58),
.B(n_49),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_L g66 ( 
.A(n_61),
.B(n_62),
.Y(n_66)
);

AOI21xp5_ASAP7_75t_L g64 ( 
.A1(n_63),
.A2(n_5),
.B(n_6),
.Y(n_64)
);

OAI21xp5_ASAP7_75t_L g68 ( 
.A1(n_64),
.A2(n_7),
.B(n_2),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_L g67 ( 
.A(n_66),
.B(n_7),
.Y(n_67)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_67),
.Y(n_69)
);

BUFx24_ASAP7_75t_SL g70 ( 
.A(n_68),
.Y(n_70)
);

AOI221xp5_ASAP7_75t_L g71 ( 
.A1(n_69),
.A2(n_65),
.B1(n_70),
.B2(n_26),
.C(n_9),
.Y(n_71)
);

XOR2xp5_ASAP7_75t_L g72 ( 
.A(n_71),
.B(n_26),
.Y(n_72)
);


endmodule