module fake_jpeg_16253_n_211 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_211);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_211;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_84;
wire n_59;
wire n_98;
wire n_178;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_207;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_57;
wire n_21;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_24;
wire n_44;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_121;
wire n_99;
wire n_130;
wire n_102;
wire n_70;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_189;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

INVx1_ASAP7_75t_L g16 ( 
.A(n_1),
.Y(n_16)
);

BUFx10_ASAP7_75t_L g17 ( 
.A(n_0),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_15),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_1),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_8),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_13),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_15),
.Y(n_22)
);

INVx5_ASAP7_75t_L g23 ( 
.A(n_6),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_5),
.Y(n_24)
);

BUFx3_ASAP7_75t_L g25 ( 
.A(n_2),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_0),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_9),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_14),
.Y(n_28)
);

BUFx5_ASAP7_75t_L g29 ( 
.A(n_3),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_1),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_14),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_0),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_3),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_SL g34 ( 
.A(n_16),
.B(n_2),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_34),
.B(n_35),
.Y(n_48)
);

INVx11_ASAP7_75t_L g35 ( 
.A(n_20),
.Y(n_35)
);

NAND2xp5_ASAP7_75t_L g36 ( 
.A(n_17),
.B(n_2),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_36),
.B(n_38),
.Y(n_55)
);

INVx2_ASAP7_75t_L g37 ( 
.A(n_20),
.Y(n_37)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_37),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g38 ( 
.A(n_17),
.B(n_3),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_L g39 ( 
.A(n_16),
.B(n_4),
.Y(n_39)
);

OAI21xp33_ASAP7_75t_L g58 ( 
.A1(n_39),
.A2(n_27),
.B(n_24),
.Y(n_58)
);

BUFx5_ASAP7_75t_L g40 ( 
.A(n_17),
.Y(n_40)
);

INVx4_ASAP7_75t_L g53 ( 
.A(n_40),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_20),
.Y(n_41)
);

INVx4_ASAP7_75t_L g57 ( 
.A(n_41),
.Y(n_57)
);

BUFx3_ASAP7_75t_L g42 ( 
.A(n_17),
.Y(n_42)
);

INVx5_ASAP7_75t_L g44 ( 
.A(n_42),
.Y(n_44)
);

INVx2_ASAP7_75t_L g43 ( 
.A(n_20),
.Y(n_43)
);

INVx3_ASAP7_75t_L g51 ( 
.A(n_43),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_L g45 ( 
.A(n_36),
.B(n_34),
.Y(n_45)
);

NAND2xp5_ASAP7_75t_L g81 ( 
.A(n_45),
.B(n_46),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_SL g46 ( 
.A(n_34),
.B(n_16),
.Y(n_46)
);

AND2x2_ASAP7_75t_SL g47 ( 
.A(n_36),
.B(n_26),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_47),
.B(n_17),
.Y(n_73)
);

OAI22xp33_ASAP7_75t_L g49 ( 
.A1(n_35),
.A2(n_43),
.B1(n_37),
.B2(n_41),
.Y(n_49)
);

OAI22xp5_ASAP7_75t_SL g70 ( 
.A1(n_49),
.A2(n_35),
.B1(n_23),
.B2(n_41),
.Y(n_70)
);

NAND2xp33_ASAP7_75t_SL g50 ( 
.A(n_38),
.B(n_17),
.Y(n_50)
);

AOI22xp5_ASAP7_75t_SL g69 ( 
.A1(n_50),
.A2(n_23),
.B1(n_19),
.B2(n_33),
.Y(n_69)
);

INVx3_ASAP7_75t_L g52 ( 
.A(n_37),
.Y(n_52)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_52),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_SL g54 ( 
.A(n_39),
.B(n_27),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_SL g62 ( 
.A(n_54),
.B(n_59),
.Y(n_62)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_58),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_L g59 ( 
.A(n_38),
.B(n_26),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_L g60 ( 
.A(n_43),
.B(n_24),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_SL g75 ( 
.A(n_60),
.B(n_61),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_SL g61 ( 
.A(n_35),
.B(n_33),
.Y(n_61)
);

INVx11_ASAP7_75t_L g64 ( 
.A(n_57),
.Y(n_64)
);

BUFx2_ASAP7_75t_L g111 ( 
.A(n_64),
.Y(n_111)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_56),
.Y(n_65)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_65),
.Y(n_104)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_56),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_66),
.B(n_71),
.Y(n_101)
);

INVx2_ASAP7_75t_L g67 ( 
.A(n_44),
.Y(n_67)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_67),
.Y(n_88)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_51),
.Y(n_68)
);

INVx2_ASAP7_75t_L g90 ( 
.A(n_68),
.Y(n_90)
);

XNOR2xp5_ASAP7_75t_L g100 ( 
.A(n_69),
.B(n_73),
.Y(n_100)
);

AOI22xp5_ASAP7_75t_L g109 ( 
.A1(n_70),
.A2(n_19),
.B1(n_30),
.B2(n_32),
.Y(n_109)
);

INVx3_ASAP7_75t_L g71 ( 
.A(n_44),
.Y(n_71)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_51),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_72),
.B(n_74),
.Y(n_102)
);

INVx5_ASAP7_75t_L g74 ( 
.A(n_53),
.Y(n_74)
);

INVxp67_ASAP7_75t_L g76 ( 
.A(n_61),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_SL g105 ( 
.A(n_76),
.B(n_78),
.Y(n_105)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_52),
.Y(n_77)
);

CKINVDCx20_ASAP7_75t_R g92 ( 
.A(n_77),
.Y(n_92)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_60),
.Y(n_78)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_48),
.Y(n_79)
);

HB1xp67_ASAP7_75t_L g99 ( 
.A(n_79),
.Y(n_99)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_48),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_SL g94 ( 
.A(n_80),
.B(n_87),
.Y(n_94)
);

INVx5_ASAP7_75t_L g83 ( 
.A(n_53),
.Y(n_83)
);

INVxp67_ASAP7_75t_L g98 ( 
.A(n_83),
.Y(n_98)
);

INVx2_ASAP7_75t_L g84 ( 
.A(n_57),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g91 ( 
.A(n_84),
.B(n_86),
.Y(n_91)
);

INVx8_ASAP7_75t_L g85 ( 
.A(n_50),
.Y(n_85)
);

AOI22xp5_ASAP7_75t_SL g107 ( 
.A1(n_85),
.A2(n_71),
.B1(n_67),
.B2(n_74),
.Y(n_107)
);

INVx3_ASAP7_75t_L g86 ( 
.A(n_47),
.Y(n_86)
);

CKINVDCx16_ASAP7_75t_R g87 ( 
.A(n_59),
.Y(n_87)
);

O2A1O1Ixp33_ASAP7_75t_SL g89 ( 
.A1(n_85),
.A2(n_55),
.B(n_45),
.C(n_46),
.Y(n_89)
);

OAI21xp5_ASAP7_75t_L g127 ( 
.A1(n_89),
.A2(n_107),
.B(n_31),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_L g93 ( 
.A(n_81),
.B(n_47),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_L g120 ( 
.A(n_93),
.B(n_96),
.Y(n_120)
);

OAI22xp5_ASAP7_75t_SL g95 ( 
.A1(n_63),
.A2(n_69),
.B1(n_86),
.B2(n_81),
.Y(n_95)
);

OAI22xp5_ASAP7_75t_SL g113 ( 
.A1(n_95),
.A2(n_97),
.B1(n_103),
.B2(n_84),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_L g96 ( 
.A(n_75),
.B(n_47),
.Y(n_96)
);

OAI22xp5_ASAP7_75t_SL g97 ( 
.A1(n_76),
.A2(n_55),
.B1(n_23),
.B2(n_41),
.Y(n_97)
);

OAI22xp5_ASAP7_75t_SL g103 ( 
.A1(n_70),
.A2(n_82),
.B1(n_62),
.B2(n_64),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_L g106 ( 
.A(n_82),
.B(n_54),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_L g129 ( 
.A(n_106),
.B(n_108),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_L g108 ( 
.A(n_68),
.B(n_25),
.Y(n_108)
);

OAI22xp5_ASAP7_75t_L g116 ( 
.A1(n_109),
.A2(n_32),
.B1(n_30),
.B2(n_28),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_L g110 ( 
.A(n_83),
.B(n_25),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_L g131 ( 
.A(n_110),
.B(n_42),
.Y(n_131)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_101),
.Y(n_112)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_112),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_SL g148 ( 
.A(n_113),
.B(n_122),
.Y(n_148)
);

INVxp67_ASAP7_75t_L g114 ( 
.A(n_90),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_L g134 ( 
.A(n_114),
.B(n_126),
.Y(n_134)
);

XOR2xp5_ASAP7_75t_L g115 ( 
.A(n_100),
.B(n_40),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_L g138 ( 
.A(n_115),
.B(n_118),
.Y(n_138)
);

AOI22xp5_ASAP7_75t_L g146 ( 
.A1(n_116),
.A2(n_121),
.B1(n_123),
.B2(n_124),
.Y(n_146)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_90),
.Y(n_117)
);

CKINVDCx20_ASAP7_75t_R g145 ( 
.A(n_117),
.Y(n_145)
);

MAJIxp5_ASAP7_75t_L g118 ( 
.A(n_100),
.B(n_42),
.C(n_40),
.Y(n_118)
);

AOI21xp5_ASAP7_75t_L g119 ( 
.A1(n_91),
.A2(n_4),
.B(n_5),
.Y(n_119)
);

A2O1A1Ixp33_ASAP7_75t_SL g144 ( 
.A1(n_119),
.A2(n_124),
.B(n_108),
.C(n_89),
.Y(n_144)
);

AOI22xp5_ASAP7_75t_L g121 ( 
.A1(n_91),
.A2(n_22),
.B1(n_28),
.B2(n_6),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_L g122 ( 
.A(n_99),
.B(n_31),
.Y(n_122)
);

AND2x2_ASAP7_75t_L g123 ( 
.A(n_93),
.B(n_4),
.Y(n_123)
);

AOI22xp5_ASAP7_75t_L g124 ( 
.A1(n_96),
.A2(n_22),
.B1(n_6),
.B2(n_7),
.Y(n_124)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_88),
.Y(n_125)
);

CKINVDCx20_ASAP7_75t_R g153 ( 
.A(n_125),
.Y(n_153)
);

CKINVDCx20_ASAP7_75t_R g126 ( 
.A(n_104),
.Y(n_126)
);

OAI22xp33_ASAP7_75t_SL g143 ( 
.A1(n_127),
.A2(n_133),
.B1(n_21),
.B2(n_92),
.Y(n_143)
);

NOR2xp33_ASAP7_75t_SL g128 ( 
.A(n_94),
.B(n_18),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_L g136 ( 
.A(n_128),
.B(n_132),
.Y(n_136)
);

MAJIxp5_ASAP7_75t_L g130 ( 
.A(n_95),
.B(n_105),
.C(n_106),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_L g141 ( 
.A(n_130),
.B(n_131),
.Y(n_141)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_88),
.Y(n_132)
);

OAI22xp5_ASAP7_75t_L g133 ( 
.A1(n_109),
.A2(n_18),
.B1(n_21),
.B2(n_25),
.Y(n_133)
);

INVxp67_ASAP7_75t_L g135 ( 
.A(n_131),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_SL g155 ( 
.A(n_135),
.B(n_137),
.Y(n_155)
);

NOR3xp33_ASAP7_75t_L g137 ( 
.A(n_119),
.B(n_89),
.C(n_107),
.Y(n_137)
);

INVxp33_ASAP7_75t_L g139 ( 
.A(n_114),
.Y(n_139)
);

CKINVDCx16_ASAP7_75t_R g160 ( 
.A(n_139),
.Y(n_160)
);

INVxp67_ASAP7_75t_L g140 ( 
.A(n_121),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_SL g157 ( 
.A(n_140),
.B(n_142),
.Y(n_157)
);

NOR2xp33_ASAP7_75t_L g142 ( 
.A(n_126),
.B(n_102),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_SL g165 ( 
.A(n_143),
.B(n_147),
.Y(n_165)
);

OAI22xp5_ASAP7_75t_L g156 ( 
.A1(n_144),
.A2(n_149),
.B1(n_129),
.B2(n_130),
.Y(n_156)
);

OR2x2_ASAP7_75t_L g147 ( 
.A(n_129),
.B(n_103),
.Y(n_147)
);

INVxp67_ASAP7_75t_L g149 ( 
.A(n_113),
.Y(n_149)
);

NOR2xp33_ASAP7_75t_L g150 ( 
.A(n_112),
.B(n_98),
.Y(n_150)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_150),
.Y(n_154)
);

O2A1O1Ixp33_ASAP7_75t_L g152 ( 
.A1(n_127),
.A2(n_110),
.B(n_98),
.C(n_97),
.Y(n_152)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_152),
.Y(n_163)
);

AOI22xp5_ASAP7_75t_L g170 ( 
.A1(n_156),
.A2(n_158),
.B1(n_140),
.B2(n_153),
.Y(n_170)
);

OAI22xp5_ASAP7_75t_L g158 ( 
.A1(n_149),
.A2(n_118),
.B1(n_125),
.B2(n_132),
.Y(n_158)
);

AOI322xp5_ASAP7_75t_L g159 ( 
.A1(n_141),
.A2(n_120),
.A3(n_123),
.B1(n_115),
.B2(n_111),
.C1(n_42),
.C2(n_117),
.Y(n_159)
);

NOR2xp33_ASAP7_75t_SL g175 ( 
.A(n_159),
.B(n_161),
.Y(n_175)
);

CKINVDCx20_ASAP7_75t_R g161 ( 
.A(n_134),
.Y(n_161)
);

MAJIxp5_ASAP7_75t_L g162 ( 
.A(n_138),
.B(n_120),
.C(n_123),
.Y(n_162)
);

MAJIxp5_ASAP7_75t_L g173 ( 
.A(n_162),
.B(n_166),
.C(n_167),
.Y(n_173)
);

BUFx2_ASAP7_75t_L g164 ( 
.A(n_145),
.Y(n_164)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_164),
.Y(n_172)
);

MAJIxp5_ASAP7_75t_L g166 ( 
.A(n_138),
.B(n_40),
.C(n_111),
.Y(n_166)
);

XNOR2xp5_ASAP7_75t_L g167 ( 
.A(n_141),
.B(n_29),
.Y(n_167)
);

MAJIxp5_ASAP7_75t_L g168 ( 
.A(n_135),
.B(n_29),
.C(n_10),
.Y(n_168)
);

MAJIxp5_ASAP7_75t_L g177 ( 
.A(n_168),
.B(n_169),
.C(n_146),
.Y(n_177)
);

MAJIxp5_ASAP7_75t_L g169 ( 
.A(n_148),
.B(n_29),
.C(n_10),
.Y(n_169)
);

OAI22xp5_ASAP7_75t_L g188 ( 
.A1(n_170),
.A2(n_171),
.B1(n_178),
.B2(n_179),
.Y(n_188)
);

AOI22xp5_ASAP7_75t_L g171 ( 
.A1(n_157),
.A2(n_153),
.B1(n_147),
.B2(n_151),
.Y(n_171)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_154),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_SL g184 ( 
.A(n_174),
.B(n_176),
.Y(n_184)
);

INVxp67_ASAP7_75t_L g176 ( 
.A(n_155),
.Y(n_176)
);

MAJIxp5_ASAP7_75t_L g186 ( 
.A(n_177),
.B(n_181),
.C(n_162),
.Y(n_186)
);

OAI22xp5_ASAP7_75t_L g178 ( 
.A1(n_165),
.A2(n_146),
.B1(n_151),
.B2(n_145),
.Y(n_178)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_154),
.Y(n_179)
);

HB1xp67_ASAP7_75t_L g180 ( 
.A(n_160),
.Y(n_180)
);

OAI21x1_ASAP7_75t_L g187 ( 
.A1(n_180),
.A2(n_172),
.B(n_136),
.Y(n_187)
);

MAJIxp5_ASAP7_75t_L g181 ( 
.A(n_166),
.B(n_144),
.C(n_152),
.Y(n_181)
);

XNOR2x1_ASAP7_75t_L g182 ( 
.A(n_181),
.B(n_167),
.Y(n_182)
);

AOI22xp5_ASAP7_75t_SL g191 ( 
.A1(n_182),
.A2(n_190),
.B1(n_173),
.B2(n_7),
.Y(n_191)
);

AOI21xp5_ASAP7_75t_SL g183 ( 
.A1(n_176),
.A2(n_163),
.B(n_144),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_L g193 ( 
.A(n_183),
.B(n_185),
.Y(n_193)
);

AOI31xp67_ASAP7_75t_L g185 ( 
.A1(n_177),
.A2(n_144),
.A3(n_163),
.B(n_164),
.Y(n_185)
);

MAJIxp5_ASAP7_75t_L g195 ( 
.A(n_186),
.B(n_189),
.C(n_8),
.Y(n_195)
);

INVx11_ASAP7_75t_L g196 ( 
.A(n_187),
.Y(n_196)
);

MAJIxp5_ASAP7_75t_L g189 ( 
.A(n_173),
.B(n_168),
.C(n_169),
.Y(n_189)
);

OA21x2_ASAP7_75t_L g190 ( 
.A1(n_175),
.A2(n_144),
.B(n_7),
.Y(n_190)
);

AND2x2_ASAP7_75t_L g202 ( 
.A(n_191),
.B(n_192),
.Y(n_202)
);

AOI22xp5_ASAP7_75t_SL g192 ( 
.A1(n_188),
.A2(n_183),
.B1(n_184),
.B2(n_190),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_L g194 ( 
.A(n_184),
.B(n_5),
.Y(n_194)
);

AOI21xp5_ASAP7_75t_L g198 ( 
.A1(n_194),
.A2(n_9),
.B(n_11),
.Y(n_198)
);

OAI221xp5_ASAP7_75t_L g201 ( 
.A1(n_195),
.A2(n_11),
.B1(n_12),
.B2(n_13),
.C(n_194),
.Y(n_201)
);

NAND2xp33_ASAP7_75t_SL g197 ( 
.A(n_185),
.B(n_8),
.Y(n_197)
);

NAND2xp33_ASAP7_75t_L g200 ( 
.A(n_197),
.B(n_9),
.Y(n_200)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_198),
.Y(n_204)
);

AOI21xp5_ASAP7_75t_L g199 ( 
.A1(n_193),
.A2(n_197),
.B(n_196),
.Y(n_199)
);

XNOR2xp5_ASAP7_75t_L g205 ( 
.A(n_199),
.B(n_201),
.Y(n_205)
);

NOR2xp33_ASAP7_75t_L g203 ( 
.A(n_200),
.B(n_193),
.Y(n_203)
);

NOR2xp33_ASAP7_75t_L g208 ( 
.A(n_203),
.B(n_206),
.Y(n_208)
);

INVxp67_ASAP7_75t_L g206 ( 
.A(n_202),
.Y(n_206)
);

INVxp67_ASAP7_75t_L g207 ( 
.A(n_206),
.Y(n_207)
);

OR2x2_ASAP7_75t_L g209 ( 
.A(n_207),
.B(n_192),
.Y(n_209)
);

XNOR2xp5_ASAP7_75t_L g211 ( 
.A(n_209),
.B(n_210),
.Y(n_211)
);

OAI321xp33_ASAP7_75t_L g210 ( 
.A1(n_208),
.A2(n_205),
.A3(n_196),
.B1(n_204),
.B2(n_191),
.C(n_195),
.Y(n_210)
);


endmodule