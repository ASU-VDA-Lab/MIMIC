module fake_jpeg_9548_n_204 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_204);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_204;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_24;
wire n_44;
wire n_143;
wire n_202;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_161;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_189;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_140;
wire n_82;
wire n_128;
wire n_118;
wire n_96;

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_10),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_14),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_12),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_10),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_0),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_12),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_9),
.Y(n_21)
);

INVx3_ASAP7_75t_L g22 ( 
.A(n_1),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_13),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_14),
.Y(n_24)
);

BUFx12_ASAP7_75t_L g25 ( 
.A(n_3),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_6),
.Y(n_26)
);

BUFx12f_ASAP7_75t_L g27 ( 
.A(n_0),
.Y(n_27)
);

CKINVDCx16_ASAP7_75t_R g28 ( 
.A(n_1),
.Y(n_28)
);

BUFx24_ASAP7_75t_L g29 ( 
.A(n_9),
.Y(n_29)
);

INVx11_ASAP7_75t_L g30 ( 
.A(n_11),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_2),
.Y(n_31)
);

NOR2xp33_ASAP7_75t_L g32 ( 
.A(n_16),
.B(n_0),
.Y(n_32)
);

NOR2xp33_ASAP7_75t_SL g62 ( 
.A(n_32),
.B(n_35),
.Y(n_62)
);

CKINVDCx12_ASAP7_75t_R g33 ( 
.A(n_20),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_L g51 ( 
.A(n_33),
.B(n_34),
.Y(n_51)
);

INVx2_ASAP7_75t_L g34 ( 
.A(n_30),
.Y(n_34)
);

NAND2xp5_ASAP7_75t_L g35 ( 
.A(n_18),
.B(n_1),
.Y(n_35)
);

BUFx10_ASAP7_75t_L g36 ( 
.A(n_27),
.Y(n_36)
);

BUFx12f_ASAP7_75t_L g50 ( 
.A(n_36),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_30),
.Y(n_37)
);

INVx3_ASAP7_75t_L g44 ( 
.A(n_37),
.Y(n_44)
);

INVx2_ASAP7_75t_L g38 ( 
.A(n_30),
.Y(n_38)
);

INVx8_ASAP7_75t_L g60 ( 
.A(n_38),
.Y(n_60)
);

BUFx3_ASAP7_75t_L g39 ( 
.A(n_29),
.Y(n_39)
);

INVx4_ASAP7_75t_L g52 ( 
.A(n_39),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g40 ( 
.A(n_16),
.B(n_2),
.Y(n_40)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_40),
.Y(n_49)
);

INVx2_ASAP7_75t_R g41 ( 
.A(n_29),
.Y(n_41)
);

AND2x2_ASAP7_75t_L g57 ( 
.A(n_41),
.B(n_3),
.Y(n_57)
);

NAND2xp33_ASAP7_75t_SL g42 ( 
.A(n_25),
.B(n_2),
.Y(n_42)
);

OR2x2_ASAP7_75t_SL g48 ( 
.A(n_42),
.B(n_41),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_37),
.Y(n_43)
);

INVx5_ASAP7_75t_L g81 ( 
.A(n_43),
.Y(n_81)
);

OAI22xp33_ASAP7_75t_SL g45 ( 
.A1(n_34),
.A2(n_22),
.B1(n_18),
.B2(n_19),
.Y(n_45)
);

AOI22xp33_ASAP7_75t_L g75 ( 
.A1(n_45),
.A2(n_29),
.B1(n_37),
.B2(n_27),
.Y(n_75)
);

AOI22xp33_ASAP7_75t_SL g46 ( 
.A1(n_41),
.A2(n_22),
.B1(n_28),
.B2(n_18),
.Y(n_46)
);

AOI22xp33_ASAP7_75t_SL g64 ( 
.A1(n_46),
.A2(n_47),
.B1(n_26),
.B2(n_21),
.Y(n_64)
);

AOI22xp33_ASAP7_75t_SL g47 ( 
.A1(n_41),
.A2(n_22),
.B1(n_28),
.B2(n_19),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_48),
.B(n_55),
.Y(n_67)
);

AOI22xp33_ASAP7_75t_L g53 ( 
.A1(n_35),
.A2(n_17),
.B1(n_16),
.B2(n_19),
.Y(n_53)
);

OAI22xp5_ASAP7_75t_L g65 ( 
.A1(n_53),
.A2(n_59),
.B1(n_61),
.B2(n_24),
.Y(n_65)
);

MAJIxp5_ASAP7_75t_L g54 ( 
.A(n_36),
.B(n_17),
.C(n_31),
.Y(n_54)
);

MAJIxp5_ASAP7_75t_L g66 ( 
.A(n_54),
.B(n_24),
.C(n_23),
.Y(n_66)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_32),
.Y(n_55)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_40),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_56),
.B(n_58),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_SL g63 ( 
.A(n_57),
.B(n_29),
.Y(n_63)
);

CKINVDCx20_ASAP7_75t_R g58 ( 
.A(n_33),
.Y(n_58)
);

AOI22xp5_ASAP7_75t_L g59 ( 
.A1(n_38),
.A2(n_17),
.B1(n_31),
.B2(n_15),
.Y(n_59)
);

OAI22xp5_ASAP7_75t_L g61 ( 
.A1(n_42),
.A2(n_15),
.B1(n_21),
.B2(n_26),
.Y(n_61)
);

AND2x2_ASAP7_75t_L g94 ( 
.A(n_63),
.B(n_66),
.Y(n_94)
);

AOI22xp33_ASAP7_75t_SL g89 ( 
.A1(n_64),
.A2(n_44),
.B1(n_81),
.B2(n_73),
.Y(n_89)
);

XNOR2xp5_ASAP7_75t_L g93 ( 
.A(n_65),
.B(n_27),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_L g68 ( 
.A(n_62),
.B(n_27),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_L g82 ( 
.A(n_68),
.B(n_70),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_L g70 ( 
.A(n_62),
.B(n_27),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_49),
.B(n_23),
.Y(n_71)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_71),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_49),
.B(n_20),
.Y(n_72)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_72),
.Y(n_86)
);

INVx2_ASAP7_75t_L g73 ( 
.A(n_60),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_73),
.B(n_76),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_55),
.B(n_11),
.Y(n_74)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_74),
.Y(n_96)
);

OAI22xp5_ASAP7_75t_SL g101 ( 
.A1(n_75),
.A2(n_36),
.B1(n_25),
.B2(n_50),
.Y(n_101)
);

CKINVDCx20_ASAP7_75t_R g76 ( 
.A(n_59),
.Y(n_76)
);

NOR3xp33_ASAP7_75t_L g77 ( 
.A(n_61),
.B(n_39),
.C(n_29),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_77),
.B(n_60),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_56),
.B(n_13),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_SL g95 ( 
.A(n_78),
.B(n_80),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_SL g79 ( 
.A(n_57),
.B(n_37),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_L g88 ( 
.A(n_79),
.B(n_57),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_54),
.B(n_25),
.Y(n_80)
);

OA22x2_ASAP7_75t_L g85 ( 
.A1(n_76),
.A2(n_44),
.B1(n_48),
.B2(n_81),
.Y(n_85)
);

AOI22xp5_ASAP7_75t_SL g114 ( 
.A1(n_85),
.A2(n_89),
.B1(n_97),
.B2(n_101),
.Y(n_114)
);

OAI21xp5_ASAP7_75t_SL g108 ( 
.A1(n_87),
.A2(n_88),
.B(n_90),
.Y(n_108)
);

NAND2x1p5_ASAP7_75t_L g90 ( 
.A(n_79),
.B(n_39),
.Y(n_90)
);

AOI22xp5_ASAP7_75t_L g91 ( 
.A1(n_67),
.A2(n_51),
.B1(n_52),
.B2(n_43),
.Y(n_91)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_91),
.Y(n_119)
);

BUFx3_ASAP7_75t_L g92 ( 
.A(n_80),
.Y(n_92)
);

INVxp67_ASAP7_75t_L g118 ( 
.A(n_92),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_SL g103 ( 
.A(n_93),
.B(n_99),
.Y(n_103)
);

AOI22xp5_ASAP7_75t_L g97 ( 
.A1(n_67),
.A2(n_52),
.B1(n_36),
.B2(n_58),
.Y(n_97)
);

AND2x2_ASAP7_75t_L g98 ( 
.A(n_63),
.B(n_36),
.Y(n_98)
);

XNOR2x1_ASAP7_75t_SL g120 ( 
.A(n_98),
.B(n_100),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_66),
.B(n_50),
.Y(n_99)
);

AND2x2_ASAP7_75t_L g100 ( 
.A(n_68),
.B(n_36),
.Y(n_100)
);

CKINVDCx20_ASAP7_75t_R g102 ( 
.A(n_69),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_L g106 ( 
.A(n_102),
.B(n_69),
.Y(n_106)
);

CKINVDCx20_ASAP7_75t_R g104 ( 
.A(n_83),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_SL g140 ( 
.A(n_104),
.B(n_105),
.Y(n_140)
);

CKINVDCx20_ASAP7_75t_R g105 ( 
.A(n_82),
.Y(n_105)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_106),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_L g107 ( 
.A(n_82),
.B(n_70),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_L g138 ( 
.A(n_107),
.B(n_110),
.Y(n_138)
);

HB1xp67_ASAP7_75t_L g109 ( 
.A(n_90),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_L g133 ( 
.A(n_109),
.B(n_111),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_L g110 ( 
.A(n_100),
.B(n_65),
.Y(n_110)
);

CKINVDCx20_ASAP7_75t_R g111 ( 
.A(n_100),
.Y(n_111)
);

CKINVDCx20_ASAP7_75t_R g112 ( 
.A(n_91),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_L g135 ( 
.A(n_112),
.B(n_113),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_SL g113 ( 
.A(n_84),
.B(n_72),
.Y(n_113)
);

AOI22xp5_ASAP7_75t_SL g115 ( 
.A1(n_90),
.A2(n_71),
.B1(n_25),
.B2(n_78),
.Y(n_115)
);

OAI22xp5_ASAP7_75t_L g131 ( 
.A1(n_115),
.A2(n_121),
.B1(n_10),
.B2(n_5),
.Y(n_131)
);

CKINVDCx20_ASAP7_75t_R g116 ( 
.A(n_97),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_L g136 ( 
.A(n_116),
.B(n_117),
.Y(n_136)
);

CKINVDCx20_ASAP7_75t_R g117 ( 
.A(n_98),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_SL g121 ( 
.A(n_86),
.B(n_74),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_L g122 ( 
.A(n_96),
.B(n_50),
.Y(n_122)
);

AOI22xp33_ASAP7_75t_L g124 ( 
.A1(n_122),
.A2(n_85),
.B1(n_88),
.B2(n_98),
.Y(n_124)
);

OAI22xp5_ASAP7_75t_L g123 ( 
.A1(n_114),
.A2(n_85),
.B1(n_92),
.B2(n_93),
.Y(n_123)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_123),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_L g142 ( 
.A(n_124),
.B(n_125),
.Y(n_142)
);

A2O1A1O1Ixp25_ASAP7_75t_L g125 ( 
.A1(n_120),
.A2(n_85),
.B(n_94),
.C(n_95),
.D(n_101),
.Y(n_125)
);

AOI21xp5_ASAP7_75t_L g126 ( 
.A1(n_120),
.A2(n_94),
.B(n_25),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_L g143 ( 
.A(n_126),
.B(n_127),
.Y(n_143)
);

INVx1_ASAP7_75t_SL g127 ( 
.A(n_110),
.Y(n_127)
);

AOI21xp5_ASAP7_75t_SL g128 ( 
.A1(n_108),
.A2(n_94),
.B(n_50),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_L g153 ( 
.A(n_128),
.B(n_132),
.Y(n_153)
);

AOI22xp5_ASAP7_75t_L g129 ( 
.A1(n_119),
.A2(n_3),
.B1(n_4),
.B2(n_5),
.Y(n_129)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_129),
.Y(n_146)
);

MAJIxp5_ASAP7_75t_L g130 ( 
.A(n_103),
.B(n_4),
.C(n_5),
.Y(n_130)
);

MAJIxp5_ASAP7_75t_L g149 ( 
.A(n_130),
.B(n_139),
.C(n_107),
.Y(n_149)
);

NOR2xp33_ASAP7_75t_SL g145 ( 
.A(n_131),
.B(n_115),
.Y(n_145)
);

AOI22xp5_ASAP7_75t_SL g132 ( 
.A1(n_119),
.A2(n_4),
.B1(n_6),
.B2(n_7),
.Y(n_132)
);

OAI22xp5_ASAP7_75t_L g134 ( 
.A1(n_114),
.A2(n_6),
.B1(n_7),
.B2(n_8),
.Y(n_134)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_134),
.Y(n_147)
);

XOR2xp5_ASAP7_75t_L g139 ( 
.A(n_108),
.B(n_9),
.Y(n_139)
);

BUFx2_ASAP7_75t_L g144 ( 
.A(n_137),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_L g157 ( 
.A(n_144),
.B(n_145),
.Y(n_157)
);

CKINVDCx20_ASAP7_75t_R g148 ( 
.A(n_140),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_L g159 ( 
.A(n_148),
.B(n_149),
.Y(n_159)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_136),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_L g162 ( 
.A(n_150),
.B(n_151),
.Y(n_162)
);

CKINVDCx20_ASAP7_75t_R g151 ( 
.A(n_135),
.Y(n_151)
);

NOR2x1_ASAP7_75t_L g152 ( 
.A(n_127),
.B(n_104),
.Y(n_152)
);

OAI21xp5_ASAP7_75t_L g166 ( 
.A1(n_152),
.A2(n_133),
.B(n_132),
.Y(n_166)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_138),
.Y(n_154)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_154),
.Y(n_156)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_138),
.Y(n_155)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_155),
.Y(n_160)
);

XNOR2xp5_ASAP7_75t_L g158 ( 
.A(n_142),
.B(n_126),
.Y(n_158)
);

MAJIxp5_ASAP7_75t_L g173 ( 
.A(n_158),
.B(n_161),
.C(n_164),
.Y(n_173)
);

XNOR2xp5_ASAP7_75t_L g161 ( 
.A(n_143),
.B(n_125),
.Y(n_161)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_152),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_SL g169 ( 
.A(n_163),
.B(n_165),
.Y(n_169)
);

XNOR2xp5_ASAP7_75t_L g164 ( 
.A(n_149),
.B(n_123),
.Y(n_164)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_144),
.Y(n_165)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_166),
.Y(n_175)
);

BUFx12f_ASAP7_75t_SL g167 ( 
.A(n_150),
.Y(n_167)
);

AOI21xp5_ASAP7_75t_L g174 ( 
.A1(n_167),
.A2(n_118),
.B(n_137),
.Y(n_174)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_148),
.Y(n_168)
);

NOR2xp33_ASAP7_75t_L g171 ( 
.A(n_168),
.B(n_151),
.Y(n_171)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_162),
.Y(n_170)
);

AOI21xp5_ASAP7_75t_L g185 ( 
.A1(n_170),
.A2(n_171),
.B(n_176),
.Y(n_185)
);

AOI22xp33_ASAP7_75t_SL g172 ( 
.A1(n_167),
.A2(n_141),
.B1(n_146),
.B2(n_112),
.Y(n_172)
);

OAI22xp5_ASAP7_75t_SL g181 ( 
.A1(n_172),
.A2(n_178),
.B1(n_156),
.B2(n_147),
.Y(n_181)
);

OAI21xp5_ASAP7_75t_L g183 ( 
.A1(n_174),
.A2(n_118),
.B(n_129),
.Y(n_183)
);

NOR2xp33_ASAP7_75t_L g176 ( 
.A(n_157),
.B(n_146),
.Y(n_176)
);

XNOR2xp5_ASAP7_75t_L g177 ( 
.A(n_164),
.B(n_128),
.Y(n_177)
);

OAI322xp33_ASAP7_75t_L g182 ( 
.A1(n_177),
.A2(n_158),
.A3(n_161),
.B1(n_111),
.B2(n_117),
.C1(n_105),
.C2(n_153),
.Y(n_182)
);

OAI22xp5_ASAP7_75t_L g178 ( 
.A1(n_166),
.A2(n_141),
.B1(n_147),
.B2(n_116),
.Y(n_178)
);

NOR2xp67_ASAP7_75t_L g179 ( 
.A(n_170),
.B(n_159),
.Y(n_179)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_179),
.Y(n_188)
);

OAI31xp33_ASAP7_75t_L g180 ( 
.A1(n_175),
.A2(n_155),
.A3(n_154),
.B(n_160),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_L g190 ( 
.A(n_180),
.B(n_186),
.Y(n_190)
);

NOR2xp33_ASAP7_75t_L g187 ( 
.A(n_181),
.B(n_184),
.Y(n_187)
);

XNOR2xp5_ASAP7_75t_L g192 ( 
.A(n_182),
.B(n_183),
.Y(n_192)
);

AOI22xp5_ASAP7_75t_L g184 ( 
.A1(n_177),
.A2(n_145),
.B1(n_139),
.B2(n_130),
.Y(n_184)
);

NAND4xp25_ASAP7_75t_L g186 ( 
.A(n_174),
.B(n_7),
.C(n_8),
.D(n_169),
.Y(n_186)
);

NOR2xp33_ASAP7_75t_L g189 ( 
.A(n_185),
.B(n_173),
.Y(n_189)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_189),
.Y(n_195)
);

HB1xp67_ASAP7_75t_L g191 ( 
.A(n_180),
.Y(n_191)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_191),
.Y(n_196)
);

INVx11_ASAP7_75t_L g193 ( 
.A(n_191),
.Y(n_193)
);

NOR2xp33_ASAP7_75t_L g199 ( 
.A(n_193),
.B(n_194),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_L g194 ( 
.A(n_190),
.B(n_188),
.Y(n_194)
);

AOI21xp5_ASAP7_75t_L g197 ( 
.A1(n_187),
.A2(n_183),
.B(n_173),
.Y(n_197)
);

XOR2xp5_ASAP7_75t_L g200 ( 
.A(n_197),
.B(n_193),
.Y(n_200)
);

AOI22xp5_ASAP7_75t_L g198 ( 
.A1(n_196),
.A2(n_192),
.B1(n_184),
.B2(n_8),
.Y(n_198)
);

OAI22xp5_ASAP7_75t_L g202 ( 
.A1(n_198),
.A2(n_195),
.B1(n_197),
.B2(n_200),
.Y(n_202)
);

NAND2xp5_ASAP7_75t_L g201 ( 
.A(n_200),
.B(n_199),
.Y(n_201)
);

INVxp67_ASAP7_75t_L g203 ( 
.A(n_201),
.Y(n_203)
);

XNOR2xp5_ASAP7_75t_L g204 ( 
.A(n_203),
.B(n_202),
.Y(n_204)
);


endmodule