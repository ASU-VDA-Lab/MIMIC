module fake_aes_3901_n_516 (n_53, n_67, n_45, n_20, n_2, n_38, n_44, n_64, n_54, n_62, n_36, n_47, n_37, n_69, n_34, n_5, n_23, n_8, n_28, n_31, n_22, n_46, n_48, n_58, n_57, n_11, n_25, n_16, n_26, n_13, n_30, n_33, n_50, n_52, n_49, n_59, n_73, n_3, n_18, n_60, n_66, n_32, n_0, n_41, n_1, n_35, n_55, n_65, n_12, n_9, n_70, n_17, n_63, n_14, n_10, n_15, n_56, n_71, n_42, n_24, n_19, n_61, n_21, n_6, n_4, n_74, n_72, n_51, n_29, n_43, n_7, n_68, n_40, n_27, n_39, n_516);
input n_53;
input n_67;
input n_45;
input n_20;
input n_2;
input n_38;
input n_44;
input n_64;
input n_54;
input n_62;
input n_36;
input n_47;
input n_37;
input n_69;
input n_34;
input n_5;
input n_23;
input n_8;
input n_28;
input n_31;
input n_22;
input n_46;
input n_48;
input n_58;
input n_57;
input n_11;
input n_25;
input n_16;
input n_26;
input n_13;
input n_30;
input n_33;
input n_50;
input n_52;
input n_49;
input n_59;
input n_73;
input n_3;
input n_18;
input n_60;
input n_66;
input n_32;
input n_0;
input n_41;
input n_1;
input n_35;
input n_55;
input n_65;
input n_12;
input n_9;
input n_70;
input n_17;
input n_63;
input n_14;
input n_10;
input n_15;
input n_56;
input n_71;
input n_42;
input n_24;
input n_19;
input n_61;
input n_21;
input n_6;
input n_4;
input n_74;
input n_72;
input n_51;
input n_29;
input n_43;
input n_7;
input n_68;
input n_40;
input n_27;
input n_39;
output n_516;
wire n_117;
wire n_361;
wire n_513;
wire n_185;
wire n_407;
wire n_284;
wire n_278;
wire n_500;
wire n_114;
wire n_94;
wire n_125;
wire n_431;
wire n_484;
wire n_161;
wire n_496;
wire n_177;
wire n_130;
wire n_189;
wire n_311;
wire n_292;
wire n_309;
wire n_160;
wire n_154;
wire n_328;
wire n_468;
wire n_229;
wire n_336;
wire n_464;
wire n_448;
wire n_348;
wire n_252;
wire n_152;
wire n_113;
wire n_353;
wire n_206;
wire n_288;
wire n_383;
wire n_400;
wire n_296;
wire n_157;
wire n_79;
wire n_202;
wire n_386;
wire n_432;
wire n_142;
wire n_232;
wire n_462;
wire n_316;
wire n_211;
wire n_334;
wire n_389;
wire n_436;
wire n_275;
wire n_463;
wire n_131;
wire n_112;
wire n_205;
wire n_330;
wire n_162;
wire n_387;
wire n_163;
wire n_476;
wire n_105;
wire n_227;
wire n_384;
wire n_434;
wire n_231;
wire n_452;
wire n_298;
wire n_411;
wire n_144;
wire n_183;
wire n_489;
wire n_199;
wire n_351;
wire n_83;
wire n_401;
wire n_100;
wire n_305;
wire n_461;
wire n_228;
wire n_345;
wire n_360;
wire n_236;
wire n_340;
wire n_481;
wire n_443;
wire n_150;
wire n_373;
wire n_301;
wire n_222;
wire n_234;
wire n_465;
wire n_366;
wire n_286;
wire n_190;
wire n_246;
wire n_321;
wire n_324;
wire n_392;
wire n_279;
wire n_303;
wire n_437;
wire n_512;
wire n_326;
wire n_289;
wire n_333;
wire n_249;
wire n_244;
wire n_119;
wire n_141;
wire n_479;
wire n_97;
wire n_167;
wire n_447;
wire n_171;
wire n_196;
wire n_192;
wire n_502;
wire n_312;
wire n_455;
wire n_137;
wire n_511;
wire n_277;
wire n_467;
wire n_367;
wire n_85;
wire n_250;
wire n_314;
wire n_237;
wire n_181;
wire n_101;
wire n_255;
wire n_426;
wire n_91;
wire n_108;
wire n_116;
wire n_230;
wire n_209;
wire n_274;
wire n_282;
wire n_319;
wire n_499;
wire n_417;
wire n_241;
wire n_95;
wire n_238;
wire n_318;
wire n_471;
wire n_293;
wire n_506;
wire n_135;
wire n_393;
wire n_247;
wire n_490;
wire n_381;
wire n_304;
wire n_399;
wire n_294;
wire n_459;
wire n_313;
wire n_210;
wire n_184;
wire n_322;
wire n_310;
wire n_191;
wire n_307;
wire n_474;
wire n_354;
wire n_402;
wire n_413;
wire n_391;
wire n_427;
wire n_460;
wire n_478;
wire n_243;
wire n_235;
wire n_415;
wire n_394;
wire n_482;
wire n_442;
wire n_331;
wire n_485;
wire n_352;
wire n_268;
wire n_174;
wire n_501;
wire n_248;
wire n_299;
wire n_89;
wire n_338;
wire n_256;
wire n_77;
wire n_404;
wire n_369;
wire n_509;
wire n_172;
wire n_329;
wire n_251;
wire n_218;
wire n_507;
wire n_271;
wire n_302;
wire n_466;
wire n_270;
wire n_362;
wire n_153;
wire n_259;
wire n_308;
wire n_93;
wire n_412;
wire n_140;
wire n_207;
wire n_224;
wire n_96;
wire n_219;
wire n_475;
wire n_133;
wire n_149;
wire n_81;
wire n_214;
wire n_204;
wire n_430;
wire n_88;
wire n_450;
wire n_107;
wire n_403;
wire n_254;
wire n_262;
wire n_239;
wire n_439;
wire n_87;
wire n_379;
wire n_98;
wire n_276;
wire n_320;
wire n_285;
wire n_195;
wire n_165;
wire n_446;
wire n_420;
wire n_342;
wire n_423;
wire n_370;
wire n_217;
wire n_139;
wire n_388;
wire n_454;
wire n_193;
wire n_273;
wire n_505;
wire n_390;
wire n_120;
wire n_514;
wire n_486;
wire n_245;
wire n_90;
wire n_357;
wire n_260;
wire n_78;
wire n_201;
wire n_197;
wire n_317;
wire n_416;
wire n_374;
wire n_111;
wire n_265;
wire n_264;
wire n_200;
wire n_208;
wire n_126;
wire n_178;
wire n_118;
wire n_365;
wire n_179;
wire n_315;
wire n_363;
wire n_409;
wire n_86;
wire n_143;
wire n_295;
wire n_263;
wire n_166;
wire n_495;
wire n_186;
wire n_364;
wire n_428;
wire n_75;
wire n_376;
wire n_344;
wire n_136;
wire n_503;
wire n_283;
wire n_76;
wire n_435;
wire n_216;
wire n_147;
wire n_148;
wire n_212;
wire n_472;
wire n_92;
wire n_419;
wire n_396;
wire n_168;
wire n_477;
wire n_508;
wire n_398;
wire n_445;
wire n_438;
wire n_134;
wire n_429;
wire n_488;
wire n_233;
wire n_82;
wire n_106;
wire n_440;
wire n_173;
wire n_422;
wire n_327;
wire n_325;
wire n_349;
wire n_498;
wire n_225;
wire n_220;
wire n_358;
wire n_267;
wire n_221;
wire n_456;
wire n_203;
wire n_102;
wire n_449;
wire n_115;
wire n_80;
wire n_300;
wire n_158;
wire n_121;
wire n_497;
wire n_339;
wire n_240;
wire n_378;
wire n_359;
wire n_346;
wire n_103;
wire n_180;
wire n_441;
wire n_104;
wire n_335;
wire n_272;
wire n_146;
wire n_397;
wire n_306;
wire n_215;
wire n_242;
wire n_155;
wire n_198;
wire n_169;
wire n_424;
wire n_156;
wire n_124;
wire n_297;
wire n_128;
wire n_129;
wire n_410;
wire n_188;
wire n_377;
wire n_510;
wire n_343;
wire n_127;
wire n_291;
wire n_170;
wire n_504;
wire n_458;
wire n_493;
wire n_418;
wire n_380;
wire n_356;
wire n_281;
wire n_341;
wire n_470;
wire n_122;
wire n_187;
wire n_375;
wire n_138;
wire n_487;
wire n_451;
wire n_371;
wire n_323;
wire n_473;
wire n_347;
wire n_258;
wire n_253;
wire n_515;
wire n_84;
wire n_266;
wire n_213;
wire n_182;
wire n_492;
wire n_368;
wire n_355;
wire n_226;
wire n_382;
wire n_159;
wire n_337;
wire n_444;
wire n_176;
wire n_469;
wire n_123;
wire n_457;
wire n_223;
wire n_494;
wire n_480;
wire n_372;
wire n_453;
wire n_194;
wire n_287;
wire n_110;
wire n_261;
wire n_425;
wire n_332;
wire n_414;
wire n_350;
wire n_433;
wire n_164;
wire n_421;
wire n_175;
wire n_145;
wire n_483;
wire n_408;
wire n_290;
wire n_405;
wire n_280;
wire n_132;
wire n_99;
wire n_109;
wire n_395;
wire n_406;
wire n_491;
wire n_151;
wire n_385;
wire n_257;
wire n_269;
INVxp33_ASAP7_75t_SL g75 ( .A(n_15), .Y(n_75) );
INVx1_ASAP7_75t_L g76 ( .A(n_39), .Y(n_76) );
INVx1_ASAP7_75t_L g77 ( .A(n_17), .Y(n_77) );
HB1xp67_ASAP7_75t_L g78 ( .A(n_24), .Y(n_78) );
INVx1_ASAP7_75t_L g79 ( .A(n_53), .Y(n_79) );
INVx2_ASAP7_75t_L g80 ( .A(n_43), .Y(n_80) );
BUFx3_ASAP7_75t_L g81 ( .A(n_17), .Y(n_81) );
INVx1_ASAP7_75t_L g82 ( .A(n_6), .Y(n_82) );
INVx1_ASAP7_75t_L g83 ( .A(n_28), .Y(n_83) );
INVx1_ASAP7_75t_L g84 ( .A(n_0), .Y(n_84) );
INVx1_ASAP7_75t_L g85 ( .A(n_71), .Y(n_85) );
INVx1_ASAP7_75t_L g86 ( .A(n_61), .Y(n_86) );
INVx1_ASAP7_75t_L g87 ( .A(n_47), .Y(n_87) );
CKINVDCx5p33_ASAP7_75t_R g88 ( .A(n_67), .Y(n_88) );
INVx1_ASAP7_75t_L g89 ( .A(n_36), .Y(n_89) );
INVx2_ASAP7_75t_L g90 ( .A(n_33), .Y(n_90) );
INVx1_ASAP7_75t_L g91 ( .A(n_13), .Y(n_91) );
INVxp67_ASAP7_75t_SL g92 ( .A(n_73), .Y(n_92) );
BUFx6f_ASAP7_75t_L g93 ( .A(n_11), .Y(n_93) );
INVx1_ASAP7_75t_L g94 ( .A(n_66), .Y(n_94) );
INVxp33_ASAP7_75t_SL g95 ( .A(n_29), .Y(n_95) );
CKINVDCx20_ASAP7_75t_R g96 ( .A(n_20), .Y(n_96) );
INVxp33_ASAP7_75t_L g97 ( .A(n_51), .Y(n_97) );
INVx1_ASAP7_75t_L g98 ( .A(n_45), .Y(n_98) );
NOR2xp67_ASAP7_75t_L g99 ( .A(n_15), .B(n_55), .Y(n_99) );
INVx2_ASAP7_75t_L g100 ( .A(n_56), .Y(n_100) );
INVx2_ASAP7_75t_L g101 ( .A(n_57), .Y(n_101) );
INVxp33_ASAP7_75t_L g102 ( .A(n_35), .Y(n_102) );
INVx1_ASAP7_75t_L g103 ( .A(n_26), .Y(n_103) );
INVx1_ASAP7_75t_L g104 ( .A(n_9), .Y(n_104) );
INVx1_ASAP7_75t_L g105 ( .A(n_30), .Y(n_105) );
INVx1_ASAP7_75t_L g106 ( .A(n_10), .Y(n_106) );
INVx1_ASAP7_75t_L g107 ( .A(n_70), .Y(n_107) );
CKINVDCx5p33_ASAP7_75t_R g108 ( .A(n_58), .Y(n_108) );
INVx2_ASAP7_75t_L g109 ( .A(n_80), .Y(n_109) );
AND2x4_ASAP7_75t_L g110 ( .A(n_81), .B(n_0), .Y(n_110) );
INVx1_ASAP7_75t_SL g111 ( .A(n_96), .Y(n_111) );
INVx2_ASAP7_75t_L g112 ( .A(n_80), .Y(n_112) );
NAND2xp5_ASAP7_75t_L g113 ( .A(n_78), .B(n_1), .Y(n_113) );
INVx3_ASAP7_75t_L g114 ( .A(n_81), .Y(n_114) );
INVx1_ASAP7_75t_L g115 ( .A(n_81), .Y(n_115) );
INVx1_ASAP7_75t_L g116 ( .A(n_76), .Y(n_116) );
NAND2xp5_ASAP7_75t_L g117 ( .A(n_77), .B(n_1), .Y(n_117) );
INVx2_ASAP7_75t_L g118 ( .A(n_90), .Y(n_118) );
INVx1_ASAP7_75t_L g119 ( .A(n_76), .Y(n_119) );
INVx1_ASAP7_75t_L g120 ( .A(n_79), .Y(n_120) );
HB1xp67_ASAP7_75t_L g121 ( .A(n_77), .Y(n_121) );
INVx3_ASAP7_75t_L g122 ( .A(n_93), .Y(n_122) );
INVx2_ASAP7_75t_L g123 ( .A(n_90), .Y(n_123) );
BUFx6f_ASAP7_75t_L g124 ( .A(n_93), .Y(n_124) );
INVx1_ASAP7_75t_L g125 ( .A(n_79), .Y(n_125) );
OA21x2_ASAP7_75t_L g126 ( .A1(n_83), .A2(n_34), .B(n_72), .Y(n_126) );
NAND2xp5_ASAP7_75t_L g127 ( .A(n_82), .B(n_2), .Y(n_127) );
OA21x2_ASAP7_75t_L g128 ( .A1(n_83), .A2(n_32), .B(n_69), .Y(n_128) );
INVx1_ASAP7_75t_L g129 ( .A(n_85), .Y(n_129) );
INVx1_ASAP7_75t_L g130 ( .A(n_85), .Y(n_130) );
BUFx6f_ASAP7_75t_L g131 ( .A(n_93), .Y(n_131) );
NAND2xp5_ASAP7_75t_L g132 ( .A(n_116), .B(n_100), .Y(n_132) );
INVx1_ASAP7_75t_L g133 ( .A(n_109), .Y(n_133) );
BUFx3_ASAP7_75t_L g134 ( .A(n_114), .Y(n_134) );
BUFx3_ASAP7_75t_L g135 ( .A(n_114), .Y(n_135) );
AND2x2_ASAP7_75t_L g136 ( .A(n_121), .B(n_97), .Y(n_136) );
NOR2xp33_ASAP7_75t_L g137 ( .A(n_116), .B(n_102), .Y(n_137) );
NOR2xp33_ASAP7_75t_L g138 ( .A(n_119), .B(n_95), .Y(n_138) );
BUFx6f_ASAP7_75t_L g139 ( .A(n_124), .Y(n_139) );
BUFx3_ASAP7_75t_L g140 ( .A(n_114), .Y(n_140) );
NAND2xp5_ASAP7_75t_L g141 ( .A(n_119), .B(n_100), .Y(n_141) );
BUFx6f_ASAP7_75t_L g142 ( .A(n_124), .Y(n_142) );
BUFx10_ASAP7_75t_L g143 ( .A(n_110), .Y(n_143) );
INVx3_ASAP7_75t_L g144 ( .A(n_110), .Y(n_144) );
AOI22xp5_ASAP7_75t_L g145 ( .A1(n_110), .A2(n_75), .B1(n_82), .B2(n_106), .Y(n_145) );
INVx1_ASAP7_75t_L g146 ( .A(n_109), .Y(n_146) );
INVx1_ASAP7_75t_L g147 ( .A(n_109), .Y(n_147) );
INVx4_ASAP7_75t_L g148 ( .A(n_110), .Y(n_148) );
NAND2xp5_ASAP7_75t_L g149 ( .A(n_120), .B(n_101), .Y(n_149) );
BUFx6f_ASAP7_75t_L g150 ( .A(n_124), .Y(n_150) );
NAND2xp5_ASAP7_75t_L g151 ( .A(n_120), .B(n_101), .Y(n_151) );
AND2x2_ASAP7_75t_L g152 ( .A(n_125), .B(n_84), .Y(n_152) );
INVx1_ASAP7_75t_L g153 ( .A(n_112), .Y(n_153) );
NAND3xp33_ASAP7_75t_L g154 ( .A(n_125), .B(n_94), .C(n_107), .Y(n_154) );
INVx1_ASAP7_75t_L g155 ( .A(n_112), .Y(n_155) );
NOR2xp33_ASAP7_75t_L g156 ( .A(n_129), .B(n_94), .Y(n_156) );
INVx2_ASAP7_75t_L g157 ( .A(n_124), .Y(n_157) );
AND2x2_ASAP7_75t_L g158 ( .A(n_136), .B(n_113), .Y(n_158) );
INVx1_ASAP7_75t_L g159 ( .A(n_133), .Y(n_159) );
INVx2_ASAP7_75t_L g160 ( .A(n_134), .Y(n_160) );
O2A1O1Ixp33_ASAP7_75t_L g161 ( .A1(n_132), .A2(n_113), .B(n_117), .C(n_127), .Y(n_161) );
INVx5_ASAP7_75t_L g162 ( .A(n_143), .Y(n_162) );
INVx1_ASAP7_75t_L g163 ( .A(n_133), .Y(n_163) );
NAND2xp5_ASAP7_75t_L g164 ( .A(n_138), .B(n_129), .Y(n_164) );
INVx3_ASAP7_75t_L g165 ( .A(n_148), .Y(n_165) );
NAND2xp5_ASAP7_75t_L g166 ( .A(n_137), .B(n_130), .Y(n_166) );
NAND2xp5_ASAP7_75t_L g167 ( .A(n_136), .B(n_130), .Y(n_167) );
BUFx3_ASAP7_75t_L g168 ( .A(n_134), .Y(n_168) );
INVx1_ASAP7_75t_L g169 ( .A(n_146), .Y(n_169) );
NAND2xp5_ASAP7_75t_L g170 ( .A(n_136), .B(n_117), .Y(n_170) );
INVx1_ASAP7_75t_L g171 ( .A(n_146), .Y(n_171) );
INVx2_ASAP7_75t_L g172 ( .A(n_134), .Y(n_172) );
AOI22xp5_ASAP7_75t_L g173 ( .A1(n_145), .A2(n_127), .B1(n_115), .B2(n_84), .Y(n_173) );
BUFx2_ASAP7_75t_L g174 ( .A(n_148), .Y(n_174) );
NAND2xp5_ASAP7_75t_L g175 ( .A(n_152), .B(n_114), .Y(n_175) );
INVx1_ASAP7_75t_L g176 ( .A(n_147), .Y(n_176) );
BUFx6f_ASAP7_75t_L g177 ( .A(n_135), .Y(n_177) );
NAND2xp5_ASAP7_75t_L g178 ( .A(n_152), .B(n_115), .Y(n_178) );
INVx2_ASAP7_75t_L g179 ( .A(n_135), .Y(n_179) );
NAND2xp5_ASAP7_75t_L g180 ( .A(n_152), .B(n_88), .Y(n_180) );
INVx1_ASAP7_75t_L g181 ( .A(n_147), .Y(n_181) );
INVxp67_ASAP7_75t_L g182 ( .A(n_132), .Y(n_182) );
OR2x6_ASAP7_75t_L g183 ( .A(n_148), .B(n_91), .Y(n_183) );
INVx1_ASAP7_75t_L g184 ( .A(n_153), .Y(n_184) );
INVx3_ASAP7_75t_L g185 ( .A(n_148), .Y(n_185) );
OR2x6_ASAP7_75t_L g186 ( .A(n_144), .B(n_91), .Y(n_186) );
INVx3_ASAP7_75t_L g187 ( .A(n_143), .Y(n_187) );
INVx2_ASAP7_75t_L g188 ( .A(n_135), .Y(n_188) );
INVx1_ASAP7_75t_L g189 ( .A(n_153), .Y(n_189) );
CKINVDCx20_ASAP7_75t_R g190 ( .A(n_145), .Y(n_190) );
BUFx3_ASAP7_75t_L g191 ( .A(n_140), .Y(n_191) );
AOI22xp33_ASAP7_75t_L g192 ( .A1(n_158), .A2(n_144), .B1(n_154), .B2(n_156), .Y(n_192) );
AND2x6_ASAP7_75t_L g193 ( .A(n_187), .B(n_144), .Y(n_193) );
O2A1O1Ixp33_ASAP7_75t_L g194 ( .A1(n_170), .A2(n_149), .B(n_141), .C(n_151), .Y(n_194) );
INVx1_ASAP7_75t_L g195 ( .A(n_182), .Y(n_195) );
INVx1_ASAP7_75t_L g196 ( .A(n_175), .Y(n_196) );
NOR2xp33_ASAP7_75t_L g197 ( .A(n_158), .B(n_144), .Y(n_197) );
CKINVDCx20_ASAP7_75t_R g198 ( .A(n_190), .Y(n_198) );
INVx4_ASAP7_75t_L g199 ( .A(n_162), .Y(n_199) );
BUFx2_ASAP7_75t_L g200 ( .A(n_183), .Y(n_200) );
BUFx2_ASAP7_75t_L g201 ( .A(n_183), .Y(n_201) );
AND2x4_ASAP7_75t_L g202 ( .A(n_162), .B(n_111), .Y(n_202) );
OR2x6_ASAP7_75t_L g203 ( .A(n_183), .B(n_141), .Y(n_203) );
AOI22xp33_ASAP7_75t_L g204 ( .A1(n_183), .A2(n_154), .B1(n_155), .B2(n_143), .Y(n_204) );
INVx3_ASAP7_75t_L g205 ( .A(n_162), .Y(n_205) );
AOI21xp5_ASAP7_75t_L g206 ( .A1(n_161), .A2(n_140), .B(n_149), .Y(n_206) );
INVx4_ASAP7_75t_L g207 ( .A(n_162), .Y(n_207) );
INVx5_ASAP7_75t_L g208 ( .A(n_183), .Y(n_208) );
NOR2xp33_ASAP7_75t_L g209 ( .A(n_167), .B(n_143), .Y(n_209) );
AOI221xp5_ASAP7_75t_L g210 ( .A1(n_173), .A2(n_111), .B1(n_151), .B2(n_106), .C(n_104), .Y(n_210) );
INVx1_ASAP7_75t_L g211 ( .A(n_178), .Y(n_211) );
AOI21xp33_ASAP7_75t_L g212 ( .A1(n_186), .A2(n_140), .B(n_92), .Y(n_212) );
INVx1_ASAP7_75t_L g213 ( .A(n_159), .Y(n_213) );
INVx1_ASAP7_75t_L g214 ( .A(n_159), .Y(n_214) );
INVx2_ASAP7_75t_L g215 ( .A(n_163), .Y(n_215) );
AOI22xp33_ASAP7_75t_L g216 ( .A1(n_186), .A2(n_155), .B1(n_112), .B2(n_118), .Y(n_216) );
INVx2_ASAP7_75t_L g217 ( .A(n_163), .Y(n_217) );
OAI22xp5_ASAP7_75t_L g218 ( .A1(n_186), .A2(n_173), .B1(n_166), .B2(n_164), .Y(n_218) );
NOR2xp33_ASAP7_75t_L g219 ( .A(n_180), .B(n_104), .Y(n_219) );
NAND2xp5_ASAP7_75t_L g220 ( .A(n_186), .B(n_123), .Y(n_220) );
BUFx12f_ASAP7_75t_L g221 ( .A(n_186), .Y(n_221) );
INVx1_ASAP7_75t_SL g222 ( .A(n_174), .Y(n_222) );
AOI22xp33_ASAP7_75t_L g223 ( .A1(n_169), .A2(n_118), .B1(n_123), .B2(n_93), .Y(n_223) );
NOR2x1_ASAP7_75t_L g224 ( .A(n_169), .B(n_99), .Y(n_224) );
AND2x2_ASAP7_75t_L g225 ( .A(n_211), .B(n_171), .Y(n_225) );
INVx2_ASAP7_75t_L g226 ( .A(n_215), .Y(n_226) );
AND2x2_ASAP7_75t_L g227 ( .A(n_195), .B(n_171), .Y(n_227) );
INVx1_ASAP7_75t_L g228 ( .A(n_215), .Y(n_228) );
AOI22xp33_ASAP7_75t_SL g229 ( .A1(n_221), .A2(n_174), .B1(n_189), .B2(n_176), .Y(n_229) );
INVx2_ASAP7_75t_L g230 ( .A(n_217), .Y(n_230) );
INVxp33_ASAP7_75t_SL g231 ( .A(n_218), .Y(n_231) );
INVx1_ASAP7_75t_L g232 ( .A(n_217), .Y(n_232) );
AOI22xp33_ASAP7_75t_L g233 ( .A1(n_221), .A2(n_185), .B1(n_165), .B2(n_189), .Y(n_233) );
INVx2_ASAP7_75t_L g234 ( .A(n_213), .Y(n_234) );
INVx1_ASAP7_75t_L g235 ( .A(n_214), .Y(n_235) );
AOI22xp33_ASAP7_75t_L g236 ( .A1(n_200), .A2(n_185), .B1(n_165), .B2(n_176), .Y(n_236) );
OAI22xp33_ASAP7_75t_L g237 ( .A1(n_208), .A2(n_184), .B1(n_181), .B2(n_162), .Y(n_237) );
CKINVDCx5p33_ASAP7_75t_R g238 ( .A(n_198), .Y(n_238) );
AOI22xp33_ASAP7_75t_L g239 ( .A1(n_201), .A2(n_165), .B1(n_185), .B2(n_181), .Y(n_239) );
AOI22xp33_ASAP7_75t_L g240 ( .A1(n_209), .A2(n_165), .B1(n_185), .B2(n_184), .Y(n_240) );
BUFx5_ASAP7_75t_L g241 ( .A(n_193), .Y(n_241) );
NAND2xp5_ASAP7_75t_L g242 ( .A(n_197), .B(n_162), .Y(n_242) );
AOI222xp33_ASAP7_75t_L g243 ( .A1(n_210), .A2(n_123), .B1(n_118), .B2(n_93), .C1(n_89), .C2(n_98), .Y(n_243) );
AND2x4_ASAP7_75t_L g244 ( .A(n_208), .B(n_187), .Y(n_244) );
INVx1_ASAP7_75t_L g245 ( .A(n_196), .Y(n_245) );
INVx1_ASAP7_75t_L g246 ( .A(n_194), .Y(n_246) );
INVx8_ASAP7_75t_L g247 ( .A(n_208), .Y(n_247) );
AO221x2_ASAP7_75t_L g248 ( .A1(n_220), .A2(n_86), .B1(n_87), .B2(n_89), .C(n_98), .Y(n_248) );
BUFx3_ASAP7_75t_L g249 ( .A(n_208), .Y(n_249) );
OAI22xp5_ASAP7_75t_L g250 ( .A1(n_231), .A2(n_203), .B1(n_216), .B2(n_222), .Y(n_250) );
OAI22xp5_ASAP7_75t_L g251 ( .A1(n_229), .A2(n_203), .B1(n_216), .B2(n_204), .Y(n_251) );
BUFx4f_ASAP7_75t_L g252 ( .A(n_247), .Y(n_252) );
INVx1_ASAP7_75t_L g253 ( .A(n_227), .Y(n_253) );
AOI222xp33_ASAP7_75t_L g254 ( .A1(n_245), .A2(n_197), .B1(n_219), .B2(n_198), .C1(n_192), .C2(n_202), .Y(n_254) );
OAI22xp5_ASAP7_75t_L g255 ( .A1(n_228), .A2(n_203), .B1(n_204), .B2(n_209), .Y(n_255) );
OAI22xp5_ASAP7_75t_L g256 ( .A1(n_228), .A2(n_192), .B1(n_202), .B2(n_219), .Y(n_256) );
AOI22xp33_ASAP7_75t_L g257 ( .A1(n_248), .A2(n_224), .B1(n_202), .B2(n_206), .Y(n_257) );
AOI21xp33_ASAP7_75t_L g258 ( .A1(n_246), .A2(n_212), .B(n_205), .Y(n_258) );
AOI22xp33_ASAP7_75t_L g259 ( .A1(n_248), .A2(n_223), .B1(n_93), .B2(n_207), .Y(n_259) );
AOI22xp33_ASAP7_75t_L g260 ( .A1(n_248), .A2(n_223), .B1(n_207), .B2(n_199), .Y(n_260) );
AND2x2_ASAP7_75t_L g261 ( .A(n_227), .B(n_199), .Y(n_261) );
NAND4xp25_ASAP7_75t_L g262 ( .A(n_243), .B(n_86), .C(n_87), .D(n_103), .Y(n_262) );
OAI211xp5_ASAP7_75t_L g263 ( .A1(n_245), .A2(n_103), .B(n_105), .C(n_107), .Y(n_263) );
INVx1_ASAP7_75t_L g264 ( .A(n_225), .Y(n_264) );
OAI22xp5_ASAP7_75t_L g265 ( .A1(n_232), .A2(n_205), .B1(n_168), .B2(n_191), .Y(n_265) );
OAI221xp5_ASAP7_75t_L g266 ( .A1(n_246), .A2(n_105), .B1(n_187), .B2(n_188), .C(n_179), .Y(n_266) );
NOR2xp33_ASAP7_75t_L g267 ( .A(n_238), .B(n_187), .Y(n_267) );
AOI222xp33_ASAP7_75t_L g268 ( .A1(n_225), .A2(n_193), .B1(n_172), .B2(n_188), .C1(n_179), .C2(n_160), .Y(n_268) );
INVx2_ASAP7_75t_L g269 ( .A(n_226), .Y(n_269) );
AOI22xp33_ASAP7_75t_L g270 ( .A1(n_248), .A2(n_193), .B1(n_128), .B2(n_126), .Y(n_270) );
OA21x2_ASAP7_75t_L g271 ( .A1(n_270), .A2(n_232), .B(n_234), .Y(n_271) );
AOI22xp33_ASAP7_75t_L g272 ( .A1(n_254), .A2(n_242), .B1(n_235), .B2(n_234), .Y(n_272) );
AOI22xp33_ASAP7_75t_L g273 ( .A1(n_251), .A2(n_235), .B1(n_234), .B2(n_247), .Y(n_273) );
INVx2_ASAP7_75t_L g274 ( .A(n_269), .Y(n_274) );
BUFx2_ASAP7_75t_L g275 ( .A(n_261), .Y(n_275) );
OAI221xp5_ASAP7_75t_L g276 ( .A1(n_259), .A2(n_240), .B1(n_239), .B2(n_236), .C(n_233), .Y(n_276) );
OAI33xp33_ASAP7_75t_L g277 ( .A1(n_262), .A2(n_237), .A3(n_226), .B1(n_230), .B2(n_108), .B3(n_6), .Y(n_277) );
NAND3xp33_ASAP7_75t_L g278 ( .A(n_257), .B(n_230), .C(n_124), .Y(n_278) );
NAND2xp5_ASAP7_75t_L g279 ( .A(n_264), .B(n_249), .Y(n_279) );
NAND2xp5_ASAP7_75t_L g280 ( .A(n_253), .B(n_249), .Y(n_280) );
AOI22xp33_ASAP7_75t_L g281 ( .A1(n_259), .A2(n_247), .B1(n_249), .B2(n_244), .Y(n_281) );
AOI222xp33_ASAP7_75t_L g282 ( .A1(n_252), .A2(n_247), .B1(n_244), .B2(n_193), .C1(n_122), .C2(n_172), .Y(n_282) );
OAI22xp5_ASAP7_75t_L g283 ( .A1(n_250), .A2(n_247), .B1(n_244), .B2(n_126), .Y(n_283) );
AOI22xp33_ASAP7_75t_L g284 ( .A1(n_252), .A2(n_244), .B1(n_241), .B2(n_193), .Y(n_284) );
INVx1_ASAP7_75t_L g285 ( .A(n_256), .Y(n_285) );
AND2x2_ASAP7_75t_L g286 ( .A(n_260), .B(n_128), .Y(n_286) );
AND2x2_ASAP7_75t_L g287 ( .A(n_260), .B(n_128), .Y(n_287) );
AOI22xp33_ASAP7_75t_L g288 ( .A1(n_255), .A2(n_241), .B1(n_177), .B2(n_191), .Y(n_288) );
AND2x2_ASAP7_75t_L g289 ( .A(n_257), .B(n_128), .Y(n_289) );
INVx1_ASAP7_75t_L g290 ( .A(n_270), .Y(n_290) );
OA21x2_ASAP7_75t_L g291 ( .A1(n_258), .A2(n_157), .B(n_172), .Y(n_291) );
AND2x4_ASAP7_75t_L g292 ( .A(n_267), .B(n_160), .Y(n_292) );
NAND2xp33_ASAP7_75t_SL g293 ( .A(n_275), .B(n_265), .Y(n_293) );
INVx1_ASAP7_75t_L g294 ( .A(n_271), .Y(n_294) );
OAI22xp5_ASAP7_75t_L g295 ( .A1(n_281), .A2(n_263), .B1(n_266), .B2(n_268), .Y(n_295) );
AND2x2_ASAP7_75t_L g296 ( .A(n_290), .B(n_126), .Y(n_296) );
AND2x4_ASAP7_75t_L g297 ( .A(n_290), .B(n_46), .Y(n_297) );
AOI22xp33_ASAP7_75t_L g298 ( .A1(n_273), .A2(n_241), .B1(n_128), .B2(n_126), .Y(n_298) );
OAI33xp33_ASAP7_75t_L g299 ( .A1(n_283), .A2(n_2), .A3(n_3), .B1(n_4), .B2(n_5), .B3(n_7), .Y(n_299) );
INVx1_ASAP7_75t_L g300 ( .A(n_271), .Y(n_300) );
INVx2_ASAP7_75t_SL g301 ( .A(n_275), .Y(n_301) );
INVx1_ASAP7_75t_L g302 ( .A(n_271), .Y(n_302) );
INVx1_ASAP7_75t_L g303 ( .A(n_271), .Y(n_303) );
AND2x2_ASAP7_75t_L g304 ( .A(n_285), .B(n_126), .Y(n_304) );
OAI22xp5_ASAP7_75t_L g305 ( .A1(n_272), .A2(n_241), .B1(n_191), .B2(n_168), .Y(n_305) );
AND2x4_ASAP7_75t_L g306 ( .A(n_285), .B(n_42), .Y(n_306) );
INVx2_ASAP7_75t_L g307 ( .A(n_274), .Y(n_307) );
NAND2xp5_ASAP7_75t_L g308 ( .A(n_279), .B(n_3), .Y(n_308) );
INVx1_ASAP7_75t_L g309 ( .A(n_271), .Y(n_309) );
INVx1_ASAP7_75t_L g310 ( .A(n_274), .Y(n_310) );
AND2x2_ASAP7_75t_L g311 ( .A(n_274), .B(n_4), .Y(n_311) );
NAND2xp5_ASAP7_75t_L g312 ( .A(n_279), .B(n_5), .Y(n_312) );
AND2x2_ASAP7_75t_L g313 ( .A(n_289), .B(n_7), .Y(n_313) );
HB1xp67_ASAP7_75t_L g314 ( .A(n_280), .Y(n_314) );
OAI33xp33_ASAP7_75t_L g315 ( .A1(n_283), .A2(n_280), .A3(n_278), .B1(n_277), .B2(n_11), .B3(n_12), .Y(n_315) );
BUFx3_ASAP7_75t_L g316 ( .A(n_292), .Y(n_316) );
OR2x2_ASAP7_75t_L g317 ( .A(n_278), .B(n_8), .Y(n_317) );
INVx2_ASAP7_75t_L g318 ( .A(n_291), .Y(n_318) );
NAND3xp33_ASAP7_75t_L g319 ( .A(n_282), .B(n_124), .C(n_131), .Y(n_319) );
AND2x4_ASAP7_75t_SL g320 ( .A(n_284), .B(n_241), .Y(n_320) );
AOI21xp5_ASAP7_75t_SL g321 ( .A1(n_286), .A2(n_241), .B(n_168), .Y(n_321) );
AND2x2_ASAP7_75t_L g322 ( .A(n_289), .B(n_8), .Y(n_322) );
HB1xp67_ASAP7_75t_L g323 ( .A(n_292), .Y(n_323) );
INVx1_ASAP7_75t_L g324 ( .A(n_310), .Y(n_324) );
HB1xp67_ASAP7_75t_L g325 ( .A(n_301), .Y(n_325) );
NAND2xp5_ASAP7_75t_L g326 ( .A(n_314), .B(n_287), .Y(n_326) );
AND2x2_ASAP7_75t_L g327 ( .A(n_310), .B(n_287), .Y(n_327) );
AND2x2_ASAP7_75t_L g328 ( .A(n_307), .B(n_286), .Y(n_328) );
OR2x6_ASAP7_75t_L g329 ( .A(n_321), .B(n_291), .Y(n_329) );
HB1xp67_ASAP7_75t_L g330 ( .A(n_301), .Y(n_330) );
BUFx3_ASAP7_75t_L g331 ( .A(n_316), .Y(n_331) );
AND2x2_ASAP7_75t_L g332 ( .A(n_307), .B(n_291), .Y(n_332) );
AOI22xp33_ASAP7_75t_L g333 ( .A1(n_295), .A2(n_277), .B1(n_276), .B2(n_292), .Y(n_333) );
AND2x2_ASAP7_75t_L g334 ( .A(n_294), .B(n_291), .Y(n_334) );
AOI21xp33_ASAP7_75t_SL g335 ( .A1(n_319), .A2(n_317), .B(n_282), .Y(n_335) );
INVx1_ASAP7_75t_L g336 ( .A(n_294), .Y(n_336) );
AND2x2_ASAP7_75t_L g337 ( .A(n_300), .B(n_291), .Y(n_337) );
AOI21xp5_ASAP7_75t_L g338 ( .A1(n_321), .A2(n_288), .B(n_276), .Y(n_338) );
NAND2xp5_ASAP7_75t_L g339 ( .A(n_313), .B(n_292), .Y(n_339) );
AND2x2_ASAP7_75t_L g340 ( .A(n_300), .B(n_124), .Y(n_340) );
HB1xp67_ASAP7_75t_L g341 ( .A(n_311), .Y(n_341) );
INVx1_ASAP7_75t_L g342 ( .A(n_302), .Y(n_342) );
NAND2xp5_ASAP7_75t_L g343 ( .A(n_313), .B(n_122), .Y(n_343) );
AOI221x1_ASAP7_75t_L g344 ( .A1(n_319), .A2(n_131), .B1(n_122), .B2(n_12), .C(n_13), .Y(n_344) );
INVx3_ASAP7_75t_L g345 ( .A(n_318), .Y(n_345) );
OAI21xp5_ASAP7_75t_L g346 ( .A1(n_317), .A2(n_122), .B(n_157), .Y(n_346) );
OAI211xp5_ASAP7_75t_L g347 ( .A1(n_293), .A2(n_131), .B(n_10), .C(n_14), .Y(n_347) );
INVx1_ASAP7_75t_L g348 ( .A(n_302), .Y(n_348) );
AND2x2_ASAP7_75t_L g349 ( .A(n_303), .B(n_131), .Y(n_349) );
INVx2_ASAP7_75t_L g350 ( .A(n_303), .Y(n_350) );
INVx1_ASAP7_75t_L g351 ( .A(n_309), .Y(n_351) );
INVx1_ASAP7_75t_L g352 ( .A(n_309), .Y(n_352) );
NOR3xp33_ASAP7_75t_L g353 ( .A(n_299), .B(n_157), .C(n_14), .Y(n_353) );
INVx1_ASAP7_75t_L g354 ( .A(n_318), .Y(n_354) );
AND2x2_ASAP7_75t_L g355 ( .A(n_322), .B(n_131), .Y(n_355) );
AND2x2_ASAP7_75t_L g356 ( .A(n_322), .B(n_131), .Y(n_356) );
NAND2xp5_ASAP7_75t_L g357 ( .A(n_323), .B(n_131), .Y(n_357) );
OR2x2_ASAP7_75t_L g358 ( .A(n_316), .B(n_9), .Y(n_358) );
INVx1_ASAP7_75t_SL g359 ( .A(n_316), .Y(n_359) );
INVx2_ASAP7_75t_L g360 ( .A(n_296), .Y(n_360) );
INVx1_ASAP7_75t_L g361 ( .A(n_311), .Y(n_361) );
AOI33xp33_ASAP7_75t_L g362 ( .A1(n_306), .A2(n_16), .A3(n_18), .B1(n_19), .B2(n_21), .B3(n_22), .Y(n_362) );
NOR2xp33_ASAP7_75t_L g363 ( .A(n_308), .B(n_16), .Y(n_363) );
NAND2xp5_ASAP7_75t_SL g364 ( .A(n_306), .B(n_241), .Y(n_364) );
AND2x2_ASAP7_75t_L g365 ( .A(n_297), .B(n_23), .Y(n_365) );
AND2x2_ASAP7_75t_L g366 ( .A(n_297), .B(n_25), .Y(n_366) );
NAND2xp5_ASAP7_75t_L g367 ( .A(n_296), .B(n_241), .Y(n_367) );
AND2x2_ASAP7_75t_L g368 ( .A(n_297), .B(n_306), .Y(n_368) );
AND2x2_ASAP7_75t_L g369 ( .A(n_297), .B(n_27), .Y(n_369) );
HB1xp67_ASAP7_75t_L g370 ( .A(n_325), .Y(n_370) );
OAI21xp33_ASAP7_75t_L g371 ( .A1(n_333), .A2(n_306), .B(n_312), .Y(n_371) );
NAND2xp5_ASAP7_75t_L g372 ( .A(n_336), .B(n_304), .Y(n_372) );
AND2x2_ASAP7_75t_L g373 ( .A(n_330), .B(n_320), .Y(n_373) );
HB1xp67_ASAP7_75t_L g374 ( .A(n_355), .Y(n_374) );
AND2x2_ASAP7_75t_L g375 ( .A(n_339), .B(n_320), .Y(n_375) );
AND2x2_ASAP7_75t_L g376 ( .A(n_339), .B(n_304), .Y(n_376) );
NAND2xp5_ASAP7_75t_L g377 ( .A(n_336), .B(n_315), .Y(n_377) );
O2A1O1Ixp33_ASAP7_75t_L g378 ( .A1(n_335), .A2(n_305), .B(n_298), .C(n_241), .Y(n_378) );
INVx1_ASAP7_75t_SL g379 ( .A(n_359), .Y(n_379) );
NAND2xp5_ASAP7_75t_L g380 ( .A(n_342), .B(n_31), .Y(n_380) );
AND2x4_ASAP7_75t_L g381 ( .A(n_331), .B(n_37), .Y(n_381) );
OR2x6_ASAP7_75t_L g382 ( .A(n_368), .B(n_38), .Y(n_382) );
AND4x1_ASAP7_75t_L g383 ( .A(n_362), .B(n_40), .C(n_41), .D(n_44), .Y(n_383) );
INVx1_ASAP7_75t_L g384 ( .A(n_324), .Y(n_384) );
NAND3xp33_ASAP7_75t_L g385 ( .A(n_363), .B(n_150), .C(n_142), .Y(n_385) );
NOR2x1_ASAP7_75t_L g386 ( .A(n_347), .B(n_48), .Y(n_386) );
AOI211xp5_ASAP7_75t_SL g387 ( .A1(n_347), .A2(n_49), .B(n_50), .C(n_52), .Y(n_387) );
INVx1_ASAP7_75t_SL g388 ( .A(n_359), .Y(n_388) );
INVx1_ASAP7_75t_L g389 ( .A(n_342), .Y(n_389) );
OR2x2_ASAP7_75t_L g390 ( .A(n_341), .B(n_54), .Y(n_390) );
NAND2xp5_ASAP7_75t_L g391 ( .A(n_348), .B(n_59), .Y(n_391) );
OR2x2_ASAP7_75t_L g392 ( .A(n_326), .B(n_60), .Y(n_392) );
NAND2xp5_ASAP7_75t_L g393 ( .A(n_348), .B(n_62), .Y(n_393) );
AND2x2_ASAP7_75t_L g394 ( .A(n_368), .B(n_63), .Y(n_394) );
INVx1_ASAP7_75t_L g395 ( .A(n_351), .Y(n_395) );
INVx1_ASAP7_75t_L g396 ( .A(n_351), .Y(n_396) );
NAND2xp5_ASAP7_75t_L g397 ( .A(n_352), .B(n_64), .Y(n_397) );
INVxp67_ASAP7_75t_L g398 ( .A(n_352), .Y(n_398) );
AND2x4_ASAP7_75t_SL g399 ( .A(n_365), .B(n_177), .Y(n_399) );
AND2x2_ASAP7_75t_L g400 ( .A(n_331), .B(n_65), .Y(n_400) );
INVx2_ASAP7_75t_L g401 ( .A(n_345), .Y(n_401) );
INVx3_ASAP7_75t_L g402 ( .A(n_331), .Y(n_402) );
AND2x4_ASAP7_75t_L g403 ( .A(n_350), .B(n_68), .Y(n_403) );
CKINVDCx16_ASAP7_75t_R g404 ( .A(n_365), .Y(n_404) );
OR2x2_ASAP7_75t_L g405 ( .A(n_326), .B(n_74), .Y(n_405) );
INVx1_ASAP7_75t_L g406 ( .A(n_358), .Y(n_406) );
INVx1_ASAP7_75t_L g407 ( .A(n_358), .Y(n_407) );
OAI21xp5_ASAP7_75t_L g408 ( .A1(n_344), .A2(n_177), .B(n_142), .Y(n_408) );
NOR3xp33_ASAP7_75t_L g409 ( .A(n_343), .B(n_139), .C(n_142), .Y(n_409) );
INVx2_ASAP7_75t_L g410 ( .A(n_345), .Y(n_410) );
OR2x2_ASAP7_75t_L g411 ( .A(n_361), .B(n_177), .Y(n_411) );
INVx1_ASAP7_75t_L g412 ( .A(n_340), .Y(n_412) );
INVx1_ASAP7_75t_L g413 ( .A(n_340), .Y(n_413) );
A2O1A1Ixp33_ASAP7_75t_L g414 ( .A1(n_335), .A2(n_177), .B(n_142), .C(n_150), .Y(n_414) );
NOR2xp67_ASAP7_75t_L g415 ( .A(n_345), .B(n_139), .Y(n_415) );
INVxp67_ASAP7_75t_L g416 ( .A(n_370), .Y(n_416) );
INVx1_ASAP7_75t_SL g417 ( .A(n_379), .Y(n_417) );
INVx1_ASAP7_75t_L g418 ( .A(n_389), .Y(n_418) );
OR2x2_ASAP7_75t_L g419 ( .A(n_374), .B(n_360), .Y(n_419) );
AND2x2_ASAP7_75t_L g420 ( .A(n_376), .B(n_360), .Y(n_420) );
OAI21x1_ASAP7_75t_L g421 ( .A1(n_377), .A2(n_334), .B(n_337), .Y(n_421) );
INVxp67_ASAP7_75t_L g422 ( .A(n_377), .Y(n_422) );
INVx1_ASAP7_75t_L g423 ( .A(n_395), .Y(n_423) );
XNOR2xp5_ASAP7_75t_L g424 ( .A(n_375), .B(n_356), .Y(n_424) );
INVx1_ASAP7_75t_L g425 ( .A(n_396), .Y(n_425) );
NAND2xp5_ASAP7_75t_L g426 ( .A(n_406), .B(n_327), .Y(n_426) );
AND2x2_ASAP7_75t_SL g427 ( .A(n_404), .B(n_369), .Y(n_427) );
NOR2xp33_ASAP7_75t_L g428 ( .A(n_371), .B(n_343), .Y(n_428) );
INVx1_ASAP7_75t_SL g429 ( .A(n_388), .Y(n_429) );
INVx1_ASAP7_75t_L g430 ( .A(n_398), .Y(n_430) );
AOI21xp5_ASAP7_75t_SL g431 ( .A1(n_382), .A2(n_364), .B(n_369), .Y(n_431) );
INVx1_ASAP7_75t_L g432 ( .A(n_398), .Y(n_432) );
NAND2xp5_ASAP7_75t_SL g433 ( .A(n_415), .B(n_354), .Y(n_433) );
INVx3_ASAP7_75t_L g434 ( .A(n_402), .Y(n_434) );
INVx1_ASAP7_75t_L g435 ( .A(n_384), .Y(n_435) );
NAND2xp5_ASAP7_75t_L g436 ( .A(n_407), .B(n_372), .Y(n_436) );
AND2x2_ASAP7_75t_L g437 ( .A(n_401), .B(n_327), .Y(n_437) );
INVx1_ASAP7_75t_SL g438 ( .A(n_399), .Y(n_438) );
INVx2_ASAP7_75t_L g439 ( .A(n_410), .Y(n_439) );
AOI22xp33_ASAP7_75t_SL g440 ( .A1(n_382), .A2(n_366), .B1(n_355), .B2(n_356), .Y(n_440) );
INVxp67_ASAP7_75t_SL g441 ( .A(n_409), .Y(n_441) );
OR2x2_ASAP7_75t_L g442 ( .A(n_372), .B(n_354), .Y(n_442) );
INVx1_ASAP7_75t_L g443 ( .A(n_412), .Y(n_443) );
OR2x2_ASAP7_75t_L g444 ( .A(n_413), .B(n_328), .Y(n_444) );
NOR2xp33_ASAP7_75t_L g445 ( .A(n_402), .B(n_357), .Y(n_445) );
AOI21xp33_ASAP7_75t_SL g446 ( .A1(n_382), .A2(n_385), .B(n_390), .Y(n_446) );
INVx1_ASAP7_75t_L g447 ( .A(n_380), .Y(n_447) );
AOI221x1_ASAP7_75t_L g448 ( .A1(n_408), .A2(n_357), .B1(n_338), .B2(n_353), .C(n_346), .Y(n_448) );
AND2x2_ASAP7_75t_L g449 ( .A(n_373), .B(n_328), .Y(n_449) );
AOI22xp5_ASAP7_75t_L g450 ( .A1(n_394), .A2(n_338), .B1(n_366), .B2(n_346), .Y(n_450) );
OR2x2_ASAP7_75t_L g451 ( .A(n_411), .B(n_349), .Y(n_451) );
NOR2xp33_ASAP7_75t_L g452 ( .A(n_392), .B(n_349), .Y(n_452) );
AOI22x1_ASAP7_75t_L g453 ( .A1(n_387), .A2(n_344), .B1(n_337), .B2(n_334), .Y(n_453) );
OAI22xp5_ASAP7_75t_L g454 ( .A1(n_386), .A2(n_329), .B1(n_367), .B2(n_332), .Y(n_454) );
XNOR2x1_ASAP7_75t_L g455 ( .A(n_405), .B(n_329), .Y(n_455) );
BUFx2_ASAP7_75t_L g456 ( .A(n_381), .Y(n_456) );
INVx1_ASAP7_75t_L g457 ( .A(n_380), .Y(n_457) );
OAI211xp5_ASAP7_75t_SL g458 ( .A1(n_387), .A2(n_367), .B(n_329), .C(n_332), .Y(n_458) );
AOI322xp5_ASAP7_75t_L g459 ( .A1(n_381), .A2(n_139), .A3(n_142), .B1(n_150), .B2(n_177), .C1(n_329), .C2(n_400), .Y(n_459) );
AOI21xp5_ASAP7_75t_L g460 ( .A1(n_414), .A2(n_329), .B(n_142), .Y(n_460) );
NOR2xp33_ASAP7_75t_L g461 ( .A(n_383), .B(n_139), .Y(n_461) );
INVxp33_ASAP7_75t_L g462 ( .A(n_403), .Y(n_462) );
AOI21xp5_ASAP7_75t_L g463 ( .A1(n_408), .A2(n_150), .B(n_378), .Y(n_463) );
NOR2xp33_ASAP7_75t_L g464 ( .A(n_391), .B(n_150), .Y(n_464) );
INVx1_ASAP7_75t_L g465 ( .A(n_391), .Y(n_465) );
INVx1_ASAP7_75t_L g466 ( .A(n_393), .Y(n_466) );
AND2x2_ASAP7_75t_L g467 ( .A(n_403), .B(n_150), .Y(n_467) );
AND2x2_ASAP7_75t_L g468 ( .A(n_393), .B(n_397), .Y(n_468) );
OAI22xp33_ASAP7_75t_L g469 ( .A1(n_397), .A2(n_404), .B1(n_382), .B2(n_335), .Y(n_469) );
INVx1_ASAP7_75t_L g470 ( .A(n_378), .Y(n_470) );
INVx1_ASAP7_75t_L g471 ( .A(n_389), .Y(n_471) );
A2O1A1Ixp33_ASAP7_75t_L g472 ( .A1(n_371), .A2(n_335), .B(n_387), .C(n_386), .Y(n_472) );
INVx1_ASAP7_75t_L g473 ( .A(n_389), .Y(n_473) );
INVx1_ASAP7_75t_L g474 ( .A(n_389), .Y(n_474) );
INVx1_ASAP7_75t_L g475 ( .A(n_389), .Y(n_475) );
O2A1O1Ixp5_ASAP7_75t_L g476 ( .A1(n_387), .A2(n_377), .B(n_347), .C(n_402), .Y(n_476) );
NOR2xp33_ASAP7_75t_L g477 ( .A(n_370), .B(n_371), .Y(n_477) );
INVx1_ASAP7_75t_L g478 ( .A(n_430), .Y(n_478) );
AOI22xp33_ASAP7_75t_L g479 ( .A1(n_469), .A2(n_427), .B1(n_428), .B2(n_470), .Y(n_479) );
INVx1_ASAP7_75t_L g480 ( .A(n_432), .Y(n_480) );
XOR2x2_ASAP7_75t_L g481 ( .A(n_427), .B(n_455), .Y(n_481) );
INVx2_ASAP7_75t_L g482 ( .A(n_439), .Y(n_482) );
AOI22xp5_ASAP7_75t_L g483 ( .A1(n_469), .A2(n_477), .B1(n_422), .B2(n_428), .Y(n_483) );
OAI21xp5_ASAP7_75t_SL g484 ( .A1(n_472), .A2(n_440), .B(n_446), .Y(n_484) );
NOR2x1_ASAP7_75t_L g485 ( .A(n_431), .B(n_472), .Y(n_485) );
NAND5xp2_ASAP7_75t_L g486 ( .A(n_459), .B(n_450), .C(n_463), .D(n_477), .E(n_461), .Y(n_486) );
OAI21xp33_ASAP7_75t_L g487 ( .A1(n_421), .A2(n_436), .B(n_431), .Y(n_487) );
INVx1_ASAP7_75t_L g488 ( .A(n_421), .Y(n_488) );
AOI211xp5_ASAP7_75t_SL g489 ( .A1(n_454), .A2(n_441), .B(n_458), .C(n_460), .Y(n_489) );
AOI221xp5_ASAP7_75t_L g490 ( .A1(n_416), .A2(n_476), .B1(n_443), .B2(n_447), .C(n_457), .Y(n_490) );
AOI22xp5_ASAP7_75t_L g491 ( .A1(n_456), .A2(n_417), .B1(n_429), .B2(n_445), .Y(n_491) );
AOI221xp5_ASAP7_75t_SL g492 ( .A1(n_426), .A2(n_424), .B1(n_449), .B2(n_420), .C(n_445), .Y(n_492) );
OAI22xp5_ASAP7_75t_L g493 ( .A1(n_434), .A2(n_438), .B1(n_453), .B2(n_419), .Y(n_493) );
NAND4xp25_ASAP7_75t_SL g494 ( .A(n_485), .B(n_448), .C(n_449), .D(n_444), .Y(n_494) );
OAI21xp33_ASAP7_75t_L g495 ( .A1(n_484), .A2(n_479), .B(n_487), .Y(n_495) );
NOR2x1p5_ASAP7_75t_L g496 ( .A(n_484), .B(n_434), .Y(n_496) );
OAI21xp5_ASAP7_75t_SL g497 ( .A1(n_489), .A2(n_434), .B(n_462), .Y(n_497) );
AOI211xp5_ASAP7_75t_L g498 ( .A1(n_493), .A2(n_466), .B(n_465), .C(n_468), .Y(n_498) );
AND2x2_ASAP7_75t_L g499 ( .A(n_492), .B(n_420), .Y(n_499) );
OAI211xp5_ASAP7_75t_SL g500 ( .A1(n_490), .A2(n_433), .B(n_461), .C(n_475), .Y(n_500) );
AOI221xp5_ASAP7_75t_L g501 ( .A1(n_488), .A2(n_418), .B1(n_423), .B2(n_473), .C(n_425), .Y(n_501) );
NOR3x2_ASAP7_75t_L g502 ( .A(n_481), .B(n_442), .C(n_451), .Y(n_502) );
NOR3xp33_ASAP7_75t_L g503 ( .A(n_495), .B(n_486), .C(n_483), .Y(n_503) );
AND4x1_ASAP7_75t_L g504 ( .A(n_498), .B(n_491), .C(n_478), .D(n_480), .Y(n_504) );
NOR4xp25_ASAP7_75t_L g505 ( .A(n_494), .B(n_482), .C(n_464), .D(n_474), .Y(n_505) );
NAND4xp25_ASAP7_75t_L g506 ( .A(n_497), .B(n_452), .C(n_464), .D(n_433), .Y(n_506) );
AOI211x1_ASAP7_75t_L g507 ( .A1(n_499), .A2(n_471), .B(n_435), .C(n_437), .Y(n_507) );
INVx1_ASAP7_75t_L g508 ( .A(n_503), .Y(n_508) );
INVx1_ASAP7_75t_L g509 ( .A(n_506), .Y(n_509) );
INVx1_ASAP7_75t_L g510 ( .A(n_507), .Y(n_510) );
INVx1_ASAP7_75t_L g511 ( .A(n_508), .Y(n_511) );
OAI221xp5_ASAP7_75t_L g512 ( .A1(n_509), .A2(n_505), .B1(n_504), .B2(n_500), .C(n_502), .Y(n_512) );
INVx4_ASAP7_75t_L g513 ( .A(n_511), .Y(n_513) );
INVx1_ASAP7_75t_L g514 ( .A(n_513), .Y(n_514) );
AOI22x1_ASAP7_75t_L g515 ( .A1(n_514), .A2(n_496), .B1(n_510), .B2(n_512), .Y(n_515) );
AOI21xp5_ASAP7_75t_L g516 ( .A1(n_515), .A2(n_501), .B(n_467), .Y(n_516) );
endmodule