module real_jpeg_7142_n_25 (n_17, n_8, n_0, n_157, n_21, n_2, n_10, n_9, n_12, n_154, n_156, n_152, n_24, n_6, n_153, n_151, n_23, n_11, n_14, n_7, n_22, n_18, n_3, n_5, n_4, n_150, n_1, n_20, n_19, n_148, n_149, n_16, n_15, n_13, n_155, n_25);

input n_17;
input n_8;
input n_0;
input n_157;
input n_21;
input n_2;
input n_10;
input n_9;
input n_12;
input n_154;
input n_156;
input n_152;
input n_24;
input n_6;
input n_153;
input n_151;
input n_23;
input n_11;
input n_14;
input n_7;
input n_22;
input n_18;
input n_3;
input n_5;
input n_4;
input n_150;
input n_1;
input n_20;
input n_19;
input n_148;
input n_149;
input n_16;
input n_15;
input n_13;
input n_155;

output n_25;

wire n_108;
wire n_54;
wire n_37;
wire n_73;
wire n_35;
wire n_38;
wire n_29;
wire n_91;
wire n_49;
wire n_114;
wire n_68;
wire n_146;
wire n_83;
wire n_78;
wire n_104;
wire n_64;
wire n_47;
wire n_131;
wire n_87;
wire n_40;
wire n_105;
wire n_115;
wire n_98;
wire n_27;
wire n_56;
wire n_48;
wire n_140;
wire n_126;
wire n_120;
wire n_113;
wire n_93;
wire n_95;
wire n_141;
wire n_139;
wire n_33;
wire n_65;
wire n_142;
wire n_76;
wire n_67;
wire n_79;
wire n_107;
wire n_66;
wire n_136;
wire n_44;
wire n_28;
wire n_62;
wire n_121;
wire n_106;
wire n_45;
wire n_112;
wire n_42;
wire n_145;
wire n_77;
wire n_109;
wire n_39;
wire n_122;
wire n_94;
wire n_26;
wire n_118;
wire n_123;
wire n_116;
wire n_50;
wire n_143;
wire n_69;
wire n_31;
wire n_137;
wire n_129;
wire n_135;
wire n_134;
wire n_72;
wire n_100;
wire n_51;
wire n_71;
wire n_90;
wire n_110;
wire n_61;
wire n_117;
wire n_99;
wire n_86;
wire n_70;
wire n_41;
wire n_80;
wire n_74;
wire n_32;
wire n_30;
wire n_144;
wire n_130;
wire n_103;
wire n_43;
wire n_57;
wire n_84;
wire n_82;
wire n_111;
wire n_132;
wire n_125;
wire n_55;
wire n_58;
wire n_52;
wire n_63;
wire n_124;
wire n_92;
wire n_97;
wire n_75;
wire n_34;
wire n_60;
wire n_46;
wire n_88;
wire n_59;
wire n_128;
wire n_133;
wire n_138;
wire n_53;
wire n_127;
wire n_119;
wire n_36;
wire n_102;
wire n_81;
wire n_85;
wire n_101;
wire n_96;
wire n_89;

INVx5_ASAP7_75t_L g33 ( 
.A(n_0),
.Y(n_33)
);

BUFx5_ASAP7_75t_L g52 ( 
.A(n_0),
.Y(n_52)
);

BUFx5_ASAP7_75t_L g58 ( 
.A(n_0),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g71 ( 
.A(n_0),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_SL g91 ( 
.A(n_0),
.B(n_92),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_SL g29 ( 
.A(n_1),
.B(n_30),
.Y(n_29)
);

NAND2xp5_ASAP7_75t_L g34 ( 
.A(n_1),
.B(n_30),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_2),
.B(n_91),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_L g93 ( 
.A(n_2),
.B(n_91),
.Y(n_93)
);

CKINVDCx20_ASAP7_75t_R g101 ( 
.A(n_3),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_SL g47 ( 
.A(n_4),
.B(n_48),
.Y(n_47)
);

NAND2xp5_ASAP7_75t_L g115 ( 
.A(n_4),
.B(n_48),
.Y(n_115)
);

CKINVDCx20_ASAP7_75t_R g79 ( 
.A(n_5),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_SL g38 ( 
.A(n_6),
.B(n_39),
.Y(n_38)
);

AND2x2_ASAP7_75t_L g116 ( 
.A(n_6),
.B(n_39),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_SL g129 ( 
.A(n_7),
.B(n_130),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_L g142 ( 
.A(n_7),
.B(n_130),
.Y(n_142)
);

CKINVDCx20_ASAP7_75t_R g135 ( 
.A(n_8),
.Y(n_135)
);

CKINVDCx20_ASAP7_75t_R g125 ( 
.A(n_9),
.Y(n_125)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_10),
.Y(n_31)
);

NOR2xp33_ASAP7_75t_L g43 ( 
.A(n_11),
.B(n_44),
.Y(n_43)
);

AND2x2_ASAP7_75t_L g118 ( 
.A(n_11),
.B(n_44),
.Y(n_118)
);

CKINVDCx20_ASAP7_75t_R g131 ( 
.A(n_12),
.Y(n_131)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_13),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_14),
.Y(n_45)
);

AND2x2_ASAP7_75t_L g82 ( 
.A(n_15),
.B(n_83),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_SL g67 ( 
.A(n_16),
.B(n_68),
.Y(n_67)
);

AND2x2_ASAP7_75t_L g97 ( 
.A(n_16),
.B(n_68),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_17),
.B(n_104),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_L g109 ( 
.A(n_17),
.B(n_104),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_18),
.B(n_54),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_L g114 ( 
.A(n_18),
.B(n_54),
.Y(n_114)
);

CKINVDCx20_ASAP7_75t_R g121 ( 
.A(n_19),
.Y(n_121)
);

OR2x2_ASAP7_75t_L g119 ( 
.A(n_20),
.B(n_120),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_L g141 ( 
.A(n_20),
.B(n_120),
.Y(n_141)
);

CKINVDCx20_ASAP7_75t_R g88 ( 
.A(n_21),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_SL g63 ( 
.A(n_22),
.B(n_64),
.Y(n_63)
);

AND2x2_ASAP7_75t_L g96 ( 
.A(n_22),
.B(n_64),
.Y(n_96)
);

CKINVDCx20_ASAP7_75t_R g127 ( 
.A(n_23),
.Y(n_127)
);

CKINVDCx20_ASAP7_75t_R g138 ( 
.A(n_24),
.Y(n_138)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_26),
.Y(n_25)
);

OAI22xp5_ASAP7_75t_L g26 ( 
.A1(n_27),
.A2(n_35),
.B1(n_145),
.B2(n_146),
.Y(n_26)
);

CKINVDCx16_ASAP7_75t_R g145 ( 
.A(n_27),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_SL g27 ( 
.A(n_28),
.B(n_34),
.Y(n_27)
);

INVxp67_ASAP7_75t_L g28 ( 
.A(n_29),
.Y(n_28)
);

NOR2xp33_ASAP7_75t_L g30 ( 
.A(n_31),
.B(n_32),
.Y(n_30)
);

INVx2_ASAP7_75t_L g32 ( 
.A(n_33),
.Y(n_32)
);

BUFx3_ASAP7_75t_L g42 ( 
.A(n_33),
.Y(n_42)
);

INVx11_ASAP7_75t_L g46 ( 
.A(n_33),
.Y(n_46)
);

INVx4_ASAP7_75t_L g66 ( 
.A(n_33),
.Y(n_66)
);

INVx5_ASAP7_75t_L g78 ( 
.A(n_33),
.Y(n_78)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_35),
.Y(n_146)
);

OAI21xp5_ASAP7_75t_SL g35 ( 
.A1(n_36),
.A2(n_123),
.B(n_139),
.Y(n_35)
);

A2O1A1Ixp33_ASAP7_75t_L g36 ( 
.A1(n_37),
.A2(n_59),
.B(n_110),
.C(n_119),
.Y(n_36)
);

NOR4xp25_ASAP7_75t_L g37 ( 
.A(n_38),
.B(n_43),
.C(n_47),
.D(n_53),
.Y(n_37)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_38),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_L g39 ( 
.A(n_40),
.B(n_41),
.Y(n_39)
);

INVx3_ASAP7_75t_L g41 ( 
.A(n_42),
.Y(n_41)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_43),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_L g44 ( 
.A(n_45),
.B(n_46),
.Y(n_44)
);

BUFx3_ASAP7_75t_L g122 ( 
.A(n_46),
.Y(n_122)
);

OAI21xp5_ASAP7_75t_L g113 ( 
.A1(n_47),
.A2(n_114),
.B(n_115),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_49),
.B(n_50),
.Y(n_48)
);

OR2x2_ASAP7_75t_L g99 ( 
.A(n_50),
.B(n_100),
.Y(n_99)
);

OR2x2_ASAP7_75t_L g126 ( 
.A(n_50),
.B(n_127),
.Y(n_126)
);

INVx4_ASAP7_75t_L g50 ( 
.A(n_51),
.Y(n_50)
);

INVx2_ASAP7_75t_L g51 ( 
.A(n_52),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_55),
.B(n_56),
.Y(n_54)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_57),
.Y(n_56)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_58),
.Y(n_57)
);

OR2x2_ASAP7_75t_L g86 ( 
.A(n_58),
.B(n_87),
.Y(n_86)
);

OAI21x1_ASAP7_75t_L g59 ( 
.A1(n_60),
.A2(n_103),
.B(n_109),
.Y(n_59)
);

AOI21xp5_ASAP7_75t_L g60 ( 
.A1(n_61),
.A2(n_98),
.B(n_102),
.Y(n_60)
);

AO221x1_ASAP7_75t_L g61 ( 
.A1(n_62),
.A2(n_72),
.B1(n_95),
.B2(n_96),
.C(n_97),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_63),
.B(n_67),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_65),
.B(n_66),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_66),
.B(n_84),
.Y(n_83)
);

INVx6_ASAP7_75t_L g108 ( 
.A(n_66),
.Y(n_108)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_67),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_69),
.B(n_70),
.Y(n_68)
);

BUFx8_ASAP7_75t_L g132 ( 
.A(n_70),
.Y(n_132)
);

INVx3_ASAP7_75t_L g137 ( 
.A(n_70),
.Y(n_137)
);

BUFx12f_ASAP7_75t_L g70 ( 
.A(n_71),
.Y(n_70)
);

AO21x1_ASAP7_75t_L g72 ( 
.A1(n_73),
.A2(n_80),
.B(n_94),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_SL g73 ( 
.A(n_74),
.B(n_79),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_74),
.B(n_79),
.Y(n_94)
);

OR2x2_ASAP7_75t_L g74 ( 
.A(n_75),
.B(n_76),
.Y(n_74)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_77),
.Y(n_76)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_78),
.Y(n_77)
);

OAI21xp5_ASAP7_75t_L g80 ( 
.A1(n_81),
.A2(n_90),
.B(n_93),
.Y(n_80)
);

AOI21xp5_ASAP7_75t_L g81 ( 
.A1(n_82),
.A2(n_85),
.B(n_89),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_SL g85 ( 
.A(n_86),
.B(n_88),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_86),
.B(n_88),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_SL g98 ( 
.A(n_99),
.B(n_101),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_99),
.B(n_101),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_105),
.B(n_106),
.Y(n_104)
);

BUFx2_ASAP7_75t_L g106 ( 
.A(n_107),
.Y(n_106)
);

INVx8_ASAP7_75t_L g107 ( 
.A(n_108),
.Y(n_107)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_111),
.Y(n_110)
);

A2O1A1O1Ixp25_ASAP7_75t_L g111 ( 
.A1(n_112),
.A2(n_113),
.B(n_116),
.C(n_117),
.D(n_118),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_L g120 ( 
.A(n_121),
.B(n_122),
.Y(n_120)
);

NAND3xp33_ASAP7_75t_L g123 ( 
.A(n_124),
.B(n_128),
.C(n_133),
.Y(n_123)
);

A2O1A1O1Ixp25_ASAP7_75t_L g139 ( 
.A1(n_124),
.A2(n_133),
.B(n_140),
.C(n_143),
.D(n_144),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_L g124 ( 
.A(n_125),
.B(n_126),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_L g144 ( 
.A(n_125),
.B(n_126),
.Y(n_144)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_129),
.Y(n_128)
);

OAI21xp5_ASAP7_75t_L g140 ( 
.A1(n_129),
.A2(n_141),
.B(n_142),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_L g130 ( 
.A(n_131),
.B(n_132),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_SL g133 ( 
.A(n_134),
.B(n_138),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_L g143 ( 
.A(n_134),
.B(n_138),
.Y(n_143)
);

OR2x2_ASAP7_75t_L g134 ( 
.A(n_135),
.B(n_136),
.Y(n_134)
);

INVx8_ASAP7_75t_L g136 ( 
.A(n_137),
.Y(n_136)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_148),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g55 ( 
.A(n_149),
.Y(n_55)
);

CKINVDCx20_ASAP7_75t_R g65 ( 
.A(n_150),
.Y(n_65)
);

CKINVDCx20_ASAP7_75t_R g69 ( 
.A(n_151),
.Y(n_69)
);

CKINVDCx20_ASAP7_75t_R g75 ( 
.A(n_152),
.Y(n_75)
);

CKINVDCx20_ASAP7_75t_R g84 ( 
.A(n_153),
.Y(n_84)
);

CKINVDCx20_ASAP7_75t_R g87 ( 
.A(n_154),
.Y(n_87)
);

CKINVDCx20_ASAP7_75t_R g92 ( 
.A(n_155),
.Y(n_92)
);

CKINVDCx20_ASAP7_75t_R g100 ( 
.A(n_156),
.Y(n_100)
);

CKINVDCx20_ASAP7_75t_R g105 ( 
.A(n_157),
.Y(n_105)
);


endmodule