module real_aes_1044_n_104 (n_17, n_28, n_76, n_56, n_34, n_98, n_90, n_82, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_83, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_91, n_100, n_43, n_103, n_96, n_54, n_35, n_42, n_99, n_15, n_9, n_23, n_72, n_95, n_44, n_102, n_7, n_4, n_80, n_6, n_12, n_68, n_79, n_69, n_46, n_59, n_25, n_73, n_77, n_81, n_48, n_37, n_97, n_70, n_50, n_89, n_26, n_86, n_93, n_13, n_24, n_2, n_55, n_62, n_84, n_67, n_92, n_33, n_88, n_14, n_11, n_85, n_16, n_94, n_39, n_5, n_45, n_60, n_38, n_87, n_0, n_78, n_101, n_63, n_1, n_53, n_36, n_104);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_98;
input n_90;
input n_82;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_83;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_91;
input n_100;
input n_43;
input n_103;
input n_96;
input n_54;
input n_35;
input n_42;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_95;
input n_44;
input n_102;
input n_7;
input n_4;
input n_80;
input n_6;
input n_12;
input n_68;
input n_79;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_81;
input n_48;
input n_37;
input n_97;
input n_70;
input n_50;
input n_89;
input n_26;
input n_86;
input n_93;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_84;
input n_67;
input n_92;
input n_33;
input n_88;
input n_14;
input n_11;
input n_85;
input n_16;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_87;
input n_0;
input n_78;
input n_101;
input n_63;
input n_1;
input n_53;
input n_36;
output n_104;
wire n_480;
wire n_113;
wire n_476;
wire n_758;
wire n_599;
wire n_187;
wire n_436;
wire n_684;
wire n_257;
wire n_390;
wire n_821;
wire n_185;
wire n_285;
wire n_624;
wire n_618;
wire n_778;
wire n_800;
wire n_522;
wire n_485;
wire n_822;
wire n_222;
wire n_750;
wire n_631;
wire n_287;
wire n_357;
wire n_503;
wire n_792;
wire n_386;
wire n_635;
wire n_673;
wire n_518;
wire n_254;
wire n_207;
wire n_665;
wire n_667;
wire n_577;
wire n_580;
wire n_469;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_759;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_718;
wire n_318;
wire n_355;
wire n_239;
wire n_669;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_761;
wire n_742;
wire n_112;
wire n_364;
wire n_319;
wire n_421;
wire n_555;
wire n_329;
wire n_766;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_169;
wire n_242;
wire n_571;
wire n_376;
wire n_549;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_752;
wire n_448;
wire n_556;
wire n_545;
wire n_341;
wire n_593;
wire n_232;
wire n_460;
wire n_773;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_537;
wire n_320;
wire n_551;
wire n_666;
wire n_560;
wire n_260;
wire n_660;
wire n_814;
wire n_594;
wire n_186;
wire n_767;
wire n_138;
wire n_696;
wire n_704;
wire n_379;
wire n_374;
wire n_453;
wire n_647;
wire n_235;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_775;
wire n_161;
wire n_763;
wire n_189;
wire n_271;
wire n_489;
wire n_548;
wire n_427;
wire n_678;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_815;
wire n_519;
wire n_564;
wire n_638;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_786;
wire n_512;
wire n_395;
wire n_332;
wire n_795;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_816;
wire n_116;
wire n_625;
wire n_289;
wire n_462;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_818;
wire n_716;
wire n_213;
wire n_478;
wire n_356;
wire n_584;
wire n_408;
wire n_553;
wire n_184;
wire n_372;
wire n_528;
wire n_578;
wire n_202;
wire n_495;
wire n_370;
wire n_384;
wire n_744;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_824;
wire n_467;
wire n_327;
wire n_774;
wire n_813;
wire n_106;
wire n_791;
wire n_559;
wire n_466;
wire n_636;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_726;
wire n_517;
wire n_683;
wire n_780;
wire n_174;
wire n_570;
wire n_675;
wire n_530;
wire n_535;
wire n_732;
wire n_784;
wire n_211;
wire n_281;
wire n_496;
wire n_693;
wire n_173;
wire n_468;
wire n_234;
wire n_746;
wire n_284;
wire n_153;
wire n_532;
wire n_316;
wire n_656;
wire n_755;
wire n_178;
wire n_409;
wire n_748;
wire n_781;
wire n_523;
wire n_298;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_796;
wire n_297;
wire n_801;
wire n_383;
wire n_529;
wire n_119;
wire n_310;
wire n_455;
wire n_504;
wire n_725;
wire n_164;
wire n_671;
wire n_231;
wire n_547;
wire n_659;
wire n_634;
wire n_682;
wire n_454;
wire n_122;
wire n_812;
wire n_817;
wire n_443;
wire n_565;
wire n_782;
wire n_760;
wire n_608;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_819;
wire n_267;
wire n_218;
wire n_737;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_808;
wire n_770;
wire n_722;
wire n_745;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_331;
wire n_449;
wire n_182;
wire n_363;
wire n_417;
wire n_607;
wire n_754;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_142;
wire n_561;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_783;
wire n_655;
wire n_654;
wire n_527;
wire n_502;
wire n_434;
wire n_505;
wire n_769;
wire n_600;
wire n_731;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_602;
wire n_402;
wire n_552;
wire n_617;
wire n_733;
wire n_171;
wire n_658;
wire n_676;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_146;
wire n_432;
wire n_807;
wire n_226;
wire n_255;
wire n_286;
wire n_416;
wire n_790;
wire n_410;
wire n_120;
wire n_799;
wire n_805;
wire n_751;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_695;
wire n_685;
wire n_165;
wire n_361;
wire n_632;
wire n_246;
wire n_176;
wire n_768;
wire n_412;
wire n_163;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_777;
wire n_501;
wire n_488;
wire n_251;
wire n_642;
wire n_613;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_702;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_734;
wire n_110;
wire n_392;
wire n_562;
wire n_150;
wire n_147;
wire n_404;
wire n_288;
wire n_598;
wire n_713;
wire n_728;
wire n_735;
wire n_756;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_569;
wire n_563;
wire n_785;
wire n_188;
wire n_269;
wire n_430;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_810;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_193;
wire n_397;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_649;
wire n_663;
wire n_749;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_707;
wire n_622;
wire n_470;
wire n_133;
wire n_494;
wire n_711;
wire n_377;
wire n_273;
wire n_723;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_265;
wire n_354;
wire n_720;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_730;
wire n_643;
wire n_747;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_779;
wire n_148;
wire n_498;
wire n_481;
wire n_691;
wire n_765;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_487;
wire n_233;
wire n_290;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_155;
wire n_243;
wire n_692;
wire n_544;
wire n_268;
wire n_789;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_738;
wire n_701;
wire n_309;
wire n_344;
wire n_107;
wire n_229;
wire n_809;
wire n_482;
wire n_520;
wire n_633;
wire n_679;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_787;
wire n_262;
wire n_630;
wire n_806;
wire n_689;
wire n_820;
wire n_715;
wire n_134;
wire n_349;
wire n_336;
wire n_420;
wire n_612;
wire n_195;
wire n_438;
wire n_764;
wire n_794;
wire n_300;
wire n_252;
wire n_283;
wire n_314;
wire n_741;
wire n_753;
wire n_249;
wire n_623;
wire n_446;
wire n_721;
wire n_221;
wire n_681;
wire n_156;
wire n_456;
wire n_359;
wire n_717;
wire n_312;
wire n_183;
wire n_266;
wire n_712;
wire n_205;
wire n_433;
wire n_335;
wire n_177;
wire n_516;
wire n_313;
wire n_627;
wire n_739;
wire n_140;
wire n_418;
wire n_521;
wire n_422;
wire n_771;
wire n_524;
wire n_219;
wire n_705;
wire n_180;
wire n_212;
wire n_210;
wire n_575;
wire n_325;
wire n_762;
wire n_338;
wire n_479;
wire n_442;
wire n_825;
wire n_698;
wire n_371;
wire n_740;
wire n_541;
wire n_166;
wire n_224;
wire n_151;
wire n_546;
wire n_587;
wire n_639;
wire n_811;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_724;
wire n_440;
wire n_525;
wire n_674;
wire n_644;
wire n_152;
wire n_198;
wire n_793;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_414;
wire n_757;
wire n_123;
wire n_279;
wire n_686;
wire n_776;
wire n_803;
wire n_543;
wire n_497;
wire n_514;
wire n_270;
wire n_507;
wire n_614;
wire n_305;
wire n_586;
wire n_772;
wire n_450;
wire n_788;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_465;
wire n_473;
wire n_719;
wire n_566;
wire n_474;
wire n_170;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_168;
wire n_175;
wire n_241;
wire n_687;
wire n_729;
wire n_646;
wire n_710;
wire n_650;
wire n_105;
wire n_743;
wire n_823;
wire n_393;
wire n_294;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_500;
wire n_307;
wire n_601;
wire n_661;
wire n_463;
wire n_396;
wire n_804;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_802;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_143;
wire n_192;
wire n_475;
wire n_554;
wire n_264;
wire n_798;
wire n_237;
wire n_668;
wire n_797;
NAND2xp5_ASAP7_75t_SL g219 ( .A(n_0), .B(n_162), .Y(n_219) );
AOI21xp5_ASAP7_75t_L g194 ( .A1(n_1), .A2(n_144), .B(n_195), .Y(n_194) );
AOI22xp33_ASAP7_75t_L g464 ( .A1(n_2), .A2(n_465), .B1(n_470), .B2(n_815), .Y(n_464) );
NAND2xp5_ASAP7_75t_L g113 ( .A(n_3), .B(n_114), .Y(n_113) );
AOI22xp5_ASAP7_75t_L g128 ( .A1(n_4), .A2(n_11), .B1(n_129), .B2(n_130), .Y(n_128) );
CKINVDCx20_ASAP7_75t_R g130 ( .A(n_4), .Y(n_130) );
NAND2xp5_ASAP7_75t_SL g208 ( .A(n_5), .B(n_152), .Y(n_208) );
INVx1_ASAP7_75t_L g149 ( .A(n_6), .Y(n_149) );
NAND2xp5_ASAP7_75t_L g172 ( .A(n_7), .B(n_152), .Y(n_172) );
AOI22xp5_ASAP7_75t_L g123 ( .A1(n_8), .A2(n_124), .B1(n_448), .B2(n_449), .Y(n_123) );
INVxp67_ASAP7_75t_L g449 ( .A(n_8), .Y(n_449) );
NAND2xp5_ASAP7_75t_SL g506 ( .A(n_8), .B(n_139), .Y(n_506) );
INVx1_ASAP7_75t_L g534 ( .A(n_9), .Y(n_534) );
CKINVDCx16_ASAP7_75t_R g114 ( .A(n_10), .Y(n_114) );
CKINVDCx20_ASAP7_75t_R g129 ( .A(n_11), .Y(n_129) );
CKINVDCx5p33_ASAP7_75t_R g549 ( .A(n_12), .Y(n_549) );
NAND2xp33_ASAP7_75t_L g189 ( .A(n_13), .B(n_156), .Y(n_189) );
INVx2_ASAP7_75t_L g141 ( .A(n_14), .Y(n_141) );
AOI221x1_ASAP7_75t_L g231 ( .A1(n_15), .A2(n_29), .B1(n_144), .B2(n_162), .C(n_232), .Y(n_231) );
NOR3xp33_ASAP7_75t_L g112 ( .A(n_16), .B(n_113), .C(n_115), .Y(n_112) );
CKINVDCx16_ASAP7_75t_R g453 ( .A(n_16), .Y(n_453) );
NAND2xp5_ASAP7_75t_SL g185 ( .A(n_17), .B(n_162), .Y(n_185) );
AO21x2_ASAP7_75t_L g182 ( .A1(n_18), .A2(n_183), .B(n_184), .Y(n_182) );
INVx1_ASAP7_75t_L g515 ( .A(n_19), .Y(n_515) );
NAND2xp5_ASAP7_75t_L g235 ( .A(n_20), .B(n_175), .Y(n_235) );
NAND2xp5_ASAP7_75t_L g151 ( .A(n_21), .B(n_152), .Y(n_151) );
AO21x1_ASAP7_75t_L g203 ( .A1(n_22), .A2(n_162), .B(n_204), .Y(n_203) );
INVx1_ASAP7_75t_L g110 ( .A(n_23), .Y(n_110) );
NAND2xp5_ASAP7_75t_L g456 ( .A(n_24), .B(n_457), .Y(n_456) );
INVx1_ASAP7_75t_L g513 ( .A(n_25), .Y(n_513) );
INVx1_ASAP7_75t_SL g499 ( .A(n_26), .Y(n_499) );
CKINVDCx20_ASAP7_75t_R g824 ( .A(n_27), .Y(n_824) );
NAND2xp5_ASAP7_75t_SL g593 ( .A(n_28), .B(n_163), .Y(n_593) );
NAND2x1_ASAP7_75t_L g217 ( .A(n_30), .B(n_152), .Y(n_217) );
AOI33xp33_ASAP7_75t_L g561 ( .A1(n_31), .A2(n_56), .A3(n_489), .B1(n_496), .B2(n_562), .B3(n_563), .Y(n_561) );
NAND2x1_ASAP7_75t_L g171 ( .A(n_32), .B(n_156), .Y(n_171) );
INVx1_ASAP7_75t_L g543 ( .A(n_33), .Y(n_543) );
OR2x2_ASAP7_75t_L g140 ( .A(n_34), .B(n_90), .Y(n_140) );
OA21x2_ASAP7_75t_L g180 ( .A1(n_34), .A2(n_90), .B(n_141), .Y(n_180) );
NAND2xp5_ASAP7_75t_L g486 ( .A(n_35), .B(n_487), .Y(n_486) );
NAND2xp5_ASAP7_75t_L g197 ( .A(n_36), .B(n_156), .Y(n_197) );
NAND2xp5_ASAP7_75t_L g188 ( .A(n_37), .B(n_152), .Y(n_188) );
NAND2xp5_ASAP7_75t_L g207 ( .A(n_38), .B(n_156), .Y(n_207) );
AOI21xp5_ASAP7_75t_L g249 ( .A1(n_39), .A2(n_144), .B(n_250), .Y(n_249) );
AND2x2_ASAP7_75t_L g145 ( .A(n_40), .B(n_146), .Y(n_145) );
AND2x2_ASAP7_75t_L g160 ( .A(n_40), .B(n_149), .Y(n_160) );
INVx1_ASAP7_75t_L g495 ( .A(n_40), .Y(n_495) );
INVxp67_ASAP7_75t_L g115 ( .A(n_41), .Y(n_115) );
OR2x6_ASAP7_75t_L g455 ( .A(n_41), .B(n_109), .Y(n_455) );
XNOR2xp5_ASAP7_75t_L g466 ( .A(n_42), .B(n_467), .Y(n_466) );
CKINVDCx20_ASAP7_75t_R g545 ( .A(n_43), .Y(n_545) );
NAND2xp5_ASAP7_75t_SL g253 ( .A(n_44), .B(n_162), .Y(n_253) );
NAND2xp5_ASAP7_75t_L g569 ( .A(n_45), .B(n_487), .Y(n_569) );
AOI22xp5_ASAP7_75t_L g586 ( .A1(n_46), .A2(n_139), .B1(n_179), .B2(n_587), .Y(n_586) );
NAND2xp5_ASAP7_75t_L g594 ( .A(n_47), .B(n_595), .Y(n_594) );
NAND2xp5_ASAP7_75t_L g501 ( .A(n_48), .B(n_163), .Y(n_501) );
CKINVDCx20_ASAP7_75t_R g165 ( .A(n_49), .Y(n_165) );
NAND2xp5_ASAP7_75t_L g251 ( .A(n_50), .B(n_156), .Y(n_251) );
NAND2xp5_ASAP7_75t_SL g536 ( .A(n_51), .B(n_183), .Y(n_536) );
NAND2xp5_ASAP7_75t_L g535 ( .A(n_52), .B(n_163), .Y(n_535) );
AOI21xp5_ASAP7_75t_L g169 ( .A1(n_53), .A2(n_144), .B(n_170), .Y(n_169) );
CKINVDCx5p33_ASAP7_75t_R g590 ( .A(n_54), .Y(n_590) );
NAND2xp5_ASAP7_75t_L g218 ( .A(n_55), .B(n_156), .Y(n_218) );
NAND2xp5_ASAP7_75t_L g573 ( .A(n_57), .B(n_163), .Y(n_573) );
INVx1_ASAP7_75t_L g148 ( .A(n_58), .Y(n_148) );
INVx1_ASAP7_75t_L g158 ( .A(n_58), .Y(n_158) );
AND2x2_ASAP7_75t_L g574 ( .A(n_59), .B(n_175), .Y(n_574) );
AOI221xp5_ASAP7_75t_L g532 ( .A1(n_60), .A2(n_77), .B1(n_487), .B2(n_493), .C(n_533), .Y(n_532) );
NAND2xp5_ASAP7_75t_L g527 ( .A(n_61), .B(n_487), .Y(n_527) );
NAND2xp5_ASAP7_75t_L g234 ( .A(n_62), .B(n_152), .Y(n_234) );
NAND2xp5_ASAP7_75t_L g551 ( .A(n_63), .B(n_179), .Y(n_551) );
AOI21xp5_ASAP7_75t_SL g523 ( .A1(n_64), .A2(n_493), .B(n_524), .Y(n_523) );
AOI21xp5_ASAP7_75t_L g215 ( .A1(n_65), .A2(n_144), .B(n_216), .Y(n_215) );
INVx1_ASAP7_75t_L g509 ( .A(n_66), .Y(n_509) );
AO21x1_ASAP7_75t_L g205 ( .A1(n_67), .A2(n_144), .B(n_206), .Y(n_205) );
NAND2xp5_ASAP7_75t_SL g193 ( .A(n_68), .B(n_162), .Y(n_193) );
INVx1_ASAP7_75t_L g572 ( .A(n_69), .Y(n_572) );
NAND2xp5_ASAP7_75t_SL g173 ( .A(n_70), .B(n_162), .Y(n_173) );
AOI21xp5_ASAP7_75t_L g570 ( .A1(n_71), .A2(n_493), .B(n_571), .Y(n_570) );
AND2x2_ASAP7_75t_L g254 ( .A(n_72), .B(n_176), .Y(n_254) );
INVx1_ASAP7_75t_L g146 ( .A(n_73), .Y(n_146) );
INVx1_ASAP7_75t_L g154 ( .A(n_73), .Y(n_154) );
AOI22xp5_ASAP7_75t_L g467 ( .A1(n_74), .A2(n_100), .B1(n_468), .B2(n_469), .Y(n_467) );
CKINVDCx20_ASAP7_75t_R g468 ( .A(n_74), .Y(n_468) );
AND2x2_ASAP7_75t_L g177 ( .A(n_75), .B(n_178), .Y(n_177) );
NAND2xp5_ASAP7_75t_L g564 ( .A(n_76), .B(n_487), .Y(n_564) );
AND2x2_ASAP7_75t_L g502 ( .A(n_78), .B(n_178), .Y(n_502) );
INVx1_ASAP7_75t_L g510 ( .A(n_79), .Y(n_510) );
AOI21xp5_ASAP7_75t_L g492 ( .A1(n_80), .A2(n_493), .B(n_498), .Y(n_492) );
A2O1A1Ixp33_ASAP7_75t_L g591 ( .A1(n_81), .A2(n_493), .B(n_556), .C(n_592), .Y(n_591) );
INVx1_ASAP7_75t_L g111 ( .A(n_82), .Y(n_111) );
NAND2xp5_ASAP7_75t_SL g161 ( .A(n_83), .B(n_162), .Y(n_161) );
AND2x2_ASAP7_75t_L g191 ( .A(n_84), .B(n_178), .Y(n_191) );
AND2x2_ASAP7_75t_SL g521 ( .A(n_85), .B(n_178), .Y(n_521) );
AOI22xp5_ASAP7_75t_L g558 ( .A1(n_86), .A2(n_493), .B1(n_559), .B2(n_560), .Y(n_558) );
OAI22xp5_ASAP7_75t_SL g125 ( .A1(n_87), .A2(n_126), .B1(n_127), .B2(n_128), .Y(n_125) );
CKINVDCx20_ASAP7_75t_R g126 ( .A(n_87), .Y(n_126) );
XNOR2xp5_ASAP7_75t_L g465 ( .A(n_88), .B(n_466), .Y(n_465) );
AND2x2_ASAP7_75t_L g204 ( .A(n_89), .B(n_139), .Y(n_204) );
NAND2xp5_ASAP7_75t_L g155 ( .A(n_91), .B(n_156), .Y(n_155) );
AND2x2_ASAP7_75t_L g221 ( .A(n_92), .B(n_178), .Y(n_221) );
INVx1_ASAP7_75t_L g525 ( .A(n_93), .Y(n_525) );
NAND2xp5_ASAP7_75t_L g252 ( .A(n_94), .B(n_152), .Y(n_252) );
AOI21xp5_ASAP7_75t_L g143 ( .A1(n_95), .A2(n_144), .B(n_150), .Y(n_143) );
NAND2xp5_ASAP7_75t_L g233 ( .A(n_96), .B(n_156), .Y(n_233) );
AND2x2_ASAP7_75t_L g565 ( .A(n_97), .B(n_178), .Y(n_565) );
NAND2xp5_ASAP7_75t_L g196 ( .A(n_98), .B(n_152), .Y(n_196) );
A2O1A1Ixp33_ASAP7_75t_L g540 ( .A1(n_99), .A2(n_541), .B(n_542), .C(n_544), .Y(n_540) );
CKINVDCx20_ASAP7_75t_R g469 ( .A(n_100), .Y(n_469) );
BUFx2_ASAP7_75t_L g121 ( .A(n_101), .Y(n_121) );
BUFx2_ASAP7_75t_SL g462 ( .A(n_101), .Y(n_462) );
AOI21xp5_ASAP7_75t_L g186 ( .A1(n_102), .A2(n_144), .B(n_187), .Y(n_186) );
NAND2xp5_ASAP7_75t_L g526 ( .A(n_103), .B(n_163), .Y(n_526) );
AOI21xp33_ASAP7_75t_SL g104 ( .A1(n_105), .A2(n_116), .B(n_823), .Y(n_104) );
CKINVDCx5p33_ASAP7_75t_R g105 ( .A(n_106), .Y(n_105) );
INVx1_ASAP7_75t_SL g825 ( .A(n_106), .Y(n_825) );
INVx2_ASAP7_75t_SL g106 ( .A(n_107), .Y(n_106) );
AND2x2_ASAP7_75t_SL g107 ( .A(n_108), .B(n_112), .Y(n_107) );
INVx1_ASAP7_75t_L g108 ( .A(n_109), .Y(n_108) );
NAND2xp5_ASAP7_75t_L g109 ( .A(n_110), .B(n_111), .Y(n_109) );
OA22x2_ASAP7_75t_L g116 ( .A1(n_117), .A2(n_122), .B1(n_459), .B2(n_463), .Y(n_116) );
INVx1_ASAP7_75t_SL g117 ( .A(n_118), .Y(n_117) );
BUFx3_ASAP7_75t_L g118 ( .A(n_119), .Y(n_118) );
CKINVDCx20_ASAP7_75t_R g119 ( .A(n_120), .Y(n_119) );
HB1xp67_ASAP7_75t_L g120 ( .A(n_121), .Y(n_120) );
OAI21xp5_ASAP7_75t_L g122 ( .A1(n_123), .A2(n_450), .B(n_456), .Y(n_122) );
INVx1_ASAP7_75t_L g448 ( .A(n_124), .Y(n_448) );
XNOR2x1_ASAP7_75t_L g124 ( .A(n_125), .B(n_131), .Y(n_124) );
CKINVDCx20_ASAP7_75t_R g127 ( .A(n_128), .Y(n_127) );
OAI22xp5_ASAP7_75t_L g470 ( .A1(n_131), .A2(n_471), .B1(n_475), .B2(n_478), .Y(n_470) );
INVx2_ASAP7_75t_L g820 ( .A(n_131), .Y(n_820) );
OR2x6_ASAP7_75t_L g131 ( .A(n_132), .B(n_346), .Y(n_131) );
NAND3xp33_ASAP7_75t_SL g132 ( .A(n_133), .B(n_258), .C(n_313), .Y(n_132) );
AOI221xp5_ASAP7_75t_L g133 ( .A1(n_134), .A2(n_198), .B1(n_222), .B2(n_226), .C(n_236), .Y(n_133) );
AND2x2_ASAP7_75t_L g134 ( .A(n_135), .B(n_181), .Y(n_134) );
AND2x2_ASAP7_75t_SL g224 ( .A(n_135), .B(n_225), .Y(n_224) );
INVx2_ASAP7_75t_L g257 ( .A(n_135), .Y(n_257) );
AND2x2_ASAP7_75t_L g302 ( .A(n_135), .B(n_239), .Y(n_302) );
AND2x4_ASAP7_75t_L g135 ( .A(n_136), .B(n_166), .Y(n_135) );
INVx1_ASAP7_75t_L g136 ( .A(n_137), .Y(n_136) );
INVx2_ASAP7_75t_L g290 ( .A(n_137), .Y(n_290) );
INVx1_ASAP7_75t_L g300 ( .A(n_137), .Y(n_300) );
AO21x2_ASAP7_75t_L g137 ( .A1(n_138), .A2(n_142), .B(n_164), .Y(n_137) );
NOR2xp33_ASAP7_75t_L g164 ( .A(n_138), .B(n_165), .Y(n_164) );
AO21x2_ASAP7_75t_L g264 ( .A1(n_138), .A2(n_142), .B(n_164), .Y(n_264) );
INVx1_ASAP7_75t_SL g138 ( .A(n_139), .Y(n_138) );
AOI21xp5_ASAP7_75t_L g184 ( .A1(n_139), .A2(n_185), .B(n_186), .Y(n_184) );
NAND2xp5_ASAP7_75t_L g209 ( .A(n_139), .B(n_210), .Y(n_209) );
NOR2xp33_ASAP7_75t_L g517 ( .A(n_139), .B(n_159), .Y(n_517) );
AOI21xp5_ASAP7_75t_L g522 ( .A1(n_139), .A2(n_523), .B(n_527), .Y(n_522) );
AND2x4_ASAP7_75t_L g139 ( .A(n_140), .B(n_141), .Y(n_139) );
AND2x2_ASAP7_75t_SL g176 ( .A(n_140), .B(n_141), .Y(n_176) );
NAND2xp5_ASAP7_75t_L g142 ( .A(n_143), .B(n_161), .Y(n_142) );
AND2x6_ASAP7_75t_L g144 ( .A(n_145), .B(n_147), .Y(n_144) );
BUFx3_ASAP7_75t_L g491 ( .A(n_145), .Y(n_491) );
AND2x6_ASAP7_75t_L g156 ( .A(n_146), .B(n_157), .Y(n_156) );
INVx2_ASAP7_75t_L g497 ( .A(n_146), .Y(n_497) );
AND2x4_ASAP7_75t_L g493 ( .A(n_147), .B(n_494), .Y(n_493) );
AND2x2_ASAP7_75t_L g147 ( .A(n_148), .B(n_149), .Y(n_147) );
AND2x4_ASAP7_75t_L g152 ( .A(n_148), .B(n_153), .Y(n_152) );
INVx2_ASAP7_75t_L g489 ( .A(n_148), .Y(n_489) );
HB1xp67_ASAP7_75t_L g490 ( .A(n_149), .Y(n_490) );
AOI21xp5_ASAP7_75t_L g150 ( .A1(n_151), .A2(n_155), .B(n_159), .Y(n_150) );
INVxp67_ASAP7_75t_L g516 ( .A(n_152), .Y(n_516) );
AND2x4_ASAP7_75t_L g163 ( .A(n_153), .B(n_157), .Y(n_163) );
INVx2_ASAP7_75t_L g153 ( .A(n_154), .Y(n_153) );
INVxp67_ASAP7_75t_L g514 ( .A(n_156), .Y(n_514) );
INVx2_ASAP7_75t_L g157 ( .A(n_158), .Y(n_157) );
AOI21xp5_ASAP7_75t_L g170 ( .A1(n_159), .A2(n_171), .B(n_172), .Y(n_170) );
AOI21xp5_ASAP7_75t_L g187 ( .A1(n_159), .A2(n_188), .B(n_189), .Y(n_187) );
AOI21xp5_ASAP7_75t_L g195 ( .A1(n_159), .A2(n_196), .B(n_197), .Y(n_195) );
AOI21xp5_ASAP7_75t_L g206 ( .A1(n_159), .A2(n_207), .B(n_208), .Y(n_206) );
AOI21xp5_ASAP7_75t_L g216 ( .A1(n_159), .A2(n_217), .B(n_218), .Y(n_216) );
AOI21xp5_ASAP7_75t_L g232 ( .A1(n_159), .A2(n_233), .B(n_234), .Y(n_232) );
AOI21xp5_ASAP7_75t_L g250 ( .A1(n_159), .A2(n_251), .B(n_252), .Y(n_250) );
O2A1O1Ixp33_ASAP7_75t_SL g498 ( .A1(n_159), .A2(n_499), .B(n_500), .C(n_501), .Y(n_498) );
O2A1O1Ixp33_ASAP7_75t_L g524 ( .A1(n_159), .A2(n_500), .B(n_525), .C(n_526), .Y(n_524) );
O2A1O1Ixp33_ASAP7_75t_SL g533 ( .A1(n_159), .A2(n_500), .B(n_534), .C(n_535), .Y(n_533) );
INVx1_ASAP7_75t_L g559 ( .A(n_159), .Y(n_559) );
O2A1O1Ixp33_ASAP7_75t_L g571 ( .A1(n_159), .A2(n_500), .B(n_572), .C(n_573), .Y(n_571) );
AOI21xp5_ASAP7_75t_L g592 ( .A1(n_159), .A2(n_593), .B(n_594), .Y(n_592) );
INVx5_ASAP7_75t_L g159 ( .A(n_160), .Y(n_159) );
AND2x4_ASAP7_75t_L g162 ( .A(n_160), .B(n_163), .Y(n_162) );
HB1xp67_ASAP7_75t_L g544 ( .A(n_160), .Y(n_544) );
INVx1_ASAP7_75t_L g511 ( .A(n_163), .Y(n_511) );
OR2x2_ASAP7_75t_L g279 ( .A(n_166), .B(n_182), .Y(n_279) );
NAND2x1p5_ASAP7_75t_L g310 ( .A(n_166), .B(n_225), .Y(n_310) );
NAND2xp5_ASAP7_75t_L g323 ( .A(n_166), .B(n_190), .Y(n_323) );
INVx2_ASAP7_75t_L g332 ( .A(n_166), .Y(n_332) );
AND2x2_ASAP7_75t_L g353 ( .A(n_166), .B(n_354), .Y(n_353) );
AND2x2_ASAP7_75t_L g437 ( .A(n_166), .B(n_256), .Y(n_437) );
INVx4_ASAP7_75t_L g166 ( .A(n_167), .Y(n_166) );
AND2x2_ASAP7_75t_L g265 ( .A(n_167), .B(n_190), .Y(n_265) );
AND2x2_ASAP7_75t_L g398 ( .A(n_167), .B(n_225), .Y(n_398) );
HB1xp67_ASAP7_75t_L g424 ( .A(n_167), .Y(n_424) );
AO21x2_ASAP7_75t_L g167 ( .A1(n_168), .A2(n_174), .B(n_177), .Y(n_167) );
NAND2xp5_ASAP7_75t_L g168 ( .A(n_169), .B(n_173), .Y(n_168) );
AO21x2_ASAP7_75t_L g484 ( .A1(n_174), .A2(n_485), .B(n_502), .Y(n_484) );
CKINVDCx5p33_ASAP7_75t_R g174 ( .A(n_175), .Y(n_174) );
AOI21xp5_ASAP7_75t_L g192 ( .A1(n_175), .A2(n_193), .B(n_194), .Y(n_192) );
OA21x2_ASAP7_75t_L g230 ( .A1(n_175), .A2(n_231), .B(n_235), .Y(n_230) );
OA21x2_ASAP7_75t_L g242 ( .A1(n_175), .A2(n_231), .B(n_235), .Y(n_242) );
BUFx6f_ASAP7_75t_L g175 ( .A(n_176), .Y(n_175) );
INVx3_ASAP7_75t_L g220 ( .A(n_178), .Y(n_220) );
OAI22xp5_ASAP7_75t_L g539 ( .A1(n_178), .A2(n_220), .B1(n_540), .B2(n_545), .Y(n_539) );
INVx4_ASAP7_75t_L g178 ( .A(n_179), .Y(n_178) );
NAND2xp5_ASAP7_75t_L g547 ( .A(n_179), .B(n_548), .Y(n_547) );
INVx3_ASAP7_75t_L g179 ( .A(n_180), .Y(n_179) );
BUFx4f_ASAP7_75t_L g183 ( .A(n_180), .Y(n_183) );
AND2x4_ASAP7_75t_L g352 ( .A(n_181), .B(n_353), .Y(n_352) );
AOI321xp33_ASAP7_75t_L g366 ( .A1(n_181), .A2(n_295), .A3(n_296), .B1(n_328), .B2(n_367), .C(n_370), .Y(n_366) );
AND2x2_ASAP7_75t_L g181 ( .A(n_182), .B(n_190), .Y(n_181) );
BUFx3_ASAP7_75t_L g223 ( .A(n_182), .Y(n_223) );
INVx2_ASAP7_75t_L g256 ( .A(n_182), .Y(n_256) );
NAND2xp5_ASAP7_75t_L g263 ( .A(n_182), .B(n_264), .Y(n_263) );
AND2x2_ASAP7_75t_L g289 ( .A(n_182), .B(n_290), .Y(n_289) );
INVx1_ASAP7_75t_L g322 ( .A(n_182), .Y(n_322) );
OA21x2_ASAP7_75t_L g531 ( .A1(n_183), .A2(n_532), .B(n_536), .Y(n_531) );
INVx2_ASAP7_75t_SL g556 ( .A(n_183), .Y(n_556) );
INVx5_ASAP7_75t_L g225 ( .A(n_190), .Y(n_225) );
NOR2x1_ASAP7_75t_SL g274 ( .A(n_190), .B(n_264), .Y(n_274) );
BUFx2_ASAP7_75t_L g369 ( .A(n_190), .Y(n_369) );
OR2x6_ASAP7_75t_L g190 ( .A(n_191), .B(n_192), .Y(n_190) );
INVxp67_ASAP7_75t_L g198 ( .A(n_199), .Y(n_198) );
NAND2xp5_ASAP7_75t_L g199 ( .A(n_200), .B(n_211), .Y(n_199) );
NOR2xp33_ASAP7_75t_SL g267 ( .A(n_200), .B(n_268), .Y(n_267) );
NOR4xp25_ASAP7_75t_L g370 ( .A(n_200), .B(n_364), .C(n_368), .D(n_371), .Y(n_370) );
INVx1_ASAP7_75t_L g408 ( .A(n_200), .Y(n_408) );
AND2x2_ASAP7_75t_L g442 ( .A(n_200), .B(n_382), .Y(n_442) );
BUFx2_ASAP7_75t_L g200 ( .A(n_201), .Y(n_200) );
INVx2_ASAP7_75t_L g243 ( .A(n_201), .Y(n_243) );
INVx2_ASAP7_75t_L g201 ( .A(n_202), .Y(n_201) );
INVx2_ASAP7_75t_L g297 ( .A(n_202), .Y(n_297) );
OAI21x1_ASAP7_75t_SL g202 ( .A1(n_203), .A2(n_205), .B(n_209), .Y(n_202) );
INVx1_ASAP7_75t_L g210 ( .A(n_204), .Y(n_210) );
AOI33xp33_ASAP7_75t_L g438 ( .A1(n_211), .A2(n_240), .A3(n_271), .B1(n_287), .B2(n_393), .B3(n_439), .Y(n_438) );
INVx1_ASAP7_75t_SL g211 ( .A(n_212), .Y(n_211) );
AND2x2_ASAP7_75t_L g228 ( .A(n_212), .B(n_229), .Y(n_228) );
AND2x4_ASAP7_75t_L g238 ( .A(n_212), .B(n_239), .Y(n_238) );
BUFx3_ASAP7_75t_L g212 ( .A(n_213), .Y(n_212) );
INVx2_ASAP7_75t_L g245 ( .A(n_213), .Y(n_245) );
INVxp67_ASAP7_75t_L g326 ( .A(n_213), .Y(n_326) );
AND2x2_ASAP7_75t_L g382 ( .A(n_213), .B(n_247), .Y(n_382) );
AO21x2_ASAP7_75t_L g213 ( .A1(n_214), .A2(n_220), .B(n_221), .Y(n_213) );
AO21x2_ASAP7_75t_L g286 ( .A1(n_214), .A2(n_220), .B(n_221), .Y(n_286) );
NAND2xp5_ASAP7_75t_L g214 ( .A(n_215), .B(n_219), .Y(n_214) );
AO21x2_ASAP7_75t_L g247 ( .A1(n_220), .A2(n_248), .B(n_254), .Y(n_247) );
AO21x2_ASAP7_75t_L g283 ( .A1(n_220), .A2(n_248), .B(n_254), .Y(n_283) );
AO21x2_ASAP7_75t_L g567 ( .A1(n_220), .A2(n_568), .B(n_574), .Y(n_567) );
AO21x2_ASAP7_75t_L g605 ( .A1(n_220), .A2(n_568), .B(n_574), .Y(n_605) );
AOI21xp5_ASAP7_75t_L g403 ( .A1(n_222), .A2(n_404), .B(n_405), .Y(n_403) );
AND2x2_ASAP7_75t_L g222 ( .A(n_223), .B(n_224), .Y(n_222) );
AND2x2_ASAP7_75t_L g391 ( .A(n_223), .B(n_265), .Y(n_391) );
AND3x2_ASAP7_75t_L g393 ( .A(n_223), .B(n_277), .C(n_332), .Y(n_393) );
INVx3_ASAP7_75t_SL g345 ( .A(n_224), .Y(n_345) );
INVx4_ASAP7_75t_L g239 ( .A(n_225), .Y(n_239) );
AND2x2_ASAP7_75t_L g277 ( .A(n_225), .B(n_264), .Y(n_277) );
INVxp67_ASAP7_75t_L g226 ( .A(n_227), .Y(n_226) );
INVx1_ASAP7_75t_L g227 ( .A(n_228), .Y(n_227) );
BUFx2_ASAP7_75t_L g271 ( .A(n_229), .Y(n_271) );
AND2x4_ASAP7_75t_L g296 ( .A(n_229), .B(n_297), .Y(n_296) );
AND2x2_ASAP7_75t_L g359 ( .A(n_229), .B(n_247), .Y(n_359) );
INVx2_ASAP7_75t_L g229 ( .A(n_230), .Y(n_229) );
INVx2_ASAP7_75t_L g329 ( .A(n_230), .Y(n_329) );
HB1xp67_ASAP7_75t_L g351 ( .A(n_230), .Y(n_351) );
O2A1O1Ixp33_ASAP7_75t_R g236 ( .A1(n_237), .A2(n_240), .B(n_244), .C(n_255), .Y(n_236) );
CKINVDCx16_ASAP7_75t_R g237 ( .A(n_238), .Y(n_237) );
AND2x2_ASAP7_75t_L g288 ( .A(n_239), .B(n_289), .Y(n_288) );
NAND2xp5_ASAP7_75t_L g299 ( .A(n_239), .B(n_300), .Y(n_299) );
NAND2xp5_ASAP7_75t_L g417 ( .A(n_239), .B(n_256), .Y(n_417) );
INVx1_ASAP7_75t_SL g240 ( .A(n_241), .Y(n_240) );
AND2x2_ASAP7_75t_L g399 ( .A(n_241), .B(n_389), .Y(n_399) );
AND2x2_ASAP7_75t_SL g241 ( .A(n_242), .B(n_243), .Y(n_241) );
AND2x2_ASAP7_75t_L g246 ( .A(n_242), .B(n_247), .Y(n_246) );
AND2x2_ASAP7_75t_L g268 ( .A(n_242), .B(n_269), .Y(n_268) );
AND2x2_ASAP7_75t_L g284 ( .A(n_242), .B(n_285), .Y(n_284) );
AND2x4_ASAP7_75t_L g317 ( .A(n_242), .B(n_297), .Y(n_317) );
AND2x4_ASAP7_75t_L g282 ( .A(n_243), .B(n_283), .Y(n_282) );
OR2x2_ASAP7_75t_L g306 ( .A(n_243), .B(n_307), .Y(n_306) );
AND2x2_ASAP7_75t_L g344 ( .A(n_243), .B(n_269), .Y(n_344) );
NAND2xp5_ASAP7_75t_L g244 ( .A(n_245), .B(n_246), .Y(n_244) );
AND2x2_ASAP7_75t_L g272 ( .A(n_245), .B(n_269), .Y(n_272) );
AND2x2_ASAP7_75t_L g287 ( .A(n_245), .B(n_247), .Y(n_287) );
BUFx2_ASAP7_75t_L g343 ( .A(n_245), .Y(n_343) );
AND2x2_ASAP7_75t_L g357 ( .A(n_245), .B(n_268), .Y(n_357) );
INVx2_ASAP7_75t_L g269 ( .A(n_247), .Y(n_269) );
NAND2xp5_ASAP7_75t_SL g248 ( .A(n_249), .B(n_253), .Y(n_248) );
OAI22xp33_ASAP7_75t_L g305 ( .A1(n_255), .A2(n_306), .B1(n_308), .B2(n_312), .Y(n_305) );
INVx2_ASAP7_75t_SL g336 ( .A(n_255), .Y(n_336) );
OR2x2_ASAP7_75t_L g255 ( .A(n_256), .B(n_257), .Y(n_255) );
AND2x2_ASAP7_75t_L g311 ( .A(n_256), .B(n_264), .Y(n_311) );
INVx1_ASAP7_75t_L g418 ( .A(n_257), .Y(n_418) );
NOR3xp33_ASAP7_75t_L g258 ( .A(n_259), .B(n_291), .C(n_305), .Y(n_258) );
OAI221xp5_ASAP7_75t_SL g259 ( .A1(n_260), .A2(n_266), .B1(n_270), .B2(n_273), .C(n_275), .Y(n_259) );
INVx1_ASAP7_75t_SL g260 ( .A(n_261), .Y(n_260) );
AND2x2_ASAP7_75t_L g261 ( .A(n_262), .B(n_265), .Y(n_261) );
INVxp67_ASAP7_75t_SL g262 ( .A(n_263), .Y(n_262) );
INVx1_ASAP7_75t_L g319 ( .A(n_263), .Y(n_319) );
INVxp67_ASAP7_75t_SL g447 ( .A(n_263), .Y(n_447) );
INVx1_ASAP7_75t_L g410 ( .A(n_265), .Y(n_410) );
AND2x2_ASAP7_75t_SL g420 ( .A(n_265), .B(n_289), .Y(n_420) );
INVxp67_ASAP7_75t_L g266 ( .A(n_267), .Y(n_266) );
NAND2xp5_ASAP7_75t_L g325 ( .A(n_269), .B(n_297), .Y(n_325) );
NAND2xp5_ASAP7_75t_L g270 ( .A(n_271), .B(n_272), .Y(n_270) );
OR2x2_ASAP7_75t_L g303 ( .A(n_271), .B(n_304), .Y(n_303) );
INVx1_ASAP7_75t_L g381 ( .A(n_271), .Y(n_381) );
AND2x2_ASAP7_75t_L g316 ( .A(n_272), .B(n_317), .Y(n_316) );
INVx1_ASAP7_75t_L g273 ( .A(n_274), .Y(n_273) );
AND2x2_ASAP7_75t_L g362 ( .A(n_274), .B(n_322), .Y(n_362) );
AND2x2_ASAP7_75t_L g439 ( .A(n_274), .B(n_437), .Y(n_439) );
AOI22xp5_ASAP7_75t_L g275 ( .A1(n_276), .A2(n_280), .B1(n_287), .B2(n_288), .Y(n_275) );
AND2x4_ASAP7_75t_L g276 ( .A(n_277), .B(n_278), .Y(n_276) );
INVx2_ASAP7_75t_L g278 ( .A(n_279), .Y(n_278) );
OR2x2_ASAP7_75t_L g298 ( .A(n_279), .B(n_299), .Y(n_298) );
INVx1_ASAP7_75t_SL g280 ( .A(n_281), .Y(n_280) );
NAND2xp5_ASAP7_75t_L g281 ( .A(n_282), .B(n_284), .Y(n_281) );
INVx2_ASAP7_75t_L g304 ( .A(n_282), .Y(n_304) );
AND2x4_ASAP7_75t_L g328 ( .A(n_282), .B(n_329), .Y(n_328) );
OAI21xp33_ASAP7_75t_SL g358 ( .A1(n_282), .A2(n_359), .B(n_360), .Y(n_358) );
AND2x2_ASAP7_75t_L g385 ( .A(n_282), .B(n_343), .Y(n_385) );
INVx2_ASAP7_75t_L g307 ( .A(n_283), .Y(n_307) );
HB1xp67_ASAP7_75t_L g340 ( .A(n_283), .Y(n_340) );
INVx1_ASAP7_75t_SL g364 ( .A(n_284), .Y(n_364) );
INVx1_ASAP7_75t_L g285 ( .A(n_286), .Y(n_285) );
BUFx2_ASAP7_75t_L g295 ( .A(n_286), .Y(n_295) );
AND2x4_ASAP7_75t_SL g389 ( .A(n_286), .B(n_307), .Y(n_389) );
AND2x2_ASAP7_75t_L g386 ( .A(n_289), .B(n_332), .Y(n_386) );
AND2x2_ASAP7_75t_L g412 ( .A(n_289), .B(n_398), .Y(n_412) );
HB1xp67_ASAP7_75t_L g334 ( .A(n_290), .Y(n_334) );
INVx1_ASAP7_75t_L g354 ( .A(n_290), .Y(n_354) );
OAI22xp33_ASAP7_75t_L g291 ( .A1(n_292), .A2(n_298), .B1(n_301), .B2(n_303), .Y(n_291) );
INVx1_ASAP7_75t_L g292 ( .A(n_293), .Y(n_292) );
AND2x2_ASAP7_75t_L g293 ( .A(n_294), .B(n_296), .Y(n_293) );
INVx2_ASAP7_75t_L g294 ( .A(n_295), .Y(n_294) );
NAND2xp5_ASAP7_75t_SL g312 ( .A(n_296), .B(n_307), .Y(n_312) );
NAND2xp5_ASAP7_75t_L g388 ( .A(n_296), .B(n_389), .Y(n_388) );
INVx1_ASAP7_75t_L g435 ( .A(n_296), .Y(n_435) );
INVx2_ASAP7_75t_SL g360 ( .A(n_298), .Y(n_360) );
AND2x2_ASAP7_75t_L g372 ( .A(n_300), .B(n_332), .Y(n_372) );
INVx2_ASAP7_75t_L g378 ( .A(n_300), .Y(n_378) );
INVxp33_ASAP7_75t_L g301 ( .A(n_302), .Y(n_301) );
INVx2_ASAP7_75t_L g337 ( .A(n_303), .Y(n_337) );
NOR2xp33_ASAP7_75t_L g363 ( .A(n_306), .B(n_364), .Y(n_363) );
INVx1_ASAP7_75t_L g428 ( .A(n_306), .Y(n_428) );
INVx1_ASAP7_75t_L g356 ( .A(n_308), .Y(n_356) );
NAND2xp5_ASAP7_75t_L g308 ( .A(n_309), .B(n_311), .Y(n_308) );
NAND2xp5_ASAP7_75t_L g375 ( .A(n_309), .B(n_376), .Y(n_375) );
INVx2_ASAP7_75t_L g309 ( .A(n_310), .Y(n_309) );
AND2x2_ASAP7_75t_L g367 ( .A(n_311), .B(n_368), .Y(n_367) );
AOI22xp5_ASAP7_75t_L g440 ( .A1(n_311), .A2(n_441), .B1(n_442), .B2(n_443), .Y(n_440) );
NOR3xp33_ASAP7_75t_L g313 ( .A(n_314), .B(n_335), .C(n_338), .Y(n_313) );
OAI221xp5_ASAP7_75t_L g314 ( .A1(n_315), .A2(n_318), .B1(n_320), .B2(n_324), .C(n_327), .Y(n_314) );
INVx1_ASAP7_75t_SL g315 ( .A(n_316), .Y(n_315) );
INVx1_ASAP7_75t_SL g433 ( .A(n_318), .Y(n_433) );
INVx1_ASAP7_75t_L g318 ( .A(n_319), .Y(n_318) );
AND2x2_ASAP7_75t_L g402 ( .A(n_319), .B(n_368), .Y(n_402) );
OR2x2_ASAP7_75t_L g320 ( .A(n_321), .B(n_323), .Y(n_320) );
INVx1_ASAP7_75t_L g321 ( .A(n_322), .Y(n_321) );
AND2x2_ASAP7_75t_L g333 ( .A(n_322), .B(n_334), .Y(n_333) );
INVx1_ASAP7_75t_L g404 ( .A(n_324), .Y(n_404) );
OR2x2_ASAP7_75t_L g324 ( .A(n_325), .B(n_326), .Y(n_324) );
INVx1_ASAP7_75t_L g401 ( .A(n_325), .Y(n_401) );
INVx1_ASAP7_75t_L g407 ( .A(n_326), .Y(n_407) );
OR2x2_ASAP7_75t_L g430 ( .A(n_326), .B(n_431), .Y(n_430) );
NAND2xp5_ASAP7_75t_L g327 ( .A(n_328), .B(n_330), .Y(n_327) );
INVx1_ASAP7_75t_SL g339 ( .A(n_329), .Y(n_339) );
AND2x2_ASAP7_75t_L g409 ( .A(n_329), .B(n_389), .Y(n_409) );
AND2x2_ASAP7_75t_SL g441 ( .A(n_329), .B(n_342), .Y(n_441) );
INVx1_ASAP7_75t_SL g330 ( .A(n_331), .Y(n_330) );
NAND2xp5_ASAP7_75t_L g331 ( .A(n_332), .B(n_333), .Y(n_331) );
INVx1_ASAP7_75t_L g446 ( .A(n_332), .Y(n_446) );
INVx1_ASAP7_75t_L g396 ( .A(n_334), .Y(n_396) );
AND2x2_ASAP7_75t_L g335 ( .A(n_336), .B(n_337), .Y(n_335) );
O2A1O1Ixp33_ASAP7_75t_L g338 ( .A1(n_339), .A2(n_340), .B(n_341), .C(n_345), .Y(n_338) );
NAND2xp5_ASAP7_75t_L g413 ( .A(n_339), .B(n_389), .Y(n_413) );
INVx1_ASAP7_75t_L g341 ( .A(n_342), .Y(n_341) );
NAND2xp5_ASAP7_75t_L g392 ( .A(n_342), .B(n_393), .Y(n_392) );
AND2x2_ASAP7_75t_L g342 ( .A(n_343), .B(n_344), .Y(n_342) );
AND2x2_ASAP7_75t_L g350 ( .A(n_344), .B(n_351), .Y(n_350) );
INVx1_ASAP7_75t_L g431 ( .A(n_344), .Y(n_431) );
NAND4xp75_ASAP7_75t_L g346 ( .A(n_347), .B(n_403), .C(n_419), .D(n_440), .Y(n_346) );
NOR3x1_ASAP7_75t_L g347 ( .A(n_348), .B(n_365), .C(n_387), .Y(n_347) );
NAND4xp75_ASAP7_75t_L g348 ( .A(n_349), .B(n_355), .C(n_358), .D(n_361), .Y(n_348) );
NAND2xp5_ASAP7_75t_SL g349 ( .A(n_350), .B(n_352), .Y(n_349) );
AND2x2_ASAP7_75t_L g400 ( .A(n_351), .B(n_401), .Y(n_400) );
INVx1_ASAP7_75t_SL g425 ( .A(n_352), .Y(n_425) );
NAND2xp5_ASAP7_75t_SL g355 ( .A(n_356), .B(n_357), .Y(n_355) );
INVx1_ASAP7_75t_SL g414 ( .A(n_357), .Y(n_414) );
NAND2xp5_ASAP7_75t_L g361 ( .A(n_362), .B(n_363), .Y(n_361) );
NAND2xp5_ASAP7_75t_L g365 ( .A(n_366), .B(n_373), .Y(n_365) );
INVx2_ASAP7_75t_L g368 ( .A(n_369), .Y(n_368) );
NAND2xp5_ASAP7_75t_L g432 ( .A(n_369), .B(n_433), .Y(n_432) );
INVx1_ASAP7_75t_SL g371 ( .A(n_372), .Y(n_371) );
AOI21xp5_ASAP7_75t_L g373 ( .A1(n_374), .A2(n_379), .B(n_383), .Y(n_373) );
INVx1_ASAP7_75t_L g374 ( .A(n_375), .Y(n_374) );
INVx1_ASAP7_75t_L g376 ( .A(n_377), .Y(n_376) );
OAI322xp33_ASAP7_75t_L g405 ( .A1(n_377), .A2(n_406), .A3(n_410), .B1(n_411), .B2(n_413), .C1(n_414), .C2(n_415), .Y(n_405) );
INVx2_ASAP7_75t_L g377 ( .A(n_378), .Y(n_377) );
NAND2xp5_ASAP7_75t_L g423 ( .A(n_378), .B(n_424), .Y(n_423) );
INVx1_ASAP7_75t_L g379 ( .A(n_380), .Y(n_379) );
NAND2xp5_ASAP7_75t_L g380 ( .A(n_381), .B(n_382), .Y(n_380) );
NAND2xp5_ASAP7_75t_L g427 ( .A(n_381), .B(n_428), .Y(n_427) );
NAND2xp5_ASAP7_75t_L g434 ( .A(n_382), .B(n_435), .Y(n_434) );
INVx1_ASAP7_75t_L g383 ( .A(n_384), .Y(n_383) );
NAND2xp5_ASAP7_75t_L g384 ( .A(n_385), .B(n_386), .Y(n_384) );
OAI211xp5_ASAP7_75t_L g387 ( .A1(n_388), .A2(n_390), .B(n_392), .C(n_394), .Y(n_387) );
INVx1_ASAP7_75t_L g390 ( .A(n_391), .Y(n_390) );
AOI22xp5_ASAP7_75t_L g394 ( .A1(n_395), .A2(n_399), .B1(n_400), .B2(n_402), .Y(n_394) );
NOR2xp33_ASAP7_75t_SL g395 ( .A(n_396), .B(n_397), .Y(n_395) );
INVx2_ASAP7_75t_SL g397 ( .A(n_398), .Y(n_397) );
AOI21xp5_ASAP7_75t_L g406 ( .A1(n_407), .A2(n_408), .B(n_409), .Y(n_406) );
INVxp67_ASAP7_75t_L g411 ( .A(n_412), .Y(n_411) );
NOR2xp33_ASAP7_75t_L g444 ( .A(n_412), .B(n_445), .Y(n_444) );
NAND2xp5_ASAP7_75t_SL g415 ( .A(n_416), .B(n_418), .Y(n_415) );
INVx1_ASAP7_75t_L g416 ( .A(n_417), .Y(n_416) );
OR2x2_ASAP7_75t_L g422 ( .A(n_417), .B(n_423), .Y(n_422) );
O2A1O1Ixp5_ASAP7_75t_L g419 ( .A1(n_420), .A2(n_421), .B(n_426), .C(n_429), .Y(n_419) );
NAND2xp5_ASAP7_75t_SL g421 ( .A(n_422), .B(n_425), .Y(n_421) );
INVx1_ASAP7_75t_L g426 ( .A(n_427), .Y(n_426) );
OAI221xp5_ASAP7_75t_SL g429 ( .A1(n_430), .A2(n_432), .B1(n_434), .B2(n_436), .C(n_438), .Y(n_429) );
INVxp67_ASAP7_75t_L g436 ( .A(n_437), .Y(n_436) );
INVx1_ASAP7_75t_L g443 ( .A(n_444), .Y(n_443) );
AND2x2_ASAP7_75t_L g445 ( .A(n_446), .B(n_447), .Y(n_445) );
INVx2_ASAP7_75t_L g450 ( .A(n_451), .Y(n_450) );
BUFx2_ASAP7_75t_L g451 ( .A(n_452), .Y(n_451) );
BUFx2_ASAP7_75t_L g458 ( .A(n_452), .Y(n_458) );
NAND2xp5_ASAP7_75t_L g452 ( .A(n_453), .B(n_454), .Y(n_452) );
AND2x6_ASAP7_75t_SL g474 ( .A(n_453), .B(n_455), .Y(n_474) );
OR2x6_ASAP7_75t_SL g477 ( .A(n_453), .B(n_454), .Y(n_477) );
OR2x2_ASAP7_75t_L g816 ( .A(n_453), .B(n_455), .Y(n_816) );
CKINVDCx5p33_ASAP7_75t_R g454 ( .A(n_455), .Y(n_454) );
NAND2xp5_ASAP7_75t_SL g459 ( .A(n_456), .B(n_460), .Y(n_459) );
INVx1_ASAP7_75t_SL g457 ( .A(n_458), .Y(n_457) );
CKINVDCx11_ASAP7_75t_R g460 ( .A(n_461), .Y(n_460) );
CKINVDCx8_ASAP7_75t_R g461 ( .A(n_462), .Y(n_461) );
NAND2xp5_ASAP7_75t_SL g463 ( .A(n_464), .B(n_817), .Y(n_463) );
INVx1_ASAP7_75t_L g818 ( .A(n_465), .Y(n_818) );
CKINVDCx6p67_ASAP7_75t_R g471 ( .A(n_472), .Y(n_471) );
INVx4_ASAP7_75t_SL g821 ( .A(n_472), .Y(n_821) );
INVx3_ASAP7_75t_SL g472 ( .A(n_473), .Y(n_472) );
CKINVDCx5p33_ASAP7_75t_R g473 ( .A(n_474), .Y(n_473) );
INVx2_ASAP7_75t_L g475 ( .A(n_476), .Y(n_475) );
CKINVDCx11_ASAP7_75t_R g476 ( .A(n_477), .Y(n_476) );
OAI22x1_ASAP7_75t_L g819 ( .A1(n_477), .A2(n_820), .B1(n_821), .B2(n_822), .Y(n_819) );
INVx1_ASAP7_75t_L g822 ( .A(n_478), .Y(n_822) );
OR3x2_ASAP7_75t_L g478 ( .A(n_479), .B(n_680), .C(n_751), .Y(n_478) );
NAND3x1_ASAP7_75t_SL g479 ( .A(n_480), .B(n_607), .C(n_629), .Y(n_479) );
AND2x2_ASAP7_75t_L g480 ( .A(n_481), .B(n_597), .Y(n_480) );
AOI22xp33_ASAP7_75t_SL g481 ( .A1(n_482), .A2(n_528), .B1(n_575), .B2(n_579), .Y(n_481) );
AOI22xp33_ASAP7_75t_L g782 ( .A1(n_482), .A2(n_783), .B1(n_784), .B2(n_786), .Y(n_782) );
AND2x2_ASAP7_75t_L g482 ( .A(n_483), .B(n_503), .Y(n_482) );
AND2x2_ASAP7_75t_L g598 ( .A(n_483), .B(n_599), .Y(n_598) );
NAND2xp5_ASAP7_75t_SL g664 ( .A(n_483), .B(n_645), .Y(n_664) );
INVx1_ASAP7_75t_L g483 ( .A(n_484), .Y(n_483) );
INVx2_ASAP7_75t_L g582 ( .A(n_484), .Y(n_582) );
AND2x2_ASAP7_75t_L g632 ( .A(n_484), .B(n_505), .Y(n_632) );
INVx1_ASAP7_75t_L g671 ( .A(n_484), .Y(n_671) );
OR2x2_ASAP7_75t_L g708 ( .A(n_484), .B(n_520), .Y(n_708) );
HB1xp67_ASAP7_75t_L g720 ( .A(n_484), .Y(n_720) );
HB1xp67_ASAP7_75t_L g744 ( .A(n_484), .Y(n_744) );
AND2x2_ASAP7_75t_L g801 ( .A(n_484), .B(n_628), .Y(n_801) );
NAND2xp5_ASAP7_75t_L g485 ( .A(n_486), .B(n_492), .Y(n_485) );
INVx1_ASAP7_75t_L g552 ( .A(n_487), .Y(n_552) );
AND2x4_ASAP7_75t_L g487 ( .A(n_488), .B(n_491), .Y(n_487) );
INVx1_ASAP7_75t_L g588 ( .A(n_488), .Y(n_588) );
AND2x2_ASAP7_75t_L g488 ( .A(n_489), .B(n_490), .Y(n_488) );
OR2x6_ASAP7_75t_L g500 ( .A(n_489), .B(n_497), .Y(n_500) );
INVxp33_ASAP7_75t_L g562 ( .A(n_489), .Y(n_562) );
INVx1_ASAP7_75t_L g589 ( .A(n_491), .Y(n_589) );
INVxp67_ASAP7_75t_L g550 ( .A(n_493), .Y(n_550) );
NOR2x1p5_ASAP7_75t_L g494 ( .A(n_495), .B(n_496), .Y(n_494) );
INVx1_ASAP7_75t_L g563 ( .A(n_496), .Y(n_563) );
INVx3_ASAP7_75t_L g496 ( .A(n_497), .Y(n_496) );
OAI22xp5_ASAP7_75t_L g508 ( .A1(n_500), .A2(n_509), .B1(n_510), .B2(n_511), .Y(n_508) );
INVxp67_ASAP7_75t_L g541 ( .A(n_500), .Y(n_541) );
INVx2_ASAP7_75t_L g595 ( .A(n_500), .Y(n_595) );
NOR2x1_ASAP7_75t_L g503 ( .A(n_504), .B(n_518), .Y(n_503) );
INVx1_ASAP7_75t_L g676 ( .A(n_504), .Y(n_676) );
AND2x2_ASAP7_75t_L g702 ( .A(n_504), .B(n_520), .Y(n_702) );
NAND2x1_ASAP7_75t_L g718 ( .A(n_504), .B(n_719), .Y(n_718) );
INVx2_ASAP7_75t_L g504 ( .A(n_505), .Y(n_504) );
AND2x2_ASAP7_75t_L g599 ( .A(n_505), .B(n_585), .Y(n_599) );
INVx3_ASAP7_75t_L g628 ( .A(n_505), .Y(n_628) );
NOR2x1_ASAP7_75t_SL g747 ( .A(n_505), .B(n_520), .Y(n_747) );
AND2x4_ASAP7_75t_L g505 ( .A(n_506), .B(n_507), .Y(n_505) );
OAI21xp5_ASAP7_75t_L g507 ( .A1(n_508), .A2(n_512), .B(n_517), .Y(n_507) );
NOR2xp33_ASAP7_75t_L g542 ( .A(n_511), .B(n_543), .Y(n_542) );
OAI22xp5_ASAP7_75t_L g512 ( .A1(n_513), .A2(n_514), .B1(n_515), .B2(n_516), .Y(n_512) );
NOR2x1_ASAP7_75t_L g655 ( .A(n_518), .B(n_656), .Y(n_655) );
INVx1_ASAP7_75t_L g518 ( .A(n_519), .Y(n_518) );
AND2x2_ASAP7_75t_L g626 ( .A(n_519), .B(n_627), .Y(n_626) );
INVx2_ASAP7_75t_L g519 ( .A(n_520), .Y(n_519) );
INVx4_ASAP7_75t_L g596 ( .A(n_520), .Y(n_596) );
BUFx6f_ASAP7_75t_L g641 ( .A(n_520), .Y(n_641) );
AND2x2_ASAP7_75t_L g713 ( .A(n_520), .B(n_585), .Y(n_713) );
AND2x4_ASAP7_75t_L g730 ( .A(n_520), .B(n_674), .Y(n_730) );
NAND2xp5_ASAP7_75t_SL g777 ( .A(n_520), .B(n_672), .Y(n_777) );
NAND2xp5_ASAP7_75t_L g806 ( .A(n_520), .B(n_581), .Y(n_806) );
OR2x6_ASAP7_75t_L g520 ( .A(n_521), .B(n_522), .Y(n_520) );
AOI22xp5_ASAP7_75t_L g735 ( .A1(n_528), .A2(n_623), .B1(n_694), .B2(n_736), .Y(n_735) );
AND2x2_ASAP7_75t_L g528 ( .A(n_529), .B(n_553), .Y(n_528) );
INVx2_ASAP7_75t_L g696 ( .A(n_529), .Y(n_696) );
AND2x2_ASAP7_75t_L g529 ( .A(n_530), .B(n_537), .Y(n_529) );
BUFx3_ASAP7_75t_L g686 ( .A(n_530), .Y(n_686) );
INVx1_ASAP7_75t_L g530 ( .A(n_531), .Y(n_530) );
NAND2xp5_ASAP7_75t_L g578 ( .A(n_531), .B(n_555), .Y(n_578) );
INVx2_ASAP7_75t_L g602 ( .A(n_531), .Y(n_602) );
INVx1_ASAP7_75t_L g614 ( .A(n_531), .Y(n_614) );
AND2x4_ASAP7_75t_L g621 ( .A(n_531), .B(n_622), .Y(n_621) );
AND2x2_ASAP7_75t_L g638 ( .A(n_531), .B(n_538), .Y(n_638) );
HB1xp67_ASAP7_75t_L g652 ( .A(n_531), .Y(n_652) );
INVxp67_ASAP7_75t_L g660 ( .A(n_531), .Y(n_660) );
AND2x2_ASAP7_75t_L g689 ( .A(n_537), .B(n_605), .Y(n_689) );
AND2x2_ASAP7_75t_L g705 ( .A(n_537), .B(n_606), .Y(n_705) );
NOR2xp67_ASAP7_75t_L g792 ( .A(n_537), .B(n_605), .Y(n_792) );
INVx2_ASAP7_75t_L g537 ( .A(n_538), .Y(n_537) );
AND2x4_ASAP7_75t_L g601 ( .A(n_538), .B(n_602), .Y(n_601) );
INVx1_ASAP7_75t_L g612 ( .A(n_538), .Y(n_612) );
INVx1_ASAP7_75t_L g625 ( .A(n_538), .Y(n_625) );
NAND2xp5_ASAP7_75t_L g662 ( .A(n_538), .B(n_567), .Y(n_662) );
OR2x2_ASAP7_75t_L g538 ( .A(n_539), .B(n_546), .Y(n_538) );
OAI22xp5_ASAP7_75t_L g546 ( .A1(n_547), .A2(n_550), .B1(n_551), .B2(n_552), .Y(n_546) );
INVx1_ASAP7_75t_L g548 ( .A(n_549), .Y(n_548) );
INVx1_ASAP7_75t_L g785 ( .A(n_553), .Y(n_785) );
AND2x4_ASAP7_75t_L g553 ( .A(n_554), .B(n_566), .Y(n_553) );
AND2x2_ASAP7_75t_L g659 ( .A(n_554), .B(n_660), .Y(n_659) );
INVx1_ASAP7_75t_L g688 ( .A(n_554), .Y(n_688) );
AND2x2_ASAP7_75t_L g790 ( .A(n_554), .B(n_605), .Y(n_790) );
INVx2_ASAP7_75t_L g554 ( .A(n_555), .Y(n_554) );
NAND2xp5_ASAP7_75t_L g650 ( .A(n_555), .B(n_567), .Y(n_650) );
AO21x2_ASAP7_75t_L g555 ( .A1(n_556), .A2(n_557), .B(n_565), .Y(n_555) );
AO21x2_ASAP7_75t_L g606 ( .A1(n_556), .A2(n_557), .B(n_565), .Y(n_606) );
NAND2xp5_ASAP7_75t_SL g557 ( .A(n_558), .B(n_564), .Y(n_557) );
INVx1_ASAP7_75t_L g560 ( .A(n_561), .Y(n_560) );
INVx3_ASAP7_75t_L g576 ( .A(n_566), .Y(n_576) );
NAND2x1p5_ASAP7_75t_L g765 ( .A(n_566), .B(n_686), .Y(n_765) );
INVx3_ASAP7_75t_L g566 ( .A(n_567), .Y(n_566) );
HB1xp67_ASAP7_75t_L g679 ( .A(n_567), .Y(n_679) );
AND2x2_ASAP7_75t_L g706 ( .A(n_567), .B(n_652), .Y(n_706) );
NAND2xp5_ASAP7_75t_L g568 ( .A(n_569), .B(n_570), .Y(n_568) );
AND2x2_ASAP7_75t_L g575 ( .A(n_576), .B(n_577), .Y(n_575) );
AND2x2_ASAP7_75t_L g620 ( .A(n_576), .B(n_621), .Y(n_620) );
INVx1_ASAP7_75t_L g636 ( .A(n_576), .Y(n_636) );
AND2x2_ASAP7_75t_L g724 ( .A(n_576), .B(n_601), .Y(n_724) );
NAND2xp5_ASAP7_75t_L g749 ( .A(n_576), .B(n_744), .Y(n_749) );
AND2x2_ASAP7_75t_L g759 ( .A(n_576), .B(n_638), .Y(n_759) );
OR2x2_ASAP7_75t_L g796 ( .A(n_576), .B(n_696), .Y(n_796) );
NAND2xp5_ASAP7_75t_L g635 ( .A(n_577), .B(n_636), .Y(n_635) );
AND2x2_ASAP7_75t_L g756 ( .A(n_577), .B(n_612), .Y(n_756) );
AND2x2_ASAP7_75t_L g772 ( .A(n_577), .B(n_773), .Y(n_772) );
INVx2_ASAP7_75t_L g577 ( .A(n_578), .Y(n_577) );
OR2x2_ASAP7_75t_L g766 ( .A(n_578), .B(n_662), .Y(n_766) );
AND2x2_ASAP7_75t_L g579 ( .A(n_580), .B(n_583), .Y(n_579) );
INVx1_ASAP7_75t_L g648 ( .A(n_580), .Y(n_648) );
NAND2xp5_ASAP7_75t_L g729 ( .A(n_580), .B(n_730), .Y(n_729) );
AND2x2_ASAP7_75t_L g746 ( .A(n_580), .B(n_747), .Y(n_746) );
NAND2xp5_ASAP7_75t_L g771 ( .A(n_580), .B(n_627), .Y(n_771) );
INVx3_ASAP7_75t_L g580 ( .A(n_581), .Y(n_580) );
HB1xp67_ASAP7_75t_L g618 ( .A(n_581), .Y(n_618) );
INVx2_ASAP7_75t_L g581 ( .A(n_582), .Y(n_581) );
HB1xp67_ASAP7_75t_L g727 ( .A(n_582), .Y(n_727) );
AOI22xp5_ASAP7_75t_L g633 ( .A1(n_583), .A2(n_616), .B1(n_634), .B2(n_637), .Y(n_633) );
NOR2xp33_ASAP7_75t_L g717 ( .A(n_583), .B(n_718), .Y(n_717) );
INVx2_ASAP7_75t_SL g750 ( .A(n_583), .Y(n_750) );
AND2x4_ASAP7_75t_SL g583 ( .A(n_584), .B(n_596), .Y(n_583) );
HB1xp67_ASAP7_75t_L g584 ( .A(n_585), .Y(n_584) );
AND2x4_ASAP7_75t_L g627 ( .A(n_585), .B(n_628), .Y(n_627) );
INVx2_ASAP7_75t_L g647 ( .A(n_585), .Y(n_647) );
INVx1_ASAP7_75t_L g674 ( .A(n_585), .Y(n_674) );
AND2x2_ASAP7_75t_L g585 ( .A(n_586), .B(n_591), .Y(n_585) );
NOR3xp33_ASAP7_75t_L g587 ( .A(n_588), .B(n_589), .C(n_590), .Y(n_587) );
HB1xp67_ASAP7_75t_L g616 ( .A(n_596), .Y(n_616) );
AND2x4_ASAP7_75t_L g673 ( .A(n_596), .B(n_674), .Y(n_673) );
NOR2x1_ASAP7_75t_L g734 ( .A(n_596), .B(n_703), .Y(n_734) );
NAND2xp5_ASAP7_75t_L g597 ( .A(n_598), .B(n_600), .Y(n_597) );
AND2x2_ASAP7_75t_L g698 ( .A(n_598), .B(n_641), .Y(n_698) );
OAI21xp5_ASAP7_75t_L g778 ( .A1(n_598), .A2(n_779), .B(n_780), .Y(n_778) );
INVx2_ASAP7_75t_L g656 ( .A(n_599), .Y(n_656) );
AOI22xp5_ASAP7_75t_L g709 ( .A1(n_600), .A2(n_710), .B1(n_714), .B2(n_717), .Y(n_709) );
AND2x2_ASAP7_75t_L g600 ( .A(n_601), .B(n_603), .Y(n_600) );
HB1xp67_ASAP7_75t_L g667 ( .A(n_601), .Y(n_667) );
AND2x2_ASAP7_75t_L g677 ( .A(n_601), .B(n_678), .Y(n_677) );
INVx3_ASAP7_75t_L g716 ( .A(n_601), .Y(n_716) );
NAND2x1_ASAP7_75t_SL g741 ( .A(n_601), .B(n_610), .Y(n_741) );
AND2x2_ASAP7_75t_L g637 ( .A(n_603), .B(n_638), .Y(n_637) );
AND2x4_ASAP7_75t_L g603 ( .A(n_604), .B(n_606), .Y(n_603) );
INVx2_ASAP7_75t_L g604 ( .A(n_605), .Y(n_604) );
NOR2x1_ASAP7_75t_L g613 ( .A(n_605), .B(n_614), .Y(n_613) );
INVx1_ASAP7_75t_L g610 ( .A(n_606), .Y(n_610) );
INVx2_ASAP7_75t_L g622 ( .A(n_606), .Y(n_622) );
AOI21xp5_ASAP7_75t_SL g607 ( .A1(n_608), .A2(n_615), .B(n_619), .Y(n_607) );
INVx1_ASAP7_75t_L g608 ( .A(n_609), .Y(n_608) );
NAND2xp5_ASAP7_75t_L g609 ( .A(n_610), .B(n_611), .Y(n_609) );
NAND2xp5_ASAP7_75t_L g803 ( .A(n_610), .B(n_804), .Y(n_803) );
AOI22xp5_ASAP7_75t_L g699 ( .A1(n_611), .A2(n_700), .B1(n_704), .B2(n_707), .Y(n_699) );
AND2x2_ASAP7_75t_L g611 ( .A(n_612), .B(n_613), .Y(n_611) );
BUFx2_ASAP7_75t_L g804 ( .A(n_612), .Y(n_804) );
INVx1_ASAP7_75t_SL g811 ( .A(n_612), .Y(n_811) );
HB1xp67_ASAP7_75t_L g774 ( .A(n_613), .Y(n_774) );
NOR2xp33_ASAP7_75t_L g615 ( .A(n_616), .B(n_617), .Y(n_615) );
HB1xp67_ASAP7_75t_L g617 ( .A(n_618), .Y(n_617) );
OA21x2_ASAP7_75t_L g619 ( .A1(n_620), .A2(n_623), .B(n_626), .Y(n_619) );
AND2x2_ASAP7_75t_L g623 ( .A(n_621), .B(n_624), .Y(n_623) );
AND2x2_ASAP7_75t_L g665 ( .A(n_621), .B(n_661), .Y(n_665) );
AND2x2_ASAP7_75t_L g780 ( .A(n_621), .B(n_678), .Y(n_780) );
AND2x2_ASAP7_75t_L g783 ( .A(n_621), .B(n_689), .Y(n_783) );
AND2x4_ASAP7_75t_L g791 ( .A(n_621), .B(n_792), .Y(n_791) );
OAI21xp33_ASAP7_75t_L g745 ( .A1(n_623), .A2(n_746), .B(n_748), .Y(n_745) );
INVx2_ASAP7_75t_L g624 ( .A(n_625), .Y(n_624) );
INVx1_ASAP7_75t_L g773 ( .A(n_625), .Y(n_773) );
AND2x2_ASAP7_75t_L g789 ( .A(n_625), .B(n_790), .Y(n_789) );
INVx4_ASAP7_75t_L g703 ( .A(n_627), .Y(n_703) );
INVx1_ASAP7_75t_L g672 ( .A(n_628), .Y(n_672) );
AND2x2_ASAP7_75t_L g694 ( .A(n_628), .B(n_647), .Y(n_694) );
NOR2x1_ASAP7_75t_L g629 ( .A(n_630), .B(n_653), .Y(n_629) );
OAI21xp5_ASAP7_75t_L g630 ( .A1(n_631), .A2(n_633), .B(n_639), .Y(n_630) );
INVx1_ASAP7_75t_L g631 ( .A(n_632), .Y(n_631) );
AND2x2_ASAP7_75t_L g640 ( .A(n_632), .B(n_641), .Y(n_640) );
AND2x2_ASAP7_75t_SL g793 ( .A(n_632), .B(n_645), .Y(n_793) );
AND2x2_ASAP7_75t_L g814 ( .A(n_632), .B(n_730), .Y(n_814) );
INVx1_ASAP7_75t_L g634 ( .A(n_635), .Y(n_634) );
INVx2_ASAP7_75t_L g740 ( .A(n_637), .Y(n_740) );
OAI21xp5_ASAP7_75t_SL g639 ( .A1(n_640), .A2(n_642), .B(n_649), .Y(n_639) );
OR2x6_ASAP7_75t_L g692 ( .A(n_641), .B(n_693), .Y(n_692) );
INVx1_ASAP7_75t_L g642 ( .A(n_643), .Y(n_642) );
NAND2xp5_ASAP7_75t_L g643 ( .A(n_644), .B(n_648), .Y(n_643) );
INVx2_ASAP7_75t_SL g644 ( .A(n_645), .Y(n_644) );
INVx2_ASAP7_75t_L g645 ( .A(n_646), .Y(n_645) );
INVx1_ASAP7_75t_L g646 ( .A(n_647), .Y(n_646) );
NOR2xp33_ASAP7_75t_L g649 ( .A(n_650), .B(n_651), .Y(n_649) );
OR2x2_ASAP7_75t_L g715 ( .A(n_650), .B(n_716), .Y(n_715) );
INVx1_ASAP7_75t_L g812 ( .A(n_650), .Y(n_812) );
NOR2xp33_ASAP7_75t_L g784 ( .A(n_651), .B(n_785), .Y(n_784) );
HB1xp67_ASAP7_75t_L g651 ( .A(n_652), .Y(n_651) );
NAND2xp5_ASAP7_75t_L g653 ( .A(n_654), .B(n_666), .Y(n_653) );
AOI22xp5_ASAP7_75t_L g654 ( .A1(n_655), .A2(n_657), .B1(n_663), .B2(n_665), .Y(n_654) );
OR2x2_ASAP7_75t_L g726 ( .A(n_656), .B(n_727), .Y(n_726) );
INVx3_ASAP7_75t_L g657 ( .A(n_658), .Y(n_657) );
HB1xp67_ASAP7_75t_L g683 ( .A(n_658), .Y(n_683) );
NAND2x1p5_ASAP7_75t_L g658 ( .A(n_659), .B(n_661), .Y(n_658) );
INVx1_ASAP7_75t_L g732 ( .A(n_661), .Y(n_732) );
INVx2_ASAP7_75t_SL g661 ( .A(n_662), .Y(n_661) );
INVxp67_ASAP7_75t_L g663 ( .A(n_664), .Y(n_663) );
AOI22xp5_ASAP7_75t_L g666 ( .A1(n_667), .A2(n_668), .B1(n_675), .B2(n_677), .Y(n_666) );
INVx1_ASAP7_75t_L g668 ( .A(n_669), .Y(n_668) );
NAND2xp5_ASAP7_75t_L g669 ( .A(n_670), .B(n_673), .Y(n_669) );
AND2x4_ASAP7_75t_SL g670 ( .A(n_671), .B(n_672), .Y(n_670) );
AND2x2_ASAP7_75t_L g675 ( .A(n_673), .B(n_676), .Y(n_675) );
AND2x2_ASAP7_75t_L g736 ( .A(n_676), .B(n_730), .Y(n_736) );
INVx1_ASAP7_75t_L g678 ( .A(n_679), .Y(n_678) );
NAND2xp5_ASAP7_75t_SL g680 ( .A(n_681), .B(n_721), .Y(n_680) );
NOR2xp67_ASAP7_75t_L g681 ( .A(n_682), .B(n_695), .Y(n_681) );
AOI21xp33_ASAP7_75t_SL g682 ( .A1(n_683), .A2(n_684), .B(n_690), .Y(n_682) );
OR2x2_ASAP7_75t_L g684 ( .A(n_685), .B(n_687), .Y(n_684) );
INVx3_ASAP7_75t_L g685 ( .A(n_686), .Y(n_685) );
NAND2x1p5_ASAP7_75t_L g687 ( .A(n_688), .B(n_689), .Y(n_687) );
INVx1_ASAP7_75t_L g690 ( .A(n_691), .Y(n_690) );
INVx2_ASAP7_75t_L g691 ( .A(n_692), .Y(n_691) );
OAI22xp33_ASAP7_75t_SL g760 ( .A1(n_692), .A2(n_761), .B1(n_763), .B2(n_766), .Y(n_760) );
NOR2x1_ASAP7_75t_L g707 ( .A(n_693), .B(n_708), .Y(n_707) );
INVx2_ASAP7_75t_L g693 ( .A(n_694), .Y(n_693) );
AND2x2_ASAP7_75t_L g743 ( .A(n_694), .B(n_744), .Y(n_743) );
OAI211xp5_ASAP7_75t_L g695 ( .A1(n_696), .A2(n_697), .B(n_699), .C(n_709), .Y(n_695) );
INVx2_ASAP7_75t_L g697 ( .A(n_698), .Y(n_697) );
NAND2xp33_ASAP7_75t_SL g700 ( .A(n_701), .B(n_703), .Y(n_700) );
INVxp33_ASAP7_75t_L g701 ( .A(n_702), .Y(n_701) );
INVx2_ASAP7_75t_L g712 ( .A(n_703), .Y(n_712) );
AOI221xp5_ASAP7_75t_L g723 ( .A1(n_704), .A2(n_724), .B1(n_725), .B2(n_728), .C(n_731), .Y(n_723) );
AND2x4_ASAP7_75t_L g704 ( .A(n_705), .B(n_706), .Y(n_704) );
INVx1_ASAP7_75t_L g764 ( .A(n_705), .Y(n_764) );
INVx2_ASAP7_75t_SL g762 ( .A(n_708), .Y(n_762) );
INVx1_ASAP7_75t_L g710 ( .A(n_711), .Y(n_710) );
NOR2xp33_ASAP7_75t_L g711 ( .A(n_712), .B(n_713), .Y(n_711) );
NAND2x1_ASAP7_75t_L g761 ( .A(n_712), .B(n_762), .Y(n_761) );
INVx1_ASAP7_75t_L g714 ( .A(n_715), .Y(n_714) );
INVx1_ASAP7_75t_L g758 ( .A(n_718), .Y(n_758) );
INVx1_ASAP7_75t_L g787 ( .A(n_719), .Y(n_787) );
INVx1_ASAP7_75t_L g719 ( .A(n_720), .Y(n_719) );
NOR2x1_ASAP7_75t_L g721 ( .A(n_722), .B(n_737), .Y(n_721) );
NAND2xp5_ASAP7_75t_L g722 ( .A(n_723), .B(n_735), .Y(n_722) );
INVx1_ASAP7_75t_L g725 ( .A(n_726), .Y(n_725) );
INVx1_ASAP7_75t_L g776 ( .A(n_727), .Y(n_776) );
INVx1_ASAP7_75t_L g728 ( .A(n_729), .Y(n_728) );
AND2x2_ASAP7_75t_L g797 ( .A(n_730), .B(n_798), .Y(n_797) );
INVx2_ASAP7_75t_L g802 ( .A(n_730), .Y(n_802) );
NOR2xp33_ASAP7_75t_L g731 ( .A(n_732), .B(n_733), .Y(n_731) );
INVxp33_ASAP7_75t_L g733 ( .A(n_734), .Y(n_733) );
BUFx2_ASAP7_75t_L g755 ( .A(n_734), .Y(n_755) );
OAI21xp5_ASAP7_75t_SL g737 ( .A1(n_738), .A2(n_742), .B(n_745), .Y(n_737) );
INVxp67_ASAP7_75t_L g738 ( .A(n_739), .Y(n_738) );
NAND2xp5_ASAP7_75t_L g739 ( .A(n_740), .B(n_741), .Y(n_739) );
INVx2_ASAP7_75t_L g742 ( .A(n_743), .Y(n_742) );
BUFx2_ASAP7_75t_L g798 ( .A(n_744), .Y(n_798) );
AND2x2_ASAP7_75t_L g786 ( .A(n_747), .B(n_787), .Y(n_786) );
NOR2xp33_ASAP7_75t_R g748 ( .A(n_749), .B(n_750), .Y(n_748) );
NAND3xp33_ASAP7_75t_L g751 ( .A(n_752), .B(n_767), .C(n_794), .Y(n_751) );
NOR2xp33_ASAP7_75t_L g752 ( .A(n_753), .B(n_760), .Y(n_752) );
NAND2xp5_ASAP7_75t_SL g753 ( .A(n_754), .B(n_757), .Y(n_753) );
NAND2xp5_ASAP7_75t_L g754 ( .A(n_755), .B(n_756), .Y(n_754) );
NAND2xp5_ASAP7_75t_L g757 ( .A(n_758), .B(n_759), .Y(n_757) );
OR2x2_ASAP7_75t_L g763 ( .A(n_764), .B(n_765), .Y(n_763) );
NOR2xp33_ASAP7_75t_L g767 ( .A(n_768), .B(n_781), .Y(n_767) );
NAND2xp5_ASAP7_75t_SL g768 ( .A(n_769), .B(n_778), .Y(n_768) );
AOI22xp33_ASAP7_75t_SL g769 ( .A1(n_770), .A2(n_772), .B1(n_774), .B2(n_775), .Y(n_769) );
INVx1_ASAP7_75t_L g770 ( .A(n_771), .Y(n_770) );
NOR2x1_ASAP7_75t_L g775 ( .A(n_776), .B(n_777), .Y(n_775) );
INVxp67_ASAP7_75t_SL g779 ( .A(n_777), .Y(n_779) );
NAND2xp5_ASAP7_75t_SL g781 ( .A(n_782), .B(n_788), .Y(n_781) );
OAI21xp5_ASAP7_75t_L g788 ( .A1(n_789), .A2(n_791), .B(n_793), .Y(n_788) );
INVx1_ASAP7_75t_L g807 ( .A(n_791), .Y(n_807) );
AOI211xp5_ASAP7_75t_L g794 ( .A1(n_795), .A2(n_797), .B(n_799), .C(n_808), .Y(n_794) );
INVx1_ASAP7_75t_L g795 ( .A(n_796), .Y(n_795) );
OAI22xp5_ASAP7_75t_L g799 ( .A1(n_800), .A2(n_803), .B1(n_805), .B2(n_807), .Y(n_799) );
NAND2xp5_ASAP7_75t_L g800 ( .A(n_801), .B(n_802), .Y(n_800) );
HB1xp67_ASAP7_75t_L g805 ( .A(n_806), .Y(n_805) );
NOR2xp33_ASAP7_75t_L g808 ( .A(n_809), .B(n_813), .Y(n_808) );
INVx1_ASAP7_75t_L g809 ( .A(n_810), .Y(n_809) );
AND2x2_ASAP7_75t_L g810 ( .A(n_811), .B(n_812), .Y(n_810) );
INVxp67_ASAP7_75t_L g813 ( .A(n_814), .Y(n_813) );
INVx2_ASAP7_75t_L g815 ( .A(n_816), .Y(n_815) );
NAND2xp5_ASAP7_75t_L g817 ( .A(n_818), .B(n_819), .Y(n_817) );
NOR2xp33_ASAP7_75t_L g823 ( .A(n_824), .B(n_825), .Y(n_823) );
endmodule