module fake_jpeg_19747_n_86 (n_13, n_21, n_1, n_10, n_6, n_14, n_19, n_18, n_20, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_86);

input n_13;
input n_21;
input n_1;
input n_10;
input n_6;
input n_14;
input n_19;
input n_18;
input n_20;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_86;

wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_73;
wire n_59;
wire n_84;
wire n_65;
wire n_42;
wire n_49;
wire n_76;
wire n_28;
wire n_38;
wire n_26;
wire n_74;
wire n_31;
wire n_29;
wire n_50;
wire n_57;
wire n_23;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_30;
wire n_24;
wire n_44;
wire n_25;
wire n_75;
wire n_37;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_68;
wire n_52;
wire n_58;
wire n_41;
wire n_60;
wire n_63;
wire n_34;
wire n_39;
wire n_72;
wire n_56;
wire n_79;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_22;
wire n_48;
wire n_35;
wire n_46;
wire n_36;
wire n_62;
wire n_43;
wire n_32;
wire n_82;

AND2x2_ASAP7_75t_L g22 ( 
.A(n_12),
.B(n_7),
.Y(n_22)
);

INVx2_ASAP7_75t_L g23 ( 
.A(n_7),
.Y(n_23)
);

INVx2_ASAP7_75t_L g24 ( 
.A(n_14),
.Y(n_24)
);

NOR2xp33_ASAP7_75t_L g25 ( 
.A(n_16),
.B(n_4),
.Y(n_25)
);

INVx4_ASAP7_75t_L g26 ( 
.A(n_19),
.Y(n_26)
);

INVx5_ASAP7_75t_L g27 ( 
.A(n_4),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_11),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_18),
.Y(n_29)
);

BUFx12f_ASAP7_75t_L g30 ( 
.A(n_15),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_21),
.Y(n_31)
);

INVx2_ASAP7_75t_L g32 ( 
.A(n_2),
.Y(n_32)
);

BUFx8_ASAP7_75t_L g33 ( 
.A(n_0),
.Y(n_33)
);

BUFx2_ASAP7_75t_L g34 ( 
.A(n_6),
.Y(n_34)
);

BUFx3_ASAP7_75t_L g35 ( 
.A(n_1),
.Y(n_35)
);

INVx3_ASAP7_75t_L g36 ( 
.A(n_2),
.Y(n_36)
);

INVx6_ASAP7_75t_L g37 ( 
.A(n_13),
.Y(n_37)
);

AOI22xp33_ASAP7_75t_L g38 ( 
.A1(n_17),
.A2(n_3),
.B1(n_10),
.B2(n_6),
.Y(n_38)
);

INVx4_ASAP7_75t_L g39 ( 
.A(n_3),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_1),
.Y(n_40)
);

BUFx2_ASAP7_75t_L g41 ( 
.A(n_9),
.Y(n_41)
);

BUFx4f_ASAP7_75t_L g42 ( 
.A(n_8),
.Y(n_42)
);

OAI22xp5_ASAP7_75t_L g43 ( 
.A1(n_37),
.A2(n_20),
.B1(n_5),
.B2(n_8),
.Y(n_43)
);

OAI22xp5_ASAP7_75t_L g64 ( 
.A1(n_43),
.A2(n_47),
.B1(n_51),
.B2(n_52),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_24),
.Y(n_44)
);

INVx6_ASAP7_75t_L g65 ( 
.A(n_44),
.Y(n_65)
);

HB1xp67_ASAP7_75t_L g45 ( 
.A(n_33),
.Y(n_45)
);

INVx13_ASAP7_75t_L g60 ( 
.A(n_45),
.Y(n_60)
);

BUFx12f_ASAP7_75t_L g46 ( 
.A(n_30),
.Y(n_46)
);

INVx13_ASAP7_75t_L g61 ( 
.A(n_46),
.Y(n_61)
);

AOI22xp33_ASAP7_75t_L g47 ( 
.A1(n_23),
.A2(n_0),
.B1(n_5),
.B2(n_32),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_40),
.B(n_22),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_48),
.B(n_49),
.Y(n_62)
);

INVx3_ASAP7_75t_L g49 ( 
.A(n_42),
.Y(n_49)
);

INVx2_ASAP7_75t_L g50 ( 
.A(n_33),
.Y(n_50)
);

AND2x2_ASAP7_75t_L g66 ( 
.A(n_50),
.B(n_53),
.Y(n_66)
);

AOI22xp33_ASAP7_75t_SL g51 ( 
.A1(n_24),
.A2(n_23),
.B1(n_32),
.B2(n_26),
.Y(n_51)
);

AOI22xp33_ASAP7_75t_SL g52 ( 
.A1(n_39),
.A2(n_27),
.B1(n_36),
.B2(n_38),
.Y(n_52)
);

AND2x2_ASAP7_75t_L g53 ( 
.A(n_30),
.B(n_25),
.Y(n_53)
);

INVx4_ASAP7_75t_L g54 ( 
.A(n_35),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_L g67 ( 
.A(n_54),
.B(n_55),
.Y(n_67)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_28),
.Y(n_55)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_34),
.Y(n_56)
);

MAJIxp5_ASAP7_75t_L g63 ( 
.A(n_56),
.B(n_57),
.C(n_58),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g57 ( 
.A(n_31),
.B(n_29),
.Y(n_57)
);

INVx4_ASAP7_75t_L g58 ( 
.A(n_41),
.Y(n_58)
);

CKINVDCx12_ASAP7_75t_R g59 ( 
.A(n_41),
.Y(n_59)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_67),
.Y(n_68)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_68),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_SL g69 ( 
.A(n_67),
.B(n_53),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_L g73 ( 
.A(n_69),
.B(n_70),
.Y(n_73)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_60),
.Y(n_70)
);

OAI22xp5_ASAP7_75t_SL g71 ( 
.A1(n_64),
.A2(n_52),
.B1(n_51),
.B2(n_47),
.Y(n_71)
);

AOI21xp5_ASAP7_75t_L g74 ( 
.A1(n_71),
.A2(n_72),
.B(n_66),
.Y(n_74)
);

MAJIxp5_ASAP7_75t_L g72 ( 
.A(n_66),
.B(n_46),
.C(n_59),
.Y(n_72)
);

OAI22xp5_ASAP7_75t_L g78 ( 
.A1(n_74),
.A2(n_75),
.B1(n_63),
.B2(n_62),
.Y(n_78)
);

NOR2xp67_ASAP7_75t_L g75 ( 
.A(n_72),
.B(n_66),
.Y(n_75)
);

HB1xp67_ASAP7_75t_L g77 ( 
.A(n_73),
.Y(n_77)
);

INVxp67_ASAP7_75t_L g79 ( 
.A(n_77),
.Y(n_79)
);

XOR2xp5_ASAP7_75t_L g80 ( 
.A(n_78),
.B(n_74),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_SL g81 ( 
.A(n_80),
.B(n_79),
.Y(n_81)
);

XOR2xp5_ASAP7_75t_L g84 ( 
.A(n_81),
.B(n_61),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_SL g82 ( 
.A(n_80),
.B(n_76),
.Y(n_82)
);

AOI311xp33_ASAP7_75t_L g83 ( 
.A1(n_82),
.A2(n_71),
.A3(n_63),
.B(n_65),
.C(n_45),
.Y(n_83)
);

AOI21xp33_ASAP7_75t_L g85 ( 
.A1(n_83),
.A2(n_84),
.B(n_61),
.Y(n_85)
);

XOR2xp5_ASAP7_75t_L g86 ( 
.A(n_85),
.B(n_60),
.Y(n_86)
);


endmodule