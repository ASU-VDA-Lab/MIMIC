module fake_ariane_3298_n_1869 (n_83, n_8, n_56, n_60, n_160, n_64, n_119, n_124, n_167, n_90, n_38, n_47, n_110, n_153, n_18, n_86, n_75, n_89, n_67, n_149, n_34, n_158, n_69, n_95, n_92, n_143, n_150, n_98, n_74, n_113, n_114, n_33, n_19, n_40, n_152, n_120, n_106, n_12, n_53, n_111, n_21, n_115, n_133, n_66, n_71, n_24, n_7, n_109, n_96, n_156, n_49, n_20, n_100, n_17, n_50, n_132, n_62, n_147, n_51, n_166, n_76, n_103, n_79, n_26, n_3, n_46, n_0, n_84, n_36, n_91, n_159, n_107, n_72, n_105, n_128, n_44, n_30, n_82, n_31, n_42, n_57, n_131, n_70, n_10, n_117, n_139, n_165, n_85, n_130, n_144, n_6, n_48, n_94, n_101, n_4, n_134, n_2, n_32, n_37, n_58, n_65, n_123, n_9, n_138, n_112, n_45, n_162, n_11, n_129, n_126, n_137, n_122, n_148, n_164, n_52, n_157, n_135, n_73, n_77, n_15, n_118, n_93, n_121, n_23, n_61, n_108, n_102, n_125, n_22, n_168, n_43, n_1, n_81, n_87, n_13, n_27, n_29, n_41, n_140, n_55, n_151, n_136, n_28, n_80, n_146, n_97, n_154, n_142, n_161, n_14, n_163, n_88, n_141, n_68, n_116, n_104, n_145, n_78, n_39, n_59, n_63, n_99, n_16, n_5, n_155, n_127, n_35, n_54, n_25, n_1869);

input n_83;
input n_8;
input n_56;
input n_60;
input n_160;
input n_64;
input n_119;
input n_124;
input n_167;
input n_90;
input n_38;
input n_47;
input n_110;
input n_153;
input n_18;
input n_86;
input n_75;
input n_89;
input n_67;
input n_149;
input n_34;
input n_158;
input n_69;
input n_95;
input n_92;
input n_143;
input n_150;
input n_98;
input n_74;
input n_113;
input n_114;
input n_33;
input n_19;
input n_40;
input n_152;
input n_120;
input n_106;
input n_12;
input n_53;
input n_111;
input n_21;
input n_115;
input n_133;
input n_66;
input n_71;
input n_24;
input n_7;
input n_109;
input n_96;
input n_156;
input n_49;
input n_20;
input n_100;
input n_17;
input n_50;
input n_132;
input n_62;
input n_147;
input n_51;
input n_166;
input n_76;
input n_103;
input n_79;
input n_26;
input n_3;
input n_46;
input n_0;
input n_84;
input n_36;
input n_91;
input n_159;
input n_107;
input n_72;
input n_105;
input n_128;
input n_44;
input n_30;
input n_82;
input n_31;
input n_42;
input n_57;
input n_131;
input n_70;
input n_10;
input n_117;
input n_139;
input n_165;
input n_85;
input n_130;
input n_144;
input n_6;
input n_48;
input n_94;
input n_101;
input n_4;
input n_134;
input n_2;
input n_32;
input n_37;
input n_58;
input n_65;
input n_123;
input n_9;
input n_138;
input n_112;
input n_45;
input n_162;
input n_11;
input n_129;
input n_126;
input n_137;
input n_122;
input n_148;
input n_164;
input n_52;
input n_157;
input n_135;
input n_73;
input n_77;
input n_15;
input n_118;
input n_93;
input n_121;
input n_23;
input n_61;
input n_108;
input n_102;
input n_125;
input n_22;
input n_168;
input n_43;
input n_1;
input n_81;
input n_87;
input n_13;
input n_27;
input n_29;
input n_41;
input n_140;
input n_55;
input n_151;
input n_136;
input n_28;
input n_80;
input n_146;
input n_97;
input n_154;
input n_142;
input n_161;
input n_14;
input n_163;
input n_88;
input n_141;
input n_68;
input n_116;
input n_104;
input n_145;
input n_78;
input n_39;
input n_59;
input n_63;
input n_99;
input n_16;
input n_5;
input n_155;
input n_127;
input n_35;
input n_54;
input n_25;

output n_1869;

wire n_913;
wire n_1681;
wire n_1507;
wire n_1486;
wire n_589;
wire n_1174;
wire n_1469;
wire n_691;
wire n_1353;
wire n_1355;
wire n_423;
wire n_1383;
wire n_603;
wire n_373;
wire n_1250;
wire n_1169;
wire n_789;
wire n_850;
wire n_610;
wire n_245;
wire n_1713;
wire n_319;
wire n_1436;
wire n_690;
wire n_416;
wire n_1109;
wire n_1430;
wire n_525;
wire n_187;
wire n_1463;
wire n_1238;
wire n_1515;
wire n_817;
wire n_1837;
wire n_924;
wire n_781;
wire n_1566;
wire n_189;
wire n_717;
wire n_952;
wire n_864;
wire n_1096;
wire n_1379;
wire n_1706;
wire n_524;
wire n_1214;
wire n_634;
wire n_1839;
wire n_1246;
wire n_1138;
wire n_214;
wire n_1853;
wire n_764;
wire n_1503;
wire n_462;
wire n_1196;
wire n_1181;
wire n_410;
wire n_1187;
wire n_1131;
wire n_1225;
wire n_737;
wire n_1298;
wire n_1745;
wire n_1366;
wire n_232;
wire n_568;
wire n_1088;
wire n_1424;
wire n_766;
wire n_1835;
wire n_1457;
wire n_377;
wire n_1682;
wire n_1836;
wire n_520;
wire n_870;
wire n_1453;
wire n_279;
wire n_958;
wire n_945;
wire n_813;
wire n_419;
wire n_270;
wire n_338;
wire n_995;
wire n_285;
wire n_1184;
wire n_202;
wire n_1535;
wire n_500;
wire n_665;
wire n_754;
wire n_903;
wire n_871;
wire n_1073;
wire n_239;
wire n_402;
wire n_1277;
wire n_1746;
wire n_829;
wire n_1761;
wire n_1062;
wire n_339;
wire n_738;
wire n_1690;
wire n_672;
wire n_740;
wire n_1283;
wire n_1736;
wire n_1018;
wire n_259;
wire n_953;
wire n_1364;
wire n_1224;
wire n_1425;
wire n_625;
wire n_557;
wire n_1107;
wire n_1688;
wire n_989;
wire n_242;
wire n_645;
wire n_331;
wire n_559;
wire n_267;
wire n_495;
wire n_350;
wire n_381;
wire n_795;
wire n_721;
wire n_1084;
wire n_1718;
wire n_1276;
wire n_200;
wire n_1428;
wire n_1284;
wire n_1241;
wire n_821;
wire n_561;
wire n_770;
wire n_1514;
wire n_1528;
wire n_507;
wire n_486;
wire n_901;
wire n_569;
wire n_1145;
wire n_971;
wire n_787;
wire n_1650;
wire n_1519;
wire n_1195;
wire n_1522;
wire n_518;
wire n_1207;
wire n_222;
wire n_786;
wire n_1404;
wire n_868;
wire n_1847;
wire n_1542;
wire n_1314;
wire n_1512;
wire n_1539;
wire n_884;
wire n_1851;
wire n_1415;
wire n_1034;
wire n_1652;
wire n_1676;
wire n_1085;
wire n_277;
wire n_1636;
wire n_432;
wire n_293;
wire n_823;
wire n_620;
wire n_1074;
wire n_859;
wire n_1765;
wire n_587;
wire n_693;
wire n_863;
wire n_303;
wire n_1254;
wire n_929;
wire n_206;
wire n_352;
wire n_899;
wire n_1703;
wire n_611;
wire n_1295;
wire n_1850;
wire n_365;
wire n_238;
wire n_1013;
wire n_1495;
wire n_1637;
wire n_334;
wire n_192;
wire n_661;
wire n_1751;
wire n_300;
wire n_533;
wire n_438;
wire n_1560;
wire n_1654;
wire n_1548;
wire n_1811;
wire n_440;
wire n_273;
wire n_1396;
wire n_1230;
wire n_612;
wire n_333;
wire n_1840;
wire n_376;
wire n_512;
wire n_1597;
wire n_1771;
wire n_1544;
wire n_579;
wire n_844;
wire n_1012;
wire n_1267;
wire n_1354;
wire n_1790;
wire n_1213;
wire n_237;
wire n_780;
wire n_1021;
wire n_1443;
wire n_491;
wire n_1465;
wire n_1595;
wire n_1142;
wire n_1140;
wire n_705;
wire n_570;
wire n_260;
wire n_942;
wire n_1437;
wire n_1378;
wire n_461;
wire n_1121;
wire n_1416;
wire n_209;
wire n_490;
wire n_1461;
wire n_1391;
wire n_225;
wire n_1599;
wire n_1006;
wire n_1830;
wire n_575;
wire n_546;
wire n_503;
wire n_1112;
wire n_700;
wire n_1159;
wire n_772;
wire n_1216;
wire n_1245;
wire n_1669;
wire n_1675;
wire n_676;
wire n_1838;
wire n_1594;
wire n_680;
wire n_287;
wire n_1716;
wire n_302;
wire n_380;
wire n_1585;
wire n_1432;
wire n_249;
wire n_1108;
wire n_355;
wire n_212;
wire n_444;
wire n_851;
wire n_1590;
wire n_1351;
wire n_1274;
wire n_257;
wire n_652;
wire n_1819;
wire n_475;
wire n_947;
wire n_930;
wire n_1260;
wire n_1179;
wire n_468;
wire n_182;
wire n_696;
wire n_1442;
wire n_482;
wire n_798;
wire n_577;
wire n_1833;
wire n_407;
wire n_1691;
wire n_916;
wire n_1386;
wire n_912;
wire n_460;
wire n_1555;
wire n_1842;
wire n_366;
wire n_762;
wire n_1253;
wire n_1468;
wire n_1661;
wire n_555;
wire n_804;
wire n_1656;
wire n_1382;
wire n_966;
wire n_992;
wire n_955;
wire n_1182;
wire n_794;
wire n_1692;
wire n_1562;
wire n_514;
wire n_418;
wire n_1376;
wire n_513;
wire n_288;
wire n_179;
wire n_1292;
wire n_1178;
wire n_1435;
wire n_1750;
wire n_1026;
wire n_1506;
wire n_1610;
wire n_306;
wire n_203;
wire n_436;
wire n_324;
wire n_669;
wire n_931;
wire n_1491;
wire n_619;
wire n_337;
wire n_437;
wire n_274;
wire n_967;
wire n_1083;
wire n_1418;
wire n_746;
wire n_1357;
wire n_292;
wire n_1079;
wire n_1787;
wire n_1389;
wire n_615;
wire n_1139;
wire n_517;
wire n_1312;
wire n_1717;
wire n_1812;
wire n_824;
wire n_428;
wire n_892;
wire n_959;
wire n_1399;
wire n_1101;
wire n_1567;
wire n_1343;
wire n_563;
wire n_1855;
wire n_990;
wire n_1623;
wire n_867;
wire n_1226;
wire n_944;
wire n_749;
wire n_1780;
wire n_815;
wire n_542;
wire n_1340;
wire n_470;
wire n_1240;
wire n_1087;
wire n_632;
wire n_477;
wire n_650;
wire n_425;
wire n_1433;
wire n_1825;
wire n_1155;
wire n_1071;
wire n_712;
wire n_976;
wire n_909;
wire n_1392;
wire n_767;
wire n_1832;
wire n_1841;
wire n_1680;
wire n_964;
wire n_1627;
wire n_382;
wire n_489;
wire n_251;
wire n_974;
wire n_506;
wire n_1731;
wire n_799;
wire n_1147;
wire n_397;
wire n_471;
wire n_351;
wire n_965;
wire n_934;
wire n_1447;
wire n_1220;
wire n_356;
wire n_698;
wire n_1674;
wire n_307;
wire n_1209;
wire n_1020;
wire n_1563;
wire n_646;
wire n_1633;
wire n_404;
wire n_172;
wire n_1058;
wire n_347;
wire n_1042;
wire n_183;
wire n_1234;
wire n_479;
wire n_1578;
wire n_1455;
wire n_299;
wire n_836;
wire n_1279;
wire n_564;
wire n_205;
wire n_1029;
wire n_1247;
wire n_760;
wire n_522;
wire n_1568;
wire n_1483;
wire n_1363;
wire n_367;
wire n_1111;
wire n_970;
wire n_1689;
wire n_713;
wire n_1255;
wire n_1646;
wire n_598;
wire n_345;
wire n_1237;
wire n_927;
wire n_261;
wire n_1095;
wire n_1728;
wire n_370;
wire n_706;
wire n_286;
wire n_1401;
wire n_1419;
wire n_1531;
wire n_776;
wire n_424;
wire n_1651;
wire n_1387;
wire n_466;
wire n_1263;
wire n_346;
wire n_1817;
wire n_348;
wire n_552;
wire n_670;
wire n_1826;
wire n_379;
wire n_264;
wire n_441;
wire n_1032;
wire n_1217;
wire n_1496;
wire n_637;
wire n_1592;
wire n_327;
wire n_1259;
wire n_1177;
wire n_1231;
wire n_980;
wire n_1618;
wire n_1743;
wire n_905;
wire n_207;
wire n_720;
wire n_926;
wire n_194;
wire n_1802;
wire n_1163;
wire n_186;
wire n_1795;
wire n_1384;
wire n_1868;
wire n_1501;
wire n_1173;
wire n_1068;
wire n_1198;
wire n_1570;
wire n_487;
wire n_1518;
wire n_1456;
wire n_1648;
wire n_1413;
wire n_855;
wire n_808;
wire n_1365;
wire n_553;
wire n_1439;
wire n_814;
wire n_578;
wire n_1665;
wire n_1287;
wire n_405;
wire n_1611;
wire n_320;
wire n_1414;
wire n_1134;
wire n_1484;
wire n_647;
wire n_1423;
wire n_481;
wire n_600;
wire n_1053;
wire n_1609;
wire n_529;
wire n_502;
wire n_218;
wire n_1467;
wire n_247;
wire n_1828;
wire n_1798;
wire n_1304;
wire n_1608;
wire n_1744;
wire n_1105;
wire n_547;
wire n_439;
wire n_677;
wire n_604;
wire n_478;
wire n_703;
wire n_1349;
wire n_1709;
wire n_1061;
wire n_326;
wire n_681;
wire n_227;
wire n_874;
wire n_1278;
wire n_707;
wire n_983;
wire n_590;
wire n_699;
wire n_727;
wire n_301;
wire n_1726;
wire n_545;
wire n_1015;
wire n_1377;
wire n_1162;
wire n_536;
wire n_1614;
wire n_325;
wire n_1740;
wire n_1602;
wire n_688;
wire n_636;
wire n_427;
wire n_1098;
wire n_1490;
wire n_442;
wire n_777;
wire n_1553;
wire n_1080;
wire n_920;
wire n_1760;
wire n_1086;
wire n_1092;
wire n_986;
wire n_1104;
wire n_729;
wire n_887;
wire n_1122;
wire n_1205;
wire n_1408;
wire n_1693;
wire n_1132;
wire n_390;
wire n_1156;
wire n_501;
wire n_314;
wire n_1823;
wire n_1120;
wire n_1202;
wire n_627;
wire n_1188;
wire n_1498;
wire n_1371;
wire n_233;
wire n_957;
wire n_388;
wire n_1402;
wire n_1242;
wire n_1607;
wire n_1489;
wire n_1218;
wire n_221;
wire n_321;
wire n_1586;
wire n_861;
wire n_1543;
wire n_1431;
wire n_877;
wire n_1119;
wire n_1863;
wire n_1763;
wire n_1666;
wire n_1500;
wire n_616;
wire n_1055;
wire n_1395;
wire n_1346;
wire n_1189;
wire n_1089;
wire n_281;
wire n_1859;
wire n_262;
wire n_1502;
wire n_1523;
wire n_1478;
wire n_735;
wire n_297;
wire n_1005;
wire n_527;
wire n_1294;
wire n_1667;
wire n_888;
wire n_845;
wire n_1649;
wire n_1677;
wire n_1297;
wire n_178;
wire n_551;
wire n_417;
wire n_1708;
wire n_343;
wire n_1222;
wire n_1844;
wire n_582;
wire n_755;
wire n_1097;
wire n_1219;
wire n_1711;
wire n_710;
wire n_534;
wire n_1791;
wire n_1460;
wire n_1239;
wire n_278;
wire n_560;
wire n_890;
wire n_842;
wire n_451;
wire n_745;
wire n_1741;
wire n_1572;
wire n_1793;
wire n_742;
wire n_1081;
wire n_1373;
wire n_1388;
wire n_1266;
wire n_1540;
wire n_1719;
wire n_769;
wire n_1797;
wire n_1753;
wire n_1372;
wire n_476;
wire n_832;
wire n_535;
wire n_744;
wire n_982;
wire n_1800;
wire n_915;
wire n_215;
wire n_1075;
wire n_454;
wire n_298;
wire n_1331;
wire n_1529;
wire n_1227;
wire n_655;
wire n_1734;
wire n_1860;
wire n_403;
wire n_1007;
wire n_1580;
wire n_1319;
wire n_657;
wire n_837;
wire n_812;
wire n_606;
wire n_951;
wire n_862;
wire n_1700;
wire n_659;
wire n_1332;
wire n_509;
wire n_1854;
wire n_666;
wire n_1747;
wire n_430;
wire n_1206;
wire n_1729;
wire n_722;
wire n_1508;
wire n_1532;
wire n_1171;
wire n_1030;
wire n_785;
wire n_1309;
wire n_999;
wire n_1766;
wire n_1338;
wire n_1342;
wire n_456;
wire n_1867;
wire n_852;
wire n_1394;
wire n_704;
wire n_1060;
wire n_1044;
wire n_1714;
wire n_521;
wire n_873;
wire n_1301;
wire n_1748;
wire n_1243;
wire n_1400;
wire n_342;
wire n_1466;
wire n_1527;
wire n_1513;
wire n_358;
wire n_1783;
wire n_608;
wire n_1538;
wire n_1037;
wire n_1329;
wire n_317;
wire n_1545;
wire n_1257;
wire n_1480;
wire n_1668;
wire n_1605;
wire n_1078;
wire n_266;
wire n_1161;
wire n_811;
wire n_624;
wire n_791;
wire n_876;
wire n_618;
wire n_1191;
wire n_736;
wire n_1025;
wire n_1215;
wire n_241;
wire n_1449;
wire n_687;
wire n_797;
wire n_1786;
wire n_480;
wire n_1327;
wire n_1475;
wire n_211;
wire n_642;
wire n_1804;
wire n_408;
wire n_1406;
wire n_595;
wire n_1405;
wire n_602;
wire n_1757;
wire n_592;
wire n_1499;
wire n_854;
wire n_1318;
wire n_393;
wire n_1632;
wire n_1769;
wire n_474;
wire n_805;
wire n_295;
wire n_1658;
wire n_190;
wire n_1072;
wire n_695;
wire n_1526;
wire n_1305;
wire n_180;
wire n_730;
wire n_386;
wire n_1596;
wire n_1281;
wire n_516;
wire n_1137;
wire n_1258;
wire n_197;
wire n_640;
wire n_463;
wire n_1476;
wire n_1524;
wire n_1733;
wire n_1856;
wire n_943;
wire n_1118;
wire n_678;
wire n_651;
wire n_1293;
wire n_961;
wire n_469;
wire n_1046;
wire n_1807;
wire n_726;
wire n_1123;
wire n_1657;
wire n_878;
wire n_1784;
wire n_771;
wire n_1321;
wire n_752;
wire n_1488;
wire n_985;
wire n_421;
wire n_1330;
wire n_906;
wire n_1180;
wire n_1697;
wire n_283;
wire n_806;
wire n_1350;
wire n_1556;
wire n_649;
wire n_1561;
wire n_374;
wire n_1352;
wire n_1824;
wire n_643;
wire n_1492;
wire n_226;
wire n_1441;
wire n_1822;
wire n_682;
wire n_1616;
wire n_819;
wire n_586;
wire n_1324;
wire n_1429;
wire n_1778;
wire n_1776;
wire n_686;
wire n_605;
wire n_1154;
wire n_584;
wire n_1557;
wire n_1759;
wire n_1829;
wire n_1130;
wire n_1450;
wire n_349;
wire n_756;
wire n_1016;
wire n_1149;
wire n_1505;
wire n_979;
wire n_1642;
wire n_1815;
wire n_897;
wire n_949;
wire n_1493;
wire n_515;
wire n_807;
wire n_891;
wire n_885;
wire n_1659;
wire n_198;
wire n_1864;
wire n_1208;
wire n_396;
wire n_802;
wire n_1151;
wire n_554;
wire n_960;
wire n_1256;
wire n_714;
wire n_790;
wire n_354;
wire n_725;
wire n_1577;
wire n_1448;
wire n_1009;
wire n_230;
wire n_1133;
wire n_883;
wire n_473;
wire n_1852;
wire n_801;
wire n_1286;
wire n_818;
wire n_1685;
wire n_779;
wire n_594;
wire n_1397;
wire n_1052;
wire n_272;
wire n_1333;
wire n_1306;
wire n_1849;
wire n_833;
wire n_1426;
wire n_879;
wire n_1117;
wire n_422;
wire n_1269;
wire n_1303;
wire n_1547;
wire n_1438;
wire n_1541;
wire n_597;
wire n_1047;
wire n_1472;
wire n_1593;
wire n_1050;
wire n_566;
wire n_169;
wire n_1201;
wire n_1288;
wire n_173;
wire n_858;
wire n_1185;
wire n_335;
wire n_1035;
wire n_1143;
wire n_344;
wire n_426;
wire n_433;
wire n_398;
wire n_210;
wire n_1090;
wire n_1367;
wire n_253;
wire n_928;
wire n_1153;
wire n_271;
wire n_465;
wire n_825;
wire n_1103;
wire n_732;
wire n_1565;
wire n_1192;
wire n_224;
wire n_894;
wire n_1380;
wire n_1624;
wire n_1801;
wire n_420;
wire n_1291;
wire n_562;
wire n_748;
wire n_510;
wire n_1045;
wire n_256;
wire n_1160;
wire n_1023;
wire n_988;
wire n_330;
wire n_914;
wire n_400;
wire n_689;
wire n_1116;
wire n_282;
wire n_328;
wire n_368;
wire n_467;
wire n_1511;
wire n_1422;
wire n_644;
wire n_1197;
wire n_276;
wire n_497;
wire n_1165;
wire n_1641;
wire n_538;
wire n_1517;
wire n_576;
wire n_843;
wire n_511;
wire n_455;
wire n_429;
wire n_588;
wire n_638;
wire n_1307;
wire n_1128;
wire n_1671;
wire n_1417;
wire n_1048;
wire n_775;
wire n_667;
wire n_1049;
wire n_869;
wire n_846;
wire n_1398;
wire n_1356;
wire n_1341;
wire n_1504;
wire n_1773;
wire n_1440;
wire n_1370;
wire n_1603;
wire n_305;
wire n_312;
wire n_728;
wire n_413;
wire n_715;
wire n_889;
wire n_1066;
wire n_1549;
wire n_935;
wire n_685;
wire n_911;
wire n_361;
wire n_623;
wire n_1712;
wire n_1403;
wire n_1065;
wire n_453;
wire n_1534;
wire n_810;
wire n_1290;
wire n_181;
wire n_617;
wire n_543;
wire n_1362;
wire n_1559;
wire n_236;
wire n_683;
wire n_601;
wire n_565;
wire n_628;
wire n_1300;
wire n_743;
wire n_1194;
wire n_1647;
wire n_1546;
wire n_1420;
wire n_907;
wire n_1454;
wire n_660;
wire n_464;
wire n_962;
wire n_941;
wire n_1210;
wire n_847;
wire n_747;
wire n_1622;
wire n_1135;
wire n_918;
wire n_639;
wire n_452;
wire n_673;
wire n_1038;
wire n_414;
wire n_571;
wire n_1521;
wire n_1694;
wire n_284;
wire n_593;
wire n_1695;
wire n_1164;
wire n_609;
wire n_1193;
wire n_1345;
wire n_613;
wire n_1022;
wire n_1336;
wire n_1033;
wire n_1774;
wire n_409;
wire n_171;
wire n_519;
wire n_384;
wire n_1166;
wire n_1056;
wire n_526;
wire n_1767;
wire n_1040;
wire n_674;
wire n_1158;
wire n_316;
wire n_1444;
wire n_1803;
wire n_820;
wire n_1749;
wire n_872;
wire n_1653;
wire n_254;
wire n_1157;
wire n_1584;
wire n_234;
wire n_848;
wire n_1664;
wire n_280;
wire n_629;
wire n_1739;
wire n_1814;
wire n_532;
wire n_1789;
wire n_763;
wire n_540;
wire n_216;
wire n_692;
wire n_1857;
wire n_984;
wire n_1687;
wire n_223;
wire n_1552;
wire n_750;
wire n_834;
wire n_1612;
wire n_800;
wire n_1816;
wire n_1756;
wire n_1606;
wire n_395;
wire n_621;
wire n_1587;
wire n_213;
wire n_1772;
wire n_1014;
wire n_724;
wire n_1427;
wire n_1481;
wire n_493;
wire n_1311;
wire n_1589;
wire n_1100;
wire n_585;
wire n_875;
wire n_1617;
wire n_827;
wire n_697;
wire n_622;
wire n_1626;
wire n_1335;
wire n_1715;
wire n_296;
wire n_880;
wire n_793;
wire n_1175;
wire n_751;
wire n_1027;
wire n_1070;
wire n_1621;
wire n_739;
wire n_1485;
wire n_1028;
wire n_1221;
wire n_530;
wire n_1785;
wire n_792;
wire n_1262;
wire n_580;
wire n_1579;
wire n_494;
wire n_434;
wire n_975;
wire n_229;
wire n_394;
wire n_923;
wire n_1645;
wire n_1124;
wire n_1381;
wire n_1494;
wire n_932;
wire n_1183;
wire n_1326;
wire n_1805;
wire n_981;
wire n_1110;
wire n_1758;
wire n_243;
wire n_1407;
wire n_185;
wire n_1204;
wire n_1554;
wire n_994;
wire n_1360;
wire n_973;
wire n_268;
wire n_972;
wire n_184;
wire n_856;
wire n_1248;
wire n_1176;
wire n_1564;
wire n_1054;
wire n_508;
wire n_1679;
wire n_1858;
wire n_353;
wire n_1678;
wire n_1482;
wire n_1361;
wire n_1601;
wire n_1057;
wire n_191;
wire n_1834;
wire n_978;
wire n_1011;
wire n_1520;
wire n_1509;
wire n_828;
wire n_322;
wire n_1411;
wire n_1359;
wire n_558;
wire n_1721;
wire n_653;
wire n_1445;
wire n_1317;
wire n_783;
wire n_556;
wire n_1127;
wire n_170;
wire n_1536;
wire n_1471;
wire n_1008;
wire n_332;
wire n_581;
wire n_294;
wire n_1024;
wire n_830;
wire n_176;
wire n_987;
wire n_936;
wire n_1620;
wire n_1385;
wire n_1525;
wire n_541;
wire n_499;
wire n_1775;
wire n_788;
wire n_908;
wire n_1036;
wire n_341;
wire n_1270;
wire n_1167;
wire n_1272;
wire n_549;
wire n_591;
wire n_969;
wire n_919;
wire n_1663;
wire n_1625;
wire n_318;
wire n_1458;
wire n_244;
wire n_679;
wire n_1630;
wire n_220;
wire n_663;
wire n_1720;
wire n_443;
wire n_1412;
wire n_1738;
wire n_1550;
wire n_528;
wire n_1358;
wire n_1200;
wire n_387;
wire n_406;
wire n_826;
wire n_1735;
wire n_1788;
wire n_391;
wire n_940;
wire n_1537;
wire n_1077;
wire n_607;
wire n_956;
wire n_445;
wire n_765;
wire n_1809;
wire n_1843;
wire n_1268;
wire n_385;
wire n_917;
wire n_1271;
wire n_372;
wire n_1530;
wire n_631;
wire n_399;
wire n_1170;
wire n_1261;
wire n_702;
wire n_898;
wire n_857;
wire n_363;
wire n_968;
wire n_1067;
wire n_1235;
wire n_1323;
wire n_1462;
wire n_1064;
wire n_633;
wire n_900;
wire n_1446;
wire n_1282;
wire n_1701;
wire n_1093;
wire n_1551;
wire n_1755;
wire n_1285;
wire n_193;
wire n_761;
wire n_733;
wire n_731;
wire n_336;
wire n_1813;
wire n_315;
wire n_311;
wire n_1452;
wire n_1573;
wire n_668;
wire n_758;
wire n_1106;
wire n_648;
wire n_784;
wire n_269;
wire n_816;
wire n_1322;
wire n_1473;
wire n_835;
wire n_446;
wire n_1076;
wire n_1348;
wire n_753;
wire n_1770;
wire n_701;
wire n_1003;
wire n_1125;
wire n_1710;
wire n_1865;
wire n_309;
wire n_1344;
wire n_1390;
wire n_401;
wire n_485;
wire n_1792;
wire n_504;
wire n_483;
wire n_435;
wire n_1141;
wire n_1629;
wire n_291;
wire n_1640;
wire n_822;
wire n_1094;
wire n_840;
wire n_1459;
wire n_1510;
wire n_1099;
wire n_839;
wire n_1754;
wire n_759;
wire n_567;
wire n_369;
wire n_240;
wire n_1727;
wire n_1575;
wire n_1848;
wire n_1172;
wire n_614;
wire n_1212;
wire n_831;
wire n_778;
wire n_1619;
wire n_188;
wire n_323;
wire n_550;
wire n_1315;
wire n_1660;
wire n_997;
wire n_635;
wire n_694;
wire n_1643;
wire n_1320;
wire n_1113;
wire n_248;
wire n_1152;
wire n_1845;
wire n_921;
wire n_1615;
wire n_1236;
wire n_228;
wire n_1265;
wire n_1576;
wire n_1470;
wire n_671;
wire n_1533;
wire n_1806;
wire n_1409;
wire n_1148;
wire n_1588;
wire n_1684;
wire n_1673;
wire n_1334;
wire n_654;
wire n_1275;
wire n_488;
wire n_904;
wire n_505;
wire n_1696;
wire n_498;
wire n_1059;
wire n_684;
wire n_1039;
wire n_539;
wire n_1150;
wire n_977;
wire n_449;
wire n_392;
wire n_1628;
wire n_1289;
wire n_1831;
wire n_1497;
wire n_1866;
wire n_459;
wire n_1136;
wire n_1782;
wire n_458;
wire n_1190;
wire n_1600;
wire n_1144;
wire n_383;
wire n_838;
wire n_1558;
wire n_1316;
wire n_175;
wire n_950;
wire n_1017;
wire n_711;
wire n_734;
wire n_723;
wire n_1393;
wire n_658;
wire n_630;
wire n_1369;
wire n_362;
wire n_310;
wire n_1781;
wire n_709;
wire n_809;
wire n_1686;
wire n_235;
wire n_881;
wire n_1019;
wire n_1477;
wire n_1777;
wire n_662;
wire n_641;
wire n_910;
wire n_290;
wire n_741;
wire n_939;
wire n_1410;
wire n_371;
wire n_199;
wire n_217;
wire n_1114;
wire n_1325;
wire n_1742;
wire n_708;
wire n_308;
wire n_1223;
wire n_201;
wire n_1768;
wire n_572;
wire n_1199;
wire n_865;
wire n_1273;
wire n_1041;
wire n_993;
wire n_1862;
wire n_948;
wire n_922;
wire n_1004;
wire n_1810;
wire n_448;
wire n_1347;
wire n_860;
wire n_1043;
wire n_255;
wire n_450;
wire n_1764;
wire n_896;
wire n_1737;
wire n_1479;
wire n_1613;
wire n_902;
wire n_1031;
wire n_1723;
wire n_1638;
wire n_853;
wire n_716;
wire n_1571;
wire n_1698;
wire n_196;
wire n_1337;
wire n_774;
wire n_933;
wire n_1779;
wire n_596;
wire n_954;
wire n_1168;
wire n_1821;
wire n_219;
wire n_1310;
wire n_231;
wire n_656;
wire n_492;
wire n_574;
wire n_252;
wire n_664;
wire n_1591;
wire n_1229;
wire n_1683;
wire n_1732;
wire n_415;
wire n_1280;
wire n_544;
wire n_1516;
wire n_1186;
wire n_1705;
wire n_599;
wire n_768;
wire n_1091;
wire n_537;
wire n_1063;
wire n_991;
wire n_389;
wire n_1724;
wire n_1670;
wire n_1707;
wire n_1799;
wire n_1126;
wire n_195;
wire n_1846;
wire n_938;
wire n_1328;
wire n_895;
wire n_304;
wire n_1639;
wire n_583;
wire n_1302;
wire n_1000;
wire n_313;
wire n_626;
wire n_378;
wire n_1581;
wire n_946;
wire n_757;
wire n_375;
wire n_1655;
wire n_1818;
wire n_1146;
wire n_1634;
wire n_1203;
wire n_998;
wire n_1699;
wire n_1598;
wire n_472;
wire n_937;
wire n_1474;
wire n_265;
wire n_1583;
wire n_1604;
wire n_208;
wire n_1631;
wire n_1702;
wire n_174;
wire n_275;
wire n_1794;
wire n_1375;
wire n_204;
wire n_1232;
wire n_996;
wire n_1211;
wire n_1368;
wire n_963;
wire n_1264;
wire n_1082;
wire n_1725;
wire n_496;
wire n_1827;
wire n_866;
wire n_246;
wire n_925;
wire n_1752;
wire n_1313;
wire n_1001;
wire n_1722;
wire n_1115;
wire n_1339;
wire n_1002;
wire n_1644;
wire n_1051;
wire n_719;
wire n_263;
wire n_1102;
wire n_360;
wire n_1129;
wire n_1252;
wire n_250;
wire n_1464;
wire n_1296;
wire n_773;
wire n_1010;
wire n_882;
wire n_1249;
wire n_803;
wire n_329;
wire n_718;
wire n_1434;
wire n_340;
wire n_1569;
wire n_289;
wire n_548;
wire n_523;
wire n_1662;
wire n_457;
wire n_1299;
wire n_177;
wire n_782;
wire n_364;
wire n_258;
wire n_431;
wire n_1861;
wire n_1228;
wire n_1244;
wire n_1796;
wire n_411;
wire n_484;
wire n_849;
wire n_1820;
wire n_357;
wire n_412;
wire n_1251;
wire n_447;
wire n_1421;
wire n_1762;
wire n_1233;
wire n_1808;
wire n_1574;
wire n_1672;
wire n_1635;
wire n_1704;
wire n_893;
wire n_1582;
wire n_841;
wire n_886;
wire n_1069;
wire n_359;
wire n_1308;
wire n_573;
wire n_796;
wire n_531;
wire n_1730;
wire n_1374;
wire n_1451;
wire n_1487;
wire n_675;

BUFx6f_ASAP7_75t_L g169 ( 
.A(n_102),
.Y(n_169)
);

CKINVDCx5p33_ASAP7_75t_R g170 ( 
.A(n_118),
.Y(n_170)
);

BUFx6f_ASAP7_75t_L g171 ( 
.A(n_68),
.Y(n_171)
);

BUFx2_ASAP7_75t_L g172 ( 
.A(n_111),
.Y(n_172)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_32),
.Y(n_173)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_90),
.Y(n_174)
);

CKINVDCx5p33_ASAP7_75t_R g175 ( 
.A(n_131),
.Y(n_175)
);

BUFx3_ASAP7_75t_L g176 ( 
.A(n_124),
.Y(n_176)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_7),
.Y(n_177)
);

CKINVDCx5p33_ASAP7_75t_R g178 ( 
.A(n_9),
.Y(n_178)
);

CKINVDCx5p33_ASAP7_75t_R g179 ( 
.A(n_24),
.Y(n_179)
);

BUFx6f_ASAP7_75t_L g180 ( 
.A(n_62),
.Y(n_180)
);

BUFx2_ASAP7_75t_SL g181 ( 
.A(n_154),
.Y(n_181)
);

CKINVDCx20_ASAP7_75t_R g182 ( 
.A(n_59),
.Y(n_182)
);

CKINVDCx5p33_ASAP7_75t_R g183 ( 
.A(n_92),
.Y(n_183)
);

CKINVDCx5p33_ASAP7_75t_R g184 ( 
.A(n_101),
.Y(n_184)
);

CKINVDCx5p33_ASAP7_75t_R g185 ( 
.A(n_159),
.Y(n_185)
);

CKINVDCx5p33_ASAP7_75t_R g186 ( 
.A(n_23),
.Y(n_186)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_46),
.Y(n_187)
);

INVx2_ASAP7_75t_L g188 ( 
.A(n_28),
.Y(n_188)
);

BUFx6f_ASAP7_75t_L g189 ( 
.A(n_126),
.Y(n_189)
);

CKINVDCx5p33_ASAP7_75t_R g190 ( 
.A(n_122),
.Y(n_190)
);

CKINVDCx20_ASAP7_75t_R g191 ( 
.A(n_32),
.Y(n_191)
);

CKINVDCx5p33_ASAP7_75t_R g192 ( 
.A(n_79),
.Y(n_192)
);

CKINVDCx20_ASAP7_75t_R g193 ( 
.A(n_24),
.Y(n_193)
);

INVx1_ASAP7_75t_SL g194 ( 
.A(n_11),
.Y(n_194)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_135),
.Y(n_195)
);

INVx2_ASAP7_75t_L g196 ( 
.A(n_140),
.Y(n_196)
);

INVx1_ASAP7_75t_SL g197 ( 
.A(n_49),
.Y(n_197)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_166),
.Y(n_198)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_73),
.Y(n_199)
);

CKINVDCx5p33_ASAP7_75t_R g200 ( 
.A(n_45),
.Y(n_200)
);

CKINVDCx5p33_ASAP7_75t_R g201 ( 
.A(n_30),
.Y(n_201)
);

CKINVDCx5p33_ASAP7_75t_R g202 ( 
.A(n_70),
.Y(n_202)
);

CKINVDCx5p33_ASAP7_75t_R g203 ( 
.A(n_147),
.Y(n_203)
);

CKINVDCx20_ASAP7_75t_R g204 ( 
.A(n_109),
.Y(n_204)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_6),
.Y(n_205)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_4),
.Y(n_206)
);

CKINVDCx5p33_ASAP7_75t_R g207 ( 
.A(n_84),
.Y(n_207)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_75),
.Y(n_208)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_23),
.Y(n_209)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_51),
.Y(n_210)
);

CKINVDCx5p33_ASAP7_75t_R g211 ( 
.A(n_42),
.Y(n_211)
);

BUFx5_ASAP7_75t_L g212 ( 
.A(n_16),
.Y(n_212)
);

INVx1_ASAP7_75t_SL g213 ( 
.A(n_83),
.Y(n_213)
);

CKINVDCx20_ASAP7_75t_R g214 ( 
.A(n_76),
.Y(n_214)
);

CKINVDCx5p33_ASAP7_75t_R g215 ( 
.A(n_34),
.Y(n_215)
);

CKINVDCx5p33_ASAP7_75t_R g216 ( 
.A(n_163),
.Y(n_216)
);

CKINVDCx5p33_ASAP7_75t_R g217 ( 
.A(n_61),
.Y(n_217)
);

CKINVDCx5p33_ASAP7_75t_R g218 ( 
.A(n_104),
.Y(n_218)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_106),
.Y(n_219)
);

BUFx3_ASAP7_75t_L g220 ( 
.A(n_33),
.Y(n_220)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_36),
.Y(n_221)
);

CKINVDCx5p33_ASAP7_75t_R g222 ( 
.A(n_161),
.Y(n_222)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_52),
.Y(n_223)
);

CKINVDCx5p33_ASAP7_75t_R g224 ( 
.A(n_26),
.Y(n_224)
);

INVx1_ASAP7_75t_SL g225 ( 
.A(n_44),
.Y(n_225)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_165),
.Y(n_226)
);

CKINVDCx5p33_ASAP7_75t_R g227 ( 
.A(n_119),
.Y(n_227)
);

CKINVDCx5p33_ASAP7_75t_R g228 ( 
.A(n_146),
.Y(n_228)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_41),
.Y(n_229)
);

BUFx3_ASAP7_75t_L g230 ( 
.A(n_29),
.Y(n_230)
);

HB1xp67_ASAP7_75t_L g231 ( 
.A(n_66),
.Y(n_231)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_128),
.Y(n_232)
);

CKINVDCx20_ASAP7_75t_R g233 ( 
.A(n_17),
.Y(n_233)
);

CKINVDCx5p33_ASAP7_75t_R g234 ( 
.A(n_120),
.Y(n_234)
);

BUFx3_ASAP7_75t_L g235 ( 
.A(n_60),
.Y(n_235)
);

CKINVDCx5p33_ASAP7_75t_R g236 ( 
.A(n_100),
.Y(n_236)
);

CKINVDCx5p33_ASAP7_75t_R g237 ( 
.A(n_108),
.Y(n_237)
);

CKINVDCx5p33_ASAP7_75t_R g238 ( 
.A(n_37),
.Y(n_238)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_21),
.Y(n_239)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_142),
.Y(n_240)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_56),
.Y(n_241)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_115),
.Y(n_242)
);

CKINVDCx20_ASAP7_75t_R g243 ( 
.A(n_36),
.Y(n_243)
);

CKINVDCx5p33_ASAP7_75t_R g244 ( 
.A(n_20),
.Y(n_244)
);

CKINVDCx5p33_ASAP7_75t_R g245 ( 
.A(n_18),
.Y(n_245)
);

CKINVDCx20_ASAP7_75t_R g246 ( 
.A(n_38),
.Y(n_246)
);

CKINVDCx5p33_ASAP7_75t_R g247 ( 
.A(n_87),
.Y(n_247)
);

INVxp67_ASAP7_75t_L g248 ( 
.A(n_139),
.Y(n_248)
);

CKINVDCx20_ASAP7_75t_R g249 ( 
.A(n_55),
.Y(n_249)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_99),
.Y(n_250)
);

CKINVDCx5p33_ASAP7_75t_R g251 ( 
.A(n_13),
.Y(n_251)
);

BUFx6f_ASAP7_75t_L g252 ( 
.A(n_143),
.Y(n_252)
);

CKINVDCx5p33_ASAP7_75t_R g253 ( 
.A(n_112),
.Y(n_253)
);

CKINVDCx5p33_ASAP7_75t_R g254 ( 
.A(n_4),
.Y(n_254)
);

CKINVDCx5p33_ASAP7_75t_R g255 ( 
.A(n_152),
.Y(n_255)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_69),
.Y(n_256)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_157),
.Y(n_257)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_82),
.Y(n_258)
);

CKINVDCx5p33_ASAP7_75t_R g259 ( 
.A(n_158),
.Y(n_259)
);

CKINVDCx5p33_ASAP7_75t_R g260 ( 
.A(n_48),
.Y(n_260)
);

CKINVDCx5p33_ASAP7_75t_R g261 ( 
.A(n_130),
.Y(n_261)
);

CKINVDCx5p33_ASAP7_75t_R g262 ( 
.A(n_103),
.Y(n_262)
);

CKINVDCx5p33_ASAP7_75t_R g263 ( 
.A(n_50),
.Y(n_263)
);

CKINVDCx16_ASAP7_75t_R g264 ( 
.A(n_21),
.Y(n_264)
);

CKINVDCx5p33_ASAP7_75t_R g265 ( 
.A(n_1),
.Y(n_265)
);

CKINVDCx5p33_ASAP7_75t_R g266 ( 
.A(n_38),
.Y(n_266)
);

INVx2_ASAP7_75t_L g267 ( 
.A(n_34),
.Y(n_267)
);

INVx2_ASAP7_75t_L g268 ( 
.A(n_86),
.Y(n_268)
);

CKINVDCx5p33_ASAP7_75t_R g269 ( 
.A(n_81),
.Y(n_269)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_18),
.Y(n_270)
);

CKINVDCx20_ASAP7_75t_R g271 ( 
.A(n_15),
.Y(n_271)
);

INVx1_ASAP7_75t_SL g272 ( 
.A(n_3),
.Y(n_272)
);

CKINVDCx5p33_ASAP7_75t_R g273 ( 
.A(n_85),
.Y(n_273)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_127),
.Y(n_274)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_96),
.Y(n_275)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_26),
.Y(n_276)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_137),
.Y(n_277)
);

CKINVDCx5p33_ASAP7_75t_R g278 ( 
.A(n_71),
.Y(n_278)
);

CKINVDCx5p33_ASAP7_75t_R g279 ( 
.A(n_29),
.Y(n_279)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_136),
.Y(n_280)
);

CKINVDCx5p33_ASAP7_75t_R g281 ( 
.A(n_155),
.Y(n_281)
);

CKINVDCx5p33_ASAP7_75t_R g282 ( 
.A(n_5),
.Y(n_282)
);

CKINVDCx16_ASAP7_75t_R g283 ( 
.A(n_11),
.Y(n_283)
);

INVxp67_ASAP7_75t_SL g284 ( 
.A(n_89),
.Y(n_284)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_63),
.Y(n_285)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_113),
.Y(n_286)
);

CKINVDCx5p33_ASAP7_75t_R g287 ( 
.A(n_141),
.Y(n_287)
);

CKINVDCx5p33_ASAP7_75t_R g288 ( 
.A(n_3),
.Y(n_288)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_145),
.Y(n_289)
);

CKINVDCx5p33_ASAP7_75t_R g290 ( 
.A(n_58),
.Y(n_290)
);

CKINVDCx5p33_ASAP7_75t_R g291 ( 
.A(n_134),
.Y(n_291)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_28),
.Y(n_292)
);

HB1xp67_ASAP7_75t_L g293 ( 
.A(n_156),
.Y(n_293)
);

CKINVDCx16_ASAP7_75t_R g294 ( 
.A(n_65),
.Y(n_294)
);

CKINVDCx5p33_ASAP7_75t_R g295 ( 
.A(n_12),
.Y(n_295)
);

CKINVDCx16_ASAP7_75t_R g296 ( 
.A(n_148),
.Y(n_296)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_20),
.Y(n_297)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_6),
.Y(n_298)
);

CKINVDCx20_ASAP7_75t_R g299 ( 
.A(n_117),
.Y(n_299)
);

CKINVDCx5p33_ASAP7_75t_R g300 ( 
.A(n_160),
.Y(n_300)
);

CKINVDCx5p33_ASAP7_75t_R g301 ( 
.A(n_25),
.Y(n_301)
);

INVx1_ASAP7_75t_SL g302 ( 
.A(n_80),
.Y(n_302)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_7),
.Y(n_303)
);

CKINVDCx20_ASAP7_75t_R g304 ( 
.A(n_150),
.Y(n_304)
);

HB1xp67_ASAP7_75t_L g305 ( 
.A(n_47),
.Y(n_305)
);

CKINVDCx5p33_ASAP7_75t_R g306 ( 
.A(n_33),
.Y(n_306)
);

INVx2_ASAP7_75t_SL g307 ( 
.A(n_149),
.Y(n_307)
);

CKINVDCx5p33_ASAP7_75t_R g308 ( 
.A(n_91),
.Y(n_308)
);

CKINVDCx5p33_ASAP7_75t_R g309 ( 
.A(n_15),
.Y(n_309)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_8),
.Y(n_310)
);

CKINVDCx5p33_ASAP7_75t_R g311 ( 
.A(n_1),
.Y(n_311)
);

CKINVDCx5p33_ASAP7_75t_R g312 ( 
.A(n_77),
.Y(n_312)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_144),
.Y(n_313)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_153),
.Y(n_314)
);

CKINVDCx5p33_ASAP7_75t_R g315 ( 
.A(n_46),
.Y(n_315)
);

CKINVDCx5p33_ASAP7_75t_R g316 ( 
.A(n_30),
.Y(n_316)
);

CKINVDCx5p33_ASAP7_75t_R g317 ( 
.A(n_167),
.Y(n_317)
);

CKINVDCx20_ASAP7_75t_R g318 ( 
.A(n_107),
.Y(n_318)
);

CKINVDCx5p33_ASAP7_75t_R g319 ( 
.A(n_5),
.Y(n_319)
);

CKINVDCx5p33_ASAP7_75t_R g320 ( 
.A(n_14),
.Y(n_320)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_45),
.Y(n_321)
);

CKINVDCx20_ASAP7_75t_R g322 ( 
.A(n_12),
.Y(n_322)
);

CKINVDCx5p33_ASAP7_75t_R g323 ( 
.A(n_22),
.Y(n_323)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_14),
.Y(n_324)
);

CKINVDCx5p33_ASAP7_75t_R g325 ( 
.A(n_168),
.Y(n_325)
);

CKINVDCx5p33_ASAP7_75t_R g326 ( 
.A(n_129),
.Y(n_326)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_39),
.Y(n_327)
);

CKINVDCx5p33_ASAP7_75t_R g328 ( 
.A(n_39),
.Y(n_328)
);

INVx1_ASAP7_75t_SL g329 ( 
.A(n_17),
.Y(n_329)
);

CKINVDCx5p33_ASAP7_75t_R g330 ( 
.A(n_138),
.Y(n_330)
);

CKINVDCx5p33_ASAP7_75t_R g331 ( 
.A(n_37),
.Y(n_331)
);

BUFx6f_ASAP7_75t_L g332 ( 
.A(n_41),
.Y(n_332)
);

CKINVDCx5p33_ASAP7_75t_R g333 ( 
.A(n_116),
.Y(n_333)
);

INVx2_ASAP7_75t_SL g334 ( 
.A(n_44),
.Y(n_334)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_110),
.Y(n_335)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_132),
.Y(n_336)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_220),
.Y(n_337)
);

INVxp33_ASAP7_75t_SL g338 ( 
.A(n_186),
.Y(n_338)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_212),
.Y(n_339)
);

CKINVDCx20_ASAP7_75t_R g340 ( 
.A(n_182),
.Y(n_340)
);

BUFx10_ASAP7_75t_L g341 ( 
.A(n_231),
.Y(n_341)
);

INVx1_ASAP7_75t_L g342 ( 
.A(n_220),
.Y(n_342)
);

CKINVDCx5p33_ASAP7_75t_R g343 ( 
.A(n_294),
.Y(n_343)
);

INVx1_ASAP7_75t_L g344 ( 
.A(n_230),
.Y(n_344)
);

INVx1_ASAP7_75t_L g345 ( 
.A(n_230),
.Y(n_345)
);

INVx1_ASAP7_75t_L g346 ( 
.A(n_212),
.Y(n_346)
);

INVx1_ASAP7_75t_L g347 ( 
.A(n_212),
.Y(n_347)
);

CKINVDCx5p33_ASAP7_75t_R g348 ( 
.A(n_296),
.Y(n_348)
);

CKINVDCx5p33_ASAP7_75t_R g349 ( 
.A(n_172),
.Y(n_349)
);

CKINVDCx5p33_ASAP7_75t_R g350 ( 
.A(n_182),
.Y(n_350)
);

BUFx3_ASAP7_75t_L g351 ( 
.A(n_176),
.Y(n_351)
);

INVx1_ASAP7_75t_L g352 ( 
.A(n_212),
.Y(n_352)
);

INVx1_ASAP7_75t_L g353 ( 
.A(n_212),
.Y(n_353)
);

INVx1_ASAP7_75t_L g354 ( 
.A(n_212),
.Y(n_354)
);

INVx1_ASAP7_75t_L g355 ( 
.A(n_212),
.Y(n_355)
);

INVx1_ASAP7_75t_L g356 ( 
.A(n_332),
.Y(n_356)
);

CKINVDCx5p33_ASAP7_75t_R g357 ( 
.A(n_204),
.Y(n_357)
);

INVx1_ASAP7_75t_L g358 ( 
.A(n_332),
.Y(n_358)
);

INVx1_ASAP7_75t_L g359 ( 
.A(n_332),
.Y(n_359)
);

INVx2_ASAP7_75t_L g360 ( 
.A(n_332),
.Y(n_360)
);

CKINVDCx14_ASAP7_75t_R g361 ( 
.A(n_204),
.Y(n_361)
);

BUFx2_ASAP7_75t_SL g362 ( 
.A(n_214),
.Y(n_362)
);

INVx2_ASAP7_75t_L g363 ( 
.A(n_176),
.Y(n_363)
);

CKINVDCx20_ASAP7_75t_R g364 ( 
.A(n_214),
.Y(n_364)
);

INVxp67_ASAP7_75t_SL g365 ( 
.A(n_188),
.Y(n_365)
);

INVx1_ASAP7_75t_L g366 ( 
.A(n_188),
.Y(n_366)
);

INVx2_ASAP7_75t_L g367 ( 
.A(n_235),
.Y(n_367)
);

INVx1_ASAP7_75t_L g368 ( 
.A(n_173),
.Y(n_368)
);

INVx1_ASAP7_75t_L g369 ( 
.A(n_177),
.Y(n_369)
);

INVx1_ASAP7_75t_L g370 ( 
.A(n_187),
.Y(n_370)
);

INVxp33_ASAP7_75t_SL g371 ( 
.A(n_186),
.Y(n_371)
);

INVx1_ASAP7_75t_L g372 ( 
.A(n_205),
.Y(n_372)
);

CKINVDCx16_ASAP7_75t_R g373 ( 
.A(n_264),
.Y(n_373)
);

INVx1_ASAP7_75t_L g374 ( 
.A(n_206),
.Y(n_374)
);

CKINVDCx20_ASAP7_75t_R g375 ( 
.A(n_249),
.Y(n_375)
);

INVx1_ASAP7_75t_L g376 ( 
.A(n_209),
.Y(n_376)
);

CKINVDCx5p33_ASAP7_75t_R g377 ( 
.A(n_249),
.Y(n_377)
);

CKINVDCx5p33_ASAP7_75t_R g378 ( 
.A(n_299),
.Y(n_378)
);

CKINVDCx5p33_ASAP7_75t_R g379 ( 
.A(n_299),
.Y(n_379)
);

INVx1_ASAP7_75t_L g380 ( 
.A(n_221),
.Y(n_380)
);

INVx1_ASAP7_75t_L g381 ( 
.A(n_229),
.Y(n_381)
);

INVx2_ASAP7_75t_L g382 ( 
.A(n_235),
.Y(n_382)
);

INVx1_ASAP7_75t_L g383 ( 
.A(n_239),
.Y(n_383)
);

INVx1_ASAP7_75t_L g384 ( 
.A(n_270),
.Y(n_384)
);

CKINVDCx16_ASAP7_75t_R g385 ( 
.A(n_283),
.Y(n_385)
);

INVx1_ASAP7_75t_L g386 ( 
.A(n_276),
.Y(n_386)
);

CKINVDCx5p33_ASAP7_75t_R g387 ( 
.A(n_304),
.Y(n_387)
);

CKINVDCx5p33_ASAP7_75t_R g388 ( 
.A(n_304),
.Y(n_388)
);

CKINVDCx20_ASAP7_75t_R g389 ( 
.A(n_318),
.Y(n_389)
);

CKINVDCx5p33_ASAP7_75t_R g390 ( 
.A(n_318),
.Y(n_390)
);

INVxp33_ASAP7_75t_L g391 ( 
.A(n_292),
.Y(n_391)
);

CKINVDCx5p33_ASAP7_75t_R g392 ( 
.A(n_183),
.Y(n_392)
);

CKINVDCx20_ASAP7_75t_R g393 ( 
.A(n_191),
.Y(n_393)
);

INVx1_ASAP7_75t_L g394 ( 
.A(n_297),
.Y(n_394)
);

INVxp67_ASAP7_75t_SL g395 ( 
.A(n_267),
.Y(n_395)
);

INVx1_ASAP7_75t_L g396 ( 
.A(n_298),
.Y(n_396)
);

INVx1_ASAP7_75t_L g397 ( 
.A(n_303),
.Y(n_397)
);

CKINVDCx5p33_ASAP7_75t_R g398 ( 
.A(n_183),
.Y(n_398)
);

INVx1_ASAP7_75t_L g399 ( 
.A(n_310),
.Y(n_399)
);

CKINVDCx5p33_ASAP7_75t_R g400 ( 
.A(n_184),
.Y(n_400)
);

INVxp67_ASAP7_75t_L g401 ( 
.A(n_334),
.Y(n_401)
);

HB1xp67_ASAP7_75t_L g402 ( 
.A(n_315),
.Y(n_402)
);

INVx1_ASAP7_75t_L g403 ( 
.A(n_321),
.Y(n_403)
);

INVxp67_ASAP7_75t_L g404 ( 
.A(n_334),
.Y(n_404)
);

INVx1_ASAP7_75t_L g405 ( 
.A(n_324),
.Y(n_405)
);

INVx1_ASAP7_75t_L g406 ( 
.A(n_267),
.Y(n_406)
);

CKINVDCx5p33_ASAP7_75t_R g407 ( 
.A(n_184),
.Y(n_407)
);

INVx1_ASAP7_75t_L g408 ( 
.A(n_196),
.Y(n_408)
);

CKINVDCx5p33_ASAP7_75t_R g409 ( 
.A(n_185),
.Y(n_409)
);

INVx1_ASAP7_75t_L g410 ( 
.A(n_196),
.Y(n_410)
);

INVx1_ASAP7_75t_L g411 ( 
.A(n_268),
.Y(n_411)
);

INVxp67_ASAP7_75t_L g412 ( 
.A(n_327),
.Y(n_412)
);

INVx1_ASAP7_75t_L g413 ( 
.A(n_268),
.Y(n_413)
);

CKINVDCx5p33_ASAP7_75t_R g414 ( 
.A(n_185),
.Y(n_414)
);

CKINVDCx20_ASAP7_75t_R g415 ( 
.A(n_191),
.Y(n_415)
);

CKINVDCx5p33_ASAP7_75t_R g416 ( 
.A(n_190),
.Y(n_416)
);

INVx2_ASAP7_75t_L g417 ( 
.A(n_174),
.Y(n_417)
);

INVxp67_ASAP7_75t_SL g418 ( 
.A(n_293),
.Y(n_418)
);

BUFx2_ASAP7_75t_L g419 ( 
.A(n_343),
.Y(n_419)
);

INVx1_ASAP7_75t_L g420 ( 
.A(n_339),
.Y(n_420)
);

NAND2xp5_ASAP7_75t_L g421 ( 
.A(n_363),
.B(n_305),
.Y(n_421)
);

AND2x2_ASAP7_75t_L g422 ( 
.A(n_365),
.B(n_315),
.Y(n_422)
);

INVx1_ASAP7_75t_L g423 ( 
.A(n_339),
.Y(n_423)
);

INVx1_ASAP7_75t_L g424 ( 
.A(n_354),
.Y(n_424)
);

INVx3_ASAP7_75t_L g425 ( 
.A(n_354),
.Y(n_425)
);

INVx1_ASAP7_75t_L g426 ( 
.A(n_355),
.Y(n_426)
);

INVx2_ASAP7_75t_SL g427 ( 
.A(n_351),
.Y(n_427)
);

INVx2_ASAP7_75t_L g428 ( 
.A(n_346),
.Y(n_428)
);

INVx1_ASAP7_75t_L g429 ( 
.A(n_355),
.Y(n_429)
);

AND2x2_ASAP7_75t_L g430 ( 
.A(n_395),
.B(n_316),
.Y(n_430)
);

NAND2xp5_ASAP7_75t_SL g431 ( 
.A(n_392),
.B(n_190),
.Y(n_431)
);

AO22x1_ASAP7_75t_L g432 ( 
.A1(n_418),
.A2(n_316),
.B1(n_319),
.B2(n_320),
.Y(n_432)
);

INVx1_ASAP7_75t_L g433 ( 
.A(n_347),
.Y(n_433)
);

INVx2_ASAP7_75t_L g434 ( 
.A(n_352),
.Y(n_434)
);

INVx4_ASAP7_75t_L g435 ( 
.A(n_417),
.Y(n_435)
);

CKINVDCx20_ASAP7_75t_R g436 ( 
.A(n_340),
.Y(n_436)
);

NAND2xp5_ASAP7_75t_L g437 ( 
.A(n_363),
.B(n_367),
.Y(n_437)
);

BUFx3_ASAP7_75t_L g438 ( 
.A(n_351),
.Y(n_438)
);

NAND2xp5_ASAP7_75t_L g439 ( 
.A(n_367),
.B(n_195),
.Y(n_439)
);

CKINVDCx5p33_ASAP7_75t_R g440 ( 
.A(n_361),
.Y(n_440)
);

NAND2xp5_ASAP7_75t_L g441 ( 
.A(n_382),
.B(n_198),
.Y(n_441)
);

CKINVDCx20_ASAP7_75t_R g442 ( 
.A(n_364),
.Y(n_442)
);

INVx2_ASAP7_75t_L g443 ( 
.A(n_353),
.Y(n_443)
);

NAND2xp5_ASAP7_75t_L g444 ( 
.A(n_382),
.B(n_199),
.Y(n_444)
);

INVx1_ASAP7_75t_L g445 ( 
.A(n_408),
.Y(n_445)
);

BUFx6f_ASAP7_75t_L g446 ( 
.A(n_360),
.Y(n_446)
);

INVx1_ASAP7_75t_L g447 ( 
.A(n_408),
.Y(n_447)
);

HB1xp67_ASAP7_75t_L g448 ( 
.A(n_402),
.Y(n_448)
);

INVx2_ASAP7_75t_L g449 ( 
.A(n_360),
.Y(n_449)
);

INVx2_ASAP7_75t_L g450 ( 
.A(n_356),
.Y(n_450)
);

OAI22xp5_ASAP7_75t_SL g451 ( 
.A1(n_393),
.A2(n_246),
.B1(n_233),
.B2(n_193),
.Y(n_451)
);

OAI22xp5_ASAP7_75t_L g452 ( 
.A1(n_391),
.A2(n_246),
.B1(n_233),
.B2(n_193),
.Y(n_452)
);

NAND2xp5_ASAP7_75t_L g453 ( 
.A(n_417),
.B(n_208),
.Y(n_453)
);

CKINVDCx5p33_ASAP7_75t_R g454 ( 
.A(n_350),
.Y(n_454)
);

INVx4_ASAP7_75t_L g455 ( 
.A(n_392),
.Y(n_455)
);

INVx2_ASAP7_75t_L g456 ( 
.A(n_356),
.Y(n_456)
);

CKINVDCx5p33_ASAP7_75t_R g457 ( 
.A(n_350),
.Y(n_457)
);

INVx1_ASAP7_75t_L g458 ( 
.A(n_410),
.Y(n_458)
);

INVx1_ASAP7_75t_L g459 ( 
.A(n_410),
.Y(n_459)
);

INVx3_ASAP7_75t_L g460 ( 
.A(n_358),
.Y(n_460)
);

INVx2_ASAP7_75t_L g461 ( 
.A(n_358),
.Y(n_461)
);

INVx1_ASAP7_75t_L g462 ( 
.A(n_411),
.Y(n_462)
);

OAI22xp5_ASAP7_75t_SL g463 ( 
.A1(n_415),
.A2(n_271),
.B1(n_322),
.B2(n_243),
.Y(n_463)
);

INVx1_ASAP7_75t_L g464 ( 
.A(n_411),
.Y(n_464)
);

INVx4_ASAP7_75t_L g465 ( 
.A(n_398),
.Y(n_465)
);

INVx2_ASAP7_75t_L g466 ( 
.A(n_359),
.Y(n_466)
);

BUFx6f_ASAP7_75t_L g467 ( 
.A(n_359),
.Y(n_467)
);

NOR2xp33_ASAP7_75t_L g468 ( 
.A(n_398),
.B(n_248),
.Y(n_468)
);

INVx2_ASAP7_75t_L g469 ( 
.A(n_413),
.Y(n_469)
);

INVx2_ASAP7_75t_L g470 ( 
.A(n_413),
.Y(n_470)
);

INVx1_ASAP7_75t_L g471 ( 
.A(n_366),
.Y(n_471)
);

BUFx3_ASAP7_75t_L g472 ( 
.A(n_337),
.Y(n_472)
);

AND2x6_ASAP7_75t_L g473 ( 
.A(n_342),
.B(n_169),
.Y(n_473)
);

BUFx6f_ASAP7_75t_L g474 ( 
.A(n_366),
.Y(n_474)
);

AND2x2_ASAP7_75t_L g475 ( 
.A(n_344),
.B(n_319),
.Y(n_475)
);

OAI22xp5_ASAP7_75t_L g476 ( 
.A1(n_349),
.A2(n_271),
.B1(n_322),
.B2(n_243),
.Y(n_476)
);

INVx1_ASAP7_75t_L g477 ( 
.A(n_406),
.Y(n_477)
);

INVx3_ASAP7_75t_L g478 ( 
.A(n_406),
.Y(n_478)
);

INVx2_ASAP7_75t_L g479 ( 
.A(n_368),
.Y(n_479)
);

INVx2_ASAP7_75t_L g480 ( 
.A(n_369),
.Y(n_480)
);

AND2x2_ASAP7_75t_L g481 ( 
.A(n_345),
.B(n_320),
.Y(n_481)
);

NOR2x1_ASAP7_75t_L g482 ( 
.A(n_370),
.B(n_181),
.Y(n_482)
);

HB1xp67_ASAP7_75t_L g483 ( 
.A(n_373),
.Y(n_483)
);

INVx1_ASAP7_75t_L g484 ( 
.A(n_372),
.Y(n_484)
);

INVx2_ASAP7_75t_L g485 ( 
.A(n_374),
.Y(n_485)
);

AND2x2_ASAP7_75t_L g486 ( 
.A(n_401),
.B(n_323),
.Y(n_486)
);

INVx1_ASAP7_75t_L g487 ( 
.A(n_376),
.Y(n_487)
);

BUFx6f_ASAP7_75t_L g488 ( 
.A(n_380),
.Y(n_488)
);

CKINVDCx8_ASAP7_75t_R g489 ( 
.A(n_362),
.Y(n_489)
);

AOI22xp5_ASAP7_75t_L g490 ( 
.A1(n_349),
.A2(n_272),
.B1(n_194),
.B2(n_225),
.Y(n_490)
);

INVx1_ASAP7_75t_L g491 ( 
.A(n_381),
.Y(n_491)
);

INVx1_ASAP7_75t_L g492 ( 
.A(n_383),
.Y(n_492)
);

INVx2_ASAP7_75t_L g493 ( 
.A(n_428),
.Y(n_493)
);

INVx1_ASAP7_75t_L g494 ( 
.A(n_428),
.Y(n_494)
);

INVx1_ASAP7_75t_L g495 ( 
.A(n_428),
.Y(n_495)
);

INVx1_ASAP7_75t_L g496 ( 
.A(n_434),
.Y(n_496)
);

NAND2xp5_ASAP7_75t_SL g497 ( 
.A(n_455),
.B(n_400),
.Y(n_497)
);

INVx2_ASAP7_75t_L g498 ( 
.A(n_434),
.Y(n_498)
);

AND3x2_ASAP7_75t_L g499 ( 
.A(n_483),
.B(n_404),
.C(n_412),
.Y(n_499)
);

NAND2xp5_ASAP7_75t_SL g500 ( 
.A(n_455),
.B(n_465),
.Y(n_500)
);

NAND2xp33_ASAP7_75t_L g501 ( 
.A(n_425),
.B(n_416),
.Y(n_501)
);

BUFx8_ASAP7_75t_SL g502 ( 
.A(n_436),
.Y(n_502)
);

BUFx6f_ASAP7_75t_SL g503 ( 
.A(n_455),
.Y(n_503)
);

AO22x2_ASAP7_75t_L g504 ( 
.A1(n_452),
.A2(n_362),
.B1(n_329),
.B2(n_307),
.Y(n_504)
);

BUFx3_ASAP7_75t_L g505 ( 
.A(n_438),
.Y(n_505)
);

INVx1_ASAP7_75t_L g506 ( 
.A(n_434),
.Y(n_506)
);

NAND2xp5_ASAP7_75t_SL g507 ( 
.A(n_455),
.B(n_400),
.Y(n_507)
);

HB1xp67_ASAP7_75t_L g508 ( 
.A(n_483),
.Y(n_508)
);

INVx2_ASAP7_75t_L g509 ( 
.A(n_443),
.Y(n_509)
);

INVx5_ASAP7_75t_L g510 ( 
.A(n_473),
.Y(n_510)
);

INVx2_ASAP7_75t_L g511 ( 
.A(n_443),
.Y(n_511)
);

INVx2_ASAP7_75t_L g512 ( 
.A(n_443),
.Y(n_512)
);

BUFx6f_ASAP7_75t_L g513 ( 
.A(n_474),
.Y(n_513)
);

INVx1_ASAP7_75t_L g514 ( 
.A(n_420),
.Y(n_514)
);

CKINVDCx5p33_ASAP7_75t_R g515 ( 
.A(n_454),
.Y(n_515)
);

NAND2xp33_ASAP7_75t_SL g516 ( 
.A(n_465),
.B(n_407),
.Y(n_516)
);

NAND2xp33_ASAP7_75t_L g517 ( 
.A(n_425),
.B(n_407),
.Y(n_517)
);

NOR2xp33_ASAP7_75t_L g518 ( 
.A(n_431),
.B(n_343),
.Y(n_518)
);

INVx2_ASAP7_75t_L g519 ( 
.A(n_425),
.Y(n_519)
);

NAND2xp5_ASAP7_75t_L g520 ( 
.A(n_427),
.B(n_468),
.Y(n_520)
);

BUFx10_ASAP7_75t_L g521 ( 
.A(n_440),
.Y(n_521)
);

INVx2_ASAP7_75t_L g522 ( 
.A(n_425),
.Y(n_522)
);

NAND2xp5_ASAP7_75t_L g523 ( 
.A(n_427),
.B(n_409),
.Y(n_523)
);

BUFx6f_ASAP7_75t_L g524 ( 
.A(n_474),
.Y(n_524)
);

NAND2xp5_ASAP7_75t_L g525 ( 
.A(n_427),
.B(n_409),
.Y(n_525)
);

BUFx3_ASAP7_75t_L g526 ( 
.A(n_438),
.Y(n_526)
);

NOR2xp33_ASAP7_75t_L g527 ( 
.A(n_465),
.B(n_348),
.Y(n_527)
);

INVx1_ASAP7_75t_L g528 ( 
.A(n_420),
.Y(n_528)
);

INVx1_ASAP7_75t_L g529 ( 
.A(n_423),
.Y(n_529)
);

NOR2xp67_ASAP7_75t_L g530 ( 
.A(n_465),
.B(n_307),
.Y(n_530)
);

INVx2_ASAP7_75t_L g531 ( 
.A(n_423),
.Y(n_531)
);

NAND2xp5_ASAP7_75t_SL g532 ( 
.A(n_489),
.B(n_414),
.Y(n_532)
);

INVx3_ASAP7_75t_L g533 ( 
.A(n_474),
.Y(n_533)
);

INVx1_ASAP7_75t_L g534 ( 
.A(n_424),
.Y(n_534)
);

INVx2_ASAP7_75t_L g535 ( 
.A(n_424),
.Y(n_535)
);

AOI22xp33_ASAP7_75t_L g536 ( 
.A1(n_435),
.A2(n_371),
.B1(n_338),
.B2(n_341),
.Y(n_536)
);

BUFx3_ASAP7_75t_L g537 ( 
.A(n_438),
.Y(n_537)
);

INVx4_ASAP7_75t_SL g538 ( 
.A(n_473),
.Y(n_538)
);

INVx2_ASAP7_75t_SL g539 ( 
.A(n_422),
.Y(n_539)
);

INVx3_ASAP7_75t_L g540 ( 
.A(n_474),
.Y(n_540)
);

AND2x6_ASAP7_75t_L g541 ( 
.A(n_482),
.B(n_169),
.Y(n_541)
);

NOR2xp33_ASAP7_75t_L g542 ( 
.A(n_435),
.B(n_348),
.Y(n_542)
);

INVx4_ASAP7_75t_L g543 ( 
.A(n_435),
.Y(n_543)
);

INVx2_ASAP7_75t_L g544 ( 
.A(n_426),
.Y(n_544)
);

INVx1_ASAP7_75t_L g545 ( 
.A(n_426),
.Y(n_545)
);

BUFx6f_ASAP7_75t_SL g546 ( 
.A(n_472),
.Y(n_546)
);

AND2x4_ASAP7_75t_L g547 ( 
.A(n_482),
.B(n_384),
.Y(n_547)
);

INVx1_ASAP7_75t_L g548 ( 
.A(n_429),
.Y(n_548)
);

NAND2xp5_ASAP7_75t_L g549 ( 
.A(n_433),
.B(n_414),
.Y(n_549)
);

BUFx6f_ASAP7_75t_L g550 ( 
.A(n_474),
.Y(n_550)
);

AOI22xp33_ASAP7_75t_L g551 ( 
.A1(n_435),
.A2(n_341),
.B1(n_405),
.B2(n_403),
.Y(n_551)
);

BUFx6f_ASAP7_75t_L g552 ( 
.A(n_474),
.Y(n_552)
);

NAND2xp5_ASAP7_75t_SL g553 ( 
.A(n_489),
.B(n_416),
.Y(n_553)
);

BUFx3_ASAP7_75t_L g554 ( 
.A(n_429),
.Y(n_554)
);

INVx2_ASAP7_75t_L g555 ( 
.A(n_460),
.Y(n_555)
);

INVx2_ASAP7_75t_L g556 ( 
.A(n_460),
.Y(n_556)
);

NOR3xp33_ASAP7_75t_L g557 ( 
.A(n_432),
.B(n_385),
.C(n_377),
.Y(n_557)
);

INVx1_ASAP7_75t_L g558 ( 
.A(n_433),
.Y(n_558)
);

INVx2_ASAP7_75t_L g559 ( 
.A(n_460),
.Y(n_559)
);

NAND3xp33_ASAP7_75t_L g560 ( 
.A(n_432),
.B(n_323),
.C(n_179),
.Y(n_560)
);

BUFx3_ASAP7_75t_L g561 ( 
.A(n_472),
.Y(n_561)
);

CKINVDCx20_ASAP7_75t_R g562 ( 
.A(n_442),
.Y(n_562)
);

INVx2_ASAP7_75t_SL g563 ( 
.A(n_422),
.Y(n_563)
);

NAND2xp5_ASAP7_75t_L g564 ( 
.A(n_475),
.B(n_341),
.Y(n_564)
);

INVx2_ASAP7_75t_L g565 ( 
.A(n_460),
.Y(n_565)
);

BUFx3_ASAP7_75t_L g566 ( 
.A(n_472),
.Y(n_566)
);

INVx3_ASAP7_75t_L g567 ( 
.A(n_474),
.Y(n_567)
);

INVx3_ASAP7_75t_L g568 ( 
.A(n_446),
.Y(n_568)
);

INVx1_ASAP7_75t_L g569 ( 
.A(n_469),
.Y(n_569)
);

NOR2xp67_ASAP7_75t_L g570 ( 
.A(n_448),
.B(n_386),
.Y(n_570)
);

BUFx6f_ASAP7_75t_L g571 ( 
.A(n_488),
.Y(n_571)
);

BUFx6f_ASAP7_75t_L g572 ( 
.A(n_488),
.Y(n_572)
);

INVx2_ASAP7_75t_L g573 ( 
.A(n_450),
.Y(n_573)
);

INVx1_ASAP7_75t_L g574 ( 
.A(n_469),
.Y(n_574)
);

NAND2xp5_ASAP7_75t_SL g575 ( 
.A(n_489),
.B(n_192),
.Y(n_575)
);

HB1xp67_ASAP7_75t_L g576 ( 
.A(n_457),
.Y(n_576)
);

INVxp33_ASAP7_75t_L g577 ( 
.A(n_452),
.Y(n_577)
);

INVx3_ASAP7_75t_L g578 ( 
.A(n_446),
.Y(n_578)
);

INVx2_ASAP7_75t_L g579 ( 
.A(n_450),
.Y(n_579)
);

INVx1_ASAP7_75t_L g580 ( 
.A(n_469),
.Y(n_580)
);

INVx1_ASAP7_75t_L g581 ( 
.A(n_470),
.Y(n_581)
);

INVxp67_ASAP7_75t_SL g582 ( 
.A(n_437),
.Y(n_582)
);

INVx1_ASAP7_75t_L g583 ( 
.A(n_470),
.Y(n_583)
);

INVx3_ASAP7_75t_L g584 ( 
.A(n_446),
.Y(n_584)
);

INVx2_ASAP7_75t_L g585 ( 
.A(n_450),
.Y(n_585)
);

AND2x2_ASAP7_75t_L g586 ( 
.A(n_479),
.B(n_399),
.Y(n_586)
);

INVx2_ASAP7_75t_L g587 ( 
.A(n_456),
.Y(n_587)
);

INVx2_ASAP7_75t_L g588 ( 
.A(n_456),
.Y(n_588)
);

BUFx8_ASAP7_75t_SL g589 ( 
.A(n_419),
.Y(n_589)
);

NOR2xp33_ASAP7_75t_L g590 ( 
.A(n_430),
.B(n_394),
.Y(n_590)
);

AND2x2_ASAP7_75t_L g591 ( 
.A(n_479),
.B(n_480),
.Y(n_591)
);

NAND2xp5_ASAP7_75t_L g592 ( 
.A(n_475),
.B(n_396),
.Y(n_592)
);

NOR2xp33_ASAP7_75t_L g593 ( 
.A(n_430),
.B(n_397),
.Y(n_593)
);

NAND2xp5_ASAP7_75t_SL g594 ( 
.A(n_481),
.B(n_192),
.Y(n_594)
);

INVx3_ASAP7_75t_L g595 ( 
.A(n_446),
.Y(n_595)
);

INVx1_ASAP7_75t_L g596 ( 
.A(n_470),
.Y(n_596)
);

INVx1_ASAP7_75t_L g597 ( 
.A(n_445),
.Y(n_597)
);

INVx2_ASAP7_75t_L g598 ( 
.A(n_456),
.Y(n_598)
);

INVx1_ASAP7_75t_L g599 ( 
.A(n_445),
.Y(n_599)
);

INVx2_ASAP7_75t_SL g600 ( 
.A(n_486),
.Y(n_600)
);

INVx2_ASAP7_75t_L g601 ( 
.A(n_461),
.Y(n_601)
);

CKINVDCx5p33_ASAP7_75t_R g602 ( 
.A(n_419),
.Y(n_602)
);

INVxp67_ASAP7_75t_L g603 ( 
.A(n_448),
.Y(n_603)
);

INVx2_ASAP7_75t_L g604 ( 
.A(n_461),
.Y(n_604)
);

AOI22xp5_ASAP7_75t_L g605 ( 
.A1(n_481),
.A2(n_238),
.B1(n_331),
.B2(n_328),
.Y(n_605)
);

INVxp33_ASAP7_75t_L g606 ( 
.A(n_476),
.Y(n_606)
);

BUFx10_ASAP7_75t_L g607 ( 
.A(n_484),
.Y(n_607)
);

INVx1_ASAP7_75t_L g608 ( 
.A(n_447),
.Y(n_608)
);

INVx1_ASAP7_75t_L g609 ( 
.A(n_447),
.Y(n_609)
);

AOI21x1_ASAP7_75t_L g610 ( 
.A1(n_453),
.A2(n_219),
.B(n_210),
.Y(n_610)
);

NAND2xp5_ASAP7_75t_SL g611 ( 
.A(n_486),
.B(n_312),
.Y(n_611)
);

INVx2_ASAP7_75t_L g612 ( 
.A(n_461),
.Y(n_612)
);

INVx1_ASAP7_75t_L g613 ( 
.A(n_458),
.Y(n_613)
);

NAND2xp5_ASAP7_75t_SL g614 ( 
.A(n_488),
.B(n_312),
.Y(n_614)
);

INVx2_ASAP7_75t_L g615 ( 
.A(n_466),
.Y(n_615)
);

INVx5_ASAP7_75t_L g616 ( 
.A(n_473),
.Y(n_616)
);

NOR2xp33_ASAP7_75t_L g617 ( 
.A(n_421),
.B(n_437),
.Y(n_617)
);

OR2x6_ASAP7_75t_L g618 ( 
.A(n_479),
.B(n_223),
.Y(n_618)
);

INVx2_ASAP7_75t_L g619 ( 
.A(n_466),
.Y(n_619)
);

NOR2x1p5_ASAP7_75t_L g620 ( 
.A(n_484),
.B(n_357),
.Y(n_620)
);

NOR2xp33_ASAP7_75t_L g621 ( 
.A(n_421),
.B(n_357),
.Y(n_621)
);

AND2x2_ASAP7_75t_L g622 ( 
.A(n_480),
.B(n_377),
.Y(n_622)
);

INVx2_ASAP7_75t_SL g623 ( 
.A(n_487),
.Y(n_623)
);

INVx2_ASAP7_75t_L g624 ( 
.A(n_466),
.Y(n_624)
);

INVx1_ASAP7_75t_L g625 ( 
.A(n_458),
.Y(n_625)
);

NAND2xp5_ASAP7_75t_L g626 ( 
.A(n_487),
.B(n_197),
.Y(n_626)
);

NAND2xp5_ASAP7_75t_SL g627 ( 
.A(n_488),
.B(n_317),
.Y(n_627)
);

INVx2_ASAP7_75t_L g628 ( 
.A(n_449),
.Y(n_628)
);

INVx2_ASAP7_75t_L g629 ( 
.A(n_449),
.Y(n_629)
);

INVx1_ASAP7_75t_L g630 ( 
.A(n_459),
.Y(n_630)
);

AND2x2_ASAP7_75t_L g631 ( 
.A(n_480),
.B(n_378),
.Y(n_631)
);

INVx2_ASAP7_75t_L g632 ( 
.A(n_449),
.Y(n_632)
);

NAND2xp5_ASAP7_75t_L g633 ( 
.A(n_491),
.B(n_213),
.Y(n_633)
);

INVx1_ASAP7_75t_L g634 ( 
.A(n_459),
.Y(n_634)
);

INVx1_ASAP7_75t_L g635 ( 
.A(n_462),
.Y(n_635)
);

INVx1_ASAP7_75t_L g636 ( 
.A(n_462),
.Y(n_636)
);

BUFx2_ASAP7_75t_L g637 ( 
.A(n_490),
.Y(n_637)
);

INVx1_ASAP7_75t_L g638 ( 
.A(n_464),
.Y(n_638)
);

INVx2_ASAP7_75t_L g639 ( 
.A(n_467),
.Y(n_639)
);

BUFx2_ASAP7_75t_L g640 ( 
.A(n_490),
.Y(n_640)
);

NAND2xp5_ASAP7_75t_L g641 ( 
.A(n_491),
.B(n_302),
.Y(n_641)
);

INVx2_ASAP7_75t_L g642 ( 
.A(n_467),
.Y(n_642)
);

INVx2_ASAP7_75t_L g643 ( 
.A(n_467),
.Y(n_643)
);

INVx2_ASAP7_75t_L g644 ( 
.A(n_493),
.Y(n_644)
);

O2A1O1Ixp5_ASAP7_75t_L g645 ( 
.A1(n_614),
.A2(n_492),
.B(n_478),
.C(n_485),
.Y(n_645)
);

AOI22xp33_ASAP7_75t_L g646 ( 
.A1(n_637),
.A2(n_488),
.B1(n_476),
.B2(n_485),
.Y(n_646)
);

INVx2_ASAP7_75t_L g647 ( 
.A(n_493),
.Y(n_647)
);

NAND2xp5_ASAP7_75t_SL g648 ( 
.A(n_607),
.B(n_488),
.Y(n_648)
);

NOR2xp33_ASAP7_75t_L g649 ( 
.A(n_520),
.B(n_492),
.Y(n_649)
);

INVx2_ASAP7_75t_SL g650 ( 
.A(n_508),
.Y(n_650)
);

INVx1_ASAP7_75t_L g651 ( 
.A(n_558),
.Y(n_651)
);

NOR2xp33_ASAP7_75t_L g652 ( 
.A(n_549),
.B(n_488),
.Y(n_652)
);

NOR2xp33_ASAP7_75t_L g653 ( 
.A(n_539),
.B(n_439),
.Y(n_653)
);

AND2x2_ASAP7_75t_L g654 ( 
.A(n_621),
.B(n_378),
.Y(n_654)
);

INVx1_ASAP7_75t_L g655 ( 
.A(n_558),
.Y(n_655)
);

AO22x2_ASAP7_75t_L g656 ( 
.A1(n_504),
.A2(n_451),
.B1(n_463),
.B2(n_389),
.Y(n_656)
);

AOI22xp5_ASAP7_75t_L g657 ( 
.A1(n_539),
.A2(n_485),
.B1(n_284),
.B2(n_390),
.Y(n_657)
);

A2O1A1Ixp33_ASAP7_75t_L g658 ( 
.A1(n_590),
.A2(n_464),
.B(n_478),
.C(n_453),
.Y(n_658)
);

NAND2xp5_ASAP7_75t_L g659 ( 
.A(n_617),
.B(n_478),
.Y(n_659)
);

NOR2xp33_ASAP7_75t_L g660 ( 
.A(n_563),
.B(n_439),
.Y(n_660)
);

NAND2xp5_ASAP7_75t_L g661 ( 
.A(n_623),
.B(n_478),
.Y(n_661)
);

INVx1_ASAP7_75t_L g662 ( 
.A(n_554),
.Y(n_662)
);

NAND2xp5_ASAP7_75t_L g663 ( 
.A(n_623),
.B(n_441),
.Y(n_663)
);

NAND2xp5_ASAP7_75t_L g664 ( 
.A(n_582),
.B(n_441),
.Y(n_664)
);

INVxp67_ASAP7_75t_L g665 ( 
.A(n_502),
.Y(n_665)
);

NOR2xp33_ASAP7_75t_L g666 ( 
.A(n_563),
.B(n_444),
.Y(n_666)
);

NAND2xp5_ASAP7_75t_L g667 ( 
.A(n_593),
.B(n_547),
.Y(n_667)
);

OAI22xp5_ASAP7_75t_L g668 ( 
.A1(n_600),
.A2(n_295),
.B1(n_200),
.B2(n_201),
.Y(n_668)
);

INVx1_ASAP7_75t_L g669 ( 
.A(n_554),
.Y(n_669)
);

INVx1_ASAP7_75t_L g670 ( 
.A(n_514),
.Y(n_670)
);

O2A1O1Ixp5_ASAP7_75t_L g671 ( 
.A1(n_627),
.A2(n_477),
.B(n_471),
.C(n_444),
.Y(n_671)
);

NAND2xp5_ASAP7_75t_L g672 ( 
.A(n_547),
.B(n_471),
.Y(n_672)
);

NAND2xp5_ASAP7_75t_L g673 ( 
.A(n_547),
.B(n_477),
.Y(n_673)
);

NOR2xp33_ASAP7_75t_L g674 ( 
.A(n_600),
.B(n_178),
.Y(n_674)
);

INVx2_ASAP7_75t_L g675 ( 
.A(n_498),
.Y(n_675)
);

INVxp33_ASAP7_75t_L g676 ( 
.A(n_589),
.Y(n_676)
);

NOR2xp33_ASAP7_75t_L g677 ( 
.A(n_532),
.B(n_553),
.Y(n_677)
);

INVx1_ASAP7_75t_L g678 ( 
.A(n_514),
.Y(n_678)
);

NAND3xp33_ASAP7_75t_L g679 ( 
.A(n_501),
.B(n_379),
.C(n_387),
.Y(n_679)
);

NAND2xp5_ASAP7_75t_SL g680 ( 
.A(n_607),
.B(n_379),
.Y(n_680)
);

OAI221xp5_ASAP7_75t_L g681 ( 
.A1(n_560),
.A2(n_605),
.B1(n_592),
.B2(n_551),
.C(n_564),
.Y(n_681)
);

NAND2xp5_ASAP7_75t_L g682 ( 
.A(n_527),
.B(n_317),
.Y(n_682)
);

INVxp67_ASAP7_75t_L g683 ( 
.A(n_576),
.Y(n_683)
);

NAND2xp5_ASAP7_75t_SL g684 ( 
.A(n_607),
.B(n_387),
.Y(n_684)
);

INVx1_ASAP7_75t_L g685 ( 
.A(n_528),
.Y(n_685)
);

AOI22xp33_ASAP7_75t_L g686 ( 
.A1(n_637),
.A2(n_388),
.B1(n_390),
.B2(n_463),
.Y(n_686)
);

NAND2xp5_ASAP7_75t_SL g687 ( 
.A(n_530),
.B(n_325),
.Y(n_687)
);

NAND2x1_ASAP7_75t_L g688 ( 
.A(n_543),
.B(n_473),
.Y(n_688)
);

AOI21xp5_ASAP7_75t_L g689 ( 
.A1(n_528),
.A2(n_258),
.B(n_286),
.Y(n_689)
);

INVx1_ASAP7_75t_L g690 ( 
.A(n_529),
.Y(n_690)
);

NAND2xp5_ASAP7_75t_L g691 ( 
.A(n_591),
.B(n_325),
.Y(n_691)
);

INVx1_ASAP7_75t_L g692 ( 
.A(n_529),
.Y(n_692)
);

INVx2_ASAP7_75t_L g693 ( 
.A(n_498),
.Y(n_693)
);

NAND2xp5_ASAP7_75t_L g694 ( 
.A(n_591),
.B(n_326),
.Y(n_694)
);

NAND3xp33_ASAP7_75t_L g695 ( 
.A(n_501),
.B(n_388),
.C(n_266),
.Y(n_695)
);

AND2x2_ASAP7_75t_L g696 ( 
.A(n_622),
.B(n_375),
.Y(n_696)
);

NAND2xp5_ASAP7_75t_L g697 ( 
.A(n_626),
.B(n_326),
.Y(n_697)
);

NAND2xp5_ASAP7_75t_SL g698 ( 
.A(n_530),
.B(n_226),
.Y(n_698)
);

NAND2xp5_ASAP7_75t_L g699 ( 
.A(n_633),
.B(n_211),
.Y(n_699)
);

INVx2_ASAP7_75t_L g700 ( 
.A(n_509),
.Y(n_700)
);

INVx2_ASAP7_75t_L g701 ( 
.A(n_509),
.Y(n_701)
);

INVx2_ASAP7_75t_L g702 ( 
.A(n_511),
.Y(n_702)
);

BUFx2_ASAP7_75t_L g703 ( 
.A(n_562),
.Y(n_703)
);

BUFx12f_ASAP7_75t_SL g704 ( 
.A(n_622),
.Y(n_704)
);

AOI22xp5_ASAP7_75t_L g705 ( 
.A1(n_517),
.A2(n_232),
.B1(n_336),
.B2(n_335),
.Y(n_705)
);

INVxp67_ASAP7_75t_SL g706 ( 
.A(n_561),
.Y(n_706)
);

OAI22xp5_ASAP7_75t_L g707 ( 
.A1(n_523),
.A2(n_251),
.B1(n_265),
.B2(n_245),
.Y(n_707)
);

AND2x4_ASAP7_75t_L g708 ( 
.A(n_561),
.B(n_240),
.Y(n_708)
);

OAI22xp5_ASAP7_75t_SL g709 ( 
.A1(n_606),
.A2(n_451),
.B1(n_244),
.B2(n_254),
.Y(n_709)
);

NAND2xp5_ASAP7_75t_L g710 ( 
.A(n_641),
.B(n_215),
.Y(n_710)
);

NAND2xp5_ASAP7_75t_SL g711 ( 
.A(n_516),
.B(n_224),
.Y(n_711)
);

NAND2xp5_ASAP7_75t_L g712 ( 
.A(n_542),
.B(n_279),
.Y(n_712)
);

INVxp67_ASAP7_75t_L g713 ( 
.A(n_602),
.Y(n_713)
);

NAND2xp5_ASAP7_75t_L g714 ( 
.A(n_586),
.B(n_282),
.Y(n_714)
);

CKINVDCx5p33_ASAP7_75t_R g715 ( 
.A(n_515),
.Y(n_715)
);

CKINVDCx5p33_ASAP7_75t_R g716 ( 
.A(n_515),
.Y(n_716)
);

O2A1O1Ixp33_ASAP7_75t_L g717 ( 
.A1(n_517),
.A2(n_314),
.B(n_242),
.C(n_250),
.Y(n_717)
);

NOR2xp33_ASAP7_75t_L g718 ( 
.A(n_525),
.B(n_288),
.Y(n_718)
);

NAND2xp5_ASAP7_75t_SL g719 ( 
.A(n_518),
.B(n_301),
.Y(n_719)
);

OAI22xp33_ASAP7_75t_L g720 ( 
.A1(n_577),
.A2(n_309),
.B1(n_306),
.B2(n_311),
.Y(n_720)
);

NOR2xp67_ASAP7_75t_SL g721 ( 
.A(n_500),
.B(n_170),
.Y(n_721)
);

INVx1_ASAP7_75t_L g722 ( 
.A(n_534),
.Y(n_722)
);

INVx2_ASAP7_75t_L g723 ( 
.A(n_511),
.Y(n_723)
);

NOR2xp33_ASAP7_75t_L g724 ( 
.A(n_611),
.B(n_241),
.Y(n_724)
);

NAND2xp5_ASAP7_75t_L g725 ( 
.A(n_586),
.B(n_175),
.Y(n_725)
);

NAND2xp5_ASAP7_75t_SL g726 ( 
.A(n_570),
.B(n_202),
.Y(n_726)
);

NAND2xp5_ASAP7_75t_L g727 ( 
.A(n_597),
.B(n_203),
.Y(n_727)
);

INVx2_ASAP7_75t_L g728 ( 
.A(n_512),
.Y(n_728)
);

INVx2_ASAP7_75t_L g729 ( 
.A(n_512),
.Y(n_729)
);

NAND2xp5_ASAP7_75t_L g730 ( 
.A(n_597),
.B(n_207),
.Y(n_730)
);

INVxp67_ASAP7_75t_L g731 ( 
.A(n_602),
.Y(n_731)
);

NAND2xp5_ASAP7_75t_SL g732 ( 
.A(n_536),
.B(n_216),
.Y(n_732)
);

NAND2xp5_ASAP7_75t_L g733 ( 
.A(n_599),
.B(n_217),
.Y(n_733)
);

AND2x2_ASAP7_75t_L g734 ( 
.A(n_631),
.B(n_467),
.Y(n_734)
);

INVx1_ASAP7_75t_L g735 ( 
.A(n_534),
.Y(n_735)
);

NAND2xp5_ASAP7_75t_L g736 ( 
.A(n_599),
.B(n_218),
.Y(n_736)
);

INVx8_ASAP7_75t_L g737 ( 
.A(n_503),
.Y(n_737)
);

OAI22xp33_ASAP7_75t_L g738 ( 
.A1(n_640),
.A2(n_274),
.B1(n_289),
.B2(n_256),
.Y(n_738)
);

INVx2_ASAP7_75t_L g739 ( 
.A(n_628),
.Y(n_739)
);

NOR2xp33_ASAP7_75t_L g740 ( 
.A(n_543),
.B(n_257),
.Y(n_740)
);

NOR2x1p5_ASAP7_75t_L g741 ( 
.A(n_631),
.B(n_521),
.Y(n_741)
);

NAND2xp5_ASAP7_75t_SL g742 ( 
.A(n_497),
.B(n_222),
.Y(n_742)
);

AOI22xp5_ASAP7_75t_L g743 ( 
.A1(n_503),
.A2(n_275),
.B1(n_277),
.B2(n_280),
.Y(n_743)
);

INVx1_ASAP7_75t_L g744 ( 
.A(n_545),
.Y(n_744)
);

NAND2xp5_ASAP7_75t_SL g745 ( 
.A(n_543),
.B(n_285),
.Y(n_745)
);

INVx1_ASAP7_75t_L g746 ( 
.A(n_545),
.Y(n_746)
);

NAND2xp5_ASAP7_75t_SL g747 ( 
.A(n_519),
.B(n_313),
.Y(n_747)
);

NAND2xp5_ASAP7_75t_L g748 ( 
.A(n_608),
.B(n_227),
.Y(n_748)
);

NAND2xp5_ASAP7_75t_L g749 ( 
.A(n_608),
.B(n_228),
.Y(n_749)
);

INVx2_ASAP7_75t_L g750 ( 
.A(n_628),
.Y(n_750)
);

INVx2_ASAP7_75t_L g751 ( 
.A(n_629),
.Y(n_751)
);

HB1xp67_ASAP7_75t_L g752 ( 
.A(n_603),
.Y(n_752)
);

NAND2xp5_ASAP7_75t_SL g753 ( 
.A(n_507),
.B(n_234),
.Y(n_753)
);

AOI22xp33_ASAP7_75t_L g754 ( 
.A1(n_640),
.A2(n_473),
.B1(n_446),
.B2(n_467),
.Y(n_754)
);

AND2x2_ASAP7_75t_L g755 ( 
.A(n_521),
.B(n_467),
.Y(n_755)
);

NOR2xp33_ASAP7_75t_L g756 ( 
.A(n_594),
.B(n_0),
.Y(n_756)
);

INVx2_ASAP7_75t_L g757 ( 
.A(n_629),
.Y(n_757)
);

NAND2xp5_ASAP7_75t_L g758 ( 
.A(n_609),
.B(n_236),
.Y(n_758)
);

BUFx3_ASAP7_75t_L g759 ( 
.A(n_505),
.Y(n_759)
);

INVxp67_ASAP7_75t_L g760 ( 
.A(n_521),
.Y(n_760)
);

NOR2xp33_ASAP7_75t_L g761 ( 
.A(n_566),
.B(n_0),
.Y(n_761)
);

INVx1_ASAP7_75t_L g762 ( 
.A(n_548),
.Y(n_762)
);

INVx2_ASAP7_75t_L g763 ( 
.A(n_632),
.Y(n_763)
);

OAI22xp33_ASAP7_75t_L g764 ( 
.A1(n_618),
.A2(n_467),
.B1(n_237),
.B2(n_247),
.Y(n_764)
);

NAND2xp5_ASAP7_75t_L g765 ( 
.A(n_609),
.B(n_269),
.Y(n_765)
);

NOR2xp33_ASAP7_75t_L g766 ( 
.A(n_566),
.B(n_2),
.Y(n_766)
);

NAND2xp5_ASAP7_75t_L g767 ( 
.A(n_613),
.B(n_625),
.Y(n_767)
);

INVx1_ASAP7_75t_L g768 ( 
.A(n_548),
.Y(n_768)
);

NAND2xp33_ASAP7_75t_L g769 ( 
.A(n_519),
.B(n_473),
.Y(n_769)
);

NAND2xp5_ASAP7_75t_L g770 ( 
.A(n_613),
.B(n_263),
.Y(n_770)
);

NOR2xp33_ASAP7_75t_L g771 ( 
.A(n_575),
.B(n_2),
.Y(n_771)
);

INVx1_ASAP7_75t_L g772 ( 
.A(n_625),
.Y(n_772)
);

BUFx3_ASAP7_75t_L g773 ( 
.A(n_505),
.Y(n_773)
);

NAND2xp5_ASAP7_75t_SL g774 ( 
.A(n_557),
.B(n_300),
.Y(n_774)
);

BUFx6f_ASAP7_75t_L g775 ( 
.A(n_571),
.Y(n_775)
);

INVx1_ASAP7_75t_L g776 ( 
.A(n_630),
.Y(n_776)
);

NAND3xp33_ASAP7_75t_L g777 ( 
.A(n_630),
.B(n_308),
.C(n_253),
.Y(n_777)
);

NAND2xp5_ASAP7_75t_SL g778 ( 
.A(n_526),
.B(n_330),
.Y(n_778)
);

INVx1_ASAP7_75t_L g779 ( 
.A(n_634),
.Y(n_779)
);

NAND2xp5_ASAP7_75t_L g780 ( 
.A(n_634),
.B(n_262),
.Y(n_780)
);

INVx2_ASAP7_75t_L g781 ( 
.A(n_632),
.Y(n_781)
);

NAND2xp5_ASAP7_75t_SL g782 ( 
.A(n_526),
.B(n_537),
.Y(n_782)
);

BUFx6f_ASAP7_75t_L g783 ( 
.A(n_571),
.Y(n_783)
);

NAND2xp5_ASAP7_75t_SL g784 ( 
.A(n_537),
.B(n_333),
.Y(n_784)
);

AOI22xp33_ASAP7_75t_L g785 ( 
.A1(n_504),
.A2(n_618),
.B1(n_535),
.B2(n_544),
.Y(n_785)
);

A2O1A1Ixp33_ASAP7_75t_L g786 ( 
.A1(n_635),
.A2(n_291),
.B(n_255),
.C(n_259),
.Y(n_786)
);

NAND2xp5_ASAP7_75t_L g787 ( 
.A(n_635),
.B(n_261),
.Y(n_787)
);

NOR2xp33_ASAP7_75t_L g788 ( 
.A(n_546),
.B(n_8),
.Y(n_788)
);

INVx2_ASAP7_75t_L g789 ( 
.A(n_531),
.Y(n_789)
);

NAND2xp5_ASAP7_75t_L g790 ( 
.A(n_636),
.B(n_273),
.Y(n_790)
);

NOR2xp33_ASAP7_75t_L g791 ( 
.A(n_546),
.B(n_9),
.Y(n_791)
);

INVxp67_ASAP7_75t_L g792 ( 
.A(n_620),
.Y(n_792)
);

AND2x2_ASAP7_75t_L g793 ( 
.A(n_504),
.B(n_446),
.Y(n_793)
);

NOR2xp67_ASAP7_75t_L g794 ( 
.A(n_636),
.B(n_260),
.Y(n_794)
);

INVx2_ASAP7_75t_L g795 ( 
.A(n_531),
.Y(n_795)
);

NAND2xp5_ASAP7_75t_L g796 ( 
.A(n_638),
.B(n_278),
.Y(n_796)
);

AOI22xp5_ASAP7_75t_L g797 ( 
.A1(n_503),
.A2(n_290),
.B1(n_287),
.B2(n_281),
.Y(n_797)
);

NAND2xp33_ASAP7_75t_L g798 ( 
.A(n_522),
.B(n_473),
.Y(n_798)
);

HB1xp67_ASAP7_75t_L g799 ( 
.A(n_620),
.Y(n_799)
);

NAND2xp33_ASAP7_75t_L g800 ( 
.A(n_522),
.B(n_473),
.Y(n_800)
);

NAND2xp5_ASAP7_75t_SL g801 ( 
.A(n_638),
.B(n_169),
.Y(n_801)
);

AOI22xp33_ASAP7_75t_L g802 ( 
.A1(n_504),
.A2(n_473),
.B1(n_446),
.B2(n_252),
.Y(n_802)
);

NOR2xp67_ASAP7_75t_L g803 ( 
.A(n_569),
.B(n_88),
.Y(n_803)
);

INVx2_ASAP7_75t_L g804 ( 
.A(n_535),
.Y(n_804)
);

NAND2xp5_ASAP7_75t_SL g805 ( 
.A(n_513),
.B(n_252),
.Y(n_805)
);

NAND2xp5_ASAP7_75t_L g806 ( 
.A(n_544),
.B(n_252),
.Y(n_806)
);

NAND2xp5_ASAP7_75t_SL g807 ( 
.A(n_513),
.B(n_252),
.Y(n_807)
);

BUFx3_ASAP7_75t_L g808 ( 
.A(n_513),
.Y(n_808)
);

INVxp67_ASAP7_75t_SL g809 ( 
.A(n_513),
.Y(n_809)
);

INVx2_ASAP7_75t_L g810 ( 
.A(n_573),
.Y(n_810)
);

HB1xp67_ASAP7_75t_L g811 ( 
.A(n_618),
.Y(n_811)
);

INVx1_ASAP7_75t_L g812 ( 
.A(n_569),
.Y(n_812)
);

NAND2xp5_ASAP7_75t_SL g813 ( 
.A(n_513),
.B(n_524),
.Y(n_813)
);

INVx1_ASAP7_75t_L g814 ( 
.A(n_574),
.Y(n_814)
);

INVx2_ASAP7_75t_L g815 ( 
.A(n_573),
.Y(n_815)
);

INVx1_ASAP7_75t_L g816 ( 
.A(n_670),
.Y(n_816)
);

INVx2_ASAP7_75t_L g817 ( 
.A(n_739),
.Y(n_817)
);

NOR3xp33_ASAP7_75t_SL g818 ( 
.A(n_715),
.B(n_574),
.C(n_596),
.Y(n_818)
);

NAND2xp5_ASAP7_75t_L g819 ( 
.A(n_649),
.B(n_580),
.Y(n_819)
);

BUFx6f_ASAP7_75t_L g820 ( 
.A(n_775),
.Y(n_820)
);

AND2x2_ASAP7_75t_L g821 ( 
.A(n_654),
.B(n_499),
.Y(n_821)
);

NOR2x2_ASAP7_75t_L g822 ( 
.A(n_716),
.B(n_618),
.Y(n_822)
);

OAI22xp5_ASAP7_75t_SL g823 ( 
.A1(n_709),
.A2(n_580),
.B1(n_596),
.B2(n_583),
.Y(n_823)
);

HB1xp67_ASAP7_75t_L g824 ( 
.A(n_704),
.Y(n_824)
);

INVx2_ASAP7_75t_SL g825 ( 
.A(n_703),
.Y(n_825)
);

NAND2xp5_ASAP7_75t_L g826 ( 
.A(n_649),
.B(n_653),
.Y(n_826)
);

INVx1_ASAP7_75t_L g827 ( 
.A(n_678),
.Y(n_827)
);

AOI22xp5_ASAP7_75t_L g828 ( 
.A1(n_667),
.A2(n_546),
.B1(n_541),
.B2(n_555),
.Y(n_828)
);

NAND2xp5_ASAP7_75t_L g829 ( 
.A(n_653),
.B(n_581),
.Y(n_829)
);

AND2x4_ASAP7_75t_L g830 ( 
.A(n_741),
.B(n_538),
.Y(n_830)
);

BUFx3_ASAP7_75t_L g831 ( 
.A(n_650),
.Y(n_831)
);

AOI22xp33_ASAP7_75t_L g832 ( 
.A1(n_656),
.A2(n_495),
.B1(n_496),
.B2(n_506),
.Y(n_832)
);

NAND2xp5_ASAP7_75t_L g833 ( 
.A(n_660),
.B(n_581),
.Y(n_833)
);

AOI22xp5_ASAP7_75t_L g834 ( 
.A1(n_771),
.A2(n_541),
.B1(n_555),
.B2(n_556),
.Y(n_834)
);

INVx2_ASAP7_75t_L g835 ( 
.A(n_750),
.Y(n_835)
);

AND2x4_ASAP7_75t_L g836 ( 
.A(n_811),
.B(n_538),
.Y(n_836)
);

NAND2xp5_ASAP7_75t_L g837 ( 
.A(n_660),
.B(n_583),
.Y(n_837)
);

OR2x2_ASAP7_75t_SL g838 ( 
.A(n_679),
.B(n_556),
.Y(n_838)
);

INVx2_ASAP7_75t_SL g839 ( 
.A(n_696),
.Y(n_839)
);

INVx2_ASAP7_75t_L g840 ( 
.A(n_751),
.Y(n_840)
);

AOI22xp5_ASAP7_75t_L g841 ( 
.A1(n_771),
.A2(n_541),
.B1(n_565),
.B2(n_559),
.Y(n_841)
);

NAND2xp5_ASAP7_75t_L g842 ( 
.A(n_666),
.B(n_494),
.Y(n_842)
);

BUFx6f_ASAP7_75t_L g843 ( 
.A(n_775),
.Y(n_843)
);

INVx2_ASAP7_75t_L g844 ( 
.A(n_751),
.Y(n_844)
);

AOI22xp5_ASAP7_75t_SL g845 ( 
.A1(n_713),
.A2(n_541),
.B1(n_495),
.B2(n_496),
.Y(n_845)
);

INVx4_ASAP7_75t_L g846 ( 
.A(n_737),
.Y(n_846)
);

INVx1_ASAP7_75t_L g847 ( 
.A(n_685),
.Y(n_847)
);

INVx1_ASAP7_75t_L g848 ( 
.A(n_690),
.Y(n_848)
);

AOI21xp5_ASAP7_75t_L g849 ( 
.A1(n_659),
.A2(n_565),
.B(n_559),
.Y(n_849)
);

NOR2xp33_ASAP7_75t_L g850 ( 
.A(n_681),
.B(n_533),
.Y(n_850)
);

NAND2xp5_ASAP7_75t_L g851 ( 
.A(n_666),
.B(n_494),
.Y(n_851)
);

INVx2_ASAP7_75t_SL g852 ( 
.A(n_752),
.Y(n_852)
);

NOR2xp33_ASAP7_75t_SL g853 ( 
.A(n_665),
.B(n_510),
.Y(n_853)
);

NAND2xp5_ASAP7_75t_L g854 ( 
.A(n_663),
.B(n_506),
.Y(n_854)
);

NOR2xp33_ASAP7_75t_L g855 ( 
.A(n_677),
.B(n_533),
.Y(n_855)
);

NOR2xp67_ASAP7_75t_L g856 ( 
.A(n_760),
.B(n_610),
.Y(n_856)
);

BUFx6f_ASAP7_75t_L g857 ( 
.A(n_775),
.Y(n_857)
);

INVx3_ASAP7_75t_L g858 ( 
.A(n_759),
.Y(n_858)
);

INVx1_ASAP7_75t_L g859 ( 
.A(n_692),
.Y(n_859)
);

OR2x6_ASAP7_75t_L g860 ( 
.A(n_737),
.B(n_579),
.Y(n_860)
);

INVx2_ASAP7_75t_L g861 ( 
.A(n_757),
.Y(n_861)
);

NAND2xp5_ASAP7_75t_SL g862 ( 
.A(n_677),
.B(n_524),
.Y(n_862)
);

NAND2xp5_ASAP7_75t_L g863 ( 
.A(n_664),
.B(n_541),
.Y(n_863)
);

INVx2_ASAP7_75t_SL g864 ( 
.A(n_799),
.Y(n_864)
);

INVx2_ASAP7_75t_SL g865 ( 
.A(n_708),
.Y(n_865)
);

NAND2xp5_ASAP7_75t_L g866 ( 
.A(n_718),
.B(n_541),
.Y(n_866)
);

NAND2xp5_ASAP7_75t_L g867 ( 
.A(n_718),
.B(n_734),
.Y(n_867)
);

NAND2xp5_ASAP7_75t_SL g868 ( 
.A(n_775),
.B(n_524),
.Y(n_868)
);

NOR2xp33_ASAP7_75t_L g869 ( 
.A(n_680),
.B(n_533),
.Y(n_869)
);

INVx2_ASAP7_75t_L g870 ( 
.A(n_757),
.Y(n_870)
);

AOI22xp5_ASAP7_75t_L g871 ( 
.A1(n_756),
.A2(n_541),
.B1(n_567),
.B2(n_540),
.Y(n_871)
);

INVx5_ASAP7_75t_L g872 ( 
.A(n_737),
.Y(n_872)
);

INVx1_ASAP7_75t_L g873 ( 
.A(n_722),
.Y(n_873)
);

INVx2_ASAP7_75t_L g874 ( 
.A(n_763),
.Y(n_874)
);

BUFx6f_ASAP7_75t_L g875 ( 
.A(n_783),
.Y(n_875)
);

INVx2_ASAP7_75t_L g876 ( 
.A(n_763),
.Y(n_876)
);

INVx1_ASAP7_75t_L g877 ( 
.A(n_735),
.Y(n_877)
);

NAND2xp5_ASAP7_75t_L g878 ( 
.A(n_672),
.B(n_579),
.Y(n_878)
);

BUFx6f_ASAP7_75t_L g879 ( 
.A(n_783),
.Y(n_879)
);

AND2x4_ASAP7_75t_L g880 ( 
.A(n_792),
.B(n_538),
.Y(n_880)
);

NOR3xp33_ASAP7_75t_SL g881 ( 
.A(n_711),
.B(n_10),
.C(n_13),
.Y(n_881)
);

INVx1_ASAP7_75t_L g882 ( 
.A(n_744),
.Y(n_882)
);

NAND3xp33_ASAP7_75t_SL g883 ( 
.A(n_712),
.B(n_643),
.C(n_642),
.Y(n_883)
);

OR2x6_ASAP7_75t_L g884 ( 
.A(n_731),
.B(n_585),
.Y(n_884)
);

INVx3_ASAP7_75t_L g885 ( 
.A(n_759),
.Y(n_885)
);

INVx2_ASAP7_75t_L g886 ( 
.A(n_781),
.Y(n_886)
);

AND2x2_ASAP7_75t_L g887 ( 
.A(n_683),
.B(n_585),
.Y(n_887)
);

INVx2_ASAP7_75t_L g888 ( 
.A(n_781),
.Y(n_888)
);

INVx4_ASAP7_75t_L g889 ( 
.A(n_773),
.Y(n_889)
);

INVx1_ASAP7_75t_L g890 ( 
.A(n_746),
.Y(n_890)
);

INVx1_ASAP7_75t_L g891 ( 
.A(n_762),
.Y(n_891)
);

NAND2xp5_ASAP7_75t_L g892 ( 
.A(n_673),
.B(n_587),
.Y(n_892)
);

NOR2xp33_ASAP7_75t_L g893 ( 
.A(n_684),
.B(n_540),
.Y(n_893)
);

AOI22xp33_ASAP7_75t_L g894 ( 
.A1(n_656),
.A2(n_604),
.B1(n_601),
.B2(n_587),
.Y(n_894)
);

INVx2_ASAP7_75t_L g895 ( 
.A(n_810),
.Y(n_895)
);

OAI21xp5_ASAP7_75t_L g896 ( 
.A1(n_658),
.A2(n_540),
.B(n_567),
.Y(n_896)
);

NAND2xp5_ASAP7_75t_L g897 ( 
.A(n_651),
.B(n_619),
.Y(n_897)
);

NOR2x1p5_ASAP7_75t_L g898 ( 
.A(n_695),
.B(n_567),
.Y(n_898)
);

INVx3_ASAP7_75t_L g899 ( 
.A(n_773),
.Y(n_899)
);

INVx2_ASAP7_75t_L g900 ( 
.A(n_810),
.Y(n_900)
);

NAND2xp5_ASAP7_75t_L g901 ( 
.A(n_655),
.B(n_612),
.Y(n_901)
);

NAND2xp5_ASAP7_75t_SL g902 ( 
.A(n_682),
.B(n_550),
.Y(n_902)
);

INVx2_ASAP7_75t_L g903 ( 
.A(n_815),
.Y(n_903)
);

AND2x6_ASAP7_75t_SL g904 ( 
.A(n_756),
.B(n_10),
.Y(n_904)
);

INVx2_ASAP7_75t_SL g905 ( 
.A(n_708),
.Y(n_905)
);

INVx1_ASAP7_75t_L g906 ( 
.A(n_768),
.Y(n_906)
);

NAND2xp5_ASAP7_75t_L g907 ( 
.A(n_674),
.B(n_612),
.Y(n_907)
);

INVxp33_ASAP7_75t_L g908 ( 
.A(n_674),
.Y(n_908)
);

INVx1_ASAP7_75t_L g909 ( 
.A(n_772),
.Y(n_909)
);

CKINVDCx5p33_ASAP7_75t_R g910 ( 
.A(n_686),
.Y(n_910)
);

BUFx6f_ASAP7_75t_L g911 ( 
.A(n_783),
.Y(n_911)
);

INVx2_ASAP7_75t_L g912 ( 
.A(n_815),
.Y(n_912)
);

AOI22xp33_ASAP7_75t_L g913 ( 
.A1(n_656),
.A2(n_619),
.B1(n_601),
.B2(n_588),
.Y(n_913)
);

INVx1_ASAP7_75t_L g914 ( 
.A(n_776),
.Y(n_914)
);

INVx1_ASAP7_75t_L g915 ( 
.A(n_779),
.Y(n_915)
);

INVx3_ASAP7_75t_L g916 ( 
.A(n_808),
.Y(n_916)
);

BUFx3_ASAP7_75t_L g917 ( 
.A(n_708),
.Y(n_917)
);

AOI22xp5_ASAP7_75t_L g918 ( 
.A1(n_705),
.A2(n_572),
.B1(n_571),
.B2(n_550),
.Y(n_918)
);

NAND2xp5_ASAP7_75t_L g919 ( 
.A(n_646),
.B(n_588),
.Y(n_919)
);

INVx2_ASAP7_75t_SL g920 ( 
.A(n_755),
.Y(n_920)
);

NAND2xp5_ASAP7_75t_SL g921 ( 
.A(n_783),
.B(n_524),
.Y(n_921)
);

BUFx2_ASAP7_75t_L g922 ( 
.A(n_788),
.Y(n_922)
);

INVx1_ASAP7_75t_L g923 ( 
.A(n_812),
.Y(n_923)
);

NAND2xp5_ASAP7_75t_L g924 ( 
.A(n_697),
.B(n_615),
.Y(n_924)
);

NAND2xp5_ASAP7_75t_L g925 ( 
.A(n_714),
.B(n_615),
.Y(n_925)
);

INVxp67_ASAP7_75t_L g926 ( 
.A(n_761),
.Y(n_926)
);

INVx1_ASAP7_75t_SL g927 ( 
.A(n_793),
.Y(n_927)
);

INVx5_ASAP7_75t_L g928 ( 
.A(n_808),
.Y(n_928)
);

BUFx4f_ASAP7_75t_SL g929 ( 
.A(n_774),
.Y(n_929)
);

AND2x2_ASAP7_75t_L g930 ( 
.A(n_657),
.B(n_598),
.Y(n_930)
);

AOI22xp33_ASAP7_75t_L g931 ( 
.A1(n_785),
.A2(n_598),
.B1(n_624),
.B2(n_604),
.Y(n_931)
);

BUFx6f_ASAP7_75t_L g932 ( 
.A(n_688),
.Y(n_932)
);

NAND2xp5_ASAP7_75t_SL g933 ( 
.A(n_767),
.B(n_789),
.Y(n_933)
);

INVx4_ASAP7_75t_L g934 ( 
.A(n_789),
.Y(n_934)
);

NAND2xp5_ASAP7_75t_SL g935 ( 
.A(n_795),
.B(n_524),
.Y(n_935)
);

INVx1_ASAP7_75t_L g936 ( 
.A(n_814),
.Y(n_936)
);

OR2x6_ASAP7_75t_L g937 ( 
.A(n_662),
.B(n_624),
.Y(n_937)
);

INVx1_ASAP7_75t_L g938 ( 
.A(n_795),
.Y(n_938)
);

NAND2xp5_ASAP7_75t_SL g939 ( 
.A(n_788),
.B(n_550),
.Y(n_939)
);

INVx2_ASAP7_75t_L g940 ( 
.A(n_644),
.Y(n_940)
);

INVx2_ASAP7_75t_SL g941 ( 
.A(n_791),
.Y(n_941)
);

INVx1_ASAP7_75t_L g942 ( 
.A(n_804),
.Y(n_942)
);

NAND2xp5_ASAP7_75t_SL g943 ( 
.A(n_804),
.B(n_550),
.Y(n_943)
);

NOR3xp33_ASAP7_75t_SL g944 ( 
.A(n_742),
.B(n_16),
.C(n_19),
.Y(n_944)
);

INVx2_ASAP7_75t_L g945 ( 
.A(n_644),
.Y(n_945)
);

NAND2xp5_ASAP7_75t_SL g946 ( 
.A(n_791),
.B(n_550),
.Y(n_946)
);

INVx1_ASAP7_75t_L g947 ( 
.A(n_669),
.Y(n_947)
);

NAND2xp5_ASAP7_75t_L g948 ( 
.A(n_691),
.B(n_552),
.Y(n_948)
);

BUFx6f_ASAP7_75t_L g949 ( 
.A(n_647),
.Y(n_949)
);

AND2x6_ASAP7_75t_L g950 ( 
.A(n_761),
.B(n_571),
.Y(n_950)
);

INVx2_ASAP7_75t_L g951 ( 
.A(n_647),
.Y(n_951)
);

INVx2_ASAP7_75t_L g952 ( 
.A(n_675),
.Y(n_952)
);

NAND2xp5_ASAP7_75t_L g953 ( 
.A(n_694),
.B(n_552),
.Y(n_953)
);

NOR2xp33_ASAP7_75t_L g954 ( 
.A(n_699),
.B(n_584),
.Y(n_954)
);

BUFx2_ASAP7_75t_L g955 ( 
.A(n_766),
.Y(n_955)
);

INVx1_ASAP7_75t_L g956 ( 
.A(n_675),
.Y(n_956)
);

AOI22xp33_ASAP7_75t_L g957 ( 
.A1(n_802),
.A2(n_571),
.B1(n_572),
.B2(n_639),
.Y(n_957)
);

INVx2_ASAP7_75t_L g958 ( 
.A(n_693),
.Y(n_958)
);

AOI22xp33_ASAP7_75t_L g959 ( 
.A1(n_724),
.A2(n_572),
.B1(n_642),
.B2(n_639),
.Y(n_959)
);

NAND2xp5_ASAP7_75t_SL g960 ( 
.A(n_794),
.B(n_552),
.Y(n_960)
);

NAND2xp5_ASAP7_75t_SL g961 ( 
.A(n_743),
.B(n_552),
.Y(n_961)
);

NOR2xp33_ASAP7_75t_L g962 ( 
.A(n_710),
.B(n_578),
.Y(n_962)
);

NAND2xp5_ASAP7_75t_L g963 ( 
.A(n_724),
.B(n_725),
.Y(n_963)
);

AND2x6_ASAP7_75t_SL g964 ( 
.A(n_676),
.B(n_19),
.Y(n_964)
);

NAND2xp5_ASAP7_75t_SL g965 ( 
.A(n_661),
.B(n_552),
.Y(n_965)
);

NAND2xp5_ASAP7_75t_L g966 ( 
.A(n_740),
.B(n_572),
.Y(n_966)
);

INVx1_ASAP7_75t_L g967 ( 
.A(n_693),
.Y(n_967)
);

INVx3_ASAP7_75t_L g968 ( 
.A(n_700),
.Y(n_968)
);

INVx1_ASAP7_75t_L g969 ( 
.A(n_700),
.Y(n_969)
);

BUFx2_ASAP7_75t_L g970 ( 
.A(n_766),
.Y(n_970)
);

INVxp67_ASAP7_75t_L g971 ( 
.A(n_740),
.Y(n_971)
);

NOR2xp33_ASAP7_75t_L g972 ( 
.A(n_719),
.B(n_595),
.Y(n_972)
);

NAND2xp5_ASAP7_75t_SL g973 ( 
.A(n_797),
.B(n_572),
.Y(n_973)
);

NAND2xp5_ASAP7_75t_L g974 ( 
.A(n_706),
.B(n_595),
.Y(n_974)
);

INVx2_ASAP7_75t_SL g975 ( 
.A(n_726),
.Y(n_975)
);

AND2x2_ASAP7_75t_L g976 ( 
.A(n_668),
.B(n_610),
.Y(n_976)
);

NOR2xp33_ASAP7_75t_L g977 ( 
.A(n_707),
.B(n_595),
.Y(n_977)
);

INVx2_ASAP7_75t_L g978 ( 
.A(n_701),
.Y(n_978)
);

INVxp67_ASAP7_75t_L g979 ( 
.A(n_745),
.Y(n_979)
);

NAND2xp5_ASAP7_75t_SL g980 ( 
.A(n_652),
.B(n_643),
.Y(n_980)
);

NAND2xp5_ASAP7_75t_L g981 ( 
.A(n_652),
.B(n_568),
.Y(n_981)
);

INVx1_ASAP7_75t_L g982 ( 
.A(n_701),
.Y(n_982)
);

INVx2_ASAP7_75t_SL g983 ( 
.A(n_778),
.Y(n_983)
);

AND2x4_ASAP7_75t_L g984 ( 
.A(n_648),
.B(n_538),
.Y(n_984)
);

INVx1_ASAP7_75t_SL g985 ( 
.A(n_732),
.Y(n_985)
);

INVx1_ASAP7_75t_SL g986 ( 
.A(n_727),
.Y(n_986)
);

INVx1_ASAP7_75t_SL g987 ( 
.A(n_730),
.Y(n_987)
);

NAND2xp5_ASAP7_75t_L g988 ( 
.A(n_738),
.B(n_568),
.Y(n_988)
);

NAND2xp5_ASAP7_75t_L g989 ( 
.A(n_733),
.B(n_568),
.Y(n_989)
);

INVx2_ASAP7_75t_L g990 ( 
.A(n_702),
.Y(n_990)
);

NAND2xp5_ASAP7_75t_L g991 ( 
.A(n_736),
.B(n_748),
.Y(n_991)
);

NAND2xp5_ASAP7_75t_L g992 ( 
.A(n_749),
.B(n_578),
.Y(n_992)
);

NOR2xp33_ASAP7_75t_L g993 ( 
.A(n_720),
.B(n_578),
.Y(n_993)
);

NAND2xp5_ASAP7_75t_L g994 ( 
.A(n_758),
.B(n_584),
.Y(n_994)
);

INVx2_ASAP7_75t_SL g995 ( 
.A(n_784),
.Y(n_995)
);

NOR2xp33_ASAP7_75t_L g996 ( 
.A(n_745),
.B(n_765),
.Y(n_996)
);

NAND2xp5_ASAP7_75t_SL g997 ( 
.A(n_717),
.B(n_584),
.Y(n_997)
);

INVx1_ASAP7_75t_L g998 ( 
.A(n_702),
.Y(n_998)
);

NAND3xp33_ASAP7_75t_SL g999 ( 
.A(n_689),
.B(n_22),
.C(n_25),
.Y(n_999)
);

INVx1_ASAP7_75t_L g1000 ( 
.A(n_723),
.Y(n_1000)
);

AOI21xp5_ASAP7_75t_L g1001 ( 
.A1(n_813),
.A2(n_189),
.B(n_180),
.Y(n_1001)
);

AND2x2_ASAP7_75t_L g1002 ( 
.A(n_770),
.B(n_787),
.Y(n_1002)
);

NAND2xp5_ASAP7_75t_SL g1003 ( 
.A(n_803),
.B(n_616),
.Y(n_1003)
);

INVx1_ASAP7_75t_L g1004 ( 
.A(n_723),
.Y(n_1004)
);

INVx2_ASAP7_75t_L g1005 ( 
.A(n_728),
.Y(n_1005)
);

BUFx2_ASAP7_75t_L g1006 ( 
.A(n_780),
.Y(n_1006)
);

INVxp67_ASAP7_75t_L g1007 ( 
.A(n_852),
.Y(n_1007)
);

AOI21xp5_ASAP7_75t_L g1008 ( 
.A1(n_826),
.A2(n_809),
.B(n_687),
.Y(n_1008)
);

INVx2_ASAP7_75t_L g1009 ( 
.A(n_817),
.Y(n_1009)
);

AOI22xp33_ASAP7_75t_L g1010 ( 
.A1(n_910),
.A2(n_790),
.B1(n_796),
.B2(n_728),
.Y(n_1010)
);

NAND2xp5_ASAP7_75t_SL g1011 ( 
.A(n_971),
.B(n_764),
.Y(n_1011)
);

O2A1O1Ixp33_ASAP7_75t_SL g1012 ( 
.A1(n_971),
.A2(n_687),
.B(n_786),
.C(n_753),
.Y(n_1012)
);

AOI22xp33_ASAP7_75t_L g1013 ( 
.A1(n_839),
.A2(n_729),
.B1(n_747),
.B2(n_777),
.Y(n_1013)
);

INVx4_ASAP7_75t_L g1014 ( 
.A(n_872),
.Y(n_1014)
);

OAI22xp5_ASAP7_75t_L g1015 ( 
.A1(n_926),
.A2(n_698),
.B1(n_782),
.B2(n_729),
.Y(n_1015)
);

INVx1_ASAP7_75t_L g1016 ( 
.A(n_816),
.Y(n_1016)
);

AOI21xp5_ASAP7_75t_L g1017 ( 
.A1(n_819),
.A2(n_698),
.B(n_645),
.Y(n_1017)
);

AND2x2_ASAP7_75t_L g1018 ( 
.A(n_922),
.B(n_747),
.Y(n_1018)
);

A2O1A1Ixp33_ASAP7_75t_L g1019 ( 
.A1(n_996),
.A2(n_671),
.B(n_806),
.C(n_721),
.Y(n_1019)
);

OAI22xp5_ASAP7_75t_L g1020 ( 
.A1(n_926),
.A2(n_754),
.B1(n_801),
.B2(n_805),
.Y(n_1020)
);

INVxp67_ASAP7_75t_L g1021 ( 
.A(n_831),
.Y(n_1021)
);

INVx3_ASAP7_75t_L g1022 ( 
.A(n_872),
.Y(n_1022)
);

NOR2xp33_ASAP7_75t_R g1023 ( 
.A(n_846),
.B(n_800),
.Y(n_1023)
);

O2A1O1Ixp33_ASAP7_75t_L g1024 ( 
.A1(n_908),
.A2(n_798),
.B(n_769),
.C(n_807),
.Y(n_1024)
);

AND2x2_ASAP7_75t_L g1025 ( 
.A(n_821),
.B(n_27),
.Y(n_1025)
);

BUFx6f_ASAP7_75t_L g1026 ( 
.A(n_872),
.Y(n_1026)
);

INVx4_ASAP7_75t_L g1027 ( 
.A(n_872),
.Y(n_1027)
);

AOI22xp5_ASAP7_75t_L g1028 ( 
.A1(n_823),
.A2(n_616),
.B1(n_510),
.B2(n_189),
.Y(n_1028)
);

AOI21xp5_ASAP7_75t_L g1029 ( 
.A1(n_966),
.A2(n_189),
.B(n_180),
.Y(n_1029)
);

O2A1O1Ixp5_ASAP7_75t_L g1030 ( 
.A1(n_902),
.A2(n_27),
.B(n_31),
.C(n_35),
.Y(n_1030)
);

INVx1_ASAP7_75t_L g1031 ( 
.A(n_827),
.Y(n_1031)
);

INVxp67_ASAP7_75t_SL g1032 ( 
.A(n_957),
.Y(n_1032)
);

A2O1A1Ixp33_ASAP7_75t_L g1033 ( 
.A1(n_996),
.A2(n_189),
.B(n_180),
.C(n_171),
.Y(n_1033)
);

A2O1A1Ixp33_ASAP7_75t_SL g1034 ( 
.A1(n_954),
.A2(n_31),
.B(n_35),
.C(n_40),
.Y(n_1034)
);

AOI21xp5_ASAP7_75t_L g1035 ( 
.A1(n_842),
.A2(n_180),
.B(n_171),
.Y(n_1035)
);

AOI21xp5_ASAP7_75t_L g1036 ( 
.A1(n_851),
.A2(n_171),
.B(n_169),
.Y(n_1036)
);

INVx1_ASAP7_75t_L g1037 ( 
.A(n_847),
.Y(n_1037)
);

NOR2xp33_ASAP7_75t_L g1038 ( 
.A(n_986),
.B(n_40),
.Y(n_1038)
);

NAND3xp33_ASAP7_75t_L g1039 ( 
.A(n_944),
.B(n_171),
.C(n_616),
.Y(n_1039)
);

NAND2xp5_ASAP7_75t_L g1040 ( 
.A(n_955),
.B(n_42),
.Y(n_1040)
);

OR2x6_ASAP7_75t_L g1041 ( 
.A(n_825),
.B(n_616),
.Y(n_1041)
);

AOI21xp5_ASAP7_75t_L g1042 ( 
.A1(n_829),
.A2(n_616),
.B(n_510),
.Y(n_1042)
);

AND2x6_ASAP7_75t_L g1043 ( 
.A(n_836),
.B(n_616),
.Y(n_1043)
);

A2O1A1Ixp33_ASAP7_75t_L g1044 ( 
.A1(n_963),
.A2(n_510),
.B(n_43),
.C(n_54),
.Y(n_1044)
);

BUFx6f_ASAP7_75t_L g1045 ( 
.A(n_820),
.Y(n_1045)
);

OAI21x1_ASAP7_75t_L g1046 ( 
.A1(n_849),
.A2(n_510),
.B(n_53),
.Y(n_1046)
);

AOI21xp5_ASAP7_75t_L g1047 ( 
.A1(n_833),
.A2(n_510),
.B(n_57),
.Y(n_1047)
);

AOI21xp5_ASAP7_75t_L g1048 ( 
.A1(n_837),
.A2(n_98),
.B(n_64),
.Y(n_1048)
);

HB1xp67_ASAP7_75t_L g1049 ( 
.A(n_824),
.Y(n_1049)
);

NAND3xp33_ASAP7_75t_SL g1050 ( 
.A(n_970),
.B(n_987),
.C(n_944),
.Y(n_1050)
);

AOI21xp5_ASAP7_75t_L g1051 ( 
.A1(n_981),
.A2(n_105),
.B(n_67),
.Y(n_1051)
);

NAND2xp5_ASAP7_75t_L g1052 ( 
.A(n_941),
.B(n_43),
.Y(n_1052)
);

AOI21xp5_ASAP7_75t_L g1053 ( 
.A1(n_991),
.A2(n_72),
.B(n_74),
.Y(n_1053)
);

OAI22xp5_ASAP7_75t_L g1054 ( 
.A1(n_867),
.A2(n_78),
.B1(n_93),
.B2(n_94),
.Y(n_1054)
);

AOI21x1_ASAP7_75t_L g1055 ( 
.A1(n_965),
.A2(n_95),
.B(n_97),
.Y(n_1055)
);

BUFx6f_ASAP7_75t_L g1056 ( 
.A(n_820),
.Y(n_1056)
);

OAI22xp5_ASAP7_75t_SL g1057 ( 
.A1(n_929),
.A2(n_114),
.B1(n_121),
.B2(n_123),
.Y(n_1057)
);

BUFx8_ASAP7_75t_L g1058 ( 
.A(n_864),
.Y(n_1058)
);

NOR3xp33_ASAP7_75t_SL g1059 ( 
.A(n_999),
.B(n_893),
.C(n_869),
.Y(n_1059)
);

INVx2_ASAP7_75t_L g1060 ( 
.A(n_835),
.Y(n_1060)
);

INVx1_ASAP7_75t_L g1061 ( 
.A(n_848),
.Y(n_1061)
);

AOI21xp5_ASAP7_75t_L g1062 ( 
.A1(n_854),
.A2(n_125),
.B(n_133),
.Y(n_1062)
);

NAND2x1p5_ASAP7_75t_L g1063 ( 
.A(n_846),
.B(n_151),
.Y(n_1063)
);

NOR2x1p5_ASAP7_75t_L g1064 ( 
.A(n_917),
.B(n_162),
.Y(n_1064)
);

AND2x4_ASAP7_75t_L g1065 ( 
.A(n_830),
.B(n_164),
.Y(n_1065)
);

NAND2xp5_ASAP7_75t_L g1066 ( 
.A(n_887),
.B(n_1002),
.Y(n_1066)
);

OAI22xp5_ASAP7_75t_L g1067 ( 
.A1(n_855),
.A2(n_882),
.B1(n_915),
.B2(n_890),
.Y(n_1067)
);

O2A1O1Ixp5_ASAP7_75t_L g1068 ( 
.A1(n_960),
.A2(n_997),
.B(n_977),
.C(n_866),
.Y(n_1068)
);

OR2x6_ASAP7_75t_L g1069 ( 
.A(n_824),
.B(n_865),
.Y(n_1069)
);

INVx1_ASAP7_75t_L g1070 ( 
.A(n_859),
.Y(n_1070)
);

A2O1A1Ixp33_ASAP7_75t_L g1071 ( 
.A1(n_850),
.A2(n_993),
.B(n_855),
.C(n_977),
.Y(n_1071)
);

AOI21xp5_ASAP7_75t_L g1072 ( 
.A1(n_965),
.A2(n_992),
.B(n_989),
.Y(n_1072)
);

NAND2xp5_ASAP7_75t_L g1073 ( 
.A(n_1006),
.B(n_905),
.Y(n_1073)
);

INVx2_ASAP7_75t_L g1074 ( 
.A(n_840),
.Y(n_1074)
);

O2A1O1Ixp33_ASAP7_75t_L g1075 ( 
.A1(n_999),
.A2(n_907),
.B(n_884),
.C(n_923),
.Y(n_1075)
);

NOR2xp33_ASAP7_75t_R g1076 ( 
.A(n_853),
.B(n_858),
.Y(n_1076)
);

NOR2xp33_ASAP7_75t_L g1077 ( 
.A(n_985),
.B(n_979),
.Y(n_1077)
);

AOI21xp5_ASAP7_75t_L g1078 ( 
.A1(n_994),
.A2(n_948),
.B(n_953),
.Y(n_1078)
);

NOR2xp33_ASAP7_75t_L g1079 ( 
.A(n_979),
.B(n_884),
.Y(n_1079)
);

INVx3_ASAP7_75t_L g1080 ( 
.A(n_860),
.Y(n_1080)
);

INVx1_ASAP7_75t_L g1081 ( 
.A(n_873),
.Y(n_1081)
);

NAND2xp5_ASAP7_75t_L g1082 ( 
.A(n_877),
.B(n_891),
.Y(n_1082)
);

AND2x2_ASAP7_75t_L g1083 ( 
.A(n_884),
.B(n_832),
.Y(n_1083)
);

INVx4_ASAP7_75t_L g1084 ( 
.A(n_928),
.Y(n_1084)
);

AOI21xp5_ASAP7_75t_L g1085 ( 
.A1(n_849),
.A2(n_980),
.B(n_933),
.Y(n_1085)
);

NAND2xp5_ASAP7_75t_L g1086 ( 
.A(n_906),
.B(n_909),
.Y(n_1086)
);

NOR2xp33_ASAP7_75t_L g1087 ( 
.A(n_983),
.B(n_995),
.Y(n_1087)
);

INVx1_ASAP7_75t_L g1088 ( 
.A(n_914),
.Y(n_1088)
);

NAND2xp5_ASAP7_75t_L g1089 ( 
.A(n_930),
.B(n_832),
.Y(n_1089)
);

OAI22xp5_ASAP7_75t_L g1090 ( 
.A1(n_936),
.A2(n_993),
.B1(n_988),
.B2(n_850),
.Y(n_1090)
);

NAND2xp5_ASAP7_75t_SL g1091 ( 
.A(n_928),
.B(n_818),
.Y(n_1091)
);

NOR2xp33_ASAP7_75t_L g1092 ( 
.A(n_975),
.B(n_929),
.Y(n_1092)
);

NOR2xp33_ASAP7_75t_L g1093 ( 
.A(n_947),
.B(n_889),
.Y(n_1093)
);

AOI21xp5_ASAP7_75t_L g1094 ( 
.A1(n_980),
.A2(n_933),
.B(n_921),
.Y(n_1094)
);

INVxp67_ASAP7_75t_L g1095 ( 
.A(n_869),
.Y(n_1095)
);

O2A1O1Ixp33_ASAP7_75t_SL g1096 ( 
.A1(n_868),
.A2(n_921),
.B(n_862),
.C(n_997),
.Y(n_1096)
);

NAND2xp5_ASAP7_75t_L g1097 ( 
.A(n_894),
.B(n_913),
.Y(n_1097)
);

BUFx6f_ASAP7_75t_L g1098 ( 
.A(n_820),
.Y(n_1098)
);

NAND2xp5_ASAP7_75t_L g1099 ( 
.A(n_894),
.B(n_913),
.Y(n_1099)
);

NAND2xp5_ASAP7_75t_L g1100 ( 
.A(n_927),
.B(n_925),
.Y(n_1100)
);

A2O1A1Ixp33_ASAP7_75t_L g1101 ( 
.A1(n_954),
.A2(n_962),
.B(n_893),
.C(n_972),
.Y(n_1101)
);

NAND2xp5_ASAP7_75t_L g1102 ( 
.A(n_858),
.B(n_885),
.Y(n_1102)
);

NOR2xp33_ASAP7_75t_L g1103 ( 
.A(n_889),
.B(n_885),
.Y(n_1103)
);

INVx8_ASAP7_75t_L g1104 ( 
.A(n_860),
.Y(n_1104)
);

AOI21xp5_ASAP7_75t_L g1105 ( 
.A1(n_868),
.A2(n_962),
.B(n_883),
.Y(n_1105)
);

HB1xp67_ASAP7_75t_L g1106 ( 
.A(n_860),
.Y(n_1106)
);

AND2x4_ASAP7_75t_L g1107 ( 
.A(n_830),
.B(n_836),
.Y(n_1107)
);

INVx2_ASAP7_75t_L g1108 ( 
.A(n_844),
.Y(n_1108)
);

INVx1_ASAP7_75t_L g1109 ( 
.A(n_938),
.Y(n_1109)
);

NAND2xp5_ASAP7_75t_L g1110 ( 
.A(n_899),
.B(n_950),
.Y(n_1110)
);

AO22x1_ASAP7_75t_L g1111 ( 
.A1(n_880),
.A2(n_950),
.B1(n_904),
.B2(n_899),
.Y(n_1111)
);

NAND2xp5_ASAP7_75t_L g1112 ( 
.A(n_950),
.B(n_878),
.Y(n_1112)
);

CKINVDCx5p33_ASAP7_75t_R g1113 ( 
.A(n_964),
.Y(n_1113)
);

INVx1_ASAP7_75t_L g1114 ( 
.A(n_942),
.Y(n_1114)
);

INVx1_ASAP7_75t_L g1115 ( 
.A(n_956),
.Y(n_1115)
);

INVx1_ASAP7_75t_L g1116 ( 
.A(n_967),
.Y(n_1116)
);

OAI21xp5_ASAP7_75t_L g1117 ( 
.A1(n_896),
.A2(n_863),
.B(n_924),
.Y(n_1117)
);

INVx2_ASAP7_75t_L g1118 ( 
.A(n_861),
.Y(n_1118)
);

AOI33xp33_ASAP7_75t_L g1119 ( 
.A1(n_976),
.A2(n_881),
.A3(n_841),
.B1(n_834),
.B2(n_931),
.B3(n_959),
.Y(n_1119)
);

NAND2xp5_ASAP7_75t_L g1120 ( 
.A(n_950),
.B(n_892),
.Y(n_1120)
);

AOI21xp5_ASAP7_75t_L g1121 ( 
.A1(n_883),
.A2(n_901),
.B(n_897),
.Y(n_1121)
);

BUFx2_ASAP7_75t_L g1122 ( 
.A(n_822),
.Y(n_1122)
);

INVx2_ASAP7_75t_L g1123 ( 
.A(n_870),
.Y(n_1123)
);

NOR2xp33_ASAP7_75t_L g1124 ( 
.A(n_880),
.B(n_939),
.Y(n_1124)
);

CKINVDCx20_ASAP7_75t_R g1125 ( 
.A(n_838),
.Y(n_1125)
);

NOR2xp33_ASAP7_75t_L g1126 ( 
.A(n_946),
.B(n_972),
.Y(n_1126)
);

AO21x1_ASAP7_75t_L g1127 ( 
.A1(n_973),
.A2(n_943),
.B(n_935),
.Y(n_1127)
);

NAND2xp5_ASAP7_75t_L g1128 ( 
.A(n_950),
.B(n_920),
.Y(n_1128)
);

NOR3xp33_ASAP7_75t_L g1129 ( 
.A(n_961),
.B(n_916),
.C(n_856),
.Y(n_1129)
);

INVx1_ASAP7_75t_L g1130 ( 
.A(n_969),
.Y(n_1130)
);

INVx1_ASAP7_75t_SL g1131 ( 
.A(n_937),
.Y(n_1131)
);

HAxp5_ASAP7_75t_L g1132 ( 
.A(n_898),
.B(n_881),
.CON(n_1132),
.SN(n_1132)
);

OAI22xp5_ASAP7_75t_L g1133 ( 
.A1(n_957),
.A2(n_959),
.B1(n_828),
.B2(n_818),
.Y(n_1133)
);

OAI22xp5_ASAP7_75t_L g1134 ( 
.A1(n_871),
.A2(n_928),
.B1(n_937),
.B2(n_974),
.Y(n_1134)
);

INVx3_ASAP7_75t_L g1135 ( 
.A(n_928),
.Y(n_1135)
);

AOI22xp5_ASAP7_75t_L g1136 ( 
.A1(n_937),
.A2(n_918),
.B1(n_934),
.B2(n_968),
.Y(n_1136)
);

NAND2xp5_ASAP7_75t_L g1137 ( 
.A(n_934),
.B(n_968),
.Y(n_1137)
);

INVx1_ASAP7_75t_L g1138 ( 
.A(n_982),
.Y(n_1138)
);

AOI21xp5_ASAP7_75t_L g1139 ( 
.A1(n_935),
.A2(n_943),
.B(n_1003),
.Y(n_1139)
);

AOI21xp5_ASAP7_75t_L g1140 ( 
.A1(n_1003),
.A2(n_820),
.B(n_843),
.Y(n_1140)
);

OR2x6_ASAP7_75t_L g1141 ( 
.A(n_984),
.B(n_916),
.Y(n_1141)
);

BUFx2_ASAP7_75t_L g1142 ( 
.A(n_843),
.Y(n_1142)
);

INVx2_ASAP7_75t_L g1143 ( 
.A(n_874),
.Y(n_1143)
);

NOR2xp33_ASAP7_75t_L g1144 ( 
.A(n_949),
.B(n_1000),
.Y(n_1144)
);

NAND2xp5_ASAP7_75t_L g1145 ( 
.A(n_998),
.B(n_1004),
.Y(n_1145)
);

AOI21xp5_ASAP7_75t_L g1146 ( 
.A1(n_843),
.A2(n_879),
.B(n_857),
.Y(n_1146)
);

O2A1O1Ixp33_ASAP7_75t_L g1147 ( 
.A1(n_1001),
.A2(n_1005),
.B(n_990),
.C(n_978),
.Y(n_1147)
);

OAI22xp5_ASAP7_75t_L g1148 ( 
.A1(n_843),
.A2(n_911),
.B1(n_857),
.B2(n_875),
.Y(n_1148)
);

NAND2xp33_ASAP7_75t_L g1149 ( 
.A(n_857),
.B(n_875),
.Y(n_1149)
);

INVx2_ASAP7_75t_L g1150 ( 
.A(n_876),
.Y(n_1150)
);

BUFx6f_ASAP7_75t_L g1151 ( 
.A(n_857),
.Y(n_1151)
);

NOR2xp33_ASAP7_75t_L g1152 ( 
.A(n_949),
.B(n_911),
.Y(n_1152)
);

CKINVDCx5p33_ASAP7_75t_R g1153 ( 
.A(n_875),
.Y(n_1153)
);

INVx4_ASAP7_75t_L g1154 ( 
.A(n_875),
.Y(n_1154)
);

NAND2xp5_ASAP7_75t_SL g1155 ( 
.A(n_879),
.B(n_911),
.Y(n_1155)
);

INVx1_ASAP7_75t_L g1156 ( 
.A(n_886),
.Y(n_1156)
);

NAND2xp5_ASAP7_75t_L g1157 ( 
.A(n_888),
.B(n_958),
.Y(n_1157)
);

AOI21xp5_ASAP7_75t_L g1158 ( 
.A1(n_879),
.A2(n_911),
.B(n_919),
.Y(n_1158)
);

INVx1_ASAP7_75t_SL g1159 ( 
.A(n_845),
.Y(n_1159)
);

NOR2xp33_ASAP7_75t_L g1160 ( 
.A(n_949),
.B(n_879),
.Y(n_1160)
);

NAND2xp5_ASAP7_75t_SL g1161 ( 
.A(n_949),
.B(n_984),
.Y(n_1161)
);

AOI21xp5_ASAP7_75t_L g1162 ( 
.A1(n_932),
.A2(n_1001),
.B(n_900),
.Y(n_1162)
);

AOI21xp5_ASAP7_75t_L g1163 ( 
.A1(n_932),
.A2(n_895),
.B(n_903),
.Y(n_1163)
);

BUFx6f_ASAP7_75t_L g1164 ( 
.A(n_1107),
.Y(n_1164)
);

AOI21xp5_ASAP7_75t_L g1165 ( 
.A1(n_1071),
.A2(n_1101),
.B(n_1105),
.Y(n_1165)
);

INVx1_ASAP7_75t_L g1166 ( 
.A(n_1016),
.Y(n_1166)
);

OAI21x1_ASAP7_75t_SL g1167 ( 
.A1(n_1075),
.A2(n_931),
.B(n_912),
.Y(n_1167)
);

O2A1O1Ixp5_ASAP7_75t_L g1168 ( 
.A1(n_1011),
.A2(n_952),
.B(n_940),
.C(n_945),
.Y(n_1168)
);

NAND2xp5_ASAP7_75t_L g1169 ( 
.A(n_1066),
.B(n_951),
.Y(n_1169)
);

OAI21x1_ASAP7_75t_L g1170 ( 
.A1(n_1085),
.A2(n_932),
.B(n_1046),
.Y(n_1170)
);

OAI21x1_ASAP7_75t_L g1171 ( 
.A1(n_1162),
.A2(n_932),
.B(n_1072),
.Y(n_1171)
);

OAI21x1_ASAP7_75t_L g1172 ( 
.A1(n_1139),
.A2(n_1094),
.B(n_1078),
.Y(n_1172)
);

INVx1_ASAP7_75t_L g1173 ( 
.A(n_1031),
.Y(n_1173)
);

AND2x2_ASAP7_75t_L g1174 ( 
.A(n_1018),
.B(n_1025),
.Y(n_1174)
);

A2O1A1Ixp33_ASAP7_75t_L g1175 ( 
.A1(n_1119),
.A2(n_1059),
.B(n_1090),
.C(n_1028),
.Y(n_1175)
);

OAI21x1_ASAP7_75t_SL g1176 ( 
.A1(n_1067),
.A2(n_1110),
.B(n_1146),
.Y(n_1176)
);

OA21x2_ASAP7_75t_L g1177 ( 
.A1(n_1068),
.A2(n_1117),
.B(n_1121),
.Y(n_1177)
);

OAI21x1_ASAP7_75t_L g1178 ( 
.A1(n_1158),
.A2(n_1029),
.B(n_1140),
.Y(n_1178)
);

OAI21x1_ASAP7_75t_L g1179 ( 
.A1(n_1055),
.A2(n_1036),
.B(n_1035),
.Y(n_1179)
);

INVx3_ASAP7_75t_L g1180 ( 
.A(n_1014),
.Y(n_1180)
);

OAI21x1_ASAP7_75t_L g1181 ( 
.A1(n_1147),
.A2(n_1127),
.B(n_1017),
.Y(n_1181)
);

OAI21x1_ASAP7_75t_L g1182 ( 
.A1(n_1163),
.A2(n_1134),
.B(n_1047),
.Y(n_1182)
);

NAND3xp33_ASAP7_75t_L g1183 ( 
.A(n_1010),
.B(n_1039),
.C(n_1038),
.Y(n_1183)
);

INVx1_ASAP7_75t_L g1184 ( 
.A(n_1037),
.Y(n_1184)
);

AO21x2_ASAP7_75t_L g1185 ( 
.A1(n_1112),
.A2(n_1120),
.B(n_1033),
.Y(n_1185)
);

OAI21xp5_ASAP7_75t_L g1186 ( 
.A1(n_1008),
.A2(n_1095),
.B(n_1019),
.Y(n_1186)
);

OAI21x1_ASAP7_75t_L g1187 ( 
.A1(n_1148),
.A2(n_1051),
.B(n_1133),
.Y(n_1187)
);

INVx1_ASAP7_75t_L g1188 ( 
.A(n_1061),
.Y(n_1188)
);

AO31x2_ASAP7_75t_L g1189 ( 
.A1(n_1097),
.A2(n_1099),
.A3(n_1144),
.B(n_1089),
.Y(n_1189)
);

OAI21xp5_ASAP7_75t_L g1190 ( 
.A1(n_1126),
.A2(n_1015),
.B(n_1096),
.Y(n_1190)
);

BUFx3_ASAP7_75t_L g1191 ( 
.A(n_1058),
.Y(n_1191)
);

BUFx6f_ASAP7_75t_L g1192 ( 
.A(n_1107),
.Y(n_1192)
);

INVx1_ASAP7_75t_L g1193 ( 
.A(n_1070),
.Y(n_1193)
);

AOI21xp5_ASAP7_75t_L g1194 ( 
.A1(n_1149),
.A2(n_1012),
.B(n_1048),
.Y(n_1194)
);

O2A1O1Ixp5_ASAP7_75t_L g1195 ( 
.A1(n_1091),
.A2(n_1155),
.B(n_1054),
.C(n_1044),
.Y(n_1195)
);

XNOR2xp5_ASAP7_75t_L g1196 ( 
.A(n_1113),
.B(n_1122),
.Y(n_1196)
);

AND2x4_ASAP7_75t_L g1197 ( 
.A(n_1065),
.B(n_1141),
.Y(n_1197)
);

BUFx10_ASAP7_75t_L g1198 ( 
.A(n_1092),
.Y(n_1198)
);

NAND2xp5_ASAP7_75t_L g1199 ( 
.A(n_1077),
.B(n_1100),
.Y(n_1199)
);

OAI21x1_ASAP7_75t_L g1200 ( 
.A1(n_1128),
.A2(n_1136),
.B(n_1062),
.Y(n_1200)
);

INVx1_ASAP7_75t_L g1201 ( 
.A(n_1081),
.Y(n_1201)
);

OAI21x1_ASAP7_75t_L g1202 ( 
.A1(n_1136),
.A2(n_1053),
.B(n_1145),
.Y(n_1202)
);

AO21x1_ASAP7_75t_L g1203 ( 
.A1(n_1129),
.A2(n_1020),
.B(n_1079),
.Y(n_1203)
);

INVx3_ASAP7_75t_L g1204 ( 
.A(n_1014),
.Y(n_1204)
);

INVx1_ASAP7_75t_SL g1205 ( 
.A(n_1073),
.Y(n_1205)
);

AOI21xp5_ASAP7_75t_L g1206 ( 
.A1(n_1082),
.A2(n_1086),
.B(n_1102),
.Y(n_1206)
);

AO32x2_ASAP7_75t_L g1207 ( 
.A1(n_1057),
.A2(n_1154),
.A3(n_1034),
.B1(n_1084),
.B2(n_1132),
.Y(n_1207)
);

AOI21x1_ASAP7_75t_L g1208 ( 
.A1(n_1137),
.A2(n_1111),
.B(n_1161),
.Y(n_1208)
);

OAI22x1_ASAP7_75t_L g1209 ( 
.A1(n_1064),
.A2(n_1159),
.B1(n_1083),
.B2(n_1093),
.Y(n_1209)
);

HB1xp67_ASAP7_75t_L g1210 ( 
.A(n_1007),
.Y(n_1210)
);

AO21x1_ASAP7_75t_L g1211 ( 
.A1(n_1152),
.A2(n_1160),
.B(n_1052),
.Y(n_1211)
);

INVx1_ASAP7_75t_L g1212 ( 
.A(n_1088),
.Y(n_1212)
);

INVx1_ASAP7_75t_L g1213 ( 
.A(n_1109),
.Y(n_1213)
);

NAND3xp33_ASAP7_75t_L g1214 ( 
.A(n_1040),
.B(n_1030),
.C(n_1013),
.Y(n_1214)
);

AO31x2_ASAP7_75t_L g1215 ( 
.A1(n_1114),
.A2(n_1130),
.A3(n_1115),
.B(n_1116),
.Y(n_1215)
);

OAI21xp33_ASAP7_75t_L g1216 ( 
.A1(n_1050),
.A2(n_1087),
.B(n_1021),
.Y(n_1216)
);

AO32x2_ASAP7_75t_L g1217 ( 
.A1(n_1154),
.A2(n_1084),
.A3(n_1027),
.B1(n_1125),
.B2(n_1032),
.Y(n_1217)
);

OAI21x1_ASAP7_75t_L g1218 ( 
.A1(n_1135),
.A2(n_1080),
.B(n_1042),
.Y(n_1218)
);

OAI22xp5_ASAP7_75t_L g1219 ( 
.A1(n_1153),
.A2(n_1141),
.B1(n_1065),
.B2(n_1131),
.Y(n_1219)
);

INVx1_ASAP7_75t_L g1220 ( 
.A(n_1138),
.Y(n_1220)
);

BUFx2_ASAP7_75t_L g1221 ( 
.A(n_1058),
.Y(n_1221)
);

HB1xp67_ASAP7_75t_L g1222 ( 
.A(n_1049),
.Y(n_1222)
);

A2O1A1Ixp33_ASAP7_75t_L g1223 ( 
.A1(n_1124),
.A2(n_1024),
.B(n_1103),
.C(n_1135),
.Y(n_1223)
);

INVx1_ASAP7_75t_L g1224 ( 
.A(n_1156),
.Y(n_1224)
);

NAND2xp33_ASAP7_75t_L g1225 ( 
.A(n_1026),
.B(n_1076),
.Y(n_1225)
);

INVx2_ASAP7_75t_L g1226 ( 
.A(n_1060),
.Y(n_1226)
);

NAND2xp5_ASAP7_75t_SL g1227 ( 
.A(n_1026),
.B(n_1098),
.Y(n_1227)
);

CKINVDCx20_ASAP7_75t_R g1228 ( 
.A(n_1104),
.Y(n_1228)
);

A2O1A1Ixp33_ASAP7_75t_L g1229 ( 
.A1(n_1080),
.A2(n_1022),
.B(n_1106),
.C(n_1142),
.Y(n_1229)
);

AO31x2_ASAP7_75t_L g1230 ( 
.A1(n_1074),
.A2(n_1108),
.A3(n_1150),
.B(n_1143),
.Y(n_1230)
);

AOI21xp5_ASAP7_75t_SL g1231 ( 
.A1(n_1041),
.A2(n_1141),
.B(n_1063),
.Y(n_1231)
);

INVx1_ASAP7_75t_L g1232 ( 
.A(n_1118),
.Y(n_1232)
);

OA21x2_ASAP7_75t_L g1233 ( 
.A1(n_1157),
.A2(n_1123),
.B(n_1151),
.Y(n_1233)
);

NAND2xp5_ASAP7_75t_L g1234 ( 
.A(n_1069),
.B(n_1104),
.Y(n_1234)
);

OAI21x1_ASAP7_75t_L g1235 ( 
.A1(n_1022),
.A2(n_1045),
.B(n_1098),
.Y(n_1235)
);

AOI21xp5_ASAP7_75t_L g1236 ( 
.A1(n_1045),
.A2(n_1151),
.B(n_1098),
.Y(n_1236)
);

NAND2xp5_ASAP7_75t_L g1237 ( 
.A(n_1151),
.B(n_1056),
.Y(n_1237)
);

NAND2xp5_ASAP7_75t_SL g1238 ( 
.A(n_1026),
.B(n_1045),
.Y(n_1238)
);

AOI21x1_ASAP7_75t_L g1239 ( 
.A1(n_1041),
.A2(n_1069),
.B(n_1056),
.Y(n_1239)
);

NAND2xp5_ASAP7_75t_L g1240 ( 
.A(n_1056),
.B(n_1027),
.Y(n_1240)
);

NAND2xp5_ASAP7_75t_L g1241 ( 
.A(n_1041),
.B(n_1043),
.Y(n_1241)
);

AO31x2_ASAP7_75t_L g1242 ( 
.A1(n_1043),
.A2(n_1127),
.A3(n_1071),
.B(n_1078),
.Y(n_1242)
);

OAI21xp5_ASAP7_75t_L g1243 ( 
.A1(n_1043),
.A2(n_1071),
.B(n_1090),
.Y(n_1243)
);

AOI21xp5_ASAP7_75t_L g1244 ( 
.A1(n_1023),
.A2(n_1071),
.B(n_826),
.Y(n_1244)
);

AOI21xp33_ASAP7_75t_L g1245 ( 
.A1(n_1090),
.A2(n_1071),
.B(n_1075),
.Y(n_1245)
);

NOR2xp33_ASAP7_75t_L g1246 ( 
.A(n_1007),
.B(n_350),
.Y(n_1246)
);

OR2x2_ASAP7_75t_L g1247 ( 
.A(n_1066),
.B(n_1073),
.Y(n_1247)
);

INVx3_ASAP7_75t_L g1248 ( 
.A(n_1014),
.Y(n_1248)
);

AOI21xp5_ASAP7_75t_L g1249 ( 
.A1(n_1071),
.A2(n_826),
.B(n_819),
.Y(n_1249)
);

BUFx2_ASAP7_75t_L g1250 ( 
.A(n_1058),
.Y(n_1250)
);

BUFx6f_ASAP7_75t_L g1251 ( 
.A(n_1107),
.Y(n_1251)
);

AOI21xp5_ASAP7_75t_L g1252 ( 
.A1(n_1071),
.A2(n_826),
.B(n_819),
.Y(n_1252)
);

AND2x4_ASAP7_75t_L g1253 ( 
.A(n_1107),
.B(n_872),
.Y(n_1253)
);

OAI21x1_ASAP7_75t_L g1254 ( 
.A1(n_1085),
.A2(n_1046),
.B(n_1162),
.Y(n_1254)
);

INVx3_ASAP7_75t_L g1255 ( 
.A(n_1014),
.Y(n_1255)
);

OAI21x1_ASAP7_75t_L g1256 ( 
.A1(n_1085),
.A2(n_1046),
.B(n_1162),
.Y(n_1256)
);

NAND2xp5_ASAP7_75t_SL g1257 ( 
.A(n_1090),
.B(n_971),
.Y(n_1257)
);

A2O1A1Ixp33_ASAP7_75t_L g1258 ( 
.A1(n_1071),
.A2(n_826),
.B(n_963),
.C(n_971),
.Y(n_1258)
);

INVx2_ASAP7_75t_L g1259 ( 
.A(n_1009),
.Y(n_1259)
);

INVx1_ASAP7_75t_L g1260 ( 
.A(n_1016),
.Y(n_1260)
);

NAND2xp5_ASAP7_75t_L g1261 ( 
.A(n_1071),
.B(n_826),
.Y(n_1261)
);

BUFx12f_ASAP7_75t_L g1262 ( 
.A(n_1058),
.Y(n_1262)
);

NAND2xp5_ASAP7_75t_L g1263 ( 
.A(n_1071),
.B(n_826),
.Y(n_1263)
);

AOI21xp5_ASAP7_75t_L g1264 ( 
.A1(n_1071),
.A2(n_826),
.B(n_819),
.Y(n_1264)
);

INVx2_ASAP7_75t_L g1265 ( 
.A(n_1009),
.Y(n_1265)
);

OAI21xp5_ASAP7_75t_L g1266 ( 
.A1(n_1071),
.A2(n_1090),
.B(n_826),
.Y(n_1266)
);

AOI21xp5_ASAP7_75t_SL g1267 ( 
.A1(n_1071),
.A2(n_1090),
.B(n_867),
.Y(n_1267)
);

OAI21xp5_ASAP7_75t_L g1268 ( 
.A1(n_1071),
.A2(n_1090),
.B(n_826),
.Y(n_1268)
);

NAND2xp5_ASAP7_75t_L g1269 ( 
.A(n_1071),
.B(n_826),
.Y(n_1269)
);

NAND2xp5_ASAP7_75t_L g1270 ( 
.A(n_1066),
.B(n_826),
.Y(n_1270)
);

INVx1_ASAP7_75t_L g1271 ( 
.A(n_1016),
.Y(n_1271)
);

NAND2xp5_ASAP7_75t_L g1272 ( 
.A(n_1066),
.B(n_826),
.Y(n_1272)
);

INVx1_ASAP7_75t_L g1273 ( 
.A(n_1016),
.Y(n_1273)
);

INVx1_ASAP7_75t_L g1274 ( 
.A(n_1016),
.Y(n_1274)
);

NAND3xp33_ASAP7_75t_L g1275 ( 
.A(n_1071),
.B(n_1059),
.C(n_826),
.Y(n_1275)
);

INVx1_ASAP7_75t_L g1276 ( 
.A(n_1016),
.Y(n_1276)
);

OAI21xp5_ASAP7_75t_L g1277 ( 
.A1(n_1071),
.A2(n_1090),
.B(n_826),
.Y(n_1277)
);

INVx3_ASAP7_75t_L g1278 ( 
.A(n_1014),
.Y(n_1278)
);

BUFx3_ASAP7_75t_L g1279 ( 
.A(n_1058),
.Y(n_1279)
);

CKINVDCx11_ASAP7_75t_R g1280 ( 
.A(n_1122),
.Y(n_1280)
);

NAND2x1p5_ASAP7_75t_L g1281 ( 
.A(n_1084),
.B(n_928),
.Y(n_1281)
);

INVx2_ASAP7_75t_L g1282 ( 
.A(n_1009),
.Y(n_1282)
);

OAI21x1_ASAP7_75t_L g1283 ( 
.A1(n_1085),
.A2(n_1046),
.B(n_1162),
.Y(n_1283)
);

AOI21xp5_ASAP7_75t_L g1284 ( 
.A1(n_1071),
.A2(n_826),
.B(n_819),
.Y(n_1284)
);

NOR2xp67_ASAP7_75t_L g1285 ( 
.A(n_1007),
.B(n_715),
.Y(n_1285)
);

AOI21x1_ASAP7_75t_L g1286 ( 
.A1(n_1105),
.A2(n_1085),
.B(n_1072),
.Y(n_1286)
);

INVx1_ASAP7_75t_SL g1287 ( 
.A(n_1073),
.Y(n_1287)
);

NAND2xp5_ASAP7_75t_L g1288 ( 
.A(n_1066),
.B(n_826),
.Y(n_1288)
);

NAND3xp33_ASAP7_75t_L g1289 ( 
.A(n_1071),
.B(n_1059),
.C(n_826),
.Y(n_1289)
);

OAI21x1_ASAP7_75t_L g1290 ( 
.A1(n_1085),
.A2(n_1046),
.B(n_1162),
.Y(n_1290)
);

INVxp67_ASAP7_75t_L g1291 ( 
.A(n_1049),
.Y(n_1291)
);

CKINVDCx5p33_ASAP7_75t_R g1292 ( 
.A(n_1058),
.Y(n_1292)
);

O2A1O1Ixp33_ASAP7_75t_L g1293 ( 
.A1(n_1071),
.A2(n_654),
.B(n_826),
.C(n_971),
.Y(n_1293)
);

AND2x6_ASAP7_75t_L g1294 ( 
.A(n_1083),
.B(n_1159),
.Y(n_1294)
);

OAI21xp5_ASAP7_75t_L g1295 ( 
.A1(n_1071),
.A2(n_1090),
.B(n_826),
.Y(n_1295)
);

OA21x2_ASAP7_75t_L g1296 ( 
.A1(n_1071),
.A2(n_1105),
.B(n_1085),
.Y(n_1296)
);

A2O1A1Ixp33_ASAP7_75t_L g1297 ( 
.A1(n_1071),
.A2(n_826),
.B(n_963),
.C(n_971),
.Y(n_1297)
);

NAND2xp5_ASAP7_75t_L g1298 ( 
.A(n_1071),
.B(n_826),
.Y(n_1298)
);

INVx2_ASAP7_75t_SL g1299 ( 
.A(n_1058),
.Y(n_1299)
);

INVx3_ASAP7_75t_SL g1300 ( 
.A(n_1153),
.Y(n_1300)
);

OAI21x1_ASAP7_75t_L g1301 ( 
.A1(n_1085),
.A2(n_1046),
.B(n_1162),
.Y(n_1301)
);

OAI21x1_ASAP7_75t_L g1302 ( 
.A1(n_1085),
.A2(n_1046),
.B(n_1162),
.Y(n_1302)
);

O2A1O1Ixp33_ASAP7_75t_SL g1303 ( 
.A1(n_1071),
.A2(n_826),
.B(n_971),
.C(n_1091),
.Y(n_1303)
);

BUFx3_ASAP7_75t_L g1304 ( 
.A(n_1058),
.Y(n_1304)
);

INVx2_ASAP7_75t_L g1305 ( 
.A(n_1009),
.Y(n_1305)
);

NAND2xp5_ASAP7_75t_L g1306 ( 
.A(n_1066),
.B(n_826),
.Y(n_1306)
);

NAND2xp5_ASAP7_75t_L g1307 ( 
.A(n_1066),
.B(n_826),
.Y(n_1307)
);

INVx1_ASAP7_75t_L g1308 ( 
.A(n_1016),
.Y(n_1308)
);

NAND2xp5_ASAP7_75t_SL g1309 ( 
.A(n_1090),
.B(n_971),
.Y(n_1309)
);

NAND3xp33_ASAP7_75t_L g1310 ( 
.A(n_1071),
.B(n_1059),
.C(n_826),
.Y(n_1310)
);

INVx4_ASAP7_75t_L g1311 ( 
.A(n_1153),
.Y(n_1311)
);

AO31x2_ASAP7_75t_L g1312 ( 
.A1(n_1127),
.A2(n_1071),
.A3(n_1078),
.B(n_1085),
.Y(n_1312)
);

OAI21xp5_ASAP7_75t_SL g1313 ( 
.A1(n_1050),
.A2(n_654),
.B(n_908),
.Y(n_1313)
);

AND2x2_ASAP7_75t_L g1314 ( 
.A(n_1018),
.B(n_696),
.Y(n_1314)
);

BUFx6f_ASAP7_75t_L g1315 ( 
.A(n_1107),
.Y(n_1315)
);

AOI21xp5_ASAP7_75t_L g1316 ( 
.A1(n_1071),
.A2(n_826),
.B(n_819),
.Y(n_1316)
);

INVx1_ASAP7_75t_L g1317 ( 
.A(n_1016),
.Y(n_1317)
);

AO21x2_ASAP7_75t_L g1318 ( 
.A1(n_1167),
.A2(n_1186),
.B(n_1176),
.Y(n_1318)
);

OAI21xp5_ASAP7_75t_L g1319 ( 
.A1(n_1266),
.A2(n_1277),
.B(n_1268),
.Y(n_1319)
);

OAI22xp33_ASAP7_75t_L g1320 ( 
.A1(n_1275),
.A2(n_1289),
.B1(n_1310),
.B2(n_1263),
.Y(n_1320)
);

INVx3_ASAP7_75t_L g1321 ( 
.A(n_1197),
.Y(n_1321)
);

AOI21x1_ASAP7_75t_L g1322 ( 
.A1(n_1194),
.A2(n_1286),
.B(n_1257),
.Y(n_1322)
);

OAI21x1_ASAP7_75t_L g1323 ( 
.A1(n_1290),
.A2(n_1302),
.B(n_1301),
.Y(n_1323)
);

AOI221xp5_ASAP7_75t_L g1324 ( 
.A1(n_1293),
.A2(n_1245),
.B1(n_1277),
.B2(n_1268),
.C(n_1295),
.Y(n_1324)
);

AOI22xp33_ASAP7_75t_L g1325 ( 
.A1(n_1183),
.A2(n_1275),
.B1(n_1289),
.B2(n_1310),
.Y(n_1325)
);

OAI21x1_ASAP7_75t_L g1326 ( 
.A1(n_1178),
.A2(n_1179),
.B(n_1181),
.Y(n_1326)
);

AO21x2_ASAP7_75t_L g1327 ( 
.A1(n_1186),
.A2(n_1211),
.B(n_1182),
.Y(n_1327)
);

INVx2_ASAP7_75t_SL g1328 ( 
.A(n_1300),
.Y(n_1328)
);

AOI21xp5_ASAP7_75t_L g1329 ( 
.A1(n_1266),
.A2(n_1295),
.B(n_1267),
.Y(n_1329)
);

BUFx2_ASAP7_75t_L g1330 ( 
.A(n_1311),
.Y(n_1330)
);

AOI21xp33_ASAP7_75t_L g1331 ( 
.A1(n_1183),
.A2(n_1214),
.B(n_1209),
.Y(n_1331)
);

OAI21x1_ASAP7_75t_L g1332 ( 
.A1(n_1172),
.A2(n_1171),
.B(n_1170),
.Y(n_1332)
);

INVx1_ASAP7_75t_L g1333 ( 
.A(n_1166),
.Y(n_1333)
);

INVx1_ASAP7_75t_L g1334 ( 
.A(n_1173),
.Y(n_1334)
);

INVx1_ASAP7_75t_L g1335 ( 
.A(n_1184),
.Y(n_1335)
);

INVx1_ASAP7_75t_SL g1336 ( 
.A(n_1198),
.Y(n_1336)
);

INVx1_ASAP7_75t_L g1337 ( 
.A(n_1188),
.Y(n_1337)
);

INVx2_ASAP7_75t_L g1338 ( 
.A(n_1233),
.Y(n_1338)
);

BUFx3_ASAP7_75t_L g1339 ( 
.A(n_1228),
.Y(n_1339)
);

AND2x2_ASAP7_75t_L g1340 ( 
.A(n_1174),
.B(n_1314),
.Y(n_1340)
);

INVx2_ASAP7_75t_L g1341 ( 
.A(n_1215),
.Y(n_1341)
);

OAI22xp33_ASAP7_75t_L g1342 ( 
.A1(n_1261),
.A2(n_1263),
.B1(n_1269),
.B2(n_1298),
.Y(n_1342)
);

AOI22xp33_ASAP7_75t_SL g1343 ( 
.A1(n_1294),
.A2(n_1243),
.B1(n_1219),
.B2(n_1214),
.Y(n_1343)
);

NAND2xp5_ASAP7_75t_L g1344 ( 
.A(n_1270),
.B(n_1272),
.Y(n_1344)
);

INVx1_ASAP7_75t_L g1345 ( 
.A(n_1193),
.Y(n_1345)
);

INVx1_ASAP7_75t_L g1346 ( 
.A(n_1201),
.Y(n_1346)
);

OAI21x1_ASAP7_75t_L g1347 ( 
.A1(n_1187),
.A2(n_1200),
.B(n_1165),
.Y(n_1347)
);

INVx2_ASAP7_75t_L g1348 ( 
.A(n_1215),
.Y(n_1348)
);

OAI22xp5_ASAP7_75t_L g1349 ( 
.A1(n_1261),
.A2(n_1298),
.B1(n_1269),
.B2(n_1175),
.Y(n_1349)
);

OAI21x1_ASAP7_75t_L g1350 ( 
.A1(n_1202),
.A2(n_1218),
.B(n_1296),
.Y(n_1350)
);

OAI21xp5_ASAP7_75t_L g1351 ( 
.A1(n_1244),
.A2(n_1284),
.B(n_1264),
.Y(n_1351)
);

OA21x2_ASAP7_75t_L g1352 ( 
.A1(n_1245),
.A2(n_1243),
.B(n_1190),
.Y(n_1352)
);

CKINVDCx5p33_ASAP7_75t_R g1353 ( 
.A(n_1262),
.Y(n_1353)
);

CKINVDCx20_ASAP7_75t_R g1354 ( 
.A(n_1280),
.Y(n_1354)
);

AOI22xp33_ASAP7_75t_L g1355 ( 
.A1(n_1309),
.A2(n_1294),
.B1(n_1288),
.B2(n_1306),
.Y(n_1355)
);

BUFx4f_ASAP7_75t_SL g1356 ( 
.A(n_1191),
.Y(n_1356)
);

OAI21x1_ASAP7_75t_L g1357 ( 
.A1(n_1296),
.A2(n_1177),
.B(n_1190),
.Y(n_1357)
);

INVx1_ASAP7_75t_L g1358 ( 
.A(n_1212),
.Y(n_1358)
);

INVx1_ASAP7_75t_L g1359 ( 
.A(n_1260),
.Y(n_1359)
);

INVx1_ASAP7_75t_L g1360 ( 
.A(n_1271),
.Y(n_1360)
);

OAI21x1_ASAP7_75t_L g1361 ( 
.A1(n_1177),
.A2(n_1195),
.B(n_1235),
.Y(n_1361)
);

INVx1_ASAP7_75t_L g1362 ( 
.A(n_1273),
.Y(n_1362)
);

AOI22xp5_ASAP7_75t_L g1363 ( 
.A1(n_1246),
.A2(n_1313),
.B1(n_1216),
.B2(n_1219),
.Y(n_1363)
);

AND2x2_ASAP7_75t_L g1364 ( 
.A(n_1247),
.B(n_1205),
.Y(n_1364)
);

INVx1_ASAP7_75t_L g1365 ( 
.A(n_1274),
.Y(n_1365)
);

AO22x2_ASAP7_75t_L g1366 ( 
.A1(n_1313),
.A2(n_1224),
.B1(n_1213),
.B2(n_1220),
.Y(n_1366)
);

AND2x2_ASAP7_75t_L g1367 ( 
.A(n_1205),
.B(n_1287),
.Y(n_1367)
);

INVx1_ASAP7_75t_L g1368 ( 
.A(n_1276),
.Y(n_1368)
);

OR2x2_ASAP7_75t_L g1369 ( 
.A(n_1199),
.B(n_1287),
.Y(n_1369)
);

OA21x2_ASAP7_75t_L g1370 ( 
.A1(n_1249),
.A2(n_1252),
.B(n_1316),
.Y(n_1370)
);

NAND2xp5_ASAP7_75t_L g1371 ( 
.A(n_1307),
.B(n_1258),
.Y(n_1371)
);

AO21x2_ASAP7_75t_L g1372 ( 
.A1(n_1185),
.A2(n_1203),
.B(n_1206),
.Y(n_1372)
);

INVx2_ASAP7_75t_L g1373 ( 
.A(n_1215),
.Y(n_1373)
);

AOI22xp33_ASAP7_75t_SL g1374 ( 
.A1(n_1294),
.A2(n_1225),
.B1(n_1169),
.B2(n_1241),
.Y(n_1374)
);

INVx2_ASAP7_75t_L g1375 ( 
.A(n_1230),
.Y(n_1375)
);

OAI21x1_ASAP7_75t_L g1376 ( 
.A1(n_1208),
.A2(n_1168),
.B(n_1236),
.Y(n_1376)
);

OAI21x1_ASAP7_75t_L g1377 ( 
.A1(n_1241),
.A2(n_1281),
.B(n_1237),
.Y(n_1377)
);

OA21x2_ASAP7_75t_L g1378 ( 
.A1(n_1297),
.A2(n_1223),
.B(n_1229),
.Y(n_1378)
);

OAI22xp5_ASAP7_75t_L g1379 ( 
.A1(n_1291),
.A2(n_1222),
.B1(n_1311),
.B2(n_1210),
.Y(n_1379)
);

OAI21x1_ASAP7_75t_L g1380 ( 
.A1(n_1281),
.A2(n_1237),
.B(n_1240),
.Y(n_1380)
);

OAI222xp33_ASAP7_75t_L g1381 ( 
.A1(n_1232),
.A2(n_1226),
.B1(n_1265),
.B2(n_1305),
.C1(n_1259),
.C2(n_1282),
.Y(n_1381)
);

AO21x2_ASAP7_75t_L g1382 ( 
.A1(n_1185),
.A2(n_1317),
.B(n_1308),
.Y(n_1382)
);

OAI21x1_ASAP7_75t_L g1383 ( 
.A1(n_1240),
.A2(n_1278),
.B(n_1180),
.Y(n_1383)
);

OAI21x1_ASAP7_75t_SL g1384 ( 
.A1(n_1234),
.A2(n_1299),
.B(n_1303),
.Y(n_1384)
);

OAI21x1_ASAP7_75t_L g1385 ( 
.A1(n_1180),
.A2(n_1255),
.B(n_1278),
.Y(n_1385)
);

BUFx6f_ASAP7_75t_L g1386 ( 
.A(n_1164),
.Y(n_1386)
);

OAI21x1_ASAP7_75t_L g1387 ( 
.A1(n_1204),
.A2(n_1255),
.B(n_1248),
.Y(n_1387)
);

OAI22xp5_ASAP7_75t_L g1388 ( 
.A1(n_1285),
.A2(n_1216),
.B1(n_1221),
.B2(n_1250),
.Y(n_1388)
);

OAI21x1_ASAP7_75t_L g1389 ( 
.A1(n_1204),
.A2(n_1248),
.B(n_1231),
.Y(n_1389)
);

AOI21x1_ASAP7_75t_L g1390 ( 
.A1(n_1227),
.A2(n_1238),
.B(n_1253),
.Y(n_1390)
);

BUFx2_ASAP7_75t_SL g1391 ( 
.A(n_1279),
.Y(n_1391)
);

INVxp67_ASAP7_75t_SL g1392 ( 
.A(n_1164),
.Y(n_1392)
);

OAI22xp33_ASAP7_75t_L g1393 ( 
.A1(n_1304),
.A2(n_1315),
.B1(n_1192),
.B2(n_1251),
.Y(n_1393)
);

OAI22xp5_ASAP7_75t_SL g1394 ( 
.A1(n_1292),
.A2(n_1196),
.B1(n_1192),
.B2(n_1251),
.Y(n_1394)
);

OAI21x1_ASAP7_75t_L g1395 ( 
.A1(n_1312),
.A2(n_1242),
.B(n_1207),
.Y(n_1395)
);

OAI21x1_ASAP7_75t_L g1396 ( 
.A1(n_1312),
.A2(n_1242),
.B(n_1207),
.Y(n_1396)
);

INVx1_ASAP7_75t_L g1397 ( 
.A(n_1230),
.Y(n_1397)
);

OAI21x1_ASAP7_75t_L g1398 ( 
.A1(n_1242),
.A2(n_1207),
.B(n_1217),
.Y(n_1398)
);

NOR2xp33_ASAP7_75t_L g1399 ( 
.A(n_1198),
.B(n_1251),
.Y(n_1399)
);

NOR2xp67_ASAP7_75t_L g1400 ( 
.A(n_1217),
.B(n_1189),
.Y(n_1400)
);

CKINVDCx20_ASAP7_75t_R g1401 ( 
.A(n_1189),
.Y(n_1401)
);

INVx5_ASAP7_75t_L g1402 ( 
.A(n_1197),
.Y(n_1402)
);

NOR2xp33_ASAP7_75t_L g1403 ( 
.A(n_1275),
.B(n_908),
.Y(n_1403)
);

AND2x2_ASAP7_75t_L g1404 ( 
.A(n_1174),
.B(n_1314),
.Y(n_1404)
);

OAI21x1_ASAP7_75t_L g1405 ( 
.A1(n_1181),
.A2(n_1256),
.B(n_1254),
.Y(n_1405)
);

INVx2_ASAP7_75t_L g1406 ( 
.A(n_1233),
.Y(n_1406)
);

INVx1_ASAP7_75t_L g1407 ( 
.A(n_1166),
.Y(n_1407)
);

AOI21xp5_ASAP7_75t_L g1408 ( 
.A1(n_1266),
.A2(n_1277),
.B(n_1268),
.Y(n_1408)
);

AND2x2_ASAP7_75t_L g1409 ( 
.A(n_1174),
.B(n_1314),
.Y(n_1409)
);

OAI21x1_ASAP7_75t_L g1410 ( 
.A1(n_1254),
.A2(n_1283),
.B(n_1256),
.Y(n_1410)
);

CKINVDCx20_ASAP7_75t_R g1411 ( 
.A(n_1280),
.Y(n_1411)
);

OAI21x1_ASAP7_75t_L g1412 ( 
.A1(n_1254),
.A2(n_1283),
.B(n_1256),
.Y(n_1412)
);

NAND2xp5_ASAP7_75t_L g1413 ( 
.A(n_1270),
.B(n_1272),
.Y(n_1413)
);

INVx2_ASAP7_75t_L g1414 ( 
.A(n_1233),
.Y(n_1414)
);

AND2x4_ASAP7_75t_L g1415 ( 
.A(n_1197),
.B(n_1239),
.Y(n_1415)
);

INVx2_ASAP7_75t_L g1416 ( 
.A(n_1233),
.Y(n_1416)
);

AND2x2_ASAP7_75t_L g1417 ( 
.A(n_1174),
.B(n_1314),
.Y(n_1417)
);

AO21x2_ASAP7_75t_L g1418 ( 
.A1(n_1167),
.A2(n_1186),
.B(n_1176),
.Y(n_1418)
);

HB1xp67_ASAP7_75t_L g1419 ( 
.A(n_1312),
.Y(n_1419)
);

INVx1_ASAP7_75t_L g1420 ( 
.A(n_1166),
.Y(n_1420)
);

INVx2_ASAP7_75t_SL g1421 ( 
.A(n_1300),
.Y(n_1421)
);

CKINVDCx16_ASAP7_75t_R g1422 ( 
.A(n_1262),
.Y(n_1422)
);

OAI21x1_ASAP7_75t_L g1423 ( 
.A1(n_1254),
.A2(n_1283),
.B(n_1256),
.Y(n_1423)
);

OAI21x1_ASAP7_75t_L g1424 ( 
.A1(n_1254),
.A2(n_1283),
.B(n_1256),
.Y(n_1424)
);

HB1xp67_ASAP7_75t_L g1425 ( 
.A(n_1312),
.Y(n_1425)
);

BUFx2_ASAP7_75t_SL g1426 ( 
.A(n_1228),
.Y(n_1426)
);

INVx3_ASAP7_75t_L g1427 ( 
.A(n_1197),
.Y(n_1427)
);

OAI21x1_ASAP7_75t_L g1428 ( 
.A1(n_1254),
.A2(n_1283),
.B(n_1256),
.Y(n_1428)
);

AO21x2_ASAP7_75t_L g1429 ( 
.A1(n_1167),
.A2(n_1186),
.B(n_1176),
.Y(n_1429)
);

INVx1_ASAP7_75t_L g1430 ( 
.A(n_1166),
.Y(n_1430)
);

AND2x4_ASAP7_75t_L g1431 ( 
.A(n_1197),
.B(n_1239),
.Y(n_1431)
);

OAI21x1_ASAP7_75t_L g1432 ( 
.A1(n_1254),
.A2(n_1283),
.B(n_1256),
.Y(n_1432)
);

NAND2xp5_ASAP7_75t_L g1433 ( 
.A(n_1270),
.B(n_1272),
.Y(n_1433)
);

INVx1_ASAP7_75t_L g1434 ( 
.A(n_1166),
.Y(n_1434)
);

NAND2x1p5_ASAP7_75t_L g1435 ( 
.A(n_1197),
.B(n_1084),
.Y(n_1435)
);

AO21x1_ASAP7_75t_L g1436 ( 
.A1(n_1257),
.A2(n_1309),
.B(n_1268),
.Y(n_1436)
);

OAI21xp5_ASAP7_75t_L g1437 ( 
.A1(n_1266),
.A2(n_1071),
.B(n_971),
.Y(n_1437)
);

AOI21xp5_ASAP7_75t_L g1438 ( 
.A1(n_1266),
.A2(n_1277),
.B(n_1268),
.Y(n_1438)
);

OAI21x1_ASAP7_75t_L g1439 ( 
.A1(n_1254),
.A2(n_1283),
.B(n_1256),
.Y(n_1439)
);

NAND2x1p5_ASAP7_75t_L g1440 ( 
.A(n_1197),
.B(n_1084),
.Y(n_1440)
);

INVx2_ASAP7_75t_SL g1441 ( 
.A(n_1300),
.Y(n_1441)
);

NOR2xp33_ASAP7_75t_L g1442 ( 
.A(n_1275),
.B(n_908),
.Y(n_1442)
);

INVx1_ASAP7_75t_L g1443 ( 
.A(n_1166),
.Y(n_1443)
);

OAI21x1_ASAP7_75t_L g1444 ( 
.A1(n_1181),
.A2(n_1256),
.B(n_1254),
.Y(n_1444)
);

OAI21x1_ASAP7_75t_L g1445 ( 
.A1(n_1181),
.A2(n_1256),
.B(n_1254),
.Y(n_1445)
);

INVx1_ASAP7_75t_L g1446 ( 
.A(n_1166),
.Y(n_1446)
);

OAI21x1_ASAP7_75t_L g1447 ( 
.A1(n_1254),
.A2(n_1283),
.B(n_1256),
.Y(n_1447)
);

NOR2xp33_ASAP7_75t_L g1448 ( 
.A(n_1275),
.B(n_908),
.Y(n_1448)
);

OAI21x1_ASAP7_75t_L g1449 ( 
.A1(n_1254),
.A2(n_1283),
.B(n_1256),
.Y(n_1449)
);

INVx1_ASAP7_75t_L g1450 ( 
.A(n_1166),
.Y(n_1450)
);

OAI21x1_ASAP7_75t_L g1451 ( 
.A1(n_1254),
.A2(n_1283),
.B(n_1256),
.Y(n_1451)
);

AND2x2_ASAP7_75t_L g1452 ( 
.A(n_1340),
.B(n_1404),
.Y(n_1452)
);

AND2x2_ASAP7_75t_L g1453 ( 
.A(n_1409),
.B(n_1417),
.Y(n_1453)
);

NAND2xp5_ASAP7_75t_L g1454 ( 
.A(n_1344),
.B(n_1413),
.Y(n_1454)
);

NAND2xp5_ASAP7_75t_L g1455 ( 
.A(n_1433),
.B(n_1364),
.Y(n_1455)
);

AND2x2_ASAP7_75t_L g1456 ( 
.A(n_1367),
.B(n_1366),
.Y(n_1456)
);

BUFx12f_ASAP7_75t_L g1457 ( 
.A(n_1353),
.Y(n_1457)
);

OAI22xp5_ASAP7_75t_L g1458 ( 
.A1(n_1325),
.A2(n_1329),
.B1(n_1408),
.B2(n_1438),
.Y(n_1458)
);

AND2x2_ASAP7_75t_L g1459 ( 
.A(n_1366),
.B(n_1363),
.Y(n_1459)
);

O2A1O1Ixp5_ASAP7_75t_L g1460 ( 
.A1(n_1319),
.A2(n_1351),
.B(n_1436),
.C(n_1320),
.Y(n_1460)
);

INVx3_ASAP7_75t_L g1461 ( 
.A(n_1389),
.Y(n_1461)
);

NAND2xp5_ASAP7_75t_L g1462 ( 
.A(n_1369),
.B(n_1349),
.Y(n_1462)
);

AND2x2_ASAP7_75t_L g1463 ( 
.A(n_1366),
.B(n_1321),
.Y(n_1463)
);

BUFx3_ASAP7_75t_L g1464 ( 
.A(n_1356),
.Y(n_1464)
);

OA21x2_ASAP7_75t_L g1465 ( 
.A1(n_1347),
.A2(n_1396),
.B(n_1395),
.Y(n_1465)
);

OAI22xp5_ASAP7_75t_L g1466 ( 
.A1(n_1325),
.A2(n_1324),
.B1(n_1320),
.B2(n_1343),
.Y(n_1466)
);

O2A1O1Ixp33_ASAP7_75t_L g1467 ( 
.A1(n_1437),
.A2(n_1448),
.B(n_1442),
.C(n_1403),
.Y(n_1467)
);

OAI31xp33_ASAP7_75t_L g1468 ( 
.A1(n_1331),
.A2(n_1403),
.A3(n_1442),
.B(n_1448),
.Y(n_1468)
);

AOI21xp5_ASAP7_75t_L g1469 ( 
.A1(n_1342),
.A2(n_1370),
.B(n_1352),
.Y(n_1469)
);

NAND2xp5_ASAP7_75t_L g1470 ( 
.A(n_1371),
.B(n_1342),
.Y(n_1470)
);

INVx6_ASAP7_75t_L g1471 ( 
.A(n_1402),
.Y(n_1471)
);

AOI21xp5_ASAP7_75t_SL g1472 ( 
.A1(n_1388),
.A2(n_1378),
.B(n_1352),
.Y(n_1472)
);

O2A1O1Ixp5_ASAP7_75t_L g1473 ( 
.A1(n_1322),
.A2(n_1379),
.B(n_1419),
.C(n_1425),
.Y(n_1473)
);

A2O1A1Ixp33_ASAP7_75t_L g1474 ( 
.A1(n_1355),
.A2(n_1398),
.B(n_1400),
.C(n_1396),
.Y(n_1474)
);

AND2x2_ASAP7_75t_L g1475 ( 
.A(n_1427),
.B(n_1355),
.Y(n_1475)
);

AOI21xp5_ASAP7_75t_L g1476 ( 
.A1(n_1370),
.A2(n_1352),
.B(n_1347),
.Y(n_1476)
);

INVx1_ASAP7_75t_L g1477 ( 
.A(n_1333),
.Y(n_1477)
);

BUFx6f_ASAP7_75t_L g1478 ( 
.A(n_1386),
.Y(n_1478)
);

OA21x2_ASAP7_75t_L g1479 ( 
.A1(n_1326),
.A2(n_1395),
.B(n_1350),
.Y(n_1479)
);

AOI21xp5_ASAP7_75t_SL g1480 ( 
.A1(n_1378),
.A2(n_1399),
.B(n_1393),
.Y(n_1480)
);

AOI21xp5_ASAP7_75t_SL g1481 ( 
.A1(n_1378),
.A2(n_1399),
.B(n_1393),
.Y(n_1481)
);

NAND2xp5_ASAP7_75t_L g1482 ( 
.A(n_1334),
.B(n_1335),
.Y(n_1482)
);

INVx1_ASAP7_75t_L g1483 ( 
.A(n_1337),
.Y(n_1483)
);

AOI21xp5_ASAP7_75t_L g1484 ( 
.A1(n_1370),
.A2(n_1327),
.B(n_1429),
.Y(n_1484)
);

AND2x2_ASAP7_75t_L g1485 ( 
.A(n_1345),
.B(n_1346),
.Y(n_1485)
);

INVx3_ASAP7_75t_L g1486 ( 
.A(n_1380),
.Y(n_1486)
);

OR2x2_ASAP7_75t_L g1487 ( 
.A(n_1358),
.B(n_1359),
.Y(n_1487)
);

INVx2_ASAP7_75t_SL g1488 ( 
.A(n_1339),
.Y(n_1488)
);

OAI22xp5_ASAP7_75t_L g1489 ( 
.A1(n_1336),
.A2(n_1339),
.B1(n_1374),
.B2(n_1330),
.Y(n_1489)
);

INVx3_ASAP7_75t_SL g1490 ( 
.A(n_1353),
.Y(n_1490)
);

NAND2xp5_ASAP7_75t_L g1491 ( 
.A(n_1360),
.B(n_1362),
.Y(n_1491)
);

OAI22xp5_ASAP7_75t_L g1492 ( 
.A1(n_1426),
.A2(n_1441),
.B1(n_1421),
.B2(n_1328),
.Y(n_1492)
);

NAND2xp5_ASAP7_75t_L g1493 ( 
.A(n_1365),
.B(n_1368),
.Y(n_1493)
);

O2A1O1Ixp33_ASAP7_75t_L g1494 ( 
.A1(n_1384),
.A2(n_1318),
.B(n_1418),
.C(n_1446),
.Y(n_1494)
);

NAND2xp5_ASAP7_75t_L g1495 ( 
.A(n_1407),
.B(n_1420),
.Y(n_1495)
);

AND2x2_ASAP7_75t_L g1496 ( 
.A(n_1430),
.B(n_1434),
.Y(n_1496)
);

NAND2xp5_ASAP7_75t_L g1497 ( 
.A(n_1443),
.B(n_1450),
.Y(n_1497)
);

AOI21xp5_ASAP7_75t_L g1498 ( 
.A1(n_1418),
.A2(n_1350),
.B(n_1323),
.Y(n_1498)
);

OAI22xp5_ASAP7_75t_L g1499 ( 
.A1(n_1356),
.A2(n_1391),
.B1(n_1402),
.B2(n_1411),
.Y(n_1499)
);

OAI22xp5_ASAP7_75t_L g1500 ( 
.A1(n_1402),
.A2(n_1411),
.B1(n_1354),
.B2(n_1422),
.Y(n_1500)
);

OAI22xp5_ASAP7_75t_L g1501 ( 
.A1(n_1402),
.A2(n_1354),
.B1(n_1435),
.B2(n_1440),
.Y(n_1501)
);

AOI21xp5_ASAP7_75t_SL g1502 ( 
.A1(n_1435),
.A2(n_1440),
.B(n_1372),
.Y(n_1502)
);

NAND2xp5_ASAP7_75t_L g1503 ( 
.A(n_1386),
.B(n_1392),
.Y(n_1503)
);

OA21x2_ASAP7_75t_L g1504 ( 
.A1(n_1326),
.A2(n_1357),
.B(n_1398),
.Y(n_1504)
);

OA22x2_ASAP7_75t_L g1505 ( 
.A1(n_1394),
.A2(n_1377),
.B1(n_1373),
.B2(n_1341),
.Y(n_1505)
);

O2A1O1Ixp5_ASAP7_75t_L g1506 ( 
.A1(n_1390),
.A2(n_1373),
.B(n_1341),
.C(n_1348),
.Y(n_1506)
);

O2A1O1Ixp33_ASAP7_75t_L g1507 ( 
.A1(n_1372),
.A2(n_1381),
.B(n_1348),
.C(n_1401),
.Y(n_1507)
);

INVx1_ASAP7_75t_L g1508 ( 
.A(n_1397),
.Y(n_1508)
);

OAI22xp5_ASAP7_75t_L g1509 ( 
.A1(n_1401),
.A2(n_1386),
.B1(n_1375),
.B2(n_1338),
.Y(n_1509)
);

AND2x2_ASAP7_75t_L g1510 ( 
.A(n_1385),
.B(n_1387),
.Y(n_1510)
);

O2A1O1Ixp33_ASAP7_75t_L g1511 ( 
.A1(n_1406),
.A2(n_1414),
.B(n_1416),
.C(n_1361),
.Y(n_1511)
);

AND2x4_ASAP7_75t_L g1512 ( 
.A(n_1383),
.B(n_1385),
.Y(n_1512)
);

BUFx6f_ASAP7_75t_L g1513 ( 
.A(n_1376),
.Y(n_1513)
);

AOI21xp5_ASAP7_75t_L g1514 ( 
.A1(n_1410),
.A2(n_1439),
.B(n_1449),
.Y(n_1514)
);

AOI211xp5_ASAP7_75t_L g1515 ( 
.A1(n_1332),
.A2(n_1405),
.B(n_1445),
.C(n_1444),
.Y(n_1515)
);

O2A1O1Ixp33_ASAP7_75t_L g1516 ( 
.A1(n_1332),
.A2(n_1412),
.B(n_1423),
.C(n_1424),
.Y(n_1516)
);

AND2x2_ASAP7_75t_L g1517 ( 
.A(n_1412),
.B(n_1423),
.Y(n_1517)
);

AOI21x1_ASAP7_75t_SL g1518 ( 
.A1(n_1424),
.A2(n_1428),
.B(n_1432),
.Y(n_1518)
);

NAND2xp5_ASAP7_75t_L g1519 ( 
.A(n_1428),
.B(n_1451),
.Y(n_1519)
);

HB1xp67_ASAP7_75t_L g1520 ( 
.A(n_1447),
.Y(n_1520)
);

AND2x2_ASAP7_75t_L g1521 ( 
.A(n_1340),
.B(n_1404),
.Y(n_1521)
);

BUFx3_ASAP7_75t_L g1522 ( 
.A(n_1356),
.Y(n_1522)
);

NAND2xp5_ASAP7_75t_L g1523 ( 
.A(n_1344),
.B(n_1413),
.Y(n_1523)
);

OA21x2_ASAP7_75t_L g1524 ( 
.A1(n_1347),
.A2(n_1396),
.B(n_1395),
.Y(n_1524)
);

AND2x6_ASAP7_75t_L g1525 ( 
.A(n_1415),
.B(n_1431),
.Y(n_1525)
);

AND2x2_ASAP7_75t_L g1526 ( 
.A(n_1340),
.B(n_1404),
.Y(n_1526)
);

NAND2x1p5_ASAP7_75t_L g1527 ( 
.A(n_1402),
.B(n_1389),
.Y(n_1527)
);

AND2x2_ASAP7_75t_L g1528 ( 
.A(n_1340),
.B(n_1404),
.Y(n_1528)
);

AND2x2_ASAP7_75t_L g1529 ( 
.A(n_1340),
.B(n_1404),
.Y(n_1529)
);

AND2x2_ASAP7_75t_L g1530 ( 
.A(n_1340),
.B(n_1404),
.Y(n_1530)
);

NAND2xp5_ASAP7_75t_L g1531 ( 
.A(n_1344),
.B(n_1413),
.Y(n_1531)
);

AND2x6_ASAP7_75t_L g1532 ( 
.A(n_1415),
.B(n_1431),
.Y(n_1532)
);

CKINVDCx16_ASAP7_75t_R g1533 ( 
.A(n_1422),
.Y(n_1533)
);

INVx1_ASAP7_75t_SL g1534 ( 
.A(n_1426),
.Y(n_1534)
);

INVx1_ASAP7_75t_L g1535 ( 
.A(n_1333),
.Y(n_1535)
);

HB1xp67_ASAP7_75t_L g1536 ( 
.A(n_1382),
.Y(n_1536)
);

OAI21xp5_ASAP7_75t_L g1537 ( 
.A1(n_1460),
.A2(n_1466),
.B(n_1458),
.Y(n_1537)
);

OAI21x1_ASAP7_75t_L g1538 ( 
.A1(n_1518),
.A2(n_1476),
.B(n_1484),
.Y(n_1538)
);

AO21x1_ASAP7_75t_SL g1539 ( 
.A1(n_1470),
.A2(n_1460),
.B(n_1519),
.Y(n_1539)
);

AND2x2_ASAP7_75t_L g1540 ( 
.A(n_1469),
.B(n_1465),
.Y(n_1540)
);

INVx2_ASAP7_75t_L g1541 ( 
.A(n_1465),
.Y(n_1541)
);

AND2x2_ASAP7_75t_L g1542 ( 
.A(n_1524),
.B(n_1510),
.Y(n_1542)
);

INVx1_ASAP7_75t_L g1543 ( 
.A(n_1508),
.Y(n_1543)
);

OR2x2_ASAP7_75t_L g1544 ( 
.A(n_1462),
.B(n_1459),
.Y(n_1544)
);

INVx2_ASAP7_75t_L g1545 ( 
.A(n_1524),
.Y(n_1545)
);

AND2x2_ASAP7_75t_L g1546 ( 
.A(n_1504),
.B(n_1520),
.Y(n_1546)
);

INVx2_ASAP7_75t_L g1547 ( 
.A(n_1504),
.Y(n_1547)
);

AO21x2_ASAP7_75t_L g1548 ( 
.A1(n_1536),
.A2(n_1498),
.B(n_1472),
.Y(n_1548)
);

OR2x6_ASAP7_75t_L g1549 ( 
.A(n_1527),
.B(n_1502),
.Y(n_1549)
);

INVx1_ASAP7_75t_L g1550 ( 
.A(n_1477),
.Y(n_1550)
);

OR2x2_ASAP7_75t_L g1551 ( 
.A(n_1456),
.B(n_1474),
.Y(n_1551)
);

AND2x2_ASAP7_75t_L g1552 ( 
.A(n_1517),
.B(n_1479),
.Y(n_1552)
);

INVx2_ASAP7_75t_L g1553 ( 
.A(n_1479),
.Y(n_1553)
);

NAND2xp5_ASAP7_75t_L g1554 ( 
.A(n_1485),
.B(n_1496),
.Y(n_1554)
);

INVx1_ASAP7_75t_L g1555 ( 
.A(n_1483),
.Y(n_1555)
);

AOI22xp5_ASAP7_75t_L g1556 ( 
.A1(n_1489),
.A2(n_1475),
.B1(n_1523),
.B2(n_1454),
.Y(n_1556)
);

INVx1_ASAP7_75t_L g1557 ( 
.A(n_1535),
.Y(n_1557)
);

AND2x4_ASAP7_75t_L g1558 ( 
.A(n_1512),
.B(n_1461),
.Y(n_1558)
);

NAND2xp5_ASAP7_75t_L g1559 ( 
.A(n_1482),
.B(n_1491),
.Y(n_1559)
);

BUFx2_ASAP7_75t_L g1560 ( 
.A(n_1512),
.Y(n_1560)
);

BUFx6f_ASAP7_75t_L g1561 ( 
.A(n_1513),
.Y(n_1561)
);

INVx1_ASAP7_75t_L g1562 ( 
.A(n_1493),
.Y(n_1562)
);

OR2x6_ASAP7_75t_L g1563 ( 
.A(n_1471),
.B(n_1507),
.Y(n_1563)
);

BUFx2_ASAP7_75t_L g1564 ( 
.A(n_1486),
.Y(n_1564)
);

OA21x2_ASAP7_75t_L g1565 ( 
.A1(n_1514),
.A2(n_1498),
.B(n_1474),
.Y(n_1565)
);

OR2x6_ASAP7_75t_L g1566 ( 
.A(n_1471),
.B(n_1507),
.Y(n_1566)
);

INVx1_ASAP7_75t_L g1567 ( 
.A(n_1495),
.Y(n_1567)
);

BUFx3_ASAP7_75t_L g1568 ( 
.A(n_1525),
.Y(n_1568)
);

INVx1_ASAP7_75t_L g1569 ( 
.A(n_1497),
.Y(n_1569)
);

INVx1_ASAP7_75t_L g1570 ( 
.A(n_1487),
.Y(n_1570)
);

CKINVDCx20_ASAP7_75t_R g1571 ( 
.A(n_1533),
.Y(n_1571)
);

INVx1_ASAP7_75t_L g1572 ( 
.A(n_1463),
.Y(n_1572)
);

INVx1_ASAP7_75t_L g1573 ( 
.A(n_1511),
.Y(n_1573)
);

NAND2xp5_ASAP7_75t_L g1574 ( 
.A(n_1531),
.B(n_1455),
.Y(n_1574)
);

AO21x2_ASAP7_75t_L g1575 ( 
.A1(n_1511),
.A2(n_1494),
.B(n_1516),
.Y(n_1575)
);

INVx1_ASAP7_75t_L g1576 ( 
.A(n_1494),
.Y(n_1576)
);

INVxp67_ASAP7_75t_L g1577 ( 
.A(n_1503),
.Y(n_1577)
);

INVx1_ASAP7_75t_L g1578 ( 
.A(n_1506),
.Y(n_1578)
);

INVx1_ASAP7_75t_L g1579 ( 
.A(n_1525),
.Y(n_1579)
);

BUFx6f_ASAP7_75t_L g1580 ( 
.A(n_1478),
.Y(n_1580)
);

NAND2xp5_ASAP7_75t_L g1581 ( 
.A(n_1467),
.B(n_1468),
.Y(n_1581)
);

INVx2_ASAP7_75t_L g1582 ( 
.A(n_1505),
.Y(n_1582)
);

HB1xp67_ASAP7_75t_L g1583 ( 
.A(n_1473),
.Y(n_1583)
);

AND2x2_ASAP7_75t_L g1584 ( 
.A(n_1542),
.B(n_1515),
.Y(n_1584)
);

HB1xp67_ASAP7_75t_L g1585 ( 
.A(n_1546),
.Y(n_1585)
);

INVx2_ASAP7_75t_L g1586 ( 
.A(n_1547),
.Y(n_1586)
);

INVx1_ASAP7_75t_L g1587 ( 
.A(n_1543),
.Y(n_1587)
);

HB1xp67_ASAP7_75t_L g1588 ( 
.A(n_1546),
.Y(n_1588)
);

AND2x2_ASAP7_75t_L g1589 ( 
.A(n_1542),
.B(n_1452),
.Y(n_1589)
);

AND2x2_ASAP7_75t_L g1590 ( 
.A(n_1542),
.B(n_1453),
.Y(n_1590)
);

OR2x2_ASAP7_75t_L g1591 ( 
.A(n_1554),
.B(n_1521),
.Y(n_1591)
);

AND2x2_ASAP7_75t_L g1592 ( 
.A(n_1552),
.B(n_1530),
.Y(n_1592)
);

BUFx2_ASAP7_75t_L g1593 ( 
.A(n_1558),
.Y(n_1593)
);

BUFx2_ASAP7_75t_L g1594 ( 
.A(n_1558),
.Y(n_1594)
);

BUFx2_ASAP7_75t_L g1595 ( 
.A(n_1558),
.Y(n_1595)
);

NOR2x1_ASAP7_75t_L g1596 ( 
.A(n_1576),
.B(n_1481),
.Y(n_1596)
);

AND2x2_ASAP7_75t_L g1597 ( 
.A(n_1552),
.B(n_1529),
.Y(n_1597)
);

CKINVDCx20_ASAP7_75t_R g1598 ( 
.A(n_1571),
.Y(n_1598)
);

INVx1_ASAP7_75t_L g1599 ( 
.A(n_1543),
.Y(n_1599)
);

INVx2_ASAP7_75t_L g1600 ( 
.A(n_1541),
.Y(n_1600)
);

AND2x2_ASAP7_75t_L g1601 ( 
.A(n_1552),
.B(n_1526),
.Y(n_1601)
);

AOI22xp5_ASAP7_75t_L g1602 ( 
.A1(n_1581),
.A2(n_1528),
.B1(n_1501),
.B2(n_1532),
.Y(n_1602)
);

BUFx6f_ASAP7_75t_L g1603 ( 
.A(n_1561),
.Y(n_1603)
);

OAI22xp5_ASAP7_75t_L g1604 ( 
.A1(n_1537),
.A2(n_1467),
.B1(n_1488),
.B2(n_1534),
.Y(n_1604)
);

OAI21xp33_ASAP7_75t_L g1605 ( 
.A1(n_1537),
.A2(n_1480),
.B(n_1499),
.Y(n_1605)
);

OR2x2_ASAP7_75t_L g1606 ( 
.A(n_1554),
.B(n_1509),
.Y(n_1606)
);

INVx1_ASAP7_75t_L g1607 ( 
.A(n_1550),
.Y(n_1607)
);

HB1xp67_ASAP7_75t_L g1608 ( 
.A(n_1546),
.Y(n_1608)
);

NOR2x1_ASAP7_75t_L g1609 ( 
.A(n_1576),
.B(n_1500),
.Y(n_1609)
);

OR2x2_ASAP7_75t_L g1610 ( 
.A(n_1551),
.B(n_1544),
.Y(n_1610)
);

BUFx3_ASAP7_75t_L g1611 ( 
.A(n_1568),
.Y(n_1611)
);

INVxp67_ASAP7_75t_L g1612 ( 
.A(n_1539),
.Y(n_1612)
);

AOI22xp33_ASAP7_75t_SL g1613 ( 
.A1(n_1604),
.A2(n_1581),
.B1(n_1582),
.B2(n_1583),
.Y(n_1613)
);

INVx1_ASAP7_75t_L g1614 ( 
.A(n_1587),
.Y(n_1614)
);

AOI221xp5_ASAP7_75t_L g1615 ( 
.A1(n_1604),
.A2(n_1583),
.B1(n_1556),
.B2(n_1540),
.C(n_1578),
.Y(n_1615)
);

OAI33xp33_ASAP7_75t_L g1616 ( 
.A1(n_1610),
.A2(n_1544),
.A3(n_1559),
.B1(n_1574),
.B2(n_1570),
.B3(n_1567),
.Y(n_1616)
);

AOI22xp33_ASAP7_75t_L g1617 ( 
.A1(n_1605),
.A2(n_1582),
.B1(n_1566),
.B2(n_1563),
.Y(n_1617)
);

NAND2xp33_ASAP7_75t_SL g1618 ( 
.A(n_1598),
.B(n_1571),
.Y(n_1618)
);

AND2x2_ASAP7_75t_L g1619 ( 
.A(n_1589),
.B(n_1560),
.Y(n_1619)
);

OR2x2_ASAP7_75t_L g1620 ( 
.A(n_1610),
.B(n_1544),
.Y(n_1620)
);

OA211x2_ASAP7_75t_L g1621 ( 
.A1(n_1605),
.A2(n_1539),
.B(n_1577),
.C(n_1559),
.Y(n_1621)
);

OAI31xp33_ASAP7_75t_L g1622 ( 
.A1(n_1584),
.A2(n_1582),
.A3(n_1540),
.B(n_1578),
.Y(n_1622)
);

OAI22xp5_ASAP7_75t_L g1623 ( 
.A1(n_1609),
.A2(n_1556),
.B1(n_1568),
.B2(n_1579),
.Y(n_1623)
);

HB1xp67_ASAP7_75t_L g1624 ( 
.A(n_1585),
.Y(n_1624)
);

BUFx3_ASAP7_75t_L g1625 ( 
.A(n_1598),
.Y(n_1625)
);

AO21x2_ASAP7_75t_L g1626 ( 
.A1(n_1586),
.A2(n_1540),
.B(n_1573),
.Y(n_1626)
);

NAND2xp5_ASAP7_75t_SL g1627 ( 
.A(n_1609),
.B(n_1574),
.Y(n_1627)
);

OA21x2_ASAP7_75t_L g1628 ( 
.A1(n_1600),
.A2(n_1538),
.B(n_1545),
.Y(n_1628)
);

OR2x2_ASAP7_75t_L g1629 ( 
.A(n_1610),
.B(n_1570),
.Y(n_1629)
);

INVx1_ASAP7_75t_L g1630 ( 
.A(n_1587),
.Y(n_1630)
);

BUFx2_ASAP7_75t_L g1631 ( 
.A(n_1612),
.Y(n_1631)
);

INVx2_ASAP7_75t_L g1632 ( 
.A(n_1600),
.Y(n_1632)
);

INVxp67_ASAP7_75t_SL g1633 ( 
.A(n_1584),
.Y(n_1633)
);

INVx1_ASAP7_75t_L g1634 ( 
.A(n_1599),
.Y(n_1634)
);

HB1xp67_ASAP7_75t_L g1635 ( 
.A(n_1585),
.Y(n_1635)
);

NAND2xp5_ASAP7_75t_L g1636 ( 
.A(n_1589),
.B(n_1562),
.Y(n_1636)
);

OAI211xp5_ASAP7_75t_L g1637 ( 
.A1(n_1612),
.A2(n_1565),
.B(n_1560),
.C(n_1564),
.Y(n_1637)
);

AOI22xp5_ASAP7_75t_L g1638 ( 
.A1(n_1596),
.A2(n_1602),
.B1(n_1532),
.B2(n_1525),
.Y(n_1638)
);

OR2x2_ASAP7_75t_L g1639 ( 
.A(n_1591),
.B(n_1577),
.Y(n_1639)
);

HB1xp67_ASAP7_75t_L g1640 ( 
.A(n_1588),
.Y(n_1640)
);

INVx2_ASAP7_75t_L g1641 ( 
.A(n_1600),
.Y(n_1641)
);

INVx1_ASAP7_75t_L g1642 ( 
.A(n_1599),
.Y(n_1642)
);

INVx4_ASAP7_75t_L g1643 ( 
.A(n_1603),
.Y(n_1643)
);

OR2x2_ASAP7_75t_L g1644 ( 
.A(n_1591),
.B(n_1562),
.Y(n_1644)
);

AOI22xp33_ASAP7_75t_L g1645 ( 
.A1(n_1584),
.A2(n_1563),
.B1(n_1566),
.B2(n_1539),
.Y(n_1645)
);

NOR4xp25_ASAP7_75t_SL g1646 ( 
.A(n_1593),
.B(n_1560),
.C(n_1564),
.D(n_1573),
.Y(n_1646)
);

INVx1_ASAP7_75t_L g1647 ( 
.A(n_1607),
.Y(n_1647)
);

NOR3xp33_ASAP7_75t_SL g1648 ( 
.A(n_1607),
.B(n_1492),
.C(n_1557),
.Y(n_1648)
);

BUFx2_ASAP7_75t_L g1649 ( 
.A(n_1593),
.Y(n_1649)
);

AOI221xp5_ASAP7_75t_L g1650 ( 
.A1(n_1588),
.A2(n_1569),
.B1(n_1567),
.B2(n_1555),
.C(n_1557),
.Y(n_1650)
);

HB1xp67_ASAP7_75t_L g1651 ( 
.A(n_1608),
.Y(n_1651)
);

OAI31xp33_ASAP7_75t_L g1652 ( 
.A1(n_1606),
.A2(n_1569),
.A3(n_1579),
.B(n_1572),
.Y(n_1652)
);

INVx2_ASAP7_75t_L g1653 ( 
.A(n_1626),
.Y(n_1653)
);

INVx1_ASAP7_75t_SL g1654 ( 
.A(n_1625),
.Y(n_1654)
);

INVx2_ASAP7_75t_L g1655 ( 
.A(n_1626),
.Y(n_1655)
);

INVx2_ASAP7_75t_L g1656 ( 
.A(n_1626),
.Y(n_1656)
);

INVx3_ASAP7_75t_L g1657 ( 
.A(n_1643),
.Y(n_1657)
);

BUFx2_ASAP7_75t_L g1658 ( 
.A(n_1633),
.Y(n_1658)
);

INVx1_ASAP7_75t_L g1659 ( 
.A(n_1614),
.Y(n_1659)
);

BUFx2_ASAP7_75t_L g1660 ( 
.A(n_1649),
.Y(n_1660)
);

INVx1_ASAP7_75t_L g1661 ( 
.A(n_1614),
.Y(n_1661)
);

HB1xp67_ASAP7_75t_L g1662 ( 
.A(n_1630),
.Y(n_1662)
);

INVx1_ASAP7_75t_L g1663 ( 
.A(n_1630),
.Y(n_1663)
);

INVx1_ASAP7_75t_L g1664 ( 
.A(n_1634),
.Y(n_1664)
);

INVx1_ASAP7_75t_L g1665 ( 
.A(n_1634),
.Y(n_1665)
);

BUFx8_ASAP7_75t_L g1666 ( 
.A(n_1625),
.Y(n_1666)
);

BUFx2_ASAP7_75t_L g1667 ( 
.A(n_1649),
.Y(n_1667)
);

NAND2xp5_ASAP7_75t_L g1668 ( 
.A(n_1627),
.B(n_1608),
.Y(n_1668)
);

AND2x2_ASAP7_75t_L g1669 ( 
.A(n_1619),
.B(n_1593),
.Y(n_1669)
);

AND2x2_ASAP7_75t_L g1670 ( 
.A(n_1619),
.B(n_1594),
.Y(n_1670)
);

INVx4_ASAP7_75t_SL g1671 ( 
.A(n_1631),
.Y(n_1671)
);

OR2x6_ASAP7_75t_L g1672 ( 
.A(n_1637),
.B(n_1549),
.Y(n_1672)
);

BUFx8_ASAP7_75t_L g1673 ( 
.A(n_1631),
.Y(n_1673)
);

OR2x6_ASAP7_75t_L g1674 ( 
.A(n_1623),
.B(n_1549),
.Y(n_1674)
);

OA21x2_ASAP7_75t_L g1675 ( 
.A1(n_1615),
.A2(n_1545),
.B(n_1553),
.Y(n_1675)
);

NAND2xp5_ASAP7_75t_L g1676 ( 
.A(n_1650),
.B(n_1590),
.Y(n_1676)
);

BUFx3_ASAP7_75t_L g1677 ( 
.A(n_1643),
.Y(n_1677)
);

AND2x6_ASAP7_75t_L g1678 ( 
.A(n_1638),
.B(n_1611),
.Y(n_1678)
);

AOI21xp33_ASAP7_75t_L g1679 ( 
.A1(n_1613),
.A2(n_1575),
.B(n_1548),
.Y(n_1679)
);

BUFx2_ASAP7_75t_L g1680 ( 
.A(n_1643),
.Y(n_1680)
);

BUFx2_ASAP7_75t_L g1681 ( 
.A(n_1624),
.Y(n_1681)
);

AO21x2_ASAP7_75t_L g1682 ( 
.A1(n_1632),
.A2(n_1548),
.B(n_1575),
.Y(n_1682)
);

AND2x2_ASAP7_75t_L g1683 ( 
.A(n_1635),
.B(n_1594),
.Y(n_1683)
);

INVx2_ASAP7_75t_L g1684 ( 
.A(n_1628),
.Y(n_1684)
);

CKINVDCx5p33_ASAP7_75t_R g1685 ( 
.A(n_1618),
.Y(n_1685)
);

INVx1_ASAP7_75t_L g1686 ( 
.A(n_1642),
.Y(n_1686)
);

INVx2_ASAP7_75t_L g1687 ( 
.A(n_1641),
.Y(n_1687)
);

INVx1_ASAP7_75t_L g1688 ( 
.A(n_1662),
.Y(n_1688)
);

AND2x2_ASAP7_75t_L g1689 ( 
.A(n_1658),
.B(n_1646),
.Y(n_1689)
);

INVx2_ASAP7_75t_L g1690 ( 
.A(n_1682),
.Y(n_1690)
);

AND2x2_ASAP7_75t_L g1691 ( 
.A(n_1658),
.B(n_1648),
.Y(n_1691)
);

AND2x2_ASAP7_75t_L g1692 ( 
.A(n_1658),
.B(n_1590),
.Y(n_1692)
);

NOR2xp33_ASAP7_75t_L g1693 ( 
.A(n_1654),
.B(n_1490),
.Y(n_1693)
);

NAND5xp2_ASAP7_75t_SL g1694 ( 
.A(n_1685),
.B(n_1622),
.C(n_1652),
.D(n_1638),
.E(n_1645),
.Y(n_1694)
);

AND2x2_ASAP7_75t_L g1695 ( 
.A(n_1671),
.B(n_1592),
.Y(n_1695)
);

OR2x2_ASAP7_75t_L g1696 ( 
.A(n_1676),
.B(n_1620),
.Y(n_1696)
);

OR2x2_ASAP7_75t_L g1697 ( 
.A(n_1676),
.B(n_1620),
.Y(n_1697)
);

INVx1_ASAP7_75t_L g1698 ( 
.A(n_1662),
.Y(n_1698)
);

NAND2xp5_ASAP7_75t_L g1699 ( 
.A(n_1654),
.B(n_1652),
.Y(n_1699)
);

NAND3x1_ASAP7_75t_L g1700 ( 
.A(n_1657),
.B(n_1621),
.C(n_1602),
.Y(n_1700)
);

INVx2_ASAP7_75t_L g1701 ( 
.A(n_1682),
.Y(n_1701)
);

OR2x2_ASAP7_75t_L g1702 ( 
.A(n_1668),
.B(n_1639),
.Y(n_1702)
);

AND2x2_ASAP7_75t_L g1703 ( 
.A(n_1671),
.B(n_1592),
.Y(n_1703)
);

NAND3xp33_ASAP7_75t_L g1704 ( 
.A(n_1679),
.B(n_1617),
.C(n_1565),
.Y(n_1704)
);

NOR2xp33_ASAP7_75t_SL g1705 ( 
.A(n_1666),
.B(n_1490),
.Y(n_1705)
);

OR2x2_ASAP7_75t_L g1706 ( 
.A(n_1668),
.B(n_1639),
.Y(n_1706)
);

AND2x2_ASAP7_75t_L g1707 ( 
.A(n_1671),
.B(n_1592),
.Y(n_1707)
);

OR2x2_ASAP7_75t_L g1708 ( 
.A(n_1659),
.B(n_1629),
.Y(n_1708)
);

INVx1_ASAP7_75t_L g1709 ( 
.A(n_1659),
.Y(n_1709)
);

AND2x2_ASAP7_75t_L g1710 ( 
.A(n_1671),
.B(n_1597),
.Y(n_1710)
);

INVx6_ASAP7_75t_L g1711 ( 
.A(n_1666),
.Y(n_1711)
);

OR2x2_ASAP7_75t_L g1712 ( 
.A(n_1661),
.B(n_1629),
.Y(n_1712)
);

INVx1_ASAP7_75t_L g1713 ( 
.A(n_1661),
.Y(n_1713)
);

INVx1_ASAP7_75t_L g1714 ( 
.A(n_1663),
.Y(n_1714)
);

INVx1_ASAP7_75t_L g1715 ( 
.A(n_1663),
.Y(n_1715)
);

NAND2xp5_ASAP7_75t_L g1716 ( 
.A(n_1681),
.B(n_1597),
.Y(n_1716)
);

NAND2xp5_ASAP7_75t_L g1717 ( 
.A(n_1681),
.B(n_1597),
.Y(n_1717)
);

INVx1_ASAP7_75t_L g1718 ( 
.A(n_1664),
.Y(n_1718)
);

OAI33xp33_ASAP7_75t_L g1719 ( 
.A1(n_1664),
.A2(n_1647),
.A3(n_1642),
.B1(n_1644),
.B2(n_1606),
.B3(n_1636),
.Y(n_1719)
);

NAND2xp5_ASAP7_75t_L g1720 ( 
.A(n_1681),
.B(n_1601),
.Y(n_1720)
);

NOR2x1_ASAP7_75t_L g1721 ( 
.A(n_1660),
.B(n_1464),
.Y(n_1721)
);

HB1xp67_ASAP7_75t_L g1722 ( 
.A(n_1665),
.Y(n_1722)
);

NAND2xp5_ASAP7_75t_L g1723 ( 
.A(n_1675),
.B(n_1601),
.Y(n_1723)
);

AND2x2_ASAP7_75t_L g1724 ( 
.A(n_1671),
.B(n_1601),
.Y(n_1724)
);

INVx1_ASAP7_75t_SL g1725 ( 
.A(n_1671),
.Y(n_1725)
);

AND2x2_ASAP7_75t_L g1726 ( 
.A(n_1669),
.B(n_1594),
.Y(n_1726)
);

OR2x2_ASAP7_75t_L g1727 ( 
.A(n_1665),
.B(n_1644),
.Y(n_1727)
);

NAND2xp5_ASAP7_75t_SL g1728 ( 
.A(n_1673),
.B(n_1640),
.Y(n_1728)
);

INVx2_ASAP7_75t_L g1729 ( 
.A(n_1682),
.Y(n_1729)
);

AND2x2_ASAP7_75t_L g1730 ( 
.A(n_1669),
.B(n_1595),
.Y(n_1730)
);

INVx1_ASAP7_75t_L g1731 ( 
.A(n_1722),
.Y(n_1731)
);

OR2x2_ASAP7_75t_L g1732 ( 
.A(n_1696),
.B(n_1686),
.Y(n_1732)
);

NAND2xp5_ASAP7_75t_L g1733 ( 
.A(n_1691),
.B(n_1660),
.Y(n_1733)
);

INVx2_ASAP7_75t_L g1734 ( 
.A(n_1692),
.Y(n_1734)
);

INVx2_ASAP7_75t_L g1735 ( 
.A(n_1692),
.Y(n_1735)
);

INVx1_ASAP7_75t_L g1736 ( 
.A(n_1709),
.Y(n_1736)
);

AND2x2_ASAP7_75t_L g1737 ( 
.A(n_1691),
.B(n_1669),
.Y(n_1737)
);

AOI22xp5_ASAP7_75t_L g1738 ( 
.A1(n_1704),
.A2(n_1679),
.B1(n_1675),
.B2(n_1621),
.Y(n_1738)
);

OR2x2_ASAP7_75t_L g1739 ( 
.A(n_1696),
.B(n_1686),
.Y(n_1739)
);

INVx3_ASAP7_75t_R g1740 ( 
.A(n_1711),
.Y(n_1740)
);

HB1xp67_ASAP7_75t_L g1741 ( 
.A(n_1688),
.Y(n_1741)
);

NAND2xp5_ASAP7_75t_L g1742 ( 
.A(n_1699),
.B(n_1660),
.Y(n_1742)
);

INVx1_ASAP7_75t_L g1743 ( 
.A(n_1713),
.Y(n_1743)
);

NAND3xp33_ASAP7_75t_L g1744 ( 
.A(n_1698),
.B(n_1675),
.C(n_1673),
.Y(n_1744)
);

NAND2xp5_ASAP7_75t_L g1745 ( 
.A(n_1697),
.B(n_1667),
.Y(n_1745)
);

INVx1_ASAP7_75t_L g1746 ( 
.A(n_1714),
.Y(n_1746)
);

INVx1_ASAP7_75t_L g1747 ( 
.A(n_1715),
.Y(n_1747)
);

INVxp67_ASAP7_75t_SL g1748 ( 
.A(n_1700),
.Y(n_1748)
);

HB1xp67_ASAP7_75t_L g1749 ( 
.A(n_1718),
.Y(n_1749)
);

NOR2xp33_ASAP7_75t_L g1750 ( 
.A(n_1711),
.B(n_1666),
.Y(n_1750)
);

INVx1_ASAP7_75t_SL g1751 ( 
.A(n_1711),
.Y(n_1751)
);

NOR2x1_ASAP7_75t_L g1752 ( 
.A(n_1721),
.B(n_1667),
.Y(n_1752)
);

INVx1_ASAP7_75t_L g1753 ( 
.A(n_1708),
.Y(n_1753)
);

INVx1_ASAP7_75t_L g1754 ( 
.A(n_1708),
.Y(n_1754)
);

INVx1_ASAP7_75t_L g1755 ( 
.A(n_1712),
.Y(n_1755)
);

HB1xp67_ASAP7_75t_L g1756 ( 
.A(n_1702),
.Y(n_1756)
);

INVx1_ASAP7_75t_L g1757 ( 
.A(n_1712),
.Y(n_1757)
);

NAND2xp5_ASAP7_75t_L g1758 ( 
.A(n_1697),
.B(n_1667),
.Y(n_1758)
);

AND2x2_ASAP7_75t_L g1759 ( 
.A(n_1695),
.B(n_1670),
.Y(n_1759)
);

NOR3xp33_ASAP7_75t_L g1760 ( 
.A(n_1725),
.B(n_1616),
.C(n_1657),
.Y(n_1760)
);

OR2x2_ASAP7_75t_L g1761 ( 
.A(n_1702),
.B(n_1675),
.Y(n_1761)
);

AND2x2_ASAP7_75t_L g1762 ( 
.A(n_1695),
.B(n_1670),
.Y(n_1762)
);

INVx1_ASAP7_75t_L g1763 ( 
.A(n_1727),
.Y(n_1763)
);

INVx1_ASAP7_75t_L g1764 ( 
.A(n_1727),
.Y(n_1764)
);

NAND2xp5_ASAP7_75t_L g1765 ( 
.A(n_1706),
.B(n_1675),
.Y(n_1765)
);

INVx2_ASAP7_75t_L g1766 ( 
.A(n_1690),
.Y(n_1766)
);

NAND2xp5_ASAP7_75t_L g1767 ( 
.A(n_1756),
.B(n_1763),
.Y(n_1767)
);

INVx1_ASAP7_75t_SL g1768 ( 
.A(n_1751),
.Y(n_1768)
);

OR2x2_ASAP7_75t_L g1769 ( 
.A(n_1732),
.B(n_1716),
.Y(n_1769)
);

INVx2_ASAP7_75t_L g1770 ( 
.A(n_1761),
.Y(n_1770)
);

NOR3xp33_ASAP7_75t_L g1771 ( 
.A(n_1748),
.B(n_1689),
.C(n_1719),
.Y(n_1771)
);

AND2x2_ASAP7_75t_L g1772 ( 
.A(n_1737),
.B(n_1703),
.Y(n_1772)
);

AND2x2_ASAP7_75t_L g1773 ( 
.A(n_1737),
.B(n_1734),
.Y(n_1773)
);

INVx1_ASAP7_75t_SL g1774 ( 
.A(n_1733),
.Y(n_1774)
);

INVx2_ASAP7_75t_L g1775 ( 
.A(n_1761),
.Y(n_1775)
);

INVx2_ASAP7_75t_L g1776 ( 
.A(n_1734),
.Y(n_1776)
);

OR2x2_ASAP7_75t_L g1777 ( 
.A(n_1732),
.B(n_1717),
.Y(n_1777)
);

INVx1_ASAP7_75t_SL g1778 ( 
.A(n_1741),
.Y(n_1778)
);

AND2x2_ASAP7_75t_L g1779 ( 
.A(n_1735),
.B(n_1703),
.Y(n_1779)
);

INVx1_ASAP7_75t_L g1780 ( 
.A(n_1749),
.Y(n_1780)
);

AOI222xp33_ASAP7_75t_L g1781 ( 
.A1(n_1765),
.A2(n_1723),
.B1(n_1689),
.B2(n_1694),
.C1(n_1653),
.C2(n_1655),
.Y(n_1781)
);

AOI22xp33_ASAP7_75t_L g1782 ( 
.A1(n_1738),
.A2(n_1672),
.B1(n_1674),
.B2(n_1678),
.Y(n_1782)
);

AND2x2_ASAP7_75t_L g1783 ( 
.A(n_1735),
.B(n_1707),
.Y(n_1783)
);

BUFx3_ASAP7_75t_L g1784 ( 
.A(n_1750),
.Y(n_1784)
);

INVx1_ASAP7_75t_L g1785 ( 
.A(n_1736),
.Y(n_1785)
);

INVx1_ASAP7_75t_L g1786 ( 
.A(n_1736),
.Y(n_1786)
);

OR2x2_ASAP7_75t_L g1787 ( 
.A(n_1739),
.B(n_1720),
.Y(n_1787)
);

NAND2xp5_ASAP7_75t_L g1788 ( 
.A(n_1763),
.B(n_1666),
.Y(n_1788)
);

INVx1_ASAP7_75t_L g1789 ( 
.A(n_1739),
.Y(n_1789)
);

NAND2xp5_ASAP7_75t_L g1790 ( 
.A(n_1764),
.B(n_1666),
.Y(n_1790)
);

NAND2xp5_ASAP7_75t_L g1791 ( 
.A(n_1764),
.B(n_1726),
.Y(n_1791)
);

NOR2x1p5_ASAP7_75t_L g1792 ( 
.A(n_1745),
.B(n_1758),
.Y(n_1792)
);

OR2x2_ASAP7_75t_L g1793 ( 
.A(n_1768),
.B(n_1742),
.Y(n_1793)
);

NAND2xp5_ASAP7_75t_L g1794 ( 
.A(n_1768),
.B(n_1753),
.Y(n_1794)
);

AOI22xp33_ASAP7_75t_L g1795 ( 
.A1(n_1781),
.A2(n_1744),
.B1(n_1760),
.B2(n_1672),
.Y(n_1795)
);

NOR2xp67_ASAP7_75t_SL g1796 ( 
.A(n_1784),
.B(n_1457),
.Y(n_1796)
);

INVx1_ASAP7_75t_L g1797 ( 
.A(n_1773),
.Y(n_1797)
);

OAI21xp5_ASAP7_75t_L g1798 ( 
.A1(n_1771),
.A2(n_1700),
.B(n_1752),
.Y(n_1798)
);

INVxp67_ASAP7_75t_L g1799 ( 
.A(n_1784),
.Y(n_1799)
);

INVx2_ASAP7_75t_L g1800 ( 
.A(n_1772),
.Y(n_1800)
);

NAND2xp5_ASAP7_75t_L g1801 ( 
.A(n_1773),
.B(n_1754),
.Y(n_1801)
);

AOI22xp5_ASAP7_75t_L g1802 ( 
.A1(n_1792),
.A2(n_1678),
.B1(n_1731),
.B2(n_1672),
.Y(n_1802)
);

OA21x2_ASAP7_75t_L g1803 ( 
.A1(n_1780),
.A2(n_1731),
.B(n_1766),
.Y(n_1803)
);

AOI21xp5_ASAP7_75t_L g1804 ( 
.A1(n_1778),
.A2(n_1728),
.B(n_1705),
.Y(n_1804)
);

INVx1_ASAP7_75t_L g1805 ( 
.A(n_1785),
.Y(n_1805)
);

OAI221xp5_ASAP7_75t_L g1806 ( 
.A1(n_1782),
.A2(n_1672),
.B1(n_1755),
.B2(n_1757),
.C(n_1655),
.Y(n_1806)
);

INVx1_ASAP7_75t_L g1807 ( 
.A(n_1785),
.Y(n_1807)
);

OR2x2_ASAP7_75t_L g1808 ( 
.A(n_1791),
.B(n_1743),
.Y(n_1808)
);

NAND3xp33_ASAP7_75t_SL g1809 ( 
.A(n_1778),
.B(n_1728),
.C(n_1759),
.Y(n_1809)
);

NOR3xp33_ASAP7_75t_L g1810 ( 
.A(n_1774),
.B(n_1747),
.C(n_1746),
.Y(n_1810)
);

AOI31xp33_ASAP7_75t_SL g1811 ( 
.A1(n_1788),
.A2(n_1740),
.A3(n_1693),
.B(n_1673),
.Y(n_1811)
);

OAI22xp33_ASAP7_75t_L g1812 ( 
.A1(n_1770),
.A2(n_1672),
.B1(n_1674),
.B2(n_1653),
.Y(n_1812)
);

AOI22xp33_ASAP7_75t_L g1813 ( 
.A1(n_1795),
.A2(n_1770),
.B1(n_1775),
.B2(n_1792),
.Y(n_1813)
);

AOI22xp5_ASAP7_75t_L g1814 ( 
.A1(n_1798),
.A2(n_1775),
.B1(n_1772),
.B2(n_1776),
.Y(n_1814)
);

AND2x2_ASAP7_75t_L g1815 ( 
.A(n_1799),
.B(n_1800),
.Y(n_1815)
);

AOI21xp5_ASAP7_75t_L g1816 ( 
.A1(n_1809),
.A2(n_1767),
.B(n_1780),
.Y(n_1816)
);

HB1xp67_ASAP7_75t_L g1817 ( 
.A(n_1803),
.Y(n_1817)
);

NAND2xp5_ASAP7_75t_L g1818 ( 
.A(n_1797),
.B(n_1810),
.Y(n_1818)
);

NAND2xp5_ASAP7_75t_L g1819 ( 
.A(n_1803),
.B(n_1789),
.Y(n_1819)
);

INVx1_ASAP7_75t_L g1820 ( 
.A(n_1794),
.Y(n_1820)
);

INVx2_ASAP7_75t_L g1821 ( 
.A(n_1793),
.Y(n_1821)
);

AND2x2_ASAP7_75t_L g1822 ( 
.A(n_1796),
.B(n_1784),
.Y(n_1822)
);

NAND2xp5_ASAP7_75t_L g1823 ( 
.A(n_1801),
.B(n_1789),
.Y(n_1823)
);

NAND2xp5_ASAP7_75t_L g1824 ( 
.A(n_1808),
.B(n_1776),
.Y(n_1824)
);

AOI221xp5_ASAP7_75t_L g1825 ( 
.A1(n_1817),
.A2(n_1806),
.B1(n_1807),
.B2(n_1805),
.C(n_1786),
.Y(n_1825)
);

AOI21xp5_ASAP7_75t_L g1826 ( 
.A1(n_1816),
.A2(n_1804),
.B(n_1790),
.Y(n_1826)
);

INVx1_ASAP7_75t_L g1827 ( 
.A(n_1824),
.Y(n_1827)
);

OAI211xp5_ASAP7_75t_L g1828 ( 
.A1(n_1814),
.A2(n_1786),
.B(n_1802),
.C(n_1779),
.Y(n_1828)
);

AOI22xp33_ASAP7_75t_SL g1829 ( 
.A1(n_1819),
.A2(n_1779),
.B1(n_1783),
.B2(n_1672),
.Y(n_1829)
);

AND2x2_ASAP7_75t_L g1830 ( 
.A(n_1822),
.B(n_1783),
.Y(n_1830)
);

AOI221xp5_ASAP7_75t_L g1831 ( 
.A1(n_1819),
.A2(n_1812),
.B1(n_1802),
.B2(n_1684),
.C(n_1690),
.Y(n_1831)
);

AOI21xp5_ASAP7_75t_L g1832 ( 
.A1(n_1818),
.A2(n_1777),
.B(n_1769),
.Y(n_1832)
);

AOI221x1_ASAP7_75t_L g1833 ( 
.A1(n_1820),
.A2(n_1740),
.B1(n_1811),
.B2(n_1766),
.C(n_1759),
.Y(n_1833)
);

INVx2_ASAP7_75t_SL g1834 ( 
.A(n_1815),
.Y(n_1834)
);

AOI21xp5_ASAP7_75t_L g1835 ( 
.A1(n_1823),
.A2(n_1777),
.B(n_1769),
.Y(n_1835)
);

OAI22xp5_ASAP7_75t_L g1836 ( 
.A1(n_1821),
.A2(n_1787),
.B1(n_1724),
.B2(n_1710),
.Y(n_1836)
);

OAI211xp5_ASAP7_75t_SL g1837 ( 
.A1(n_1826),
.A2(n_1813),
.B(n_1787),
.C(n_1729),
.Y(n_1837)
);

INVx2_ASAP7_75t_SL g1838 ( 
.A(n_1830),
.Y(n_1838)
);

OAI21xp5_ASAP7_75t_L g1839 ( 
.A1(n_1832),
.A2(n_1762),
.B(n_1710),
.Y(n_1839)
);

XOR2xp5_ASAP7_75t_L g1840 ( 
.A(n_1834),
.B(n_1522),
.Y(n_1840)
);

AOI221x1_ASAP7_75t_L g1841 ( 
.A1(n_1827),
.A2(n_1762),
.B1(n_1657),
.B2(n_1653),
.C(n_1655),
.Y(n_1841)
);

OR2x2_ASAP7_75t_L g1842 ( 
.A(n_1838),
.B(n_1835),
.Y(n_1842)
);

NAND3xp33_ASAP7_75t_L g1843 ( 
.A(n_1837),
.B(n_1833),
.C(n_1825),
.Y(n_1843)
);

AND2x4_ASAP7_75t_L g1844 ( 
.A(n_1839),
.B(n_1707),
.Y(n_1844)
);

NAND3xp33_ASAP7_75t_L g1845 ( 
.A(n_1841),
.B(n_1828),
.C(n_1829),
.Y(n_1845)
);

AOI221xp5_ASAP7_75t_L g1846 ( 
.A1(n_1840),
.A2(n_1831),
.B1(n_1836),
.B2(n_1701),
.C(n_1729),
.Y(n_1846)
);

INVx2_ASAP7_75t_SL g1847 ( 
.A(n_1838),
.Y(n_1847)
);

AOI22xp5_ASAP7_75t_L g1848 ( 
.A1(n_1843),
.A2(n_1724),
.B1(n_1673),
.B2(n_1684),
.Y(n_1848)
);

NOR2xp33_ASAP7_75t_R g1849 ( 
.A(n_1842),
.B(n_1673),
.Y(n_1849)
);

INVx1_ASAP7_75t_L g1850 ( 
.A(n_1847),
.Y(n_1850)
);

INVx1_ASAP7_75t_L g1851 ( 
.A(n_1845),
.Y(n_1851)
);

NAND2xp5_ASAP7_75t_L g1852 ( 
.A(n_1844),
.B(n_1680),
.Y(n_1852)
);

OR2x6_ASAP7_75t_L g1853 ( 
.A(n_1850),
.B(n_1674),
.Y(n_1853)
);

INVx1_ASAP7_75t_L g1854 ( 
.A(n_1851),
.Y(n_1854)
);

AOI221xp5_ASAP7_75t_L g1855 ( 
.A1(n_1848),
.A2(n_1846),
.B1(n_1701),
.B2(n_1684),
.C(n_1656),
.Y(n_1855)
);

NAND2xp5_ASAP7_75t_L g1856 ( 
.A(n_1854),
.B(n_1852),
.Y(n_1856)
);

OAI322xp33_ASAP7_75t_L g1857 ( 
.A1(n_1856),
.A2(n_1849),
.A3(n_1855),
.B1(n_1853),
.B2(n_1656),
.C1(n_1657),
.C2(n_1680),
.Y(n_1857)
);

INVx3_ASAP7_75t_L g1858 ( 
.A(n_1857),
.Y(n_1858)
);

INVx1_ASAP7_75t_L g1859 ( 
.A(n_1857),
.Y(n_1859)
);

INVx1_ASAP7_75t_L g1860 ( 
.A(n_1858),
.Y(n_1860)
);

AO22x2_ASAP7_75t_L g1861 ( 
.A1(n_1858),
.A2(n_1656),
.B1(n_1726),
.B2(n_1730),
.Y(n_1861)
);

INVx2_ASAP7_75t_SL g1862 ( 
.A(n_1861),
.Y(n_1862)
);

OA21x2_ASAP7_75t_L g1863 ( 
.A1(n_1860),
.A2(n_1859),
.B(n_1858),
.Y(n_1863)
);

NAND5xp2_ASAP7_75t_SL g1864 ( 
.A(n_1863),
.B(n_1730),
.C(n_1683),
.D(n_1670),
.E(n_1680),
.Y(n_1864)
);

A2O1A1O1Ixp25_ASAP7_75t_L g1865 ( 
.A1(n_1864),
.A2(n_1862),
.B(n_1678),
.C(n_1672),
.D(n_1677),
.Y(n_1865)
);

AOI22xp33_ASAP7_75t_R g1866 ( 
.A1(n_1865),
.A2(n_1651),
.B1(n_1687),
.B2(n_1677),
.Y(n_1866)
);

HB1xp67_ASAP7_75t_L g1867 ( 
.A(n_1866),
.Y(n_1867)
);

AOI22xp5_ASAP7_75t_L g1868 ( 
.A1(n_1867),
.A2(n_1677),
.B1(n_1657),
.B2(n_1678),
.Y(n_1868)
);

AOI211xp5_ASAP7_75t_L g1869 ( 
.A1(n_1868),
.A2(n_1677),
.B(n_1683),
.C(n_1580),
.Y(n_1869)
);


endmodule