module fake_jpeg_23154_n_231 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_231);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_231;

wire n_159;
wire n_117;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_84;
wire n_59;
wire n_98;
wire n_178;
wire n_228;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_16;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_223;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_24;
wire n_44;
wire n_143;
wire n_202;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_131;
wire n_56;
wire n_212;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_216;
wire n_217;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

BUFx6f_ASAP7_75t_L g16 ( 
.A(n_7),
.Y(n_16)
);

INVx13_ASAP7_75t_L g17 ( 
.A(n_10),
.Y(n_17)
);

BUFx12f_ASAP7_75t_L g18 ( 
.A(n_2),
.Y(n_18)
);

BUFx12f_ASAP7_75t_L g19 ( 
.A(n_11),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_8),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_10),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_5),
.Y(n_22)
);

BUFx12f_ASAP7_75t_L g23 ( 
.A(n_10),
.Y(n_23)
);

BUFx12f_ASAP7_75t_L g24 ( 
.A(n_7),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_5),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_9),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_5),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_14),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_11),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_0),
.Y(n_30)
);

INVx6_ASAP7_75t_L g31 ( 
.A(n_0),
.Y(n_31)
);

INVx2_ASAP7_75t_L g32 ( 
.A(n_8),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_15),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_18),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_L g45 ( 
.A(n_34),
.B(n_35),
.Y(n_45)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_18),
.Y(n_35)
);

INVx2_ASAP7_75t_SL g36 ( 
.A(n_18),
.Y(n_36)
);

INVx4_ASAP7_75t_SL g52 ( 
.A(n_36),
.Y(n_52)
);

INVx2_ASAP7_75t_L g37 ( 
.A(n_19),
.Y(n_37)
);

INVx6_ASAP7_75t_L g43 ( 
.A(n_37),
.Y(n_43)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_25),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_38),
.B(n_39),
.Y(n_58)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_19),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_19),
.Y(n_40)
);

INVx3_ASAP7_75t_L g47 ( 
.A(n_40),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g41 ( 
.A(n_17),
.B(n_0),
.Y(n_41)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_41),
.Y(n_44)
);

INVx3_ASAP7_75t_L g42 ( 
.A(n_19),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_42),
.B(n_23),
.Y(n_59)
);

INVx2_ASAP7_75t_L g46 ( 
.A(n_40),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_46),
.B(n_49),
.Y(n_62)
);

OAI22xp33_ASAP7_75t_SL g48 ( 
.A1(n_38),
.A2(n_32),
.B1(n_31),
.B2(n_17),
.Y(n_48)
);

AOI22xp33_ASAP7_75t_L g61 ( 
.A1(n_48),
.A2(n_23),
.B1(n_24),
.B2(n_22),
.Y(n_61)
);

INVx3_ASAP7_75t_L g49 ( 
.A(n_40),
.Y(n_49)
);

INVx2_ASAP7_75t_L g50 ( 
.A(n_40),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_50),
.B(n_56),
.Y(n_74)
);

AND2x2_ASAP7_75t_L g51 ( 
.A(n_42),
.B(n_24),
.Y(n_51)
);

A2O1A1Ixp33_ASAP7_75t_L g64 ( 
.A1(n_51),
.A2(n_24),
.B(n_16),
.C(n_21),
.Y(n_64)
);

AOI21xp5_ASAP7_75t_L g53 ( 
.A1(n_37),
.A2(n_32),
.B(n_18),
.Y(n_53)
);

AOI21xp5_ASAP7_75t_L g60 ( 
.A1(n_53),
.A2(n_24),
.B(n_23),
.Y(n_60)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_41),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_SL g75 ( 
.A(n_54),
.B(n_55),
.Y(n_75)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_37),
.Y(n_55)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_42),
.Y(n_56)
);

AOI22xp33_ASAP7_75t_L g57 ( 
.A1(n_39),
.A2(n_31),
.B1(n_30),
.B2(n_25),
.Y(n_57)
);

OAI22xp5_ASAP7_75t_L g81 ( 
.A1(n_57),
.A2(n_20),
.B1(n_26),
.B2(n_27),
.Y(n_81)
);

CKINVDCx16_ASAP7_75t_R g76 ( 
.A(n_59),
.Y(n_76)
);

OAI22xp5_ASAP7_75t_L g112 ( 
.A1(n_60),
.A2(n_61),
.B1(n_64),
.B2(n_80),
.Y(n_112)
);

OAI22xp5_ASAP7_75t_SL g63 ( 
.A1(n_53),
.A2(n_35),
.B1(n_34),
.B2(n_23),
.Y(n_63)
);

AOI22xp5_ASAP7_75t_L g96 ( 
.A1(n_63),
.A2(n_81),
.B1(n_82),
.B2(n_75),
.Y(n_96)
);

BUFx12_ASAP7_75t_L g65 ( 
.A(n_52),
.Y(n_65)
);

CKINVDCx16_ASAP7_75t_R g95 ( 
.A(n_65),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g66 ( 
.A(n_44),
.B(n_35),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_L g100 ( 
.A(n_66),
.B(n_69),
.Y(n_100)
);

CKINVDCx20_ASAP7_75t_R g67 ( 
.A(n_58),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_67),
.B(n_68),
.Y(n_90)
);

INVx2_ASAP7_75t_L g68 ( 
.A(n_46),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_L g69 ( 
.A(n_44),
.B(n_34),
.Y(n_69)
);

AOI22xp5_ASAP7_75t_L g70 ( 
.A1(n_43),
.A2(n_54),
.B1(n_36),
.B2(n_55),
.Y(n_70)
);

OAI22xp5_ASAP7_75t_SL g104 ( 
.A1(n_70),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_104)
);

INVx4_ASAP7_75t_L g71 ( 
.A(n_47),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_71),
.B(n_72),
.Y(n_92)
);

INVx8_ASAP7_75t_L g72 ( 
.A(n_47),
.Y(n_72)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_45),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_73),
.B(n_78),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_SL g77 ( 
.A(n_56),
.B(n_33),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_SL g98 ( 
.A(n_77),
.B(n_67),
.Y(n_98)
);

INVxp33_ASAP7_75t_L g78 ( 
.A(n_49),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_43),
.B(n_33),
.Y(n_79)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_79),
.Y(n_103)
);

AOI22xp33_ASAP7_75t_L g80 ( 
.A1(n_51),
.A2(n_30),
.B1(n_26),
.B2(n_22),
.Y(n_80)
);

O2A1O1Ixp33_ASAP7_75t_L g82 ( 
.A1(n_51),
.A2(n_36),
.B(n_21),
.C(n_16),
.Y(n_82)
);

AND2x2_ASAP7_75t_SL g83 ( 
.A(n_52),
.B(n_36),
.Y(n_83)
);

AOI21xp33_ASAP7_75t_L g93 ( 
.A1(n_83),
.A2(n_69),
.B(n_66),
.Y(n_93)
);

BUFx6f_ASAP7_75t_L g84 ( 
.A(n_50),
.Y(n_84)
);

BUFx6f_ASAP7_75t_L g89 ( 
.A(n_84),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_SL g85 ( 
.A(n_52),
.B(n_20),
.Y(n_85)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_85),
.Y(n_105)
);

INVx2_ASAP7_75t_L g86 ( 
.A(n_46),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_86),
.B(n_1),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_58),
.B(n_27),
.Y(n_87)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_87),
.Y(n_108)
);

AOI22xp5_ASAP7_75t_SL g88 ( 
.A1(n_44),
.A2(n_29),
.B1(n_28),
.B2(n_3),
.Y(n_88)
);

INVxp67_ASAP7_75t_L g91 ( 
.A(n_88),
.Y(n_91)
);

A2O1A1Ixp33_ASAP7_75t_L g130 ( 
.A1(n_93),
.A2(n_65),
.B(n_6),
.C(n_7),
.Y(n_130)
);

NOR2x1_ASAP7_75t_L g94 ( 
.A(n_83),
.B(n_1),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_SL g135 ( 
.A(n_94),
.B(n_4),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_L g132 ( 
.A(n_96),
.B(n_97),
.Y(n_132)
);

INVx3_ASAP7_75t_L g97 ( 
.A(n_84),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g120 ( 
.A(n_98),
.B(n_111),
.Y(n_120)
);

OAI22xp33_ASAP7_75t_L g99 ( 
.A1(n_60),
.A2(n_29),
.B1(n_28),
.B2(n_3),
.Y(n_99)
);

AOI22xp5_ASAP7_75t_L g119 ( 
.A1(n_99),
.A2(n_104),
.B1(n_106),
.B2(n_109),
.Y(n_119)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_102),
.Y(n_115)
);

OAI22xp5_ASAP7_75t_SL g106 ( 
.A1(n_64),
.A2(n_15),
.B1(n_14),
.B2(n_13),
.Y(n_106)
);

CKINVDCx20_ASAP7_75t_R g107 ( 
.A(n_74),
.Y(n_107)
);

CKINVDCx20_ASAP7_75t_R g126 ( 
.A(n_107),
.Y(n_126)
);

OAI22xp5_ASAP7_75t_SL g109 ( 
.A1(n_70),
.A2(n_13),
.B1(n_12),
.B2(n_6),
.Y(n_109)
);

BUFx6f_ASAP7_75t_L g110 ( 
.A(n_84),
.Y(n_110)
);

INVx13_ASAP7_75t_L g134 ( 
.A(n_110),
.Y(n_134)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_62),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_L g113 ( 
.A(n_73),
.B(n_12),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_L g122 ( 
.A(n_113),
.B(n_2),
.Y(n_122)
);

AOI21xp5_ASAP7_75t_L g114 ( 
.A1(n_91),
.A2(n_63),
.B(n_75),
.Y(n_114)
);

OAI21xp5_ASAP7_75t_SL g155 ( 
.A1(n_114),
.A2(n_116),
.B(n_117),
.Y(n_155)
);

OAI21xp5_ASAP7_75t_L g116 ( 
.A1(n_100),
.A2(n_85),
.B(n_83),
.Y(n_116)
);

AOI21xp5_ASAP7_75t_L g117 ( 
.A1(n_91),
.A2(n_76),
.B(n_71),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_L g118 ( 
.A(n_100),
.B(n_76),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_L g153 ( 
.A(n_118),
.B(n_121),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_L g121 ( 
.A(n_105),
.B(n_77),
.Y(n_121)
);

CKINVDCx14_ASAP7_75t_R g151 ( 
.A(n_122),
.Y(n_151)
);

OAI21xp5_ASAP7_75t_L g123 ( 
.A1(n_94),
.A2(n_82),
.B(n_88),
.Y(n_123)
);

XNOR2xp5_ASAP7_75t_L g138 ( 
.A(n_123),
.B(n_96),
.Y(n_138)
);

AND2x2_ASAP7_75t_L g124 ( 
.A(n_106),
.B(n_4),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_L g154 ( 
.A(n_124),
.B(n_131),
.Y(n_154)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_90),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_SL g143 ( 
.A(n_125),
.B(n_135),
.Y(n_143)
);

CKINVDCx20_ASAP7_75t_R g127 ( 
.A(n_92),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_L g140 ( 
.A(n_127),
.B(n_129),
.Y(n_140)
);

AOI22xp5_ASAP7_75t_L g128 ( 
.A1(n_112),
.A2(n_81),
.B1(n_72),
.B2(n_86),
.Y(n_128)
);

OAI22xp5_ASAP7_75t_L g152 ( 
.A1(n_128),
.A2(n_68),
.B1(n_97),
.B2(n_103),
.Y(n_152)
);

CKINVDCx20_ASAP7_75t_R g129 ( 
.A(n_98),
.Y(n_129)
);

AOI221xp5_ASAP7_75t_L g149 ( 
.A1(n_130),
.A2(n_108),
.B1(n_103),
.B2(n_8),
.C(n_9),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_L g131 ( 
.A(n_105),
.B(n_65),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g133 ( 
.A(n_107),
.B(n_65),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_L g157 ( 
.A(n_133),
.B(n_116),
.Y(n_157)
);

CKINVDCx20_ASAP7_75t_R g136 ( 
.A(n_101),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_L g145 ( 
.A(n_136),
.B(n_137),
.Y(n_145)
);

CKINVDCx20_ASAP7_75t_R g137 ( 
.A(n_109),
.Y(n_137)
);

XOR2xp5_ASAP7_75t_L g165 ( 
.A(n_138),
.B(n_119),
.Y(n_165)
);

MAJIxp5_ASAP7_75t_L g139 ( 
.A(n_118),
.B(n_95),
.C(n_111),
.Y(n_139)
);

MAJIxp5_ASAP7_75t_L g174 ( 
.A(n_139),
.B(n_115),
.C(n_130),
.Y(n_174)
);

OA21x2_ASAP7_75t_L g141 ( 
.A1(n_137),
.A2(n_99),
.B(n_104),
.Y(n_141)
);

OAI21xp5_ASAP7_75t_SL g178 ( 
.A1(n_141),
.A2(n_149),
.B(n_135),
.Y(n_178)
);

INVx4_ASAP7_75t_L g142 ( 
.A(n_134),
.Y(n_142)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_142),
.Y(n_162)
);

CKINVDCx16_ASAP7_75t_R g144 ( 
.A(n_120),
.Y(n_144)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_144),
.Y(n_163)
);

AO22x2_ASAP7_75t_L g146 ( 
.A1(n_114),
.A2(n_132),
.B1(n_117),
.B2(n_123),
.Y(n_146)
);

AOI22xp5_ASAP7_75t_L g169 ( 
.A1(n_146),
.A2(n_152),
.B1(n_157),
.B2(n_154),
.Y(n_169)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_120),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_L g167 ( 
.A(n_147),
.B(n_148),
.Y(n_167)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_133),
.Y(n_148)
);

NOR2xp33_ASAP7_75t_L g150 ( 
.A(n_126),
.B(n_108),
.Y(n_150)
);

CKINVDCx16_ASAP7_75t_R g166 ( 
.A(n_150),
.Y(n_166)
);

INVx2_ASAP7_75t_L g156 ( 
.A(n_134),
.Y(n_156)
);

INVx6_ASAP7_75t_L g175 ( 
.A(n_156),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_L g170 ( 
.A(n_157),
.B(n_158),
.Y(n_170)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_131),
.Y(n_158)
);

NOR2xp33_ASAP7_75t_L g159 ( 
.A(n_126),
.B(n_4),
.Y(n_159)
);

CKINVDCx20_ASAP7_75t_R g161 ( 
.A(n_159),
.Y(n_161)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_121),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_L g171 ( 
.A(n_160),
.B(n_125),
.Y(n_171)
);

OAI22xp5_ASAP7_75t_L g164 ( 
.A1(n_145),
.A2(n_128),
.B1(n_119),
.B2(n_129),
.Y(n_164)
);

AOI22xp5_ASAP7_75t_L g185 ( 
.A1(n_164),
.A2(n_146),
.B1(n_160),
.B2(n_154),
.Y(n_185)
);

XNOR2xp5_ASAP7_75t_L g186 ( 
.A(n_165),
.B(n_138),
.Y(n_186)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_140),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_L g180 ( 
.A(n_168),
.B(n_172),
.Y(n_180)
);

OAI22xp5_ASAP7_75t_L g191 ( 
.A1(n_169),
.A2(n_178),
.B1(n_179),
.B2(n_141),
.Y(n_191)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_171),
.Y(n_181)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_153),
.Y(n_172)
);

OA21x2_ASAP7_75t_L g173 ( 
.A1(n_146),
.A2(n_136),
.B(n_127),
.Y(n_173)
);

OAI21xp5_ASAP7_75t_L g190 ( 
.A1(n_173),
.A2(n_141),
.B(n_151),
.Y(n_190)
);

MAJIxp5_ASAP7_75t_L g183 ( 
.A(n_174),
.B(n_176),
.C(n_155),
.Y(n_183)
);

MAJIxp5_ASAP7_75t_L g176 ( 
.A(n_155),
.B(n_139),
.C(n_158),
.Y(n_176)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_153),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_L g187 ( 
.A(n_177),
.B(n_148),
.Y(n_187)
);

AOI22xp5_ASAP7_75t_L g179 ( 
.A1(n_146),
.A2(n_124),
.B1(n_115),
.B2(n_134),
.Y(n_179)
);

BUFx12_ASAP7_75t_L g182 ( 
.A(n_162),
.Y(n_182)
);

CKINVDCx20_ASAP7_75t_R g204 ( 
.A(n_182),
.Y(n_204)
);

MAJIxp5_ASAP7_75t_L g196 ( 
.A(n_183),
.B(n_186),
.C(n_189),
.Y(n_196)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_167),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_SL g201 ( 
.A(n_184),
.B(n_187),
.Y(n_201)
);

OAI22xp5_ASAP7_75t_L g202 ( 
.A1(n_185),
.A2(n_170),
.B1(n_181),
.B2(n_172),
.Y(n_202)
);

NAND2xp5_ASAP7_75t_L g188 ( 
.A(n_167),
.B(n_147),
.Y(n_188)
);

OAI21xp5_ASAP7_75t_L g197 ( 
.A1(n_188),
.A2(n_192),
.B(n_171),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_SL g189 ( 
.A(n_168),
.B(n_143),
.Y(n_189)
);

AOI21xp5_ASAP7_75t_SL g198 ( 
.A1(n_190),
.A2(n_178),
.B(n_173),
.Y(n_198)
);

AOI22xp5_ASAP7_75t_L g195 ( 
.A1(n_191),
.A2(n_193),
.B1(n_170),
.B2(n_177),
.Y(n_195)
);

MAJIxp5_ASAP7_75t_L g192 ( 
.A(n_176),
.B(n_156),
.C(n_122),
.Y(n_192)
);

OAI22xp5_ASAP7_75t_L g193 ( 
.A1(n_169),
.A2(n_124),
.B1(n_142),
.B2(n_89),
.Y(n_193)
);

OR2x2_ASAP7_75t_L g194 ( 
.A(n_188),
.B(n_161),
.Y(n_194)
);

NOR2xp33_ASAP7_75t_L g208 ( 
.A(n_194),
.B(n_195),
.Y(n_208)
);

OAI21xp5_ASAP7_75t_L g213 ( 
.A1(n_197),
.A2(n_179),
.B(n_163),
.Y(n_213)
);

AOI21xp5_ASAP7_75t_L g210 ( 
.A1(n_198),
.A2(n_200),
.B(n_174),
.Y(n_210)
);

HB1xp67_ASAP7_75t_L g199 ( 
.A(n_182),
.Y(n_199)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_199),
.Y(n_206)
);

AND2x2_ASAP7_75t_L g200 ( 
.A(n_180),
.B(n_165),
.Y(n_200)
);

AOI22xp5_ASAP7_75t_L g211 ( 
.A1(n_202),
.A2(n_203),
.B1(n_163),
.B2(n_162),
.Y(n_211)
);

HB1xp67_ASAP7_75t_L g203 ( 
.A(n_182),
.Y(n_203)
);

MAJIxp5_ASAP7_75t_L g205 ( 
.A(n_196),
.B(n_183),
.C(n_192),
.Y(n_205)
);

NAND2xp5_ASAP7_75t_L g218 ( 
.A(n_205),
.B(n_207),
.Y(n_218)
);

MAJIxp5_ASAP7_75t_L g207 ( 
.A(n_204),
.B(n_180),
.C(n_187),
.Y(n_207)
);

AO22x1_ASAP7_75t_L g209 ( 
.A1(n_201),
.A2(n_190),
.B1(n_173),
.B2(n_185),
.Y(n_209)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_209),
.Y(n_217)
);

NAND4xp25_ASAP7_75t_L g214 ( 
.A(n_210),
.B(n_199),
.C(n_201),
.D(n_161),
.Y(n_214)
);

NOR2xp33_ASAP7_75t_L g215 ( 
.A(n_211),
.B(n_212),
.Y(n_215)
);

XNOR2xp5_ASAP7_75t_L g212 ( 
.A(n_200),
.B(n_186),
.Y(n_212)
);

NOR2xp33_ASAP7_75t_L g216 ( 
.A(n_213),
.B(n_166),
.Y(n_216)
);

AO21x1_ASAP7_75t_L g222 ( 
.A1(n_214),
.A2(n_212),
.B(n_175),
.Y(n_222)
);

NOR2xp33_ASAP7_75t_SL g220 ( 
.A(n_216),
.B(n_208),
.Y(n_220)
);

INVxp67_ASAP7_75t_L g219 ( 
.A(n_207),
.Y(n_219)
);

NOR2xp33_ASAP7_75t_L g223 ( 
.A(n_219),
.B(n_175),
.Y(n_223)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_220),
.Y(n_225)
);

AOI22xp5_ASAP7_75t_L g221 ( 
.A1(n_217),
.A2(n_209),
.B1(n_206),
.B2(n_205),
.Y(n_221)
);

XNOR2xp5_ASAP7_75t_L g226 ( 
.A(n_221),
.B(n_222),
.Y(n_226)
);

HB1xp67_ASAP7_75t_L g227 ( 
.A(n_223),
.Y(n_227)
);

NOR2xp33_ASAP7_75t_L g224 ( 
.A(n_219),
.B(n_6),
.Y(n_224)
);

CKINVDCx20_ASAP7_75t_R g228 ( 
.A(n_227),
.Y(n_228)
);

AOI322xp5_ASAP7_75t_L g230 ( 
.A1(n_228),
.A2(n_229),
.A3(n_223),
.B1(n_224),
.B2(n_215),
.C1(n_225),
.C2(n_89),
.Y(n_230)
);

XOR2xp5_ASAP7_75t_L g229 ( 
.A(n_226),
.B(n_218),
.Y(n_229)
);

XOR2xp5_ASAP7_75t_L g231 ( 
.A(n_230),
.B(n_110),
.Y(n_231)
);


endmodule