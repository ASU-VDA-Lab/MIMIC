module fake_netlist_1_2158_n_23 (n_1, n_2, n_6, n_4, n_3, n_5, n_0, n_23);
input n_1;
input n_2;
input n_6;
input n_4;
input n_3;
input n_5;
input n_0;
output n_23;
wire n_20;
wire n_8;
wire n_22;
wire n_11;
wire n_16;
wire n_13;
wire n_18;
wire n_12;
wire n_9;
wire n_17;
wire n_14;
wire n_10;
wire n_15;
wire n_19;
wire n_21;
wire n_7;
NAND2xp5_ASAP7_75t_L g7 ( .A(n_3), .B(n_6), .Y(n_7) );
INVx2_ASAP7_75t_L g8 ( .A(n_4), .Y(n_8) );
INVx1_ASAP7_75t_L g9 ( .A(n_0), .Y(n_9) );
INVx1_ASAP7_75t_L g10 ( .A(n_5), .Y(n_10) );
INVx2_ASAP7_75t_L g11 ( .A(n_1), .Y(n_11) );
CKINVDCx8_ASAP7_75t_R g12 ( .A(n_7), .Y(n_12) );
NOR2xp67_ASAP7_75t_SL g13 ( .A(n_7), .B(n_0), .Y(n_13) );
BUFx2_ASAP7_75t_L g14 ( .A(n_9), .Y(n_14) );
INVx2_ASAP7_75t_L g15 ( .A(n_14), .Y(n_15) );
INVx3_ASAP7_75t_L g16 ( .A(n_12), .Y(n_16) );
INVx2_ASAP7_75t_L g17 ( .A(n_15), .Y(n_17) );
INVx2_ASAP7_75t_L g18 ( .A(n_16), .Y(n_18) );
OAI221xp5_ASAP7_75t_SL g19 ( .A1(n_17), .A2(n_16), .B1(n_11), .B2(n_10), .C(n_8), .Y(n_19) );
INVx1_ASAP7_75t_SL g20 ( .A(n_19), .Y(n_20) );
NAND3xp33_ASAP7_75t_SL g21 ( .A(n_19), .B(n_12), .C(n_18), .Y(n_21) );
OAI22xp5_ASAP7_75t_L g22 ( .A1(n_20), .A2(n_13), .B1(n_1), .B2(n_2), .Y(n_22) );
NAND2xp33_ASAP7_75t_L g23 ( .A(n_22), .B(n_21), .Y(n_23) );
endmodule