module real_jpeg_23015_n_18 (n_17, n_8, n_0, n_2, n_10, n_9, n_12, n_369, n_6, n_11, n_14, n_7, n_3, n_5, n_4, n_1, n_16, n_15, n_13, n_18);

input n_17;
input n_8;
input n_0;
input n_2;
input n_10;
input n_9;
input n_12;
input n_369;
input n_6;
input n_11;
input n_14;
input n_7;
input n_3;
input n_5;
input n_4;
input n_1;
input n_16;
input n_15;
input n_13;

output n_18;

wire n_37;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_300;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_199;
wire n_95;
wire n_238;
wire n_67;
wire n_350;
wire n_235;
wire n_107;
wire n_354;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_355;
wire n_123;
wire n_50;
wire n_186;
wire n_137;
wire n_72;
wire n_171;
wire n_151;
wire n_272;
wire n_198;
wire n_203;
wire n_23;
wire n_362;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_326;
wire n_339;
wire n_80;
wire n_30;
wire n_332;
wire n_149;
wire n_366;
wire n_328;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_353;
wire n_230;
wire n_128;
wire n_202;
wire n_216;
wire n_127;
wire n_365;
wire n_356;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_348;
wire n_252;
wire n_363;
wire n_310;
wire n_345;
wire n_78;
wire n_83;
wire n_288;
wire n_221;
wire n_104;
wire n_153;
wire n_337;
wire n_131;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_200;
wire n_335;
wire n_214;
wire n_113;
wire n_251;
wire n_139;
wire n_33;
wire n_175;
wire n_338;
wire n_156;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_77;
wire n_219;
wire n_122;
wire n_19;
wire n_262;
wire n_334;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_20;
wire n_278;
wire n_314;
wire n_103;
wire n_232;
wire n_212;
wire n_284;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_213;
wire n_25;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_341;
wire n_331;
wire n_49;
wire n_68;
wire n_146;
wire n_323;
wire n_166;
wire n_176;
wire n_215;
wire n_286;
wire n_312;
wire n_325;
wire n_307;
wire n_316;
wire n_161;
wire n_207;
wire n_357;
wire n_237;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_140;
wire n_126;
wire n_342;
wire n_120;
wire n_155;
wire n_319;
wire n_93;
wire n_242;
wire n_142;
wire n_76;
wire n_79;
wire n_282;
wire n_147;
wire n_359;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_145;
wire n_266;
wire n_109;
wire n_148;
wire n_196;
wire n_298;
wire n_330;
wire n_333;
wire n_152;
wire n_270;
wire n_159;
wire n_347;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_336;
wire n_258;
wire n_150;
wire n_41;
wire n_74;
wire n_204;
wire n_158;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_75;
wire n_346;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_119;
wire n_283;
wire n_181;
wire n_358;
wire n_256;
wire n_253;
wire n_273;
wire n_54;
wire n_168;
wire n_38;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_349;
wire n_292;
wire n_343;
wire n_64;
wire n_291;
wire n_236;
wire n_276;
wire n_287;
wire n_174;
wire n_255;
wire n_243;
wire n_299;
wire n_352;
wire n_56;
wire n_293;
wire n_275;
wire n_227;
wire n_229;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_360;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_45;
wire n_268;
wire n_42;
wire n_313;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_143;
wire n_351;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_303;
wire n_321;
wire n_100;
wire n_51;
wire n_205;
wire n_361;
wire n_261;
wire n_86;
wire n_324;
wire n_70;
wire n_32;
wire n_228;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_133;
wire n_257;
wire n_344;
wire n_210;
wire n_206;
wire n_85;
wire n_96;
wire n_308;
wire n_364;

BUFx6f_ASAP7_75t_L g114 ( 
.A(n_0),
.Y(n_114)
);

AOI22xp33_ASAP7_75t_L g34 ( 
.A1(n_1),
.A2(n_35),
.B1(n_36),
.B2(n_38),
.Y(n_34)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_1),
.Y(n_38)
);

AOI21xp5_ASAP7_75t_L g53 ( 
.A1(n_1),
.A2(n_42),
.B(n_47),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_L g57 ( 
.A(n_1),
.B(n_58),
.Y(n_57)
);

OAI22xp5_ASAP7_75t_SL g98 ( 
.A1(n_1),
.A2(n_68),
.B1(n_93),
.B2(n_99),
.Y(n_98)
);

AOI21xp5_ASAP7_75t_L g110 ( 
.A1(n_1),
.A2(n_111),
.B(n_115),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_L g148 ( 
.A(n_1),
.B(n_149),
.Y(n_148)
);

OAI22xp5_ASAP7_75t_L g75 ( 
.A1(n_2),
.A2(n_46),
.B1(n_47),
.B2(n_76),
.Y(n_75)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_2),
.Y(n_76)
);

OAI22xp5_ASAP7_75t_L g167 ( 
.A1(n_2),
.A2(n_35),
.B1(n_36),
.B2(n_76),
.Y(n_167)
);

AOI22xp5_ASAP7_75t_L g219 ( 
.A1(n_2),
.A2(n_76),
.B1(n_111),
.B2(n_112),
.Y(n_219)
);

OAI22xp5_ASAP7_75t_SL g266 ( 
.A1(n_2),
.A2(n_76),
.B1(n_181),
.B2(n_267),
.Y(n_266)
);

BUFx12f_ASAP7_75t_L g43 ( 
.A(n_3),
.Y(n_43)
);

AOI22xp33_ASAP7_75t_L g18 ( 
.A1(n_4),
.A2(n_13),
.B1(n_19),
.B2(n_20),
.Y(n_18)
);

CKINVDCx12_ASAP7_75t_R g19 ( 
.A(n_4),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_5),
.Y(n_48)
);

OAI22xp5_ASAP7_75t_L g50 ( 
.A1(n_6),
.A2(n_35),
.B1(n_36),
.B2(n_51),
.Y(n_50)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_6),
.Y(n_51)
);

AOI22xp33_ASAP7_75t_L g93 ( 
.A1(n_6),
.A2(n_46),
.B1(n_47),
.B2(n_51),
.Y(n_93)
);

AOI22xp33_ASAP7_75t_L g120 ( 
.A1(n_6),
.A2(n_51),
.B1(n_111),
.B2(n_112),
.Y(n_120)
);

OAI22xp5_ASAP7_75t_SL g208 ( 
.A1(n_6),
.A2(n_51),
.B1(n_179),
.B2(n_207),
.Y(n_208)
);

INVx8_ASAP7_75t_SL g153 ( 
.A(n_7),
.Y(n_153)
);

OAI22xp5_ASAP7_75t_L g186 ( 
.A1(n_8),
.A2(n_46),
.B1(n_47),
.B2(n_187),
.Y(n_186)
);

CKINVDCx20_ASAP7_75t_R g187 ( 
.A(n_8),
.Y(n_187)
);

AOI22xp5_ASAP7_75t_L g247 ( 
.A1(n_8),
.A2(n_35),
.B1(n_36),
.B2(n_187),
.Y(n_247)
);

OAI22xp5_ASAP7_75t_L g284 ( 
.A1(n_8),
.A2(n_111),
.B1(n_112),
.B2(n_187),
.Y(n_284)
);

OAI22xp5_ASAP7_75t_L g333 ( 
.A1(n_8),
.A2(n_177),
.B1(n_187),
.B2(n_297),
.Y(n_333)
);

AOI22xp5_ASAP7_75t_L g72 ( 
.A1(n_9),
.A2(n_46),
.B1(n_47),
.B2(n_73),
.Y(n_72)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_9),
.Y(n_73)
);

OAI22xp5_ASAP7_75t_L g122 ( 
.A1(n_9),
.A2(n_35),
.B1(n_36),
.B2(n_73),
.Y(n_122)
);

OAI22xp5_ASAP7_75t_L g196 ( 
.A1(n_9),
.A2(n_73),
.B1(n_111),
.B2(n_112),
.Y(n_196)
);

AOI22xp5_ASAP7_75t_SL g239 ( 
.A1(n_9),
.A2(n_73),
.B1(n_179),
.B2(n_207),
.Y(n_239)
);

OAI22xp5_ASAP7_75t_SL g133 ( 
.A1(n_10),
.A2(n_46),
.B1(n_47),
.B2(n_134),
.Y(n_133)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_10),
.Y(n_134)
);

AOI22xp5_ASAP7_75t_L g199 ( 
.A1(n_10),
.A2(n_35),
.B1(n_36),
.B2(n_134),
.Y(n_199)
);

OAI22xp5_ASAP7_75t_SL g242 ( 
.A1(n_10),
.A2(n_111),
.B1(n_112),
.B2(n_134),
.Y(n_242)
);

OAI22xp5_ASAP7_75t_SL g295 ( 
.A1(n_10),
.A2(n_134),
.B1(n_207),
.B2(n_296),
.Y(n_295)
);

BUFx12f_ASAP7_75t_L g60 ( 
.A(n_11),
.Y(n_60)
);

OAI22xp5_ASAP7_75t_L g64 ( 
.A1(n_12),
.A2(n_35),
.B1(n_36),
.B2(n_65),
.Y(n_64)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_12),
.Y(n_65)
);

AOI22xp33_ASAP7_75t_L g83 ( 
.A1(n_12),
.A2(n_46),
.B1(n_47),
.B2(n_65),
.Y(n_83)
);

OAI22xp5_ASAP7_75t_L g145 ( 
.A1(n_12),
.A2(n_65),
.B1(n_111),
.B2(n_112),
.Y(n_145)
);

AOI22xp33_ASAP7_75t_SL g222 ( 
.A1(n_12),
.A2(n_65),
.B1(n_204),
.B2(n_207),
.Y(n_222)
);

AOI22xp33_ASAP7_75t_L g158 ( 
.A1(n_14),
.A2(n_46),
.B1(n_47),
.B2(n_159),
.Y(n_158)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_14),
.Y(n_159)
);

AOI22xp5_ASAP7_75t_SL g228 ( 
.A1(n_14),
.A2(n_35),
.B1(n_36),
.B2(n_159),
.Y(n_228)
);

AOI22xp33_ASAP7_75t_SL g269 ( 
.A1(n_14),
.A2(n_111),
.B1(n_112),
.B2(n_159),
.Y(n_269)
);

AOI22xp33_ASAP7_75t_SL g317 ( 
.A1(n_14),
.A2(n_159),
.B1(n_181),
.B2(n_296),
.Y(n_317)
);

INVx13_ASAP7_75t_L g179 ( 
.A(n_15),
.Y(n_179)
);

BUFx12f_ASAP7_75t_L g37 ( 
.A(n_16),
.Y(n_37)
);

INVx3_ASAP7_75t_L g71 ( 
.A(n_17),
.Y(n_71)
);

INVx2_ASAP7_75t_L g78 ( 
.A(n_17),
.Y(n_78)
);

INVx6_ASAP7_75t_L g86 ( 
.A(n_17),
.Y(n_86)
);

INVx6_ASAP7_75t_L g96 ( 
.A(n_17),
.Y(n_96)
);

MAJIxp5_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_365),
.C(n_366),
.Y(n_20)
);

OAI21xp5_ASAP7_75t_SL g21 ( 
.A1(n_22),
.A2(n_361),
.B(n_364),
.Y(n_21)
);

AOI21xp5_ASAP7_75t_L g22 ( 
.A1(n_23),
.A2(n_347),
.B(n_360),
.Y(n_22)
);

OAI321xp33_ASAP7_75t_L g23 ( 
.A1(n_24),
.A2(n_312),
.A3(n_340),
.B1(n_345),
.B2(n_346),
.C(n_369),
.Y(n_23)
);

AOI311xp33_ASAP7_75t_L g24 ( 
.A1(n_25),
.A2(n_257),
.A3(n_302),
.B(n_306),
.C(n_307),
.Y(n_24)
);

NOR3xp33_ASAP7_75t_L g25 ( 
.A(n_26),
.B(n_210),
.C(n_252),
.Y(n_25)
);

AOI21xp5_ASAP7_75t_L g26 ( 
.A1(n_27),
.A2(n_171),
.B(n_209),
.Y(n_26)
);

OAI21xp5_ASAP7_75t_SL g27 ( 
.A1(n_28),
.A2(n_138),
.B(n_170),
.Y(n_27)
);

AOI21xp5_ASAP7_75t_L g28 ( 
.A1(n_29),
.A2(n_105),
.B(n_137),
.Y(n_28)
);

OAI21xp5_ASAP7_75t_SL g29 ( 
.A1(n_30),
.A2(n_79),
.B(n_104),
.Y(n_29)
);

NOR2xp33_ASAP7_75t_L g30 ( 
.A(n_31),
.B(n_54),
.Y(n_30)
);

NAND2xp5_ASAP7_75t_SL g104 ( 
.A(n_31),
.B(n_54),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_SL g31 ( 
.A(n_32),
.B(n_52),
.Y(n_31)
);

AOI22xp5_ASAP7_75t_SL g87 ( 
.A1(n_32),
.A2(n_33),
.B1(n_52),
.B2(n_88),
.Y(n_87)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_33),
.Y(n_32)
);

OAI22xp5_ASAP7_75t_L g33 ( 
.A1(n_34),
.A2(n_39),
.B1(n_45),
.B2(n_49),
.Y(n_33)
);

OAI22xp33_ASAP7_75t_L g41 ( 
.A1(n_35),
.A2(n_36),
.B1(n_42),
.B2(n_44),
.Y(n_41)
);

AOI22xp5_ASAP7_75t_L g59 ( 
.A1(n_35),
.A2(n_36),
.B1(n_60),
.B2(n_61),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_SL g127 ( 
.A(n_35),
.B(n_61),
.Y(n_127)
);

INVx8_ASAP7_75t_L g35 ( 
.A(n_36),
.Y(n_35)
);

A2O1A1Ixp33_ASAP7_75t_SL g52 ( 
.A1(n_36),
.A2(n_38),
.B(n_44),
.C(n_53),
.Y(n_52)
);

OAI32xp33_ASAP7_75t_L g126 ( 
.A1(n_36),
.A2(n_60),
.A3(n_111),
.B1(n_116),
.B2(n_127),
.Y(n_126)
);

BUFx12f_ASAP7_75t_L g36 ( 
.A(n_37),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_SL g91 ( 
.A(n_38),
.B(n_45),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_38),
.B(n_78),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_L g116 ( 
.A(n_38),
.B(n_112),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_L g180 ( 
.A(n_38),
.B(n_181),
.Y(n_180)
);

OAI21xp33_ASAP7_75t_L g206 ( 
.A1(n_38),
.A2(n_180),
.B(n_207),
.Y(n_206)
);

OAI21xp5_ASAP7_75t_SL g164 ( 
.A1(n_39),
.A2(n_165),
.B(n_166),
.Y(n_164)
);

OAI22xp5_ASAP7_75t_L g246 ( 
.A1(n_39),
.A2(n_45),
.B1(n_228),
.B2(n_247),
.Y(n_246)
);

OAI21xp5_ASAP7_75t_SL g275 ( 
.A1(n_39),
.A2(n_247),
.B(n_276),
.Y(n_275)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_40),
.Y(n_39)
);

AOI22xp5_ASAP7_75t_L g62 ( 
.A1(n_40),
.A2(n_50),
.B1(n_63),
.B2(n_64),
.Y(n_62)
);

AOI22xp5_ASAP7_75t_L g121 ( 
.A1(n_40),
.A2(n_63),
.B1(n_64),
.B2(n_122),
.Y(n_121)
);

AOI21xp5_ASAP7_75t_L g197 ( 
.A1(n_40),
.A2(n_167),
.B(n_198),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_L g229 ( 
.A(n_40),
.B(n_230),
.Y(n_229)
);

OAI21xp5_ASAP7_75t_SL g321 ( 
.A1(n_40),
.A2(n_63),
.B(n_167),
.Y(n_321)
);

AND2x2_ASAP7_75t_L g40 ( 
.A(n_41),
.B(n_45),
.Y(n_40)
);

INVx13_ASAP7_75t_L g44 ( 
.A(n_42),
.Y(n_44)
);

AOI22xp5_ASAP7_75t_L g45 ( 
.A1(n_42),
.A2(n_44),
.B1(n_46),
.B2(n_47),
.Y(n_45)
);

BUFx24_ASAP7_75t_L g42 ( 
.A(n_43),
.Y(n_42)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_45),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g198 ( 
.A(n_45),
.B(n_199),
.Y(n_198)
);

OAI21xp5_ASAP7_75t_L g227 ( 
.A1(n_45),
.A2(n_228),
.B(n_229),
.Y(n_227)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_46),
.B(n_70),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_SL g100 ( 
.A(n_46),
.B(n_101),
.Y(n_100)
);

INVx5_ASAP7_75t_L g46 ( 
.A(n_47),
.Y(n_46)
);

BUFx12f_ASAP7_75t_L g47 ( 
.A(n_48),
.Y(n_47)
);

CKINVDCx16_ASAP7_75t_R g49 ( 
.A(n_50),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g88 ( 
.A(n_52),
.Y(n_88)
);

XNOR2xp5_ASAP7_75t_L g54 ( 
.A(n_55),
.B(n_67),
.Y(n_54)
);

AOI22xp5_ASAP7_75t_L g55 ( 
.A1(n_56),
.A2(n_57),
.B1(n_62),
.B2(n_66),
.Y(n_55)
);

MAJIxp5_ASAP7_75t_L g106 ( 
.A(n_56),
.B(n_66),
.C(n_67),
.Y(n_106)
);

CKINVDCx14_ASAP7_75t_R g56 ( 
.A(n_57),
.Y(n_56)
);

AOI22xp5_ASAP7_75t_L g143 ( 
.A1(n_58),
.A2(n_118),
.B1(n_144),
.B2(n_145),
.Y(n_143)
);

AOI22xp5_ASAP7_75t_L g195 ( 
.A1(n_58),
.A2(n_118),
.B1(n_145),
.B2(n_196),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_L g241 ( 
.A(n_58),
.B(n_242),
.Y(n_241)
);

AOI22xp5_ASAP7_75t_L g282 ( 
.A1(n_58),
.A2(n_118),
.B1(n_283),
.B2(n_284),
.Y(n_282)
);

OAI21xp5_ASAP7_75t_L g356 ( 
.A1(n_58),
.A2(n_118),
.B(n_357),
.Y(n_356)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_59),
.Y(n_58)
);

OAI22xp5_ASAP7_75t_L g109 ( 
.A1(n_59),
.A2(n_110),
.B1(n_117),
.B2(n_120),
.Y(n_109)
);

AND2x2_ASAP7_75t_L g118 ( 
.A(n_59),
.B(n_119),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_L g218 ( 
.A(n_59),
.B(n_219),
.Y(n_218)
);

OAI21xp5_ASAP7_75t_L g268 ( 
.A1(n_59),
.A2(n_269),
.B(n_270),
.Y(n_268)
);

INVx5_ASAP7_75t_L g61 ( 
.A(n_60),
.Y(n_61)
);

OAI22xp5_ASAP7_75t_L g119 ( 
.A1(n_60),
.A2(n_61),
.B1(n_111),
.B2(n_112),
.Y(n_119)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_62),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_SL g166 ( 
.A(n_63),
.B(n_167),
.Y(n_166)
);

OAI21xp5_ASAP7_75t_L g67 ( 
.A1(n_68),
.A2(n_72),
.B(n_74),
.Y(n_67)
);

OAI22xp5_ASAP7_75t_SL g92 ( 
.A1(n_68),
.A2(n_83),
.B1(n_93),
.B2(n_94),
.Y(n_92)
);

OAI21xp5_ASAP7_75t_L g128 ( 
.A1(n_68),
.A2(n_129),
.B(n_130),
.Y(n_128)
);

OAI21xp5_ASAP7_75t_L g225 ( 
.A1(n_68),
.A2(n_130),
.B(n_226),
.Y(n_225)
);

AOI21xp5_ASAP7_75t_L g273 ( 
.A1(n_68),
.A2(n_94),
.B(n_129),
.Y(n_273)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_69),
.Y(n_68)
);

AOI22xp5_ASAP7_75t_SL g81 ( 
.A1(n_69),
.A2(n_82),
.B1(n_84),
.B2(n_85),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_SL g160 ( 
.A(n_69),
.B(n_133),
.Y(n_160)
);

AOI22xp5_ASAP7_75t_L g183 ( 
.A1(n_69),
.A2(n_184),
.B1(n_185),
.B2(n_186),
.Y(n_183)
);

INVx3_ASAP7_75t_L g70 ( 
.A(n_71),
.Y(n_70)
);

CKINVDCx20_ASAP7_75t_R g84 ( 
.A(n_72),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g245 ( 
.A(n_74),
.B(n_160),
.Y(n_245)
);

NAND2xp5_ASAP7_75t_SL g74 ( 
.A(n_75),
.B(n_77),
.Y(n_74)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_75),
.Y(n_129)
);

INVx2_ASAP7_75t_L g77 ( 
.A(n_78),
.Y(n_77)
);

BUFx2_ASAP7_75t_L g132 ( 
.A(n_78),
.Y(n_132)
);

AOI21xp5_ASAP7_75t_L g79 ( 
.A1(n_80),
.A2(n_89),
.B(n_103),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_L g80 ( 
.A(n_81),
.B(n_87),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_SL g103 ( 
.A(n_81),
.B(n_87),
.Y(n_103)
);

CKINVDCx16_ASAP7_75t_R g82 ( 
.A(n_83),
.Y(n_82)
);

INVx5_ASAP7_75t_L g99 ( 
.A(n_85),
.Y(n_99)
);

INVx5_ASAP7_75t_L g85 ( 
.A(n_86),
.Y(n_85)
);

OAI21xp5_ASAP7_75t_SL g89 ( 
.A1(n_90),
.A2(n_97),
.B(n_102),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_91),
.B(n_92),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_SL g102 ( 
.A(n_91),
.B(n_92),
.Y(n_102)
);

INVx3_ASAP7_75t_L g185 ( 
.A(n_94),
.Y(n_185)
);

INVx5_ASAP7_75t_L g94 ( 
.A(n_95),
.Y(n_94)
);

INVx8_ASAP7_75t_L g95 ( 
.A(n_96),
.Y(n_95)
);

INVx5_ASAP7_75t_L g157 ( 
.A(n_96),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_SL g97 ( 
.A(n_98),
.B(n_100),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g105 ( 
.A(n_106),
.B(n_107),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_SL g137 ( 
.A(n_106),
.B(n_107),
.Y(n_137)
);

AOI22xp5_ASAP7_75t_SL g107 ( 
.A1(n_108),
.A2(n_125),
.B1(n_135),
.B2(n_136),
.Y(n_107)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_108),
.Y(n_136)
);

AOI22xp5_ASAP7_75t_L g108 ( 
.A1(n_109),
.A2(n_121),
.B1(n_123),
.B2(n_124),
.Y(n_108)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_109),
.Y(n_124)
);

AOI22xp5_ASAP7_75t_L g150 ( 
.A1(n_111),
.A2(n_112),
.B1(n_151),
.B2(n_152),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_L g182 ( 
.A(n_111),
.B(n_152),
.Y(n_182)
);

CKINVDCx20_ASAP7_75t_R g111 ( 
.A(n_112),
.Y(n_111)
);

OAI32xp33_ASAP7_75t_L g176 ( 
.A1(n_112),
.A2(n_151),
.A3(n_177),
.B1(n_180),
.B2(n_182),
.Y(n_176)
);

BUFx12f_ASAP7_75t_L g112 ( 
.A(n_113),
.Y(n_112)
);

BUFx12f_ASAP7_75t_L g113 ( 
.A(n_114),
.Y(n_113)
);

CKINVDCx20_ASAP7_75t_R g115 ( 
.A(n_116),
.Y(n_115)
);

OAI21xp5_ASAP7_75t_SL g240 ( 
.A1(n_117),
.A2(n_219),
.B(n_241),
.Y(n_240)
);

CKINVDCx20_ASAP7_75t_R g117 ( 
.A(n_118),
.Y(n_117)
);

AOI21xp5_ASAP7_75t_L g217 ( 
.A1(n_118),
.A2(n_196),
.B(n_218),
.Y(n_217)
);

NAND2xp5_ASAP7_75t_SL g270 ( 
.A(n_118),
.B(n_242),
.Y(n_270)
);

AOI21xp5_ASAP7_75t_L g322 ( 
.A1(n_118),
.A2(n_284),
.B(n_323),
.Y(n_322)
);

CKINVDCx14_ASAP7_75t_R g144 ( 
.A(n_120),
.Y(n_144)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_121),
.Y(n_123)
);

MAJIxp5_ASAP7_75t_L g139 ( 
.A(n_121),
.B(n_124),
.C(n_135),
.Y(n_139)
);

CKINVDCx20_ASAP7_75t_R g165 ( 
.A(n_122),
.Y(n_165)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_125),
.Y(n_135)
);

XOR2xp5_ASAP7_75t_L g125 ( 
.A(n_126),
.B(n_128),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_L g163 ( 
.A(n_126),
.B(n_128),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_L g130 ( 
.A(n_131),
.B(n_133),
.Y(n_130)
);

CKINVDCx20_ASAP7_75t_R g131 ( 
.A(n_132),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_L g138 ( 
.A(n_139),
.B(n_140),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_SL g170 ( 
.A(n_139),
.B(n_140),
.Y(n_170)
);

OAI22xp5_ASAP7_75t_SL g140 ( 
.A1(n_141),
.A2(n_142),
.B1(n_161),
.B2(n_162),
.Y(n_140)
);

MAJIxp5_ASAP7_75t_L g172 ( 
.A(n_141),
.B(n_164),
.C(n_168),
.Y(n_172)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_142),
.Y(n_141)
);

XNOR2xp5_ASAP7_75t_SL g142 ( 
.A(n_143),
.B(n_146),
.Y(n_142)
);

MAJIxp5_ASAP7_75t_L g190 ( 
.A(n_143),
.B(n_148),
.C(n_154),
.Y(n_190)
);

AOI22xp5_ASAP7_75t_L g146 ( 
.A1(n_147),
.A2(n_148),
.B1(n_154),
.B2(n_155),
.Y(n_146)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_148),
.Y(n_147)
);

AOI22xp5_ASAP7_75t_SL g200 ( 
.A1(n_149),
.A2(n_201),
.B1(n_206),
.B2(n_208),
.Y(n_200)
);

AOI22xp5_ASAP7_75t_L g220 ( 
.A1(n_149),
.A2(n_201),
.B1(n_208),
.B2(n_221),
.Y(n_220)
);

NAND2xp5_ASAP7_75t_SL g265 ( 
.A(n_149),
.B(n_266),
.Y(n_265)
);

NAND2xp5_ASAP7_75t_SL g294 ( 
.A(n_149),
.B(n_295),
.Y(n_294)
);

AOI22xp5_ASAP7_75t_L g331 ( 
.A1(n_149),
.A2(n_201),
.B1(n_332),
.B2(n_333),
.Y(n_331)
);

OAI21xp5_ASAP7_75t_SL g365 ( 
.A1(n_149),
.A2(n_201),
.B(n_266),
.Y(n_365)
);

CKINVDCx16_ASAP7_75t_R g149 ( 
.A(n_150),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_SL g202 ( 
.A(n_150),
.B(n_203),
.Y(n_202)
);

OAI22xp5_ASAP7_75t_SL g238 ( 
.A1(n_150),
.A2(n_202),
.B1(n_222),
.B2(n_239),
.Y(n_238)
);

OAI21xp5_ASAP7_75t_L g316 ( 
.A1(n_150),
.A2(n_317),
.B(n_318),
.Y(n_316)
);

OAI22xp33_ASAP7_75t_L g203 ( 
.A1(n_151),
.A2(n_152),
.B1(n_204),
.B2(n_205),
.Y(n_203)
);

INVx4_ASAP7_75t_L g151 ( 
.A(n_152),
.Y(n_151)
);

BUFx6f_ASAP7_75t_L g152 ( 
.A(n_153),
.Y(n_152)
);

CKINVDCx16_ASAP7_75t_R g154 ( 
.A(n_155),
.Y(n_154)
);

OAI21xp5_ASAP7_75t_L g155 ( 
.A1(n_156),
.A2(n_158),
.B(n_160),
.Y(n_155)
);

INVx2_ASAP7_75t_L g156 ( 
.A(n_157),
.Y(n_156)
);

INVxp67_ASAP7_75t_L g184 ( 
.A(n_158),
.Y(n_184)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_162),
.Y(n_161)
);

OAI22xp5_ASAP7_75t_SL g162 ( 
.A1(n_163),
.A2(n_164),
.B1(n_168),
.B2(n_169),
.Y(n_162)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_163),
.Y(n_168)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_164),
.Y(n_169)
);

AND2x2_ASAP7_75t_L g285 ( 
.A(n_166),
.B(n_229),
.Y(n_285)
);

NAND2xp5_ASAP7_75t_L g171 ( 
.A(n_172),
.B(n_173),
.Y(n_171)
);

NOR2xp33_ASAP7_75t_SL g209 ( 
.A(n_172),
.B(n_173),
.Y(n_209)
);

XOR2xp5_ASAP7_75t_L g173 ( 
.A(n_174),
.B(n_193),
.Y(n_173)
);

OAI22xp5_ASAP7_75t_L g174 ( 
.A1(n_175),
.A2(n_190),
.B1(n_191),
.B2(n_192),
.Y(n_174)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_175),
.Y(n_191)
);

MAJIxp5_ASAP7_75t_L g253 ( 
.A(n_175),
.B(n_192),
.C(n_193),
.Y(n_253)
);

AOI22xp5_ASAP7_75t_L g175 ( 
.A1(n_176),
.A2(n_183),
.B1(n_188),
.B2(n_189),
.Y(n_175)
);

CKINVDCx14_ASAP7_75t_R g189 ( 
.A(n_176),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_L g215 ( 
.A(n_176),
.B(n_188),
.Y(n_215)
);

INVx8_ASAP7_75t_L g207 ( 
.A(n_177),
.Y(n_207)
);

INVx8_ASAP7_75t_L g177 ( 
.A(n_178),
.Y(n_177)
);

INVx6_ASAP7_75t_L g178 ( 
.A(n_179),
.Y(n_178)
);

INVx11_ASAP7_75t_L g181 ( 
.A(n_179),
.Y(n_181)
);

INVx8_ASAP7_75t_L g205 ( 
.A(n_179),
.Y(n_205)
);

INVx8_ASAP7_75t_L g297 ( 
.A(n_179),
.Y(n_297)
);

INVx8_ASAP7_75t_L g267 ( 
.A(n_181),
.Y(n_267)
);

CKINVDCx20_ASAP7_75t_R g188 ( 
.A(n_183),
.Y(n_188)
);

INVxp67_ASAP7_75t_L g226 ( 
.A(n_186),
.Y(n_226)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_190),
.Y(n_192)
);

XOR2xp5_ASAP7_75t_L g193 ( 
.A(n_194),
.B(n_200),
.Y(n_193)
);

XOR2xp5_ASAP7_75t_L g194 ( 
.A(n_195),
.B(n_197),
.Y(n_194)
);

MAJIxp5_ASAP7_75t_L g223 ( 
.A(n_195),
.B(n_197),
.C(n_200),
.Y(n_223)
);

INVxp67_ASAP7_75t_L g276 ( 
.A(n_198),
.Y(n_276)
);

CKINVDCx20_ASAP7_75t_R g230 ( 
.A(n_199),
.Y(n_230)
);

NAND2xp5_ASAP7_75t_L g318 ( 
.A(n_201),
.B(n_295),
.Y(n_318)
);

AOI21xp5_ASAP7_75t_L g353 ( 
.A1(n_201),
.A2(n_333),
.B(n_354),
.Y(n_353)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_202),
.Y(n_201)
);

OAI21xp5_ASAP7_75t_SL g264 ( 
.A1(n_202),
.A2(n_239),
.B(n_265),
.Y(n_264)
);

OAI21xp5_ASAP7_75t_SL g292 ( 
.A1(n_202),
.A2(n_293),
.B(n_294),
.Y(n_292)
);

INVx4_ASAP7_75t_L g204 ( 
.A(n_205),
.Y(n_204)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_211),
.Y(n_210)
);

AOI21xp33_ASAP7_75t_L g308 ( 
.A1(n_211),
.A2(n_309),
.B(n_310),
.Y(n_308)
);

NAND2xp5_ASAP7_75t_L g211 ( 
.A(n_212),
.B(n_231),
.Y(n_211)
);

NOR2xp33_ASAP7_75t_SL g310 ( 
.A(n_212),
.B(n_231),
.Y(n_310)
);

MAJIxp5_ASAP7_75t_L g212 ( 
.A(n_213),
.B(n_223),
.C(n_224),
.Y(n_212)
);

OAI22xp5_ASAP7_75t_L g254 ( 
.A1(n_213),
.A2(n_214),
.B1(n_255),
.B2(n_256),
.Y(n_254)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_214),
.Y(n_213)
);

XOR2xp5_ASAP7_75t_L g214 ( 
.A(n_215),
.B(n_216),
.Y(n_214)
);

MAJIxp5_ASAP7_75t_L g249 ( 
.A(n_215),
.B(n_217),
.C(n_220),
.Y(n_249)
);

XOR2xp5_ASAP7_75t_L g216 ( 
.A(n_217),
.B(n_220),
.Y(n_216)
);

INVxp67_ASAP7_75t_L g337 ( 
.A(n_218),
.Y(n_337)
);

CKINVDCx16_ASAP7_75t_R g357 ( 
.A(n_219),
.Y(n_357)
);

INVxp67_ASAP7_75t_L g221 ( 
.A(n_222),
.Y(n_221)
);

XNOR2xp5_ASAP7_75t_SL g256 ( 
.A(n_223),
.B(n_224),
.Y(n_256)
);

XOR2xp5_ASAP7_75t_L g224 ( 
.A(n_225),
.B(n_227),
.Y(n_224)
);

NAND2xp5_ASAP7_75t_L g235 ( 
.A(n_225),
.B(n_227),
.Y(n_235)
);

AOI22xp5_ASAP7_75t_SL g231 ( 
.A1(n_232),
.A2(n_249),
.B1(n_250),
.B2(n_251),
.Y(n_231)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_232),
.Y(n_250)
);

AOI22xp5_ASAP7_75t_SL g232 ( 
.A1(n_233),
.A2(n_234),
.B1(n_244),
.B2(n_248),
.Y(n_232)
);

MAJIxp5_ASAP7_75t_L g304 ( 
.A(n_233),
.B(n_248),
.C(n_251),
.Y(n_304)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_234),
.Y(n_233)
);

OAI22xp5_ASAP7_75t_L g234 ( 
.A1(n_235),
.A2(n_236),
.B1(n_237),
.B2(n_243),
.Y(n_234)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_235),
.Y(n_243)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_237),
.Y(n_236)
);

XNOR2xp5_ASAP7_75t_SL g237 ( 
.A(n_238),
.B(n_240),
.Y(n_237)
);

MAJIxp5_ASAP7_75t_L g278 ( 
.A(n_238),
.B(n_240),
.C(n_243),
.Y(n_278)
);

INVxp67_ASAP7_75t_L g323 ( 
.A(n_241),
.Y(n_323)
);

CKINVDCx16_ASAP7_75t_R g248 ( 
.A(n_244),
.Y(n_248)
);

XOR2xp5_ASAP7_75t_L g244 ( 
.A(n_245),
.B(n_246),
.Y(n_244)
);

NAND2xp5_ASAP7_75t_L g262 ( 
.A(n_245),
.B(n_246),
.Y(n_262)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_249),
.Y(n_251)
);

NOR2xp33_ASAP7_75t_L g252 ( 
.A(n_253),
.B(n_254),
.Y(n_252)
);

AND2x2_ASAP7_75t_L g309 ( 
.A(n_253),
.B(n_254),
.Y(n_309)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_256),
.Y(n_255)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_258),
.Y(n_257)
);

O2A1O1Ixp33_ASAP7_75t_SL g307 ( 
.A1(n_258),
.A2(n_303),
.B(n_308),
.C(n_311),
.Y(n_307)
);

NOR2xp33_ASAP7_75t_L g258 ( 
.A(n_259),
.B(n_279),
.Y(n_258)
);

AND2x2_ASAP7_75t_L g306 ( 
.A(n_259),
.B(n_279),
.Y(n_306)
);

MAJIxp5_ASAP7_75t_L g259 ( 
.A(n_260),
.B(n_272),
.C(n_278),
.Y(n_259)
);

FAx1_ASAP7_75t_SL g305 ( 
.A(n_260),
.B(n_272),
.CI(n_278),
.CON(n_305),
.SN(n_305)
);

AOI22xp5_ASAP7_75t_L g260 ( 
.A1(n_261),
.A2(n_262),
.B1(n_263),
.B2(n_271),
.Y(n_260)
);

MAJIxp5_ASAP7_75t_L g301 ( 
.A(n_261),
.B(n_264),
.C(n_268),
.Y(n_301)
);

CKINVDCx14_ASAP7_75t_R g261 ( 
.A(n_262),
.Y(n_261)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_263),
.Y(n_271)
);

XNOR2xp5_ASAP7_75t_SL g263 ( 
.A(n_264),
.B(n_268),
.Y(n_263)
);

AND2x2_ASAP7_75t_L g362 ( 
.A(n_265),
.B(n_318),
.Y(n_362)
);

CKINVDCx16_ASAP7_75t_R g293 ( 
.A(n_266),
.Y(n_293)
);

CKINVDCx14_ASAP7_75t_R g283 ( 
.A(n_269),
.Y(n_283)
);

NAND2xp5_ASAP7_75t_L g336 ( 
.A(n_270),
.B(n_337),
.Y(n_336)
);

AOI22xp5_ASAP7_75t_L g272 ( 
.A1(n_273),
.A2(n_274),
.B1(n_275),
.B2(n_277),
.Y(n_272)
);

CKINVDCx16_ASAP7_75t_R g277 ( 
.A(n_273),
.Y(n_277)
);

NAND2xp5_ASAP7_75t_L g289 ( 
.A(n_273),
.B(n_275),
.Y(n_289)
);

AOI22xp5_ASAP7_75t_L g290 ( 
.A1(n_273),
.A2(n_277),
.B1(n_291),
.B2(n_292),
.Y(n_290)
);

INVxp67_ASAP7_75t_L g274 ( 
.A(n_275),
.Y(n_274)
);

OAI21xp5_ASAP7_75t_L g327 ( 
.A1(n_277),
.A2(n_288),
.B(n_292),
.Y(n_327)
);

XOR2xp5_ASAP7_75t_L g279 ( 
.A(n_280),
.B(n_301),
.Y(n_279)
);

AOI22xp5_ASAP7_75t_L g280 ( 
.A1(n_281),
.A2(n_287),
.B1(n_299),
.B2(n_300),
.Y(n_280)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_281),
.Y(n_299)
);

OAI21xp5_ASAP7_75t_L g281 ( 
.A1(n_282),
.A2(n_285),
.B(n_286),
.Y(n_281)
);

NAND2xp5_ASAP7_75t_SL g286 ( 
.A(n_282),
.B(n_285),
.Y(n_286)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_286),
.Y(n_326)
);

AOI22xp5_ASAP7_75t_L g343 ( 
.A1(n_286),
.A2(n_314),
.B1(n_326),
.B2(n_344),
.Y(n_343)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_287),
.Y(n_300)
);

MAJIxp5_ASAP7_75t_L g341 ( 
.A(n_287),
.B(n_299),
.C(n_301),
.Y(n_341)
);

AOI22xp5_ASAP7_75t_L g287 ( 
.A1(n_288),
.A2(n_289),
.B1(n_290),
.B2(n_298),
.Y(n_287)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_289),
.Y(n_288)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_290),
.Y(n_298)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_292),
.Y(n_291)
);

INVxp67_ASAP7_75t_L g354 ( 
.A(n_294),
.Y(n_354)
);

INVx11_ASAP7_75t_L g296 ( 
.A(n_297),
.Y(n_296)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_303),
.Y(n_302)
);

NOR2xp33_ASAP7_75t_L g303 ( 
.A(n_304),
.B(n_305),
.Y(n_303)
);

NAND2xp5_ASAP7_75t_SL g311 ( 
.A(n_304),
.B(n_305),
.Y(n_311)
);

BUFx24_ASAP7_75t_SL g367 ( 
.A(n_305),
.Y(n_367)
);

NOR2xp33_ASAP7_75t_L g312 ( 
.A(n_313),
.B(n_328),
.Y(n_312)
);

NAND2xp5_ASAP7_75t_SL g346 ( 
.A(n_313),
.B(n_328),
.Y(n_346)
);

MAJIxp5_ASAP7_75t_L g313 ( 
.A(n_314),
.B(n_326),
.C(n_327),
.Y(n_313)
);

INVx1_ASAP7_75t_L g344 ( 
.A(n_314),
.Y(n_344)
);

AOI22xp5_ASAP7_75t_L g314 ( 
.A1(n_315),
.A2(n_316),
.B1(n_319),
.B2(n_325),
.Y(n_314)
);

AOI22xp5_ASAP7_75t_L g329 ( 
.A1(n_315),
.A2(n_316),
.B1(n_330),
.B2(n_338),
.Y(n_329)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_316),
.Y(n_315)
);

MAJIxp5_ASAP7_75t_L g339 ( 
.A(n_316),
.B(n_321),
.C(n_322),
.Y(n_339)
);

MAJIxp5_ASAP7_75t_L g359 ( 
.A(n_316),
.B(n_338),
.C(n_339),
.Y(n_359)
);

CKINVDCx20_ASAP7_75t_R g332 ( 
.A(n_317),
.Y(n_332)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_319),
.Y(n_325)
);

AOI22xp5_ASAP7_75t_L g319 ( 
.A1(n_320),
.A2(n_321),
.B1(n_322),
.B2(n_324),
.Y(n_319)
);

AOI22xp5_ASAP7_75t_L g334 ( 
.A1(n_320),
.A2(n_321),
.B1(n_335),
.B2(n_336),
.Y(n_334)
);

MAJIxp5_ASAP7_75t_L g350 ( 
.A(n_320),
.B(n_331),
.C(n_335),
.Y(n_350)
);

CKINVDCx16_ASAP7_75t_R g320 ( 
.A(n_321),
.Y(n_320)
);

CKINVDCx20_ASAP7_75t_R g324 ( 
.A(n_322),
.Y(n_324)
);

XOR2xp5_ASAP7_75t_L g342 ( 
.A(n_327),
.B(n_343),
.Y(n_342)
);

XNOR2xp5_ASAP7_75t_L g328 ( 
.A(n_329),
.B(n_339),
.Y(n_328)
);

INVx1_ASAP7_75t_L g338 ( 
.A(n_330),
.Y(n_338)
);

XNOR2xp5_ASAP7_75t_SL g330 ( 
.A(n_331),
.B(n_334),
.Y(n_330)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_336),
.Y(n_335)
);

NOR2xp33_ASAP7_75t_L g340 ( 
.A(n_341),
.B(n_342),
.Y(n_340)
);

NAND2xp5_ASAP7_75t_SL g345 ( 
.A(n_341),
.B(n_342),
.Y(n_345)
);

NAND2xp5_ASAP7_75t_L g347 ( 
.A(n_348),
.B(n_359),
.Y(n_347)
);

NOR2xp33_ASAP7_75t_SL g360 ( 
.A(n_348),
.B(n_359),
.Y(n_360)
);

AOI22xp5_ASAP7_75t_SL g348 ( 
.A1(n_349),
.A2(n_350),
.B1(n_351),
.B2(n_358),
.Y(n_348)
);

MAJIxp5_ASAP7_75t_L g363 ( 
.A(n_349),
.B(n_353),
.C(n_355),
.Y(n_363)
);

CKINVDCx20_ASAP7_75t_R g349 ( 
.A(n_350),
.Y(n_349)
);

INVx1_ASAP7_75t_L g358 ( 
.A(n_351),
.Y(n_358)
);

OAI22xp5_ASAP7_75t_L g351 ( 
.A1(n_352),
.A2(n_353),
.B1(n_355),
.B2(n_356),
.Y(n_351)
);

CKINVDCx20_ASAP7_75t_R g352 ( 
.A(n_353),
.Y(n_352)
);

CKINVDCx20_ASAP7_75t_R g355 ( 
.A(n_356),
.Y(n_355)
);

NOR2xp33_ASAP7_75t_L g361 ( 
.A(n_362),
.B(n_363),
.Y(n_361)
);

NAND2xp5_ASAP7_75t_SL g364 ( 
.A(n_362),
.B(n_363),
.Y(n_364)
);

CKINVDCx20_ASAP7_75t_R g366 ( 
.A(n_362),
.Y(n_366)
);


endmodule