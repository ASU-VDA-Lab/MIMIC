module fake_jpeg_20035_n_292 (n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_292);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_292;

wire n_159;
wire n_117;
wire n_253;
wire n_286;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_14;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_84;
wire n_59;
wire n_98;
wire n_251;
wire n_252;
wire n_273;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_279;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_278;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_281;
wire n_31;
wire n_155;
wire n_207;
wire n_277;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_291;
wire n_236;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_13;
wire n_175;
wire n_223;
wire n_21;
wire n_57;
wire n_187;
wire n_234;
wire n_284;
wire n_272;
wire n_288;
wire n_280;
wire n_171;
wire n_263;
wire n_119;
wire n_23;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_289;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_267;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_274;
wire n_186;
wire n_24;
wire n_44;
wire n_276;
wire n_143;
wire n_202;
wire n_25;
wire n_17;
wire n_269;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_287;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_266;
wire n_34;
wire n_283;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_285;
wire n_215;
wire n_262;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_271;
wire n_217;
wire n_216;
wire n_264;
wire n_184;
wire n_53;
wire n_268;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_265;
wire n_176;
wire n_199;
wire n_112;
wire n_260;
wire n_270;
wire n_222;
wire n_95;
wire n_275;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_290;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_258;
wire n_282;
wire n_96;

BUFx3_ASAP7_75t_L g13 ( 
.A(n_4),
.Y(n_13)
);

CKINVDCx20_ASAP7_75t_R g14 ( 
.A(n_2),
.Y(n_14)
);

INVx4_ASAP7_75t_L g15 ( 
.A(n_2),
.Y(n_15)
);

INVx6_ASAP7_75t_L g16 ( 
.A(n_3),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_12),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_10),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_1),
.Y(n_19)
);

INVx2_ASAP7_75t_L g20 ( 
.A(n_9),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_8),
.Y(n_21)
);

BUFx12f_ASAP7_75t_L g22 ( 
.A(n_12),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_11),
.Y(n_23)
);

BUFx12_ASAP7_75t_L g24 ( 
.A(n_12),
.Y(n_24)
);

INVx13_ASAP7_75t_L g25 ( 
.A(n_6),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_7),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_22),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_27),
.Y(n_40)
);

INVx2_ASAP7_75t_L g28 ( 
.A(n_22),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_28),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g29 ( 
.A(n_24),
.B(n_0),
.Y(n_29)
);

NOR2xp33_ASAP7_75t_L g37 ( 
.A(n_29),
.B(n_31),
.Y(n_37)
);

INVx8_ASAP7_75t_L g30 ( 
.A(n_22),
.Y(n_30)
);

INVx6_ASAP7_75t_L g48 ( 
.A(n_30),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_L g31 ( 
.A(n_20),
.B(n_13),
.Y(n_31)
);

INVx2_ASAP7_75t_L g32 ( 
.A(n_22),
.Y(n_32)
);

INVx4_ASAP7_75t_L g39 ( 
.A(n_32),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_22),
.Y(n_33)
);

INVx2_ASAP7_75t_SL g46 ( 
.A(n_33),
.Y(n_46)
);

INVx8_ASAP7_75t_L g34 ( 
.A(n_22),
.Y(n_34)
);

INVx3_ASAP7_75t_L g42 ( 
.A(n_34),
.Y(n_42)
);

BUFx5_ASAP7_75t_L g35 ( 
.A(n_24),
.Y(n_35)
);

BUFx3_ASAP7_75t_L g45 ( 
.A(n_35),
.Y(n_45)
);

BUFx3_ASAP7_75t_L g36 ( 
.A(n_25),
.Y(n_36)
);

INVx2_ASAP7_75t_L g49 ( 
.A(n_36),
.Y(n_49)
);

INVx2_ASAP7_75t_L g38 ( 
.A(n_36),
.Y(n_38)
);

INVx4_ASAP7_75t_L g65 ( 
.A(n_38),
.Y(n_65)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_36),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_41),
.B(n_44),
.Y(n_67)
);

A2O1A1Ixp33_ASAP7_75t_L g44 ( 
.A1(n_31),
.A2(n_17),
.B(n_20),
.C(n_21),
.Y(n_44)
);

INVx2_ASAP7_75t_L g47 ( 
.A(n_36),
.Y(n_47)
);

INVx3_ASAP7_75t_L g61 ( 
.A(n_47),
.Y(n_61)
);

OAI22xp33_ASAP7_75t_SL g50 ( 
.A1(n_44),
.A2(n_32),
.B1(n_28),
.B2(n_31),
.Y(n_50)
);

AOI22xp33_ASAP7_75t_L g75 ( 
.A1(n_50),
.A2(n_46),
.B1(n_48),
.B2(n_47),
.Y(n_75)
);

INVx2_ASAP7_75t_L g51 ( 
.A(n_43),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g73 ( 
.A(n_51),
.Y(n_73)
);

INVx2_ASAP7_75t_L g52 ( 
.A(n_43),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g90 ( 
.A(n_52),
.Y(n_90)
);

OAI22xp5_ASAP7_75t_L g53 ( 
.A1(n_37),
.A2(n_28),
.B1(n_32),
.B2(n_16),
.Y(n_53)
);

OAI22xp5_ASAP7_75t_L g86 ( 
.A1(n_53),
.A2(n_54),
.B1(n_57),
.B2(n_59),
.Y(n_86)
);

OAI22xp5_ASAP7_75t_L g54 ( 
.A1(n_37),
.A2(n_16),
.B1(n_20),
.B2(n_15),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_L g55 ( 
.A(n_43),
.B(n_29),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_L g76 ( 
.A(n_55),
.B(n_63),
.Y(n_76)
);

AOI22xp5_ASAP7_75t_SL g56 ( 
.A1(n_39),
.A2(n_16),
.B1(n_15),
.B2(n_17),
.Y(n_56)
);

INVxp67_ASAP7_75t_L g85 ( 
.A(n_56),
.Y(n_85)
);

AOI22xp5_ASAP7_75t_L g57 ( 
.A1(n_39),
.A2(n_34),
.B1(n_30),
.B2(n_16),
.Y(n_57)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_40),
.Y(n_58)
);

INVx4_ASAP7_75t_L g82 ( 
.A(n_58),
.Y(n_82)
);

AOI22xp33_ASAP7_75t_SL g59 ( 
.A1(n_48),
.A2(n_16),
.B1(n_15),
.B2(n_30),
.Y(n_59)
);

BUFx3_ASAP7_75t_L g60 ( 
.A(n_45),
.Y(n_60)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_60),
.Y(n_83)
);

INVx3_ASAP7_75t_L g62 ( 
.A(n_49),
.Y(n_62)
);

INVx5_ASAP7_75t_L g70 ( 
.A(n_62),
.Y(n_70)
);

OAI22xp5_ASAP7_75t_L g63 ( 
.A1(n_46),
.A2(n_15),
.B1(n_30),
.B2(n_34),
.Y(n_63)
);

AOI22xp33_ASAP7_75t_SL g64 ( 
.A1(n_48),
.A2(n_34),
.B1(n_17),
.B2(n_26),
.Y(n_64)
);

AOI22xp5_ASAP7_75t_SL g79 ( 
.A1(n_64),
.A2(n_46),
.B1(n_49),
.B2(n_38),
.Y(n_79)
);

INVx6_ASAP7_75t_L g66 ( 
.A(n_40),
.Y(n_66)
);

BUFx10_ASAP7_75t_L g74 ( 
.A(n_66),
.Y(n_74)
);

INVx2_ASAP7_75t_L g68 ( 
.A(n_40),
.Y(n_68)
);

INVx3_ASAP7_75t_L g89 ( 
.A(n_68),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_41),
.B(n_14),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_69),
.B(n_26),
.Y(n_72)
);

CKINVDCx20_ASAP7_75t_R g71 ( 
.A(n_69),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_SL g91 ( 
.A(n_71),
.B(n_72),
.Y(n_91)
);

AOI22xp5_ASAP7_75t_L g96 ( 
.A1(n_75),
.A2(n_54),
.B1(n_63),
.B2(n_51),
.Y(n_96)
);

CKINVDCx20_ASAP7_75t_R g77 ( 
.A(n_57),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_L g98 ( 
.A(n_77),
.B(n_88),
.Y(n_98)
);

MAJIxp5_ASAP7_75t_L g78 ( 
.A(n_67),
.B(n_27),
.C(n_33),
.Y(n_78)
);

MAJIxp5_ASAP7_75t_L g110 ( 
.A(n_78),
.B(n_81),
.C(n_77),
.Y(n_110)
);

OAI22xp5_ASAP7_75t_SL g104 ( 
.A1(n_79),
.A2(n_59),
.B1(n_66),
.B2(n_58),
.Y(n_104)
);

NOR2x1_ASAP7_75t_L g80 ( 
.A(n_67),
.B(n_50),
.Y(n_80)
);

CKINVDCx14_ASAP7_75t_R g95 ( 
.A(n_80),
.Y(n_95)
);

MAJIxp5_ASAP7_75t_L g81 ( 
.A(n_53),
.B(n_33),
.C(n_27),
.Y(n_81)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_65),
.Y(n_84)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_84),
.Y(n_93)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_65),
.Y(n_87)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_87),
.Y(n_94)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_65),
.Y(n_88)
);

AOI22xp5_ASAP7_75t_SL g92 ( 
.A1(n_78),
.A2(n_64),
.B1(n_56),
.B2(n_52),
.Y(n_92)
);

OAI21xp5_ASAP7_75t_L g131 ( 
.A1(n_92),
.A2(n_97),
.B(n_106),
.Y(n_131)
);

AOI22xp33_ASAP7_75t_L g128 ( 
.A1(n_96),
.A2(n_95),
.B1(n_108),
.B2(n_106),
.Y(n_128)
);

AOI21xp5_ASAP7_75t_L g97 ( 
.A1(n_85),
.A2(n_55),
.B(n_57),
.Y(n_97)
);

INVx2_ASAP7_75t_L g99 ( 
.A(n_73),
.Y(n_99)
);

INVx2_ASAP7_75t_L g123 ( 
.A(n_99),
.Y(n_123)
);

INVx2_ASAP7_75t_L g100 ( 
.A(n_73),
.Y(n_100)
);

AOI22xp33_ASAP7_75t_SL g119 ( 
.A1(n_100),
.A2(n_101),
.B1(n_99),
.B2(n_70),
.Y(n_119)
);

INVx8_ASAP7_75t_L g101 ( 
.A(n_89),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_L g102 ( 
.A(n_76),
.B(n_56),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_L g126 ( 
.A(n_102),
.B(n_107),
.Y(n_126)
);

BUFx6f_ASAP7_75t_L g103 ( 
.A(n_73),
.Y(n_103)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_103),
.Y(n_113)
);

AOI22xp5_ASAP7_75t_L g125 ( 
.A1(n_104),
.A2(n_83),
.B1(n_87),
.B2(n_84),
.Y(n_125)
);

INVxp67_ASAP7_75t_L g105 ( 
.A(n_79),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_SL g112 ( 
.A(n_105),
.B(n_109),
.Y(n_112)
);

AND2x2_ASAP7_75t_L g106 ( 
.A(n_86),
.B(n_33),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_L g107 ( 
.A(n_76),
.B(n_27),
.Y(n_107)
);

AOI22xp5_ASAP7_75t_L g108 ( 
.A1(n_86),
.A2(n_68),
.B1(n_66),
.B2(n_62),
.Y(n_108)
);

OAI22xp5_ASAP7_75t_SL g127 ( 
.A1(n_108),
.A2(n_70),
.B1(n_82),
.B2(n_62),
.Y(n_127)
);

INVxp67_ASAP7_75t_L g109 ( 
.A(n_81),
.Y(n_109)
);

XNOR2xp5_ASAP7_75t_L g116 ( 
.A(n_110),
.B(n_80),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_SL g111 ( 
.A(n_91),
.B(n_71),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_L g152 ( 
.A(n_111),
.B(n_114),
.Y(n_152)
);

CKINVDCx16_ASAP7_75t_R g114 ( 
.A(n_98),
.Y(n_114)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_98),
.Y(n_115)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_115),
.Y(n_160)
);

MAJIxp5_ASAP7_75t_L g138 ( 
.A(n_116),
.B(n_110),
.C(n_92),
.Y(n_138)
);

CKINVDCx20_ASAP7_75t_R g117 ( 
.A(n_93),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_L g158 ( 
.A(n_117),
.B(n_120),
.Y(n_158)
);

OAI22xp5_ASAP7_75t_L g118 ( 
.A1(n_97),
.A2(n_85),
.B1(n_80),
.B2(n_88),
.Y(n_118)
);

AOI22xp5_ASAP7_75t_L g147 ( 
.A1(n_118),
.A2(n_127),
.B1(n_128),
.B2(n_130),
.Y(n_147)
);

INVxp67_ASAP7_75t_L g159 ( 
.A(n_119),
.Y(n_159)
);

CKINVDCx20_ASAP7_75t_R g120 ( 
.A(n_93),
.Y(n_120)
);

CKINVDCx20_ASAP7_75t_R g121 ( 
.A(n_94),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_L g141 ( 
.A(n_121),
.B(n_122),
.Y(n_141)
);

CKINVDCx20_ASAP7_75t_R g122 ( 
.A(n_94),
.Y(n_122)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_107),
.Y(n_124)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_124),
.Y(n_135)
);

OAI22xp5_ASAP7_75t_SL g139 ( 
.A1(n_125),
.A2(n_133),
.B1(n_96),
.B2(n_92),
.Y(n_139)
);

CKINVDCx20_ASAP7_75t_R g129 ( 
.A(n_91),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_L g137 ( 
.A(n_129),
.B(n_134),
.Y(n_137)
);

OAI22xp5_ASAP7_75t_SL g130 ( 
.A1(n_95),
.A2(n_82),
.B1(n_61),
.B2(n_89),
.Y(n_130)
);

AOI22xp5_ASAP7_75t_SL g132 ( 
.A1(n_110),
.A2(n_83),
.B1(n_61),
.B2(n_42),
.Y(n_132)
);

OAI21xp5_ASAP7_75t_L g142 ( 
.A1(n_132),
.A2(n_106),
.B(n_104),
.Y(n_142)
);

AOI22xp5_ASAP7_75t_L g133 ( 
.A1(n_106),
.A2(n_61),
.B1(n_42),
.B2(n_74),
.Y(n_133)
);

OAI22xp5_ASAP7_75t_SL g134 ( 
.A1(n_102),
.A2(n_74),
.B1(n_21),
.B2(n_19),
.Y(n_134)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_115),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_L g176 ( 
.A(n_136),
.B(n_143),
.Y(n_176)
);

MAJIxp5_ASAP7_75t_L g163 ( 
.A(n_138),
.B(n_154),
.C(n_131),
.Y(n_163)
);

AOI22xp5_ASAP7_75t_L g165 ( 
.A1(n_139),
.A2(n_153),
.B1(n_127),
.B2(n_126),
.Y(n_165)
);

HB1xp67_ASAP7_75t_L g140 ( 
.A(n_132),
.Y(n_140)
);

CKINVDCx20_ASAP7_75t_R g161 ( 
.A(n_140),
.Y(n_161)
);

AOI22xp5_ASAP7_75t_SL g173 ( 
.A1(n_142),
.A2(n_155),
.B1(n_157),
.B2(n_18),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_L g143 ( 
.A(n_114),
.B(n_101),
.Y(n_143)
);

CKINVDCx16_ASAP7_75t_R g144 ( 
.A(n_111),
.Y(n_144)
);

NOR2xp33_ASAP7_75t_L g166 ( 
.A(n_144),
.B(n_149),
.Y(n_166)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_130),
.Y(n_145)
);

CKINVDCx20_ASAP7_75t_R g164 ( 
.A(n_145),
.Y(n_164)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_113),
.Y(n_146)
);

CKINVDCx20_ASAP7_75t_R g167 ( 
.A(n_146),
.Y(n_167)
);

AOI22xp33_ASAP7_75t_SL g148 ( 
.A1(n_129),
.A2(n_101),
.B1(n_100),
.B2(n_60),
.Y(n_148)
);

OAI22xp5_ASAP7_75t_SL g174 ( 
.A1(n_148),
.A2(n_45),
.B1(n_90),
.B2(n_35),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_L g149 ( 
.A(n_126),
.B(n_90),
.Y(n_149)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_113),
.Y(n_150)
);

CKINVDCx20_ASAP7_75t_R g177 ( 
.A(n_150),
.Y(n_177)
);

INVx2_ASAP7_75t_L g151 ( 
.A(n_123),
.Y(n_151)
);

CKINVDCx20_ASAP7_75t_R g182 ( 
.A(n_151),
.Y(n_182)
);

OAI22xp5_ASAP7_75t_SL g153 ( 
.A1(n_131),
.A2(n_74),
.B1(n_103),
.B2(n_90),
.Y(n_153)
);

MAJIxp5_ASAP7_75t_L g154 ( 
.A(n_116),
.B(n_118),
.C(n_112),
.Y(n_154)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_124),
.Y(n_155)
);

OAI21xp5_ASAP7_75t_SL g156 ( 
.A1(n_125),
.A2(n_60),
.B(n_18),
.Y(n_156)
);

OAI21xp5_ASAP7_75t_L g162 ( 
.A1(n_156),
.A2(n_121),
.B(n_122),
.Y(n_162)
);

CKINVDCx20_ASAP7_75t_R g157 ( 
.A(n_117),
.Y(n_157)
);

MAJIxp5_ASAP7_75t_SL g202 ( 
.A(n_162),
.B(n_170),
.C(n_174),
.Y(n_202)
);

XNOR2xp5_ASAP7_75t_L g187 ( 
.A(n_163),
.B(n_171),
.Y(n_187)
);

OAI22xp5_ASAP7_75t_SL g207 ( 
.A1(n_165),
.A2(n_168),
.B1(n_169),
.B2(n_179),
.Y(n_207)
);

AOI22xp5_ASAP7_75t_L g168 ( 
.A1(n_139),
.A2(n_120),
.B1(n_134),
.B2(n_133),
.Y(n_168)
);

AOI22xp5_ASAP7_75t_L g169 ( 
.A1(n_153),
.A2(n_123),
.B1(n_103),
.B2(n_74),
.Y(n_169)
);

OAI21xp33_ASAP7_75t_SL g170 ( 
.A1(n_144),
.A2(n_147),
.B(n_137),
.Y(n_170)
);

XOR2xp5_ASAP7_75t_L g171 ( 
.A(n_138),
.B(n_35),
.Y(n_171)
);

OAI22xp5_ASAP7_75t_L g172 ( 
.A1(n_159),
.A2(n_14),
.B1(n_26),
.B2(n_23),
.Y(n_172)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_172),
.Y(n_191)
);

OAI21xp5_ASAP7_75t_L g200 ( 
.A1(n_173),
.A2(n_135),
.B(n_150),
.Y(n_200)
);

XNOR2xp5_ASAP7_75t_L g175 ( 
.A(n_154),
.B(n_24),
.Y(n_175)
);

XNOR2xp5_ASAP7_75t_L g190 ( 
.A(n_175),
.B(n_180),
.Y(n_190)
);

NAND2xp33_ASAP7_75t_SL g178 ( 
.A(n_157),
.B(n_22),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_SL g196 ( 
.A(n_178),
.B(n_181),
.Y(n_196)
);

AOI22xp5_ASAP7_75t_L g179 ( 
.A1(n_145),
.A2(n_160),
.B1(n_136),
.B2(n_147),
.Y(n_179)
);

XNOR2xp5_ASAP7_75t_L g180 ( 
.A(n_142),
.B(n_24),
.Y(n_180)
);

XNOR2xp5_ASAP7_75t_SL g181 ( 
.A(n_152),
.B(n_24),
.Y(n_181)
);

XNOR2xp5_ASAP7_75t_L g183 ( 
.A(n_152),
.B(n_24),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_SL g203 ( 
.A(n_183),
.B(n_184),
.Y(n_203)
);

XNOR2xp5_ASAP7_75t_SL g184 ( 
.A(n_137),
.B(n_24),
.Y(n_184)
);

XNOR2xp5_ASAP7_75t_L g185 ( 
.A(n_160),
.B(n_13),
.Y(n_185)
);

NOR2xp33_ASAP7_75t_L g204 ( 
.A(n_185),
.B(n_25),
.Y(n_204)
);

INVx2_ASAP7_75t_SL g186 ( 
.A(n_167),
.Y(n_186)
);

INVx1_ASAP7_75t_SL g209 ( 
.A(n_186),
.Y(n_209)
);

CKINVDCx16_ASAP7_75t_R g188 ( 
.A(n_166),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_L g208 ( 
.A(n_188),
.B(n_192),
.Y(n_208)
);

NAND2xp5_ASAP7_75t_L g189 ( 
.A(n_177),
.B(n_158),
.Y(n_189)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_189),
.Y(n_218)
);

OAI22xp5_ASAP7_75t_L g192 ( 
.A1(n_168),
.A2(n_161),
.B1(n_162),
.B2(n_164),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_L g193 ( 
.A(n_176),
.B(n_158),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_L g213 ( 
.A(n_193),
.B(n_198),
.Y(n_213)
);

OAI21xp5_ASAP7_75t_SL g194 ( 
.A1(n_179),
.A2(n_141),
.B(n_156),
.Y(n_194)
);

OAI21xp5_ASAP7_75t_SL g225 ( 
.A1(n_194),
.A2(n_195),
.B(n_197),
.Y(n_225)
);

OAI21xp5_ASAP7_75t_SL g195 ( 
.A1(n_173),
.A2(n_143),
.B(n_155),
.Y(n_195)
);

AOI21xp5_ASAP7_75t_L g197 ( 
.A1(n_169),
.A2(n_135),
.B(n_149),
.Y(n_197)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_181),
.Y(n_198)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_184),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_L g226 ( 
.A(n_199),
.B(n_201),
.Y(n_226)
);

OAI22xp5_ASAP7_75t_L g210 ( 
.A1(n_200),
.A2(n_183),
.B1(n_185),
.B2(n_23),
.Y(n_210)
);

OAI22xp5_ASAP7_75t_L g201 ( 
.A1(n_163),
.A2(n_146),
.B1(n_151),
.B2(n_23),
.Y(n_201)
);

XNOR2xp5_ASAP7_75t_L g219 ( 
.A(n_204),
.B(n_206),
.Y(n_219)
);

INVx1_ASAP7_75t_SL g205 ( 
.A(n_182),
.Y(n_205)
);

CKINVDCx16_ASAP7_75t_R g224 ( 
.A(n_205),
.Y(n_224)
);

OAI21xp5_ASAP7_75t_SL g206 ( 
.A1(n_180),
.A2(n_21),
.B(n_19),
.Y(n_206)
);

AOI22xp5_ASAP7_75t_L g239 ( 
.A1(n_210),
.A2(n_215),
.B1(n_223),
.B2(n_4),
.Y(n_239)
);

MAJIxp5_ASAP7_75t_L g211 ( 
.A(n_187),
.B(n_171),
.C(n_175),
.Y(n_211)
);

MAJIxp5_ASAP7_75t_L g234 ( 
.A(n_211),
.B(n_214),
.C(n_217),
.Y(n_234)
);

NOR2xp33_ASAP7_75t_SL g212 ( 
.A(n_193),
.B(n_14),
.Y(n_212)
);

NAND2xp5_ASAP7_75t_L g240 ( 
.A(n_212),
.B(n_209),
.Y(n_240)
);

MAJIxp5_ASAP7_75t_L g214 ( 
.A(n_187),
.B(n_19),
.C(n_18),
.Y(n_214)
);

OAI22xp5_ASAP7_75t_SL g215 ( 
.A1(n_197),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_215)
);

AOI21xp33_ASAP7_75t_L g216 ( 
.A1(n_189),
.A2(n_0),
.B(n_1),
.Y(n_216)
);

OAI21xp5_ASAP7_75t_SL g230 ( 
.A1(n_216),
.A2(n_205),
.B(n_206),
.Y(n_230)
);

MAJIxp5_ASAP7_75t_L g217 ( 
.A(n_190),
.B(n_13),
.C(n_25),
.Y(n_217)
);

MAJIxp5_ASAP7_75t_L g220 ( 
.A(n_190),
.B(n_13),
.C(n_25),
.Y(n_220)
);

MAJIxp5_ASAP7_75t_L g242 ( 
.A(n_220),
.B(n_221),
.C(n_222),
.Y(n_242)
);

MAJIxp5_ASAP7_75t_L g221 ( 
.A(n_194),
.B(n_195),
.C(n_203),
.Y(n_221)
);

MAJIxp5_ASAP7_75t_L g222 ( 
.A(n_200),
.B(n_25),
.C(n_1),
.Y(n_222)
);

OAI22xp5_ASAP7_75t_L g223 ( 
.A1(n_191),
.A2(n_0),
.B1(n_2),
.B2(n_3),
.Y(n_223)
);

OAI21xp5_ASAP7_75t_L g227 ( 
.A1(n_225),
.A2(n_202),
.B(n_196),
.Y(n_227)
);

AOI21xp5_ASAP7_75t_L g248 ( 
.A1(n_227),
.A2(n_232),
.B(n_236),
.Y(n_248)
);

XNOR2xp5_ASAP7_75t_SL g228 ( 
.A(n_221),
.B(n_211),
.Y(n_228)
);

XOR2xp5_ASAP7_75t_L g250 ( 
.A(n_228),
.B(n_233),
.Y(n_250)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_218),
.Y(n_229)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_229),
.Y(n_245)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_230),
.Y(n_253)
);

AOI21xp5_ASAP7_75t_L g231 ( 
.A1(n_208),
.A2(n_202),
.B(n_186),
.Y(n_231)
);

OAI21xp5_ASAP7_75t_SL g246 ( 
.A1(n_231),
.A2(n_238),
.B(n_222),
.Y(n_246)
);

NOR2xp33_ASAP7_75t_L g232 ( 
.A(n_224),
.B(n_186),
.Y(n_232)
);

XOR2xp5_ASAP7_75t_L g233 ( 
.A(n_213),
.B(n_207),
.Y(n_233)
);

XOR2xp5_ASAP7_75t_L g235 ( 
.A(n_225),
.B(n_207),
.Y(n_235)
);

XOR2xp5_ASAP7_75t_L g252 ( 
.A(n_235),
.B(n_237),
.Y(n_252)
);

NAND2xp5_ASAP7_75t_SL g236 ( 
.A(n_226),
.B(n_3),
.Y(n_236)
);

XNOR2xp5_ASAP7_75t_SL g237 ( 
.A(n_219),
.B(n_11),
.Y(n_237)
);

OAI21xp5_ASAP7_75t_SL g238 ( 
.A1(n_209),
.A2(n_3),
.B(n_4),
.Y(n_238)
);

OAI22xp5_ASAP7_75t_SL g249 ( 
.A1(n_239),
.A2(n_220),
.B1(n_217),
.B2(n_215),
.Y(n_249)
);

HB1xp67_ASAP7_75t_L g244 ( 
.A(n_240),
.Y(n_244)
);

HB1xp67_ASAP7_75t_L g241 ( 
.A(n_214),
.Y(n_241)
);

XNOR2xp5_ASAP7_75t_L g243 ( 
.A(n_241),
.B(n_219),
.Y(n_243)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_243),
.Y(n_260)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_246),
.Y(n_263)
);

INVxp33_ASAP7_75t_L g247 ( 
.A(n_227),
.Y(n_247)
);

NOR2xp33_ASAP7_75t_L g262 ( 
.A(n_247),
.B(n_249),
.Y(n_262)
);

FAx1_ASAP7_75t_SL g251 ( 
.A(n_235),
.B(n_4),
.CI(n_5),
.CON(n_251),
.SN(n_251)
);

NAND2xp5_ASAP7_75t_SL g258 ( 
.A(n_251),
.B(n_234),
.Y(n_258)
);

MAJIxp5_ASAP7_75t_L g254 ( 
.A(n_242),
.B(n_5),
.C(n_6),
.Y(n_254)
);

MAJIxp5_ASAP7_75t_L g265 ( 
.A(n_254),
.B(n_255),
.C(n_5),
.Y(n_265)
);

MAJIxp5_ASAP7_75t_L g255 ( 
.A(n_242),
.B(n_5),
.C(n_6),
.Y(n_255)
);

BUFx6f_ASAP7_75t_L g256 ( 
.A(n_247),
.Y(n_256)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_256),
.Y(n_270)
);

XOR2xp5_ASAP7_75t_L g257 ( 
.A(n_250),
.B(n_228),
.Y(n_257)
);

MAJIxp5_ASAP7_75t_L g273 ( 
.A(n_257),
.B(n_264),
.C(n_266),
.Y(n_273)
);

NOR2xp33_ASAP7_75t_L g268 ( 
.A(n_258),
.B(n_259),
.Y(n_268)
);

NAND2xp5_ASAP7_75t_SL g259 ( 
.A(n_248),
.B(n_233),
.Y(n_259)
);

OAI22xp5_ASAP7_75t_SL g261 ( 
.A1(n_253),
.A2(n_234),
.B1(n_237),
.B2(n_7),
.Y(n_261)
);

NOR2xp33_ASAP7_75t_L g271 ( 
.A(n_261),
.B(n_265),
.Y(n_271)
);

XOR2xp5_ASAP7_75t_L g264 ( 
.A(n_250),
.B(n_11),
.Y(n_264)
);

OAI22xp5_ASAP7_75t_SL g266 ( 
.A1(n_251),
.A2(n_252),
.B1(n_245),
.B2(n_255),
.Y(n_266)
);

XNOR2xp5_ASAP7_75t_SL g267 ( 
.A(n_257),
.B(n_243),
.Y(n_267)
);

AOI22xp5_ASAP7_75t_SL g277 ( 
.A1(n_267),
.A2(n_264),
.B1(n_266),
.B2(n_265),
.Y(n_277)
);

NOR2x1_ASAP7_75t_L g269 ( 
.A(n_256),
.B(n_244),
.Y(n_269)
);

NAND2xp5_ASAP7_75t_SL g280 ( 
.A(n_269),
.B(n_7),
.Y(n_280)
);

BUFx4f_ASAP7_75t_SL g272 ( 
.A(n_262),
.Y(n_272)
);

NAND2xp5_ASAP7_75t_L g276 ( 
.A(n_272),
.B(n_275),
.Y(n_276)
);

NOR2xp67_ASAP7_75t_L g274 ( 
.A(n_263),
.B(n_251),
.Y(n_274)
);

OAI22xp5_ASAP7_75t_SL g281 ( 
.A1(n_274),
.A2(n_11),
.B1(n_8),
.B2(n_9),
.Y(n_281)
);

OAI21xp5_ASAP7_75t_L g275 ( 
.A1(n_260),
.A2(n_254),
.B(n_252),
.Y(n_275)
);

XNOR2xp5_ASAP7_75t_L g283 ( 
.A(n_277),
.B(n_279),
.Y(n_283)
);

INVxp67_ASAP7_75t_L g278 ( 
.A(n_268),
.Y(n_278)
);

OAI21xp5_ASAP7_75t_L g282 ( 
.A1(n_278),
.A2(n_280),
.B(n_271),
.Y(n_282)
);

NAND2xp5_ASAP7_75t_L g279 ( 
.A(n_270),
.B(n_6),
.Y(n_279)
);

AOI21x1_ASAP7_75t_L g284 ( 
.A1(n_281),
.A2(n_274),
.B(n_272),
.Y(n_284)
);

MAJIxp5_ASAP7_75t_L g286 ( 
.A(n_282),
.B(n_284),
.C(n_273),
.Y(n_286)
);

OAI21xp5_ASAP7_75t_SL g285 ( 
.A1(n_283),
.A2(n_276),
.B(n_278),
.Y(n_285)
);

OAI21xp5_ASAP7_75t_SL g287 ( 
.A1(n_285),
.A2(n_286),
.B(n_7),
.Y(n_287)
);

XOR2xp5_ASAP7_75t_L g288 ( 
.A(n_287),
.B(n_10),
.Y(n_288)
);

AOI21xp5_ASAP7_75t_L g289 ( 
.A1(n_288),
.A2(n_8),
.B(n_9),
.Y(n_289)
);

OAI21xp5_ASAP7_75t_L g290 ( 
.A1(n_289),
.A2(n_8),
.B(n_9),
.Y(n_290)
);

AND2x2_ASAP7_75t_L g291 ( 
.A(n_290),
.B(n_10),
.Y(n_291)
);

XNOR2xp5_ASAP7_75t_L g292 ( 
.A(n_291),
.B(n_10),
.Y(n_292)
);


endmodule