module fake_jpeg_2931_n_680 (n_13, n_1, n_10, n_6, n_14, n_19, n_18, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_680);

input n_13;
input n_1;
input n_10;
input n_6;
input n_14;
input n_19;
input n_18;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_680;

wire n_529;
wire n_595;
wire n_390;
wire n_552;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_252;
wire n_525;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_586;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_657;
wire n_27;
wire n_664;
wire n_365;
wire n_179;
wire n_620;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_678;
wire n_611;
wire n_44;
wire n_355;
wire n_519;
wire n_276;
wire n_143;
wire n_431;
wire n_102;
wire n_549;
wire n_196;
wire n_66;
wire n_374;
wire n_566;
wire n_142;
wire n_417;
wire n_362;
wire n_470;
wire n_597;
wire n_172;
wire n_547;
wire n_345;
wire n_591;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_513;
wire n_283;
wire n_107;
wire n_490;
wire n_635;
wire n_517;
wire n_629;
wire n_415;
wire n_479;
wire n_543;
wire n_357;
wire n_89;
wire n_131;
wire n_607;
wire n_294;
wire n_230;
wire n_643;
wire n_170;
wire n_602;
wire n_313;
wire n_542;
wire n_574;
wire n_264;
wire n_647;
wire n_437;
wire n_93;
wire n_227;
wire n_559;
wire n_641;
wire n_48;
wire n_465;
wire n_638;
wire n_200;
wire n_582;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_623;
wire n_579;
wire n_416;
wire n_221;
wire n_256;
wire n_454;
wire n_540;
wire n_292;
wire n_213;
wire n_135;
wire n_435;
wire n_189;
wire n_637;
wire n_370;
wire n_410;
wire n_571;
wire n_82;
wire n_155;
wire n_508;
wire n_672;
wire n_309;
wire n_624;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_606;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_596;
wire n_569;
wire n_400;
wire n_646;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_544;
wire n_31;
wire n_277;
wire n_663;
wire n_255;
wire n_605;
wire n_601;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_393;
wire n_349;
wire n_234;
wire n_530;
wire n_634;
wire n_23;
wire n_69;
wire n_658;
wire n_195;
wire n_450;
wire n_557;
wire n_408;
wire n_80;
wire n_562;
wire n_204;
wire n_666;
wire n_639;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_645;
wire n_298;
wire n_106;
wire n_545;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_584;
wire n_254;
wire n_608;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_622;
wire n_463;
wire n_667;
wire n_92;
wire n_332;
wire n_640;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_653;
wire n_474;
wire n_539;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_626;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_668;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_575;
wire n_268;
wire n_404;
wire n_91;
wire n_511;
wire n_486;
wire n_305;
wire n_161;
wire n_441;
wire n_555;
wire n_342;
wire n_642;
wire n_101;
wire n_226;
wire n_509;
wire n_644;
wire n_149;
wire n_87;
wire n_46;
wire n_578;
wire n_656;
wire n_589;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_614;
wire n_97;
wire n_649;
wire n_573;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_610;
wire n_174;
wire n_198;
wire n_422;
wire n_560;
wire n_190;
wire n_510;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_536;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_679;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_537;
wire n_110;
wire n_594;
wire n_590;
wire n_531;
wire n_76;
wire n_278;
wire n_343;
wire n_577;
wire n_26;
wire n_88;
wire n_397;
wire n_592;
wire n_363;
wire n_570;
wire n_238;
wire n_598;
wire n_615;
wire n_29;
wire n_103;
wire n_150;
wire n_352;
wire n_350;
wire n_488;
wire n_662;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_554;
wire n_301;
wire n_609;
wire n_201;
wire n_420;
wire n_676;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_648;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_523;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_533;
wire n_612;
wire n_296;
wire n_384;
wire n_588;
wire n_168;
wire n_670;
wire n_459;
wire n_274;
wire n_485;
wire n_585;
wire n_491;
wire n_24;
wire n_526;
wire n_467;
wire n_269;
wire n_572;
wire n_546;
wire n_287;
wire n_219;
wire n_452;
wire n_631;
wire n_433;
wire n_636;
wire n_77;
wire n_473;
wire n_45;
wire n_520;
wire n_476;
wire n_337;
wire n_317;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_344;
wire n_328;
wire n_650;
wire n_218;
wire n_63;
wire n_652;
wire n_599;
wire n_239;
wire n_674;
wire n_243;
wire n_481;
wire n_628;
wire n_619;
wire n_348;
wire n_587;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_583;
wire n_522;
wire n_333;
wire n_518;
wire n_132;
wire n_133;
wire n_419;
wire n_378;
wire n_565;
wire n_302;
wire n_216;
wire n_528;
wire n_184;
wire n_655;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_260;
wire n_199;
wire n_550;
wire n_413;
wire n_275;
wire n_494;
wire n_604;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_551;
wire n_36;
wire n_62;
wire n_600;
wire n_492;
wire n_603;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_567;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_515;
wire n_347;
wire n_521;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_538;
wire n_625;
wire n_147;
wire n_449;
wire n_627;
wire n_98;
wire n_251;
wire n_534;
wire n_472;
wire n_279;
wire n_593;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_618;
wire n_356;
wire n_119;
wire n_484;
wire n_568;
wire n_83;
wire n_395;
wire n_659;
wire n_125;
wire n_661;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_576;
wire n_469;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_553;
wire n_257;
wire n_61;
wire n_173;
wire n_561;
wire n_244;
wire n_232;
wire n_527;
wire n_482;
wire n_673;
wire n_58;
wire n_41;
wire n_613;
wire n_630;
wire n_266;
wire n_548;
wire n_665;
wire n_72;
wire n_512;
wire n_654;
wire n_445;
wire n_443;
wire n_677;
wire n_617;
wire n_215;
wire n_212;
wire n_516;
wire n_183;
wire n_409;
wire n_532;
wire n_249;
wire n_412;
wire n_581;
wire n_217;
wire n_471;
wire n_580;
wire n_541;
wire n_53;
wire n_372;
wire n_558;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_535;
wire n_671;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_556;
wire n_669;
wire n_524;
wire n_402;
wire n_563;
wire n_504;
wire n_438;
wire n_475;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_660;
wire n_373;
wire n_633;
wire n_112;
wire n_632;
wire n_616;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_514;
wire n_651;
wire n_564;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_675;
wire n_335;
wire n_120;
wire n_621;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_8),
.Y(n_20)
);

INVx2_ASAP7_75t_L g21 ( 
.A(n_17),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_4),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_14),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_19),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_19),
.Y(n_25)
);

NOR2xp33_ASAP7_75t_L g26 ( 
.A(n_17),
.B(n_3),
.Y(n_26)
);

INVx8_ASAP7_75t_L g27 ( 
.A(n_17),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_18),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_11),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_5),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_13),
.Y(n_31)
);

BUFx12f_ASAP7_75t_L g32 ( 
.A(n_0),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_17),
.Y(n_33)
);

INVxp67_ASAP7_75t_L g34 ( 
.A(n_7),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_5),
.Y(n_35)
);

BUFx3_ASAP7_75t_L g36 ( 
.A(n_0),
.Y(n_36)
);

BUFx5_ASAP7_75t_L g37 ( 
.A(n_13),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_13),
.Y(n_38)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_5),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_11),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_19),
.Y(n_41)
);

BUFx12f_ASAP7_75t_L g42 ( 
.A(n_8),
.Y(n_42)
);

INVx6_ASAP7_75t_L g43 ( 
.A(n_13),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_SL g44 ( 
.A(n_5),
.B(n_7),
.Y(n_44)
);

INVx13_ASAP7_75t_L g45 ( 
.A(n_7),
.Y(n_45)
);

INVx3_ASAP7_75t_L g46 ( 
.A(n_14),
.Y(n_46)
);

BUFx12_ASAP7_75t_L g47 ( 
.A(n_14),
.Y(n_47)
);

BUFx4f_ASAP7_75t_L g48 ( 
.A(n_1),
.Y(n_48)
);

INVx11_ASAP7_75t_L g49 ( 
.A(n_1),
.Y(n_49)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_15),
.Y(n_50)
);

INVx5_ASAP7_75t_L g51 ( 
.A(n_6),
.Y(n_51)
);

BUFx12_ASAP7_75t_L g52 ( 
.A(n_9),
.Y(n_52)
);

BUFx3_ASAP7_75t_L g53 ( 
.A(n_12),
.Y(n_53)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_4),
.Y(n_54)
);

BUFx3_ASAP7_75t_L g55 ( 
.A(n_6),
.Y(n_55)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_18),
.Y(n_56)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_1),
.Y(n_57)
);

CKINVDCx20_ASAP7_75t_R g58 ( 
.A(n_0),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_44),
.B(n_18),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g161 ( 
.A(n_59),
.B(n_71),
.Y(n_161)
);

INVx8_ASAP7_75t_L g60 ( 
.A(n_32),
.Y(n_60)
);

BUFx2_ASAP7_75t_L g160 ( 
.A(n_60),
.Y(n_160)
);

BUFx4f_ASAP7_75t_L g61 ( 
.A(n_21),
.Y(n_61)
);

INVx1_ASAP7_75t_SL g224 ( 
.A(n_61),
.Y(n_224)
);

BUFx12f_ASAP7_75t_L g62 ( 
.A(n_47),
.Y(n_62)
);

BUFx4f_ASAP7_75t_SL g137 ( 
.A(n_62),
.Y(n_137)
);

INVx3_ASAP7_75t_L g63 ( 
.A(n_51),
.Y(n_63)
);

INVx3_ASAP7_75t_L g139 ( 
.A(n_63),
.Y(n_139)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_23),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g148 ( 
.A(n_64),
.Y(n_148)
);

BUFx3_ASAP7_75t_L g65 ( 
.A(n_51),
.Y(n_65)
);

BUFx2_ASAP7_75t_L g177 ( 
.A(n_65),
.Y(n_177)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_23),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g184 ( 
.A(n_66),
.Y(n_184)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_23),
.Y(n_67)
);

BUFx6f_ASAP7_75t_L g186 ( 
.A(n_67),
.Y(n_186)
);

INVx4_ASAP7_75t_SL g68 ( 
.A(n_32),
.Y(n_68)
);

BUFx3_ASAP7_75t_L g165 ( 
.A(n_68),
.Y(n_165)
);

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_31),
.Y(n_69)
);

BUFx6f_ASAP7_75t_L g188 ( 
.A(n_69),
.Y(n_188)
);

INVx3_ASAP7_75t_SL g70 ( 
.A(n_27),
.Y(n_70)
);

BUFx2_ASAP7_75t_L g193 ( 
.A(n_70),
.Y(n_193)
);

CKINVDCx20_ASAP7_75t_R g71 ( 
.A(n_24),
.Y(n_71)
);

INVx3_ASAP7_75t_L g72 ( 
.A(n_51),
.Y(n_72)
);

INVx3_ASAP7_75t_L g152 ( 
.A(n_72),
.Y(n_152)
);

INVx3_ASAP7_75t_L g73 ( 
.A(n_36),
.Y(n_73)
);

INVx3_ASAP7_75t_L g179 ( 
.A(n_73),
.Y(n_179)
);

BUFx6f_ASAP7_75t_L g74 ( 
.A(n_31),
.Y(n_74)
);

BUFx6f_ASAP7_75t_L g196 ( 
.A(n_74),
.Y(n_196)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_28),
.Y(n_75)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_75),
.Y(n_144)
);

BUFx12f_ASAP7_75t_L g76 ( 
.A(n_47),
.Y(n_76)
);

BUFx4f_ASAP7_75t_SL g149 ( 
.A(n_76),
.Y(n_149)
);

INVx5_ASAP7_75t_L g77 ( 
.A(n_27),
.Y(n_77)
);

BUFx3_ASAP7_75t_L g181 ( 
.A(n_77),
.Y(n_181)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_28),
.Y(n_78)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_78),
.Y(n_150)
);

BUFx6f_ASAP7_75t_L g79 ( 
.A(n_31),
.Y(n_79)
);

BUFx6f_ASAP7_75t_L g199 ( 
.A(n_79),
.Y(n_199)
);

INVx6_ASAP7_75t_SL g80 ( 
.A(n_45),
.Y(n_80)
);

CKINVDCx9p33_ASAP7_75t_R g221 ( 
.A(n_80),
.Y(n_221)
);

INVx2_ASAP7_75t_L g81 ( 
.A(n_21),
.Y(n_81)
);

INVx2_ASAP7_75t_L g136 ( 
.A(n_81),
.Y(n_136)
);

INVx2_ASAP7_75t_R g82 ( 
.A(n_44),
.Y(n_82)
);

AND2x2_ASAP7_75t_L g167 ( 
.A(n_82),
.B(n_58),
.Y(n_167)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_26),
.B(n_0),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g169 ( 
.A(n_83),
.B(n_89),
.Y(n_169)
);

BUFx6f_ASAP7_75t_L g84 ( 
.A(n_40),
.Y(n_84)
);

BUFx6f_ASAP7_75t_L g231 ( 
.A(n_84),
.Y(n_231)
);

BUFx6f_ASAP7_75t_L g85 ( 
.A(n_40),
.Y(n_85)
);

BUFx6f_ASAP7_75t_L g206 ( 
.A(n_85),
.Y(n_206)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_56),
.Y(n_86)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_86),
.Y(n_151)
);

INVx6_ASAP7_75t_L g87 ( 
.A(n_40),
.Y(n_87)
);

BUFx6f_ASAP7_75t_L g207 ( 
.A(n_87),
.Y(n_207)
);

BUFx6f_ASAP7_75t_L g88 ( 
.A(n_43),
.Y(n_88)
);

INVx6_ASAP7_75t_L g133 ( 
.A(n_88),
.Y(n_133)
);

CKINVDCx20_ASAP7_75t_R g89 ( 
.A(n_24),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_SL g90 ( 
.A(n_26),
.B(n_1),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g180 ( 
.A(n_90),
.B(n_92),
.Y(n_180)
);

BUFx3_ASAP7_75t_L g91 ( 
.A(n_36),
.Y(n_91)
);

BUFx3_ASAP7_75t_L g183 ( 
.A(n_91),
.Y(n_183)
);

CKINVDCx20_ASAP7_75t_R g92 ( 
.A(n_24),
.Y(n_92)
);

INVx4_ASAP7_75t_L g93 ( 
.A(n_37),
.Y(n_93)
);

INVx3_ASAP7_75t_L g194 ( 
.A(n_93),
.Y(n_194)
);

INVx5_ASAP7_75t_L g94 ( 
.A(n_27),
.Y(n_94)
);

INVx4_ASAP7_75t_L g166 ( 
.A(n_94),
.Y(n_166)
);

BUFx4f_ASAP7_75t_L g95 ( 
.A(n_45),
.Y(n_95)
);

INVx2_ASAP7_75t_L g230 ( 
.A(n_95),
.Y(n_230)
);

BUFx5_ASAP7_75t_L g96 ( 
.A(n_37),
.Y(n_96)
);

INVx4_ASAP7_75t_L g178 ( 
.A(n_96),
.Y(n_178)
);

INVx3_ASAP7_75t_L g97 ( 
.A(n_36),
.Y(n_97)
);

INVx4_ASAP7_75t_L g187 ( 
.A(n_97),
.Y(n_187)
);

INVx3_ASAP7_75t_L g98 ( 
.A(n_53),
.Y(n_98)
);

INVx4_ASAP7_75t_L g189 ( 
.A(n_98),
.Y(n_189)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_56),
.Y(n_99)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_99),
.Y(n_162)
);

INVx11_ASAP7_75t_L g100 ( 
.A(n_32),
.Y(n_100)
);

INVx11_ASAP7_75t_L g211 ( 
.A(n_100),
.Y(n_211)
);

INVx2_ASAP7_75t_L g101 ( 
.A(n_46),
.Y(n_101)
);

INVx2_ASAP7_75t_L g141 ( 
.A(n_101),
.Y(n_141)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_29),
.Y(n_102)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_102),
.Y(n_170)
);

BUFx12_ASAP7_75t_L g103 ( 
.A(n_34),
.Y(n_103)
);

BUFx12f_ASAP7_75t_L g140 ( 
.A(n_103),
.Y(n_140)
);

BUFx6f_ASAP7_75t_L g104 ( 
.A(n_43),
.Y(n_104)
);

INVx6_ASAP7_75t_L g135 ( 
.A(n_104),
.Y(n_135)
);

INVx8_ASAP7_75t_L g105 ( 
.A(n_32),
.Y(n_105)
);

INVx5_ASAP7_75t_L g138 ( 
.A(n_105),
.Y(n_138)
);

BUFx6f_ASAP7_75t_L g106 ( 
.A(n_43),
.Y(n_106)
);

INVx6_ASAP7_75t_L g164 ( 
.A(n_106),
.Y(n_164)
);

BUFx8_ASAP7_75t_L g107 ( 
.A(n_45),
.Y(n_107)
);

BUFx24_ASAP7_75t_L g220 ( 
.A(n_107),
.Y(n_220)
);

BUFx6f_ASAP7_75t_L g108 ( 
.A(n_25),
.Y(n_108)
);

INVx6_ASAP7_75t_L g174 ( 
.A(n_108),
.Y(n_174)
);

BUFx3_ASAP7_75t_L g109 ( 
.A(n_53),
.Y(n_109)
);

INVx5_ASAP7_75t_L g145 ( 
.A(n_109),
.Y(n_145)
);

CKINVDCx20_ASAP7_75t_R g110 ( 
.A(n_25),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_L g198 ( 
.A(n_110),
.B(n_111),
.Y(n_198)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_20),
.B(n_2),
.Y(n_111)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_29),
.Y(n_112)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_112),
.Y(n_185)
);

BUFx6f_ASAP7_75t_L g113 ( 
.A(n_25),
.Y(n_113)
);

INVx6_ASAP7_75t_L g215 ( 
.A(n_113),
.Y(n_215)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_30),
.Y(n_114)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_114),
.Y(n_202)
);

INVx3_ASAP7_75t_L g115 ( 
.A(n_53),
.Y(n_115)
);

INVx4_ASAP7_75t_L g201 ( 
.A(n_115),
.Y(n_201)
);

BUFx6f_ASAP7_75t_L g116 ( 
.A(n_41),
.Y(n_116)
);

INVx6_ASAP7_75t_L g218 ( 
.A(n_116),
.Y(n_218)
);

CKINVDCx20_ASAP7_75t_R g117 ( 
.A(n_41),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_L g214 ( 
.A(n_117),
.B(n_119),
.Y(n_214)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_30),
.Y(n_118)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_118),
.Y(n_212)
);

CKINVDCx20_ASAP7_75t_R g119 ( 
.A(n_41),
.Y(n_119)
);

INVx4_ASAP7_75t_L g120 ( 
.A(n_37),
.Y(n_120)
);

INVx4_ASAP7_75t_L g213 ( 
.A(n_120),
.Y(n_213)
);

INVx4_ASAP7_75t_L g121 ( 
.A(n_46),
.Y(n_121)
);

INVx4_ASAP7_75t_L g217 ( 
.A(n_121),
.Y(n_217)
);

NAND2xp5_ASAP7_75t_L g122 ( 
.A(n_20),
.B(n_16),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_L g226 ( 
.A(n_122),
.B(n_123),
.Y(n_226)
);

CKINVDCx20_ASAP7_75t_R g123 ( 
.A(n_48),
.Y(n_123)
);

BUFx6f_ASAP7_75t_L g124 ( 
.A(n_55),
.Y(n_124)
);

INVx5_ASAP7_75t_L g158 ( 
.A(n_124),
.Y(n_158)
);

NOR2xp33_ASAP7_75t_L g125 ( 
.A(n_22),
.B(n_2),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_SL g219 ( 
.A(n_125),
.B(n_58),
.Y(n_219)
);

INVx2_ASAP7_75t_L g126 ( 
.A(n_46),
.Y(n_126)
);

INVx2_ASAP7_75t_L g142 ( 
.A(n_126),
.Y(n_142)
);

INVx5_ASAP7_75t_L g127 ( 
.A(n_55),
.Y(n_127)
);

INVx4_ASAP7_75t_L g225 ( 
.A(n_127),
.Y(n_225)
);

INVx6_ASAP7_75t_L g128 ( 
.A(n_32),
.Y(n_128)
);

INVx2_ASAP7_75t_L g143 ( 
.A(n_128),
.Y(n_143)
);

BUFx3_ASAP7_75t_L g129 ( 
.A(n_55),
.Y(n_129)
);

INVx5_ASAP7_75t_L g176 ( 
.A(n_129),
.Y(n_176)
);

INVx8_ASAP7_75t_L g130 ( 
.A(n_42),
.Y(n_130)
);

INVx5_ASAP7_75t_L g203 ( 
.A(n_130),
.Y(n_203)
);

INVx3_ASAP7_75t_L g131 ( 
.A(n_42),
.Y(n_131)
);

BUFx12f_ASAP7_75t_L g147 ( 
.A(n_131),
.Y(n_147)
);

INVx4_ASAP7_75t_SL g132 ( 
.A(n_42),
.Y(n_132)
);

INVx13_ASAP7_75t_L g159 ( 
.A(n_132),
.Y(n_159)
);

BUFx12_ASAP7_75t_L g134 ( 
.A(n_107),
.Y(n_134)
);

INVx13_ASAP7_75t_L g313 ( 
.A(n_134),
.Y(n_313)
);

BUFx10_ASAP7_75t_L g146 ( 
.A(n_62),
.Y(n_146)
);

BUFx24_ASAP7_75t_L g295 ( 
.A(n_146),
.Y(n_295)
);

OAI22xp5_ASAP7_75t_SL g153 ( 
.A1(n_83),
.A2(n_48),
.B1(n_42),
.B2(n_22),
.Y(n_153)
);

AOI22xp5_ASAP7_75t_SL g281 ( 
.A1(n_153),
.A2(n_79),
.B1(n_52),
.B2(n_47),
.Y(n_281)
);

CKINVDCx20_ASAP7_75t_R g154 ( 
.A(n_128),
.Y(n_154)
);

NOR2xp33_ASAP7_75t_SL g254 ( 
.A(n_154),
.B(n_167),
.Y(n_254)
);

INVx2_ASAP7_75t_L g155 ( 
.A(n_61),
.Y(n_155)
);

INVx2_ASAP7_75t_L g248 ( 
.A(n_155),
.Y(n_248)
);

AOI22xp33_ASAP7_75t_SL g156 ( 
.A1(n_68),
.A2(n_49),
.B1(n_48),
.B2(n_42),
.Y(n_156)
);

AOI22xp33_ASAP7_75t_SL g263 ( 
.A1(n_156),
.A2(n_209),
.B1(n_91),
.B2(n_33),
.Y(n_263)
);

INVx2_ASAP7_75t_L g157 ( 
.A(n_95),
.Y(n_157)
);

INVx2_ASAP7_75t_L g262 ( 
.A(n_157),
.Y(n_262)
);

AOI22xp33_ASAP7_75t_L g163 ( 
.A1(n_64),
.A2(n_48),
.B1(n_49),
.B2(n_35),
.Y(n_163)
);

OAI22xp5_ASAP7_75t_SL g279 ( 
.A1(n_163),
.A2(n_171),
.B1(n_38),
.B2(n_33),
.Y(n_279)
);

INVx2_ASAP7_75t_L g168 ( 
.A(n_87),
.Y(n_168)
);

INVx2_ASAP7_75t_L g243 ( 
.A(n_168),
.Y(n_243)
);

AOI22xp33_ASAP7_75t_L g171 ( 
.A1(n_66),
.A2(n_49),
.B1(n_57),
.B2(n_35),
.Y(n_171)
);

INVx2_ASAP7_75t_L g172 ( 
.A(n_88),
.Y(n_172)
);

INVx2_ASAP7_75t_L g245 ( 
.A(n_172),
.Y(n_245)
);

INVx2_ASAP7_75t_L g173 ( 
.A(n_104),
.Y(n_173)
);

INVx2_ASAP7_75t_L g275 ( 
.A(n_173),
.Y(n_275)
);

BUFx5_ASAP7_75t_L g175 ( 
.A(n_103),
.Y(n_175)
);

INVx2_ASAP7_75t_SL g246 ( 
.A(n_175),
.Y(n_246)
);

CKINVDCx20_ASAP7_75t_R g182 ( 
.A(n_106),
.Y(n_182)
);

NOR2xp33_ASAP7_75t_SL g304 ( 
.A(n_182),
.B(n_205),
.Y(n_304)
);

BUFx12f_ASAP7_75t_L g190 ( 
.A(n_60),
.Y(n_190)
);

INVx5_ASAP7_75t_L g265 ( 
.A(n_190),
.Y(n_265)
);

BUFx12f_ASAP7_75t_L g191 ( 
.A(n_105),
.Y(n_191)
);

INVx8_ASAP7_75t_L g297 ( 
.A(n_191),
.Y(n_297)
);

BUFx12f_ASAP7_75t_L g192 ( 
.A(n_130),
.Y(n_192)
);

INVx8_ASAP7_75t_L g307 ( 
.A(n_192),
.Y(n_307)
);

CKINVDCx16_ASAP7_75t_R g195 ( 
.A(n_132),
.Y(n_195)
);

AND2x2_ASAP7_75t_L g238 ( 
.A(n_195),
.B(n_210),
.Y(n_238)
);

INVx2_ASAP7_75t_L g197 ( 
.A(n_108),
.Y(n_197)
);

INVx2_ASAP7_75t_L g285 ( 
.A(n_197),
.Y(n_285)
);

INVx2_ASAP7_75t_L g200 ( 
.A(n_113),
.Y(n_200)
);

INVx2_ASAP7_75t_L g289 ( 
.A(n_200),
.Y(n_289)
);

INVx2_ASAP7_75t_L g204 ( 
.A(n_116),
.Y(n_204)
);

INVx2_ASAP7_75t_L g290 ( 
.A(n_204),
.Y(n_290)
);

CKINVDCx20_ASAP7_75t_R g205 ( 
.A(n_124),
.Y(n_205)
);

INVx5_ASAP7_75t_L g208 ( 
.A(n_62),
.Y(n_208)
);

INVx4_ASAP7_75t_L g274 ( 
.A(n_208),
.Y(n_274)
);

AOI22xp33_ASAP7_75t_SL g209 ( 
.A1(n_93),
.A2(n_50),
.B1(n_57),
.B2(n_39),
.Y(n_209)
);

CKINVDCx16_ASAP7_75t_R g210 ( 
.A(n_70),
.Y(n_210)
);

INVx2_ASAP7_75t_L g216 ( 
.A(n_67),
.Y(n_216)
);

INVx2_ASAP7_75t_L g299 ( 
.A(n_216),
.Y(n_299)
);

NAND2xp5_ASAP7_75t_SL g241 ( 
.A(n_219),
.B(n_228),
.Y(n_241)
);

INVx2_ASAP7_75t_L g222 ( 
.A(n_69),
.Y(n_222)
);

INVx2_ASAP7_75t_L g300 ( 
.A(n_222),
.Y(n_300)
);

MAJIxp5_ASAP7_75t_L g223 ( 
.A(n_59),
.B(n_50),
.C(n_39),
.Y(n_223)
);

MAJIxp5_ASAP7_75t_L g303 ( 
.A(n_223),
.B(n_52),
.C(n_7),
.Y(n_303)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_111),
.Y(n_227)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_227),
.Y(n_233)
);

NAND2xp5_ASAP7_75t_SL g228 ( 
.A(n_82),
.B(n_54),
.Y(n_228)
);

INVx2_ASAP7_75t_L g229 ( 
.A(n_74),
.Y(n_229)
);

INVx2_ASAP7_75t_L g301 ( 
.A(n_229),
.Y(n_301)
);

CKINVDCx20_ASAP7_75t_R g232 ( 
.A(n_221),
.Y(n_232)
);

NAND2xp5_ASAP7_75t_SL g322 ( 
.A(n_232),
.B(n_240),
.Y(n_322)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_144),
.Y(n_234)
);

INVx1_ASAP7_75t_SL g370 ( 
.A(n_234),
.Y(n_370)
);

BUFx6f_ASAP7_75t_L g235 ( 
.A(n_148),
.Y(n_235)
);

INVx5_ASAP7_75t_L g323 ( 
.A(n_235),
.Y(n_323)
);

AOI21xp33_ASAP7_75t_L g236 ( 
.A1(n_226),
.A2(n_125),
.B(n_76),
.Y(n_236)
);

OAI21xp33_ASAP7_75t_L g330 ( 
.A1(n_236),
.A2(n_269),
.B(n_270),
.Y(n_330)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_150),
.Y(n_237)
);

HB1xp67_ASAP7_75t_L g339 ( 
.A(n_237),
.Y(n_339)
);

NOR2xp33_ASAP7_75t_L g239 ( 
.A(n_180),
.B(n_129),
.Y(n_239)
);

NOR2xp33_ASAP7_75t_SL g344 ( 
.A(n_239),
.B(n_250),
.Y(n_344)
);

CKINVDCx20_ASAP7_75t_R g240 ( 
.A(n_214),
.Y(n_240)
);

NAND2xp5_ASAP7_75t_L g242 ( 
.A(n_226),
.B(n_54),
.Y(n_242)
);

NOR2xp33_ASAP7_75t_SL g325 ( 
.A(n_242),
.B(n_251),
.Y(n_325)
);

INVx3_ASAP7_75t_L g244 ( 
.A(n_165),
.Y(n_244)
);

INVx3_ASAP7_75t_L g337 ( 
.A(n_244),
.Y(n_337)
);

AND2x2_ASAP7_75t_L g247 ( 
.A(n_195),
.B(n_76),
.Y(n_247)
);

CKINVDCx14_ASAP7_75t_R g378 ( 
.A(n_247),
.Y(n_378)
);

BUFx2_ASAP7_75t_L g249 ( 
.A(n_193),
.Y(n_249)
);

BUFx3_ASAP7_75t_L g342 ( 
.A(n_249),
.Y(n_342)
);

NAND2xp5_ASAP7_75t_SL g250 ( 
.A(n_169),
.B(n_180),
.Y(n_250)
);

NAND2xp5_ASAP7_75t_SL g251 ( 
.A(n_169),
.B(n_161),
.Y(n_251)
);

CKINVDCx20_ASAP7_75t_R g252 ( 
.A(n_214),
.Y(n_252)
);

NAND2xp5_ASAP7_75t_SL g364 ( 
.A(n_252),
.B(n_253),
.Y(n_364)
);

CKINVDCx20_ASAP7_75t_R g253 ( 
.A(n_193),
.Y(n_253)
);

BUFx6f_ASAP7_75t_L g255 ( 
.A(n_148),
.Y(n_255)
);

INVx8_ASAP7_75t_L g318 ( 
.A(n_255),
.Y(n_318)
);

NOR2xp33_ASAP7_75t_L g256 ( 
.A(n_161),
.B(n_109),
.Y(n_256)
);

NOR2xp33_ASAP7_75t_L g328 ( 
.A(n_256),
.B(n_258),
.Y(n_328)
);

BUFx2_ASAP7_75t_L g257 ( 
.A(n_230),
.Y(n_257)
);

BUFx3_ASAP7_75t_L g345 ( 
.A(n_257),
.Y(n_345)
);

CKINVDCx20_ASAP7_75t_R g258 ( 
.A(n_160),
.Y(n_258)
);

CKINVDCx16_ASAP7_75t_R g259 ( 
.A(n_137),
.Y(n_259)
);

NOR2xp33_ASAP7_75t_L g334 ( 
.A(n_259),
.B(n_267),
.Y(n_334)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_151),
.Y(n_260)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_260),
.Y(n_321)
);

INVx3_ASAP7_75t_L g261 ( 
.A(n_138),
.Y(n_261)
);

INVx2_ASAP7_75t_L g353 ( 
.A(n_261),
.Y(n_353)
);

INVxp67_ASAP7_75t_L g348 ( 
.A(n_263),
.Y(n_348)
);

INVxp67_ASAP7_75t_L g264 ( 
.A(n_209),
.Y(n_264)
);

INVxp67_ASAP7_75t_L g350 ( 
.A(n_264),
.Y(n_350)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_162),
.Y(n_266)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_266),
.Y(n_324)
);

NOR2xp33_ASAP7_75t_L g267 ( 
.A(n_228),
.B(n_167),
.Y(n_267)
);

INVx6_ASAP7_75t_L g268 ( 
.A(n_184),
.Y(n_268)
);

INVx2_ASAP7_75t_L g354 ( 
.A(n_268),
.Y(n_354)
);

NAND2xp5_ASAP7_75t_SL g269 ( 
.A(n_198),
.B(n_38),
.Y(n_269)
);

NAND2x1p5_ASAP7_75t_L g270 ( 
.A(n_198),
.B(n_85),
.Y(n_270)
);

NOR2xp33_ASAP7_75t_L g271 ( 
.A(n_170),
.B(n_185),
.Y(n_271)
);

NOR2xp33_ASAP7_75t_L g341 ( 
.A(n_271),
.B(n_284),
.Y(n_341)
);

BUFx6f_ASAP7_75t_L g272 ( 
.A(n_184),
.Y(n_272)
);

INVx2_ASAP7_75t_L g356 ( 
.A(n_272),
.Y(n_356)
);

AND2x2_ASAP7_75t_SL g273 ( 
.A(n_136),
.B(n_141),
.Y(n_273)
);

CKINVDCx16_ASAP7_75t_R g355 ( 
.A(n_273),
.Y(n_355)
);

INVx3_ASAP7_75t_L g276 ( 
.A(n_203),
.Y(n_276)
);

INVx2_ASAP7_75t_L g358 ( 
.A(n_276),
.Y(n_358)
);

INVx3_ASAP7_75t_L g277 ( 
.A(n_145),
.Y(n_277)
);

INVx2_ASAP7_75t_L g362 ( 
.A(n_277),
.Y(n_362)
);

INVx6_ASAP7_75t_L g278 ( 
.A(n_186),
.Y(n_278)
);

INVx2_ASAP7_75t_L g372 ( 
.A(n_278),
.Y(n_372)
);

AOI22xp33_ASAP7_75t_SL g332 ( 
.A1(n_279),
.A2(n_283),
.B1(n_309),
.B2(n_220),
.Y(n_332)
);

OAI21xp5_ASAP7_75t_L g280 ( 
.A1(n_202),
.A2(n_65),
.B(n_84),
.Y(n_280)
);

OAI21xp5_ASAP7_75t_L g336 ( 
.A1(n_280),
.A2(n_220),
.B(n_177),
.Y(n_336)
);

OAI22xp5_ASAP7_75t_L g366 ( 
.A1(n_281),
.A2(n_306),
.B1(n_218),
.B2(n_215),
.Y(n_366)
);

NAND2xp5_ASAP7_75t_L g282 ( 
.A(n_212),
.B(n_2),
.Y(n_282)
);

AOI21xp33_ASAP7_75t_L g367 ( 
.A1(n_282),
.A2(n_286),
.B(n_288),
.Y(n_367)
);

AOI22xp33_ASAP7_75t_SL g283 ( 
.A1(n_178),
.A2(n_52),
.B1(n_47),
.B2(n_4),
.Y(n_283)
);

NOR2xp33_ASAP7_75t_L g284 ( 
.A(n_140),
.B(n_2),
.Y(n_284)
);

NAND2xp5_ASAP7_75t_SL g286 ( 
.A(n_142),
.B(n_3),
.Y(n_286)
);

INVx4_ASAP7_75t_L g287 ( 
.A(n_166),
.Y(n_287)
);

INVx2_ASAP7_75t_L g376 ( 
.A(n_287),
.Y(n_376)
);

NAND2xp5_ASAP7_75t_L g288 ( 
.A(n_224),
.B(n_3),
.Y(n_288)
);

NOR2xp33_ASAP7_75t_L g291 ( 
.A(n_140),
.B(n_3),
.Y(n_291)
);

NOR2xp33_ASAP7_75t_L g346 ( 
.A(n_291),
.B(n_293),
.Y(n_346)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_143),
.Y(n_292)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_292),
.Y(n_331)
);

NAND2xp5_ASAP7_75t_L g293 ( 
.A(n_194),
.B(n_4),
.Y(n_293)
);

OAI22xp33_ASAP7_75t_L g294 ( 
.A1(n_156),
.A2(n_52),
.B1(n_47),
.B2(n_8),
.Y(n_294)
);

AOI22xp5_ASAP7_75t_L g359 ( 
.A1(n_294),
.A2(n_137),
.B1(n_149),
.B2(n_158),
.Y(n_359)
);

NOR2xp33_ASAP7_75t_L g296 ( 
.A(n_179),
.B(n_6),
.Y(n_296)
);

NOR2xp33_ASAP7_75t_L g352 ( 
.A(n_296),
.B(n_303),
.Y(n_352)
);

INVx6_ASAP7_75t_L g298 ( 
.A(n_231),
.Y(n_298)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_298),
.Y(n_335)
);

INVx2_ASAP7_75t_L g302 ( 
.A(n_207),
.Y(n_302)
);

INVx1_ASAP7_75t_L g343 ( 
.A(n_302),
.Y(n_343)
);

BUFx6f_ASAP7_75t_L g305 ( 
.A(n_186),
.Y(n_305)
);

INVx1_ASAP7_75t_L g349 ( 
.A(n_305),
.Y(n_349)
);

AOI22xp33_ASAP7_75t_L g306 ( 
.A1(n_163),
.A2(n_52),
.B1(n_8),
.B2(n_9),
.Y(n_306)
);

INVx3_ASAP7_75t_L g308 ( 
.A(n_176),
.Y(n_308)
);

INVx1_ASAP7_75t_L g351 ( 
.A(n_308),
.Y(n_351)
);

AOI22xp33_ASAP7_75t_SL g309 ( 
.A1(n_225),
.A2(n_6),
.B1(n_9),
.B2(n_10),
.Y(n_309)
);

NOR2xp33_ASAP7_75t_L g310 ( 
.A(n_139),
.B(n_9),
.Y(n_310)
);

CKINVDCx20_ASAP7_75t_R g320 ( 
.A(n_310),
.Y(n_320)
);

NOR2xp33_ASAP7_75t_SL g311 ( 
.A(n_213),
.B(n_10),
.Y(n_311)
);

INVx1_ASAP7_75t_L g360 ( 
.A(n_311),
.Y(n_360)
);

INVx6_ASAP7_75t_L g312 ( 
.A(n_188),
.Y(n_312)
);

INVx1_ASAP7_75t_L g361 ( 
.A(n_312),
.Y(n_361)
);

OR2x2_ASAP7_75t_SL g314 ( 
.A(n_159),
.B(n_10),
.Y(n_314)
);

MAJIxp5_ASAP7_75t_L g340 ( 
.A(n_314),
.B(n_177),
.C(n_160),
.Y(n_340)
);

NOR2xp33_ASAP7_75t_L g315 ( 
.A(n_152),
.B(n_10),
.Y(n_315)
);

NAND2xp5_ASAP7_75t_L g327 ( 
.A(n_315),
.B(n_316),
.Y(n_327)
);

NAND2xp5_ASAP7_75t_L g316 ( 
.A(n_210),
.B(n_11),
.Y(n_316)
);

INVx2_ASAP7_75t_L g317 ( 
.A(n_174),
.Y(n_317)
);

INVx1_ASAP7_75t_L g379 ( 
.A(n_317),
.Y(n_379)
);

INVx13_ASAP7_75t_L g319 ( 
.A(n_313),
.Y(n_319)
);

INVx1_ASAP7_75t_SL g426 ( 
.A(n_319),
.Y(n_426)
);

BUFx8_ASAP7_75t_L g326 ( 
.A(n_313),
.Y(n_326)
);

INVx13_ASAP7_75t_L g411 ( 
.A(n_326),
.Y(n_411)
);

AOI22xp33_ASAP7_75t_L g329 ( 
.A1(n_264),
.A2(n_171),
.B1(n_187),
.B2(n_189),
.Y(n_329)
);

OA22x2_ASAP7_75t_L g421 ( 
.A1(n_329),
.A2(n_357),
.B1(n_373),
.B2(n_287),
.Y(n_421)
);

INVxp67_ASAP7_75t_L g424 ( 
.A(n_332),
.Y(n_424)
);

OAI22xp5_ASAP7_75t_SL g333 ( 
.A1(n_281),
.A2(n_164),
.B1(n_135),
.B2(n_133),
.Y(n_333)
);

AOI22xp5_ASAP7_75t_L g394 ( 
.A1(n_333),
.A2(n_359),
.B1(n_368),
.B2(n_247),
.Y(n_394)
);

CKINVDCx16_ASAP7_75t_R g416 ( 
.A(n_336),
.Y(n_416)
);

O2A1O1Ixp33_ASAP7_75t_L g338 ( 
.A1(n_280),
.A2(n_181),
.B(n_183),
.C(n_134),
.Y(n_338)
);

AOI21xp5_ASAP7_75t_L g428 ( 
.A1(n_338),
.A2(n_274),
.B(n_249),
.Y(n_428)
);

CKINVDCx14_ASAP7_75t_R g406 ( 
.A(n_340),
.Y(n_406)
);

NAND2xp5_ASAP7_75t_L g347 ( 
.A(n_270),
.B(n_201),
.Y(n_347)
);

NAND2xp5_ASAP7_75t_L g382 ( 
.A(n_347),
.B(n_371),
.Y(n_382)
);

AOI22xp33_ASAP7_75t_L g357 ( 
.A1(n_279),
.A2(n_231),
.B1(n_199),
.B2(n_188),
.Y(n_357)
);

AOI22xp33_ASAP7_75t_SL g363 ( 
.A1(n_238),
.A2(n_217),
.B1(n_191),
.B2(n_190),
.Y(n_363)
);

AOI22xp33_ASAP7_75t_SL g407 ( 
.A1(n_363),
.A2(n_366),
.B1(n_369),
.B2(n_246),
.Y(n_407)
);

XNOR2xp5_ASAP7_75t_L g365 ( 
.A(n_233),
.B(n_149),
.Y(n_365)
);

XNOR2xp5_ASAP7_75t_L g417 ( 
.A(n_365),
.B(n_275),
.Y(n_417)
);

OAI22xp33_ASAP7_75t_L g368 ( 
.A1(n_294),
.A2(n_206),
.B1(n_199),
.B2(n_196),
.Y(n_368)
);

AOI22xp33_ASAP7_75t_SL g369 ( 
.A1(n_238),
.A2(n_192),
.B1(n_147),
.B2(n_211),
.Y(n_369)
);

NAND2xp5_ASAP7_75t_L g371 ( 
.A(n_270),
.B(n_196),
.Y(n_371)
);

AOI22xp33_ASAP7_75t_L g373 ( 
.A1(n_317),
.A2(n_147),
.B1(n_12),
.B2(n_14),
.Y(n_373)
);

NAND2xp5_ASAP7_75t_L g374 ( 
.A(n_273),
.B(n_11),
.Y(n_374)
);

NAND2xp5_ASAP7_75t_L g383 ( 
.A(n_374),
.B(n_273),
.Y(n_383)
);

INVx13_ASAP7_75t_L g375 ( 
.A(n_246),
.Y(n_375)
);

BUFx16f_ASAP7_75t_L g404 ( 
.A(n_375),
.Y(n_404)
);

AOI32xp33_ASAP7_75t_L g377 ( 
.A1(n_254),
.A2(n_146),
.A3(n_15),
.B1(n_16),
.B2(n_12),
.Y(n_377)
);

NOR2xp33_ASAP7_75t_L g398 ( 
.A(n_377),
.B(n_297),
.Y(n_398)
);

BUFx6f_ASAP7_75t_L g380 ( 
.A(n_356),
.Y(n_380)
);

INVxp67_ASAP7_75t_L g431 ( 
.A(n_380),
.Y(n_431)
);

INVx1_ASAP7_75t_L g381 ( 
.A(n_343),
.Y(n_381)
);

INVx1_ASAP7_75t_L g434 ( 
.A(n_381),
.Y(n_434)
);

NAND2xp5_ASAP7_75t_SL g445 ( 
.A(n_383),
.B(n_403),
.Y(n_445)
);

CKINVDCx20_ASAP7_75t_R g384 ( 
.A(n_339),
.Y(n_384)
);

NOR2xp33_ASAP7_75t_SL g429 ( 
.A(n_384),
.B(n_388),
.Y(n_429)
);

INVx3_ASAP7_75t_L g385 ( 
.A(n_323),
.Y(n_385)
);

INVx1_ASAP7_75t_L g439 ( 
.A(n_385),
.Y(n_439)
);

NAND2xp5_ASAP7_75t_L g386 ( 
.A(n_352),
.B(n_304),
.Y(n_386)
);

NAND2xp5_ASAP7_75t_L g430 ( 
.A(n_386),
.B(n_413),
.Y(n_430)
);

INVx1_ASAP7_75t_L g387 ( 
.A(n_343),
.Y(n_387)
);

INVx1_ASAP7_75t_L g441 ( 
.A(n_387),
.Y(n_441)
);

NAND2xp5_ASAP7_75t_SL g388 ( 
.A(n_325),
.B(n_241),
.Y(n_388)
);

INVx1_ASAP7_75t_L g389 ( 
.A(n_379),
.Y(n_389)
);

INVx1_ASAP7_75t_L g442 ( 
.A(n_389),
.Y(n_442)
);

NAND2xp5_ASAP7_75t_SL g390 ( 
.A(n_325),
.B(n_303),
.Y(n_390)
);

NOR2xp33_ASAP7_75t_SL g435 ( 
.A(n_390),
.B(n_393),
.Y(n_435)
);

AND2x2_ASAP7_75t_SL g391 ( 
.A(n_347),
.B(n_238),
.Y(n_391)
);

AND2x2_ASAP7_75t_L g444 ( 
.A(n_391),
.B(n_394),
.Y(n_444)
);

OAI21xp5_ASAP7_75t_SL g392 ( 
.A1(n_371),
.A2(n_314),
.B(n_247),
.Y(n_392)
);

OAI21xp5_ASAP7_75t_L g432 ( 
.A1(n_392),
.A2(n_414),
.B(n_336),
.Y(n_432)
);

CKINVDCx20_ASAP7_75t_R g393 ( 
.A(n_322),
.Y(n_393)
);

OAI22xp5_ASAP7_75t_L g395 ( 
.A1(n_348),
.A2(n_302),
.B1(n_278),
.B2(n_312),
.Y(n_395)
);

AOI22xp5_ASAP7_75t_L g447 ( 
.A1(n_395),
.A2(n_397),
.B1(n_408),
.B2(n_410),
.Y(n_447)
);

NAND2xp5_ASAP7_75t_SL g396 ( 
.A(n_344),
.B(n_248),
.Y(n_396)
);

NAND2xp5_ASAP7_75t_SL g457 ( 
.A(n_396),
.B(n_402),
.Y(n_457)
);

OAI22xp5_ASAP7_75t_L g397 ( 
.A1(n_348),
.A2(n_298),
.B1(n_268),
.B2(n_272),
.Y(n_397)
);

INVxp67_ASAP7_75t_L g433 ( 
.A(n_398),
.Y(n_433)
);

INVx1_ASAP7_75t_L g399 ( 
.A(n_379),
.Y(n_399)
);

INVx1_ASAP7_75t_L g464 ( 
.A(n_399),
.Y(n_464)
);

BUFx3_ASAP7_75t_L g400 ( 
.A(n_326),
.Y(n_400)
);

INVx1_ASAP7_75t_L g470 ( 
.A(n_400),
.Y(n_470)
);

INVx1_ASAP7_75t_L g401 ( 
.A(n_331),
.Y(n_401)
);

AND2x2_ASAP7_75t_L g448 ( 
.A(n_401),
.B(n_409),
.Y(n_448)
);

NAND2xp5_ASAP7_75t_SL g402 ( 
.A(n_327),
.B(n_262),
.Y(n_402)
);

NOR2xp33_ASAP7_75t_L g403 ( 
.A(n_320),
.B(n_341),
.Y(n_403)
);

AOI22xp5_ASAP7_75t_L g405 ( 
.A1(n_333),
.A2(n_290),
.B1(n_285),
.B2(n_301),
.Y(n_405)
);

OAI22xp5_ASAP7_75t_L g452 ( 
.A1(n_405),
.A2(n_422),
.B1(n_335),
.B2(n_361),
.Y(n_452)
);

AOI22xp33_ASAP7_75t_SL g463 ( 
.A1(n_407),
.A2(n_420),
.B1(n_427),
.B2(n_342),
.Y(n_463)
);

OAI22xp5_ASAP7_75t_SL g408 ( 
.A1(n_355),
.A2(n_275),
.B1(n_245),
.B2(n_243),
.Y(n_408)
);

INVx1_ASAP7_75t_L g409 ( 
.A(n_331),
.Y(n_409)
);

OAI22xp5_ASAP7_75t_L g410 ( 
.A1(n_330),
.A2(n_305),
.B1(n_235),
.B2(n_255),
.Y(n_410)
);

INVx1_ASAP7_75t_L g412 ( 
.A(n_321),
.Y(n_412)
);

NAND2xp5_ASAP7_75t_SL g467 ( 
.A(n_412),
.B(n_415),
.Y(n_467)
);

CKINVDCx20_ASAP7_75t_R g413 ( 
.A(n_364),
.Y(n_413)
);

OAI21xp5_ASAP7_75t_L g414 ( 
.A1(n_350),
.A2(n_244),
.B(n_307),
.Y(n_414)
);

NOR2xp33_ASAP7_75t_SL g415 ( 
.A(n_346),
.B(n_276),
.Y(n_415)
);

XOR2xp5_ASAP7_75t_L g443 ( 
.A(n_417),
.B(n_365),
.Y(n_443)
);

AOI21xp5_ASAP7_75t_L g418 ( 
.A1(n_350),
.A2(n_308),
.B(n_277),
.Y(n_418)
);

AOI21xp5_ASAP7_75t_L g436 ( 
.A1(n_418),
.A2(n_428),
.B(n_338),
.Y(n_436)
);

AND2x6_ASAP7_75t_L g419 ( 
.A(n_328),
.B(n_295),
.Y(n_419)
);

NAND2xp5_ASAP7_75t_L g446 ( 
.A(n_419),
.B(n_423),
.Y(n_446)
);

AOI22xp33_ASAP7_75t_L g420 ( 
.A1(n_378),
.A2(n_261),
.B1(n_301),
.B2(n_300),
.Y(n_420)
);

CKINVDCx16_ASAP7_75t_R g437 ( 
.A(n_421),
.Y(n_437)
);

AOI22xp5_ASAP7_75t_L g422 ( 
.A1(n_368),
.A2(n_289),
.B1(n_300),
.B2(n_299),
.Y(n_422)
);

NAND2xp5_ASAP7_75t_SL g423 ( 
.A(n_327),
.B(n_243),
.Y(n_423)
);

INVx1_ASAP7_75t_L g425 ( 
.A(n_321),
.Y(n_425)
);

NAND2xp5_ASAP7_75t_L g449 ( 
.A(n_425),
.B(n_370),
.Y(n_449)
);

INVx2_ASAP7_75t_L g427 ( 
.A(n_354),
.Y(n_427)
);

INVx1_ASAP7_75t_SL g499 ( 
.A(n_432),
.Y(n_499)
);

AND2x2_ASAP7_75t_L g474 ( 
.A(n_436),
.B(n_469),
.Y(n_474)
);

OAI22xp5_ASAP7_75t_SL g438 ( 
.A1(n_382),
.A2(n_320),
.B1(n_374),
.B2(n_359),
.Y(n_438)
);

NAND2xp5_ASAP7_75t_L g472 ( 
.A(n_438),
.B(n_450),
.Y(n_472)
);

CKINVDCx20_ASAP7_75t_R g440 ( 
.A(n_404),
.Y(n_440)
);

INVx13_ASAP7_75t_L g473 ( 
.A(n_440),
.Y(n_473)
);

XOR2xp5_ASAP7_75t_L g476 ( 
.A(n_443),
.B(n_462),
.Y(n_476)
);

INVx1_ASAP7_75t_L g471 ( 
.A(n_449),
.Y(n_471)
);

NAND2xp5_ASAP7_75t_L g450 ( 
.A(n_382),
.B(n_367),
.Y(n_450)
);

AOI22xp5_ASAP7_75t_L g451 ( 
.A1(n_416),
.A2(n_340),
.B1(n_360),
.B2(n_361),
.Y(n_451)
);

OAI22xp5_ASAP7_75t_SL g477 ( 
.A1(n_451),
.A2(n_386),
.B1(n_418),
.B2(n_414),
.Y(n_477)
);

AOI22xp33_ASAP7_75t_L g505 ( 
.A1(n_452),
.A2(n_456),
.B1(n_458),
.B2(n_463),
.Y(n_505)
);

AOI21xp5_ASAP7_75t_L g453 ( 
.A1(n_428),
.A2(n_326),
.B(n_319),
.Y(n_453)
);

OAI21xp5_ASAP7_75t_L g479 ( 
.A1(n_453),
.A2(n_461),
.B(n_426),
.Y(n_479)
);

OAI32xp33_ASAP7_75t_L g454 ( 
.A1(n_383),
.A2(n_360),
.A3(n_334),
.B1(n_370),
.B2(n_324),
.Y(n_454)
);

INVxp67_ASAP7_75t_L g486 ( 
.A(n_454),
.Y(n_486)
);

MAJIxp5_ASAP7_75t_L g455 ( 
.A(n_406),
.B(n_324),
.C(n_351),
.Y(n_455)
);

XNOR2xp5_ASAP7_75t_L g488 ( 
.A(n_455),
.B(n_401),
.Y(n_488)
);

OAI22xp5_ASAP7_75t_L g456 ( 
.A1(n_416),
.A2(n_335),
.B1(n_349),
.B2(n_372),
.Y(n_456)
);

OAI22xp5_ASAP7_75t_L g458 ( 
.A1(n_394),
.A2(n_349),
.B1(n_372),
.B2(n_354),
.Y(n_458)
);

NAND2xp5_ASAP7_75t_L g459 ( 
.A(n_423),
.B(n_351),
.Y(n_459)
);

NAND2xp5_ASAP7_75t_L g475 ( 
.A(n_459),
.B(n_460),
.Y(n_475)
);

NAND2xp5_ASAP7_75t_L g460 ( 
.A(n_417),
.B(n_358),
.Y(n_460)
);

OAI21xp5_ASAP7_75t_L g461 ( 
.A1(n_392),
.A2(n_353),
.B(n_358),
.Y(n_461)
);

XNOR2xp5_ASAP7_75t_L g462 ( 
.A(n_391),
.B(n_362),
.Y(n_462)
);

XOR2xp5_ASAP7_75t_L g465 ( 
.A(n_391),
.B(n_353),
.Y(n_465)
);

XOR2xp5_ASAP7_75t_L g480 ( 
.A(n_465),
.B(n_408),
.Y(n_480)
);

NAND2xp5_ASAP7_75t_L g466 ( 
.A(n_413),
.B(n_362),
.Y(n_466)
);

NAND2xp5_ASAP7_75t_L g484 ( 
.A(n_466),
.B(n_468),
.Y(n_484)
);

OAI22xp5_ASAP7_75t_L g468 ( 
.A1(n_424),
.A2(n_356),
.B1(n_323),
.B2(n_318),
.Y(n_468)
);

CKINVDCx20_ASAP7_75t_R g469 ( 
.A(n_404),
.Y(n_469)
);

NAND2xp5_ASAP7_75t_SL g513 ( 
.A(n_477),
.B(n_451),
.Y(n_513)
);

NOR2xp33_ASAP7_75t_SL g478 ( 
.A(n_430),
.B(n_393),
.Y(n_478)
);

NOR2xp33_ASAP7_75t_L g523 ( 
.A(n_478),
.B(n_493),
.Y(n_523)
);

OAI21xp5_ASAP7_75t_SL g520 ( 
.A1(n_479),
.A2(n_506),
.B(n_456),
.Y(n_520)
);

XOR2xp5_ASAP7_75t_L g514 ( 
.A(n_480),
.B(n_488),
.Y(n_514)
);

CKINVDCx20_ASAP7_75t_R g481 ( 
.A(n_448),
.Y(n_481)
);

CKINVDCx5p33_ASAP7_75t_R g541 ( 
.A(n_481),
.Y(n_541)
);

OAI22xp5_ASAP7_75t_SL g482 ( 
.A1(n_444),
.A2(n_424),
.B1(n_422),
.B2(n_405),
.Y(n_482)
);

AOI22xp5_ASAP7_75t_L g512 ( 
.A1(n_482),
.A2(n_495),
.B1(n_496),
.B2(n_503),
.Y(n_512)
);

AND2x2_ASAP7_75t_L g483 ( 
.A(n_461),
.B(n_436),
.Y(n_483)
);

AND2x2_ASAP7_75t_L g538 ( 
.A(n_483),
.B(n_490),
.Y(n_538)
);

INVx1_ASAP7_75t_L g485 ( 
.A(n_448),
.Y(n_485)
);

INVx1_ASAP7_75t_L g516 ( 
.A(n_485),
.Y(n_516)
);

NAND2xp5_ASAP7_75t_L g487 ( 
.A(n_467),
.B(n_409),
.Y(n_487)
);

INVx1_ASAP7_75t_L g519 ( 
.A(n_487),
.Y(n_519)
);

XNOR2xp5_ASAP7_75t_L g489 ( 
.A(n_445),
.B(n_415),
.Y(n_489)
);

XOR2xp5_ASAP7_75t_L g529 ( 
.A(n_489),
.B(n_460),
.Y(n_529)
);

OAI21xp33_ASAP7_75t_L g490 ( 
.A1(n_430),
.A2(n_388),
.B(n_419),
.Y(n_490)
);

NAND2xp5_ASAP7_75t_L g491 ( 
.A(n_467),
.B(n_384),
.Y(n_491)
);

INVx1_ASAP7_75t_L g532 ( 
.A(n_491),
.Y(n_532)
);

AND2x6_ASAP7_75t_L g492 ( 
.A(n_446),
.B(n_410),
.Y(n_492)
);

NAND2xp5_ASAP7_75t_L g517 ( 
.A(n_492),
.B(n_497),
.Y(n_517)
);

NAND2xp5_ASAP7_75t_SL g493 ( 
.A(n_435),
.B(n_412),
.Y(n_493)
);

NOR2xp33_ASAP7_75t_L g494 ( 
.A(n_435),
.B(n_337),
.Y(n_494)
);

NOR2xp33_ASAP7_75t_L g521 ( 
.A(n_494),
.B(n_501),
.Y(n_521)
);

OAI22xp5_ASAP7_75t_SL g495 ( 
.A1(n_444),
.A2(n_421),
.B1(n_425),
.B2(n_389),
.Y(n_495)
);

OAI22xp5_ASAP7_75t_SL g496 ( 
.A1(n_444),
.A2(n_421),
.B1(n_399),
.B2(n_387),
.Y(n_496)
);

NAND2xp5_ASAP7_75t_L g497 ( 
.A(n_459),
.B(n_466),
.Y(n_497)
);

NAND2xp5_ASAP7_75t_SL g498 ( 
.A(n_429),
.B(n_381),
.Y(n_498)
);

NOR2xp33_ASAP7_75t_L g524 ( 
.A(n_498),
.B(n_507),
.Y(n_524)
);

NAND2xp5_ASAP7_75t_L g500 ( 
.A(n_429),
.B(n_427),
.Y(n_500)
);

NAND2xp5_ASAP7_75t_L g525 ( 
.A(n_500),
.B(n_504),
.Y(n_525)
);

NOR2xp33_ASAP7_75t_L g501 ( 
.A(n_457),
.B(n_337),
.Y(n_501)
);

XOR2xp5_ASAP7_75t_L g502 ( 
.A(n_443),
.B(n_404),
.Y(n_502)
);

MAJIxp5_ASAP7_75t_L g518 ( 
.A(n_502),
.B(n_455),
.C(n_465),
.Y(n_518)
);

OAI22xp5_ASAP7_75t_SL g503 ( 
.A1(n_437),
.A2(n_421),
.B1(n_397),
.B2(n_385),
.Y(n_503)
);

INVx1_ASAP7_75t_L g504 ( 
.A(n_448),
.Y(n_504)
);

OA21x2_ASAP7_75t_L g506 ( 
.A1(n_446),
.A2(n_395),
.B(n_376),
.Y(n_506)
);

INVx1_ASAP7_75t_L g507 ( 
.A(n_434),
.Y(n_507)
);

CKINVDCx20_ASAP7_75t_R g508 ( 
.A(n_449),
.Y(n_508)
);

NOR2xp33_ASAP7_75t_L g544 ( 
.A(n_508),
.B(n_245),
.Y(n_544)
);

NAND2xp5_ASAP7_75t_L g509 ( 
.A(n_445),
.B(n_380),
.Y(n_509)
);

NAND2xp5_ASAP7_75t_L g536 ( 
.A(n_509),
.B(n_439),
.Y(n_536)
);

AOI21xp5_ASAP7_75t_L g510 ( 
.A1(n_483),
.A2(n_453),
.B(n_432),
.Y(n_510)
);

OAI21xp5_ASAP7_75t_SL g571 ( 
.A1(n_510),
.A2(n_513),
.B(n_520),
.Y(n_571)
);

CKINVDCx20_ASAP7_75t_R g511 ( 
.A(n_491),
.Y(n_511)
);

NOR2xp33_ASAP7_75t_L g549 ( 
.A(n_511),
.B(n_527),
.Y(n_549)
);

OAI22xp5_ASAP7_75t_L g515 ( 
.A1(n_471),
.A2(n_437),
.B1(n_447),
.B2(n_458),
.Y(n_515)
);

OAI22xp5_ASAP7_75t_L g561 ( 
.A1(n_515),
.A2(n_526),
.B1(n_540),
.B2(n_542),
.Y(n_561)
);

XOR2xp5_ASAP7_75t_L g552 ( 
.A(n_518),
.B(n_489),
.Y(n_552)
);

NAND2xp5_ASAP7_75t_SL g522 ( 
.A(n_504),
.B(n_450),
.Y(n_522)
);

INVx1_ASAP7_75t_L g554 ( 
.A(n_522),
.Y(n_554)
);

AOI22xp5_ASAP7_75t_L g526 ( 
.A1(n_486),
.A2(n_438),
.B1(n_433),
.B2(n_447),
.Y(n_526)
);

AOI21xp5_ASAP7_75t_SL g527 ( 
.A1(n_486),
.A2(n_454),
.B(n_462),
.Y(n_527)
);

OAI21xp5_ASAP7_75t_L g528 ( 
.A1(n_499),
.A2(n_434),
.B(n_441),
.Y(n_528)
);

INVx1_ASAP7_75t_SL g556 ( 
.A(n_528),
.Y(n_556)
);

XNOR2xp5_ASAP7_75t_SL g553 ( 
.A(n_529),
.B(n_477),
.Y(n_553)
);

MAJIxp5_ASAP7_75t_L g530 ( 
.A(n_476),
.B(n_441),
.C(n_464),
.Y(n_530)
);

MAJIxp5_ASAP7_75t_L g548 ( 
.A(n_530),
.B(n_537),
.C(n_502),
.Y(n_548)
);

OAI21xp5_ASAP7_75t_SL g531 ( 
.A1(n_483),
.A2(n_468),
.B(n_469),
.Y(n_531)
);

NAND2xp5_ASAP7_75t_SL g560 ( 
.A(n_531),
.B(n_474),
.Y(n_560)
);

INVx13_ASAP7_75t_L g533 ( 
.A(n_473),
.Y(n_533)
);

INVx1_ASAP7_75t_SL g574 ( 
.A(n_533),
.Y(n_574)
);

OAI21xp5_ASAP7_75t_L g534 ( 
.A1(n_499),
.A2(n_464),
.B(n_442),
.Y(n_534)
);

CKINVDCx16_ASAP7_75t_R g568 ( 
.A(n_534),
.Y(n_568)
);

OAI22xp5_ASAP7_75t_SL g535 ( 
.A1(n_472),
.A2(n_442),
.B1(n_439),
.B2(n_452),
.Y(n_535)
);

AOI22xp5_ASAP7_75t_L g576 ( 
.A1(n_535),
.A2(n_484),
.B1(n_482),
.B2(n_473),
.Y(n_576)
);

INVx1_ASAP7_75t_L g562 ( 
.A(n_536),
.Y(n_562)
);

MAJIxp5_ASAP7_75t_L g537 ( 
.A(n_476),
.B(n_440),
.C(n_470),
.Y(n_537)
);

NAND2xp5_ASAP7_75t_L g539 ( 
.A(n_487),
.B(n_431),
.Y(n_539)
);

INVx1_ASAP7_75t_L g563 ( 
.A(n_539),
.Y(n_563)
);

OAI22xp5_ASAP7_75t_L g540 ( 
.A1(n_471),
.A2(n_470),
.B1(n_426),
.B2(n_380),
.Y(n_540)
);

OAI22xp5_ASAP7_75t_L g542 ( 
.A1(n_505),
.A2(n_318),
.B1(n_400),
.B2(n_376),
.Y(n_542)
);

OR2x2_ASAP7_75t_L g543 ( 
.A(n_479),
.B(n_411),
.Y(n_543)
);

INVx1_ASAP7_75t_L g564 ( 
.A(n_543),
.Y(n_564)
);

INVx1_ASAP7_75t_L g555 ( 
.A(n_544),
.Y(n_555)
);

NAND2xp5_ASAP7_75t_L g545 ( 
.A(n_497),
.B(n_475),
.Y(n_545)
);

INVx1_ASAP7_75t_L g557 ( 
.A(n_545),
.Y(n_557)
);

NAND2xp5_ASAP7_75t_L g546 ( 
.A(n_475),
.B(n_290),
.Y(n_546)
);

INVx1_ASAP7_75t_L g558 ( 
.A(n_546),
.Y(n_558)
);

OR2x2_ASAP7_75t_L g547 ( 
.A(n_474),
.B(n_411),
.Y(n_547)
);

INVx1_ASAP7_75t_L g569 ( 
.A(n_547),
.Y(n_569)
);

XNOR2xp5_ASAP7_75t_L g580 ( 
.A(n_548),
.B(n_551),
.Y(n_580)
);

MAJIxp5_ASAP7_75t_L g550 ( 
.A(n_530),
.B(n_488),
.C(n_480),
.Y(n_550)
);

MAJIxp5_ASAP7_75t_L g584 ( 
.A(n_550),
.B(n_570),
.C(n_575),
.Y(n_584)
);

XNOR2xp5_ASAP7_75t_L g551 ( 
.A(n_514),
.B(n_472),
.Y(n_551)
);

XOR2xp5_ASAP7_75t_L g586 ( 
.A(n_552),
.B(n_565),
.Y(n_586)
);

XNOR2xp5_ASAP7_75t_SL g583 ( 
.A(n_553),
.B(n_538),
.Y(n_583)
);

XNOR2xp5_ASAP7_75t_L g559 ( 
.A(n_514),
.B(n_509),
.Y(n_559)
);

XNOR2xp5_ASAP7_75t_L g588 ( 
.A(n_559),
.B(n_535),
.Y(n_588)
);

NAND2xp5_ASAP7_75t_L g599 ( 
.A(n_560),
.B(n_541),
.Y(n_599)
);

XOR2xp5_ASAP7_75t_L g565 ( 
.A(n_518),
.B(n_537),
.Y(n_565)
);

XOR2xp5_ASAP7_75t_L g566 ( 
.A(n_527),
.B(n_474),
.Y(n_566)
);

XOR2xp5_ASAP7_75t_L g587 ( 
.A(n_566),
.B(n_572),
.Y(n_587)
);

OAI22xp5_ASAP7_75t_L g567 ( 
.A1(n_523),
.A2(n_526),
.B1(n_517),
.B2(n_512),
.Y(n_567)
);

AOI22xp5_ASAP7_75t_L g594 ( 
.A1(n_567),
.A2(n_573),
.B1(n_515),
.B2(n_519),
.Y(n_594)
);

MAJIxp5_ASAP7_75t_L g570 ( 
.A(n_529),
.B(n_500),
.C(n_506),
.Y(n_570)
);

XOR2xp5_ASAP7_75t_L g572 ( 
.A(n_522),
.B(n_506),
.Y(n_572)
);

OAI22xp5_ASAP7_75t_L g573 ( 
.A1(n_517),
.A2(n_484),
.B1(n_492),
.B2(n_503),
.Y(n_573)
);

MAJIxp5_ASAP7_75t_SL g575 ( 
.A(n_538),
.B(n_496),
.C(n_495),
.Y(n_575)
);

OAI22xp5_ASAP7_75t_SL g581 ( 
.A1(n_576),
.A2(n_512),
.B1(n_516),
.B2(n_511),
.Y(n_581)
);

XOR2xp5_ASAP7_75t_L g577 ( 
.A(n_513),
.B(n_375),
.Y(n_577)
);

XOR2xp5_ASAP7_75t_L g595 ( 
.A(n_577),
.B(n_540),
.Y(n_595)
);

INVx1_ASAP7_75t_L g578 ( 
.A(n_539),
.Y(n_578)
);

INVx1_ASAP7_75t_L g591 ( 
.A(n_578),
.Y(n_591)
);

OAI21xp5_ASAP7_75t_L g579 ( 
.A1(n_548),
.A2(n_538),
.B(n_516),
.Y(n_579)
);

OAI21x1_ASAP7_75t_L g610 ( 
.A1(n_579),
.A2(n_598),
.B(n_566),
.Y(n_610)
);

AOI22xp5_ASAP7_75t_L g605 ( 
.A1(n_581),
.A2(n_556),
.B1(n_568),
.B2(n_562),
.Y(n_605)
);

OAI21xp5_ASAP7_75t_L g582 ( 
.A1(n_571),
.A2(n_510),
.B(n_543),
.Y(n_582)
);

AOI21xp5_ASAP7_75t_L g623 ( 
.A1(n_582),
.A2(n_585),
.B(n_564),
.Y(n_623)
);

XNOR2xp5_ASAP7_75t_L g604 ( 
.A(n_583),
.B(n_588),
.Y(n_604)
);

OAI21xp5_ASAP7_75t_L g585 ( 
.A1(n_571),
.A2(n_543),
.B(n_520),
.Y(n_585)
);

XNOR2xp5_ASAP7_75t_L g589 ( 
.A(n_552),
.B(n_534),
.Y(n_589)
);

XNOR2xp5_ASAP7_75t_L g607 ( 
.A(n_589),
.B(n_592),
.Y(n_607)
);

CKINVDCx14_ASAP7_75t_R g590 ( 
.A(n_549),
.Y(n_590)
);

NAND2xp5_ASAP7_75t_L g613 ( 
.A(n_590),
.B(n_593),
.Y(n_613)
);

XNOR2xp5_ASAP7_75t_L g592 ( 
.A(n_565),
.B(n_528),
.Y(n_592)
);

MAJIxp5_ASAP7_75t_L g593 ( 
.A(n_550),
.B(n_547),
.C(n_531),
.Y(n_593)
);

OAI22xp5_ASAP7_75t_SL g620 ( 
.A1(n_594),
.A2(n_564),
.B1(n_558),
.B2(n_574),
.Y(n_620)
);

INVx1_ASAP7_75t_SL g608 ( 
.A(n_595),
.Y(n_608)
);

MAJIxp5_ASAP7_75t_L g596 ( 
.A(n_551),
.B(n_547),
.C(n_525),
.Y(n_596)
);

NAND2xp5_ASAP7_75t_L g615 ( 
.A(n_596),
.B(n_600),
.Y(n_615)
);

OAI22xp5_ASAP7_75t_SL g597 ( 
.A1(n_554),
.A2(n_532),
.B1(n_519),
.B2(n_524),
.Y(n_597)
);

HB1xp67_ASAP7_75t_L g619 ( 
.A(n_597),
.Y(n_619)
);

XOR2xp5_ASAP7_75t_L g598 ( 
.A(n_553),
.B(n_525),
.Y(n_598)
);

MAJIxp5_ASAP7_75t_L g616 ( 
.A(n_598),
.B(n_572),
.C(n_575),
.Y(n_616)
);

INVx1_ASAP7_75t_L g614 ( 
.A(n_599),
.Y(n_614)
);

NAND2xp5_ASAP7_75t_L g600 ( 
.A(n_555),
.B(n_521),
.Y(n_600)
);

AOI22xp5_ASAP7_75t_L g601 ( 
.A1(n_561),
.A2(n_557),
.B1(n_542),
.B2(n_563),
.Y(n_601)
);

INVxp67_ASAP7_75t_L g624 ( 
.A(n_601),
.Y(n_624)
);

XNOR2xp5_ASAP7_75t_SL g602 ( 
.A(n_559),
.B(n_545),
.Y(n_602)
);

NOR2xp33_ASAP7_75t_L g611 ( 
.A(n_602),
.B(n_592),
.Y(n_611)
);

OAI22xp5_ASAP7_75t_SL g603 ( 
.A1(n_576),
.A2(n_532),
.B1(n_521),
.B2(n_536),
.Y(n_603)
);

NAND2xp5_ASAP7_75t_SL g606 ( 
.A(n_603),
.B(n_541),
.Y(n_606)
);

INVx1_ASAP7_75t_L g634 ( 
.A(n_605),
.Y(n_634)
);

INVx1_ASAP7_75t_L g628 ( 
.A(n_606),
.Y(n_628)
);

BUFx12_ASAP7_75t_L g609 ( 
.A(n_602),
.Y(n_609)
);

INVx1_ASAP7_75t_L g637 ( 
.A(n_609),
.Y(n_637)
);

INVxp33_ASAP7_75t_L g627 ( 
.A(n_610),
.Y(n_627)
);

NOR2xp33_ASAP7_75t_L g632 ( 
.A(n_611),
.B(n_622),
.Y(n_632)
);

NOR2xp33_ASAP7_75t_L g612 ( 
.A(n_580),
.B(n_570),
.Y(n_612)
);

NOR2xp33_ASAP7_75t_SL g631 ( 
.A(n_612),
.B(n_617),
.Y(n_631)
);

XOR2xp5_ASAP7_75t_L g638 ( 
.A(n_616),
.B(n_623),
.Y(n_638)
);

NAND2xp5_ASAP7_75t_L g617 ( 
.A(n_591),
.B(n_563),
.Y(n_617)
);

AOI22xp5_ASAP7_75t_L g618 ( 
.A1(n_585),
.A2(n_556),
.B1(n_562),
.B2(n_569),
.Y(n_618)
);

OAI22xp5_ASAP7_75t_SL g629 ( 
.A1(n_618),
.A2(n_582),
.B1(n_595),
.B2(n_587),
.Y(n_629)
);

AOI22xp5_ASAP7_75t_L g640 ( 
.A1(n_620),
.A2(n_583),
.B1(n_533),
.B2(n_411),
.Y(n_640)
);

MAJIxp5_ASAP7_75t_L g621 ( 
.A(n_580),
.B(n_577),
.C(n_574),
.Y(n_621)
);

MAJIxp5_ASAP7_75t_L g625 ( 
.A(n_621),
.B(n_586),
.C(n_593),
.Y(n_625)
);

NOR2xp33_ASAP7_75t_SL g622 ( 
.A(n_589),
.B(n_546),
.Y(n_622)
);

NOR2xp33_ASAP7_75t_L g644 ( 
.A(n_625),
.B(n_608),
.Y(n_644)
);

NAND2xp5_ASAP7_75t_L g626 ( 
.A(n_614),
.B(n_588),
.Y(n_626)
);

AOI22xp5_ASAP7_75t_L g643 ( 
.A1(n_626),
.A2(n_629),
.B1(n_633),
.B2(n_635),
.Y(n_643)
);

AOI22xp33_ASAP7_75t_SL g630 ( 
.A1(n_619),
.A2(n_596),
.B1(n_584),
.B2(n_533),
.Y(n_630)
);

OAI22xp5_ASAP7_75t_SL g652 ( 
.A1(n_630),
.A2(n_640),
.B1(n_637),
.B2(n_634),
.Y(n_652)
);

NOR2xp33_ASAP7_75t_L g633 ( 
.A(n_624),
.B(n_584),
.Y(n_633)
);

INVx1_ASAP7_75t_L g635 ( 
.A(n_620),
.Y(n_635)
);

MAJIxp5_ASAP7_75t_L g636 ( 
.A(n_607),
.B(n_586),
.C(n_613),
.Y(n_636)
);

MAJIxp5_ASAP7_75t_L g653 ( 
.A(n_636),
.B(n_285),
.C(n_299),
.Y(n_653)
);

NAND2xp5_ASAP7_75t_L g639 ( 
.A(n_615),
.B(n_587),
.Y(n_639)
);

AOI21xp5_ASAP7_75t_L g646 ( 
.A1(n_639),
.A2(n_642),
.B(n_604),
.Y(n_646)
);

XOR2xp5_ASAP7_75t_L g641 ( 
.A(n_607),
.B(n_289),
.Y(n_641)
);

XOR2xp5_ASAP7_75t_L g645 ( 
.A(n_641),
.B(n_621),
.Y(n_645)
);

NOR2xp33_ASAP7_75t_L g642 ( 
.A(n_624),
.B(n_345),
.Y(n_642)
);

NAND2xp5_ASAP7_75t_L g663 ( 
.A(n_644),
.B(n_648),
.Y(n_663)
);

XNOR2xp5_ASAP7_75t_L g661 ( 
.A(n_645),
.B(n_651),
.Y(n_661)
);

INVx1_ASAP7_75t_L g658 ( 
.A(n_646),
.Y(n_658)
);

OAI21xp33_ASAP7_75t_L g647 ( 
.A1(n_627),
.A2(n_618),
.B(n_605),
.Y(n_647)
);

INVx1_ASAP7_75t_L g662 ( 
.A(n_647),
.Y(n_662)
);

AOI22xp5_ASAP7_75t_SL g648 ( 
.A1(n_628),
.A2(n_608),
.B1(n_609),
.B2(n_616),
.Y(n_648)
);

NOR2xp33_ASAP7_75t_L g649 ( 
.A(n_631),
.B(n_627),
.Y(n_649)
);

AOI21xp5_ASAP7_75t_L g664 ( 
.A1(n_649),
.A2(n_650),
.B(n_653),
.Y(n_664)
);

NOR2xp33_ASAP7_75t_L g650 ( 
.A(n_632),
.B(n_604),
.Y(n_650)
);

XOR2xp5_ASAP7_75t_L g651 ( 
.A(n_629),
.B(n_609),
.Y(n_651)
);

AOI22xp5_ASAP7_75t_L g656 ( 
.A1(n_652),
.A2(n_655),
.B1(n_640),
.B2(n_635),
.Y(n_656)
);

NOR2xp33_ASAP7_75t_L g654 ( 
.A(n_639),
.B(n_345),
.Y(n_654)
);

AOI22xp5_ASAP7_75t_L g659 ( 
.A1(n_654),
.A2(n_641),
.B1(n_638),
.B2(n_625),
.Y(n_659)
);

A2O1A1Ixp33_ASAP7_75t_SL g655 ( 
.A1(n_634),
.A2(n_307),
.B(n_297),
.C(n_295),
.Y(n_655)
);

OAI22xp5_ASAP7_75t_SL g667 ( 
.A1(n_656),
.A2(n_655),
.B1(n_265),
.B2(n_342),
.Y(n_667)
);

AOI21x1_ASAP7_75t_L g657 ( 
.A1(n_647),
.A2(n_626),
.B(n_636),
.Y(n_657)
);

HB1xp67_ASAP7_75t_L g666 ( 
.A(n_657),
.Y(n_666)
);

NAND2xp5_ASAP7_75t_L g669 ( 
.A(n_659),
.B(n_660),
.Y(n_669)
);

MAJIxp5_ASAP7_75t_L g660 ( 
.A(n_643),
.B(n_638),
.C(n_274),
.Y(n_660)
);

AOI322xp5_ASAP7_75t_L g665 ( 
.A1(n_658),
.A2(n_655),
.A3(n_651),
.B1(n_653),
.B2(n_645),
.C1(n_265),
.C2(n_295),
.Y(n_665)
);

INVx1_ASAP7_75t_L g673 ( 
.A(n_665),
.Y(n_673)
);

NOR2x1_ASAP7_75t_SL g672 ( 
.A(n_667),
.B(n_668),
.Y(n_672)
);

AND2x2_ASAP7_75t_L g668 ( 
.A(n_663),
.B(n_655),
.Y(n_668)
);

A2O1A1Ixp33_ASAP7_75t_L g670 ( 
.A1(n_662),
.A2(n_257),
.B(n_15),
.C(n_16),
.Y(n_670)
);

OAI21xp5_ASAP7_75t_SL g671 ( 
.A1(n_670),
.A2(n_656),
.B(n_664),
.Y(n_671)
);

NOR2xp33_ASAP7_75t_SL g675 ( 
.A(n_671),
.B(n_660),
.Y(n_675)
);

OAI21xp5_ASAP7_75t_L g674 ( 
.A1(n_673),
.A2(n_666),
.B(n_669),
.Y(n_674)
);

AOI21x1_ASAP7_75t_L g676 ( 
.A1(n_674),
.A2(n_675),
.B(n_672),
.Y(n_676)
);

INVx1_ASAP7_75t_L g677 ( 
.A(n_676),
.Y(n_677)
);

AOI21x1_ASAP7_75t_L g678 ( 
.A1(n_677),
.A2(n_661),
.B(n_15),
.Y(n_678)
);

MAJIxp5_ASAP7_75t_L g679 ( 
.A(n_678),
.B(n_12),
.C(n_16),
.Y(n_679)
);

NOR2xp33_ASAP7_75t_L g680 ( 
.A(n_679),
.B(n_661),
.Y(n_680)
);


endmodule