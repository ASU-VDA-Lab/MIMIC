module fake_jpeg_6346_n_308 (n_13, n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_308);

input n_13;
input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_308;

wire n_253;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_15;
wire n_141;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_286;
wire n_225;
wire n_105;
wire n_51;
wire n_84;
wire n_59;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_14;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_20;
wire n_18;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_208;
wire n_297;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_247;
wire n_157;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVx1_ASAP7_75t_L g14 ( 
.A(n_4),
.Y(n_14)
);

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_3),
.Y(n_15)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_9),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_11),
.Y(n_17)
);

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_12),
.Y(n_18)
);

BUFx5_ASAP7_75t_L g19 ( 
.A(n_9),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_1),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_7),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_10),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_4),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_3),
.Y(n_24)
);

NOR2xp33_ASAP7_75t_L g25 ( 
.A(n_0),
.B(n_8),
.Y(n_25)
);

AOI21xp5_ASAP7_75t_L g26 ( 
.A1(n_6),
.A2(n_3),
.B(n_13),
.Y(n_26)
);

INVx8_ASAP7_75t_L g27 ( 
.A(n_10),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_7),
.Y(n_28)
);

INVx4_ASAP7_75t_L g29 ( 
.A(n_7),
.Y(n_29)
);

INVx2_ASAP7_75t_L g30 ( 
.A(n_9),
.Y(n_30)
);

INVx13_ASAP7_75t_L g31 ( 
.A(n_11),
.Y(n_31)
);

BUFx3_ASAP7_75t_L g32 ( 
.A(n_12),
.Y(n_32)
);

INVx3_ASAP7_75t_L g33 ( 
.A(n_12),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_1),
.Y(n_34)
);

NAND2xp5_ASAP7_75t_SL g35 ( 
.A(n_14),
.B(n_0),
.Y(n_35)
);

NAND2xp5_ASAP7_75t_L g51 ( 
.A(n_35),
.B(n_37),
.Y(n_51)
);

BUFx5_ASAP7_75t_L g36 ( 
.A(n_19),
.Y(n_36)
);

BUFx3_ASAP7_75t_L g83 ( 
.A(n_36),
.Y(n_83)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_32),
.Y(n_37)
);

INVx8_ASAP7_75t_L g38 ( 
.A(n_32),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_38),
.B(n_42),
.Y(n_50)
);

AOI22xp5_ASAP7_75t_L g39 ( 
.A1(n_30),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_39)
);

OAI22xp5_ASAP7_75t_SL g52 ( 
.A1(n_39),
.A2(n_20),
.B1(n_16),
.B2(n_14),
.Y(n_52)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_17),
.Y(n_40)
);

NAND2xp5_ASAP7_75t_L g67 ( 
.A(n_40),
.B(n_41),
.Y(n_67)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_17),
.Y(n_41)
);

INVx2_ASAP7_75t_L g42 ( 
.A(n_32),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g43 ( 
.A(n_22),
.B(n_13),
.Y(n_43)
);

NAND2xp5_ASAP7_75t_SL g53 ( 
.A(n_43),
.B(n_22),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_19),
.Y(n_44)
);

BUFx3_ASAP7_75t_L g95 ( 
.A(n_44),
.Y(n_95)
);

BUFx3_ASAP7_75t_L g45 ( 
.A(n_18),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_45),
.B(n_31),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_L g46 ( 
.A(n_14),
.B(n_0),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_L g87 ( 
.A(n_46),
.B(n_20),
.Y(n_87)
);

AOI21xp5_ASAP7_75t_L g47 ( 
.A1(n_26),
.A2(n_1),
.B(n_2),
.Y(n_47)
);

MAJIxp5_ASAP7_75t_L g91 ( 
.A(n_47),
.B(n_20),
.C(n_16),
.Y(n_91)
);

INVx5_ASAP7_75t_L g48 ( 
.A(n_19),
.Y(n_48)
);

INVx5_ASAP7_75t_L g54 ( 
.A(n_48),
.Y(n_54)
);

INVx2_ASAP7_75t_L g49 ( 
.A(n_45),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_49),
.B(n_55),
.Y(n_110)
);

AND2x2_ASAP7_75t_L g109 ( 
.A(n_52),
.B(n_81),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_SL g120 ( 
.A(n_53),
.B(n_61),
.Y(n_120)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_45),
.Y(n_55)
);

CKINVDCx20_ASAP7_75t_R g56 ( 
.A(n_40),
.Y(n_56)
);

CKINVDCx20_ASAP7_75t_R g112 ( 
.A(n_56),
.Y(n_112)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_45),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g122 ( 
.A(n_57),
.B(n_58),
.Y(n_122)
);

INVx3_ASAP7_75t_L g58 ( 
.A(n_48),
.Y(n_58)
);

INVx4_ASAP7_75t_L g59 ( 
.A(n_48),
.Y(n_59)
);

INVx5_ASAP7_75t_L g118 ( 
.A(n_59),
.Y(n_118)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_48),
.Y(n_60)
);

INVx6_ASAP7_75t_L g117 ( 
.A(n_60),
.Y(n_117)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_46),
.Y(n_61)
);

OAI22xp33_ASAP7_75t_SL g62 ( 
.A1(n_40),
.A2(n_30),
.B1(n_33),
.B2(n_27),
.Y(n_62)
);

OAI22xp5_ASAP7_75t_SL g125 ( 
.A1(n_62),
.A2(n_72),
.B1(n_86),
.B2(n_31),
.Y(n_125)
);

CKINVDCx5p33_ASAP7_75t_R g63 ( 
.A(n_36),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_SL g121 ( 
.A(n_63),
.B(n_66),
.Y(n_121)
);

AOI22xp33_ASAP7_75t_L g64 ( 
.A1(n_47),
.A2(n_26),
.B1(n_33),
.B2(n_27),
.Y(n_64)
);

OAI22xp5_ASAP7_75t_L g103 ( 
.A1(n_64),
.A2(n_73),
.B1(n_90),
.B2(n_98),
.Y(n_103)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_36),
.Y(n_65)
);

BUFx3_ASAP7_75t_L g114 ( 
.A(n_65),
.Y(n_114)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_46),
.Y(n_66)
);

HB1xp67_ASAP7_75t_L g68 ( 
.A(n_42),
.Y(n_68)
);

CKINVDCx16_ASAP7_75t_R g104 ( 
.A(n_68),
.Y(n_104)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_43),
.Y(n_69)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_69),
.Y(n_102)
);

INVx4_ASAP7_75t_L g70 ( 
.A(n_42),
.Y(n_70)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_70),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_SL g71 ( 
.A(n_41),
.B(n_25),
.Y(n_71)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_71),
.Y(n_116)
);

AOI22xp5_ASAP7_75t_L g72 ( 
.A1(n_47),
.A2(n_30),
.B1(n_33),
.B2(n_27),
.Y(n_72)
);

AOI22xp33_ASAP7_75t_L g73 ( 
.A1(n_41),
.A2(n_26),
.B1(n_27),
.B2(n_29),
.Y(n_73)
);

HB1xp67_ASAP7_75t_L g74 ( 
.A(n_38),
.Y(n_74)
);

OR2x2_ASAP7_75t_L g108 ( 
.A(n_74),
.B(n_75),
.Y(n_108)
);

BUFx6f_ASAP7_75t_L g75 ( 
.A(n_38),
.Y(n_75)
);

BUFx12f_ASAP7_75t_L g76 ( 
.A(n_44),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_L g100 ( 
.A(n_76),
.B(n_78),
.Y(n_100)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_39),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_SL g107 ( 
.A(n_77),
.B(n_80),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_44),
.B(n_25),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_L g105 ( 
.A(n_79),
.B(n_82),
.Y(n_105)
);

INVx5_ASAP7_75t_L g80 ( 
.A(n_38),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_L g81 ( 
.A(n_35),
.B(n_22),
.Y(n_81)
);

INVxp67_ASAP7_75t_L g82 ( 
.A(n_39),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_44),
.B(n_15),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g111 ( 
.A(n_84),
.B(n_85),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_L g85 ( 
.A(n_37),
.B(n_15),
.Y(n_85)
);

OAI22xp5_ASAP7_75t_SL g86 ( 
.A1(n_37),
.A2(n_29),
.B1(n_23),
.B2(n_34),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_L g119 ( 
.A(n_87),
.B(n_88),
.Y(n_119)
);

BUFx6f_ASAP7_75t_L g88 ( 
.A(n_48),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_43),
.B(n_34),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g126 ( 
.A(n_89),
.B(n_92),
.Y(n_126)
);

OAI22xp5_ASAP7_75t_L g90 ( 
.A1(n_47),
.A2(n_23),
.B1(n_21),
.B2(n_28),
.Y(n_90)
);

AOI21xp5_ASAP7_75t_L g106 ( 
.A1(n_91),
.A2(n_97),
.B(n_99),
.Y(n_106)
);

INVx2_ASAP7_75t_L g92 ( 
.A(n_45),
.Y(n_92)
);

INVxp67_ASAP7_75t_L g93 ( 
.A(n_48),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_93),
.B(n_94),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_L g94 ( 
.A(n_46),
.B(n_28),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_SL g96 ( 
.A(n_43),
.B(n_21),
.Y(n_96)
);

XNOR2xp5_ASAP7_75t_L g113 ( 
.A(n_96),
.B(n_31),
.Y(n_113)
);

BUFx6f_ASAP7_75t_L g97 ( 
.A(n_48),
.Y(n_97)
);

OAI22xp5_ASAP7_75t_L g98 ( 
.A1(n_47),
.A2(n_16),
.B1(n_24),
.B2(n_18),
.Y(n_98)
);

INVx2_ASAP7_75t_L g99 ( 
.A(n_45),
.Y(n_99)
);

MAJIxp5_ASAP7_75t_L g101 ( 
.A(n_72),
.B(n_29),
.C(n_24),
.Y(n_101)
);

AND2x2_ASAP7_75t_L g134 ( 
.A(n_101),
.B(n_125),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_SL g137 ( 
.A(n_113),
.B(n_109),
.Y(n_137)
);

AO22x1_ASAP7_75t_SL g115 ( 
.A1(n_82),
.A2(n_24),
.B1(n_18),
.B2(n_4),
.Y(n_115)
);

OAI22xp5_ASAP7_75t_L g151 ( 
.A1(n_115),
.A2(n_124),
.B1(n_57),
.B2(n_92),
.Y(n_151)
);

XNOR2xp5_ASAP7_75t_L g123 ( 
.A(n_91),
.B(n_31),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_L g130 ( 
.A(n_123),
.B(n_51),
.Y(n_130)
);

AO22x1_ASAP7_75t_SL g124 ( 
.A1(n_52),
.A2(n_24),
.B1(n_18),
.B2(n_4),
.Y(n_124)
);

INVx2_ASAP7_75t_L g129 ( 
.A(n_114),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_L g169 ( 
.A(n_129),
.B(n_132),
.Y(n_169)
);

XNOR2xp5_ASAP7_75t_SL g187 ( 
.A(n_130),
.B(n_104),
.Y(n_187)
);

CKINVDCx20_ASAP7_75t_R g131 ( 
.A(n_112),
.Y(n_131)
);

CKINVDCx20_ASAP7_75t_R g185 ( 
.A(n_131),
.Y(n_185)
);

CKINVDCx14_ASAP7_75t_R g132 ( 
.A(n_118),
.Y(n_132)
);

INVx1_ASAP7_75t_SL g133 ( 
.A(n_107),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_L g170 ( 
.A(n_133),
.B(n_143),
.Y(n_170)
);

NOR2xp33_ASAP7_75t_SL g135 ( 
.A(n_109),
.B(n_87),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_SL g167 ( 
.A(n_135),
.B(n_147),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_L g136 ( 
.A(n_119),
.B(n_51),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_L g176 ( 
.A(n_136),
.B(n_155),
.Y(n_176)
);

XOR2xp5_ASAP7_75t_L g200 ( 
.A(n_137),
.B(n_6),
.Y(n_200)
);

AND2x2_ASAP7_75t_L g138 ( 
.A(n_123),
.B(n_86),
.Y(n_138)
);

AOI21xp5_ASAP7_75t_SL g171 ( 
.A1(n_138),
.A2(n_157),
.B(n_130),
.Y(n_171)
);

NOR2xp33_ASAP7_75t_L g139 ( 
.A(n_112),
.B(n_58),
.Y(n_139)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_139),
.Y(n_175)
);

NOR2xp33_ASAP7_75t_L g140 ( 
.A(n_107),
.B(n_59),
.Y(n_140)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_140),
.Y(n_183)
);

OAI22xp33_ASAP7_75t_L g141 ( 
.A1(n_115),
.A2(n_80),
.B1(n_54),
.B2(n_93),
.Y(n_141)
);

OAI22xp5_ASAP7_75t_L g188 ( 
.A1(n_141),
.A2(n_160),
.B1(n_128),
.B2(n_3),
.Y(n_188)
);

AO21x2_ASAP7_75t_L g142 ( 
.A1(n_115),
.A2(n_54),
.B(n_60),
.Y(n_142)
);

OA22x2_ASAP7_75t_L g193 ( 
.A1(n_142),
.A2(n_154),
.B1(n_76),
.B2(n_83),
.Y(n_193)
);

INVx2_ASAP7_75t_L g143 ( 
.A(n_114),
.Y(n_143)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_122),
.Y(n_144)
);

NOR2xp33_ASAP7_75t_L g174 ( 
.A(n_144),
.B(n_145),
.Y(n_174)
);

INVx2_ASAP7_75t_L g145 ( 
.A(n_118),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_SL g146 ( 
.A(n_109),
.B(n_67),
.Y(n_146)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_146),
.Y(n_189)
);

NOR2xp33_ASAP7_75t_SL g147 ( 
.A(n_116),
.B(n_50),
.Y(n_147)
);

INVx3_ASAP7_75t_L g148 ( 
.A(n_117),
.Y(n_148)
);

NOR2xp33_ASAP7_75t_L g180 ( 
.A(n_148),
.B(n_150),
.Y(n_180)
);

NOR2xp33_ASAP7_75t_SL g149 ( 
.A(n_116),
.B(n_70),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_SL g195 ( 
.A(n_149),
.B(n_153),
.Y(n_195)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_119),
.Y(n_150)
);

AOI22xp5_ASAP7_75t_L g190 ( 
.A1(n_151),
.A2(n_152),
.B1(n_162),
.B2(n_164),
.Y(n_190)
);

OAI22xp5_ASAP7_75t_L g152 ( 
.A1(n_101),
.A2(n_49),
.B1(n_99),
.B2(n_75),
.Y(n_152)
);

CKINVDCx16_ASAP7_75t_R g153 ( 
.A(n_110),
.Y(n_153)
);

OA22x2_ASAP7_75t_L g154 ( 
.A1(n_115),
.A2(n_124),
.B1(n_108),
.B2(n_125),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_L g155 ( 
.A(n_127),
.B(n_63),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_L g156 ( 
.A(n_117),
.B(n_97),
.Y(n_156)
);

NOR2xp33_ASAP7_75t_SL g179 ( 
.A(n_156),
.B(n_163),
.Y(n_179)
);

AND2x2_ASAP7_75t_L g157 ( 
.A(n_113),
.B(n_88),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_SL g158 ( 
.A(n_111),
.B(n_10),
.Y(n_158)
);

CKINVDCx16_ASAP7_75t_R g172 ( 
.A(n_158),
.Y(n_172)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_127),
.Y(n_159)
);

INVx13_ASAP7_75t_L g194 ( 
.A(n_159),
.Y(n_194)
);

AOI22xp33_ASAP7_75t_L g160 ( 
.A1(n_124),
.A2(n_95),
.B1(n_13),
.B2(n_11),
.Y(n_160)
);

CKINVDCx20_ASAP7_75t_R g161 ( 
.A(n_126),
.Y(n_161)
);

MAJIxp5_ASAP7_75t_SL g197 ( 
.A(n_161),
.B(n_2),
.C(n_5),
.Y(n_197)
);

OAI22xp5_ASAP7_75t_L g162 ( 
.A1(n_103),
.A2(n_124),
.B1(n_105),
.B2(n_106),
.Y(n_162)
);

NOR2xp33_ASAP7_75t_L g163 ( 
.A(n_104),
.B(n_95),
.Y(n_163)
);

OAI22xp5_ASAP7_75t_L g164 ( 
.A1(n_103),
.A2(n_76),
.B1(n_65),
.B2(n_83),
.Y(n_164)
);

INVx3_ASAP7_75t_L g165 ( 
.A(n_129),
.Y(n_165)
);

NOR2xp33_ASAP7_75t_L g209 ( 
.A(n_165),
.B(n_166),
.Y(n_209)
);

BUFx6f_ASAP7_75t_L g166 ( 
.A(n_143),
.Y(n_166)
);

INVx8_ASAP7_75t_L g168 ( 
.A(n_142),
.Y(n_168)
);

OAI21xp5_ASAP7_75t_L g218 ( 
.A1(n_171),
.A2(n_191),
.B(n_6),
.Y(n_218)
);

MAJIxp5_ASAP7_75t_L g173 ( 
.A(n_150),
.B(n_106),
.C(n_121),
.Y(n_173)
);

MAJIxp5_ASAP7_75t_L g204 ( 
.A(n_173),
.B(n_182),
.C(n_187),
.Y(n_204)
);

NAND2xp5_ASAP7_75t_L g177 ( 
.A(n_136),
.B(n_105),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_L g202 ( 
.A(n_177),
.B(n_178),
.Y(n_202)
);

OAI32xp33_ASAP7_75t_L g178 ( 
.A1(n_154),
.A2(n_108),
.A3(n_111),
.B1(n_126),
.B2(n_100),
.Y(n_178)
);

AOI21xp5_ASAP7_75t_L g181 ( 
.A1(n_154),
.A2(n_100),
.B(n_108),
.Y(n_181)
);

AOI21xp5_ASAP7_75t_L g201 ( 
.A1(n_181),
.A2(n_196),
.B(n_186),
.Y(n_201)
);

MAJIxp5_ASAP7_75t_L g182 ( 
.A(n_159),
.B(n_162),
.C(n_155),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_L g184 ( 
.A(n_133),
.B(n_120),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_L g206 ( 
.A(n_184),
.B(n_186),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_L g186 ( 
.A(n_138),
.B(n_102),
.Y(n_186)
);

AOI22xp5_ASAP7_75t_L g208 ( 
.A1(n_188),
.A2(n_193),
.B1(n_142),
.B2(n_152),
.Y(n_208)
);

OAI21xp33_ASAP7_75t_L g191 ( 
.A1(n_154),
.A2(n_2),
.B(n_5),
.Y(n_191)
);

XNOR2xp5_ASAP7_75t_L g192 ( 
.A(n_138),
.B(n_157),
.Y(n_192)
);

OAI21xp5_ASAP7_75t_L g196 ( 
.A1(n_135),
.A2(n_128),
.B(n_5),
.Y(n_196)
);

CKINVDCx20_ASAP7_75t_R g207 ( 
.A(n_197),
.Y(n_207)
);

XNOR2xp5_ASAP7_75t_SL g198 ( 
.A(n_157),
.B(n_5),
.Y(n_198)
);

MAJIxp5_ASAP7_75t_L g199 ( 
.A(n_161),
.B(n_6),
.C(n_7),
.Y(n_199)
);

MAJIxp5_ASAP7_75t_L g211 ( 
.A(n_200),
.B(n_149),
.C(n_147),
.Y(n_211)
);

AOI21xp5_ASAP7_75t_L g240 ( 
.A1(n_201),
.A2(n_210),
.B(n_218),
.Y(n_240)
);

INVx2_ASAP7_75t_SL g203 ( 
.A(n_193),
.Y(n_203)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_203),
.Y(n_225)
);

OAI22xp5_ASAP7_75t_L g205 ( 
.A1(n_190),
.A2(n_142),
.B1(n_151),
.B2(n_164),
.Y(n_205)
);

CKINVDCx16_ASAP7_75t_R g236 ( 
.A(n_205),
.Y(n_236)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_208),
.Y(n_227)
);

XOR2xp5_ASAP7_75t_SL g210 ( 
.A(n_181),
.B(n_134),
.Y(n_210)
);

XNOR2xp5_ASAP7_75t_L g241 ( 
.A(n_211),
.B(n_220),
.Y(n_241)
);

NAND2xp5_ASAP7_75t_L g212 ( 
.A(n_176),
.B(n_134),
.Y(n_212)
);

NAND2xp5_ASAP7_75t_L g242 ( 
.A(n_212),
.B(n_214),
.Y(n_242)
);

NAND3xp33_ASAP7_75t_L g213 ( 
.A(n_198),
.B(n_142),
.C(n_134),
.Y(n_213)
);

AOI22xp5_ASAP7_75t_SL g237 ( 
.A1(n_213),
.A2(n_165),
.B1(n_166),
.B2(n_219),
.Y(n_237)
);

NAND2xp5_ASAP7_75t_SL g214 ( 
.A(n_177),
.B(n_144),
.Y(n_214)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_180),
.Y(n_215)
);

NAND2xp5_ASAP7_75t_L g243 ( 
.A(n_215),
.B(n_216),
.Y(n_243)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_174),
.Y(n_216)
);

NAND2xp5_ASAP7_75t_SL g217 ( 
.A(n_184),
.B(n_141),
.Y(n_217)
);

NAND2xp5_ASAP7_75t_L g246 ( 
.A(n_217),
.B(n_219),
.Y(n_246)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_176),
.Y(n_219)
);

AOI21xp5_ASAP7_75t_L g220 ( 
.A1(n_193),
.A2(n_145),
.B(n_148),
.Y(n_220)
);

AOI322xp5_ASAP7_75t_L g221 ( 
.A1(n_193),
.A2(n_8),
.A3(n_9),
.B1(n_191),
.B2(n_171),
.C1(n_192),
.C2(n_178),
.Y(n_221)
);

AOI322xp5_ASAP7_75t_L g231 ( 
.A1(n_221),
.A2(n_196),
.A3(n_167),
.B1(n_189),
.B2(n_195),
.C1(n_197),
.C2(n_185),
.Y(n_231)
);

NAND2xp5_ASAP7_75t_L g222 ( 
.A(n_182),
.B(n_8),
.Y(n_222)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_222),
.Y(n_228)
);

NAND2xp5_ASAP7_75t_SL g223 ( 
.A(n_183),
.B(n_8),
.Y(n_223)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_223),
.Y(n_233)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_170),
.Y(n_224)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_224),
.Y(n_234)
);

CKINVDCx20_ASAP7_75t_R g226 ( 
.A(n_209),
.Y(n_226)
);

NAND2xp5_ASAP7_75t_L g248 ( 
.A(n_226),
.B(n_216),
.Y(n_248)
);

MAJIxp5_ASAP7_75t_L g229 ( 
.A(n_204),
.B(n_187),
.C(n_173),
.Y(n_229)
);

MAJIxp5_ASAP7_75t_L g257 ( 
.A(n_229),
.B(n_230),
.C(n_232),
.Y(n_257)
);

MAJIxp5_ASAP7_75t_L g230 ( 
.A(n_204),
.B(n_190),
.C(n_200),
.Y(n_230)
);

XNOR2xp5_ASAP7_75t_SL g250 ( 
.A(n_231),
.B(n_222),
.Y(n_250)
);

MAJIxp5_ASAP7_75t_L g232 ( 
.A(n_212),
.B(n_194),
.C(n_199),
.Y(n_232)
);

AOI322xp5_ASAP7_75t_L g235 ( 
.A1(n_210),
.A2(n_168),
.A3(n_179),
.B1(n_175),
.B2(n_194),
.C1(n_172),
.C2(n_169),
.Y(n_235)
);

XNOR2xp5_ASAP7_75t_L g261 ( 
.A(n_235),
.B(n_232),
.Y(n_261)
);

XOR2xp5_ASAP7_75t_L g252 ( 
.A(n_237),
.B(n_239),
.Y(n_252)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_209),
.Y(n_238)
);

NOR2xp33_ASAP7_75t_L g247 ( 
.A(n_238),
.B(n_244),
.Y(n_247)
);

XOR2xp5_ASAP7_75t_L g239 ( 
.A(n_210),
.B(n_202),
.Y(n_239)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_214),
.Y(n_244)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_206),
.Y(n_245)
);

NOR2xp33_ASAP7_75t_L g258 ( 
.A(n_245),
.B(n_246),
.Y(n_258)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_248),
.Y(n_272)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_243),
.Y(n_249)
);

NAND2xp5_ASAP7_75t_SL g264 ( 
.A(n_249),
.B(n_260),
.Y(n_264)
);

XNOR2xp5_ASAP7_75t_L g276 ( 
.A(n_250),
.B(n_230),
.Y(n_276)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_242),
.Y(n_251)
);

NOR2xp33_ASAP7_75t_L g268 ( 
.A(n_251),
.B(n_261),
.Y(n_268)
);

NAND2xp5_ASAP7_75t_L g253 ( 
.A(n_244),
.B(n_206),
.Y(n_253)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_253),
.Y(n_271)
);

NAND2xp5_ASAP7_75t_L g254 ( 
.A(n_245),
.B(n_202),
.Y(n_254)
);

OAI21xp5_ASAP7_75t_L g275 ( 
.A1(n_254),
.A2(n_255),
.B(n_256),
.Y(n_275)
);

NAND2xp5_ASAP7_75t_L g255 ( 
.A(n_242),
.B(n_207),
.Y(n_255)
);

NAND2xp5_ASAP7_75t_L g256 ( 
.A(n_246),
.B(n_207),
.Y(n_256)
);

CKINVDCx14_ASAP7_75t_R g267 ( 
.A(n_258),
.Y(n_267)
);

XOR2xp5_ASAP7_75t_L g259 ( 
.A(n_239),
.B(n_201),
.Y(n_259)
);

XOR2xp5_ASAP7_75t_L g266 ( 
.A(n_259),
.B(n_240),
.Y(n_266)
);

NOR2xp33_ASAP7_75t_L g260 ( 
.A(n_226),
.B(n_215),
.Y(n_260)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_243),
.Y(n_262)
);

NAND2xp5_ASAP7_75t_SL g270 ( 
.A(n_262),
.B(n_263),
.Y(n_270)
);

INVx13_ASAP7_75t_L g263 ( 
.A(n_238),
.Y(n_263)
);

OAI22xp33_ASAP7_75t_SL g265 ( 
.A1(n_262),
.A2(n_227),
.B1(n_236),
.B2(n_225),
.Y(n_265)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_265),
.Y(n_286)
);

MAJIxp5_ASAP7_75t_L g287 ( 
.A(n_266),
.B(n_257),
.C(n_259),
.Y(n_287)
);

AOI22xp5_ASAP7_75t_L g269 ( 
.A1(n_256),
.A2(n_227),
.B1(n_205),
.B2(n_203),
.Y(n_269)
);

AOI22xp5_ASAP7_75t_L g282 ( 
.A1(n_269),
.A2(n_273),
.B1(n_274),
.B2(n_253),
.Y(n_282)
);

AOI22xp5_ASAP7_75t_L g273 ( 
.A1(n_251),
.A2(n_203),
.B1(n_225),
.B2(n_218),
.Y(n_273)
);

AOI22xp5_ASAP7_75t_L g274 ( 
.A1(n_255),
.A2(n_237),
.B1(n_217),
.B2(n_213),
.Y(n_274)
);

NOR2xp33_ASAP7_75t_L g280 ( 
.A(n_276),
.B(n_257),
.Y(n_280)
);

INVx1_ASAP7_75t_SL g277 ( 
.A(n_267),
.Y(n_277)
);

NAND2xp5_ASAP7_75t_L g295 ( 
.A(n_277),
.B(n_281),
.Y(n_295)
);

NAND2xp5_ASAP7_75t_L g278 ( 
.A(n_270),
.B(n_234),
.Y(n_278)
);

OAI21xp5_ASAP7_75t_SL g288 ( 
.A1(n_278),
.A2(n_279),
.B(n_283),
.Y(n_288)
);

NAND2xp5_ASAP7_75t_L g279 ( 
.A(n_264),
.B(n_234),
.Y(n_279)
);

MAJIxp5_ASAP7_75t_L g291 ( 
.A(n_280),
.B(n_252),
.C(n_268),
.Y(n_291)
);

NOR2xp33_ASAP7_75t_L g281 ( 
.A(n_272),
.B(n_263),
.Y(n_281)
);

OAI22xp5_ASAP7_75t_L g289 ( 
.A1(n_282),
.A2(n_284),
.B1(n_269),
.B2(n_273),
.Y(n_289)
);

NAND2xp5_ASAP7_75t_SL g283 ( 
.A(n_275),
.B(n_224),
.Y(n_283)
);

AOI21xp5_ASAP7_75t_L g284 ( 
.A1(n_272),
.A2(n_247),
.B(n_248),
.Y(n_284)
);

NOR2xp33_ASAP7_75t_L g285 ( 
.A(n_275),
.B(n_228),
.Y(n_285)
);

NOR2xp33_ASAP7_75t_SL g293 ( 
.A(n_285),
.B(n_233),
.Y(n_293)
);

NAND2xp5_ASAP7_75t_SL g298 ( 
.A(n_289),
.B(n_292),
.Y(n_298)
);

MAJIxp5_ASAP7_75t_L g290 ( 
.A(n_287),
.B(n_229),
.C(n_266),
.Y(n_290)
);

NOR2xp33_ASAP7_75t_L g297 ( 
.A(n_290),
.B(n_291),
.Y(n_297)
);

NOR2xp67_ASAP7_75t_L g292 ( 
.A(n_284),
.B(n_250),
.Y(n_292)
);

NOR2xp33_ASAP7_75t_L g299 ( 
.A(n_293),
.B(n_294),
.Y(n_299)
);

MAJIxp5_ASAP7_75t_L g294 ( 
.A(n_282),
.B(n_271),
.C(n_228),
.Y(n_294)
);

OAI22xp5_ASAP7_75t_SL g296 ( 
.A1(n_294),
.A2(n_286),
.B1(n_274),
.B2(n_254),
.Y(n_296)
);

OAI22xp5_ASAP7_75t_L g302 ( 
.A1(n_296),
.A2(n_240),
.B1(n_221),
.B2(n_241),
.Y(n_302)
);

NOR2xp33_ASAP7_75t_L g300 ( 
.A(n_295),
.B(n_233),
.Y(n_300)
);

NAND2xp5_ASAP7_75t_L g303 ( 
.A(n_300),
.B(n_277),
.Y(n_303)
);

OAI21xp5_ASAP7_75t_L g301 ( 
.A1(n_298),
.A2(n_288),
.B(n_290),
.Y(n_301)
);

MAJIxp5_ASAP7_75t_L g305 ( 
.A(n_301),
.B(n_303),
.C(n_304),
.Y(n_305)
);

XOR2xp5_ASAP7_75t_L g306 ( 
.A(n_302),
.B(n_296),
.Y(n_306)
);

OAI22xp5_ASAP7_75t_L g304 ( 
.A1(n_299),
.A2(n_208),
.B1(n_220),
.B2(n_241),
.Y(n_304)
);

NAND2xp5_ASAP7_75t_L g307 ( 
.A(n_306),
.B(n_297),
.Y(n_307)
);

XOR2xp5_ASAP7_75t_L g308 ( 
.A(n_307),
.B(n_305),
.Y(n_308)
);


endmodule