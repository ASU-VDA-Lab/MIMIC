module fake_netlist_5_2083_n_757 (n_137, n_91, n_82, n_122, n_142, n_10, n_140, n_24, n_124, n_86, n_136, n_146, n_143, n_83, n_132, n_61, n_90, n_127, n_75, n_101, n_65, n_78, n_74, n_144, n_114, n_57, n_96, n_37, n_111, n_108, n_129, n_31, n_13, n_66, n_98, n_60, n_16, n_43, n_107, n_0, n_58, n_9, n_69, n_18, n_116, n_42, n_22, n_1, n_45, n_117, n_46, n_21, n_94, n_113, n_38, n_123, n_139, n_105, n_80, n_4, n_125, n_35, n_128, n_73, n_17, n_92, n_19, n_149, n_120, n_135, n_30, n_5, n_33, n_126, n_14, n_84, n_23, n_130, n_29, n_79, n_131, n_151, n_47, n_25, n_53, n_8, n_44, n_40, n_34, n_100, n_62, n_138, n_148, n_71, n_109, n_112, n_85, n_95, n_119, n_59, n_26, n_133, n_55, n_99, n_2, n_3, n_49, n_20, n_6, n_39, n_54, n_147, n_12, n_67, n_121, n_36, n_76, n_87, n_150, n_27, n_64, n_77, n_102, n_106, n_81, n_118, n_28, n_89, n_70, n_115, n_68, n_93, n_72, n_134, n_32, n_41, n_104, n_103, n_56, n_51, n_63, n_97, n_141, n_11, n_7, n_15, n_145, n_48, n_50, n_52, n_88, n_110, n_757);

input n_137;
input n_91;
input n_82;
input n_122;
input n_142;
input n_10;
input n_140;
input n_24;
input n_124;
input n_86;
input n_136;
input n_146;
input n_143;
input n_83;
input n_132;
input n_61;
input n_90;
input n_127;
input n_75;
input n_101;
input n_65;
input n_78;
input n_74;
input n_144;
input n_114;
input n_57;
input n_96;
input n_37;
input n_111;
input n_108;
input n_129;
input n_31;
input n_13;
input n_66;
input n_98;
input n_60;
input n_16;
input n_43;
input n_107;
input n_0;
input n_58;
input n_9;
input n_69;
input n_18;
input n_116;
input n_42;
input n_22;
input n_1;
input n_45;
input n_117;
input n_46;
input n_21;
input n_94;
input n_113;
input n_38;
input n_123;
input n_139;
input n_105;
input n_80;
input n_4;
input n_125;
input n_35;
input n_128;
input n_73;
input n_17;
input n_92;
input n_19;
input n_149;
input n_120;
input n_135;
input n_30;
input n_5;
input n_33;
input n_126;
input n_14;
input n_84;
input n_23;
input n_130;
input n_29;
input n_79;
input n_131;
input n_151;
input n_47;
input n_25;
input n_53;
input n_8;
input n_44;
input n_40;
input n_34;
input n_100;
input n_62;
input n_138;
input n_148;
input n_71;
input n_109;
input n_112;
input n_85;
input n_95;
input n_119;
input n_59;
input n_26;
input n_133;
input n_55;
input n_99;
input n_2;
input n_3;
input n_49;
input n_20;
input n_6;
input n_39;
input n_54;
input n_147;
input n_12;
input n_67;
input n_121;
input n_36;
input n_76;
input n_87;
input n_150;
input n_27;
input n_64;
input n_77;
input n_102;
input n_106;
input n_81;
input n_118;
input n_28;
input n_89;
input n_70;
input n_115;
input n_68;
input n_93;
input n_72;
input n_134;
input n_32;
input n_41;
input n_104;
input n_103;
input n_56;
input n_51;
input n_63;
input n_97;
input n_141;
input n_11;
input n_7;
input n_15;
input n_145;
input n_48;
input n_50;
input n_52;
input n_88;
input n_110;

output n_757;

wire n_676;
wire n_294;
wire n_431;
wire n_318;
wire n_419;
wire n_380;
wire n_653;
wire n_611;
wire n_444;
wire n_642;
wire n_469;
wire n_615;
wire n_194;
wire n_316;
wire n_389;
wire n_549;
wire n_684;
wire n_418;
wire n_248;
wire n_315;
wire n_268;
wire n_523;
wire n_451;
wire n_532;
wire n_705;
wire n_619;
wire n_408;
wire n_678;
wire n_664;
wire n_376;
wire n_697;
wire n_503;
wire n_235;
wire n_226;
wire n_605;
wire n_667;
wire n_515;
wire n_353;
wire n_351;
wire n_367;
wire n_620;
wire n_643;
wire n_452;
wire n_397;
wire n_525;
wire n_493;
wire n_703;
wire n_698;
wire n_483;
wire n_544;
wire n_683;
wire n_155;
wire n_649;
wire n_552;
wire n_547;
wire n_721;
wire n_467;
wire n_564;
wire n_423;
wire n_284;
wire n_245;
wire n_501;
wire n_725;
wire n_280;
wire n_744;
wire n_590;
wire n_629;
wire n_672;
wire n_378;
wire n_551;
wire n_688;
wire n_581;
wire n_382;
wire n_554;
wire n_254;
wire n_690;
wire n_583;
wire n_671;
wire n_718;
wire n_302;
wire n_265;
wire n_526;
wire n_719;
wire n_293;
wire n_372;
wire n_443;
wire n_244;
wire n_677;
wire n_173;
wire n_198;
wire n_714;
wire n_447;
wire n_247;
wire n_314;
wire n_368;
wire n_433;
wire n_604;
wire n_321;
wire n_292;
wire n_625;
wire n_621;
wire n_753;
wire n_455;
wire n_674;
wire n_417;
wire n_612;
wire n_212;
wire n_385;
wire n_516;
wire n_498;
wire n_507;
wire n_497;
wire n_689;
wire n_738;
wire n_606;
wire n_559;
wire n_275;
wire n_640;
wire n_252;
wire n_624;
wire n_295;
wire n_330;
wire n_508;
wire n_739;
wire n_506;
wire n_737;
wire n_610;
wire n_692;
wire n_755;
wire n_568;
wire n_509;
wire n_373;
wire n_307;
wire n_633;
wire n_439;
wire n_530;
wire n_556;
wire n_209;
wire n_259;
wire n_448;
wire n_668;
wire n_733;
wire n_375;
wire n_301;
wire n_576;
wire n_186;
wire n_537;
wire n_191;
wire n_587;
wire n_659;
wire n_492;
wire n_563;
wire n_171;
wire n_153;
wire n_756;
wire n_524;
wire n_399;
wire n_341;
wire n_204;
wire n_394;
wire n_250;
wire n_579;
wire n_741;
wire n_548;
wire n_543;
wire n_260;
wire n_298;
wire n_650;
wire n_320;
wire n_694;
wire n_518;
wire n_505;
wire n_286;
wire n_282;
wire n_752;
wire n_331;
wire n_406;
wire n_519;
wire n_470;
wire n_325;
wire n_449;
wire n_724;
wire n_546;
wire n_658;
wire n_281;
wire n_240;
wire n_381;
wire n_189;
wire n_220;
wire n_291;
wire n_231;
wire n_257;
wire n_390;
wire n_731;
wire n_456;
wire n_371;
wire n_481;
wire n_535;
wire n_709;
wire n_152;
wire n_540;
wire n_317;
wire n_618;
wire n_323;
wire n_569;
wire n_195;
wire n_356;
wire n_227;
wire n_592;
wire n_271;
wire n_335;
wire n_654;
wire n_370;
wire n_167;
wire n_234;
wire n_343;
wire n_308;
wire n_379;
wire n_428;
wire n_267;
wire n_514;
wire n_457;
wire n_570;
wire n_297;
wire n_156;
wire n_603;
wire n_225;
wire n_377;
wire n_751;
wire n_484;
wire n_219;
wire n_442;
wire n_157;
wire n_192;
wire n_636;
wire n_600;
wire n_660;
wire n_223;
wire n_392;
wire n_158;
wire n_655;
wire n_704;
wire n_264;
wire n_669;
wire n_472;
wire n_742;
wire n_750;
wire n_454;
wire n_387;
wire n_374;
wire n_163;
wire n_276;
wire n_339;
wire n_183;
wire n_185;
wire n_243;
wire n_398;
wire n_396;
wire n_635;
wire n_347;
wire n_169;
wire n_522;
wire n_550;
wire n_255;
wire n_696;
wire n_215;
wire n_350;
wire n_196;
wire n_662;
wire n_459;
wire n_646;
wire n_211;
wire n_218;
wire n_400;
wire n_181;
wire n_436;
wire n_290;
wire n_580;
wire n_221;
wire n_178;
wire n_622;
wire n_723;
wire n_386;
wire n_578;
wire n_287;
wire n_344;
wire n_555;
wire n_473;
wire n_422;
wire n_475;
wire n_661;
wire n_682;
wire n_415;
wire n_485;
wire n_496;
wire n_355;
wire n_486;
wire n_670;
wire n_336;
wire n_584;
wire n_681;
wire n_591;
wire n_521;
wire n_614;
wire n_663;
wire n_337;
wire n_430;
wire n_313;
wire n_673;
wire n_631;
wire n_479;
wire n_528;
wire n_510;
wire n_216;
wire n_680;
wire n_168;
wire n_395;
wire n_164;
wire n_432;
wire n_553;
wire n_727;
wire n_311;
wire n_208;
wire n_743;
wire n_214;
wire n_328;
wire n_299;
wire n_303;
wire n_369;
wire n_675;
wire n_296;
wire n_613;
wire n_241;
wire n_637;
wire n_357;
wire n_598;
wire n_685;
wire n_608;
wire n_184;
wire n_446;
wire n_445;
wire n_749;
wire n_691;
wire n_717;
wire n_165;
wire n_468;
wire n_499;
wire n_213;
wire n_342;
wire n_482;
wire n_517;
wire n_588;
wire n_361;
wire n_464;
wire n_363;
wire n_413;
wire n_402;
wire n_734;
wire n_638;
wire n_700;
wire n_197;
wire n_573;
wire n_236;
wire n_388;
wire n_249;
wire n_740;
wire n_304;
wire n_329;
wire n_203;
wire n_274;
wire n_577;
wire n_384;
wire n_582;
wire n_460;
wire n_277;
wire n_338;
wire n_477;
wire n_461;
wire n_333;
wire n_571;
wire n_693;
wire n_309;
wire n_512;
wire n_462;
wire n_322;
wire n_567;
wire n_258;
wire n_652;
wire n_306;
wire n_722;
wire n_458;
wire n_288;
wire n_188;
wire n_190;
wire n_201;
wire n_263;
wire n_471;
wire n_609;
wire n_224;
wire n_228;
wire n_283;
wire n_383;
wire n_711;
wire n_474;
wire n_542;
wire n_463;
wire n_488;
wire n_595;
wire n_736;
wire n_502;
wire n_239;
wire n_466;
wire n_420;
wire n_630;
wire n_489;
wire n_632;
wire n_699;
wire n_617;
wire n_310;
wire n_593;
wire n_504;
wire n_511;
wire n_748;
wire n_586;
wire n_465;
wire n_358;
wire n_362;
wire n_170;
wire n_332;
wire n_161;
wire n_273;
wire n_349;
wire n_585;
wire n_270;
wire n_616;
wire n_230;
wire n_601;
wire n_279;
wire n_253;
wire n_261;
wire n_174;
wire n_289;
wire n_745;
wire n_627;
wire n_172;
wire n_206;
wire n_217;
wire n_440;
wire n_726;
wire n_478;
wire n_545;
wire n_441;
wire n_450;
wire n_648;
wire n_312;
wire n_476;
wire n_429;
wire n_534;
wire n_345;
wire n_210;
wire n_494;
wire n_641;
wire n_628;
wire n_365;
wire n_729;
wire n_730;
wire n_176;
wire n_557;
wire n_182;
wire n_354;
wire n_575;
wire n_607;
wire n_480;
wire n_647;
wire n_237;
wire n_425;
wire n_513;
wire n_407;
wire n_527;
wire n_679;
wire n_707;
wire n_710;
wire n_695;
wire n_180;
wire n_560;
wire n_656;
wire n_340;
wire n_207;
wire n_561;
wire n_346;
wire n_393;
wire n_229;
wire n_495;
wire n_487;
wire n_602;
wire n_665;
wire n_574;
wire n_437;
wire n_177;
wire n_403;
wire n_453;
wire n_421;
wire n_720;
wire n_623;
wire n_405;
wire n_359;
wire n_490;
wire n_326;
wire n_233;
wire n_404;
wire n_686;
wire n_205;
wire n_366;
wire n_572;
wire n_712;
wire n_754;
wire n_246;
wire n_596;
wire n_179;
wire n_410;
wire n_558;
wire n_708;
wire n_269;
wire n_529;
wire n_735;
wire n_702;
wire n_285;
wire n_412;
wire n_232;
wire n_327;
wire n_657;
wire n_644;
wire n_728;
wire n_202;
wire n_266;
wire n_272;
wire n_491;
wire n_427;
wire n_732;
wire n_193;
wire n_251;
wire n_352;
wire n_160;
wire n_565;
wire n_426;
wire n_520;
wire n_566;
wire n_409;
wire n_589;
wire n_716;
wire n_597;
wire n_500;
wire n_562;
wire n_154;
wire n_300;
wire n_651;
wire n_435;
wire n_159;
wire n_334;
wire n_599;
wire n_541;
wire n_391;
wire n_701;
wire n_434;
wire n_645;
wire n_539;
wire n_175;
wire n_538;
wire n_666;
wire n_262;
wire n_238;
wire n_639;
wire n_687;
wire n_715;
wire n_411;
wire n_414;
wire n_319;
wire n_364;
wire n_536;
wire n_531;
wire n_242;
wire n_360;
wire n_594;
wire n_200;
wire n_162;
wire n_222;
wire n_438;
wire n_713;
wire n_324;
wire n_634;
wire n_416;
wire n_199;
wire n_187;
wire n_401;
wire n_348;
wire n_166;
wire n_626;
wire n_424;
wire n_706;
wire n_746;
wire n_256;
wire n_305;
wire n_533;
wire n_747;
wire n_278;

BUFx3_ASAP7_75t_L g152 ( 
.A(n_68),
.Y(n_152)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_44),
.Y(n_153)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_69),
.Y(n_154)
);

CKINVDCx5p33_ASAP7_75t_R g155 ( 
.A(n_122),
.Y(n_155)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_0),
.Y(n_156)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_105),
.Y(n_157)
);

HB1xp67_ASAP7_75t_L g158 ( 
.A(n_58),
.Y(n_158)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_85),
.Y(n_159)
);

CKINVDCx20_ASAP7_75t_R g160 ( 
.A(n_118),
.Y(n_160)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_99),
.Y(n_161)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_48),
.Y(n_162)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_127),
.Y(n_163)
);

CKINVDCx5p33_ASAP7_75t_R g164 ( 
.A(n_40),
.Y(n_164)
);

CKINVDCx5p33_ASAP7_75t_R g165 ( 
.A(n_106),
.Y(n_165)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_43),
.Y(n_166)
);

BUFx5_ASAP7_75t_L g167 ( 
.A(n_72),
.Y(n_167)
);

CKINVDCx5p33_ASAP7_75t_R g168 ( 
.A(n_28),
.Y(n_168)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_67),
.Y(n_169)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_146),
.Y(n_170)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_148),
.Y(n_171)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_98),
.Y(n_172)
);

CKINVDCx5p33_ASAP7_75t_R g173 ( 
.A(n_60),
.Y(n_173)
);

CKINVDCx5p33_ASAP7_75t_R g174 ( 
.A(n_83),
.Y(n_174)
);

INVx2_ASAP7_75t_L g175 ( 
.A(n_59),
.Y(n_175)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_41),
.Y(n_176)
);

CKINVDCx5p33_ASAP7_75t_R g177 ( 
.A(n_22),
.Y(n_177)
);

CKINVDCx20_ASAP7_75t_R g178 ( 
.A(n_75),
.Y(n_178)
);

CKINVDCx5p33_ASAP7_75t_R g179 ( 
.A(n_120),
.Y(n_179)
);

CKINVDCx5p33_ASAP7_75t_R g180 ( 
.A(n_24),
.Y(n_180)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_128),
.Y(n_181)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_23),
.Y(n_182)
);

INVx2_ASAP7_75t_L g183 ( 
.A(n_130),
.Y(n_183)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_91),
.Y(n_184)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_143),
.Y(n_185)
);

CKINVDCx5p33_ASAP7_75t_R g186 ( 
.A(n_136),
.Y(n_186)
);

CKINVDCx5p33_ASAP7_75t_R g187 ( 
.A(n_13),
.Y(n_187)
);

BUFx3_ASAP7_75t_L g188 ( 
.A(n_33),
.Y(n_188)
);

CKINVDCx5p33_ASAP7_75t_R g189 ( 
.A(n_151),
.Y(n_189)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_117),
.Y(n_190)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_129),
.Y(n_191)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_78),
.Y(n_192)
);

CKINVDCx5p33_ASAP7_75t_R g193 ( 
.A(n_45),
.Y(n_193)
);

BUFx6f_ASAP7_75t_L g194 ( 
.A(n_124),
.Y(n_194)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_81),
.Y(n_195)
);

INVx3_ASAP7_75t_L g196 ( 
.A(n_31),
.Y(n_196)
);

CKINVDCx5p33_ASAP7_75t_R g197 ( 
.A(n_11),
.Y(n_197)
);

INVx2_ASAP7_75t_SL g198 ( 
.A(n_14),
.Y(n_198)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_84),
.Y(n_199)
);

CKINVDCx16_ASAP7_75t_R g200 ( 
.A(n_116),
.Y(n_200)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_61),
.Y(n_201)
);

HB1xp67_ASAP7_75t_L g202 ( 
.A(n_19),
.Y(n_202)
);

CKINVDCx5p33_ASAP7_75t_R g203 ( 
.A(n_39),
.Y(n_203)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_55),
.Y(n_204)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_4),
.Y(n_205)
);

CKINVDCx5p33_ASAP7_75t_R g206 ( 
.A(n_88),
.Y(n_206)
);

CKINVDCx6p67_ASAP7_75t_R g207 ( 
.A(n_200),
.Y(n_207)
);

BUFx6f_ASAP7_75t_L g208 ( 
.A(n_194),
.Y(n_208)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_156),
.Y(n_209)
);

INVxp67_ASAP7_75t_L g210 ( 
.A(n_205),
.Y(n_210)
);

AND2x4_ASAP7_75t_L g211 ( 
.A(n_152),
.B(n_20),
.Y(n_211)
);

INVx2_ASAP7_75t_L g212 ( 
.A(n_167),
.Y(n_212)
);

NAND2xp5_ASAP7_75t_SL g213 ( 
.A(n_198),
.B(n_0),
.Y(n_213)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_152),
.Y(n_214)
);

BUFx6f_ASAP7_75t_L g215 ( 
.A(n_194),
.Y(n_215)
);

NAND2xp5_ASAP7_75t_L g216 ( 
.A(n_196),
.B(n_1),
.Y(n_216)
);

BUFx6f_ASAP7_75t_L g217 ( 
.A(n_194),
.Y(n_217)
);

BUFx6f_ASAP7_75t_L g218 ( 
.A(n_194),
.Y(n_218)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_188),
.Y(n_219)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_188),
.Y(n_220)
);

INVxp33_ASAP7_75t_SL g221 ( 
.A(n_158),
.Y(n_221)
);

BUFx6f_ASAP7_75t_L g222 ( 
.A(n_175),
.Y(n_222)
);

AND2x4_ASAP7_75t_L g223 ( 
.A(n_196),
.B(n_21),
.Y(n_223)
);

INVx2_ASAP7_75t_L g224 ( 
.A(n_167),
.Y(n_224)
);

CKINVDCx5p33_ASAP7_75t_R g225 ( 
.A(n_187),
.Y(n_225)
);

AND2x2_ASAP7_75t_L g226 ( 
.A(n_202),
.B(n_197),
.Y(n_226)
);

INVx2_ASAP7_75t_L g227 ( 
.A(n_167),
.Y(n_227)
);

BUFx6f_ASAP7_75t_L g228 ( 
.A(n_175),
.Y(n_228)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_153),
.Y(n_229)
);

INVx5_ASAP7_75t_L g230 ( 
.A(n_183),
.Y(n_230)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_154),
.Y(n_231)
);

INVx2_ASAP7_75t_L g232 ( 
.A(n_167),
.Y(n_232)
);

INVx2_ASAP7_75t_L g233 ( 
.A(n_167),
.Y(n_233)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_157),
.Y(n_234)
);

CKINVDCx5p33_ASAP7_75t_R g235 ( 
.A(n_155),
.Y(n_235)
);

BUFx6f_ASAP7_75t_L g236 ( 
.A(n_183),
.Y(n_236)
);

BUFx6f_ASAP7_75t_L g237 ( 
.A(n_159),
.Y(n_237)
);

HB1xp67_ASAP7_75t_L g238 ( 
.A(n_161),
.Y(n_238)
);

AND2x4_ASAP7_75t_L g239 ( 
.A(n_162),
.B(n_25),
.Y(n_239)
);

BUFx6f_ASAP7_75t_L g240 ( 
.A(n_163),
.Y(n_240)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_166),
.Y(n_241)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_169),
.Y(n_242)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_170),
.Y(n_243)
);

BUFx6f_ASAP7_75t_L g244 ( 
.A(n_171),
.Y(n_244)
);

BUFx6f_ASAP7_75t_L g245 ( 
.A(n_172),
.Y(n_245)
);

BUFx6f_ASAP7_75t_L g246 ( 
.A(n_176),
.Y(n_246)
);

CKINVDCx16_ASAP7_75t_R g247 ( 
.A(n_160),
.Y(n_247)
);

INVx3_ASAP7_75t_L g248 ( 
.A(n_180),
.Y(n_248)
);

INVx2_ASAP7_75t_L g249 ( 
.A(n_167),
.Y(n_249)
);

NAND2xp5_ASAP7_75t_L g250 ( 
.A(n_235),
.B(n_181),
.Y(n_250)
);

INVxp33_ASAP7_75t_L g251 ( 
.A(n_226),
.Y(n_251)
);

NAND2xp5_ASAP7_75t_SL g252 ( 
.A(n_221),
.B(n_225),
.Y(n_252)
);

INVx2_ASAP7_75t_L g253 ( 
.A(n_222),
.Y(n_253)
);

NAND3xp33_ASAP7_75t_L g254 ( 
.A(n_216),
.B(n_203),
.C(n_180),
.Y(n_254)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_222),
.Y(n_255)
);

NAND2xp5_ASAP7_75t_SL g256 ( 
.A(n_221),
.B(n_225),
.Y(n_256)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_222),
.Y(n_257)
);

INVx2_ASAP7_75t_L g258 ( 
.A(n_222),
.Y(n_258)
);

INVx2_ASAP7_75t_L g259 ( 
.A(n_228),
.Y(n_259)
);

NOR2xp33_ASAP7_75t_L g260 ( 
.A(n_248),
.B(n_203),
.Y(n_260)
);

OR2x6_ASAP7_75t_L g261 ( 
.A(n_213),
.B(n_182),
.Y(n_261)
);

INVx3_ASAP7_75t_L g262 ( 
.A(n_208),
.Y(n_262)
);

INVx2_ASAP7_75t_L g263 ( 
.A(n_228),
.Y(n_263)
);

AO21x2_ASAP7_75t_L g264 ( 
.A1(n_213),
.A2(n_184),
.B(n_204),
.Y(n_264)
);

INVx2_ASAP7_75t_L g265 ( 
.A(n_228),
.Y(n_265)
);

NOR2x1p5_ASAP7_75t_L g266 ( 
.A(n_207),
.B(n_206),
.Y(n_266)
);

INVx3_ASAP7_75t_L g267 ( 
.A(n_208),
.Y(n_267)
);

INVx2_ASAP7_75t_L g268 ( 
.A(n_228),
.Y(n_268)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_236),
.Y(n_269)
);

INVx2_ASAP7_75t_L g270 ( 
.A(n_236),
.Y(n_270)
);

INVx2_ASAP7_75t_L g271 ( 
.A(n_236),
.Y(n_271)
);

NAND2xp5_ASAP7_75t_L g272 ( 
.A(n_248),
.B(n_185),
.Y(n_272)
);

CKINVDCx16_ASAP7_75t_R g273 ( 
.A(n_247),
.Y(n_273)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_236),
.Y(n_274)
);

INVx2_ASAP7_75t_L g275 ( 
.A(n_208),
.Y(n_275)
);

NAND2xp5_ASAP7_75t_SL g276 ( 
.A(n_223),
.B(n_160),
.Y(n_276)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_208),
.Y(n_277)
);

NAND2xp33_ASAP7_75t_SL g278 ( 
.A(n_223),
.B(n_178),
.Y(n_278)
);

INVx3_ASAP7_75t_L g279 ( 
.A(n_215),
.Y(n_279)
);

INVx2_ASAP7_75t_L g280 ( 
.A(n_215),
.Y(n_280)
);

INVx2_ASAP7_75t_L g281 ( 
.A(n_215),
.Y(n_281)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_229),
.Y(n_282)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_215),
.Y(n_283)
);

INVx1_ASAP7_75t_SL g284 ( 
.A(n_214),
.Y(n_284)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_217),
.Y(n_285)
);

BUFx10_ASAP7_75t_L g286 ( 
.A(n_223),
.Y(n_286)
);

INVx2_ASAP7_75t_L g287 ( 
.A(n_217),
.Y(n_287)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_217),
.Y(n_288)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_217),
.Y(n_289)
);

INVx2_ASAP7_75t_L g290 ( 
.A(n_218),
.Y(n_290)
);

NAND2xp5_ASAP7_75t_L g291 ( 
.A(n_211),
.B(n_190),
.Y(n_291)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_218),
.Y(n_292)
);

INVx1_ASAP7_75t_SL g293 ( 
.A(n_219),
.Y(n_293)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_218),
.Y(n_294)
);

INVx3_ASAP7_75t_L g295 ( 
.A(n_218),
.Y(n_295)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_231),
.Y(n_296)
);

BUFx6f_ASAP7_75t_L g297 ( 
.A(n_237),
.Y(n_297)
);

BUFx3_ASAP7_75t_L g298 ( 
.A(n_211),
.Y(n_298)
);

NAND2xp5_ASAP7_75t_L g299 ( 
.A(n_298),
.B(n_211),
.Y(n_299)
);

NAND2xp5_ASAP7_75t_L g300 ( 
.A(n_298),
.B(n_239),
.Y(n_300)
);

NAND2xp5_ASAP7_75t_L g301 ( 
.A(n_260),
.B(n_239),
.Y(n_301)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_282),
.Y(n_302)
);

NAND2xp5_ASAP7_75t_L g303 ( 
.A(n_264),
.B(n_250),
.Y(n_303)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_296),
.Y(n_304)
);

INVx3_ASAP7_75t_L g305 ( 
.A(n_297),
.Y(n_305)
);

A2O1A1Ixp33_ASAP7_75t_L g306 ( 
.A1(n_291),
.A2(n_239),
.B(n_234),
.C(n_241),
.Y(n_306)
);

NAND2xp5_ASAP7_75t_L g307 ( 
.A(n_264),
.B(n_230),
.Y(n_307)
);

NOR2xp33_ASAP7_75t_L g308 ( 
.A(n_251),
.B(n_220),
.Y(n_308)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_255),
.Y(n_309)
);

HB1xp67_ASAP7_75t_L g310 ( 
.A(n_284),
.Y(n_310)
);

NAND2xp5_ASAP7_75t_L g311 ( 
.A(n_264),
.B(n_230),
.Y(n_311)
);

NOR2xp33_ASAP7_75t_L g312 ( 
.A(n_254),
.B(n_242),
.Y(n_312)
);

HB1xp67_ASAP7_75t_L g313 ( 
.A(n_293),
.Y(n_313)
);

NAND2xp5_ASAP7_75t_L g314 ( 
.A(n_286),
.B(n_230),
.Y(n_314)
);

NAND2xp5_ASAP7_75t_L g315 ( 
.A(n_286),
.B(n_243),
.Y(n_315)
);

OAI22xp5_ASAP7_75t_L g316 ( 
.A1(n_261),
.A2(n_178),
.B1(n_238),
.B2(n_210),
.Y(n_316)
);

NAND2xp5_ASAP7_75t_SL g317 ( 
.A(n_276),
.B(n_206),
.Y(n_317)
);

NAND2xp5_ASAP7_75t_L g318 ( 
.A(n_272),
.B(n_237),
.Y(n_318)
);

AOI221xp5_ASAP7_75t_L g319 ( 
.A1(n_278),
.A2(n_238),
.B1(n_209),
.B2(n_192),
.C(n_199),
.Y(n_319)
);

AND2x6_ASAP7_75t_L g320 ( 
.A(n_253),
.B(n_191),
.Y(n_320)
);

NAND2xp5_ASAP7_75t_L g321 ( 
.A(n_255),
.B(n_237),
.Y(n_321)
);

INVx2_ASAP7_75t_L g322 ( 
.A(n_253),
.Y(n_322)
);

NAND2xp5_ASAP7_75t_L g323 ( 
.A(n_257),
.B(n_237),
.Y(n_323)
);

INVxp67_ASAP7_75t_L g324 ( 
.A(n_252),
.Y(n_324)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_257),
.Y(n_325)
);

NAND2xp5_ASAP7_75t_SL g326 ( 
.A(n_278),
.B(n_164),
.Y(n_326)
);

INVx1_ASAP7_75t_SL g327 ( 
.A(n_273),
.Y(n_327)
);

NOR2xp67_ASAP7_75t_L g328 ( 
.A(n_256),
.B(n_165),
.Y(n_328)
);

INVx2_ASAP7_75t_L g329 ( 
.A(n_258),
.Y(n_329)
);

INVxp67_ASAP7_75t_L g330 ( 
.A(n_261),
.Y(n_330)
);

NAND3xp33_ASAP7_75t_L g331 ( 
.A(n_261),
.B(n_240),
.C(n_246),
.Y(n_331)
);

AOI22xp33_ASAP7_75t_L g332 ( 
.A1(n_261),
.A2(n_240),
.B1(n_246),
.B2(n_245),
.Y(n_332)
);

BUFx6f_ASAP7_75t_L g333 ( 
.A(n_297),
.Y(n_333)
);

NAND2xp5_ASAP7_75t_SL g334 ( 
.A(n_297),
.B(n_168),
.Y(n_334)
);

NOR2xp33_ASAP7_75t_L g335 ( 
.A(n_269),
.B(n_240),
.Y(n_335)
);

NOR2xp33_ASAP7_75t_L g336 ( 
.A(n_269),
.B(n_274),
.Y(n_336)
);

INVxp67_ASAP7_75t_L g337 ( 
.A(n_266),
.Y(n_337)
);

INVx1_ASAP7_75t_L g338 ( 
.A(n_277),
.Y(n_338)
);

NAND2xp5_ASAP7_75t_L g339 ( 
.A(n_259),
.B(n_240),
.Y(n_339)
);

NAND2xp5_ASAP7_75t_SL g340 ( 
.A(n_297),
.B(n_173),
.Y(n_340)
);

NAND2xp5_ASAP7_75t_L g341 ( 
.A(n_259),
.B(n_244),
.Y(n_341)
);

NAND2xp5_ASAP7_75t_SL g342 ( 
.A(n_297),
.B(n_174),
.Y(n_342)
);

HB1xp67_ASAP7_75t_L g343 ( 
.A(n_263),
.Y(n_343)
);

OAI21xp33_ASAP7_75t_L g344 ( 
.A1(n_263),
.A2(n_201),
.B(n_195),
.Y(n_344)
);

AOI22xp33_ASAP7_75t_L g345 ( 
.A1(n_265),
.A2(n_244),
.B1(n_246),
.B2(n_245),
.Y(n_345)
);

NAND2xp5_ASAP7_75t_L g346 ( 
.A(n_265),
.B(n_244),
.Y(n_346)
);

INVx2_ASAP7_75t_L g347 ( 
.A(n_268),
.Y(n_347)
);

AND2x6_ASAP7_75t_L g348 ( 
.A(n_268),
.B(n_212),
.Y(n_348)
);

NAND2xp5_ASAP7_75t_L g349 ( 
.A(n_270),
.B(n_244),
.Y(n_349)
);

NAND2xp5_ASAP7_75t_L g350 ( 
.A(n_270),
.B(n_245),
.Y(n_350)
);

A2O1A1Ixp33_ASAP7_75t_L g351 ( 
.A1(n_271),
.A2(n_249),
.B(n_212),
.C(n_224),
.Y(n_351)
);

BUFx8_ASAP7_75t_L g352 ( 
.A(n_271),
.Y(n_352)
);

NOR2xp33_ASAP7_75t_L g353 ( 
.A(n_262),
.B(n_245),
.Y(n_353)
);

NAND2xp5_ASAP7_75t_SL g354 ( 
.A(n_275),
.B(n_177),
.Y(n_354)
);

NAND2xp5_ASAP7_75t_SL g355 ( 
.A(n_275),
.B(n_179),
.Y(n_355)
);

NOR2xp33_ASAP7_75t_L g356 ( 
.A(n_262),
.B(n_246),
.Y(n_356)
);

INVx1_ASAP7_75t_L g357 ( 
.A(n_277),
.Y(n_357)
);

NOR2xp67_ASAP7_75t_SL g358 ( 
.A(n_267),
.B(n_224),
.Y(n_358)
);

AND2x4_ASAP7_75t_L g359 ( 
.A(n_280),
.B(n_227),
.Y(n_359)
);

AO22x1_ASAP7_75t_L g360 ( 
.A1(n_283),
.A2(n_193),
.B1(n_189),
.B2(n_186),
.Y(n_360)
);

NOR3xp33_ASAP7_75t_L g361 ( 
.A(n_324),
.B(n_227),
.C(n_232),
.Y(n_361)
);

AOI22xp5_ASAP7_75t_L g362 ( 
.A1(n_330),
.A2(n_232),
.B1(n_233),
.B2(n_249),
.Y(n_362)
);

AOI21xp5_ASAP7_75t_L g363 ( 
.A1(n_299),
.A2(n_300),
.B(n_301),
.Y(n_363)
);

NAND2xp5_ASAP7_75t_L g364 ( 
.A(n_303),
.B(n_280),
.Y(n_364)
);

A2O1A1Ixp33_ASAP7_75t_L g365 ( 
.A1(n_312),
.A2(n_233),
.B(n_287),
.C(n_281),
.Y(n_365)
);

INVx3_ASAP7_75t_L g366 ( 
.A(n_359),
.Y(n_366)
);

NAND3xp33_ASAP7_75t_L g367 ( 
.A(n_308),
.B(n_289),
.C(n_294),
.Y(n_367)
);

OAI21xp5_ASAP7_75t_L g368 ( 
.A1(n_307),
.A2(n_289),
.B(n_294),
.Y(n_368)
);

NAND2xp5_ASAP7_75t_L g369 ( 
.A(n_343),
.B(n_281),
.Y(n_369)
);

INVx2_ASAP7_75t_L g370 ( 
.A(n_359),
.Y(n_370)
);

AOI21xp5_ASAP7_75t_L g371 ( 
.A1(n_311),
.A2(n_318),
.B(n_315),
.Y(n_371)
);

NAND2xp5_ASAP7_75t_L g372 ( 
.A(n_306),
.B(n_287),
.Y(n_372)
);

NOR2x1_ASAP7_75t_L g373 ( 
.A(n_328),
.B(n_267),
.Y(n_373)
);

A2O1A1Ixp33_ASAP7_75t_L g374 ( 
.A1(n_319),
.A2(n_290),
.B(n_292),
.C(n_288),
.Y(n_374)
);

NAND3xp33_ASAP7_75t_SL g375 ( 
.A(n_316),
.B(n_283),
.C(n_285),
.Y(n_375)
);

AND2x2_ASAP7_75t_L g376 ( 
.A(n_310),
.B(n_279),
.Y(n_376)
);

INVx1_ASAP7_75t_L g377 ( 
.A(n_302),
.Y(n_377)
);

NAND2xp5_ASAP7_75t_SL g378 ( 
.A(n_313),
.B(n_295),
.Y(n_378)
);

O2A1O1Ixp33_ASAP7_75t_L g379 ( 
.A1(n_351),
.A2(n_1),
.B(n_2),
.C(n_3),
.Y(n_379)
);

O2A1O1Ixp33_ASAP7_75t_L g380 ( 
.A1(n_326),
.A2(n_2),
.B(n_3),
.C(n_4),
.Y(n_380)
);

AOI21xp5_ASAP7_75t_L g381 ( 
.A1(n_314),
.A2(n_86),
.B(n_149),
.Y(n_381)
);

O2A1O1Ixp33_ASAP7_75t_L g382 ( 
.A1(n_317),
.A2(n_5),
.B(n_6),
.C(n_7),
.Y(n_382)
);

OAI21xp5_ASAP7_75t_L g383 ( 
.A1(n_336),
.A2(n_82),
.B(n_147),
.Y(n_383)
);

NAND2xp5_ASAP7_75t_L g384 ( 
.A(n_309),
.B(n_26),
.Y(n_384)
);

NOR2xp33_ASAP7_75t_L g385 ( 
.A(n_304),
.B(n_5),
.Y(n_385)
);

NAND2xp5_ASAP7_75t_L g386 ( 
.A(n_325),
.B(n_338),
.Y(n_386)
);

AOI21xp5_ASAP7_75t_L g387 ( 
.A1(n_321),
.A2(n_87),
.B(n_145),
.Y(n_387)
);

AOI21xp5_ASAP7_75t_L g388 ( 
.A1(n_323),
.A2(n_80),
.B(n_144),
.Y(n_388)
);

NAND2xp5_ASAP7_75t_L g389 ( 
.A(n_357),
.B(n_27),
.Y(n_389)
);

INVx1_ASAP7_75t_L g390 ( 
.A(n_339),
.Y(n_390)
);

INVx1_ASAP7_75t_L g391 ( 
.A(n_341),
.Y(n_391)
);

INVx2_ASAP7_75t_L g392 ( 
.A(n_322),
.Y(n_392)
);

HB1xp67_ASAP7_75t_L g393 ( 
.A(n_327),
.Y(n_393)
);

AOI21xp5_ASAP7_75t_L g394 ( 
.A1(n_346),
.A2(n_79),
.B(n_142),
.Y(n_394)
);

AOI21xp5_ASAP7_75t_L g395 ( 
.A1(n_349),
.A2(n_350),
.B(n_354),
.Y(n_395)
);

NAND2xp5_ASAP7_75t_L g396 ( 
.A(n_332),
.B(n_29),
.Y(n_396)
);

BUFx3_ASAP7_75t_L g397 ( 
.A(n_352),
.Y(n_397)
);

AOI21x1_ASAP7_75t_L g398 ( 
.A1(n_358),
.A2(n_89),
.B(n_141),
.Y(n_398)
);

AOI21x1_ASAP7_75t_L g399 ( 
.A1(n_329),
.A2(n_77),
.B(n_140),
.Y(n_399)
);

INVx1_ASAP7_75t_L g400 ( 
.A(n_347),
.Y(n_400)
);

INVx3_ASAP7_75t_L g401 ( 
.A(n_348),
.Y(n_401)
);

INVx1_ASAP7_75t_L g402 ( 
.A(n_348),
.Y(n_402)
);

NOR2xp33_ASAP7_75t_L g403 ( 
.A(n_316),
.B(n_6),
.Y(n_403)
);

AOI21xp5_ASAP7_75t_L g404 ( 
.A1(n_355),
.A2(n_76),
.B(n_139),
.Y(n_404)
);

AOI21xp5_ASAP7_75t_L g405 ( 
.A1(n_334),
.A2(n_74),
.B(n_138),
.Y(n_405)
);

INVx2_ASAP7_75t_L g406 ( 
.A(n_333),
.Y(n_406)
);

AOI21xp5_ASAP7_75t_L g407 ( 
.A1(n_340),
.A2(n_73),
.B(n_137),
.Y(n_407)
);

AOI21xp33_ASAP7_75t_L g408 ( 
.A1(n_337),
.A2(n_7),
.B(n_8),
.Y(n_408)
);

NAND2xp5_ASAP7_75t_L g409 ( 
.A(n_305),
.B(n_30),
.Y(n_409)
);

AND2x2_ASAP7_75t_L g410 ( 
.A(n_327),
.B(n_8),
.Y(n_410)
);

INVxp67_ASAP7_75t_L g411 ( 
.A(n_352),
.Y(n_411)
);

NAND2xp5_ASAP7_75t_L g412 ( 
.A(n_305),
.B(n_32),
.Y(n_412)
);

BUFx5_ASAP7_75t_L g413 ( 
.A(n_348),
.Y(n_413)
);

NAND2xp5_ASAP7_75t_L g414 ( 
.A(n_360),
.B(n_34),
.Y(n_414)
);

NOR2xp67_ASAP7_75t_L g415 ( 
.A(n_331),
.B(n_35),
.Y(n_415)
);

AOI22xp5_ASAP7_75t_L g416 ( 
.A1(n_342),
.A2(n_93),
.B1(n_135),
.B2(n_134),
.Y(n_416)
);

INVx2_ASAP7_75t_L g417 ( 
.A(n_333),
.Y(n_417)
);

NOR2x1_ASAP7_75t_L g418 ( 
.A(n_353),
.B(n_36),
.Y(n_418)
);

AOI21xp5_ASAP7_75t_L g419 ( 
.A1(n_335),
.A2(n_356),
.B(n_344),
.Y(n_419)
);

BUFx4f_ASAP7_75t_L g420 ( 
.A(n_320),
.Y(n_420)
);

AOI21xp5_ASAP7_75t_L g421 ( 
.A1(n_333),
.A2(n_92),
.B(n_133),
.Y(n_421)
);

INVx3_ASAP7_75t_L g422 ( 
.A(n_348),
.Y(n_422)
);

NAND2xp5_ASAP7_75t_SL g423 ( 
.A(n_345),
.B(n_9),
.Y(n_423)
);

NAND2xp5_ASAP7_75t_L g424 ( 
.A(n_320),
.B(n_90),
.Y(n_424)
);

NAND2xp5_ASAP7_75t_L g425 ( 
.A(n_320),
.B(n_94),
.Y(n_425)
);

INVx3_ASAP7_75t_L g426 ( 
.A(n_320),
.Y(n_426)
);

OAI21x1_ASAP7_75t_L g427 ( 
.A1(n_395),
.A2(n_150),
.B(n_71),
.Y(n_427)
);

OR2x6_ASAP7_75t_L g428 ( 
.A(n_397),
.B(n_9),
.Y(n_428)
);

OAI21xp5_ASAP7_75t_L g429 ( 
.A1(n_363),
.A2(n_95),
.B(n_131),
.Y(n_429)
);

NOR4xp25_ASAP7_75t_L g430 ( 
.A(n_382),
.B(n_10),
.C(n_11),
.D(n_12),
.Y(n_430)
);

OAI21xp5_ASAP7_75t_L g431 ( 
.A1(n_364),
.A2(n_70),
.B(n_126),
.Y(n_431)
);

AO31x2_ASAP7_75t_L g432 ( 
.A1(n_365),
.A2(n_10),
.A3(n_12),
.B(n_13),
.Y(n_432)
);

BUFx2_ASAP7_75t_L g433 ( 
.A(n_393),
.Y(n_433)
);

OAI21x1_ASAP7_75t_SL g434 ( 
.A1(n_383),
.A2(n_97),
.B(n_125),
.Y(n_434)
);

A2O1A1Ixp33_ASAP7_75t_L g435 ( 
.A1(n_371),
.A2(n_14),
.B(n_15),
.C(n_16),
.Y(n_435)
);

INVx2_ASAP7_75t_L g436 ( 
.A(n_366),
.Y(n_436)
);

OAI21xp33_ASAP7_75t_L g437 ( 
.A1(n_403),
.A2(n_15),
.B(n_16),
.Y(n_437)
);

NAND2xp33_ASAP7_75t_L g438 ( 
.A(n_413),
.B(n_100),
.Y(n_438)
);

NAND2xp5_ASAP7_75t_L g439 ( 
.A(n_390),
.B(n_17),
.Y(n_439)
);

A2O1A1Ixp33_ASAP7_75t_L g440 ( 
.A1(n_368),
.A2(n_17),
.B(n_18),
.C(n_37),
.Y(n_440)
);

NAND2xp5_ASAP7_75t_L g441 ( 
.A(n_391),
.B(n_377),
.Y(n_441)
);

AOI221x1_ASAP7_75t_L g442 ( 
.A1(n_419),
.A2(n_101),
.B1(n_38),
.B2(n_42),
.C(n_46),
.Y(n_442)
);

AOI21xp5_ASAP7_75t_L g443 ( 
.A1(n_372),
.A2(n_103),
.B(n_47),
.Y(n_443)
);

INVx1_ASAP7_75t_L g444 ( 
.A(n_370),
.Y(n_444)
);

NAND2x1_ASAP7_75t_L g445 ( 
.A(n_401),
.B(n_104),
.Y(n_445)
);

OAI21xp5_ASAP7_75t_L g446 ( 
.A1(n_402),
.A2(n_102),
.B(n_49),
.Y(n_446)
);

INVx1_ASAP7_75t_L g447 ( 
.A(n_366),
.Y(n_447)
);

AO31x2_ASAP7_75t_L g448 ( 
.A1(n_374),
.A2(n_18),
.A3(n_50),
.B(n_51),
.Y(n_448)
);

OAI22xp5_ASAP7_75t_L g449 ( 
.A1(n_386),
.A2(n_52),
.B1(n_53),
.B2(n_54),
.Y(n_449)
);

AOI21xp5_ASAP7_75t_L g450 ( 
.A1(n_369),
.A2(n_56),
.B(n_57),
.Y(n_450)
);

AOI21xp5_ASAP7_75t_L g451 ( 
.A1(n_401),
.A2(n_62),
.B(n_63),
.Y(n_451)
);

NAND3xp33_ASAP7_75t_SL g452 ( 
.A(n_380),
.B(n_64),
.C(n_65),
.Y(n_452)
);

OAI21x1_ASAP7_75t_L g453 ( 
.A1(n_422),
.A2(n_132),
.B(n_96),
.Y(n_453)
);

NAND2xp5_ASAP7_75t_SL g454 ( 
.A(n_376),
.B(n_66),
.Y(n_454)
);

BUFx2_ASAP7_75t_L g455 ( 
.A(n_410),
.Y(n_455)
);

AOI21xp5_ASAP7_75t_SL g456 ( 
.A1(n_409),
.A2(n_107),
.B(n_108),
.Y(n_456)
);

NAND2xp5_ASAP7_75t_L g457 ( 
.A(n_361),
.B(n_109),
.Y(n_457)
);

AND2x2_ASAP7_75t_L g458 ( 
.A(n_378),
.B(n_110),
.Y(n_458)
);

NAND2xp5_ASAP7_75t_L g459 ( 
.A(n_362),
.B(n_111),
.Y(n_459)
);

AOI22xp33_ASAP7_75t_L g460 ( 
.A1(n_375),
.A2(n_112),
.B1(n_113),
.B2(n_114),
.Y(n_460)
);

INVx1_ASAP7_75t_L g461 ( 
.A(n_400),
.Y(n_461)
);

NAND2xp5_ASAP7_75t_L g462 ( 
.A(n_362),
.B(n_115),
.Y(n_462)
);

INVx2_ASAP7_75t_L g463 ( 
.A(n_392),
.Y(n_463)
);

BUFx10_ASAP7_75t_L g464 ( 
.A(n_385),
.Y(n_464)
);

OAI21x1_ASAP7_75t_L g465 ( 
.A1(n_412),
.A2(n_119),
.B(n_121),
.Y(n_465)
);

OAI21x1_ASAP7_75t_L g466 ( 
.A1(n_399),
.A2(n_426),
.B(n_398),
.Y(n_466)
);

OAI21x1_ASAP7_75t_L g467 ( 
.A1(n_426),
.A2(n_123),
.B(n_389),
.Y(n_467)
);

CKINVDCx11_ASAP7_75t_R g468 ( 
.A(n_411),
.Y(n_468)
);

INVx2_ASAP7_75t_L g469 ( 
.A(n_406),
.Y(n_469)
);

A2O1A1Ixp33_ASAP7_75t_L g470 ( 
.A1(n_367),
.A2(n_396),
.B(n_408),
.C(n_420),
.Y(n_470)
);

INVxp67_ASAP7_75t_L g471 ( 
.A(n_423),
.Y(n_471)
);

OAI21x1_ASAP7_75t_L g472 ( 
.A1(n_384),
.A2(n_417),
.B(n_373),
.Y(n_472)
);

NAND2xp5_ASAP7_75t_L g473 ( 
.A(n_415),
.B(n_413),
.Y(n_473)
);

NAND2xp5_ASAP7_75t_L g474 ( 
.A(n_413),
.B(n_414),
.Y(n_474)
);

OAI21x1_ASAP7_75t_L g475 ( 
.A1(n_405),
.A2(n_407),
.B(n_404),
.Y(n_475)
);

NAND2xp5_ASAP7_75t_L g476 ( 
.A(n_413),
.B(n_418),
.Y(n_476)
);

OAI21x1_ASAP7_75t_L g477 ( 
.A1(n_387),
.A2(n_388),
.B(n_394),
.Y(n_477)
);

A2O1A1Ixp33_ASAP7_75t_L g478 ( 
.A1(n_420),
.A2(n_379),
.B(n_416),
.C(n_381),
.Y(n_478)
);

INVx4_ASAP7_75t_L g479 ( 
.A(n_413),
.Y(n_479)
);

NAND2xp5_ASAP7_75t_L g480 ( 
.A(n_425),
.B(n_424),
.Y(n_480)
);

INVx4_ASAP7_75t_L g481 ( 
.A(n_421),
.Y(n_481)
);

INVx5_ASAP7_75t_L g482 ( 
.A(n_426),
.Y(n_482)
);

AO21x1_ASAP7_75t_L g483 ( 
.A1(n_429),
.A2(n_431),
.B(n_446),
.Y(n_483)
);

INVx2_ASAP7_75t_L g484 ( 
.A(n_436),
.Y(n_484)
);

AOI21xp33_ASAP7_75t_SL g485 ( 
.A1(n_428),
.A2(n_437),
.B(n_433),
.Y(n_485)
);

CKINVDCx16_ASAP7_75t_R g486 ( 
.A(n_464),
.Y(n_486)
);

AOI22xp33_ASAP7_75t_L g487 ( 
.A1(n_437),
.A2(n_452),
.B1(n_471),
.B2(n_454),
.Y(n_487)
);

INVx1_ASAP7_75t_L g488 ( 
.A(n_447),
.Y(n_488)
);

OAI221xp5_ASAP7_75t_L g489 ( 
.A1(n_455),
.A2(n_441),
.B1(n_460),
.B2(n_440),
.C(n_430),
.Y(n_489)
);

AO21x2_ASAP7_75t_L g490 ( 
.A1(n_434),
.A2(n_429),
.B(n_478),
.Y(n_490)
);

OAI21x1_ASAP7_75t_L g491 ( 
.A1(n_427),
.A2(n_477),
.B(n_475),
.Y(n_491)
);

AOI22xp33_ASAP7_75t_L g492 ( 
.A1(n_444),
.A2(n_458),
.B1(n_439),
.B2(n_463),
.Y(n_492)
);

CKINVDCx16_ASAP7_75t_R g493 ( 
.A(n_464),
.Y(n_493)
);

INVx2_ASAP7_75t_L g494 ( 
.A(n_469),
.Y(n_494)
);

INVx1_ASAP7_75t_L g495 ( 
.A(n_461),
.Y(n_495)
);

AOI22xp33_ASAP7_75t_SL g496 ( 
.A1(n_431),
.A2(n_459),
.B1(n_462),
.B2(n_428),
.Y(n_496)
);

AND2x4_ASAP7_75t_L g497 ( 
.A(n_482),
.B(n_481),
.Y(n_497)
);

INVx2_ASAP7_75t_L g498 ( 
.A(n_482),
.Y(n_498)
);

NAND2xp5_ASAP7_75t_L g499 ( 
.A(n_470),
.B(n_474),
.Y(n_499)
);

INVx3_ASAP7_75t_L g500 ( 
.A(n_479),
.Y(n_500)
);

OAI21xp5_ASAP7_75t_L g501 ( 
.A1(n_480),
.A2(n_476),
.B(n_473),
.Y(n_501)
);

AO21x2_ASAP7_75t_L g502 ( 
.A1(n_435),
.A2(n_443),
.B(n_430),
.Y(n_502)
);

OAI21x1_ASAP7_75t_L g503 ( 
.A1(n_453),
.A2(n_465),
.B(n_445),
.Y(n_503)
);

INVx2_ASAP7_75t_L g504 ( 
.A(n_482),
.Y(n_504)
);

AO21x2_ASAP7_75t_L g505 ( 
.A1(n_457),
.A2(n_438),
.B(n_450),
.Y(n_505)
);

INVx2_ASAP7_75t_L g506 ( 
.A(n_432),
.Y(n_506)
);

OA21x2_ASAP7_75t_L g507 ( 
.A1(n_442),
.A2(n_451),
.B(n_449),
.Y(n_507)
);

CKINVDCx16_ASAP7_75t_R g508 ( 
.A(n_428),
.Y(n_508)
);

BUFx3_ASAP7_75t_L g509 ( 
.A(n_468),
.Y(n_509)
);

INVx2_ASAP7_75t_L g510 ( 
.A(n_432),
.Y(n_510)
);

OAI21x1_ASAP7_75t_L g511 ( 
.A1(n_456),
.A2(n_479),
.B(n_481),
.Y(n_511)
);

INVx5_ASAP7_75t_L g512 ( 
.A(n_448),
.Y(n_512)
);

CKINVDCx5p33_ASAP7_75t_R g513 ( 
.A(n_432),
.Y(n_513)
);

INVx1_ASAP7_75t_L g514 ( 
.A(n_448),
.Y(n_514)
);

INVx3_ASAP7_75t_L g515 ( 
.A(n_448),
.Y(n_515)
);

O2A1O1Ixp33_ASAP7_75t_L g516 ( 
.A1(n_437),
.A2(n_403),
.B(n_439),
.C(n_440),
.Y(n_516)
);

CKINVDCx11_ASAP7_75t_R g517 ( 
.A(n_468),
.Y(n_517)
);

AND2x4_ASAP7_75t_L g518 ( 
.A(n_436),
.B(n_447),
.Y(n_518)
);

OAI21x1_ASAP7_75t_L g519 ( 
.A1(n_466),
.A2(n_472),
.B(n_467),
.Y(n_519)
);

INVx1_ASAP7_75t_L g520 ( 
.A(n_447),
.Y(n_520)
);

AO21x1_ASAP7_75t_L g521 ( 
.A1(n_429),
.A2(n_431),
.B(n_383),
.Y(n_521)
);

INVx1_ASAP7_75t_L g522 ( 
.A(n_447),
.Y(n_522)
);

CKINVDCx5p33_ASAP7_75t_R g523 ( 
.A(n_468),
.Y(n_523)
);

INVx2_ASAP7_75t_L g524 ( 
.A(n_436),
.Y(n_524)
);

O2A1O1Ixp33_ASAP7_75t_L g525 ( 
.A1(n_437),
.A2(n_403),
.B(n_439),
.C(n_440),
.Y(n_525)
);

HB1xp67_ASAP7_75t_L g526 ( 
.A(n_433),
.Y(n_526)
);

AND2x2_ASAP7_75t_L g527 ( 
.A(n_455),
.B(n_441),
.Y(n_527)
);

INVx1_ASAP7_75t_L g528 ( 
.A(n_495),
.Y(n_528)
);

OA21x2_ASAP7_75t_L g529 ( 
.A1(n_514),
.A2(n_510),
.B(n_506),
.Y(n_529)
);

INVx1_ASAP7_75t_L g530 ( 
.A(n_495),
.Y(n_530)
);

INVx2_ASAP7_75t_L g531 ( 
.A(n_494),
.Y(n_531)
);

INVx2_ASAP7_75t_SL g532 ( 
.A(n_526),
.Y(n_532)
);

AND2x4_ASAP7_75t_L g533 ( 
.A(n_497),
.B(n_518),
.Y(n_533)
);

A2O1A1Ixp33_ASAP7_75t_L g534 ( 
.A1(n_516),
.A2(n_525),
.B(n_496),
.C(n_487),
.Y(n_534)
);

INVx2_ASAP7_75t_L g535 ( 
.A(n_506),
.Y(n_535)
);

OR2x2_ASAP7_75t_L g536 ( 
.A(n_499),
.B(n_489),
.Y(n_536)
);

AND2x2_ASAP7_75t_L g537 ( 
.A(n_527),
.B(n_484),
.Y(n_537)
);

INVx1_ASAP7_75t_L g538 ( 
.A(n_494),
.Y(n_538)
);

AND2x2_ASAP7_75t_L g539 ( 
.A(n_527),
.B(n_484),
.Y(n_539)
);

OAI221xp5_ASAP7_75t_L g540 ( 
.A1(n_485),
.A2(n_492),
.B1(n_501),
.B2(n_488),
.C(n_522),
.Y(n_540)
);

INVx2_ASAP7_75t_L g541 ( 
.A(n_524),
.Y(n_541)
);

AO21x2_ASAP7_75t_L g542 ( 
.A1(n_521),
.A2(n_483),
.B(n_491),
.Y(n_542)
);

INVx3_ASAP7_75t_L g543 ( 
.A(n_500),
.Y(n_543)
);

NAND2x1p5_ASAP7_75t_L g544 ( 
.A(n_500),
.B(n_497),
.Y(n_544)
);

BUFx2_ASAP7_75t_L g545 ( 
.A(n_518),
.Y(n_545)
);

INVx1_ASAP7_75t_L g546 ( 
.A(n_488),
.Y(n_546)
);

OR2x2_ASAP7_75t_L g547 ( 
.A(n_486),
.B(n_493),
.Y(n_547)
);

HB1xp67_ASAP7_75t_L g548 ( 
.A(n_524),
.Y(n_548)
);

INVx1_ASAP7_75t_L g549 ( 
.A(n_520),
.Y(n_549)
);

INVx1_ASAP7_75t_L g550 ( 
.A(n_522),
.Y(n_550)
);

OR2x6_ASAP7_75t_L g551 ( 
.A(n_521),
.B(n_483),
.Y(n_551)
);

INVx1_ASAP7_75t_L g552 ( 
.A(n_510),
.Y(n_552)
);

INVx2_ASAP7_75t_SL g553 ( 
.A(n_498),
.Y(n_553)
);

INVx2_ASAP7_75t_L g554 ( 
.A(n_518),
.Y(n_554)
);

INVx2_ASAP7_75t_L g555 ( 
.A(n_498),
.Y(n_555)
);

INVx2_ASAP7_75t_L g556 ( 
.A(n_504),
.Y(n_556)
);

INVx1_ASAP7_75t_L g557 ( 
.A(n_514),
.Y(n_557)
);

INVx2_ASAP7_75t_L g558 ( 
.A(n_504),
.Y(n_558)
);

INVx2_ASAP7_75t_SL g559 ( 
.A(n_497),
.Y(n_559)
);

INVx1_ASAP7_75t_L g560 ( 
.A(n_515),
.Y(n_560)
);

INVx1_ASAP7_75t_L g561 ( 
.A(n_515),
.Y(n_561)
);

AND2x2_ASAP7_75t_L g562 ( 
.A(n_537),
.B(n_513),
.Y(n_562)
);

AND2x2_ASAP7_75t_L g563 ( 
.A(n_537),
.B(n_513),
.Y(n_563)
);

INVx3_ASAP7_75t_L g564 ( 
.A(n_543),
.Y(n_564)
);

OR2x2_ASAP7_75t_L g565 ( 
.A(n_536),
.B(n_502),
.Y(n_565)
);

INVx1_ASAP7_75t_L g566 ( 
.A(n_557),
.Y(n_566)
);

AND2x2_ASAP7_75t_L g567 ( 
.A(n_539),
.B(n_502),
.Y(n_567)
);

HB1xp67_ASAP7_75t_L g568 ( 
.A(n_532),
.Y(n_568)
);

OR2x2_ASAP7_75t_L g569 ( 
.A(n_536),
.B(n_502),
.Y(n_569)
);

INVxp67_ASAP7_75t_SL g570 ( 
.A(n_539),
.Y(n_570)
);

INVx1_ASAP7_75t_L g571 ( 
.A(n_557),
.Y(n_571)
);

INVx1_ASAP7_75t_L g572 ( 
.A(n_552),
.Y(n_572)
);

OR2x2_ASAP7_75t_L g573 ( 
.A(n_551),
.B(n_490),
.Y(n_573)
);

INVx1_ASAP7_75t_L g574 ( 
.A(n_552),
.Y(n_574)
);

HB1xp67_ASAP7_75t_L g575 ( 
.A(n_532),
.Y(n_575)
);

INVx2_ASAP7_75t_SL g576 ( 
.A(n_533),
.Y(n_576)
);

AND2x2_ASAP7_75t_L g577 ( 
.A(n_554),
.B(n_490),
.Y(n_577)
);

AND2x2_ASAP7_75t_L g578 ( 
.A(n_554),
.B(n_490),
.Y(n_578)
);

BUFx3_ASAP7_75t_L g579 ( 
.A(n_533),
.Y(n_579)
);

INVx1_ASAP7_75t_L g580 ( 
.A(n_535),
.Y(n_580)
);

INVx2_ASAP7_75t_L g581 ( 
.A(n_531),
.Y(n_581)
);

NAND2xp5_ASAP7_75t_L g582 ( 
.A(n_545),
.B(n_486),
.Y(n_582)
);

NAND2xp5_ASAP7_75t_L g583 ( 
.A(n_545),
.B(n_493),
.Y(n_583)
);

OR2x2_ASAP7_75t_L g584 ( 
.A(n_551),
.B(n_534),
.Y(n_584)
);

NAND2xp5_ASAP7_75t_L g585 ( 
.A(n_533),
.B(n_508),
.Y(n_585)
);

NOR2xp33_ASAP7_75t_L g586 ( 
.A(n_547),
.B(n_508),
.Y(n_586)
);

INVx1_ASAP7_75t_L g587 ( 
.A(n_529),
.Y(n_587)
);

NOR2xp67_ASAP7_75t_L g588 ( 
.A(n_540),
.B(n_512),
.Y(n_588)
);

AND2x2_ASAP7_75t_L g589 ( 
.A(n_538),
.B(n_541),
.Y(n_589)
);

HB1xp67_ASAP7_75t_L g590 ( 
.A(n_548),
.Y(n_590)
);

OR2x2_ASAP7_75t_L g591 ( 
.A(n_551),
.B(n_507),
.Y(n_591)
);

HB1xp67_ASAP7_75t_L g592 ( 
.A(n_555),
.Y(n_592)
);

AND2x4_ASAP7_75t_L g593 ( 
.A(n_533),
.B(n_511),
.Y(n_593)
);

INVx2_ASAP7_75t_L g594 ( 
.A(n_529),
.Y(n_594)
);

INVx1_ASAP7_75t_L g595 ( 
.A(n_529),
.Y(n_595)
);

BUFx6f_ASAP7_75t_L g596 ( 
.A(n_559),
.Y(n_596)
);

NOR2xp33_ASAP7_75t_L g597 ( 
.A(n_547),
.B(n_523),
.Y(n_597)
);

INVx2_ASAP7_75t_L g598 ( 
.A(n_529),
.Y(n_598)
);

AND2x2_ASAP7_75t_L g599 ( 
.A(n_528),
.B(n_512),
.Y(n_599)
);

INVx1_ASAP7_75t_L g600 ( 
.A(n_560),
.Y(n_600)
);

INVx2_ASAP7_75t_L g601 ( 
.A(n_528),
.Y(n_601)
);

INVx1_ASAP7_75t_L g602 ( 
.A(n_560),
.Y(n_602)
);

BUFx2_ASAP7_75t_L g603 ( 
.A(n_577),
.Y(n_603)
);

INVx1_ASAP7_75t_L g604 ( 
.A(n_587),
.Y(n_604)
);

AND2x2_ASAP7_75t_L g605 ( 
.A(n_567),
.B(n_551),
.Y(n_605)
);

AND2x2_ASAP7_75t_L g606 ( 
.A(n_567),
.B(n_551),
.Y(n_606)
);

INVx2_ASAP7_75t_SL g607 ( 
.A(n_590),
.Y(n_607)
);

HB1xp67_ASAP7_75t_L g608 ( 
.A(n_568),
.Y(n_608)
);

OR2x2_ASAP7_75t_L g609 ( 
.A(n_565),
.B(n_542),
.Y(n_609)
);

NAND2xp5_ASAP7_75t_L g610 ( 
.A(n_570),
.B(n_530),
.Y(n_610)
);

INVx1_ASAP7_75t_L g611 ( 
.A(n_587),
.Y(n_611)
);

INVx1_ASAP7_75t_L g612 ( 
.A(n_595),
.Y(n_612)
);

AND2x2_ASAP7_75t_L g613 ( 
.A(n_562),
.B(n_542),
.Y(n_613)
);

AND2x2_ASAP7_75t_L g614 ( 
.A(n_562),
.B(n_542),
.Y(n_614)
);

INVx2_ASAP7_75t_L g615 ( 
.A(n_594),
.Y(n_615)
);

INVx2_ASAP7_75t_L g616 ( 
.A(n_594),
.Y(n_616)
);

AND2x2_ASAP7_75t_L g617 ( 
.A(n_563),
.B(n_530),
.Y(n_617)
);

INVx2_ASAP7_75t_L g618 ( 
.A(n_601),
.Y(n_618)
);

INVx1_ASAP7_75t_SL g619 ( 
.A(n_575),
.Y(n_619)
);

AND2x2_ASAP7_75t_L g620 ( 
.A(n_563),
.B(n_577),
.Y(n_620)
);

INVx2_ASAP7_75t_L g621 ( 
.A(n_601),
.Y(n_621)
);

INVxp67_ASAP7_75t_SL g622 ( 
.A(n_592),
.Y(n_622)
);

HB1xp67_ASAP7_75t_L g623 ( 
.A(n_589),
.Y(n_623)
);

AND2x2_ASAP7_75t_SL g624 ( 
.A(n_584),
.B(n_507),
.Y(n_624)
);

INVx1_ASAP7_75t_L g625 ( 
.A(n_595),
.Y(n_625)
);

AND2x4_ASAP7_75t_L g626 ( 
.A(n_593),
.B(n_561),
.Y(n_626)
);

AND2x2_ASAP7_75t_L g627 ( 
.A(n_578),
.B(n_556),
.Y(n_627)
);

AND2x2_ASAP7_75t_L g628 ( 
.A(n_578),
.B(n_556),
.Y(n_628)
);

NAND2xp5_ASAP7_75t_L g629 ( 
.A(n_582),
.B(n_583),
.Y(n_629)
);

AND2x2_ASAP7_75t_L g630 ( 
.A(n_584),
.B(n_558),
.Y(n_630)
);

INVx1_ASAP7_75t_L g631 ( 
.A(n_598),
.Y(n_631)
);

INVx2_ASAP7_75t_L g632 ( 
.A(n_566),
.Y(n_632)
);

INVx1_ASAP7_75t_L g633 ( 
.A(n_566),
.Y(n_633)
);

AND2x2_ASAP7_75t_L g634 ( 
.A(n_565),
.B(n_558),
.Y(n_634)
);

AND2x2_ASAP7_75t_L g635 ( 
.A(n_569),
.B(n_571),
.Y(n_635)
);

OR2x2_ASAP7_75t_L g636 ( 
.A(n_569),
.B(n_561),
.Y(n_636)
);

AND2x2_ASAP7_75t_L g637 ( 
.A(n_571),
.B(n_555),
.Y(n_637)
);

AND2x2_ASAP7_75t_L g638 ( 
.A(n_573),
.B(n_550),
.Y(n_638)
);

AOI22xp33_ASAP7_75t_L g639 ( 
.A1(n_588),
.A2(n_505),
.B1(n_559),
.B2(n_509),
.Y(n_639)
);

INVx1_ASAP7_75t_L g640 ( 
.A(n_572),
.Y(n_640)
);

NAND2xp5_ASAP7_75t_L g641 ( 
.A(n_629),
.B(n_572),
.Y(n_641)
);

AND2x2_ASAP7_75t_L g642 ( 
.A(n_620),
.B(n_586),
.Y(n_642)
);

INVx1_ASAP7_75t_L g643 ( 
.A(n_633),
.Y(n_643)
);

INVx1_ASAP7_75t_L g644 ( 
.A(n_633),
.Y(n_644)
);

INVx1_ASAP7_75t_L g645 ( 
.A(n_632),
.Y(n_645)
);

INVx1_ASAP7_75t_L g646 ( 
.A(n_632),
.Y(n_646)
);

AND2x2_ASAP7_75t_L g647 ( 
.A(n_605),
.B(n_573),
.Y(n_647)
);

INVx1_ASAP7_75t_L g648 ( 
.A(n_632),
.Y(n_648)
);

AND2x2_ASAP7_75t_L g649 ( 
.A(n_620),
.B(n_579),
.Y(n_649)
);

OR2x2_ASAP7_75t_L g650 ( 
.A(n_603),
.B(n_591),
.Y(n_650)
);

OR2x2_ASAP7_75t_L g651 ( 
.A(n_603),
.B(n_591),
.Y(n_651)
);

AND2x2_ASAP7_75t_L g652 ( 
.A(n_605),
.B(n_593),
.Y(n_652)
);

OR2x2_ASAP7_75t_L g653 ( 
.A(n_606),
.B(n_593),
.Y(n_653)
);

AND2x2_ASAP7_75t_L g654 ( 
.A(n_606),
.B(n_593),
.Y(n_654)
);

NOR2xp67_ASAP7_75t_L g655 ( 
.A(n_607),
.B(n_597),
.Y(n_655)
);

INVx1_ASAP7_75t_L g656 ( 
.A(n_640),
.Y(n_656)
);

INVx1_ASAP7_75t_L g657 ( 
.A(n_640),
.Y(n_657)
);

INVx1_ASAP7_75t_L g658 ( 
.A(n_604),
.Y(n_658)
);

NAND2xp5_ASAP7_75t_L g659 ( 
.A(n_608),
.B(n_574),
.Y(n_659)
);

AND2x2_ASAP7_75t_L g660 ( 
.A(n_613),
.B(n_599),
.Y(n_660)
);

AND2x2_ASAP7_75t_L g661 ( 
.A(n_613),
.B(n_599),
.Y(n_661)
);

OAI21xp33_ASAP7_75t_L g662 ( 
.A1(n_639),
.A2(n_588),
.B(n_585),
.Y(n_662)
);

NOR2xp33_ASAP7_75t_L g663 ( 
.A(n_619),
.B(n_579),
.Y(n_663)
);

AND2x4_ASAP7_75t_L g664 ( 
.A(n_626),
.B(n_602),
.Y(n_664)
);

NOR2xp33_ASAP7_75t_L g665 ( 
.A(n_607),
.B(n_579),
.Y(n_665)
);

NAND2xp5_ASAP7_75t_L g666 ( 
.A(n_617),
.B(n_623),
.Y(n_666)
);

INVx1_ASAP7_75t_L g667 ( 
.A(n_643),
.Y(n_667)
);

INVx1_ASAP7_75t_L g668 ( 
.A(n_644),
.Y(n_668)
);

INVx2_ASAP7_75t_L g669 ( 
.A(n_664),
.Y(n_669)
);

HB1xp67_ASAP7_75t_L g670 ( 
.A(n_650),
.Y(n_670)
);

OR2x2_ASAP7_75t_L g671 ( 
.A(n_651),
.B(n_609),
.Y(n_671)
);

OAI21xp33_ASAP7_75t_L g672 ( 
.A1(n_662),
.A2(n_630),
.B(n_614),
.Y(n_672)
);

INVx1_ASAP7_75t_L g673 ( 
.A(n_656),
.Y(n_673)
);

INVx1_ASAP7_75t_L g674 ( 
.A(n_657),
.Y(n_674)
);

NAND2xp5_ASAP7_75t_L g675 ( 
.A(n_641),
.B(n_634),
.Y(n_675)
);

OR2x2_ASAP7_75t_L g676 ( 
.A(n_653),
.B(n_609),
.Y(n_676)
);

AND2x4_ASAP7_75t_L g677 ( 
.A(n_652),
.B(n_626),
.Y(n_677)
);

NAND2xp5_ASAP7_75t_L g678 ( 
.A(n_642),
.B(n_634),
.Y(n_678)
);

AND2x4_ASAP7_75t_L g679 ( 
.A(n_652),
.B(n_626),
.Y(n_679)
);

NAND2x2_ASAP7_75t_L g680 ( 
.A(n_659),
.B(n_509),
.Y(n_680)
);

INVx1_ASAP7_75t_L g681 ( 
.A(n_658),
.Y(n_681)
);

NAND2xp5_ASAP7_75t_R g682 ( 
.A(n_663),
.B(n_614),
.Y(n_682)
);

NAND2xp5_ASAP7_75t_L g683 ( 
.A(n_670),
.B(n_647),
.Y(n_683)
);

INVx1_ASAP7_75t_L g684 ( 
.A(n_667),
.Y(n_684)
);

NAND2xp5_ASAP7_75t_L g685 ( 
.A(n_675),
.B(n_647),
.Y(n_685)
);

AND2x2_ASAP7_75t_L g686 ( 
.A(n_677),
.B(n_654),
.Y(n_686)
);

INVx1_ASAP7_75t_L g687 ( 
.A(n_667),
.Y(n_687)
);

AOI22xp5_ASAP7_75t_L g688 ( 
.A1(n_672),
.A2(n_655),
.B1(n_624),
.B2(n_663),
.Y(n_688)
);

OR2x2_ASAP7_75t_L g689 ( 
.A(n_676),
.B(n_660),
.Y(n_689)
);

OR2x2_ASAP7_75t_L g690 ( 
.A(n_671),
.B(n_660),
.Y(n_690)
);

INVx1_ASAP7_75t_L g691 ( 
.A(n_668),
.Y(n_691)
);

NOR2xp33_ASAP7_75t_L g692 ( 
.A(n_678),
.B(n_654),
.Y(n_692)
);

AND2x2_ASAP7_75t_L g693 ( 
.A(n_677),
.B(n_661),
.Y(n_693)
);

AOI21xp33_ASAP7_75t_L g694 ( 
.A1(n_673),
.A2(n_665),
.B(n_664),
.Y(n_694)
);

OR2x2_ASAP7_75t_L g695 ( 
.A(n_690),
.B(n_669),
.Y(n_695)
);

AOI221xp5_ASAP7_75t_L g696 ( 
.A1(n_694),
.A2(n_681),
.B1(n_674),
.B2(n_665),
.C(n_666),
.Y(n_696)
);

INVx1_ASAP7_75t_L g697 ( 
.A(n_684),
.Y(n_697)
);

AOI22xp33_ASAP7_75t_L g698 ( 
.A1(n_688),
.A2(n_680),
.B1(n_624),
.B2(n_664),
.Y(n_698)
);

OR2x2_ASAP7_75t_L g699 ( 
.A(n_689),
.B(n_661),
.Y(n_699)
);

INVx2_ASAP7_75t_L g700 ( 
.A(n_695),
.Y(n_700)
);

NAND2xp5_ASAP7_75t_L g701 ( 
.A(n_696),
.B(n_692),
.Y(n_701)
);

AOI22xp5_ASAP7_75t_L g702 ( 
.A1(n_698),
.A2(n_688),
.B1(n_679),
.B2(n_683),
.Y(n_702)
);

NAND4xp25_ASAP7_75t_L g703 ( 
.A(n_697),
.B(n_691),
.C(n_617),
.D(n_630),
.Y(n_703)
);

OAI321xp33_ASAP7_75t_L g704 ( 
.A1(n_702),
.A2(n_687),
.A3(n_699),
.B1(n_685),
.B2(n_682),
.C(n_610),
.Y(n_704)
);

NAND2xp5_ASAP7_75t_L g705 ( 
.A(n_701),
.B(n_693),
.Y(n_705)
);

AOI21xp5_ASAP7_75t_L g706 ( 
.A1(n_703),
.A2(n_523),
.B(n_679),
.Y(n_706)
);

INVx1_ASAP7_75t_L g707 ( 
.A(n_705),
.Y(n_707)
);

NOR3xp33_ASAP7_75t_L g708 ( 
.A(n_704),
.B(n_517),
.C(n_700),
.Y(n_708)
);

NAND3xp33_ASAP7_75t_SL g709 ( 
.A(n_708),
.B(n_706),
.C(n_686),
.Y(n_709)
);

OAI22xp5_ASAP7_75t_L g710 ( 
.A1(n_707),
.A2(n_624),
.B1(n_649),
.B2(n_648),
.Y(n_710)
);

INVx1_ASAP7_75t_L g711 ( 
.A(n_707),
.Y(n_711)
);

OAI21xp5_ASAP7_75t_L g712 ( 
.A1(n_709),
.A2(n_622),
.B(n_576),
.Y(n_712)
);

AND2x4_ASAP7_75t_L g713 ( 
.A(n_711),
.B(n_635),
.Y(n_713)
);

XNOR2xp5_ASAP7_75t_L g714 ( 
.A(n_710),
.B(n_576),
.Y(n_714)
);

XNOR2xp5_ASAP7_75t_L g715 ( 
.A(n_709),
.B(n_626),
.Y(n_715)
);

XNOR2xp5_ASAP7_75t_L g716 ( 
.A(n_709),
.B(n_638),
.Y(n_716)
);

XOR2x2_ASAP7_75t_L g717 ( 
.A(n_709),
.B(n_507),
.Y(n_717)
);

A2O1A1Ixp33_ASAP7_75t_L g718 ( 
.A1(n_712),
.A2(n_646),
.B(n_645),
.C(n_638),
.Y(n_718)
);

OAI22xp5_ASAP7_75t_L g719 ( 
.A1(n_716),
.A2(n_636),
.B1(n_635),
.B2(n_604),
.Y(n_719)
);

INVx1_ASAP7_75t_L g720 ( 
.A(n_713),
.Y(n_720)
);

NAND2xp33_ASAP7_75t_SL g721 ( 
.A(n_715),
.B(n_596),
.Y(n_721)
);

INVx1_ASAP7_75t_L g722 ( 
.A(n_717),
.Y(n_722)
);

NOR2x1_ASAP7_75t_L g723 ( 
.A(n_714),
.B(n_549),
.Y(n_723)
);

NOR3xp33_ASAP7_75t_L g724 ( 
.A(n_712),
.B(n_553),
.C(n_550),
.Y(n_724)
);

XNOR2xp5_ASAP7_75t_L g725 ( 
.A(n_720),
.B(n_553),
.Y(n_725)
);

AND2x2_ASAP7_75t_L g726 ( 
.A(n_722),
.B(n_723),
.Y(n_726)
);

NAND2xp5_ASAP7_75t_L g727 ( 
.A(n_724),
.B(n_718),
.Y(n_727)
);

NOR3xp33_ASAP7_75t_L g728 ( 
.A(n_721),
.B(n_549),
.C(n_546),
.Y(n_728)
);

INVx1_ASAP7_75t_L g729 ( 
.A(n_719),
.Y(n_729)
);

OAI211xp5_ASAP7_75t_L g730 ( 
.A1(n_722),
.A2(n_546),
.B(n_507),
.C(n_596),
.Y(n_730)
);

AOI22xp5_ASAP7_75t_L g731 ( 
.A1(n_721),
.A2(n_596),
.B1(n_637),
.B2(n_574),
.Y(n_731)
);

AOI22xp5_ASAP7_75t_L g732 ( 
.A1(n_729),
.A2(n_596),
.B1(n_637),
.B2(n_600),
.Y(n_732)
);

NAND3xp33_ASAP7_75t_L g733 ( 
.A(n_726),
.B(n_596),
.C(n_621),
.Y(n_733)
);

OAI22xp5_ASAP7_75t_L g734 ( 
.A1(n_731),
.A2(n_636),
.B1(n_611),
.B2(n_612),
.Y(n_734)
);

CKINVDCx20_ASAP7_75t_R g735 ( 
.A(n_725),
.Y(n_735)
);

AOI22xp5_ASAP7_75t_L g736 ( 
.A1(n_728),
.A2(n_602),
.B1(n_600),
.B2(n_628),
.Y(n_736)
);

INVx3_ASAP7_75t_L g737 ( 
.A(n_727),
.Y(n_737)
);

AO22x2_ASAP7_75t_L g738 ( 
.A1(n_730),
.A2(n_611),
.B1(n_612),
.B2(n_625),
.Y(n_738)
);

NOR2xp33_ASAP7_75t_L g739 ( 
.A(n_729),
.B(n_618),
.Y(n_739)
);

XNOR2xp5_ASAP7_75t_L g740 ( 
.A(n_725),
.B(n_544),
.Y(n_740)
);

INVx2_ASAP7_75t_L g741 ( 
.A(n_735),
.Y(n_741)
);

AOI22xp5_ASAP7_75t_L g742 ( 
.A1(n_737),
.A2(n_628),
.B1(n_627),
.B2(n_625),
.Y(n_742)
);

OAI22x1_ASAP7_75t_L g743 ( 
.A1(n_732),
.A2(n_544),
.B1(n_621),
.B2(n_618),
.Y(n_743)
);

OAI21x1_ASAP7_75t_L g744 ( 
.A1(n_733),
.A2(n_740),
.B(n_739),
.Y(n_744)
);

NAND2xp5_ASAP7_75t_L g745 ( 
.A(n_736),
.B(n_627),
.Y(n_745)
);

OAI22xp33_ASAP7_75t_L g746 ( 
.A1(n_734),
.A2(n_631),
.B1(n_580),
.B2(n_564),
.Y(n_746)
);

INVxp67_ASAP7_75t_SL g747 ( 
.A(n_738),
.Y(n_747)
);

OAI22xp5_ASAP7_75t_L g748 ( 
.A1(n_735),
.A2(n_631),
.B1(n_616),
.B2(n_615),
.Y(n_748)
);

AOI21xp5_ASAP7_75t_L g749 ( 
.A1(n_747),
.A2(n_505),
.B(n_503),
.Y(n_749)
);

AOI21xp5_ASAP7_75t_L g750 ( 
.A1(n_741),
.A2(n_505),
.B(n_503),
.Y(n_750)
);

AOI22xp33_ASAP7_75t_SL g751 ( 
.A1(n_744),
.A2(n_748),
.B1(n_745),
.B2(n_743),
.Y(n_751)
);

AOI21xp33_ASAP7_75t_SL g752 ( 
.A1(n_746),
.A2(n_544),
.B(n_511),
.Y(n_752)
);

XNOR2x1_ASAP7_75t_L g753 ( 
.A(n_742),
.B(n_543),
.Y(n_753)
);

NAND2xp5_ASAP7_75t_L g754 ( 
.A(n_751),
.B(n_753),
.Y(n_754)
);

AO21x2_ASAP7_75t_L g755 ( 
.A1(n_749),
.A2(n_752),
.B(n_750),
.Y(n_755)
);

NOR2xp33_ASAP7_75t_L g756 ( 
.A(n_754),
.B(n_581),
.Y(n_756)
);

AOI21xp5_ASAP7_75t_L g757 ( 
.A1(n_756),
.A2(n_755),
.B(n_519),
.Y(n_757)
);


endmodule