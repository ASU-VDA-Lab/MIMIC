module fake_jpeg_17375_n_249 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_249);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_249;

wire n_159;
wire n_117;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_84;
wire n_59;
wire n_98;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_16;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_223;
wire n_234;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_24;
wire n_44;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_216;
wire n_217;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

INVx1_ASAP7_75t_L g16 ( 
.A(n_15),
.Y(n_16)
);

INVx13_ASAP7_75t_L g17 ( 
.A(n_6),
.Y(n_17)
);

INVx2_ASAP7_75t_L g18 ( 
.A(n_12),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_2),
.Y(n_19)
);

INVx2_ASAP7_75t_L g20 ( 
.A(n_5),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_6),
.Y(n_21)
);

NOR2xp33_ASAP7_75t_L g22 ( 
.A(n_11),
.B(n_9),
.Y(n_22)
);

BUFx12f_ASAP7_75t_L g23 ( 
.A(n_10),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_5),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_12),
.Y(n_25)
);

INVx11_ASAP7_75t_SL g26 ( 
.A(n_7),
.Y(n_26)
);

BUFx3_ASAP7_75t_L g27 ( 
.A(n_13),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_6),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_10),
.Y(n_29)
);

NOR2xp33_ASAP7_75t_L g30 ( 
.A(n_4),
.B(n_15),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_7),
.Y(n_31)
);

NOR2xp33_ASAP7_75t_L g32 ( 
.A(n_11),
.B(n_13),
.Y(n_32)
);

NOR2xp33_ASAP7_75t_L g33 ( 
.A(n_22),
.B(n_15),
.Y(n_33)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_33),
.Y(n_51)
);

INVx11_ASAP7_75t_L g34 ( 
.A(n_17),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_34),
.Y(n_55)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_21),
.Y(n_35)
);

NAND2xp5_ASAP7_75t_SL g61 ( 
.A(n_35),
.B(n_43),
.Y(n_61)
);

INVx8_ASAP7_75t_L g36 ( 
.A(n_17),
.Y(n_36)
);

INVx4_ASAP7_75t_L g44 ( 
.A(n_36),
.Y(n_44)
);

INVx11_ASAP7_75t_L g37 ( 
.A(n_17),
.Y(n_37)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_37),
.Y(n_64)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_23),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_38),
.Y(n_45)
);

BUFx12f_ASAP7_75t_L g39 ( 
.A(n_23),
.Y(n_39)
);

BUFx3_ASAP7_75t_L g50 ( 
.A(n_39),
.Y(n_50)
);

INVx2_ASAP7_75t_L g40 ( 
.A(n_23),
.Y(n_40)
);

INVx2_ASAP7_75t_L g49 ( 
.A(n_40),
.Y(n_49)
);

BUFx8_ASAP7_75t_L g41 ( 
.A(n_26),
.Y(n_41)
);

INVx4_ASAP7_75t_L g53 ( 
.A(n_41),
.Y(n_53)
);

INVx5_ASAP7_75t_L g42 ( 
.A(n_23),
.Y(n_42)
);

INVx3_ASAP7_75t_L g48 ( 
.A(n_42),
.Y(n_48)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_21),
.Y(n_43)
);

OAI22xp33_ASAP7_75t_SL g46 ( 
.A1(n_35),
.A2(n_17),
.B1(n_26),
.B2(n_28),
.Y(n_46)
);

OAI22xp33_ASAP7_75t_SL g86 ( 
.A1(n_46),
.A2(n_25),
.B1(n_37),
.B2(n_36),
.Y(n_86)
);

AOI22xp33_ASAP7_75t_SL g47 ( 
.A1(n_42),
.A2(n_20),
.B1(n_18),
.B2(n_21),
.Y(n_47)
);

AOI22xp33_ASAP7_75t_SL g66 ( 
.A1(n_47),
.A2(n_52),
.B1(n_34),
.B2(n_37),
.Y(n_66)
);

AOI22xp33_ASAP7_75t_SL g52 ( 
.A1(n_42),
.A2(n_20),
.B1(n_18),
.B2(n_19),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_L g54 ( 
.A(n_43),
.B(n_20),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_L g73 ( 
.A(n_54),
.B(n_43),
.Y(n_73)
);

AND2x2_ASAP7_75t_L g56 ( 
.A(n_38),
.B(n_19),
.Y(n_56)
);

OAI21xp33_ASAP7_75t_L g85 ( 
.A1(n_56),
.A2(n_62),
.B(n_31),
.Y(n_85)
);

INVx4_ASAP7_75t_L g57 ( 
.A(n_36),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_57),
.B(n_60),
.Y(n_70)
);

INVx3_ASAP7_75t_L g58 ( 
.A(n_40),
.Y(n_58)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_58),
.Y(n_82)
);

AOI22xp5_ASAP7_75t_L g59 ( 
.A1(n_42),
.A2(n_18),
.B1(n_19),
.B2(n_31),
.Y(n_59)
);

OAI22xp5_ASAP7_75t_SL g81 ( 
.A1(n_59),
.A2(n_63),
.B1(n_29),
.B2(n_24),
.Y(n_81)
);

INVx3_ASAP7_75t_L g60 ( 
.A(n_40),
.Y(n_60)
);

AND2x2_ASAP7_75t_L g62 ( 
.A(n_38),
.B(n_0),
.Y(n_62)
);

OAI22xp5_ASAP7_75t_L g63 ( 
.A1(n_34),
.A2(n_24),
.B1(n_29),
.B2(n_28),
.Y(n_63)
);

INVx2_ASAP7_75t_L g65 ( 
.A(n_39),
.Y(n_65)
);

INVx2_ASAP7_75t_L g69 ( 
.A(n_65),
.Y(n_69)
);

AOI22xp33_ASAP7_75t_SL g97 ( 
.A1(n_66),
.A2(n_53),
.B1(n_44),
.B2(n_57),
.Y(n_97)
);

INVx13_ASAP7_75t_L g67 ( 
.A(n_53),
.Y(n_67)
);

INVx11_ASAP7_75t_L g88 ( 
.A(n_67),
.Y(n_88)
);

OAI22xp5_ASAP7_75t_L g68 ( 
.A1(n_54),
.A2(n_34),
.B1(n_37),
.B2(n_36),
.Y(n_68)
);

AOI22xp5_ASAP7_75t_L g105 ( 
.A1(n_68),
.A2(n_75),
.B1(n_56),
.B2(n_80),
.Y(n_105)
);

INVx2_ASAP7_75t_L g71 ( 
.A(n_49),
.Y(n_71)
);

BUFx2_ASAP7_75t_L g91 ( 
.A(n_71),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_51),
.B(n_33),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_72),
.B(n_76),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_L g108 ( 
.A(n_73),
.B(n_74),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_L g74 ( 
.A(n_56),
.B(n_61),
.Y(n_74)
);

AOI32xp33_ASAP7_75t_L g75 ( 
.A1(n_45),
.A2(n_32),
.A3(n_22),
.B1(n_30),
.B2(n_39),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_SL g76 ( 
.A(n_51),
.B(n_35),
.Y(n_76)
);

INVx4_ASAP7_75t_L g77 ( 
.A(n_55),
.Y(n_77)
);

INVx4_ASAP7_75t_SL g95 ( 
.A(n_77),
.Y(n_95)
);

BUFx12f_ASAP7_75t_L g78 ( 
.A(n_55),
.Y(n_78)
);

INVx5_ASAP7_75t_L g109 ( 
.A(n_78),
.Y(n_109)
);

INVx2_ASAP7_75t_L g79 ( 
.A(n_49),
.Y(n_79)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_79),
.Y(n_93)
);

AND2x4_ASAP7_75t_SL g80 ( 
.A(n_62),
.B(n_39),
.Y(n_80)
);

NAND2xp33_ASAP7_75t_SL g111 ( 
.A(n_80),
.B(n_39),
.Y(n_111)
);

OAI22xp33_ASAP7_75t_SL g101 ( 
.A1(n_81),
.A2(n_85),
.B1(n_86),
.B2(n_62),
.Y(n_101)
);

INVxp67_ASAP7_75t_L g83 ( 
.A(n_65),
.Y(n_83)
);

INVxp67_ASAP7_75t_L g89 ( 
.A(n_83),
.Y(n_89)
);

BUFx12f_ASAP7_75t_L g84 ( 
.A(n_55),
.Y(n_84)
);

INVx8_ASAP7_75t_L g100 ( 
.A(n_84),
.Y(n_100)
);

AOI22xp33_ASAP7_75t_L g87 ( 
.A1(n_63),
.A2(n_25),
.B1(n_16),
.B2(n_30),
.Y(n_87)
);

OAI22xp5_ASAP7_75t_SL g96 ( 
.A1(n_87),
.A2(n_16),
.B1(n_32),
.B2(n_59),
.Y(n_96)
);

MAJIxp5_ASAP7_75t_L g90 ( 
.A(n_74),
.B(n_45),
.C(n_39),
.Y(n_90)
);

MAJIxp5_ASAP7_75t_L g132 ( 
.A(n_90),
.B(n_41),
.C(n_1),
.Y(n_132)
);

CKINVDCx20_ASAP7_75t_R g92 ( 
.A(n_82),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_SL g126 ( 
.A(n_92),
.B(n_96),
.Y(n_126)
);

OAI22xp5_ASAP7_75t_L g127 ( 
.A1(n_97),
.A2(n_105),
.B1(n_110),
.B2(n_27),
.Y(n_127)
);

CKINVDCx20_ASAP7_75t_R g98 ( 
.A(n_82),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g123 ( 
.A(n_98),
.B(n_99),
.Y(n_123)
);

INVx4_ASAP7_75t_L g99 ( 
.A(n_78),
.Y(n_99)
);

NOR2x1_ASAP7_75t_L g134 ( 
.A(n_101),
.B(n_41),
.Y(n_134)
);

INVx2_ASAP7_75t_L g102 ( 
.A(n_69),
.Y(n_102)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_102),
.Y(n_124)
);

INVxp67_ASAP7_75t_L g103 ( 
.A(n_70),
.Y(n_103)
);

INVx1_ASAP7_75t_SL g112 ( 
.A(n_103),
.Y(n_112)
);

BUFx6f_ASAP7_75t_L g104 ( 
.A(n_78),
.Y(n_104)
);

BUFx6f_ASAP7_75t_L g133 ( 
.A(n_104),
.Y(n_133)
);

OAI22xp5_ASAP7_75t_L g106 ( 
.A1(n_73),
.A2(n_60),
.B1(n_58),
.B2(n_48),
.Y(n_106)
);

AOI22xp5_ASAP7_75t_L g128 ( 
.A1(n_106),
.A2(n_41),
.B1(n_84),
.B2(n_2),
.Y(n_128)
);

CKINVDCx20_ASAP7_75t_R g107 ( 
.A(n_78),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_SL g116 ( 
.A(n_107),
.B(n_64),
.Y(n_116)
);

AOI22xp33_ASAP7_75t_SL g110 ( 
.A1(n_80),
.A2(n_48),
.B1(n_44),
.B2(n_64),
.Y(n_110)
);

AND2x2_ASAP7_75t_L g120 ( 
.A(n_111),
.B(n_67),
.Y(n_120)
);

OAI21xp5_ASAP7_75t_L g113 ( 
.A1(n_90),
.A2(n_80),
.B(n_75),
.Y(n_113)
);

OAI21xp5_ASAP7_75t_L g138 ( 
.A1(n_113),
.A2(n_93),
.B(n_91),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_L g114 ( 
.A(n_108),
.B(n_81),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g149 ( 
.A(n_114),
.B(n_115),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_L g115 ( 
.A(n_108),
.B(n_68),
.Y(n_115)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_116),
.Y(n_135)
);

A2O1A1O1Ixp25_ASAP7_75t_L g117 ( 
.A1(n_111),
.A2(n_83),
.B(n_71),
.C(n_79),
.D(n_50),
.Y(n_117)
);

A2O1A1O1Ixp25_ASAP7_75t_L g145 ( 
.A1(n_117),
.A2(n_95),
.B(n_91),
.C(n_88),
.D(n_100),
.Y(n_145)
);

OAI22xp5_ASAP7_75t_L g118 ( 
.A1(n_105),
.A2(n_77),
.B1(n_69),
.B2(n_50),
.Y(n_118)
);

AOI22xp5_ASAP7_75t_L g148 ( 
.A1(n_118),
.A2(n_119),
.B1(n_127),
.B2(n_99),
.Y(n_148)
);

OAI22xp5_ASAP7_75t_L g119 ( 
.A1(n_106),
.A2(n_84),
.B1(n_23),
.B2(n_27),
.Y(n_119)
);

OAI21xp5_ASAP7_75t_SL g152 ( 
.A1(n_120),
.A2(n_134),
.B(n_0),
.Y(n_152)
);

OAI22xp5_ASAP7_75t_SL g121 ( 
.A1(n_96),
.A2(n_23),
.B1(n_27),
.B2(n_84),
.Y(n_121)
);

OAI22xp5_ASAP7_75t_SL g142 ( 
.A1(n_121),
.A2(n_128),
.B1(n_129),
.B2(n_130),
.Y(n_142)
);

NAND3xp33_ASAP7_75t_L g122 ( 
.A(n_94),
.B(n_9),
.C(n_14),
.Y(n_122)
);

INVxp67_ASAP7_75t_L g139 ( 
.A(n_122),
.Y(n_139)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_102),
.Y(n_125)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_125),
.Y(n_140)
);

OAI22xp5_ASAP7_75t_SL g129 ( 
.A1(n_94),
.A2(n_41),
.B1(n_1),
.B2(n_2),
.Y(n_129)
);

OAI22xp5_ASAP7_75t_SL g130 ( 
.A1(n_92),
.A2(n_41),
.B1(n_1),
.B2(n_2),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_SL g131 ( 
.A(n_98),
.B(n_9),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_L g144 ( 
.A(n_131),
.B(n_12),
.Y(n_144)
);

MAJIxp5_ASAP7_75t_L g141 ( 
.A(n_132),
.B(n_93),
.C(n_104),
.Y(n_141)
);

AOI21xp5_ASAP7_75t_L g136 ( 
.A1(n_120),
.A2(n_89),
.B(n_107),
.Y(n_136)
);

OAI21xp5_ASAP7_75t_SL g175 ( 
.A1(n_136),
.A2(n_145),
.B(n_148),
.Y(n_175)
);

XNOR2xp5_ASAP7_75t_SL g137 ( 
.A(n_113),
.B(n_114),
.Y(n_137)
);

XNOR2xp5_ASAP7_75t_SL g172 ( 
.A(n_137),
.B(n_138),
.Y(n_172)
);

XNOR2xp5_ASAP7_75t_L g160 ( 
.A(n_141),
.B(n_152),
.Y(n_160)
);

OAI22xp5_ASAP7_75t_SL g143 ( 
.A1(n_115),
.A2(n_95),
.B1(n_100),
.B2(n_109),
.Y(n_143)
);

OAI22xp5_ASAP7_75t_SL g169 ( 
.A1(n_143),
.A2(n_146),
.B1(n_133),
.B2(n_4),
.Y(n_169)
);

NOR2xp33_ASAP7_75t_SL g166 ( 
.A(n_144),
.B(n_130),
.Y(n_166)
);

OAI22xp5_ASAP7_75t_SL g146 ( 
.A1(n_134),
.A2(n_95),
.B1(n_100),
.B2(n_109),
.Y(n_146)
);

XOR2xp5_ASAP7_75t_L g147 ( 
.A(n_120),
.B(n_91),
.Y(n_147)
);

MAJIxp5_ASAP7_75t_L g163 ( 
.A(n_147),
.B(n_117),
.C(n_112),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_L g150 ( 
.A(n_126),
.B(n_88),
.Y(n_150)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_150),
.Y(n_170)
);

NOR2xp33_ASAP7_75t_L g151 ( 
.A(n_116),
.B(n_104),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_L g178 ( 
.A(n_151),
.B(n_157),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_L g153 ( 
.A(n_132),
.B(n_0),
.Y(n_153)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_153),
.Y(n_177)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_123),
.Y(n_154)
);

CKINVDCx20_ASAP7_75t_R g161 ( 
.A(n_154),
.Y(n_161)
);

CKINVDCx16_ASAP7_75t_R g155 ( 
.A(n_124),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_L g162 ( 
.A(n_155),
.B(n_125),
.Y(n_162)
);

AOI21xp5_ASAP7_75t_L g156 ( 
.A1(n_118),
.A2(n_0),
.B(n_1),
.Y(n_156)
);

AOI21xp5_ASAP7_75t_L g158 ( 
.A1(n_156),
.A2(n_131),
.B(n_152),
.Y(n_158)
);

NOR2xp33_ASAP7_75t_L g157 ( 
.A(n_112),
.B(n_3),
.Y(n_157)
);

OAI22xp5_ASAP7_75t_SL g195 ( 
.A1(n_158),
.A2(n_167),
.B1(n_168),
.B2(n_171),
.Y(n_195)
);

INVxp67_ASAP7_75t_L g159 ( 
.A(n_143),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_L g185 ( 
.A(n_159),
.B(n_176),
.Y(n_185)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_162),
.Y(n_179)
);

MAJIxp5_ASAP7_75t_L g180 ( 
.A(n_163),
.B(n_138),
.C(n_141),
.Y(n_180)
);

XNOR2x1_ASAP7_75t_L g164 ( 
.A(n_137),
.B(n_129),
.Y(n_164)
);

XOR2xp5_ASAP7_75t_L g182 ( 
.A(n_164),
.B(n_142),
.Y(n_182)
);

NOR2xp33_ASAP7_75t_L g165 ( 
.A(n_150),
.B(n_154),
.Y(n_165)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_165),
.Y(n_189)
);

NOR2xp33_ASAP7_75t_SL g194 ( 
.A(n_166),
.B(n_142),
.Y(n_194)
);

AOI22xp5_ASAP7_75t_SL g167 ( 
.A1(n_145),
.A2(n_121),
.B1(n_128),
.B2(n_119),
.Y(n_167)
);

AOI22xp5_ASAP7_75t_L g168 ( 
.A1(n_149),
.A2(n_124),
.B1(n_133),
.B2(n_5),
.Y(n_168)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_169),
.Y(n_192)
);

OAI22xp5_ASAP7_75t_SL g171 ( 
.A1(n_148),
.A2(n_133),
.B1(n_4),
.B2(n_7),
.Y(n_171)
);

AND2x2_ASAP7_75t_SL g173 ( 
.A(n_147),
.B(n_3),
.Y(n_173)
);

AOI22xp5_ASAP7_75t_L g183 ( 
.A1(n_173),
.A2(n_174),
.B1(n_144),
.B2(n_157),
.Y(n_183)
);

AND2x2_ASAP7_75t_L g174 ( 
.A(n_136),
.B(n_3),
.Y(n_174)
);

CKINVDCx20_ASAP7_75t_R g176 ( 
.A(n_140),
.Y(n_176)
);

XNOR2xp5_ASAP7_75t_L g202 ( 
.A(n_180),
.B(n_183),
.Y(n_202)
);

MAJIxp5_ASAP7_75t_L g181 ( 
.A(n_160),
.B(n_149),
.C(n_153),
.Y(n_181)
);

MAJIxp5_ASAP7_75t_L g205 ( 
.A(n_181),
.B(n_184),
.C(n_188),
.Y(n_205)
);

XOR2xp5_ASAP7_75t_L g200 ( 
.A(n_182),
.B(n_191),
.Y(n_200)
);

MAJIxp5_ASAP7_75t_L g184 ( 
.A(n_160),
.B(n_146),
.C(n_140),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_L g186 ( 
.A(n_170),
.B(n_135),
.Y(n_186)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_186),
.Y(n_196)
);

NAND2xp5_ASAP7_75t_L g187 ( 
.A(n_170),
.B(n_135),
.Y(n_187)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_187),
.Y(n_197)
);

MAJIxp5_ASAP7_75t_L g188 ( 
.A(n_172),
.B(n_151),
.C(n_155),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_L g190 ( 
.A(n_161),
.B(n_139),
.Y(n_190)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_190),
.Y(n_199)
);

XNOR2xp5_ASAP7_75t_L g191 ( 
.A(n_172),
.B(n_156),
.Y(n_191)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_168),
.Y(n_193)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_193),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_SL g201 ( 
.A(n_194),
.B(n_159),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_L g198 ( 
.A(n_179),
.B(n_161),
.Y(n_198)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_198),
.Y(n_214)
);

NAND2xp5_ASAP7_75t_L g219 ( 
.A(n_201),
.B(n_206),
.Y(n_219)
);

OAI21xp5_ASAP7_75t_L g204 ( 
.A1(n_185),
.A2(n_158),
.B(n_164),
.Y(n_204)
);

AOI21xp5_ASAP7_75t_L g218 ( 
.A1(n_204),
.A2(n_174),
.B(n_173),
.Y(n_218)
);

AOI22xp5_ASAP7_75t_L g206 ( 
.A1(n_192),
.A2(n_184),
.B1(n_189),
.B2(n_177),
.Y(n_206)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_186),
.Y(n_207)
);

CKINVDCx20_ASAP7_75t_R g212 ( 
.A(n_207),
.Y(n_212)
);

XNOR2xp5_ASAP7_75t_L g208 ( 
.A(n_188),
.B(n_163),
.Y(n_208)
);

MAJIxp5_ASAP7_75t_L g210 ( 
.A(n_208),
.B(n_209),
.C(n_191),
.Y(n_210)
);

XNOR2xp5_ASAP7_75t_L g209 ( 
.A(n_180),
.B(n_175),
.Y(n_209)
);

XOR2xp5_ASAP7_75t_L g221 ( 
.A(n_210),
.B(n_218),
.Y(n_221)
);

AOI22xp5_ASAP7_75t_L g211 ( 
.A1(n_196),
.A2(n_195),
.B1(n_187),
.B2(n_182),
.Y(n_211)
);

NAND2xp5_ASAP7_75t_SL g228 ( 
.A(n_211),
.B(n_216),
.Y(n_228)
);

MAJIxp5_ASAP7_75t_L g213 ( 
.A(n_205),
.B(n_181),
.C(n_177),
.Y(n_213)
);

MAJIxp5_ASAP7_75t_L g222 ( 
.A(n_213),
.B(n_215),
.C(n_217),
.Y(n_222)
);

XNOR2xp5_ASAP7_75t_L g215 ( 
.A(n_202),
.B(n_175),
.Y(n_215)
);

CKINVDCx20_ASAP7_75t_R g216 ( 
.A(n_197),
.Y(n_216)
);

MAJIxp5_ASAP7_75t_L g217 ( 
.A(n_205),
.B(n_173),
.C(n_195),
.Y(n_217)
);

AOI21xp5_ASAP7_75t_L g220 ( 
.A1(n_204),
.A2(n_176),
.B(n_174),
.Y(n_220)
);

XNOR2xp5_ASAP7_75t_L g223 ( 
.A(n_220),
.B(n_169),
.Y(n_223)
);

XOR2xp5_ASAP7_75t_L g230 ( 
.A(n_223),
.B(n_218),
.Y(n_230)
);

AOI21xp5_ASAP7_75t_L g224 ( 
.A1(n_214),
.A2(n_209),
.B(n_199),
.Y(n_224)
);

OAI21xp5_ASAP7_75t_L g234 ( 
.A1(n_224),
.A2(n_210),
.B(n_213),
.Y(n_234)
);

NAND2xp5_ASAP7_75t_L g225 ( 
.A(n_212),
.B(n_178),
.Y(n_225)
);

NAND2xp5_ASAP7_75t_SL g231 ( 
.A(n_225),
.B(n_227),
.Y(n_231)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_211),
.Y(n_226)
);

NAND2xp5_ASAP7_75t_L g233 ( 
.A(n_226),
.B(n_215),
.Y(n_233)
);

NOR2xp33_ASAP7_75t_SL g227 ( 
.A(n_219),
.B(n_183),
.Y(n_227)
);

OAI22xp5_ASAP7_75t_SL g229 ( 
.A1(n_228),
.A2(n_203),
.B1(n_220),
.B2(n_217),
.Y(n_229)
);

NOR2xp33_ASAP7_75t_L g239 ( 
.A(n_229),
.B(n_233),
.Y(n_239)
);

XOR2xp5_ASAP7_75t_L g240 ( 
.A(n_230),
.B(n_200),
.Y(n_240)
);

NOR2xp33_ASAP7_75t_L g232 ( 
.A(n_223),
.B(n_178),
.Y(n_232)
);

NOR2xp33_ASAP7_75t_SL g238 ( 
.A(n_232),
.B(n_235),
.Y(n_238)
);

AOI21xp33_ASAP7_75t_L g237 ( 
.A1(n_234),
.A2(n_221),
.B(n_230),
.Y(n_237)
);

NAND2xp5_ASAP7_75t_L g235 ( 
.A(n_222),
.B(n_202),
.Y(n_235)
);

OAI21xp5_ASAP7_75t_L g236 ( 
.A1(n_234),
.A2(n_222),
.B(n_221),
.Y(n_236)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_236),
.Y(n_243)
);

AOI21xp5_ASAP7_75t_L g244 ( 
.A1(n_237),
.A2(n_240),
.B(n_8),
.Y(n_244)
);

A2O1A1Ixp33_ASAP7_75t_L g241 ( 
.A1(n_239),
.A2(n_231),
.B(n_229),
.C(n_208),
.Y(n_241)
);

HB1xp67_ASAP7_75t_L g245 ( 
.A(n_241),
.Y(n_245)
);

AOI322xp5_ASAP7_75t_L g242 ( 
.A1(n_238),
.A2(n_171),
.A3(n_200),
.B1(n_167),
.B2(n_13),
.C1(n_8),
.C2(n_11),
.Y(n_242)
);

INVxp67_ASAP7_75t_L g246 ( 
.A(n_242),
.Y(n_246)
);

AOI321xp33_ASAP7_75t_L g247 ( 
.A1(n_245),
.A2(n_243),
.A3(n_244),
.B1(n_240),
.B2(n_14),
.C(n_8),
.Y(n_247)
);

NAND3xp33_ASAP7_75t_L g248 ( 
.A(n_247),
.B(n_10),
.C(n_14),
.Y(n_248)
);

XNOR2xp5_ASAP7_75t_L g249 ( 
.A(n_248),
.B(n_246),
.Y(n_249)
);


endmodule