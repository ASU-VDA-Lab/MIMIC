module fake_netlist_6_394_n_981 (n_52, n_16, n_1, n_91, n_119, n_46, n_146, n_163, n_18, n_21, n_147, n_154, n_88, n_3, n_98, n_113, n_39, n_63, n_73, n_4, n_148, n_138, n_22, n_161, n_68, n_166, n_28, n_184, n_50, n_158, n_49, n_7, n_83, n_5, n_101, n_167, n_144, n_174, n_127, n_125, n_153, n_168, n_178, n_77, n_156, n_149, n_152, n_106, n_92, n_145, n_42, n_133, n_96, n_8, n_90, n_160, n_24, n_105, n_131, n_54, n_132, n_188, n_102, n_186, n_0, n_87, n_189, n_32, n_66, n_85, n_99, n_78, n_84, n_130, n_164, n_100, n_129, n_13, n_121, n_11, n_137, n_17, n_23, n_142, n_20, n_143, n_2, n_180, n_19, n_47, n_62, n_29, n_155, n_75, n_109, n_150, n_122, n_45, n_34, n_140, n_70, n_120, n_37, n_15, n_67, n_33, n_82, n_27, n_38, n_110, n_151, n_61, n_112, n_172, n_81, n_59, n_181, n_76, n_36, n_182, n_26, n_124, n_55, n_126, n_94, n_97, n_108, n_58, n_116, n_64, n_117, n_118, n_175, n_48, n_65, n_25, n_40, n_93, n_80, n_141, n_135, n_165, n_139, n_41, n_134, n_177, n_176, n_114, n_86, n_104, n_95, n_179, n_9, n_107, n_10, n_71, n_74, n_6, n_14, n_123, n_136, n_72, n_187, n_89, n_173, n_103, n_111, n_60, n_159, n_157, n_162, n_170, n_185, n_35, n_183, n_115, n_12, n_69, n_128, n_30, n_79, n_43, n_171, n_31, n_57, n_169, n_53, n_51, n_44, n_56, n_981);

input n_52;
input n_16;
input n_1;
input n_91;
input n_119;
input n_46;
input n_146;
input n_163;
input n_18;
input n_21;
input n_147;
input n_154;
input n_88;
input n_3;
input n_98;
input n_113;
input n_39;
input n_63;
input n_73;
input n_4;
input n_148;
input n_138;
input n_22;
input n_161;
input n_68;
input n_166;
input n_28;
input n_184;
input n_50;
input n_158;
input n_49;
input n_7;
input n_83;
input n_5;
input n_101;
input n_167;
input n_144;
input n_174;
input n_127;
input n_125;
input n_153;
input n_168;
input n_178;
input n_77;
input n_156;
input n_149;
input n_152;
input n_106;
input n_92;
input n_145;
input n_42;
input n_133;
input n_96;
input n_8;
input n_90;
input n_160;
input n_24;
input n_105;
input n_131;
input n_54;
input n_132;
input n_188;
input n_102;
input n_186;
input n_0;
input n_87;
input n_189;
input n_32;
input n_66;
input n_85;
input n_99;
input n_78;
input n_84;
input n_130;
input n_164;
input n_100;
input n_129;
input n_13;
input n_121;
input n_11;
input n_137;
input n_17;
input n_23;
input n_142;
input n_20;
input n_143;
input n_2;
input n_180;
input n_19;
input n_47;
input n_62;
input n_29;
input n_155;
input n_75;
input n_109;
input n_150;
input n_122;
input n_45;
input n_34;
input n_140;
input n_70;
input n_120;
input n_37;
input n_15;
input n_67;
input n_33;
input n_82;
input n_27;
input n_38;
input n_110;
input n_151;
input n_61;
input n_112;
input n_172;
input n_81;
input n_59;
input n_181;
input n_76;
input n_36;
input n_182;
input n_26;
input n_124;
input n_55;
input n_126;
input n_94;
input n_97;
input n_108;
input n_58;
input n_116;
input n_64;
input n_117;
input n_118;
input n_175;
input n_48;
input n_65;
input n_25;
input n_40;
input n_93;
input n_80;
input n_141;
input n_135;
input n_165;
input n_139;
input n_41;
input n_134;
input n_177;
input n_176;
input n_114;
input n_86;
input n_104;
input n_95;
input n_179;
input n_9;
input n_107;
input n_10;
input n_71;
input n_74;
input n_6;
input n_14;
input n_123;
input n_136;
input n_72;
input n_187;
input n_89;
input n_173;
input n_103;
input n_111;
input n_60;
input n_159;
input n_157;
input n_162;
input n_170;
input n_185;
input n_35;
input n_183;
input n_115;
input n_12;
input n_69;
input n_128;
input n_30;
input n_79;
input n_43;
input n_171;
input n_31;
input n_57;
input n_169;
input n_53;
input n_51;
input n_44;
input n_56;

output n_981;

wire n_591;
wire n_435;
wire n_793;
wire n_326;
wire n_801;
wire n_256;
wire n_853;
wire n_440;
wire n_587;
wire n_695;
wire n_507;
wire n_968;
wire n_909;
wire n_580;
wire n_762;
wire n_881;
wire n_875;
wire n_209;
wire n_367;
wire n_465;
wire n_680;
wire n_741;
wire n_760;
wire n_590;
wire n_625;
wire n_661;
wire n_223;
wire n_278;
wire n_362;
wire n_341;
wire n_226;
wire n_828;
wire n_208;
wire n_462;
wire n_671;
wire n_726;
wire n_607;
wire n_316;
wire n_419;
wire n_304;
wire n_212;
wire n_700;
wire n_694;
wire n_933;
wire n_740;
wire n_578;
wire n_703;
wire n_365;
wire n_978;
wire n_384;
wire n_297;
wire n_595;
wire n_627;
wire n_524;
wire n_342;
wire n_820;
wire n_951;
wire n_783;
wire n_725;
wire n_952;
wire n_358;
wire n_751;
wire n_449;
wire n_749;
wire n_798;
wire n_310;
wire n_509;
wire n_245;
wire n_368;
wire n_575;
wire n_677;
wire n_969;
wire n_805;
wire n_396;
wire n_495;
wire n_815;
wire n_350;
wire n_585;
wire n_732;
wire n_974;
wire n_568;
wire n_392;
wire n_840;
wire n_442;
wire n_480;
wire n_874;
wire n_724;
wire n_382;
wire n_673;
wire n_628;
wire n_883;
wire n_557;
wire n_823;
wire n_349;
wire n_643;
wire n_233;
wire n_617;
wire n_698;
wire n_898;
wire n_845;
wire n_255;
wire n_807;
wire n_739;
wire n_400;
wire n_284;
wire n_955;
wire n_337;
wire n_865;
wire n_893;
wire n_214;
wire n_925;
wire n_485;
wire n_443;
wire n_246;
wire n_892;
wire n_768;
wire n_471;
wire n_289;
wire n_935;
wire n_421;
wire n_781;
wire n_424;
wire n_789;
wire n_615;
wire n_238;
wire n_573;
wire n_769;
wire n_202;
wire n_320;
wire n_639;
wire n_676;
wire n_327;
wire n_794;
wire n_963;
wire n_727;
wire n_894;
wire n_369;
wire n_597;
wire n_685;
wire n_280;
wire n_287;
wire n_832;
wire n_353;
wire n_610;
wire n_555;
wire n_389;
wire n_814;
wire n_415;
wire n_830;
wire n_230;
wire n_605;
wire n_461;
wire n_873;
wire n_383;
wire n_826;
wire n_669;
wire n_200;
wire n_447;
wire n_872;
wire n_198;
wire n_300;
wire n_222;
wire n_718;
wire n_248;
wire n_517;
wire n_747;
wire n_852;
wire n_667;
wire n_229;
wire n_542;
wire n_847;
wire n_644;
wire n_682;
wire n_851;
wire n_621;
wire n_305;
wire n_721;
wire n_750;
wire n_742;
wire n_532;
wire n_535;
wire n_691;
wire n_250;
wire n_372;
wire n_468;
wire n_544;
wire n_901;
wire n_504;
wire n_923;
wire n_314;
wire n_378;
wire n_413;
wire n_377;
wire n_791;
wire n_510;
wire n_837;
wire n_836;
wire n_863;
wire n_375;
wire n_601;
wire n_338;
wire n_522;
wire n_948;
wire n_466;
wire n_704;
wire n_918;
wire n_748;
wire n_506;
wire n_763;
wire n_360;
wire n_945;
wire n_977;
wire n_603;
wire n_957;
wire n_235;
wire n_536;
wire n_895;
wire n_866;
wire n_622;
wire n_191;
wire n_340;
wire n_710;
wire n_387;
wire n_452;
wire n_616;
wire n_658;
wire n_744;
wire n_971;
wire n_946;
wire n_344;
wire n_581;
wire n_428;
wire n_761;
wire n_785;
wire n_746;
wire n_609;
wire n_765;
wire n_432;
wire n_641;
wire n_822;
wire n_693;
wire n_631;
wire n_516;
wire n_720;
wire n_758;
wire n_842;
wire n_525;
wire n_611;
wire n_943;
wire n_491;
wire n_878;
wire n_656;
wire n_772;
wire n_843;
wire n_797;
wire n_666;
wire n_371;
wire n_795;
wire n_770;
wire n_940;
wire n_567;
wire n_899;
wire n_738;
wire n_405;
wire n_213;
wire n_538;
wire n_294;
wire n_302;
wire n_499;
wire n_380;
wire n_838;
wire n_705;
wire n_647;
wire n_197;
wire n_844;
wire n_343;
wire n_448;
wire n_886;
wire n_953;
wire n_494;
wire n_539;
wire n_493;
wire n_397;
wire n_614;
wire n_529;
wire n_445;
wire n_425;
wire n_684;
wire n_930;
wire n_888;
wire n_454;
wire n_218;
wire n_638;
wire n_234;
wire n_910;
wire n_486;
wire n_911;
wire n_381;
wire n_947;
wire n_236;
wire n_653;
wire n_887;
wire n_752;
wire n_908;
wire n_944;
wire n_713;
wire n_648;
wire n_657;
wire n_576;
wire n_472;
wire n_270;
wire n_239;
wire n_414;
wire n_563;
wire n_782;
wire n_976;
wire n_490;
wire n_803;
wire n_290;
wire n_220;
wire n_809;
wire n_224;
wire n_926;
wire n_927;
wire n_839;
wire n_734;
wire n_708;
wire n_196;
wire n_919;
wire n_402;
wire n_352;
wire n_917;
wire n_668;
wire n_478;
wire n_626;
wire n_574;
wire n_779;
wire n_800;
wire n_929;
wire n_460;
wire n_907;
wire n_854;
wire n_417;
wire n_446;
wire n_498;
wire n_662;
wire n_374;
wire n_659;
wire n_709;
wire n_870;
wire n_366;
wire n_904;
wire n_777;
wire n_407;
wire n_913;
wire n_450;
wire n_808;
wire n_867;
wire n_272;
wire n_526;
wire n_921;
wire n_712;
wire n_348;
wire n_711;
wire n_579;
wire n_376;
wire n_937;
wire n_390;
wire n_473;
wire n_293;
wire n_334;
wire n_559;
wire n_370;
wire n_458;
wire n_232;
wire n_650;
wire n_717;
wire n_330;
wire n_771;
wire n_470;
wire n_475;
wire n_924;
wire n_298;
wire n_492;
wire n_972;
wire n_281;
wire n_258;
wire n_551;
wire n_699;
wire n_456;
wire n_564;
wire n_260;
wire n_265;
wire n_313;
wire n_451;
wire n_624;
wire n_824;
wire n_962;
wire n_279;
wire n_686;
wire n_796;
wire n_252;
wire n_757;
wire n_228;
wire n_594;
wire n_565;
wire n_719;
wire n_356;
wire n_577;
wire n_936;
wire n_552;
wire n_619;
wire n_885;
wire n_216;
wire n_455;
wire n_896;
wire n_521;
wire n_363;
wire n_572;
wire n_912;
wire n_395;
wire n_813;
wire n_592;
wire n_745;
wire n_654;
wire n_323;
wire n_829;
wire n_606;
wire n_393;
wire n_818;
wire n_411;
wire n_503;
wire n_716;
wire n_623;
wire n_884;
wire n_599;
wire n_513;
wire n_855;
wire n_776;
wire n_321;
wire n_645;
wire n_331;
wire n_916;
wire n_227;
wire n_868;
wire n_570;
wire n_731;
wire n_859;
wire n_406;
wire n_483;
wire n_735;
wire n_204;
wire n_482;
wire n_934;
wire n_755;
wire n_931;
wire n_474;
wire n_608;
wire n_261;
wire n_683;
wire n_620;
wire n_420;
wire n_527;
wire n_630;
wire n_312;
wire n_394;
wire n_519;
wire n_541;
wire n_512;
wire n_958;
wire n_292;
wire n_307;
wire n_469;
wire n_433;
wire n_500;
wire n_942;
wire n_792;
wire n_880;
wire n_476;
wire n_714;
wire n_291;
wire n_219;
wire n_543;
wire n_889;
wire n_357;
wire n_264;
wire n_263;
wire n_589;
wire n_860;
wire n_481;
wire n_788;
wire n_819;
wire n_939;
wire n_821;
wire n_325;
wire n_938;
wire n_767;
wire n_804;
wire n_329;
wire n_600;
wire n_464;
wire n_831;
wire n_802;
wire n_964;
wire n_561;
wire n_477;
wire n_549;
wire n_980;
wire n_533;
wire n_954;
wire n_408;
wire n_932;
wire n_806;
wire n_864;
wire n_879;
wire n_959;
wire n_237;
wire n_584;
wire n_244;
wire n_399;
wire n_243;
wire n_979;
wire n_548;
wire n_905;
wire n_282;
wire n_436;
wire n_833;
wire n_211;
wire n_523;
wire n_322;
wire n_707;
wire n_345;
wire n_409;
wire n_231;
wire n_354;
wire n_689;
wire n_799;
wire n_505;
wire n_240;
wire n_756;
wire n_319;
wire n_547;
wire n_537;
wire n_273;
wire n_558;
wire n_810;
wire n_635;
wire n_787;
wire n_311;
wire n_403;
wire n_723;
wire n_253;
wire n_634;
wire n_583;
wire n_596;
wire n_966;
wire n_546;
wire n_562;
wire n_249;
wire n_201;
wire n_386;
wire n_764;
wire n_556;
wire n_692;
wire n_733;
wire n_754;
wire n_941;
wire n_975;
wire n_487;
wire n_550;
wire n_241;
wire n_275;
wire n_553;
wire n_652;
wire n_849;
wire n_970;
wire n_560;
wire n_753;
wire n_642;
wire n_276;
wire n_569;
wire n_441;
wire n_221;
wire n_811;
wire n_882;
wire n_444;
wire n_586;
wire n_423;
wire n_737;
wire n_318;
wire n_303;
wire n_511;
wire n_715;
wire n_467;
wire n_306;
wire n_193;
wire n_269;
wire n_359;
wire n_973;
wire n_346;
wire n_416;
wire n_530;
wire n_277;
wire n_520;
wire n_418;
wire n_618;
wire n_790;
wire n_582;
wire n_199;
wire n_266;
wire n_296;
wire n_861;
wire n_674;
wire n_857;
wire n_871;
wire n_967;
wire n_775;
wire n_922;
wire n_571;
wire n_268;
wire n_271;
wire n_404;
wire n_651;
wire n_439;
wire n_217;
wire n_210;
wire n_299;
wire n_518;
wire n_206;
wire n_679;
wire n_453;
wire n_612;
wire n_633;
wire n_665;
wire n_902;
wire n_333;
wire n_588;
wire n_215;
wire n_247;
wire n_225;
wire n_308;
wire n_309;
wire n_914;
wire n_759;
wire n_355;
wire n_426;
wire n_317;
wire n_915;
wire n_632;
wire n_702;
wire n_431;
wire n_347;
wire n_812;
wire n_459;
wire n_502;
wire n_328;
wire n_672;
wire n_534;
wire n_488;
wire n_429;
wire n_373;
wire n_195;
wire n_497;
wire n_285;
wire n_780;
wire n_773;
wire n_675;
wire n_903;
wire n_257;
wire n_920;
wire n_730;
wire n_655;
wire n_706;
wire n_786;
wire n_670;
wire n_203;
wire n_286;
wire n_254;
wire n_207;
wire n_834;
wire n_242;
wire n_835;
wire n_928;
wire n_690;
wire n_850;
wire n_401;
wire n_324;
wire n_766;
wire n_743;
wire n_816;
wire n_335;
wire n_430;
wire n_463;
wire n_545;
wire n_489;
wire n_877;
wire n_205;
wire n_604;
wire n_848;
wire n_251;
wire n_301;
wire n_274;
wire n_636;
wire n_825;
wire n_728;
wire n_681;
wire n_729;
wire n_876;
wire n_774;
wire n_412;
wire n_640;
wire n_660;
wire n_965;
wire n_267;
wire n_438;
wire n_339;
wire n_784;
wire n_434;
wire n_315;
wire n_515;
wire n_288;
wire n_427;
wire n_479;
wire n_598;
wire n_496;
wire n_422;
wire n_696;
wire n_906;
wire n_688;
wire n_722;
wire n_961;
wire n_862;
wire n_869;
wire n_351;
wire n_437;
wire n_259;
wire n_540;
wire n_593;
wire n_514;
wire n_646;
wire n_528;
wire n_457;
wire n_391;
wire n_687;
wire n_697;
wire n_364;
wire n_890;
wire n_637;
wire n_295;
wire n_385;
wire n_701;
wire n_817;
wire n_950;
wire n_629;
wire n_388;
wire n_190;
wire n_858;
wire n_262;
wire n_484;
wire n_613;
wire n_736;
wire n_897;
wire n_900;
wire n_846;
wire n_501;
wire n_841;
wire n_956;
wire n_960;
wire n_531;
wire n_827;
wire n_361;
wire n_508;
wire n_663;
wire n_856;
wire n_379;
wire n_778;
wire n_332;
wire n_891;
wire n_336;
wire n_410;
wire n_398;
wire n_566;
wire n_554;
wire n_602;
wire n_194;
wire n_664;
wire n_949;
wire n_678;
wire n_192;
wire n_649;
wire n_283;

CKINVDCx5p33_ASAP7_75t_R g190 ( 
.A(n_171),
.Y(n_190)
);

CKINVDCx5p33_ASAP7_75t_R g191 ( 
.A(n_133),
.Y(n_191)
);

CKINVDCx5p33_ASAP7_75t_R g192 ( 
.A(n_186),
.Y(n_192)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_105),
.Y(n_193)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_129),
.Y(n_194)
);

CKINVDCx5p33_ASAP7_75t_R g195 ( 
.A(n_163),
.Y(n_195)
);

CKINVDCx16_ASAP7_75t_R g196 ( 
.A(n_147),
.Y(n_196)
);

INVx2_ASAP7_75t_L g197 ( 
.A(n_126),
.Y(n_197)
);

INVx1_ASAP7_75t_SL g198 ( 
.A(n_150),
.Y(n_198)
);

CKINVDCx16_ASAP7_75t_R g199 ( 
.A(n_13),
.Y(n_199)
);

CKINVDCx5p33_ASAP7_75t_R g200 ( 
.A(n_178),
.Y(n_200)
);

CKINVDCx5p33_ASAP7_75t_R g201 ( 
.A(n_76),
.Y(n_201)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_56),
.Y(n_202)
);

CKINVDCx5p33_ASAP7_75t_R g203 ( 
.A(n_48),
.Y(n_203)
);

CKINVDCx20_ASAP7_75t_R g204 ( 
.A(n_155),
.Y(n_204)
);

CKINVDCx20_ASAP7_75t_R g205 ( 
.A(n_93),
.Y(n_205)
);

CKINVDCx5p33_ASAP7_75t_R g206 ( 
.A(n_19),
.Y(n_206)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_44),
.Y(n_207)
);

CKINVDCx5p33_ASAP7_75t_R g208 ( 
.A(n_5),
.Y(n_208)
);

CKINVDCx5p33_ASAP7_75t_R g209 ( 
.A(n_91),
.Y(n_209)
);

CKINVDCx20_ASAP7_75t_R g210 ( 
.A(n_54),
.Y(n_210)
);

CKINVDCx5p33_ASAP7_75t_R g211 ( 
.A(n_99),
.Y(n_211)
);

BUFx3_ASAP7_75t_L g212 ( 
.A(n_11),
.Y(n_212)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_162),
.Y(n_213)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_73),
.Y(n_214)
);

CKINVDCx5p33_ASAP7_75t_R g215 ( 
.A(n_117),
.Y(n_215)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_128),
.Y(n_216)
);

CKINVDCx5p33_ASAP7_75t_R g217 ( 
.A(n_4),
.Y(n_217)
);

CKINVDCx5p33_ASAP7_75t_R g218 ( 
.A(n_0),
.Y(n_218)
);

CKINVDCx5p33_ASAP7_75t_R g219 ( 
.A(n_113),
.Y(n_219)
);

CKINVDCx5p33_ASAP7_75t_R g220 ( 
.A(n_119),
.Y(n_220)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_106),
.Y(n_221)
);

INVx2_ASAP7_75t_L g222 ( 
.A(n_45),
.Y(n_222)
);

CKINVDCx5p33_ASAP7_75t_R g223 ( 
.A(n_176),
.Y(n_223)
);

BUFx3_ASAP7_75t_L g224 ( 
.A(n_71),
.Y(n_224)
);

CKINVDCx5p33_ASAP7_75t_R g225 ( 
.A(n_185),
.Y(n_225)
);

CKINVDCx14_ASAP7_75t_R g226 ( 
.A(n_86),
.Y(n_226)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_77),
.Y(n_227)
);

BUFx2_ASAP7_75t_SL g228 ( 
.A(n_121),
.Y(n_228)
);

CKINVDCx5p33_ASAP7_75t_R g229 ( 
.A(n_85),
.Y(n_229)
);

CKINVDCx5p33_ASAP7_75t_R g230 ( 
.A(n_154),
.Y(n_230)
);

BUFx3_ASAP7_75t_L g231 ( 
.A(n_35),
.Y(n_231)
);

HB1xp67_ASAP7_75t_L g232 ( 
.A(n_90),
.Y(n_232)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_120),
.Y(n_233)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_5),
.Y(n_234)
);

INVx2_ASAP7_75t_L g235 ( 
.A(n_27),
.Y(n_235)
);

BUFx3_ASAP7_75t_L g236 ( 
.A(n_34),
.Y(n_236)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_167),
.Y(n_237)
);

CKINVDCx5p33_ASAP7_75t_R g238 ( 
.A(n_7),
.Y(n_238)
);

CKINVDCx5p33_ASAP7_75t_R g239 ( 
.A(n_123),
.Y(n_239)
);

CKINVDCx5p33_ASAP7_75t_R g240 ( 
.A(n_166),
.Y(n_240)
);

CKINVDCx5p33_ASAP7_75t_R g241 ( 
.A(n_25),
.Y(n_241)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_64),
.Y(n_242)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_18),
.Y(n_243)
);

INVx2_ASAP7_75t_L g244 ( 
.A(n_144),
.Y(n_244)
);

CKINVDCx20_ASAP7_75t_R g245 ( 
.A(n_78),
.Y(n_245)
);

CKINVDCx5p33_ASAP7_75t_R g246 ( 
.A(n_125),
.Y(n_246)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_40),
.Y(n_247)
);

CKINVDCx5p33_ASAP7_75t_R g248 ( 
.A(n_39),
.Y(n_248)
);

CKINVDCx5p33_ASAP7_75t_R g249 ( 
.A(n_189),
.Y(n_249)
);

CKINVDCx20_ASAP7_75t_R g250 ( 
.A(n_100),
.Y(n_250)
);

CKINVDCx5p33_ASAP7_75t_R g251 ( 
.A(n_160),
.Y(n_251)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_110),
.Y(n_252)
);

CKINVDCx5p33_ASAP7_75t_R g253 ( 
.A(n_1),
.Y(n_253)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_49),
.Y(n_254)
);

CKINVDCx5p33_ASAP7_75t_R g255 ( 
.A(n_188),
.Y(n_255)
);

INVx4_ASAP7_75t_R g256 ( 
.A(n_65),
.Y(n_256)
);

CKINVDCx5p33_ASAP7_75t_R g257 ( 
.A(n_169),
.Y(n_257)
);

BUFx6f_ASAP7_75t_L g258 ( 
.A(n_43),
.Y(n_258)
);

CKINVDCx5p33_ASAP7_75t_R g259 ( 
.A(n_28),
.Y(n_259)
);

CKINVDCx5p33_ASAP7_75t_R g260 ( 
.A(n_34),
.Y(n_260)
);

CKINVDCx20_ASAP7_75t_R g261 ( 
.A(n_41),
.Y(n_261)
);

CKINVDCx5p33_ASAP7_75t_R g262 ( 
.A(n_15),
.Y(n_262)
);

BUFx3_ASAP7_75t_L g263 ( 
.A(n_24),
.Y(n_263)
);

CKINVDCx20_ASAP7_75t_R g264 ( 
.A(n_177),
.Y(n_264)
);

CKINVDCx5p33_ASAP7_75t_R g265 ( 
.A(n_13),
.Y(n_265)
);

INVx2_ASAP7_75t_L g266 ( 
.A(n_173),
.Y(n_266)
);

CKINVDCx5p33_ASAP7_75t_R g267 ( 
.A(n_55),
.Y(n_267)
);

CKINVDCx5p33_ASAP7_75t_R g268 ( 
.A(n_7),
.Y(n_268)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_170),
.Y(n_269)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_175),
.Y(n_270)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_142),
.Y(n_271)
);

CKINVDCx5p33_ASAP7_75t_R g272 ( 
.A(n_33),
.Y(n_272)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_148),
.Y(n_273)
);

CKINVDCx20_ASAP7_75t_R g274 ( 
.A(n_67),
.Y(n_274)
);

BUFx12f_ASAP7_75t_L g275 ( 
.A(n_253),
.Y(n_275)
);

INVx5_ASAP7_75t_L g276 ( 
.A(n_258),
.Y(n_276)
);

NOR2xp33_ASAP7_75t_L g277 ( 
.A(n_232),
.B(n_0),
.Y(n_277)
);

NAND2xp5_ASAP7_75t_L g278 ( 
.A(n_197),
.B(n_1),
.Y(n_278)
);

AND2x2_ASAP7_75t_L g279 ( 
.A(n_212),
.B(n_2),
.Y(n_279)
);

AND2x4_ASAP7_75t_L g280 ( 
.A(n_224),
.B(n_2),
.Y(n_280)
);

BUFx12f_ASAP7_75t_L g281 ( 
.A(n_253),
.Y(n_281)
);

AND2x4_ASAP7_75t_L g282 ( 
.A(n_224),
.B(n_3),
.Y(n_282)
);

AND2x4_ASAP7_75t_L g283 ( 
.A(n_197),
.B(n_3),
.Y(n_283)
);

INVx5_ASAP7_75t_L g284 ( 
.A(n_258),
.Y(n_284)
);

BUFx6f_ASAP7_75t_L g285 ( 
.A(n_258),
.Y(n_285)
);

AND2x4_ASAP7_75t_L g286 ( 
.A(n_222),
.B(n_4),
.Y(n_286)
);

INVx5_ASAP7_75t_L g287 ( 
.A(n_258),
.Y(n_287)
);

BUFx6f_ASAP7_75t_L g288 ( 
.A(n_258),
.Y(n_288)
);

BUFx6f_ASAP7_75t_L g289 ( 
.A(n_222),
.Y(n_289)
);

CKINVDCx20_ASAP7_75t_R g290 ( 
.A(n_199),
.Y(n_290)
);

NAND2xp5_ASAP7_75t_L g291 ( 
.A(n_244),
.B(n_266),
.Y(n_291)
);

BUFx3_ASAP7_75t_L g292 ( 
.A(n_193),
.Y(n_292)
);

BUFx6f_ASAP7_75t_L g293 ( 
.A(n_244),
.Y(n_293)
);

CKINVDCx5p33_ASAP7_75t_R g294 ( 
.A(n_209),
.Y(n_294)
);

INVxp67_ASAP7_75t_L g295 ( 
.A(n_234),
.Y(n_295)
);

BUFx8_ASAP7_75t_SL g296 ( 
.A(n_259),
.Y(n_296)
);

INVx3_ASAP7_75t_L g297 ( 
.A(n_212),
.Y(n_297)
);

NOR2xp33_ASAP7_75t_L g298 ( 
.A(n_198),
.B(n_6),
.Y(n_298)
);

INVx5_ASAP7_75t_L g299 ( 
.A(n_196),
.Y(n_299)
);

INVxp67_ASAP7_75t_L g300 ( 
.A(n_243),
.Y(n_300)
);

BUFx6f_ASAP7_75t_L g301 ( 
.A(n_266),
.Y(n_301)
);

NAND2xp5_ASAP7_75t_L g302 ( 
.A(n_226),
.B(n_6),
.Y(n_302)
);

AND2x4_ASAP7_75t_L g303 ( 
.A(n_194),
.B(n_8),
.Y(n_303)
);

AND2x6_ASAP7_75t_L g304 ( 
.A(n_202),
.B(n_42),
.Y(n_304)
);

AND2x4_ASAP7_75t_L g305 ( 
.A(n_207),
.B(n_8),
.Y(n_305)
);

NAND2xp5_ASAP7_75t_L g306 ( 
.A(n_213),
.B(n_9),
.Y(n_306)
);

BUFx6f_ASAP7_75t_L g307 ( 
.A(n_214),
.Y(n_307)
);

BUFx12f_ASAP7_75t_L g308 ( 
.A(n_259),
.Y(n_308)
);

INVxp67_ASAP7_75t_L g309 ( 
.A(n_231),
.Y(n_309)
);

XNOR2xp5_ASAP7_75t_L g310 ( 
.A(n_260),
.B(n_9),
.Y(n_310)
);

NAND2xp5_ASAP7_75t_L g311 ( 
.A(n_216),
.B(n_221),
.Y(n_311)
);

INVx5_ASAP7_75t_L g312 ( 
.A(n_231),
.Y(n_312)
);

BUFx6f_ASAP7_75t_L g313 ( 
.A(n_227),
.Y(n_313)
);

BUFx6f_ASAP7_75t_L g314 ( 
.A(n_233),
.Y(n_314)
);

BUFx6f_ASAP7_75t_L g315 ( 
.A(n_237),
.Y(n_315)
);

BUFx6f_ASAP7_75t_L g316 ( 
.A(n_242),
.Y(n_316)
);

NAND2xp5_ASAP7_75t_L g317 ( 
.A(n_247),
.B(n_10),
.Y(n_317)
);

BUFx3_ASAP7_75t_L g318 ( 
.A(n_252),
.Y(n_318)
);

NAND2xp5_ASAP7_75t_L g319 ( 
.A(n_254),
.B(n_10),
.Y(n_319)
);

AND2x6_ASAP7_75t_L g320 ( 
.A(n_269),
.B(n_46),
.Y(n_320)
);

NOR2xp33_ASAP7_75t_SL g321 ( 
.A(n_236),
.B(n_263),
.Y(n_321)
);

AND2x2_ASAP7_75t_L g322 ( 
.A(n_236),
.B(n_11),
.Y(n_322)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_263),
.Y(n_323)
);

BUFx12f_ASAP7_75t_L g324 ( 
.A(n_260),
.Y(n_324)
);

BUFx2_ASAP7_75t_L g325 ( 
.A(n_262),
.Y(n_325)
);

INVx5_ASAP7_75t_L g326 ( 
.A(n_235),
.Y(n_326)
);

BUFx12f_ASAP7_75t_L g327 ( 
.A(n_262),
.Y(n_327)
);

INVx2_ASAP7_75t_L g328 ( 
.A(n_235),
.Y(n_328)
);

NOR2xp33_ASAP7_75t_L g329 ( 
.A(n_299),
.B(n_190),
.Y(n_329)
);

AOI22xp5_ASAP7_75t_L g330 ( 
.A1(n_290),
.A2(n_265),
.B1(n_204),
.B2(n_210),
.Y(n_330)
);

OR2x6_ASAP7_75t_L g331 ( 
.A(n_324),
.B(n_228),
.Y(n_331)
);

AOI22xp5_ASAP7_75t_L g332 ( 
.A1(n_290),
.A2(n_265),
.B1(n_205),
.B2(n_261),
.Y(n_332)
);

OAI22xp33_ASAP7_75t_L g333 ( 
.A1(n_321),
.A2(n_302),
.B1(n_278),
.B2(n_325),
.Y(n_333)
);

INVx2_ASAP7_75t_L g334 ( 
.A(n_285),
.Y(n_334)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_289),
.Y(n_335)
);

AND2x2_ASAP7_75t_L g336 ( 
.A(n_299),
.B(n_190),
.Y(n_336)
);

INVx2_ASAP7_75t_SL g337 ( 
.A(n_275),
.Y(n_337)
);

AO22x2_ASAP7_75t_L g338 ( 
.A1(n_280),
.A2(n_270),
.B1(n_271),
.B2(n_273),
.Y(n_338)
);

OAI22xp33_ASAP7_75t_L g339 ( 
.A1(n_306),
.A2(n_217),
.B1(n_272),
.B2(n_268),
.Y(n_339)
);

AOI22xp5_ASAP7_75t_L g340 ( 
.A1(n_277),
.A2(n_274),
.B1(n_245),
.B2(n_264),
.Y(n_340)
);

BUFx6f_ASAP7_75t_L g341 ( 
.A(n_289),
.Y(n_341)
);

OAI22xp33_ASAP7_75t_SL g342 ( 
.A1(n_277),
.A2(n_248),
.B1(n_208),
.B2(n_238),
.Y(n_342)
);

OAI22xp5_ASAP7_75t_L g343 ( 
.A1(n_298),
.A2(n_218),
.B1(n_206),
.B2(n_241),
.Y(n_343)
);

OAI22xp5_ASAP7_75t_SL g344 ( 
.A1(n_310),
.A2(n_250),
.B1(n_257),
.B2(n_255),
.Y(n_344)
);

OAI22xp33_ASAP7_75t_SL g345 ( 
.A1(n_280),
.A2(n_191),
.B1(n_257),
.B2(n_192),
.Y(n_345)
);

AOI22xp5_ASAP7_75t_L g346 ( 
.A1(n_298),
.A2(n_191),
.B1(n_192),
.B2(n_255),
.Y(n_346)
);

INVx1_ASAP7_75t_L g347 ( 
.A(n_289),
.Y(n_347)
);

OA22x2_ASAP7_75t_L g348 ( 
.A1(n_309),
.A2(n_195),
.B1(n_251),
.B2(n_200),
.Y(n_348)
);

AND2x2_ASAP7_75t_L g349 ( 
.A(n_299),
.B(n_195),
.Y(n_349)
);

INVx2_ASAP7_75t_L g350 ( 
.A(n_285),
.Y(n_350)
);

INVx1_ASAP7_75t_L g351 ( 
.A(n_289),
.Y(n_351)
);

AO22x2_ASAP7_75t_L g352 ( 
.A1(n_282),
.A2(n_256),
.B1(n_14),
.B2(n_15),
.Y(n_352)
);

OAI22xp33_ASAP7_75t_SL g353 ( 
.A1(n_282),
.A2(n_200),
.B1(n_251),
.B2(n_201),
.Y(n_353)
);

INVx1_ASAP7_75t_L g354 ( 
.A(n_293),
.Y(n_354)
);

NOR2xp33_ASAP7_75t_L g355 ( 
.A(n_299),
.B(n_201),
.Y(n_355)
);

AND2x2_ASAP7_75t_L g356 ( 
.A(n_294),
.B(n_203),
.Y(n_356)
);

AOI22xp5_ASAP7_75t_L g357 ( 
.A1(n_283),
.A2(n_203),
.B1(n_249),
.B2(n_246),
.Y(n_357)
);

OAI22xp33_ASAP7_75t_L g358 ( 
.A1(n_317),
.A2(n_267),
.B1(n_240),
.B2(n_239),
.Y(n_358)
);

INVx1_ASAP7_75t_L g359 ( 
.A(n_293),
.Y(n_359)
);

OAI22xp33_ASAP7_75t_SL g360 ( 
.A1(n_291),
.A2(n_230),
.B1(n_229),
.B2(n_225),
.Y(n_360)
);

OAI22xp5_ASAP7_75t_SL g361 ( 
.A1(n_275),
.A2(n_223),
.B1(n_220),
.B2(n_219),
.Y(n_361)
);

AND2x2_ASAP7_75t_L g362 ( 
.A(n_309),
.B(n_211),
.Y(n_362)
);

OAI22xp33_ASAP7_75t_L g363 ( 
.A1(n_319),
.A2(n_215),
.B1(n_14),
.B2(n_16),
.Y(n_363)
);

INVx2_ASAP7_75t_L g364 ( 
.A(n_285),
.Y(n_364)
);

AOI22xp5_ASAP7_75t_L g365 ( 
.A1(n_283),
.A2(n_12),
.B1(n_16),
.B2(n_17),
.Y(n_365)
);

INVx1_ASAP7_75t_L g366 ( 
.A(n_293),
.Y(n_366)
);

OR2x6_ASAP7_75t_L g367 ( 
.A(n_281),
.B(n_12),
.Y(n_367)
);

NAND2xp5_ASAP7_75t_L g368 ( 
.A(n_312),
.B(n_47),
.Y(n_368)
);

NAND2xp5_ASAP7_75t_SL g369 ( 
.A(n_286),
.B(n_312),
.Y(n_369)
);

INVx2_ASAP7_75t_SL g370 ( 
.A(n_281),
.Y(n_370)
);

AOI22xp5_ASAP7_75t_L g371 ( 
.A1(n_308),
.A2(n_327),
.B1(n_303),
.B2(n_305),
.Y(n_371)
);

INVx1_ASAP7_75t_L g372 ( 
.A(n_293),
.Y(n_372)
);

NOR2xp33_ASAP7_75t_L g373 ( 
.A(n_311),
.B(n_17),
.Y(n_373)
);

AND2x2_ASAP7_75t_L g374 ( 
.A(n_297),
.B(n_50),
.Y(n_374)
);

OAI22xp33_ASAP7_75t_L g375 ( 
.A1(n_308),
.A2(n_327),
.B1(n_295),
.B2(n_300),
.Y(n_375)
);

INVx1_ASAP7_75t_L g376 ( 
.A(n_301),
.Y(n_376)
);

OAI22xp33_ASAP7_75t_L g377 ( 
.A1(n_295),
.A2(n_18),
.B1(n_19),
.B2(n_20),
.Y(n_377)
);

AND2x2_ASAP7_75t_L g378 ( 
.A(n_297),
.B(n_51),
.Y(n_378)
);

NOR2xp33_ASAP7_75t_L g379 ( 
.A(n_303),
.B(n_20),
.Y(n_379)
);

INVx2_ASAP7_75t_L g380 ( 
.A(n_285),
.Y(n_380)
);

INVx2_ASAP7_75t_L g381 ( 
.A(n_288),
.Y(n_381)
);

OAI22xp33_ASAP7_75t_L g382 ( 
.A1(n_300),
.A2(n_21),
.B1(n_22),
.B2(n_23),
.Y(n_382)
);

INVx1_ASAP7_75t_L g383 ( 
.A(n_301),
.Y(n_383)
);

AO22x2_ASAP7_75t_L g384 ( 
.A1(n_286),
.A2(n_21),
.B1(n_22),
.B2(n_23),
.Y(n_384)
);

INVx2_ASAP7_75t_SL g385 ( 
.A(n_362),
.Y(n_385)
);

AND2x2_ASAP7_75t_SL g386 ( 
.A(n_365),
.B(n_305),
.Y(n_386)
);

INVx2_ASAP7_75t_L g387 ( 
.A(n_334),
.Y(n_387)
);

INVx1_ASAP7_75t_L g388 ( 
.A(n_335),
.Y(n_388)
);

INVx1_ASAP7_75t_L g389 ( 
.A(n_347),
.Y(n_389)
);

INVx1_ASAP7_75t_L g390 ( 
.A(n_351),
.Y(n_390)
);

INVx1_ASAP7_75t_L g391 ( 
.A(n_354),
.Y(n_391)
);

CKINVDCx20_ASAP7_75t_R g392 ( 
.A(n_330),
.Y(n_392)
);

INVx2_ASAP7_75t_L g393 ( 
.A(n_350),
.Y(n_393)
);

NOR2xp33_ASAP7_75t_L g394 ( 
.A(n_346),
.B(n_312),
.Y(n_394)
);

NAND2xp5_ASAP7_75t_L g395 ( 
.A(n_336),
.B(n_276),
.Y(n_395)
);

INVx1_ASAP7_75t_L g396 ( 
.A(n_359),
.Y(n_396)
);

INVx1_ASAP7_75t_L g397 ( 
.A(n_366),
.Y(n_397)
);

INVx1_ASAP7_75t_L g398 ( 
.A(n_372),
.Y(n_398)
);

XOR2xp5_ASAP7_75t_L g399 ( 
.A(n_330),
.B(n_52),
.Y(n_399)
);

OR2x6_ASAP7_75t_L g400 ( 
.A(n_384),
.B(n_323),
.Y(n_400)
);

INVx1_ASAP7_75t_L g401 ( 
.A(n_376),
.Y(n_401)
);

NAND2xp5_ASAP7_75t_L g402 ( 
.A(n_349),
.B(n_276),
.Y(n_402)
);

AND2x4_ASAP7_75t_L g403 ( 
.A(n_369),
.B(n_328),
.Y(n_403)
);

INVx1_ASAP7_75t_L g404 ( 
.A(n_383),
.Y(n_404)
);

INVx1_ASAP7_75t_L g405 ( 
.A(n_364),
.Y(n_405)
);

NOR2xp33_ASAP7_75t_L g406 ( 
.A(n_346),
.B(n_312),
.Y(n_406)
);

INVx1_ASAP7_75t_L g407 ( 
.A(n_380),
.Y(n_407)
);

INVx1_ASAP7_75t_L g408 ( 
.A(n_381),
.Y(n_408)
);

XNOR2x2_ASAP7_75t_L g409 ( 
.A(n_384),
.B(n_279),
.Y(n_409)
);

INVx1_ASAP7_75t_L g410 ( 
.A(n_341),
.Y(n_410)
);

HB1xp67_ASAP7_75t_L g411 ( 
.A(n_348),
.Y(n_411)
);

AND2x4_ASAP7_75t_L g412 ( 
.A(n_374),
.B(n_328),
.Y(n_412)
);

INVx1_ASAP7_75t_L g413 ( 
.A(n_341),
.Y(n_413)
);

INVx1_ASAP7_75t_L g414 ( 
.A(n_341),
.Y(n_414)
);

INVx1_ASAP7_75t_L g415 ( 
.A(n_378),
.Y(n_415)
);

NOR2xp33_ASAP7_75t_SL g416 ( 
.A(n_337),
.B(n_296),
.Y(n_416)
);

CKINVDCx20_ASAP7_75t_R g417 ( 
.A(n_332),
.Y(n_417)
);

NOR2xp33_ASAP7_75t_L g418 ( 
.A(n_333),
.B(n_357),
.Y(n_418)
);

XNOR2xp5_ASAP7_75t_SL g419 ( 
.A(n_332),
.B(n_296),
.Y(n_419)
);

INVx1_ASAP7_75t_L g420 ( 
.A(n_379),
.Y(n_420)
);

AND2x2_ASAP7_75t_L g421 ( 
.A(n_356),
.B(n_292),
.Y(n_421)
);

INVx1_ASAP7_75t_L g422 ( 
.A(n_338),
.Y(n_422)
);

AND2x2_ASAP7_75t_L g423 ( 
.A(n_357),
.B(n_292),
.Y(n_423)
);

AND2x2_ASAP7_75t_L g424 ( 
.A(n_329),
.B(n_318),
.Y(n_424)
);

AND2x2_ASAP7_75t_L g425 ( 
.A(n_355),
.B(n_318),
.Y(n_425)
);

BUFx2_ASAP7_75t_L g426 ( 
.A(n_367),
.Y(n_426)
);

XOR2xp5_ASAP7_75t_L g427 ( 
.A(n_340),
.B(n_53),
.Y(n_427)
);

AND2x2_ASAP7_75t_L g428 ( 
.A(n_343),
.B(n_322),
.Y(n_428)
);

CKINVDCx20_ASAP7_75t_R g429 ( 
.A(n_344),
.Y(n_429)
);

INVx1_ASAP7_75t_L g430 ( 
.A(n_338),
.Y(n_430)
);

NAND2xp5_ASAP7_75t_SL g431 ( 
.A(n_360),
.B(n_301),
.Y(n_431)
);

INVx1_ASAP7_75t_L g432 ( 
.A(n_373),
.Y(n_432)
);

INVx1_ASAP7_75t_L g433 ( 
.A(n_368),
.Y(n_433)
);

INVx1_ASAP7_75t_L g434 ( 
.A(n_352),
.Y(n_434)
);

INVx1_ASAP7_75t_L g435 ( 
.A(n_352),
.Y(n_435)
);

INVx1_ASAP7_75t_SL g436 ( 
.A(n_361),
.Y(n_436)
);

XOR2xp5_ASAP7_75t_L g437 ( 
.A(n_340),
.B(n_57),
.Y(n_437)
);

INVxp33_ASAP7_75t_L g438 ( 
.A(n_371),
.Y(n_438)
);

XOR2xp5_ASAP7_75t_L g439 ( 
.A(n_342),
.B(n_58),
.Y(n_439)
);

NAND2x1p5_ASAP7_75t_L g440 ( 
.A(n_365),
.B(n_301),
.Y(n_440)
);

INVx2_ASAP7_75t_L g441 ( 
.A(n_367),
.Y(n_441)
);

CKINVDCx20_ASAP7_75t_R g442 ( 
.A(n_331),
.Y(n_442)
);

NOR2xp33_ASAP7_75t_L g443 ( 
.A(n_345),
.B(n_307),
.Y(n_443)
);

BUFx5_ASAP7_75t_L g444 ( 
.A(n_377),
.Y(n_444)
);

XNOR2x2_ASAP7_75t_L g445 ( 
.A(n_382),
.B(n_24),
.Y(n_445)
);

AND2x2_ASAP7_75t_L g446 ( 
.A(n_370),
.B(n_326),
.Y(n_446)
);

INVx1_ASAP7_75t_L g447 ( 
.A(n_353),
.Y(n_447)
);

INVx2_ASAP7_75t_L g448 ( 
.A(n_367),
.Y(n_448)
);

INVx1_ASAP7_75t_L g449 ( 
.A(n_363),
.Y(n_449)
);

NAND2xp33_ASAP7_75t_SL g450 ( 
.A(n_339),
.B(n_307),
.Y(n_450)
);

INVx1_ASAP7_75t_L g451 ( 
.A(n_358),
.Y(n_451)
);

INVx1_ASAP7_75t_L g452 ( 
.A(n_331),
.Y(n_452)
);

INVx1_ASAP7_75t_L g453 ( 
.A(n_331),
.Y(n_453)
);

INVx1_ASAP7_75t_L g454 ( 
.A(n_375),
.Y(n_454)
);

INVx1_ASAP7_75t_L g455 ( 
.A(n_335),
.Y(n_455)
);

CKINVDCx20_ASAP7_75t_R g456 ( 
.A(n_330),
.Y(n_456)
);

INVx1_ASAP7_75t_L g457 ( 
.A(n_335),
.Y(n_457)
);

INVx1_ASAP7_75t_L g458 ( 
.A(n_335),
.Y(n_458)
);

CKINVDCx5p33_ASAP7_75t_R g459 ( 
.A(n_361),
.Y(n_459)
);

AND2x2_ASAP7_75t_L g460 ( 
.A(n_432),
.B(n_420),
.Y(n_460)
);

AND2x6_ASAP7_75t_L g461 ( 
.A(n_434),
.B(n_304),
.Y(n_461)
);

OAI21xp5_ASAP7_75t_L g462 ( 
.A1(n_433),
.A2(n_320),
.B(n_304),
.Y(n_462)
);

NAND2xp5_ASAP7_75t_L g463 ( 
.A(n_412),
.B(n_304),
.Y(n_463)
);

OAI21xp5_ASAP7_75t_L g464 ( 
.A1(n_415),
.A2(n_320),
.B(n_304),
.Y(n_464)
);

INVx4_ASAP7_75t_L g465 ( 
.A(n_412),
.Y(n_465)
);

BUFx4_ASAP7_75t_SL g466 ( 
.A(n_442),
.Y(n_466)
);

NAND2xp5_ASAP7_75t_L g467 ( 
.A(n_412),
.B(n_304),
.Y(n_467)
);

AND2x2_ASAP7_75t_SL g468 ( 
.A(n_386),
.B(n_320),
.Y(n_468)
);

AND2x2_ASAP7_75t_L g469 ( 
.A(n_424),
.B(n_425),
.Y(n_469)
);

INVx2_ASAP7_75t_L g470 ( 
.A(n_387),
.Y(n_470)
);

NAND2xp5_ASAP7_75t_L g471 ( 
.A(n_385),
.B(n_421),
.Y(n_471)
);

AND2x2_ASAP7_75t_L g472 ( 
.A(n_428),
.B(n_307),
.Y(n_472)
);

INVx2_ASAP7_75t_L g473 ( 
.A(n_387),
.Y(n_473)
);

INVx1_ASAP7_75t_L g474 ( 
.A(n_393),
.Y(n_474)
);

NAND2xp5_ASAP7_75t_SL g475 ( 
.A(n_394),
.B(n_307),
.Y(n_475)
);

AND2x2_ASAP7_75t_L g476 ( 
.A(n_423),
.B(n_313),
.Y(n_476)
);

INVx1_ASAP7_75t_SL g477 ( 
.A(n_411),
.Y(n_477)
);

AND2x4_ASAP7_75t_L g478 ( 
.A(n_403),
.B(n_320),
.Y(n_478)
);

AND2x2_ASAP7_75t_L g479 ( 
.A(n_403),
.B(n_440),
.Y(n_479)
);

INVx1_ASAP7_75t_L g480 ( 
.A(n_393),
.Y(n_480)
);

INVx1_ASAP7_75t_SL g481 ( 
.A(n_411),
.Y(n_481)
);

INVx3_ASAP7_75t_SL g482 ( 
.A(n_459),
.Y(n_482)
);

INVx2_ASAP7_75t_L g483 ( 
.A(n_405),
.Y(n_483)
);

AND2x4_ASAP7_75t_L g484 ( 
.A(n_403),
.B(n_320),
.Y(n_484)
);

INVx1_ASAP7_75t_L g485 ( 
.A(n_407),
.Y(n_485)
);

HB1xp67_ASAP7_75t_L g486 ( 
.A(n_440),
.Y(n_486)
);

INVx1_ASAP7_75t_L g487 ( 
.A(n_408),
.Y(n_487)
);

INVx2_ASAP7_75t_L g488 ( 
.A(n_388),
.Y(n_488)
);

INVx2_ASAP7_75t_L g489 ( 
.A(n_458),
.Y(n_489)
);

NAND2xp5_ASAP7_75t_L g490 ( 
.A(n_451),
.B(n_313),
.Y(n_490)
);

OAI21xp5_ASAP7_75t_L g491 ( 
.A1(n_395),
.A2(n_402),
.B(n_394),
.Y(n_491)
);

INVx2_ASAP7_75t_SL g492 ( 
.A(n_431),
.Y(n_492)
);

INVx1_ASAP7_75t_L g493 ( 
.A(n_389),
.Y(n_493)
);

NAND2xp5_ASAP7_75t_L g494 ( 
.A(n_406),
.B(n_313),
.Y(n_494)
);

INVx2_ASAP7_75t_L g495 ( 
.A(n_457),
.Y(n_495)
);

NAND2xp5_ASAP7_75t_SL g496 ( 
.A(n_406),
.B(n_313),
.Y(n_496)
);

INVx2_ASAP7_75t_SL g497 ( 
.A(n_431),
.Y(n_497)
);

NAND2xp5_ASAP7_75t_L g498 ( 
.A(n_390),
.B(n_314),
.Y(n_498)
);

NAND2xp5_ASAP7_75t_SL g499 ( 
.A(n_386),
.B(n_314),
.Y(n_499)
);

BUFx3_ASAP7_75t_L g500 ( 
.A(n_410),
.Y(n_500)
);

AOI22xp5_ASAP7_75t_L g501 ( 
.A1(n_418),
.A2(n_316),
.B1(n_315),
.B2(n_314),
.Y(n_501)
);

NAND2xp5_ASAP7_75t_L g502 ( 
.A(n_391),
.B(n_396),
.Y(n_502)
);

INVx2_ASAP7_75t_L g503 ( 
.A(n_397),
.Y(n_503)
);

NAND2xp5_ASAP7_75t_L g504 ( 
.A(n_398),
.B(n_314),
.Y(n_504)
);

INVx2_ASAP7_75t_L g505 ( 
.A(n_401),
.Y(n_505)
);

INVx3_ASAP7_75t_L g506 ( 
.A(n_404),
.Y(n_506)
);

BUFx3_ASAP7_75t_L g507 ( 
.A(n_413),
.Y(n_507)
);

INVx2_ASAP7_75t_SL g508 ( 
.A(n_422),
.Y(n_508)
);

BUFx6f_ASAP7_75t_L g509 ( 
.A(n_414),
.Y(n_509)
);

HB1xp67_ASAP7_75t_L g510 ( 
.A(n_430),
.Y(n_510)
);

AND2x2_ASAP7_75t_L g511 ( 
.A(n_435),
.B(n_315),
.Y(n_511)
);

CKINVDCx20_ASAP7_75t_R g512 ( 
.A(n_419),
.Y(n_512)
);

INVx1_ASAP7_75t_L g513 ( 
.A(n_455),
.Y(n_513)
);

AND2x2_ASAP7_75t_L g514 ( 
.A(n_443),
.B(n_315),
.Y(n_514)
);

INVx2_ASAP7_75t_L g515 ( 
.A(n_444),
.Y(n_515)
);

INVx1_ASAP7_75t_L g516 ( 
.A(n_443),
.Y(n_516)
);

INVx1_ASAP7_75t_SL g517 ( 
.A(n_392),
.Y(n_517)
);

NAND2xp5_ASAP7_75t_SL g518 ( 
.A(n_418),
.B(n_447),
.Y(n_518)
);

AND2x2_ASAP7_75t_L g519 ( 
.A(n_449),
.B(n_315),
.Y(n_519)
);

NOR2xp33_ASAP7_75t_L g520 ( 
.A(n_438),
.B(n_454),
.Y(n_520)
);

INVx1_ASAP7_75t_SL g521 ( 
.A(n_392),
.Y(n_521)
);

AND2x6_ASAP7_75t_L g522 ( 
.A(n_441),
.B(n_288),
.Y(n_522)
);

NOR2xp33_ASAP7_75t_L g523 ( 
.A(n_438),
.B(n_316),
.Y(n_523)
);

INVx1_ASAP7_75t_L g524 ( 
.A(n_450),
.Y(n_524)
);

INVx1_ASAP7_75t_L g525 ( 
.A(n_450),
.Y(n_525)
);

NAND2xp5_ASAP7_75t_SL g526 ( 
.A(n_436),
.B(n_316),
.Y(n_526)
);

NAND2xp5_ASAP7_75t_L g527 ( 
.A(n_446),
.B(n_316),
.Y(n_527)
);

INVx1_ASAP7_75t_L g528 ( 
.A(n_409),
.Y(n_528)
);

INVx1_ASAP7_75t_SL g529 ( 
.A(n_417),
.Y(n_529)
);

INVx2_ASAP7_75t_L g530 ( 
.A(n_444),
.Y(n_530)
);

HB1xp67_ASAP7_75t_L g531 ( 
.A(n_400),
.Y(n_531)
);

NAND2xp5_ASAP7_75t_L g532 ( 
.A(n_444),
.B(n_276),
.Y(n_532)
);

AND2x4_ASAP7_75t_L g533 ( 
.A(n_441),
.B(n_59),
.Y(n_533)
);

INVx2_ASAP7_75t_L g534 ( 
.A(n_444),
.Y(n_534)
);

NOR2xp33_ASAP7_75t_L g535 ( 
.A(n_400),
.B(n_25),
.Y(n_535)
);

CKINVDCx20_ASAP7_75t_R g536 ( 
.A(n_417),
.Y(n_536)
);

NAND2xp5_ASAP7_75t_L g537 ( 
.A(n_444),
.B(n_276),
.Y(n_537)
);

INVx2_ASAP7_75t_SL g538 ( 
.A(n_400),
.Y(n_538)
);

INVxp67_ASAP7_75t_L g539 ( 
.A(n_427),
.Y(n_539)
);

NAND2xp5_ASAP7_75t_L g540 ( 
.A(n_444),
.B(n_284),
.Y(n_540)
);

HB1xp67_ASAP7_75t_L g541 ( 
.A(n_445),
.Y(n_541)
);

INVx1_ASAP7_75t_L g542 ( 
.A(n_448),
.Y(n_542)
);

AND2x2_ASAP7_75t_L g543 ( 
.A(n_448),
.B(n_326),
.Y(n_543)
);

AND2x2_ASAP7_75t_L g544 ( 
.A(n_515),
.B(n_426),
.Y(n_544)
);

INVx1_ASAP7_75t_L g545 ( 
.A(n_493),
.Y(n_545)
);

NAND2xp5_ASAP7_75t_L g546 ( 
.A(n_469),
.B(n_452),
.Y(n_546)
);

INVx2_ASAP7_75t_L g547 ( 
.A(n_470),
.Y(n_547)
);

NOR2xp33_ASAP7_75t_L g548 ( 
.A(n_520),
.B(n_456),
.Y(n_548)
);

NAND2xp5_ASAP7_75t_L g549 ( 
.A(n_469),
.B(n_472),
.Y(n_549)
);

INVx1_ASAP7_75t_L g550 ( 
.A(n_493),
.Y(n_550)
);

INVx1_ASAP7_75t_L g551 ( 
.A(n_474),
.Y(n_551)
);

INVx1_ASAP7_75t_L g552 ( 
.A(n_513),
.Y(n_552)
);

OR2x2_ASAP7_75t_L g553 ( 
.A(n_517),
.B(n_453),
.Y(n_553)
);

INVx2_ASAP7_75t_L g554 ( 
.A(n_470),
.Y(n_554)
);

AND2x2_ASAP7_75t_L g555 ( 
.A(n_515),
.B(n_437),
.Y(n_555)
);

BUFx2_ASAP7_75t_SL g556 ( 
.A(n_465),
.Y(n_556)
);

HB1xp67_ASAP7_75t_L g557 ( 
.A(n_510),
.Y(n_557)
);

INVx3_ASAP7_75t_L g558 ( 
.A(n_465),
.Y(n_558)
);

INVx5_ASAP7_75t_L g559 ( 
.A(n_461),
.Y(n_559)
);

OR2x2_ASAP7_75t_L g560 ( 
.A(n_521),
.B(n_399),
.Y(n_560)
);

NAND2x1_ASAP7_75t_L g561 ( 
.A(n_465),
.B(n_288),
.Y(n_561)
);

INVx3_ASAP7_75t_L g562 ( 
.A(n_509),
.Y(n_562)
);

INVx3_ASAP7_75t_L g563 ( 
.A(n_509),
.Y(n_563)
);

BUFx3_ASAP7_75t_L g564 ( 
.A(n_479),
.Y(n_564)
);

NAND2xp5_ASAP7_75t_L g565 ( 
.A(n_472),
.B(n_439),
.Y(n_565)
);

NAND2xp5_ASAP7_75t_SL g566 ( 
.A(n_479),
.B(n_416),
.Y(n_566)
);

INVx4_ASAP7_75t_L g567 ( 
.A(n_509),
.Y(n_567)
);

INVx1_ASAP7_75t_L g568 ( 
.A(n_513),
.Y(n_568)
);

BUFx3_ASAP7_75t_L g569 ( 
.A(n_533),
.Y(n_569)
);

NAND2xp5_ASAP7_75t_L g570 ( 
.A(n_516),
.B(n_326),
.Y(n_570)
);

BUFx3_ASAP7_75t_L g571 ( 
.A(n_533),
.Y(n_571)
);

AND2x4_ASAP7_75t_L g572 ( 
.A(n_533),
.B(n_486),
.Y(n_572)
);

NAND2xp5_ASAP7_75t_L g573 ( 
.A(n_516),
.B(n_326),
.Y(n_573)
);

INVx3_ASAP7_75t_L g574 ( 
.A(n_509),
.Y(n_574)
);

INVx2_ASAP7_75t_L g575 ( 
.A(n_473),
.Y(n_575)
);

INVx1_ASAP7_75t_L g576 ( 
.A(n_474),
.Y(n_576)
);

NAND2xp5_ASAP7_75t_L g577 ( 
.A(n_476),
.B(n_288),
.Y(n_577)
);

AND2x2_ASAP7_75t_L g578 ( 
.A(n_530),
.B(n_456),
.Y(n_578)
);

NAND2xp5_ASAP7_75t_L g579 ( 
.A(n_476),
.B(n_284),
.Y(n_579)
);

NAND2x1p5_ASAP7_75t_L g580 ( 
.A(n_530),
.B(n_284),
.Y(n_580)
);

OR2x6_ASAP7_75t_L g581 ( 
.A(n_534),
.B(n_429),
.Y(n_581)
);

NAND2xp5_ASAP7_75t_L g582 ( 
.A(n_524),
.B(n_525),
.Y(n_582)
);

INVx2_ASAP7_75t_L g583 ( 
.A(n_473),
.Y(n_583)
);

AND2x4_ASAP7_75t_L g584 ( 
.A(n_538),
.B(n_429),
.Y(n_584)
);

BUFx2_ASAP7_75t_L g585 ( 
.A(n_541),
.Y(n_585)
);

AND2x6_ASAP7_75t_L g586 ( 
.A(n_534),
.B(n_60),
.Y(n_586)
);

BUFx6f_ASAP7_75t_L g587 ( 
.A(n_468),
.Y(n_587)
);

BUFx2_ASAP7_75t_L g588 ( 
.A(n_528),
.Y(n_588)
);

AND2x4_ASAP7_75t_L g589 ( 
.A(n_538),
.B(n_508),
.Y(n_589)
);

BUFx2_ASAP7_75t_L g590 ( 
.A(n_528),
.Y(n_590)
);

NOR2xp33_ASAP7_75t_L g591 ( 
.A(n_471),
.B(n_442),
.Y(n_591)
);

AND2x4_ASAP7_75t_L g592 ( 
.A(n_508),
.B(n_61),
.Y(n_592)
);

INVx5_ASAP7_75t_L g593 ( 
.A(n_461),
.Y(n_593)
);

INVx2_ASAP7_75t_L g594 ( 
.A(n_480),
.Y(n_594)
);

AND2x4_ASAP7_75t_L g595 ( 
.A(n_492),
.B(n_497),
.Y(n_595)
);

OR2x6_ASAP7_75t_L g596 ( 
.A(n_492),
.B(n_62),
.Y(n_596)
);

AND2x4_ASAP7_75t_L g597 ( 
.A(n_497),
.B(n_63),
.Y(n_597)
);

INVx2_ASAP7_75t_L g598 ( 
.A(n_480),
.Y(n_598)
);

NAND2x1p5_ASAP7_75t_L g599 ( 
.A(n_468),
.B(n_284),
.Y(n_599)
);

INVx1_ASAP7_75t_L g600 ( 
.A(n_485),
.Y(n_600)
);

AND2x2_ASAP7_75t_L g601 ( 
.A(n_519),
.B(n_66),
.Y(n_601)
);

AND2x4_ASAP7_75t_L g602 ( 
.A(n_542),
.B(n_68),
.Y(n_602)
);

BUFx2_ASAP7_75t_L g603 ( 
.A(n_531),
.Y(n_603)
);

NAND2xp5_ASAP7_75t_L g604 ( 
.A(n_524),
.B(n_287),
.Y(n_604)
);

AND2x2_ASAP7_75t_L g605 ( 
.A(n_519),
.B(n_69),
.Y(n_605)
);

BUFx2_ASAP7_75t_L g606 ( 
.A(n_525),
.Y(n_606)
);

INVx5_ASAP7_75t_L g607 ( 
.A(n_461),
.Y(n_607)
);

INVx1_ASAP7_75t_L g608 ( 
.A(n_485),
.Y(n_608)
);

INVx1_ASAP7_75t_L g609 ( 
.A(n_506),
.Y(n_609)
);

INVx1_ASAP7_75t_L g610 ( 
.A(n_551),
.Y(n_610)
);

AND2x4_ASAP7_75t_L g611 ( 
.A(n_564),
.B(n_542),
.Y(n_611)
);

CKINVDCx20_ASAP7_75t_R g612 ( 
.A(n_585),
.Y(n_612)
);

INVxp67_ASAP7_75t_SL g613 ( 
.A(n_569),
.Y(n_613)
);

INVx2_ASAP7_75t_L g614 ( 
.A(n_594),
.Y(n_614)
);

NAND2xp5_ASAP7_75t_L g615 ( 
.A(n_549),
.B(n_460),
.Y(n_615)
);

INVx5_ASAP7_75t_SL g616 ( 
.A(n_596),
.Y(n_616)
);

BUFx3_ASAP7_75t_L g617 ( 
.A(n_603),
.Y(n_617)
);

BUFx2_ASAP7_75t_R g618 ( 
.A(n_565),
.Y(n_618)
);

INVx3_ASAP7_75t_L g619 ( 
.A(n_567),
.Y(n_619)
);

INVxp67_ASAP7_75t_SL g620 ( 
.A(n_569),
.Y(n_620)
);

INVx3_ASAP7_75t_L g621 ( 
.A(n_567),
.Y(n_621)
);

INVx1_ASAP7_75t_L g622 ( 
.A(n_551),
.Y(n_622)
);

BUFx5_ASAP7_75t_L g623 ( 
.A(n_586),
.Y(n_623)
);

NOR2xp33_ASAP7_75t_L g624 ( 
.A(n_548),
.B(n_518),
.Y(n_624)
);

INVx1_ASAP7_75t_L g625 ( 
.A(n_594),
.Y(n_625)
);

BUFx12f_ASAP7_75t_L g626 ( 
.A(n_553),
.Y(n_626)
);

OR2x2_ASAP7_75t_L g627 ( 
.A(n_578),
.B(n_529),
.Y(n_627)
);

AND2x2_ASAP7_75t_L g628 ( 
.A(n_578),
.B(n_460),
.Y(n_628)
);

BUFx2_ASAP7_75t_L g629 ( 
.A(n_581),
.Y(n_629)
);

BUFx6f_ASAP7_75t_L g630 ( 
.A(n_571),
.Y(n_630)
);

INVx6_ASAP7_75t_L g631 ( 
.A(n_572),
.Y(n_631)
);

NAND2xp5_ASAP7_75t_L g632 ( 
.A(n_595),
.B(n_523),
.Y(n_632)
);

INVx1_ASAP7_75t_SL g633 ( 
.A(n_553),
.Y(n_633)
);

BUFx3_ASAP7_75t_L g634 ( 
.A(n_603),
.Y(n_634)
);

NAND2x1p5_ASAP7_75t_L g635 ( 
.A(n_571),
.B(n_468),
.Y(n_635)
);

INVx1_ASAP7_75t_L g636 ( 
.A(n_598),
.Y(n_636)
);

BUFx3_ASAP7_75t_L g637 ( 
.A(n_585),
.Y(n_637)
);

INVx6_ASAP7_75t_SL g638 ( 
.A(n_596),
.Y(n_638)
);

INVx2_ASAP7_75t_SL g639 ( 
.A(n_572),
.Y(n_639)
);

BUFx5_ASAP7_75t_L g640 ( 
.A(n_586),
.Y(n_640)
);

INVx1_ASAP7_75t_L g641 ( 
.A(n_598),
.Y(n_641)
);

BUFx3_ASAP7_75t_L g642 ( 
.A(n_564),
.Y(n_642)
);

INVxp67_ASAP7_75t_SL g643 ( 
.A(n_558),
.Y(n_643)
);

BUFx12f_ASAP7_75t_L g644 ( 
.A(n_584),
.Y(n_644)
);

AND2x4_ASAP7_75t_L g645 ( 
.A(n_572),
.B(n_511),
.Y(n_645)
);

INVx3_ASAP7_75t_L g646 ( 
.A(n_567),
.Y(n_646)
);

INVx2_ASAP7_75t_L g647 ( 
.A(n_547),
.Y(n_647)
);

BUFx3_ASAP7_75t_L g648 ( 
.A(n_589),
.Y(n_648)
);

CKINVDCx14_ASAP7_75t_R g649 ( 
.A(n_560),
.Y(n_649)
);

INVx2_ASAP7_75t_SL g650 ( 
.A(n_557),
.Y(n_650)
);

NAND2x1p5_ASAP7_75t_L g651 ( 
.A(n_558),
.B(n_478),
.Y(n_651)
);

NAND2x1p5_ASAP7_75t_L g652 ( 
.A(n_558),
.B(n_478),
.Y(n_652)
);

BUFx10_ASAP7_75t_L g653 ( 
.A(n_591),
.Y(n_653)
);

AO21x1_ASAP7_75t_L g654 ( 
.A1(n_601),
.A2(n_491),
.B(n_494),
.Y(n_654)
);

BUFx3_ASAP7_75t_L g655 ( 
.A(n_589),
.Y(n_655)
);

BUFx3_ASAP7_75t_L g656 ( 
.A(n_589),
.Y(n_656)
);

BUFx4f_ASAP7_75t_SL g657 ( 
.A(n_566),
.Y(n_657)
);

BUFx5_ASAP7_75t_L g658 ( 
.A(n_586),
.Y(n_658)
);

INVx5_ASAP7_75t_L g659 ( 
.A(n_586),
.Y(n_659)
);

CKINVDCx20_ASAP7_75t_R g660 ( 
.A(n_560),
.Y(n_660)
);

AND2x2_ASAP7_75t_L g661 ( 
.A(n_555),
.B(n_482),
.Y(n_661)
);

NAND2x1p5_ASAP7_75t_L g662 ( 
.A(n_587),
.B(n_478),
.Y(n_662)
);

NAND2x1p5_ASAP7_75t_L g663 ( 
.A(n_587),
.B(n_484),
.Y(n_663)
);

OR2x2_ASAP7_75t_L g664 ( 
.A(n_581),
.B(n_477),
.Y(n_664)
);

INVx2_ASAP7_75t_L g665 ( 
.A(n_547),
.Y(n_665)
);

INVx2_ASAP7_75t_SL g666 ( 
.A(n_595),
.Y(n_666)
);

BUFx3_ASAP7_75t_L g667 ( 
.A(n_544),
.Y(n_667)
);

HB1xp67_ASAP7_75t_L g668 ( 
.A(n_633),
.Y(n_668)
);

INVx1_ASAP7_75t_L g669 ( 
.A(n_610),
.Y(n_669)
);

INVx1_ASAP7_75t_SL g670 ( 
.A(n_612),
.Y(n_670)
);

OAI22x1_ASAP7_75t_L g671 ( 
.A1(n_624),
.A2(n_588),
.B1(n_590),
.B2(n_606),
.Y(n_671)
);

BUFx6f_ASAP7_75t_L g672 ( 
.A(n_630),
.Y(n_672)
);

BUFx2_ASAP7_75t_L g673 ( 
.A(n_626),
.Y(n_673)
);

OAI22xp33_ASAP7_75t_L g674 ( 
.A1(n_615),
.A2(n_581),
.B1(n_590),
.B2(n_588),
.Y(n_674)
);

OAI22xp5_ASAP7_75t_L g675 ( 
.A1(n_624),
.A2(n_581),
.B1(n_587),
.B2(n_555),
.Y(n_675)
);

INVx1_ASAP7_75t_L g676 ( 
.A(n_622),
.Y(n_676)
);

AOI22xp33_ASAP7_75t_L g677 ( 
.A1(n_628),
.A2(n_596),
.B1(n_514),
.B2(n_606),
.Y(n_677)
);

OAI22xp33_ASAP7_75t_L g678 ( 
.A1(n_657),
.A2(n_587),
.B1(n_596),
.B2(n_568),
.Y(n_678)
);

INVx1_ASAP7_75t_SL g679 ( 
.A(n_612),
.Y(n_679)
);

INVx6_ASAP7_75t_L g680 ( 
.A(n_626),
.Y(n_680)
);

INVx1_ASAP7_75t_L g681 ( 
.A(n_625),
.Y(n_681)
);

BUFx5_ASAP7_75t_L g682 ( 
.A(n_636),
.Y(n_682)
);

INVx2_ASAP7_75t_L g683 ( 
.A(n_614),
.Y(n_683)
);

BUFx3_ASAP7_75t_L g684 ( 
.A(n_617),
.Y(n_684)
);

OAI21xp5_ASAP7_75t_L g685 ( 
.A1(n_632),
.A2(n_605),
.B(n_601),
.Y(n_685)
);

INVx1_ASAP7_75t_L g686 ( 
.A(n_641),
.Y(n_686)
);

INVx3_ASAP7_75t_SL g687 ( 
.A(n_627),
.Y(n_687)
);

AOI22xp33_ASAP7_75t_SL g688 ( 
.A1(n_616),
.A2(n_587),
.B1(n_535),
.B2(n_597),
.Y(n_688)
);

CKINVDCx8_ASAP7_75t_R g689 ( 
.A(n_629),
.Y(n_689)
);

INVx1_ASAP7_75t_L g690 ( 
.A(n_614),
.Y(n_690)
);

BUFx12f_ASAP7_75t_L g691 ( 
.A(n_644),
.Y(n_691)
);

INVx2_ASAP7_75t_L g692 ( 
.A(n_647),
.Y(n_692)
);

OAI22xp5_ASAP7_75t_L g693 ( 
.A1(n_635),
.A2(n_595),
.B1(n_552),
.B2(n_545),
.Y(n_693)
);

AND2x2_ASAP7_75t_L g694 ( 
.A(n_661),
.B(n_544),
.Y(n_694)
);

AOI22xp33_ASAP7_75t_L g695 ( 
.A1(n_657),
.A2(n_514),
.B1(n_550),
.B2(n_608),
.Y(n_695)
);

AOI22xp33_ASAP7_75t_L g696 ( 
.A1(n_667),
.A2(n_499),
.B1(n_597),
.B2(n_584),
.Y(n_696)
);

INVx1_ASAP7_75t_L g697 ( 
.A(n_647),
.Y(n_697)
);

AOI22xp33_ASAP7_75t_L g698 ( 
.A1(n_638),
.A2(n_600),
.B1(n_605),
.B2(n_597),
.Y(n_698)
);

AOI22xp33_ASAP7_75t_L g699 ( 
.A1(n_638),
.A2(n_586),
.B1(n_582),
.B2(n_490),
.Y(n_699)
);

CKINVDCx5p33_ASAP7_75t_R g700 ( 
.A(n_649),
.Y(n_700)
);

INVx1_ASAP7_75t_L g701 ( 
.A(n_665),
.Y(n_701)
);

INVx1_ASAP7_75t_L g702 ( 
.A(n_665),
.Y(n_702)
);

INVx1_ASAP7_75t_SL g703 ( 
.A(n_617),
.Y(n_703)
);

CKINVDCx11_ASAP7_75t_R g704 ( 
.A(n_660),
.Y(n_704)
);

NAND2xp5_ASAP7_75t_L g705 ( 
.A(n_667),
.B(n_511),
.Y(n_705)
);

INVx2_ASAP7_75t_L g706 ( 
.A(n_611),
.Y(n_706)
);

INVx1_ASAP7_75t_SL g707 ( 
.A(n_634),
.Y(n_707)
);

INVx5_ASAP7_75t_L g708 ( 
.A(n_619),
.Y(n_708)
);

BUFx3_ASAP7_75t_L g709 ( 
.A(n_634),
.Y(n_709)
);

BUFx3_ASAP7_75t_L g710 ( 
.A(n_637),
.Y(n_710)
);

OAI22xp33_ASAP7_75t_L g711 ( 
.A1(n_664),
.A2(n_638),
.B1(n_637),
.B2(n_659),
.Y(n_711)
);

INVx5_ASAP7_75t_L g712 ( 
.A(n_619),
.Y(n_712)
);

CKINVDCx11_ASAP7_75t_R g713 ( 
.A(n_660),
.Y(n_713)
);

INVx1_ASAP7_75t_L g714 ( 
.A(n_611),
.Y(n_714)
);

OAI22xp5_ASAP7_75t_L g715 ( 
.A1(n_635),
.A2(n_556),
.B1(n_599),
.B2(n_559),
.Y(n_715)
);

AOI22xp33_ASAP7_75t_L g716 ( 
.A1(n_616),
.A2(n_586),
.B1(n_475),
.B2(n_496),
.Y(n_716)
);

CKINVDCx20_ASAP7_75t_R g717 ( 
.A(n_649),
.Y(n_717)
);

BUFx3_ASAP7_75t_L g718 ( 
.A(n_650),
.Y(n_718)
);

INVx1_ASAP7_75t_L g719 ( 
.A(n_611),
.Y(n_719)
);

AOI22xp33_ASAP7_75t_SL g720 ( 
.A1(n_616),
.A2(n_512),
.B1(n_536),
.B2(n_592),
.Y(n_720)
);

CKINVDCx20_ASAP7_75t_R g721 ( 
.A(n_653),
.Y(n_721)
);

NAND2xp5_ASAP7_75t_L g722 ( 
.A(n_694),
.B(n_645),
.Y(n_722)
);

INVx1_ASAP7_75t_L g723 ( 
.A(n_669),
.Y(n_723)
);

AOI222xp33_ASAP7_75t_L g724 ( 
.A1(n_675),
.A2(n_539),
.B1(n_546),
.B2(n_644),
.C1(n_526),
.C2(n_584),
.Y(n_724)
);

AND2x2_ASAP7_75t_L g725 ( 
.A(n_687),
.B(n_481),
.Y(n_725)
);

INVx1_ASAP7_75t_L g726 ( 
.A(n_676),
.Y(n_726)
);

AOI22xp5_ASAP7_75t_L g727 ( 
.A1(n_717),
.A2(n_536),
.B1(n_482),
.B2(n_653),
.Y(n_727)
);

INVx1_ASAP7_75t_L g728 ( 
.A(n_681),
.Y(n_728)
);

OAI22xp5_ASAP7_75t_L g729 ( 
.A1(n_698),
.A2(n_618),
.B1(n_482),
.B2(n_642),
.Y(n_729)
);

OAI22xp5_ASAP7_75t_L g730 ( 
.A1(n_698),
.A2(n_642),
.B1(n_659),
.B2(n_620),
.Y(n_730)
);

AOI22xp33_ASAP7_75t_SL g731 ( 
.A1(n_680),
.A2(n_659),
.B1(n_640),
.B2(n_658),
.Y(n_731)
);

NOR2x1_ASAP7_75t_R g732 ( 
.A(n_691),
.B(n_704),
.Y(n_732)
);

AOI22xp33_ASAP7_75t_SL g733 ( 
.A1(n_680),
.A2(n_659),
.B1(n_640),
.B2(n_658),
.Y(n_733)
);

AOI22xp33_ASAP7_75t_L g734 ( 
.A1(n_687),
.A2(n_653),
.B1(n_645),
.B2(n_666),
.Y(n_734)
);

HB1xp67_ASAP7_75t_L g735 ( 
.A(n_668),
.Y(n_735)
);

AOI22xp33_ASAP7_75t_L g736 ( 
.A1(n_674),
.A2(n_645),
.B1(n_666),
.B2(n_602),
.Y(n_736)
);

AO22x1_ASAP7_75t_L g737 ( 
.A1(n_700),
.A2(n_592),
.B1(n_602),
.B2(n_613),
.Y(n_737)
);

INVx2_ASAP7_75t_L g738 ( 
.A(n_683),
.Y(n_738)
);

INVx1_ASAP7_75t_L g739 ( 
.A(n_686),
.Y(n_739)
);

OAI22xp33_ASAP7_75t_L g740 ( 
.A1(n_674),
.A2(n_501),
.B1(n_655),
.B2(n_648),
.Y(n_740)
);

AOI22xp33_ASAP7_75t_L g741 ( 
.A1(n_678),
.A2(n_602),
.B1(n_639),
.B2(n_656),
.Y(n_741)
);

OAI22xp5_ASAP7_75t_L g742 ( 
.A1(n_695),
.A2(n_720),
.B1(n_696),
.B2(n_677),
.Y(n_742)
);

NAND2xp5_ASAP7_75t_L g743 ( 
.A(n_705),
.B(n_650),
.Y(n_743)
);

BUFx12f_ASAP7_75t_SL g744 ( 
.A(n_672),
.Y(n_744)
);

AOI21xp33_ASAP7_75t_L g745 ( 
.A1(n_685),
.A2(n_654),
.B(n_577),
.Y(n_745)
);

OAI22xp33_ASAP7_75t_L g746 ( 
.A1(n_671),
.A2(n_648),
.B1(n_656),
.B2(n_655),
.Y(n_746)
);

AOI22xp5_ASAP7_75t_L g747 ( 
.A1(n_720),
.A2(n_512),
.B1(n_631),
.B2(n_639),
.Y(n_747)
);

INVx1_ASAP7_75t_L g748 ( 
.A(n_690),
.Y(n_748)
);

CKINVDCx5p33_ASAP7_75t_R g749 ( 
.A(n_713),
.Y(n_749)
);

INVx3_ASAP7_75t_L g750 ( 
.A(n_672),
.Y(n_750)
);

NAND2xp5_ASAP7_75t_L g751 ( 
.A(n_668),
.B(n_631),
.Y(n_751)
);

AOI22xp33_ASAP7_75t_SL g752 ( 
.A1(n_680),
.A2(n_623),
.B1(n_658),
.B2(n_640),
.Y(n_752)
);

OAI21xp5_ASAP7_75t_L g753 ( 
.A1(n_699),
.A2(n_579),
.B(n_502),
.Y(n_753)
);

BUFx6f_ASAP7_75t_L g754 ( 
.A(n_672),
.Y(n_754)
);

AOI22xp33_ASAP7_75t_L g755 ( 
.A1(n_678),
.A2(n_631),
.B1(n_592),
.B2(n_503),
.Y(n_755)
);

INVx1_ASAP7_75t_L g756 ( 
.A(n_697),
.Y(n_756)
);

INVx2_ASAP7_75t_L g757 ( 
.A(n_692),
.Y(n_757)
);

NAND2xp5_ASAP7_75t_L g758 ( 
.A(n_706),
.B(n_630),
.Y(n_758)
);

AOI22xp33_ASAP7_75t_SL g759 ( 
.A1(n_721),
.A2(n_623),
.B1(n_640),
.B2(n_658),
.Y(n_759)
);

INVx3_ASAP7_75t_L g760 ( 
.A(n_672),
.Y(n_760)
);

OR2x2_ASAP7_75t_SL g761 ( 
.A(n_714),
.B(n_466),
.Y(n_761)
);

INVx1_ASAP7_75t_L g762 ( 
.A(n_701),
.Y(n_762)
);

AOI22xp33_ASAP7_75t_L g763 ( 
.A1(n_688),
.A2(n_495),
.B1(n_503),
.B2(n_488),
.Y(n_763)
);

INVx2_ASAP7_75t_L g764 ( 
.A(n_702),
.Y(n_764)
);

INVx1_ASAP7_75t_L g765 ( 
.A(n_719),
.Y(n_765)
);

OAI22xp5_ASAP7_75t_L g766 ( 
.A1(n_695),
.A2(n_677),
.B1(n_688),
.B2(n_699),
.Y(n_766)
);

INVx1_ASAP7_75t_L g767 ( 
.A(n_682),
.Y(n_767)
);

AOI22xp33_ASAP7_75t_L g768 ( 
.A1(n_670),
.A2(n_679),
.B1(n_673),
.B2(n_693),
.Y(n_768)
);

AOI22xp33_ASAP7_75t_L g769 ( 
.A1(n_718),
.A2(n_505),
.B1(n_489),
.B2(n_488),
.Y(n_769)
);

INVx2_ASAP7_75t_L g770 ( 
.A(n_682),
.Y(n_770)
);

AND2x2_ASAP7_75t_L g771 ( 
.A(n_703),
.B(n_543),
.Y(n_771)
);

OAI22xp33_ASAP7_75t_L g772 ( 
.A1(n_689),
.A2(n_576),
.B1(n_609),
.B2(n_630),
.Y(n_772)
);

NAND2xp5_ASAP7_75t_L g773 ( 
.A(n_707),
.B(n_630),
.Y(n_773)
);

AOI22xp33_ASAP7_75t_L g774 ( 
.A1(n_711),
.A2(n_505),
.B1(n_489),
.B2(n_495),
.Y(n_774)
);

NAND2xp5_ASAP7_75t_L g775 ( 
.A(n_684),
.B(n_543),
.Y(n_775)
);

OAI22xp5_ASAP7_75t_L g776 ( 
.A1(n_716),
.A2(n_556),
.B1(n_662),
.B2(n_663),
.Y(n_776)
);

CKINVDCx5p33_ASAP7_75t_R g777 ( 
.A(n_709),
.Y(n_777)
);

HB1xp67_ASAP7_75t_L g778 ( 
.A(n_708),
.Y(n_778)
);

AOI22xp33_ASAP7_75t_SL g779 ( 
.A1(n_710),
.A2(n_658),
.B1(n_623),
.B2(n_640),
.Y(n_779)
);

INVx2_ASAP7_75t_SL g780 ( 
.A(n_708),
.Y(n_780)
);

BUFx6f_ASAP7_75t_L g781 ( 
.A(n_708),
.Y(n_781)
);

INVx1_ASAP7_75t_L g782 ( 
.A(n_682),
.Y(n_782)
);

AOI222xp33_ASAP7_75t_L g783 ( 
.A1(n_742),
.A2(n_716),
.B1(n_711),
.B2(n_487),
.C1(n_462),
.C2(n_464),
.Y(n_783)
);

OAI21xp5_ASAP7_75t_SL g784 ( 
.A1(n_724),
.A2(n_663),
.B(n_662),
.Y(n_784)
);

OAI22xp33_ASAP7_75t_L g785 ( 
.A1(n_766),
.A2(n_712),
.B1(n_708),
.B2(n_609),
.Y(n_785)
);

AOI22xp5_ASAP7_75t_L g786 ( 
.A1(n_729),
.A2(n_640),
.B1(n_623),
.B2(n_658),
.Y(n_786)
);

AOI221xp5_ASAP7_75t_L g787 ( 
.A1(n_745),
.A2(n_487),
.B1(n_483),
.B2(n_573),
.C(n_570),
.Y(n_787)
);

OAI22xp5_ASAP7_75t_L g788 ( 
.A1(n_768),
.A2(n_599),
.B1(n_712),
.B2(n_643),
.Y(n_788)
);

AOI22xp5_ASAP7_75t_L g789 ( 
.A1(n_747),
.A2(n_727),
.B1(n_734),
.B2(n_725),
.Y(n_789)
);

OAI21xp5_ASAP7_75t_SL g790 ( 
.A1(n_759),
.A2(n_484),
.B(n_715),
.Y(n_790)
);

AOI22xp5_ASAP7_75t_L g791 ( 
.A1(n_749),
.A2(n_623),
.B1(n_483),
.B2(n_461),
.Y(n_791)
);

AOI22xp33_ASAP7_75t_L g792 ( 
.A1(n_736),
.A2(n_506),
.B1(n_623),
.B2(n_500),
.Y(n_792)
);

OAI21xp5_ASAP7_75t_L g793 ( 
.A1(n_753),
.A2(n_527),
.B(n_504),
.Y(n_793)
);

AOI22xp33_ASAP7_75t_L g794 ( 
.A1(n_722),
.A2(n_746),
.B1(n_771),
.B2(n_741),
.Y(n_794)
);

AND2x6_ASAP7_75t_L g795 ( 
.A(n_781),
.B(n_619),
.Y(n_795)
);

AOI22xp33_ASAP7_75t_L g796 ( 
.A1(n_755),
.A2(n_506),
.B1(n_507),
.B2(n_500),
.Y(n_796)
);

AOI21xp5_ASAP7_75t_SL g797 ( 
.A1(n_781),
.A2(n_599),
.B(n_652),
.Y(n_797)
);

AOI22xp33_ASAP7_75t_SL g798 ( 
.A1(n_730),
.A2(n_776),
.B1(n_781),
.B2(n_735),
.Y(n_798)
);

AOI22xp33_ASAP7_75t_SL g799 ( 
.A1(n_781),
.A2(n_735),
.B1(n_751),
.B2(n_743),
.Y(n_799)
);

AOI22xp33_ASAP7_75t_L g800 ( 
.A1(n_740),
.A2(n_507),
.B1(n_682),
.B2(n_461),
.Y(n_800)
);

INVx1_ASAP7_75t_L g801 ( 
.A(n_723),
.Y(n_801)
);

OAI22xp5_ASAP7_75t_L g802 ( 
.A1(n_761),
.A2(n_712),
.B1(n_652),
.B2(n_651),
.Y(n_802)
);

AOI22xp33_ASAP7_75t_L g803 ( 
.A1(n_740),
.A2(n_682),
.B1(n_461),
.B2(n_509),
.Y(n_803)
);

AOI22xp33_ASAP7_75t_L g804 ( 
.A1(n_759),
.A2(n_682),
.B1(n_461),
.B2(n_522),
.Y(n_804)
);

NOR3xp33_ASAP7_75t_L g805 ( 
.A(n_737),
.B(n_498),
.C(n_604),
.Y(n_805)
);

AOI22xp33_ASAP7_75t_L g806 ( 
.A1(n_763),
.A2(n_775),
.B1(n_774),
.B2(n_772),
.Y(n_806)
);

AOI22xp33_ASAP7_75t_L g807 ( 
.A1(n_726),
.A2(n_575),
.B1(n_554),
.B2(n_583),
.Y(n_807)
);

AOI22xp33_ASAP7_75t_L g808 ( 
.A1(n_772),
.A2(n_522),
.B1(n_562),
.B2(n_563),
.Y(n_808)
);

AOI22xp33_ASAP7_75t_SL g809 ( 
.A1(n_778),
.A2(n_712),
.B1(n_621),
.B2(n_646),
.Y(n_809)
);

AND2x2_ASAP7_75t_L g810 ( 
.A(n_758),
.B(n_562),
.Y(n_810)
);

INVx2_ASAP7_75t_L g811 ( 
.A(n_738),
.Y(n_811)
);

OAI22xp5_ASAP7_75t_L g812 ( 
.A1(n_769),
.A2(n_773),
.B1(n_777),
.B2(n_779),
.Y(n_812)
);

OAI22xp5_ASAP7_75t_L g813 ( 
.A1(n_779),
.A2(n_651),
.B1(n_646),
.B2(n_621),
.Y(n_813)
);

OAI221xp5_ASAP7_75t_L g814 ( 
.A1(n_731),
.A2(n_532),
.B1(n_537),
.B2(n_540),
.C(n_467),
.Y(n_814)
);

INVxp67_ASAP7_75t_SL g815 ( 
.A(n_778),
.Y(n_815)
);

OAI22xp5_ASAP7_75t_L g816 ( 
.A1(n_731),
.A2(n_733),
.B1(n_752),
.B2(n_739),
.Y(n_816)
);

AOI21xp33_ASAP7_75t_L g817 ( 
.A1(n_765),
.A2(n_554),
.B(n_575),
.Y(n_817)
);

NAND2xp5_ASAP7_75t_L g818 ( 
.A(n_757),
.B(n_583),
.Y(n_818)
);

AOI22xp33_ASAP7_75t_L g819 ( 
.A1(n_752),
.A2(n_522),
.B1(n_562),
.B2(n_563),
.Y(n_819)
);

OAI22xp5_ASAP7_75t_L g820 ( 
.A1(n_733),
.A2(n_621),
.B1(n_574),
.B2(n_563),
.Y(n_820)
);

AOI22xp33_ASAP7_75t_L g821 ( 
.A1(n_728),
.A2(n_522),
.B1(n_574),
.B2(n_484),
.Y(n_821)
);

INVx1_ASAP7_75t_SL g822 ( 
.A(n_750),
.Y(n_822)
);

INVxp67_ASAP7_75t_SL g823 ( 
.A(n_764),
.Y(n_823)
);

NAND3xp33_ASAP7_75t_L g824 ( 
.A(n_748),
.B(n_762),
.C(n_756),
.Y(n_824)
);

NOR2xp33_ASAP7_75t_L g825 ( 
.A(n_732),
.B(n_750),
.Y(n_825)
);

INVx1_ASAP7_75t_L g826 ( 
.A(n_767),
.Y(n_826)
);

AOI22xp33_ASAP7_75t_L g827 ( 
.A1(n_782),
.A2(n_522),
.B1(n_574),
.B2(n_463),
.Y(n_827)
);

AOI22xp33_ASAP7_75t_L g828 ( 
.A1(n_770),
.A2(n_522),
.B1(n_561),
.B2(n_580),
.Y(n_828)
);

AOI22xp33_ASAP7_75t_L g829 ( 
.A1(n_760),
.A2(n_522),
.B1(n_561),
.B2(n_580),
.Y(n_829)
);

AOI22xp33_ASAP7_75t_L g830 ( 
.A1(n_744),
.A2(n_26),
.B1(n_27),
.B2(n_28),
.Y(n_830)
);

AOI22xp33_ASAP7_75t_L g831 ( 
.A1(n_760),
.A2(n_780),
.B1(n_754),
.B2(n_30),
.Y(n_831)
);

NAND2xp5_ASAP7_75t_L g832 ( 
.A(n_823),
.B(n_754),
.Y(n_832)
);

INVx1_ASAP7_75t_L g833 ( 
.A(n_826),
.Y(n_833)
);

NAND2xp5_ASAP7_75t_L g834 ( 
.A(n_801),
.B(n_754),
.Y(n_834)
);

NAND3xp33_ASAP7_75t_L g835 ( 
.A(n_830),
.B(n_754),
.C(n_29),
.Y(n_835)
);

AOI221xp5_ASAP7_75t_L g836 ( 
.A1(n_830),
.A2(n_26),
.B1(n_29),
.B2(n_30),
.C(n_31),
.Y(n_836)
);

AND2x2_ASAP7_75t_L g837 ( 
.A(n_816),
.B(n_31),
.Y(n_837)
);

AOI211xp5_ASAP7_75t_L g838 ( 
.A1(n_785),
.A2(n_32),
.B(n_33),
.C(n_35),
.Y(n_838)
);

AND2x2_ASAP7_75t_L g839 ( 
.A(n_815),
.B(n_32),
.Y(n_839)
);

NAND2xp5_ASAP7_75t_L g840 ( 
.A(n_811),
.B(n_36),
.Y(n_840)
);

NAND2xp5_ASAP7_75t_L g841 ( 
.A(n_799),
.B(n_36),
.Y(n_841)
);

NAND2xp5_ASAP7_75t_L g842 ( 
.A(n_824),
.B(n_37),
.Y(n_842)
);

OAI22xp5_ASAP7_75t_L g843 ( 
.A1(n_789),
.A2(n_607),
.B1(n_593),
.B2(n_559),
.Y(n_843)
);

AND2x2_ASAP7_75t_L g844 ( 
.A(n_810),
.B(n_798),
.Y(n_844)
);

AND2x2_ASAP7_75t_L g845 ( 
.A(n_803),
.B(n_37),
.Y(n_845)
);

AOI22xp33_ASAP7_75t_L g846 ( 
.A1(n_794),
.A2(n_607),
.B1(n_593),
.B2(n_559),
.Y(n_846)
);

AND2x2_ASAP7_75t_L g847 ( 
.A(n_822),
.B(n_38),
.Y(n_847)
);

NAND3xp33_ASAP7_75t_L g848 ( 
.A(n_831),
.B(n_38),
.C(n_39),
.Y(n_848)
);

OAI22xp5_ASAP7_75t_L g849 ( 
.A1(n_806),
.A2(n_607),
.B1(n_593),
.B2(n_559),
.Y(n_849)
);

NAND2xp5_ASAP7_75t_L g850 ( 
.A(n_785),
.B(n_70),
.Y(n_850)
);

NAND4xp25_ASAP7_75t_L g851 ( 
.A(n_831),
.B(n_72),
.C(n_74),
.D(n_75),
.Y(n_851)
);

NAND2xp5_ASAP7_75t_L g852 ( 
.A(n_812),
.B(n_79),
.Y(n_852)
);

OAI221xp5_ASAP7_75t_L g853 ( 
.A1(n_784),
.A2(n_580),
.B1(n_607),
.B2(n_593),
.C(n_559),
.Y(n_853)
);

NAND2xp5_ASAP7_75t_L g854 ( 
.A(n_818),
.B(n_783),
.Y(n_854)
);

OAI22xp5_ASAP7_75t_L g855 ( 
.A1(n_800),
.A2(n_607),
.B1(n_593),
.B2(n_287),
.Y(n_855)
);

AND2x2_ASAP7_75t_L g856 ( 
.A(n_786),
.B(n_80),
.Y(n_856)
);

AOI21xp5_ASAP7_75t_SL g857 ( 
.A1(n_788),
.A2(n_81),
.B(n_82),
.Y(n_857)
);

NAND4xp25_ASAP7_75t_L g858 ( 
.A(n_825),
.B(n_83),
.C(n_84),
.D(n_87),
.Y(n_858)
);

OAI211xp5_ASAP7_75t_L g859 ( 
.A1(n_790),
.A2(n_287),
.B(n_89),
.C(n_92),
.Y(n_859)
);

NAND2xp5_ASAP7_75t_L g860 ( 
.A(n_802),
.B(n_88),
.Y(n_860)
);

AND2x2_ASAP7_75t_L g861 ( 
.A(n_804),
.B(n_94),
.Y(n_861)
);

NAND2xp5_ASAP7_75t_L g862 ( 
.A(n_792),
.B(n_95),
.Y(n_862)
);

AOI22xp33_ASAP7_75t_L g863 ( 
.A1(n_805),
.A2(n_287),
.B1(n_97),
.B2(n_98),
.Y(n_863)
);

NAND2xp5_ASAP7_75t_L g864 ( 
.A(n_787),
.B(n_96),
.Y(n_864)
);

AND2x2_ASAP7_75t_L g865 ( 
.A(n_819),
.B(n_101),
.Y(n_865)
);

NAND2xp5_ASAP7_75t_L g866 ( 
.A(n_807),
.B(n_102),
.Y(n_866)
);

AND2x2_ASAP7_75t_L g867 ( 
.A(n_791),
.B(n_793),
.Y(n_867)
);

OAI21xp5_ASAP7_75t_SL g868 ( 
.A1(n_808),
.A2(n_103),
.B(n_104),
.Y(n_868)
);

NAND3xp33_ASAP7_75t_L g869 ( 
.A(n_838),
.B(n_809),
.C(n_821),
.Y(n_869)
);

OR2x2_ASAP7_75t_L g870 ( 
.A(n_833),
.B(n_832),
.Y(n_870)
);

AND2x2_ASAP7_75t_L g871 ( 
.A(n_844),
.B(n_833),
.Y(n_871)
);

OR2x2_ASAP7_75t_L g872 ( 
.A(n_834),
.B(n_817),
.Y(n_872)
);

NAND3xp33_ASAP7_75t_L g873 ( 
.A(n_838),
.B(n_827),
.C(n_796),
.Y(n_873)
);

AND2x2_ASAP7_75t_L g874 ( 
.A(n_844),
.B(n_813),
.Y(n_874)
);

NOR3xp33_ASAP7_75t_L g875 ( 
.A(n_835),
.B(n_814),
.C(n_820),
.Y(n_875)
);

OAI221xp5_ASAP7_75t_L g876 ( 
.A1(n_835),
.A2(n_829),
.B1(n_807),
.B2(n_828),
.C(n_797),
.Y(n_876)
);

AO21x2_ASAP7_75t_L g877 ( 
.A1(n_842),
.A2(n_857),
.B(n_852),
.Y(n_877)
);

NAND3xp33_ASAP7_75t_L g878 ( 
.A(n_836),
.B(n_795),
.C(n_108),
.Y(n_878)
);

OR2x2_ASAP7_75t_L g879 ( 
.A(n_867),
.B(n_854),
.Y(n_879)
);

NOR3xp33_ASAP7_75t_L g880 ( 
.A(n_848),
.B(n_795),
.C(n_109),
.Y(n_880)
);

AND2x2_ASAP7_75t_L g881 ( 
.A(n_839),
.B(n_795),
.Y(n_881)
);

BUFx2_ASAP7_75t_L g882 ( 
.A(n_839),
.Y(n_882)
);

NAND3xp33_ASAP7_75t_L g883 ( 
.A(n_848),
.B(n_795),
.C(n_111),
.Y(n_883)
);

NOR2xp33_ASAP7_75t_L g884 ( 
.A(n_837),
.B(n_795),
.Y(n_884)
);

NAND3xp33_ASAP7_75t_SL g885 ( 
.A(n_837),
.B(n_107),
.C(n_112),
.Y(n_885)
);

AOI22xp5_ASAP7_75t_L g886 ( 
.A1(n_851),
.A2(n_114),
.B1(n_115),
.B2(n_116),
.Y(n_886)
);

INVx1_ASAP7_75t_L g887 ( 
.A(n_840),
.Y(n_887)
);

INVx2_ASAP7_75t_L g888 ( 
.A(n_867),
.Y(n_888)
);

AND2x2_ASAP7_75t_L g889 ( 
.A(n_847),
.B(n_118),
.Y(n_889)
);

AND2x2_ASAP7_75t_L g890 ( 
.A(n_847),
.B(n_122),
.Y(n_890)
);

NAND4xp75_ASAP7_75t_L g891 ( 
.A(n_841),
.B(n_124),
.C(n_127),
.D(n_130),
.Y(n_891)
);

NAND3xp33_ASAP7_75t_L g892 ( 
.A(n_863),
.B(n_131),
.C(n_132),
.Y(n_892)
);

NOR3xp33_ASAP7_75t_L g893 ( 
.A(n_859),
.B(n_134),
.C(n_135),
.Y(n_893)
);

NAND3xp33_ASAP7_75t_L g894 ( 
.A(n_864),
.B(n_136),
.C(n_137),
.Y(n_894)
);

INVx1_ASAP7_75t_L g895 ( 
.A(n_870),
.Y(n_895)
);

NAND4xp75_ASAP7_75t_L g896 ( 
.A(n_886),
.B(n_845),
.C(n_850),
.D(n_856),
.Y(n_896)
);

INVxp67_ASAP7_75t_L g897 ( 
.A(n_871),
.Y(n_897)
);

XNOR2x2_ASAP7_75t_L g898 ( 
.A(n_883),
.B(n_858),
.Y(n_898)
);

NOR4xp25_ASAP7_75t_L g899 ( 
.A(n_879),
.B(n_853),
.C(n_845),
.D(n_868),
.Y(n_899)
);

NOR4xp25_ASAP7_75t_L g900 ( 
.A(n_878),
.B(n_856),
.C(n_860),
.D(n_865),
.Y(n_900)
);

AND2x2_ASAP7_75t_L g901 ( 
.A(n_888),
.B(n_857),
.Y(n_901)
);

AND2x2_ASAP7_75t_L g902 ( 
.A(n_888),
.B(n_861),
.Y(n_902)
);

NAND3xp33_ASAP7_75t_SL g903 ( 
.A(n_880),
.B(n_846),
.C(n_862),
.Y(n_903)
);

XOR2x2_ASAP7_75t_L g904 ( 
.A(n_882),
.B(n_865),
.Y(n_904)
);

INVx1_ASAP7_75t_L g905 ( 
.A(n_887),
.Y(n_905)
);

NOR3xp33_ASAP7_75t_L g906 ( 
.A(n_880),
.B(n_866),
.C(n_843),
.Y(n_906)
);

INVx2_ASAP7_75t_L g907 ( 
.A(n_872),
.Y(n_907)
);

NAND2xp5_ASAP7_75t_L g908 ( 
.A(n_874),
.B(n_849),
.Y(n_908)
);

XNOR2xp5_ASAP7_75t_L g909 ( 
.A(n_889),
.B(n_861),
.Y(n_909)
);

NAND2xp5_ASAP7_75t_SL g910 ( 
.A(n_874),
.B(n_855),
.Y(n_910)
);

INVx1_ASAP7_75t_L g911 ( 
.A(n_905),
.Y(n_911)
);

INVx1_ASAP7_75t_L g912 ( 
.A(n_905),
.Y(n_912)
);

INVx2_ASAP7_75t_SL g913 ( 
.A(n_895),
.Y(n_913)
);

XOR2x2_ASAP7_75t_L g914 ( 
.A(n_904),
.B(n_891),
.Y(n_914)
);

XOR2xp5_ASAP7_75t_L g915 ( 
.A(n_909),
.B(n_890),
.Y(n_915)
);

AND2x2_ASAP7_75t_L g916 ( 
.A(n_907),
.B(n_881),
.Y(n_916)
);

INVx3_ASAP7_75t_L g917 ( 
.A(n_907),
.Y(n_917)
);

XOR2x2_ASAP7_75t_L g918 ( 
.A(n_904),
.B(n_869),
.Y(n_918)
);

INVx1_ASAP7_75t_L g919 ( 
.A(n_897),
.Y(n_919)
);

AOI22xp5_ASAP7_75t_L g920 ( 
.A1(n_918),
.A2(n_896),
.B1(n_877),
.B2(n_906),
.Y(n_920)
);

AOI22xp5_ASAP7_75t_L g921 ( 
.A1(n_918),
.A2(n_896),
.B1(n_877),
.B2(n_875),
.Y(n_921)
);

INVx1_ASAP7_75t_L g922 ( 
.A(n_911),
.Y(n_922)
);

OA22x2_ASAP7_75t_L g923 ( 
.A1(n_915),
.A2(n_909),
.B1(n_919),
.B2(n_913),
.Y(n_923)
);

OAI22xp33_ASAP7_75t_L g924 ( 
.A1(n_914),
.A2(n_908),
.B1(n_903),
.B2(n_873),
.Y(n_924)
);

AOI22xp5_ASAP7_75t_L g925 ( 
.A1(n_914),
.A2(n_875),
.B1(n_899),
.B2(n_893),
.Y(n_925)
);

INVx1_ASAP7_75t_L g926 ( 
.A(n_912),
.Y(n_926)
);

AOI22xp5_ASAP7_75t_SL g927 ( 
.A1(n_917),
.A2(n_901),
.B1(n_889),
.B2(n_884),
.Y(n_927)
);

OA22x2_ASAP7_75t_L g928 ( 
.A1(n_913),
.A2(n_901),
.B1(n_902),
.B2(n_910),
.Y(n_928)
);

INVx1_ASAP7_75t_L g929 ( 
.A(n_922),
.Y(n_929)
);

INVxp67_ASAP7_75t_SL g930 ( 
.A(n_925),
.Y(n_930)
);

INVxp67_ASAP7_75t_L g931 ( 
.A(n_923),
.Y(n_931)
);

INVx1_ASAP7_75t_L g932 ( 
.A(n_926),
.Y(n_932)
);

INVx2_ASAP7_75t_L g933 ( 
.A(n_928),
.Y(n_933)
);

INVx1_ASAP7_75t_L g934 ( 
.A(n_921),
.Y(n_934)
);

INVx1_ASAP7_75t_L g935 ( 
.A(n_929),
.Y(n_935)
);

INVx1_ASAP7_75t_L g936 ( 
.A(n_929),
.Y(n_936)
);

BUFx4_ASAP7_75t_R g937 ( 
.A(n_933),
.Y(n_937)
);

INVx1_ASAP7_75t_L g938 ( 
.A(n_935),
.Y(n_938)
);

INVx1_ASAP7_75t_L g939 ( 
.A(n_936),
.Y(n_939)
);

INVx1_ASAP7_75t_L g940 ( 
.A(n_937),
.Y(n_940)
);

INVx1_ASAP7_75t_L g941 ( 
.A(n_935),
.Y(n_941)
);

INVx1_ASAP7_75t_L g942 ( 
.A(n_938),
.Y(n_942)
);

INVx1_ASAP7_75t_L g943 ( 
.A(n_939),
.Y(n_943)
);

NOR2xp33_ASAP7_75t_L g944 ( 
.A(n_940),
.B(n_930),
.Y(n_944)
);

NOR2xp33_ASAP7_75t_L g945 ( 
.A(n_941),
.B(n_931),
.Y(n_945)
);

NOR2xp33_ASAP7_75t_L g946 ( 
.A(n_940),
.B(n_934),
.Y(n_946)
);

NOR2x1_ASAP7_75t_L g947 ( 
.A(n_940),
.B(n_924),
.Y(n_947)
);

AOI22xp5_ASAP7_75t_L g948 ( 
.A1(n_947),
.A2(n_920),
.B1(n_933),
.B2(n_932),
.Y(n_948)
);

INVx2_ASAP7_75t_L g949 ( 
.A(n_942),
.Y(n_949)
);

NOR2x1_ASAP7_75t_L g950 ( 
.A(n_944),
.B(n_917),
.Y(n_950)
);

INVx1_ASAP7_75t_L g951 ( 
.A(n_946),
.Y(n_951)
);

AOI22xp5_ASAP7_75t_L g952 ( 
.A1(n_945),
.A2(n_943),
.B1(n_900),
.B2(n_917),
.Y(n_952)
);

INVx2_ASAP7_75t_L g953 ( 
.A(n_942),
.Y(n_953)
);

OAI22xp5_ASAP7_75t_L g954 ( 
.A1(n_948),
.A2(n_927),
.B1(n_916),
.B2(n_884),
.Y(n_954)
);

NAND4xp75_ASAP7_75t_L g955 ( 
.A(n_950),
.B(n_951),
.C(n_953),
.D(n_949),
.Y(n_955)
);

NOR2xp67_ASAP7_75t_L g956 ( 
.A(n_952),
.B(n_916),
.Y(n_956)
);

INVx1_ASAP7_75t_L g957 ( 
.A(n_951),
.Y(n_957)
);

INVx2_ASAP7_75t_L g958 ( 
.A(n_950),
.Y(n_958)
);

INVx1_ASAP7_75t_L g959 ( 
.A(n_957),
.Y(n_959)
);

INVx2_ASAP7_75t_L g960 ( 
.A(n_958),
.Y(n_960)
);

INVx1_ASAP7_75t_L g961 ( 
.A(n_955),
.Y(n_961)
);

INVx2_ASAP7_75t_L g962 ( 
.A(n_954),
.Y(n_962)
);

OAI22xp5_ASAP7_75t_SL g963 ( 
.A1(n_956),
.A2(n_892),
.B1(n_894),
.B2(n_898),
.Y(n_963)
);

AOI221xp5_ASAP7_75t_SL g964 ( 
.A1(n_961),
.A2(n_898),
.B1(n_876),
.B2(n_902),
.C(n_893),
.Y(n_964)
);

AOI22xp33_ASAP7_75t_SL g965 ( 
.A1(n_963),
.A2(n_885),
.B1(n_139),
.B2(n_140),
.Y(n_965)
);

OAI22xp33_ASAP7_75t_L g966 ( 
.A1(n_962),
.A2(n_138),
.B1(n_141),
.B2(n_143),
.Y(n_966)
);

NAND4xp75_ASAP7_75t_L g967 ( 
.A(n_960),
.B(n_145),
.C(n_146),
.D(n_149),
.Y(n_967)
);

AOI22xp5_ASAP7_75t_L g968 ( 
.A1(n_963),
.A2(n_151),
.B1(n_152),
.B2(n_153),
.Y(n_968)
);

OAI22xp5_ASAP7_75t_SL g969 ( 
.A1(n_959),
.A2(n_156),
.B1(n_157),
.B2(n_158),
.Y(n_969)
);

INVx2_ASAP7_75t_L g970 ( 
.A(n_967),
.Y(n_970)
);

INVx1_ASAP7_75t_L g971 ( 
.A(n_968),
.Y(n_971)
);

INVx1_ASAP7_75t_L g972 ( 
.A(n_969),
.Y(n_972)
);

OAI22xp33_ASAP7_75t_L g973 ( 
.A1(n_972),
.A2(n_966),
.B1(n_964),
.B2(n_965),
.Y(n_973)
);

OAI22xp5_ASAP7_75t_L g974 ( 
.A1(n_970),
.A2(n_159),
.B1(n_161),
.B2(n_164),
.Y(n_974)
);

INVx1_ASAP7_75t_L g975 ( 
.A(n_973),
.Y(n_975)
);

INVx1_ASAP7_75t_L g976 ( 
.A(n_974),
.Y(n_976)
);

AOI22xp5_ASAP7_75t_L g977 ( 
.A1(n_975),
.A2(n_971),
.B1(n_168),
.B2(n_172),
.Y(n_977)
);

AOI22xp5_ASAP7_75t_SL g978 ( 
.A1(n_976),
.A2(n_165),
.B1(n_174),
.B2(n_179),
.Y(n_978)
);

INVx1_ASAP7_75t_L g979 ( 
.A(n_977),
.Y(n_979)
);

AOI221x1_ASAP7_75t_L g980 ( 
.A1(n_979),
.A2(n_978),
.B1(n_181),
.B2(n_182),
.C(n_183),
.Y(n_980)
);

AOI211xp5_ASAP7_75t_L g981 ( 
.A1(n_980),
.A2(n_180),
.B(n_184),
.C(n_187),
.Y(n_981)
);


endmodule