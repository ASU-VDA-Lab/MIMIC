module real_aes_515_n_104 (n_17, n_28, n_76, n_56, n_34, n_98, n_90, n_82, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_83, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_91, n_100, n_43, n_103, n_96, n_54, n_35, n_42, n_99, n_15, n_9, n_23, n_72, n_95, n_44, n_102, n_7, n_4, n_80, n_6, n_12, n_68, n_79, n_69, n_46, n_59, n_25, n_73, n_77, n_81, n_48, n_37, n_97, n_70, n_50, n_89, n_26, n_86, n_93, n_13, n_24, n_2, n_55, n_62, n_84, n_67, n_92, n_33, n_88, n_14, n_11, n_85, n_16, n_94, n_39, n_5, n_45, n_60, n_38, n_87, n_0, n_78, n_101, n_63, n_1, n_53, n_36, n_104);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_98;
input n_90;
input n_82;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_83;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_91;
input n_100;
input n_43;
input n_103;
input n_96;
input n_54;
input n_35;
input n_42;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_95;
input n_44;
input n_102;
input n_7;
input n_4;
input n_80;
input n_6;
input n_12;
input n_68;
input n_79;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_81;
input n_48;
input n_37;
input n_97;
input n_70;
input n_50;
input n_89;
input n_26;
input n_86;
input n_93;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_84;
input n_67;
input n_92;
input n_33;
input n_88;
input n_14;
input n_11;
input n_85;
input n_16;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_87;
input n_0;
input n_78;
input n_101;
input n_63;
input n_1;
input n_53;
input n_36;
output n_104;
wire n_480;
wire n_113;
wire n_476;
wire n_758;
wire n_599;
wire n_187;
wire n_436;
wire n_684;
wire n_257;
wire n_390;
wire n_185;
wire n_285;
wire n_624;
wire n_618;
wire n_778;
wire n_800;
wire n_522;
wire n_485;
wire n_222;
wire n_750;
wire n_631;
wire n_287;
wire n_357;
wire n_503;
wire n_792;
wire n_386;
wire n_635;
wire n_673;
wire n_518;
wire n_254;
wire n_207;
wire n_665;
wire n_667;
wire n_577;
wire n_580;
wire n_469;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_759;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_718;
wire n_318;
wire n_355;
wire n_239;
wire n_669;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_761;
wire n_742;
wire n_112;
wire n_319;
wire n_364;
wire n_421;
wire n_555;
wire n_329;
wire n_766;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_169;
wire n_242;
wire n_376;
wire n_549;
wire n_571;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_752;
wire n_448;
wire n_545;
wire n_556;
wire n_341;
wire n_593;
wire n_232;
wire n_460;
wire n_773;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_537;
wire n_320;
wire n_551;
wire n_666;
wire n_560;
wire n_260;
wire n_660;
wire n_594;
wire n_186;
wire n_767;
wire n_138;
wire n_696;
wire n_704;
wire n_379;
wire n_374;
wire n_453;
wire n_647;
wire n_235;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_775;
wire n_161;
wire n_763;
wire n_189;
wire n_271;
wire n_489;
wire n_548;
wire n_427;
wire n_678;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_519;
wire n_564;
wire n_638;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_786;
wire n_512;
wire n_395;
wire n_332;
wire n_795;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_116;
wire n_625;
wire n_462;
wire n_289;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_716;
wire n_213;
wire n_478;
wire n_356;
wire n_584;
wire n_408;
wire n_553;
wire n_184;
wire n_372;
wire n_528;
wire n_578;
wire n_202;
wire n_495;
wire n_370;
wire n_384;
wire n_744;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_467;
wire n_327;
wire n_774;
wire n_106;
wire n_791;
wire n_466;
wire n_559;
wire n_636;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_726;
wire n_517;
wire n_683;
wire n_780;
wire n_174;
wire n_570;
wire n_675;
wire n_530;
wire n_535;
wire n_732;
wire n_784;
wire n_211;
wire n_281;
wire n_693;
wire n_496;
wire n_173;
wire n_468;
wire n_234;
wire n_746;
wire n_284;
wire n_153;
wire n_316;
wire n_532;
wire n_656;
wire n_755;
wire n_178;
wire n_409;
wire n_748;
wire n_781;
wire n_298;
wire n_523;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_796;
wire n_297;
wire n_801;
wire n_383;
wire n_529;
wire n_119;
wire n_310;
wire n_455;
wire n_504;
wire n_725;
wire n_164;
wire n_671;
wire n_231;
wire n_547;
wire n_659;
wire n_634;
wire n_682;
wire n_454;
wire n_122;
wire n_782;
wire n_443;
wire n_565;
wire n_760;
wire n_608;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_267;
wire n_218;
wire n_737;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_770;
wire n_745;
wire n_722;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_331;
wire n_182;
wire n_363;
wire n_417;
wire n_449;
wire n_607;
wire n_754;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_142;
wire n_561;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_783;
wire n_655;
wire n_654;
wire n_502;
wire n_527;
wire n_434;
wire n_505;
wire n_769;
wire n_600;
wire n_731;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_602;
wire n_402;
wire n_552;
wire n_617;
wire n_733;
wire n_171;
wire n_658;
wire n_676;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_146;
wire n_432;
wire n_226;
wire n_255;
wire n_286;
wire n_416;
wire n_790;
wire n_410;
wire n_120;
wire n_799;
wire n_751;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_695;
wire n_685;
wire n_165;
wire n_361;
wire n_632;
wire n_246;
wire n_176;
wire n_768;
wire n_412;
wire n_163;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_777;
wire n_501;
wire n_488;
wire n_251;
wire n_642;
wire n_613;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_702;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_734;
wire n_110;
wire n_392;
wire n_562;
wire n_150;
wire n_147;
wire n_288;
wire n_404;
wire n_598;
wire n_713;
wire n_735;
wire n_728;
wire n_756;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_569;
wire n_563;
wire n_785;
wire n_188;
wire n_269;
wire n_430;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_193;
wire n_397;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_649;
wire n_663;
wire n_749;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_707;
wire n_622;
wire n_470;
wire n_133;
wire n_494;
wire n_711;
wire n_377;
wire n_273;
wire n_723;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_265;
wire n_354;
wire n_720;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_730;
wire n_643;
wire n_747;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_779;
wire n_481;
wire n_148;
wire n_498;
wire n_691;
wire n_765;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_233;
wire n_487;
wire n_290;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_155;
wire n_243;
wire n_692;
wire n_789;
wire n_544;
wire n_268;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_738;
wire n_701;
wire n_309;
wire n_344;
wire n_229;
wire n_107;
wire n_482;
wire n_520;
wire n_633;
wire n_679;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_787;
wire n_262;
wire n_630;
wire n_689;
wire n_715;
wire n_134;
wire n_420;
wire n_336;
wire n_349;
wire n_612;
wire n_195;
wire n_438;
wire n_764;
wire n_794;
wire n_300;
wire n_252;
wire n_314;
wire n_283;
wire n_741;
wire n_753;
wire n_249;
wire n_623;
wire n_446;
wire n_721;
wire n_221;
wire n_681;
wire n_156;
wire n_359;
wire n_456;
wire n_717;
wire n_312;
wire n_183;
wire n_266;
wire n_712;
wire n_205;
wire n_433;
wire n_516;
wire n_177;
wire n_335;
wire n_313;
wire n_627;
wire n_739;
wire n_140;
wire n_418;
wire n_521;
wire n_422;
wire n_771;
wire n_219;
wire n_524;
wire n_705;
wire n_180;
wire n_212;
wire n_210;
wire n_575;
wire n_325;
wire n_762;
wire n_479;
wire n_338;
wire n_442;
wire n_740;
wire n_371;
wire n_698;
wire n_166;
wire n_541;
wire n_224;
wire n_151;
wire n_546;
wire n_587;
wire n_639;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_724;
wire n_440;
wire n_525;
wire n_644;
wire n_674;
wire n_152;
wire n_198;
wire n_793;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_414;
wire n_757;
wire n_123;
wire n_279;
wire n_686;
wire n_776;
wire n_543;
wire n_497;
wire n_514;
wire n_270;
wire n_507;
wire n_614;
wire n_305;
wire n_586;
wire n_772;
wire n_450;
wire n_788;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_465;
wire n_473;
wire n_719;
wire n_566;
wire n_474;
wire n_170;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_168;
wire n_175;
wire n_241;
wire n_687;
wire n_729;
wire n_646;
wire n_650;
wire n_710;
wire n_105;
wire n_743;
wire n_294;
wire n_393;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_500;
wire n_307;
wire n_601;
wire n_661;
wire n_463;
wire n_396;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_143;
wire n_192;
wire n_475;
wire n_554;
wire n_264;
wire n_798;
wire n_237;
wire n_668;
wire n_797;
NAND2xp5_ASAP7_75t_L g235 ( .A(n_0), .B(n_156), .Y(n_235) );
NAND2xp5_ASAP7_75t_L g117 ( .A(n_1), .B(n_118), .Y(n_117) );
NAND2xp5_ASAP7_75t_L g539 ( .A(n_2), .B(n_140), .Y(n_539) );
NAND2xp5_ASAP7_75t_L g510 ( .A(n_3), .B(n_158), .Y(n_510) );
INVx1_ASAP7_75t_L g147 ( .A(n_4), .Y(n_147) );
NAND2xp5_ASAP7_75t_L g139 ( .A(n_5), .B(n_140), .Y(n_139) );
NAND2xp33_ASAP7_75t_SL g226 ( .A(n_6), .B(n_146), .Y(n_226) );
INVx1_ASAP7_75t_L g207 ( .A(n_7), .Y(n_207) );
CKINVDCx16_ASAP7_75t_R g118 ( .A(n_8), .Y(n_118) );
AND2x2_ASAP7_75t_L g134 ( .A(n_9), .B(n_135), .Y(n_134) );
XNOR2xp5_ASAP7_75t_L g125 ( .A(n_10), .B(n_126), .Y(n_125) );
AND2x2_ASAP7_75t_L g520 ( .A(n_10), .B(n_223), .Y(n_520) );
AND2x2_ASAP7_75t_L g512 ( .A(n_11), .B(n_197), .Y(n_512) );
INVx2_ASAP7_75t_L g136 ( .A(n_12), .Y(n_136) );
NAND2xp5_ASAP7_75t_L g529 ( .A(n_13), .B(n_158), .Y(n_529) );
XNOR2xp5_ASAP7_75t_L g481 ( .A(n_14), .B(n_482), .Y(n_481) );
CKINVDCx16_ASAP7_75t_R g111 ( .A(n_15), .Y(n_111) );
AOI221x1_ASAP7_75t_L g220 ( .A1(n_16), .A2(n_149), .B1(n_221), .B2(n_223), .C(n_225), .Y(n_220) );
NAND2xp5_ASAP7_75t_SL g192 ( .A(n_17), .B(n_140), .Y(n_192) );
NAND2xp5_ASAP7_75t_SL g543 ( .A(n_18), .B(n_140), .Y(n_543) );
INVx1_ASAP7_75t_L g114 ( .A(n_19), .Y(n_114) );
AOI22xp33_ASAP7_75t_L g581 ( .A1(n_20), .A2(n_91), .B1(n_140), .B2(n_208), .Y(n_581) );
AOI21xp5_ASAP7_75t_L g148 ( .A1(n_21), .A2(n_149), .B(n_154), .Y(n_148) );
AOI221xp5_ASAP7_75t_SL g184 ( .A1(n_22), .A2(n_35), .B1(n_140), .B2(n_149), .C(n_185), .Y(n_184) );
NAND2xp5_ASAP7_75t_L g155 ( .A(n_23), .B(n_156), .Y(n_155) );
OR2x2_ASAP7_75t_L g137 ( .A(n_24), .B(n_90), .Y(n_137) );
OA21x2_ASAP7_75t_L g198 ( .A1(n_24), .A2(n_90), .B(n_136), .Y(n_198) );
NAND2xp5_ASAP7_75t_L g196 ( .A(n_25), .B(n_158), .Y(n_196) );
INVxp67_ASAP7_75t_L g219 ( .A(n_26), .Y(n_219) );
AND2x2_ASAP7_75t_L g180 ( .A(n_27), .B(n_170), .Y(n_180) );
AOI21xp5_ASAP7_75t_L g233 ( .A1(n_28), .A2(n_149), .B(n_234), .Y(n_233) );
AO21x2_ASAP7_75t_L g524 ( .A1(n_29), .A2(n_223), .B(n_525), .Y(n_524) );
NAND2xp5_ASAP7_75t_L g186 ( .A(n_30), .B(n_158), .Y(n_186) );
AOI21xp5_ASAP7_75t_L g507 ( .A1(n_31), .A2(n_149), .B(n_508), .Y(n_507) );
NAND2xp5_ASAP7_75t_L g538 ( .A(n_32), .B(n_158), .Y(n_538) );
AND2x2_ASAP7_75t_L g146 ( .A(n_33), .B(n_147), .Y(n_146) );
AND2x2_ASAP7_75t_L g150 ( .A(n_33), .B(n_151), .Y(n_150) );
INVx1_ASAP7_75t_L g215 ( .A(n_33), .Y(n_215) );
OR2x6_ASAP7_75t_L g112 ( .A(n_34), .B(n_113), .Y(n_112) );
XOR2xp5_ASAP7_75t_L g480 ( .A(n_36), .B(n_481), .Y(n_480) );
NAND2xp5_ASAP7_75t_L g511 ( .A(n_37), .B(n_140), .Y(n_511) );
AOI22xp5_ASAP7_75t_L g250 ( .A1(n_38), .A2(n_82), .B1(n_149), .B2(n_213), .Y(n_250) );
NAND2xp5_ASAP7_75t_L g559 ( .A(n_39), .B(n_158), .Y(n_559) );
AOI22xp5_ASAP7_75t_L g464 ( .A1(n_40), .A2(n_74), .B1(n_465), .B2(n_466), .Y(n_464) );
CKINVDCx20_ASAP7_75t_R g466 ( .A(n_40), .Y(n_466) );
NAND2xp5_ASAP7_75t_L g498 ( .A(n_41), .B(n_140), .Y(n_498) );
NAND2xp5_ASAP7_75t_L g178 ( .A(n_42), .B(n_156), .Y(n_178) );
CKINVDCx20_ASAP7_75t_R g796 ( .A(n_43), .Y(n_796) );
AOI21xp5_ASAP7_75t_L g515 ( .A1(n_44), .A2(n_149), .B(n_516), .Y(n_515) );
NAND2xp5_ASAP7_75t_SL g474 ( .A(n_45), .B(n_475), .Y(n_474) );
AND2x2_ASAP7_75t_L g238 ( .A(n_46), .B(n_170), .Y(n_238) );
NAND2xp5_ASAP7_75t_L g502 ( .A(n_47), .B(n_156), .Y(n_502) );
NAND2xp5_ASAP7_75t_L g188 ( .A(n_48), .B(n_170), .Y(n_188) );
NAND2xp5_ASAP7_75t_SL g526 ( .A(n_49), .B(n_140), .Y(n_526) );
OAI22xp5_ASAP7_75t_SL g462 ( .A1(n_50), .A2(n_463), .B1(n_464), .B2(n_467), .Y(n_462) );
CKINVDCx20_ASAP7_75t_R g467 ( .A(n_50), .Y(n_467) );
INVx1_ASAP7_75t_L g143 ( .A(n_51), .Y(n_143) );
INVx1_ASAP7_75t_L g153 ( .A(n_51), .Y(n_153) );
NAND2xp5_ASAP7_75t_L g518 ( .A(n_52), .B(n_158), .Y(n_518) );
AND2x2_ASAP7_75t_L g554 ( .A(n_53), .B(n_170), .Y(n_554) );
NAND2xp5_ASAP7_75t_SL g179 ( .A(n_54), .B(n_140), .Y(n_179) );
NAND2xp5_ASAP7_75t_L g517 ( .A(n_55), .B(n_156), .Y(n_517) );
NAND2xp5_ASAP7_75t_L g537 ( .A(n_56), .B(n_156), .Y(n_537) );
AND2x2_ASAP7_75t_L g171 ( .A(n_57), .B(n_170), .Y(n_171) );
NAND2xp5_ASAP7_75t_SL g519 ( .A(n_58), .B(n_140), .Y(n_519) );
NAND2xp5_ASAP7_75t_L g236 ( .A(n_59), .B(n_158), .Y(n_236) );
NAND2xp5_ASAP7_75t_SL g556 ( .A(n_60), .B(n_140), .Y(n_556) );
AOI21xp5_ASAP7_75t_L g535 ( .A1(n_61), .A2(n_149), .B(n_536), .Y(n_535) );
NAND2xp5_ASAP7_75t_L g167 ( .A(n_62), .B(n_156), .Y(n_167) );
AND2x2_ASAP7_75t_SL g199 ( .A(n_63), .B(n_135), .Y(n_199) );
AND2x2_ASAP7_75t_L g549 ( .A(n_64), .B(n_135), .Y(n_549) );
AOI21xp5_ASAP7_75t_L g175 ( .A1(n_65), .A2(n_149), .B(n_176), .Y(n_175) );
NAND2xp5_ASAP7_75t_L g157 ( .A(n_66), .B(n_158), .Y(n_157) );
AND2x2_ASAP7_75t_SL g251 ( .A(n_67), .B(n_197), .Y(n_251) );
NAND2xp5_ASAP7_75t_L g560 ( .A(n_68), .B(n_156), .Y(n_560) );
NAND2xp5_ASAP7_75t_L g530 ( .A(n_69), .B(n_156), .Y(n_530) );
AOI22xp5_ASAP7_75t_L g582 ( .A1(n_70), .A2(n_94), .B1(n_149), .B2(n_213), .Y(n_582) );
NAND2xp5_ASAP7_75t_L g546 ( .A(n_71), .B(n_158), .Y(n_546) );
INVx1_ASAP7_75t_L g145 ( .A(n_72), .Y(n_145) );
INVx1_ASAP7_75t_L g151 ( .A(n_72), .Y(n_151) );
NAND2xp5_ASAP7_75t_L g509 ( .A(n_73), .B(n_156), .Y(n_509) );
CKINVDCx20_ASAP7_75t_R g465 ( .A(n_74), .Y(n_465) );
AOI21xp5_ASAP7_75t_L g557 ( .A1(n_75), .A2(n_149), .B(n_558), .Y(n_557) );
AOI21xp5_ASAP7_75t_L g499 ( .A1(n_76), .A2(n_149), .B(n_500), .Y(n_499) );
AOI21xp5_ASAP7_75t_L g527 ( .A1(n_77), .A2(n_149), .B(n_528), .Y(n_527) );
AND2x2_ASAP7_75t_L g540 ( .A(n_78), .B(n_135), .Y(n_540) );
NAND2xp5_ASAP7_75t_SL g579 ( .A(n_79), .B(n_170), .Y(n_579) );
NAND2xp5_ASAP7_75t_SL g168 ( .A(n_80), .B(n_140), .Y(n_168) );
AOI22xp5_ASAP7_75t_L g249 ( .A1(n_81), .A2(n_84), .B1(n_140), .B2(n_208), .Y(n_249) );
INVx1_ASAP7_75t_L g115 ( .A(n_83), .Y(n_115) );
NAND2xp5_ASAP7_75t_L g195 ( .A(n_85), .B(n_156), .Y(n_195) );
NAND2xp5_ASAP7_75t_L g187 ( .A(n_86), .B(n_156), .Y(n_187) );
AND2x2_ASAP7_75t_L g503 ( .A(n_87), .B(n_197), .Y(n_503) );
CKINVDCx20_ASAP7_75t_R g799 ( .A(n_88), .Y(n_799) );
AOI21xp5_ASAP7_75t_L g164 ( .A1(n_89), .A2(n_149), .B(n_165), .Y(n_164) );
NAND2xp5_ASAP7_75t_L g166 ( .A(n_92), .B(n_158), .Y(n_166) );
AOI21xp5_ASAP7_75t_L g544 ( .A1(n_93), .A2(n_149), .B(n_545), .Y(n_544) );
NAND2xp5_ASAP7_75t_L g501 ( .A(n_95), .B(n_158), .Y(n_501) );
AOI22xp5_ASAP7_75t_L g482 ( .A1(n_96), .A2(n_103), .B1(n_483), .B2(n_484), .Y(n_482) );
CKINVDCx20_ASAP7_75t_R g483 ( .A(n_96), .Y(n_483) );
INVxp67_ASAP7_75t_L g222 ( .A(n_97), .Y(n_222) );
NAND2xp5_ASAP7_75t_L g237 ( .A(n_98), .B(n_140), .Y(n_237) );
NAND2xp5_ASAP7_75t_L g177 ( .A(n_99), .B(n_158), .Y(n_177) );
AOI21xp5_ASAP7_75t_L g193 ( .A1(n_100), .A2(n_149), .B(n_194), .Y(n_193) );
BUFx2_ASAP7_75t_L g548 ( .A(n_101), .Y(n_548) );
BUFx2_ASAP7_75t_L g123 ( .A(n_102), .Y(n_123) );
NAND2xp5_ASAP7_75t_L g478 ( .A(n_102), .B(n_474), .Y(n_478) );
CKINVDCx20_ASAP7_75t_R g484 ( .A(n_103), .Y(n_484) );
AOI21xp5_ASAP7_75t_L g104 ( .A1(n_105), .A2(n_119), .B(n_798), .Y(n_104) );
HB1xp67_ASAP7_75t_L g105 ( .A(n_106), .Y(n_105) );
BUFx3_ASAP7_75t_L g106 ( .A(n_107), .Y(n_106) );
INVx3_ASAP7_75t_L g801 ( .A(n_107), .Y(n_801) );
INVx2_ASAP7_75t_SL g107 ( .A(n_108), .Y(n_107) );
NAND2xp5_ASAP7_75t_SL g108 ( .A(n_109), .B(n_116), .Y(n_108) );
INVx3_ASAP7_75t_L g109 ( .A(n_110), .Y(n_109) );
BUFx2_ASAP7_75t_L g797 ( .A(n_110), .Y(n_797) );
OR2x2_ASAP7_75t_L g110 ( .A(n_111), .B(n_112), .Y(n_110) );
NAND2xp5_ASAP7_75t_L g472 ( .A(n_111), .B(n_473), .Y(n_472) );
AND2x6_ASAP7_75t_SL g489 ( .A(n_111), .B(n_112), .Y(n_489) );
OR2x6_ASAP7_75t_SL g791 ( .A(n_111), .B(n_473), .Y(n_791) );
CKINVDCx5p33_ASAP7_75t_R g473 ( .A(n_112), .Y(n_473) );
NAND2xp5_ASAP7_75t_L g113 ( .A(n_114), .B(n_115), .Y(n_113) );
INVx2_ASAP7_75t_L g116 ( .A(n_117), .Y(n_116) );
OA22x2_ASAP7_75t_L g119 ( .A1(n_120), .A2(n_124), .B1(n_478), .B2(n_479), .Y(n_119) );
CKINVDCx11_ASAP7_75t_R g120 ( .A(n_121), .Y(n_120) );
CKINVDCx20_ASAP7_75t_R g121 ( .A(n_122), .Y(n_121) );
HB1xp67_ASAP7_75t_L g122 ( .A(n_123), .Y(n_122) );
OAI21xp5_ASAP7_75t_L g124 ( .A1(n_125), .A2(n_468), .B(n_474), .Y(n_124) );
OAI22x1_ASAP7_75t_L g126 ( .A1(n_127), .A2(n_128), .B1(n_461), .B2(n_462), .Y(n_126) );
OAI22x1_ASAP7_75t_L g793 ( .A1(n_127), .A2(n_486), .B1(n_791), .B2(n_794), .Y(n_793) );
INVx4_ASAP7_75t_L g127 ( .A(n_128), .Y(n_127) );
OAI22xp5_ASAP7_75t_L g485 ( .A1(n_128), .A2(n_486), .B1(n_490), .B2(n_789), .Y(n_485) );
AND2x4_ASAP7_75t_L g128 ( .A(n_129), .B(n_372), .Y(n_128) );
NOR3xp33_ASAP7_75t_L g129 ( .A(n_130), .B(n_294), .C(n_344), .Y(n_129) );
NAND2xp5_ASAP7_75t_L g130 ( .A(n_131), .B(n_261), .Y(n_130) );
AOI221xp5_ASAP7_75t_L g131 ( .A1(n_132), .A2(n_181), .B1(n_200), .B2(n_243), .C(n_253), .Y(n_131) );
INVx1_ASAP7_75t_SL g343 ( .A(n_132), .Y(n_343) );
AND2x4_ASAP7_75t_SL g132 ( .A(n_133), .B(n_161), .Y(n_132) );
INVx2_ASAP7_75t_L g265 ( .A(n_133), .Y(n_265) );
OR2x2_ASAP7_75t_L g287 ( .A(n_133), .B(n_278), .Y(n_287) );
HB1xp67_ASAP7_75t_L g302 ( .A(n_133), .Y(n_302) );
INVx5_ASAP7_75t_L g309 ( .A(n_133), .Y(n_309) );
AND2x4_ASAP7_75t_L g315 ( .A(n_133), .B(n_173), .Y(n_315) );
AND2x2_ASAP7_75t_SL g318 ( .A(n_133), .B(n_245), .Y(n_318) );
OR2x2_ASAP7_75t_L g327 ( .A(n_133), .B(n_328), .Y(n_327) );
AND2x2_ASAP7_75t_L g334 ( .A(n_133), .B(n_162), .Y(n_334) );
AND2x2_ASAP7_75t_L g435 ( .A(n_133), .B(n_172), .Y(n_435) );
OR2x6_ASAP7_75t_L g133 ( .A(n_134), .B(n_138), .Y(n_133) );
BUFx6f_ASAP7_75t_L g170 ( .A(n_135), .Y(n_170) );
AND2x2_ASAP7_75t_SL g135 ( .A(n_136), .B(n_137), .Y(n_135) );
AND2x4_ASAP7_75t_L g160 ( .A(n_136), .B(n_137), .Y(n_160) );
AOI21xp5_ASAP7_75t_L g138 ( .A1(n_139), .A2(n_148), .B(n_160), .Y(n_138) );
AND2x4_ASAP7_75t_L g140 ( .A(n_141), .B(n_146), .Y(n_140) );
INVx1_ASAP7_75t_L g227 ( .A(n_141), .Y(n_227) );
AND2x4_ASAP7_75t_L g141 ( .A(n_142), .B(n_144), .Y(n_141) );
AND2x6_ASAP7_75t_L g156 ( .A(n_142), .B(n_151), .Y(n_156) );
INVx2_ASAP7_75t_L g142 ( .A(n_143), .Y(n_142) );
AND2x4_ASAP7_75t_L g158 ( .A(n_144), .B(n_153), .Y(n_158) );
INVx2_ASAP7_75t_L g144 ( .A(n_145), .Y(n_144) );
INVx5_ASAP7_75t_L g159 ( .A(n_146), .Y(n_159) );
AND2x2_ASAP7_75t_L g152 ( .A(n_147), .B(n_153), .Y(n_152) );
HB1xp67_ASAP7_75t_L g211 ( .A(n_147), .Y(n_211) );
AND2x6_ASAP7_75t_L g149 ( .A(n_150), .B(n_152), .Y(n_149) );
BUFx3_ASAP7_75t_L g212 ( .A(n_150), .Y(n_212) );
INVx2_ASAP7_75t_L g217 ( .A(n_151), .Y(n_217) );
AND2x4_ASAP7_75t_L g213 ( .A(n_152), .B(n_214), .Y(n_213) );
INVx2_ASAP7_75t_L g210 ( .A(n_153), .Y(n_210) );
AOI21xp5_ASAP7_75t_L g154 ( .A1(n_155), .A2(n_157), .B(n_159), .Y(n_154) );
NAND2xp5_ASAP7_75t_L g547 ( .A(n_156), .B(n_548), .Y(n_547) );
AOI21xp5_ASAP7_75t_L g165 ( .A1(n_159), .A2(n_166), .B(n_167), .Y(n_165) );
AOI21xp5_ASAP7_75t_L g176 ( .A1(n_159), .A2(n_177), .B(n_178), .Y(n_176) );
AOI21xp5_ASAP7_75t_L g185 ( .A1(n_159), .A2(n_186), .B(n_187), .Y(n_185) );
AOI21xp5_ASAP7_75t_L g194 ( .A1(n_159), .A2(n_195), .B(n_196), .Y(n_194) );
AOI21xp5_ASAP7_75t_L g234 ( .A1(n_159), .A2(n_235), .B(n_236), .Y(n_234) );
AOI21xp5_ASAP7_75t_L g500 ( .A1(n_159), .A2(n_501), .B(n_502), .Y(n_500) );
AOI21xp5_ASAP7_75t_L g508 ( .A1(n_159), .A2(n_509), .B(n_510), .Y(n_508) );
AOI21xp5_ASAP7_75t_L g516 ( .A1(n_159), .A2(n_517), .B(n_518), .Y(n_516) );
AOI21xp5_ASAP7_75t_L g528 ( .A1(n_159), .A2(n_529), .B(n_530), .Y(n_528) );
AOI21xp5_ASAP7_75t_L g536 ( .A1(n_159), .A2(n_537), .B(n_538), .Y(n_536) );
AOI21xp5_ASAP7_75t_L g545 ( .A1(n_159), .A2(n_546), .B(n_547), .Y(n_545) );
AOI21xp5_ASAP7_75t_L g558 ( .A1(n_159), .A2(n_559), .B(n_560), .Y(n_558) );
NOR2xp33_ASAP7_75t_L g206 ( .A(n_160), .B(n_207), .Y(n_206) );
NOR2xp33_ASAP7_75t_L g218 ( .A(n_160), .B(n_219), .Y(n_218) );
NOR2xp33_ASAP7_75t_L g221 ( .A(n_160), .B(n_222), .Y(n_221) );
NOR3xp33_ASAP7_75t_L g225 ( .A(n_160), .B(n_226), .C(n_227), .Y(n_225) );
AOI21xp5_ASAP7_75t_L g525 ( .A1(n_160), .A2(n_526), .B(n_527), .Y(n_525) );
AOI21xp5_ASAP7_75t_L g555 ( .A1(n_160), .A2(n_556), .B(n_557), .Y(n_555) );
INVx3_ASAP7_75t_SL g286 ( .A(n_161), .Y(n_286) );
AND2x2_ASAP7_75t_L g330 ( .A(n_161), .B(n_245), .Y(n_330) );
OAI21xp5_ASAP7_75t_L g333 ( .A1(n_161), .A2(n_334), .B(n_335), .Y(n_333) );
AND2x2_ASAP7_75t_L g371 ( .A(n_161), .B(n_309), .Y(n_371) );
AND2x4_ASAP7_75t_L g161 ( .A(n_162), .B(n_172), .Y(n_161) );
NAND2xp5_ASAP7_75t_L g252 ( .A(n_162), .B(n_173), .Y(n_252) );
OR2x2_ASAP7_75t_L g256 ( .A(n_162), .B(n_173), .Y(n_256) );
INVx1_ASAP7_75t_L g264 ( .A(n_162), .Y(n_264) );
HB1xp67_ASAP7_75t_L g276 ( .A(n_162), .Y(n_276) );
INVx2_ASAP7_75t_L g284 ( .A(n_162), .Y(n_284) );
NAND2xp5_ASAP7_75t_L g308 ( .A(n_162), .B(n_309), .Y(n_308) );
AND2x2_ASAP7_75t_L g393 ( .A(n_162), .B(n_278), .Y(n_393) );
AND2x2_ASAP7_75t_L g408 ( .A(n_162), .B(n_245), .Y(n_408) );
AO21x2_ASAP7_75t_L g162 ( .A1(n_163), .A2(n_169), .B(n_171), .Y(n_162) );
NAND2xp5_ASAP7_75t_L g163 ( .A(n_164), .B(n_168), .Y(n_163) );
AO21x2_ASAP7_75t_L g173 ( .A1(n_169), .A2(n_174), .B(n_180), .Y(n_173) );
AO21x2_ASAP7_75t_L g328 ( .A1(n_169), .A2(n_174), .B(n_180), .Y(n_328) );
AOI21x1_ASAP7_75t_L g505 ( .A1(n_169), .A2(n_506), .B(n_512), .Y(n_505) );
CKINVDCx5p33_ASAP7_75t_R g169 ( .A(n_170), .Y(n_169) );
OA21x2_ASAP7_75t_L g183 ( .A1(n_170), .A2(n_184), .B(n_188), .Y(n_183) );
AOI21xp5_ASAP7_75t_L g497 ( .A1(n_170), .A2(n_498), .B(n_499), .Y(n_497) );
AO21x2_ASAP7_75t_L g580 ( .A1(n_170), .A2(n_581), .B(n_582), .Y(n_580) );
INVx2_ASAP7_75t_L g172 ( .A(n_173), .Y(n_172) );
AND2x2_ASAP7_75t_L g277 ( .A(n_173), .B(n_278), .Y(n_277) );
HB1xp67_ASAP7_75t_L g348 ( .A(n_173), .Y(n_348) );
NAND2xp5_ASAP7_75t_L g174 ( .A(n_175), .B(n_179), .Y(n_174) );
NAND2xp5_ASAP7_75t_L g400 ( .A(n_181), .B(n_401), .Y(n_400) );
NOR2x1p5_ASAP7_75t_L g181 ( .A(n_182), .B(n_189), .Y(n_181) );
BUFx3_ASAP7_75t_L g182 ( .A(n_183), .Y(n_182) );
AND2x2_ASAP7_75t_L g229 ( .A(n_183), .B(n_230), .Y(n_229) );
NAND2xp5_ASAP7_75t_L g259 ( .A(n_183), .B(n_190), .Y(n_259) );
INVx1_ASAP7_75t_L g269 ( .A(n_183), .Y(n_269) );
INVx2_ASAP7_75t_L g292 ( .A(n_183), .Y(n_292) );
INVx2_ASAP7_75t_L g298 ( .A(n_183), .Y(n_298) );
HB1xp67_ASAP7_75t_L g368 ( .A(n_183), .Y(n_368) );
OR2x2_ASAP7_75t_L g399 ( .A(n_183), .B(n_190), .Y(n_399) );
OR2x2_ASAP7_75t_L g415 ( .A(n_189), .B(n_416), .Y(n_415) );
INVx2_ASAP7_75t_L g189 ( .A(n_190), .Y(n_189) );
AND2x4_ASAP7_75t_SL g203 ( .A(n_190), .B(n_204), .Y(n_203) );
AND2x4_ASAP7_75t_L g241 ( .A(n_190), .B(n_242), .Y(n_241) );
OR2x2_ASAP7_75t_L g279 ( .A(n_190), .B(n_280), .Y(n_279) );
OR2x2_ASAP7_75t_L g291 ( .A(n_190), .B(n_292), .Y(n_291) );
AND2x2_ASAP7_75t_L g304 ( .A(n_190), .B(n_270), .Y(n_304) );
OR2x2_ASAP7_75t_L g312 ( .A(n_190), .B(n_204), .Y(n_312) );
INVx2_ASAP7_75t_L g339 ( .A(n_190), .Y(n_339) );
INVx1_ASAP7_75t_L g357 ( .A(n_190), .Y(n_357) );
NOR2xp33_ASAP7_75t_R g390 ( .A(n_190), .B(n_230), .Y(n_390) );
OR2x6_ASAP7_75t_L g190 ( .A(n_191), .B(n_199), .Y(n_190) );
AOI21xp5_ASAP7_75t_L g191 ( .A1(n_192), .A2(n_193), .B(n_197), .Y(n_191) );
INVx2_ASAP7_75t_SL g247 ( .A(n_197), .Y(n_247) );
AOI21xp5_ASAP7_75t_L g542 ( .A1(n_197), .A2(n_543), .B(n_544), .Y(n_542) );
BUFx4f_ASAP7_75t_L g197 ( .A(n_198), .Y(n_197) );
INVx3_ASAP7_75t_L g224 ( .A(n_198), .Y(n_224) );
NAND2xp5_ASAP7_75t_SL g200 ( .A(n_201), .B(n_239), .Y(n_200) );
OAI22xp5_ASAP7_75t_L g281 ( .A1(n_201), .A2(n_282), .B1(n_285), .B2(n_288), .Y(n_281) );
OR2x2_ASAP7_75t_L g201 ( .A(n_202), .B(n_228), .Y(n_201) );
INVx1_ASAP7_75t_SL g202 ( .A(n_203), .Y(n_202) );
AND2x2_ASAP7_75t_L g296 ( .A(n_203), .B(n_297), .Y(n_296) );
AND2x2_ASAP7_75t_L g331 ( .A(n_203), .B(n_332), .Y(n_331) );
AND2x4_ASAP7_75t_L g410 ( .A(n_203), .B(n_388), .Y(n_410) );
INVx3_ASAP7_75t_L g242 ( .A(n_204), .Y(n_242) );
AND2x4_ASAP7_75t_L g270 ( .A(n_204), .B(n_271), .Y(n_270) );
NAND2xp5_ASAP7_75t_L g325 ( .A(n_204), .B(n_230), .Y(n_325) );
NAND2xp5_ASAP7_75t_L g337 ( .A(n_204), .B(n_292), .Y(n_337) );
AND2x2_ASAP7_75t_L g342 ( .A(n_204), .B(n_339), .Y(n_342) );
NAND2xp5_ASAP7_75t_L g379 ( .A(n_204), .B(n_229), .Y(n_379) );
INVx1_ASAP7_75t_L g449 ( .A(n_204), .Y(n_449) );
NAND2xp5_ASAP7_75t_L g460 ( .A(n_204), .B(n_367), .Y(n_460) );
AND2x4_ASAP7_75t_L g204 ( .A(n_205), .B(n_220), .Y(n_204) );
AOI22xp5_ASAP7_75t_L g205 ( .A1(n_206), .A2(n_208), .B1(n_213), .B2(n_218), .Y(n_205) );
AND2x4_ASAP7_75t_L g208 ( .A(n_209), .B(n_212), .Y(n_208) );
AND2x2_ASAP7_75t_L g209 ( .A(n_210), .B(n_211), .Y(n_209) );
NOR2x1p5_ASAP7_75t_L g214 ( .A(n_215), .B(n_216), .Y(n_214) );
INVx3_ASAP7_75t_L g216 ( .A(n_217), .Y(n_216) );
INVx3_ASAP7_75t_L g533 ( .A(n_223), .Y(n_533) );
INVx4_ASAP7_75t_L g223 ( .A(n_224), .Y(n_223) );
AOI21x1_ASAP7_75t_L g231 ( .A1(n_224), .A2(n_232), .B(n_238), .Y(n_231) );
AO21x2_ASAP7_75t_L g513 ( .A1(n_224), .A2(n_514), .B(n_520), .Y(n_513) );
INVx2_ASAP7_75t_L g228 ( .A(n_229), .Y(n_228) );
INVx1_ASAP7_75t_L g240 ( .A(n_230), .Y(n_240) );
NAND2xp5_ASAP7_75t_L g260 ( .A(n_230), .B(n_242), .Y(n_260) );
INVx2_ASAP7_75t_L g271 ( .A(n_230), .Y(n_271) );
AND2x2_ASAP7_75t_L g297 ( .A(n_230), .B(n_298), .Y(n_297) );
OR2x2_ASAP7_75t_L g313 ( .A(n_230), .B(n_292), .Y(n_313) );
HB1xp67_ASAP7_75t_L g332 ( .A(n_230), .Y(n_332) );
NAND2xp5_ASAP7_75t_L g338 ( .A(n_230), .B(n_339), .Y(n_338) );
INVx1_ASAP7_75t_L g402 ( .A(n_230), .Y(n_402) );
INVx3_ASAP7_75t_L g230 ( .A(n_231), .Y(n_230) );
NAND2xp5_ASAP7_75t_L g232 ( .A(n_233), .B(n_237), .Y(n_232) );
NAND2xp5_ASAP7_75t_L g239 ( .A(n_240), .B(n_241), .Y(n_239) );
NAND2xp5_ASAP7_75t_L g280 ( .A(n_240), .B(n_269), .Y(n_280) );
AOI221x1_ASAP7_75t_SL g374 ( .A1(n_241), .A2(n_375), .B1(n_378), .B2(n_380), .C(n_384), .Y(n_374) );
NAND2xp5_ASAP7_75t_L g422 ( .A(n_241), .B(n_423), .Y(n_422) );
AND2x2_ASAP7_75t_L g432 ( .A(n_241), .B(n_297), .Y(n_432) );
NAND2xp5_ASAP7_75t_L g453 ( .A(n_241), .B(n_454), .Y(n_453) );
OR2x2_ASAP7_75t_L g363 ( .A(n_242), .B(n_291), .Y(n_363) );
AND2x2_ASAP7_75t_L g401 ( .A(n_242), .B(n_402), .Y(n_401) );
INVx1_ASAP7_75t_SL g243 ( .A(n_244), .Y(n_243) );
OR2x2_ASAP7_75t_L g244 ( .A(n_245), .B(n_252), .Y(n_244) );
AND2x2_ASAP7_75t_L g254 ( .A(n_245), .B(n_255), .Y(n_254) );
INVx2_ASAP7_75t_L g349 ( .A(n_245), .Y(n_349) );
NOR2xp33_ASAP7_75t_L g354 ( .A(n_245), .B(n_265), .Y(n_354) );
AND2x4_ASAP7_75t_L g383 ( .A(n_245), .B(n_284), .Y(n_383) );
NAND2xp5_ASAP7_75t_SL g419 ( .A(n_245), .B(n_315), .Y(n_419) );
OR2x2_ASAP7_75t_L g437 ( .A(n_245), .B(n_368), .Y(n_437) );
NOR2xp33_ASAP7_75t_L g447 ( .A(n_245), .B(n_328), .Y(n_447) );
BUFx6f_ASAP7_75t_L g245 ( .A(n_246), .Y(n_245) );
INVx2_ASAP7_75t_L g278 ( .A(n_246), .Y(n_278) );
AOI21x1_ASAP7_75t_L g246 ( .A1(n_247), .A2(n_248), .B(n_251), .Y(n_246) );
NAND2xp5_ASAP7_75t_L g248 ( .A(n_249), .B(n_250), .Y(n_248) );
INVx1_ASAP7_75t_L g303 ( .A(n_252), .Y(n_303) );
OAI22xp5_ASAP7_75t_L g310 ( .A1(n_252), .A2(n_311), .B1(n_314), .B2(n_316), .Y(n_310) );
AND2x2_ASAP7_75t_L g253 ( .A(n_254), .B(n_257), .Y(n_253) );
INVx2_ASAP7_75t_L g266 ( .A(n_254), .Y(n_266) );
AND2x2_ASAP7_75t_L g405 ( .A(n_255), .B(n_265), .Y(n_405) );
AND2x2_ASAP7_75t_L g451 ( .A(n_255), .B(n_318), .Y(n_451) );
AND2x2_ASAP7_75t_L g456 ( .A(n_255), .B(n_307), .Y(n_456) );
INVx2_ASAP7_75t_L g255 ( .A(n_256), .Y(n_255) );
AOI32xp33_ASAP7_75t_L g425 ( .A1(n_257), .A2(n_327), .A3(n_407), .B1(n_426), .B2(n_428), .Y(n_425) );
INVx2_ASAP7_75t_L g257 ( .A(n_258), .Y(n_257) );
OR2x2_ASAP7_75t_L g258 ( .A(n_259), .B(n_260), .Y(n_258) );
INVx1_ASAP7_75t_L g293 ( .A(n_260), .Y(n_293) );
AOI211xp5_ASAP7_75t_SL g261 ( .A1(n_262), .A2(n_267), .B(n_272), .C(n_281), .Y(n_261) );
OAI21xp5_ASAP7_75t_L g262 ( .A1(n_263), .A2(n_265), .B(n_266), .Y(n_262) );
INVx1_ASAP7_75t_L g263 ( .A(n_264), .Y(n_263) );
NAND2xp5_ASAP7_75t_L g314 ( .A(n_264), .B(n_315), .Y(n_314) );
NAND2xp5_ASAP7_75t_L g282 ( .A(n_265), .B(n_283), .Y(n_282) );
INVx2_ASAP7_75t_L g445 ( .A(n_265), .Y(n_445) );
AND2x2_ASAP7_75t_L g355 ( .A(n_267), .B(n_356), .Y(n_355) );
AND2x2_ASAP7_75t_SL g267 ( .A(n_268), .B(n_270), .Y(n_267) );
HB1xp67_ASAP7_75t_L g455 ( .A(n_268), .Y(n_455) );
INVx1_ASAP7_75t_L g268 ( .A(n_269), .Y(n_268) );
INVxp67_ASAP7_75t_SL g324 ( .A(n_269), .Y(n_324) );
HB1xp67_ASAP7_75t_L g424 ( .A(n_269), .Y(n_424) );
INVx1_ASAP7_75t_L g321 ( .A(n_270), .Y(n_321) );
AND2x2_ASAP7_75t_L g387 ( .A(n_270), .B(n_388), .Y(n_387) );
NAND2xp5_ASAP7_75t_L g427 ( .A(n_270), .B(n_398), .Y(n_427) );
NOR2xp33_ASAP7_75t_L g272 ( .A(n_273), .B(n_279), .Y(n_272) );
INVx1_ASAP7_75t_L g273 ( .A(n_274), .Y(n_273) );
OAI21xp33_ASAP7_75t_L g353 ( .A1(n_274), .A2(n_354), .B(n_355), .Y(n_353) );
AND2x2_ASAP7_75t_SL g274 ( .A(n_275), .B(n_277), .Y(n_274) );
INVx1_ASAP7_75t_L g275 ( .A(n_276), .Y(n_275) );
AND2x2_ASAP7_75t_L g283 ( .A(n_278), .B(n_284), .Y(n_283) );
BUFx2_ASAP7_75t_L g307 ( .A(n_278), .Y(n_307) );
NAND2xp5_ASAP7_75t_L g376 ( .A(n_283), .B(n_377), .Y(n_376) );
INVx1_ASAP7_75t_L g414 ( .A(n_283), .Y(n_414) );
AND2x2_ASAP7_75t_L g444 ( .A(n_283), .B(n_445), .Y(n_444) );
HB1xp67_ASAP7_75t_L g421 ( .A(n_284), .Y(n_421) );
OR2x2_ASAP7_75t_L g285 ( .A(n_286), .B(n_287), .Y(n_285) );
NAND2xp5_ASAP7_75t_L g433 ( .A(n_286), .B(n_434), .Y(n_433) );
INVx1_ASAP7_75t_SL g361 ( .A(n_287), .Y(n_361) );
INVx1_ASAP7_75t_L g288 ( .A(n_289), .Y(n_288) );
AND2x4_ASAP7_75t_L g289 ( .A(n_290), .B(n_293), .Y(n_289) );
INVx2_ASAP7_75t_L g290 ( .A(n_291), .Y(n_290) );
OR2x2_ASAP7_75t_L g320 ( .A(n_291), .B(n_321), .Y(n_320) );
HB1xp67_ASAP7_75t_L g388 ( .A(n_292), .Y(n_388) );
AND2x2_ASAP7_75t_L g397 ( .A(n_293), .B(n_398), .Y(n_397) );
NAND2xp5_ASAP7_75t_L g294 ( .A(n_295), .B(n_317), .Y(n_294) );
AOI221xp5_ASAP7_75t_L g295 ( .A1(n_296), .A2(n_299), .B1(n_304), .B2(n_305), .C(n_310), .Y(n_295) );
INVx1_ASAP7_75t_L g416 ( .A(n_297), .Y(n_416) );
INVxp33_ASAP7_75t_SL g448 ( .A(n_297), .Y(n_448) );
AOI21xp5_ASAP7_75t_L g394 ( .A1(n_299), .A2(n_395), .B(n_403), .Y(n_394) );
INVx2_ASAP7_75t_L g299 ( .A(n_300), .Y(n_299) );
NAND2xp5_ASAP7_75t_SL g300 ( .A(n_301), .B(n_303), .Y(n_300) );
INVx1_ASAP7_75t_L g301 ( .A(n_302), .Y(n_301) );
NAND2xp5_ASAP7_75t_L g360 ( .A(n_303), .B(n_361), .Y(n_360) );
INVx2_ASAP7_75t_L g316 ( .A(n_304), .Y(n_316) );
AND2x2_ASAP7_75t_L g351 ( .A(n_304), .B(n_352), .Y(n_351) );
AND2x2_ASAP7_75t_L g370 ( .A(n_304), .B(n_371), .Y(n_370) );
AOI22xp33_ASAP7_75t_SL g431 ( .A1(n_304), .A2(n_432), .B1(n_433), .B2(n_436), .Y(n_431) );
INVx1_ASAP7_75t_L g305 ( .A(n_306), .Y(n_305) );
OR2x2_ASAP7_75t_L g306 ( .A(n_307), .B(n_308), .Y(n_306) );
OR2x2_ASAP7_75t_L g326 ( .A(n_307), .B(n_327), .Y(n_326) );
NAND2xp5_ASAP7_75t_L g365 ( .A(n_307), .B(n_315), .Y(n_365) );
AND2x4_ASAP7_75t_L g382 ( .A(n_309), .B(n_328), .Y(n_382) );
NAND2xp5_ASAP7_75t_L g429 ( .A(n_309), .B(n_383), .Y(n_429) );
AND2x2_ASAP7_75t_L g441 ( .A(n_309), .B(n_393), .Y(n_441) );
NAND2xp33_ASAP7_75t_L g426 ( .A(n_311), .B(n_427), .Y(n_426) );
OR2x2_ASAP7_75t_L g311 ( .A(n_312), .B(n_313), .Y(n_311) );
INVx1_ASAP7_75t_SL g369 ( .A(n_312), .Y(n_369) );
INVx1_ASAP7_75t_L g440 ( .A(n_313), .Y(n_440) );
INVx2_ASAP7_75t_SL g392 ( .A(n_315), .Y(n_392) );
AOI211xp5_ASAP7_75t_SL g317 ( .A1(n_318), .A2(n_319), .B(n_322), .C(n_340), .Y(n_317) );
INVx1_ASAP7_75t_L g319 ( .A(n_320), .Y(n_319) );
OAI211xp5_ASAP7_75t_L g322 ( .A1(n_323), .A2(n_326), .B(n_329), .C(n_333), .Y(n_322) );
OR2x6_ASAP7_75t_SL g323 ( .A(n_324), .B(n_325), .Y(n_323) );
INVx1_ASAP7_75t_L g352 ( .A(n_324), .Y(n_352) );
INVx1_ASAP7_75t_SL g377 ( .A(n_327), .Y(n_377) );
NOR2xp33_ASAP7_75t_L g436 ( .A(n_327), .B(n_437), .Y(n_436) );
NAND2xp5_ASAP7_75t_L g329 ( .A(n_330), .B(n_331), .Y(n_329) );
NAND2xp5_ASAP7_75t_L g341 ( .A(n_332), .B(n_342), .Y(n_341) );
INVx2_ASAP7_75t_SL g335 ( .A(n_336), .Y(n_335) );
OAI22xp33_ASAP7_75t_L g418 ( .A1(n_336), .A2(n_419), .B1(n_420), .B2(n_422), .Y(n_418) );
OR2x2_ASAP7_75t_L g336 ( .A(n_337), .B(n_338), .Y(n_336) );
NOR2xp33_ASAP7_75t_L g340 ( .A(n_341), .B(n_343), .Y(n_340) );
OAI211xp5_ASAP7_75t_SL g344 ( .A1(n_345), .A2(n_350), .B(n_353), .C(n_358), .Y(n_344) );
INVxp67_ASAP7_75t_L g345 ( .A(n_346), .Y(n_345) );
NOR2xp33_ASAP7_75t_L g346 ( .A(n_347), .B(n_349), .Y(n_346) );
INVx1_ASAP7_75t_L g347 ( .A(n_348), .Y(n_347) );
INVx1_ASAP7_75t_L g350 ( .A(n_351), .Y(n_350) );
INVx1_ASAP7_75t_L g356 ( .A(n_357), .Y(n_356) );
AOI221xp5_ASAP7_75t_L g358 ( .A1(n_359), .A2(n_362), .B1(n_364), .B2(n_366), .C(n_370), .Y(n_358) );
INVx1_ASAP7_75t_L g359 ( .A(n_360), .Y(n_359) );
INVx1_ASAP7_75t_SL g362 ( .A(n_363), .Y(n_362) );
INVx1_ASAP7_75t_L g364 ( .A(n_365), .Y(n_364) );
AND2x2_ASAP7_75t_L g366 ( .A(n_367), .B(n_369), .Y(n_366) );
HB1xp67_ASAP7_75t_L g367 ( .A(n_368), .Y(n_367) );
AOI222xp33_ASAP7_75t_L g450 ( .A1(n_369), .A2(n_451), .B1(n_452), .B2(n_456), .C1(n_457), .C2(n_459), .Y(n_450) );
INVx2_ASAP7_75t_L g385 ( .A(n_371), .Y(n_385) );
NOR3xp33_ASAP7_75t_L g372 ( .A(n_373), .B(n_411), .C(n_430), .Y(n_372) );
NAND2xp5_ASAP7_75t_L g373 ( .A(n_374), .B(n_394), .Y(n_373) );
INVx1_ASAP7_75t_L g375 ( .A(n_376), .Y(n_375) );
INVxp67_ASAP7_75t_L g378 ( .A(n_379), .Y(n_378) );
INVx1_ASAP7_75t_L g380 ( .A(n_381), .Y(n_380) );
NAND2xp5_ASAP7_75t_L g381 ( .A(n_382), .B(n_383), .Y(n_381) );
NAND2xp5_ASAP7_75t_L g420 ( .A(n_382), .B(n_421), .Y(n_420) );
NAND2xp5_ASAP7_75t_L g458 ( .A(n_383), .B(n_445), .Y(n_458) );
OAI22xp33_ASAP7_75t_L g384 ( .A1(n_385), .A2(n_386), .B1(n_389), .B2(n_391), .Y(n_384) );
INVx1_ASAP7_75t_SL g386 ( .A(n_387), .Y(n_386) );
INVxp33_ASAP7_75t_L g389 ( .A(n_390), .Y(n_389) );
NAND2xp5_ASAP7_75t_L g391 ( .A(n_392), .B(n_393), .Y(n_391) );
NOR2xp33_ASAP7_75t_L g413 ( .A(n_392), .B(n_414), .Y(n_413) );
NAND2xp5_ASAP7_75t_L g395 ( .A(n_396), .B(n_400), .Y(n_395) );
INVx1_ASAP7_75t_L g396 ( .A(n_397), .Y(n_396) );
INVx1_ASAP7_75t_SL g398 ( .A(n_399), .Y(n_398) );
OAI22xp5_ASAP7_75t_L g403 ( .A1(n_400), .A2(n_404), .B1(n_406), .B2(n_409), .Y(n_403) );
INVx2_ASAP7_75t_L g404 ( .A(n_405), .Y(n_404) );
INVx1_ASAP7_75t_L g406 ( .A(n_407), .Y(n_406) );
BUFx2_ASAP7_75t_L g407 ( .A(n_408), .Y(n_407) );
CKINVDCx16_ASAP7_75t_R g409 ( .A(n_410), .Y(n_409) );
OAI211xp5_ASAP7_75t_SL g411 ( .A1(n_412), .A2(n_415), .B(n_417), .C(n_425), .Y(n_411) );
INVx1_ASAP7_75t_L g412 ( .A(n_413), .Y(n_412) );
INVx1_ASAP7_75t_L g417 ( .A(n_418), .Y(n_417) );
INVxp67_ASAP7_75t_L g423 ( .A(n_424), .Y(n_423) );
INVx1_ASAP7_75t_L g428 ( .A(n_429), .Y(n_428) );
NAND3xp33_ASAP7_75t_L g430 ( .A(n_431), .B(n_438), .C(n_450), .Y(n_430) );
INVx2_ASAP7_75t_L g434 ( .A(n_435), .Y(n_434) );
OAI21xp5_ASAP7_75t_L g438 ( .A1(n_439), .A2(n_442), .B(n_449), .Y(n_438) );
AND2x2_ASAP7_75t_L g439 ( .A(n_440), .B(n_441), .Y(n_439) );
AOI21xp5_ASAP7_75t_L g442 ( .A1(n_443), .A2(n_446), .B(n_448), .Y(n_442) );
INVx1_ASAP7_75t_L g443 ( .A(n_444), .Y(n_443) );
INVx1_ASAP7_75t_L g446 ( .A(n_447), .Y(n_446) );
INVx1_ASAP7_75t_L g452 ( .A(n_453), .Y(n_452) );
INVx1_ASAP7_75t_L g454 ( .A(n_455), .Y(n_454) );
INVx1_ASAP7_75t_L g457 ( .A(n_458), .Y(n_457) );
INVx1_ASAP7_75t_L g459 ( .A(n_460), .Y(n_459) );
INVxp33_ASAP7_75t_SL g461 ( .A(n_462), .Y(n_461) );
CKINVDCx20_ASAP7_75t_R g463 ( .A(n_464), .Y(n_463) );
CKINVDCx11_ASAP7_75t_R g468 ( .A(n_469), .Y(n_468) );
INVx1_ASAP7_75t_SL g469 ( .A(n_470), .Y(n_469) );
INVx1_ASAP7_75t_SL g470 ( .A(n_471), .Y(n_470) );
BUFx2_ASAP7_75t_L g471 ( .A(n_472), .Y(n_471) );
BUFx3_ASAP7_75t_L g477 ( .A(n_472), .Y(n_477) );
BUFx2_ASAP7_75t_L g475 ( .A(n_476), .Y(n_475) );
CKINVDCx20_ASAP7_75t_R g476 ( .A(n_477), .Y(n_476) );
AO221x1_ASAP7_75t_L g479 ( .A1(n_480), .A2(n_485), .B1(n_792), .B2(n_793), .C(n_795), .Y(n_479) );
INVx1_ASAP7_75t_L g792 ( .A(n_480), .Y(n_792) );
CKINVDCx11_ASAP7_75t_R g486 ( .A(n_487), .Y(n_486) );
INVx3_ASAP7_75t_SL g487 ( .A(n_488), .Y(n_487) );
CKINVDCx5p33_ASAP7_75t_R g488 ( .A(n_489), .Y(n_488) );
INVx5_ASAP7_75t_L g794 ( .A(n_490), .Y(n_794) );
AND2x4_ASAP7_75t_L g490 ( .A(n_491), .B(n_693), .Y(n_490) );
NOR3xp33_ASAP7_75t_L g491 ( .A(n_492), .B(n_618), .C(n_654), .Y(n_491) );
NAND2xp5_ASAP7_75t_L g492 ( .A(n_493), .B(n_592), .Y(n_492) );
AOI211xp5_ASAP7_75t_L g493 ( .A1(n_494), .A2(n_521), .B(n_550), .C(n_575), .Y(n_493) );
AND2x2_ASAP7_75t_L g683 ( .A(n_494), .B(n_552), .Y(n_683) );
AND2x2_ASAP7_75t_L g494 ( .A(n_495), .B(n_504), .Y(n_494) );
NAND2xp5_ASAP7_75t_L g664 ( .A(n_495), .B(n_665), .Y(n_664) );
AND2x2_ASAP7_75t_L g716 ( .A(n_495), .B(n_598), .Y(n_716) );
AND2x2_ASAP7_75t_L g732 ( .A(n_495), .B(n_567), .Y(n_732) );
NAND2xp5_ASAP7_75t_L g741 ( .A(n_495), .B(n_742), .Y(n_741) );
NAND2x1p5_ASAP7_75t_L g765 ( .A(n_495), .B(n_766), .Y(n_765) );
INVx4_ASAP7_75t_L g495 ( .A(n_496), .Y(n_495) );
AND2x4_ASAP7_75t_SL g562 ( .A(n_496), .B(n_563), .Y(n_562) );
INVx1_ASAP7_75t_L g587 ( .A(n_496), .Y(n_587) );
AND2x2_ASAP7_75t_L g634 ( .A(n_496), .B(n_577), .Y(n_634) );
AND2x2_ASAP7_75t_L g653 ( .A(n_496), .B(n_504), .Y(n_653) );
BUFx2_ASAP7_75t_L g658 ( .A(n_496), .Y(n_658) );
AND2x2_ASAP7_75t_L g702 ( .A(n_496), .B(n_513), .Y(n_702) );
AND2x4_ASAP7_75t_L g774 ( .A(n_496), .B(n_775), .Y(n_774) );
NOR2x1_ASAP7_75t_L g786 ( .A(n_496), .B(n_566), .Y(n_786) );
OR2x6_ASAP7_75t_L g496 ( .A(n_497), .B(n_503), .Y(n_496) );
NAND2xp5_ASAP7_75t_L g612 ( .A(n_504), .B(n_613), .Y(n_612) );
INVx1_ASAP7_75t_L g705 ( .A(n_504), .Y(n_705) );
BUFx2_ASAP7_75t_L g754 ( .A(n_504), .Y(n_754) );
INVx1_ASAP7_75t_L g776 ( .A(n_504), .Y(n_776) );
AND2x2_ASAP7_75t_L g504 ( .A(n_505), .B(n_513), .Y(n_504) );
INVx3_ASAP7_75t_L g563 ( .A(n_505), .Y(n_563) );
HB1xp67_ASAP7_75t_L g742 ( .A(n_505), .Y(n_742) );
NAND2xp5_ASAP7_75t_L g506 ( .A(n_507), .B(n_511), .Y(n_506) );
INVx2_ASAP7_75t_L g566 ( .A(n_513), .Y(n_566) );
AND2x2_ASAP7_75t_L g567 ( .A(n_513), .B(n_563), .Y(n_567) );
INVx2_ASAP7_75t_L g642 ( .A(n_513), .Y(n_642) );
OR2x2_ASAP7_75t_L g649 ( .A(n_513), .B(n_598), .Y(n_649) );
NAND2xp5_ASAP7_75t_L g514 ( .A(n_515), .B(n_519), .Y(n_514) );
AND2x2_ASAP7_75t_L g604 ( .A(n_521), .B(n_605), .Y(n_604) );
AND2x2_ASAP7_75t_L g638 ( .A(n_521), .B(n_601), .Y(n_638) );
AND2x2_ASAP7_75t_L g521 ( .A(n_522), .B(n_531), .Y(n_521) );
AND2x2_ASAP7_75t_L g674 ( .A(n_522), .B(n_573), .Y(n_674) );
INVx1_ASAP7_75t_L g522 ( .A(n_523), .Y(n_522) );
AND2x2_ASAP7_75t_L g631 ( .A(n_523), .B(n_532), .Y(n_631) );
AND2x2_ASAP7_75t_L g750 ( .A(n_523), .B(n_541), .Y(n_750) );
INVx2_ASAP7_75t_L g523 ( .A(n_524), .Y(n_523) );
INVx1_ASAP7_75t_L g572 ( .A(n_524), .Y(n_572) );
INVx1_ASAP7_75t_L g590 ( .A(n_524), .Y(n_590) );
AND2x2_ASAP7_75t_L g646 ( .A(n_524), .B(n_532), .Y(n_646) );
AND2x2_ASAP7_75t_L g651 ( .A(n_524), .B(n_553), .Y(n_651) );
OR2x2_ASAP7_75t_L g714 ( .A(n_524), .B(n_541), .Y(n_714) );
HB1xp67_ASAP7_75t_L g723 ( .A(n_524), .Y(n_723) );
AND2x2_ASAP7_75t_L g552 ( .A(n_531), .B(n_553), .Y(n_552) );
INVx2_ASAP7_75t_L g591 ( .A(n_531), .Y(n_591) );
NOR2x1_ASAP7_75t_SL g531 ( .A(n_532), .B(n_541), .Y(n_531) );
AO21x1_ASAP7_75t_SL g532 ( .A1(n_533), .A2(n_534), .B(n_540), .Y(n_532) );
AO21x2_ASAP7_75t_L g574 ( .A1(n_533), .A2(n_534), .B(n_540), .Y(n_574) );
NAND2xp5_ASAP7_75t_L g534 ( .A(n_535), .B(n_539), .Y(n_534) );
AND2x2_ASAP7_75t_L g569 ( .A(n_541), .B(n_570), .Y(n_569) );
INVx2_ASAP7_75t_SL g617 ( .A(n_541), .Y(n_617) );
NAND2x1_ASAP7_75t_L g627 ( .A(n_541), .B(n_553), .Y(n_627) );
OR2x2_ASAP7_75t_L g632 ( .A(n_541), .B(n_570), .Y(n_632) );
BUFx2_ASAP7_75t_L g688 ( .A(n_541), .Y(n_688) );
AND2x2_ASAP7_75t_L g724 ( .A(n_541), .B(n_603), .Y(n_724) );
AND2x2_ASAP7_75t_L g735 ( .A(n_541), .B(n_573), .Y(n_735) );
OR2x6_ASAP7_75t_L g541 ( .A(n_542), .B(n_549), .Y(n_541) );
INVx1_ASAP7_75t_L g550 ( .A(n_551), .Y(n_550) );
AOI22xp5_ASAP7_75t_L g551 ( .A1(n_552), .A2(n_561), .B1(n_567), .B2(n_568), .Y(n_551) );
AOI22xp5_ASAP7_75t_L g781 ( .A1(n_552), .A2(n_732), .B1(n_782), .B2(n_787), .Y(n_781) );
INVx4_ASAP7_75t_L g570 ( .A(n_553), .Y(n_570) );
INVx2_ASAP7_75t_L g601 ( .A(n_553), .Y(n_601) );
HB1xp67_ASAP7_75t_L g672 ( .A(n_553), .Y(n_672) );
OR2x2_ASAP7_75t_L g687 ( .A(n_553), .B(n_573), .Y(n_687) );
OR2x2_ASAP7_75t_SL g713 ( .A(n_553), .B(n_714), .Y(n_713) );
OR2x6_ASAP7_75t_L g553 ( .A(n_554), .B(n_555), .Y(n_553) );
AND2x2_ASAP7_75t_SL g561 ( .A(n_562), .B(n_564), .Y(n_561) );
INVx2_ASAP7_75t_SL g594 ( .A(n_562), .Y(n_594) );
NAND2xp5_ASAP7_75t_L g647 ( .A(n_562), .B(n_648), .Y(n_647) );
AND2x2_ASAP7_75t_L g662 ( .A(n_562), .B(n_610), .Y(n_662) );
NAND2xp5_ASAP7_75t_L g699 ( .A(n_562), .B(n_700), .Y(n_699) );
INVx2_ASAP7_75t_L g584 ( .A(n_563), .Y(n_584) );
HB1xp67_ASAP7_75t_L g609 ( .A(n_563), .Y(n_609) );
AND2x2_ASAP7_75t_L g665 ( .A(n_563), .B(n_642), .Y(n_665) );
INVx1_ASAP7_75t_L g775 ( .A(n_563), .Y(n_775) );
INVx1_ASAP7_75t_L g564 ( .A(n_565), .Y(n_564) );
NOR2xp33_ASAP7_75t_L g586 ( .A(n_565), .B(n_587), .Y(n_586) );
NAND2xp5_ASAP7_75t_L g596 ( .A(n_565), .B(n_597), .Y(n_596) );
INVx1_ASAP7_75t_L g565 ( .A(n_566), .Y(n_565) );
AND2x2_ASAP7_75t_L g583 ( .A(n_566), .B(n_584), .Y(n_583) );
NAND2xp5_ASAP7_75t_L g715 ( .A(n_567), .B(n_716), .Y(n_715) );
AOI321xp33_ASAP7_75t_L g737 ( .A1(n_568), .A2(n_639), .A3(n_707), .B1(n_738), .B2(n_739), .C(n_743), .Y(n_737) );
AND2x2_ASAP7_75t_L g568 ( .A(n_569), .B(n_571), .Y(n_568) );
INVxp67_ASAP7_75t_SL g636 ( .A(n_569), .Y(n_636) );
AND2x2_ASAP7_75t_L g661 ( .A(n_569), .B(n_590), .Y(n_661) );
AND2x2_ASAP7_75t_L g736 ( .A(n_569), .B(n_646), .Y(n_736) );
INVx1_ASAP7_75t_L g605 ( .A(n_570), .Y(n_605) );
BUFx2_ASAP7_75t_L g615 ( .A(n_570), .Y(n_615) );
NOR2xp67_ASAP7_75t_L g722 ( .A(n_570), .B(n_723), .Y(n_722) );
INVx1_ASAP7_75t_SL g660 ( .A(n_571), .Y(n_660) );
AND2x2_ASAP7_75t_L g571 ( .A(n_572), .B(n_573), .Y(n_571) );
BUFx2_ASAP7_75t_L g667 ( .A(n_572), .Y(n_667) );
INVx2_ASAP7_75t_L g603 ( .A(n_573), .Y(n_603) );
HB1xp67_ASAP7_75t_L g626 ( .A(n_573), .Y(n_626) );
INVx3_ASAP7_75t_L g573 ( .A(n_574), .Y(n_573) );
AOI21xp33_ASAP7_75t_SL g575 ( .A1(n_576), .A2(n_585), .B(n_588), .Y(n_575) );
NOR2xp67_ASAP7_75t_L g719 ( .A(n_576), .B(n_720), .Y(n_719) );
INVx2_ASAP7_75t_L g576 ( .A(n_577), .Y(n_576) );
AND2x2_ASAP7_75t_L g577 ( .A(n_578), .B(n_583), .Y(n_577) );
INVx3_ASAP7_75t_L g610 ( .A(n_578), .Y(n_610) );
AND2x2_ASAP7_75t_L g641 ( .A(n_578), .B(n_642), .Y(n_641) );
AND2x4_ASAP7_75t_L g578 ( .A(n_579), .B(n_580), .Y(n_578) );
AND2x4_ASAP7_75t_L g598 ( .A(n_579), .B(n_580), .Y(n_598) );
INVx1_ASAP7_75t_L g681 ( .A(n_583), .Y(n_681) );
INVx1_ASAP7_75t_SL g766 ( .A(n_584), .Y(n_766) );
INVxp33_ASAP7_75t_L g585 ( .A(n_586), .Y(n_585) );
NAND2xp5_ASAP7_75t_SL g640 ( .A(n_587), .B(n_641), .Y(n_640) );
OR2x2_ASAP7_75t_L g692 ( .A(n_587), .B(n_649), .Y(n_692) );
OR2x2_ASAP7_75t_L g588 ( .A(n_589), .B(n_591), .Y(n_588) );
AND2x2_ASAP7_75t_L g696 ( .A(n_589), .B(n_697), .Y(n_696) );
NAND2xp5_ASAP7_75t_L g710 ( .A(n_589), .B(n_711), .Y(n_710) );
INVx3_ASAP7_75t_L g589 ( .A(n_590), .Y(n_589) );
NOR2xp33_ASAP7_75t_L g682 ( .A(n_590), .B(n_627), .Y(n_682) );
NOR4xp25_ASAP7_75t_L g777 ( .A(n_590), .B(n_621), .C(n_778), .D(n_779), .Y(n_777) );
OR2x2_ASAP7_75t_L g745 ( .A(n_591), .B(n_746), .Y(n_745) );
AOI221xp5_ASAP7_75t_L g592 ( .A1(n_593), .A2(n_599), .B1(n_604), .B2(n_606), .C(n_611), .Y(n_592) );
AND2x2_ASAP7_75t_L g593 ( .A(n_594), .B(n_595), .Y(n_593) );
AND2x2_ASAP7_75t_L g620 ( .A(n_595), .B(n_621), .Y(n_620) );
INVx2_ASAP7_75t_L g595 ( .A(n_596), .Y(n_595) );
OR2x2_ASAP7_75t_L g657 ( .A(n_596), .B(n_658), .Y(n_657) );
INVx2_ASAP7_75t_L g677 ( .A(n_597), .Y(n_677) );
INVx2_ASAP7_75t_L g597 ( .A(n_598), .Y(n_597) );
BUFx3_ASAP7_75t_L g700 ( .A(n_598), .Y(n_700) );
AND2x2_ASAP7_75t_L g707 ( .A(n_598), .B(n_708), .Y(n_707) );
INVxp67_ASAP7_75t_L g599 ( .A(n_600), .Y(n_599) );
NAND2xp5_ASAP7_75t_L g600 ( .A(n_601), .B(n_602), .Y(n_600) );
OR2x2_ASAP7_75t_L g644 ( .A(n_601), .B(n_645), .Y(n_644) );
INVxp67_ASAP7_75t_L g602 ( .A(n_603), .Y(n_602) );
NAND2xp5_ASAP7_75t_L g616 ( .A(n_603), .B(n_617), .Y(n_616) );
INVxp67_ASAP7_75t_L g606 ( .A(n_607), .Y(n_606) );
OR2x2_ASAP7_75t_L g607 ( .A(n_608), .B(n_610), .Y(n_607) );
INVx2_ASAP7_75t_L g621 ( .A(n_608), .Y(n_621) );
NAND2xp5_ASAP7_75t_L g690 ( .A(n_608), .B(n_691), .Y(n_690) );
INVx2_ASAP7_75t_L g608 ( .A(n_609), .Y(n_608) );
INVx2_ASAP7_75t_L g613 ( .A(n_610), .Y(n_613) );
OAI321xp33_ASAP7_75t_L g725 ( .A1(n_610), .A2(n_718), .A3(n_726), .B1(n_731), .B2(n_733), .C(n_737), .Y(n_725) );
NOR2xp33_ASAP7_75t_L g611 ( .A(n_612), .B(n_614), .Y(n_611) );
OR2x2_ASAP7_75t_L g680 ( .A(n_613), .B(n_681), .Y(n_680) );
OR2x2_ASAP7_75t_L g614 ( .A(n_615), .B(n_616), .Y(n_614) );
INVx1_ASAP7_75t_L g780 ( .A(n_616), .Y(n_780) );
NOR2xp33_ASAP7_75t_L g659 ( .A(n_617), .B(n_660), .Y(n_659) );
NAND2xp33_ASAP7_75t_SL g760 ( .A(n_617), .B(n_631), .Y(n_760) );
OAI211xp5_ASAP7_75t_L g618 ( .A1(n_619), .A2(n_622), .B(n_633), .C(n_637), .Y(n_618) );
INVxp67_ASAP7_75t_L g619 ( .A(n_620), .Y(n_619) );
NOR2x1_ASAP7_75t_L g622 ( .A(n_623), .B(n_628), .Y(n_622) );
INVx1_ASAP7_75t_L g623 ( .A(n_624), .Y(n_623) );
OR2x2_ASAP7_75t_L g624 ( .A(n_625), .B(n_627), .Y(n_624) );
INVx1_ASAP7_75t_L g625 ( .A(n_626), .Y(n_625) );
INVx1_ASAP7_75t_L g729 ( .A(n_626), .Y(n_729) );
INVx3_ASAP7_75t_L g668 ( .A(n_627), .Y(n_668) );
OR2x2_ASAP7_75t_L g771 ( .A(n_627), .B(n_645), .Y(n_771) );
INVx2_ASAP7_75t_L g628 ( .A(n_629), .Y(n_628) );
OAI22xp5_ASAP7_75t_L g712 ( .A1(n_629), .A2(n_713), .B1(n_715), .B2(n_717), .Y(n_712) );
OR2x2_ASAP7_75t_L g629 ( .A(n_630), .B(n_632), .Y(n_629) );
INVx1_ASAP7_75t_L g630 ( .A(n_631), .Y(n_630) );
INVx2_ASAP7_75t_SL g711 ( .A(n_632), .Y(n_711) );
OR2x2_ASAP7_75t_L g788 ( .A(n_632), .B(n_645), .Y(n_788) );
NAND2xp5_ASAP7_75t_L g633 ( .A(n_634), .B(n_635), .Y(n_633) );
INVx1_ASAP7_75t_L g635 ( .A(n_636), .Y(n_635) );
AOI21xp5_ASAP7_75t_SL g637 ( .A1(n_638), .A2(n_639), .B(n_643), .Y(n_637) );
INVx1_ASAP7_75t_L g639 ( .A(n_640), .Y(n_639) );
NAND2xp5_ASAP7_75t_L g757 ( .A(n_641), .B(n_658), .Y(n_757) );
AND2x2_ASAP7_75t_L g763 ( .A(n_641), .B(n_764), .Y(n_763) );
INVx1_ASAP7_75t_L g708 ( .A(n_642), .Y(n_708) );
OAI22xp5_ASAP7_75t_L g643 ( .A1(n_644), .A2(n_647), .B1(n_650), .B2(n_652), .Y(n_643) );
A2O1A1Ixp33_ASAP7_75t_L g689 ( .A1(n_645), .A2(n_688), .B(n_690), .C(n_692), .Y(n_689) );
INVx2_ASAP7_75t_SL g645 ( .A(n_646), .Y(n_645) );
NAND2xp5_ASAP7_75t_L g717 ( .A(n_648), .B(n_718), .Y(n_717) );
NAND2xp5_ASAP7_75t_L g762 ( .A(n_648), .B(n_740), .Y(n_762) );
INVx2_ASAP7_75t_SL g648 ( .A(n_649), .Y(n_648) );
INVx1_ASAP7_75t_L g650 ( .A(n_651), .Y(n_650) );
AND2x2_ASAP7_75t_L g734 ( .A(n_651), .B(n_735), .Y(n_734) );
INVx2_ASAP7_75t_SL g652 ( .A(n_653), .Y(n_652) );
A2O1A1Ixp33_ASAP7_75t_L g684 ( .A1(n_653), .A2(n_685), .B(n_688), .C(n_689), .Y(n_684) );
NAND3xp33_ASAP7_75t_SL g654 ( .A(n_655), .B(n_669), .C(n_684), .Y(n_654) );
AOI222xp33_ASAP7_75t_L g655 ( .A1(n_656), .A2(n_659), .B1(n_661), .B2(n_662), .C1(n_663), .C2(n_666), .Y(n_655) );
INVx1_ASAP7_75t_L g656 ( .A(n_657), .Y(n_656) );
INVx2_ASAP7_75t_L g718 ( .A(n_658), .Y(n_718) );
NAND2xp5_ASAP7_75t_L g744 ( .A(n_658), .B(n_691), .Y(n_744) );
INVx1_ASAP7_75t_L g663 ( .A(n_664), .Y(n_663) );
INVx1_ASAP7_75t_SL g678 ( .A(n_665), .Y(n_678) );
AND2x2_ASAP7_75t_L g666 ( .A(n_667), .B(n_668), .Y(n_666) );
OR2x2_ASAP7_75t_L g783 ( .A(n_667), .B(n_700), .Y(n_783) );
AOI22xp5_ASAP7_75t_L g758 ( .A1(n_668), .A2(n_759), .B1(n_761), .B2(n_763), .Y(n_758) );
AOI221xp5_ASAP7_75t_L g669 ( .A1(n_670), .A2(n_675), .B1(n_679), .B2(n_682), .C(n_683), .Y(n_669) );
INVx2_ASAP7_75t_SL g670 ( .A(n_671), .Y(n_670) );
OR2x2_ASAP7_75t_L g671 ( .A(n_672), .B(n_673), .Y(n_671) );
INVx1_ASAP7_75t_L g673 ( .A(n_674), .Y(n_673) );
INVx1_ASAP7_75t_L g675 ( .A(n_676), .Y(n_675) );
AOI21xp5_ASAP7_75t_SL g743 ( .A1(n_676), .A2(n_744), .B(n_745), .Y(n_743) );
OR2x2_ASAP7_75t_L g676 ( .A(n_677), .B(n_678), .Y(n_676) );
INVx2_ASAP7_75t_L g691 ( .A(n_677), .Y(n_691) );
AND2x2_ASAP7_75t_L g785 ( .A(n_677), .B(n_786), .Y(n_785) );
INVx1_ASAP7_75t_L g679 ( .A(n_680), .Y(n_679) );
INVx2_ASAP7_75t_L g769 ( .A(n_681), .Y(n_769) );
INVx1_ASAP7_75t_L g685 ( .A(n_686), .Y(n_685) );
HB1xp67_ASAP7_75t_L g686 ( .A(n_687), .Y(n_686) );
OR2x2_ASAP7_75t_L g698 ( .A(n_687), .B(n_688), .Y(n_698) );
INVx1_ASAP7_75t_L g751 ( .A(n_687), .Y(n_751) );
NOR3xp33_ASAP7_75t_L g693 ( .A(n_694), .B(n_725), .C(n_747), .Y(n_693) );
OAI211xp5_ASAP7_75t_L g694 ( .A1(n_695), .A2(n_699), .B(n_701), .C(n_706), .Y(n_694) );
INVx1_ASAP7_75t_L g695 ( .A(n_696), .Y(n_695) );
OAI21xp33_ASAP7_75t_L g701 ( .A1(n_696), .A2(n_702), .B(n_703), .Y(n_701) );
INVx1_ASAP7_75t_SL g697 ( .A(n_698), .Y(n_697) );
INVx1_ASAP7_75t_L g703 ( .A(n_704), .Y(n_703) );
HB1xp67_ASAP7_75t_L g704 ( .A(n_705), .Y(n_704) );
AOI211xp5_ASAP7_75t_L g706 ( .A1(n_707), .A2(n_709), .B(n_712), .C(n_719), .Y(n_706) );
INVx1_ASAP7_75t_L g709 ( .A(n_710), .Y(n_709) );
INVx2_ASAP7_75t_L g730 ( .A(n_713), .Y(n_730) );
INVxp67_ASAP7_75t_SL g755 ( .A(n_714), .Y(n_755) );
NAND2xp5_ASAP7_75t_L g753 ( .A(n_716), .B(n_754), .Y(n_753) );
INVx1_ASAP7_75t_L g778 ( .A(n_716), .Y(n_778) );
AND2x2_ASAP7_75t_L g768 ( .A(n_718), .B(n_769), .Y(n_768) );
INVx1_ASAP7_75t_L g738 ( .A(n_720), .Y(n_738) );
INVx2_ASAP7_75t_L g720 ( .A(n_721), .Y(n_720) );
AND2x2_ASAP7_75t_L g721 ( .A(n_722), .B(n_724), .Y(n_721) );
INVx1_ASAP7_75t_L g746 ( .A(n_722), .Y(n_746) );
INVx2_ASAP7_75t_SL g726 ( .A(n_727), .Y(n_726) );
AND2x4_ASAP7_75t_L g727 ( .A(n_728), .B(n_730), .Y(n_727) );
INVx1_ASAP7_75t_L g728 ( .A(n_729), .Y(n_728) );
INVx1_ASAP7_75t_SL g731 ( .A(n_732), .Y(n_731) );
NOR2xp33_ASAP7_75t_L g733 ( .A(n_734), .B(n_736), .Y(n_733) );
AOI221xp5_ASAP7_75t_L g767 ( .A1(n_734), .A2(n_768), .B1(n_770), .B2(n_772), .C(n_777), .Y(n_767) );
OAI21xp33_ASAP7_75t_SL g782 ( .A1(n_739), .A2(n_783), .B(n_784), .Y(n_782) );
INVx2_ASAP7_75t_SL g739 ( .A(n_740), .Y(n_739) );
INVx1_ASAP7_75t_L g740 ( .A(n_741), .Y(n_740) );
NAND4xp25_ASAP7_75t_L g747 ( .A(n_748), .B(n_758), .C(n_767), .D(n_781), .Y(n_747) );
AOI22xp5_ASAP7_75t_L g748 ( .A1(n_749), .A2(n_752), .B1(n_755), .B2(n_756), .Y(n_748) );
AND2x4_ASAP7_75t_L g749 ( .A(n_750), .B(n_751), .Y(n_749) );
INVx1_ASAP7_75t_L g752 ( .A(n_753), .Y(n_752) );
INVx1_ASAP7_75t_SL g756 ( .A(n_757), .Y(n_756) );
INVxp67_ASAP7_75t_L g759 ( .A(n_760), .Y(n_759) );
INVx1_ASAP7_75t_SL g761 ( .A(n_762), .Y(n_761) );
INVx1_ASAP7_75t_L g764 ( .A(n_765), .Y(n_764) );
INVx2_ASAP7_75t_L g770 ( .A(n_771), .Y(n_770) );
NAND2xp5_ASAP7_75t_L g772 ( .A(n_773), .B(n_776), .Y(n_772) );
INVx2_ASAP7_75t_L g773 ( .A(n_774), .Y(n_773) );
INVx1_ASAP7_75t_L g779 ( .A(n_780), .Y(n_779) );
INVx1_ASAP7_75t_L g784 ( .A(n_785), .Y(n_784) );
INVx2_ASAP7_75t_L g787 ( .A(n_788), .Y(n_787) );
INVx1_ASAP7_75t_SL g789 ( .A(n_790), .Y(n_789) );
CKINVDCx11_ASAP7_75t_R g790 ( .A(n_791), .Y(n_790) );
NOR2xp33_ASAP7_75t_L g795 ( .A(n_796), .B(n_797), .Y(n_795) );
NOR2xp33_ASAP7_75t_L g798 ( .A(n_799), .B(n_800), .Y(n_798) );
INVx1_ASAP7_75t_L g800 ( .A(n_801), .Y(n_800) );
endmodule