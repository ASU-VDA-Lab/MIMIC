module fake_jpeg_16170_n_148 (n_13, n_21, n_33, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_40, n_19, n_18, n_20, n_35, n_41, n_4, n_34, n_30, n_39, n_42, n_16, n_3, n_0, n_24, n_28, n_38, n_26, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_43, n_12, n_32, n_8, n_15, n_7, n_148);

input n_13;
input n_21;
input n_33;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_42;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_43;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_148;

wire n_117;
wire n_144;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_147;
wire n_73;
wire n_84;
wire n_59;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_49;
wire n_76;
wire n_127;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_103;
wire n_50;
wire n_124;
wire n_141;
wire n_57;
wire n_119;
wire n_69;
wire n_83;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_106;
wire n_111;
wire n_44;
wire n_143;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_78;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_54;
wire n_93;
wire n_91;
wire n_138;
wire n_101;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_97;
wire n_135;
wire n_62;
wire n_120;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

BUFx12f_ASAP7_75t_L g44 ( 
.A(n_14),
.Y(n_44)
);

BUFx5_ASAP7_75t_L g45 ( 
.A(n_7),
.Y(n_45)
);

INVx5_ASAP7_75t_L g46 ( 
.A(n_5),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_8),
.Y(n_47)
);

INVx2_ASAP7_75t_L g48 ( 
.A(n_27),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_41),
.Y(n_49)
);

INVx13_ASAP7_75t_L g50 ( 
.A(n_30),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_34),
.Y(n_51)
);

INVx6_ASAP7_75t_L g52 ( 
.A(n_2),
.Y(n_52)
);

INVx11_ASAP7_75t_L g53 ( 
.A(n_2),
.Y(n_53)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_38),
.Y(n_54)
);

BUFx12f_ASAP7_75t_L g55 ( 
.A(n_12),
.Y(n_55)
);

BUFx16f_ASAP7_75t_L g56 ( 
.A(n_11),
.Y(n_56)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_37),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_42),
.Y(n_58)
);

CKINVDCx20_ASAP7_75t_R g59 ( 
.A(n_10),
.Y(n_59)
);

BUFx2_ASAP7_75t_L g60 ( 
.A(n_25),
.Y(n_60)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_21),
.Y(n_61)
);

CKINVDCx20_ASAP7_75t_R g62 ( 
.A(n_3),
.Y(n_62)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_54),
.Y(n_63)
);

INVx4_ASAP7_75t_L g84 ( 
.A(n_63),
.Y(n_84)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_49),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g74 ( 
.A(n_64),
.Y(n_74)
);

INVx3_ASAP7_75t_L g65 ( 
.A(n_47),
.Y(n_65)
);

INVx3_ASAP7_75t_L g75 ( 
.A(n_65),
.Y(n_75)
);

INVx6_ASAP7_75t_L g66 ( 
.A(n_50),
.Y(n_66)
);

INVx5_ASAP7_75t_L g77 ( 
.A(n_66),
.Y(n_77)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_57),
.Y(n_67)
);

INVx2_ASAP7_75t_L g80 ( 
.A(n_67),
.Y(n_80)
);

INVx6_ASAP7_75t_L g68 ( 
.A(n_50),
.Y(n_68)
);

INVx5_ASAP7_75t_L g82 ( 
.A(n_68),
.Y(n_82)
);

INVx4_ASAP7_75t_L g69 ( 
.A(n_44),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_69),
.B(n_60),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_L g70 ( 
.A(n_62),
.B(n_0),
.Y(n_70)
);

AND2x2_ASAP7_75t_L g86 ( 
.A(n_70),
.B(n_0),
.Y(n_86)
);

CKINVDCx14_ASAP7_75t_R g71 ( 
.A(n_66),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_L g95 ( 
.A(n_71),
.B(n_55),
.Y(n_95)
);

AOI22xp5_ASAP7_75t_SL g72 ( 
.A1(n_65),
.A2(n_52),
.B1(n_46),
.B2(n_48),
.Y(n_72)
);

OAI22xp5_ASAP7_75t_SL g92 ( 
.A1(n_72),
.A2(n_78),
.B1(n_81),
.B2(n_55),
.Y(n_92)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_73),
.Y(n_87)
);

INVx6_ASAP7_75t_L g76 ( 
.A(n_64),
.Y(n_76)
);

INVx2_ASAP7_75t_L g101 ( 
.A(n_76),
.Y(n_101)
);

AOI22xp33_ASAP7_75t_L g78 ( 
.A1(n_69),
.A2(n_52),
.B1(n_53),
.B2(n_56),
.Y(n_78)
);

BUFx6f_ASAP7_75t_L g79 ( 
.A(n_68),
.Y(n_79)
);

INVx3_ASAP7_75t_L g91 ( 
.A(n_79),
.Y(n_91)
);

AOI22xp33_ASAP7_75t_SL g81 ( 
.A1(n_65),
.A2(n_56),
.B1(n_60),
.B2(n_47),
.Y(n_81)
);

HB1xp67_ASAP7_75t_L g83 ( 
.A(n_63),
.Y(n_83)
);

CKINVDCx20_ASAP7_75t_R g94 ( 
.A(n_83),
.Y(n_94)
);

BUFx6f_ASAP7_75t_L g85 ( 
.A(n_64),
.Y(n_85)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_85),
.Y(n_93)
);

AND2x2_ASAP7_75t_L g88 ( 
.A(n_86),
.B(n_1),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_L g106 ( 
.A(n_88),
.B(n_95),
.Y(n_106)
);

INVx2_ASAP7_75t_SL g89 ( 
.A(n_77),
.Y(n_89)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_89),
.Y(n_105)
);

AOI22xp33_ASAP7_75t_SL g90 ( 
.A1(n_75),
.A2(n_82),
.B1(n_49),
.B2(n_51),
.Y(n_90)
);

OAI22xp5_ASAP7_75t_SL g109 ( 
.A1(n_90),
.A2(n_97),
.B1(n_100),
.B2(n_104),
.Y(n_109)
);

CKINVDCx14_ASAP7_75t_R g111 ( 
.A(n_92),
.Y(n_111)
);

CKINVDCx16_ASAP7_75t_R g96 ( 
.A(n_73),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g113 ( 
.A(n_96),
.B(n_102),
.Y(n_113)
);

AOI22xp33_ASAP7_75t_L g97 ( 
.A1(n_74),
.A2(n_58),
.B1(n_51),
.B2(n_44),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_SL g98 ( 
.A(n_86),
.B(n_59),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_SL g112 ( 
.A(n_98),
.B(n_99),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_80),
.B(n_61),
.Y(n_99)
);

OAI22xp5_ASAP7_75t_L g100 ( 
.A1(n_84),
.A2(n_58),
.B1(n_22),
.B2(n_23),
.Y(n_100)
);

INVxp67_ASAP7_75t_L g102 ( 
.A(n_71),
.Y(n_102)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_83),
.Y(n_103)
);

CKINVDCx20_ASAP7_75t_R g108 ( 
.A(n_103),
.Y(n_108)
);

AOI22xp33_ASAP7_75t_SL g104 ( 
.A1(n_76),
.A2(n_45),
.B1(n_3),
.B2(n_4),
.Y(n_104)
);

OAI22xp5_ASAP7_75t_SL g107 ( 
.A1(n_97),
.A2(n_20),
.B1(n_43),
.B2(n_40),
.Y(n_107)
);

AOI22xp5_ASAP7_75t_L g117 ( 
.A1(n_107),
.A2(n_110),
.B1(n_115),
.B2(n_88),
.Y(n_117)
);

OAI22xp5_ASAP7_75t_SL g110 ( 
.A1(n_90),
.A2(n_18),
.B1(n_39),
.B2(n_36),
.Y(n_110)
);

INVx2_ASAP7_75t_L g114 ( 
.A(n_101),
.Y(n_114)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_114),
.Y(n_119)
);

OAI22xp5_ASAP7_75t_SL g115 ( 
.A1(n_87),
.A2(n_17),
.B1(n_35),
.B2(n_33),
.Y(n_115)
);

INVx5_ASAP7_75t_L g116 ( 
.A(n_105),
.Y(n_116)
);

AOI22xp5_ASAP7_75t_L g123 ( 
.A1(n_116),
.A2(n_117),
.B1(n_121),
.B2(n_89),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_L g118 ( 
.A(n_108),
.B(n_94),
.Y(n_118)
);

CKINVDCx20_ASAP7_75t_R g124 ( 
.A(n_118),
.Y(n_124)
);

CKINVDCx20_ASAP7_75t_R g120 ( 
.A(n_113),
.Y(n_120)
);

OAI21xp5_ASAP7_75t_L g126 ( 
.A1(n_120),
.A2(n_93),
.B(n_91),
.Y(n_126)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_112),
.Y(n_121)
);

MAJIxp5_ASAP7_75t_L g122 ( 
.A(n_117),
.B(n_111),
.C(n_106),
.Y(n_122)
);

MAJIxp5_ASAP7_75t_L g128 ( 
.A(n_122),
.B(n_125),
.C(n_107),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_123),
.B(n_126),
.Y(n_127)
);

XOR2xp5_ASAP7_75t_L g125 ( 
.A(n_116),
.B(n_109),
.Y(n_125)
);

XOR2xp5_ASAP7_75t_L g132 ( 
.A(n_128),
.B(n_129),
.Y(n_132)
);

XNOR2xp5_ASAP7_75t_SL g129 ( 
.A(n_125),
.B(n_110),
.Y(n_129)
);

CKINVDCx20_ASAP7_75t_R g130 ( 
.A(n_124),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_L g135 ( 
.A(n_130),
.B(n_131),
.Y(n_135)
);

CKINVDCx16_ASAP7_75t_R g131 ( 
.A(n_126),
.Y(n_131)
);

AO22x2_ASAP7_75t_SL g133 ( 
.A1(n_129),
.A2(n_127),
.B1(n_104),
.B2(n_119),
.Y(n_133)
);

OAI22xp5_ASAP7_75t_SL g137 ( 
.A1(n_133),
.A2(n_1),
.B1(n_5),
.B2(n_6),
.Y(n_137)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_130),
.Y(n_134)
);

OAI21xp5_ASAP7_75t_SL g136 ( 
.A1(n_134),
.A2(n_115),
.B(n_4),
.Y(n_136)
);

FAx1_ASAP7_75t_SL g138 ( 
.A(n_136),
.B(n_137),
.CI(n_135),
.CON(n_138),
.SN(n_138)
);

NAND2xp5_ASAP7_75t_L g139 ( 
.A(n_138),
.B(n_133),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_L g140 ( 
.A(n_139),
.B(n_138),
.Y(n_140)
);

MAJIxp5_ASAP7_75t_L g141 ( 
.A(n_140),
.B(n_132),
.C(n_19),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_L g142 ( 
.A(n_141),
.B(n_16),
.Y(n_142)
);

OAI21xp5_ASAP7_75t_L g143 ( 
.A1(n_142),
.A2(n_24),
.B(n_32),
.Y(n_143)
);

AOI21xp5_ASAP7_75t_SL g144 ( 
.A1(n_143),
.A2(n_15),
.B(n_31),
.Y(n_144)
);

INVxp67_ASAP7_75t_L g145 ( 
.A(n_144),
.Y(n_145)
);

A2O1A1Ixp33_ASAP7_75t_L g146 ( 
.A1(n_145),
.A2(n_13),
.B(n_29),
.C(n_28),
.Y(n_146)
);

XNOR2xp5_ASAP7_75t_L g147 ( 
.A(n_146),
.B(n_9),
.Y(n_147)
);

XOR2xp5_ASAP7_75t_L g148 ( 
.A(n_147),
.B(n_26),
.Y(n_148)
);


endmodule