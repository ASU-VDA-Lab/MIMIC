module real_jpeg_12761_n_12 (n_5, n_4, n_8, n_0, n_1, n_11, n_2, n_6, n_7, n_3, n_10, n_9, n_12);

input n_5;
input n_4;
input n_8;
input n_0;
input n_1;
input n_11;
input n_2;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_12;

wire n_108;
wire n_54;
wire n_37;
wire n_168;
wire n_73;
wire n_35;
wire n_38;
wire n_29;
wire n_91;
wire n_49;
wire n_114;
wire n_68;
wire n_146;
wire n_83;
wire n_78;
wire n_166;
wire n_176;
wire n_104;
wire n_194;
wire n_153;
wire n_161;
wire n_64;
wire n_177;
wire n_47;
wire n_131;
wire n_163;
wire n_22;
wire n_174;
wire n_87;
wire n_197;
wire n_40;
wire n_105;
wire n_173;
wire n_115;
wire n_98;
wire n_27;
wire n_56;
wire n_184;
wire n_48;
wire n_164;
wire n_140;
wire n_126;
wire n_13;
wire n_113;
wire n_120;
wire n_155;
wire n_93;
wire n_95;
wire n_141;
wire n_65;
wire n_33;
wire n_188;
wire n_139;
wire n_142;
wire n_175;
wire n_76;
wire n_178;
wire n_67;
wire n_79;
wire n_107;
wire n_156;
wire n_147;
wire n_189;
wire n_170;
wire n_66;
wire n_136;
wire n_28;
wire n_44;
wire n_62;
wire n_162;
wire n_121;
wire n_106;
wire n_160;
wire n_172;
wire n_45;
wire n_112;
wire n_42;
wire n_18;
wire n_145;
wire n_77;
wire n_109;
wire n_39;
wire n_122;
wire n_94;
wire n_26;
wire n_19;
wire n_148;
wire n_118;
wire n_17;
wire n_123;
wire n_116;
wire n_21;
wire n_50;
wire n_143;
wire n_196;
wire n_69;
wire n_186;
wire n_31;
wire n_137;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_165;
wire n_134;
wire n_72;
wire n_159;
wire n_171;
wire n_151;
wire n_183;
wire n_198;
wire n_192;
wire n_100;
wire n_23;
wire n_51;
wire n_14;
wire n_71;
wire n_90;
wire n_61;
wire n_110;
wire n_195;
wire n_117;
wire n_99;
wire n_193;
wire n_86;
wire n_70;
wire n_41;
wire n_74;
wire n_80;
wire n_32;
wire n_20;
wire n_150;
wire n_30;
wire n_158;
wire n_149;
wire n_15;
wire n_144;
wire n_130;
wire n_103;
wire n_43;
wire n_57;
wire n_157;
wire n_84;
wire n_82;
wire n_111;
wire n_132;
wire n_125;
wire n_185;
wire n_55;
wire n_180;
wire n_58;
wire n_52;
wire n_191;
wire n_63;
wire n_124;
wire n_24;
wire n_92;
wire n_75;
wire n_97;
wire n_187;
wire n_34;
wire n_190;
wire n_60;
wire n_46;
wire n_169;
wire n_88;
wire n_59;
wire n_128;
wire n_167;
wire n_179;
wire n_133;
wire n_138;
wire n_25;
wire n_53;
wire n_127;
wire n_119;
wire n_36;
wire n_102;
wire n_81;
wire n_85;
wire n_181;
wire n_101;
wire n_182;
wire n_96;
wire n_89;
wire n_16;

INVx4_ASAP7_75t_L g32 ( 
.A(n_0),
.Y(n_32)
);

INVx4_ASAP7_75t_L g29 ( 
.A(n_1),
.Y(n_29)
);

AOI22xp5_ASAP7_75t_SL g33 ( 
.A1(n_2),
.A2(n_34),
.B1(n_35),
.B2(n_38),
.Y(n_33)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_2),
.Y(n_38)
);

BUFx16f_ASAP7_75t_L g84 ( 
.A(n_3),
.Y(n_84)
);

OAI22xp5_ASAP7_75t_L g51 ( 
.A1(n_4),
.A2(n_28),
.B1(n_47),
.B2(n_52),
.Y(n_51)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_4),
.Y(n_52)
);

OAI22xp33_ASAP7_75t_SL g68 ( 
.A1(n_4),
.A2(n_24),
.B1(n_25),
.B2(n_52),
.Y(n_68)
);

AOI22xp5_ASAP7_75t_L g129 ( 
.A1(n_4),
.A2(n_34),
.B1(n_35),
.B2(n_52),
.Y(n_129)
);

OAI22xp5_ASAP7_75t_L g134 ( 
.A1(n_4),
.A2(n_52),
.B1(n_58),
.B2(n_59),
.Y(n_134)
);

INVx3_ASAP7_75t_L g60 ( 
.A(n_5),
.Y(n_60)
);

BUFx12f_ASAP7_75t_L g25 ( 
.A(n_6),
.Y(n_25)
);

AOI22xp5_ASAP7_75t_L g40 ( 
.A1(n_7),
.A2(n_34),
.B1(n_35),
.B2(n_41),
.Y(n_40)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_7),
.Y(n_41)
);

OAI22xp5_ASAP7_75t_SL g46 ( 
.A1(n_7),
.A2(n_28),
.B1(n_41),
.B2(n_47),
.Y(n_46)
);

AOI22xp33_ASAP7_75t_L g90 ( 
.A1(n_7),
.A2(n_24),
.B1(n_25),
.B2(n_41),
.Y(n_90)
);

OAI22xp5_ASAP7_75t_L g101 ( 
.A1(n_7),
.A2(n_41),
.B1(n_58),
.B2(n_59),
.Y(n_101)
);

BUFx12_ASAP7_75t_L g61 ( 
.A(n_8),
.Y(n_61)
);

BUFx2_ASAP7_75t_L g27 ( 
.A(n_9),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_10),
.Y(n_23)
);

OAI22xp5_ASAP7_75t_L g55 ( 
.A1(n_10),
.A2(n_23),
.B1(n_24),
.B2(n_25),
.Y(n_55)
);

AOI22xp5_ASAP7_75t_SL g77 ( 
.A1(n_10),
.A2(n_23),
.B1(n_28),
.B2(n_47),
.Y(n_77)
);

AOI22xp5_ASAP7_75t_L g87 ( 
.A1(n_10),
.A2(n_23),
.B1(n_58),
.B2(n_59),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_L g111 ( 
.A(n_10),
.B(n_45),
.Y(n_111)
);

AOI22xp5_ASAP7_75t_L g114 ( 
.A1(n_10),
.A2(n_23),
.B1(n_34),
.B2(n_35),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g135 ( 
.A(n_10),
.B(n_56),
.Y(n_135)
);

MAJIxp5_ASAP7_75t_L g142 ( 
.A(n_10),
.B(n_35),
.C(n_84),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_SL g149 ( 
.A(n_10),
.B(n_126),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_L g154 ( 
.A(n_10),
.B(n_85),
.Y(n_154)
);

O2A1O1Ixp33_ASAP7_75t_L g175 ( 
.A1(n_10),
.A2(n_24),
.B(n_61),
.C(n_176),
.Y(n_175)
);

INVx11_ASAP7_75t_L g37 ( 
.A(n_11),
.Y(n_37)
);

INVx1_ASAP7_75t_L g12 ( 
.A(n_13),
.Y(n_12)
);

OAI22xp5_ASAP7_75t_L g13 ( 
.A1(n_14),
.A2(n_117),
.B1(n_197),
.B2(n_198),
.Y(n_13)
);

CKINVDCx20_ASAP7_75t_R g197 ( 
.A(n_14),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_L g14 ( 
.A(n_15),
.B(n_115),
.Y(n_14)
);

NAND2xp5_ASAP7_75t_SL g15 ( 
.A(n_16),
.B(n_102),
.Y(n_15)
);

NOR2xp33_ASAP7_75t_L g116 ( 
.A(n_16),
.B(n_102),
.Y(n_116)
);

AOI22xp5_ASAP7_75t_L g16 ( 
.A1(n_17),
.A2(n_18),
.B1(n_69),
.B2(n_70),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_18),
.Y(n_17)
);

BUFx24_ASAP7_75t_SL g199 ( 
.A(n_18),
.Y(n_199)
);

FAx1_ASAP7_75t_SL g18 ( 
.A(n_19),
.B(n_43),
.CI(n_53),
.CON(n_18),
.SN(n_18)
);

NOR2xp33_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_30),
.Y(n_19)
);

OAI22xp5_ASAP7_75t_L g107 ( 
.A1(n_20),
.A2(n_21),
.B1(n_30),
.B2(n_31),
.Y(n_107)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_21),
.Y(n_20)
);

NOR2xp33_ASAP7_75t_SL g21 ( 
.A(n_22),
.B(n_28),
.Y(n_21)
);

MAJIxp5_ASAP7_75t_L g22 ( 
.A(n_23),
.B(n_24),
.C(n_26),
.Y(n_22)
);

OAI21xp33_ASAP7_75t_L g176 ( 
.A1(n_23),
.A2(n_58),
.B(n_62),
.Y(n_176)
);

OAI22xp5_ASAP7_75t_SL g45 ( 
.A1(n_24),
.A2(n_25),
.B1(n_26),
.B2(n_27),
.Y(n_45)
);

OAI22xp5_ASAP7_75t_L g66 ( 
.A1(n_24),
.A2(n_25),
.B1(n_61),
.B2(n_62),
.Y(n_66)
);

INVx8_ASAP7_75t_L g24 ( 
.A(n_25),
.Y(n_24)
);

AOI22xp33_ASAP7_75t_L g50 ( 
.A1(n_26),
.A2(n_27),
.B1(n_28),
.B2(n_47),
.Y(n_50)
);

INVx2_ASAP7_75t_L g26 ( 
.A(n_27),
.Y(n_26)
);

INVx13_ASAP7_75t_L g47 ( 
.A(n_28),
.Y(n_47)
);

BUFx12f_ASAP7_75t_L g28 ( 
.A(n_29),
.Y(n_28)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_31),
.Y(n_30)
);

OAI21xp5_ASAP7_75t_L g31 ( 
.A1(n_32),
.A2(n_33),
.B(n_39),
.Y(n_31)
);

NAND2xp5_ASAP7_75t_L g42 ( 
.A(n_32),
.B(n_35),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_32),
.B(n_40),
.Y(n_96)
);

INVx2_ASAP7_75t_L g126 ( 
.A(n_32),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_L g151 ( 
.A(n_32),
.B(n_129),
.Y(n_151)
);

AOI21xp5_ASAP7_75t_L g174 ( 
.A1(n_32),
.A2(n_42),
.B(n_114),
.Y(n_174)
);

OAI21xp5_ASAP7_75t_SL g94 ( 
.A1(n_33),
.A2(n_42),
.B(n_95),
.Y(n_94)
);

AO22x1_ASAP7_75t_L g85 ( 
.A1(n_34),
.A2(n_35),
.B1(n_83),
.B2(n_84),
.Y(n_85)
);

INVx4_ASAP7_75t_L g34 ( 
.A(n_35),
.Y(n_34)
);

NAND2xp5_ASAP7_75t_L g148 ( 
.A(n_35),
.B(n_149),
.Y(n_148)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_36),
.Y(n_35)
);

INVx5_ASAP7_75t_L g36 ( 
.A(n_37),
.Y(n_36)
);

NAND2xp5_ASAP7_75t_L g159 ( 
.A(n_39),
.B(n_160),
.Y(n_159)
);

OR2x2_ASAP7_75t_L g39 ( 
.A(n_40),
.B(n_42),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g113 ( 
.A(n_42),
.B(n_114),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_42),
.B(n_129),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_L g43 ( 
.A(n_44),
.B(n_48),
.Y(n_43)
);

NAND2xp5_ASAP7_75t_L g44 ( 
.A(n_45),
.B(n_46),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g49 ( 
.A(n_45),
.B(n_50),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_L g74 ( 
.A(n_45),
.B(n_51),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_SL g48 ( 
.A(n_49),
.B(n_51),
.Y(n_48)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_49),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_L g53 ( 
.A(n_54),
.B(n_63),
.Y(n_53)
);

NAND2x1_ASAP7_75t_SL g54 ( 
.A(n_55),
.B(n_56),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_SL g168 ( 
.A(n_55),
.B(n_169),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_L g92 ( 
.A(n_56),
.B(n_68),
.Y(n_92)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_57),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_L g65 ( 
.A(n_57),
.B(n_66),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_SL g110 ( 
.A(n_57),
.B(n_90),
.Y(n_110)
);

AOI22xp5_ASAP7_75t_SL g57 ( 
.A1(n_58),
.A2(n_59),
.B1(n_61),
.B2(n_62),
.Y(n_57)
);

AOI22xp33_ASAP7_75t_L g82 ( 
.A1(n_58),
.A2(n_59),
.B1(n_83),
.B2(n_84),
.Y(n_82)
);

INVx3_ASAP7_75t_L g58 ( 
.A(n_59),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_L g141 ( 
.A(n_59),
.B(n_142),
.Y(n_141)
);

INVx6_ASAP7_75t_L g59 ( 
.A(n_60),
.Y(n_59)
);

INVx8_ASAP7_75t_L g62 ( 
.A(n_61),
.Y(n_62)
);

INVxp67_ASAP7_75t_L g63 ( 
.A(n_64),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_64),
.B(n_110),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_SL g64 ( 
.A(n_65),
.B(n_67),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_SL g89 ( 
.A(n_65),
.B(n_90),
.Y(n_89)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_65),
.Y(n_169)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_68),
.Y(n_67)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_70),
.Y(n_69)
);

XOR2xp5_ASAP7_75t_L g70 ( 
.A(n_71),
.B(n_93),
.Y(n_70)
);

MAJIxp5_ASAP7_75t_L g71 ( 
.A(n_72),
.B(n_78),
.C(n_88),
.Y(n_71)
);

XOR2xp5_ASAP7_75t_L g104 ( 
.A(n_72),
.B(n_105),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_73),
.B(n_75),
.Y(n_72)
);

INVxp33_ASAP7_75t_L g73 ( 
.A(n_74),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_SL g75 ( 
.A(n_76),
.B(n_77),
.Y(n_75)
);

OAI22xp5_ASAP7_75t_SL g105 ( 
.A1(n_78),
.A2(n_79),
.B1(n_88),
.B2(n_106),
.Y(n_105)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_79),
.Y(n_78)
);

AOI21xp5_ASAP7_75t_L g79 ( 
.A1(n_80),
.A2(n_86),
.B(n_87),
.Y(n_79)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_81),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_L g98 ( 
.A(n_81),
.B(n_99),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_SL g133 ( 
.A(n_81),
.B(n_134),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_SL g171 ( 
.A(n_81),
.B(n_101),
.Y(n_171)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_82),
.B(n_85),
.Y(n_81)
);

INVx6_ASAP7_75t_L g83 ( 
.A(n_84),
.Y(n_83)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_85),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_SL g100 ( 
.A(n_85),
.B(n_101),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_SL g144 ( 
.A(n_85),
.B(n_134),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_SL g183 ( 
.A(n_85),
.B(n_99),
.Y(n_183)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_87),
.Y(n_99)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_88),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_SL g88 ( 
.A(n_89),
.B(n_91),
.Y(n_88)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_92),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_L g167 ( 
.A(n_92),
.B(n_168),
.Y(n_167)
);

XOR2xp5_ASAP7_75t_L g93 ( 
.A(n_94),
.B(n_97),
.Y(n_93)
);

INVxp67_ASAP7_75t_L g95 ( 
.A(n_96),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g112 ( 
.A(n_96),
.B(n_113),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_L g153 ( 
.A(n_96),
.B(n_128),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_SL g97 ( 
.A(n_98),
.B(n_100),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g143 ( 
.A(n_98),
.B(n_144),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_L g132 ( 
.A(n_100),
.B(n_133),
.Y(n_132)
);

MAJIxp5_ASAP7_75t_L g102 ( 
.A(n_103),
.B(n_107),
.C(n_108),
.Y(n_102)
);

OAI22xp5_ASAP7_75t_SL g193 ( 
.A1(n_103),
.A2(n_104),
.B1(n_194),
.B2(n_195),
.Y(n_193)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_104),
.Y(n_103)
);

XOR2xp5_ASAP7_75t_L g195 ( 
.A(n_107),
.B(n_108),
.Y(n_195)
);

MAJIxp5_ASAP7_75t_L g108 ( 
.A(n_109),
.B(n_111),
.C(n_112),
.Y(n_108)
);

XOR2xp5_ASAP7_75t_L g187 ( 
.A(n_109),
.B(n_188),
.Y(n_187)
);

XOR2xp5_ASAP7_75t_L g188 ( 
.A(n_111),
.B(n_112),
.Y(n_188)
);

NOR2xp33_ASAP7_75t_SL g150 ( 
.A(n_113),
.B(n_151),
.Y(n_150)
);

INVxp67_ASAP7_75t_L g125 ( 
.A(n_114),
.Y(n_125)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_116),
.Y(n_115)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_117),
.Y(n_198)
);

OAI21xp5_ASAP7_75t_SL g117 ( 
.A1(n_118),
.A2(n_191),
.B(n_196),
.Y(n_117)
);

AOI21xp5_ASAP7_75t_SL g118 ( 
.A1(n_119),
.A2(n_179),
.B(n_190),
.Y(n_118)
);

OAI21xp5_ASAP7_75t_SL g119 ( 
.A1(n_120),
.A2(n_163),
.B(n_178),
.Y(n_119)
);

AOI21xp5_ASAP7_75t_L g120 ( 
.A1(n_121),
.A2(n_145),
.B(n_162),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_SL g121 ( 
.A(n_122),
.B(n_139),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_L g162 ( 
.A(n_122),
.B(n_139),
.Y(n_162)
);

AOI22xp5_ASAP7_75t_L g122 ( 
.A1(n_123),
.A2(n_130),
.B1(n_131),
.B2(n_138),
.Y(n_122)
);

CKINVDCx16_ASAP7_75t_R g138 ( 
.A(n_123),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_L g123 ( 
.A(n_124),
.B(n_127),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_SL g124 ( 
.A(n_125),
.B(n_126),
.Y(n_124)
);

INVxp67_ASAP7_75t_L g127 ( 
.A(n_128),
.Y(n_127)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_131),
.Y(n_130)
);

OAI22xp5_ASAP7_75t_SL g131 ( 
.A1(n_132),
.A2(n_135),
.B1(n_136),
.B2(n_137),
.Y(n_131)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_132),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_L g182 ( 
.A(n_133),
.B(n_183),
.Y(n_182)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_135),
.Y(n_137)
);

MAJIxp5_ASAP7_75t_L g164 ( 
.A(n_135),
.B(n_136),
.C(n_138),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_L g139 ( 
.A(n_140),
.B(n_143),
.Y(n_139)
);

OAI22xp5_ASAP7_75t_SL g157 ( 
.A1(n_140),
.A2(n_141),
.B1(n_143),
.B2(n_158),
.Y(n_157)
);

CKINVDCx20_ASAP7_75t_R g140 ( 
.A(n_141),
.Y(n_140)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_143),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_L g170 ( 
.A(n_144),
.B(n_171),
.Y(n_170)
);

OAI21xp5_ASAP7_75t_L g145 ( 
.A1(n_146),
.A2(n_156),
.B(n_161),
.Y(n_145)
);

AOI21xp5_ASAP7_75t_L g146 ( 
.A1(n_147),
.A2(n_152),
.B(n_155),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_L g147 ( 
.A(n_148),
.B(n_150),
.Y(n_147)
);

INVxp67_ASAP7_75t_L g160 ( 
.A(n_151),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_SL g152 ( 
.A(n_153),
.B(n_154),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_L g155 ( 
.A(n_153),
.B(n_154),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_SL g156 ( 
.A(n_157),
.B(n_159),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_L g161 ( 
.A(n_157),
.B(n_159),
.Y(n_161)
);

NOR2xp33_ASAP7_75t_L g163 ( 
.A(n_164),
.B(n_165),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_L g178 ( 
.A(n_164),
.B(n_165),
.Y(n_178)
);

XOR2xp5_ASAP7_75t_L g165 ( 
.A(n_166),
.B(n_172),
.Y(n_165)
);

XOR2xp5_ASAP7_75t_L g166 ( 
.A(n_167),
.B(n_170),
.Y(n_166)
);

MAJIxp5_ASAP7_75t_L g189 ( 
.A(n_167),
.B(n_170),
.C(n_172),
.Y(n_189)
);

OAI22xp5_ASAP7_75t_L g172 ( 
.A1(n_173),
.A2(n_174),
.B1(n_175),
.B2(n_177),
.Y(n_172)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_174),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_L g184 ( 
.A(n_174),
.B(n_175),
.Y(n_184)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_175),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_SL g179 ( 
.A(n_180),
.B(n_189),
.Y(n_179)
);

NOR2xp33_ASAP7_75t_L g190 ( 
.A(n_180),
.B(n_189),
.Y(n_190)
);

XOR2xp5_ASAP7_75t_L g180 ( 
.A(n_181),
.B(n_187),
.Y(n_180)
);

OAI22xp5_ASAP7_75t_SL g181 ( 
.A1(n_182),
.A2(n_184),
.B1(n_185),
.B2(n_186),
.Y(n_181)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_182),
.Y(n_185)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_184),
.Y(n_186)
);

MAJIxp5_ASAP7_75t_L g192 ( 
.A(n_184),
.B(n_185),
.C(n_187),
.Y(n_192)
);

NOR2xp33_ASAP7_75t_L g191 ( 
.A(n_192),
.B(n_193),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_L g196 ( 
.A(n_192),
.B(n_193),
.Y(n_196)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_195),
.Y(n_194)
);


endmodule