module fake_netlist_6_2287_n_1909 (n_52, n_16, n_1, n_91, n_119, n_46, n_146, n_163, n_18, n_21, n_147, n_154, n_88, n_3, n_98, n_113, n_39, n_63, n_73, n_4, n_148, n_138, n_22, n_161, n_68, n_166, n_28, n_50, n_158, n_49, n_7, n_83, n_5, n_101, n_167, n_144, n_174, n_127, n_125, n_153, n_168, n_77, n_156, n_149, n_152, n_106, n_92, n_145, n_42, n_133, n_96, n_8, n_90, n_160, n_24, n_105, n_131, n_54, n_132, n_102, n_0, n_87, n_32, n_66, n_85, n_99, n_78, n_84, n_130, n_164, n_100, n_129, n_13, n_121, n_11, n_137, n_17, n_23, n_142, n_20, n_143, n_2, n_19, n_47, n_62, n_29, n_155, n_75, n_109, n_150, n_122, n_45, n_34, n_140, n_70, n_120, n_37, n_15, n_67, n_33, n_82, n_27, n_38, n_110, n_151, n_61, n_112, n_172, n_81, n_59, n_76, n_36, n_26, n_124, n_55, n_126, n_94, n_97, n_108, n_58, n_116, n_64, n_117, n_118, n_175, n_48, n_65, n_25, n_40, n_93, n_80, n_141, n_135, n_165, n_139, n_41, n_134, n_176, n_114, n_86, n_104, n_95, n_9, n_107, n_10, n_71, n_74, n_6, n_14, n_123, n_136, n_72, n_89, n_173, n_103, n_111, n_60, n_159, n_157, n_162, n_170, n_35, n_115, n_12, n_69, n_128, n_30, n_79, n_43, n_171, n_31, n_57, n_169, n_53, n_51, n_44, n_56, n_1909);

input n_52;
input n_16;
input n_1;
input n_91;
input n_119;
input n_46;
input n_146;
input n_163;
input n_18;
input n_21;
input n_147;
input n_154;
input n_88;
input n_3;
input n_98;
input n_113;
input n_39;
input n_63;
input n_73;
input n_4;
input n_148;
input n_138;
input n_22;
input n_161;
input n_68;
input n_166;
input n_28;
input n_50;
input n_158;
input n_49;
input n_7;
input n_83;
input n_5;
input n_101;
input n_167;
input n_144;
input n_174;
input n_127;
input n_125;
input n_153;
input n_168;
input n_77;
input n_156;
input n_149;
input n_152;
input n_106;
input n_92;
input n_145;
input n_42;
input n_133;
input n_96;
input n_8;
input n_90;
input n_160;
input n_24;
input n_105;
input n_131;
input n_54;
input n_132;
input n_102;
input n_0;
input n_87;
input n_32;
input n_66;
input n_85;
input n_99;
input n_78;
input n_84;
input n_130;
input n_164;
input n_100;
input n_129;
input n_13;
input n_121;
input n_11;
input n_137;
input n_17;
input n_23;
input n_142;
input n_20;
input n_143;
input n_2;
input n_19;
input n_47;
input n_62;
input n_29;
input n_155;
input n_75;
input n_109;
input n_150;
input n_122;
input n_45;
input n_34;
input n_140;
input n_70;
input n_120;
input n_37;
input n_15;
input n_67;
input n_33;
input n_82;
input n_27;
input n_38;
input n_110;
input n_151;
input n_61;
input n_112;
input n_172;
input n_81;
input n_59;
input n_76;
input n_36;
input n_26;
input n_124;
input n_55;
input n_126;
input n_94;
input n_97;
input n_108;
input n_58;
input n_116;
input n_64;
input n_117;
input n_118;
input n_175;
input n_48;
input n_65;
input n_25;
input n_40;
input n_93;
input n_80;
input n_141;
input n_135;
input n_165;
input n_139;
input n_41;
input n_134;
input n_176;
input n_114;
input n_86;
input n_104;
input n_95;
input n_9;
input n_107;
input n_10;
input n_71;
input n_74;
input n_6;
input n_14;
input n_123;
input n_136;
input n_72;
input n_89;
input n_173;
input n_103;
input n_111;
input n_60;
input n_159;
input n_157;
input n_162;
input n_170;
input n_35;
input n_115;
input n_12;
input n_69;
input n_128;
input n_30;
input n_79;
input n_43;
input n_171;
input n_31;
input n_57;
input n_169;
input n_53;
input n_51;
input n_44;
input n_56;

output n_1909;

wire n_992;
wire n_1671;
wire n_801;
wire n_1613;
wire n_1234;
wire n_1458;
wire n_1199;
wire n_1674;
wire n_741;
wire n_1027;
wire n_1351;
wire n_625;
wire n_1189;
wire n_223;
wire n_1212;
wire n_226;
wire n_208;
wire n_726;
wire n_212;
wire n_700;
wire n_1307;
wire n_1038;
wire n_578;
wire n_1581;
wire n_1003;
wire n_365;
wire n_1237;
wire n_1061;
wire n_1357;
wire n_1853;
wire n_783;
wire n_1738;
wire n_798;
wire n_188;
wire n_1575;
wire n_1854;
wire n_509;
wire n_1342;
wire n_245;
wire n_1209;
wire n_1348;
wire n_1387;
wire n_677;
wire n_1708;
wire n_805;
wire n_1151;
wire n_396;
wire n_1739;
wire n_350;
wire n_1380;
wire n_442;
wire n_480;
wire n_1402;
wire n_1691;
wire n_1688;
wire n_1009;
wire n_1743;
wire n_1160;
wire n_883;
wire n_1238;
wire n_1724;
wire n_1032;
wire n_1247;
wire n_1547;
wire n_1553;
wire n_893;
wire n_1099;
wire n_1264;
wire n_1192;
wire n_471;
wire n_1844;
wire n_424;
wire n_1700;
wire n_1555;
wire n_1415;
wire n_1370;
wire n_1786;
wire n_369;
wire n_287;
wire n_415;
wire n_830;
wire n_230;
wire n_461;
wire n_873;
wire n_383;
wire n_1285;
wire n_1371;
wire n_200;
wire n_447;
wire n_1803;
wire n_1172;
wire n_852;
wire n_229;
wire n_1590;
wire n_1532;
wire n_1393;
wire n_1517;
wire n_1867;
wire n_1704;
wire n_1078;
wire n_250;
wire n_544;
wire n_1711;
wire n_1140;
wire n_1444;
wire n_1670;
wire n_1603;
wire n_1579;
wire n_1263;
wire n_836;
wire n_375;
wire n_522;
wire n_1261;
wire n_945;
wire n_1649;
wire n_1903;
wire n_1511;
wire n_1143;
wire n_1422;
wire n_1232;
wire n_1772;
wire n_1572;
wire n_616;
wire n_658;
wire n_1874;
wire n_1119;
wire n_428;
wire n_1433;
wire n_1902;
wire n_1842;
wire n_1620;
wire n_1735;
wire n_1541;
wire n_1300;
wire n_641;
wire n_822;
wire n_693;
wire n_1313;
wire n_1056;
wire n_758;
wire n_516;
wire n_1455;
wire n_1163;
wire n_1180;
wire n_943;
wire n_1798;
wire n_1550;
wire n_491;
wire n_1591;
wire n_772;
wire n_1344;
wire n_666;
wire n_371;
wire n_940;
wire n_770;
wire n_567;
wire n_1781;
wire n_405;
wire n_213;
wire n_538;
wire n_1106;
wire n_886;
wire n_1471;
wire n_343;
wire n_953;
wire n_1094;
wire n_1345;
wire n_1820;
wire n_494;
wire n_539;
wire n_493;
wire n_454;
wire n_1421;
wire n_638;
wire n_1404;
wire n_1211;
wire n_381;
wire n_887;
wire n_1660;
wire n_1280;
wire n_713;
wire n_1400;
wire n_1467;
wire n_976;
wire n_224;
wire n_1445;
wire n_1526;
wire n_1560;
wire n_734;
wire n_1088;
wire n_1894;
wire n_196;
wire n_1231;
wire n_917;
wire n_574;
wire n_907;
wire n_1446;
wire n_659;
wire n_1815;
wire n_407;
wire n_913;
wire n_1658;
wire n_808;
wire n_867;
wire n_1230;
wire n_473;
wire n_1193;
wire n_1054;
wire n_559;
wire n_1333;
wire n_1648;
wire n_1644;
wire n_1558;
wire n_1732;
wire n_281;
wire n_551;
wire n_699;
wire n_564;
wire n_451;
wire n_824;
wire n_279;
wire n_686;
wire n_757;
wire n_594;
wire n_1641;
wire n_577;
wire n_1843;
wire n_619;
wire n_1367;
wire n_1336;
wire n_521;
wire n_572;
wire n_395;
wire n_813;
wire n_1481;
wire n_323;
wire n_606;
wire n_1441;
wire n_818;
wire n_1123;
wire n_1309;
wire n_513;
wire n_645;
wire n_1381;
wire n_331;
wire n_1699;
wire n_916;
wire n_483;
wire n_608;
wire n_261;
wire n_630;
wire n_541;
wire n_512;
wire n_433;
wire n_792;
wire n_476;
wire n_1328;
wire n_219;
wire n_1907;
wire n_264;
wire n_263;
wire n_1162;
wire n_860;
wire n_1530;
wire n_788;
wire n_939;
wire n_1543;
wire n_821;
wire n_938;
wire n_1302;
wire n_1068;
wire n_1599;
wire n_329;
wire n_982;
wire n_549;
wire n_1762;
wire n_1075;
wire n_408;
wire n_932;
wire n_237;
wire n_1876;
wire n_1895;
wire n_1697;
wire n_243;
wire n_979;
wire n_1873;
wire n_905;
wire n_1866;
wire n_1680;
wire n_322;
wire n_993;
wire n_689;
wire n_354;
wire n_1330;
wire n_1413;
wire n_1605;
wire n_1278;
wire n_547;
wire n_558;
wire n_1064;
wire n_1396;
wire n_634;
wire n_966;
wire n_764;
wire n_1663;
wire n_692;
wire n_733;
wire n_1793;
wire n_1233;
wire n_1289;
wire n_487;
wire n_241;
wire n_1107;
wire n_1014;
wire n_1290;
wire n_1703;
wire n_882;
wire n_1354;
wire n_586;
wire n_423;
wire n_1865;
wire n_1875;
wire n_1701;
wire n_318;
wire n_1111;
wire n_1713;
wire n_715;
wire n_1251;
wire n_1265;
wire n_1726;
wire n_530;
wire n_1563;
wire n_277;
wire n_618;
wire n_1297;
wire n_1662;
wire n_1312;
wire n_199;
wire n_1167;
wire n_1359;
wire n_674;
wire n_871;
wire n_922;
wire n_268;
wire n_1335;
wire n_1760;
wire n_210;
wire n_1069;
wire n_1664;
wire n_1722;
wire n_612;
wire n_178;
wire n_247;
wire n_1165;
wire n_355;
wire n_702;
wire n_347;
wire n_1175;
wire n_328;
wire n_1386;
wire n_1896;
wire n_429;
wire n_1747;
wire n_1012;
wire n_195;
wire n_780;
wire n_675;
wire n_903;
wire n_1540;
wire n_1802;
wire n_1504;
wire n_286;
wire n_254;
wire n_1655;
wire n_242;
wire n_835;
wire n_928;
wire n_1214;
wire n_690;
wire n_850;
wire n_1801;
wire n_1886;
wire n_1654;
wire n_816;
wire n_1157;
wire n_1750;
wire n_1462;
wire n_1188;
wire n_1752;
wire n_877;
wire n_1813;
wire n_604;
wire n_825;
wire n_728;
wire n_1063;
wire n_1588;
wire n_267;
wire n_1124;
wire n_1624;
wire n_515;
wire n_598;
wire n_696;
wire n_1515;
wire n_961;
wire n_437;
wire n_1082;
wire n_1317;
wire n_593;
wire n_514;
wire n_687;
wire n_697;
wire n_890;
wire n_637;
wire n_701;
wire n_295;
wire n_950;
wire n_388;
wire n_190;
wire n_484;
wire n_1709;
wire n_1825;
wire n_1757;
wire n_1796;
wire n_1792;
wire n_891;
wire n_1412;
wire n_949;
wire n_1630;
wire n_678;
wire n_283;
wire n_507;
wire n_968;
wire n_909;
wire n_1369;
wire n_881;
wire n_1008;
wire n_760;
wire n_1546;
wire n_590;
wire n_362;
wire n_462;
wire n_1033;
wire n_1052;
wire n_1296;
wire n_304;
wire n_694;
wire n_1294;
wire n_1420;
wire n_1634;
wire n_595;
wire n_627;
wire n_297;
wire n_1767;
wire n_1779;
wire n_524;
wire n_1465;
wire n_342;
wire n_1858;
wire n_1044;
wire n_1712;
wire n_1391;
wire n_449;
wire n_1523;
wire n_1208;
wire n_1164;
wire n_1295;
wire n_1627;
wire n_1072;
wire n_1527;
wire n_1495;
wire n_1438;
wire n_495;
wire n_815;
wire n_1100;
wire n_585;
wire n_1487;
wire n_840;
wire n_874;
wire n_1756;
wire n_1128;
wire n_382;
wire n_673;
wire n_1071;
wire n_1067;
wire n_1565;
wire n_1493;
wire n_898;
wire n_255;
wire n_284;
wire n_865;
wire n_925;
wire n_1101;
wire n_1026;
wire n_1880;
wire n_289;
wire n_1364;
wire n_615;
wire n_1249;
wire n_1293;
wire n_1127;
wire n_1512;
wire n_1451;
wire n_320;
wire n_639;
wire n_963;
wire n_794;
wire n_727;
wire n_894;
wire n_1839;
wire n_685;
wire n_1765;
wire n_353;
wire n_605;
wire n_1514;
wire n_1863;
wire n_826;
wire n_1646;
wire n_872;
wire n_1139;
wire n_1714;
wire n_718;
wire n_1018;
wire n_1521;
wire n_1366;
wire n_542;
wire n_847;
wire n_644;
wire n_682;
wire n_851;
wire n_305;
wire n_996;
wire n_532;
wire n_1308;
wire n_1376;
wire n_1513;
wire n_413;
wire n_791;
wire n_510;
wire n_837;
wire n_1488;
wire n_1808;
wire n_948;
wire n_704;
wire n_977;
wire n_1005;
wire n_536;
wire n_1788;
wire n_622;
wire n_1469;
wire n_1838;
wire n_1835;
wire n_1776;
wire n_1766;
wire n_581;
wire n_765;
wire n_432;
wire n_987;
wire n_1492;
wire n_1340;
wire n_1771;
wire n_631;
wire n_720;
wire n_842;
wire n_1707;
wire n_1432;
wire n_843;
wire n_656;
wire n_989;
wire n_1277;
wire n_797;
wire n_1473;
wire n_1723;
wire n_1246;
wire n_1878;
wire n_899;
wire n_189;
wire n_738;
wire n_1304;
wire n_1035;
wire n_294;
wire n_499;
wire n_1426;
wire n_705;
wire n_1004;
wire n_1176;
wire n_1529;
wire n_1022;
wire n_614;
wire n_529;
wire n_425;
wire n_684;
wire n_1431;
wire n_1615;
wire n_1474;
wire n_1571;
wire n_1809;
wire n_1577;
wire n_1181;
wire n_1822;
wire n_486;
wire n_947;
wire n_1117;
wire n_1087;
wire n_1448;
wire n_648;
wire n_657;
wire n_1049;
wire n_1666;
wire n_1505;
wire n_803;
wire n_290;
wire n_1717;
wire n_926;
wire n_1817;
wire n_927;
wire n_1849;
wire n_919;
wire n_1698;
wire n_478;
wire n_929;
wire n_1228;
wire n_417;
wire n_446;
wire n_1568;
wire n_1490;
wire n_777;
wire n_1299;
wire n_272;
wire n_526;
wire n_1183;
wire n_1436;
wire n_1384;
wire n_293;
wire n_458;
wire n_1070;
wire n_998;
wire n_717;
wire n_1665;
wire n_1383;
wire n_1178;
wire n_1424;
wire n_1073;
wire n_1000;
wire n_796;
wire n_252;
wire n_1195;
wire n_1626;
wire n_1507;
wire n_184;
wire n_552;
wire n_1358;
wire n_1811;
wire n_1388;
wire n_216;
wire n_912;
wire n_1857;
wire n_1519;
wire n_745;
wire n_1284;
wire n_1604;
wire n_1142;
wire n_716;
wire n_1475;
wire n_623;
wire n_1048;
wire n_1201;
wire n_1398;
wire n_884;
wire n_1774;
wire n_1395;
wire n_731;
wire n_1502;
wire n_1659;
wire n_755;
wire n_931;
wire n_1021;
wire n_474;
wire n_683;
wire n_527;
wire n_811;
wire n_1207;
wire n_312;
wire n_1791;
wire n_1368;
wire n_1418;
wire n_958;
wire n_292;
wire n_1250;
wire n_1137;
wire n_1897;
wire n_880;
wire n_889;
wire n_1478;
wire n_589;
wire n_1310;
wire n_819;
wire n_1363;
wire n_1334;
wire n_767;
wire n_1314;
wire n_600;
wire n_964;
wire n_831;
wire n_1837;
wire n_477;
wire n_954;
wire n_864;
wire n_1110;
wire n_1410;
wire n_399;
wire n_1440;
wire n_1382;
wire n_1534;
wire n_1564;
wire n_1736;
wire n_211;
wire n_1483;
wire n_1834;
wire n_1372;
wire n_231;
wire n_1457;
wire n_505;
wire n_1719;
wire n_319;
wire n_1339;
wire n_1787;
wire n_537;
wire n_1427;
wire n_311;
wire n_1466;
wire n_403;
wire n_1080;
wire n_723;
wire n_1877;
wire n_596;
wire n_546;
wire n_562;
wire n_1141;
wire n_1268;
wire n_386;
wire n_1769;
wire n_1220;
wire n_1893;
wire n_556;
wire n_1755;
wire n_1602;
wire n_1136;
wire n_1125;
wire n_970;
wire n_642;
wire n_995;
wire n_276;
wire n_1159;
wire n_1092;
wire n_441;
wire n_221;
wire n_1060;
wire n_444;
wire n_1252;
wire n_1784;
wire n_1223;
wire n_303;
wire n_511;
wire n_193;
wire n_1286;
wire n_1773;
wire n_1775;
wire n_1053;
wire n_416;
wire n_1681;
wire n_520;
wire n_418;
wire n_1093;
wire n_1783;
wire n_1533;
wire n_1597;
wire n_266;
wire n_296;
wire n_775;
wire n_651;
wire n_1153;
wire n_439;
wire n_1618;
wire n_217;
wire n_518;
wire n_1531;
wire n_1185;
wire n_453;
wire n_215;
wire n_1745;
wire n_914;
wire n_759;
wire n_1831;
wire n_426;
wire n_317;
wire n_1653;
wire n_1679;
wire n_1625;
wire n_1453;
wire n_488;
wire n_497;
wire n_773;
wire n_1901;
wire n_920;
wire n_1374;
wire n_1315;
wire n_1647;
wire n_1224;
wire n_1614;
wire n_1459;
wire n_1892;
wire n_1135;
wire n_1179;
wire n_1169;
wire n_401;
wire n_324;
wire n_1617;
wire n_335;
wire n_1470;
wire n_463;
wire n_1243;
wire n_848;
wire n_301;
wire n_274;
wire n_1096;
wire n_1091;
wire n_1580;
wire n_1425;
wire n_1881;
wire n_1281;
wire n_1267;
wire n_1806;
wire n_983;
wire n_427;
wire n_1520;
wire n_496;
wire n_906;
wire n_1390;
wire n_688;
wire n_1077;
wire n_1733;
wire n_1419;
wire n_351;
wire n_259;
wire n_1731;
wire n_177;
wire n_1855;
wire n_1636;
wire n_1437;
wire n_1645;
wire n_1832;
wire n_385;
wire n_1687;
wire n_1439;
wire n_1323;
wire n_858;
wire n_1331;
wire n_613;
wire n_736;
wire n_501;
wire n_956;
wire n_960;
wire n_663;
wire n_856;
wire n_379;
wire n_778;
wire n_1668;
wire n_1134;
wire n_410;
wire n_1129;
wire n_554;
wire n_602;
wire n_1696;
wire n_1594;
wire n_664;
wire n_1869;
wire n_1764;
wire n_1429;
wire n_1610;
wire n_1889;
wire n_435;
wire n_1905;
wire n_793;
wire n_326;
wire n_587;
wire n_1593;
wire n_580;
wire n_762;
wire n_1030;
wire n_1202;
wire n_465;
wire n_1790;
wire n_1778;
wire n_1635;
wire n_1079;
wire n_341;
wire n_1744;
wire n_828;
wire n_607;
wire n_316;
wire n_419;
wire n_1551;
wire n_1103;
wire n_1203;
wire n_820;
wire n_951;
wire n_725;
wire n_952;
wire n_999;
wire n_358;
wire n_1254;
wire n_186;
wire n_368;
wire n_575;
wire n_994;
wire n_1508;
wire n_732;
wire n_974;
wire n_392;
wire n_724;
wire n_1020;
wire n_1042;
wire n_628;
wire n_1273;
wire n_1434;
wire n_1573;
wire n_1728;
wire n_557;
wire n_1871;
wire n_349;
wire n_617;
wire n_845;
wire n_807;
wire n_1036;
wire n_1138;
wire n_1661;
wire n_1275;
wire n_485;
wire n_1549;
wire n_443;
wire n_1510;
wire n_892;
wire n_768;
wire n_421;
wire n_1468;
wire n_1859;
wire n_238;
wire n_1095;
wire n_1595;
wire n_202;
wire n_1718;
wire n_1749;
wire n_1683;
wire n_597;
wire n_280;
wire n_1270;
wire n_1187;
wire n_610;
wire n_1403;
wire n_1669;
wire n_1852;
wire n_1024;
wire n_1768;
wire n_198;
wire n_1847;
wire n_179;
wire n_248;
wire n_517;
wire n_1667;
wire n_667;
wire n_1206;
wire n_621;
wire n_1037;
wire n_1397;
wire n_1279;
wire n_1115;
wire n_750;
wire n_901;
wire n_1499;
wire n_468;
wire n_923;
wire n_504;
wire n_1409;
wire n_1841;
wire n_1639;
wire n_1623;
wire n_183;
wire n_1015;
wire n_1503;
wire n_466;
wire n_1057;
wire n_603;
wire n_991;
wire n_1657;
wire n_235;
wire n_1126;
wire n_340;
wire n_710;
wire n_1108;
wire n_1818;
wire n_1182;
wire n_1298;
wire n_1611;
wire n_785;
wire n_746;
wire n_609;
wire n_1601;
wire n_1686;
wire n_1356;
wire n_1589;
wire n_1740;
wire n_1497;
wire n_1168;
wire n_1216;
wire n_1320;
wire n_1430;
wire n_1316;
wire n_1287;
wire n_1452;
wire n_1622;
wire n_1586;
wire n_302;
wire n_1694;
wire n_380;
wire n_1535;
wire n_1596;
wire n_1190;
wire n_1734;
wire n_397;
wire n_1262;
wire n_218;
wire n_1891;
wire n_1213;
wire n_1350;
wire n_1673;
wire n_1715;
wire n_1443;
wire n_1272;
wire n_239;
wire n_782;
wire n_1539;
wire n_490;
wire n_220;
wire n_809;
wire n_1043;
wire n_1797;
wire n_1608;
wire n_986;
wire n_1472;
wire n_1081;
wire n_402;
wire n_1870;
wire n_352;
wire n_1692;
wire n_800;
wire n_1084;
wire n_1171;
wire n_460;
wire n_1827;
wire n_1361;
wire n_1864;
wire n_1491;
wire n_662;
wire n_374;
wire n_1152;
wire n_1840;
wire n_1705;
wire n_450;
wire n_1684;
wire n_921;
wire n_1346;
wire n_711;
wire n_1642;
wire n_579;
wire n_1352;
wire n_937;
wire n_1682;
wire n_370;
wire n_1695;
wire n_1828;
wire n_650;
wire n_1046;
wire n_1145;
wire n_330;
wire n_1121;
wire n_1102;
wire n_972;
wire n_1405;
wire n_258;
wire n_1406;
wire n_456;
wire n_1332;
wire n_260;
wire n_313;
wire n_624;
wire n_962;
wire n_1041;
wire n_565;
wire n_356;
wire n_1569;
wire n_936;
wire n_1883;
wire n_1288;
wire n_1186;
wire n_1062;
wire n_885;
wire n_896;
wire n_654;
wire n_411;
wire n_1222;
wire n_599;
wire n_776;
wire n_321;
wire n_1823;
wire n_227;
wire n_1720;
wire n_204;
wire n_482;
wire n_934;
wire n_1637;
wire n_1407;
wire n_1795;
wire n_420;
wire n_1341;
wire n_394;
wire n_1456;
wire n_1845;
wire n_1489;
wire n_942;
wire n_1524;
wire n_543;
wire n_1496;
wire n_1271;
wire n_1545;
wire n_1355;
wire n_1225;
wire n_1544;
wire n_1485;
wire n_325;
wire n_1640;
wire n_804;
wire n_464;
wire n_1846;
wire n_533;
wire n_806;
wire n_959;
wire n_879;
wire n_584;
wire n_244;
wire n_1343;
wire n_1522;
wire n_548;
wire n_1782;
wire n_282;
wire n_1676;
wire n_833;
wire n_1830;
wire n_1567;
wire n_523;
wire n_1319;
wire n_707;
wire n_345;
wire n_1900;
wire n_799;
wire n_1548;
wire n_1155;
wire n_273;
wire n_1633;
wire n_787;
wire n_1416;
wire n_1528;
wire n_1146;
wire n_1086;
wire n_1066;
wire n_1282;
wire n_550;
wire n_275;
wire n_652;
wire n_560;
wire n_1906;
wire n_1484;
wire n_1321;
wire n_1241;
wire n_1672;
wire n_569;
wire n_1758;
wire n_737;
wire n_1318;
wire n_1235;
wire n_1229;
wire n_306;
wire n_1292;
wire n_1373;
wire n_346;
wire n_1029;
wire n_1447;
wire n_790;
wire n_1706;
wire n_1498;
wire n_1210;
wire n_299;
wire n_1248;
wire n_1556;
wire n_902;
wire n_333;
wire n_1047;
wire n_1385;
wire n_431;
wire n_459;
wire n_1269;
wire n_502;
wire n_672;
wire n_1257;
wire n_1751;
wire n_285;
wire n_1375;
wire n_655;
wire n_706;
wire n_1045;
wire n_1650;
wire n_786;
wire n_1794;
wire n_1236;
wire n_1559;
wire n_1725;
wire n_1872;
wire n_834;
wire n_743;
wire n_766;
wire n_430;
wire n_1746;
wire n_1325;
wire n_1002;
wire n_1741;
wire n_545;
wire n_489;
wire n_1804;
wire n_1727;
wire n_251;
wire n_1019;
wire n_636;
wire n_729;
wire n_876;
wire n_774;
wire n_1337;
wire n_660;
wire n_438;
wire n_1477;
wire n_1360;
wire n_1860;
wire n_1904;
wire n_1200;
wire n_479;
wire n_1607;
wire n_1353;
wire n_1777;
wire n_1908;
wire n_1454;
wire n_869;
wire n_1154;
wire n_1113;
wire n_1600;
wire n_646;
wire n_528;
wire n_391;
wire n_1098;
wire n_1329;
wire n_817;
wire n_262;
wire n_187;
wire n_897;
wire n_846;
wire n_841;
wire n_1476;
wire n_1001;
wire n_508;
wire n_1800;
wire n_1050;
wire n_1411;
wire n_1463;
wire n_1177;
wire n_332;
wire n_1150;
wire n_1742;
wire n_1562;
wire n_1690;
wire n_398;
wire n_1191;
wire n_1826;
wire n_566;
wire n_1023;
wire n_1882;
wire n_1076;
wire n_1118;
wire n_194;
wire n_1007;
wire n_1807;
wire n_1378;
wire n_855;
wire n_1592;
wire n_1759;
wire n_1814;
wire n_1631;
wire n_591;
wire n_1377;
wire n_1879;
wire n_256;
wire n_853;
wire n_440;
wire n_695;
wire n_1542;
wire n_875;
wire n_209;
wire n_367;
wire n_680;
wire n_1678;
wire n_661;
wire n_1716;
wire n_278;
wire n_1256;
wire n_671;
wire n_933;
wire n_740;
wire n_703;
wire n_978;
wire n_384;
wire n_1291;
wire n_1217;
wire n_751;
wire n_749;
wire n_1824;
wire n_310;
wire n_1628;
wire n_1324;
wire n_1399;
wire n_1435;
wire n_969;
wire n_988;
wire n_1065;
wire n_1401;
wire n_1255;
wire n_568;
wire n_1516;
wire n_1536;
wire n_180;
wire n_1204;
wire n_823;
wire n_1132;
wire n_643;
wire n_233;
wire n_698;
wire n_1074;
wire n_1394;
wire n_1327;
wire n_1326;
wire n_739;
wire n_400;
wire n_955;
wire n_337;
wire n_1379;
wire n_214;
wire n_246;
wire n_1338;
wire n_1097;
wire n_935;
wire n_781;
wire n_789;
wire n_1554;
wire n_1130;
wire n_181;
wire n_1810;
wire n_182;
wire n_573;
wire n_769;
wire n_676;
wire n_327;
wire n_1120;
wire n_832;
wire n_1583;
wire n_1730;
wire n_555;
wire n_389;
wire n_814;
wire n_1643;
wire n_1729;
wire n_669;
wire n_300;
wire n_222;
wire n_747;
wire n_1389;
wire n_1105;
wire n_721;
wire n_1461;
wire n_742;
wire n_535;
wire n_691;
wire n_372;
wire n_314;
wire n_1408;
wire n_378;
wire n_1196;
wire n_377;
wire n_1598;
wire n_863;
wire n_601;
wire n_338;
wire n_1283;
wire n_918;
wire n_748;
wire n_506;
wire n_1114;
wire n_1785;
wire n_763;
wire n_1147;
wire n_1848;
wire n_360;
wire n_1754;
wire n_1506;
wire n_1652;
wire n_1812;
wire n_957;
wire n_895;
wire n_866;
wire n_1227;
wire n_191;
wire n_387;
wire n_452;
wire n_744;
wire n_971;
wire n_946;
wire n_344;
wire n_761;
wire n_1303;
wire n_1205;
wire n_1258;
wire n_1392;
wire n_1173;
wire n_525;
wire n_1677;
wire n_1116;
wire n_611;
wire n_1702;
wire n_1570;
wire n_1219;
wire n_1780;
wire n_1689;
wire n_1174;
wire n_1016;
wire n_1347;
wire n_795;
wire n_1501;
wire n_1221;
wire n_1245;
wire n_838;
wire n_647;
wire n_197;
wire n_844;
wire n_448;
wire n_1017;
wire n_1083;
wire n_445;
wire n_1561;
wire n_930;
wire n_888;
wire n_1112;
wire n_234;
wire n_910;
wire n_1656;
wire n_1721;
wire n_1460;
wire n_911;
wire n_1464;
wire n_236;
wire n_653;
wire n_1737;
wire n_1414;
wire n_752;
wire n_908;
wire n_944;
wire n_576;
wire n_1028;
wire n_472;
wire n_270;
wire n_414;
wire n_563;
wire n_1011;
wire n_1566;
wire n_1215;
wire n_839;
wire n_708;
wire n_668;
wire n_626;
wire n_990;
wire n_1500;
wire n_779;
wire n_1537;
wire n_1821;
wire n_1104;
wire n_854;
wire n_1058;
wire n_498;
wire n_1122;
wire n_870;
wire n_904;
wire n_1253;
wire n_709;
wire n_1266;
wire n_366;
wire n_1509;
wire n_1693;
wire n_1109;
wire n_185;
wire n_712;
wire n_348;
wire n_1276;
wire n_376;
wire n_390;
wire n_1148;
wire n_334;
wire n_1161;
wire n_1085;
wire n_232;
wire n_1239;
wire n_771;
wire n_1584;
wire n_470;
wire n_475;
wire n_924;
wire n_298;
wire n_1582;
wire n_492;
wire n_1149;
wire n_265;
wire n_1184;
wire n_228;
wire n_719;
wire n_1525;
wire n_455;
wire n_1585;
wire n_1851;
wire n_363;
wire n_1799;
wire n_1090;
wire n_592;
wire n_1816;
wire n_1518;
wire n_829;
wire n_1156;
wire n_1362;
wire n_393;
wire n_984;
wire n_1829;
wire n_503;
wire n_1450;
wire n_1638;
wire n_868;
wire n_570;
wire n_859;
wire n_406;
wire n_735;
wire n_1789;
wire n_1770;
wire n_878;
wire n_620;
wire n_519;
wire n_307;
wire n_469;
wire n_1218;
wire n_500;
wire n_1482;
wire n_981;
wire n_714;
wire n_1349;
wire n_291;
wire n_1144;
wire n_357;
wire n_985;
wire n_481;
wire n_997;
wire n_1710;
wire n_1301;
wire n_802;
wire n_561;
wire n_980;
wire n_1306;
wire n_1651;
wire n_1198;
wire n_1609;
wire n_436;
wire n_409;
wire n_1244;
wire n_1685;
wire n_1763;
wire n_1574;
wire n_240;
wire n_756;
wire n_1619;
wire n_1606;
wire n_810;
wire n_1133;
wire n_635;
wire n_1194;
wire n_1051;
wire n_253;
wire n_1552;
wire n_583;
wire n_249;
wire n_201;
wire n_1039;
wire n_1442;
wire n_1034;
wire n_1480;
wire n_1158;
wire n_754;
wire n_941;
wire n_975;
wire n_1031;
wire n_1305;
wire n_553;
wire n_849;
wire n_753;
wire n_1753;
wire n_467;
wire n_269;
wire n_359;
wire n_973;
wire n_1479;
wire n_1055;
wire n_1675;
wire n_582;
wire n_861;
wire n_857;
wire n_967;
wire n_571;
wire n_404;
wire n_271;
wire n_1884;
wire n_206;
wire n_679;
wire n_633;
wire n_1170;
wire n_665;
wire n_1629;
wire n_588;
wire n_225;
wire n_1260;
wire n_308;
wire n_309;
wire n_1819;
wire n_1010;
wire n_1040;
wire n_915;
wire n_632;
wire n_1166;
wire n_812;
wire n_1131;
wire n_1761;
wire n_534;
wire n_1578;
wire n_1006;
wire n_1861;
wire n_373;
wire n_1632;
wire n_1890;
wire n_1805;
wire n_257;
wire n_1557;
wire n_1888;
wire n_1833;
wire n_730;
wire n_1311;
wire n_1494;
wire n_670;
wire n_203;
wire n_1850;
wire n_1898;
wire n_1868;
wire n_207;
wire n_1089;
wire n_1887;
wire n_1587;
wire n_1365;
wire n_1417;
wire n_205;
wire n_1242;
wire n_1836;
wire n_681;
wire n_1226;
wire n_1274;
wire n_1486;
wire n_412;
wire n_640;
wire n_1322;
wire n_965;
wire n_1899;
wire n_1428;
wire n_1616;
wire n_1576;
wire n_1856;
wire n_1862;
wire n_339;
wire n_784;
wire n_434;
wire n_315;
wire n_288;
wire n_1059;
wire n_1197;
wire n_422;
wire n_722;
wire n_862;
wire n_540;
wire n_1423;
wire n_457;
wire n_364;
wire n_629;
wire n_1621;
wire n_1748;
wire n_900;
wire n_1449;
wire n_531;
wire n_827;
wire n_361;
wire n_1025;
wire n_336;
wire n_1885;
wire n_1013;
wire n_1259;
wire n_192;
wire n_1538;
wire n_649;
wire n_1612;
wire n_1240;

INVx2_ASAP7_75t_L g177 ( 
.A(n_73),
.Y(n_177)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_121),
.Y(n_178)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_94),
.Y(n_179)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_123),
.Y(n_180)
);

BUFx2_ASAP7_75t_L g181 ( 
.A(n_14),
.Y(n_181)
);

CKINVDCx5p33_ASAP7_75t_R g182 ( 
.A(n_21),
.Y(n_182)
);

CKINVDCx5p33_ASAP7_75t_R g183 ( 
.A(n_162),
.Y(n_183)
);

CKINVDCx5p33_ASAP7_75t_R g184 ( 
.A(n_44),
.Y(n_184)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_90),
.Y(n_185)
);

CKINVDCx5p33_ASAP7_75t_R g186 ( 
.A(n_127),
.Y(n_186)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_49),
.Y(n_187)
);

CKINVDCx5p33_ASAP7_75t_R g188 ( 
.A(n_18),
.Y(n_188)
);

CKINVDCx5p33_ASAP7_75t_R g189 ( 
.A(n_19),
.Y(n_189)
);

CKINVDCx5p33_ASAP7_75t_R g190 ( 
.A(n_125),
.Y(n_190)
);

CKINVDCx5p33_ASAP7_75t_R g191 ( 
.A(n_21),
.Y(n_191)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_145),
.Y(n_192)
);

CKINVDCx5p33_ASAP7_75t_R g193 ( 
.A(n_157),
.Y(n_193)
);

CKINVDCx5p33_ASAP7_75t_R g194 ( 
.A(n_141),
.Y(n_194)
);

CKINVDCx20_ASAP7_75t_R g195 ( 
.A(n_31),
.Y(n_195)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_142),
.Y(n_196)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_55),
.Y(n_197)
);

CKINVDCx5p33_ASAP7_75t_R g198 ( 
.A(n_130),
.Y(n_198)
);

HB1xp67_ASAP7_75t_L g199 ( 
.A(n_92),
.Y(n_199)
);

CKINVDCx5p33_ASAP7_75t_R g200 ( 
.A(n_33),
.Y(n_200)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_132),
.Y(n_201)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_65),
.Y(n_202)
);

CKINVDCx14_ASAP7_75t_R g203 ( 
.A(n_107),
.Y(n_203)
);

CKINVDCx5p33_ASAP7_75t_R g204 ( 
.A(n_64),
.Y(n_204)
);

CKINVDCx20_ASAP7_75t_R g205 ( 
.A(n_15),
.Y(n_205)
);

CKINVDCx5p33_ASAP7_75t_R g206 ( 
.A(n_75),
.Y(n_206)
);

CKINVDCx5p33_ASAP7_75t_R g207 ( 
.A(n_67),
.Y(n_207)
);

INVx1_ASAP7_75t_SL g208 ( 
.A(n_151),
.Y(n_208)
);

CKINVDCx5p33_ASAP7_75t_R g209 ( 
.A(n_61),
.Y(n_209)
);

BUFx6f_ASAP7_75t_L g210 ( 
.A(n_126),
.Y(n_210)
);

CKINVDCx5p33_ASAP7_75t_R g211 ( 
.A(n_39),
.Y(n_211)
);

CKINVDCx20_ASAP7_75t_R g212 ( 
.A(n_91),
.Y(n_212)
);

CKINVDCx5p33_ASAP7_75t_R g213 ( 
.A(n_0),
.Y(n_213)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_80),
.Y(n_214)
);

CKINVDCx20_ASAP7_75t_R g215 ( 
.A(n_10),
.Y(n_215)
);

CKINVDCx5p33_ASAP7_75t_R g216 ( 
.A(n_77),
.Y(n_216)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_38),
.Y(n_217)
);

CKINVDCx5p33_ASAP7_75t_R g218 ( 
.A(n_116),
.Y(n_218)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_39),
.Y(n_219)
);

CKINVDCx20_ASAP7_75t_R g220 ( 
.A(n_117),
.Y(n_220)
);

INVx1_ASAP7_75t_SL g221 ( 
.A(n_9),
.Y(n_221)
);

CKINVDCx5p33_ASAP7_75t_R g222 ( 
.A(n_138),
.Y(n_222)
);

CKINVDCx5p33_ASAP7_75t_R g223 ( 
.A(n_26),
.Y(n_223)
);

CKINVDCx5p33_ASAP7_75t_R g224 ( 
.A(n_143),
.Y(n_224)
);

CKINVDCx5p33_ASAP7_75t_R g225 ( 
.A(n_83),
.Y(n_225)
);

CKINVDCx5p33_ASAP7_75t_R g226 ( 
.A(n_86),
.Y(n_226)
);

CKINVDCx5p33_ASAP7_75t_R g227 ( 
.A(n_152),
.Y(n_227)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_59),
.Y(n_228)
);

CKINVDCx5p33_ASAP7_75t_R g229 ( 
.A(n_109),
.Y(n_229)
);

CKINVDCx5p33_ASAP7_75t_R g230 ( 
.A(n_164),
.Y(n_230)
);

CKINVDCx5p33_ASAP7_75t_R g231 ( 
.A(n_78),
.Y(n_231)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_166),
.Y(n_232)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_52),
.Y(n_233)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_135),
.Y(n_234)
);

BUFx10_ASAP7_75t_L g235 ( 
.A(n_170),
.Y(n_235)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_108),
.Y(n_236)
);

CKINVDCx5p33_ASAP7_75t_R g237 ( 
.A(n_71),
.Y(n_237)
);

INVxp67_ASAP7_75t_L g238 ( 
.A(n_31),
.Y(n_238)
);

CKINVDCx5p33_ASAP7_75t_R g239 ( 
.A(n_24),
.Y(n_239)
);

CKINVDCx5p33_ASAP7_75t_R g240 ( 
.A(n_167),
.Y(n_240)
);

CKINVDCx5p33_ASAP7_75t_R g241 ( 
.A(n_44),
.Y(n_241)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_136),
.Y(n_242)
);

BUFx6f_ASAP7_75t_L g243 ( 
.A(n_76),
.Y(n_243)
);

CKINVDCx5p33_ASAP7_75t_R g244 ( 
.A(n_124),
.Y(n_244)
);

CKINVDCx20_ASAP7_75t_R g245 ( 
.A(n_22),
.Y(n_245)
);

CKINVDCx5p33_ASAP7_75t_R g246 ( 
.A(n_59),
.Y(n_246)
);

BUFx10_ASAP7_75t_L g247 ( 
.A(n_100),
.Y(n_247)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_23),
.Y(n_248)
);

HB1xp67_ASAP7_75t_L g249 ( 
.A(n_58),
.Y(n_249)
);

BUFx3_ASAP7_75t_L g250 ( 
.A(n_99),
.Y(n_250)
);

CKINVDCx5p33_ASAP7_75t_R g251 ( 
.A(n_171),
.Y(n_251)
);

CKINVDCx5p33_ASAP7_75t_R g252 ( 
.A(n_95),
.Y(n_252)
);

BUFx3_ASAP7_75t_L g253 ( 
.A(n_63),
.Y(n_253)
);

BUFx3_ASAP7_75t_L g254 ( 
.A(n_98),
.Y(n_254)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_133),
.Y(n_255)
);

CKINVDCx5p33_ASAP7_75t_R g256 ( 
.A(n_104),
.Y(n_256)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_40),
.Y(n_257)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_175),
.Y(n_258)
);

CKINVDCx5p33_ASAP7_75t_R g259 ( 
.A(n_96),
.Y(n_259)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_69),
.Y(n_260)
);

CKINVDCx5p33_ASAP7_75t_R g261 ( 
.A(n_103),
.Y(n_261)
);

INVxp67_ASAP7_75t_L g262 ( 
.A(n_49),
.Y(n_262)
);

CKINVDCx5p33_ASAP7_75t_R g263 ( 
.A(n_154),
.Y(n_263)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_160),
.Y(n_264)
);

CKINVDCx5p33_ASAP7_75t_R g265 ( 
.A(n_150),
.Y(n_265)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_4),
.Y(n_266)
);

CKINVDCx5p33_ASAP7_75t_R g267 ( 
.A(n_66),
.Y(n_267)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_56),
.Y(n_268)
);

CKINVDCx5p33_ASAP7_75t_R g269 ( 
.A(n_33),
.Y(n_269)
);

BUFx10_ASAP7_75t_L g270 ( 
.A(n_32),
.Y(n_270)
);

BUFx6f_ASAP7_75t_L g271 ( 
.A(n_137),
.Y(n_271)
);

INVx1_ASAP7_75t_SL g272 ( 
.A(n_176),
.Y(n_272)
);

CKINVDCx5p33_ASAP7_75t_R g273 ( 
.A(n_12),
.Y(n_273)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_35),
.Y(n_274)
);

BUFx3_ASAP7_75t_L g275 ( 
.A(n_29),
.Y(n_275)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_82),
.Y(n_276)
);

CKINVDCx5p33_ASAP7_75t_R g277 ( 
.A(n_23),
.Y(n_277)
);

CKINVDCx20_ASAP7_75t_R g278 ( 
.A(n_155),
.Y(n_278)
);

CKINVDCx5p33_ASAP7_75t_R g279 ( 
.A(n_140),
.Y(n_279)
);

INVx2_ASAP7_75t_SL g280 ( 
.A(n_11),
.Y(n_280)
);

BUFx10_ASAP7_75t_L g281 ( 
.A(n_113),
.Y(n_281)
);

CKINVDCx5p33_ASAP7_75t_R g282 ( 
.A(n_84),
.Y(n_282)
);

CKINVDCx5p33_ASAP7_75t_R g283 ( 
.A(n_16),
.Y(n_283)
);

CKINVDCx5p33_ASAP7_75t_R g284 ( 
.A(n_70),
.Y(n_284)
);

BUFx3_ASAP7_75t_L g285 ( 
.A(n_36),
.Y(n_285)
);

CKINVDCx5p33_ASAP7_75t_R g286 ( 
.A(n_56),
.Y(n_286)
);

INVx1_ASAP7_75t_SL g287 ( 
.A(n_102),
.Y(n_287)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_14),
.Y(n_288)
);

CKINVDCx5p33_ASAP7_75t_R g289 ( 
.A(n_40),
.Y(n_289)
);

BUFx2_ASAP7_75t_R g290 ( 
.A(n_146),
.Y(n_290)
);

BUFx2_ASAP7_75t_SL g291 ( 
.A(n_30),
.Y(n_291)
);

CKINVDCx5p33_ASAP7_75t_R g292 ( 
.A(n_89),
.Y(n_292)
);

INVx2_ASAP7_75t_L g293 ( 
.A(n_147),
.Y(n_293)
);

CKINVDCx20_ASAP7_75t_R g294 ( 
.A(n_52),
.Y(n_294)
);

CKINVDCx5p33_ASAP7_75t_R g295 ( 
.A(n_22),
.Y(n_295)
);

INVxp67_ASAP7_75t_SL g296 ( 
.A(n_38),
.Y(n_296)
);

CKINVDCx5p33_ASAP7_75t_R g297 ( 
.A(n_97),
.Y(n_297)
);

CKINVDCx5p33_ASAP7_75t_R g298 ( 
.A(n_101),
.Y(n_298)
);

INVx1_ASAP7_75t_SL g299 ( 
.A(n_149),
.Y(n_299)
);

INVx1_ASAP7_75t_SL g300 ( 
.A(n_159),
.Y(n_300)
);

INVx1_ASAP7_75t_SL g301 ( 
.A(n_122),
.Y(n_301)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_74),
.Y(n_302)
);

INVxp67_ASAP7_75t_L g303 ( 
.A(n_60),
.Y(n_303)
);

CKINVDCx5p33_ASAP7_75t_R g304 ( 
.A(n_62),
.Y(n_304)
);

BUFx8_ASAP7_75t_SL g305 ( 
.A(n_13),
.Y(n_305)
);

CKINVDCx5p33_ASAP7_75t_R g306 ( 
.A(n_88),
.Y(n_306)
);

CKINVDCx5p33_ASAP7_75t_R g307 ( 
.A(n_106),
.Y(n_307)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_17),
.Y(n_308)
);

CKINVDCx5p33_ASAP7_75t_R g309 ( 
.A(n_87),
.Y(n_309)
);

BUFx3_ASAP7_75t_L g310 ( 
.A(n_156),
.Y(n_310)
);

BUFx3_ASAP7_75t_L g311 ( 
.A(n_12),
.Y(n_311)
);

CKINVDCx5p33_ASAP7_75t_R g312 ( 
.A(n_118),
.Y(n_312)
);

INVx1_ASAP7_75t_SL g313 ( 
.A(n_48),
.Y(n_313)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_41),
.Y(n_314)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_153),
.Y(n_315)
);

CKINVDCx20_ASAP7_75t_R g316 ( 
.A(n_62),
.Y(n_316)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_18),
.Y(n_317)
);

CKINVDCx5p33_ASAP7_75t_R g318 ( 
.A(n_45),
.Y(n_318)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_36),
.Y(n_319)
);

CKINVDCx5p33_ASAP7_75t_R g320 ( 
.A(n_15),
.Y(n_320)
);

CKINVDCx20_ASAP7_75t_R g321 ( 
.A(n_172),
.Y(n_321)
);

CKINVDCx5p33_ASAP7_75t_R g322 ( 
.A(n_131),
.Y(n_322)
);

CKINVDCx5p33_ASAP7_75t_R g323 ( 
.A(n_8),
.Y(n_323)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_19),
.Y(n_324)
);

INVx2_ASAP7_75t_L g325 ( 
.A(n_120),
.Y(n_325)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_29),
.Y(n_326)
);

CKINVDCx5p33_ASAP7_75t_R g327 ( 
.A(n_105),
.Y(n_327)
);

BUFx3_ASAP7_75t_L g328 ( 
.A(n_7),
.Y(n_328)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_148),
.Y(n_329)
);

CKINVDCx5p33_ASAP7_75t_R g330 ( 
.A(n_169),
.Y(n_330)
);

CKINVDCx5p33_ASAP7_75t_R g331 ( 
.A(n_119),
.Y(n_331)
);

CKINVDCx5p33_ASAP7_75t_R g332 ( 
.A(n_60),
.Y(n_332)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_111),
.Y(n_333)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_24),
.Y(n_334)
);

INVxp67_ASAP7_75t_L g335 ( 
.A(n_144),
.Y(n_335)
);

CKINVDCx5p33_ASAP7_75t_R g336 ( 
.A(n_32),
.Y(n_336)
);

CKINVDCx5p33_ASAP7_75t_R g337 ( 
.A(n_168),
.Y(n_337)
);

INVx2_ASAP7_75t_SL g338 ( 
.A(n_58),
.Y(n_338)
);

CKINVDCx5p33_ASAP7_75t_R g339 ( 
.A(n_8),
.Y(n_339)
);

CKINVDCx5p33_ASAP7_75t_R g340 ( 
.A(n_85),
.Y(n_340)
);

CKINVDCx5p33_ASAP7_75t_R g341 ( 
.A(n_81),
.Y(n_341)
);

INVx2_ASAP7_75t_L g342 ( 
.A(n_7),
.Y(n_342)
);

CKINVDCx5p33_ASAP7_75t_R g343 ( 
.A(n_5),
.Y(n_343)
);

CKINVDCx5p33_ASAP7_75t_R g344 ( 
.A(n_28),
.Y(n_344)
);

CKINVDCx5p33_ASAP7_75t_R g345 ( 
.A(n_174),
.Y(n_345)
);

CKINVDCx5p33_ASAP7_75t_R g346 ( 
.A(n_112),
.Y(n_346)
);

CKINVDCx20_ASAP7_75t_R g347 ( 
.A(n_42),
.Y(n_347)
);

CKINVDCx5p33_ASAP7_75t_R g348 ( 
.A(n_30),
.Y(n_348)
);

INVx1_ASAP7_75t_L g349 ( 
.A(n_26),
.Y(n_349)
);

BUFx5_ASAP7_75t_L g350 ( 
.A(n_68),
.Y(n_350)
);

INVx2_ASAP7_75t_SL g351 ( 
.A(n_10),
.Y(n_351)
);

CKINVDCx5p33_ASAP7_75t_R g352 ( 
.A(n_50),
.Y(n_352)
);

INVx1_ASAP7_75t_L g353 ( 
.A(n_28),
.Y(n_353)
);

BUFx10_ASAP7_75t_L g354 ( 
.A(n_43),
.Y(n_354)
);

INVx1_ASAP7_75t_L g355 ( 
.A(n_342),
.Y(n_355)
);

NAND2xp5_ASAP7_75t_L g356 ( 
.A(n_280),
.B(n_0),
.Y(n_356)
);

INVx1_ASAP7_75t_L g357 ( 
.A(n_342),
.Y(n_357)
);

INVx1_ASAP7_75t_L g358 ( 
.A(n_275),
.Y(n_358)
);

HB1xp67_ASAP7_75t_L g359 ( 
.A(n_249),
.Y(n_359)
);

HB1xp67_ASAP7_75t_L g360 ( 
.A(n_181),
.Y(n_360)
);

INVxp67_ASAP7_75t_L g361 ( 
.A(n_305),
.Y(n_361)
);

INVx1_ASAP7_75t_L g362 ( 
.A(n_275),
.Y(n_362)
);

INVxp67_ASAP7_75t_L g363 ( 
.A(n_270),
.Y(n_363)
);

INVx1_ASAP7_75t_L g364 ( 
.A(n_285),
.Y(n_364)
);

CKINVDCx5p33_ASAP7_75t_R g365 ( 
.A(n_224),
.Y(n_365)
);

CKINVDCx5p33_ASAP7_75t_R g366 ( 
.A(n_225),
.Y(n_366)
);

INVx1_ASAP7_75t_L g367 ( 
.A(n_285),
.Y(n_367)
);

CKINVDCx14_ASAP7_75t_R g368 ( 
.A(n_203),
.Y(n_368)
);

HB1xp67_ASAP7_75t_L g369 ( 
.A(n_182),
.Y(n_369)
);

CKINVDCx20_ASAP7_75t_R g370 ( 
.A(n_212),
.Y(n_370)
);

INVxp67_ASAP7_75t_SL g371 ( 
.A(n_199),
.Y(n_371)
);

INVxp67_ASAP7_75t_SL g372 ( 
.A(n_250),
.Y(n_372)
);

INVx1_ASAP7_75t_SL g373 ( 
.A(n_221),
.Y(n_373)
);

CKINVDCx20_ASAP7_75t_R g374 ( 
.A(n_220),
.Y(n_374)
);

NOR2xp33_ASAP7_75t_L g375 ( 
.A(n_335),
.B(n_177),
.Y(n_375)
);

CKINVDCx5p33_ASAP7_75t_R g376 ( 
.A(n_226),
.Y(n_376)
);

NAND2xp5_ASAP7_75t_L g377 ( 
.A(n_280),
.B(n_1),
.Y(n_377)
);

CKINVDCx5p33_ASAP7_75t_R g378 ( 
.A(n_227),
.Y(n_378)
);

CKINVDCx20_ASAP7_75t_R g379 ( 
.A(n_278),
.Y(n_379)
);

INVx1_ASAP7_75t_L g380 ( 
.A(n_311),
.Y(n_380)
);

CKINVDCx5p33_ASAP7_75t_R g381 ( 
.A(n_229),
.Y(n_381)
);

INVx1_ASAP7_75t_L g382 ( 
.A(n_311),
.Y(n_382)
);

HB1xp67_ASAP7_75t_L g383 ( 
.A(n_182),
.Y(n_383)
);

CKINVDCx5p33_ASAP7_75t_R g384 ( 
.A(n_230),
.Y(n_384)
);

INVx1_ASAP7_75t_L g385 ( 
.A(n_328),
.Y(n_385)
);

NOR2xp33_ASAP7_75t_L g386 ( 
.A(n_177),
.B(n_1),
.Y(n_386)
);

INVx1_ASAP7_75t_L g387 ( 
.A(n_328),
.Y(n_387)
);

INVx1_ASAP7_75t_L g388 ( 
.A(n_187),
.Y(n_388)
);

INVx1_ASAP7_75t_L g389 ( 
.A(n_197),
.Y(n_389)
);

CKINVDCx5p33_ASAP7_75t_R g390 ( 
.A(n_231),
.Y(n_390)
);

CKINVDCx5p33_ASAP7_75t_R g391 ( 
.A(n_237),
.Y(n_391)
);

NOR2xp33_ASAP7_75t_L g392 ( 
.A(n_293),
.B(n_2),
.Y(n_392)
);

INVx1_ASAP7_75t_L g393 ( 
.A(n_217),
.Y(n_393)
);

INVx1_ASAP7_75t_L g394 ( 
.A(n_219),
.Y(n_394)
);

CKINVDCx5p33_ASAP7_75t_R g395 ( 
.A(n_240),
.Y(n_395)
);

INVx1_ASAP7_75t_L g396 ( 
.A(n_228),
.Y(n_396)
);

CKINVDCx5p33_ASAP7_75t_R g397 ( 
.A(n_244),
.Y(n_397)
);

NOR2xp33_ASAP7_75t_L g398 ( 
.A(n_293),
.B(n_325),
.Y(n_398)
);

CKINVDCx16_ASAP7_75t_R g399 ( 
.A(n_235),
.Y(n_399)
);

NAND2xp5_ASAP7_75t_L g400 ( 
.A(n_338),
.B(n_2),
.Y(n_400)
);

INVx2_ASAP7_75t_L g401 ( 
.A(n_350),
.Y(n_401)
);

CKINVDCx5p33_ASAP7_75t_R g402 ( 
.A(n_251),
.Y(n_402)
);

CKINVDCx5p33_ASAP7_75t_R g403 ( 
.A(n_252),
.Y(n_403)
);

CKINVDCx16_ASAP7_75t_R g404 ( 
.A(n_235),
.Y(n_404)
);

CKINVDCx14_ASAP7_75t_R g405 ( 
.A(n_270),
.Y(n_405)
);

CKINVDCx20_ASAP7_75t_R g406 ( 
.A(n_321),
.Y(n_406)
);

CKINVDCx20_ASAP7_75t_R g407 ( 
.A(n_256),
.Y(n_407)
);

INVx1_ASAP7_75t_L g408 ( 
.A(n_233),
.Y(n_408)
);

INVxp67_ASAP7_75t_SL g409 ( 
.A(n_250),
.Y(n_409)
);

INVx1_ASAP7_75t_L g410 ( 
.A(n_248),
.Y(n_410)
);

CKINVDCx20_ASAP7_75t_R g411 ( 
.A(n_263),
.Y(n_411)
);

NAND2xp5_ASAP7_75t_L g412 ( 
.A(n_338),
.B(n_3),
.Y(n_412)
);

INVx1_ASAP7_75t_L g413 ( 
.A(n_257),
.Y(n_413)
);

CKINVDCx20_ASAP7_75t_R g414 ( 
.A(n_265),
.Y(n_414)
);

NOR2xp33_ASAP7_75t_L g415 ( 
.A(n_325),
.B(n_3),
.Y(n_415)
);

CKINVDCx5p33_ASAP7_75t_R g416 ( 
.A(n_267),
.Y(n_416)
);

CKINVDCx20_ASAP7_75t_R g417 ( 
.A(n_279),
.Y(n_417)
);

CKINVDCx5p33_ASAP7_75t_R g418 ( 
.A(n_322),
.Y(n_418)
);

CKINVDCx5p33_ASAP7_75t_R g419 ( 
.A(n_327),
.Y(n_419)
);

CKINVDCx5p33_ASAP7_75t_R g420 ( 
.A(n_330),
.Y(n_420)
);

CKINVDCx14_ASAP7_75t_R g421 ( 
.A(n_354),
.Y(n_421)
);

NAND2xp5_ASAP7_75t_L g422 ( 
.A(n_351),
.B(n_4),
.Y(n_422)
);

INVx1_ASAP7_75t_L g423 ( 
.A(n_266),
.Y(n_423)
);

INVx1_ASAP7_75t_L g424 ( 
.A(n_268),
.Y(n_424)
);

CKINVDCx5p33_ASAP7_75t_R g425 ( 
.A(n_331),
.Y(n_425)
);

INVx1_ASAP7_75t_L g426 ( 
.A(n_274),
.Y(n_426)
);

CKINVDCx5p33_ASAP7_75t_R g427 ( 
.A(n_337),
.Y(n_427)
);

CKINVDCx5p33_ASAP7_75t_R g428 ( 
.A(n_223),
.Y(n_428)
);

HB1xp67_ASAP7_75t_L g429 ( 
.A(n_184),
.Y(n_429)
);

INVx1_ASAP7_75t_L g430 ( 
.A(n_288),
.Y(n_430)
);

INVx1_ASAP7_75t_L g431 ( 
.A(n_308),
.Y(n_431)
);

INVx1_ASAP7_75t_L g432 ( 
.A(n_314),
.Y(n_432)
);

INVx1_ASAP7_75t_L g433 ( 
.A(n_317),
.Y(n_433)
);

OR2x2_ASAP7_75t_L g434 ( 
.A(n_319),
.B(n_5),
.Y(n_434)
);

INVxp67_ASAP7_75t_SL g435 ( 
.A(n_253),
.Y(n_435)
);

INVx1_ASAP7_75t_L g436 ( 
.A(n_324),
.Y(n_436)
);

CKINVDCx5p33_ASAP7_75t_R g437 ( 
.A(n_241),
.Y(n_437)
);

CKINVDCx20_ASAP7_75t_R g438 ( 
.A(n_183),
.Y(n_438)
);

INVx2_ASAP7_75t_L g439 ( 
.A(n_350),
.Y(n_439)
);

CKINVDCx5p33_ASAP7_75t_R g440 ( 
.A(n_246),
.Y(n_440)
);

CKINVDCx5p33_ASAP7_75t_R g441 ( 
.A(n_269),
.Y(n_441)
);

NAND2xp5_ASAP7_75t_L g442 ( 
.A(n_351),
.B(n_6),
.Y(n_442)
);

CKINVDCx5p33_ASAP7_75t_R g443 ( 
.A(n_273),
.Y(n_443)
);

INVx1_ASAP7_75t_L g444 ( 
.A(n_326),
.Y(n_444)
);

AND2x2_ASAP7_75t_L g445 ( 
.A(n_372),
.B(n_253),
.Y(n_445)
);

INVx1_ASAP7_75t_L g446 ( 
.A(n_388),
.Y(n_446)
);

INVx1_ASAP7_75t_L g447 ( 
.A(n_388),
.Y(n_447)
);

INVx1_ASAP7_75t_L g448 ( 
.A(n_389),
.Y(n_448)
);

NOR2xp33_ASAP7_75t_SL g449 ( 
.A(n_373),
.B(n_290),
.Y(n_449)
);

NAND2xp5_ASAP7_75t_L g450 ( 
.A(n_365),
.B(n_254),
.Y(n_450)
);

OAI21x1_ASAP7_75t_L g451 ( 
.A1(n_401),
.A2(n_439),
.B(n_377),
.Y(n_451)
);

INVx2_ASAP7_75t_L g452 ( 
.A(n_401),
.Y(n_452)
);

AND2x6_ASAP7_75t_L g453 ( 
.A(n_398),
.B(n_210),
.Y(n_453)
);

NOR2xp33_ASAP7_75t_L g454 ( 
.A(n_375),
.B(n_208),
.Y(n_454)
);

AND2x4_ASAP7_75t_L g455 ( 
.A(n_409),
.B(n_254),
.Y(n_455)
);

INVx1_ASAP7_75t_L g456 ( 
.A(n_389),
.Y(n_456)
);

NAND2xp5_ASAP7_75t_SL g457 ( 
.A(n_399),
.B(n_235),
.Y(n_457)
);

HB1xp67_ASAP7_75t_L g458 ( 
.A(n_428),
.Y(n_458)
);

BUFx6f_ASAP7_75t_L g459 ( 
.A(n_401),
.Y(n_459)
);

NOR2xp33_ASAP7_75t_L g460 ( 
.A(n_437),
.B(n_272),
.Y(n_460)
);

BUFx3_ASAP7_75t_L g461 ( 
.A(n_358),
.Y(n_461)
);

BUFx6f_ASAP7_75t_L g462 ( 
.A(n_439),
.Y(n_462)
);

NAND2xp5_ASAP7_75t_L g463 ( 
.A(n_366),
.B(n_310),
.Y(n_463)
);

HB1xp67_ASAP7_75t_L g464 ( 
.A(n_440),
.Y(n_464)
);

INVx5_ASAP7_75t_L g465 ( 
.A(n_439),
.Y(n_465)
);

INVx3_ASAP7_75t_L g466 ( 
.A(n_355),
.Y(n_466)
);

INVx1_ASAP7_75t_L g467 ( 
.A(n_393),
.Y(n_467)
);

BUFx6f_ASAP7_75t_L g468 ( 
.A(n_355),
.Y(n_468)
);

AND2x4_ASAP7_75t_L g469 ( 
.A(n_435),
.B(n_310),
.Y(n_469)
);

INVx1_ASAP7_75t_L g470 ( 
.A(n_393),
.Y(n_470)
);

NAND2xp5_ASAP7_75t_L g471 ( 
.A(n_376),
.B(n_378),
.Y(n_471)
);

INVx1_ASAP7_75t_L g472 ( 
.A(n_394),
.Y(n_472)
);

INVx3_ASAP7_75t_L g473 ( 
.A(n_357),
.Y(n_473)
);

NOR2x1_ASAP7_75t_L g474 ( 
.A(n_386),
.B(n_178),
.Y(n_474)
);

INVxp67_ASAP7_75t_L g475 ( 
.A(n_373),
.Y(n_475)
);

BUFx2_ASAP7_75t_L g476 ( 
.A(n_441),
.Y(n_476)
);

INVx1_ASAP7_75t_L g477 ( 
.A(n_394),
.Y(n_477)
);

NAND2xp5_ASAP7_75t_L g478 ( 
.A(n_381),
.B(n_179),
.Y(n_478)
);

NOR2xp33_ASAP7_75t_SL g479 ( 
.A(n_399),
.B(n_354),
.Y(n_479)
);

INVx1_ASAP7_75t_L g480 ( 
.A(n_396),
.Y(n_480)
);

BUFx2_ASAP7_75t_L g481 ( 
.A(n_443),
.Y(n_481)
);

BUFx6f_ASAP7_75t_L g482 ( 
.A(n_357),
.Y(n_482)
);

AND2x6_ASAP7_75t_L g483 ( 
.A(n_392),
.B(n_210),
.Y(n_483)
);

NAND2xp5_ASAP7_75t_L g484 ( 
.A(n_415),
.B(n_183),
.Y(n_484)
);

BUFx6f_ASAP7_75t_L g485 ( 
.A(n_396),
.Y(n_485)
);

INVx2_ASAP7_75t_L g486 ( 
.A(n_408),
.Y(n_486)
);

INVx1_ASAP7_75t_L g487 ( 
.A(n_408),
.Y(n_487)
);

INVx3_ASAP7_75t_L g488 ( 
.A(n_410),
.Y(n_488)
);

AND2x4_ASAP7_75t_L g489 ( 
.A(n_358),
.B(n_180),
.Y(n_489)
);

NOR2xp33_ASAP7_75t_L g490 ( 
.A(n_384),
.B(n_287),
.Y(n_490)
);

AND2x4_ASAP7_75t_L g491 ( 
.A(n_362),
.B(n_185),
.Y(n_491)
);

NAND2x1p5_ASAP7_75t_L g492 ( 
.A(n_434),
.B(n_299),
.Y(n_492)
);

INVx1_ASAP7_75t_L g493 ( 
.A(n_410),
.Y(n_493)
);

INVx1_ASAP7_75t_L g494 ( 
.A(n_413),
.Y(n_494)
);

NAND2xp5_ASAP7_75t_SL g495 ( 
.A(n_404),
.B(n_247),
.Y(n_495)
);

OA21x2_ASAP7_75t_L g496 ( 
.A1(n_356),
.A2(n_196),
.B(n_192),
.Y(n_496)
);

INVx1_ASAP7_75t_L g497 ( 
.A(n_413),
.Y(n_497)
);

NAND2xp5_ASAP7_75t_L g498 ( 
.A(n_390),
.B(n_201),
.Y(n_498)
);

AND2x4_ASAP7_75t_L g499 ( 
.A(n_362),
.B(n_202),
.Y(n_499)
);

INVx1_ASAP7_75t_L g500 ( 
.A(n_423),
.Y(n_500)
);

INVx2_ASAP7_75t_L g501 ( 
.A(n_423),
.Y(n_501)
);

NOR2xp33_ASAP7_75t_L g502 ( 
.A(n_391),
.B(n_300),
.Y(n_502)
);

INVx1_ASAP7_75t_L g503 ( 
.A(n_424),
.Y(n_503)
);

BUFx3_ASAP7_75t_L g504 ( 
.A(n_364),
.Y(n_504)
);

INVx1_ASAP7_75t_L g505 ( 
.A(n_424),
.Y(n_505)
);

INVx2_ASAP7_75t_L g506 ( 
.A(n_426),
.Y(n_506)
);

NAND2xp5_ASAP7_75t_L g507 ( 
.A(n_395),
.B(n_214),
.Y(n_507)
);

INVx1_ASAP7_75t_L g508 ( 
.A(n_426),
.Y(n_508)
);

INVx1_ASAP7_75t_L g509 ( 
.A(n_430),
.Y(n_509)
);

BUFx6f_ASAP7_75t_L g510 ( 
.A(n_430),
.Y(n_510)
);

AND2x2_ASAP7_75t_SL g511 ( 
.A(n_356),
.B(n_210),
.Y(n_511)
);

INVx2_ASAP7_75t_L g512 ( 
.A(n_431),
.Y(n_512)
);

INVx1_ASAP7_75t_L g513 ( 
.A(n_431),
.Y(n_513)
);

INVx3_ASAP7_75t_L g514 ( 
.A(n_432),
.Y(n_514)
);

BUFx6f_ASAP7_75t_L g515 ( 
.A(n_432),
.Y(n_515)
);

INVx1_ASAP7_75t_L g516 ( 
.A(n_433),
.Y(n_516)
);

INVx2_ASAP7_75t_L g517 ( 
.A(n_433),
.Y(n_517)
);

AND3x2_ASAP7_75t_L g518 ( 
.A(n_360),
.B(n_262),
.C(n_238),
.Y(n_518)
);

INVx1_ASAP7_75t_L g519 ( 
.A(n_436),
.Y(n_519)
);

NAND2xp5_ASAP7_75t_SL g520 ( 
.A(n_404),
.B(n_397),
.Y(n_520)
);

HB1xp67_ASAP7_75t_L g521 ( 
.A(n_405),
.Y(n_521)
);

BUFx6f_ASAP7_75t_L g522 ( 
.A(n_436),
.Y(n_522)
);

INVx1_ASAP7_75t_L g523 ( 
.A(n_485),
.Y(n_523)
);

INVx1_ASAP7_75t_L g524 ( 
.A(n_485),
.Y(n_524)
);

INVx1_ASAP7_75t_L g525 ( 
.A(n_485),
.Y(n_525)
);

INVx4_ASAP7_75t_L g526 ( 
.A(n_459),
.Y(n_526)
);

INVx3_ASAP7_75t_L g527 ( 
.A(n_459),
.Y(n_527)
);

INVx1_ASAP7_75t_L g528 ( 
.A(n_485),
.Y(n_528)
);

INVx2_ASAP7_75t_L g529 ( 
.A(n_452),
.Y(n_529)
);

OAI22xp5_ASAP7_75t_L g530 ( 
.A1(n_492),
.A2(n_371),
.B1(n_417),
.B2(n_407),
.Y(n_530)
);

INVx2_ASAP7_75t_L g531 ( 
.A(n_452),
.Y(n_531)
);

NAND2xp5_ASAP7_75t_L g532 ( 
.A(n_454),
.B(n_402),
.Y(n_532)
);

INVx1_ASAP7_75t_L g533 ( 
.A(n_485),
.Y(n_533)
);

INVx2_ASAP7_75t_L g534 ( 
.A(n_452),
.Y(n_534)
);

INVx2_ASAP7_75t_L g535 ( 
.A(n_468),
.Y(n_535)
);

AOI22xp5_ASAP7_75t_L g536 ( 
.A1(n_460),
.A2(n_414),
.B1(n_411),
.B2(n_438),
.Y(n_536)
);

NAND2xp33_ASAP7_75t_SL g537 ( 
.A(n_457),
.B(n_377),
.Y(n_537)
);

INVx2_ASAP7_75t_L g538 ( 
.A(n_468),
.Y(n_538)
);

OAI22xp33_ASAP7_75t_L g539 ( 
.A1(n_475),
.A2(n_400),
.B1(n_442),
.B2(n_412),
.Y(n_539)
);

BUFx3_ASAP7_75t_L g540 ( 
.A(n_461),
.Y(n_540)
);

INVx1_ASAP7_75t_L g541 ( 
.A(n_485),
.Y(n_541)
);

AND3x2_ASAP7_75t_L g542 ( 
.A(n_479),
.B(n_303),
.C(n_296),
.Y(n_542)
);

OAI22xp5_ASAP7_75t_SL g543 ( 
.A1(n_492),
.A2(n_195),
.B1(n_205),
.B2(n_215),
.Y(n_543)
);

INVx2_ASAP7_75t_L g544 ( 
.A(n_468),
.Y(n_544)
);

INVx1_ASAP7_75t_L g545 ( 
.A(n_510),
.Y(n_545)
);

INVx2_ASAP7_75t_L g546 ( 
.A(n_468),
.Y(n_546)
);

NAND2xp33_ASAP7_75t_L g547 ( 
.A(n_483),
.B(n_453),
.Y(n_547)
);

INVx2_ASAP7_75t_L g548 ( 
.A(n_468),
.Y(n_548)
);

INVx2_ASAP7_75t_L g549 ( 
.A(n_468),
.Y(n_549)
);

AOI22xp33_ASAP7_75t_L g550 ( 
.A1(n_511),
.A2(n_400),
.B1(n_442),
.B2(n_412),
.Y(n_550)
);

INVx2_ASAP7_75t_L g551 ( 
.A(n_482),
.Y(n_551)
);

INVx1_ASAP7_75t_L g552 ( 
.A(n_510),
.Y(n_552)
);

INVx1_ASAP7_75t_L g553 ( 
.A(n_510),
.Y(n_553)
);

INVx6_ASAP7_75t_L g554 ( 
.A(n_489),
.Y(n_554)
);

INVx1_ASAP7_75t_L g555 ( 
.A(n_510),
.Y(n_555)
);

INVx3_ASAP7_75t_L g556 ( 
.A(n_459),
.Y(n_556)
);

INVx3_ASAP7_75t_L g557 ( 
.A(n_459),
.Y(n_557)
);

NAND2xp5_ASAP7_75t_L g558 ( 
.A(n_490),
.B(n_403),
.Y(n_558)
);

INVx2_ASAP7_75t_L g559 ( 
.A(n_482),
.Y(n_559)
);

CKINVDCx20_ASAP7_75t_R g560 ( 
.A(n_476),
.Y(n_560)
);

INVx1_ASAP7_75t_L g561 ( 
.A(n_510),
.Y(n_561)
);

NOR2xp33_ASAP7_75t_L g562 ( 
.A(n_502),
.B(n_416),
.Y(n_562)
);

NAND2xp5_ASAP7_75t_SL g563 ( 
.A(n_479),
.B(n_418),
.Y(n_563)
);

NAND2xp5_ASAP7_75t_L g564 ( 
.A(n_455),
.B(n_419),
.Y(n_564)
);

INVx1_ASAP7_75t_L g565 ( 
.A(n_510),
.Y(n_565)
);

OR2x2_ASAP7_75t_L g566 ( 
.A(n_492),
.B(n_369),
.Y(n_566)
);

OAI22xp33_ASAP7_75t_L g567 ( 
.A1(n_484),
.A2(n_422),
.B1(n_313),
.B2(n_434),
.Y(n_567)
);

NAND2xp5_ASAP7_75t_L g568 ( 
.A(n_455),
.B(n_469),
.Y(n_568)
);

INVx1_ASAP7_75t_L g569 ( 
.A(n_515),
.Y(n_569)
);

NAND2xp5_ASAP7_75t_SL g570 ( 
.A(n_450),
.B(n_420),
.Y(n_570)
);

NOR2xp33_ASAP7_75t_L g571 ( 
.A(n_463),
.B(n_425),
.Y(n_571)
);

INVx1_ASAP7_75t_L g572 ( 
.A(n_515),
.Y(n_572)
);

AOI22xp33_ASAP7_75t_L g573 ( 
.A1(n_511),
.A2(n_422),
.B1(n_359),
.B2(n_353),
.Y(n_573)
);

NAND2xp5_ASAP7_75t_L g574 ( 
.A(n_455),
.B(n_427),
.Y(n_574)
);

INVx2_ASAP7_75t_L g575 ( 
.A(n_482),
.Y(n_575)
);

INVx1_ASAP7_75t_L g576 ( 
.A(n_515),
.Y(n_576)
);

CKINVDCx20_ASAP7_75t_R g577 ( 
.A(n_476),
.Y(n_577)
);

NAND3xp33_ASAP7_75t_L g578 ( 
.A(n_474),
.B(n_429),
.C(n_383),
.Y(n_578)
);

AND2x6_ASAP7_75t_L g579 ( 
.A(n_474),
.B(n_210),
.Y(n_579)
);

NAND2xp5_ASAP7_75t_L g580 ( 
.A(n_455),
.B(n_368),
.Y(n_580)
);

BUFx6f_ASAP7_75t_L g581 ( 
.A(n_459),
.Y(n_581)
);

INVx1_ASAP7_75t_L g582 ( 
.A(n_461),
.Y(n_582)
);

BUFx6f_ASAP7_75t_L g583 ( 
.A(n_459),
.Y(n_583)
);

INVx1_ASAP7_75t_L g584 ( 
.A(n_461),
.Y(n_584)
);

INVx1_ASAP7_75t_L g585 ( 
.A(n_504),
.Y(n_585)
);

BUFx3_ASAP7_75t_L g586 ( 
.A(n_504),
.Y(n_586)
);

INVx1_ASAP7_75t_L g587 ( 
.A(n_504),
.Y(n_587)
);

INVx2_ASAP7_75t_L g588 ( 
.A(n_482),
.Y(n_588)
);

NAND2xp33_ASAP7_75t_SL g589 ( 
.A(n_495),
.B(n_245),
.Y(n_589)
);

AND3x1_ASAP7_75t_L g590 ( 
.A(n_449),
.B(n_349),
.C(n_334),
.Y(n_590)
);

BUFx3_ASAP7_75t_L g591 ( 
.A(n_469),
.Y(n_591)
);

BUFx2_ASAP7_75t_L g592 ( 
.A(n_469),
.Y(n_592)
);

NAND2xp33_ASAP7_75t_L g593 ( 
.A(n_483),
.B(n_210),
.Y(n_593)
);

AOI22xp33_ASAP7_75t_L g594 ( 
.A1(n_511),
.A2(n_483),
.B1(n_484),
.B2(n_496),
.Y(n_594)
);

INVx1_ASAP7_75t_L g595 ( 
.A(n_515),
.Y(n_595)
);

BUFx6f_ASAP7_75t_L g596 ( 
.A(n_462),
.Y(n_596)
);

INVx2_ASAP7_75t_SL g597 ( 
.A(n_469),
.Y(n_597)
);

INVx1_ASAP7_75t_L g598 ( 
.A(n_515),
.Y(n_598)
);

INVx1_ASAP7_75t_L g599 ( 
.A(n_515),
.Y(n_599)
);

INVx1_ASAP7_75t_L g600 ( 
.A(n_522),
.Y(n_600)
);

NOR2xp33_ASAP7_75t_L g601 ( 
.A(n_478),
.B(n_421),
.Y(n_601)
);

INVx2_ASAP7_75t_L g602 ( 
.A(n_482),
.Y(n_602)
);

BUFx3_ASAP7_75t_L g603 ( 
.A(n_451),
.Y(n_603)
);

INVx5_ASAP7_75t_L g604 ( 
.A(n_453),
.Y(n_604)
);

INVx1_ASAP7_75t_L g605 ( 
.A(n_522),
.Y(n_605)
);

INVx4_ASAP7_75t_L g606 ( 
.A(n_462),
.Y(n_606)
);

INVx2_ASAP7_75t_L g607 ( 
.A(n_482),
.Y(n_607)
);

INVx2_ASAP7_75t_L g608 ( 
.A(n_462),
.Y(n_608)
);

INVx1_ASAP7_75t_L g609 ( 
.A(n_522),
.Y(n_609)
);

INVx1_ASAP7_75t_L g610 ( 
.A(n_522),
.Y(n_610)
);

INVx2_ASAP7_75t_L g611 ( 
.A(n_462),
.Y(n_611)
);

NAND2xp5_ASAP7_75t_SL g612 ( 
.A(n_481),
.B(n_363),
.Y(n_612)
);

INVx1_ASAP7_75t_SL g613 ( 
.A(n_481),
.Y(n_613)
);

NAND3xp33_ASAP7_75t_L g614 ( 
.A(n_445),
.B(n_367),
.C(n_364),
.Y(n_614)
);

NAND2xp5_ASAP7_75t_L g615 ( 
.A(n_498),
.B(n_301),
.Y(n_615)
);

BUFx4f_ASAP7_75t_L g616 ( 
.A(n_496),
.Y(n_616)
);

INVx5_ASAP7_75t_L g617 ( 
.A(n_453),
.Y(n_617)
);

AND2x2_ASAP7_75t_L g618 ( 
.A(n_445),
.B(n_489),
.Y(n_618)
);

INVx4_ASAP7_75t_L g619 ( 
.A(n_462),
.Y(n_619)
);

INVx2_ASAP7_75t_L g620 ( 
.A(n_462),
.Y(n_620)
);

INVx1_ASAP7_75t_L g621 ( 
.A(n_522),
.Y(n_621)
);

INVx2_ASAP7_75t_L g622 ( 
.A(n_466),
.Y(n_622)
);

BUFx3_ASAP7_75t_L g623 ( 
.A(n_451),
.Y(n_623)
);

OR2x6_ASAP7_75t_L g624 ( 
.A(n_471),
.B(n_291),
.Y(n_624)
);

INVx2_ASAP7_75t_L g625 ( 
.A(n_466),
.Y(n_625)
);

INVx4_ASAP7_75t_L g626 ( 
.A(n_465),
.Y(n_626)
);

INVx1_ASAP7_75t_L g627 ( 
.A(n_522),
.Y(n_627)
);

NAND2xp5_ASAP7_75t_SL g628 ( 
.A(n_507),
.B(n_247),
.Y(n_628)
);

NAND2xp5_ASAP7_75t_L g629 ( 
.A(n_483),
.B(n_232),
.Y(n_629)
);

OR2x2_ASAP7_75t_L g630 ( 
.A(n_489),
.B(n_367),
.Y(n_630)
);

INVx1_ASAP7_75t_L g631 ( 
.A(n_488),
.Y(n_631)
);

NAND2xp5_ASAP7_75t_SL g632 ( 
.A(n_521),
.B(n_247),
.Y(n_632)
);

NOR2xp33_ASAP7_75t_L g633 ( 
.A(n_458),
.B(n_361),
.Y(n_633)
);

AND3x2_ASAP7_75t_L g634 ( 
.A(n_449),
.B(n_234),
.C(n_333),
.Y(n_634)
);

BUFx6f_ASAP7_75t_L g635 ( 
.A(n_488),
.Y(n_635)
);

INVx1_ASAP7_75t_SL g636 ( 
.A(n_464),
.Y(n_636)
);

AND2x2_ASAP7_75t_L g637 ( 
.A(n_489),
.B(n_380),
.Y(n_637)
);

INVx1_ASAP7_75t_L g638 ( 
.A(n_488),
.Y(n_638)
);

BUFx10_ASAP7_75t_L g639 ( 
.A(n_491),
.Y(n_639)
);

INVx1_ASAP7_75t_L g640 ( 
.A(n_488),
.Y(n_640)
);

INVx2_ASAP7_75t_L g641 ( 
.A(n_466),
.Y(n_641)
);

INVx1_ASAP7_75t_L g642 ( 
.A(n_514),
.Y(n_642)
);

NAND2xp5_ASAP7_75t_L g643 ( 
.A(n_483),
.B(n_236),
.Y(n_643)
);

INVx5_ASAP7_75t_L g644 ( 
.A(n_453),
.Y(n_644)
);

INVx1_ASAP7_75t_SL g645 ( 
.A(n_520),
.Y(n_645)
);

INVx2_ASAP7_75t_L g646 ( 
.A(n_466),
.Y(n_646)
);

NAND2xp5_ASAP7_75t_SL g647 ( 
.A(n_491),
.B(n_281),
.Y(n_647)
);

BUFx6f_ASAP7_75t_L g648 ( 
.A(n_514),
.Y(n_648)
);

NAND2xp5_ASAP7_75t_SL g649 ( 
.A(n_491),
.B(n_281),
.Y(n_649)
);

AND2x2_ASAP7_75t_L g650 ( 
.A(n_491),
.B(n_380),
.Y(n_650)
);

NAND3xp33_ASAP7_75t_L g651 ( 
.A(n_499),
.B(n_382),
.C(n_387),
.Y(n_651)
);

INVx2_ASAP7_75t_L g652 ( 
.A(n_473),
.Y(n_652)
);

INVx1_ASAP7_75t_L g653 ( 
.A(n_514),
.Y(n_653)
);

INVx2_ASAP7_75t_L g654 ( 
.A(n_473),
.Y(n_654)
);

INVx1_ASAP7_75t_L g655 ( 
.A(n_514),
.Y(n_655)
);

INVx2_ASAP7_75t_L g656 ( 
.A(n_473),
.Y(n_656)
);

BUFx6f_ASAP7_75t_L g657 ( 
.A(n_465),
.Y(n_657)
);

BUFx10_ASAP7_75t_L g658 ( 
.A(n_499),
.Y(n_658)
);

INVx5_ASAP7_75t_L g659 ( 
.A(n_453),
.Y(n_659)
);

INVx2_ASAP7_75t_SL g660 ( 
.A(n_496),
.Y(n_660)
);

INVx1_ASAP7_75t_L g661 ( 
.A(n_486),
.Y(n_661)
);

AOI22xp33_ASAP7_75t_L g662 ( 
.A1(n_483),
.A2(n_271),
.B1(n_243),
.B2(n_385),
.Y(n_662)
);

CKINVDCx20_ASAP7_75t_R g663 ( 
.A(n_496),
.Y(n_663)
);

INVx4_ASAP7_75t_L g664 ( 
.A(n_465),
.Y(n_664)
);

INVx2_ASAP7_75t_L g665 ( 
.A(n_473),
.Y(n_665)
);

AND2x2_ASAP7_75t_SL g666 ( 
.A(n_499),
.B(n_243),
.Y(n_666)
);

AOI22xp33_ASAP7_75t_L g667 ( 
.A1(n_483),
.A2(n_271),
.B1(n_243),
.B2(n_385),
.Y(n_667)
);

BUFx3_ASAP7_75t_L g668 ( 
.A(n_499),
.Y(n_668)
);

INVx2_ASAP7_75t_SL g669 ( 
.A(n_518),
.Y(n_669)
);

NAND3xp33_ASAP7_75t_L g670 ( 
.A(n_446),
.B(n_382),
.C(n_387),
.Y(n_670)
);

CKINVDCx16_ASAP7_75t_R g671 ( 
.A(n_483),
.Y(n_671)
);

INVx2_ASAP7_75t_L g672 ( 
.A(n_486),
.Y(n_672)
);

INVx1_ASAP7_75t_L g673 ( 
.A(n_486),
.Y(n_673)
);

INVx2_ASAP7_75t_L g674 ( 
.A(n_501),
.Y(n_674)
);

INVx1_ASAP7_75t_L g675 ( 
.A(n_501),
.Y(n_675)
);

OR2x6_ASAP7_75t_L g676 ( 
.A(n_592),
.B(n_242),
.Y(n_676)
);

NOR2xp33_ASAP7_75t_L g677 ( 
.A(n_532),
.B(n_370),
.Y(n_677)
);

INVx2_ASAP7_75t_SL g678 ( 
.A(n_591),
.Y(n_678)
);

AOI22xp33_ASAP7_75t_L g679 ( 
.A1(n_550),
.A2(n_539),
.B1(n_618),
.B2(n_567),
.Y(n_679)
);

NAND2xp5_ASAP7_75t_SL g680 ( 
.A(n_558),
.B(n_186),
.Y(n_680)
);

NAND2xp5_ASAP7_75t_SL g681 ( 
.A(n_592),
.B(n_186),
.Y(n_681)
);

INVx1_ASAP7_75t_L g682 ( 
.A(n_631),
.Y(n_682)
);

NAND2xp33_ASAP7_75t_L g683 ( 
.A(n_594),
.B(n_662),
.Y(n_683)
);

AOI22xp33_ASAP7_75t_L g684 ( 
.A1(n_618),
.A2(n_453),
.B1(n_255),
.B2(n_258),
.Y(n_684)
);

AOI22xp5_ASAP7_75t_L g685 ( 
.A1(n_537),
.A2(n_374),
.B1(n_406),
.B2(n_379),
.Y(n_685)
);

OR2x2_ASAP7_75t_L g686 ( 
.A(n_566),
.B(n_444),
.Y(n_686)
);

NAND2xp5_ASAP7_75t_L g687 ( 
.A(n_597),
.B(n_453),
.Y(n_687)
);

INVxp67_ASAP7_75t_L g688 ( 
.A(n_566),
.Y(n_688)
);

NAND2xp5_ASAP7_75t_L g689 ( 
.A(n_597),
.B(n_453),
.Y(n_689)
);

NAND2xp5_ASAP7_75t_L g690 ( 
.A(n_568),
.B(n_501),
.Y(n_690)
);

NAND2xp5_ASAP7_75t_SL g691 ( 
.A(n_562),
.B(n_190),
.Y(n_691)
);

NAND2xp5_ASAP7_75t_SL g692 ( 
.A(n_615),
.B(n_190),
.Y(n_692)
);

OAI22xp33_ASAP7_75t_L g693 ( 
.A1(n_624),
.A2(n_329),
.B1(n_302),
.B2(n_276),
.Y(n_693)
);

NAND2xp5_ASAP7_75t_SL g694 ( 
.A(n_571),
.B(n_193),
.Y(n_694)
);

INVx2_ASAP7_75t_L g695 ( 
.A(n_672),
.Y(n_695)
);

NAND2xp33_ASAP7_75t_L g696 ( 
.A(n_667),
.B(n_350),
.Y(n_696)
);

NAND2xp5_ASAP7_75t_SL g697 ( 
.A(n_591),
.B(n_193),
.Y(n_697)
);

NAND2xp5_ASAP7_75t_L g698 ( 
.A(n_582),
.B(n_506),
.Y(n_698)
);

NAND2xp5_ASAP7_75t_L g699 ( 
.A(n_584),
.B(n_506),
.Y(n_699)
);

INVx1_ASAP7_75t_L g700 ( 
.A(n_585),
.Y(n_700)
);

AOI22xp33_ASAP7_75t_L g701 ( 
.A1(n_573),
.A2(n_264),
.B1(n_260),
.B2(n_315),
.Y(n_701)
);

NAND2xp5_ASAP7_75t_L g702 ( 
.A(n_587),
.B(n_506),
.Y(n_702)
);

INVx1_ASAP7_75t_L g703 ( 
.A(n_631),
.Y(n_703)
);

OR2x2_ASAP7_75t_L g704 ( 
.A(n_613),
.B(n_444),
.Y(n_704)
);

NAND2xp5_ASAP7_75t_L g705 ( 
.A(n_666),
.B(n_512),
.Y(n_705)
);

NAND3xp33_ASAP7_75t_L g706 ( 
.A(n_578),
.B(n_277),
.C(n_318),
.Y(n_706)
);

NAND2xp5_ASAP7_75t_L g707 ( 
.A(n_666),
.B(n_668),
.Y(n_707)
);

NAND2xp5_ASAP7_75t_L g708 ( 
.A(n_668),
.B(n_512),
.Y(n_708)
);

NAND2xp5_ASAP7_75t_L g709 ( 
.A(n_637),
.B(n_512),
.Y(n_709)
);

INVx4_ASAP7_75t_L g710 ( 
.A(n_604),
.Y(n_710)
);

BUFx2_ASAP7_75t_L g711 ( 
.A(n_590),
.Y(n_711)
);

BUFx3_ASAP7_75t_L g712 ( 
.A(n_540),
.Y(n_712)
);

INVx2_ASAP7_75t_L g713 ( 
.A(n_672),
.Y(n_713)
);

NOR2xp33_ASAP7_75t_L g714 ( 
.A(n_564),
.B(n_194),
.Y(n_714)
);

AOI22xp5_ASAP7_75t_L g715 ( 
.A1(n_663),
.A2(n_346),
.B1(n_194),
.B2(n_204),
.Y(n_715)
);

OAI22xp33_ASAP7_75t_L g716 ( 
.A1(n_624),
.A2(n_347),
.B1(n_294),
.B2(n_316),
.Y(n_716)
);

NAND2xp33_ASAP7_75t_L g717 ( 
.A(n_660),
.B(n_350),
.Y(n_717)
);

INVx2_ASAP7_75t_L g718 ( 
.A(n_674),
.Y(n_718)
);

NAND2xp5_ASAP7_75t_L g719 ( 
.A(n_637),
.B(n_517),
.Y(n_719)
);

INVx1_ASAP7_75t_L g720 ( 
.A(n_638),
.Y(n_720)
);

INVx1_ASAP7_75t_L g721 ( 
.A(n_638),
.Y(n_721)
);

INVx2_ASAP7_75t_L g722 ( 
.A(n_674),
.Y(n_722)
);

NOR2xp33_ASAP7_75t_L g723 ( 
.A(n_574),
.B(n_198),
.Y(n_723)
);

NAND2xp5_ASAP7_75t_SL g724 ( 
.A(n_601),
.B(n_198),
.Y(n_724)
);

BUFx6f_ASAP7_75t_SL g725 ( 
.A(n_669),
.Y(n_725)
);

NAND2xp5_ASAP7_75t_L g726 ( 
.A(n_650),
.B(n_517),
.Y(n_726)
);

INVxp67_ASAP7_75t_L g727 ( 
.A(n_612),
.Y(n_727)
);

OR2x2_ASAP7_75t_L g728 ( 
.A(n_624),
.B(n_446),
.Y(n_728)
);

INVx1_ASAP7_75t_L g729 ( 
.A(n_640),
.Y(n_729)
);

INVx2_ASAP7_75t_L g730 ( 
.A(n_622),
.Y(n_730)
);

BUFx3_ASAP7_75t_L g731 ( 
.A(n_540),
.Y(n_731)
);

NAND2xp5_ASAP7_75t_L g732 ( 
.A(n_650),
.B(n_517),
.Y(n_732)
);

NAND2xp5_ASAP7_75t_L g733 ( 
.A(n_640),
.B(n_447),
.Y(n_733)
);

INVx1_ASAP7_75t_L g734 ( 
.A(n_642),
.Y(n_734)
);

INVx2_ASAP7_75t_L g735 ( 
.A(n_622),
.Y(n_735)
);

INVx1_ASAP7_75t_L g736 ( 
.A(n_642),
.Y(n_736)
);

AND2x6_ASAP7_75t_SL g737 ( 
.A(n_633),
.B(n_447),
.Y(n_737)
);

BUFx3_ASAP7_75t_L g738 ( 
.A(n_586),
.Y(n_738)
);

CKINVDCx5p33_ASAP7_75t_R g739 ( 
.A(n_560),
.Y(n_739)
);

NOR3xp33_ASAP7_75t_L g740 ( 
.A(n_589),
.B(n_480),
.C(n_516),
.Y(n_740)
);

INVx1_ASAP7_75t_L g741 ( 
.A(n_653),
.Y(n_741)
);

NOR2xp33_ASAP7_75t_L g742 ( 
.A(n_570),
.B(n_204),
.Y(n_742)
);

NAND2xp5_ASAP7_75t_L g743 ( 
.A(n_653),
.B(n_655),
.Y(n_743)
);

INVx2_ASAP7_75t_L g744 ( 
.A(n_625),
.Y(n_744)
);

INVx2_ASAP7_75t_L g745 ( 
.A(n_625),
.Y(n_745)
);

NAND2xp5_ASAP7_75t_SL g746 ( 
.A(n_530),
.B(n_206),
.Y(n_746)
);

INVx2_ASAP7_75t_SL g747 ( 
.A(n_630),
.Y(n_747)
);

INVx2_ASAP7_75t_L g748 ( 
.A(n_641),
.Y(n_748)
);

NAND2xp5_ASAP7_75t_L g749 ( 
.A(n_655),
.B(n_448),
.Y(n_749)
);

INVx2_ASAP7_75t_L g750 ( 
.A(n_641),
.Y(n_750)
);

AOI22xp33_ASAP7_75t_L g751 ( 
.A1(n_663),
.A2(n_350),
.B1(n_243),
.B2(n_271),
.Y(n_751)
);

O2A1O1Ixp33_ASAP7_75t_L g752 ( 
.A1(n_660),
.A2(n_519),
.B(n_516),
.C(n_513),
.Y(n_752)
);

BUFx6f_ASAP7_75t_L g753 ( 
.A(n_635),
.Y(n_753)
);

INVx1_ASAP7_75t_L g754 ( 
.A(n_630),
.Y(n_754)
);

NAND3xp33_ASAP7_75t_L g755 ( 
.A(n_614),
.B(n_323),
.C(n_320),
.Y(n_755)
);

INVx2_ASAP7_75t_L g756 ( 
.A(n_646),
.Y(n_756)
);

INVxp67_ASAP7_75t_L g757 ( 
.A(n_636),
.Y(n_757)
);

INVx2_ASAP7_75t_L g758 ( 
.A(n_646),
.Y(n_758)
);

NAND2xp5_ASAP7_75t_L g759 ( 
.A(n_586),
.B(n_448),
.Y(n_759)
);

NAND2xp5_ASAP7_75t_SL g760 ( 
.A(n_604),
.B(n_206),
.Y(n_760)
);

NAND2xp5_ASAP7_75t_SL g761 ( 
.A(n_604),
.B(n_207),
.Y(n_761)
);

INVx2_ASAP7_75t_L g762 ( 
.A(n_652),
.Y(n_762)
);

AND2x2_ASAP7_75t_L g763 ( 
.A(n_580),
.B(n_456),
.Y(n_763)
);

BUFx8_ASAP7_75t_L g764 ( 
.A(n_669),
.Y(n_764)
);

INVx1_ASAP7_75t_L g765 ( 
.A(n_652),
.Y(n_765)
);

OR2x2_ASAP7_75t_L g766 ( 
.A(n_624),
.B(n_456),
.Y(n_766)
);

NAND2xp5_ASAP7_75t_L g767 ( 
.A(n_554),
.B(n_467),
.Y(n_767)
);

NAND2xp5_ASAP7_75t_L g768 ( 
.A(n_554),
.B(n_467),
.Y(n_768)
);

NAND2xp5_ASAP7_75t_L g769 ( 
.A(n_554),
.B(n_470),
.Y(n_769)
);

INVx2_ASAP7_75t_L g770 ( 
.A(n_654),
.Y(n_770)
);

NAND2xp5_ASAP7_75t_SL g771 ( 
.A(n_604),
.B(n_207),
.Y(n_771)
);

NAND2xp5_ASAP7_75t_L g772 ( 
.A(n_554),
.B(n_470),
.Y(n_772)
);

NAND2xp5_ASAP7_75t_SL g773 ( 
.A(n_604),
.B(n_216),
.Y(n_773)
);

NAND2xp5_ASAP7_75t_L g774 ( 
.A(n_671),
.B(n_472),
.Y(n_774)
);

AOI22xp33_ASAP7_75t_L g775 ( 
.A1(n_579),
.A2(n_350),
.B1(n_271),
.B2(n_243),
.Y(n_775)
);

INVxp33_ASAP7_75t_L g776 ( 
.A(n_543),
.Y(n_776)
);

BUFx6f_ASAP7_75t_L g777 ( 
.A(n_635),
.Y(n_777)
);

INVxp67_ASAP7_75t_SL g778 ( 
.A(n_635),
.Y(n_778)
);

INVx2_ASAP7_75t_L g779 ( 
.A(n_654),
.Y(n_779)
);

NOR3xp33_ASAP7_75t_L g780 ( 
.A(n_563),
.B(n_519),
.C(n_513),
.Y(n_780)
);

NAND2xp5_ASAP7_75t_L g781 ( 
.A(n_635),
.B(n_472),
.Y(n_781)
);

INVx1_ASAP7_75t_L g782 ( 
.A(n_656),
.Y(n_782)
);

NAND2xp5_ASAP7_75t_L g783 ( 
.A(n_635),
.B(n_477),
.Y(n_783)
);

INVx1_ASAP7_75t_L g784 ( 
.A(n_656),
.Y(n_784)
);

NAND2xp5_ASAP7_75t_L g785 ( 
.A(n_648),
.B(n_477),
.Y(n_785)
);

NOR2xp33_ASAP7_75t_L g786 ( 
.A(n_628),
.B(n_216),
.Y(n_786)
);

INVx2_ASAP7_75t_SL g787 ( 
.A(n_616),
.Y(n_787)
);

NAND2xp5_ASAP7_75t_L g788 ( 
.A(n_648),
.B(n_480),
.Y(n_788)
);

NAND2xp5_ASAP7_75t_L g789 ( 
.A(n_648),
.B(n_487),
.Y(n_789)
);

AND2x2_ASAP7_75t_L g790 ( 
.A(n_639),
.B(n_487),
.Y(n_790)
);

NAND2xp5_ASAP7_75t_SL g791 ( 
.A(n_617),
.B(n_218),
.Y(n_791)
);

INVx2_ASAP7_75t_L g792 ( 
.A(n_665),
.Y(n_792)
);

NAND2xp5_ASAP7_75t_L g793 ( 
.A(n_648),
.B(n_493),
.Y(n_793)
);

NAND2xp5_ASAP7_75t_L g794 ( 
.A(n_579),
.B(n_493),
.Y(n_794)
);

NOR2xp33_ASAP7_75t_L g795 ( 
.A(n_647),
.B(n_218),
.Y(n_795)
);

BUFx6f_ASAP7_75t_SL g796 ( 
.A(n_579),
.Y(n_796)
);

O2A1O1Ixp33_ASAP7_75t_L g797 ( 
.A1(n_629),
.A2(n_509),
.B(n_508),
.C(n_505),
.Y(n_797)
);

HB1xp67_ASAP7_75t_L g798 ( 
.A(n_645),
.Y(n_798)
);

NOR2xp33_ASAP7_75t_L g799 ( 
.A(n_649),
.B(n_222),
.Y(n_799)
);

AND2x6_ASAP7_75t_SL g800 ( 
.A(n_560),
.B(n_494),
.Y(n_800)
);

INVx1_ASAP7_75t_L g801 ( 
.A(n_665),
.Y(n_801)
);

INVx2_ASAP7_75t_L g802 ( 
.A(n_529),
.Y(n_802)
);

INVx1_ASAP7_75t_L g803 ( 
.A(n_661),
.Y(n_803)
);

NAND2xp5_ASAP7_75t_SL g804 ( 
.A(n_617),
.B(n_222),
.Y(n_804)
);

OAI21xp5_ASAP7_75t_L g805 ( 
.A1(n_616),
.A2(n_465),
.B(n_508),
.Y(n_805)
);

NAND2xp5_ASAP7_75t_SL g806 ( 
.A(n_617),
.B(n_259),
.Y(n_806)
);

O2A1O1Ixp33_ASAP7_75t_L g807 ( 
.A1(n_643),
.A2(n_509),
.B(n_505),
.C(n_503),
.Y(n_807)
);

NAND2xp5_ASAP7_75t_L g808 ( 
.A(n_579),
.B(n_494),
.Y(n_808)
);

NOR2xp33_ASAP7_75t_SL g809 ( 
.A(n_542),
.B(n_281),
.Y(n_809)
);

AND2x2_ASAP7_75t_L g810 ( 
.A(n_639),
.B(n_497),
.Y(n_810)
);

CKINVDCx5p33_ASAP7_75t_R g811 ( 
.A(n_577),
.Y(n_811)
);

INVx2_ASAP7_75t_SL g812 ( 
.A(n_616),
.Y(n_812)
);

AOI22xp33_ASAP7_75t_L g813 ( 
.A1(n_579),
.A2(n_350),
.B1(n_271),
.B2(n_503),
.Y(n_813)
);

INVx1_ASAP7_75t_L g814 ( 
.A(n_661),
.Y(n_814)
);

INVx1_ASAP7_75t_L g815 ( 
.A(n_673),
.Y(n_815)
);

OAI22xp5_ASAP7_75t_L g816 ( 
.A1(n_603),
.A2(n_298),
.B1(n_259),
.B2(n_261),
.Y(n_816)
);

INVx2_ASAP7_75t_L g817 ( 
.A(n_529),
.Y(n_817)
);

INVx2_ASAP7_75t_L g818 ( 
.A(n_531),
.Y(n_818)
);

NOR2xp33_ASAP7_75t_L g819 ( 
.A(n_536),
.B(n_261),
.Y(n_819)
);

INVx2_ASAP7_75t_L g820 ( 
.A(n_531),
.Y(n_820)
);

NOR2xp67_ASAP7_75t_L g821 ( 
.A(n_670),
.B(n_500),
.Y(n_821)
);

HB1xp67_ASAP7_75t_L g822 ( 
.A(n_577),
.Y(n_822)
);

INVx1_ASAP7_75t_L g823 ( 
.A(n_673),
.Y(n_823)
);

INVx2_ASAP7_75t_L g824 ( 
.A(n_534),
.Y(n_824)
);

INVx2_ASAP7_75t_L g825 ( 
.A(n_534),
.Y(n_825)
);

INVxp33_ASAP7_75t_L g826 ( 
.A(n_632),
.Y(n_826)
);

OR2x6_ASAP7_75t_L g827 ( 
.A(n_651),
.B(n_603),
.Y(n_827)
);

INVx2_ASAP7_75t_L g828 ( 
.A(n_675),
.Y(n_828)
);

INVx2_ASAP7_75t_SL g829 ( 
.A(n_639),
.Y(n_829)
);

INVx1_ASAP7_75t_L g830 ( 
.A(n_675),
.Y(n_830)
);

NOR2xp33_ASAP7_75t_L g831 ( 
.A(n_634),
.B(n_282),
.Y(n_831)
);

NOR2xp33_ASAP7_75t_L g832 ( 
.A(n_658),
.B(n_282),
.Y(n_832)
);

INVx4_ASAP7_75t_L g833 ( 
.A(n_617),
.Y(n_833)
);

NAND2xp5_ASAP7_75t_L g834 ( 
.A(n_608),
.B(n_497),
.Y(n_834)
);

NAND2xp5_ASAP7_75t_L g835 ( 
.A(n_608),
.B(n_500),
.Y(n_835)
);

NAND2xp33_ASAP7_75t_L g836 ( 
.A(n_617),
.B(n_350),
.Y(n_836)
);

NAND2xp5_ASAP7_75t_SL g837 ( 
.A(n_644),
.B(n_284),
.Y(n_837)
);

NOR2xp33_ASAP7_75t_L g838 ( 
.A(n_658),
.B(n_284),
.Y(n_838)
);

NOR2xp33_ASAP7_75t_L g839 ( 
.A(n_658),
.B(n_292),
.Y(n_839)
);

INVx2_ASAP7_75t_L g840 ( 
.A(n_623),
.Y(n_840)
);

INVx1_ASAP7_75t_L g841 ( 
.A(n_623),
.Y(n_841)
);

INVx1_ASAP7_75t_L g842 ( 
.A(n_523),
.Y(n_842)
);

INVx1_ASAP7_75t_L g843 ( 
.A(n_523),
.Y(n_843)
);

INVx2_ASAP7_75t_L g844 ( 
.A(n_611),
.Y(n_844)
);

NAND2xp5_ASAP7_75t_L g845 ( 
.A(n_611),
.B(n_465),
.Y(n_845)
);

INVxp67_ASAP7_75t_SL g846 ( 
.A(n_581),
.Y(n_846)
);

INVx3_ASAP7_75t_L g847 ( 
.A(n_753),
.Y(n_847)
);

INVx2_ASAP7_75t_L g848 ( 
.A(n_730),
.Y(n_848)
);

INVx1_ASAP7_75t_L g849 ( 
.A(n_682),
.Y(n_849)
);

O2A1O1Ixp33_ASAP7_75t_L g850 ( 
.A1(n_683),
.A2(n_707),
.B(n_774),
.C(n_754),
.Y(n_850)
);

AOI21xp5_ASAP7_75t_L g851 ( 
.A1(n_690),
.A2(n_547),
.B(n_644),
.Y(n_851)
);

INVx2_ASAP7_75t_L g852 ( 
.A(n_730),
.Y(n_852)
);

AOI21xp5_ASAP7_75t_L g853 ( 
.A1(n_710),
.A2(n_547),
.B(n_644),
.Y(n_853)
);

AND2x2_ASAP7_75t_L g854 ( 
.A(n_704),
.B(n_270),
.Y(n_854)
);

CKINVDCx5p33_ASAP7_75t_R g855 ( 
.A(n_739),
.Y(n_855)
);

HB1xp67_ASAP7_75t_L g856 ( 
.A(n_757),
.Y(n_856)
);

AOI21xp33_ASAP7_75t_L g857 ( 
.A1(n_819),
.A2(n_742),
.B(n_677),
.Y(n_857)
);

AOI21xp5_ASAP7_75t_L g858 ( 
.A1(n_710),
.A2(n_659),
.B(n_644),
.Y(n_858)
);

NAND2xp5_ASAP7_75t_SL g859 ( 
.A(n_787),
.B(n_644),
.Y(n_859)
);

OAI21xp5_ASAP7_75t_L g860 ( 
.A1(n_683),
.A2(n_620),
.B(n_556),
.Y(n_860)
);

AOI22xp5_ASAP7_75t_L g861 ( 
.A1(n_763),
.A2(n_541),
.B1(n_524),
.B2(n_627),
.Y(n_861)
);

AOI22xp5_ASAP7_75t_L g862 ( 
.A1(n_763),
.A2(n_541),
.B1(n_524),
.B2(n_627),
.Y(n_862)
);

NAND2xp5_ASAP7_75t_L g863 ( 
.A(n_790),
.B(n_620),
.Y(n_863)
);

AOI21xp5_ASAP7_75t_L g864 ( 
.A1(n_710),
.A2(n_659),
.B(n_606),
.Y(n_864)
);

HB1xp67_ASAP7_75t_L g865 ( 
.A(n_798),
.Y(n_865)
);

AND2x2_ASAP7_75t_L g866 ( 
.A(n_704),
.B(n_354),
.Y(n_866)
);

NAND2xp5_ASAP7_75t_SL g867 ( 
.A(n_787),
.B(n_659),
.Y(n_867)
);

NAND2xp5_ASAP7_75t_L g868 ( 
.A(n_790),
.B(n_810),
.Y(n_868)
);

OAI21xp5_ASAP7_75t_L g869 ( 
.A1(n_805),
.A2(n_527),
.B(n_556),
.Y(n_869)
);

NAND2xp5_ASAP7_75t_SL g870 ( 
.A(n_812),
.B(n_659),
.Y(n_870)
);

NAND2xp5_ASAP7_75t_SL g871 ( 
.A(n_812),
.B(n_659),
.Y(n_871)
);

AO21x1_ASAP7_75t_L g872 ( 
.A1(n_841),
.A2(n_593),
.B(n_525),
.Y(n_872)
);

OAI21xp5_ASAP7_75t_L g873 ( 
.A1(n_717),
.A2(n_705),
.B(n_689),
.Y(n_873)
);

NAND2xp5_ASAP7_75t_L g874 ( 
.A(n_810),
.B(n_527),
.Y(n_874)
);

OAI21xp5_ASAP7_75t_L g875 ( 
.A1(n_717),
.A2(n_687),
.B(n_752),
.Y(n_875)
);

A2O1A1Ixp33_ASAP7_75t_L g876 ( 
.A1(n_679),
.A2(n_593),
.B(n_348),
.C(n_286),
.Y(n_876)
);

NAND2xp5_ASAP7_75t_SL g877 ( 
.A(n_833),
.B(n_581),
.Y(n_877)
);

NAND2xp5_ASAP7_75t_L g878 ( 
.A(n_751),
.B(n_527),
.Y(n_878)
);

AOI21x1_ASAP7_75t_L g879 ( 
.A1(n_708),
.A2(n_572),
.B(n_555),
.Y(n_879)
);

NAND2xp5_ASAP7_75t_L g880 ( 
.A(n_714),
.B(n_556),
.Y(n_880)
);

NOR2x1p5_ASAP7_75t_SL g881 ( 
.A(n_840),
.B(n_535),
.Y(n_881)
);

HB1xp67_ASAP7_75t_L g882 ( 
.A(n_688),
.Y(n_882)
);

OR2x6_ASAP7_75t_L g883 ( 
.A(n_676),
.B(n_535),
.Y(n_883)
);

NAND2xp5_ASAP7_75t_L g884 ( 
.A(n_723),
.B(n_557),
.Y(n_884)
);

NAND2xp5_ASAP7_75t_L g885 ( 
.A(n_678),
.B(n_557),
.Y(n_885)
);

AOI21xp5_ASAP7_75t_L g886 ( 
.A1(n_833),
.A2(n_619),
.B(n_526),
.Y(n_886)
);

INVx1_ASAP7_75t_L g887 ( 
.A(n_703),
.Y(n_887)
);

AOI21xp5_ASAP7_75t_L g888 ( 
.A1(n_833),
.A2(n_619),
.B(n_526),
.Y(n_888)
);

INVx1_ASAP7_75t_L g889 ( 
.A(n_729),
.Y(n_889)
);

NOR2xp33_ASAP7_75t_L g890 ( 
.A(n_727),
.B(n_557),
.Y(n_890)
);

AOI21xp5_ASAP7_75t_L g891 ( 
.A1(n_778),
.A2(n_526),
.B(n_619),
.Y(n_891)
);

INVxp67_ASAP7_75t_L g892 ( 
.A(n_686),
.Y(n_892)
);

INVx2_ASAP7_75t_SL g893 ( 
.A(n_686),
.Y(n_893)
);

NOR2xp33_ASAP7_75t_L g894 ( 
.A(n_747),
.B(n_525),
.Y(n_894)
);

INVx1_ASAP7_75t_L g895 ( 
.A(n_729),
.Y(n_895)
);

INVxp67_ASAP7_75t_L g896 ( 
.A(n_822),
.Y(n_896)
);

AND2x2_ASAP7_75t_L g897 ( 
.A(n_747),
.B(n_184),
.Y(n_897)
);

NAND2xp5_ASAP7_75t_L g898 ( 
.A(n_678),
.B(n_709),
.Y(n_898)
);

NAND2xp5_ASAP7_75t_SL g899 ( 
.A(n_829),
.B(n_840),
.Y(n_899)
);

INVx2_ASAP7_75t_L g900 ( 
.A(n_735),
.Y(n_900)
);

AOI21xp5_ASAP7_75t_L g901 ( 
.A1(n_846),
.A2(n_726),
.B(n_719),
.Y(n_901)
);

NAND2xp5_ASAP7_75t_L g902 ( 
.A(n_732),
.B(n_528),
.Y(n_902)
);

NAND2xp5_ASAP7_75t_L g903 ( 
.A(n_759),
.B(n_528),
.Y(n_903)
);

OAI21xp5_ASAP7_75t_L g904 ( 
.A1(n_743),
.A2(n_552),
.B(n_545),
.Y(n_904)
);

AOI21xp5_ASAP7_75t_L g905 ( 
.A1(n_767),
.A2(n_606),
.B(n_581),
.Y(n_905)
);

INVx2_ASAP7_75t_L g906 ( 
.A(n_735),
.Y(n_906)
);

NAND2xp5_ASAP7_75t_L g907 ( 
.A(n_700),
.B(n_533),
.Y(n_907)
);

INVx2_ASAP7_75t_SL g908 ( 
.A(n_728),
.Y(n_908)
);

BUFx2_ASAP7_75t_L g909 ( 
.A(n_739),
.Y(n_909)
);

AOI21xp5_ASAP7_75t_L g910 ( 
.A1(n_768),
.A2(n_581),
.B(n_583),
.Y(n_910)
);

HB1xp67_ASAP7_75t_L g911 ( 
.A(n_676),
.Y(n_911)
);

BUFx2_ASAP7_75t_L g912 ( 
.A(n_811),
.Y(n_912)
);

INVx2_ASAP7_75t_L g913 ( 
.A(n_744),
.Y(n_913)
);

NAND2xp5_ASAP7_75t_L g914 ( 
.A(n_736),
.B(n_533),
.Y(n_914)
);

AOI21xp5_ASAP7_75t_L g915 ( 
.A1(n_769),
.A2(n_583),
.B(n_596),
.Y(n_915)
);

NAND2xp5_ASAP7_75t_L g916 ( 
.A(n_720),
.B(n_545),
.Y(n_916)
);

BUFx2_ASAP7_75t_L g917 ( 
.A(n_811),
.Y(n_917)
);

A2O1A1Ixp33_ASAP7_75t_L g918 ( 
.A1(n_701),
.A2(n_289),
.B(n_304),
.C(n_295),
.Y(n_918)
);

INVx2_ASAP7_75t_L g919 ( 
.A(n_744),
.Y(n_919)
);

NAND2xp5_ASAP7_75t_L g920 ( 
.A(n_721),
.B(n_552),
.Y(n_920)
);

NAND2xp5_ASAP7_75t_L g921 ( 
.A(n_734),
.B(n_553),
.Y(n_921)
);

NAND2xp5_ASAP7_75t_L g922 ( 
.A(n_741),
.B(n_553),
.Y(n_922)
);

OAI21xp5_ASAP7_75t_L g923 ( 
.A1(n_841),
.A2(n_576),
.B(n_555),
.Y(n_923)
);

NAND2xp5_ASAP7_75t_L g924 ( 
.A(n_772),
.B(n_561),
.Y(n_924)
);

NAND2xp5_ASAP7_75t_SL g925 ( 
.A(n_829),
.B(n_583),
.Y(n_925)
);

BUFx12f_ASAP7_75t_L g926 ( 
.A(n_800),
.Y(n_926)
);

OAI21xp5_ASAP7_75t_L g927 ( 
.A1(n_765),
.A2(n_561),
.B(n_565),
.Y(n_927)
);

OAI22xp5_ASAP7_75t_L g928 ( 
.A1(n_827),
.A2(n_565),
.B1(n_621),
.B2(n_610),
.Y(n_928)
);

INVx2_ASAP7_75t_L g929 ( 
.A(n_745),
.Y(n_929)
);

AOI21xp5_ASAP7_75t_L g930 ( 
.A1(n_836),
.A2(n_583),
.B(n_596),
.Y(n_930)
);

A2O1A1Ixp33_ASAP7_75t_L g931 ( 
.A1(n_795),
.A2(n_283),
.B(n_343),
.C(n_344),
.Y(n_931)
);

AND2x2_ASAP7_75t_L g932 ( 
.A(n_711),
.B(n_188),
.Y(n_932)
);

NOR2x1_ASAP7_75t_R g933 ( 
.A(n_711),
.B(n_188),
.Y(n_933)
);

BUFx3_ASAP7_75t_L g934 ( 
.A(n_712),
.Y(n_934)
);

NAND2xp5_ASAP7_75t_SL g935 ( 
.A(n_753),
.B(n_583),
.Y(n_935)
);

NOR2xp33_ASAP7_75t_L g936 ( 
.A(n_715),
.B(n_569),
.Y(n_936)
);

NOR2xp33_ASAP7_75t_L g937 ( 
.A(n_826),
.B(n_569),
.Y(n_937)
);

NAND2xp5_ASAP7_75t_L g938 ( 
.A(n_832),
.B(n_572),
.Y(n_938)
);

AOI21x1_ASAP7_75t_L g939 ( 
.A1(n_733),
.A2(n_599),
.B(n_576),
.Y(n_939)
);

INVx3_ASAP7_75t_L g940 ( 
.A(n_753),
.Y(n_940)
);

NAND2xp5_ASAP7_75t_SL g941 ( 
.A(n_753),
.B(n_596),
.Y(n_941)
);

BUFx3_ASAP7_75t_L g942 ( 
.A(n_712),
.Y(n_942)
);

NOR2xp33_ASAP7_75t_L g943 ( 
.A(n_826),
.B(n_716),
.Y(n_943)
);

OAI21xp5_ASAP7_75t_L g944 ( 
.A1(n_765),
.A2(n_598),
.B(n_595),
.Y(n_944)
);

A2O1A1Ixp33_ASAP7_75t_L g945 ( 
.A1(n_799),
.A2(n_213),
.B(n_239),
.C(n_283),
.Y(n_945)
);

NAND2xp5_ASAP7_75t_SL g946 ( 
.A(n_753),
.B(n_596),
.Y(n_946)
);

AOI21xp5_ASAP7_75t_L g947 ( 
.A1(n_836),
.A2(n_596),
.B(n_465),
.Y(n_947)
);

AND2x4_ASAP7_75t_L g948 ( 
.A(n_731),
.B(n_595),
.Y(n_948)
);

NAND2xp5_ASAP7_75t_L g949 ( 
.A(n_838),
.B(n_598),
.Y(n_949)
);

INVx1_ASAP7_75t_SL g950 ( 
.A(n_728),
.Y(n_950)
);

BUFx6f_ASAP7_75t_L g951 ( 
.A(n_777),
.Y(n_951)
);

NAND2xp5_ASAP7_75t_SL g952 ( 
.A(n_777),
.B(n_599),
.Y(n_952)
);

INVx1_ASAP7_75t_SL g953 ( 
.A(n_766),
.Y(n_953)
);

NAND2xp5_ASAP7_75t_L g954 ( 
.A(n_839),
.B(n_600),
.Y(n_954)
);

AOI21xp5_ASAP7_75t_L g955 ( 
.A1(n_781),
.A2(n_664),
.B(n_626),
.Y(n_955)
);

NAND2xp5_ASAP7_75t_L g956 ( 
.A(n_694),
.B(n_749),
.Y(n_956)
);

CKINVDCx6p67_ASAP7_75t_R g957 ( 
.A(n_725),
.Y(n_957)
);

NAND2xp5_ASAP7_75t_SL g958 ( 
.A(n_777),
.B(n_600),
.Y(n_958)
);

INVx2_ASAP7_75t_L g959 ( 
.A(n_745),
.Y(n_959)
);

AOI21xp5_ASAP7_75t_L g960 ( 
.A1(n_783),
.A2(n_788),
.B(n_785),
.Y(n_960)
);

BUFx8_ASAP7_75t_L g961 ( 
.A(n_725),
.Y(n_961)
);

AOI21xp5_ASAP7_75t_L g962 ( 
.A1(n_789),
.A2(n_664),
.B(n_626),
.Y(n_962)
);

INVx2_ASAP7_75t_L g963 ( 
.A(n_748),
.Y(n_963)
);

AOI22xp33_ASAP7_75t_L g964 ( 
.A1(n_696),
.A2(n_200),
.B1(n_191),
.B2(n_209),
.Y(n_964)
);

O2A1O1Ixp5_ASAP7_75t_L g965 ( 
.A1(n_691),
.A2(n_605),
.B(n_609),
.C(n_621),
.Y(n_965)
);

INVx2_ASAP7_75t_L g966 ( 
.A(n_750),
.Y(n_966)
);

AOI22x1_ASAP7_75t_L g967 ( 
.A1(n_844),
.A2(n_605),
.B1(n_609),
.B2(n_610),
.Y(n_967)
);

NAND2xp5_ASAP7_75t_L g968 ( 
.A(n_842),
.B(n_538),
.Y(n_968)
);

A2O1A1Ixp33_ASAP7_75t_L g969 ( 
.A1(n_786),
.A2(n_189),
.B(n_200),
.C(n_209),
.Y(n_969)
);

O2A1O1Ixp33_ASAP7_75t_L g970 ( 
.A1(n_746),
.A2(n_549),
.B(n_538),
.C(n_544),
.Y(n_970)
);

OR2x2_ASAP7_75t_L g971 ( 
.A(n_766),
.B(n_189),
.Y(n_971)
);

NAND2xp5_ASAP7_75t_L g972 ( 
.A(n_842),
.B(n_544),
.Y(n_972)
);

O2A1O1Ixp33_ASAP7_75t_L g973 ( 
.A1(n_680),
.A2(n_692),
.B(n_696),
.C(n_740),
.Y(n_973)
);

BUFx6f_ASAP7_75t_L g974 ( 
.A(n_777),
.Y(n_974)
);

NOR2xp33_ASAP7_75t_L g975 ( 
.A(n_809),
.B(n_332),
.Y(n_975)
);

NAND2x1p5_ASAP7_75t_L g976 ( 
.A(n_731),
.B(n_546),
.Y(n_976)
);

AOI21x1_ASAP7_75t_L g977 ( 
.A1(n_793),
.A2(n_546),
.B(n_548),
.Y(n_977)
);

HB1xp67_ASAP7_75t_L g978 ( 
.A(n_676),
.Y(n_978)
);

NOR2xp33_ASAP7_75t_R g979 ( 
.A(n_737),
.B(n_292),
.Y(n_979)
);

BUFx3_ASAP7_75t_L g980 ( 
.A(n_738),
.Y(n_980)
);

NAND2xp5_ASAP7_75t_L g981 ( 
.A(n_780),
.B(n_548),
.Y(n_981)
);

NAND2xp5_ASAP7_75t_L g982 ( 
.A(n_803),
.B(n_815),
.Y(n_982)
);

NAND2xp5_ASAP7_75t_SL g983 ( 
.A(n_777),
.B(n_549),
.Y(n_983)
);

NAND2xp5_ASAP7_75t_L g984 ( 
.A(n_803),
.B(n_551),
.Y(n_984)
);

NAND2xp5_ASAP7_75t_SL g985 ( 
.A(n_750),
.B(n_551),
.Y(n_985)
);

AND2x4_ASAP7_75t_L g986 ( 
.A(n_738),
.B(n_559),
.Y(n_986)
);

OAI21xp5_ASAP7_75t_L g987 ( 
.A1(n_782),
.A2(n_559),
.B(n_607),
.Y(n_987)
);

INVx2_ASAP7_75t_L g988 ( 
.A(n_756),
.Y(n_988)
);

NAND2xp5_ASAP7_75t_L g989 ( 
.A(n_815),
.B(n_575),
.Y(n_989)
);

NAND2xp5_ASAP7_75t_L g990 ( 
.A(n_823),
.B(n_575),
.Y(n_990)
);

OAI22xp5_ASAP7_75t_L g991 ( 
.A1(n_827),
.A2(n_588),
.B1(n_602),
.B2(n_607),
.Y(n_991)
);

NOR2xp33_ASAP7_75t_L g992 ( 
.A(n_681),
.B(n_336),
.Y(n_992)
);

NOR2xp33_ASAP7_75t_L g993 ( 
.A(n_724),
.B(n_339),
.Y(n_993)
);

A2O1A1Ixp33_ASAP7_75t_L g994 ( 
.A1(n_776),
.A2(n_295),
.B(n_289),
.C(n_286),
.Y(n_994)
);

INVx4_ASAP7_75t_L g995 ( 
.A(n_827),
.Y(n_995)
);

AOI21xp5_ASAP7_75t_L g996 ( 
.A1(n_698),
.A2(n_664),
.B(n_626),
.Y(n_996)
);

INVxp67_ASAP7_75t_L g997 ( 
.A(n_831),
.Y(n_997)
);

NOR2xp33_ASAP7_75t_L g998 ( 
.A(n_816),
.B(n_191),
.Y(n_998)
);

OAI321xp33_ASAP7_75t_L g999 ( 
.A1(n_693),
.A2(n_239),
.A3(n_213),
.B1(n_211),
.B2(n_304),
.C(n_343),
.Y(n_999)
);

INVx1_ASAP7_75t_SL g1000 ( 
.A(n_685),
.Y(n_1000)
);

CKINVDCx5p33_ASAP7_75t_R g1001 ( 
.A(n_725),
.Y(n_1001)
);

A2O1A1Ixp33_ASAP7_75t_L g1002 ( 
.A1(n_776),
.A2(n_211),
.B(n_352),
.C(n_348),
.Y(n_1002)
);

NAND2xp5_ASAP7_75t_L g1003 ( 
.A(n_823),
.B(n_588),
.Y(n_1003)
);

NAND2xp5_ASAP7_75t_L g1004 ( 
.A(n_814),
.B(n_602),
.Y(n_1004)
);

AOI21xp5_ASAP7_75t_L g1005 ( 
.A1(n_699),
.A2(n_657),
.B(n_340),
.Y(n_1005)
);

NAND2xp5_ASAP7_75t_L g1006 ( 
.A(n_830),
.B(n_340),
.Y(n_1006)
);

NAND2xp5_ASAP7_75t_L g1007 ( 
.A(n_782),
.B(n_312),
.Y(n_1007)
);

NAND2xp5_ASAP7_75t_L g1008 ( 
.A(n_834),
.B(n_312),
.Y(n_1008)
);

NAND2xp5_ASAP7_75t_L g1009 ( 
.A(n_835),
.B(n_341),
.Y(n_1009)
);

BUFx3_ASAP7_75t_L g1010 ( 
.A(n_764),
.Y(n_1010)
);

NOR2xp33_ASAP7_75t_L g1011 ( 
.A(n_706),
.B(n_697),
.Y(n_1011)
);

NAND2xp5_ASAP7_75t_SL g1012 ( 
.A(n_756),
.B(n_341),
.Y(n_1012)
);

NAND2xp5_ASAP7_75t_L g1013 ( 
.A(n_828),
.B(n_309),
.Y(n_1013)
);

BUFx4f_ASAP7_75t_L g1014 ( 
.A(n_827),
.Y(n_1014)
);

NAND2xp5_ASAP7_75t_SL g1015 ( 
.A(n_758),
.B(n_309),
.Y(n_1015)
);

AND2x2_ASAP7_75t_L g1016 ( 
.A(n_821),
.B(n_344),
.Y(n_1016)
);

INVx2_ASAP7_75t_L g1017 ( 
.A(n_758),
.Y(n_1017)
);

NOR2xp33_ASAP7_75t_L g1018 ( 
.A(n_755),
.B(n_843),
.Y(n_1018)
);

AOI21xp5_ASAP7_75t_L g1019 ( 
.A1(n_702),
.A2(n_657),
.B(n_307),
.Y(n_1019)
);

OAI22xp5_ASAP7_75t_L g1020 ( 
.A1(n_684),
.A2(n_796),
.B1(n_813),
.B2(n_775),
.Y(n_1020)
);

NAND2xp5_ASAP7_75t_L g1021 ( 
.A(n_762),
.B(n_307),
.Y(n_1021)
);

INVx3_ASAP7_75t_L g1022 ( 
.A(n_762),
.Y(n_1022)
);

INVx2_ASAP7_75t_L g1023 ( 
.A(n_695),
.Y(n_1023)
);

NOR2xp33_ASAP7_75t_L g1024 ( 
.A(n_784),
.B(n_352),
.Y(n_1024)
);

NAND2xp5_ASAP7_75t_SL g1025 ( 
.A(n_770),
.B(n_346),
.Y(n_1025)
);

NAND2xp5_ASAP7_75t_L g1026 ( 
.A(n_770),
.B(n_779),
.Y(n_1026)
);

NAND2xp5_ASAP7_75t_L g1027 ( 
.A(n_779),
.B(n_345),
.Y(n_1027)
);

AOI21xp5_ASAP7_75t_L g1028 ( 
.A1(n_845),
.A2(n_657),
.B(n_345),
.Y(n_1028)
);

OR2x6_ASAP7_75t_L g1029 ( 
.A(n_797),
.B(n_657),
.Y(n_1029)
);

NAND2xp5_ASAP7_75t_L g1030 ( 
.A(n_792),
.B(n_306),
.Y(n_1030)
);

BUFx8_ASAP7_75t_L g1031 ( 
.A(n_796),
.Y(n_1031)
);

A2O1A1Ixp33_ASAP7_75t_L g1032 ( 
.A1(n_807),
.A2(n_306),
.B(n_298),
.C(n_297),
.Y(n_1032)
);

OAI321xp33_ASAP7_75t_L g1033 ( 
.A1(n_794),
.A2(n_6),
.A3(n_9),
.B1(n_11),
.B2(n_13),
.C(n_16),
.Y(n_1033)
);

INVx5_ASAP7_75t_L g1034 ( 
.A(n_951),
.Y(n_1034)
);

INVx4_ASAP7_75t_L g1035 ( 
.A(n_951),
.Y(n_1035)
);

AOI21x1_ASAP7_75t_L g1036 ( 
.A1(n_925),
.A2(n_801),
.B(n_844),
.Y(n_1036)
);

INVx2_ASAP7_75t_L g1037 ( 
.A(n_1023),
.Y(n_1037)
);

A2O1A1Ixp33_ASAP7_75t_L g1038 ( 
.A1(n_857),
.A2(n_850),
.B(n_973),
.C(n_993),
.Y(n_1038)
);

NOR2xp33_ASAP7_75t_R g1039 ( 
.A(n_855),
.B(n_764),
.Y(n_1039)
);

INVx1_ASAP7_75t_L g1040 ( 
.A(n_849),
.Y(n_1040)
);

BUFx2_ASAP7_75t_L g1041 ( 
.A(n_856),
.Y(n_1041)
);

NAND2xp5_ASAP7_75t_L g1042 ( 
.A(n_868),
.B(n_792),
.Y(n_1042)
);

AOI21xp5_ASAP7_75t_L g1043 ( 
.A1(n_901),
.A2(n_808),
.B(n_791),
.Y(n_1043)
);

O2A1O1Ixp33_ASAP7_75t_L g1044 ( 
.A1(n_969),
.A2(n_837),
.B(n_760),
.C(n_761),
.Y(n_1044)
);

INVx1_ASAP7_75t_SL g1045 ( 
.A(n_865),
.Y(n_1045)
);

BUFx3_ASAP7_75t_L g1046 ( 
.A(n_961),
.Y(n_1046)
);

AND2x4_ASAP7_75t_SL g1047 ( 
.A(n_957),
.B(n_695),
.Y(n_1047)
);

AOI21xp5_ASAP7_75t_L g1048 ( 
.A1(n_960),
.A2(n_771),
.B(n_773),
.Y(n_1048)
);

OA22x2_ASAP7_75t_L g1049 ( 
.A1(n_893),
.A2(n_764),
.B1(n_297),
.B2(n_718),
.Y(n_1049)
);

O2A1O1Ixp33_ASAP7_75t_L g1050 ( 
.A1(n_969),
.A2(n_806),
.B(n_804),
.C(n_713),
.Y(n_1050)
);

AOI221x1_ASAP7_75t_L g1051 ( 
.A1(n_1032),
.A2(n_722),
.B1(n_718),
.B2(n_713),
.C(n_818),
.Y(n_1051)
);

NOR2xp33_ASAP7_75t_L g1052 ( 
.A(n_1000),
.B(n_722),
.Y(n_1052)
);

A2O1A1Ixp33_ASAP7_75t_L g1053 ( 
.A1(n_993),
.A2(n_1011),
.B(n_1018),
.C(n_992),
.Y(n_1053)
);

BUFx6f_ASAP7_75t_L g1054 ( 
.A(n_951),
.Y(n_1054)
);

OAI21xp33_ASAP7_75t_SL g1055 ( 
.A1(n_923),
.A2(n_878),
.B(n_982),
.Y(n_1055)
);

A2O1A1Ixp33_ASAP7_75t_L g1056 ( 
.A1(n_1011),
.A2(n_1018),
.B(n_992),
.C(n_936),
.Y(n_1056)
);

NAND2xp5_ASAP7_75t_L g1057 ( 
.A(n_898),
.B(n_825),
.Y(n_1057)
);

HB1xp67_ASAP7_75t_L g1058 ( 
.A(n_950),
.Y(n_1058)
);

INVx4_ASAP7_75t_L g1059 ( 
.A(n_951),
.Y(n_1059)
);

NOR2xp33_ASAP7_75t_L g1060 ( 
.A(n_892),
.B(n_824),
.Y(n_1060)
);

NOR2xp33_ASAP7_75t_L g1061 ( 
.A(n_997),
.B(n_820),
.Y(n_1061)
);

INVx1_ASAP7_75t_SL g1062 ( 
.A(n_953),
.Y(n_1062)
);

A2O1A1Ixp33_ASAP7_75t_L g1063 ( 
.A1(n_936),
.A2(n_818),
.B(n_817),
.C(n_802),
.Y(n_1063)
);

INVx2_ASAP7_75t_L g1064 ( 
.A(n_1022),
.Y(n_1064)
);

NAND2x1p5_ASAP7_75t_L g1065 ( 
.A(n_974),
.B(n_817),
.Y(n_1065)
);

OAI22x1_ASAP7_75t_L g1066 ( 
.A1(n_943),
.A2(n_802),
.B1(n_20),
.B2(n_25),
.Y(n_1066)
);

AOI21xp5_ASAP7_75t_L g1067 ( 
.A1(n_873),
.A2(n_657),
.B(n_796),
.Y(n_1067)
);

NAND2xp5_ASAP7_75t_SL g1068 ( 
.A(n_1014),
.B(n_173),
.Y(n_1068)
);

OAI22xp5_ASAP7_75t_L g1069 ( 
.A1(n_1014),
.A2(n_17),
.B1(n_20),
.B2(n_25),
.Y(n_1069)
);

AOI21xp5_ASAP7_75t_L g1070 ( 
.A1(n_875),
.A2(n_165),
.B(n_163),
.Y(n_1070)
);

INVxp67_ASAP7_75t_L g1071 ( 
.A(n_882),
.Y(n_1071)
);

BUFx3_ASAP7_75t_L g1072 ( 
.A(n_961),
.Y(n_1072)
);

NOR2xp33_ASAP7_75t_L g1073 ( 
.A(n_943),
.B(n_27),
.Y(n_1073)
);

BUFx6f_ASAP7_75t_L g1074 ( 
.A(n_974),
.Y(n_1074)
);

INVx1_ASAP7_75t_L g1075 ( 
.A(n_887),
.Y(n_1075)
);

NAND2xp5_ASAP7_75t_SL g1076 ( 
.A(n_908),
.B(n_161),
.Y(n_1076)
);

AND2x2_ASAP7_75t_L g1077 ( 
.A(n_854),
.B(n_27),
.Y(n_1077)
);

INVx1_ASAP7_75t_L g1078 ( 
.A(n_889),
.Y(n_1078)
);

AOI33xp33_ASAP7_75t_L g1079 ( 
.A1(n_964),
.A2(n_34),
.A3(n_35),
.B1(n_37),
.B2(n_41),
.B3(n_42),
.Y(n_1079)
);

INVx1_ASAP7_75t_L g1080 ( 
.A(n_895),
.Y(n_1080)
);

NAND2xp5_ASAP7_75t_L g1081 ( 
.A(n_956),
.B(n_34),
.Y(n_1081)
);

INVx2_ASAP7_75t_L g1082 ( 
.A(n_1022),
.Y(n_1082)
);

INVx1_ASAP7_75t_L g1083 ( 
.A(n_848),
.Y(n_1083)
);

INVx1_ASAP7_75t_L g1084 ( 
.A(n_852),
.Y(n_1084)
);

AOI21xp5_ASAP7_75t_L g1085 ( 
.A1(n_902),
.A2(n_158),
.B(n_139),
.Y(n_1085)
);

NAND2x1p5_ASAP7_75t_L g1086 ( 
.A(n_974),
.B(n_995),
.Y(n_1086)
);

NOR3xp33_ASAP7_75t_L g1087 ( 
.A(n_975),
.B(n_37),
.C(n_43),
.Y(n_1087)
);

AOI21xp5_ASAP7_75t_L g1088 ( 
.A1(n_927),
.A2(n_134),
.B(n_129),
.Y(n_1088)
);

BUFx6f_ASAP7_75t_L g1089 ( 
.A(n_974),
.Y(n_1089)
);

AOI21xp5_ASAP7_75t_L g1090 ( 
.A1(n_944),
.A2(n_128),
.B(n_115),
.Y(n_1090)
);

INVx1_ASAP7_75t_L g1091 ( 
.A(n_900),
.Y(n_1091)
);

NOR2xp33_ASAP7_75t_L g1092 ( 
.A(n_896),
.B(n_975),
.Y(n_1092)
);

INVx1_ASAP7_75t_L g1093 ( 
.A(n_906),
.Y(n_1093)
);

O2A1O1Ixp33_ASAP7_75t_L g1094 ( 
.A1(n_931),
.A2(n_45),
.B(n_46),
.C(n_47),
.Y(n_1094)
);

NAND2xp5_ASAP7_75t_L g1095 ( 
.A(n_937),
.B(n_890),
.Y(n_1095)
);

NOR2xp33_ASAP7_75t_L g1096 ( 
.A(n_998),
.B(n_46),
.Y(n_1096)
);

AOI33xp33_ASAP7_75t_L g1097 ( 
.A1(n_964),
.A2(n_47),
.A3(n_48),
.B1(n_50),
.B2(n_51),
.B3(n_53),
.Y(n_1097)
);

CKINVDCx5p33_ASAP7_75t_R g1098 ( 
.A(n_909),
.Y(n_1098)
);

BUFx6f_ASAP7_75t_L g1099 ( 
.A(n_934),
.Y(n_1099)
);

NAND2xp5_ASAP7_75t_SL g1100 ( 
.A(n_937),
.B(n_114),
.Y(n_1100)
);

BUFx4f_ASAP7_75t_L g1101 ( 
.A(n_912),
.Y(n_1101)
);

BUFx6f_ASAP7_75t_L g1102 ( 
.A(n_942),
.Y(n_1102)
);

NAND2xp5_ASAP7_75t_L g1103 ( 
.A(n_890),
.B(n_894),
.Y(n_1103)
);

AOI21xp5_ASAP7_75t_L g1104 ( 
.A1(n_891),
.A2(n_110),
.B(n_93),
.Y(n_1104)
);

OR2x6_ASAP7_75t_SL g1105 ( 
.A(n_1001),
.B(n_51),
.Y(n_1105)
);

INVx1_ASAP7_75t_L g1106 ( 
.A(n_913),
.Y(n_1106)
);

O2A1O1Ixp33_ASAP7_75t_L g1107 ( 
.A1(n_931),
.A2(n_53),
.B(n_54),
.C(n_55),
.Y(n_1107)
);

INVx1_ASAP7_75t_L g1108 ( 
.A(n_919),
.Y(n_1108)
);

NAND2xp5_ASAP7_75t_L g1109 ( 
.A(n_894),
.B(n_54),
.Y(n_1109)
);

NOR2xp33_ASAP7_75t_R g1110 ( 
.A(n_1031),
.B(n_72),
.Y(n_1110)
);

A2O1A1Ixp33_ASAP7_75t_L g1111 ( 
.A1(n_998),
.A2(n_57),
.B(n_61),
.C(n_79),
.Y(n_1111)
);

NOR2xp67_ASAP7_75t_L g1112 ( 
.A(n_1006),
.B(n_57),
.Y(n_1112)
);

OAI22xp5_ASAP7_75t_L g1113 ( 
.A1(n_876),
.A2(n_1020),
.B1(n_862),
.B2(n_861),
.Y(n_1113)
);

INVx8_ASAP7_75t_L g1114 ( 
.A(n_883),
.Y(n_1114)
);

AOI21xp5_ASAP7_75t_L g1115 ( 
.A1(n_880),
.A2(n_884),
.B(n_869),
.Y(n_1115)
);

NAND2xp5_ASAP7_75t_L g1116 ( 
.A(n_1016),
.B(n_863),
.Y(n_1116)
);

OAI22xp5_ASAP7_75t_L g1117 ( 
.A1(n_876),
.A2(n_995),
.B1(n_918),
.B2(n_945),
.Y(n_1117)
);

INVx1_ASAP7_75t_L g1118 ( 
.A(n_929),
.Y(n_1118)
);

AOI21xp5_ASAP7_75t_L g1119 ( 
.A1(n_904),
.A2(n_851),
.B(n_905),
.Y(n_1119)
);

NAND2xp5_ASAP7_75t_SL g1120 ( 
.A(n_942),
.B(n_980),
.Y(n_1120)
);

O2A1O1Ixp33_ASAP7_75t_L g1121 ( 
.A1(n_945),
.A2(n_999),
.B(n_994),
.C(n_1002),
.Y(n_1121)
);

NOR2xp33_ASAP7_75t_R g1122 ( 
.A(n_1031),
.B(n_917),
.Y(n_1122)
);

BUFx12f_ASAP7_75t_L g1123 ( 
.A(n_926),
.Y(n_1123)
);

INVx1_ASAP7_75t_SL g1124 ( 
.A(n_971),
.Y(n_1124)
);

BUFx6f_ASAP7_75t_L g1125 ( 
.A(n_980),
.Y(n_1125)
);

AO32x1_ASAP7_75t_L g1126 ( 
.A1(n_991),
.A2(n_928),
.A3(n_963),
.B1(n_988),
.B2(n_1017),
.Y(n_1126)
);

NOR3xp33_ASAP7_75t_L g1127 ( 
.A(n_933),
.B(n_866),
.C(n_932),
.Y(n_1127)
);

NAND2xp5_ASAP7_75t_L g1128 ( 
.A(n_938),
.B(n_949),
.Y(n_1128)
);

INVx1_ASAP7_75t_L g1129 ( 
.A(n_959),
.Y(n_1129)
);

OAI22xp5_ASAP7_75t_SL g1130 ( 
.A1(n_1010),
.A2(n_978),
.B1(n_911),
.B2(n_1033),
.Y(n_1130)
);

NOR2xp33_ASAP7_75t_L g1131 ( 
.A(n_897),
.B(n_954),
.Y(n_1131)
);

BUFx3_ASAP7_75t_L g1132 ( 
.A(n_1010),
.Y(n_1132)
);

OAI22xp5_ASAP7_75t_L g1133 ( 
.A1(n_918),
.A2(n_883),
.B1(n_874),
.B2(n_1002),
.Y(n_1133)
);

NAND2xp5_ASAP7_75t_SL g1134 ( 
.A(n_948),
.B(n_986),
.Y(n_1134)
);

BUFx6f_ASAP7_75t_L g1135 ( 
.A(n_883),
.Y(n_1135)
);

A2O1A1Ixp33_ASAP7_75t_L g1136 ( 
.A1(n_1024),
.A2(n_981),
.B(n_1015),
.C(n_1012),
.Y(n_1136)
);

NAND2xp5_ASAP7_75t_L g1137 ( 
.A(n_1024),
.B(n_948),
.Y(n_1137)
);

INVx5_ASAP7_75t_L g1138 ( 
.A(n_847),
.Y(n_1138)
);

INVx2_ASAP7_75t_L g1139 ( 
.A(n_966),
.Y(n_1139)
);

NAND2xp5_ASAP7_75t_SL g1140 ( 
.A(n_986),
.B(n_1013),
.Y(n_1140)
);

NAND2xp5_ASAP7_75t_SL g1141 ( 
.A(n_1008),
.B(n_1009),
.Y(n_1141)
);

O2A1O1Ixp33_ASAP7_75t_L g1142 ( 
.A1(n_994),
.A2(n_1032),
.B(n_1025),
.C(n_1012),
.Y(n_1142)
);

AND2x4_ASAP7_75t_L g1143 ( 
.A(n_899),
.B(n_847),
.Y(n_1143)
);

INVx1_ASAP7_75t_L g1144 ( 
.A(n_907),
.Y(n_1144)
);

AOI21xp5_ASAP7_75t_L g1145 ( 
.A1(n_930),
.A2(n_886),
.B(n_888),
.Y(n_1145)
);

BUFx6f_ASAP7_75t_L g1146 ( 
.A(n_940),
.Y(n_1146)
);

O2A1O1Ixp33_ASAP7_75t_L g1147 ( 
.A1(n_1015),
.A2(n_1025),
.B(n_1007),
.C(n_1030),
.Y(n_1147)
);

AND2x4_ASAP7_75t_L g1148 ( 
.A(n_899),
.B(n_940),
.Y(n_1148)
);

BUFx6f_ASAP7_75t_L g1149 ( 
.A(n_976),
.Y(n_1149)
);

AOI22xp33_ASAP7_75t_L g1150 ( 
.A1(n_1021),
.A2(n_1027),
.B1(n_872),
.B2(n_903),
.Y(n_1150)
);

NOR2xp33_ASAP7_75t_L g1151 ( 
.A(n_925),
.B(n_921),
.Y(n_1151)
);

NAND2xp5_ASAP7_75t_L g1152 ( 
.A(n_914),
.B(n_924),
.Y(n_1152)
);

INVx2_ASAP7_75t_L g1153 ( 
.A(n_1026),
.Y(n_1153)
);

NOR2xp33_ASAP7_75t_L g1154 ( 
.A(n_916),
.B(n_922),
.Y(n_1154)
);

BUFx2_ASAP7_75t_L g1155 ( 
.A(n_979),
.Y(n_1155)
);

INVx1_ASAP7_75t_L g1156 ( 
.A(n_920),
.Y(n_1156)
);

A2O1A1Ixp33_ASAP7_75t_L g1157 ( 
.A1(n_965),
.A2(n_970),
.B(n_881),
.C(n_860),
.Y(n_1157)
);

CKINVDCx16_ASAP7_75t_R g1158 ( 
.A(n_979),
.Y(n_1158)
);

NOR2xp33_ASAP7_75t_R g1159 ( 
.A(n_939),
.B(n_879),
.Y(n_1159)
);

INVx3_ASAP7_75t_SL g1160 ( 
.A(n_952),
.Y(n_1160)
);

AOI21xp5_ASAP7_75t_L g1161 ( 
.A1(n_859),
.A2(n_870),
.B(n_867),
.Y(n_1161)
);

NAND2xp5_ASAP7_75t_L g1162 ( 
.A(n_984),
.B(n_989),
.Y(n_1162)
);

O2A1O1Ixp33_ASAP7_75t_L g1163 ( 
.A1(n_1004),
.A2(n_990),
.B(n_1003),
.C(n_968),
.Y(n_1163)
);

INVx2_ASAP7_75t_L g1164 ( 
.A(n_972),
.Y(n_1164)
);

NAND2xp5_ASAP7_75t_L g1165 ( 
.A(n_885),
.B(n_952),
.Y(n_1165)
);

NAND2xp5_ASAP7_75t_L g1166 ( 
.A(n_976),
.B(n_985),
.Y(n_1166)
);

NAND2xp5_ASAP7_75t_L g1167 ( 
.A(n_985),
.B(n_958),
.Y(n_1167)
);

NOR2xp33_ASAP7_75t_L g1168 ( 
.A(n_983),
.B(n_870),
.Y(n_1168)
);

AND2x2_ASAP7_75t_SL g1169 ( 
.A(n_859),
.B(n_871),
.Y(n_1169)
);

INVx1_ASAP7_75t_L g1170 ( 
.A(n_983),
.Y(n_1170)
);

INVx1_ASAP7_75t_L g1171 ( 
.A(n_935),
.Y(n_1171)
);

AOI22xp5_ASAP7_75t_L g1172 ( 
.A1(n_935),
.A2(n_946),
.B1(n_941),
.B2(n_867),
.Y(n_1172)
);

O2A1O1Ixp33_ASAP7_75t_L g1173 ( 
.A1(n_987),
.A2(n_946),
.B(n_941),
.C(n_871),
.Y(n_1173)
);

INVx2_ASAP7_75t_L g1174 ( 
.A(n_967),
.Y(n_1174)
);

AO21x1_ASAP7_75t_L g1175 ( 
.A1(n_977),
.A2(n_915),
.B(n_910),
.Y(n_1175)
);

NAND2xp5_ASAP7_75t_L g1176 ( 
.A(n_1005),
.B(n_1019),
.Y(n_1176)
);

CKINVDCx8_ASAP7_75t_R g1177 ( 
.A(n_1029),
.Y(n_1177)
);

NAND2xp5_ASAP7_75t_SL g1178 ( 
.A(n_1028),
.B(n_877),
.Y(n_1178)
);

NAND2xp5_ASAP7_75t_L g1179 ( 
.A(n_877),
.B(n_1029),
.Y(n_1179)
);

NAND2xp5_ASAP7_75t_SL g1180 ( 
.A(n_996),
.B(n_955),
.Y(n_1180)
);

A2O1A1Ixp33_ASAP7_75t_L g1181 ( 
.A1(n_962),
.A2(n_853),
.B(n_947),
.C(n_864),
.Y(n_1181)
);

NAND2xp5_ASAP7_75t_L g1182 ( 
.A(n_1029),
.B(n_858),
.Y(n_1182)
);

BUFx2_ASAP7_75t_L g1183 ( 
.A(n_856),
.Y(n_1183)
);

CKINVDCx11_ASAP7_75t_R g1184 ( 
.A(n_926),
.Y(n_1184)
);

INVx1_ASAP7_75t_SL g1185 ( 
.A(n_856),
.Y(n_1185)
);

AOI21xp5_ASAP7_75t_L g1186 ( 
.A1(n_1119),
.A2(n_1115),
.B(n_1152),
.Y(n_1186)
);

OA21x2_ASAP7_75t_L g1187 ( 
.A1(n_1051),
.A2(n_1157),
.B(n_1038),
.Y(n_1187)
);

INVxp67_ASAP7_75t_SL g1188 ( 
.A(n_1058),
.Y(n_1188)
);

O2A1O1Ixp33_ASAP7_75t_SL g1189 ( 
.A1(n_1053),
.A2(n_1056),
.B(n_1136),
.C(n_1096),
.Y(n_1189)
);

INVx4_ASAP7_75t_SL g1190 ( 
.A(n_1123),
.Y(n_1190)
);

OA21x2_ASAP7_75t_L g1191 ( 
.A1(n_1150),
.A2(n_1174),
.B(n_1175),
.Y(n_1191)
);

AOI21xp5_ASAP7_75t_L g1192 ( 
.A1(n_1180),
.A2(n_1128),
.B(n_1043),
.Y(n_1192)
);

INVx1_ASAP7_75t_L g1193 ( 
.A(n_1040),
.Y(n_1193)
);

AO31x2_ASAP7_75t_L g1194 ( 
.A1(n_1113),
.A2(n_1117),
.A3(n_1181),
.B(n_1133),
.Y(n_1194)
);

O2A1O1Ixp33_ASAP7_75t_L g1195 ( 
.A1(n_1073),
.A2(n_1111),
.B(n_1087),
.C(n_1069),
.Y(n_1195)
);

INVx2_ASAP7_75t_L g1196 ( 
.A(n_1037),
.Y(n_1196)
);

AND2x2_ASAP7_75t_L g1197 ( 
.A(n_1131),
.B(n_1124),
.Y(n_1197)
);

NAND2xp5_ASAP7_75t_L g1198 ( 
.A(n_1144),
.B(n_1156),
.Y(n_1198)
);

BUFx6f_ASAP7_75t_L g1199 ( 
.A(n_1099),
.Y(n_1199)
);

AO32x2_ASAP7_75t_L g1200 ( 
.A1(n_1117),
.A2(n_1113),
.A3(n_1130),
.B1(n_1133),
.B2(n_1069),
.Y(n_1200)
);

NAND2xp5_ASAP7_75t_L g1201 ( 
.A(n_1154),
.B(n_1116),
.Y(n_1201)
);

CKINVDCx5p33_ASAP7_75t_R g1202 ( 
.A(n_1098),
.Y(n_1202)
);

NAND2xp5_ASAP7_75t_L g1203 ( 
.A(n_1137),
.B(n_1052),
.Y(n_1203)
);

OAI21x1_ASAP7_75t_L g1204 ( 
.A1(n_1145),
.A2(n_1036),
.B(n_1161),
.Y(n_1204)
);

O2A1O1Ixp33_ASAP7_75t_SL g1205 ( 
.A1(n_1100),
.A2(n_1068),
.B(n_1179),
.C(n_1076),
.Y(n_1205)
);

OAI21xp33_ASAP7_75t_L g1206 ( 
.A1(n_1092),
.A2(n_1079),
.B(n_1097),
.Y(n_1206)
);

OAI21x1_ASAP7_75t_L g1207 ( 
.A1(n_1048),
.A2(n_1067),
.B(n_1173),
.Y(n_1207)
);

AO31x2_ASAP7_75t_L g1208 ( 
.A1(n_1063),
.A2(n_1182),
.A3(n_1168),
.B(n_1151),
.Y(n_1208)
);

OAI22xp5_ASAP7_75t_L g1209 ( 
.A1(n_1177),
.A2(n_1103),
.B1(n_1095),
.B2(n_1078),
.Y(n_1209)
);

CKINVDCx6p67_ASAP7_75t_R g1210 ( 
.A(n_1046),
.Y(n_1210)
);

AO31x2_ASAP7_75t_L g1211 ( 
.A1(n_1176),
.A2(n_1070),
.A3(n_1088),
.B(n_1090),
.Y(n_1211)
);

BUFx6f_ASAP7_75t_L g1212 ( 
.A(n_1099),
.Y(n_1212)
);

AOI21x1_ASAP7_75t_L g1213 ( 
.A1(n_1178),
.A2(n_1162),
.B(n_1081),
.Y(n_1213)
);

AND2x4_ASAP7_75t_L g1214 ( 
.A(n_1135),
.B(n_1099),
.Y(n_1214)
);

BUFx2_ASAP7_75t_L g1215 ( 
.A(n_1041),
.Y(n_1215)
);

AO31x2_ASAP7_75t_L g1216 ( 
.A1(n_1066),
.A2(n_1109),
.A3(n_1165),
.B(n_1171),
.Y(n_1216)
);

AO31x2_ASAP7_75t_L g1217 ( 
.A1(n_1165),
.A2(n_1166),
.A3(n_1170),
.B(n_1167),
.Y(n_1217)
);

O2A1O1Ixp33_ASAP7_75t_L g1218 ( 
.A1(n_1141),
.A2(n_1121),
.B(n_1094),
.C(n_1107),
.Y(n_1218)
);

AOI21xp5_ASAP7_75t_L g1219 ( 
.A1(n_1055),
.A2(n_1163),
.B(n_1147),
.Y(n_1219)
);

NAND2xp5_ASAP7_75t_L g1220 ( 
.A(n_1164),
.B(n_1061),
.Y(n_1220)
);

BUFx12f_ASAP7_75t_L g1221 ( 
.A(n_1184),
.Y(n_1221)
);

AOI21xp5_ASAP7_75t_L g1222 ( 
.A1(n_1042),
.A2(n_1140),
.B(n_1057),
.Y(n_1222)
);

INVx1_ASAP7_75t_L g1223 ( 
.A(n_1075),
.Y(n_1223)
);

HB1xp67_ASAP7_75t_L g1224 ( 
.A(n_1045),
.Y(n_1224)
);

INVx1_ASAP7_75t_L g1225 ( 
.A(n_1080),
.Y(n_1225)
);

INVx2_ASAP7_75t_SL g1226 ( 
.A(n_1101),
.Y(n_1226)
);

AOI21xp5_ASAP7_75t_L g1227 ( 
.A1(n_1044),
.A2(n_1153),
.B(n_1050),
.Y(n_1227)
);

AND2x2_ASAP7_75t_L g1228 ( 
.A(n_1124),
.B(n_1077),
.Y(n_1228)
);

CKINVDCx6p67_ASAP7_75t_R g1229 ( 
.A(n_1072),
.Y(n_1229)
);

OA21x2_ASAP7_75t_L g1230 ( 
.A1(n_1172),
.A2(n_1104),
.B(n_1085),
.Y(n_1230)
);

NAND2xp5_ASAP7_75t_L g1231 ( 
.A(n_1060),
.B(n_1185),
.Y(n_1231)
);

O2A1O1Ixp33_ASAP7_75t_L g1232 ( 
.A1(n_1142),
.A2(n_1127),
.B(n_1071),
.C(n_1062),
.Y(n_1232)
);

CKINVDCx11_ASAP7_75t_R g1233 ( 
.A(n_1105),
.Y(n_1233)
);

AOI22xp33_ASAP7_75t_L g1234 ( 
.A1(n_1130),
.A2(n_1114),
.B1(n_1112),
.B2(n_1135),
.Y(n_1234)
);

OAI21x1_ASAP7_75t_L g1235 ( 
.A1(n_1065),
.A2(n_1086),
.B(n_1172),
.Y(n_1235)
);

INVx2_ASAP7_75t_SL g1236 ( 
.A(n_1101),
.Y(n_1236)
);

OAI21xp5_ASAP7_75t_L g1237 ( 
.A1(n_1169),
.A2(n_1083),
.B(n_1118),
.Y(n_1237)
);

BUFx3_ASAP7_75t_L g1238 ( 
.A(n_1183),
.Y(n_1238)
);

BUFx8_ASAP7_75t_SL g1239 ( 
.A(n_1155),
.Y(n_1239)
);

INVx4_ASAP7_75t_L g1240 ( 
.A(n_1034),
.Y(n_1240)
);

OAI21x1_ASAP7_75t_L g1241 ( 
.A1(n_1065),
.A2(n_1086),
.B(n_1129),
.Y(n_1241)
);

INVx3_ASAP7_75t_L g1242 ( 
.A(n_1149),
.Y(n_1242)
);

INVxp67_ASAP7_75t_SL g1243 ( 
.A(n_1134),
.Y(n_1243)
);

NOR2xp33_ASAP7_75t_L g1244 ( 
.A(n_1062),
.B(n_1185),
.Y(n_1244)
);

AOI21xp5_ASAP7_75t_L g1245 ( 
.A1(n_1034),
.A2(n_1126),
.B(n_1138),
.Y(n_1245)
);

NAND2xp5_ASAP7_75t_L g1246 ( 
.A(n_1045),
.B(n_1160),
.Y(n_1246)
);

OAI21x1_ASAP7_75t_L g1247 ( 
.A1(n_1084),
.A2(n_1108),
.B(n_1106),
.Y(n_1247)
);

NAND3xp33_ASAP7_75t_L g1248 ( 
.A(n_1091),
.B(n_1093),
.C(n_1120),
.Y(n_1248)
);

O2A1O1Ixp33_ASAP7_75t_L g1249 ( 
.A1(n_1139),
.A2(n_1064),
.B(n_1082),
.C(n_1143),
.Y(n_1249)
);

A2O1A1Ixp33_ASAP7_75t_L g1250 ( 
.A1(n_1143),
.A2(n_1148),
.B(n_1114),
.C(n_1135),
.Y(n_1250)
);

O2A1O1Ixp5_ASAP7_75t_L g1251 ( 
.A1(n_1148),
.A2(n_1035),
.B(n_1059),
.C(n_1126),
.Y(n_1251)
);

AOI21xp5_ASAP7_75t_SL g1252 ( 
.A1(n_1149),
.A2(n_1059),
.B(n_1035),
.Y(n_1252)
);

OAI22xp5_ASAP7_75t_L g1253 ( 
.A1(n_1114),
.A2(n_1034),
.B1(n_1138),
.B2(n_1149),
.Y(n_1253)
);

AO31x2_ASAP7_75t_L g1254 ( 
.A1(n_1126),
.A2(n_1159),
.A3(n_1049),
.B(n_1138),
.Y(n_1254)
);

AOI21xp5_ASAP7_75t_L g1255 ( 
.A1(n_1054),
.A2(n_1089),
.B(n_1074),
.Y(n_1255)
);

A2O1A1Ixp33_ASAP7_75t_L g1256 ( 
.A1(n_1047),
.A2(n_1146),
.B(n_1132),
.C(n_1125),
.Y(n_1256)
);

NAND3x1_ASAP7_75t_L g1257 ( 
.A(n_1039),
.B(n_1158),
.C(n_1110),
.Y(n_1257)
);

AOI21xp5_ASAP7_75t_SL g1258 ( 
.A1(n_1054),
.A2(n_1074),
.B(n_1089),
.Y(n_1258)
);

AOI221x1_ASAP7_75t_L g1259 ( 
.A1(n_1054),
.A2(n_1074),
.B1(n_1089),
.B2(n_1146),
.C(n_1125),
.Y(n_1259)
);

AOI21xp5_ASAP7_75t_L g1260 ( 
.A1(n_1146),
.A2(n_1102),
.B(n_1125),
.Y(n_1260)
);

AOI21xp5_ASAP7_75t_L g1261 ( 
.A1(n_1102),
.A2(n_1119),
.B(n_1115),
.Y(n_1261)
);

OAI22xp5_ASAP7_75t_L g1262 ( 
.A1(n_1102),
.A2(n_1056),
.B1(n_1053),
.B2(n_857),
.Y(n_1262)
);

OAI21xp5_ASAP7_75t_L g1263 ( 
.A1(n_1122),
.A2(n_1056),
.B(n_1053),
.Y(n_1263)
);

BUFx2_ASAP7_75t_L g1264 ( 
.A(n_1041),
.Y(n_1264)
);

AOI21xp5_ASAP7_75t_L g1265 ( 
.A1(n_1119),
.A2(n_1115),
.B(n_1152),
.Y(n_1265)
);

NAND3x1_ASAP7_75t_L g1266 ( 
.A(n_1096),
.B(n_1127),
.C(n_1073),
.Y(n_1266)
);

BUFx2_ASAP7_75t_SL g1267 ( 
.A(n_1185),
.Y(n_1267)
);

AO21x2_ASAP7_75t_L g1268 ( 
.A1(n_1119),
.A2(n_1159),
.B(n_1038),
.Y(n_1268)
);

AO31x2_ASAP7_75t_L g1269 ( 
.A1(n_1051),
.A2(n_1175),
.A3(n_1157),
.B(n_1038),
.Y(n_1269)
);

AO21x2_ASAP7_75t_L g1270 ( 
.A1(n_1119),
.A2(n_1159),
.B(n_1038),
.Y(n_1270)
);

INVxp67_ASAP7_75t_SL g1271 ( 
.A(n_1058),
.Y(n_1271)
);

NOR2xp33_ASAP7_75t_L g1272 ( 
.A(n_1053),
.B(n_857),
.Y(n_1272)
);

BUFx5_ASAP7_75t_L g1273 ( 
.A(n_1169),
.Y(n_1273)
);

AND2x6_ASAP7_75t_L g1274 ( 
.A(n_1149),
.B(n_1135),
.Y(n_1274)
);

OAI21xp5_ASAP7_75t_SL g1275 ( 
.A1(n_1096),
.A2(n_857),
.B(n_776),
.Y(n_1275)
);

NOR2xp33_ASAP7_75t_L g1276 ( 
.A(n_1053),
.B(n_857),
.Y(n_1276)
);

NAND2xp5_ASAP7_75t_L g1277 ( 
.A(n_1131),
.B(n_1056),
.Y(n_1277)
);

A2O1A1Ixp33_ASAP7_75t_L g1278 ( 
.A1(n_1056),
.A2(n_1053),
.B(n_857),
.C(n_1073),
.Y(n_1278)
);

OAI21x1_ASAP7_75t_L g1279 ( 
.A1(n_1145),
.A2(n_977),
.B(n_1119),
.Y(n_1279)
);

AOI21xp5_ASAP7_75t_L g1280 ( 
.A1(n_1119),
.A2(n_1115),
.B(n_1152),
.Y(n_1280)
);

AOI22xp5_ASAP7_75t_L g1281 ( 
.A1(n_1073),
.A2(n_1096),
.B1(n_1056),
.B2(n_1053),
.Y(n_1281)
);

INVx1_ASAP7_75t_L g1282 ( 
.A(n_1040),
.Y(n_1282)
);

AOI21xp5_ASAP7_75t_L g1283 ( 
.A1(n_1119),
.A2(n_1115),
.B(n_1152),
.Y(n_1283)
);

BUFx4f_ASAP7_75t_SL g1284 ( 
.A(n_1123),
.Y(n_1284)
);

OAI21x1_ASAP7_75t_L g1285 ( 
.A1(n_1145),
.A2(n_977),
.B(n_1119),
.Y(n_1285)
);

AOI21xp5_ASAP7_75t_L g1286 ( 
.A1(n_1119),
.A2(n_1115),
.B(n_1152),
.Y(n_1286)
);

OAI22xp5_ASAP7_75t_L g1287 ( 
.A1(n_1056),
.A2(n_1053),
.B1(n_751),
.B2(n_1096),
.Y(n_1287)
);

OAI22xp5_ASAP7_75t_L g1288 ( 
.A1(n_1056),
.A2(n_1053),
.B1(n_751),
.B2(n_1096),
.Y(n_1288)
);

OAI22xp5_ASAP7_75t_L g1289 ( 
.A1(n_1056),
.A2(n_1053),
.B1(n_751),
.B2(n_1096),
.Y(n_1289)
);

AOI21xp5_ASAP7_75t_SL g1290 ( 
.A1(n_1056),
.A2(n_1053),
.B(n_1038),
.Y(n_1290)
);

INVx1_ASAP7_75t_L g1291 ( 
.A(n_1040),
.Y(n_1291)
);

OAI21x1_ASAP7_75t_L g1292 ( 
.A1(n_1145),
.A2(n_977),
.B(n_1119),
.Y(n_1292)
);

BUFx2_ASAP7_75t_L g1293 ( 
.A(n_1041),
.Y(n_1293)
);

OAI21x1_ASAP7_75t_L g1294 ( 
.A1(n_1145),
.A2(n_977),
.B(n_1119),
.Y(n_1294)
);

OAI22x1_ASAP7_75t_L g1295 ( 
.A1(n_1096),
.A2(n_1073),
.B1(n_943),
.B2(n_998),
.Y(n_1295)
);

NAND2xp5_ASAP7_75t_L g1296 ( 
.A(n_1131),
.B(n_1056),
.Y(n_1296)
);

AND2x4_ASAP7_75t_L g1297 ( 
.A(n_1135),
.B(n_934),
.Y(n_1297)
);

OAI22xp5_ASAP7_75t_L g1298 ( 
.A1(n_1056),
.A2(n_1053),
.B1(n_751),
.B2(n_1096),
.Y(n_1298)
);

AOI21xp5_ASAP7_75t_L g1299 ( 
.A1(n_1119),
.A2(n_1115),
.B(n_1152),
.Y(n_1299)
);

OA21x2_ASAP7_75t_L g1300 ( 
.A1(n_1051),
.A2(n_1157),
.B(n_1119),
.Y(n_1300)
);

OAI22xp5_ASAP7_75t_L g1301 ( 
.A1(n_1056),
.A2(n_1053),
.B1(n_751),
.B2(n_1096),
.Y(n_1301)
);

A2O1A1Ixp33_ASAP7_75t_L g1302 ( 
.A1(n_1056),
.A2(n_1053),
.B(n_857),
.C(n_1073),
.Y(n_1302)
);

AOI21xp5_ASAP7_75t_L g1303 ( 
.A1(n_1119),
.A2(n_1115),
.B(n_1152),
.Y(n_1303)
);

BUFx2_ASAP7_75t_L g1304 ( 
.A(n_1041),
.Y(n_1304)
);

AOI21xp5_ASAP7_75t_L g1305 ( 
.A1(n_1119),
.A2(n_1115),
.B(n_1152),
.Y(n_1305)
);

AOI22xp5_ASAP7_75t_L g1306 ( 
.A1(n_1073),
.A2(n_1096),
.B1(n_1056),
.B2(n_1053),
.Y(n_1306)
);

OAI21x1_ASAP7_75t_L g1307 ( 
.A1(n_1145),
.A2(n_977),
.B(n_1119),
.Y(n_1307)
);

AND2x4_ASAP7_75t_L g1308 ( 
.A(n_1135),
.B(n_934),
.Y(n_1308)
);

OA21x2_ASAP7_75t_L g1309 ( 
.A1(n_1051),
.A2(n_1157),
.B(n_1119),
.Y(n_1309)
);

INVx2_ASAP7_75t_L g1310 ( 
.A(n_1037),
.Y(n_1310)
);

NAND2xp5_ASAP7_75t_L g1311 ( 
.A(n_1131),
.B(n_1056),
.Y(n_1311)
);

NAND2xp5_ASAP7_75t_L g1312 ( 
.A(n_1131),
.B(n_1056),
.Y(n_1312)
);

BUFx6f_ASAP7_75t_L g1313 ( 
.A(n_1099),
.Y(n_1313)
);

INVxp67_ASAP7_75t_L g1314 ( 
.A(n_1041),
.Y(n_1314)
);

NAND2xp5_ASAP7_75t_L g1315 ( 
.A(n_1131),
.B(n_1056),
.Y(n_1315)
);

NAND2xp5_ASAP7_75t_L g1316 ( 
.A(n_1131),
.B(n_1056),
.Y(n_1316)
);

O2A1O1Ixp5_ASAP7_75t_SL g1317 ( 
.A1(n_1180),
.A2(n_857),
.B(n_1117),
.C(n_1069),
.Y(n_1317)
);

OAI21xp5_ASAP7_75t_L g1318 ( 
.A1(n_1056),
.A2(n_1053),
.B(n_1038),
.Y(n_1318)
);

AOI22xp33_ASAP7_75t_L g1319 ( 
.A1(n_1073),
.A2(n_857),
.B1(n_1096),
.B2(n_943),
.Y(n_1319)
);

OAI21xp5_ASAP7_75t_L g1320 ( 
.A1(n_1056),
.A2(n_1053),
.B(n_1038),
.Y(n_1320)
);

NAND2xp5_ASAP7_75t_L g1321 ( 
.A(n_1131),
.B(n_1056),
.Y(n_1321)
);

O2A1O1Ixp33_ASAP7_75t_SL g1322 ( 
.A1(n_1053),
.A2(n_1056),
.B(n_857),
.C(n_1038),
.Y(n_1322)
);

AOI221xp5_ASAP7_75t_L g1323 ( 
.A1(n_1096),
.A2(n_857),
.B1(n_539),
.B2(n_1073),
.C(n_567),
.Y(n_1323)
);

INVx4_ASAP7_75t_SL g1324 ( 
.A(n_1123),
.Y(n_1324)
);

BUFx12f_ASAP7_75t_L g1325 ( 
.A(n_1184),
.Y(n_1325)
);

BUFx10_ASAP7_75t_L g1326 ( 
.A(n_1092),
.Y(n_1326)
);

OAI22x1_ASAP7_75t_L g1327 ( 
.A1(n_1096),
.A2(n_1073),
.B1(n_943),
.B2(n_998),
.Y(n_1327)
);

AO31x2_ASAP7_75t_L g1328 ( 
.A1(n_1051),
.A2(n_1175),
.A3(n_1157),
.B(n_1038),
.Y(n_1328)
);

OAI22xp5_ASAP7_75t_L g1329 ( 
.A1(n_1056),
.A2(n_1053),
.B1(n_751),
.B2(n_1096),
.Y(n_1329)
);

OAI21xp5_ASAP7_75t_L g1330 ( 
.A1(n_1056),
.A2(n_1053),
.B(n_1038),
.Y(n_1330)
);

BUFx8_ASAP7_75t_SL g1331 ( 
.A(n_1123),
.Y(n_1331)
);

INVxp67_ASAP7_75t_L g1332 ( 
.A(n_1041),
.Y(n_1332)
);

NOR2xp33_ASAP7_75t_L g1333 ( 
.A(n_1053),
.B(n_857),
.Y(n_1333)
);

INVx1_ASAP7_75t_L g1334 ( 
.A(n_1040),
.Y(n_1334)
);

INVx1_ASAP7_75t_L g1335 ( 
.A(n_1040),
.Y(n_1335)
);

AOI21xp5_ASAP7_75t_L g1336 ( 
.A1(n_1119),
.A2(n_1115),
.B(n_1152),
.Y(n_1336)
);

OAI22xp5_ASAP7_75t_L g1337 ( 
.A1(n_1056),
.A2(n_1053),
.B1(n_751),
.B2(n_1096),
.Y(n_1337)
);

OAI22xp33_ASAP7_75t_L g1338 ( 
.A1(n_1281),
.A2(n_1306),
.B1(n_1295),
.B2(n_1327),
.Y(n_1338)
);

HB1xp67_ASAP7_75t_L g1339 ( 
.A(n_1208),
.Y(n_1339)
);

INVx6_ASAP7_75t_L g1340 ( 
.A(n_1199),
.Y(n_1340)
);

CKINVDCx11_ASAP7_75t_R g1341 ( 
.A(n_1221),
.Y(n_1341)
);

BUFx3_ASAP7_75t_L g1342 ( 
.A(n_1238),
.Y(n_1342)
);

BUFx4f_ASAP7_75t_SL g1343 ( 
.A(n_1325),
.Y(n_1343)
);

INVx1_ASAP7_75t_SL g1344 ( 
.A(n_1267),
.Y(n_1344)
);

AOI22xp33_ASAP7_75t_L g1345 ( 
.A1(n_1323),
.A2(n_1319),
.B1(n_1272),
.B2(n_1276),
.Y(n_1345)
);

INVx11_ASAP7_75t_L g1346 ( 
.A(n_1274),
.Y(n_1346)
);

AOI22xp33_ASAP7_75t_L g1347 ( 
.A1(n_1333),
.A2(n_1281),
.B1(n_1306),
.B2(n_1301),
.Y(n_1347)
);

INVx3_ASAP7_75t_L g1348 ( 
.A(n_1199),
.Y(n_1348)
);

OAI22x1_ASAP7_75t_L g1349 ( 
.A1(n_1277),
.A2(n_1316),
.B1(n_1296),
.B2(n_1315),
.Y(n_1349)
);

NAND2xp5_ASAP7_75t_L g1350 ( 
.A(n_1201),
.B(n_1203),
.Y(n_1350)
);

AND2x2_ASAP7_75t_L g1351 ( 
.A(n_1197),
.B(n_1228),
.Y(n_1351)
);

CKINVDCx11_ASAP7_75t_R g1352 ( 
.A(n_1190),
.Y(n_1352)
);

AOI22xp33_ASAP7_75t_L g1353 ( 
.A1(n_1287),
.A2(n_1337),
.B1(n_1329),
.B2(n_1288),
.Y(n_1353)
);

INVx6_ASAP7_75t_L g1354 ( 
.A(n_1199),
.Y(n_1354)
);

AOI22xp33_ASAP7_75t_L g1355 ( 
.A1(n_1287),
.A2(n_1337),
.B1(n_1329),
.B2(n_1288),
.Y(n_1355)
);

CKINVDCx5p33_ASAP7_75t_R g1356 ( 
.A(n_1202),
.Y(n_1356)
);

INVx6_ASAP7_75t_L g1357 ( 
.A(n_1212),
.Y(n_1357)
);

INVx2_ASAP7_75t_L g1358 ( 
.A(n_1193),
.Y(n_1358)
);

CKINVDCx5p33_ASAP7_75t_R g1359 ( 
.A(n_1331),
.Y(n_1359)
);

CKINVDCx11_ASAP7_75t_R g1360 ( 
.A(n_1190),
.Y(n_1360)
);

NAND2xp5_ASAP7_75t_L g1361 ( 
.A(n_1220),
.B(n_1198),
.Y(n_1361)
);

CKINVDCx11_ASAP7_75t_R g1362 ( 
.A(n_1324),
.Y(n_1362)
);

AOI22xp33_ASAP7_75t_L g1363 ( 
.A1(n_1289),
.A2(n_1298),
.B1(n_1301),
.B2(n_1330),
.Y(n_1363)
);

OAI21xp33_ASAP7_75t_L g1364 ( 
.A1(n_1275),
.A2(n_1302),
.B(n_1278),
.Y(n_1364)
);

AOI22xp33_ASAP7_75t_L g1365 ( 
.A1(n_1289),
.A2(n_1298),
.B1(n_1320),
.B2(n_1330),
.Y(n_1365)
);

BUFx3_ASAP7_75t_L g1366 ( 
.A(n_1215),
.Y(n_1366)
);

AOI22xp33_ASAP7_75t_L g1367 ( 
.A1(n_1318),
.A2(n_1320),
.B1(n_1321),
.B2(n_1312),
.Y(n_1367)
);

INVx1_ASAP7_75t_L g1368 ( 
.A(n_1223),
.Y(n_1368)
);

CKINVDCx11_ASAP7_75t_R g1369 ( 
.A(n_1324),
.Y(n_1369)
);

CKINVDCx11_ASAP7_75t_R g1370 ( 
.A(n_1210),
.Y(n_1370)
);

BUFx6f_ASAP7_75t_L g1371 ( 
.A(n_1212),
.Y(n_1371)
);

INVx1_ASAP7_75t_L g1372 ( 
.A(n_1225),
.Y(n_1372)
);

OAI22xp5_ASAP7_75t_L g1373 ( 
.A1(n_1275),
.A2(n_1266),
.B1(n_1311),
.B2(n_1209),
.Y(n_1373)
);

CKINVDCx11_ASAP7_75t_R g1374 ( 
.A(n_1229),
.Y(n_1374)
);

AOI22xp33_ASAP7_75t_SL g1375 ( 
.A1(n_1318),
.A2(n_1263),
.B1(n_1262),
.B2(n_1209),
.Y(n_1375)
);

BUFx8_ASAP7_75t_SL g1376 ( 
.A(n_1239),
.Y(n_1376)
);

OAI21xp5_ASAP7_75t_SL g1377 ( 
.A1(n_1195),
.A2(n_1263),
.B(n_1218),
.Y(n_1377)
);

OAI22xp5_ASAP7_75t_L g1378 ( 
.A1(n_1231),
.A2(n_1234),
.B1(n_1246),
.B2(n_1243),
.Y(n_1378)
);

AOI22xp33_ASAP7_75t_L g1379 ( 
.A1(n_1206),
.A2(n_1219),
.B1(n_1326),
.B2(n_1270),
.Y(n_1379)
);

INVx6_ASAP7_75t_L g1380 ( 
.A(n_1313),
.Y(n_1380)
);

BUFx3_ASAP7_75t_L g1381 ( 
.A(n_1264),
.Y(n_1381)
);

INVx3_ASAP7_75t_L g1382 ( 
.A(n_1313),
.Y(n_1382)
);

BUFx4_ASAP7_75t_SL g1383 ( 
.A(n_1293),
.Y(n_1383)
);

INVx2_ASAP7_75t_L g1384 ( 
.A(n_1282),
.Y(n_1384)
);

AOI22xp33_ASAP7_75t_L g1385 ( 
.A1(n_1206),
.A2(n_1326),
.B1(n_1268),
.B2(n_1270),
.Y(n_1385)
);

INVx6_ASAP7_75t_L g1386 ( 
.A(n_1313),
.Y(n_1386)
);

CKINVDCx11_ASAP7_75t_R g1387 ( 
.A(n_1233),
.Y(n_1387)
);

AOI22xp5_ASAP7_75t_L g1388 ( 
.A1(n_1189),
.A2(n_1322),
.B1(n_1244),
.B2(n_1236),
.Y(n_1388)
);

INVx1_ASAP7_75t_L g1389 ( 
.A(n_1291),
.Y(n_1389)
);

AOI22xp33_ASAP7_75t_L g1390 ( 
.A1(n_1268),
.A2(n_1224),
.B1(n_1237),
.B2(n_1273),
.Y(n_1390)
);

NAND2xp5_ASAP7_75t_L g1391 ( 
.A(n_1188),
.B(n_1271),
.Y(n_1391)
);

BUFx12f_ASAP7_75t_L g1392 ( 
.A(n_1304),
.Y(n_1392)
);

OAI21xp5_ASAP7_75t_SL g1393 ( 
.A1(n_1232),
.A2(n_1227),
.B(n_1250),
.Y(n_1393)
);

AOI22xp33_ASAP7_75t_L g1394 ( 
.A1(n_1237),
.A2(n_1273),
.B1(n_1187),
.B2(n_1222),
.Y(n_1394)
);

AOI22xp33_ASAP7_75t_L g1395 ( 
.A1(n_1273),
.A2(n_1187),
.B1(n_1335),
.B2(n_1334),
.Y(n_1395)
);

AND2x2_ASAP7_75t_L g1396 ( 
.A(n_1297),
.B(n_1308),
.Y(n_1396)
);

BUFx10_ASAP7_75t_L g1397 ( 
.A(n_1214),
.Y(n_1397)
);

CKINVDCx11_ASAP7_75t_R g1398 ( 
.A(n_1284),
.Y(n_1398)
);

INVx2_ASAP7_75t_L g1399 ( 
.A(n_1196),
.Y(n_1399)
);

AOI22xp33_ASAP7_75t_L g1400 ( 
.A1(n_1273),
.A2(n_1230),
.B1(n_1290),
.B2(n_1248),
.Y(n_1400)
);

CKINVDCx11_ASAP7_75t_R g1401 ( 
.A(n_1214),
.Y(n_1401)
);

AOI22xp5_ASAP7_75t_SL g1402 ( 
.A1(n_1226),
.A2(n_1332),
.B1(n_1314),
.B2(n_1297),
.Y(n_1402)
);

BUFx6f_ASAP7_75t_L g1403 ( 
.A(n_1274),
.Y(n_1403)
);

OAI22xp5_ASAP7_75t_L g1404 ( 
.A1(n_1256),
.A2(n_1253),
.B1(n_1257),
.B2(n_1308),
.Y(n_1404)
);

INVx1_ASAP7_75t_L g1405 ( 
.A(n_1310),
.Y(n_1405)
);

INVx1_ASAP7_75t_SL g1406 ( 
.A(n_1242),
.Y(n_1406)
);

AOI22xp5_ASAP7_75t_L g1407 ( 
.A1(n_1205),
.A2(n_1273),
.B1(n_1274),
.B2(n_1253),
.Y(n_1407)
);

INVx1_ASAP7_75t_SL g1408 ( 
.A(n_1242),
.Y(n_1408)
);

AOI22xp5_ASAP7_75t_L g1409 ( 
.A1(n_1274),
.A2(n_1230),
.B1(n_1261),
.B2(n_1260),
.Y(n_1409)
);

AOI22xp33_ASAP7_75t_SL g1410 ( 
.A1(n_1200),
.A2(n_1309),
.B1(n_1300),
.B2(n_1317),
.Y(n_1410)
);

BUFx2_ASAP7_75t_SL g1411 ( 
.A(n_1240),
.Y(n_1411)
);

INVx3_ASAP7_75t_L g1412 ( 
.A(n_1240),
.Y(n_1412)
);

AND2x2_ASAP7_75t_L g1413 ( 
.A(n_1216),
.B(n_1247),
.Y(n_1413)
);

INVx3_ASAP7_75t_L g1414 ( 
.A(n_1241),
.Y(n_1414)
);

BUFx6f_ASAP7_75t_L g1415 ( 
.A(n_1235),
.Y(n_1415)
);

BUFx6f_ASAP7_75t_L g1416 ( 
.A(n_1207),
.Y(n_1416)
);

INVx1_ASAP7_75t_L g1417 ( 
.A(n_1217),
.Y(n_1417)
);

AOI22xp5_ASAP7_75t_L g1418 ( 
.A1(n_1186),
.A2(n_1265),
.B1(n_1305),
.B2(n_1303),
.Y(n_1418)
);

INVx1_ASAP7_75t_L g1419 ( 
.A(n_1217),
.Y(n_1419)
);

BUFx10_ASAP7_75t_L g1420 ( 
.A(n_1258),
.Y(n_1420)
);

OAI22xp5_ASAP7_75t_L g1421 ( 
.A1(n_1249),
.A2(n_1245),
.B1(n_1300),
.B2(n_1309),
.Y(n_1421)
);

INVx1_ASAP7_75t_L g1422 ( 
.A(n_1217),
.Y(n_1422)
);

AOI21xp33_ASAP7_75t_L g1423 ( 
.A1(n_1191),
.A2(n_1336),
.B(n_1299),
.Y(n_1423)
);

NAND2xp33_ASAP7_75t_L g1424 ( 
.A(n_1255),
.B(n_1192),
.Y(n_1424)
);

BUFx8_ASAP7_75t_L g1425 ( 
.A(n_1200),
.Y(n_1425)
);

CKINVDCx14_ASAP7_75t_R g1426 ( 
.A(n_1200),
.Y(n_1426)
);

OAI22xp33_ASAP7_75t_L g1427 ( 
.A1(n_1259),
.A2(n_1213),
.B1(n_1280),
.B2(n_1286),
.Y(n_1427)
);

CKINVDCx11_ASAP7_75t_R g1428 ( 
.A(n_1252),
.Y(n_1428)
);

AND2x2_ASAP7_75t_L g1429 ( 
.A(n_1216),
.B(n_1208),
.Y(n_1429)
);

AOI22xp33_ASAP7_75t_L g1430 ( 
.A1(n_1283),
.A2(n_1194),
.B1(n_1204),
.B2(n_1294),
.Y(n_1430)
);

BUFx2_ASAP7_75t_L g1431 ( 
.A(n_1254),
.Y(n_1431)
);

INVx3_ASAP7_75t_SL g1432 ( 
.A(n_1254),
.Y(n_1432)
);

BUFx3_ASAP7_75t_L g1433 ( 
.A(n_1194),
.Y(n_1433)
);

OAI21xp5_ASAP7_75t_SL g1434 ( 
.A1(n_1194),
.A2(n_1211),
.B(n_1328),
.Y(n_1434)
);

AOI22xp5_ASAP7_75t_L g1435 ( 
.A1(n_1279),
.A2(n_1285),
.B1(n_1292),
.B2(n_1307),
.Y(n_1435)
);

OAI22xp5_ASAP7_75t_L g1436 ( 
.A1(n_1211),
.A2(n_1328),
.B1(n_1269),
.B2(n_1251),
.Y(n_1436)
);

INVx6_ASAP7_75t_L g1437 ( 
.A(n_1269),
.Y(n_1437)
);

CKINVDCx11_ASAP7_75t_R g1438 ( 
.A(n_1221),
.Y(n_1438)
);

AOI22xp33_ASAP7_75t_L g1439 ( 
.A1(n_1323),
.A2(n_1319),
.B1(n_1327),
.B2(n_1295),
.Y(n_1439)
);

AOI22xp33_ASAP7_75t_L g1440 ( 
.A1(n_1323),
.A2(n_1319),
.B1(n_1327),
.B2(n_1295),
.Y(n_1440)
);

CKINVDCx11_ASAP7_75t_R g1441 ( 
.A(n_1221),
.Y(n_1441)
);

BUFx3_ASAP7_75t_L g1442 ( 
.A(n_1238),
.Y(n_1442)
);

CKINVDCx20_ASAP7_75t_R g1443 ( 
.A(n_1331),
.Y(n_1443)
);

INVx6_ASAP7_75t_L g1444 ( 
.A(n_1199),
.Y(n_1444)
);

INVx6_ASAP7_75t_L g1445 ( 
.A(n_1199),
.Y(n_1445)
);

NAND2xp5_ASAP7_75t_L g1446 ( 
.A(n_1201),
.B(n_1203),
.Y(n_1446)
);

INVx6_ASAP7_75t_L g1447 ( 
.A(n_1199),
.Y(n_1447)
);

OAI22xp33_ASAP7_75t_L g1448 ( 
.A1(n_1281),
.A2(n_1306),
.B1(n_1327),
.B2(n_1295),
.Y(n_1448)
);

INVx3_ASAP7_75t_L g1449 ( 
.A(n_1199),
.Y(n_1449)
);

INVx6_ASAP7_75t_L g1450 ( 
.A(n_1199),
.Y(n_1450)
);

AOI22xp33_ASAP7_75t_SL g1451 ( 
.A1(n_1287),
.A2(n_1096),
.B1(n_449),
.B2(n_479),
.Y(n_1451)
);

AOI22xp33_ASAP7_75t_L g1452 ( 
.A1(n_1323),
.A2(n_1319),
.B1(n_1327),
.B2(n_1295),
.Y(n_1452)
);

BUFx2_ASAP7_75t_SL g1453 ( 
.A(n_1226),
.Y(n_1453)
);

BUFx12f_ASAP7_75t_L g1454 ( 
.A(n_1221),
.Y(n_1454)
);

OAI21xp5_ASAP7_75t_SL g1455 ( 
.A1(n_1275),
.A2(n_857),
.B(n_1319),
.Y(n_1455)
);

NAND2xp5_ASAP7_75t_L g1456 ( 
.A(n_1201),
.B(n_1203),
.Y(n_1456)
);

HB1xp67_ASAP7_75t_L g1457 ( 
.A(n_1208),
.Y(n_1457)
);

AOI22xp33_ASAP7_75t_L g1458 ( 
.A1(n_1323),
.A2(n_1319),
.B1(n_1327),
.B2(n_1295),
.Y(n_1458)
);

OAI22xp5_ASAP7_75t_L g1459 ( 
.A1(n_1319),
.A2(n_1306),
.B1(n_1281),
.B2(n_1056),
.Y(n_1459)
);

BUFx12f_ASAP7_75t_L g1460 ( 
.A(n_1221),
.Y(n_1460)
);

BUFx2_ASAP7_75t_SL g1461 ( 
.A(n_1226),
.Y(n_1461)
);

INVx2_ASAP7_75t_SL g1462 ( 
.A(n_1238),
.Y(n_1462)
);

BUFx3_ASAP7_75t_L g1463 ( 
.A(n_1238),
.Y(n_1463)
);

INVx6_ASAP7_75t_L g1464 ( 
.A(n_1199),
.Y(n_1464)
);

CKINVDCx20_ASAP7_75t_R g1465 ( 
.A(n_1331),
.Y(n_1465)
);

NAND2xp5_ASAP7_75t_L g1466 ( 
.A(n_1201),
.B(n_1203),
.Y(n_1466)
);

BUFx12f_ASAP7_75t_L g1467 ( 
.A(n_1221),
.Y(n_1467)
);

INVx6_ASAP7_75t_L g1468 ( 
.A(n_1199),
.Y(n_1468)
);

BUFx2_ASAP7_75t_L g1469 ( 
.A(n_1433),
.Y(n_1469)
);

O2A1O1Ixp5_ASAP7_75t_L g1470 ( 
.A1(n_1459),
.A2(n_1338),
.B(n_1448),
.C(n_1373),
.Y(n_1470)
);

HB1xp67_ASAP7_75t_L g1471 ( 
.A(n_1391),
.Y(n_1471)
);

AND2x4_ASAP7_75t_L g1472 ( 
.A(n_1415),
.B(n_1414),
.Y(n_1472)
);

INVx1_ASAP7_75t_L g1473 ( 
.A(n_1417),
.Y(n_1473)
);

AND2x2_ASAP7_75t_L g1474 ( 
.A(n_1426),
.B(n_1429),
.Y(n_1474)
);

AND2x2_ASAP7_75t_L g1475 ( 
.A(n_1426),
.B(n_1347),
.Y(n_1475)
);

HB1xp67_ASAP7_75t_L g1476 ( 
.A(n_1358),
.Y(n_1476)
);

INVx1_ASAP7_75t_L g1477 ( 
.A(n_1419),
.Y(n_1477)
);

INVx1_ASAP7_75t_L g1478 ( 
.A(n_1422),
.Y(n_1478)
);

INVx1_ASAP7_75t_L g1479 ( 
.A(n_1413),
.Y(n_1479)
);

AND2x2_ASAP7_75t_L g1480 ( 
.A(n_1347),
.B(n_1375),
.Y(n_1480)
);

INVx1_ASAP7_75t_L g1481 ( 
.A(n_1339),
.Y(n_1481)
);

OAI21xp5_ASAP7_75t_L g1482 ( 
.A1(n_1345),
.A2(n_1455),
.B(n_1377),
.Y(n_1482)
);

BUFx2_ASAP7_75t_L g1483 ( 
.A(n_1339),
.Y(n_1483)
);

INVx2_ASAP7_75t_SL g1484 ( 
.A(n_1397),
.Y(n_1484)
);

INVx2_ASAP7_75t_L g1485 ( 
.A(n_1384),
.Y(n_1485)
);

INVx1_ASAP7_75t_L g1486 ( 
.A(n_1457),
.Y(n_1486)
);

OR2x2_ASAP7_75t_L g1487 ( 
.A(n_1457),
.B(n_1434),
.Y(n_1487)
);

OAI21x1_ASAP7_75t_L g1488 ( 
.A1(n_1430),
.A2(n_1435),
.B(n_1414),
.Y(n_1488)
);

INVx2_ASAP7_75t_L g1489 ( 
.A(n_1437),
.Y(n_1489)
);

INVxp67_ASAP7_75t_SL g1490 ( 
.A(n_1361),
.Y(n_1490)
);

INVxp67_ASAP7_75t_L g1491 ( 
.A(n_1351),
.Y(n_1491)
);

AND2x4_ASAP7_75t_L g1492 ( 
.A(n_1409),
.B(n_1416),
.Y(n_1492)
);

NAND2xp5_ASAP7_75t_L g1493 ( 
.A(n_1350),
.B(n_1446),
.Y(n_1493)
);

INVx1_ASAP7_75t_L g1494 ( 
.A(n_1431),
.Y(n_1494)
);

INVx1_ASAP7_75t_L g1495 ( 
.A(n_1436),
.Y(n_1495)
);

BUFx3_ASAP7_75t_L g1496 ( 
.A(n_1428),
.Y(n_1496)
);

NOR2xp33_ASAP7_75t_L g1497 ( 
.A(n_1456),
.B(n_1466),
.Y(n_1497)
);

INVx1_ASAP7_75t_L g1498 ( 
.A(n_1368),
.Y(n_1498)
);

INVx1_ASAP7_75t_L g1499 ( 
.A(n_1372),
.Y(n_1499)
);

INVx1_ASAP7_75t_L g1500 ( 
.A(n_1389),
.Y(n_1500)
);

AND2x2_ASAP7_75t_L g1501 ( 
.A(n_1375),
.B(n_1353),
.Y(n_1501)
);

AOI22xp33_ASAP7_75t_L g1502 ( 
.A1(n_1345),
.A2(n_1451),
.B1(n_1364),
.B2(n_1452),
.Y(n_1502)
);

AND2x4_ASAP7_75t_L g1503 ( 
.A(n_1416),
.B(n_1400),
.Y(n_1503)
);

OAI21x1_ASAP7_75t_L g1504 ( 
.A1(n_1430),
.A2(n_1418),
.B(n_1421),
.Y(n_1504)
);

AND2x2_ASAP7_75t_L g1505 ( 
.A(n_1353),
.B(n_1355),
.Y(n_1505)
);

BUFx2_ASAP7_75t_L g1506 ( 
.A(n_1425),
.Y(n_1506)
);

INVx2_ASAP7_75t_SL g1507 ( 
.A(n_1397),
.Y(n_1507)
);

OAI21x1_ASAP7_75t_L g1508 ( 
.A1(n_1400),
.A2(n_1394),
.B(n_1355),
.Y(n_1508)
);

INVx1_ASAP7_75t_L g1509 ( 
.A(n_1432),
.Y(n_1509)
);

INVx1_ASAP7_75t_L g1510 ( 
.A(n_1349),
.Y(n_1510)
);

INVx2_ASAP7_75t_SL g1511 ( 
.A(n_1340),
.Y(n_1511)
);

AOI22xp33_ASAP7_75t_SL g1512 ( 
.A1(n_1425),
.A2(n_1451),
.B1(n_1402),
.B2(n_1378),
.Y(n_1512)
);

INVx1_ASAP7_75t_L g1513 ( 
.A(n_1410),
.Y(n_1513)
);

BUFx3_ASAP7_75t_L g1514 ( 
.A(n_1403),
.Y(n_1514)
);

AO31x2_ASAP7_75t_L g1515 ( 
.A1(n_1410),
.A2(n_1363),
.A3(n_1365),
.B(n_1427),
.Y(n_1515)
);

INVx1_ASAP7_75t_L g1516 ( 
.A(n_1405),
.Y(n_1516)
);

INVx2_ASAP7_75t_L g1517 ( 
.A(n_1399),
.Y(n_1517)
);

NAND2x1p5_ASAP7_75t_L g1518 ( 
.A(n_1407),
.B(n_1403),
.Y(n_1518)
);

AND2x2_ASAP7_75t_L g1519 ( 
.A(n_1363),
.B(n_1365),
.Y(n_1519)
);

INVx4_ASAP7_75t_L g1520 ( 
.A(n_1403),
.Y(n_1520)
);

INVx1_ASAP7_75t_L g1521 ( 
.A(n_1395),
.Y(n_1521)
);

AND2x6_ASAP7_75t_L g1522 ( 
.A(n_1388),
.B(n_1412),
.Y(n_1522)
);

HB1xp67_ASAP7_75t_L g1523 ( 
.A(n_1344),
.Y(n_1523)
);

INVx1_ASAP7_75t_L g1524 ( 
.A(n_1395),
.Y(n_1524)
);

INVx1_ASAP7_75t_L g1525 ( 
.A(n_1424),
.Y(n_1525)
);

INVx1_ASAP7_75t_L g1526 ( 
.A(n_1427),
.Y(n_1526)
);

NOR2xp67_ASAP7_75t_SL g1527 ( 
.A(n_1411),
.B(n_1393),
.Y(n_1527)
);

INVx3_ASAP7_75t_L g1528 ( 
.A(n_1420),
.Y(n_1528)
);

INVx1_ASAP7_75t_L g1529 ( 
.A(n_1394),
.Y(n_1529)
);

INVx1_ASAP7_75t_L g1530 ( 
.A(n_1338),
.Y(n_1530)
);

INVx1_ASAP7_75t_L g1531 ( 
.A(n_1448),
.Y(n_1531)
);

BUFx2_ASAP7_75t_L g1532 ( 
.A(n_1366),
.Y(n_1532)
);

AND2x2_ASAP7_75t_L g1533 ( 
.A(n_1367),
.B(n_1452),
.Y(n_1533)
);

INVx1_ASAP7_75t_L g1534 ( 
.A(n_1390),
.Y(n_1534)
);

INVx3_ASAP7_75t_L g1535 ( 
.A(n_1346),
.Y(n_1535)
);

INVx1_ASAP7_75t_L g1536 ( 
.A(n_1390),
.Y(n_1536)
);

BUFx4f_ASAP7_75t_SL g1537 ( 
.A(n_1454),
.Y(n_1537)
);

INVx1_ASAP7_75t_L g1538 ( 
.A(n_1367),
.Y(n_1538)
);

INVxp67_ASAP7_75t_L g1539 ( 
.A(n_1381),
.Y(n_1539)
);

AND2x2_ASAP7_75t_L g1540 ( 
.A(n_1439),
.B(n_1440),
.Y(n_1540)
);

INVx2_ASAP7_75t_SL g1541 ( 
.A(n_1340),
.Y(n_1541)
);

AOI22xp33_ASAP7_75t_L g1542 ( 
.A1(n_1439),
.A2(n_1458),
.B1(n_1440),
.B2(n_1379),
.Y(n_1542)
);

AND2x2_ASAP7_75t_L g1543 ( 
.A(n_1458),
.B(n_1385),
.Y(n_1543)
);

AND2x2_ASAP7_75t_L g1544 ( 
.A(n_1385),
.B(n_1379),
.Y(n_1544)
);

AND2x2_ASAP7_75t_L g1545 ( 
.A(n_1396),
.B(n_1423),
.Y(n_1545)
);

INVx1_ASAP7_75t_L g1546 ( 
.A(n_1404),
.Y(n_1546)
);

HB1xp67_ASAP7_75t_L g1547 ( 
.A(n_1406),
.Y(n_1547)
);

BUFx2_ASAP7_75t_L g1548 ( 
.A(n_1392),
.Y(n_1548)
);

AND2x4_ASAP7_75t_L g1549 ( 
.A(n_1348),
.B(n_1382),
.Y(n_1549)
);

OA21x2_ASAP7_75t_L g1550 ( 
.A1(n_1408),
.A2(n_1462),
.B(n_1371),
.Y(n_1550)
);

BUFx2_ASAP7_75t_L g1551 ( 
.A(n_1342),
.Y(n_1551)
);

AND2x2_ASAP7_75t_L g1552 ( 
.A(n_1348),
.B(n_1449),
.Y(n_1552)
);

OR2x2_ASAP7_75t_L g1553 ( 
.A(n_1342),
.B(n_1463),
.Y(n_1553)
);

AND2x4_ASAP7_75t_L g1554 ( 
.A(n_1551),
.B(n_1463),
.Y(n_1554)
);

OR2x2_ASAP7_75t_L g1555 ( 
.A(n_1471),
.B(n_1442),
.Y(n_1555)
);

NAND2xp5_ASAP7_75t_L g1556 ( 
.A(n_1490),
.B(n_1442),
.Y(n_1556)
);

AND2x2_ASAP7_75t_L g1557 ( 
.A(n_1474),
.B(n_1401),
.Y(n_1557)
);

CKINVDCx6p67_ASAP7_75t_R g1558 ( 
.A(n_1496),
.Y(n_1558)
);

AOI22xp5_ASAP7_75t_L g1559 ( 
.A1(n_1502),
.A2(n_1482),
.B1(n_1540),
.B2(n_1480),
.Y(n_1559)
);

OAI22xp5_ASAP7_75t_L g1560 ( 
.A1(n_1512),
.A2(n_1461),
.B1(n_1453),
.B2(n_1356),
.Y(n_1560)
);

AOI211xp5_ASAP7_75t_SL g1561 ( 
.A1(n_1480),
.A2(n_1382),
.B(n_1449),
.C(n_1343),
.Y(n_1561)
);

NOR2xp33_ASAP7_75t_L g1562 ( 
.A(n_1497),
.B(n_1387),
.Y(n_1562)
);

NOR2xp33_ASAP7_75t_L g1563 ( 
.A(n_1493),
.B(n_1376),
.Y(n_1563)
);

INVxp67_ASAP7_75t_L g1564 ( 
.A(n_1523),
.Y(n_1564)
);

AND2x2_ASAP7_75t_L g1565 ( 
.A(n_1491),
.B(n_1340),
.Y(n_1565)
);

OR2x6_ASAP7_75t_L g1566 ( 
.A(n_1508),
.B(n_1467),
.Y(n_1566)
);

AND2x2_ASAP7_75t_L g1567 ( 
.A(n_1545),
.B(n_1386),
.Y(n_1567)
);

AND2x2_ASAP7_75t_L g1568 ( 
.A(n_1545),
.B(n_1386),
.Y(n_1568)
);

AO21x1_ASAP7_75t_L g1569 ( 
.A1(n_1540),
.A2(n_1383),
.B(n_1468),
.Y(n_1569)
);

NAND2xp5_ASAP7_75t_L g1570 ( 
.A(n_1476),
.B(n_1386),
.Y(n_1570)
);

AND2x2_ASAP7_75t_L g1571 ( 
.A(n_1506),
.B(n_1468),
.Y(n_1571)
);

OR2x2_ASAP7_75t_L g1572 ( 
.A(n_1479),
.B(n_1359),
.Y(n_1572)
);

OR2x2_ASAP7_75t_L g1573 ( 
.A(n_1510),
.B(n_1383),
.Y(n_1573)
);

NOR2xp33_ASAP7_75t_L g1574 ( 
.A(n_1539),
.B(n_1374),
.Y(n_1574)
);

AO21x1_ASAP7_75t_L g1575 ( 
.A1(n_1546),
.A2(n_1464),
.B(n_1445),
.Y(n_1575)
);

A2O1A1Ixp33_ASAP7_75t_L g1576 ( 
.A1(n_1470),
.A2(n_1352),
.B(n_1369),
.C(n_1360),
.Y(n_1576)
);

INVx2_ASAP7_75t_L g1577 ( 
.A(n_1485),
.Y(n_1577)
);

OAI22xp5_ASAP7_75t_L g1578 ( 
.A1(n_1542),
.A2(n_1445),
.B1(n_1354),
.B2(n_1357),
.Y(n_1578)
);

OAI21xp5_ASAP7_75t_L g1579 ( 
.A1(n_1533),
.A2(n_1465),
.B(n_1443),
.Y(n_1579)
);

AOI21xp5_ASAP7_75t_L g1580 ( 
.A1(n_1525),
.A2(n_1450),
.B(n_1354),
.Y(n_1580)
);

OAI21xp5_ASAP7_75t_L g1581 ( 
.A1(n_1533),
.A2(n_1362),
.B(n_1354),
.Y(n_1581)
);

CKINVDCx14_ASAP7_75t_R g1582 ( 
.A(n_1548),
.Y(n_1582)
);

OR2x2_ASAP7_75t_L g1583 ( 
.A(n_1510),
.B(n_1341),
.Y(n_1583)
);

NAND2xp5_ASAP7_75t_L g1584 ( 
.A(n_1530),
.B(n_1357),
.Y(n_1584)
);

OR2x2_ASAP7_75t_L g1585 ( 
.A(n_1534),
.B(n_1441),
.Y(n_1585)
);

OR2x2_ASAP7_75t_L g1586 ( 
.A(n_1534),
.B(n_1438),
.Y(n_1586)
);

AOI221xp5_ASAP7_75t_L g1587 ( 
.A1(n_1501),
.A2(n_1370),
.B1(n_1460),
.B2(n_1380),
.C(n_1357),
.Y(n_1587)
);

OR2x2_ASAP7_75t_L g1588 ( 
.A(n_1536),
.B(n_1380),
.Y(n_1588)
);

AOI211xp5_ASAP7_75t_L g1589 ( 
.A1(n_1501),
.A2(n_1398),
.B(n_1444),
.C(n_1447),
.Y(n_1589)
);

INVx1_ASAP7_75t_L g1590 ( 
.A(n_1498),
.Y(n_1590)
);

INVxp67_ASAP7_75t_L g1591 ( 
.A(n_1547),
.Y(n_1591)
);

OAI21xp5_ASAP7_75t_L g1592 ( 
.A1(n_1527),
.A2(n_1450),
.B(n_1505),
.Y(n_1592)
);

AOI21xp5_ASAP7_75t_SL g1593 ( 
.A1(n_1496),
.A2(n_1450),
.B(n_1550),
.Y(n_1593)
);

A2O1A1Ixp33_ASAP7_75t_L g1594 ( 
.A1(n_1527),
.A2(n_1505),
.B(n_1508),
.C(n_1519),
.Y(n_1594)
);

INVx3_ASAP7_75t_L g1595 ( 
.A(n_1550),
.Y(n_1595)
);

NOR2xp33_ASAP7_75t_L g1596 ( 
.A(n_1553),
.B(n_1532),
.Y(n_1596)
);

OR2x2_ASAP7_75t_L g1597 ( 
.A(n_1536),
.B(n_1487),
.Y(n_1597)
);

OAI22xp5_ASAP7_75t_L g1598 ( 
.A1(n_1546),
.A2(n_1496),
.B1(n_1519),
.B2(n_1530),
.Y(n_1598)
);

A2O1A1Ixp33_ASAP7_75t_L g1599 ( 
.A1(n_1543),
.A2(n_1531),
.B(n_1538),
.C(n_1544),
.Y(n_1599)
);

NAND2xp5_ASAP7_75t_L g1600 ( 
.A(n_1531),
.B(n_1516),
.Y(n_1600)
);

NOR2xp33_ASAP7_75t_L g1601 ( 
.A(n_1532),
.B(n_1548),
.Y(n_1601)
);

INVxp67_ASAP7_75t_L g1602 ( 
.A(n_1552),
.Y(n_1602)
);

AND2x4_ASAP7_75t_L g1603 ( 
.A(n_1469),
.B(n_1489),
.Y(n_1603)
);

NOR2xp33_ASAP7_75t_L g1604 ( 
.A(n_1537),
.B(n_1549),
.Y(n_1604)
);

AO21x2_ASAP7_75t_L g1605 ( 
.A1(n_1526),
.A2(n_1488),
.B(n_1504),
.Y(n_1605)
);

AOI22xp5_ASAP7_75t_L g1606 ( 
.A1(n_1543),
.A2(n_1538),
.B1(n_1475),
.B2(n_1544),
.Y(n_1606)
);

BUFx12f_ASAP7_75t_L g1607 ( 
.A(n_1511),
.Y(n_1607)
);

OAI22xp5_ASAP7_75t_L g1608 ( 
.A1(n_1518),
.A2(n_1535),
.B1(n_1520),
.B2(n_1514),
.Y(n_1608)
);

AO32x2_ASAP7_75t_L g1609 ( 
.A1(n_1513),
.A2(n_1520),
.A3(n_1507),
.B1(n_1484),
.B2(n_1541),
.Y(n_1609)
);

NAND2x1_ASAP7_75t_L g1610 ( 
.A(n_1528),
.B(n_1550),
.Y(n_1610)
);

NAND2xp5_ASAP7_75t_L g1611 ( 
.A(n_1516),
.B(n_1498),
.Y(n_1611)
);

NOR2x1_ASAP7_75t_SL g1612 ( 
.A(n_1487),
.B(n_1525),
.Y(n_1612)
);

AO32x2_ASAP7_75t_L g1613 ( 
.A1(n_1513),
.A2(n_1520),
.A3(n_1507),
.B1(n_1484),
.B2(n_1511),
.Y(n_1613)
);

NAND2xp5_ASAP7_75t_L g1614 ( 
.A(n_1499),
.B(n_1500),
.Y(n_1614)
);

AOI22xp5_ASAP7_75t_L g1615 ( 
.A1(n_1522),
.A2(n_1529),
.B1(n_1518),
.B2(n_1526),
.Y(n_1615)
);

AO32x2_ASAP7_75t_L g1616 ( 
.A1(n_1520),
.A2(n_1541),
.A3(n_1483),
.B1(n_1515),
.B2(n_1495),
.Y(n_1616)
);

INVx2_ASAP7_75t_L g1617 ( 
.A(n_1517),
.Y(n_1617)
);

AOI22xp5_ASAP7_75t_L g1618 ( 
.A1(n_1522),
.A2(n_1529),
.B1(n_1518),
.B2(n_1524),
.Y(n_1618)
);

NAND2x1_ASAP7_75t_L g1619 ( 
.A(n_1528),
.B(n_1550),
.Y(n_1619)
);

NAND2xp5_ASAP7_75t_L g1620 ( 
.A(n_1499),
.B(n_1500),
.Y(n_1620)
);

OR2x2_ASAP7_75t_L g1621 ( 
.A(n_1597),
.B(n_1495),
.Y(n_1621)
);

AND2x4_ASAP7_75t_L g1622 ( 
.A(n_1595),
.B(n_1472),
.Y(n_1622)
);

INVx3_ASAP7_75t_L g1623 ( 
.A(n_1595),
.Y(n_1623)
);

INVx2_ASAP7_75t_L g1624 ( 
.A(n_1617),
.Y(n_1624)
);

INVx3_ASAP7_75t_L g1625 ( 
.A(n_1610),
.Y(n_1625)
);

HB1xp67_ASAP7_75t_L g1626 ( 
.A(n_1619),
.Y(n_1626)
);

INVx1_ASAP7_75t_L g1627 ( 
.A(n_1590),
.Y(n_1627)
);

AOI22xp33_ASAP7_75t_L g1628 ( 
.A1(n_1559),
.A2(n_1522),
.B1(n_1492),
.B2(n_1503),
.Y(n_1628)
);

INVxp67_ASAP7_75t_SL g1629 ( 
.A(n_1600),
.Y(n_1629)
);

AND2x2_ASAP7_75t_L g1630 ( 
.A(n_1616),
.B(n_1488),
.Y(n_1630)
);

AND2x2_ASAP7_75t_L g1631 ( 
.A(n_1616),
.B(n_1605),
.Y(n_1631)
);

AND2x2_ASAP7_75t_L g1632 ( 
.A(n_1605),
.B(n_1618),
.Y(n_1632)
);

INVx1_ASAP7_75t_L g1633 ( 
.A(n_1614),
.Y(n_1633)
);

BUFx2_ASAP7_75t_L g1634 ( 
.A(n_1609),
.Y(n_1634)
);

INVx1_ASAP7_75t_L g1635 ( 
.A(n_1620),
.Y(n_1635)
);

INVx2_ASAP7_75t_L g1636 ( 
.A(n_1577),
.Y(n_1636)
);

INVx2_ASAP7_75t_L g1637 ( 
.A(n_1611),
.Y(n_1637)
);

BUFx3_ASAP7_75t_L g1638 ( 
.A(n_1558),
.Y(n_1638)
);

AND2x2_ASAP7_75t_L g1639 ( 
.A(n_1615),
.B(n_1503),
.Y(n_1639)
);

AND2x2_ASAP7_75t_L g1640 ( 
.A(n_1615),
.B(n_1503),
.Y(n_1640)
);

INVx1_ASAP7_75t_L g1641 ( 
.A(n_1609),
.Y(n_1641)
);

INVx1_ASAP7_75t_L g1642 ( 
.A(n_1613),
.Y(n_1642)
);

INVx1_ASAP7_75t_L g1643 ( 
.A(n_1613),
.Y(n_1643)
);

INVxp67_ASAP7_75t_L g1644 ( 
.A(n_1612),
.Y(n_1644)
);

BUFx2_ASAP7_75t_L g1645 ( 
.A(n_1603),
.Y(n_1645)
);

AOI21xp33_ASAP7_75t_L g1646 ( 
.A1(n_1559),
.A2(n_1524),
.B(n_1521),
.Y(n_1646)
);

INVx1_ASAP7_75t_SL g1647 ( 
.A(n_1555),
.Y(n_1647)
);

INVxp67_ASAP7_75t_L g1648 ( 
.A(n_1596),
.Y(n_1648)
);

NAND2xp5_ASAP7_75t_L g1649 ( 
.A(n_1606),
.B(n_1521),
.Y(n_1649)
);

INVxp67_ASAP7_75t_SL g1650 ( 
.A(n_1591),
.Y(n_1650)
);

INVxp67_ASAP7_75t_L g1651 ( 
.A(n_1556),
.Y(n_1651)
);

AND2x2_ASAP7_75t_L g1652 ( 
.A(n_1566),
.B(n_1492),
.Y(n_1652)
);

NOR2x1_ASAP7_75t_L g1653 ( 
.A(n_1593),
.B(n_1509),
.Y(n_1653)
);

BUFx2_ASAP7_75t_L g1654 ( 
.A(n_1566),
.Y(n_1654)
);

INVx2_ASAP7_75t_L g1655 ( 
.A(n_1588),
.Y(n_1655)
);

INVx1_ASAP7_75t_L g1656 ( 
.A(n_1602),
.Y(n_1656)
);

OR2x2_ASAP7_75t_L g1657 ( 
.A(n_1564),
.B(n_1483),
.Y(n_1657)
);

AOI22xp33_ASAP7_75t_L g1658 ( 
.A1(n_1649),
.A2(n_1569),
.B1(n_1560),
.B2(n_1585),
.Y(n_1658)
);

INVx1_ASAP7_75t_L g1659 ( 
.A(n_1627),
.Y(n_1659)
);

INVx2_ASAP7_75t_L g1660 ( 
.A(n_1623),
.Y(n_1660)
);

OR2x2_ASAP7_75t_L g1661 ( 
.A(n_1657),
.B(n_1494),
.Y(n_1661)
);

INVx2_ASAP7_75t_L g1662 ( 
.A(n_1623),
.Y(n_1662)
);

NAND2xp5_ASAP7_75t_L g1663 ( 
.A(n_1629),
.B(n_1481),
.Y(n_1663)
);

OAI33xp33_ASAP7_75t_L g1664 ( 
.A1(n_1649),
.A2(n_1598),
.A3(n_1584),
.B1(n_1586),
.B2(n_1572),
.B3(n_1573),
.Y(n_1664)
);

INVx1_ASAP7_75t_L g1665 ( 
.A(n_1624),
.Y(n_1665)
);

INVx2_ASAP7_75t_L g1666 ( 
.A(n_1623),
.Y(n_1666)
);

HB1xp67_ASAP7_75t_L g1667 ( 
.A(n_1641),
.Y(n_1667)
);

INVx2_ASAP7_75t_L g1668 ( 
.A(n_1623),
.Y(n_1668)
);

INVx3_ASAP7_75t_L g1669 ( 
.A(n_1622),
.Y(n_1669)
);

NAND2xp5_ASAP7_75t_L g1670 ( 
.A(n_1629),
.B(n_1637),
.Y(n_1670)
);

AOI211xp5_ASAP7_75t_L g1671 ( 
.A1(n_1646),
.A2(n_1576),
.B(n_1581),
.C(n_1587),
.Y(n_1671)
);

AND2x2_ASAP7_75t_L g1672 ( 
.A(n_1630),
.B(n_1567),
.Y(n_1672)
);

BUFx3_ASAP7_75t_L g1673 ( 
.A(n_1638),
.Y(n_1673)
);

OR2x2_ASAP7_75t_L g1674 ( 
.A(n_1657),
.B(n_1486),
.Y(n_1674)
);

INVx1_ASAP7_75t_L g1675 ( 
.A(n_1624),
.Y(n_1675)
);

OR2x2_ASAP7_75t_L g1676 ( 
.A(n_1657),
.B(n_1594),
.Y(n_1676)
);

OAI31xp33_ASAP7_75t_SL g1677 ( 
.A1(n_1646),
.A2(n_1581),
.A3(n_1592),
.B(n_1579),
.Y(n_1677)
);

INVx1_ASAP7_75t_SL g1678 ( 
.A(n_1645),
.Y(n_1678)
);

OAI221xp5_ASAP7_75t_L g1679 ( 
.A1(n_1628),
.A2(n_1589),
.B1(n_1599),
.B2(n_1583),
.C(n_1561),
.Y(n_1679)
);

OA21x2_ASAP7_75t_L g1680 ( 
.A1(n_1631),
.A2(n_1575),
.B(n_1478),
.Y(n_1680)
);

AND2x2_ASAP7_75t_L g1681 ( 
.A(n_1630),
.B(n_1568),
.Y(n_1681)
);

OR2x2_ASAP7_75t_L g1682 ( 
.A(n_1621),
.B(n_1473),
.Y(n_1682)
);

BUFx3_ASAP7_75t_L g1683 ( 
.A(n_1638),
.Y(n_1683)
);

NAND2xp33_ASAP7_75t_SL g1684 ( 
.A(n_1654),
.B(n_1557),
.Y(n_1684)
);

INVx2_ASAP7_75t_L g1685 ( 
.A(n_1636),
.Y(n_1685)
);

BUFx2_ASAP7_75t_L g1686 ( 
.A(n_1644),
.Y(n_1686)
);

OR2x2_ASAP7_75t_L g1687 ( 
.A(n_1621),
.B(n_1477),
.Y(n_1687)
);

OAI22xp5_ASAP7_75t_L g1688 ( 
.A1(n_1634),
.A2(n_1589),
.B1(n_1582),
.B2(n_1601),
.Y(n_1688)
);

OAI31xp33_ASAP7_75t_L g1689 ( 
.A1(n_1638),
.A2(n_1561),
.A3(n_1578),
.B(n_1608),
.Y(n_1689)
);

NAND2xp5_ASAP7_75t_L g1690 ( 
.A(n_1633),
.B(n_1635),
.Y(n_1690)
);

NAND2xp5_ASAP7_75t_L g1691 ( 
.A(n_1670),
.B(n_1635),
.Y(n_1691)
);

INVx1_ASAP7_75t_L g1692 ( 
.A(n_1685),
.Y(n_1692)
);

INVx2_ASAP7_75t_L g1693 ( 
.A(n_1680),
.Y(n_1693)
);

INVxp67_ASAP7_75t_L g1694 ( 
.A(n_1686),
.Y(n_1694)
);

NAND2xp5_ASAP7_75t_L g1695 ( 
.A(n_1670),
.B(n_1651),
.Y(n_1695)
);

NAND2xp5_ASAP7_75t_L g1696 ( 
.A(n_1690),
.B(n_1651),
.Y(n_1696)
);

AND2x2_ASAP7_75t_L g1697 ( 
.A(n_1669),
.B(n_1631),
.Y(n_1697)
);

AND2x2_ASAP7_75t_L g1698 ( 
.A(n_1669),
.B(n_1631),
.Y(n_1698)
);

AND2x2_ASAP7_75t_L g1699 ( 
.A(n_1660),
.B(n_1632),
.Y(n_1699)
);

AND2x2_ASAP7_75t_L g1700 ( 
.A(n_1660),
.B(n_1632),
.Y(n_1700)
);

INVx2_ASAP7_75t_L g1701 ( 
.A(n_1680),
.Y(n_1701)
);

AND2x2_ASAP7_75t_L g1702 ( 
.A(n_1660),
.B(n_1632),
.Y(n_1702)
);

INVx1_ASAP7_75t_L g1703 ( 
.A(n_1685),
.Y(n_1703)
);

AND2x2_ASAP7_75t_L g1704 ( 
.A(n_1662),
.B(n_1641),
.Y(n_1704)
);

INVx2_ASAP7_75t_L g1705 ( 
.A(n_1680),
.Y(n_1705)
);

INVx2_ASAP7_75t_L g1706 ( 
.A(n_1680),
.Y(n_1706)
);

INVx1_ASAP7_75t_L g1707 ( 
.A(n_1685),
.Y(n_1707)
);

NAND2xp5_ASAP7_75t_L g1708 ( 
.A(n_1690),
.B(n_1656),
.Y(n_1708)
);

NAND2xp5_ASAP7_75t_L g1709 ( 
.A(n_1659),
.B(n_1656),
.Y(n_1709)
);

NAND3xp33_ASAP7_75t_L g1710 ( 
.A(n_1677),
.B(n_1650),
.C(n_1653),
.Y(n_1710)
);

NAND2x1p5_ASAP7_75t_L g1711 ( 
.A(n_1680),
.B(n_1653),
.Y(n_1711)
);

AND2x2_ASAP7_75t_L g1712 ( 
.A(n_1667),
.B(n_1642),
.Y(n_1712)
);

INVx2_ASAP7_75t_L g1713 ( 
.A(n_1666),
.Y(n_1713)
);

INVx1_ASAP7_75t_L g1714 ( 
.A(n_1665),
.Y(n_1714)
);

INVx2_ASAP7_75t_L g1715 ( 
.A(n_1666),
.Y(n_1715)
);

INVx1_ASAP7_75t_L g1716 ( 
.A(n_1665),
.Y(n_1716)
);

AND2x2_ASAP7_75t_L g1717 ( 
.A(n_1667),
.B(n_1642),
.Y(n_1717)
);

INVx2_ASAP7_75t_SL g1718 ( 
.A(n_1666),
.Y(n_1718)
);

INVx1_ASAP7_75t_L g1719 ( 
.A(n_1675),
.Y(n_1719)
);

NAND2xp5_ASAP7_75t_SL g1720 ( 
.A(n_1677),
.B(n_1644),
.Y(n_1720)
);

NAND2xp5_ASAP7_75t_L g1721 ( 
.A(n_1659),
.B(n_1650),
.Y(n_1721)
);

INVx2_ASAP7_75t_L g1722 ( 
.A(n_1668),
.Y(n_1722)
);

INVx2_ASAP7_75t_L g1723 ( 
.A(n_1668),
.Y(n_1723)
);

NAND2xp67_ASAP7_75t_L g1724 ( 
.A(n_1663),
.B(n_1565),
.Y(n_1724)
);

AND2x2_ASAP7_75t_L g1725 ( 
.A(n_1672),
.B(n_1643),
.Y(n_1725)
);

AND2x2_ASAP7_75t_L g1726 ( 
.A(n_1725),
.B(n_1686),
.Y(n_1726)
);

INVx1_ASAP7_75t_SL g1727 ( 
.A(n_1720),
.Y(n_1727)
);

INVx2_ASAP7_75t_L g1728 ( 
.A(n_1718),
.Y(n_1728)
);

NOR2xp33_ASAP7_75t_L g1729 ( 
.A(n_1720),
.B(n_1664),
.Y(n_1729)
);

NAND2xp5_ASAP7_75t_L g1730 ( 
.A(n_1724),
.B(n_1676),
.Y(n_1730)
);

INVx1_ASAP7_75t_L g1731 ( 
.A(n_1721),
.Y(n_1731)
);

OR2x2_ASAP7_75t_L g1732 ( 
.A(n_1695),
.B(n_1676),
.Y(n_1732)
);

INVx1_ASAP7_75t_SL g1733 ( 
.A(n_1696),
.Y(n_1733)
);

INVx2_ASAP7_75t_L g1734 ( 
.A(n_1718),
.Y(n_1734)
);

NAND2xp5_ASAP7_75t_L g1735 ( 
.A(n_1724),
.B(n_1647),
.Y(n_1735)
);

INVx1_ASAP7_75t_L g1736 ( 
.A(n_1721),
.Y(n_1736)
);

INVx1_ASAP7_75t_L g1737 ( 
.A(n_1709),
.Y(n_1737)
);

OR2x2_ASAP7_75t_L g1738 ( 
.A(n_1695),
.B(n_1674),
.Y(n_1738)
);

AND2x2_ASAP7_75t_L g1739 ( 
.A(n_1725),
.B(n_1672),
.Y(n_1739)
);

INVx1_ASAP7_75t_L g1740 ( 
.A(n_1709),
.Y(n_1740)
);

AND2x4_ASAP7_75t_L g1741 ( 
.A(n_1694),
.B(n_1673),
.Y(n_1741)
);

INVx1_ASAP7_75t_L g1742 ( 
.A(n_1714),
.Y(n_1742)
);

AND2x2_ASAP7_75t_L g1743 ( 
.A(n_1725),
.B(n_1672),
.Y(n_1743)
);

INVx1_ASAP7_75t_L g1744 ( 
.A(n_1714),
.Y(n_1744)
);

AND2x2_ASAP7_75t_L g1745 ( 
.A(n_1699),
.B(n_1681),
.Y(n_1745)
);

OR2x2_ASAP7_75t_L g1746 ( 
.A(n_1696),
.B(n_1691),
.Y(n_1746)
);

NAND2xp5_ASAP7_75t_L g1747 ( 
.A(n_1724),
.B(n_1647),
.Y(n_1747)
);

AOI22xp5_ASAP7_75t_L g1748 ( 
.A1(n_1710),
.A2(n_1684),
.B1(n_1664),
.B2(n_1688),
.Y(n_1748)
);

INVx1_ASAP7_75t_L g1749 ( 
.A(n_1714),
.Y(n_1749)
);

NAND2xp5_ASAP7_75t_L g1750 ( 
.A(n_1710),
.B(n_1648),
.Y(n_1750)
);

OR2x2_ASAP7_75t_L g1751 ( 
.A(n_1691),
.B(n_1674),
.Y(n_1751)
);

AND2x4_ASAP7_75t_L g1752 ( 
.A(n_1694),
.B(n_1673),
.Y(n_1752)
);

OR2x2_ASAP7_75t_L g1753 ( 
.A(n_1708),
.B(n_1655),
.Y(n_1753)
);

INVx1_ASAP7_75t_L g1754 ( 
.A(n_1716),
.Y(n_1754)
);

INVx1_ASAP7_75t_L g1755 ( 
.A(n_1716),
.Y(n_1755)
);

INVx2_ASAP7_75t_L g1756 ( 
.A(n_1718),
.Y(n_1756)
);

HB1xp67_ASAP7_75t_L g1757 ( 
.A(n_1708),
.Y(n_1757)
);

NAND2xp5_ASAP7_75t_L g1758 ( 
.A(n_1699),
.B(n_1648),
.Y(n_1758)
);

INVx1_ASAP7_75t_L g1759 ( 
.A(n_1716),
.Y(n_1759)
);

INVxp67_ASAP7_75t_L g1760 ( 
.A(n_1712),
.Y(n_1760)
);

INVx1_ASAP7_75t_L g1761 ( 
.A(n_1719),
.Y(n_1761)
);

INVx2_ASAP7_75t_SL g1762 ( 
.A(n_1718),
.Y(n_1762)
);

NAND2xp5_ASAP7_75t_SL g1763 ( 
.A(n_1711),
.B(n_1688),
.Y(n_1763)
);

INVx1_ASAP7_75t_L g1764 ( 
.A(n_1719),
.Y(n_1764)
);

NOR3xp33_ASAP7_75t_L g1765 ( 
.A(n_1693),
.B(n_1671),
.C(n_1679),
.Y(n_1765)
);

INVx1_ASAP7_75t_L g1766 ( 
.A(n_1719),
.Y(n_1766)
);

INVx2_ASAP7_75t_SL g1767 ( 
.A(n_1711),
.Y(n_1767)
);

INVx1_ASAP7_75t_L g1768 ( 
.A(n_1704),
.Y(n_1768)
);

INVx1_ASAP7_75t_L g1769 ( 
.A(n_1742),
.Y(n_1769)
);

OR2x2_ASAP7_75t_L g1770 ( 
.A(n_1732),
.B(n_1661),
.Y(n_1770)
);

NAND2xp5_ASAP7_75t_L g1771 ( 
.A(n_1727),
.B(n_1681),
.Y(n_1771)
);

AND2x2_ASAP7_75t_L g1772 ( 
.A(n_1726),
.B(n_1699),
.Y(n_1772)
);

INVx1_ASAP7_75t_L g1773 ( 
.A(n_1744),
.Y(n_1773)
);

NOR3xp33_ASAP7_75t_SL g1774 ( 
.A(n_1729),
.B(n_1679),
.C(n_1689),
.Y(n_1774)
);

NAND2xp5_ASAP7_75t_L g1775 ( 
.A(n_1729),
.B(n_1681),
.Y(n_1775)
);

AND2x2_ASAP7_75t_L g1776 ( 
.A(n_1726),
.B(n_1699),
.Y(n_1776)
);

OR2x2_ASAP7_75t_L g1777 ( 
.A(n_1732),
.B(n_1661),
.Y(n_1777)
);

INVx1_ASAP7_75t_L g1778 ( 
.A(n_1749),
.Y(n_1778)
);

AND2x2_ASAP7_75t_L g1779 ( 
.A(n_1739),
.B(n_1700),
.Y(n_1779)
);

NOR2xp33_ASAP7_75t_SL g1780 ( 
.A(n_1765),
.B(n_1689),
.Y(n_1780)
);

NAND2xp5_ASAP7_75t_L g1781 ( 
.A(n_1750),
.B(n_1733),
.Y(n_1781)
);

NAND2x1p5_ASAP7_75t_L g1782 ( 
.A(n_1763),
.B(n_1673),
.Y(n_1782)
);

INVx1_ASAP7_75t_L g1783 ( 
.A(n_1754),
.Y(n_1783)
);

AND2x2_ASAP7_75t_L g1784 ( 
.A(n_1739),
.B(n_1700),
.Y(n_1784)
);

OR2x2_ASAP7_75t_L g1785 ( 
.A(n_1746),
.B(n_1682),
.Y(n_1785)
);

HB1xp67_ASAP7_75t_L g1786 ( 
.A(n_1741),
.Y(n_1786)
);

OAI21xp5_ASAP7_75t_L g1787 ( 
.A1(n_1748),
.A2(n_1711),
.B(n_1671),
.Y(n_1787)
);

OR2x2_ASAP7_75t_L g1788 ( 
.A(n_1746),
.B(n_1682),
.Y(n_1788)
);

OR2x2_ASAP7_75t_L g1789 ( 
.A(n_1738),
.B(n_1687),
.Y(n_1789)
);

AND2x4_ASAP7_75t_L g1790 ( 
.A(n_1741),
.B(n_1752),
.Y(n_1790)
);

INVx1_ASAP7_75t_L g1791 ( 
.A(n_1755),
.Y(n_1791)
);

OR2x2_ASAP7_75t_L g1792 ( 
.A(n_1738),
.B(n_1687),
.Y(n_1792)
);

OR2x2_ASAP7_75t_L g1793 ( 
.A(n_1758),
.B(n_1663),
.Y(n_1793)
);

NAND2xp5_ASAP7_75t_L g1794 ( 
.A(n_1730),
.B(n_1683),
.Y(n_1794)
);

NAND2xp5_ASAP7_75t_L g1795 ( 
.A(n_1741),
.B(n_1683),
.Y(n_1795)
);

INVx1_ASAP7_75t_L g1796 ( 
.A(n_1759),
.Y(n_1796)
);

AND2x2_ASAP7_75t_L g1797 ( 
.A(n_1743),
.B(n_1700),
.Y(n_1797)
);

INVx2_ASAP7_75t_L g1798 ( 
.A(n_1762),
.Y(n_1798)
);

INVx2_ASAP7_75t_L g1799 ( 
.A(n_1762),
.Y(n_1799)
);

INVx1_ASAP7_75t_L g1800 ( 
.A(n_1761),
.Y(n_1800)
);

AND2x2_ASAP7_75t_L g1801 ( 
.A(n_1743),
.B(n_1700),
.Y(n_1801)
);

AND2x2_ASAP7_75t_L g1802 ( 
.A(n_1752),
.B(n_1702),
.Y(n_1802)
);

INVx1_ASAP7_75t_L g1803 ( 
.A(n_1764),
.Y(n_1803)
);

AND2x2_ASAP7_75t_L g1804 ( 
.A(n_1752),
.B(n_1702),
.Y(n_1804)
);

INVx1_ASAP7_75t_L g1805 ( 
.A(n_1769),
.Y(n_1805)
);

OAI21xp5_ASAP7_75t_L g1806 ( 
.A1(n_1787),
.A2(n_1763),
.B(n_1711),
.Y(n_1806)
);

AND2x2_ASAP7_75t_L g1807 ( 
.A(n_1790),
.B(n_1745),
.Y(n_1807)
);

OAI22xp5_ASAP7_75t_L g1808 ( 
.A1(n_1782),
.A2(n_1658),
.B1(n_1711),
.B2(n_1735),
.Y(n_1808)
);

INVx1_ASAP7_75t_L g1809 ( 
.A(n_1769),
.Y(n_1809)
);

AOI31xp33_ASAP7_75t_L g1810 ( 
.A1(n_1782),
.A2(n_1562),
.A3(n_1747),
.B(n_1563),
.Y(n_1810)
);

O2A1O1Ixp33_ASAP7_75t_L g1811 ( 
.A1(n_1780),
.A2(n_1757),
.B(n_1767),
.C(n_1731),
.Y(n_1811)
);

OAI22xp5_ASAP7_75t_L g1812 ( 
.A1(n_1782),
.A2(n_1683),
.B1(n_1760),
.B2(n_1654),
.Y(n_1812)
);

INVx1_ASAP7_75t_L g1813 ( 
.A(n_1773),
.Y(n_1813)
);

AOI22xp5_ASAP7_75t_L g1814 ( 
.A1(n_1774),
.A2(n_1736),
.B1(n_1740),
.B2(n_1737),
.Y(n_1814)
);

INVx1_ASAP7_75t_L g1815 ( 
.A(n_1773),
.Y(n_1815)
);

OR2x2_ASAP7_75t_L g1816 ( 
.A(n_1775),
.B(n_1751),
.Y(n_1816)
);

OAI22xp5_ASAP7_75t_L g1817 ( 
.A1(n_1781),
.A2(n_1745),
.B1(n_1678),
.B2(n_1693),
.Y(n_1817)
);

AOI322xp5_ASAP7_75t_L g1818 ( 
.A1(n_1771),
.A2(n_1797),
.A3(n_1784),
.B1(n_1779),
.B2(n_1801),
.C1(n_1776),
.C2(n_1772),
.Y(n_1818)
);

NAND2xp5_ASAP7_75t_L g1819 ( 
.A(n_1786),
.B(n_1751),
.Y(n_1819)
);

AOI21xp5_ASAP7_75t_L g1820 ( 
.A1(n_1794),
.A2(n_1701),
.B(n_1693),
.Y(n_1820)
);

INVx2_ASAP7_75t_L g1821 ( 
.A(n_1790),
.Y(n_1821)
);

INVx1_ASAP7_75t_L g1822 ( 
.A(n_1783),
.Y(n_1822)
);

AOI222xp33_ASAP7_75t_L g1823 ( 
.A1(n_1790),
.A2(n_1705),
.B1(n_1693),
.B2(n_1701),
.C1(n_1706),
.C2(n_1712),
.Y(n_1823)
);

OAI22xp5_ASAP7_75t_SL g1824 ( 
.A1(n_1795),
.A2(n_1574),
.B1(n_1604),
.B2(n_1767),
.Y(n_1824)
);

INVxp67_ASAP7_75t_SL g1825 ( 
.A(n_1798),
.Y(n_1825)
);

AOI22xp5_ASAP7_75t_L g1826 ( 
.A1(n_1802),
.A2(n_1652),
.B1(n_1639),
.B2(n_1640),
.Y(n_1826)
);

INVx1_ASAP7_75t_SL g1827 ( 
.A(n_1802),
.Y(n_1827)
);

AND2x2_ASAP7_75t_L g1828 ( 
.A(n_1804),
.B(n_1768),
.Y(n_1828)
);

OAI22xp33_ASAP7_75t_SL g1829 ( 
.A1(n_1770),
.A2(n_1706),
.B1(n_1705),
.B2(n_1701),
.Y(n_1829)
);

NAND2xp5_ASAP7_75t_L g1830 ( 
.A(n_1804),
.B(n_1753),
.Y(n_1830)
);

INVx1_ASAP7_75t_SL g1831 ( 
.A(n_1827),
.Y(n_1831)
);

INVx1_ASAP7_75t_L g1832 ( 
.A(n_1825),
.Y(n_1832)
);

INVx3_ASAP7_75t_L g1833 ( 
.A(n_1821),
.Y(n_1833)
);

INVx1_ASAP7_75t_SL g1834 ( 
.A(n_1807),
.Y(n_1834)
);

OA22x2_ASAP7_75t_L g1835 ( 
.A1(n_1806),
.A2(n_1799),
.B1(n_1798),
.B2(n_1701),
.Y(n_1835)
);

OR2x2_ASAP7_75t_L g1836 ( 
.A(n_1819),
.B(n_1770),
.Y(n_1836)
);

AOI211xp5_ASAP7_75t_L g1837 ( 
.A1(n_1808),
.A2(n_1778),
.B(n_1796),
.C(n_1800),
.Y(n_1837)
);

AND2x2_ASAP7_75t_L g1838 ( 
.A(n_1807),
.B(n_1772),
.Y(n_1838)
);

INVx1_ASAP7_75t_L g1839 ( 
.A(n_1825),
.Y(n_1839)
);

OAI21xp5_ASAP7_75t_L g1840 ( 
.A1(n_1811),
.A2(n_1799),
.B(n_1793),
.Y(n_1840)
);

HB1xp67_ASAP7_75t_L g1841 ( 
.A(n_1821),
.Y(n_1841)
);

INVx1_ASAP7_75t_L g1842 ( 
.A(n_1805),
.Y(n_1842)
);

INVx1_ASAP7_75t_L g1843 ( 
.A(n_1809),
.Y(n_1843)
);

INVx1_ASAP7_75t_L g1844 ( 
.A(n_1813),
.Y(n_1844)
);

INVx1_ASAP7_75t_L g1845 ( 
.A(n_1815),
.Y(n_1845)
);

INVx1_ASAP7_75t_L g1846 ( 
.A(n_1822),
.Y(n_1846)
);

OAI22xp33_ASAP7_75t_L g1847 ( 
.A1(n_1810),
.A2(n_1814),
.B1(n_1812),
.B2(n_1826),
.Y(n_1847)
);

OAI22xp33_ASAP7_75t_L g1848 ( 
.A1(n_1817),
.A2(n_1706),
.B1(n_1705),
.B2(n_1777),
.Y(n_1848)
);

AOI22xp5_ASAP7_75t_L g1849 ( 
.A1(n_1824),
.A2(n_1776),
.B1(n_1803),
.B2(n_1800),
.Y(n_1849)
);

OAI221xp5_ASAP7_75t_SL g1850 ( 
.A1(n_1818),
.A2(n_1706),
.B1(n_1705),
.B2(n_1777),
.C(n_1793),
.Y(n_1850)
);

A2O1A1Ixp33_ASAP7_75t_L g1851 ( 
.A1(n_1849),
.A2(n_1820),
.B(n_1816),
.C(n_1783),
.Y(n_1851)
);

INVx1_ASAP7_75t_L g1852 ( 
.A(n_1841),
.Y(n_1852)
);

AOI21xp5_ASAP7_75t_L g1853 ( 
.A1(n_1847),
.A2(n_1829),
.B(n_1823),
.Y(n_1853)
);

XNOR2xp5_ASAP7_75t_L g1854 ( 
.A(n_1834),
.B(n_1830),
.Y(n_1854)
);

NAND2xp5_ASAP7_75t_L g1855 ( 
.A(n_1831),
.B(n_1828),
.Y(n_1855)
);

INVx1_ASAP7_75t_L g1856 ( 
.A(n_1841),
.Y(n_1856)
);

INVx1_ASAP7_75t_L g1857 ( 
.A(n_1832),
.Y(n_1857)
);

NAND2xp5_ASAP7_75t_L g1858 ( 
.A(n_1833),
.B(n_1828),
.Y(n_1858)
);

INVx1_ASAP7_75t_L g1859 ( 
.A(n_1839),
.Y(n_1859)
);

INVx2_ASAP7_75t_L g1860 ( 
.A(n_1833),
.Y(n_1860)
);

NOR2xp33_ASAP7_75t_L g1861 ( 
.A(n_1836),
.B(n_1785),
.Y(n_1861)
);

INVx1_ASAP7_75t_L g1862 ( 
.A(n_1842),
.Y(n_1862)
);

OAI211xp5_ASAP7_75t_L g1863 ( 
.A1(n_1853),
.A2(n_1837),
.B(n_1850),
.C(n_1840),
.Y(n_1863)
);

INVxp67_ASAP7_75t_L g1864 ( 
.A(n_1852),
.Y(n_1864)
);

INVx1_ASAP7_75t_L g1865 ( 
.A(n_1856),
.Y(n_1865)
);

NOR2x1_ASAP7_75t_L g1866 ( 
.A(n_1860),
.B(n_1843),
.Y(n_1866)
);

AND2x2_ASAP7_75t_L g1867 ( 
.A(n_1861),
.B(n_1838),
.Y(n_1867)
);

NAND2xp5_ASAP7_75t_L g1868 ( 
.A(n_1854),
.B(n_1844),
.Y(n_1868)
);

INVx1_ASAP7_75t_L g1869 ( 
.A(n_1855),
.Y(n_1869)
);

NOR2xp33_ASAP7_75t_L g1870 ( 
.A(n_1861),
.B(n_1845),
.Y(n_1870)
);

AOI21xp5_ASAP7_75t_L g1871 ( 
.A1(n_1851),
.A2(n_1850),
.B(n_1835),
.Y(n_1871)
);

NAND2xp5_ASAP7_75t_L g1872 ( 
.A(n_1858),
.B(n_1846),
.Y(n_1872)
);

OAI211xp5_ASAP7_75t_L g1873 ( 
.A1(n_1851),
.A2(n_1835),
.B(n_1791),
.C(n_1803),
.Y(n_1873)
);

INVx1_ASAP7_75t_SL g1874 ( 
.A(n_1857),
.Y(n_1874)
);

AOI31xp33_ASAP7_75t_L g1875 ( 
.A1(n_1868),
.A2(n_1859),
.A3(n_1862),
.B(n_1848),
.Y(n_1875)
);

AND2x4_ASAP7_75t_L g1876 ( 
.A(n_1867),
.B(n_1779),
.Y(n_1876)
);

AOI222xp33_ASAP7_75t_L g1877 ( 
.A1(n_1863),
.A2(n_1848),
.B1(n_1791),
.B2(n_1801),
.C1(n_1797),
.C2(n_1784),
.Y(n_1877)
);

AOI211xp5_ASAP7_75t_L g1878 ( 
.A1(n_1871),
.A2(n_1788),
.B(n_1785),
.C(n_1792),
.Y(n_1878)
);

AOI221xp5_ASAP7_75t_L g1879 ( 
.A1(n_1870),
.A2(n_1766),
.B1(n_1788),
.B2(n_1756),
.C(n_1734),
.Y(n_1879)
);

OAI211xp5_ASAP7_75t_L g1880 ( 
.A1(n_1873),
.A2(n_1864),
.B(n_1866),
.C(n_1874),
.Y(n_1880)
);

OAI22xp33_ASAP7_75t_L g1881 ( 
.A1(n_1869),
.A2(n_1792),
.B1(n_1789),
.B2(n_1756),
.Y(n_1881)
);

AOI221x1_ASAP7_75t_L g1882 ( 
.A1(n_1876),
.A2(n_1865),
.B1(n_1872),
.B2(n_1864),
.C(n_1734),
.Y(n_1882)
);

OAI211xp5_ASAP7_75t_SL g1883 ( 
.A1(n_1880),
.A2(n_1789),
.B(n_1728),
.C(n_1678),
.Y(n_1883)
);

INVx1_ASAP7_75t_SL g1884 ( 
.A(n_1875),
.Y(n_1884)
);

OAI211xp5_ASAP7_75t_L g1885 ( 
.A1(n_1878),
.A2(n_1728),
.B(n_1626),
.C(n_1580),
.Y(n_1885)
);

OAI211xp5_ASAP7_75t_L g1886 ( 
.A1(n_1877),
.A2(n_1626),
.B(n_1712),
.C(n_1717),
.Y(n_1886)
);

O2A1O1Ixp33_ASAP7_75t_L g1887 ( 
.A1(n_1881),
.A2(n_1717),
.B(n_1702),
.C(n_1698),
.Y(n_1887)
);

NOR3xp33_ASAP7_75t_L g1888 ( 
.A(n_1879),
.B(n_1625),
.C(n_1570),
.Y(n_1888)
);

INVx2_ASAP7_75t_SL g1889 ( 
.A(n_1884),
.Y(n_1889)
);

XOR2xp5_ASAP7_75t_L g1890 ( 
.A(n_1883),
.B(n_1554),
.Y(n_1890)
);

INVx1_ASAP7_75t_SL g1891 ( 
.A(n_1882),
.Y(n_1891)
);

NAND3xp33_ASAP7_75t_L g1892 ( 
.A(n_1886),
.B(n_1717),
.C(n_1692),
.Y(n_1892)
);

INVx1_ASAP7_75t_L g1893 ( 
.A(n_1885),
.Y(n_1893)
);

NOR3xp33_ASAP7_75t_L g1894 ( 
.A(n_1889),
.B(n_1888),
.C(n_1887),
.Y(n_1894)
);

AND2x2_ASAP7_75t_L g1895 ( 
.A(n_1893),
.B(n_1697),
.Y(n_1895)
);

OAI211xp5_ASAP7_75t_L g1896 ( 
.A1(n_1891),
.A2(n_1890),
.B(n_1892),
.C(n_1702),
.Y(n_1896)
);

INVxp33_ASAP7_75t_L g1897 ( 
.A(n_1894),
.Y(n_1897)
);

OAI22xp5_ASAP7_75t_L g1898 ( 
.A1(n_1897),
.A2(n_1896),
.B1(n_1895),
.B2(n_1723),
.Y(n_1898)
);

INVx1_ASAP7_75t_L g1899 ( 
.A(n_1898),
.Y(n_1899)
);

AO22x1_ASAP7_75t_L g1900 ( 
.A1(n_1898),
.A2(n_1698),
.B1(n_1697),
.B2(n_1722),
.Y(n_1900)
);

XNOR2xp5_ASAP7_75t_L g1901 ( 
.A(n_1899),
.B(n_1571),
.Y(n_1901)
);

OAI22xp5_ASAP7_75t_SL g1902 ( 
.A1(n_1900),
.A2(n_1607),
.B1(n_1722),
.B2(n_1715),
.Y(n_1902)
);

OAI21xp33_ASAP7_75t_SL g1903 ( 
.A1(n_1901),
.A2(n_1713),
.B(n_1722),
.Y(n_1903)
);

AOI22x1_ASAP7_75t_L g1904 ( 
.A1(n_1902),
.A2(n_1723),
.B1(n_1713),
.B2(n_1722),
.Y(n_1904)
);

AOI21xp5_ASAP7_75t_L g1905 ( 
.A1(n_1904),
.A2(n_1723),
.B(n_1713),
.Y(n_1905)
);

AND2x2_ASAP7_75t_L g1906 ( 
.A(n_1905),
.B(n_1903),
.Y(n_1906)
);

OAI22xp5_ASAP7_75t_L g1907 ( 
.A1(n_1906),
.A2(n_1723),
.B1(n_1715),
.B2(n_1713),
.Y(n_1907)
);

AOI221xp5_ASAP7_75t_L g1908 ( 
.A1(n_1907),
.A2(n_1692),
.B1(n_1703),
.B2(n_1707),
.C(n_1715),
.Y(n_1908)
);

AOI211xp5_ASAP7_75t_L g1909 ( 
.A1(n_1908),
.A2(n_1707),
.B(n_1692),
.C(n_1703),
.Y(n_1909)
);


endmodule