module real_jpeg_760_n_6 (n_5, n_4, n_0, n_1, n_2, n_3, n_6);

input n_5;
input n_4;
input n_0;
input n_1;
input n_2;
input n_3;

output n_6;

wire n_17;
wire n_8;
wire n_43;
wire n_37;
wire n_21;
wire n_35;
wire n_33;
wire n_50;
wire n_38;
wire n_29;
wire n_49;
wire n_10;
wire n_31;
wire n_9;
wire n_12;
wire n_24;
wire n_34;
wire n_28;
wire n_44;
wire n_46;
wire n_23;
wire n_11;
wire n_14;
wire n_47;
wire n_45;
wire n_25;
wire n_42;
wire n_7;
wire n_22;
wire n_18;
wire n_40;
wire n_36;
wire n_39;
wire n_41;
wire n_26;
wire n_27;
wire n_20;
wire n_48;
wire n_19;
wire n_32;
wire n_30;
wire n_16;
wire n_15;
wire n_13;

NAND2xp5_ASAP7_75t_L g8 ( 
.A(n_0),
.B(n_9),
.Y(n_8)
);

INVx1_ASAP7_75t_SL g22 ( 
.A(n_0),
.Y(n_22)
);

NOR2xp33_ASAP7_75t_L g33 ( 
.A(n_0),
.B(n_10),
.Y(n_33)
);

NAND2xp5_ASAP7_75t_L g45 ( 
.A(n_0),
.B(n_40),
.Y(n_45)
);

NAND2xp5_ASAP7_75t_L g49 ( 
.A(n_0),
.B(n_48),
.Y(n_49)
);

INVx1_ASAP7_75t_SL g11 ( 
.A(n_1),
.Y(n_11)
);

OR2x4_ASAP7_75t_L g24 ( 
.A(n_1),
.B(n_25),
.Y(n_24)
);

AND2x2_ASAP7_75t_SL g40 ( 
.A(n_1),
.B(n_41),
.Y(n_40)
);

OA22x2_ASAP7_75t_L g13 ( 
.A1(n_2),
.A2(n_14),
.B1(n_15),
.B2(n_16),
.Y(n_13)
);

CKINVDCx20_ASAP7_75t_R g14 ( 
.A(n_2),
.Y(n_14)
);

AO21x1_ASAP7_75t_L g27 ( 
.A1(n_2),
.A2(n_28),
.B(n_30),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_3),
.Y(n_19)
);

NOR2xp33_ASAP7_75t_L g29 ( 
.A(n_3),
.B(n_4),
.Y(n_29)
);

NAND2xp5_ASAP7_75t_L g31 ( 
.A(n_3),
.B(n_4),
.Y(n_31)
);

NOR2xp33_ASAP7_75t_L g18 ( 
.A(n_4),
.B(n_19),
.Y(n_18)
);

NAND2x1_ASAP7_75t_SL g20 ( 
.A(n_4),
.B(n_19),
.Y(n_20)
);

OR2x2_ASAP7_75t_L g10 ( 
.A(n_5),
.B(n_11),
.Y(n_10)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_5),
.Y(n_25)
);

NOR4xp25_ASAP7_75t_L g6 ( 
.A(n_7),
.B(n_26),
.C(n_37),
.D(n_46),
.Y(n_6)
);

OAI22xp5_ASAP7_75t_L g7 ( 
.A1(n_8),
.A2(n_12),
.B1(n_13),
.B2(n_21),
.Y(n_7)
);

INVx1_ASAP7_75t_SL g9 ( 
.A(n_10),
.Y(n_9)
);

AND2x2_ASAP7_75t_SL g48 ( 
.A(n_11),
.B(n_25),
.Y(n_48)
);

CKINVDCx20_ASAP7_75t_R g12 ( 
.A(n_13),
.Y(n_12)
);

NOR2xp33_ASAP7_75t_SL g38 ( 
.A(n_14),
.B(n_22),
.Y(n_38)
);

OA21x2_ASAP7_75t_L g43 ( 
.A1(n_14),
.A2(n_18),
.B(n_20),
.Y(n_43)
);

O2A1O1Ixp33_ASAP7_75t_SL g46 ( 
.A1(n_14),
.A2(n_47),
.B(n_49),
.C(n_50),
.Y(n_46)
);

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_16),
.Y(n_15)
);

AND2x2_ASAP7_75t_L g16 ( 
.A(n_17),
.B(n_20),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_18),
.Y(n_17)
);

NAND2xp5_ASAP7_75t_L g21 ( 
.A(n_22),
.B(n_23),
.Y(n_21)
);

NOR2xp33_ASAP7_75t_L g36 ( 
.A(n_22),
.B(n_24),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_SL g50 ( 
.A(n_22),
.B(n_43),
.Y(n_50)
);

INVx1_ASAP7_75t_SL g23 ( 
.A(n_24),
.Y(n_23)
);

CKINVDCx16_ASAP7_75t_R g41 ( 
.A(n_25),
.Y(n_41)
);

OAI22xp5_ASAP7_75t_L g26 ( 
.A1(n_27),
.A2(n_32),
.B1(n_34),
.B2(n_35),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_27),
.Y(n_34)
);

INVxp67_ASAP7_75t_L g28 ( 
.A(n_29),
.Y(n_28)
);

CKINVDCx16_ASAP7_75t_R g30 ( 
.A(n_31),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_33),
.Y(n_32)
);

CKINVDCx16_ASAP7_75t_R g35 ( 
.A(n_36),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g37 ( 
.A(n_38),
.B(n_39),
.Y(n_37)
);

AOI21xp5_ASAP7_75t_L g39 ( 
.A1(n_40),
.A2(n_42),
.B(n_44),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_43),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_45),
.Y(n_44)
);

INVx1_ASAP7_75t_SL g47 ( 
.A(n_48),
.Y(n_47)
);


endmodule