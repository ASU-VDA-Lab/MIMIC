module fake_jpeg_2491_n_290 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_290);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_290;

wire n_159;
wire n_117;
wire n_253;
wire n_286;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_182;
wire n_19;
wire n_152;
wire n_59;
wire n_84;
wire n_98;
wire n_252;
wire n_251;
wire n_273;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_279;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_127;
wire n_76;
wire n_154;
wire n_278;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_281;
wire n_31;
wire n_155;
wire n_207;
wire n_277;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_223;
wire n_187;
wire n_57;
wire n_21;
wire n_175;
wire n_234;
wire n_284;
wire n_272;
wire n_288;
wire n_280;
wire n_171;
wire n_263;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_289;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_267;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_274;
wire n_186;
wire n_44;
wire n_24;
wire n_276;
wire n_143;
wire n_202;
wire n_25;
wire n_17;
wire n_269;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_287;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_266;
wire n_34;
wire n_283;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_285;
wire n_215;
wire n_262;
wire n_131;
wire n_56;
wire n_240;
wire n_212;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_271;
wire n_216;
wire n_217;
wire n_264;
wire n_184;
wire n_53;
wire n_268;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_48;
wire n_35;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_270;
wire n_176;
wire n_199;
wire n_112;
wire n_260;
wire n_265;
wire n_222;
wire n_95;
wire n_275;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_258;
wire n_282;
wire n_96;

INVx1_ASAP7_75t_L g17 ( 
.A(n_6),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_11),
.Y(n_18)
);

BUFx12f_ASAP7_75t_L g19 ( 
.A(n_16),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_10),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_11),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_4),
.Y(n_22)
);

INVx2_ASAP7_75t_L g23 ( 
.A(n_15),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_0),
.Y(n_24)
);

BUFx16f_ASAP7_75t_L g25 ( 
.A(n_1),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_1),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_3),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_11),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_0),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_6),
.Y(n_30)
);

CKINVDCx16_ASAP7_75t_R g31 ( 
.A(n_16),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_9),
.Y(n_32)
);

BUFx3_ASAP7_75t_L g33 ( 
.A(n_8),
.Y(n_33)
);

INVx5_ASAP7_75t_L g34 ( 
.A(n_12),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_1),
.Y(n_35)
);

BUFx3_ASAP7_75t_L g36 ( 
.A(n_8),
.Y(n_36)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_14),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_8),
.Y(n_38)
);

INVx4_ASAP7_75t_L g39 ( 
.A(n_2),
.Y(n_39)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_16),
.Y(n_40)
);

INVx2_ASAP7_75t_L g41 ( 
.A(n_23),
.Y(n_41)
);

INVx2_ASAP7_75t_L g99 ( 
.A(n_41),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_SL g42 ( 
.A(n_18),
.B(n_7),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_42),
.B(n_31),
.Y(n_72)
);

INVx2_ASAP7_75t_SL g43 ( 
.A(n_25),
.Y(n_43)
);

INVx2_ASAP7_75t_SL g66 ( 
.A(n_43),
.Y(n_66)
);

CKINVDCx6p67_ASAP7_75t_R g44 ( 
.A(n_25),
.Y(n_44)
);

CKINVDCx9p33_ASAP7_75t_R g65 ( 
.A(n_44),
.Y(n_65)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_32),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_45),
.Y(n_68)
);

INVx2_ASAP7_75t_L g46 ( 
.A(n_23),
.Y(n_46)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_46),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_L g47 ( 
.A(n_39),
.B(n_0),
.Y(n_47)
);

NAND2xp5_ASAP7_75t_L g82 ( 
.A(n_47),
.B(n_49),
.Y(n_82)
);

INVx11_ASAP7_75t_L g48 ( 
.A(n_25),
.Y(n_48)
);

INVx4_ASAP7_75t_L g74 ( 
.A(n_48),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_SL g49 ( 
.A(n_17),
.B(n_15),
.Y(n_49)
);

INVx8_ASAP7_75t_L g50 ( 
.A(n_25),
.Y(n_50)
);

INVx5_ASAP7_75t_L g70 ( 
.A(n_50),
.Y(n_70)
);

INVx6_ASAP7_75t_L g51 ( 
.A(n_32),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g94 ( 
.A(n_51),
.Y(n_94)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_32),
.Y(n_52)
);

INVx6_ASAP7_75t_L g80 ( 
.A(n_52),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_18),
.B(n_7),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_L g83 ( 
.A(n_53),
.B(n_57),
.Y(n_83)
);

INVx3_ASAP7_75t_L g54 ( 
.A(n_39),
.Y(n_54)
);

INVx3_ASAP7_75t_L g71 ( 
.A(n_54),
.Y(n_71)
);

INVx3_ASAP7_75t_L g55 ( 
.A(n_39),
.Y(n_55)
);

INVx3_ASAP7_75t_L g76 ( 
.A(n_55),
.Y(n_76)
);

INVx3_ASAP7_75t_L g56 ( 
.A(n_19),
.Y(n_56)
);

INVx3_ASAP7_75t_L g98 ( 
.A(n_56),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g57 ( 
.A(n_21),
.B(n_7),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_35),
.Y(n_58)
);

INVx8_ASAP7_75t_L g81 ( 
.A(n_58),
.Y(n_81)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_35),
.Y(n_59)
);

INVx5_ASAP7_75t_L g89 ( 
.A(n_59),
.Y(n_89)
);

INVx3_ASAP7_75t_L g60 ( 
.A(n_19),
.Y(n_60)
);

INVx3_ASAP7_75t_L g106 ( 
.A(n_60),
.Y(n_106)
);

INVx6_ASAP7_75t_L g61 ( 
.A(n_35),
.Y(n_61)
);

INVx5_ASAP7_75t_L g102 ( 
.A(n_61),
.Y(n_102)
);

INVx2_ASAP7_75t_SL g62 ( 
.A(n_19),
.Y(n_62)
);

INVx4_ASAP7_75t_L g90 ( 
.A(n_62),
.Y(n_90)
);

INVx4_ASAP7_75t_L g63 ( 
.A(n_19),
.Y(n_63)
);

INVx3_ASAP7_75t_L g78 ( 
.A(n_63),
.Y(n_78)
);

BUFx12f_ASAP7_75t_L g67 ( 
.A(n_50),
.Y(n_67)
);

BUFx4f_ASAP7_75t_SL g122 ( 
.A(n_67),
.Y(n_122)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_43),
.Y(n_69)
);

INVx1_ASAP7_75t_SL g112 ( 
.A(n_69),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_L g130 ( 
.A(n_72),
.B(n_75),
.Y(n_130)
);

HB1xp67_ASAP7_75t_L g73 ( 
.A(n_62),
.Y(n_73)
);

INVxp67_ASAP7_75t_L g111 ( 
.A(n_73),
.Y(n_111)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_43),
.Y(n_75)
);

OAI22xp5_ASAP7_75t_SL g77 ( 
.A1(n_47),
.A2(n_41),
.B1(n_46),
.B2(n_51),
.Y(n_77)
);

AOI22xp5_ASAP7_75t_L g128 ( 
.A1(n_77),
.A2(n_79),
.B1(n_107),
.B2(n_4),
.Y(n_128)
);

OAI22xp5_ASAP7_75t_SL g79 ( 
.A1(n_61),
.A2(n_38),
.B1(n_36),
.B2(n_33),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_SL g84 ( 
.A(n_44),
.B(n_21),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_SL g120 ( 
.A(n_84),
.B(n_86),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_56),
.B(n_22),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g135 ( 
.A(n_85),
.B(n_95),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_SL g86 ( 
.A(n_44),
.B(n_22),
.Y(n_86)
);

BUFx12_ASAP7_75t_L g87 ( 
.A(n_44),
.Y(n_87)
);

BUFx5_ASAP7_75t_L g110 ( 
.A(n_87),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_L g88 ( 
.A(n_54),
.B(n_40),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_SL g123 ( 
.A(n_88),
.B(n_91),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_L g91 ( 
.A(n_55),
.B(n_28),
.Y(n_91)
);

AOI22xp33_ASAP7_75t_SL g92 ( 
.A1(n_62),
.A2(n_34),
.B1(n_36),
.B2(n_33),
.Y(n_92)
);

AOI22xp33_ASAP7_75t_SL g113 ( 
.A1(n_92),
.A2(n_96),
.B1(n_100),
.B2(n_29),
.Y(n_113)
);

AOI21xp33_ASAP7_75t_L g93 ( 
.A1(n_48),
.A2(n_40),
.B(n_20),
.Y(n_93)
);

AOI21xp33_ASAP7_75t_L g138 ( 
.A1(n_93),
.A2(n_6),
.B(n_9),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_60),
.B(n_20),
.Y(n_95)
);

AOI22xp33_ASAP7_75t_SL g96 ( 
.A1(n_63),
.A2(n_34),
.B1(n_36),
.B2(n_33),
.Y(n_96)
);

BUFx3_ASAP7_75t_L g97 ( 
.A(n_45),
.Y(n_97)
);

BUFx2_ASAP7_75t_L g119 ( 
.A(n_97),
.Y(n_119)
);

AOI22xp33_ASAP7_75t_SL g100 ( 
.A1(n_52),
.A2(n_34),
.B1(n_38),
.B2(n_37),
.Y(n_100)
);

AND2x2_ASAP7_75t_SL g101 ( 
.A(n_58),
.B(n_38),
.Y(n_101)
);

AND2x2_ASAP7_75t_L g139 ( 
.A(n_101),
.B(n_80),
.Y(n_139)
);

OR2x2_ASAP7_75t_L g103 ( 
.A(n_59),
.B(n_37),
.Y(n_103)
);

OR2x2_ASAP7_75t_L g136 ( 
.A(n_103),
.B(n_5),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_42),
.B(n_27),
.Y(n_104)
);

CKINVDCx16_ASAP7_75t_R g137 ( 
.A(n_104),
.Y(n_137)
);

INVx3_ASAP7_75t_L g105 ( 
.A(n_50),
.Y(n_105)
);

INVx4_ASAP7_75t_L g140 ( 
.A(n_105),
.Y(n_140)
);

AOI22xp33_ASAP7_75t_L g107 ( 
.A1(n_47),
.A2(n_24),
.B1(n_29),
.B2(n_30),
.Y(n_107)
);

CKINVDCx20_ASAP7_75t_R g108 ( 
.A(n_65),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_SL g166 ( 
.A(n_108),
.B(n_118),
.Y(n_166)
);

AO22x2_ASAP7_75t_L g109 ( 
.A1(n_102),
.A2(n_24),
.B1(n_30),
.B2(n_28),
.Y(n_109)
);

AND2x2_ASAP7_75t_L g141 ( 
.A(n_109),
.B(n_125),
.Y(n_141)
);

INVxp67_ASAP7_75t_L g145 ( 
.A(n_113),
.Y(n_145)
);

AO22x1_ASAP7_75t_SL g114 ( 
.A1(n_99),
.A2(n_27),
.B1(n_26),
.B2(n_17),
.Y(n_114)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_114),
.Y(n_147)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_90),
.Y(n_115)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_115),
.Y(n_157)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_90),
.Y(n_116)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_116),
.Y(n_170)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_64),
.Y(n_117)
);

INVx1_ASAP7_75t_SL g159 ( 
.A(n_117),
.Y(n_159)
);

CKINVDCx20_ASAP7_75t_R g118 ( 
.A(n_70),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_L g121 ( 
.A(n_82),
.B(n_107),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_L g151 ( 
.A(n_121),
.B(n_126),
.Y(n_151)
);

AOI22xp33_ASAP7_75t_L g124 ( 
.A1(n_89),
.A2(n_26),
.B1(n_31),
.B2(n_0),
.Y(n_124)
);

OAI22xp5_ASAP7_75t_L g160 ( 
.A1(n_124),
.A2(n_128),
.B1(n_81),
.B2(n_106),
.Y(n_160)
);

AO22x1_ASAP7_75t_SL g125 ( 
.A1(n_101),
.A2(n_2),
.B1(n_3),
.B2(n_4),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_L g126 ( 
.A(n_103),
.B(n_83),
.Y(n_126)
);

MAJIxp5_ASAP7_75t_L g127 ( 
.A(n_71),
.B(n_2),
.C(n_3),
.Y(n_127)
);

MAJIxp5_ASAP7_75t_L g161 ( 
.A(n_127),
.B(n_87),
.C(n_12),
.Y(n_161)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_66),
.Y(n_129)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_129),
.Y(n_155)
);

INVx2_ASAP7_75t_L g131 ( 
.A(n_94),
.Y(n_131)
);

INVx2_ASAP7_75t_L g152 ( 
.A(n_131),
.Y(n_152)
);

INVx2_ASAP7_75t_L g132 ( 
.A(n_94),
.Y(n_132)
);

INVx2_ASAP7_75t_L g163 ( 
.A(n_132),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_L g133 ( 
.A(n_66),
.B(n_5),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_L g158 ( 
.A(n_133),
.B(n_134),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_L g134 ( 
.A(n_102),
.B(n_5),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_L g143 ( 
.A(n_136),
.B(n_9),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_L g164 ( 
.A(n_138),
.B(n_10),
.Y(n_164)
);

AOI22xp5_ASAP7_75t_L g149 ( 
.A1(n_139),
.A2(n_74),
.B1(n_78),
.B2(n_76),
.Y(n_149)
);

BUFx6f_ASAP7_75t_L g142 ( 
.A(n_131),
.Y(n_142)
);

BUFx2_ASAP7_75t_L g175 ( 
.A(n_142),
.Y(n_175)
);

NOR2xp33_ASAP7_75t_L g190 ( 
.A(n_143),
.B(n_154),
.Y(n_190)
);

OAI22xp5_ASAP7_75t_SL g144 ( 
.A1(n_128),
.A2(n_100),
.B1(n_96),
.B2(n_92),
.Y(n_144)
);

AOI22xp5_ASAP7_75t_L g184 ( 
.A1(n_144),
.A2(n_146),
.B1(n_148),
.B2(n_122),
.Y(n_184)
);

OAI22xp5_ASAP7_75t_SL g146 ( 
.A1(n_121),
.A2(n_80),
.B1(n_68),
.B2(n_97),
.Y(n_146)
);

OAI22xp5_ASAP7_75t_SL g148 ( 
.A1(n_123),
.A2(n_68),
.B1(n_89),
.B2(n_81),
.Y(n_148)
);

INVxp67_ASAP7_75t_L g174 ( 
.A(n_149),
.Y(n_174)
);

XOR2xp5_ASAP7_75t_L g150 ( 
.A(n_126),
.B(n_78),
.Y(n_150)
);

MAJIxp5_ASAP7_75t_L g198 ( 
.A(n_150),
.B(n_110),
.C(n_14),
.Y(n_198)
);

AOI21xp5_ASAP7_75t_L g153 ( 
.A1(n_139),
.A2(n_74),
.B(n_105),
.Y(n_153)
);

AOI21xp5_ASAP7_75t_L g194 ( 
.A1(n_153),
.A2(n_169),
.B(n_122),
.Y(n_194)
);

NOR2xp33_ASAP7_75t_L g154 ( 
.A(n_137),
.B(n_98),
.Y(n_154)
);

CKINVDCx20_ASAP7_75t_R g156 ( 
.A(n_111),
.Y(n_156)
);

NOR2xp33_ASAP7_75t_L g195 ( 
.A(n_156),
.B(n_164),
.Y(n_195)
);

OAI22xp5_ASAP7_75t_L g176 ( 
.A1(n_160),
.A2(n_172),
.B1(n_112),
.B2(n_117),
.Y(n_176)
);

XNOR2xp5_ASAP7_75t_L g173 ( 
.A(n_161),
.B(n_127),
.Y(n_173)
);

A2O1A1Ixp33_ASAP7_75t_L g162 ( 
.A1(n_120),
.A2(n_87),
.B(n_12),
.C(n_13),
.Y(n_162)
);

OAI21xp5_ASAP7_75t_L g178 ( 
.A1(n_162),
.A2(n_125),
.B(n_134),
.Y(n_178)
);

INVx3_ASAP7_75t_L g165 ( 
.A(n_140),
.Y(n_165)
);

INVxp67_ASAP7_75t_L g188 ( 
.A(n_165),
.Y(n_188)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_129),
.Y(n_167)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_167),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_L g168 ( 
.A(n_133),
.B(n_70),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_L g179 ( 
.A(n_168),
.B(n_125),
.Y(n_179)
);

AOI21xp5_ASAP7_75t_L g169 ( 
.A1(n_139),
.A2(n_67),
.B(n_13),
.Y(n_169)
);

NOR2xp33_ASAP7_75t_L g171 ( 
.A(n_130),
.B(n_67),
.Y(n_171)
);

NOR2xp33_ASAP7_75t_L g197 ( 
.A(n_171),
.B(n_122),
.Y(n_197)
);

AOI22xp5_ASAP7_75t_L g172 ( 
.A1(n_136),
.A2(n_10),
.B1(n_13),
.B2(n_14),
.Y(n_172)
);

XOR2xp5_ASAP7_75t_L g217 ( 
.A(n_173),
.B(n_198),
.Y(n_217)
);

AND2x2_ASAP7_75t_L g214 ( 
.A(n_176),
.B(n_183),
.Y(n_214)
);

OAI21xp5_ASAP7_75t_SL g177 ( 
.A1(n_147),
.A2(n_135),
.B(n_112),
.Y(n_177)
);

OAI21xp5_ASAP7_75t_L g203 ( 
.A1(n_177),
.A2(n_193),
.B(n_200),
.Y(n_203)
);

NOR2xp33_ASAP7_75t_L g212 ( 
.A(n_178),
.B(n_191),
.Y(n_212)
);

NAND2xp5_ASAP7_75t_L g211 ( 
.A(n_179),
.B(n_194),
.Y(n_211)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_155),
.Y(n_181)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_181),
.Y(n_205)
);

AOI22xp33_ASAP7_75t_L g182 ( 
.A1(n_147),
.A2(n_109),
.B1(n_114),
.B2(n_132),
.Y(n_182)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_182),
.Y(n_218)
);

AO22x1_ASAP7_75t_L g183 ( 
.A1(n_141),
.A2(n_109),
.B1(n_114),
.B2(n_116),
.Y(n_183)
);

AOI22xp5_ASAP7_75t_L g207 ( 
.A1(n_184),
.A2(n_187),
.B1(n_201),
.B2(n_169),
.Y(n_207)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_159),
.Y(n_185)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_185),
.Y(n_202)
);

XOR2xp5_ASAP7_75t_L g186 ( 
.A(n_150),
.B(n_115),
.Y(n_186)
);

XNOR2xp5_ASAP7_75t_L g204 ( 
.A(n_186),
.B(n_149),
.Y(n_204)
);

OAI22xp5_ASAP7_75t_L g187 ( 
.A1(n_151),
.A2(n_109),
.B1(n_140),
.B2(n_119),
.Y(n_187)
);

INVxp67_ASAP7_75t_L g189 ( 
.A(n_153),
.Y(n_189)
);

HB1xp67_ASAP7_75t_L g208 ( 
.A(n_189),
.Y(n_208)
);

INVxp67_ASAP7_75t_L g191 ( 
.A(n_165),
.Y(n_191)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_159),
.Y(n_192)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_192),
.Y(n_209)
);

AOI21xp5_ASAP7_75t_SL g193 ( 
.A1(n_141),
.A2(n_111),
.B(n_119),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_L g196 ( 
.A(n_158),
.B(n_151),
.Y(n_196)
);

NAND2xp5_ASAP7_75t_L g216 ( 
.A(n_196),
.B(n_157),
.Y(n_216)
);

NAND2xp5_ASAP7_75t_SL g213 ( 
.A(n_197),
.B(n_199),
.Y(n_213)
);

NOR2xp33_ASAP7_75t_L g199 ( 
.A(n_164),
.B(n_15),
.Y(n_199)
);

AOI22xp33_ASAP7_75t_SL g200 ( 
.A1(n_145),
.A2(n_110),
.B1(n_144),
.B2(n_148),
.Y(n_200)
);

OAI22xp5_ASAP7_75t_SL g201 ( 
.A1(n_141),
.A2(n_145),
.B1(n_168),
.B2(n_158),
.Y(n_201)
);

XOR2xp5_ASAP7_75t_L g225 ( 
.A(n_204),
.B(n_186),
.Y(n_225)
);

CKINVDCx20_ASAP7_75t_R g206 ( 
.A(n_188),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_L g231 ( 
.A(n_206),
.B(n_216),
.Y(n_231)
);

AOI22xp5_ASAP7_75t_L g224 ( 
.A1(n_207),
.A2(n_215),
.B1(n_220),
.B2(n_183),
.Y(n_224)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_180),
.Y(n_210)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_210),
.Y(n_226)
);

AOI22xp5_ASAP7_75t_L g215 ( 
.A1(n_201),
.A2(n_146),
.B1(n_162),
.B2(n_166),
.Y(n_215)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_180),
.Y(n_219)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_219),
.Y(n_232)
);

OAI22xp5_ASAP7_75t_SL g220 ( 
.A1(n_184),
.A2(n_172),
.B1(n_152),
.B2(n_163),
.Y(n_220)
);

NAND2xp5_ASAP7_75t_L g221 ( 
.A(n_196),
.B(n_161),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_L g227 ( 
.A(n_221),
.B(n_223),
.Y(n_227)
);

NAND2xp5_ASAP7_75t_SL g222 ( 
.A(n_177),
.B(n_157),
.Y(n_222)
);

INVxp67_ASAP7_75t_SL g239 ( 
.A(n_222),
.Y(n_239)
);

NAND2xp5_ASAP7_75t_L g223 ( 
.A(n_179),
.B(n_170),
.Y(n_223)
);

HB1xp67_ASAP7_75t_L g242 ( 
.A(n_224),
.Y(n_242)
);

XNOR2xp5_ASAP7_75t_SL g249 ( 
.A(n_225),
.B(n_235),
.Y(n_249)
);

OAI21xp5_ASAP7_75t_SL g228 ( 
.A1(n_203),
.A2(n_193),
.B(n_194),
.Y(n_228)
);

NAND2xp5_ASAP7_75t_SL g254 ( 
.A(n_228),
.B(n_241),
.Y(n_254)
);

AOI22xp5_ASAP7_75t_L g229 ( 
.A1(n_214),
.A2(n_183),
.B1(n_174),
.B2(n_189),
.Y(n_229)
);

OAI22xp5_ASAP7_75t_SL g247 ( 
.A1(n_229),
.A2(n_234),
.B1(n_240),
.B2(n_215),
.Y(n_247)
);

AOI21xp5_ASAP7_75t_L g230 ( 
.A1(n_203),
.A2(n_178),
.B(n_174),
.Y(n_230)
);

NAND2xp5_ASAP7_75t_L g251 ( 
.A(n_230),
.B(n_236),
.Y(n_251)
);

XOR2xp5_ASAP7_75t_L g233 ( 
.A(n_217),
.B(n_221),
.Y(n_233)
);

MAJIxp5_ASAP7_75t_L g244 ( 
.A(n_233),
.B(n_235),
.C(n_237),
.Y(n_244)
);

AOI22xp5_ASAP7_75t_L g234 ( 
.A1(n_214),
.A2(n_173),
.B1(n_195),
.B2(n_192),
.Y(n_234)
);

XOR2xp5_ASAP7_75t_L g235 ( 
.A(n_217),
.B(n_198),
.Y(n_235)
);

AOI21xp5_ASAP7_75t_L g236 ( 
.A1(n_211),
.A2(n_191),
.B(n_188),
.Y(n_236)
);

MAJIxp5_ASAP7_75t_L g237 ( 
.A(n_204),
.B(n_181),
.C(n_185),
.Y(n_237)
);

INVxp67_ASAP7_75t_L g238 ( 
.A(n_208),
.Y(n_238)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_238),
.Y(n_243)
);

AOI22xp5_ASAP7_75t_L g240 ( 
.A1(n_214),
.A2(n_190),
.B1(n_175),
.B2(n_170),
.Y(n_240)
);

OAI21xp5_ASAP7_75t_SL g241 ( 
.A1(n_211),
.A2(n_152),
.B(n_163),
.Y(n_241)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_226),
.Y(n_245)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_245),
.Y(n_256)
);

MAJIxp5_ASAP7_75t_L g246 ( 
.A(n_233),
.B(n_216),
.C(n_223),
.Y(n_246)
);

MAJIxp5_ASAP7_75t_L g257 ( 
.A(n_246),
.B(n_250),
.C(n_237),
.Y(n_257)
);

NOR2xp33_ASAP7_75t_L g263 ( 
.A(n_247),
.B(n_207),
.Y(n_263)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_232),
.Y(n_248)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_248),
.Y(n_259)
);

XNOR2x1_ASAP7_75t_L g258 ( 
.A(n_249),
.B(n_253),
.Y(n_258)
);

XOR2xp5_ASAP7_75t_L g250 ( 
.A(n_225),
.B(n_234),
.Y(n_250)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_231),
.Y(n_252)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_252),
.Y(n_261)
);

AOI22xp5_ASAP7_75t_SL g253 ( 
.A1(n_239),
.A2(n_212),
.B1(n_218),
.B2(n_220),
.Y(n_253)
);

NAND4xp25_ASAP7_75t_L g255 ( 
.A(n_251),
.B(n_230),
.C(n_240),
.D(n_224),
.Y(n_255)
);

NOR2xp33_ASAP7_75t_L g265 ( 
.A(n_255),
.B(n_264),
.Y(n_265)
);

XNOR2xp5_ASAP7_75t_L g271 ( 
.A(n_257),
.B(n_241),
.Y(n_271)
);

MAJIxp5_ASAP7_75t_L g260 ( 
.A(n_244),
.B(n_227),
.C(n_236),
.Y(n_260)
);

MAJIxp5_ASAP7_75t_L g267 ( 
.A(n_260),
.B(n_244),
.C(n_250),
.Y(n_267)
);

AOI31xp67_ASAP7_75t_L g262 ( 
.A1(n_246),
.A2(n_229),
.A3(n_227),
.B(n_228),
.Y(n_262)
);

AOI22xp5_ASAP7_75t_L g272 ( 
.A1(n_262),
.A2(n_263),
.B1(n_254),
.B2(n_238),
.Y(n_272)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_243),
.Y(n_264)
);

BUFx6f_ASAP7_75t_L g266 ( 
.A(n_261),
.Y(n_266)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_266),
.Y(n_277)
);

MAJIxp5_ASAP7_75t_L g274 ( 
.A(n_267),
.B(n_271),
.C(n_272),
.Y(n_274)
);

MAJIxp5_ASAP7_75t_L g268 ( 
.A(n_257),
.B(n_249),
.C(n_213),
.Y(n_268)
);

NAND2xp5_ASAP7_75t_L g276 ( 
.A(n_268),
.B(n_269),
.Y(n_276)
);

NOR2xp33_ASAP7_75t_L g269 ( 
.A(n_260),
.B(n_247),
.Y(n_269)
);

OAI22x1_ASAP7_75t_L g270 ( 
.A1(n_262),
.A2(n_242),
.B1(n_251),
.B2(n_253),
.Y(n_270)
);

AOI22xp33_ASAP7_75t_SL g273 ( 
.A1(n_270),
.A2(n_255),
.B1(n_258),
.B2(n_256),
.Y(n_273)
);

NOR2xp33_ASAP7_75t_L g281 ( 
.A(n_273),
.B(n_270),
.Y(n_281)
);

MAJIxp5_ASAP7_75t_L g275 ( 
.A(n_267),
.B(n_258),
.C(n_209),
.Y(n_275)
);

NAND2xp5_ASAP7_75t_SL g280 ( 
.A(n_275),
.B(n_278),
.Y(n_280)
);

NOR2xp33_ASAP7_75t_SL g278 ( 
.A(n_265),
.B(n_259),
.Y(n_278)
);

NOR2xp33_ASAP7_75t_SL g279 ( 
.A(n_276),
.B(n_266),
.Y(n_279)
);

NOR2xp33_ASAP7_75t_L g285 ( 
.A(n_279),
.B(n_219),
.Y(n_285)
);

OAI21x1_ASAP7_75t_L g283 ( 
.A1(n_281),
.A2(n_282),
.B(n_277),
.Y(n_283)
);

OR2x2_ASAP7_75t_L g282 ( 
.A(n_274),
.B(n_210),
.Y(n_282)
);

NAND2xp5_ASAP7_75t_L g286 ( 
.A(n_283),
.B(n_284),
.Y(n_286)
);

OAI21x1_ASAP7_75t_L g284 ( 
.A1(n_282),
.A2(n_273),
.B(n_202),
.Y(n_284)
);

NAND2xp5_ASAP7_75t_SL g287 ( 
.A(n_285),
.B(n_205),
.Y(n_287)
);

INVxp67_ASAP7_75t_L g288 ( 
.A(n_287),
.Y(n_288)
);

AOI22xp5_ASAP7_75t_L g289 ( 
.A1(n_288),
.A2(n_286),
.B1(n_280),
.B2(n_202),
.Y(n_289)
);

XOR2xp5_ASAP7_75t_L g290 ( 
.A(n_289),
.B(n_209),
.Y(n_290)
);


endmodule