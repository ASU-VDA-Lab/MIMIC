module real_jpeg_4531_n_29 (n_17, n_8, n_0, n_157, n_21, n_2, n_10, n_9, n_12, n_156, n_24, n_6, n_159, n_28, n_161, n_162, n_23, n_11, n_14, n_160, n_25, n_163, n_7, n_22, n_18, n_3, n_5, n_4, n_1, n_26, n_27, n_20, n_19, n_164, n_158, n_16, n_15, n_13, n_155, n_29);

input n_17;
input n_8;
input n_0;
input n_157;
input n_21;
input n_2;
input n_10;
input n_9;
input n_12;
input n_156;
input n_24;
input n_6;
input n_159;
input n_28;
input n_161;
input n_162;
input n_23;
input n_11;
input n_14;
input n_160;
input n_25;
input n_163;
input n_7;
input n_22;
input n_18;
input n_3;
input n_5;
input n_4;
input n_1;
input n_26;
input n_27;
input n_20;
input n_19;
input n_164;
input n_158;
input n_16;
input n_15;
input n_13;
input n_155;

output n_29;

wire n_108;
wire n_54;
wire n_37;
wire n_73;
wire n_35;
wire n_38;
wire n_91;
wire n_49;
wire n_114;
wire n_68;
wire n_146;
wire n_83;
wire n_78;
wire n_104;
wire n_153;
wire n_64;
wire n_47;
wire n_131;
wire n_87;
wire n_40;
wire n_105;
wire n_115;
wire n_98;
wire n_56;
wire n_48;
wire n_140;
wire n_126;
wire n_113;
wire n_120;
wire n_93;
wire n_141;
wire n_95;
wire n_65;
wire n_33;
wire n_139;
wire n_142;
wire n_76;
wire n_67;
wire n_79;
wire n_107;
wire n_147;
wire n_66;
wire n_136;
wire n_44;
wire n_62;
wire n_121;
wire n_106;
wire n_45;
wire n_112;
wire n_42;
wire n_145;
wire n_77;
wire n_109;
wire n_39;
wire n_122;
wire n_94;
wire n_148;
wire n_118;
wire n_123;
wire n_116;
wire n_50;
wire n_143;
wire n_69;
wire n_31;
wire n_137;
wire n_129;
wire n_135;
wire n_152;
wire n_134;
wire n_72;
wire n_151;
wire n_100;
wire n_51;
wire n_71;
wire n_90;
wire n_61;
wire n_110;
wire n_117;
wire n_99;
wire n_86;
wire n_70;
wire n_41;
wire n_74;
wire n_80;
wire n_32;
wire n_150;
wire n_30;
wire n_149;
wire n_144;
wire n_130;
wire n_103;
wire n_43;
wire n_57;
wire n_84;
wire n_82;
wire n_111;
wire n_132;
wire n_125;
wire n_55;
wire n_58;
wire n_52;
wire n_63;
wire n_124;
wire n_92;
wire n_75;
wire n_97;
wire n_34;
wire n_60;
wire n_46;
wire n_88;
wire n_59;
wire n_128;
wire n_133;
wire n_138;
wire n_53;
wire n_127;
wire n_119;
wire n_36;
wire n_102;
wire n_81;
wire n_85;
wire n_101;
wire n_96;
wire n_89;

BUFx5_ASAP7_75t_L g39 ( 
.A(n_0),
.Y(n_39)
);

INVx5_ASAP7_75t_L g44 ( 
.A(n_0),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_0),
.Y(n_62)
);

BUFx5_ASAP7_75t_L g66 ( 
.A(n_0),
.Y(n_66)
);

OR2x2_ASAP7_75t_L g78 ( 
.A(n_0),
.B(n_79),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_SL g45 ( 
.A(n_1),
.B(n_46),
.Y(n_45)
);

NAND2xp5_ASAP7_75t_L g108 ( 
.A(n_1),
.B(n_46),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_SL g63 ( 
.A(n_2),
.B(n_64),
.Y(n_63)
);

AND2x2_ASAP7_75t_L g91 ( 
.A(n_2),
.B(n_64),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_3),
.B(n_51),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_L g107 ( 
.A(n_3),
.B(n_51),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_4),
.B(n_100),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g102 ( 
.A(n_4),
.B(n_100),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_SL g123 ( 
.A(n_5),
.B(n_124),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_L g133 ( 
.A(n_5),
.B(n_124),
.Y(n_133)
);

CKINVDCx20_ASAP7_75t_R g128 ( 
.A(n_6),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_SL g140 ( 
.A(n_7),
.B(n_141),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_L g145 ( 
.A(n_7),
.B(n_141),
.Y(n_145)
);

CKINVDCx20_ASAP7_75t_R g121 ( 
.A(n_8),
.Y(n_121)
);

AND2x2_ASAP7_75t_L g74 ( 
.A(n_9),
.B(n_75),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_SL g34 ( 
.A(n_10),
.B(n_35),
.Y(n_34)
);

AND2x2_ASAP7_75t_L g109 ( 
.A(n_10),
.B(n_35),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_11),
.B(n_83),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_L g87 ( 
.A(n_11),
.B(n_83),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g147 ( 
.A(n_12),
.B(n_148),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_L g153 ( 
.A(n_12),
.B(n_148),
.Y(n_153)
);

OR2x2_ASAP7_75t_L g112 ( 
.A(n_13),
.B(n_113),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_L g132 ( 
.A(n_13),
.B(n_113),
.Y(n_132)
);

CKINVDCx20_ASAP7_75t_R g142 ( 
.A(n_14),
.Y(n_142)
);

CKINVDCx20_ASAP7_75t_R g114 ( 
.A(n_15),
.Y(n_114)
);

CKINVDCx20_ASAP7_75t_R g125 ( 
.A(n_16),
.Y(n_125)
);

CKINVDCx20_ASAP7_75t_R g97 ( 
.A(n_17),
.Y(n_97)
);

CKINVDCx20_ASAP7_75t_R g149 ( 
.A(n_18),
.Y(n_149)
);

CKINVDCx20_ASAP7_75t_R g139 ( 
.A(n_19),
.Y(n_139)
);

CKINVDCx20_ASAP7_75t_R g129 ( 
.A(n_20),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_SL g137 ( 
.A(n_21),
.B(n_138),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_L g144 ( 
.A(n_21),
.B(n_138),
.Y(n_144)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_22),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_23),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g40 ( 
.A(n_24),
.B(n_41),
.Y(n_40)
);

AND2x2_ASAP7_75t_L g111 ( 
.A(n_24),
.B(n_41),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_SL g58 ( 
.A(n_25),
.B(n_59),
.Y(n_58)
);

AND2x2_ASAP7_75t_L g90 ( 
.A(n_25),
.B(n_59),
.Y(n_90)
);

CKINVDCx20_ASAP7_75t_R g71 ( 
.A(n_26),
.Y(n_71)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_27),
.Y(n_80)
);

CKINVDCx20_ASAP7_75t_R g119 ( 
.A(n_28),
.Y(n_119)
);

XOR2xp5_ASAP7_75t_L g29 ( 
.A(n_30),
.B(n_146),
.Y(n_29)
);

AOI21xp5_ASAP7_75t_L g30 ( 
.A1(n_31),
.A2(n_136),
.B(n_143),
.Y(n_30)
);

OAI21xp5_ASAP7_75t_SL g31 ( 
.A1(n_32),
.A2(n_117),
.B(n_130),
.Y(n_31)
);

A2O1A1Ixp33_ASAP7_75t_L g32 ( 
.A1(n_33),
.A2(n_54),
.B(n_103),
.C(n_112),
.Y(n_32)
);

NOR4xp25_ASAP7_75t_L g33 ( 
.A(n_34),
.B(n_40),
.C(n_45),
.D(n_50),
.Y(n_33)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_34),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g35 ( 
.A(n_36),
.B(n_37),
.Y(n_35)
);

INVx4_ASAP7_75t_L g37 ( 
.A(n_38),
.Y(n_37)
);

INVx2_ASAP7_75t_L g38 ( 
.A(n_39),
.Y(n_38)
);

OR2x2_ASAP7_75t_L g69 ( 
.A(n_39),
.B(n_70),
.Y(n_69)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_40),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_L g41 ( 
.A(n_42),
.B(n_43),
.Y(n_41)
);

BUFx3_ASAP7_75t_L g53 ( 
.A(n_43),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_43),
.B(n_76),
.Y(n_75)
);

INVx11_ASAP7_75t_L g43 ( 
.A(n_44),
.Y(n_43)
);

BUFx3_ASAP7_75t_L g49 ( 
.A(n_44),
.Y(n_49)
);

INVx5_ASAP7_75t_L g96 ( 
.A(n_44),
.Y(n_96)
);

OAI21xp5_ASAP7_75t_L g106 ( 
.A1(n_45),
.A2(n_107),
.B(n_108),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g46 ( 
.A(n_47),
.B(n_48),
.Y(n_46)
);

INVx3_ASAP7_75t_L g48 ( 
.A(n_49),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g51 ( 
.A(n_52),
.B(n_53),
.Y(n_51)
);

CKINVDCx20_ASAP7_75t_R g151 ( 
.A(n_53),
.Y(n_151)
);

OAI21x1_ASAP7_75t_L g54 ( 
.A1(n_55),
.A2(n_99),
.B(n_102),
.Y(n_54)
);

AOI21xp5_ASAP7_75t_L g55 ( 
.A1(n_56),
.A2(n_92),
.B(n_98),
.Y(n_55)
);

AO221x1_ASAP7_75t_L g56 ( 
.A1(n_57),
.A2(n_67),
.B1(n_89),
.B2(n_90),
.C(n_91),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g57 ( 
.A(n_58),
.B(n_63),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_60),
.B(n_61),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_61),
.B(n_101),
.Y(n_100)
);

INVx3_ASAP7_75t_L g116 ( 
.A(n_61),
.Y(n_116)
);

BUFx12f_ASAP7_75t_L g61 ( 
.A(n_62),
.Y(n_61)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_63),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_65),
.B(n_66),
.Y(n_64)
);

INVx2_ASAP7_75t_L g85 ( 
.A(n_66),
.Y(n_85)
);

AO21x1_ASAP7_75t_L g67 ( 
.A1(n_68),
.A2(n_72),
.B(n_88),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_SL g68 ( 
.A(n_69),
.B(n_71),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_69),
.B(n_71),
.Y(n_88)
);

OAI21xp5_ASAP7_75t_SL g72 ( 
.A1(n_73),
.A2(n_82),
.B(n_87),
.Y(n_72)
);

AOI21xp5_ASAP7_75t_L g73 ( 
.A1(n_74),
.A2(n_77),
.B(n_81),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_SL g77 ( 
.A(n_78),
.B(n_80),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_78),
.B(n_80),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_SL g83 ( 
.A(n_84),
.B(n_86),
.Y(n_83)
);

INVx3_ASAP7_75t_L g84 ( 
.A(n_85),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_SL g92 ( 
.A(n_93),
.B(n_97),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_93),
.B(n_97),
.Y(n_98)
);

OR2x2_ASAP7_75t_L g93 ( 
.A(n_94),
.B(n_95),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_95),
.B(n_125),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_L g138 ( 
.A(n_95),
.B(n_139),
.Y(n_138)
);

BUFx12_ASAP7_75t_L g95 ( 
.A(n_96),
.Y(n_95)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_104),
.Y(n_103)
);

A2O1A1O1Ixp25_ASAP7_75t_L g104 ( 
.A1(n_105),
.A2(n_106),
.B(n_109),
.C(n_110),
.D(n_111),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_L g113 ( 
.A(n_114),
.B(n_115),
.Y(n_113)
);

OR2x2_ASAP7_75t_L g120 ( 
.A(n_115),
.B(n_121),
.Y(n_120)
);

OR2x2_ASAP7_75t_L g127 ( 
.A(n_115),
.B(n_128),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_L g141 ( 
.A(n_115),
.B(n_142),
.Y(n_141)
);

INVx8_ASAP7_75t_L g115 ( 
.A(n_116),
.Y(n_115)
);

NAND3xp33_ASAP7_75t_L g117 ( 
.A(n_118),
.B(n_122),
.C(n_126),
.Y(n_117)
);

A2O1A1O1Ixp25_ASAP7_75t_L g130 ( 
.A1(n_118),
.A2(n_126),
.B(n_131),
.C(n_134),
.D(n_135),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_L g118 ( 
.A(n_119),
.B(n_120),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_L g135 ( 
.A(n_119),
.B(n_120),
.Y(n_135)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_123),
.Y(n_122)
);

OAI21xp5_ASAP7_75t_L g131 ( 
.A1(n_123),
.A2(n_132),
.B(n_133),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_SL g126 ( 
.A(n_127),
.B(n_129),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_L g134 ( 
.A(n_127),
.B(n_129),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_L g136 ( 
.A(n_137),
.B(n_140),
.Y(n_136)
);

OAI21xp5_ASAP7_75t_L g143 ( 
.A1(n_140),
.A2(n_144),
.B(n_145),
.Y(n_143)
);

NOR2xp33_ASAP7_75t_L g146 ( 
.A(n_147),
.B(n_152),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_L g148 ( 
.A(n_149),
.B(n_150),
.Y(n_148)
);

INVx3_ASAP7_75t_L g150 ( 
.A(n_151),
.Y(n_150)
);

INVxp33_ASAP7_75t_L g152 ( 
.A(n_153),
.Y(n_152)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_155),
.Y(n_47)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_156),
.Y(n_52)
);

CKINVDCx20_ASAP7_75t_R g60 ( 
.A(n_157),
.Y(n_60)
);

CKINVDCx20_ASAP7_75t_R g65 ( 
.A(n_158),
.Y(n_65)
);

CKINVDCx20_ASAP7_75t_R g70 ( 
.A(n_159),
.Y(n_70)
);

CKINVDCx20_ASAP7_75t_R g76 ( 
.A(n_160),
.Y(n_76)
);

CKINVDCx20_ASAP7_75t_R g79 ( 
.A(n_161),
.Y(n_79)
);

CKINVDCx20_ASAP7_75t_R g86 ( 
.A(n_162),
.Y(n_86)
);

CKINVDCx20_ASAP7_75t_R g94 ( 
.A(n_163),
.Y(n_94)
);

CKINVDCx20_ASAP7_75t_R g101 ( 
.A(n_164),
.Y(n_101)
);


endmodule