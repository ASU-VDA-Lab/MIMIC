module fake_aes_4709_n_39 (n_1, n_2, n_6, n_4, n_3, n_9, n_5, n_7, n_10, n_8, n_0, n_39);
input n_1;
input n_2;
input n_6;
input n_4;
input n_3;
input n_9;
input n_5;
input n_7;
input n_10;
input n_8;
input n_0;
output n_39;
wire n_20;
wire n_38;
wire n_36;
wire n_37;
wire n_34;
wire n_23;
wire n_28;
wire n_31;
wire n_22;
wire n_11;
wire n_25;
wire n_16;
wire n_26;
wire n_13;
wire n_33;
wire n_30;
wire n_18;
wire n_32;
wire n_35;
wire n_12;
wire n_17;
wire n_14;
wire n_15;
wire n_24;
wire n_19;
wire n_21;
wire n_29;
wire n_27;
NAND2xp5_ASAP7_75t_L g11 ( .A(n_2), .B(n_4), .Y(n_11) );
INVx1_ASAP7_75t_L g12 ( .A(n_0), .Y(n_12) );
CKINVDCx5p33_ASAP7_75t_R g13 ( .A(n_2), .Y(n_13) );
INVx1_ASAP7_75t_L g14 ( .A(n_7), .Y(n_14) );
NAND2xp5_ASAP7_75t_L g15 ( .A(n_5), .B(n_6), .Y(n_15) );
INVx1_ASAP7_75t_L g16 ( .A(n_10), .Y(n_16) );
CKINVDCx5p33_ASAP7_75t_R g17 ( .A(n_3), .Y(n_17) );
INVx2_ASAP7_75t_L g18 ( .A(n_6), .Y(n_18) );
INVx2_ASAP7_75t_SL g19 ( .A(n_14), .Y(n_19) );
BUFx2_ASAP7_75t_L g20 ( .A(n_13), .Y(n_20) );
INVx2_ASAP7_75t_L g21 ( .A(n_16), .Y(n_21) );
AND2x2_ASAP7_75t_L g22 ( .A(n_18), .B(n_0), .Y(n_22) );
BUFx4f_ASAP7_75t_L g23 ( .A(n_12), .Y(n_23) );
BUFx8_ASAP7_75t_L g24 ( .A(n_18), .Y(n_24) );
AOI221xp5_ASAP7_75t_L g25 ( .A1(n_20), .A2(n_13), .B1(n_17), .B2(n_12), .C(n_15), .Y(n_25) );
OAI22xp5_ASAP7_75t_L g26 ( .A1(n_23), .A2(n_17), .B1(n_11), .B2(n_4), .Y(n_26) );
HB1xp67_ASAP7_75t_L g27 ( .A(n_24), .Y(n_27) );
OAI22xp33_ASAP7_75t_L g28 ( .A1(n_27), .A2(n_23), .B1(n_19), .B2(n_21), .Y(n_28) );
OAI322xp33_ASAP7_75t_L g29 ( .A1(n_26), .A2(n_19), .A3(n_21), .B1(n_22), .B2(n_23), .C1(n_24), .C2(n_5), .Y(n_29) );
INVx1_ASAP7_75t_L g30 ( .A(n_29), .Y(n_30) );
AND2x2_ASAP7_75t_SL g31 ( .A(n_28), .B(n_25), .Y(n_31) );
AOI21xp33_ASAP7_75t_L g32 ( .A1(n_31), .A2(n_24), .B(n_3), .Y(n_32) );
NOR2xp33_ASAP7_75t_L g33 ( .A(n_31), .B(n_1), .Y(n_33) );
XOR2xp5_ASAP7_75t_L g34 ( .A(n_33), .B(n_30), .Y(n_34) );
NOR2x1_ASAP7_75t_L g35 ( .A(n_32), .B(n_30), .Y(n_35) );
XNOR2x1_ASAP7_75t_L g36 ( .A(n_34), .B(n_35), .Y(n_36) );
CKINVDCx14_ASAP7_75t_R g37 ( .A(n_34), .Y(n_37) );
OR2x2_ASAP7_75t_L g38 ( .A(n_36), .B(n_1), .Y(n_38) );
OAI221xp5_ASAP7_75t_R g39 ( .A1(n_38), .A2(n_37), .B1(n_31), .B2(n_9), .C(n_8), .Y(n_39) );
endmodule