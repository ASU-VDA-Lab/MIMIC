module real_jpeg_4012_n_18 (n_17, n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_16, n_3, n_10, n_9, n_18);

input n_17;
input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_16;
input n_3;
input n_10;
input n_9;

output n_18;

wire n_384;
wire n_37;
wire n_430;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_460;
wire n_300;
wire n_415;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_446;
wire n_199;
wire n_95;
wire n_441;
wire n_238;
wire n_67;
wire n_350;
wire n_235;
wire n_107;
wire n_369;
wire n_498;
wire n_471;
wire n_376;
wire n_354;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_490;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_355;
wire n_123;
wire n_463;
wire n_425;
wire n_455;
wire n_462;
wire n_50;
wire n_409;
wire n_485;
wire n_186;
wire n_137;
wire n_491;
wire n_72;
wire n_440;
wire n_171;
wire n_151;
wire n_272;
wire n_461;
wire n_198;
wire n_203;
wire n_500;
wire n_23;
wire n_362;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_326;
wire n_339;
wire n_80;
wire n_30;
wire n_332;
wire n_149;
wire n_366;
wire n_328;
wire n_456;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_499;
wire n_58;
wire n_52;
wire n_466;
wire n_353;
wire n_453;
wire n_230;
wire n_417;
wire n_428;
wire n_128;
wire n_202;
wire n_216;
wire n_483;
wire n_367;
wire n_127;
wire n_356;
wire n_365;
wire n_464;
wire n_423;
wire n_36;
wire n_102;
wire n_81;
wire n_101;
wire n_422;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_348;
wire n_473;
wire n_252;
wire n_363;
wire n_310;
wire n_345;
wire n_78;
wire n_83;
wire n_288;
wire n_221;
wire n_393;
wire n_489;
wire n_104;
wire n_153;
wire n_443;
wire n_337;
wire n_131;
wire n_439;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_378;
wire n_469;
wire n_200;
wire n_432;
wire n_465;
wire n_335;
wire n_214;
wire n_113;
wire n_251;
wire n_459;
wire n_139;
wire n_33;
wire n_175;
wire n_338;
wire n_488;
wire n_156;
wire n_387;
wire n_434;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_390;
wire n_77;
wire n_399;
wire n_219;
wire n_470;
wire n_372;
wire n_122;
wire n_19;
wire n_262;
wire n_334;
wire n_383;
wire n_246;
wire n_21;
wire n_476;
wire n_69;
wire n_31;
wire n_426;
wire n_154;
wire n_495;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_371;
wire n_410;
wire n_421;
wire n_195;
wire n_110;
wire n_289;
wire n_117;
wire n_193;
wire n_382;
wire n_411;
wire n_20;
wire n_314;
wire n_278;
wire n_103;
wire n_232;
wire n_448;
wire n_212;
wire n_284;
wire n_402;
wire n_478;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_452;
wire n_213;
wire n_25;
wire n_480;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_407;
wire n_419;
wire n_386;
wire n_341;
wire n_331;
wire n_49;
wire n_68;
wire n_497;
wire n_395;
wire n_146;
wire n_496;
wire n_286;
wire n_166;
wire n_215;
wire n_176;
wire n_323;
wire n_312;
wire n_325;
wire n_316;
wire n_307;
wire n_161;
wire n_207;
wire n_431;
wire n_420;
wire n_357;
wire n_237;
wire n_445;
wire n_173;
wire n_115;
wire n_474;
wire n_184;
wire n_164;
wire n_380;
wire n_414;
wire n_140;
wire n_126;
wire n_342;
wire n_120;
wire n_155;
wire n_412;
wire n_405;
wire n_319;
wire n_93;
wire n_487;
wire n_242;
wire n_493;
wire n_142;
wire n_397;
wire n_76;
wire n_403;
wire n_79;
wire n_282;
wire n_147;
wire n_359;
wire n_265;
wire n_231;
wire n_44;
wire n_482;
wire n_208;
wire n_162;
wire n_449;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_145;
wire n_266;
wire n_377;
wire n_109;
wire n_391;
wire n_427;
wire n_401;
wire n_148;
wire n_373;
wire n_396;
wire n_501;
wire n_392;
wire n_196;
wire n_375;
wire n_298;
wire n_330;
wire n_333;
wire n_450;
wire n_492;
wire n_152;
wire n_270;
wire n_159;
wire n_429;
wire n_347;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_336;
wire n_258;
wire n_458;
wire n_150;
wire n_41;
wire n_74;
wire n_475;
wire n_404;
wire n_158;
wire n_204;
wire n_241;
wire n_111;
wire n_479;
wire n_226;
wire n_125;
wire n_297;
wire n_413;
wire n_494;
wire n_75;
wire n_346;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_457;
wire n_119;
wire n_283;
wire n_181;
wire n_358;
wire n_256;
wire n_253;
wire n_273;
wire n_54;
wire n_168;
wire n_38;
wire n_442;
wire n_385;
wire n_201;
wire n_484;
wire n_260;
wire n_247;
wire n_249;
wire n_349;
wire n_418;
wire n_472;
wire n_292;
wire n_343;
wire n_486;
wire n_64;
wire n_291;
wire n_236;
wire n_370;
wire n_276;
wire n_374;
wire n_287;
wire n_388;
wire n_174;
wire n_400;
wire n_255;
wire n_243;
wire n_299;
wire n_352;
wire n_477;
wire n_56;
wire n_293;
wire n_275;
wire n_381;
wire n_227;
wire n_229;
wire n_454;
wire n_379;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_444;
wire n_360;
wire n_398;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_451;
wire n_45;
wire n_437;
wire n_313;
wire n_42;
wire n_268;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_416;
wire n_143;
wire n_351;
wire n_467;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_406;
wire n_303;
wire n_321;
wire n_100;
wire n_368;
wire n_51;
wire n_205;
wire n_361;
wire n_261;
wire n_86;
wire n_324;
wire n_70;
wire n_435;
wire n_32;
wire n_228;
wire n_389;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_438;
wire n_82;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_481;
wire n_191;
wire n_394;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_436;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_424;
wire n_133;
wire n_468;
wire n_257;
wire n_447;
wire n_344;
wire n_210;
wire n_206;
wire n_408;
wire n_85;
wire n_96;
wire n_308;
wire n_433;
wire n_364;

NAND2xp5_ASAP7_75t_L g41 ( 
.A(n_0),
.B(n_42),
.Y(n_41)
);

NAND2xp5_ASAP7_75t_L g72 ( 
.A(n_0),
.B(n_73),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_L g83 ( 
.A(n_0),
.B(n_84),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g122 ( 
.A(n_0),
.B(n_123),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_L g128 ( 
.A(n_0),
.B(n_129),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_L g180 ( 
.A(n_0),
.B(n_181),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_L g222 ( 
.A(n_0),
.B(n_223),
.Y(n_222)
);

INVx2_ASAP7_75t_L g285 ( 
.A(n_0),
.Y(n_285)
);

INVx8_ASAP7_75t_L g47 ( 
.A(n_1),
.Y(n_47)
);

CKINVDCx20_ASAP7_75t_R g501 ( 
.A(n_2),
.Y(n_501)
);

AND2x2_ASAP7_75t_L g184 ( 
.A(n_3),
.B(n_185),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_L g260 ( 
.A(n_3),
.B(n_261),
.Y(n_260)
);

NAND2xp5_ASAP7_75t_L g291 ( 
.A(n_3),
.B(n_292),
.Y(n_291)
);

NAND2xp5_ASAP7_75t_SL g308 ( 
.A(n_3),
.B(n_309),
.Y(n_308)
);

INVx1_ASAP7_75t_L g373 ( 
.A(n_3),
.Y(n_373)
);

NAND2xp5_ASAP7_75t_L g399 ( 
.A(n_3),
.B(n_290),
.Y(n_399)
);

NAND2xp5_ASAP7_75t_L g432 ( 
.A(n_3),
.B(n_433),
.Y(n_432)
);

AND2x2_ASAP7_75t_L g235 ( 
.A(n_4),
.B(n_236),
.Y(n_235)
);

AOI21xp5_ASAP7_75t_L g281 ( 
.A1(n_4),
.A2(n_282),
.B(n_284),
.Y(n_281)
);

INVx1_ASAP7_75t_L g344 ( 
.A(n_4),
.Y(n_344)
);

NAND2xp5_ASAP7_75t_L g353 ( 
.A(n_4),
.B(n_354),
.Y(n_353)
);

NAND2xp5_ASAP7_75t_L g376 ( 
.A(n_4),
.B(n_377),
.Y(n_376)
);

NAND2xp5_ASAP7_75t_L g393 ( 
.A(n_4),
.B(n_394),
.Y(n_393)
);

NAND2xp5_ASAP7_75t_L g429 ( 
.A(n_4),
.B(n_430),
.Y(n_429)
);

NAND2xp5_ASAP7_75t_L g441 ( 
.A(n_4),
.B(n_442),
.Y(n_441)
);

INVx2_ASAP7_75t_L g118 ( 
.A(n_5),
.Y(n_118)
);

BUFx3_ASAP7_75t_L g196 ( 
.A(n_5),
.Y(n_196)
);

BUFx6f_ASAP7_75t_L g268 ( 
.A(n_5),
.Y(n_268)
);

AND2x2_ASAP7_75t_L g152 ( 
.A(n_6),
.B(n_153),
.Y(n_152)
);

AND2x2_ASAP7_75t_L g219 ( 
.A(n_6),
.B(n_220),
.Y(n_219)
);

NAND2xp5_ASAP7_75t_L g242 ( 
.A(n_6),
.B(n_243),
.Y(n_242)
);

NAND2xp5_ASAP7_75t_L g271 ( 
.A(n_6),
.B(n_272),
.Y(n_271)
);

NAND2xp5_ASAP7_75t_L g304 ( 
.A(n_6),
.B(n_305),
.Y(n_304)
);

INVx1_ASAP7_75t_L g409 ( 
.A(n_6),
.Y(n_409)
);

NAND2xp5_ASAP7_75t_L g414 ( 
.A(n_6),
.B(n_415),
.Y(n_414)
);

NAND2xp5_ASAP7_75t_L g455 ( 
.A(n_6),
.B(n_456),
.Y(n_455)
);

CKINVDCx20_ASAP7_75t_R g276 ( 
.A(n_7),
.Y(n_276)
);

NAND2xp5_ASAP7_75t_L g313 ( 
.A(n_7),
.B(n_314),
.Y(n_313)
);

NAND2xp5_ASAP7_75t_L g369 ( 
.A(n_7),
.B(n_370),
.Y(n_369)
);

NAND2xp5_ASAP7_75t_L g400 ( 
.A(n_7),
.B(n_401),
.Y(n_400)
);

NAND2xp5_ASAP7_75t_L g424 ( 
.A(n_7),
.B(n_305),
.Y(n_424)
);

NAND2xp5_ASAP7_75t_L g435 ( 
.A(n_7),
.B(n_290),
.Y(n_435)
);

NAND2xp5_ASAP7_75t_L g437 ( 
.A(n_7),
.B(n_438),
.Y(n_437)
);

INVx6_ASAP7_75t_L g31 ( 
.A(n_8),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g147 ( 
.A(n_9),
.Y(n_147)
);

INVx8_ASAP7_75t_L g234 ( 
.A(n_9),
.Y(n_234)
);

INVx2_ASAP7_75t_L g288 ( 
.A(n_9),
.Y(n_288)
);

BUFx5_ASAP7_75t_L g442 ( 
.A(n_9),
.Y(n_442)
);

BUFx5_ASAP7_75t_L g39 ( 
.A(n_10),
.Y(n_39)
);

BUFx5_ASAP7_75t_L g58 ( 
.A(n_10),
.Y(n_58)
);

INVx3_ASAP7_75t_L g76 ( 
.A(n_10),
.Y(n_76)
);

BUFx6f_ASAP7_75t_L g283 ( 
.A(n_10),
.Y(n_283)
);

AND2x2_ASAP7_75t_SL g38 ( 
.A(n_11),
.B(n_39),
.Y(n_38)
);

NAND2xp5_ASAP7_75t_L g49 ( 
.A(n_11),
.B(n_50),
.Y(n_49)
);

AND2x2_ASAP7_75t_L g60 ( 
.A(n_11),
.B(n_61),
.Y(n_60)
);

AND2x2_ASAP7_75t_L g88 ( 
.A(n_11),
.B(n_89),
.Y(n_88)
);

AND2x2_ASAP7_75t_SL g134 ( 
.A(n_11),
.B(n_135),
.Y(n_134)
);

INVxp67_ASAP7_75t_L g149 ( 
.A(n_11),
.Y(n_149)
);

AND2x2_ASAP7_75t_L g194 ( 
.A(n_11),
.B(n_195),
.Y(n_194)
);

AND2x2_ASAP7_75t_L g230 ( 
.A(n_11),
.B(n_231),
.Y(n_230)
);

INVx8_ASAP7_75t_L g36 ( 
.A(n_12),
.Y(n_36)
);

INVx2_ASAP7_75t_L g43 ( 
.A(n_13),
.Y(n_43)
);

INVx6_ASAP7_75t_L g79 ( 
.A(n_13),
.Y(n_79)
);

BUFx6f_ASAP7_75t_L g114 ( 
.A(n_13),
.Y(n_114)
);

BUFx6f_ASAP7_75t_L g153 ( 
.A(n_13),
.Y(n_153)
);

BUFx5_ASAP7_75t_L g185 ( 
.A(n_13),
.Y(n_185)
);

BUFx6f_ASAP7_75t_L g236 ( 
.A(n_13),
.Y(n_236)
);

BUFx6f_ASAP7_75t_L g278 ( 
.A(n_13),
.Y(n_278)
);

NAND2xp5_ASAP7_75t_L g77 ( 
.A(n_14),
.B(n_78),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_L g91 ( 
.A(n_14),
.B(n_92),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_L g154 ( 
.A(n_14),
.B(n_155),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_L g197 ( 
.A(n_14),
.B(n_198),
.Y(n_197)
);

AND2x2_ASAP7_75t_L g237 ( 
.A(n_14),
.B(n_238),
.Y(n_237)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_14),
.Y(n_265)
);

NAND2xp5_ASAP7_75t_L g289 ( 
.A(n_14),
.B(n_290),
.Y(n_289)
);

NAND2xp5_ASAP7_75t_L g350 ( 
.A(n_14),
.B(n_351),
.Y(n_350)
);

INVx3_ASAP7_75t_L g498 ( 
.A(n_15),
.Y(n_498)
);

INVx1_ASAP7_75t_SL g29 ( 
.A(n_16),
.Y(n_29)
);

NAND2xp5_ASAP7_75t_SL g33 ( 
.A(n_16),
.B(n_34),
.Y(n_33)
);

AND2x2_ASAP7_75t_L g57 ( 
.A(n_16),
.B(n_58),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_L g68 ( 
.A(n_16),
.B(n_69),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_L g113 ( 
.A(n_16),
.B(n_114),
.Y(n_113)
);

AND2x2_ASAP7_75t_SL g115 ( 
.A(n_16),
.B(n_116),
.Y(n_115)
);

AND2x2_ASAP7_75t_SL g146 ( 
.A(n_16),
.B(n_147),
.Y(n_146)
);

BUFx3_ASAP7_75t_L g70 ( 
.A(n_17),
.Y(n_70)
);

BUFx5_ASAP7_75t_L g151 ( 
.A(n_17),
.Y(n_151)
);

INVx2_ASAP7_75t_L g183 ( 
.A(n_17),
.Y(n_183)
);

BUFx6f_ASAP7_75t_L g290 ( 
.A(n_17),
.Y(n_290)
);

AOI21xp5_ASAP7_75t_L g18 ( 
.A1(n_19),
.A2(n_497),
.B(n_499),
.Y(n_18)
);

XNOR2xp5_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_103),
.Y(n_19)
);

OAI21xp33_ASAP7_75t_L g20 ( 
.A1(n_21),
.A2(n_63),
.B(n_102),
.Y(n_20)
);

NAND2xp5_ASAP7_75t_SL g102 ( 
.A(n_21),
.B(n_63),
.Y(n_102)
);

BUFx24_ASAP7_75t_SL g503 ( 
.A(n_21),
.Y(n_503)
);

FAx1_ASAP7_75t_SL g21 ( 
.A(n_22),
.B(n_53),
.CI(n_54),
.CON(n_21),
.SN(n_21)
);

MAJIxp5_ASAP7_75t_L g22 ( 
.A(n_23),
.B(n_40),
.C(n_44),
.Y(n_22)
);

AOI22xp5_ASAP7_75t_L g98 ( 
.A1(n_23),
.A2(n_24),
.B1(n_99),
.B2(n_100),
.Y(n_98)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_24),
.Y(n_23)
);

OAI22xp5_ASAP7_75t_SL g24 ( 
.A1(n_25),
.A2(n_26),
.B1(n_37),
.B2(n_38),
.Y(n_24)
);

CKINVDCx16_ASAP7_75t_R g25 ( 
.A(n_26),
.Y(n_25)
);

AOI22xp5_ASAP7_75t_L g26 ( 
.A1(n_27),
.A2(n_28),
.B1(n_32),
.B2(n_33),
.Y(n_26)
);

MAJIxp5_ASAP7_75t_L g44 ( 
.A(n_27),
.B(n_45),
.C(n_48),
.Y(n_44)
);

AOI22xp5_ASAP7_75t_L g95 ( 
.A1(n_27),
.A2(n_28),
.B1(n_45),
.B2(n_96),
.Y(n_95)
);

AOI22xp5_ASAP7_75t_L g316 ( 
.A1(n_27),
.A2(n_28),
.B1(n_317),
.B2(n_318),
.Y(n_316)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_28),
.Y(n_27)
);

MAJIxp5_ASAP7_75t_L g53 ( 
.A(n_28),
.B(n_32),
.C(n_38),
.Y(n_53)
);

MAJIxp5_ASAP7_75t_L g228 ( 
.A(n_28),
.B(n_229),
.C(n_235),
.Y(n_228)
);

OR2x2_ASAP7_75t_L g28 ( 
.A(n_29),
.B(n_30),
.Y(n_28)
);

OR2x2_ASAP7_75t_L g45 ( 
.A(n_29),
.B(n_46),
.Y(n_45)
);

BUFx3_ASAP7_75t_L g30 ( 
.A(n_31),
.Y(n_30)
);

INVx3_ASAP7_75t_L g90 ( 
.A(n_31),
.Y(n_90)
);

INVx3_ASAP7_75t_L g133 ( 
.A(n_31),
.Y(n_133)
);

INVx3_ASAP7_75t_L g309 ( 
.A(n_31),
.Y(n_309)
);

AOI22xp5_ASAP7_75t_L g56 ( 
.A1(n_32),
.A2(n_33),
.B1(n_57),
.B2(n_59),
.Y(n_56)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_33),
.Y(n_32)
);

MAJIxp5_ASAP7_75t_L g179 ( 
.A(n_33),
.B(n_180),
.C(n_184),
.Y(n_179)
);

XNOR2xp5_ASAP7_75t_L g225 ( 
.A(n_33),
.B(n_226),
.Y(n_225)
);

INVx4_ASAP7_75t_L g34 ( 
.A(n_35),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_36),
.Y(n_35)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_36),
.Y(n_52)
);

INVx2_ASAP7_75t_L g86 ( 
.A(n_36),
.Y(n_86)
);

INVx6_ASAP7_75t_L g157 ( 
.A(n_36),
.Y(n_157)
);

BUFx5_ASAP7_75t_L g221 ( 
.A(n_36),
.Y(n_221)
);

BUFx6f_ASAP7_75t_L g371 ( 
.A(n_36),
.Y(n_371)
);

OAI22xp5_ASAP7_75t_SL g125 ( 
.A1(n_37),
.A2(n_38),
.B1(n_126),
.B2(n_127),
.Y(n_125)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_38),
.Y(n_37)
);

MAJIxp5_ASAP7_75t_L g163 ( 
.A(n_38),
.B(n_134),
.C(n_137),
.Y(n_163)
);

INVx1_ASAP7_75t_L g345 ( 
.A(n_39),
.Y(n_345)
);

OAI22xp5_ASAP7_75t_SL g100 ( 
.A1(n_40),
.A2(n_41),
.B1(n_44),
.B2(n_101),
.Y(n_100)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_41),
.Y(n_40)
);

INVx3_ASAP7_75t_L g42 ( 
.A(n_43),
.Y(n_42)
);

INVx3_ASAP7_75t_L g61 ( 
.A(n_43),
.Y(n_61)
);

CKINVDCx16_ASAP7_75t_R g101 ( 
.A(n_44),
.Y(n_101)
);

MAJIxp5_ASAP7_75t_L g66 ( 
.A(n_45),
.B(n_60),
.C(n_67),
.Y(n_66)
);

CKINVDCx20_ASAP7_75t_R g96 ( 
.A(n_45),
.Y(n_96)
);

AOI22xp5_ASAP7_75t_L g160 ( 
.A1(n_45),
.A2(n_96),
.B1(n_161),
.B2(n_162),
.Y(n_160)
);

AOI22xp5_ASAP7_75t_L g302 ( 
.A1(n_45),
.A2(n_96),
.B1(n_259),
.B2(n_260),
.Y(n_302)
);

BUFx3_ASAP7_75t_L g46 ( 
.A(n_47),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g124 ( 
.A(n_47),
.Y(n_124)
);

INVx3_ASAP7_75t_L g136 ( 
.A(n_47),
.Y(n_136)
);

INVx11_ASAP7_75t_L g240 ( 
.A(n_47),
.Y(n_240)
);

INVx2_ASAP7_75t_L g307 ( 
.A(n_47),
.Y(n_307)
);

BUFx3_ASAP7_75t_L g397 ( 
.A(n_47),
.Y(n_397)
);

OAI22xp5_ASAP7_75t_SL g93 ( 
.A1(n_48),
.A2(n_49),
.B1(n_94),
.B2(n_95),
.Y(n_93)
);

AOI22xp5_ASAP7_75t_L g177 ( 
.A1(n_48),
.A2(n_49),
.B1(n_122),
.B2(n_178),
.Y(n_177)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_49),
.Y(n_48)
);

MAJIxp5_ASAP7_75t_L g121 ( 
.A(n_49),
.B(n_120),
.C(n_122),
.Y(n_121)
);

INVx4_ASAP7_75t_L g50 ( 
.A(n_51),
.Y(n_50)
);

INVx3_ASAP7_75t_L g51 ( 
.A(n_52),
.Y(n_51)
);

OAI22xp5_ASAP7_75t_SL g54 ( 
.A1(n_55),
.A2(n_56),
.B1(n_60),
.B2(n_62),
.Y(n_54)
);

CKINVDCx20_ASAP7_75t_R g55 ( 
.A(n_56),
.Y(n_55)
);

CKINVDCx16_ASAP7_75t_R g59 ( 
.A(n_57),
.Y(n_59)
);

MAJx2_ASAP7_75t_L g192 ( 
.A(n_57),
.B(n_193),
.C(n_197),
.Y(n_192)
);

AOI22xp5_ASAP7_75t_L g202 ( 
.A1(n_57),
.A2(n_59),
.B1(n_154),
.B2(n_203),
.Y(n_202)
);

OAI22xp5_ASAP7_75t_SL g246 ( 
.A1(n_57),
.A2(n_59),
.B1(n_197),
.B2(n_247),
.Y(n_246)
);

MAJIxp5_ASAP7_75t_L g143 ( 
.A(n_59),
.B(n_144),
.C(n_154),
.Y(n_143)
);

CKINVDCx20_ASAP7_75t_R g62 ( 
.A(n_60),
.Y(n_62)
);

OAI22xp5_ASAP7_75t_SL g162 ( 
.A1(n_60),
.A2(n_62),
.B1(n_67),
.B2(n_68),
.Y(n_162)
);

MAJIxp5_ASAP7_75t_L g63 ( 
.A(n_64),
.B(n_97),
.C(n_98),
.Y(n_63)
);

XNOR2xp5_ASAP7_75t_L g494 ( 
.A(n_64),
.B(n_495),
.Y(n_494)
);

MAJIxp5_ASAP7_75t_L g64 ( 
.A(n_65),
.B(n_82),
.C(n_93),
.Y(n_64)
);

XNOR2xp5_ASAP7_75t_L g165 ( 
.A(n_65),
.B(n_166),
.Y(n_165)
);

XOR2xp5_ASAP7_75t_L g65 ( 
.A(n_66),
.B(n_71),
.Y(n_65)
);

MAJIxp5_ASAP7_75t_L g97 ( 
.A(n_66),
.B(n_77),
.C(n_80),
.Y(n_97)
);

OAI22xp5_ASAP7_75t_SL g110 ( 
.A1(n_67),
.A2(n_68),
.B1(n_111),
.B2(n_112),
.Y(n_110)
);

MAJIxp5_ASAP7_75t_L g164 ( 
.A(n_67),
.B(n_113),
.C(n_120),
.Y(n_164)
);

AOI22xp5_ASAP7_75t_L g365 ( 
.A1(n_67),
.A2(n_68),
.B1(n_308),
.B2(n_366),
.Y(n_365)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_68),
.Y(n_67)
);

MAJIxp5_ASAP7_75t_L g303 ( 
.A(n_68),
.B(n_304),
.C(n_308),
.Y(n_303)
);

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_70),
.Y(n_69)
);

OAI22xp5_ASAP7_75t_SL g71 ( 
.A1(n_72),
.A2(n_77),
.B1(n_80),
.B2(n_81),
.Y(n_71)
);

CKINVDCx20_ASAP7_75t_R g80 ( 
.A(n_72),
.Y(n_80)
);

INVx3_ASAP7_75t_L g73 ( 
.A(n_74),
.Y(n_73)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_74),
.Y(n_92)
);

INVx6_ASAP7_75t_L g74 ( 
.A(n_75),
.Y(n_74)
);

INVx5_ASAP7_75t_L g75 ( 
.A(n_76),
.Y(n_75)
);

BUFx6f_ASAP7_75t_L g244 ( 
.A(n_76),
.Y(n_244)
);

INVx3_ASAP7_75t_L g292 ( 
.A(n_76),
.Y(n_292)
);

CKINVDCx20_ASAP7_75t_R g81 ( 
.A(n_77),
.Y(n_81)
);

INVx8_ASAP7_75t_L g78 ( 
.A(n_79),
.Y(n_78)
);

XNOR2xp5_ASAP7_75t_L g166 ( 
.A(n_82),
.B(n_93),
.Y(n_166)
);

MAJIxp5_ASAP7_75t_L g82 ( 
.A(n_83),
.B(n_87),
.C(n_91),
.Y(n_82)
);

AOI22xp5_ASAP7_75t_L g140 ( 
.A1(n_83),
.A2(n_87),
.B1(n_88),
.B2(n_141),
.Y(n_140)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_83),
.Y(n_141)
);

INVx2_ASAP7_75t_L g84 ( 
.A(n_85),
.Y(n_84)
);

INVx6_ASAP7_75t_L g85 ( 
.A(n_86),
.Y(n_85)
);

OAI22xp5_ASAP7_75t_L g213 ( 
.A1(n_87),
.A2(n_88),
.B1(n_214),
.B2(n_215),
.Y(n_213)
);

CKINVDCx20_ASAP7_75t_R g87 ( 
.A(n_88),
.Y(n_87)
);

MAJIxp5_ASAP7_75t_L g193 ( 
.A(n_88),
.B(n_146),
.C(n_194),
.Y(n_193)
);

BUFx6f_ASAP7_75t_L g89 ( 
.A(n_90),
.Y(n_89)
);

INVx4_ASAP7_75t_L g200 ( 
.A(n_90),
.Y(n_200)
);

XNOR2xp5_ASAP7_75t_L g139 ( 
.A(n_91),
.B(n_140),
.Y(n_139)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_95),
.Y(n_94)
);

MAJIxp5_ASAP7_75t_L g258 ( 
.A(n_96),
.B(n_259),
.C(n_264),
.Y(n_258)
);

XNOR2xp5_ASAP7_75t_L g495 ( 
.A(n_97),
.B(n_98),
.Y(n_495)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_100),
.Y(n_99)
);

AO21x1_ASAP7_75t_SL g103 ( 
.A1(n_104),
.A2(n_492),
.B(n_496),
.Y(n_103)
);

OAI21xp33_ASAP7_75t_L g104 ( 
.A1(n_105),
.A2(n_249),
.B(n_489),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_L g105 ( 
.A(n_106),
.B(n_205),
.Y(n_105)
);

AOI21xp33_ASAP7_75t_SL g489 ( 
.A1(n_106),
.A2(n_490),
.B(n_491),
.Y(n_489)
);

NAND2xp5_ASAP7_75t_SL g106 ( 
.A(n_107),
.B(n_167),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g491 ( 
.A(n_107),
.B(n_167),
.Y(n_491)
);

XOR2xp5_ASAP7_75t_L g107 ( 
.A(n_108),
.B(n_158),
.Y(n_107)
);

MAJIxp5_ASAP7_75t_L g493 ( 
.A(n_108),
.B(n_159),
.C(n_165),
.Y(n_493)
);

MAJIxp5_ASAP7_75t_L g108 ( 
.A(n_109),
.B(n_139),
.C(n_142),
.Y(n_108)
);

XNOR2xp5_ASAP7_75t_SL g168 ( 
.A(n_109),
.B(n_169),
.Y(n_168)
);

MAJIxp5_ASAP7_75t_L g109 ( 
.A(n_110),
.B(n_121),
.C(n_125),
.Y(n_109)
);

XNOR2xp5_ASAP7_75t_L g209 ( 
.A(n_110),
.B(n_210),
.Y(n_209)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_112),
.Y(n_111)
);

AOI22xp5_ASAP7_75t_L g112 ( 
.A1(n_113),
.A2(n_115),
.B1(n_119),
.B2(n_120),
.Y(n_112)
);

CKINVDCx14_ASAP7_75t_R g119 ( 
.A(n_113),
.Y(n_119)
);

INVx1_ASAP7_75t_SL g120 ( 
.A(n_115),
.Y(n_120)
);

OAI22xp5_ASAP7_75t_L g175 ( 
.A1(n_115),
.A2(n_120),
.B1(n_176),
.B2(n_177),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_SL g348 ( 
.A(n_115),
.B(n_230),
.Y(n_348)
);

AOI22xp5_ASAP7_75t_L g457 ( 
.A1(n_115),
.A2(n_120),
.B1(n_229),
.B2(n_230),
.Y(n_457)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_116),
.Y(n_224)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_117),
.Y(n_116)
);

BUFx3_ASAP7_75t_L g117 ( 
.A(n_118),
.Y(n_117)
);

XNOR2xp5_ASAP7_75t_L g210 ( 
.A(n_121),
.B(n_125),
.Y(n_210)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_122),
.Y(n_178)
);

INVx5_ASAP7_75t_L g123 ( 
.A(n_124),
.Y(n_123)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_127),
.Y(n_126)
);

AOI22xp5_ASAP7_75t_L g127 ( 
.A1(n_128),
.A2(n_134),
.B1(n_137),
.B2(n_138),
.Y(n_127)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_128),
.Y(n_137)
);

INVx2_ASAP7_75t_L g129 ( 
.A(n_130),
.Y(n_129)
);

INVx4_ASAP7_75t_L g130 ( 
.A(n_131),
.Y(n_130)
);

INVx8_ASAP7_75t_L g131 ( 
.A(n_132),
.Y(n_131)
);

INVx6_ASAP7_75t_L g274 ( 
.A(n_132),
.Y(n_274)
);

INVx4_ASAP7_75t_L g132 ( 
.A(n_133),
.Y(n_132)
);

BUFx6f_ASAP7_75t_L g402 ( 
.A(n_133),
.Y(n_402)
);

INVx1_ASAP7_75t_SL g138 ( 
.A(n_134),
.Y(n_138)
);

XNOR2xp5_ASAP7_75t_L g257 ( 
.A(n_134),
.B(n_219),
.Y(n_257)
);

BUFx6f_ASAP7_75t_L g135 ( 
.A(n_136),
.Y(n_135)
);

MAJIxp5_ASAP7_75t_L g217 ( 
.A(n_138),
.B(n_218),
.C(n_222),
.Y(n_217)
);

OAI22xp5_ASAP7_75t_SL g169 ( 
.A1(n_139),
.A2(n_142),
.B1(n_143),
.B2(n_170),
.Y(n_169)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_139),
.Y(n_170)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_143),
.Y(n_142)
);

OA22x2_ASAP7_75t_L g201 ( 
.A1(n_144),
.A2(n_145),
.B1(n_202),
.B2(n_204),
.Y(n_201)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_145),
.Y(n_144)
);

MAJIxp5_ASAP7_75t_L g145 ( 
.A(n_146),
.B(n_148),
.C(n_152),
.Y(n_145)
);

OAI22xp5_ASAP7_75t_L g187 ( 
.A1(n_146),
.A2(n_152),
.B1(n_188),
.B2(n_189),
.Y(n_187)
);

CKINVDCx20_ASAP7_75t_R g188 ( 
.A(n_146),
.Y(n_188)
);

AOI22xp5_ASAP7_75t_L g215 ( 
.A1(n_146),
.A2(n_188),
.B1(n_194),
.B2(n_216),
.Y(n_215)
);

AOI22xp5_ASAP7_75t_L g413 ( 
.A1(n_146),
.A2(n_188),
.B1(n_414),
.B2(n_416),
.Y(n_413)
);

NAND2xp5_ASAP7_75t_SL g458 ( 
.A(n_146),
.B(n_416),
.Y(n_458)
);

INVx4_ASAP7_75t_L g434 ( 
.A(n_147),
.Y(n_434)
);

OAI22xp5_ASAP7_75t_L g186 ( 
.A1(n_148),
.A2(n_187),
.B1(n_190),
.B2(n_191),
.Y(n_186)
);

CKINVDCx20_ASAP7_75t_R g190 ( 
.A(n_148),
.Y(n_190)
);

MAJIxp5_ASAP7_75t_L g270 ( 
.A(n_148),
.B(n_271),
.C(n_275),
.Y(n_270)
);

OAI22xp5_ASAP7_75t_SL g340 ( 
.A1(n_148),
.A2(n_190),
.B1(n_271),
.B2(n_341),
.Y(n_340)
);

OR2x2_ASAP7_75t_L g148 ( 
.A(n_149),
.B(n_150),
.Y(n_148)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_151),
.Y(n_150)
);

CKINVDCx20_ASAP7_75t_R g189 ( 
.A(n_152),
.Y(n_189)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_154),
.Y(n_203)
);

BUFx12f_ASAP7_75t_L g155 ( 
.A(n_156),
.Y(n_155)
);

BUFx6f_ASAP7_75t_L g156 ( 
.A(n_157),
.Y(n_156)
);

BUFx6f_ASAP7_75t_L g263 ( 
.A(n_157),
.Y(n_263)
);

XNOR2xp5_ASAP7_75t_L g158 ( 
.A(n_159),
.B(n_165),
.Y(n_158)
);

MAJIxp5_ASAP7_75t_L g159 ( 
.A(n_160),
.B(n_163),
.C(n_164),
.Y(n_159)
);

XOR2xp5_ASAP7_75t_L g171 ( 
.A(n_160),
.B(n_172),
.Y(n_171)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_162),
.Y(n_161)
);

XNOR2xp5_ASAP7_75t_L g172 ( 
.A(n_163),
.B(n_164),
.Y(n_172)
);

MAJIxp5_ASAP7_75t_L g167 ( 
.A(n_168),
.B(n_171),
.C(n_173),
.Y(n_167)
);

FAx1_ASAP7_75t_SL g248 ( 
.A(n_168),
.B(n_171),
.CI(n_173),
.CON(n_248),
.SN(n_248)
);

MAJIxp5_ASAP7_75t_L g173 ( 
.A(n_174),
.B(n_192),
.C(n_201),
.Y(n_173)
);

XOR2xp5_ASAP7_75t_L g207 ( 
.A(n_174),
.B(n_208),
.Y(n_207)
);

MAJIxp5_ASAP7_75t_L g174 ( 
.A(n_175),
.B(n_179),
.C(n_186),
.Y(n_174)
);

XNOR2xp5_ASAP7_75t_L g325 ( 
.A(n_175),
.B(n_179),
.Y(n_325)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_177),
.Y(n_176)
);

XOR2xp5_ASAP7_75t_L g226 ( 
.A(n_180),
.B(n_184),
.Y(n_226)
);

INVx2_ASAP7_75t_L g181 ( 
.A(n_182),
.Y(n_181)
);

BUFx3_ASAP7_75t_L g182 ( 
.A(n_183),
.Y(n_182)
);

BUFx6f_ASAP7_75t_L g422 ( 
.A(n_183),
.Y(n_422)
);

XOR2xp5_ASAP7_75t_L g324 ( 
.A(n_186),
.B(n_325),
.Y(n_324)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_187),
.Y(n_191)
);

XNOR2xp5_ASAP7_75t_L g208 ( 
.A(n_192),
.B(n_201),
.Y(n_208)
);

XOR2xp5_ASAP7_75t_L g245 ( 
.A(n_193),
.B(n_246),
.Y(n_245)
);

CKINVDCx16_ASAP7_75t_R g216 ( 
.A(n_194),
.Y(n_216)
);

NAND2xp5_ASAP7_75t_L g311 ( 
.A(n_194),
.B(n_312),
.Y(n_311)
);

OAI22xp5_ASAP7_75t_SL g380 ( 
.A1(n_194),
.A2(n_216),
.B1(n_312),
.B2(n_313),
.Y(n_380)
);

BUFx2_ASAP7_75t_L g407 ( 
.A(n_195),
.Y(n_407)
);

INVx8_ASAP7_75t_L g431 ( 
.A(n_195),
.Y(n_431)
);

BUFx8_ASAP7_75t_L g195 ( 
.A(n_196),
.Y(n_195)
);

BUFx5_ASAP7_75t_L g440 ( 
.A(n_196),
.Y(n_440)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_197),
.Y(n_247)
);

INVx3_ASAP7_75t_L g198 ( 
.A(n_199),
.Y(n_198)
);

BUFx6f_ASAP7_75t_L g199 ( 
.A(n_200),
.Y(n_199)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_202),
.Y(n_204)
);

NAND2xp5_ASAP7_75t_L g205 ( 
.A(n_206),
.B(n_248),
.Y(n_205)
);

NOR2xp33_ASAP7_75t_L g490 ( 
.A(n_206),
.B(n_248),
.Y(n_490)
);

MAJIxp5_ASAP7_75t_L g206 ( 
.A(n_207),
.B(n_209),
.C(n_211),
.Y(n_206)
);

XNOR2xp5_ASAP7_75t_L g332 ( 
.A(n_207),
.B(n_209),
.Y(n_332)
);

XNOR2xp5_ASAP7_75t_L g331 ( 
.A(n_211),
.B(n_332),
.Y(n_331)
);

MAJIxp5_ASAP7_75t_L g211 ( 
.A(n_212),
.B(n_227),
.C(n_245),
.Y(n_211)
);

XNOR2xp5_ASAP7_75t_SL g326 ( 
.A(n_212),
.B(n_327),
.Y(n_326)
);

MAJIxp5_ASAP7_75t_L g212 ( 
.A(n_213),
.B(n_217),
.C(n_225),
.Y(n_212)
);

HB1xp67_ASAP7_75t_L g297 ( 
.A(n_213),
.Y(n_297)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_215),
.Y(n_214)
);

XNOR2xp5_ASAP7_75t_L g298 ( 
.A(n_217),
.B(n_225),
.Y(n_298)
);

INVxp67_ASAP7_75t_L g218 ( 
.A(n_219),
.Y(n_218)
);

INVx5_ASAP7_75t_L g220 ( 
.A(n_221),
.Y(n_220)
);

XOR2xp5_ASAP7_75t_L g256 ( 
.A(n_222),
.B(n_257),
.Y(n_256)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_224),
.Y(n_223)
);

XNOR2xp5_ASAP7_75t_L g327 ( 
.A(n_227),
.B(n_245),
.Y(n_327)
);

MAJIxp5_ASAP7_75t_L g227 ( 
.A(n_228),
.B(n_237),
.C(n_241),
.Y(n_227)
);

XNOR2xp5_ASAP7_75t_L g293 ( 
.A(n_228),
.B(n_294),
.Y(n_293)
);

OAI22xp5_ASAP7_75t_SL g318 ( 
.A1(n_229),
.A2(n_230),
.B1(n_235),
.B2(n_319),
.Y(n_318)
);

INVx1_ASAP7_75t_SL g229 ( 
.A(n_230),
.Y(n_229)
);

INVx2_ASAP7_75t_L g231 ( 
.A(n_232),
.Y(n_231)
);

INVx3_ASAP7_75t_L g232 ( 
.A(n_233),
.Y(n_232)
);

INVx3_ASAP7_75t_L g233 ( 
.A(n_234),
.Y(n_233)
);

INVx4_ASAP7_75t_L g351 ( 
.A(n_234),
.Y(n_351)
);

BUFx6f_ASAP7_75t_L g412 ( 
.A(n_234),
.Y(n_412)
);

CKINVDCx20_ASAP7_75t_R g319 ( 
.A(n_235),
.Y(n_319)
);

AOI22xp5_ASAP7_75t_SL g294 ( 
.A1(n_237),
.A2(n_241),
.B1(n_242),
.B2(n_295),
.Y(n_294)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_237),
.Y(n_295)
);

INVx4_ASAP7_75t_L g238 ( 
.A(n_239),
.Y(n_238)
);

INVx5_ASAP7_75t_L g239 ( 
.A(n_240),
.Y(n_239)
);

INVx6_ASAP7_75t_L g374 ( 
.A(n_240),
.Y(n_374)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_242),
.Y(n_241)
);

INVx6_ASAP7_75t_L g243 ( 
.A(n_244),
.Y(n_243)
);

BUFx24_ASAP7_75t_SL g504 ( 
.A(n_248),
.Y(n_504)
);

AOI221xp5_ASAP7_75t_L g249 ( 
.A1(n_250),
.A2(n_386),
.B1(n_482),
.B2(n_487),
.C(n_488),
.Y(n_249)
);

NOR3xp33_ASAP7_75t_SL g250 ( 
.A(n_251),
.B(n_329),
.C(n_333),
.Y(n_250)
);

OAI21xp5_ASAP7_75t_SL g482 ( 
.A1(n_251),
.A2(n_483),
.B(n_486),
.Y(n_482)
);

AND2x2_ASAP7_75t_L g251 ( 
.A(n_252),
.B(n_322),
.Y(n_251)
);

OR2x2_ASAP7_75t_L g486 ( 
.A(n_252),
.B(n_322),
.Y(n_486)
);

MAJIxp5_ASAP7_75t_L g252 ( 
.A(n_253),
.B(n_296),
.C(n_299),
.Y(n_252)
);

XNOR2xp5_ASAP7_75t_L g358 ( 
.A(n_253),
.B(n_296),
.Y(n_358)
);

XNOR2xp5_ASAP7_75t_SL g253 ( 
.A(n_254),
.B(n_279),
.Y(n_253)
);

MAJIxp5_ASAP7_75t_L g328 ( 
.A(n_254),
.B(n_280),
.C(n_293),
.Y(n_328)
);

MAJIxp5_ASAP7_75t_L g254 ( 
.A(n_255),
.B(n_258),
.C(n_269),
.Y(n_254)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_256),
.Y(n_255)
);

XNOR2xp5_ASAP7_75t_L g356 ( 
.A(n_256),
.B(n_270),
.Y(n_356)
);

XOR2xp5_ASAP7_75t_L g355 ( 
.A(n_258),
.B(n_356),
.Y(n_355)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_260),
.Y(n_259)
);

INVx6_ASAP7_75t_L g261 ( 
.A(n_262),
.Y(n_261)
);

INVx5_ASAP7_75t_L g262 ( 
.A(n_263),
.Y(n_262)
);

BUFx6f_ASAP7_75t_L g354 ( 
.A(n_263),
.Y(n_354)
);

XNOR2xp5_ASAP7_75t_SL g301 ( 
.A(n_264),
.B(n_302),
.Y(n_301)
);

NOR2xp33_ASAP7_75t_L g264 ( 
.A(n_265),
.B(n_266),
.Y(n_264)
);

INVx5_ASAP7_75t_L g266 ( 
.A(n_267),
.Y(n_266)
);

BUFx6f_ASAP7_75t_L g267 ( 
.A(n_268),
.Y(n_267)
);

BUFx5_ASAP7_75t_L g415 ( 
.A(n_268),
.Y(n_415)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_270),
.Y(n_269)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_271),
.Y(n_341)
);

INVx2_ASAP7_75t_L g272 ( 
.A(n_273),
.Y(n_272)
);

INVx3_ASAP7_75t_L g273 ( 
.A(n_274),
.Y(n_273)
);

XOR2xp5_ASAP7_75t_L g339 ( 
.A(n_275),
.B(n_340),
.Y(n_339)
);

NOR2xp33_ASAP7_75t_L g275 ( 
.A(n_276),
.B(n_277),
.Y(n_275)
);

INVx2_ASAP7_75t_L g277 ( 
.A(n_278),
.Y(n_277)
);

XNOR2xp5_ASAP7_75t_L g279 ( 
.A(n_280),
.B(n_293),
.Y(n_279)
);

MAJIxp5_ASAP7_75t_L g280 ( 
.A(n_281),
.B(n_289),
.C(n_291),
.Y(n_280)
);

XNOR2xp5_ASAP7_75t_L g320 ( 
.A(n_281),
.B(n_321),
.Y(n_320)
);

AOI21xp5_ASAP7_75t_L g342 ( 
.A1(n_281),
.A2(n_284),
.B(n_343),
.Y(n_342)
);

BUFx6f_ASAP7_75t_L g282 ( 
.A(n_283),
.Y(n_282)
);

INVx4_ASAP7_75t_L g315 ( 
.A(n_283),
.Y(n_315)
);

NOR2xp33_ASAP7_75t_L g284 ( 
.A(n_285),
.B(n_286),
.Y(n_284)
);

INVx5_ASAP7_75t_L g286 ( 
.A(n_287),
.Y(n_286)
);

INVx2_ASAP7_75t_L g287 ( 
.A(n_288),
.Y(n_287)
);

XNOR2xp5_ASAP7_75t_L g321 ( 
.A(n_289),
.B(n_291),
.Y(n_321)
);

XNOR2xp5_ASAP7_75t_L g296 ( 
.A(n_297),
.B(n_298),
.Y(n_296)
);

XOR2xp5_ASAP7_75t_L g357 ( 
.A(n_299),
.B(n_358),
.Y(n_357)
);

MAJIxp5_ASAP7_75t_L g299 ( 
.A(n_300),
.B(n_316),
.C(n_320),
.Y(n_299)
);

XOR2xp5_ASAP7_75t_L g336 ( 
.A(n_300),
.B(n_337),
.Y(n_336)
);

MAJIxp5_ASAP7_75t_L g300 ( 
.A(n_301),
.B(n_303),
.C(n_310),
.Y(n_300)
);

XNOR2xp5_ASAP7_75t_L g381 ( 
.A(n_301),
.B(n_382),
.Y(n_381)
);

AOI22xp5_ASAP7_75t_L g382 ( 
.A1(n_303),
.A2(n_310),
.B1(n_311),
.B2(n_383),
.Y(n_382)
);

INVx1_ASAP7_75t_L g383 ( 
.A(n_303),
.Y(n_383)
);

XNOR2xp5_ASAP7_75t_SL g364 ( 
.A(n_304),
.B(n_365),
.Y(n_364)
);

INVx2_ASAP7_75t_L g305 ( 
.A(n_306),
.Y(n_305)
);

INVx4_ASAP7_75t_L g306 ( 
.A(n_307),
.Y(n_306)
);

INVxp67_ASAP7_75t_L g366 ( 
.A(n_308),
.Y(n_366)
);

INVx6_ASAP7_75t_L g378 ( 
.A(n_309),
.Y(n_378)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_311),
.Y(n_310)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_313),
.Y(n_312)
);

INVx6_ASAP7_75t_L g314 ( 
.A(n_315),
.Y(n_314)
);

XNOR2xp5_ASAP7_75t_L g337 ( 
.A(n_316),
.B(n_320),
.Y(n_337)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_318),
.Y(n_317)
);

XNOR2xp5_ASAP7_75t_L g322 ( 
.A(n_323),
.B(n_328),
.Y(n_322)
);

XNOR2xp5_ASAP7_75t_L g323 ( 
.A(n_324),
.B(n_326),
.Y(n_323)
);

MAJIxp5_ASAP7_75t_L g330 ( 
.A(n_324),
.B(n_326),
.C(n_328),
.Y(n_330)
);

INVx1_ASAP7_75t_L g487 ( 
.A(n_329),
.Y(n_487)
);

NOR2xp33_ASAP7_75t_L g329 ( 
.A(n_330),
.B(n_331),
.Y(n_329)
);

AND2x2_ASAP7_75t_L g488 ( 
.A(n_330),
.B(n_331),
.Y(n_488)
);

NAND2xp5_ASAP7_75t_SL g333 ( 
.A(n_334),
.B(n_359),
.Y(n_333)
);

AOI21xp5_ASAP7_75t_L g483 ( 
.A1(n_334),
.A2(n_484),
.B(n_485),
.Y(n_483)
);

NAND2xp5_ASAP7_75t_L g334 ( 
.A(n_335),
.B(n_357),
.Y(n_334)
);

NOR2xp33_ASAP7_75t_L g485 ( 
.A(n_335),
.B(n_357),
.Y(n_485)
);

MAJIxp5_ASAP7_75t_L g335 ( 
.A(n_336),
.B(n_338),
.C(n_355),
.Y(n_335)
);

XOR2xp5_ASAP7_75t_L g384 ( 
.A(n_336),
.B(n_385),
.Y(n_384)
);

XNOR2xp5_ASAP7_75t_L g385 ( 
.A(n_338),
.B(n_355),
.Y(n_385)
);

MAJIxp5_ASAP7_75t_L g338 ( 
.A(n_339),
.B(n_342),
.C(n_346),
.Y(n_338)
);

XNOR2xp5_ASAP7_75t_L g362 ( 
.A(n_339),
.B(n_342),
.Y(n_362)
);

NOR2xp33_ASAP7_75t_L g343 ( 
.A(n_344),
.B(n_345),
.Y(n_343)
);

NOR2xp33_ASAP7_75t_L g419 ( 
.A(n_344),
.B(n_420),
.Y(n_419)
);

XOR2xp5_ASAP7_75t_L g361 ( 
.A(n_346),
.B(n_362),
.Y(n_361)
);

MAJIxp5_ASAP7_75t_L g346 ( 
.A(n_347),
.B(n_349),
.C(n_352),
.Y(n_346)
);

AOI22xp5_ASAP7_75t_L g469 ( 
.A1(n_347),
.A2(n_348),
.B1(n_470),
.B2(n_471),
.Y(n_469)
);

INVx1_ASAP7_75t_L g347 ( 
.A(n_348),
.Y(n_347)
);

AOI22xp5_ASAP7_75t_L g470 ( 
.A1(n_349),
.A2(n_350),
.B1(n_352),
.B2(n_353),
.Y(n_470)
);

CKINVDCx14_ASAP7_75t_R g349 ( 
.A(n_350),
.Y(n_349)
);

INVx1_ASAP7_75t_L g352 ( 
.A(n_353),
.Y(n_352)
);

NAND2xp5_ASAP7_75t_L g359 ( 
.A(n_360),
.B(n_384),
.Y(n_359)
);

NOR2xp33_ASAP7_75t_L g484 ( 
.A(n_360),
.B(n_384),
.Y(n_484)
);

MAJIxp5_ASAP7_75t_L g360 ( 
.A(n_361),
.B(n_363),
.C(n_381),
.Y(n_360)
);

XNOR2xp5_ASAP7_75t_L g479 ( 
.A(n_361),
.B(n_480),
.Y(n_479)
);

XNOR2xp5_ASAP7_75t_L g480 ( 
.A(n_363),
.B(n_381),
.Y(n_480)
);

MAJIxp5_ASAP7_75t_L g363 ( 
.A(n_364),
.B(n_367),
.C(n_379),
.Y(n_363)
);

XNOR2xp5_ASAP7_75t_SL g472 ( 
.A(n_364),
.B(n_473),
.Y(n_472)
);

AOI22xp5_ASAP7_75t_L g473 ( 
.A1(n_367),
.A2(n_379),
.B1(n_380),
.B2(n_474),
.Y(n_473)
);

INVx1_ASAP7_75t_L g474 ( 
.A(n_367),
.Y(n_474)
);

MAJIxp5_ASAP7_75t_L g367 ( 
.A(n_368),
.B(n_372),
.C(n_375),
.Y(n_367)
);

AOI22xp5_ASAP7_75t_L g462 ( 
.A1(n_368),
.A2(n_369),
.B1(n_375),
.B2(n_376),
.Y(n_462)
);

INVx1_ASAP7_75t_L g368 ( 
.A(n_369),
.Y(n_368)
);

INVx1_ASAP7_75t_L g370 ( 
.A(n_371),
.Y(n_370)
);

XNOR2xp5_ASAP7_75t_L g461 ( 
.A(n_372),
.B(n_462),
.Y(n_461)
);

NOR2xp33_ASAP7_75t_L g372 ( 
.A(n_373),
.B(n_374),
.Y(n_372)
);

NOR2xp33_ASAP7_75t_L g405 ( 
.A(n_373),
.B(n_406),
.Y(n_405)
);

INVx1_ASAP7_75t_L g375 ( 
.A(n_376),
.Y(n_375)
);

INVx4_ASAP7_75t_L g377 ( 
.A(n_378),
.Y(n_377)
);

INVx1_ASAP7_75t_L g379 ( 
.A(n_380),
.Y(n_379)
);

OAI21xp5_ASAP7_75t_SL g386 ( 
.A1(n_387),
.A2(n_477),
.B(n_481),
.Y(n_386)
);

AOI21xp5_ASAP7_75t_L g387 ( 
.A1(n_388),
.A2(n_464),
.B(n_476),
.Y(n_387)
);

OAI21xp5_ASAP7_75t_L g388 ( 
.A1(n_389),
.A2(n_451),
.B(n_463),
.Y(n_388)
);

AOI21xp5_ASAP7_75t_L g389 ( 
.A1(n_390),
.A2(n_425),
.B(n_450),
.Y(n_389)
);

NAND2xp5_ASAP7_75t_SL g390 ( 
.A(n_391),
.B(n_417),
.Y(n_390)
);

NOR2xp33_ASAP7_75t_L g450 ( 
.A(n_391),
.B(n_417),
.Y(n_450)
);

XNOR2xp5_ASAP7_75t_L g391 ( 
.A(n_392),
.B(n_403),
.Y(n_391)
);

MAJIxp5_ASAP7_75t_L g452 ( 
.A(n_392),
.B(n_404),
.C(n_413),
.Y(n_452)
);

XOR2xp5_ASAP7_75t_L g392 ( 
.A(n_393),
.B(n_398),
.Y(n_392)
);

MAJIxp5_ASAP7_75t_L g460 ( 
.A(n_393),
.B(n_399),
.C(n_400),
.Y(n_460)
);

INVx1_ASAP7_75t_L g394 ( 
.A(n_395),
.Y(n_394)
);

INVx2_ASAP7_75t_L g395 ( 
.A(n_396),
.Y(n_395)
);

INVx3_ASAP7_75t_L g396 ( 
.A(n_397),
.Y(n_396)
);

XOR2xp5_ASAP7_75t_L g398 ( 
.A(n_399),
.B(n_400),
.Y(n_398)
);

BUFx2_ASAP7_75t_L g401 ( 
.A(n_402),
.Y(n_401)
);

XNOR2xp5_ASAP7_75t_L g403 ( 
.A(n_404),
.B(n_413),
.Y(n_403)
);

NAND2xp5_ASAP7_75t_L g404 ( 
.A(n_405),
.B(n_408),
.Y(n_404)
);

XOR2xp5_ASAP7_75t_L g418 ( 
.A(n_405),
.B(n_408),
.Y(n_418)
);

INVx2_ASAP7_75t_L g406 ( 
.A(n_407),
.Y(n_406)
);

NOR2xp33_ASAP7_75t_L g408 ( 
.A(n_409),
.B(n_410),
.Y(n_408)
);

INVx2_ASAP7_75t_L g410 ( 
.A(n_411),
.Y(n_410)
);

INVx8_ASAP7_75t_L g411 ( 
.A(n_412),
.Y(n_411)
);

INVx1_ASAP7_75t_L g416 ( 
.A(n_414),
.Y(n_416)
);

MAJIxp5_ASAP7_75t_L g417 ( 
.A(n_418),
.B(n_419),
.C(n_423),
.Y(n_417)
);

XOR2xp5_ASAP7_75t_L g446 ( 
.A(n_418),
.B(n_447),
.Y(n_446)
);

OAI22xp5_ASAP7_75t_L g447 ( 
.A1(n_419),
.A2(n_423),
.B1(n_424),
.B2(n_448),
.Y(n_447)
);

INVx1_ASAP7_75t_L g448 ( 
.A(n_419),
.Y(n_448)
);

INVx2_ASAP7_75t_L g420 ( 
.A(n_421),
.Y(n_420)
);

INVx3_ASAP7_75t_L g421 ( 
.A(n_422),
.Y(n_421)
);

INVx3_ASAP7_75t_L g456 ( 
.A(n_422),
.Y(n_456)
);

INVx1_ASAP7_75t_L g423 ( 
.A(n_424),
.Y(n_423)
);

OAI21xp5_ASAP7_75t_L g425 ( 
.A1(n_426),
.A2(n_444),
.B(n_449),
.Y(n_425)
);

AOI21xp5_ASAP7_75t_L g426 ( 
.A1(n_427),
.A2(n_436),
.B(n_443),
.Y(n_426)
);

NAND2xp5_ASAP7_75t_SL g427 ( 
.A(n_428),
.B(n_435),
.Y(n_427)
);

NOR2xp33_ASAP7_75t_L g443 ( 
.A(n_428),
.B(n_435),
.Y(n_443)
);

XNOR2xp5_ASAP7_75t_L g428 ( 
.A(n_429),
.B(n_432),
.Y(n_428)
);

NOR2xp33_ASAP7_75t_L g445 ( 
.A(n_429),
.B(n_432),
.Y(n_445)
);

INVx2_ASAP7_75t_L g430 ( 
.A(n_431),
.Y(n_430)
);

INVx3_ASAP7_75t_SL g433 ( 
.A(n_434),
.Y(n_433)
);

NOR2xp33_ASAP7_75t_L g436 ( 
.A(n_437),
.B(n_441),
.Y(n_436)
);

INVx1_ASAP7_75t_SL g438 ( 
.A(n_439),
.Y(n_438)
);

INVx3_ASAP7_75t_L g439 ( 
.A(n_440),
.Y(n_439)
);

NOR2xp33_ASAP7_75t_L g444 ( 
.A(n_445),
.B(n_446),
.Y(n_444)
);

NAND2xp5_ASAP7_75t_L g449 ( 
.A(n_445),
.B(n_446),
.Y(n_449)
);

NOR2xp33_ASAP7_75t_L g451 ( 
.A(n_452),
.B(n_453),
.Y(n_451)
);

NAND2xp5_ASAP7_75t_L g463 ( 
.A(n_452),
.B(n_453),
.Y(n_463)
);

XNOR2xp5_ASAP7_75t_L g453 ( 
.A(n_454),
.B(n_459),
.Y(n_453)
);

OAI22xp5_ASAP7_75t_SL g466 ( 
.A1(n_454),
.A2(n_467),
.B1(n_468),
.B2(n_469),
.Y(n_466)
);

INVx1_ASAP7_75t_L g467 ( 
.A(n_454),
.Y(n_467)
);

MAJIxp5_ASAP7_75t_L g475 ( 
.A(n_454),
.B(n_460),
.C(n_461),
.Y(n_475)
);

FAx1_ASAP7_75t_SL g454 ( 
.A(n_455),
.B(n_457),
.CI(n_458),
.CON(n_454),
.SN(n_454)
);

XNOR2xp5_ASAP7_75t_L g459 ( 
.A(n_460),
.B(n_461),
.Y(n_459)
);

NAND2xp5_ASAP7_75t_SL g464 ( 
.A(n_465),
.B(n_475),
.Y(n_464)
);

NOR2xp33_ASAP7_75t_L g476 ( 
.A(n_465),
.B(n_475),
.Y(n_476)
);

XOR2xp5_ASAP7_75t_L g465 ( 
.A(n_466),
.B(n_472),
.Y(n_465)
);

MAJIxp5_ASAP7_75t_L g478 ( 
.A(n_467),
.B(n_469),
.C(n_472),
.Y(n_478)
);

INVx1_ASAP7_75t_L g468 ( 
.A(n_469),
.Y(n_468)
);

INVx1_ASAP7_75t_L g471 ( 
.A(n_470),
.Y(n_471)
);

NOR2xp33_ASAP7_75t_L g477 ( 
.A(n_478),
.B(n_479),
.Y(n_477)
);

NAND2xp5_ASAP7_75t_L g481 ( 
.A(n_478),
.B(n_479),
.Y(n_481)
);

NAND2xp5_ASAP7_75t_L g492 ( 
.A(n_493),
.B(n_494),
.Y(n_492)
);

NOR2xp33_ASAP7_75t_L g496 ( 
.A(n_493),
.B(n_494),
.Y(n_496)
);

INVx6_ASAP7_75t_L g497 ( 
.A(n_498),
.Y(n_497)
);

INVx6_ASAP7_75t_L g500 ( 
.A(n_498),
.Y(n_500)
);

NOR2xp33_ASAP7_75t_L g499 ( 
.A(n_500),
.B(n_501),
.Y(n_499)
);


endmodule