module fake_jpeg_30046_n_457 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_457);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_457;

wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_385;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_377;
wire n_291;
wire n_236;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_17;
wire n_431;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_415;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_256;
wire n_221;
wire n_454;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_349;
wire n_21;
wire n_288;
wire n_393;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_429;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_305;
wire n_161;
wire n_441;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_382;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_389;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_384;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_199;
wire n_260;
wire n_413;
wire n_275;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_379;
wire n_114;
wire n_444;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_183;
wire n_409;
wire n_249;
wire n_412;
wire n_217;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_391;
wire n_209;
wire n_22;
wire n_138;
wire n_402;
wire n_438;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_4),
.Y(n_17)
);

BUFx12f_ASAP7_75t_L g18 ( 
.A(n_5),
.Y(n_18)
);

CKINVDCx16_ASAP7_75t_R g19 ( 
.A(n_15),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_7),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_3),
.Y(n_21)
);

BUFx12f_ASAP7_75t_L g22 ( 
.A(n_5),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_12),
.Y(n_23)
);

BUFx4f_ASAP7_75t_SL g24 ( 
.A(n_2),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_14),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_10),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_11),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_14),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_12),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_2),
.Y(n_30)
);

HB1xp67_ASAP7_75t_L g31 ( 
.A(n_16),
.Y(n_31)
);

INVx2_ASAP7_75t_L g32 ( 
.A(n_11),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_16),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_3),
.Y(n_34)
);

BUFx4f_ASAP7_75t_SL g35 ( 
.A(n_11),
.Y(n_35)
);

BUFx8_ASAP7_75t_L g36 ( 
.A(n_13),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_4),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_15),
.Y(n_38)
);

BUFx3_ASAP7_75t_L g39 ( 
.A(n_5),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_8),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_8),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_7),
.Y(n_42)
);

INVx2_ASAP7_75t_L g43 ( 
.A(n_7),
.Y(n_43)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_9),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_10),
.Y(n_45)
);

BUFx3_ASAP7_75t_L g46 ( 
.A(n_39),
.Y(n_46)
);

INVx4_ASAP7_75t_L g95 ( 
.A(n_46),
.Y(n_95)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_21),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g100 ( 
.A(n_47),
.Y(n_100)
);

INVx11_ASAP7_75t_L g48 ( 
.A(n_21),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g102 ( 
.A(n_48),
.Y(n_102)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_31),
.Y(n_49)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_49),
.Y(n_93)
);

INVx3_ASAP7_75t_L g50 ( 
.A(n_39),
.Y(n_50)
);

INVx3_ASAP7_75t_L g94 ( 
.A(n_50),
.Y(n_94)
);

BUFx10_ASAP7_75t_L g51 ( 
.A(n_24),
.Y(n_51)
);

INVx2_ASAP7_75t_SL g96 ( 
.A(n_51),
.Y(n_96)
);

INVx3_ASAP7_75t_L g52 ( 
.A(n_39),
.Y(n_52)
);

INVx3_ASAP7_75t_L g118 ( 
.A(n_52),
.Y(n_118)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_21),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g103 ( 
.A(n_53),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_33),
.B(n_16),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g113 ( 
.A(n_54),
.B(n_63),
.Y(n_113)
);

INVx2_ASAP7_75t_L g55 ( 
.A(n_32),
.Y(n_55)
);

INVx2_ASAP7_75t_L g104 ( 
.A(n_55),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_L g56 ( 
.A(n_33),
.B(n_15),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_L g108 ( 
.A(n_56),
.B(n_78),
.Y(n_108)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_42),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g106 ( 
.A(n_57),
.Y(n_106)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_42),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g115 ( 
.A(n_58),
.Y(n_115)
);

INVx5_ASAP7_75t_L g59 ( 
.A(n_42),
.Y(n_59)
);

INVx5_ASAP7_75t_L g129 ( 
.A(n_59),
.Y(n_129)
);

INVx8_ASAP7_75t_L g60 ( 
.A(n_36),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g131 ( 
.A(n_60),
.Y(n_131)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_31),
.Y(n_61)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_61),
.Y(n_124)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_23),
.Y(n_62)
);

INVx5_ASAP7_75t_L g148 ( 
.A(n_62),
.Y(n_148)
);

CKINVDCx20_ASAP7_75t_R g63 ( 
.A(n_36),
.Y(n_63)
);

INVx4_ASAP7_75t_SL g64 ( 
.A(n_32),
.Y(n_64)
);

CKINVDCx14_ASAP7_75t_R g97 ( 
.A(n_64),
.Y(n_97)
);

BUFx12_ASAP7_75t_L g65 ( 
.A(n_24),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g139 ( 
.A(n_65),
.B(n_68),
.Y(n_139)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_23),
.Y(n_66)
);

INVx3_ASAP7_75t_L g125 ( 
.A(n_66),
.Y(n_125)
);

INVx3_ASAP7_75t_L g67 ( 
.A(n_18),
.Y(n_67)
);

INVx3_ASAP7_75t_L g126 ( 
.A(n_67),
.Y(n_126)
);

CKINVDCx20_ASAP7_75t_R g68 ( 
.A(n_36),
.Y(n_68)
);

INVx3_ASAP7_75t_L g69 ( 
.A(n_18),
.Y(n_69)
);

INVx3_ASAP7_75t_L g128 ( 
.A(n_69),
.Y(n_128)
);

BUFx12f_ASAP7_75t_L g70 ( 
.A(n_23),
.Y(n_70)
);

BUFx12f_ASAP7_75t_L g119 ( 
.A(n_70),
.Y(n_119)
);

CKINVDCx20_ASAP7_75t_R g71 ( 
.A(n_36),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_SL g146 ( 
.A(n_71),
.B(n_75),
.Y(n_146)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_25),
.Y(n_72)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_72),
.Y(n_130)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_25),
.Y(n_73)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_73),
.Y(n_132)
);

INVx1_ASAP7_75t_SL g74 ( 
.A(n_43),
.Y(n_74)
);

CKINVDCx14_ASAP7_75t_R g123 ( 
.A(n_74),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_19),
.B(n_14),
.Y(n_75)
);

BUFx6f_ASAP7_75t_L g76 ( 
.A(n_29),
.Y(n_76)
);

BUFx3_ASAP7_75t_L g134 ( 
.A(n_76),
.Y(n_134)
);

BUFx4f_ASAP7_75t_L g77 ( 
.A(n_24),
.Y(n_77)
);

INVx4_ASAP7_75t_L g101 ( 
.A(n_77),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_19),
.B(n_13),
.Y(n_78)
);

BUFx16f_ASAP7_75t_L g79 ( 
.A(n_24),
.Y(n_79)
);

BUFx12f_ASAP7_75t_L g136 ( 
.A(n_79),
.Y(n_136)
);

CKINVDCx20_ASAP7_75t_R g80 ( 
.A(n_36),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_L g110 ( 
.A(n_80),
.B(n_84),
.Y(n_110)
);

BUFx6f_ASAP7_75t_L g81 ( 
.A(n_29),
.Y(n_81)
);

INVx4_ASAP7_75t_L g120 ( 
.A(n_81),
.Y(n_120)
);

INVx2_ASAP7_75t_L g82 ( 
.A(n_43),
.Y(n_82)
);

INVx2_ASAP7_75t_L g116 ( 
.A(n_82),
.Y(n_116)
);

INVx3_ASAP7_75t_L g83 ( 
.A(n_18),
.Y(n_83)
);

INVx4_ASAP7_75t_L g141 ( 
.A(n_83),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_SL g84 ( 
.A(n_28),
.B(n_13),
.Y(n_84)
);

INVx3_ASAP7_75t_L g85 ( 
.A(n_18),
.Y(n_85)
);

INVx4_ASAP7_75t_L g142 ( 
.A(n_85),
.Y(n_142)
);

INVx3_ASAP7_75t_SL g86 ( 
.A(n_29),
.Y(n_86)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_86),
.Y(n_133)
);

INVx5_ASAP7_75t_L g87 ( 
.A(n_38),
.Y(n_87)
);

INVx4_ASAP7_75t_L g145 ( 
.A(n_87),
.Y(n_145)
);

INVx1_ASAP7_75t_SL g88 ( 
.A(n_27),
.Y(n_88)
);

INVx1_ASAP7_75t_SL g99 ( 
.A(n_88),
.Y(n_99)
);

INVx11_ASAP7_75t_SL g89 ( 
.A(n_35),
.Y(n_89)
);

INVx4_ASAP7_75t_L g147 ( 
.A(n_89),
.Y(n_147)
);

BUFx6f_ASAP7_75t_L g90 ( 
.A(n_38),
.Y(n_90)
);

INVx2_ASAP7_75t_L g121 ( 
.A(n_90),
.Y(n_121)
);

BUFx6f_ASAP7_75t_L g91 ( 
.A(n_38),
.Y(n_91)
);

INVx2_ASAP7_75t_L g140 ( 
.A(n_91),
.Y(n_140)
);

CKINVDCx20_ASAP7_75t_R g92 ( 
.A(n_28),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_L g117 ( 
.A(n_92),
.B(n_30),
.Y(n_117)
);

AOI22xp33_ASAP7_75t_SL g98 ( 
.A1(n_86),
.A2(n_18),
.B1(n_22),
.B2(n_44),
.Y(n_98)
);

OAI22xp5_ASAP7_75t_L g149 ( 
.A1(n_98),
.A2(n_109),
.B1(n_111),
.B2(n_112),
.Y(n_149)
);

AOI22xp5_ASAP7_75t_SL g105 ( 
.A1(n_74),
.A2(n_34),
.B1(n_40),
.B2(n_37),
.Y(n_105)
);

AND2x2_ASAP7_75t_L g182 ( 
.A(n_105),
.B(n_46),
.Y(n_182)
);

A2O1A1Ixp33_ASAP7_75t_L g107 ( 
.A1(n_79),
.A2(n_44),
.B(n_27),
.C(n_45),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_SL g167 ( 
.A(n_107),
.B(n_12),
.Y(n_167)
);

AOI22xp33_ASAP7_75t_SL g109 ( 
.A1(n_60),
.A2(n_22),
.B1(n_41),
.B2(n_40),
.Y(n_109)
);

OAI22xp5_ASAP7_75t_L g111 ( 
.A1(n_62),
.A2(n_45),
.B1(n_41),
.B2(n_37),
.Y(n_111)
);

OAI22xp5_ASAP7_75t_L g112 ( 
.A1(n_66),
.A2(n_34),
.B1(n_30),
.B2(n_26),
.Y(n_112)
);

OA22x2_ASAP7_75t_L g114 ( 
.A1(n_88),
.A2(n_35),
.B1(n_22),
.B2(n_26),
.Y(n_114)
);

AOI22x1_ASAP7_75t_L g201 ( 
.A1(n_114),
.A2(n_137),
.B1(n_4),
.B2(n_5),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_L g153 ( 
.A(n_117),
.B(n_108),
.Y(n_153)
);

AOI22xp33_ASAP7_75t_L g122 ( 
.A1(n_76),
.A2(n_22),
.B1(n_20),
.B2(n_17),
.Y(n_122)
);

AOI22xp33_ASAP7_75t_L g151 ( 
.A1(n_122),
.A2(n_91),
.B1(n_90),
.B2(n_58),
.Y(n_151)
);

AO22x1_ASAP7_75t_L g127 ( 
.A1(n_77),
.A2(n_79),
.B1(n_89),
.B2(n_64),
.Y(n_127)
);

O2A1O1Ixp33_ASAP7_75t_L g197 ( 
.A1(n_127),
.A2(n_0),
.B(n_1),
.C(n_3),
.Y(n_197)
);

AOI22xp33_ASAP7_75t_SL g135 ( 
.A1(n_87),
.A2(n_22),
.B1(n_20),
.B2(n_17),
.Y(n_135)
);

AOI22xp33_ASAP7_75t_SL g155 ( 
.A1(n_135),
.A2(n_143),
.B1(n_144),
.B2(n_59),
.Y(n_155)
);

OAI22xp33_ASAP7_75t_SL g137 ( 
.A1(n_81),
.A2(n_35),
.B1(n_1),
.B2(n_2),
.Y(n_137)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_67),
.Y(n_138)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_138),
.Y(n_165)
);

AOI22xp33_ASAP7_75t_SL g143 ( 
.A1(n_70),
.A2(n_35),
.B1(n_1),
.B2(n_2),
.Y(n_143)
);

AOI22xp33_ASAP7_75t_SL g144 ( 
.A1(n_70),
.A2(n_0),
.B1(n_1),
.B2(n_3),
.Y(n_144)
);

INVx11_ASAP7_75t_L g150 ( 
.A(n_131),
.Y(n_150)
);

INVx2_ASAP7_75t_L g207 ( 
.A(n_150),
.Y(n_207)
);

OAI22xp5_ASAP7_75t_SL g241 ( 
.A1(n_151),
.A2(n_181),
.B1(n_185),
.B2(n_6),
.Y(n_241)
);

O2A1O1Ixp33_ASAP7_75t_SL g152 ( 
.A1(n_114),
.A2(n_77),
.B(n_51),
.C(n_65),
.Y(n_152)
);

AOI21xp5_ASAP7_75t_L g216 ( 
.A1(n_152),
.A2(n_168),
.B(n_6),
.Y(n_216)
);

NAND2xp5_ASAP7_75t_SL g217 ( 
.A(n_153),
.B(n_154),
.Y(n_217)
);

CKINVDCx20_ASAP7_75t_R g154 ( 
.A(n_139),
.Y(n_154)
);

INVxp67_ASAP7_75t_L g225 ( 
.A(n_155),
.Y(n_225)
);

INVx2_ASAP7_75t_L g156 ( 
.A(n_126),
.Y(n_156)
);

INVx2_ASAP7_75t_L g222 ( 
.A(n_156),
.Y(n_222)
);

INVxp67_ASAP7_75t_L g157 ( 
.A(n_127),
.Y(n_157)
);

NOR2xp33_ASAP7_75t_L g204 ( 
.A(n_157),
.B(n_169),
.Y(n_204)
);

INVxp33_ASAP7_75t_L g158 ( 
.A(n_123),
.Y(n_158)
);

INVxp67_ASAP7_75t_L g234 ( 
.A(n_158),
.Y(n_234)
);

INVx2_ASAP7_75t_SL g159 ( 
.A(n_94),
.Y(n_159)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_159),
.Y(n_211)
);

INVx8_ASAP7_75t_L g160 ( 
.A(n_131),
.Y(n_160)
);

BUFx2_ASAP7_75t_L g244 ( 
.A(n_160),
.Y(n_244)
);

NAND2xp5_ASAP7_75t_L g161 ( 
.A(n_130),
.B(n_53),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_L g209 ( 
.A(n_161),
.B(n_170),
.Y(n_209)
);

CKINVDCx20_ASAP7_75t_R g162 ( 
.A(n_134),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_SL g219 ( 
.A(n_162),
.B(n_167),
.Y(n_219)
);

HB1xp67_ASAP7_75t_L g163 ( 
.A(n_118),
.Y(n_163)
);

INVx2_ASAP7_75t_L g236 ( 
.A(n_163),
.Y(n_236)
);

INVx2_ASAP7_75t_L g164 ( 
.A(n_128),
.Y(n_164)
);

INVx4_ASAP7_75t_L g238 ( 
.A(n_164),
.Y(n_238)
);

INVxp33_ASAP7_75t_L g166 ( 
.A(n_123),
.Y(n_166)
);

CKINVDCx16_ASAP7_75t_R g226 ( 
.A(n_166),
.Y(n_226)
);

NAND2x1_ASAP7_75t_SL g168 ( 
.A(n_114),
.B(n_99),
.Y(n_168)
);

CKINVDCx16_ASAP7_75t_R g169 ( 
.A(n_132),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_L g170 ( 
.A(n_110),
.B(n_47),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_L g171 ( 
.A(n_93),
.B(n_57),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_L g215 ( 
.A(n_171),
.B(n_179),
.Y(n_215)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_124),
.Y(n_172)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_172),
.Y(n_220)
);

NOR2xp33_ASAP7_75t_L g173 ( 
.A(n_146),
.B(n_65),
.Y(n_173)
);

NOR2xp33_ASAP7_75t_L g210 ( 
.A(n_173),
.B(n_177),
.Y(n_210)
);

CKINVDCx20_ASAP7_75t_R g174 ( 
.A(n_134),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_SL g224 ( 
.A(n_174),
.B(n_178),
.Y(n_224)
);

BUFx12f_ASAP7_75t_L g175 ( 
.A(n_129),
.Y(n_175)
);

INVx3_ASAP7_75t_L g242 ( 
.A(n_175),
.Y(n_242)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_104),
.Y(n_176)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_176),
.Y(n_237)
);

INVxp67_ASAP7_75t_L g177 ( 
.A(n_143),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_L g178 ( 
.A(n_113),
.B(n_51),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_L g179 ( 
.A(n_116),
.B(n_85),
.Y(n_179)
);

CKINVDCx16_ASAP7_75t_R g180 ( 
.A(n_109),
.Y(n_180)
);

NOR2xp33_ASAP7_75t_L g212 ( 
.A(n_180),
.B(n_183),
.Y(n_212)
);

AOI22xp33_ASAP7_75t_SL g181 ( 
.A1(n_97),
.A2(n_50),
.B1(n_52),
.B2(n_133),
.Y(n_181)
);

OAI21xp5_ASAP7_75t_L g227 ( 
.A1(n_182),
.A2(n_197),
.B(n_136),
.Y(n_227)
);

INVxp67_ASAP7_75t_L g183 ( 
.A(n_98),
.Y(n_183)
);

INVx2_ASAP7_75t_L g184 ( 
.A(n_141),
.Y(n_184)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_184),
.Y(n_240)
);

AOI22xp33_ASAP7_75t_SL g185 ( 
.A1(n_97),
.A2(n_83),
.B1(n_69),
.B2(n_48),
.Y(n_185)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_142),
.Y(n_186)
);

NOR2xp33_ASAP7_75t_L g246 ( 
.A(n_186),
.B(n_187),
.Y(n_246)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_121),
.Y(n_187)
);

AND2x2_ASAP7_75t_L g188 ( 
.A(n_101),
.B(n_0),
.Y(n_188)
);

MAJIxp5_ASAP7_75t_L g247 ( 
.A(n_188),
.B(n_11),
.C(n_9),
.Y(n_247)
);

INVx4_ASAP7_75t_L g189 ( 
.A(n_147),
.Y(n_189)
);

HB1xp67_ASAP7_75t_L g206 ( 
.A(n_189),
.Y(n_206)
);

BUFx2_ASAP7_75t_L g190 ( 
.A(n_95),
.Y(n_190)
);

CKINVDCx20_ASAP7_75t_R g203 ( 
.A(n_190),
.Y(n_203)
);

INVx3_ASAP7_75t_L g191 ( 
.A(n_119),
.Y(n_191)
);

INVx8_ASAP7_75t_L g228 ( 
.A(n_191),
.Y(n_228)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_140),
.Y(n_192)
);

CKINVDCx20_ASAP7_75t_R g221 ( 
.A(n_192),
.Y(n_221)
);

INVx2_ASAP7_75t_L g193 ( 
.A(n_125),
.Y(n_193)
);

CKINVDCx20_ASAP7_75t_R g235 ( 
.A(n_193),
.Y(n_235)
);

BUFx6f_ASAP7_75t_L g194 ( 
.A(n_100),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_L g218 ( 
.A(n_194),
.B(n_195),
.Y(n_218)
);

NAND2xp5_ASAP7_75t_L g195 ( 
.A(n_137),
.B(n_0),
.Y(n_195)
);

INVx3_ASAP7_75t_L g196 ( 
.A(n_119),
.Y(n_196)
);

NAND2xp5_ASAP7_75t_L g231 ( 
.A(n_196),
.B(n_198),
.Y(n_231)
);

INVx3_ASAP7_75t_L g198 ( 
.A(n_119),
.Y(n_198)
);

INVx3_ASAP7_75t_L g199 ( 
.A(n_136),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_L g245 ( 
.A(n_199),
.B(n_200),
.Y(n_245)
);

INVx3_ASAP7_75t_SL g200 ( 
.A(n_145),
.Y(n_200)
);

AOI22xp5_ASAP7_75t_L g205 ( 
.A1(n_201),
.A2(n_96),
.B1(n_144),
.B2(n_148),
.Y(n_205)
);

NAND2xp5_ASAP7_75t_L g202 ( 
.A(n_96),
.B(n_4),
.Y(n_202)
);

NOR2xp33_ASAP7_75t_SL g229 ( 
.A(n_202),
.B(n_6),
.Y(n_229)
);

AND2x2_ASAP7_75t_L g250 ( 
.A(n_205),
.B(n_216),
.Y(n_250)
);

AOI22xp5_ASAP7_75t_L g208 ( 
.A1(n_149),
.A2(n_120),
.B1(n_103),
.B2(n_115),
.Y(n_208)
);

OAI22xp5_ASAP7_75t_L g252 ( 
.A1(n_208),
.A2(n_223),
.B1(n_159),
.B2(n_188),
.Y(n_252)
);

AO22x2_ASAP7_75t_L g213 ( 
.A1(n_183),
.A2(n_135),
.B1(n_115),
.B2(n_106),
.Y(n_213)
);

NAND2xp5_ASAP7_75t_L g258 ( 
.A(n_213),
.B(n_197),
.Y(n_258)
);

AOI32xp33_ASAP7_75t_L g214 ( 
.A1(n_177),
.A2(n_122),
.A3(n_136),
.B1(n_100),
.B2(n_106),
.Y(n_214)
);

NOR2xp33_ASAP7_75t_L g249 ( 
.A(n_214),
.B(n_230),
.Y(n_249)
);

AOI22xp5_ASAP7_75t_L g223 ( 
.A1(n_152),
.A2(n_103),
.B1(n_102),
.B2(n_8),
.Y(n_223)
);

AND2x2_ASAP7_75t_L g282 ( 
.A(n_227),
.B(n_233),
.Y(n_282)
);

NAND2xp5_ASAP7_75t_SL g251 ( 
.A(n_229),
.B(n_232),
.Y(n_251)
);

OAI32xp33_ASAP7_75t_L g230 ( 
.A1(n_195),
.A2(n_170),
.A3(n_168),
.B1(n_161),
.B2(n_201),
.Y(n_230)
);

NOR2xp33_ASAP7_75t_SL g232 ( 
.A(n_158),
.B(n_6),
.Y(n_232)
);

OA21x2_ASAP7_75t_L g233 ( 
.A1(n_201),
.A2(n_102),
.B(n_7),
.Y(n_233)
);

NOR2xp33_ASAP7_75t_SL g239 ( 
.A(n_166),
.B(n_157),
.Y(n_239)
);

NAND2xp5_ASAP7_75t_SL g283 ( 
.A(n_239),
.B(n_243),
.Y(n_283)
);

INVxp67_ASAP7_75t_L g269 ( 
.A(n_241),
.Y(n_269)
);

NOR2xp33_ASAP7_75t_SL g243 ( 
.A(n_171),
.B(n_8),
.Y(n_243)
);

MAJx2_ASAP7_75t_L g275 ( 
.A(n_247),
.B(n_9),
.C(n_10),
.Y(n_275)
);

AOI22xp5_ASAP7_75t_L g248 ( 
.A1(n_216),
.A2(n_182),
.B1(n_188),
.B2(n_193),
.Y(n_248)
);

OAI22xp5_ASAP7_75t_SL g303 ( 
.A1(n_248),
.A2(n_256),
.B1(n_260),
.B2(n_266),
.Y(n_303)
);

AOI22xp5_ASAP7_75t_L g293 ( 
.A1(n_252),
.A2(n_262),
.B1(n_234),
.B2(n_203),
.Y(n_293)
);

NOR2xp33_ASAP7_75t_L g253 ( 
.A(n_224),
.B(n_165),
.Y(n_253)
);

CKINVDCx14_ASAP7_75t_R g297 ( 
.A(n_253),
.Y(n_297)
);

HAxp5_ASAP7_75t_SL g254 ( 
.A(n_219),
.B(n_182),
.CON(n_254),
.SN(n_254)
);

INVxp67_ASAP7_75t_L g309 ( 
.A(n_254),
.Y(n_309)
);

CKINVDCx20_ASAP7_75t_R g255 ( 
.A(n_231),
.Y(n_255)
);

OR2x2_ASAP7_75t_L g294 ( 
.A(n_255),
.B(n_263),
.Y(n_294)
);

AOI22xp5_ASAP7_75t_L g256 ( 
.A1(n_225),
.A2(n_159),
.B1(n_160),
.B2(n_194),
.Y(n_256)
);

MAJIxp5_ASAP7_75t_L g257 ( 
.A(n_209),
.B(n_164),
.C(n_156),
.Y(n_257)
);

MAJIxp5_ASAP7_75t_L g318 ( 
.A(n_257),
.B(n_277),
.C(n_248),
.Y(n_318)
);

OAI21xp5_ASAP7_75t_SL g289 ( 
.A1(n_258),
.A2(n_213),
.B(n_234),
.Y(n_289)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_211),
.Y(n_259)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_259),
.Y(n_288)
);

AOI22xp5_ASAP7_75t_L g260 ( 
.A1(n_225),
.A2(n_200),
.B1(n_150),
.B2(n_184),
.Y(n_260)
);

INVx2_ASAP7_75t_L g261 ( 
.A(n_222),
.Y(n_261)
);

INVx1_ASAP7_75t_SL g319 ( 
.A(n_261),
.Y(n_319)
);

OAI22xp5_ASAP7_75t_L g262 ( 
.A1(n_205),
.A2(n_190),
.B1(n_189),
.B2(n_196),
.Y(n_262)
);

CKINVDCx20_ASAP7_75t_R g263 ( 
.A(n_231),
.Y(n_263)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_211),
.Y(n_264)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_264),
.Y(n_308)
);

NAND2xp5_ASAP7_75t_L g265 ( 
.A(n_209),
.B(n_175),
.Y(n_265)
);

NAND2xp5_ASAP7_75t_L g317 ( 
.A(n_265),
.B(n_271),
.Y(n_317)
);

AOI22xp5_ASAP7_75t_L g266 ( 
.A1(n_230),
.A2(n_191),
.B1(n_198),
.B2(n_199),
.Y(n_266)
);

CKINVDCx20_ASAP7_75t_R g267 ( 
.A(n_245),
.Y(n_267)
);

NAND2xp5_ASAP7_75t_SL g312 ( 
.A(n_267),
.B(n_280),
.Y(n_312)
);

INVx2_ASAP7_75t_L g268 ( 
.A(n_222),
.Y(n_268)
);

HB1xp67_ASAP7_75t_L g300 ( 
.A(n_268),
.Y(n_300)
);

BUFx2_ASAP7_75t_L g270 ( 
.A(n_228),
.Y(n_270)
);

INVx3_ASAP7_75t_L g306 ( 
.A(n_270),
.Y(n_306)
);

NAND2xp5_ASAP7_75t_L g271 ( 
.A(n_215),
.B(n_243),
.Y(n_271)
);

NAND2xp5_ASAP7_75t_L g272 ( 
.A(n_215),
.B(n_175),
.Y(n_272)
);

NAND2xp5_ASAP7_75t_L g322 ( 
.A(n_272),
.B(n_284),
.Y(n_322)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_237),
.Y(n_273)
);

CKINVDCx16_ASAP7_75t_R g299 ( 
.A(n_273),
.Y(n_299)
);

OAI21xp5_ASAP7_75t_L g274 ( 
.A1(n_227),
.A2(n_9),
.B(n_10),
.Y(n_274)
);

OAI21xp5_ASAP7_75t_L g304 ( 
.A1(n_274),
.A2(n_281),
.B(n_282),
.Y(n_304)
);

XNOR2xp5_ASAP7_75t_L g307 ( 
.A(n_275),
.B(n_206),
.Y(n_307)
);

NOR2xp33_ASAP7_75t_L g276 ( 
.A(n_217),
.B(n_204),
.Y(n_276)
);

NOR2xp33_ASAP7_75t_SL g311 ( 
.A(n_276),
.B(n_286),
.Y(n_311)
);

MAJIxp5_ASAP7_75t_L g277 ( 
.A(n_210),
.B(n_212),
.C(n_239),
.Y(n_277)
);

CKINVDCx5p33_ASAP7_75t_R g278 ( 
.A(n_226),
.Y(n_278)
);

NOR2xp33_ASAP7_75t_L g290 ( 
.A(n_278),
.B(n_285),
.Y(n_290)
);

AOI22xp5_ASAP7_75t_L g279 ( 
.A1(n_241),
.A2(n_233),
.B1(n_213),
.B2(n_208),
.Y(n_279)
);

OAI22xp5_ASAP7_75t_SL g314 ( 
.A1(n_279),
.A2(n_207),
.B1(n_242),
.B2(n_228),
.Y(n_314)
);

INVxp67_ASAP7_75t_L g280 ( 
.A(n_245),
.Y(n_280)
);

OAI21xp5_ASAP7_75t_L g281 ( 
.A1(n_233),
.A2(n_232),
.B(n_218),
.Y(n_281)
);

NAND2xp5_ASAP7_75t_L g284 ( 
.A(n_218),
.B(n_229),
.Y(n_284)
);

INVxp33_ASAP7_75t_L g285 ( 
.A(n_246),
.Y(n_285)
);

NOR2xp33_ASAP7_75t_L g286 ( 
.A(n_220),
.B(n_221),
.Y(n_286)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_237),
.Y(n_287)
);

NOR2xp33_ASAP7_75t_L g291 ( 
.A(n_287),
.B(n_221),
.Y(n_291)
);

NAND2xp5_ASAP7_75t_SL g337 ( 
.A(n_289),
.B(n_256),
.Y(n_337)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_291),
.Y(n_326)
);

AOI22xp33_ASAP7_75t_L g292 ( 
.A1(n_262),
.A2(n_252),
.B1(n_269),
.B2(n_281),
.Y(n_292)
);

INVxp67_ASAP7_75t_L g331 ( 
.A(n_292),
.Y(n_331)
);

OA22x2_ASAP7_75t_L g338 ( 
.A1(n_293),
.A2(n_295),
.B1(n_310),
.B2(n_260),
.Y(n_338)
);

AOI22xp5_ASAP7_75t_L g295 ( 
.A1(n_269),
.A2(n_213),
.B1(n_223),
.B2(n_220),
.Y(n_295)
);

OAI22xp5_ASAP7_75t_L g296 ( 
.A1(n_279),
.A2(n_213),
.B1(n_247),
.B2(n_244),
.Y(n_296)
);

AOI22xp5_ASAP7_75t_L g325 ( 
.A1(n_296),
.A2(n_302),
.B1(n_314),
.B2(n_303),
.Y(n_325)
);

CKINVDCx20_ASAP7_75t_R g298 ( 
.A(n_270),
.Y(n_298)
);

CKINVDCx20_ASAP7_75t_R g323 ( 
.A(n_298),
.Y(n_323)
);

AO22x1_ASAP7_75t_SL g301 ( 
.A1(n_258),
.A2(n_240),
.B1(n_238),
.B2(n_236),
.Y(n_301)
);

NAND2xp5_ASAP7_75t_L g329 ( 
.A(n_301),
.B(n_267),
.Y(n_329)
);

OAI22xp5_ASAP7_75t_L g302 ( 
.A1(n_249),
.A2(n_244),
.B1(n_235),
.B2(n_203),
.Y(n_302)
);

INVxp67_ASAP7_75t_L g347 ( 
.A(n_304),
.Y(n_347)
);

XOR2xp5_ASAP7_75t_L g305 ( 
.A(n_265),
.B(n_271),
.Y(n_305)
);

MAJIxp5_ASAP7_75t_L g327 ( 
.A(n_305),
.B(n_316),
.C(n_272),
.Y(n_327)
);

XNOR2xp5_ASAP7_75t_SL g340 ( 
.A(n_307),
.B(n_313),
.Y(n_340)
);

AOI22xp5_ASAP7_75t_L g310 ( 
.A1(n_250),
.A2(n_235),
.B1(n_236),
.B2(n_240),
.Y(n_310)
);

XNOR2xp5_ASAP7_75t_L g313 ( 
.A(n_284),
.B(n_238),
.Y(n_313)
);

AOI22xp5_ASAP7_75t_SL g315 ( 
.A1(n_282),
.A2(n_207),
.B1(n_242),
.B2(n_250),
.Y(n_315)
);

OAI21xp5_ASAP7_75t_SL g324 ( 
.A1(n_315),
.A2(n_320),
.B(n_280),
.Y(n_324)
);

XOR2xp5_ASAP7_75t_L g316 ( 
.A(n_277),
.B(n_257),
.Y(n_316)
);

XNOR2x1_ASAP7_75t_L g342 ( 
.A(n_318),
.B(n_251),
.Y(n_342)
);

AOI22xp5_ASAP7_75t_SL g320 ( 
.A1(n_282),
.A2(n_250),
.B1(n_263),
.B2(n_255),
.Y(n_320)
);

CKINVDCx20_ASAP7_75t_R g321 ( 
.A(n_270),
.Y(n_321)
);

CKINVDCx20_ASAP7_75t_R g346 ( 
.A(n_321),
.Y(n_346)
);

AOI21xp5_ASAP7_75t_L g357 ( 
.A1(n_324),
.A2(n_328),
.B(n_337),
.Y(n_357)
);

OAI22xp5_ASAP7_75t_L g367 ( 
.A1(n_325),
.A2(n_349),
.B1(n_350),
.B2(n_351),
.Y(n_367)
);

MAJIxp5_ASAP7_75t_L g368 ( 
.A(n_327),
.B(n_342),
.C(n_309),
.Y(n_368)
);

OAI21xp5_ASAP7_75t_SL g328 ( 
.A1(n_315),
.A2(n_274),
.B(n_283),
.Y(n_328)
);

NAND2xp5_ASAP7_75t_L g356 ( 
.A(n_329),
.B(n_334),
.Y(n_356)
);

AOI22xp5_ASAP7_75t_L g330 ( 
.A1(n_314),
.A2(n_266),
.B1(n_264),
.B2(n_259),
.Y(n_330)
);

OAI22xp5_ASAP7_75t_SL g355 ( 
.A1(n_330),
.A2(n_343),
.B1(n_293),
.B2(n_295),
.Y(n_355)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_288),
.Y(n_332)
);

INVx1_ASAP7_75t_L g354 ( 
.A(n_332),
.Y(n_354)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_288),
.Y(n_333)
);

INVx1_ASAP7_75t_L g360 ( 
.A(n_333),
.Y(n_360)
);

NAND2xp5_ASAP7_75t_L g334 ( 
.A(n_294),
.B(n_287),
.Y(n_334)
);

CKINVDCx20_ASAP7_75t_R g335 ( 
.A(n_294),
.Y(n_335)
);

NAND2xp5_ASAP7_75t_L g366 ( 
.A(n_335),
.B(n_341),
.Y(n_366)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_308),
.Y(n_336)
);

INVx1_ASAP7_75t_L g361 ( 
.A(n_336),
.Y(n_361)
);

INVx2_ASAP7_75t_SL g370 ( 
.A(n_338),
.Y(n_370)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_308),
.Y(n_339)
);

INVx1_ASAP7_75t_L g369 ( 
.A(n_339),
.Y(n_369)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_312),
.Y(n_341)
);

AOI22xp5_ASAP7_75t_L g343 ( 
.A1(n_303),
.A2(n_273),
.B1(n_278),
.B2(n_261),
.Y(n_343)
);

INVx1_ASAP7_75t_L g344 ( 
.A(n_300),
.Y(n_344)
);

CKINVDCx16_ASAP7_75t_R g372 ( 
.A(n_344),
.Y(n_372)
);

XNOR2xp5_ASAP7_75t_SL g345 ( 
.A(n_305),
.B(n_275),
.Y(n_345)
);

XOR2xp5_ASAP7_75t_L g364 ( 
.A(n_345),
.B(n_307),
.Y(n_364)
);

OAI21xp5_ASAP7_75t_SL g348 ( 
.A1(n_309),
.A2(n_268),
.B(n_304),
.Y(n_348)
);

CKINVDCx20_ASAP7_75t_R g359 ( 
.A(n_348),
.Y(n_359)
);

NOR2xp33_ASAP7_75t_SL g349 ( 
.A(n_297),
.B(n_311),
.Y(n_349)
);

INVx1_ASAP7_75t_L g350 ( 
.A(n_301),
.Y(n_350)
);

INVx1_ASAP7_75t_L g351 ( 
.A(n_301),
.Y(n_351)
);

XNOR2xp5_ASAP7_75t_L g352 ( 
.A(n_340),
.B(n_327),
.Y(n_352)
);

XNOR2xp5_ASAP7_75t_L g382 ( 
.A(n_352),
.B(n_358),
.Y(n_382)
);

FAx1_ASAP7_75t_SL g353 ( 
.A(n_334),
.B(n_322),
.CI(n_317),
.CON(n_353),
.SN(n_353)
);

NAND2xp5_ASAP7_75t_L g380 ( 
.A(n_353),
.B(n_355),
.Y(n_380)
);

XNOR2xp5_ASAP7_75t_L g358 ( 
.A(n_340),
.B(n_316),
.Y(n_358)
);

OAI22xp5_ASAP7_75t_SL g362 ( 
.A1(n_331),
.A2(n_320),
.B1(n_322),
.B2(n_317),
.Y(n_362)
);

INVx1_ASAP7_75t_L g383 ( 
.A(n_362),
.Y(n_383)
);

XNOR2xp5_ASAP7_75t_L g363 ( 
.A(n_342),
.B(n_318),
.Y(n_363)
);

XNOR2xp5_ASAP7_75t_L g397 ( 
.A(n_363),
.B(n_365),
.Y(n_397)
);

XNOR2xp5_ASAP7_75t_SL g389 ( 
.A(n_364),
.B(n_375),
.Y(n_389)
);

XNOR2xp5_ASAP7_75t_L g365 ( 
.A(n_345),
.B(n_313),
.Y(n_365)
);

XOR2xp5_ASAP7_75t_L g384 ( 
.A(n_368),
.B(n_374),
.Y(n_384)
);

AOI22xp5_ASAP7_75t_SL g371 ( 
.A1(n_331),
.A2(n_289),
.B1(n_310),
.B2(n_298),
.Y(n_371)
);

OAI22xp5_ASAP7_75t_SL g393 ( 
.A1(n_371),
.A2(n_330),
.B1(n_343),
.B2(n_351),
.Y(n_393)
);

MAJIxp5_ASAP7_75t_L g373 ( 
.A(n_347),
.B(n_299),
.C(n_290),
.Y(n_373)
);

MAJIxp5_ASAP7_75t_L g377 ( 
.A(n_373),
.B(n_376),
.C(n_328),
.Y(n_377)
);

XNOR2xp5_ASAP7_75t_L g374 ( 
.A(n_348),
.B(n_319),
.Y(n_374)
);

XOR2xp5_ASAP7_75t_L g375 ( 
.A(n_324),
.B(n_319),
.Y(n_375)
);

MAJIxp5_ASAP7_75t_L g376 ( 
.A(n_347),
.B(n_321),
.C(n_306),
.Y(n_376)
);

XNOR2xp5_ASAP7_75t_L g404 ( 
.A(n_377),
.B(n_375),
.Y(n_404)
);

CKINVDCx14_ASAP7_75t_R g378 ( 
.A(n_366),
.Y(n_378)
);

NAND2xp5_ASAP7_75t_L g407 ( 
.A(n_378),
.B(n_379),
.Y(n_407)
);

NOR2xp33_ASAP7_75t_SL g379 ( 
.A(n_353),
.B(n_341),
.Y(n_379)
);

NOR2xp33_ASAP7_75t_L g381 ( 
.A(n_353),
.B(n_326),
.Y(n_381)
);

NAND2xp5_ASAP7_75t_L g411 ( 
.A(n_381),
.B(n_387),
.Y(n_411)
);

MAJIxp5_ASAP7_75t_L g385 ( 
.A(n_363),
.B(n_325),
.C(n_338),
.Y(n_385)
);

MAJIxp5_ASAP7_75t_L g401 ( 
.A(n_385),
.B(n_388),
.C(n_390),
.Y(n_401)
);

INVx1_ASAP7_75t_L g386 ( 
.A(n_354),
.Y(n_386)
);

INVx1_ASAP7_75t_L g405 ( 
.A(n_386),
.Y(n_405)
);

HB1xp67_ASAP7_75t_L g387 ( 
.A(n_367),
.Y(n_387)
);

MAJIxp5_ASAP7_75t_L g388 ( 
.A(n_352),
.B(n_338),
.C(n_329),
.Y(n_388)
);

MAJIxp5_ASAP7_75t_L g390 ( 
.A(n_358),
.B(n_338),
.C(n_326),
.Y(n_390)
);

CKINVDCx20_ASAP7_75t_R g391 ( 
.A(n_356),
.Y(n_391)
);

NAND2xp5_ASAP7_75t_SL g399 ( 
.A(n_391),
.B(n_396),
.Y(n_399)
);

XNOR2xp5_ASAP7_75t_SL g392 ( 
.A(n_365),
.B(n_364),
.Y(n_392)
);

XOR2xp5_ASAP7_75t_L g409 ( 
.A(n_392),
.B(n_357),
.Y(n_409)
);

NAND2xp5_ASAP7_75t_L g406 ( 
.A(n_393),
.B(n_355),
.Y(n_406)
);

INVx1_ASAP7_75t_L g394 ( 
.A(n_360),
.Y(n_394)
);

INVx1_ASAP7_75t_SL g402 ( 
.A(n_394),
.Y(n_402)
);

MAJIxp5_ASAP7_75t_L g395 ( 
.A(n_368),
.B(n_350),
.C(n_344),
.Y(n_395)
);

MAJIxp5_ASAP7_75t_L g403 ( 
.A(n_395),
.B(n_397),
.C(n_384),
.Y(n_403)
);

AOI21xp5_ASAP7_75t_L g396 ( 
.A1(n_374),
.A2(n_323),
.B(n_346),
.Y(n_396)
);

OAI22xp5_ASAP7_75t_L g398 ( 
.A1(n_380),
.A2(n_370),
.B1(n_359),
.B2(n_357),
.Y(n_398)
);

INVx1_ASAP7_75t_L g418 ( 
.A(n_398),
.Y(n_418)
);

NAND2xp5_ASAP7_75t_SL g400 ( 
.A(n_388),
.B(n_373),
.Y(n_400)
);

NOR2xp33_ASAP7_75t_L g421 ( 
.A(n_400),
.B(n_389),
.Y(n_421)
);

MAJIxp5_ASAP7_75t_L g417 ( 
.A(n_403),
.B(n_382),
.C(n_397),
.Y(n_417)
);

XNOR2xp5_ASAP7_75t_L g423 ( 
.A(n_404),
.B(n_392),
.Y(n_423)
);

NAND2xp5_ASAP7_75t_L g422 ( 
.A(n_406),
.B(n_408),
.Y(n_422)
);

NOR2xp33_ASAP7_75t_L g408 ( 
.A(n_383),
.B(n_362),
.Y(n_408)
);

XOR2xp5_ASAP7_75t_L g424 ( 
.A(n_409),
.B(n_369),
.Y(n_424)
);

OAI22xp5_ASAP7_75t_SL g410 ( 
.A1(n_385),
.A2(n_370),
.B1(n_371),
.B2(n_376),
.Y(n_410)
);

AOI22xp5_ASAP7_75t_L g419 ( 
.A1(n_410),
.A2(n_389),
.B1(n_382),
.B2(n_361),
.Y(n_419)
);

HB1xp67_ASAP7_75t_L g412 ( 
.A(n_384),
.Y(n_412)
);

INVx1_ASAP7_75t_L g425 ( 
.A(n_412),
.Y(n_425)
);

NOR2xp33_ASAP7_75t_L g413 ( 
.A(n_395),
.B(n_372),
.Y(n_413)
);

CKINVDCx20_ASAP7_75t_R g420 ( 
.A(n_413),
.Y(n_420)
);

INVx2_ASAP7_75t_L g414 ( 
.A(n_393),
.Y(n_414)
);

NOR2xp33_ASAP7_75t_L g427 ( 
.A(n_414),
.B(n_333),
.Y(n_427)
);

OAI21xp5_ASAP7_75t_SL g415 ( 
.A1(n_399),
.A2(n_390),
.B(n_377),
.Y(n_415)
);

INVxp67_ASAP7_75t_L g429 ( 
.A(n_415),
.Y(n_429)
);

OAI21xp5_ASAP7_75t_L g416 ( 
.A1(n_406),
.A2(n_346),
.B(n_323),
.Y(n_416)
);

AOI21xp5_ASAP7_75t_SL g437 ( 
.A1(n_416),
.A2(n_402),
.B(n_336),
.Y(n_437)
);

MAJIxp5_ASAP7_75t_L g433 ( 
.A(n_417),
.B(n_401),
.C(n_411),
.Y(n_433)
);

XOR2xp5_ASAP7_75t_L g436 ( 
.A(n_419),
.B(n_423),
.Y(n_436)
);

NOR2xp33_ASAP7_75t_L g431 ( 
.A(n_421),
.B(n_404),
.Y(n_431)
);

XNOR2x1_ASAP7_75t_L g428 ( 
.A(n_424),
.B(n_409),
.Y(n_428)
);

XNOR2xp5_ASAP7_75t_L g426 ( 
.A(n_401),
.B(n_332),
.Y(n_426)
);

XOR2xp5_ASAP7_75t_L g435 ( 
.A(n_426),
.B(n_407),
.Y(n_435)
);

INVx1_ASAP7_75t_L g434 ( 
.A(n_427),
.Y(n_434)
);

XNOR2xp5_ASAP7_75t_L g441 ( 
.A(n_428),
.B(n_435),
.Y(n_441)
);

XNOR2xp5_ASAP7_75t_L g430 ( 
.A(n_417),
.B(n_403),
.Y(n_430)
);

NAND2xp5_ASAP7_75t_L g444 ( 
.A(n_430),
.B(n_423),
.Y(n_444)
);

NAND2xp5_ASAP7_75t_L g442 ( 
.A(n_431),
.B(n_432),
.Y(n_442)
);

AOI22xp5_ASAP7_75t_L g432 ( 
.A1(n_418),
.A2(n_414),
.B1(n_410),
.B2(n_402),
.Y(n_432)
);

MAJIxp5_ASAP7_75t_L g443 ( 
.A(n_433),
.B(n_426),
.C(n_415),
.Y(n_443)
);

OAI21x1_ASAP7_75t_L g440 ( 
.A1(n_437),
.A2(n_422),
.B(n_339),
.Y(n_440)
);

NOR2xp33_ASAP7_75t_SL g438 ( 
.A(n_429),
.B(n_420),
.Y(n_438)
);

NOR2xp33_ASAP7_75t_L g447 ( 
.A(n_438),
.B(n_440),
.Y(n_447)
);

OR2x2_ASAP7_75t_L g439 ( 
.A(n_434),
.B(n_416),
.Y(n_439)
);

INVx1_ASAP7_75t_L g446 ( 
.A(n_439),
.Y(n_446)
);

NOR2xp33_ASAP7_75t_L g448 ( 
.A(n_443),
.B(n_444),
.Y(n_448)
);

OA21x2_ASAP7_75t_SL g445 ( 
.A1(n_442),
.A2(n_429),
.B(n_422),
.Y(n_445)
);

INVxp33_ASAP7_75t_L g451 ( 
.A(n_445),
.Y(n_451)
);

MAJIxp5_ASAP7_75t_L g449 ( 
.A(n_448),
.B(n_441),
.C(n_439),
.Y(n_449)
);

NAND2xp5_ASAP7_75t_SL g453 ( 
.A(n_449),
.B(n_447),
.Y(n_453)
);

NAND4xp25_ASAP7_75t_SL g450 ( 
.A(n_446),
.B(n_419),
.C(n_425),
.D(n_405),
.Y(n_450)
);

NAND2xp5_ASAP7_75t_L g452 ( 
.A(n_450),
.B(n_446),
.Y(n_452)
);

OAI21xp5_ASAP7_75t_L g454 ( 
.A1(n_452),
.A2(n_453),
.B(n_437),
.Y(n_454)
);

OAI321xp33_ASAP7_75t_L g455 ( 
.A1(n_454),
.A2(n_451),
.A3(n_428),
.B1(n_424),
.B2(n_436),
.C(n_306),
.Y(n_455)
);

INVx1_ASAP7_75t_L g456 ( 
.A(n_455),
.Y(n_456)
);

NOR2xp33_ASAP7_75t_L g457 ( 
.A(n_456),
.B(n_436),
.Y(n_457)
);


endmodule