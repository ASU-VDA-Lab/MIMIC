module fake_jpeg_22811_n_328 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_328);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_328;

wire n_253;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_260;
wire n_199;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_7),
.Y(n_17)
);

NOR2xp33_ASAP7_75t_L g18 ( 
.A(n_9),
.B(n_14),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_6),
.Y(n_19)
);

INVx6_ASAP7_75t_L g20 ( 
.A(n_7),
.Y(n_20)
);

BUFx5_ASAP7_75t_L g21 ( 
.A(n_2),
.Y(n_21)
);

BUFx16f_ASAP7_75t_L g22 ( 
.A(n_6),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_8),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_3),
.Y(n_24)
);

NOR2xp33_ASAP7_75t_L g25 ( 
.A(n_9),
.B(n_15),
.Y(n_25)
);

INVx13_ASAP7_75t_L g26 ( 
.A(n_10),
.Y(n_26)
);

BUFx5_ASAP7_75t_L g27 ( 
.A(n_2),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_6),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_4),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_1),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_5),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_1),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_10),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_12),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_11),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_16),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_14),
.Y(n_37)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_14),
.Y(n_38)
);

INVx11_ASAP7_75t_L g39 ( 
.A(n_26),
.Y(n_39)
);

INVx11_ASAP7_75t_L g62 ( 
.A(n_39),
.Y(n_62)
);

BUFx2_ASAP7_75t_L g40 ( 
.A(n_22),
.Y(n_40)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_40),
.Y(n_75)
);

INVx2_ASAP7_75t_L g41 ( 
.A(n_22),
.Y(n_41)
);

INVx6_ASAP7_75t_L g59 ( 
.A(n_41),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_L g42 ( 
.A(n_32),
.B(n_0),
.Y(n_42)
);

AND2x2_ASAP7_75t_L g76 ( 
.A(n_42),
.B(n_0),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g43 ( 
.A(n_18),
.B(n_8),
.Y(n_43)
);

OAI21xp5_ASAP7_75t_L g69 ( 
.A1(n_43),
.A2(n_45),
.B(n_38),
.Y(n_69)
);

INVx2_ASAP7_75t_L g44 ( 
.A(n_22),
.Y(n_44)
);

INVx6_ASAP7_75t_L g63 ( 
.A(n_44),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_SL g45 ( 
.A(n_18),
.B(n_25),
.Y(n_45)
);

INVx4_ASAP7_75t_L g46 ( 
.A(n_26),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_46),
.B(n_49),
.Y(n_53)
);

INVx2_ASAP7_75t_SL g47 ( 
.A(n_21),
.Y(n_47)
);

AOI22xp33_ASAP7_75t_SL g54 ( 
.A1(n_47),
.A2(n_20),
.B1(n_26),
.B2(n_27),
.Y(n_54)
);

INVx5_ASAP7_75t_L g48 ( 
.A(n_20),
.Y(n_48)
);

INVx5_ASAP7_75t_L g61 ( 
.A(n_48),
.Y(n_61)
);

BUFx8_ASAP7_75t_L g49 ( 
.A(n_21),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_21),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_50),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_L g52 ( 
.A(n_45),
.B(n_34),
.Y(n_52)
);

AND2x2_ASAP7_75t_L g117 ( 
.A(n_52),
.B(n_55),
.Y(n_117)
);

CKINVDCx14_ASAP7_75t_R g91 ( 
.A(n_54),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_L g55 ( 
.A(n_42),
.B(n_34),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_48),
.Y(n_56)
);

CKINVDCx16_ASAP7_75t_R g100 ( 
.A(n_56),
.Y(n_100)
);

OAI22xp5_ASAP7_75t_L g57 ( 
.A1(n_42),
.A2(n_20),
.B1(n_26),
.B2(n_38),
.Y(n_57)
);

AOI22xp5_ASAP7_75t_L g99 ( 
.A1(n_57),
.A2(n_23),
.B1(n_29),
.B2(n_33),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_43),
.B(n_25),
.Y(n_58)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_58),
.Y(n_93)
);

BUFx3_ASAP7_75t_L g60 ( 
.A(n_40),
.Y(n_60)
);

CKINVDCx14_ASAP7_75t_R g108 ( 
.A(n_60),
.Y(n_108)
);

INVx2_ASAP7_75t_L g64 ( 
.A(n_48),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_64),
.B(n_65),
.Y(n_82)
);

INVx3_ASAP7_75t_L g65 ( 
.A(n_39),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_41),
.B(n_22),
.Y(n_66)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_66),
.Y(n_97)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_48),
.Y(n_67)
);

BUFx2_ASAP7_75t_L g111 ( 
.A(n_67),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_L g68 ( 
.A(n_50),
.B(n_34),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_SL g86 ( 
.A(n_68),
.B(n_71),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_SL g114 ( 
.A(n_69),
.B(n_17),
.Y(n_114)
);

BUFx12f_ASAP7_75t_L g70 ( 
.A(n_40),
.Y(n_70)
);

BUFx3_ASAP7_75t_L g109 ( 
.A(n_70),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_L g71 ( 
.A(n_50),
.B(n_38),
.Y(n_71)
);

BUFx3_ASAP7_75t_L g72 ( 
.A(n_40),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_72),
.B(n_74),
.Y(n_84)
);

AOI22xp5_ASAP7_75t_L g73 ( 
.A1(n_47),
.A2(n_20),
.B1(n_17),
.B2(n_31),
.Y(n_73)
);

OAI22xp5_ASAP7_75t_SL g87 ( 
.A1(n_73),
.A2(n_23),
.B1(n_29),
.B2(n_33),
.Y(n_87)
);

INVx2_ASAP7_75t_L g74 ( 
.A(n_50),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_L g83 ( 
.A(n_76),
.B(n_23),
.Y(n_83)
);

BUFx6f_ASAP7_75t_L g77 ( 
.A(n_47),
.Y(n_77)
);

INVx4_ASAP7_75t_L g106 ( 
.A(n_77),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_41),
.B(n_22),
.Y(n_78)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_78),
.Y(n_105)
);

BUFx6f_ASAP7_75t_L g79 ( 
.A(n_47),
.Y(n_79)
);

INVx2_ASAP7_75t_L g88 ( 
.A(n_79),
.Y(n_88)
);

BUFx3_ASAP7_75t_L g80 ( 
.A(n_47),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_80),
.B(n_81),
.Y(n_92)
);

INVx3_ASAP7_75t_L g81 ( 
.A(n_39),
.Y(n_81)
);

NOR2x1_ASAP7_75t_R g150 ( 
.A(n_83),
.B(n_49),
.Y(n_150)
);

CKINVDCx20_ASAP7_75t_R g85 ( 
.A(n_60),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_SL g130 ( 
.A(n_85),
.B(n_101),
.Y(n_130)
);

OAI22xp33_ASAP7_75t_SL g132 ( 
.A1(n_87),
.A2(n_36),
.B1(n_35),
.B2(n_30),
.Y(n_132)
);

AOI22xp33_ASAP7_75t_L g89 ( 
.A1(n_76),
.A2(n_27),
.B1(n_17),
.B2(n_35),
.Y(n_89)
);

OAI22xp5_ASAP7_75t_L g122 ( 
.A1(n_89),
.A2(n_90),
.B1(n_99),
.B2(n_104),
.Y(n_122)
);

OAI22xp5_ASAP7_75t_L g90 ( 
.A1(n_54),
.A2(n_44),
.B1(n_39),
.B2(n_27),
.Y(n_90)
);

MAJIxp5_ASAP7_75t_L g94 ( 
.A(n_75),
.B(n_44),
.C(n_49),
.Y(n_94)
);

MAJIxp5_ASAP7_75t_L g153 ( 
.A(n_94),
.B(n_119),
.C(n_79),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_59),
.B(n_36),
.Y(n_95)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_95),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_L g96 ( 
.A(n_69),
.B(n_59),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g123 ( 
.A(n_96),
.B(n_113),
.Y(n_123)
);

INVx2_ASAP7_75t_L g98 ( 
.A(n_80),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g146 ( 
.A(n_98),
.B(n_103),
.Y(n_146)
);

CKINVDCx20_ASAP7_75t_R g101 ( 
.A(n_72),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_63),
.B(n_31),
.Y(n_102)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_102),
.Y(n_121)
);

INVx2_ASAP7_75t_L g103 ( 
.A(n_70),
.Y(n_103)
);

AOI22xp33_ASAP7_75t_SL g104 ( 
.A1(n_61),
.A2(n_29),
.B1(n_33),
.B2(n_32),
.Y(n_104)
);

INVx2_ASAP7_75t_L g107 ( 
.A(n_70),
.Y(n_107)
);

INVx1_ASAP7_75t_SL g128 ( 
.A(n_107),
.Y(n_128)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_53),
.Y(n_110)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_110),
.Y(n_131)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_65),
.Y(n_112)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_112),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_L g113 ( 
.A(n_63),
.B(n_32),
.Y(n_113)
);

CKINVDCx14_ASAP7_75t_R g148 ( 
.A(n_114),
.Y(n_148)
);

OAI22xp5_ASAP7_75t_L g115 ( 
.A1(n_61),
.A2(n_46),
.B1(n_19),
.B2(n_37),
.Y(n_115)
);

OAI22xp5_ASAP7_75t_L g140 ( 
.A1(n_115),
.A2(n_116),
.B1(n_24),
.B2(n_19),
.Y(n_140)
);

OAI22xp5_ASAP7_75t_L g116 ( 
.A1(n_81),
.A2(n_46),
.B1(n_19),
.B2(n_37),
.Y(n_116)
);

INVx2_ASAP7_75t_L g118 ( 
.A(n_51),
.Y(n_118)
);

INVx2_ASAP7_75t_L g136 ( 
.A(n_118),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_L g119 ( 
.A(n_62),
.B(n_37),
.Y(n_119)
);

AOI21xp33_ASAP7_75t_L g124 ( 
.A1(n_96),
.A2(n_83),
.B(n_114),
.Y(n_124)
);

OAI21xp5_ASAP7_75t_SL g169 ( 
.A1(n_124),
.A2(n_125),
.B(n_134),
.Y(n_169)
);

OAI21xp5_ASAP7_75t_L g125 ( 
.A1(n_91),
.A2(n_30),
.B(n_28),
.Y(n_125)
);

INVxp67_ASAP7_75t_L g126 ( 
.A(n_92),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_L g158 ( 
.A(n_126),
.B(n_129),
.Y(n_158)
);

AOI22xp33_ASAP7_75t_SL g127 ( 
.A1(n_110),
.A2(n_62),
.B1(n_46),
.B2(n_28),
.Y(n_127)
);

AOI21xp5_ASAP7_75t_L g170 ( 
.A1(n_127),
.A2(n_106),
.B(n_88),
.Y(n_170)
);

INVx13_ASAP7_75t_L g129 ( 
.A(n_109),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_SL g174 ( 
.A(n_132),
.B(n_138),
.Y(n_174)
);

AOI32xp33_ASAP7_75t_L g134 ( 
.A1(n_94),
.A2(n_49),
.A3(n_67),
.B1(n_56),
.B2(n_51),
.Y(n_134)
);

OAI22xp5_ASAP7_75t_SL g135 ( 
.A1(n_99),
.A2(n_37),
.B1(n_24),
.B2(n_19),
.Y(n_135)
);

AOI22xp5_ASAP7_75t_L g160 ( 
.A1(n_135),
.A2(n_140),
.B1(n_100),
.B2(n_118),
.Y(n_160)
);

INVxp67_ASAP7_75t_L g137 ( 
.A(n_109),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_L g173 ( 
.A(n_137),
.B(n_141),
.Y(n_173)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_113),
.Y(n_138)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_82),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_SL g159 ( 
.A(n_139),
.B(n_152),
.Y(n_159)
);

INVx2_ASAP7_75t_L g141 ( 
.A(n_116),
.Y(n_141)
);

AND2x2_ASAP7_75t_SL g142 ( 
.A(n_119),
.B(n_49),
.Y(n_142)
);

MAJIxp5_ASAP7_75t_L g157 ( 
.A(n_142),
.B(n_86),
.C(n_112),
.Y(n_157)
);

INVxp67_ASAP7_75t_L g143 ( 
.A(n_84),
.Y(n_143)
);

NOR2xp33_ASAP7_75t_L g179 ( 
.A(n_143),
.B(n_144),
.Y(n_179)
);

INVx2_ASAP7_75t_L g144 ( 
.A(n_115),
.Y(n_144)
);

INVxp67_ASAP7_75t_L g145 ( 
.A(n_90),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_L g181 ( 
.A(n_145),
.B(n_147),
.Y(n_181)
);

INVx13_ASAP7_75t_L g147 ( 
.A(n_103),
.Y(n_147)
);

INVx2_ASAP7_75t_L g149 ( 
.A(n_98),
.Y(n_149)
);

NOR2xp33_ASAP7_75t_L g182 ( 
.A(n_149),
.B(n_151),
.Y(n_182)
);

OAI21xp5_ASAP7_75t_SL g180 ( 
.A1(n_150),
.A2(n_49),
.B(n_108),
.Y(n_180)
);

CKINVDCx20_ASAP7_75t_R g151 ( 
.A(n_85),
.Y(n_151)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_111),
.Y(n_152)
);

XNOR2xp5_ASAP7_75t_L g187 ( 
.A(n_153),
.B(n_24),
.Y(n_187)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_111),
.Y(n_154)
);

NOR2xp33_ASAP7_75t_L g185 ( 
.A(n_154),
.B(n_111),
.Y(n_185)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_130),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_L g199 ( 
.A(n_155),
.B(n_177),
.Y(n_199)
);

AND2x2_ASAP7_75t_L g156 ( 
.A(n_123),
.B(n_87),
.Y(n_156)
);

OAI21xp5_ASAP7_75t_SL g214 ( 
.A1(n_156),
.A2(n_180),
.B(n_0),
.Y(n_214)
);

XNOR2xp5_ASAP7_75t_L g193 ( 
.A(n_157),
.B(n_125),
.Y(n_193)
);

OAI22xp5_ASAP7_75t_L g202 ( 
.A1(n_160),
.A2(n_167),
.B1(n_136),
.B2(n_133),
.Y(n_202)
);

NAND2xp5_ASAP7_75t_L g161 ( 
.A(n_123),
.B(n_117),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_L g189 ( 
.A(n_161),
.B(n_162),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_L g162 ( 
.A(n_138),
.B(n_117),
.Y(n_162)
);

OAI22xp5_ASAP7_75t_SL g163 ( 
.A1(n_145),
.A2(n_97),
.B1(n_105),
.B2(n_117),
.Y(n_163)
);

OAI22xp5_ASAP7_75t_SL g195 ( 
.A1(n_163),
.A2(n_186),
.B1(n_154),
.B2(n_152),
.Y(n_195)
);

CKINVDCx16_ASAP7_75t_R g164 ( 
.A(n_146),
.Y(n_164)
);

AOI22xp33_ASAP7_75t_SL g188 ( 
.A1(n_164),
.A2(n_165),
.B1(n_171),
.B2(n_178),
.Y(n_188)
);

INVx5_ASAP7_75t_L g165 ( 
.A(n_128),
.Y(n_165)
);

MAJIxp5_ASAP7_75t_L g166 ( 
.A(n_153),
.B(n_105),
.C(n_97),
.Y(n_166)
);

XOR2xp5_ASAP7_75t_L g190 ( 
.A(n_166),
.B(n_187),
.Y(n_190)
);

OAI22xp5_ASAP7_75t_L g167 ( 
.A1(n_144),
.A2(n_100),
.B1(n_106),
.B2(n_88),
.Y(n_167)
);

BUFx12f_ASAP7_75t_L g168 ( 
.A(n_128),
.Y(n_168)
);

INVx3_ASAP7_75t_L g203 ( 
.A(n_168),
.Y(n_203)
);

AOI22xp33_ASAP7_75t_L g211 ( 
.A1(n_170),
.A2(n_129),
.B1(n_149),
.B2(n_137),
.Y(n_211)
);

CKINVDCx16_ASAP7_75t_R g171 ( 
.A(n_142),
.Y(n_171)
);

OR2x2_ASAP7_75t_L g172 ( 
.A(n_150),
.B(n_101),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_L g206 ( 
.A(n_172),
.B(n_176),
.Y(n_206)
);

CKINVDCx20_ASAP7_75t_R g175 ( 
.A(n_151),
.Y(n_175)
);

CKINVDCx20_ASAP7_75t_R g191 ( 
.A(n_175),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_L g176 ( 
.A(n_142),
.B(n_93),
.Y(n_176)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_133),
.Y(n_177)
);

CKINVDCx16_ASAP7_75t_R g178 ( 
.A(n_135),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_L g183 ( 
.A(n_148),
.B(n_93),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_L g210 ( 
.A(n_183),
.B(n_147),
.Y(n_210)
);

NOR2xp33_ASAP7_75t_SL g184 ( 
.A(n_131),
.B(n_10),
.Y(n_184)
);

NOR2xp33_ASAP7_75t_SL g213 ( 
.A(n_184),
.B(n_8),
.Y(n_213)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_185),
.Y(n_194)
);

OAI22xp5_ASAP7_75t_SL g186 ( 
.A1(n_141),
.A2(n_24),
.B1(n_107),
.B2(n_77),
.Y(n_186)
);

XOR2xp5_ASAP7_75t_L g192 ( 
.A(n_187),
.B(n_122),
.Y(n_192)
);

MAJIxp5_ASAP7_75t_L g241 ( 
.A(n_192),
.B(n_155),
.C(n_3),
.Y(n_241)
);

XNOR2xp5_ASAP7_75t_L g221 ( 
.A(n_193),
.B(n_157),
.Y(n_221)
);

AOI22xp5_ASAP7_75t_L g239 ( 
.A1(n_195),
.A2(n_202),
.B1(n_207),
.B2(n_177),
.Y(n_239)
);

CKINVDCx14_ASAP7_75t_R g196 ( 
.A(n_173),
.Y(n_196)
);

NAND2xp5_ASAP7_75t_L g234 ( 
.A(n_196),
.B(n_197),
.Y(n_234)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_182),
.Y(n_197)
);

OAI22x1_ASAP7_75t_SL g198 ( 
.A1(n_172),
.A2(n_126),
.B1(n_143),
.B2(n_131),
.Y(n_198)
);

OAI22xp5_ASAP7_75t_L g222 ( 
.A1(n_198),
.A2(n_211),
.B1(n_170),
.B2(n_179),
.Y(n_222)
);

NOR2x1_ASAP7_75t_L g200 ( 
.A(n_172),
.B(n_139),
.Y(n_200)
);

NAND2xp5_ASAP7_75t_L g238 ( 
.A(n_200),
.B(n_204),
.Y(n_238)
);

NOR2xp33_ASAP7_75t_L g201 ( 
.A(n_175),
.B(n_120),
.Y(n_201)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_201),
.Y(n_225)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_159),
.Y(n_204)
);

CKINVDCx20_ASAP7_75t_R g205 ( 
.A(n_168),
.Y(n_205)
);

CKINVDCx20_ASAP7_75t_R g224 ( 
.A(n_205),
.Y(n_224)
);

OAI22xp5_ASAP7_75t_SL g207 ( 
.A1(n_178),
.A2(n_136),
.B1(n_121),
.B2(n_120),
.Y(n_207)
);

CKINVDCx20_ASAP7_75t_R g208 ( 
.A(n_168),
.Y(n_208)
);

CKINVDCx20_ASAP7_75t_R g226 ( 
.A(n_208),
.Y(n_226)
);

OR2x2_ASAP7_75t_SL g209 ( 
.A(n_171),
.B(n_121),
.Y(n_209)
);

OAI21xp5_ASAP7_75t_L g235 ( 
.A1(n_209),
.A2(n_215),
.B(n_184),
.Y(n_235)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_210),
.Y(n_229)
);

INVxp33_ASAP7_75t_L g212 ( 
.A(n_168),
.Y(n_212)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_212),
.Y(n_237)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_213),
.Y(n_242)
);

OAI21xp5_ASAP7_75t_SL g219 ( 
.A1(n_214),
.A2(n_217),
.B(n_218),
.Y(n_219)
);

AND2x2_ASAP7_75t_SL g215 ( 
.A(n_176),
.B(n_0),
.Y(n_215)
);

CKINVDCx20_ASAP7_75t_R g216 ( 
.A(n_159),
.Y(n_216)
);

CKINVDCx20_ASAP7_75t_R g230 ( 
.A(n_216),
.Y(n_230)
);

NAND2xp5_ASAP7_75t_L g217 ( 
.A(n_161),
.B(n_1),
.Y(n_217)
);

NAND2xp5_ASAP7_75t_L g218 ( 
.A(n_156),
.B(n_1),
.Y(n_218)
);

AOI21xp5_ASAP7_75t_L g220 ( 
.A1(n_206),
.A2(n_181),
.B(n_180),
.Y(n_220)
);

OAI22xp5_ASAP7_75t_L g247 ( 
.A1(n_220),
.A2(n_227),
.B1(n_231),
.B2(n_239),
.Y(n_247)
);

XOR2xp5_ASAP7_75t_L g262 ( 
.A(n_221),
.B(n_228),
.Y(n_262)
);

AOI22xp5_ASAP7_75t_L g253 ( 
.A1(n_222),
.A2(n_223),
.B1(n_236),
.B2(n_243),
.Y(n_253)
);

OAI22xp5_ASAP7_75t_SL g223 ( 
.A1(n_188),
.A2(n_169),
.B1(n_160),
.B2(n_166),
.Y(n_223)
);

OAI21xp5_ASAP7_75t_SL g227 ( 
.A1(n_206),
.A2(n_169),
.B(n_164),
.Y(n_227)
);

XNOR2xp5_ASAP7_75t_L g228 ( 
.A(n_190),
.B(n_163),
.Y(n_228)
);

OAI21xp5_ASAP7_75t_SL g231 ( 
.A1(n_214),
.A2(n_162),
.B(n_158),
.Y(n_231)
);

XNOR2xp5_ASAP7_75t_L g232 ( 
.A(n_190),
.B(n_183),
.Y(n_232)
);

XNOR2xp5_ASAP7_75t_L g245 ( 
.A(n_232),
.B(n_240),
.Y(n_245)
);

XOR2xp5_ASAP7_75t_L g233 ( 
.A(n_192),
.B(n_156),
.Y(n_233)
);

MAJIxp5_ASAP7_75t_L g250 ( 
.A(n_233),
.B(n_241),
.C(n_215),
.Y(n_250)
);

CKINVDCx14_ASAP7_75t_R g258 ( 
.A(n_235),
.Y(n_258)
);

A2O1A1Ixp33_ASAP7_75t_SL g236 ( 
.A1(n_200),
.A2(n_167),
.B(n_186),
.C(n_165),
.Y(n_236)
);

XNOR2xp5_ASAP7_75t_L g240 ( 
.A(n_193),
.B(n_174),
.Y(n_240)
);

AOI22xp5_ASAP7_75t_L g243 ( 
.A1(n_195),
.A2(n_2),
.B1(n_3),
.B2(n_4),
.Y(n_243)
);

NOR2xp33_ASAP7_75t_L g244 ( 
.A(n_224),
.B(n_191),
.Y(n_244)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_244),
.Y(n_265)
);

INVxp67_ASAP7_75t_SL g246 ( 
.A(n_236),
.Y(n_246)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_246),
.Y(n_272)
);

NAND2xp5_ASAP7_75t_L g248 ( 
.A(n_238),
.B(n_189),
.Y(n_248)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_248),
.Y(n_278)
);

NAND2xp5_ASAP7_75t_L g249 ( 
.A(n_226),
.B(n_191),
.Y(n_249)
);

NAND2xp5_ASAP7_75t_L g277 ( 
.A(n_249),
.B(n_251),
.Y(n_277)
);

MAJIxp5_ASAP7_75t_L g264 ( 
.A(n_250),
.B(n_252),
.C(n_241),
.Y(n_264)
);

NAND2xp5_ASAP7_75t_L g251 ( 
.A(n_225),
.B(n_210),
.Y(n_251)
);

MAJIxp5_ASAP7_75t_L g252 ( 
.A(n_233),
.B(n_189),
.C(n_218),
.Y(n_252)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_234),
.Y(n_254)
);

NAND2xp5_ASAP7_75t_L g279 ( 
.A(n_254),
.B(n_255),
.Y(n_279)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_238),
.Y(n_255)
);

AOI22xp5_ASAP7_75t_L g256 ( 
.A1(n_223),
.A2(n_198),
.B1(n_207),
.B2(n_216),
.Y(n_256)
);

OAI22xp5_ASAP7_75t_SL g273 ( 
.A1(n_256),
.A2(n_263),
.B1(n_219),
.B2(n_243),
.Y(n_273)
);

NOR2xp33_ASAP7_75t_L g257 ( 
.A(n_230),
.B(n_203),
.Y(n_257)
);

NAND2xp5_ASAP7_75t_L g270 ( 
.A(n_257),
.B(n_261),
.Y(n_270)
);

AND2x6_ASAP7_75t_L g259 ( 
.A(n_227),
.B(n_232),
.Y(n_259)
);

OAI21xp5_ASAP7_75t_L g281 ( 
.A1(n_259),
.A2(n_209),
.B(n_217),
.Y(n_281)
);

INVx2_ASAP7_75t_L g260 ( 
.A(n_237),
.Y(n_260)
);

AOI21xp5_ASAP7_75t_L g266 ( 
.A1(n_260),
.A2(n_205),
.B(n_194),
.Y(n_266)
);

HB1xp67_ASAP7_75t_L g261 ( 
.A(n_236),
.Y(n_261)
);

AOI22xp5_ASAP7_75t_L g263 ( 
.A1(n_229),
.A2(n_204),
.B1(n_197),
.B2(n_208),
.Y(n_263)
);

MAJIxp5_ASAP7_75t_L g282 ( 
.A(n_264),
.B(n_267),
.C(n_280),
.Y(n_282)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_266),
.Y(n_289)
);

MAJIxp5_ASAP7_75t_L g267 ( 
.A(n_262),
.B(n_231),
.C(n_221),
.Y(n_267)
);

AOI22xp5_ASAP7_75t_L g268 ( 
.A1(n_247),
.A2(n_236),
.B1(n_239),
.B2(n_203),
.Y(n_268)
);

OAI22xp5_ASAP7_75t_SL g287 ( 
.A1(n_268),
.A2(n_271),
.B1(n_281),
.B2(n_253),
.Y(n_287)
);

XOR2xp5_ASAP7_75t_L g269 ( 
.A(n_262),
.B(n_228),
.Y(n_269)
);

XOR2xp5_ASAP7_75t_L g292 ( 
.A(n_269),
.B(n_275),
.Y(n_292)
);

AOI22xp5_ASAP7_75t_L g271 ( 
.A1(n_258),
.A2(n_220),
.B1(n_219),
.B2(n_194),
.Y(n_271)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_273),
.Y(n_290)
);

NAND2xp5_ASAP7_75t_L g274 ( 
.A(n_248),
.B(n_215),
.Y(n_274)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_274),
.Y(n_291)
);

XOR2xp5_ASAP7_75t_L g275 ( 
.A(n_245),
.B(n_252),
.Y(n_275)
);

XNOR2xp5_ASAP7_75t_L g276 ( 
.A(n_245),
.B(n_250),
.Y(n_276)
);

XNOR2xp5_ASAP7_75t_L g284 ( 
.A(n_276),
.B(n_256),
.Y(n_284)
);

MAJIxp5_ASAP7_75t_L g280 ( 
.A(n_259),
.B(n_240),
.C(n_235),
.Y(n_280)
);

NAND2xp5_ASAP7_75t_L g283 ( 
.A(n_265),
.B(n_199),
.Y(n_283)
);

NAND2xp5_ASAP7_75t_L g300 ( 
.A(n_283),
.B(n_273),
.Y(n_300)
);

MAJIxp5_ASAP7_75t_L g296 ( 
.A(n_284),
.B(n_295),
.C(n_264),
.Y(n_296)
);

OAI22xp5_ASAP7_75t_L g285 ( 
.A1(n_268),
.A2(n_272),
.B1(n_253),
.B2(n_270),
.Y(n_285)
);

CKINVDCx14_ASAP7_75t_R g299 ( 
.A(n_285),
.Y(n_299)
);

HB1xp67_ASAP7_75t_L g286 ( 
.A(n_266),
.Y(n_286)
);

INVxp67_ASAP7_75t_L g305 ( 
.A(n_286),
.Y(n_305)
);

NAND2xp5_ASAP7_75t_SL g303 ( 
.A(n_287),
.B(n_293),
.Y(n_303)
);

AOI22xp5_ASAP7_75t_SL g288 ( 
.A1(n_270),
.A2(n_260),
.B1(n_263),
.B2(n_242),
.Y(n_288)
);

AOI22xp5_ASAP7_75t_SL g302 ( 
.A1(n_288),
.A2(n_294),
.B1(n_9),
.B2(n_11),
.Y(n_302)
);

NOR2xp33_ASAP7_75t_SL g293 ( 
.A(n_277),
.B(n_4),
.Y(n_293)
);

XOR2x1_ASAP7_75t_SL g294 ( 
.A(n_271),
.B(n_5),
.Y(n_294)
);

MAJIxp5_ASAP7_75t_L g295 ( 
.A(n_275),
.B(n_5),
.C(n_7),
.Y(n_295)
);

XNOR2xp5_ASAP7_75t_L g312 ( 
.A(n_296),
.B(n_297),
.Y(n_312)
);

OAI322xp33_ASAP7_75t_L g297 ( 
.A1(n_294),
.A2(n_279),
.A3(n_281),
.B1(n_280),
.B2(n_274),
.C1(n_267),
.C2(n_276),
.Y(n_297)
);

NOR2xp33_ASAP7_75t_L g298 ( 
.A(n_288),
.B(n_278),
.Y(n_298)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_298),
.Y(n_310)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_300),
.Y(n_313)
);

MAJIxp5_ASAP7_75t_L g301 ( 
.A(n_292),
.B(n_282),
.C(n_269),
.Y(n_301)
);

NAND2xp5_ASAP7_75t_L g306 ( 
.A(n_301),
.B(n_292),
.Y(n_306)
);

NOR2xp33_ASAP7_75t_SL g307 ( 
.A(n_302),
.B(n_12),
.Y(n_307)
);

OA21x2_ASAP7_75t_SL g304 ( 
.A1(n_295),
.A2(n_11),
.B(n_12),
.Y(n_304)
);

AOI21x1_ASAP7_75t_SL g308 ( 
.A1(n_304),
.A2(n_13),
.B(n_15),
.Y(n_308)
);

AOI21xp5_ASAP7_75t_L g314 ( 
.A1(n_306),
.A2(n_301),
.B(n_296),
.Y(n_314)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_307),
.Y(n_315)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_308),
.Y(n_317)
);

OR2x2_ASAP7_75t_L g309 ( 
.A(n_302),
.B(n_291),
.Y(n_309)
);

AOI21x1_ASAP7_75t_L g316 ( 
.A1(n_309),
.A2(n_311),
.B(n_305),
.Y(n_316)
);

OR2x2_ASAP7_75t_L g311 ( 
.A(n_305),
.B(n_289),
.Y(n_311)
);

XOR2xp5_ASAP7_75t_L g320 ( 
.A(n_314),
.B(n_318),
.Y(n_320)
);

OAI31xp33_ASAP7_75t_L g321 ( 
.A1(n_316),
.A2(n_309),
.A3(n_311),
.B(n_315),
.Y(n_321)
);

AOI21xp5_ASAP7_75t_L g318 ( 
.A1(n_313),
.A2(n_299),
.B(n_290),
.Y(n_318)
);

NOR2xp33_ASAP7_75t_L g319 ( 
.A(n_310),
.B(n_303),
.Y(n_319)
);

XOR2xp5_ASAP7_75t_L g322 ( 
.A(n_319),
.B(n_312),
.Y(n_322)
);

NAND2xp5_ASAP7_75t_SL g323 ( 
.A(n_321),
.B(n_322),
.Y(n_323)
);

XOR2xp5_ASAP7_75t_L g324 ( 
.A(n_320),
.B(n_282),
.Y(n_324)
);

AOI21xp5_ASAP7_75t_L g325 ( 
.A1(n_324),
.A2(n_284),
.B(n_317),
.Y(n_325)
);

AOI22xp5_ASAP7_75t_SL g326 ( 
.A1(n_325),
.A2(n_323),
.B1(n_15),
.B2(n_16),
.Y(n_326)
);

OAI21xp5_ASAP7_75t_SL g327 ( 
.A1(n_326),
.A2(n_13),
.B(n_16),
.Y(n_327)
);

XNOR2xp5_ASAP7_75t_L g328 ( 
.A(n_327),
.B(n_13),
.Y(n_328)
);


endmodule