module real_aes_6643_n_99 (n_17, n_28, n_76, n_56, n_34, n_98, n_90, n_82, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_83, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_91, n_43, n_96, n_54, n_35, n_42, n_15, n_9, n_23, n_72, n_95, n_44, n_7, n_4, n_80, n_6, n_12, n_68, n_79, n_69, n_46, n_59, n_25, n_73, n_77, n_81, n_48, n_37, n_97, n_70, n_50, n_89, n_26, n_86, n_93, n_13, n_24, n_2, n_55, n_62, n_84, n_67, n_92, n_33, n_88, n_14, n_11, n_85, n_16, n_94, n_39, n_5, n_45, n_60, n_38, n_87, n_0, n_78, n_63, n_1, n_53, n_36, n_99);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_98;
input n_90;
input n_82;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_83;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_91;
input n_43;
input n_96;
input n_54;
input n_35;
input n_42;
input n_15;
input n_9;
input n_23;
input n_72;
input n_95;
input n_44;
input n_7;
input n_4;
input n_80;
input n_6;
input n_12;
input n_68;
input n_79;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_81;
input n_48;
input n_37;
input n_97;
input n_70;
input n_50;
input n_89;
input n_26;
input n_86;
input n_93;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_84;
input n_67;
input n_92;
input n_33;
input n_88;
input n_14;
input n_11;
input n_85;
input n_16;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_87;
input n_0;
input n_78;
input n_63;
input n_1;
input n_53;
input n_36;
output n_99;
wire n_480;
wire n_113;
wire n_476;
wire n_599;
wire n_187;
wire n_436;
wire n_684;
wire n_257;
wire n_390;
wire n_185;
wire n_285;
wire n_624;
wire n_618;
wire n_522;
wire n_485;
wire n_222;
wire n_631;
wire n_503;
wire n_357;
wire n_287;
wire n_635;
wire n_386;
wire n_673;
wire n_518;
wire n_254;
wire n_207;
wire n_665;
wire n_667;
wire n_577;
wire n_580;
wire n_469;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_718;
wire n_318;
wire n_355;
wire n_239;
wire n_669;
wire n_100;
wire n_423;
wire n_458;
wire n_444;
wire n_112;
wire n_319;
wire n_364;
wire n_421;
wire n_555;
wire n_329;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_169;
wire n_242;
wire n_376;
wire n_549;
wire n_571;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_448;
wire n_545;
wire n_341;
wire n_556;
wire n_593;
wire n_232;
wire n_460;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_537;
wire n_320;
wire n_551;
wire n_666;
wire n_560;
wire n_260;
wire n_660;
wire n_594;
wire n_186;
wire n_138;
wire n_696;
wire n_704;
wire n_453;
wire n_374;
wire n_379;
wire n_647;
wire n_235;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_161;
wire n_189;
wire n_271;
wire n_489;
wire n_427;
wire n_548;
wire n_678;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_519;
wire n_564;
wire n_638;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_512;
wire n_395;
wire n_332;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_116;
wire n_625;
wire n_462;
wire n_289;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_716;
wire n_213;
wire n_356;
wire n_478;
wire n_584;
wire n_408;
wire n_553;
wire n_184;
wire n_372;
wire n_528;
wire n_578;
wire n_202;
wire n_495;
wire n_370;
wire n_384;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_467;
wire n_327;
wire n_106;
wire n_466;
wire n_559;
wire n_636;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_517;
wire n_683;
wire n_174;
wire n_570;
wire n_675;
wire n_530;
wire n_104;
wire n_535;
wire n_211;
wire n_281;
wire n_496;
wire n_693;
wire n_173;
wire n_468;
wire n_234;
wire n_284;
wire n_153;
wire n_532;
wire n_316;
wire n_656;
wire n_178;
wire n_409;
wire n_298;
wire n_523;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_297;
wire n_383;
wire n_529;
wire n_119;
wire n_455;
wire n_310;
wire n_504;
wire n_164;
wire n_671;
wire n_231;
wire n_102;
wire n_547;
wire n_659;
wire n_634;
wire n_682;
wire n_454;
wire n_122;
wire n_443;
wire n_565;
wire n_608;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_267;
wire n_218;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_722;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_331;
wire n_182;
wire n_363;
wire n_449;
wire n_417;
wire n_607;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_142;
wire n_561;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_655;
wire n_654;
wire n_505;
wire n_434;
wire n_502;
wire n_527;
wire n_600;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_602;
wire n_402;
wire n_552;
wire n_617;
wire n_171;
wire n_658;
wire n_676;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_432;
wire n_146;
wire n_255;
wire n_226;
wire n_286;
wire n_416;
wire n_410;
wire n_120;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_695;
wire n_685;
wire n_165;
wire n_361;
wire n_632;
wire n_246;
wire n_176;
wire n_412;
wire n_163;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_501;
wire n_488;
wire n_251;
wire n_642;
wire n_613;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_702;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_110;
wire n_392;
wire n_562;
wire n_150;
wire n_147;
wire n_288;
wire n_404;
wire n_598;
wire n_713;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_569;
wire n_563;
wire n_188;
wire n_269;
wire n_430;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_193;
wire n_397;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_649;
wire n_663;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_707;
wire n_622;
wire n_470;
wire n_133;
wire n_494;
wire n_711;
wire n_377;
wire n_273;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_265;
wire n_354;
wire n_720;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_643;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_148;
wire n_481;
wire n_498;
wire n_691;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_487;
wire n_233;
wire n_290;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_155;
wire n_243;
wire n_692;
wire n_544;
wire n_268;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_101;
wire n_701;
wire n_309;
wire n_344;
wire n_107;
wire n_229;
wire n_482;
wire n_520;
wire n_679;
wire n_633;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_262;
wire n_630;
wire n_689;
wire n_715;
wire n_134;
wire n_349;
wire n_336;
wire n_420;
wire n_612;
wire n_195;
wire n_438;
wire n_300;
wire n_252;
wire n_283;
wire n_314;
wire n_249;
wire n_623;
wire n_446;
wire n_721;
wire n_221;
wire n_681;
wire n_156;
wire n_359;
wire n_717;
wire n_456;
wire n_312;
wire n_183;
wire n_266;
wire n_712;
wire n_205;
wire n_433;
wire n_335;
wire n_177;
wire n_516;
wire n_313;
wire n_627;
wire n_140;
wire n_418;
wire n_521;
wire n_422;
wire n_219;
wire n_524;
wire n_705;
wire n_180;
wire n_212;
wire n_210;
wire n_575;
wire n_325;
wire n_338;
wire n_479;
wire n_442;
wire n_698;
wire n_371;
wire n_103;
wire n_166;
wire n_541;
wire n_224;
wire n_151;
wire n_546;
wire n_587;
wire n_639;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_440;
wire n_525;
wire n_644;
wire n_674;
wire n_152;
wire n_198;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_414;
wire n_123;
wire n_279;
wire n_686;
wire n_543;
wire n_497;
wire n_514;
wire n_507;
wire n_270;
wire n_614;
wire n_305;
wire n_586;
wire n_450;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_465;
wire n_473;
wire n_719;
wire n_566;
wire n_474;
wire n_170;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_168;
wire n_175;
wire n_241;
wire n_687;
wire n_646;
wire n_710;
wire n_650;
wire n_105;
wire n_294;
wire n_393;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_500;
wire n_307;
wire n_601;
wire n_661;
wire n_463;
wire n_396;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_143;
wire n_192;
wire n_475;
wire n_554;
wire n_264;
wire n_237;
wire n_668;
AOI222xp33_ASAP7_75t_L g438 ( .A1(n_0), .A2(n_7), .B1(n_439), .B2(n_711), .C1(n_716), .C2(n_717), .Y(n_438) );
INVx1_ASAP7_75t_L g107 ( .A(n_1), .Y(n_107) );
A2O1A1Ixp33_ASAP7_75t_L g181 ( .A1(n_2), .A2(n_140), .B(n_145), .C(n_182), .Y(n_181) );
AOI21xp5_ASAP7_75t_L g204 ( .A1(n_3), .A2(n_135), .B(n_205), .Y(n_204) );
INVx1_ASAP7_75t_L g451 ( .A(n_4), .Y(n_451) );
NAND2xp5_ASAP7_75t_L g212 ( .A(n_5), .B(n_159), .Y(n_212) );
NAND2xp5_ASAP7_75t_SL g434 ( .A(n_6), .B(n_435), .Y(n_434) );
CKINVDCx20_ASAP7_75t_R g716 ( .A(n_7), .Y(n_716) );
AOI21xp33_ASAP7_75t_L g468 ( .A1(n_8), .A2(n_135), .B(n_469), .Y(n_468) );
AND2x6_ASAP7_75t_L g140 ( .A(n_9), .B(n_141), .Y(n_140) );
INVx1_ASAP7_75t_L g169 ( .A(n_10), .Y(n_169) );
INVx1_ASAP7_75t_L g105 ( .A(n_11), .Y(n_105) );
NOR2xp33_ASAP7_75t_L g433 ( .A(n_11), .B(n_44), .Y(n_433) );
AOI21xp5_ASAP7_75t_L g528 ( .A1(n_12), .A2(n_247), .B(n_529), .Y(n_528) );
NAND2xp5_ASAP7_75t_SL g186 ( .A(n_13), .B(n_150), .Y(n_186) );
INVx1_ASAP7_75t_L g473 ( .A(n_14), .Y(n_473) );
NAND2xp5_ASAP7_75t_L g521 ( .A(n_15), .B(n_149), .Y(n_521) );
INVx1_ASAP7_75t_L g133 ( .A(n_16), .Y(n_133) );
INVx1_ASAP7_75t_L g533 ( .A(n_17), .Y(n_533) );
A2O1A1Ixp33_ASAP7_75t_L g194 ( .A1(n_18), .A2(n_170), .B(n_195), .C(n_197), .Y(n_194) );
NAND2xp5_ASAP7_75t_L g198 ( .A(n_19), .B(n_159), .Y(n_198) );
NAND2xp5_ASAP7_75t_L g512 ( .A(n_20), .B(n_462), .Y(n_512) );
NAND2xp5_ASAP7_75t_SL g499 ( .A(n_21), .B(n_135), .Y(n_499) );
NAND2xp5_ASAP7_75t_L g254 ( .A(n_22), .B(n_255), .Y(n_254) );
A2O1A1Ixp33_ASAP7_75t_L g148 ( .A1(n_23), .A2(n_149), .B(n_151), .C(n_155), .Y(n_148) );
AOI22xp5_ASAP7_75t_L g99 ( .A1(n_24), .A2(n_100), .B1(n_111), .B2(n_722), .Y(n_99) );
NAND2xp5_ASAP7_75t_L g465 ( .A(n_25), .B(n_159), .Y(n_465) );
NAND2xp5_ASAP7_75t_SL g219 ( .A(n_26), .B(n_150), .Y(n_219) );
A2O1A1Ixp33_ASAP7_75t_L g531 ( .A1(n_27), .A2(n_153), .B(n_197), .C(n_532), .Y(n_531) );
NAND2xp5_ASAP7_75t_SL g231 ( .A(n_28), .B(n_150), .Y(n_231) );
CKINVDCx16_ASAP7_75t_R g215 ( .A(n_29), .Y(n_215) );
INVx1_ASAP7_75t_L g229 ( .A(n_30), .Y(n_229) );
BUFx6f_ASAP7_75t_L g139 ( .A(n_31), .Y(n_139) );
CKINVDCx20_ASAP7_75t_R g179 ( .A(n_32), .Y(n_179) );
NAND2xp5_ASAP7_75t_L g452 ( .A(n_33), .B(n_150), .Y(n_452) );
INVx1_ASAP7_75t_L g252 ( .A(n_34), .Y(n_252) );
INVx1_ASAP7_75t_L g486 ( .A(n_35), .Y(n_486) );
INVx2_ASAP7_75t_L g138 ( .A(n_36), .Y(n_138) );
CKINVDCx20_ASAP7_75t_R g189 ( .A(n_37), .Y(n_189) );
A2O1A1Ixp33_ASAP7_75t_L g207 ( .A1(n_38), .A2(n_149), .B(n_208), .C(n_210), .Y(n_207) );
INVxp67_ASAP7_75t_L g253 ( .A(n_39), .Y(n_253) );
CKINVDCx14_ASAP7_75t_R g206 ( .A(n_40), .Y(n_206) );
A2O1A1Ixp33_ASAP7_75t_L g227 ( .A1(n_41), .A2(n_145), .B(n_228), .C(n_234), .Y(n_227) );
A2O1A1Ixp33_ASAP7_75t_L g500 ( .A1(n_42), .A2(n_140), .B(n_145), .C(n_501), .Y(n_500) );
AOI22xp33_ASAP7_75t_L g117 ( .A1(n_43), .A2(n_118), .B1(n_119), .B2(n_426), .Y(n_117) );
CKINVDCx20_ASAP7_75t_R g426 ( .A(n_43), .Y(n_426) );
NAND2xp5_ASAP7_75t_L g104 ( .A(n_44), .B(n_105), .Y(n_104) );
INVx1_ASAP7_75t_L g485 ( .A(n_45), .Y(n_485) );
A2O1A1Ixp33_ASAP7_75t_L g166 ( .A1(n_46), .A2(n_167), .B(n_168), .C(n_171), .Y(n_166) );
NAND2xp5_ASAP7_75t_SL g511 ( .A(n_47), .B(n_150), .Y(n_511) );
CKINVDCx20_ASAP7_75t_R g236 ( .A(n_48), .Y(n_236) );
CKINVDCx20_ASAP7_75t_R g249 ( .A(n_49), .Y(n_249) );
INVx1_ASAP7_75t_L g143 ( .A(n_50), .Y(n_143) );
CKINVDCx16_ASAP7_75t_R g487 ( .A(n_51), .Y(n_487) );
NAND2xp5_ASAP7_75t_L g523 ( .A(n_52), .B(n_135), .Y(n_523) );
AOI22xp5_ASAP7_75t_L g483 ( .A1(n_53), .A2(n_145), .B1(n_155), .B2(n_484), .Y(n_483) );
CKINVDCx20_ASAP7_75t_R g505 ( .A(n_54), .Y(n_505) );
CKINVDCx16_ASAP7_75t_R g448 ( .A(n_55), .Y(n_448) );
CKINVDCx14_ASAP7_75t_R g165 ( .A(n_56), .Y(n_165) );
A2O1A1Ixp33_ASAP7_75t_L g471 ( .A1(n_57), .A2(n_167), .B(n_210), .C(n_472), .Y(n_471) );
CKINVDCx20_ASAP7_75t_R g514 ( .A(n_58), .Y(n_514) );
INVx1_ASAP7_75t_L g470 ( .A(n_59), .Y(n_470) );
INVx1_ASAP7_75t_L g141 ( .A(n_60), .Y(n_141) );
INVx1_ASAP7_75t_L g132 ( .A(n_61), .Y(n_132) );
INVx1_ASAP7_75t_SL g209 ( .A(n_62), .Y(n_209) );
CKINVDCx20_ASAP7_75t_R g115 ( .A(n_63), .Y(n_115) );
NAND2xp5_ASAP7_75t_L g158 ( .A(n_64), .B(n_159), .Y(n_158) );
INVx1_ASAP7_75t_L g218 ( .A(n_65), .Y(n_218) );
A2O1A1Ixp33_ASAP7_75t_SL g461 ( .A1(n_66), .A2(n_210), .B(n_462), .C(n_463), .Y(n_461) );
INVxp67_ASAP7_75t_L g464 ( .A(n_67), .Y(n_464) );
INVx1_ASAP7_75t_L g110 ( .A(n_68), .Y(n_110) );
AOI21xp5_ASAP7_75t_L g163 ( .A1(n_69), .A2(n_135), .B(n_164), .Y(n_163) );
CKINVDCx20_ASAP7_75t_R g222 ( .A(n_70), .Y(n_222) );
AOI21xp5_ASAP7_75t_L g191 ( .A1(n_71), .A2(n_135), .B(n_192), .Y(n_191) );
CKINVDCx20_ASAP7_75t_R g489 ( .A(n_72), .Y(n_489) );
INVx1_ASAP7_75t_L g508 ( .A(n_73), .Y(n_508) );
AOI21xp5_ASAP7_75t_L g246 ( .A1(n_74), .A2(n_247), .B(n_248), .Y(n_246) );
INVx1_ASAP7_75t_L g193 ( .A(n_75), .Y(n_193) );
CKINVDCx16_ASAP7_75t_R g226 ( .A(n_76), .Y(n_226) );
A2O1A1Ixp33_ASAP7_75t_L g509 ( .A1(n_77), .A2(n_140), .B(n_145), .C(n_510), .Y(n_509) );
AOI21xp5_ASAP7_75t_L g134 ( .A1(n_78), .A2(n_135), .B(n_142), .Y(n_134) );
INVx1_ASAP7_75t_L g196 ( .A(n_79), .Y(n_196) );
NAND2xp5_ASAP7_75t_SL g502 ( .A(n_80), .B(n_230), .Y(n_502) );
INVx2_ASAP7_75t_L g130 ( .A(n_81), .Y(n_130) );
INVx1_ASAP7_75t_L g183 ( .A(n_82), .Y(n_183) );
NAND2xp5_ASAP7_75t_L g503 ( .A(n_83), .B(n_462), .Y(n_503) );
A2O1A1Ixp33_ASAP7_75t_L g449 ( .A1(n_84), .A2(n_140), .B(n_145), .C(n_450), .Y(n_449) );
NAND3xp33_ASAP7_75t_SL g106 ( .A(n_85), .B(n_107), .C(n_108), .Y(n_106) );
OR2x2_ASAP7_75t_L g430 ( .A(n_85), .B(n_431), .Y(n_430) );
INVx2_ASAP7_75t_L g709 ( .A(n_85), .Y(n_709) );
OR2x2_ASAP7_75t_L g710 ( .A(n_85), .B(n_432), .Y(n_710) );
A2O1A1Ixp33_ASAP7_75t_L g216 ( .A1(n_86), .A2(n_145), .B(n_217), .C(n_220), .Y(n_216) );
NAND2xp5_ASAP7_75t_L g474 ( .A(n_87), .B(n_162), .Y(n_474) );
CKINVDCx20_ASAP7_75t_R g455 ( .A(n_88), .Y(n_455) );
A2O1A1Ixp33_ASAP7_75t_L g518 ( .A1(n_89), .A2(n_140), .B(n_145), .C(n_519), .Y(n_518) );
CKINVDCx20_ASAP7_75t_R g525 ( .A(n_90), .Y(n_525) );
INVx1_ASAP7_75t_L g460 ( .A(n_91), .Y(n_460) );
CKINVDCx16_ASAP7_75t_R g530 ( .A(n_92), .Y(n_530) );
NAND2xp5_ASAP7_75t_SL g520 ( .A(n_93), .B(n_230), .Y(n_520) );
NAND2xp5_ASAP7_75t_L g173 ( .A(n_94), .B(n_128), .Y(n_173) );
NAND2xp5_ASAP7_75t_L g534 ( .A(n_95), .B(n_128), .Y(n_534) );
NAND2xp5_ASAP7_75t_L g109 ( .A(n_96), .B(n_110), .Y(n_109) );
INVx2_ASAP7_75t_L g152 ( .A(n_97), .Y(n_152) );
AOI21xp5_ASAP7_75t_L g458 ( .A1(n_98), .A2(n_135), .B(n_459), .Y(n_458) );
CKINVDCx20_ASAP7_75t_R g100 ( .A(n_101), .Y(n_100) );
INVx5_ASAP7_75t_SL g101 ( .A(n_102), .Y(n_101) );
CKINVDCx9p33_ASAP7_75t_R g102 ( .A(n_103), .Y(n_102) );
BUFx2_ASAP7_75t_L g722 ( .A(n_103), .Y(n_722) );
OR2x4_ASAP7_75t_L g103 ( .A(n_104), .B(n_106), .Y(n_103) );
AND2x2_ASAP7_75t_L g432 ( .A(n_107), .B(n_433), .Y(n_432) );
INVx1_ASAP7_75t_SL g108 ( .A(n_109), .Y(n_108) );
AO21x2_ASAP7_75t_L g111 ( .A1(n_112), .A2(n_116), .B(n_437), .Y(n_111) );
HB1xp67_ASAP7_75t_L g112 ( .A(n_113), .Y(n_112) );
INVx2_ASAP7_75t_SL g113 ( .A(n_114), .Y(n_113) );
INVx2_ASAP7_75t_L g114 ( .A(n_115), .Y(n_114) );
INVx1_ASAP7_75t_L g721 ( .A(n_115), .Y(n_721) );
OAI21xp5_ASAP7_75t_SL g116 ( .A1(n_117), .A2(n_427), .B(n_434), .Y(n_116) );
INVx1_ASAP7_75t_L g118 ( .A(n_119), .Y(n_118) );
HB1xp67_ASAP7_75t_L g119 ( .A(n_120), .Y(n_119) );
OAI22xp5_ASAP7_75t_SL g439 ( .A1(n_120), .A2(n_440), .B1(n_708), .B2(n_710), .Y(n_439) );
INVx1_ASAP7_75t_L g120 ( .A(n_121), .Y(n_120) );
BUFx2_ASAP7_75t_L g715 ( .A(n_121), .Y(n_715) );
AND2x2_ASAP7_75t_L g121 ( .A(n_122), .B(n_352), .Y(n_121) );
NOR4xp25_ASAP7_75t_L g122 ( .A(n_123), .B(n_294), .C(n_324), .D(n_334), .Y(n_122) );
OAI211xp5_ASAP7_75t_L g123 ( .A1(n_124), .A2(n_199), .B(n_257), .C(n_284), .Y(n_123) );
OAI222xp33_ASAP7_75t_L g379 ( .A1(n_124), .A2(n_299), .B1(n_380), .B2(n_381), .C1(n_382), .C2(n_383), .Y(n_379) );
OR2x2_ASAP7_75t_L g124 ( .A(n_125), .B(n_174), .Y(n_124) );
AOI33xp33_ASAP7_75t_L g305 ( .A1(n_125), .A2(n_292), .A3(n_293), .B1(n_306), .B2(n_311), .B3(n_313), .Y(n_305) );
OAI211xp5_ASAP7_75t_SL g362 ( .A1(n_125), .A2(n_363), .B(n_365), .C(n_367), .Y(n_362) );
OR2x2_ASAP7_75t_L g378 ( .A(n_125), .B(n_364), .Y(n_378) );
INVx1_ASAP7_75t_L g411 ( .A(n_125), .Y(n_411) );
OR2x2_ASAP7_75t_L g125 ( .A(n_126), .B(n_161), .Y(n_125) );
INVx2_ASAP7_75t_L g288 ( .A(n_126), .Y(n_288) );
AND2x2_ASAP7_75t_L g304 ( .A(n_126), .B(n_190), .Y(n_304) );
HB1xp67_ASAP7_75t_L g339 ( .A(n_126), .Y(n_339) );
AND2x2_ASAP7_75t_L g368 ( .A(n_126), .B(n_161), .Y(n_368) );
OA21x2_ASAP7_75t_L g126 ( .A1(n_127), .A2(n_134), .B(n_158), .Y(n_126) );
OA21x2_ASAP7_75t_L g190 ( .A1(n_127), .A2(n_191), .B(n_198), .Y(n_190) );
OA21x2_ASAP7_75t_L g203 ( .A1(n_127), .A2(n_204), .B(n_212), .Y(n_203) );
HB1xp67_ASAP7_75t_L g127 ( .A(n_128), .Y(n_127) );
INVx4_ASAP7_75t_L g160 ( .A(n_128), .Y(n_160) );
OA21x2_ASAP7_75t_L g457 ( .A1(n_128), .A2(n_458), .B(n_465), .Y(n_457) );
BUFx6f_ASAP7_75t_L g128 ( .A(n_129), .Y(n_128) );
INVx1_ASAP7_75t_L g245 ( .A(n_129), .Y(n_245) );
AND2x2_ASAP7_75t_L g129 ( .A(n_130), .B(n_131), .Y(n_129) );
AND2x2_ASAP7_75t_SL g162 ( .A(n_130), .B(n_131), .Y(n_162) );
NAND2xp5_ASAP7_75t_L g131 ( .A(n_132), .B(n_133), .Y(n_131) );
BUFx2_ASAP7_75t_L g247 ( .A(n_135), .Y(n_247) );
AND2x4_ASAP7_75t_L g135 ( .A(n_136), .B(n_140), .Y(n_135) );
NAND2x1p5_ASAP7_75t_L g180 ( .A(n_136), .B(n_140), .Y(n_180) );
AND2x2_ASAP7_75t_L g136 ( .A(n_137), .B(n_139), .Y(n_136) );
INVx1_ASAP7_75t_L g233 ( .A(n_137), .Y(n_233) );
INVx1_ASAP7_75t_L g137 ( .A(n_138), .Y(n_137) );
INVx2_ASAP7_75t_L g146 ( .A(n_138), .Y(n_146) );
INVx1_ASAP7_75t_L g156 ( .A(n_138), .Y(n_156) );
INVx1_ASAP7_75t_L g147 ( .A(n_139), .Y(n_147) );
BUFx6f_ASAP7_75t_L g150 ( .A(n_139), .Y(n_150) );
BUFx6f_ASAP7_75t_L g154 ( .A(n_139), .Y(n_154) );
INVx3_ASAP7_75t_L g170 ( .A(n_139), .Y(n_170) );
INVx1_ASAP7_75t_L g462 ( .A(n_139), .Y(n_462) );
INVx4_ASAP7_75t_SL g157 ( .A(n_140), .Y(n_157) );
BUFx3_ASAP7_75t_L g234 ( .A(n_140), .Y(n_234) );
O2A1O1Ixp33_ASAP7_75t_SL g142 ( .A1(n_143), .A2(n_144), .B(n_148), .C(n_157), .Y(n_142) );
O2A1O1Ixp33_ASAP7_75t_SL g164 ( .A1(n_144), .A2(n_157), .B(n_165), .C(n_166), .Y(n_164) );
O2A1O1Ixp33_ASAP7_75t_SL g192 ( .A1(n_144), .A2(n_157), .B(n_193), .C(n_194), .Y(n_192) );
O2A1O1Ixp33_ASAP7_75t_L g205 ( .A1(n_144), .A2(n_157), .B(n_206), .C(n_207), .Y(n_205) );
O2A1O1Ixp33_ASAP7_75t_SL g248 ( .A1(n_144), .A2(n_157), .B(n_249), .C(n_250), .Y(n_248) );
O2A1O1Ixp33_ASAP7_75t_L g459 ( .A1(n_144), .A2(n_157), .B(n_460), .C(n_461), .Y(n_459) );
O2A1O1Ixp33_ASAP7_75t_L g469 ( .A1(n_144), .A2(n_157), .B(n_470), .C(n_471), .Y(n_469) );
O2A1O1Ixp33_ASAP7_75t_L g529 ( .A1(n_144), .A2(n_157), .B(n_530), .C(n_531), .Y(n_529) );
INVx5_ASAP7_75t_L g144 ( .A(n_145), .Y(n_144) );
AND2x6_ASAP7_75t_L g145 ( .A(n_146), .B(n_147), .Y(n_145) );
BUFx3_ASAP7_75t_L g172 ( .A(n_146), .Y(n_172) );
BUFx6f_ASAP7_75t_L g211 ( .A(n_146), .Y(n_211) );
NOR2xp33_ASAP7_75t_L g208 ( .A(n_149), .B(n_209), .Y(n_208) );
INVx4_ASAP7_75t_L g149 ( .A(n_150), .Y(n_149) );
INVx2_ASAP7_75t_L g167 ( .A(n_150), .Y(n_167) );
NOR2xp33_ASAP7_75t_L g151 ( .A(n_152), .B(n_153), .Y(n_151) );
NOR2xp33_ASAP7_75t_L g195 ( .A(n_153), .B(n_196), .Y(n_195) );
OAI22xp33_ASAP7_75t_L g251 ( .A1(n_153), .A2(n_230), .B1(n_252), .B2(n_253), .Y(n_251) );
NOR2xp33_ASAP7_75t_L g532 ( .A(n_153), .B(n_533), .Y(n_532) );
INVx4_ASAP7_75t_L g153 ( .A(n_154), .Y(n_153) );
INVx2_ASAP7_75t_L g185 ( .A(n_154), .Y(n_185) );
OAI22xp5_ASAP7_75t_SL g484 ( .A1(n_154), .A2(n_185), .B1(n_485), .B2(n_486), .Y(n_484) );
INVx2_ASAP7_75t_L g453 ( .A(n_155), .Y(n_453) );
INVx3_ASAP7_75t_L g155 ( .A(n_156), .Y(n_155) );
INVx1_ASAP7_75t_L g220 ( .A(n_157), .Y(n_220) );
OAI22xp33_ASAP7_75t_L g482 ( .A1(n_157), .A2(n_180), .B1(n_483), .B2(n_487), .Y(n_482) );
OA21x2_ASAP7_75t_L g467 ( .A1(n_159), .A2(n_468), .B(n_474), .Y(n_467) );
INVx3_ASAP7_75t_L g159 ( .A(n_160), .Y(n_159) );
NOR2xp33_ASAP7_75t_L g188 ( .A(n_160), .B(n_189), .Y(n_188) );
AO21x2_ASAP7_75t_L g213 ( .A1(n_160), .A2(n_214), .B(n_221), .Y(n_213) );
NOR2xp33_ASAP7_75t_L g235 ( .A(n_160), .B(n_236), .Y(n_235) );
NOR2xp33_ASAP7_75t_SL g504 ( .A(n_160), .B(n_505), .Y(n_504) );
INVx2_ASAP7_75t_L g268 ( .A(n_161), .Y(n_268) );
BUFx3_ASAP7_75t_L g276 ( .A(n_161), .Y(n_276) );
NAND2xp5_ASAP7_75t_L g278 ( .A(n_161), .B(n_279), .Y(n_278) );
AND2x2_ASAP7_75t_L g287 ( .A(n_161), .B(n_288), .Y(n_287) );
NOR2xp33_ASAP7_75t_L g316 ( .A(n_161), .B(n_175), .Y(n_316) );
AND2x2_ASAP7_75t_L g385 ( .A(n_161), .B(n_319), .Y(n_385) );
OA21x2_ASAP7_75t_L g161 ( .A1(n_162), .A2(n_163), .B(n_173), .Y(n_161) );
INVx1_ASAP7_75t_L g177 ( .A(n_162), .Y(n_177) );
INVx2_ASAP7_75t_L g223 ( .A(n_162), .Y(n_223) );
O2A1O1Ixp33_ASAP7_75t_L g225 ( .A1(n_162), .A2(n_180), .B(n_226), .C(n_227), .Y(n_225) );
OA21x2_ASAP7_75t_L g527 ( .A1(n_162), .A2(n_528), .B(n_534), .Y(n_527) );
NOR2xp33_ASAP7_75t_L g168 ( .A(n_169), .B(n_170), .Y(n_168) );
INVx5_ASAP7_75t_L g230 ( .A(n_170), .Y(n_230) );
NOR2xp33_ASAP7_75t_L g463 ( .A(n_170), .B(n_464), .Y(n_463) );
NOR2xp33_ASAP7_75t_L g472 ( .A(n_170), .B(n_473), .Y(n_472) );
INVx2_ASAP7_75t_L g187 ( .A(n_171), .Y(n_187) );
INVx2_ASAP7_75t_L g171 ( .A(n_172), .Y(n_171) );
INVx1_ASAP7_75t_L g197 ( .A(n_172), .Y(n_197) );
INVx2_ASAP7_75t_SL g279 ( .A(n_174), .Y(n_279) );
OR2x2_ASAP7_75t_L g174 ( .A(n_175), .B(n_190), .Y(n_174) );
NAND2xp5_ASAP7_75t_L g267 ( .A(n_175), .B(n_268), .Y(n_267) );
INVx1_ASAP7_75t_L g321 ( .A(n_175), .Y(n_321) );
AND2x2_ASAP7_75t_L g332 ( .A(n_175), .B(n_288), .Y(n_332) );
NAND2xp5_ASAP7_75t_L g348 ( .A(n_175), .B(n_317), .Y(n_348) );
NAND2xp5_ASAP7_75t_L g364 ( .A(n_175), .B(n_319), .Y(n_364) );
AND2x2_ASAP7_75t_L g423 ( .A(n_175), .B(n_368), .Y(n_423) );
INVx4_ASAP7_75t_L g175 ( .A(n_176), .Y(n_175) );
AND2x2_ASAP7_75t_L g293 ( .A(n_176), .B(n_190), .Y(n_293) );
AND2x2_ASAP7_75t_L g303 ( .A(n_176), .B(n_304), .Y(n_303) );
BUFx3_ASAP7_75t_L g325 ( .A(n_176), .Y(n_325) );
AND3x2_ASAP7_75t_L g384 ( .A(n_176), .B(n_385), .C(n_386), .Y(n_384) );
AO21x2_ASAP7_75t_L g176 ( .A1(n_177), .A2(n_178), .B(n_188), .Y(n_176) );
NOR2xp33_ASAP7_75t_L g454 ( .A(n_177), .B(n_455), .Y(n_454) );
NOR2xp33_ASAP7_75t_L g513 ( .A(n_177), .B(n_514), .Y(n_513) );
NOR2xp33_ASAP7_75t_L g524 ( .A(n_177), .B(n_525), .Y(n_524) );
OAI21xp5_ASAP7_75t_L g178 ( .A1(n_179), .A2(n_180), .B(n_181), .Y(n_178) );
OAI21xp5_ASAP7_75t_L g214 ( .A1(n_180), .A2(n_215), .B(n_216), .Y(n_214) );
OAI21xp5_ASAP7_75t_L g447 ( .A1(n_180), .A2(n_448), .B(n_449), .Y(n_447) );
OAI21xp5_ASAP7_75t_L g507 ( .A1(n_180), .A2(n_508), .B(n_509), .Y(n_507) );
O2A1O1Ixp5_ASAP7_75t_L g182 ( .A1(n_183), .A2(n_184), .B(n_186), .C(n_187), .Y(n_182) );
O2A1O1Ixp33_ASAP7_75t_L g217 ( .A1(n_184), .A2(n_187), .B(n_218), .C(n_219), .Y(n_217) );
INVx2_ASAP7_75t_L g184 ( .A(n_185), .Y(n_184) );
AOI21xp5_ASAP7_75t_L g501 ( .A1(n_187), .A2(n_502), .B(n_503), .Y(n_501) );
AOI21xp5_ASAP7_75t_L g510 ( .A1(n_187), .A2(n_511), .B(n_512), .Y(n_510) );
HB1xp67_ASAP7_75t_L g275 ( .A(n_190), .Y(n_275) );
INVx1_ASAP7_75t_SL g319 ( .A(n_190), .Y(n_319) );
NAND3xp33_ASAP7_75t_L g331 ( .A(n_190), .B(n_268), .C(n_332), .Y(n_331) );
NOR2xp33_ASAP7_75t_L g199 ( .A(n_200), .B(n_237), .Y(n_199) );
A2O1A1Ixp33_ASAP7_75t_L g354 ( .A1(n_200), .A2(n_303), .B(n_355), .C(n_357), .Y(n_354) );
INVx1_ASAP7_75t_L g200 ( .A(n_201), .Y(n_200) );
NAND2xp5_ASAP7_75t_SL g201 ( .A(n_202), .B(n_224), .Y(n_201) );
NAND2xp5_ASAP7_75t_L g360 ( .A(n_202), .B(n_361), .Y(n_360) );
INVx2_ASAP7_75t_SL g371 ( .A(n_202), .Y(n_371) );
AND2x2_ASAP7_75t_L g392 ( .A(n_202), .B(n_239), .Y(n_392) );
NOR2xp33_ASAP7_75t_L g420 ( .A(n_202), .B(n_301), .Y(n_420) );
AND2x2_ASAP7_75t_L g202 ( .A(n_203), .B(n_213), .Y(n_202) );
AND2x2_ASAP7_75t_L g265 ( .A(n_203), .B(n_256), .Y(n_265) );
INVx2_ASAP7_75t_L g272 ( .A(n_203), .Y(n_272) );
AND2x2_ASAP7_75t_L g292 ( .A(n_203), .B(n_239), .Y(n_292) );
AND2x2_ASAP7_75t_L g342 ( .A(n_203), .B(n_224), .Y(n_342) );
INVx1_ASAP7_75t_L g346 ( .A(n_203), .Y(n_346) );
INVx3_ASAP7_75t_L g210 ( .A(n_211), .Y(n_210) );
HB1xp67_ASAP7_75t_L g522 ( .A(n_211), .Y(n_522) );
INVx2_ASAP7_75t_SL g256 ( .A(n_213), .Y(n_256) );
BUFx2_ASAP7_75t_L g282 ( .A(n_213), .Y(n_282) );
AND2x2_ASAP7_75t_L g409 ( .A(n_213), .B(n_224), .Y(n_409) );
NOR2xp33_ASAP7_75t_L g221 ( .A(n_222), .B(n_223), .Y(n_221) );
INVx1_ASAP7_75t_L g255 ( .A(n_223), .Y(n_255) );
AO21x2_ASAP7_75t_L g516 ( .A1(n_223), .A2(n_517), .B(n_524), .Y(n_516) );
INVx3_ASAP7_75t_SL g239 ( .A(n_224), .Y(n_239) );
AND2x2_ASAP7_75t_L g264 ( .A(n_224), .B(n_265), .Y(n_264) );
AND2x4_ASAP7_75t_L g271 ( .A(n_224), .B(n_272), .Y(n_271) );
OR2x2_ASAP7_75t_L g301 ( .A(n_224), .B(n_261), .Y(n_301) );
OR2x2_ASAP7_75t_L g310 ( .A(n_224), .B(n_256), .Y(n_310) );
HB1xp67_ASAP7_75t_L g328 ( .A(n_224), .Y(n_328) );
AND2x2_ASAP7_75t_L g333 ( .A(n_224), .B(n_286), .Y(n_333) );
AND2x2_ASAP7_75t_L g361 ( .A(n_224), .B(n_241), .Y(n_361) );
NAND2xp5_ASAP7_75t_L g396 ( .A(n_224), .B(n_397), .Y(n_396) );
OR2x2_ASAP7_75t_L g399 ( .A(n_224), .B(n_240), .Y(n_399) );
OR2x6_ASAP7_75t_L g224 ( .A(n_225), .B(n_235), .Y(n_224) );
O2A1O1Ixp33_ASAP7_75t_L g228 ( .A1(n_229), .A2(n_230), .B(n_231), .C(n_232), .Y(n_228) );
O2A1O1Ixp33_ASAP7_75t_L g450 ( .A1(n_230), .A2(n_451), .B(n_452), .C(n_453), .Y(n_450) );
INVx2_ASAP7_75t_L g232 ( .A(n_233), .Y(n_232) );
NAND2xp5_ASAP7_75t_SL g250 ( .A(n_233), .B(n_251), .Y(n_250) );
INVx1_ASAP7_75t_L g237 ( .A(n_238), .Y(n_237) );
OR2x2_ASAP7_75t_L g238 ( .A(n_239), .B(n_240), .Y(n_238) );
AND2x2_ASAP7_75t_L g323 ( .A(n_239), .B(n_272), .Y(n_323) );
NAND2xp5_ASAP7_75t_L g351 ( .A(n_239), .B(n_265), .Y(n_351) );
AND2x2_ASAP7_75t_L g369 ( .A(n_239), .B(n_286), .Y(n_369) );
OR2x2_ASAP7_75t_L g240 ( .A(n_241), .B(n_256), .Y(n_240) );
AND2x2_ASAP7_75t_L g270 ( .A(n_241), .B(n_256), .Y(n_270) );
NAND2xp5_ASAP7_75t_L g298 ( .A(n_241), .B(n_299), .Y(n_298) );
BUFx3_ASAP7_75t_L g308 ( .A(n_241), .Y(n_308) );
OR2x2_ASAP7_75t_L g356 ( .A(n_241), .B(n_276), .Y(n_356) );
OA21x2_ASAP7_75t_L g241 ( .A1(n_242), .A2(n_246), .B(n_254), .Y(n_241) );
INVx1_ASAP7_75t_L g242 ( .A(n_243), .Y(n_242) );
AO21x2_ASAP7_75t_L g261 ( .A1(n_243), .A2(n_262), .B(n_263), .Y(n_261) );
AO21x2_ASAP7_75t_L g506 ( .A1(n_243), .A2(n_507), .B(n_513), .Y(n_506) );
INVx1_ASAP7_75t_L g243 ( .A(n_244), .Y(n_243) );
AOI21xp5_ASAP7_75t_SL g498 ( .A1(n_244), .A2(n_499), .B(n_500), .Y(n_498) );
INVx2_ASAP7_75t_L g244 ( .A(n_245), .Y(n_244) );
AO21x2_ASAP7_75t_L g446 ( .A1(n_245), .A2(n_447), .B(n_454), .Y(n_446) );
AO21x2_ASAP7_75t_L g481 ( .A1(n_245), .A2(n_482), .B(n_488), .Y(n_481) );
NOR2xp33_ASAP7_75t_L g488 ( .A(n_245), .B(n_489), .Y(n_488) );
INVx1_ASAP7_75t_L g262 ( .A(n_246), .Y(n_262) );
INVx1_ASAP7_75t_L g263 ( .A(n_254), .Y(n_263) );
AND2x2_ASAP7_75t_L g291 ( .A(n_256), .B(n_261), .Y(n_291) );
INVx1_ASAP7_75t_L g299 ( .A(n_256), .Y(n_299) );
AND2x2_ASAP7_75t_L g394 ( .A(n_256), .B(n_272), .Y(n_394) );
AOI222xp33_ASAP7_75t_L g257 ( .A1(n_258), .A2(n_266), .B1(n_269), .B2(n_273), .C1(n_277), .C2(n_280), .Y(n_257) );
INVx1_ASAP7_75t_L g389 ( .A(n_258), .Y(n_389) );
AND2x2_ASAP7_75t_L g258 ( .A(n_259), .B(n_264), .Y(n_258) );
AND2x2_ASAP7_75t_L g285 ( .A(n_259), .B(n_286), .Y(n_285) );
AND2x2_ASAP7_75t_L g296 ( .A(n_259), .B(n_265), .Y(n_296) );
NAND2xp5_ASAP7_75t_L g312 ( .A(n_259), .B(n_287), .Y(n_312) );
OAI222xp33_ASAP7_75t_L g334 ( .A1(n_259), .A2(n_335), .B1(n_340), .B2(n_341), .C1(n_349), .C2(n_351), .Y(n_334) );
INVx2_ASAP7_75t_L g259 ( .A(n_260), .Y(n_259) );
INVx1_ASAP7_75t_SL g260 ( .A(n_261), .Y(n_260) );
AND2x2_ASAP7_75t_L g322 ( .A(n_261), .B(n_323), .Y(n_322) );
NAND2xp5_ASAP7_75t_L g382 ( .A(n_261), .B(n_342), .Y(n_382) );
AND2x2_ASAP7_75t_L g393 ( .A(n_261), .B(n_394), .Y(n_393) );
INVx1_ASAP7_75t_L g401 ( .A(n_264), .Y(n_401) );
NAND2xp5_ASAP7_75t_SL g380 ( .A(n_266), .B(n_317), .Y(n_380) );
INVx1_ASAP7_75t_L g266 ( .A(n_267), .Y(n_266) );
NOR2xp33_ASAP7_75t_L g320 ( .A(n_268), .B(n_321), .Y(n_320) );
AND2x2_ASAP7_75t_L g338 ( .A(n_268), .B(n_339), .Y(n_338) );
AND2x2_ASAP7_75t_L g269 ( .A(n_270), .B(n_271), .Y(n_269) );
INVx3_ASAP7_75t_L g283 ( .A(n_271), .Y(n_283) );
O2A1O1Ixp33_ASAP7_75t_L g373 ( .A1(n_271), .A2(n_374), .B(n_377), .C(n_379), .Y(n_373) );
NAND2xp5_ASAP7_75t_L g388 ( .A(n_271), .B(n_308), .Y(n_388) );
NAND2xp5_ASAP7_75t_L g413 ( .A(n_271), .B(n_291), .Y(n_413) );
AND2x2_ASAP7_75t_L g286 ( .A(n_272), .B(n_282), .Y(n_286) );
INVx1_ASAP7_75t_L g273 ( .A(n_274), .Y(n_273) );
NAND2xp5_ASAP7_75t_L g274 ( .A(n_275), .B(n_276), .Y(n_274) );
INVx1_ASAP7_75t_L g313 ( .A(n_275), .Y(n_313) );
NAND2xp5_ASAP7_75t_SL g302 ( .A(n_276), .B(n_303), .Y(n_302) );
OR2x2_ASAP7_75t_L g365 ( .A(n_276), .B(n_366), .Y(n_365) );
AND2x2_ASAP7_75t_L g404 ( .A(n_276), .B(n_304), .Y(n_404) );
INVx1_ASAP7_75t_L g416 ( .A(n_276), .Y(n_416) );
INVx1_ASAP7_75t_L g277 ( .A(n_278), .Y(n_277) );
NAND2xp5_ASAP7_75t_L g417 ( .A(n_279), .B(n_418), .Y(n_417) );
INVx1_ASAP7_75t_L g280 ( .A(n_281), .Y(n_280) );
OR2x2_ASAP7_75t_L g281 ( .A(n_282), .B(n_283), .Y(n_281) );
INVx1_ASAP7_75t_L g397 ( .A(n_282), .Y(n_397) );
A2O1A1Ixp33_ASAP7_75t_SL g284 ( .A1(n_285), .A2(n_287), .B(n_289), .C(n_293), .Y(n_284) );
AOI22xp33_ASAP7_75t_L g329 ( .A1(n_285), .A2(n_315), .B1(n_330), .B2(n_333), .Y(n_329) );
NAND2xp5_ASAP7_75t_L g340 ( .A(n_286), .B(n_300), .Y(n_340) );
NAND2xp5_ASAP7_75t_L g425 ( .A(n_286), .B(n_308), .Y(n_425) );
NAND2xp5_ASAP7_75t_L g344 ( .A(n_287), .B(n_345), .Y(n_344) );
INVx1_ASAP7_75t_SL g350 ( .A(n_287), .Y(n_350) );
AND2x2_ASAP7_75t_L g357 ( .A(n_287), .B(n_337), .Y(n_357) );
INVx2_ASAP7_75t_L g318 ( .A(n_288), .Y(n_318) );
INVxp67_ASAP7_75t_L g289 ( .A(n_290), .Y(n_289) );
NAND2xp5_ASAP7_75t_L g290 ( .A(n_291), .B(n_292), .Y(n_290) );
NOR4xp25_ASAP7_75t_L g295 ( .A(n_292), .B(n_296), .C(n_297), .D(n_300), .Y(n_295) );
INVx1_ASAP7_75t_SL g366 ( .A(n_293), .Y(n_366) );
AND2x2_ASAP7_75t_L g410 ( .A(n_293), .B(n_411), .Y(n_410) );
OAI211xp5_ASAP7_75t_SL g294 ( .A1(n_295), .A2(n_302), .B(n_305), .C(n_314), .Y(n_294) );
INVx1_ASAP7_75t_L g297 ( .A(n_298), .Y(n_297) );
INVx1_ASAP7_75t_SL g300 ( .A(n_301), .Y(n_300) );
NOR2xp33_ASAP7_75t_L g422 ( .A(n_301), .B(n_371), .Y(n_422) );
AOI22xp5_ASAP7_75t_L g421 ( .A1(n_303), .A2(n_422), .B1(n_423), .B2(n_424), .Y(n_421) );
INVx1_ASAP7_75t_SL g376 ( .A(n_304), .Y(n_376) );
AND2x2_ASAP7_75t_L g415 ( .A(n_304), .B(n_416), .Y(n_415) );
INVx1_ASAP7_75t_L g306 ( .A(n_307), .Y(n_306) );
NAND2xp5_ASAP7_75t_L g307 ( .A(n_308), .B(n_309), .Y(n_307) );
NAND2xp5_ASAP7_75t_SL g408 ( .A(n_308), .B(n_409), .Y(n_408) );
INVx1_ASAP7_75t_L g309 ( .A(n_310), .Y(n_309) );
INVx1_ASAP7_75t_L g311 ( .A(n_312), .Y(n_311) );
NOR2xp33_ASAP7_75t_L g327 ( .A(n_312), .B(n_328), .Y(n_327) );
NAND2xp5_ASAP7_75t_L g398 ( .A(n_313), .B(n_338), .Y(n_398) );
OAI21xp5_ASAP7_75t_SL g314 ( .A1(n_315), .A2(n_320), .B(n_322), .Y(n_314) );
AND2x2_ASAP7_75t_L g315 ( .A(n_316), .B(n_317), .Y(n_315) );
INVx1_ASAP7_75t_L g390 ( .A(n_317), .Y(n_390) );
AND2x2_ASAP7_75t_L g317 ( .A(n_318), .B(n_319), .Y(n_317) );
INVx2_ASAP7_75t_L g418 ( .A(n_318), .Y(n_418) );
HB1xp67_ASAP7_75t_L g345 ( .A(n_319), .Y(n_345) );
OAI21xp33_ASAP7_75t_L g324 ( .A1(n_325), .A2(n_326), .B(n_329), .Y(n_324) );
CKINVDCx16_ASAP7_75t_R g337 ( .A(n_325), .Y(n_337) );
OR2x2_ASAP7_75t_L g375 ( .A(n_325), .B(n_376), .Y(n_375) );
INVx1_ASAP7_75t_L g326 ( .A(n_327), .Y(n_326) );
AOI21xp33_ASAP7_75t_SL g370 ( .A1(n_328), .A2(n_371), .B(n_372), .Y(n_370) );
INVx1_ASAP7_75t_L g330 ( .A(n_331), .Y(n_330) );
AOI221xp5_ASAP7_75t_L g358 ( .A1(n_332), .A2(n_359), .B1(n_362), .B2(n_369), .C(n_370), .Y(n_358) );
INVx1_ASAP7_75t_SL g402 ( .A(n_333), .Y(n_402) );
INVx1_ASAP7_75t_L g335 ( .A(n_336), .Y(n_335) );
AND2x2_ASAP7_75t_L g336 ( .A(n_337), .B(n_338), .Y(n_336) );
OR2x2_ASAP7_75t_L g349 ( .A(n_337), .B(n_350), .Y(n_349) );
INVxp67_ASAP7_75t_L g386 ( .A(n_339), .Y(n_386) );
AOI22xp5_ASAP7_75t_L g341 ( .A1(n_342), .A2(n_343), .B1(n_346), .B2(n_347), .Y(n_341) );
INVx1_ASAP7_75t_L g381 ( .A(n_342), .Y(n_381) );
INVxp67_ASAP7_75t_L g343 ( .A(n_344), .Y(n_343) );
NAND2xp5_ASAP7_75t_L g367 ( .A(n_345), .B(n_368), .Y(n_367) );
INVx1_ASAP7_75t_L g347 ( .A(n_348), .Y(n_347) );
NOR4xp25_ASAP7_75t_L g352 ( .A(n_353), .B(n_387), .C(n_400), .D(n_412), .Y(n_352) );
NAND3xp33_ASAP7_75t_SL g353 ( .A(n_354), .B(n_358), .C(n_373), .Y(n_353) );
INVx1_ASAP7_75t_L g355 ( .A(n_356), .Y(n_355) );
NOR2xp33_ASAP7_75t_L g374 ( .A(n_356), .B(n_375), .Y(n_374) );
INVx1_ASAP7_75t_L g359 ( .A(n_360), .Y(n_359) );
NAND2xp5_ASAP7_75t_L g372 ( .A(n_363), .B(n_368), .Y(n_372) );
INVx1_ASAP7_75t_L g363 ( .A(n_364), .Y(n_363) );
OAI221xp5_ASAP7_75t_SL g400 ( .A1(n_375), .A2(n_401), .B1(n_402), .B2(n_403), .C(n_405), .Y(n_400) );
O2A1O1Ixp33_ASAP7_75t_L g391 ( .A1(n_377), .A2(n_392), .B(n_393), .C(n_395), .Y(n_391) );
INVx2_ASAP7_75t_L g377 ( .A(n_378), .Y(n_377) );
OAI22xp5_ASAP7_75t_L g395 ( .A1(n_378), .A2(n_396), .B1(n_398), .B2(n_399), .Y(n_395) );
INVx2_ASAP7_75t_SL g383 ( .A(n_384), .Y(n_383) );
A2O1A1Ixp33_ASAP7_75t_L g387 ( .A1(n_388), .A2(n_389), .B(n_390), .C(n_391), .Y(n_387) );
INVx1_ASAP7_75t_L g406 ( .A(n_399), .Y(n_406) );
INVx1_ASAP7_75t_L g403 ( .A(n_404), .Y(n_403) );
OAI21xp5_ASAP7_75t_SL g405 ( .A1(n_406), .A2(n_407), .B(n_410), .Y(n_405) );
INVx1_ASAP7_75t_L g407 ( .A(n_408), .Y(n_407) );
OAI221xp5_ASAP7_75t_SL g412 ( .A1(n_413), .A2(n_414), .B1(n_417), .B2(n_419), .C(n_421), .Y(n_412) );
INVx1_ASAP7_75t_L g414 ( .A(n_415), .Y(n_414) );
INVxp67_ASAP7_75t_L g419 ( .A(n_420), .Y(n_419) );
INVx1_ASAP7_75t_L g424 ( .A(n_425), .Y(n_424) );
INVx1_ASAP7_75t_L g427 ( .A(n_428), .Y(n_427) );
INVx1_ASAP7_75t_SL g428 ( .A(n_429), .Y(n_428) );
INVx1_ASAP7_75t_SL g429 ( .A(n_430), .Y(n_429) );
HB1xp67_ASAP7_75t_L g436 ( .A(n_430), .Y(n_436) );
NOR2x2_ASAP7_75t_L g719 ( .A(n_431), .B(n_709), .Y(n_719) );
INVx2_ASAP7_75t_L g431 ( .A(n_432), .Y(n_431) );
OR2x2_ASAP7_75t_L g708 ( .A(n_432), .B(n_709), .Y(n_708) );
AOI21xp33_ASAP7_75t_L g437 ( .A1(n_434), .A2(n_438), .B(n_720), .Y(n_437) );
INVx1_ASAP7_75t_L g435 ( .A(n_436), .Y(n_435) );
INVx1_ASAP7_75t_L g712 ( .A(n_440), .Y(n_712) );
NAND2x1_ASAP7_75t_L g440 ( .A(n_441), .B(n_624), .Y(n_440) );
NOR5xp2_ASAP7_75t_L g441 ( .A(n_442), .B(n_547), .C(n_579), .D(n_594), .E(n_611), .Y(n_441) );
A2O1A1Ixp33_ASAP7_75t_L g442 ( .A1(n_443), .A2(n_475), .B(n_494), .C(n_535), .Y(n_442) );
NAND2xp5_ASAP7_75t_L g443 ( .A(n_444), .B(n_456), .Y(n_443) );
NAND2xp5_ASAP7_75t_L g646 ( .A(n_444), .B(n_647), .Y(n_646) );
NAND2xp5_ASAP7_75t_L g662 ( .A(n_444), .B(n_599), .Y(n_662) );
INVx1_ASAP7_75t_L g444 ( .A(n_445), .Y(n_444) );
NAND2xp5_ASAP7_75t_L g543 ( .A(n_445), .B(n_544), .Y(n_543) );
NAND2xp5_ASAP7_75t_L g548 ( .A(n_445), .B(n_491), .Y(n_548) );
AND2x2_ASAP7_75t_L g589 ( .A(n_445), .B(n_590), .Y(n_589) );
NAND2xp5_ASAP7_75t_L g593 ( .A(n_445), .B(n_558), .Y(n_593) );
OR2x2_ASAP7_75t_L g630 ( .A(n_445), .B(n_481), .Y(n_630) );
INVx3_ASAP7_75t_L g445 ( .A(n_446), .Y(n_445) );
AND2x2_ASAP7_75t_L g480 ( .A(n_446), .B(n_481), .Y(n_480) );
INVx3_ASAP7_75t_L g538 ( .A(n_446), .Y(n_538) );
OR2x2_ASAP7_75t_L g701 ( .A(n_446), .B(n_541), .Y(n_701) );
AOI22xp5_ASAP7_75t_L g603 ( .A1(n_456), .A2(n_604), .B1(n_605), .B2(n_608), .Y(n_603) );
NAND2xp5_ASAP7_75t_L g687 ( .A(n_456), .B(n_538), .Y(n_687) );
AND2x2_ASAP7_75t_L g456 ( .A(n_457), .B(n_466), .Y(n_456) );
AND2x2_ASAP7_75t_L g493 ( .A(n_457), .B(n_481), .Y(n_493) );
AND2x2_ASAP7_75t_L g540 ( .A(n_457), .B(n_541), .Y(n_540) );
INVx1_ASAP7_75t_L g545 ( .A(n_457), .Y(n_545) );
INVx3_ASAP7_75t_L g558 ( .A(n_457), .Y(n_558) );
OR2x2_ASAP7_75t_L g578 ( .A(n_457), .B(n_541), .Y(n_578) );
AND2x2_ASAP7_75t_L g597 ( .A(n_457), .B(n_467), .Y(n_597) );
BUFx2_ASAP7_75t_L g629 ( .A(n_457), .Y(n_629) );
AND2x4_ASAP7_75t_L g544 ( .A(n_466), .B(n_545), .Y(n_544) );
INVx1_ASAP7_75t_SL g466 ( .A(n_467), .Y(n_466) );
BUFx2_ASAP7_75t_L g479 ( .A(n_467), .Y(n_479) );
INVx2_ASAP7_75t_L g492 ( .A(n_467), .Y(n_492) );
OR2x2_ASAP7_75t_L g560 ( .A(n_467), .B(n_541), .Y(n_560) );
AND2x2_ASAP7_75t_L g590 ( .A(n_467), .B(n_481), .Y(n_590) );
AND2x2_ASAP7_75t_L g607 ( .A(n_467), .B(n_538), .Y(n_607) );
AND2x2_ASAP7_75t_L g647 ( .A(n_467), .B(n_558), .Y(n_647) );
AND2x2_ASAP7_75t_SL g683 ( .A(n_467), .B(n_493), .Y(n_683) );
INVx1_ASAP7_75t_L g475 ( .A(n_476), .Y(n_475) );
NAND2xp33_ASAP7_75t_SL g476 ( .A(n_477), .B(n_490), .Y(n_476) );
NAND2xp5_ASAP7_75t_L g477 ( .A(n_478), .B(n_480), .Y(n_477) );
NOR2xp33_ASAP7_75t_L g661 ( .A(n_478), .B(n_662), .Y(n_661) );
INVx1_ASAP7_75t_SL g478 ( .A(n_479), .Y(n_478) );
OAI21xp33_ASAP7_75t_L g621 ( .A1(n_479), .A2(n_493), .B(n_622), .Y(n_621) );
NOR2xp33_ASAP7_75t_L g677 ( .A(n_479), .B(n_481), .Y(n_677) );
AND2x2_ASAP7_75t_L g613 ( .A(n_480), .B(n_614), .Y(n_613) );
INVx3_ASAP7_75t_L g541 ( .A(n_481), .Y(n_541) );
HB1xp67_ASAP7_75t_L g639 ( .A(n_481), .Y(n_639) );
NOR2xp33_ASAP7_75t_L g706 ( .A(n_490), .B(n_538), .Y(n_706) );
INVx2_ASAP7_75t_L g490 ( .A(n_491), .Y(n_490) );
AOI22xp33_ASAP7_75t_L g648 ( .A1(n_491), .A2(n_649), .B1(n_650), .B2(n_655), .Y(n_648) );
AND2x2_ASAP7_75t_L g491 ( .A(n_492), .B(n_493), .Y(n_491) );
AND2x2_ASAP7_75t_L g539 ( .A(n_492), .B(n_540), .Y(n_539) );
OR2x2_ASAP7_75t_L g577 ( .A(n_492), .B(n_578), .Y(n_577) );
INVx1_ASAP7_75t_SL g614 ( .A(n_492), .Y(n_614) );
NAND2xp5_ASAP7_75t_L g606 ( .A(n_493), .B(n_607), .Y(n_606) );
INVx1_ASAP7_75t_L g668 ( .A(n_493), .Y(n_668) );
CKINVDCx16_ASAP7_75t_R g494 ( .A(n_495), .Y(n_494) );
AND2x2_ASAP7_75t_L g495 ( .A(n_496), .B(n_515), .Y(n_495) );
INVx4_ASAP7_75t_L g554 ( .A(n_496), .Y(n_554) );
AND2x2_ASAP7_75t_L g632 ( .A(n_496), .B(n_599), .Y(n_632) );
AND2x2_ASAP7_75t_L g496 ( .A(n_497), .B(n_506), .Y(n_496) );
INVx3_ASAP7_75t_L g551 ( .A(n_497), .Y(n_551) );
AND2x2_ASAP7_75t_L g565 ( .A(n_497), .B(n_566), .Y(n_565) );
INVx1_ASAP7_75t_L g569 ( .A(n_497), .Y(n_569) );
INVx2_ASAP7_75t_L g583 ( .A(n_497), .Y(n_583) );
NAND2xp5_ASAP7_75t_L g598 ( .A(n_497), .B(n_599), .Y(n_598) );
AND2x2_ASAP7_75t_L g640 ( .A(n_497), .B(n_635), .Y(n_640) );
AND2x2_ASAP7_75t_L g705 ( .A(n_497), .B(n_675), .Y(n_705) );
OR2x6_ASAP7_75t_L g497 ( .A(n_498), .B(n_504), .Y(n_497) );
AND2x2_ASAP7_75t_L g546 ( .A(n_506), .B(n_527), .Y(n_546) );
INVx2_ASAP7_75t_L g566 ( .A(n_506), .Y(n_566) );
INVx1_ASAP7_75t_L g571 ( .A(n_515), .Y(n_571) );
AND2x2_ASAP7_75t_L g617 ( .A(n_515), .B(n_565), .Y(n_617) );
AND2x2_ASAP7_75t_L g515 ( .A(n_516), .B(n_526), .Y(n_515) );
INVx2_ASAP7_75t_L g556 ( .A(n_516), .Y(n_556) );
INVx1_ASAP7_75t_L g564 ( .A(n_516), .Y(n_564) );
AND2x2_ASAP7_75t_L g582 ( .A(n_516), .B(n_583), .Y(n_582) );
NAND2xp5_ASAP7_75t_L g620 ( .A(n_516), .B(n_566), .Y(n_620) );
NAND2xp5_ASAP7_75t_L g517 ( .A(n_518), .B(n_523), .Y(n_517) );
AOI21xp5_ASAP7_75t_L g519 ( .A1(n_520), .A2(n_521), .B(n_522), .Y(n_519) );
AND2x2_ASAP7_75t_L g599 ( .A(n_526), .B(n_556), .Y(n_599) );
INVx1_ASAP7_75t_L g526 ( .A(n_527), .Y(n_526) );
INVx2_ASAP7_75t_L g552 ( .A(n_527), .Y(n_552) );
AND2x2_ASAP7_75t_L g635 ( .A(n_527), .B(n_566), .Y(n_635) );
OAI21xp5_ASAP7_75t_SL g535 ( .A1(n_536), .A2(n_542), .B(n_546), .Y(n_535) );
INVx1_ASAP7_75t_SL g580 ( .A(n_536), .Y(n_580) );
AND2x2_ASAP7_75t_L g536 ( .A(n_537), .B(n_539), .Y(n_536) );
NAND2xp5_ASAP7_75t_L g637 ( .A(n_537), .B(n_544), .Y(n_637) );
INVx1_ASAP7_75t_SL g537 ( .A(n_538), .Y(n_537) );
AND2x2_ASAP7_75t_L g586 ( .A(n_538), .B(n_541), .Y(n_586) );
AND2x2_ASAP7_75t_L g615 ( .A(n_538), .B(n_559), .Y(n_615) );
OR2x2_ASAP7_75t_L g618 ( .A(n_538), .B(n_578), .Y(n_618) );
AOI222xp33_ASAP7_75t_L g682 ( .A1(n_539), .A2(n_631), .B1(n_683), .B2(n_684), .C1(n_686), .C2(n_688), .Y(n_682) );
BUFx2_ASAP7_75t_L g596 ( .A(n_541), .Y(n_596) );
INVx1_ASAP7_75t_L g542 ( .A(n_543), .Y(n_542) );
AND2x2_ASAP7_75t_L g585 ( .A(n_544), .B(n_586), .Y(n_585) );
INVx3_ASAP7_75t_SL g602 ( .A(n_544), .Y(n_602) );
NAND2xp5_ASAP7_75t_L g656 ( .A(n_544), .B(n_596), .Y(n_656) );
AND2x2_ASAP7_75t_L g591 ( .A(n_546), .B(n_551), .Y(n_591) );
INVx1_ASAP7_75t_L g610 ( .A(n_546), .Y(n_610) );
OAI221xp5_ASAP7_75t_SL g547 ( .A1(n_548), .A2(n_549), .B1(n_553), .B2(n_557), .C(n_561), .Y(n_547) );
OR2x2_ASAP7_75t_L g619 ( .A(n_549), .B(n_620), .Y(n_619) );
INVx1_ASAP7_75t_L g549 ( .A(n_550), .Y(n_549) );
AND2x2_ASAP7_75t_L g550 ( .A(n_551), .B(n_552), .Y(n_550) );
AND2x2_ASAP7_75t_L g604 ( .A(n_551), .B(n_574), .Y(n_604) );
NAND2xp5_ASAP7_75t_L g644 ( .A(n_551), .B(n_564), .Y(n_644) );
AND2x2_ASAP7_75t_L g649 ( .A(n_551), .B(n_599), .Y(n_649) );
HB1xp67_ASAP7_75t_L g659 ( .A(n_551), .Y(n_659) );
NAND2x1_ASAP7_75t_SL g670 ( .A(n_551), .B(n_671), .Y(n_670) );
OR2x2_ASAP7_75t_L g555 ( .A(n_552), .B(n_556), .Y(n_555) );
INVx2_ASAP7_75t_L g575 ( .A(n_552), .Y(n_575) );
NAND2xp5_ASAP7_75t_L g601 ( .A(n_552), .B(n_570), .Y(n_601) );
INVx1_ASAP7_75t_L g667 ( .A(n_552), .Y(n_667) );
INVx1_ASAP7_75t_L g642 ( .A(n_553), .Y(n_642) );
OR2x2_ASAP7_75t_L g553 ( .A(n_554), .B(n_555), .Y(n_553) );
INVx1_ASAP7_75t_L g654 ( .A(n_554), .Y(n_654) );
NOR2xp67_ASAP7_75t_L g666 ( .A(n_554), .B(n_667), .Y(n_666) );
INVx2_ASAP7_75t_L g671 ( .A(n_555), .Y(n_671) );
NOR2xp33_ASAP7_75t_L g678 ( .A(n_555), .B(n_679), .Y(n_678) );
AND2x2_ASAP7_75t_L g574 ( .A(n_556), .B(n_575), .Y(n_574) );
NAND2xp5_ASAP7_75t_L g587 ( .A(n_556), .B(n_566), .Y(n_587) );
INVx1_ASAP7_75t_L g653 ( .A(n_556), .Y(n_653) );
INVx1_ASAP7_75t_L g674 ( .A(n_557), .Y(n_674) );
NAND2xp5_ASAP7_75t_L g557 ( .A(n_558), .B(n_559), .Y(n_557) );
INVx1_ASAP7_75t_L g559 ( .A(n_560), .Y(n_559) );
OAI21xp5_ASAP7_75t_SL g561 ( .A1(n_562), .A2(n_567), .B(n_576), .Y(n_561) );
AND2x2_ASAP7_75t_L g562 ( .A(n_563), .B(n_565), .Y(n_562) );
AND2x2_ASAP7_75t_L g707 ( .A(n_563), .B(n_640), .Y(n_707) );
INVx1_ASAP7_75t_L g563 ( .A(n_564), .Y(n_563) );
AND2x2_ASAP7_75t_L g675 ( .A(n_564), .B(n_635), .Y(n_675) );
AOI32xp33_ASAP7_75t_L g588 ( .A1(n_565), .A2(n_571), .A3(n_589), .B1(n_591), .B2(n_592), .Y(n_588) );
AOI322xp5_ASAP7_75t_L g690 ( .A1(n_565), .A2(n_597), .A3(n_680), .B1(n_691), .B2(n_692), .C1(n_693), .C2(n_695), .Y(n_690) );
INVx2_ASAP7_75t_L g570 ( .A(n_566), .Y(n_570) );
INVx1_ASAP7_75t_L g680 ( .A(n_566), .Y(n_680) );
OAI22xp5_ASAP7_75t_L g567 ( .A1(n_568), .A2(n_571), .B1(n_572), .B2(n_573), .Y(n_567) );
NAND2xp5_ASAP7_75t_L g623 ( .A(n_568), .B(n_574), .Y(n_623) );
AND2x2_ASAP7_75t_L g568 ( .A(n_569), .B(n_570), .Y(n_568) );
NAND2xp5_ASAP7_75t_L g685 ( .A(n_569), .B(n_635), .Y(n_685) );
INVx1_ASAP7_75t_L g572 ( .A(n_570), .Y(n_572) );
NAND2xp5_ASAP7_75t_L g689 ( .A(n_570), .B(n_599), .Y(n_689) );
INVx1_ASAP7_75t_L g573 ( .A(n_574), .Y(n_573) );
INVx1_ASAP7_75t_SL g576 ( .A(n_577), .Y(n_576) );
NOR2xp33_ASAP7_75t_L g672 ( .A(n_578), .B(n_673), .Y(n_672) );
OAI221xp5_ASAP7_75t_SL g579 ( .A1(n_580), .A2(n_581), .B1(n_584), .B2(n_587), .C(n_588), .Y(n_579) );
OR2x2_ASAP7_75t_L g600 ( .A(n_581), .B(n_601), .Y(n_600) );
OR2x2_ASAP7_75t_L g609 ( .A(n_581), .B(n_610), .Y(n_609) );
INVx1_ASAP7_75t_L g581 ( .A(n_582), .Y(n_581) );
AND2x2_ASAP7_75t_L g634 ( .A(n_582), .B(n_635), .Y(n_634) );
INVx2_ASAP7_75t_L g584 ( .A(n_585), .Y(n_584) );
AND2x2_ASAP7_75t_L g638 ( .A(n_592), .B(n_639), .Y(n_638) );
INVx1_ASAP7_75t_L g592 ( .A(n_593), .Y(n_592) );
OAI221xp5_ASAP7_75t_L g594 ( .A1(n_595), .A2(n_598), .B1(n_600), .B2(n_602), .C(n_603), .Y(n_594) );
NAND2xp5_ASAP7_75t_L g595 ( .A(n_596), .B(n_597), .Y(n_595) );
AOI22xp5_ASAP7_75t_L g626 ( .A1(n_596), .A2(n_627), .B1(n_631), .B2(n_632), .Y(n_626) );
NAND2xp5_ASAP7_75t_L g697 ( .A(n_597), .B(n_698), .Y(n_697) );
INVx1_ASAP7_75t_L g702 ( .A(n_597), .Y(n_702) );
INVx1_ASAP7_75t_L g696 ( .A(n_599), .Y(n_696) );
INVx1_ASAP7_75t_SL g631 ( .A(n_600), .Y(n_631) );
NOR2xp33_ASAP7_75t_L g692 ( .A(n_602), .B(n_630), .Y(n_692) );
INVx1_ASAP7_75t_L g605 ( .A(n_606), .Y(n_605) );
NAND2xp5_ASAP7_75t_L g665 ( .A(n_607), .B(n_666), .Y(n_665) );
INVx1_ASAP7_75t_SL g673 ( .A(n_607), .Y(n_673) );
INVx1_ASAP7_75t_SL g608 ( .A(n_609), .Y(n_608) );
OAI221xp5_ASAP7_75t_SL g611 ( .A1(n_612), .A2(n_616), .B1(n_618), .B2(n_619), .C(n_621), .Y(n_611) );
NOR2xp33_ASAP7_75t_SL g612 ( .A(n_613), .B(n_615), .Y(n_612) );
AOI22xp5_ASAP7_75t_L g676 ( .A1(n_613), .A2(n_631), .B1(n_677), .B2(n_678), .Y(n_676) );
CKINVDCx14_ASAP7_75t_R g616 ( .A(n_617), .Y(n_616) );
OAI21xp33_ASAP7_75t_L g695 ( .A1(n_618), .A2(n_696), .B(n_697), .Y(n_695) );
INVx1_ASAP7_75t_L g622 ( .A(n_623), .Y(n_622) );
NOR3xp33_ASAP7_75t_SL g624 ( .A(n_625), .B(n_657), .C(n_681), .Y(n_624) );
NAND4xp25_ASAP7_75t_L g625 ( .A(n_626), .B(n_633), .C(n_641), .D(n_648), .Y(n_625) );
INVx1_ASAP7_75t_L g627 ( .A(n_628), .Y(n_627) );
OR2x2_ASAP7_75t_L g628 ( .A(n_629), .B(n_630), .Y(n_628) );
INVx1_ASAP7_75t_L g704 ( .A(n_629), .Y(n_704) );
INVx3_ASAP7_75t_SL g698 ( .A(n_630), .Y(n_698) );
OR2x2_ASAP7_75t_L g703 ( .A(n_630), .B(n_704), .Y(n_703) );
AOI22xp5_ASAP7_75t_L g633 ( .A1(n_634), .A2(n_636), .B1(n_638), .B2(n_640), .Y(n_633) );
NAND2xp5_ASAP7_75t_L g694 ( .A(n_635), .B(n_653), .Y(n_694) );
INVxp67_ASAP7_75t_L g636 ( .A(n_637), .Y(n_636) );
OAI21xp5_ASAP7_75t_SL g641 ( .A1(n_642), .A2(n_643), .B(n_645), .Y(n_641) );
INVxp67_ASAP7_75t_L g643 ( .A(n_644), .Y(n_643) );
INVx1_ASAP7_75t_L g645 ( .A(n_646), .Y(n_645) );
INVx1_ASAP7_75t_L g650 ( .A(n_651), .Y(n_650) );
NAND2xp5_ASAP7_75t_L g651 ( .A(n_652), .B(n_654), .Y(n_651) );
INVxp67_ASAP7_75t_L g652 ( .A(n_653), .Y(n_652) );
INVx1_ASAP7_75t_L g655 ( .A(n_656), .Y(n_655) );
OAI211xp5_ASAP7_75t_SL g657 ( .A1(n_658), .A2(n_660), .B(n_663), .C(n_676), .Y(n_657) );
INVx1_ASAP7_75t_L g658 ( .A(n_659), .Y(n_658) );
INVx1_ASAP7_75t_L g660 ( .A(n_661), .Y(n_660) );
INVx1_ASAP7_75t_L g691 ( .A(n_662), .Y(n_691) );
AOI222xp33_ASAP7_75t_L g663 ( .A1(n_664), .A2(n_668), .B1(n_669), .B2(n_672), .C1(n_674), .C2(n_675), .Y(n_663) );
INVxp67_ASAP7_75t_L g664 ( .A(n_665), .Y(n_664) );
INVx1_ASAP7_75t_L g669 ( .A(n_670), .Y(n_669) );
NAND4xp25_ASAP7_75t_SL g700 ( .A(n_673), .B(n_701), .C(n_702), .D(n_703), .Y(n_700) );
INVx1_ASAP7_75t_L g679 ( .A(n_680), .Y(n_679) );
NAND3xp33_ASAP7_75t_SL g681 ( .A(n_682), .B(n_690), .C(n_699), .Y(n_681) );
INVx1_ASAP7_75t_L g684 ( .A(n_685), .Y(n_684) );
INVx1_ASAP7_75t_L g686 ( .A(n_687), .Y(n_686) );
INVx1_ASAP7_75t_L g688 ( .A(n_689), .Y(n_688) );
INVx1_ASAP7_75t_L g693 ( .A(n_694), .Y(n_693) );
AOI22xp33_ASAP7_75t_L g699 ( .A1(n_700), .A2(n_705), .B1(n_706), .B2(n_707), .Y(n_699) );
OAI22xp5_ASAP7_75t_L g711 ( .A1(n_708), .A2(n_712), .B1(n_713), .B2(n_715), .Y(n_711) );
INVx1_ASAP7_75t_L g714 ( .A(n_710), .Y(n_714) );
INVx2_ASAP7_75t_L g713 ( .A(n_714), .Y(n_713) );
INVx1_ASAP7_75t_SL g717 ( .A(n_718), .Y(n_717) );
INVx2_ASAP7_75t_L g718 ( .A(n_719), .Y(n_718) );
INVx1_ASAP7_75t_L g720 ( .A(n_721), .Y(n_720) );
endmodule