module fake_jpeg_3888_n_162 (n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_162);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_162;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_147;
wire n_158;
wire n_14;
wire n_73;
wire n_152;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_106;
wire n_111;
wire n_24;
wire n_44;
wire n_143;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_78;
wire n_20;
wire n_18;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_161;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_153;
wire n_135;
wire n_36;
wire n_62;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

INVx1_ASAP7_75t_L g13 ( 
.A(n_8),
.Y(n_13)
);

INVx8_ASAP7_75t_L g14 ( 
.A(n_9),
.Y(n_14)
);

BUFx6f_ASAP7_75t_L g15 ( 
.A(n_12),
.Y(n_15)
);

INVx3_ASAP7_75t_L g16 ( 
.A(n_7),
.Y(n_16)
);

BUFx8_ASAP7_75t_L g17 ( 
.A(n_10),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_4),
.Y(n_18)
);

BUFx10_ASAP7_75t_L g19 ( 
.A(n_0),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_5),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_0),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_2),
.Y(n_22)
);

BUFx3_ASAP7_75t_L g23 ( 
.A(n_0),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_12),
.Y(n_24)
);

INVx8_ASAP7_75t_L g25 ( 
.A(n_4),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_10),
.Y(n_26)
);

BUFx2_ASAP7_75t_L g27 ( 
.A(n_4),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_6),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_2),
.Y(n_29)
);

INVx3_ASAP7_75t_L g30 ( 
.A(n_27),
.Y(n_30)
);

NOR2xp33_ASAP7_75t_L g46 ( 
.A(n_30),
.B(n_31),
.Y(n_46)
);

BUFx3_ASAP7_75t_L g31 ( 
.A(n_15),
.Y(n_31)
);

NOR2xp33_ASAP7_75t_L g32 ( 
.A(n_13),
.B(n_1),
.Y(n_32)
);

NOR2xp33_ASAP7_75t_SL g64 ( 
.A(n_32),
.B(n_16),
.Y(n_64)
);

INVx3_ASAP7_75t_L g33 ( 
.A(n_27),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_33),
.B(n_38),
.Y(n_52)
);

INVx8_ASAP7_75t_L g34 ( 
.A(n_23),
.Y(n_34)
);

AOI22xp33_ASAP7_75t_SL g69 ( 
.A1(n_34),
.A2(n_36),
.B1(n_41),
.B2(n_14),
.Y(n_69)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_15),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_35),
.Y(n_55)
);

INVx6_ASAP7_75t_L g36 ( 
.A(n_15),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_26),
.Y(n_37)
);

BUFx3_ASAP7_75t_L g44 ( 
.A(n_37),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_26),
.Y(n_38)
);

BUFx3_ASAP7_75t_L g39 ( 
.A(n_26),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_39),
.B(n_40),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_25),
.Y(n_40)
);

INVx8_ASAP7_75t_L g41 ( 
.A(n_23),
.Y(n_41)
);

NAND3xp33_ASAP7_75t_L g42 ( 
.A(n_20),
.B(n_21),
.C(n_28),
.Y(n_42)
);

AND2x2_ASAP7_75t_L g56 ( 
.A(n_42),
.B(n_20),
.Y(n_56)
);

AOI21xp33_ASAP7_75t_L g43 ( 
.A1(n_19),
.A2(n_28),
.B(n_22),
.Y(n_43)
);

OAI21xp5_ASAP7_75t_SL g66 ( 
.A1(n_43),
.A2(n_19),
.B(n_16),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_L g45 ( 
.A(n_31),
.B(n_29),
.Y(n_45)
);

NAND2xp5_ASAP7_75t_SL g83 ( 
.A(n_45),
.B(n_49),
.Y(n_83)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_39),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_47),
.B(n_48),
.Y(n_72)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_30),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_SL g49 ( 
.A(n_36),
.B(n_24),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_L g50 ( 
.A(n_35),
.B(n_29),
.Y(n_50)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_50),
.Y(n_85)
);

CKINVDCx16_ASAP7_75t_R g51 ( 
.A(n_34),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_51),
.B(n_54),
.Y(n_79)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_41),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_56),
.B(n_58),
.Y(n_81)
);

OAI32xp33_ASAP7_75t_L g57 ( 
.A1(n_40),
.A2(n_24),
.A3(n_13),
.B1(n_18),
.B2(n_17),
.Y(n_57)
);

OAI22xp5_ASAP7_75t_SL g78 ( 
.A1(n_57),
.A2(n_59),
.B1(n_67),
.B2(n_17),
.Y(n_78)
);

CKINVDCx12_ASAP7_75t_R g58 ( 
.A(n_37),
.Y(n_58)
);

A2O1A1Ixp33_ASAP7_75t_SL g59 ( 
.A1(n_38),
.A2(n_19),
.B(n_27),
.C(n_25),
.Y(n_59)
);

MAJIxp5_ASAP7_75t_L g60 ( 
.A(n_43),
.B(n_22),
.C(n_21),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_60),
.B(n_61),
.Y(n_87)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_31),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_32),
.B(n_18),
.Y(n_62)
);

CKINVDCx16_ASAP7_75t_R g73 ( 
.A(n_62),
.Y(n_73)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_31),
.Y(n_63)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_63),
.Y(n_86)
);

CKINVDCx20_ASAP7_75t_R g82 ( 
.A(n_64),
.Y(n_82)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_31),
.Y(n_65)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_65),
.Y(n_89)
);

NAND2xp33_ASAP7_75t_SL g92 ( 
.A(n_66),
.B(n_70),
.Y(n_92)
);

AOI22xp5_ASAP7_75t_L g67 ( 
.A1(n_43),
.A2(n_16),
.B1(n_25),
.B2(n_14),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_32),
.B(n_23),
.Y(n_68)
);

CKINVDCx20_ASAP7_75t_R g91 ( 
.A(n_68),
.Y(n_91)
);

INVxp67_ASAP7_75t_L g76 ( 
.A(n_69),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_L g70 ( 
.A(n_32),
.B(n_19),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_SL g71 ( 
.A(n_32),
.B(n_14),
.Y(n_71)
);

OAI22xp33_ASAP7_75t_SL g77 ( 
.A1(n_71),
.A2(n_17),
.B1(n_11),
.B2(n_9),
.Y(n_77)
);

BUFx6f_ASAP7_75t_L g74 ( 
.A(n_55),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_74),
.B(n_80),
.Y(n_94)
);

OAI22x1_ASAP7_75t_L g75 ( 
.A1(n_57),
.A2(n_19),
.B1(n_17),
.B2(n_3),
.Y(n_75)
);

AOI22xp33_ASAP7_75t_L g102 ( 
.A1(n_75),
.A2(n_59),
.B1(n_65),
.B2(n_63),
.Y(n_102)
);

NOR3xp33_ASAP7_75t_L g104 ( 
.A(n_77),
.B(n_75),
.C(n_81),
.Y(n_104)
);

XOR2xp5_ASAP7_75t_L g96 ( 
.A(n_78),
.B(n_60),
.Y(n_96)
);

INVx5_ASAP7_75t_L g80 ( 
.A(n_44),
.Y(n_80)
);

AOI22xp33_ASAP7_75t_SL g84 ( 
.A1(n_54),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_84)
);

AOI21xp5_ASAP7_75t_L g109 ( 
.A1(n_84),
.A2(n_52),
.B(n_46),
.Y(n_109)
);

AO22x1_ASAP7_75t_SL g88 ( 
.A1(n_66),
.A2(n_1),
.B1(n_3),
.B2(n_5),
.Y(n_88)
);

OAI22xp5_ASAP7_75t_SL g98 ( 
.A1(n_88),
.A2(n_90),
.B1(n_59),
.B2(n_71),
.Y(n_98)
);

OAI22xp5_ASAP7_75t_SL g90 ( 
.A1(n_67),
.A2(n_5),
.B1(n_6),
.B2(n_7),
.Y(n_90)
);

INVx2_ASAP7_75t_L g93 ( 
.A(n_44),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_93),
.B(n_55),
.Y(n_95)
);

CKINVDCx20_ASAP7_75t_R g121 ( 
.A(n_95),
.Y(n_121)
);

MAJIxp5_ASAP7_75t_L g118 ( 
.A(n_96),
.B(n_97),
.C(n_100),
.Y(n_118)
);

AND2x6_ASAP7_75t_L g97 ( 
.A(n_92),
.B(n_88),
.Y(n_97)
);

XNOR2xp5_ASAP7_75t_SL g125 ( 
.A(n_98),
.B(n_101),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_82),
.B(n_56),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_SL g114 ( 
.A(n_99),
.B(n_110),
.Y(n_114)
);

MAJIxp5_ASAP7_75t_L g100 ( 
.A(n_87),
.B(n_45),
.C(n_48),
.Y(n_100)
);

XOR2xp5_ASAP7_75t_SL g101 ( 
.A(n_92),
.B(n_56),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_L g120 ( 
.A(n_102),
.B(n_104),
.Y(n_120)
);

AND2x6_ASAP7_75t_L g103 ( 
.A(n_88),
.B(n_59),
.Y(n_103)
);

MAJIxp5_ASAP7_75t_L g119 ( 
.A(n_103),
.B(n_107),
.C(n_90),
.Y(n_119)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_72),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_SL g123 ( 
.A(n_105),
.B(n_106),
.Y(n_123)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_79),
.Y(n_106)
);

AND2x6_ASAP7_75t_L g107 ( 
.A(n_78),
.B(n_59),
.Y(n_107)
);

OAI21xp5_ASAP7_75t_SL g108 ( 
.A1(n_85),
.A2(n_50),
.B(n_70),
.Y(n_108)
);

AOI21xp5_ASAP7_75t_L g122 ( 
.A1(n_108),
.A2(n_109),
.B(n_111),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_82),
.B(n_6),
.Y(n_110)
);

OAI21xp33_ASAP7_75t_L g111 ( 
.A1(n_83),
.A2(n_53),
.B(n_7),
.Y(n_111)
);

CKINVDCx16_ASAP7_75t_R g112 ( 
.A(n_94),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_L g131 ( 
.A(n_112),
.B(n_113),
.Y(n_131)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_98),
.Y(n_113)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_100),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_L g134 ( 
.A(n_115),
.B(n_89),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_L g116 ( 
.A(n_96),
.B(n_85),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_L g128 ( 
.A(n_116),
.B(n_108),
.Y(n_128)
);

INVxp67_ASAP7_75t_L g117 ( 
.A(n_109),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_SL g132 ( 
.A(n_117),
.B(n_106),
.Y(n_132)
);

AOI22xp5_ASAP7_75t_L g130 ( 
.A1(n_119),
.A2(n_124),
.B1(n_99),
.B2(n_110),
.Y(n_130)
);

AOI22xp5_ASAP7_75t_L g124 ( 
.A1(n_107),
.A2(n_76),
.B1(n_91),
.B2(n_61),
.Y(n_124)
);

AOI21xp5_ASAP7_75t_L g126 ( 
.A1(n_103),
.A2(n_76),
.B(n_91),
.Y(n_126)
);

OAI21xp5_ASAP7_75t_SL g127 ( 
.A1(n_126),
.A2(n_97),
.B(n_101),
.Y(n_127)
);

XNOR2xp5_ASAP7_75t_L g140 ( 
.A(n_127),
.B(n_130),
.Y(n_140)
);

MAJIxp5_ASAP7_75t_L g138 ( 
.A(n_128),
.B(n_133),
.C(n_125),
.Y(n_138)
);

CKINVDCx20_ASAP7_75t_R g129 ( 
.A(n_123),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_SL g141 ( 
.A(n_129),
.B(n_136),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_L g143 ( 
.A(n_132),
.B(n_135),
.Y(n_143)
);

MAJIxp5_ASAP7_75t_L g133 ( 
.A(n_116),
.B(n_105),
.C(n_73),
.Y(n_133)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_134),
.Y(n_144)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_120),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_L g136 ( 
.A(n_121),
.B(n_89),
.Y(n_136)
);

OAI21x1_ASAP7_75t_L g137 ( 
.A1(n_131),
.A2(n_117),
.B(n_125),
.Y(n_137)
);

OAI21xp5_ASAP7_75t_L g149 ( 
.A1(n_137),
.A2(n_122),
.B(n_114),
.Y(n_149)
);

MAJIxp5_ASAP7_75t_L g147 ( 
.A(n_138),
.B(n_142),
.C(n_127),
.Y(n_147)
);

CKINVDCx20_ASAP7_75t_R g139 ( 
.A(n_130),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_L g151 ( 
.A(n_139),
.B(n_145),
.Y(n_151)
);

MAJIxp5_ASAP7_75t_L g142 ( 
.A(n_128),
.B(n_118),
.C(n_115),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_L g145 ( 
.A(n_133),
.B(n_121),
.Y(n_145)
);

XOR2xp5_ASAP7_75t_L g146 ( 
.A(n_140),
.B(n_118),
.Y(n_146)
);

MAJIxp5_ASAP7_75t_L g154 ( 
.A(n_146),
.B(n_147),
.C(n_149),
.Y(n_154)
);

AO22x1_ASAP7_75t_L g148 ( 
.A1(n_143),
.A2(n_124),
.B1(n_126),
.B2(n_113),
.Y(n_148)
);

NOR2xp33_ASAP7_75t_L g152 ( 
.A(n_148),
.B(n_122),
.Y(n_152)
);

AND2x2_ASAP7_75t_L g150 ( 
.A(n_140),
.B(n_119),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_L g155 ( 
.A(n_150),
.B(n_141),
.Y(n_155)
);

AO21x1_ASAP7_75t_L g158 ( 
.A1(n_152),
.A2(n_153),
.B(n_150),
.Y(n_158)
);

NAND5xp2_ASAP7_75t_L g153 ( 
.A(n_148),
.B(n_142),
.C(n_138),
.D(n_144),
.E(n_114),
.Y(n_153)
);

MAJIxp5_ASAP7_75t_L g156 ( 
.A(n_155),
.B(n_147),
.C(n_146),
.Y(n_156)
);

INVxp67_ASAP7_75t_L g160 ( 
.A(n_156),
.Y(n_160)
);

NOR2xp33_ASAP7_75t_L g157 ( 
.A(n_152),
.B(n_151),
.Y(n_157)
);

AOI21xp5_ASAP7_75t_SL g159 ( 
.A1(n_157),
.A2(n_158),
.B(n_154),
.Y(n_159)
);

AOI21xp5_ASAP7_75t_L g161 ( 
.A1(n_159),
.A2(n_160),
.B(n_86),
.Y(n_161)
);

XOR2xp5_ASAP7_75t_L g162 ( 
.A(n_161),
.B(n_80),
.Y(n_162)
);


endmodule