module fake_netlist_5_1331_n_1660 (n_137, n_91, n_82, n_122, n_142, n_10, n_140, n_24, n_124, n_86, n_136, n_146, n_143, n_83, n_132, n_61, n_90, n_127, n_75, n_101, n_65, n_78, n_74, n_144, n_114, n_57, n_96, n_37, n_111, n_108, n_129, n_31, n_13, n_66, n_98, n_60, n_152, n_16, n_43, n_107, n_0, n_58, n_9, n_69, n_18, n_116, n_42, n_22, n_1, n_45, n_117, n_46, n_21, n_94, n_113, n_38, n_123, n_139, n_105, n_80, n_4, n_125, n_35, n_128, n_73, n_17, n_92, n_19, n_149, n_120, n_135, n_30, n_5, n_33, n_126, n_14, n_84, n_23, n_130, n_29, n_79, n_131, n_151, n_47, n_25, n_53, n_8, n_44, n_40, n_34, n_100, n_62, n_138, n_148, n_71, n_109, n_112, n_85, n_95, n_119, n_59, n_26, n_133, n_55, n_99, n_2, n_3, n_49, n_20, n_6, n_39, n_54, n_147, n_12, n_67, n_121, n_36, n_76, n_87, n_150, n_27, n_64, n_77, n_102, n_106, n_81, n_118, n_28, n_89, n_70, n_115, n_68, n_93, n_72, n_134, n_32, n_41, n_104, n_103, n_56, n_51, n_63, n_97, n_141, n_11, n_153, n_7, n_15, n_145, n_48, n_50, n_52, n_88, n_110, n_1660);

input n_137;
input n_91;
input n_82;
input n_122;
input n_142;
input n_10;
input n_140;
input n_24;
input n_124;
input n_86;
input n_136;
input n_146;
input n_143;
input n_83;
input n_132;
input n_61;
input n_90;
input n_127;
input n_75;
input n_101;
input n_65;
input n_78;
input n_74;
input n_144;
input n_114;
input n_57;
input n_96;
input n_37;
input n_111;
input n_108;
input n_129;
input n_31;
input n_13;
input n_66;
input n_98;
input n_60;
input n_152;
input n_16;
input n_43;
input n_107;
input n_0;
input n_58;
input n_9;
input n_69;
input n_18;
input n_116;
input n_42;
input n_22;
input n_1;
input n_45;
input n_117;
input n_46;
input n_21;
input n_94;
input n_113;
input n_38;
input n_123;
input n_139;
input n_105;
input n_80;
input n_4;
input n_125;
input n_35;
input n_128;
input n_73;
input n_17;
input n_92;
input n_19;
input n_149;
input n_120;
input n_135;
input n_30;
input n_5;
input n_33;
input n_126;
input n_14;
input n_84;
input n_23;
input n_130;
input n_29;
input n_79;
input n_131;
input n_151;
input n_47;
input n_25;
input n_53;
input n_8;
input n_44;
input n_40;
input n_34;
input n_100;
input n_62;
input n_138;
input n_148;
input n_71;
input n_109;
input n_112;
input n_85;
input n_95;
input n_119;
input n_59;
input n_26;
input n_133;
input n_55;
input n_99;
input n_2;
input n_3;
input n_49;
input n_20;
input n_6;
input n_39;
input n_54;
input n_147;
input n_12;
input n_67;
input n_121;
input n_36;
input n_76;
input n_87;
input n_150;
input n_27;
input n_64;
input n_77;
input n_102;
input n_106;
input n_81;
input n_118;
input n_28;
input n_89;
input n_70;
input n_115;
input n_68;
input n_93;
input n_72;
input n_134;
input n_32;
input n_41;
input n_104;
input n_103;
input n_56;
input n_51;
input n_63;
input n_97;
input n_141;
input n_11;
input n_153;
input n_7;
input n_15;
input n_145;
input n_48;
input n_50;
input n_52;
input n_88;
input n_110;

output n_1660;

wire n_924;
wire n_1263;
wire n_977;
wire n_1378;
wire n_611;
wire n_1126;
wire n_1423;
wire n_1166;
wire n_469;
wire n_1508;
wire n_785;
wire n_549;
wire n_532;
wire n_1161;
wire n_1150;
wire n_226;
wire n_1488;
wire n_667;
wire n_790;
wire n_1055;
wire n_1501;
wire n_880;
wire n_544;
wire n_1007;
wire n_155;
wire n_552;
wire n_1528;
wire n_1370;
wire n_1292;
wire n_1198;
wire n_1360;
wire n_1099;
wire n_956;
wire n_564;
wire n_423;
wire n_1021;
wire n_551;
wire n_1323;
wire n_1466;
wire n_688;
wire n_1353;
wire n_800;
wire n_1347;
wire n_1535;
wire n_671;
wire n_819;
wire n_1451;
wire n_1022;
wire n_915;
wire n_1545;
wire n_864;
wire n_173;
wire n_859;
wire n_951;
wire n_1264;
wire n_447;
wire n_247;
wire n_1494;
wire n_292;
wire n_625;
wire n_854;
wire n_1462;
wire n_1580;
wire n_674;
wire n_417;
wire n_516;
wire n_933;
wire n_1152;
wire n_497;
wire n_1607;
wire n_1563;
wire n_606;
wire n_275;
wire n_877;
wire n_755;
wire n_1118;
wire n_947;
wire n_1285;
wire n_373;
wire n_307;
wire n_1359;
wire n_530;
wire n_1107;
wire n_556;
wire n_1230;
wire n_668;
wire n_375;
wire n_301;
wire n_929;
wire n_1124;
wire n_902;
wire n_1576;
wire n_191;
wire n_1104;
wire n_1294;
wire n_659;
wire n_1257;
wire n_171;
wire n_1182;
wire n_579;
wire n_1261;
wire n_938;
wire n_1098;
wire n_320;
wire n_1154;
wire n_1242;
wire n_1135;
wire n_406;
wire n_519;
wire n_1016;
wire n_1243;
wire n_546;
wire n_1280;
wire n_281;
wire n_240;
wire n_291;
wire n_231;
wire n_257;
wire n_731;
wire n_371;
wire n_1483;
wire n_1314;
wire n_1512;
wire n_709;
wire n_1490;
wire n_317;
wire n_1236;
wire n_1633;
wire n_569;
wire n_227;
wire n_920;
wire n_1289;
wire n_1517;
wire n_335;
wire n_370;
wire n_976;
wire n_343;
wire n_1449;
wire n_308;
wire n_1566;
wire n_297;
wire n_156;
wire n_1078;
wire n_775;
wire n_219;
wire n_157;
wire n_600;
wire n_1484;
wire n_1374;
wire n_1328;
wire n_223;
wire n_264;
wire n_1598;
wire n_955;
wire n_163;
wire n_339;
wire n_1146;
wire n_882;
wire n_183;
wire n_243;
wire n_1036;
wire n_1097;
wire n_347;
wire n_550;
wire n_696;
wire n_897;
wire n_215;
wire n_350;
wire n_196;
wire n_798;
wire n_646;
wire n_1428;
wire n_436;
wire n_1394;
wire n_1414;
wire n_1216;
wire n_290;
wire n_580;
wire n_1040;
wire n_578;
wire n_926;
wire n_344;
wire n_1218;
wire n_422;
wire n_475;
wire n_777;
wire n_1070;
wire n_1547;
wire n_1030;
wire n_415;
wire n_1071;
wire n_485;
wire n_1165;
wire n_1267;
wire n_1561;
wire n_496;
wire n_1391;
wire n_958;
wire n_1034;
wire n_670;
wire n_1513;
wire n_1600;
wire n_521;
wire n_663;
wire n_845;
wire n_673;
wire n_837;
wire n_1239;
wire n_528;
wire n_680;
wire n_1473;
wire n_1587;
wire n_395;
wire n_164;
wire n_553;
wire n_901;
wire n_813;
wire n_1521;
wire n_1284;
wire n_1590;
wire n_214;
wire n_675;
wire n_888;
wire n_1167;
wire n_1626;
wire n_637;
wire n_1384;
wire n_1556;
wire n_184;
wire n_446;
wire n_1064;
wire n_858;
wire n_923;
wire n_691;
wire n_1151;
wire n_881;
wire n_1405;
wire n_468;
wire n_213;
wire n_342;
wire n_464;
wire n_363;
wire n_1582;
wire n_197;
wire n_1069;
wire n_1075;
wire n_1450;
wire n_1322;
wire n_1471;
wire n_1459;
wire n_460;
wire n_889;
wire n_973;
wire n_477;
wire n_571;
wire n_1585;
wire n_461;
wire n_1599;
wire n_1211;
wire n_1197;
wire n_1523;
wire n_907;
wire n_1447;
wire n_1377;
wire n_190;
wire n_989;
wire n_1039;
wire n_228;
wire n_283;
wire n_1403;
wire n_488;
wire n_736;
wire n_892;
wire n_1000;
wire n_1202;
wire n_1278;
wire n_1002;
wire n_1463;
wire n_1581;
wire n_310;
wire n_593;
wire n_748;
wire n_586;
wire n_1058;
wire n_838;
wire n_332;
wire n_1053;
wire n_1224;
wire n_349;
wire n_1248;
wire n_230;
wire n_1331;
wire n_953;
wire n_279;
wire n_1014;
wire n_1241;
wire n_289;
wire n_963;
wire n_1052;
wire n_954;
wire n_627;
wire n_1385;
wire n_440;
wire n_793;
wire n_478;
wire n_476;
wire n_1527;
wire n_534;
wire n_884;
wire n_345;
wire n_944;
wire n_1623;
wire n_1565;
wire n_182;
wire n_647;
wire n_237;
wire n_407;
wire n_1072;
wire n_832;
wire n_857;
wire n_207;
wire n_561;
wire n_1319;
wire n_1387;
wire n_1532;
wire n_1027;
wire n_971;
wire n_1156;
wire n_326;
wire n_794;
wire n_404;
wire n_686;
wire n_847;
wire n_1393;
wire n_596;
wire n_1368;
wire n_558;
wire n_702;
wire n_1276;
wire n_822;
wire n_1412;
wire n_728;
wire n_266;
wire n_1162;
wire n_272;
wire n_1538;
wire n_1199;
wire n_352;
wire n_1038;
wire n_520;
wire n_1369;
wire n_409;
wire n_887;
wire n_154;
wire n_300;
wire n_809;
wire n_870;
wire n_931;
wire n_599;
wire n_1481;
wire n_434;
wire n_1544;
wire n_868;
wire n_639;
wire n_914;
wire n_411;
wire n_414;
wire n_1629;
wire n_1293;
wire n_965;
wire n_935;
wire n_1175;
wire n_817;
wire n_360;
wire n_1479;
wire n_759;
wire n_806;
wire n_1477;
wire n_324;
wire n_1635;
wire n_1571;
wire n_187;
wire n_1189;
wire n_1259;
wire n_706;
wire n_746;
wire n_1649;
wire n_747;
wire n_784;
wire n_1244;
wire n_431;
wire n_1194;
wire n_615;
wire n_851;
wire n_843;
wire n_523;
wire n_913;
wire n_1537;
wire n_705;
wire n_865;
wire n_678;
wire n_697;
wire n_1222;
wire n_776;
wire n_1415;
wire n_367;
wire n_452;
wire n_525;
wire n_1260;
wire n_1647;
wire n_1464;
wire n_649;
wire n_547;
wire n_1444;
wire n_1191;
wire n_284;
wire n_1128;
wire n_744;
wire n_629;
wire n_590;
wire n_1308;
wire n_254;
wire n_1233;
wire n_1615;
wire n_1529;
wire n_526;
wire n_372;
wire n_293;
wire n_677;
wire n_244;
wire n_1333;
wire n_1121;
wire n_314;
wire n_368;
wire n_433;
wire n_604;
wire n_949;
wire n_1443;
wire n_1008;
wire n_946;
wire n_1539;
wire n_1001;
wire n_1503;
wire n_498;
wire n_1468;
wire n_1559;
wire n_689;
wire n_738;
wire n_1624;
wire n_640;
wire n_1510;
wire n_252;
wire n_624;
wire n_1380;
wire n_1617;
wire n_295;
wire n_1010;
wire n_1231;
wire n_739;
wire n_1279;
wire n_1406;
wire n_1195;
wire n_610;
wire n_936;
wire n_568;
wire n_1500;
wire n_1090;
wire n_757;
wire n_633;
wire n_439;
wire n_259;
wire n_448;
wire n_758;
wire n_999;
wire n_1656;
wire n_1158;
wire n_1509;
wire n_563;
wire n_1145;
wire n_878;
wire n_524;
wire n_204;
wire n_394;
wire n_1049;
wire n_1153;
wire n_741;
wire n_1639;
wire n_1306;
wire n_1068;
wire n_331;
wire n_906;
wire n_1163;
wire n_1207;
wire n_919;
wire n_908;
wire n_724;
wire n_658;
wire n_1362;
wire n_1586;
wire n_456;
wire n_959;
wire n_535;
wire n_940;
wire n_1445;
wire n_1492;
wire n_592;
wire n_1169;
wire n_1596;
wire n_1017;
wire n_978;
wire n_1434;
wire n_1054;
wire n_1474;
wire n_1269;
wire n_1095;
wire n_1614;
wire n_267;
wire n_514;
wire n_457;
wire n_1079;
wire n_1045;
wire n_1208;
wire n_603;
wire n_1431;
wire n_484;
wire n_1593;
wire n_1033;
wire n_442;
wire n_636;
wire n_660;
wire n_1640;
wire n_1009;
wire n_1148;
wire n_742;
wire n_750;
wire n_995;
wire n_454;
wire n_1609;
wire n_374;
wire n_185;
wire n_396;
wire n_1383;
wire n_1073;
wire n_255;
wire n_662;
wire n_459;
wire n_218;
wire n_962;
wire n_1215;
wire n_1171;
wire n_1578;
wire n_723;
wire n_1065;
wire n_1592;
wire n_1336;
wire n_1574;
wire n_473;
wire n_1309;
wire n_1426;
wire n_1043;
wire n_355;
wire n_486;
wire n_1548;
wire n_614;
wire n_337;
wire n_1421;
wire n_1286;
wire n_1177;
wire n_1355;
wire n_168;
wire n_974;
wire n_727;
wire n_1159;
wire n_957;
wire n_773;
wire n_208;
wire n_743;
wire n_299;
wire n_303;
wire n_296;
wire n_613;
wire n_1119;
wire n_1240;
wire n_829;
wire n_1612;
wire n_1416;
wire n_361;
wire n_700;
wire n_1237;
wire n_573;
wire n_1420;
wire n_1132;
wire n_388;
wire n_1366;
wire n_1300;
wire n_1127;
wire n_761;
wire n_1568;
wire n_1006;
wire n_329;
wire n_274;
wire n_1270;
wire n_1486;
wire n_582;
wire n_1332;
wire n_1390;
wire n_309;
wire n_512;
wire n_1591;
wire n_322;
wire n_1249;
wire n_652;
wire n_1111;
wire n_1365;
wire n_1349;
wire n_1093;
wire n_288;
wire n_1031;
wire n_263;
wire n_609;
wire n_1041;
wire n_1265;
wire n_224;
wire n_1562;
wire n_383;
wire n_834;
wire n_765;
wire n_893;
wire n_1015;
wire n_1140;
wire n_891;
wire n_1651;
wire n_239;
wire n_630;
wire n_504;
wire n_511;
wire n_874;
wire n_358;
wire n_1101;
wire n_1106;
wire n_1456;
wire n_1304;
wire n_1324;
wire n_987;
wire n_261;
wire n_174;
wire n_1455;
wire n_767;
wire n_993;
wire n_1407;
wire n_1551;
wire n_545;
wire n_441;
wire n_860;
wire n_450;
wire n_429;
wire n_948;
wire n_1217;
wire n_628;
wire n_365;
wire n_729;
wire n_1131;
wire n_1084;
wire n_970;
wire n_911;
wire n_1430;
wire n_513;
wire n_1094;
wire n_1354;
wire n_560;
wire n_1534;
wire n_340;
wire n_1351;
wire n_1044;
wire n_1205;
wire n_346;
wire n_1209;
wire n_1552;
wire n_495;
wire n_602;
wire n_574;
wire n_1435;
wire n_879;
wire n_623;
wire n_405;
wire n_824;
wire n_359;
wire n_1645;
wire n_490;
wire n_1327;
wire n_996;
wire n_921;
wire n_233;
wire n_572;
wire n_366;
wire n_815;
wire n_327;
wire n_1381;
wire n_1611;
wire n_1037;
wire n_1080;
wire n_1274;
wire n_1316;
wire n_426;
wire n_1438;
wire n_1082;
wire n_589;
wire n_716;
wire n_1630;
wire n_562;
wire n_1436;
wire n_952;
wire n_1229;
wire n_391;
wire n_701;
wire n_1437;
wire n_1023;
wire n_645;
wire n_539;
wire n_803;
wire n_1092;
wire n_238;
wire n_531;
wire n_890;
wire n_764;
wire n_1056;
wire n_1424;
wire n_162;
wire n_960;
wire n_222;
wire n_1290;
wire n_1123;
wire n_1467;
wire n_1047;
wire n_634;
wire n_199;
wire n_1252;
wire n_348;
wire n_1382;
wire n_1029;
wire n_925;
wire n_1206;
wire n_424;
wire n_1311;
wire n_1519;
wire n_256;
wire n_950;
wire n_1553;
wire n_380;
wire n_419;
wire n_1346;
wire n_444;
wire n_1299;
wire n_1060;
wire n_1141;
wire n_316;
wire n_389;
wire n_418;
wire n_248;
wire n_912;
wire n_315;
wire n_968;
wire n_451;
wire n_619;
wire n_408;
wire n_1386;
wire n_376;
wire n_967;
wire n_1442;
wire n_1139;
wire n_515;
wire n_351;
wire n_885;
wire n_397;
wire n_1432;
wire n_1357;
wire n_483;
wire n_683;
wire n_1632;
wire n_1057;
wire n_1051;
wire n_1085;
wire n_1066;
wire n_721;
wire n_1157;
wire n_841;
wire n_1050;
wire n_802;
wire n_1608;
wire n_983;
wire n_280;
wire n_1305;
wire n_873;
wire n_378;
wire n_1112;
wire n_762;
wire n_1283;
wire n_1644;
wire n_690;
wire n_583;
wire n_302;
wire n_1343;
wire n_1203;
wire n_1631;
wire n_821;
wire n_321;
wire n_1179;
wire n_621;
wire n_753;
wire n_455;
wire n_1048;
wire n_1288;
wire n_385;
wire n_212;
wire n_507;
wire n_1560;
wire n_1605;
wire n_330;
wire n_1228;
wire n_972;
wire n_692;
wire n_820;
wire n_1200;
wire n_1301;
wire n_1363;
wire n_1185;
wire n_991;
wire n_828;
wire n_779;
wire n_576;
wire n_1143;
wire n_1579;
wire n_1329;
wire n_1312;
wire n_1439;
wire n_804;
wire n_537;
wire n_945;
wire n_492;
wire n_1504;
wire n_943;
wire n_341;
wire n_250;
wire n_992;
wire n_543;
wire n_260;
wire n_842;
wire n_650;
wire n_984;
wire n_694;
wire n_286;
wire n_1643;
wire n_883;
wire n_470;
wire n_325;
wire n_449;
wire n_1594;
wire n_1214;
wire n_1342;
wire n_1400;
wire n_900;
wire n_856;
wire n_918;
wire n_942;
wire n_189;
wire n_1147;
wire n_1557;
wire n_1610;
wire n_1077;
wire n_1422;
wire n_540;
wire n_618;
wire n_896;
wire n_323;
wire n_195;
wire n_356;
wire n_894;
wire n_1636;
wire n_831;
wire n_964;
wire n_1373;
wire n_1350;
wire n_1511;
wire n_1470;
wire n_1096;
wire n_234;
wire n_1575;
wire n_833;
wire n_1646;
wire n_225;
wire n_1307;
wire n_988;
wire n_814;
wire n_192;
wire n_1549;
wire n_1201;
wire n_1114;
wire n_655;
wire n_1616;
wire n_1446;
wire n_669;
wire n_472;
wire n_1458;
wire n_1176;
wire n_1472;
wire n_387;
wire n_1149;
wire n_398;
wire n_635;
wire n_763;
wire n_1020;
wire n_1062;
wire n_211;
wire n_1219;
wire n_1204;
wire n_178;
wire n_1035;
wire n_287;
wire n_555;
wire n_783;
wire n_1188;
wire n_661;
wire n_849;
wire n_336;
wire n_584;
wire n_681;
wire n_1638;
wire n_430;
wire n_510;
wire n_216;
wire n_311;
wire n_830;
wire n_1296;
wire n_1413;
wire n_801;
wire n_241;
wire n_875;
wire n_357;
wire n_1110;
wire n_1655;
wire n_445;
wire n_749;
wire n_1134;
wire n_1358;
wire n_717;
wire n_165;
wire n_939;
wire n_482;
wire n_1088;
wire n_588;
wire n_1173;
wire n_789;
wire n_1232;
wire n_1603;
wire n_734;
wire n_638;
wire n_866;
wire n_969;
wire n_1401;
wire n_1019;
wire n_1105;
wire n_249;
wire n_304;
wire n_1338;
wire n_577;
wire n_1522;
wire n_1637;
wire n_1419;
wire n_338;
wire n_1653;
wire n_693;
wire n_1506;
wire n_836;
wire n_990;
wire n_1389;
wire n_975;
wire n_1256;
wire n_567;
wire n_1465;
wire n_778;
wire n_1122;
wire n_306;
wire n_458;
wire n_770;
wire n_1375;
wire n_1102;
wire n_711;
wire n_1499;
wire n_1187;
wire n_1441;
wire n_1392;
wire n_1597;
wire n_1164;
wire n_1659;
wire n_489;
wire n_1174;
wire n_1371;
wire n_617;
wire n_1303;
wire n_1572;
wire n_876;
wire n_1516;
wire n_1190;
wire n_601;
wire n_917;
wire n_966;
wire n_253;
wire n_1116;
wire n_1212;
wire n_1541;
wire n_206;
wire n_172;
wire n_217;
wire n_726;
wire n_982;
wire n_1573;
wire n_1453;
wire n_818;
wire n_861;
wire n_1183;
wire n_1658;
wire n_899;
wire n_1253;
wire n_210;
wire n_774;
wire n_1628;
wire n_1335;
wire n_1514;
wire n_1059;
wire n_1345;
wire n_176;
wire n_1133;
wire n_557;
wire n_1410;
wire n_1005;
wire n_607;
wire n_1003;
wire n_679;
wire n_710;
wire n_527;
wire n_1168;
wire n_707;
wire n_937;
wire n_1427;
wire n_393;
wire n_487;
wire n_1584;
wire n_665;
wire n_1440;
wire n_177;
wire n_421;
wire n_1356;
wire n_910;
wire n_1657;
wire n_768;
wire n_1475;
wire n_1302;
wire n_205;
wire n_1136;
wire n_1313;
wire n_1491;
wire n_754;
wire n_1496;
wire n_179;
wire n_1125;
wire n_410;
wire n_708;
wire n_529;
wire n_735;
wire n_232;
wire n_1109;
wire n_895;
wire n_1310;
wire n_202;
wire n_427;
wire n_1399;
wire n_1543;
wire n_791;
wire n_732;
wire n_1533;
wire n_193;
wire n_808;
wire n_797;
wire n_1025;
wire n_500;
wire n_1067;
wire n_435;
wire n_159;
wire n_766;
wire n_1457;
wire n_541;
wire n_538;
wire n_1117;
wire n_799;
wire n_687;
wire n_715;
wire n_1480;
wire n_1482;
wire n_1213;
wire n_1266;
wire n_536;
wire n_872;
wire n_594;
wire n_200;
wire n_1291;
wire n_1297;
wire n_1155;
wire n_1418;
wire n_1524;
wire n_1485;
wire n_1011;
wire n_1184;
wire n_985;
wire n_869;
wire n_810;
wire n_416;
wire n_827;
wire n_401;
wire n_1352;
wire n_626;
wire n_1650;
wire n_1144;
wire n_1137;
wire n_1570;
wire n_1170;
wire n_305;
wire n_676;
wire n_294;
wire n_318;
wire n_653;
wire n_642;
wire n_1602;
wire n_194;
wire n_855;
wire n_1178;
wire n_1461;
wire n_850;
wire n_684;
wire n_268;
wire n_664;
wire n_503;
wire n_235;
wire n_1372;
wire n_605;
wire n_1273;
wire n_353;
wire n_620;
wire n_643;
wire n_916;
wire n_1081;
wire n_493;
wire n_1235;
wire n_703;
wire n_698;
wire n_980;
wire n_1115;
wire n_1282;
wire n_1318;
wire n_780;
wire n_998;
wire n_1454;
wire n_467;
wire n_1227;
wire n_1531;
wire n_840;
wire n_1334;
wire n_501;
wire n_823;
wire n_245;
wire n_725;
wire n_1388;
wire n_1417;
wire n_1295;
wire n_672;
wire n_581;
wire n_382;
wire n_554;
wire n_1625;
wire n_898;
wire n_1013;
wire n_1452;
wire n_718;
wire n_265;
wire n_1120;
wire n_719;
wire n_443;
wire n_198;
wire n_714;
wire n_909;
wire n_1497;
wire n_1530;
wire n_997;
wire n_932;
wire n_612;
wire n_1409;
wire n_788;
wire n_1326;
wire n_1268;
wire n_559;
wire n_825;
wire n_508;
wire n_506;
wire n_1320;
wire n_737;
wire n_986;
wire n_509;
wire n_1317;
wire n_1518;
wire n_1281;
wire n_1192;
wire n_1024;
wire n_1063;
wire n_209;
wire n_1564;
wire n_1613;
wire n_733;
wire n_1489;
wire n_1376;
wire n_941;
wire n_981;
wire n_1569;
wire n_867;
wire n_186;
wire n_587;
wire n_792;
wire n_756;
wire n_1429;
wire n_399;
wire n_1238;
wire n_548;
wire n_812;
wire n_298;
wire n_518;
wire n_505;
wire n_282;
wire n_752;
wire n_905;
wire n_1476;
wire n_1108;
wire n_782;
wire n_1100;
wire n_1395;
wire n_862;
wire n_1425;
wire n_760;
wire n_1620;
wire n_381;
wire n_220;
wire n_390;
wire n_1330;
wire n_481;
wire n_1554;
wire n_769;
wire n_1046;
wire n_271;
wire n_934;
wire n_1618;
wire n_826;
wire n_886;
wire n_1221;
wire n_654;
wire n_1172;
wire n_167;
wire n_428;
wire n_379;
wire n_1341;
wire n_570;
wire n_1641;
wire n_1361;
wire n_853;
wire n_377;
wire n_751;
wire n_786;
wire n_1083;
wire n_1142;
wire n_1129;
wire n_392;
wire n_158;
wire n_704;
wire n_787;
wire n_961;
wire n_771;
wire n_276;
wire n_1225;
wire n_1520;
wire n_169;
wire n_522;
wire n_1287;
wire n_1262;
wire n_400;
wire n_930;
wire n_181;
wire n_1411;
wire n_221;
wire n_622;
wire n_1577;
wire n_1087;
wire n_386;
wire n_994;
wire n_848;
wire n_1550;
wire n_1498;
wire n_1223;
wire n_1272;
wire n_682;
wire n_1567;
wire n_1247;
wire n_922;
wire n_816;
wire n_1648;
wire n_591;
wire n_1536;
wire n_1344;
wire n_313;
wire n_631;
wire n_479;
wire n_1246;
wire n_1478;
wire n_1339;
wire n_432;
wire n_839;
wire n_1210;
wire n_1364;
wire n_328;
wire n_1250;
wire n_369;
wire n_871;
wire n_598;
wire n_685;
wire n_928;
wire n_608;
wire n_1367;
wire n_1460;
wire n_772;
wire n_1555;
wire n_499;
wire n_1589;
wire n_517;
wire n_413;
wire n_402;
wire n_1086;
wire n_796;
wire n_1619;
wire n_236;
wire n_1502;
wire n_1469;
wire n_1012;
wire n_1396;
wire n_1348;
wire n_903;
wire n_1525;
wire n_740;
wire n_203;
wire n_384;
wire n_1404;
wire n_1315;
wire n_277;
wire n_1061;
wire n_333;
wire n_1298;
wire n_1652;
wire n_462;
wire n_1193;
wire n_1255;
wire n_258;
wire n_1113;
wire n_1226;
wire n_722;
wire n_1277;
wire n_188;
wire n_844;
wire n_201;
wire n_471;
wire n_852;
wire n_1487;
wire n_1028;
wire n_1601;
wire n_781;
wire n_474;
wire n_542;
wire n_463;
wire n_1546;
wire n_595;
wire n_502;
wire n_466;
wire n_420;
wire n_1337;
wire n_1495;
wire n_632;
wire n_699;
wire n_979;
wire n_1515;
wire n_1627;
wire n_1245;
wire n_846;
wire n_465;
wire n_362;
wire n_1321;
wire n_170;
wire n_161;
wire n_273;
wire n_585;
wire n_270;
wire n_616;
wire n_745;
wire n_1654;
wire n_1103;
wire n_648;
wire n_1379;
wire n_312;
wire n_1076;
wire n_1091;
wire n_1408;
wire n_494;
wire n_641;
wire n_730;
wire n_1325;
wire n_1595;
wire n_354;
wire n_575;
wire n_480;
wire n_425;
wire n_795;
wire n_695;
wire n_180;
wire n_656;
wire n_1606;
wire n_1220;
wire n_1540;
wire n_229;
wire n_437;
wire n_1642;
wire n_403;
wire n_453;
wire n_1130;
wire n_720;
wire n_1526;
wire n_863;
wire n_805;
wire n_1604;
wire n_1275;
wire n_712;
wire n_246;
wire n_1583;
wire n_1042;
wire n_1402;
wire n_269;
wire n_285;
wire n_412;
wire n_1493;
wire n_657;
wire n_644;
wire n_1160;
wire n_1397;
wire n_491;
wire n_1258;
wire n_1074;
wire n_1621;
wire n_251;
wire n_160;
wire n_566;
wire n_565;
wire n_1448;
wire n_1507;
wire n_1398;
wire n_597;
wire n_1181;
wire n_1505;
wire n_1634;
wire n_1196;
wire n_651;
wire n_1340;
wire n_334;
wire n_811;
wire n_1558;
wire n_807;
wire n_835;
wire n_175;
wire n_666;
wire n_262;
wire n_1433;
wire n_1254;
wire n_1026;
wire n_1234;
wire n_319;
wire n_364;
wire n_1138;
wire n_927;
wire n_1089;
wire n_1004;
wire n_1186;
wire n_1032;
wire n_242;
wire n_1018;
wire n_438;
wire n_713;
wire n_904;
wire n_1588;
wire n_1622;
wire n_166;
wire n_1180;
wire n_1271;
wire n_533;
wire n_1542;
wire n_1251;
wire n_278;

BUFx10_ASAP7_75t_L g154 ( 
.A(n_109),
.Y(n_154)
);

CKINVDCx5p33_ASAP7_75t_R g155 ( 
.A(n_104),
.Y(n_155)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_131),
.Y(n_156)
);

CKINVDCx5p33_ASAP7_75t_R g157 ( 
.A(n_150),
.Y(n_157)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_61),
.Y(n_158)
);

CKINVDCx5p33_ASAP7_75t_R g159 ( 
.A(n_84),
.Y(n_159)
);

CKINVDCx5p33_ASAP7_75t_R g160 ( 
.A(n_29),
.Y(n_160)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_143),
.Y(n_161)
);

CKINVDCx5p33_ASAP7_75t_R g162 ( 
.A(n_75),
.Y(n_162)
);

BUFx2_ASAP7_75t_L g163 ( 
.A(n_135),
.Y(n_163)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_106),
.Y(n_164)
);

INVx2_ASAP7_75t_SL g165 ( 
.A(n_87),
.Y(n_165)
);

CKINVDCx5p33_ASAP7_75t_R g166 ( 
.A(n_132),
.Y(n_166)
);

CKINVDCx5p33_ASAP7_75t_R g167 ( 
.A(n_39),
.Y(n_167)
);

CKINVDCx14_ASAP7_75t_R g168 ( 
.A(n_120),
.Y(n_168)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_27),
.Y(n_169)
);

BUFx10_ASAP7_75t_L g170 ( 
.A(n_38),
.Y(n_170)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_97),
.Y(n_171)
);

CKINVDCx5p33_ASAP7_75t_R g172 ( 
.A(n_58),
.Y(n_172)
);

CKINVDCx5p33_ASAP7_75t_R g173 ( 
.A(n_9),
.Y(n_173)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_153),
.Y(n_174)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_79),
.Y(n_175)
);

BUFx10_ASAP7_75t_L g176 ( 
.A(n_43),
.Y(n_176)
);

CKINVDCx5p33_ASAP7_75t_R g177 ( 
.A(n_134),
.Y(n_177)
);

BUFx2_ASAP7_75t_L g178 ( 
.A(n_43),
.Y(n_178)
);

INVx2_ASAP7_75t_L g179 ( 
.A(n_12),
.Y(n_179)
);

CKINVDCx5p33_ASAP7_75t_R g180 ( 
.A(n_21),
.Y(n_180)
);

CKINVDCx14_ASAP7_75t_R g181 ( 
.A(n_81),
.Y(n_181)
);

CKINVDCx5p33_ASAP7_75t_R g182 ( 
.A(n_86),
.Y(n_182)
);

CKINVDCx5p33_ASAP7_75t_R g183 ( 
.A(n_98),
.Y(n_183)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_68),
.Y(n_184)
);

INVx2_ASAP7_75t_L g185 ( 
.A(n_6),
.Y(n_185)
);

INVx1_ASAP7_75t_SL g186 ( 
.A(n_46),
.Y(n_186)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_63),
.Y(n_187)
);

INVx1_ASAP7_75t_SL g188 ( 
.A(n_50),
.Y(n_188)
);

CKINVDCx5p33_ASAP7_75t_R g189 ( 
.A(n_74),
.Y(n_189)
);

INVx1_ASAP7_75t_SL g190 ( 
.A(n_93),
.Y(n_190)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_4),
.Y(n_191)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_56),
.Y(n_192)
);

BUFx2_ASAP7_75t_SL g193 ( 
.A(n_59),
.Y(n_193)
);

CKINVDCx5p33_ASAP7_75t_R g194 ( 
.A(n_57),
.Y(n_194)
);

BUFx8_ASAP7_75t_SL g195 ( 
.A(n_39),
.Y(n_195)
);

CKINVDCx5p33_ASAP7_75t_R g196 ( 
.A(n_85),
.Y(n_196)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_112),
.Y(n_197)
);

INVx2_ASAP7_75t_L g198 ( 
.A(n_78),
.Y(n_198)
);

CKINVDCx5p33_ASAP7_75t_R g199 ( 
.A(n_105),
.Y(n_199)
);

BUFx6f_ASAP7_75t_L g200 ( 
.A(n_71),
.Y(n_200)
);

CKINVDCx5p33_ASAP7_75t_R g201 ( 
.A(n_5),
.Y(n_201)
);

INVx2_ASAP7_75t_L g202 ( 
.A(n_14),
.Y(n_202)
);

CKINVDCx5p33_ASAP7_75t_R g203 ( 
.A(n_13),
.Y(n_203)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_10),
.Y(n_204)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_89),
.Y(n_205)
);

INVxp67_ASAP7_75t_L g206 ( 
.A(n_45),
.Y(n_206)
);

CKINVDCx5p33_ASAP7_75t_R g207 ( 
.A(n_88),
.Y(n_207)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_141),
.Y(n_208)
);

CKINVDCx5p33_ASAP7_75t_R g209 ( 
.A(n_10),
.Y(n_209)
);

INVx2_ASAP7_75t_L g210 ( 
.A(n_91),
.Y(n_210)
);

CKINVDCx5p33_ASAP7_75t_R g211 ( 
.A(n_46),
.Y(n_211)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_62),
.Y(n_212)
);

CKINVDCx5p33_ASAP7_75t_R g213 ( 
.A(n_44),
.Y(n_213)
);

CKINVDCx5p33_ASAP7_75t_R g214 ( 
.A(n_52),
.Y(n_214)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_139),
.Y(n_215)
);

BUFx3_ASAP7_75t_L g216 ( 
.A(n_142),
.Y(n_216)
);

CKINVDCx5p33_ASAP7_75t_R g217 ( 
.A(n_42),
.Y(n_217)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_15),
.Y(n_218)
);

CKINVDCx5p33_ASAP7_75t_R g219 ( 
.A(n_7),
.Y(n_219)
);

CKINVDCx20_ASAP7_75t_R g220 ( 
.A(n_64),
.Y(n_220)
);

CKINVDCx5p33_ASAP7_75t_R g221 ( 
.A(n_11),
.Y(n_221)
);

CKINVDCx20_ASAP7_75t_R g222 ( 
.A(n_144),
.Y(n_222)
);

CKINVDCx5p33_ASAP7_75t_R g223 ( 
.A(n_9),
.Y(n_223)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_49),
.Y(n_224)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_48),
.Y(n_225)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_65),
.Y(n_226)
);

CKINVDCx5p33_ASAP7_75t_R g227 ( 
.A(n_130),
.Y(n_227)
);

INVx2_ASAP7_75t_SL g228 ( 
.A(n_70),
.Y(n_228)
);

CKINVDCx20_ASAP7_75t_R g229 ( 
.A(n_60),
.Y(n_229)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_138),
.Y(n_230)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_123),
.Y(n_231)
);

CKINVDCx5p33_ASAP7_75t_R g232 ( 
.A(n_99),
.Y(n_232)
);

CKINVDCx5p33_ASAP7_75t_R g233 ( 
.A(n_102),
.Y(n_233)
);

CKINVDCx5p33_ASAP7_75t_R g234 ( 
.A(n_145),
.Y(n_234)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_3),
.Y(n_235)
);

BUFx3_ASAP7_75t_L g236 ( 
.A(n_111),
.Y(n_236)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_77),
.Y(n_237)
);

CKINVDCx5p33_ASAP7_75t_R g238 ( 
.A(n_121),
.Y(n_238)
);

CKINVDCx5p33_ASAP7_75t_R g239 ( 
.A(n_129),
.Y(n_239)
);

CKINVDCx5p33_ASAP7_75t_R g240 ( 
.A(n_80),
.Y(n_240)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_14),
.Y(n_241)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_16),
.Y(n_242)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_19),
.Y(n_243)
);

CKINVDCx5p33_ASAP7_75t_R g244 ( 
.A(n_31),
.Y(n_244)
);

CKINVDCx5p33_ASAP7_75t_R g245 ( 
.A(n_76),
.Y(n_245)
);

CKINVDCx5p33_ASAP7_75t_R g246 ( 
.A(n_90),
.Y(n_246)
);

CKINVDCx5p33_ASAP7_75t_R g247 ( 
.A(n_94),
.Y(n_247)
);

BUFx3_ASAP7_75t_L g248 ( 
.A(n_8),
.Y(n_248)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_11),
.Y(n_249)
);

CKINVDCx5p33_ASAP7_75t_R g250 ( 
.A(n_152),
.Y(n_250)
);

CKINVDCx5p33_ASAP7_75t_R g251 ( 
.A(n_2),
.Y(n_251)
);

CKINVDCx5p33_ASAP7_75t_R g252 ( 
.A(n_25),
.Y(n_252)
);

CKINVDCx20_ASAP7_75t_R g253 ( 
.A(n_22),
.Y(n_253)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_18),
.Y(n_254)
);

INVx2_ASAP7_75t_L g255 ( 
.A(n_100),
.Y(n_255)
);

BUFx3_ASAP7_75t_L g256 ( 
.A(n_117),
.Y(n_256)
);

CKINVDCx5p33_ASAP7_75t_R g257 ( 
.A(n_47),
.Y(n_257)
);

CKINVDCx5p33_ASAP7_75t_R g258 ( 
.A(n_54),
.Y(n_258)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_32),
.Y(n_259)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_95),
.Y(n_260)
);

INVx2_ASAP7_75t_L g261 ( 
.A(n_33),
.Y(n_261)
);

CKINVDCx5p33_ASAP7_75t_R g262 ( 
.A(n_125),
.Y(n_262)
);

CKINVDCx5p33_ASAP7_75t_R g263 ( 
.A(n_37),
.Y(n_263)
);

CKINVDCx5p33_ASAP7_75t_R g264 ( 
.A(n_4),
.Y(n_264)
);

CKINVDCx5p33_ASAP7_75t_R g265 ( 
.A(n_137),
.Y(n_265)
);

CKINVDCx5p33_ASAP7_75t_R g266 ( 
.A(n_119),
.Y(n_266)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_110),
.Y(n_267)
);

CKINVDCx5p33_ASAP7_75t_R g268 ( 
.A(n_149),
.Y(n_268)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_25),
.Y(n_269)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_151),
.Y(n_270)
);

BUFx10_ASAP7_75t_L g271 ( 
.A(n_27),
.Y(n_271)
);

CKINVDCx5p33_ASAP7_75t_R g272 ( 
.A(n_5),
.Y(n_272)
);

CKINVDCx20_ASAP7_75t_R g273 ( 
.A(n_136),
.Y(n_273)
);

CKINVDCx5p33_ASAP7_75t_R g274 ( 
.A(n_22),
.Y(n_274)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_69),
.Y(n_275)
);

CKINVDCx5p33_ASAP7_75t_R g276 ( 
.A(n_146),
.Y(n_276)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_35),
.Y(n_277)
);

BUFx10_ASAP7_75t_L g278 ( 
.A(n_16),
.Y(n_278)
);

CKINVDCx5p33_ASAP7_75t_R g279 ( 
.A(n_128),
.Y(n_279)
);

CKINVDCx5p33_ASAP7_75t_R g280 ( 
.A(n_148),
.Y(n_280)
);

CKINVDCx5p33_ASAP7_75t_R g281 ( 
.A(n_126),
.Y(n_281)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_51),
.Y(n_282)
);

CKINVDCx5p33_ASAP7_75t_R g283 ( 
.A(n_33),
.Y(n_283)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_118),
.Y(n_284)
);

INVx2_ASAP7_75t_SL g285 ( 
.A(n_24),
.Y(n_285)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_72),
.Y(n_286)
);

CKINVDCx5p33_ASAP7_75t_R g287 ( 
.A(n_20),
.Y(n_287)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_36),
.Y(n_288)
);

INVx2_ASAP7_75t_SL g289 ( 
.A(n_28),
.Y(n_289)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_32),
.Y(n_290)
);

CKINVDCx5p33_ASAP7_75t_R g291 ( 
.A(n_17),
.Y(n_291)
);

INVx2_ASAP7_75t_SL g292 ( 
.A(n_114),
.Y(n_292)
);

CKINVDCx5p33_ASAP7_75t_R g293 ( 
.A(n_19),
.Y(n_293)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_83),
.Y(n_294)
);

CKINVDCx5p33_ASAP7_75t_R g295 ( 
.A(n_73),
.Y(n_295)
);

BUFx6f_ASAP7_75t_L g296 ( 
.A(n_42),
.Y(n_296)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_82),
.Y(n_297)
);

CKINVDCx5p33_ASAP7_75t_R g298 ( 
.A(n_24),
.Y(n_298)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_29),
.Y(n_299)
);

INVx1_ASAP7_75t_SL g300 ( 
.A(n_55),
.Y(n_300)
);

CKINVDCx5p33_ASAP7_75t_R g301 ( 
.A(n_195),
.Y(n_301)
);

INVxp67_ASAP7_75t_SL g302 ( 
.A(n_163),
.Y(n_302)
);

CKINVDCx20_ASAP7_75t_R g303 ( 
.A(n_220),
.Y(n_303)
);

INVx2_ASAP7_75t_L g304 ( 
.A(n_200),
.Y(n_304)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_296),
.Y(n_305)
);

INVx2_ASAP7_75t_L g306 ( 
.A(n_200),
.Y(n_306)
);

CKINVDCx5p33_ASAP7_75t_R g307 ( 
.A(n_189),
.Y(n_307)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_296),
.Y(n_308)
);

INVx2_ASAP7_75t_L g309 ( 
.A(n_200),
.Y(n_309)
);

INVxp67_ASAP7_75t_L g310 ( 
.A(n_178),
.Y(n_310)
);

CKINVDCx16_ASAP7_75t_R g311 ( 
.A(n_168),
.Y(n_311)
);

CKINVDCx5p33_ASAP7_75t_R g312 ( 
.A(n_194),
.Y(n_312)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_296),
.Y(n_313)
);

INVxp67_ASAP7_75t_SL g314 ( 
.A(n_216),
.Y(n_314)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_296),
.Y(n_315)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_296),
.Y(n_316)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_179),
.Y(n_317)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_179),
.Y(n_318)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_185),
.Y(n_319)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_185),
.Y(n_320)
);

CKINVDCx20_ASAP7_75t_R g321 ( 
.A(n_222),
.Y(n_321)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_202),
.Y(n_322)
);

INVxp33_ASAP7_75t_SL g323 ( 
.A(n_160),
.Y(n_323)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_202),
.Y(n_324)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_261),
.Y(n_325)
);

INVxp67_ASAP7_75t_SL g326 ( 
.A(n_216),
.Y(n_326)
);

CKINVDCx5p33_ASAP7_75t_R g327 ( 
.A(n_196),
.Y(n_327)
);

CKINVDCx16_ASAP7_75t_R g328 ( 
.A(n_181),
.Y(n_328)
);

CKINVDCx16_ASAP7_75t_R g329 ( 
.A(n_154),
.Y(n_329)
);

INVx2_ASAP7_75t_L g330 ( 
.A(n_261),
.Y(n_330)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_248),
.Y(n_331)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_248),
.Y(n_332)
);

INVxp67_ASAP7_75t_SL g333 ( 
.A(n_236),
.Y(n_333)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_169),
.Y(n_334)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_191),
.Y(n_335)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_204),
.Y(n_336)
);

CKINVDCx16_ASAP7_75t_R g337 ( 
.A(n_154),
.Y(n_337)
);

INVx1_ASAP7_75t_L g338 ( 
.A(n_218),
.Y(n_338)
);

CKINVDCx5p33_ASAP7_75t_R g339 ( 
.A(n_199),
.Y(n_339)
);

CKINVDCx5p33_ASAP7_75t_R g340 ( 
.A(n_207),
.Y(n_340)
);

HB1xp67_ASAP7_75t_L g341 ( 
.A(n_160),
.Y(n_341)
);

INVx1_ASAP7_75t_L g342 ( 
.A(n_235),
.Y(n_342)
);

INVx2_ASAP7_75t_L g343 ( 
.A(n_200),
.Y(n_343)
);

INVx1_ASAP7_75t_L g344 ( 
.A(n_241),
.Y(n_344)
);

INVx1_ASAP7_75t_L g345 ( 
.A(n_242),
.Y(n_345)
);

INVx1_ASAP7_75t_L g346 ( 
.A(n_243),
.Y(n_346)
);

INVx1_ASAP7_75t_L g347 ( 
.A(n_249),
.Y(n_347)
);

BUFx2_ASAP7_75t_L g348 ( 
.A(n_167),
.Y(n_348)
);

INVxp67_ASAP7_75t_SL g349 ( 
.A(n_236),
.Y(n_349)
);

INVxp67_ASAP7_75t_L g350 ( 
.A(n_170),
.Y(n_350)
);

INVxp67_ASAP7_75t_SL g351 ( 
.A(n_256),
.Y(n_351)
);

INVx1_ASAP7_75t_L g352 ( 
.A(n_254),
.Y(n_352)
);

INVx1_ASAP7_75t_L g353 ( 
.A(n_259),
.Y(n_353)
);

CKINVDCx5p33_ASAP7_75t_R g354 ( 
.A(n_227),
.Y(n_354)
);

CKINVDCx20_ASAP7_75t_R g355 ( 
.A(n_229),
.Y(n_355)
);

INVxp67_ASAP7_75t_SL g356 ( 
.A(n_256),
.Y(n_356)
);

INVxp67_ASAP7_75t_SL g357 ( 
.A(n_156),
.Y(n_357)
);

INVx1_ASAP7_75t_L g358 ( 
.A(n_269),
.Y(n_358)
);

CKINVDCx5p33_ASAP7_75t_R g359 ( 
.A(n_232),
.Y(n_359)
);

INVx1_ASAP7_75t_L g360 ( 
.A(n_277),
.Y(n_360)
);

INVx1_ASAP7_75t_L g361 ( 
.A(n_288),
.Y(n_361)
);

INVx1_ASAP7_75t_L g362 ( 
.A(n_290),
.Y(n_362)
);

INVx1_ASAP7_75t_L g363 ( 
.A(n_299),
.Y(n_363)
);

CKINVDCx20_ASAP7_75t_R g364 ( 
.A(n_273),
.Y(n_364)
);

BUFx3_ASAP7_75t_L g365 ( 
.A(n_158),
.Y(n_365)
);

INVx1_ASAP7_75t_L g366 ( 
.A(n_285),
.Y(n_366)
);

INVxp67_ASAP7_75t_SL g367 ( 
.A(n_161),
.Y(n_367)
);

INVxp67_ASAP7_75t_L g368 ( 
.A(n_170),
.Y(n_368)
);

INVx1_ASAP7_75t_L g369 ( 
.A(n_285),
.Y(n_369)
);

INVx1_ASAP7_75t_L g370 ( 
.A(n_289),
.Y(n_370)
);

CKINVDCx5p33_ASAP7_75t_R g371 ( 
.A(n_233),
.Y(n_371)
);

CKINVDCx5p33_ASAP7_75t_R g372 ( 
.A(n_234),
.Y(n_372)
);

INVx2_ASAP7_75t_L g373 ( 
.A(n_200),
.Y(n_373)
);

AND2x2_ASAP7_75t_L g374 ( 
.A(n_314),
.B(n_289),
.Y(n_374)
);

AND2x4_ASAP7_75t_L g375 ( 
.A(n_365),
.B(n_165),
.Y(n_375)
);

OAI22xp5_ASAP7_75t_SL g376 ( 
.A1(n_329),
.A2(n_253),
.B1(n_298),
.B2(n_173),
.Y(n_376)
);

BUFx6f_ASAP7_75t_L g377 ( 
.A(n_304),
.Y(n_377)
);

NOR2xp33_ASAP7_75t_R g378 ( 
.A(n_307),
.B(n_238),
.Y(n_378)
);

OA21x2_ASAP7_75t_L g379 ( 
.A1(n_304),
.A2(n_210),
.B(n_198),
.Y(n_379)
);

CKINVDCx5p33_ASAP7_75t_R g380 ( 
.A(n_312),
.Y(n_380)
);

INVx1_ASAP7_75t_L g381 ( 
.A(n_305),
.Y(n_381)
);

NAND2xp5_ASAP7_75t_L g382 ( 
.A(n_327),
.B(n_165),
.Y(n_382)
);

CKINVDCx5p33_ASAP7_75t_R g383 ( 
.A(n_339),
.Y(n_383)
);

NAND2xp5_ASAP7_75t_L g384 ( 
.A(n_340),
.B(n_228),
.Y(n_384)
);

INVx1_ASAP7_75t_L g385 ( 
.A(n_305),
.Y(n_385)
);

INVx1_ASAP7_75t_L g386 ( 
.A(n_308),
.Y(n_386)
);

BUFx6f_ASAP7_75t_L g387 ( 
.A(n_304),
.Y(n_387)
);

NOR2xp33_ASAP7_75t_SL g388 ( 
.A(n_329),
.B(n_154),
.Y(n_388)
);

HB1xp67_ASAP7_75t_L g389 ( 
.A(n_341),
.Y(n_389)
);

BUFx6f_ASAP7_75t_L g390 ( 
.A(n_306),
.Y(n_390)
);

INVx1_ASAP7_75t_L g391 ( 
.A(n_308),
.Y(n_391)
);

BUFx8_ASAP7_75t_L g392 ( 
.A(n_348),
.Y(n_392)
);

BUFx6f_ASAP7_75t_L g393 ( 
.A(n_306),
.Y(n_393)
);

OR2x2_ASAP7_75t_L g394 ( 
.A(n_348),
.B(n_186),
.Y(n_394)
);

INVx1_ASAP7_75t_L g395 ( 
.A(n_313),
.Y(n_395)
);

INVx1_ASAP7_75t_L g396 ( 
.A(n_313),
.Y(n_396)
);

INVx1_ASAP7_75t_L g397 ( 
.A(n_315),
.Y(n_397)
);

INVx1_ASAP7_75t_L g398 ( 
.A(n_315),
.Y(n_398)
);

INVx2_ASAP7_75t_L g399 ( 
.A(n_316),
.Y(n_399)
);

BUFx6f_ASAP7_75t_L g400 ( 
.A(n_306),
.Y(n_400)
);

INVx2_ASAP7_75t_L g401 ( 
.A(n_309),
.Y(n_401)
);

INVx2_ASAP7_75t_L g402 ( 
.A(n_309),
.Y(n_402)
);

INVx2_ASAP7_75t_L g403 ( 
.A(n_316),
.Y(n_403)
);

INVx3_ASAP7_75t_L g404 ( 
.A(n_309),
.Y(n_404)
);

BUFx2_ASAP7_75t_L g405 ( 
.A(n_350),
.Y(n_405)
);

NAND2xp5_ASAP7_75t_L g406 ( 
.A(n_354),
.B(n_359),
.Y(n_406)
);

AND2x4_ASAP7_75t_L g407 ( 
.A(n_365),
.B(n_292),
.Y(n_407)
);

INVx3_ASAP7_75t_L g408 ( 
.A(n_343),
.Y(n_408)
);

NAND2xp5_ASAP7_75t_L g409 ( 
.A(n_371),
.B(n_292),
.Y(n_409)
);

INVx1_ASAP7_75t_L g410 ( 
.A(n_330),
.Y(n_410)
);

NOR2xp33_ASAP7_75t_L g411 ( 
.A(n_372),
.B(n_188),
.Y(n_411)
);

INVx1_ASAP7_75t_L g412 ( 
.A(n_330),
.Y(n_412)
);

AND2x4_ASAP7_75t_L g413 ( 
.A(n_365),
.B(n_198),
.Y(n_413)
);

INVx1_ASAP7_75t_L g414 ( 
.A(n_343),
.Y(n_414)
);

AOI22xp5_ASAP7_75t_L g415 ( 
.A1(n_310),
.A2(n_167),
.B1(n_298),
.B2(n_293),
.Y(n_415)
);

BUFx6f_ASAP7_75t_L g416 ( 
.A(n_343),
.Y(n_416)
);

AND2x2_ASAP7_75t_L g417 ( 
.A(n_326),
.B(n_333),
.Y(n_417)
);

INVx1_ASAP7_75t_L g418 ( 
.A(n_373),
.Y(n_418)
);

INVx1_ASAP7_75t_L g419 ( 
.A(n_373),
.Y(n_419)
);

NOR2xp33_ASAP7_75t_R g420 ( 
.A(n_311),
.B(n_239),
.Y(n_420)
);

INVx2_ASAP7_75t_L g421 ( 
.A(n_373),
.Y(n_421)
);

CKINVDCx20_ASAP7_75t_R g422 ( 
.A(n_303),
.Y(n_422)
);

CKINVDCx5p33_ASAP7_75t_R g423 ( 
.A(n_301),
.Y(n_423)
);

BUFx3_ASAP7_75t_L g424 ( 
.A(n_331),
.Y(n_424)
);

AND2x2_ASAP7_75t_SL g425 ( 
.A(n_311),
.B(n_210),
.Y(n_425)
);

INVx1_ASAP7_75t_L g426 ( 
.A(n_334),
.Y(n_426)
);

CKINVDCx5p33_ASAP7_75t_R g427 ( 
.A(n_321),
.Y(n_427)
);

CKINVDCx5p33_ASAP7_75t_R g428 ( 
.A(n_355),
.Y(n_428)
);

INVx1_ASAP7_75t_L g429 ( 
.A(n_334),
.Y(n_429)
);

INVx2_ASAP7_75t_L g430 ( 
.A(n_317),
.Y(n_430)
);

OA21x2_ASAP7_75t_L g431 ( 
.A1(n_317),
.A2(n_255),
.B(n_171),
.Y(n_431)
);

BUFx6f_ASAP7_75t_L g432 ( 
.A(n_318),
.Y(n_432)
);

INVx1_ASAP7_75t_L g433 ( 
.A(n_335),
.Y(n_433)
);

INVx1_ASAP7_75t_L g434 ( 
.A(n_335),
.Y(n_434)
);

INVx1_ASAP7_75t_L g435 ( 
.A(n_336),
.Y(n_435)
);

AND2x2_ASAP7_75t_L g436 ( 
.A(n_349),
.B(n_351),
.Y(n_436)
);

INVx3_ASAP7_75t_L g437 ( 
.A(n_318),
.Y(n_437)
);

INVx1_ASAP7_75t_L g438 ( 
.A(n_336),
.Y(n_438)
);

BUFx6f_ASAP7_75t_L g439 ( 
.A(n_319),
.Y(n_439)
);

BUFx6f_ASAP7_75t_L g440 ( 
.A(n_319),
.Y(n_440)
);

INVx2_ASAP7_75t_L g441 ( 
.A(n_399),
.Y(n_441)
);

NAND2xp5_ASAP7_75t_SL g442 ( 
.A(n_425),
.B(n_337),
.Y(n_442)
);

OAI21xp33_ASAP7_75t_SL g443 ( 
.A1(n_374),
.A2(n_425),
.B(n_302),
.Y(n_443)
);

INVx1_ASAP7_75t_L g444 ( 
.A(n_381),
.Y(n_444)
);

NAND2xp5_ASAP7_75t_SL g445 ( 
.A(n_425),
.B(n_337),
.Y(n_445)
);

INVx2_ASAP7_75t_L g446 ( 
.A(n_399),
.Y(n_446)
);

INVx2_ASAP7_75t_L g447 ( 
.A(n_403),
.Y(n_447)
);

BUFx6f_ASAP7_75t_L g448 ( 
.A(n_377),
.Y(n_448)
);

INVx2_ASAP7_75t_L g449 ( 
.A(n_403),
.Y(n_449)
);

NAND2xp5_ASAP7_75t_SL g450 ( 
.A(n_411),
.B(n_328),
.Y(n_450)
);

CKINVDCx5p33_ASAP7_75t_R g451 ( 
.A(n_427),
.Y(n_451)
);

BUFx3_ASAP7_75t_L g452 ( 
.A(n_424),
.Y(n_452)
);

INVx2_ASAP7_75t_L g453 ( 
.A(n_432),
.Y(n_453)
);

INVx3_ASAP7_75t_L g454 ( 
.A(n_377),
.Y(n_454)
);

AND2x2_ASAP7_75t_L g455 ( 
.A(n_417),
.B(n_356),
.Y(n_455)
);

INVx1_ASAP7_75t_L g456 ( 
.A(n_381),
.Y(n_456)
);

INVx2_ASAP7_75t_L g457 ( 
.A(n_432),
.Y(n_457)
);

AND2x4_ASAP7_75t_L g458 ( 
.A(n_413),
.B(n_255),
.Y(n_458)
);

INVx1_ASAP7_75t_L g459 ( 
.A(n_385),
.Y(n_459)
);

INVx4_ASAP7_75t_L g460 ( 
.A(n_431),
.Y(n_460)
);

NOR2xp33_ASAP7_75t_L g461 ( 
.A(n_382),
.B(n_323),
.Y(n_461)
);

INVx2_ASAP7_75t_L g462 ( 
.A(n_432),
.Y(n_462)
);

INVx3_ASAP7_75t_L g463 ( 
.A(n_377),
.Y(n_463)
);

INVx1_ASAP7_75t_L g464 ( 
.A(n_385),
.Y(n_464)
);

OAI22xp5_ASAP7_75t_L g465 ( 
.A1(n_406),
.A2(n_328),
.B1(n_206),
.B2(n_367),
.Y(n_465)
);

INVx2_ASAP7_75t_L g466 ( 
.A(n_432),
.Y(n_466)
);

NAND2xp5_ASAP7_75t_SL g467 ( 
.A(n_388),
.B(n_368),
.Y(n_467)
);

INVx2_ASAP7_75t_L g468 ( 
.A(n_432),
.Y(n_468)
);

INVx1_ASAP7_75t_L g469 ( 
.A(n_386),
.Y(n_469)
);

INVxp67_ASAP7_75t_L g470 ( 
.A(n_405),
.Y(n_470)
);

BUFx3_ASAP7_75t_L g471 ( 
.A(n_424),
.Y(n_471)
);

OR2x2_ASAP7_75t_L g472 ( 
.A(n_394),
.B(n_331),
.Y(n_472)
);

AOI22xp33_ASAP7_75t_L g473 ( 
.A1(n_374),
.A2(n_357),
.B1(n_193),
.B2(n_332),
.Y(n_473)
);

NAND2xp5_ASAP7_75t_SL g474 ( 
.A(n_420),
.B(n_155),
.Y(n_474)
);

INVx2_ASAP7_75t_L g475 ( 
.A(n_432),
.Y(n_475)
);

CKINVDCx5p33_ASAP7_75t_R g476 ( 
.A(n_428),
.Y(n_476)
);

CKINVDCx5p33_ASAP7_75t_R g477 ( 
.A(n_378),
.Y(n_477)
);

NAND2xp5_ASAP7_75t_SL g478 ( 
.A(n_380),
.B(n_383),
.Y(n_478)
);

INVx2_ASAP7_75t_L g479 ( 
.A(n_439),
.Y(n_479)
);

INVx2_ASAP7_75t_L g480 ( 
.A(n_439),
.Y(n_480)
);

NAND2xp5_ASAP7_75t_L g481 ( 
.A(n_417),
.B(n_190),
.Y(n_481)
);

AOI22xp5_ASAP7_75t_L g482 ( 
.A1(n_376),
.A2(n_180),
.B1(n_173),
.B2(n_221),
.Y(n_482)
);

INVx2_ASAP7_75t_L g483 ( 
.A(n_439),
.Y(n_483)
);

INVx2_ASAP7_75t_L g484 ( 
.A(n_439),
.Y(n_484)
);

NAND2xp5_ASAP7_75t_L g485 ( 
.A(n_436),
.B(n_300),
.Y(n_485)
);

INVx2_ASAP7_75t_L g486 ( 
.A(n_439),
.Y(n_486)
);

INVxp67_ASAP7_75t_SL g487 ( 
.A(n_436),
.Y(n_487)
);

INVxp33_ASAP7_75t_L g488 ( 
.A(n_394),
.Y(n_488)
);

CKINVDCx6p67_ASAP7_75t_R g489 ( 
.A(n_422),
.Y(n_489)
);

OAI22xp33_ASAP7_75t_L g490 ( 
.A1(n_415),
.A2(n_219),
.B1(n_217),
.B2(n_213),
.Y(n_490)
);

INVx3_ASAP7_75t_L g491 ( 
.A(n_377),
.Y(n_491)
);

INVx2_ASAP7_75t_L g492 ( 
.A(n_439),
.Y(n_492)
);

CKINVDCx5p33_ASAP7_75t_R g493 ( 
.A(n_392),
.Y(n_493)
);

INVx2_ASAP7_75t_SL g494 ( 
.A(n_375),
.Y(n_494)
);

INVx2_ASAP7_75t_L g495 ( 
.A(n_440),
.Y(n_495)
);

INVx2_ASAP7_75t_L g496 ( 
.A(n_440),
.Y(n_496)
);

NOR2xp33_ASAP7_75t_L g497 ( 
.A(n_384),
.B(n_409),
.Y(n_497)
);

INVx2_ASAP7_75t_SL g498 ( 
.A(n_375),
.Y(n_498)
);

INVx1_ASAP7_75t_L g499 ( 
.A(n_386),
.Y(n_499)
);

INVx2_ASAP7_75t_L g500 ( 
.A(n_440),
.Y(n_500)
);

INVx1_ASAP7_75t_L g501 ( 
.A(n_391),
.Y(n_501)
);

NAND2xp5_ASAP7_75t_SL g502 ( 
.A(n_405),
.B(n_157),
.Y(n_502)
);

NAND2xp5_ASAP7_75t_L g503 ( 
.A(n_375),
.B(n_240),
.Y(n_503)
);

INVx2_ASAP7_75t_L g504 ( 
.A(n_440),
.Y(n_504)
);

INVx5_ASAP7_75t_L g505 ( 
.A(n_377),
.Y(n_505)
);

NAND2xp5_ASAP7_75t_SL g506 ( 
.A(n_415),
.B(n_159),
.Y(n_506)
);

INVx2_ASAP7_75t_L g507 ( 
.A(n_440),
.Y(n_507)
);

INVx2_ASAP7_75t_L g508 ( 
.A(n_440),
.Y(n_508)
);

INVx1_ASAP7_75t_L g509 ( 
.A(n_391),
.Y(n_509)
);

AOI22xp5_ASAP7_75t_L g510 ( 
.A1(n_389),
.A2(n_251),
.B1(n_180),
.B2(n_221),
.Y(n_510)
);

OAI22xp33_ASAP7_75t_L g511 ( 
.A1(n_424),
.A2(n_244),
.B1(n_211),
.B2(n_209),
.Y(n_511)
);

INVx1_ASAP7_75t_L g512 ( 
.A(n_395),
.Y(n_512)
);

NAND2xp5_ASAP7_75t_SL g513 ( 
.A(n_375),
.B(n_407),
.Y(n_513)
);

INVx2_ASAP7_75t_L g514 ( 
.A(n_395),
.Y(n_514)
);

INVx1_ASAP7_75t_L g515 ( 
.A(n_396),
.Y(n_515)
);

NOR2x1p5_ASAP7_75t_L g516 ( 
.A(n_423),
.B(n_251),
.Y(n_516)
);

INVx2_ASAP7_75t_SL g517 ( 
.A(n_407),
.Y(n_517)
);

INVx1_ASAP7_75t_L g518 ( 
.A(n_396),
.Y(n_518)
);

INVx2_ASAP7_75t_L g519 ( 
.A(n_397),
.Y(n_519)
);

INVx1_ASAP7_75t_L g520 ( 
.A(n_397),
.Y(n_520)
);

INVx1_ASAP7_75t_L g521 ( 
.A(n_398),
.Y(n_521)
);

NAND3xp33_ASAP7_75t_L g522 ( 
.A(n_413),
.B(n_431),
.C(n_407),
.Y(n_522)
);

OA22x2_ASAP7_75t_L g523 ( 
.A1(n_407),
.A2(n_370),
.B1(n_369),
.B2(n_366),
.Y(n_523)
);

INVx3_ASAP7_75t_L g524 ( 
.A(n_377),
.Y(n_524)
);

INVx4_ASAP7_75t_L g525 ( 
.A(n_431),
.Y(n_525)
);

INVx2_ASAP7_75t_SL g526 ( 
.A(n_413),
.Y(n_526)
);

OAI22xp33_ASAP7_75t_L g527 ( 
.A1(n_426),
.A2(n_203),
.B1(n_201),
.B2(n_223),
.Y(n_527)
);

NAND2xp5_ASAP7_75t_SL g528 ( 
.A(n_392),
.B(n_159),
.Y(n_528)
);

INVx1_ASAP7_75t_L g529 ( 
.A(n_398),
.Y(n_529)
);

INVx3_ASAP7_75t_L g530 ( 
.A(n_387),
.Y(n_530)
);

NOR2xp33_ASAP7_75t_L g531 ( 
.A(n_429),
.B(n_332),
.Y(n_531)
);

INVx2_ASAP7_75t_L g532 ( 
.A(n_401),
.Y(n_532)
);

INVx1_ASAP7_75t_L g533 ( 
.A(n_431),
.Y(n_533)
);

NAND3xp33_ASAP7_75t_L g534 ( 
.A(n_413),
.B(n_338),
.C(n_363),
.Y(n_534)
);

NOR2xp33_ASAP7_75t_L g535 ( 
.A(n_429),
.B(n_364),
.Y(n_535)
);

INVx2_ASAP7_75t_L g536 ( 
.A(n_401),
.Y(n_536)
);

NOR2xp33_ASAP7_75t_L g537 ( 
.A(n_433),
.B(n_366),
.Y(n_537)
);

INVx1_ASAP7_75t_L g538 ( 
.A(n_433),
.Y(n_538)
);

NAND2xp5_ASAP7_75t_SL g539 ( 
.A(n_392),
.B(n_162),
.Y(n_539)
);

INVx1_ASAP7_75t_L g540 ( 
.A(n_434),
.Y(n_540)
);

INVx2_ASAP7_75t_L g541 ( 
.A(n_401),
.Y(n_541)
);

INVx2_ASAP7_75t_L g542 ( 
.A(n_402),
.Y(n_542)
);

INVx2_ASAP7_75t_L g543 ( 
.A(n_402),
.Y(n_543)
);

INVx2_ASAP7_75t_L g544 ( 
.A(n_402),
.Y(n_544)
);

INVx1_ASAP7_75t_L g545 ( 
.A(n_434),
.Y(n_545)
);

CKINVDCx11_ASAP7_75t_R g546 ( 
.A(n_392),
.Y(n_546)
);

INVx2_ASAP7_75t_L g547 ( 
.A(n_421),
.Y(n_547)
);

BUFx2_ASAP7_75t_L g548 ( 
.A(n_435),
.Y(n_548)
);

INVx1_ASAP7_75t_L g549 ( 
.A(n_435),
.Y(n_549)
);

NOR2xp33_ASAP7_75t_L g550 ( 
.A(n_438),
.B(n_369),
.Y(n_550)
);

INVxp67_ASAP7_75t_SL g551 ( 
.A(n_387),
.Y(n_551)
);

INVx2_ASAP7_75t_L g552 ( 
.A(n_421),
.Y(n_552)
);

INVx1_ASAP7_75t_L g553 ( 
.A(n_438),
.Y(n_553)
);

INVx3_ASAP7_75t_L g554 ( 
.A(n_387),
.Y(n_554)
);

AOI22xp33_ASAP7_75t_L g555 ( 
.A1(n_379),
.A2(n_338),
.B1(n_363),
.B2(n_362),
.Y(n_555)
);

INVx2_ASAP7_75t_L g556 ( 
.A(n_421),
.Y(n_556)
);

INVx1_ASAP7_75t_L g557 ( 
.A(n_414),
.Y(n_557)
);

INVx2_ASAP7_75t_L g558 ( 
.A(n_414),
.Y(n_558)
);

NAND2xp33_ASAP7_75t_L g559 ( 
.A(n_387),
.B(n_162),
.Y(n_559)
);

BUFx6f_ASAP7_75t_L g560 ( 
.A(n_387),
.Y(n_560)
);

INVx2_ASAP7_75t_SL g561 ( 
.A(n_379),
.Y(n_561)
);

OAI22xp33_ASAP7_75t_L g562 ( 
.A1(n_430),
.A2(n_291),
.B1(n_283),
.B2(n_287),
.Y(n_562)
);

OAI21xp33_ASAP7_75t_SL g563 ( 
.A1(n_410),
.A2(n_370),
.B(n_362),
.Y(n_563)
);

NOR2xp33_ASAP7_75t_L g564 ( 
.A(n_430),
.B(n_166),
.Y(n_564)
);

INVx2_ASAP7_75t_L g565 ( 
.A(n_418),
.Y(n_565)
);

INVx2_ASAP7_75t_L g566 ( 
.A(n_418),
.Y(n_566)
);

INVx2_ASAP7_75t_L g567 ( 
.A(n_419),
.Y(n_567)
);

INVx1_ASAP7_75t_L g568 ( 
.A(n_379),
.Y(n_568)
);

BUFx6f_ASAP7_75t_L g569 ( 
.A(n_387),
.Y(n_569)
);

INVx1_ASAP7_75t_L g570 ( 
.A(n_379),
.Y(n_570)
);

INVx2_ASAP7_75t_L g571 ( 
.A(n_404),
.Y(n_571)
);

NAND2xp5_ASAP7_75t_SL g572 ( 
.A(n_437),
.B(n_166),
.Y(n_572)
);

INVx2_ASAP7_75t_L g573 ( 
.A(n_404),
.Y(n_573)
);

INVx3_ASAP7_75t_L g574 ( 
.A(n_390),
.Y(n_574)
);

INVx1_ASAP7_75t_L g575 ( 
.A(n_410),
.Y(n_575)
);

INVx2_ASAP7_75t_L g576 ( 
.A(n_404),
.Y(n_576)
);

CKINVDCx5p33_ASAP7_75t_R g577 ( 
.A(n_437),
.Y(n_577)
);

NAND2xp33_ASAP7_75t_SL g578 ( 
.A(n_437),
.B(n_252),
.Y(n_578)
);

NAND2xp5_ASAP7_75t_L g579 ( 
.A(n_437),
.B(n_245),
.Y(n_579)
);

NAND2xp5_ASAP7_75t_SL g580 ( 
.A(n_412),
.B(n_172),
.Y(n_580)
);

INVx1_ASAP7_75t_L g581 ( 
.A(n_412),
.Y(n_581)
);

INVx2_ASAP7_75t_L g582 ( 
.A(n_404),
.Y(n_582)
);

INVx2_ASAP7_75t_SL g583 ( 
.A(n_416),
.Y(n_583)
);

NAND2xp5_ASAP7_75t_L g584 ( 
.A(n_408),
.B(n_390),
.Y(n_584)
);

INVx1_ASAP7_75t_L g585 ( 
.A(n_408),
.Y(n_585)
);

INVx2_ASAP7_75t_L g586 ( 
.A(n_408),
.Y(n_586)
);

INVx1_ASAP7_75t_L g587 ( 
.A(n_526),
.Y(n_587)
);

INVx2_ASAP7_75t_L g588 ( 
.A(n_514),
.Y(n_588)
);

INVx4_ASAP7_75t_L g589 ( 
.A(n_452),
.Y(n_589)
);

NAND2xp33_ASAP7_75t_SL g590 ( 
.A(n_488),
.B(n_252),
.Y(n_590)
);

NAND2xp5_ASAP7_75t_SL g591 ( 
.A(n_494),
.B(n_164),
.Y(n_591)
);

INVx1_ASAP7_75t_L g592 ( 
.A(n_526),
.Y(n_592)
);

INVx1_ASAP7_75t_L g593 ( 
.A(n_538),
.Y(n_593)
);

INVx1_ASAP7_75t_L g594 ( 
.A(n_538),
.Y(n_594)
);

BUFx5_ASAP7_75t_L g595 ( 
.A(n_568),
.Y(n_595)
);

INVx2_ASAP7_75t_L g596 ( 
.A(n_514),
.Y(n_596)
);

NAND2xp5_ASAP7_75t_SL g597 ( 
.A(n_494),
.B(n_174),
.Y(n_597)
);

INVx1_ASAP7_75t_L g598 ( 
.A(n_540),
.Y(n_598)
);

INVx2_ASAP7_75t_L g599 ( 
.A(n_519),
.Y(n_599)
);

NOR2xp33_ASAP7_75t_L g600 ( 
.A(n_497),
.B(n_172),
.Y(n_600)
);

NAND2xp5_ASAP7_75t_L g601 ( 
.A(n_498),
.B(n_175),
.Y(n_601)
);

NAND2xp5_ASAP7_75t_L g602 ( 
.A(n_498),
.B(n_517),
.Y(n_602)
);

INVx1_ASAP7_75t_L g603 ( 
.A(n_545),
.Y(n_603)
);

BUFx6f_ASAP7_75t_L g604 ( 
.A(n_452),
.Y(n_604)
);

INVx1_ASAP7_75t_L g605 ( 
.A(n_545),
.Y(n_605)
);

INVx2_ASAP7_75t_L g606 ( 
.A(n_519),
.Y(n_606)
);

AOI22xp5_ASAP7_75t_L g607 ( 
.A1(n_443),
.A2(n_281),
.B1(n_279),
.B2(n_246),
.Y(n_607)
);

NAND2xp5_ASAP7_75t_SL g608 ( 
.A(n_517),
.B(n_184),
.Y(n_608)
);

INVx2_ASAP7_75t_L g609 ( 
.A(n_571),
.Y(n_609)
);

NAND2xp5_ASAP7_75t_SL g610 ( 
.A(n_443),
.B(n_187),
.Y(n_610)
);

BUFx6f_ASAP7_75t_L g611 ( 
.A(n_452),
.Y(n_611)
);

INVx2_ASAP7_75t_L g612 ( 
.A(n_571),
.Y(n_612)
);

BUFx6f_ASAP7_75t_SL g613 ( 
.A(n_546),
.Y(n_613)
);

NAND2xp5_ASAP7_75t_SL g614 ( 
.A(n_577),
.B(n_192),
.Y(n_614)
);

NAND2xp5_ASAP7_75t_L g615 ( 
.A(n_487),
.B(n_197),
.Y(n_615)
);

NAND2xp5_ASAP7_75t_SL g616 ( 
.A(n_577),
.B(n_205),
.Y(n_616)
);

NAND2xp5_ASAP7_75t_L g617 ( 
.A(n_513),
.B(n_208),
.Y(n_617)
);

NAND2xp5_ASAP7_75t_L g618 ( 
.A(n_455),
.B(n_212),
.Y(n_618)
);

NOR2xp33_ASAP7_75t_L g619 ( 
.A(n_461),
.B(n_177),
.Y(n_619)
);

NAND2xp5_ASAP7_75t_L g620 ( 
.A(n_455),
.B(n_215),
.Y(n_620)
);

AOI21xp5_ASAP7_75t_L g621 ( 
.A1(n_561),
.A2(n_416),
.B(n_400),
.Y(n_621)
);

INVx3_ASAP7_75t_L g622 ( 
.A(n_471),
.Y(n_622)
);

AND2x2_ASAP7_75t_L g623 ( 
.A(n_548),
.B(n_170),
.Y(n_623)
);

AOI22xp5_ASAP7_75t_L g624 ( 
.A1(n_442),
.A2(n_214),
.B1(n_183),
.B2(n_182),
.Y(n_624)
);

INVx1_ASAP7_75t_L g625 ( 
.A(n_549),
.Y(n_625)
);

NOR2xp33_ASAP7_75t_L g626 ( 
.A(n_481),
.B(n_177),
.Y(n_626)
);

INVxp67_ASAP7_75t_L g627 ( 
.A(n_535),
.Y(n_627)
);

NAND2xp5_ASAP7_75t_L g628 ( 
.A(n_549),
.B(n_224),
.Y(n_628)
);

INVxp67_ASAP7_75t_L g629 ( 
.A(n_472),
.Y(n_629)
);

AND2x2_ASAP7_75t_L g630 ( 
.A(n_548),
.B(n_176),
.Y(n_630)
);

INVx2_ASAP7_75t_L g631 ( 
.A(n_573),
.Y(n_631)
);

INVx3_ASAP7_75t_L g632 ( 
.A(n_471),
.Y(n_632)
);

AOI22xp33_ASAP7_75t_L g633 ( 
.A1(n_522),
.A2(n_231),
.B1(n_237),
.B2(n_230),
.Y(n_633)
);

INVx1_ASAP7_75t_L g634 ( 
.A(n_553),
.Y(n_634)
);

NOR2xp33_ASAP7_75t_L g635 ( 
.A(n_485),
.B(n_182),
.Y(n_635)
);

AOI22xp33_ASAP7_75t_L g636 ( 
.A1(n_522),
.A2(n_260),
.B1(n_275),
.B2(n_270),
.Y(n_636)
);

INVx2_ASAP7_75t_L g637 ( 
.A(n_573),
.Y(n_637)
);

INVx2_ASAP7_75t_L g638 ( 
.A(n_576),
.Y(n_638)
);

BUFx3_ASAP7_75t_L g639 ( 
.A(n_471),
.Y(n_639)
);

NAND2xp5_ASAP7_75t_L g640 ( 
.A(n_561),
.B(n_533),
.Y(n_640)
);

INVx2_ASAP7_75t_L g641 ( 
.A(n_576),
.Y(n_641)
);

INVx1_ASAP7_75t_L g642 ( 
.A(n_444),
.Y(n_642)
);

NOR2xp33_ASAP7_75t_L g643 ( 
.A(n_472),
.B(n_445),
.Y(n_643)
);

INVx1_ASAP7_75t_L g644 ( 
.A(n_444),
.Y(n_644)
);

INVx3_ASAP7_75t_L g645 ( 
.A(n_460),
.Y(n_645)
);

NAND2xp5_ASAP7_75t_L g646 ( 
.A(n_533),
.B(n_225),
.Y(n_646)
);

NAND2xp5_ASAP7_75t_L g647 ( 
.A(n_458),
.B(n_226),
.Y(n_647)
);

NAND2xp5_ASAP7_75t_L g648 ( 
.A(n_458),
.B(n_267),
.Y(n_648)
);

INVx2_ASAP7_75t_SL g649 ( 
.A(n_523),
.Y(n_649)
);

NAND2xp5_ASAP7_75t_SL g650 ( 
.A(n_460),
.B(n_282),
.Y(n_650)
);

NAND2xp5_ASAP7_75t_L g651 ( 
.A(n_458),
.B(n_284),
.Y(n_651)
);

NAND2xp33_ASAP7_75t_L g652 ( 
.A(n_503),
.B(n_183),
.Y(n_652)
);

INVx1_ASAP7_75t_L g653 ( 
.A(n_456),
.Y(n_653)
);

INVxp67_ASAP7_75t_L g654 ( 
.A(n_502),
.Y(n_654)
);

INVx1_ASAP7_75t_L g655 ( 
.A(n_456),
.Y(n_655)
);

NAND2xp33_ASAP7_75t_L g656 ( 
.A(n_555),
.B(n_214),
.Y(n_656)
);

OR2x2_ASAP7_75t_L g657 ( 
.A(n_470),
.B(n_342),
.Y(n_657)
);

INVxp67_ASAP7_75t_L g658 ( 
.A(n_467),
.Y(n_658)
);

A2O1A1Ixp33_ASAP7_75t_L g659 ( 
.A1(n_563),
.A2(n_531),
.B(n_550),
.C(n_537),
.Y(n_659)
);

NAND2xp5_ASAP7_75t_L g660 ( 
.A(n_458),
.B(n_286),
.Y(n_660)
);

NAND2xp5_ASAP7_75t_SL g661 ( 
.A(n_460),
.B(n_294),
.Y(n_661)
);

NAND2xp33_ASAP7_75t_L g662 ( 
.A(n_568),
.B(n_247),
.Y(n_662)
);

NOR2xp67_ASAP7_75t_L g663 ( 
.A(n_477),
.B(n_250),
.Y(n_663)
);

BUFx8_ASAP7_75t_L g664 ( 
.A(n_489),
.Y(n_664)
);

NOR3xp33_ASAP7_75t_L g665 ( 
.A(n_506),
.B(n_347),
.C(n_342),
.Y(n_665)
);

NAND2xp5_ASAP7_75t_SL g666 ( 
.A(n_460),
.B(n_297),
.Y(n_666)
);

AOI22xp33_ASAP7_75t_L g667 ( 
.A1(n_525),
.A2(n_523),
.B1(n_570),
.B2(n_534),
.Y(n_667)
);

AO22x2_ASAP7_75t_L g668 ( 
.A1(n_465),
.A2(n_352),
.B1(n_361),
.B2(n_360),
.Y(n_668)
);

AND2x2_ASAP7_75t_L g669 ( 
.A(n_450),
.B(n_176),
.Y(n_669)
);

NAND2xp5_ASAP7_75t_SL g670 ( 
.A(n_525),
.B(n_250),
.Y(n_670)
);

NAND2xp5_ASAP7_75t_L g671 ( 
.A(n_570),
.B(n_390),
.Y(n_671)
);

INVx1_ASAP7_75t_L g672 ( 
.A(n_459),
.Y(n_672)
);

NAND2xp5_ASAP7_75t_L g673 ( 
.A(n_459),
.B(n_390),
.Y(n_673)
);

AND2x2_ASAP7_75t_L g674 ( 
.A(n_510),
.B(n_176),
.Y(n_674)
);

INVx2_ASAP7_75t_L g675 ( 
.A(n_582),
.Y(n_675)
);

AND2x2_ASAP7_75t_L g676 ( 
.A(n_510),
.B(n_271),
.Y(n_676)
);

NAND2xp5_ASAP7_75t_L g677 ( 
.A(n_464),
.B(n_390),
.Y(n_677)
);

NAND2xp5_ASAP7_75t_SL g678 ( 
.A(n_525),
.B(n_579),
.Y(n_678)
);

NAND2xp5_ASAP7_75t_L g679 ( 
.A(n_464),
.B(n_390),
.Y(n_679)
);

NAND2xp5_ASAP7_75t_L g680 ( 
.A(n_469),
.B(n_393),
.Y(n_680)
);

INVx4_ASAP7_75t_L g681 ( 
.A(n_448),
.Y(n_681)
);

INVx2_ASAP7_75t_L g682 ( 
.A(n_575),
.Y(n_682)
);

AND2x2_ASAP7_75t_L g683 ( 
.A(n_473),
.B(n_271),
.Y(n_683)
);

INVx2_ASAP7_75t_SL g684 ( 
.A(n_523),
.Y(n_684)
);

NAND2xp5_ASAP7_75t_L g685 ( 
.A(n_469),
.B(n_393),
.Y(n_685)
);

AOI221xp5_ASAP7_75t_L g686 ( 
.A1(n_490),
.A2(n_293),
.B1(n_263),
.B2(n_264),
.C(n_272),
.Y(n_686)
);

A2O1A1Ixp33_ASAP7_75t_L g687 ( 
.A1(n_563),
.A2(n_347),
.B(n_344),
.C(n_345),
.Y(n_687)
);

AOI22xp33_ASAP7_75t_L g688 ( 
.A1(n_525),
.A2(n_263),
.B1(n_264),
.B2(n_274),
.Y(n_688)
);

NAND2xp5_ASAP7_75t_SL g689 ( 
.A(n_499),
.B(n_257),
.Y(n_689)
);

AOI22xp5_ASAP7_75t_L g690 ( 
.A1(n_572),
.A2(n_257),
.B1(n_258),
.B2(n_262),
.Y(n_690)
);

INVx1_ASAP7_75t_L g691 ( 
.A(n_499),
.Y(n_691)
);

NAND2xp5_ASAP7_75t_L g692 ( 
.A(n_501),
.B(n_393),
.Y(n_692)
);

NOR2xp67_ASAP7_75t_L g693 ( 
.A(n_478),
.B(n_258),
.Y(n_693)
);

INVx1_ASAP7_75t_L g694 ( 
.A(n_501),
.Y(n_694)
);

INVxp67_ASAP7_75t_L g695 ( 
.A(n_578),
.Y(n_695)
);

BUFx6f_ASAP7_75t_SL g696 ( 
.A(n_489),
.Y(n_696)
);

INVx2_ASAP7_75t_L g697 ( 
.A(n_586),
.Y(n_697)
);

INVxp67_ASAP7_75t_L g698 ( 
.A(n_580),
.Y(n_698)
);

NAND2xp5_ASAP7_75t_L g699 ( 
.A(n_509),
.B(n_393),
.Y(n_699)
);

AOI21xp5_ASAP7_75t_L g700 ( 
.A1(n_551),
.A2(n_416),
.B(n_400),
.Y(n_700)
);

NAND2xp5_ASAP7_75t_L g701 ( 
.A(n_509),
.B(n_393),
.Y(n_701)
);

INVx1_ASAP7_75t_SL g702 ( 
.A(n_451),
.Y(n_702)
);

INVx1_ASAP7_75t_L g703 ( 
.A(n_512),
.Y(n_703)
);

NAND2xp5_ASAP7_75t_L g704 ( 
.A(n_512),
.B(n_393),
.Y(n_704)
);

NOR2xp33_ASAP7_75t_L g705 ( 
.A(n_474),
.B(n_262),
.Y(n_705)
);

NAND2xp5_ASAP7_75t_L g706 ( 
.A(n_515),
.B(n_400),
.Y(n_706)
);

NAND2xp5_ASAP7_75t_L g707 ( 
.A(n_515),
.B(n_400),
.Y(n_707)
);

NAND2xp5_ASAP7_75t_L g708 ( 
.A(n_518),
.B(n_400),
.Y(n_708)
);

NAND2xp5_ASAP7_75t_L g709 ( 
.A(n_518),
.B(n_400),
.Y(n_709)
);

NAND2xp5_ASAP7_75t_L g710 ( 
.A(n_520),
.B(n_416),
.Y(n_710)
);

AOI22xp33_ASAP7_75t_L g711 ( 
.A1(n_534),
.A2(n_278),
.B1(n_271),
.B2(n_361),
.Y(n_711)
);

INVx1_ASAP7_75t_L g712 ( 
.A(n_520),
.Y(n_712)
);

NOR2xp33_ASAP7_75t_L g713 ( 
.A(n_511),
.B(n_265),
.Y(n_713)
);

AND2x2_ASAP7_75t_L g714 ( 
.A(n_516),
.B(n_278),
.Y(n_714)
);

INVx1_ASAP7_75t_L g715 ( 
.A(n_521),
.Y(n_715)
);

NAND2xp5_ASAP7_75t_L g716 ( 
.A(n_521),
.B(n_416),
.Y(n_716)
);

INVx2_ASAP7_75t_L g717 ( 
.A(n_575),
.Y(n_717)
);

INVx1_ASAP7_75t_L g718 ( 
.A(n_529),
.Y(n_718)
);

NAND2xp5_ASAP7_75t_SL g719 ( 
.A(n_529),
.B(n_265),
.Y(n_719)
);

NAND2xp5_ASAP7_75t_L g720 ( 
.A(n_564),
.B(n_416),
.Y(n_720)
);

NAND2xp5_ASAP7_75t_SL g721 ( 
.A(n_453),
.B(n_266),
.Y(n_721)
);

NOR2xp33_ASAP7_75t_L g722 ( 
.A(n_527),
.B(n_266),
.Y(n_722)
);

CKINVDCx20_ASAP7_75t_R g723 ( 
.A(n_451),
.Y(n_723)
);

CKINVDCx5p33_ASAP7_75t_R g724 ( 
.A(n_476),
.Y(n_724)
);

INVx1_ASAP7_75t_L g725 ( 
.A(n_581),
.Y(n_725)
);

INVx1_ASAP7_75t_L g726 ( 
.A(n_581),
.Y(n_726)
);

INVx1_ASAP7_75t_L g727 ( 
.A(n_557),
.Y(n_727)
);

AOI22xp33_ASAP7_75t_L g728 ( 
.A1(n_557),
.A2(n_278),
.B1(n_360),
.B2(n_358),
.Y(n_728)
);

NOR2xp33_ASAP7_75t_L g729 ( 
.A(n_562),
.B(n_268),
.Y(n_729)
);

NAND2xp5_ASAP7_75t_L g730 ( 
.A(n_583),
.B(n_268),
.Y(n_730)
);

INVx1_ASAP7_75t_L g731 ( 
.A(n_558),
.Y(n_731)
);

INVx2_ASAP7_75t_SL g732 ( 
.A(n_516),
.Y(n_732)
);

INVx2_ASAP7_75t_SL g733 ( 
.A(n_476),
.Y(n_733)
);

INVx2_ASAP7_75t_SL g734 ( 
.A(n_528),
.Y(n_734)
);

NOR2xp33_ASAP7_75t_L g735 ( 
.A(n_539),
.B(n_276),
.Y(n_735)
);

NAND2xp5_ASAP7_75t_L g736 ( 
.A(n_583),
.B(n_454),
.Y(n_736)
);

NAND2xp5_ASAP7_75t_L g737 ( 
.A(n_454),
.B(n_276),
.Y(n_737)
);

INVx2_ASAP7_75t_L g738 ( 
.A(n_558),
.Y(n_738)
);

BUFx6f_ASAP7_75t_SL g739 ( 
.A(n_493),
.Y(n_739)
);

BUFx6f_ASAP7_75t_L g740 ( 
.A(n_448),
.Y(n_740)
);

NAND2xp5_ASAP7_75t_L g741 ( 
.A(n_454),
.B(n_280),
.Y(n_741)
);

NAND2xp5_ASAP7_75t_L g742 ( 
.A(n_454),
.B(n_280),
.Y(n_742)
);

INVx2_ASAP7_75t_L g743 ( 
.A(n_532),
.Y(n_743)
);

INVx2_ASAP7_75t_L g744 ( 
.A(n_565),
.Y(n_744)
);

INVx1_ASAP7_75t_L g745 ( 
.A(n_565),
.Y(n_745)
);

AOI22xp5_ASAP7_75t_L g746 ( 
.A1(n_559),
.A2(n_295),
.B1(n_353),
.B2(n_352),
.Y(n_746)
);

NOR3xp33_ASAP7_75t_L g747 ( 
.A(n_482),
.B(n_358),
.C(n_353),
.Y(n_747)
);

NAND2xp5_ASAP7_75t_L g748 ( 
.A(n_463),
.B(n_295),
.Y(n_748)
);

OAI22xp5_ASAP7_75t_SL g749 ( 
.A1(n_723),
.A2(n_482),
.B1(n_493),
.B2(n_345),
.Y(n_749)
);

AOI22xp33_ASAP7_75t_L g750 ( 
.A1(n_649),
.A2(n_684),
.B1(n_600),
.B2(n_610),
.Y(n_750)
);

OAI22xp5_ASAP7_75t_L g751 ( 
.A1(n_633),
.A2(n_344),
.B1(n_346),
.B2(n_320),
.Y(n_751)
);

INVx5_ASAP7_75t_L g752 ( 
.A(n_645),
.Y(n_752)
);

BUFx6f_ASAP7_75t_L g753 ( 
.A(n_604),
.Y(n_753)
);

AOI211xp5_ASAP7_75t_L g754 ( 
.A1(n_619),
.A2(n_346),
.B(n_325),
.C(n_324),
.Y(n_754)
);

INVx1_ASAP7_75t_L g755 ( 
.A(n_682),
.Y(n_755)
);

AND2x4_ASAP7_75t_L g756 ( 
.A(n_639),
.B(n_453),
.Y(n_756)
);

BUFx6f_ASAP7_75t_L g757 ( 
.A(n_604),
.Y(n_757)
);

INVx5_ASAP7_75t_L g758 ( 
.A(n_645),
.Y(n_758)
);

NAND2xp33_ASAP7_75t_L g759 ( 
.A(n_595),
.B(n_448),
.Y(n_759)
);

NOR2xp33_ASAP7_75t_L g760 ( 
.A(n_627),
.B(n_524),
.Y(n_760)
);

INVx1_ASAP7_75t_L g761 ( 
.A(n_717),
.Y(n_761)
);

INVx3_ASAP7_75t_L g762 ( 
.A(n_604),
.Y(n_762)
);

INVxp67_ASAP7_75t_SL g763 ( 
.A(n_622),
.Y(n_763)
);

AOI22xp5_ASAP7_75t_L g764 ( 
.A1(n_619),
.A2(n_500),
.B1(n_457),
.B2(n_496),
.Y(n_764)
);

INVx2_ASAP7_75t_L g765 ( 
.A(n_738),
.Y(n_765)
);

NAND2xp5_ASAP7_75t_L g766 ( 
.A(n_595),
.B(n_640),
.Y(n_766)
);

INVx2_ASAP7_75t_L g767 ( 
.A(n_738),
.Y(n_767)
);

NAND2xp5_ASAP7_75t_L g768 ( 
.A(n_595),
.B(n_457),
.Y(n_768)
);

NAND2xp5_ASAP7_75t_L g769 ( 
.A(n_595),
.B(n_462),
.Y(n_769)
);

O2A1O1Ixp33_ASAP7_75t_L g770 ( 
.A1(n_659),
.A2(n_567),
.B(n_566),
.C(n_441),
.Y(n_770)
);

NAND2x1p5_ASAP7_75t_L g771 ( 
.A(n_589),
.B(n_463),
.Y(n_771)
);

INVx5_ASAP7_75t_L g772 ( 
.A(n_740),
.Y(n_772)
);

INVx2_ASAP7_75t_L g773 ( 
.A(n_744),
.Y(n_773)
);

AND2x4_ASAP7_75t_L g774 ( 
.A(n_639),
.B(n_462),
.Y(n_774)
);

NOR2xp33_ASAP7_75t_L g775 ( 
.A(n_600),
.B(n_524),
.Y(n_775)
);

INVx1_ASAP7_75t_L g776 ( 
.A(n_588),
.Y(n_776)
);

AOI22xp33_ASAP7_75t_L g777 ( 
.A1(n_610),
.A2(n_446),
.B1(n_447),
.B2(n_449),
.Y(n_777)
);

INVx1_ASAP7_75t_L g778 ( 
.A(n_588),
.Y(n_778)
);

NOR2xp33_ASAP7_75t_L g779 ( 
.A(n_654),
.B(n_524),
.Y(n_779)
);

OAI21xp5_ASAP7_75t_L g780 ( 
.A1(n_667),
.A2(n_584),
.B(n_504),
.Y(n_780)
);

NOR2xp67_ASAP7_75t_L g781 ( 
.A(n_724),
.B(n_733),
.Y(n_781)
);

CKINVDCx5p33_ASAP7_75t_R g782 ( 
.A(n_696),
.Y(n_782)
);

O2A1O1Ixp33_ASAP7_75t_L g783 ( 
.A1(n_659),
.A2(n_567),
.B(n_566),
.C(n_449),
.Y(n_783)
);

INVx1_ASAP7_75t_L g784 ( 
.A(n_596),
.Y(n_784)
);

AND2x4_ASAP7_75t_L g785 ( 
.A(n_732),
.B(n_466),
.Y(n_785)
);

AND2x6_ASAP7_75t_SL g786 ( 
.A(n_722),
.B(n_322),
.Y(n_786)
);

BUFx4f_ASAP7_75t_L g787 ( 
.A(n_734),
.Y(n_787)
);

INVx4_ASAP7_75t_L g788 ( 
.A(n_604),
.Y(n_788)
);

INVx1_ASAP7_75t_L g789 ( 
.A(n_596),
.Y(n_789)
);

BUFx8_ASAP7_75t_L g790 ( 
.A(n_696),
.Y(n_790)
);

NOR2xp33_ASAP7_75t_L g791 ( 
.A(n_629),
.B(n_530),
.Y(n_791)
);

INVx1_ASAP7_75t_L g792 ( 
.A(n_599),
.Y(n_792)
);

BUFx3_ASAP7_75t_L g793 ( 
.A(n_664),
.Y(n_793)
);

NAND2xp5_ASAP7_75t_L g794 ( 
.A(n_595),
.B(n_468),
.Y(n_794)
);

NAND2xp5_ASAP7_75t_L g795 ( 
.A(n_595),
.B(n_468),
.Y(n_795)
);

BUFx3_ASAP7_75t_L g796 ( 
.A(n_664),
.Y(n_796)
);

INVx1_ASAP7_75t_L g797 ( 
.A(n_606),
.Y(n_797)
);

NAND2xp33_ASAP7_75t_L g798 ( 
.A(n_633),
.B(n_448),
.Y(n_798)
);

INVx1_ASAP7_75t_L g799 ( 
.A(n_727),
.Y(n_799)
);

NAND2x1p5_ASAP7_75t_L g800 ( 
.A(n_589),
.B(n_611),
.Y(n_800)
);

INVx2_ASAP7_75t_SL g801 ( 
.A(n_657),
.Y(n_801)
);

INVx2_ASAP7_75t_SL g802 ( 
.A(n_623),
.Y(n_802)
);

INVx1_ASAP7_75t_L g803 ( 
.A(n_725),
.Y(n_803)
);

NAND2xp5_ASAP7_75t_L g804 ( 
.A(n_636),
.B(n_475),
.Y(n_804)
);

NAND2xp5_ASAP7_75t_SL g805 ( 
.A(n_643),
.B(n_479),
.Y(n_805)
);

INVx2_ASAP7_75t_SL g806 ( 
.A(n_630),
.Y(n_806)
);

NAND2xp5_ASAP7_75t_L g807 ( 
.A(n_636),
.B(n_593),
.Y(n_807)
);

NAND2xp5_ASAP7_75t_L g808 ( 
.A(n_594),
.B(n_479),
.Y(n_808)
);

INVx1_ASAP7_75t_L g809 ( 
.A(n_726),
.Y(n_809)
);

BUFx6f_ASAP7_75t_L g810 ( 
.A(n_611),
.Y(n_810)
);

INVx1_ASAP7_75t_L g811 ( 
.A(n_598),
.Y(n_811)
);

INVx2_ASAP7_75t_L g812 ( 
.A(n_609),
.Y(n_812)
);

BUFx2_ASAP7_75t_L g813 ( 
.A(n_695),
.Y(n_813)
);

AOI22xp33_ASAP7_75t_L g814 ( 
.A1(n_643),
.A2(n_447),
.B1(n_446),
.B2(n_507),
.Y(n_814)
);

AOI22xp33_ASAP7_75t_L g815 ( 
.A1(n_729),
.A2(n_507),
.B1(n_480),
.B2(n_483),
.Y(n_815)
);

BUFx6f_ASAP7_75t_L g816 ( 
.A(n_611),
.Y(n_816)
);

NAND2xp5_ASAP7_75t_L g817 ( 
.A(n_603),
.B(n_480),
.Y(n_817)
);

NOR2xp33_ASAP7_75t_L g818 ( 
.A(n_658),
.B(n_626),
.Y(n_818)
);

AOI22xp5_ASAP7_75t_L g819 ( 
.A1(n_626),
.A2(n_635),
.B1(n_607),
.B2(n_592),
.Y(n_819)
);

NAND2xp5_ASAP7_75t_L g820 ( 
.A(n_605),
.B(n_625),
.Y(n_820)
);

NAND2xp5_ASAP7_75t_SL g821 ( 
.A(n_635),
.B(n_483),
.Y(n_821)
);

INVx2_ASAP7_75t_SL g822 ( 
.A(n_669),
.Y(n_822)
);

HB1xp67_ASAP7_75t_L g823 ( 
.A(n_634),
.Y(n_823)
);

INVx3_ASAP7_75t_L g824 ( 
.A(n_611),
.Y(n_824)
);

INVx1_ASAP7_75t_L g825 ( 
.A(n_642),
.Y(n_825)
);

INVx3_ASAP7_75t_L g826 ( 
.A(n_622),
.Y(n_826)
);

NAND2xp5_ASAP7_75t_L g827 ( 
.A(n_644),
.B(n_484),
.Y(n_827)
);

INVx3_ASAP7_75t_L g828 ( 
.A(n_632),
.Y(n_828)
);

AOI21x1_ASAP7_75t_L g829 ( 
.A1(n_678),
.A2(n_508),
.B(n_484),
.Y(n_829)
);

AND2x2_ASAP7_75t_L g830 ( 
.A(n_674),
.B(n_322),
.Y(n_830)
);

INVx1_ASAP7_75t_L g831 ( 
.A(n_653),
.Y(n_831)
);

HB1xp67_ASAP7_75t_L g832 ( 
.A(n_655),
.Y(n_832)
);

INVx2_ASAP7_75t_L g833 ( 
.A(n_612),
.Y(n_833)
);

AND2x2_ASAP7_75t_L g834 ( 
.A(n_676),
.B(n_325),
.Y(n_834)
);

NAND2xp5_ASAP7_75t_SL g835 ( 
.A(n_618),
.B(n_486),
.Y(n_835)
);

AND2x2_ASAP7_75t_L g836 ( 
.A(n_683),
.B(n_486),
.Y(n_836)
);

INVx2_ASAP7_75t_L g837 ( 
.A(n_631),
.Y(n_837)
);

BUFx6f_ASAP7_75t_L g838 ( 
.A(n_740),
.Y(n_838)
);

HB1xp67_ASAP7_75t_L g839 ( 
.A(n_672),
.Y(n_839)
);

INVxp67_ASAP7_75t_L g840 ( 
.A(n_590),
.Y(n_840)
);

INVx1_ASAP7_75t_L g841 ( 
.A(n_691),
.Y(n_841)
);

NAND2xp5_ASAP7_75t_L g842 ( 
.A(n_694),
.B(n_492),
.Y(n_842)
);

AND2x6_ASAP7_75t_SL g843 ( 
.A(n_722),
.B(n_0),
.Y(n_843)
);

INVx1_ASAP7_75t_L g844 ( 
.A(n_703),
.Y(n_844)
);

AOI22xp5_ASAP7_75t_L g845 ( 
.A1(n_587),
.A2(n_495),
.B1(n_508),
.B2(n_504),
.Y(n_845)
);

INVx4_ASAP7_75t_L g846 ( 
.A(n_740),
.Y(n_846)
);

NAND2xp33_ASAP7_75t_SL g847 ( 
.A(n_714),
.B(n_739),
.Y(n_847)
);

INVx1_ASAP7_75t_SL g848 ( 
.A(n_702),
.Y(n_848)
);

OAI22xp33_ASAP7_75t_L g849 ( 
.A1(n_620),
.A2(n_500),
.B1(n_496),
.B2(n_495),
.Y(n_849)
);

INVx1_ASAP7_75t_L g850 ( 
.A(n_712),
.Y(n_850)
);

INVx2_ASAP7_75t_L g851 ( 
.A(n_637),
.Y(n_851)
);

NAND2xp5_ASAP7_75t_L g852 ( 
.A(n_715),
.B(n_492),
.Y(n_852)
);

OAI21xp33_ASAP7_75t_L g853 ( 
.A1(n_688),
.A2(n_585),
.B(n_544),
.Y(n_853)
);

BUFx4f_ASAP7_75t_L g854 ( 
.A(n_718),
.Y(n_854)
);

NAND2xp5_ASAP7_75t_L g855 ( 
.A(n_667),
.B(n_463),
.Y(n_855)
);

INVx2_ASAP7_75t_SL g856 ( 
.A(n_668),
.Y(n_856)
);

NAND2xp5_ASAP7_75t_L g857 ( 
.A(n_615),
.B(n_463),
.Y(n_857)
);

BUFx8_ASAP7_75t_L g858 ( 
.A(n_613),
.Y(n_858)
);

NAND2xp5_ASAP7_75t_L g859 ( 
.A(n_632),
.B(n_574),
.Y(n_859)
);

NOR2xp33_ASAP7_75t_L g860 ( 
.A(n_698),
.B(n_530),
.Y(n_860)
);

NAND2xp5_ASAP7_75t_L g861 ( 
.A(n_646),
.B(n_574),
.Y(n_861)
);

AOI22xp5_ASAP7_75t_L g862 ( 
.A1(n_670),
.A2(n_530),
.B1(n_491),
.B2(n_574),
.Y(n_862)
);

INVx3_ASAP7_75t_L g863 ( 
.A(n_740),
.Y(n_863)
);

INVx1_ASAP7_75t_L g864 ( 
.A(n_731),
.Y(n_864)
);

INVx8_ASAP7_75t_L g865 ( 
.A(n_739),
.Y(n_865)
);

OAI21xp5_ASAP7_75t_L g866 ( 
.A1(n_678),
.A2(n_543),
.B(n_536),
.Y(n_866)
);

INVx4_ASAP7_75t_L g867 ( 
.A(n_681),
.Y(n_867)
);

OR2x6_ASAP7_75t_L g868 ( 
.A(n_668),
.B(n_569),
.Y(n_868)
);

NAND2xp5_ASAP7_75t_L g869 ( 
.A(n_671),
.B(n_554),
.Y(n_869)
);

NOR2x1_ASAP7_75t_L g870 ( 
.A(n_663),
.B(n_554),
.Y(n_870)
);

NAND2xp5_ASAP7_75t_SL g871 ( 
.A(n_705),
.B(n_569),
.Y(n_871)
);

INVx2_ASAP7_75t_SL g872 ( 
.A(n_668),
.Y(n_872)
);

OAI22xp33_ASAP7_75t_L g873 ( 
.A1(n_602),
.A2(n_554),
.B1(n_491),
.B2(n_556),
.Y(n_873)
);

INVx1_ASAP7_75t_L g874 ( 
.A(n_745),
.Y(n_874)
);

INVx2_ASAP7_75t_L g875 ( 
.A(n_638),
.Y(n_875)
);

NAND2xp5_ASAP7_75t_SL g876 ( 
.A(n_705),
.B(n_569),
.Y(n_876)
);

INVx2_ASAP7_75t_SL g877 ( 
.A(n_689),
.Y(n_877)
);

AOI22xp33_ASAP7_75t_L g878 ( 
.A1(n_729),
.A2(n_554),
.B1(n_491),
.B2(n_556),
.Y(n_878)
);

CKINVDCx5p33_ASAP7_75t_R g879 ( 
.A(n_613),
.Y(n_879)
);

A2O1A1Ixp33_ASAP7_75t_L g880 ( 
.A1(n_713),
.A2(n_543),
.B(n_536),
.C(n_552),
.Y(n_880)
);

OR2x6_ASAP7_75t_L g881 ( 
.A(n_693),
.B(n_569),
.Y(n_881)
);

INVx2_ASAP7_75t_L g882 ( 
.A(n_641),
.Y(n_882)
);

INVx1_ASAP7_75t_L g883 ( 
.A(n_675),
.Y(n_883)
);

NAND2xp5_ASAP7_75t_L g884 ( 
.A(n_650),
.B(n_542),
.Y(n_884)
);

NAND2xp5_ASAP7_75t_L g885 ( 
.A(n_650),
.B(n_542),
.Y(n_885)
);

AND2x4_ASAP7_75t_L g886 ( 
.A(n_665),
.B(n_560),
.Y(n_886)
);

NAND2xp33_ASAP7_75t_L g887 ( 
.A(n_647),
.B(n_560),
.Y(n_887)
);

HB1xp67_ASAP7_75t_L g888 ( 
.A(n_721),
.Y(n_888)
);

INVx3_ASAP7_75t_L g889 ( 
.A(n_681),
.Y(n_889)
);

INVx2_ASAP7_75t_SL g890 ( 
.A(n_719),
.Y(n_890)
);

AOI22xp5_ASAP7_75t_L g891 ( 
.A1(n_670),
.A2(n_560),
.B1(n_448),
.B2(n_547),
.Y(n_891)
);

INVx3_ASAP7_75t_L g892 ( 
.A(n_697),
.Y(n_892)
);

NAND2xp5_ASAP7_75t_L g893 ( 
.A(n_661),
.B(n_552),
.Y(n_893)
);

INVx2_ASAP7_75t_SL g894 ( 
.A(n_719),
.Y(n_894)
);

NAND2xp5_ASAP7_75t_SL g895 ( 
.A(n_735),
.B(n_560),
.Y(n_895)
);

HB1xp67_ASAP7_75t_L g896 ( 
.A(n_721),
.Y(n_896)
);

NAND2xp5_ASAP7_75t_L g897 ( 
.A(n_661),
.B(n_547),
.Y(n_897)
);

AND2x4_ASAP7_75t_L g898 ( 
.A(n_747),
.B(n_614),
.Y(n_898)
);

NAND2xp5_ASAP7_75t_SL g899 ( 
.A(n_735),
.B(n_560),
.Y(n_899)
);

NAND2xp5_ASAP7_75t_L g900 ( 
.A(n_666),
.B(n_688),
.Y(n_900)
);

INVxp67_ASAP7_75t_L g901 ( 
.A(n_624),
.Y(n_901)
);

INVx1_ASAP7_75t_L g902 ( 
.A(n_673),
.Y(n_902)
);

NAND2xp5_ASAP7_75t_SL g903 ( 
.A(n_614),
.B(n_541),
.Y(n_903)
);

OAI22xp5_ASAP7_75t_SL g904 ( 
.A1(n_711),
.A2(n_0),
.B1(n_1),
.B2(n_6),
.Y(n_904)
);

NAND2xp5_ASAP7_75t_L g905 ( 
.A(n_666),
.B(n_544),
.Y(n_905)
);

NAND2xp5_ASAP7_75t_L g906 ( 
.A(n_628),
.B(n_541),
.Y(n_906)
);

INVx1_ASAP7_75t_L g907 ( 
.A(n_677),
.Y(n_907)
);

INVx1_ASAP7_75t_L g908 ( 
.A(n_679),
.Y(n_908)
);

NAND2xp5_ASAP7_75t_L g909 ( 
.A(n_743),
.B(n_505),
.Y(n_909)
);

NOR2xp33_ASAP7_75t_L g910 ( 
.A(n_616),
.B(n_690),
.Y(n_910)
);

AOI22xp5_ASAP7_75t_L g911 ( 
.A1(n_591),
.A2(n_505),
.B1(n_147),
.B2(n_140),
.Y(n_911)
);

AOI22xp5_ASAP7_75t_L g912 ( 
.A1(n_591),
.A2(n_505),
.B1(n_133),
.B2(n_127),
.Y(n_912)
);

INVx1_ASAP7_75t_SL g913 ( 
.A(n_616),
.Y(n_913)
);

NAND2xp5_ASAP7_75t_SL g914 ( 
.A(n_746),
.B(n_505),
.Y(n_914)
);

INVx1_ASAP7_75t_L g915 ( 
.A(n_680),
.Y(n_915)
);

BUFx3_ASAP7_75t_L g916 ( 
.A(n_730),
.Y(n_916)
);

NAND2xp5_ASAP7_75t_SL g917 ( 
.A(n_728),
.B(n_601),
.Y(n_917)
);

AOI21xp5_ASAP7_75t_L g918 ( 
.A1(n_720),
.A2(n_505),
.B(n_124),
.Y(n_918)
);

AO22x1_ASAP7_75t_L g919 ( 
.A1(n_617),
.A2(n_1),
.B1(n_8),
.B2(n_13),
.Y(n_919)
);

BUFx6f_ASAP7_75t_L g920 ( 
.A(n_838),
.Y(n_920)
);

INVx1_ASAP7_75t_L g921 ( 
.A(n_755),
.Y(n_921)
);

OR2x2_ASAP7_75t_L g922 ( 
.A(n_848),
.B(n_648),
.Y(n_922)
);

INVx6_ASAP7_75t_L g923 ( 
.A(n_790),
.Y(n_923)
);

AND2x2_ASAP7_75t_L g924 ( 
.A(n_830),
.B(n_728),
.Y(n_924)
);

NAND2xp5_ASAP7_75t_L g925 ( 
.A(n_818),
.B(n_597),
.Y(n_925)
);

OAI22xp5_ASAP7_75t_L g926 ( 
.A1(n_819),
.A2(n_651),
.B1(n_660),
.B2(n_597),
.Y(n_926)
);

INVx1_ASAP7_75t_L g927 ( 
.A(n_761),
.Y(n_927)
);

AOI21xp5_ASAP7_75t_L g928 ( 
.A1(n_752),
.A2(n_662),
.B(n_621),
.Y(n_928)
);

NOR2xp33_ASAP7_75t_SL g929 ( 
.A(n_781),
.B(n_687),
.Y(n_929)
);

O2A1O1Ixp33_ASAP7_75t_L g930 ( 
.A1(n_910),
.A2(n_652),
.B(n_608),
.C(n_687),
.Y(n_930)
);

NOR2xp33_ASAP7_75t_L g931 ( 
.A(n_901),
.B(n_608),
.Y(n_931)
);

AND2x2_ASAP7_75t_L g932 ( 
.A(n_834),
.B(n_711),
.Y(n_932)
);

NOR2xp33_ASAP7_75t_SL g933 ( 
.A(n_848),
.B(n_748),
.Y(n_933)
);

INVx2_ASAP7_75t_L g934 ( 
.A(n_765),
.Y(n_934)
);

AND2x2_ASAP7_75t_L g935 ( 
.A(n_801),
.B(n_742),
.Y(n_935)
);

BUFx6f_ASAP7_75t_L g936 ( 
.A(n_838),
.Y(n_936)
);

NAND2xp5_ASAP7_75t_SL g937 ( 
.A(n_854),
.B(n_741),
.Y(n_937)
);

OAI22xp5_ASAP7_75t_L g938 ( 
.A1(n_900),
.A2(n_736),
.B1(n_737),
.B2(n_706),
.Y(n_938)
);

OAI22xp5_ASAP7_75t_L g939 ( 
.A1(n_900),
.A2(n_704),
.B1(n_716),
.B2(n_710),
.Y(n_939)
);

NAND2xp5_ASAP7_75t_L g940 ( 
.A(n_836),
.B(n_656),
.Y(n_940)
);

O2A1O1Ixp33_ASAP7_75t_L g941 ( 
.A1(n_917),
.A2(n_701),
.B(n_709),
.C(n_708),
.Y(n_941)
);

INVx2_ASAP7_75t_L g942 ( 
.A(n_767),
.Y(n_942)
);

NAND3xp33_ASAP7_75t_SL g943 ( 
.A(n_913),
.B(n_707),
.C(n_699),
.Y(n_943)
);

CKINVDCx5p33_ASAP7_75t_R g944 ( 
.A(n_790),
.Y(n_944)
);

AOI21xp5_ASAP7_75t_L g945 ( 
.A1(n_752),
.A2(n_700),
.B(n_692),
.Y(n_945)
);

BUFx6f_ASAP7_75t_L g946 ( 
.A(n_838),
.Y(n_946)
);

NOR2xp33_ASAP7_75t_L g947 ( 
.A(n_913),
.B(n_685),
.Y(n_947)
);

INVxp67_ASAP7_75t_L g948 ( 
.A(n_813),
.Y(n_948)
);

INVx1_ASAP7_75t_L g949 ( 
.A(n_799),
.Y(n_949)
);

NAND2xp5_ASAP7_75t_L g950 ( 
.A(n_820),
.B(n_916),
.Y(n_950)
);

O2A1O1Ixp33_ASAP7_75t_L g951 ( 
.A1(n_840),
.A2(n_15),
.B(n_18),
.C(n_20),
.Y(n_951)
);

AND2x4_ASAP7_75t_L g952 ( 
.A(n_785),
.B(n_122),
.Y(n_952)
);

AND2x2_ASAP7_75t_L g953 ( 
.A(n_802),
.B(n_21),
.Y(n_953)
);

NAND2xp5_ASAP7_75t_L g954 ( 
.A(n_820),
.B(n_23),
.Y(n_954)
);

INVx2_ASAP7_75t_SL g955 ( 
.A(n_787),
.Y(n_955)
);

HB1xp67_ASAP7_75t_L g956 ( 
.A(n_856),
.Y(n_956)
);

AOI21xp5_ASAP7_75t_L g957 ( 
.A1(n_752),
.A2(n_116),
.B(n_115),
.Y(n_957)
);

CKINVDCx5p33_ASAP7_75t_R g958 ( 
.A(n_879),
.Y(n_958)
);

BUFx6f_ASAP7_75t_L g959 ( 
.A(n_753),
.Y(n_959)
);

NAND2xp5_ASAP7_75t_L g960 ( 
.A(n_750),
.B(n_26),
.Y(n_960)
);

AO32x1_ASAP7_75t_L g961 ( 
.A1(n_872),
.A2(n_28),
.A3(n_30),
.B1(n_31),
.B2(n_34),
.Y(n_961)
);

NOR3xp33_ASAP7_75t_SL g962 ( 
.A(n_749),
.B(n_30),
.C(n_34),
.Y(n_962)
);

INVx1_ASAP7_75t_L g963 ( 
.A(n_803),
.Y(n_963)
);

OR2x6_ASAP7_75t_L g964 ( 
.A(n_865),
.B(n_35),
.Y(n_964)
);

O2A1O1Ixp33_ASAP7_75t_L g965 ( 
.A1(n_888),
.A2(n_36),
.B(n_37),
.C(n_38),
.Y(n_965)
);

BUFx8_ASAP7_75t_L g966 ( 
.A(n_793),
.Y(n_966)
);

A2O1A1Ixp33_ASAP7_75t_L g967 ( 
.A1(n_898),
.A2(n_40),
.B(n_41),
.C(n_44),
.Y(n_967)
);

BUFx6f_ASAP7_75t_L g968 ( 
.A(n_757),
.Y(n_968)
);

OAI21x1_ASAP7_75t_L g969 ( 
.A1(n_829),
.A2(n_92),
.B(n_108),
.Y(n_969)
);

AOI33xp33_ASAP7_75t_L g970 ( 
.A1(n_806),
.A2(n_40),
.A3(n_41),
.B1(n_45),
.B2(n_53),
.B3(n_66),
.Y(n_970)
);

A2O1A1Ixp33_ASAP7_75t_SL g971 ( 
.A1(n_775),
.A2(n_67),
.B(n_96),
.C(n_101),
.Y(n_971)
);

INVx2_ASAP7_75t_SL g972 ( 
.A(n_787),
.Y(n_972)
);

CKINVDCx5p33_ASAP7_75t_R g973 ( 
.A(n_858),
.Y(n_973)
);

NOR2xp67_ASAP7_75t_L g974 ( 
.A(n_822),
.B(n_103),
.Y(n_974)
);

INVx1_ASAP7_75t_L g975 ( 
.A(n_809),
.Y(n_975)
);

A2O1A1Ixp33_ASAP7_75t_L g976 ( 
.A1(n_877),
.A2(n_107),
.B(n_113),
.C(n_890),
.Y(n_976)
);

AND2x2_ASAP7_75t_L g977 ( 
.A(n_894),
.B(n_823),
.Y(n_977)
);

INVx5_ASAP7_75t_L g978 ( 
.A(n_865),
.Y(n_978)
);

INVx1_ASAP7_75t_L g979 ( 
.A(n_811),
.Y(n_979)
);

NAND2xp5_ASAP7_75t_SL g980 ( 
.A(n_854),
.B(n_752),
.Y(n_980)
);

INVx1_ASAP7_75t_L g981 ( 
.A(n_825),
.Y(n_981)
);

OAI22xp5_ASAP7_75t_L g982 ( 
.A1(n_807),
.A2(n_766),
.B1(n_758),
.B2(n_868),
.Y(n_982)
);

AOI21xp5_ASAP7_75t_L g983 ( 
.A1(n_758),
.A2(n_759),
.B(n_798),
.Y(n_983)
);

AOI21xp5_ASAP7_75t_L g984 ( 
.A1(n_758),
.A2(n_772),
.B(n_766),
.Y(n_984)
);

NAND2xp5_ASAP7_75t_L g985 ( 
.A(n_831),
.B(n_841),
.Y(n_985)
);

BUFx6f_ASAP7_75t_L g986 ( 
.A(n_757),
.Y(n_986)
);

NOR2xp33_ASAP7_75t_SL g987 ( 
.A(n_782),
.B(n_865),
.Y(n_987)
);

AOI21xp5_ASAP7_75t_L g988 ( 
.A1(n_758),
.A2(n_772),
.B(n_887),
.Y(n_988)
);

NOR2xp33_ASAP7_75t_L g989 ( 
.A(n_896),
.B(n_832),
.Y(n_989)
);

AOI21xp5_ASAP7_75t_L g990 ( 
.A1(n_772),
.A2(n_861),
.B(n_795),
.Y(n_990)
);

BUFx6f_ASAP7_75t_L g991 ( 
.A(n_757),
.Y(n_991)
);

OAI22xp5_ASAP7_75t_L g992 ( 
.A1(n_807),
.A2(n_868),
.B1(n_804),
.B2(n_763),
.Y(n_992)
);

AOI22xp5_ASAP7_75t_L g993 ( 
.A1(n_785),
.A2(n_839),
.B1(n_847),
.B2(n_850),
.Y(n_993)
);

INVx1_ASAP7_75t_L g994 ( 
.A(n_844),
.Y(n_994)
);

OR2x6_ASAP7_75t_L g995 ( 
.A(n_796),
.B(n_868),
.Y(n_995)
);

BUFx2_ASAP7_75t_SL g996 ( 
.A(n_810),
.Y(n_996)
);

NAND2xp5_ASAP7_75t_L g997 ( 
.A(n_902),
.B(n_907),
.Y(n_997)
);

INVx1_ASAP7_75t_L g998 ( 
.A(n_776),
.Y(n_998)
);

BUFx3_ASAP7_75t_L g999 ( 
.A(n_816),
.Y(n_999)
);

AOI21xp5_ASAP7_75t_L g1000 ( 
.A1(n_861),
.A2(n_768),
.B(n_795),
.Y(n_1000)
);

NAND2xp5_ASAP7_75t_L g1001 ( 
.A(n_908),
.B(n_915),
.Y(n_1001)
);

NAND2xp5_ASAP7_75t_L g1002 ( 
.A(n_760),
.B(n_779),
.Y(n_1002)
);

INVx1_ASAP7_75t_L g1003 ( 
.A(n_778),
.Y(n_1003)
);

INVx4_ASAP7_75t_L g1004 ( 
.A(n_816),
.Y(n_1004)
);

INVx1_ASAP7_75t_L g1005 ( 
.A(n_784),
.Y(n_1005)
);

HB1xp67_ASAP7_75t_L g1006 ( 
.A(n_791),
.Y(n_1006)
);

BUFx6f_ASAP7_75t_L g1007 ( 
.A(n_762),
.Y(n_1007)
);

BUFx12f_ASAP7_75t_L g1008 ( 
.A(n_786),
.Y(n_1008)
);

INVx5_ASAP7_75t_L g1009 ( 
.A(n_846),
.Y(n_1009)
);

O2A1O1Ixp5_ASAP7_75t_L g1010 ( 
.A1(n_895),
.A2(n_899),
.B(n_876),
.C(n_871),
.Y(n_1010)
);

NAND2xp5_ASAP7_75t_L g1011 ( 
.A(n_860),
.B(n_864),
.Y(n_1011)
);

OAI22xp5_ASAP7_75t_L g1012 ( 
.A1(n_804),
.A2(n_855),
.B1(n_828),
.B2(n_826),
.Y(n_1012)
);

AND2x2_ASAP7_75t_L g1013 ( 
.A(n_754),
.B(n_874),
.Y(n_1013)
);

AOI21xp5_ASAP7_75t_L g1014 ( 
.A1(n_768),
.A2(n_794),
.B(n_769),
.Y(n_1014)
);

INVx1_ASAP7_75t_SL g1015 ( 
.A(n_843),
.Y(n_1015)
);

AOI221xp5_ASAP7_75t_L g1016 ( 
.A1(n_904),
.A2(n_919),
.B1(n_751),
.B2(n_853),
.C(n_855),
.Y(n_1016)
);

OAI22xp5_ASAP7_75t_L g1017 ( 
.A1(n_826),
.A2(n_828),
.B1(n_878),
.B2(n_815),
.Y(n_1017)
);

O2A1O1Ixp33_ASAP7_75t_L g1018 ( 
.A1(n_805),
.A2(n_903),
.B(n_821),
.C(n_880),
.Y(n_1018)
);

INVx6_ASAP7_75t_L g1019 ( 
.A(n_788),
.Y(n_1019)
);

INVx2_ASAP7_75t_SL g1020 ( 
.A(n_756),
.Y(n_1020)
);

AOI21xp5_ASAP7_75t_L g1021 ( 
.A1(n_769),
.A2(n_794),
.B(n_857),
.Y(n_1021)
);

BUFx6f_ASAP7_75t_L g1022 ( 
.A(n_762),
.Y(n_1022)
);

CKINVDCx11_ASAP7_75t_R g1023 ( 
.A(n_881),
.Y(n_1023)
);

OAI22xp5_ASAP7_75t_L g1024 ( 
.A1(n_857),
.A2(n_814),
.B1(n_800),
.B2(n_889),
.Y(n_1024)
);

O2A1O1Ixp33_ASAP7_75t_L g1025 ( 
.A1(n_835),
.A2(n_808),
.B(n_817),
.C(n_827),
.Y(n_1025)
);

OAI22xp5_ASAP7_75t_L g1026 ( 
.A1(n_800),
.A2(n_889),
.B1(n_852),
.B2(n_842),
.Y(n_1026)
);

INVx2_ASAP7_75t_L g1027 ( 
.A(n_773),
.Y(n_1027)
);

INVx1_ASAP7_75t_L g1028 ( 
.A(n_789),
.Y(n_1028)
);

NAND2xp5_ASAP7_75t_L g1029 ( 
.A(n_869),
.B(n_797),
.Y(n_1029)
);

A2O1A1Ixp33_ASAP7_75t_L g1030 ( 
.A1(n_783),
.A2(n_770),
.B(n_780),
.C(n_918),
.Y(n_1030)
);

AOI21xp5_ASAP7_75t_L g1031 ( 
.A1(n_869),
.A2(n_859),
.B(n_906),
.Y(n_1031)
);

NOR2xp33_ASAP7_75t_L g1032 ( 
.A(n_892),
.B(n_883),
.Y(n_1032)
);

OR2x6_ASAP7_75t_L g1033 ( 
.A(n_881),
.B(n_886),
.Y(n_1033)
);

INVx5_ASAP7_75t_L g1034 ( 
.A(n_846),
.Y(n_1034)
);

O2A1O1Ixp33_ASAP7_75t_L g1035 ( 
.A1(n_808),
.A2(n_852),
.B(n_827),
.C(n_842),
.Y(n_1035)
);

NAND2xp5_ASAP7_75t_L g1036 ( 
.A(n_792),
.B(n_906),
.Y(n_1036)
);

OAI22xp5_ASAP7_75t_L g1037 ( 
.A1(n_817),
.A2(n_764),
.B1(n_862),
.B2(n_891),
.Y(n_1037)
);

NAND2xp5_ASAP7_75t_SL g1038 ( 
.A(n_867),
.B(n_774),
.Y(n_1038)
);

AOI21xp5_ASAP7_75t_L g1039 ( 
.A1(n_859),
.A2(n_897),
.B(n_905),
.Y(n_1039)
);

AND2x4_ASAP7_75t_L g1040 ( 
.A(n_824),
.B(n_870),
.Y(n_1040)
);

AOI21xp5_ASAP7_75t_L g1041 ( 
.A1(n_884),
.A2(n_905),
.B(n_897),
.Y(n_1041)
);

INVx2_ASAP7_75t_L g1042 ( 
.A(n_812),
.Y(n_1042)
);

NAND2xp5_ASAP7_75t_L g1043 ( 
.A(n_833),
.B(n_837),
.Y(n_1043)
);

INVx2_ASAP7_75t_SL g1044 ( 
.A(n_851),
.Y(n_1044)
);

OR2x2_ASAP7_75t_L g1045 ( 
.A(n_875),
.B(n_882),
.Y(n_1045)
);

OAI21xp33_ASAP7_75t_SL g1046 ( 
.A1(n_884),
.A2(n_885),
.B(n_893),
.Y(n_1046)
);

AO22x1_ASAP7_75t_L g1047 ( 
.A1(n_780),
.A2(n_863),
.B1(n_893),
.B2(n_885),
.Y(n_1047)
);

NOR2xp33_ASAP7_75t_L g1048 ( 
.A(n_863),
.B(n_849),
.Y(n_1048)
);

OAI22x1_ASAP7_75t_L g1049 ( 
.A1(n_911),
.A2(n_912),
.B1(n_845),
.B2(n_914),
.Y(n_1049)
);

A2O1A1Ixp33_ASAP7_75t_L g1050 ( 
.A1(n_770),
.A2(n_918),
.B(n_866),
.C(n_777),
.Y(n_1050)
);

AOI21xp5_ASAP7_75t_SL g1051 ( 
.A1(n_983),
.A2(n_771),
.B(n_873),
.Y(n_1051)
);

INVx3_ASAP7_75t_L g1052 ( 
.A(n_1007),
.Y(n_1052)
);

NAND2xp5_ASAP7_75t_L g1053 ( 
.A(n_950),
.B(n_771),
.Y(n_1053)
);

INVx1_ASAP7_75t_L g1054 ( 
.A(n_949),
.Y(n_1054)
);

AOI21xp5_ASAP7_75t_L g1055 ( 
.A1(n_1021),
.A2(n_909),
.B(n_1000),
.Y(n_1055)
);

NAND2xp5_ASAP7_75t_L g1056 ( 
.A(n_931),
.B(n_925),
.Y(n_1056)
);

AOI21xp5_ASAP7_75t_L g1057 ( 
.A1(n_1031),
.A2(n_1030),
.B(n_928),
.Y(n_1057)
);

INVx2_ASAP7_75t_L g1058 ( 
.A(n_1045),
.Y(n_1058)
);

BUFx3_ASAP7_75t_L g1059 ( 
.A(n_978),
.Y(n_1059)
);

OAI21xp5_ASAP7_75t_L g1060 ( 
.A1(n_1050),
.A2(n_1046),
.B(n_1014),
.Y(n_1060)
);

NAND2x1p5_ASAP7_75t_L g1061 ( 
.A(n_1009),
.B(n_1034),
.Y(n_1061)
);

AND2x2_ASAP7_75t_L g1062 ( 
.A(n_932),
.B(n_924),
.Y(n_1062)
);

AOI21xp5_ASAP7_75t_L g1063 ( 
.A1(n_926),
.A2(n_1035),
.B(n_988),
.Y(n_1063)
);

BUFx3_ASAP7_75t_L g1064 ( 
.A(n_978),
.Y(n_1064)
);

INVx2_ASAP7_75t_L g1065 ( 
.A(n_963),
.Y(n_1065)
);

OAI21x1_ASAP7_75t_L g1066 ( 
.A1(n_1039),
.A2(n_969),
.B(n_945),
.Y(n_1066)
);

OAI21xp5_ASAP7_75t_L g1067 ( 
.A1(n_1018),
.A2(n_1010),
.B(n_938),
.Y(n_1067)
);

AOI21xp5_ASAP7_75t_L g1068 ( 
.A1(n_990),
.A2(n_1025),
.B(n_1037),
.Y(n_1068)
);

OAI21x1_ASAP7_75t_L g1069 ( 
.A1(n_1041),
.A2(n_984),
.B(n_1012),
.Y(n_1069)
);

AOI21xp5_ASAP7_75t_L g1070 ( 
.A1(n_1024),
.A2(n_940),
.B(n_1049),
.Y(n_1070)
);

NAND2xp5_ASAP7_75t_L g1071 ( 
.A(n_997),
.B(n_1001),
.Y(n_1071)
);

INVx1_ASAP7_75t_L g1072 ( 
.A(n_975),
.Y(n_1072)
);

AO31x2_ASAP7_75t_L g1073 ( 
.A1(n_939),
.A2(n_1026),
.A3(n_1048),
.B(n_1017),
.Y(n_1073)
);

AO22x2_ASAP7_75t_L g1074 ( 
.A1(n_960),
.A2(n_943),
.B1(n_954),
.B2(n_1013),
.Y(n_1074)
);

INVx1_ASAP7_75t_L g1075 ( 
.A(n_979),
.Y(n_1075)
);

NAND3xp33_ASAP7_75t_L g1076 ( 
.A(n_962),
.B(n_929),
.C(n_1016),
.Y(n_1076)
);

INVx1_ASAP7_75t_SL g1077 ( 
.A(n_922),
.Y(n_1077)
);

OR2x6_ASAP7_75t_L g1078 ( 
.A(n_1033),
.B(n_996),
.Y(n_1078)
);

INVx1_ASAP7_75t_L g1079 ( 
.A(n_981),
.Y(n_1079)
);

AND2x2_ASAP7_75t_L g1080 ( 
.A(n_977),
.B(n_935),
.Y(n_1080)
);

NAND2xp5_ASAP7_75t_L g1081 ( 
.A(n_947),
.B(n_1006),
.Y(n_1081)
);

AOI21x1_ASAP7_75t_L g1082 ( 
.A1(n_1047),
.A2(n_1002),
.B(n_937),
.Y(n_1082)
);

OAI21x1_ASAP7_75t_L g1083 ( 
.A1(n_941),
.A2(n_1029),
.B(n_1036),
.Y(n_1083)
);

AOI21xp5_ASAP7_75t_L g1084 ( 
.A1(n_1011),
.A2(n_1034),
.B(n_1009),
.Y(n_1084)
);

NAND2xp5_ASAP7_75t_L g1085 ( 
.A(n_989),
.B(n_985),
.Y(n_1085)
);

CKINVDCx20_ASAP7_75t_R g1086 ( 
.A(n_958),
.Y(n_1086)
);

NAND2xp5_ASAP7_75t_L g1087 ( 
.A(n_994),
.B(n_933),
.Y(n_1087)
);

OAI21xp5_ASAP7_75t_SL g1088 ( 
.A1(n_951),
.A2(n_967),
.B(n_965),
.Y(n_1088)
);

INVx1_ASAP7_75t_L g1089 ( 
.A(n_998),
.Y(n_1089)
);

AOI21xp5_ASAP7_75t_L g1090 ( 
.A1(n_1038),
.A2(n_980),
.B(n_1032),
.Y(n_1090)
);

OAI21x1_ASAP7_75t_L g1091 ( 
.A1(n_921),
.A2(n_927),
.B(n_1003),
.Y(n_1091)
);

INVx2_ASAP7_75t_L g1092 ( 
.A(n_934),
.Y(n_1092)
);

OAI21x1_ASAP7_75t_SL g1093 ( 
.A1(n_957),
.A2(n_993),
.B(n_1005),
.Y(n_1093)
);

O2A1O1Ixp33_ASAP7_75t_SL g1094 ( 
.A1(n_976),
.A2(n_956),
.B(n_1043),
.C(n_1028),
.Y(n_1094)
);

NAND2x1p5_ASAP7_75t_L g1095 ( 
.A(n_978),
.B(n_1004),
.Y(n_1095)
);

BUFx6f_ASAP7_75t_L g1096 ( 
.A(n_920),
.Y(n_1096)
);

AOI21xp5_ASAP7_75t_L g1097 ( 
.A1(n_1040),
.A2(n_1020),
.B(n_952),
.Y(n_1097)
);

AOI21xp5_ASAP7_75t_SL g1098 ( 
.A1(n_952),
.A2(n_1040),
.B(n_959),
.Y(n_1098)
);

NAND2xp5_ASAP7_75t_L g1099 ( 
.A(n_1044),
.B(n_1042),
.Y(n_1099)
);

AOI21xp5_ASAP7_75t_L g1100 ( 
.A1(n_1027),
.A2(n_942),
.B(n_974),
.Y(n_1100)
);

BUFx4f_ASAP7_75t_L g1101 ( 
.A(n_923),
.Y(n_1101)
);

NAND2xp5_ASAP7_75t_L g1102 ( 
.A(n_953),
.B(n_970),
.Y(n_1102)
);

OAI21xp5_ASAP7_75t_L g1103 ( 
.A1(n_995),
.A2(n_1004),
.B(n_972),
.Y(n_1103)
);

AOI21xp5_ASAP7_75t_L g1104 ( 
.A1(n_1007),
.A2(n_1022),
.B(n_991),
.Y(n_1104)
);

OAI21x1_ASAP7_75t_SL g1105 ( 
.A1(n_955),
.A2(n_1023),
.B(n_961),
.Y(n_1105)
);

CKINVDCx5p33_ASAP7_75t_R g1106 ( 
.A(n_973),
.Y(n_1106)
);

INVx4_ASAP7_75t_L g1107 ( 
.A(n_1019),
.Y(n_1107)
);

NAND2xp5_ASAP7_75t_L g1108 ( 
.A(n_999),
.B(n_1022),
.Y(n_1108)
);

OAI21x1_ASAP7_75t_L g1109 ( 
.A1(n_1007),
.A2(n_1022),
.B(n_968),
.Y(n_1109)
);

OAI21x1_ASAP7_75t_L g1110 ( 
.A1(n_959),
.A2(n_968),
.B(n_991),
.Y(n_1110)
);

AOI21xp33_ASAP7_75t_L g1111 ( 
.A1(n_995),
.A2(n_987),
.B(n_964),
.Y(n_1111)
);

OAI21xp5_ASAP7_75t_L g1112 ( 
.A1(n_964),
.A2(n_961),
.B(n_1015),
.Y(n_1112)
);

AO32x2_ASAP7_75t_L g1113 ( 
.A1(n_961),
.A2(n_986),
.A3(n_936),
.B1(n_946),
.B2(n_920),
.Y(n_1113)
);

OA21x2_ASAP7_75t_L g1114 ( 
.A1(n_986),
.A2(n_920),
.B(n_936),
.Y(n_1114)
);

INVx1_ASAP7_75t_L g1115 ( 
.A(n_936),
.Y(n_1115)
);

CKINVDCx5p33_ASAP7_75t_R g1116 ( 
.A(n_944),
.Y(n_1116)
);

NOR2xp33_ASAP7_75t_L g1117 ( 
.A(n_1008),
.B(n_986),
.Y(n_1117)
);

AOI21xp5_ASAP7_75t_L g1118 ( 
.A1(n_946),
.A2(n_758),
.B(n_752),
.Y(n_1118)
);

OAI21x1_ASAP7_75t_SL g1119 ( 
.A1(n_946),
.A2(n_872),
.B(n_856),
.Y(n_1119)
);

INVx1_ASAP7_75t_L g1120 ( 
.A(n_966),
.Y(n_1120)
);

AO31x2_ASAP7_75t_L g1121 ( 
.A1(n_1030),
.A2(n_1050),
.A3(n_982),
.B(n_1037),
.Y(n_1121)
);

A2O1A1Ixp33_ASAP7_75t_L g1122 ( 
.A1(n_930),
.A2(n_910),
.B(n_600),
.C(n_619),
.Y(n_1122)
);

OR2x2_ASAP7_75t_L g1123 ( 
.A(n_922),
.B(n_950),
.Y(n_1123)
);

AOI21x1_ASAP7_75t_L g1124 ( 
.A1(n_1047),
.A2(n_1031),
.B(n_990),
.Y(n_1124)
);

INVx2_ASAP7_75t_L g1125 ( 
.A(n_1045),
.Y(n_1125)
);

OR2x2_ASAP7_75t_L g1126 ( 
.A(n_922),
.B(n_950),
.Y(n_1126)
);

BUFx6f_ASAP7_75t_L g1127 ( 
.A(n_920),
.Y(n_1127)
);

INVx1_ASAP7_75t_L g1128 ( 
.A(n_949),
.Y(n_1128)
);

INVx1_ASAP7_75t_SL g1129 ( 
.A(n_922),
.Y(n_1129)
);

NOR2xp33_ASAP7_75t_L g1130 ( 
.A(n_931),
.B(n_627),
.Y(n_1130)
);

CKINVDCx9p33_ASAP7_75t_R g1131 ( 
.A(n_989),
.Y(n_1131)
);

NAND2xp5_ASAP7_75t_L g1132 ( 
.A(n_950),
.B(n_818),
.Y(n_1132)
);

AND2x2_ASAP7_75t_L g1133 ( 
.A(n_932),
.B(n_924),
.Y(n_1133)
);

INVx1_ASAP7_75t_L g1134 ( 
.A(n_949),
.Y(n_1134)
);

OAI21x1_ASAP7_75t_L g1135 ( 
.A1(n_1014),
.A2(n_829),
.B(n_1039),
.Y(n_1135)
);

AND2x4_ASAP7_75t_L g1136 ( 
.A(n_978),
.B(n_977),
.Y(n_1136)
);

OAI22xp5_ASAP7_75t_L g1137 ( 
.A1(n_931),
.A2(n_600),
.B1(n_910),
.B2(n_819),
.Y(n_1137)
);

AO31x2_ASAP7_75t_L g1138 ( 
.A1(n_1030),
.A2(n_1050),
.A3(n_982),
.B(n_1037),
.Y(n_1138)
);

INVx1_ASAP7_75t_L g1139 ( 
.A(n_949),
.Y(n_1139)
);

AND2x2_ASAP7_75t_L g1140 ( 
.A(n_932),
.B(n_924),
.Y(n_1140)
);

CKINVDCx5p33_ASAP7_75t_R g1141 ( 
.A(n_958),
.Y(n_1141)
);

INVx2_ASAP7_75t_SL g1142 ( 
.A(n_955),
.Y(n_1142)
);

OAI21x1_ASAP7_75t_L g1143 ( 
.A1(n_1014),
.A2(n_829),
.B(n_1039),
.Y(n_1143)
);

A2O1A1Ixp33_ASAP7_75t_L g1144 ( 
.A1(n_930),
.A2(n_910),
.B(n_600),
.C(n_619),
.Y(n_1144)
);

AND2x4_ASAP7_75t_L g1145 ( 
.A(n_978),
.B(n_977),
.Y(n_1145)
);

AO31x2_ASAP7_75t_L g1146 ( 
.A1(n_1030),
.A2(n_1050),
.A3(n_982),
.B(n_1037),
.Y(n_1146)
);

OAI21x1_ASAP7_75t_L g1147 ( 
.A1(n_1014),
.A2(n_829),
.B(n_1039),
.Y(n_1147)
);

NAND2xp5_ASAP7_75t_L g1148 ( 
.A(n_950),
.B(n_818),
.Y(n_1148)
);

BUFx6f_ASAP7_75t_L g1149 ( 
.A(n_920),
.Y(n_1149)
);

INVx6_ASAP7_75t_L g1150 ( 
.A(n_978),
.Y(n_1150)
);

INVxp67_ASAP7_75t_SL g1151 ( 
.A(n_950),
.Y(n_1151)
);

INVx1_ASAP7_75t_L g1152 ( 
.A(n_949),
.Y(n_1152)
);

NAND3x1_ASAP7_75t_L g1153 ( 
.A(n_993),
.B(n_482),
.C(n_686),
.Y(n_1153)
);

O2A1O1Ixp33_ASAP7_75t_SL g1154 ( 
.A1(n_976),
.A2(n_900),
.B(n_971),
.C(n_967),
.Y(n_1154)
);

OAI21xp5_ASAP7_75t_L g1155 ( 
.A1(n_1030),
.A2(n_1050),
.B(n_1031),
.Y(n_1155)
);

BUFx2_ASAP7_75t_L g1156 ( 
.A(n_948),
.Y(n_1156)
);

INVx1_ASAP7_75t_L g1157 ( 
.A(n_949),
.Y(n_1157)
);

INVx1_ASAP7_75t_L g1158 ( 
.A(n_949),
.Y(n_1158)
);

OR2x2_ASAP7_75t_L g1159 ( 
.A(n_922),
.B(n_950),
.Y(n_1159)
);

NAND2xp5_ASAP7_75t_L g1160 ( 
.A(n_950),
.B(n_818),
.Y(n_1160)
);

OAI22xp5_ASAP7_75t_L g1161 ( 
.A1(n_931),
.A2(n_600),
.B1(n_910),
.B2(n_819),
.Y(n_1161)
);

AO21x2_ASAP7_75t_L g1162 ( 
.A1(n_1030),
.A2(n_1050),
.B(n_982),
.Y(n_1162)
);

OAI21x1_ASAP7_75t_L g1163 ( 
.A1(n_1014),
.A2(n_829),
.B(n_1039),
.Y(n_1163)
);

NAND2xp5_ASAP7_75t_L g1164 ( 
.A(n_950),
.B(n_818),
.Y(n_1164)
);

AND2x4_ASAP7_75t_L g1165 ( 
.A(n_978),
.B(n_977),
.Y(n_1165)
);

OAI21x1_ASAP7_75t_L g1166 ( 
.A1(n_1014),
.A2(n_829),
.B(n_1039),
.Y(n_1166)
);

AOI21xp5_ASAP7_75t_L g1167 ( 
.A1(n_983),
.A2(n_758),
.B(n_752),
.Y(n_1167)
);

OAI22xp5_ASAP7_75t_L g1168 ( 
.A1(n_931),
.A2(n_600),
.B1(n_910),
.B2(n_819),
.Y(n_1168)
);

OA21x2_ASAP7_75t_L g1169 ( 
.A1(n_1030),
.A2(n_1050),
.B(n_1010),
.Y(n_1169)
);

OAI21xp5_ASAP7_75t_L g1170 ( 
.A1(n_1030),
.A2(n_1050),
.B(n_1031),
.Y(n_1170)
);

NAND2xp5_ASAP7_75t_L g1171 ( 
.A(n_950),
.B(n_818),
.Y(n_1171)
);

AOI21x1_ASAP7_75t_L g1172 ( 
.A1(n_1047),
.A2(n_1031),
.B(n_990),
.Y(n_1172)
);

BUFx2_ASAP7_75t_L g1173 ( 
.A(n_948),
.Y(n_1173)
);

INVx1_ASAP7_75t_L g1174 ( 
.A(n_949),
.Y(n_1174)
);

OAI21x1_ASAP7_75t_SL g1175 ( 
.A1(n_983),
.A2(n_872),
.B(n_856),
.Y(n_1175)
);

NAND2xp5_ASAP7_75t_L g1176 ( 
.A(n_950),
.B(n_818),
.Y(n_1176)
);

AO32x2_ASAP7_75t_L g1177 ( 
.A1(n_982),
.A2(n_992),
.A3(n_856),
.B1(n_872),
.B2(n_1012),
.Y(n_1177)
);

OAI21x1_ASAP7_75t_L g1178 ( 
.A1(n_1014),
.A2(n_829),
.B(n_1039),
.Y(n_1178)
);

OAI21xp5_ASAP7_75t_L g1179 ( 
.A1(n_1030),
.A2(n_1050),
.B(n_1031),
.Y(n_1179)
);

INVx1_ASAP7_75t_L g1180 ( 
.A(n_949),
.Y(n_1180)
);

OAI22xp5_ASAP7_75t_L g1181 ( 
.A1(n_931),
.A2(n_600),
.B1(n_910),
.B2(n_819),
.Y(n_1181)
);

AOI21xp5_ASAP7_75t_L g1182 ( 
.A1(n_983),
.A2(n_758),
.B(n_752),
.Y(n_1182)
);

OAI21x1_ASAP7_75t_L g1183 ( 
.A1(n_1014),
.A2(n_829),
.B(n_1039),
.Y(n_1183)
);

INVx4_ASAP7_75t_L g1184 ( 
.A(n_1009),
.Y(n_1184)
);

NAND2xp5_ASAP7_75t_L g1185 ( 
.A(n_950),
.B(n_818),
.Y(n_1185)
);

OAI21x1_ASAP7_75t_L g1186 ( 
.A1(n_1014),
.A2(n_829),
.B(n_1039),
.Y(n_1186)
);

OAI21x1_ASAP7_75t_L g1187 ( 
.A1(n_1147),
.A2(n_1166),
.B(n_1163),
.Y(n_1187)
);

OAI21x1_ASAP7_75t_L g1188 ( 
.A1(n_1178),
.A2(n_1186),
.B(n_1183),
.Y(n_1188)
);

NOR2xp33_ASAP7_75t_L g1189 ( 
.A(n_1137),
.B(n_1161),
.Y(n_1189)
);

OA21x2_ASAP7_75t_L g1190 ( 
.A1(n_1063),
.A2(n_1060),
.B(n_1068),
.Y(n_1190)
);

HB1xp67_ASAP7_75t_L g1191 ( 
.A(n_1077),
.Y(n_1191)
);

INVx2_ASAP7_75t_L g1192 ( 
.A(n_1065),
.Y(n_1192)
);

INVx1_ASAP7_75t_L g1193 ( 
.A(n_1054),
.Y(n_1193)
);

OAI21xp5_ASAP7_75t_L g1194 ( 
.A1(n_1122),
.A2(n_1144),
.B(n_1168),
.Y(n_1194)
);

BUFx2_ASAP7_75t_L g1195 ( 
.A(n_1156),
.Y(n_1195)
);

AND2x4_ASAP7_75t_L g1196 ( 
.A(n_1103),
.B(n_1078),
.Y(n_1196)
);

AOI21xp5_ASAP7_75t_L g1197 ( 
.A1(n_1057),
.A2(n_1170),
.B(n_1155),
.Y(n_1197)
);

OA21x2_ASAP7_75t_L g1198 ( 
.A1(n_1060),
.A2(n_1067),
.B(n_1155),
.Y(n_1198)
);

OAI21x1_ASAP7_75t_L g1199 ( 
.A1(n_1055),
.A2(n_1069),
.B(n_1172),
.Y(n_1199)
);

AND2x2_ASAP7_75t_L g1200 ( 
.A(n_1062),
.B(n_1133),
.Y(n_1200)
);

OAI22xp5_ASAP7_75t_L g1201 ( 
.A1(n_1181),
.A2(n_1130),
.B1(n_1071),
.B2(n_1056),
.Y(n_1201)
);

INVx1_ASAP7_75t_L g1202 ( 
.A(n_1072),
.Y(n_1202)
);

INVx1_ASAP7_75t_SL g1203 ( 
.A(n_1129),
.Y(n_1203)
);

OAI21x1_ASAP7_75t_L g1204 ( 
.A1(n_1124),
.A2(n_1170),
.B(n_1179),
.Y(n_1204)
);

BUFx12f_ASAP7_75t_L g1205 ( 
.A(n_1141),
.Y(n_1205)
);

OAI21x1_ASAP7_75t_L g1206 ( 
.A1(n_1179),
.A2(n_1070),
.B(n_1067),
.Y(n_1206)
);

OAI22xp5_ASAP7_75t_L g1207 ( 
.A1(n_1076),
.A2(n_1085),
.B1(n_1185),
.B2(n_1176),
.Y(n_1207)
);

NAND2x1p5_ASAP7_75t_L g1208 ( 
.A(n_1184),
.B(n_1107),
.Y(n_1208)
);

NAND3xp33_ASAP7_75t_L g1209 ( 
.A(n_1076),
.B(n_1088),
.C(n_1160),
.Y(n_1209)
);

INVx1_ASAP7_75t_L g1210 ( 
.A(n_1075),
.Y(n_1210)
);

AND2x2_ASAP7_75t_L g1211 ( 
.A(n_1140),
.B(n_1080),
.Y(n_1211)
);

AOI22xp33_ASAP7_75t_L g1212 ( 
.A1(n_1132),
.A2(n_1171),
.B1(n_1148),
.B2(n_1164),
.Y(n_1212)
);

NAND2xp5_ASAP7_75t_L g1213 ( 
.A(n_1151),
.B(n_1123),
.Y(n_1213)
);

INVx2_ASAP7_75t_L g1214 ( 
.A(n_1079),
.Y(n_1214)
);

AOI21xp5_ASAP7_75t_L g1215 ( 
.A1(n_1167),
.A2(n_1182),
.B(n_1051),
.Y(n_1215)
);

INVx2_ASAP7_75t_L g1216 ( 
.A(n_1128),
.Y(n_1216)
);

INVx1_ASAP7_75t_L g1217 ( 
.A(n_1134),
.Y(n_1217)
);

OAI21x1_ASAP7_75t_L g1218 ( 
.A1(n_1083),
.A2(n_1082),
.B(n_1169),
.Y(n_1218)
);

HB1xp67_ASAP7_75t_L g1219 ( 
.A(n_1173),
.Y(n_1219)
);

INVx1_ASAP7_75t_L g1220 ( 
.A(n_1139),
.Y(n_1220)
);

INVx4_ASAP7_75t_SL g1221 ( 
.A(n_1150),
.Y(n_1221)
);

OAI21xp5_ASAP7_75t_L g1222 ( 
.A1(n_1153),
.A2(n_1090),
.B(n_1088),
.Y(n_1222)
);

AOI22x1_ASAP7_75t_L g1223 ( 
.A1(n_1074),
.A2(n_1100),
.B1(n_1084),
.B2(n_1105),
.Y(n_1223)
);

OAI22xp33_ASAP7_75t_L g1224 ( 
.A1(n_1081),
.A2(n_1087),
.B1(n_1159),
.B2(n_1126),
.Y(n_1224)
);

INVx1_ASAP7_75t_L g1225 ( 
.A(n_1152),
.Y(n_1225)
);

CKINVDCx16_ASAP7_75t_R g1226 ( 
.A(n_1086),
.Y(n_1226)
);

INVx2_ASAP7_75t_L g1227 ( 
.A(n_1157),
.Y(n_1227)
);

OA21x2_ASAP7_75t_L g1228 ( 
.A1(n_1053),
.A2(n_1102),
.B(n_1112),
.Y(n_1228)
);

OA21x2_ASAP7_75t_L g1229 ( 
.A1(n_1112),
.A2(n_1089),
.B(n_1158),
.Y(n_1229)
);

OAI21x1_ASAP7_75t_L g1230 ( 
.A1(n_1118),
.A2(n_1109),
.B(n_1103),
.Y(n_1230)
);

OAI21x1_ASAP7_75t_L g1231 ( 
.A1(n_1110),
.A2(n_1097),
.B(n_1104),
.Y(n_1231)
);

INVx2_ASAP7_75t_L g1232 ( 
.A(n_1174),
.Y(n_1232)
);

OAI22xp5_ASAP7_75t_L g1233 ( 
.A1(n_1074),
.A2(n_1098),
.B1(n_1078),
.B2(n_1145),
.Y(n_1233)
);

OAI21xp5_ASAP7_75t_L g1234 ( 
.A1(n_1154),
.A2(n_1094),
.B(n_1058),
.Y(n_1234)
);

NAND2xp5_ASAP7_75t_L g1235 ( 
.A(n_1125),
.B(n_1145),
.Y(n_1235)
);

INVx2_ASAP7_75t_L g1236 ( 
.A(n_1180),
.Y(n_1236)
);

INVx2_ASAP7_75t_L g1237 ( 
.A(n_1092),
.Y(n_1237)
);

INVx2_ASAP7_75t_L g1238 ( 
.A(n_1121),
.Y(n_1238)
);

AOI22xp33_ASAP7_75t_L g1239 ( 
.A1(n_1162),
.A2(n_1111),
.B1(n_1136),
.B2(n_1165),
.Y(n_1239)
);

AND2x4_ASAP7_75t_L g1240 ( 
.A(n_1078),
.B(n_1052),
.Y(n_1240)
);

OAI21xp5_ASAP7_75t_L g1241 ( 
.A1(n_1099),
.A2(n_1061),
.B(n_1108),
.Y(n_1241)
);

AOI22xp33_ASAP7_75t_L g1242 ( 
.A1(n_1120),
.A2(n_1101),
.B1(n_1150),
.B2(n_1064),
.Y(n_1242)
);

INVx2_ASAP7_75t_L g1243 ( 
.A(n_1121),
.Y(n_1243)
);

OA21x2_ASAP7_75t_L g1244 ( 
.A1(n_1177),
.A2(n_1146),
.B(n_1138),
.Y(n_1244)
);

HB1xp67_ASAP7_75t_L g1245 ( 
.A(n_1142),
.Y(n_1245)
);

AND2x4_ASAP7_75t_L g1246 ( 
.A(n_1052),
.B(n_1115),
.Y(n_1246)
);

AOI221xp5_ASAP7_75t_L g1247 ( 
.A1(n_1117),
.A2(n_1101),
.B1(n_1116),
.B2(n_1106),
.C(n_1059),
.Y(n_1247)
);

AOI22xp33_ASAP7_75t_L g1248 ( 
.A1(n_1184),
.A2(n_1131),
.B1(n_1096),
.B2(n_1149),
.Y(n_1248)
);

AOI22xp33_ASAP7_75t_L g1249 ( 
.A1(n_1096),
.A2(n_1149),
.B1(n_1127),
.B2(n_1095),
.Y(n_1249)
);

OAI21x1_ASAP7_75t_L g1250 ( 
.A1(n_1114),
.A2(n_1146),
.B(n_1138),
.Y(n_1250)
);

OAI21x1_ASAP7_75t_L g1251 ( 
.A1(n_1114),
.A2(n_1146),
.B(n_1138),
.Y(n_1251)
);

BUFx3_ASAP7_75t_L g1252 ( 
.A(n_1127),
.Y(n_1252)
);

INVx1_ASAP7_75t_L g1253 ( 
.A(n_1177),
.Y(n_1253)
);

AOI21xp5_ASAP7_75t_L g1254 ( 
.A1(n_1073),
.A2(n_1177),
.B(n_1113),
.Y(n_1254)
);

INVx1_ASAP7_75t_L g1255 ( 
.A(n_1073),
.Y(n_1255)
);

OAI21x1_ASAP7_75t_SL g1256 ( 
.A1(n_1113),
.A2(n_1175),
.B(n_1119),
.Y(n_1256)
);

INVx2_ASAP7_75t_L g1257 ( 
.A(n_1091),
.Y(n_1257)
);

INVx4_ASAP7_75t_L g1258 ( 
.A(n_1184),
.Y(n_1258)
);

INVx2_ASAP7_75t_SL g1259 ( 
.A(n_1150),
.Y(n_1259)
);

OAI21x1_ASAP7_75t_L g1260 ( 
.A1(n_1066),
.A2(n_1143),
.B(n_1135),
.Y(n_1260)
);

OAI22xp5_ASAP7_75t_L g1261 ( 
.A1(n_1137),
.A2(n_1168),
.B1(n_1181),
.B2(n_1161),
.Y(n_1261)
);

OAI21x1_ASAP7_75t_L g1262 ( 
.A1(n_1066),
.A2(n_1143),
.B(n_1135),
.Y(n_1262)
);

AND2x4_ASAP7_75t_L g1263 ( 
.A(n_1103),
.B(n_1078),
.Y(n_1263)
);

AO21x2_ASAP7_75t_L g1264 ( 
.A1(n_1063),
.A2(n_1068),
.B(n_1057),
.Y(n_1264)
);

BUFx2_ASAP7_75t_L g1265 ( 
.A(n_1156),
.Y(n_1265)
);

AO32x2_ASAP7_75t_L g1266 ( 
.A1(n_1137),
.A2(n_1168),
.A3(n_1181),
.B1(n_1161),
.B2(n_904),
.Y(n_1266)
);

OAI21x1_ASAP7_75t_L g1267 ( 
.A1(n_1066),
.A2(n_1143),
.B(n_1135),
.Y(n_1267)
);

AND2x2_ASAP7_75t_L g1268 ( 
.A(n_1062),
.B(n_1133),
.Y(n_1268)
);

AOI22xp5_ASAP7_75t_L g1269 ( 
.A1(n_1137),
.A2(n_1168),
.B1(n_1181),
.B2(n_1161),
.Y(n_1269)
);

NAND2x1_ASAP7_75t_L g1270 ( 
.A(n_1184),
.B(n_1175),
.Y(n_1270)
);

OR2x2_ASAP7_75t_L g1271 ( 
.A(n_1077),
.B(n_1129),
.Y(n_1271)
);

AND2x4_ASAP7_75t_L g1272 ( 
.A(n_1103),
.B(n_1078),
.Y(n_1272)
);

AOI222xp33_ASAP7_75t_L g1273 ( 
.A1(n_1137),
.A2(n_904),
.B1(n_674),
.B2(n_676),
.C1(n_1168),
.C2(n_1161),
.Y(n_1273)
);

OAI21x1_ASAP7_75t_SL g1274 ( 
.A1(n_1175),
.A2(n_1119),
.B(n_1093),
.Y(n_1274)
);

AOI22xp33_ASAP7_75t_L g1275 ( 
.A1(n_1137),
.A2(n_1161),
.B1(n_1181),
.B2(n_1168),
.Y(n_1275)
);

INVx1_ASAP7_75t_L g1276 ( 
.A(n_1065),
.Y(n_1276)
);

INVx1_ASAP7_75t_L g1277 ( 
.A(n_1065),
.Y(n_1277)
);

BUFx3_ASAP7_75t_L g1278 ( 
.A(n_1136),
.Y(n_1278)
);

AND2x4_ASAP7_75t_L g1279 ( 
.A(n_1103),
.B(n_1078),
.Y(n_1279)
);

AND3x2_ASAP7_75t_L g1280 ( 
.A(n_1130),
.B(n_388),
.C(n_627),
.Y(n_1280)
);

INVx3_ASAP7_75t_L g1281 ( 
.A(n_1184),
.Y(n_1281)
);

OAI21xp5_ASAP7_75t_L g1282 ( 
.A1(n_1122),
.A2(n_1144),
.B(n_1137),
.Y(n_1282)
);

BUFx3_ASAP7_75t_L g1283 ( 
.A(n_1136),
.Y(n_1283)
);

INVx4_ASAP7_75t_L g1284 ( 
.A(n_1184),
.Y(n_1284)
);

INVx1_ASAP7_75t_L g1285 ( 
.A(n_1065),
.Y(n_1285)
);

AND2x4_ASAP7_75t_L g1286 ( 
.A(n_1103),
.B(n_1078),
.Y(n_1286)
);

O2A1O1Ixp33_ASAP7_75t_L g1287 ( 
.A1(n_1137),
.A2(n_1168),
.B(n_1181),
.C(n_1161),
.Y(n_1287)
);

OAI21xp5_ASAP7_75t_L g1288 ( 
.A1(n_1122),
.A2(n_1144),
.B(n_1137),
.Y(n_1288)
);

OAI21xp5_ASAP7_75t_L g1289 ( 
.A1(n_1122),
.A2(n_1144),
.B(n_1137),
.Y(n_1289)
);

AOI22xp33_ASAP7_75t_L g1290 ( 
.A1(n_1137),
.A2(n_1161),
.B1(n_1181),
.B2(n_1168),
.Y(n_1290)
);

AND2x2_ASAP7_75t_L g1291 ( 
.A(n_1062),
.B(n_1133),
.Y(n_1291)
);

INVx2_ASAP7_75t_L g1292 ( 
.A(n_1091),
.Y(n_1292)
);

NAND2x1p5_ASAP7_75t_L g1293 ( 
.A(n_1184),
.B(n_1009),
.Y(n_1293)
);

AND2x4_ASAP7_75t_L g1294 ( 
.A(n_1103),
.B(n_1078),
.Y(n_1294)
);

AND2x4_ASAP7_75t_L g1295 ( 
.A(n_1103),
.B(n_1078),
.Y(n_1295)
);

BUFx6f_ASAP7_75t_L g1296 ( 
.A(n_1096),
.Y(n_1296)
);

INVx1_ASAP7_75t_L g1297 ( 
.A(n_1065),
.Y(n_1297)
);

BUFx3_ASAP7_75t_L g1298 ( 
.A(n_1136),
.Y(n_1298)
);

OAI22xp5_ASAP7_75t_L g1299 ( 
.A1(n_1275),
.A2(n_1290),
.B1(n_1269),
.B2(n_1209),
.Y(n_1299)
);

AND2x2_ASAP7_75t_L g1300 ( 
.A(n_1268),
.B(n_1200),
.Y(n_1300)
);

AND2x4_ASAP7_75t_L g1301 ( 
.A(n_1196),
.B(n_1263),
.Y(n_1301)
);

OAI22xp5_ASAP7_75t_L g1302 ( 
.A1(n_1275),
.A2(n_1290),
.B1(n_1212),
.B2(n_1189),
.Y(n_1302)
);

NAND2xp5_ASAP7_75t_L g1303 ( 
.A(n_1207),
.B(n_1213),
.Y(n_1303)
);

AOI221x1_ASAP7_75t_SL g1304 ( 
.A1(n_1261),
.A2(n_1224),
.B1(n_1233),
.B2(n_1235),
.C(n_1266),
.Y(n_1304)
);

AOI21x1_ASAP7_75t_SL g1305 ( 
.A1(n_1196),
.A2(n_1272),
.B(n_1263),
.Y(n_1305)
);

O2A1O1Ixp33_ASAP7_75t_L g1306 ( 
.A1(n_1273),
.A2(n_1287),
.B(n_1222),
.C(n_1289),
.Y(n_1306)
);

INVx2_ASAP7_75t_L g1307 ( 
.A(n_1214),
.Y(n_1307)
);

AOI21xp5_ASAP7_75t_SL g1308 ( 
.A1(n_1197),
.A2(n_1282),
.B(n_1194),
.Y(n_1308)
);

OAI22xp5_ASAP7_75t_L g1309 ( 
.A1(n_1248),
.A2(n_1242),
.B1(n_1239),
.B2(n_1203),
.Y(n_1309)
);

AOI21xp5_ASAP7_75t_L g1310 ( 
.A1(n_1198),
.A2(n_1215),
.B(n_1190),
.Y(n_1310)
);

CKINVDCx20_ASAP7_75t_R g1311 ( 
.A(n_1226),
.Y(n_1311)
);

NAND2xp5_ASAP7_75t_L g1312 ( 
.A(n_1268),
.B(n_1291),
.Y(n_1312)
);

O2A1O1Ixp5_ASAP7_75t_L g1313 ( 
.A1(n_1288),
.A2(n_1234),
.B(n_1254),
.C(n_1255),
.Y(n_1313)
);

OR2x2_ASAP7_75t_L g1314 ( 
.A(n_1271),
.B(n_1191),
.Y(n_1314)
);

OAI22xp5_ASAP7_75t_L g1315 ( 
.A1(n_1195),
.A2(n_1265),
.B1(n_1219),
.B2(n_1272),
.Y(n_1315)
);

CKINVDCx20_ASAP7_75t_R g1316 ( 
.A(n_1205),
.Y(n_1316)
);

NAND2xp5_ASAP7_75t_L g1317 ( 
.A(n_1211),
.B(n_1192),
.Y(n_1317)
);

AOI21x1_ASAP7_75t_SL g1318 ( 
.A1(n_1196),
.A2(n_1263),
.B(n_1279),
.Y(n_1318)
);

OAI22xp5_ASAP7_75t_L g1319 ( 
.A1(n_1272),
.A2(n_1294),
.B1(n_1279),
.B2(n_1286),
.Y(n_1319)
);

OAI22xp5_ASAP7_75t_L g1320 ( 
.A1(n_1279),
.A2(n_1294),
.B1(n_1286),
.B2(n_1295),
.Y(n_1320)
);

OA21x2_ASAP7_75t_L g1321 ( 
.A1(n_1218),
.A2(n_1204),
.B(n_1206),
.Y(n_1321)
);

INVxp67_ASAP7_75t_L g1322 ( 
.A(n_1216),
.Y(n_1322)
);

OR2x2_ASAP7_75t_L g1323 ( 
.A(n_1216),
.B(n_1227),
.Y(n_1323)
);

OAI22xp5_ASAP7_75t_L g1324 ( 
.A1(n_1286),
.A2(n_1294),
.B1(n_1295),
.B2(n_1245),
.Y(n_1324)
);

AND2x4_ASAP7_75t_L g1325 ( 
.A(n_1295),
.B(n_1240),
.Y(n_1325)
);

OAI22xp5_ASAP7_75t_L g1326 ( 
.A1(n_1249),
.A2(n_1283),
.B1(n_1298),
.B2(n_1278),
.Y(n_1326)
);

AOI221xp5_ASAP7_75t_L g1327 ( 
.A1(n_1266),
.A2(n_1220),
.B1(n_1217),
.B2(n_1210),
.C(n_1225),
.Y(n_1327)
);

CKINVDCx5p33_ASAP7_75t_R g1328 ( 
.A(n_1205),
.Y(n_1328)
);

INVx1_ASAP7_75t_L g1329 ( 
.A(n_1232),
.Y(n_1329)
);

CKINVDCx5p33_ASAP7_75t_R g1330 ( 
.A(n_1298),
.Y(n_1330)
);

NAND2xp5_ASAP7_75t_L g1331 ( 
.A(n_1192),
.B(n_1276),
.Y(n_1331)
);

OA21x2_ASAP7_75t_L g1332 ( 
.A1(n_1218),
.A2(n_1204),
.B(n_1206),
.Y(n_1332)
);

OAI22xp5_ASAP7_75t_L g1333 ( 
.A1(n_1249),
.A2(n_1240),
.B1(n_1259),
.B2(n_1202),
.Y(n_1333)
);

OR2x2_ASAP7_75t_L g1334 ( 
.A(n_1236),
.B(n_1229),
.Y(n_1334)
);

NAND2xp5_ASAP7_75t_L g1335 ( 
.A(n_1277),
.B(n_1285),
.Y(n_1335)
);

OAI22xp5_ASAP7_75t_L g1336 ( 
.A1(n_1259),
.A2(n_1193),
.B1(n_1198),
.B2(n_1247),
.Y(n_1336)
);

OA22x2_ASAP7_75t_L g1337 ( 
.A1(n_1280),
.A2(n_1241),
.B1(n_1256),
.B2(n_1274),
.Y(n_1337)
);

NOR2xp33_ASAP7_75t_L g1338 ( 
.A(n_1246),
.B(n_1297),
.Y(n_1338)
);

BUFx12f_ASAP7_75t_L g1339 ( 
.A(n_1296),
.Y(n_1339)
);

INVx1_ASAP7_75t_L g1340 ( 
.A(n_1229),
.Y(n_1340)
);

OAI22xp5_ASAP7_75t_L g1341 ( 
.A1(n_1208),
.A2(n_1223),
.B1(n_1293),
.B2(n_1228),
.Y(n_1341)
);

AND2x2_ASAP7_75t_L g1342 ( 
.A(n_1237),
.B(n_1246),
.Y(n_1342)
);

OR2x2_ASAP7_75t_L g1343 ( 
.A(n_1229),
.B(n_1228),
.Y(n_1343)
);

AOI21xp5_ASAP7_75t_SL g1344 ( 
.A1(n_1258),
.A2(n_1284),
.B(n_1190),
.Y(n_1344)
);

AOI21xp5_ASAP7_75t_L g1345 ( 
.A1(n_1190),
.A2(n_1264),
.B(n_1199),
.Y(n_1345)
);

CKINVDCx20_ASAP7_75t_R g1346 ( 
.A(n_1221),
.Y(n_1346)
);

CKINVDCx5p33_ASAP7_75t_R g1347 ( 
.A(n_1252),
.Y(n_1347)
);

AND2x4_ASAP7_75t_L g1348 ( 
.A(n_1221),
.B(n_1281),
.Y(n_1348)
);

O2A1O1Ixp5_ASAP7_75t_L g1349 ( 
.A1(n_1238),
.A2(n_1243),
.B(n_1270),
.C(n_1257),
.Y(n_1349)
);

OR2x2_ASAP7_75t_SL g1350 ( 
.A(n_1296),
.B(n_1244),
.Y(n_1350)
);

OR2x2_ASAP7_75t_L g1351 ( 
.A(n_1238),
.B(n_1243),
.Y(n_1351)
);

AND2x4_ASAP7_75t_L g1352 ( 
.A(n_1258),
.B(n_1284),
.Y(n_1352)
);

HB1xp67_ASAP7_75t_L g1353 ( 
.A(n_1250),
.Y(n_1353)
);

OR2x2_ASAP7_75t_L g1354 ( 
.A(n_1244),
.B(n_1253),
.Y(n_1354)
);

AND2x2_ASAP7_75t_L g1355 ( 
.A(n_1250),
.B(n_1251),
.Y(n_1355)
);

HB1xp67_ASAP7_75t_L g1356 ( 
.A(n_1251),
.Y(n_1356)
);

NOR2xp33_ASAP7_75t_L g1357 ( 
.A(n_1230),
.B(n_1292),
.Y(n_1357)
);

INVx1_ASAP7_75t_SL g1358 ( 
.A(n_1231),
.Y(n_1358)
);

OA21x2_ASAP7_75t_L g1359 ( 
.A1(n_1187),
.A2(n_1188),
.B(n_1267),
.Y(n_1359)
);

INVx2_ASAP7_75t_L g1360 ( 
.A(n_1231),
.Y(n_1360)
);

AND2x2_ASAP7_75t_SL g1361 ( 
.A(n_1260),
.B(n_1262),
.Y(n_1361)
);

OA21x2_ASAP7_75t_L g1362 ( 
.A1(n_1218),
.A2(n_1204),
.B(n_1206),
.Y(n_1362)
);

BUFx3_ASAP7_75t_L g1363 ( 
.A(n_1195),
.Y(n_1363)
);

AND2x2_ASAP7_75t_L g1364 ( 
.A(n_1268),
.B(n_1200),
.Y(n_1364)
);

NAND2xp5_ASAP7_75t_L g1365 ( 
.A(n_1201),
.B(n_1212),
.Y(n_1365)
);

OAI22xp5_ASAP7_75t_L g1366 ( 
.A1(n_1275),
.A2(n_1130),
.B1(n_1290),
.B2(n_1076),
.Y(n_1366)
);

AOI21xp5_ASAP7_75t_L g1367 ( 
.A1(n_1197),
.A2(n_1144),
.B(n_1122),
.Y(n_1367)
);

HB1xp67_ASAP7_75t_L g1368 ( 
.A(n_1191),
.Y(n_1368)
);

AOI21xp5_ASAP7_75t_L g1369 ( 
.A1(n_1197),
.A2(n_1144),
.B(n_1122),
.Y(n_1369)
);

NAND2xp5_ASAP7_75t_L g1370 ( 
.A(n_1201),
.B(n_1212),
.Y(n_1370)
);

AOI221x1_ASAP7_75t_SL g1371 ( 
.A1(n_1261),
.A2(n_1130),
.B1(n_1168),
.B2(n_1161),
.C(n_1137),
.Y(n_1371)
);

AND2x2_ASAP7_75t_SL g1372 ( 
.A(n_1189),
.B(n_1275),
.Y(n_1372)
);

O2A1O1Ixp5_ASAP7_75t_L g1373 ( 
.A1(n_1194),
.A2(n_1288),
.B(n_1289),
.C(n_1282),
.Y(n_1373)
);

BUFx2_ASAP7_75t_L g1374 ( 
.A(n_1350),
.Y(n_1374)
);

AO21x2_ASAP7_75t_L g1375 ( 
.A1(n_1345),
.A2(n_1310),
.B(n_1367),
.Y(n_1375)
);

INVx2_ASAP7_75t_L g1376 ( 
.A(n_1340),
.Y(n_1376)
);

INVx1_ASAP7_75t_L g1377 ( 
.A(n_1334),
.Y(n_1377)
);

NOR2xp33_ASAP7_75t_L g1378 ( 
.A(n_1372),
.B(n_1303),
.Y(n_1378)
);

OAI21xp5_ASAP7_75t_L g1379 ( 
.A1(n_1373),
.A2(n_1308),
.B(n_1306),
.Y(n_1379)
);

INVx2_ASAP7_75t_L g1380 ( 
.A(n_1343),
.Y(n_1380)
);

OA21x2_ASAP7_75t_L g1381 ( 
.A1(n_1313),
.A2(n_1367),
.B(n_1369),
.Y(n_1381)
);

INVx2_ASAP7_75t_SL g1382 ( 
.A(n_1301),
.Y(n_1382)
);

INVx1_ASAP7_75t_L g1383 ( 
.A(n_1329),
.Y(n_1383)
);

AOI21xp5_ASAP7_75t_SL g1384 ( 
.A1(n_1306),
.A2(n_1299),
.B(n_1366),
.Y(n_1384)
);

INVx1_ASAP7_75t_L g1385 ( 
.A(n_1354),
.Y(n_1385)
);

INVx1_ASAP7_75t_L g1386 ( 
.A(n_1351),
.Y(n_1386)
);

INVx1_ASAP7_75t_L g1387 ( 
.A(n_1323),
.Y(n_1387)
);

INVx1_ASAP7_75t_L g1388 ( 
.A(n_1322),
.Y(n_1388)
);

INVx1_ASAP7_75t_L g1389 ( 
.A(n_1322),
.Y(n_1389)
);

AO21x2_ASAP7_75t_L g1390 ( 
.A1(n_1356),
.A2(n_1360),
.B(n_1353),
.Y(n_1390)
);

AND2x6_ASAP7_75t_L g1391 ( 
.A(n_1325),
.B(n_1348),
.Y(n_1391)
);

CKINVDCx5p33_ASAP7_75t_R g1392 ( 
.A(n_1311),
.Y(n_1392)
);

BUFx2_ASAP7_75t_SL g1393 ( 
.A(n_1346),
.Y(n_1393)
);

AND2x2_ASAP7_75t_L g1394 ( 
.A(n_1355),
.B(n_1357),
.Y(n_1394)
);

INVx1_ASAP7_75t_L g1395 ( 
.A(n_1307),
.Y(n_1395)
);

INVx1_ASAP7_75t_L g1396 ( 
.A(n_1349),
.Y(n_1396)
);

AND2x2_ASAP7_75t_L g1397 ( 
.A(n_1321),
.B(n_1332),
.Y(n_1397)
);

INVx1_ASAP7_75t_L g1398 ( 
.A(n_1349),
.Y(n_1398)
);

OR2x6_ASAP7_75t_L g1399 ( 
.A(n_1344),
.B(n_1320),
.Y(n_1399)
);

AND2x2_ASAP7_75t_L g1400 ( 
.A(n_1362),
.B(n_1358),
.Y(n_1400)
);

AO21x2_ASAP7_75t_L g1401 ( 
.A1(n_1341),
.A2(n_1365),
.B(n_1370),
.Y(n_1401)
);

INVx1_ASAP7_75t_L g1402 ( 
.A(n_1331),
.Y(n_1402)
);

OR2x2_ASAP7_75t_L g1403 ( 
.A(n_1362),
.B(n_1319),
.Y(n_1403)
);

OA21x2_ASAP7_75t_L g1404 ( 
.A1(n_1327),
.A2(n_1336),
.B(n_1335),
.Y(n_1404)
);

NAND2xp5_ASAP7_75t_L g1405 ( 
.A(n_1302),
.B(n_1371),
.Y(n_1405)
);

BUFx5_ASAP7_75t_L g1406 ( 
.A(n_1361),
.Y(n_1406)
);

INVx1_ASAP7_75t_L g1407 ( 
.A(n_1324),
.Y(n_1407)
);

NAND2xp5_ASAP7_75t_L g1408 ( 
.A(n_1368),
.B(n_1304),
.Y(n_1408)
);

BUFx3_ASAP7_75t_L g1409 ( 
.A(n_1337),
.Y(n_1409)
);

INVx2_ASAP7_75t_SL g1410 ( 
.A(n_1359),
.Y(n_1410)
);

AND2x2_ASAP7_75t_L g1411 ( 
.A(n_1342),
.B(n_1300),
.Y(n_1411)
);

INVx1_ASAP7_75t_L g1412 ( 
.A(n_1317),
.Y(n_1412)
);

BUFx2_ASAP7_75t_L g1413 ( 
.A(n_1337),
.Y(n_1413)
);

OA21x2_ASAP7_75t_L g1414 ( 
.A1(n_1338),
.A2(n_1309),
.B(n_1315),
.Y(n_1414)
);

BUFx2_ASAP7_75t_L g1415 ( 
.A(n_1374),
.Y(n_1415)
);

NAND2xp5_ASAP7_75t_L g1416 ( 
.A(n_1377),
.B(n_1380),
.Y(n_1416)
);

INVx1_ASAP7_75t_L g1417 ( 
.A(n_1376),
.Y(n_1417)
);

INVx1_ASAP7_75t_L g1418 ( 
.A(n_1376),
.Y(n_1418)
);

OR2x6_ASAP7_75t_L g1419 ( 
.A(n_1399),
.B(n_1305),
.Y(n_1419)
);

INVx1_ASAP7_75t_L g1420 ( 
.A(n_1376),
.Y(n_1420)
);

AND2x2_ASAP7_75t_L g1421 ( 
.A(n_1394),
.B(n_1364),
.Y(n_1421)
);

NAND2xp5_ASAP7_75t_L g1422 ( 
.A(n_1377),
.B(n_1314),
.Y(n_1422)
);

AND2x2_ASAP7_75t_L g1423 ( 
.A(n_1394),
.B(n_1312),
.Y(n_1423)
);

OR2x2_ASAP7_75t_L g1424 ( 
.A(n_1380),
.B(n_1363),
.Y(n_1424)
);

OR2x2_ASAP7_75t_L g1425 ( 
.A(n_1374),
.B(n_1385),
.Y(n_1425)
);

HB1xp67_ASAP7_75t_L g1426 ( 
.A(n_1385),
.Y(n_1426)
);

NAND2xp5_ASAP7_75t_L g1427 ( 
.A(n_1401),
.B(n_1388),
.Y(n_1427)
);

AND2x2_ASAP7_75t_L g1428 ( 
.A(n_1374),
.B(n_1305),
.Y(n_1428)
);

OAI21xp33_ASAP7_75t_L g1429 ( 
.A1(n_1384),
.A2(n_1333),
.B(n_1326),
.Y(n_1429)
);

BUFx3_ASAP7_75t_L g1430 ( 
.A(n_1391),
.Y(n_1430)
);

AND2x2_ASAP7_75t_L g1431 ( 
.A(n_1400),
.B(n_1318),
.Y(n_1431)
);

OR2x2_ASAP7_75t_L g1432 ( 
.A(n_1403),
.B(n_1330),
.Y(n_1432)
);

NAND2xp5_ASAP7_75t_L g1433 ( 
.A(n_1401),
.B(n_1347),
.Y(n_1433)
);

INVx2_ASAP7_75t_L g1434 ( 
.A(n_1410),
.Y(n_1434)
);

AOI22xp33_ASAP7_75t_L g1435 ( 
.A1(n_1378),
.A2(n_1316),
.B1(n_1328),
.B2(n_1348),
.Y(n_1435)
);

AND2x2_ASAP7_75t_L g1436 ( 
.A(n_1397),
.B(n_1352),
.Y(n_1436)
);

BUFx2_ASAP7_75t_L g1437 ( 
.A(n_1390),
.Y(n_1437)
);

AOI221xp5_ASAP7_75t_L g1438 ( 
.A1(n_1429),
.A2(n_1378),
.B1(n_1379),
.B2(n_1405),
.C(n_1408),
.Y(n_1438)
);

OR2x6_ASAP7_75t_L g1439 ( 
.A(n_1419),
.B(n_1399),
.Y(n_1439)
);

AOI221xp5_ASAP7_75t_L g1440 ( 
.A1(n_1429),
.A2(n_1379),
.B1(n_1405),
.B2(n_1408),
.C(n_1413),
.Y(n_1440)
);

BUFx2_ASAP7_75t_L g1441 ( 
.A(n_1430),
.Y(n_1441)
);

INVx1_ASAP7_75t_L g1442 ( 
.A(n_1417),
.Y(n_1442)
);

AOI22xp33_ASAP7_75t_L g1443 ( 
.A1(n_1419),
.A2(n_1401),
.B1(n_1409),
.B2(n_1413),
.Y(n_1443)
);

NAND2xp5_ASAP7_75t_L g1444 ( 
.A(n_1423),
.B(n_1401),
.Y(n_1444)
);

OR2x2_ASAP7_75t_L g1445 ( 
.A(n_1425),
.B(n_1403),
.Y(n_1445)
);

AOI33xp33_ASAP7_75t_L g1446 ( 
.A1(n_1435),
.A2(n_1412),
.A3(n_1407),
.B1(n_1402),
.B2(n_1387),
.B3(n_1389),
.Y(n_1446)
);

AOI22xp5_ASAP7_75t_L g1447 ( 
.A1(n_1435),
.A2(n_1413),
.B1(n_1409),
.B2(n_1401),
.Y(n_1447)
);

BUFx2_ASAP7_75t_L g1448 ( 
.A(n_1430),
.Y(n_1448)
);

AND2x2_ASAP7_75t_L g1449 ( 
.A(n_1415),
.B(n_1406),
.Y(n_1449)
);

INVx1_ASAP7_75t_L g1450 ( 
.A(n_1418),
.Y(n_1450)
);

INVxp67_ASAP7_75t_SL g1451 ( 
.A(n_1427),
.Y(n_1451)
);

AND2x4_ASAP7_75t_L g1452 ( 
.A(n_1430),
.B(n_1399),
.Y(n_1452)
);

AOI322xp5_ASAP7_75t_L g1453 ( 
.A1(n_1433),
.A2(n_1392),
.A3(n_1411),
.B1(n_1396),
.B2(n_1398),
.C1(n_1382),
.C2(n_1387),
.Y(n_1453)
);

AOI211xp5_ASAP7_75t_L g1454 ( 
.A1(n_1433),
.A2(n_1403),
.B(n_1398),
.C(n_1386),
.Y(n_1454)
);

AO21x2_ASAP7_75t_L g1455 ( 
.A1(n_1434),
.A2(n_1397),
.B(n_1375),
.Y(n_1455)
);

OAI211xp5_ASAP7_75t_SL g1456 ( 
.A1(n_1432),
.A2(n_1386),
.B(n_1383),
.C(n_1395),
.Y(n_1456)
);

HB1xp67_ASAP7_75t_L g1457 ( 
.A(n_1425),
.Y(n_1457)
);

INVx1_ASAP7_75t_L g1458 ( 
.A(n_1418),
.Y(n_1458)
);

AND2x2_ASAP7_75t_L g1459 ( 
.A(n_1415),
.B(n_1406),
.Y(n_1459)
);

BUFx3_ASAP7_75t_L g1460 ( 
.A(n_1424),
.Y(n_1460)
);

AND2x2_ASAP7_75t_L g1461 ( 
.A(n_1415),
.B(n_1406),
.Y(n_1461)
);

AND2x2_ASAP7_75t_L g1462 ( 
.A(n_1436),
.B(n_1406),
.Y(n_1462)
);

AOI22xp33_ASAP7_75t_L g1463 ( 
.A1(n_1419),
.A2(n_1428),
.B1(n_1414),
.B2(n_1432),
.Y(n_1463)
);

AND2x6_ASAP7_75t_SL g1464 ( 
.A(n_1419),
.B(n_1393),
.Y(n_1464)
);

HB1xp67_ASAP7_75t_L g1465 ( 
.A(n_1425),
.Y(n_1465)
);

NAND3xp33_ASAP7_75t_L g1466 ( 
.A(n_1432),
.B(n_1381),
.C(n_1404),
.Y(n_1466)
);

INVx1_ASAP7_75t_L g1467 ( 
.A(n_1420),
.Y(n_1467)
);

OR2x2_ASAP7_75t_L g1468 ( 
.A(n_1424),
.B(n_1416),
.Y(n_1468)
);

NAND4xp75_ASAP7_75t_L g1469 ( 
.A(n_1428),
.B(n_1381),
.C(n_1414),
.D(n_1404),
.Y(n_1469)
);

BUFx2_ASAP7_75t_L g1470 ( 
.A(n_1464),
.Y(n_1470)
);

INVx2_ASAP7_75t_L g1471 ( 
.A(n_1455),
.Y(n_1471)
);

INVx2_ASAP7_75t_L g1472 ( 
.A(n_1455),
.Y(n_1472)
);

INVx2_ASAP7_75t_SL g1473 ( 
.A(n_1441),
.Y(n_1473)
);

NAND2xp5_ASAP7_75t_L g1474 ( 
.A(n_1451),
.B(n_1426),
.Y(n_1474)
);

INVx4_ASAP7_75t_SL g1475 ( 
.A(n_1439),
.Y(n_1475)
);

INVx1_ASAP7_75t_L g1476 ( 
.A(n_1442),
.Y(n_1476)
);

NAND2xp5_ASAP7_75t_SL g1477 ( 
.A(n_1446),
.B(n_1428),
.Y(n_1477)
);

BUFx2_ASAP7_75t_L g1478 ( 
.A(n_1464),
.Y(n_1478)
);

NAND2xp5_ASAP7_75t_L g1479 ( 
.A(n_1444),
.B(n_1423),
.Y(n_1479)
);

INVx2_ASAP7_75t_SL g1480 ( 
.A(n_1441),
.Y(n_1480)
);

BUFx2_ASAP7_75t_L g1481 ( 
.A(n_1439),
.Y(n_1481)
);

HB1xp67_ASAP7_75t_L g1482 ( 
.A(n_1457),
.Y(n_1482)
);

NAND2xp5_ASAP7_75t_L g1483 ( 
.A(n_1454),
.B(n_1468),
.Y(n_1483)
);

HB1xp67_ASAP7_75t_L g1484 ( 
.A(n_1465),
.Y(n_1484)
);

OA21x2_ASAP7_75t_L g1485 ( 
.A1(n_1469),
.A2(n_1437),
.B(n_1434),
.Y(n_1485)
);

HB1xp67_ASAP7_75t_L g1486 ( 
.A(n_1450),
.Y(n_1486)
);

NAND2xp5_ASAP7_75t_SL g1487 ( 
.A(n_1447),
.B(n_1431),
.Y(n_1487)
);

HB1xp67_ASAP7_75t_L g1488 ( 
.A(n_1450),
.Y(n_1488)
);

AND2x2_ASAP7_75t_L g1489 ( 
.A(n_1449),
.B(n_1459),
.Y(n_1489)
);

NOR2xp33_ASAP7_75t_L g1490 ( 
.A(n_1438),
.B(n_1421),
.Y(n_1490)
);

INVx1_ASAP7_75t_L g1491 ( 
.A(n_1486),
.Y(n_1491)
);

NAND2xp5_ASAP7_75t_L g1492 ( 
.A(n_1490),
.B(n_1445),
.Y(n_1492)
);

AND2x4_ASAP7_75t_SL g1493 ( 
.A(n_1482),
.B(n_1439),
.Y(n_1493)
);

AND2x2_ASAP7_75t_L g1494 ( 
.A(n_1470),
.B(n_1462),
.Y(n_1494)
);

INVx1_ASAP7_75t_L g1495 ( 
.A(n_1486),
.Y(n_1495)
);

AND2x2_ASAP7_75t_L g1496 ( 
.A(n_1470),
.B(n_1462),
.Y(n_1496)
);

INVx1_ASAP7_75t_L g1497 ( 
.A(n_1488),
.Y(n_1497)
);

INVx1_ASAP7_75t_L g1498 ( 
.A(n_1488),
.Y(n_1498)
);

INVx1_ASAP7_75t_L g1499 ( 
.A(n_1476),
.Y(n_1499)
);

INVx2_ASAP7_75t_L g1500 ( 
.A(n_1471),
.Y(n_1500)
);

AND2x4_ASAP7_75t_L g1501 ( 
.A(n_1475),
.B(n_1452),
.Y(n_1501)
);

INVx2_ASAP7_75t_L g1502 ( 
.A(n_1471),
.Y(n_1502)
);

INVx2_ASAP7_75t_L g1503 ( 
.A(n_1471),
.Y(n_1503)
);

AND2x2_ASAP7_75t_L g1504 ( 
.A(n_1470),
.B(n_1448),
.Y(n_1504)
);

HB1xp67_ASAP7_75t_L g1505 ( 
.A(n_1482),
.Y(n_1505)
);

AND2x2_ASAP7_75t_L g1506 ( 
.A(n_1478),
.B(n_1452),
.Y(n_1506)
);

OR2x2_ASAP7_75t_L g1507 ( 
.A(n_1483),
.B(n_1445),
.Y(n_1507)
);

NAND2xp5_ASAP7_75t_L g1508 ( 
.A(n_1490),
.B(n_1453),
.Y(n_1508)
);

AND2x2_ASAP7_75t_L g1509 ( 
.A(n_1478),
.B(n_1452),
.Y(n_1509)
);

OR2x2_ASAP7_75t_L g1510 ( 
.A(n_1483),
.B(n_1468),
.Y(n_1510)
);

INVxp67_ASAP7_75t_SL g1511 ( 
.A(n_1484),
.Y(n_1511)
);

AND2x2_ASAP7_75t_L g1512 ( 
.A(n_1478),
.B(n_1459),
.Y(n_1512)
);

OAI33xp33_ASAP7_75t_L g1513 ( 
.A1(n_1487),
.A2(n_1466),
.A3(n_1456),
.B1(n_1422),
.B2(n_1458),
.B3(n_1467),
.Y(n_1513)
);

INVx1_ASAP7_75t_L g1514 ( 
.A(n_1476),
.Y(n_1514)
);

AND2x2_ASAP7_75t_L g1515 ( 
.A(n_1481),
.B(n_1461),
.Y(n_1515)
);

AND2x2_ASAP7_75t_L g1516 ( 
.A(n_1481),
.B(n_1461),
.Y(n_1516)
);

INVx2_ASAP7_75t_L g1517 ( 
.A(n_1471),
.Y(n_1517)
);

NAND2xp5_ASAP7_75t_SL g1518 ( 
.A(n_1477),
.B(n_1453),
.Y(n_1518)
);

INVx2_ASAP7_75t_L g1519 ( 
.A(n_1472),
.Y(n_1519)
);

INVx1_ASAP7_75t_SL g1520 ( 
.A(n_1473),
.Y(n_1520)
);

NOR2xp33_ASAP7_75t_R g1521 ( 
.A(n_1473),
.B(n_1339),
.Y(n_1521)
);

INVx6_ASAP7_75t_L g1522 ( 
.A(n_1475),
.Y(n_1522)
);

OR2x2_ASAP7_75t_L g1523 ( 
.A(n_1479),
.B(n_1460),
.Y(n_1523)
);

NAND2xp5_ASAP7_75t_L g1524 ( 
.A(n_1477),
.B(n_1421),
.Y(n_1524)
);

NAND3xp33_ASAP7_75t_L g1525 ( 
.A(n_1487),
.B(n_1440),
.C(n_1447),
.Y(n_1525)
);

INVx2_ASAP7_75t_L g1526 ( 
.A(n_1472),
.Y(n_1526)
);

INVx1_ASAP7_75t_L g1527 ( 
.A(n_1505),
.Y(n_1527)
);

INVx1_ASAP7_75t_L g1528 ( 
.A(n_1505),
.Y(n_1528)
);

AND2x2_ASAP7_75t_L g1529 ( 
.A(n_1504),
.B(n_1489),
.Y(n_1529)
);

INVx1_ASAP7_75t_L g1530 ( 
.A(n_1499),
.Y(n_1530)
);

OR2x2_ASAP7_75t_L g1531 ( 
.A(n_1507),
.B(n_1484),
.Y(n_1531)
);

NAND2xp5_ASAP7_75t_L g1532 ( 
.A(n_1508),
.B(n_1489),
.Y(n_1532)
);

NAND2xp5_ASAP7_75t_L g1533 ( 
.A(n_1508),
.B(n_1489),
.Y(n_1533)
);

INVx1_ASAP7_75t_L g1534 ( 
.A(n_1499),
.Y(n_1534)
);

NAND2xp5_ASAP7_75t_L g1535 ( 
.A(n_1518),
.B(n_1473),
.Y(n_1535)
);

INVx1_ASAP7_75t_L g1536 ( 
.A(n_1514),
.Y(n_1536)
);

INVx1_ASAP7_75t_L g1537 ( 
.A(n_1514),
.Y(n_1537)
);

AND2x2_ASAP7_75t_L g1538 ( 
.A(n_1504),
.B(n_1481),
.Y(n_1538)
);

INVx1_ASAP7_75t_L g1539 ( 
.A(n_1511),
.Y(n_1539)
);

INVx1_ASAP7_75t_L g1540 ( 
.A(n_1511),
.Y(n_1540)
);

OR2x2_ASAP7_75t_L g1541 ( 
.A(n_1507),
.B(n_1474),
.Y(n_1541)
);

INVx2_ASAP7_75t_L g1542 ( 
.A(n_1520),
.Y(n_1542)
);

INVx1_ASAP7_75t_L g1543 ( 
.A(n_1491),
.Y(n_1543)
);

AND2x2_ASAP7_75t_L g1544 ( 
.A(n_1494),
.B(n_1475),
.Y(n_1544)
);

AND2x2_ASAP7_75t_L g1545 ( 
.A(n_1494),
.B(n_1475),
.Y(n_1545)
);

INVx1_ASAP7_75t_L g1546 ( 
.A(n_1491),
.Y(n_1546)
);

INVx1_ASAP7_75t_L g1547 ( 
.A(n_1495),
.Y(n_1547)
);

AND2x4_ASAP7_75t_L g1548 ( 
.A(n_1506),
.B(n_1475),
.Y(n_1548)
);

OAI21xp33_ASAP7_75t_L g1549 ( 
.A1(n_1525),
.A2(n_1443),
.B(n_1463),
.Y(n_1549)
);

INVx1_ASAP7_75t_L g1550 ( 
.A(n_1495),
.Y(n_1550)
);

NAND2xp5_ASAP7_75t_L g1551 ( 
.A(n_1512),
.B(n_1480),
.Y(n_1551)
);

INVx2_ASAP7_75t_L g1552 ( 
.A(n_1520),
.Y(n_1552)
);

INVx1_ASAP7_75t_L g1553 ( 
.A(n_1497),
.Y(n_1553)
);

INVx2_ASAP7_75t_SL g1554 ( 
.A(n_1522),
.Y(n_1554)
);

INVx1_ASAP7_75t_SL g1555 ( 
.A(n_1506),
.Y(n_1555)
);

NAND2xp5_ASAP7_75t_L g1556 ( 
.A(n_1512),
.B(n_1480),
.Y(n_1556)
);

INVx1_ASAP7_75t_L g1557 ( 
.A(n_1497),
.Y(n_1557)
);

AND2x2_ASAP7_75t_L g1558 ( 
.A(n_1494),
.B(n_1475),
.Y(n_1558)
);

OAI211xp5_ASAP7_75t_L g1559 ( 
.A1(n_1525),
.A2(n_1492),
.B(n_1496),
.C(n_1485),
.Y(n_1559)
);

INVx1_ASAP7_75t_L g1560 ( 
.A(n_1498),
.Y(n_1560)
);

INVx2_ASAP7_75t_L g1561 ( 
.A(n_1526),
.Y(n_1561)
);

OAI22xp5_ASAP7_75t_L g1562 ( 
.A1(n_1549),
.A2(n_1524),
.B1(n_1522),
.B2(n_1492),
.Y(n_1562)
);

INVx1_ASAP7_75t_SL g1563 ( 
.A(n_1538),
.Y(n_1563)
);

AND2x4_ASAP7_75t_L g1564 ( 
.A(n_1544),
.B(n_1509),
.Y(n_1564)
);

INVx1_ASAP7_75t_L g1565 ( 
.A(n_1539),
.Y(n_1565)
);

HB1xp67_ASAP7_75t_L g1566 ( 
.A(n_1529),
.Y(n_1566)
);

INVx2_ASAP7_75t_L g1567 ( 
.A(n_1529),
.Y(n_1567)
);

OR2x2_ASAP7_75t_L g1568 ( 
.A(n_1531),
.B(n_1510),
.Y(n_1568)
);

INVx1_ASAP7_75t_L g1569 ( 
.A(n_1539),
.Y(n_1569)
);

INVx1_ASAP7_75t_L g1570 ( 
.A(n_1540),
.Y(n_1570)
);

AND2x2_ASAP7_75t_L g1571 ( 
.A(n_1538),
.B(n_1544),
.Y(n_1571)
);

INVx3_ASAP7_75t_L g1572 ( 
.A(n_1548),
.Y(n_1572)
);

NAND2xp5_ASAP7_75t_L g1573 ( 
.A(n_1555),
.B(n_1512),
.Y(n_1573)
);

HB1xp67_ASAP7_75t_L g1574 ( 
.A(n_1531),
.Y(n_1574)
);

NAND2xp5_ASAP7_75t_L g1575 ( 
.A(n_1535),
.B(n_1496),
.Y(n_1575)
);

INVx2_ASAP7_75t_L g1576 ( 
.A(n_1545),
.Y(n_1576)
);

INVx2_ASAP7_75t_L g1577 ( 
.A(n_1545),
.Y(n_1577)
);

INVxp67_ASAP7_75t_L g1578 ( 
.A(n_1554),
.Y(n_1578)
);

CKINVDCx16_ASAP7_75t_R g1579 ( 
.A(n_1558),
.Y(n_1579)
);

INVx1_ASAP7_75t_L g1580 ( 
.A(n_1540),
.Y(n_1580)
);

NOR2x1_ASAP7_75t_L g1581 ( 
.A(n_1559),
.B(n_1498),
.Y(n_1581)
);

AND2x2_ASAP7_75t_L g1582 ( 
.A(n_1558),
.B(n_1496),
.Y(n_1582)
);

BUFx2_ASAP7_75t_L g1583 ( 
.A(n_1548),
.Y(n_1583)
);

OAI22xp5_ASAP7_75t_L g1584 ( 
.A1(n_1532),
.A2(n_1524),
.B1(n_1522),
.B2(n_1469),
.Y(n_1584)
);

OR2x2_ASAP7_75t_L g1585 ( 
.A(n_1528),
.B(n_1510),
.Y(n_1585)
);

INVx1_ASAP7_75t_L g1586 ( 
.A(n_1527),
.Y(n_1586)
);

NAND2xp5_ASAP7_75t_L g1587 ( 
.A(n_1579),
.B(n_1533),
.Y(n_1587)
);

OAI22xp33_ASAP7_75t_SL g1588 ( 
.A1(n_1581),
.A2(n_1522),
.B1(n_1554),
.B2(n_1548),
.Y(n_1588)
);

INVxp67_ASAP7_75t_SL g1589 ( 
.A(n_1581),
.Y(n_1589)
);

INVx1_ASAP7_75t_L g1590 ( 
.A(n_1574),
.Y(n_1590)
);

INVx1_ASAP7_75t_L g1591 ( 
.A(n_1566),
.Y(n_1591)
);

INVx1_ASAP7_75t_L g1592 ( 
.A(n_1565),
.Y(n_1592)
);

INVx1_ASAP7_75t_L g1593 ( 
.A(n_1565),
.Y(n_1593)
);

AOI21xp5_ASAP7_75t_L g1594 ( 
.A1(n_1562),
.A2(n_1513),
.B(n_1551),
.Y(n_1594)
);

AND2x2_ASAP7_75t_L g1595 ( 
.A(n_1571),
.B(n_1509),
.Y(n_1595)
);

AO21x1_ASAP7_75t_L g1596 ( 
.A1(n_1569),
.A2(n_1527),
.B(n_1542),
.Y(n_1596)
);

INVx1_ASAP7_75t_L g1597 ( 
.A(n_1569),
.Y(n_1597)
);

NAND2xp5_ASAP7_75t_L g1598 ( 
.A(n_1579),
.B(n_1542),
.Y(n_1598)
);

AOI22xp33_ASAP7_75t_L g1599 ( 
.A1(n_1584),
.A2(n_1522),
.B1(n_1513),
.B2(n_1501),
.Y(n_1599)
);

AOI22xp5_ASAP7_75t_L g1600 ( 
.A1(n_1571),
.A2(n_1501),
.B1(n_1556),
.B2(n_1552),
.Y(n_1600)
);

AOI22xp33_ASAP7_75t_L g1601 ( 
.A1(n_1575),
.A2(n_1552),
.B1(n_1485),
.B2(n_1557),
.Y(n_1601)
);

OAI31xp33_ASAP7_75t_L g1602 ( 
.A1(n_1563),
.A2(n_1493),
.A3(n_1541),
.B(n_1501),
.Y(n_1602)
);

NOR3xp33_ASAP7_75t_SL g1603 ( 
.A(n_1586),
.B(n_1546),
.C(n_1543),
.Y(n_1603)
);

NAND2xp5_ASAP7_75t_L g1604 ( 
.A(n_1576),
.B(n_1547),
.Y(n_1604)
);

INVx1_ASAP7_75t_L g1605 ( 
.A(n_1570),
.Y(n_1605)
);

NAND2xp33_ASAP7_75t_R g1606 ( 
.A(n_1603),
.B(n_1583),
.Y(n_1606)
);

AND2x4_ASAP7_75t_L g1607 ( 
.A(n_1590),
.B(n_1583),
.Y(n_1607)
);

OR2x2_ASAP7_75t_L g1608 ( 
.A(n_1587),
.B(n_1598),
.Y(n_1608)
);

INVx1_ASAP7_75t_SL g1609 ( 
.A(n_1595),
.Y(n_1609)
);

INVx2_ASAP7_75t_L g1610 ( 
.A(n_1591),
.Y(n_1610)
);

NAND2xp5_ASAP7_75t_L g1611 ( 
.A(n_1589),
.B(n_1576),
.Y(n_1611)
);

NOR2xp33_ASAP7_75t_L g1612 ( 
.A(n_1600),
.B(n_1577),
.Y(n_1612)
);

INVx1_ASAP7_75t_L g1613 ( 
.A(n_1589),
.Y(n_1613)
);

AND2x2_ASAP7_75t_L g1614 ( 
.A(n_1602),
.B(n_1564),
.Y(n_1614)
);

OR2x2_ASAP7_75t_L g1615 ( 
.A(n_1604),
.B(n_1568),
.Y(n_1615)
);

NAND2xp5_ASAP7_75t_L g1616 ( 
.A(n_1594),
.B(n_1577),
.Y(n_1616)
);

NOR2xp33_ASAP7_75t_L g1617 ( 
.A(n_1588),
.B(n_1572),
.Y(n_1617)
);

NOR2x1_ASAP7_75t_L g1618 ( 
.A(n_1613),
.B(n_1592),
.Y(n_1618)
);

AOI22xp5_ASAP7_75t_L g1619 ( 
.A1(n_1606),
.A2(n_1564),
.B1(n_1596),
.B2(n_1614),
.Y(n_1619)
);

O2A1O1Ixp33_ASAP7_75t_SL g1620 ( 
.A1(n_1616),
.A2(n_1578),
.B(n_1572),
.C(n_1586),
.Y(n_1620)
);

O2A1O1Ixp33_ASAP7_75t_L g1621 ( 
.A1(n_1611),
.A2(n_1603),
.B(n_1605),
.C(n_1593),
.Y(n_1621)
);

AOI31xp33_ASAP7_75t_L g1622 ( 
.A1(n_1608),
.A2(n_1599),
.A3(n_1568),
.B(n_1597),
.Y(n_1622)
);

NAND2xp33_ASAP7_75t_SL g1623 ( 
.A(n_1615),
.B(n_1572),
.Y(n_1623)
);

OAI211xp5_ASAP7_75t_SL g1624 ( 
.A1(n_1609),
.A2(n_1601),
.B(n_1570),
.C(n_1580),
.Y(n_1624)
);

O2A1O1Ixp33_ASAP7_75t_L g1625 ( 
.A1(n_1617),
.A2(n_1580),
.B(n_1601),
.C(n_1585),
.Y(n_1625)
);

AOI22xp33_ASAP7_75t_L g1626 ( 
.A1(n_1612),
.A2(n_1564),
.B1(n_1582),
.B2(n_1567),
.Y(n_1626)
);

NAND2xp33_ASAP7_75t_L g1627 ( 
.A(n_1610),
.B(n_1585),
.Y(n_1627)
);

A2O1A1Ixp33_ASAP7_75t_L g1628 ( 
.A1(n_1621),
.A2(n_1607),
.B(n_1582),
.C(n_1573),
.Y(n_1628)
);

AOI322xp5_ASAP7_75t_L g1629 ( 
.A1(n_1619),
.A2(n_1607),
.A3(n_1567),
.B1(n_1550),
.B2(n_1560),
.C1(n_1553),
.C2(n_1516),
.Y(n_1629)
);

INVx1_ASAP7_75t_SL g1630 ( 
.A(n_1623),
.Y(n_1630)
);

INVx1_ASAP7_75t_L g1631 ( 
.A(n_1627),
.Y(n_1631)
);

OAI21xp5_ASAP7_75t_L g1632 ( 
.A1(n_1625),
.A2(n_1622),
.B(n_1624),
.Y(n_1632)
);

INVxp67_ASAP7_75t_L g1633 ( 
.A(n_1631),
.Y(n_1633)
);

INVxp67_ASAP7_75t_L g1634 ( 
.A(n_1630),
.Y(n_1634)
);

INVx1_ASAP7_75t_L g1635 ( 
.A(n_1628),
.Y(n_1635)
);

AND2x2_ASAP7_75t_L g1636 ( 
.A(n_1629),
.B(n_1626),
.Y(n_1636)
);

INVx1_ASAP7_75t_L g1637 ( 
.A(n_1632),
.Y(n_1637)
);

AND2x2_ASAP7_75t_L g1638 ( 
.A(n_1631),
.B(n_1618),
.Y(n_1638)
);

INVx1_ASAP7_75t_L g1639 ( 
.A(n_1638),
.Y(n_1639)
);

INVx1_ASAP7_75t_L g1640 ( 
.A(n_1634),
.Y(n_1640)
);

OAI211xp5_ASAP7_75t_SL g1641 ( 
.A1(n_1637),
.A2(n_1620),
.B(n_1541),
.C(n_1561),
.Y(n_1641)
);

AOI21xp33_ASAP7_75t_L g1642 ( 
.A1(n_1635),
.A2(n_1536),
.B(n_1534),
.Y(n_1642)
);

INVx1_ASAP7_75t_SL g1643 ( 
.A(n_1636),
.Y(n_1643)
);

O2A1O1Ixp33_ASAP7_75t_SL g1644 ( 
.A1(n_1643),
.A2(n_1633),
.B(n_1534),
.C(n_1537),
.Y(n_1644)
);

NAND3xp33_ASAP7_75t_SL g1645 ( 
.A(n_1640),
.B(n_1633),
.C(n_1521),
.Y(n_1645)
);

INVx2_ASAP7_75t_L g1646 ( 
.A(n_1639),
.Y(n_1646)
);

NAND4xp75_ASAP7_75t_L g1647 ( 
.A(n_1646),
.B(n_1642),
.C(n_1645),
.D(n_1644),
.Y(n_1647)
);

HB1xp67_ASAP7_75t_L g1648 ( 
.A(n_1647),
.Y(n_1648)
);

INVx2_ASAP7_75t_L g1649 ( 
.A(n_1648),
.Y(n_1649)
);

NOR3xp33_ASAP7_75t_L g1650 ( 
.A(n_1648),
.B(n_1641),
.C(n_1537),
.Y(n_1650)
);

NAND2xp5_ASAP7_75t_L g1651 ( 
.A(n_1650),
.B(n_1530),
.Y(n_1651)
);

INVx2_ASAP7_75t_L g1652 ( 
.A(n_1649),
.Y(n_1652)
);

AOI22xp5_ASAP7_75t_L g1653 ( 
.A1(n_1652),
.A2(n_1561),
.B1(n_1536),
.B2(n_1501),
.Y(n_1653)
);

INVx1_ASAP7_75t_L g1654 ( 
.A(n_1651),
.Y(n_1654)
);

XOR2xp5_ASAP7_75t_L g1655 ( 
.A(n_1654),
.B(n_1523),
.Y(n_1655)
);

AOI22xp5_ASAP7_75t_L g1656 ( 
.A1(n_1655),
.A2(n_1653),
.B1(n_1526),
.B2(n_1502),
.Y(n_1656)
);

NAND2xp33_ASAP7_75t_L g1657 ( 
.A(n_1656),
.B(n_1515),
.Y(n_1657)
);

XNOR2xp5_ASAP7_75t_L g1658 ( 
.A(n_1657),
.B(n_1515),
.Y(n_1658)
);

AOI221xp5_ASAP7_75t_SL g1659 ( 
.A1(n_1658),
.A2(n_1526),
.B1(n_1519),
.B2(n_1500),
.C(n_1502),
.Y(n_1659)
);

AOI211xp5_ASAP7_75t_L g1660 ( 
.A1(n_1659),
.A2(n_1502),
.B(n_1503),
.C(n_1517),
.Y(n_1660)
);


endmodule