module fake_jpeg_25311_n_197 (n_3, n_2, n_1, n_0, n_10, n_4, n_8, n_9, n_6, n_5, n_7, n_197);

input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_197;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_14;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_84;
wire n_59;
wire n_98;
wire n_178;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_13;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_186;
wire n_24;
wire n_44;
wire n_143;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_11;
wire n_131;
wire n_56;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_12;
wire n_132;
wire n_133;
wire n_67;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_161;
wire n_22;
wire n_138;
wire n_101;
wire n_48;
wire n_35;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_189;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

INVx1_ASAP7_75t_L g11 ( 
.A(n_10),
.Y(n_11)
);

CKINVDCx20_ASAP7_75t_R g12 ( 
.A(n_4),
.Y(n_12)
);

BUFx5_ASAP7_75t_L g13 ( 
.A(n_5),
.Y(n_13)
);

BUFx10_ASAP7_75t_L g14 ( 
.A(n_2),
.Y(n_14)
);

BUFx6f_ASAP7_75t_L g15 ( 
.A(n_0),
.Y(n_15)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_6),
.Y(n_16)
);

INVx2_ASAP7_75t_L g17 ( 
.A(n_10),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_6),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_0),
.Y(n_19)
);

INVx2_ASAP7_75t_L g20 ( 
.A(n_10),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_2),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_9),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_22),
.Y(n_23)
);

NAND2xp5_ASAP7_75t_SL g36 ( 
.A(n_23),
.B(n_25),
.Y(n_36)
);

NAND2xp5_ASAP7_75t_L g24 ( 
.A(n_17),
.B(n_0),
.Y(n_24)
);

NAND2xp5_ASAP7_75t_L g41 ( 
.A(n_24),
.B(n_14),
.Y(n_41)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_14),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_14),
.Y(n_26)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_26),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_22),
.Y(n_27)
);

OR2x2_ASAP7_75t_L g33 ( 
.A(n_27),
.B(n_28),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_L g28 ( 
.A(n_17),
.B(n_9),
.Y(n_28)
);

INVx5_ASAP7_75t_L g29 ( 
.A(n_14),
.Y(n_29)
);

INVx4_ASAP7_75t_L g40 ( 
.A(n_29),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_17),
.Y(n_30)
);

INVx2_ASAP7_75t_L g35 ( 
.A(n_30),
.Y(n_35)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_14),
.Y(n_31)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_31),
.Y(n_42)
);

A2O1A1Ixp33_ASAP7_75t_L g32 ( 
.A1(n_24),
.A2(n_11),
.B(n_16),
.C(n_19),
.Y(n_32)
);

NOR2xp33_ASAP7_75t_L g43 ( 
.A(n_32),
.B(n_28),
.Y(n_43)
);

NAND2xp33_ASAP7_75t_SL g34 ( 
.A(n_24),
.B(n_13),
.Y(n_34)
);

OR2x2_ASAP7_75t_L g57 ( 
.A(n_34),
.B(n_13),
.Y(n_57)
);

AOI22xp33_ASAP7_75t_SL g38 ( 
.A1(n_29),
.A2(n_20),
.B1(n_12),
.B2(n_11),
.Y(n_38)
);

AOI22xp33_ASAP7_75t_SL g52 ( 
.A1(n_38),
.A2(n_16),
.B1(n_11),
.B2(n_12),
.Y(n_52)
);

OAI22xp33_ASAP7_75t_SL g39 ( 
.A1(n_29),
.A2(n_20),
.B1(n_21),
.B2(n_15),
.Y(n_39)
);

OAI22xp5_ASAP7_75t_L g47 ( 
.A1(n_39),
.A2(n_31),
.B1(n_25),
.B2(n_26),
.Y(n_47)
);

NAND2xp5_ASAP7_75t_L g44 ( 
.A(n_41),
.B(n_30),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_SL g61 ( 
.A(n_43),
.B(n_50),
.Y(n_61)
);

AND2x2_ASAP7_75t_L g78 ( 
.A(n_44),
.B(n_47),
.Y(n_78)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_36),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_45),
.B(n_56),
.Y(n_67)
);

HB1xp67_ASAP7_75t_L g46 ( 
.A(n_40),
.Y(n_46)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_46),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_L g48 ( 
.A(n_41),
.B(n_30),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_SL g62 ( 
.A(n_48),
.B(n_33),
.Y(n_62)
);

OAI22xp5_ASAP7_75t_L g49 ( 
.A1(n_41),
.A2(n_20),
.B1(n_31),
.B2(n_26),
.Y(n_49)
);

OAI22xp5_ASAP7_75t_SL g68 ( 
.A1(n_49),
.A2(n_51),
.B1(n_54),
.B2(n_33),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_33),
.B(n_27),
.Y(n_50)
);

OAI22xp5_ASAP7_75t_L g51 ( 
.A1(n_38),
.A2(n_25),
.B1(n_27),
.B2(n_23),
.Y(n_51)
);

OAI22xp5_ASAP7_75t_L g66 ( 
.A1(n_52),
.A2(n_18),
.B1(n_42),
.B2(n_37),
.Y(n_66)
);

INVx4_ASAP7_75t_L g53 ( 
.A(n_40),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_53),
.Y(n_65)
);

AOI22xp33_ASAP7_75t_SL g54 ( 
.A1(n_40),
.A2(n_16),
.B1(n_18),
.B2(n_19),
.Y(n_54)
);

INVx6_ASAP7_75t_L g55 ( 
.A(n_35),
.Y(n_55)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_55),
.Y(n_76)
);

INVx4_ASAP7_75t_SL g56 ( 
.A(n_37),
.Y(n_56)
);

AOI21xp5_ASAP7_75t_L g64 ( 
.A1(n_57),
.A2(n_32),
.B(n_33),
.Y(n_64)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_35),
.Y(n_58)
);

BUFx3_ASAP7_75t_L g73 ( 
.A(n_58),
.Y(n_73)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_36),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_59),
.B(n_60),
.Y(n_69)
);

INVx1_ASAP7_75t_SL g60 ( 
.A(n_37),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_L g94 ( 
.A(n_62),
.B(n_30),
.Y(n_94)
);

OAI21xp5_ASAP7_75t_L g100 ( 
.A1(n_64),
.A2(n_75),
.B(n_61),
.Y(n_100)
);

AOI22xp5_ASAP7_75t_L g86 ( 
.A1(n_66),
.A2(n_68),
.B1(n_74),
.B2(n_49),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_45),
.B(n_23),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_SL g95 ( 
.A(n_70),
.B(n_71),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_50),
.B(n_42),
.Y(n_71)
);

INVxp67_ASAP7_75t_L g72 ( 
.A(n_54),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_72),
.B(n_79),
.Y(n_83)
);

OAI22xp5_ASAP7_75t_SL g74 ( 
.A1(n_44),
.A2(n_35),
.B1(n_42),
.B2(n_39),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_SL g75 ( 
.A(n_43),
.B(n_32),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_SL g91 ( 
.A(n_75),
.B(n_77),
.Y(n_91)
);

CKINVDCx20_ASAP7_75t_R g77 ( 
.A(n_46),
.Y(n_77)
);

CKINVDCx20_ASAP7_75t_R g79 ( 
.A(n_47),
.Y(n_79)
);

BUFx3_ASAP7_75t_L g80 ( 
.A(n_53),
.Y(n_80)
);

INVx11_ASAP7_75t_L g102 ( 
.A(n_80),
.Y(n_102)
);

INVx4_ASAP7_75t_L g81 ( 
.A(n_53),
.Y(n_81)
);

CKINVDCx14_ASAP7_75t_R g98 ( 
.A(n_81),
.Y(n_98)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_67),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_L g112 ( 
.A(n_82),
.B(n_87),
.Y(n_112)
);

OAI22xp5_ASAP7_75t_L g84 ( 
.A1(n_79),
.A2(n_52),
.B1(n_59),
.B2(n_51),
.Y(n_84)
);

AOI22xp5_ASAP7_75t_L g125 ( 
.A1(n_84),
.A2(n_96),
.B1(n_0),
.B2(n_1),
.Y(n_125)
);

MAJx2_ASAP7_75t_L g85 ( 
.A(n_64),
.B(n_57),
.C(n_48),
.Y(n_85)
);

MAJIxp5_ASAP7_75t_L g122 ( 
.A(n_85),
.B(n_88),
.C(n_73),
.Y(n_122)
);

OAI22xp5_ASAP7_75t_L g115 ( 
.A1(n_86),
.A2(n_90),
.B1(n_101),
.B2(n_89),
.Y(n_115)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_67),
.Y(n_87)
);

MAJIxp5_ASAP7_75t_L g88 ( 
.A(n_62),
.B(n_57),
.C(n_60),
.Y(n_88)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_74),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g116 ( 
.A(n_89),
.B(n_92),
.Y(n_116)
);

AOI22xp5_ASAP7_75t_L g90 ( 
.A1(n_78),
.A2(n_56),
.B1(n_60),
.B2(n_55),
.Y(n_90)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_69),
.Y(n_92)
);

NAND2xp33_ASAP7_75t_SL g93 ( 
.A(n_68),
.B(n_56),
.Y(n_93)
);

OAI21xp5_ASAP7_75t_SL g108 ( 
.A1(n_93),
.A2(n_103),
.B(n_104),
.Y(n_108)
);

AO21x1_ASAP7_75t_L g124 ( 
.A1(n_94),
.A2(n_100),
.B(n_73),
.Y(n_124)
);

OAI22xp5_ASAP7_75t_L g96 ( 
.A1(n_61),
.A2(n_55),
.B1(n_58),
.B2(n_21),
.Y(n_96)
);

INVxp67_ASAP7_75t_L g97 ( 
.A(n_66),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g119 ( 
.A(n_97),
.B(n_99),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_78),
.B(n_14),
.Y(n_99)
);

AOI22xp5_ASAP7_75t_L g101 ( 
.A1(n_78),
.A2(n_21),
.B1(n_15),
.B2(n_13),
.Y(n_101)
);

AOI22xp5_ASAP7_75t_SL g103 ( 
.A1(n_70),
.A2(n_21),
.B1(n_15),
.B2(n_9),
.Y(n_103)
);

INVxp67_ASAP7_75t_L g104 ( 
.A(n_69),
.Y(n_104)
);

INVx3_ASAP7_75t_L g105 ( 
.A(n_65),
.Y(n_105)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_105),
.Y(n_113)
);

XOR2xp5_ASAP7_75t_L g106 ( 
.A(n_88),
.B(n_100),
.Y(n_106)
);

XOR2xp5_ASAP7_75t_L g131 ( 
.A(n_106),
.B(n_107),
.Y(n_131)
);

XNOR2xp5_ASAP7_75t_SL g107 ( 
.A(n_85),
.B(n_99),
.Y(n_107)
);

OAI21xp5_ASAP7_75t_L g109 ( 
.A1(n_83),
.A2(n_71),
.B(n_77),
.Y(n_109)
);

AOI21xp5_ASAP7_75t_SL g139 ( 
.A1(n_109),
.A2(n_110),
.B(n_117),
.Y(n_139)
);

OAI21xp5_ASAP7_75t_SL g110 ( 
.A1(n_97),
.A2(n_63),
.B(n_76),
.Y(n_110)
);

XOR2xp5_ASAP7_75t_L g111 ( 
.A(n_86),
.B(n_63),
.Y(n_111)
);

XOR2xp5_ASAP7_75t_L g134 ( 
.A(n_111),
.B(n_122),
.Y(n_134)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_90),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_L g136 ( 
.A(n_114),
.B(n_126),
.Y(n_136)
);

AOI22xp5_ASAP7_75t_L g145 ( 
.A1(n_115),
.A2(n_118),
.B1(n_128),
.B2(n_102),
.Y(n_145)
);

AOI21xp5_ASAP7_75t_L g117 ( 
.A1(n_82),
.A2(n_76),
.B(n_80),
.Y(n_117)
);

OAI22xp5_ASAP7_75t_L g118 ( 
.A1(n_87),
.A2(n_81),
.B1(n_15),
.B2(n_65),
.Y(n_118)
);

OA21x2_ASAP7_75t_L g120 ( 
.A1(n_93),
.A2(n_80),
.B(n_65),
.Y(n_120)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_120),
.Y(n_132)
);

CKINVDCx20_ASAP7_75t_R g121 ( 
.A(n_91),
.Y(n_121)
);

CKINVDCx20_ASAP7_75t_R g143 ( 
.A(n_121),
.Y(n_143)
);

MAJIxp5_ASAP7_75t_L g123 ( 
.A(n_94),
.B(n_73),
.C(n_8),
.Y(n_123)
);

MAJIxp5_ASAP7_75t_L g142 ( 
.A(n_123),
.B(n_98),
.C(n_8),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_L g133 ( 
.A(n_124),
.B(n_127),
.Y(n_133)
);

OAI22xp5_ASAP7_75t_SL g135 ( 
.A1(n_125),
.A2(n_103),
.B1(n_92),
.B2(n_105),
.Y(n_135)
);

AOI22xp5_ASAP7_75t_SL g126 ( 
.A1(n_104),
.A2(n_8),
.B1(n_7),
.B2(n_3),
.Y(n_126)
);

OAI21xp5_ASAP7_75t_L g127 ( 
.A1(n_95),
.A2(n_1),
.B(n_2),
.Y(n_127)
);

AOI22x1_ASAP7_75t_L g128 ( 
.A1(n_101),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_128)
);

INVx13_ASAP7_75t_L g129 ( 
.A(n_113),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_L g152 ( 
.A(n_129),
.B(n_130),
.Y(n_152)
);

CKINVDCx20_ASAP7_75t_R g130 ( 
.A(n_112),
.Y(n_130)
);

AOI22xp5_ASAP7_75t_L g149 ( 
.A1(n_135),
.A2(n_145),
.B1(n_119),
.B2(n_125),
.Y(n_149)
);

A2O1A1O1Ixp25_ASAP7_75t_L g137 ( 
.A1(n_107),
.A2(n_106),
.B(n_109),
.C(n_124),
.D(n_111),
.Y(n_137)
);

XNOR2xp5_ASAP7_75t_SL g148 ( 
.A(n_137),
.B(n_122),
.Y(n_148)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_112),
.Y(n_138)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_138),
.Y(n_157)
);

BUFx2_ASAP7_75t_L g140 ( 
.A(n_128),
.Y(n_140)
);

INVxp67_ASAP7_75t_SL g158 ( 
.A(n_140),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_L g141 ( 
.A(n_116),
.B(n_95),
.Y(n_141)
);

INVxp67_ASAP7_75t_L g150 ( 
.A(n_141),
.Y(n_150)
);

XNOR2xp5_ASAP7_75t_L g155 ( 
.A(n_142),
.B(n_144),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_L g144 ( 
.A(n_116),
.B(n_1),
.Y(n_144)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_110),
.Y(n_146)
);

AOI22xp5_ASAP7_75t_SL g147 ( 
.A1(n_146),
.A2(n_120),
.B1(n_117),
.B2(n_128),
.Y(n_147)
);

XNOR2xp5_ASAP7_75t_L g162 ( 
.A(n_147),
.B(n_139),
.Y(n_162)
);

XOR2xp5_ASAP7_75t_L g161 ( 
.A(n_148),
.B(n_156),
.Y(n_161)
);

OAI22xp5_ASAP7_75t_L g163 ( 
.A1(n_149),
.A2(n_153),
.B1(n_154),
.B2(n_145),
.Y(n_163)
);

MAJIxp5_ASAP7_75t_L g151 ( 
.A(n_134),
.B(n_120),
.C(n_108),
.Y(n_151)
);

MAJIxp5_ASAP7_75t_L g164 ( 
.A(n_151),
.B(n_131),
.C(n_133),
.Y(n_164)
);

AOI22xp5_ASAP7_75t_L g153 ( 
.A1(n_135),
.A2(n_108),
.B1(n_123),
.B2(n_102),
.Y(n_153)
);

AOI22xp5_ASAP7_75t_L g154 ( 
.A1(n_146),
.A2(n_127),
.B1(n_126),
.B2(n_7),
.Y(n_154)
);

XOR2xp5_ASAP7_75t_L g156 ( 
.A(n_134),
.B(n_7),
.Y(n_156)
);

AOI22xp5_ASAP7_75t_L g159 ( 
.A1(n_157),
.A2(n_132),
.B1(n_138),
.B2(n_130),
.Y(n_159)
);

OAI22xp5_ASAP7_75t_SL g169 ( 
.A1(n_159),
.A2(n_132),
.B1(n_139),
.B2(n_150),
.Y(n_169)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_152),
.Y(n_160)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_160),
.Y(n_170)
);

XNOR2xp5_ASAP7_75t_L g176 ( 
.A(n_162),
.B(n_164),
.Y(n_176)
);

CKINVDCx14_ASAP7_75t_R g173 ( 
.A(n_163),
.Y(n_173)
);

INVx13_ASAP7_75t_L g165 ( 
.A(n_158),
.Y(n_165)
);

OAI22xp5_ASAP7_75t_L g174 ( 
.A1(n_165),
.A2(n_167),
.B1(n_168),
.B2(n_136),
.Y(n_174)
);

MAJIxp5_ASAP7_75t_L g166 ( 
.A(n_148),
.B(n_131),
.C(n_141),
.Y(n_166)
);

MAJIxp5_ASAP7_75t_L g172 ( 
.A(n_166),
.B(n_151),
.C(n_155),
.Y(n_172)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_147),
.Y(n_167)
);

NAND3xp33_ASAP7_75t_L g168 ( 
.A(n_156),
.B(n_143),
.C(n_133),
.Y(n_168)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_169),
.Y(n_178)
);

INVxp67_ASAP7_75t_SL g171 ( 
.A(n_160),
.Y(n_171)
);

NOR2xp33_ASAP7_75t_L g180 ( 
.A(n_171),
.B(n_129),
.Y(n_180)
);

MAJIxp5_ASAP7_75t_L g181 ( 
.A(n_172),
.B(n_166),
.C(n_161),
.Y(n_181)
);

XNOR2xp5_ASAP7_75t_L g183 ( 
.A(n_174),
.B(n_142),
.Y(n_183)
);

OAI22xp5_ASAP7_75t_SL g175 ( 
.A1(n_167),
.A2(n_150),
.B1(n_137),
.B2(n_140),
.Y(n_175)
);

AOI22xp5_ASAP7_75t_L g177 ( 
.A1(n_175),
.A2(n_162),
.B1(n_165),
.B2(n_159),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_SL g186 ( 
.A(n_177),
.B(n_181),
.Y(n_186)
);

OA21x2_ASAP7_75t_L g179 ( 
.A1(n_169),
.A2(n_144),
.B(n_164),
.Y(n_179)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_179),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_L g185 ( 
.A(n_180),
.B(n_183),
.Y(n_185)
);

AOI21xp5_ASAP7_75t_SL g182 ( 
.A1(n_170),
.A2(n_155),
.B(n_161),
.Y(n_182)
);

OAI21xp5_ASAP7_75t_SL g187 ( 
.A1(n_182),
.A2(n_170),
.B(n_172),
.Y(n_187)
);

MAJIxp5_ASAP7_75t_L g189 ( 
.A(n_187),
.B(n_184),
.C(n_185),
.Y(n_189)
);

OAI21xp5_ASAP7_75t_L g188 ( 
.A1(n_179),
.A2(n_173),
.B(n_176),
.Y(n_188)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_188),
.Y(n_190)
);

MAJIxp5_ASAP7_75t_L g193 ( 
.A(n_189),
.B(n_191),
.C(n_3),
.Y(n_193)
);

MAJIxp5_ASAP7_75t_L g191 ( 
.A(n_186),
.B(n_176),
.C(n_178),
.Y(n_191)
);

AOI322xp5_ASAP7_75t_L g192 ( 
.A1(n_190),
.A2(n_180),
.A3(n_175),
.B1(n_5),
.B2(n_6),
.C1(n_4),
.C2(n_3),
.Y(n_192)
);

AOI22xp33_ASAP7_75t_L g194 ( 
.A1(n_192),
.A2(n_193),
.B1(n_4),
.B2(n_5),
.Y(n_194)
);

INVxp67_ASAP7_75t_L g195 ( 
.A(n_194),
.Y(n_195)
);

MAJIxp5_ASAP7_75t_L g196 ( 
.A(n_195),
.B(n_4),
.C(n_5),
.Y(n_196)
);

XNOR2xp5_ASAP7_75t_L g197 ( 
.A(n_196),
.B(n_6),
.Y(n_197)
);


endmodule