module fake_jpeg_8474_n_314 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_314);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_314;

wire n_253;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_51;
wire n_84;
wire n_59;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_145;
wire n_18;
wire n_20;
wire n_303;
wire n_259;
wire n_90;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_208;
wire n_308;
wire n_297;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

BUFx6f_ASAP7_75t_L g16 ( 
.A(n_5),
.Y(n_16)
);

INVx2_ASAP7_75t_L g17 ( 
.A(n_7),
.Y(n_17)
);

BUFx3_ASAP7_75t_L g18 ( 
.A(n_2),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_12),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_8),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_0),
.Y(n_21)
);

BUFx12f_ASAP7_75t_L g22 ( 
.A(n_3),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_11),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_13),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_14),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_5),
.Y(n_26)
);

BUFx12f_ASAP7_75t_L g27 ( 
.A(n_9),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_3),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_11),
.Y(n_29)
);

INVx13_ASAP7_75t_L g30 ( 
.A(n_10),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_14),
.Y(n_31)
);

INVx6_ASAP7_75t_L g32 ( 
.A(n_2),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_3),
.Y(n_33)
);

INVx4_ASAP7_75t_L g34 ( 
.A(n_22),
.Y(n_34)
);

INVx11_ASAP7_75t_L g55 ( 
.A(n_34),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_22),
.Y(n_35)
);

INVx11_ASAP7_75t_L g61 ( 
.A(n_35),
.Y(n_61)
);

BUFx5_ASAP7_75t_L g36 ( 
.A(n_22),
.Y(n_36)
);

BUFx4f_ASAP7_75t_SL g60 ( 
.A(n_36),
.Y(n_60)
);

INVx5_ASAP7_75t_L g37 ( 
.A(n_30),
.Y(n_37)
);

INVx5_ASAP7_75t_L g44 ( 
.A(n_37),
.Y(n_44)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_17),
.Y(n_38)
);

NAND2xp5_ASAP7_75t_L g49 ( 
.A(n_38),
.B(n_29),
.Y(n_49)
);

BUFx5_ASAP7_75t_L g39 ( 
.A(n_22),
.Y(n_39)
);

CKINVDCx6p67_ASAP7_75t_R g67 ( 
.A(n_39),
.Y(n_67)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_22),
.Y(n_40)
);

INVx3_ASAP7_75t_L g62 ( 
.A(n_40),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_27),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_41),
.Y(n_57)
);

INVx11_ASAP7_75t_L g42 ( 
.A(n_16),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_42),
.Y(n_59)
);

INVx8_ASAP7_75t_L g43 ( 
.A(n_16),
.Y(n_43)
);

INVx8_ASAP7_75t_L g56 ( 
.A(n_43),
.Y(n_56)
);

AOI22xp33_ASAP7_75t_SL g45 ( 
.A1(n_43),
.A2(n_32),
.B1(n_17),
.B2(n_30),
.Y(n_45)
);

OAI22xp5_ASAP7_75t_L g71 ( 
.A1(n_45),
.A2(n_47),
.B1(n_53),
.B2(n_65),
.Y(n_71)
);

INVxp67_ASAP7_75t_L g46 ( 
.A(n_36),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_SL g85 ( 
.A(n_46),
.B(n_66),
.Y(n_85)
);

AOI22xp33_ASAP7_75t_SL g47 ( 
.A1(n_43),
.A2(n_32),
.B1(n_17),
.B2(n_30),
.Y(n_47)
);

A2O1A1Ixp33_ASAP7_75t_L g48 ( 
.A1(n_37),
.A2(n_32),
.B(n_28),
.C(n_31),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_48),
.B(n_52),
.Y(n_89)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_49),
.Y(n_91)
);

BUFx12f_ASAP7_75t_L g50 ( 
.A(n_36),
.Y(n_50)
);

CKINVDCx16_ASAP7_75t_R g82 ( 
.A(n_50),
.Y(n_82)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_36),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_L g76 ( 
.A(n_51),
.B(n_64),
.Y(n_76)
);

INVx13_ASAP7_75t_L g52 ( 
.A(n_39),
.Y(n_52)
);

AOI22xp33_ASAP7_75t_L g53 ( 
.A1(n_42),
.A2(n_31),
.B1(n_23),
.B2(n_28),
.Y(n_53)
);

BUFx3_ASAP7_75t_L g54 ( 
.A(n_39),
.Y(n_54)
);

INVx3_ASAP7_75t_L g86 ( 
.A(n_54),
.Y(n_86)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_42),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_58),
.B(n_27),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_34),
.B(n_23),
.Y(n_63)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_63),
.Y(n_94)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_39),
.Y(n_64)
);

AOI22xp33_ASAP7_75t_SL g65 ( 
.A1(n_43),
.A2(n_19),
.B1(n_33),
.B2(n_25),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_34),
.B(n_26),
.Y(n_66)
);

CKINVDCx20_ASAP7_75t_R g68 ( 
.A(n_42),
.Y(n_68)
);

NOR3xp33_ASAP7_75t_L g87 ( 
.A(n_68),
.B(n_37),
.C(n_21),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_L g69 ( 
.A(n_38),
.B(n_27),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_SL g92 ( 
.A(n_69),
.B(n_41),
.Y(n_92)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_55),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_70),
.B(n_72),
.Y(n_117)
);

INVx2_ASAP7_75t_L g72 ( 
.A(n_55),
.Y(n_72)
);

BUFx6f_ASAP7_75t_L g73 ( 
.A(n_61),
.Y(n_73)
);

INVx4_ASAP7_75t_L g118 ( 
.A(n_73),
.Y(n_118)
);

OAI22xp5_ASAP7_75t_L g74 ( 
.A1(n_49),
.A2(n_43),
.B1(n_38),
.B2(n_34),
.Y(n_74)
);

O2A1O1Ixp33_ASAP7_75t_L g113 ( 
.A1(n_74),
.A2(n_93),
.B(n_46),
.C(n_29),
.Y(n_113)
);

BUFx6f_ASAP7_75t_L g75 ( 
.A(n_61),
.Y(n_75)
);

CKINVDCx16_ASAP7_75t_R g111 ( 
.A(n_75),
.Y(n_111)
);

HB1xp67_ASAP7_75t_L g77 ( 
.A(n_67),
.Y(n_77)
);

INVx2_ASAP7_75t_L g121 ( 
.A(n_77),
.Y(n_121)
);

AOI22xp5_ASAP7_75t_L g78 ( 
.A1(n_58),
.A2(n_34),
.B1(n_37),
.B2(n_19),
.Y(n_78)
);

XNOR2xp5_ASAP7_75t_L g119 ( 
.A(n_78),
.B(n_88),
.Y(n_119)
);

INVx2_ASAP7_75t_L g79 ( 
.A(n_44),
.Y(n_79)
);

CKINVDCx16_ASAP7_75t_R g105 ( 
.A(n_79),
.Y(n_105)
);

INVx13_ASAP7_75t_L g80 ( 
.A(n_67),
.Y(n_80)
);

CKINVDCx14_ASAP7_75t_R g114 ( 
.A(n_80),
.Y(n_114)
);

OR2x2_ASAP7_75t_L g81 ( 
.A(n_68),
.B(n_26),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_SL g112 ( 
.A(n_81),
.B(n_84),
.Y(n_112)
);

INVxp67_ASAP7_75t_L g83 ( 
.A(n_67),
.Y(n_83)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_83),
.Y(n_98)
);

CKINVDCx20_ASAP7_75t_R g84 ( 
.A(n_69),
.Y(n_84)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_87),
.Y(n_100)
);

AOI22xp5_ASAP7_75t_L g88 ( 
.A1(n_56),
.A2(n_19),
.B1(n_25),
.B2(n_24),
.Y(n_88)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_90),
.Y(n_103)
);

AND2x2_ASAP7_75t_L g97 ( 
.A(n_92),
.B(n_52),
.Y(n_97)
);

OAI22xp5_ASAP7_75t_SL g93 ( 
.A1(n_48),
.A2(n_21),
.B1(n_33),
.B2(n_24),
.Y(n_93)
);

CKINVDCx16_ASAP7_75t_R g95 ( 
.A(n_50),
.Y(n_95)
);

AOI22xp33_ASAP7_75t_SL g106 ( 
.A1(n_95),
.A2(n_79),
.B1(n_80),
.B2(n_56),
.Y(n_106)
);

MAJIxp5_ASAP7_75t_L g96 ( 
.A(n_84),
.B(n_91),
.C(n_76),
.Y(n_96)
);

MAJIxp5_ASAP7_75t_L g127 ( 
.A(n_96),
.B(n_88),
.C(n_94),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_SL g128 ( 
.A(n_97),
.B(n_101),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_91),
.B(n_64),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g136 ( 
.A(n_99),
.B(n_107),
.Y(n_136)
);

CKINVDCx20_ASAP7_75t_R g101 ( 
.A(n_76),
.Y(n_101)
);

AOI21xp5_ASAP7_75t_L g102 ( 
.A1(n_89),
.A2(n_44),
.B(n_60),
.Y(n_102)
);

XNOR2xp5_ASAP7_75t_L g143 ( 
.A(n_102),
.B(n_108),
.Y(n_143)
);

BUFx3_ASAP7_75t_L g104 ( 
.A(n_95),
.Y(n_104)
);

INVx11_ASAP7_75t_L g123 ( 
.A(n_104),
.Y(n_123)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_106),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_L g107 ( 
.A(n_93),
.B(n_51),
.Y(n_107)
);

AOI21xp5_ASAP7_75t_SL g108 ( 
.A1(n_85),
.A2(n_67),
.B(n_27),
.Y(n_108)
);

AOI22xp33_ASAP7_75t_SL g109 ( 
.A1(n_71),
.A2(n_52),
.B1(n_62),
.B2(n_86),
.Y(n_109)
);

OAI22xp5_ASAP7_75t_SL g124 ( 
.A1(n_109),
.A2(n_115),
.B1(n_116),
.B2(n_83),
.Y(n_124)
);

CKINVDCx20_ASAP7_75t_R g110 ( 
.A(n_81),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_SL g144 ( 
.A(n_110),
.B(n_116),
.Y(n_144)
);

AOI22xp5_ASAP7_75t_L g133 ( 
.A1(n_113),
.A2(n_70),
.B1(n_72),
.B2(n_86),
.Y(n_133)
);

AOI22xp33_ASAP7_75t_SL g115 ( 
.A1(n_71),
.A2(n_62),
.B1(n_1),
.B2(n_2),
.Y(n_115)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_74),
.Y(n_116)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_78),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_SL g148 ( 
.A(n_120),
.B(n_59),
.Y(n_148)
);

AND2x2_ASAP7_75t_L g122 ( 
.A(n_94),
.B(n_0),
.Y(n_122)
);

AND2x2_ASAP7_75t_L g130 ( 
.A(n_122),
.B(n_10),
.Y(n_130)
);

AOI22xp5_ASAP7_75t_SL g156 ( 
.A1(n_124),
.A2(n_139),
.B1(n_142),
.B2(n_110),
.Y(n_156)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_117),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_L g153 ( 
.A(n_125),
.B(n_131),
.Y(n_153)
);

INVx5_ASAP7_75t_L g126 ( 
.A(n_104),
.Y(n_126)
);

AOI22xp33_ASAP7_75t_SL g157 ( 
.A1(n_126),
.A2(n_118),
.B1(n_111),
.B2(n_105),
.Y(n_157)
);

MAJIxp5_ASAP7_75t_L g170 ( 
.A(n_127),
.B(n_135),
.C(n_102),
.Y(n_170)
);

XNOR2xp5_ASAP7_75t_SL g162 ( 
.A(n_130),
.B(n_132),
.Y(n_162)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_99),
.Y(n_131)
);

AND2x2_ASAP7_75t_L g132 ( 
.A(n_119),
.B(n_0),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_L g168 ( 
.A(n_133),
.B(n_137),
.Y(n_168)
);

NOR2xp33_ASAP7_75t_L g134 ( 
.A(n_121),
.B(n_81),
.Y(n_134)
);

CKINVDCx16_ASAP7_75t_R g149 ( 
.A(n_134),
.Y(n_149)
);

MAJIxp5_ASAP7_75t_L g135 ( 
.A(n_96),
.B(n_82),
.C(n_60),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_L g137 ( 
.A(n_121),
.B(n_50),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_L g138 ( 
.A(n_103),
.B(n_50),
.Y(n_138)
);

INVxp67_ASAP7_75t_L g155 ( 
.A(n_138),
.Y(n_155)
);

XNOR2x2_ASAP7_75t_L g139 ( 
.A(n_97),
.B(n_60),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_L g140 ( 
.A(n_101),
.B(n_60),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_L g158 ( 
.A(n_140),
.B(n_141),
.Y(n_158)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_119),
.Y(n_141)
);

AND2x2_ASAP7_75t_L g142 ( 
.A(n_120),
.B(n_0),
.Y(n_142)
);

AOI22xp5_ASAP7_75t_L g145 ( 
.A1(n_113),
.A2(n_40),
.B1(n_35),
.B2(n_41),
.Y(n_145)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_145),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_L g146 ( 
.A(n_103),
.B(n_27),
.Y(n_146)
);

INVxp67_ASAP7_75t_L g171 ( 
.A(n_146),
.Y(n_171)
);

OAI22xp5_ASAP7_75t_SL g147 ( 
.A1(n_107),
.A2(n_59),
.B1(n_35),
.B2(n_40),
.Y(n_147)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_147),
.Y(n_154)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_148),
.Y(n_159)
);

INVx2_ASAP7_75t_SL g150 ( 
.A(n_126),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_L g181 ( 
.A(n_150),
.B(n_160),
.Y(n_181)
);

OR2x2_ASAP7_75t_L g151 ( 
.A(n_144),
.B(n_112),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_L g180 ( 
.A(n_151),
.B(n_163),
.Y(n_180)
);

OAI21xp5_ASAP7_75t_L g196 ( 
.A1(n_156),
.A2(n_130),
.B(n_122),
.Y(n_196)
);

AOI22xp33_ASAP7_75t_L g192 ( 
.A1(n_157),
.A2(n_167),
.B1(n_114),
.B2(n_73),
.Y(n_192)
);

CKINVDCx20_ASAP7_75t_R g160 ( 
.A(n_123),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_L g161 ( 
.A(n_136),
.B(n_112),
.Y(n_161)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_161),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_L g163 ( 
.A(n_136),
.B(n_97),
.Y(n_163)
);

INVx2_ASAP7_75t_SL g164 ( 
.A(n_123),
.Y(n_164)
);

NOR2xp33_ASAP7_75t_L g191 ( 
.A(n_164),
.B(n_75),
.Y(n_191)
);

HB1xp67_ASAP7_75t_L g165 ( 
.A(n_139),
.Y(n_165)
);

INVx2_ASAP7_75t_L g193 ( 
.A(n_165),
.Y(n_193)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_140),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_L g187 ( 
.A(n_166),
.B(n_169),
.Y(n_187)
);

AOI22xp33_ASAP7_75t_SL g167 ( 
.A1(n_129),
.A2(n_98),
.B1(n_118),
.B2(n_105),
.Y(n_167)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_147),
.Y(n_169)
);

MAJIxp5_ASAP7_75t_L g183 ( 
.A(n_170),
.B(n_172),
.C(n_173),
.Y(n_183)
);

MAJIxp5_ASAP7_75t_L g172 ( 
.A(n_141),
.B(n_98),
.C(n_100),
.Y(n_172)
);

XOR2xp5_ASAP7_75t_L g173 ( 
.A(n_135),
.B(n_108),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_L g174 ( 
.A(n_131),
.B(n_132),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_L g188 ( 
.A(n_174),
.B(n_142),
.Y(n_188)
);

INVx11_ASAP7_75t_L g175 ( 
.A(n_133),
.Y(n_175)
);

INVx2_ASAP7_75t_L g195 ( 
.A(n_175),
.Y(n_195)
);

AOI221xp5_ASAP7_75t_L g177 ( 
.A1(n_174),
.A2(n_124),
.B1(n_143),
.B2(n_100),
.C(n_132),
.Y(n_177)
);

XOR2xp5_ASAP7_75t_L g211 ( 
.A(n_177),
.B(n_149),
.Y(n_211)
);

OAI22xp5_ASAP7_75t_SL g178 ( 
.A1(n_175),
.A2(n_129),
.B1(n_145),
.B2(n_127),
.Y(n_178)
);

AOI22xp5_ASAP7_75t_L g210 ( 
.A1(n_178),
.A2(n_154),
.B1(n_166),
.B2(n_159),
.Y(n_210)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_153),
.Y(n_179)
);

NOR2xp33_ASAP7_75t_L g206 ( 
.A(n_179),
.B(n_184),
.Y(n_206)
);

XOR2xp5_ASAP7_75t_L g182 ( 
.A(n_173),
.B(n_143),
.Y(n_182)
);

MAJIxp5_ASAP7_75t_L g202 ( 
.A(n_182),
.B(n_185),
.C(n_197),
.Y(n_202)
);

CKINVDCx20_ASAP7_75t_R g184 ( 
.A(n_151),
.Y(n_184)
);

XNOR2xp5_ASAP7_75t_L g185 ( 
.A(n_170),
.B(n_128),
.Y(n_185)
);

BUFx5_ASAP7_75t_L g186 ( 
.A(n_150),
.Y(n_186)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_186),
.Y(n_207)
);

NAND2xp5_ASAP7_75t_L g212 ( 
.A(n_188),
.B(n_176),
.Y(n_212)
);

NOR2x1_ASAP7_75t_R g189 ( 
.A(n_156),
.B(n_142),
.Y(n_189)
);

AOI22xp5_ASAP7_75t_SL g225 ( 
.A1(n_189),
.A2(n_18),
.B1(n_16),
.B2(n_20),
.Y(n_225)
);

NAND2xp5_ASAP7_75t_L g190 ( 
.A(n_161),
.B(n_130),
.Y(n_190)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_190),
.Y(n_216)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_191),
.Y(n_218)
);

OAI22xp5_ASAP7_75t_L g203 ( 
.A1(n_192),
.A2(n_152),
.B1(n_150),
.B2(n_164),
.Y(n_203)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_168),
.Y(n_194)
);

NOR2xp33_ASAP7_75t_L g213 ( 
.A(n_194),
.B(n_198),
.Y(n_213)
);

XNOR2xp5_ASAP7_75t_SL g204 ( 
.A(n_196),
.B(n_162),
.Y(n_204)
);

XNOR2xp5_ASAP7_75t_L g197 ( 
.A(n_162),
.B(n_122),
.Y(n_197)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_158),
.Y(n_198)
);

CKINVDCx20_ASAP7_75t_R g199 ( 
.A(n_160),
.Y(n_199)
);

NOR2xp33_ASAP7_75t_L g215 ( 
.A(n_199),
.B(n_200),
.Y(n_215)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_158),
.Y(n_200)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_164),
.Y(n_201)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_201),
.Y(n_220)
);

OAI22xp5_ASAP7_75t_L g238 ( 
.A1(n_203),
.A2(n_210),
.B1(n_221),
.B2(n_225),
.Y(n_238)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_204),
.Y(n_229)
);

MAJIxp5_ASAP7_75t_L g205 ( 
.A(n_183),
.B(n_172),
.C(n_163),
.Y(n_205)
);

MAJIxp5_ASAP7_75t_L g227 ( 
.A(n_205),
.B(n_211),
.C(n_219),
.Y(n_227)
);

OAI22xp5_ASAP7_75t_L g208 ( 
.A1(n_195),
.A2(n_169),
.B1(n_154),
.B2(n_152),
.Y(n_208)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_208),
.Y(n_240)
);

INVx2_ASAP7_75t_L g209 ( 
.A(n_186),
.Y(n_209)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_209),
.Y(n_243)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_212),
.Y(n_231)
);

CKINVDCx20_ASAP7_75t_R g214 ( 
.A(n_181),
.Y(n_214)
);

NOR2xp33_ASAP7_75t_L g237 ( 
.A(n_214),
.B(n_223),
.Y(n_237)
);

AND2x2_ASAP7_75t_L g217 ( 
.A(n_182),
.B(n_189),
.Y(n_217)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_217),
.Y(n_233)
);

MAJIxp5_ASAP7_75t_L g219 ( 
.A(n_183),
.B(n_159),
.C(n_155),
.Y(n_219)
);

AOI21xp5_ASAP7_75t_L g221 ( 
.A1(n_187),
.A2(n_155),
.B(n_171),
.Y(n_221)
);

XNOR2xp5_ASAP7_75t_L g222 ( 
.A(n_185),
.B(n_171),
.Y(n_222)
);

MAJIxp5_ASAP7_75t_L g235 ( 
.A(n_222),
.B(n_202),
.C(n_204),
.Y(n_235)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_187),
.Y(n_223)
);

CKINVDCx20_ASAP7_75t_R g224 ( 
.A(n_180),
.Y(n_224)
);

NOR2xp33_ASAP7_75t_L g245 ( 
.A(n_224),
.B(n_1),
.Y(n_245)
);

CKINVDCx16_ASAP7_75t_R g226 ( 
.A(n_215),
.Y(n_226)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_226),
.Y(n_257)
);

CKINVDCx20_ASAP7_75t_R g228 ( 
.A(n_206),
.Y(n_228)
);

NAND2xp5_ASAP7_75t_SL g250 ( 
.A(n_228),
.B(n_242),
.Y(n_250)
);

NAND2xp5_ASAP7_75t_L g230 ( 
.A(n_212),
.B(n_176),
.Y(n_230)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_230),
.Y(n_259)
);

AOI22xp5_ASAP7_75t_L g232 ( 
.A1(n_216),
.A2(n_195),
.B1(n_178),
.B2(n_193),
.Y(n_232)
);

OAI22xp5_ASAP7_75t_SL g255 ( 
.A1(n_232),
.A2(n_239),
.B1(n_40),
.B2(n_35),
.Y(n_255)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_213),
.Y(n_234)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_234),
.Y(n_261)
);

XNOR2xp5_ASAP7_75t_L g246 ( 
.A(n_235),
.B(n_222),
.Y(n_246)
);

MAJIxp5_ASAP7_75t_L g236 ( 
.A(n_205),
.B(n_188),
.C(n_180),
.Y(n_236)
);

MAJIxp5_ASAP7_75t_L g249 ( 
.A(n_236),
.B(n_241),
.C(n_244),
.Y(n_249)
);

AOI22xp5_ASAP7_75t_L g239 ( 
.A1(n_210),
.A2(n_193),
.B1(n_196),
.B2(n_190),
.Y(n_239)
);

MAJIxp5_ASAP7_75t_L g241 ( 
.A(n_219),
.B(n_197),
.C(n_54),
.Y(n_241)
);

CKINVDCx20_ASAP7_75t_R g242 ( 
.A(n_221),
.Y(n_242)
);

MAJIxp5_ASAP7_75t_L g244 ( 
.A(n_202),
.B(n_40),
.C(n_35),
.Y(n_244)
);

NAND2xp5_ASAP7_75t_SL g262 ( 
.A(n_245),
.B(n_4),
.Y(n_262)
);

XNOR2xp5_ASAP7_75t_L g273 ( 
.A(n_246),
.B(n_247),
.Y(n_273)
);

AOI22xp5_ASAP7_75t_SL g247 ( 
.A1(n_233),
.A2(n_217),
.B1(n_220),
.B2(n_211),
.Y(n_247)
);

AOI22xp5_ASAP7_75t_L g248 ( 
.A1(n_240),
.A2(n_218),
.B1(n_209),
.B2(n_217),
.Y(n_248)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_248),
.Y(n_263)
);

XNOR2xp5_ASAP7_75t_SL g251 ( 
.A(n_239),
.B(n_225),
.Y(n_251)
);

XNOR2xp5_ASAP7_75t_SL g269 ( 
.A(n_251),
.B(n_230),
.Y(n_269)
);

AOI22xp5_ASAP7_75t_L g252 ( 
.A1(n_233),
.A2(n_207),
.B1(n_16),
.B2(n_20),
.Y(n_252)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_252),
.Y(n_268)
);

AOI22xp5_ASAP7_75t_L g253 ( 
.A1(n_237),
.A2(n_20),
.B1(n_29),
.B2(n_18),
.Y(n_253)
);

AOI22xp5_ASAP7_75t_L g272 ( 
.A1(n_253),
.A2(n_255),
.B1(n_229),
.B2(n_73),
.Y(n_272)
);

XNOR2xp5_ASAP7_75t_L g254 ( 
.A(n_244),
.B(n_41),
.Y(n_254)
);

NAND2xp5_ASAP7_75t_L g266 ( 
.A(n_254),
.B(n_260),
.Y(n_266)
);

HB1xp67_ASAP7_75t_L g256 ( 
.A(n_243),
.Y(n_256)
);

NOR2xp33_ASAP7_75t_L g265 ( 
.A(n_256),
.B(n_231),
.Y(n_265)
);

MAJIxp5_ASAP7_75t_L g258 ( 
.A(n_236),
.B(n_57),
.C(n_75),
.Y(n_258)
);

MAJIxp5_ASAP7_75t_L g271 ( 
.A(n_258),
.B(n_227),
.C(n_241),
.Y(n_271)
);

NOR2xp33_ASAP7_75t_L g260 ( 
.A(n_234),
.B(n_1),
.Y(n_260)
);

NAND2xp5_ASAP7_75t_SL g264 ( 
.A(n_262),
.B(n_4),
.Y(n_264)
);

CKINVDCx20_ASAP7_75t_R g283 ( 
.A(n_264),
.Y(n_283)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_265),
.Y(n_285)
);

AOI22xp5_ASAP7_75t_L g267 ( 
.A1(n_259),
.A2(n_231),
.B1(n_238),
.B2(n_232),
.Y(n_267)
);

AOI22xp5_ASAP7_75t_L g280 ( 
.A1(n_267),
.A2(n_269),
.B1(n_247),
.B2(n_261),
.Y(n_280)
);

NOR2xp33_ASAP7_75t_L g270 ( 
.A(n_256),
.B(n_227),
.Y(n_270)
);

OR2x2_ASAP7_75t_L g281 ( 
.A(n_270),
.B(n_258),
.Y(n_281)
);

MAJIxp5_ASAP7_75t_L g278 ( 
.A(n_271),
.B(n_274),
.C(n_275),
.Y(n_278)
);

NOR2xp33_ASAP7_75t_L g284 ( 
.A(n_272),
.B(n_249),
.Y(n_284)
);

MAJIxp5_ASAP7_75t_L g274 ( 
.A(n_249),
.B(n_235),
.C(n_57),
.Y(n_274)
);

AOI21xp5_ASAP7_75t_L g275 ( 
.A1(n_250),
.A2(n_4),
.B(n_5),
.Y(n_275)
);

FAx1_ASAP7_75t_SL g276 ( 
.A(n_251),
.B(n_18),
.CI(n_29),
.CON(n_276),
.SN(n_276)
);

NOR2xp33_ASAP7_75t_L g279 ( 
.A(n_276),
.B(n_266),
.Y(n_279)
);

AND2x2_ASAP7_75t_L g277 ( 
.A(n_273),
.B(n_263),
.Y(n_277)
);

AOI21xp5_ASAP7_75t_L g289 ( 
.A1(n_277),
.A2(n_286),
.B(n_287),
.Y(n_289)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_279),
.Y(n_297)
);

CKINVDCx14_ASAP7_75t_R g293 ( 
.A(n_280),
.Y(n_293)
);

NAND2xp5_ASAP7_75t_SL g294 ( 
.A(n_281),
.B(n_282),
.Y(n_294)
);

NAND2xp5_ASAP7_75t_L g282 ( 
.A(n_267),
.B(n_257),
.Y(n_282)
);

AOI322xp5_ASAP7_75t_L g290 ( 
.A1(n_284),
.A2(n_271),
.A3(n_273),
.B1(n_269),
.B2(n_59),
.C1(n_10),
.C2(n_11),
.Y(n_290)
);

NAND2xp5_ASAP7_75t_L g286 ( 
.A(n_268),
.B(n_57),
.Y(n_286)
);

NOR2xp33_ASAP7_75t_L g287 ( 
.A(n_276),
.B(n_6),
.Y(n_287)
);

MAJIxp5_ASAP7_75t_L g288 ( 
.A(n_274),
.B(n_41),
.C(n_20),
.Y(n_288)
);

MAJIxp5_ASAP7_75t_L g296 ( 
.A(n_288),
.B(n_6),
.C(n_7),
.Y(n_296)
);

AOI31xp67_ASAP7_75t_L g301 ( 
.A1(n_290),
.A2(n_12),
.A3(n_13),
.B(n_14),
.Y(n_301)
);

AOI22xp5_ASAP7_75t_L g291 ( 
.A1(n_285),
.A2(n_277),
.B1(n_279),
.B2(n_287),
.Y(n_291)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_291),
.Y(n_298)
);

NOR2xp33_ASAP7_75t_L g292 ( 
.A(n_283),
.B(n_278),
.Y(n_292)
);

NOR2xp33_ASAP7_75t_SL g303 ( 
.A(n_292),
.B(n_295),
.Y(n_303)
);

NOR2xp33_ASAP7_75t_L g295 ( 
.A(n_281),
.B(n_6),
.Y(n_295)
);

NOR2xp33_ASAP7_75t_L g302 ( 
.A(n_296),
.B(n_13),
.Y(n_302)
);

NAND4xp25_ASAP7_75t_L g299 ( 
.A(n_291),
.B(n_7),
.C(n_8),
.D(n_9),
.Y(n_299)
);

AND2x2_ASAP7_75t_L g307 ( 
.A(n_299),
.B(n_15),
.Y(n_307)
);

AOI22xp5_ASAP7_75t_SL g300 ( 
.A1(n_297),
.A2(n_8),
.B1(n_9),
.B2(n_12),
.Y(n_300)
);

NAND2xp5_ASAP7_75t_SL g306 ( 
.A(n_300),
.B(n_301),
.Y(n_306)
);

NAND2xp5_ASAP7_75t_SL g308 ( 
.A(n_302),
.B(n_303),
.Y(n_308)
);

NOR2xp33_ASAP7_75t_L g304 ( 
.A(n_289),
.B(n_15),
.Y(n_304)
);

AOI21xp5_ASAP7_75t_L g305 ( 
.A1(n_304),
.A2(n_296),
.B(n_294),
.Y(n_305)
);

NAND2xp5_ASAP7_75t_L g311 ( 
.A(n_305),
.B(n_307),
.Y(n_311)
);

BUFx24_ASAP7_75t_SL g310 ( 
.A(n_308),
.Y(n_310)
);

INVxp33_ASAP7_75t_L g309 ( 
.A(n_304),
.Y(n_309)
);

OAI21xp5_ASAP7_75t_SL g312 ( 
.A1(n_311),
.A2(n_298),
.B(n_306),
.Y(n_312)
);

OAI21xp5_ASAP7_75t_SL g313 ( 
.A1(n_312),
.A2(n_293),
.B(n_309),
.Y(n_313)
);

XNOR2xp5_ASAP7_75t_L g314 ( 
.A(n_313),
.B(n_310),
.Y(n_314)
);


endmodule