module fake_jpeg_23200_n_305 (n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_305);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_305;

wire n_159;
wire n_117;
wire n_253;
wire n_286;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_14;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_251;
wire n_252;
wire n_273;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_279;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_16;
wire n_76;
wire n_127;
wire n_154;
wire n_278;
wire n_205;
wire n_295;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_293;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_281;
wire n_31;
wire n_155;
wire n_207;
wire n_277;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_291;
wire n_236;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_13;
wire n_175;
wire n_187;
wire n_57;
wire n_223;
wire n_21;
wire n_234;
wire n_288;
wire n_272;
wire n_284;
wire n_280;
wire n_171;
wire n_263;
wire n_119;
wire n_23;
wire n_301;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_289;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_267;
wire n_248;
wire n_30;
wire n_296;
wire n_168;
wire n_298;
wire n_106;
wire n_111;
wire n_197;
wire n_274;
wire n_186;
wire n_44;
wire n_24;
wire n_276;
wire n_143;
wire n_202;
wire n_25;
wire n_17;
wire n_269;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_287;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_303;
wire n_90;
wire n_304;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_266;
wire n_34;
wire n_283;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_285;
wire n_215;
wire n_262;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_294;
wire n_300;
wire n_211;
wire n_299;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_249;
wire n_302;
wire n_67;
wire n_271;
wire n_216;
wire n_217;
wire n_264;
wire n_184;
wire n_53;
wire n_268;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_297;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_265;
wire n_176;
wire n_199;
wire n_112;
wire n_260;
wire n_270;
wire n_222;
wire n_95;
wire n_275;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_290;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_292;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_140;
wire n_82;
wire n_128;
wire n_118;
wire n_258;
wire n_282;
wire n_96;

BUFx12_ASAP7_75t_L g13 ( 
.A(n_12),
.Y(n_13)
);

INVx11_ASAP7_75t_L g14 ( 
.A(n_8),
.Y(n_14)
);

INVx1_ASAP7_75t_L g15 ( 
.A(n_7),
.Y(n_15)
);

INVx4_ASAP7_75t_L g16 ( 
.A(n_5),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_6),
.Y(n_17)
);

INVx2_ASAP7_75t_L g18 ( 
.A(n_12),
.Y(n_18)
);

NOR2xp33_ASAP7_75t_SL g19 ( 
.A(n_12),
.B(n_4),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_4),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_0),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_3),
.Y(n_22)
);

INVx2_ASAP7_75t_L g23 ( 
.A(n_2),
.Y(n_23)
);

INVx2_ASAP7_75t_L g24 ( 
.A(n_6),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_7),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_6),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_10),
.Y(n_27)
);

INVx2_ASAP7_75t_L g28 ( 
.A(n_13),
.Y(n_28)
);

INVx6_ASAP7_75t_L g52 ( 
.A(n_28),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_27),
.Y(n_29)
);

INVx8_ASAP7_75t_L g40 ( 
.A(n_29),
.Y(n_40)
);

AND2x2_ASAP7_75t_L g30 ( 
.A(n_20),
.B(n_0),
.Y(n_30)
);

AND2x2_ASAP7_75t_L g47 ( 
.A(n_30),
.B(n_0),
.Y(n_47)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_25),
.Y(n_31)
);

NOR2xp33_ASAP7_75t_L g38 ( 
.A(n_31),
.B(n_35),
.Y(n_38)
);

INVx6_ASAP7_75t_L g32 ( 
.A(n_27),
.Y(n_32)
);

INVx5_ASAP7_75t_L g46 ( 
.A(n_32),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_27),
.Y(n_33)
);

INVx6_ASAP7_75t_L g53 ( 
.A(n_33),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_27),
.Y(n_34)
);

INVx3_ASAP7_75t_L g42 ( 
.A(n_34),
.Y(n_42)
);

INVx2_ASAP7_75t_SL g35 ( 
.A(n_26),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_25),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g44 ( 
.A(n_36),
.B(n_37),
.Y(n_44)
);

INVx4_ASAP7_75t_SL g37 ( 
.A(n_26),
.Y(n_37)
);

INVx2_ASAP7_75t_L g39 ( 
.A(n_29),
.Y(n_39)
);

HB1xp67_ASAP7_75t_L g58 ( 
.A(n_39),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_L g41 ( 
.A(n_30),
.B(n_15),
.Y(n_41)
);

NAND2xp5_ASAP7_75t_L g69 ( 
.A(n_41),
.B(n_45),
.Y(n_69)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_31),
.Y(n_43)
);

CKINVDCx20_ASAP7_75t_R g57 ( 
.A(n_43),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_L g45 ( 
.A(n_30),
.B(n_15),
.Y(n_45)
);

NAND2xp5_ASAP7_75t_L g71 ( 
.A(n_47),
.B(n_30),
.Y(n_71)
);

INVx2_ASAP7_75t_L g48 ( 
.A(n_29),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_48),
.B(n_49),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_SL g49 ( 
.A(n_31),
.B(n_19),
.Y(n_49)
);

INVx2_ASAP7_75t_L g50 ( 
.A(n_29),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_50),
.B(n_51),
.Y(n_63)
);

INVx2_ASAP7_75t_L g51 ( 
.A(n_29),
.Y(n_51)
);

INVx3_ASAP7_75t_L g54 ( 
.A(n_33),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_54),
.B(n_32),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_L g55 ( 
.A(n_41),
.B(n_30),
.Y(n_55)
);

XNOR2xp5_ASAP7_75t_L g89 ( 
.A(n_55),
.B(n_61),
.Y(n_89)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_38),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_59),
.B(n_66),
.Y(n_76)
);

INVx4_ASAP7_75t_L g60 ( 
.A(n_46),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_60),
.B(n_68),
.Y(n_88)
);

OAI21xp5_ASAP7_75t_L g61 ( 
.A1(n_45),
.A2(n_30),
.B(n_15),
.Y(n_61)
);

AOI22xp33_ASAP7_75t_SL g62 ( 
.A1(n_46),
.A2(n_14),
.B1(n_16),
.B2(n_18),
.Y(n_62)
);

AOI22xp33_ASAP7_75t_SL g80 ( 
.A1(n_62),
.A2(n_32),
.B1(n_37),
.B2(n_35),
.Y(n_80)
);

AOI22xp5_ASAP7_75t_L g64 ( 
.A1(n_46),
.A2(n_32),
.B1(n_37),
.B2(n_35),
.Y(n_64)
);

OAI22xp5_ASAP7_75t_SL g91 ( 
.A1(n_64),
.A2(n_53),
.B1(n_54),
.B2(n_42),
.Y(n_91)
);

CKINVDCx12_ASAP7_75t_R g65 ( 
.A(n_43),
.Y(n_65)
);

CKINVDCx16_ASAP7_75t_R g86 ( 
.A(n_65),
.Y(n_86)
);

CKINVDCx20_ASAP7_75t_R g66 ( 
.A(n_38),
.Y(n_66)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_67),
.Y(n_78)
);

BUFx16f_ASAP7_75t_L g68 ( 
.A(n_52),
.Y(n_68)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_44),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_70),
.B(n_74),
.Y(n_95)
);

AND2x2_ASAP7_75t_SL g94 ( 
.A(n_71),
.B(n_72),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_L g72 ( 
.A(n_47),
.B(n_44),
.Y(n_72)
);

BUFx12f_ASAP7_75t_L g73 ( 
.A(n_52),
.Y(n_73)
);

INVx13_ASAP7_75t_L g90 ( 
.A(n_73),
.Y(n_90)
);

INVx13_ASAP7_75t_L g74 ( 
.A(n_52),
.Y(n_74)
);

INVx2_ASAP7_75t_SL g75 ( 
.A(n_42),
.Y(n_75)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_75),
.Y(n_85)
);

NAND2x1_ASAP7_75t_SL g77 ( 
.A(n_66),
.B(n_47),
.Y(n_77)
);

A2O1A1Ixp33_ASAP7_75t_L g106 ( 
.A1(n_77),
.A2(n_71),
.B(n_72),
.C(n_55),
.Y(n_106)
);

INVx2_ASAP7_75t_L g79 ( 
.A(n_68),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_79),
.B(n_84),
.Y(n_98)
);

INVxp67_ASAP7_75t_L g109 ( 
.A(n_80),
.Y(n_109)
);

CKINVDCx20_ASAP7_75t_R g81 ( 
.A(n_57),
.Y(n_81)
);

CKINVDCx20_ASAP7_75t_R g110 ( 
.A(n_81),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_SL g82 ( 
.A(n_57),
.B(n_49),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_SL g113 ( 
.A(n_82),
.B(n_61),
.Y(n_113)
);

HB1xp67_ASAP7_75t_L g83 ( 
.A(n_73),
.Y(n_83)
);

INVx3_ASAP7_75t_SL g107 ( 
.A(n_83),
.Y(n_107)
);

INVx2_ASAP7_75t_L g84 ( 
.A(n_68),
.Y(n_84)
);

INVx6_ASAP7_75t_L g87 ( 
.A(n_73),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g115 ( 
.A(n_87),
.B(n_92),
.Y(n_115)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_91),
.Y(n_111)
);

INVx2_ASAP7_75t_L g92 ( 
.A(n_68),
.Y(n_92)
);

INVx3_ASAP7_75t_L g93 ( 
.A(n_73),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g118 ( 
.A(n_93),
.B(n_96),
.Y(n_118)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_63),
.Y(n_96)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_63),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g103 ( 
.A(n_97),
.B(n_56),
.Y(n_103)
);

INVx2_ASAP7_75t_L g99 ( 
.A(n_79),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g139 ( 
.A(n_99),
.B(n_104),
.Y(n_139)
);

INVx13_ASAP7_75t_L g100 ( 
.A(n_84),
.Y(n_100)
);

INVx4_ASAP7_75t_L g131 ( 
.A(n_100),
.Y(n_131)
);

MAJIxp5_ASAP7_75t_L g101 ( 
.A(n_94),
.B(n_69),
.C(n_55),
.Y(n_101)
);

MAJIxp5_ASAP7_75t_L g130 ( 
.A(n_101),
.B(n_114),
.C(n_77),
.Y(n_130)
);

OR2x2_ASAP7_75t_L g102 ( 
.A(n_76),
.B(n_56),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_L g120 ( 
.A(n_102),
.B(n_117),
.Y(n_120)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_103),
.Y(n_122)
);

INVx13_ASAP7_75t_L g104 ( 
.A(n_92),
.Y(n_104)
);

INVx4_ASAP7_75t_L g105 ( 
.A(n_90),
.Y(n_105)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_105),
.Y(n_123)
);

OAI21xp5_ASAP7_75t_SL g143 ( 
.A1(n_106),
.A2(n_114),
.B(n_113),
.Y(n_143)
);

OAI22xp5_ASAP7_75t_SL g108 ( 
.A1(n_76),
.A2(n_64),
.B1(n_69),
.B2(n_62),
.Y(n_108)
);

AOI22xp5_ASAP7_75t_L g133 ( 
.A1(n_108),
.A2(n_91),
.B1(n_77),
.B2(n_78),
.Y(n_133)
);

INVx2_ASAP7_75t_L g112 ( 
.A(n_93),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_L g121 ( 
.A(n_112),
.B(n_116),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_SL g126 ( 
.A(n_113),
.B(n_119),
.Y(n_126)
);

MAJIxp5_ASAP7_75t_L g114 ( 
.A(n_94),
.B(n_61),
.C(n_70),
.Y(n_114)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_95),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_L g117 ( 
.A(n_89),
.B(n_59),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_SL g119 ( 
.A(n_82),
.B(n_65),
.Y(n_119)
);

XNOR2xp5_ASAP7_75t_L g124 ( 
.A(n_117),
.B(n_89),
.Y(n_124)
);

XNOR2xp5_ASAP7_75t_L g156 ( 
.A(n_124),
.B(n_67),
.Y(n_156)
);

CKINVDCx16_ASAP7_75t_R g125 ( 
.A(n_98),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_L g144 ( 
.A(n_125),
.B(n_134),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_SL g127 ( 
.A(n_103),
.B(n_81),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_L g155 ( 
.A(n_127),
.B(n_129),
.Y(n_155)
);

CKINVDCx20_ASAP7_75t_R g128 ( 
.A(n_110),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_SL g148 ( 
.A(n_128),
.B(n_132),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_L g129 ( 
.A(n_102),
.B(n_94),
.Y(n_129)
);

MAJIxp5_ASAP7_75t_L g152 ( 
.A(n_130),
.B(n_140),
.C(n_108),
.Y(n_152)
);

CKINVDCx20_ASAP7_75t_R g132 ( 
.A(n_110),
.Y(n_132)
);

OAI22xp5_ASAP7_75t_L g145 ( 
.A1(n_133),
.A2(n_138),
.B1(n_37),
.B2(n_109),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_L g134 ( 
.A(n_116),
.B(n_97),
.Y(n_134)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_118),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_L g151 ( 
.A(n_135),
.B(n_142),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_L g136 ( 
.A(n_102),
.B(n_96),
.Y(n_136)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_136),
.Y(n_162)
);

OAI22xp5_ASAP7_75t_SL g137 ( 
.A1(n_111),
.A2(n_78),
.B1(n_64),
.B2(n_60),
.Y(n_137)
);

AOI22xp5_ASAP7_75t_L g154 ( 
.A1(n_137),
.A2(n_122),
.B1(n_37),
.B2(n_138),
.Y(n_154)
);

AOI22xp5_ASAP7_75t_L g138 ( 
.A1(n_111),
.A2(n_60),
.B1(n_32),
.B2(n_74),
.Y(n_138)
);

MAJIxp5_ASAP7_75t_L g140 ( 
.A(n_101),
.B(n_86),
.C(n_88),
.Y(n_140)
);

HB1xp67_ASAP7_75t_L g141 ( 
.A(n_100),
.Y(n_141)
);

INVx1_ASAP7_75t_SL g158 ( 
.A(n_141),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_L g142 ( 
.A(n_101),
.B(n_47),
.Y(n_142)
);

MAJIxp5_ASAP7_75t_SL g149 ( 
.A(n_143),
.B(n_114),
.C(n_108),
.Y(n_149)
);

AOI22xp5_ASAP7_75t_L g172 ( 
.A1(n_145),
.A2(n_168),
.B1(n_107),
.B2(n_85),
.Y(n_172)
);

AOI21xp5_ASAP7_75t_L g146 ( 
.A1(n_129),
.A2(n_118),
.B(n_106),
.Y(n_146)
);

AOI21xp5_ASAP7_75t_L g188 ( 
.A1(n_146),
.A2(n_147),
.B(n_150),
.Y(n_188)
);

AOI21xp5_ASAP7_75t_SL g147 ( 
.A1(n_143),
.A2(n_106),
.B(n_119),
.Y(n_147)
);

XOR2xp5_ASAP7_75t_L g173 ( 
.A(n_149),
.B(n_156),
.Y(n_173)
);

AOI21xp5_ASAP7_75t_L g150 ( 
.A1(n_136),
.A2(n_115),
.B(n_98),
.Y(n_150)
);

MAJIxp5_ASAP7_75t_L g177 ( 
.A(n_152),
.B(n_140),
.C(n_142),
.Y(n_177)
);

INVx2_ASAP7_75t_L g153 ( 
.A(n_131),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_L g170 ( 
.A(n_153),
.B(n_169),
.Y(n_170)
);

OAI22xp5_ASAP7_75t_SL g176 ( 
.A1(n_154),
.A2(n_165),
.B1(n_53),
.B2(n_40),
.Y(n_176)
);

CKINVDCx16_ASAP7_75t_R g157 ( 
.A(n_139),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_SL g182 ( 
.A(n_157),
.B(n_121),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_L g159 ( 
.A(n_127),
.B(n_86),
.Y(n_159)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_159),
.Y(n_181)
);

BUFx12f_ASAP7_75t_L g160 ( 
.A(n_131),
.Y(n_160)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_160),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_L g161 ( 
.A(n_128),
.B(n_115),
.Y(n_161)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_161),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_SL g163 ( 
.A(n_132),
.B(n_112),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_L g192 ( 
.A(n_163),
.B(n_104),
.Y(n_192)
);

NOR2xp33_ASAP7_75t_L g164 ( 
.A(n_123),
.B(n_105),
.Y(n_164)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_164),
.Y(n_194)
);

AOI22xp5_ASAP7_75t_L g165 ( 
.A1(n_137),
.A2(n_107),
.B1(n_74),
.B2(n_105),
.Y(n_165)
);

XNOR2xp5_ASAP7_75t_L g166 ( 
.A(n_130),
.B(n_73),
.Y(n_166)
);

XOR2xp5_ASAP7_75t_L g175 ( 
.A(n_166),
.B(n_152),
.Y(n_175)
);

AOI22xp5_ASAP7_75t_SL g167 ( 
.A1(n_122),
.A2(n_120),
.B1(n_133),
.B2(n_135),
.Y(n_167)
);

OAI22xp5_ASAP7_75t_SL g193 ( 
.A1(n_167),
.A2(n_90),
.B1(n_28),
.B2(n_18),
.Y(n_193)
);

OAI22xp5_ASAP7_75t_L g168 ( 
.A1(n_125),
.A2(n_85),
.B1(n_18),
.B2(n_87),
.Y(n_168)
);

INVx2_ASAP7_75t_L g169 ( 
.A(n_123),
.Y(n_169)
);

AO22x2_ASAP7_75t_L g171 ( 
.A1(n_149),
.A2(n_167),
.B1(n_162),
.B2(n_154),
.Y(n_171)
);

AOI22x1_ASAP7_75t_L g202 ( 
.A1(n_171),
.A2(n_160),
.B1(n_58),
.B2(n_26),
.Y(n_202)
);

OAI22xp5_ASAP7_75t_L g199 ( 
.A1(n_172),
.A2(n_171),
.B1(n_194),
.B2(n_191),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_L g174 ( 
.A(n_155),
.B(n_120),
.Y(n_174)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_174),
.Y(n_207)
);

MAJIxp5_ASAP7_75t_L g196 ( 
.A(n_175),
.B(n_177),
.C(n_179),
.Y(n_196)
);

AOI22xp5_ASAP7_75t_L g205 ( 
.A1(n_176),
.A2(n_178),
.B1(n_193),
.B2(n_90),
.Y(n_205)
);

OAI22xp5_ASAP7_75t_SL g178 ( 
.A1(n_155),
.A2(n_134),
.B1(n_121),
.B2(n_126),
.Y(n_178)
);

XOR2xp5_ASAP7_75t_L g179 ( 
.A(n_166),
.B(n_124),
.Y(n_179)
);

AND2x2_ASAP7_75t_L g180 ( 
.A(n_144),
.B(n_126),
.Y(n_180)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_180),
.Y(n_215)
);

NAND2xp5_ASAP7_75t_L g206 ( 
.A(n_182),
.B(n_185),
.Y(n_206)
);

NAND3xp33_ASAP7_75t_L g184 ( 
.A(n_151),
.B(n_11),
.C(n_10),
.Y(n_184)
);

XNOR2xp5_ASAP7_75t_L g204 ( 
.A(n_184),
.B(n_192),
.Y(n_204)
);

NAND2xp5_ASAP7_75t_SL g185 ( 
.A(n_148),
.B(n_99),
.Y(n_185)
);

NOR2xp33_ASAP7_75t_L g186 ( 
.A(n_158),
.B(n_107),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_L g213 ( 
.A(n_186),
.B(n_187),
.Y(n_213)
);

NAND2xp5_ASAP7_75t_SL g187 ( 
.A(n_158),
.B(n_169),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_SL g189 ( 
.A(n_153),
.B(n_107),
.Y(n_189)
);

CKINVDCx20_ASAP7_75t_R g212 ( 
.A(n_189),
.Y(n_212)
);

NOR2xp33_ASAP7_75t_L g190 ( 
.A(n_165),
.B(n_104),
.Y(n_190)
);

CKINVDCx20_ASAP7_75t_R g214 ( 
.A(n_190),
.Y(n_214)
);

BUFx4f_ASAP7_75t_SL g195 ( 
.A(n_171),
.Y(n_195)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_195),
.Y(n_226)
);

MAJIxp5_ASAP7_75t_L g197 ( 
.A(n_175),
.B(n_146),
.C(n_150),
.Y(n_197)
);

MAJIxp5_ASAP7_75t_L g219 ( 
.A(n_197),
.B(n_203),
.C(n_181),
.Y(n_219)
);

XNOR2xp5_ASAP7_75t_L g198 ( 
.A(n_173),
.B(n_156),
.Y(n_198)
);

XOR2xp5_ASAP7_75t_L g216 ( 
.A(n_198),
.B(n_174),
.Y(n_216)
);

AOI22xp5_ASAP7_75t_L g225 ( 
.A1(n_199),
.A2(n_53),
.B1(n_40),
.B2(n_24),
.Y(n_225)
);

AND2x2_ASAP7_75t_L g200 ( 
.A(n_171),
.B(n_147),
.Y(n_200)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_200),
.Y(n_235)
);

MAJx2_ASAP7_75t_L g201 ( 
.A(n_173),
.B(n_160),
.C(n_58),
.Y(n_201)
);

XNOR2xp5_ASAP7_75t_SL g232 ( 
.A(n_201),
.B(n_26),
.Y(n_232)
);

OAI22xp5_ASAP7_75t_SL g227 ( 
.A1(n_202),
.A2(n_205),
.B1(n_208),
.B2(n_211),
.Y(n_227)
);

MAJIxp5_ASAP7_75t_L g203 ( 
.A(n_177),
.B(n_179),
.C(n_188),
.Y(n_203)
);

AOI22xp5_ASAP7_75t_L g208 ( 
.A1(n_176),
.A2(n_100),
.B1(n_16),
.B2(n_23),
.Y(n_208)
);

XNOR2x1_ASAP7_75t_L g209 ( 
.A(n_188),
.B(n_24),
.Y(n_209)
);

XNOR2x1_ASAP7_75t_L g223 ( 
.A(n_209),
.B(n_23),
.Y(n_223)
);

XNOR2xp5_ASAP7_75t_L g210 ( 
.A(n_193),
.B(n_28),
.Y(n_210)
);

XNOR2xp5_ASAP7_75t_L g218 ( 
.A(n_210),
.B(n_172),
.Y(n_218)
);

AOI22xp5_ASAP7_75t_L g211 ( 
.A1(n_178),
.A2(n_16),
.B1(n_23),
.B2(n_24),
.Y(n_211)
);

XOR2xp5_ASAP7_75t_L g236 ( 
.A(n_216),
.B(n_217),
.Y(n_236)
);

XOR2xp5_ASAP7_75t_L g217 ( 
.A(n_196),
.B(n_180),
.Y(n_217)
);

XNOR2xp5_ASAP7_75t_L g244 ( 
.A(n_218),
.B(n_222),
.Y(n_244)
);

MAJIxp5_ASAP7_75t_L g241 ( 
.A(n_219),
.B(n_221),
.C(n_216),
.Y(n_241)
);

OAI21xp5_ASAP7_75t_L g220 ( 
.A1(n_195),
.A2(n_170),
.B(n_183),
.Y(n_220)
);

AOI21xp5_ASAP7_75t_L g242 ( 
.A1(n_220),
.A2(n_201),
.B(n_198),
.Y(n_242)
);

MAJIxp5_ASAP7_75t_L g221 ( 
.A(n_196),
.B(n_180),
.C(n_40),
.Y(n_221)
);

XNOR2xp5_ASAP7_75t_L g222 ( 
.A(n_197),
.B(n_28),
.Y(n_222)
);

AO21x1_ASAP7_75t_L g252 ( 
.A1(n_223),
.A2(n_228),
.B(n_75),
.Y(n_252)
);

NAND2xp5_ASAP7_75t_SL g224 ( 
.A(n_206),
.B(n_214),
.Y(n_224)
);

NAND2xp5_ASAP7_75t_L g239 ( 
.A(n_224),
.B(n_229),
.Y(n_239)
);

OAI22xp5_ASAP7_75t_SL g245 ( 
.A1(n_225),
.A2(n_48),
.B1(n_39),
.B2(n_17),
.Y(n_245)
);

A2O1A1Ixp33_ASAP7_75t_SL g228 ( 
.A1(n_195),
.A2(n_75),
.B(n_51),
.C(n_50),
.Y(n_228)
);

CKINVDCx20_ASAP7_75t_R g229 ( 
.A(n_213),
.Y(n_229)
);

OAI22xp5_ASAP7_75t_SL g230 ( 
.A1(n_215),
.A2(n_14),
.B1(n_36),
.B2(n_17),
.Y(n_230)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_230),
.Y(n_238)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_202),
.Y(n_231)
);

NAND2xp5_ASAP7_75t_L g240 ( 
.A(n_231),
.B(n_204),
.Y(n_240)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_232),
.Y(n_248)
);

OAI22xp5_ASAP7_75t_SL g233 ( 
.A1(n_209),
.A2(n_14),
.B1(n_36),
.B2(n_17),
.Y(n_233)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_233),
.Y(n_250)
);

OAI22xp5_ASAP7_75t_SL g234 ( 
.A1(n_200),
.A2(n_207),
.B1(n_212),
.B2(n_203),
.Y(n_234)
);

NAND2xp5_ASAP7_75t_SL g246 ( 
.A(n_234),
.B(n_9),
.Y(n_246)
);

HB1xp67_ASAP7_75t_L g237 ( 
.A(n_228),
.Y(n_237)
);

CKINVDCx14_ASAP7_75t_R g265 ( 
.A(n_237),
.Y(n_265)
);

NAND2xp5_ASAP7_75t_L g266 ( 
.A(n_240),
.B(n_246),
.Y(n_266)
);

MAJIxp5_ASAP7_75t_L g263 ( 
.A(n_241),
.B(n_243),
.C(n_251),
.Y(n_263)
);

AOI21xp5_ASAP7_75t_L g264 ( 
.A1(n_242),
.A2(n_252),
.B(n_22),
.Y(n_264)
);

A2O1A1O1Ixp25_ASAP7_75t_L g243 ( 
.A1(n_235),
.A2(n_19),
.B(n_11),
.C(n_10),
.D(n_9),
.Y(n_243)
);

AOI22xp5_ASAP7_75t_L g262 ( 
.A1(n_245),
.A2(n_35),
.B1(n_21),
.B2(n_22),
.Y(n_262)
);

BUFx12_ASAP7_75t_L g247 ( 
.A(n_226),
.Y(n_247)
);

NAND2xp5_ASAP7_75t_SL g259 ( 
.A(n_247),
.B(n_249),
.Y(n_259)
);

XNOR2xp5_ASAP7_75t_L g249 ( 
.A(n_232),
.B(n_13),
.Y(n_249)
);

XNOR2xp5_ASAP7_75t_L g251 ( 
.A(n_219),
.B(n_222),
.Y(n_251)
);

MAJIxp5_ASAP7_75t_L g253 ( 
.A(n_236),
.B(n_221),
.C(n_217),
.Y(n_253)
);

MAJIxp5_ASAP7_75t_L g271 ( 
.A(n_253),
.B(n_256),
.C(n_257),
.Y(n_271)
);

OAI22xp5_ASAP7_75t_L g254 ( 
.A1(n_237),
.A2(n_239),
.B1(n_250),
.B2(n_238),
.Y(n_254)
);

AOI22xp5_ASAP7_75t_L g268 ( 
.A1(n_254),
.A2(n_35),
.B1(n_21),
.B2(n_20),
.Y(n_268)
);

OAI21xp5_ASAP7_75t_SL g255 ( 
.A1(n_247),
.A2(n_228),
.B(n_227),
.Y(n_255)
);

OAI21xp5_ASAP7_75t_SL g273 ( 
.A1(n_255),
.A2(n_261),
.B(n_20),
.Y(n_273)
);

XOR2xp5_ASAP7_75t_L g256 ( 
.A(n_236),
.B(n_223),
.Y(n_256)
);

MAJIxp5_ASAP7_75t_L g257 ( 
.A(n_247),
.B(n_228),
.C(n_75),
.Y(n_257)
);

MAJIxp5_ASAP7_75t_L g258 ( 
.A(n_248),
.B(n_33),
.C(n_34),
.Y(n_258)
);

MAJIxp5_ASAP7_75t_L g275 ( 
.A(n_258),
.B(n_267),
.C(n_34),
.Y(n_275)
);

XNOR2xp5_ASAP7_75t_SL g260 ( 
.A(n_252),
.B(n_9),
.Y(n_260)
);

XOR2xp5_ASAP7_75t_L g274 ( 
.A(n_260),
.B(n_264),
.Y(n_274)
);

OAI21xp5_ASAP7_75t_SL g261 ( 
.A1(n_244),
.A2(n_22),
.B(n_21),
.Y(n_261)
);

NAND2xp5_ASAP7_75t_L g272 ( 
.A(n_262),
.B(n_0),
.Y(n_272)
);

MAJIxp5_ASAP7_75t_L g267 ( 
.A(n_243),
.B(n_34),
.C(n_33),
.Y(n_267)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_268),
.Y(n_286)
);

NAND2xp5_ASAP7_75t_SL g269 ( 
.A(n_266),
.B(n_11),
.Y(n_269)
);

NAND2xp5_ASAP7_75t_L g284 ( 
.A(n_269),
.B(n_272),
.Y(n_284)
);

HB1xp67_ASAP7_75t_L g270 ( 
.A(n_265),
.Y(n_270)
);

OA21x2_ASAP7_75t_L g288 ( 
.A1(n_270),
.A2(n_279),
.B(n_1),
.Y(n_288)
);

OAI22xp5_ASAP7_75t_SL g281 ( 
.A1(n_273),
.A2(n_263),
.B1(n_258),
.B2(n_3),
.Y(n_281)
);

AOI22xp5_ASAP7_75t_L g289 ( 
.A1(n_275),
.A2(n_35),
.B1(n_2),
.B2(n_3),
.Y(n_289)
);

OR2x2_ASAP7_75t_L g276 ( 
.A(n_267),
.B(n_34),
.Y(n_276)
);

NAND2xp5_ASAP7_75t_L g285 ( 
.A(n_276),
.B(n_278),
.Y(n_285)
);

CKINVDCx14_ASAP7_75t_R g277 ( 
.A(n_260),
.Y(n_277)
);

OAI21xp5_ASAP7_75t_L g280 ( 
.A1(n_277),
.A2(n_279),
.B(n_259),
.Y(n_280)
);

MAJIxp5_ASAP7_75t_L g278 ( 
.A(n_253),
.B(n_1),
.C(n_2),
.Y(n_278)
);

HB1xp67_ASAP7_75t_L g279 ( 
.A(n_257),
.Y(n_279)
);

NAND2xp5_ASAP7_75t_SL g294 ( 
.A(n_280),
.B(n_282),
.Y(n_294)
);

NAND2xp5_ASAP7_75t_L g295 ( 
.A(n_281),
.B(n_287),
.Y(n_295)
);

CKINVDCx16_ASAP7_75t_R g282 ( 
.A(n_270),
.Y(n_282)
);

A2O1A1Ixp33_ASAP7_75t_L g283 ( 
.A1(n_277),
.A2(n_256),
.B(n_33),
.C(n_3),
.Y(n_283)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_283),
.Y(n_290)
);

OAI21xp5_ASAP7_75t_L g287 ( 
.A1(n_271),
.A2(n_1),
.B(n_2),
.Y(n_287)
);

MAJx2_ASAP7_75t_L g293 ( 
.A(n_288),
.B(n_1),
.C(n_4),
.Y(n_293)
);

OAI22xp5_ASAP7_75t_SL g292 ( 
.A1(n_289),
.A2(n_283),
.B1(n_286),
.B2(n_285),
.Y(n_292)
);

NAND4xp25_ASAP7_75t_SL g291 ( 
.A(n_288),
.B(n_274),
.C(n_13),
.D(n_5),
.Y(n_291)
);

MAJIxp5_ASAP7_75t_L g298 ( 
.A(n_291),
.B(n_290),
.C(n_294),
.Y(n_298)
);

MAJIxp5_ASAP7_75t_L g296 ( 
.A(n_292),
.B(n_293),
.C(n_295),
.Y(n_296)
);

NAND2xp5_ASAP7_75t_L g299 ( 
.A(n_296),
.B(n_297),
.Y(n_299)
);

MAJIxp5_ASAP7_75t_L g297 ( 
.A(n_294),
.B(n_280),
.C(n_284),
.Y(n_297)
);

NAND2xp5_ASAP7_75t_L g300 ( 
.A(n_298),
.B(n_4),
.Y(n_300)
);

AOI21x1_ASAP7_75t_SL g301 ( 
.A1(n_300),
.A2(n_5),
.B(n_6),
.Y(n_301)
);

AOI322xp5_ASAP7_75t_L g302 ( 
.A1(n_301),
.A2(n_5),
.A3(n_7),
.B1(n_8),
.B2(n_13),
.C1(n_299),
.C2(n_237),
.Y(n_302)
);

INVx2_ASAP7_75t_L g303 ( 
.A(n_302),
.Y(n_303)
);

AO21x1_ASAP7_75t_L g304 ( 
.A1(n_303),
.A2(n_13),
.B(n_7),
.Y(n_304)
);

AOI21xp5_ASAP7_75t_L g305 ( 
.A1(n_304),
.A2(n_8),
.B(n_13),
.Y(n_305)
);


endmodule