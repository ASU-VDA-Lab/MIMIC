module fake_jpeg_29118_n_235 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_235);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_235;

wire n_159;
wire n_117;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_16;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_57;
wire n_21;
wire n_223;
wire n_234;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_44;
wire n_24;
wire n_143;
wire n_202;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_37;
wire n_233;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_232;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_131;
wire n_56;
wire n_212;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_216;
wire n_217;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_48;
wire n_35;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

INVx1_ASAP7_75t_L g15 ( 
.A(n_13),
.Y(n_15)
);

BUFx8_ASAP7_75t_L g16 ( 
.A(n_3),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_9),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_2),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_10),
.Y(n_19)
);

INVx4_ASAP7_75t_L g20 ( 
.A(n_5),
.Y(n_20)
);

BUFx3_ASAP7_75t_L g21 ( 
.A(n_9),
.Y(n_21)
);

BUFx2_ASAP7_75t_L g22 ( 
.A(n_10),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_4),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_0),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_11),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_11),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_13),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_4),
.Y(n_28)
);

INVx3_ASAP7_75t_L g29 ( 
.A(n_5),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_2),
.Y(n_30)
);

BUFx12f_ASAP7_75t_L g31 ( 
.A(n_4),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_10),
.Y(n_32)
);

BUFx5_ASAP7_75t_L g33 ( 
.A(n_6),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_0),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_8),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_2),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_23),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g76 ( 
.A(n_37),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g38 ( 
.A(n_26),
.B(n_14),
.Y(n_38)
);

AND2x2_ASAP7_75t_L g94 ( 
.A(n_38),
.B(n_47),
.Y(n_94)
);

INVx4_ASAP7_75t_L g39 ( 
.A(n_20),
.Y(n_39)
);

INVx4_ASAP7_75t_L g70 ( 
.A(n_39),
.Y(n_70)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_23),
.Y(n_40)
);

INVx6_ASAP7_75t_L g72 ( 
.A(n_40),
.Y(n_72)
);

INVx2_ASAP7_75t_L g41 ( 
.A(n_22),
.Y(n_41)
);

INVx2_ASAP7_75t_L g69 ( 
.A(n_41),
.Y(n_69)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_22),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_42),
.B(n_55),
.Y(n_60)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_28),
.Y(n_43)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_43),
.Y(n_68)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_28),
.Y(n_44)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_44),
.Y(n_81)
);

INVx13_ASAP7_75t_L g45 ( 
.A(n_29),
.Y(n_45)
);

BUFx12f_ASAP7_75t_L g61 ( 
.A(n_45),
.Y(n_61)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_30),
.Y(n_46)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_46),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g47 ( 
.A(n_26),
.B(n_14),
.Y(n_47)
);

INVx3_ASAP7_75t_L g48 ( 
.A(n_31),
.Y(n_48)
);

INVx3_ASAP7_75t_L g77 ( 
.A(n_48),
.Y(n_77)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_23),
.Y(n_49)
);

INVx6_ASAP7_75t_L g96 ( 
.A(n_49),
.Y(n_96)
);

INVx2_ASAP7_75t_L g50 ( 
.A(n_22),
.Y(n_50)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_50),
.Y(n_85)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_30),
.Y(n_51)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_51),
.Y(n_87)
);

BUFx12f_ASAP7_75t_L g52 ( 
.A(n_35),
.Y(n_52)
);

INVx3_ASAP7_75t_L g80 ( 
.A(n_52),
.Y(n_80)
);

INVx3_ASAP7_75t_L g53 ( 
.A(n_31),
.Y(n_53)
);

INVx3_ASAP7_75t_L g88 ( 
.A(n_53),
.Y(n_88)
);

BUFx3_ASAP7_75t_L g54 ( 
.A(n_33),
.Y(n_54)
);

INVx5_ASAP7_75t_L g90 ( 
.A(n_54),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_15),
.B(n_12),
.Y(n_55)
);

INVx6_ASAP7_75t_L g56 ( 
.A(n_35),
.Y(n_56)
);

INVx8_ASAP7_75t_L g86 ( 
.A(n_56),
.Y(n_86)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_35),
.Y(n_57)
);

BUFx3_ASAP7_75t_L g67 ( 
.A(n_57),
.Y(n_67)
);

INVx8_ASAP7_75t_L g58 ( 
.A(n_16),
.Y(n_58)
);

INVx3_ASAP7_75t_L g93 ( 
.A(n_58),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_15),
.B(n_12),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_59),
.B(n_25),
.Y(n_71)
);

INVx2_ASAP7_75t_SL g62 ( 
.A(n_48),
.Y(n_62)
);

INVx13_ASAP7_75t_L g111 ( 
.A(n_62),
.Y(n_111)
);

CKINVDCx16_ASAP7_75t_R g63 ( 
.A(n_43),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_63),
.B(n_65),
.Y(n_103)
);

NOR3xp33_ASAP7_75t_L g64 ( 
.A(n_44),
.B(n_19),
.C(n_32),
.Y(n_64)
);

NAND3xp33_ASAP7_75t_L g104 ( 
.A(n_64),
.B(n_34),
.C(n_1),
.Y(n_104)
);

CKINVDCx20_ASAP7_75t_R g65 ( 
.A(n_54),
.Y(n_65)
);

AOI22xp33_ASAP7_75t_SL g66 ( 
.A1(n_58),
.A2(n_20),
.B1(n_29),
.B2(n_21),
.Y(n_66)
);

AOI22xp33_ASAP7_75t_SL g106 ( 
.A1(n_66),
.A2(n_91),
.B1(n_95),
.B2(n_61),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g115 ( 
.A(n_71),
.B(n_73),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_46),
.B(n_25),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_L g74 ( 
.A(n_51),
.B(n_18),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_SL g124 ( 
.A(n_74),
.B(n_82),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_45),
.B(n_18),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g118 ( 
.A(n_75),
.B(n_84),
.Y(n_118)
);

OAI22xp5_ASAP7_75t_L g78 ( 
.A1(n_56),
.A2(n_27),
.B1(n_36),
.B2(n_19),
.Y(n_78)
);

AOI22xp33_ASAP7_75t_L g107 ( 
.A1(n_78),
.A2(n_52),
.B1(n_16),
.B2(n_3),
.Y(n_107)
);

OR2x2_ASAP7_75t_L g79 ( 
.A(n_42),
.B(n_32),
.Y(n_79)
);

OR2x2_ASAP7_75t_L g97 ( 
.A(n_79),
.B(n_17),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g82 ( 
.A(n_41),
.B(n_36),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_53),
.B(n_24),
.Y(n_84)
);

CKINVDCx20_ASAP7_75t_R g89 ( 
.A(n_50),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g127 ( 
.A(n_89),
.B(n_92),
.Y(n_127)
);

AOI22xp33_ASAP7_75t_SL g91 ( 
.A1(n_52),
.A2(n_21),
.B1(n_31),
.B2(n_33),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_SL g92 ( 
.A(n_39),
.B(n_24),
.Y(n_92)
);

AOI22xp33_ASAP7_75t_SL g95 ( 
.A1(n_52),
.A2(n_31),
.B1(n_27),
.B2(n_17),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g145 ( 
.A(n_97),
.B(n_102),
.Y(n_145)
);

INVx2_ASAP7_75t_L g98 ( 
.A(n_69),
.Y(n_98)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_98),
.Y(n_140)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_68),
.Y(n_99)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_99),
.Y(n_141)
);

OAI22xp5_ASAP7_75t_L g100 ( 
.A1(n_95),
.A2(n_57),
.B1(n_49),
.B2(n_40),
.Y(n_100)
);

OAI22xp5_ASAP7_75t_L g135 ( 
.A1(n_100),
.A2(n_107),
.B1(n_122),
.B2(n_72),
.Y(n_135)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_81),
.Y(n_101)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_101),
.Y(n_147)
);

CKINVDCx16_ASAP7_75t_R g102 ( 
.A(n_83),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_L g132 ( 
.A(n_104),
.B(n_116),
.Y(n_132)
);

OAI22xp33_ASAP7_75t_SL g105 ( 
.A1(n_87),
.A2(n_37),
.B1(n_27),
.B2(n_34),
.Y(n_105)
);

AOI22xp5_ASAP7_75t_SL g136 ( 
.A1(n_105),
.A2(n_106),
.B1(n_86),
.B2(n_88),
.Y(n_136)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_85),
.Y(n_108)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_108),
.Y(n_150)
);

AOI22xp33_ASAP7_75t_SL g109 ( 
.A1(n_66),
.A2(n_16),
.B1(n_1),
.B2(n_3),
.Y(n_109)
);

CKINVDCx16_ASAP7_75t_R g138 ( 
.A(n_109),
.Y(n_138)
);

INVx11_ASAP7_75t_L g110 ( 
.A(n_90),
.Y(n_110)
);

INVx3_ASAP7_75t_SL g151 ( 
.A(n_110),
.Y(n_151)
);

BUFx6f_ASAP7_75t_L g112 ( 
.A(n_76),
.Y(n_112)
);

HB1xp67_ASAP7_75t_L g131 ( 
.A(n_112),
.Y(n_131)
);

AOI22xp33_ASAP7_75t_SL g113 ( 
.A1(n_90),
.A2(n_16),
.B1(n_1),
.B2(n_5),
.Y(n_113)
);

OAI21xp5_ASAP7_75t_SL g149 ( 
.A1(n_113),
.A2(n_122),
.B(n_100),
.Y(n_149)
);

INVx8_ASAP7_75t_L g114 ( 
.A(n_80),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_L g152 ( 
.A(n_114),
.B(n_110),
.Y(n_152)
);

INVx3_ASAP7_75t_L g116 ( 
.A(n_77),
.Y(n_116)
);

OAI32xp33_ASAP7_75t_L g117 ( 
.A1(n_60),
.A2(n_0),
.A3(n_6),
.B1(n_7),
.B2(n_8),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_L g137 ( 
.A(n_117),
.B(n_121),
.Y(n_137)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_69),
.Y(n_119)
);

AND2x2_ASAP7_75t_L g144 ( 
.A(n_119),
.B(n_120),
.Y(n_144)
);

AOI22xp5_ASAP7_75t_SL g120 ( 
.A1(n_94),
.A2(n_6),
.B1(n_7),
.B2(n_8),
.Y(n_120)
);

INVx13_ASAP7_75t_L g121 ( 
.A(n_93),
.Y(n_121)
);

OAI22xp5_ASAP7_75t_L g122 ( 
.A1(n_91),
.A2(n_7),
.B1(n_9),
.B2(n_96),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_L g123 ( 
.A(n_79),
.B(n_94),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_L g139 ( 
.A(n_123),
.B(n_126),
.Y(n_139)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_77),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_SL g133 ( 
.A(n_125),
.B(n_70),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_L g126 ( 
.A(n_72),
.B(n_96),
.Y(n_126)
);

INVx3_ASAP7_75t_L g128 ( 
.A(n_88),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_L g142 ( 
.A(n_128),
.B(n_61),
.Y(n_142)
);

AND2x2_ASAP7_75t_L g129 ( 
.A(n_70),
.B(n_80),
.Y(n_129)
);

MAJIxp5_ASAP7_75t_L g134 ( 
.A(n_129),
.B(n_93),
.C(n_62),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_SL g130 ( 
.A(n_123),
.B(n_61),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_SL g158 ( 
.A(n_130),
.B(n_148),
.Y(n_158)
);

CKINVDCx16_ASAP7_75t_R g162 ( 
.A(n_133),
.Y(n_162)
);

MAJIxp5_ASAP7_75t_L g165 ( 
.A(n_134),
.B(n_129),
.C(n_125),
.Y(n_165)
);

OAI22xp5_ASAP7_75t_L g163 ( 
.A1(n_135),
.A2(n_136),
.B1(n_143),
.B2(n_126),
.Y(n_163)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_142),
.Y(n_153)
);

OAI22xp5_ASAP7_75t_L g143 ( 
.A1(n_124),
.A2(n_76),
.B1(n_86),
.B2(n_67),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_SL g146 ( 
.A(n_127),
.B(n_67),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_L g161 ( 
.A(n_146),
.B(n_120),
.Y(n_161)
);

NOR2xp33_ASAP7_75t_SL g148 ( 
.A(n_118),
.B(n_115),
.Y(n_148)
);

INVx4_ASAP7_75t_SL g170 ( 
.A(n_149),
.Y(n_170)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_152),
.Y(n_156)
);

CKINVDCx20_ASAP7_75t_R g154 ( 
.A(n_146),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_SL g181 ( 
.A(n_154),
.B(n_157),
.Y(n_181)
);

AND2x6_ASAP7_75t_L g155 ( 
.A(n_137),
.B(n_117),
.Y(n_155)
);

NOR3xp33_ASAP7_75t_SL g184 ( 
.A(n_155),
.B(n_138),
.C(n_143),
.Y(n_184)
);

CKINVDCx20_ASAP7_75t_R g157 ( 
.A(n_133),
.Y(n_157)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_141),
.Y(n_159)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_159),
.Y(n_172)
);

OAI21xp5_ASAP7_75t_SL g160 ( 
.A1(n_139),
.A2(n_103),
.B(n_99),
.Y(n_160)
);

XNOR2xp5_ASAP7_75t_L g185 ( 
.A(n_160),
.B(n_165),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_L g174 ( 
.A(n_161),
.B(n_164),
.Y(n_174)
);

OAI22xp5_ASAP7_75t_L g177 ( 
.A1(n_163),
.A2(n_154),
.B1(n_162),
.B2(n_136),
.Y(n_177)
);

NOR2xp33_ASAP7_75t_SL g164 ( 
.A(n_145),
.B(n_101),
.Y(n_164)
);

INVx13_ASAP7_75t_L g166 ( 
.A(n_151),
.Y(n_166)
);

INVx3_ASAP7_75t_L g171 ( 
.A(n_166),
.Y(n_171)
);

INVx2_ASAP7_75t_L g167 ( 
.A(n_140),
.Y(n_167)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_167),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_SL g168 ( 
.A(n_148),
.B(n_97),
.Y(n_168)
);

NOR2xp33_ASAP7_75t_L g186 ( 
.A(n_168),
.B(n_169),
.Y(n_186)
);

NOR2xp33_ASAP7_75t_L g169 ( 
.A(n_145),
.B(n_102),
.Y(n_169)
);

XOR2xp5_ASAP7_75t_L g175 ( 
.A(n_160),
.B(n_139),
.Y(n_175)
);

MAJIxp5_ASAP7_75t_L g190 ( 
.A(n_175),
.B(n_178),
.C(n_179),
.Y(n_190)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_159),
.Y(n_176)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_176),
.Y(n_187)
);

AOI22xp5_ASAP7_75t_SL g192 ( 
.A1(n_177),
.A2(n_180),
.B1(n_163),
.B2(n_135),
.Y(n_192)
);

MAJIxp5_ASAP7_75t_L g178 ( 
.A(n_165),
.B(n_134),
.C(n_130),
.Y(n_178)
);

MAJIxp5_ASAP7_75t_L g179 ( 
.A(n_156),
.B(n_144),
.C(n_141),
.Y(n_179)
);

OAI22xp5_ASAP7_75t_L g180 ( 
.A1(n_170),
.A2(n_138),
.B1(n_149),
.B2(n_144),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_L g182 ( 
.A(n_157),
.B(n_147),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_L g193 ( 
.A(n_182),
.B(n_162),
.Y(n_193)
);

AOI21xp5_ASAP7_75t_SL g183 ( 
.A1(n_170),
.A2(n_132),
.B(n_144),
.Y(n_183)
);

OAI21xp5_ASAP7_75t_SL g189 ( 
.A1(n_183),
.A2(n_181),
.B(n_174),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_SL g188 ( 
.A(n_184),
.B(n_161),
.Y(n_188)
);

OAI21xp5_ASAP7_75t_SL g200 ( 
.A1(n_188),
.A2(n_199),
.B(n_183),
.Y(n_200)
);

NAND2xp5_ASAP7_75t_SL g209 ( 
.A(n_189),
.B(n_193),
.Y(n_209)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_172),
.Y(n_191)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_191),
.Y(n_202)
);

NOR2xp33_ASAP7_75t_L g205 ( 
.A(n_192),
.B(n_194),
.Y(n_205)
);

NAND2xp5_ASAP7_75t_SL g194 ( 
.A(n_174),
.B(n_164),
.Y(n_194)
);

NOR2xp33_ASAP7_75t_L g195 ( 
.A(n_186),
.B(n_158),
.Y(n_195)
);

CKINVDCx16_ASAP7_75t_R g201 ( 
.A(n_195),
.Y(n_201)
);

HB1xp67_ASAP7_75t_L g196 ( 
.A(n_171),
.Y(n_196)
);

NOR2xp33_ASAP7_75t_L g206 ( 
.A(n_196),
.B(n_197),
.Y(n_206)
);

NOR2xp33_ASAP7_75t_L g197 ( 
.A(n_175),
.B(n_158),
.Y(n_197)
);

NOR2xp33_ASAP7_75t_L g198 ( 
.A(n_179),
.B(n_153),
.Y(n_198)
);

BUFx3_ASAP7_75t_L g207 ( 
.A(n_198),
.Y(n_207)
);

MAJIxp5_ASAP7_75t_L g199 ( 
.A(n_185),
.B(n_156),
.C(n_153),
.Y(n_199)
);

NOR2xp33_ASAP7_75t_L g213 ( 
.A(n_200),
.B(n_150),
.Y(n_213)
);

AOI22xp5_ASAP7_75t_L g203 ( 
.A1(n_192),
.A2(n_170),
.B1(n_184),
.B2(n_185),
.Y(n_203)
);

AOI22xp33_ASAP7_75t_L g210 ( 
.A1(n_203),
.A2(n_190),
.B1(n_199),
.B2(n_131),
.Y(n_210)
);

NAND5xp2_ASAP7_75t_L g204 ( 
.A(n_189),
.B(n_182),
.C(n_155),
.D(n_178),
.E(n_173),
.Y(n_204)
);

NAND2xp5_ASAP7_75t_L g214 ( 
.A(n_204),
.B(n_129),
.Y(n_214)
);

AOI22xp5_ASAP7_75t_SL g208 ( 
.A1(n_187),
.A2(n_171),
.B1(n_147),
.B2(n_167),
.Y(n_208)
);

OAI21xp5_ASAP7_75t_L g216 ( 
.A1(n_208),
.A2(n_116),
.B(n_128),
.Y(n_216)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_210),
.Y(n_219)
);

MAJIxp5_ASAP7_75t_L g211 ( 
.A(n_200),
.B(n_190),
.C(n_140),
.Y(n_211)
);

MAJIxp5_ASAP7_75t_L g221 ( 
.A(n_211),
.B(n_215),
.C(n_202),
.Y(n_221)
);

OAI21xp5_ASAP7_75t_SL g212 ( 
.A1(n_209),
.A2(n_150),
.B(n_151),
.Y(n_212)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_212),
.Y(n_223)
);

NOR2xp33_ASAP7_75t_SL g218 ( 
.A(n_213),
.B(n_205),
.Y(n_218)
);

NAND2xp5_ASAP7_75t_SL g220 ( 
.A(n_214),
.B(n_216),
.Y(n_220)
);

MAJIxp5_ASAP7_75t_L g215 ( 
.A(n_207),
.B(n_108),
.C(n_119),
.Y(n_215)
);

XOR2xp5_ASAP7_75t_L g217 ( 
.A(n_203),
.B(n_121),
.Y(n_217)
);

MAJIxp5_ASAP7_75t_L g222 ( 
.A(n_217),
.B(n_206),
.C(n_208),
.Y(n_222)
);

AOI22xp5_ASAP7_75t_SL g226 ( 
.A1(n_218),
.A2(n_98),
.B1(n_151),
.B2(n_114),
.Y(n_226)
);

XNOR2xp5_ASAP7_75t_L g227 ( 
.A(n_221),
.B(n_166),
.Y(n_227)
);

XOR2xp5_ASAP7_75t_L g225 ( 
.A(n_222),
.B(n_207),
.Y(n_225)
);

AOI322xp5_ASAP7_75t_L g224 ( 
.A1(n_219),
.A2(n_204),
.A3(n_217),
.B1(n_201),
.B2(n_210),
.C1(n_211),
.C2(n_202),
.Y(n_224)
);

AOI22xp5_ASAP7_75t_SL g229 ( 
.A1(n_224),
.A2(n_227),
.B1(n_223),
.B2(n_220),
.Y(n_229)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_225),
.Y(n_228)
);

AOI31xp67_ASAP7_75t_SL g230 ( 
.A1(n_226),
.A2(n_166),
.A3(n_220),
.B(n_224),
.Y(n_230)
);

CKINVDCx20_ASAP7_75t_R g231 ( 
.A(n_229),
.Y(n_231)
);

NOR2xp33_ASAP7_75t_SL g232 ( 
.A(n_230),
.B(n_112),
.Y(n_232)
);

AOI22xp5_ASAP7_75t_L g233 ( 
.A1(n_232),
.A2(n_112),
.B1(n_228),
.B2(n_111),
.Y(n_233)
);

NAND2xp5_ASAP7_75t_SL g234 ( 
.A(n_233),
.B(n_231),
.Y(n_234)
);

XNOR2xp5_ASAP7_75t_L g235 ( 
.A(n_234),
.B(n_111),
.Y(n_235)
);


endmodule