module fake_jpeg_17307_n_319 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_319);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_319;

wire n_253;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_15;
wire n_141;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_51;
wire n_84;
wire n_59;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

BUFx6f_ASAP7_75t_L g15 ( 
.A(n_3),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_11),
.Y(n_16)
);

INVx1_ASAP7_75t_SL g17 ( 
.A(n_0),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_13),
.Y(n_18)
);

INVx6_ASAP7_75t_SL g19 ( 
.A(n_12),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_11),
.Y(n_20)
);

INVx11_ASAP7_75t_L g21 ( 
.A(n_12),
.Y(n_21)
);

BUFx12f_ASAP7_75t_L g22 ( 
.A(n_11),
.Y(n_22)
);

INVx13_ASAP7_75t_L g23 ( 
.A(n_10),
.Y(n_23)
);

CKINVDCx16_ASAP7_75t_R g24 ( 
.A(n_8),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_1),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_13),
.Y(n_26)
);

BUFx5_ASAP7_75t_L g27 ( 
.A(n_2),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_5),
.Y(n_28)
);

BUFx5_ASAP7_75t_L g29 ( 
.A(n_12),
.Y(n_29)
);

INVx3_ASAP7_75t_L g30 ( 
.A(n_0),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_6),
.Y(n_31)
);

INVx4_ASAP7_75t_L g32 ( 
.A(n_22),
.Y(n_32)
);

BUFx3_ASAP7_75t_L g55 ( 
.A(n_32),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_SL g33 ( 
.A(n_16),
.B(n_6),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_SL g44 ( 
.A(n_33),
.B(n_34),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g34 ( 
.A(n_17),
.B(n_6),
.Y(n_34)
);

BUFx4f_ASAP7_75t_SL g35 ( 
.A(n_22),
.Y(n_35)
);

INVx1_ASAP7_75t_SL g51 ( 
.A(n_35),
.Y(n_51)
);

BUFx12f_ASAP7_75t_L g36 ( 
.A(n_22),
.Y(n_36)
);

BUFx12f_ASAP7_75t_L g47 ( 
.A(n_36),
.Y(n_47)
);

INVx11_ASAP7_75t_L g37 ( 
.A(n_23),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_37),
.Y(n_46)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_30),
.Y(n_38)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_38),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_15),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_39),
.Y(n_48)
);

INVx4_ASAP7_75t_L g40 ( 
.A(n_22),
.Y(n_40)
);

INVx4_ASAP7_75t_L g53 ( 
.A(n_40),
.Y(n_53)
);

INVx2_ASAP7_75t_L g41 ( 
.A(n_38),
.Y(n_41)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_41),
.Y(n_61)
);

INVx2_ASAP7_75t_L g42 ( 
.A(n_38),
.Y(n_42)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_42),
.Y(n_69)
);

AND2x2_ASAP7_75t_L g43 ( 
.A(n_34),
.B(n_23),
.Y(n_43)
);

AOI21xp5_ASAP7_75t_L g80 ( 
.A1(n_43),
.A2(n_17),
.B(n_24),
.Y(n_80)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_33),
.Y(n_45)
);

NAND2xp5_ASAP7_75t_L g56 ( 
.A(n_45),
.B(n_34),
.Y(n_56)
);

MAJIxp5_ASAP7_75t_L g49 ( 
.A(n_35),
.B(n_22),
.C(n_29),
.Y(n_49)
);

AND2x2_ASAP7_75t_L g58 ( 
.A(n_49),
.B(n_54),
.Y(n_58)
);

INVx5_ASAP7_75t_L g52 ( 
.A(n_36),
.Y(n_52)
);

INVx5_ASAP7_75t_L g60 ( 
.A(n_52),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_SL g54 ( 
.A(n_33),
.B(n_18),
.Y(n_54)
);

OR2x2_ASAP7_75t_L g105 ( 
.A(n_56),
.B(n_20),
.Y(n_105)
);

A2O1A1Ixp33_ASAP7_75t_L g57 ( 
.A1(n_45),
.A2(n_20),
.B(n_31),
.C(n_28),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_L g90 ( 
.A(n_57),
.B(n_44),
.Y(n_90)
);

INVx8_ASAP7_75t_L g59 ( 
.A(n_47),
.Y(n_59)
);

INVx5_ASAP7_75t_L g99 ( 
.A(n_59),
.Y(n_99)
);

INVxp67_ASAP7_75t_L g62 ( 
.A(n_41),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_62),
.B(n_63),
.Y(n_87)
);

INVx6_ASAP7_75t_SL g63 ( 
.A(n_46),
.Y(n_63)
);

BUFx12_ASAP7_75t_L g64 ( 
.A(n_55),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_64),
.B(n_68),
.Y(n_102)
);

INVx5_ASAP7_75t_L g65 ( 
.A(n_52),
.Y(n_65)
);

INVx3_ASAP7_75t_L g101 ( 
.A(n_65),
.Y(n_101)
);

INVx4_ASAP7_75t_L g66 ( 
.A(n_46),
.Y(n_66)
);

BUFx3_ASAP7_75t_L g97 ( 
.A(n_66),
.Y(n_97)
);

BUFx12f_ASAP7_75t_L g67 ( 
.A(n_47),
.Y(n_67)
);

INVx4_ASAP7_75t_L g92 ( 
.A(n_67),
.Y(n_92)
);

INVx4_ASAP7_75t_L g68 ( 
.A(n_46),
.Y(n_68)
);

CKINVDCx12_ASAP7_75t_R g70 ( 
.A(n_55),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_70),
.B(n_71),
.Y(n_109)
);

INVx3_ASAP7_75t_SL g71 ( 
.A(n_48),
.Y(n_71)
);

INVx2_ASAP7_75t_L g72 ( 
.A(n_42),
.Y(n_72)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_72),
.Y(n_89)
);

AOI22xp5_ASAP7_75t_L g73 ( 
.A1(n_43),
.A2(n_30),
.B1(n_40),
.B2(n_32),
.Y(n_73)
);

OAI22xp5_ASAP7_75t_SL g95 ( 
.A1(n_73),
.A2(n_79),
.B1(n_37),
.B2(n_17),
.Y(n_95)
);

CKINVDCx20_ASAP7_75t_R g74 ( 
.A(n_50),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_74),
.B(n_75),
.Y(n_111)
);

INVx1_ASAP7_75t_SL g75 ( 
.A(n_43),
.Y(n_75)
);

INVx4_ASAP7_75t_L g76 ( 
.A(n_48),
.Y(n_76)
);

INVx4_ASAP7_75t_SL g86 ( 
.A(n_76),
.Y(n_86)
);

OAI22xp5_ASAP7_75t_SL g77 ( 
.A1(n_54),
.A2(n_30),
.B1(n_21),
.B2(n_31),
.Y(n_77)
);

OAI22xp5_ASAP7_75t_L g100 ( 
.A1(n_77),
.A2(n_18),
.B1(n_17),
.B2(n_20),
.Y(n_100)
);

INVx8_ASAP7_75t_L g78 ( 
.A(n_47),
.Y(n_78)
);

OAI22xp33_ASAP7_75t_SL g108 ( 
.A1(n_78),
.A2(n_37),
.B1(n_51),
.B2(n_53),
.Y(n_108)
);

AOI22xp33_ASAP7_75t_L g79 ( 
.A1(n_49),
.A2(n_30),
.B1(n_21),
.B2(n_32),
.Y(n_79)
);

AND2x2_ASAP7_75t_L g103 ( 
.A(n_80),
.B(n_18),
.Y(n_103)
);

INVx3_ASAP7_75t_L g81 ( 
.A(n_48),
.Y(n_81)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_81),
.Y(n_110)
);

INVx2_ASAP7_75t_L g82 ( 
.A(n_50),
.Y(n_82)
);

INVx2_ASAP7_75t_L g98 ( 
.A(n_82),
.Y(n_98)
);

BUFx6f_ASAP7_75t_L g83 ( 
.A(n_47),
.Y(n_83)
);

BUFx6f_ASAP7_75t_L g88 ( 
.A(n_83),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_44),
.B(n_31),
.Y(n_84)
);

INVxp67_ASAP7_75t_L g85 ( 
.A(n_84),
.Y(n_85)
);

OR2x2_ASAP7_75t_L g126 ( 
.A(n_90),
.B(n_105),
.Y(n_126)
);

MAJIxp5_ASAP7_75t_L g91 ( 
.A(n_75),
.B(n_35),
.C(n_36),
.Y(n_91)
);

MAJIxp5_ASAP7_75t_L g124 ( 
.A(n_91),
.B(n_35),
.C(n_36),
.Y(n_124)
);

AOI22xp33_ASAP7_75t_L g93 ( 
.A1(n_79),
.A2(n_21),
.B1(n_23),
.B2(n_40),
.Y(n_93)
);

OAI22xp5_ASAP7_75t_SL g118 ( 
.A1(n_93),
.A2(n_94),
.B1(n_96),
.B2(n_66),
.Y(n_118)
);

AOI22xp5_ASAP7_75t_L g94 ( 
.A1(n_58),
.A2(n_32),
.B1(n_40),
.B2(n_53),
.Y(n_94)
);

AOI22xp5_ASAP7_75t_L g137 ( 
.A1(n_95),
.A2(n_100),
.B1(n_24),
.B2(n_68),
.Y(n_137)
);

AOI22xp33_ASAP7_75t_L g96 ( 
.A1(n_73),
.A2(n_21),
.B1(n_23),
.B2(n_37),
.Y(n_96)
);

AND2x2_ASAP7_75t_L g134 ( 
.A(n_103),
.B(n_106),
.Y(n_134)
);

INVx13_ASAP7_75t_L g104 ( 
.A(n_64),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_L g138 ( 
.A(n_104),
.B(n_64),
.Y(n_138)
);

AND2x2_ASAP7_75t_L g106 ( 
.A(n_58),
.B(n_69),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_L g107 ( 
.A(n_57),
.B(n_53),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_L g128 ( 
.A(n_107),
.B(n_112),
.Y(n_128)
);

INVxp67_ASAP7_75t_L g129 ( 
.A(n_108),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_L g112 ( 
.A(n_62),
.B(n_51),
.Y(n_112)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_61),
.Y(n_113)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_113),
.Y(n_125)
);

AO22x2_ASAP7_75t_SL g114 ( 
.A1(n_95),
.A2(n_39),
.B1(n_35),
.B2(n_71),
.Y(n_114)
);

OAI22xp5_ASAP7_75t_SL g149 ( 
.A1(n_114),
.A2(n_86),
.B1(n_76),
.B2(n_99),
.Y(n_149)
);

AND2x6_ASAP7_75t_L g115 ( 
.A(n_106),
.B(n_14),
.Y(n_115)
);

CKINVDCx20_ASAP7_75t_R g146 ( 
.A(n_115),
.Y(n_146)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_113),
.Y(n_116)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_116),
.Y(n_153)
);

AOI22xp33_ASAP7_75t_SL g117 ( 
.A1(n_101),
.A2(n_60),
.B1(n_65),
.B2(n_51),
.Y(n_117)
);

OAI22xp5_ASAP7_75t_L g145 ( 
.A1(n_117),
.A2(n_118),
.B1(n_137),
.B2(n_86),
.Y(n_145)
);

CKINVDCx12_ASAP7_75t_R g119 ( 
.A(n_104),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_L g156 ( 
.A(n_119),
.B(n_133),
.Y(n_156)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_98),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_SL g142 ( 
.A(n_120),
.B(n_121),
.Y(n_142)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_98),
.Y(n_121)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_89),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_SL g151 ( 
.A(n_122),
.B(n_123),
.Y(n_151)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_87),
.Y(n_123)
);

MAJIxp5_ASAP7_75t_L g161 ( 
.A(n_124),
.B(n_127),
.C(n_36),
.Y(n_161)
);

MAJIxp5_ASAP7_75t_L g127 ( 
.A(n_91),
.B(n_35),
.C(n_36),
.Y(n_127)
);

INVx3_ASAP7_75t_L g130 ( 
.A(n_101),
.Y(n_130)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_130),
.Y(n_147)
);

CKINVDCx20_ASAP7_75t_R g131 ( 
.A(n_110),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_SL g155 ( 
.A(n_131),
.B(n_132),
.Y(n_155)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_110),
.Y(n_132)
);

NOR3xp33_ASAP7_75t_L g133 ( 
.A(n_90),
.B(n_60),
.C(n_28),
.Y(n_133)
);

INVx5_ASAP7_75t_L g135 ( 
.A(n_99),
.Y(n_135)
);

INVx5_ASAP7_75t_L g173 ( 
.A(n_135),
.Y(n_173)
);

AND2x2_ASAP7_75t_L g136 ( 
.A(n_94),
.B(n_0),
.Y(n_136)
);

OAI21xp5_ASAP7_75t_SL g165 ( 
.A1(n_136),
.A2(n_16),
.B(n_26),
.Y(n_165)
);

INVxp67_ASAP7_75t_L g171 ( 
.A(n_138),
.Y(n_171)
);

NOR2xp33_ASAP7_75t_L g139 ( 
.A(n_85),
.B(n_59),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_SL g169 ( 
.A(n_139),
.B(n_140),
.Y(n_169)
);

NOR2xp33_ASAP7_75t_L g140 ( 
.A(n_85),
.B(n_78),
.Y(n_140)
);

AOI21xp5_ASAP7_75t_L g141 ( 
.A1(n_128),
.A2(n_107),
.B(n_106),
.Y(n_141)
);

OAI21xp5_ASAP7_75t_SL g178 ( 
.A1(n_141),
.A2(n_144),
.B(n_165),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_L g143 ( 
.A(n_128),
.B(n_111),
.Y(n_143)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_143),
.Y(n_181)
);

AOI21xp5_ASAP7_75t_L g144 ( 
.A1(n_134),
.A2(n_136),
.B(n_129),
.Y(n_144)
);

AOI22xp5_ASAP7_75t_L g200 ( 
.A1(n_145),
.A2(n_19),
.B1(n_1),
.B2(n_2),
.Y(n_200)
);

AOI22xp5_ASAP7_75t_L g148 ( 
.A1(n_134),
.A2(n_103),
.B1(n_112),
.B2(n_81),
.Y(n_148)
);

OAI22xp5_ASAP7_75t_L g183 ( 
.A1(n_148),
.A2(n_149),
.B1(n_166),
.B2(n_92),
.Y(n_183)
);

XOR2x1_ASAP7_75t_SL g150 ( 
.A(n_134),
.B(n_103),
.Y(n_150)
);

OAI21xp5_ASAP7_75t_L g191 ( 
.A1(n_150),
.A2(n_157),
.B(n_158),
.Y(n_191)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_125),
.Y(n_152)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_152),
.Y(n_186)
);

OAI22xp5_ASAP7_75t_SL g154 ( 
.A1(n_114),
.A2(n_39),
.B1(n_105),
.B2(n_102),
.Y(n_154)
);

OAI22xp5_ASAP7_75t_SL g199 ( 
.A1(n_154),
.A2(n_148),
.B1(n_167),
.B2(n_166),
.Y(n_199)
);

OAI21xp5_ASAP7_75t_L g157 ( 
.A1(n_136),
.A2(n_109),
.B(n_24),
.Y(n_157)
);

OAI21xp5_ASAP7_75t_L g158 ( 
.A1(n_126),
.A2(n_26),
.B(n_28),
.Y(n_158)
);

XOR2xp5_ASAP7_75t_L g159 ( 
.A(n_124),
.B(n_35),
.Y(n_159)
);

MAJIxp5_ASAP7_75t_L g187 ( 
.A(n_159),
.B(n_161),
.C(n_162),
.Y(n_187)
);

CKINVDCx16_ASAP7_75t_R g160 ( 
.A(n_125),
.Y(n_160)
);

NOR2xp33_ASAP7_75t_L g175 ( 
.A(n_160),
.B(n_164),
.Y(n_175)
);

MAJIxp5_ASAP7_75t_L g162 ( 
.A(n_127),
.B(n_55),
.C(n_36),
.Y(n_162)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_130),
.Y(n_163)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_163),
.Y(n_188)
);

CKINVDCx20_ASAP7_75t_R g164 ( 
.A(n_126),
.Y(n_164)
);

AOI22xp5_ASAP7_75t_L g166 ( 
.A1(n_114),
.A2(n_39),
.B1(n_19),
.B2(n_25),
.Y(n_166)
);

MAJIxp5_ASAP7_75t_L g167 ( 
.A(n_118),
.B(n_67),
.C(n_83),
.Y(n_167)
);

MAJIxp5_ASAP7_75t_L g197 ( 
.A(n_167),
.B(n_97),
.C(n_22),
.Y(n_197)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_137),
.Y(n_168)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_168),
.Y(n_194)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_135),
.Y(n_170)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_170),
.Y(n_196)
);

CKINVDCx20_ASAP7_75t_R g172 ( 
.A(n_115),
.Y(n_172)
);

NOR2xp33_ASAP7_75t_L g190 ( 
.A(n_172),
.B(n_15),
.Y(n_190)
);

CKINVDCx20_ASAP7_75t_R g174 ( 
.A(n_155),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_L g218 ( 
.A(n_174),
.B(n_180),
.Y(n_218)
);

XNOR2xp5_ASAP7_75t_L g176 ( 
.A(n_141),
.B(n_129),
.Y(n_176)
);

MAJIxp5_ASAP7_75t_L g210 ( 
.A(n_176),
.B(n_185),
.C(n_189),
.Y(n_210)
);

NOR2xp33_ASAP7_75t_SL g177 ( 
.A(n_151),
.B(n_26),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_SL g211 ( 
.A(n_177),
.B(n_184),
.Y(n_211)
);

OR2x2_ASAP7_75t_L g179 ( 
.A(n_143),
.B(n_25),
.Y(n_179)
);

OAI21xp5_ASAP7_75t_L g207 ( 
.A1(n_179),
.A2(n_205),
.B(n_158),
.Y(n_207)
);

CKINVDCx20_ASAP7_75t_R g180 ( 
.A(n_142),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_L g182 ( 
.A(n_152),
.B(n_169),
.Y(n_182)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_182),
.Y(n_213)
);

A2O1A1Ixp33_ASAP7_75t_SL g224 ( 
.A1(n_183),
.A2(n_156),
.B(n_15),
.C(n_27),
.Y(n_224)
);

CKINVDCx20_ASAP7_75t_R g184 ( 
.A(n_153),
.Y(n_184)
);

XOR2xp5_ASAP7_75t_L g185 ( 
.A(n_150),
.B(n_92),
.Y(n_185)
);

XOR2xp5_ASAP7_75t_L g189 ( 
.A(n_161),
.B(n_67),
.Y(n_189)
);

OAI22xp5_ASAP7_75t_L g223 ( 
.A1(n_190),
.A2(n_193),
.B1(n_200),
.B2(n_173),
.Y(n_223)
);

OAI21xp5_ASAP7_75t_SL g192 ( 
.A1(n_144),
.A2(n_25),
.B(n_16),
.Y(n_192)
);

AOI21xp5_ASAP7_75t_L g214 ( 
.A1(n_192),
.A2(n_165),
.B(n_178),
.Y(n_214)
);

OAI22xp5_ASAP7_75t_L g193 ( 
.A1(n_168),
.A2(n_19),
.B1(n_15),
.B2(n_39),
.Y(n_193)
);

NOR2xp33_ASAP7_75t_L g195 ( 
.A(n_147),
.B(n_97),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_SL g221 ( 
.A(n_195),
.B(n_198),
.Y(n_221)
);

MAJIxp5_ASAP7_75t_L g222 ( 
.A(n_197),
.B(n_162),
.C(n_149),
.Y(n_222)
);

NOR2xp33_ASAP7_75t_L g198 ( 
.A(n_147),
.B(n_88),
.Y(n_198)
);

NOR2xp33_ASAP7_75t_L g209 ( 
.A(n_199),
.B(n_201),
.Y(n_209)
);

CKINVDCx20_ASAP7_75t_R g201 ( 
.A(n_163),
.Y(n_201)
);

NOR2xp33_ASAP7_75t_L g202 ( 
.A(n_171),
.B(n_88),
.Y(n_202)
);

NOR2xp33_ASAP7_75t_L g216 ( 
.A(n_202),
.B(n_203),
.Y(n_216)
);

NAND2xp5_ASAP7_75t_L g203 ( 
.A(n_171),
.B(n_22),
.Y(n_203)
);

XNOR2xp5_ASAP7_75t_SL g204 ( 
.A(n_157),
.B(n_29),
.Y(n_204)
);

XOR2xp5_ASAP7_75t_L g220 ( 
.A(n_204),
.B(n_192),
.Y(n_220)
);

OAI21xp5_ASAP7_75t_L g205 ( 
.A1(n_146),
.A2(n_29),
.B(n_27),
.Y(n_205)
);

CKINVDCx20_ASAP7_75t_R g206 ( 
.A(n_170),
.Y(n_206)
);

NOR2xp33_ASAP7_75t_L g217 ( 
.A(n_206),
.B(n_173),
.Y(n_217)
);

NAND2xp5_ASAP7_75t_SL g237 ( 
.A(n_207),
.B(n_208),
.Y(n_237)
);

CKINVDCx20_ASAP7_75t_R g208 ( 
.A(n_186),
.Y(n_208)
);

AND2x2_ASAP7_75t_L g212 ( 
.A(n_185),
.B(n_159),
.Y(n_212)
);

OAI21xp5_ASAP7_75t_SL g242 ( 
.A1(n_212),
.A2(n_214),
.B(n_178),
.Y(n_242)
);

HB1xp67_ASAP7_75t_L g215 ( 
.A(n_188),
.Y(n_215)
);

BUFx2_ASAP7_75t_L g246 ( 
.A(n_215),
.Y(n_246)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_217),
.Y(n_238)
);

NOR2xp33_ASAP7_75t_L g219 ( 
.A(n_206),
.B(n_154),
.Y(n_219)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_219),
.Y(n_251)
);

MAJIxp5_ASAP7_75t_L g234 ( 
.A(n_220),
.B(n_222),
.C(n_226),
.Y(n_234)
);

CKINVDCx16_ASAP7_75t_R g233 ( 
.A(n_223),
.Y(n_233)
);

OAI22xp5_ASAP7_75t_SL g239 ( 
.A1(n_224),
.A2(n_194),
.B1(n_203),
.B2(n_196),
.Y(n_239)
);

BUFx12_ASAP7_75t_L g225 ( 
.A(n_188),
.Y(n_225)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_225),
.Y(n_235)
);

MAJIxp5_ASAP7_75t_L g226 ( 
.A(n_187),
.B(n_27),
.C(n_0),
.Y(n_226)
);

NOR2xp33_ASAP7_75t_L g227 ( 
.A(n_175),
.B(n_1),
.Y(n_227)
);

NAND2xp5_ASAP7_75t_SL g249 ( 
.A(n_227),
.B(n_228),
.Y(n_249)
);

OAI22xp5_ASAP7_75t_L g228 ( 
.A1(n_200),
.A2(n_2),
.B1(n_3),
.B2(n_4),
.Y(n_228)
);

NOR2xp33_ASAP7_75t_L g229 ( 
.A(n_181),
.B(n_3),
.Y(n_229)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_229),
.Y(n_236)
);

MAJIxp5_ASAP7_75t_L g230 ( 
.A(n_187),
.B(n_4),
.C(n_5),
.Y(n_230)
);

MAJIxp5_ASAP7_75t_L g240 ( 
.A(n_230),
.B(n_231),
.C(n_191),
.Y(n_240)
);

XNOR2xp5_ASAP7_75t_L g231 ( 
.A(n_176),
.B(n_4),
.Y(n_231)
);

NAND2xp5_ASAP7_75t_L g232 ( 
.A(n_213),
.B(n_181),
.Y(n_232)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_232),
.Y(n_266)
);

CKINVDCx14_ASAP7_75t_R g257 ( 
.A(n_239),
.Y(n_257)
);

MAJIxp5_ASAP7_75t_L g261 ( 
.A(n_240),
.B(n_220),
.C(n_204),
.Y(n_261)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_221),
.Y(n_241)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_241),
.Y(n_267)
);

AO21x1_ASAP7_75t_L g268 ( 
.A1(n_242),
.A2(n_250),
.B(n_191),
.Y(n_268)
);

AOI22xp5_ASAP7_75t_L g243 ( 
.A1(n_209),
.A2(n_212),
.B1(n_222),
.B2(n_194),
.Y(n_243)
);

AOI22xp5_ASAP7_75t_L g256 ( 
.A1(n_243),
.A2(n_212),
.B1(n_197),
.B2(n_230),
.Y(n_256)
);

INVx1_ASAP7_75t_SL g244 ( 
.A(n_225),
.Y(n_244)
);

NOR2xp33_ASAP7_75t_L g258 ( 
.A(n_244),
.B(n_248),
.Y(n_258)
);

NAND2xp5_ASAP7_75t_L g245 ( 
.A(n_216),
.B(n_182),
.Y(n_245)
);

CKINVDCx20_ASAP7_75t_R g260 ( 
.A(n_245),
.Y(n_260)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_218),
.Y(n_247)
);

CKINVDCx20_ASAP7_75t_R g265 ( 
.A(n_247),
.Y(n_265)
);

NAND2xp5_ASAP7_75t_L g248 ( 
.A(n_207),
.B(n_186),
.Y(n_248)
);

OR2x2_ASAP7_75t_L g250 ( 
.A(n_225),
.B(n_196),
.Y(n_250)
);

XOR2xp5_ASAP7_75t_L g252 ( 
.A(n_242),
.B(n_210),
.Y(n_252)
);

XOR2xp5_ASAP7_75t_L g271 ( 
.A(n_252),
.B(n_253),
.Y(n_271)
);

XOR2xp5_ASAP7_75t_L g253 ( 
.A(n_243),
.B(n_210),
.Y(n_253)
);

HB1xp67_ASAP7_75t_L g254 ( 
.A(n_233),
.Y(n_254)
);

BUFx2_ASAP7_75t_L g269 ( 
.A(n_254),
.Y(n_269)
);

MAJIxp5_ASAP7_75t_L g255 ( 
.A(n_234),
.B(n_189),
.C(n_226),
.Y(n_255)
);

MAJIxp5_ASAP7_75t_L g273 ( 
.A(n_255),
.B(n_259),
.C(n_240),
.Y(n_273)
);

XOR2xp5_ASAP7_75t_L g276 ( 
.A(n_256),
.B(n_264),
.Y(n_276)
);

MAJIxp5_ASAP7_75t_L g259 ( 
.A(n_234),
.B(n_231),
.C(n_199),
.Y(n_259)
);

MAJIxp5_ASAP7_75t_L g280 ( 
.A(n_261),
.B(n_262),
.C(n_263),
.Y(n_280)
);

XNOR2xp5_ASAP7_75t_L g262 ( 
.A(n_237),
.B(n_214),
.Y(n_262)
);

MAJIxp5_ASAP7_75t_L g263 ( 
.A(n_241),
.B(n_247),
.C(n_238),
.Y(n_263)
);

XOR2xp5_ASAP7_75t_L g264 ( 
.A(n_248),
.B(n_205),
.Y(n_264)
);

NAND2xp5_ASAP7_75t_L g282 ( 
.A(n_268),
.B(n_179),
.Y(n_282)
);

NOR2xp33_ASAP7_75t_L g270 ( 
.A(n_265),
.B(n_244),
.Y(n_270)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_270),
.Y(n_284)
);

AOI22xp5_ASAP7_75t_L g272 ( 
.A1(n_257),
.A2(n_251),
.B1(n_235),
.B2(n_245),
.Y(n_272)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_272),
.Y(n_289)
);

MAJIxp5_ASAP7_75t_L g292 ( 
.A(n_273),
.B(n_5),
.C(n_7),
.Y(n_292)
);

AOI322xp5_ASAP7_75t_L g274 ( 
.A1(n_267),
.A2(n_246),
.A3(n_249),
.B1(n_235),
.B2(n_232),
.C1(n_224),
.C2(n_236),
.Y(n_274)
);

NOR2xp33_ASAP7_75t_L g286 ( 
.A(n_274),
.B(n_279),
.Y(n_286)
);

NOR2xp33_ASAP7_75t_L g275 ( 
.A(n_260),
.B(n_246),
.Y(n_275)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_275),
.Y(n_290)
);

NOR2xp33_ASAP7_75t_L g277 ( 
.A(n_258),
.B(n_236),
.Y(n_277)
);

NAND2xp5_ASAP7_75t_L g288 ( 
.A(n_277),
.B(n_278),
.Y(n_288)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_266),
.Y(n_278)
);

AOI22xp5_ASAP7_75t_L g279 ( 
.A1(n_259),
.A2(n_250),
.B1(n_224),
.B2(n_239),
.Y(n_279)
);

AND2x2_ASAP7_75t_L g281 ( 
.A(n_264),
.B(n_224),
.Y(n_281)
);

AOI21xp5_ASAP7_75t_L g287 ( 
.A1(n_281),
.A2(n_282),
.B(n_253),
.Y(n_287)
);

INVx6_ASAP7_75t_L g283 ( 
.A(n_269),
.Y(n_283)
);

NAND2xp5_ASAP7_75t_L g303 ( 
.A(n_283),
.B(n_293),
.Y(n_303)
);

AOI22xp5_ASAP7_75t_L g285 ( 
.A1(n_281),
.A2(n_268),
.B1(n_255),
.B2(n_252),
.Y(n_285)
);

AND2x2_ASAP7_75t_L g299 ( 
.A(n_285),
.B(n_271),
.Y(n_299)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_287),
.Y(n_298)
);

XNOR2xp5_ASAP7_75t_L g291 ( 
.A(n_273),
.B(n_211),
.Y(n_291)
);

XOR2xp5_ASAP7_75t_L g300 ( 
.A(n_291),
.B(n_292),
.Y(n_300)
);

NAND2xp5_ASAP7_75t_L g293 ( 
.A(n_280),
.B(n_7),
.Y(n_293)
);

OAI21xp5_ASAP7_75t_SL g294 ( 
.A1(n_269),
.A2(n_7),
.B(n_8),
.Y(n_294)
);

XOR2xp5_ASAP7_75t_L g301 ( 
.A(n_294),
.B(n_288),
.Y(n_301)
);

XNOR2xp5_ASAP7_75t_L g295 ( 
.A(n_291),
.B(n_276),
.Y(n_295)
);

NAND2xp5_ASAP7_75t_SL g305 ( 
.A(n_295),
.B(n_297),
.Y(n_305)
);

INVxp67_ASAP7_75t_L g296 ( 
.A(n_286),
.Y(n_296)
);

NAND2xp5_ASAP7_75t_L g306 ( 
.A(n_296),
.B(n_301),
.Y(n_306)
);

NOR2xp33_ASAP7_75t_SL g297 ( 
.A(n_284),
.B(n_276),
.Y(n_297)
);

OAI21xp5_ASAP7_75t_L g309 ( 
.A1(n_299),
.A2(n_283),
.B(n_9),
.Y(n_309)
);

AOI22xp5_ASAP7_75t_L g302 ( 
.A1(n_289),
.A2(n_271),
.B1(n_9),
.B2(n_10),
.Y(n_302)
);

INVxp33_ASAP7_75t_L g307 ( 
.A(n_302),
.Y(n_307)
);

AOI31xp67_ASAP7_75t_L g304 ( 
.A1(n_300),
.A2(n_292),
.A3(n_290),
.B(n_287),
.Y(n_304)
);

NAND2xp5_ASAP7_75t_L g311 ( 
.A(n_304),
.B(n_308),
.Y(n_311)
);

NOR2xp33_ASAP7_75t_SL g308 ( 
.A(n_303),
.B(n_285),
.Y(n_308)
);

XNOR2xp5_ASAP7_75t_L g312 ( 
.A(n_309),
.B(n_298),
.Y(n_312)
);

HB1xp67_ASAP7_75t_L g310 ( 
.A(n_306),
.Y(n_310)
);

NAND2xp5_ASAP7_75t_L g313 ( 
.A(n_310),
.B(n_312),
.Y(n_313)
);

AOI322xp5_ASAP7_75t_L g314 ( 
.A1(n_313),
.A2(n_311),
.A3(n_305),
.B1(n_307),
.B2(n_299),
.C1(n_296),
.C2(n_14),
.Y(n_314)
);

OAI21xp5_ASAP7_75t_L g315 ( 
.A1(n_314),
.A2(n_8),
.B(n_9),
.Y(n_315)
);

AND2x2_ASAP7_75t_L g316 ( 
.A(n_315),
.B(n_10),
.Y(n_316)
);

AOI21xp5_ASAP7_75t_SL g317 ( 
.A1(n_316),
.A2(n_13),
.B(n_14),
.Y(n_317)
);

BUFx24_ASAP7_75t_SL g318 ( 
.A(n_317),
.Y(n_318)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_318),
.Y(n_319)
);


endmodule