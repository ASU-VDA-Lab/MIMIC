module fake_netlist_6_2637_n_1054 (n_52, n_16, n_1, n_91, n_119, n_46, n_146, n_163, n_18, n_21, n_193, n_147, n_154, n_191, n_88, n_3, n_98, n_113, n_39, n_63, n_73, n_4, n_148, n_199, n_138, n_22, n_161, n_68, n_166, n_28, n_184, n_50, n_158, n_49, n_7, n_83, n_5, n_101, n_167, n_144, n_174, n_127, n_125, n_153, n_168, n_178, n_77, n_156, n_149, n_152, n_106, n_92, n_145, n_42, n_133, n_96, n_8, n_90, n_160, n_24, n_105, n_131, n_54, n_132, n_188, n_102, n_186, n_0, n_87, n_195, n_189, n_32, n_66, n_85, n_99, n_78, n_84, n_130, n_164, n_100, n_129, n_13, n_121, n_197, n_11, n_137, n_17, n_23, n_142, n_20, n_143, n_2, n_180, n_19, n_47, n_62, n_29, n_155, n_75, n_109, n_150, n_122, n_45, n_34, n_140, n_70, n_120, n_37, n_15, n_67, n_33, n_82, n_27, n_38, n_110, n_151, n_61, n_112, n_172, n_81, n_59, n_181, n_76, n_36, n_182, n_26, n_124, n_55, n_126, n_94, n_97, n_108, n_58, n_116, n_64, n_117, n_118, n_175, n_48, n_65, n_25, n_40, n_93, n_80, n_141, n_135, n_196, n_200, n_165, n_139, n_41, n_134, n_177, n_176, n_114, n_86, n_198, n_104, n_95, n_179, n_9, n_107, n_10, n_71, n_74, n_6, n_190, n_14, n_123, n_136, n_72, n_187, n_89, n_173, n_103, n_111, n_60, n_159, n_157, n_162, n_170, n_185, n_35, n_183, n_115, n_12, n_69, n_128, n_30, n_79, n_43, n_194, n_171, n_31, n_192, n_57, n_169, n_53, n_51, n_44, n_56, n_1054);

input n_52;
input n_16;
input n_1;
input n_91;
input n_119;
input n_46;
input n_146;
input n_163;
input n_18;
input n_21;
input n_193;
input n_147;
input n_154;
input n_191;
input n_88;
input n_3;
input n_98;
input n_113;
input n_39;
input n_63;
input n_73;
input n_4;
input n_148;
input n_199;
input n_138;
input n_22;
input n_161;
input n_68;
input n_166;
input n_28;
input n_184;
input n_50;
input n_158;
input n_49;
input n_7;
input n_83;
input n_5;
input n_101;
input n_167;
input n_144;
input n_174;
input n_127;
input n_125;
input n_153;
input n_168;
input n_178;
input n_77;
input n_156;
input n_149;
input n_152;
input n_106;
input n_92;
input n_145;
input n_42;
input n_133;
input n_96;
input n_8;
input n_90;
input n_160;
input n_24;
input n_105;
input n_131;
input n_54;
input n_132;
input n_188;
input n_102;
input n_186;
input n_0;
input n_87;
input n_195;
input n_189;
input n_32;
input n_66;
input n_85;
input n_99;
input n_78;
input n_84;
input n_130;
input n_164;
input n_100;
input n_129;
input n_13;
input n_121;
input n_197;
input n_11;
input n_137;
input n_17;
input n_23;
input n_142;
input n_20;
input n_143;
input n_2;
input n_180;
input n_19;
input n_47;
input n_62;
input n_29;
input n_155;
input n_75;
input n_109;
input n_150;
input n_122;
input n_45;
input n_34;
input n_140;
input n_70;
input n_120;
input n_37;
input n_15;
input n_67;
input n_33;
input n_82;
input n_27;
input n_38;
input n_110;
input n_151;
input n_61;
input n_112;
input n_172;
input n_81;
input n_59;
input n_181;
input n_76;
input n_36;
input n_182;
input n_26;
input n_124;
input n_55;
input n_126;
input n_94;
input n_97;
input n_108;
input n_58;
input n_116;
input n_64;
input n_117;
input n_118;
input n_175;
input n_48;
input n_65;
input n_25;
input n_40;
input n_93;
input n_80;
input n_141;
input n_135;
input n_196;
input n_200;
input n_165;
input n_139;
input n_41;
input n_134;
input n_177;
input n_176;
input n_114;
input n_86;
input n_198;
input n_104;
input n_95;
input n_179;
input n_9;
input n_107;
input n_10;
input n_71;
input n_74;
input n_6;
input n_190;
input n_14;
input n_123;
input n_136;
input n_72;
input n_187;
input n_89;
input n_173;
input n_103;
input n_111;
input n_60;
input n_159;
input n_157;
input n_162;
input n_170;
input n_185;
input n_35;
input n_183;
input n_115;
input n_12;
input n_69;
input n_128;
input n_30;
input n_79;
input n_43;
input n_194;
input n_171;
input n_31;
input n_192;
input n_57;
input n_169;
input n_53;
input n_51;
input n_44;
input n_56;

output n_1054;

wire n_992;
wire n_591;
wire n_435;
wire n_793;
wire n_326;
wire n_801;
wire n_256;
wire n_853;
wire n_440;
wire n_587;
wire n_695;
wire n_507;
wire n_968;
wire n_909;
wire n_580;
wire n_762;
wire n_1030;
wire n_881;
wire n_875;
wire n_209;
wire n_367;
wire n_465;
wire n_680;
wire n_741;
wire n_760;
wire n_1008;
wire n_1027;
wire n_590;
wire n_625;
wire n_661;
wire n_223;
wire n_278;
wire n_362;
wire n_341;
wire n_226;
wire n_828;
wire n_208;
wire n_462;
wire n_607;
wire n_671;
wire n_726;
wire n_1033;
wire n_316;
wire n_419;
wire n_304;
wire n_212;
wire n_700;
wire n_694;
wire n_933;
wire n_740;
wire n_1038;
wire n_578;
wire n_703;
wire n_1003;
wire n_365;
wire n_978;
wire n_384;
wire n_297;
wire n_627;
wire n_595;
wire n_524;
wire n_342;
wire n_820;
wire n_1044;
wire n_951;
wire n_783;
wire n_725;
wire n_952;
wire n_999;
wire n_358;
wire n_751;
wire n_449;
wire n_749;
wire n_798;
wire n_310;
wire n_509;
wire n_245;
wire n_368;
wire n_575;
wire n_994;
wire n_677;
wire n_969;
wire n_988;
wire n_805;
wire n_396;
wire n_495;
wire n_815;
wire n_350;
wire n_585;
wire n_732;
wire n_974;
wire n_568;
wire n_392;
wire n_840;
wire n_442;
wire n_480;
wire n_874;
wire n_724;
wire n_382;
wire n_673;
wire n_1020;
wire n_1009;
wire n_1042;
wire n_628;
wire n_883;
wire n_557;
wire n_823;
wire n_349;
wire n_643;
wire n_233;
wire n_617;
wire n_698;
wire n_898;
wire n_1032;
wire n_845;
wire n_255;
wire n_807;
wire n_1036;
wire n_739;
wire n_284;
wire n_400;
wire n_955;
wire n_337;
wire n_865;
wire n_893;
wire n_214;
wire n_925;
wire n_485;
wire n_1026;
wire n_443;
wire n_246;
wire n_892;
wire n_768;
wire n_471;
wire n_289;
wire n_935;
wire n_421;
wire n_781;
wire n_424;
wire n_789;
wire n_615;
wire n_238;
wire n_573;
wire n_769;
wire n_202;
wire n_320;
wire n_639;
wire n_676;
wire n_327;
wire n_794;
wire n_963;
wire n_727;
wire n_894;
wire n_369;
wire n_597;
wire n_685;
wire n_280;
wire n_287;
wire n_832;
wire n_353;
wire n_610;
wire n_555;
wire n_389;
wire n_814;
wire n_415;
wire n_830;
wire n_230;
wire n_605;
wire n_461;
wire n_873;
wire n_383;
wire n_826;
wire n_1024;
wire n_669;
wire n_447;
wire n_872;
wire n_300;
wire n_222;
wire n_248;
wire n_517;
wire n_718;
wire n_1018;
wire n_852;
wire n_747;
wire n_667;
wire n_229;
wire n_542;
wire n_847;
wire n_644;
wire n_682;
wire n_851;
wire n_621;
wire n_305;
wire n_1037;
wire n_721;
wire n_996;
wire n_750;
wire n_532;
wire n_742;
wire n_535;
wire n_691;
wire n_250;
wire n_372;
wire n_468;
wire n_544;
wire n_901;
wire n_504;
wire n_923;
wire n_314;
wire n_378;
wire n_413;
wire n_377;
wire n_791;
wire n_510;
wire n_837;
wire n_836;
wire n_1015;
wire n_863;
wire n_375;
wire n_601;
wire n_338;
wire n_522;
wire n_948;
wire n_466;
wire n_704;
wire n_918;
wire n_748;
wire n_506;
wire n_763;
wire n_360;
wire n_945;
wire n_977;
wire n_603;
wire n_1005;
wire n_991;
wire n_957;
wire n_235;
wire n_536;
wire n_895;
wire n_866;
wire n_622;
wire n_340;
wire n_710;
wire n_387;
wire n_452;
wire n_616;
wire n_658;
wire n_744;
wire n_971;
wire n_946;
wire n_344;
wire n_581;
wire n_428;
wire n_785;
wire n_761;
wire n_746;
wire n_609;
wire n_765;
wire n_432;
wire n_987;
wire n_641;
wire n_822;
wire n_693;
wire n_631;
wire n_516;
wire n_720;
wire n_758;
wire n_525;
wire n_842;
wire n_611;
wire n_943;
wire n_491;
wire n_878;
wire n_656;
wire n_772;
wire n_843;
wire n_989;
wire n_797;
wire n_666;
wire n_1016;
wire n_371;
wire n_795;
wire n_940;
wire n_770;
wire n_567;
wire n_899;
wire n_738;
wire n_405;
wire n_213;
wire n_538;
wire n_1035;
wire n_294;
wire n_302;
wire n_499;
wire n_380;
wire n_838;
wire n_705;
wire n_647;
wire n_844;
wire n_343;
wire n_953;
wire n_448;
wire n_886;
wire n_1004;
wire n_1017;
wire n_494;
wire n_539;
wire n_493;
wire n_397;
wire n_1022;
wire n_614;
wire n_529;
wire n_445;
wire n_425;
wire n_684;
wire n_930;
wire n_888;
wire n_454;
wire n_218;
wire n_638;
wire n_234;
wire n_910;
wire n_486;
wire n_911;
wire n_381;
wire n_947;
wire n_236;
wire n_653;
wire n_887;
wire n_752;
wire n_908;
wire n_944;
wire n_713;
wire n_648;
wire n_657;
wire n_1049;
wire n_576;
wire n_1028;
wire n_472;
wire n_270;
wire n_239;
wire n_414;
wire n_563;
wire n_782;
wire n_976;
wire n_490;
wire n_803;
wire n_290;
wire n_220;
wire n_809;
wire n_1043;
wire n_1011;
wire n_224;
wire n_926;
wire n_927;
wire n_839;
wire n_986;
wire n_734;
wire n_708;
wire n_919;
wire n_402;
wire n_352;
wire n_917;
wire n_668;
wire n_478;
wire n_626;
wire n_990;
wire n_574;
wire n_800;
wire n_779;
wire n_929;
wire n_460;
wire n_907;
wire n_854;
wire n_417;
wire n_446;
wire n_498;
wire n_662;
wire n_374;
wire n_659;
wire n_709;
wire n_904;
wire n_366;
wire n_870;
wire n_777;
wire n_407;
wire n_913;
wire n_450;
wire n_808;
wire n_867;
wire n_272;
wire n_526;
wire n_921;
wire n_712;
wire n_348;
wire n_711;
wire n_579;
wire n_376;
wire n_937;
wire n_390;
wire n_473;
wire n_293;
wire n_334;
wire n_559;
wire n_370;
wire n_458;
wire n_232;
wire n_650;
wire n_998;
wire n_1046;
wire n_717;
wire n_330;
wire n_771;
wire n_470;
wire n_475;
wire n_924;
wire n_298;
wire n_492;
wire n_972;
wire n_281;
wire n_258;
wire n_551;
wire n_699;
wire n_456;
wire n_564;
wire n_260;
wire n_265;
wire n_313;
wire n_451;
wire n_624;
wire n_824;
wire n_962;
wire n_1000;
wire n_279;
wire n_686;
wire n_796;
wire n_1041;
wire n_252;
wire n_757;
wire n_228;
wire n_565;
wire n_594;
wire n_719;
wire n_356;
wire n_577;
wire n_936;
wire n_552;
wire n_619;
wire n_885;
wire n_216;
wire n_455;
wire n_896;
wire n_521;
wire n_363;
wire n_572;
wire n_912;
wire n_395;
wire n_813;
wire n_592;
wire n_745;
wire n_654;
wire n_323;
wire n_829;
wire n_606;
wire n_393;
wire n_818;
wire n_984;
wire n_411;
wire n_503;
wire n_716;
wire n_623;
wire n_1048;
wire n_884;
wire n_599;
wire n_513;
wire n_855;
wire n_776;
wire n_321;
wire n_645;
wire n_331;
wire n_916;
wire n_227;
wire n_868;
wire n_570;
wire n_731;
wire n_859;
wire n_406;
wire n_483;
wire n_735;
wire n_204;
wire n_482;
wire n_934;
wire n_755;
wire n_931;
wire n_1021;
wire n_474;
wire n_527;
wire n_261;
wire n_608;
wire n_620;
wire n_420;
wire n_683;
wire n_630;
wire n_394;
wire n_312;
wire n_519;
wire n_541;
wire n_512;
wire n_958;
wire n_292;
wire n_307;
wire n_469;
wire n_433;
wire n_500;
wire n_942;
wire n_792;
wire n_880;
wire n_476;
wire n_981;
wire n_714;
wire n_291;
wire n_219;
wire n_543;
wire n_889;
wire n_357;
wire n_264;
wire n_263;
wire n_985;
wire n_589;
wire n_860;
wire n_481;
wire n_788;
wire n_819;
wire n_939;
wire n_997;
wire n_821;
wire n_325;
wire n_938;
wire n_767;
wire n_804;
wire n_329;
wire n_464;
wire n_600;
wire n_831;
wire n_802;
wire n_964;
wire n_982;
wire n_561;
wire n_477;
wire n_549;
wire n_980;
wire n_533;
wire n_954;
wire n_408;
wire n_932;
wire n_806;
wire n_864;
wire n_879;
wire n_959;
wire n_237;
wire n_584;
wire n_244;
wire n_399;
wire n_243;
wire n_979;
wire n_548;
wire n_905;
wire n_282;
wire n_436;
wire n_833;
wire n_211;
wire n_523;
wire n_322;
wire n_707;
wire n_993;
wire n_345;
wire n_409;
wire n_231;
wire n_354;
wire n_689;
wire n_799;
wire n_505;
wire n_240;
wire n_756;
wire n_319;
wire n_547;
wire n_537;
wire n_273;
wire n_558;
wire n_810;
wire n_635;
wire n_787;
wire n_311;
wire n_403;
wire n_723;
wire n_253;
wire n_634;
wire n_1051;
wire n_583;
wire n_596;
wire n_966;
wire n_546;
wire n_562;
wire n_249;
wire n_201;
wire n_386;
wire n_764;
wire n_1039;
wire n_556;
wire n_1034;
wire n_692;
wire n_733;
wire n_754;
wire n_941;
wire n_975;
wire n_1031;
wire n_487;
wire n_550;
wire n_241;
wire n_275;
wire n_553;
wire n_652;
wire n_970;
wire n_849;
wire n_560;
wire n_1014;
wire n_753;
wire n_642;
wire n_995;
wire n_276;
wire n_569;
wire n_441;
wire n_221;
wire n_811;
wire n_882;
wire n_444;
wire n_586;
wire n_423;
wire n_737;
wire n_318;
wire n_303;
wire n_511;
wire n_715;
wire n_467;
wire n_306;
wire n_269;
wire n_359;
wire n_973;
wire n_346;
wire n_416;
wire n_1053;
wire n_530;
wire n_277;
wire n_520;
wire n_1029;
wire n_418;
wire n_618;
wire n_790;
wire n_582;
wire n_266;
wire n_296;
wire n_861;
wire n_674;
wire n_857;
wire n_871;
wire n_967;
wire n_775;
wire n_922;
wire n_571;
wire n_268;
wire n_271;
wire n_404;
wire n_651;
wire n_439;
wire n_217;
wire n_210;
wire n_299;
wire n_518;
wire n_206;
wire n_679;
wire n_453;
wire n_612;
wire n_633;
wire n_665;
wire n_902;
wire n_333;
wire n_588;
wire n_215;
wire n_247;
wire n_225;
wire n_308;
wire n_309;
wire n_914;
wire n_759;
wire n_1047;
wire n_1010;
wire n_355;
wire n_426;
wire n_317;
wire n_1040;
wire n_915;
wire n_632;
wire n_702;
wire n_431;
wire n_347;
wire n_812;
wire n_459;
wire n_1052;
wire n_502;
wire n_328;
wire n_672;
wire n_534;
wire n_488;
wire n_429;
wire n_1006;
wire n_373;
wire n_1012;
wire n_285;
wire n_497;
wire n_780;
wire n_773;
wire n_675;
wire n_903;
wire n_257;
wire n_920;
wire n_730;
wire n_655;
wire n_706;
wire n_1045;
wire n_786;
wire n_670;
wire n_203;
wire n_286;
wire n_254;
wire n_207;
wire n_834;
wire n_242;
wire n_928;
wire n_835;
wire n_690;
wire n_850;
wire n_401;
wire n_324;
wire n_743;
wire n_766;
wire n_816;
wire n_335;
wire n_430;
wire n_1002;
wire n_463;
wire n_545;
wire n_489;
wire n_877;
wire n_205;
wire n_604;
wire n_848;
wire n_251;
wire n_1019;
wire n_301;
wire n_274;
wire n_636;
wire n_825;
wire n_728;
wire n_681;
wire n_729;
wire n_876;
wire n_774;
wire n_412;
wire n_640;
wire n_660;
wire n_965;
wire n_267;
wire n_438;
wire n_339;
wire n_784;
wire n_315;
wire n_434;
wire n_515;
wire n_983;
wire n_288;
wire n_427;
wire n_479;
wire n_496;
wire n_598;
wire n_422;
wire n_696;
wire n_906;
wire n_722;
wire n_688;
wire n_961;
wire n_862;
wire n_351;
wire n_869;
wire n_437;
wire n_259;
wire n_540;
wire n_593;
wire n_514;
wire n_646;
wire n_528;
wire n_391;
wire n_457;
wire n_687;
wire n_697;
wire n_364;
wire n_890;
wire n_637;
wire n_295;
wire n_385;
wire n_701;
wire n_817;
wire n_950;
wire n_629;
wire n_388;
wire n_858;
wire n_262;
wire n_484;
wire n_613;
wire n_736;
wire n_897;
wire n_900;
wire n_846;
wire n_501;
wire n_956;
wire n_960;
wire n_841;
wire n_531;
wire n_827;
wire n_1001;
wire n_508;
wire n_361;
wire n_663;
wire n_856;
wire n_1050;
wire n_379;
wire n_778;
wire n_1025;
wire n_332;
wire n_891;
wire n_336;
wire n_398;
wire n_410;
wire n_566;
wire n_554;
wire n_602;
wire n_1013;
wire n_1023;
wire n_664;
wire n_949;
wire n_678;
wire n_1007;
wire n_649;
wire n_283;

CKINVDCx5p33_ASAP7_75t_R g201 ( 
.A(n_195),
.Y(n_201)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_99),
.Y(n_202)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_154),
.Y(n_203)
);

CKINVDCx14_ASAP7_75t_R g204 ( 
.A(n_179),
.Y(n_204)
);

BUFx10_ASAP7_75t_L g205 ( 
.A(n_33),
.Y(n_205)
);

CKINVDCx5p33_ASAP7_75t_R g206 ( 
.A(n_24),
.Y(n_206)
);

INVx2_ASAP7_75t_SL g207 ( 
.A(n_17),
.Y(n_207)
);

CKINVDCx20_ASAP7_75t_R g208 ( 
.A(n_188),
.Y(n_208)
);

BUFx3_ASAP7_75t_L g209 ( 
.A(n_101),
.Y(n_209)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_1),
.Y(n_210)
);

CKINVDCx20_ASAP7_75t_R g211 ( 
.A(n_42),
.Y(n_211)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_199),
.Y(n_212)
);

CKINVDCx20_ASAP7_75t_R g213 ( 
.A(n_190),
.Y(n_213)
);

HB1xp67_ASAP7_75t_SL g214 ( 
.A(n_69),
.Y(n_214)
);

CKINVDCx5p33_ASAP7_75t_R g215 ( 
.A(n_3),
.Y(n_215)
);

CKINVDCx5p33_ASAP7_75t_R g216 ( 
.A(n_108),
.Y(n_216)
);

CKINVDCx5p33_ASAP7_75t_R g217 ( 
.A(n_44),
.Y(n_217)
);

CKINVDCx5p33_ASAP7_75t_R g218 ( 
.A(n_100),
.Y(n_218)
);

CKINVDCx5p33_ASAP7_75t_R g219 ( 
.A(n_139),
.Y(n_219)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_176),
.Y(n_220)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_192),
.Y(n_221)
);

CKINVDCx5p33_ASAP7_75t_R g222 ( 
.A(n_66),
.Y(n_222)
);

INVx2_ASAP7_75t_L g223 ( 
.A(n_162),
.Y(n_223)
);

CKINVDCx5p33_ASAP7_75t_R g224 ( 
.A(n_62),
.Y(n_224)
);

CKINVDCx5p33_ASAP7_75t_R g225 ( 
.A(n_160),
.Y(n_225)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_186),
.Y(n_226)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_114),
.Y(n_227)
);

BUFx8_ASAP7_75t_SL g228 ( 
.A(n_12),
.Y(n_228)
);

BUFx3_ASAP7_75t_L g229 ( 
.A(n_127),
.Y(n_229)
);

INVx1_ASAP7_75t_SL g230 ( 
.A(n_89),
.Y(n_230)
);

BUFx6f_ASAP7_75t_L g231 ( 
.A(n_61),
.Y(n_231)
);

CKINVDCx5p33_ASAP7_75t_R g232 ( 
.A(n_38),
.Y(n_232)
);

CKINVDCx5p33_ASAP7_75t_R g233 ( 
.A(n_94),
.Y(n_233)
);

BUFx2_ASAP7_75t_L g234 ( 
.A(n_65),
.Y(n_234)
);

CKINVDCx5p33_ASAP7_75t_R g235 ( 
.A(n_83),
.Y(n_235)
);

CKINVDCx5p33_ASAP7_75t_R g236 ( 
.A(n_12),
.Y(n_236)
);

BUFx3_ASAP7_75t_L g237 ( 
.A(n_35),
.Y(n_237)
);

CKINVDCx5p33_ASAP7_75t_R g238 ( 
.A(n_194),
.Y(n_238)
);

BUFx6f_ASAP7_75t_L g239 ( 
.A(n_73),
.Y(n_239)
);

CKINVDCx5p33_ASAP7_75t_R g240 ( 
.A(n_16),
.Y(n_240)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_163),
.Y(n_241)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_0),
.Y(n_242)
);

CKINVDCx20_ASAP7_75t_R g243 ( 
.A(n_130),
.Y(n_243)
);

BUFx10_ASAP7_75t_L g244 ( 
.A(n_178),
.Y(n_244)
);

INVx2_ASAP7_75t_L g245 ( 
.A(n_167),
.Y(n_245)
);

BUFx6f_ASAP7_75t_L g246 ( 
.A(n_147),
.Y(n_246)
);

CKINVDCx20_ASAP7_75t_R g247 ( 
.A(n_43),
.Y(n_247)
);

BUFx10_ASAP7_75t_L g248 ( 
.A(n_136),
.Y(n_248)
);

CKINVDCx5p33_ASAP7_75t_R g249 ( 
.A(n_68),
.Y(n_249)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_189),
.Y(n_250)
);

CKINVDCx5p33_ASAP7_75t_R g251 ( 
.A(n_32),
.Y(n_251)
);

CKINVDCx5p33_ASAP7_75t_R g252 ( 
.A(n_70),
.Y(n_252)
);

CKINVDCx5p33_ASAP7_75t_R g253 ( 
.A(n_150),
.Y(n_253)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_166),
.Y(n_254)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_16),
.Y(n_255)
);

BUFx10_ASAP7_75t_L g256 ( 
.A(n_141),
.Y(n_256)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_78),
.Y(n_257)
);

INVx2_ASAP7_75t_L g258 ( 
.A(n_168),
.Y(n_258)
);

CKINVDCx5p33_ASAP7_75t_R g259 ( 
.A(n_138),
.Y(n_259)
);

CKINVDCx20_ASAP7_75t_R g260 ( 
.A(n_92),
.Y(n_260)
);

CKINVDCx5p33_ASAP7_75t_R g261 ( 
.A(n_87),
.Y(n_261)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_143),
.Y(n_262)
);

BUFx2_ASAP7_75t_L g263 ( 
.A(n_181),
.Y(n_263)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_133),
.Y(n_264)
);

CKINVDCx5p33_ASAP7_75t_R g265 ( 
.A(n_161),
.Y(n_265)
);

CKINVDCx5p33_ASAP7_75t_R g266 ( 
.A(n_151),
.Y(n_266)
);

CKINVDCx20_ASAP7_75t_R g267 ( 
.A(n_228),
.Y(n_267)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_210),
.Y(n_268)
);

INVxp67_ASAP7_75t_L g269 ( 
.A(n_228),
.Y(n_269)
);

INVx2_ASAP7_75t_L g270 ( 
.A(n_242),
.Y(n_270)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_255),
.Y(n_271)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_209),
.Y(n_272)
);

CKINVDCx16_ASAP7_75t_R g273 ( 
.A(n_204),
.Y(n_273)
);

CKINVDCx20_ASAP7_75t_R g274 ( 
.A(n_206),
.Y(n_274)
);

INVxp67_ASAP7_75t_L g275 ( 
.A(n_207),
.Y(n_275)
);

CKINVDCx5p33_ASAP7_75t_R g276 ( 
.A(n_215),
.Y(n_276)
);

HB1xp67_ASAP7_75t_L g277 ( 
.A(n_236),
.Y(n_277)
);

CKINVDCx20_ASAP7_75t_R g278 ( 
.A(n_240),
.Y(n_278)
);

INVxp67_ASAP7_75t_SL g279 ( 
.A(n_234),
.Y(n_279)
);

CKINVDCx5p33_ASAP7_75t_R g280 ( 
.A(n_201),
.Y(n_280)
);

INVx2_ASAP7_75t_L g281 ( 
.A(n_231),
.Y(n_281)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_223),
.Y(n_282)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_223),
.Y(n_283)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_209),
.Y(n_284)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_229),
.Y(n_285)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_229),
.Y(n_286)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_237),
.Y(n_287)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_237),
.Y(n_288)
);

INVx2_ASAP7_75t_L g289 ( 
.A(n_231),
.Y(n_289)
);

CKINVDCx5p33_ASAP7_75t_R g290 ( 
.A(n_216),
.Y(n_290)
);

INVxp67_ASAP7_75t_SL g291 ( 
.A(n_263),
.Y(n_291)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_245),
.Y(n_292)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_202),
.Y(n_293)
);

CKINVDCx20_ASAP7_75t_R g294 ( 
.A(n_208),
.Y(n_294)
);

CKINVDCx16_ASAP7_75t_R g295 ( 
.A(n_204),
.Y(n_295)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_203),
.Y(n_296)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_245),
.Y(n_297)
);

BUFx3_ASAP7_75t_L g298 ( 
.A(n_205),
.Y(n_298)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_212),
.Y(n_299)
);

HB1xp67_ASAP7_75t_L g300 ( 
.A(n_220),
.Y(n_300)
);

CKINVDCx5p33_ASAP7_75t_R g301 ( 
.A(n_217),
.Y(n_301)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_221),
.Y(n_302)
);

BUFx6f_ASAP7_75t_L g303 ( 
.A(n_231),
.Y(n_303)
);

HB1xp67_ASAP7_75t_L g304 ( 
.A(n_226),
.Y(n_304)
);

INVx2_ASAP7_75t_L g305 ( 
.A(n_231),
.Y(n_305)
);

CKINVDCx16_ASAP7_75t_R g306 ( 
.A(n_214),
.Y(n_306)
);

HB1xp67_ASAP7_75t_L g307 ( 
.A(n_227),
.Y(n_307)
);

INVx2_ASAP7_75t_L g308 ( 
.A(n_239),
.Y(n_308)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_258),
.Y(n_309)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_258),
.Y(n_310)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_241),
.Y(n_311)
);

BUFx2_ASAP7_75t_L g312 ( 
.A(n_250),
.Y(n_312)
);

CKINVDCx5p33_ASAP7_75t_R g313 ( 
.A(n_218),
.Y(n_313)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_254),
.Y(n_314)
);

INVxp67_ASAP7_75t_SL g315 ( 
.A(n_257),
.Y(n_315)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_281),
.Y(n_316)
);

INVx3_ASAP7_75t_L g317 ( 
.A(n_303),
.Y(n_317)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_293),
.Y(n_318)
);

BUFx6f_ASAP7_75t_L g319 ( 
.A(n_303),
.Y(n_319)
);

AND2x2_ASAP7_75t_L g320 ( 
.A(n_272),
.B(n_205),
.Y(n_320)
);

OAI22xp5_ASAP7_75t_SL g321 ( 
.A1(n_274),
.A2(n_278),
.B1(n_267),
.B2(n_294),
.Y(n_321)
);

INVx3_ASAP7_75t_L g322 ( 
.A(n_303),
.Y(n_322)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_281),
.Y(n_323)
);

INVx3_ASAP7_75t_L g324 ( 
.A(n_303),
.Y(n_324)
);

NAND2xp5_ASAP7_75t_L g325 ( 
.A(n_280),
.B(n_262),
.Y(n_325)
);

AND2x2_ASAP7_75t_L g326 ( 
.A(n_284),
.B(n_244),
.Y(n_326)
);

INVx4_ASAP7_75t_L g327 ( 
.A(n_303),
.Y(n_327)
);

INVx6_ASAP7_75t_L g328 ( 
.A(n_273),
.Y(n_328)
);

CKINVDCx5p33_ASAP7_75t_R g329 ( 
.A(n_306),
.Y(n_329)
);

INVx3_ASAP7_75t_L g330 ( 
.A(n_289),
.Y(n_330)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_289),
.Y(n_331)
);

NOR2xp33_ASAP7_75t_L g332 ( 
.A(n_280),
.B(n_230),
.Y(n_332)
);

BUFx3_ASAP7_75t_L g333 ( 
.A(n_285),
.Y(n_333)
);

NAND2xp5_ASAP7_75t_L g334 ( 
.A(n_290),
.B(n_264),
.Y(n_334)
);

INVx2_ASAP7_75t_L g335 ( 
.A(n_305),
.Y(n_335)
);

NAND2xp5_ASAP7_75t_L g336 ( 
.A(n_290),
.B(n_219),
.Y(n_336)
);

AND2x4_ASAP7_75t_L g337 ( 
.A(n_315),
.B(n_286),
.Y(n_337)
);

INVx1_ASAP7_75t_L g338 ( 
.A(n_296),
.Y(n_338)
);

BUFx6f_ASAP7_75t_L g339 ( 
.A(n_305),
.Y(n_339)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_308),
.Y(n_340)
);

BUFx6f_ASAP7_75t_L g341 ( 
.A(n_308),
.Y(n_341)
);

BUFx3_ASAP7_75t_L g342 ( 
.A(n_287),
.Y(n_342)
);

INVx1_ASAP7_75t_L g343 ( 
.A(n_270),
.Y(n_343)
);

NAND2xp5_ASAP7_75t_L g344 ( 
.A(n_301),
.B(n_266),
.Y(n_344)
);

INVx1_ASAP7_75t_L g345 ( 
.A(n_299),
.Y(n_345)
);

INVx3_ASAP7_75t_L g346 ( 
.A(n_282),
.Y(n_346)
);

BUFx6f_ASAP7_75t_L g347 ( 
.A(n_282),
.Y(n_347)
);

INVx5_ASAP7_75t_L g348 ( 
.A(n_312),
.Y(n_348)
);

AND2x4_ASAP7_75t_L g349 ( 
.A(n_288),
.B(n_239),
.Y(n_349)
);

INVx2_ASAP7_75t_L g350 ( 
.A(n_283),
.Y(n_350)
);

INVx1_ASAP7_75t_L g351 ( 
.A(n_270),
.Y(n_351)
);

AND2x2_ASAP7_75t_L g352 ( 
.A(n_312),
.B(n_244),
.Y(n_352)
);

INVx2_ASAP7_75t_L g353 ( 
.A(n_283),
.Y(n_353)
);

AOI22xp5_ASAP7_75t_L g354 ( 
.A1(n_279),
.A2(n_243),
.B1(n_213),
.B2(n_260),
.Y(n_354)
);

INVxp67_ASAP7_75t_L g355 ( 
.A(n_277),
.Y(n_355)
);

INVx2_ASAP7_75t_L g356 ( 
.A(n_292),
.Y(n_356)
);

INVx1_ASAP7_75t_L g357 ( 
.A(n_292),
.Y(n_357)
);

AND2x2_ASAP7_75t_SL g358 ( 
.A(n_295),
.B(n_239),
.Y(n_358)
);

INVx1_ASAP7_75t_L g359 ( 
.A(n_297),
.Y(n_359)
);

OAI22xp5_ASAP7_75t_L g360 ( 
.A1(n_291),
.A2(n_211),
.B1(n_247),
.B2(n_259),
.Y(n_360)
);

INVx1_ASAP7_75t_L g361 ( 
.A(n_297),
.Y(n_361)
);

INVx1_ASAP7_75t_L g362 ( 
.A(n_309),
.Y(n_362)
);

INVx1_ASAP7_75t_L g363 ( 
.A(n_309),
.Y(n_363)
);

NAND2xp5_ASAP7_75t_L g364 ( 
.A(n_301),
.B(n_265),
.Y(n_364)
);

INVx2_ASAP7_75t_L g365 ( 
.A(n_310),
.Y(n_365)
);

NAND2xp5_ASAP7_75t_L g366 ( 
.A(n_313),
.B(n_222),
.Y(n_366)
);

INVx1_ASAP7_75t_L g367 ( 
.A(n_302),
.Y(n_367)
);

INVx3_ASAP7_75t_L g368 ( 
.A(n_310),
.Y(n_368)
);

AND2x4_ASAP7_75t_L g369 ( 
.A(n_311),
.B(n_239),
.Y(n_369)
);

NOR2xp33_ASAP7_75t_L g370 ( 
.A(n_332),
.B(n_313),
.Y(n_370)
);

INVx2_ASAP7_75t_L g371 ( 
.A(n_335),
.Y(n_371)
);

INVx1_ASAP7_75t_L g372 ( 
.A(n_335),
.Y(n_372)
);

INVx2_ASAP7_75t_SL g373 ( 
.A(n_348),
.Y(n_373)
);

INVx2_ASAP7_75t_L g374 ( 
.A(n_316),
.Y(n_374)
);

BUFx3_ASAP7_75t_L g375 ( 
.A(n_333),
.Y(n_375)
);

AND2x2_ASAP7_75t_L g376 ( 
.A(n_337),
.B(n_300),
.Y(n_376)
);

NAND2xp33_ASAP7_75t_L g377 ( 
.A(n_325),
.B(n_276),
.Y(n_377)
);

NAND2xp5_ASAP7_75t_L g378 ( 
.A(n_337),
.B(n_314),
.Y(n_378)
);

INVx3_ASAP7_75t_L g379 ( 
.A(n_319),
.Y(n_379)
);

NAND2xp33_ASAP7_75t_L g380 ( 
.A(n_334),
.B(n_276),
.Y(n_380)
);

INVx2_ASAP7_75t_L g381 ( 
.A(n_316),
.Y(n_381)
);

NOR2xp33_ASAP7_75t_L g382 ( 
.A(n_336),
.B(n_298),
.Y(n_382)
);

INVx1_ASAP7_75t_L g383 ( 
.A(n_318),
.Y(n_383)
);

CKINVDCx5p33_ASAP7_75t_R g384 ( 
.A(n_329),
.Y(n_384)
);

INVx2_ASAP7_75t_L g385 ( 
.A(n_323),
.Y(n_385)
);

INVx2_ASAP7_75t_L g386 ( 
.A(n_323),
.Y(n_386)
);

HB1xp67_ASAP7_75t_L g387 ( 
.A(n_348),
.Y(n_387)
);

INVx11_ASAP7_75t_L g388 ( 
.A(n_328),
.Y(n_388)
);

INVx2_ASAP7_75t_L g389 ( 
.A(n_331),
.Y(n_389)
);

AND2x2_ASAP7_75t_L g390 ( 
.A(n_348),
.B(n_304),
.Y(n_390)
);

NOR2x1p5_ASAP7_75t_L g391 ( 
.A(n_329),
.B(n_298),
.Y(n_391)
);

INVx1_ASAP7_75t_L g392 ( 
.A(n_338),
.Y(n_392)
);

AND2x2_ASAP7_75t_L g393 ( 
.A(n_348),
.B(n_307),
.Y(n_393)
);

INVx2_ASAP7_75t_L g394 ( 
.A(n_331),
.Y(n_394)
);

NAND2xp5_ASAP7_75t_SL g395 ( 
.A(n_358),
.B(n_269),
.Y(n_395)
);

INVxp33_ASAP7_75t_L g396 ( 
.A(n_321),
.Y(n_396)
);

HB1xp67_ASAP7_75t_L g397 ( 
.A(n_348),
.Y(n_397)
);

XNOR2xp5_ASAP7_75t_L g398 ( 
.A(n_354),
.B(n_294),
.Y(n_398)
);

AND2x2_ASAP7_75t_L g399 ( 
.A(n_349),
.B(n_268),
.Y(n_399)
);

INVx2_ASAP7_75t_L g400 ( 
.A(n_340),
.Y(n_400)
);

INVx1_ASAP7_75t_L g401 ( 
.A(n_345),
.Y(n_401)
);

INVx2_ASAP7_75t_L g402 ( 
.A(n_340),
.Y(n_402)
);

NAND2xp5_ASAP7_75t_SL g403 ( 
.A(n_358),
.B(n_352),
.Y(n_403)
);

INVx2_ASAP7_75t_L g404 ( 
.A(n_347),
.Y(n_404)
);

INVx2_ASAP7_75t_L g405 ( 
.A(n_347),
.Y(n_405)
);

INVx2_ASAP7_75t_L g406 ( 
.A(n_347),
.Y(n_406)
);

INVx2_ASAP7_75t_L g407 ( 
.A(n_347),
.Y(n_407)
);

NAND2xp5_ASAP7_75t_L g408 ( 
.A(n_344),
.B(n_224),
.Y(n_408)
);

INVx2_ASAP7_75t_L g409 ( 
.A(n_347),
.Y(n_409)
);

INVx1_ASAP7_75t_L g410 ( 
.A(n_367),
.Y(n_410)
);

NAND3x1_ASAP7_75t_L g411 ( 
.A(n_352),
.B(n_271),
.C(n_256),
.Y(n_411)
);

INVx2_ASAP7_75t_L g412 ( 
.A(n_339),
.Y(n_412)
);

INVx2_ASAP7_75t_SL g413 ( 
.A(n_320),
.Y(n_413)
);

INVx6_ASAP7_75t_L g414 ( 
.A(n_327),
.Y(n_414)
);

INVx2_ASAP7_75t_L g415 ( 
.A(n_339),
.Y(n_415)
);

INVx1_ASAP7_75t_L g416 ( 
.A(n_357),
.Y(n_416)
);

NOR2xp33_ASAP7_75t_L g417 ( 
.A(n_364),
.B(n_366),
.Y(n_417)
);

INVx1_ASAP7_75t_L g418 ( 
.A(n_357),
.Y(n_418)
);

OR2x2_ASAP7_75t_L g419 ( 
.A(n_360),
.B(n_320),
.Y(n_419)
);

INVx1_ASAP7_75t_L g420 ( 
.A(n_359),
.Y(n_420)
);

INVx1_ASAP7_75t_L g421 ( 
.A(n_359),
.Y(n_421)
);

AO21x2_ASAP7_75t_L g422 ( 
.A1(n_369),
.A2(n_275),
.B(n_246),
.Y(n_422)
);

INVx2_ASAP7_75t_L g423 ( 
.A(n_339),
.Y(n_423)
);

BUFx6f_ASAP7_75t_SL g424 ( 
.A(n_349),
.Y(n_424)
);

INVx2_ASAP7_75t_L g425 ( 
.A(n_339),
.Y(n_425)
);

INVx4_ASAP7_75t_L g426 ( 
.A(n_319),
.Y(n_426)
);

INVx1_ASAP7_75t_L g427 ( 
.A(n_361),
.Y(n_427)
);

INVx2_ASAP7_75t_L g428 ( 
.A(n_330),
.Y(n_428)
);

INVx1_ASAP7_75t_L g429 ( 
.A(n_361),
.Y(n_429)
);

NAND2xp5_ASAP7_75t_SL g430 ( 
.A(n_355),
.B(n_326),
.Y(n_430)
);

INVxp33_ASAP7_75t_L g431 ( 
.A(n_326),
.Y(n_431)
);

NOR2x1p5_ASAP7_75t_L g432 ( 
.A(n_333),
.B(n_225),
.Y(n_432)
);

INVx2_ASAP7_75t_L g433 ( 
.A(n_339),
.Y(n_433)
);

INVx1_ASAP7_75t_L g434 ( 
.A(n_362),
.Y(n_434)
);

INVx2_ASAP7_75t_L g435 ( 
.A(n_341),
.Y(n_435)
);

INVx2_ASAP7_75t_L g436 ( 
.A(n_341),
.Y(n_436)
);

BUFx3_ASAP7_75t_L g437 ( 
.A(n_342),
.Y(n_437)
);

INVx2_ASAP7_75t_L g438 ( 
.A(n_341),
.Y(n_438)
);

INVx3_ASAP7_75t_L g439 ( 
.A(n_319),
.Y(n_439)
);

NAND2xp33_ASAP7_75t_L g440 ( 
.A(n_341),
.B(n_246),
.Y(n_440)
);

NAND2xp5_ASAP7_75t_L g441 ( 
.A(n_369),
.B(n_317),
.Y(n_441)
);

NOR2xp33_ASAP7_75t_SL g442 ( 
.A(n_370),
.B(n_248),
.Y(n_442)
);

INVx1_ASAP7_75t_L g443 ( 
.A(n_383),
.Y(n_443)
);

INVx1_ASAP7_75t_L g444 ( 
.A(n_383),
.Y(n_444)
);

XOR2xp5_ASAP7_75t_L g445 ( 
.A(n_398),
.B(n_384),
.Y(n_445)
);

INVx1_ASAP7_75t_L g446 ( 
.A(n_392),
.Y(n_446)
);

NAND2xp5_ASAP7_75t_L g447 ( 
.A(n_417),
.B(n_346),
.Y(n_447)
);

NAND2xp33_ASAP7_75t_SL g448 ( 
.A(n_403),
.B(n_274),
.Y(n_448)
);

INVx1_ASAP7_75t_L g449 ( 
.A(n_392),
.Y(n_449)
);

INVxp67_ASAP7_75t_L g450 ( 
.A(n_376),
.Y(n_450)
);

CKINVDCx20_ASAP7_75t_R g451 ( 
.A(n_395),
.Y(n_451)
);

INVx1_ASAP7_75t_L g452 ( 
.A(n_401),
.Y(n_452)
);

INVxp67_ASAP7_75t_SL g453 ( 
.A(n_416),
.Y(n_453)
);

INVx1_ASAP7_75t_L g454 ( 
.A(n_401),
.Y(n_454)
);

INVx1_ASAP7_75t_L g455 ( 
.A(n_410),
.Y(n_455)
);

INVx1_ASAP7_75t_L g456 ( 
.A(n_410),
.Y(n_456)
);

AND2x4_ASAP7_75t_L g457 ( 
.A(n_375),
.B(n_342),
.Y(n_457)
);

AND2x2_ASAP7_75t_L g458 ( 
.A(n_431),
.B(n_328),
.Y(n_458)
);

XNOR2xp5_ASAP7_75t_L g459 ( 
.A(n_391),
.B(n_267),
.Y(n_459)
);

INVx1_ASAP7_75t_L g460 ( 
.A(n_416),
.Y(n_460)
);

CKINVDCx20_ASAP7_75t_R g461 ( 
.A(n_375),
.Y(n_461)
);

INVx1_ASAP7_75t_L g462 ( 
.A(n_418),
.Y(n_462)
);

BUFx3_ASAP7_75t_L g463 ( 
.A(n_375),
.Y(n_463)
);

INVx1_ASAP7_75t_L g464 ( 
.A(n_418),
.Y(n_464)
);

INVx2_ASAP7_75t_SL g465 ( 
.A(n_376),
.Y(n_465)
);

INVx1_ASAP7_75t_L g466 ( 
.A(n_420),
.Y(n_466)
);

INVx1_ASAP7_75t_L g467 ( 
.A(n_420),
.Y(n_467)
);

AND2x2_ASAP7_75t_L g468 ( 
.A(n_413),
.B(n_328),
.Y(n_468)
);

INVx1_ASAP7_75t_L g469 ( 
.A(n_421),
.Y(n_469)
);

XNOR2xp5_ASAP7_75t_L g470 ( 
.A(n_391),
.B(n_411),
.Y(n_470)
);

INVx1_ASAP7_75t_L g471 ( 
.A(n_427),
.Y(n_471)
);

NOR2xp67_ASAP7_75t_L g472 ( 
.A(n_413),
.B(n_346),
.Y(n_472)
);

INVx2_ASAP7_75t_L g473 ( 
.A(n_428),
.Y(n_473)
);

INVx1_ASAP7_75t_L g474 ( 
.A(n_429),
.Y(n_474)
);

NAND2xp33_ASAP7_75t_SL g475 ( 
.A(n_419),
.B(n_278),
.Y(n_475)
);

INVx1_ASAP7_75t_L g476 ( 
.A(n_434),
.Y(n_476)
);

INVx2_ASAP7_75t_L g477 ( 
.A(n_428),
.Y(n_477)
);

INVx1_ASAP7_75t_L g478 ( 
.A(n_434),
.Y(n_478)
);

INVx1_ASAP7_75t_L g479 ( 
.A(n_441),
.Y(n_479)
);

INVx4_ASAP7_75t_SL g480 ( 
.A(n_424),
.Y(n_480)
);

XOR2xp5_ASAP7_75t_L g481 ( 
.A(n_396),
.B(n_232),
.Y(n_481)
);

INVx1_ASAP7_75t_L g482 ( 
.A(n_374),
.Y(n_482)
);

INVx1_ASAP7_75t_L g483 ( 
.A(n_381),
.Y(n_483)
);

XOR2xp5_ASAP7_75t_L g484 ( 
.A(n_419),
.B(n_233),
.Y(n_484)
);

INVx1_ASAP7_75t_L g485 ( 
.A(n_381),
.Y(n_485)
);

INVx1_ASAP7_75t_L g486 ( 
.A(n_400),
.Y(n_486)
);

AND2x2_ASAP7_75t_L g487 ( 
.A(n_390),
.B(n_328),
.Y(n_487)
);

INVx1_ASAP7_75t_L g488 ( 
.A(n_400),
.Y(n_488)
);

INVx1_ASAP7_75t_L g489 ( 
.A(n_402),
.Y(n_489)
);

INVx1_ASAP7_75t_L g490 ( 
.A(n_402),
.Y(n_490)
);

INVx1_ASAP7_75t_L g491 ( 
.A(n_399),
.Y(n_491)
);

CKINVDCx20_ASAP7_75t_R g492 ( 
.A(n_437),
.Y(n_492)
);

AND2x2_ASAP7_75t_L g493 ( 
.A(n_393),
.B(n_382),
.Y(n_493)
);

XOR2xp5_ASAP7_75t_L g494 ( 
.A(n_408),
.B(n_235),
.Y(n_494)
);

INVx1_ASAP7_75t_L g495 ( 
.A(n_399),
.Y(n_495)
);

AND2x2_ASAP7_75t_L g496 ( 
.A(n_393),
.B(n_343),
.Y(n_496)
);

INVx2_ASAP7_75t_L g497 ( 
.A(n_371),
.Y(n_497)
);

CKINVDCx16_ASAP7_75t_R g498 ( 
.A(n_424),
.Y(n_498)
);

AND2x4_ASAP7_75t_L g499 ( 
.A(n_437),
.B(n_362),
.Y(n_499)
);

NOR2xp33_ASAP7_75t_L g500 ( 
.A(n_430),
.B(n_369),
.Y(n_500)
);

INVx1_ASAP7_75t_SL g501 ( 
.A(n_437),
.Y(n_501)
);

NOR2xp33_ASAP7_75t_L g502 ( 
.A(n_378),
.B(n_238),
.Y(n_502)
);

NAND2xp5_ASAP7_75t_L g503 ( 
.A(n_422),
.B(n_368),
.Y(n_503)
);

INVx2_ASAP7_75t_SL g504 ( 
.A(n_432),
.Y(n_504)
);

INVx1_ASAP7_75t_L g505 ( 
.A(n_385),
.Y(n_505)
);

NOR2xp33_ASAP7_75t_L g506 ( 
.A(n_377),
.B(n_380),
.Y(n_506)
);

BUFx6f_ASAP7_75t_L g507 ( 
.A(n_405),
.Y(n_507)
);

XOR2xp5_ASAP7_75t_L g508 ( 
.A(n_387),
.B(n_249),
.Y(n_508)
);

INVx1_ASAP7_75t_L g509 ( 
.A(n_385),
.Y(n_509)
);

INVx1_ASAP7_75t_L g510 ( 
.A(n_385),
.Y(n_510)
);

NOR2xp33_ASAP7_75t_L g511 ( 
.A(n_397),
.B(n_251),
.Y(n_511)
);

INVx2_ASAP7_75t_L g512 ( 
.A(n_371),
.Y(n_512)
);

INVx2_ASAP7_75t_L g513 ( 
.A(n_386),
.Y(n_513)
);

INVx1_ASAP7_75t_L g514 ( 
.A(n_386),
.Y(n_514)
);

INVx1_ASAP7_75t_L g515 ( 
.A(n_386),
.Y(n_515)
);

OR2x2_ASAP7_75t_L g516 ( 
.A(n_432),
.B(n_363),
.Y(n_516)
);

BUFx2_ASAP7_75t_L g517 ( 
.A(n_461),
.Y(n_517)
);

NAND2xp5_ASAP7_75t_SL g518 ( 
.A(n_493),
.B(n_373),
.Y(n_518)
);

NAND3xp33_ASAP7_75t_SL g519 ( 
.A(n_442),
.B(n_253),
.C(n_252),
.Y(n_519)
);

AOI22xp5_ASAP7_75t_L g520 ( 
.A1(n_506),
.A2(n_424),
.B1(n_373),
.B2(n_411),
.Y(n_520)
);

INVx2_ASAP7_75t_L g521 ( 
.A(n_497),
.Y(n_521)
);

NAND2xp5_ASAP7_75t_L g522 ( 
.A(n_447),
.B(n_453),
.Y(n_522)
);

AOI22xp33_ASAP7_75t_L g523 ( 
.A1(n_479),
.A2(n_422),
.B1(n_394),
.B2(n_389),
.Y(n_523)
);

AND2x2_ASAP7_75t_L g524 ( 
.A(n_450),
.B(n_422),
.Y(n_524)
);

NAND2xp5_ASAP7_75t_L g525 ( 
.A(n_447),
.B(n_404),
.Y(n_525)
);

NOR2x2_ASAP7_75t_L g526 ( 
.A(n_484),
.B(n_388),
.Y(n_526)
);

NAND2xp5_ASAP7_75t_SL g527 ( 
.A(n_501),
.B(n_406),
.Y(n_527)
);

AOI22xp33_ASAP7_75t_L g528 ( 
.A1(n_491),
.A2(n_407),
.B1(n_409),
.B2(n_406),
.Y(n_528)
);

NAND2xp5_ASAP7_75t_SL g529 ( 
.A(n_501),
.B(n_409),
.Y(n_529)
);

INVx2_ASAP7_75t_SL g530 ( 
.A(n_465),
.Y(n_530)
);

NAND2xp5_ASAP7_75t_SL g531 ( 
.A(n_506),
.B(n_405),
.Y(n_531)
);

AND2x2_ASAP7_75t_SL g532 ( 
.A(n_503),
.B(n_246),
.Y(n_532)
);

AND2x4_ASAP7_75t_L g533 ( 
.A(n_463),
.B(n_405),
.Y(n_533)
);

AOI22xp5_ASAP7_75t_L g534 ( 
.A1(n_448),
.A2(n_414),
.B1(n_415),
.B2(n_412),
.Y(n_534)
);

AND2x2_ASAP7_75t_L g535 ( 
.A(n_468),
.B(n_351),
.Y(n_535)
);

A2O1A1Ixp33_ASAP7_75t_L g536 ( 
.A1(n_500),
.A2(n_394),
.B(n_389),
.C(n_412),
.Y(n_536)
);

AND2x4_ASAP7_75t_L g537 ( 
.A(n_480),
.B(n_457),
.Y(n_537)
);

NAND2xp5_ASAP7_75t_L g538 ( 
.A(n_496),
.B(n_379),
.Y(n_538)
);

NAND2xp5_ASAP7_75t_L g539 ( 
.A(n_460),
.B(n_379),
.Y(n_539)
);

INVx1_ASAP7_75t_L g540 ( 
.A(n_482),
.Y(n_540)
);

AOI22xp33_ASAP7_75t_L g541 ( 
.A1(n_462),
.A2(n_394),
.B1(n_389),
.B2(n_372),
.Y(n_541)
);

AOI22xp33_ASAP7_75t_L g542 ( 
.A1(n_464),
.A2(n_466),
.B1(n_469),
.B2(n_467),
.Y(n_542)
);

NAND2xp5_ASAP7_75t_SL g543 ( 
.A(n_487),
.B(n_261),
.Y(n_543)
);

NOR2xp33_ASAP7_75t_L g544 ( 
.A(n_494),
.B(n_414),
.Y(n_544)
);

O2A1O1Ixp33_ASAP7_75t_L g545 ( 
.A1(n_495),
.A2(n_372),
.B(n_440),
.C(n_368),
.Y(n_545)
);

AND2x6_ASAP7_75t_L g546 ( 
.A(n_503),
.B(n_415),
.Y(n_546)
);

INVx2_ASAP7_75t_L g547 ( 
.A(n_512),
.Y(n_547)
);

INVxp67_ASAP7_75t_L g548 ( 
.A(n_500),
.Y(n_548)
);

INVx2_ASAP7_75t_SL g549 ( 
.A(n_458),
.Y(n_549)
);

NAND2xp5_ASAP7_75t_L g550 ( 
.A(n_471),
.B(n_379),
.Y(n_550)
);

INVx1_ASAP7_75t_L g551 ( 
.A(n_483),
.Y(n_551)
);

NAND2xp5_ASAP7_75t_L g552 ( 
.A(n_474),
.B(n_379),
.Y(n_552)
);

NAND2xp5_ASAP7_75t_SL g553 ( 
.A(n_472),
.B(n_248),
.Y(n_553)
);

INVx2_ASAP7_75t_SL g554 ( 
.A(n_516),
.Y(n_554)
);

NOR3xp33_ASAP7_75t_L g555 ( 
.A(n_475),
.B(n_351),
.C(n_368),
.Y(n_555)
);

AOI22xp5_ASAP7_75t_L g556 ( 
.A1(n_448),
.A2(n_414),
.B1(n_438),
.B2(n_436),
.Y(n_556)
);

NAND2xp5_ASAP7_75t_SL g557 ( 
.A(n_457),
.B(n_256),
.Y(n_557)
);

NAND2xp5_ASAP7_75t_L g558 ( 
.A(n_476),
.B(n_439),
.Y(n_558)
);

INVx2_ASAP7_75t_L g559 ( 
.A(n_513),
.Y(n_559)
);

NAND2xp5_ASAP7_75t_L g560 ( 
.A(n_478),
.B(n_439),
.Y(n_560)
);

NAND2xp5_ASAP7_75t_L g561 ( 
.A(n_443),
.B(n_439),
.Y(n_561)
);

NAND2xp5_ASAP7_75t_L g562 ( 
.A(n_444),
.B(n_439),
.Y(n_562)
);

AOI22xp33_ASAP7_75t_L g563 ( 
.A1(n_446),
.A2(n_246),
.B1(n_436),
.B2(n_435),
.Y(n_563)
);

INVx1_ASAP7_75t_L g564 ( 
.A(n_485),
.Y(n_564)
);

NAND2xp5_ASAP7_75t_SL g565 ( 
.A(n_499),
.B(n_423),
.Y(n_565)
);

INVx2_ASAP7_75t_L g566 ( 
.A(n_486),
.Y(n_566)
);

HB1xp67_ASAP7_75t_L g567 ( 
.A(n_499),
.Y(n_567)
);

NAND2xp5_ASAP7_75t_L g568 ( 
.A(n_449),
.B(n_423),
.Y(n_568)
);

NOR3xp33_ASAP7_75t_L g569 ( 
.A(n_498),
.B(n_353),
.C(n_350),
.Y(n_569)
);

NOR2xp33_ASAP7_75t_L g570 ( 
.A(n_481),
.B(n_426),
.Y(n_570)
);

OAI22xp33_ASAP7_75t_SL g571 ( 
.A1(n_504),
.A2(n_350),
.B1(n_353),
.B2(n_356),
.Y(n_571)
);

NAND2xp5_ASAP7_75t_SL g572 ( 
.A(n_502),
.B(n_425),
.Y(n_572)
);

AND2x2_ASAP7_75t_L g573 ( 
.A(n_452),
.B(n_356),
.Y(n_573)
);

NOR2xp33_ASAP7_75t_L g574 ( 
.A(n_451),
.B(n_426),
.Y(n_574)
);

INVx1_ASAP7_75t_L g575 ( 
.A(n_488),
.Y(n_575)
);

NOR3xp33_ASAP7_75t_SL g576 ( 
.A(n_519),
.B(n_470),
.C(n_459),
.Y(n_576)
);

NOR2xp33_ASAP7_75t_R g577 ( 
.A(n_519),
.B(n_492),
.Y(n_577)
);

BUFx3_ASAP7_75t_L g578 ( 
.A(n_517),
.Y(n_578)
);

AND2x4_ASAP7_75t_L g579 ( 
.A(n_537),
.B(n_549),
.Y(n_579)
);

NAND2xp5_ASAP7_75t_L g580 ( 
.A(n_522),
.B(n_548),
.Y(n_580)
);

INVx2_ASAP7_75t_L g581 ( 
.A(n_559),
.Y(n_581)
);

CKINVDCx5p33_ASAP7_75t_R g582 ( 
.A(n_544),
.Y(n_582)
);

INVx2_ASAP7_75t_L g583 ( 
.A(n_566),
.Y(n_583)
);

NAND2xp5_ASAP7_75t_L g584 ( 
.A(n_535),
.B(n_454),
.Y(n_584)
);

INVx1_ASAP7_75t_L g585 ( 
.A(n_573),
.Y(n_585)
);

NOR2xp33_ASAP7_75t_L g586 ( 
.A(n_574),
.B(n_445),
.Y(n_586)
);

BUFx6f_ASAP7_75t_L g587 ( 
.A(n_537),
.Y(n_587)
);

BUFx2_ASAP7_75t_L g588 ( 
.A(n_554),
.Y(n_588)
);

BUFx6f_ASAP7_75t_L g589 ( 
.A(n_533),
.Y(n_589)
);

OR2x6_ASAP7_75t_L g590 ( 
.A(n_530),
.B(n_455),
.Y(n_590)
);

AND2x6_ASAP7_75t_L g591 ( 
.A(n_524),
.B(n_456),
.Y(n_591)
);

INVx5_ASAP7_75t_L g592 ( 
.A(n_546),
.Y(n_592)
);

NOR2xp33_ASAP7_75t_R g593 ( 
.A(n_570),
.B(n_511),
.Y(n_593)
);

BUFx6f_ASAP7_75t_L g594 ( 
.A(n_533),
.Y(n_594)
);

HB1xp67_ASAP7_75t_L g595 ( 
.A(n_567),
.Y(n_595)
);

NAND3xp33_ASAP7_75t_SL g596 ( 
.A(n_569),
.B(n_508),
.C(n_511),
.Y(n_596)
);

CKINVDCx5p33_ASAP7_75t_R g597 ( 
.A(n_520),
.Y(n_597)
);

INVx1_ASAP7_75t_L g598 ( 
.A(n_540),
.Y(n_598)
);

INVx1_ASAP7_75t_L g599 ( 
.A(n_551),
.Y(n_599)
);

AOI22xp33_ASAP7_75t_L g600 ( 
.A1(n_555),
.A2(n_532),
.B1(n_569),
.B2(n_567),
.Y(n_600)
);

INVx2_ASAP7_75t_SL g601 ( 
.A(n_557),
.Y(n_601)
);

INVx1_ASAP7_75t_L g602 ( 
.A(n_564),
.Y(n_602)
);

INVx1_ASAP7_75t_SL g603 ( 
.A(n_543),
.Y(n_603)
);

BUFx4f_ASAP7_75t_L g604 ( 
.A(n_575),
.Y(n_604)
);

INVx1_ASAP7_75t_L g605 ( 
.A(n_568),
.Y(n_605)
);

AND2x4_ASAP7_75t_L g606 ( 
.A(n_555),
.B(n_480),
.Y(n_606)
);

INVx3_ASAP7_75t_L g607 ( 
.A(n_521),
.Y(n_607)
);

CKINVDCx14_ASAP7_75t_R g608 ( 
.A(n_526),
.Y(n_608)
);

NAND2xp5_ASAP7_75t_L g609 ( 
.A(n_542),
.B(n_489),
.Y(n_609)
);

HB1xp67_ASAP7_75t_L g610 ( 
.A(n_547),
.Y(n_610)
);

OR2x4_ASAP7_75t_L g611 ( 
.A(n_553),
.B(n_507),
.Y(n_611)
);

BUFx6f_ASAP7_75t_L g612 ( 
.A(n_527),
.Y(n_612)
);

INVx2_ASAP7_75t_L g613 ( 
.A(n_539),
.Y(n_613)
);

NAND2xp5_ASAP7_75t_SL g614 ( 
.A(n_542),
.B(n_507),
.Y(n_614)
);

INVx1_ASAP7_75t_L g615 ( 
.A(n_561),
.Y(n_615)
);

INVx2_ASAP7_75t_L g616 ( 
.A(n_550),
.Y(n_616)
);

OAI22xp33_ASAP7_75t_L g617 ( 
.A1(n_538),
.A2(n_490),
.B1(n_514),
.B2(n_510),
.Y(n_617)
);

INVx1_ASAP7_75t_L g618 ( 
.A(n_562),
.Y(n_618)
);

AND2x4_ASAP7_75t_L g619 ( 
.A(n_565),
.B(n_505),
.Y(n_619)
);

NAND2xp5_ASAP7_75t_L g620 ( 
.A(n_525),
.B(n_509),
.Y(n_620)
);

BUFx2_ASAP7_75t_L g621 ( 
.A(n_546),
.Y(n_621)
);

NAND2xp5_ASAP7_75t_L g622 ( 
.A(n_532),
.B(n_515),
.Y(n_622)
);

BUFx2_ASAP7_75t_L g623 ( 
.A(n_546),
.Y(n_623)
);

CKINVDCx6p67_ASAP7_75t_R g624 ( 
.A(n_546),
.Y(n_624)
);

CKINVDCx20_ASAP7_75t_R g625 ( 
.A(n_518),
.Y(n_625)
);

INVx1_ASAP7_75t_L g626 ( 
.A(n_552),
.Y(n_626)
);

NAND2xp5_ASAP7_75t_SL g627 ( 
.A(n_571),
.B(n_473),
.Y(n_627)
);

AO31x2_ASAP7_75t_L g628 ( 
.A1(n_621),
.A2(n_536),
.A3(n_560),
.B(n_558),
.Y(n_628)
);

NAND2xp5_ASAP7_75t_L g629 ( 
.A(n_580),
.B(n_546),
.Y(n_629)
);

OA21x2_ASAP7_75t_L g630 ( 
.A1(n_622),
.A2(n_523),
.B(n_531),
.Y(n_630)
);

NAND2xp5_ASAP7_75t_L g631 ( 
.A(n_585),
.B(n_529),
.Y(n_631)
);

AND2x4_ASAP7_75t_L g632 ( 
.A(n_587),
.B(n_579),
.Y(n_632)
);

AOI21xp5_ASAP7_75t_L g633 ( 
.A1(n_620),
.A2(n_572),
.B(n_523),
.Y(n_633)
);

OAI21x1_ASAP7_75t_L g634 ( 
.A1(n_627),
.A2(n_541),
.B(n_545),
.Y(n_634)
);

INVx3_ASAP7_75t_L g635 ( 
.A(n_587),
.Y(n_635)
);

NAND2xp5_ASAP7_75t_L g636 ( 
.A(n_584),
.B(n_541),
.Y(n_636)
);

AND2x2_ASAP7_75t_L g637 ( 
.A(n_593),
.B(n_528),
.Y(n_637)
);

OA22x2_ASAP7_75t_L g638 ( 
.A1(n_597),
.A2(n_534),
.B1(n_556),
.B2(n_477),
.Y(n_638)
);

O2A1O1Ixp33_ASAP7_75t_L g639 ( 
.A1(n_596),
.A2(n_365),
.B(n_438),
.C(n_435),
.Y(n_639)
);

BUFx3_ASAP7_75t_L g640 ( 
.A(n_578),
.Y(n_640)
);

OAI21xp5_ASAP7_75t_L g641 ( 
.A1(n_622),
.A2(n_563),
.B(n_433),
.Y(n_641)
);

AOI21xp5_ASAP7_75t_L g642 ( 
.A1(n_614),
.A2(n_426),
.B(n_327),
.Y(n_642)
);

INVx1_ASAP7_75t_L g643 ( 
.A(n_598),
.Y(n_643)
);

INVx4_ASAP7_75t_L g644 ( 
.A(n_587),
.Y(n_644)
);

AOI21xp5_ASAP7_75t_L g645 ( 
.A1(n_617),
.A2(n_327),
.B(n_319),
.Y(n_645)
);

BUFx3_ASAP7_75t_L g646 ( 
.A(n_588),
.Y(n_646)
);

INVx2_ASAP7_75t_L g647 ( 
.A(n_599),
.Y(n_647)
);

NAND2xp5_ASAP7_75t_L g648 ( 
.A(n_605),
.B(n_330),
.Y(n_648)
);

BUFx5_ASAP7_75t_L g649 ( 
.A(n_591),
.Y(n_649)
);

INVx2_ASAP7_75t_L g650 ( 
.A(n_602),
.Y(n_650)
);

INVx1_ASAP7_75t_L g651 ( 
.A(n_610),
.Y(n_651)
);

OAI21x1_ASAP7_75t_L g652 ( 
.A1(n_609),
.A2(n_322),
.B(n_317),
.Y(n_652)
);

NAND2xp5_ASAP7_75t_L g653 ( 
.A(n_626),
.B(n_330),
.Y(n_653)
);

OAI21xp5_ASAP7_75t_L g654 ( 
.A1(n_615),
.A2(n_618),
.B(n_600),
.Y(n_654)
);

OAI21xp5_ASAP7_75t_L g655 ( 
.A1(n_613),
.A2(n_322),
.B(n_317),
.Y(n_655)
);

OAI22xp5_ASAP7_75t_L g656 ( 
.A1(n_604),
.A2(n_603),
.B1(n_589),
.B2(n_594),
.Y(n_656)
);

NAND2xp5_ASAP7_75t_L g657 ( 
.A(n_616),
.B(n_0),
.Y(n_657)
);

NAND2xp5_ASAP7_75t_L g658 ( 
.A(n_603),
.B(n_1),
.Y(n_658)
);

A2O1A1Ixp33_ASAP7_75t_L g659 ( 
.A1(n_604),
.A2(n_324),
.B(n_341),
.C(n_319),
.Y(n_659)
);

OAI21xp5_ASAP7_75t_L g660 ( 
.A1(n_619),
.A2(n_324),
.B(n_31),
.Y(n_660)
);

BUFx6f_ASAP7_75t_L g661 ( 
.A(n_589),
.Y(n_661)
);

BUFx2_ASAP7_75t_L g662 ( 
.A(n_625),
.Y(n_662)
);

NAND2xp5_ASAP7_75t_L g663 ( 
.A(n_583),
.B(n_2),
.Y(n_663)
);

NOR2x1_ASAP7_75t_L g664 ( 
.A(n_590),
.B(n_324),
.Y(n_664)
);

AO31x2_ASAP7_75t_L g665 ( 
.A1(n_623),
.A2(n_2),
.A3(n_3),
.B(n_4),
.Y(n_665)
);

AOI21x1_ASAP7_75t_L g666 ( 
.A1(n_606),
.A2(n_36),
.B(n_34),
.Y(n_666)
);

NAND2xp5_ASAP7_75t_L g667 ( 
.A(n_589),
.B(n_4),
.Y(n_667)
);

AO31x2_ASAP7_75t_L g668 ( 
.A1(n_581),
.A2(n_5),
.A3(n_6),
.B(n_7),
.Y(n_668)
);

AND2x2_ASAP7_75t_L g669 ( 
.A(n_595),
.B(n_5),
.Y(n_669)
);

NAND2xp5_ASAP7_75t_L g670 ( 
.A(n_594),
.B(n_6),
.Y(n_670)
);

BUFx10_ASAP7_75t_L g671 ( 
.A(n_579),
.Y(n_671)
);

NAND2x1_ASAP7_75t_L g672 ( 
.A(n_591),
.B(n_37),
.Y(n_672)
);

A2O1A1Ixp33_ASAP7_75t_L g673 ( 
.A1(n_601),
.A2(n_8),
.B(n_9),
.C(n_10),
.Y(n_673)
);

OAI21x1_ASAP7_75t_L g674 ( 
.A1(n_607),
.A2(n_40),
.B(n_39),
.Y(n_674)
);

NOR2xp33_ASAP7_75t_L g675 ( 
.A(n_586),
.B(n_10),
.Y(n_675)
);

AOI21xp33_ASAP7_75t_L g676 ( 
.A1(n_582),
.A2(n_590),
.B(n_612),
.Y(n_676)
);

NAND2xp5_ASAP7_75t_L g677 ( 
.A(n_607),
.B(n_11),
.Y(n_677)
);

OAI21x1_ASAP7_75t_L g678 ( 
.A1(n_624),
.A2(n_45),
.B(n_41),
.Y(n_678)
);

AOI21xp5_ASAP7_75t_L g679 ( 
.A1(n_592),
.A2(n_47),
.B(n_46),
.Y(n_679)
);

NAND2x1p5_ASAP7_75t_L g680 ( 
.A(n_592),
.B(n_48),
.Y(n_680)
);

OA21x2_ASAP7_75t_L g681 ( 
.A1(n_619),
.A2(n_50),
.B(n_49),
.Y(n_681)
);

BUFx6f_ASAP7_75t_L g682 ( 
.A(n_590),
.Y(n_682)
);

OA21x2_ASAP7_75t_L g683 ( 
.A1(n_652),
.A2(n_606),
.B(n_592),
.Y(n_683)
);

CKINVDCx5p33_ASAP7_75t_R g684 ( 
.A(n_640),
.Y(n_684)
);

O2A1O1Ixp33_ASAP7_75t_SL g685 ( 
.A1(n_660),
.A2(n_611),
.B(n_576),
.C(n_591),
.Y(n_685)
);

NAND2xp5_ASAP7_75t_SL g686 ( 
.A(n_637),
.B(n_577),
.Y(n_686)
);

INVx1_ASAP7_75t_L g687 ( 
.A(n_647),
.Y(n_687)
);

NOR2xp33_ASAP7_75t_L g688 ( 
.A(n_675),
.B(n_608),
.Y(n_688)
);

AOI21xp5_ASAP7_75t_L g689 ( 
.A1(n_633),
.A2(n_612),
.B(n_52),
.Y(n_689)
);

A2O1A1Ixp33_ASAP7_75t_L g690 ( 
.A1(n_654),
.A2(n_11),
.B(n_13),
.C(n_14),
.Y(n_690)
);

NAND2xp5_ASAP7_75t_SL g691 ( 
.A(n_656),
.B(n_13),
.Y(n_691)
);

NAND2xp5_ASAP7_75t_L g692 ( 
.A(n_651),
.B(n_14),
.Y(n_692)
);

INVx1_ASAP7_75t_L g693 ( 
.A(n_650),
.Y(n_693)
);

NAND2xp5_ASAP7_75t_SL g694 ( 
.A(n_676),
.B(n_15),
.Y(n_694)
);

A2O1A1Ixp33_ASAP7_75t_L g695 ( 
.A1(n_673),
.A2(n_15),
.B(n_17),
.C(n_18),
.Y(n_695)
);

NOR2xp33_ASAP7_75t_SL g696 ( 
.A(n_646),
.B(n_51),
.Y(n_696)
);

OAI22xp5_ASAP7_75t_L g697 ( 
.A1(n_636),
.A2(n_18),
.B1(n_19),
.B2(n_20),
.Y(n_697)
);

AO31x2_ASAP7_75t_L g698 ( 
.A1(n_659),
.A2(n_117),
.A3(n_198),
.B(n_197),
.Y(n_698)
);

AOI21xp5_ASAP7_75t_L g699 ( 
.A1(n_629),
.A2(n_116),
.B(n_196),
.Y(n_699)
);

NAND2xp5_ASAP7_75t_L g700 ( 
.A(n_631),
.B(n_19),
.Y(n_700)
);

AOI21xp5_ASAP7_75t_L g701 ( 
.A1(n_642),
.A2(n_200),
.B(n_115),
.Y(n_701)
);

AOI21xp5_ASAP7_75t_L g702 ( 
.A1(n_641),
.A2(n_193),
.B(n_113),
.Y(n_702)
);

INVx1_ASAP7_75t_L g703 ( 
.A(n_643),
.Y(n_703)
);

A2O1A1Ixp33_ASAP7_75t_L g704 ( 
.A1(n_657),
.A2(n_20),
.B(n_21),
.C(n_22),
.Y(n_704)
);

OAI22xp5_ASAP7_75t_L g705 ( 
.A1(n_682),
.A2(n_658),
.B1(n_662),
.B2(n_638),
.Y(n_705)
);

NAND2xp5_ASAP7_75t_L g706 ( 
.A(n_632),
.B(n_21),
.Y(n_706)
);

AND2x6_ASAP7_75t_L g707 ( 
.A(n_661),
.B(n_53),
.Y(n_707)
);

AOI21xp5_ASAP7_75t_L g708 ( 
.A1(n_630),
.A2(n_119),
.B(n_191),
.Y(n_708)
);

OAI21x1_ASAP7_75t_L g709 ( 
.A1(n_634),
.A2(n_118),
.B(n_187),
.Y(n_709)
);

OR2x2_ASAP7_75t_L g710 ( 
.A(n_663),
.B(n_22),
.Y(n_710)
);

NAND2xp5_ASAP7_75t_L g711 ( 
.A(n_632),
.B(n_23),
.Y(n_711)
);

AO31x2_ASAP7_75t_L g712 ( 
.A1(n_645),
.A2(n_23),
.A3(n_24),
.B(n_25),
.Y(n_712)
);

INVx1_ASAP7_75t_L g713 ( 
.A(n_677),
.Y(n_713)
);

HB1xp67_ASAP7_75t_L g714 ( 
.A(n_661),
.Y(n_714)
);

OAI21xp5_ASAP7_75t_L g715 ( 
.A1(n_639),
.A2(n_25),
.B(n_26),
.Y(n_715)
);

OAI21x1_ASAP7_75t_L g716 ( 
.A1(n_674),
.A2(n_121),
.B(n_184),
.Y(n_716)
);

AOI21xp5_ASAP7_75t_L g717 ( 
.A1(n_655),
.A2(n_120),
.B(n_183),
.Y(n_717)
);

AOI21xp5_ASAP7_75t_L g718 ( 
.A1(n_672),
.A2(n_112),
.B(n_182),
.Y(n_718)
);

AOI21xp5_ASAP7_75t_L g719 ( 
.A1(n_672),
.A2(n_111),
.B(n_180),
.Y(n_719)
);

NAND2xp5_ASAP7_75t_L g720 ( 
.A(n_669),
.B(n_26),
.Y(n_720)
);

NOR2xp67_ASAP7_75t_L g721 ( 
.A(n_635),
.B(n_54),
.Y(n_721)
);

BUFx6f_ASAP7_75t_L g722 ( 
.A(n_682),
.Y(n_722)
);

NOR2x1_ASAP7_75t_SL g723 ( 
.A(n_682),
.B(n_55),
.Y(n_723)
);

AOI21xp5_ASAP7_75t_L g724 ( 
.A1(n_681),
.A2(n_185),
.B(n_122),
.Y(n_724)
);

OAI22xp5_ASAP7_75t_L g725 ( 
.A1(n_664),
.A2(n_667),
.B1(n_670),
.B2(n_644),
.Y(n_725)
);

OAI21x1_ASAP7_75t_L g726 ( 
.A1(n_666),
.A2(n_110),
.B(n_177),
.Y(n_726)
);

AOI21xp5_ASAP7_75t_L g727 ( 
.A1(n_679),
.A2(n_175),
.B(n_109),
.Y(n_727)
);

OR2x2_ASAP7_75t_L g728 ( 
.A(n_648),
.B(n_27),
.Y(n_728)
);

INVx3_ASAP7_75t_L g729 ( 
.A(n_671),
.Y(n_729)
);

AOI21xp5_ASAP7_75t_L g730 ( 
.A1(n_653),
.A2(n_123),
.B(n_173),
.Y(n_730)
);

OAI21xp5_ASAP7_75t_L g731 ( 
.A1(n_678),
.A2(n_680),
.B(n_644),
.Y(n_731)
);

OR2x6_ASAP7_75t_L g732 ( 
.A(n_661),
.B(n_56),
.Y(n_732)
);

OAI21x1_ASAP7_75t_L g733 ( 
.A1(n_649),
.A2(n_107),
.B(n_172),
.Y(n_733)
);

AO21x2_ASAP7_75t_L g734 ( 
.A1(n_628),
.A2(n_106),
.B(n_171),
.Y(n_734)
);

AOI21xp5_ASAP7_75t_L g735 ( 
.A1(n_649),
.A2(n_174),
.B(n_105),
.Y(n_735)
);

AO31x2_ASAP7_75t_L g736 ( 
.A1(n_628),
.A2(n_104),
.A3(n_170),
.B(n_169),
.Y(n_736)
);

AOI21xp5_ASAP7_75t_L g737 ( 
.A1(n_649),
.A2(n_103),
.B(n_165),
.Y(n_737)
);

INVx5_ASAP7_75t_L g738 ( 
.A(n_671),
.Y(n_738)
);

OAI21x1_ASAP7_75t_L g739 ( 
.A1(n_649),
.A2(n_102),
.B(n_164),
.Y(n_739)
);

INVx3_ASAP7_75t_L g740 ( 
.A(n_665),
.Y(n_740)
);

AND2x2_ASAP7_75t_L g741 ( 
.A(n_665),
.B(n_28),
.Y(n_741)
);

INVx3_ASAP7_75t_L g742 ( 
.A(n_722),
.Y(n_742)
);

CKINVDCx6p67_ASAP7_75t_R g743 ( 
.A(n_738),
.Y(n_743)
);

BUFx2_ASAP7_75t_L g744 ( 
.A(n_722),
.Y(n_744)
);

INVx2_ASAP7_75t_L g745 ( 
.A(n_687),
.Y(n_745)
);

CKINVDCx16_ASAP7_75t_R g746 ( 
.A(n_696),
.Y(n_746)
);

INVx8_ASAP7_75t_L g747 ( 
.A(n_707),
.Y(n_747)
);

AOI22xp33_ASAP7_75t_SL g748 ( 
.A1(n_715),
.A2(n_668),
.B1(n_30),
.B2(n_29),
.Y(n_748)
);

INVx1_ASAP7_75t_L g749 ( 
.A(n_703),
.Y(n_749)
);

INVx6_ASAP7_75t_L g750 ( 
.A(n_738),
.Y(n_750)
);

BUFx3_ASAP7_75t_L g751 ( 
.A(n_684),
.Y(n_751)
);

INVx2_ASAP7_75t_SL g752 ( 
.A(n_738),
.Y(n_752)
);

INVx2_ASAP7_75t_L g753 ( 
.A(n_693),
.Y(n_753)
);

INVx1_ASAP7_75t_SL g754 ( 
.A(n_713),
.Y(n_754)
);

AOI22xp33_ASAP7_75t_L g755 ( 
.A1(n_686),
.A2(n_57),
.B1(n_58),
.B2(n_59),
.Y(n_755)
);

INVx8_ASAP7_75t_L g756 ( 
.A(n_707),
.Y(n_756)
);

BUFx2_ASAP7_75t_R g757 ( 
.A(n_694),
.Y(n_757)
);

INVx1_ASAP7_75t_L g758 ( 
.A(n_740),
.Y(n_758)
);

INVx1_ASAP7_75t_SL g759 ( 
.A(n_714),
.Y(n_759)
);

BUFx2_ASAP7_75t_SL g760 ( 
.A(n_729),
.Y(n_760)
);

CKINVDCx20_ASAP7_75t_R g761 ( 
.A(n_705),
.Y(n_761)
);

INVx6_ASAP7_75t_L g762 ( 
.A(n_732),
.Y(n_762)
);

CKINVDCx11_ASAP7_75t_R g763 ( 
.A(n_732),
.Y(n_763)
);

AOI22xp33_ASAP7_75t_L g764 ( 
.A1(n_691),
.A2(n_60),
.B1(n_63),
.B2(n_64),
.Y(n_764)
);

AOI22xp33_ASAP7_75t_L g765 ( 
.A1(n_697),
.A2(n_67),
.B1(n_71),
.B2(n_72),
.Y(n_765)
);

AOI22xp33_ASAP7_75t_L g766 ( 
.A1(n_688),
.A2(n_74),
.B1(n_75),
.B2(n_76),
.Y(n_766)
);

INVx2_ASAP7_75t_L g767 ( 
.A(n_728),
.Y(n_767)
);

AOI22xp33_ASAP7_75t_L g768 ( 
.A1(n_741),
.A2(n_77),
.B1(n_79),
.B2(n_80),
.Y(n_768)
);

INVx2_ASAP7_75t_SL g769 ( 
.A(n_692),
.Y(n_769)
);

BUFx4f_ASAP7_75t_SL g770 ( 
.A(n_707),
.Y(n_770)
);

INVx3_ASAP7_75t_SL g771 ( 
.A(n_710),
.Y(n_771)
);

INVx1_ASAP7_75t_SL g772 ( 
.A(n_706),
.Y(n_772)
);

INVx1_ASAP7_75t_L g773 ( 
.A(n_712),
.Y(n_773)
);

BUFx4f_ASAP7_75t_SL g774 ( 
.A(n_723),
.Y(n_774)
);

INVx2_ASAP7_75t_SL g775 ( 
.A(n_711),
.Y(n_775)
);

NAND2xp5_ASAP7_75t_L g776 ( 
.A(n_700),
.B(n_81),
.Y(n_776)
);

CKINVDCx5p33_ASAP7_75t_R g777 ( 
.A(n_720),
.Y(n_777)
);

AOI22xp33_ASAP7_75t_SL g778 ( 
.A1(n_702),
.A2(n_82),
.B1(n_84),
.B2(n_85),
.Y(n_778)
);

AOI22xp33_ASAP7_75t_L g779 ( 
.A1(n_725),
.A2(n_86),
.B1(n_88),
.B2(n_90),
.Y(n_779)
);

OAI22xp33_ASAP7_75t_L g780 ( 
.A1(n_735),
.A2(n_737),
.B1(n_689),
.B2(n_717),
.Y(n_780)
);

BUFx4f_ASAP7_75t_SL g781 ( 
.A(n_721),
.Y(n_781)
);

INVx1_ASAP7_75t_L g782 ( 
.A(n_712),
.Y(n_782)
);

INVx1_ASAP7_75t_L g783 ( 
.A(n_712),
.Y(n_783)
);

CKINVDCx11_ASAP7_75t_R g784 ( 
.A(n_685),
.Y(n_784)
);

BUFx10_ASAP7_75t_L g785 ( 
.A(n_690),
.Y(n_785)
);

INVx6_ASAP7_75t_L g786 ( 
.A(n_731),
.Y(n_786)
);

HB1xp67_ASAP7_75t_L g787 ( 
.A(n_736),
.Y(n_787)
);

CKINVDCx11_ASAP7_75t_R g788 ( 
.A(n_704),
.Y(n_788)
);

INVx1_ASAP7_75t_L g789 ( 
.A(n_736),
.Y(n_789)
);

INVx1_ASAP7_75t_L g790 ( 
.A(n_734),
.Y(n_790)
);

INVx3_ASAP7_75t_L g791 ( 
.A(n_733),
.Y(n_791)
);

BUFx2_ASAP7_75t_L g792 ( 
.A(n_739),
.Y(n_792)
);

BUFx3_ASAP7_75t_L g793 ( 
.A(n_709),
.Y(n_793)
);

INVx4_ASAP7_75t_L g794 ( 
.A(n_683),
.Y(n_794)
);

CKINVDCx6p67_ASAP7_75t_R g795 ( 
.A(n_695),
.Y(n_795)
);

AOI22xp33_ASAP7_75t_SL g796 ( 
.A1(n_724),
.A2(n_91),
.B1(n_93),
.B2(n_95),
.Y(n_796)
);

INVx1_ASAP7_75t_SL g797 ( 
.A(n_683),
.Y(n_797)
);

BUFx6f_ASAP7_75t_SL g798 ( 
.A(n_699),
.Y(n_798)
);

NAND2xp5_ASAP7_75t_L g799 ( 
.A(n_754),
.B(n_708),
.Y(n_799)
);

INVx1_ASAP7_75t_L g800 ( 
.A(n_773),
.Y(n_800)
);

INVx1_ASAP7_75t_L g801 ( 
.A(n_782),
.Y(n_801)
);

AOI22xp33_ASAP7_75t_L g802 ( 
.A1(n_788),
.A2(n_730),
.B1(n_727),
.B2(n_718),
.Y(n_802)
);

INVx3_ASAP7_75t_L g803 ( 
.A(n_794),
.Y(n_803)
);

INVx1_ASAP7_75t_L g804 ( 
.A(n_783),
.Y(n_804)
);

AOI22xp33_ASAP7_75t_SL g805 ( 
.A1(n_785),
.A2(n_701),
.B1(n_719),
.B2(n_716),
.Y(n_805)
);

INVx2_ASAP7_75t_L g806 ( 
.A(n_749),
.Y(n_806)
);

INVx1_ASAP7_75t_L g807 ( 
.A(n_789),
.Y(n_807)
);

INVx3_ASAP7_75t_L g808 ( 
.A(n_794),
.Y(n_808)
);

CKINVDCx14_ASAP7_75t_R g809 ( 
.A(n_763),
.Y(n_809)
);

INVx1_ASAP7_75t_L g810 ( 
.A(n_758),
.Y(n_810)
);

INVx2_ASAP7_75t_L g811 ( 
.A(n_797),
.Y(n_811)
);

OAI21x1_ASAP7_75t_L g812 ( 
.A1(n_791),
.A2(n_726),
.B(n_698),
.Y(n_812)
);

INVx2_ASAP7_75t_L g813 ( 
.A(n_797),
.Y(n_813)
);

INVx1_ASAP7_75t_L g814 ( 
.A(n_745),
.Y(n_814)
);

INVx2_ASAP7_75t_L g815 ( 
.A(n_753),
.Y(n_815)
);

INVx1_ASAP7_75t_L g816 ( 
.A(n_787),
.Y(n_816)
);

HB1xp67_ASAP7_75t_L g817 ( 
.A(n_754),
.Y(n_817)
);

INVx1_ASAP7_75t_L g818 ( 
.A(n_790),
.Y(n_818)
);

INVx1_ASAP7_75t_SL g819 ( 
.A(n_771),
.Y(n_819)
);

AOI22xp33_ASAP7_75t_L g820 ( 
.A1(n_795),
.A2(n_698),
.B1(n_97),
.B2(n_98),
.Y(n_820)
);

INVx1_ASAP7_75t_L g821 ( 
.A(n_786),
.Y(n_821)
);

INVx1_ASAP7_75t_L g822 ( 
.A(n_786),
.Y(n_822)
);

INVx2_ASAP7_75t_L g823 ( 
.A(n_786),
.Y(n_823)
);

AOI21xp5_ASAP7_75t_L g824 ( 
.A1(n_780),
.A2(n_96),
.B(n_124),
.Y(n_824)
);

INVx3_ASAP7_75t_L g825 ( 
.A(n_793),
.Y(n_825)
);

INVxp67_ASAP7_75t_L g826 ( 
.A(n_769),
.Y(n_826)
);

AND2x2_ASAP7_75t_L g827 ( 
.A(n_772),
.B(n_125),
.Y(n_827)
);

OR2x2_ASAP7_75t_L g828 ( 
.A(n_772),
.B(n_126),
.Y(n_828)
);

INVx2_ASAP7_75t_L g829 ( 
.A(n_792),
.Y(n_829)
);

INVx2_ASAP7_75t_L g830 ( 
.A(n_759),
.Y(n_830)
);

INVx2_ASAP7_75t_SL g831 ( 
.A(n_750),
.Y(n_831)
);

INVx2_ASAP7_75t_L g832 ( 
.A(n_759),
.Y(n_832)
);

INVx1_ASAP7_75t_L g833 ( 
.A(n_767),
.Y(n_833)
);

INVx1_ASAP7_75t_L g834 ( 
.A(n_750),
.Y(n_834)
);

INVxp67_ASAP7_75t_L g835 ( 
.A(n_744),
.Y(n_835)
);

INVxp67_ASAP7_75t_L g836 ( 
.A(n_775),
.Y(n_836)
);

INVx2_ASAP7_75t_L g837 ( 
.A(n_750),
.Y(n_837)
);

AOI22xp33_ASAP7_75t_L g838 ( 
.A1(n_785),
.A2(n_128),
.B1(n_129),
.B2(n_131),
.Y(n_838)
);

INVx2_ASAP7_75t_L g839 ( 
.A(n_752),
.Y(n_839)
);

INVx1_ASAP7_75t_L g840 ( 
.A(n_776),
.Y(n_840)
);

INVx2_ASAP7_75t_L g841 ( 
.A(n_742),
.Y(n_841)
);

INVx1_ASAP7_75t_L g842 ( 
.A(n_776),
.Y(n_842)
);

INVx1_ASAP7_75t_L g843 ( 
.A(n_800),
.Y(n_843)
);

BUFx6f_ASAP7_75t_L g844 ( 
.A(n_831),
.Y(n_844)
);

AND2x2_ASAP7_75t_L g845 ( 
.A(n_811),
.B(n_777),
.Y(n_845)
);

INVx3_ASAP7_75t_SL g846 ( 
.A(n_819),
.Y(n_846)
);

HB1xp67_ASAP7_75t_L g847 ( 
.A(n_817),
.Y(n_847)
);

INVx1_ASAP7_75t_L g848 ( 
.A(n_800),
.Y(n_848)
);

AO31x2_ASAP7_75t_L g849 ( 
.A1(n_801),
.A2(n_748),
.A3(n_798),
.B(n_796),
.Y(n_849)
);

INVx1_ASAP7_75t_L g850 ( 
.A(n_801),
.Y(n_850)
);

INVx1_ASAP7_75t_L g851 ( 
.A(n_804),
.Y(n_851)
);

BUFx12f_ASAP7_75t_L g852 ( 
.A(n_828),
.Y(n_852)
);

OR2x2_ASAP7_75t_L g853 ( 
.A(n_811),
.B(n_813),
.Y(n_853)
);

INVx3_ASAP7_75t_L g854 ( 
.A(n_803),
.Y(n_854)
);

INVx2_ASAP7_75t_L g855 ( 
.A(n_806),
.Y(n_855)
);

CKINVDCx5p33_ASAP7_75t_R g856 ( 
.A(n_809),
.Y(n_856)
);

AND2x2_ASAP7_75t_L g857 ( 
.A(n_811),
.B(n_742),
.Y(n_857)
);

AOI22xp5_ASAP7_75t_L g858 ( 
.A1(n_802),
.A2(n_798),
.B1(n_761),
.B2(n_762),
.Y(n_858)
);

INVx1_ASAP7_75t_L g859 ( 
.A(n_804),
.Y(n_859)
);

INVx2_ASAP7_75t_L g860 ( 
.A(n_815),
.Y(n_860)
);

AND2x2_ASAP7_75t_L g861 ( 
.A(n_813),
.B(n_760),
.Y(n_861)
);

INVx1_ASAP7_75t_L g862 ( 
.A(n_818),
.Y(n_862)
);

AND2x2_ASAP7_75t_L g863 ( 
.A(n_813),
.B(n_746),
.Y(n_863)
);

AO21x1_ASAP7_75t_SL g864 ( 
.A1(n_799),
.A2(n_768),
.B(n_779),
.Y(n_864)
);

HB1xp67_ASAP7_75t_L g865 ( 
.A(n_830),
.Y(n_865)
);

OR2x6_ASAP7_75t_L g866 ( 
.A(n_829),
.B(n_756),
.Y(n_866)
);

AOI21x1_ASAP7_75t_L g867 ( 
.A1(n_818),
.A2(n_784),
.B(n_743),
.Y(n_867)
);

AO21x2_ASAP7_75t_L g868 ( 
.A1(n_812),
.A2(n_778),
.B(n_796),
.Y(n_868)
);

AND2x2_ASAP7_75t_L g869 ( 
.A(n_829),
.B(n_762),
.Y(n_869)
);

INVx2_ASAP7_75t_L g870 ( 
.A(n_815),
.Y(n_870)
);

NAND2xp5_ASAP7_75t_L g871 ( 
.A(n_840),
.B(n_762),
.Y(n_871)
);

HB1xp67_ASAP7_75t_L g872 ( 
.A(n_830),
.Y(n_872)
);

OR2x2_ASAP7_75t_L g873 ( 
.A(n_832),
.B(n_756),
.Y(n_873)
);

AND2x2_ASAP7_75t_L g874 ( 
.A(n_810),
.B(n_778),
.Y(n_874)
);

INVx1_ASAP7_75t_L g875 ( 
.A(n_807),
.Y(n_875)
);

INVx1_ASAP7_75t_L g876 ( 
.A(n_807),
.Y(n_876)
);

OA21x2_ASAP7_75t_L g877 ( 
.A1(n_812),
.A2(n_765),
.B(n_764),
.Y(n_877)
);

INVx1_ASAP7_75t_L g878 ( 
.A(n_862),
.Y(n_878)
);

BUFx2_ASAP7_75t_L g879 ( 
.A(n_854),
.Y(n_879)
);

INVx1_ASAP7_75t_L g880 ( 
.A(n_862),
.Y(n_880)
);

INVx2_ASAP7_75t_L g881 ( 
.A(n_853),
.Y(n_881)
);

NAND2xp5_ASAP7_75t_L g882 ( 
.A(n_847),
.B(n_832),
.Y(n_882)
);

INVx1_ASAP7_75t_L g883 ( 
.A(n_875),
.Y(n_883)
);

AND2x2_ASAP7_75t_L g884 ( 
.A(n_869),
.B(n_803),
.Y(n_884)
);

AND2x6_ASAP7_75t_L g885 ( 
.A(n_874),
.B(n_822),
.Y(n_885)
);

INVx2_ASAP7_75t_L g886 ( 
.A(n_853),
.Y(n_886)
);

NAND2xp5_ASAP7_75t_L g887 ( 
.A(n_871),
.B(n_842),
.Y(n_887)
);

AOI21xp5_ASAP7_75t_L g888 ( 
.A1(n_868),
.A2(n_824),
.B(n_756),
.Y(n_888)
);

INVxp67_ASAP7_75t_SL g889 ( 
.A(n_865),
.Y(n_889)
);

INVx1_ASAP7_75t_L g890 ( 
.A(n_875),
.Y(n_890)
);

NAND2xp5_ASAP7_75t_L g891 ( 
.A(n_845),
.B(n_842),
.Y(n_891)
);

HB1xp67_ASAP7_75t_L g892 ( 
.A(n_872),
.Y(n_892)
);

NOR2xp33_ASAP7_75t_L g893 ( 
.A(n_846),
.B(n_826),
.Y(n_893)
);

AND2x2_ASAP7_75t_L g894 ( 
.A(n_869),
.B(n_803),
.Y(n_894)
);

AND2x2_ASAP7_75t_L g895 ( 
.A(n_845),
.B(n_803),
.Y(n_895)
);

INVx2_ASAP7_75t_SL g896 ( 
.A(n_844),
.Y(n_896)
);

AND2x2_ASAP7_75t_L g897 ( 
.A(n_863),
.B(n_808),
.Y(n_897)
);

INVx2_ASAP7_75t_L g898 ( 
.A(n_876),
.Y(n_898)
);

INVx2_ASAP7_75t_L g899 ( 
.A(n_876),
.Y(n_899)
);

INVx2_ASAP7_75t_L g900 ( 
.A(n_843),
.Y(n_900)
);

INVx2_ASAP7_75t_L g901 ( 
.A(n_843),
.Y(n_901)
);

OR2x2_ASAP7_75t_L g902 ( 
.A(n_891),
.B(n_882),
.Y(n_902)
);

OR2x2_ASAP7_75t_L g903 ( 
.A(n_892),
.B(n_863),
.Y(n_903)
);

AND2x2_ASAP7_75t_L g904 ( 
.A(n_884),
.B(n_861),
.Y(n_904)
);

NAND2xp5_ASAP7_75t_L g905 ( 
.A(n_887),
.B(n_861),
.Y(n_905)
);

AND2x2_ASAP7_75t_L g906 ( 
.A(n_884),
.B(n_857),
.Y(n_906)
);

AND2x2_ASAP7_75t_L g907 ( 
.A(n_894),
.B(n_857),
.Y(n_907)
);

INVx4_ASAP7_75t_L g908 ( 
.A(n_885),
.Y(n_908)
);

AND2x2_ASAP7_75t_L g909 ( 
.A(n_894),
.B(n_846),
.Y(n_909)
);

NAND2xp5_ASAP7_75t_L g910 ( 
.A(n_889),
.B(n_874),
.Y(n_910)
);

INVx1_ASAP7_75t_L g911 ( 
.A(n_883),
.Y(n_911)
);

NAND2x1_ASAP7_75t_L g912 ( 
.A(n_885),
.B(n_854),
.Y(n_912)
);

AND2x2_ASAP7_75t_L g913 ( 
.A(n_897),
.B(n_846),
.Y(n_913)
);

BUFx2_ASAP7_75t_L g914 ( 
.A(n_885),
.Y(n_914)
);

INVx1_ASAP7_75t_SL g915 ( 
.A(n_895),
.Y(n_915)
);

INVx1_ASAP7_75t_L g916 ( 
.A(n_883),
.Y(n_916)
);

AND2x2_ASAP7_75t_L g917 ( 
.A(n_909),
.B(n_895),
.Y(n_917)
);

INVx2_ASAP7_75t_L g918 ( 
.A(n_911),
.Y(n_918)
);

INVx1_ASAP7_75t_L g919 ( 
.A(n_916),
.Y(n_919)
);

HB1xp67_ASAP7_75t_L g920 ( 
.A(n_910),
.Y(n_920)
);

INVx1_ASAP7_75t_L g921 ( 
.A(n_903),
.Y(n_921)
);

OR2x2_ASAP7_75t_L g922 ( 
.A(n_902),
.B(n_881),
.Y(n_922)
);

AND2x2_ASAP7_75t_L g923 ( 
.A(n_909),
.B(n_897),
.Y(n_923)
);

NAND2x1_ASAP7_75t_L g924 ( 
.A(n_908),
.B(n_885),
.Y(n_924)
);

AND2x2_ASAP7_75t_L g925 ( 
.A(n_913),
.B(n_893),
.Y(n_925)
);

INVx2_ASAP7_75t_L g926 ( 
.A(n_913),
.Y(n_926)
);

NAND2xp5_ASAP7_75t_L g927 ( 
.A(n_905),
.B(n_878),
.Y(n_927)
);

OR2x2_ASAP7_75t_L g928 ( 
.A(n_915),
.B(n_881),
.Y(n_928)
);

NAND2xp5_ASAP7_75t_L g929 ( 
.A(n_920),
.B(n_904),
.Y(n_929)
);

AND2x2_ASAP7_75t_L g930 ( 
.A(n_925),
.B(n_926),
.Y(n_930)
);

INVx3_ASAP7_75t_SL g931 ( 
.A(n_928),
.Y(n_931)
);

INVx1_ASAP7_75t_L g932 ( 
.A(n_918),
.Y(n_932)
);

OR2x2_ASAP7_75t_L g933 ( 
.A(n_921),
.B(n_904),
.Y(n_933)
);

INVx1_ASAP7_75t_L g934 ( 
.A(n_919),
.Y(n_934)
);

INVx2_ASAP7_75t_L g935 ( 
.A(n_923),
.Y(n_935)
);

INVx1_ASAP7_75t_L g936 ( 
.A(n_918),
.Y(n_936)
);

INVx2_ASAP7_75t_L g937 ( 
.A(n_917),
.Y(n_937)
);

NAND2xp33_ASAP7_75t_R g938 ( 
.A(n_930),
.B(n_856),
.Y(n_938)
);

OR2x2_ASAP7_75t_L g939 ( 
.A(n_931),
.B(n_920),
.Y(n_939)
);

AOI22xp5_ASAP7_75t_L g940 ( 
.A1(n_935),
.A2(n_908),
.B1(n_914),
.B2(n_924),
.Y(n_940)
);

AO221x2_ASAP7_75t_L g941 ( 
.A1(n_934),
.A2(n_856),
.B1(n_927),
.B2(n_908),
.C(n_821),
.Y(n_941)
);

INVx1_ASAP7_75t_L g942 ( 
.A(n_932),
.Y(n_942)
);

AOI22xp5_ASAP7_75t_L g943 ( 
.A1(n_937),
.A2(n_885),
.B1(n_888),
.B2(n_858),
.Y(n_943)
);

NAND2xp5_ASAP7_75t_L g944 ( 
.A(n_929),
.B(n_927),
.Y(n_944)
);

NAND2xp5_ASAP7_75t_L g945 ( 
.A(n_933),
.B(n_932),
.Y(n_945)
);

OR2x2_ASAP7_75t_L g946 ( 
.A(n_939),
.B(n_922),
.Y(n_946)
);

INVx1_ASAP7_75t_SL g947 ( 
.A(n_945),
.Y(n_947)
);

AOI22xp5_ASAP7_75t_L g948 ( 
.A1(n_938),
.A2(n_941),
.B1(n_943),
.B2(n_940),
.Y(n_948)
);

NAND2xp5_ASAP7_75t_L g949 ( 
.A(n_942),
.B(n_936),
.Y(n_949)
);

NAND2xp5_ASAP7_75t_SL g950 ( 
.A(n_944),
.B(n_936),
.Y(n_950)
);

INVx1_ASAP7_75t_SL g951 ( 
.A(n_941),
.Y(n_951)
);

INVx1_ASAP7_75t_L g952 ( 
.A(n_942),
.Y(n_952)
);

NOR3xp33_ASAP7_75t_L g953 ( 
.A(n_939),
.B(n_867),
.C(n_827),
.Y(n_953)
);

HB1xp67_ASAP7_75t_L g954 ( 
.A(n_939),
.Y(n_954)
);

INVx1_ASAP7_75t_L g955 ( 
.A(n_942),
.Y(n_955)
);

AND2x2_ASAP7_75t_L g956 ( 
.A(n_939),
.B(n_906),
.Y(n_956)
);

NAND4xp25_ASAP7_75t_L g957 ( 
.A(n_948),
.B(n_751),
.C(n_836),
.D(n_766),
.Y(n_957)
);

OAI32xp33_ASAP7_75t_L g958 ( 
.A1(n_951),
.A2(n_896),
.A3(n_873),
.B1(n_828),
.B2(n_840),
.Y(n_958)
);

AOI21xp33_ASAP7_75t_L g959 ( 
.A1(n_954),
.A2(n_912),
.B(n_839),
.Y(n_959)
);

NAND2xp5_ASAP7_75t_SL g960 ( 
.A(n_946),
.B(n_867),
.Y(n_960)
);

NOR2xp33_ASAP7_75t_L g961 ( 
.A(n_947),
.B(n_852),
.Y(n_961)
);

AND2x2_ASAP7_75t_L g962 ( 
.A(n_956),
.B(n_906),
.Y(n_962)
);

NAND2xp5_ASAP7_75t_L g963 ( 
.A(n_950),
.B(n_907),
.Y(n_963)
);

AOI22xp33_ASAP7_75t_L g964 ( 
.A1(n_953),
.A2(n_868),
.B1(n_864),
.B2(n_885),
.Y(n_964)
);

AOI322xp5_ASAP7_75t_L g965 ( 
.A1(n_955),
.A2(n_852),
.A3(n_907),
.B1(n_827),
.B2(n_896),
.C1(n_879),
.C2(n_820),
.Y(n_965)
);

INVx1_ASAP7_75t_L g966 ( 
.A(n_963),
.Y(n_966)
);

INVx1_ASAP7_75t_L g967 ( 
.A(n_962),
.Y(n_967)
);

INVx1_ASAP7_75t_SL g968 ( 
.A(n_960),
.Y(n_968)
);

NAND2xp5_ASAP7_75t_L g969 ( 
.A(n_961),
.B(n_952),
.Y(n_969)
);

AOI21xp5_ASAP7_75t_L g970 ( 
.A1(n_957),
.A2(n_949),
.B(n_747),
.Y(n_970)
);

NAND2xp5_ASAP7_75t_L g971 ( 
.A(n_965),
.B(n_949),
.Y(n_971)
);

AND2x2_ASAP7_75t_L g972 ( 
.A(n_964),
.B(n_886),
.Y(n_972)
);

INVx2_ASAP7_75t_L g973 ( 
.A(n_959),
.Y(n_973)
);

OAI21xp33_ASAP7_75t_L g974 ( 
.A1(n_971),
.A2(n_958),
.B(n_821),
.Y(n_974)
);

INVxp67_ASAP7_75t_L g975 ( 
.A(n_967),
.Y(n_975)
);

AOI221x1_ASAP7_75t_L g976 ( 
.A1(n_969),
.A2(n_839),
.B1(n_890),
.B2(n_880),
.C(n_834),
.Y(n_976)
);

OAI211xp5_ASAP7_75t_SL g977 ( 
.A1(n_966),
.A2(n_838),
.B(n_835),
.C(n_755),
.Y(n_977)
);

OAI22xp5_ASAP7_75t_L g978 ( 
.A1(n_968),
.A2(n_770),
.B1(n_879),
.B2(n_774),
.Y(n_978)
);

INVx2_ASAP7_75t_L g979 ( 
.A(n_975),
.Y(n_979)
);

INVx2_ASAP7_75t_L g980 ( 
.A(n_978),
.Y(n_980)
);

INVx1_ASAP7_75t_L g981 ( 
.A(n_974),
.Y(n_981)
);

INVx1_ASAP7_75t_L g982 ( 
.A(n_976),
.Y(n_982)
);

INVx1_ASAP7_75t_L g983 ( 
.A(n_977),
.Y(n_983)
);

INVx1_ASAP7_75t_L g984 ( 
.A(n_975),
.Y(n_984)
);

NOR2x1_ASAP7_75t_L g985 ( 
.A(n_979),
.B(n_968),
.Y(n_985)
);

HB1xp67_ASAP7_75t_L g986 ( 
.A(n_982),
.Y(n_986)
);

NOR2xp33_ASAP7_75t_L g987 ( 
.A(n_981),
.B(n_984),
.Y(n_987)
);

NOR3xp33_ASAP7_75t_L g988 ( 
.A(n_980),
.B(n_970),
.C(n_973),
.Y(n_988)
);

OAI322xp33_ASAP7_75t_L g989 ( 
.A1(n_981),
.A2(n_972),
.A3(n_873),
.B1(n_822),
.B2(n_841),
.C1(n_831),
.C2(n_833),
.Y(n_989)
);

NOR2x1_ASAP7_75t_L g990 ( 
.A(n_983),
.B(n_868),
.Y(n_990)
);

AOI22x1_ASAP7_75t_L g991 ( 
.A1(n_986),
.A2(n_823),
.B1(n_837),
.B2(n_834),
.Y(n_991)
);

NOR2xp67_ASAP7_75t_L g992 ( 
.A(n_987),
.B(n_132),
.Y(n_992)
);

NAND2xp5_ASAP7_75t_L g993 ( 
.A(n_985),
.B(n_833),
.Y(n_993)
);

NAND2xp5_ASAP7_75t_L g994 ( 
.A(n_988),
.B(n_901),
.Y(n_994)
);

NAND2xp5_ASAP7_75t_L g995 ( 
.A(n_992),
.B(n_993),
.Y(n_995)
);

BUFx6f_ASAP7_75t_L g996 ( 
.A(n_994),
.Y(n_996)
);

AOI211xp5_ASAP7_75t_L g997 ( 
.A1(n_991),
.A2(n_989),
.B(n_990),
.C(n_844),
.Y(n_997)
);

NAND4xp25_ASAP7_75t_L g998 ( 
.A(n_994),
.B(n_823),
.C(n_805),
.D(n_837),
.Y(n_998)
);

XNOR2xp5_ASAP7_75t_L g999 ( 
.A(n_992),
.B(n_134),
.Y(n_999)
);

OAI221xp5_ASAP7_75t_L g1000 ( 
.A1(n_994),
.A2(n_866),
.B1(n_844),
.B2(n_886),
.C(n_841),
.Y(n_1000)
);

OAI211xp5_ASAP7_75t_L g1001 ( 
.A1(n_992),
.A2(n_747),
.B(n_844),
.C(n_854),
.Y(n_1001)
);

NOR4xp25_ASAP7_75t_L g1002 ( 
.A(n_994),
.B(n_901),
.C(n_900),
.D(n_899),
.Y(n_1002)
);

INVx2_ASAP7_75t_L g1003 ( 
.A(n_999),
.Y(n_1003)
);

NOR3xp33_ASAP7_75t_SL g1004 ( 
.A(n_995),
.B(n_747),
.C(n_781),
.Y(n_1004)
);

INVxp67_ASAP7_75t_SL g1005 ( 
.A(n_996),
.Y(n_1005)
);

NAND2xp5_ASAP7_75t_L g1006 ( 
.A(n_996),
.B(n_900),
.Y(n_1006)
);

AND4x1_ASAP7_75t_L g1007 ( 
.A(n_997),
.B(n_757),
.C(n_137),
.D(n_140),
.Y(n_1007)
);

AND3x2_ASAP7_75t_L g1008 ( 
.A(n_1002),
.B(n_757),
.C(n_142),
.Y(n_1008)
);

OAI322xp33_ASAP7_75t_L g1009 ( 
.A1(n_1000),
.A2(n_1001),
.A3(n_998),
.B1(n_844),
.B2(n_898),
.C1(n_899),
.C2(n_816),
.Y(n_1009)
);

INVx1_ASAP7_75t_L g1010 ( 
.A(n_999),
.Y(n_1010)
);

AOI22xp33_ASAP7_75t_L g1011 ( 
.A1(n_996),
.A2(n_864),
.B1(n_877),
.B2(n_866),
.Y(n_1011)
);

AND2x4_ASAP7_75t_L g1012 ( 
.A(n_1004),
.B(n_866),
.Y(n_1012)
);

OR2x2_ASAP7_75t_L g1013 ( 
.A(n_1005),
.B(n_849),
.Y(n_1013)
);

BUFx3_ASAP7_75t_L g1014 ( 
.A(n_1003),
.Y(n_1014)
);

NAND2xp5_ASAP7_75t_L g1015 ( 
.A(n_1008),
.B(n_898),
.Y(n_1015)
);

INVx2_ASAP7_75t_L g1016 ( 
.A(n_1010),
.Y(n_1016)
);

INVx4_ASAP7_75t_L g1017 ( 
.A(n_1007),
.Y(n_1017)
);

NAND3xp33_ASAP7_75t_L g1018 ( 
.A(n_1006),
.B(n_866),
.C(n_816),
.Y(n_1018)
);

INVx3_ASAP7_75t_SL g1019 ( 
.A(n_1009),
.Y(n_1019)
);

INVx1_ASAP7_75t_L g1020 ( 
.A(n_1011),
.Y(n_1020)
);

INVx1_ASAP7_75t_L g1021 ( 
.A(n_1005),
.Y(n_1021)
);

AND2x2_ASAP7_75t_L g1022 ( 
.A(n_1004),
.B(n_849),
.Y(n_1022)
);

AND2x4_ASAP7_75t_L g1023 ( 
.A(n_1004),
.B(n_849),
.Y(n_1023)
);

AND2x2_ASAP7_75t_L g1024 ( 
.A(n_1004),
.B(n_849),
.Y(n_1024)
);

OA21x2_ASAP7_75t_L g1025 ( 
.A1(n_1021),
.A2(n_1020),
.B(n_1016),
.Y(n_1025)
);

AND2x2_ASAP7_75t_L g1026 ( 
.A(n_1012),
.B(n_849),
.Y(n_1026)
);

XOR2xp5_ASAP7_75t_L g1027 ( 
.A(n_1014),
.B(n_135),
.Y(n_1027)
);

AO22x2_ASAP7_75t_L g1028 ( 
.A1(n_1017),
.A2(n_851),
.B1(n_850),
.B2(n_848),
.Y(n_1028)
);

INVxp67_ASAP7_75t_L g1029 ( 
.A(n_1013),
.Y(n_1029)
);

NAND2xp5_ASAP7_75t_L g1030 ( 
.A(n_1019),
.B(n_814),
.Y(n_1030)
);

OAI221xp5_ASAP7_75t_L g1031 ( 
.A1(n_1015),
.A2(n_825),
.B1(n_808),
.B2(n_814),
.C(n_877),
.Y(n_1031)
);

CKINVDCx20_ASAP7_75t_R g1032 ( 
.A(n_1022),
.Y(n_1032)
);

NAND2xp33_ASAP7_75t_SL g1033 ( 
.A(n_1024),
.B(n_825),
.Y(n_1033)
);

AOI22xp5_ASAP7_75t_L g1034 ( 
.A1(n_1032),
.A2(n_1024),
.B1(n_1023),
.B2(n_1018),
.Y(n_1034)
);

INVx1_ASAP7_75t_L g1035 ( 
.A(n_1025),
.Y(n_1035)
);

AO22x2_ASAP7_75t_L g1036 ( 
.A1(n_1029),
.A2(n_825),
.B1(n_808),
.B2(n_848),
.Y(n_1036)
);

AO22x2_ASAP7_75t_L g1037 ( 
.A1(n_1027),
.A2(n_825),
.B1(n_808),
.B2(n_859),
.Y(n_1037)
);

INVx1_ASAP7_75t_L g1038 ( 
.A(n_1030),
.Y(n_1038)
);

NAND4xp25_ASAP7_75t_L g1039 ( 
.A(n_1033),
.B(n_144),
.C(n_145),
.D(n_146),
.Y(n_1039)
);

AND2x2_ASAP7_75t_L g1040 ( 
.A(n_1034),
.B(n_1026),
.Y(n_1040)
);

OAI22xp5_ASAP7_75t_L g1041 ( 
.A1(n_1035),
.A2(n_1031),
.B1(n_1028),
.B2(n_851),
.Y(n_1041)
);

XNOR2xp5_ASAP7_75t_L g1042 ( 
.A(n_1038),
.B(n_1039),
.Y(n_1042)
);

AOI22xp33_ASAP7_75t_SL g1043 ( 
.A1(n_1040),
.A2(n_1037),
.B1(n_1036),
.B2(n_1028),
.Y(n_1043)
);

NOR2xp67_ASAP7_75t_L g1044 ( 
.A(n_1043),
.B(n_1042),
.Y(n_1044)
);

AOI21xp5_ASAP7_75t_L g1045 ( 
.A1(n_1044),
.A2(n_1041),
.B(n_149),
.Y(n_1045)
);

AOI22xp5_ASAP7_75t_L g1046 ( 
.A1(n_1045),
.A2(n_877),
.B1(n_850),
.B2(n_859),
.Y(n_1046)
);

AOI22xp33_ASAP7_75t_L g1047 ( 
.A1(n_1045),
.A2(n_870),
.B1(n_860),
.B2(n_877),
.Y(n_1047)
);

OAI22xp5_ASAP7_75t_L g1048 ( 
.A1(n_1045),
.A2(n_870),
.B1(n_860),
.B2(n_855),
.Y(n_1048)
);

HB1xp67_ASAP7_75t_L g1049 ( 
.A(n_1048),
.Y(n_1049)
);

NAND2xp5_ASAP7_75t_L g1050 ( 
.A(n_1046),
.B(n_148),
.Y(n_1050)
);

AND2x2_ASAP7_75t_L g1051 ( 
.A(n_1047),
.B(n_855),
.Y(n_1051)
);

OA21x2_ASAP7_75t_L g1052 ( 
.A1(n_1049),
.A2(n_152),
.B(n_153),
.Y(n_1052)
);

AOI221xp5_ASAP7_75t_L g1053 ( 
.A1(n_1052),
.A2(n_1050),
.B1(n_1051),
.B2(n_157),
.C(n_158),
.Y(n_1053)
);

AOI211xp5_ASAP7_75t_L g1054 ( 
.A1(n_1053),
.A2(n_155),
.B(n_156),
.C(n_159),
.Y(n_1054)
);


endmodule