module fake_jpeg_7464_n_95 (n_13, n_21, n_33, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_19, n_18, n_20, n_35, n_4, n_34, n_30, n_16, n_3, n_0, n_24, n_28, n_26, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_12, n_32, n_8, n_15, n_7, n_95);

input n_13;
input n_21;
input n_33;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_35;
input n_4;
input n_34;
input n_30;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_26;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_95;

wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_73;
wire n_59;
wire n_84;
wire n_65;
wire n_42;
wire n_49;
wire n_76;
wire n_38;
wire n_88;
wire n_74;
wire n_50;
wire n_57;
wire n_69;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_44;
wire n_75;
wire n_37;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_39;
wire n_72;
wire n_89;
wire n_56;
wire n_79;
wire n_67;
wire n_53;
wire n_91;
wire n_54;
wire n_93;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_62;
wire n_43;
wire n_82;

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_11),
.Y(n_37)
);

BUFx5_ASAP7_75t_L g38 ( 
.A(n_29),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_32),
.Y(n_39)
);

BUFx5_ASAP7_75t_L g40 ( 
.A(n_0),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_14),
.Y(n_41)
);

HB1xp67_ASAP7_75t_L g42 ( 
.A(n_13),
.Y(n_42)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_2),
.Y(n_43)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_19),
.Y(n_44)
);

INVxp33_ASAP7_75t_L g45 ( 
.A(n_36),
.Y(n_45)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_10),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_2),
.Y(n_47)
);

INVx4_ASAP7_75t_L g48 ( 
.A(n_23),
.Y(n_48)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_12),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_SL g50 ( 
.A(n_43),
.B(n_0),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_L g60 ( 
.A(n_50),
.B(n_3),
.Y(n_60)
);

INVx3_ASAP7_75t_L g51 ( 
.A(n_47),
.Y(n_51)
);

INVx4_ASAP7_75t_L g57 ( 
.A(n_51),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_37),
.B(n_1),
.Y(n_52)
);

BUFx12f_ASAP7_75t_L g53 ( 
.A(n_38),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_SL g54 ( 
.A(n_46),
.B(n_1),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_SL g64 ( 
.A(n_54),
.B(n_4),
.Y(n_64)
);

BUFx24_ASAP7_75t_L g55 ( 
.A(n_40),
.Y(n_55)
);

CKINVDCx20_ASAP7_75t_R g56 ( 
.A(n_49),
.Y(n_56)
);

AOI22xp33_ASAP7_75t_SL g58 ( 
.A1(n_55),
.A2(n_48),
.B1(n_47),
.B2(n_45),
.Y(n_58)
);

OAI22xp5_ASAP7_75t_L g77 ( 
.A1(n_58),
.A2(n_62),
.B1(n_69),
.B2(n_17),
.Y(n_77)
);

AOI21xp33_ASAP7_75t_L g59 ( 
.A1(n_53),
.A2(n_44),
.B(n_41),
.Y(n_59)
);

OR2x2_ASAP7_75t_L g72 ( 
.A(n_59),
.B(n_15),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_60),
.B(n_64),
.Y(n_74)
);

CKINVDCx20_ASAP7_75t_R g61 ( 
.A(n_52),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_61),
.B(n_66),
.Y(n_76)
);

OAI22xp5_ASAP7_75t_SL g62 ( 
.A1(n_51),
.A2(n_39),
.B1(n_42),
.B2(n_45),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_54),
.B(n_42),
.Y(n_63)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_63),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_54),
.B(n_5),
.Y(n_65)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_65),
.Y(n_81)
);

CKINVDCx12_ASAP7_75t_R g66 ( 
.A(n_56),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_54),
.B(n_6),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_L g75 ( 
.A(n_67),
.B(n_16),
.Y(n_75)
);

INVx5_ASAP7_75t_L g68 ( 
.A(n_51),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_68),
.B(n_70),
.Y(n_78)
);

AOI22xp33_ASAP7_75t_SL g69 ( 
.A1(n_51),
.A2(n_7),
.B1(n_8),
.B2(n_9),
.Y(n_69)
);

CKINVDCx20_ASAP7_75t_R g70 ( 
.A(n_52),
.Y(n_70)
);

INVx5_ASAP7_75t_L g71 ( 
.A(n_51),
.Y(n_71)
);

AOI22xp33_ASAP7_75t_SL g80 ( 
.A1(n_71),
.A2(n_20),
.B1(n_21),
.B2(n_22),
.Y(n_80)
);

AND2x2_ASAP7_75t_L g82 ( 
.A(n_72),
.B(n_75),
.Y(n_82)
);

AOI22xp33_ASAP7_75t_SL g83 ( 
.A1(n_77),
.A2(n_79),
.B1(n_80),
.B2(n_57),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g79 ( 
.A(n_64),
.B(n_18),
.Y(n_79)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_83),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_84),
.B(n_73),
.Y(n_85)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_85),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_L g87 ( 
.A(n_86),
.B(n_74),
.Y(n_87)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_87),
.Y(n_88)
);

XOR2xp5_ASAP7_75t_L g89 ( 
.A(n_88),
.B(n_76),
.Y(n_89)
);

MAJIxp5_ASAP7_75t_L g90 ( 
.A(n_89),
.B(n_81),
.C(n_78),
.Y(n_90)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_90),
.Y(n_91)
);

INVxp67_ASAP7_75t_L g92 ( 
.A(n_91),
.Y(n_92)
);

AOI322xp5_ASAP7_75t_L g93 ( 
.A1(n_92),
.A2(n_82),
.A3(n_25),
.B1(n_26),
.B2(n_27),
.C1(n_28),
.C2(n_30),
.Y(n_93)
);

OAI321xp33_ASAP7_75t_L g94 ( 
.A1(n_93),
.A2(n_24),
.A3(n_31),
.B1(n_33),
.B2(n_34),
.C(n_35),
.Y(n_94)
);

XOR2xp5_ASAP7_75t_L g95 ( 
.A(n_94),
.B(n_78),
.Y(n_95)
);


endmodule