module fake_ariane_1055_n_1722 (n_83, n_8, n_56, n_60, n_64, n_119, n_124, n_90, n_38, n_47, n_110, n_153, n_18, n_86, n_75, n_89, n_67, n_149, n_34, n_69, n_95, n_92, n_143, n_150, n_98, n_74, n_113, n_114, n_33, n_19, n_40, n_152, n_120, n_106, n_12, n_53, n_111, n_21, n_115, n_133, n_66, n_71, n_24, n_7, n_109, n_96, n_156, n_49, n_20, n_100, n_17, n_50, n_132, n_62, n_147, n_51, n_76, n_103, n_79, n_26, n_3, n_46, n_0, n_84, n_36, n_91, n_107, n_72, n_105, n_128, n_44, n_30, n_82, n_31, n_42, n_57, n_131, n_70, n_10, n_117, n_139, n_85, n_130, n_144, n_6, n_48, n_94, n_101, n_4, n_134, n_2, n_32, n_37, n_58, n_65, n_123, n_9, n_138, n_112, n_45, n_11, n_129, n_126, n_137, n_122, n_148, n_52, n_135, n_73, n_77, n_15, n_118, n_93, n_121, n_23, n_61, n_108, n_102, n_125, n_22, n_43, n_1, n_81, n_87, n_13, n_27, n_29, n_41, n_140, n_55, n_151, n_136, n_28, n_80, n_146, n_97, n_154, n_142, n_14, n_88, n_141, n_68, n_116, n_104, n_145, n_78, n_39, n_59, n_63, n_99, n_16, n_5, n_155, n_127, n_35, n_54, n_25, n_1722);

input n_83;
input n_8;
input n_56;
input n_60;
input n_64;
input n_119;
input n_124;
input n_90;
input n_38;
input n_47;
input n_110;
input n_153;
input n_18;
input n_86;
input n_75;
input n_89;
input n_67;
input n_149;
input n_34;
input n_69;
input n_95;
input n_92;
input n_143;
input n_150;
input n_98;
input n_74;
input n_113;
input n_114;
input n_33;
input n_19;
input n_40;
input n_152;
input n_120;
input n_106;
input n_12;
input n_53;
input n_111;
input n_21;
input n_115;
input n_133;
input n_66;
input n_71;
input n_24;
input n_7;
input n_109;
input n_96;
input n_156;
input n_49;
input n_20;
input n_100;
input n_17;
input n_50;
input n_132;
input n_62;
input n_147;
input n_51;
input n_76;
input n_103;
input n_79;
input n_26;
input n_3;
input n_46;
input n_0;
input n_84;
input n_36;
input n_91;
input n_107;
input n_72;
input n_105;
input n_128;
input n_44;
input n_30;
input n_82;
input n_31;
input n_42;
input n_57;
input n_131;
input n_70;
input n_10;
input n_117;
input n_139;
input n_85;
input n_130;
input n_144;
input n_6;
input n_48;
input n_94;
input n_101;
input n_4;
input n_134;
input n_2;
input n_32;
input n_37;
input n_58;
input n_65;
input n_123;
input n_9;
input n_138;
input n_112;
input n_45;
input n_11;
input n_129;
input n_126;
input n_137;
input n_122;
input n_148;
input n_52;
input n_135;
input n_73;
input n_77;
input n_15;
input n_118;
input n_93;
input n_121;
input n_23;
input n_61;
input n_108;
input n_102;
input n_125;
input n_22;
input n_43;
input n_1;
input n_81;
input n_87;
input n_13;
input n_27;
input n_29;
input n_41;
input n_140;
input n_55;
input n_151;
input n_136;
input n_28;
input n_80;
input n_146;
input n_97;
input n_154;
input n_142;
input n_14;
input n_88;
input n_141;
input n_68;
input n_116;
input n_104;
input n_145;
input n_78;
input n_39;
input n_59;
input n_63;
input n_99;
input n_16;
input n_5;
input n_155;
input n_127;
input n_35;
input n_54;
input n_25;

output n_1722;

wire n_913;
wire n_1681;
wire n_1486;
wire n_1507;
wire n_589;
wire n_1174;
wire n_1469;
wire n_691;
wire n_1353;
wire n_1355;
wire n_423;
wire n_1383;
wire n_603;
wire n_373;
wire n_1250;
wire n_1169;
wire n_789;
wire n_850;
wire n_610;
wire n_245;
wire n_1713;
wire n_319;
wire n_1436;
wire n_690;
wire n_416;
wire n_1109;
wire n_1430;
wire n_525;
wire n_187;
wire n_1463;
wire n_1238;
wire n_1515;
wire n_817;
wire n_924;
wire n_781;
wire n_1566;
wire n_189;
wire n_717;
wire n_952;
wire n_864;
wire n_1096;
wire n_1379;
wire n_1706;
wire n_524;
wire n_1214;
wire n_634;
wire n_1246;
wire n_1138;
wire n_214;
wire n_764;
wire n_1503;
wire n_462;
wire n_1196;
wire n_1181;
wire n_410;
wire n_1187;
wire n_1131;
wire n_1225;
wire n_737;
wire n_1298;
wire n_1366;
wire n_232;
wire n_568;
wire n_1088;
wire n_1424;
wire n_766;
wire n_1457;
wire n_377;
wire n_1682;
wire n_520;
wire n_870;
wire n_1453;
wire n_279;
wire n_945;
wire n_958;
wire n_813;
wire n_419;
wire n_270;
wire n_338;
wire n_995;
wire n_285;
wire n_1184;
wire n_202;
wire n_1535;
wire n_500;
wire n_754;
wire n_665;
wire n_903;
wire n_871;
wire n_1073;
wire n_239;
wire n_402;
wire n_1277;
wire n_829;
wire n_1062;
wire n_339;
wire n_738;
wire n_1690;
wire n_672;
wire n_740;
wire n_1283;
wire n_167;
wire n_1018;
wire n_259;
wire n_953;
wire n_1364;
wire n_1224;
wire n_1425;
wire n_625;
wire n_557;
wire n_1107;
wire n_1688;
wire n_989;
wire n_242;
wire n_645;
wire n_331;
wire n_559;
wire n_267;
wire n_495;
wire n_350;
wire n_381;
wire n_795;
wire n_721;
wire n_1084;
wire n_1718;
wire n_1276;
wire n_200;
wire n_1428;
wire n_1284;
wire n_1241;
wire n_821;
wire n_561;
wire n_770;
wire n_1514;
wire n_1528;
wire n_507;
wire n_486;
wire n_901;
wire n_569;
wire n_1145;
wire n_971;
wire n_787;
wire n_1650;
wire n_1519;
wire n_1195;
wire n_1522;
wire n_518;
wire n_1207;
wire n_222;
wire n_786;
wire n_1404;
wire n_868;
wire n_1542;
wire n_1314;
wire n_1512;
wire n_1539;
wire n_884;
wire n_1415;
wire n_1034;
wire n_1652;
wire n_1676;
wire n_1085;
wire n_277;
wire n_1636;
wire n_432;
wire n_293;
wire n_823;
wire n_620;
wire n_1074;
wire n_859;
wire n_587;
wire n_693;
wire n_863;
wire n_303;
wire n_1254;
wire n_929;
wire n_352;
wire n_206;
wire n_899;
wire n_1703;
wire n_611;
wire n_1295;
wire n_365;
wire n_238;
wire n_1013;
wire n_1495;
wire n_1637;
wire n_334;
wire n_192;
wire n_661;
wire n_300;
wire n_533;
wire n_438;
wire n_1560;
wire n_1654;
wire n_1548;
wire n_440;
wire n_273;
wire n_1396;
wire n_1230;
wire n_612;
wire n_333;
wire n_376;
wire n_512;
wire n_1597;
wire n_1544;
wire n_579;
wire n_844;
wire n_1012;
wire n_1267;
wire n_1354;
wire n_1213;
wire n_237;
wire n_780;
wire n_1021;
wire n_1443;
wire n_491;
wire n_1465;
wire n_1595;
wire n_1142;
wire n_1140;
wire n_705;
wire n_570;
wire n_260;
wire n_942;
wire n_1437;
wire n_1378;
wire n_461;
wire n_1121;
wire n_1416;
wire n_209;
wire n_490;
wire n_1461;
wire n_1391;
wire n_225;
wire n_1599;
wire n_1006;
wire n_575;
wire n_546;
wire n_503;
wire n_1112;
wire n_700;
wire n_1159;
wire n_772;
wire n_1216;
wire n_1245;
wire n_1669;
wire n_1675;
wire n_676;
wire n_1594;
wire n_680;
wire n_287;
wire n_1716;
wire n_302;
wire n_380;
wire n_1585;
wire n_1432;
wire n_249;
wire n_1108;
wire n_355;
wire n_212;
wire n_444;
wire n_851;
wire n_1590;
wire n_1351;
wire n_1274;
wire n_257;
wire n_652;
wire n_475;
wire n_947;
wire n_930;
wire n_1260;
wire n_1179;
wire n_468;
wire n_182;
wire n_696;
wire n_1442;
wire n_482;
wire n_798;
wire n_577;
wire n_407;
wire n_1691;
wire n_916;
wire n_1386;
wire n_912;
wire n_460;
wire n_1555;
wire n_366;
wire n_762;
wire n_1253;
wire n_1468;
wire n_1661;
wire n_555;
wire n_804;
wire n_1656;
wire n_1382;
wire n_992;
wire n_966;
wire n_955;
wire n_1182;
wire n_794;
wire n_1692;
wire n_1562;
wire n_514;
wire n_418;
wire n_1376;
wire n_513;
wire n_288;
wire n_179;
wire n_1292;
wire n_1178;
wire n_1435;
wire n_1026;
wire n_1506;
wire n_1610;
wire n_306;
wire n_203;
wire n_436;
wire n_324;
wire n_669;
wire n_931;
wire n_1491;
wire n_619;
wire n_337;
wire n_437;
wire n_274;
wire n_967;
wire n_1083;
wire n_1418;
wire n_746;
wire n_1357;
wire n_292;
wire n_1079;
wire n_1389;
wire n_615;
wire n_1139;
wire n_517;
wire n_1312;
wire n_1717;
wire n_824;
wire n_428;
wire n_159;
wire n_892;
wire n_959;
wire n_1399;
wire n_1101;
wire n_1567;
wire n_1343;
wire n_563;
wire n_990;
wire n_1623;
wire n_867;
wire n_1226;
wire n_944;
wire n_749;
wire n_815;
wire n_542;
wire n_1340;
wire n_470;
wire n_1240;
wire n_1087;
wire n_632;
wire n_477;
wire n_650;
wire n_425;
wire n_1433;
wire n_1155;
wire n_1071;
wire n_712;
wire n_976;
wire n_909;
wire n_1392;
wire n_767;
wire n_1680;
wire n_964;
wire n_1627;
wire n_382;
wire n_489;
wire n_251;
wire n_974;
wire n_506;
wire n_799;
wire n_1147;
wire n_397;
wire n_471;
wire n_351;
wire n_965;
wire n_934;
wire n_1447;
wire n_1220;
wire n_356;
wire n_698;
wire n_1674;
wire n_307;
wire n_1209;
wire n_1020;
wire n_1563;
wire n_646;
wire n_1633;
wire n_404;
wire n_172;
wire n_1058;
wire n_347;
wire n_1042;
wire n_183;
wire n_1234;
wire n_479;
wire n_1578;
wire n_1455;
wire n_299;
wire n_836;
wire n_1279;
wire n_564;
wire n_205;
wire n_1029;
wire n_1247;
wire n_760;
wire n_522;
wire n_1568;
wire n_1483;
wire n_1363;
wire n_367;
wire n_1111;
wire n_970;
wire n_1689;
wire n_713;
wire n_1255;
wire n_1646;
wire n_598;
wire n_345;
wire n_1237;
wire n_927;
wire n_261;
wire n_1095;
wire n_370;
wire n_706;
wire n_286;
wire n_1401;
wire n_1419;
wire n_1531;
wire n_776;
wire n_424;
wire n_1651;
wire n_1387;
wire n_466;
wire n_1263;
wire n_346;
wire n_348;
wire n_552;
wire n_670;
wire n_379;
wire n_162;
wire n_264;
wire n_441;
wire n_1032;
wire n_1217;
wire n_1496;
wire n_637;
wire n_1592;
wire n_327;
wire n_1259;
wire n_1177;
wire n_1231;
wire n_980;
wire n_1618;
wire n_905;
wire n_207;
wire n_720;
wire n_926;
wire n_194;
wire n_1163;
wire n_186;
wire n_1384;
wire n_1501;
wire n_1173;
wire n_1068;
wire n_1198;
wire n_1570;
wire n_487;
wire n_1518;
wire n_1456;
wire n_1648;
wire n_1413;
wire n_855;
wire n_158;
wire n_808;
wire n_1365;
wire n_553;
wire n_1439;
wire n_814;
wire n_578;
wire n_1665;
wire n_1287;
wire n_405;
wire n_1611;
wire n_320;
wire n_1414;
wire n_1134;
wire n_1484;
wire n_647;
wire n_1423;
wire n_481;
wire n_600;
wire n_1053;
wire n_1609;
wire n_529;
wire n_502;
wire n_218;
wire n_1467;
wire n_247;
wire n_1304;
wire n_1608;
wire n_1105;
wire n_547;
wire n_439;
wire n_604;
wire n_677;
wire n_478;
wire n_703;
wire n_1349;
wire n_1709;
wire n_1061;
wire n_326;
wire n_681;
wire n_227;
wire n_874;
wire n_1278;
wire n_707;
wire n_983;
wire n_590;
wire n_699;
wire n_727;
wire n_301;
wire n_545;
wire n_1015;
wire n_1377;
wire n_1162;
wire n_536;
wire n_1614;
wire n_325;
wire n_1602;
wire n_688;
wire n_636;
wire n_427;
wire n_1098;
wire n_1490;
wire n_442;
wire n_777;
wire n_1553;
wire n_1080;
wire n_920;
wire n_1086;
wire n_1092;
wire n_986;
wire n_1104;
wire n_729;
wire n_887;
wire n_1122;
wire n_1205;
wire n_1408;
wire n_163;
wire n_1693;
wire n_1132;
wire n_390;
wire n_1156;
wire n_501;
wire n_314;
wire n_1120;
wire n_1202;
wire n_627;
wire n_1188;
wire n_1498;
wire n_1371;
wire n_233;
wire n_957;
wire n_388;
wire n_1402;
wire n_1242;
wire n_1607;
wire n_1489;
wire n_1218;
wire n_321;
wire n_221;
wire n_1586;
wire n_861;
wire n_1543;
wire n_1431;
wire n_877;
wire n_1119;
wire n_1666;
wire n_1500;
wire n_616;
wire n_1055;
wire n_1395;
wire n_1346;
wire n_1189;
wire n_1089;
wire n_281;
wire n_262;
wire n_1502;
wire n_1523;
wire n_1478;
wire n_735;
wire n_297;
wire n_1005;
wire n_527;
wire n_1294;
wire n_1667;
wire n_888;
wire n_845;
wire n_1649;
wire n_1677;
wire n_1297;
wire n_178;
wire n_551;
wire n_417;
wire n_1708;
wire n_343;
wire n_1222;
wire n_582;
wire n_755;
wire n_1097;
wire n_1219;
wire n_1711;
wire n_710;
wire n_534;
wire n_1460;
wire n_1239;
wire n_278;
wire n_560;
wire n_890;
wire n_842;
wire n_451;
wire n_745;
wire n_1572;
wire n_742;
wire n_1081;
wire n_1373;
wire n_1388;
wire n_1266;
wire n_1540;
wire n_1719;
wire n_769;
wire n_1372;
wire n_476;
wire n_832;
wire n_535;
wire n_744;
wire n_982;
wire n_915;
wire n_215;
wire n_1075;
wire n_454;
wire n_298;
wire n_1331;
wire n_1529;
wire n_1227;
wire n_655;
wire n_403;
wire n_1007;
wire n_1580;
wire n_1319;
wire n_657;
wire n_837;
wire n_812;
wire n_606;
wire n_951;
wire n_862;
wire n_1700;
wire n_659;
wire n_1332;
wire n_509;
wire n_666;
wire n_430;
wire n_1206;
wire n_722;
wire n_1508;
wire n_1532;
wire n_1171;
wire n_1030;
wire n_785;
wire n_1309;
wire n_999;
wire n_1338;
wire n_1342;
wire n_456;
wire n_852;
wire n_1394;
wire n_704;
wire n_1060;
wire n_1044;
wire n_1714;
wire n_521;
wire n_873;
wire n_1301;
wire n_1243;
wire n_1400;
wire n_342;
wire n_1466;
wire n_1513;
wire n_1527;
wire n_358;
wire n_608;
wire n_1538;
wire n_1037;
wire n_1329;
wire n_317;
wire n_1545;
wire n_1257;
wire n_1480;
wire n_1668;
wire n_1605;
wire n_1078;
wire n_266;
wire n_157;
wire n_1161;
wire n_811;
wire n_624;
wire n_791;
wire n_876;
wire n_618;
wire n_1191;
wire n_736;
wire n_1025;
wire n_1215;
wire n_241;
wire n_1449;
wire n_687;
wire n_797;
wire n_480;
wire n_1327;
wire n_1475;
wire n_211;
wire n_642;
wire n_408;
wire n_1406;
wire n_595;
wire n_1405;
wire n_602;
wire n_592;
wire n_1499;
wire n_854;
wire n_1318;
wire n_393;
wire n_1632;
wire n_474;
wire n_805;
wire n_295;
wire n_1658;
wire n_190;
wire n_1072;
wire n_695;
wire n_1526;
wire n_1305;
wire n_180;
wire n_730;
wire n_386;
wire n_1596;
wire n_1281;
wire n_516;
wire n_1137;
wire n_1258;
wire n_197;
wire n_640;
wire n_463;
wire n_1476;
wire n_1524;
wire n_943;
wire n_1118;
wire n_678;
wire n_651;
wire n_1293;
wire n_961;
wire n_469;
wire n_1046;
wire n_726;
wire n_1123;
wire n_1657;
wire n_878;
wire n_771;
wire n_1321;
wire n_752;
wire n_1488;
wire n_985;
wire n_421;
wire n_1330;
wire n_906;
wire n_1180;
wire n_1697;
wire n_283;
wire n_806;
wire n_1350;
wire n_1556;
wire n_649;
wire n_1561;
wire n_374;
wire n_1352;
wire n_643;
wire n_1492;
wire n_226;
wire n_1441;
wire n_682;
wire n_1616;
wire n_819;
wire n_586;
wire n_1324;
wire n_1429;
wire n_686;
wire n_605;
wire n_1154;
wire n_584;
wire n_1557;
wire n_1130;
wire n_1450;
wire n_349;
wire n_756;
wire n_1016;
wire n_1149;
wire n_1505;
wire n_979;
wire n_1642;
wire n_897;
wire n_949;
wire n_1493;
wire n_515;
wire n_807;
wire n_891;
wire n_885;
wire n_1659;
wire n_198;
wire n_1208;
wire n_396;
wire n_802;
wire n_1151;
wire n_554;
wire n_960;
wire n_1256;
wire n_714;
wire n_790;
wire n_354;
wire n_725;
wire n_1577;
wire n_1448;
wire n_1009;
wire n_230;
wire n_1133;
wire n_883;
wire n_473;
wire n_801;
wire n_1286;
wire n_818;
wire n_1685;
wire n_779;
wire n_594;
wire n_1397;
wire n_1052;
wire n_272;
wire n_1333;
wire n_1306;
wire n_833;
wire n_1426;
wire n_879;
wire n_1117;
wire n_422;
wire n_1269;
wire n_1303;
wire n_1547;
wire n_1438;
wire n_1541;
wire n_597;
wire n_1047;
wire n_1472;
wire n_1593;
wire n_1050;
wire n_566;
wire n_169;
wire n_1201;
wire n_1288;
wire n_173;
wire n_858;
wire n_1185;
wire n_335;
wire n_1035;
wire n_1143;
wire n_344;
wire n_426;
wire n_433;
wire n_398;
wire n_210;
wire n_1090;
wire n_1367;
wire n_166;
wire n_253;
wire n_928;
wire n_1153;
wire n_271;
wire n_465;
wire n_825;
wire n_1103;
wire n_732;
wire n_1565;
wire n_1192;
wire n_224;
wire n_894;
wire n_1380;
wire n_1624;
wire n_420;
wire n_1291;
wire n_562;
wire n_748;
wire n_510;
wire n_1045;
wire n_256;
wire n_1160;
wire n_1023;
wire n_988;
wire n_330;
wire n_914;
wire n_400;
wire n_689;
wire n_1116;
wire n_282;
wire n_328;
wire n_368;
wire n_467;
wire n_1511;
wire n_1422;
wire n_644;
wire n_1197;
wire n_276;
wire n_497;
wire n_1165;
wire n_1641;
wire n_168;
wire n_538;
wire n_1517;
wire n_576;
wire n_843;
wire n_511;
wire n_455;
wire n_429;
wire n_588;
wire n_638;
wire n_1307;
wire n_1128;
wire n_1671;
wire n_1417;
wire n_1048;
wire n_775;
wire n_667;
wire n_1049;
wire n_869;
wire n_846;
wire n_1398;
wire n_1356;
wire n_1341;
wire n_1504;
wire n_1440;
wire n_1370;
wire n_1603;
wire n_305;
wire n_312;
wire n_728;
wire n_413;
wire n_715;
wire n_889;
wire n_1066;
wire n_1549;
wire n_935;
wire n_685;
wire n_911;
wire n_361;
wire n_623;
wire n_1712;
wire n_1403;
wire n_1065;
wire n_453;
wire n_1534;
wire n_810;
wire n_1290;
wire n_181;
wire n_617;
wire n_543;
wire n_1362;
wire n_1559;
wire n_236;
wire n_683;
wire n_601;
wire n_565;
wire n_628;
wire n_1300;
wire n_743;
wire n_1194;
wire n_1647;
wire n_1546;
wire n_1420;
wire n_907;
wire n_1454;
wire n_660;
wire n_464;
wire n_962;
wire n_941;
wire n_1210;
wire n_847;
wire n_747;
wire n_1622;
wire n_1135;
wire n_918;
wire n_639;
wire n_452;
wire n_673;
wire n_1038;
wire n_414;
wire n_571;
wire n_1521;
wire n_1694;
wire n_284;
wire n_593;
wire n_1695;
wire n_1164;
wire n_609;
wire n_1193;
wire n_1345;
wire n_613;
wire n_1022;
wire n_1336;
wire n_1033;
wire n_409;
wire n_171;
wire n_519;
wire n_384;
wire n_1166;
wire n_1056;
wire n_526;
wire n_1040;
wire n_674;
wire n_1158;
wire n_316;
wire n_1444;
wire n_820;
wire n_872;
wire n_1653;
wire n_254;
wire n_1157;
wire n_1584;
wire n_234;
wire n_848;
wire n_1664;
wire n_280;
wire n_629;
wire n_161;
wire n_532;
wire n_763;
wire n_540;
wire n_216;
wire n_692;
wire n_984;
wire n_1687;
wire n_223;
wire n_1552;
wire n_750;
wire n_834;
wire n_1612;
wire n_800;
wire n_1606;
wire n_395;
wire n_621;
wire n_1587;
wire n_213;
wire n_1014;
wire n_724;
wire n_1427;
wire n_1481;
wire n_493;
wire n_1311;
wire n_1589;
wire n_1100;
wire n_585;
wire n_875;
wire n_1617;
wire n_827;
wire n_697;
wire n_622;
wire n_1626;
wire n_1335;
wire n_1715;
wire n_296;
wire n_880;
wire n_793;
wire n_1175;
wire n_751;
wire n_1027;
wire n_1070;
wire n_1621;
wire n_739;
wire n_1485;
wire n_1028;
wire n_1221;
wire n_530;
wire n_792;
wire n_1262;
wire n_580;
wire n_1579;
wire n_494;
wire n_434;
wire n_975;
wire n_229;
wire n_394;
wire n_923;
wire n_1645;
wire n_1124;
wire n_1381;
wire n_1494;
wire n_932;
wire n_1183;
wire n_1326;
wire n_981;
wire n_1110;
wire n_243;
wire n_1407;
wire n_185;
wire n_1204;
wire n_1554;
wire n_994;
wire n_1360;
wire n_973;
wire n_268;
wire n_972;
wire n_164;
wire n_184;
wire n_856;
wire n_1248;
wire n_1176;
wire n_1564;
wire n_1054;
wire n_508;
wire n_1679;
wire n_353;
wire n_1678;
wire n_1482;
wire n_1361;
wire n_1601;
wire n_1057;
wire n_191;
wire n_1011;
wire n_978;
wire n_1520;
wire n_1509;
wire n_828;
wire n_322;
wire n_1411;
wire n_1359;
wire n_558;
wire n_1721;
wire n_653;
wire n_1445;
wire n_1317;
wire n_783;
wire n_556;
wire n_1127;
wire n_170;
wire n_1536;
wire n_1471;
wire n_160;
wire n_1008;
wire n_332;
wire n_581;
wire n_294;
wire n_1024;
wire n_830;
wire n_176;
wire n_987;
wire n_936;
wire n_1620;
wire n_1385;
wire n_1525;
wire n_541;
wire n_499;
wire n_788;
wire n_908;
wire n_1036;
wire n_341;
wire n_1270;
wire n_1167;
wire n_1272;
wire n_549;
wire n_591;
wire n_969;
wire n_919;
wire n_1663;
wire n_1625;
wire n_318;
wire n_1458;
wire n_244;
wire n_679;
wire n_1630;
wire n_220;
wire n_663;
wire n_1720;
wire n_443;
wire n_1412;
wire n_1550;
wire n_528;
wire n_1358;
wire n_1200;
wire n_387;
wire n_406;
wire n_826;
wire n_391;
wire n_940;
wire n_1537;
wire n_1077;
wire n_607;
wire n_956;
wire n_445;
wire n_765;
wire n_1268;
wire n_385;
wire n_917;
wire n_1271;
wire n_372;
wire n_1530;
wire n_631;
wire n_399;
wire n_1170;
wire n_1261;
wire n_702;
wire n_898;
wire n_857;
wire n_363;
wire n_968;
wire n_1067;
wire n_1235;
wire n_1323;
wire n_1462;
wire n_1064;
wire n_633;
wire n_900;
wire n_1446;
wire n_1282;
wire n_1701;
wire n_1093;
wire n_1551;
wire n_1285;
wire n_193;
wire n_761;
wire n_733;
wire n_731;
wire n_336;
wire n_315;
wire n_311;
wire n_1452;
wire n_1573;
wire n_668;
wire n_758;
wire n_1106;
wire n_648;
wire n_784;
wire n_269;
wire n_816;
wire n_1322;
wire n_1473;
wire n_835;
wire n_446;
wire n_1076;
wire n_1348;
wire n_753;
wire n_701;
wire n_1003;
wire n_1125;
wire n_1710;
wire n_309;
wire n_1344;
wire n_1390;
wire n_401;
wire n_485;
wire n_504;
wire n_483;
wire n_435;
wire n_1141;
wire n_1629;
wire n_291;
wire n_1640;
wire n_822;
wire n_1094;
wire n_840;
wire n_1459;
wire n_1510;
wire n_1099;
wire n_839;
wire n_759;
wire n_567;
wire n_369;
wire n_240;
wire n_1575;
wire n_1172;
wire n_614;
wire n_1212;
wire n_831;
wire n_778;
wire n_1619;
wire n_188;
wire n_323;
wire n_550;
wire n_1315;
wire n_1660;
wire n_997;
wire n_635;
wire n_694;
wire n_1643;
wire n_1320;
wire n_1113;
wire n_248;
wire n_1152;
wire n_921;
wire n_1615;
wire n_1236;
wire n_228;
wire n_1265;
wire n_1576;
wire n_1470;
wire n_671;
wire n_1533;
wire n_1409;
wire n_1148;
wire n_1588;
wire n_1684;
wire n_1673;
wire n_1334;
wire n_654;
wire n_1275;
wire n_488;
wire n_904;
wire n_505;
wire n_1696;
wire n_498;
wire n_1059;
wire n_684;
wire n_1039;
wire n_539;
wire n_1150;
wire n_977;
wire n_449;
wire n_392;
wire n_1628;
wire n_1289;
wire n_1497;
wire n_459;
wire n_1136;
wire n_458;
wire n_1190;
wire n_1600;
wire n_1144;
wire n_383;
wire n_838;
wire n_1558;
wire n_1316;
wire n_175;
wire n_950;
wire n_1017;
wire n_711;
wire n_734;
wire n_723;
wire n_1393;
wire n_658;
wire n_630;
wire n_1369;
wire n_362;
wire n_310;
wire n_709;
wire n_809;
wire n_1686;
wire n_235;
wire n_881;
wire n_1019;
wire n_1477;
wire n_662;
wire n_641;
wire n_910;
wire n_290;
wire n_741;
wire n_939;
wire n_1410;
wire n_371;
wire n_199;
wire n_217;
wire n_1114;
wire n_1325;
wire n_708;
wire n_308;
wire n_1223;
wire n_201;
wire n_572;
wire n_1199;
wire n_865;
wire n_1273;
wire n_1041;
wire n_993;
wire n_948;
wire n_922;
wire n_1004;
wire n_448;
wire n_1347;
wire n_860;
wire n_1043;
wire n_255;
wire n_450;
wire n_896;
wire n_1479;
wire n_1613;
wire n_902;
wire n_1031;
wire n_1638;
wire n_853;
wire n_716;
wire n_1571;
wire n_1698;
wire n_196;
wire n_1337;
wire n_774;
wire n_933;
wire n_596;
wire n_954;
wire n_1168;
wire n_219;
wire n_1310;
wire n_231;
wire n_656;
wire n_492;
wire n_574;
wire n_252;
wire n_664;
wire n_1591;
wire n_1229;
wire n_1683;
wire n_415;
wire n_1280;
wire n_544;
wire n_1516;
wire n_1186;
wire n_1705;
wire n_599;
wire n_768;
wire n_1091;
wire n_537;
wire n_1063;
wire n_991;
wire n_389;
wire n_1670;
wire n_1707;
wire n_1126;
wire n_195;
wire n_938;
wire n_1328;
wire n_895;
wire n_304;
wire n_1639;
wire n_583;
wire n_1302;
wire n_1000;
wire n_313;
wire n_626;
wire n_378;
wire n_1581;
wire n_946;
wire n_757;
wire n_375;
wire n_1655;
wire n_1146;
wire n_1634;
wire n_1203;
wire n_998;
wire n_1699;
wire n_1598;
wire n_472;
wire n_937;
wire n_1474;
wire n_265;
wire n_1583;
wire n_1604;
wire n_208;
wire n_1631;
wire n_1702;
wire n_174;
wire n_275;
wire n_1375;
wire n_204;
wire n_1232;
wire n_996;
wire n_1211;
wire n_1368;
wire n_963;
wire n_1264;
wire n_1082;
wire n_496;
wire n_866;
wire n_246;
wire n_925;
wire n_1313;
wire n_1001;
wire n_1115;
wire n_1339;
wire n_1002;
wire n_1644;
wire n_1051;
wire n_719;
wire n_263;
wire n_1102;
wire n_360;
wire n_1129;
wire n_1252;
wire n_250;
wire n_1464;
wire n_1296;
wire n_773;
wire n_165;
wire n_1010;
wire n_882;
wire n_1249;
wire n_803;
wire n_329;
wire n_718;
wire n_1434;
wire n_340;
wire n_1569;
wire n_289;
wire n_548;
wire n_523;
wire n_1662;
wire n_457;
wire n_1299;
wire n_177;
wire n_782;
wire n_364;
wire n_258;
wire n_431;
wire n_1228;
wire n_1244;
wire n_411;
wire n_484;
wire n_849;
wire n_357;
wire n_412;
wire n_1251;
wire n_447;
wire n_1421;
wire n_1233;
wire n_1574;
wire n_1672;
wire n_1635;
wire n_1704;
wire n_893;
wire n_1582;
wire n_841;
wire n_886;
wire n_1069;
wire n_359;
wire n_1308;
wire n_573;
wire n_796;
wire n_531;
wire n_1374;
wire n_1451;
wire n_1487;
wire n_675;

INVx1_ASAP7_75t_L g157 ( 
.A(n_37),
.Y(n_157)
);

CKINVDCx5p33_ASAP7_75t_R g158 ( 
.A(n_17),
.Y(n_158)
);

INVx2_ASAP7_75t_L g159 ( 
.A(n_49),
.Y(n_159)
);

BUFx3_ASAP7_75t_L g160 ( 
.A(n_60),
.Y(n_160)
);

CKINVDCx5p33_ASAP7_75t_R g161 ( 
.A(n_30),
.Y(n_161)
);

CKINVDCx20_ASAP7_75t_R g162 ( 
.A(n_37),
.Y(n_162)
);

CKINVDCx16_ASAP7_75t_R g163 ( 
.A(n_10),
.Y(n_163)
);

CKINVDCx5p33_ASAP7_75t_R g164 ( 
.A(n_94),
.Y(n_164)
);

CKINVDCx5p33_ASAP7_75t_R g165 ( 
.A(n_118),
.Y(n_165)
);

CKINVDCx5p33_ASAP7_75t_R g166 ( 
.A(n_76),
.Y(n_166)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_133),
.Y(n_167)
);

CKINVDCx5p33_ASAP7_75t_R g168 ( 
.A(n_48),
.Y(n_168)
);

CKINVDCx5p33_ASAP7_75t_R g169 ( 
.A(n_122),
.Y(n_169)
);

CKINVDCx5p33_ASAP7_75t_R g170 ( 
.A(n_29),
.Y(n_170)
);

CKINVDCx20_ASAP7_75t_R g171 ( 
.A(n_25),
.Y(n_171)
);

HB1xp67_ASAP7_75t_L g172 ( 
.A(n_18),
.Y(n_172)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_78),
.Y(n_173)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_85),
.Y(n_174)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_17),
.Y(n_175)
);

CKINVDCx5p33_ASAP7_75t_R g176 ( 
.A(n_145),
.Y(n_176)
);

CKINVDCx5p33_ASAP7_75t_R g177 ( 
.A(n_30),
.Y(n_177)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_123),
.Y(n_178)
);

CKINVDCx5p33_ASAP7_75t_R g179 ( 
.A(n_38),
.Y(n_179)
);

CKINVDCx5p33_ASAP7_75t_R g180 ( 
.A(n_32),
.Y(n_180)
);

CKINVDCx5p33_ASAP7_75t_R g181 ( 
.A(n_46),
.Y(n_181)
);

CKINVDCx5p33_ASAP7_75t_R g182 ( 
.A(n_147),
.Y(n_182)
);

CKINVDCx5p33_ASAP7_75t_R g183 ( 
.A(n_137),
.Y(n_183)
);

CKINVDCx5p33_ASAP7_75t_R g184 ( 
.A(n_126),
.Y(n_184)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_150),
.Y(n_185)
);

CKINVDCx5p33_ASAP7_75t_R g186 ( 
.A(n_72),
.Y(n_186)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_18),
.Y(n_187)
);

CKINVDCx20_ASAP7_75t_R g188 ( 
.A(n_24),
.Y(n_188)
);

CKINVDCx5p33_ASAP7_75t_R g189 ( 
.A(n_36),
.Y(n_189)
);

CKINVDCx5p33_ASAP7_75t_R g190 ( 
.A(n_25),
.Y(n_190)
);

CKINVDCx20_ASAP7_75t_R g191 ( 
.A(n_7),
.Y(n_191)
);

BUFx3_ASAP7_75t_L g192 ( 
.A(n_21),
.Y(n_192)
);

CKINVDCx5p33_ASAP7_75t_R g193 ( 
.A(n_61),
.Y(n_193)
);

CKINVDCx5p33_ASAP7_75t_R g194 ( 
.A(n_66),
.Y(n_194)
);

CKINVDCx5p33_ASAP7_75t_R g195 ( 
.A(n_132),
.Y(n_195)
);

CKINVDCx5p33_ASAP7_75t_R g196 ( 
.A(n_121),
.Y(n_196)
);

CKINVDCx5p33_ASAP7_75t_R g197 ( 
.A(n_105),
.Y(n_197)
);

CKINVDCx5p33_ASAP7_75t_R g198 ( 
.A(n_127),
.Y(n_198)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_97),
.Y(n_199)
);

INVx2_ASAP7_75t_L g200 ( 
.A(n_44),
.Y(n_200)
);

CKINVDCx5p33_ASAP7_75t_R g201 ( 
.A(n_31),
.Y(n_201)
);

CKINVDCx5p33_ASAP7_75t_R g202 ( 
.A(n_146),
.Y(n_202)
);

CKINVDCx5p33_ASAP7_75t_R g203 ( 
.A(n_59),
.Y(n_203)
);

CKINVDCx5p33_ASAP7_75t_R g204 ( 
.A(n_80),
.Y(n_204)
);

CKINVDCx5p33_ASAP7_75t_R g205 ( 
.A(n_138),
.Y(n_205)
);

CKINVDCx5p33_ASAP7_75t_R g206 ( 
.A(n_87),
.Y(n_206)
);

CKINVDCx5p33_ASAP7_75t_R g207 ( 
.A(n_141),
.Y(n_207)
);

INVx1_ASAP7_75t_SL g208 ( 
.A(n_53),
.Y(n_208)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_98),
.Y(n_209)
);

BUFx3_ASAP7_75t_L g210 ( 
.A(n_41),
.Y(n_210)
);

CKINVDCx5p33_ASAP7_75t_R g211 ( 
.A(n_108),
.Y(n_211)
);

CKINVDCx20_ASAP7_75t_R g212 ( 
.A(n_142),
.Y(n_212)
);

INVxp33_ASAP7_75t_L g213 ( 
.A(n_13),
.Y(n_213)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_9),
.Y(n_214)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_88),
.Y(n_215)
);

CKINVDCx20_ASAP7_75t_R g216 ( 
.A(n_111),
.Y(n_216)
);

INVx1_ASAP7_75t_SL g217 ( 
.A(n_117),
.Y(n_217)
);

CKINVDCx5p33_ASAP7_75t_R g218 ( 
.A(n_129),
.Y(n_218)
);

CKINVDCx5p33_ASAP7_75t_R g219 ( 
.A(n_48),
.Y(n_219)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_9),
.Y(n_220)
);

BUFx3_ASAP7_75t_L g221 ( 
.A(n_135),
.Y(n_221)
);

CKINVDCx5p33_ASAP7_75t_R g222 ( 
.A(n_54),
.Y(n_222)
);

CKINVDCx5p33_ASAP7_75t_R g223 ( 
.A(n_23),
.Y(n_223)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_54),
.Y(n_224)
);

CKINVDCx5p33_ASAP7_75t_R g225 ( 
.A(n_45),
.Y(n_225)
);

CKINVDCx5p33_ASAP7_75t_R g226 ( 
.A(n_22),
.Y(n_226)
);

CKINVDCx5p33_ASAP7_75t_R g227 ( 
.A(n_53),
.Y(n_227)
);

BUFx10_ASAP7_75t_L g228 ( 
.A(n_45),
.Y(n_228)
);

CKINVDCx5p33_ASAP7_75t_R g229 ( 
.A(n_51),
.Y(n_229)
);

CKINVDCx5p33_ASAP7_75t_R g230 ( 
.A(n_62),
.Y(n_230)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_39),
.Y(n_231)
);

CKINVDCx5p33_ASAP7_75t_R g232 ( 
.A(n_134),
.Y(n_232)
);

CKINVDCx5p33_ASAP7_75t_R g233 ( 
.A(n_130),
.Y(n_233)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_99),
.Y(n_234)
);

CKINVDCx5p33_ASAP7_75t_R g235 ( 
.A(n_4),
.Y(n_235)
);

INVx2_ASAP7_75t_L g236 ( 
.A(n_41),
.Y(n_236)
);

HB1xp67_ASAP7_75t_L g237 ( 
.A(n_93),
.Y(n_237)
);

CKINVDCx5p33_ASAP7_75t_R g238 ( 
.A(n_81),
.Y(n_238)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_31),
.Y(n_239)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_50),
.Y(n_240)
);

CKINVDCx5p33_ASAP7_75t_R g241 ( 
.A(n_35),
.Y(n_241)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_153),
.Y(n_242)
);

CKINVDCx5p33_ASAP7_75t_R g243 ( 
.A(n_35),
.Y(n_243)
);

CKINVDCx5p33_ASAP7_75t_R g244 ( 
.A(n_149),
.Y(n_244)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_82),
.Y(n_245)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_2),
.Y(n_246)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_3),
.Y(n_247)
);

CKINVDCx5p33_ASAP7_75t_R g248 ( 
.A(n_11),
.Y(n_248)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_131),
.Y(n_249)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_46),
.Y(n_250)
);

CKINVDCx20_ASAP7_75t_R g251 ( 
.A(n_75),
.Y(n_251)
);

CKINVDCx5p33_ASAP7_75t_R g252 ( 
.A(n_32),
.Y(n_252)
);

CKINVDCx5p33_ASAP7_75t_R g253 ( 
.A(n_42),
.Y(n_253)
);

CKINVDCx20_ASAP7_75t_R g254 ( 
.A(n_79),
.Y(n_254)
);

CKINVDCx5p33_ASAP7_75t_R g255 ( 
.A(n_110),
.Y(n_255)
);

CKINVDCx5p33_ASAP7_75t_R g256 ( 
.A(n_63),
.Y(n_256)
);

CKINVDCx5p33_ASAP7_75t_R g257 ( 
.A(n_128),
.Y(n_257)
);

INVx2_ASAP7_75t_L g258 ( 
.A(n_33),
.Y(n_258)
);

CKINVDCx5p33_ASAP7_75t_R g259 ( 
.A(n_143),
.Y(n_259)
);

CKINVDCx20_ASAP7_75t_R g260 ( 
.A(n_64),
.Y(n_260)
);

CKINVDCx5p33_ASAP7_75t_R g261 ( 
.A(n_34),
.Y(n_261)
);

CKINVDCx5p33_ASAP7_75t_R g262 ( 
.A(n_100),
.Y(n_262)
);

CKINVDCx5p33_ASAP7_75t_R g263 ( 
.A(n_43),
.Y(n_263)
);

BUFx3_ASAP7_75t_L g264 ( 
.A(n_70),
.Y(n_264)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_5),
.Y(n_265)
);

CKINVDCx5p33_ASAP7_75t_R g266 ( 
.A(n_90),
.Y(n_266)
);

CKINVDCx5p33_ASAP7_75t_R g267 ( 
.A(n_120),
.Y(n_267)
);

INVx2_ASAP7_75t_L g268 ( 
.A(n_52),
.Y(n_268)
);

CKINVDCx5p33_ASAP7_75t_R g269 ( 
.A(n_22),
.Y(n_269)
);

CKINVDCx20_ASAP7_75t_R g270 ( 
.A(n_67),
.Y(n_270)
);

CKINVDCx5p33_ASAP7_75t_R g271 ( 
.A(n_109),
.Y(n_271)
);

CKINVDCx5p33_ASAP7_75t_R g272 ( 
.A(n_77),
.Y(n_272)
);

CKINVDCx5p33_ASAP7_75t_R g273 ( 
.A(n_2),
.Y(n_273)
);

CKINVDCx16_ASAP7_75t_R g274 ( 
.A(n_95),
.Y(n_274)
);

INVx2_ASAP7_75t_L g275 ( 
.A(n_19),
.Y(n_275)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_3),
.Y(n_276)
);

CKINVDCx20_ASAP7_75t_R g277 ( 
.A(n_27),
.Y(n_277)
);

CKINVDCx11_ASAP7_75t_R g278 ( 
.A(n_27),
.Y(n_278)
);

INVx1_ASAP7_75t_SL g279 ( 
.A(n_155),
.Y(n_279)
);

CKINVDCx5p33_ASAP7_75t_R g280 ( 
.A(n_50),
.Y(n_280)
);

CKINVDCx5p33_ASAP7_75t_R g281 ( 
.A(n_116),
.Y(n_281)
);

CKINVDCx5p33_ASAP7_75t_R g282 ( 
.A(n_56),
.Y(n_282)
);

BUFx6f_ASAP7_75t_L g283 ( 
.A(n_36),
.Y(n_283)
);

INVx4_ASAP7_75t_R g284 ( 
.A(n_104),
.Y(n_284)
);

BUFx5_ASAP7_75t_L g285 ( 
.A(n_39),
.Y(n_285)
);

CKINVDCx5p33_ASAP7_75t_R g286 ( 
.A(n_52),
.Y(n_286)
);

CKINVDCx5p33_ASAP7_75t_R g287 ( 
.A(n_89),
.Y(n_287)
);

CKINVDCx16_ASAP7_75t_R g288 ( 
.A(n_8),
.Y(n_288)
);

CKINVDCx5p33_ASAP7_75t_R g289 ( 
.A(n_34),
.Y(n_289)
);

BUFx6f_ASAP7_75t_L g290 ( 
.A(n_83),
.Y(n_290)
);

CKINVDCx5p33_ASAP7_75t_R g291 ( 
.A(n_4),
.Y(n_291)
);

CKINVDCx5p33_ASAP7_75t_R g292 ( 
.A(n_152),
.Y(n_292)
);

CKINVDCx5p33_ASAP7_75t_R g293 ( 
.A(n_101),
.Y(n_293)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_1),
.Y(n_294)
);

CKINVDCx5p33_ASAP7_75t_R g295 ( 
.A(n_24),
.Y(n_295)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_28),
.Y(n_296)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_114),
.Y(n_297)
);

BUFx6f_ASAP7_75t_L g298 ( 
.A(n_144),
.Y(n_298)
);

CKINVDCx5p33_ASAP7_75t_R g299 ( 
.A(n_29),
.Y(n_299)
);

CKINVDCx5p33_ASAP7_75t_R g300 ( 
.A(n_10),
.Y(n_300)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_119),
.Y(n_301)
);

INVx2_ASAP7_75t_L g302 ( 
.A(n_40),
.Y(n_302)
);

CKINVDCx5p33_ASAP7_75t_R g303 ( 
.A(n_43),
.Y(n_303)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_21),
.Y(n_304)
);

CKINVDCx20_ASAP7_75t_R g305 ( 
.A(n_65),
.Y(n_305)
);

CKINVDCx5p33_ASAP7_75t_R g306 ( 
.A(n_136),
.Y(n_306)
);

CKINVDCx20_ASAP7_75t_R g307 ( 
.A(n_154),
.Y(n_307)
);

CKINVDCx5p33_ASAP7_75t_R g308 ( 
.A(n_26),
.Y(n_308)
);

CKINVDCx5p33_ASAP7_75t_R g309 ( 
.A(n_151),
.Y(n_309)
);

BUFx3_ASAP7_75t_L g310 ( 
.A(n_13),
.Y(n_310)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_156),
.Y(n_311)
);

CKINVDCx20_ASAP7_75t_R g312 ( 
.A(n_278),
.Y(n_312)
);

INVxp67_ASAP7_75t_SL g313 ( 
.A(n_157),
.Y(n_313)
);

NAND2xp5_ASAP7_75t_L g314 ( 
.A(n_285),
.B(n_0),
.Y(n_314)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_285),
.Y(n_315)
);

NOR2xp33_ASAP7_75t_L g316 ( 
.A(n_213),
.B(n_0),
.Y(n_316)
);

INVxp33_ASAP7_75t_SL g317 ( 
.A(n_172),
.Y(n_317)
);

INVxp67_ASAP7_75t_L g318 ( 
.A(n_159),
.Y(n_318)
);

INVx2_ASAP7_75t_L g319 ( 
.A(n_285),
.Y(n_319)
);

AND2x2_ASAP7_75t_L g320 ( 
.A(n_163),
.B(n_288),
.Y(n_320)
);

INVxp33_ASAP7_75t_SL g321 ( 
.A(n_158),
.Y(n_321)
);

CKINVDCx20_ASAP7_75t_R g322 ( 
.A(n_212),
.Y(n_322)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_285),
.Y(n_323)
);

CKINVDCx5p33_ASAP7_75t_R g324 ( 
.A(n_216),
.Y(n_324)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_285),
.Y(n_325)
);

HB1xp67_ASAP7_75t_L g326 ( 
.A(n_163),
.Y(n_326)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_285),
.Y(n_327)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_285),
.Y(n_328)
);

CKINVDCx20_ASAP7_75t_R g329 ( 
.A(n_251),
.Y(n_329)
);

CKINVDCx5p33_ASAP7_75t_R g330 ( 
.A(n_254),
.Y(n_330)
);

CKINVDCx5p33_ASAP7_75t_R g331 ( 
.A(n_260),
.Y(n_331)
);

INVxp67_ASAP7_75t_SL g332 ( 
.A(n_175),
.Y(n_332)
);

HB1xp67_ASAP7_75t_L g333 ( 
.A(n_288),
.Y(n_333)
);

CKINVDCx16_ASAP7_75t_R g334 ( 
.A(n_274),
.Y(n_334)
);

CKINVDCx5p33_ASAP7_75t_R g335 ( 
.A(n_270),
.Y(n_335)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_285),
.Y(n_336)
);

CKINVDCx20_ASAP7_75t_R g337 ( 
.A(n_305),
.Y(n_337)
);

INVx1_ASAP7_75t_L g338 ( 
.A(n_285),
.Y(n_338)
);

NOR2xp67_ASAP7_75t_L g339 ( 
.A(n_159),
.B(n_1),
.Y(n_339)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_167),
.Y(n_340)
);

CKINVDCx20_ASAP7_75t_R g341 ( 
.A(n_307),
.Y(n_341)
);

INVx1_ASAP7_75t_L g342 ( 
.A(n_167),
.Y(n_342)
);

CKINVDCx5p33_ASAP7_75t_R g343 ( 
.A(n_161),
.Y(n_343)
);

CKINVDCx20_ASAP7_75t_R g344 ( 
.A(n_162),
.Y(n_344)
);

INVx1_ASAP7_75t_L g345 ( 
.A(n_173),
.Y(n_345)
);

INVx1_ASAP7_75t_L g346 ( 
.A(n_173),
.Y(n_346)
);

NAND2xp5_ASAP7_75t_L g347 ( 
.A(n_237),
.B(n_5),
.Y(n_347)
);

INVx1_ASAP7_75t_L g348 ( 
.A(n_174),
.Y(n_348)
);

INVx1_ASAP7_75t_L g349 ( 
.A(n_174),
.Y(n_349)
);

CKINVDCx5p33_ASAP7_75t_R g350 ( 
.A(n_168),
.Y(n_350)
);

HB1xp67_ASAP7_75t_L g351 ( 
.A(n_175),
.Y(n_351)
);

INVx1_ASAP7_75t_L g352 ( 
.A(n_178),
.Y(n_352)
);

INVx1_ASAP7_75t_L g353 ( 
.A(n_178),
.Y(n_353)
);

NOR2xp33_ASAP7_75t_L g354 ( 
.A(n_185),
.B(n_6),
.Y(n_354)
);

HB1xp67_ASAP7_75t_L g355 ( 
.A(n_210),
.Y(n_355)
);

INVx1_ASAP7_75t_L g356 ( 
.A(n_185),
.Y(n_356)
);

INVx1_ASAP7_75t_L g357 ( 
.A(n_199),
.Y(n_357)
);

HB1xp67_ASAP7_75t_L g358 ( 
.A(n_187),
.Y(n_358)
);

CKINVDCx5p33_ASAP7_75t_R g359 ( 
.A(n_170),
.Y(n_359)
);

INVx2_ASAP7_75t_L g360 ( 
.A(n_283),
.Y(n_360)
);

HB1xp67_ASAP7_75t_L g361 ( 
.A(n_187),
.Y(n_361)
);

CKINVDCx5p33_ASAP7_75t_R g362 ( 
.A(n_177),
.Y(n_362)
);

INVx1_ASAP7_75t_L g363 ( 
.A(n_199),
.Y(n_363)
);

CKINVDCx20_ASAP7_75t_R g364 ( 
.A(n_171),
.Y(n_364)
);

INVxp67_ASAP7_75t_SL g365 ( 
.A(n_214),
.Y(n_365)
);

INVx1_ASAP7_75t_L g366 ( 
.A(n_209),
.Y(n_366)
);

CKINVDCx20_ASAP7_75t_R g367 ( 
.A(n_188),
.Y(n_367)
);

INVx1_ASAP7_75t_L g368 ( 
.A(n_209),
.Y(n_368)
);

CKINVDCx5p33_ASAP7_75t_R g369 ( 
.A(n_179),
.Y(n_369)
);

NOR2xp33_ASAP7_75t_L g370 ( 
.A(n_311),
.B(n_6),
.Y(n_370)
);

CKINVDCx5p33_ASAP7_75t_R g371 ( 
.A(n_180),
.Y(n_371)
);

INVx1_ASAP7_75t_L g372 ( 
.A(n_215),
.Y(n_372)
);

CKINVDCx5p33_ASAP7_75t_R g373 ( 
.A(n_181),
.Y(n_373)
);

NOR2xp67_ASAP7_75t_L g374 ( 
.A(n_200),
.B(n_7),
.Y(n_374)
);

CKINVDCx5p33_ASAP7_75t_R g375 ( 
.A(n_189),
.Y(n_375)
);

CKINVDCx20_ASAP7_75t_R g376 ( 
.A(n_191),
.Y(n_376)
);

INVx1_ASAP7_75t_L g377 ( 
.A(n_215),
.Y(n_377)
);

CKINVDCx5p33_ASAP7_75t_R g378 ( 
.A(n_190),
.Y(n_378)
);

NOR2xp67_ASAP7_75t_L g379 ( 
.A(n_200),
.B(n_8),
.Y(n_379)
);

CKINVDCx5p33_ASAP7_75t_R g380 ( 
.A(n_201),
.Y(n_380)
);

INVxp67_ASAP7_75t_SL g381 ( 
.A(n_214),
.Y(n_381)
);

INVx1_ASAP7_75t_L g382 ( 
.A(n_234),
.Y(n_382)
);

INVxp67_ASAP7_75t_SL g383 ( 
.A(n_220),
.Y(n_383)
);

CKINVDCx5p33_ASAP7_75t_R g384 ( 
.A(n_219),
.Y(n_384)
);

CKINVDCx5p33_ASAP7_75t_R g385 ( 
.A(n_222),
.Y(n_385)
);

INVx1_ASAP7_75t_L g386 ( 
.A(n_234),
.Y(n_386)
);

INVx3_ASAP7_75t_L g387 ( 
.A(n_360),
.Y(n_387)
);

NAND2xp5_ASAP7_75t_SL g388 ( 
.A(n_334),
.B(n_274),
.Y(n_388)
);

INVx2_ASAP7_75t_L g389 ( 
.A(n_319),
.Y(n_389)
);

INVx1_ASAP7_75t_L g390 ( 
.A(n_315),
.Y(n_390)
);

CKINVDCx5p33_ASAP7_75t_R g391 ( 
.A(n_324),
.Y(n_391)
);

NOR2xp67_ASAP7_75t_L g392 ( 
.A(n_340),
.B(n_164),
.Y(n_392)
);

INVx1_ASAP7_75t_L g393 ( 
.A(n_315),
.Y(n_393)
);

INVx1_ASAP7_75t_L g394 ( 
.A(n_323),
.Y(n_394)
);

BUFx6f_ASAP7_75t_L g395 ( 
.A(n_319),
.Y(n_395)
);

INVx3_ASAP7_75t_L g396 ( 
.A(n_360),
.Y(n_396)
);

INVx3_ASAP7_75t_L g397 ( 
.A(n_360),
.Y(n_397)
);

CKINVDCx5p33_ASAP7_75t_R g398 ( 
.A(n_330),
.Y(n_398)
);

AND2x4_ASAP7_75t_L g399 ( 
.A(n_340),
.B(n_192),
.Y(n_399)
);

CKINVDCx5p33_ASAP7_75t_R g400 ( 
.A(n_331),
.Y(n_400)
);

NOR2xp33_ASAP7_75t_L g401 ( 
.A(n_321),
.B(n_242),
.Y(n_401)
);

HB1xp67_ASAP7_75t_L g402 ( 
.A(n_326),
.Y(n_402)
);

CKINVDCx5p33_ASAP7_75t_R g403 ( 
.A(n_335),
.Y(n_403)
);

BUFx6f_ASAP7_75t_L g404 ( 
.A(n_319),
.Y(n_404)
);

AND2x2_ASAP7_75t_L g405 ( 
.A(n_342),
.B(n_192),
.Y(n_405)
);

INVx1_ASAP7_75t_L g406 ( 
.A(n_323),
.Y(n_406)
);

INVx1_ASAP7_75t_L g407 ( 
.A(n_325),
.Y(n_407)
);

AND2x2_ASAP7_75t_L g408 ( 
.A(n_342),
.B(n_345),
.Y(n_408)
);

INVx1_ASAP7_75t_L g409 ( 
.A(n_325),
.Y(n_409)
);

BUFx8_ASAP7_75t_L g410 ( 
.A(n_320),
.Y(n_410)
);

INVx1_ASAP7_75t_L g411 ( 
.A(n_327),
.Y(n_411)
);

CKINVDCx5p33_ASAP7_75t_R g412 ( 
.A(n_322),
.Y(n_412)
);

INVx2_ASAP7_75t_L g413 ( 
.A(n_327),
.Y(n_413)
);

INVx1_ASAP7_75t_L g414 ( 
.A(n_328),
.Y(n_414)
);

INVx2_ASAP7_75t_L g415 ( 
.A(n_328),
.Y(n_415)
);

CKINVDCx5p33_ASAP7_75t_R g416 ( 
.A(n_329),
.Y(n_416)
);

AND2x2_ASAP7_75t_L g417 ( 
.A(n_345),
.B(n_346),
.Y(n_417)
);

OAI21x1_ASAP7_75t_L g418 ( 
.A1(n_314),
.A2(n_245),
.B(n_242),
.Y(n_418)
);

CKINVDCx20_ASAP7_75t_R g419 ( 
.A(n_344),
.Y(n_419)
);

CKINVDCx20_ASAP7_75t_R g420 ( 
.A(n_364),
.Y(n_420)
);

BUFx8_ASAP7_75t_L g421 ( 
.A(n_320),
.Y(n_421)
);

OA21x2_ASAP7_75t_L g422 ( 
.A1(n_314),
.A2(n_249),
.B(n_245),
.Y(n_422)
);

INVx1_ASAP7_75t_L g423 ( 
.A(n_336),
.Y(n_423)
);

CKINVDCx5p33_ASAP7_75t_R g424 ( 
.A(n_337),
.Y(n_424)
);

CKINVDCx20_ASAP7_75t_R g425 ( 
.A(n_367),
.Y(n_425)
);

CKINVDCx5p33_ASAP7_75t_R g426 ( 
.A(n_341),
.Y(n_426)
);

INVx3_ASAP7_75t_L g427 ( 
.A(n_336),
.Y(n_427)
);

INVx1_ASAP7_75t_L g428 ( 
.A(n_338),
.Y(n_428)
);

BUFx2_ASAP7_75t_L g429 ( 
.A(n_333),
.Y(n_429)
);

HB1xp67_ASAP7_75t_L g430 ( 
.A(n_326),
.Y(n_430)
);

AND2x2_ASAP7_75t_L g431 ( 
.A(n_346),
.B(n_192),
.Y(n_431)
);

INVx1_ASAP7_75t_L g432 ( 
.A(n_338),
.Y(n_432)
);

INVx1_ASAP7_75t_L g433 ( 
.A(n_348),
.Y(n_433)
);

CKINVDCx5p33_ASAP7_75t_R g434 ( 
.A(n_343),
.Y(n_434)
);

CKINVDCx5p33_ASAP7_75t_R g435 ( 
.A(n_350),
.Y(n_435)
);

INVx1_ASAP7_75t_L g436 ( 
.A(n_348),
.Y(n_436)
);

NAND2xp5_ASAP7_75t_L g437 ( 
.A(n_349),
.B(n_249),
.Y(n_437)
);

INVx1_ASAP7_75t_L g438 ( 
.A(n_349),
.Y(n_438)
);

NAND2xp5_ASAP7_75t_L g439 ( 
.A(n_352),
.B(n_297),
.Y(n_439)
);

CKINVDCx20_ASAP7_75t_R g440 ( 
.A(n_376),
.Y(n_440)
);

NOR2xp33_ASAP7_75t_L g441 ( 
.A(n_347),
.B(n_297),
.Y(n_441)
);

CKINVDCx5p33_ASAP7_75t_R g442 ( 
.A(n_359),
.Y(n_442)
);

CKINVDCx20_ASAP7_75t_R g443 ( 
.A(n_334),
.Y(n_443)
);

HB1xp67_ASAP7_75t_L g444 ( 
.A(n_355),
.Y(n_444)
);

CKINVDCx5p33_ASAP7_75t_R g445 ( 
.A(n_362),
.Y(n_445)
);

CKINVDCx5p33_ASAP7_75t_R g446 ( 
.A(n_369),
.Y(n_446)
);

NOR2xp33_ASAP7_75t_R g447 ( 
.A(n_371),
.B(n_165),
.Y(n_447)
);

NOR2xp33_ASAP7_75t_SL g448 ( 
.A(n_316),
.B(n_228),
.Y(n_448)
);

INVx2_ASAP7_75t_L g449 ( 
.A(n_352),
.Y(n_449)
);

CKINVDCx20_ASAP7_75t_R g450 ( 
.A(n_312),
.Y(n_450)
);

INVx2_ASAP7_75t_L g451 ( 
.A(n_353),
.Y(n_451)
);

NOR2xp67_ASAP7_75t_L g452 ( 
.A(n_353),
.B(n_356),
.Y(n_452)
);

INVx1_ASAP7_75t_L g453 ( 
.A(n_356),
.Y(n_453)
);

CKINVDCx5p33_ASAP7_75t_R g454 ( 
.A(n_373),
.Y(n_454)
);

INVx1_ASAP7_75t_L g455 ( 
.A(n_357),
.Y(n_455)
);

INVx1_ASAP7_75t_L g456 ( 
.A(n_357),
.Y(n_456)
);

NAND2xp5_ASAP7_75t_L g457 ( 
.A(n_363),
.B(n_301),
.Y(n_457)
);

CKINVDCx5p33_ASAP7_75t_R g458 ( 
.A(n_375),
.Y(n_458)
);

NAND2xp5_ASAP7_75t_SL g459 ( 
.A(n_448),
.B(n_441),
.Y(n_459)
);

NAND2xp5_ASAP7_75t_SL g460 ( 
.A(n_448),
.B(n_378),
.Y(n_460)
);

OAI22xp33_ASAP7_75t_SL g461 ( 
.A1(n_441),
.A2(n_347),
.B1(n_317),
.B2(n_365),
.Y(n_461)
);

INVx1_ASAP7_75t_L g462 ( 
.A(n_433),
.Y(n_462)
);

INVx2_ASAP7_75t_L g463 ( 
.A(n_389),
.Y(n_463)
);

AND2x6_ASAP7_75t_L g464 ( 
.A(n_408),
.B(n_301),
.Y(n_464)
);

NOR2xp33_ASAP7_75t_L g465 ( 
.A(n_401),
.B(n_380),
.Y(n_465)
);

INVx4_ASAP7_75t_L g466 ( 
.A(n_427),
.Y(n_466)
);

AOI22xp5_ASAP7_75t_L g467 ( 
.A1(n_401),
.A2(n_385),
.B1(n_384),
.B2(n_370),
.Y(n_467)
);

OR2x6_ASAP7_75t_L g468 ( 
.A(n_388),
.B(n_339),
.Y(n_468)
);

INVx2_ASAP7_75t_L g469 ( 
.A(n_389),
.Y(n_469)
);

BUFx4f_ASAP7_75t_L g470 ( 
.A(n_422),
.Y(n_470)
);

NAND2xp5_ASAP7_75t_L g471 ( 
.A(n_408),
.B(n_417),
.Y(n_471)
);

BUFx3_ASAP7_75t_L g472 ( 
.A(n_390),
.Y(n_472)
);

NAND2xp5_ASAP7_75t_L g473 ( 
.A(n_408),
.B(n_417),
.Y(n_473)
);

BUFx6f_ASAP7_75t_SL g474 ( 
.A(n_399),
.Y(n_474)
);

INVx1_ASAP7_75t_L g475 ( 
.A(n_433),
.Y(n_475)
);

INVx3_ASAP7_75t_L g476 ( 
.A(n_427),
.Y(n_476)
);

INVx1_ASAP7_75t_L g477 ( 
.A(n_436),
.Y(n_477)
);

BUFx2_ASAP7_75t_L g478 ( 
.A(n_443),
.Y(n_478)
);

NAND2xp5_ASAP7_75t_L g479 ( 
.A(n_417),
.B(n_436),
.Y(n_479)
);

NOR2xp33_ASAP7_75t_L g480 ( 
.A(n_438),
.B(n_363),
.Y(n_480)
);

NOR2xp33_ASAP7_75t_L g481 ( 
.A(n_453),
.B(n_366),
.Y(n_481)
);

NOR2xp33_ASAP7_75t_L g482 ( 
.A(n_453),
.B(n_366),
.Y(n_482)
);

NOR2x1p5_ASAP7_75t_L g483 ( 
.A(n_434),
.B(n_313),
.Y(n_483)
);

AO22x2_ASAP7_75t_L g484 ( 
.A1(n_421),
.A2(n_365),
.B1(n_383),
.B2(n_332),
.Y(n_484)
);

INVx6_ASAP7_75t_L g485 ( 
.A(n_421),
.Y(n_485)
);

NAND2xp5_ASAP7_75t_L g486 ( 
.A(n_455),
.B(n_368),
.Y(n_486)
);

HB1xp67_ASAP7_75t_L g487 ( 
.A(n_429),
.Y(n_487)
);

AOI22xp5_ASAP7_75t_L g488 ( 
.A1(n_421),
.A2(n_354),
.B1(n_383),
.B2(n_381),
.Y(n_488)
);

NAND2xp5_ASAP7_75t_L g489 ( 
.A(n_455),
.B(n_368),
.Y(n_489)
);

INVx4_ASAP7_75t_L g490 ( 
.A(n_427),
.Y(n_490)
);

BUFx3_ASAP7_75t_L g491 ( 
.A(n_390),
.Y(n_491)
);

AOI22xp33_ASAP7_75t_L g492 ( 
.A1(n_422),
.A2(n_374),
.B1(n_339),
.B2(n_379),
.Y(n_492)
);

NAND2xp5_ASAP7_75t_SL g493 ( 
.A(n_427),
.B(n_311),
.Y(n_493)
);

AND2x2_ASAP7_75t_L g494 ( 
.A(n_405),
.B(n_313),
.Y(n_494)
);

NAND2xp5_ASAP7_75t_L g495 ( 
.A(n_456),
.B(n_372),
.Y(n_495)
);

NAND2xp5_ASAP7_75t_L g496 ( 
.A(n_456),
.B(n_372),
.Y(n_496)
);

INVx4_ASAP7_75t_SL g497 ( 
.A(n_395),
.Y(n_497)
);

NAND2xp5_ASAP7_75t_SL g498 ( 
.A(n_447),
.B(n_377),
.Y(n_498)
);

INVx2_ASAP7_75t_L g499 ( 
.A(n_389),
.Y(n_499)
);

INVx3_ASAP7_75t_L g500 ( 
.A(n_413),
.Y(n_500)
);

INVxp67_ASAP7_75t_SL g501 ( 
.A(n_452),
.Y(n_501)
);

INVx1_ASAP7_75t_L g502 ( 
.A(n_449),
.Y(n_502)
);

OAI21xp33_ASAP7_75t_SL g503 ( 
.A1(n_418),
.A2(n_382),
.B(n_377),
.Y(n_503)
);

INVx1_ASAP7_75t_L g504 ( 
.A(n_449),
.Y(n_504)
);

AOI22xp33_ASAP7_75t_L g505 ( 
.A1(n_422),
.A2(n_379),
.B1(n_374),
.B2(n_386),
.Y(n_505)
);

INVx1_ASAP7_75t_L g506 ( 
.A(n_449),
.Y(n_506)
);

AOI22xp33_ASAP7_75t_L g507 ( 
.A1(n_422),
.A2(n_386),
.B1(n_382),
.B2(n_381),
.Y(n_507)
);

NAND2xp5_ASAP7_75t_SL g508 ( 
.A(n_447),
.B(n_166),
.Y(n_508)
);

INVx2_ASAP7_75t_L g509 ( 
.A(n_413),
.Y(n_509)
);

INVx1_ASAP7_75t_L g510 ( 
.A(n_451),
.Y(n_510)
);

INVx3_ASAP7_75t_L g511 ( 
.A(n_413),
.Y(n_511)
);

INVx5_ASAP7_75t_L g512 ( 
.A(n_395),
.Y(n_512)
);

INVx2_ASAP7_75t_SL g513 ( 
.A(n_444),
.Y(n_513)
);

INVx1_ASAP7_75t_L g514 ( 
.A(n_451),
.Y(n_514)
);

NAND2xp5_ASAP7_75t_L g515 ( 
.A(n_392),
.B(n_332),
.Y(n_515)
);

NAND2xp5_ASAP7_75t_L g516 ( 
.A(n_392),
.B(n_318),
.Y(n_516)
);

INVx1_ASAP7_75t_L g517 ( 
.A(n_451),
.Y(n_517)
);

HB1xp67_ASAP7_75t_L g518 ( 
.A(n_429),
.Y(n_518)
);

INVx1_ASAP7_75t_L g519 ( 
.A(n_452),
.Y(n_519)
);

INVx2_ASAP7_75t_L g520 ( 
.A(n_415),
.Y(n_520)
);

NOR2xp33_ASAP7_75t_L g521 ( 
.A(n_435),
.B(n_361),
.Y(n_521)
);

NAND2xp5_ASAP7_75t_L g522 ( 
.A(n_393),
.B(n_318),
.Y(n_522)
);

INVx2_ASAP7_75t_SL g523 ( 
.A(n_444),
.Y(n_523)
);

AND2x4_ASAP7_75t_L g524 ( 
.A(n_399),
.B(n_351),
.Y(n_524)
);

INVx3_ASAP7_75t_L g525 ( 
.A(n_415),
.Y(n_525)
);

INVx6_ASAP7_75t_L g526 ( 
.A(n_421),
.Y(n_526)
);

BUFx2_ASAP7_75t_L g527 ( 
.A(n_442),
.Y(n_527)
);

INVx1_ASAP7_75t_L g528 ( 
.A(n_415),
.Y(n_528)
);

INVx1_ASAP7_75t_L g529 ( 
.A(n_405),
.Y(n_529)
);

BUFx6f_ASAP7_75t_L g530 ( 
.A(n_395),
.Y(n_530)
);

BUFx4_ASAP7_75t_L g531 ( 
.A(n_419),
.Y(n_531)
);

INVx2_ASAP7_75t_L g532 ( 
.A(n_395),
.Y(n_532)
);

INVx2_ASAP7_75t_L g533 ( 
.A(n_395),
.Y(n_533)
);

NAND2xp33_ASAP7_75t_L g534 ( 
.A(n_393),
.B(n_283),
.Y(n_534)
);

NAND2xp5_ASAP7_75t_SL g535 ( 
.A(n_394),
.B(n_169),
.Y(n_535)
);

CKINVDCx5p33_ASAP7_75t_R g536 ( 
.A(n_391),
.Y(n_536)
);

AOI22xp5_ASAP7_75t_L g537 ( 
.A1(n_421),
.A2(n_208),
.B1(n_277),
.B2(n_303),
.Y(n_537)
);

NOR2x1p5_ASAP7_75t_L g538 ( 
.A(n_445),
.B(n_210),
.Y(n_538)
);

AND2x2_ASAP7_75t_L g539 ( 
.A(n_431),
.B(n_351),
.Y(n_539)
);

INVx1_ASAP7_75t_L g540 ( 
.A(n_431),
.Y(n_540)
);

BUFx8_ASAP7_75t_SL g541 ( 
.A(n_450),
.Y(n_541)
);

AND2x2_ASAP7_75t_L g542 ( 
.A(n_399),
.B(n_358),
.Y(n_542)
);

NAND2xp5_ASAP7_75t_SL g543 ( 
.A(n_394),
.B(n_176),
.Y(n_543)
);

AND2x2_ASAP7_75t_L g544 ( 
.A(n_399),
.B(n_358),
.Y(n_544)
);

BUFx8_ASAP7_75t_SL g545 ( 
.A(n_420),
.Y(n_545)
);

NOR2x1p5_ASAP7_75t_L g546 ( 
.A(n_446),
.B(n_310),
.Y(n_546)
);

CKINVDCx16_ASAP7_75t_R g547 ( 
.A(n_425),
.Y(n_547)
);

BUFx3_ASAP7_75t_L g548 ( 
.A(n_406),
.Y(n_548)
);

INVx5_ASAP7_75t_L g549 ( 
.A(n_395),
.Y(n_549)
);

NAND2xp5_ASAP7_75t_L g550 ( 
.A(n_406),
.B(n_217),
.Y(n_550)
);

AND2x2_ASAP7_75t_L g551 ( 
.A(n_399),
.B(n_361),
.Y(n_551)
);

INVx2_ASAP7_75t_L g552 ( 
.A(n_395),
.Y(n_552)
);

INVx2_ASAP7_75t_L g553 ( 
.A(n_404),
.Y(n_553)
);

BUFx3_ASAP7_75t_L g554 ( 
.A(n_407),
.Y(n_554)
);

INVx2_ASAP7_75t_L g555 ( 
.A(n_404),
.Y(n_555)
);

INVxp33_ASAP7_75t_L g556 ( 
.A(n_402),
.Y(n_556)
);

INVx1_ASAP7_75t_L g557 ( 
.A(n_407),
.Y(n_557)
);

BUFx4f_ASAP7_75t_L g558 ( 
.A(n_422),
.Y(n_558)
);

NAND2xp5_ASAP7_75t_L g559 ( 
.A(n_409),
.B(n_279),
.Y(n_559)
);

NAND2xp5_ASAP7_75t_L g560 ( 
.A(n_409),
.B(n_182),
.Y(n_560)
);

OR2x2_ASAP7_75t_L g561 ( 
.A(n_402),
.B(n_430),
.Y(n_561)
);

BUFx2_ASAP7_75t_L g562 ( 
.A(n_454),
.Y(n_562)
);

INVx2_ASAP7_75t_SL g563 ( 
.A(n_410),
.Y(n_563)
);

NOR2xp33_ASAP7_75t_L g564 ( 
.A(n_458),
.B(n_310),
.Y(n_564)
);

INVx3_ASAP7_75t_L g565 ( 
.A(n_404),
.Y(n_565)
);

NAND2xp5_ASAP7_75t_L g566 ( 
.A(n_411),
.B(n_414),
.Y(n_566)
);

NOR2xp33_ASAP7_75t_L g567 ( 
.A(n_430),
.B(n_223),
.Y(n_567)
);

INVx5_ASAP7_75t_L g568 ( 
.A(n_404),
.Y(n_568)
);

BUFx3_ASAP7_75t_L g569 ( 
.A(n_411),
.Y(n_569)
);

INVx1_ASAP7_75t_L g570 ( 
.A(n_414),
.Y(n_570)
);

INVxp67_ASAP7_75t_SL g571 ( 
.A(n_404),
.Y(n_571)
);

NAND2xp5_ASAP7_75t_L g572 ( 
.A(n_423),
.B(n_183),
.Y(n_572)
);

NAND2xp5_ASAP7_75t_SL g573 ( 
.A(n_423),
.B(n_184),
.Y(n_573)
);

NAND2xp5_ASAP7_75t_L g574 ( 
.A(n_428),
.B(n_186),
.Y(n_574)
);

NAND2xp5_ASAP7_75t_SL g575 ( 
.A(n_428),
.B(n_193),
.Y(n_575)
);

INVx1_ASAP7_75t_SL g576 ( 
.A(n_440),
.Y(n_576)
);

INVx2_ASAP7_75t_L g577 ( 
.A(n_404),
.Y(n_577)
);

NAND2xp33_ASAP7_75t_L g578 ( 
.A(n_432),
.B(n_283),
.Y(n_578)
);

INVx2_ASAP7_75t_L g579 ( 
.A(n_404),
.Y(n_579)
);

NOR2xp33_ASAP7_75t_L g580 ( 
.A(n_432),
.B(n_225),
.Y(n_580)
);

INVx3_ASAP7_75t_L g581 ( 
.A(n_387),
.Y(n_581)
);

INVx2_ASAP7_75t_SL g582 ( 
.A(n_410),
.Y(n_582)
);

INVx1_ASAP7_75t_L g583 ( 
.A(n_437),
.Y(n_583)
);

NOR2xp33_ASAP7_75t_L g584 ( 
.A(n_437),
.B(n_226),
.Y(n_584)
);

INVx1_ASAP7_75t_L g585 ( 
.A(n_439),
.Y(n_585)
);

AOI22xp5_ASAP7_75t_L g586 ( 
.A1(n_410),
.A2(n_229),
.B1(n_308),
.B2(n_227),
.Y(n_586)
);

OR2x2_ASAP7_75t_L g587 ( 
.A(n_398),
.B(n_220),
.Y(n_587)
);

INVx1_ASAP7_75t_L g588 ( 
.A(n_439),
.Y(n_588)
);

NOR2xp33_ASAP7_75t_L g589 ( 
.A(n_457),
.B(n_235),
.Y(n_589)
);

INVx1_ASAP7_75t_L g590 ( 
.A(n_457),
.Y(n_590)
);

AND2x4_ASAP7_75t_L g591 ( 
.A(n_418),
.B(n_224),
.Y(n_591)
);

OR2x6_ASAP7_75t_L g592 ( 
.A(n_410),
.B(n_236),
.Y(n_592)
);

INVx1_ASAP7_75t_L g593 ( 
.A(n_387),
.Y(n_593)
);

BUFx4f_ASAP7_75t_L g594 ( 
.A(n_387),
.Y(n_594)
);

NAND2xp5_ASAP7_75t_L g595 ( 
.A(n_387),
.B(n_194),
.Y(n_595)
);

OR2x2_ASAP7_75t_L g596 ( 
.A(n_400),
.B(n_224),
.Y(n_596)
);

INVx2_ASAP7_75t_L g597 ( 
.A(n_396),
.Y(n_597)
);

INVxp67_ASAP7_75t_SL g598 ( 
.A(n_418),
.Y(n_598)
);

BUFx3_ASAP7_75t_L g599 ( 
.A(n_403),
.Y(n_599)
);

NOR2xp33_ASAP7_75t_L g600 ( 
.A(n_396),
.B(n_241),
.Y(n_600)
);

INVx2_ASAP7_75t_L g601 ( 
.A(n_396),
.Y(n_601)
);

NAND2xp5_ASAP7_75t_L g602 ( 
.A(n_396),
.B(n_195),
.Y(n_602)
);

INVx1_ASAP7_75t_SL g603 ( 
.A(n_412),
.Y(n_603)
);

OAI22xp5_ASAP7_75t_L g604 ( 
.A1(n_416),
.A2(n_261),
.B1(n_280),
.B2(n_263),
.Y(n_604)
);

INVx2_ASAP7_75t_L g605 ( 
.A(n_397),
.Y(n_605)
);

NAND3xp33_ASAP7_75t_L g606 ( 
.A(n_397),
.B(n_289),
.C(n_243),
.Y(n_606)
);

NAND2xp5_ASAP7_75t_SL g607 ( 
.A(n_459),
.B(n_290),
.Y(n_607)
);

A2O1A1Ixp33_ASAP7_75t_L g608 ( 
.A1(n_459),
.A2(n_265),
.B(n_240),
.C(n_250),
.Y(n_608)
);

INVx1_ASAP7_75t_L g609 ( 
.A(n_472),
.Y(n_609)
);

NAND2xp5_ASAP7_75t_L g610 ( 
.A(n_583),
.B(n_397),
.Y(n_610)
);

NAND2xp5_ASAP7_75t_L g611 ( 
.A(n_585),
.B(n_397),
.Y(n_611)
);

CKINVDCx11_ASAP7_75t_R g612 ( 
.A(n_547),
.Y(n_612)
);

CKINVDCx20_ASAP7_75t_R g613 ( 
.A(n_545),
.Y(n_613)
);

NAND2xp5_ASAP7_75t_L g614 ( 
.A(n_588),
.B(n_236),
.Y(n_614)
);

NOR2xp33_ASAP7_75t_L g615 ( 
.A(n_465),
.B(n_248),
.Y(n_615)
);

CKINVDCx5p33_ASAP7_75t_R g616 ( 
.A(n_536),
.Y(n_616)
);

NAND2xp5_ASAP7_75t_L g617 ( 
.A(n_590),
.B(n_258),
.Y(n_617)
);

NOR2xp33_ASAP7_75t_L g618 ( 
.A(n_460),
.B(n_252),
.Y(n_618)
);

NAND2xp5_ASAP7_75t_L g619 ( 
.A(n_584),
.B(n_258),
.Y(n_619)
);

INVxp67_ASAP7_75t_L g620 ( 
.A(n_521),
.Y(n_620)
);

NOR2xp33_ASAP7_75t_L g621 ( 
.A(n_460),
.B(n_253),
.Y(n_621)
);

AOI22xp5_ASAP7_75t_L g622 ( 
.A1(n_464),
.A2(n_211),
.B1(n_309),
.B2(n_306),
.Y(n_622)
);

NAND2xp5_ASAP7_75t_SL g623 ( 
.A(n_470),
.B(n_290),
.Y(n_623)
);

NAND2xp5_ASAP7_75t_L g624 ( 
.A(n_589),
.B(n_268),
.Y(n_624)
);

INVx2_ASAP7_75t_L g625 ( 
.A(n_500),
.Y(n_625)
);

NAND2xp5_ASAP7_75t_SL g626 ( 
.A(n_470),
.B(n_290),
.Y(n_626)
);

INVx2_ASAP7_75t_L g627 ( 
.A(n_500),
.Y(n_627)
);

NAND2xp33_ASAP7_75t_L g628 ( 
.A(n_464),
.B(n_476),
.Y(n_628)
);

INVx1_ASAP7_75t_L g629 ( 
.A(n_472),
.Y(n_629)
);

NOR3xp33_ASAP7_75t_L g630 ( 
.A(n_527),
.B(n_426),
.C(n_424),
.Y(n_630)
);

AND2x2_ASAP7_75t_L g631 ( 
.A(n_513),
.B(n_228),
.Y(n_631)
);

NAND2xp5_ASAP7_75t_SL g632 ( 
.A(n_470),
.B(n_290),
.Y(n_632)
);

AOI22xp33_ASAP7_75t_L g633 ( 
.A1(n_464),
.A2(n_268),
.B1(n_302),
.B2(n_275),
.Y(n_633)
);

INVx8_ASAP7_75t_L g634 ( 
.A(n_592),
.Y(n_634)
);

INVx2_ASAP7_75t_L g635 ( 
.A(n_500),
.Y(n_635)
);

OR2x6_ASAP7_75t_L g636 ( 
.A(n_592),
.B(n_302),
.Y(n_636)
);

NAND2xp5_ASAP7_75t_SL g637 ( 
.A(n_558),
.B(n_290),
.Y(n_637)
);

NAND2xp5_ASAP7_75t_L g638 ( 
.A(n_515),
.B(n_231),
.Y(n_638)
);

NOR3xp33_ASAP7_75t_L g639 ( 
.A(n_562),
.B(n_304),
.C(n_239),
.Y(n_639)
);

INVx1_ASAP7_75t_L g640 ( 
.A(n_491),
.Y(n_640)
);

NAND2xp5_ASAP7_75t_L g641 ( 
.A(n_494),
.B(n_231),
.Y(n_641)
);

INVx3_ASAP7_75t_L g642 ( 
.A(n_491),
.Y(n_642)
);

NAND2xp5_ASAP7_75t_L g643 ( 
.A(n_494),
.B(n_239),
.Y(n_643)
);

AND2x2_ASAP7_75t_L g644 ( 
.A(n_513),
.B(n_228),
.Y(n_644)
);

NAND2xp5_ASAP7_75t_L g645 ( 
.A(n_580),
.B(n_240),
.Y(n_645)
);

AOI22xp5_ASAP7_75t_L g646 ( 
.A1(n_464),
.A2(n_203),
.B1(n_196),
.B2(n_197),
.Y(n_646)
);

NAND2xp5_ASAP7_75t_SL g647 ( 
.A(n_558),
.B(n_298),
.Y(n_647)
);

NAND2xp5_ASAP7_75t_L g648 ( 
.A(n_480),
.B(n_246),
.Y(n_648)
);

AOI221xp5_ASAP7_75t_L g649 ( 
.A1(n_461),
.A2(n_304),
.B1(n_250),
.B2(n_265),
.C(n_296),
.Y(n_649)
);

NAND2xp5_ASAP7_75t_SL g650 ( 
.A(n_558),
.B(n_466),
.Y(n_650)
);

INVx2_ASAP7_75t_L g651 ( 
.A(n_511),
.Y(n_651)
);

AOI22xp33_ASAP7_75t_L g652 ( 
.A1(n_464),
.A2(n_276),
.B1(n_246),
.B2(n_296),
.Y(n_652)
);

AOI22xp5_ASAP7_75t_L g653 ( 
.A1(n_464),
.A2(n_198),
.B1(n_202),
.B2(n_204),
.Y(n_653)
);

INVx2_ASAP7_75t_L g654 ( 
.A(n_511),
.Y(n_654)
);

AND2x2_ASAP7_75t_L g655 ( 
.A(n_523),
.B(n_228),
.Y(n_655)
);

AOI22xp5_ASAP7_75t_L g656 ( 
.A1(n_498),
.A2(n_266),
.B1(n_238),
.B2(n_205),
.Y(n_656)
);

NAND2xp5_ASAP7_75t_L g657 ( 
.A(n_481),
.B(n_247),
.Y(n_657)
);

INVx2_ASAP7_75t_L g658 ( 
.A(n_511),
.Y(n_658)
);

NAND2xp5_ASAP7_75t_L g659 ( 
.A(n_482),
.B(n_247),
.Y(n_659)
);

INVx1_ASAP7_75t_L g660 ( 
.A(n_548),
.Y(n_660)
);

HB1xp67_ASAP7_75t_L g661 ( 
.A(n_487),
.Y(n_661)
);

INVx2_ASAP7_75t_L g662 ( 
.A(n_525),
.Y(n_662)
);

NAND2xp5_ASAP7_75t_SL g663 ( 
.A(n_466),
.B(n_298),
.Y(n_663)
);

AOI22xp5_ASAP7_75t_L g664 ( 
.A1(n_498),
.A2(n_230),
.B1(n_244),
.B2(n_206),
.Y(n_664)
);

AND2x2_ASAP7_75t_L g665 ( 
.A(n_523),
.B(n_276),
.Y(n_665)
);

AND2x2_ASAP7_75t_L g666 ( 
.A(n_556),
.B(n_294),
.Y(n_666)
);

BUFx6f_ASAP7_75t_SL g667 ( 
.A(n_599),
.Y(n_667)
);

INVx2_ASAP7_75t_SL g668 ( 
.A(n_518),
.Y(n_668)
);

NOR2xp33_ASAP7_75t_L g669 ( 
.A(n_467),
.B(n_471),
.Y(n_669)
);

INVx2_ASAP7_75t_L g670 ( 
.A(n_525),
.Y(n_670)
);

NOR2xp33_ASAP7_75t_L g671 ( 
.A(n_473),
.B(n_269),
.Y(n_671)
);

NOR2xp33_ASAP7_75t_L g672 ( 
.A(n_535),
.B(n_543),
.Y(n_672)
);

NAND2xp5_ASAP7_75t_SL g673 ( 
.A(n_466),
.B(n_298),
.Y(n_673)
);

NOR2xp33_ASAP7_75t_L g674 ( 
.A(n_535),
.B(n_273),
.Y(n_674)
);

AOI22xp33_ASAP7_75t_L g675 ( 
.A1(n_484),
.A2(n_294),
.B1(n_160),
.B2(n_264),
.Y(n_675)
);

NAND2xp5_ASAP7_75t_SL g676 ( 
.A(n_490),
.B(n_298),
.Y(n_676)
);

BUFx8_ASAP7_75t_L g677 ( 
.A(n_478),
.Y(n_677)
);

NAND2xp5_ASAP7_75t_SL g678 ( 
.A(n_490),
.B(n_298),
.Y(n_678)
);

OR2x6_ASAP7_75t_L g679 ( 
.A(n_592),
.B(n_221),
.Y(n_679)
);

NOR2xp33_ASAP7_75t_L g680 ( 
.A(n_543),
.B(n_286),
.Y(n_680)
);

INVx1_ASAP7_75t_L g681 ( 
.A(n_548),
.Y(n_681)
);

INVx1_ASAP7_75t_L g682 ( 
.A(n_554),
.Y(n_682)
);

AOI22xp33_ASAP7_75t_L g683 ( 
.A1(n_484),
.A2(n_505),
.B1(n_591),
.B2(n_507),
.Y(n_683)
);

NAND2xp5_ASAP7_75t_L g684 ( 
.A(n_501),
.B(n_291),
.Y(n_684)
);

NOR2xp33_ASAP7_75t_L g685 ( 
.A(n_573),
.B(n_295),
.Y(n_685)
);

O2A1O1Ixp33_ASAP7_75t_L g686 ( 
.A1(n_479),
.A2(n_160),
.B(n_264),
.C(n_221),
.Y(n_686)
);

NAND2xp5_ASAP7_75t_L g687 ( 
.A(n_550),
.B(n_299),
.Y(n_687)
);

NAND2xp5_ASAP7_75t_SL g688 ( 
.A(n_490),
.B(n_283),
.Y(n_688)
);

AND2x2_ASAP7_75t_L g689 ( 
.A(n_556),
.B(n_300),
.Y(n_689)
);

NOR2xp33_ASAP7_75t_L g690 ( 
.A(n_573),
.B(n_11),
.Y(n_690)
);

NOR2xp33_ASAP7_75t_L g691 ( 
.A(n_575),
.B(n_12),
.Y(n_691)
);

NAND2xp5_ASAP7_75t_L g692 ( 
.A(n_559),
.B(n_207),
.Y(n_692)
);

INVx2_ASAP7_75t_SL g693 ( 
.A(n_483),
.Y(n_693)
);

INVx1_ASAP7_75t_L g694 ( 
.A(n_554),
.Y(n_694)
);

NOR2xp33_ASAP7_75t_L g695 ( 
.A(n_575),
.B(n_12),
.Y(n_695)
);

AO221x1_ASAP7_75t_L g696 ( 
.A1(n_484),
.A2(n_284),
.B1(n_15),
.B2(n_16),
.C(n_19),
.Y(n_696)
);

INVx1_ASAP7_75t_L g697 ( 
.A(n_569),
.Y(n_697)
);

INVx2_ASAP7_75t_L g698 ( 
.A(n_525),
.Y(n_698)
);

NOR2xp33_ASAP7_75t_L g699 ( 
.A(n_529),
.B(n_14),
.Y(n_699)
);

AOI221xp5_ASAP7_75t_L g700 ( 
.A1(n_567),
.A2(n_293),
.B1(n_292),
.B2(n_287),
.C(n_282),
.Y(n_700)
);

NOR2xp33_ASAP7_75t_SL g701 ( 
.A(n_536),
.B(n_160),
.Y(n_701)
);

AOI22xp5_ASAP7_75t_L g702 ( 
.A1(n_474),
.A2(n_257),
.B1(n_281),
.B2(n_272),
.Y(n_702)
);

OAI21xp5_ASAP7_75t_L g703 ( 
.A1(n_503),
.A2(n_256),
.B(n_271),
.Y(n_703)
);

INVx1_ASAP7_75t_L g704 ( 
.A(n_569),
.Y(n_704)
);

OR2x6_ASAP7_75t_L g705 ( 
.A(n_592),
.B(n_284),
.Y(n_705)
);

INVx1_ASAP7_75t_L g706 ( 
.A(n_557),
.Y(n_706)
);

INVx1_ASAP7_75t_L g707 ( 
.A(n_570),
.Y(n_707)
);

INVx2_ASAP7_75t_L g708 ( 
.A(n_463),
.Y(n_708)
);

OAI21xp5_ASAP7_75t_L g709 ( 
.A1(n_598),
.A2(n_255),
.B(n_267),
.Y(n_709)
);

AND2x2_ASAP7_75t_L g710 ( 
.A(n_539),
.B(n_14),
.Y(n_710)
);

INVx1_ASAP7_75t_L g711 ( 
.A(n_462),
.Y(n_711)
);

NOR2xp33_ASAP7_75t_L g712 ( 
.A(n_540),
.B(n_15),
.Y(n_712)
);

INVx1_ASAP7_75t_L g713 ( 
.A(n_475),
.Y(n_713)
);

AND2x6_ASAP7_75t_L g714 ( 
.A(n_485),
.B(n_86),
.Y(n_714)
);

INVx2_ASAP7_75t_SL g715 ( 
.A(n_561),
.Y(n_715)
);

INVx1_ASAP7_75t_L g716 ( 
.A(n_477),
.Y(n_716)
);

INVxp67_ASAP7_75t_L g717 ( 
.A(n_545),
.Y(n_717)
);

INVx2_ASAP7_75t_SL g718 ( 
.A(n_561),
.Y(n_718)
);

NAND2xp5_ASAP7_75t_L g719 ( 
.A(n_519),
.B(n_262),
.Y(n_719)
);

AND2x2_ASAP7_75t_L g720 ( 
.A(n_539),
.B(n_16),
.Y(n_720)
);

NOR2xp33_ASAP7_75t_L g721 ( 
.A(n_468),
.B(n_20),
.Y(n_721)
);

INVx1_ASAP7_75t_L g722 ( 
.A(n_476),
.Y(n_722)
);

NAND2xp5_ASAP7_75t_L g723 ( 
.A(n_522),
.B(n_259),
.Y(n_723)
);

INVx2_ASAP7_75t_SL g724 ( 
.A(n_587),
.Y(n_724)
);

BUFx6f_ASAP7_75t_SL g725 ( 
.A(n_599),
.Y(n_725)
);

AND2x2_ASAP7_75t_L g726 ( 
.A(n_524),
.B(n_20),
.Y(n_726)
);

NAND2xp33_ASAP7_75t_L g727 ( 
.A(n_566),
.B(n_233),
.Y(n_727)
);

OR2x6_ASAP7_75t_L g728 ( 
.A(n_563),
.B(n_23),
.Y(n_728)
);

NOR2xp33_ASAP7_75t_L g729 ( 
.A(n_468),
.B(n_26),
.Y(n_729)
);

INVx1_ASAP7_75t_L g730 ( 
.A(n_502),
.Y(n_730)
);

NAND2xp5_ASAP7_75t_L g731 ( 
.A(n_564),
.B(n_232),
.Y(n_731)
);

NAND2xp5_ASAP7_75t_L g732 ( 
.A(n_524),
.B(n_218),
.Y(n_732)
);

NAND2xp33_ASAP7_75t_L g733 ( 
.A(n_530),
.B(n_28),
.Y(n_733)
);

NAND2xp5_ASAP7_75t_L g734 ( 
.A(n_524),
.B(n_33),
.Y(n_734)
);

NAND2xp33_ASAP7_75t_L g735 ( 
.A(n_530),
.B(n_38),
.Y(n_735)
);

INVx2_ASAP7_75t_L g736 ( 
.A(n_463),
.Y(n_736)
);

NAND2xp5_ASAP7_75t_L g737 ( 
.A(n_516),
.B(n_40),
.Y(n_737)
);

NAND2xp5_ASAP7_75t_L g738 ( 
.A(n_542),
.B(n_42),
.Y(n_738)
);

INVx2_ASAP7_75t_L g739 ( 
.A(n_469),
.Y(n_739)
);

NAND2xp5_ASAP7_75t_L g740 ( 
.A(n_542),
.B(n_44),
.Y(n_740)
);

HB1xp67_ASAP7_75t_L g741 ( 
.A(n_576),
.Y(n_741)
);

BUFx12f_ASAP7_75t_L g742 ( 
.A(n_538),
.Y(n_742)
);

NAND2xp33_ASAP7_75t_L g743 ( 
.A(n_530),
.B(n_47),
.Y(n_743)
);

NOR2xp33_ASAP7_75t_L g744 ( 
.A(n_468),
.B(n_47),
.Y(n_744)
);

BUFx6f_ASAP7_75t_L g745 ( 
.A(n_485),
.Y(n_745)
);

INVx2_ASAP7_75t_L g746 ( 
.A(n_469),
.Y(n_746)
);

NAND2xp5_ASAP7_75t_SL g747 ( 
.A(n_591),
.B(n_49),
.Y(n_747)
);

INVx2_ASAP7_75t_L g748 ( 
.A(n_499),
.Y(n_748)
);

NAND2xp5_ASAP7_75t_SL g749 ( 
.A(n_591),
.B(n_51),
.Y(n_749)
);

A2O1A1Ixp33_ASAP7_75t_L g750 ( 
.A1(n_544),
.A2(n_55),
.B(n_57),
.C(n_58),
.Y(n_750)
);

NAND2xp5_ASAP7_75t_L g751 ( 
.A(n_544),
.B(n_148),
.Y(n_751)
);

NOR2xp33_ASAP7_75t_L g752 ( 
.A(n_468),
.B(n_488),
.Y(n_752)
);

NAND2xp5_ASAP7_75t_L g753 ( 
.A(n_551),
.B(n_68),
.Y(n_753)
);

INVx1_ASAP7_75t_L g754 ( 
.A(n_504),
.Y(n_754)
);

INVx2_ASAP7_75t_L g755 ( 
.A(n_499),
.Y(n_755)
);

AOI21xp5_ASAP7_75t_L g756 ( 
.A1(n_571),
.A2(n_69),
.B(n_71),
.Y(n_756)
);

NAND2xp5_ASAP7_75t_SL g757 ( 
.A(n_530),
.B(n_73),
.Y(n_757)
);

INVx1_ASAP7_75t_L g758 ( 
.A(n_506),
.Y(n_758)
);

INVx2_ASAP7_75t_L g759 ( 
.A(n_509),
.Y(n_759)
);

OR2x6_ASAP7_75t_L g760 ( 
.A(n_563),
.B(n_74),
.Y(n_760)
);

INVx1_ASAP7_75t_L g761 ( 
.A(n_510),
.Y(n_761)
);

AND2x2_ASAP7_75t_L g762 ( 
.A(n_551),
.B(n_84),
.Y(n_762)
);

AND2x2_ASAP7_75t_L g763 ( 
.A(n_587),
.B(n_91),
.Y(n_763)
);

INVx2_ASAP7_75t_L g764 ( 
.A(n_509),
.Y(n_764)
);

AOI22xp33_ASAP7_75t_L g765 ( 
.A1(n_492),
.A2(n_92),
.B1(n_96),
.B2(n_102),
.Y(n_765)
);

NAND2xp5_ASAP7_75t_L g766 ( 
.A(n_486),
.B(n_103),
.Y(n_766)
);

OAI22xp5_ASAP7_75t_L g767 ( 
.A1(n_560),
.A2(n_106),
.B1(n_107),
.B2(n_112),
.Y(n_767)
);

NAND2xp5_ASAP7_75t_SL g768 ( 
.A(n_594),
.B(n_113),
.Y(n_768)
);

INVx1_ASAP7_75t_L g769 ( 
.A(n_514),
.Y(n_769)
);

INVx2_ASAP7_75t_L g770 ( 
.A(n_520),
.Y(n_770)
);

BUFx4_ASAP7_75t_L g771 ( 
.A(n_531),
.Y(n_771)
);

O2A1O1Ixp5_ASAP7_75t_L g772 ( 
.A1(n_493),
.A2(n_115),
.B(n_124),
.C(n_125),
.Y(n_772)
);

NAND2xp5_ASAP7_75t_L g773 ( 
.A(n_489),
.B(n_139),
.Y(n_773)
);

NAND2xp5_ASAP7_75t_SL g774 ( 
.A(n_594),
.B(n_140),
.Y(n_774)
);

INVx1_ASAP7_75t_L g775 ( 
.A(n_517),
.Y(n_775)
);

INVx2_ASAP7_75t_L g776 ( 
.A(n_748),
.Y(n_776)
);

NAND3xp33_ASAP7_75t_L g777 ( 
.A(n_615),
.B(n_604),
.C(n_596),
.Y(n_777)
);

AOI22xp33_ASAP7_75t_L g778 ( 
.A1(n_752),
.A2(n_675),
.B1(n_683),
.B2(n_669),
.Y(n_778)
);

OAI21xp33_ASAP7_75t_L g779 ( 
.A1(n_615),
.A2(n_596),
.B(n_574),
.Y(n_779)
);

BUFx2_ASAP7_75t_L g780 ( 
.A(n_741),
.Y(n_780)
);

INVx1_ASAP7_75t_L g781 ( 
.A(n_706),
.Y(n_781)
);

AOI22xp5_ASAP7_75t_L g782 ( 
.A1(n_669),
.A2(n_474),
.B1(n_537),
.B2(n_508),
.Y(n_782)
);

INVx2_ASAP7_75t_L g783 ( 
.A(n_748),
.Y(n_783)
);

INVx2_ASAP7_75t_L g784 ( 
.A(n_755),
.Y(n_784)
);

NOR2x1_ASAP7_75t_L g785 ( 
.A(n_642),
.B(n_546),
.Y(n_785)
);

AOI22xp5_ASAP7_75t_L g786 ( 
.A1(n_752),
.A2(n_474),
.B1(n_508),
.B2(n_603),
.Y(n_786)
);

AOI22xp5_ASAP7_75t_L g787 ( 
.A1(n_620),
.A2(n_582),
.B1(n_586),
.B2(n_600),
.Y(n_787)
);

NAND2xp5_ASAP7_75t_L g788 ( 
.A(n_707),
.B(n_520),
.Y(n_788)
);

NAND2xp5_ASAP7_75t_L g789 ( 
.A(n_711),
.B(n_528),
.Y(n_789)
);

AOI21xp5_ASAP7_75t_L g790 ( 
.A1(n_650),
.A2(n_565),
.B(n_553),
.Y(n_790)
);

CKINVDCx20_ASAP7_75t_R g791 ( 
.A(n_613),
.Y(n_791)
);

AOI21xp5_ASAP7_75t_L g792 ( 
.A1(n_650),
.A2(n_565),
.B(n_553),
.Y(n_792)
);

NOR2xp33_ASAP7_75t_SL g793 ( 
.A(n_616),
.B(n_541),
.Y(n_793)
);

BUFx3_ASAP7_75t_L g794 ( 
.A(n_677),
.Y(n_794)
);

AOI21xp5_ASAP7_75t_L g795 ( 
.A1(n_628),
.A2(n_565),
.B(n_552),
.Y(n_795)
);

AO32x2_ASAP7_75t_L g796 ( 
.A1(n_767),
.A2(n_582),
.A3(n_493),
.B1(n_496),
.B2(n_495),
.Y(n_796)
);

INVx1_ASAP7_75t_L g797 ( 
.A(n_713),
.Y(n_797)
);

NAND2xp5_ASAP7_75t_L g798 ( 
.A(n_716),
.B(n_581),
.Y(n_798)
);

NAND2xp5_ASAP7_75t_L g799 ( 
.A(n_672),
.B(n_581),
.Y(n_799)
);

AOI21xp5_ASAP7_75t_L g800 ( 
.A1(n_610),
.A2(n_577),
.B(n_579),
.Y(n_800)
);

O2A1O1Ixp33_ASAP7_75t_SL g801 ( 
.A1(n_768),
.A2(n_572),
.B(n_593),
.C(n_602),
.Y(n_801)
);

AOI21xp5_ASAP7_75t_L g802 ( 
.A1(n_611),
.A2(n_579),
.B(n_552),
.Y(n_802)
);

AND2x4_ASAP7_75t_L g803 ( 
.A(n_636),
.B(n_581),
.Y(n_803)
);

INVx1_ASAP7_75t_L g804 ( 
.A(n_730),
.Y(n_804)
);

O2A1O1Ixp33_ASAP7_75t_L g805 ( 
.A1(n_747),
.A2(n_595),
.B(n_605),
.C(n_601),
.Y(n_805)
);

AOI21xp33_ASAP7_75t_L g806 ( 
.A1(n_690),
.A2(n_606),
.B(n_605),
.Y(n_806)
);

OAI21xp5_ASAP7_75t_L g807 ( 
.A1(n_703),
.A2(n_532),
.B(n_533),
.Y(n_807)
);

AOI22xp5_ASAP7_75t_L g808 ( 
.A1(n_618),
.A2(n_526),
.B1(n_594),
.B2(n_577),
.Y(n_808)
);

AOI21xp5_ASAP7_75t_L g809 ( 
.A1(n_623),
.A2(n_555),
.B(n_532),
.Y(n_809)
);

INVx1_ASAP7_75t_L g810 ( 
.A(n_754),
.Y(n_810)
);

BUFx8_ASAP7_75t_L g811 ( 
.A(n_667),
.Y(n_811)
);

NAND2xp5_ASAP7_75t_L g812 ( 
.A(n_671),
.B(n_526),
.Y(n_812)
);

NAND2xp5_ASAP7_75t_L g813 ( 
.A(n_671),
.B(n_526),
.Y(n_813)
);

CKINVDCx10_ASAP7_75t_R g814 ( 
.A(n_667),
.Y(n_814)
);

A2O1A1Ixp33_ASAP7_75t_L g815 ( 
.A1(n_672),
.A2(n_601),
.B(n_597),
.C(n_533),
.Y(n_815)
);

AOI21xp5_ASAP7_75t_L g816 ( 
.A1(n_623),
.A2(n_555),
.B(n_512),
.Y(n_816)
);

INVx4_ASAP7_75t_L g817 ( 
.A(n_634),
.Y(n_817)
);

O2A1O1Ixp33_ASAP7_75t_L g818 ( 
.A1(n_747),
.A2(n_597),
.B(n_578),
.C(n_534),
.Y(n_818)
);

NAND2xp5_ASAP7_75t_SL g819 ( 
.A(n_701),
.B(n_512),
.Y(n_819)
);

NOR2x1_ASAP7_75t_R g820 ( 
.A(n_612),
.B(n_742),
.Y(n_820)
);

NAND2xp5_ASAP7_75t_L g821 ( 
.A(n_631),
.B(n_512),
.Y(n_821)
);

NAND2xp5_ASAP7_75t_SL g822 ( 
.A(n_642),
.B(n_512),
.Y(n_822)
);

NAND2xp5_ASAP7_75t_L g823 ( 
.A(n_722),
.B(n_549),
.Y(n_823)
);

CKINVDCx6p67_ASAP7_75t_R g824 ( 
.A(n_725),
.Y(n_824)
);

NOR2x1_ASAP7_75t_L g825 ( 
.A(n_636),
.B(n_534),
.Y(n_825)
);

NOR3xp33_ASAP7_75t_L g826 ( 
.A(n_724),
.B(n_541),
.C(n_578),
.Y(n_826)
);

AOI22xp33_ASAP7_75t_L g827 ( 
.A1(n_675),
.A2(n_497),
.B1(n_549),
.B2(n_568),
.Y(n_827)
);

OAI21xp5_ASAP7_75t_L g828 ( 
.A1(n_626),
.A2(n_549),
.B(n_568),
.Y(n_828)
);

A2O1A1Ixp33_ASAP7_75t_L g829 ( 
.A1(n_690),
.A2(n_549),
.B(n_568),
.C(n_497),
.Y(n_829)
);

NAND2xp5_ASAP7_75t_SL g830 ( 
.A(n_763),
.B(n_549),
.Y(n_830)
);

AND2x2_ASAP7_75t_L g831 ( 
.A(n_715),
.B(n_497),
.Y(n_831)
);

AOI21xp5_ASAP7_75t_L g832 ( 
.A1(n_626),
.A2(n_637),
.B(n_632),
.Y(n_832)
);

AOI21xp5_ASAP7_75t_L g833 ( 
.A1(n_632),
.A2(n_568),
.B(n_497),
.Y(n_833)
);

OAI21xp33_ASAP7_75t_L g834 ( 
.A1(n_645),
.A2(n_695),
.B(n_691),
.Y(n_834)
);

A2O1A1Ixp33_ASAP7_75t_L g835 ( 
.A1(n_691),
.A2(n_695),
.B(n_621),
.C(n_618),
.Y(n_835)
);

A2O1A1Ixp33_ASAP7_75t_L g836 ( 
.A1(n_621),
.A2(n_568),
.B(n_729),
.C(n_721),
.Y(n_836)
);

BUFx6f_ASAP7_75t_L g837 ( 
.A(n_745),
.Y(n_837)
);

INVx1_ASAP7_75t_L g838 ( 
.A(n_775),
.Y(n_838)
);

NOR2xp33_ASAP7_75t_R g839 ( 
.A(n_725),
.B(n_677),
.Y(n_839)
);

INVx1_ASAP7_75t_L g840 ( 
.A(n_758),
.Y(n_840)
);

AND2x2_ASAP7_75t_L g841 ( 
.A(n_718),
.B(n_689),
.Y(n_841)
);

AOI21xp5_ASAP7_75t_L g842 ( 
.A1(n_637),
.A2(n_647),
.B(n_676),
.Y(n_842)
);

OAI22xp5_ASAP7_75t_L g843 ( 
.A1(n_652),
.A2(n_683),
.B1(n_633),
.B2(n_749),
.Y(n_843)
);

NAND2xp5_ASAP7_75t_L g844 ( 
.A(n_644),
.B(n_655),
.Y(n_844)
);

AOI21xp5_ASAP7_75t_L g845 ( 
.A1(n_647),
.A2(n_663),
.B(n_673),
.Y(n_845)
);

INVx2_ASAP7_75t_L g846 ( 
.A(n_755),
.Y(n_846)
);

AND2x4_ASAP7_75t_L g847 ( 
.A(n_636),
.B(n_705),
.Y(n_847)
);

NAND2xp5_ASAP7_75t_L g848 ( 
.A(n_710),
.B(n_720),
.Y(n_848)
);

INVx2_ASAP7_75t_L g849 ( 
.A(n_708),
.Y(n_849)
);

AOI21xp5_ASAP7_75t_L g850 ( 
.A1(n_663),
.A2(n_673),
.B(n_676),
.Y(n_850)
);

OAI22xp5_ASAP7_75t_L g851 ( 
.A1(n_652),
.A2(n_633),
.B1(n_749),
.B2(n_734),
.Y(n_851)
);

NAND2xp5_ASAP7_75t_L g852 ( 
.A(n_761),
.B(n_769),
.Y(n_852)
);

NAND2xp5_ASAP7_75t_L g853 ( 
.A(n_619),
.B(n_624),
.Y(n_853)
);

AOI21xp5_ASAP7_75t_L g854 ( 
.A1(n_678),
.A2(n_688),
.B(n_773),
.Y(n_854)
);

NAND2xp5_ASAP7_75t_L g855 ( 
.A(n_762),
.B(n_614),
.Y(n_855)
);

OAI21x1_ASAP7_75t_L g856 ( 
.A1(n_766),
.A2(n_607),
.B(n_678),
.Y(n_856)
);

NAND2xp5_ASAP7_75t_L g857 ( 
.A(n_617),
.B(n_638),
.Y(n_857)
);

AOI21xp5_ASAP7_75t_L g858 ( 
.A1(n_688),
.A2(n_698),
.B(n_651),
.Y(n_858)
);

AOI21xp5_ASAP7_75t_L g859 ( 
.A1(n_625),
.A2(n_670),
.B(n_635),
.Y(n_859)
);

INVx1_ASAP7_75t_L g860 ( 
.A(n_609),
.Y(n_860)
);

AOI21xp5_ASAP7_75t_L g861 ( 
.A1(n_627),
.A2(n_662),
.B(n_658),
.Y(n_861)
);

INVx1_ASAP7_75t_SL g862 ( 
.A(n_668),
.Y(n_862)
);

AOI21xp5_ASAP7_75t_L g863 ( 
.A1(n_654),
.A2(n_753),
.B(n_751),
.Y(n_863)
);

INVx4_ASAP7_75t_L g864 ( 
.A(n_634),
.Y(n_864)
);

BUFx8_ASAP7_75t_L g865 ( 
.A(n_693),
.Y(n_865)
);

AOI21xp5_ASAP7_75t_L g866 ( 
.A1(n_607),
.A2(n_768),
.B(n_774),
.Y(n_866)
);

INVx2_ASAP7_75t_L g867 ( 
.A(n_736),
.Y(n_867)
);

O2A1O1Ixp33_ASAP7_75t_SL g868 ( 
.A1(n_774),
.A2(n_709),
.B(n_750),
.C(n_757),
.Y(n_868)
);

NAND2xp5_ASAP7_75t_L g869 ( 
.A(n_665),
.B(n_699),
.Y(n_869)
);

AOI21x1_ASAP7_75t_L g870 ( 
.A1(n_759),
.A2(n_770),
.B(n_764),
.Y(n_870)
);

AOI21xp5_ASAP7_75t_L g871 ( 
.A1(n_684),
.A2(n_723),
.B(n_727),
.Y(n_871)
);

NAND2xp5_ASAP7_75t_L g872 ( 
.A(n_699),
.B(n_712),
.Y(n_872)
);

NAND2xp5_ASAP7_75t_L g873 ( 
.A(n_712),
.B(n_641),
.Y(n_873)
);

AOI21xp5_ASAP7_75t_L g874 ( 
.A1(n_692),
.A2(n_719),
.B(n_731),
.Y(n_874)
);

AOI21xp5_ASAP7_75t_L g875 ( 
.A1(n_629),
.A2(n_640),
.B(n_704),
.Y(n_875)
);

AND2x2_ASAP7_75t_L g876 ( 
.A(n_666),
.B(n_661),
.Y(n_876)
);

NOR2xp33_ASAP7_75t_L g877 ( 
.A(n_674),
.B(n_680),
.Y(n_877)
);

AOI21xp5_ASAP7_75t_L g878 ( 
.A1(n_660),
.A2(n_681),
.B(n_694),
.Y(n_878)
);

INVx1_ASAP7_75t_L g879 ( 
.A(n_682),
.Y(n_879)
);

INVx2_ASAP7_75t_L g880 ( 
.A(n_739),
.Y(n_880)
);

NOR2xp33_ASAP7_75t_L g881 ( 
.A(n_674),
.B(n_680),
.Y(n_881)
);

INVx1_ASAP7_75t_L g882 ( 
.A(n_697),
.Y(n_882)
);

INVx1_ASAP7_75t_SL g883 ( 
.A(n_771),
.Y(n_883)
);

NAND2x1p5_ASAP7_75t_L g884 ( 
.A(n_745),
.B(n_726),
.Y(n_884)
);

INVx1_ASAP7_75t_L g885 ( 
.A(n_746),
.Y(n_885)
);

INVx2_ASAP7_75t_L g886 ( 
.A(n_643),
.Y(n_886)
);

INVx2_ASAP7_75t_L g887 ( 
.A(n_737),
.Y(n_887)
);

NAND2xp5_ASAP7_75t_L g888 ( 
.A(n_608),
.B(n_738),
.Y(n_888)
);

CKINVDCx16_ASAP7_75t_R g889 ( 
.A(n_728),
.Y(n_889)
);

INVx2_ASAP7_75t_L g890 ( 
.A(n_740),
.Y(n_890)
);

AOI21xp5_ASAP7_75t_L g891 ( 
.A1(n_687),
.A2(n_732),
.B(n_657),
.Y(n_891)
);

AOI21xp5_ASAP7_75t_L g892 ( 
.A1(n_648),
.A2(n_659),
.B(n_757),
.Y(n_892)
);

INVx4_ASAP7_75t_L g893 ( 
.A(n_634),
.Y(n_893)
);

NAND2xp5_ASAP7_75t_L g894 ( 
.A(n_685),
.B(n_608),
.Y(n_894)
);

INVx1_ASAP7_75t_L g895 ( 
.A(n_728),
.Y(n_895)
);

OAI21xp33_ASAP7_75t_L g896 ( 
.A1(n_685),
.A2(n_700),
.B(n_639),
.Y(n_896)
);

INVx1_ASAP7_75t_L g897 ( 
.A(n_728),
.Y(n_897)
);

INVx4_ASAP7_75t_L g898 ( 
.A(n_745),
.Y(n_898)
);

AOI22xp33_ASAP7_75t_SL g899 ( 
.A1(n_721),
.A2(n_729),
.B1(n_744),
.B2(n_696),
.Y(n_899)
);

AOI21xp5_ASAP7_75t_L g900 ( 
.A1(n_750),
.A2(n_743),
.B(n_735),
.Y(n_900)
);

BUFx12f_ASAP7_75t_L g901 ( 
.A(n_679),
.Y(n_901)
);

NOR2x1_ASAP7_75t_L g902 ( 
.A(n_760),
.B(n_679),
.Y(n_902)
);

NAND2xp5_ASAP7_75t_L g903 ( 
.A(n_744),
.B(n_649),
.Y(n_903)
);

O2A1O1Ixp33_ASAP7_75t_L g904 ( 
.A1(n_733),
.A2(n_686),
.B(n_630),
.C(n_760),
.Y(n_904)
);

A2O1A1Ixp33_ASAP7_75t_L g905 ( 
.A1(n_622),
.A2(n_646),
.B(n_653),
.C(n_765),
.Y(n_905)
);

NOR2xp33_ASAP7_75t_L g906 ( 
.A(n_679),
.B(n_656),
.Y(n_906)
);

INVx2_ASAP7_75t_L g907 ( 
.A(n_745),
.Y(n_907)
);

BUFx2_ASAP7_75t_L g908 ( 
.A(n_717),
.Y(n_908)
);

OAI21xp33_ASAP7_75t_L g909 ( 
.A1(n_664),
.A2(n_702),
.B(n_760),
.Y(n_909)
);

BUFx6f_ASAP7_75t_L g910 ( 
.A(n_714),
.Y(n_910)
);

NOR2xp67_ASAP7_75t_L g911 ( 
.A(n_765),
.B(n_756),
.Y(n_911)
);

INVx1_ASAP7_75t_L g912 ( 
.A(n_714),
.Y(n_912)
);

NAND2xp5_ASAP7_75t_L g913 ( 
.A(n_714),
.B(n_705),
.Y(n_913)
);

A2O1A1Ixp33_ASAP7_75t_L g914 ( 
.A1(n_772),
.A2(n_669),
.B(n_459),
.C(n_615),
.Y(n_914)
);

AOI21x1_ASAP7_75t_L g915 ( 
.A1(n_705),
.A2(n_626),
.B(n_623),
.Y(n_915)
);

NOR2xp33_ASAP7_75t_R g916 ( 
.A(n_714),
.B(n_536),
.Y(n_916)
);

INVx2_ASAP7_75t_L g917 ( 
.A(n_748),
.Y(n_917)
);

INVx2_ASAP7_75t_L g918 ( 
.A(n_748),
.Y(n_918)
);

AOI21xp5_ASAP7_75t_L g919 ( 
.A1(n_650),
.A2(n_628),
.B(n_598),
.Y(n_919)
);

OAI22xp5_ASAP7_75t_L g920 ( 
.A1(n_669),
.A2(n_459),
.B1(n_652),
.B2(n_441),
.Y(n_920)
);

AOI21xp5_ASAP7_75t_L g921 ( 
.A1(n_650),
.A2(n_628),
.B(n_598),
.Y(n_921)
);

OAI22xp5_ASAP7_75t_L g922 ( 
.A1(n_669),
.A2(n_459),
.B1(n_652),
.B2(n_441),
.Y(n_922)
);

INVx1_ASAP7_75t_L g923 ( 
.A(n_706),
.Y(n_923)
);

NAND2xp5_ASAP7_75t_SL g924 ( 
.A(n_669),
.B(n_599),
.Y(n_924)
);

AO21x1_ASAP7_75t_L g925 ( 
.A1(n_623),
.A2(n_459),
.B(n_626),
.Y(n_925)
);

NAND2xp5_ASAP7_75t_L g926 ( 
.A(n_615),
.B(n_669),
.Y(n_926)
);

INVx2_ASAP7_75t_SL g927 ( 
.A(n_741),
.Y(n_927)
);

OAI21xp5_ASAP7_75t_L g928 ( 
.A1(n_650),
.A2(n_558),
.B(n_470),
.Y(n_928)
);

INVx4_ASAP7_75t_L g929 ( 
.A(n_634),
.Y(n_929)
);

INVx3_ASAP7_75t_L g930 ( 
.A(n_745),
.Y(n_930)
);

A2O1A1Ixp33_ASAP7_75t_L g931 ( 
.A1(n_669),
.A2(n_459),
.B(n_615),
.C(n_672),
.Y(n_931)
);

NOR2xp33_ASAP7_75t_L g932 ( 
.A(n_620),
.B(n_324),
.Y(n_932)
);

INVx2_ASAP7_75t_SL g933 ( 
.A(n_741),
.Y(n_933)
);

AND2x2_ASAP7_75t_L g934 ( 
.A(n_620),
.B(n_715),
.Y(n_934)
);

NAND2xp5_ASAP7_75t_L g935 ( 
.A(n_615),
.B(n_669),
.Y(n_935)
);

A2O1A1Ixp33_ASAP7_75t_L g936 ( 
.A1(n_669),
.A2(n_459),
.B(n_615),
.C(n_672),
.Y(n_936)
);

AOI21xp5_ASAP7_75t_L g937 ( 
.A1(n_650),
.A2(n_628),
.B(n_598),
.Y(n_937)
);

AOI22xp5_ASAP7_75t_L g938 ( 
.A1(n_615),
.A2(n_669),
.B1(n_448),
.B2(n_465),
.Y(n_938)
);

NAND2xp5_ASAP7_75t_L g939 ( 
.A(n_615),
.B(n_669),
.Y(n_939)
);

NOR2xp33_ASAP7_75t_L g940 ( 
.A(n_620),
.B(n_324),
.Y(n_940)
);

NAND2xp5_ASAP7_75t_L g941 ( 
.A(n_615),
.B(n_669),
.Y(n_941)
);

NAND2xp5_ASAP7_75t_L g942 ( 
.A(n_615),
.B(n_669),
.Y(n_942)
);

AOI21xp5_ASAP7_75t_L g943 ( 
.A1(n_650),
.A2(n_628),
.B(n_598),
.Y(n_943)
);

NOR2xp33_ASAP7_75t_L g944 ( 
.A(n_620),
.B(n_324),
.Y(n_944)
);

NAND2xp5_ASAP7_75t_L g945 ( 
.A(n_615),
.B(n_669),
.Y(n_945)
);

BUFx6f_ASAP7_75t_L g946 ( 
.A(n_745),
.Y(n_946)
);

AOI21xp5_ASAP7_75t_L g947 ( 
.A1(n_650),
.A2(n_628),
.B(n_598),
.Y(n_947)
);

NAND2xp5_ASAP7_75t_L g948 ( 
.A(n_669),
.B(n_583),
.Y(n_948)
);

NAND2xp5_ASAP7_75t_L g949 ( 
.A(n_669),
.B(n_583),
.Y(n_949)
);

BUFx6f_ASAP7_75t_L g950 ( 
.A(n_745),
.Y(n_950)
);

AOI21x1_ASAP7_75t_L g951 ( 
.A1(n_623),
.A2(n_632),
.B(n_626),
.Y(n_951)
);

OAI22xp5_ASAP7_75t_L g952 ( 
.A1(n_669),
.A2(n_459),
.B1(n_652),
.B2(n_441),
.Y(n_952)
);

AOI21xp5_ASAP7_75t_L g953 ( 
.A1(n_650),
.A2(n_628),
.B(n_598),
.Y(n_953)
);

INVx1_ASAP7_75t_L g954 ( 
.A(n_706),
.Y(n_954)
);

A2O1A1Ixp33_ASAP7_75t_L g955 ( 
.A1(n_669),
.A2(n_459),
.B(n_615),
.C(n_672),
.Y(n_955)
);

NOR2xp33_ASAP7_75t_L g956 ( 
.A(n_620),
.B(n_324),
.Y(n_956)
);

INVx1_ASAP7_75t_L g957 ( 
.A(n_706),
.Y(n_957)
);

OAI21xp33_ASAP7_75t_L g958 ( 
.A1(n_615),
.A2(n_465),
.B(n_521),
.Y(n_958)
);

NAND2xp5_ASAP7_75t_L g959 ( 
.A(n_615),
.B(n_669),
.Y(n_959)
);

INVx1_ASAP7_75t_L g960 ( 
.A(n_706),
.Y(n_960)
);

OAI21x1_ASAP7_75t_L g961 ( 
.A1(n_650),
.A2(n_598),
.B(n_623),
.Y(n_961)
);

NAND2xp5_ASAP7_75t_L g962 ( 
.A(n_615),
.B(n_669),
.Y(n_962)
);

NAND2xp5_ASAP7_75t_L g963 ( 
.A(n_669),
.B(n_583),
.Y(n_963)
);

OAI21xp5_ASAP7_75t_L g964 ( 
.A1(n_650),
.A2(n_558),
.B(n_470),
.Y(n_964)
);

INVx2_ASAP7_75t_L g965 ( 
.A(n_748),
.Y(n_965)
);

OAI21x1_ASAP7_75t_L g966 ( 
.A1(n_961),
.A2(n_856),
.B(n_866),
.Y(n_966)
);

INVx1_ASAP7_75t_L g967 ( 
.A(n_781),
.Y(n_967)
);

INVx1_ASAP7_75t_L g968 ( 
.A(n_797),
.Y(n_968)
);

NAND2xp5_ASAP7_75t_L g969 ( 
.A(n_926),
.B(n_935),
.Y(n_969)
);

OAI22xp5_ASAP7_75t_L g970 ( 
.A1(n_939),
.A2(n_962),
.B1(n_945),
.B2(n_959),
.Y(n_970)
);

NAND2xp5_ASAP7_75t_L g971 ( 
.A(n_941),
.B(n_942),
.Y(n_971)
);

NAND3xp33_ASAP7_75t_L g972 ( 
.A(n_938),
.B(n_958),
.C(n_881),
.Y(n_972)
);

NAND2x1_ASAP7_75t_L g973 ( 
.A(n_898),
.B(n_930),
.Y(n_973)
);

BUFx2_ASAP7_75t_L g974 ( 
.A(n_780),
.Y(n_974)
);

BUFx2_ASAP7_75t_SL g975 ( 
.A(n_791),
.Y(n_975)
);

NAND2xp5_ASAP7_75t_L g976 ( 
.A(n_948),
.B(n_949),
.Y(n_976)
);

NAND2xp5_ASAP7_75t_SL g977 ( 
.A(n_877),
.B(n_931),
.Y(n_977)
);

OAI21x1_ASAP7_75t_L g978 ( 
.A1(n_951),
.A2(n_832),
.B(n_863),
.Y(n_978)
);

OAI21xp5_ASAP7_75t_L g979 ( 
.A1(n_936),
.A2(n_955),
.B(n_914),
.Y(n_979)
);

BUFx6f_ASAP7_75t_L g980 ( 
.A(n_910),
.Y(n_980)
);

O2A1O1Ixp33_ASAP7_75t_SL g981 ( 
.A1(n_835),
.A2(n_872),
.B(n_963),
.C(n_905),
.Y(n_981)
);

NOR2xp67_ASAP7_75t_L g982 ( 
.A(n_927),
.B(n_933),
.Y(n_982)
);

NOR2x1_ASAP7_75t_SL g983 ( 
.A(n_910),
.B(n_963),
.Y(n_983)
);

AO31x2_ASAP7_75t_L g984 ( 
.A1(n_925),
.A2(n_843),
.A3(n_829),
.B(n_892),
.Y(n_984)
);

AOI21xp5_ASAP7_75t_L g985 ( 
.A1(n_868),
.A2(n_855),
.B(n_874),
.Y(n_985)
);

BUFx2_ASAP7_75t_SL g986 ( 
.A(n_794),
.Y(n_986)
);

AO31x2_ASAP7_75t_L g987 ( 
.A1(n_843),
.A2(n_815),
.A3(n_888),
.B(n_952),
.Y(n_987)
);

OAI21xp5_ASAP7_75t_L g988 ( 
.A1(n_920),
.A2(n_952),
.B(n_922),
.Y(n_988)
);

AOI21x1_ASAP7_75t_L g989 ( 
.A1(n_900),
.A2(n_915),
.B(n_911),
.Y(n_989)
);

BUFx2_ASAP7_75t_L g990 ( 
.A(n_862),
.Y(n_990)
);

NAND2xp5_ASAP7_75t_SL g991 ( 
.A(n_920),
.B(n_922),
.Y(n_991)
);

AOI21xp5_ASAP7_75t_L g992 ( 
.A1(n_855),
.A2(n_921),
.B(n_919),
.Y(n_992)
);

AOI221x1_ASAP7_75t_L g993 ( 
.A1(n_834),
.A2(n_896),
.B1(n_851),
.B2(n_894),
.C(n_909),
.Y(n_993)
);

OAI22xp5_ASAP7_75t_L g994 ( 
.A1(n_778),
.A2(n_873),
.B1(n_777),
.B2(n_869),
.Y(n_994)
);

A2O1A1Ixp33_ASAP7_75t_L g995 ( 
.A1(n_779),
.A2(n_903),
.B(n_888),
.C(n_891),
.Y(n_995)
);

OAI21xp5_ASAP7_75t_L g996 ( 
.A1(n_799),
.A2(n_845),
.B(n_842),
.Y(n_996)
);

AOI21x1_ASAP7_75t_L g997 ( 
.A1(n_854),
.A2(n_830),
.B(n_937),
.Y(n_997)
);

OAI21xp5_ASAP7_75t_L g998 ( 
.A1(n_799),
.A2(n_928),
.B(n_964),
.Y(n_998)
);

NAND2xp5_ASAP7_75t_L g999 ( 
.A(n_886),
.B(n_934),
.Y(n_999)
);

NAND2xp5_ASAP7_75t_SL g1000 ( 
.A(n_928),
.B(n_964),
.Y(n_1000)
);

AOI21x1_ASAP7_75t_L g1001 ( 
.A1(n_943),
.A2(n_953),
.B(n_947),
.Y(n_1001)
);

INVx3_ASAP7_75t_L g1002 ( 
.A(n_817),
.Y(n_1002)
);

A2O1A1Ixp33_ASAP7_75t_L g1003 ( 
.A1(n_782),
.A2(n_787),
.B(n_836),
.C(n_899),
.Y(n_1003)
);

A2O1A1Ixp33_ASAP7_75t_L g1004 ( 
.A1(n_851),
.A2(n_848),
.B(n_904),
.C(n_924),
.Y(n_1004)
);

AO31x2_ASAP7_75t_L g1005 ( 
.A1(n_853),
.A2(n_809),
.A3(n_802),
.B(n_800),
.Y(n_1005)
);

BUFx6f_ASAP7_75t_L g1006 ( 
.A(n_910),
.Y(n_1006)
);

NAND2xp5_ASAP7_75t_L g1007 ( 
.A(n_876),
.B(n_848),
.Y(n_1007)
);

BUFx6f_ASAP7_75t_L g1008 ( 
.A(n_837),
.Y(n_1008)
);

AOI21xp5_ASAP7_75t_L g1009 ( 
.A1(n_801),
.A2(n_813),
.B(n_812),
.Y(n_1009)
);

NAND2xp5_ASAP7_75t_L g1010 ( 
.A(n_844),
.B(n_932),
.Y(n_1010)
);

OAI22xp5_ASAP7_75t_L g1011 ( 
.A1(n_852),
.A2(n_956),
.B1(n_940),
.B2(n_944),
.Y(n_1011)
);

OAI21xp5_ASAP7_75t_L g1012 ( 
.A1(n_850),
.A2(n_807),
.B(n_878),
.Y(n_1012)
);

BUFx2_ASAP7_75t_L g1013 ( 
.A(n_839),
.Y(n_1013)
);

BUFx3_ASAP7_75t_L g1014 ( 
.A(n_811),
.Y(n_1014)
);

A2O1A1Ixp33_ASAP7_75t_L g1015 ( 
.A1(n_890),
.A2(n_906),
.B(n_857),
.C(n_853),
.Y(n_1015)
);

AOI21xp5_ASAP7_75t_L g1016 ( 
.A1(n_871),
.A2(n_795),
.B(n_792),
.Y(n_1016)
);

OAI21x1_ASAP7_75t_L g1017 ( 
.A1(n_807),
.A2(n_870),
.B(n_790),
.Y(n_1017)
);

BUFx2_ASAP7_75t_L g1018 ( 
.A(n_916),
.Y(n_1018)
);

AND2x2_ASAP7_75t_L g1019 ( 
.A(n_841),
.B(n_889),
.Y(n_1019)
);

OAI21xp5_ASAP7_75t_L g1020 ( 
.A1(n_875),
.A2(n_798),
.B(n_859),
.Y(n_1020)
);

NAND2xp33_ASAP7_75t_L g1021 ( 
.A(n_798),
.B(n_912),
.Y(n_1021)
);

AO31x2_ASAP7_75t_L g1022 ( 
.A1(n_887),
.A2(n_816),
.A3(n_857),
.B(n_858),
.Y(n_1022)
);

OAI21xp5_ASAP7_75t_L g1023 ( 
.A1(n_861),
.A2(n_805),
.B(n_788),
.Y(n_1023)
);

NAND2xp5_ASAP7_75t_L g1024 ( 
.A(n_786),
.B(n_923),
.Y(n_1024)
);

OAI21x1_ASAP7_75t_L g1025 ( 
.A1(n_828),
.A2(n_833),
.B(n_913),
.Y(n_1025)
);

BUFx10_ASAP7_75t_L g1026 ( 
.A(n_803),
.Y(n_1026)
);

NAND2xp5_ASAP7_75t_L g1027 ( 
.A(n_954),
.B(n_960),
.Y(n_1027)
);

NAND2xp5_ASAP7_75t_L g1028 ( 
.A(n_957),
.B(n_852),
.Y(n_1028)
);

NAND2xp5_ASAP7_75t_L g1029 ( 
.A(n_804),
.B(n_840),
.Y(n_1029)
);

NAND2xp5_ASAP7_75t_L g1030 ( 
.A(n_810),
.B(n_838),
.Y(n_1030)
);

INVx2_ASAP7_75t_L g1031 ( 
.A(n_783),
.Y(n_1031)
);

OAI21xp5_ASAP7_75t_L g1032 ( 
.A1(n_788),
.A2(n_806),
.B(n_789),
.Y(n_1032)
);

AOI21xp5_ASAP7_75t_L g1033 ( 
.A1(n_828),
.A2(n_823),
.B(n_789),
.Y(n_1033)
);

O2A1O1Ixp33_ASAP7_75t_L g1034 ( 
.A1(n_806),
.A2(n_860),
.B(n_879),
.C(n_882),
.Y(n_1034)
);

AND2x2_ASAP7_75t_L g1035 ( 
.A(n_847),
.B(n_824),
.Y(n_1035)
);

OAI21xp5_ASAP7_75t_L g1036 ( 
.A1(n_818),
.A2(n_821),
.B(n_823),
.Y(n_1036)
);

NAND2x1p5_ASAP7_75t_L g1037 ( 
.A(n_817),
.B(n_929),
.Y(n_1037)
);

AO21x2_ASAP7_75t_L g1038 ( 
.A1(n_808),
.A2(n_822),
.B(n_965),
.Y(n_1038)
);

INVx5_ASAP7_75t_L g1039 ( 
.A(n_864),
.Y(n_1039)
);

AOI21x1_ASAP7_75t_SL g1040 ( 
.A1(n_796),
.A2(n_803),
.B(n_831),
.Y(n_1040)
);

INVx1_ASAP7_75t_L g1041 ( 
.A(n_885),
.Y(n_1041)
);

NAND2xp5_ASAP7_75t_L g1042 ( 
.A(n_902),
.B(n_929),
.Y(n_1042)
);

AND2x2_ASAP7_75t_L g1043 ( 
.A(n_847),
.B(n_793),
.Y(n_1043)
);

AOI221xp5_ASAP7_75t_SL g1044 ( 
.A1(n_895),
.A2(n_897),
.B1(n_908),
.B2(n_827),
.C(n_819),
.Y(n_1044)
);

AND2x2_ASAP7_75t_L g1045 ( 
.A(n_826),
.B(n_901),
.Y(n_1045)
);

AOI21xp33_ASAP7_75t_L g1046 ( 
.A1(n_849),
.A2(n_867),
.B(n_880),
.Y(n_1046)
);

OAI22xp5_ASAP7_75t_L g1047 ( 
.A1(n_884),
.A2(n_785),
.B1(n_864),
.B2(n_893),
.Y(n_1047)
);

NAND2xp5_ASAP7_75t_L g1048 ( 
.A(n_893),
.B(n_784),
.Y(n_1048)
);

INVx2_ASAP7_75t_L g1049 ( 
.A(n_846),
.Y(n_1049)
);

OAI21x1_ASAP7_75t_L g1050 ( 
.A1(n_917),
.A2(n_918),
.B(n_825),
.Y(n_1050)
);

AOI21x1_ASAP7_75t_L g1051 ( 
.A1(n_907),
.A2(n_796),
.B(n_884),
.Y(n_1051)
);

AOI21xp5_ASAP7_75t_L g1052 ( 
.A1(n_930),
.A2(n_950),
.B(n_946),
.Y(n_1052)
);

OAI21xp5_ASAP7_75t_L g1053 ( 
.A1(n_898),
.A2(n_796),
.B(n_837),
.Y(n_1053)
);

AOI21xp33_ASAP7_75t_L g1054 ( 
.A1(n_837),
.A2(n_946),
.B(n_950),
.Y(n_1054)
);

OAI21x1_ASAP7_75t_L g1055 ( 
.A1(n_946),
.A2(n_950),
.B(n_811),
.Y(n_1055)
);

A2O1A1Ixp33_ASAP7_75t_L g1056 ( 
.A1(n_883),
.A2(n_814),
.B(n_865),
.C(n_820),
.Y(n_1056)
);

AOI221xp5_ASAP7_75t_L g1057 ( 
.A1(n_865),
.A2(n_935),
.B1(n_941),
.B2(n_939),
.C(n_926),
.Y(n_1057)
);

OAI21x1_ASAP7_75t_L g1058 ( 
.A1(n_961),
.A2(n_856),
.B(n_866),
.Y(n_1058)
);

OAI21x1_ASAP7_75t_L g1059 ( 
.A1(n_961),
.A2(n_856),
.B(n_866),
.Y(n_1059)
);

OA21x2_ASAP7_75t_L g1060 ( 
.A1(n_807),
.A2(n_961),
.B(n_914),
.Y(n_1060)
);

AOI21xp5_ASAP7_75t_L g1061 ( 
.A1(n_926),
.A2(n_939),
.B(n_935),
.Y(n_1061)
);

NAND2xp5_ASAP7_75t_L g1062 ( 
.A(n_926),
.B(n_935),
.Y(n_1062)
);

INVx3_ASAP7_75t_L g1063 ( 
.A(n_817),
.Y(n_1063)
);

NOR2xp67_ASAP7_75t_SL g1064 ( 
.A(n_926),
.B(n_599),
.Y(n_1064)
);

NAND2xp5_ASAP7_75t_L g1065 ( 
.A(n_926),
.B(n_935),
.Y(n_1065)
);

AND2x4_ASAP7_75t_L g1066 ( 
.A(n_817),
.B(n_864),
.Y(n_1066)
);

NAND2xp5_ASAP7_75t_L g1067 ( 
.A(n_926),
.B(n_935),
.Y(n_1067)
);

OAI21x1_ASAP7_75t_L g1068 ( 
.A1(n_961),
.A2(n_856),
.B(n_866),
.Y(n_1068)
);

A2O1A1Ixp33_ASAP7_75t_L g1069 ( 
.A1(n_926),
.A2(n_939),
.B(n_941),
.C(n_935),
.Y(n_1069)
);

OAI21x1_ASAP7_75t_L g1070 ( 
.A1(n_961),
.A2(n_921),
.B(n_919),
.Y(n_1070)
);

NAND2xp5_ASAP7_75t_L g1071 ( 
.A(n_926),
.B(n_935),
.Y(n_1071)
);

OAI21x1_ASAP7_75t_L g1072 ( 
.A1(n_961),
.A2(n_921),
.B(n_919),
.Y(n_1072)
);

OAI22x1_ASAP7_75t_L g1073 ( 
.A1(n_938),
.A2(n_537),
.B1(n_881),
.B2(n_877),
.Y(n_1073)
);

INVx1_ASAP7_75t_L g1074 ( 
.A(n_781),
.Y(n_1074)
);

AO21x1_ASAP7_75t_L g1075 ( 
.A1(n_877),
.A2(n_881),
.B(n_926),
.Y(n_1075)
);

AOI21x1_ASAP7_75t_L g1076 ( 
.A1(n_900),
.A2(n_866),
.B(n_951),
.Y(n_1076)
);

BUFx2_ASAP7_75t_L g1077 ( 
.A(n_780),
.Y(n_1077)
);

NOR2x1_ASAP7_75t_L g1078 ( 
.A(n_794),
.B(n_599),
.Y(n_1078)
);

OAI21x1_ASAP7_75t_L g1079 ( 
.A1(n_961),
.A2(n_921),
.B(n_919),
.Y(n_1079)
);

A2O1A1Ixp33_ASAP7_75t_SL g1080 ( 
.A1(n_877),
.A2(n_881),
.B(n_938),
.C(n_615),
.Y(n_1080)
);

INVx2_ASAP7_75t_L g1081 ( 
.A(n_776),
.Y(n_1081)
);

INVx2_ASAP7_75t_SL g1082 ( 
.A(n_794),
.Y(n_1082)
);

BUFx2_ASAP7_75t_L g1083 ( 
.A(n_780),
.Y(n_1083)
);

NAND2xp5_ASAP7_75t_L g1084 ( 
.A(n_926),
.B(n_935),
.Y(n_1084)
);

INVx3_ASAP7_75t_L g1085 ( 
.A(n_817),
.Y(n_1085)
);

OA21x2_ASAP7_75t_L g1086 ( 
.A1(n_807),
.A2(n_961),
.B(n_914),
.Y(n_1086)
);

INVx3_ASAP7_75t_L g1087 ( 
.A(n_817),
.Y(n_1087)
);

NAND2xp5_ASAP7_75t_L g1088 ( 
.A(n_926),
.B(n_935),
.Y(n_1088)
);

AND2x4_ASAP7_75t_L g1089 ( 
.A(n_817),
.B(n_864),
.Y(n_1089)
);

NAND2xp5_ASAP7_75t_L g1090 ( 
.A(n_926),
.B(n_935),
.Y(n_1090)
);

INVx1_ASAP7_75t_L g1091 ( 
.A(n_781),
.Y(n_1091)
);

NAND2xp5_ASAP7_75t_L g1092 ( 
.A(n_926),
.B(n_935),
.Y(n_1092)
);

OAI22x1_ASAP7_75t_L g1093 ( 
.A1(n_938),
.A2(n_537),
.B1(n_881),
.B2(n_877),
.Y(n_1093)
);

OAI21x1_ASAP7_75t_L g1094 ( 
.A1(n_961),
.A2(n_856),
.B(n_866),
.Y(n_1094)
);

AO21x1_ASAP7_75t_L g1095 ( 
.A1(n_877),
.A2(n_881),
.B(n_926),
.Y(n_1095)
);

NOR2xp33_ASAP7_75t_L g1096 ( 
.A(n_926),
.B(n_935),
.Y(n_1096)
);

OAI21x1_ASAP7_75t_L g1097 ( 
.A1(n_961),
.A2(n_856),
.B(n_866),
.Y(n_1097)
);

NOR2x1_ASAP7_75t_SL g1098 ( 
.A(n_910),
.B(n_636),
.Y(n_1098)
);

NAND2xp5_ASAP7_75t_L g1099 ( 
.A(n_926),
.B(n_935),
.Y(n_1099)
);

AOI21xp5_ASAP7_75t_L g1100 ( 
.A1(n_926),
.A2(n_939),
.B(n_935),
.Y(n_1100)
);

INVx1_ASAP7_75t_L g1101 ( 
.A(n_781),
.Y(n_1101)
);

AOI21x1_ASAP7_75t_L g1102 ( 
.A1(n_900),
.A2(n_866),
.B(n_951),
.Y(n_1102)
);

AND2x2_ASAP7_75t_L g1103 ( 
.A(n_876),
.B(n_620),
.Y(n_1103)
);

AOI21xp5_ASAP7_75t_L g1104 ( 
.A1(n_926),
.A2(n_939),
.B(n_935),
.Y(n_1104)
);

INVx1_ASAP7_75t_L g1105 ( 
.A(n_781),
.Y(n_1105)
);

OAI21xp5_ASAP7_75t_L g1106 ( 
.A1(n_926),
.A2(n_959),
.B(n_935),
.Y(n_1106)
);

AOI21x1_ASAP7_75t_L g1107 ( 
.A1(n_900),
.A2(n_866),
.B(n_951),
.Y(n_1107)
);

O2A1O1Ixp5_ASAP7_75t_L g1108 ( 
.A1(n_926),
.A2(n_939),
.B(n_942),
.C(n_941),
.Y(n_1108)
);

NAND2xp5_ASAP7_75t_L g1109 ( 
.A(n_926),
.B(n_935),
.Y(n_1109)
);

OAI21xp5_ASAP7_75t_L g1110 ( 
.A1(n_926),
.A2(n_959),
.B(n_935),
.Y(n_1110)
);

AO21x2_ASAP7_75t_L g1111 ( 
.A1(n_807),
.A2(n_925),
.B(n_832),
.Y(n_1111)
);

OAI21x1_ASAP7_75t_L g1112 ( 
.A1(n_961),
.A2(n_856),
.B(n_866),
.Y(n_1112)
);

AOI22xp33_ASAP7_75t_L g1113 ( 
.A1(n_1073),
.A2(n_1093),
.B1(n_988),
.B2(n_1096),
.Y(n_1113)
);

INVx1_ASAP7_75t_L g1114 ( 
.A(n_967),
.Y(n_1114)
);

INVx1_ASAP7_75t_L g1115 ( 
.A(n_968),
.Y(n_1115)
);

HB1xp67_ASAP7_75t_L g1116 ( 
.A(n_974),
.Y(n_1116)
);

INVx3_ASAP7_75t_L g1117 ( 
.A(n_980),
.Y(n_1117)
);

OAI33xp33_ASAP7_75t_L g1118 ( 
.A1(n_1011),
.A2(n_970),
.A3(n_1010),
.B1(n_969),
.B2(n_971),
.B3(n_1071),
.Y(n_1118)
);

AND2x2_ASAP7_75t_L g1119 ( 
.A(n_1103),
.B(n_1019),
.Y(n_1119)
);

O2A1O1Ixp33_ASAP7_75t_L g1120 ( 
.A1(n_1080),
.A2(n_977),
.B(n_1069),
.C(n_1096),
.Y(n_1120)
);

OAI321xp33_ASAP7_75t_L g1121 ( 
.A1(n_991),
.A2(n_977),
.A3(n_979),
.B1(n_972),
.B2(n_994),
.C(n_1003),
.Y(n_1121)
);

INVx1_ASAP7_75t_SL g1122 ( 
.A(n_990),
.Y(n_1122)
);

NAND2xp5_ASAP7_75t_L g1123 ( 
.A(n_1062),
.B(n_1065),
.Y(n_1123)
);

NAND2xp5_ASAP7_75t_L g1124 ( 
.A(n_1067),
.B(n_1084),
.Y(n_1124)
);

INVx1_ASAP7_75t_SL g1125 ( 
.A(n_1077),
.Y(n_1125)
);

AND2x4_ASAP7_75t_L g1126 ( 
.A(n_1066),
.B(n_1089),
.Y(n_1126)
);

AOI22xp5_ASAP7_75t_L g1127 ( 
.A1(n_991),
.A2(n_1099),
.B1(n_1088),
.B2(n_1109),
.Y(n_1127)
);

INVx3_ASAP7_75t_L g1128 ( 
.A(n_980),
.Y(n_1128)
);

OAI21xp5_ASAP7_75t_L g1129 ( 
.A1(n_1061),
.A2(n_1100),
.B(n_1104),
.Y(n_1129)
);

NAND3xp33_ASAP7_75t_L g1130 ( 
.A(n_1080),
.B(n_1069),
.C(n_1003),
.Y(n_1130)
);

AND2x2_ASAP7_75t_L g1131 ( 
.A(n_1083),
.B(n_1007),
.Y(n_1131)
);

NAND2xp5_ASAP7_75t_L g1132 ( 
.A(n_1090),
.B(n_1092),
.Y(n_1132)
);

AOI21xp5_ASAP7_75t_SL g1133 ( 
.A1(n_1015),
.A2(n_976),
.B(n_995),
.Y(n_1133)
);

NAND2xp5_ASAP7_75t_L g1134 ( 
.A(n_1106),
.B(n_1110),
.Y(n_1134)
);

OA21x2_ASAP7_75t_L g1135 ( 
.A1(n_978),
.A2(n_1017),
.B(n_1112),
.Y(n_1135)
);

AOI22xp33_ASAP7_75t_L g1136 ( 
.A1(n_1075),
.A2(n_1095),
.B1(n_1024),
.B2(n_1057),
.Y(n_1136)
);

INVx3_ASAP7_75t_L g1137 ( 
.A(n_980),
.Y(n_1137)
);

INVx1_ASAP7_75t_L g1138 ( 
.A(n_1074),
.Y(n_1138)
);

AND2x4_ASAP7_75t_L g1139 ( 
.A(n_1089),
.B(n_1098),
.Y(n_1139)
);

INVx1_ASAP7_75t_L g1140 ( 
.A(n_1091),
.Y(n_1140)
);

INVxp67_ASAP7_75t_L g1141 ( 
.A(n_982),
.Y(n_1141)
);

OAI22xp5_ASAP7_75t_L g1142 ( 
.A1(n_1004),
.A2(n_1028),
.B1(n_995),
.B2(n_1015),
.Y(n_1142)
);

A2O1A1Ixp33_ASAP7_75t_L g1143 ( 
.A1(n_1108),
.A2(n_1004),
.B(n_1034),
.C(n_1032),
.Y(n_1143)
);

NOR2xp33_ASAP7_75t_R g1144 ( 
.A(n_1013),
.B(n_1018),
.Y(n_1144)
);

O2A1O1Ixp33_ASAP7_75t_L g1145 ( 
.A1(n_981),
.A2(n_1108),
.B(n_985),
.C(n_1029),
.Y(n_1145)
);

INVx3_ASAP7_75t_L g1146 ( 
.A(n_1006),
.Y(n_1146)
);

NAND2xp5_ASAP7_75t_L g1147 ( 
.A(n_999),
.B(n_1027),
.Y(n_1147)
);

INVx1_ASAP7_75t_L g1148 ( 
.A(n_1101),
.Y(n_1148)
);

NAND2xp5_ASAP7_75t_L g1149 ( 
.A(n_1030),
.B(n_1105),
.Y(n_1149)
);

OR2x6_ASAP7_75t_L g1150 ( 
.A(n_986),
.B(n_1035),
.Y(n_1150)
);

NOR2x1_ASAP7_75t_L g1151 ( 
.A(n_1014),
.B(n_975),
.Y(n_1151)
);

NOR2xp67_ASAP7_75t_L g1152 ( 
.A(n_1039),
.B(n_1052),
.Y(n_1152)
);

OAI22xp33_ASAP7_75t_L g1153 ( 
.A1(n_993),
.A2(n_1082),
.B1(n_1014),
.B2(n_1043),
.Y(n_1153)
);

INVx1_ASAP7_75t_L g1154 ( 
.A(n_1041),
.Y(n_1154)
);

AND2x4_ASAP7_75t_L g1155 ( 
.A(n_1039),
.B(n_1002),
.Y(n_1155)
);

AOI21xp5_ASAP7_75t_L g1156 ( 
.A1(n_981),
.A2(n_1009),
.B(n_1033),
.Y(n_1156)
);

AND2x2_ASAP7_75t_L g1157 ( 
.A(n_1045),
.B(n_1026),
.Y(n_1157)
);

INVx3_ASAP7_75t_L g1158 ( 
.A(n_1006),
.Y(n_1158)
);

NAND2xp5_ASAP7_75t_L g1159 ( 
.A(n_1064),
.B(n_1002),
.Y(n_1159)
);

INVx2_ASAP7_75t_SL g1160 ( 
.A(n_1078),
.Y(n_1160)
);

AOI21xp5_ASAP7_75t_L g1161 ( 
.A1(n_1016),
.A2(n_992),
.B(n_1020),
.Y(n_1161)
);

AND2x4_ASAP7_75t_L g1162 ( 
.A(n_1063),
.B(n_1085),
.Y(n_1162)
);

BUFx4f_ASAP7_75t_SL g1163 ( 
.A(n_1026),
.Y(n_1163)
);

INVx1_ASAP7_75t_L g1164 ( 
.A(n_1031),
.Y(n_1164)
);

BUFx12f_ASAP7_75t_L g1165 ( 
.A(n_1026),
.Y(n_1165)
);

BUFx6f_ASAP7_75t_L g1166 ( 
.A(n_1008),
.Y(n_1166)
);

AND2x2_ASAP7_75t_L g1167 ( 
.A(n_1056),
.B(n_1037),
.Y(n_1167)
);

HB1xp67_ASAP7_75t_L g1168 ( 
.A(n_1008),
.Y(n_1168)
);

INVx1_ASAP7_75t_L g1169 ( 
.A(n_1049),
.Y(n_1169)
);

CKINVDCx5p33_ASAP7_75t_R g1170 ( 
.A(n_1008),
.Y(n_1170)
);

OAI21xp33_ASAP7_75t_SL g1171 ( 
.A1(n_1000),
.A2(n_998),
.B(n_1036),
.Y(n_1171)
);

OAI21x1_ASAP7_75t_SL g1172 ( 
.A1(n_983),
.A2(n_1053),
.B(n_996),
.Y(n_1172)
);

CKINVDCx5p33_ASAP7_75t_R g1173 ( 
.A(n_1047),
.Y(n_1173)
);

AO21x1_ASAP7_75t_L g1174 ( 
.A1(n_1021),
.A2(n_1023),
.B(n_1000),
.Y(n_1174)
);

AOI21xp5_ASAP7_75t_L g1175 ( 
.A1(n_1021),
.A2(n_1012),
.B(n_1060),
.Y(n_1175)
);

NAND2xp5_ASAP7_75t_L g1176 ( 
.A(n_1087),
.B(n_1042),
.Y(n_1176)
);

AOI21xp5_ASAP7_75t_L g1177 ( 
.A1(n_1060),
.A2(n_1086),
.B(n_1079),
.Y(n_1177)
);

AND2x4_ASAP7_75t_L g1178 ( 
.A(n_1087),
.B(n_1055),
.Y(n_1178)
);

AND2x4_ASAP7_75t_L g1179 ( 
.A(n_1048),
.B(n_1081),
.Y(n_1179)
);

BUFx6f_ASAP7_75t_L g1180 ( 
.A(n_973),
.Y(n_1180)
);

INVx1_ASAP7_75t_L g1181 ( 
.A(n_1081),
.Y(n_1181)
);

O2A1O1Ixp33_ASAP7_75t_L g1182 ( 
.A1(n_1056),
.A2(n_1054),
.B(n_1086),
.C(n_1060),
.Y(n_1182)
);

INVx1_ASAP7_75t_L g1183 ( 
.A(n_1022),
.Y(n_1183)
);

AOI221xp5_ASAP7_75t_L g1184 ( 
.A1(n_1044),
.A2(n_1046),
.B1(n_1111),
.B2(n_987),
.C(n_1038),
.Y(n_1184)
);

NAND2x1p5_ASAP7_75t_L g1185 ( 
.A(n_1050),
.B(n_1025),
.Y(n_1185)
);

INVx5_ASAP7_75t_L g1186 ( 
.A(n_1040),
.Y(n_1186)
);

AND2x2_ASAP7_75t_L g1187 ( 
.A(n_987),
.B(n_1051),
.Y(n_1187)
);

INVx1_ASAP7_75t_L g1188 ( 
.A(n_1022),
.Y(n_1188)
);

OAI22xp5_ASAP7_75t_L g1189 ( 
.A1(n_1086),
.A2(n_989),
.B1(n_1076),
.B2(n_1102),
.Y(n_1189)
);

INVx1_ASAP7_75t_L g1190 ( 
.A(n_1022),
.Y(n_1190)
);

AND2x4_ASAP7_75t_L g1191 ( 
.A(n_987),
.B(n_1038),
.Y(n_1191)
);

NAND2xp5_ASAP7_75t_L g1192 ( 
.A(n_987),
.B(n_984),
.Y(n_1192)
);

NOR2xp33_ASAP7_75t_L g1193 ( 
.A(n_1107),
.B(n_997),
.Y(n_1193)
);

NAND2xp5_ASAP7_75t_L g1194 ( 
.A(n_984),
.B(n_1022),
.Y(n_1194)
);

NAND3xp33_ASAP7_75t_L g1195 ( 
.A(n_1040),
.B(n_984),
.C(n_1005),
.Y(n_1195)
);

NAND2xp5_ASAP7_75t_SL g1196 ( 
.A(n_1001),
.B(n_1017),
.Y(n_1196)
);

INVx3_ASAP7_75t_SL g1197 ( 
.A(n_1005),
.Y(n_1197)
);

AOI21xp5_ASAP7_75t_L g1198 ( 
.A1(n_1070),
.A2(n_1072),
.B(n_1068),
.Y(n_1198)
);

NAND2xp5_ASAP7_75t_L g1199 ( 
.A(n_1005),
.B(n_978),
.Y(n_1199)
);

BUFx12f_ASAP7_75t_L g1200 ( 
.A(n_966),
.Y(n_1200)
);

INVx1_ASAP7_75t_L g1201 ( 
.A(n_966),
.Y(n_1201)
);

AOI22xp5_ASAP7_75t_L g1202 ( 
.A1(n_1058),
.A2(n_1059),
.B1(n_1068),
.B2(n_1094),
.Y(n_1202)
);

AND2x2_ASAP7_75t_L g1203 ( 
.A(n_1058),
.B(n_1059),
.Y(n_1203)
);

OAI22xp5_ASAP7_75t_SL g1204 ( 
.A1(n_1094),
.A2(n_938),
.B1(n_1011),
.B2(n_935),
.Y(n_1204)
);

NOR2xp33_ASAP7_75t_L g1205 ( 
.A(n_1097),
.B(n_1112),
.Y(n_1205)
);

AOI21xp5_ASAP7_75t_SL g1206 ( 
.A1(n_1097),
.A2(n_835),
.B(n_926),
.Y(n_1206)
);

CKINVDCx5p33_ASAP7_75t_R g1207 ( 
.A(n_975),
.Y(n_1207)
);

INVx1_ASAP7_75t_L g1208 ( 
.A(n_967),
.Y(n_1208)
);

OR2x6_ASAP7_75t_L g1209 ( 
.A(n_986),
.B(n_634),
.Y(n_1209)
);

AOI22xp5_ASAP7_75t_L g1210 ( 
.A1(n_1096),
.A2(n_935),
.B1(n_939),
.B2(n_926),
.Y(n_1210)
);

CKINVDCx5p33_ASAP7_75t_R g1211 ( 
.A(n_975),
.Y(n_1211)
);

CKINVDCx11_ASAP7_75t_R g1212 ( 
.A(n_1014),
.Y(n_1212)
);

NOR2xp67_ASAP7_75t_SL g1213 ( 
.A(n_975),
.B(n_599),
.Y(n_1213)
);

OAI22xp5_ASAP7_75t_L g1214 ( 
.A1(n_988),
.A2(n_926),
.B1(n_939),
.B2(n_935),
.Y(n_1214)
);

BUFx2_ASAP7_75t_L g1215 ( 
.A(n_974),
.Y(n_1215)
);

NOR2xp33_ASAP7_75t_SL g1216 ( 
.A(n_988),
.B(n_877),
.Y(n_1216)
);

INVx5_ASAP7_75t_L g1217 ( 
.A(n_980),
.Y(n_1217)
);

AOI211xp5_ASAP7_75t_L g1218 ( 
.A1(n_1011),
.A2(n_958),
.B(n_935),
.C(n_941),
.Y(n_1218)
);

AOI21xp5_ASAP7_75t_L g1219 ( 
.A1(n_977),
.A2(n_935),
.B(n_926),
.Y(n_1219)
);

INVx2_ASAP7_75t_SL g1220 ( 
.A(n_1013),
.Y(n_1220)
);

NAND2xp5_ASAP7_75t_L g1221 ( 
.A(n_1096),
.B(n_969),
.Y(n_1221)
);

OAI22xp5_ASAP7_75t_L g1222 ( 
.A1(n_1096),
.A2(n_926),
.B1(n_939),
.B2(n_935),
.Y(n_1222)
);

AOI21xp5_ASAP7_75t_L g1223 ( 
.A1(n_977),
.A2(n_935),
.B(n_926),
.Y(n_1223)
);

BUFx3_ASAP7_75t_L g1224 ( 
.A(n_1013),
.Y(n_1224)
);

NAND2xp5_ASAP7_75t_L g1225 ( 
.A(n_1096),
.B(n_969),
.Y(n_1225)
);

AND2x4_ASAP7_75t_L g1226 ( 
.A(n_1066),
.B(n_1089),
.Y(n_1226)
);

OR2x2_ASAP7_75t_L g1227 ( 
.A(n_1007),
.B(n_715),
.Y(n_1227)
);

AOI22xp5_ASAP7_75t_L g1228 ( 
.A1(n_1096),
.A2(n_935),
.B1(n_939),
.B2(n_926),
.Y(n_1228)
);

AND2x2_ASAP7_75t_L g1229 ( 
.A(n_1103),
.B(n_876),
.Y(n_1229)
);

INVx1_ASAP7_75t_SL g1230 ( 
.A(n_990),
.Y(n_1230)
);

BUFx2_ASAP7_75t_L g1231 ( 
.A(n_974),
.Y(n_1231)
);

INVx3_ASAP7_75t_L g1232 ( 
.A(n_980),
.Y(n_1232)
);

O2A1O1Ixp5_ASAP7_75t_SL g1233 ( 
.A1(n_991),
.A2(n_977),
.B(n_988),
.C(n_979),
.Y(n_1233)
);

O2A1O1Ixp5_ASAP7_75t_SL g1234 ( 
.A1(n_991),
.A2(n_977),
.B(n_988),
.C(n_979),
.Y(n_1234)
);

INVx1_ASAP7_75t_L g1235 ( 
.A(n_967),
.Y(n_1235)
);

OR2x6_ASAP7_75t_L g1236 ( 
.A(n_986),
.B(n_634),
.Y(n_1236)
);

INVx5_ASAP7_75t_L g1237 ( 
.A(n_980),
.Y(n_1237)
);

INVx1_ASAP7_75t_L g1238 ( 
.A(n_967),
.Y(n_1238)
);

INVx1_ASAP7_75t_L g1239 ( 
.A(n_967),
.Y(n_1239)
);

AND2x2_ASAP7_75t_L g1240 ( 
.A(n_1103),
.B(n_876),
.Y(n_1240)
);

NAND2xp5_ASAP7_75t_L g1241 ( 
.A(n_1096),
.B(n_969),
.Y(n_1241)
);

NAND3xp33_ASAP7_75t_L g1242 ( 
.A(n_972),
.B(n_938),
.C(n_935),
.Y(n_1242)
);

CKINVDCx5p33_ASAP7_75t_R g1243 ( 
.A(n_975),
.Y(n_1243)
);

AOI21xp33_ASAP7_75t_SL g1244 ( 
.A1(n_1222),
.A2(n_1225),
.B(n_1221),
.Y(n_1244)
);

AOI22xp33_ASAP7_75t_L g1245 ( 
.A1(n_1216),
.A2(n_1214),
.B1(n_1113),
.B2(n_1130),
.Y(n_1245)
);

OAI21x1_ASAP7_75t_L g1246 ( 
.A1(n_1198),
.A2(n_1161),
.B(n_1177),
.Y(n_1246)
);

INVx1_ASAP7_75t_L g1247 ( 
.A(n_1114),
.Y(n_1247)
);

OA21x2_ASAP7_75t_L g1248 ( 
.A1(n_1156),
.A2(n_1175),
.B(n_1129),
.Y(n_1248)
);

INVx3_ASAP7_75t_L g1249 ( 
.A(n_1200),
.Y(n_1249)
);

AND2x4_ASAP7_75t_L g1250 ( 
.A(n_1139),
.B(n_1126),
.Y(n_1250)
);

OAI21x1_ASAP7_75t_L g1251 ( 
.A1(n_1189),
.A2(n_1196),
.B(n_1199),
.Y(n_1251)
);

INVx1_ASAP7_75t_L g1252 ( 
.A(n_1115),
.Y(n_1252)
);

HB1xp67_ASAP7_75t_L g1253 ( 
.A(n_1116),
.Y(n_1253)
);

OR2x6_ASAP7_75t_L g1254 ( 
.A(n_1182),
.B(n_1133),
.Y(n_1254)
);

INVx1_ASAP7_75t_SL g1255 ( 
.A(n_1144),
.Y(n_1255)
);

BUFx2_ASAP7_75t_R g1256 ( 
.A(n_1173),
.Y(n_1256)
);

OAI22xp33_ASAP7_75t_L g1257 ( 
.A1(n_1210),
.A2(n_1228),
.B1(n_1216),
.B2(n_1241),
.Y(n_1257)
);

INVx1_ASAP7_75t_L g1258 ( 
.A(n_1138),
.Y(n_1258)
);

NAND2xp33_ASAP7_75t_SL g1259 ( 
.A(n_1204),
.B(n_1134),
.Y(n_1259)
);

OAI22xp5_ASAP7_75t_L g1260 ( 
.A1(n_1210),
.A2(n_1218),
.B1(n_1242),
.B2(n_1136),
.Y(n_1260)
);

OR2x2_ASAP7_75t_L g1261 ( 
.A(n_1192),
.B(n_1194),
.Y(n_1261)
);

AOI22xp33_ASAP7_75t_L g1262 ( 
.A1(n_1229),
.A2(n_1240),
.B1(n_1204),
.B2(n_1119),
.Y(n_1262)
);

INVx1_ASAP7_75t_L g1263 ( 
.A(n_1140),
.Y(n_1263)
);

INVx1_ASAP7_75t_L g1264 ( 
.A(n_1148),
.Y(n_1264)
);

AOI22xp33_ASAP7_75t_L g1265 ( 
.A1(n_1118),
.A2(n_1153),
.B1(n_1179),
.B2(n_1142),
.Y(n_1265)
);

AO21x1_ASAP7_75t_SL g1266 ( 
.A1(n_1129),
.A2(n_1190),
.B(n_1188),
.Y(n_1266)
);

INVx3_ASAP7_75t_L g1267 ( 
.A(n_1186),
.Y(n_1267)
);

INVx1_ASAP7_75t_L g1268 ( 
.A(n_1208),
.Y(n_1268)
);

INVx1_ASAP7_75t_L g1269 ( 
.A(n_1235),
.Y(n_1269)
);

NAND2xp5_ASAP7_75t_L g1270 ( 
.A(n_1123),
.B(n_1124),
.Y(n_1270)
);

HB1xp67_ASAP7_75t_L g1271 ( 
.A(n_1125),
.Y(n_1271)
);

CKINVDCx20_ASAP7_75t_R g1272 ( 
.A(n_1212),
.Y(n_1272)
);

AOI222xp33_ASAP7_75t_L g1273 ( 
.A1(n_1121),
.A2(n_1132),
.B1(n_1147),
.B2(n_1131),
.C1(n_1238),
.C2(n_1239),
.Y(n_1273)
);

HB1xp67_ASAP7_75t_L g1274 ( 
.A(n_1125),
.Y(n_1274)
);

AO21x1_ASAP7_75t_L g1275 ( 
.A1(n_1218),
.A2(n_1120),
.B(n_1223),
.Y(n_1275)
);

INVx1_ASAP7_75t_SL g1276 ( 
.A(n_1122),
.Y(n_1276)
);

INVx1_ASAP7_75t_L g1277 ( 
.A(n_1154),
.Y(n_1277)
);

AOI22xp33_ASAP7_75t_L g1278 ( 
.A1(n_1179),
.A2(n_1219),
.B1(n_1230),
.B2(n_1122),
.Y(n_1278)
);

AND2x2_ASAP7_75t_L g1279 ( 
.A(n_1233),
.B(n_1234),
.Y(n_1279)
);

BUFx2_ASAP7_75t_L g1280 ( 
.A(n_1191),
.Y(n_1280)
);

HB1xp67_ASAP7_75t_L g1281 ( 
.A(n_1215),
.Y(n_1281)
);

INVxp67_ASAP7_75t_L g1282 ( 
.A(n_1231),
.Y(n_1282)
);

AND2x2_ASAP7_75t_L g1283 ( 
.A(n_1127),
.B(n_1187),
.Y(n_1283)
);

AOI22xp33_ASAP7_75t_L g1284 ( 
.A1(n_1230),
.A2(n_1127),
.B1(n_1181),
.B2(n_1169),
.Y(n_1284)
);

INVx1_ASAP7_75t_L g1285 ( 
.A(n_1164),
.Y(n_1285)
);

BUFx2_ASAP7_75t_L g1286 ( 
.A(n_1185),
.Y(n_1286)
);

CKINVDCx6p67_ASAP7_75t_R g1287 ( 
.A(n_1150),
.Y(n_1287)
);

INVx1_ASAP7_75t_L g1288 ( 
.A(n_1149),
.Y(n_1288)
);

NAND2xp5_ASAP7_75t_L g1289 ( 
.A(n_1227),
.B(n_1126),
.Y(n_1289)
);

OAI22xp5_ASAP7_75t_SL g1290 ( 
.A1(n_1150),
.A2(n_1243),
.B1(n_1207),
.B2(n_1211),
.Y(n_1290)
);

OR2x2_ASAP7_75t_L g1291 ( 
.A(n_1195),
.B(n_1197),
.Y(n_1291)
);

AOI22xp33_ASAP7_75t_L g1292 ( 
.A1(n_1167),
.A2(n_1184),
.B1(n_1157),
.B2(n_1141),
.Y(n_1292)
);

AOI22xp33_ASAP7_75t_L g1293 ( 
.A1(n_1150),
.A2(n_1160),
.B1(n_1213),
.B2(n_1165),
.Y(n_1293)
);

AOI222xp33_ASAP7_75t_L g1294 ( 
.A1(n_1121),
.A2(n_1143),
.B1(n_1171),
.B2(n_1163),
.C1(n_1195),
.C2(n_1176),
.Y(n_1294)
);

AOI22xp33_ASAP7_75t_L g1295 ( 
.A1(n_1178),
.A2(n_1186),
.B1(n_1236),
.B2(n_1209),
.Y(n_1295)
);

BUFx3_ASAP7_75t_L g1296 ( 
.A(n_1224),
.Y(n_1296)
);

OAI22xp5_ASAP7_75t_L g1297 ( 
.A1(n_1220),
.A2(n_1206),
.B1(n_1226),
.B2(n_1151),
.Y(n_1297)
);

AOI22xp33_ASAP7_75t_L g1298 ( 
.A1(n_1186),
.A2(n_1209),
.B1(n_1236),
.B2(n_1172),
.Y(n_1298)
);

INVx11_ASAP7_75t_L g1299 ( 
.A(n_1170),
.Y(n_1299)
);

INVx1_ASAP7_75t_L g1300 ( 
.A(n_1168),
.Y(n_1300)
);

INVx1_ASAP7_75t_L g1301 ( 
.A(n_1159),
.Y(n_1301)
);

OR2x2_ASAP7_75t_L g1302 ( 
.A(n_1174),
.B(n_1201),
.Y(n_1302)
);

INVx2_ASAP7_75t_L g1303 ( 
.A(n_1135),
.Y(n_1303)
);

BUFx2_ASAP7_75t_L g1304 ( 
.A(n_1171),
.Y(n_1304)
);

INVx2_ASAP7_75t_L g1305 ( 
.A(n_1135),
.Y(n_1305)
);

OAI21x1_ASAP7_75t_L g1306 ( 
.A1(n_1202),
.A2(n_1145),
.B(n_1203),
.Y(n_1306)
);

INVx1_ASAP7_75t_L g1307 ( 
.A(n_1166),
.Y(n_1307)
);

INVx1_ASAP7_75t_L g1308 ( 
.A(n_1117),
.Y(n_1308)
);

INVx2_ASAP7_75t_L g1309 ( 
.A(n_1193),
.Y(n_1309)
);

BUFx2_ASAP7_75t_L g1310 ( 
.A(n_1205),
.Y(n_1310)
);

BUFx2_ASAP7_75t_L g1311 ( 
.A(n_1128),
.Y(n_1311)
);

INVx2_ASAP7_75t_L g1312 ( 
.A(n_1137),
.Y(n_1312)
);

INVx1_ASAP7_75t_L g1313 ( 
.A(n_1137),
.Y(n_1313)
);

AOI21x1_ASAP7_75t_L g1314 ( 
.A1(n_1152),
.A2(n_1162),
.B(n_1155),
.Y(n_1314)
);

INVx1_ASAP7_75t_L g1315 ( 
.A(n_1146),
.Y(n_1315)
);

INVx3_ASAP7_75t_L g1316 ( 
.A(n_1158),
.Y(n_1316)
);

AND2x2_ASAP7_75t_L g1317 ( 
.A(n_1232),
.B(n_1217),
.Y(n_1317)
);

HB1xp67_ASAP7_75t_L g1318 ( 
.A(n_1217),
.Y(n_1318)
);

INVx1_ASAP7_75t_L g1319 ( 
.A(n_1237),
.Y(n_1319)
);

INVx1_ASAP7_75t_L g1320 ( 
.A(n_1152),
.Y(n_1320)
);

NAND2xp5_ASAP7_75t_L g1321 ( 
.A(n_1180),
.B(n_1221),
.Y(n_1321)
);

OAI21xp5_ASAP7_75t_L g1322 ( 
.A1(n_1216),
.A2(n_938),
.B(n_935),
.Y(n_1322)
);

AOI22xp33_ASAP7_75t_L g1323 ( 
.A1(n_1216),
.A2(n_877),
.B1(n_881),
.B2(n_752),
.Y(n_1323)
);

OAI22xp33_ASAP7_75t_L g1324 ( 
.A1(n_1210),
.A2(n_938),
.B1(n_926),
.B2(n_935),
.Y(n_1324)
);

BUFx8_ASAP7_75t_L g1325 ( 
.A(n_1215),
.Y(n_1325)
);

CKINVDCx20_ASAP7_75t_R g1326 ( 
.A(n_1212),
.Y(n_1326)
);

HB1xp67_ASAP7_75t_L g1327 ( 
.A(n_1116),
.Y(n_1327)
);

CKINVDCx6p67_ASAP7_75t_R g1328 ( 
.A(n_1212),
.Y(n_1328)
);

INVx1_ASAP7_75t_L g1329 ( 
.A(n_1114),
.Y(n_1329)
);

INVx1_ASAP7_75t_L g1330 ( 
.A(n_1114),
.Y(n_1330)
);

BUFx2_ASAP7_75t_L g1331 ( 
.A(n_1200),
.Y(n_1331)
);

INVx1_ASAP7_75t_L g1332 ( 
.A(n_1183),
.Y(n_1332)
);

OAI21xp5_ASAP7_75t_L g1333 ( 
.A1(n_1216),
.A2(n_938),
.B(n_935),
.Y(n_1333)
);

CKINVDCx14_ASAP7_75t_R g1334 ( 
.A(n_1144),
.Y(n_1334)
);

AND2x4_ASAP7_75t_L g1335 ( 
.A(n_1139),
.B(n_1126),
.Y(n_1335)
);

INVx3_ASAP7_75t_L g1336 ( 
.A(n_1200),
.Y(n_1336)
);

INVx1_ASAP7_75t_L g1337 ( 
.A(n_1114),
.Y(n_1337)
);

INVx1_ASAP7_75t_L g1338 ( 
.A(n_1114),
.Y(n_1338)
);

INVx3_ASAP7_75t_L g1339 ( 
.A(n_1200),
.Y(n_1339)
);

INVx1_ASAP7_75t_SL g1340 ( 
.A(n_1144),
.Y(n_1340)
);

AOI22xp33_ASAP7_75t_L g1341 ( 
.A1(n_1216),
.A2(n_877),
.B1(n_881),
.B2(n_752),
.Y(n_1341)
);

OR2x2_ASAP7_75t_L g1342 ( 
.A(n_1192),
.B(n_1113),
.Y(n_1342)
);

AO21x2_ASAP7_75t_L g1343 ( 
.A1(n_1303),
.A2(n_1305),
.B(n_1309),
.Y(n_1343)
);

OA21x2_ASAP7_75t_L g1344 ( 
.A1(n_1246),
.A2(n_1306),
.B(n_1251),
.Y(n_1344)
);

INVx1_ASAP7_75t_L g1345 ( 
.A(n_1332),
.Y(n_1345)
);

BUFx6f_ASAP7_75t_L g1346 ( 
.A(n_1266),
.Y(n_1346)
);

OR2x2_ASAP7_75t_L g1347 ( 
.A(n_1261),
.B(n_1283),
.Y(n_1347)
);

INVx2_ASAP7_75t_L g1348 ( 
.A(n_1302),
.Y(n_1348)
);

NAND2xp5_ASAP7_75t_L g1349 ( 
.A(n_1270),
.B(n_1244),
.Y(n_1349)
);

INVx1_ASAP7_75t_L g1350 ( 
.A(n_1261),
.Y(n_1350)
);

OR2x2_ASAP7_75t_L g1351 ( 
.A(n_1283),
.B(n_1304),
.Y(n_1351)
);

INVx2_ASAP7_75t_L g1352 ( 
.A(n_1302),
.Y(n_1352)
);

AND2x2_ASAP7_75t_L g1353 ( 
.A(n_1304),
.B(n_1310),
.Y(n_1353)
);

INVx1_ASAP7_75t_L g1354 ( 
.A(n_1285),
.Y(n_1354)
);

HB1xp67_ASAP7_75t_L g1355 ( 
.A(n_1271),
.Y(n_1355)
);

NOR2xp33_ASAP7_75t_L g1356 ( 
.A(n_1256),
.B(n_1296),
.Y(n_1356)
);

INVx1_ASAP7_75t_SL g1357 ( 
.A(n_1255),
.Y(n_1357)
);

INVx1_ASAP7_75t_L g1358 ( 
.A(n_1247),
.Y(n_1358)
);

NAND2xp5_ASAP7_75t_L g1359 ( 
.A(n_1257),
.B(n_1288),
.Y(n_1359)
);

HB1xp67_ASAP7_75t_L g1360 ( 
.A(n_1274),
.Y(n_1360)
);

INVx1_ASAP7_75t_L g1361 ( 
.A(n_1252),
.Y(n_1361)
);

INVx2_ASAP7_75t_SL g1362 ( 
.A(n_1249),
.Y(n_1362)
);

HB1xp67_ASAP7_75t_L g1363 ( 
.A(n_1253),
.Y(n_1363)
);

AND2x2_ASAP7_75t_L g1364 ( 
.A(n_1310),
.B(n_1280),
.Y(n_1364)
);

OR2x2_ASAP7_75t_L g1365 ( 
.A(n_1342),
.B(n_1291),
.Y(n_1365)
);

AND2x2_ASAP7_75t_L g1366 ( 
.A(n_1280),
.B(n_1258),
.Y(n_1366)
);

INVx1_ASAP7_75t_L g1367 ( 
.A(n_1263),
.Y(n_1367)
);

NAND2xp5_ASAP7_75t_L g1368 ( 
.A(n_1273),
.B(n_1276),
.Y(n_1368)
);

INVx1_ASAP7_75t_L g1369 ( 
.A(n_1264),
.Y(n_1369)
);

NAND2xp5_ASAP7_75t_L g1370 ( 
.A(n_1327),
.B(n_1321),
.Y(n_1370)
);

INVx3_ASAP7_75t_L g1371 ( 
.A(n_1248),
.Y(n_1371)
);

INVx1_ASAP7_75t_L g1372 ( 
.A(n_1268),
.Y(n_1372)
);

INVx1_ASAP7_75t_L g1373 ( 
.A(n_1269),
.Y(n_1373)
);

NOR2xp33_ASAP7_75t_L g1374 ( 
.A(n_1296),
.B(n_1340),
.Y(n_1374)
);

INVx1_ASAP7_75t_L g1375 ( 
.A(n_1277),
.Y(n_1375)
);

OR2x2_ASAP7_75t_L g1376 ( 
.A(n_1342),
.B(n_1291),
.Y(n_1376)
);

HB1xp67_ASAP7_75t_L g1377 ( 
.A(n_1300),
.Y(n_1377)
);

AND2x2_ASAP7_75t_L g1378 ( 
.A(n_1329),
.B(n_1330),
.Y(n_1378)
);

INVx1_ASAP7_75t_L g1379 ( 
.A(n_1337),
.Y(n_1379)
);

INVx1_ASAP7_75t_L g1380 ( 
.A(n_1338),
.Y(n_1380)
);

INVx1_ASAP7_75t_L g1381 ( 
.A(n_1320),
.Y(n_1381)
);

INVx4_ASAP7_75t_SL g1382 ( 
.A(n_1254),
.Y(n_1382)
);

INVxp67_ASAP7_75t_L g1383 ( 
.A(n_1281),
.Y(n_1383)
);

OR2x2_ASAP7_75t_L g1384 ( 
.A(n_1260),
.B(n_1245),
.Y(n_1384)
);

OR2x6_ASAP7_75t_L g1385 ( 
.A(n_1254),
.B(n_1331),
.Y(n_1385)
);

INVx1_ASAP7_75t_L g1386 ( 
.A(n_1320),
.Y(n_1386)
);

INVx1_ASAP7_75t_SL g1387 ( 
.A(n_1290),
.Y(n_1387)
);

BUFx6f_ASAP7_75t_L g1388 ( 
.A(n_1266),
.Y(n_1388)
);

INVx3_ASAP7_75t_L g1389 ( 
.A(n_1248),
.Y(n_1389)
);

INVx3_ASAP7_75t_L g1390 ( 
.A(n_1248),
.Y(n_1390)
);

NOR2xp67_ASAP7_75t_R g1391 ( 
.A(n_1259),
.B(n_1267),
.Y(n_1391)
);

OAI21x1_ASAP7_75t_L g1392 ( 
.A1(n_1314),
.A2(n_1275),
.B(n_1298),
.Y(n_1392)
);

BUFx3_ASAP7_75t_L g1393 ( 
.A(n_1249),
.Y(n_1393)
);

OR2x6_ASAP7_75t_L g1394 ( 
.A(n_1254),
.B(n_1331),
.Y(n_1394)
);

AND2x2_ASAP7_75t_L g1395 ( 
.A(n_1286),
.B(n_1262),
.Y(n_1395)
);

INVx1_ASAP7_75t_L g1396 ( 
.A(n_1286),
.Y(n_1396)
);

NAND2xp5_ASAP7_75t_L g1397 ( 
.A(n_1324),
.B(n_1282),
.Y(n_1397)
);

INVx1_ASAP7_75t_L g1398 ( 
.A(n_1313),
.Y(n_1398)
);

INVx1_ASAP7_75t_L g1399 ( 
.A(n_1313),
.Y(n_1399)
);

INVx1_ASAP7_75t_L g1400 ( 
.A(n_1315),
.Y(n_1400)
);

AOI21x1_ASAP7_75t_L g1401 ( 
.A1(n_1279),
.A2(n_1275),
.B(n_1254),
.Y(n_1401)
);

INVxp33_ASAP7_75t_L g1402 ( 
.A(n_1289),
.Y(n_1402)
);

INVx1_ASAP7_75t_L g1403 ( 
.A(n_1315),
.Y(n_1403)
);

BUFx2_ASAP7_75t_L g1404 ( 
.A(n_1336),
.Y(n_1404)
);

BUFx2_ASAP7_75t_L g1405 ( 
.A(n_1336),
.Y(n_1405)
);

INVx1_ASAP7_75t_L g1406 ( 
.A(n_1301),
.Y(n_1406)
);

NAND2x1p5_ASAP7_75t_L g1407 ( 
.A(n_1336),
.B(n_1339),
.Y(n_1407)
);

HB1xp67_ASAP7_75t_L g1408 ( 
.A(n_1311),
.Y(n_1408)
);

OAI21x1_ASAP7_75t_L g1409 ( 
.A1(n_1314),
.A2(n_1339),
.B(n_1295),
.Y(n_1409)
);

BUFx3_ASAP7_75t_L g1410 ( 
.A(n_1287),
.Y(n_1410)
);

CKINVDCx20_ASAP7_75t_R g1411 ( 
.A(n_1272),
.Y(n_1411)
);

NOR2xp33_ASAP7_75t_L g1412 ( 
.A(n_1334),
.B(n_1299),
.Y(n_1412)
);

AND2x2_ASAP7_75t_L g1413 ( 
.A(n_1353),
.B(n_1294),
.Y(n_1413)
);

AND2x2_ASAP7_75t_L g1414 ( 
.A(n_1353),
.B(n_1333),
.Y(n_1414)
);

HB1xp67_ASAP7_75t_L g1415 ( 
.A(n_1343),
.Y(n_1415)
);

AOI22xp33_ASAP7_75t_L g1416 ( 
.A1(n_1384),
.A2(n_1341),
.B1(n_1323),
.B2(n_1259),
.Y(n_1416)
);

OR2x2_ASAP7_75t_L g1417 ( 
.A(n_1351),
.B(n_1278),
.Y(n_1417)
);

INVx2_ASAP7_75t_SL g1418 ( 
.A(n_1346),
.Y(n_1418)
);

NAND2xp5_ASAP7_75t_L g1419 ( 
.A(n_1350),
.B(n_1322),
.Y(n_1419)
);

BUFx2_ASAP7_75t_L g1420 ( 
.A(n_1346),
.Y(n_1420)
);

BUFx6f_ASAP7_75t_L g1421 ( 
.A(n_1344),
.Y(n_1421)
);

NAND2xp5_ASAP7_75t_L g1422 ( 
.A(n_1350),
.B(n_1265),
.Y(n_1422)
);

OR2x2_ASAP7_75t_L g1423 ( 
.A(n_1351),
.B(n_1292),
.Y(n_1423)
);

AND2x2_ASAP7_75t_L g1424 ( 
.A(n_1371),
.B(n_1312),
.Y(n_1424)
);

AOI22xp5_ASAP7_75t_L g1425 ( 
.A1(n_1384),
.A2(n_1368),
.B1(n_1359),
.B2(n_1349),
.Y(n_1425)
);

INVx1_ASAP7_75t_L g1426 ( 
.A(n_1345),
.Y(n_1426)
);

OAI22xp5_ASAP7_75t_L g1427 ( 
.A1(n_1397),
.A2(n_1287),
.B1(n_1284),
.B2(n_1334),
.Y(n_1427)
);

INVx1_ASAP7_75t_L g1428 ( 
.A(n_1354),
.Y(n_1428)
);

OR2x2_ASAP7_75t_L g1429 ( 
.A(n_1347),
.B(n_1365),
.Y(n_1429)
);

AND2x2_ASAP7_75t_L g1430 ( 
.A(n_1371),
.B(n_1308),
.Y(n_1430)
);

INVx1_ASAP7_75t_L g1431 ( 
.A(n_1354),
.Y(n_1431)
);

NAND2xp5_ASAP7_75t_L g1432 ( 
.A(n_1348),
.B(n_1316),
.Y(n_1432)
);

INVx1_ASAP7_75t_L g1433 ( 
.A(n_1358),
.Y(n_1433)
);

NAND3xp33_ASAP7_75t_L g1434 ( 
.A(n_1355),
.B(n_1293),
.C(n_1325),
.Y(n_1434)
);

AND2x2_ASAP7_75t_L g1435 ( 
.A(n_1389),
.B(n_1307),
.Y(n_1435)
);

NAND2xp5_ASAP7_75t_L g1436 ( 
.A(n_1352),
.B(n_1318),
.Y(n_1436)
);

NOR2x1_ASAP7_75t_L g1437 ( 
.A(n_1393),
.B(n_1297),
.Y(n_1437)
);

AOI22xp33_ASAP7_75t_L g1438 ( 
.A1(n_1395),
.A2(n_1335),
.B1(n_1250),
.B2(n_1328),
.Y(n_1438)
);

OR2x2_ASAP7_75t_L g1439 ( 
.A(n_1347),
.B(n_1365),
.Y(n_1439)
);

AND2x2_ASAP7_75t_L g1440 ( 
.A(n_1390),
.B(n_1317),
.Y(n_1440)
);

AND2x2_ASAP7_75t_L g1441 ( 
.A(n_1390),
.B(n_1364),
.Y(n_1441)
);

OR2x2_ASAP7_75t_L g1442 ( 
.A(n_1376),
.B(n_1319),
.Y(n_1442)
);

INVx1_ASAP7_75t_L g1443 ( 
.A(n_1358),
.Y(n_1443)
);

INVx1_ASAP7_75t_L g1444 ( 
.A(n_1361),
.Y(n_1444)
);

INVx1_ASAP7_75t_L g1445 ( 
.A(n_1361),
.Y(n_1445)
);

AND2x4_ASAP7_75t_L g1446 ( 
.A(n_1382),
.B(n_1335),
.Y(n_1446)
);

NAND2xp5_ASAP7_75t_L g1447 ( 
.A(n_1414),
.B(n_1360),
.Y(n_1447)
);

AND2x2_ASAP7_75t_L g1448 ( 
.A(n_1414),
.B(n_1441),
.Y(n_1448)
);

AND2x2_ASAP7_75t_L g1449 ( 
.A(n_1414),
.B(n_1366),
.Y(n_1449)
);

NAND3xp33_ASAP7_75t_L g1450 ( 
.A(n_1416),
.B(n_1381),
.C(n_1386),
.Y(n_1450)
);

INVx1_ASAP7_75t_L g1451 ( 
.A(n_1429),
.Y(n_1451)
);

NAND2xp5_ASAP7_75t_SL g1452 ( 
.A(n_1437),
.B(n_1413),
.Y(n_1452)
);

OAI21xp5_ASAP7_75t_SL g1453 ( 
.A1(n_1416),
.A2(n_1387),
.B(n_1401),
.Y(n_1453)
);

NAND2xp5_ASAP7_75t_L g1454 ( 
.A(n_1413),
.B(n_1363),
.Y(n_1454)
);

NAND3xp33_ASAP7_75t_L g1455 ( 
.A(n_1425),
.B(n_1386),
.C(n_1396),
.Y(n_1455)
);

NAND2xp5_ASAP7_75t_L g1456 ( 
.A(n_1419),
.B(n_1383),
.Y(n_1456)
);

INVx1_ASAP7_75t_L g1457 ( 
.A(n_1426),
.Y(n_1457)
);

NAND3xp33_ASAP7_75t_L g1458 ( 
.A(n_1425),
.B(n_1396),
.C(n_1406),
.Y(n_1458)
);

NAND2xp5_ASAP7_75t_SL g1459 ( 
.A(n_1437),
.B(n_1388),
.Y(n_1459)
);

NAND3xp33_ASAP7_75t_L g1460 ( 
.A(n_1436),
.B(n_1406),
.C(n_1377),
.Y(n_1460)
);

NAND2xp5_ASAP7_75t_L g1461 ( 
.A(n_1429),
.B(n_1370),
.Y(n_1461)
);

NAND2xp5_ASAP7_75t_L g1462 ( 
.A(n_1439),
.B(n_1378),
.Y(n_1462)
);

AND2x2_ASAP7_75t_L g1463 ( 
.A(n_1441),
.B(n_1366),
.Y(n_1463)
);

NAND2xp5_ASAP7_75t_L g1464 ( 
.A(n_1439),
.B(n_1378),
.Y(n_1464)
);

NAND3xp33_ASAP7_75t_L g1465 ( 
.A(n_1436),
.B(n_1430),
.C(n_1435),
.Y(n_1465)
);

NAND2xp5_ASAP7_75t_L g1466 ( 
.A(n_1439),
.B(n_1367),
.Y(n_1466)
);

NAND2xp5_ASAP7_75t_SL g1467 ( 
.A(n_1438),
.B(n_1388),
.Y(n_1467)
);

OAI21xp5_ASAP7_75t_SL g1468 ( 
.A1(n_1434),
.A2(n_1401),
.B(n_1412),
.Y(n_1468)
);

OAI21xp5_ASAP7_75t_SL g1469 ( 
.A1(n_1434),
.A2(n_1356),
.B(n_1404),
.Y(n_1469)
);

OAI221xp5_ASAP7_75t_SL g1470 ( 
.A1(n_1423),
.A2(n_1395),
.B1(n_1394),
.B2(n_1385),
.C(n_1404),
.Y(n_1470)
);

NAND2xp5_ASAP7_75t_L g1471 ( 
.A(n_1442),
.B(n_1369),
.Y(n_1471)
);

AOI21xp5_ASAP7_75t_SL g1472 ( 
.A1(n_1446),
.A2(n_1385),
.B(n_1394),
.Y(n_1472)
);

NAND2xp5_ASAP7_75t_L g1473 ( 
.A(n_1428),
.B(n_1372),
.Y(n_1473)
);

OAI22xp5_ASAP7_75t_L g1474 ( 
.A1(n_1438),
.A2(n_1427),
.B1(n_1423),
.B2(n_1385),
.Y(n_1474)
);

AND2x2_ASAP7_75t_L g1475 ( 
.A(n_1440),
.B(n_1388),
.Y(n_1475)
);

NAND2xp5_ASAP7_75t_L g1476 ( 
.A(n_1428),
.B(n_1372),
.Y(n_1476)
);

OAI21xp5_ASAP7_75t_L g1477 ( 
.A1(n_1427),
.A2(n_1392),
.B(n_1409),
.Y(n_1477)
);

NAND2xp5_ASAP7_75t_L g1478 ( 
.A(n_1431),
.B(n_1373),
.Y(n_1478)
);

NAND3xp33_ASAP7_75t_L g1479 ( 
.A(n_1430),
.B(n_1408),
.C(n_1398),
.Y(n_1479)
);

NAND2xp5_ASAP7_75t_L g1480 ( 
.A(n_1431),
.B(n_1373),
.Y(n_1480)
);

NAND2xp5_ASAP7_75t_L g1481 ( 
.A(n_1433),
.B(n_1375),
.Y(n_1481)
);

NAND2xp5_ASAP7_75t_L g1482 ( 
.A(n_1433),
.B(n_1375),
.Y(n_1482)
);

NAND3xp33_ASAP7_75t_L g1483 ( 
.A(n_1430),
.B(n_1398),
.C(n_1399),
.Y(n_1483)
);

AOI221xp5_ASAP7_75t_L g1484 ( 
.A1(n_1423),
.A2(n_1379),
.B1(n_1380),
.B2(n_1402),
.C(n_1357),
.Y(n_1484)
);

NAND3xp33_ASAP7_75t_L g1485 ( 
.A(n_1435),
.B(n_1399),
.C(n_1400),
.Y(n_1485)
);

OAI221xp5_ASAP7_75t_L g1486 ( 
.A1(n_1422),
.A2(n_1362),
.B1(n_1407),
.B2(n_1405),
.C(n_1379),
.Y(n_1486)
);

NAND3xp33_ASAP7_75t_L g1487 ( 
.A(n_1435),
.B(n_1400),
.C(n_1403),
.Y(n_1487)
);

BUFx2_ASAP7_75t_L g1488 ( 
.A(n_1448),
.Y(n_1488)
);

AND3x1_ASAP7_75t_L g1489 ( 
.A(n_1453),
.B(n_1374),
.C(n_1418),
.Y(n_1489)
);

INVx1_ASAP7_75t_L g1490 ( 
.A(n_1457),
.Y(n_1490)
);

NOR2xp67_ASAP7_75t_L g1491 ( 
.A(n_1465),
.B(n_1415),
.Y(n_1491)
);

INVx2_ASAP7_75t_L g1492 ( 
.A(n_1457),
.Y(n_1492)
);

HB1xp67_ASAP7_75t_L g1493 ( 
.A(n_1485),
.Y(n_1493)
);

OR2x2_ASAP7_75t_L g1494 ( 
.A(n_1454),
.B(n_1432),
.Y(n_1494)
);

NAND2xp5_ASAP7_75t_L g1495 ( 
.A(n_1451),
.B(n_1443),
.Y(n_1495)
);

INVx2_ASAP7_75t_L g1496 ( 
.A(n_1463),
.Y(n_1496)
);

INVx1_ASAP7_75t_L g1497 ( 
.A(n_1483),
.Y(n_1497)
);

NAND2xp5_ASAP7_75t_L g1498 ( 
.A(n_1449),
.B(n_1443),
.Y(n_1498)
);

NAND2xp5_ASAP7_75t_L g1499 ( 
.A(n_1456),
.B(n_1444),
.Y(n_1499)
);

OR2x2_ASAP7_75t_L g1500 ( 
.A(n_1447),
.B(n_1417),
.Y(n_1500)
);

INVx5_ASAP7_75t_L g1501 ( 
.A(n_1475),
.Y(n_1501)
);

INVx2_ASAP7_75t_L g1502 ( 
.A(n_1487),
.Y(n_1502)
);

HB1xp67_ASAP7_75t_L g1503 ( 
.A(n_1460),
.Y(n_1503)
);

NOR2xp33_ASAP7_75t_L g1504 ( 
.A(n_1469),
.B(n_1362),
.Y(n_1504)
);

NAND2xp5_ASAP7_75t_L g1505 ( 
.A(n_1471),
.B(n_1466),
.Y(n_1505)
);

INVx1_ASAP7_75t_L g1506 ( 
.A(n_1473),
.Y(n_1506)
);

NAND2xp5_ASAP7_75t_L g1507 ( 
.A(n_1461),
.B(n_1445),
.Y(n_1507)
);

INVx1_ASAP7_75t_L g1508 ( 
.A(n_1476),
.Y(n_1508)
);

BUFx3_ASAP7_75t_L g1509 ( 
.A(n_1486),
.Y(n_1509)
);

HB1xp67_ASAP7_75t_L g1510 ( 
.A(n_1479),
.Y(n_1510)
);

AND2x2_ASAP7_75t_L g1511 ( 
.A(n_1462),
.B(n_1464),
.Y(n_1511)
);

HB1xp67_ASAP7_75t_L g1512 ( 
.A(n_1478),
.Y(n_1512)
);

AND2x2_ASAP7_75t_L g1513 ( 
.A(n_1477),
.B(n_1424),
.Y(n_1513)
);

AND3x2_ASAP7_75t_L g1514 ( 
.A(n_1503),
.B(n_1472),
.C(n_1484),
.Y(n_1514)
);

INVx2_ASAP7_75t_SL g1515 ( 
.A(n_1501),
.Y(n_1515)
);

OAI22xp5_ASAP7_75t_L g1516 ( 
.A1(n_1489),
.A2(n_1450),
.B1(n_1455),
.B2(n_1458),
.Y(n_1516)
);

HB1xp67_ASAP7_75t_L g1517 ( 
.A(n_1493),
.Y(n_1517)
);

OAI221xp5_ASAP7_75t_SL g1518 ( 
.A1(n_1489),
.A2(n_1468),
.B1(n_1417),
.B2(n_1394),
.C(n_1391),
.Y(n_1518)
);

AND2x2_ASAP7_75t_L g1519 ( 
.A(n_1488),
.B(n_1459),
.Y(n_1519)
);

AND2x2_ASAP7_75t_L g1520 ( 
.A(n_1488),
.B(n_1452),
.Y(n_1520)
);

INVx2_ASAP7_75t_L g1521 ( 
.A(n_1492),
.Y(n_1521)
);

NAND2xp5_ASAP7_75t_L g1522 ( 
.A(n_1497),
.B(n_1452),
.Y(n_1522)
);

NAND2xp5_ASAP7_75t_L g1523 ( 
.A(n_1497),
.B(n_1480),
.Y(n_1523)
);

BUFx2_ASAP7_75t_L g1524 ( 
.A(n_1493),
.Y(n_1524)
);

NOR2xp33_ASAP7_75t_L g1525 ( 
.A(n_1503),
.B(n_1411),
.Y(n_1525)
);

NAND2xp5_ASAP7_75t_L g1526 ( 
.A(n_1497),
.B(n_1481),
.Y(n_1526)
);

NOR2x1_ASAP7_75t_L g1527 ( 
.A(n_1509),
.B(n_1393),
.Y(n_1527)
);

OR2x2_ASAP7_75t_L g1528 ( 
.A(n_1500),
.B(n_1482),
.Y(n_1528)
);

INVx2_ASAP7_75t_L g1529 ( 
.A(n_1492),
.Y(n_1529)
);

HB1xp67_ASAP7_75t_L g1530 ( 
.A(n_1502),
.Y(n_1530)
);

OAI21xp33_ASAP7_75t_L g1531 ( 
.A1(n_1510),
.A2(n_1467),
.B(n_1421),
.Y(n_1531)
);

OR2x2_ASAP7_75t_L g1532 ( 
.A(n_1500),
.B(n_1417),
.Y(n_1532)
);

INVx1_ASAP7_75t_L g1533 ( 
.A(n_1490),
.Y(n_1533)
);

INVx1_ASAP7_75t_L g1534 ( 
.A(n_1490),
.Y(n_1534)
);

NOR2xp33_ASAP7_75t_L g1535 ( 
.A(n_1509),
.B(n_1272),
.Y(n_1535)
);

NAND2xp5_ASAP7_75t_L g1536 ( 
.A(n_1502),
.B(n_1512),
.Y(n_1536)
);

INVx2_ASAP7_75t_L g1537 ( 
.A(n_1492),
.Y(n_1537)
);

INVx1_ASAP7_75t_L g1538 ( 
.A(n_1490),
.Y(n_1538)
);

AOI211xp5_ASAP7_75t_L g1539 ( 
.A1(n_1509),
.A2(n_1467),
.B(n_1474),
.C(n_1470),
.Y(n_1539)
);

INVx1_ASAP7_75t_L g1540 ( 
.A(n_1512),
.Y(n_1540)
);

NAND2xp5_ASAP7_75t_SL g1541 ( 
.A(n_1509),
.B(n_1501),
.Y(n_1541)
);

AND2x2_ASAP7_75t_L g1542 ( 
.A(n_1488),
.B(n_1420),
.Y(n_1542)
);

NAND2xp5_ASAP7_75t_L g1543 ( 
.A(n_1502),
.B(n_1510),
.Y(n_1543)
);

INVx1_ASAP7_75t_L g1544 ( 
.A(n_1506),
.Y(n_1544)
);

INVx1_ASAP7_75t_L g1545 ( 
.A(n_1506),
.Y(n_1545)
);

INVx2_ASAP7_75t_L g1546 ( 
.A(n_1496),
.Y(n_1546)
);

INVx1_ASAP7_75t_L g1547 ( 
.A(n_1495),
.Y(n_1547)
);

INVx1_ASAP7_75t_L g1548 ( 
.A(n_1495),
.Y(n_1548)
);

INVx2_ASAP7_75t_L g1549 ( 
.A(n_1546),
.Y(n_1549)
);

AOI221xp5_ASAP7_75t_L g1550 ( 
.A1(n_1516),
.A2(n_1502),
.B1(n_1513),
.B2(n_1504),
.C(n_1499),
.Y(n_1550)
);

INVx2_ASAP7_75t_L g1551 ( 
.A(n_1546),
.Y(n_1551)
);

AND2x2_ASAP7_75t_L g1552 ( 
.A(n_1520),
.B(n_1501),
.Y(n_1552)
);

NAND2xp5_ASAP7_75t_L g1553 ( 
.A(n_1524),
.B(n_1500),
.Y(n_1553)
);

NOR2xp33_ASAP7_75t_L g1554 ( 
.A(n_1535),
.B(n_1326),
.Y(n_1554)
);

INVx2_ASAP7_75t_SL g1555 ( 
.A(n_1520),
.Y(n_1555)
);

AND2x2_ASAP7_75t_L g1556 ( 
.A(n_1519),
.B(n_1501),
.Y(n_1556)
);

AOI21xp33_ASAP7_75t_L g1557 ( 
.A1(n_1543),
.A2(n_1504),
.B(n_1499),
.Y(n_1557)
);

INVx1_ASAP7_75t_L g1558 ( 
.A(n_1533),
.Y(n_1558)
);

INVx1_ASAP7_75t_L g1559 ( 
.A(n_1533),
.Y(n_1559)
);

INVx1_ASAP7_75t_L g1560 ( 
.A(n_1534),
.Y(n_1560)
);

INVx1_ASAP7_75t_L g1561 ( 
.A(n_1534),
.Y(n_1561)
);

INVx1_ASAP7_75t_L g1562 ( 
.A(n_1538),
.Y(n_1562)
);

NAND2xp33_ASAP7_75t_L g1563 ( 
.A(n_1516),
.B(n_1326),
.Y(n_1563)
);

AND2x2_ASAP7_75t_L g1564 ( 
.A(n_1519),
.B(n_1501),
.Y(n_1564)
);

OR2x2_ASAP7_75t_L g1565 ( 
.A(n_1543),
.B(n_1505),
.Y(n_1565)
);

OR2x2_ASAP7_75t_L g1566 ( 
.A(n_1536),
.B(n_1505),
.Y(n_1566)
);

INVx3_ASAP7_75t_L g1567 ( 
.A(n_1515),
.Y(n_1567)
);

HB1xp67_ASAP7_75t_L g1568 ( 
.A(n_1530),
.Y(n_1568)
);

INVx1_ASAP7_75t_L g1569 ( 
.A(n_1538),
.Y(n_1569)
);

INVx1_ASAP7_75t_L g1570 ( 
.A(n_1544),
.Y(n_1570)
);

AND2x2_ASAP7_75t_L g1571 ( 
.A(n_1541),
.B(n_1501),
.Y(n_1571)
);

NAND2xp5_ASAP7_75t_L g1572 ( 
.A(n_1524),
.B(n_1508),
.Y(n_1572)
);

INVxp67_ASAP7_75t_L g1573 ( 
.A(n_1525),
.Y(n_1573)
);

INVx2_ASAP7_75t_L g1574 ( 
.A(n_1546),
.Y(n_1574)
);

OR2x2_ASAP7_75t_L g1575 ( 
.A(n_1536),
.B(n_1494),
.Y(n_1575)
);

INVx1_ASAP7_75t_L g1576 ( 
.A(n_1544),
.Y(n_1576)
);

INVx1_ASAP7_75t_L g1577 ( 
.A(n_1545),
.Y(n_1577)
);

NAND2xp5_ASAP7_75t_L g1578 ( 
.A(n_1517),
.B(n_1508),
.Y(n_1578)
);

NOR2x1p5_ASAP7_75t_SL g1579 ( 
.A(n_1521),
.B(n_1508),
.Y(n_1579)
);

INVx1_ASAP7_75t_L g1580 ( 
.A(n_1545),
.Y(n_1580)
);

NAND2xp5_ASAP7_75t_L g1581 ( 
.A(n_1517),
.B(n_1511),
.Y(n_1581)
);

NOR2xp33_ASAP7_75t_L g1582 ( 
.A(n_1522),
.B(n_1507),
.Y(n_1582)
);

NOR2xp33_ASAP7_75t_L g1583 ( 
.A(n_1522),
.B(n_1507),
.Y(n_1583)
);

AND2x2_ASAP7_75t_L g1584 ( 
.A(n_1542),
.B(n_1501),
.Y(n_1584)
);

BUFx8_ASAP7_75t_SL g1585 ( 
.A(n_1523),
.Y(n_1585)
);

INVx2_ASAP7_75t_L g1586 ( 
.A(n_1521),
.Y(n_1586)
);

INVx1_ASAP7_75t_L g1587 ( 
.A(n_1540),
.Y(n_1587)
);

OR2x2_ASAP7_75t_L g1588 ( 
.A(n_1523),
.B(n_1494),
.Y(n_1588)
);

NOR2xp33_ASAP7_75t_L g1589 ( 
.A(n_1526),
.B(n_1498),
.Y(n_1589)
);

AND2x2_ASAP7_75t_L g1590 ( 
.A(n_1542),
.B(n_1501),
.Y(n_1590)
);

AND2x2_ASAP7_75t_L g1591 ( 
.A(n_1515),
.B(n_1501),
.Y(n_1591)
);

INVx2_ASAP7_75t_L g1592 ( 
.A(n_1555),
.Y(n_1592)
);

INVx1_ASAP7_75t_SL g1593 ( 
.A(n_1585),
.Y(n_1593)
);

INVx2_ASAP7_75t_SL g1594 ( 
.A(n_1555),
.Y(n_1594)
);

INVx1_ASAP7_75t_L g1595 ( 
.A(n_1558),
.Y(n_1595)
);

AOI222xp33_ASAP7_75t_L g1596 ( 
.A1(n_1563),
.A2(n_1531),
.B1(n_1530),
.B2(n_1491),
.C1(n_1526),
.C2(n_1513),
.Y(n_1596)
);

OR2x2_ASAP7_75t_L g1597 ( 
.A(n_1565),
.B(n_1575),
.Y(n_1597)
);

NAND2xp5_ASAP7_75t_L g1598 ( 
.A(n_1582),
.B(n_1540),
.Y(n_1598)
);

INVx1_ASAP7_75t_SL g1599 ( 
.A(n_1554),
.Y(n_1599)
);

INVx3_ASAP7_75t_L g1600 ( 
.A(n_1567),
.Y(n_1600)
);

INVx1_ASAP7_75t_L g1601 ( 
.A(n_1558),
.Y(n_1601)
);

AND2x2_ASAP7_75t_L g1602 ( 
.A(n_1552),
.B(n_1515),
.Y(n_1602)
);

NAND2xp5_ASAP7_75t_L g1603 ( 
.A(n_1583),
.B(n_1528),
.Y(n_1603)
);

NAND2xp5_ASAP7_75t_L g1604 ( 
.A(n_1589),
.B(n_1528),
.Y(n_1604)
);

NAND2xp5_ASAP7_75t_L g1605 ( 
.A(n_1565),
.B(n_1547),
.Y(n_1605)
);

OR2x2_ASAP7_75t_L g1606 ( 
.A(n_1575),
.B(n_1547),
.Y(n_1606)
);

INVx1_ASAP7_75t_L g1607 ( 
.A(n_1559),
.Y(n_1607)
);

AND2x2_ASAP7_75t_L g1608 ( 
.A(n_1552),
.B(n_1527),
.Y(n_1608)
);

INVx1_ASAP7_75t_L g1609 ( 
.A(n_1559),
.Y(n_1609)
);

OA21x2_ASAP7_75t_L g1610 ( 
.A1(n_1550),
.A2(n_1531),
.B(n_1529),
.Y(n_1610)
);

NAND2xp5_ASAP7_75t_L g1611 ( 
.A(n_1581),
.B(n_1548),
.Y(n_1611)
);

INVx2_ASAP7_75t_L g1612 ( 
.A(n_1549),
.Y(n_1612)
);

INVx1_ASAP7_75t_SL g1613 ( 
.A(n_1553),
.Y(n_1613)
);

INVx2_ASAP7_75t_L g1614 ( 
.A(n_1549),
.Y(n_1614)
);

INVx4_ASAP7_75t_L g1615 ( 
.A(n_1568),
.Y(n_1615)
);

CKINVDCx16_ASAP7_75t_R g1616 ( 
.A(n_1571),
.Y(n_1616)
);

NAND3xp33_ASAP7_75t_L g1617 ( 
.A(n_1572),
.B(n_1539),
.C(n_1518),
.Y(n_1617)
);

NAND2xp5_ASAP7_75t_L g1618 ( 
.A(n_1566),
.B(n_1548),
.Y(n_1618)
);

INVx2_ASAP7_75t_L g1619 ( 
.A(n_1551),
.Y(n_1619)
);

OR2x2_ASAP7_75t_L g1620 ( 
.A(n_1588),
.B(n_1532),
.Y(n_1620)
);

INVxp67_ASAP7_75t_SL g1621 ( 
.A(n_1573),
.Y(n_1621)
);

NOR2xp33_ASAP7_75t_L g1622 ( 
.A(n_1566),
.B(n_1527),
.Y(n_1622)
);

HB1xp67_ASAP7_75t_L g1623 ( 
.A(n_1587),
.Y(n_1623)
);

INVx1_ASAP7_75t_L g1624 ( 
.A(n_1560),
.Y(n_1624)
);

NAND2xp5_ASAP7_75t_L g1625 ( 
.A(n_1588),
.B(n_1539),
.Y(n_1625)
);

INVx1_ASAP7_75t_L g1626 ( 
.A(n_1560),
.Y(n_1626)
);

INVx1_ASAP7_75t_SL g1627 ( 
.A(n_1587),
.Y(n_1627)
);

OAI22xp5_ASAP7_75t_L g1628 ( 
.A1(n_1617),
.A2(n_1518),
.B1(n_1491),
.B2(n_1557),
.Y(n_1628)
);

INVx4_ASAP7_75t_L g1629 ( 
.A(n_1615),
.Y(n_1629)
);

AOI22xp5_ASAP7_75t_L g1630 ( 
.A1(n_1617),
.A2(n_1514),
.B1(n_1513),
.B2(n_1532),
.Y(n_1630)
);

INVx1_ASAP7_75t_L g1631 ( 
.A(n_1623),
.Y(n_1631)
);

BUFx2_ASAP7_75t_SL g1632 ( 
.A(n_1593),
.Y(n_1632)
);

OAI22xp33_ASAP7_75t_L g1633 ( 
.A1(n_1625),
.A2(n_1578),
.B1(n_1514),
.B2(n_1576),
.Y(n_1633)
);

INVx1_ASAP7_75t_L g1634 ( 
.A(n_1595),
.Y(n_1634)
);

NAND2xp5_ASAP7_75t_L g1635 ( 
.A(n_1627),
.B(n_1570),
.Y(n_1635)
);

NOR2xp67_ASAP7_75t_L g1636 ( 
.A(n_1594),
.B(n_1571),
.Y(n_1636)
);

AND2x2_ASAP7_75t_L g1637 ( 
.A(n_1593),
.B(n_1556),
.Y(n_1637)
);

AND2x4_ASAP7_75t_L g1638 ( 
.A(n_1594),
.B(n_1556),
.Y(n_1638)
);

INVx1_ASAP7_75t_L g1639 ( 
.A(n_1595),
.Y(n_1639)
);

OAI21xp5_ASAP7_75t_L g1640 ( 
.A1(n_1621),
.A2(n_1576),
.B(n_1570),
.Y(n_1640)
);

INVx1_ASAP7_75t_L g1641 ( 
.A(n_1601),
.Y(n_1641)
);

INVx2_ASAP7_75t_L g1642 ( 
.A(n_1600),
.Y(n_1642)
);

INVx1_ASAP7_75t_L g1643 ( 
.A(n_1601),
.Y(n_1643)
);

INVx1_ASAP7_75t_L g1644 ( 
.A(n_1607),
.Y(n_1644)
);

INVx1_ASAP7_75t_L g1645 ( 
.A(n_1607),
.Y(n_1645)
);

INVx2_ASAP7_75t_L g1646 ( 
.A(n_1600),
.Y(n_1646)
);

OAI22xp33_ASAP7_75t_SL g1647 ( 
.A1(n_1616),
.A2(n_1579),
.B1(n_1551),
.B2(n_1574),
.Y(n_1647)
);

OAI221xp5_ASAP7_75t_L g1648 ( 
.A1(n_1610),
.A2(n_1586),
.B1(n_1577),
.B2(n_1580),
.C(n_1574),
.Y(n_1648)
);

AOI222xp33_ASAP7_75t_L g1649 ( 
.A1(n_1613),
.A2(n_1579),
.B1(n_1580),
.B2(n_1577),
.C1(n_1586),
.C2(n_1562),
.Y(n_1649)
);

OAI21xp5_ASAP7_75t_SL g1650 ( 
.A1(n_1596),
.A2(n_1564),
.B(n_1591),
.Y(n_1650)
);

AND2x2_ASAP7_75t_L g1651 ( 
.A(n_1616),
.B(n_1564),
.Y(n_1651)
);

AOI22xp5_ASAP7_75t_L g1652 ( 
.A1(n_1610),
.A2(n_1599),
.B1(n_1622),
.B2(n_1614),
.Y(n_1652)
);

AOI211xp5_ASAP7_75t_L g1653 ( 
.A1(n_1627),
.A2(n_1591),
.B(n_1569),
.C(n_1562),
.Y(n_1653)
);

NAND2xp33_ASAP7_75t_SL g1654 ( 
.A(n_1637),
.B(n_1615),
.Y(n_1654)
);

OR2x6_ASAP7_75t_L g1655 ( 
.A(n_1632),
.B(n_1592),
.Y(n_1655)
);

NOR2xp33_ASAP7_75t_L g1656 ( 
.A(n_1629),
.B(n_1599),
.Y(n_1656)
);

INVx1_ASAP7_75t_L g1657 ( 
.A(n_1635),
.Y(n_1657)
);

INVxp67_ASAP7_75t_L g1658 ( 
.A(n_1651),
.Y(n_1658)
);

HB1xp67_ASAP7_75t_L g1659 ( 
.A(n_1642),
.Y(n_1659)
);

NAND2xp5_ASAP7_75t_L g1660 ( 
.A(n_1631),
.B(n_1592),
.Y(n_1660)
);

NAND2xp5_ASAP7_75t_L g1661 ( 
.A(n_1653),
.B(n_1597),
.Y(n_1661)
);

NAND2xp5_ASAP7_75t_L g1662 ( 
.A(n_1652),
.B(n_1597),
.Y(n_1662)
);

AND2x2_ASAP7_75t_L g1663 ( 
.A(n_1638),
.B(n_1608),
.Y(n_1663)
);

AND2x2_ASAP7_75t_L g1664 ( 
.A(n_1638),
.B(n_1608),
.Y(n_1664)
);

INVx1_ASAP7_75t_L g1665 ( 
.A(n_1634),
.Y(n_1665)
);

AND2x2_ASAP7_75t_L g1666 ( 
.A(n_1636),
.B(n_1602),
.Y(n_1666)
);

INVx1_ASAP7_75t_L g1667 ( 
.A(n_1639),
.Y(n_1667)
);

HB1xp67_ASAP7_75t_L g1668 ( 
.A(n_1646),
.Y(n_1668)
);

INVxp67_ASAP7_75t_SL g1669 ( 
.A(n_1647),
.Y(n_1669)
);

HB1xp67_ASAP7_75t_L g1670 ( 
.A(n_1629),
.Y(n_1670)
);

INVx1_ASAP7_75t_L g1671 ( 
.A(n_1641),
.Y(n_1671)
);

INVx1_ASAP7_75t_L g1672 ( 
.A(n_1635),
.Y(n_1672)
);

NAND3xp33_ASAP7_75t_L g1673 ( 
.A(n_1669),
.B(n_1648),
.C(n_1649),
.Y(n_1673)
);

AOI321xp33_ASAP7_75t_L g1674 ( 
.A1(n_1662),
.A2(n_1648),
.A3(n_1633),
.B1(n_1630),
.B2(n_1628),
.C(n_1643),
.Y(n_1674)
);

NAND4xp25_ASAP7_75t_L g1675 ( 
.A(n_1656),
.B(n_1640),
.C(n_1650),
.D(n_1615),
.Y(n_1675)
);

NOR2xp33_ASAP7_75t_SL g1676 ( 
.A(n_1658),
.B(n_1615),
.Y(n_1676)
);

NAND3xp33_ASAP7_75t_L g1677 ( 
.A(n_1655),
.B(n_1628),
.C(n_1640),
.Y(n_1677)
);

OR2x2_ASAP7_75t_L g1678 ( 
.A(n_1661),
.B(n_1655),
.Y(n_1678)
);

NAND3xp33_ASAP7_75t_L g1679 ( 
.A(n_1655),
.B(n_1610),
.C(n_1633),
.Y(n_1679)
);

OAI21xp5_ASAP7_75t_L g1680 ( 
.A1(n_1655),
.A2(n_1610),
.B(n_1598),
.Y(n_1680)
);

OAI21xp5_ASAP7_75t_SL g1681 ( 
.A1(n_1666),
.A2(n_1602),
.B(n_1600),
.Y(n_1681)
);

NOR4xp25_ASAP7_75t_L g1682 ( 
.A(n_1657),
.B(n_1645),
.C(n_1644),
.D(n_1626),
.Y(n_1682)
);

NOR2x1_ASAP7_75t_SL g1683 ( 
.A(n_1679),
.B(n_1663),
.Y(n_1683)
);

NAND3xp33_ASAP7_75t_L g1684 ( 
.A(n_1674),
.B(n_1673),
.C(n_1677),
.Y(n_1684)
);

NAND5xp2_ASAP7_75t_L g1685 ( 
.A(n_1680),
.B(n_1666),
.C(n_1664),
.D(n_1663),
.E(n_1657),
.Y(n_1685)
);

OR2x2_ASAP7_75t_L g1686 ( 
.A(n_1678),
.B(n_1660),
.Y(n_1686)
);

AOI211xp5_ASAP7_75t_L g1687 ( 
.A1(n_1682),
.A2(n_1672),
.B(n_1659),
.C(n_1668),
.Y(n_1687)
);

A2O1A1Ixp33_ASAP7_75t_L g1688 ( 
.A1(n_1675),
.A2(n_1672),
.B(n_1654),
.C(n_1671),
.Y(n_1688)
);

AND5x1_ASAP7_75t_L g1689 ( 
.A(n_1676),
.B(n_1654),
.C(n_1664),
.D(n_1670),
.E(n_1665),
.Y(n_1689)
);

INVx1_ASAP7_75t_L g1690 ( 
.A(n_1681),
.Y(n_1690)
);

NAND2xp5_ASAP7_75t_L g1691 ( 
.A(n_1676),
.B(n_1667),
.Y(n_1691)
);

AOI221x1_ASAP7_75t_L g1692 ( 
.A1(n_1684),
.A2(n_1626),
.B1(n_1624),
.B2(n_1609),
.C(n_1619),
.Y(n_1692)
);

NAND4xp25_ASAP7_75t_L g1693 ( 
.A(n_1685),
.B(n_1624),
.C(n_1609),
.D(n_1605),
.Y(n_1693)
);

NAND3xp33_ASAP7_75t_L g1694 ( 
.A(n_1687),
.B(n_1618),
.C(n_1620),
.Y(n_1694)
);

NOR4xp25_ASAP7_75t_L g1695 ( 
.A(n_1688),
.B(n_1690),
.C(n_1686),
.D(n_1691),
.Y(n_1695)
);

NOR3xp33_ASAP7_75t_L g1696 ( 
.A(n_1683),
.B(n_1614),
.C(n_1612),
.Y(n_1696)
);

AOI22xp5_ASAP7_75t_L g1697 ( 
.A1(n_1696),
.A2(n_1619),
.B1(n_1612),
.B2(n_1620),
.Y(n_1697)
);

CKINVDCx20_ASAP7_75t_R g1698 ( 
.A(n_1694),
.Y(n_1698)
);

INVxp67_ASAP7_75t_L g1699 ( 
.A(n_1692),
.Y(n_1699)
);

INVx1_ASAP7_75t_L g1700 ( 
.A(n_1693),
.Y(n_1700)
);

INVx1_ASAP7_75t_L g1701 ( 
.A(n_1695),
.Y(n_1701)
);

INVxp67_ASAP7_75t_SL g1702 ( 
.A(n_1696),
.Y(n_1702)
);

AOI32xp33_ASAP7_75t_L g1703 ( 
.A1(n_1701),
.A2(n_1689),
.A3(n_1567),
.B1(n_1611),
.B2(n_1603),
.Y(n_1703)
);

NOR3xp33_ASAP7_75t_L g1704 ( 
.A(n_1702),
.B(n_1606),
.C(n_1604),
.Y(n_1704)
);

OAI211xp5_ASAP7_75t_SL g1705 ( 
.A1(n_1699),
.A2(n_1606),
.B(n_1567),
.C(n_1561),
.Y(n_1705)
);

INVx1_ASAP7_75t_L g1706 ( 
.A(n_1697),
.Y(n_1706)
);

INVx1_ASAP7_75t_L g1707 ( 
.A(n_1698),
.Y(n_1707)
);

INVx2_ASAP7_75t_L g1708 ( 
.A(n_1707),
.Y(n_1708)
);

BUFx6f_ASAP7_75t_L g1709 ( 
.A(n_1706),
.Y(n_1709)
);

INVx3_ASAP7_75t_L g1710 ( 
.A(n_1705),
.Y(n_1710)
);

OAI22xp33_ASAP7_75t_L g1711 ( 
.A1(n_1710),
.A2(n_1700),
.B1(n_1704),
.B2(n_1703),
.Y(n_1711)
);

OAI211xp5_ASAP7_75t_L g1712 ( 
.A1(n_1711),
.A2(n_1708),
.B(n_1710),
.C(n_1709),
.Y(n_1712)
);

HB1xp67_ASAP7_75t_L g1713 ( 
.A(n_1712),
.Y(n_1713)
);

INVx2_ASAP7_75t_L g1714 ( 
.A(n_1712),
.Y(n_1714)
);

INVx2_ASAP7_75t_L g1715 ( 
.A(n_1714),
.Y(n_1715)
);

AOI21xp5_ASAP7_75t_SL g1716 ( 
.A1(n_1713),
.A2(n_1708),
.B(n_1709),
.Y(n_1716)
);

OAI22xp5_ASAP7_75t_L g1717 ( 
.A1(n_1715),
.A2(n_1710),
.B1(n_1709),
.B2(n_1567),
.Y(n_1717)
);

OAI21xp5_ASAP7_75t_L g1718 ( 
.A1(n_1716),
.A2(n_1709),
.B(n_1569),
.Y(n_1718)
);

HB1xp67_ASAP7_75t_L g1719 ( 
.A(n_1717),
.Y(n_1719)
);

OAI22xp33_ASAP7_75t_L g1720 ( 
.A1(n_1719),
.A2(n_1718),
.B1(n_1561),
.B2(n_1537),
.Y(n_1720)
);

OAI221xp5_ASAP7_75t_R g1721 ( 
.A1(n_1720),
.A2(n_1325),
.B1(n_1584),
.B2(n_1590),
.C(n_1299),
.Y(n_1721)
);

AOI211xp5_ASAP7_75t_L g1722 ( 
.A1(n_1721),
.A2(n_1410),
.B(n_1590),
.C(n_1584),
.Y(n_1722)
);


endmodule