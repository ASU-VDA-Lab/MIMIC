module fake_netlist_1_11139_n_309 (n_44, n_81, n_69, n_22, n_57, n_88, n_52, n_26, n_50, n_33, n_102, n_73, n_49, n_97, n_80, n_60, n_41, n_35, n_94, n_65, n_9, n_10, n_103, n_19, n_87, n_98, n_74, n_7, n_29, n_45, n_85, n_101, n_62, n_36, n_47, n_37, n_34, n_5, n_23, n_8, n_91, n_16, n_13, n_95, n_70, n_17, n_63, n_14, n_71, n_90, n_56, n_42, n_24, n_78, n_6, n_4, n_40, n_79, n_38, n_64, n_46, n_31, n_58, n_32, n_0, n_84, n_55, n_12, n_86, n_75, n_72, n_43, n_76, n_89, n_68, n_27, n_53, n_67, n_77, n_20, n_2, n_54, n_83, n_28, n_48, n_100, n_92, n_11, n_25, n_30, n_59, n_3, n_18, n_66, n_1, n_82, n_15, n_61, n_21, n_99, n_93, n_51, n_96, n_39, n_309);
input n_44;
input n_81;
input n_69;
input n_22;
input n_57;
input n_88;
input n_52;
input n_26;
input n_50;
input n_33;
input n_102;
input n_73;
input n_49;
input n_97;
input n_80;
input n_60;
input n_41;
input n_35;
input n_94;
input n_65;
input n_9;
input n_10;
input n_103;
input n_19;
input n_87;
input n_98;
input n_74;
input n_7;
input n_29;
input n_45;
input n_85;
input n_101;
input n_62;
input n_36;
input n_47;
input n_37;
input n_34;
input n_5;
input n_23;
input n_8;
input n_91;
input n_16;
input n_13;
input n_95;
input n_70;
input n_17;
input n_63;
input n_14;
input n_71;
input n_90;
input n_56;
input n_42;
input n_24;
input n_78;
input n_6;
input n_4;
input n_40;
input n_79;
input n_38;
input n_64;
input n_46;
input n_31;
input n_58;
input n_32;
input n_0;
input n_84;
input n_55;
input n_12;
input n_86;
input n_75;
input n_72;
input n_43;
input n_76;
input n_89;
input n_68;
input n_27;
input n_53;
input n_67;
input n_77;
input n_20;
input n_2;
input n_54;
input n_83;
input n_28;
input n_48;
input n_100;
input n_92;
input n_11;
input n_25;
input n_30;
input n_59;
input n_3;
input n_18;
input n_66;
input n_1;
input n_82;
input n_15;
input n_61;
input n_21;
input n_99;
input n_93;
input n_51;
input n_96;
input n_39;
output n_309;
wire n_117;
wire n_185;
wire n_284;
wire n_278;
wire n_114;
wire n_125;
wire n_161;
wire n_177;
wire n_130;
wire n_189;
wire n_292;
wire n_160;
wire n_154;
wire n_229;
wire n_252;
wire n_152;
wire n_113;
wire n_206;
wire n_288;
wire n_296;
wire n_157;
wire n_202;
wire n_142;
wire n_232;
wire n_211;
wire n_275;
wire n_131;
wire n_112;
wire n_205;
wire n_162;
wire n_163;
wire n_105;
wire n_227;
wire n_231;
wire n_298;
wire n_144;
wire n_183;
wire n_199;
wire n_305;
wire n_228;
wire n_236;
wire n_150;
wire n_301;
wire n_222;
wire n_234;
wire n_286;
wire n_190;
wire n_246;
wire n_279;
wire n_303;
wire n_289;
wire n_249;
wire n_244;
wire n_141;
wire n_119;
wire n_167;
wire n_171;
wire n_196;
wire n_192;
wire n_137;
wire n_277;
wire n_250;
wire n_237;
wire n_181;
wire n_255;
wire n_108;
wire n_116;
wire n_230;
wire n_209;
wire n_274;
wire n_282;
wire n_241;
wire n_238;
wire n_293;
wire n_135;
wire n_247;
wire n_304;
wire n_294;
wire n_210;
wire n_184;
wire n_191;
wire n_307;
wire n_235;
wire n_243;
wire n_268;
wire n_174;
wire n_248;
wire n_299;
wire n_256;
wire n_172;
wire n_251;
wire n_218;
wire n_271;
wire n_302;
wire n_270;
wire n_153;
wire n_259;
wire n_308;
wire n_140;
wire n_207;
wire n_224;
wire n_219;
wire n_133;
wire n_149;
wire n_214;
wire n_204;
wire n_107;
wire n_254;
wire n_262;
wire n_239;
wire n_276;
wire n_285;
wire n_195;
wire n_165;
wire n_217;
wire n_139;
wire n_193;
wire n_273;
wire n_120;
wire n_245;
wire n_260;
wire n_201;
wire n_197;
wire n_111;
wire n_265;
wire n_264;
wire n_200;
wire n_208;
wire n_126;
wire n_178;
wire n_118;
wire n_179;
wire n_143;
wire n_295;
wire n_263;
wire n_166;
wire n_186;
wire n_136;
wire n_283;
wire n_216;
wire n_147;
wire n_148;
wire n_212;
wire n_168;
wire n_134;
wire n_233;
wire n_106;
wire n_173;
wire n_225;
wire n_220;
wire n_267;
wire n_221;
wire n_203;
wire n_115;
wire n_300;
wire n_158;
wire n_121;
wire n_240;
wire n_180;
wire n_104;
wire n_272;
wire n_146;
wire n_306;
wire n_215;
wire n_242;
wire n_155;
wire n_198;
wire n_169;
wire n_156;
wire n_124;
wire n_297;
wire n_128;
wire n_129;
wire n_188;
wire n_127;
wire n_291;
wire n_170;
wire n_281;
wire n_122;
wire n_187;
wire n_138;
wire n_258;
wire n_253;
wire n_266;
wire n_213;
wire n_182;
wire n_226;
wire n_159;
wire n_176;
wire n_123;
wire n_223;
wire n_194;
wire n_287;
wire n_110;
wire n_261;
wire n_164;
wire n_175;
wire n_145;
wire n_290;
wire n_280;
wire n_132;
wire n_109;
wire n_151;
wire n_257;
wire n_269;
INVxp67_ASAP7_75t_L g104 ( .A(n_91), .Y(n_104) );
CKINVDCx20_ASAP7_75t_R g105 ( .A(n_90), .Y(n_105) );
INVx2_ASAP7_75t_L g106 ( .A(n_73), .Y(n_106) );
CKINVDCx5p33_ASAP7_75t_R g107 ( .A(n_67), .Y(n_107) );
INVx1_ASAP7_75t_L g108 ( .A(n_34), .Y(n_108) );
HB1xp67_ASAP7_75t_L g109 ( .A(n_97), .Y(n_109) );
INVx1_ASAP7_75t_L g110 ( .A(n_32), .Y(n_110) );
INVx3_ASAP7_75t_L g111 ( .A(n_72), .Y(n_111) );
BUFx6f_ASAP7_75t_L g112 ( .A(n_39), .Y(n_112) );
INVx1_ASAP7_75t_L g113 ( .A(n_35), .Y(n_113) );
INVx1_ASAP7_75t_L g114 ( .A(n_59), .Y(n_114) );
INVx2_ASAP7_75t_L g115 ( .A(n_30), .Y(n_115) );
NOR2xp33_ASAP7_75t_L g116 ( .A(n_33), .B(n_41), .Y(n_116) );
CKINVDCx5p33_ASAP7_75t_R g117 ( .A(n_49), .Y(n_117) );
BUFx6f_ASAP7_75t_L g118 ( .A(n_84), .Y(n_118) );
CKINVDCx5p33_ASAP7_75t_R g119 ( .A(n_61), .Y(n_119) );
INVx2_ASAP7_75t_SL g120 ( .A(n_54), .Y(n_120) );
CKINVDCx5p33_ASAP7_75t_R g121 ( .A(n_66), .Y(n_121) );
CKINVDCx5p33_ASAP7_75t_R g122 ( .A(n_75), .Y(n_122) );
INVx1_ASAP7_75t_L g123 ( .A(n_55), .Y(n_123) );
INVx1_ASAP7_75t_L g124 ( .A(n_95), .Y(n_124) );
INVx1_ASAP7_75t_L g125 ( .A(n_71), .Y(n_125) );
CKINVDCx20_ASAP7_75t_R g126 ( .A(n_83), .Y(n_126) );
BUFx6f_ASAP7_75t_L g127 ( .A(n_4), .Y(n_127) );
CKINVDCx20_ASAP7_75t_R g128 ( .A(n_68), .Y(n_128) );
BUFx6f_ASAP7_75t_L g129 ( .A(n_93), .Y(n_129) );
BUFx6f_ASAP7_75t_L g130 ( .A(n_102), .Y(n_130) );
INVx1_ASAP7_75t_L g131 ( .A(n_12), .Y(n_131) );
INVx3_ASAP7_75t_L g132 ( .A(n_11), .Y(n_132) );
INVx1_ASAP7_75t_L g133 ( .A(n_18), .Y(n_133) );
INVx2_ASAP7_75t_L g134 ( .A(n_100), .Y(n_134) );
INVx2_ASAP7_75t_L g135 ( .A(n_92), .Y(n_135) );
BUFx2_ASAP7_75t_L g136 ( .A(n_53), .Y(n_136) );
INVx2_ASAP7_75t_L g137 ( .A(n_81), .Y(n_137) );
INVx1_ASAP7_75t_L g138 ( .A(n_10), .Y(n_138) );
BUFx6f_ASAP7_75t_L g139 ( .A(n_26), .Y(n_139) );
INVx1_ASAP7_75t_L g140 ( .A(n_87), .Y(n_140) );
HB1xp67_ASAP7_75t_L g141 ( .A(n_99), .Y(n_141) );
INVx1_ASAP7_75t_L g142 ( .A(n_70), .Y(n_142) );
INVx1_ASAP7_75t_L g143 ( .A(n_56), .Y(n_143) );
CKINVDCx16_ASAP7_75t_R g144 ( .A(n_15), .Y(n_144) );
INVx3_ASAP7_75t_L g145 ( .A(n_103), .Y(n_145) );
INVx1_ASAP7_75t_L g146 ( .A(n_31), .Y(n_146) );
INVx4_ASAP7_75t_R g147 ( .A(n_80), .Y(n_147) );
INVx1_ASAP7_75t_L g148 ( .A(n_42), .Y(n_148) );
INVx1_ASAP7_75t_L g149 ( .A(n_74), .Y(n_149) );
INVxp67_ASAP7_75t_SL g150 ( .A(n_82), .Y(n_150) );
BUFx6f_ASAP7_75t_L g151 ( .A(n_112), .Y(n_151) );
BUFx2_ASAP7_75t_L g152 ( .A(n_109), .Y(n_152) );
OA21x2_ASAP7_75t_L g153 ( .A1(n_108), .A2(n_24), .B(n_23), .Y(n_153) );
BUFx3_ASAP7_75t_L g154 ( .A(n_111), .Y(n_154) );
OAI21x1_ASAP7_75t_L g155 ( .A1(n_111), .A2(n_27), .B(n_25), .Y(n_155) );
OAI21x1_ASAP7_75t_L g156 ( .A1(n_145), .A2(n_29), .B(n_28), .Y(n_156) );
NAND2xp5_ASAP7_75t_L g157 ( .A(n_141), .B(n_0), .Y(n_157) );
INVx5_ASAP7_75t_L g158 ( .A(n_145), .Y(n_158) );
INVx2_ASAP7_75t_L g159 ( .A(n_106), .Y(n_159) );
INVx3_ASAP7_75t_L g160 ( .A(n_132), .Y(n_160) );
INVx2_ASAP7_75t_L g161 ( .A(n_115), .Y(n_161) );
AND2x4_ASAP7_75t_L g162 ( .A(n_132), .B(n_1), .Y(n_162) );
BUFx6f_ASAP7_75t_L g163 ( .A(n_112), .Y(n_163) );
INVx1_ASAP7_75t_L g164 ( .A(n_136), .Y(n_164) );
INVx3_ASAP7_75t_L g165 ( .A(n_127), .Y(n_165) );
BUFx6f_ASAP7_75t_L g166 ( .A(n_112), .Y(n_166) );
NOR2xp33_ASAP7_75t_L g167 ( .A(n_120), .B(n_2), .Y(n_167) );
INVx6_ASAP7_75t_L g168 ( .A(n_112), .Y(n_168) );
BUFx6f_ASAP7_75t_L g169 ( .A(n_118), .Y(n_169) );
INVx2_ASAP7_75t_L g170 ( .A(n_163), .Y(n_170) );
OAI22xp5_ASAP7_75t_L g171 ( .A1(n_152), .A2(n_144), .B1(n_105), .B2(n_128), .Y(n_171) );
INVx2_ASAP7_75t_SL g172 ( .A(n_154), .Y(n_172) );
INVx3_ASAP7_75t_L g173 ( .A(n_162), .Y(n_173) );
INVx2_ASAP7_75t_L g174 ( .A(n_163), .Y(n_174) );
BUFx4f_ASAP7_75t_L g175 ( .A(n_153), .Y(n_175) );
INVx1_ASAP7_75t_L g176 ( .A(n_165), .Y(n_176) );
INVx2_ASAP7_75t_SL g177 ( .A(n_158), .Y(n_177) );
INVx2_ASAP7_75t_L g178 ( .A(n_166), .Y(n_178) );
INVx3_ASAP7_75t_L g179 ( .A(n_160), .Y(n_179) );
INVx2_ASAP7_75t_L g180 ( .A(n_166), .Y(n_180) );
NAND2xp5_ASAP7_75t_SL g181 ( .A(n_164), .B(n_104), .Y(n_181) );
AOI22xp33_ASAP7_75t_L g182 ( .A1(n_157), .A2(n_133), .B1(n_138), .B2(n_131), .Y(n_182) );
INVx2_ASAP7_75t_SL g183 ( .A(n_179), .Y(n_183) );
NOR2xp33_ASAP7_75t_L g184 ( .A(n_181), .B(n_167), .Y(n_184) );
NOR2x1_ASAP7_75t_L g185 ( .A(n_171), .B(n_126), .Y(n_185) );
NAND2xp5_ASAP7_75t_L g186 ( .A(n_172), .B(n_160), .Y(n_186) );
INVx2_ASAP7_75t_L g187 ( .A(n_173), .Y(n_187) );
INVx1_ASAP7_75t_L g188 ( .A(n_176), .Y(n_188) );
NOR2xp33_ASAP7_75t_L g189 ( .A(n_182), .B(n_159), .Y(n_189) );
A2O1A1Ixp33_ASAP7_75t_L g190 ( .A1(n_175), .A2(n_155), .B(n_156), .C(n_161), .Y(n_190) );
NOR2xp33_ASAP7_75t_L g191 ( .A(n_177), .B(n_150), .Y(n_191) );
NAND2xp5_ASAP7_75t_L g192 ( .A(n_170), .B(n_107), .Y(n_192) );
BUFx8_ASAP7_75t_L g193 ( .A(n_174), .Y(n_193) );
NAND2x1p5_ASAP7_75t_L g194 ( .A(n_185), .B(n_155), .Y(n_194) );
AO32x2_ASAP7_75t_L g195 ( .A1(n_190), .A2(n_151), .A3(n_169), .B1(n_166), .B2(n_168), .Y(n_195) );
A2O1A1Ixp33_ASAP7_75t_L g196 ( .A1(n_189), .A2(n_110), .B(n_114), .C(n_113), .Y(n_196) );
A2O1A1Ixp33_ASAP7_75t_L g197 ( .A1(n_184), .A2(n_123), .B(n_125), .C(n_124), .Y(n_197) );
INVx2_ASAP7_75t_L g198 ( .A(n_187), .Y(n_198) );
BUFx12f_ASAP7_75t_L g199 ( .A(n_193), .Y(n_199) );
AO32x1_ASAP7_75t_L g200 ( .A1(n_183), .A2(n_143), .A3(n_146), .B1(n_142), .B2(n_140), .Y(n_200) );
INVx1_ASAP7_75t_L g201 ( .A(n_186), .Y(n_201) );
AOI21xp5_ASAP7_75t_L g202 ( .A1(n_188), .A2(n_149), .B(n_148), .Y(n_202) );
OAI22xp5_ASAP7_75t_L g203 ( .A1(n_191), .A2(n_117), .B1(n_121), .B2(n_119), .Y(n_203) );
NOR3xp33_ASAP7_75t_L g204 ( .A(n_192), .B(n_116), .C(n_122), .Y(n_204) );
AO31x2_ASAP7_75t_L g205 ( .A1(n_196), .A2(n_134), .A3(n_137), .B(n_135), .Y(n_205) );
INVx1_ASAP7_75t_L g206 ( .A(n_201), .Y(n_206) );
INVx3_ASAP7_75t_L g207 ( .A(n_199), .Y(n_207) );
AO31x2_ASAP7_75t_L g208 ( .A1(n_197), .A2(n_116), .A3(n_180), .B(n_178), .Y(n_208) );
OAI21xp5_ASAP7_75t_SL g209 ( .A1(n_194), .A2(n_129), .B(n_118), .Y(n_209) );
INVx1_ASAP7_75t_L g210 ( .A(n_198), .Y(n_210) );
INVx1_ASAP7_75t_L g211 ( .A(n_202), .Y(n_211) );
AOI221x1_ASAP7_75t_L g212 ( .A1(n_204), .A2(n_151), .B1(n_169), .B2(n_130), .C(n_139), .Y(n_212) );
AO32x2_ASAP7_75t_L g213 ( .A1(n_195), .A2(n_168), .A3(n_151), .B1(n_169), .B2(n_147), .Y(n_213) );
NAND2xp5_ASAP7_75t_SL g214 ( .A(n_203), .B(n_139), .Y(n_214) );
OAI22xp5_ASAP7_75t_L g215 ( .A1(n_200), .A2(n_6), .B1(n_3), .B2(n_5), .Y(n_215) );
INVx5_ASAP7_75t_L g216 ( .A(n_199), .Y(n_216) );
OR2x6_ASAP7_75t_L g217 ( .A(n_207), .B(n_7), .Y(n_217) );
INVx1_ASAP7_75t_L g218 ( .A(n_206), .Y(n_218) );
INVx1_ASAP7_75t_L g219 ( .A(n_211), .Y(n_219) );
BUFx5_ASAP7_75t_L g220 ( .A(n_210), .Y(n_220) );
OR3x4_ASAP7_75t_SL g221 ( .A(n_216), .B(n_8), .C(n_9), .Y(n_221) );
AO21x2_ASAP7_75t_L g222 ( .A1(n_209), .A2(n_37), .B(n_36), .Y(n_222) );
OA21x2_ASAP7_75t_L g223 ( .A1(n_212), .A2(n_40), .B(n_38), .Y(n_223) );
INVx2_ASAP7_75t_SL g224 ( .A(n_205), .Y(n_224) );
BUFx2_ASAP7_75t_R g225 ( .A(n_214), .Y(n_225) );
INVx2_ASAP7_75t_L g226 ( .A(n_205), .Y(n_226) );
INVx3_ASAP7_75t_L g227 ( .A(n_205), .Y(n_227) );
OA21x2_ASAP7_75t_L g228 ( .A1(n_213), .A2(n_44), .B(n_43), .Y(n_228) );
INVx1_ASAP7_75t_L g229 ( .A(n_208), .Y(n_229) );
OA21x2_ASAP7_75t_L g230 ( .A1(n_213), .A2(n_46), .B(n_45), .Y(n_230) );
AO31x2_ASAP7_75t_L g231 ( .A1(n_215), .A2(n_12), .A3(n_13), .B(n_14), .Y(n_231) );
OAI21x1_ASAP7_75t_L g232 ( .A1(n_208), .A2(n_48), .B(n_47), .Y(n_232) );
INVx2_ASAP7_75t_L g233 ( .A(n_219), .Y(n_233) );
INVx1_ASAP7_75t_L g234 ( .A(n_218), .Y(n_234) );
INVx2_ASAP7_75t_L g235 ( .A(n_219), .Y(n_235) );
AO21x2_ASAP7_75t_L g236 ( .A1(n_229), .A2(n_16), .B(n_17), .Y(n_236) );
INVx2_ASAP7_75t_L g237 ( .A(n_220), .Y(n_237) );
HB1xp67_ASAP7_75t_L g238 ( .A(n_224), .Y(n_238) );
AND2x2_ASAP7_75t_L g239 ( .A(n_217), .B(n_19), .Y(n_239) );
INVx1_ASAP7_75t_L g240 ( .A(n_231), .Y(n_240) );
INVx2_ASAP7_75t_L g241 ( .A(n_231), .Y(n_241) );
OA21x2_ASAP7_75t_L g242 ( .A1(n_226), .A2(n_51), .B(n_50), .Y(n_242) );
AO21x2_ASAP7_75t_L g243 ( .A1(n_232), .A2(n_20), .B(n_21), .Y(n_243) );
NAND2xp5_ASAP7_75t_L g244 ( .A(n_227), .B(n_22), .Y(n_244) );
INVx2_ASAP7_75t_L g245 ( .A(n_228), .Y(n_245) );
INVx1_ASAP7_75t_SL g246 ( .A(n_225), .Y(n_246) );
BUFx2_ASAP7_75t_L g247 ( .A(n_222), .Y(n_247) );
AND2x2_ASAP7_75t_L g248 ( .A(n_221), .B(n_52), .Y(n_248) );
HB1xp67_ASAP7_75t_L g249 ( .A(n_230), .Y(n_249) );
INVx1_ASAP7_75t_L g250 ( .A(n_223), .Y(n_250) );
AO21x2_ASAP7_75t_L g251 ( .A1(n_250), .A2(n_57), .B(n_58), .Y(n_251) );
INVx1_ASAP7_75t_L g252 ( .A(n_233), .Y(n_252) );
INVx1_ASAP7_75t_L g253 ( .A(n_235), .Y(n_253) );
INVx1_ASAP7_75t_L g254 ( .A(n_240), .Y(n_254) );
INVx1_ASAP7_75t_L g255 ( .A(n_234), .Y(n_255) );
AND2x6_ASAP7_75t_L g256 ( .A(n_237), .B(n_60), .Y(n_256) );
AOI211x1_ASAP7_75t_L g257 ( .A1(n_239), .A2(n_62), .B(n_63), .C(n_64), .Y(n_257) );
INVx2_ASAP7_75t_L g258 ( .A(n_236), .Y(n_258) );
OR2x2_ASAP7_75t_L g259 ( .A(n_246), .B(n_65), .Y(n_259) );
INVx1_ASAP7_75t_L g260 ( .A(n_241), .Y(n_260) );
AND2x2_ASAP7_75t_L g261 ( .A(n_248), .B(n_69), .Y(n_261) );
INVx1_ASAP7_75t_L g262 ( .A(n_244), .Y(n_262) );
INVx1_ASAP7_75t_L g263 ( .A(n_238), .Y(n_263) );
INVx1_ASAP7_75t_L g264 ( .A(n_238), .Y(n_264) );
INVx2_ASAP7_75t_L g265 ( .A(n_243), .Y(n_265) );
INVx1_ASAP7_75t_L g266 ( .A(n_249), .Y(n_266) );
INVx1_ASAP7_75t_L g267 ( .A(n_249), .Y(n_267) );
INVx3_ASAP7_75t_L g268 ( .A(n_242), .Y(n_268) );
OR2x2_ASAP7_75t_L g269 ( .A(n_245), .B(n_101), .Y(n_269) );
AOI22xp33_ASAP7_75t_L g270 ( .A1(n_247), .A2(n_76), .B1(n_77), .B2(n_78), .Y(n_270) );
INVx1_ASAP7_75t_L g271 ( .A(n_255), .Y(n_271) );
INVx1_ASAP7_75t_L g272 ( .A(n_252), .Y(n_272) );
INVx1_ASAP7_75t_L g273 ( .A(n_253), .Y(n_273) );
AND2x4_ASAP7_75t_L g274 ( .A(n_254), .B(n_79), .Y(n_274) );
HB1xp67_ASAP7_75t_L g275 ( .A(n_263), .Y(n_275) );
HB1xp67_ASAP7_75t_L g276 ( .A(n_264), .Y(n_276) );
INVx1_ASAP7_75t_L g277 ( .A(n_262), .Y(n_277) );
INVx2_ASAP7_75t_L g278 ( .A(n_260), .Y(n_278) );
AND2x4_ASAP7_75t_L g279 ( .A(n_266), .B(n_85), .Y(n_279) );
AOI21xp33_ASAP7_75t_SL g280 ( .A1(n_259), .A2(n_86), .B(n_88), .Y(n_280) );
NAND2xp5_ASAP7_75t_L g281 ( .A(n_261), .B(n_89), .Y(n_281) );
INVx2_ASAP7_75t_L g282 ( .A(n_267), .Y(n_282) );
HB1xp67_ASAP7_75t_L g283 ( .A(n_258), .Y(n_283) );
INVx2_ASAP7_75t_L g284 ( .A(n_268), .Y(n_284) );
OR2x2_ASAP7_75t_L g285 ( .A(n_269), .B(n_94), .Y(n_285) );
NAND2xp5_ASAP7_75t_L g286 ( .A(n_277), .B(n_265), .Y(n_286) );
INVx1_ASAP7_75t_L g287 ( .A(n_275), .Y(n_287) );
INVx1_ASAP7_75t_L g288 ( .A(n_276), .Y(n_288) );
INVx1_ASAP7_75t_L g289 ( .A(n_271), .Y(n_289) );
NAND2xp5_ASAP7_75t_L g290 ( .A(n_282), .B(n_257), .Y(n_290) );
NAND2xp5_ASAP7_75t_L g291 ( .A(n_272), .B(n_251), .Y(n_291) );
NAND2xp5_ASAP7_75t_L g292 ( .A(n_273), .B(n_251), .Y(n_292) );
INVx1_ASAP7_75t_L g293 ( .A(n_289), .Y(n_293) );
NAND2xp5_ASAP7_75t_L g294 ( .A(n_287), .B(n_278), .Y(n_294) );
NAND2xp5_ASAP7_75t_L g295 ( .A(n_288), .B(n_278), .Y(n_295) );
O2A1O1Ixp33_ASAP7_75t_L g296 ( .A1(n_293), .A2(n_280), .B(n_290), .C(n_281), .Y(n_296) );
INVxp67_ASAP7_75t_L g297 ( .A(n_296), .Y(n_297) );
NAND3xp33_ASAP7_75t_L g298 ( .A(n_297), .B(n_295), .C(n_294), .Y(n_298) );
INVx2_ASAP7_75t_L g299 ( .A(n_298), .Y(n_299) );
NAND2xp5_ASAP7_75t_SL g300 ( .A(n_299), .B(n_279), .Y(n_300) );
INVx1_ASAP7_75t_L g301 ( .A(n_300), .Y(n_301) );
INVx2_ASAP7_75t_L g302 ( .A(n_301), .Y(n_302) );
INVx2_ASAP7_75t_L g303 ( .A(n_302), .Y(n_303) );
OAI22xp5_ASAP7_75t_L g304 ( .A1(n_303), .A2(n_292), .B1(n_291), .B2(n_286), .Y(n_304) );
OAI22xp5_ASAP7_75t_L g305 ( .A1(n_304), .A2(n_292), .B1(n_291), .B2(n_285), .Y(n_305) );
AOI21xp33_ASAP7_75t_SL g306 ( .A1(n_305), .A2(n_96), .B(n_98), .Y(n_306) );
OAI21xp5_ASAP7_75t_L g307 ( .A1(n_306), .A2(n_256), .B(n_270), .Y(n_307) );
INVx1_ASAP7_75t_L g308 ( .A(n_307), .Y(n_308) );
AOI22xp33_ASAP7_75t_L g309 ( .A1(n_308), .A2(n_284), .B1(n_283), .B2(n_274), .Y(n_309) );
endmodule