module fake_jpeg_24934_n_51 (n_13, n_21, n_1, n_10, n_23, n_6, n_22, n_14, n_19, n_18, n_20, n_4, n_16, n_3, n_0, n_24, n_9, n_5, n_11, n_17, n_25, n_2, n_12, n_8, n_15, n_7, n_51);

input n_13;
input n_21;
input n_1;
input n_10;
input n_23;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_4;
input n_16;
input n_3;
input n_0;
input n_24;
input n_9;
input n_5;
input n_11;
input n_17;
input n_25;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_51;

wire n_33;
wire n_45;
wire n_27;
wire n_47;
wire n_40;
wire n_35;
wire n_48;
wire n_46;
wire n_41;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_49;
wire n_28;
wire n_38;
wire n_26;
wire n_44;
wire n_36;
wire n_31;
wire n_29;
wire n_37;
wire n_43;
wire n_50;
wire n_32;

INVx4_ASAP7_75t_L g26 ( 
.A(n_13),
.Y(n_26)
);

NOR2xp33_ASAP7_75t_L g27 ( 
.A(n_14),
.B(n_16),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_8),
.Y(n_28)
);

INVx2_ASAP7_75t_L g29 ( 
.A(n_24),
.Y(n_29)
);

INVx3_ASAP7_75t_SL g30 ( 
.A(n_15),
.Y(n_30)
);

NAND2xp5_ASAP7_75t_L g31 ( 
.A(n_20),
.B(n_9),
.Y(n_31)
);

OAI21xp33_ASAP7_75t_L g32 ( 
.A1(n_31),
.A2(n_11),
.B(n_23),
.Y(n_32)
);

AO21x1_ASAP7_75t_L g40 ( 
.A1(n_32),
.A2(n_12),
.B(n_18),
.Y(n_40)
);

OAI32xp33_ASAP7_75t_L g33 ( 
.A1(n_27),
.A2(n_10),
.A3(n_22),
.B1(n_21),
.B2(n_3),
.Y(n_33)
);

AOI22xp5_ASAP7_75t_SL g39 ( 
.A1(n_33),
.A2(n_7),
.B1(n_19),
.B2(n_4),
.Y(n_39)
);

INVx2_ASAP7_75t_L g34 ( 
.A(n_28),
.Y(n_34)
);

NAND2xp5_ASAP7_75t_SL g36 ( 
.A(n_34),
.B(n_0),
.Y(n_36)
);

AOI22xp5_ASAP7_75t_L g35 ( 
.A1(n_32),
.A2(n_30),
.B1(n_26),
.B2(n_29),
.Y(n_35)
);

OAI22xp5_ASAP7_75t_SL g41 ( 
.A1(n_35),
.A2(n_1),
.B1(n_2),
.B2(n_5),
.Y(n_41)
);

NAND2xp5_ASAP7_75t_L g42 ( 
.A(n_36),
.B(n_39),
.Y(n_42)
);

MAJIxp5_ASAP7_75t_L g37 ( 
.A(n_34),
.B(n_30),
.C(n_26),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g43 ( 
.A(n_37),
.B(n_38),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_SL g38 ( 
.A(n_32),
.B(n_0),
.Y(n_38)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_40),
.Y(n_44)
);

MAJIxp5_ASAP7_75t_L g45 ( 
.A(n_41),
.B(n_36),
.C(n_40),
.Y(n_45)
);

OAI21xp33_ASAP7_75t_L g47 ( 
.A1(n_45),
.A2(n_46),
.B(n_42),
.Y(n_47)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_43),
.Y(n_46)
);

CKINVDCx16_ASAP7_75t_R g48 ( 
.A(n_47),
.Y(n_48)
);

OAI21xp5_ASAP7_75t_L g49 ( 
.A1(n_48),
.A2(n_44),
.B(n_41),
.Y(n_49)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_49),
.Y(n_50)
);

AOI221xp5_ASAP7_75t_L g51 ( 
.A1(n_50),
.A2(n_6),
.B1(n_17),
.B2(n_25),
.C(n_2),
.Y(n_51)
);


endmodule