module fake_netlist_6_945_n_2346 (n_52, n_435, n_1, n_91, n_326, n_256, n_440, n_507, n_209, n_367, n_465, n_63, n_223, n_278, n_341, n_362, n_148, n_226, n_161, n_22, n_208, n_462, n_68, n_316, n_419, n_28, n_304, n_212, n_50, n_7, n_144, n_365, n_125, n_168, n_384, n_297, n_524, n_342, n_77, n_106, n_358, n_160, n_449, n_131, n_188, n_310, n_509, n_186, n_245, n_0, n_368, n_396, n_495, n_350, n_78, n_84, n_392, n_442, n_480, n_142, n_143, n_382, n_180, n_62, n_349, n_233, n_255, n_284, n_400, n_140, n_337, n_214, n_485, n_67, n_15, n_443, n_246, n_38, n_471, n_289, n_421, n_424, n_59, n_181, n_182, n_238, n_202, n_320, n_108, n_327, n_369, n_280, n_287, n_353, n_389, n_415, n_65, n_230, n_461, n_141, n_383, n_200, n_447, n_176, n_114, n_86, n_198, n_104, n_222, n_179, n_248, n_300, n_517, n_71, n_74, n_229, n_542, n_305, n_72, n_532, n_173, n_535, n_250, n_372, n_468, n_544, n_111, n_504, n_314, n_378, n_413, n_377, n_35, n_183, n_510, n_79, n_375, n_338, n_522, n_466, n_506, n_56, n_360, n_119, n_235, n_536, n_147, n_191, n_340, n_387, n_452, n_39, n_344, n_73, n_428, n_432, n_101, n_167, n_174, n_127, n_516, n_153, n_525, n_156, n_491, n_145, n_42, n_133, n_96, n_8, n_371, n_189, n_405, n_213, n_538, n_294, n_302, n_499, n_380, n_129, n_197, n_11, n_137, n_17, n_343, n_448, n_20, n_494, n_539, n_493, n_397, n_155, n_109, n_529, n_445, n_425, n_122, n_45, n_454, n_34, n_218, n_70, n_234, n_37, n_486, n_381, n_82, n_27, n_236, n_112, n_172, n_472, n_270, n_239, n_126, n_414, n_97, n_58, n_490, n_290, n_220, n_118, n_224, n_48, n_25, n_93, n_80, n_196, n_402, n_352, n_478, n_9, n_460, n_107, n_6, n_417, n_14, n_446, n_498, n_89, n_374, n_366, n_407, n_450, n_103, n_272, n_526, n_185, n_348, n_69, n_376, n_390, n_473, n_293, n_31, n_334, n_53, n_370, n_44, n_458, n_232, n_16, n_163, n_46, n_330, n_470, n_475, n_298, n_18, n_492, n_281, n_258, n_551, n_154, n_456, n_98, n_260, n_265, n_313, n_451, n_279, n_252, n_228, n_356, n_166, n_184, n_552, n_216, n_455, n_83, n_521, n_363, n_395, n_323, n_393, n_411, n_503, n_152, n_92, n_513, n_321, n_331, n_105, n_227, n_132, n_406, n_483, n_102, n_204, n_482, n_474, n_527, n_261, n_420, n_312, n_394, n_32, n_66, n_130, n_519, n_541, n_512, n_164, n_292, n_100, n_121, n_307, n_469, n_433, n_500, n_23, n_476, n_2, n_291, n_219, n_543, n_357, n_150, n_264, n_263, n_481, n_325, n_329, n_464, n_33, n_477, n_549, n_533, n_408, n_61, n_237, n_244, n_399, n_76, n_243, n_124, n_548, n_94, n_282, n_436, n_116, n_211, n_523, n_117, n_175, n_322, n_345, n_409, n_231, n_354, n_40, n_505, n_240, n_139, n_319, n_41, n_134, n_547, n_537, n_273, n_95, n_311, n_10, n_403, n_253, n_123, n_136, n_546, n_249, n_201, n_386, n_159, n_157, n_162, n_115, n_487, n_550, n_128, n_241, n_30, n_275, n_553, n_43, n_276, n_441, n_221, n_444, n_423, n_146, n_318, n_303, n_511, n_467, n_306, n_21, n_193, n_269, n_359, n_346, n_88, n_3, n_416, n_530, n_277, n_520, n_418, n_113, n_4, n_199, n_138, n_266, n_296, n_268, n_271, n_404, n_439, n_158, n_217, n_49, n_210, n_299, n_518, n_206, n_5, n_453, n_333, n_215, n_178, n_247, n_225, n_308, n_309, n_355, n_426, n_317, n_149, n_431, n_90, n_347, n_24, n_459, n_54, n_502, n_328, n_534, n_488, n_429, n_373, n_87, n_195, n_285, n_497, n_85, n_99, n_257, n_13, n_203, n_286, n_254, n_207, n_242, n_19, n_47, n_29, n_75, n_401, n_324, n_335, n_430, n_463, n_545, n_489, n_205, n_120, n_251, n_301, n_274, n_110, n_151, n_412, n_81, n_36, n_26, n_55, n_267, n_438, n_339, n_315, n_434, n_515, n_64, n_288, n_427, n_479, n_496, n_422, n_135, n_165, n_351, n_437, n_259, n_177, n_540, n_514, n_528, n_391, n_457, n_364, n_295, n_385, n_388, n_190, n_262, n_484, n_187, n_501, n_531, n_60, n_361, n_508, n_379, n_170, n_332, n_336, n_12, n_398, n_410, n_554, n_194, n_171, n_192, n_57, n_169, n_51, n_283, n_2346);

input n_52;
input n_435;
input n_1;
input n_91;
input n_326;
input n_256;
input n_440;
input n_507;
input n_209;
input n_367;
input n_465;
input n_63;
input n_223;
input n_278;
input n_341;
input n_362;
input n_148;
input n_226;
input n_161;
input n_22;
input n_208;
input n_462;
input n_68;
input n_316;
input n_419;
input n_28;
input n_304;
input n_212;
input n_50;
input n_7;
input n_144;
input n_365;
input n_125;
input n_168;
input n_384;
input n_297;
input n_524;
input n_342;
input n_77;
input n_106;
input n_358;
input n_160;
input n_449;
input n_131;
input n_188;
input n_310;
input n_509;
input n_186;
input n_245;
input n_0;
input n_368;
input n_396;
input n_495;
input n_350;
input n_78;
input n_84;
input n_392;
input n_442;
input n_480;
input n_142;
input n_143;
input n_382;
input n_180;
input n_62;
input n_349;
input n_233;
input n_255;
input n_284;
input n_400;
input n_140;
input n_337;
input n_214;
input n_485;
input n_67;
input n_15;
input n_443;
input n_246;
input n_38;
input n_471;
input n_289;
input n_421;
input n_424;
input n_59;
input n_181;
input n_182;
input n_238;
input n_202;
input n_320;
input n_108;
input n_327;
input n_369;
input n_280;
input n_287;
input n_353;
input n_389;
input n_415;
input n_65;
input n_230;
input n_461;
input n_141;
input n_383;
input n_200;
input n_447;
input n_176;
input n_114;
input n_86;
input n_198;
input n_104;
input n_222;
input n_179;
input n_248;
input n_300;
input n_517;
input n_71;
input n_74;
input n_229;
input n_542;
input n_305;
input n_72;
input n_532;
input n_173;
input n_535;
input n_250;
input n_372;
input n_468;
input n_544;
input n_111;
input n_504;
input n_314;
input n_378;
input n_413;
input n_377;
input n_35;
input n_183;
input n_510;
input n_79;
input n_375;
input n_338;
input n_522;
input n_466;
input n_506;
input n_56;
input n_360;
input n_119;
input n_235;
input n_536;
input n_147;
input n_191;
input n_340;
input n_387;
input n_452;
input n_39;
input n_344;
input n_73;
input n_428;
input n_432;
input n_101;
input n_167;
input n_174;
input n_127;
input n_516;
input n_153;
input n_525;
input n_156;
input n_491;
input n_145;
input n_42;
input n_133;
input n_96;
input n_8;
input n_371;
input n_189;
input n_405;
input n_213;
input n_538;
input n_294;
input n_302;
input n_499;
input n_380;
input n_129;
input n_197;
input n_11;
input n_137;
input n_17;
input n_343;
input n_448;
input n_20;
input n_494;
input n_539;
input n_493;
input n_397;
input n_155;
input n_109;
input n_529;
input n_445;
input n_425;
input n_122;
input n_45;
input n_454;
input n_34;
input n_218;
input n_70;
input n_234;
input n_37;
input n_486;
input n_381;
input n_82;
input n_27;
input n_236;
input n_112;
input n_172;
input n_472;
input n_270;
input n_239;
input n_126;
input n_414;
input n_97;
input n_58;
input n_490;
input n_290;
input n_220;
input n_118;
input n_224;
input n_48;
input n_25;
input n_93;
input n_80;
input n_196;
input n_402;
input n_352;
input n_478;
input n_9;
input n_460;
input n_107;
input n_6;
input n_417;
input n_14;
input n_446;
input n_498;
input n_89;
input n_374;
input n_366;
input n_407;
input n_450;
input n_103;
input n_272;
input n_526;
input n_185;
input n_348;
input n_69;
input n_376;
input n_390;
input n_473;
input n_293;
input n_31;
input n_334;
input n_53;
input n_370;
input n_44;
input n_458;
input n_232;
input n_16;
input n_163;
input n_46;
input n_330;
input n_470;
input n_475;
input n_298;
input n_18;
input n_492;
input n_281;
input n_258;
input n_551;
input n_154;
input n_456;
input n_98;
input n_260;
input n_265;
input n_313;
input n_451;
input n_279;
input n_252;
input n_228;
input n_356;
input n_166;
input n_184;
input n_552;
input n_216;
input n_455;
input n_83;
input n_521;
input n_363;
input n_395;
input n_323;
input n_393;
input n_411;
input n_503;
input n_152;
input n_92;
input n_513;
input n_321;
input n_331;
input n_105;
input n_227;
input n_132;
input n_406;
input n_483;
input n_102;
input n_204;
input n_482;
input n_474;
input n_527;
input n_261;
input n_420;
input n_312;
input n_394;
input n_32;
input n_66;
input n_130;
input n_519;
input n_541;
input n_512;
input n_164;
input n_292;
input n_100;
input n_121;
input n_307;
input n_469;
input n_433;
input n_500;
input n_23;
input n_476;
input n_2;
input n_291;
input n_219;
input n_543;
input n_357;
input n_150;
input n_264;
input n_263;
input n_481;
input n_325;
input n_329;
input n_464;
input n_33;
input n_477;
input n_549;
input n_533;
input n_408;
input n_61;
input n_237;
input n_244;
input n_399;
input n_76;
input n_243;
input n_124;
input n_548;
input n_94;
input n_282;
input n_436;
input n_116;
input n_211;
input n_523;
input n_117;
input n_175;
input n_322;
input n_345;
input n_409;
input n_231;
input n_354;
input n_40;
input n_505;
input n_240;
input n_139;
input n_319;
input n_41;
input n_134;
input n_547;
input n_537;
input n_273;
input n_95;
input n_311;
input n_10;
input n_403;
input n_253;
input n_123;
input n_136;
input n_546;
input n_249;
input n_201;
input n_386;
input n_159;
input n_157;
input n_162;
input n_115;
input n_487;
input n_550;
input n_128;
input n_241;
input n_30;
input n_275;
input n_553;
input n_43;
input n_276;
input n_441;
input n_221;
input n_444;
input n_423;
input n_146;
input n_318;
input n_303;
input n_511;
input n_467;
input n_306;
input n_21;
input n_193;
input n_269;
input n_359;
input n_346;
input n_88;
input n_3;
input n_416;
input n_530;
input n_277;
input n_520;
input n_418;
input n_113;
input n_4;
input n_199;
input n_138;
input n_266;
input n_296;
input n_268;
input n_271;
input n_404;
input n_439;
input n_158;
input n_217;
input n_49;
input n_210;
input n_299;
input n_518;
input n_206;
input n_5;
input n_453;
input n_333;
input n_215;
input n_178;
input n_247;
input n_225;
input n_308;
input n_309;
input n_355;
input n_426;
input n_317;
input n_149;
input n_431;
input n_90;
input n_347;
input n_24;
input n_459;
input n_54;
input n_502;
input n_328;
input n_534;
input n_488;
input n_429;
input n_373;
input n_87;
input n_195;
input n_285;
input n_497;
input n_85;
input n_99;
input n_257;
input n_13;
input n_203;
input n_286;
input n_254;
input n_207;
input n_242;
input n_19;
input n_47;
input n_29;
input n_75;
input n_401;
input n_324;
input n_335;
input n_430;
input n_463;
input n_545;
input n_489;
input n_205;
input n_120;
input n_251;
input n_301;
input n_274;
input n_110;
input n_151;
input n_412;
input n_81;
input n_36;
input n_26;
input n_55;
input n_267;
input n_438;
input n_339;
input n_315;
input n_434;
input n_515;
input n_64;
input n_288;
input n_427;
input n_479;
input n_496;
input n_422;
input n_135;
input n_165;
input n_351;
input n_437;
input n_259;
input n_177;
input n_540;
input n_514;
input n_528;
input n_391;
input n_457;
input n_364;
input n_295;
input n_385;
input n_388;
input n_190;
input n_262;
input n_484;
input n_187;
input n_501;
input n_531;
input n_60;
input n_361;
input n_508;
input n_379;
input n_170;
input n_332;
input n_336;
input n_12;
input n_398;
input n_410;
input n_554;
input n_194;
input n_171;
input n_192;
input n_57;
input n_169;
input n_51;
input n_283;

output n_2346;

wire n_992;
wire n_1671;
wire n_801;
wire n_1613;
wire n_1234;
wire n_1458;
wire n_1199;
wire n_1674;
wire n_741;
wire n_1027;
wire n_1351;
wire n_625;
wire n_1189;
wire n_1212;
wire n_726;
wire n_2157;
wire n_2332;
wire n_700;
wire n_1307;
wire n_2003;
wire n_1038;
wire n_578;
wire n_1581;
wire n_1003;
wire n_1237;
wire n_1061;
wire n_1357;
wire n_1853;
wire n_783;
wire n_1738;
wire n_2243;
wire n_798;
wire n_1575;
wire n_1854;
wire n_2324;
wire n_1923;
wire n_1342;
wire n_1209;
wire n_1348;
wire n_1387;
wire n_2260;
wire n_677;
wire n_1708;
wire n_805;
wire n_1151;
wire n_1739;
wire n_2051;
wire n_2317;
wire n_1380;
wire n_1402;
wire n_1688;
wire n_1691;
wire n_1975;
wire n_1009;
wire n_1743;
wire n_1930;
wire n_1160;
wire n_883;
wire n_1238;
wire n_1991;
wire n_2179;
wire n_1724;
wire n_1032;
wire n_2336;
wire n_1247;
wire n_1547;
wire n_1553;
wire n_893;
wire n_1099;
wire n_1264;
wire n_1192;
wire n_1844;
wire n_1700;
wire n_1555;
wire n_1415;
wire n_2211;
wire n_1370;
wire n_1786;
wire n_2291;
wire n_830;
wire n_2299;
wire n_873;
wire n_1371;
wire n_1285;
wire n_1985;
wire n_2184;
wire n_1803;
wire n_1172;
wire n_852;
wire n_1590;
wire n_1532;
wire n_2313;
wire n_1393;
wire n_1517;
wire n_1867;
wire n_1704;
wire n_1078;
wire n_1711;
wire n_2247;
wire n_1140;
wire n_1444;
wire n_1670;
wire n_1603;
wire n_2344;
wire n_1579;
wire n_2321;
wire n_1263;
wire n_2019;
wire n_836;
wire n_2074;
wire n_2129;
wire n_2340;
wire n_1261;
wire n_945;
wire n_2286;
wire n_1649;
wire n_2018;
wire n_2094;
wire n_1903;
wire n_1511;
wire n_1143;
wire n_1422;
wire n_1232;
wire n_1772;
wire n_1572;
wire n_616;
wire n_658;
wire n_1874;
wire n_1119;
wire n_2013;
wire n_1433;
wire n_1902;
wire n_1842;
wire n_1620;
wire n_2044;
wire n_1954;
wire n_1735;
wire n_1541;
wire n_1300;
wire n_641;
wire n_822;
wire n_693;
wire n_1313;
wire n_1056;
wire n_2212;
wire n_758;
wire n_1455;
wire n_1163;
wire n_1180;
wire n_2256;
wire n_943;
wire n_1798;
wire n_1550;
wire n_1591;
wire n_772;
wire n_1344;
wire n_666;
wire n_940;
wire n_770;
wire n_567;
wire n_1781;
wire n_1971;
wire n_2058;
wire n_2090;
wire n_2173;
wire n_2004;
wire n_1106;
wire n_886;
wire n_1471;
wire n_953;
wire n_1094;
wire n_1345;
wire n_1820;
wire n_2108;
wire n_1421;
wire n_1936;
wire n_638;
wire n_1404;
wire n_1211;
wire n_2124;
wire n_887;
wire n_1660;
wire n_1961;
wire n_1280;
wire n_713;
wire n_1400;
wire n_1467;
wire n_976;
wire n_2155;
wire n_1445;
wire n_1560;
wire n_1526;
wire n_734;
wire n_1088;
wire n_1894;
wire n_1231;
wire n_1978;
wire n_2085;
wire n_917;
wire n_574;
wire n_907;
wire n_1446;
wire n_659;
wire n_1815;
wire n_2214;
wire n_913;
wire n_1658;
wire n_808;
wire n_867;
wire n_1230;
wire n_1193;
wire n_1967;
wire n_1054;
wire n_559;
wire n_1333;
wire n_1648;
wire n_1911;
wire n_1956;
wire n_1644;
wire n_2011;
wire n_2277;
wire n_1558;
wire n_1732;
wire n_699;
wire n_1986;
wire n_2300;
wire n_564;
wire n_824;
wire n_686;
wire n_757;
wire n_594;
wire n_1641;
wire n_2113;
wire n_1918;
wire n_2190;
wire n_577;
wire n_1843;
wire n_619;
wire n_2268;
wire n_1367;
wire n_1336;
wire n_572;
wire n_813;
wire n_1909;
wire n_2080;
wire n_1481;
wire n_606;
wire n_1441;
wire n_818;
wire n_1123;
wire n_1309;
wire n_2104;
wire n_645;
wire n_1381;
wire n_1699;
wire n_916;
wire n_2093;
wire n_2207;
wire n_1970;
wire n_608;
wire n_2101;
wire n_630;
wire n_2059;
wire n_2198;
wire n_2073;
wire n_2273;
wire n_792;
wire n_1328;
wire n_1957;
wire n_1907;
wire n_1162;
wire n_860;
wire n_1530;
wire n_788;
wire n_939;
wire n_1543;
wire n_821;
wire n_938;
wire n_1302;
wire n_1068;
wire n_1599;
wire n_982;
wire n_1762;
wire n_1910;
wire n_1075;
wire n_932;
wire n_1876;
wire n_1895;
wire n_2123;
wire n_1697;
wire n_2143;
wire n_979;
wire n_1873;
wire n_905;
wire n_1866;
wire n_1680;
wire n_993;
wire n_689;
wire n_2031;
wire n_2130;
wire n_1330;
wire n_1413;
wire n_1605;
wire n_2228;
wire n_1988;
wire n_1278;
wire n_558;
wire n_1064;
wire n_1396;
wire n_634;
wire n_966;
wire n_764;
wire n_1663;
wire n_2009;
wire n_692;
wire n_733;
wire n_1793;
wire n_1233;
wire n_1289;
wire n_2245;
wire n_2068;
wire n_1107;
wire n_1014;
wire n_1290;
wire n_1703;
wire n_882;
wire n_2176;
wire n_2072;
wire n_1354;
wire n_586;
wire n_1865;
wire n_1875;
wire n_1701;
wire n_1111;
wire n_1713;
wire n_715;
wire n_1251;
wire n_1265;
wire n_1726;
wire n_1950;
wire n_1563;
wire n_1912;
wire n_1982;
wire n_618;
wire n_1297;
wire n_1662;
wire n_1312;
wire n_1167;
wire n_1359;
wire n_674;
wire n_871;
wire n_922;
wire n_1335;
wire n_1760;
wire n_1927;
wire n_2028;
wire n_1069;
wire n_1664;
wire n_1722;
wire n_612;
wire n_1165;
wire n_702;
wire n_2008;
wire n_2192;
wire n_2254;
wire n_2345;
wire n_1926;
wire n_1175;
wire n_1386;
wire n_2311;
wire n_1896;
wire n_1747;
wire n_1012;
wire n_780;
wire n_675;
wire n_903;
wire n_1540;
wire n_1977;
wire n_1802;
wire n_1504;
wire n_2193;
wire n_1655;
wire n_835;
wire n_928;
wire n_1214;
wire n_1801;
wire n_850;
wire n_690;
wire n_1886;
wire n_2092;
wire n_1654;
wire n_816;
wire n_1157;
wire n_1750;
wire n_1462;
wire n_1188;
wire n_1752;
wire n_877;
wire n_1813;
wire n_2206;
wire n_604;
wire n_2319;
wire n_825;
wire n_728;
wire n_1063;
wire n_1588;
wire n_1124;
wire n_1624;
wire n_2096;
wire n_1965;
wire n_598;
wire n_696;
wire n_1515;
wire n_961;
wire n_1082;
wire n_1317;
wire n_593;
wire n_697;
wire n_687;
wire n_890;
wire n_637;
wire n_701;
wire n_2178;
wire n_950;
wire n_2036;
wire n_2152;
wire n_1709;
wire n_1825;
wire n_1796;
wire n_1757;
wire n_1792;
wire n_891;
wire n_2067;
wire n_2136;
wire n_2082;
wire n_2252;
wire n_1412;
wire n_949;
wire n_1630;
wire n_678;
wire n_2075;
wire n_2194;
wire n_1987;
wire n_968;
wire n_909;
wire n_1369;
wire n_881;
wire n_2271;
wire n_1008;
wire n_760;
wire n_1546;
wire n_590;
wire n_2279;
wire n_1033;
wire n_1052;
wire n_1296;
wire n_1990;
wire n_694;
wire n_2150;
wire n_1294;
wire n_1420;
wire n_1634;
wire n_2078;
wire n_595;
wire n_627;
wire n_1767;
wire n_1779;
wire n_1465;
wire n_1858;
wire n_1044;
wire n_2165;
wire n_2133;
wire n_1712;
wire n_1391;
wire n_1523;
wire n_1208;
wire n_1164;
wire n_1295;
wire n_1627;
wire n_1072;
wire n_1527;
wire n_1495;
wire n_1438;
wire n_815;
wire n_1100;
wire n_585;
wire n_1487;
wire n_840;
wire n_874;
wire n_1756;
wire n_1128;
wire n_673;
wire n_2230;
wire n_1969;
wire n_1071;
wire n_1067;
wire n_1565;
wire n_1493;
wire n_2145;
wire n_1968;
wire n_898;
wire n_1952;
wire n_865;
wire n_925;
wire n_1932;
wire n_1101;
wire n_1026;
wire n_1880;
wire n_1364;
wire n_615;
wire n_1249;
wire n_1293;
wire n_1127;
wire n_1512;
wire n_2151;
wire n_1451;
wire n_639;
wire n_963;
wire n_794;
wire n_727;
wire n_894;
wire n_1839;
wire n_2341;
wire n_685;
wire n_1765;
wire n_605;
wire n_1514;
wire n_1863;
wire n_826;
wire n_1646;
wire n_872;
wire n_1139;
wire n_1714;
wire n_718;
wire n_1018;
wire n_1521;
wire n_1366;
wire n_847;
wire n_851;
wire n_682;
wire n_644;
wire n_996;
wire n_1308;
wire n_2089;
wire n_1376;
wire n_1513;
wire n_791;
wire n_1913;
wire n_837;
wire n_2097;
wire n_2170;
wire n_1488;
wire n_1808;
wire n_948;
wire n_704;
wire n_2148;
wire n_977;
wire n_2339;
wire n_1005;
wire n_1947;
wire n_1788;
wire n_1999;
wire n_622;
wire n_1469;
wire n_2060;
wire n_1838;
wire n_1835;
wire n_1766;
wire n_1776;
wire n_1959;
wire n_2002;
wire n_581;
wire n_2138;
wire n_765;
wire n_987;
wire n_1492;
wire n_1340;
wire n_1771;
wire n_2316;
wire n_631;
wire n_720;
wire n_842;
wire n_2262;
wire n_1707;
wire n_2239;
wire n_1432;
wire n_2208;
wire n_843;
wire n_656;
wire n_989;
wire n_1277;
wire n_797;
wire n_1473;
wire n_2191;
wire n_1723;
wire n_1246;
wire n_1878;
wire n_899;
wire n_738;
wire n_2012;
wire n_1304;
wire n_1035;
wire n_1426;
wire n_705;
wire n_1004;
wire n_1176;
wire n_2134;
wire n_1529;
wire n_2335;
wire n_1022;
wire n_614;
wire n_2069;
wire n_2307;
wire n_684;
wire n_1431;
wire n_1615;
wire n_1474;
wire n_1571;
wire n_1809;
wire n_1577;
wire n_2297;
wire n_1181;
wire n_2119;
wire n_1822;
wire n_947;
wire n_1117;
wire n_1087;
wire n_1448;
wire n_1992;
wire n_648;
wire n_657;
wire n_1049;
wire n_2057;
wire n_2103;
wire n_1666;
wire n_1505;
wire n_803;
wire n_1717;
wire n_926;
wire n_1817;
wire n_927;
wire n_1849;
wire n_919;
wire n_1698;
wire n_2231;
wire n_929;
wire n_1228;
wire n_1568;
wire n_1490;
wire n_777;
wire n_1299;
wire n_1183;
wire n_1436;
wire n_2251;
wire n_1384;
wire n_2238;
wire n_1070;
wire n_998;
wire n_717;
wire n_1665;
wire n_1383;
wire n_1178;
wire n_2127;
wire n_1424;
wire n_2338;
wire n_1073;
wire n_1000;
wire n_796;
wire n_1195;
wire n_2137;
wire n_1626;
wire n_1507;
wire n_1358;
wire n_1811;
wire n_1388;
wire n_912;
wire n_1857;
wire n_1519;
wire n_2144;
wire n_745;
wire n_1284;
wire n_1604;
wire n_2296;
wire n_1142;
wire n_716;
wire n_1475;
wire n_623;
wire n_1048;
wire n_1201;
wire n_1398;
wire n_884;
wire n_1774;
wire n_1395;
wire n_2110;
wire n_2199;
wire n_731;
wire n_1502;
wire n_1659;
wire n_1955;
wire n_755;
wire n_1021;
wire n_931;
wire n_811;
wire n_683;
wire n_1207;
wire n_1791;
wire n_1368;
wire n_1418;
wire n_958;
wire n_1250;
wire n_1137;
wire n_1897;
wire n_2064;
wire n_880;
wire n_2053;
wire n_2259;
wire n_2121;
wire n_889;
wire n_1478;
wire n_589;
wire n_1310;
wire n_819;
wire n_2294;
wire n_1363;
wire n_1334;
wire n_1966;
wire n_1942;
wire n_767;
wire n_1314;
wire n_600;
wire n_964;
wire n_831;
wire n_1837;
wire n_2218;
wire n_954;
wire n_864;
wire n_1110;
wire n_2213;
wire n_1410;
wire n_1440;
wire n_2132;
wire n_2063;
wire n_1382;
wire n_1534;
wire n_1564;
wire n_1736;
wire n_1483;
wire n_1834;
wire n_2331;
wire n_1372;
wire n_2292;
wire n_2330;
wire n_1457;
wire n_1719;
wire n_1339;
wire n_1787;
wire n_1993;
wire n_2281;
wire n_1427;
wire n_1466;
wire n_1919;
wire n_1080;
wire n_723;
wire n_1877;
wire n_596;
wire n_562;
wire n_1141;
wire n_1268;
wire n_1939;
wire n_2030;
wire n_1769;
wire n_1220;
wire n_2323;
wire n_1893;
wire n_556;
wire n_2209;
wire n_2301;
wire n_1755;
wire n_1602;
wire n_1136;
wire n_2025;
wire n_1125;
wire n_970;
wire n_2224;
wire n_1980;
wire n_1159;
wire n_995;
wire n_642;
wire n_2329;
wire n_1092;
wire n_2237;
wire n_1060;
wire n_1951;
wire n_2250;
wire n_1252;
wire n_1784;
wire n_1223;
wire n_1286;
wire n_1773;
wire n_1775;
wire n_2115;
wire n_1053;
wire n_1681;
wire n_1093;
wire n_1783;
wire n_1533;
wire n_1597;
wire n_2274;
wire n_775;
wire n_651;
wire n_1153;
wire n_1618;
wire n_1531;
wire n_1185;
wire n_1745;
wire n_914;
wire n_759;
wire n_1831;
wire n_1653;
wire n_1679;
wire n_1625;
wire n_2160;
wire n_1453;
wire n_2146;
wire n_2226;
wire n_2131;
wire n_773;
wire n_1901;
wire n_920;
wire n_1374;
wire n_1315;
wire n_1647;
wire n_1224;
wire n_2306;
wire n_1614;
wire n_1459;
wire n_1892;
wire n_1933;
wire n_1135;
wire n_1179;
wire n_1169;
wire n_1617;
wire n_1470;
wire n_1243;
wire n_848;
wire n_1096;
wire n_2249;
wire n_1091;
wire n_1917;
wire n_2000;
wire n_1580;
wire n_2227;
wire n_2270;
wire n_1425;
wire n_1881;
wire n_1267;
wire n_1281;
wire n_1806;
wire n_983;
wire n_2023;
wire n_2204;
wire n_1520;
wire n_2159;
wire n_906;
wire n_1390;
wire n_688;
wire n_2289;
wire n_1077;
wire n_1733;
wire n_2315;
wire n_1419;
wire n_1731;
wire n_2158;
wire n_2087;
wire n_1855;
wire n_1636;
wire n_1437;
wire n_2135;
wire n_1645;
wire n_1832;
wire n_1687;
wire n_1439;
wire n_2328;
wire n_1323;
wire n_2202;
wire n_858;
wire n_2049;
wire n_1331;
wire n_736;
wire n_613;
wire n_956;
wire n_960;
wire n_2276;
wire n_663;
wire n_856;
wire n_2100;
wire n_778;
wire n_1668;
wire n_1134;
wire n_1129;
wire n_602;
wire n_1696;
wire n_1995;
wire n_1594;
wire n_2181;
wire n_664;
wire n_1869;
wire n_1764;
wire n_1429;
wire n_1610;
wire n_1889;
wire n_1905;
wire n_2016;
wire n_2343;
wire n_793;
wire n_587;
wire n_1593;
wire n_580;
wire n_762;
wire n_1030;
wire n_1202;
wire n_1937;
wire n_1790;
wire n_1778;
wire n_1635;
wire n_1079;
wire n_1744;
wire n_828;
wire n_2139;
wire n_2142;
wire n_607;
wire n_1551;
wire n_1103;
wire n_2219;
wire n_1203;
wire n_820;
wire n_2327;
wire n_951;
wire n_2201;
wire n_725;
wire n_952;
wire n_999;
wire n_1254;
wire n_575;
wire n_994;
wire n_2263;
wire n_2304;
wire n_1508;
wire n_732;
wire n_974;
wire n_2240;
wire n_2278;
wire n_724;
wire n_1934;
wire n_1020;
wire n_1042;
wire n_628;
wire n_1273;
wire n_1434;
wire n_1573;
wire n_1728;
wire n_557;
wire n_1871;
wire n_617;
wire n_845;
wire n_807;
wire n_1036;
wire n_1138;
wire n_1661;
wire n_1275;
wire n_1549;
wire n_1510;
wire n_892;
wire n_768;
wire n_1468;
wire n_1859;
wire n_2102;
wire n_1095;
wire n_2024;
wire n_1595;
wire n_2156;
wire n_1718;
wire n_1749;
wire n_1683;
wire n_1916;
wire n_597;
wire n_1270;
wire n_1187;
wire n_610;
wire n_1403;
wire n_1669;
wire n_1852;
wire n_1024;
wire n_1768;
wire n_2153;
wire n_2052;
wire n_1847;
wire n_2302;
wire n_1667;
wire n_667;
wire n_1206;
wire n_1037;
wire n_621;
wire n_1397;
wire n_1279;
wire n_1115;
wire n_750;
wire n_901;
wire n_1499;
wire n_923;
wire n_1409;
wire n_1841;
wire n_1639;
wire n_1623;
wire n_1015;
wire n_1503;
wire n_1057;
wire n_603;
wire n_991;
wire n_1657;
wire n_1126;
wire n_1997;
wire n_710;
wire n_1108;
wire n_1818;
wire n_1182;
wire n_1298;
wire n_2177;
wire n_2088;
wire n_1611;
wire n_785;
wire n_746;
wire n_609;
wire n_1601;
wire n_1960;
wire n_2061;
wire n_1686;
wire n_2337;
wire n_1356;
wire n_1589;
wire n_2309;
wire n_1740;
wire n_1497;
wire n_1168;
wire n_1216;
wire n_1943;
wire n_1320;
wire n_1430;
wire n_1316;
wire n_1287;
wire n_1452;
wire n_1622;
wire n_1586;
wire n_2264;
wire n_1694;
wire n_1535;
wire n_1596;
wire n_1190;
wire n_1734;
wire n_1983;
wire n_1938;
wire n_2220;
wire n_1262;
wire n_1891;
wire n_2171;
wire n_1213;
wire n_2235;
wire n_1350;
wire n_1673;
wire n_2232;
wire n_1715;
wire n_1443;
wire n_1272;
wire n_2037;
wire n_2298;
wire n_782;
wire n_2326;
wire n_1539;
wire n_809;
wire n_1043;
wire n_1797;
wire n_1608;
wire n_986;
wire n_2305;
wire n_2120;
wire n_1472;
wire n_2050;
wire n_2164;
wire n_2225;
wire n_1081;
wire n_1870;
wire n_1692;
wire n_800;
wire n_1084;
wire n_1171;
wire n_2169;
wire n_1827;
wire n_1361;
wire n_1864;
wire n_2006;
wire n_1491;
wire n_2187;
wire n_662;
wire n_1152;
wire n_1840;
wire n_1705;
wire n_2244;
wire n_1684;
wire n_921;
wire n_1346;
wire n_711;
wire n_1642;
wire n_579;
wire n_1352;
wire n_937;
wire n_2257;
wire n_1682;
wire n_2017;
wire n_1695;
wire n_1828;
wire n_2046;
wire n_2272;
wire n_2200;
wire n_650;
wire n_1046;
wire n_1940;
wire n_1979;
wire n_1145;
wire n_1121;
wire n_1102;
wire n_1963;
wire n_972;
wire n_1405;
wire n_1406;
wire n_1332;
wire n_624;
wire n_962;
wire n_1041;
wire n_565;
wire n_1569;
wire n_936;
wire n_1883;
wire n_1288;
wire n_1186;
wire n_1062;
wire n_885;
wire n_896;
wire n_2342;
wire n_2167;
wire n_2084;
wire n_654;
wire n_1222;
wire n_599;
wire n_776;
wire n_1823;
wire n_1974;
wire n_1720;
wire n_934;
wire n_1637;
wire n_1407;
wire n_1795;
wire n_1341;
wire n_1456;
wire n_1845;
wire n_1489;
wire n_2314;
wire n_942;
wire n_1524;
wire n_2229;
wire n_1964;
wire n_2288;
wire n_1920;
wire n_2099;
wire n_1496;
wire n_1271;
wire n_1545;
wire n_2007;
wire n_2039;
wire n_1946;
wire n_1355;
wire n_1225;
wire n_1544;
wire n_1485;
wire n_2258;
wire n_1640;
wire n_804;
wire n_1846;
wire n_806;
wire n_959;
wire n_879;
wire n_2310;
wire n_584;
wire n_2141;
wire n_1343;
wire n_1522;
wire n_1782;
wire n_1676;
wire n_833;
wire n_1830;
wire n_1567;
wire n_1319;
wire n_707;
wire n_1900;
wire n_799;
wire n_1548;
wire n_1155;
wire n_2196;
wire n_1633;
wire n_2195;
wire n_787;
wire n_2172;
wire n_1416;
wire n_1528;
wire n_2293;
wire n_1146;
wire n_2021;
wire n_2114;
wire n_1086;
wire n_1066;
wire n_1948;
wire n_2125;
wire n_2026;
wire n_1282;
wire n_2322;
wire n_652;
wire n_2154;
wire n_560;
wire n_1906;
wire n_1484;
wire n_1321;
wire n_1241;
wire n_1672;
wire n_569;
wire n_1758;
wire n_2283;
wire n_1925;
wire n_737;
wire n_1318;
wire n_1914;
wire n_1235;
wire n_1229;
wire n_1292;
wire n_1373;
wire n_2266;
wire n_1029;
wire n_1447;
wire n_2056;
wire n_790;
wire n_1706;
wire n_1498;
wire n_1210;
wire n_1248;
wire n_1556;
wire n_902;
wire n_2189;
wire n_2246;
wire n_1047;
wire n_1984;
wire n_2236;
wire n_1385;
wire n_1269;
wire n_1931;
wire n_2083;
wire n_672;
wire n_1257;
wire n_1751;
wire n_1375;
wire n_1941;
wire n_2128;
wire n_655;
wire n_1045;
wire n_706;
wire n_1650;
wire n_786;
wire n_1794;
wire n_1236;
wire n_1962;
wire n_1559;
wire n_1725;
wire n_1928;
wire n_1872;
wire n_834;
wire n_743;
wire n_766;
wire n_1746;
wire n_1325;
wire n_1002;
wire n_1741;
wire n_1949;
wire n_1804;
wire n_1727;
wire n_1019;
wire n_636;
wire n_2054;
wire n_729;
wire n_876;
wire n_774;
wire n_1337;
wire n_660;
wire n_2062;
wire n_2041;
wire n_1477;
wire n_1360;
wire n_1860;
wire n_1904;
wire n_1200;
wire n_2070;
wire n_1607;
wire n_1353;
wire n_1777;
wire n_1908;
wire n_1454;
wire n_2126;
wire n_869;
wire n_1154;
wire n_1113;
wire n_1600;
wire n_2253;
wire n_646;
wire n_1098;
wire n_1329;
wire n_2045;
wire n_817;
wire n_2261;
wire n_2216;
wire n_2210;
wire n_897;
wire n_846;
wire n_2066;
wire n_841;
wire n_1476;
wire n_1001;
wire n_1800;
wire n_2241;
wire n_1050;
wire n_1411;
wire n_1463;
wire n_1177;
wire n_1150;
wire n_1742;
wire n_1562;
wire n_1690;
wire n_1191;
wire n_1826;
wire n_566;
wire n_1023;
wire n_1882;
wire n_1076;
wire n_1118;
wire n_1007;
wire n_1807;
wire n_1929;
wire n_1378;
wire n_855;
wire n_1592;
wire n_1759;
wire n_1814;
wire n_1631;
wire n_591;
wire n_1377;
wire n_1879;
wire n_853;
wire n_695;
wire n_1542;
wire n_875;
wire n_680;
wire n_1678;
wire n_661;
wire n_1716;
wire n_1256;
wire n_671;
wire n_1953;
wire n_933;
wire n_740;
wire n_703;
wire n_978;
wire n_1976;
wire n_1291;
wire n_1217;
wire n_751;
wire n_749;
wire n_1824;
wire n_1628;
wire n_1324;
wire n_1399;
wire n_2122;
wire n_2109;
wire n_1435;
wire n_969;
wire n_988;
wire n_2140;
wire n_1065;
wire n_1401;
wire n_1255;
wire n_568;
wire n_1516;
wire n_1536;
wire n_2163;
wire n_2186;
wire n_2029;
wire n_1204;
wire n_823;
wire n_1132;
wire n_643;
wire n_1074;
wire n_698;
wire n_1394;
wire n_1327;
wire n_1326;
wire n_955;
wire n_739;
wire n_1379;
wire n_1338;
wire n_1097;
wire n_935;
wire n_781;
wire n_789;
wire n_1554;
wire n_1130;
wire n_1810;
wire n_573;
wire n_769;
wire n_676;
wire n_1120;
wire n_832;
wire n_1583;
wire n_1730;
wire n_2295;
wire n_555;
wire n_814;
wire n_1643;
wire n_2020;
wire n_2269;
wire n_1729;
wire n_669;
wire n_2290;
wire n_2048;
wire n_2005;
wire n_747;
wire n_1389;
wire n_1105;
wire n_721;
wire n_1461;
wire n_742;
wire n_691;
wire n_2076;
wire n_1408;
wire n_1196;
wire n_1598;
wire n_863;
wire n_2175;
wire n_601;
wire n_2182;
wire n_1283;
wire n_918;
wire n_748;
wire n_1114;
wire n_1785;
wire n_1147;
wire n_763;
wire n_1848;
wire n_1754;
wire n_2149;
wire n_1506;
wire n_1652;
wire n_1812;
wire n_957;
wire n_1994;
wire n_895;
wire n_866;
wire n_1227;
wire n_2284;
wire n_2287;
wire n_744;
wire n_971;
wire n_946;
wire n_761;
wire n_1303;
wire n_1205;
wire n_1258;
wire n_1392;
wire n_1173;
wire n_1924;
wire n_1677;
wire n_1116;
wire n_611;
wire n_1570;
wire n_1702;
wire n_1219;
wire n_1780;
wire n_1689;
wire n_2180;
wire n_1174;
wire n_1944;
wire n_1016;
wire n_1347;
wire n_795;
wire n_1501;
wire n_1221;
wire n_1245;
wire n_838;
wire n_647;
wire n_844;
wire n_1017;
wire n_2117;
wire n_2234;
wire n_1083;
wire n_1561;
wire n_930;
wire n_888;
wire n_2275;
wire n_1112;
wire n_2081;
wire n_2168;
wire n_2022;
wire n_1945;
wire n_2203;
wire n_910;
wire n_1656;
wire n_1721;
wire n_1460;
wire n_911;
wire n_2112;
wire n_2255;
wire n_1464;
wire n_653;
wire n_1737;
wire n_1414;
wire n_908;
wire n_752;
wire n_944;
wire n_2034;
wire n_1028;
wire n_576;
wire n_2106;
wire n_2265;
wire n_1922;
wire n_563;
wire n_2032;
wire n_1011;
wire n_1566;
wire n_1215;
wire n_839;
wire n_708;
wire n_1973;
wire n_2267;
wire n_668;
wire n_626;
wire n_990;
wire n_1500;
wire n_779;
wire n_1537;
wire n_1821;
wire n_2205;
wire n_1104;
wire n_1058;
wire n_854;
wire n_2312;
wire n_1122;
wire n_870;
wire n_904;
wire n_1253;
wire n_709;
wire n_1266;
wire n_2242;
wire n_1509;
wire n_1693;
wire n_1109;
wire n_2222;
wire n_712;
wire n_1276;
wire n_2015;
wire n_2118;
wire n_2111;
wire n_1148;
wire n_2188;
wire n_1989;
wire n_1161;
wire n_1085;
wire n_2014;
wire n_2042;
wire n_1239;
wire n_771;
wire n_1584;
wire n_924;
wire n_1582;
wire n_2318;
wire n_1149;
wire n_1184;
wire n_719;
wire n_1972;
wire n_1525;
wire n_1585;
wire n_1851;
wire n_1799;
wire n_1090;
wire n_2147;
wire n_592;
wire n_1816;
wire n_1518;
wire n_829;
wire n_1156;
wire n_1362;
wire n_984;
wire n_1829;
wire n_2035;
wire n_1450;
wire n_1638;
wire n_868;
wire n_570;
wire n_859;
wire n_2033;
wire n_735;
wire n_1789;
wire n_1770;
wire n_878;
wire n_620;
wire n_1218;
wire n_1482;
wire n_981;
wire n_714;
wire n_1349;
wire n_1144;
wire n_2071;
wire n_985;
wire n_2233;
wire n_997;
wire n_1710;
wire n_2161;
wire n_1301;
wire n_802;
wire n_561;
wire n_980;
wire n_1306;
wire n_2010;
wire n_2282;
wire n_1651;
wire n_1198;
wire n_2047;
wire n_2095;
wire n_1609;
wire n_2174;
wire n_2334;
wire n_1244;
wire n_1685;
wire n_1763;
wire n_1998;
wire n_1574;
wire n_756;
wire n_2303;
wire n_1619;
wire n_1981;
wire n_2285;
wire n_1606;
wire n_810;
wire n_1133;
wire n_635;
wire n_1194;
wire n_1051;
wire n_1552;
wire n_583;
wire n_1996;
wire n_1039;
wire n_1442;
wire n_1034;
wire n_2043;
wire n_1480;
wire n_1158;
wire n_2248;
wire n_754;
wire n_941;
wire n_975;
wire n_1031;
wire n_1305;
wire n_849;
wire n_753;
wire n_1753;
wire n_973;
wire n_1921;
wire n_1479;
wire n_1055;
wire n_1675;
wire n_2197;
wire n_2217;
wire n_582;
wire n_2065;
wire n_861;
wire n_857;
wire n_967;
wire n_571;
wire n_2215;
wire n_2001;
wire n_2107;
wire n_1884;
wire n_2040;
wire n_679;
wire n_633;
wire n_1170;
wire n_665;
wire n_1629;
wire n_2221;
wire n_588;
wire n_1260;
wire n_1819;
wire n_2055;
wire n_1010;
wire n_1040;
wire n_915;
wire n_632;
wire n_1166;
wire n_2038;
wire n_812;
wire n_1131;
wire n_1761;
wire n_1578;
wire n_1006;
wire n_1861;
wire n_1632;
wire n_1890;
wire n_1805;
wire n_1888;
wire n_1557;
wire n_2280;
wire n_1833;
wire n_730;
wire n_1311;
wire n_1494;
wire n_2325;
wire n_670;
wire n_1850;
wire n_1898;
wire n_2308;
wire n_2162;
wire n_1868;
wire n_2333;
wire n_2079;
wire n_1089;
wire n_1887;
wire n_1587;
wire n_1365;
wire n_1417;
wire n_1242;
wire n_2086;
wire n_2185;
wire n_1836;
wire n_681;
wire n_1226;
wire n_1274;
wire n_1486;
wire n_2166;
wire n_640;
wire n_1322;
wire n_965;
wire n_1899;
wire n_1428;
wire n_1616;
wire n_1576;
wire n_1862;
wire n_1856;
wire n_1958;
wire n_2077;
wire n_784;
wire n_1059;
wire n_1197;
wire n_722;
wire n_862;
wire n_2105;
wire n_2098;
wire n_1423;
wire n_1935;
wire n_2027;
wire n_2223;
wire n_2091;
wire n_1915;
wire n_629;
wire n_1621;
wire n_1748;
wire n_900;
wire n_1449;
wire n_827;
wire n_1025;
wire n_2116;
wire n_2320;
wire n_1885;
wire n_1013;
wire n_1259;
wire n_2183;
wire n_1538;
wire n_649;
wire n_1612;
wire n_1240;

INVx1_ASAP7_75t_SL g555 ( 
.A(n_392),
.Y(n_555)
);

CKINVDCx5p33_ASAP7_75t_R g556 ( 
.A(n_491),
.Y(n_556)
);

BUFx5_ASAP7_75t_L g557 ( 
.A(n_165),
.Y(n_557)
);

CKINVDCx5p33_ASAP7_75t_R g558 ( 
.A(n_203),
.Y(n_558)
);

INVx1_ASAP7_75t_L g559 ( 
.A(n_335),
.Y(n_559)
);

CKINVDCx5p33_ASAP7_75t_R g560 ( 
.A(n_409),
.Y(n_560)
);

CKINVDCx5p33_ASAP7_75t_R g561 ( 
.A(n_388),
.Y(n_561)
);

INVx1_ASAP7_75t_L g562 ( 
.A(n_261),
.Y(n_562)
);

CKINVDCx5p33_ASAP7_75t_R g563 ( 
.A(n_267),
.Y(n_563)
);

CKINVDCx5p33_ASAP7_75t_R g564 ( 
.A(n_291),
.Y(n_564)
);

CKINVDCx5p33_ASAP7_75t_R g565 ( 
.A(n_278),
.Y(n_565)
);

CKINVDCx5p33_ASAP7_75t_R g566 ( 
.A(n_432),
.Y(n_566)
);

CKINVDCx5p33_ASAP7_75t_R g567 ( 
.A(n_532),
.Y(n_567)
);

CKINVDCx20_ASAP7_75t_R g568 ( 
.A(n_49),
.Y(n_568)
);

CKINVDCx5p33_ASAP7_75t_R g569 ( 
.A(n_449),
.Y(n_569)
);

INVx1_ASAP7_75t_L g570 ( 
.A(n_351),
.Y(n_570)
);

CKINVDCx5p33_ASAP7_75t_R g571 ( 
.A(n_322),
.Y(n_571)
);

CKINVDCx5p33_ASAP7_75t_R g572 ( 
.A(n_273),
.Y(n_572)
);

CKINVDCx5p33_ASAP7_75t_R g573 ( 
.A(n_55),
.Y(n_573)
);

INVx2_ASAP7_75t_SL g574 ( 
.A(n_540),
.Y(n_574)
);

INVx1_ASAP7_75t_SL g575 ( 
.A(n_208),
.Y(n_575)
);

CKINVDCx5p33_ASAP7_75t_R g576 ( 
.A(n_412),
.Y(n_576)
);

INVx1_ASAP7_75t_L g577 ( 
.A(n_157),
.Y(n_577)
);

INVx1_ASAP7_75t_SL g578 ( 
.A(n_179),
.Y(n_578)
);

CKINVDCx5p33_ASAP7_75t_R g579 ( 
.A(n_51),
.Y(n_579)
);

INVx1_ASAP7_75t_SL g580 ( 
.A(n_293),
.Y(n_580)
);

CKINVDCx20_ASAP7_75t_R g581 ( 
.A(n_210),
.Y(n_581)
);

CKINVDCx20_ASAP7_75t_R g582 ( 
.A(n_519),
.Y(n_582)
);

CKINVDCx5p33_ASAP7_75t_R g583 ( 
.A(n_144),
.Y(n_583)
);

CKINVDCx20_ASAP7_75t_R g584 ( 
.A(n_44),
.Y(n_584)
);

BUFx8_ASAP7_75t_SL g585 ( 
.A(n_165),
.Y(n_585)
);

CKINVDCx5p33_ASAP7_75t_R g586 ( 
.A(n_475),
.Y(n_586)
);

CKINVDCx5p33_ASAP7_75t_R g587 ( 
.A(n_50),
.Y(n_587)
);

CKINVDCx5p33_ASAP7_75t_R g588 ( 
.A(n_92),
.Y(n_588)
);

INVx1_ASAP7_75t_L g589 ( 
.A(n_468),
.Y(n_589)
);

INVx1_ASAP7_75t_SL g590 ( 
.A(n_292),
.Y(n_590)
);

CKINVDCx5p33_ASAP7_75t_R g591 ( 
.A(n_450),
.Y(n_591)
);

CKINVDCx5p33_ASAP7_75t_R g592 ( 
.A(n_477),
.Y(n_592)
);

CKINVDCx5p33_ASAP7_75t_R g593 ( 
.A(n_533),
.Y(n_593)
);

BUFx3_ASAP7_75t_L g594 ( 
.A(n_90),
.Y(n_594)
);

INVx2_ASAP7_75t_L g595 ( 
.A(n_365),
.Y(n_595)
);

CKINVDCx5p33_ASAP7_75t_R g596 ( 
.A(n_219),
.Y(n_596)
);

CKINVDCx5p33_ASAP7_75t_R g597 ( 
.A(n_265),
.Y(n_597)
);

CKINVDCx5p33_ASAP7_75t_R g598 ( 
.A(n_536),
.Y(n_598)
);

CKINVDCx5p33_ASAP7_75t_R g599 ( 
.A(n_467),
.Y(n_599)
);

CKINVDCx5p33_ASAP7_75t_R g600 ( 
.A(n_83),
.Y(n_600)
);

CKINVDCx5p33_ASAP7_75t_R g601 ( 
.A(n_124),
.Y(n_601)
);

CKINVDCx5p33_ASAP7_75t_R g602 ( 
.A(n_359),
.Y(n_602)
);

CKINVDCx5p33_ASAP7_75t_R g603 ( 
.A(n_405),
.Y(n_603)
);

CKINVDCx5p33_ASAP7_75t_R g604 ( 
.A(n_430),
.Y(n_604)
);

INVx1_ASAP7_75t_L g605 ( 
.A(n_129),
.Y(n_605)
);

INVx1_ASAP7_75t_L g606 ( 
.A(n_462),
.Y(n_606)
);

CKINVDCx5p33_ASAP7_75t_R g607 ( 
.A(n_59),
.Y(n_607)
);

CKINVDCx5p33_ASAP7_75t_R g608 ( 
.A(n_400),
.Y(n_608)
);

INVx1_ASAP7_75t_L g609 ( 
.A(n_184),
.Y(n_609)
);

INVx1_ASAP7_75t_L g610 ( 
.A(n_385),
.Y(n_610)
);

CKINVDCx5p33_ASAP7_75t_R g611 ( 
.A(n_547),
.Y(n_611)
);

BUFx6f_ASAP7_75t_L g612 ( 
.A(n_360),
.Y(n_612)
);

CKINVDCx5p33_ASAP7_75t_R g613 ( 
.A(n_256),
.Y(n_613)
);

INVx2_ASAP7_75t_SL g614 ( 
.A(n_245),
.Y(n_614)
);

CKINVDCx5p33_ASAP7_75t_R g615 ( 
.A(n_310),
.Y(n_615)
);

CKINVDCx20_ASAP7_75t_R g616 ( 
.A(n_490),
.Y(n_616)
);

INVx2_ASAP7_75t_L g617 ( 
.A(n_444),
.Y(n_617)
);

INVx1_ASAP7_75t_L g618 ( 
.A(n_204),
.Y(n_618)
);

INVx2_ASAP7_75t_L g619 ( 
.A(n_320),
.Y(n_619)
);

CKINVDCx5p33_ASAP7_75t_R g620 ( 
.A(n_266),
.Y(n_620)
);

CKINVDCx5p33_ASAP7_75t_R g621 ( 
.A(n_384),
.Y(n_621)
);

CKINVDCx5p33_ASAP7_75t_R g622 ( 
.A(n_47),
.Y(n_622)
);

CKINVDCx5p33_ASAP7_75t_R g623 ( 
.A(n_288),
.Y(n_623)
);

INVx1_ASAP7_75t_L g624 ( 
.A(n_448),
.Y(n_624)
);

INVx1_ASAP7_75t_L g625 ( 
.A(n_158),
.Y(n_625)
);

CKINVDCx20_ASAP7_75t_R g626 ( 
.A(n_493),
.Y(n_626)
);

BUFx3_ASAP7_75t_L g627 ( 
.A(n_258),
.Y(n_627)
);

INVx1_ASAP7_75t_L g628 ( 
.A(n_81),
.Y(n_628)
);

CKINVDCx5p33_ASAP7_75t_R g629 ( 
.A(n_381),
.Y(n_629)
);

INVx1_ASAP7_75t_L g630 ( 
.A(n_123),
.Y(n_630)
);

CKINVDCx5p33_ASAP7_75t_R g631 ( 
.A(n_29),
.Y(n_631)
);

CKINVDCx5p33_ASAP7_75t_R g632 ( 
.A(n_114),
.Y(n_632)
);

CKINVDCx5p33_ASAP7_75t_R g633 ( 
.A(n_184),
.Y(n_633)
);

BUFx2_ASAP7_75t_L g634 ( 
.A(n_267),
.Y(n_634)
);

CKINVDCx5p33_ASAP7_75t_R g635 ( 
.A(n_537),
.Y(n_635)
);

CKINVDCx5p33_ASAP7_75t_R g636 ( 
.A(n_482),
.Y(n_636)
);

INVx2_ASAP7_75t_L g637 ( 
.A(n_176),
.Y(n_637)
);

INVx1_ASAP7_75t_L g638 ( 
.A(n_256),
.Y(n_638)
);

INVx1_ASAP7_75t_L g639 ( 
.A(n_344),
.Y(n_639)
);

CKINVDCx5p33_ASAP7_75t_R g640 ( 
.A(n_509),
.Y(n_640)
);

INVx1_ASAP7_75t_L g641 ( 
.A(n_301),
.Y(n_641)
);

CKINVDCx5p33_ASAP7_75t_R g642 ( 
.A(n_49),
.Y(n_642)
);

INVx1_ASAP7_75t_L g643 ( 
.A(n_382),
.Y(n_643)
);

CKINVDCx5p33_ASAP7_75t_R g644 ( 
.A(n_162),
.Y(n_644)
);

CKINVDCx5p33_ASAP7_75t_R g645 ( 
.A(n_92),
.Y(n_645)
);

INVx1_ASAP7_75t_L g646 ( 
.A(n_70),
.Y(n_646)
);

CKINVDCx5p33_ASAP7_75t_R g647 ( 
.A(n_445),
.Y(n_647)
);

CKINVDCx5p33_ASAP7_75t_R g648 ( 
.A(n_473),
.Y(n_648)
);

CKINVDCx14_ASAP7_75t_R g649 ( 
.A(n_288),
.Y(n_649)
);

CKINVDCx5p33_ASAP7_75t_R g650 ( 
.A(n_99),
.Y(n_650)
);

BUFx3_ASAP7_75t_L g651 ( 
.A(n_423),
.Y(n_651)
);

CKINVDCx5p33_ASAP7_75t_R g652 ( 
.A(n_208),
.Y(n_652)
);

INVx1_ASAP7_75t_L g653 ( 
.A(n_387),
.Y(n_653)
);

CKINVDCx5p33_ASAP7_75t_R g654 ( 
.A(n_525),
.Y(n_654)
);

CKINVDCx5p33_ASAP7_75t_R g655 ( 
.A(n_251),
.Y(n_655)
);

BUFx6f_ASAP7_75t_L g656 ( 
.A(n_270),
.Y(n_656)
);

INVx1_ASAP7_75t_L g657 ( 
.A(n_188),
.Y(n_657)
);

CKINVDCx5p33_ASAP7_75t_R g658 ( 
.A(n_183),
.Y(n_658)
);

INVx1_ASAP7_75t_L g659 ( 
.A(n_124),
.Y(n_659)
);

BUFx6f_ASAP7_75t_L g660 ( 
.A(n_127),
.Y(n_660)
);

INVx1_ASAP7_75t_L g661 ( 
.A(n_41),
.Y(n_661)
);

INVx3_ASAP7_75t_L g662 ( 
.A(n_336),
.Y(n_662)
);

BUFx3_ASAP7_75t_L g663 ( 
.A(n_499),
.Y(n_663)
);

CKINVDCx5p33_ASAP7_75t_R g664 ( 
.A(n_485),
.Y(n_664)
);

INVx1_ASAP7_75t_L g665 ( 
.A(n_406),
.Y(n_665)
);

BUFx3_ASAP7_75t_L g666 ( 
.A(n_345),
.Y(n_666)
);

INVx1_ASAP7_75t_SL g667 ( 
.A(n_386),
.Y(n_667)
);

CKINVDCx20_ASAP7_75t_R g668 ( 
.A(n_197),
.Y(n_668)
);

INVx2_ASAP7_75t_L g669 ( 
.A(n_218),
.Y(n_669)
);

INVx2_ASAP7_75t_L g670 ( 
.A(n_281),
.Y(n_670)
);

CKINVDCx5p33_ASAP7_75t_R g671 ( 
.A(n_441),
.Y(n_671)
);

CKINVDCx5p33_ASAP7_75t_R g672 ( 
.A(n_128),
.Y(n_672)
);

CKINVDCx5p33_ASAP7_75t_R g673 ( 
.A(n_17),
.Y(n_673)
);

INVx1_ASAP7_75t_L g674 ( 
.A(n_394),
.Y(n_674)
);

CKINVDCx20_ASAP7_75t_R g675 ( 
.A(n_380),
.Y(n_675)
);

CKINVDCx5p33_ASAP7_75t_R g676 ( 
.A(n_422),
.Y(n_676)
);

INVx1_ASAP7_75t_L g677 ( 
.A(n_401),
.Y(n_677)
);

CKINVDCx5p33_ASAP7_75t_R g678 ( 
.A(n_93),
.Y(n_678)
);

CKINVDCx5p33_ASAP7_75t_R g679 ( 
.A(n_58),
.Y(n_679)
);

INVx3_ASAP7_75t_L g680 ( 
.A(n_363),
.Y(n_680)
);

INVx1_ASAP7_75t_L g681 ( 
.A(n_548),
.Y(n_681)
);

BUFx3_ASAP7_75t_L g682 ( 
.A(n_489),
.Y(n_682)
);

INVx2_ASAP7_75t_SL g683 ( 
.A(n_40),
.Y(n_683)
);

CKINVDCx5p33_ASAP7_75t_R g684 ( 
.A(n_495),
.Y(n_684)
);

CKINVDCx5p33_ASAP7_75t_R g685 ( 
.A(n_252),
.Y(n_685)
);

CKINVDCx16_ASAP7_75t_R g686 ( 
.A(n_246),
.Y(n_686)
);

CKINVDCx5p33_ASAP7_75t_R g687 ( 
.A(n_369),
.Y(n_687)
);

CKINVDCx5p33_ASAP7_75t_R g688 ( 
.A(n_178),
.Y(n_688)
);

CKINVDCx5p33_ASAP7_75t_R g689 ( 
.A(n_64),
.Y(n_689)
);

INVx1_ASAP7_75t_L g690 ( 
.A(n_159),
.Y(n_690)
);

INVx1_ASAP7_75t_L g691 ( 
.A(n_22),
.Y(n_691)
);

CKINVDCx5p33_ASAP7_75t_R g692 ( 
.A(n_29),
.Y(n_692)
);

CKINVDCx5p33_ASAP7_75t_R g693 ( 
.A(n_133),
.Y(n_693)
);

CKINVDCx5p33_ASAP7_75t_R g694 ( 
.A(n_10),
.Y(n_694)
);

CKINVDCx5p33_ASAP7_75t_R g695 ( 
.A(n_113),
.Y(n_695)
);

CKINVDCx5p33_ASAP7_75t_R g696 ( 
.A(n_425),
.Y(n_696)
);

CKINVDCx5p33_ASAP7_75t_R g697 ( 
.A(n_510),
.Y(n_697)
);

CKINVDCx5p33_ASAP7_75t_R g698 ( 
.A(n_35),
.Y(n_698)
);

INVx1_ASAP7_75t_L g699 ( 
.A(n_118),
.Y(n_699)
);

INVx1_ASAP7_75t_L g700 ( 
.A(n_358),
.Y(n_700)
);

CKINVDCx16_ASAP7_75t_R g701 ( 
.A(n_33),
.Y(n_701)
);

INVx1_ASAP7_75t_L g702 ( 
.A(n_201),
.Y(n_702)
);

CKINVDCx5p33_ASAP7_75t_R g703 ( 
.A(n_14),
.Y(n_703)
);

BUFx6f_ASAP7_75t_L g704 ( 
.A(n_69),
.Y(n_704)
);

BUFx3_ASAP7_75t_L g705 ( 
.A(n_90),
.Y(n_705)
);

INVx1_ASAP7_75t_L g706 ( 
.A(n_361),
.Y(n_706)
);

INVx1_ASAP7_75t_L g707 ( 
.A(n_501),
.Y(n_707)
);

INVx1_ASAP7_75t_L g708 ( 
.A(n_96),
.Y(n_708)
);

BUFx5_ASAP7_75t_L g709 ( 
.A(n_544),
.Y(n_709)
);

INVx1_ASAP7_75t_L g710 ( 
.A(n_238),
.Y(n_710)
);

INVx1_ASAP7_75t_L g711 ( 
.A(n_170),
.Y(n_711)
);

INVx1_ASAP7_75t_L g712 ( 
.A(n_378),
.Y(n_712)
);

INVx1_ASAP7_75t_L g713 ( 
.A(n_442),
.Y(n_713)
);

CKINVDCx5p33_ASAP7_75t_R g714 ( 
.A(n_167),
.Y(n_714)
);

CKINVDCx5p33_ASAP7_75t_R g715 ( 
.A(n_237),
.Y(n_715)
);

INVx1_ASAP7_75t_L g716 ( 
.A(n_438),
.Y(n_716)
);

CKINVDCx5p33_ASAP7_75t_R g717 ( 
.A(n_223),
.Y(n_717)
);

INVx1_ASAP7_75t_L g718 ( 
.A(n_177),
.Y(n_718)
);

INVx1_ASAP7_75t_L g719 ( 
.A(n_465),
.Y(n_719)
);

CKINVDCx5p33_ASAP7_75t_R g720 ( 
.A(n_421),
.Y(n_720)
);

INVx1_ASAP7_75t_L g721 ( 
.A(n_487),
.Y(n_721)
);

INVx2_ASAP7_75t_L g722 ( 
.A(n_161),
.Y(n_722)
);

CKINVDCx5p33_ASAP7_75t_R g723 ( 
.A(n_188),
.Y(n_723)
);

INVx1_ASAP7_75t_L g724 ( 
.A(n_177),
.Y(n_724)
);

BUFx6f_ASAP7_75t_L g725 ( 
.A(n_43),
.Y(n_725)
);

INVx2_ASAP7_75t_L g726 ( 
.A(n_120),
.Y(n_726)
);

CKINVDCx5p33_ASAP7_75t_R g727 ( 
.A(n_393),
.Y(n_727)
);

INVxp67_ASAP7_75t_L g728 ( 
.A(n_484),
.Y(n_728)
);

INVxp67_ASAP7_75t_L g729 ( 
.A(n_30),
.Y(n_729)
);

INVx1_ASAP7_75t_L g730 ( 
.A(n_186),
.Y(n_730)
);

CKINVDCx5p33_ASAP7_75t_R g731 ( 
.A(n_217),
.Y(n_731)
);

CKINVDCx5p33_ASAP7_75t_R g732 ( 
.A(n_77),
.Y(n_732)
);

CKINVDCx5p33_ASAP7_75t_R g733 ( 
.A(n_455),
.Y(n_733)
);

INVx1_ASAP7_75t_L g734 ( 
.A(n_543),
.Y(n_734)
);

CKINVDCx5p33_ASAP7_75t_R g735 ( 
.A(n_327),
.Y(n_735)
);

CKINVDCx20_ASAP7_75t_R g736 ( 
.A(n_371),
.Y(n_736)
);

CKINVDCx5p33_ASAP7_75t_R g737 ( 
.A(n_179),
.Y(n_737)
);

CKINVDCx5p33_ASAP7_75t_R g738 ( 
.A(n_194),
.Y(n_738)
);

INVx1_ASAP7_75t_L g739 ( 
.A(n_513),
.Y(n_739)
);

CKINVDCx5p33_ASAP7_75t_R g740 ( 
.A(n_443),
.Y(n_740)
);

CKINVDCx5p33_ASAP7_75t_R g741 ( 
.A(n_300),
.Y(n_741)
);

INVx2_ASAP7_75t_L g742 ( 
.A(n_204),
.Y(n_742)
);

CKINVDCx5p33_ASAP7_75t_R g743 ( 
.A(n_542),
.Y(n_743)
);

CKINVDCx5p33_ASAP7_75t_R g744 ( 
.A(n_18),
.Y(n_744)
);

CKINVDCx5p33_ASAP7_75t_R g745 ( 
.A(n_447),
.Y(n_745)
);

CKINVDCx5p33_ASAP7_75t_R g746 ( 
.A(n_13),
.Y(n_746)
);

INVx1_ASAP7_75t_L g747 ( 
.A(n_138),
.Y(n_747)
);

CKINVDCx5p33_ASAP7_75t_R g748 ( 
.A(n_306),
.Y(n_748)
);

INVxp67_ASAP7_75t_SL g749 ( 
.A(n_117),
.Y(n_749)
);

CKINVDCx5p33_ASAP7_75t_R g750 ( 
.A(n_494),
.Y(n_750)
);

INVx1_ASAP7_75t_L g751 ( 
.A(n_81),
.Y(n_751)
);

CKINVDCx5p33_ASAP7_75t_R g752 ( 
.A(n_359),
.Y(n_752)
);

INVx1_ASAP7_75t_L g753 ( 
.A(n_316),
.Y(n_753)
);

CKINVDCx5p33_ASAP7_75t_R g754 ( 
.A(n_123),
.Y(n_754)
);

BUFx2_ASAP7_75t_L g755 ( 
.A(n_105),
.Y(n_755)
);

INVx1_ASAP7_75t_L g756 ( 
.A(n_209),
.Y(n_756)
);

INVx1_ASAP7_75t_L g757 ( 
.A(n_379),
.Y(n_757)
);

INVx2_ASAP7_75t_L g758 ( 
.A(n_125),
.Y(n_758)
);

CKINVDCx5p33_ASAP7_75t_R g759 ( 
.A(n_48),
.Y(n_759)
);

CKINVDCx14_ASAP7_75t_R g760 ( 
.A(n_315),
.Y(n_760)
);

INVx1_ASAP7_75t_L g761 ( 
.A(n_186),
.Y(n_761)
);

CKINVDCx5p33_ASAP7_75t_R g762 ( 
.A(n_301),
.Y(n_762)
);

CKINVDCx5p33_ASAP7_75t_R g763 ( 
.A(n_481),
.Y(n_763)
);

CKINVDCx5p33_ASAP7_75t_R g764 ( 
.A(n_427),
.Y(n_764)
);

INVx1_ASAP7_75t_L g765 ( 
.A(n_75),
.Y(n_765)
);

CKINVDCx5p33_ASAP7_75t_R g766 ( 
.A(n_45),
.Y(n_766)
);

BUFx2_ASAP7_75t_L g767 ( 
.A(n_500),
.Y(n_767)
);

CKINVDCx5p33_ASAP7_75t_R g768 ( 
.A(n_239),
.Y(n_768)
);

CKINVDCx5p33_ASAP7_75t_R g769 ( 
.A(n_357),
.Y(n_769)
);

BUFx3_ASAP7_75t_L g770 ( 
.A(n_296),
.Y(n_770)
);

CKINVDCx5p33_ASAP7_75t_R g771 ( 
.A(n_59),
.Y(n_771)
);

CKINVDCx5p33_ASAP7_75t_R g772 ( 
.A(n_13),
.Y(n_772)
);

CKINVDCx5p33_ASAP7_75t_R g773 ( 
.A(n_372),
.Y(n_773)
);

CKINVDCx20_ASAP7_75t_R g774 ( 
.A(n_418),
.Y(n_774)
);

CKINVDCx5p33_ASAP7_75t_R g775 ( 
.A(n_140),
.Y(n_775)
);

INVx1_ASAP7_75t_L g776 ( 
.A(n_146),
.Y(n_776)
);

CKINVDCx5p33_ASAP7_75t_R g777 ( 
.A(n_143),
.Y(n_777)
);

INVxp33_ASAP7_75t_SL g778 ( 
.A(n_565),
.Y(n_778)
);

CKINVDCx5p33_ASAP7_75t_R g779 ( 
.A(n_585),
.Y(n_779)
);

INVx2_ASAP7_75t_L g780 ( 
.A(n_557),
.Y(n_780)
);

INVx1_ASAP7_75t_L g781 ( 
.A(n_557),
.Y(n_781)
);

INVx1_ASAP7_75t_L g782 ( 
.A(n_557),
.Y(n_782)
);

INVx1_ASAP7_75t_L g783 ( 
.A(n_557),
.Y(n_783)
);

INVx1_ASAP7_75t_L g784 ( 
.A(n_557),
.Y(n_784)
);

INVx2_ASAP7_75t_L g785 ( 
.A(n_557),
.Y(n_785)
);

INVx1_ASAP7_75t_L g786 ( 
.A(n_557),
.Y(n_786)
);

CKINVDCx20_ASAP7_75t_R g787 ( 
.A(n_585),
.Y(n_787)
);

INVx1_ASAP7_75t_L g788 ( 
.A(n_662),
.Y(n_788)
);

CKINVDCx5p33_ASAP7_75t_R g789 ( 
.A(n_556),
.Y(n_789)
);

INVx3_ASAP7_75t_L g790 ( 
.A(n_612),
.Y(n_790)
);

INVx1_ASAP7_75t_L g791 ( 
.A(n_662),
.Y(n_791)
);

INVxp33_ASAP7_75t_SL g792 ( 
.A(n_565),
.Y(n_792)
);

CKINVDCx16_ASAP7_75t_R g793 ( 
.A(n_686),
.Y(n_793)
);

INVx1_ASAP7_75t_L g794 ( 
.A(n_662),
.Y(n_794)
);

INVx1_ASAP7_75t_L g795 ( 
.A(n_680),
.Y(n_795)
);

INVx1_ASAP7_75t_L g796 ( 
.A(n_680),
.Y(n_796)
);

INVx3_ASAP7_75t_L g797 ( 
.A(n_612),
.Y(n_797)
);

INVxp33_ASAP7_75t_SL g798 ( 
.A(n_571),
.Y(n_798)
);

INVx2_ASAP7_75t_L g799 ( 
.A(n_680),
.Y(n_799)
);

INVx1_ASAP7_75t_L g800 ( 
.A(n_594),
.Y(n_800)
);

INVxp33_ASAP7_75t_SL g801 ( 
.A(n_571),
.Y(n_801)
);

INVxp33_ASAP7_75t_L g802 ( 
.A(n_634),
.Y(n_802)
);

INVxp67_ASAP7_75t_L g803 ( 
.A(n_755),
.Y(n_803)
);

INVxp67_ASAP7_75t_SL g804 ( 
.A(n_767),
.Y(n_804)
);

INVx1_ASAP7_75t_L g805 ( 
.A(n_594),
.Y(n_805)
);

INVx1_ASAP7_75t_L g806 ( 
.A(n_627),
.Y(n_806)
);

INVxp67_ASAP7_75t_L g807 ( 
.A(n_559),
.Y(n_807)
);

INVxp67_ASAP7_75t_SL g808 ( 
.A(n_651),
.Y(n_808)
);

BUFx3_ASAP7_75t_L g809 ( 
.A(n_651),
.Y(n_809)
);

INVxp33_ASAP7_75t_L g810 ( 
.A(n_595),
.Y(n_810)
);

INVx1_ASAP7_75t_L g811 ( 
.A(n_627),
.Y(n_811)
);

INVxp67_ASAP7_75t_SL g812 ( 
.A(n_663),
.Y(n_812)
);

INVx2_ASAP7_75t_L g813 ( 
.A(n_709),
.Y(n_813)
);

INVx1_ASAP7_75t_L g814 ( 
.A(n_666),
.Y(n_814)
);

INVx1_ASAP7_75t_L g815 ( 
.A(n_666),
.Y(n_815)
);

INVx1_ASAP7_75t_L g816 ( 
.A(n_705),
.Y(n_816)
);

INVx1_ASAP7_75t_L g817 ( 
.A(n_705),
.Y(n_817)
);

INVx1_ASAP7_75t_L g818 ( 
.A(n_770),
.Y(n_818)
);

INVx1_ASAP7_75t_L g819 ( 
.A(n_770),
.Y(n_819)
);

INVxp67_ASAP7_75t_SL g820 ( 
.A(n_663),
.Y(n_820)
);

INVx1_ASAP7_75t_L g821 ( 
.A(n_612),
.Y(n_821)
);

INVx1_ASAP7_75t_L g822 ( 
.A(n_612),
.Y(n_822)
);

INVx1_ASAP7_75t_SL g823 ( 
.A(n_701),
.Y(n_823)
);

INVx1_ASAP7_75t_L g824 ( 
.A(n_656),
.Y(n_824)
);

INVx1_ASAP7_75t_L g825 ( 
.A(n_656),
.Y(n_825)
);

BUFx6f_ASAP7_75t_L g826 ( 
.A(n_682),
.Y(n_826)
);

INVx1_ASAP7_75t_L g827 ( 
.A(n_656),
.Y(n_827)
);

INVx1_ASAP7_75t_L g828 ( 
.A(n_656),
.Y(n_828)
);

INVx1_ASAP7_75t_L g829 ( 
.A(n_660),
.Y(n_829)
);

INVx1_ASAP7_75t_L g830 ( 
.A(n_660),
.Y(n_830)
);

CKINVDCx16_ASAP7_75t_R g831 ( 
.A(n_649),
.Y(n_831)
);

INVxp67_ASAP7_75t_L g832 ( 
.A(n_562),
.Y(n_832)
);

INVxp67_ASAP7_75t_SL g833 ( 
.A(n_682),
.Y(n_833)
);

INVx1_ASAP7_75t_L g834 ( 
.A(n_660),
.Y(n_834)
);

INVx1_ASAP7_75t_L g835 ( 
.A(n_660),
.Y(n_835)
);

BUFx5_ASAP7_75t_L g836 ( 
.A(n_589),
.Y(n_836)
);

INVxp67_ASAP7_75t_SL g837 ( 
.A(n_728),
.Y(n_837)
);

INVx1_ASAP7_75t_L g838 ( 
.A(n_704),
.Y(n_838)
);

CKINVDCx5p33_ASAP7_75t_R g839 ( 
.A(n_760),
.Y(n_839)
);

CKINVDCx5p33_ASAP7_75t_R g840 ( 
.A(n_560),
.Y(n_840)
);

CKINVDCx5p33_ASAP7_75t_R g841 ( 
.A(n_558),
.Y(n_841)
);

INVx1_ASAP7_75t_L g842 ( 
.A(n_704),
.Y(n_842)
);

NOR2xp67_ASAP7_75t_L g843 ( 
.A(n_729),
.B(n_0),
.Y(n_843)
);

INVx1_ASAP7_75t_L g844 ( 
.A(n_704),
.Y(n_844)
);

BUFx5_ASAP7_75t_L g845 ( 
.A(n_606),
.Y(n_845)
);

BUFx2_ASAP7_75t_L g846 ( 
.A(n_572),
.Y(n_846)
);

INVx1_ASAP7_75t_L g847 ( 
.A(n_704),
.Y(n_847)
);

INVx1_ASAP7_75t_L g848 ( 
.A(n_725),
.Y(n_848)
);

INVxp67_ASAP7_75t_L g849 ( 
.A(n_570),
.Y(n_849)
);

CKINVDCx5p33_ASAP7_75t_R g850 ( 
.A(n_563),
.Y(n_850)
);

INVxp33_ASAP7_75t_L g851 ( 
.A(n_595),
.Y(n_851)
);

INVx1_ASAP7_75t_L g852 ( 
.A(n_725),
.Y(n_852)
);

CKINVDCx5p33_ASAP7_75t_R g853 ( 
.A(n_564),
.Y(n_853)
);

INVx1_ASAP7_75t_L g854 ( 
.A(n_725),
.Y(n_854)
);

BUFx2_ASAP7_75t_L g855 ( 
.A(n_572),
.Y(n_855)
);

CKINVDCx5p33_ASAP7_75t_R g856 ( 
.A(n_587),
.Y(n_856)
);

INVx1_ASAP7_75t_L g857 ( 
.A(n_725),
.Y(n_857)
);

INVxp67_ASAP7_75t_L g858 ( 
.A(n_577),
.Y(n_858)
);

INVxp67_ASAP7_75t_SL g859 ( 
.A(n_610),
.Y(n_859)
);

INVxp67_ASAP7_75t_SL g860 ( 
.A(n_624),
.Y(n_860)
);

INVx1_ASAP7_75t_L g861 ( 
.A(n_605),
.Y(n_861)
);

CKINVDCx14_ASAP7_75t_R g862 ( 
.A(n_566),
.Y(n_862)
);

CKINVDCx5p33_ASAP7_75t_R g863 ( 
.A(n_588),
.Y(n_863)
);

CKINVDCx20_ASAP7_75t_R g864 ( 
.A(n_568),
.Y(n_864)
);

INVx1_ASAP7_75t_L g865 ( 
.A(n_609),
.Y(n_865)
);

INVx1_ASAP7_75t_L g866 ( 
.A(n_618),
.Y(n_866)
);

INVxp67_ASAP7_75t_SL g867 ( 
.A(n_643),
.Y(n_867)
);

INVxp33_ASAP7_75t_L g868 ( 
.A(n_619),
.Y(n_868)
);

INVx1_ASAP7_75t_L g869 ( 
.A(n_625),
.Y(n_869)
);

INVxp67_ASAP7_75t_SL g870 ( 
.A(n_653),
.Y(n_870)
);

INVxp33_ASAP7_75t_SL g871 ( 
.A(n_573),
.Y(n_871)
);

INVxp33_ASAP7_75t_L g872 ( 
.A(n_619),
.Y(n_872)
);

INVxp33_ASAP7_75t_L g873 ( 
.A(n_637),
.Y(n_873)
);

INVx1_ASAP7_75t_L g874 ( 
.A(n_628),
.Y(n_874)
);

INVxp67_ASAP7_75t_SL g875 ( 
.A(n_665),
.Y(n_875)
);

CKINVDCx20_ASAP7_75t_R g876 ( 
.A(n_568),
.Y(n_876)
);

INVx1_ASAP7_75t_L g877 ( 
.A(n_630),
.Y(n_877)
);

INVx1_ASAP7_75t_L g878 ( 
.A(n_638),
.Y(n_878)
);

INVx1_ASAP7_75t_L g879 ( 
.A(n_639),
.Y(n_879)
);

BUFx12f_ASAP7_75t_L g880 ( 
.A(n_839),
.Y(n_880)
);

INVx2_ASAP7_75t_SL g881 ( 
.A(n_809),
.Y(n_881)
);

AND2x6_ASAP7_75t_L g882 ( 
.A(n_780),
.B(n_617),
.Y(n_882)
);

INVx1_ASAP7_75t_L g883 ( 
.A(n_790),
.Y(n_883)
);

INVx1_ASAP7_75t_L g884 ( 
.A(n_790),
.Y(n_884)
);

NAND2xp5_ASAP7_75t_L g885 ( 
.A(n_789),
.B(n_574),
.Y(n_885)
);

BUFx6f_ASAP7_75t_L g886 ( 
.A(n_790),
.Y(n_886)
);

INVx1_ASAP7_75t_L g887 ( 
.A(n_797),
.Y(n_887)
);

INVx2_ASAP7_75t_L g888 ( 
.A(n_797),
.Y(n_888)
);

AND2x4_ASAP7_75t_L g889 ( 
.A(n_799),
.B(n_574),
.Y(n_889)
);

INVx3_ASAP7_75t_L g890 ( 
.A(n_780),
.Y(n_890)
);

HB1xp67_ASAP7_75t_L g891 ( 
.A(n_823),
.Y(n_891)
);

CKINVDCx5p33_ASAP7_75t_R g892 ( 
.A(n_840),
.Y(n_892)
);

HB1xp67_ASAP7_75t_L g893 ( 
.A(n_841),
.Y(n_893)
);

INVx2_ASAP7_75t_L g894 ( 
.A(n_797),
.Y(n_894)
);

BUFx6f_ASAP7_75t_L g895 ( 
.A(n_799),
.Y(n_895)
);

CKINVDCx5p33_ASAP7_75t_R g896 ( 
.A(n_862),
.Y(n_896)
);

CKINVDCx6p67_ASAP7_75t_R g897 ( 
.A(n_831),
.Y(n_897)
);

INVx2_ASAP7_75t_L g898 ( 
.A(n_785),
.Y(n_898)
);

NAND2xp5_ASAP7_75t_L g899 ( 
.A(n_808),
.B(n_617),
.Y(n_899)
);

INVx1_ASAP7_75t_L g900 ( 
.A(n_821),
.Y(n_900)
);

INVx2_ASAP7_75t_L g901 ( 
.A(n_785),
.Y(n_901)
);

BUFx8_ASAP7_75t_L g902 ( 
.A(n_846),
.Y(n_902)
);

CKINVDCx6p67_ASAP7_75t_R g903 ( 
.A(n_787),
.Y(n_903)
);

INVx1_ASAP7_75t_L g904 ( 
.A(n_822),
.Y(n_904)
);

AND2x4_ASAP7_75t_L g905 ( 
.A(n_788),
.B(n_674),
.Y(n_905)
);

AND2x2_ASAP7_75t_SL g906 ( 
.A(n_826),
.B(n_677),
.Y(n_906)
);

CKINVDCx5p33_ASAP7_75t_R g907 ( 
.A(n_862),
.Y(n_907)
);

BUFx12f_ASAP7_75t_L g908 ( 
.A(n_839),
.Y(n_908)
);

NAND2xp5_ASAP7_75t_L g909 ( 
.A(n_812),
.B(n_681),
.Y(n_909)
);

INVx1_ASAP7_75t_L g910 ( 
.A(n_824),
.Y(n_910)
);

AND2x2_ASAP7_75t_L g911 ( 
.A(n_820),
.B(n_614),
.Y(n_911)
);

BUFx6f_ASAP7_75t_L g912 ( 
.A(n_825),
.Y(n_912)
);

NAND2xp5_ASAP7_75t_L g913 ( 
.A(n_833),
.B(n_707),
.Y(n_913)
);

INVx2_ASAP7_75t_L g914 ( 
.A(n_781),
.Y(n_914)
);

AND2x4_ASAP7_75t_L g915 ( 
.A(n_791),
.B(n_712),
.Y(n_915)
);

INVx1_ASAP7_75t_L g916 ( 
.A(n_827),
.Y(n_916)
);

INVx1_ASAP7_75t_L g917 ( 
.A(n_828),
.Y(n_917)
);

BUFx12f_ASAP7_75t_L g918 ( 
.A(n_779),
.Y(n_918)
);

INVx2_ASAP7_75t_L g919 ( 
.A(n_782),
.Y(n_919)
);

OAI22xp5_ASAP7_75t_SL g920 ( 
.A1(n_864),
.A2(n_581),
.B1(n_668),
.B2(n_584),
.Y(n_920)
);

INVx3_ASAP7_75t_L g921 ( 
.A(n_783),
.Y(n_921)
);

INVx1_ASAP7_75t_L g922 ( 
.A(n_829),
.Y(n_922)
);

INVxp33_ASAP7_75t_L g923 ( 
.A(n_855),
.Y(n_923)
);

AND2x4_ASAP7_75t_SL g924 ( 
.A(n_787),
.B(n_582),
.Y(n_924)
);

INVx3_ASAP7_75t_L g925 ( 
.A(n_784),
.Y(n_925)
);

AOI22x1_ASAP7_75t_SL g926 ( 
.A1(n_864),
.A2(n_584),
.B1(n_668),
.B2(n_581),
.Y(n_926)
);

INVx5_ASAP7_75t_L g927 ( 
.A(n_826),
.Y(n_927)
);

AND2x4_ASAP7_75t_L g928 ( 
.A(n_794),
.B(n_713),
.Y(n_928)
);

AOI22xp5_ASAP7_75t_L g929 ( 
.A1(n_803),
.A2(n_736),
.B1(n_616),
.B2(n_626),
.Y(n_929)
);

BUFx8_ASAP7_75t_SL g930 ( 
.A(n_876),
.Y(n_930)
);

INVx1_ASAP7_75t_L g931 ( 
.A(n_830),
.Y(n_931)
);

INVx2_ASAP7_75t_L g932 ( 
.A(n_786),
.Y(n_932)
);

INVxp67_ASAP7_75t_L g933 ( 
.A(n_841),
.Y(n_933)
);

BUFx2_ASAP7_75t_L g934 ( 
.A(n_850),
.Y(n_934)
);

INVx1_ASAP7_75t_L g935 ( 
.A(n_834),
.Y(n_935)
);

BUFx6f_ASAP7_75t_L g936 ( 
.A(n_835),
.Y(n_936)
);

BUFx2_ASAP7_75t_L g937 ( 
.A(n_850),
.Y(n_937)
);

INVx3_ASAP7_75t_L g938 ( 
.A(n_813),
.Y(n_938)
);

NOR2xp33_ASAP7_75t_SL g939 ( 
.A(n_793),
.B(n_582),
.Y(n_939)
);

INVx5_ASAP7_75t_L g940 ( 
.A(n_826),
.Y(n_940)
);

BUFx2_ASAP7_75t_L g941 ( 
.A(n_853),
.Y(n_941)
);

NAND2xp5_ASAP7_75t_L g942 ( 
.A(n_837),
.B(n_716),
.Y(n_942)
);

BUFx6f_ASAP7_75t_L g943 ( 
.A(n_838),
.Y(n_943)
);

BUFx6f_ASAP7_75t_L g944 ( 
.A(n_842),
.Y(n_944)
);

INVx2_ASAP7_75t_L g945 ( 
.A(n_844),
.Y(n_945)
);

INVx4_ASAP7_75t_L g946 ( 
.A(n_927),
.Y(n_946)
);

INVx1_ASAP7_75t_L g947 ( 
.A(n_898),
.Y(n_947)
);

INVx1_ASAP7_75t_L g948 ( 
.A(n_898),
.Y(n_948)
);

CKINVDCx5p33_ASAP7_75t_R g949 ( 
.A(n_930),
.Y(n_949)
);

BUFx2_ASAP7_75t_L g950 ( 
.A(n_891),
.Y(n_950)
);

CKINVDCx20_ASAP7_75t_R g951 ( 
.A(n_897),
.Y(n_951)
);

CKINVDCx5p33_ASAP7_75t_R g952 ( 
.A(n_896),
.Y(n_952)
);

INVx1_ASAP7_75t_L g953 ( 
.A(n_914),
.Y(n_953)
);

INVx3_ASAP7_75t_L g954 ( 
.A(n_938),
.Y(n_954)
);

NAND2xp5_ASAP7_75t_L g955 ( 
.A(n_906),
.B(n_859),
.Y(n_955)
);

INVxp67_ASAP7_75t_L g956 ( 
.A(n_934),
.Y(n_956)
);

INVx1_ASAP7_75t_L g957 ( 
.A(n_914),
.Y(n_957)
);

XNOR2xp5_ASAP7_75t_L g958 ( 
.A(n_929),
.B(n_876),
.Y(n_958)
);

INVx1_ASAP7_75t_L g959 ( 
.A(n_901),
.Y(n_959)
);

CKINVDCx5p33_ASAP7_75t_R g960 ( 
.A(n_896),
.Y(n_960)
);

INVx1_ASAP7_75t_L g961 ( 
.A(n_901),
.Y(n_961)
);

INVx2_ASAP7_75t_L g962 ( 
.A(n_890),
.Y(n_962)
);

NOR2xp33_ASAP7_75t_L g963 ( 
.A(n_885),
.B(n_778),
.Y(n_963)
);

INVx1_ASAP7_75t_L g964 ( 
.A(n_919),
.Y(n_964)
);

INVx1_ASAP7_75t_L g965 ( 
.A(n_919),
.Y(n_965)
);

HB1xp67_ASAP7_75t_L g966 ( 
.A(n_881),
.Y(n_966)
);

HB1xp67_ASAP7_75t_L g967 ( 
.A(n_881),
.Y(n_967)
);

INVx4_ASAP7_75t_L g968 ( 
.A(n_927),
.Y(n_968)
);

INVx1_ASAP7_75t_L g969 ( 
.A(n_932),
.Y(n_969)
);

XNOR2xp5_ASAP7_75t_L g970 ( 
.A(n_929),
.B(n_736),
.Y(n_970)
);

BUFx6f_ASAP7_75t_L g971 ( 
.A(n_886),
.Y(n_971)
);

INVx3_ASAP7_75t_L g972 ( 
.A(n_938),
.Y(n_972)
);

NAND2xp5_ASAP7_75t_SL g973 ( 
.A(n_907),
.B(n_853),
.Y(n_973)
);

CKINVDCx20_ASAP7_75t_R g974 ( 
.A(n_892),
.Y(n_974)
);

CKINVDCx5p33_ASAP7_75t_R g975 ( 
.A(n_907),
.Y(n_975)
);

INVx1_ASAP7_75t_L g976 ( 
.A(n_932),
.Y(n_976)
);

INVx2_ASAP7_75t_L g977 ( 
.A(n_890),
.Y(n_977)
);

INVx2_ASAP7_75t_L g978 ( 
.A(n_890),
.Y(n_978)
);

BUFx6f_ASAP7_75t_L g979 ( 
.A(n_886),
.Y(n_979)
);

INVx1_ASAP7_75t_L g980 ( 
.A(n_921),
.Y(n_980)
);

NAND2xp5_ASAP7_75t_L g981 ( 
.A(n_906),
.B(n_911),
.Y(n_981)
);

INVx1_ASAP7_75t_L g982 ( 
.A(n_921),
.Y(n_982)
);

INVx1_ASAP7_75t_L g983 ( 
.A(n_921),
.Y(n_983)
);

INVx2_ASAP7_75t_L g984 ( 
.A(n_895),
.Y(n_984)
);

BUFx2_ASAP7_75t_L g985 ( 
.A(n_934),
.Y(n_985)
);

INVx1_ASAP7_75t_L g986 ( 
.A(n_925),
.Y(n_986)
);

INVx1_ASAP7_75t_L g987 ( 
.A(n_925),
.Y(n_987)
);

BUFx2_ASAP7_75t_L g988 ( 
.A(n_937),
.Y(n_988)
);

CKINVDCx5p33_ASAP7_75t_R g989 ( 
.A(n_880),
.Y(n_989)
);

CKINVDCx5p33_ASAP7_75t_R g990 ( 
.A(n_880),
.Y(n_990)
);

INVx2_ASAP7_75t_L g991 ( 
.A(n_895),
.Y(n_991)
);

INVx2_ASAP7_75t_L g992 ( 
.A(n_895),
.Y(n_992)
);

CKINVDCx5p33_ASAP7_75t_R g993 ( 
.A(n_908),
.Y(n_993)
);

AND2x2_ASAP7_75t_SL g994 ( 
.A(n_906),
.B(n_719),
.Y(n_994)
);

INVx1_ASAP7_75t_L g995 ( 
.A(n_925),
.Y(n_995)
);

NOR2xp33_ASAP7_75t_SL g996 ( 
.A(n_908),
.B(n_616),
.Y(n_996)
);

INVx1_ASAP7_75t_L g997 ( 
.A(n_938),
.Y(n_997)
);

OA21x2_ASAP7_75t_L g998 ( 
.A1(n_899),
.A2(n_796),
.B(n_795),
.Y(n_998)
);

INVx1_ASAP7_75t_L g999 ( 
.A(n_883),
.Y(n_999)
);

CKINVDCx20_ASAP7_75t_R g1000 ( 
.A(n_892),
.Y(n_1000)
);

NAND2xp5_ASAP7_75t_L g1001 ( 
.A(n_911),
.B(n_860),
.Y(n_1001)
);

CKINVDCx5p33_ASAP7_75t_R g1002 ( 
.A(n_902),
.Y(n_1002)
);

INVx1_ASAP7_75t_L g1003 ( 
.A(n_883),
.Y(n_1003)
);

INVx1_ASAP7_75t_L g1004 ( 
.A(n_884),
.Y(n_1004)
);

INVx2_ASAP7_75t_L g1005 ( 
.A(n_895),
.Y(n_1005)
);

INVx1_ASAP7_75t_L g1006 ( 
.A(n_884),
.Y(n_1006)
);

INVx3_ASAP7_75t_L g1007 ( 
.A(n_895),
.Y(n_1007)
);

INVx2_ASAP7_75t_L g1008 ( 
.A(n_888),
.Y(n_1008)
);

INVx3_ASAP7_75t_L g1009 ( 
.A(n_886),
.Y(n_1009)
);

AND2x2_ASAP7_75t_L g1010 ( 
.A(n_905),
.B(n_809),
.Y(n_1010)
);

HB1xp67_ASAP7_75t_L g1011 ( 
.A(n_893),
.Y(n_1011)
);

INVxp67_ASAP7_75t_L g1012 ( 
.A(n_937),
.Y(n_1012)
);

INVx2_ASAP7_75t_L g1013 ( 
.A(n_888),
.Y(n_1013)
);

INVx2_ASAP7_75t_L g1014 ( 
.A(n_894),
.Y(n_1014)
);

INVx2_ASAP7_75t_L g1015 ( 
.A(n_894),
.Y(n_1015)
);

INVx1_ASAP7_75t_L g1016 ( 
.A(n_887),
.Y(n_1016)
);

INVx1_ASAP7_75t_L g1017 ( 
.A(n_887),
.Y(n_1017)
);

INVx1_ASAP7_75t_L g1018 ( 
.A(n_900),
.Y(n_1018)
);

INVx2_ASAP7_75t_L g1019 ( 
.A(n_945),
.Y(n_1019)
);

NAND2xp5_ASAP7_75t_L g1020 ( 
.A(n_909),
.B(n_867),
.Y(n_1020)
);

INVx2_ASAP7_75t_L g1021 ( 
.A(n_945),
.Y(n_1021)
);

CKINVDCx5p33_ASAP7_75t_R g1022 ( 
.A(n_902),
.Y(n_1022)
);

NAND2xp5_ASAP7_75t_L g1023 ( 
.A(n_913),
.B(n_870),
.Y(n_1023)
);

INVx3_ASAP7_75t_L g1024 ( 
.A(n_886),
.Y(n_1024)
);

HB1xp67_ASAP7_75t_L g1025 ( 
.A(n_941),
.Y(n_1025)
);

NAND2xp5_ASAP7_75t_SL g1026 ( 
.A(n_941),
.B(n_856),
.Y(n_1026)
);

CKINVDCx5p33_ASAP7_75t_R g1027 ( 
.A(n_902),
.Y(n_1027)
);

NAND2xp5_ASAP7_75t_L g1028 ( 
.A(n_886),
.B(n_875),
.Y(n_1028)
);

INVx3_ASAP7_75t_L g1029 ( 
.A(n_912),
.Y(n_1029)
);

BUFx2_ASAP7_75t_L g1030 ( 
.A(n_902),
.Y(n_1030)
);

INVx1_ASAP7_75t_L g1031 ( 
.A(n_900),
.Y(n_1031)
);

CKINVDCx20_ASAP7_75t_R g1032 ( 
.A(n_924),
.Y(n_1032)
);

CKINVDCx5p33_ASAP7_75t_R g1033 ( 
.A(n_903),
.Y(n_1033)
);

OAI22xp33_ASAP7_75t_L g1034 ( 
.A1(n_981),
.A2(n_939),
.B1(n_802),
.B2(n_851),
.Y(n_1034)
);

INVx2_ASAP7_75t_L g1035 ( 
.A(n_1019),
.Y(n_1035)
);

INVx1_ASAP7_75t_L g1036 ( 
.A(n_1018),
.Y(n_1036)
);

INVx2_ASAP7_75t_L g1037 ( 
.A(n_1019),
.Y(n_1037)
);

INVx2_ASAP7_75t_L g1038 ( 
.A(n_1021),
.Y(n_1038)
);

AND2x2_ASAP7_75t_L g1039 ( 
.A(n_950),
.B(n_923),
.Y(n_1039)
);

INVx2_ASAP7_75t_L g1040 ( 
.A(n_999),
.Y(n_1040)
);

INVx3_ASAP7_75t_L g1041 ( 
.A(n_954),
.Y(n_1041)
);

BUFx6f_ASAP7_75t_SL g1042 ( 
.A(n_994),
.Y(n_1042)
);

NAND2xp5_ASAP7_75t_L g1043 ( 
.A(n_994),
.B(n_942),
.Y(n_1043)
);

INVx1_ASAP7_75t_L g1044 ( 
.A(n_1018),
.Y(n_1044)
);

INVxp33_ASAP7_75t_L g1045 ( 
.A(n_950),
.Y(n_1045)
);

NAND2xp5_ASAP7_75t_SL g1046 ( 
.A(n_994),
.B(n_955),
.Y(n_1046)
);

INVx1_ASAP7_75t_L g1047 ( 
.A(n_1031),
.Y(n_1047)
);

NAND3xp33_ASAP7_75t_L g1048 ( 
.A(n_963),
.B(n_863),
.C(n_856),
.Y(n_1048)
);

INVx4_ASAP7_75t_L g1049 ( 
.A(n_971),
.Y(n_1049)
);

INVx2_ASAP7_75t_L g1050 ( 
.A(n_999),
.Y(n_1050)
);

NAND2xp5_ASAP7_75t_SL g1051 ( 
.A(n_1001),
.B(n_980),
.Y(n_1051)
);

INVx2_ASAP7_75t_L g1052 ( 
.A(n_1003),
.Y(n_1052)
);

INVx4_ASAP7_75t_L g1053 ( 
.A(n_971),
.Y(n_1053)
);

NAND2xp5_ASAP7_75t_SL g1054 ( 
.A(n_980),
.B(n_982),
.Y(n_1054)
);

BUFx10_ASAP7_75t_L g1055 ( 
.A(n_949),
.Y(n_1055)
);

OAI22xp33_ASAP7_75t_L g1056 ( 
.A1(n_1020),
.A2(n_802),
.B1(n_851),
.B2(n_810),
.Y(n_1056)
);

INVx2_ASAP7_75t_L g1057 ( 
.A(n_1003),
.Y(n_1057)
);

INVx2_ASAP7_75t_L g1058 ( 
.A(n_1004),
.Y(n_1058)
);

NAND2xp5_ASAP7_75t_SL g1059 ( 
.A(n_982),
.B(n_933),
.Y(n_1059)
);

INVx1_ASAP7_75t_SL g1060 ( 
.A(n_985),
.Y(n_1060)
);

INVx2_ASAP7_75t_L g1061 ( 
.A(n_1004),
.Y(n_1061)
);

BUFx4f_ASAP7_75t_L g1062 ( 
.A(n_985),
.Y(n_1062)
);

NAND2xp5_ASAP7_75t_L g1063 ( 
.A(n_1028),
.B(n_905),
.Y(n_1063)
);

AOI22xp5_ASAP7_75t_L g1064 ( 
.A1(n_1010),
.A2(n_626),
.B1(n_774),
.B2(n_675),
.Y(n_1064)
);

INVx2_ASAP7_75t_L g1065 ( 
.A(n_1016),
.Y(n_1065)
);

NAND3xp33_ASAP7_75t_L g1066 ( 
.A(n_1023),
.B(n_863),
.C(n_1010),
.Y(n_1066)
);

BUFx3_ASAP7_75t_L g1067 ( 
.A(n_966),
.Y(n_1067)
);

INVx2_ASAP7_75t_L g1068 ( 
.A(n_1016),
.Y(n_1068)
);

NAND2xp5_ASAP7_75t_SL g1069 ( 
.A(n_995),
.B(n_905),
.Y(n_1069)
);

AND2x4_ASAP7_75t_L g1070 ( 
.A(n_1031),
.B(n_905),
.Y(n_1070)
);

INVx3_ASAP7_75t_L g1071 ( 
.A(n_954),
.Y(n_1071)
);

BUFx10_ASAP7_75t_L g1072 ( 
.A(n_949),
.Y(n_1072)
);

INVx2_ASAP7_75t_L g1073 ( 
.A(n_1017),
.Y(n_1073)
);

INVx2_ASAP7_75t_L g1074 ( 
.A(n_1017),
.Y(n_1074)
);

INVx1_ASAP7_75t_L g1075 ( 
.A(n_995),
.Y(n_1075)
);

BUFx6f_ASAP7_75t_L g1076 ( 
.A(n_971),
.Y(n_1076)
);

NOR2xp33_ASAP7_75t_L g1077 ( 
.A(n_967),
.B(n_778),
.Y(n_1077)
);

INVx1_ASAP7_75t_L g1078 ( 
.A(n_1006),
.Y(n_1078)
);

INVx2_ASAP7_75t_L g1079 ( 
.A(n_947),
.Y(n_1079)
);

NOR2xp33_ASAP7_75t_L g1080 ( 
.A(n_973),
.B(n_792),
.Y(n_1080)
);

INVx4_ASAP7_75t_L g1081 ( 
.A(n_971),
.Y(n_1081)
);

BUFx2_ASAP7_75t_L g1082 ( 
.A(n_988),
.Y(n_1082)
);

NOR2xp33_ASAP7_75t_L g1083 ( 
.A(n_1026),
.B(n_792),
.Y(n_1083)
);

NOR2x1p5_ASAP7_75t_L g1084 ( 
.A(n_1002),
.B(n_903),
.Y(n_1084)
);

INVx5_ASAP7_75t_L g1085 ( 
.A(n_971),
.Y(n_1085)
);

INVx1_ASAP7_75t_L g1086 ( 
.A(n_983),
.Y(n_1086)
);

INVx1_ASAP7_75t_L g1087 ( 
.A(n_986),
.Y(n_1087)
);

NAND2xp5_ASAP7_75t_L g1088 ( 
.A(n_987),
.B(n_928),
.Y(n_1088)
);

BUFx10_ASAP7_75t_L g1089 ( 
.A(n_952),
.Y(n_1089)
);

INVx2_ASAP7_75t_L g1090 ( 
.A(n_947),
.Y(n_1090)
);

NAND2xp5_ASAP7_75t_L g1091 ( 
.A(n_972),
.B(n_928),
.Y(n_1091)
);

INVx2_ASAP7_75t_L g1092 ( 
.A(n_948),
.Y(n_1092)
);

OR2x6_ASAP7_75t_L g1093 ( 
.A(n_1030),
.B(n_918),
.Y(n_1093)
);

NAND2xp5_ASAP7_75t_SL g1094 ( 
.A(n_964),
.B(n_915),
.Y(n_1094)
);

NAND2xp33_ASAP7_75t_L g1095 ( 
.A(n_979),
.B(n_709),
.Y(n_1095)
);

BUFx3_ASAP7_75t_L g1096 ( 
.A(n_988),
.Y(n_1096)
);

OAI22xp5_ASAP7_75t_L g1097 ( 
.A1(n_956),
.A2(n_1012),
.B1(n_774),
.B2(n_675),
.Y(n_1097)
);

INVx1_ASAP7_75t_L g1098 ( 
.A(n_965),
.Y(n_1098)
);

INVx1_ASAP7_75t_L g1099 ( 
.A(n_965),
.Y(n_1099)
);

CKINVDCx20_ASAP7_75t_R g1100 ( 
.A(n_1032),
.Y(n_1100)
);

AO21x2_ASAP7_75t_L g1101 ( 
.A1(n_984),
.A2(n_734),
.B(n_721),
.Y(n_1101)
);

INVx1_ASAP7_75t_L g1102 ( 
.A(n_969),
.Y(n_1102)
);

BUFx6f_ASAP7_75t_L g1103 ( 
.A(n_979),
.Y(n_1103)
);

INVx2_ASAP7_75t_SL g1104 ( 
.A(n_1025),
.Y(n_1104)
);

INVx1_ASAP7_75t_L g1105 ( 
.A(n_969),
.Y(n_1105)
);

INVx2_ASAP7_75t_L g1106 ( 
.A(n_959),
.Y(n_1106)
);

AOI22xp33_ASAP7_75t_L g1107 ( 
.A1(n_998),
.A2(n_637),
.B1(n_670),
.B2(n_669),
.Y(n_1107)
);

INVx1_ASAP7_75t_L g1108 ( 
.A(n_976),
.Y(n_1108)
);

NOR2xp33_ASAP7_75t_L g1109 ( 
.A(n_953),
.B(n_798),
.Y(n_1109)
);

INVx1_ASAP7_75t_L g1110 ( 
.A(n_976),
.Y(n_1110)
);

NOR2x1p5_ASAP7_75t_L g1111 ( 
.A(n_1002),
.B(n_918),
.Y(n_1111)
);

INVx2_ASAP7_75t_L g1112 ( 
.A(n_959),
.Y(n_1112)
);

INVx3_ASAP7_75t_L g1113 ( 
.A(n_1009),
.Y(n_1113)
);

NOR2xp33_ASAP7_75t_L g1114 ( 
.A(n_957),
.B(n_798),
.Y(n_1114)
);

NAND2xp5_ASAP7_75t_L g1115 ( 
.A(n_997),
.B(n_915),
.Y(n_1115)
);

AOI22xp33_ASAP7_75t_SL g1116 ( 
.A1(n_996),
.A2(n_920),
.B1(n_926),
.B2(n_924),
.Y(n_1116)
);

INVx2_ASAP7_75t_SL g1117 ( 
.A(n_1011),
.Y(n_1117)
);

INVx1_ASAP7_75t_L g1118 ( 
.A(n_1008),
.Y(n_1118)
);

NAND3xp33_ASAP7_75t_L g1119 ( 
.A(n_998),
.B(n_804),
.C(n_807),
.Y(n_1119)
);

INVx2_ASAP7_75t_L g1120 ( 
.A(n_961),
.Y(n_1120)
);

BUFx3_ASAP7_75t_L g1121 ( 
.A(n_974),
.Y(n_1121)
);

NOR2xp33_ASAP7_75t_L g1122 ( 
.A(n_998),
.B(n_801),
.Y(n_1122)
);

XOR2xp5_ASAP7_75t_L g1123 ( 
.A(n_1000),
.B(n_926),
.Y(n_1123)
);

INVx2_ASAP7_75t_L g1124 ( 
.A(n_961),
.Y(n_1124)
);

INVx1_ASAP7_75t_L g1125 ( 
.A(n_1008),
.Y(n_1125)
);

AO21x2_ASAP7_75t_L g1126 ( 
.A1(n_984),
.A2(n_757),
.B(n_739),
.Y(n_1126)
);

BUFx6f_ASAP7_75t_L g1127 ( 
.A(n_979),
.Y(n_1127)
);

AOI22xp5_ASAP7_75t_L g1128 ( 
.A1(n_998),
.A2(n_915),
.B1(n_667),
.B2(n_555),
.Y(n_1128)
);

NAND2xp5_ASAP7_75t_SL g1129 ( 
.A(n_991),
.B(n_709),
.Y(n_1129)
);

NAND2xp5_ASAP7_75t_SL g1130 ( 
.A(n_991),
.B(n_709),
.Y(n_1130)
);

INVx3_ASAP7_75t_L g1131 ( 
.A(n_1009),
.Y(n_1131)
);

NAND3xp33_ASAP7_75t_L g1132 ( 
.A(n_952),
.B(n_849),
.C(n_832),
.Y(n_1132)
);

INVx1_ASAP7_75t_L g1133 ( 
.A(n_1013),
.Y(n_1133)
);

NOR2xp33_ASAP7_75t_L g1134 ( 
.A(n_1007),
.B(n_871),
.Y(n_1134)
);

INVx2_ASAP7_75t_L g1135 ( 
.A(n_1014),
.Y(n_1135)
);

INVx3_ASAP7_75t_L g1136 ( 
.A(n_1009),
.Y(n_1136)
);

INVx1_ASAP7_75t_L g1137 ( 
.A(n_1014),
.Y(n_1137)
);

HB1xp67_ASAP7_75t_L g1138 ( 
.A(n_958),
.Y(n_1138)
);

INVx1_ASAP7_75t_SL g1139 ( 
.A(n_960),
.Y(n_1139)
);

INVx1_ASAP7_75t_L g1140 ( 
.A(n_1015),
.Y(n_1140)
);

INVx1_ASAP7_75t_L g1141 ( 
.A(n_1015),
.Y(n_1141)
);

NOR2xp33_ASAP7_75t_L g1142 ( 
.A(n_1007),
.B(n_810),
.Y(n_1142)
);

INVx2_ASAP7_75t_L g1143 ( 
.A(n_962),
.Y(n_1143)
);

INVx2_ASAP7_75t_L g1144 ( 
.A(n_977),
.Y(n_1144)
);

INVx2_ASAP7_75t_L g1145 ( 
.A(n_977),
.Y(n_1145)
);

NAND2xp33_ASAP7_75t_SL g1146 ( 
.A(n_970),
.B(n_614),
.Y(n_1146)
);

BUFx2_ASAP7_75t_L g1147 ( 
.A(n_975),
.Y(n_1147)
);

AOI21x1_ASAP7_75t_L g1148 ( 
.A1(n_992),
.A2(n_935),
.B(n_931),
.Y(n_1148)
);

INVx1_ASAP7_75t_L g1149 ( 
.A(n_978),
.Y(n_1149)
);

OR2x2_ASAP7_75t_L g1150 ( 
.A(n_970),
.B(n_800),
.Y(n_1150)
);

INVx2_ASAP7_75t_L g1151 ( 
.A(n_992),
.Y(n_1151)
);

AND2x2_ASAP7_75t_SL g1152 ( 
.A(n_1030),
.B(n_889),
.Y(n_1152)
);

BUFx3_ASAP7_75t_L g1153 ( 
.A(n_951),
.Y(n_1153)
);

INVx1_ASAP7_75t_L g1154 ( 
.A(n_1005),
.Y(n_1154)
);

INVx2_ASAP7_75t_L g1155 ( 
.A(n_1005),
.Y(n_1155)
);

INVx1_ASAP7_75t_L g1156 ( 
.A(n_1024),
.Y(n_1156)
);

OAI22xp5_ASAP7_75t_L g1157 ( 
.A1(n_1024),
.A2(n_566),
.B1(n_569),
.B2(n_567),
.Y(n_1157)
);

INVx1_ASAP7_75t_L g1158 ( 
.A(n_1024),
.Y(n_1158)
);

INVx1_ASAP7_75t_L g1159 ( 
.A(n_1040),
.Y(n_1159)
);

NAND2xp33_ASAP7_75t_L g1160 ( 
.A(n_1043),
.B(n_1022),
.Y(n_1160)
);

INVx2_ASAP7_75t_L g1161 ( 
.A(n_1040),
.Y(n_1161)
);

INVx1_ASAP7_75t_SL g1162 ( 
.A(n_1060),
.Y(n_1162)
);

INVxp67_ASAP7_75t_L g1163 ( 
.A(n_1039),
.Y(n_1163)
);

NAND2xp33_ASAP7_75t_L g1164 ( 
.A(n_1076),
.B(n_1022),
.Y(n_1164)
);

NAND2xp5_ASAP7_75t_SL g1165 ( 
.A(n_1067),
.B(n_1027),
.Y(n_1165)
);

NAND2xp5_ASAP7_75t_L g1166 ( 
.A(n_1046),
.B(n_1029),
.Y(n_1166)
);

NOR3xp33_ASAP7_75t_L g1167 ( 
.A(n_1097),
.B(n_990),
.C(n_989),
.Y(n_1167)
);

BUFx6f_ASAP7_75t_SL g1168 ( 
.A(n_1089),
.Y(n_1168)
);

NOR2xp33_ASAP7_75t_L g1169 ( 
.A(n_1045),
.B(n_958),
.Y(n_1169)
);

NOR2xp33_ASAP7_75t_L g1170 ( 
.A(n_1045),
.B(n_1033),
.Y(n_1170)
);

INVx1_ASAP7_75t_L g1171 ( 
.A(n_1050),
.Y(n_1171)
);

INVx2_ASAP7_75t_L g1172 ( 
.A(n_1050),
.Y(n_1172)
);

NOR2xp33_ASAP7_75t_L g1173 ( 
.A(n_1077),
.B(n_1033),
.Y(n_1173)
);

NAND2xp5_ASAP7_75t_L g1174 ( 
.A(n_1046),
.B(n_1029),
.Y(n_1174)
);

INVx2_ASAP7_75t_SL g1175 ( 
.A(n_1096),
.Y(n_1175)
);

NOR2xp67_ASAP7_75t_L g1176 ( 
.A(n_1132),
.B(n_1048),
.Y(n_1176)
);

NOR2xp33_ASAP7_75t_L g1177 ( 
.A(n_1083),
.B(n_989),
.Y(n_1177)
);

NAND2xp5_ASAP7_75t_L g1178 ( 
.A(n_1051),
.B(n_1029),
.Y(n_1178)
);

INVx1_ASAP7_75t_L g1179 ( 
.A(n_1052),
.Y(n_1179)
);

OR2x6_ASAP7_75t_L g1180 ( 
.A(n_1093),
.B(n_1096),
.Y(n_1180)
);

INVx2_ASAP7_75t_L g1181 ( 
.A(n_1057),
.Y(n_1181)
);

BUFx3_ASAP7_75t_L g1182 ( 
.A(n_1082),
.Y(n_1182)
);

INVx1_ASAP7_75t_L g1183 ( 
.A(n_1057),
.Y(n_1183)
);

NAND2xp5_ASAP7_75t_L g1184 ( 
.A(n_1051),
.B(n_836),
.Y(n_1184)
);

INVx1_ASAP7_75t_L g1185 ( 
.A(n_1058),
.Y(n_1185)
);

INVx1_ASAP7_75t_L g1186 ( 
.A(n_1058),
.Y(n_1186)
);

NAND2xp5_ASAP7_75t_SL g1187 ( 
.A(n_1067),
.B(n_993),
.Y(n_1187)
);

NAND2xp5_ASAP7_75t_L g1188 ( 
.A(n_1142),
.B(n_979),
.Y(n_1188)
);

INVx2_ASAP7_75t_L g1189 ( 
.A(n_1061),
.Y(n_1189)
);

INVx3_ASAP7_75t_R g1190 ( 
.A(n_1150),
.Y(n_1190)
);

NAND2xp5_ASAP7_75t_L g1191 ( 
.A(n_1142),
.B(n_979),
.Y(n_1191)
);

BUFx5_ASAP7_75t_L g1192 ( 
.A(n_1075),
.Y(n_1192)
);

OAI22xp33_ASAP7_75t_L g1193 ( 
.A1(n_1064),
.A2(n_993),
.B1(n_868),
.B2(n_873),
.Y(n_1193)
);

NAND2xp5_ASAP7_75t_L g1194 ( 
.A(n_1036),
.B(n_889),
.Y(n_1194)
);

INVx2_ASAP7_75t_L g1195 ( 
.A(n_1061),
.Y(n_1195)
);

NAND2xp5_ASAP7_75t_L g1196 ( 
.A(n_1044),
.B(n_889),
.Y(n_1196)
);

INVx2_ASAP7_75t_L g1197 ( 
.A(n_1065),
.Y(n_1197)
);

INVx2_ASAP7_75t_L g1198 ( 
.A(n_1065),
.Y(n_1198)
);

NOR3xp33_ASAP7_75t_L g1199 ( 
.A(n_1080),
.B(n_858),
.C(n_749),
.Y(n_1199)
);

INVx4_ASAP7_75t_L g1200 ( 
.A(n_1076),
.Y(n_1200)
);

INVx3_ASAP7_75t_L g1201 ( 
.A(n_1041),
.Y(n_1201)
);

INVx1_ASAP7_75t_L g1202 ( 
.A(n_1068),
.Y(n_1202)
);

INVx2_ASAP7_75t_SL g1203 ( 
.A(n_1062),
.Y(n_1203)
);

NOR2xp67_ASAP7_75t_L g1204 ( 
.A(n_1119),
.B(n_805),
.Y(n_1204)
);

NAND2xp5_ASAP7_75t_SL g1205 ( 
.A(n_1152),
.B(n_567),
.Y(n_1205)
);

INVx2_ASAP7_75t_L g1206 ( 
.A(n_1068),
.Y(n_1206)
);

NAND2xp5_ASAP7_75t_L g1207 ( 
.A(n_1073),
.B(n_1074),
.Y(n_1207)
);

INVx1_ASAP7_75t_L g1208 ( 
.A(n_1074),
.Y(n_1208)
);

BUFx6f_ASAP7_75t_L g1209 ( 
.A(n_1076),
.Y(n_1209)
);

NAND2xp5_ASAP7_75t_L g1210 ( 
.A(n_1047),
.B(n_889),
.Y(n_1210)
);

NAND2xp5_ASAP7_75t_L g1211 ( 
.A(n_1122),
.B(n_836),
.Y(n_1211)
);

INVx1_ASAP7_75t_L g1212 ( 
.A(n_1079),
.Y(n_1212)
);

INVx2_ASAP7_75t_SL g1213 ( 
.A(n_1062),
.Y(n_1213)
);

NAND2xp5_ASAP7_75t_L g1214 ( 
.A(n_1122),
.B(n_836),
.Y(n_1214)
);

NAND2xp5_ASAP7_75t_L g1215 ( 
.A(n_1134),
.B(n_836),
.Y(n_1215)
);

BUFx6f_ASAP7_75t_L g1216 ( 
.A(n_1076),
.Y(n_1216)
);

INVx1_ASAP7_75t_L g1217 ( 
.A(n_1079),
.Y(n_1217)
);

INVx1_ASAP7_75t_SL g1218 ( 
.A(n_1104),
.Y(n_1218)
);

NAND2xp5_ASAP7_75t_L g1219 ( 
.A(n_1063),
.B(n_836),
.Y(n_1219)
);

AOI221xp5_ASAP7_75t_L g1220 ( 
.A1(n_1034),
.A2(n_580),
.B1(n_590),
.B2(n_578),
.C(n_575),
.Y(n_1220)
);

INVx1_ASAP7_75t_L g1221 ( 
.A(n_1090),
.Y(n_1221)
);

INVx8_ASAP7_75t_L g1222 ( 
.A(n_1093),
.Y(n_1222)
);

NAND2xp33_ASAP7_75t_L g1223 ( 
.A(n_1103),
.B(n_709),
.Y(n_1223)
);

NAND2xp5_ASAP7_75t_SL g1224 ( 
.A(n_1152),
.B(n_569),
.Y(n_1224)
);

NOR2xp33_ASAP7_75t_L g1225 ( 
.A(n_1080),
.B(n_868),
.Y(n_1225)
);

NOR3xp33_ASAP7_75t_L g1226 ( 
.A(n_1034),
.B(n_811),
.C(n_806),
.Y(n_1226)
);

NAND2xp5_ASAP7_75t_L g1227 ( 
.A(n_1107),
.B(n_836),
.Y(n_1227)
);

NOR2xp33_ASAP7_75t_L g1228 ( 
.A(n_1117),
.B(n_872),
.Y(n_1228)
);

BUFx6f_ASAP7_75t_SL g1229 ( 
.A(n_1089),
.Y(n_1229)
);

NAND2xp5_ASAP7_75t_L g1230 ( 
.A(n_1107),
.B(n_836),
.Y(n_1230)
);

INVx1_ASAP7_75t_L g1231 ( 
.A(n_1090),
.Y(n_1231)
);

CKINVDCx20_ASAP7_75t_R g1232 ( 
.A(n_1100),
.Y(n_1232)
);

NAND2xp5_ASAP7_75t_L g1233 ( 
.A(n_1041),
.B(n_845),
.Y(n_1233)
);

NOR2xp33_ASAP7_75t_L g1234 ( 
.A(n_1066),
.B(n_872),
.Y(n_1234)
);

INVx2_ASAP7_75t_L g1235 ( 
.A(n_1135),
.Y(n_1235)
);

NAND3xp33_ASAP7_75t_L g1236 ( 
.A(n_1109),
.B(n_843),
.C(n_597),
.Y(n_1236)
);

AOI221xp5_ASAP7_75t_L g1237 ( 
.A1(n_1146),
.A2(n_873),
.B1(n_772),
.B2(n_573),
.C(n_583),
.Y(n_1237)
);

NAND2xp5_ASAP7_75t_L g1238 ( 
.A(n_1071),
.B(n_845),
.Y(n_1238)
);

INVxp67_ASAP7_75t_SL g1239 ( 
.A(n_1103),
.Y(n_1239)
);

NOR2xp33_ASAP7_75t_L g1240 ( 
.A(n_1139),
.B(n_576),
.Y(n_1240)
);

INVx3_ASAP7_75t_L g1241 ( 
.A(n_1071),
.Y(n_1241)
);

INVx2_ASAP7_75t_L g1242 ( 
.A(n_1092),
.Y(n_1242)
);

NAND2xp5_ASAP7_75t_SL g1243 ( 
.A(n_1114),
.B(n_576),
.Y(n_1243)
);

NAND2xp5_ASAP7_75t_L g1244 ( 
.A(n_1092),
.B(n_845),
.Y(n_1244)
);

NAND2xp5_ASAP7_75t_L g1245 ( 
.A(n_1106),
.B(n_845),
.Y(n_1245)
);

BUFx3_ASAP7_75t_L g1246 ( 
.A(n_1121),
.Y(n_1246)
);

NAND2xp5_ASAP7_75t_L g1247 ( 
.A(n_1106),
.B(n_845),
.Y(n_1247)
);

NAND2xp5_ASAP7_75t_L g1248 ( 
.A(n_1112),
.B(n_882),
.Y(n_1248)
);

NAND2xp5_ASAP7_75t_L g1249 ( 
.A(n_1070),
.B(n_882),
.Y(n_1249)
);

CKINVDCx5p33_ASAP7_75t_R g1250 ( 
.A(n_1055),
.Y(n_1250)
);

BUFx6f_ASAP7_75t_L g1251 ( 
.A(n_1103),
.Y(n_1251)
);

NAND2xp5_ASAP7_75t_SL g1252 ( 
.A(n_1070),
.B(n_561),
.Y(n_1252)
);

NAND3xp33_ASAP7_75t_L g1253 ( 
.A(n_1059),
.B(n_600),
.C(n_596),
.Y(n_1253)
);

NAND2xp5_ASAP7_75t_L g1254 ( 
.A(n_1078),
.B(n_882),
.Y(n_1254)
);

INVx2_ASAP7_75t_SL g1255 ( 
.A(n_1121),
.Y(n_1255)
);

AND2x2_ASAP7_75t_L g1256 ( 
.A(n_1147),
.B(n_814),
.Y(n_1256)
);

OR2x6_ASAP7_75t_L g1257 ( 
.A(n_1093),
.B(n_683),
.Y(n_1257)
);

INVx2_ASAP7_75t_L g1258 ( 
.A(n_1120),
.Y(n_1258)
);

INVx2_ASAP7_75t_SL g1259 ( 
.A(n_1059),
.Y(n_1259)
);

INVx2_ASAP7_75t_SL g1260 ( 
.A(n_1153),
.Y(n_1260)
);

NOR2xp33_ASAP7_75t_L g1261 ( 
.A(n_1056),
.B(n_601),
.Y(n_1261)
);

NAND2xp5_ASAP7_75t_L g1262 ( 
.A(n_1124),
.B(n_882),
.Y(n_1262)
);

NAND2xp5_ASAP7_75t_L g1263 ( 
.A(n_1124),
.B(n_882),
.Y(n_1263)
);

INVx1_ASAP7_75t_L g1264 ( 
.A(n_1035),
.Y(n_1264)
);

AND2x2_ASAP7_75t_SL g1265 ( 
.A(n_1138),
.B(n_669),
.Y(n_1265)
);

NAND2xp5_ASAP7_75t_SL g1266 ( 
.A(n_1056),
.B(n_586),
.Y(n_1266)
);

INVx1_ASAP7_75t_L g1267 ( 
.A(n_1035),
.Y(n_1267)
);

INVx3_ASAP7_75t_L g1268 ( 
.A(n_1113),
.Y(n_1268)
);

NAND2xp5_ASAP7_75t_L g1269 ( 
.A(n_1098),
.B(n_813),
.Y(n_1269)
);

NAND2xp5_ASAP7_75t_L g1270 ( 
.A(n_1099),
.B(n_1102),
.Y(n_1270)
);

NAND2xp5_ASAP7_75t_SL g1271 ( 
.A(n_1128),
.B(n_591),
.Y(n_1271)
);

NAND2xp5_ASAP7_75t_SL g1272 ( 
.A(n_1103),
.B(n_592),
.Y(n_1272)
);

NAND2xp5_ASAP7_75t_L g1273 ( 
.A(n_1105),
.B(n_904),
.Y(n_1273)
);

NAND2xp5_ASAP7_75t_SL g1274 ( 
.A(n_1127),
.B(n_593),
.Y(n_1274)
);

INVx1_ASAP7_75t_L g1275 ( 
.A(n_1037),
.Y(n_1275)
);

NAND2xp5_ASAP7_75t_L g1276 ( 
.A(n_1108),
.B(n_904),
.Y(n_1276)
);

NAND2xp5_ASAP7_75t_L g1277 ( 
.A(n_1110),
.B(n_910),
.Y(n_1277)
);

NAND2xp5_ASAP7_75t_L g1278 ( 
.A(n_1038),
.B(n_910),
.Y(n_1278)
);

XOR2xp5_ASAP7_75t_L g1279 ( 
.A(n_1153),
.B(n_598),
.Y(n_1279)
);

AOI22xp5_ASAP7_75t_L g1280 ( 
.A1(n_1042),
.A2(n_603),
.B1(n_604),
.B2(n_599),
.Y(n_1280)
);

NOR2xp33_ASAP7_75t_L g1281 ( 
.A(n_1042),
.B(n_602),
.Y(n_1281)
);

INVx2_ASAP7_75t_L g1282 ( 
.A(n_1143),
.Y(n_1282)
);

NAND2xp5_ASAP7_75t_L g1283 ( 
.A(n_1086),
.B(n_916),
.Y(n_1283)
);

NOR3xp33_ASAP7_75t_L g1284 ( 
.A(n_1146),
.B(n_816),
.C(n_815),
.Y(n_1284)
);

NAND2xp5_ASAP7_75t_SL g1285 ( 
.A(n_1127),
.B(n_608),
.Y(n_1285)
);

NAND2xp5_ASAP7_75t_L g1286 ( 
.A(n_1087),
.B(n_916),
.Y(n_1286)
);

NOR2xp67_ASAP7_75t_L g1287 ( 
.A(n_1149),
.B(n_817),
.Y(n_1287)
);

NAND2xp33_ASAP7_75t_L g1288 ( 
.A(n_1127),
.B(n_709),
.Y(n_1288)
);

NAND2xp5_ASAP7_75t_L g1289 ( 
.A(n_1054),
.B(n_917),
.Y(n_1289)
);

INVx2_ASAP7_75t_L g1290 ( 
.A(n_1144),
.Y(n_1290)
);

NAND2xp5_ASAP7_75t_L g1291 ( 
.A(n_1118),
.B(n_917),
.Y(n_1291)
);

NAND2xp5_ASAP7_75t_SL g1292 ( 
.A(n_1088),
.B(n_611),
.Y(n_1292)
);

BUFx8_ASAP7_75t_L g1293 ( 
.A(n_1055),
.Y(n_1293)
);

NOR2xp33_ASAP7_75t_SL g1294 ( 
.A(n_1072),
.B(n_621),
.Y(n_1294)
);

AND2x4_ASAP7_75t_L g1295 ( 
.A(n_1084),
.B(n_861),
.Y(n_1295)
);

INVxp33_ASAP7_75t_L g1296 ( 
.A(n_1116),
.Y(n_1296)
);

INVx1_ASAP7_75t_L g1297 ( 
.A(n_1145),
.Y(n_1297)
);

AO221x1_ASAP7_75t_L g1298 ( 
.A1(n_1157),
.A2(n_641),
.B1(n_659),
.B2(n_657),
.C(n_646),
.Y(n_1298)
);

NOR2xp33_ASAP7_75t_L g1299 ( 
.A(n_1069),
.B(n_607),
.Y(n_1299)
);

NAND2xp5_ASAP7_75t_L g1300 ( 
.A(n_1069),
.B(n_922),
.Y(n_1300)
);

NAND3xp33_ASAP7_75t_SL g1301 ( 
.A(n_1123),
.B(n_583),
.C(n_579),
.Y(n_1301)
);

INVx2_ASAP7_75t_SL g1302 ( 
.A(n_1072),
.Y(n_1302)
);

AND2x2_ASAP7_75t_L g1303 ( 
.A(n_1111),
.B(n_818),
.Y(n_1303)
);

INVx1_ASAP7_75t_L g1304 ( 
.A(n_1125),
.Y(n_1304)
);

INVx1_ASAP7_75t_L g1305 ( 
.A(n_1133),
.Y(n_1305)
);

AND2x2_ASAP7_75t_L g1306 ( 
.A(n_1094),
.B(n_819),
.Y(n_1306)
);

INVx1_ASAP7_75t_L g1307 ( 
.A(n_1137),
.Y(n_1307)
);

INVx1_ASAP7_75t_L g1308 ( 
.A(n_1140),
.Y(n_1308)
);

INVx1_ASAP7_75t_L g1309 ( 
.A(n_1141),
.Y(n_1309)
);

NAND2xp5_ASAP7_75t_SL g1310 ( 
.A(n_1085),
.B(n_629),
.Y(n_1310)
);

NAND2xp5_ASAP7_75t_L g1311 ( 
.A(n_1151),
.B(n_922),
.Y(n_1311)
);

NAND2xp5_ASAP7_75t_L g1312 ( 
.A(n_1155),
.B(n_931),
.Y(n_1312)
);

INVx2_ASAP7_75t_SL g1313 ( 
.A(n_1101),
.Y(n_1313)
);

NAND3xp33_ASAP7_75t_L g1314 ( 
.A(n_1115),
.B(n_615),
.C(n_613),
.Y(n_1314)
);

NAND2xp5_ASAP7_75t_L g1315 ( 
.A(n_1155),
.B(n_935),
.Y(n_1315)
);

INVx1_ASAP7_75t_L g1316 ( 
.A(n_1154),
.Y(n_1316)
);

NAND2xp5_ASAP7_75t_L g1317 ( 
.A(n_1091),
.B(n_826),
.Y(n_1317)
);

INVxp67_ASAP7_75t_L g1318 ( 
.A(n_1129),
.Y(n_1318)
);

NAND2xp5_ASAP7_75t_SL g1319 ( 
.A(n_1085),
.B(n_635),
.Y(n_1319)
);

INVx1_ASAP7_75t_L g1320 ( 
.A(n_1156),
.Y(n_1320)
);

INVx2_ASAP7_75t_SL g1321 ( 
.A(n_1101),
.Y(n_1321)
);

INVx2_ASAP7_75t_L g1322 ( 
.A(n_1148),
.Y(n_1322)
);

INVx1_ASAP7_75t_L g1323 ( 
.A(n_1158),
.Y(n_1323)
);

NAND2xp5_ASAP7_75t_SL g1324 ( 
.A(n_1085),
.B(n_636),
.Y(n_1324)
);

HB1xp67_ASAP7_75t_L g1325 ( 
.A(n_1162),
.Y(n_1325)
);

INVx1_ASAP7_75t_L g1326 ( 
.A(n_1159),
.Y(n_1326)
);

NOR2xp67_ASAP7_75t_L g1327 ( 
.A(n_1236),
.B(n_1129),
.Y(n_1327)
);

BUFx3_ASAP7_75t_L g1328 ( 
.A(n_1182),
.Y(n_1328)
);

AO22x2_ASAP7_75t_L g1329 ( 
.A1(n_1266),
.A2(n_683),
.B1(n_722),
.B2(n_670),
.Y(n_1329)
);

AND2x2_ASAP7_75t_L g1330 ( 
.A(n_1225),
.B(n_1228),
.Y(n_1330)
);

NOR2xp67_ASAP7_75t_L g1331 ( 
.A(n_1250),
.B(n_1130),
.Y(n_1331)
);

INVx2_ASAP7_75t_L g1332 ( 
.A(n_1161),
.Y(n_1332)
);

AO22x2_ASAP7_75t_L g1333 ( 
.A1(n_1205),
.A2(n_726),
.B1(n_742),
.B2(n_722),
.Y(n_1333)
);

AO22x2_ASAP7_75t_L g1334 ( 
.A1(n_1224),
.A2(n_742),
.B1(n_758),
.B2(n_726),
.Y(n_1334)
);

INVx3_ASAP7_75t_L g1335 ( 
.A(n_1246),
.Y(n_1335)
);

NAND2x1p5_ASAP7_75t_L g1336 ( 
.A(n_1218),
.B(n_1049),
.Y(n_1336)
);

AND2x2_ASAP7_75t_L g1337 ( 
.A(n_1256),
.B(n_865),
.Y(n_1337)
);

INVx1_ASAP7_75t_L g1338 ( 
.A(n_1171),
.Y(n_1338)
);

AND2x4_ASAP7_75t_L g1339 ( 
.A(n_1175),
.B(n_1113),
.Y(n_1339)
);

INVx1_ASAP7_75t_L g1340 ( 
.A(n_1179),
.Y(n_1340)
);

INVx2_ASAP7_75t_SL g1341 ( 
.A(n_1162),
.Y(n_1341)
);

INVx1_ASAP7_75t_L g1342 ( 
.A(n_1183),
.Y(n_1342)
);

AND2x2_ASAP7_75t_L g1343 ( 
.A(n_1265),
.B(n_866),
.Y(n_1343)
);

INVx1_ASAP7_75t_L g1344 ( 
.A(n_1185),
.Y(n_1344)
);

INVx1_ASAP7_75t_L g1345 ( 
.A(n_1186),
.Y(n_1345)
);

INVx2_ASAP7_75t_L g1346 ( 
.A(n_1172),
.Y(n_1346)
);

INVx2_ASAP7_75t_L g1347 ( 
.A(n_1181),
.Y(n_1347)
);

INVx1_ASAP7_75t_L g1348 ( 
.A(n_1202),
.Y(n_1348)
);

INVx1_ASAP7_75t_L g1349 ( 
.A(n_1208),
.Y(n_1349)
);

NAND3xp33_ASAP7_75t_SL g1350 ( 
.A(n_1177),
.B(n_672),
.C(n_579),
.Y(n_1350)
);

AO22x2_ASAP7_75t_L g1351 ( 
.A1(n_1259),
.A2(n_758),
.B1(n_690),
.B2(n_691),
.Y(n_1351)
);

OAI221xp5_ASAP7_75t_L g1352 ( 
.A1(n_1220),
.A2(n_773),
.B1(n_775),
.B2(n_772),
.C(n_672),
.Y(n_1352)
);

AND2x6_ASAP7_75t_SL g1353 ( 
.A(n_1169),
.B(n_661),
.Y(n_1353)
);

INVx2_ASAP7_75t_L g1354 ( 
.A(n_1189),
.Y(n_1354)
);

AND2x4_ASAP7_75t_L g1355 ( 
.A(n_1203),
.B(n_1131),
.Y(n_1355)
);

INVx2_ASAP7_75t_L g1356 ( 
.A(n_1195),
.Y(n_1356)
);

NAND2xp5_ASAP7_75t_L g1357 ( 
.A(n_1306),
.B(n_1136),
.Y(n_1357)
);

AOI22xp33_ASAP7_75t_L g1358 ( 
.A1(n_1261),
.A2(n_1130),
.B1(n_1126),
.B2(n_1095),
.Y(n_1358)
);

INVx1_ASAP7_75t_L g1359 ( 
.A(n_1212),
.Y(n_1359)
);

INVx2_ASAP7_75t_L g1360 ( 
.A(n_1197),
.Y(n_1360)
);

AND2x2_ASAP7_75t_L g1361 ( 
.A(n_1163),
.B(n_869),
.Y(n_1361)
);

INVx2_ASAP7_75t_L g1362 ( 
.A(n_1198),
.Y(n_1362)
);

INVx1_ASAP7_75t_L g1363 ( 
.A(n_1217),
.Y(n_1363)
);

INVxp67_ASAP7_75t_L g1364 ( 
.A(n_1218),
.Y(n_1364)
);

NOR2xp33_ASAP7_75t_SL g1365 ( 
.A(n_1232),
.B(n_773),
.Y(n_1365)
);

CKINVDCx16_ASAP7_75t_R g1366 ( 
.A(n_1168),
.Y(n_1366)
);

AO22x2_ASAP7_75t_L g1367 ( 
.A1(n_1199),
.A2(n_700),
.B1(n_702),
.B2(n_699),
.Y(n_1367)
);

INVx1_ASAP7_75t_L g1368 ( 
.A(n_1221),
.Y(n_1368)
);

INVx1_ASAP7_75t_L g1369 ( 
.A(n_1231),
.Y(n_1369)
);

AND2x2_ASAP7_75t_L g1370 ( 
.A(n_1234),
.B(n_874),
.Y(n_1370)
);

AND2x2_ASAP7_75t_L g1371 ( 
.A(n_1173),
.B(n_877),
.Y(n_1371)
);

AO22x2_ASAP7_75t_L g1372 ( 
.A1(n_1301),
.A2(n_708),
.B1(n_710),
.B2(n_706),
.Y(n_1372)
);

AOI22xp5_ASAP7_75t_L g1373 ( 
.A1(n_1176),
.A2(n_647),
.B1(n_648),
.B2(n_640),
.Y(n_1373)
);

AO22x2_ASAP7_75t_L g1374 ( 
.A1(n_1243),
.A2(n_718),
.B1(n_724),
.B2(n_711),
.Y(n_1374)
);

NAND2xp33_ASAP7_75t_L g1375 ( 
.A(n_1192),
.B(n_1209),
.Y(n_1375)
);

NAND2x1p5_ASAP7_75t_L g1376 ( 
.A(n_1213),
.B(n_1053),
.Y(n_1376)
);

INVxp67_ASAP7_75t_L g1377 ( 
.A(n_1170),
.Y(n_1377)
);

AO22x2_ASAP7_75t_L g1378 ( 
.A1(n_1226),
.A2(n_747),
.B1(n_751),
.B2(n_730),
.Y(n_1378)
);

AO22x2_ASAP7_75t_L g1379 ( 
.A1(n_1313),
.A2(n_756),
.B1(n_761),
.B2(n_753),
.Y(n_1379)
);

INVx1_ASAP7_75t_L g1380 ( 
.A(n_1206),
.Y(n_1380)
);

AOI22xp5_ASAP7_75t_L g1381 ( 
.A1(n_1299),
.A2(n_664),
.B1(n_671),
.B2(n_654),
.Y(n_1381)
);

NAND2x1p5_ASAP7_75t_L g1382 ( 
.A(n_1200),
.B(n_1081),
.Y(n_1382)
);

BUFx3_ASAP7_75t_L g1383 ( 
.A(n_1255),
.Y(n_1383)
);

BUFx8_ASAP7_75t_L g1384 ( 
.A(n_1168),
.Y(n_1384)
);

INVx1_ASAP7_75t_L g1385 ( 
.A(n_1242),
.Y(n_1385)
);

BUFx6f_ASAP7_75t_L g1386 ( 
.A(n_1180),
.Y(n_1386)
);

INVxp67_ASAP7_75t_L g1387 ( 
.A(n_1240),
.Y(n_1387)
);

INVx1_ASAP7_75t_L g1388 ( 
.A(n_1258),
.Y(n_1388)
);

AO22x2_ASAP7_75t_L g1389 ( 
.A1(n_1321),
.A2(n_776),
.B1(n_765),
.B2(n_878),
.Y(n_1389)
);

INVx1_ASAP7_75t_L g1390 ( 
.A(n_1264),
.Y(n_1390)
);

INVx1_ASAP7_75t_L g1391 ( 
.A(n_1267),
.Y(n_1391)
);

NAND2xp33_ASAP7_75t_R g1392 ( 
.A(n_1281),
.B(n_676),
.Y(n_1392)
);

AO22x2_ASAP7_75t_L g1393 ( 
.A1(n_1167),
.A2(n_879),
.B1(n_2),
.B2(n_0),
.Y(n_1393)
);

NAND2xp5_ASAP7_75t_SL g1394 ( 
.A(n_1294),
.B(n_1085),
.Y(n_1394)
);

NAND2xp5_ASAP7_75t_L g1395 ( 
.A(n_1270),
.B(n_1126),
.Y(n_1395)
);

NAND2xp5_ASAP7_75t_L g1396 ( 
.A(n_1270),
.B(n_684),
.Y(n_1396)
);

AOI22xp5_ASAP7_75t_L g1397 ( 
.A1(n_1160),
.A2(n_697),
.B1(n_720),
.B2(n_696),
.Y(n_1397)
);

AO22x2_ASAP7_75t_L g1398 ( 
.A1(n_1279),
.A2(n_1253),
.B1(n_1174),
.B2(n_1166),
.Y(n_1398)
);

AO22x2_ASAP7_75t_L g1399 ( 
.A1(n_1166),
.A2(n_3),
.B1(n_1),
.B2(n_2),
.Y(n_1399)
);

INVx2_ASAP7_75t_L g1400 ( 
.A(n_1282),
.Y(n_1400)
);

INVx1_ASAP7_75t_L g1401 ( 
.A(n_1275),
.Y(n_1401)
);

AO22x2_ASAP7_75t_L g1402 ( 
.A1(n_1174),
.A2(n_4),
.B1(n_1),
.B2(n_3),
.Y(n_1402)
);

INVx1_ASAP7_75t_L g1403 ( 
.A(n_1297),
.Y(n_1403)
);

INVx1_ASAP7_75t_L g1404 ( 
.A(n_1278),
.Y(n_1404)
);

INVx1_ASAP7_75t_L g1405 ( 
.A(n_1278),
.Y(n_1405)
);

INVx1_ASAP7_75t_L g1406 ( 
.A(n_1311),
.Y(n_1406)
);

NAND2x1p5_ASAP7_75t_L g1407 ( 
.A(n_1200),
.B(n_927),
.Y(n_1407)
);

CKINVDCx16_ASAP7_75t_R g1408 ( 
.A(n_1229),
.Y(n_1408)
);

NAND2xp5_ASAP7_75t_SL g1409 ( 
.A(n_1294),
.B(n_727),
.Y(n_1409)
);

AO22x2_ASAP7_75t_L g1410 ( 
.A1(n_1260),
.A2(n_1271),
.B1(n_1165),
.B2(n_1298),
.Y(n_1410)
);

INVx1_ASAP7_75t_L g1411 ( 
.A(n_1311),
.Y(n_1411)
);

AOI22xp5_ASAP7_75t_L g1412 ( 
.A1(n_1296),
.A2(n_740),
.B1(n_743),
.B2(n_733),
.Y(n_1412)
);

INVx1_ASAP7_75t_L g1413 ( 
.A(n_1312),
.Y(n_1413)
);

BUFx3_ASAP7_75t_L g1414 ( 
.A(n_1293),
.Y(n_1414)
);

AND2x4_ASAP7_75t_L g1415 ( 
.A(n_1180),
.B(n_375),
.Y(n_1415)
);

INVx1_ASAP7_75t_L g1416 ( 
.A(n_1312),
.Y(n_1416)
);

INVx2_ASAP7_75t_L g1417 ( 
.A(n_1290),
.Y(n_1417)
);

INVx1_ASAP7_75t_L g1418 ( 
.A(n_1315),
.Y(n_1418)
);

INVx1_ASAP7_75t_L g1419 ( 
.A(n_1315),
.Y(n_1419)
);

AO22x2_ASAP7_75t_L g1420 ( 
.A1(n_1187),
.A2(n_7),
.B1(n_5),
.B2(n_6),
.Y(n_1420)
);

INVx1_ASAP7_75t_L g1421 ( 
.A(n_1235),
.Y(n_1421)
);

NAND2x1p5_ASAP7_75t_L g1422 ( 
.A(n_1209),
.B(n_927),
.Y(n_1422)
);

OAI22xp5_ASAP7_75t_L g1423 ( 
.A1(n_1207),
.A2(n_750),
.B1(n_763),
.B2(n_745),
.Y(n_1423)
);

AO22x2_ASAP7_75t_L g1424 ( 
.A1(n_1211),
.A2(n_1214),
.B1(n_1305),
.B2(n_1304),
.Y(n_1424)
);

NOR2xp33_ASAP7_75t_L g1425 ( 
.A(n_1193),
.B(n_620),
.Y(n_1425)
);

NAND2xp5_ASAP7_75t_L g1426 ( 
.A(n_1194),
.B(n_764),
.Y(n_1426)
);

AO22x2_ASAP7_75t_L g1427 ( 
.A1(n_1307),
.A2(n_7),
.B1(n_5),
.B2(n_6),
.Y(n_1427)
);

AO22x2_ASAP7_75t_L g1428 ( 
.A1(n_1308),
.A2(n_10),
.B1(n_8),
.B2(n_9),
.Y(n_1428)
);

NAND2xp5_ASAP7_75t_L g1429 ( 
.A(n_1196),
.B(n_622),
.Y(n_1429)
);

INVx1_ASAP7_75t_L g1430 ( 
.A(n_1309),
.Y(n_1430)
);

INVx2_ASAP7_75t_SL g1431 ( 
.A(n_1295),
.Y(n_1431)
);

NAND2xp5_ASAP7_75t_L g1432 ( 
.A(n_1210),
.B(n_623),
.Y(n_1432)
);

NAND2xp5_ASAP7_75t_SL g1433 ( 
.A(n_1192),
.B(n_927),
.Y(n_1433)
);

AO22x2_ASAP7_75t_L g1434 ( 
.A1(n_1316),
.A2(n_11),
.B1(n_8),
.B2(n_9),
.Y(n_1434)
);

AO22x2_ASAP7_75t_L g1435 ( 
.A1(n_1178),
.A2(n_14),
.B1(n_11),
.B2(n_12),
.Y(n_1435)
);

AOI22xp5_ASAP7_75t_L g1436 ( 
.A1(n_1314),
.A2(n_936),
.B1(n_943),
.B2(n_912),
.Y(n_1436)
);

INVx1_ASAP7_75t_L g1437 ( 
.A(n_1291),
.Y(n_1437)
);

AO22x2_ASAP7_75t_L g1438 ( 
.A1(n_1178),
.A2(n_17),
.B1(n_15),
.B2(n_16),
.Y(n_1438)
);

AND2x4_ASAP7_75t_L g1439 ( 
.A(n_1180),
.B(n_376),
.Y(n_1439)
);

INVx1_ASAP7_75t_L g1440 ( 
.A(n_1273),
.Y(n_1440)
);

NAND2xp5_ASAP7_75t_L g1441 ( 
.A(n_1188),
.B(n_631),
.Y(n_1441)
);

CKINVDCx5p33_ASAP7_75t_R g1442 ( 
.A(n_1293),
.Y(n_1442)
);

INVx1_ASAP7_75t_L g1443 ( 
.A(n_1276),
.Y(n_1443)
);

AO22x2_ASAP7_75t_L g1444 ( 
.A1(n_1284),
.A2(n_1323),
.B1(n_1320),
.B2(n_1322),
.Y(n_1444)
);

AOI22xp5_ASAP7_75t_L g1445 ( 
.A1(n_1252),
.A2(n_936),
.B1(n_943),
.B2(n_912),
.Y(n_1445)
);

INVx2_ASAP7_75t_L g1446 ( 
.A(n_1268),
.Y(n_1446)
);

INVx1_ASAP7_75t_L g1447 ( 
.A(n_1277),
.Y(n_1447)
);

AO22x2_ASAP7_75t_L g1448 ( 
.A1(n_1302),
.A2(n_18),
.B1(n_15),
.B2(n_16),
.Y(n_1448)
);

INVx1_ASAP7_75t_L g1449 ( 
.A(n_1283),
.Y(n_1449)
);

BUFx8_ASAP7_75t_L g1450 ( 
.A(n_1229),
.Y(n_1450)
);

AND2x4_ASAP7_75t_L g1451 ( 
.A(n_1295),
.B(n_377),
.Y(n_1451)
);

AO22x2_ASAP7_75t_L g1452 ( 
.A1(n_1191),
.A2(n_21),
.B1(n_19),
.B2(n_20),
.Y(n_1452)
);

NAND2xp5_ASAP7_75t_L g1453 ( 
.A(n_1192),
.B(n_632),
.Y(n_1453)
);

AO22x2_ASAP7_75t_L g1454 ( 
.A1(n_1318),
.A2(n_21),
.B1(n_19),
.B2(n_20),
.Y(n_1454)
);

NAND2xp5_ASAP7_75t_L g1455 ( 
.A(n_1192),
.B(n_1201),
.Y(n_1455)
);

AOI22xp5_ASAP7_75t_L g1456 ( 
.A1(n_1292),
.A2(n_936),
.B1(n_943),
.B2(n_912),
.Y(n_1456)
);

AO22x2_ASAP7_75t_L g1457 ( 
.A1(n_1227),
.A2(n_24),
.B1(n_22),
.B2(n_23),
.Y(n_1457)
);

AO22x2_ASAP7_75t_L g1458 ( 
.A1(n_1227),
.A2(n_25),
.B1(n_23),
.B2(n_24),
.Y(n_1458)
);

AO22x2_ASAP7_75t_L g1459 ( 
.A1(n_1230),
.A2(n_27),
.B1(n_25),
.B2(n_26),
.Y(n_1459)
);

NAND2x1p5_ASAP7_75t_L g1460 ( 
.A(n_1209),
.B(n_927),
.Y(n_1460)
);

CKINVDCx20_ASAP7_75t_R g1461 ( 
.A(n_1190),
.Y(n_1461)
);

BUFx6f_ASAP7_75t_L g1462 ( 
.A(n_1222),
.Y(n_1462)
);

BUFx2_ASAP7_75t_L g1463 ( 
.A(n_1216),
.Y(n_1463)
);

CKINVDCx11_ASAP7_75t_R g1464 ( 
.A(n_1222),
.Y(n_1464)
);

NAND2xp5_ASAP7_75t_L g1465 ( 
.A(n_1201),
.B(n_633),
.Y(n_1465)
);

NAND2x1_ASAP7_75t_L g1466 ( 
.A(n_1268),
.B(n_946),
.Y(n_1466)
);

NAND2x1p5_ASAP7_75t_L g1467 ( 
.A(n_1216),
.B(n_940),
.Y(n_1467)
);

INVx1_ASAP7_75t_L g1468 ( 
.A(n_1286),
.Y(n_1468)
);

NAND2x1p5_ASAP7_75t_L g1469 ( 
.A(n_1216),
.B(n_940),
.Y(n_1469)
);

INVx1_ASAP7_75t_L g1470 ( 
.A(n_1269),
.Y(n_1470)
);

INVx1_ASAP7_75t_L g1471 ( 
.A(n_1300),
.Y(n_1471)
);

AO22x2_ASAP7_75t_L g1472 ( 
.A1(n_1230),
.A2(n_28),
.B1(n_26),
.B2(n_27),
.Y(n_1472)
);

INVx3_ASAP7_75t_L g1473 ( 
.A(n_1222),
.Y(n_1473)
);

CKINVDCx5p33_ASAP7_75t_R g1474 ( 
.A(n_1257),
.Y(n_1474)
);

NAND2x1p5_ASAP7_75t_L g1475 ( 
.A(n_1251),
.B(n_1241),
.Y(n_1475)
);

INVx1_ASAP7_75t_L g1476 ( 
.A(n_1300),
.Y(n_1476)
);

OAI221xp5_ASAP7_75t_L g1477 ( 
.A1(n_1237),
.A2(n_775),
.B1(n_645),
.B2(n_650),
.C(n_644),
.Y(n_1477)
);

OAI221xp5_ASAP7_75t_L g1478 ( 
.A1(n_1280),
.A2(n_655),
.B1(n_658),
.B2(n_652),
.C(n_642),
.Y(n_1478)
);

INVx1_ASAP7_75t_L g1479 ( 
.A(n_1289),
.Y(n_1479)
);

INVx1_ASAP7_75t_L g1480 ( 
.A(n_1289),
.Y(n_1480)
);

INVx2_ASAP7_75t_L g1481 ( 
.A(n_1241),
.Y(n_1481)
);

INVx2_ASAP7_75t_SL g1482 ( 
.A(n_1303),
.Y(n_1482)
);

INVx2_ASAP7_75t_L g1483 ( 
.A(n_1248),
.Y(n_1483)
);

INVxp67_ASAP7_75t_L g1484 ( 
.A(n_1257),
.Y(n_1484)
);

INVx1_ASAP7_75t_L g1485 ( 
.A(n_1244),
.Y(n_1485)
);

AOI22xp5_ASAP7_75t_L g1486 ( 
.A1(n_1204),
.A2(n_1285),
.B1(n_1272),
.B2(n_1274),
.Y(n_1486)
);

INVx1_ASAP7_75t_L g1487 ( 
.A(n_1244),
.Y(n_1487)
);

AO22x2_ASAP7_75t_L g1488 ( 
.A1(n_1184),
.A2(n_31),
.B1(n_28),
.B2(n_30),
.Y(n_1488)
);

INVx2_ASAP7_75t_L g1489 ( 
.A(n_1248),
.Y(n_1489)
);

INVx1_ASAP7_75t_L g1490 ( 
.A(n_1245),
.Y(n_1490)
);

AOI22xp5_ASAP7_75t_L g1491 ( 
.A1(n_1249),
.A2(n_943),
.B1(n_944),
.B2(n_936),
.Y(n_1491)
);

OAI22xp5_ASAP7_75t_L g1492 ( 
.A1(n_1215),
.A2(n_678),
.B1(n_679),
.B2(n_673),
.Y(n_1492)
);

INVx1_ASAP7_75t_L g1493 ( 
.A(n_1245),
.Y(n_1493)
);

INVx1_ASAP7_75t_L g1494 ( 
.A(n_1247),
.Y(n_1494)
);

OR2x2_ASAP7_75t_SL g1495 ( 
.A(n_1257),
.B(n_685),
.Y(n_1495)
);

INVx1_ASAP7_75t_L g1496 ( 
.A(n_1287),
.Y(n_1496)
);

NAND2xp5_ASAP7_75t_L g1497 ( 
.A(n_1219),
.B(n_687),
.Y(n_1497)
);

NAND2xp5_ASAP7_75t_L g1498 ( 
.A(n_1330),
.B(n_1219),
.Y(n_1498)
);

NAND2xp5_ASAP7_75t_L g1499 ( 
.A(n_1449),
.B(n_1317),
.Y(n_1499)
);

BUFx2_ASAP7_75t_L g1500 ( 
.A(n_1325),
.Y(n_1500)
);

NAND2xp5_ASAP7_75t_SL g1501 ( 
.A(n_1387),
.B(n_1254),
.Y(n_1501)
);

INVx2_ASAP7_75t_L g1502 ( 
.A(n_1430),
.Y(n_1502)
);

NAND2xp5_ASAP7_75t_L g1503 ( 
.A(n_1468),
.B(n_1233),
.Y(n_1503)
);

NAND2xp5_ASAP7_75t_L g1504 ( 
.A(n_1440),
.B(n_1233),
.Y(n_1504)
);

NAND2xp5_ASAP7_75t_L g1505 ( 
.A(n_1443),
.B(n_1238),
.Y(n_1505)
);

AND2x2_ASAP7_75t_L g1506 ( 
.A(n_1371),
.B(n_1164),
.Y(n_1506)
);

HB1xp67_ASAP7_75t_L g1507 ( 
.A(n_1341),
.Y(n_1507)
);

AND2x4_ASAP7_75t_L g1508 ( 
.A(n_1473),
.B(n_1239),
.Y(n_1508)
);

AOI21xp5_ASAP7_75t_L g1509 ( 
.A1(n_1375),
.A2(n_1319),
.B(n_1310),
.Y(n_1509)
);

NAND3xp33_ASAP7_75t_L g1510 ( 
.A(n_1425),
.B(n_1288),
.C(n_1223),
.Y(n_1510)
);

AND2x4_ASAP7_75t_L g1511 ( 
.A(n_1462),
.B(n_1431),
.Y(n_1511)
);

AOI21xp5_ASAP7_75t_L g1512 ( 
.A1(n_1395),
.A2(n_1324),
.B(n_1262),
.Y(n_1512)
);

NAND2xp5_ASAP7_75t_L g1513 ( 
.A(n_1447),
.B(n_1263),
.Y(n_1513)
);

AOI22xp5_ASAP7_75t_L g1514 ( 
.A1(n_1398),
.A2(n_1263),
.B1(n_689),
.B2(n_692),
.Y(n_1514)
);

INVx4_ASAP7_75t_L g1515 ( 
.A(n_1328),
.Y(n_1515)
);

AOI21xp5_ASAP7_75t_L g1516 ( 
.A1(n_1404),
.A2(n_1406),
.B(n_1405),
.Y(n_1516)
);

AOI21xp5_ASAP7_75t_L g1517 ( 
.A1(n_1411),
.A2(n_940),
.B(n_946),
.Y(n_1517)
);

OAI321xp33_ASAP7_75t_L g1518 ( 
.A1(n_1352),
.A2(n_854),
.A3(n_848),
.B1(n_857),
.B2(n_852),
.C(n_847),
.Y(n_1518)
);

NAND2xp5_ASAP7_75t_L g1519 ( 
.A(n_1437),
.B(n_688),
.Y(n_1519)
);

INVx1_ASAP7_75t_L g1520 ( 
.A(n_1390),
.Y(n_1520)
);

NOR2xp33_ASAP7_75t_L g1521 ( 
.A(n_1377),
.B(n_693),
.Y(n_1521)
);

NOR2xp33_ASAP7_75t_L g1522 ( 
.A(n_1364),
.B(n_694),
.Y(n_1522)
);

AOI21xp5_ASAP7_75t_L g1523 ( 
.A1(n_1413),
.A2(n_940),
.B(n_968),
.Y(n_1523)
);

A2O1A1Ixp33_ASAP7_75t_L g1524 ( 
.A1(n_1478),
.A2(n_698),
.B(n_703),
.C(n_695),
.Y(n_1524)
);

NAND2xp5_ASAP7_75t_L g1525 ( 
.A(n_1479),
.B(n_714),
.Y(n_1525)
);

AO21x1_ASAP7_75t_L g1526 ( 
.A1(n_1394),
.A2(n_31),
.B(n_32),
.Y(n_1526)
);

A2O1A1Ixp33_ASAP7_75t_L g1527 ( 
.A1(n_1327),
.A2(n_717),
.B(n_723),
.C(n_715),
.Y(n_1527)
);

AOI21xp5_ASAP7_75t_L g1528 ( 
.A1(n_1416),
.A2(n_968),
.B(n_944),
.Y(n_1528)
);

AOI21x1_ASAP7_75t_L g1529 ( 
.A1(n_1444),
.A2(n_944),
.B(n_968),
.Y(n_1529)
);

O2A1O1Ixp33_ASAP7_75t_L g1530 ( 
.A1(n_1350),
.A2(n_732),
.B(n_735),
.C(n_731),
.Y(n_1530)
);

AND2x2_ASAP7_75t_L g1531 ( 
.A(n_1343),
.B(n_737),
.Y(n_1531)
);

INVx1_ASAP7_75t_L g1532 ( 
.A(n_1391),
.Y(n_1532)
);

OAI21xp33_ASAP7_75t_L g1533 ( 
.A1(n_1367),
.A2(n_741),
.B(n_738),
.Y(n_1533)
);

NAND2xp5_ASAP7_75t_SL g1534 ( 
.A(n_1482),
.B(n_744),
.Y(n_1534)
);

NAND2xp5_ASAP7_75t_L g1535 ( 
.A(n_1480),
.B(n_746),
.Y(n_1535)
);

OAI21xp33_ASAP7_75t_L g1536 ( 
.A1(n_1367),
.A2(n_752),
.B(n_748),
.Y(n_1536)
);

O2A1O1Ixp33_ASAP7_75t_L g1537 ( 
.A1(n_1477),
.A2(n_759),
.B(n_762),
.C(n_754),
.Y(n_1537)
);

AOI21xp5_ASAP7_75t_L g1538 ( 
.A1(n_1418),
.A2(n_944),
.B(n_389),
.Y(n_1538)
);

AOI21xp33_ASAP7_75t_L g1539 ( 
.A1(n_1392),
.A2(n_768),
.B(n_766),
.Y(n_1539)
);

CKINVDCx8_ASAP7_75t_R g1540 ( 
.A(n_1366),
.Y(n_1540)
);

OAI21x1_ASAP7_75t_L g1541 ( 
.A1(n_1455),
.A2(n_390),
.B(n_383),
.Y(n_1541)
);

AND2x2_ASAP7_75t_L g1542 ( 
.A(n_1337),
.B(n_1370),
.Y(n_1542)
);

BUFx6f_ASAP7_75t_L g1543 ( 
.A(n_1462),
.Y(n_1543)
);

OAI22xp5_ASAP7_75t_L g1544 ( 
.A1(n_1419),
.A2(n_771),
.B1(n_777),
.B2(n_769),
.Y(n_1544)
);

NAND2xp5_ASAP7_75t_L g1545 ( 
.A(n_1471),
.B(n_32),
.Y(n_1545)
);

AOI22x1_ASAP7_75t_L g1546 ( 
.A1(n_1424),
.A2(n_944),
.B1(n_395),
.B2(n_396),
.Y(n_1546)
);

NAND2xp5_ASAP7_75t_L g1547 ( 
.A(n_1476),
.B(n_33),
.Y(n_1547)
);

A2O1A1Ixp33_ASAP7_75t_L g1548 ( 
.A1(n_1486),
.A2(n_36),
.B(n_34),
.C(n_35),
.Y(n_1548)
);

BUFx6f_ASAP7_75t_L g1549 ( 
.A(n_1464),
.Y(n_1549)
);

NOR2xp33_ASAP7_75t_L g1550 ( 
.A(n_1396),
.B(n_1365),
.Y(n_1550)
);

HB1xp67_ASAP7_75t_L g1551 ( 
.A(n_1335),
.Y(n_1551)
);

AND2x2_ASAP7_75t_L g1552 ( 
.A(n_1361),
.B(n_34),
.Y(n_1552)
);

OAI21xp33_ASAP7_75t_L g1553 ( 
.A1(n_1374),
.A2(n_36),
.B(n_37),
.Y(n_1553)
);

BUFx6f_ASAP7_75t_L g1554 ( 
.A(n_1386),
.Y(n_1554)
);

BUFx8_ASAP7_75t_SL g1555 ( 
.A(n_1461),
.Y(n_1555)
);

INVx2_ASAP7_75t_L g1556 ( 
.A(n_1400),
.Y(n_1556)
);

NOR3xp33_ASAP7_75t_L g1557 ( 
.A(n_1409),
.B(n_37),
.C(n_38),
.Y(n_1557)
);

AOI21xp5_ASAP7_75t_L g1558 ( 
.A1(n_1424),
.A2(n_397),
.B(n_391),
.Y(n_1558)
);

AND2x4_ASAP7_75t_L g1559 ( 
.A(n_1386),
.B(n_554),
.Y(n_1559)
);

INVx1_ASAP7_75t_L g1560 ( 
.A(n_1401),
.Y(n_1560)
);

AOI21xp5_ASAP7_75t_L g1561 ( 
.A1(n_1357),
.A2(n_399),
.B(n_398),
.Y(n_1561)
);

NAND2xp5_ASAP7_75t_SL g1562 ( 
.A(n_1383),
.B(n_38),
.Y(n_1562)
);

INVx2_ASAP7_75t_SL g1563 ( 
.A(n_1415),
.Y(n_1563)
);

INVx1_ASAP7_75t_L g1564 ( 
.A(n_1403),
.Y(n_1564)
);

OAI21x1_ASAP7_75t_L g1565 ( 
.A1(n_1433),
.A2(n_1483),
.B(n_1489),
.Y(n_1565)
);

OAI321xp33_ASAP7_75t_L g1566 ( 
.A1(n_1492),
.A2(n_41),
.A3(n_43),
.B1(n_39),
.B2(n_40),
.C(n_42),
.Y(n_1566)
);

NAND2xp5_ASAP7_75t_SL g1567 ( 
.A(n_1412),
.B(n_42),
.Y(n_1567)
);

AOI21xp5_ASAP7_75t_L g1568 ( 
.A1(n_1485),
.A2(n_1490),
.B(n_1487),
.Y(n_1568)
);

NAND2xp5_ASAP7_75t_L g1569 ( 
.A(n_1470),
.B(n_44),
.Y(n_1569)
);

NAND2xp5_ASAP7_75t_L g1570 ( 
.A(n_1493),
.B(n_45),
.Y(n_1570)
);

NAND2xp5_ASAP7_75t_L g1571 ( 
.A(n_1494),
.B(n_46),
.Y(n_1571)
);

AOI21xp5_ASAP7_75t_L g1572 ( 
.A1(n_1426),
.A2(n_403),
.B(n_402),
.Y(n_1572)
);

INVx2_ASAP7_75t_L g1573 ( 
.A(n_1417),
.Y(n_1573)
);

BUFx12f_ASAP7_75t_L g1574 ( 
.A(n_1450),
.Y(n_1574)
);

AOI21xp5_ASAP7_75t_L g1575 ( 
.A1(n_1358),
.A2(n_407),
.B(n_404),
.Y(n_1575)
);

AOI21x1_ASAP7_75t_L g1576 ( 
.A1(n_1453),
.A2(n_1441),
.B(n_1497),
.Y(n_1576)
);

NOR2xp33_ASAP7_75t_L g1577 ( 
.A(n_1429),
.B(n_46),
.Y(n_1577)
);

INVxp67_ASAP7_75t_L g1578 ( 
.A(n_1398),
.Y(n_1578)
);

NOR2xp33_ASAP7_75t_L g1579 ( 
.A(n_1432),
.B(n_47),
.Y(n_1579)
);

OAI22xp5_ASAP7_75t_L g1580 ( 
.A1(n_1326),
.A2(n_51),
.B1(n_48),
.B2(n_50),
.Y(n_1580)
);

INVx1_ASAP7_75t_L g1581 ( 
.A(n_1338),
.Y(n_1581)
);

OAI21xp5_ASAP7_75t_L g1582 ( 
.A1(n_1465),
.A2(n_410),
.B(n_408),
.Y(n_1582)
);

NAND2xp5_ASAP7_75t_L g1583 ( 
.A(n_1374),
.B(n_52),
.Y(n_1583)
);

OAI21xp33_ASAP7_75t_L g1584 ( 
.A1(n_1378),
.A2(n_52),
.B(n_53),
.Y(n_1584)
);

NAND2xp5_ASAP7_75t_L g1585 ( 
.A(n_1355),
.B(n_53),
.Y(n_1585)
);

AND2x4_ASAP7_75t_L g1586 ( 
.A(n_1415),
.B(n_411),
.Y(n_1586)
);

BUFx6f_ASAP7_75t_L g1587 ( 
.A(n_1463),
.Y(n_1587)
);

NAND2xp5_ASAP7_75t_L g1588 ( 
.A(n_1355),
.B(n_54),
.Y(n_1588)
);

AND2x6_ASAP7_75t_SL g1589 ( 
.A(n_1439),
.B(n_54),
.Y(n_1589)
);

AOI21xp5_ASAP7_75t_L g1590 ( 
.A1(n_1382),
.A2(n_414),
.B(n_413),
.Y(n_1590)
);

AOI21xp5_ASAP7_75t_L g1591 ( 
.A1(n_1466),
.A2(n_416),
.B(n_415),
.Y(n_1591)
);

INVx2_ASAP7_75t_SL g1592 ( 
.A(n_1439),
.Y(n_1592)
);

AOI21xp5_ASAP7_75t_L g1593 ( 
.A1(n_1340),
.A2(n_1344),
.B(n_1342),
.Y(n_1593)
);

BUFx3_ASAP7_75t_L g1594 ( 
.A(n_1384),
.Y(n_1594)
);

NAND2xp5_ASAP7_75t_L g1595 ( 
.A(n_1339),
.B(n_55),
.Y(n_1595)
);

BUFx12f_ASAP7_75t_L g1596 ( 
.A(n_1384),
.Y(n_1596)
);

NOR3xp33_ASAP7_75t_L g1597 ( 
.A(n_1484),
.B(n_56),
.C(n_57),
.Y(n_1597)
);

INVx2_ASAP7_75t_SL g1598 ( 
.A(n_1474),
.Y(n_1598)
);

O2A1O1Ixp33_ASAP7_75t_L g1599 ( 
.A1(n_1496),
.A2(n_58),
.B(n_56),
.C(n_57),
.Y(n_1599)
);

INVx2_ASAP7_75t_L g1600 ( 
.A(n_1345),
.Y(n_1600)
);

NOR2xp33_ASAP7_75t_SL g1601 ( 
.A(n_1442),
.B(n_417),
.Y(n_1601)
);

NAND2xp5_ASAP7_75t_L g1602 ( 
.A(n_1339),
.B(n_60),
.Y(n_1602)
);

NOR2xp33_ASAP7_75t_R g1603 ( 
.A(n_1408),
.B(n_419),
.Y(n_1603)
);

OAI21xp5_ASAP7_75t_L g1604 ( 
.A1(n_1380),
.A2(n_424),
.B(n_420),
.Y(n_1604)
);

INVx3_ASAP7_75t_L g1605 ( 
.A(n_1475),
.Y(n_1605)
);

INVx2_ASAP7_75t_L g1606 ( 
.A(n_1348),
.Y(n_1606)
);

AOI21xp5_ASAP7_75t_L g1607 ( 
.A1(n_1349),
.A2(n_428),
.B(n_426),
.Y(n_1607)
);

NAND2xp5_ASAP7_75t_L g1608 ( 
.A(n_1359),
.B(n_1363),
.Y(n_1608)
);

CKINVDCx20_ASAP7_75t_R g1609 ( 
.A(n_1414),
.Y(n_1609)
);

INVx2_ASAP7_75t_L g1610 ( 
.A(n_1368),
.Y(n_1610)
);

INVxp67_ASAP7_75t_L g1611 ( 
.A(n_1372),
.Y(n_1611)
);

BUFx6f_ASAP7_75t_L g1612 ( 
.A(n_1463),
.Y(n_1612)
);

AOI21xp5_ASAP7_75t_L g1613 ( 
.A1(n_1369),
.A2(n_431),
.B(n_429),
.Y(n_1613)
);

NAND2xp5_ASAP7_75t_L g1614 ( 
.A(n_1333),
.B(n_60),
.Y(n_1614)
);

NAND2x1p5_ASAP7_75t_L g1615 ( 
.A(n_1451),
.B(n_433),
.Y(n_1615)
);

AOI21x1_ASAP7_75t_L g1616 ( 
.A1(n_1333),
.A2(n_435),
.B(n_434),
.Y(n_1616)
);

NAND2xp5_ASAP7_75t_L g1617 ( 
.A(n_1334),
.B(n_61),
.Y(n_1617)
);

CKINVDCx5p33_ASAP7_75t_R g1618 ( 
.A(n_1353),
.Y(n_1618)
);

NAND2xp5_ASAP7_75t_SL g1619 ( 
.A(n_1331),
.B(n_61),
.Y(n_1619)
);

NAND2xp5_ASAP7_75t_L g1620 ( 
.A(n_1334),
.B(n_62),
.Y(n_1620)
);

OAI21xp5_ASAP7_75t_L g1621 ( 
.A1(n_1385),
.A2(n_437),
.B(n_436),
.Y(n_1621)
);

AOI21xp5_ASAP7_75t_L g1622 ( 
.A1(n_1388),
.A2(n_440),
.B(n_439),
.Y(n_1622)
);

O2A1O1Ixp5_ASAP7_75t_L g1623 ( 
.A1(n_1423),
.A2(n_64),
.B(n_62),
.C(n_63),
.Y(n_1623)
);

NAND2xp5_ASAP7_75t_SL g1624 ( 
.A(n_1451),
.B(n_63),
.Y(n_1624)
);

INVx4_ASAP7_75t_L g1625 ( 
.A(n_1376),
.Y(n_1625)
);

BUFx3_ASAP7_75t_L g1626 ( 
.A(n_1495),
.Y(n_1626)
);

BUFx2_ASAP7_75t_L g1627 ( 
.A(n_1410),
.Y(n_1627)
);

NOR2xp33_ASAP7_75t_SL g1628 ( 
.A(n_1336),
.B(n_446),
.Y(n_1628)
);

NAND2xp5_ASAP7_75t_SL g1629 ( 
.A(n_1373),
.B(n_65),
.Y(n_1629)
);

INVx1_ASAP7_75t_L g1630 ( 
.A(n_1421),
.Y(n_1630)
);

HB1xp67_ASAP7_75t_L g1631 ( 
.A(n_1446),
.Y(n_1631)
);

AOI22xp5_ASAP7_75t_L g1632 ( 
.A1(n_1378),
.A2(n_67),
.B1(n_65),
.B2(n_66),
.Y(n_1632)
);

BUFx6f_ASAP7_75t_L g1633 ( 
.A(n_1481),
.Y(n_1633)
);

NOR2xp67_ASAP7_75t_SL g1634 ( 
.A(n_1332),
.B(n_66),
.Y(n_1634)
);

NAND2xp5_ASAP7_75t_L g1635 ( 
.A(n_1346),
.B(n_67),
.Y(n_1635)
);

A2O1A1Ixp33_ASAP7_75t_L g1636 ( 
.A1(n_1381),
.A2(n_70),
.B(n_68),
.C(n_69),
.Y(n_1636)
);

NAND2xp5_ASAP7_75t_L g1637 ( 
.A(n_1347),
.B(n_68),
.Y(n_1637)
);

AND2x4_ASAP7_75t_L g1638 ( 
.A(n_1354),
.B(n_553),
.Y(n_1638)
);

BUFx3_ASAP7_75t_L g1639 ( 
.A(n_1356),
.Y(n_1639)
);

AOI21xp5_ASAP7_75t_L g1640 ( 
.A1(n_1491),
.A2(n_452),
.B(n_451),
.Y(n_1640)
);

AND2x4_ASAP7_75t_L g1641 ( 
.A(n_1360),
.B(n_453),
.Y(n_1641)
);

INVx2_ASAP7_75t_SL g1642 ( 
.A(n_1362),
.Y(n_1642)
);

AND2x4_ASAP7_75t_L g1643 ( 
.A(n_1445),
.B(n_552),
.Y(n_1643)
);

INVx1_ASAP7_75t_L g1644 ( 
.A(n_1389),
.Y(n_1644)
);

O2A1O1Ixp5_ASAP7_75t_L g1645 ( 
.A1(n_1329),
.A2(n_73),
.B(n_71),
.C(n_72),
.Y(n_1645)
);

NAND2xp5_ASAP7_75t_L g1646 ( 
.A(n_1329),
.B(n_74),
.Y(n_1646)
);

BUFx6f_ASAP7_75t_L g1647 ( 
.A(n_1422),
.Y(n_1647)
);

AOI21xp5_ASAP7_75t_L g1648 ( 
.A1(n_1456),
.A2(n_456),
.B(n_454),
.Y(n_1648)
);

AOI21xp5_ASAP7_75t_L g1649 ( 
.A1(n_1407),
.A2(n_458),
.B(n_457),
.Y(n_1649)
);

NAND2xp5_ASAP7_75t_L g1650 ( 
.A(n_1351),
.B(n_74),
.Y(n_1650)
);

A2O1A1Ixp33_ASAP7_75t_L g1651 ( 
.A1(n_1397),
.A2(n_77),
.B(n_75),
.C(n_76),
.Y(n_1651)
);

NAND2xp5_ASAP7_75t_L g1652 ( 
.A(n_1379),
.B(n_76),
.Y(n_1652)
);

NAND2xp5_ASAP7_75t_L g1653 ( 
.A(n_1393),
.B(n_78),
.Y(n_1653)
);

OAI21xp5_ASAP7_75t_L g1654 ( 
.A1(n_1436),
.A2(n_460),
.B(n_459),
.Y(n_1654)
);

AOI21xp5_ASAP7_75t_L g1655 ( 
.A1(n_1460),
.A2(n_463),
.B(n_461),
.Y(n_1655)
);

INVxp67_ASAP7_75t_L g1656 ( 
.A(n_1420),
.Y(n_1656)
);

INVx2_ASAP7_75t_L g1657 ( 
.A(n_1467),
.Y(n_1657)
);

AOI21xp5_ASAP7_75t_L g1658 ( 
.A1(n_1469),
.A2(n_466),
.B(n_464),
.Y(n_1658)
);

AOI21xp5_ASAP7_75t_L g1659 ( 
.A1(n_1516),
.A2(n_1428),
.B(n_1427),
.Y(n_1659)
);

OAI21xp5_ASAP7_75t_L g1660 ( 
.A1(n_1577),
.A2(n_1452),
.B(n_1420),
.Y(n_1660)
);

HB1xp67_ASAP7_75t_L g1661 ( 
.A(n_1500),
.Y(n_1661)
);

O2A1O1Ixp33_ASAP7_75t_SL g1662 ( 
.A1(n_1524),
.A2(n_1457),
.B(n_1459),
.C(n_1458),
.Y(n_1662)
);

A2O1A1Ixp33_ASAP7_75t_L g1663 ( 
.A1(n_1537),
.A2(n_1454),
.B(n_1428),
.C(n_1434),
.Y(n_1663)
);

AOI22xp5_ASAP7_75t_L g1664 ( 
.A1(n_1550),
.A2(n_1448),
.B1(n_1458),
.B2(n_1457),
.Y(n_1664)
);

AO32x1_ASAP7_75t_L g1665 ( 
.A1(n_1644),
.A2(n_1435),
.A3(n_1438),
.B1(n_1402),
.B2(n_1399),
.Y(n_1665)
);

A2O1A1Ixp33_ASAP7_75t_L g1666 ( 
.A1(n_1579),
.A2(n_1472),
.B(n_1459),
.C(n_1488),
.Y(n_1666)
);

AOI21xp5_ASAP7_75t_L g1667 ( 
.A1(n_1568),
.A2(n_1472),
.B(n_1488),
.Y(n_1667)
);

HB1xp67_ASAP7_75t_L g1668 ( 
.A(n_1507),
.Y(n_1668)
);

NAND2xp5_ASAP7_75t_L g1669 ( 
.A(n_1542),
.B(n_1448),
.Y(n_1669)
);

AOI21xp5_ASAP7_75t_L g1670 ( 
.A1(n_1498),
.A2(n_1438),
.B(n_1435),
.Y(n_1670)
);

BUFx2_ASAP7_75t_L g1671 ( 
.A(n_1587),
.Y(n_1671)
);

AOI21xp5_ASAP7_75t_L g1672 ( 
.A1(n_1503),
.A2(n_551),
.B(n_470),
.Y(n_1672)
);

NOR2x1_ASAP7_75t_SL g1673 ( 
.A(n_1529),
.B(n_469),
.Y(n_1673)
);

NAND2xp5_ASAP7_75t_L g1674 ( 
.A(n_1506),
.B(n_78),
.Y(n_1674)
);

INVx2_ASAP7_75t_L g1675 ( 
.A(n_1502),
.Y(n_1675)
);

CKINVDCx20_ASAP7_75t_R g1676 ( 
.A(n_1555),
.Y(n_1676)
);

AOI21xp5_ASAP7_75t_L g1677 ( 
.A1(n_1504),
.A2(n_550),
.B(n_472),
.Y(n_1677)
);

AO21x1_ASAP7_75t_L g1678 ( 
.A1(n_1654),
.A2(n_79),
.B(n_80),
.Y(n_1678)
);

AO21x1_ASAP7_75t_L g1679 ( 
.A1(n_1558),
.A2(n_79),
.B(n_80),
.Y(n_1679)
);

AND2x2_ASAP7_75t_L g1680 ( 
.A(n_1531),
.B(n_82),
.Y(n_1680)
);

INVx1_ASAP7_75t_L g1681 ( 
.A(n_1608),
.Y(n_1681)
);

INVx1_ASAP7_75t_L g1682 ( 
.A(n_1600),
.Y(n_1682)
);

AOI21xp5_ASAP7_75t_L g1683 ( 
.A1(n_1505),
.A2(n_549),
.B(n_474),
.Y(n_1683)
);

CKINVDCx5p33_ASAP7_75t_R g1684 ( 
.A(n_1574),
.Y(n_1684)
);

AND2x4_ASAP7_75t_L g1685 ( 
.A(n_1563),
.B(n_471),
.Y(n_1685)
);

OAI21xp5_ASAP7_75t_L g1686 ( 
.A1(n_1510),
.A2(n_82),
.B(n_83),
.Y(n_1686)
);

AOI22xp33_ASAP7_75t_L g1687 ( 
.A1(n_1567),
.A2(n_86),
.B1(n_84),
.B2(n_85),
.Y(n_1687)
);

INVx2_ASAP7_75t_L g1688 ( 
.A(n_1606),
.Y(n_1688)
);

NOR2xp33_ASAP7_75t_L g1689 ( 
.A(n_1624),
.B(n_476),
.Y(n_1689)
);

NAND2xp5_ASAP7_75t_L g1690 ( 
.A(n_1521),
.B(n_84),
.Y(n_1690)
);

CKINVDCx5p33_ASAP7_75t_R g1691 ( 
.A(n_1596),
.Y(n_1691)
);

OAI22xp5_ASAP7_75t_L g1692 ( 
.A1(n_1592),
.A2(n_1578),
.B1(n_1514),
.B2(n_1519),
.Y(n_1692)
);

OAI22xp5_ASAP7_75t_L g1693 ( 
.A1(n_1514),
.A2(n_87),
.B1(n_85),
.B2(n_86),
.Y(n_1693)
);

OR2x6_ASAP7_75t_L g1694 ( 
.A(n_1549),
.B(n_478),
.Y(n_1694)
);

AOI21x1_ASAP7_75t_L g1695 ( 
.A1(n_1576),
.A2(n_480),
.B(n_479),
.Y(n_1695)
);

BUFx3_ASAP7_75t_L g1696 ( 
.A(n_1543),
.Y(n_1696)
);

INVx3_ASAP7_75t_L g1697 ( 
.A(n_1587),
.Y(n_1697)
);

INVx1_ASAP7_75t_SL g1698 ( 
.A(n_1551),
.Y(n_1698)
);

INVx5_ASAP7_75t_L g1699 ( 
.A(n_1549),
.Y(n_1699)
);

AOI21xp5_ASAP7_75t_L g1700 ( 
.A1(n_1499),
.A2(n_546),
.B(n_486),
.Y(n_1700)
);

INVx1_ASAP7_75t_L g1701 ( 
.A(n_1610),
.Y(n_1701)
);

INVx1_ASAP7_75t_L g1702 ( 
.A(n_1520),
.Y(n_1702)
);

O2A1O1Ixp33_ASAP7_75t_SL g1703 ( 
.A1(n_1548),
.A2(n_89),
.B(n_87),
.C(n_88),
.Y(n_1703)
);

INVxp67_ASAP7_75t_L g1704 ( 
.A(n_1522),
.Y(n_1704)
);

O2A1O1Ixp33_ASAP7_75t_L g1705 ( 
.A1(n_1539),
.A2(n_91),
.B(n_88),
.C(n_89),
.Y(n_1705)
);

A2O1A1Ixp33_ASAP7_75t_L g1706 ( 
.A1(n_1643),
.A2(n_94),
.B(n_91),
.C(n_93),
.Y(n_1706)
);

NOR2xp33_ASAP7_75t_L g1707 ( 
.A(n_1619),
.B(n_483),
.Y(n_1707)
);

AND2x4_ASAP7_75t_L g1708 ( 
.A(n_1511),
.B(n_488),
.Y(n_1708)
);

OAI22xp5_ASAP7_75t_L g1709 ( 
.A1(n_1510),
.A2(n_96),
.B1(n_94),
.B2(n_95),
.Y(n_1709)
);

O2A1O1Ixp33_ASAP7_75t_L g1710 ( 
.A1(n_1629),
.A2(n_98),
.B(n_95),
.C(n_97),
.Y(n_1710)
);

OAI22xp5_ASAP7_75t_L g1711 ( 
.A1(n_1525),
.A2(n_99),
.B1(n_97),
.B2(n_98),
.Y(n_1711)
);

BUFx6f_ASAP7_75t_L g1712 ( 
.A(n_1612),
.Y(n_1712)
);

AOI22xp33_ASAP7_75t_L g1713 ( 
.A1(n_1557),
.A2(n_102),
.B1(n_100),
.B2(n_101),
.Y(n_1713)
);

NAND2xp5_ASAP7_75t_SL g1714 ( 
.A(n_1643),
.B(n_100),
.Y(n_1714)
);

AOI21xp5_ASAP7_75t_L g1715 ( 
.A1(n_1512),
.A2(n_545),
.B(n_496),
.Y(n_1715)
);

INVxp67_ASAP7_75t_SL g1716 ( 
.A(n_1631),
.Y(n_1716)
);

INVx1_ASAP7_75t_L g1717 ( 
.A(n_1532),
.Y(n_1717)
);

AND2x2_ASAP7_75t_L g1718 ( 
.A(n_1552),
.B(n_101),
.Y(n_1718)
);

OR2x6_ASAP7_75t_SL g1719 ( 
.A(n_1618),
.B(n_1653),
.Y(n_1719)
);

NAND2xp5_ASAP7_75t_L g1720 ( 
.A(n_1535),
.B(n_102),
.Y(n_1720)
);

NOR3xp33_ASAP7_75t_L g1721 ( 
.A(n_1584),
.B(n_103),
.C(n_104),
.Y(n_1721)
);

CKINVDCx5p33_ASAP7_75t_R g1722 ( 
.A(n_1540),
.Y(n_1722)
);

INVx3_ASAP7_75t_SL g1723 ( 
.A(n_1515),
.Y(n_1723)
);

NAND3xp33_ASAP7_75t_SL g1724 ( 
.A(n_1530),
.B(n_103),
.C(n_104),
.Y(n_1724)
);

HB1xp67_ASAP7_75t_L g1725 ( 
.A(n_1612),
.Y(n_1725)
);

AOI21xp5_ASAP7_75t_L g1726 ( 
.A1(n_1509),
.A2(n_541),
.B(n_497),
.Y(n_1726)
);

INVx2_ASAP7_75t_SL g1727 ( 
.A(n_1543),
.Y(n_1727)
);

OAI22xp5_ASAP7_75t_L g1728 ( 
.A1(n_1656),
.A2(n_107),
.B1(n_105),
.B2(n_106),
.Y(n_1728)
);

O2A1O1Ixp33_ASAP7_75t_L g1729 ( 
.A1(n_1636),
.A2(n_108),
.B(n_106),
.C(n_107),
.Y(n_1729)
);

AND2x4_ASAP7_75t_L g1730 ( 
.A(n_1511),
.B(n_492),
.Y(n_1730)
);

AND2x4_ASAP7_75t_L g1731 ( 
.A(n_1586),
.B(n_498),
.Y(n_1731)
);

A2O1A1Ixp33_ASAP7_75t_SL g1732 ( 
.A1(n_1634),
.A2(n_110),
.B(n_108),
.C(n_109),
.Y(n_1732)
);

INVx1_ASAP7_75t_L g1733 ( 
.A(n_1560),
.Y(n_1733)
);

BUFx4f_ASAP7_75t_SL g1734 ( 
.A(n_1609),
.Y(n_1734)
);

NOR2xp33_ASAP7_75t_R g1735 ( 
.A(n_1543),
.B(n_502),
.Y(n_1735)
);

NOR2xp33_ASAP7_75t_L g1736 ( 
.A(n_1586),
.B(n_503),
.Y(n_1736)
);

INVx1_ASAP7_75t_L g1737 ( 
.A(n_1564),
.Y(n_1737)
);

AOI21xp5_ASAP7_75t_L g1738 ( 
.A1(n_1575),
.A2(n_539),
.B(n_505),
.Y(n_1738)
);

AOI21xp5_ASAP7_75t_L g1739 ( 
.A1(n_1582),
.A2(n_1538),
.B(n_1604),
.Y(n_1739)
);

INVx1_ASAP7_75t_SL g1740 ( 
.A(n_1515),
.Y(n_1740)
);

NOR2xp33_ASAP7_75t_L g1741 ( 
.A(n_1639),
.B(n_504),
.Y(n_1741)
);

INVx2_ASAP7_75t_L g1742 ( 
.A(n_1556),
.Y(n_1742)
);

BUFx6f_ASAP7_75t_L g1743 ( 
.A(n_1554),
.Y(n_1743)
);

NOR2xp33_ASAP7_75t_L g1744 ( 
.A(n_1611),
.B(n_506),
.Y(n_1744)
);

AOI21xp5_ASAP7_75t_L g1745 ( 
.A1(n_1621),
.A2(n_538),
.B(n_508),
.Y(n_1745)
);

NAND2xp5_ASAP7_75t_L g1746 ( 
.A(n_1545),
.B(n_109),
.Y(n_1746)
);

INVx2_ASAP7_75t_L g1747 ( 
.A(n_1573),
.Y(n_1747)
);

BUFx6f_ASAP7_75t_L g1748 ( 
.A(n_1554),
.Y(n_1748)
);

OR2x2_ASAP7_75t_L g1749 ( 
.A(n_1547),
.B(n_110),
.Y(n_1749)
);

AND2x4_ASAP7_75t_L g1750 ( 
.A(n_1605),
.B(n_507),
.Y(n_1750)
);

XNOR2xp5_ASAP7_75t_L g1751 ( 
.A(n_1598),
.B(n_511),
.Y(n_1751)
);

BUFx3_ASAP7_75t_L g1752 ( 
.A(n_1549),
.Y(n_1752)
);

NOR2xp33_ASAP7_75t_SL g1753 ( 
.A(n_1601),
.B(n_512),
.Y(n_1753)
);

INVx1_ASAP7_75t_L g1754 ( 
.A(n_1581),
.Y(n_1754)
);

INVx1_ASAP7_75t_SL g1755 ( 
.A(n_1595),
.Y(n_1755)
);

NAND2xp5_ASAP7_75t_L g1756 ( 
.A(n_1569),
.B(n_111),
.Y(n_1756)
);

NAND2xp5_ASAP7_75t_SL g1757 ( 
.A(n_1638),
.B(n_112),
.Y(n_1757)
);

HB1xp67_ASAP7_75t_L g1758 ( 
.A(n_1642),
.Y(n_1758)
);

NAND2xp5_ASAP7_75t_L g1759 ( 
.A(n_1570),
.B(n_114),
.Y(n_1759)
);

OAI22xp5_ASAP7_75t_L g1760 ( 
.A1(n_1571),
.A2(n_117),
.B1(n_115),
.B2(n_116),
.Y(n_1760)
);

AOI21xp5_ASAP7_75t_L g1761 ( 
.A1(n_1528),
.A2(n_535),
.B(n_515),
.Y(n_1761)
);

NAND2xp5_ASAP7_75t_L g1762 ( 
.A(n_1513),
.B(n_115),
.Y(n_1762)
);

NOR2xp33_ASAP7_75t_R g1763 ( 
.A(n_1605),
.B(n_514),
.Y(n_1763)
);

OAI22xp5_ASAP7_75t_L g1764 ( 
.A1(n_1630),
.A2(n_119),
.B1(n_116),
.B2(n_118),
.Y(n_1764)
);

INVx1_ASAP7_75t_L g1765 ( 
.A(n_1635),
.Y(n_1765)
);

AND2x2_ASAP7_75t_L g1766 ( 
.A(n_1585),
.B(n_119),
.Y(n_1766)
);

NAND2xp5_ASAP7_75t_L g1767 ( 
.A(n_1544),
.B(n_120),
.Y(n_1767)
);

AOI21xp5_ASAP7_75t_L g1768 ( 
.A1(n_1628),
.A2(n_534),
.B(n_517),
.Y(n_1768)
);

OAI21xp5_ASAP7_75t_L g1769 ( 
.A1(n_1527),
.A2(n_121),
.B(n_122),
.Y(n_1769)
);

INVx1_ASAP7_75t_L g1770 ( 
.A(n_1637),
.Y(n_1770)
);

CKINVDCx5p33_ASAP7_75t_R g1771 ( 
.A(n_1594),
.Y(n_1771)
);

AOI22xp5_ASAP7_75t_L g1772 ( 
.A1(n_1584),
.A2(n_125),
.B1(n_121),
.B2(n_122),
.Y(n_1772)
);

INVx1_ASAP7_75t_L g1773 ( 
.A(n_1593),
.Y(n_1773)
);

NAND2xp5_ASAP7_75t_L g1774 ( 
.A(n_1588),
.B(n_126),
.Y(n_1774)
);

AND2x2_ASAP7_75t_L g1775 ( 
.A(n_1602),
.B(n_1559),
.Y(n_1775)
);

BUFx2_ASAP7_75t_L g1776 ( 
.A(n_1633),
.Y(n_1776)
);

AOI21xp5_ASAP7_75t_L g1777 ( 
.A1(n_1572),
.A2(n_518),
.B(n_516),
.Y(n_1777)
);

A2O1A1Ixp33_ASAP7_75t_L g1778 ( 
.A1(n_1553),
.A2(n_128),
.B(n_126),
.C(n_127),
.Y(n_1778)
);

NAND2xp5_ASAP7_75t_L g1779 ( 
.A(n_1533),
.B(n_129),
.Y(n_1779)
);

BUFx6f_ASAP7_75t_L g1780 ( 
.A(n_1647),
.Y(n_1780)
);

AOI21xp5_ASAP7_75t_L g1781 ( 
.A1(n_1517),
.A2(n_521),
.B(n_520),
.Y(n_1781)
);

BUFx6f_ASAP7_75t_L g1782 ( 
.A(n_1647),
.Y(n_1782)
);

OAI21xp33_ASAP7_75t_L g1783 ( 
.A1(n_1533),
.A2(n_130),
.B(n_131),
.Y(n_1783)
);

INVx2_ASAP7_75t_SL g1784 ( 
.A(n_1626),
.Y(n_1784)
);

AOI21xp33_ASAP7_75t_L g1785 ( 
.A1(n_1536),
.A2(n_130),
.B(n_131),
.Y(n_1785)
);

AND2x4_ASAP7_75t_L g1786 ( 
.A(n_1508),
.B(n_522),
.Y(n_1786)
);

INVx1_ASAP7_75t_L g1787 ( 
.A(n_1633),
.Y(n_1787)
);

NAND2xp5_ASAP7_75t_L g1788 ( 
.A(n_1536),
.B(n_132),
.Y(n_1788)
);

AOI21xp5_ASAP7_75t_L g1789 ( 
.A1(n_1523),
.A2(n_531),
.B(n_524),
.Y(n_1789)
);

INVx1_ASAP7_75t_L g1790 ( 
.A(n_1565),
.Y(n_1790)
);

BUFx2_ASAP7_75t_L g1791 ( 
.A(n_1559),
.Y(n_1791)
);

NAND2xp5_ASAP7_75t_L g1792 ( 
.A(n_1508),
.B(n_134),
.Y(n_1792)
);

AOI221xp5_ASAP7_75t_L g1793 ( 
.A1(n_1566),
.A2(n_135),
.B1(n_136),
.B2(n_137),
.C(n_138),
.Y(n_1793)
);

BUFx8_ASAP7_75t_L g1794 ( 
.A(n_1647),
.Y(n_1794)
);

AOI21xp5_ASAP7_75t_L g1795 ( 
.A1(n_1501),
.A2(n_530),
.B(n_526),
.Y(n_1795)
);

BUFx12f_ASAP7_75t_L g1796 ( 
.A(n_1589),
.Y(n_1796)
);

A2O1A1Ixp33_ASAP7_75t_SL g1797 ( 
.A1(n_1599),
.A2(n_137),
.B(n_135),
.C(n_136),
.Y(n_1797)
);

CKINVDCx5p33_ASAP7_75t_R g1798 ( 
.A(n_1603),
.Y(n_1798)
);

INVx2_ASAP7_75t_SL g1799 ( 
.A(n_1657),
.Y(n_1799)
);

AOI21xp5_ASAP7_75t_L g1800 ( 
.A1(n_1648),
.A2(n_527),
.B(n_523),
.Y(n_1800)
);

BUFx6f_ASAP7_75t_L g1801 ( 
.A(n_1615),
.Y(n_1801)
);

BUFx12f_ASAP7_75t_L g1802 ( 
.A(n_1589),
.Y(n_1802)
);

BUFx12f_ASAP7_75t_L g1803 ( 
.A(n_1638),
.Y(n_1803)
);

AOI31xp67_ASAP7_75t_L g1804 ( 
.A1(n_1664),
.A2(n_1617),
.A3(n_1620),
.B(n_1614),
.Y(n_1804)
);

OAI22x1_ASAP7_75t_L g1805 ( 
.A1(n_1772),
.A2(n_1632),
.B1(n_1627),
.B2(n_1546),
.Y(n_1805)
);

NAND3xp33_ASAP7_75t_L g1806 ( 
.A(n_1769),
.B(n_1632),
.C(n_1651),
.Y(n_1806)
);

A2O1A1Ixp33_ASAP7_75t_L g1807 ( 
.A1(n_1739),
.A2(n_1623),
.B(n_1645),
.C(n_1640),
.Y(n_1807)
);

NAND2xp5_ASAP7_75t_L g1808 ( 
.A(n_1681),
.B(n_1765),
.Y(n_1808)
);

INVx1_ASAP7_75t_L g1809 ( 
.A(n_1702),
.Y(n_1809)
);

OAI21xp5_ASAP7_75t_L g1810 ( 
.A1(n_1745),
.A2(n_1561),
.B(n_1518),
.Y(n_1810)
);

OAI21x1_ASAP7_75t_L g1811 ( 
.A1(n_1695),
.A2(n_1541),
.B(n_1616),
.Y(n_1811)
);

OA22x2_ASAP7_75t_L g1812 ( 
.A1(n_1772),
.A2(n_1562),
.B1(n_1583),
.B2(n_1652),
.Y(n_1812)
);

OR2x6_ASAP7_75t_L g1813 ( 
.A(n_1694),
.B(n_1625),
.Y(n_1813)
);

BUFx4f_ASAP7_75t_SL g1814 ( 
.A(n_1676),
.Y(n_1814)
);

AO21x1_ASAP7_75t_L g1815 ( 
.A1(n_1721),
.A2(n_1646),
.B(n_1650),
.Y(n_1815)
);

BUFx3_ASAP7_75t_L g1816 ( 
.A(n_1723),
.Y(n_1816)
);

INVx1_ASAP7_75t_L g1817 ( 
.A(n_1717),
.Y(n_1817)
);

OA22x2_ASAP7_75t_L g1818 ( 
.A1(n_1660),
.A2(n_1580),
.B1(n_1641),
.B2(n_1534),
.Y(n_1818)
);

BUFx4f_ASAP7_75t_L g1819 ( 
.A(n_1694),
.Y(n_1819)
);

NOR2x1_ASAP7_75t_SL g1820 ( 
.A(n_1773),
.B(n_1625),
.Y(n_1820)
);

CKINVDCx16_ASAP7_75t_R g1821 ( 
.A(n_1752),
.Y(n_1821)
);

OAI21x1_ASAP7_75t_L g1822 ( 
.A1(n_1715),
.A2(n_1591),
.B(n_1622),
.Y(n_1822)
);

AND2x2_ASAP7_75t_L g1823 ( 
.A(n_1775),
.B(n_1597),
.Y(n_1823)
);

INVxp67_ASAP7_75t_SL g1824 ( 
.A(n_1716),
.Y(n_1824)
);

AOI21xp5_ASAP7_75t_L g1825 ( 
.A1(n_1738),
.A2(n_1613),
.B(n_1607),
.Y(n_1825)
);

NAND2xp5_ASAP7_75t_L g1826 ( 
.A(n_1770),
.B(n_1526),
.Y(n_1826)
);

OR2x6_ASAP7_75t_L g1827 ( 
.A(n_1803),
.B(n_1590),
.Y(n_1827)
);

HB1xp67_ASAP7_75t_L g1828 ( 
.A(n_1661),
.Y(n_1828)
);

INVx3_ASAP7_75t_L g1829 ( 
.A(n_1712),
.Y(n_1829)
);

BUFx6f_ASAP7_75t_L g1830 ( 
.A(n_1712),
.Y(n_1830)
);

AND2x4_ASAP7_75t_L g1831 ( 
.A(n_1671),
.B(n_1655),
.Y(n_1831)
);

OAI21xp5_ASAP7_75t_SL g1832 ( 
.A1(n_1713),
.A2(n_1658),
.B(n_1649),
.Y(n_1832)
);

NOR3xp33_ASAP7_75t_L g1833 ( 
.A(n_1724),
.B(n_139),
.C(n_140),
.Y(n_1833)
);

NAND2xp5_ASAP7_75t_SL g1834 ( 
.A(n_1801),
.B(n_528),
.Y(n_1834)
);

BUFx2_ASAP7_75t_L g1835 ( 
.A(n_1712),
.Y(n_1835)
);

AOI21xp5_ASAP7_75t_L g1836 ( 
.A1(n_1800),
.A2(n_529),
.B(n_141),
.Y(n_1836)
);

OAI21x1_ASAP7_75t_L g1837 ( 
.A1(n_1790),
.A2(n_141),
.B(n_142),
.Y(n_1837)
);

OAI21x1_ASAP7_75t_L g1838 ( 
.A1(n_1726),
.A2(n_142),
.B(n_143),
.Y(n_1838)
);

NOR2xp67_ASAP7_75t_SL g1839 ( 
.A(n_1699),
.B(n_144),
.Y(n_1839)
);

AOI21xp5_ASAP7_75t_L g1840 ( 
.A1(n_1768),
.A2(n_145),
.B(n_147),
.Y(n_1840)
);

CKINVDCx5p33_ASAP7_75t_R g1841 ( 
.A(n_1722),
.Y(n_1841)
);

AOI21xp5_ASAP7_75t_L g1842 ( 
.A1(n_1777),
.A2(n_145),
.B(n_147),
.Y(n_1842)
);

AOI21xp5_ASAP7_75t_L g1843 ( 
.A1(n_1673),
.A2(n_148),
.B(n_149),
.Y(n_1843)
);

NAND2xp5_ASAP7_75t_SL g1844 ( 
.A(n_1801),
.B(n_148),
.Y(n_1844)
);

AO21x2_ASAP7_75t_L g1845 ( 
.A1(n_1667),
.A2(n_150),
.B(n_151),
.Y(n_1845)
);

OA21x2_ASAP7_75t_L g1846 ( 
.A1(n_1659),
.A2(n_151),
.B(n_152),
.Y(n_1846)
);

NAND2xp5_ASAP7_75t_L g1847 ( 
.A(n_1755),
.B(n_152),
.Y(n_1847)
);

NAND2xp5_ASAP7_75t_L g1848 ( 
.A(n_1668),
.B(n_374),
.Y(n_1848)
);

INVx1_ASAP7_75t_L g1849 ( 
.A(n_1733),
.Y(n_1849)
);

O2A1O1Ixp33_ASAP7_75t_L g1850 ( 
.A1(n_1706),
.A2(n_155),
.B(n_153),
.C(n_154),
.Y(n_1850)
);

OAI21x1_ASAP7_75t_SL g1851 ( 
.A1(n_1678),
.A2(n_1686),
.B(n_1679),
.Y(n_1851)
);

AOI21xp5_ASAP7_75t_L g1852 ( 
.A1(n_1753),
.A2(n_1714),
.B(n_1761),
.Y(n_1852)
);

NAND2xp5_ASAP7_75t_L g1853 ( 
.A(n_1762),
.B(n_374),
.Y(n_1853)
);

INVx1_ASAP7_75t_L g1854 ( 
.A(n_1737),
.Y(n_1854)
);

AOI21xp5_ASAP7_75t_L g1855 ( 
.A1(n_1781),
.A2(n_153),
.B(n_154),
.Y(n_1855)
);

NOR4xp25_ASAP7_75t_L g1856 ( 
.A(n_1666),
.B(n_157),
.C(n_155),
.D(n_156),
.Y(n_1856)
);

AOI221x1_ASAP7_75t_L g1857 ( 
.A1(n_1663),
.A2(n_156),
.B1(n_158),
.B2(n_159),
.C(n_160),
.Y(n_1857)
);

NAND2xp5_ASAP7_75t_L g1858 ( 
.A(n_1675),
.B(n_1688),
.Y(n_1858)
);

OA21x2_ASAP7_75t_L g1859 ( 
.A1(n_1670),
.A2(n_161),
.B(n_162),
.Y(n_1859)
);

AOI21xp5_ASAP7_75t_L g1860 ( 
.A1(n_1789),
.A2(n_1662),
.B(n_1672),
.Y(n_1860)
);

AND2x2_ASAP7_75t_L g1861 ( 
.A(n_1766),
.B(n_163),
.Y(n_1861)
);

AOI21x1_ASAP7_75t_L g1862 ( 
.A1(n_1692),
.A2(n_164),
.B(n_166),
.Y(n_1862)
);

A2O1A1Ixp33_ASAP7_75t_L g1863 ( 
.A1(n_1729),
.A2(n_168),
.B(n_166),
.C(n_167),
.Y(n_1863)
);

BUFx3_ASAP7_75t_L g1864 ( 
.A(n_1696),
.Y(n_1864)
);

AOI21xp5_ASAP7_75t_L g1865 ( 
.A1(n_1677),
.A2(n_168),
.B(n_169),
.Y(n_1865)
);

AND2x4_ASAP7_75t_L g1866 ( 
.A(n_1697),
.B(n_169),
.Y(n_1866)
);

A2O1A1Ixp33_ASAP7_75t_L g1867 ( 
.A1(n_1783),
.A2(n_172),
.B(n_170),
.C(n_171),
.Y(n_1867)
);

AOI21xp5_ASAP7_75t_L g1868 ( 
.A1(n_1683),
.A2(n_171),
.B(n_172),
.Y(n_1868)
);

NOR2xp67_ASAP7_75t_L g1869 ( 
.A(n_1704),
.B(n_173),
.Y(n_1869)
);

AOI22xp5_ASAP7_75t_L g1870 ( 
.A1(n_1689),
.A2(n_175),
.B1(n_173),
.B2(n_174),
.Y(n_1870)
);

A2O1A1Ixp33_ASAP7_75t_L g1871 ( 
.A1(n_1785),
.A2(n_176),
.B(n_174),
.C(n_175),
.Y(n_1871)
);

OAI21xp5_ASAP7_75t_L g1872 ( 
.A1(n_1710),
.A2(n_178),
.B(n_180),
.Y(n_1872)
);

AOI21xp5_ASAP7_75t_L g1873 ( 
.A1(n_1700),
.A2(n_180),
.B(n_181),
.Y(n_1873)
);

INVx1_ASAP7_75t_L g1874 ( 
.A(n_1754),
.Y(n_1874)
);

OAI21x1_ASAP7_75t_L g1875 ( 
.A1(n_1795),
.A2(n_182),
.B(n_185),
.Y(n_1875)
);

NAND3xp33_ASAP7_75t_L g1876 ( 
.A(n_1687),
.B(n_1693),
.C(n_1690),
.Y(n_1876)
);

INVx1_ASAP7_75t_L g1877 ( 
.A(n_1682),
.Y(n_1877)
);

NAND2xp5_ASAP7_75t_L g1878 ( 
.A(n_1701),
.B(n_187),
.Y(n_1878)
);

AOI21xp5_ASAP7_75t_L g1879 ( 
.A1(n_1778),
.A2(n_189),
.B(n_190),
.Y(n_1879)
);

INVxp67_ASAP7_75t_SL g1880 ( 
.A(n_1758),
.Y(n_1880)
);

A2O1A1Ixp33_ASAP7_75t_L g1881 ( 
.A1(n_1707),
.A2(n_189),
.B(n_190),
.C(n_191),
.Y(n_1881)
);

OAI21xp5_ASAP7_75t_L g1882 ( 
.A1(n_1793),
.A2(n_192),
.B(n_193),
.Y(n_1882)
);

INVx3_ASAP7_75t_L g1883 ( 
.A(n_1786),
.Y(n_1883)
);

OAI21x1_ASAP7_75t_L g1884 ( 
.A1(n_1742),
.A2(n_194),
.B(n_195),
.Y(n_1884)
);

AOI21xp5_ASAP7_75t_L g1885 ( 
.A1(n_1703),
.A2(n_1732),
.B(n_1665),
.Y(n_1885)
);

INVx1_ASAP7_75t_L g1886 ( 
.A(n_1747),
.Y(n_1886)
);

AND2x6_ASAP7_75t_L g1887 ( 
.A(n_1801),
.B(n_195),
.Y(n_1887)
);

INVx1_ASAP7_75t_L g1888 ( 
.A(n_1665),
.Y(n_1888)
);

AOI21xp5_ASAP7_75t_L g1889 ( 
.A1(n_1665),
.A2(n_196),
.B(n_197),
.Y(n_1889)
);

CKINVDCx20_ASAP7_75t_R g1890 ( 
.A(n_1734),
.Y(n_1890)
);

NAND2xp5_ASAP7_75t_L g1891 ( 
.A(n_1779),
.B(n_373),
.Y(n_1891)
);

BUFx2_ASAP7_75t_L g1892 ( 
.A(n_1697),
.Y(n_1892)
);

NOR2xp67_ASAP7_75t_SL g1893 ( 
.A(n_1699),
.B(n_196),
.Y(n_1893)
);

INVx3_ASAP7_75t_L g1894 ( 
.A(n_1809),
.Y(n_1894)
);

INVx2_ASAP7_75t_SL g1895 ( 
.A(n_1817),
.Y(n_1895)
);

OAI21x1_ASAP7_75t_L g1896 ( 
.A1(n_1811),
.A2(n_1788),
.B(n_1705),
.Y(n_1896)
);

OA21x2_ASAP7_75t_L g1897 ( 
.A1(n_1807),
.A2(n_1669),
.B(n_1746),
.Y(n_1897)
);

CKINVDCx11_ASAP7_75t_R g1898 ( 
.A(n_1890),
.Y(n_1898)
);

INVxp67_ASAP7_75t_SL g1899 ( 
.A(n_1824),
.Y(n_1899)
);

INVx1_ASAP7_75t_L g1900 ( 
.A(n_1849),
.Y(n_1900)
);

NAND2x1p5_ASAP7_75t_L g1901 ( 
.A(n_1819),
.B(n_1699),
.Y(n_1901)
);

INVx1_ASAP7_75t_L g1902 ( 
.A(n_1854),
.Y(n_1902)
);

AOI21x1_ASAP7_75t_L g1903 ( 
.A1(n_1862),
.A2(n_1709),
.B(n_1760),
.Y(n_1903)
);

OAI22xp5_ASAP7_75t_L g1904 ( 
.A1(n_1806),
.A2(n_1767),
.B1(n_1719),
.B2(n_1796),
.Y(n_1904)
);

OAI21x1_ASAP7_75t_L g1905 ( 
.A1(n_1822),
.A2(n_1792),
.B(n_1787),
.Y(n_1905)
);

OR2x2_ASAP7_75t_L g1906 ( 
.A(n_1828),
.B(n_1674),
.Y(n_1906)
);

BUFx8_ASAP7_75t_L g1907 ( 
.A(n_1887),
.Y(n_1907)
);

NAND2xp5_ASAP7_75t_L g1908 ( 
.A(n_1808),
.B(n_1880),
.Y(n_1908)
);

AOI222xp33_ASAP7_75t_L g1909 ( 
.A1(n_1882),
.A2(n_1711),
.B1(n_1802),
.B2(n_1720),
.C1(n_1728),
.C2(n_1756),
.Y(n_1909)
);

NOR2xp33_ASAP7_75t_L g1910 ( 
.A(n_1826),
.B(n_1759),
.Y(n_1910)
);

HB1xp67_ASAP7_75t_L g1911 ( 
.A(n_1874),
.Y(n_1911)
);

A2O1A1Ixp33_ASAP7_75t_L g1912 ( 
.A1(n_1850),
.A2(n_1757),
.B(n_1731),
.C(n_1736),
.Y(n_1912)
);

BUFx2_ASAP7_75t_L g1913 ( 
.A(n_1892),
.Y(n_1913)
);

OAI21x1_ASAP7_75t_SL g1914 ( 
.A1(n_1815),
.A2(n_1764),
.B(n_1774),
.Y(n_1914)
);

INVx1_ASAP7_75t_L g1915 ( 
.A(n_1877),
.Y(n_1915)
);

BUFx3_ASAP7_75t_L g1916 ( 
.A(n_1816),
.Y(n_1916)
);

OAI21xp5_ASAP7_75t_L g1917 ( 
.A1(n_1860),
.A2(n_1797),
.B(n_1741),
.Y(n_1917)
);

NOR2xp67_ASAP7_75t_L g1918 ( 
.A(n_1853),
.B(n_1784),
.Y(n_1918)
);

NOR2xp67_ASAP7_75t_L g1919 ( 
.A(n_1886),
.B(n_1749),
.Y(n_1919)
);

AO21x2_ASAP7_75t_L g1920 ( 
.A1(n_1851),
.A2(n_1744),
.B(n_1763),
.Y(n_1920)
);

OAI21x1_ASAP7_75t_L g1921 ( 
.A1(n_1825),
.A2(n_1725),
.B(n_1680),
.Y(n_1921)
);

AND2x2_ASAP7_75t_L g1922 ( 
.A(n_1888),
.B(n_1718),
.Y(n_1922)
);

NAND2xp5_ASAP7_75t_L g1923 ( 
.A(n_1858),
.B(n_1891),
.Y(n_1923)
);

OA21x2_ASAP7_75t_L g1924 ( 
.A1(n_1885),
.A2(n_1776),
.B(n_1685),
.Y(n_1924)
);

AOI22xp33_ASAP7_75t_L g1925 ( 
.A1(n_1876),
.A2(n_1791),
.B1(n_1731),
.B2(n_1685),
.Y(n_1925)
);

AOI22xp33_ASAP7_75t_SL g1926 ( 
.A1(n_1812),
.A2(n_1735),
.B1(n_1786),
.B2(n_1708),
.Y(n_1926)
);

AND2x4_ASAP7_75t_L g1927 ( 
.A(n_1831),
.B(n_1780),
.Y(n_1927)
);

AND2x2_ASAP7_75t_L g1928 ( 
.A(n_1823),
.B(n_1698),
.Y(n_1928)
);

NOR2x1_ASAP7_75t_SL g1929 ( 
.A(n_1813),
.B(n_1743),
.Y(n_1929)
);

OR2x6_ASAP7_75t_L g1930 ( 
.A(n_1813),
.B(n_1852),
.Y(n_1930)
);

NAND2xp5_ASAP7_75t_L g1931 ( 
.A(n_1856),
.B(n_1751),
.Y(n_1931)
);

AO21x2_ASAP7_75t_L g1932 ( 
.A1(n_1810),
.A2(n_1750),
.B(n_1730),
.Y(n_1932)
);

AO21x2_ASAP7_75t_L g1933 ( 
.A1(n_1820),
.A2(n_1730),
.B(n_1740),
.Y(n_1933)
);

INVx1_ASAP7_75t_L g1934 ( 
.A(n_1804),
.Y(n_1934)
);

NAND2xp5_ASAP7_75t_L g1935 ( 
.A(n_1878),
.B(n_1799),
.Y(n_1935)
);

NAND2xp5_ASAP7_75t_SL g1936 ( 
.A(n_1833),
.B(n_1780),
.Y(n_1936)
);

AND2x2_ASAP7_75t_L g1937 ( 
.A(n_1846),
.B(n_1743),
.Y(n_1937)
);

INVx3_ASAP7_75t_SL g1938 ( 
.A(n_1841),
.Y(n_1938)
);

INVx2_ASAP7_75t_SL g1939 ( 
.A(n_1830),
.Y(n_1939)
);

AO21x2_ASAP7_75t_L g1940 ( 
.A1(n_1872),
.A2(n_1794),
.B(n_1748),
.Y(n_1940)
);

INVx2_ASAP7_75t_SL g1941 ( 
.A(n_1830),
.Y(n_1941)
);

OAI21x1_ASAP7_75t_SL g1942 ( 
.A1(n_1889),
.A2(n_1727),
.B(n_1691),
.Y(n_1942)
);

OA21x2_ASAP7_75t_L g1943 ( 
.A1(n_1838),
.A2(n_1798),
.B(n_1771),
.Y(n_1943)
);

INVx2_ASAP7_75t_SL g1944 ( 
.A(n_1830),
.Y(n_1944)
);

INVx1_ASAP7_75t_L g1945 ( 
.A(n_1846),
.Y(n_1945)
);

NOR2xp33_ASAP7_75t_L g1946 ( 
.A(n_1818),
.B(n_1780),
.Y(n_1946)
);

AND2x4_ASAP7_75t_L g1947 ( 
.A(n_1894),
.B(n_1831),
.Y(n_1947)
);

BUFx6f_ASAP7_75t_L g1948 ( 
.A(n_1930),
.Y(n_1948)
);

HB1xp67_ASAP7_75t_L g1949 ( 
.A(n_1937),
.Y(n_1949)
);

BUFx3_ASAP7_75t_L g1950 ( 
.A(n_1907),
.Y(n_1950)
);

INVx1_ASAP7_75t_L g1951 ( 
.A(n_1911),
.Y(n_1951)
);

INVx3_ASAP7_75t_L g1952 ( 
.A(n_1894),
.Y(n_1952)
);

INVx6_ASAP7_75t_L g1953 ( 
.A(n_1907),
.Y(n_1953)
);

OAI22xp33_ASAP7_75t_L g1954 ( 
.A1(n_1931),
.A2(n_1857),
.B1(n_1870),
.B2(n_1805),
.Y(n_1954)
);

INVx2_ASAP7_75t_L g1955 ( 
.A(n_1895),
.Y(n_1955)
);

AND2x4_ASAP7_75t_L g1956 ( 
.A(n_1895),
.B(n_1835),
.Y(n_1956)
);

NAND2x1p5_ASAP7_75t_L g1957 ( 
.A(n_1924),
.B(n_1859),
.Y(n_1957)
);

OAI21xp5_ASAP7_75t_SL g1958 ( 
.A1(n_1909),
.A2(n_1881),
.B(n_1879),
.Y(n_1958)
);

INVx1_ASAP7_75t_L g1959 ( 
.A(n_1900),
.Y(n_1959)
);

INVx2_ASAP7_75t_L g1960 ( 
.A(n_1902),
.Y(n_1960)
);

INVx1_ASAP7_75t_L g1961 ( 
.A(n_1915),
.Y(n_1961)
);

BUFx2_ASAP7_75t_SL g1962 ( 
.A(n_1919),
.Y(n_1962)
);

INVx1_ASAP7_75t_SL g1963 ( 
.A(n_1898),
.Y(n_1963)
);

AOI22xp5_ASAP7_75t_L g1964 ( 
.A1(n_1940),
.A2(n_1863),
.B1(n_1867),
.B2(n_1871),
.Y(n_1964)
);

INVx1_ASAP7_75t_L g1965 ( 
.A(n_1945),
.Y(n_1965)
);

BUFx8_ASAP7_75t_L g1966 ( 
.A(n_1916),
.Y(n_1966)
);

INVx2_ASAP7_75t_L g1967 ( 
.A(n_1905),
.Y(n_1967)
);

INVx1_ASAP7_75t_L g1968 ( 
.A(n_1934),
.Y(n_1968)
);

INVx1_ASAP7_75t_L g1969 ( 
.A(n_1937),
.Y(n_1969)
);

BUFx6f_ASAP7_75t_L g1970 ( 
.A(n_1930),
.Y(n_1970)
);

INVxp67_ASAP7_75t_SL g1971 ( 
.A(n_1899),
.Y(n_1971)
);

OAI21xp5_ASAP7_75t_L g1972 ( 
.A1(n_1917),
.A2(n_1868),
.B(n_1865),
.Y(n_1972)
);

INVx2_ASAP7_75t_L g1973 ( 
.A(n_1905),
.Y(n_1973)
);

CKINVDCx5p33_ASAP7_75t_R g1974 ( 
.A(n_1898),
.Y(n_1974)
);

OAI22xp5_ASAP7_75t_L g1975 ( 
.A1(n_1926),
.A2(n_1883),
.B1(n_1827),
.B2(n_1832),
.Y(n_1975)
);

INVxp67_ASAP7_75t_L g1976 ( 
.A(n_1951),
.Y(n_1976)
);

OAI22xp5_ASAP7_75t_L g1977 ( 
.A1(n_1964),
.A2(n_1912),
.B1(n_1904),
.B2(n_1925),
.Y(n_1977)
);

HB1xp67_ASAP7_75t_L g1978 ( 
.A(n_1965),
.Y(n_1978)
);

AOI22xp33_ASAP7_75t_L g1979 ( 
.A1(n_1972),
.A2(n_1940),
.B1(n_1920),
.B2(n_1897),
.Y(n_1979)
);

OAI22xp5_ASAP7_75t_L g1980 ( 
.A1(n_1964),
.A2(n_1912),
.B1(n_1946),
.B2(n_1936),
.Y(n_1980)
);

OAI21xp5_ASAP7_75t_L g1981 ( 
.A1(n_1958),
.A2(n_1873),
.B(n_1840),
.Y(n_1981)
);

OAI22xp5_ASAP7_75t_L g1982 ( 
.A1(n_1954),
.A2(n_1953),
.B1(n_1975),
.B2(n_1946),
.Y(n_1982)
);

INVx1_ASAP7_75t_L g1983 ( 
.A(n_1960),
.Y(n_1983)
);

INVx1_ASAP7_75t_L g1984 ( 
.A(n_1960),
.Y(n_1984)
);

INVx3_ASAP7_75t_L g1985 ( 
.A(n_1952),
.Y(n_1985)
);

INVx1_ASAP7_75t_L g1986 ( 
.A(n_1960),
.Y(n_1986)
);

BUFx6f_ASAP7_75t_L g1987 ( 
.A(n_1950),
.Y(n_1987)
);

OAI22xp33_ASAP7_75t_L g1988 ( 
.A1(n_1950),
.A2(n_1936),
.B1(n_1930),
.B2(n_1859),
.Y(n_1988)
);

INVx3_ASAP7_75t_L g1989 ( 
.A(n_1952),
.Y(n_1989)
);

AOI22xp33_ASAP7_75t_SL g1990 ( 
.A1(n_1953),
.A2(n_1907),
.B1(n_1920),
.B2(n_1914),
.Y(n_1990)
);

AOI22xp33_ASAP7_75t_SL g1991 ( 
.A1(n_1953),
.A2(n_1920),
.B1(n_1932),
.B2(n_1897),
.Y(n_1991)
);

AOI22xp33_ASAP7_75t_L g1992 ( 
.A1(n_1962),
.A2(n_1897),
.B1(n_1932),
.B2(n_1930),
.Y(n_1992)
);

BUFx4f_ASAP7_75t_SL g1993 ( 
.A(n_1963),
.Y(n_1993)
);

BUFx4f_ASAP7_75t_SL g1994 ( 
.A(n_1966),
.Y(n_1994)
);

AOI22xp33_ASAP7_75t_SL g1995 ( 
.A1(n_1953),
.A2(n_1887),
.B1(n_1845),
.B2(n_1942),
.Y(n_1995)
);

OAI22xp5_ASAP7_75t_L g1996 ( 
.A1(n_1950),
.A2(n_1901),
.B1(n_1918),
.B2(n_1910),
.Y(n_1996)
);

XNOR2xp5_ASAP7_75t_L g1997 ( 
.A(n_1982),
.B(n_1974),
.Y(n_1997)
);

NAND2xp5_ASAP7_75t_L g1998 ( 
.A(n_1976),
.B(n_1951),
.Y(n_1998)
);

INVx8_ASAP7_75t_L g1999 ( 
.A(n_1987),
.Y(n_1999)
);

AND2x2_ASAP7_75t_L g2000 ( 
.A(n_1987),
.B(n_1949),
.Y(n_2000)
);

INVx2_ASAP7_75t_L g2001 ( 
.A(n_1985),
.Y(n_2001)
);

INVx1_ASAP7_75t_L g2002 ( 
.A(n_1978),
.Y(n_2002)
);

AND2x2_ASAP7_75t_L g2003 ( 
.A(n_1987),
.B(n_1969),
.Y(n_2003)
);

INVx8_ASAP7_75t_L g2004 ( 
.A(n_1987),
.Y(n_2004)
);

NAND2xp33_ASAP7_75t_R g2005 ( 
.A(n_1981),
.B(n_1943),
.Y(n_2005)
);

INVx2_ASAP7_75t_L g2006 ( 
.A(n_1985),
.Y(n_2006)
);

NAND2xp5_ASAP7_75t_L g2007 ( 
.A(n_1998),
.B(n_1980),
.Y(n_2007)
);

NAND2xp5_ASAP7_75t_L g2008 ( 
.A(n_1998),
.B(n_1969),
.Y(n_2008)
);

AND2x2_ASAP7_75t_L g2009 ( 
.A(n_2000),
.B(n_1948),
.Y(n_2009)
);

NAND2xp5_ASAP7_75t_L g2010 ( 
.A(n_2003),
.B(n_1910),
.Y(n_2010)
);

AOI22xp33_ASAP7_75t_L g2011 ( 
.A1(n_1997),
.A2(n_1977),
.B1(n_1990),
.B2(n_1991),
.Y(n_2011)
);

BUFx2_ASAP7_75t_L g2012 ( 
.A(n_1999),
.Y(n_2012)
);

AND2x2_ASAP7_75t_L g2013 ( 
.A(n_2009),
.B(n_2001),
.Y(n_2013)
);

AND2x2_ASAP7_75t_L g2014 ( 
.A(n_2012),
.B(n_2006),
.Y(n_2014)
);

BUFx2_ASAP7_75t_SL g2015 ( 
.A(n_2011),
.Y(n_2015)
);

INVxp67_ASAP7_75t_L g2016 ( 
.A(n_2007),
.Y(n_2016)
);

AND2x4_ASAP7_75t_L g2017 ( 
.A(n_2010),
.B(n_2002),
.Y(n_2017)
);

AOI22xp5_ASAP7_75t_L g2018 ( 
.A1(n_2008),
.A2(n_2005),
.B1(n_1979),
.B2(n_1988),
.Y(n_2018)
);

HB1xp67_ASAP7_75t_L g2019 ( 
.A(n_2012),
.Y(n_2019)
);

NOR2xp33_ASAP7_75t_L g2020 ( 
.A(n_2007),
.B(n_1993),
.Y(n_2020)
);

INVxp67_ASAP7_75t_SL g2021 ( 
.A(n_2007),
.Y(n_2021)
);

OAI22xp5_ASAP7_75t_L g2022 ( 
.A1(n_2011),
.A2(n_1995),
.B1(n_1992),
.B2(n_1988),
.Y(n_2022)
);

AND2x2_ASAP7_75t_L g2023 ( 
.A(n_2019),
.B(n_1916),
.Y(n_2023)
);

HB1xp67_ASAP7_75t_L g2024 ( 
.A(n_2016),
.Y(n_2024)
);

INVx1_ASAP7_75t_L g2025 ( 
.A(n_2017),
.Y(n_2025)
);

OR2x2_ASAP7_75t_L g2026 ( 
.A(n_2021),
.B(n_1906),
.Y(n_2026)
);

HB1xp67_ASAP7_75t_L g2027 ( 
.A(n_2017),
.Y(n_2027)
);

AND2x2_ASAP7_75t_L g2028 ( 
.A(n_2014),
.B(n_2013),
.Y(n_2028)
);

INVx1_ASAP7_75t_L g2029 ( 
.A(n_2015),
.Y(n_2029)
);

NAND2xp5_ASAP7_75t_L g2030 ( 
.A(n_2020),
.B(n_1928),
.Y(n_2030)
);

NAND2xp5_ASAP7_75t_L g2031 ( 
.A(n_2018),
.B(n_1928),
.Y(n_2031)
);

AND2x4_ASAP7_75t_L g2032 ( 
.A(n_2022),
.B(n_1989),
.Y(n_2032)
);

INVx2_ASAP7_75t_L g2033 ( 
.A(n_2022),
.Y(n_2033)
);

AND2x2_ASAP7_75t_L g2034 ( 
.A(n_2028),
.B(n_1938),
.Y(n_2034)
);

NAND2xp5_ASAP7_75t_L g2035 ( 
.A(n_2029),
.B(n_1999),
.Y(n_2035)
);

INVx1_ASAP7_75t_L g2036 ( 
.A(n_2027),
.Y(n_2036)
);

INVx1_ASAP7_75t_L g2037 ( 
.A(n_2027),
.Y(n_2037)
);

NAND2xp5_ASAP7_75t_L g2038 ( 
.A(n_2024),
.B(n_1978),
.Y(n_2038)
);

INVx3_ASAP7_75t_L g2039 ( 
.A(n_2023),
.Y(n_2039)
);

INVx1_ASAP7_75t_L g2040 ( 
.A(n_2024),
.Y(n_2040)
);

OR2x2_ASAP7_75t_L g2041 ( 
.A(n_2025),
.B(n_1999),
.Y(n_2041)
);

AND2x4_ASAP7_75t_L g2042 ( 
.A(n_2026),
.B(n_1684),
.Y(n_2042)
);

NAND2xp5_ASAP7_75t_L g2043 ( 
.A(n_2039),
.B(n_2033),
.Y(n_2043)
);

NOR2xp33_ASAP7_75t_L g2044 ( 
.A(n_2042),
.B(n_2030),
.Y(n_2044)
);

NAND2xp5_ASAP7_75t_L g2045 ( 
.A(n_2039),
.B(n_2033),
.Y(n_2045)
);

OR2x2_ASAP7_75t_L g2046 ( 
.A(n_2040),
.B(n_2031),
.Y(n_2046)
);

AND2x2_ASAP7_75t_L g2047 ( 
.A(n_2044),
.B(n_2034),
.Y(n_2047)
);

INVx1_ASAP7_75t_L g2048 ( 
.A(n_2043),
.Y(n_2048)
);

INVx1_ASAP7_75t_L g2049 ( 
.A(n_2045),
.Y(n_2049)
);

INVx1_ASAP7_75t_L g2050 ( 
.A(n_2046),
.Y(n_2050)
);

INVx1_ASAP7_75t_L g2051 ( 
.A(n_2050),
.Y(n_2051)
);

INVx1_ASAP7_75t_L g2052 ( 
.A(n_2048),
.Y(n_2052)
);

INVx1_ASAP7_75t_SL g2053 ( 
.A(n_2047),
.Y(n_2053)
);

INVx2_ASAP7_75t_SL g2054 ( 
.A(n_2047),
.Y(n_2054)
);

NOR2xp33_ASAP7_75t_L g2055 ( 
.A(n_2049),
.B(n_2042),
.Y(n_2055)
);

AOI22xp5_ASAP7_75t_L g2056 ( 
.A1(n_2047),
.A2(n_2032),
.B1(n_2035),
.B2(n_2036),
.Y(n_2056)
);

INVx1_ASAP7_75t_L g2057 ( 
.A(n_2054),
.Y(n_2057)
);

NOR2xp33_ASAP7_75t_L g2058 ( 
.A(n_2053),
.B(n_2056),
.Y(n_2058)
);

AOI22xp33_ASAP7_75t_L g2059 ( 
.A1(n_2055),
.A2(n_2032),
.B1(n_2037),
.B2(n_2051),
.Y(n_2059)
);

INVx2_ASAP7_75t_SL g2060 ( 
.A(n_2052),
.Y(n_2060)
);

INVxp67_ASAP7_75t_L g2061 ( 
.A(n_2054),
.Y(n_2061)
);

AOI22xp33_ASAP7_75t_SL g2062 ( 
.A1(n_2053),
.A2(n_2038),
.B1(n_2041),
.B2(n_1994),
.Y(n_2062)
);

INVx1_ASAP7_75t_SL g2063 ( 
.A(n_2053),
.Y(n_2063)
);

AOI22xp5_ASAP7_75t_L g2064 ( 
.A1(n_2053),
.A2(n_2038),
.B1(n_2005),
.B2(n_2004),
.Y(n_2064)
);

O2A1O1Ixp33_ASAP7_75t_L g2065 ( 
.A1(n_2054),
.A2(n_1847),
.B(n_1844),
.C(n_1869),
.Y(n_2065)
);

INVx1_ASAP7_75t_L g2066 ( 
.A(n_2054),
.Y(n_2066)
);

A2O1A1Ixp33_ASAP7_75t_L g2067 ( 
.A1(n_2058),
.A2(n_2061),
.B(n_2063),
.C(n_2057),
.Y(n_2067)
);

NAND2xp5_ASAP7_75t_L g2068 ( 
.A(n_2066),
.B(n_1938),
.Y(n_2068)
);

INVx1_ASAP7_75t_L g2069 ( 
.A(n_2060),
.Y(n_2069)
);

NOR2xp33_ASAP7_75t_L g2070 ( 
.A(n_2059),
.B(n_1814),
.Y(n_2070)
);

O2A1O1Ixp33_ASAP7_75t_L g2071 ( 
.A1(n_2065),
.A2(n_1848),
.B(n_1861),
.C(n_1842),
.Y(n_2071)
);

INVx1_ASAP7_75t_L g2072 ( 
.A(n_2062),
.Y(n_2072)
);

INVx1_ASAP7_75t_L g2073 ( 
.A(n_2064),
.Y(n_2073)
);

INVx1_ASAP7_75t_L g2074 ( 
.A(n_2057),
.Y(n_2074)
);

OAI321xp33_ASAP7_75t_L g2075 ( 
.A1(n_2061),
.A2(n_1996),
.A3(n_1901),
.B1(n_1827),
.B2(n_1948),
.C(n_1970),
.Y(n_2075)
);

OAI22xp5_ASAP7_75t_L g2076 ( 
.A1(n_2059),
.A2(n_2004),
.B1(n_1821),
.B2(n_1962),
.Y(n_2076)
);

O2A1O1Ixp33_ASAP7_75t_L g2077 ( 
.A1(n_2061),
.A2(n_1855),
.B(n_1836),
.C(n_1843),
.Y(n_2077)
);

AND2x2_ASAP7_75t_L g2078 ( 
.A(n_2063),
.B(n_2004),
.Y(n_2078)
);

INVx1_ASAP7_75t_L g2079 ( 
.A(n_2057),
.Y(n_2079)
);

NOR2xp67_ASAP7_75t_SL g2080 ( 
.A(n_2069),
.B(n_1743),
.Y(n_2080)
);

INVx2_ASAP7_75t_L g2081 ( 
.A(n_2078),
.Y(n_2081)
);

AO22x2_ASAP7_75t_L g2082 ( 
.A1(n_2074),
.A2(n_2079),
.B1(n_2072),
.B2(n_2073),
.Y(n_2082)
);

NOR3xp33_ASAP7_75t_SL g2083 ( 
.A(n_2067),
.B(n_1834),
.C(n_1935),
.Y(n_2083)
);

NAND2xp5_ASAP7_75t_L g2084 ( 
.A(n_2070),
.B(n_1983),
.Y(n_2084)
);

INVx1_ASAP7_75t_L g2085 ( 
.A(n_2068),
.Y(n_2085)
);

NAND2xp5_ASAP7_75t_L g2086 ( 
.A(n_2076),
.B(n_1984),
.Y(n_2086)
);

NAND2xp5_ASAP7_75t_L g2087 ( 
.A(n_2071),
.B(n_1986),
.Y(n_2087)
);

NOR2xp33_ASAP7_75t_L g2088 ( 
.A(n_2075),
.B(n_1966),
.Y(n_2088)
);

AND2x2_ASAP7_75t_L g2089 ( 
.A(n_2077),
.B(n_1922),
.Y(n_2089)
);

INVx1_ASAP7_75t_L g2090 ( 
.A(n_2074),
.Y(n_2090)
);

INVx1_ASAP7_75t_L g2091 ( 
.A(n_2074),
.Y(n_2091)
);

AOI21xp5_ASAP7_75t_L g2092 ( 
.A1(n_2067),
.A2(n_1923),
.B(n_1866),
.Y(n_2092)
);

HB1xp67_ASAP7_75t_L g2093 ( 
.A(n_2078),
.Y(n_2093)
);

NOR3xp33_ASAP7_75t_L g2094 ( 
.A(n_2067),
.B(n_1866),
.C(n_1875),
.Y(n_2094)
);

OA21x2_ASAP7_75t_L g2095 ( 
.A1(n_2090),
.A2(n_2091),
.B(n_2081),
.Y(n_2095)
);

AOI221x1_ASAP7_75t_L g2096 ( 
.A1(n_2082),
.A2(n_1748),
.B1(n_199),
.B2(n_200),
.C(n_201),
.Y(n_2096)
);

AOI211xp5_ASAP7_75t_L g2097 ( 
.A1(n_2093),
.A2(n_2088),
.B(n_2085),
.C(n_2080),
.Y(n_2097)
);

OAI211xp5_ASAP7_75t_L g2098 ( 
.A1(n_2086),
.A2(n_1748),
.B(n_1864),
.C(n_200),
.Y(n_2098)
);

AOI221xp5_ASAP7_75t_L g2099 ( 
.A1(n_2082),
.A2(n_1839),
.B1(n_1893),
.B2(n_1782),
.C(n_1971),
.Y(n_2099)
);

AOI221xp5_ASAP7_75t_L g2100 ( 
.A1(n_2094),
.A2(n_1782),
.B1(n_1970),
.B2(n_1948),
.C(n_1965),
.Y(n_2100)
);

OAI21xp5_ASAP7_75t_L g2101 ( 
.A1(n_2092),
.A2(n_1887),
.B(n_1837),
.Y(n_2101)
);

OAI221xp5_ASAP7_75t_SL g2102 ( 
.A1(n_2084),
.A2(n_1887),
.B1(n_1966),
.B2(n_1922),
.C(n_1908),
.Y(n_2102)
);

AOI221xp5_ASAP7_75t_L g2103 ( 
.A1(n_2083),
.A2(n_1970),
.B1(n_1948),
.B2(n_1989),
.C(n_1968),
.Y(n_2103)
);

OAI21xp33_ASAP7_75t_L g2104 ( 
.A1(n_2089),
.A2(n_1970),
.B(n_1948),
.Y(n_2104)
);

OAI21xp33_ASAP7_75t_SL g2105 ( 
.A1(n_2087),
.A2(n_1966),
.B(n_1968),
.Y(n_2105)
);

AOI21xp33_ASAP7_75t_L g2106 ( 
.A1(n_2093),
.A2(n_198),
.B(n_199),
.Y(n_2106)
);

AOI221xp5_ASAP7_75t_L g2107 ( 
.A1(n_2082),
.A2(n_1970),
.B1(n_1948),
.B2(n_203),
.C(n_205),
.Y(n_2107)
);

AOI21xp5_ASAP7_75t_L g2108 ( 
.A1(n_2093),
.A2(n_1943),
.B(n_1896),
.Y(n_2108)
);

AOI22xp5_ASAP7_75t_L g2109 ( 
.A1(n_2107),
.A2(n_2097),
.B1(n_2104),
.B2(n_2099),
.Y(n_2109)
);

AOI211xp5_ASAP7_75t_L g2110 ( 
.A1(n_2098),
.A2(n_205),
.B(n_198),
.C(n_202),
.Y(n_2110)
);

OAI221xp5_ASAP7_75t_L g2111 ( 
.A1(n_2105),
.A2(n_1970),
.B1(n_1943),
.B2(n_1957),
.C(n_1913),
.Y(n_2111)
);

NAND2xp5_ASAP7_75t_L g2112 ( 
.A(n_2096),
.B(n_202),
.Y(n_2112)
);

NAND2xp5_ASAP7_75t_L g2113 ( 
.A(n_2095),
.B(n_206),
.Y(n_2113)
);

NOR2x1_ASAP7_75t_L g2114 ( 
.A(n_2095),
.B(n_206),
.Y(n_2114)
);

NAND2xp5_ASAP7_75t_SL g2115 ( 
.A(n_2106),
.B(n_1829),
.Y(n_2115)
);

AOI22xp5_ASAP7_75t_L g2116 ( 
.A1(n_2100),
.A2(n_1939),
.B1(n_1944),
.B2(n_1941),
.Y(n_2116)
);

OAI221xp5_ASAP7_75t_L g2117 ( 
.A1(n_2103),
.A2(n_1957),
.B1(n_1903),
.B2(n_1967),
.C(n_1973),
.Y(n_2117)
);

OAI211xp5_ASAP7_75t_SL g2118 ( 
.A1(n_2101),
.A2(n_210),
.B(n_207),
.C(n_209),
.Y(n_2118)
);

AOI22xp5_ASAP7_75t_L g2119 ( 
.A1(n_2108),
.A2(n_1939),
.B1(n_1944),
.B2(n_1941),
.Y(n_2119)
);

AOI221xp5_ASAP7_75t_L g2120 ( 
.A1(n_2102),
.A2(n_207),
.B1(n_211),
.B2(n_212),
.C(n_213),
.Y(n_2120)
);

OR2x2_ASAP7_75t_L g2121 ( 
.A(n_2095),
.B(n_211),
.Y(n_2121)
);

AND2x2_ASAP7_75t_L g2122 ( 
.A(n_2095),
.B(n_1929),
.Y(n_2122)
);

AOI21xp33_ASAP7_75t_SL g2123 ( 
.A1(n_2095),
.A2(n_212),
.B(n_213),
.Y(n_2123)
);

OAI21xp5_ASAP7_75t_L g2124 ( 
.A1(n_2105),
.A2(n_1884),
.B(n_1921),
.Y(n_2124)
);

OAI21xp5_ASAP7_75t_SL g2125 ( 
.A1(n_2107),
.A2(n_214),
.B(n_215),
.Y(n_2125)
);

OAI221xp5_ASAP7_75t_L g2126 ( 
.A1(n_2107),
.A2(n_1957),
.B1(n_1967),
.B2(n_1973),
.C(n_1829),
.Y(n_2126)
);

AOI211xp5_ASAP7_75t_L g2127 ( 
.A1(n_2107),
.A2(n_214),
.B(n_215),
.C(n_216),
.Y(n_2127)
);

NAND3xp33_ASAP7_75t_L g2128 ( 
.A(n_2096),
.B(n_216),
.C(n_217),
.Y(n_2128)
);

AOI221x1_ASAP7_75t_L g2129 ( 
.A1(n_2106),
.A2(n_218),
.B1(n_219),
.B2(n_220),
.C(n_221),
.Y(n_2129)
);

OAI211xp5_ASAP7_75t_L g2130 ( 
.A1(n_2123),
.A2(n_220),
.B(n_221),
.C(n_222),
.Y(n_2130)
);

AOI322xp5_ASAP7_75t_L g2131 ( 
.A1(n_2114),
.A2(n_1956),
.A3(n_1955),
.B1(n_1927),
.B2(n_1947),
.C1(n_1961),
.C2(n_1959),
.Y(n_2131)
);

AND2x2_ASAP7_75t_L g2132 ( 
.A(n_2122),
.B(n_1956),
.Y(n_2132)
);

AOI21xp33_ASAP7_75t_SL g2133 ( 
.A1(n_2128),
.A2(n_2112),
.B(n_2121),
.Y(n_2133)
);

NAND2xp5_ASAP7_75t_L g2134 ( 
.A(n_2129),
.B(n_222),
.Y(n_2134)
);

NOR3xp33_ASAP7_75t_L g2135 ( 
.A(n_2125),
.B(n_223),
.C(n_224),
.Y(n_2135)
);

AOI22xp5_ASAP7_75t_L g2136 ( 
.A1(n_2109),
.A2(n_1956),
.B1(n_1927),
.B2(n_1933),
.Y(n_2136)
);

NOR2xp33_ASAP7_75t_L g2137 ( 
.A(n_2118),
.B(n_224),
.Y(n_2137)
);

A2O1A1Ixp33_ASAP7_75t_L g2138 ( 
.A1(n_2120),
.A2(n_225),
.B(n_226),
.C(n_227),
.Y(n_2138)
);

INVx1_ASAP7_75t_L g2139 ( 
.A(n_2113),
.Y(n_2139)
);

INVx1_ASAP7_75t_L g2140 ( 
.A(n_2127),
.Y(n_2140)
);

AOI221xp5_ASAP7_75t_SL g2141 ( 
.A1(n_2126),
.A2(n_225),
.B1(n_226),
.B2(n_227),
.C(n_228),
.Y(n_2141)
);

AOI221xp5_ASAP7_75t_SL g2142 ( 
.A1(n_2110),
.A2(n_228),
.B1(n_229),
.B2(n_230),
.C(n_231),
.Y(n_2142)
);

XNOR2xp5_ASAP7_75t_L g2143 ( 
.A(n_2115),
.B(n_229),
.Y(n_2143)
);

OAI221xp5_ASAP7_75t_L g2144 ( 
.A1(n_2111),
.A2(n_230),
.B1(n_231),
.B2(n_232),
.C(n_233),
.Y(n_2144)
);

AOI211xp5_ASAP7_75t_L g2145 ( 
.A1(n_2117),
.A2(n_232),
.B(n_233),
.C(n_234),
.Y(n_2145)
);

NOR4xp25_ASAP7_75t_L g2146 ( 
.A(n_2124),
.B(n_234),
.C(n_235),
.D(n_236),
.Y(n_2146)
);

INVx1_ASAP7_75t_L g2147 ( 
.A(n_2119),
.Y(n_2147)
);

NAND2xp5_ASAP7_75t_L g2148 ( 
.A(n_2116),
.B(n_235),
.Y(n_2148)
);

AOI221xp5_ASAP7_75t_L g2149 ( 
.A1(n_2123),
.A2(n_236),
.B1(n_237),
.B2(n_238),
.C(n_239),
.Y(n_2149)
);

NAND2xp5_ASAP7_75t_L g2150 ( 
.A(n_2122),
.B(n_240),
.Y(n_2150)
);

OAI211xp5_ASAP7_75t_L g2151 ( 
.A1(n_2123),
.A2(n_241),
.B(n_242),
.C(n_243),
.Y(n_2151)
);

AOI21xp5_ASAP7_75t_L g2152 ( 
.A1(n_2113),
.A2(n_241),
.B(n_242),
.Y(n_2152)
);

AOI322xp5_ASAP7_75t_L g2153 ( 
.A1(n_2114),
.A2(n_1956),
.A3(n_1955),
.B1(n_1927),
.B2(n_1947),
.C1(n_1961),
.C2(n_1959),
.Y(n_2153)
);

AOI211xp5_ASAP7_75t_L g2154 ( 
.A1(n_2123),
.A2(n_243),
.B(n_244),
.C(n_245),
.Y(n_2154)
);

AND3x1_ASAP7_75t_L g2155 ( 
.A(n_2127),
.B(n_244),
.C(n_246),
.Y(n_2155)
);

O2A1O1Ixp5_ASAP7_75t_L g2156 ( 
.A1(n_2113),
.A2(n_247),
.B(n_248),
.C(n_249),
.Y(n_2156)
);

NOR4xp25_ASAP7_75t_L g2157 ( 
.A(n_2113),
.B(n_247),
.C(n_248),
.D(n_249),
.Y(n_2157)
);

NAND4xp25_ASAP7_75t_L g2158 ( 
.A(n_2120),
.B(n_250),
.C(n_251),
.D(n_252),
.Y(n_2158)
);

AOI211xp5_ASAP7_75t_L g2159 ( 
.A1(n_2123),
.A2(n_250),
.B(n_253),
.C(n_254),
.Y(n_2159)
);

INVx3_ASAP7_75t_L g2160 ( 
.A(n_2121),
.Y(n_2160)
);

AOI211x1_ASAP7_75t_SL g2161 ( 
.A1(n_2118),
.A2(n_253),
.B(n_254),
.C(n_255),
.Y(n_2161)
);

AOI211xp5_ASAP7_75t_L g2162 ( 
.A1(n_2123),
.A2(n_255),
.B(n_257),
.C(n_258),
.Y(n_2162)
);

AOI221x1_ASAP7_75t_L g2163 ( 
.A1(n_2123),
.A2(n_257),
.B1(n_259),
.B2(n_260),
.C(n_261),
.Y(n_2163)
);

HB1xp67_ASAP7_75t_L g2164 ( 
.A(n_2134),
.Y(n_2164)
);

NOR2x1_ASAP7_75t_L g2165 ( 
.A(n_2160),
.B(n_259),
.Y(n_2165)
);

NOR2x1_ASAP7_75t_L g2166 ( 
.A(n_2160),
.B(n_260),
.Y(n_2166)
);

NAND2xp5_ASAP7_75t_L g2167 ( 
.A(n_2157),
.B(n_262),
.Y(n_2167)
);

INVx1_ASAP7_75t_L g2168 ( 
.A(n_2150),
.Y(n_2168)
);

NAND3xp33_ASAP7_75t_L g2169 ( 
.A(n_2154),
.B(n_262),
.C(n_263),
.Y(n_2169)
);

NAND4xp75_ASAP7_75t_L g2170 ( 
.A(n_2142),
.B(n_263),
.C(n_264),
.D(n_265),
.Y(n_2170)
);

HB1xp67_ASAP7_75t_L g2171 ( 
.A(n_2163),
.Y(n_2171)
);

INVx1_ASAP7_75t_L g2172 ( 
.A(n_2130),
.Y(n_2172)
);

NOR2x1_ASAP7_75t_L g2173 ( 
.A(n_2151),
.B(n_264),
.Y(n_2173)
);

NAND4xp75_ASAP7_75t_L g2174 ( 
.A(n_2155),
.B(n_266),
.C(n_268),
.D(n_269),
.Y(n_2174)
);

NOR4xp75_ASAP7_75t_L g2175 ( 
.A(n_2144),
.B(n_268),
.C(n_269),
.D(n_270),
.Y(n_2175)
);

INVx1_ASAP7_75t_L g2176 ( 
.A(n_2143),
.Y(n_2176)
);

NAND4xp75_ASAP7_75t_L g2177 ( 
.A(n_2140),
.B(n_271),
.C(n_272),
.D(n_273),
.Y(n_2177)
);

XNOR2xp5_ASAP7_75t_L g2178 ( 
.A(n_2161),
.B(n_271),
.Y(n_2178)
);

INVx1_ASAP7_75t_L g2179 ( 
.A(n_2156),
.Y(n_2179)
);

INVx1_ASAP7_75t_L g2180 ( 
.A(n_2137),
.Y(n_2180)
);

NOR2xp33_ASAP7_75t_L g2181 ( 
.A(n_2158),
.B(n_272),
.Y(n_2181)
);

INVx1_ASAP7_75t_L g2182 ( 
.A(n_2148),
.Y(n_2182)
);

AND2x2_ASAP7_75t_L g2183 ( 
.A(n_2132),
.B(n_1947),
.Y(n_2183)
);

NOR2xp33_ASAP7_75t_L g2184 ( 
.A(n_2133),
.B(n_274),
.Y(n_2184)
);

NOR2xp33_ASAP7_75t_L g2185 ( 
.A(n_2139),
.B(n_274),
.Y(n_2185)
);

INVx1_ASAP7_75t_L g2186 ( 
.A(n_2159),
.Y(n_2186)
);

NAND4xp75_ASAP7_75t_L g2187 ( 
.A(n_2152),
.B(n_275),
.C(n_276),
.D(n_277),
.Y(n_2187)
);

INVx1_ASAP7_75t_L g2188 ( 
.A(n_2162),
.Y(n_2188)
);

OA21x2_ASAP7_75t_L g2189 ( 
.A1(n_2147),
.A2(n_275),
.B(n_276),
.Y(n_2189)
);

NOR2x1_ASAP7_75t_L g2190 ( 
.A(n_2138),
.B(n_277),
.Y(n_2190)
);

NOR2x1_ASAP7_75t_L g2191 ( 
.A(n_2149),
.B(n_2146),
.Y(n_2191)
);

INVxp33_ASAP7_75t_L g2192 ( 
.A(n_2178),
.Y(n_2192)
);

INVx1_ASAP7_75t_L g2193 ( 
.A(n_2165),
.Y(n_2193)
);

OR2x2_ASAP7_75t_L g2194 ( 
.A(n_2167),
.B(n_2135),
.Y(n_2194)
);

AOI31xp33_ASAP7_75t_L g2195 ( 
.A1(n_2171),
.A2(n_2141),
.A3(n_2145),
.B(n_2136),
.Y(n_2195)
);

NOR2x1_ASAP7_75t_L g2196 ( 
.A(n_2166),
.B(n_2131),
.Y(n_2196)
);

XNOR2xp5_ASAP7_75t_L g2197 ( 
.A(n_2175),
.B(n_278),
.Y(n_2197)
);

NOR2x1_ASAP7_75t_L g2198 ( 
.A(n_2177),
.B(n_2153),
.Y(n_2198)
);

INVx1_ASAP7_75t_L g2199 ( 
.A(n_2189),
.Y(n_2199)
);

BUFx12f_ASAP7_75t_L g2200 ( 
.A(n_2164),
.Y(n_2200)
);

NAND4xp75_ASAP7_75t_L g2201 ( 
.A(n_2184),
.B(n_279),
.C(n_280),
.D(n_281),
.Y(n_2201)
);

AND3x4_ASAP7_75t_L g2202 ( 
.A(n_2173),
.B(n_2191),
.C(n_2190),
.Y(n_2202)
);

INVxp67_ASAP7_75t_L g2203 ( 
.A(n_2185),
.Y(n_2203)
);

INVx2_ASAP7_75t_L g2204 ( 
.A(n_2189),
.Y(n_2204)
);

NOR3xp33_ASAP7_75t_L g2205 ( 
.A(n_2179),
.B(n_279),
.C(n_280),
.Y(n_2205)
);

INVx2_ASAP7_75t_L g2206 ( 
.A(n_2174),
.Y(n_2206)
);

INVx2_ASAP7_75t_SL g2207 ( 
.A(n_2176),
.Y(n_2207)
);

NOR3xp33_ASAP7_75t_L g2208 ( 
.A(n_2172),
.B(n_282),
.C(n_283),
.Y(n_2208)
);

AND2x4_ASAP7_75t_L g2209 ( 
.A(n_2168),
.B(n_282),
.Y(n_2209)
);

AND2x2_ASAP7_75t_L g2210 ( 
.A(n_2181),
.B(n_1947),
.Y(n_2210)
);

INVx3_ASAP7_75t_L g2211 ( 
.A(n_2187),
.Y(n_2211)
);

NOR3xp33_ASAP7_75t_L g2212 ( 
.A(n_2186),
.B(n_283),
.C(n_284),
.Y(n_2212)
);

CKINVDCx5p33_ASAP7_75t_R g2213 ( 
.A(n_2180),
.Y(n_2213)
);

INVx1_ASAP7_75t_L g2214 ( 
.A(n_2170),
.Y(n_2214)
);

NAND3x1_ASAP7_75t_L g2215 ( 
.A(n_2188),
.B(n_284),
.C(n_285),
.Y(n_2215)
);

INVx1_ASAP7_75t_L g2216 ( 
.A(n_2169),
.Y(n_2216)
);

NOR2xp33_ASAP7_75t_L g2217 ( 
.A(n_2182),
.B(n_285),
.Y(n_2217)
);

NOR3xp33_ASAP7_75t_L g2218 ( 
.A(n_2183),
.B(n_286),
.C(n_287),
.Y(n_2218)
);

NAND3x2_ASAP7_75t_L g2219 ( 
.A(n_2172),
.B(n_286),
.C(n_287),
.Y(n_2219)
);

AND2x4_ASAP7_75t_L g2220 ( 
.A(n_2165),
.B(n_289),
.Y(n_2220)
);

INVx1_ASAP7_75t_L g2221 ( 
.A(n_2165),
.Y(n_2221)
);

HB1xp67_ASAP7_75t_L g2222 ( 
.A(n_2189),
.Y(n_2222)
);

NAND2xp5_ASAP7_75t_L g2223 ( 
.A(n_2185),
.B(n_289),
.Y(n_2223)
);

NOR2x1p5_ASAP7_75t_L g2224 ( 
.A(n_2170),
.B(n_290),
.Y(n_2224)
);

NAND2x1p5_ASAP7_75t_L g2225 ( 
.A(n_2165),
.B(n_290),
.Y(n_2225)
);

NOR3x1_ASAP7_75t_L g2226 ( 
.A(n_2174),
.B(n_291),
.C(n_292),
.Y(n_2226)
);

AND3x4_ASAP7_75t_L g2227 ( 
.A(n_2175),
.B(n_293),
.C(n_294),
.Y(n_2227)
);

INVx1_ASAP7_75t_L g2228 ( 
.A(n_2222),
.Y(n_2228)
);

XNOR2x1_ASAP7_75t_L g2229 ( 
.A(n_2227),
.B(n_294),
.Y(n_2229)
);

INVx1_ASAP7_75t_L g2230 ( 
.A(n_2199),
.Y(n_2230)
);

HB1xp67_ASAP7_75t_L g2231 ( 
.A(n_2204),
.Y(n_2231)
);

NAND2xp5_ASAP7_75t_L g2232 ( 
.A(n_2220),
.B(n_295),
.Y(n_2232)
);

OAI221xp5_ASAP7_75t_L g2233 ( 
.A1(n_2225),
.A2(n_295),
.B1(n_296),
.B2(n_297),
.C(n_298),
.Y(n_2233)
);

AOI22xp33_ASAP7_75t_SL g2234 ( 
.A1(n_2200),
.A2(n_1952),
.B1(n_298),
.B2(n_299),
.Y(n_2234)
);

NOR3x1_ASAP7_75t_L g2235 ( 
.A(n_2201),
.B(n_297),
.C(n_299),
.Y(n_2235)
);

OAI31xp33_ASAP7_75t_L g2236 ( 
.A1(n_2224),
.A2(n_300),
.A3(n_302),
.B(n_303),
.Y(n_2236)
);

NAND2xp5_ASAP7_75t_L g2237 ( 
.A(n_2197),
.B(n_302),
.Y(n_2237)
);

INVx1_ASAP7_75t_L g2238 ( 
.A(n_2197),
.Y(n_2238)
);

INVx1_ASAP7_75t_L g2239 ( 
.A(n_2215),
.Y(n_2239)
);

NOR4xp25_ASAP7_75t_L g2240 ( 
.A(n_2214),
.B(n_303),
.C(n_304),
.D(n_305),
.Y(n_2240)
);

OR2x2_ASAP7_75t_L g2241 ( 
.A(n_2219),
.B(n_304),
.Y(n_2241)
);

NAND3x1_ASAP7_75t_SL g2242 ( 
.A(n_2196),
.B(n_305),
.C(n_306),
.Y(n_2242)
);

CKINVDCx16_ASAP7_75t_R g2243 ( 
.A(n_2194),
.Y(n_2243)
);

NAND2xp5_ASAP7_75t_L g2244 ( 
.A(n_2218),
.B(n_307),
.Y(n_2244)
);

AND2x4_ASAP7_75t_L g2245 ( 
.A(n_2193),
.B(n_307),
.Y(n_2245)
);

OAI221xp5_ASAP7_75t_L g2246 ( 
.A1(n_2205),
.A2(n_308),
.B1(n_309),
.B2(n_310),
.C(n_311),
.Y(n_2246)
);

NAND4xp75_ASAP7_75t_L g2247 ( 
.A(n_2226),
.B(n_308),
.C(n_309),
.D(n_311),
.Y(n_2247)
);

OR2x2_ASAP7_75t_L g2248 ( 
.A(n_2221),
.B(n_312),
.Y(n_2248)
);

OAI221xp5_ASAP7_75t_L g2249 ( 
.A1(n_2207),
.A2(n_312),
.B1(n_313),
.B2(n_314),
.C(n_315),
.Y(n_2249)
);

OR2x2_ASAP7_75t_L g2250 ( 
.A(n_2223),
.B(n_313),
.Y(n_2250)
);

NAND2xp5_ASAP7_75t_L g2251 ( 
.A(n_2212),
.B(n_2208),
.Y(n_2251)
);

BUFx3_ASAP7_75t_L g2252 ( 
.A(n_2202),
.Y(n_2252)
);

OAI311xp33_ASAP7_75t_L g2253 ( 
.A1(n_2211),
.A2(n_2216),
.A3(n_2203),
.B1(n_2210),
.C1(n_2195),
.Y(n_2253)
);

HB1xp67_ASAP7_75t_L g2254 ( 
.A(n_2209),
.Y(n_2254)
);

NOR3xp33_ASAP7_75t_L g2255 ( 
.A(n_2206),
.B(n_314),
.C(n_316),
.Y(n_2255)
);

BUFx2_ASAP7_75t_L g2256 ( 
.A(n_2198),
.Y(n_2256)
);

NAND3xp33_ASAP7_75t_L g2257 ( 
.A(n_2236),
.B(n_2213),
.C(n_2192),
.Y(n_2257)
);

NAND2xp33_ASAP7_75t_SL g2258 ( 
.A(n_2239),
.B(n_2229),
.Y(n_2258)
);

NAND3xp33_ASAP7_75t_L g2259 ( 
.A(n_2255),
.B(n_2256),
.C(n_2237),
.Y(n_2259)
);

NAND2xp33_ASAP7_75t_SL g2260 ( 
.A(n_2232),
.B(n_2217),
.Y(n_2260)
);

NAND2xp5_ASAP7_75t_L g2261 ( 
.A(n_2240),
.B(n_317),
.Y(n_2261)
);

NAND2xp33_ASAP7_75t_SL g2262 ( 
.A(n_2241),
.B(n_317),
.Y(n_2262)
);

NAND2xp5_ASAP7_75t_SL g2263 ( 
.A(n_2234),
.B(n_2243),
.Y(n_2263)
);

NAND2xp5_ASAP7_75t_SL g2264 ( 
.A(n_2252),
.B(n_318),
.Y(n_2264)
);

NAND2xp33_ASAP7_75t_SL g2265 ( 
.A(n_2250),
.B(n_318),
.Y(n_2265)
);

XNOR2x1_ASAP7_75t_L g2266 ( 
.A(n_2247),
.B(n_319),
.Y(n_2266)
);

XNOR2xp5_ASAP7_75t_L g2267 ( 
.A(n_2242),
.B(n_319),
.Y(n_2267)
);

NOR2xp33_ASAP7_75t_R g2268 ( 
.A(n_2238),
.B(n_320),
.Y(n_2268)
);

NAND2xp33_ASAP7_75t_SL g2269 ( 
.A(n_2244),
.B(n_321),
.Y(n_2269)
);

NAND2xp33_ASAP7_75t_SL g2270 ( 
.A(n_2254),
.B(n_321),
.Y(n_2270)
);

NAND2xp5_ASAP7_75t_SL g2271 ( 
.A(n_2228),
.B(n_322),
.Y(n_2271)
);

NAND2xp5_ASAP7_75t_L g2272 ( 
.A(n_2231),
.B(n_323),
.Y(n_2272)
);

NAND2xp5_ASAP7_75t_SL g2273 ( 
.A(n_2230),
.B(n_323),
.Y(n_2273)
);

XNOR2x1_ASAP7_75t_L g2274 ( 
.A(n_2251),
.B(n_324),
.Y(n_2274)
);

NOR2xp33_ASAP7_75t_L g2275 ( 
.A(n_2233),
.B(n_324),
.Y(n_2275)
);

NAND2xp5_ASAP7_75t_SL g2276 ( 
.A(n_2248),
.B(n_325),
.Y(n_2276)
);

NOR2xp33_ASAP7_75t_R g2277 ( 
.A(n_2245),
.B(n_325),
.Y(n_2277)
);

NAND3xp33_ASAP7_75t_L g2278 ( 
.A(n_2246),
.B(n_326),
.C(n_327),
.Y(n_2278)
);

NAND2xp5_ASAP7_75t_L g2279 ( 
.A(n_2235),
.B(n_326),
.Y(n_2279)
);

NOR2xp33_ASAP7_75t_L g2280 ( 
.A(n_2249),
.B(n_328),
.Y(n_2280)
);

NOR2xp33_ASAP7_75t_R g2281 ( 
.A(n_2245),
.B(n_328),
.Y(n_2281)
);

NAND2xp33_ASAP7_75t_SL g2282 ( 
.A(n_2253),
.B(n_329),
.Y(n_2282)
);

NAND2xp5_ASAP7_75t_SL g2283 ( 
.A(n_2240),
.B(n_329),
.Y(n_2283)
);

NAND2xp5_ASAP7_75t_L g2284 ( 
.A(n_2240),
.B(n_330),
.Y(n_2284)
);

NOR2xp33_ASAP7_75t_R g2285 ( 
.A(n_2239),
.B(n_330),
.Y(n_2285)
);

XNOR2xp5_ASAP7_75t_L g2286 ( 
.A(n_2229),
.B(n_331),
.Y(n_2286)
);

INVx1_ASAP7_75t_L g2287 ( 
.A(n_2272),
.Y(n_2287)
);

INVx1_ASAP7_75t_L g2288 ( 
.A(n_2267),
.Y(n_2288)
);

INVx1_ASAP7_75t_SL g2289 ( 
.A(n_2277),
.Y(n_2289)
);

INVx1_ASAP7_75t_L g2290 ( 
.A(n_2274),
.Y(n_2290)
);

INVx1_ASAP7_75t_L g2291 ( 
.A(n_2261),
.Y(n_2291)
);

INVx1_ASAP7_75t_L g2292 ( 
.A(n_2284),
.Y(n_2292)
);

OAI22xp5_ASAP7_75t_L g2293 ( 
.A1(n_2259),
.A2(n_2279),
.B1(n_2257),
.B2(n_2278),
.Y(n_2293)
);

NAND2x1_ASAP7_75t_L g2294 ( 
.A(n_2275),
.B(n_331),
.Y(n_2294)
);

AND3x4_ASAP7_75t_L g2295 ( 
.A(n_2282),
.B(n_332),
.C(n_333),
.Y(n_2295)
);

INVx1_ASAP7_75t_L g2296 ( 
.A(n_2266),
.Y(n_2296)
);

INVx1_ASAP7_75t_L g2297 ( 
.A(n_2286),
.Y(n_2297)
);

BUFx4f_ASAP7_75t_SL g2298 ( 
.A(n_2263),
.Y(n_2298)
);

AOI22xp5_ASAP7_75t_L g2299 ( 
.A1(n_2258),
.A2(n_2270),
.B1(n_2262),
.B2(n_2280),
.Y(n_2299)
);

INVx1_ASAP7_75t_L g2300 ( 
.A(n_2264),
.Y(n_2300)
);

AOI22xp5_ASAP7_75t_L g2301 ( 
.A1(n_2265),
.A2(n_1933),
.B1(n_333),
.B2(n_334),
.Y(n_2301)
);

AOI22xp5_ASAP7_75t_L g2302 ( 
.A1(n_2260),
.A2(n_332),
.B1(n_334),
.B2(n_335),
.Y(n_2302)
);

INVx1_ASAP7_75t_L g2303 ( 
.A(n_2273),
.Y(n_2303)
);

INVx1_ASAP7_75t_L g2304 ( 
.A(n_2271),
.Y(n_2304)
);

OA22x2_ASAP7_75t_L g2305 ( 
.A1(n_2283),
.A2(n_336),
.B1(n_337),
.B2(n_338),
.Y(n_2305)
);

XNOR2x1_ASAP7_75t_L g2306 ( 
.A(n_2295),
.B(n_2281),
.Y(n_2306)
);

AO22x2_ASAP7_75t_L g2307 ( 
.A1(n_2289),
.A2(n_2276),
.B1(n_2285),
.B2(n_2269),
.Y(n_2307)
);

INVx1_ASAP7_75t_L g2308 ( 
.A(n_2305),
.Y(n_2308)
);

INVx1_ASAP7_75t_L g2309 ( 
.A(n_2294),
.Y(n_2309)
);

XNOR2xp5_ASAP7_75t_L g2310 ( 
.A(n_2293),
.B(n_2268),
.Y(n_2310)
);

NOR2xp33_ASAP7_75t_L g2311 ( 
.A(n_2298),
.B(n_337),
.Y(n_2311)
);

AOI22xp5_ASAP7_75t_L g2312 ( 
.A1(n_2288),
.A2(n_338),
.B1(n_339),
.B2(n_340),
.Y(n_2312)
);

INVx1_ASAP7_75t_L g2313 ( 
.A(n_2299),
.Y(n_2313)
);

INVx2_ASAP7_75t_L g2314 ( 
.A(n_2291),
.Y(n_2314)
);

NAND2xp5_ASAP7_75t_L g2315 ( 
.A(n_2302),
.B(n_339),
.Y(n_2315)
);

HB1xp67_ASAP7_75t_L g2316 ( 
.A(n_2304),
.Y(n_2316)
);

INVxp67_ASAP7_75t_L g2317 ( 
.A(n_2300),
.Y(n_2317)
);

AOI21xp5_ASAP7_75t_L g2318 ( 
.A1(n_2306),
.A2(n_2303),
.B(n_2290),
.Y(n_2318)
);

NOR3x1_ASAP7_75t_L g2319 ( 
.A(n_2313),
.B(n_2296),
.C(n_2292),
.Y(n_2319)
);

AOI22x1_ASAP7_75t_L g2320 ( 
.A1(n_2316),
.A2(n_2297),
.B1(n_2287),
.B2(n_2301),
.Y(n_2320)
);

OAI22x1_ASAP7_75t_L g2321 ( 
.A1(n_2310),
.A2(n_340),
.B1(n_341),
.B2(n_342),
.Y(n_2321)
);

NAND2xp5_ASAP7_75t_L g2322 ( 
.A(n_2311),
.B(n_341),
.Y(n_2322)
);

OR2x2_ASAP7_75t_SL g2323 ( 
.A(n_2315),
.B(n_342),
.Y(n_2323)
);

OAI22xp5_ASAP7_75t_SL g2324 ( 
.A1(n_2309),
.A2(n_343),
.B1(n_344),
.B2(n_345),
.Y(n_2324)
);

INVx1_ASAP7_75t_L g2325 ( 
.A(n_2307),
.Y(n_2325)
);

OR3x1_ASAP7_75t_L g2326 ( 
.A(n_2308),
.B(n_343),
.C(n_346),
.Y(n_2326)
);

OAI22xp5_ASAP7_75t_L g2327 ( 
.A1(n_2326),
.A2(n_2317),
.B1(n_2314),
.B2(n_2307),
.Y(n_2327)
);

OAI22xp5_ASAP7_75t_SL g2328 ( 
.A1(n_2323),
.A2(n_2312),
.B1(n_347),
.B2(n_348),
.Y(n_2328)
);

OAI21xp5_ASAP7_75t_SL g2329 ( 
.A1(n_2325),
.A2(n_346),
.B(n_347),
.Y(n_2329)
);

OAI21xp5_ASAP7_75t_L g2330 ( 
.A1(n_2318),
.A2(n_348),
.B(n_349),
.Y(n_2330)
);

OAI22xp5_ASAP7_75t_SL g2331 ( 
.A1(n_2328),
.A2(n_2322),
.B1(n_2324),
.B2(n_2321),
.Y(n_2331)
);

AOI22x1_ASAP7_75t_L g2332 ( 
.A1(n_2330),
.A2(n_2319),
.B1(n_2320),
.B2(n_351),
.Y(n_2332)
);

HB1xp67_ASAP7_75t_L g2333 ( 
.A(n_2329),
.Y(n_2333)
);

OAI22xp5_ASAP7_75t_SL g2334 ( 
.A1(n_2327),
.A2(n_349),
.B1(n_350),
.B2(n_352),
.Y(n_2334)
);

AOI22xp33_ASAP7_75t_L g2335 ( 
.A1(n_2332),
.A2(n_350),
.B1(n_352),
.B2(n_353),
.Y(n_2335)
);

OAI22xp5_ASAP7_75t_L g2336 ( 
.A1(n_2334),
.A2(n_353),
.B1(n_354),
.B2(n_355),
.Y(n_2336)
);

OAI331xp33_ASAP7_75t_L g2337 ( 
.A1(n_2333),
.A2(n_354),
.A3(n_355),
.B1(n_356),
.B2(n_357),
.B3(n_358),
.C1(n_360),
.Y(n_2337)
);

OR3x1_ASAP7_75t_L g2338 ( 
.A(n_2335),
.B(n_2331),
.C(n_361),
.Y(n_2338)
);

AOI221x1_ASAP7_75t_L g2339 ( 
.A1(n_2336),
.A2(n_356),
.B1(n_362),
.B2(n_363),
.C(n_364),
.Y(n_2339)
);

INVx1_ASAP7_75t_L g2340 ( 
.A(n_2338),
.Y(n_2340)
);

XOR2xp5_ASAP7_75t_L g2341 ( 
.A(n_2339),
.B(n_2337),
.Y(n_2341)
);

AOI21xp5_ASAP7_75t_L g2342 ( 
.A1(n_2341),
.A2(n_362),
.B(n_364),
.Y(n_2342)
);

AOI22xp33_ASAP7_75t_L g2343 ( 
.A1(n_2342),
.A2(n_2340),
.B1(n_366),
.B2(n_367),
.Y(n_2343)
);

OR2x6_ASAP7_75t_L g2344 ( 
.A(n_2343),
.B(n_365),
.Y(n_2344)
);

AOI221xp5_ASAP7_75t_L g2345 ( 
.A1(n_2344),
.A2(n_366),
.B1(n_367),
.B2(n_368),
.C(n_369),
.Y(n_2345)
);

AOI211xp5_ASAP7_75t_L g2346 ( 
.A1(n_2345),
.A2(n_368),
.B(n_370),
.C(n_371),
.Y(n_2346)
);


endmodule