module fake_jpeg_21985_n_318 (n_13, n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_318);

input n_13;
input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_318;

wire n_253;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_15;
wire n_141;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_14;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_317;
wire n_20;
wire n_145;
wire n_18;
wire n_303;
wire n_259;
wire n_90;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_247;
wire n_157;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

CKINVDCx20_ASAP7_75t_R g14 ( 
.A(n_3),
.Y(n_14)
);

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_5),
.Y(n_15)
);

INVx4_ASAP7_75t_L g16 ( 
.A(n_1),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_4),
.Y(n_17)
);

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_11),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_9),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_4),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_9),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_9),
.Y(n_22)
);

BUFx6f_ASAP7_75t_SL g23 ( 
.A(n_13),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_7),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_0),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_4),
.Y(n_26)
);

CKINVDCx5p33_ASAP7_75t_R g27 ( 
.A(n_3),
.Y(n_27)
);

INVx4_ASAP7_75t_L g28 ( 
.A(n_10),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_14),
.Y(n_29)
);

NOR2xp33_ASAP7_75t_L g42 ( 
.A(n_29),
.B(n_31),
.Y(n_42)
);

INVx3_ASAP7_75t_L g30 ( 
.A(n_23),
.Y(n_30)
);

INVx8_ASAP7_75t_L g48 ( 
.A(n_30),
.Y(n_48)
);

INVx6_ASAP7_75t_L g31 ( 
.A(n_20),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_23),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_32),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_14),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_L g44 ( 
.A(n_33),
.B(n_29),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_23),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_34),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_23),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_35),
.Y(n_47)
);

INVx2_ASAP7_75t_L g36 ( 
.A(n_20),
.Y(n_36)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_36),
.Y(n_52)
);

BUFx12f_ASAP7_75t_L g37 ( 
.A(n_20),
.Y(n_37)
);

BUFx12f_ASAP7_75t_L g40 ( 
.A(n_37),
.Y(n_40)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_16),
.Y(n_38)
);

NAND2xp5_ASAP7_75t_SL g43 ( 
.A(n_38),
.B(n_27),
.Y(n_43)
);

OAI22xp5_ASAP7_75t_L g39 ( 
.A1(n_31),
.A2(n_28),
.B1(n_16),
.B2(n_25),
.Y(n_39)
);

OAI22xp5_ASAP7_75t_L g75 ( 
.A1(n_39),
.A2(n_31),
.B1(n_30),
.B2(n_36),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_43),
.B(n_44),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_L g45 ( 
.A(n_38),
.B(n_27),
.Y(n_45)
);

AND2x2_ASAP7_75t_L g73 ( 
.A(n_45),
.B(n_33),
.Y(n_73)
);

INVx2_ASAP7_75t_L g49 ( 
.A(n_37),
.Y(n_49)
);

INVx11_ASAP7_75t_L g65 ( 
.A(n_49),
.Y(n_65)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_37),
.Y(n_50)
);

INVx8_ASAP7_75t_L g67 ( 
.A(n_50),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_SL g51 ( 
.A(n_29),
.B(n_27),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_L g62 ( 
.A(n_51),
.B(n_56),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_37),
.Y(n_53)
);

INVx4_ASAP7_75t_L g69 ( 
.A(n_53),
.Y(n_69)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_37),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_54),
.B(n_55),
.Y(n_76)
);

INVx2_ASAP7_75t_L g55 ( 
.A(n_37),
.Y(n_55)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_37),
.Y(n_56)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_42),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_57),
.B(n_58),
.Y(n_83)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_42),
.Y(n_58)
);

INVx2_ASAP7_75t_L g59 ( 
.A(n_48),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_59),
.B(n_61),
.Y(n_88)
);

AOI22xp33_ASAP7_75t_L g60 ( 
.A1(n_48),
.A2(n_31),
.B1(n_16),
.B2(n_28),
.Y(n_60)
);

OAI22xp5_ASAP7_75t_L g99 ( 
.A1(n_60),
.A2(n_16),
.B1(n_28),
.B2(n_55),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_SL g61 ( 
.A(n_44),
.B(n_33),
.Y(n_61)
);

INVx2_ASAP7_75t_L g63 ( 
.A(n_48),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_63),
.B(n_64),
.Y(n_91)
);

INVx2_ASAP7_75t_SL g64 ( 
.A(n_40),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_L g66 ( 
.A(n_45),
.B(n_38),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_L g80 ( 
.A(n_66),
.B(n_73),
.Y(n_80)
);

INVx2_ASAP7_75t_L g68 ( 
.A(n_40),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_68),
.B(n_71),
.Y(n_98)
);

INVx2_ASAP7_75t_L g71 ( 
.A(n_40),
.Y(n_71)
);

INVx4_ASAP7_75t_L g72 ( 
.A(n_40),
.Y(n_72)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_72),
.Y(n_82)
);

INVx2_ASAP7_75t_L g74 ( 
.A(n_40),
.Y(n_74)
);

INVx2_ASAP7_75t_L g84 ( 
.A(n_74),
.Y(n_84)
);

AOI22xp5_ASAP7_75t_L g79 ( 
.A1(n_75),
.A2(n_30),
.B1(n_39),
.B2(n_36),
.Y(n_79)
);

CKINVDCx20_ASAP7_75t_R g77 ( 
.A(n_51),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_L g81 ( 
.A(n_77),
.B(n_43),
.Y(n_81)
);

OR2x2_ASAP7_75t_L g78 ( 
.A(n_70),
.B(n_40),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_L g101 ( 
.A(n_78),
.B(n_85),
.Y(n_101)
);

OAI22xp5_ASAP7_75t_L g111 ( 
.A1(n_79),
.A2(n_100),
.B1(n_59),
.B2(n_67),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_SL g113 ( 
.A(n_81),
.B(n_49),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_L g85 ( 
.A(n_66),
.B(n_56),
.Y(n_85)
);

OAI21xp5_ASAP7_75t_SL g86 ( 
.A1(n_62),
.A2(n_52),
.B(n_54),
.Y(n_86)
);

OAI22xp5_ASAP7_75t_SL g103 ( 
.A1(n_86),
.A2(n_58),
.B1(n_70),
.B2(n_73),
.Y(n_103)
);

OAI32xp33_ASAP7_75t_L g87 ( 
.A1(n_62),
.A2(n_30),
.A3(n_52),
.B1(n_35),
.B2(n_34),
.Y(n_87)
);

AOI22xp5_ASAP7_75t_L g108 ( 
.A1(n_87),
.A2(n_90),
.B1(n_99),
.B2(n_63),
.Y(n_108)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_76),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g121 ( 
.A(n_89),
.B(n_92),
.Y(n_121)
);

OAI22xp5_ASAP7_75t_SL g90 ( 
.A1(n_57),
.A2(n_16),
.B1(n_28),
.B2(n_55),
.Y(n_90)
);

INVx2_ASAP7_75t_L g92 ( 
.A(n_67),
.Y(n_92)
);

INVx2_ASAP7_75t_L g93 ( 
.A(n_67),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g122 ( 
.A(n_93),
.B(n_94),
.Y(n_122)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_76),
.Y(n_94)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_61),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g106 ( 
.A(n_95),
.B(n_96),
.Y(n_106)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_73),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g97 ( 
.A(n_73),
.B(n_53),
.Y(n_97)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_97),
.Y(n_104)
);

AOI22xp5_ASAP7_75t_L g100 ( 
.A1(n_75),
.A2(n_28),
.B1(n_35),
.B2(n_34),
.Y(n_100)
);

AND2x2_ASAP7_75t_SL g102 ( 
.A(n_97),
.B(n_77),
.Y(n_102)
);

OAI21xp5_ASAP7_75t_SL g133 ( 
.A1(n_102),
.A2(n_103),
.B(n_109),
.Y(n_133)
);

CKINVDCx20_ASAP7_75t_R g105 ( 
.A(n_98),
.Y(n_105)
);

CKINVDCx20_ASAP7_75t_R g127 ( 
.A(n_105),
.Y(n_127)
);

BUFx3_ASAP7_75t_L g107 ( 
.A(n_84),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_L g134 ( 
.A(n_107),
.B(n_110),
.Y(n_134)
);

OAI22xp5_ASAP7_75t_L g126 ( 
.A1(n_108),
.A2(n_116),
.B1(n_120),
.B2(n_100),
.Y(n_126)
);

AND2x2_ASAP7_75t_L g109 ( 
.A(n_80),
.B(n_34),
.Y(n_109)
);

INVx2_ASAP7_75t_L g110 ( 
.A(n_84),
.Y(n_110)
);

AOI22xp5_ASAP7_75t_L g140 ( 
.A1(n_111),
.A2(n_114),
.B1(n_99),
.B2(n_90),
.Y(n_140)
);

OAI22xp33_ASAP7_75t_SL g112 ( 
.A1(n_87),
.A2(n_65),
.B1(n_49),
.B2(n_69),
.Y(n_112)
);

AOI22xp33_ASAP7_75t_L g141 ( 
.A1(n_112),
.A2(n_118),
.B1(n_91),
.B2(n_94),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_L g129 ( 
.A(n_113),
.B(n_115),
.Y(n_129)
);

OAI22xp5_ASAP7_75t_L g114 ( 
.A1(n_79),
.A2(n_65),
.B1(n_69),
.B2(n_71),
.Y(n_114)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_91),
.Y(n_115)
);

AOI22xp33_ASAP7_75t_L g116 ( 
.A1(n_79),
.A2(n_65),
.B1(n_69),
.B2(n_72),
.Y(n_116)
);

AOI22xp5_ASAP7_75t_SL g117 ( 
.A1(n_96),
.A2(n_72),
.B1(n_64),
.B2(n_68),
.Y(n_117)
);

INVxp67_ASAP7_75t_L g136 ( 
.A(n_117),
.Y(n_136)
);

CKINVDCx16_ASAP7_75t_R g118 ( 
.A(n_98),
.Y(n_118)
);

BUFx6f_ASAP7_75t_L g119 ( 
.A(n_92),
.Y(n_119)
);

CKINVDCx16_ASAP7_75t_R g131 ( 
.A(n_119),
.Y(n_131)
);

AOI22xp5_ASAP7_75t_L g120 ( 
.A1(n_80),
.A2(n_35),
.B1(n_32),
.B2(n_64),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_SL g123 ( 
.A(n_95),
.B(n_24),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_L g143 ( 
.A(n_123),
.B(n_88),
.Y(n_143)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_121),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_L g167 ( 
.A(n_124),
.B(n_128),
.Y(n_167)
);

AO22x1_ASAP7_75t_L g125 ( 
.A1(n_112),
.A2(n_87),
.B1(n_108),
.B2(n_116),
.Y(n_125)
);

OAI21xp5_ASAP7_75t_L g160 ( 
.A1(n_125),
.A2(n_139),
.B(n_102),
.Y(n_160)
);

AOI22xp5_ASAP7_75t_L g168 ( 
.A1(n_126),
.A2(n_135),
.B1(n_144),
.B2(n_145),
.Y(n_168)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_121),
.Y(n_128)
);

INVxp33_ASAP7_75t_L g130 ( 
.A(n_107),
.Y(n_130)
);

CKINVDCx16_ASAP7_75t_R g153 ( 
.A(n_130),
.Y(n_153)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_122),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_L g150 ( 
.A(n_132),
.B(n_142),
.Y(n_150)
);

OAI22xp5_ASAP7_75t_L g135 ( 
.A1(n_104),
.A2(n_100),
.B1(n_86),
.B2(n_83),
.Y(n_135)
);

CKINVDCx16_ASAP7_75t_R g137 ( 
.A(n_122),
.Y(n_137)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_137),
.Y(n_155)
);

INVxp67_ASAP7_75t_L g138 ( 
.A(n_107),
.Y(n_138)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_138),
.Y(n_154)
);

AND2x4_ASAP7_75t_L g139 ( 
.A(n_109),
.B(n_78),
.Y(n_139)
);

OAI22xp5_ASAP7_75t_SL g152 ( 
.A1(n_140),
.A2(n_148),
.B1(n_120),
.B2(n_117),
.Y(n_152)
);

INVxp67_ASAP7_75t_L g157 ( 
.A(n_141),
.Y(n_157)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_113),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_L g162 ( 
.A(n_143),
.B(n_123),
.Y(n_162)
);

O2A1O1Ixp33_ASAP7_75t_L g144 ( 
.A1(n_101),
.A2(n_90),
.B(n_83),
.C(n_88),
.Y(n_144)
);

OAI22x1_ASAP7_75t_L g145 ( 
.A1(n_117),
.A2(n_78),
.B1(n_89),
.B2(n_93),
.Y(n_145)
);

XNOR2xp5_ASAP7_75t_L g146 ( 
.A(n_103),
.B(n_85),
.Y(n_146)
);

XNOR2xp5_ASAP7_75t_L g169 ( 
.A(n_146),
.B(n_27),
.Y(n_169)
);

CKINVDCx20_ASAP7_75t_R g147 ( 
.A(n_105),
.Y(n_147)
);

CKINVDCx20_ASAP7_75t_R g165 ( 
.A(n_147),
.Y(n_165)
);

AOI22xp33_ASAP7_75t_L g148 ( 
.A1(n_111),
.A2(n_114),
.B1(n_118),
.B2(n_109),
.Y(n_148)
);

XOR2xp5_ASAP7_75t_SL g149 ( 
.A(n_139),
.B(n_101),
.Y(n_149)
);

XNOR2xp5_ASAP7_75t_L g189 ( 
.A(n_149),
.B(n_169),
.Y(n_189)
);

BUFx8_ASAP7_75t_L g151 ( 
.A(n_145),
.Y(n_151)
);

NOR2xp33_ASAP7_75t_L g177 ( 
.A(n_151),
.B(n_147),
.Y(n_177)
);

AOI22xp5_ASAP7_75t_L g192 ( 
.A1(n_152),
.A2(n_156),
.B1(n_161),
.B2(n_32),
.Y(n_192)
);

OAI22xp5_ASAP7_75t_SL g156 ( 
.A1(n_125),
.A2(n_104),
.B1(n_106),
.B2(n_102),
.Y(n_156)
);

AOI21xp5_ASAP7_75t_L g158 ( 
.A1(n_133),
.A2(n_115),
.B(n_106),
.Y(n_158)
);

AOI21xp5_ASAP7_75t_L g180 ( 
.A1(n_158),
.A2(n_137),
.B(n_127),
.Y(n_180)
);

AND2x6_ASAP7_75t_L g159 ( 
.A(n_139),
.B(n_145),
.Y(n_159)
);

OAI21xp5_ASAP7_75t_L g176 ( 
.A1(n_159),
.A2(n_173),
.B(n_136),
.Y(n_176)
);

AO21x1_ASAP7_75t_L g201 ( 
.A1(n_160),
.A2(n_21),
.B(n_25),
.Y(n_201)
);

OAI22xp5_ASAP7_75t_SL g161 ( 
.A1(n_125),
.A2(n_102),
.B1(n_109),
.B2(n_81),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_L g197 ( 
.A(n_162),
.B(n_163),
.Y(n_197)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_129),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_L g164 ( 
.A(n_129),
.B(n_119),
.Y(n_164)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_164),
.Y(n_186)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_134),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_SL g178 ( 
.A(n_166),
.B(n_132),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_L g170 ( 
.A(n_142),
.B(n_119),
.Y(n_170)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_170),
.Y(n_193)
);

INVx4_ASAP7_75t_L g171 ( 
.A(n_131),
.Y(n_171)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_171),
.Y(n_190)
);

MAJIxp5_ASAP7_75t_L g172 ( 
.A(n_133),
.B(n_82),
.C(n_110),
.Y(n_172)
);

MAJIxp5_ASAP7_75t_L g198 ( 
.A(n_172),
.B(n_174),
.C(n_32),
.Y(n_198)
);

OAI21xp5_ASAP7_75t_L g173 ( 
.A1(n_139),
.A2(n_21),
.B(n_26),
.Y(n_173)
);

MAJIxp5_ASAP7_75t_L g174 ( 
.A(n_139),
.B(n_82),
.C(n_74),
.Y(n_174)
);

OAI21xp33_ASAP7_75t_L g175 ( 
.A1(n_143),
.A2(n_0),
.B(n_1),
.Y(n_175)
);

XNOR2xp5_ASAP7_75t_L g195 ( 
.A(n_175),
.B(n_173),
.Y(n_195)
);

OAI22xp5_ASAP7_75t_SL g210 ( 
.A1(n_176),
.A2(n_180),
.B1(n_187),
.B2(n_192),
.Y(n_210)
);

OR2x2_ASAP7_75t_L g213 ( 
.A(n_177),
.B(n_157),
.Y(n_213)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_178),
.Y(n_214)
);

NAND2xp5_ASAP7_75t_SL g179 ( 
.A(n_165),
.B(n_144),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_L g215 ( 
.A(n_179),
.B(n_181),
.Y(n_215)
);

NAND2xp5_ASAP7_75t_SL g181 ( 
.A(n_153),
.B(n_144),
.Y(n_181)
);

OAI22xp5_ASAP7_75t_SL g182 ( 
.A1(n_168),
.A2(n_140),
.B1(n_127),
.B2(n_126),
.Y(n_182)
);

AOI22xp5_ASAP7_75t_L g203 ( 
.A1(n_182),
.A2(n_183),
.B1(n_196),
.B2(n_152),
.Y(n_203)
);

OAI22xp5_ASAP7_75t_L g183 ( 
.A1(n_168),
.A2(n_124),
.B1(n_128),
.B2(n_135),
.Y(n_183)
);

NOR2xp33_ASAP7_75t_L g184 ( 
.A(n_171),
.B(n_131),
.Y(n_184)
);

CKINVDCx16_ASAP7_75t_R g209 ( 
.A(n_184),
.Y(n_209)
);

INVxp67_ASAP7_75t_L g185 ( 
.A(n_170),
.Y(n_185)
);

NOR2xp33_ASAP7_75t_L g206 ( 
.A(n_185),
.B(n_188),
.Y(n_206)
);

OAI22x1_ASAP7_75t_L g187 ( 
.A1(n_151),
.A2(n_149),
.B1(n_159),
.B2(n_157),
.Y(n_187)
);

NOR2xp33_ASAP7_75t_L g188 ( 
.A(n_156),
.B(n_146),
.Y(n_188)
);

CKINVDCx16_ASAP7_75t_R g191 ( 
.A(n_167),
.Y(n_191)
);

NOR2xp33_ASAP7_75t_L g207 ( 
.A(n_191),
.B(n_194),
.Y(n_207)
);

INVx2_ASAP7_75t_L g194 ( 
.A(n_154),
.Y(n_194)
);

XOR2xp5_ASAP7_75t_SL g223 ( 
.A(n_195),
.B(n_201),
.Y(n_223)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_164),
.Y(n_196)
);

MAJIxp5_ASAP7_75t_L g204 ( 
.A(n_198),
.B(n_174),
.C(n_193),
.Y(n_204)
);

NOR2xp33_ASAP7_75t_L g199 ( 
.A(n_163),
.B(n_64),
.Y(n_199)
);

CKINVDCx20_ASAP7_75t_R g211 ( 
.A(n_199),
.Y(n_211)
);

XNOR2xp5_ASAP7_75t_L g200 ( 
.A(n_160),
.B(n_172),
.Y(n_200)
);

XOR2xp5_ASAP7_75t_L g202 ( 
.A(n_200),
.B(n_158),
.Y(n_202)
);

XOR2xp5_ASAP7_75t_L g229 ( 
.A(n_202),
.B(n_205),
.Y(n_229)
);

OAI22xp5_ASAP7_75t_L g241 ( 
.A1(n_203),
.A2(n_14),
.B1(n_17),
.B2(n_19),
.Y(n_241)
);

MAJIxp5_ASAP7_75t_L g227 ( 
.A(n_204),
.B(n_208),
.C(n_212),
.Y(n_227)
);

XOR2xp5_ASAP7_75t_L g205 ( 
.A(n_200),
.B(n_161),
.Y(n_205)
);

MAJIxp5_ASAP7_75t_L g208 ( 
.A(n_198),
.B(n_150),
.C(n_155),
.Y(n_208)
);

MAJIxp5_ASAP7_75t_L g212 ( 
.A(n_193),
.B(n_150),
.C(n_155),
.Y(n_212)
);

CKINVDCx20_ASAP7_75t_R g230 ( 
.A(n_213),
.Y(n_230)
);

CKINVDCx20_ASAP7_75t_R g216 ( 
.A(n_197),
.Y(n_216)
);

NAND2xp5_ASAP7_75t_L g224 ( 
.A(n_216),
.B(n_185),
.Y(n_224)
);

INVxp33_ASAP7_75t_L g217 ( 
.A(n_197),
.Y(n_217)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_217),
.Y(n_225)
);

MAJIxp5_ASAP7_75t_L g218 ( 
.A(n_186),
.B(n_169),
.C(n_162),
.Y(n_218)
);

MAJIxp5_ASAP7_75t_L g231 ( 
.A(n_218),
.B(n_220),
.C(n_221),
.Y(n_231)
);

XOR2xp5_ASAP7_75t_L g219 ( 
.A(n_187),
.B(n_151),
.Y(n_219)
);

MAJIxp5_ASAP7_75t_L g236 ( 
.A(n_219),
.B(n_222),
.C(n_21),
.Y(n_236)
);

MAJIxp5_ASAP7_75t_L g220 ( 
.A(n_186),
.B(n_53),
.C(n_50),
.Y(n_220)
);

MAJIxp5_ASAP7_75t_L g221 ( 
.A(n_196),
.B(n_53),
.C(n_50),
.Y(n_221)
);

XNOR2xp5_ASAP7_75t_SL g222 ( 
.A(n_192),
.B(n_18),
.Y(n_222)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_224),
.Y(n_247)
);

AOI22xp5_ASAP7_75t_SL g226 ( 
.A1(n_214),
.A2(n_190),
.B1(n_194),
.B2(n_182),
.Y(n_226)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_226),
.Y(n_248)
);

AOI22xp5_ASAP7_75t_L g228 ( 
.A1(n_210),
.A2(n_180),
.B1(n_176),
.B2(n_201),
.Y(n_228)
);

OAI22xp5_ASAP7_75t_L g251 ( 
.A1(n_228),
.A2(n_223),
.B1(n_215),
.B2(n_222),
.Y(n_251)
);

XNOR2xp5_ASAP7_75t_L g232 ( 
.A(n_208),
.B(n_189),
.Y(n_232)
);

NOR2xp33_ASAP7_75t_L g262 ( 
.A(n_232),
.B(n_233),
.Y(n_262)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_207),
.Y(n_233)
);

MAJIxp5_ASAP7_75t_L g234 ( 
.A(n_204),
.B(n_189),
.C(n_195),
.Y(n_234)
);

NOR2xp33_ASAP7_75t_SL g257 ( 
.A(n_234),
.B(n_237),
.Y(n_257)
);

AND2x2_ASAP7_75t_L g235 ( 
.A(n_219),
.B(n_0),
.Y(n_235)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_235),
.Y(n_249)
);

CKINVDCx14_ASAP7_75t_R g246 ( 
.A(n_236),
.Y(n_246)
);

MAJIxp5_ASAP7_75t_L g237 ( 
.A(n_212),
.B(n_50),
.C(n_41),
.Y(n_237)
);

MAJIxp5_ASAP7_75t_L g238 ( 
.A(n_202),
.B(n_21),
.C(n_26),
.Y(n_238)
);

NAND2xp5_ASAP7_75t_L g258 ( 
.A(n_238),
.B(n_239),
.Y(n_258)
);

XNOR2xp5_ASAP7_75t_L g239 ( 
.A(n_205),
.B(n_206),
.Y(n_239)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_217),
.Y(n_240)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_240),
.Y(n_250)
);

AOI22xp5_ASAP7_75t_L g245 ( 
.A1(n_241),
.A2(n_242),
.B1(n_26),
.B2(n_25),
.Y(n_245)
);

MAJIxp5_ASAP7_75t_L g242 ( 
.A(n_218),
.B(n_25),
.C(n_26),
.Y(n_242)
);

NOR2xp33_ASAP7_75t_L g243 ( 
.A(n_211),
.B(n_0),
.Y(n_243)
);

AOI22xp5_ASAP7_75t_SL g259 ( 
.A1(n_243),
.A2(n_24),
.B1(n_19),
.B2(n_17),
.Y(n_259)
);

MAJIxp5_ASAP7_75t_L g244 ( 
.A(n_220),
.B(n_41),
.C(n_32),
.Y(n_244)
);

OAI21xp5_ASAP7_75t_SL g261 ( 
.A1(n_244),
.A2(n_20),
.B(n_46),
.Y(n_261)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_245),
.Y(n_269)
);

AOI22xp5_ASAP7_75t_L g266 ( 
.A1(n_251),
.A2(n_252),
.B1(n_253),
.B2(n_256),
.Y(n_266)
);

OAI22xp5_ASAP7_75t_SL g252 ( 
.A1(n_225),
.A2(n_230),
.B1(n_227),
.B2(n_231),
.Y(n_252)
);

OAI22xp5_ASAP7_75t_SL g253 ( 
.A1(n_227),
.A2(n_213),
.B1(n_221),
.B2(n_223),
.Y(n_253)
);

AOI22xp5_ASAP7_75t_L g254 ( 
.A1(n_231),
.A2(n_209),
.B1(n_14),
.B2(n_19),
.Y(n_254)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_254),
.Y(n_277)
);

AOI21xp5_ASAP7_75t_L g255 ( 
.A1(n_235),
.A2(n_24),
.B(n_19),
.Y(n_255)
);

OAI21xp5_ASAP7_75t_L g264 ( 
.A1(n_255),
.A2(n_15),
.B(n_244),
.Y(n_264)
);

OAI22xp5_ASAP7_75t_SL g256 ( 
.A1(n_234),
.A2(n_15),
.B1(n_17),
.B2(n_24),
.Y(n_256)
);

NAND2xp5_ASAP7_75t_L g267 ( 
.A(n_259),
.B(n_15),
.Y(n_267)
);

OAI322xp33_ASAP7_75t_L g260 ( 
.A1(n_229),
.A2(n_17),
.A3(n_15),
.B1(n_3),
.B2(n_4),
.C1(n_5),
.C2(n_6),
.Y(n_260)
);

AOI21xp5_ASAP7_75t_L g276 ( 
.A1(n_260),
.A2(n_261),
.B(n_5),
.Y(n_276)
);

MAJIxp5_ASAP7_75t_L g263 ( 
.A(n_257),
.B(n_237),
.C(n_229),
.Y(n_263)
);

MAJIxp5_ASAP7_75t_L g279 ( 
.A(n_263),
.B(n_273),
.C(n_275),
.Y(n_279)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_264),
.Y(n_285)
);

XOR2xp5_ASAP7_75t_L g265 ( 
.A(n_252),
.B(n_1),
.Y(n_265)
);

MAJIxp5_ASAP7_75t_L g288 ( 
.A(n_265),
.B(n_274),
.C(n_5),
.Y(n_288)
);

NAND2xp5_ASAP7_75t_L g286 ( 
.A(n_267),
.B(n_270),
.Y(n_286)
);

AOI22xp5_ASAP7_75t_SL g268 ( 
.A1(n_248),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_268)
);

OAI22xp5_ASAP7_75t_SL g280 ( 
.A1(n_268),
.A2(n_276),
.B1(n_259),
.B2(n_255),
.Y(n_280)
);

NAND2xp5_ASAP7_75t_SL g270 ( 
.A(n_262),
.B(n_2),
.Y(n_270)
);

NAND2xp5_ASAP7_75t_SL g271 ( 
.A(n_249),
.B(n_2),
.Y(n_271)
);

NOR2xp33_ASAP7_75t_L g284 ( 
.A(n_271),
.B(n_272),
.Y(n_284)
);

NAND2xp5_ASAP7_75t_SL g272 ( 
.A(n_249),
.B(n_2),
.Y(n_272)
);

MAJIxp5_ASAP7_75t_L g273 ( 
.A(n_250),
.B(n_41),
.C(n_46),
.Y(n_273)
);

XOR2xp5_ASAP7_75t_L g274 ( 
.A(n_253),
.B(n_258),
.Y(n_274)
);

MAJIxp5_ASAP7_75t_L g275 ( 
.A(n_250),
.B(n_41),
.C(n_46),
.Y(n_275)
);

AOI21xp33_ASAP7_75t_SL g278 ( 
.A1(n_274),
.A2(n_246),
.B(n_258),
.Y(n_278)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_278),
.Y(n_295)
);

NAND2xp5_ASAP7_75t_L g294 ( 
.A(n_280),
.B(n_22),
.Y(n_294)
);

OAI22xp5_ASAP7_75t_L g281 ( 
.A1(n_266),
.A2(n_247),
.B1(n_254),
.B2(n_261),
.Y(n_281)
);

AOI22xp5_ASAP7_75t_L g296 ( 
.A1(n_281),
.A2(n_22),
.B1(n_18),
.B2(n_20),
.Y(n_296)
);

BUFx2_ASAP7_75t_L g282 ( 
.A(n_273),
.Y(n_282)
);

NOR2xp33_ASAP7_75t_L g300 ( 
.A(n_282),
.B(n_6),
.Y(n_300)
);

AOI21xp5_ASAP7_75t_SL g283 ( 
.A1(n_277),
.A2(n_247),
.B(n_256),
.Y(n_283)
);

MAJx2_ASAP7_75t_L g292 ( 
.A(n_283),
.B(n_268),
.C(n_7),
.Y(n_292)
);

AOI22xp5_ASAP7_75t_L g287 ( 
.A1(n_263),
.A2(n_245),
.B1(n_22),
.B2(n_18),
.Y(n_287)
);

MAJIxp5_ASAP7_75t_L g293 ( 
.A(n_287),
.B(n_288),
.C(n_289),
.Y(n_293)
);

MAJIxp5_ASAP7_75t_L g289 ( 
.A(n_265),
.B(n_22),
.C(n_18),
.Y(n_289)
);

MAJIxp5_ASAP7_75t_L g290 ( 
.A(n_275),
.B(n_269),
.C(n_264),
.Y(n_290)
);

OAI21xp5_ASAP7_75t_L g299 ( 
.A1(n_290),
.A2(n_6),
.B(n_7),
.Y(n_299)
);

INVx2_ASAP7_75t_L g291 ( 
.A(n_282),
.Y(n_291)
);

NOR2xp33_ASAP7_75t_L g303 ( 
.A(n_291),
.B(n_279),
.Y(n_303)
);

AOI22xp33_ASAP7_75t_L g301 ( 
.A1(n_292),
.A2(n_300),
.B1(n_284),
.B2(n_285),
.Y(n_301)
);

NAND2xp5_ASAP7_75t_L g302 ( 
.A(n_294),
.B(n_296),
.Y(n_302)
);

AOI22xp5_ASAP7_75t_L g297 ( 
.A1(n_290),
.A2(n_22),
.B1(n_18),
.B2(n_20),
.Y(n_297)
);

MAJIxp5_ASAP7_75t_L g304 ( 
.A(n_297),
.B(n_299),
.C(n_300),
.Y(n_304)
);

AOI21x1_ASAP7_75t_L g298 ( 
.A1(n_283),
.A2(n_6),
.B(n_7),
.Y(n_298)
);

AOI322xp5_ASAP7_75t_L g306 ( 
.A1(n_298),
.A2(n_286),
.A3(n_9),
.B1(n_10),
.B2(n_11),
.C1(n_12),
.C2(n_8),
.Y(n_306)
);

NAND2xp5_ASAP7_75t_SL g309 ( 
.A(n_301),
.B(n_303),
.Y(n_309)
);

HB1xp67_ASAP7_75t_L g305 ( 
.A(n_292),
.Y(n_305)
);

MAJIxp5_ASAP7_75t_L g308 ( 
.A(n_305),
.B(n_307),
.C(n_8),
.Y(n_308)
);

NAND2xp5_ASAP7_75t_L g311 ( 
.A(n_306),
.B(n_8),
.Y(n_311)
);

AOI22xp5_ASAP7_75t_L g307 ( 
.A1(n_295),
.A2(n_293),
.B1(n_279),
.B2(n_47),
.Y(n_307)
);

AOI322xp5_ASAP7_75t_L g313 ( 
.A1(n_308),
.A2(n_310),
.A3(n_311),
.B1(n_302),
.B2(n_304),
.C1(n_47),
.C2(n_12),
.Y(n_313)
);

MAJIxp5_ASAP7_75t_L g310 ( 
.A(n_305),
.B(n_46),
.C(n_47),
.Y(n_310)
);

BUFx24_ASAP7_75t_SL g312 ( 
.A(n_309),
.Y(n_312)
);

NOR2xp67_ASAP7_75t_L g314 ( 
.A(n_312),
.B(n_313),
.Y(n_314)
);

AOI322xp5_ASAP7_75t_L g315 ( 
.A1(n_314),
.A2(n_47),
.A3(n_10),
.B1(n_11),
.B2(n_12),
.C1(n_13),
.C2(n_8),
.Y(n_315)
);

A2O1A1Ixp33_ASAP7_75t_SL g316 ( 
.A1(n_315),
.A2(n_10),
.B(n_11),
.C(n_12),
.Y(n_316)
);

BUFx24_ASAP7_75t_SL g317 ( 
.A(n_316),
.Y(n_317)
);

AOI21xp5_ASAP7_75t_L g318 ( 
.A1(n_317),
.A2(n_13),
.B(n_303),
.Y(n_318)
);


endmodule