module fake_jpeg_22950_n_131 (n_11, n_3, n_2, n_1, n_0, n_10, n_4, n_8, n_9, n_6, n_5, n_7, n_131);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_131;

wire n_117;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_31;
wire n_29;
wire n_103;
wire n_50;
wire n_15;
wire n_124;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_30;
wire n_106;
wire n_111;
wire n_24;
wire n_44;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_20;
wire n_18;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_56;
wire n_79;
wire n_12;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_22;
wire n_101;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_97;
wire n_36;
wire n_62;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_96;

CKINVDCx5p33_ASAP7_75t_R g12 ( 
.A(n_5),
.Y(n_12)
);

INVx6_ASAP7_75t_SL g13 ( 
.A(n_10),
.Y(n_13)
);

CKINVDCx20_ASAP7_75t_R g14 ( 
.A(n_8),
.Y(n_14)
);

INVx1_ASAP7_75t_L g15 ( 
.A(n_5),
.Y(n_15)
);

BUFx6f_ASAP7_75t_L g16 ( 
.A(n_7),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_9),
.Y(n_17)
);

BUFx3_ASAP7_75t_L g18 ( 
.A(n_11),
.Y(n_18)
);

INVx4_ASAP7_75t_L g19 ( 
.A(n_3),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_3),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_9),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_11),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_7),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_1),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_2),
.Y(n_25)
);

BUFx12f_ASAP7_75t_L g26 ( 
.A(n_2),
.Y(n_26)
);

NOR2xp33_ASAP7_75t_L g27 ( 
.A(n_14),
.B(n_0),
.Y(n_27)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_27),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g28 ( 
.A(n_20),
.B(n_0),
.Y(n_28)
);

NAND2xp5_ASAP7_75t_L g40 ( 
.A(n_28),
.B(n_31),
.Y(n_40)
);

BUFx3_ASAP7_75t_L g29 ( 
.A(n_26),
.Y(n_29)
);

CKINVDCx16_ASAP7_75t_R g43 ( 
.A(n_29),
.Y(n_43)
);

BUFx12f_ASAP7_75t_L g30 ( 
.A(n_26),
.Y(n_30)
);

CKINVDCx5p33_ASAP7_75t_R g36 ( 
.A(n_30),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g31 ( 
.A(n_20),
.B(n_21),
.Y(n_31)
);

BUFx4f_ASAP7_75t_SL g32 ( 
.A(n_26),
.Y(n_32)
);

INVx2_ASAP7_75t_L g38 ( 
.A(n_32),
.Y(n_38)
);

INVx6_ASAP7_75t_L g33 ( 
.A(n_16),
.Y(n_33)
);

AOI22xp33_ASAP7_75t_SL g46 ( 
.A1(n_33),
.A2(n_19),
.B1(n_16),
.B2(n_22),
.Y(n_46)
);

BUFx3_ASAP7_75t_L g34 ( 
.A(n_26),
.Y(n_34)
);

INVx2_ASAP7_75t_L g41 ( 
.A(n_34),
.Y(n_41)
);

BUFx12f_ASAP7_75t_L g35 ( 
.A(n_18),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_35),
.Y(n_39)
);

AND2x2_ASAP7_75t_L g37 ( 
.A(n_32),
.B(n_18),
.Y(n_37)
);

BUFx24_ASAP7_75t_SL g54 ( 
.A(n_37),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_L g42 ( 
.A(n_33),
.B(n_15),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_42),
.B(n_17),
.Y(n_50)
);

AND2x2_ASAP7_75t_L g45 ( 
.A(n_32),
.B(n_25),
.Y(n_45)
);

NAND2xp5_ASAP7_75t_L g47 ( 
.A(n_45),
.B(n_12),
.Y(n_47)
);

OAI22xp5_ASAP7_75t_L g48 ( 
.A1(n_46),
.A2(n_19),
.B1(n_35),
.B2(n_22),
.Y(n_48)
);

CKINVDCx14_ASAP7_75t_R g69 ( 
.A(n_47),
.Y(n_69)
);

AOI22xp5_ASAP7_75t_L g75 ( 
.A1(n_48),
.A2(n_56),
.B1(n_13),
.B2(n_24),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_L g49 ( 
.A(n_45),
.B(n_15),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_L g74 ( 
.A(n_49),
.B(n_53),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_50),
.B(n_52),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g51 ( 
.A(n_41),
.B(n_12),
.Y(n_51)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_51),
.Y(n_82)
);

INVx2_ASAP7_75t_L g52 ( 
.A(n_41),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_L g53 ( 
.A(n_36),
.B(n_17),
.Y(n_53)
);

CKINVDCx20_ASAP7_75t_R g55 ( 
.A(n_37),
.Y(n_55)
);

CKINVDCx20_ASAP7_75t_R g70 ( 
.A(n_55),
.Y(n_70)
);

OAI22xp5_ASAP7_75t_SL g56 ( 
.A1(n_46),
.A2(n_35),
.B1(n_30),
.B2(n_34),
.Y(n_56)
);

INVxp67_ASAP7_75t_L g57 ( 
.A(n_36),
.Y(n_57)
);

CKINVDCx16_ASAP7_75t_R g83 ( 
.A(n_57),
.Y(n_83)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_40),
.Y(n_58)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_58),
.Y(n_68)
);

INVx5_ASAP7_75t_L g59 ( 
.A(n_39),
.Y(n_59)
);

INVxp67_ASAP7_75t_L g77 ( 
.A(n_59),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_44),
.B(n_25),
.Y(n_60)
);

CKINVDCx20_ASAP7_75t_R g71 ( 
.A(n_60),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_L g61 ( 
.A(n_39),
.B(n_30),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_L g76 ( 
.A(n_61),
.B(n_63),
.Y(n_76)
);

INVx5_ASAP7_75t_L g62 ( 
.A(n_43),
.Y(n_62)
);

CKINVDCx12_ASAP7_75t_R g80 ( 
.A(n_62),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_38),
.B(n_23),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_38),
.B(n_23),
.Y(n_64)
);

XNOR2xp5_ASAP7_75t_L g81 ( 
.A(n_64),
.B(n_66),
.Y(n_81)
);

INVxp67_ASAP7_75t_L g65 ( 
.A(n_46),
.Y(n_65)
);

OAI21xp5_ASAP7_75t_L g78 ( 
.A1(n_65),
.A2(n_67),
.B(n_24),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_L g66 ( 
.A(n_42),
.B(n_30),
.Y(n_66)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_42),
.Y(n_67)
);

OAI22xp5_ASAP7_75t_SL g73 ( 
.A1(n_65),
.A2(n_35),
.B1(n_29),
.B2(n_21),
.Y(n_73)
);

OAI22xp5_ASAP7_75t_SL g84 ( 
.A1(n_73),
.A2(n_75),
.B1(n_79),
.B2(n_47),
.Y(n_84)
);

OAI21xp5_ASAP7_75t_L g92 ( 
.A1(n_78),
.A2(n_53),
.B(n_49),
.Y(n_92)
);

AOI22xp5_ASAP7_75t_L g79 ( 
.A1(n_56),
.A2(n_13),
.B1(n_1),
.B2(n_0),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_84),
.B(n_88),
.Y(n_98)
);

BUFx6f_ASAP7_75t_L g85 ( 
.A(n_80),
.Y(n_85)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_85),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_SL g86 ( 
.A(n_70),
.B(n_54),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_86),
.B(n_90),
.Y(n_99)
);

XNOR2x1_ASAP7_75t_SL g87 ( 
.A(n_81),
.B(n_66),
.Y(n_87)
);

XOR2xp5_ASAP7_75t_L g106 ( 
.A(n_87),
.B(n_75),
.Y(n_106)
);

INVx1_ASAP7_75t_SL g88 ( 
.A(n_77),
.Y(n_88)
);

INVx2_ASAP7_75t_L g89 ( 
.A(n_77),
.Y(n_89)
);

CKINVDCx20_ASAP7_75t_R g104 ( 
.A(n_89),
.Y(n_104)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_72),
.Y(n_90)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_76),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_L g103 ( 
.A(n_91),
.B(n_95),
.Y(n_103)
);

AOI21xp5_ASAP7_75t_L g105 ( 
.A1(n_92),
.A2(n_94),
.B(n_82),
.Y(n_105)
);

MAJIxp5_ASAP7_75t_L g93 ( 
.A(n_74),
.B(n_61),
.C(n_57),
.Y(n_93)
);

MAJIxp5_ASAP7_75t_L g100 ( 
.A(n_93),
.B(n_87),
.C(n_92),
.Y(n_100)
);

AND2x2_ASAP7_75t_L g94 ( 
.A(n_74),
.B(n_69),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_L g95 ( 
.A(n_76),
.B(n_62),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g96 ( 
.A(n_81),
.B(n_1),
.Y(n_96)
);

XNOR2xp5_ASAP7_75t_L g97 ( 
.A(n_96),
.B(n_78),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g111 ( 
.A(n_97),
.B(n_100),
.Y(n_111)
);

MAJIxp5_ASAP7_75t_L g102 ( 
.A(n_93),
.B(n_68),
.C(n_83),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_L g113 ( 
.A(n_102),
.B(n_106),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_105),
.B(n_84),
.Y(n_107)
);

AOI22xp5_ASAP7_75t_SL g114 ( 
.A1(n_107),
.A2(n_110),
.B1(n_104),
.B2(n_94),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_SL g108 ( 
.A(n_99),
.B(n_68),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_L g117 ( 
.A(n_108),
.B(n_109),
.Y(n_117)
);

CKINVDCx16_ASAP7_75t_R g109 ( 
.A(n_103),
.Y(n_109)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_98),
.Y(n_110)
);

AOI21xp5_ASAP7_75t_L g112 ( 
.A1(n_100),
.A2(n_89),
.B(n_52),
.Y(n_112)
);

AOI22xp33_ASAP7_75t_L g118 ( 
.A1(n_112),
.A2(n_88),
.B1(n_97),
.B2(n_59),
.Y(n_118)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_114),
.Y(n_120)
);

XOR2xp5_ASAP7_75t_L g115 ( 
.A(n_113),
.B(n_106),
.Y(n_115)
);

XOR2xp5_ASAP7_75t_L g122 ( 
.A(n_115),
.B(n_111),
.Y(n_122)
);

AOI22xp5_ASAP7_75t_L g116 ( 
.A1(n_113),
.A2(n_102),
.B1(n_73),
.B2(n_101),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_L g121 ( 
.A(n_116),
.B(n_119),
.Y(n_121)
);

MAJIxp5_ASAP7_75t_L g123 ( 
.A(n_118),
.B(n_79),
.C(n_85),
.Y(n_123)
);

CKINVDCx16_ASAP7_75t_R g119 ( 
.A(n_112),
.Y(n_119)
);

MAJIxp5_ASAP7_75t_L g124 ( 
.A(n_122),
.B(n_123),
.C(n_115),
.Y(n_124)
);

XOR2xp5_ASAP7_75t_L g129 ( 
.A(n_124),
.B(n_125),
.Y(n_129)
);

MAJIxp5_ASAP7_75t_L g125 ( 
.A(n_122),
.B(n_120),
.C(n_121),
.Y(n_125)
);

OAI31xp33_ASAP7_75t_L g126 ( 
.A1(n_120),
.A2(n_117),
.A3(n_118),
.B(n_71),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_L g128 ( 
.A(n_126),
.B(n_127),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_SL g127 ( 
.A(n_120),
.B(n_4),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_L g130 ( 
.A(n_128),
.B(n_129),
.Y(n_130)
);

AOI21xp5_ASAP7_75t_L g131 ( 
.A1(n_130),
.A2(n_4),
.B(n_6),
.Y(n_131)
);


endmodule