module fake_jpeg_20875_n_334 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_334);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_334;

wire n_253;
wire n_330;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_15;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

BUFx6f_ASAP7_75t_L g15 ( 
.A(n_11),
.Y(n_15)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_12),
.Y(n_16)
);

BUFx6f_ASAP7_75t_L g17 ( 
.A(n_11),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_13),
.Y(n_18)
);

INVxp67_ASAP7_75t_L g19 ( 
.A(n_13),
.Y(n_19)
);

BUFx5_ASAP7_75t_L g20 ( 
.A(n_5),
.Y(n_20)
);

BUFx3_ASAP7_75t_L g21 ( 
.A(n_2),
.Y(n_21)
);

INVx8_ASAP7_75t_L g22 ( 
.A(n_7),
.Y(n_22)
);

BUFx12f_ASAP7_75t_L g23 ( 
.A(n_12),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_10),
.Y(n_24)
);

INVx11_ASAP7_75t_L g25 ( 
.A(n_1),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_8),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_12),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_12),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_8),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_3),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_8),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_13),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_14),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_2),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_23),
.Y(n_35)
);

INVx6_ASAP7_75t_L g52 ( 
.A(n_35),
.Y(n_52)
);

CKINVDCx16_ASAP7_75t_R g36 ( 
.A(n_21),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g45 ( 
.A(n_36),
.B(n_37),
.Y(n_45)
);

INVx2_ASAP7_75t_L g37 ( 
.A(n_23),
.Y(n_37)
);

INVx2_ASAP7_75t_L g38 ( 
.A(n_23),
.Y(n_38)
);

INVx6_ASAP7_75t_L g53 ( 
.A(n_38),
.Y(n_53)
);

BUFx12f_ASAP7_75t_L g39 ( 
.A(n_23),
.Y(n_39)
);

INVx2_ASAP7_75t_SL g48 ( 
.A(n_39),
.Y(n_48)
);

INVx4_ASAP7_75t_L g40 ( 
.A(n_23),
.Y(n_40)
);

INVx3_ASAP7_75t_L g51 ( 
.A(n_40),
.Y(n_51)
);

BUFx3_ASAP7_75t_L g41 ( 
.A(n_21),
.Y(n_41)
);

INVx2_ASAP7_75t_L g47 ( 
.A(n_41),
.Y(n_47)
);

INVx3_ASAP7_75t_L g42 ( 
.A(n_22),
.Y(n_42)
);

INVx2_ASAP7_75t_L g50 ( 
.A(n_42),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_15),
.Y(n_43)
);

INVx6_ASAP7_75t_L g54 ( 
.A(n_43),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_15),
.Y(n_44)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_44),
.Y(n_58)
);

OAI22xp5_ASAP7_75t_L g46 ( 
.A1(n_38),
.A2(n_22),
.B1(n_25),
.B2(n_19),
.Y(n_46)
);

AOI22xp5_ASAP7_75t_L g63 ( 
.A1(n_46),
.A2(n_40),
.B1(n_36),
.B2(n_22),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_L g49 ( 
.A(n_39),
.B(n_29),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_L g80 ( 
.A(n_49),
.B(n_57),
.Y(n_80)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_40),
.Y(n_55)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_55),
.Y(n_69)
);

HB1xp67_ASAP7_75t_L g56 ( 
.A(n_38),
.Y(n_56)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_56),
.Y(n_71)
);

MAJIxp5_ASAP7_75t_L g57 ( 
.A(n_39),
.B(n_17),
.C(n_33),
.Y(n_57)
);

INVx2_ASAP7_75t_L g59 ( 
.A(n_35),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g93 ( 
.A(n_59),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_49),
.B(n_37),
.Y(n_60)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_60),
.Y(n_105)
);

INVx8_ASAP7_75t_L g61 ( 
.A(n_52),
.Y(n_61)
);

INVx3_ASAP7_75t_L g118 ( 
.A(n_61),
.Y(n_118)
);

INVx8_ASAP7_75t_L g62 ( 
.A(n_52),
.Y(n_62)
);

AOI22xp33_ASAP7_75t_SL g132 ( 
.A1(n_62),
.A2(n_82),
.B1(n_99),
.B2(n_101),
.Y(n_132)
);

OAI22xp5_ASAP7_75t_L g119 ( 
.A1(n_63),
.A2(n_65),
.B1(n_66),
.B2(n_83),
.Y(n_119)
);

INVxp67_ASAP7_75t_L g64 ( 
.A(n_45),
.Y(n_64)
);

INVxp67_ASAP7_75t_L g109 ( 
.A(n_64),
.Y(n_109)
);

AOI22xp5_ASAP7_75t_L g65 ( 
.A1(n_46),
.A2(n_42),
.B1(n_43),
.B2(n_44),
.Y(n_65)
);

OAI22xp5_ASAP7_75t_SL g124 ( 
.A1(n_65),
.A2(n_66),
.B1(n_74),
.B2(n_34),
.Y(n_124)
);

AOI22xp5_ASAP7_75t_L g66 ( 
.A1(n_58),
.A2(n_42),
.B1(n_43),
.B2(n_44),
.Y(n_66)
);

INVx2_ASAP7_75t_L g67 ( 
.A(n_51),
.Y(n_67)
);

BUFx12f_ASAP7_75t_L g128 ( 
.A(n_67),
.Y(n_128)
);

INVx5_ASAP7_75t_L g68 ( 
.A(n_51),
.Y(n_68)
);

BUFx6f_ASAP7_75t_L g121 ( 
.A(n_68),
.Y(n_121)
);

CKINVDCx20_ASAP7_75t_R g70 ( 
.A(n_56),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_70),
.B(n_73),
.Y(n_102)
);

INVx2_ASAP7_75t_L g72 ( 
.A(n_51),
.Y(n_72)
);

BUFx6f_ASAP7_75t_L g127 ( 
.A(n_72),
.Y(n_127)
);

INVx5_ASAP7_75t_SL g73 ( 
.A(n_48),
.Y(n_73)
);

OAI22xp5_ASAP7_75t_SL g74 ( 
.A1(n_57),
.A2(n_44),
.B1(n_43),
.B2(n_29),
.Y(n_74)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_45),
.Y(n_75)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_75),
.Y(n_131)
);

CKINVDCx16_ASAP7_75t_R g76 ( 
.A(n_55),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g116 ( 
.A(n_76),
.B(n_85),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_47),
.B(n_18),
.Y(n_77)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_77),
.Y(n_113)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_53),
.Y(n_78)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_78),
.Y(n_122)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_53),
.Y(n_79)
);

CKINVDCx20_ASAP7_75t_R g130 ( 
.A(n_79),
.Y(n_130)
);

INVx6_ASAP7_75t_L g81 ( 
.A(n_59),
.Y(n_81)
);

INVx4_ASAP7_75t_L g120 ( 
.A(n_81),
.Y(n_120)
);

INVx6_ASAP7_75t_L g82 ( 
.A(n_50),
.Y(n_82)
);

OR2x2_ASAP7_75t_SL g83 ( 
.A(n_48),
.B(n_20),
.Y(n_83)
);

FAx1_ASAP7_75t_SL g110 ( 
.A(n_83),
.B(n_95),
.CI(n_96),
.CON(n_110),
.SN(n_110)
);

NAND2xp5_ASAP7_75t_L g84 ( 
.A(n_53),
.B(n_39),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g107 ( 
.A(n_84),
.B(n_92),
.Y(n_107)
);

CKINVDCx14_ASAP7_75t_R g85 ( 
.A(n_47),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_50),
.B(n_18),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g133 ( 
.A(n_86),
.B(n_88),
.Y(n_133)
);

BUFx3_ASAP7_75t_L g87 ( 
.A(n_48),
.Y(n_87)
);

INVx2_ASAP7_75t_L g103 ( 
.A(n_87),
.Y(n_103)
);

INVx2_ASAP7_75t_L g88 ( 
.A(n_52),
.Y(n_88)
);

CKINVDCx20_ASAP7_75t_R g89 ( 
.A(n_58),
.Y(n_89)
);

AOI22xp5_ASAP7_75t_SL g112 ( 
.A1(n_89),
.A2(n_97),
.B1(n_82),
.B2(n_73),
.Y(n_112)
);

INVx2_ASAP7_75t_L g90 ( 
.A(n_54),
.Y(n_90)
);

INVx2_ASAP7_75t_L g106 ( 
.A(n_90),
.Y(n_106)
);

INVxp67_ASAP7_75t_L g91 ( 
.A(n_54),
.Y(n_91)
);

INVxp67_ASAP7_75t_L g115 ( 
.A(n_91),
.Y(n_115)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_54),
.Y(n_92)
);

BUFx2_ASAP7_75t_SL g94 ( 
.A(n_48),
.Y(n_94)
);

INVxp67_ASAP7_75t_L g125 ( 
.A(n_94),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_49),
.B(n_27),
.Y(n_95)
);

NAND2xp67_ASAP7_75t_SL g96 ( 
.A(n_49),
.B(n_20),
.Y(n_96)
);

CKINVDCx20_ASAP7_75t_R g97 ( 
.A(n_56),
.Y(n_97)
);

INVx2_ASAP7_75t_SL g98 ( 
.A(n_51),
.Y(n_98)
);

OA22x2_ASAP7_75t_L g129 ( 
.A1(n_98),
.A2(n_33),
.B1(n_32),
.B2(n_31),
.Y(n_129)
);

HB1xp67_ASAP7_75t_L g99 ( 
.A(n_56),
.Y(n_99)
);

AOI32xp33_ASAP7_75t_L g100 ( 
.A1(n_45),
.A2(n_25),
.A3(n_39),
.B1(n_41),
.B2(n_16),
.Y(n_100)
);

XNOR2xp5_ASAP7_75t_L g126 ( 
.A(n_100),
.B(n_21),
.Y(n_126)
);

INVx5_ASAP7_75t_L g101 ( 
.A(n_51),
.Y(n_101)
);

MAJIxp5_ASAP7_75t_L g104 ( 
.A(n_80),
.B(n_39),
.C(n_35),
.Y(n_104)
);

MAJIxp5_ASAP7_75t_L g145 ( 
.A(n_104),
.B(n_79),
.C(n_78),
.Y(n_145)
);

AO22x2_ASAP7_75t_L g108 ( 
.A1(n_96),
.A2(n_35),
.B1(n_41),
.B2(n_34),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_L g134 ( 
.A(n_108),
.B(n_117),
.Y(n_134)
);

AOI22xp33_ASAP7_75t_L g111 ( 
.A1(n_75),
.A2(n_25),
.B1(n_28),
.B2(n_24),
.Y(n_111)
);

AOI22xp5_ASAP7_75t_L g138 ( 
.A1(n_111),
.A2(n_119),
.B1(n_124),
.B2(n_126),
.Y(n_138)
);

OAI21xp5_ASAP7_75t_L g143 ( 
.A1(n_112),
.A2(n_71),
.B(n_91),
.Y(n_143)
);

AO21x2_ASAP7_75t_SL g114 ( 
.A1(n_80),
.A2(n_34),
.B(n_33),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_SL g158 ( 
.A(n_114),
.B(n_93),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_L g117 ( 
.A(n_64),
.B(n_27),
.Y(n_117)
);

O2A1O1Ixp33_ASAP7_75t_L g123 ( 
.A1(n_74),
.A2(n_16),
.B(n_24),
.C(n_28),
.Y(n_123)
);

OAI21xp5_ASAP7_75t_SL g152 ( 
.A1(n_123),
.A2(n_129),
.B(n_117),
.Y(n_152)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_122),
.Y(n_135)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_135),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_L g136 ( 
.A(n_107),
.B(n_84),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_L g162 ( 
.A(n_136),
.B(n_144),
.Y(n_162)
);

XOR2xp5_ASAP7_75t_L g137 ( 
.A(n_104),
.B(n_63),
.Y(n_137)
);

XNOR2xp5_ASAP7_75t_L g184 ( 
.A(n_137),
.B(n_140),
.Y(n_184)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_107),
.Y(n_139)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_139),
.Y(n_189)
);

XOR2xp5_ASAP7_75t_L g140 ( 
.A(n_126),
.B(n_70),
.Y(n_140)
);

OAI22xp5_ASAP7_75t_SL g141 ( 
.A1(n_114),
.A2(n_124),
.B1(n_131),
.B2(n_105),
.Y(n_141)
);

AOI22xp5_ASAP7_75t_L g164 ( 
.A1(n_141),
.A2(n_158),
.B1(n_123),
.B2(n_108),
.Y(n_164)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_102),
.Y(n_142)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_142),
.Y(n_166)
);

AOI22xp5_ASAP7_75t_SL g191 ( 
.A1(n_143),
.A2(n_32),
.B1(n_31),
.B2(n_30),
.Y(n_191)
);

NOR2xp33_ASAP7_75t_L g144 ( 
.A(n_131),
.B(n_69),
.Y(n_144)
);

XOR2xp5_ASAP7_75t_L g163 ( 
.A(n_145),
.B(n_133),
.Y(n_163)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_127),
.Y(n_146)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_146),
.Y(n_171)
);

INVx3_ASAP7_75t_L g147 ( 
.A(n_128),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_L g173 ( 
.A(n_147),
.B(n_153),
.Y(n_173)
);

AOI22xp5_ASAP7_75t_SL g148 ( 
.A1(n_108),
.A2(n_69),
.B1(n_71),
.B2(n_92),
.Y(n_148)
);

OAI21xp5_ASAP7_75t_SL g167 ( 
.A1(n_148),
.A2(n_152),
.B(n_155),
.Y(n_167)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_127),
.Y(n_149)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_149),
.Y(n_172)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_112),
.Y(n_150)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_150),
.Y(n_181)
);

OR2x2_ASAP7_75t_L g151 ( 
.A(n_110),
.B(n_67),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_L g169 ( 
.A(n_151),
.B(n_154),
.Y(n_169)
);

NOR2xp33_ASAP7_75t_SL g153 ( 
.A(n_110),
.B(n_72),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_L g154 ( 
.A(n_109),
.B(n_93),
.Y(n_154)
);

OAI21xp33_ASAP7_75t_SL g155 ( 
.A1(n_108),
.A2(n_114),
.B(n_110),
.Y(n_155)
);

AOI22xp5_ASAP7_75t_L g156 ( 
.A1(n_114),
.A2(n_90),
.B1(n_81),
.B2(n_88),
.Y(n_156)
);

OAI22xp5_ASAP7_75t_SL g194 ( 
.A1(n_156),
.A2(n_30),
.B1(n_26),
.B2(n_17),
.Y(n_194)
);

AOI21xp5_ASAP7_75t_L g157 ( 
.A1(n_109),
.A2(n_14),
.B(n_1),
.Y(n_157)
);

OAI21xp5_ASAP7_75t_SL g168 ( 
.A1(n_157),
.A2(n_129),
.B(n_115),
.Y(n_168)
);

HB1xp67_ASAP7_75t_L g159 ( 
.A(n_128),
.Y(n_159)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_159),
.Y(n_183)
);

CKINVDCx20_ASAP7_75t_R g160 ( 
.A(n_128),
.Y(n_160)
);

NOR2xp33_ASAP7_75t_L g186 ( 
.A(n_160),
.B(n_87),
.Y(n_186)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_116),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_L g175 ( 
.A(n_161),
.B(n_125),
.Y(n_175)
);

MAJIxp5_ASAP7_75t_L g198 ( 
.A(n_163),
.B(n_153),
.C(n_151),
.Y(n_198)
);

OAI22xp5_ASAP7_75t_SL g219 ( 
.A1(n_164),
.A2(n_170),
.B1(n_174),
.B2(n_178),
.Y(n_219)
);

AOI22xp33_ASAP7_75t_SL g165 ( 
.A1(n_150),
.A2(n_118),
.B1(n_103),
.B2(n_113),
.Y(n_165)
);

OAI22xp5_ASAP7_75t_L g197 ( 
.A1(n_165),
.A2(n_176),
.B1(n_147),
.B2(n_146),
.Y(n_197)
);

OAI21xp5_ASAP7_75t_SL g207 ( 
.A1(n_168),
.A2(n_180),
.B(n_136),
.Y(n_207)
);

AOI22xp5_ASAP7_75t_L g170 ( 
.A1(n_141),
.A2(n_130),
.B1(n_129),
.B2(n_120),
.Y(n_170)
);

AOI22xp5_ASAP7_75t_L g174 ( 
.A1(n_158),
.A2(n_129),
.B1(n_120),
.B2(n_115),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_SL g199 ( 
.A(n_175),
.B(n_144),
.Y(n_199)
);

AOI22xp33_ASAP7_75t_SL g176 ( 
.A1(n_142),
.A2(n_118),
.B1(n_103),
.B2(n_101),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_L g177 ( 
.A(n_139),
.B(n_125),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_L g200 ( 
.A(n_177),
.B(n_154),
.Y(n_200)
);

AOI22xp5_ASAP7_75t_L g178 ( 
.A1(n_155),
.A2(n_62),
.B1(n_61),
.B2(n_106),
.Y(n_178)
);

AOI22xp5_ASAP7_75t_L g179 ( 
.A1(n_134),
.A2(n_106),
.B1(n_132),
.B2(n_98),
.Y(n_179)
);

OAI22xp5_ASAP7_75t_SL g222 ( 
.A1(n_179),
.A2(n_185),
.B1(n_187),
.B2(n_193),
.Y(n_222)
);

OAI21xp5_ASAP7_75t_SL g180 ( 
.A1(n_134),
.A2(n_121),
.B(n_98),
.Y(n_180)
);

OAI22xp5_ASAP7_75t_L g182 ( 
.A1(n_138),
.A2(n_68),
.B1(n_30),
.B2(n_32),
.Y(n_182)
);

AOI22xp5_ASAP7_75t_L g203 ( 
.A1(n_182),
.A2(n_194),
.B1(n_149),
.B2(n_135),
.Y(n_203)
);

AOI22xp5_ASAP7_75t_L g185 ( 
.A1(n_138),
.A2(n_121),
.B1(n_0),
.B2(n_2),
.Y(n_185)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_186),
.Y(n_195)
);

AOI22xp5_ASAP7_75t_L g187 ( 
.A1(n_152),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_187)
);

XNOR2xp5_ASAP7_75t_L g190 ( 
.A(n_140),
.B(n_31),
.Y(n_190)
);

XNOR2xp5_ASAP7_75t_L g214 ( 
.A(n_190),
.B(n_192),
.Y(n_214)
);

OAI21xp5_ASAP7_75t_L g206 ( 
.A1(n_191),
.A2(n_157),
.B(n_159),
.Y(n_206)
);

XNOR2xp5_ASAP7_75t_L g192 ( 
.A(n_145),
.B(n_26),
.Y(n_192)
);

AOI22xp5_ASAP7_75t_L g193 ( 
.A1(n_156),
.A2(n_0),
.B1(n_1),
.B2(n_3),
.Y(n_193)
);

AOI21xp5_ASAP7_75t_L g196 ( 
.A1(n_167),
.A2(n_143),
.B(n_151),
.Y(n_196)
);

OAI21xp5_ASAP7_75t_SL g239 ( 
.A1(n_196),
.A2(n_197),
.B(n_201),
.Y(n_239)
);

MAJIxp5_ASAP7_75t_L g232 ( 
.A(n_198),
.B(n_205),
.C(n_211),
.Y(n_232)
);

NAND2xp5_ASAP7_75t_SL g230 ( 
.A(n_199),
.B(n_216),
.Y(n_230)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_200),
.Y(n_229)
);

AOI21xp5_ASAP7_75t_L g201 ( 
.A1(n_167),
.A2(n_148),
.B(n_160),
.Y(n_201)
);

INVx2_ASAP7_75t_L g202 ( 
.A(n_183),
.Y(n_202)
);

NOR2xp33_ASAP7_75t_L g228 ( 
.A(n_202),
.B(n_209),
.Y(n_228)
);

OAI22xp5_ASAP7_75t_L g227 ( 
.A1(n_203),
.A2(n_206),
.B1(n_212),
.B2(n_221),
.Y(n_227)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_188),
.Y(n_204)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_204),
.Y(n_231)
);

MAJIxp5_ASAP7_75t_L g205 ( 
.A(n_163),
.B(n_184),
.C(n_192),
.Y(n_205)
);

AOI21xp5_ASAP7_75t_L g226 ( 
.A1(n_207),
.A2(n_223),
.B(n_224),
.Y(n_226)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_171),
.Y(n_208)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_208),
.Y(n_245)
);

INVxp33_ASAP7_75t_L g209 ( 
.A(n_175),
.Y(n_209)
);

XNOR2x2_ASAP7_75t_L g210 ( 
.A(n_169),
.B(n_137),
.Y(n_210)
);

A2O1A1O1Ixp25_ASAP7_75t_L g243 ( 
.A1(n_210),
.A2(n_217),
.B(n_191),
.C(n_168),
.D(n_194),
.Y(n_243)
);

MAJIxp5_ASAP7_75t_L g211 ( 
.A(n_184),
.B(n_161),
.C(n_147),
.Y(n_211)
);

AOI22xp5_ASAP7_75t_L g212 ( 
.A1(n_181),
.A2(n_0),
.B1(n_3),
.B2(n_4),
.Y(n_212)
);

MAJIxp5_ASAP7_75t_L g213 ( 
.A(n_190),
.B(n_189),
.C(n_162),
.Y(n_213)
);

MAJIxp5_ASAP7_75t_L g244 ( 
.A(n_213),
.B(n_183),
.C(n_172),
.Y(n_244)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_171),
.Y(n_215)
);

CKINVDCx20_ASAP7_75t_R g235 ( 
.A(n_215),
.Y(n_235)
);

NAND2xp5_ASAP7_75t_L g216 ( 
.A(n_162),
.B(n_26),
.Y(n_216)
);

FAx1_ASAP7_75t_SL g217 ( 
.A(n_173),
.B(n_17),
.CI(n_15),
.CON(n_217),
.SN(n_217)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_172),
.Y(n_218)
);

CKINVDCx20_ASAP7_75t_R g241 ( 
.A(n_218),
.Y(n_241)
);

CKINVDCx16_ASAP7_75t_R g220 ( 
.A(n_166),
.Y(n_220)
);

HB1xp67_ASAP7_75t_L g238 ( 
.A(n_220),
.Y(n_238)
);

NAND2xp5_ASAP7_75t_L g221 ( 
.A(n_177),
.B(n_0),
.Y(n_221)
);

CKINVDCx20_ASAP7_75t_R g223 ( 
.A(n_166),
.Y(n_223)
);

AND2x2_ASAP7_75t_SL g224 ( 
.A(n_169),
.B(n_3),
.Y(n_224)
);

OAI21xp5_ASAP7_75t_SL g225 ( 
.A1(n_181),
.A2(n_4),
.B(n_5),
.Y(n_225)
);

XNOR2xp5_ASAP7_75t_L g233 ( 
.A(n_225),
.B(n_187),
.Y(n_233)
);

XNOR2xp5_ASAP7_75t_SL g262 ( 
.A(n_233),
.B(n_222),
.Y(n_262)
);

XOR2xp5_ASAP7_75t_L g234 ( 
.A(n_205),
.B(n_180),
.Y(n_234)
);

XOR2xp5_ASAP7_75t_L g256 ( 
.A(n_234),
.B(n_240),
.Y(n_256)
);

OAI22xp5_ASAP7_75t_L g236 ( 
.A1(n_203),
.A2(n_185),
.B1(n_170),
.B2(n_164),
.Y(n_236)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_236),
.Y(n_257)
);

INVx2_ASAP7_75t_L g237 ( 
.A(n_224),
.Y(n_237)
);

NAND2xp5_ASAP7_75t_L g255 ( 
.A(n_237),
.B(n_228),
.Y(n_255)
);

XNOR2xp5_ASAP7_75t_SL g240 ( 
.A(n_210),
.B(n_178),
.Y(n_240)
);

OAI22xp5_ASAP7_75t_L g242 ( 
.A1(n_223),
.A2(n_174),
.B1(n_179),
.B2(n_193),
.Y(n_242)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_242),
.Y(n_266)
);

OAI21xp5_ASAP7_75t_SL g251 ( 
.A1(n_243),
.A2(n_196),
.B(n_201),
.Y(n_251)
);

MAJIxp5_ASAP7_75t_L g252 ( 
.A(n_244),
.B(n_247),
.C(n_248),
.Y(n_252)
);

NAND3xp33_ASAP7_75t_L g246 ( 
.A(n_225),
.B(n_4),
.C(n_5),
.Y(n_246)
);

CKINVDCx20_ASAP7_75t_R g269 ( 
.A(n_246),
.Y(n_269)
);

MAJIxp5_ASAP7_75t_L g247 ( 
.A(n_211),
.B(n_4),
.C(n_5),
.Y(n_247)
);

MAJIxp5_ASAP7_75t_L g248 ( 
.A(n_210),
.B(n_6),
.C(n_7),
.Y(n_248)
);

OAI22xp5_ASAP7_75t_L g249 ( 
.A1(n_206),
.A2(n_6),
.B1(n_7),
.B2(n_8),
.Y(n_249)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_249),
.Y(n_270)
);

XNOR2xp5_ASAP7_75t_L g250 ( 
.A(n_214),
.B(n_6),
.Y(n_250)
);

XNOR2xp5_ASAP7_75t_L g253 ( 
.A(n_250),
.B(n_214),
.Y(n_253)
);

XNOR2xp5_ASAP7_75t_L g280 ( 
.A(n_251),
.B(n_253),
.Y(n_280)
);

AOI21xp5_ASAP7_75t_L g254 ( 
.A1(n_239),
.A2(n_207),
.B(n_219),
.Y(n_254)
);

AOI21xp5_ASAP7_75t_SL g272 ( 
.A1(n_254),
.A2(n_267),
.B(n_226),
.Y(n_272)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_255),
.Y(n_277)
);

AOI22xp5_ASAP7_75t_L g258 ( 
.A1(n_227),
.A2(n_219),
.B1(n_222),
.B2(n_200),
.Y(n_258)
);

OAI22xp5_ASAP7_75t_SL g278 ( 
.A1(n_258),
.A2(n_259),
.B1(n_237),
.B2(n_229),
.Y(n_278)
);

AOI22xp5_ASAP7_75t_SL g259 ( 
.A1(n_248),
.A2(n_198),
.B1(n_195),
.B2(n_213),
.Y(n_259)
);

MAJIxp5_ASAP7_75t_L g260 ( 
.A(n_244),
.B(n_195),
.C(n_216),
.Y(n_260)
);

MAJIxp5_ASAP7_75t_L g273 ( 
.A(n_260),
.B(n_261),
.C(n_247),
.Y(n_273)
);

MAJIxp5_ASAP7_75t_L g261 ( 
.A(n_232),
.B(n_234),
.C(n_240),
.Y(n_261)
);

XOR2xp5_ASAP7_75t_L g285 ( 
.A(n_262),
.B(n_250),
.Y(n_285)
);

NAND2xp5_ASAP7_75t_L g263 ( 
.A(n_235),
.B(n_221),
.Y(n_263)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_263),
.Y(n_279)
);

INVx2_ASAP7_75t_L g264 ( 
.A(n_238),
.Y(n_264)
);

NAND2xp5_ASAP7_75t_L g284 ( 
.A(n_264),
.B(n_231),
.Y(n_284)
);

OAI22x1_ASAP7_75t_L g265 ( 
.A1(n_239),
.A2(n_217),
.B1(n_224),
.B2(n_202),
.Y(n_265)
);

OAI22xp5_ASAP7_75t_L g283 ( 
.A1(n_265),
.A2(n_245),
.B1(n_229),
.B2(n_231),
.Y(n_283)
);

NOR2x1_ASAP7_75t_R g267 ( 
.A(n_243),
.B(n_217),
.Y(n_267)
);

NAND2xp5_ASAP7_75t_L g268 ( 
.A(n_235),
.B(n_218),
.Y(n_268)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_268),
.Y(n_281)
);

FAx1_ASAP7_75t_SL g271 ( 
.A(n_256),
.B(n_233),
.CI(n_232),
.CON(n_271),
.SN(n_271)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_271),
.Y(n_289)
);

XNOR2xp5_ASAP7_75t_L g296 ( 
.A(n_272),
.B(n_273),
.Y(n_296)
);

NAND2xp5_ASAP7_75t_SL g274 ( 
.A(n_269),
.B(n_230),
.Y(n_274)
);

NOR2xp33_ASAP7_75t_L g299 ( 
.A(n_274),
.B(n_278),
.Y(n_299)
);

NAND2xp5_ASAP7_75t_L g275 ( 
.A(n_263),
.B(n_241),
.Y(n_275)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_275),
.Y(n_294)
);

XNOR2x1_ASAP7_75t_SL g276 ( 
.A(n_265),
.B(n_226),
.Y(n_276)
);

AOI21xp5_ASAP7_75t_L g293 ( 
.A1(n_276),
.A2(n_251),
.B(n_268),
.Y(n_293)
);

MAJIxp5_ASAP7_75t_L g282 ( 
.A(n_260),
.B(n_245),
.C(n_241),
.Y(n_282)
);

MAJIxp5_ASAP7_75t_L g290 ( 
.A(n_282),
.B(n_286),
.C(n_288),
.Y(n_290)
);

NAND2xp5_ASAP7_75t_L g302 ( 
.A(n_283),
.B(n_285),
.Y(n_302)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_284),
.Y(n_300)
);

XOR2xp5_ASAP7_75t_L g286 ( 
.A(n_256),
.B(n_212),
.Y(n_286)
);

AOI22xp5_ASAP7_75t_L g287 ( 
.A1(n_266),
.A2(n_215),
.B1(n_208),
.B2(n_204),
.Y(n_287)
);

OAI22xp5_ASAP7_75t_SL g295 ( 
.A1(n_287),
.A2(n_258),
.B1(n_254),
.B2(n_255),
.Y(n_295)
);

MAJIxp5_ASAP7_75t_L g288 ( 
.A(n_261),
.B(n_6),
.C(n_7),
.Y(n_288)
);

OAI22xp5_ASAP7_75t_L g291 ( 
.A1(n_276),
.A2(n_257),
.B1(n_270),
.B2(n_267),
.Y(n_291)
);

AOI22xp5_ASAP7_75t_L g307 ( 
.A1(n_291),
.A2(n_280),
.B1(n_286),
.B2(n_285),
.Y(n_307)
);

MAJIxp5_ASAP7_75t_L g292 ( 
.A(n_282),
.B(n_252),
.C(n_259),
.Y(n_292)
);

MAJIxp5_ASAP7_75t_L g310 ( 
.A(n_292),
.B(n_298),
.C(n_14),
.Y(n_310)
);

XOR2xp5_ASAP7_75t_L g304 ( 
.A(n_293),
.B(n_272),
.Y(n_304)
);

AOI22xp5_ASAP7_75t_L g303 ( 
.A1(n_295),
.A2(n_278),
.B1(n_279),
.B2(n_277),
.Y(n_303)
);

INVx1_ASAP7_75t_SL g297 ( 
.A(n_281),
.Y(n_297)
);

NAND2xp5_ASAP7_75t_L g309 ( 
.A(n_297),
.B(n_253),
.Y(n_309)
);

MAJIxp5_ASAP7_75t_L g298 ( 
.A(n_273),
.B(n_252),
.C(n_262),
.Y(n_298)
);

INVx11_ASAP7_75t_L g301 ( 
.A(n_275),
.Y(n_301)
);

NOR2xp33_ASAP7_75t_L g305 ( 
.A(n_301),
.B(n_287),
.Y(n_305)
);

NAND2xp5_ASAP7_75t_L g313 ( 
.A(n_303),
.B(n_308),
.Y(n_313)
);

NAND2xp5_ASAP7_75t_SL g316 ( 
.A(n_304),
.B(n_307),
.Y(n_316)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_305),
.Y(n_320)
);

OAI21xp5_ASAP7_75t_SL g306 ( 
.A1(n_289),
.A2(n_271),
.B(n_288),
.Y(n_306)
);

CKINVDCx14_ASAP7_75t_R g319 ( 
.A(n_306),
.Y(n_319)
);

AOI22xp5_ASAP7_75t_L g308 ( 
.A1(n_299),
.A2(n_280),
.B1(n_264),
.B2(n_271),
.Y(n_308)
);

NAND2xp5_ASAP7_75t_L g315 ( 
.A(n_309),
.B(n_311),
.Y(n_315)
);

MAJIxp5_ASAP7_75t_L g317 ( 
.A(n_310),
.B(n_292),
.C(n_298),
.Y(n_317)
);

NAND2xp5_ASAP7_75t_SL g311 ( 
.A(n_296),
.B(n_9),
.Y(n_311)
);

XOR2xp5_ASAP7_75t_L g312 ( 
.A(n_296),
.B(n_290),
.Y(n_312)
);

NOR2xp33_ASAP7_75t_L g314 ( 
.A(n_312),
.B(n_290),
.Y(n_314)
);

AOI21xp5_ASAP7_75t_L g325 ( 
.A1(n_314),
.A2(n_318),
.B(n_302),
.Y(n_325)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_317),
.Y(n_323)
);

OAI21xp5_ASAP7_75t_SL g318 ( 
.A1(n_304),
.A2(n_293),
.B(n_294),
.Y(n_318)
);

NOR2xp33_ASAP7_75t_SL g321 ( 
.A(n_317),
.B(n_310),
.Y(n_321)
);

MAJIxp5_ASAP7_75t_L g326 ( 
.A(n_321),
.B(n_324),
.C(n_325),
.Y(n_326)
);

OAI21x1_ASAP7_75t_L g322 ( 
.A1(n_319),
.A2(n_312),
.B(n_316),
.Y(n_322)
);

OAI21xp33_ASAP7_75t_SL g328 ( 
.A1(n_322),
.A2(n_303),
.B(n_302),
.Y(n_328)
);

OAI21xp5_ASAP7_75t_L g324 ( 
.A1(n_318),
.A2(n_294),
.B(n_300),
.Y(n_324)
);

MAJIxp5_ASAP7_75t_L g327 ( 
.A(n_323),
.B(n_313),
.C(n_320),
.Y(n_327)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_327),
.Y(n_329)
);

AOI21xp5_ASAP7_75t_L g330 ( 
.A1(n_329),
.A2(n_328),
.B(n_326),
.Y(n_330)
);

FAx1_ASAP7_75t_SL g331 ( 
.A(n_330),
.B(n_295),
.CI(n_301),
.CON(n_331),
.SN(n_331)
);

NAND2xp5_ASAP7_75t_SL g332 ( 
.A(n_331),
.B(n_297),
.Y(n_332)
);

OAI22xp5_ASAP7_75t_L g333 ( 
.A1(n_332),
.A2(n_300),
.B1(n_315),
.B2(n_331),
.Y(n_333)
);

AOI21xp5_ASAP7_75t_L g334 ( 
.A1(n_333),
.A2(n_9),
.B(n_10),
.Y(n_334)
);


endmodule