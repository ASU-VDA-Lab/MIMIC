module fake_netlist_6_3099_n_776 (n_52, n_16, n_1, n_91, n_119, n_46, n_146, n_18, n_21, n_147, n_154, n_88, n_3, n_98, n_113, n_39, n_63, n_73, n_4, n_148, n_138, n_22, n_68, n_28, n_50, n_158, n_49, n_7, n_83, n_5, n_101, n_144, n_127, n_125, n_153, n_77, n_156, n_149, n_152, n_106, n_92, n_145, n_42, n_133, n_96, n_8, n_90, n_24, n_105, n_131, n_54, n_132, n_102, n_0, n_87, n_32, n_66, n_85, n_99, n_78, n_84, n_130, n_100, n_129, n_13, n_121, n_11, n_137, n_17, n_23, n_142, n_20, n_143, n_2, n_19, n_47, n_62, n_29, n_155, n_75, n_109, n_150, n_122, n_45, n_34, n_140, n_70, n_120, n_37, n_15, n_67, n_33, n_82, n_27, n_38, n_110, n_151, n_61, n_112, n_81, n_59, n_76, n_36, n_26, n_124, n_55, n_126, n_94, n_97, n_108, n_58, n_116, n_64, n_117, n_118, n_48, n_65, n_25, n_40, n_93, n_80, n_141, n_135, n_139, n_41, n_134, n_114, n_86, n_104, n_95, n_9, n_107, n_10, n_71, n_74, n_6, n_14, n_123, n_136, n_72, n_89, n_103, n_111, n_60, n_157, n_35, n_115, n_12, n_69, n_128, n_30, n_79, n_43, n_31, n_57, n_53, n_51, n_44, n_56, n_776);

input n_52;
input n_16;
input n_1;
input n_91;
input n_119;
input n_46;
input n_146;
input n_18;
input n_21;
input n_147;
input n_154;
input n_88;
input n_3;
input n_98;
input n_113;
input n_39;
input n_63;
input n_73;
input n_4;
input n_148;
input n_138;
input n_22;
input n_68;
input n_28;
input n_50;
input n_158;
input n_49;
input n_7;
input n_83;
input n_5;
input n_101;
input n_144;
input n_127;
input n_125;
input n_153;
input n_77;
input n_156;
input n_149;
input n_152;
input n_106;
input n_92;
input n_145;
input n_42;
input n_133;
input n_96;
input n_8;
input n_90;
input n_24;
input n_105;
input n_131;
input n_54;
input n_132;
input n_102;
input n_0;
input n_87;
input n_32;
input n_66;
input n_85;
input n_99;
input n_78;
input n_84;
input n_130;
input n_100;
input n_129;
input n_13;
input n_121;
input n_11;
input n_137;
input n_17;
input n_23;
input n_142;
input n_20;
input n_143;
input n_2;
input n_19;
input n_47;
input n_62;
input n_29;
input n_155;
input n_75;
input n_109;
input n_150;
input n_122;
input n_45;
input n_34;
input n_140;
input n_70;
input n_120;
input n_37;
input n_15;
input n_67;
input n_33;
input n_82;
input n_27;
input n_38;
input n_110;
input n_151;
input n_61;
input n_112;
input n_81;
input n_59;
input n_76;
input n_36;
input n_26;
input n_124;
input n_55;
input n_126;
input n_94;
input n_97;
input n_108;
input n_58;
input n_116;
input n_64;
input n_117;
input n_118;
input n_48;
input n_65;
input n_25;
input n_40;
input n_93;
input n_80;
input n_141;
input n_135;
input n_139;
input n_41;
input n_134;
input n_114;
input n_86;
input n_104;
input n_95;
input n_9;
input n_107;
input n_10;
input n_71;
input n_74;
input n_6;
input n_14;
input n_123;
input n_136;
input n_72;
input n_89;
input n_103;
input n_111;
input n_60;
input n_157;
input n_35;
input n_115;
input n_12;
input n_69;
input n_128;
input n_30;
input n_79;
input n_43;
input n_31;
input n_57;
input n_53;
input n_51;
input n_44;
input n_56;

output n_776;

wire n_591;
wire n_435;
wire n_326;
wire n_256;
wire n_440;
wire n_587;
wire n_695;
wire n_507;
wire n_580;
wire n_762;
wire n_209;
wire n_367;
wire n_465;
wire n_680;
wire n_741;
wire n_760;
wire n_590;
wire n_625;
wire n_661;
wire n_223;
wire n_278;
wire n_341;
wire n_362;
wire n_226;
wire n_161;
wire n_208;
wire n_462;
wire n_607;
wire n_671;
wire n_726;
wire n_316;
wire n_419;
wire n_304;
wire n_212;
wire n_700;
wire n_694;
wire n_740;
wire n_578;
wire n_703;
wire n_365;
wire n_168;
wire n_384;
wire n_297;
wire n_595;
wire n_627;
wire n_524;
wire n_342;
wire n_725;
wire n_358;
wire n_160;
wire n_751;
wire n_449;
wire n_749;
wire n_188;
wire n_310;
wire n_509;
wire n_186;
wire n_245;
wire n_368;
wire n_575;
wire n_677;
wire n_396;
wire n_495;
wire n_350;
wire n_585;
wire n_732;
wire n_568;
wire n_392;
wire n_442;
wire n_480;
wire n_724;
wire n_382;
wire n_673;
wire n_180;
wire n_628;
wire n_557;
wire n_349;
wire n_643;
wire n_233;
wire n_698;
wire n_617;
wire n_255;
wire n_739;
wire n_284;
wire n_400;
wire n_337;
wire n_214;
wire n_485;
wire n_443;
wire n_246;
wire n_768;
wire n_471;
wire n_289;
wire n_421;
wire n_424;
wire n_615;
wire n_181;
wire n_182;
wire n_238;
wire n_573;
wire n_769;
wire n_202;
wire n_320;
wire n_639;
wire n_676;
wire n_327;
wire n_727;
wire n_369;
wire n_597;
wire n_685;
wire n_280;
wire n_287;
wire n_353;
wire n_610;
wire n_555;
wire n_389;
wire n_415;
wire n_230;
wire n_605;
wire n_461;
wire n_383;
wire n_669;
wire n_200;
wire n_447;
wire n_176;
wire n_198;
wire n_300;
wire n_222;
wire n_179;
wire n_248;
wire n_517;
wire n_718;
wire n_747;
wire n_667;
wire n_229;
wire n_542;
wire n_644;
wire n_682;
wire n_621;
wire n_305;
wire n_721;
wire n_750;
wire n_532;
wire n_742;
wire n_173;
wire n_535;
wire n_691;
wire n_250;
wire n_372;
wire n_468;
wire n_544;
wire n_504;
wire n_314;
wire n_378;
wire n_413;
wire n_377;
wire n_183;
wire n_510;
wire n_375;
wire n_601;
wire n_338;
wire n_522;
wire n_466;
wire n_704;
wire n_748;
wire n_506;
wire n_763;
wire n_360;
wire n_603;
wire n_235;
wire n_536;
wire n_622;
wire n_191;
wire n_340;
wire n_710;
wire n_387;
wire n_452;
wire n_616;
wire n_658;
wire n_744;
wire n_344;
wire n_581;
wire n_428;
wire n_761;
wire n_746;
wire n_609;
wire n_765;
wire n_432;
wire n_641;
wire n_693;
wire n_167;
wire n_631;
wire n_174;
wire n_516;
wire n_720;
wire n_525;
wire n_758;
wire n_611;
wire n_491;
wire n_656;
wire n_772;
wire n_666;
wire n_371;
wire n_770;
wire n_567;
wire n_189;
wire n_738;
wire n_405;
wire n_213;
wire n_538;
wire n_294;
wire n_302;
wire n_499;
wire n_380;
wire n_705;
wire n_647;
wire n_197;
wire n_343;
wire n_448;
wire n_494;
wire n_539;
wire n_493;
wire n_397;
wire n_614;
wire n_529;
wire n_445;
wire n_425;
wire n_684;
wire n_454;
wire n_218;
wire n_638;
wire n_234;
wire n_486;
wire n_381;
wire n_236;
wire n_653;
wire n_752;
wire n_172;
wire n_713;
wire n_648;
wire n_657;
wire n_576;
wire n_472;
wire n_270;
wire n_239;
wire n_414;
wire n_563;
wire n_490;
wire n_290;
wire n_220;
wire n_224;
wire n_734;
wire n_708;
wire n_196;
wire n_402;
wire n_352;
wire n_668;
wire n_478;
wire n_626;
wire n_574;
wire n_460;
wire n_417;
wire n_446;
wire n_498;
wire n_662;
wire n_374;
wire n_659;
wire n_709;
wire n_366;
wire n_407;
wire n_450;
wire n_272;
wire n_526;
wire n_185;
wire n_712;
wire n_348;
wire n_711;
wire n_579;
wire n_376;
wire n_390;
wire n_473;
wire n_293;
wire n_334;
wire n_559;
wire n_370;
wire n_458;
wire n_232;
wire n_650;
wire n_163;
wire n_717;
wire n_330;
wire n_771;
wire n_470;
wire n_475;
wire n_298;
wire n_492;
wire n_281;
wire n_258;
wire n_551;
wire n_699;
wire n_456;
wire n_564;
wire n_260;
wire n_265;
wire n_313;
wire n_451;
wire n_624;
wire n_279;
wire n_686;
wire n_252;
wire n_757;
wire n_228;
wire n_565;
wire n_594;
wire n_719;
wire n_356;
wire n_577;
wire n_166;
wire n_184;
wire n_552;
wire n_619;
wire n_216;
wire n_455;
wire n_521;
wire n_363;
wire n_572;
wire n_395;
wire n_592;
wire n_745;
wire n_654;
wire n_323;
wire n_606;
wire n_393;
wire n_411;
wire n_503;
wire n_716;
wire n_623;
wire n_599;
wire n_513;
wire n_321;
wire n_645;
wire n_331;
wire n_227;
wire n_570;
wire n_731;
wire n_406;
wire n_483;
wire n_735;
wire n_204;
wire n_482;
wire n_755;
wire n_474;
wire n_527;
wire n_261;
wire n_608;
wire n_620;
wire n_420;
wire n_683;
wire n_630;
wire n_312;
wire n_394;
wire n_519;
wire n_541;
wire n_512;
wire n_292;
wire n_164;
wire n_307;
wire n_469;
wire n_433;
wire n_500;
wire n_476;
wire n_714;
wire n_291;
wire n_219;
wire n_543;
wire n_357;
wire n_264;
wire n_263;
wire n_589;
wire n_481;
wire n_325;
wire n_767;
wire n_329;
wire n_464;
wire n_600;
wire n_561;
wire n_477;
wire n_549;
wire n_533;
wire n_408;
wire n_237;
wire n_584;
wire n_244;
wire n_399;
wire n_243;
wire n_548;
wire n_282;
wire n_436;
wire n_211;
wire n_523;
wire n_175;
wire n_322;
wire n_707;
wire n_345;
wire n_409;
wire n_231;
wire n_354;
wire n_689;
wire n_505;
wire n_240;
wire n_756;
wire n_319;
wire n_547;
wire n_537;
wire n_273;
wire n_558;
wire n_635;
wire n_311;
wire n_403;
wire n_723;
wire n_253;
wire n_634;
wire n_583;
wire n_596;
wire n_546;
wire n_562;
wire n_249;
wire n_201;
wire n_386;
wire n_764;
wire n_556;
wire n_159;
wire n_162;
wire n_692;
wire n_733;
wire n_754;
wire n_487;
wire n_550;
wire n_241;
wire n_275;
wire n_553;
wire n_652;
wire n_560;
wire n_753;
wire n_642;
wire n_276;
wire n_569;
wire n_441;
wire n_221;
wire n_444;
wire n_586;
wire n_423;
wire n_737;
wire n_318;
wire n_303;
wire n_511;
wire n_715;
wire n_467;
wire n_306;
wire n_193;
wire n_269;
wire n_359;
wire n_346;
wire n_416;
wire n_530;
wire n_277;
wire n_520;
wire n_418;
wire n_618;
wire n_582;
wire n_199;
wire n_266;
wire n_296;
wire n_674;
wire n_775;
wire n_571;
wire n_268;
wire n_271;
wire n_404;
wire n_651;
wire n_439;
wire n_217;
wire n_210;
wire n_299;
wire n_518;
wire n_206;
wire n_679;
wire n_453;
wire n_612;
wire n_633;
wire n_665;
wire n_333;
wire n_588;
wire n_215;
wire n_178;
wire n_247;
wire n_225;
wire n_308;
wire n_309;
wire n_759;
wire n_355;
wire n_426;
wire n_317;
wire n_632;
wire n_702;
wire n_431;
wire n_347;
wire n_459;
wire n_502;
wire n_328;
wire n_672;
wire n_534;
wire n_488;
wire n_429;
wire n_373;
wire n_195;
wire n_285;
wire n_497;
wire n_773;
wire n_675;
wire n_257;
wire n_730;
wire n_655;
wire n_706;
wire n_670;
wire n_203;
wire n_286;
wire n_254;
wire n_207;
wire n_242;
wire n_690;
wire n_401;
wire n_324;
wire n_743;
wire n_766;
wire n_335;
wire n_430;
wire n_463;
wire n_545;
wire n_489;
wire n_205;
wire n_604;
wire n_251;
wire n_301;
wire n_274;
wire n_636;
wire n_728;
wire n_681;
wire n_729;
wire n_774;
wire n_412;
wire n_640;
wire n_660;
wire n_267;
wire n_438;
wire n_339;
wire n_315;
wire n_434;
wire n_515;
wire n_288;
wire n_427;
wire n_479;
wire n_496;
wire n_598;
wire n_422;
wire n_696;
wire n_722;
wire n_688;
wire n_165;
wire n_351;
wire n_437;
wire n_259;
wire n_177;
wire n_540;
wire n_593;
wire n_514;
wire n_646;
wire n_528;
wire n_391;
wire n_457;
wire n_687;
wire n_697;
wire n_364;
wire n_637;
wire n_295;
wire n_385;
wire n_701;
wire n_629;
wire n_388;
wire n_190;
wire n_262;
wire n_484;
wire n_613;
wire n_736;
wire n_187;
wire n_501;
wire n_531;
wire n_361;
wire n_508;
wire n_663;
wire n_379;
wire n_170;
wire n_332;
wire n_336;
wire n_410;
wire n_398;
wire n_566;
wire n_554;
wire n_602;
wire n_194;
wire n_664;
wire n_171;
wire n_678;
wire n_192;
wire n_169;
wire n_649;
wire n_283;

CKINVDCx5p33_ASAP7_75t_R g159 ( 
.A(n_22),
.Y(n_159)
);

CKINVDCx5p33_ASAP7_75t_R g160 ( 
.A(n_15),
.Y(n_160)
);

CKINVDCx5p33_ASAP7_75t_R g161 ( 
.A(n_127),
.Y(n_161)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_146),
.Y(n_162)
);

BUFx3_ASAP7_75t_L g163 ( 
.A(n_21),
.Y(n_163)
);

CKINVDCx5p33_ASAP7_75t_R g164 ( 
.A(n_40),
.Y(n_164)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_136),
.Y(n_165)
);

INVx2_ASAP7_75t_L g166 ( 
.A(n_64),
.Y(n_166)
);

INVxp67_ASAP7_75t_L g167 ( 
.A(n_30),
.Y(n_167)
);

BUFx10_ASAP7_75t_L g168 ( 
.A(n_125),
.Y(n_168)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_119),
.Y(n_169)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_138),
.Y(n_170)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_42),
.Y(n_171)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_72),
.Y(n_172)
);

CKINVDCx5p33_ASAP7_75t_R g173 ( 
.A(n_26),
.Y(n_173)
);

CKINVDCx5p33_ASAP7_75t_R g174 ( 
.A(n_32),
.Y(n_174)
);

CKINVDCx16_ASAP7_75t_R g175 ( 
.A(n_139),
.Y(n_175)
);

CKINVDCx5p33_ASAP7_75t_R g176 ( 
.A(n_106),
.Y(n_176)
);

BUFx6f_ASAP7_75t_L g177 ( 
.A(n_110),
.Y(n_177)
);

BUFx10_ASAP7_75t_L g178 ( 
.A(n_149),
.Y(n_178)
);

INVx2_ASAP7_75t_L g179 ( 
.A(n_38),
.Y(n_179)
);

HB1xp67_ASAP7_75t_L g180 ( 
.A(n_142),
.Y(n_180)
);

CKINVDCx5p33_ASAP7_75t_R g181 ( 
.A(n_111),
.Y(n_181)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_47),
.Y(n_182)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_61),
.Y(n_183)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_66),
.Y(n_184)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_23),
.Y(n_185)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_140),
.Y(n_186)
);

CKINVDCx5p33_ASAP7_75t_R g187 ( 
.A(n_59),
.Y(n_187)
);

BUFx6f_ASAP7_75t_L g188 ( 
.A(n_25),
.Y(n_188)
);

CKINVDCx5p33_ASAP7_75t_R g189 ( 
.A(n_17),
.Y(n_189)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_87),
.Y(n_190)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_46),
.Y(n_191)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_117),
.Y(n_192)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_93),
.Y(n_193)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_68),
.Y(n_194)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_133),
.Y(n_195)
);

INVxp33_ASAP7_75t_SL g196 ( 
.A(n_152),
.Y(n_196)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_33),
.Y(n_197)
);

CKINVDCx20_ASAP7_75t_R g198 ( 
.A(n_12),
.Y(n_198)
);

INVx2_ASAP7_75t_SL g199 ( 
.A(n_67),
.Y(n_199)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_8),
.Y(n_200)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_101),
.Y(n_201)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_55),
.Y(n_202)
);

BUFx2_ASAP7_75t_L g203 ( 
.A(n_92),
.Y(n_203)
);

CKINVDCx16_ASAP7_75t_R g204 ( 
.A(n_102),
.Y(n_204)
);

CKINVDCx5p33_ASAP7_75t_R g205 ( 
.A(n_24),
.Y(n_205)
);

CKINVDCx5p33_ASAP7_75t_R g206 ( 
.A(n_105),
.Y(n_206)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_108),
.Y(n_207)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_88),
.Y(n_208)
);

CKINVDCx5p33_ASAP7_75t_R g209 ( 
.A(n_113),
.Y(n_209)
);

CKINVDCx5p33_ASAP7_75t_R g210 ( 
.A(n_37),
.Y(n_210)
);

INVx2_ASAP7_75t_L g211 ( 
.A(n_71),
.Y(n_211)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_95),
.Y(n_212)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_137),
.Y(n_213)
);

CKINVDCx5p33_ASAP7_75t_R g214 ( 
.A(n_6),
.Y(n_214)
);

NAND2xp5_ASAP7_75t_L g215 ( 
.A(n_180),
.B(n_0),
.Y(n_215)
);

BUFx6f_ASAP7_75t_L g216 ( 
.A(n_177),
.Y(n_216)
);

NAND2xp5_ASAP7_75t_L g217 ( 
.A(n_180),
.B(n_203),
.Y(n_217)
);

OAI21x1_ASAP7_75t_L g218 ( 
.A1(n_211),
.A2(n_79),
.B(n_157),
.Y(n_218)
);

BUFx3_ASAP7_75t_L g219 ( 
.A(n_163),
.Y(n_219)
);

HB1xp67_ASAP7_75t_L g220 ( 
.A(n_200),
.Y(n_220)
);

INVx2_ASAP7_75t_SL g221 ( 
.A(n_168),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_SL g222 ( 
.A(n_175),
.B(n_0),
.Y(n_222)
);

INVx5_ASAP7_75t_L g223 ( 
.A(n_177),
.Y(n_223)
);

AND2x4_ASAP7_75t_L g224 ( 
.A(n_163),
.B(n_1),
.Y(n_224)
);

INVx2_ASAP7_75t_L g225 ( 
.A(n_177),
.Y(n_225)
);

AND2x4_ASAP7_75t_L g226 ( 
.A(n_166),
.B(n_1),
.Y(n_226)
);

OAI22xp5_ASAP7_75t_SL g227 ( 
.A1(n_198),
.A2(n_2),
.B1(n_3),
.B2(n_4),
.Y(n_227)
);

BUFx6f_ASAP7_75t_L g228 ( 
.A(n_177),
.Y(n_228)
);

BUFx6f_ASAP7_75t_L g229 ( 
.A(n_188),
.Y(n_229)
);

AND2x2_ASAP7_75t_L g230 ( 
.A(n_204),
.B(n_2),
.Y(n_230)
);

OA21x2_ASAP7_75t_L g231 ( 
.A1(n_166),
.A2(n_179),
.B(n_165),
.Y(n_231)
);

CKINVDCx20_ASAP7_75t_R g232 ( 
.A(n_198),
.Y(n_232)
);

OAI22x1_ASAP7_75t_SL g233 ( 
.A1(n_214),
.A2(n_3),
.B1(n_4),
.B2(n_5),
.Y(n_233)
);

INVx6_ASAP7_75t_L g234 ( 
.A(n_168),
.Y(n_234)
);

BUFx6f_ASAP7_75t_L g235 ( 
.A(n_188),
.Y(n_235)
);

HB1xp67_ASAP7_75t_L g236 ( 
.A(n_167),
.Y(n_236)
);

AND2x2_ASAP7_75t_L g237 ( 
.A(n_178),
.B(n_5),
.Y(n_237)
);

OAI22x1_ASAP7_75t_L g238 ( 
.A1(n_167),
.A2(n_6),
.B1(n_7),
.B2(n_8),
.Y(n_238)
);

HB1xp67_ASAP7_75t_L g239 ( 
.A(n_162),
.Y(n_239)
);

AOI22x1_ASAP7_75t_SL g240 ( 
.A1(n_169),
.A2(n_7),
.B1(n_9),
.B2(n_10),
.Y(n_240)
);

NOR2xp33_ASAP7_75t_L g241 ( 
.A(n_179),
.B(n_9),
.Y(n_241)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_170),
.Y(n_242)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_171),
.Y(n_243)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_172),
.Y(n_244)
);

INVx2_ASAP7_75t_L g245 ( 
.A(n_188),
.Y(n_245)
);

INVx2_ASAP7_75t_L g246 ( 
.A(n_188),
.Y(n_246)
);

BUFx2_ASAP7_75t_L g247 ( 
.A(n_182),
.Y(n_247)
);

OA21x2_ASAP7_75t_L g248 ( 
.A1(n_183),
.A2(n_10),
.B(n_11),
.Y(n_248)
);

INVx2_ASAP7_75t_L g249 ( 
.A(n_184),
.Y(n_249)
);

INVx6_ASAP7_75t_L g250 ( 
.A(n_178),
.Y(n_250)
);

BUFx6f_ASAP7_75t_L g251 ( 
.A(n_185),
.Y(n_251)
);

BUFx6f_ASAP7_75t_L g252 ( 
.A(n_186),
.Y(n_252)
);

INVx2_ASAP7_75t_L g253 ( 
.A(n_190),
.Y(n_253)
);

BUFx2_ASAP7_75t_L g254 ( 
.A(n_191),
.Y(n_254)
);

BUFx6f_ASAP7_75t_L g255 ( 
.A(n_192),
.Y(n_255)
);

INVx3_ASAP7_75t_L g256 ( 
.A(n_193),
.Y(n_256)
);

HB1xp67_ASAP7_75t_L g257 ( 
.A(n_194),
.Y(n_257)
);

AND2x4_ASAP7_75t_L g258 ( 
.A(n_199),
.B(n_16),
.Y(n_258)
);

INVx3_ASAP7_75t_L g259 ( 
.A(n_216),
.Y(n_259)
);

INVx2_ASAP7_75t_L g260 ( 
.A(n_225),
.Y(n_260)
);

NAND2xp5_ASAP7_75t_SL g261 ( 
.A(n_230),
.B(n_196),
.Y(n_261)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_249),
.Y(n_262)
);

NOR2xp33_ASAP7_75t_L g263 ( 
.A(n_217),
.B(n_234),
.Y(n_263)
);

NAND2xp5_ASAP7_75t_L g264 ( 
.A(n_258),
.B(n_195),
.Y(n_264)
);

INVx2_ASAP7_75t_L g265 ( 
.A(n_225),
.Y(n_265)
);

INVx2_ASAP7_75t_L g266 ( 
.A(n_245),
.Y(n_266)
);

INVx4_ASAP7_75t_L g267 ( 
.A(n_251),
.Y(n_267)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_249),
.Y(n_268)
);

BUFx6f_ASAP7_75t_L g269 ( 
.A(n_216),
.Y(n_269)
);

INVx2_ASAP7_75t_SL g270 ( 
.A(n_234),
.Y(n_270)
);

INVx2_ASAP7_75t_L g271 ( 
.A(n_245),
.Y(n_271)
);

INVx3_ASAP7_75t_L g272 ( 
.A(n_216),
.Y(n_272)
);

BUFx10_ASAP7_75t_L g273 ( 
.A(n_234),
.Y(n_273)
);

NOR2xp33_ASAP7_75t_L g274 ( 
.A(n_250),
.B(n_197),
.Y(n_274)
);

NAND2xp5_ASAP7_75t_SL g275 ( 
.A(n_237),
.B(n_159),
.Y(n_275)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_253),
.Y(n_276)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_253),
.Y(n_277)
);

NAND2xp5_ASAP7_75t_L g278 ( 
.A(n_258),
.B(n_201),
.Y(n_278)
);

INVx2_ASAP7_75t_L g279 ( 
.A(n_246),
.Y(n_279)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_242),
.Y(n_280)
);

OAI22xp33_ASAP7_75t_L g281 ( 
.A1(n_215),
.A2(n_213),
.B1(n_212),
.B2(n_202),
.Y(n_281)
);

AND2x2_ASAP7_75t_L g282 ( 
.A(n_219),
.B(n_160),
.Y(n_282)
);

INVx2_ASAP7_75t_L g283 ( 
.A(n_246),
.Y(n_283)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_243),
.Y(n_284)
);

INVx2_ASAP7_75t_SL g285 ( 
.A(n_250),
.Y(n_285)
);

NAND2xp33_ASAP7_75t_SL g286 ( 
.A(n_222),
.B(n_207),
.Y(n_286)
);

INVx2_ASAP7_75t_L g287 ( 
.A(n_216),
.Y(n_287)
);

AND2x2_ASAP7_75t_L g288 ( 
.A(n_219),
.B(n_221),
.Y(n_288)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_244),
.Y(n_289)
);

INVx2_ASAP7_75t_L g290 ( 
.A(n_228),
.Y(n_290)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_251),
.Y(n_291)
);

NAND2xp5_ASAP7_75t_SL g292 ( 
.A(n_222),
.B(n_161),
.Y(n_292)
);

INVx3_ASAP7_75t_L g293 ( 
.A(n_228),
.Y(n_293)
);

AOI21x1_ASAP7_75t_L g294 ( 
.A1(n_258),
.A2(n_208),
.B(n_209),
.Y(n_294)
);

INVx2_ASAP7_75t_L g295 ( 
.A(n_228),
.Y(n_295)
);

INVx2_ASAP7_75t_L g296 ( 
.A(n_228),
.Y(n_296)
);

INVx2_ASAP7_75t_L g297 ( 
.A(n_229),
.Y(n_297)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_251),
.Y(n_298)
);

INVx2_ASAP7_75t_L g299 ( 
.A(n_229),
.Y(n_299)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_251),
.Y(n_300)
);

OAI22xp33_ASAP7_75t_L g301 ( 
.A1(n_236),
.A2(n_210),
.B1(n_206),
.B2(n_205),
.Y(n_301)
);

INVx2_ASAP7_75t_L g302 ( 
.A(n_229),
.Y(n_302)
);

INVxp33_ASAP7_75t_SL g303 ( 
.A(n_236),
.Y(n_303)
);

INVx2_ASAP7_75t_L g304 ( 
.A(n_229),
.Y(n_304)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_252),
.Y(n_305)
);

NAND2xp5_ASAP7_75t_L g306 ( 
.A(n_247),
.B(n_189),
.Y(n_306)
);

INVx2_ASAP7_75t_L g307 ( 
.A(n_235),
.Y(n_307)
);

NAND2xp5_ASAP7_75t_L g308 ( 
.A(n_263),
.B(n_223),
.Y(n_308)
);

INVxp67_ASAP7_75t_L g309 ( 
.A(n_288),
.Y(n_309)
);

NOR2xp67_ASAP7_75t_SL g310 ( 
.A(n_261),
.B(n_223),
.Y(n_310)
);

INVx2_ASAP7_75t_L g311 ( 
.A(n_259),
.Y(n_311)
);

NAND2xp5_ASAP7_75t_SL g312 ( 
.A(n_286),
.B(n_226),
.Y(n_312)
);

INVx2_ASAP7_75t_L g313 ( 
.A(n_259),
.Y(n_313)
);

NOR2xp33_ASAP7_75t_L g314 ( 
.A(n_261),
.B(n_292),
.Y(n_314)
);

OAI221xp5_ASAP7_75t_L g315 ( 
.A1(n_286),
.A2(n_241),
.B1(n_239),
.B2(n_257),
.C(n_254),
.Y(n_315)
);

AND2x2_ASAP7_75t_L g316 ( 
.A(n_282),
.B(n_273),
.Y(n_316)
);

NAND2xp5_ASAP7_75t_L g317 ( 
.A(n_275),
.B(n_223),
.Y(n_317)
);

NOR2xp67_ASAP7_75t_L g318 ( 
.A(n_270),
.B(n_223),
.Y(n_318)
);

NAND2xp5_ASAP7_75t_L g319 ( 
.A(n_275),
.B(n_224),
.Y(n_319)
);

NAND2xp5_ASAP7_75t_L g320 ( 
.A(n_264),
.B(n_224),
.Y(n_320)
);

NAND2xp5_ASAP7_75t_L g321 ( 
.A(n_278),
.B(n_231),
.Y(n_321)
);

INVx2_ASAP7_75t_L g322 ( 
.A(n_259),
.Y(n_322)
);

NAND2xp5_ASAP7_75t_SL g323 ( 
.A(n_292),
.B(n_226),
.Y(n_323)
);

INVx1_ASAP7_75t_SL g324 ( 
.A(n_303),
.Y(n_324)
);

INVx2_ASAP7_75t_L g325 ( 
.A(n_272),
.Y(n_325)
);

NAND2xp5_ASAP7_75t_L g326 ( 
.A(n_291),
.B(n_231),
.Y(n_326)
);

BUFx6f_ASAP7_75t_L g327 ( 
.A(n_269),
.Y(n_327)
);

NAND2xp5_ASAP7_75t_L g328 ( 
.A(n_298),
.B(n_231),
.Y(n_328)
);

BUFx3_ASAP7_75t_L g329 ( 
.A(n_300),
.Y(n_329)
);

NAND2xp5_ASAP7_75t_SL g330 ( 
.A(n_281),
.B(n_164),
.Y(n_330)
);

NOR2xp33_ASAP7_75t_L g331 ( 
.A(n_306),
.B(n_250),
.Y(n_331)
);

OAI221xp5_ASAP7_75t_L g332 ( 
.A1(n_280),
.A2(n_241),
.B1(n_239),
.B2(n_257),
.C(n_220),
.Y(n_332)
);

BUFx3_ASAP7_75t_L g333 ( 
.A(n_305),
.Y(n_333)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_284),
.Y(n_334)
);

NAND2xp5_ASAP7_75t_L g335 ( 
.A(n_267),
.B(n_256),
.Y(n_335)
);

INVx2_ASAP7_75t_L g336 ( 
.A(n_272),
.Y(n_336)
);

BUFx6f_ASAP7_75t_L g337 ( 
.A(n_269),
.Y(n_337)
);

INVx1_ASAP7_75t_L g338 ( 
.A(n_289),
.Y(n_338)
);

AOI22xp5_ASAP7_75t_L g339 ( 
.A1(n_301),
.A2(n_238),
.B1(n_174),
.B2(n_176),
.Y(n_339)
);

INVx2_ASAP7_75t_L g340 ( 
.A(n_272),
.Y(n_340)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_293),
.Y(n_341)
);

INVx2_ASAP7_75t_L g342 ( 
.A(n_293),
.Y(n_342)
);

INVx2_ASAP7_75t_SL g343 ( 
.A(n_273),
.Y(n_343)
);

NAND2xp33_ASAP7_75t_L g344 ( 
.A(n_260),
.B(n_235),
.Y(n_344)
);

NAND2xp5_ASAP7_75t_L g345 ( 
.A(n_267),
.B(n_293),
.Y(n_345)
);

NAND2xp5_ASAP7_75t_L g346 ( 
.A(n_267),
.B(n_256),
.Y(n_346)
);

INVx1_ASAP7_75t_L g347 ( 
.A(n_287),
.Y(n_347)
);

NAND2xp5_ASAP7_75t_L g348 ( 
.A(n_287),
.B(n_252),
.Y(n_348)
);

INVx1_ASAP7_75t_L g349 ( 
.A(n_290),
.Y(n_349)
);

INVx1_ASAP7_75t_L g350 ( 
.A(n_295),
.Y(n_350)
);

NAND2xp5_ASAP7_75t_L g351 ( 
.A(n_295),
.B(n_252),
.Y(n_351)
);

INVx2_ASAP7_75t_L g352 ( 
.A(n_296),
.Y(n_352)
);

INVx1_ASAP7_75t_L g353 ( 
.A(n_296),
.Y(n_353)
);

INVx1_ASAP7_75t_L g354 ( 
.A(n_297),
.Y(n_354)
);

AND2x2_ASAP7_75t_L g355 ( 
.A(n_273),
.B(n_220),
.Y(n_355)
);

NOR2xp33_ASAP7_75t_R g356 ( 
.A(n_294),
.B(n_173),
.Y(n_356)
);

INVx1_ASAP7_75t_L g357 ( 
.A(n_297),
.Y(n_357)
);

OAI22xp33_ASAP7_75t_L g358 ( 
.A1(n_303),
.A2(n_248),
.B1(n_233),
.B2(n_240),
.Y(n_358)
);

INVx1_ASAP7_75t_L g359 ( 
.A(n_299),
.Y(n_359)
);

NAND2xp5_ASAP7_75t_L g360 ( 
.A(n_299),
.B(n_252),
.Y(n_360)
);

NAND2xp5_ASAP7_75t_L g361 ( 
.A(n_302),
.B(n_255),
.Y(n_361)
);

INVx2_ASAP7_75t_L g362 ( 
.A(n_302),
.Y(n_362)
);

INVxp33_ASAP7_75t_L g363 ( 
.A(n_274),
.Y(n_363)
);

BUFx6f_ASAP7_75t_SL g364 ( 
.A(n_270),
.Y(n_364)
);

INVx2_ASAP7_75t_L g365 ( 
.A(n_304),
.Y(n_365)
);

NAND2xp5_ASAP7_75t_L g366 ( 
.A(n_304),
.B(n_255),
.Y(n_366)
);

NAND2xp5_ASAP7_75t_L g367 ( 
.A(n_307),
.B(n_255),
.Y(n_367)
);

NAND3xp33_ASAP7_75t_L g368 ( 
.A(n_285),
.B(n_255),
.C(n_187),
.Y(n_368)
);

NAND2xp5_ASAP7_75t_L g369 ( 
.A(n_307),
.B(n_260),
.Y(n_369)
);

NAND2xp5_ASAP7_75t_SL g370 ( 
.A(n_285),
.B(n_181),
.Y(n_370)
);

NAND2xp5_ASAP7_75t_L g371 ( 
.A(n_265),
.B(n_235),
.Y(n_371)
);

OAI22xp5_ASAP7_75t_L g372 ( 
.A1(n_314),
.A2(n_248),
.B1(n_262),
.B2(n_277),
.Y(n_372)
);

AOI21xp5_ASAP7_75t_L g373 ( 
.A1(n_321),
.A2(n_328),
.B(n_326),
.Y(n_373)
);

NAND2xp5_ASAP7_75t_L g374 ( 
.A(n_320),
.B(n_268),
.Y(n_374)
);

NAND2xp5_ASAP7_75t_SL g375 ( 
.A(n_363),
.B(n_276),
.Y(n_375)
);

NAND2xp5_ASAP7_75t_L g376 ( 
.A(n_319),
.B(n_265),
.Y(n_376)
);

NOR2xp33_ASAP7_75t_L g377 ( 
.A(n_363),
.B(n_232),
.Y(n_377)
);

AOI21xp5_ASAP7_75t_L g378 ( 
.A1(n_345),
.A2(n_346),
.B(n_335),
.Y(n_378)
);

AOI21xp5_ASAP7_75t_L g379 ( 
.A1(n_323),
.A2(n_312),
.B(n_317),
.Y(n_379)
);

AOI21xp5_ASAP7_75t_L g380 ( 
.A1(n_323),
.A2(n_312),
.B(n_369),
.Y(n_380)
);

AND2x2_ASAP7_75t_L g381 ( 
.A(n_309),
.B(n_232),
.Y(n_381)
);

NAND2xp5_ASAP7_75t_L g382 ( 
.A(n_309),
.B(n_266),
.Y(n_382)
);

NAND2xp5_ASAP7_75t_L g383 ( 
.A(n_331),
.B(n_266),
.Y(n_383)
);

INVx1_ASAP7_75t_L g384 ( 
.A(n_334),
.Y(n_384)
);

NAND2xp5_ASAP7_75t_L g385 ( 
.A(n_331),
.B(n_271),
.Y(n_385)
);

AOI21xp5_ASAP7_75t_L g386 ( 
.A1(n_308),
.A2(n_269),
.B(n_279),
.Y(n_386)
);

NAND2xp5_ASAP7_75t_L g387 ( 
.A(n_314),
.B(n_271),
.Y(n_387)
);

AOI21xp5_ASAP7_75t_L g388 ( 
.A1(n_348),
.A2(n_269),
.B(n_279),
.Y(n_388)
);

NAND2xp5_ASAP7_75t_L g389 ( 
.A(n_338),
.B(n_283),
.Y(n_389)
);

NAND2xp5_ASAP7_75t_L g390 ( 
.A(n_329),
.B(n_283),
.Y(n_390)
);

NAND2xp5_ASAP7_75t_L g391 ( 
.A(n_329),
.B(n_248),
.Y(n_391)
);

NAND2xp5_ASAP7_75t_L g392 ( 
.A(n_333),
.B(n_316),
.Y(n_392)
);

AOI21xp33_ASAP7_75t_L g393 ( 
.A1(n_315),
.A2(n_227),
.B(n_12),
.Y(n_393)
);

OAI21xp5_ASAP7_75t_L g394 ( 
.A1(n_339),
.A2(n_218),
.B(n_235),
.Y(n_394)
);

NAND2xp5_ASAP7_75t_L g395 ( 
.A(n_333),
.B(n_18),
.Y(n_395)
);

INVx1_ASAP7_75t_L g396 ( 
.A(n_347),
.Y(n_396)
);

AND2x2_ASAP7_75t_L g397 ( 
.A(n_355),
.B(n_11),
.Y(n_397)
);

NAND2xp5_ASAP7_75t_SL g398 ( 
.A(n_343),
.B(n_324),
.Y(n_398)
);

AOI21xp5_ASAP7_75t_L g399 ( 
.A1(n_351),
.A2(n_361),
.B(n_360),
.Y(n_399)
);

O2A1O1Ixp33_ASAP7_75t_L g400 ( 
.A1(n_332),
.A2(n_13),
.B(n_14),
.C(n_19),
.Y(n_400)
);

NAND2xp5_ASAP7_75t_L g401 ( 
.A(n_341),
.B(n_20),
.Y(n_401)
);

AOI21xp5_ASAP7_75t_L g402 ( 
.A1(n_366),
.A2(n_89),
.B(n_156),
.Y(n_402)
);

OAI21xp5_ASAP7_75t_L g403 ( 
.A1(n_349),
.A2(n_86),
.B(n_155),
.Y(n_403)
);

AOI21x1_ASAP7_75t_L g404 ( 
.A1(n_350),
.A2(n_85),
.B(n_154),
.Y(n_404)
);

AOI21xp5_ASAP7_75t_L g405 ( 
.A1(n_367),
.A2(n_84),
.B(n_153),
.Y(n_405)
);

BUFx6f_ASAP7_75t_L g406 ( 
.A(n_327),
.Y(n_406)
);

AOI21xp5_ASAP7_75t_L g407 ( 
.A1(n_371),
.A2(n_340),
.B(n_311),
.Y(n_407)
);

AOI21xp5_ASAP7_75t_L g408 ( 
.A1(n_313),
.A2(n_83),
.B(n_151),
.Y(n_408)
);

INVx5_ASAP7_75t_L g409 ( 
.A(n_327),
.Y(n_409)
);

NAND2xp5_ASAP7_75t_SL g410 ( 
.A(n_356),
.B(n_13),
.Y(n_410)
);

BUFx8_ASAP7_75t_SL g411 ( 
.A(n_364),
.Y(n_411)
);

INVx3_ASAP7_75t_L g412 ( 
.A(n_352),
.Y(n_412)
);

INVx11_ASAP7_75t_L g413 ( 
.A(n_364),
.Y(n_413)
);

O2A1O1Ixp5_ASAP7_75t_L g414 ( 
.A1(n_310),
.A2(n_90),
.B(n_27),
.C(n_28),
.Y(n_414)
);

AO21x1_ASAP7_75t_L g415 ( 
.A1(n_330),
.A2(n_14),
.B(n_29),
.Y(n_415)
);

INVx1_ASAP7_75t_L g416 ( 
.A(n_353),
.Y(n_416)
);

INVxp67_ASAP7_75t_SL g417 ( 
.A(n_327),
.Y(n_417)
);

OAI22xp5_ASAP7_75t_L g418 ( 
.A1(n_330),
.A2(n_31),
.B1(n_34),
.B2(n_35),
.Y(n_418)
);

BUFx6f_ASAP7_75t_L g419 ( 
.A(n_327),
.Y(n_419)
);

AOI21xp5_ASAP7_75t_L g420 ( 
.A1(n_322),
.A2(n_36),
.B(n_39),
.Y(n_420)
);

NAND2xp5_ASAP7_75t_L g421 ( 
.A(n_362),
.B(n_41),
.Y(n_421)
);

INVx3_ASAP7_75t_L g422 ( 
.A(n_365),
.Y(n_422)
);

AOI21xp5_ASAP7_75t_L g423 ( 
.A1(n_325),
.A2(n_43),
.B(n_44),
.Y(n_423)
);

NAND2xp5_ASAP7_75t_L g424 ( 
.A(n_336),
.B(n_45),
.Y(n_424)
);

INVx1_ASAP7_75t_L g425 ( 
.A(n_354),
.Y(n_425)
);

O2A1O1Ixp33_ASAP7_75t_L g426 ( 
.A1(n_370),
.A2(n_344),
.B(n_358),
.C(n_359),
.Y(n_426)
);

AOI21xp5_ASAP7_75t_L g427 ( 
.A1(n_342),
.A2(n_48),
.B(n_49),
.Y(n_427)
);

NAND2xp5_ASAP7_75t_L g428 ( 
.A(n_357),
.B(n_50),
.Y(n_428)
);

INVxp67_ASAP7_75t_L g429 ( 
.A(n_370),
.Y(n_429)
);

INVx1_ASAP7_75t_L g430 ( 
.A(n_344),
.Y(n_430)
);

NAND2xp5_ASAP7_75t_SL g431 ( 
.A(n_356),
.B(n_51),
.Y(n_431)
);

INVx3_ASAP7_75t_L g432 ( 
.A(n_337),
.Y(n_432)
);

NOR2xp33_ASAP7_75t_L g433 ( 
.A(n_368),
.B(n_52),
.Y(n_433)
);

NAND2xp5_ASAP7_75t_L g434 ( 
.A(n_337),
.B(n_53),
.Y(n_434)
);

AOI21xp5_ASAP7_75t_L g435 ( 
.A1(n_337),
.A2(n_54),
.B(n_56),
.Y(n_435)
);

AOI21xp33_ASAP7_75t_L g436 ( 
.A1(n_358),
.A2(n_337),
.B(n_318),
.Y(n_436)
);

BUFx6f_ASAP7_75t_L g437 ( 
.A(n_329),
.Y(n_437)
);

O2A1O1Ixp33_ASAP7_75t_L g438 ( 
.A1(n_323),
.A2(n_57),
.B(n_58),
.C(n_60),
.Y(n_438)
);

NAND2xp5_ASAP7_75t_L g439 ( 
.A(n_320),
.B(n_62),
.Y(n_439)
);

NOR2xp33_ASAP7_75t_L g440 ( 
.A(n_377),
.B(n_63),
.Y(n_440)
);

NAND2xp5_ASAP7_75t_L g441 ( 
.A(n_374),
.B(n_65),
.Y(n_441)
);

OAI21x1_ASAP7_75t_L g442 ( 
.A1(n_373),
.A2(n_69),
.B(n_70),
.Y(n_442)
);

NAND2xp5_ASAP7_75t_L g443 ( 
.A(n_387),
.B(n_73),
.Y(n_443)
);

AO21x1_ASAP7_75t_L g444 ( 
.A1(n_372),
.A2(n_74),
.B(n_75),
.Y(n_444)
);

AOI21xp5_ASAP7_75t_L g445 ( 
.A1(n_379),
.A2(n_76),
.B(n_77),
.Y(n_445)
);

OAI21xp5_ASAP7_75t_L g446 ( 
.A1(n_380),
.A2(n_78),
.B(n_80),
.Y(n_446)
);

OAI22xp5_ASAP7_75t_L g447 ( 
.A1(n_429),
.A2(n_81),
.B1(n_82),
.B2(n_91),
.Y(n_447)
);

NOR2xp33_ASAP7_75t_L g448 ( 
.A(n_392),
.B(n_94),
.Y(n_448)
);

INVx1_ASAP7_75t_L g449 ( 
.A(n_384),
.Y(n_449)
);

AOI21xp5_ASAP7_75t_L g450 ( 
.A1(n_378),
.A2(n_96),
.B(n_97),
.Y(n_450)
);

INVx1_ASAP7_75t_L g451 ( 
.A(n_389),
.Y(n_451)
);

AND2x4_ASAP7_75t_L g452 ( 
.A(n_437),
.B(n_98),
.Y(n_452)
);

NAND2xp5_ASAP7_75t_L g453 ( 
.A(n_383),
.B(n_99),
.Y(n_453)
);

NAND2xp5_ASAP7_75t_L g454 ( 
.A(n_385),
.B(n_100),
.Y(n_454)
);

AOI21xp5_ASAP7_75t_L g455 ( 
.A1(n_376),
.A2(n_103),
.B(n_104),
.Y(n_455)
);

OAI21x1_ASAP7_75t_L g456 ( 
.A1(n_399),
.A2(n_107),
.B(n_109),
.Y(n_456)
);

INVx2_ASAP7_75t_L g457 ( 
.A(n_396),
.Y(n_457)
);

O2A1O1Ixp5_ASAP7_75t_L g458 ( 
.A1(n_394),
.A2(n_112),
.B(n_114),
.C(n_115),
.Y(n_458)
);

A2O1A1Ixp33_ASAP7_75t_L g459 ( 
.A1(n_426),
.A2(n_116),
.B(n_118),
.C(n_120),
.Y(n_459)
);

AND2x2_ASAP7_75t_L g460 ( 
.A(n_397),
.B(n_121),
.Y(n_460)
);

OAI21x1_ASAP7_75t_L g461 ( 
.A1(n_407),
.A2(n_158),
.B(n_123),
.Y(n_461)
);

NAND2xp5_ASAP7_75t_SL g462 ( 
.A(n_437),
.B(n_436),
.Y(n_462)
);

NAND2xp5_ASAP7_75t_L g463 ( 
.A(n_382),
.B(n_122),
.Y(n_463)
);

AOI21x1_ASAP7_75t_L g464 ( 
.A1(n_391),
.A2(n_124),
.B(n_126),
.Y(n_464)
);

OAI21x1_ASAP7_75t_L g465 ( 
.A1(n_386),
.A2(n_128),
.B(n_129),
.Y(n_465)
);

AND2x2_ASAP7_75t_L g466 ( 
.A(n_381),
.B(n_130),
.Y(n_466)
);

OAI21xp5_ASAP7_75t_L g467 ( 
.A1(n_439),
.A2(n_131),
.B(n_132),
.Y(n_467)
);

INVx2_ASAP7_75t_L g468 ( 
.A(n_416),
.Y(n_468)
);

OAI21xp5_ASAP7_75t_L g469 ( 
.A1(n_403),
.A2(n_134),
.B(n_135),
.Y(n_469)
);

HB1xp67_ASAP7_75t_L g470 ( 
.A(n_437),
.Y(n_470)
);

OAI21x1_ASAP7_75t_L g471 ( 
.A1(n_388),
.A2(n_401),
.B(n_424),
.Y(n_471)
);

BUFx6f_ASAP7_75t_L g472 ( 
.A(n_406),
.Y(n_472)
);

OAI21xp5_ASAP7_75t_L g473 ( 
.A1(n_430),
.A2(n_141),
.B(n_143),
.Y(n_473)
);

OAI21x1_ASAP7_75t_SL g474 ( 
.A1(n_415),
.A2(n_144),
.B(n_145),
.Y(n_474)
);

AOI21x1_ASAP7_75t_L g475 ( 
.A1(n_390),
.A2(n_395),
.B(n_425),
.Y(n_475)
);

NAND2xp5_ASAP7_75t_L g476 ( 
.A(n_375),
.B(n_147),
.Y(n_476)
);

AOI21xp5_ASAP7_75t_L g477 ( 
.A1(n_409),
.A2(n_148),
.B(n_150),
.Y(n_477)
);

AOI22xp33_ASAP7_75t_L g478 ( 
.A1(n_393),
.A2(n_431),
.B1(n_410),
.B2(n_433),
.Y(n_478)
);

OAI21x1_ASAP7_75t_L g479 ( 
.A1(n_421),
.A2(n_432),
.B(n_434),
.Y(n_479)
);

NAND2xp5_ASAP7_75t_L g480 ( 
.A(n_412),
.B(n_422),
.Y(n_480)
);

NAND2xp5_ASAP7_75t_L g481 ( 
.A(n_412),
.B(n_422),
.Y(n_481)
);

OAI21xp5_ASAP7_75t_L g482 ( 
.A1(n_414),
.A2(n_438),
.B(n_400),
.Y(n_482)
);

OAI21x1_ASAP7_75t_SL g483 ( 
.A1(n_404),
.A2(n_418),
.B(n_428),
.Y(n_483)
);

OAI21x1_ASAP7_75t_L g484 ( 
.A1(n_432),
.A2(n_408),
.B(n_420),
.Y(n_484)
);

AOI21xp5_ASAP7_75t_L g485 ( 
.A1(n_409),
.A2(n_417),
.B(n_419),
.Y(n_485)
);

INVx1_ASAP7_75t_L g486 ( 
.A(n_406),
.Y(n_486)
);

OAI21xp5_ASAP7_75t_L g487 ( 
.A1(n_402),
.A2(n_405),
.B(n_427),
.Y(n_487)
);

INVx2_ASAP7_75t_SL g488 ( 
.A(n_398),
.Y(n_488)
);

AO31x2_ASAP7_75t_L g489 ( 
.A1(n_423),
.A2(n_435),
.A3(n_419),
.B(n_406),
.Y(n_489)
);

AOI21xp5_ASAP7_75t_L g490 ( 
.A1(n_409),
.A2(n_419),
.B(n_413),
.Y(n_490)
);

OAI21xp5_ASAP7_75t_L g491 ( 
.A1(n_411),
.A2(n_373),
.B(n_321),
.Y(n_491)
);

INVx1_ASAP7_75t_SL g492 ( 
.A(n_381),
.Y(n_492)
);

BUFx3_ASAP7_75t_L g493 ( 
.A(n_411),
.Y(n_493)
);

INVx4_ASAP7_75t_L g494 ( 
.A(n_437),
.Y(n_494)
);

BUFx6f_ASAP7_75t_L g495 ( 
.A(n_437),
.Y(n_495)
);

OAI21x1_ASAP7_75t_L g496 ( 
.A1(n_373),
.A2(n_378),
.B(n_399),
.Y(n_496)
);

BUFx3_ASAP7_75t_L g497 ( 
.A(n_495),
.Y(n_497)
);

HB1xp67_ASAP7_75t_L g498 ( 
.A(n_492),
.Y(n_498)
);

INVx1_ASAP7_75t_L g499 ( 
.A(n_449),
.Y(n_499)
);

AO21x1_ASAP7_75t_L g500 ( 
.A1(n_469),
.A2(n_446),
.B(n_482),
.Y(n_500)
);

INVx3_ASAP7_75t_L g501 ( 
.A(n_489),
.Y(n_501)
);

BUFx2_ASAP7_75t_L g502 ( 
.A(n_495),
.Y(n_502)
);

INVx1_ASAP7_75t_L g503 ( 
.A(n_457),
.Y(n_503)
);

OAI21x1_ASAP7_75t_L g504 ( 
.A1(n_496),
.A2(n_479),
.B(n_471),
.Y(n_504)
);

OAI21x1_ASAP7_75t_L g505 ( 
.A1(n_484),
.A2(n_456),
.B(n_442),
.Y(n_505)
);

AO21x2_ASAP7_75t_L g506 ( 
.A1(n_482),
.A2(n_483),
.B(n_444),
.Y(n_506)
);

AND2x2_ASAP7_75t_L g507 ( 
.A(n_451),
.B(n_466),
.Y(n_507)
);

INVx1_ASAP7_75t_L g508 ( 
.A(n_468),
.Y(n_508)
);

OAI21x1_ASAP7_75t_L g509 ( 
.A1(n_461),
.A2(n_475),
.B(n_487),
.Y(n_509)
);

BUFx2_ASAP7_75t_SL g510 ( 
.A(n_495),
.Y(n_510)
);

OA21x2_ASAP7_75t_L g511 ( 
.A1(n_469),
.A2(n_458),
.B(n_487),
.Y(n_511)
);

AO21x2_ASAP7_75t_L g512 ( 
.A1(n_443),
.A2(n_453),
.B(n_454),
.Y(n_512)
);

BUFx2_ASAP7_75t_L g513 ( 
.A(n_470),
.Y(n_513)
);

BUFx3_ASAP7_75t_L g514 ( 
.A(n_452),
.Y(n_514)
);

AND2x2_ASAP7_75t_L g515 ( 
.A(n_492),
.B(n_452),
.Y(n_515)
);

OAI21x1_ASAP7_75t_L g516 ( 
.A1(n_465),
.A2(n_464),
.B(n_445),
.Y(n_516)
);

INVx1_ASAP7_75t_L g517 ( 
.A(n_480),
.Y(n_517)
);

AOI22xp33_ASAP7_75t_SL g518 ( 
.A1(n_440),
.A2(n_488),
.B1(n_460),
.B2(n_448),
.Y(n_518)
);

OA21x2_ASAP7_75t_L g519 ( 
.A1(n_467),
.A2(n_473),
.B(n_459),
.Y(n_519)
);

OAI21x1_ASAP7_75t_L g520 ( 
.A1(n_450),
.A2(n_474),
.B(n_463),
.Y(n_520)
);

OAI21x1_ASAP7_75t_L g521 ( 
.A1(n_485),
.A2(n_467),
.B(n_473),
.Y(n_521)
);

INVx6_ASAP7_75t_L g522 ( 
.A(n_494),
.Y(n_522)
);

OR2x6_ASAP7_75t_L g523 ( 
.A(n_462),
.B(n_494),
.Y(n_523)
);

OAI21x1_ASAP7_75t_L g524 ( 
.A1(n_491),
.A2(n_455),
.B(n_441),
.Y(n_524)
);

INVx1_ASAP7_75t_L g525 ( 
.A(n_481),
.Y(n_525)
);

OAI21x1_ASAP7_75t_L g526 ( 
.A1(n_476),
.A2(n_477),
.B(n_490),
.Y(n_526)
);

OAI21x1_ASAP7_75t_L g527 ( 
.A1(n_486),
.A2(n_447),
.B(n_478),
.Y(n_527)
);

AO21x2_ASAP7_75t_L g528 ( 
.A1(n_489),
.A2(n_472),
.B(n_493),
.Y(n_528)
);

AO21x2_ASAP7_75t_L g529 ( 
.A1(n_472),
.A2(n_482),
.B(n_483),
.Y(n_529)
);

AO21x2_ASAP7_75t_L g530 ( 
.A1(n_472),
.A2(n_482),
.B(n_483),
.Y(n_530)
);

BUFx4f_ASAP7_75t_L g531 ( 
.A(n_495),
.Y(n_531)
);

OA21x2_ASAP7_75t_L g532 ( 
.A1(n_496),
.A2(n_469),
.B(n_482),
.Y(n_532)
);

BUFx2_ASAP7_75t_L g533 ( 
.A(n_495),
.Y(n_533)
);

CKINVDCx5p33_ASAP7_75t_R g534 ( 
.A(n_493),
.Y(n_534)
);

BUFx8_ASAP7_75t_SL g535 ( 
.A(n_493),
.Y(n_535)
);

NOR2xp67_ASAP7_75t_R g536 ( 
.A(n_494),
.B(n_495),
.Y(n_536)
);

OAI21x1_ASAP7_75t_L g537 ( 
.A1(n_496),
.A2(n_479),
.B(n_471),
.Y(n_537)
);

AOI22xp33_ASAP7_75t_L g538 ( 
.A1(n_478),
.A2(n_314),
.B1(n_286),
.B2(n_440),
.Y(n_538)
);

NOR2xp33_ASAP7_75t_L g539 ( 
.A(n_492),
.B(n_324),
.Y(n_539)
);

AND2x2_ASAP7_75t_L g540 ( 
.A(n_451),
.B(n_466),
.Y(n_540)
);

OAI22xp33_ASAP7_75t_L g541 ( 
.A1(n_492),
.A2(n_363),
.B1(n_314),
.B2(n_339),
.Y(n_541)
);

AO21x2_ASAP7_75t_L g542 ( 
.A1(n_482),
.A2(n_483),
.B(n_444),
.Y(n_542)
);

NOR2xp67_ASAP7_75t_L g543 ( 
.A(n_488),
.B(n_343),
.Y(n_543)
);

INVx1_ASAP7_75t_L g544 ( 
.A(n_449),
.Y(n_544)
);

OAI21x1_ASAP7_75t_L g545 ( 
.A1(n_496),
.A2(n_479),
.B(n_471),
.Y(n_545)
);

AO21x2_ASAP7_75t_L g546 ( 
.A1(n_482),
.A2(n_483),
.B(n_444),
.Y(n_546)
);

INVx1_ASAP7_75t_L g547 ( 
.A(n_499),
.Y(n_547)
);

BUFx2_ASAP7_75t_L g548 ( 
.A(n_498),
.Y(n_548)
);

AOI22xp33_ASAP7_75t_L g549 ( 
.A1(n_538),
.A2(n_500),
.B1(n_518),
.B2(n_515),
.Y(n_549)
);

HB1xp67_ASAP7_75t_L g550 ( 
.A(n_515),
.Y(n_550)
);

INVx3_ASAP7_75t_L g551 ( 
.A(n_529),
.Y(n_551)
);

INVx1_ASAP7_75t_L g552 ( 
.A(n_544),
.Y(n_552)
);

INVx1_ASAP7_75t_L g553 ( 
.A(n_517),
.Y(n_553)
);

INVx1_ASAP7_75t_L g554 ( 
.A(n_525),
.Y(n_554)
);

AOI21x1_ASAP7_75t_L g555 ( 
.A1(n_509),
.A2(n_500),
.B(n_505),
.Y(n_555)
);

AOI22xp33_ASAP7_75t_L g556 ( 
.A1(n_541),
.A2(n_514),
.B1(n_507),
.B2(n_540),
.Y(n_556)
);

INVx1_ASAP7_75t_L g557 ( 
.A(n_503),
.Y(n_557)
);

BUFx2_ASAP7_75t_L g558 ( 
.A(n_513),
.Y(n_558)
);

OR2x2_ASAP7_75t_L g559 ( 
.A(n_507),
.B(n_540),
.Y(n_559)
);

INVx1_ASAP7_75t_L g560 ( 
.A(n_508),
.Y(n_560)
);

INVx4_ASAP7_75t_L g561 ( 
.A(n_531),
.Y(n_561)
);

INVx1_ASAP7_75t_L g562 ( 
.A(n_514),
.Y(n_562)
);

INVx1_ASAP7_75t_L g563 ( 
.A(n_523),
.Y(n_563)
);

BUFx2_ASAP7_75t_L g564 ( 
.A(n_497),
.Y(n_564)
);

INVxp67_ASAP7_75t_L g565 ( 
.A(n_539),
.Y(n_565)
);

INVx1_ASAP7_75t_L g566 ( 
.A(n_523),
.Y(n_566)
);

INVx1_ASAP7_75t_L g567 ( 
.A(n_523),
.Y(n_567)
);

BUFx2_ASAP7_75t_L g568 ( 
.A(n_497),
.Y(n_568)
);

AND2x2_ASAP7_75t_L g569 ( 
.A(n_528),
.B(n_523),
.Y(n_569)
);

OR2x2_ASAP7_75t_L g570 ( 
.A(n_528),
.B(n_529),
.Y(n_570)
);

AOI21x1_ASAP7_75t_L g571 ( 
.A1(n_509),
.A2(n_545),
.B(n_504),
.Y(n_571)
);

INVx2_ASAP7_75t_L g572 ( 
.A(n_501),
.Y(n_572)
);

AOI22xp33_ASAP7_75t_L g573 ( 
.A1(n_519),
.A2(n_528),
.B1(n_532),
.B2(n_506),
.Y(n_573)
);

AO21x2_ASAP7_75t_L g574 ( 
.A1(n_537),
.A2(n_545),
.B(n_546),
.Y(n_574)
);

INVx1_ASAP7_75t_L g575 ( 
.A(n_529),
.Y(n_575)
);

INVx2_ASAP7_75t_L g576 ( 
.A(n_530),
.Y(n_576)
);

HB1xp67_ASAP7_75t_L g577 ( 
.A(n_502),
.Y(n_577)
);

AOI21x1_ASAP7_75t_L g578 ( 
.A1(n_511),
.A2(n_516),
.B(n_520),
.Y(n_578)
);

INVx2_ASAP7_75t_L g579 ( 
.A(n_530),
.Y(n_579)
);

CKINVDCx5p33_ASAP7_75t_R g580 ( 
.A(n_535),
.Y(n_580)
);

INVx2_ASAP7_75t_L g581 ( 
.A(n_530),
.Y(n_581)
);

INVx2_ASAP7_75t_L g582 ( 
.A(n_527),
.Y(n_582)
);

INVx1_ASAP7_75t_L g583 ( 
.A(n_531),
.Y(n_583)
);

OAI21xp5_ASAP7_75t_L g584 ( 
.A1(n_527),
.A2(n_521),
.B(n_524),
.Y(n_584)
);

CKINVDCx9p33_ASAP7_75t_R g585 ( 
.A(n_533),
.Y(n_585)
);

AND2x2_ASAP7_75t_L g586 ( 
.A(n_559),
.B(n_506),
.Y(n_586)
);

AND2x2_ASAP7_75t_L g587 ( 
.A(n_559),
.B(n_506),
.Y(n_587)
);

INVx5_ASAP7_75t_L g588 ( 
.A(n_561),
.Y(n_588)
);

INVx4_ASAP7_75t_L g589 ( 
.A(n_561),
.Y(n_589)
);

AND2x2_ASAP7_75t_L g590 ( 
.A(n_553),
.B(n_546),
.Y(n_590)
);

HB1xp67_ASAP7_75t_L g591 ( 
.A(n_558),
.Y(n_591)
);

AOI222xp33_ASAP7_75t_L g592 ( 
.A1(n_565),
.A2(n_543),
.B1(n_521),
.B2(n_534),
.C1(n_531),
.C2(n_536),
.Y(n_592)
);

OR2x2_ASAP7_75t_L g593 ( 
.A(n_570),
.B(n_532),
.Y(n_593)
);

AND2x2_ASAP7_75t_L g594 ( 
.A(n_553),
.B(n_546),
.Y(n_594)
);

AND2x2_ASAP7_75t_L g595 ( 
.A(n_554),
.B(n_542),
.Y(n_595)
);

AND2x2_ASAP7_75t_L g596 ( 
.A(n_554),
.B(n_542),
.Y(n_596)
);

INVx2_ASAP7_75t_L g597 ( 
.A(n_547),
.Y(n_597)
);

INVx2_ASAP7_75t_L g598 ( 
.A(n_547),
.Y(n_598)
);

HB1xp67_ASAP7_75t_L g599 ( 
.A(n_558),
.Y(n_599)
);

BUFx3_ASAP7_75t_L g600 ( 
.A(n_564),
.Y(n_600)
);

AO31x2_ASAP7_75t_L g601 ( 
.A1(n_582),
.A2(n_575),
.A3(n_581),
.B(n_576),
.Y(n_601)
);

AOI22xp33_ASAP7_75t_L g602 ( 
.A1(n_549),
.A2(n_519),
.B1(n_532),
.B2(n_542),
.Y(n_602)
);

INVx3_ASAP7_75t_L g603 ( 
.A(n_561),
.Y(n_603)
);

INVx1_ASAP7_75t_L g604 ( 
.A(n_575),
.Y(n_604)
);

INVx2_ASAP7_75t_L g605 ( 
.A(n_552),
.Y(n_605)
);

AND2x2_ASAP7_75t_L g606 ( 
.A(n_550),
.B(n_519),
.Y(n_606)
);

INVx1_ASAP7_75t_L g607 ( 
.A(n_576),
.Y(n_607)
);

BUFx2_ASAP7_75t_L g608 ( 
.A(n_548),
.Y(n_608)
);

INVx2_ASAP7_75t_SL g609 ( 
.A(n_564),
.Y(n_609)
);

INVx1_ASAP7_75t_L g610 ( 
.A(n_579),
.Y(n_610)
);

INVx2_ASAP7_75t_L g611 ( 
.A(n_557),
.Y(n_611)
);

INVx2_ASAP7_75t_L g612 ( 
.A(n_557),
.Y(n_612)
);

INVx2_ASAP7_75t_L g613 ( 
.A(n_560),
.Y(n_613)
);

INVx1_ASAP7_75t_L g614 ( 
.A(n_548),
.Y(n_614)
);

OR2x2_ASAP7_75t_L g615 ( 
.A(n_570),
.B(n_511),
.Y(n_615)
);

BUFx2_ASAP7_75t_L g616 ( 
.A(n_563),
.Y(n_616)
);

BUFx3_ASAP7_75t_L g617 ( 
.A(n_568),
.Y(n_617)
);

INVxp67_ASAP7_75t_SL g618 ( 
.A(n_577),
.Y(n_618)
);

AND2x2_ASAP7_75t_L g619 ( 
.A(n_556),
.B(n_511),
.Y(n_619)
);

NOR2xp33_ASAP7_75t_L g620 ( 
.A(n_562),
.B(n_534),
.Y(n_620)
);

AND2x2_ASAP7_75t_L g621 ( 
.A(n_569),
.B(n_526),
.Y(n_621)
);

BUFx3_ASAP7_75t_L g622 ( 
.A(n_568),
.Y(n_622)
);

OR2x2_ASAP7_75t_SL g623 ( 
.A(n_566),
.B(n_522),
.Y(n_623)
);

HB1xp67_ASAP7_75t_L g624 ( 
.A(n_567),
.Y(n_624)
);

INVx2_ASAP7_75t_L g625 ( 
.A(n_597),
.Y(n_625)
);

OAI22xp5_ASAP7_75t_L g626 ( 
.A1(n_623),
.A2(n_583),
.B1(n_569),
.B2(n_522),
.Y(n_626)
);

INVx1_ASAP7_75t_L g627 ( 
.A(n_604),
.Y(n_627)
);

INVx1_ASAP7_75t_L g628 ( 
.A(n_604),
.Y(n_628)
);

NAND2xp5_ASAP7_75t_SL g629 ( 
.A(n_588),
.B(n_551),
.Y(n_629)
);

INVx3_ASAP7_75t_L g630 ( 
.A(n_601),
.Y(n_630)
);

INVx1_ASAP7_75t_L g631 ( 
.A(n_601),
.Y(n_631)
);

AOI22xp33_ASAP7_75t_L g632 ( 
.A1(n_592),
.A2(n_582),
.B1(n_512),
.B2(n_584),
.Y(n_632)
);

AND2x2_ASAP7_75t_L g633 ( 
.A(n_586),
.B(n_573),
.Y(n_633)
);

NAND2xp5_ASAP7_75t_L g634 ( 
.A(n_591),
.B(n_599),
.Y(n_634)
);

AND2x2_ASAP7_75t_L g635 ( 
.A(n_586),
.B(n_551),
.Y(n_635)
);

BUFx2_ASAP7_75t_SL g636 ( 
.A(n_609),
.Y(n_636)
);

AND2x2_ASAP7_75t_L g637 ( 
.A(n_587),
.B(n_551),
.Y(n_637)
);

BUFx3_ASAP7_75t_L g638 ( 
.A(n_600),
.Y(n_638)
);

AND2x2_ASAP7_75t_L g639 ( 
.A(n_587),
.B(n_572),
.Y(n_639)
);

BUFx3_ASAP7_75t_L g640 ( 
.A(n_600),
.Y(n_640)
);

AND2x2_ASAP7_75t_L g641 ( 
.A(n_606),
.B(n_572),
.Y(n_641)
);

CKINVDCx20_ASAP7_75t_R g642 ( 
.A(n_623),
.Y(n_642)
);

AOI22xp33_ASAP7_75t_L g643 ( 
.A1(n_608),
.A2(n_512),
.B1(n_524),
.B2(n_522),
.Y(n_643)
);

INVx2_ASAP7_75t_L g644 ( 
.A(n_598),
.Y(n_644)
);

HB1xp67_ASAP7_75t_L g645 ( 
.A(n_608),
.Y(n_645)
);

AND2x4_ASAP7_75t_L g646 ( 
.A(n_598),
.B(n_555),
.Y(n_646)
);

AND2x2_ASAP7_75t_L g647 ( 
.A(n_590),
.B(n_574),
.Y(n_647)
);

AND2x2_ASAP7_75t_L g648 ( 
.A(n_594),
.B(n_574),
.Y(n_648)
);

INVxp67_ASAP7_75t_SL g649 ( 
.A(n_618),
.Y(n_649)
);

NAND2xp5_ASAP7_75t_L g650 ( 
.A(n_614),
.B(n_510),
.Y(n_650)
);

INVx1_ASAP7_75t_L g651 ( 
.A(n_607),
.Y(n_651)
);

BUFx2_ASAP7_75t_L g652 ( 
.A(n_616),
.Y(n_652)
);

INVx1_ASAP7_75t_L g653 ( 
.A(n_607),
.Y(n_653)
);

OR2x2_ASAP7_75t_L g654 ( 
.A(n_593),
.B(n_574),
.Y(n_654)
);

BUFx2_ASAP7_75t_L g655 ( 
.A(n_616),
.Y(n_655)
);

AND2x2_ASAP7_75t_L g656 ( 
.A(n_595),
.B(n_578),
.Y(n_656)
);

INVx4_ASAP7_75t_L g657 ( 
.A(n_588),
.Y(n_657)
);

AND2x2_ASAP7_75t_L g658 ( 
.A(n_595),
.B(n_571),
.Y(n_658)
);

AND2x2_ASAP7_75t_L g659 ( 
.A(n_596),
.B(n_619),
.Y(n_659)
);

INVx1_ASAP7_75t_L g660 ( 
.A(n_627),
.Y(n_660)
);

INVx1_ASAP7_75t_L g661 ( 
.A(n_627),
.Y(n_661)
);

INVx2_ASAP7_75t_L g662 ( 
.A(n_628),
.Y(n_662)
);

HB1xp67_ASAP7_75t_L g663 ( 
.A(n_652),
.Y(n_663)
);

NAND2xp5_ASAP7_75t_L g664 ( 
.A(n_649),
.B(n_624),
.Y(n_664)
);

INVx1_ASAP7_75t_L g665 ( 
.A(n_628),
.Y(n_665)
);

INVx1_ASAP7_75t_L g666 ( 
.A(n_651),
.Y(n_666)
);

NAND2xp5_ASAP7_75t_L g667 ( 
.A(n_634),
.B(n_605),
.Y(n_667)
);

AND2x4_ASAP7_75t_L g668 ( 
.A(n_646),
.B(n_621),
.Y(n_668)
);

AND2x2_ASAP7_75t_L g669 ( 
.A(n_659),
.B(n_621),
.Y(n_669)
);

NAND2xp5_ASAP7_75t_L g670 ( 
.A(n_645),
.B(n_605),
.Y(n_670)
);

AOI22xp33_ASAP7_75t_L g671 ( 
.A1(n_642),
.A2(n_619),
.B1(n_602),
.B2(n_613),
.Y(n_671)
);

INVx1_ASAP7_75t_L g672 ( 
.A(n_651),
.Y(n_672)
);

AND2x2_ASAP7_75t_L g673 ( 
.A(n_659),
.B(n_593),
.Y(n_673)
);

NAND2xp5_ASAP7_75t_L g674 ( 
.A(n_639),
.B(n_613),
.Y(n_674)
);

AND2x2_ASAP7_75t_L g675 ( 
.A(n_633),
.B(n_596),
.Y(n_675)
);

HB1xp67_ASAP7_75t_L g676 ( 
.A(n_652),
.Y(n_676)
);

AND2x2_ASAP7_75t_L g677 ( 
.A(n_633),
.B(n_635),
.Y(n_677)
);

INVx3_ASAP7_75t_L g678 ( 
.A(n_646),
.Y(n_678)
);

INVx1_ASAP7_75t_L g679 ( 
.A(n_653),
.Y(n_679)
);

NAND2xp5_ASAP7_75t_L g680 ( 
.A(n_639),
.B(n_612),
.Y(n_680)
);

AND2x4_ASAP7_75t_L g681 ( 
.A(n_646),
.B(n_610),
.Y(n_681)
);

INVx1_ASAP7_75t_L g682 ( 
.A(n_655),
.Y(n_682)
);

NAND2xp5_ASAP7_75t_L g683 ( 
.A(n_641),
.B(n_612),
.Y(n_683)
);

INVx1_ASAP7_75t_L g684 ( 
.A(n_655),
.Y(n_684)
);

AND2x2_ASAP7_75t_L g685 ( 
.A(n_635),
.B(n_637),
.Y(n_685)
);

HB1xp67_ASAP7_75t_L g686 ( 
.A(n_638),
.Y(n_686)
);

NAND2xp5_ASAP7_75t_L g687 ( 
.A(n_641),
.B(n_611),
.Y(n_687)
);

INVx1_ASAP7_75t_L g688 ( 
.A(n_625),
.Y(n_688)
);

AND2x2_ASAP7_75t_L g689 ( 
.A(n_637),
.B(n_615),
.Y(n_689)
);

INVx1_ASAP7_75t_L g690 ( 
.A(n_644),
.Y(n_690)
);

AND3x2_ASAP7_75t_L g691 ( 
.A(n_686),
.B(n_611),
.C(n_620),
.Y(n_691)
);

AND2x2_ASAP7_75t_L g692 ( 
.A(n_677),
.B(n_647),
.Y(n_692)
);

INVx1_ASAP7_75t_L g693 ( 
.A(n_662),
.Y(n_693)
);

OR2x2_ASAP7_75t_L g694 ( 
.A(n_677),
.B(n_654),
.Y(n_694)
);

AND2x2_ASAP7_75t_L g695 ( 
.A(n_685),
.B(n_648),
.Y(n_695)
);

AND2x2_ASAP7_75t_L g696 ( 
.A(n_685),
.B(n_648),
.Y(n_696)
);

AND2x2_ASAP7_75t_L g697 ( 
.A(n_669),
.B(n_647),
.Y(n_697)
);

INVx1_ASAP7_75t_L g698 ( 
.A(n_662),
.Y(n_698)
);

NAND2xp5_ASAP7_75t_L g699 ( 
.A(n_667),
.B(n_658),
.Y(n_699)
);

NAND2xp5_ASAP7_75t_L g700 ( 
.A(n_664),
.B(n_658),
.Y(n_700)
);

AND2x4_ASAP7_75t_L g701 ( 
.A(n_678),
.B(n_630),
.Y(n_701)
);

INVx1_ASAP7_75t_L g702 ( 
.A(n_660),
.Y(n_702)
);

AND2x2_ASAP7_75t_L g703 ( 
.A(n_669),
.B(n_640),
.Y(n_703)
);

AND2x2_ASAP7_75t_L g704 ( 
.A(n_673),
.B(n_656),
.Y(n_704)
);

AND2x2_ASAP7_75t_L g705 ( 
.A(n_673),
.B(n_640),
.Y(n_705)
);

OR2x2_ASAP7_75t_L g706 ( 
.A(n_689),
.B(n_654),
.Y(n_706)
);

INVx1_ASAP7_75t_L g707 ( 
.A(n_661),
.Y(n_707)
);

AND2x2_ASAP7_75t_L g708 ( 
.A(n_675),
.B(n_689),
.Y(n_708)
);

OR2x2_ASAP7_75t_L g709 ( 
.A(n_675),
.B(n_656),
.Y(n_709)
);

AND2x2_ASAP7_75t_L g710 ( 
.A(n_668),
.B(n_678),
.Y(n_710)
);

NAND2xp5_ASAP7_75t_SL g711 ( 
.A(n_700),
.B(n_638),
.Y(n_711)
);

NAND3xp33_ASAP7_75t_SL g712 ( 
.A(n_691),
.B(n_671),
.C(n_632),
.Y(n_712)
);

OA222x2_ASAP7_75t_L g713 ( 
.A1(n_691),
.A2(n_678),
.B1(n_682),
.B2(n_684),
.C1(n_630),
.C2(n_631),
.Y(n_713)
);

INVxp67_ASAP7_75t_L g714 ( 
.A(n_702),
.Y(n_714)
);

AOI22xp33_ASAP7_75t_L g715 ( 
.A1(n_705),
.A2(n_671),
.B1(n_626),
.B2(n_668),
.Y(n_715)
);

AO21x1_ASAP7_75t_L g716 ( 
.A1(n_707),
.A2(n_698),
.B(n_693),
.Y(n_716)
);

OAI22xp5_ASAP7_75t_L g717 ( 
.A1(n_699),
.A2(n_709),
.B1(n_694),
.B2(n_706),
.Y(n_717)
);

OAI22xp5_ASAP7_75t_L g718 ( 
.A1(n_703),
.A2(n_603),
.B1(n_668),
.B2(n_663),
.Y(n_718)
);

NAND2xp5_ASAP7_75t_L g719 ( 
.A(n_708),
.B(n_676),
.Y(n_719)
);

INVx1_ASAP7_75t_L g720 ( 
.A(n_704),
.Y(n_720)
);

AND2x2_ASAP7_75t_L g721 ( 
.A(n_692),
.B(n_681),
.Y(n_721)
);

AOI21xp5_ASAP7_75t_L g722 ( 
.A1(n_701),
.A2(n_629),
.B(n_643),
.Y(n_722)
);

INVx2_ASAP7_75t_L g723 ( 
.A(n_710),
.Y(n_723)
);

INVx1_ASAP7_75t_L g724 ( 
.A(n_704),
.Y(n_724)
);

OAI21xp33_ASAP7_75t_L g725 ( 
.A1(n_712),
.A2(n_674),
.B(n_670),
.Y(n_725)
);

INVx1_ASAP7_75t_L g726 ( 
.A(n_714),
.Y(n_726)
);

NAND2xp5_ASAP7_75t_L g727 ( 
.A(n_717),
.B(n_695),
.Y(n_727)
);

O2A1O1Ixp33_ASAP7_75t_L g728 ( 
.A1(n_712),
.A2(n_650),
.B(n_609),
.C(n_680),
.Y(n_728)
);

AOI22x1_ASAP7_75t_L g729 ( 
.A1(n_722),
.A2(n_580),
.B1(n_636),
.B2(n_710),
.Y(n_729)
);

AOI22xp5_ASAP7_75t_L g730 ( 
.A1(n_711),
.A2(n_701),
.B1(n_603),
.B2(n_589),
.Y(n_730)
);

OAI221xp5_ASAP7_75t_L g731 ( 
.A1(n_715),
.A2(n_683),
.B1(n_687),
.B2(n_665),
.C(n_672),
.Y(n_731)
);

BUFx3_ASAP7_75t_L g732 ( 
.A(n_726),
.Y(n_732)
);

AOI21xp5_ASAP7_75t_L g733 ( 
.A1(n_725),
.A2(n_716),
.B(n_714),
.Y(n_733)
);

AOI211xp5_ASAP7_75t_SL g734 ( 
.A1(n_731),
.A2(n_718),
.B(n_713),
.C(n_719),
.Y(n_734)
);

AOI21xp33_ASAP7_75t_SL g735 ( 
.A1(n_729),
.A2(n_728),
.B(n_727),
.Y(n_735)
);

OAI21xp5_ASAP7_75t_SL g736 ( 
.A1(n_730),
.A2(n_724),
.B(n_720),
.Y(n_736)
);

AOI22xp5_ASAP7_75t_L g737 ( 
.A1(n_725),
.A2(n_701),
.B1(n_723),
.B2(n_681),
.Y(n_737)
);

NAND3xp33_ASAP7_75t_SL g738 ( 
.A(n_734),
.B(n_580),
.C(n_721),
.Y(n_738)
);

NAND2xp5_ASAP7_75t_L g739 ( 
.A(n_732),
.B(n_696),
.Y(n_739)
);

AOI21xp5_ASAP7_75t_L g740 ( 
.A1(n_733),
.A2(n_666),
.B(n_679),
.Y(n_740)
);

NAND3xp33_ASAP7_75t_L g741 ( 
.A(n_735),
.B(n_688),
.C(n_690),
.Y(n_741)
);

INVx1_ASAP7_75t_L g742 ( 
.A(n_737),
.Y(n_742)
);

NOR2x1_ASAP7_75t_L g743 ( 
.A(n_741),
.B(n_736),
.Y(n_743)
);

NOR2xp33_ASAP7_75t_L g744 ( 
.A(n_738),
.B(n_535),
.Y(n_744)
);

INVx1_ASAP7_75t_L g745 ( 
.A(n_739),
.Y(n_745)
);

NAND3xp33_ASAP7_75t_L g746 ( 
.A(n_743),
.B(n_740),
.C(n_742),
.Y(n_746)
);

NAND4xp25_ASAP7_75t_L g747 ( 
.A(n_744),
.B(n_622),
.C(n_617),
.D(n_589),
.Y(n_747)
);

INVx1_ASAP7_75t_L g748 ( 
.A(n_745),
.Y(n_748)
);

INVx2_ASAP7_75t_L g749 ( 
.A(n_748),
.Y(n_749)
);

NAND2x1p5_ASAP7_75t_L g750 ( 
.A(n_747),
.B(n_588),
.Y(n_750)
);

INVx1_ASAP7_75t_L g751 ( 
.A(n_746),
.Y(n_751)
);

INVx1_ASAP7_75t_L g752 ( 
.A(n_748),
.Y(n_752)
);

AOI22xp5_ASAP7_75t_L g753 ( 
.A1(n_746),
.A2(n_636),
.B1(n_681),
.B2(n_589),
.Y(n_753)
);

INVxp67_ASAP7_75t_L g754 ( 
.A(n_746),
.Y(n_754)
);

INVx2_ASAP7_75t_L g755 ( 
.A(n_750),
.Y(n_755)
);

OAI22xp5_ASAP7_75t_SL g756 ( 
.A1(n_754),
.A2(n_588),
.B1(n_585),
.B2(n_657),
.Y(n_756)
);

OR2x2_ASAP7_75t_L g757 ( 
.A(n_751),
.B(n_749),
.Y(n_757)
);

XNOR2x1_ASAP7_75t_L g758 ( 
.A(n_752),
.B(n_603),
.Y(n_758)
);

INVx5_ASAP7_75t_L g759 ( 
.A(n_753),
.Y(n_759)
);

OAI22xp5_ASAP7_75t_L g760 ( 
.A1(n_754),
.A2(n_697),
.B1(n_696),
.B2(n_695),
.Y(n_760)
);

INVx2_ASAP7_75t_L g761 ( 
.A(n_757),
.Y(n_761)
);

NAND2xp5_ASAP7_75t_L g762 ( 
.A(n_758),
.B(n_697),
.Y(n_762)
);

INVx1_ASAP7_75t_L g763 ( 
.A(n_759),
.Y(n_763)
);

XNOR2x1_ASAP7_75t_L g764 ( 
.A(n_755),
.B(n_617),
.Y(n_764)
);

INVx1_ASAP7_75t_L g765 ( 
.A(n_761),
.Y(n_765)
);

INVx1_ASAP7_75t_L g766 ( 
.A(n_763),
.Y(n_766)
);

AND2x4_ASAP7_75t_L g767 ( 
.A(n_762),
.B(n_756),
.Y(n_767)
);

INVx1_ASAP7_75t_L g768 ( 
.A(n_766),
.Y(n_768)
);

INVx1_ASAP7_75t_L g769 ( 
.A(n_765),
.Y(n_769)
);

HB1xp67_ASAP7_75t_L g770 ( 
.A(n_767),
.Y(n_770)
);

OA22x2_ASAP7_75t_L g771 ( 
.A1(n_770),
.A2(n_764),
.B1(n_760),
.B2(n_657),
.Y(n_771)
);

INVx2_ASAP7_75t_L g772 ( 
.A(n_768),
.Y(n_772)
);

AND2x2_ASAP7_75t_L g773 ( 
.A(n_772),
.B(n_769),
.Y(n_773)
);

INVx1_ASAP7_75t_L g774 ( 
.A(n_773),
.Y(n_774)
);

NAND2xp5_ASAP7_75t_L g775 ( 
.A(n_774),
.B(n_771),
.Y(n_775)
);

AOI22xp33_ASAP7_75t_L g776 ( 
.A1(n_775),
.A2(n_622),
.B1(n_588),
.B2(n_522),
.Y(n_776)
);


endmodule