module real_aes_6236_n_102 (n_17, n_28, n_76, n_56, n_34, n_98, n_90, n_82, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_83, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_91, n_100, n_43, n_96, n_54, n_35, n_42, n_99, n_15, n_9, n_23, n_72, n_95, n_44, n_7, n_4, n_80, n_6, n_12, n_68, n_79, n_69, n_46, n_59, n_25, n_73, n_77, n_81, n_48, n_37, n_97, n_70, n_50, n_89, n_26, n_86, n_93, n_13, n_24, n_2, n_55, n_62, n_84, n_67, n_92, n_33, n_88, n_14, n_11, n_85, n_16, n_94, n_39, n_5, n_45, n_60, n_38, n_87, n_0, n_78, n_101, n_63, n_1, n_53, n_36, n_102);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_98;
input n_90;
input n_82;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_83;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_91;
input n_100;
input n_43;
input n_96;
input n_54;
input n_35;
input n_42;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_95;
input n_44;
input n_7;
input n_4;
input n_80;
input n_6;
input n_12;
input n_68;
input n_79;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_81;
input n_48;
input n_37;
input n_97;
input n_70;
input n_50;
input n_89;
input n_26;
input n_86;
input n_93;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_84;
input n_67;
input n_92;
input n_33;
input n_88;
input n_14;
input n_11;
input n_85;
input n_16;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_87;
input n_0;
input n_78;
input n_101;
input n_63;
input n_1;
input n_53;
input n_36;
output n_102;
wire n_480;
wire n_113;
wire n_476;
wire n_758;
wire n_599;
wire n_187;
wire n_436;
wire n_684;
wire n_257;
wire n_390;
wire n_185;
wire n_285;
wire n_624;
wire n_618;
wire n_522;
wire n_485;
wire n_222;
wire n_750;
wire n_631;
wire n_503;
wire n_287;
wire n_357;
wire n_635;
wire n_386;
wire n_673;
wire n_518;
wire n_254;
wire n_207;
wire n_665;
wire n_667;
wire n_577;
wire n_580;
wire n_469;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_759;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_718;
wire n_318;
wire n_355;
wire n_239;
wire n_669;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_761;
wire n_742;
wire n_112;
wire n_319;
wire n_364;
wire n_421;
wire n_555;
wire n_329;
wire n_766;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_169;
wire n_242;
wire n_376;
wire n_549;
wire n_571;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_752;
wire n_448;
wire n_556;
wire n_545;
wire n_341;
wire n_593;
wire n_232;
wire n_460;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_537;
wire n_320;
wire n_551;
wire n_666;
wire n_560;
wire n_260;
wire n_660;
wire n_594;
wire n_186;
wire n_767;
wire n_138;
wire n_696;
wire n_704;
wire n_379;
wire n_374;
wire n_453;
wire n_647;
wire n_235;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_161;
wire n_763;
wire n_189;
wire n_271;
wire n_489;
wire n_548;
wire n_427;
wire n_678;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_519;
wire n_564;
wire n_638;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_512;
wire n_395;
wire n_332;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_116;
wire n_625;
wire n_289;
wire n_462;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_716;
wire n_213;
wire n_356;
wire n_478;
wire n_584;
wire n_408;
wire n_553;
wire n_184;
wire n_372;
wire n_528;
wire n_578;
wire n_202;
wire n_495;
wire n_370;
wire n_384;
wire n_744;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_467;
wire n_327;
wire n_106;
wire n_559;
wire n_466;
wire n_636;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_726;
wire n_517;
wire n_683;
wire n_174;
wire n_570;
wire n_675;
wire n_530;
wire n_104;
wire n_535;
wire n_732;
wire n_211;
wire n_281;
wire n_496;
wire n_693;
wire n_173;
wire n_468;
wire n_234;
wire n_746;
wire n_284;
wire n_153;
wire n_316;
wire n_532;
wire n_656;
wire n_755;
wire n_178;
wire n_409;
wire n_748;
wire n_523;
wire n_298;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_297;
wire n_383;
wire n_529;
wire n_119;
wire n_310;
wire n_455;
wire n_504;
wire n_725;
wire n_164;
wire n_671;
wire n_231;
wire n_547;
wire n_659;
wire n_682;
wire n_634;
wire n_454;
wire n_122;
wire n_443;
wire n_565;
wire n_760;
wire n_608;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_267;
wire n_218;
wire n_737;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_745;
wire n_722;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_331;
wire n_182;
wire n_417;
wire n_363;
wire n_754;
wire n_449;
wire n_607;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_142;
wire n_561;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_655;
wire n_654;
wire n_505;
wire n_434;
wire n_502;
wire n_527;
wire n_769;
wire n_600;
wire n_731;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_733;
wire n_552;
wire n_402;
wire n_602;
wire n_617;
wire n_171;
wire n_658;
wire n_676;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_146;
wire n_432;
wire n_226;
wire n_255;
wire n_286;
wire n_416;
wire n_410;
wire n_120;
wire n_751;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_695;
wire n_685;
wire n_165;
wire n_361;
wire n_632;
wire n_246;
wire n_176;
wire n_768;
wire n_412;
wire n_163;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_501;
wire n_488;
wire n_251;
wire n_642;
wire n_613;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_702;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_734;
wire n_110;
wire n_392;
wire n_562;
wire n_150;
wire n_288;
wire n_147;
wire n_404;
wire n_598;
wire n_713;
wire n_728;
wire n_735;
wire n_756;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_569;
wire n_563;
wire n_188;
wire n_269;
wire n_430;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_193;
wire n_397;
wire n_293;
wire n_162;
wire n_749;
wire n_358;
wire n_275;
wire n_214;
wire n_385;
wire n_649;
wire n_663;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_707;
wire n_622;
wire n_470;
wire n_133;
wire n_494;
wire n_711;
wire n_377;
wire n_273;
wire n_723;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_265;
wire n_354;
wire n_720;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_730;
wire n_643;
wire n_747;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_148;
wire n_498;
wire n_481;
wire n_691;
wire n_765;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_233;
wire n_487;
wire n_290;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_155;
wire n_243;
wire n_692;
wire n_544;
wire n_268;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_738;
wire n_701;
wire n_309;
wire n_344;
wire n_107;
wire n_229;
wire n_482;
wire n_520;
wire n_633;
wire n_679;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_262;
wire n_630;
wire n_689;
wire n_715;
wire n_134;
wire n_420;
wire n_336;
wire n_349;
wire n_612;
wire n_195;
wire n_438;
wire n_764;
wire n_300;
wire n_753;
wire n_252;
wire n_314;
wire n_283;
wire n_741;
wire n_249;
wire n_623;
wire n_446;
wire n_721;
wire n_221;
wire n_681;
wire n_156;
wire n_359;
wire n_456;
wire n_717;
wire n_312;
wire n_183;
wire n_266;
wire n_712;
wire n_205;
wire n_433;
wire n_335;
wire n_177;
wire n_516;
wire n_313;
wire n_627;
wire n_739;
wire n_140;
wire n_418;
wire n_521;
wire n_422;
wire n_524;
wire n_219;
wire n_705;
wire n_180;
wire n_762;
wire n_212;
wire n_210;
wire n_325;
wire n_575;
wire n_338;
wire n_479;
wire n_442;
wire n_698;
wire n_371;
wire n_740;
wire n_166;
wire n_103;
wire n_541;
wire n_224;
wire n_546;
wire n_151;
wire n_587;
wire n_639;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_724;
wire n_440;
wire n_525;
wire n_674;
wire n_644;
wire n_152;
wire n_198;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_414;
wire n_757;
wire n_123;
wire n_279;
wire n_686;
wire n_543;
wire n_497;
wire n_514;
wire n_270;
wire n_507;
wire n_614;
wire n_305;
wire n_586;
wire n_450;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_473;
wire n_465;
wire n_719;
wire n_566;
wire n_474;
wire n_170;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_168;
wire n_241;
wire n_175;
wire n_687;
wire n_729;
wire n_646;
wire n_650;
wire n_710;
wire n_105;
wire n_743;
wire n_294;
wire n_393;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_307;
wire n_601;
wire n_500;
wire n_661;
wire n_463;
wire n_396;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_143;
wire n_192;
wire n_475;
wire n_554;
wire n_264;
wire n_237;
wire n_668;
A2O1A1Ixp33_ASAP7_75t_SL g485 ( .A1(n_0), .A2(n_189), .B(n_486), .C(n_489), .Y(n_485) );
NAND2xp5_ASAP7_75t_L g491 ( .A(n_1), .B(n_480), .Y(n_491) );
INVx1_ASAP7_75t_L g112 ( .A(n_2), .Y(n_112) );
INVx1_ASAP7_75t_L g238 ( .A(n_3), .Y(n_238) );
NAND2xp5_ASAP7_75t_SL g514 ( .A(n_4), .B(n_177), .Y(n_514) );
AOI21xp5_ASAP7_75t_L g533 ( .A1(n_5), .A2(n_464), .B(n_534), .Y(n_533) );
OAI22xp5_ASAP7_75t_SL g761 ( .A1(n_6), .A2(n_9), .B1(n_447), .B2(n_762), .Y(n_761) );
CKINVDCx20_ASAP7_75t_R g762 ( .A(n_6), .Y(n_762) );
AO21x2_ASAP7_75t_L g542 ( .A1(n_7), .A2(n_194), .B(n_543), .Y(n_542) );
AOI22xp33_ASAP7_75t_L g188 ( .A1(n_8), .A2(n_40), .B1(n_150), .B2(n_162), .Y(n_188) );
AOI22xp5_ASAP7_75t_L g133 ( .A1(n_9), .A2(n_134), .B1(n_135), .B2(n_447), .Y(n_133) );
CKINVDCx20_ASAP7_75t_R g447 ( .A(n_9), .Y(n_447) );
NAND2xp5_ASAP7_75t_L g227 ( .A(n_10), .B(n_194), .Y(n_227) );
AND2x6_ASAP7_75t_L g165 ( .A(n_11), .B(n_166), .Y(n_165) );
A2O1A1Ixp33_ASAP7_75t_L g555 ( .A1(n_12), .A2(n_165), .B(n_467), .C(n_556), .Y(n_555) );
CKINVDCx20_ASAP7_75t_R g750 ( .A(n_13), .Y(n_750) );
INVx1_ASAP7_75t_L g109 ( .A(n_14), .Y(n_109) );
NOR2xp33_ASAP7_75t_L g124 ( .A(n_14), .B(n_41), .Y(n_124) );
INVx1_ASAP7_75t_L g146 ( .A(n_15), .Y(n_146) );
NAND2xp5_ASAP7_75t_L g153 ( .A(n_16), .B(n_154), .Y(n_153) );
INVx1_ASAP7_75t_L g232 ( .A(n_17), .Y(n_232) );
NAND2xp5_ASAP7_75t_SL g548 ( .A(n_18), .B(n_177), .Y(n_548) );
NAND2xp5_ASAP7_75t_L g210 ( .A(n_19), .B(n_192), .Y(n_210) );
AO32x2_ASAP7_75t_L g186 ( .A1(n_20), .A2(n_187), .A3(n_191), .B1(n_193), .B2(n_194), .Y(n_186) );
OAI22xp5_ASAP7_75t_L g127 ( .A1(n_21), .A2(n_100), .B1(n_128), .B2(n_129), .Y(n_127) );
CKINVDCx20_ASAP7_75t_R g129 ( .A(n_21), .Y(n_129) );
AND2x2_ASAP7_75t_L g528 ( .A(n_22), .B(n_142), .Y(n_528) );
NAND2xp5_ASAP7_75t_SL g160 ( .A(n_23), .B(n_150), .Y(n_160) );
NAND2xp5_ASAP7_75t_L g240 ( .A(n_24), .B(n_192), .Y(n_240) );
AOI22xp33_ASAP7_75t_L g190 ( .A1(n_25), .A2(n_56), .B1(n_150), .B2(n_162), .Y(n_190) );
AOI22xp33_ASAP7_75t_SL g203 ( .A1(n_26), .A2(n_82), .B1(n_150), .B2(n_154), .Y(n_203) );
NAND2xp5_ASAP7_75t_SL g180 ( .A(n_27), .B(n_150), .Y(n_180) );
A2O1A1Ixp33_ASAP7_75t_L g466 ( .A1(n_28), .A2(n_193), .B(n_467), .C(n_469), .Y(n_466) );
A2O1A1Ixp33_ASAP7_75t_L g545 ( .A1(n_29), .A2(n_193), .B(n_467), .C(n_546), .Y(n_545) );
BUFx6f_ASAP7_75t_L g158 ( .A(n_30), .Y(n_158) );
NAND2xp5_ASAP7_75t_L g252 ( .A(n_31), .B(n_142), .Y(n_252) );
AOI22xp33_ASAP7_75t_L g102 ( .A1(n_32), .A2(n_103), .B1(n_117), .B2(n_767), .Y(n_102) );
AOI21xp5_ASAP7_75t_L g481 ( .A1(n_33), .A2(n_464), .B(n_482), .Y(n_481) );
NAND2xp5_ASAP7_75t_L g184 ( .A(n_34), .B(n_142), .Y(n_184) );
INVx2_ASAP7_75t_L g152 ( .A(n_35), .Y(n_152) );
A2O1A1Ixp33_ASAP7_75t_L g497 ( .A1(n_36), .A2(n_498), .B(n_499), .C(n_503), .Y(n_497) );
NAND2xp5_ASAP7_75t_SL g247 ( .A(n_37), .B(n_150), .Y(n_247) );
NAND2xp5_ASAP7_75t_L g167 ( .A(n_38), .B(n_142), .Y(n_167) );
NAND2xp5_ASAP7_75t_L g547 ( .A(n_39), .B(n_157), .Y(n_547) );
NAND2xp5_ASAP7_75t_L g108 ( .A(n_41), .B(n_109), .Y(n_108) );
NAND2xp5_ASAP7_75t_L g462 ( .A(n_42), .B(n_463), .Y(n_462) );
CKINVDCx20_ASAP7_75t_R g560 ( .A(n_43), .Y(n_560) );
NAND2xp5_ASAP7_75t_L g527 ( .A(n_44), .B(n_177), .Y(n_527) );
NAND2xp5_ASAP7_75t_L g544 ( .A(n_45), .B(n_464), .Y(n_544) );
A2O1A1Ixp33_ASAP7_75t_L g524 ( .A1(n_46), .A2(n_498), .B(n_503), .C(n_525), .Y(n_524) );
NAND2xp5_ASAP7_75t_SL g220 ( .A(n_47), .B(n_150), .Y(n_220) );
NAND2xp5_ASAP7_75t_SL g119 ( .A(n_48), .B(n_120), .Y(n_119) );
INVx1_ASAP7_75t_L g487 ( .A(n_49), .Y(n_487) );
AOI22xp33_ASAP7_75t_L g201 ( .A1(n_50), .A2(n_91), .B1(n_162), .B2(n_202), .Y(n_201) );
INVx1_ASAP7_75t_L g526 ( .A(n_51), .Y(n_526) );
NAND2xp5_ASAP7_75t_SL g223 ( .A(n_52), .B(n_150), .Y(n_223) );
NAND2xp5_ASAP7_75t_L g234 ( .A(n_53), .B(n_150), .Y(n_234) );
NAND2xp5_ASAP7_75t_L g523 ( .A(n_54), .B(n_464), .Y(n_523) );
NAND2xp5_ASAP7_75t_L g224 ( .A(n_55), .B(n_225), .Y(n_224) );
AOI22xp33_ASAP7_75t_SL g214 ( .A1(n_57), .A2(n_61), .B1(n_150), .B2(n_154), .Y(n_214) );
CKINVDCx20_ASAP7_75t_R g476 ( .A(n_58), .Y(n_476) );
NAND2xp5_ASAP7_75t_SL g149 ( .A(n_59), .B(n_150), .Y(n_149) );
NAND2xp5_ASAP7_75t_SL g251 ( .A(n_60), .B(n_150), .Y(n_251) );
INVx1_ASAP7_75t_L g166 ( .A(n_62), .Y(n_166) );
NAND2xp5_ASAP7_75t_L g516 ( .A(n_63), .B(n_464), .Y(n_516) );
NAND2xp5_ASAP7_75t_L g539 ( .A(n_64), .B(n_480), .Y(n_539) );
A2O1A1Ixp33_ASAP7_75t_L g536 ( .A1(n_65), .A2(n_225), .B(n_235), .C(n_537), .Y(n_536) );
NAND2xp5_ASAP7_75t_L g239 ( .A(n_66), .B(n_150), .Y(n_239) );
INVx1_ASAP7_75t_L g145 ( .A(n_67), .Y(n_145) );
CKINVDCx20_ASAP7_75t_R g756 ( .A(n_68), .Y(n_756) );
NAND2xp5_ASAP7_75t_SL g501 ( .A(n_69), .B(n_177), .Y(n_501) );
AO32x2_ASAP7_75t_L g199 ( .A1(n_70), .A2(n_193), .A3(n_194), .B1(n_200), .B2(n_204), .Y(n_199) );
NAND2xp5_ASAP7_75t_L g557 ( .A(n_71), .B(n_178), .Y(n_557) );
INVx1_ASAP7_75t_L g250 ( .A(n_72), .Y(n_250) );
INVx1_ASAP7_75t_L g175 ( .A(n_73), .Y(n_175) );
CKINVDCx16_ASAP7_75t_R g483 ( .A(n_74), .Y(n_483) );
NAND2xp5_ASAP7_75t_L g470 ( .A(n_75), .B(n_471), .Y(n_470) );
A2O1A1Ixp33_ASAP7_75t_L g511 ( .A1(n_76), .A2(n_467), .B(n_503), .C(n_512), .Y(n_511) );
NOR2xp33_ASAP7_75t_L g758 ( .A(n_77), .B(n_759), .Y(n_758) );
CKINVDCx20_ASAP7_75t_R g764 ( .A(n_77), .Y(n_764) );
NAND2xp5_ASAP7_75t_SL g176 ( .A(n_78), .B(n_154), .Y(n_176) );
CKINVDCx16_ASAP7_75t_R g535 ( .A(n_79), .Y(n_535) );
INVx1_ASAP7_75t_L g116 ( .A(n_80), .Y(n_116) );
NAND2xp5_ASAP7_75t_SL g472 ( .A(n_81), .B(n_473), .Y(n_472) );
NAND2xp5_ASAP7_75t_L g161 ( .A(n_83), .B(n_162), .Y(n_161) );
CKINVDCx20_ASAP7_75t_R g505 ( .A(n_84), .Y(n_505) );
NAND2xp5_ASAP7_75t_SL g181 ( .A(n_85), .B(n_154), .Y(n_181) );
INVx2_ASAP7_75t_L g143 ( .A(n_86), .Y(n_143) );
CKINVDCx20_ASAP7_75t_R g518 ( .A(n_87), .Y(n_518) );
NAND2xp5_ASAP7_75t_SL g558 ( .A(n_88), .B(n_164), .Y(n_558) );
NAND2xp5_ASAP7_75t_L g221 ( .A(n_89), .B(n_154), .Y(n_221) );
INVx2_ASAP7_75t_L g113 ( .A(n_90), .Y(n_113) );
OR2x2_ASAP7_75t_L g121 ( .A(n_90), .B(n_122), .Y(n_121) );
OR2x2_ASAP7_75t_L g450 ( .A(n_90), .B(n_123), .Y(n_450) );
AOI22xp33_ASAP7_75t_L g213 ( .A1(n_92), .A2(n_101), .B1(n_154), .B2(n_155), .Y(n_213) );
NAND2xp5_ASAP7_75t_L g496 ( .A(n_93), .B(n_464), .Y(n_496) );
INVx1_ASAP7_75t_L g500 ( .A(n_94), .Y(n_500) );
INVxp67_ASAP7_75t_L g538 ( .A(n_95), .Y(n_538) );
NAND2xp5_ASAP7_75t_L g248 ( .A(n_96), .B(n_154), .Y(n_248) );
NAND2xp5_ASAP7_75t_L g115 ( .A(n_97), .B(n_116), .Y(n_115) );
INVx1_ASAP7_75t_L g513 ( .A(n_98), .Y(n_513) );
INVx1_ASAP7_75t_L g553 ( .A(n_99), .Y(n_553) );
CKINVDCx20_ASAP7_75t_R g128 ( .A(n_100), .Y(n_128) );
BUFx4f_ASAP7_75t_SL g103 ( .A(n_104), .Y(n_103) );
CKINVDCx20_ASAP7_75t_R g104 ( .A(n_105), .Y(n_104) );
CKINVDCx16_ASAP7_75t_R g105 ( .A(n_106), .Y(n_105) );
INVx2_ASAP7_75t_L g769 ( .A(n_106), .Y(n_769) );
AND2x2_ASAP7_75t_L g106 ( .A(n_107), .B(n_110), .Y(n_106) );
INVx1_ASAP7_75t_L g107 ( .A(n_108), .Y(n_107) );
CKINVDCx14_ASAP7_75t_R g110 ( .A(n_111), .Y(n_110) );
NAND3xp33_ASAP7_75t_SL g111 ( .A(n_112), .B(n_113), .C(n_114), .Y(n_111) );
AND2x2_ASAP7_75t_L g123 ( .A(n_112), .B(n_124), .Y(n_123) );
OR2x2_ASAP7_75t_L g744 ( .A(n_113), .B(n_123), .Y(n_744) );
NOR2x2_ASAP7_75t_L g752 ( .A(n_113), .B(n_122), .Y(n_752) );
INVx1_ASAP7_75t_SL g114 ( .A(n_115), .Y(n_114) );
BUFx3_ASAP7_75t_L g117 ( .A(n_118), .Y(n_117) );
NAND2xp5_ASAP7_75t_L g118 ( .A(n_119), .B(n_125), .Y(n_118) );
INVx1_ASAP7_75t_SL g120 ( .A(n_121), .Y(n_120) );
INVx1_ASAP7_75t_SL g766 ( .A(n_121), .Y(n_766) );
INVx2_ASAP7_75t_L g122 ( .A(n_123), .Y(n_122) );
OAI32xp33_ASAP7_75t_L g125 ( .A1(n_126), .A2(n_749), .A3(n_753), .B1(n_754), .B2(n_757), .Y(n_125) );
OAI22xp5_ASAP7_75t_L g126 ( .A1(n_127), .A2(n_130), .B1(n_745), .B2(n_746), .Y(n_126) );
INVx1_ASAP7_75t_L g745 ( .A(n_127), .Y(n_745) );
INVx1_ASAP7_75t_L g130 ( .A(n_131), .Y(n_130) );
OAI22x1_ASAP7_75t_SL g131 ( .A1(n_132), .A2(n_448), .B1(n_451), .B2(n_742), .Y(n_131) );
INVx1_ASAP7_75t_L g132 ( .A(n_133), .Y(n_132) );
OAI22xp5_ASAP7_75t_SL g747 ( .A1(n_133), .A2(n_452), .B1(n_742), .B2(n_748), .Y(n_747) );
OAI22xp5_ASAP7_75t_SL g759 ( .A1(n_134), .A2(n_135), .B1(n_760), .B2(n_761), .Y(n_759) );
INVx1_ASAP7_75t_L g134 ( .A(n_135), .Y(n_134) );
OR2x2_ASAP7_75t_L g135 ( .A(n_136), .B(n_369), .Y(n_135) );
NAND5xp2_ASAP7_75t_L g136 ( .A(n_137), .B(n_288), .C(n_303), .D(n_329), .E(n_351), .Y(n_136) );
NOR2xp33_ASAP7_75t_SL g137 ( .A(n_138), .B(n_268), .Y(n_137) );
OAI221xp5_ASAP7_75t_L g138 ( .A1(n_139), .A2(n_205), .B1(n_241), .B2(n_257), .C(n_258), .Y(n_138) );
NOR2xp33_ASAP7_75t_SL g139 ( .A(n_140), .B(n_195), .Y(n_139) );
NAND2xp5_ASAP7_75t_L g317 ( .A(n_140), .B(n_318), .Y(n_317) );
INVx1_ASAP7_75t_SL g445 ( .A(n_140), .Y(n_445) );
AND2x2_ASAP7_75t_L g140 ( .A(n_141), .B(n_168), .Y(n_140) );
INVx1_ASAP7_75t_L g285 ( .A(n_141), .Y(n_285) );
AND2x2_ASAP7_75t_L g287 ( .A(n_141), .B(n_186), .Y(n_287) );
AND2x2_ASAP7_75t_L g297 ( .A(n_141), .B(n_185), .Y(n_297) );
HB1xp67_ASAP7_75t_L g315 ( .A(n_141), .Y(n_315) );
INVx1_ASAP7_75t_L g325 ( .A(n_141), .Y(n_325) );
OR2x2_ASAP7_75t_L g363 ( .A(n_141), .B(n_262), .Y(n_363) );
INVx2_ASAP7_75t_L g413 ( .A(n_141), .Y(n_413) );
NAND2xp5_ASAP7_75t_L g430 ( .A(n_141), .B(n_261), .Y(n_430) );
OA21x2_ASAP7_75t_L g141 ( .A1(n_142), .A2(n_147), .B(n_167), .Y(n_141) );
OA21x2_ASAP7_75t_L g171 ( .A1(n_142), .A2(n_172), .B(n_184), .Y(n_171) );
INVx2_ASAP7_75t_L g204 ( .A(n_142), .Y(n_204) );
INVx1_ASAP7_75t_L g477 ( .A(n_142), .Y(n_477) );
AOI21xp5_ASAP7_75t_L g495 ( .A1(n_142), .A2(n_496), .B(n_497), .Y(n_495) );
AOI21xp5_ASAP7_75t_L g522 ( .A1(n_142), .A2(n_523), .B(n_524), .Y(n_522) );
AND2x2_ASAP7_75t_SL g142 ( .A(n_143), .B(n_144), .Y(n_142) );
AND2x2_ASAP7_75t_L g192 ( .A(n_143), .B(n_144), .Y(n_192) );
NAND2xp5_ASAP7_75t_L g144 ( .A(n_145), .B(n_146), .Y(n_144) );
OAI21xp5_ASAP7_75t_L g147 ( .A1(n_148), .A2(n_159), .B(n_165), .Y(n_147) );
AOI21xp5_ASAP7_75t_L g148 ( .A1(n_149), .A2(n_153), .B(n_156), .Y(n_148) );
INVx3_ASAP7_75t_L g174 ( .A(n_150), .Y(n_174) );
HB1xp67_ASAP7_75t_L g515 ( .A(n_150), .Y(n_515) );
BUFx6f_ASAP7_75t_L g150 ( .A(n_151), .Y(n_150) );
INVx1_ASAP7_75t_L g162 ( .A(n_151), .Y(n_162) );
BUFx3_ASAP7_75t_L g202 ( .A(n_151), .Y(n_202) );
AND2x6_ASAP7_75t_L g467 ( .A(n_151), .B(n_468), .Y(n_467) );
INVx2_ASAP7_75t_L g151 ( .A(n_152), .Y(n_151) );
INVx1_ASAP7_75t_L g155 ( .A(n_152), .Y(n_155) );
INVx1_ASAP7_75t_L g226 ( .A(n_152), .Y(n_226) );
INVx2_ASAP7_75t_L g233 ( .A(n_154), .Y(n_233) );
INVx3_ASAP7_75t_L g154 ( .A(n_155), .Y(n_154) );
INVx1_ASAP7_75t_L g156 ( .A(n_157), .Y(n_156) );
INVx1_ASAP7_75t_L g157 ( .A(n_158), .Y(n_157) );
BUFx6f_ASAP7_75t_L g164 ( .A(n_158), .Y(n_164) );
INVx3_ASAP7_75t_L g178 ( .A(n_158), .Y(n_178) );
BUFx6f_ASAP7_75t_L g183 ( .A(n_158), .Y(n_183) );
AND2x2_ASAP7_75t_L g465 ( .A(n_158), .B(n_226), .Y(n_465) );
INVx1_ASAP7_75t_L g468 ( .A(n_158), .Y(n_468) );
AOI21xp5_ASAP7_75t_L g159 ( .A1(n_160), .A2(n_161), .B(n_163), .Y(n_159) );
O2A1O1Ixp5_ASAP7_75t_L g249 ( .A1(n_163), .A2(n_237), .B(n_250), .C(n_251), .Y(n_249) );
INVx2_ASAP7_75t_L g163 ( .A(n_164), .Y(n_163) );
OAI22xp5_ASAP7_75t_L g187 ( .A1(n_164), .A2(n_188), .B1(n_189), .B2(n_190), .Y(n_187) );
OAI22xp5_ASAP7_75t_SL g200 ( .A1(n_164), .A2(n_178), .B1(n_201), .B2(n_203), .Y(n_200) );
OAI22xp5_ASAP7_75t_L g212 ( .A1(n_164), .A2(n_189), .B1(n_213), .B2(n_214), .Y(n_212) );
INVx4_ASAP7_75t_L g488 ( .A(n_164), .Y(n_488) );
OAI21xp5_ASAP7_75t_L g172 ( .A1(n_165), .A2(n_173), .B(n_179), .Y(n_172) );
BUFx3_ASAP7_75t_L g193 ( .A(n_165), .Y(n_193) );
OAI21xp5_ASAP7_75t_L g218 ( .A1(n_165), .A2(n_219), .B(n_222), .Y(n_218) );
OAI21xp5_ASAP7_75t_L g230 ( .A1(n_165), .A2(n_231), .B(n_236), .Y(n_230) );
AND2x4_ASAP7_75t_L g464 ( .A(n_165), .B(n_465), .Y(n_464) );
INVx4_ASAP7_75t_SL g490 ( .A(n_165), .Y(n_490) );
NAND2x1p5_ASAP7_75t_L g554 ( .A(n_165), .B(n_465), .Y(n_554) );
NOR2xp67_ASAP7_75t_L g168 ( .A(n_169), .B(n_185), .Y(n_168) );
INVx1_ASAP7_75t_L g169 ( .A(n_170), .Y(n_169) );
HB1xp67_ASAP7_75t_L g279 ( .A(n_170), .Y(n_279) );
NAND2xp5_ASAP7_75t_L g295 ( .A(n_170), .B(n_296), .Y(n_295) );
AND2x2_ASAP7_75t_SL g345 ( .A(n_170), .B(n_285), .Y(n_345) );
INVx2_ASAP7_75t_L g170 ( .A(n_171), .Y(n_170) );
HB1xp67_ASAP7_75t_L g197 ( .A(n_171), .Y(n_197) );
INVx2_ASAP7_75t_L g262 ( .A(n_171), .Y(n_262) );
OR2x2_ASAP7_75t_L g324 ( .A(n_171), .B(n_325), .Y(n_324) );
O2A1O1Ixp5_ASAP7_75t_SL g173 ( .A1(n_174), .A2(n_175), .B(n_176), .C(n_177), .Y(n_173) );
INVx2_ASAP7_75t_L g189 ( .A(n_177), .Y(n_189) );
AOI21xp5_ASAP7_75t_L g219 ( .A1(n_177), .A2(n_220), .B(n_221), .Y(n_219) );
AOI21xp5_ASAP7_75t_L g246 ( .A1(n_177), .A2(n_247), .B(n_248), .Y(n_246) );
NOR2xp33_ASAP7_75t_L g537 ( .A(n_177), .B(n_538), .Y(n_537) );
INVx5_ASAP7_75t_L g177 ( .A(n_178), .Y(n_177) );
AOI21xp5_ASAP7_75t_L g179 ( .A1(n_180), .A2(n_181), .B(n_182), .Y(n_179) );
INVx1_ASAP7_75t_L g235 ( .A(n_182), .Y(n_235) );
INVx4_ASAP7_75t_L g182 ( .A(n_183), .Y(n_182) );
INVx2_ASAP7_75t_L g471 ( .A(n_183), .Y(n_471) );
AND2x2_ASAP7_75t_L g263 ( .A(n_185), .B(n_199), .Y(n_263) );
AND2x2_ASAP7_75t_L g280 ( .A(n_185), .B(n_260), .Y(n_280) );
INVx2_ASAP7_75t_L g185 ( .A(n_186), .Y(n_185) );
AND2x2_ASAP7_75t_L g198 ( .A(n_186), .B(n_199), .Y(n_198) );
BUFx2_ASAP7_75t_L g283 ( .A(n_186), .Y(n_283) );
AND2x2_ASAP7_75t_L g412 ( .A(n_186), .B(n_413), .Y(n_412) );
AOI21xp5_ASAP7_75t_L g222 ( .A1(n_189), .A2(n_223), .B(n_224), .Y(n_222) );
O2A1O1Ixp33_ASAP7_75t_L g236 ( .A1(n_189), .A2(n_237), .B(n_238), .C(n_239), .Y(n_236) );
INVx2_ASAP7_75t_L g229 ( .A(n_191), .Y(n_229) );
NOR2xp33_ASAP7_75t_L g559 ( .A(n_191), .B(n_560), .Y(n_559) );
INVx1_ASAP7_75t_L g191 ( .A(n_192), .Y(n_191) );
BUFx6f_ASAP7_75t_L g194 ( .A(n_192), .Y(n_194) );
NAND3xp33_ASAP7_75t_L g211 ( .A(n_193), .B(n_212), .C(n_215), .Y(n_211) );
OAI21xp5_ASAP7_75t_L g245 ( .A1(n_193), .A2(n_246), .B(n_249), .Y(n_245) );
INVx4_ASAP7_75t_L g215 ( .A(n_194), .Y(n_215) );
OA21x2_ASAP7_75t_L g217 ( .A1(n_194), .A2(n_218), .B(n_227), .Y(n_217) );
HB1xp67_ASAP7_75t_L g532 ( .A(n_194), .Y(n_532) );
AOI21xp5_ASAP7_75t_L g543 ( .A1(n_194), .A2(n_544), .B(n_545), .Y(n_543) );
INVx1_ASAP7_75t_L g257 ( .A(n_195), .Y(n_257) );
AND2x2_ASAP7_75t_L g195 ( .A(n_196), .B(n_198), .Y(n_195) );
AND2x2_ASAP7_75t_L g375 ( .A(n_196), .B(n_263), .Y(n_375) );
INVx1_ASAP7_75t_L g196 ( .A(n_197), .Y(n_196) );
AND2x2_ASAP7_75t_L g376 ( .A(n_197), .B(n_287), .Y(n_376) );
O2A1O1Ixp33_ASAP7_75t_L g343 ( .A1(n_198), .A2(n_344), .B(n_346), .C(n_348), .Y(n_343) );
NAND2xp5_ASAP7_75t_L g353 ( .A(n_198), .B(n_344), .Y(n_353) );
AOI221xp5_ASAP7_75t_L g416 ( .A1(n_198), .A2(n_274), .B1(n_417), .B2(n_418), .C(n_420), .Y(n_416) );
INVx1_ASAP7_75t_L g260 ( .A(n_199), .Y(n_260) );
INVx1_ASAP7_75t_L g296 ( .A(n_199), .Y(n_296) );
BUFx6f_ASAP7_75t_L g305 ( .A(n_199), .Y(n_305) );
INVx2_ASAP7_75t_L g489 ( .A(n_202), .Y(n_489) );
HB1xp67_ASAP7_75t_L g502 ( .A(n_202), .Y(n_502) );
INVx1_ASAP7_75t_L g474 ( .A(n_204), .Y(n_474) );
INVx1_ASAP7_75t_SL g205 ( .A(n_206), .Y(n_205) );
AND2x2_ASAP7_75t_L g206 ( .A(n_207), .B(n_216), .Y(n_206) );
AND2x2_ASAP7_75t_L g322 ( .A(n_207), .B(n_267), .Y(n_322) );
NAND2xp5_ASAP7_75t_L g341 ( .A(n_207), .B(n_342), .Y(n_341) );
INVx2_ASAP7_75t_L g207 ( .A(n_208), .Y(n_207) );
NOR2xp33_ASAP7_75t_L g290 ( .A(n_208), .B(n_291), .Y(n_290) );
OR2x2_ASAP7_75t_L g414 ( .A(n_208), .B(n_415), .Y(n_414) );
INVx1_ASAP7_75t_L g446 ( .A(n_208), .Y(n_446) );
INVx2_ASAP7_75t_L g208 ( .A(n_209), .Y(n_208) );
INVx3_ASAP7_75t_L g276 ( .A(n_209), .Y(n_276) );
AND2x2_ASAP7_75t_L g302 ( .A(n_209), .B(n_256), .Y(n_302) );
NOR2x1_ASAP7_75t_L g311 ( .A(n_209), .B(n_312), .Y(n_311) );
AND2x2_ASAP7_75t_L g318 ( .A(n_209), .B(n_319), .Y(n_318) );
AND2x4_ASAP7_75t_L g209 ( .A(n_210), .B(n_211), .Y(n_209) );
INVx1_ASAP7_75t_L g254 ( .A(n_210), .Y(n_254) );
AO21x1_ASAP7_75t_L g253 ( .A1(n_212), .A2(n_215), .B(n_254), .Y(n_253) );
INVx3_ASAP7_75t_L g480 ( .A(n_215), .Y(n_480) );
NOR2xp33_ASAP7_75t_L g504 ( .A(n_215), .B(n_505), .Y(n_504) );
AO21x2_ASAP7_75t_L g509 ( .A1(n_215), .A2(n_510), .B(n_517), .Y(n_509) );
NOR2xp33_ASAP7_75t_L g517 ( .A(n_215), .B(n_518), .Y(n_517) );
AO21x2_ASAP7_75t_L g551 ( .A1(n_215), .A2(n_552), .B(n_559), .Y(n_551) );
NAND2xp5_ASAP7_75t_L g393 ( .A(n_216), .B(n_358), .Y(n_393) );
INVx1_ASAP7_75t_SL g397 ( .A(n_216), .Y(n_397) );
AND2x2_ASAP7_75t_L g216 ( .A(n_217), .B(n_228), .Y(n_216) );
INVx3_ASAP7_75t_L g256 ( .A(n_217), .Y(n_256) );
AND2x2_ASAP7_75t_L g267 ( .A(n_217), .B(n_244), .Y(n_267) );
AND2x2_ASAP7_75t_L g289 ( .A(n_217), .B(n_290), .Y(n_289) );
AND2x2_ASAP7_75t_L g334 ( .A(n_217), .B(n_328), .Y(n_334) );
NAND2xp5_ASAP7_75t_L g415 ( .A(n_217), .B(n_266), .Y(n_415) );
INVx2_ASAP7_75t_L g237 ( .A(n_225), .Y(n_237) );
INVx1_ASAP7_75t_L g225 ( .A(n_226), .Y(n_225) );
AND2x2_ASAP7_75t_L g255 ( .A(n_228), .B(n_256), .Y(n_255) );
INVx2_ASAP7_75t_L g266 ( .A(n_228), .Y(n_266) );
NAND2xp5_ASAP7_75t_L g291 ( .A(n_228), .B(n_244), .Y(n_291) );
AND2x2_ASAP7_75t_L g327 ( .A(n_228), .B(n_328), .Y(n_327) );
OA21x2_ASAP7_75t_L g228 ( .A1(n_229), .A2(n_230), .B(n_240), .Y(n_228) );
OA21x2_ASAP7_75t_L g244 ( .A1(n_229), .A2(n_245), .B(n_252), .Y(n_244) );
O2A1O1Ixp33_ASAP7_75t_L g231 ( .A1(n_232), .A2(n_233), .B(n_234), .C(n_235), .Y(n_231) );
AOI21xp5_ASAP7_75t_L g546 ( .A1(n_233), .A2(n_547), .B(n_548), .Y(n_546) );
AOI21xp5_ASAP7_75t_L g556 ( .A1(n_233), .A2(n_557), .B(n_558), .Y(n_556) );
O2A1O1Ixp33_ASAP7_75t_L g512 ( .A1(n_235), .A2(n_513), .B(n_514), .C(n_515), .Y(n_512) );
AOI21xp5_ASAP7_75t_L g469 ( .A1(n_237), .A2(n_470), .B(n_472), .Y(n_469) );
INVx1_ASAP7_75t_L g241 ( .A(n_242), .Y(n_241) );
AND2x2_ASAP7_75t_L g242 ( .A(n_243), .B(n_255), .Y(n_242) );
INVx1_ASAP7_75t_L g307 ( .A(n_243), .Y(n_307) );
AND2x2_ASAP7_75t_L g349 ( .A(n_243), .B(n_350), .Y(n_349) );
NAND2xp5_ASAP7_75t_SL g355 ( .A(n_243), .B(n_270), .Y(n_355) );
AOI21xp5_ASAP7_75t_SL g429 ( .A1(n_243), .A2(n_261), .B(n_284), .Y(n_429) );
AND2x2_ASAP7_75t_L g243 ( .A(n_244), .B(n_253), .Y(n_243) );
OR2x2_ASAP7_75t_L g272 ( .A(n_244), .B(n_253), .Y(n_272) );
AND2x2_ASAP7_75t_L g319 ( .A(n_244), .B(n_256), .Y(n_319) );
INVx2_ASAP7_75t_L g328 ( .A(n_244), .Y(n_328) );
INVx1_ASAP7_75t_L g434 ( .A(n_244), .Y(n_434) );
AND2x2_ASAP7_75t_L g358 ( .A(n_253), .B(n_328), .Y(n_358) );
INVx1_ASAP7_75t_L g383 ( .A(n_253), .Y(n_383) );
AND2x2_ASAP7_75t_L g292 ( .A(n_255), .B(n_276), .Y(n_292) );
AND2x2_ASAP7_75t_L g304 ( .A(n_255), .B(n_305), .Y(n_304) );
INVx2_ASAP7_75t_SL g422 ( .A(n_255), .Y(n_422) );
INVx2_ASAP7_75t_L g312 ( .A(n_256), .Y(n_312) );
AND2x2_ASAP7_75t_L g350 ( .A(n_256), .B(n_266), .Y(n_350) );
NAND2xp5_ASAP7_75t_L g433 ( .A(n_256), .B(n_434), .Y(n_433) );
OAI21xp33_ASAP7_75t_L g258 ( .A1(n_259), .A2(n_263), .B(n_264), .Y(n_258) );
AND2x2_ASAP7_75t_L g365 ( .A(n_259), .B(n_366), .Y(n_365) );
INVx1_ASAP7_75t_L g419 ( .A(n_259), .Y(n_419) );
AND2x2_ASAP7_75t_L g259 ( .A(n_260), .B(n_261), .Y(n_259) );
INVx1_ASAP7_75t_L g339 ( .A(n_260), .Y(n_339) );
BUFx2_ASAP7_75t_L g438 ( .A(n_260), .Y(n_438) );
BUFx2_ASAP7_75t_L g309 ( .A(n_261), .Y(n_309) );
AND2x2_ASAP7_75t_L g411 ( .A(n_261), .B(n_412), .Y(n_411) );
INVx2_ASAP7_75t_L g261 ( .A(n_262), .Y(n_261) );
INVx1_ASAP7_75t_L g394 ( .A(n_262), .Y(n_394) );
AND2x4_ASAP7_75t_L g321 ( .A(n_263), .B(n_284), .Y(n_321) );
NAND2xp5_ASAP7_75t_SL g357 ( .A(n_263), .B(n_345), .Y(n_357) );
AOI32xp33_ASAP7_75t_L g281 ( .A1(n_264), .A2(n_282), .A3(n_284), .B1(n_286), .B2(n_287), .Y(n_281) );
AND2x2_ASAP7_75t_L g264 ( .A(n_265), .B(n_267), .Y(n_264) );
INVx3_ASAP7_75t_L g270 ( .A(n_265), .Y(n_270) );
OR2x2_ASAP7_75t_L g406 ( .A(n_265), .B(n_362), .Y(n_406) );
INVx2_ASAP7_75t_L g265 ( .A(n_266), .Y(n_265) );
AND2x2_ASAP7_75t_L g275 ( .A(n_266), .B(n_276), .Y(n_275) );
AND2x2_ASAP7_75t_L g382 ( .A(n_266), .B(n_383), .Y(n_382) );
AND2x2_ASAP7_75t_L g274 ( .A(n_267), .B(n_275), .Y(n_274) );
AND2x2_ASAP7_75t_L g286 ( .A(n_267), .B(n_276), .Y(n_286) );
INVx1_ASAP7_75t_L g407 ( .A(n_267), .Y(n_407) );
NAND2xp5_ASAP7_75t_L g440 ( .A(n_267), .B(n_382), .Y(n_440) );
A2O1A1Ixp33_ASAP7_75t_L g268 ( .A1(n_269), .A2(n_273), .B(n_277), .C(n_281), .Y(n_268) );
OAI322xp33_ASAP7_75t_L g377 ( .A1(n_269), .A2(n_314), .A3(n_378), .B1(n_380), .B2(n_384), .C1(n_385), .C2(n_389), .Y(n_377) );
NAND2xp5_ASAP7_75t_L g269 ( .A(n_270), .B(n_271), .Y(n_269) );
INVxp67_ASAP7_75t_L g342 ( .A(n_270), .Y(n_342) );
INVx1_ASAP7_75t_SL g271 ( .A(n_272), .Y(n_271) );
OR2x2_ASAP7_75t_L g396 ( .A(n_272), .B(n_397), .Y(n_396) );
NOR2xp33_ASAP7_75t_L g443 ( .A(n_272), .B(n_312), .Y(n_443) );
INVxp67_ASAP7_75t_L g273 ( .A(n_274), .Y(n_273) );
INVx1_ASAP7_75t_L g335 ( .A(n_275), .Y(n_335) );
OR2x2_ASAP7_75t_L g421 ( .A(n_276), .B(n_422), .Y(n_421) );
INVx1_ASAP7_75t_L g277 ( .A(n_278), .Y(n_277) );
AND2x2_ASAP7_75t_L g278 ( .A(n_279), .B(n_280), .Y(n_278) );
NAND2xp5_ASAP7_75t_L g337 ( .A(n_279), .B(n_338), .Y(n_337) );
AND2x2_ASAP7_75t_L g330 ( .A(n_280), .B(n_309), .Y(n_330) );
AND2x2_ASAP7_75t_L g401 ( .A(n_280), .B(n_314), .Y(n_401) );
NAND2xp5_ASAP7_75t_L g423 ( .A(n_280), .B(n_388), .Y(n_423) );
AOI221xp5_ASAP7_75t_L g288 ( .A1(n_282), .A2(n_289), .B1(n_292), .B2(n_293), .C(n_298), .Y(n_288) );
OR2x2_ASAP7_75t_L g299 ( .A(n_282), .B(n_295), .Y(n_299) );
AND2x2_ASAP7_75t_L g387 ( .A(n_282), .B(n_388), .Y(n_387) );
AOI32xp33_ASAP7_75t_L g426 ( .A1(n_282), .A2(n_312), .A3(n_427), .B1(n_428), .B2(n_431), .Y(n_426) );
INVx2_ASAP7_75t_L g282 ( .A(n_283), .Y(n_282) );
NAND3xp33_ASAP7_75t_L g360 ( .A(n_283), .B(n_319), .C(n_342), .Y(n_360) );
AND2x2_ASAP7_75t_L g386 ( .A(n_283), .B(n_379), .Y(n_386) );
INVxp67_ASAP7_75t_L g366 ( .A(n_284), .Y(n_366) );
BUFx3_ASAP7_75t_L g284 ( .A(n_285), .Y(n_284) );
NAND2xp5_ASAP7_75t_SL g395 ( .A(n_287), .B(n_339), .Y(n_395) );
INVx2_ASAP7_75t_L g405 ( .A(n_287), .Y(n_405) );
NOR2xp33_ASAP7_75t_L g418 ( .A(n_287), .B(n_419), .Y(n_418) );
INVx1_ASAP7_75t_L g374 ( .A(n_290), .Y(n_374) );
OR2x2_ASAP7_75t_L g300 ( .A(n_291), .B(n_301), .Y(n_300) );
NOR2xp33_ASAP7_75t_L g410 ( .A(n_293), .B(n_411), .Y(n_410) );
AND2x2_ASAP7_75t_L g293 ( .A(n_294), .B(n_297), .Y(n_293) );
INVx1_ASAP7_75t_SL g294 ( .A(n_295), .Y(n_294) );
HB1xp67_ASAP7_75t_L g379 ( .A(n_296), .Y(n_379) );
AND2x2_ASAP7_75t_L g338 ( .A(n_297), .B(n_339), .Y(n_338) );
INVx1_ASAP7_75t_L g384 ( .A(n_297), .Y(n_384) );
HB1xp67_ASAP7_75t_L g409 ( .A(n_297), .Y(n_409) );
NOR2xp33_ASAP7_75t_L g298 ( .A(n_299), .B(n_300), .Y(n_298) );
AOI21xp33_ASAP7_75t_SL g323 ( .A1(n_299), .A2(n_324), .B(n_326), .Y(n_323) );
INVx1_ASAP7_75t_L g301 ( .A(n_302), .Y(n_301) );
AND2x2_ASAP7_75t_L g417 ( .A(n_302), .B(n_327), .Y(n_417) );
AOI211xp5_ASAP7_75t_L g303 ( .A1(n_304), .A2(n_306), .B(n_316), .C(n_323), .Y(n_303) );
AND2x2_ASAP7_75t_L g347 ( .A(n_305), .B(n_315), .Y(n_347) );
INVx2_ASAP7_75t_L g362 ( .A(n_305), .Y(n_362) );
OR2x2_ASAP7_75t_L g400 ( .A(n_305), .B(n_363), .Y(n_400) );
NAND2xp5_ASAP7_75t_L g442 ( .A(n_305), .B(n_443), .Y(n_442) );
AOI211xp5_ASAP7_75t_SL g306 ( .A1(n_307), .A2(n_308), .B(n_310), .C(n_313), .Y(n_306) );
INVxp67_ASAP7_75t_L g308 ( .A(n_309), .Y(n_308) );
NAND2xp5_ASAP7_75t_L g346 ( .A(n_309), .B(n_347), .Y(n_346) );
OAI211xp5_ASAP7_75t_L g428 ( .A1(n_310), .A2(n_405), .B(n_429), .C(n_430), .Y(n_428) );
INVx1_ASAP7_75t_L g310 ( .A(n_311), .Y(n_310) );
NAND2x1p5_ASAP7_75t_L g326 ( .A(n_311), .B(n_327), .Y(n_326) );
AND2x2_ASAP7_75t_L g368 ( .A(n_312), .B(n_358), .Y(n_368) );
INVx1_ASAP7_75t_L g373 ( .A(n_312), .Y(n_373) );
INVx1_ASAP7_75t_L g313 ( .A(n_314), .Y(n_313) );
INVx1_ASAP7_75t_L g314 ( .A(n_315), .Y(n_314) );
NAND2xp5_ASAP7_75t_SL g316 ( .A(n_317), .B(n_320), .Y(n_316) );
INVxp33_ASAP7_75t_L g424 ( .A(n_318), .Y(n_424) );
AND2x2_ASAP7_75t_L g403 ( .A(n_319), .B(n_382), .Y(n_403) );
NAND2xp5_ASAP7_75t_L g320 ( .A(n_321), .B(n_322), .Y(n_320) );
AOI21xp5_ASAP7_75t_L g385 ( .A1(n_324), .A2(n_386), .B(n_387), .Y(n_385) );
OAI322xp33_ASAP7_75t_L g404 ( .A1(n_326), .A2(n_405), .A3(n_406), .B1(n_407), .B2(n_408), .C1(n_410), .C2(n_414), .Y(n_404) );
AOI221xp5_ASAP7_75t_L g329 ( .A1(n_330), .A2(n_331), .B1(n_336), .B2(n_340), .C(n_343), .Y(n_329) );
INVx2_ASAP7_75t_L g331 ( .A(n_332), .Y(n_331) );
OR2x2_ASAP7_75t_L g332 ( .A(n_333), .B(n_335), .Y(n_332) );
INVx1_ASAP7_75t_L g333 ( .A(n_334), .Y(n_333) );
AND2x2_ASAP7_75t_L g381 ( .A(n_334), .B(n_382), .Y(n_381) );
INVx1_ASAP7_75t_L g336 ( .A(n_337), .Y(n_336) );
INVx1_ASAP7_75t_L g425 ( .A(n_338), .Y(n_425) );
INVxp67_ASAP7_75t_L g340 ( .A(n_341), .Y(n_340) );
NOR2xp33_ASAP7_75t_L g427 ( .A(n_341), .B(n_361), .Y(n_427) );
INVx2_ASAP7_75t_L g344 ( .A(n_345), .Y(n_344) );
INVx1_ASAP7_75t_SL g348 ( .A(n_349), .Y(n_348) );
AND2x2_ASAP7_75t_L g390 ( .A(n_350), .B(n_358), .Y(n_390) );
AOI221xp5_ASAP7_75t_L g351 ( .A1(n_352), .A2(n_354), .B1(n_356), .B2(n_358), .C(n_359), .Y(n_351) );
INVx1_ASAP7_75t_L g352 ( .A(n_353), .Y(n_352) );
AOI221xp5_ASAP7_75t_L g370 ( .A1(n_354), .A2(n_371), .B1(n_375), .B2(n_376), .C(n_377), .Y(n_370) );
INVx1_ASAP7_75t_L g354 ( .A(n_355), .Y(n_354) );
INVxp67_ASAP7_75t_L g356 ( .A(n_357), .Y(n_356) );
NAND2xp5_ASAP7_75t_L g372 ( .A(n_358), .B(n_373), .Y(n_372) );
OAI22xp5_ASAP7_75t_L g359 ( .A1(n_360), .A2(n_361), .B1(n_364), .B2(n_367), .Y(n_359) );
OR2x2_ASAP7_75t_L g361 ( .A(n_362), .B(n_363), .Y(n_361) );
INVx2_ASAP7_75t_SL g388 ( .A(n_363), .Y(n_388) );
INVxp67_ASAP7_75t_L g364 ( .A(n_365), .Y(n_364) );
INVx1_ASAP7_75t_L g367 ( .A(n_368), .Y(n_367) );
NAND5xp2_ASAP7_75t_L g369 ( .A(n_370), .B(n_391), .C(n_416), .D(n_426), .E(n_436), .Y(n_369) );
NAND2xp5_ASAP7_75t_SL g371 ( .A(n_372), .B(n_374), .Y(n_371) );
NOR4xp25_ASAP7_75t_L g444 ( .A(n_373), .B(n_379), .C(n_445), .D(n_446), .Y(n_444) );
AOI221xp5_ASAP7_75t_L g436 ( .A1(n_376), .A2(n_437), .B1(n_439), .B2(n_441), .C(n_444), .Y(n_436) );
INVx1_ASAP7_75t_L g378 ( .A(n_379), .Y(n_378) );
INVx1_ASAP7_75t_L g380 ( .A(n_381), .Y(n_380) );
INVx1_ASAP7_75t_L g435 ( .A(n_382), .Y(n_435) );
OAI322xp33_ASAP7_75t_L g392 ( .A1(n_386), .A2(n_393), .A3(n_394), .B1(n_395), .B2(n_396), .C1(n_398), .C2(n_402), .Y(n_392) );
INVx1_ASAP7_75t_SL g389 ( .A(n_390), .Y(n_389) );
NOR2xp33_ASAP7_75t_L g391 ( .A(n_392), .B(n_404), .Y(n_391) );
NOR2xp33_ASAP7_75t_L g398 ( .A(n_399), .B(n_401), .Y(n_398) );
INVx2_ASAP7_75t_L g399 ( .A(n_400), .Y(n_399) );
INVx1_ASAP7_75t_L g402 ( .A(n_403), .Y(n_402) );
INVx1_ASAP7_75t_L g408 ( .A(n_409), .Y(n_408) );
AND2x2_ASAP7_75t_L g437 ( .A(n_412), .B(n_438), .Y(n_437) );
OAI22xp33_ASAP7_75t_L g420 ( .A1(n_421), .A2(n_423), .B1(n_424), .B2(n_425), .Y(n_420) );
INVx1_ASAP7_75t_L g431 ( .A(n_432), .Y(n_431) );
OR2x2_ASAP7_75t_L g432 ( .A(n_433), .B(n_435), .Y(n_432) );
INVx1_ASAP7_75t_L g439 ( .A(n_440), .Y(n_439) );
INVxp67_ASAP7_75t_L g441 ( .A(n_442), .Y(n_441) );
INVx2_ASAP7_75t_L g448 ( .A(n_449), .Y(n_448) );
INVx2_ASAP7_75t_L g748 ( .A(n_449), .Y(n_748) );
INVx1_ASAP7_75t_L g449 ( .A(n_450), .Y(n_449) );
INVx2_ASAP7_75t_L g451 ( .A(n_452), .Y(n_451) );
AND2x2_ASAP7_75t_SL g452 ( .A(n_453), .B(n_697), .Y(n_452) );
NOR2xp33_ASAP7_75t_L g453 ( .A(n_454), .B(n_632), .Y(n_453) );
NAND4xp25_ASAP7_75t_SL g454 ( .A(n_455), .B(n_577), .C(n_601), .D(n_624), .Y(n_454) );
AOI221xp5_ASAP7_75t_L g455 ( .A1(n_456), .A2(n_519), .B1(n_549), .B2(n_561), .C(n_564), .Y(n_455) );
INVx1_ASAP7_75t_L g456 ( .A(n_457), .Y(n_456) );
NAND2xp5_ASAP7_75t_L g457 ( .A(n_458), .B(n_492), .Y(n_457) );
AOI22xp33_ASAP7_75t_L g567 ( .A1(n_458), .A2(n_478), .B1(n_520), .B2(n_568), .Y(n_567) );
NAND2xp5_ASAP7_75t_L g635 ( .A(n_458), .B(n_493), .Y(n_635) );
AND2x2_ASAP7_75t_L g654 ( .A(n_458), .B(n_655), .Y(n_654) );
NAND2xp5_ASAP7_75t_L g724 ( .A(n_458), .B(n_638), .Y(n_724) );
AND2x4_ASAP7_75t_L g458 ( .A(n_459), .B(n_478), .Y(n_458) );
AND2x2_ASAP7_75t_L g592 ( .A(n_459), .B(n_493), .Y(n_592) );
NAND2xp5_ASAP7_75t_L g606 ( .A(n_459), .B(n_607), .Y(n_606) );
OR2x2_ASAP7_75t_L g615 ( .A(n_459), .B(n_616), .Y(n_615) );
AND2x2_ASAP7_75t_L g620 ( .A(n_459), .B(n_479), .Y(n_620) );
INVx2_ASAP7_75t_L g652 ( .A(n_459), .Y(n_652) );
HB1xp67_ASAP7_75t_L g696 ( .A(n_459), .Y(n_696) );
AND2x2_ASAP7_75t_L g713 ( .A(n_459), .B(n_590), .Y(n_713) );
INVx5_ASAP7_75t_L g459 ( .A(n_460), .Y(n_459) );
AND2x2_ASAP7_75t_L g631 ( .A(n_460), .B(n_590), .Y(n_631) );
AND2x4_ASAP7_75t_L g645 ( .A(n_460), .B(n_478), .Y(n_645) );
HB1xp67_ASAP7_75t_L g649 ( .A(n_460), .Y(n_649) );
AND2x2_ASAP7_75t_L g669 ( .A(n_460), .B(n_584), .Y(n_669) );
AND2x2_ASAP7_75t_L g719 ( .A(n_460), .B(n_494), .Y(n_719) );
AND2x2_ASAP7_75t_L g729 ( .A(n_460), .B(n_479), .Y(n_729) );
OR2x6_ASAP7_75t_L g460 ( .A(n_461), .B(n_475), .Y(n_460) );
AOI21xp5_ASAP7_75t_SL g461 ( .A1(n_462), .A2(n_466), .B(n_474), .Y(n_461) );
BUFx2_ASAP7_75t_L g463 ( .A(n_464), .Y(n_463) );
INVx5_ASAP7_75t_L g484 ( .A(n_467), .Y(n_484) );
INVx2_ASAP7_75t_L g473 ( .A(n_471), .Y(n_473) );
O2A1O1Ixp33_ASAP7_75t_L g499 ( .A1(n_473), .A2(n_500), .B(n_501), .C(n_502), .Y(n_499) );
O2A1O1Ixp33_ASAP7_75t_L g525 ( .A1(n_473), .A2(n_502), .B(n_526), .C(n_527), .Y(n_525) );
NOR2xp33_ASAP7_75t_L g475 ( .A(n_476), .B(n_477), .Y(n_475) );
AND2x2_ASAP7_75t_L g585 ( .A(n_478), .B(n_493), .Y(n_585) );
HB1xp67_ASAP7_75t_L g600 ( .A(n_478), .Y(n_600) );
NAND2xp5_ASAP7_75t_L g626 ( .A(n_478), .B(n_627), .Y(n_626) );
INVx1_ASAP7_75t_L g675 ( .A(n_478), .Y(n_675) );
INVx2_ASAP7_75t_L g478 ( .A(n_479), .Y(n_478) );
AND2x2_ASAP7_75t_L g563 ( .A(n_479), .B(n_508), .Y(n_563) );
AND2x2_ASAP7_75t_L g590 ( .A(n_479), .B(n_509), .Y(n_590) );
OA21x2_ASAP7_75t_L g479 ( .A1(n_480), .A2(n_481), .B(n_491), .Y(n_479) );
O2A1O1Ixp33_ASAP7_75t_SL g482 ( .A1(n_483), .A2(n_484), .B(n_485), .C(n_490), .Y(n_482) );
INVx2_ASAP7_75t_L g498 ( .A(n_484), .Y(n_498) );
O2A1O1Ixp33_ASAP7_75t_L g534 ( .A1(n_484), .A2(n_490), .B(n_535), .C(n_536), .Y(n_534) );
NOR2xp33_ASAP7_75t_L g486 ( .A(n_487), .B(n_488), .Y(n_486) );
INVx1_ASAP7_75t_L g503 ( .A(n_490), .Y(n_503) );
NAND2xp5_ASAP7_75t_L g648 ( .A(n_492), .B(n_649), .Y(n_648) );
AND2x2_ASAP7_75t_L g492 ( .A(n_493), .B(n_506), .Y(n_492) );
OR2x2_ASAP7_75t_L g616 ( .A(n_493), .B(n_507), .Y(n_616) );
AND2x2_ASAP7_75t_L g653 ( .A(n_493), .B(n_563), .Y(n_653) );
NAND2xp5_ASAP7_75t_L g664 ( .A(n_493), .B(n_584), .Y(n_664) );
HB1xp67_ASAP7_75t_L g668 ( .A(n_493), .Y(n_668) );
NAND2xp5_ASAP7_75t_L g737 ( .A(n_493), .B(n_620), .Y(n_737) );
INVx5_ASAP7_75t_L g493 ( .A(n_494), .Y(n_493) );
BUFx2_ASAP7_75t_L g562 ( .A(n_494), .Y(n_562) );
AND2x2_ASAP7_75t_L g571 ( .A(n_494), .B(n_507), .Y(n_571) );
AND2x2_ASAP7_75t_L g687 ( .A(n_494), .B(n_582), .Y(n_687) );
NAND2xp5_ASAP7_75t_L g709 ( .A(n_494), .B(n_620), .Y(n_709) );
OR2x6_ASAP7_75t_L g494 ( .A(n_495), .B(n_504), .Y(n_494) );
INVx1_ASAP7_75t_L g506 ( .A(n_507), .Y(n_506) );
HB1xp67_ASAP7_75t_L g655 ( .A(n_507), .Y(n_655) );
INVx2_ASAP7_75t_L g507 ( .A(n_508), .Y(n_507) );
HB1xp67_ASAP7_75t_L g607 ( .A(n_508), .Y(n_607) );
INVx2_ASAP7_75t_L g508 ( .A(n_509), .Y(n_508) );
BUFx2_ASAP7_75t_L g584 ( .A(n_509), .Y(n_584) );
NAND2xp5_ASAP7_75t_L g510 ( .A(n_511), .B(n_516), .Y(n_510) );
NOR2xp33_ASAP7_75t_L g519 ( .A(n_520), .B(n_529), .Y(n_519) );
NOR2xp33_ASAP7_75t_L g716 ( .A(n_520), .B(n_597), .Y(n_716) );
HB1xp67_ASAP7_75t_L g520 ( .A(n_521), .Y(n_520) );
NOR2xp33_ASAP7_75t_L g549 ( .A(n_521), .B(n_550), .Y(n_549) );
AND2x2_ASAP7_75t_L g568 ( .A(n_521), .B(n_569), .Y(n_568) );
INVx5_ASAP7_75t_SL g576 ( .A(n_521), .Y(n_576) );
OR2x2_ASAP7_75t_L g599 ( .A(n_521), .B(n_569), .Y(n_599) );
OR2x2_ASAP7_75t_L g609 ( .A(n_521), .B(n_610), .Y(n_609) );
AND2x2_ASAP7_75t_L g672 ( .A(n_521), .B(n_531), .Y(n_672) );
AND2x2_ASAP7_75t_SL g710 ( .A(n_521), .B(n_530), .Y(n_710) );
NOR4xp25_ASAP7_75t_L g731 ( .A(n_521), .B(n_652), .C(n_732), .D(n_733), .Y(n_731) );
AND2x2_ASAP7_75t_L g741 ( .A(n_521), .B(n_573), .Y(n_741) );
OR2x6_ASAP7_75t_L g521 ( .A(n_522), .B(n_528), .Y(n_521) );
INVx2_ASAP7_75t_L g529 ( .A(n_530), .Y(n_529) );
AND2x2_ASAP7_75t_L g566 ( .A(n_530), .B(n_562), .Y(n_566) );
NAND2xp5_ASAP7_75t_L g735 ( .A(n_530), .B(n_568), .Y(n_735) );
AND2x2_ASAP7_75t_L g530 ( .A(n_531), .B(n_540), .Y(n_530) );
OR2x2_ASAP7_75t_L g575 ( .A(n_531), .B(n_576), .Y(n_575) );
INVx3_ASAP7_75t_L g582 ( .A(n_531), .Y(n_582) );
NAND2xp5_ASAP7_75t_L g594 ( .A(n_531), .B(n_551), .Y(n_594) );
INVxp67_ASAP7_75t_L g597 ( .A(n_531), .Y(n_597) );
NAND2xp5_ASAP7_75t_L g610 ( .A(n_531), .B(n_569), .Y(n_610) );
NAND2xp5_ASAP7_75t_L g663 ( .A(n_531), .B(n_541), .Y(n_663) );
AND2x2_ASAP7_75t_L g678 ( .A(n_531), .B(n_573), .Y(n_678) );
OR2x2_ASAP7_75t_L g707 ( .A(n_531), .B(n_541), .Y(n_707) );
OA21x2_ASAP7_75t_L g531 ( .A1(n_532), .A2(n_533), .B(n_539), .Y(n_531) );
NAND2xp5_ASAP7_75t_L g611 ( .A(n_540), .B(n_612), .Y(n_611) );
NOR2xp33_ASAP7_75t_L g715 ( .A(n_540), .B(n_576), .Y(n_715) );
OR2x2_ASAP7_75t_L g736 ( .A(n_540), .B(n_613), .Y(n_736) );
INVx1_ASAP7_75t_SL g540 ( .A(n_541), .Y(n_540) );
OR2x2_ASAP7_75t_L g550 ( .A(n_541), .B(n_551), .Y(n_550) );
AND2x2_ASAP7_75t_L g573 ( .A(n_541), .B(n_569), .Y(n_573) );
NAND2xp5_ASAP7_75t_SL g588 ( .A(n_541), .B(n_551), .Y(n_588) );
AND2x2_ASAP7_75t_L g658 ( .A(n_541), .B(n_582), .Y(n_658) );
AND2x2_ASAP7_75t_L g692 ( .A(n_541), .B(n_576), .Y(n_692) );
INVx2_ASAP7_75t_L g541 ( .A(n_542), .Y(n_541) );
NAND2xp5_ASAP7_75t_L g595 ( .A(n_542), .B(n_576), .Y(n_595) );
AND2x2_ASAP7_75t_L g623 ( .A(n_542), .B(n_551), .Y(n_623) );
NAND2xp5_ASAP7_75t_L g630 ( .A(n_549), .B(n_631), .Y(n_630) );
AOI221xp5_ASAP7_75t_L g690 ( .A1(n_550), .A2(n_638), .B1(n_674), .B2(n_691), .C(n_693), .Y(n_690) );
INVx5_ASAP7_75t_SL g569 ( .A(n_551), .Y(n_569) );
OAI21xp5_ASAP7_75t_L g552 ( .A1(n_553), .A2(n_554), .B(n_555), .Y(n_552) );
AND2x2_ASAP7_75t_L g561 ( .A(n_562), .B(n_563), .Y(n_561) );
OAI33xp33_ASAP7_75t_L g589 ( .A1(n_562), .A2(n_590), .A3(n_591), .B1(n_593), .B2(n_596), .B3(n_600), .Y(n_589) );
OR2x2_ASAP7_75t_L g605 ( .A(n_562), .B(n_606), .Y(n_605) );
AOI322xp5_ASAP7_75t_L g714 ( .A1(n_562), .A2(n_631), .A3(n_638), .B1(n_715), .B2(n_716), .C1(n_717), .C2(n_720), .Y(n_714) );
NAND2xp5_ASAP7_75t_L g732 ( .A(n_562), .B(n_590), .Y(n_732) );
A2O1A1Ixp33_ASAP7_75t_SL g738 ( .A1(n_562), .A2(n_590), .B(n_739), .C(n_741), .Y(n_738) );
AOI221xp5_ASAP7_75t_L g577 ( .A1(n_563), .A2(n_578), .B1(n_583), .B2(n_586), .C(n_589), .Y(n_577) );
INVx1_ASAP7_75t_L g670 ( .A(n_563), .Y(n_670) );
NAND2xp5_ASAP7_75t_L g718 ( .A(n_563), .B(n_719), .Y(n_718) );
OAI22xp33_ASAP7_75t_L g564 ( .A1(n_565), .A2(n_567), .B1(n_570), .B2(n_572), .Y(n_564) );
INVx1_ASAP7_75t_SL g565 ( .A(n_566), .Y(n_565) );
AND2x2_ASAP7_75t_L g647 ( .A(n_568), .B(n_582), .Y(n_647) );
AND2x2_ASAP7_75t_L g705 ( .A(n_568), .B(n_706), .Y(n_705) );
OR2x2_ASAP7_75t_L g613 ( .A(n_569), .B(n_576), .Y(n_613) );
NAND2xp5_ASAP7_75t_L g641 ( .A(n_569), .B(n_582), .Y(n_641) );
INVx1_ASAP7_75t_L g570 ( .A(n_571), .Y(n_570) );
NAND2xp5_ASAP7_75t_L g643 ( .A(n_571), .B(n_644), .Y(n_643) );
NAND2xp5_ASAP7_75t_L g703 ( .A(n_571), .B(n_649), .Y(n_703) );
OAI321xp33_ASAP7_75t_L g722 ( .A1(n_571), .A2(n_644), .A3(n_723), .B1(n_724), .B2(n_725), .C(n_726), .Y(n_722) );
INVx1_ASAP7_75t_L g689 ( .A(n_572), .Y(n_689) );
NAND2xp5_ASAP7_75t_L g572 ( .A(n_573), .B(n_574), .Y(n_572) );
NAND2xp5_ASAP7_75t_L g579 ( .A(n_573), .B(n_580), .Y(n_579) );
AND2x2_ASAP7_75t_L g628 ( .A(n_573), .B(n_576), .Y(n_628) );
AOI321xp33_ASAP7_75t_L g686 ( .A1(n_573), .A2(n_590), .A3(n_687), .B1(n_688), .B2(n_689), .C(n_690), .Y(n_686) );
INVx1_ASAP7_75t_L g574 ( .A(n_575), .Y(n_574) );
OR2x2_ASAP7_75t_L g603 ( .A(n_575), .B(n_588), .Y(n_603) );
NAND2xp5_ASAP7_75t_L g581 ( .A(n_576), .B(n_582), .Y(n_581) );
NAND2xp5_ASAP7_75t_L g657 ( .A(n_576), .B(n_658), .Y(n_657) );
NAND2xp5_ASAP7_75t_L g699 ( .A(n_576), .B(n_662), .Y(n_699) );
INVx1_ASAP7_75t_L g578 ( .A(n_579), .Y(n_578) );
AND2x4_ASAP7_75t_L g622 ( .A(n_580), .B(n_623), .Y(n_622) );
INVx2_ASAP7_75t_L g580 ( .A(n_581), .Y(n_580) );
OR2x2_ASAP7_75t_L g587 ( .A(n_581), .B(n_588), .Y(n_587) );
INVx1_ASAP7_75t_L g695 ( .A(n_582), .Y(n_695) );
AND2x2_ASAP7_75t_L g583 ( .A(n_584), .B(n_585), .Y(n_583) );
NAND2xp5_ASAP7_75t_L g637 ( .A(n_585), .B(n_638), .Y(n_637) );
INVx2_ASAP7_75t_L g586 ( .A(n_587), .Y(n_586) );
INVx1_ASAP7_75t_L g618 ( .A(n_590), .Y(n_618) );
INVx1_ASAP7_75t_L g591 ( .A(n_592), .Y(n_591) );
NOR2xp33_ASAP7_75t_L g676 ( .A(n_592), .B(n_627), .Y(n_676) );
OR2x2_ASAP7_75t_L g593 ( .A(n_594), .B(n_595), .Y(n_593) );
OR2x2_ASAP7_75t_L g640 ( .A(n_595), .B(n_641), .Y(n_640) );
INVx1_ASAP7_75t_SL g685 ( .A(n_595), .Y(n_685) );
OAI22xp5_ASAP7_75t_L g642 ( .A1(n_596), .A2(n_643), .B1(n_646), .B2(n_648), .Y(n_642) );
NAND2xp5_ASAP7_75t_L g596 ( .A(n_597), .B(n_598), .Y(n_596) );
INVx1_ASAP7_75t_SL g598 ( .A(n_599), .Y(n_598) );
OR2x2_ASAP7_75t_L g740 ( .A(n_599), .B(n_663), .Y(n_740) );
AOI221xp5_ASAP7_75t_L g601 ( .A1(n_602), .A2(n_604), .B1(n_608), .B2(n_614), .C(n_617), .Y(n_601) );
INVx1_ASAP7_75t_SL g602 ( .A(n_603), .Y(n_602) );
INVx2_ASAP7_75t_L g604 ( .A(n_605), .Y(n_604) );
BUFx2_ASAP7_75t_L g638 ( .A(n_607), .Y(n_638) );
NAND2xp5_ASAP7_75t_L g608 ( .A(n_609), .B(n_611), .Y(n_608) );
INVx1_ASAP7_75t_SL g684 ( .A(n_610), .Y(n_684) );
NAND2xp5_ASAP7_75t_L g661 ( .A(n_612), .B(n_662), .Y(n_661) );
AOI21xp5_ASAP7_75t_L g679 ( .A1(n_612), .A2(n_680), .B(n_682), .Y(n_679) );
INVx2_ASAP7_75t_L g612 ( .A(n_613), .Y(n_612) );
OR2x2_ASAP7_75t_L g725 ( .A(n_613), .B(n_707), .Y(n_725) );
INVx1_ASAP7_75t_L g614 ( .A(n_615), .Y(n_614) );
INVx2_ASAP7_75t_SL g627 ( .A(n_616), .Y(n_627) );
AOI21xp33_ASAP7_75t_L g617 ( .A1(n_618), .A2(n_619), .B(n_621), .Y(n_617) );
INVx1_ASAP7_75t_L g619 ( .A(n_620), .Y(n_619) );
INVx2_ASAP7_75t_SL g621 ( .A(n_622), .Y(n_621) );
AND2x2_ASAP7_75t_L g671 ( .A(n_623), .B(n_672), .Y(n_671) );
INVxp67_ASAP7_75t_L g733 ( .A(n_623), .Y(n_733) );
AOI21xp5_ASAP7_75t_L g624 ( .A1(n_625), .A2(n_628), .B(n_629), .Y(n_624) );
INVx1_ASAP7_75t_L g625 ( .A(n_626), .Y(n_625) );
NAND2xp5_ASAP7_75t_L g681 ( .A(n_627), .B(n_645), .Y(n_681) );
INVxp67_ASAP7_75t_L g629 ( .A(n_630), .Y(n_629) );
INVx1_ASAP7_75t_L g702 ( .A(n_631), .Y(n_702) );
NAND5xp2_ASAP7_75t_L g632 ( .A(n_633), .B(n_650), .C(n_659), .D(n_679), .E(n_686), .Y(n_632) );
O2A1O1Ixp33_ASAP7_75t_L g633 ( .A1(n_634), .A2(n_636), .B(n_639), .C(n_642), .Y(n_633) );
INVx1_ASAP7_75t_L g634 ( .A(n_635), .Y(n_634) );
INVx1_ASAP7_75t_L g636 ( .A(n_637), .Y(n_636) );
INVx1_ASAP7_75t_L g674 ( .A(n_638), .Y(n_674) );
CKINVDCx16_ASAP7_75t_R g639 ( .A(n_640), .Y(n_639) );
INVx1_ASAP7_75t_SL g644 ( .A(n_645), .Y(n_644) );
NOR2xp33_ASAP7_75t_L g711 ( .A(n_646), .B(n_712), .Y(n_711) );
INVx1_ASAP7_75t_L g646 ( .A(n_647), .Y(n_646) );
INVx1_ASAP7_75t_L g688 ( .A(n_648), .Y(n_688) );
OAI21xp5_ASAP7_75t_SL g650 ( .A1(n_651), .A2(n_654), .B(n_656), .Y(n_650) );
AOI221xp5_ASAP7_75t_L g704 ( .A1(n_651), .A2(n_705), .B1(n_708), .B2(n_710), .C(n_711), .Y(n_704) );
AND2x2_ASAP7_75t_L g651 ( .A(n_652), .B(n_653), .Y(n_651) );
AOI321xp33_ASAP7_75t_L g659 ( .A1(n_652), .A2(n_660), .A3(n_664), .B1(n_665), .B2(n_671), .C(n_673), .Y(n_659) );
INVx1_ASAP7_75t_L g656 ( .A(n_657), .Y(n_656) );
INVx1_ASAP7_75t_L g660 ( .A(n_661), .Y(n_660) );
INVx1_ASAP7_75t_SL g662 ( .A(n_663), .Y(n_662) );
INVx1_ASAP7_75t_L g730 ( .A(n_664), .Y(n_730) );
NAND2xp5_ASAP7_75t_SL g665 ( .A(n_666), .B(n_670), .Y(n_665) );
INVx1_ASAP7_75t_L g666 ( .A(n_667), .Y(n_666) );
AND2x2_ASAP7_75t_L g682 ( .A(n_667), .B(n_683), .Y(n_682) );
AND2x2_ASAP7_75t_L g667 ( .A(n_668), .B(n_669), .Y(n_667) );
NOR2xp67_ASAP7_75t_SL g694 ( .A(n_668), .B(n_675), .Y(n_694) );
AOI321xp33_ASAP7_75t_SL g726 ( .A1(n_671), .A2(n_727), .A3(n_728), .B1(n_729), .B2(n_730), .C(n_731), .Y(n_726) );
O2A1O1Ixp33_ASAP7_75t_L g673 ( .A1(n_674), .A2(n_675), .B(n_676), .C(n_677), .Y(n_673) );
INVx1_ASAP7_75t_SL g677 ( .A(n_678), .Y(n_677) );
INVx1_ASAP7_75t_L g680 ( .A(n_681), .Y(n_680) );
AND2x2_ASAP7_75t_L g683 ( .A(n_684), .B(n_685), .Y(n_683) );
NAND2xp5_ASAP7_75t_L g721 ( .A(n_684), .B(n_692), .Y(n_721) );
INVx1_ASAP7_75t_L g691 ( .A(n_692), .Y(n_691) );
NAND3xp33_ASAP7_75t_L g693 ( .A(n_694), .B(n_695), .C(n_696), .Y(n_693) );
NOR3xp33_ASAP7_75t_L g697 ( .A(n_698), .B(n_722), .C(n_734), .Y(n_697) );
OAI211xp5_ASAP7_75t_SL g698 ( .A1(n_699), .A2(n_700), .B(n_704), .C(n_714), .Y(n_698) );
INVxp67_ASAP7_75t_L g700 ( .A(n_701), .Y(n_700) );
NAND2xp5_ASAP7_75t_SL g701 ( .A(n_702), .B(n_703), .Y(n_701) );
OAI221xp5_ASAP7_75t_L g734 ( .A1(n_703), .A2(n_735), .B1(n_736), .B2(n_737), .C(n_738), .Y(n_734) );
INVx1_ASAP7_75t_L g723 ( .A(n_705), .Y(n_723) );
INVx1_ASAP7_75t_SL g706 ( .A(n_707), .Y(n_706) );
INVx1_ASAP7_75t_L g708 ( .A(n_709), .Y(n_708) );
INVx1_ASAP7_75t_SL g712 ( .A(n_713), .Y(n_712) );
INVx1_ASAP7_75t_L g717 ( .A(n_718), .Y(n_717) );
INVx1_ASAP7_75t_L g720 ( .A(n_721), .Y(n_720) );
INVx1_ASAP7_75t_SL g727 ( .A(n_725), .Y(n_727) );
INVx1_ASAP7_75t_L g728 ( .A(n_729), .Y(n_728) );
CKINVDCx14_ASAP7_75t_R g739 ( .A(n_740), .Y(n_739) );
INVx2_ASAP7_75t_L g742 ( .A(n_743), .Y(n_742) );
INVx1_ASAP7_75t_L g743 ( .A(n_744), .Y(n_743) );
INVx1_ASAP7_75t_L g746 ( .A(n_747), .Y(n_746) );
NOR2xp33_ASAP7_75t_L g749 ( .A(n_750), .B(n_751), .Y(n_749) );
INVx3_ASAP7_75t_SL g751 ( .A(n_752), .Y(n_751) );
INVx1_ASAP7_75t_SL g753 ( .A(n_754), .Y(n_753) );
BUFx2_ASAP7_75t_L g754 ( .A(n_755), .Y(n_754) );
INVx2_ASAP7_75t_L g755 ( .A(n_756), .Y(n_755) );
NOR3xp33_ASAP7_75t_L g757 ( .A(n_758), .B(n_763), .C(n_766), .Y(n_757) );
INVx1_ASAP7_75t_L g765 ( .A(n_759), .Y(n_765) );
INVx1_ASAP7_75t_L g760 ( .A(n_761), .Y(n_760) );
NOR2xp33_ASAP7_75t_L g763 ( .A(n_764), .B(n_765), .Y(n_763) );
INVx1_ASAP7_75t_L g767 ( .A(n_768), .Y(n_767) );
INVx1_ASAP7_75t_L g768 ( .A(n_769), .Y(n_768) );
endmodule