module real_aes_8210_n_99 (n_17, n_28, n_76, n_56, n_34, n_98, n_90, n_82, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_83, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_91, n_43, n_96, n_54, n_35, n_42, n_15, n_9, n_23, n_72, n_95, n_44, n_7, n_4, n_80, n_6, n_12, n_68, n_79, n_69, n_46, n_59, n_25, n_73, n_77, n_81, n_48, n_37, n_97, n_70, n_50, n_89, n_26, n_86, n_93, n_13, n_24, n_2, n_55, n_62, n_84, n_67, n_92, n_33, n_88, n_14, n_11, n_85, n_16, n_94, n_39, n_5, n_45, n_60, n_38, n_87, n_0, n_78, n_63, n_1, n_53, n_36, n_99);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_98;
input n_90;
input n_82;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_83;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_91;
input n_43;
input n_96;
input n_54;
input n_35;
input n_42;
input n_15;
input n_9;
input n_23;
input n_72;
input n_95;
input n_44;
input n_7;
input n_4;
input n_80;
input n_6;
input n_12;
input n_68;
input n_79;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_81;
input n_48;
input n_37;
input n_97;
input n_70;
input n_50;
input n_89;
input n_26;
input n_86;
input n_93;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_84;
input n_67;
input n_92;
input n_33;
input n_88;
input n_14;
input n_11;
input n_85;
input n_16;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_87;
input n_0;
input n_78;
input n_63;
input n_1;
input n_53;
input n_36;
output n_99;
wire n_480;
wire n_113;
wire n_476;
wire n_599;
wire n_187;
wire n_436;
wire n_684;
wire n_257;
wire n_390;
wire n_185;
wire n_285;
wire n_624;
wire n_618;
wire n_522;
wire n_485;
wire n_222;
wire n_631;
wire n_287;
wire n_357;
wire n_503;
wire n_635;
wire n_386;
wire n_673;
wire n_518;
wire n_254;
wire n_207;
wire n_665;
wire n_667;
wire n_580;
wire n_577;
wire n_469;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_718;
wire n_318;
wire n_355;
wire n_239;
wire n_669;
wire n_100;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_742;
wire n_112;
wire n_319;
wire n_421;
wire n_364;
wire n_555;
wire n_329;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_169;
wire n_242;
wire n_376;
wire n_549;
wire n_571;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_448;
wire n_556;
wire n_341;
wire n_545;
wire n_593;
wire n_232;
wire n_460;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_537;
wire n_551;
wire n_320;
wire n_666;
wire n_560;
wire n_260;
wire n_660;
wire n_594;
wire n_186;
wire n_138;
wire n_696;
wire n_704;
wire n_453;
wire n_374;
wire n_379;
wire n_647;
wire n_235;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_161;
wire n_189;
wire n_271;
wire n_489;
wire n_548;
wire n_427;
wire n_678;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_519;
wire n_564;
wire n_638;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_512;
wire n_395;
wire n_332;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_116;
wire n_625;
wire n_462;
wire n_289;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_716;
wire n_213;
wire n_478;
wire n_356;
wire n_584;
wire n_408;
wire n_553;
wire n_184;
wire n_372;
wire n_528;
wire n_578;
wire n_202;
wire n_495;
wire n_370;
wire n_384;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_467;
wire n_327;
wire n_106;
wire n_466;
wire n_559;
wire n_636;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_726;
wire n_343;
wire n_369;
wire n_517;
wire n_683;
wire n_174;
wire n_570;
wire n_675;
wire n_530;
wire n_104;
wire n_535;
wire n_732;
wire n_211;
wire n_281;
wire n_496;
wire n_693;
wire n_173;
wire n_468;
wire n_234;
wire n_284;
wire n_153;
wire n_316;
wire n_532;
wire n_656;
wire n_178;
wire n_409;
wire n_523;
wire n_298;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_297;
wire n_383;
wire n_529;
wire n_119;
wire n_310;
wire n_455;
wire n_504;
wire n_725;
wire n_164;
wire n_671;
wire n_231;
wire n_547;
wire n_102;
wire n_659;
wire n_634;
wire n_682;
wire n_454;
wire n_122;
wire n_443;
wire n_565;
wire n_608;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_267;
wire n_218;
wire n_737;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_722;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_331;
wire n_182;
wire n_417;
wire n_363;
wire n_449;
wire n_607;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_142;
wire n_561;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_655;
wire n_654;
wire n_527;
wire n_505;
wire n_434;
wire n_502;
wire n_600;
wire n_731;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_733;
wire n_552;
wire n_402;
wire n_602;
wire n_617;
wire n_171;
wire n_676;
wire n_658;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_146;
wire n_432;
wire n_255;
wire n_226;
wire n_286;
wire n_416;
wire n_410;
wire n_120;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_695;
wire n_685;
wire n_165;
wire n_361;
wire n_632;
wire n_246;
wire n_176;
wire n_412;
wire n_542;
wire n_163;
wire n_645;
wire n_557;
wire n_714;
wire n_488;
wire n_501;
wire n_251;
wire n_642;
wire n_613;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_702;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_734;
wire n_110;
wire n_392;
wire n_562;
wire n_150;
wire n_147;
wire n_288;
wire n_404;
wire n_713;
wire n_598;
wire n_735;
wire n_728;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_569;
wire n_563;
wire n_188;
wire n_269;
wire n_430;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_193;
wire n_397;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_649;
wire n_663;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_707;
wire n_622;
wire n_470;
wire n_133;
wire n_494;
wire n_711;
wire n_377;
wire n_273;
wire n_723;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_265;
wire n_354;
wire n_720;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_730;
wire n_643;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_148;
wire n_498;
wire n_481;
wire n_691;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_487;
wire n_233;
wire n_290;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_155;
wire n_243;
wire n_692;
wire n_544;
wire n_268;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_101;
wire n_738;
wire n_701;
wire n_309;
wire n_344;
wire n_107;
wire n_229;
wire n_482;
wire n_520;
wire n_633;
wire n_679;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_262;
wire n_630;
wire n_689;
wire n_715;
wire n_134;
wire n_420;
wire n_336;
wire n_349;
wire n_612;
wire n_195;
wire n_438;
wire n_300;
wire n_252;
wire n_741;
wire n_283;
wire n_314;
wire n_249;
wire n_623;
wire n_446;
wire n_721;
wire n_221;
wire n_681;
wire n_156;
wire n_359;
wire n_456;
wire n_717;
wire n_312;
wire n_266;
wire n_183;
wire n_712;
wire n_205;
wire n_433;
wire n_335;
wire n_177;
wire n_516;
wire n_313;
wire n_627;
wire n_739;
wire n_140;
wire n_521;
wire n_418;
wire n_422;
wire n_524;
wire n_219;
wire n_705;
wire n_180;
wire n_212;
wire n_210;
wire n_575;
wire n_325;
wire n_479;
wire n_338;
wire n_442;
wire n_740;
wire n_371;
wire n_698;
wire n_103;
wire n_541;
wire n_166;
wire n_224;
wire n_151;
wire n_546;
wire n_587;
wire n_639;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_724;
wire n_440;
wire n_525;
wire n_674;
wire n_644;
wire n_152;
wire n_198;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_414;
wire n_123;
wire n_279;
wire n_686;
wire n_543;
wire n_497;
wire n_514;
wire n_507;
wire n_270;
wire n_614;
wire n_305;
wire n_586;
wire n_450;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_465;
wire n_473;
wire n_719;
wire n_566;
wire n_474;
wire n_170;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_729;
wire n_168;
wire n_175;
wire n_241;
wire n_687;
wire n_646;
wire n_650;
wire n_710;
wire n_743;
wire n_105;
wire n_294;
wire n_393;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_500;
wire n_307;
wire n_601;
wire n_661;
wire n_463;
wire n_396;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_143;
wire n_192;
wire n_475;
wire n_554;
wire n_264;
wire n_237;
wire n_668;
A2O1A1Ixp33_ASAP7_75t_SL g262 ( .A1(n_0), .A2(n_263), .B(n_264), .C(n_267), .Y(n_262) );
NAND2xp5_ASAP7_75t_L g268 ( .A(n_1), .B(n_251), .Y(n_268) );
INVx1_ASAP7_75t_L g106 ( .A(n_2), .Y(n_106) );
NAND2xp5_ASAP7_75t_SL g178 ( .A(n_3), .B(n_179), .Y(n_178) );
A2O1A1Ixp33_ASAP7_75t_L g522 ( .A1(n_4), .A2(n_140), .B(n_143), .C(n_523), .Y(n_522) );
AOI21xp5_ASAP7_75t_L g546 ( .A1(n_5), .A2(n_135), .B(n_547), .Y(n_546) );
AOI21xp5_ASAP7_75t_L g244 ( .A1(n_6), .A2(n_135), .B(n_245), .Y(n_244) );
AOI222xp33_ASAP7_75t_SL g123 ( .A1(n_7), .A2(n_62), .B1(n_124), .B2(n_730), .C1(n_731), .C2(n_735), .Y(n_123) );
NAND2xp5_ASAP7_75t_L g553 ( .A(n_8), .B(n_251), .Y(n_553) );
AO21x2_ASAP7_75t_L g206 ( .A1(n_9), .A2(n_170), .B(n_207), .Y(n_206) );
AOI22xp33_ASAP7_75t_L g99 ( .A1(n_10), .A2(n_100), .B1(n_110), .B2(n_743), .Y(n_99) );
AND2x6_ASAP7_75t_L g140 ( .A(n_11), .B(n_141), .Y(n_140) );
A2O1A1Ixp33_ASAP7_75t_L g223 ( .A1(n_12), .A2(n_140), .B(n_143), .C(n_224), .Y(n_223) );
INVx1_ASAP7_75t_L g491 ( .A(n_13), .Y(n_491) );
NAND2xp5_ASAP7_75t_L g104 ( .A(n_14), .B(n_40), .Y(n_104) );
NOR2xp33_ASAP7_75t_L g121 ( .A(n_14), .B(n_40), .Y(n_121) );
NAND2xp5_ASAP7_75t_SL g525 ( .A(n_15), .B(n_227), .Y(n_525) );
INVx1_ASAP7_75t_L g161 ( .A(n_16), .Y(n_161) );
NAND2xp5_ASAP7_75t_SL g213 ( .A(n_17), .B(n_179), .Y(n_213) );
A2O1A1Ixp33_ASAP7_75t_L g508 ( .A1(n_18), .A2(n_180), .B(n_509), .C(n_511), .Y(n_508) );
NAND2xp5_ASAP7_75t_L g512 ( .A(n_19), .B(n_251), .Y(n_512) );
NAND2xp5_ASAP7_75t_L g482 ( .A(n_20), .B(n_155), .Y(n_482) );
A2O1A1Ixp33_ASAP7_75t_L g142 ( .A1(n_21), .A2(n_143), .B(n_146), .C(n_154), .Y(n_142) );
A2O1A1Ixp33_ASAP7_75t_L g498 ( .A1(n_22), .A2(n_215), .B(n_266), .C(n_499), .Y(n_498) );
NAND2xp5_ASAP7_75t_SL g542 ( .A(n_23), .B(n_227), .Y(n_542) );
NAND2xp5_ASAP7_75t_SL g464 ( .A(n_24), .B(n_227), .Y(n_464) );
CKINVDCx16_ASAP7_75t_R g538 ( .A(n_25), .Y(n_538) );
INVx1_ASAP7_75t_L g463 ( .A(n_26), .Y(n_463) );
A2O1A1Ixp33_ASAP7_75t_L g209 ( .A1(n_27), .A2(n_143), .B(n_154), .C(n_210), .Y(n_209) );
BUFx6f_ASAP7_75t_L g139 ( .A(n_28), .Y(n_139) );
CKINVDCx20_ASAP7_75t_R g521 ( .A(n_29), .Y(n_521) );
INVx1_ASAP7_75t_L g479 ( .A(n_30), .Y(n_479) );
AOI21xp5_ASAP7_75t_L g259 ( .A1(n_31), .A2(n_135), .B(n_260), .Y(n_259) );
INVx2_ASAP7_75t_L g138 ( .A(n_32), .Y(n_138) );
A2O1A1Ixp33_ASAP7_75t_L g191 ( .A1(n_33), .A2(n_183), .B(n_192), .C(n_194), .Y(n_191) );
CKINVDCx20_ASAP7_75t_R g528 ( .A(n_34), .Y(n_528) );
A2O1A1Ixp33_ASAP7_75t_L g549 ( .A1(n_35), .A2(n_266), .B(n_550), .C(n_552), .Y(n_549) );
INVxp67_ASAP7_75t_L g480 ( .A(n_36), .Y(n_480) );
NAND2xp5_ASAP7_75t_L g211 ( .A(n_37), .B(n_212), .Y(n_211) );
A2O1A1Ixp33_ASAP7_75t_L g461 ( .A1(n_38), .A2(n_143), .B(n_154), .C(n_462), .Y(n_461) );
CKINVDCx14_ASAP7_75t_R g548 ( .A(n_39), .Y(n_548) );
A2O1A1Ixp33_ASAP7_75t_L g488 ( .A1(n_41), .A2(n_267), .B(n_489), .C(n_490), .Y(n_488) );
NAND2xp5_ASAP7_75t_L g133 ( .A(n_42), .B(n_134), .Y(n_133) );
CKINVDCx20_ASAP7_75t_R g229 ( .A(n_43), .Y(n_229) );
NAND2xp5_ASAP7_75t_L g238 ( .A(n_44), .B(n_179), .Y(n_238) );
NAND2xp5_ASAP7_75t_L g208 ( .A(n_45), .B(n_135), .Y(n_208) );
CKINVDCx20_ASAP7_75t_R g466 ( .A(n_46), .Y(n_466) );
CKINVDCx20_ASAP7_75t_R g476 ( .A(n_47), .Y(n_476) );
A2O1A1Ixp33_ASAP7_75t_L g235 ( .A1(n_48), .A2(n_183), .B(n_192), .C(n_236), .Y(n_235) );
INVx1_ASAP7_75t_L g265 ( .A(n_49), .Y(n_265) );
OAI22xp5_ASAP7_75t_L g741 ( .A1(n_50), .A2(n_125), .B1(n_733), .B2(n_742), .Y(n_741) );
CKINVDCx16_ASAP7_75t_R g742 ( .A(n_50), .Y(n_742) );
INVx1_ASAP7_75t_L g237 ( .A(n_51), .Y(n_237) );
INVx1_ASAP7_75t_L g497 ( .A(n_52), .Y(n_497) );
NAND2xp5_ASAP7_75t_L g234 ( .A(n_53), .B(n_135), .Y(n_234) );
CKINVDCx20_ASAP7_75t_R g163 ( .A(n_54), .Y(n_163) );
CKINVDCx14_ASAP7_75t_R g487 ( .A(n_55), .Y(n_487) );
INVx1_ASAP7_75t_L g141 ( .A(n_56), .Y(n_141) );
NAND2xp5_ASAP7_75t_L g185 ( .A(n_57), .B(n_135), .Y(n_185) );
NAND2xp5_ASAP7_75t_L g250 ( .A(n_58), .B(n_251), .Y(n_250) );
A2O1A1Ixp33_ASAP7_75t_L g247 ( .A1(n_59), .A2(n_153), .B(n_176), .C(n_248), .Y(n_247) );
CKINVDCx20_ASAP7_75t_R g122 ( .A(n_60), .Y(n_122) );
INVx1_ASAP7_75t_L g160 ( .A(n_61), .Y(n_160) );
CKINVDCx20_ASAP7_75t_R g730 ( .A(n_62), .Y(n_730) );
INVx1_ASAP7_75t_SL g551 ( .A(n_63), .Y(n_551) );
CKINVDCx20_ASAP7_75t_R g114 ( .A(n_64), .Y(n_114) );
NAND2xp5_ASAP7_75t_SL g196 ( .A(n_65), .B(n_179), .Y(n_196) );
NAND2xp5_ASAP7_75t_L g501 ( .A(n_66), .B(n_251), .Y(n_501) );
NAND2xp5_ASAP7_75t_L g225 ( .A(n_67), .B(n_180), .Y(n_225) );
INVx1_ASAP7_75t_L g541 ( .A(n_68), .Y(n_541) );
CKINVDCx16_ASAP7_75t_R g261 ( .A(n_69), .Y(n_261) );
NAND2xp5_ASAP7_75t_L g147 ( .A(n_70), .B(n_148), .Y(n_147) );
A2O1A1Ixp33_ASAP7_75t_L g173 ( .A1(n_71), .A2(n_143), .B(n_174), .C(n_183), .Y(n_173) );
CKINVDCx16_ASAP7_75t_R g246 ( .A(n_72), .Y(n_246) );
INVx1_ASAP7_75t_L g109 ( .A(n_73), .Y(n_109) );
AOI21xp5_ASAP7_75t_L g485 ( .A1(n_74), .A2(n_135), .B(n_486), .Y(n_485) );
CKINVDCx20_ASAP7_75t_R g544 ( .A(n_75), .Y(n_544) );
AOI21xp5_ASAP7_75t_L g505 ( .A1(n_76), .A2(n_135), .B(n_506), .Y(n_505) );
AOI21xp5_ASAP7_75t_L g474 ( .A1(n_77), .A2(n_134), .B(n_475), .Y(n_474) );
CKINVDCx16_ASAP7_75t_R g460 ( .A(n_78), .Y(n_460) );
INVx1_ASAP7_75t_L g507 ( .A(n_79), .Y(n_507) );
NAND2xp5_ASAP7_75t_SL g150 ( .A(n_80), .B(n_151), .Y(n_150) );
CKINVDCx20_ASAP7_75t_R g200 ( .A(n_81), .Y(n_200) );
AOI21xp5_ASAP7_75t_L g495 ( .A1(n_82), .A2(n_135), .B(n_496), .Y(n_495) );
INVx1_ASAP7_75t_L g510 ( .A(n_83), .Y(n_510) );
INVx2_ASAP7_75t_L g158 ( .A(n_84), .Y(n_158) );
INVx1_ASAP7_75t_L g524 ( .A(n_85), .Y(n_524) );
CKINVDCx20_ASAP7_75t_R g187 ( .A(n_86), .Y(n_187) );
NAND2xp5_ASAP7_75t_SL g226 ( .A(n_87), .B(n_227), .Y(n_226) );
NAND3xp33_ASAP7_75t_SL g105 ( .A(n_88), .B(n_106), .C(n_107), .Y(n_105) );
OR2x2_ASAP7_75t_L g118 ( .A(n_88), .B(n_119), .Y(n_118) );
OR2x2_ASAP7_75t_L g452 ( .A(n_88), .B(n_120), .Y(n_452) );
INVx2_ASAP7_75t_L g729 ( .A(n_88), .Y(n_729) );
A2O1A1Ixp33_ASAP7_75t_L g539 ( .A1(n_89), .A2(n_143), .B(n_183), .C(n_540), .Y(n_539) );
NAND2xp5_ASAP7_75t_L g190 ( .A(n_90), .B(n_135), .Y(n_190) );
INVx1_ASAP7_75t_L g195 ( .A(n_91), .Y(n_195) );
INVxp67_ASAP7_75t_L g249 ( .A(n_92), .Y(n_249) );
NAND2xp5_ASAP7_75t_L g492 ( .A(n_93), .B(n_170), .Y(n_492) );
INVx2_ASAP7_75t_L g500 ( .A(n_94), .Y(n_500) );
NAND2xp5_ASAP7_75t_L g108 ( .A(n_95), .B(n_109), .Y(n_108) );
INVx1_ASAP7_75t_L g175 ( .A(n_96), .Y(n_175) );
INVx1_ASAP7_75t_L g221 ( .A(n_97), .Y(n_221) );
AND2x2_ASAP7_75t_L g239 ( .A(n_98), .B(n_157), .Y(n_239) );
INVx1_ASAP7_75t_L g100 ( .A(n_101), .Y(n_100) );
INVx1_ASAP7_75t_L g101 ( .A(n_102), .Y(n_101) );
CKINVDCx20_ASAP7_75t_R g743 ( .A(n_102), .Y(n_743) );
CKINVDCx12_ASAP7_75t_R g102 ( .A(n_103), .Y(n_102) );
OR2x2_ASAP7_75t_L g103 ( .A(n_104), .B(n_105), .Y(n_103) );
AND2x2_ASAP7_75t_L g120 ( .A(n_106), .B(n_121), .Y(n_120) );
INVx1_ASAP7_75t_SL g107 ( .A(n_108), .Y(n_107) );
AOI22x1_ASAP7_75t_L g110 ( .A1(n_111), .A2(n_123), .B1(n_738), .B2(n_740), .Y(n_110) );
NOR2xp33_ASAP7_75t_L g111 ( .A(n_112), .B(n_115), .Y(n_111) );
INVx1_ASAP7_75t_L g112 ( .A(n_113), .Y(n_112) );
INVx1_ASAP7_75t_L g113 ( .A(n_114), .Y(n_113) );
INVx2_ASAP7_75t_L g739 ( .A(n_114), .Y(n_739) );
AOI21xp5_ASAP7_75t_L g740 ( .A1(n_115), .A2(n_118), .B(n_741), .Y(n_740) );
NOR2xp33_ASAP7_75t_SL g115 ( .A(n_116), .B(n_122), .Y(n_115) );
INVx1_ASAP7_75t_SL g116 ( .A(n_117), .Y(n_116) );
INVx1_ASAP7_75t_SL g117 ( .A(n_118), .Y(n_117) );
NOR2x2_ASAP7_75t_L g737 ( .A(n_119), .B(n_729), .Y(n_737) );
INVx2_ASAP7_75t_L g119 ( .A(n_120), .Y(n_119) );
OR2x2_ASAP7_75t_L g728 ( .A(n_120), .B(n_729), .Y(n_728) );
OAI22xp5_ASAP7_75t_SL g124 ( .A1(n_125), .A2(n_450), .B1(n_453), .B2(n_726), .Y(n_124) );
INVx1_ASAP7_75t_L g125 ( .A(n_126), .Y(n_125) );
BUFx2_ASAP7_75t_L g733 ( .A(n_126), .Y(n_733) );
AND3x1_ASAP7_75t_L g126 ( .A(n_127), .B(n_354), .C(n_411), .Y(n_126) );
NOR3xp33_ASAP7_75t_L g127 ( .A(n_128), .B(n_299), .C(n_335), .Y(n_127) );
OAI211xp5_ASAP7_75t_L g128 ( .A1(n_129), .A2(n_201), .B(n_253), .C(n_286), .Y(n_128) );
NAND2xp5_ASAP7_75t_L g129 ( .A(n_130), .B(n_165), .Y(n_129) );
HB1xp67_ASAP7_75t_L g130 ( .A(n_131), .Y(n_130) );
AND2x4_ASAP7_75t_L g256 ( .A(n_131), .B(n_257), .Y(n_256) );
INVx5_ASAP7_75t_L g285 ( .A(n_131), .Y(n_285) );
AND2x2_ASAP7_75t_L g358 ( .A(n_131), .B(n_274), .Y(n_358) );
AND2x2_ASAP7_75t_L g396 ( .A(n_131), .B(n_302), .Y(n_396) );
AND2x2_ASAP7_75t_L g416 ( .A(n_131), .B(n_258), .Y(n_416) );
OR2x6_ASAP7_75t_L g131 ( .A(n_132), .B(n_162), .Y(n_131) );
AOI21xp5_ASAP7_75t_SL g132 ( .A1(n_133), .A2(n_142), .B(n_155), .Y(n_132) );
BUFx2_ASAP7_75t_L g134 ( .A(n_135), .Y(n_134) );
AND2x4_ASAP7_75t_L g135 ( .A(n_136), .B(n_140), .Y(n_135) );
NAND2x1p5_ASAP7_75t_L g222 ( .A(n_136), .B(n_140), .Y(n_222) );
AND2x2_ASAP7_75t_L g136 ( .A(n_137), .B(n_139), .Y(n_136) );
INVx1_ASAP7_75t_L g153 ( .A(n_137), .Y(n_153) );
INVx1_ASAP7_75t_L g137 ( .A(n_138), .Y(n_137) );
INVx2_ASAP7_75t_L g144 ( .A(n_138), .Y(n_144) );
INVx1_ASAP7_75t_L g216 ( .A(n_138), .Y(n_216) );
INVx1_ASAP7_75t_L g145 ( .A(n_139), .Y(n_145) );
BUFx6f_ASAP7_75t_L g149 ( .A(n_139), .Y(n_149) );
INVx3_ASAP7_75t_L g180 ( .A(n_139), .Y(n_180) );
INVx1_ASAP7_75t_L g212 ( .A(n_139), .Y(n_212) );
BUFx6f_ASAP7_75t_L g227 ( .A(n_139), .Y(n_227) );
BUFx3_ASAP7_75t_L g154 ( .A(n_140), .Y(n_154) );
INVx4_ASAP7_75t_SL g184 ( .A(n_140), .Y(n_184) );
INVx5_ASAP7_75t_L g193 ( .A(n_143), .Y(n_193) );
AND2x6_ASAP7_75t_L g143 ( .A(n_144), .B(n_145), .Y(n_143) );
BUFx6f_ASAP7_75t_L g182 ( .A(n_144), .Y(n_182) );
BUFx3_ASAP7_75t_L g198 ( .A(n_144), .Y(n_198) );
AOI21xp5_ASAP7_75t_L g146 ( .A1(n_147), .A2(n_150), .B(n_152), .Y(n_146) );
INVx2_ASAP7_75t_L g151 ( .A(n_148), .Y(n_151) );
INVx2_ASAP7_75t_L g148 ( .A(n_149), .Y(n_148) );
INVx4_ASAP7_75t_L g177 ( .A(n_149), .Y(n_177) );
O2A1O1Ixp33_ASAP7_75t_L g194 ( .A1(n_151), .A2(n_195), .B(n_196), .C(n_197), .Y(n_194) );
O2A1O1Ixp33_ASAP7_75t_L g236 ( .A1(n_151), .A2(n_197), .B(n_237), .C(n_238), .Y(n_236) );
O2A1O1Ixp5_ASAP7_75t_L g523 ( .A1(n_151), .A2(n_524), .B(n_525), .C(n_526), .Y(n_523) );
O2A1O1Ixp33_ASAP7_75t_L g540 ( .A1(n_151), .A2(n_526), .B(n_541), .C(n_542), .Y(n_540) );
O2A1O1Ixp33_ASAP7_75t_L g462 ( .A1(n_152), .A2(n_179), .B(n_463), .C(n_464), .Y(n_462) );
INVx2_ASAP7_75t_L g152 ( .A(n_153), .Y(n_152) );
NAND2xp5_ASAP7_75t_SL g477 ( .A(n_153), .B(n_478), .Y(n_477) );
INVx1_ASAP7_75t_L g155 ( .A(n_156), .Y(n_155) );
NOR2xp33_ASAP7_75t_L g543 ( .A(n_156), .B(n_544), .Y(n_543) );
INVx2_ASAP7_75t_L g156 ( .A(n_157), .Y(n_156) );
INVx1_ASAP7_75t_L g164 ( .A(n_157), .Y(n_164) );
AOI21xp5_ASAP7_75t_L g189 ( .A1(n_157), .A2(n_190), .B(n_191), .Y(n_189) );
AOI21xp5_ASAP7_75t_L g233 ( .A1(n_157), .A2(n_234), .B(n_235), .Y(n_233) );
O2A1O1Ixp33_ASAP7_75t_L g459 ( .A1(n_157), .A2(n_222), .B(n_460), .C(n_461), .Y(n_459) );
OA21x2_ASAP7_75t_L g484 ( .A1(n_157), .A2(n_485), .B(n_492), .Y(n_484) );
AND2x2_ASAP7_75t_SL g157 ( .A(n_158), .B(n_159), .Y(n_157) );
AND2x2_ASAP7_75t_L g171 ( .A(n_158), .B(n_159), .Y(n_171) );
NAND2xp5_ASAP7_75t_L g159 ( .A(n_160), .B(n_161), .Y(n_159) );
NOR2xp33_ASAP7_75t_L g162 ( .A(n_163), .B(n_164), .Y(n_162) );
AO21x2_ASAP7_75t_L g519 ( .A1(n_164), .A2(n_520), .B(n_527), .Y(n_519) );
NAND2xp5_ASAP7_75t_L g288 ( .A(n_165), .B(n_289), .Y(n_288) );
AND2x2_ASAP7_75t_L g165 ( .A(n_166), .B(n_188), .Y(n_165) );
HB1xp67_ASAP7_75t_L g297 ( .A(n_166), .Y(n_297) );
AND2x2_ASAP7_75t_L g311 ( .A(n_166), .B(n_257), .Y(n_311) );
INVx1_ASAP7_75t_L g334 ( .A(n_166), .Y(n_334) );
NAND2xp5_ASAP7_75t_L g373 ( .A(n_166), .B(n_285), .Y(n_373) );
OR2x2_ASAP7_75t_L g410 ( .A(n_166), .B(n_255), .Y(n_410) );
INVx2_ASAP7_75t_L g166 ( .A(n_167), .Y(n_166) );
HB1xp67_ASAP7_75t_L g346 ( .A(n_167), .Y(n_346) );
AND2x2_ASAP7_75t_L g353 ( .A(n_167), .B(n_258), .Y(n_353) );
INVx2_ASAP7_75t_L g167 ( .A(n_168), .Y(n_167) );
AND2x2_ASAP7_75t_L g274 ( .A(n_168), .B(n_258), .Y(n_274) );
BUFx2_ASAP7_75t_L g302 ( .A(n_168), .Y(n_302) );
AO21x2_ASAP7_75t_L g168 ( .A1(n_169), .A2(n_172), .B(n_186), .Y(n_168) );
NOR2xp33_ASAP7_75t_L g186 ( .A(n_169), .B(n_187), .Y(n_186) );
NOR2xp33_ASAP7_75t_L g199 ( .A(n_169), .B(n_200), .Y(n_199) );
AO21x2_ASAP7_75t_L g219 ( .A1(n_169), .A2(n_220), .B(n_228), .Y(n_219) );
INVx3_ASAP7_75t_L g251 ( .A(n_169), .Y(n_251) );
NOR2xp33_ASAP7_75t_L g465 ( .A(n_169), .B(n_466), .Y(n_465) );
NOR2xp33_ASAP7_75t_L g527 ( .A(n_169), .B(n_528), .Y(n_527) );
AO21x2_ASAP7_75t_L g536 ( .A1(n_169), .A2(n_537), .B(n_543), .Y(n_536) );
INVx4_ASAP7_75t_L g169 ( .A(n_170), .Y(n_169) );
AOI21xp5_ASAP7_75t_L g207 ( .A1(n_170), .A2(n_208), .B(n_209), .Y(n_207) );
HB1xp67_ASAP7_75t_L g243 ( .A(n_170), .Y(n_243) );
BUFx6f_ASAP7_75t_L g170 ( .A(n_171), .Y(n_170) );
INVx1_ASAP7_75t_L g230 ( .A(n_171), .Y(n_230) );
NAND2xp5_ASAP7_75t_L g172 ( .A(n_173), .B(n_185), .Y(n_172) );
O2A1O1Ixp33_ASAP7_75t_L g174 ( .A1(n_175), .A2(n_176), .B(n_178), .C(n_181), .Y(n_174) );
INVx1_ASAP7_75t_L g176 ( .A(n_177), .Y(n_176) );
OAI22xp33_ASAP7_75t_L g478 ( .A1(n_177), .A2(n_179), .B1(n_479), .B2(n_480), .Y(n_478) );
NOR2xp33_ASAP7_75t_L g499 ( .A(n_177), .B(n_500), .Y(n_499) );
NOR2xp33_ASAP7_75t_L g509 ( .A(n_177), .B(n_510), .Y(n_509) );
NOR2xp33_ASAP7_75t_L g248 ( .A(n_179), .B(n_249), .Y(n_248) );
INVx2_ASAP7_75t_L g263 ( .A(n_179), .Y(n_263) );
INVx5_ASAP7_75t_L g179 ( .A(n_180), .Y(n_179) );
NOR2xp33_ASAP7_75t_L g490 ( .A(n_180), .B(n_491), .Y(n_490) );
HB1xp67_ASAP7_75t_L g181 ( .A(n_182), .Y(n_181) );
INVx3_ASAP7_75t_L g552 ( .A(n_182), .Y(n_552) );
INVx1_ASAP7_75t_L g183 ( .A(n_184), .Y(n_183) );
O2A1O1Ixp33_ASAP7_75t_L g245 ( .A1(n_184), .A2(n_193), .B(n_246), .C(n_247), .Y(n_245) );
O2A1O1Ixp33_ASAP7_75t_SL g260 ( .A1(n_184), .A2(n_193), .B(n_261), .C(n_262), .Y(n_260) );
O2A1O1Ixp33_ASAP7_75t_SL g475 ( .A1(n_184), .A2(n_193), .B(n_476), .C(n_477), .Y(n_475) );
O2A1O1Ixp33_ASAP7_75t_SL g486 ( .A1(n_184), .A2(n_193), .B(n_487), .C(n_488), .Y(n_486) );
O2A1O1Ixp33_ASAP7_75t_SL g496 ( .A1(n_184), .A2(n_193), .B(n_497), .C(n_498), .Y(n_496) );
O2A1O1Ixp33_ASAP7_75t_SL g506 ( .A1(n_184), .A2(n_193), .B(n_507), .C(n_508), .Y(n_506) );
O2A1O1Ixp33_ASAP7_75t_L g547 ( .A1(n_184), .A2(n_193), .B(n_548), .C(n_549), .Y(n_547) );
INVx5_ASAP7_75t_L g255 ( .A(n_188), .Y(n_255) );
BUFx2_ASAP7_75t_L g278 ( .A(n_188), .Y(n_278) );
AND2x2_ASAP7_75t_L g435 ( .A(n_188), .B(n_289), .Y(n_435) );
OR2x6_ASAP7_75t_L g188 ( .A(n_189), .B(n_199), .Y(n_188) );
INVx2_ASAP7_75t_L g192 ( .A(n_193), .Y(n_192) );
HB1xp67_ASAP7_75t_L g197 ( .A(n_198), .Y(n_197) );
INVx2_ASAP7_75t_L g267 ( .A(n_198), .Y(n_267) );
INVx1_ASAP7_75t_L g511 ( .A(n_198), .Y(n_511) );
INVx1_ASAP7_75t_L g201 ( .A(n_202), .Y(n_201) );
NAND2xp33_ASAP7_75t_L g202 ( .A(n_203), .B(n_240), .Y(n_202) );
OAI221xp5_ASAP7_75t_L g335 ( .A1(n_203), .A2(n_336), .B1(n_343), .B2(n_344), .C(n_347), .Y(n_335) );
OR2x2_ASAP7_75t_L g203 ( .A(n_204), .B(n_217), .Y(n_203) );
AND2x2_ASAP7_75t_L g241 ( .A(n_204), .B(n_242), .Y(n_241) );
NAND2xp5_ASAP7_75t_L g329 ( .A(n_204), .B(n_330), .Y(n_329) );
INVx1_ASAP7_75t_SL g204 ( .A(n_205), .Y(n_204) );
AND2x2_ASAP7_75t_L g270 ( .A(n_205), .B(n_218), .Y(n_270) );
NAND2xp5_ASAP7_75t_SL g280 ( .A(n_205), .B(n_219), .Y(n_280) );
OR2x2_ASAP7_75t_L g291 ( .A(n_205), .B(n_242), .Y(n_291) );
AND2x2_ASAP7_75t_L g294 ( .A(n_205), .B(n_282), .Y(n_294) );
AND2x2_ASAP7_75t_L g310 ( .A(n_205), .B(n_231), .Y(n_310) );
OR2x2_ASAP7_75t_L g326 ( .A(n_205), .B(n_219), .Y(n_326) );
NAND2xp5_ASAP7_75t_L g388 ( .A(n_205), .B(n_242), .Y(n_388) );
INVx2_ASAP7_75t_L g205 ( .A(n_206), .Y(n_205) );
NAND2xp5_ASAP7_75t_L g380 ( .A(n_206), .B(n_231), .Y(n_380) );
AND2x2_ASAP7_75t_L g383 ( .A(n_206), .B(n_219), .Y(n_383) );
AOI21xp5_ASAP7_75t_L g210 ( .A1(n_211), .A2(n_213), .B(n_214), .Y(n_210) );
AOI21xp5_ASAP7_75t_L g224 ( .A1(n_214), .A2(n_225), .B(n_226), .Y(n_224) );
INVx2_ASAP7_75t_L g214 ( .A(n_215), .Y(n_214) );
INVx3_ASAP7_75t_L g215 ( .A(n_216), .Y(n_215) );
OR2x2_ASAP7_75t_L g304 ( .A(n_217), .B(n_291), .Y(n_304) );
INVx2_ASAP7_75t_L g330 ( .A(n_217), .Y(n_330) );
OR2x2_ASAP7_75t_L g217 ( .A(n_218), .B(n_231), .Y(n_217) );
AND2x2_ASAP7_75t_L g252 ( .A(n_218), .B(n_232), .Y(n_252) );
NAND2xp5_ASAP7_75t_L g309 ( .A(n_218), .B(n_242), .Y(n_309) );
OR2x2_ASAP7_75t_L g320 ( .A(n_218), .B(n_232), .Y(n_320) );
NAND2xp5_ASAP7_75t_L g379 ( .A(n_218), .B(n_282), .Y(n_379) );
OAI221xp5_ASAP7_75t_L g412 ( .A1(n_218), .A2(n_413), .B1(n_415), .B2(n_417), .C(n_420), .Y(n_412) );
INVx5_ASAP7_75t_SL g218 ( .A(n_219), .Y(n_218) );
NAND2xp5_ASAP7_75t_L g351 ( .A(n_219), .B(n_242), .Y(n_351) );
OAI21xp5_ASAP7_75t_L g220 ( .A1(n_221), .A2(n_222), .B(n_223), .Y(n_220) );
OAI21xp5_ASAP7_75t_L g520 ( .A1(n_222), .A2(n_521), .B(n_522), .Y(n_520) );
OAI21xp5_ASAP7_75t_L g537 ( .A1(n_222), .A2(n_538), .B(n_539), .Y(n_537) );
INVx4_ASAP7_75t_L g266 ( .A(n_227), .Y(n_266) );
INVx2_ASAP7_75t_L g489 ( .A(n_227), .Y(n_489) );
NOR2xp33_ASAP7_75t_L g228 ( .A(n_229), .B(n_230), .Y(n_228) );
INVx2_ASAP7_75t_L g472 ( .A(n_230), .Y(n_472) );
NAND2xp5_ASAP7_75t_L g281 ( .A(n_231), .B(n_282), .Y(n_281) );
NOR2xp33_ASAP7_75t_L g292 ( .A(n_231), .B(n_293), .Y(n_292) );
AND2x2_ASAP7_75t_L g298 ( .A(n_231), .B(n_270), .Y(n_298) );
OR2x2_ASAP7_75t_L g342 ( .A(n_231), .B(n_242), .Y(n_342) );
NAND2xp5_ASAP7_75t_L g361 ( .A(n_231), .B(n_294), .Y(n_361) );
NAND2xp5_ASAP7_75t_L g386 ( .A(n_231), .B(n_387), .Y(n_386) );
AND2x2_ASAP7_75t_L g407 ( .A(n_231), .B(n_408), .Y(n_407) );
INVx5_ASAP7_75t_SL g231 ( .A(n_232), .Y(n_231) );
AND2x2_ASAP7_75t_SL g271 ( .A(n_232), .B(n_241), .Y(n_271) );
O2A1O1Ixp33_ASAP7_75t_SL g275 ( .A1(n_232), .A2(n_276), .B(n_279), .C(n_283), .Y(n_275) );
OR2x2_ASAP7_75t_L g313 ( .A(n_232), .B(n_309), .Y(n_313) );
OR2x2_ASAP7_75t_L g349 ( .A(n_232), .B(n_291), .Y(n_349) );
OAI311xp33_ASAP7_75t_L g355 ( .A1(n_232), .A2(n_294), .A3(n_356), .B1(n_359), .C1(n_366), .Y(n_355) );
AND2x2_ASAP7_75t_L g406 ( .A(n_232), .B(n_242), .Y(n_406) );
AND2x2_ASAP7_75t_L g414 ( .A(n_232), .B(n_269), .Y(n_414) );
HB1xp67_ASAP7_75t_L g432 ( .A(n_232), .Y(n_432) );
AND2x2_ASAP7_75t_L g449 ( .A(n_232), .B(n_270), .Y(n_449) );
OR2x6_ASAP7_75t_L g232 ( .A(n_233), .B(n_239), .Y(n_232) );
NAND2xp5_ASAP7_75t_L g240 ( .A(n_241), .B(n_252), .Y(n_240) );
AND2x2_ASAP7_75t_L g277 ( .A(n_241), .B(n_278), .Y(n_277) );
INVx2_ASAP7_75t_L g433 ( .A(n_241), .Y(n_433) );
AND2x2_ASAP7_75t_L g269 ( .A(n_242), .B(n_270), .Y(n_269) );
INVx3_ASAP7_75t_L g282 ( .A(n_242), .Y(n_282) );
HB1xp67_ASAP7_75t_L g325 ( .A(n_242), .Y(n_325) );
INVxp67_ASAP7_75t_L g364 ( .A(n_242), .Y(n_364) );
OA21x2_ASAP7_75t_L g242 ( .A1(n_243), .A2(n_244), .B(n_250), .Y(n_242) );
OA21x2_ASAP7_75t_L g494 ( .A1(n_243), .A2(n_495), .B(n_501), .Y(n_494) );
OA21x2_ASAP7_75t_L g504 ( .A1(n_243), .A2(n_505), .B(n_512), .Y(n_504) );
OA21x2_ASAP7_75t_L g545 ( .A1(n_243), .A2(n_546), .B(n_553), .Y(n_545) );
OA21x2_ASAP7_75t_L g258 ( .A1(n_251), .A2(n_259), .B(n_268), .Y(n_258) );
AND2x2_ASAP7_75t_L g442 ( .A(n_252), .B(n_290), .Y(n_442) );
AOI221xp5_ASAP7_75t_L g253 ( .A1(n_254), .A2(n_269), .B1(n_271), .B2(n_272), .C(n_275), .Y(n_253) );
AND2x2_ASAP7_75t_L g254 ( .A(n_255), .B(n_256), .Y(n_254) );
NAND2xp5_ASAP7_75t_L g273 ( .A(n_255), .B(n_274), .Y(n_273) );
AND2x2_ASAP7_75t_L g295 ( .A(n_255), .B(n_285), .Y(n_295) );
AND2x2_ASAP7_75t_L g303 ( .A(n_255), .B(n_257), .Y(n_303) );
OR2x2_ASAP7_75t_L g315 ( .A(n_255), .B(n_316), .Y(n_315) );
AND2x2_ASAP7_75t_L g333 ( .A(n_255), .B(n_334), .Y(n_333) );
AND2x2_ASAP7_75t_L g357 ( .A(n_255), .B(n_358), .Y(n_357) );
HB1xp67_ASAP7_75t_L g377 ( .A(n_255), .Y(n_377) );
AND2x2_ASAP7_75t_L g429 ( .A(n_255), .B(n_353), .Y(n_429) );
OAI31xp33_ASAP7_75t_L g437 ( .A1(n_255), .A2(n_306), .A3(n_405), .B(n_438), .Y(n_437) );
NAND2xp5_ASAP7_75t_L g332 ( .A(n_256), .B(n_333), .Y(n_332) );
INVx1_ASAP7_75t_SL g401 ( .A(n_256), .Y(n_401) );
NOR2xp33_ASAP7_75t_L g409 ( .A(n_256), .B(n_410), .Y(n_409) );
AND2x4_ASAP7_75t_L g289 ( .A(n_257), .B(n_285), .Y(n_289) );
INVx1_ASAP7_75t_L g376 ( .A(n_257), .Y(n_376) );
INVx2_ASAP7_75t_L g257 ( .A(n_258), .Y(n_257) );
AND2x2_ASAP7_75t_L g426 ( .A(n_258), .B(n_285), .Y(n_426) );
NOR2xp33_ASAP7_75t_L g264 ( .A(n_265), .B(n_266), .Y(n_264) );
NOR2xp33_ASAP7_75t_L g550 ( .A(n_266), .B(n_551), .Y(n_550) );
INVx2_ASAP7_75t_L g526 ( .A(n_267), .Y(n_526) );
INVx1_ASAP7_75t_SL g436 ( .A(n_269), .Y(n_436) );
NAND2xp5_ASAP7_75t_L g340 ( .A(n_270), .B(n_341), .Y(n_340) );
AOI22xp5_ASAP7_75t_L g420 ( .A1(n_271), .A2(n_383), .B1(n_421), .B2(n_424), .Y(n_420) );
INVx1_ASAP7_75t_L g272 ( .A(n_273), .Y(n_272) );
AND2x2_ASAP7_75t_L g284 ( .A(n_274), .B(n_285), .Y(n_284) );
INVx1_ASAP7_75t_L g343 ( .A(n_274), .Y(n_343) );
NAND2xp5_ASAP7_75t_L g448 ( .A(n_274), .B(n_295), .Y(n_448) );
INVx1_ASAP7_75t_SL g276 ( .A(n_277), .Y(n_276) );
AND2x2_ASAP7_75t_L g418 ( .A(n_277), .B(n_419), .Y(n_418) );
AOI21xp5_ASAP7_75t_L g336 ( .A1(n_278), .A2(n_337), .B(n_339), .Y(n_336) );
OR2x2_ASAP7_75t_L g344 ( .A(n_278), .B(n_345), .Y(n_344) );
AND2x2_ASAP7_75t_L g365 ( .A(n_278), .B(n_353), .Y(n_365) );
NAND2xp5_ASAP7_75t_L g404 ( .A(n_278), .B(n_376), .Y(n_404) );
NAND2xp5_ASAP7_75t_L g415 ( .A(n_278), .B(n_416), .Y(n_415) );
OAI221xp5_ASAP7_75t_SL g392 ( .A1(n_279), .A2(n_393), .B1(n_398), .B2(n_401), .C(n_402), .Y(n_392) );
OR2x2_ASAP7_75t_L g279 ( .A(n_280), .B(n_281), .Y(n_279) );
OR2x2_ASAP7_75t_L g369 ( .A(n_280), .B(n_342), .Y(n_369) );
INVx1_ASAP7_75t_L g408 ( .A(n_280), .Y(n_408) );
INVx2_ASAP7_75t_L g384 ( .A(n_281), .Y(n_384) );
INVx1_ASAP7_75t_L g318 ( .A(n_282), .Y(n_318) );
INVx1_ASAP7_75t_SL g283 ( .A(n_284), .Y(n_283) );
INVx2_ASAP7_75t_L g323 ( .A(n_285), .Y(n_323) );
NAND2xp5_ASAP7_75t_L g345 ( .A(n_285), .B(n_346), .Y(n_345) );
AND2x2_ASAP7_75t_L g352 ( .A(n_285), .B(n_353), .Y(n_352) );
OR2x2_ASAP7_75t_L g440 ( .A(n_285), .B(n_410), .Y(n_440) );
AOI222xp33_ASAP7_75t_L g286 ( .A1(n_287), .A2(n_290), .B1(n_292), .B2(n_295), .C1(n_296), .C2(n_298), .Y(n_286) );
INVxp67_ASAP7_75t_L g287 ( .A(n_288), .Y(n_287) );
AND2x2_ASAP7_75t_L g296 ( .A(n_289), .B(n_297), .Y(n_296) );
AOI22xp33_ASAP7_75t_L g366 ( .A1(n_289), .A2(n_339), .B1(n_367), .B2(n_368), .Y(n_366) );
NAND2xp5_ASAP7_75t_L g422 ( .A(n_289), .B(n_423), .Y(n_422) );
INVx1_ASAP7_75t_SL g290 ( .A(n_291), .Y(n_290) );
INVx1_ASAP7_75t_SL g293 ( .A(n_294), .Y(n_293) );
OAI21xp33_ASAP7_75t_SL g327 ( .A1(n_298), .A2(n_328), .B(n_331), .Y(n_327) );
OAI211xp5_ASAP7_75t_SL g299 ( .A1(n_300), .A2(n_304), .B(n_305), .C(n_327), .Y(n_299) );
INVxp67_ASAP7_75t_L g300 ( .A(n_301), .Y(n_300) );
AND2x2_ASAP7_75t_L g301 ( .A(n_302), .B(n_303), .Y(n_301) );
AOI221xp5_ASAP7_75t_L g305 ( .A1(n_303), .A2(n_306), .B1(n_311), .B2(n_312), .C(n_314), .Y(n_305) );
NAND2xp5_ASAP7_75t_L g390 ( .A(n_303), .B(n_391), .Y(n_390) );
INVxp67_ASAP7_75t_L g397 ( .A(n_303), .Y(n_397) );
INVx1_ASAP7_75t_L g306 ( .A(n_307), .Y(n_306) );
NAND2xp5_ASAP7_75t_L g307 ( .A(n_308), .B(n_310), .Y(n_307) );
AND2x2_ASAP7_75t_L g399 ( .A(n_308), .B(n_400), .Y(n_399) );
INVx1_ASAP7_75t_SL g308 ( .A(n_309), .Y(n_308) );
INVx1_ASAP7_75t_L g316 ( .A(n_311), .Y(n_316) );
AND2x2_ASAP7_75t_L g322 ( .A(n_311), .B(n_323), .Y(n_322) );
INVx1_ASAP7_75t_L g312 ( .A(n_313), .Y(n_312) );
OAI22xp5_ASAP7_75t_L g314 ( .A1(n_315), .A2(n_317), .B1(n_321), .B2(n_324), .Y(n_314) );
NAND2xp5_ASAP7_75t_L g317 ( .A(n_318), .B(n_319), .Y(n_317) );
NAND2xp5_ASAP7_75t_L g338 ( .A(n_318), .B(n_330), .Y(n_338) );
NAND2xp5_ASAP7_75t_L g363 ( .A(n_319), .B(n_364), .Y(n_363) );
INVx1_ASAP7_75t_SL g319 ( .A(n_320), .Y(n_319) );
INVx1_ASAP7_75t_L g321 ( .A(n_322), .Y(n_321) );
INVx1_ASAP7_75t_L g419 ( .A(n_323), .Y(n_419) );
AND2x2_ASAP7_75t_L g438 ( .A(n_323), .B(n_353), .Y(n_438) );
OR2x2_ASAP7_75t_L g324 ( .A(n_325), .B(n_326), .Y(n_324) );
INVx1_ASAP7_75t_L g328 ( .A(n_329), .Y(n_328) );
NAND2xp5_ASAP7_75t_L g446 ( .A(n_330), .B(n_387), .Y(n_446) );
INVx1_ASAP7_75t_L g331 ( .A(n_332), .Y(n_331) );
NOR2xp33_ASAP7_75t_L g444 ( .A(n_333), .B(n_401), .Y(n_444) );
INVx1_ASAP7_75t_L g337 ( .A(n_338), .Y(n_337) );
INVx1_ASAP7_75t_L g339 ( .A(n_340), .Y(n_339) );
INVx1_ASAP7_75t_L g341 ( .A(n_342), .Y(n_341) );
INVx1_ASAP7_75t_L g367 ( .A(n_345), .Y(n_367) );
BUFx2_ASAP7_75t_L g391 ( .A(n_346), .Y(n_391) );
OAI21xp5_ASAP7_75t_SL g347 ( .A1(n_348), .A2(n_350), .B(n_352), .Y(n_347) );
INVx1_ASAP7_75t_L g348 ( .A(n_349), .Y(n_348) );
INVx1_ASAP7_75t_L g350 ( .A(n_351), .Y(n_350) );
NOR3xp33_ASAP7_75t_L g354 ( .A(n_355), .B(n_370), .C(n_392), .Y(n_354) );
INVx1_ASAP7_75t_L g356 ( .A(n_357), .Y(n_356) );
OAI21xp5_ASAP7_75t_L g359 ( .A1(n_360), .A2(n_362), .B(n_365), .Y(n_359) );
INVx1_ASAP7_75t_L g360 ( .A(n_361), .Y(n_360) );
INVx1_ASAP7_75t_L g362 ( .A(n_363), .Y(n_362) );
INVx1_ASAP7_75t_SL g368 ( .A(n_369), .Y(n_368) );
A2O1A1Ixp33_ASAP7_75t_SL g370 ( .A1(n_371), .A2(n_374), .B(n_378), .C(n_381), .Y(n_370) );
NAND2xp5_ASAP7_75t_SL g403 ( .A(n_371), .B(n_404), .Y(n_403) );
INVx1_ASAP7_75t_L g371 ( .A(n_372), .Y(n_371) );
INVx1_ASAP7_75t_L g372 ( .A(n_373), .Y(n_372) );
INVx1_ASAP7_75t_L g374 ( .A(n_375), .Y(n_374) );
NOR2xp67_ASAP7_75t_SL g375 ( .A(n_376), .B(n_377), .Y(n_375) );
OR2x2_ASAP7_75t_L g378 ( .A(n_379), .B(n_380), .Y(n_378) );
INVx1_ASAP7_75t_SL g400 ( .A(n_380), .Y(n_400) );
OAI21xp5_ASAP7_75t_L g381 ( .A1(n_382), .A2(n_385), .B(n_389), .Y(n_381) );
AND2x4_ASAP7_75t_L g382 ( .A(n_383), .B(n_384), .Y(n_382) );
AND2x2_ASAP7_75t_L g405 ( .A(n_383), .B(n_406), .Y(n_405) );
INVx1_ASAP7_75t_L g385 ( .A(n_386), .Y(n_385) );
INVx1_ASAP7_75t_SL g387 ( .A(n_388), .Y(n_387) );
INVx1_ASAP7_75t_L g389 ( .A(n_390), .Y(n_389) );
INVx1_ASAP7_75t_L g393 ( .A(n_394), .Y(n_393) );
NOR2xp33_ASAP7_75t_L g394 ( .A(n_395), .B(n_397), .Y(n_394) );
INVx2_ASAP7_75t_L g395 ( .A(n_396), .Y(n_395) );
INVx1_ASAP7_75t_L g398 ( .A(n_399), .Y(n_398) );
AOI22xp33_ASAP7_75t_L g402 ( .A1(n_403), .A2(n_405), .B1(n_407), .B2(n_409), .Y(n_402) );
INVx2_ASAP7_75t_SL g423 ( .A(n_410), .Y(n_423) );
NOR3xp33_ASAP7_75t_L g411 ( .A(n_412), .B(n_427), .C(n_439), .Y(n_411) );
INVx1_ASAP7_75t_L g413 ( .A(n_414), .Y(n_413) );
INVxp67_ASAP7_75t_L g417 ( .A(n_418), .Y(n_417) );
INVxp67_ASAP7_75t_L g421 ( .A(n_422), .Y(n_421) );
NAND2xp5_ASAP7_75t_L g425 ( .A(n_423), .B(n_426), .Y(n_425) );
INVx1_ASAP7_75t_L g424 ( .A(n_425), .Y(n_424) );
OAI221xp5_ASAP7_75t_L g427 ( .A1(n_428), .A2(n_430), .B1(n_434), .B2(n_436), .C(n_437), .Y(n_427) );
A2O1A1Ixp33_ASAP7_75t_L g439 ( .A1(n_428), .A2(n_440), .B(n_441), .C(n_443), .Y(n_439) );
INVx1_ASAP7_75t_SL g428 ( .A(n_429), .Y(n_428) );
INVxp67_ASAP7_75t_L g430 ( .A(n_431), .Y(n_430) );
NOR2xp33_ASAP7_75t_L g431 ( .A(n_432), .B(n_433), .Y(n_431) );
INVx1_ASAP7_75t_L g434 ( .A(n_435), .Y(n_434) );
INVx1_ASAP7_75t_L g441 ( .A(n_442), .Y(n_441) );
AOI22xp5_ASAP7_75t_L g443 ( .A1(n_444), .A2(n_445), .B1(n_447), .B2(n_449), .Y(n_443) );
INVx1_ASAP7_75t_L g445 ( .A(n_446), .Y(n_445) );
INVx1_ASAP7_75t_L g447 ( .A(n_448), .Y(n_447) );
INVx2_ASAP7_75t_L g450 ( .A(n_451), .Y(n_450) );
INVx2_ASAP7_75t_L g732 ( .A(n_451), .Y(n_732) );
INVx1_ASAP7_75t_L g451 ( .A(n_452), .Y(n_451) );
INVx1_ASAP7_75t_SL g734 ( .A(n_453), .Y(n_734) );
OR5x1_ASAP7_75t_L g453 ( .A(n_454), .B(n_620), .C(n_684), .D(n_700), .E(n_715), .Y(n_453) );
NAND4xp25_ASAP7_75t_L g454 ( .A(n_455), .B(n_554), .C(n_581), .D(n_604), .Y(n_454) );
AOI21xp5_ASAP7_75t_L g455 ( .A1(n_456), .A2(n_502), .B(n_513), .Y(n_455) );
NOR2xp33_ASAP7_75t_L g456 ( .A(n_457), .B(n_467), .Y(n_456) );
HB1xp67_ASAP7_75t_L g457 ( .A(n_458), .Y(n_457) );
INVx3_ASAP7_75t_SL g533 ( .A(n_458), .Y(n_533) );
AND2x4_ASAP7_75t_L g567 ( .A(n_458), .B(n_556), .Y(n_567) );
OR2x2_ASAP7_75t_L g577 ( .A(n_458), .B(n_535), .Y(n_577) );
OR2x2_ASAP7_75t_L g623 ( .A(n_458), .B(n_470), .Y(n_623) );
AND2x2_ASAP7_75t_L g637 ( .A(n_458), .B(n_534), .Y(n_637) );
AND2x2_ASAP7_75t_L g680 ( .A(n_458), .B(n_570), .Y(n_680) );
AND2x2_ASAP7_75t_L g687 ( .A(n_458), .B(n_545), .Y(n_687) );
AND2x2_ASAP7_75t_L g706 ( .A(n_458), .B(n_596), .Y(n_706) );
AND2x2_ASAP7_75t_L g724 ( .A(n_458), .B(n_566), .Y(n_724) );
OR2x6_ASAP7_75t_L g458 ( .A(n_459), .B(n_465), .Y(n_458) );
INVx1_ASAP7_75t_L g689 ( .A(n_467), .Y(n_689) );
NAND2xp5_ASAP7_75t_L g467 ( .A(n_468), .B(n_483), .Y(n_467) );
AND2x2_ASAP7_75t_L g599 ( .A(n_468), .B(n_534), .Y(n_599) );
NAND2xp5_ASAP7_75t_L g618 ( .A(n_468), .B(n_619), .Y(n_618) );
AOI32xp33_ASAP7_75t_L g632 ( .A1(n_468), .A2(n_633), .A3(n_636), .B1(n_638), .B2(n_642), .Y(n_632) );
AND2x2_ASAP7_75t_L g702 ( .A(n_468), .B(n_596), .Y(n_702) );
INVx2_ASAP7_75t_L g468 ( .A(n_469), .Y(n_468) );
INVx1_ASAP7_75t_SL g469 ( .A(n_470), .Y(n_469) );
AND2x2_ASAP7_75t_L g566 ( .A(n_470), .B(n_535), .Y(n_566) );
NAND2xp5_ASAP7_75t_L g575 ( .A(n_470), .B(n_576), .Y(n_575) );
AND2x2_ASAP7_75t_L g608 ( .A(n_470), .B(n_555), .Y(n_608) );
NAND2xp5_ASAP7_75t_L g686 ( .A(n_470), .B(n_687), .Y(n_686) );
AO21x2_ASAP7_75t_L g470 ( .A1(n_471), .A2(n_473), .B(n_481), .Y(n_470) );
INVx1_ASAP7_75t_L g571 ( .A(n_471), .Y(n_571) );
INVx1_ASAP7_75t_L g471 ( .A(n_472), .Y(n_471) );
INVx1_ASAP7_75t_L g473 ( .A(n_474), .Y(n_473) );
OA21x2_ASAP7_75t_L g570 ( .A1(n_474), .A2(n_482), .B(n_571), .Y(n_570) );
INVx1_ASAP7_75t_L g481 ( .A(n_482), .Y(n_481) );
AND2x2_ASAP7_75t_L g573 ( .A(n_483), .B(n_517), .Y(n_573) );
AND2x2_ASAP7_75t_L g649 ( .A(n_483), .B(n_650), .Y(n_649) );
INVx1_ASAP7_75t_SL g721 ( .A(n_483), .Y(n_721) );
AND2x2_ASAP7_75t_L g483 ( .A(n_484), .B(n_493), .Y(n_483) );
OR2x2_ASAP7_75t_L g516 ( .A(n_484), .B(n_494), .Y(n_516) );
AND2x2_ASAP7_75t_L g530 ( .A(n_484), .B(n_531), .Y(n_530) );
NOR2xp33_ASAP7_75t_L g558 ( .A(n_484), .B(n_559), .Y(n_558) );
INVx2_ASAP7_75t_L g580 ( .A(n_484), .Y(n_580) );
AND2x2_ASAP7_75t_L g607 ( .A(n_484), .B(n_494), .Y(n_607) );
BUFx3_ASAP7_75t_L g610 ( .A(n_484), .Y(n_610) );
NAND2xp5_ASAP7_75t_L g617 ( .A(n_484), .B(n_585), .Y(n_617) );
NAND2xp5_ASAP7_75t_L g703 ( .A(n_484), .B(n_704), .Y(n_703) );
INVx2_ASAP7_75t_L g561 ( .A(n_493), .Y(n_561) );
AND2x2_ASAP7_75t_L g579 ( .A(n_493), .B(n_559), .Y(n_579) );
INVx2_ASAP7_75t_L g493 ( .A(n_494), .Y(n_493) );
AND2x2_ASAP7_75t_L g590 ( .A(n_494), .B(n_504), .Y(n_590) );
HB1xp67_ASAP7_75t_L g603 ( .A(n_494), .Y(n_603) );
INVx1_ASAP7_75t_L g502 ( .A(n_503), .Y(n_502) );
NAND2xp5_ASAP7_75t_L g660 ( .A(n_503), .B(n_610), .Y(n_660) );
HB1xp67_ASAP7_75t_L g503 ( .A(n_504), .Y(n_503) );
INVx1_ASAP7_75t_SL g531 ( .A(n_504), .Y(n_531) );
NAND3xp33_ASAP7_75t_L g578 ( .A(n_504), .B(n_579), .C(n_580), .Y(n_578) );
OR2x2_ASAP7_75t_L g586 ( .A(n_504), .B(n_559), .Y(n_586) );
AND2x2_ASAP7_75t_L g606 ( .A(n_504), .B(n_559), .Y(n_606) );
AND2x2_ASAP7_75t_L g650 ( .A(n_504), .B(n_519), .Y(n_650) );
AOI21xp5_ASAP7_75t_L g513 ( .A1(n_514), .A2(n_529), .B(n_532), .Y(n_513) );
NAND2xp5_ASAP7_75t_SL g514 ( .A(n_515), .B(n_517), .Y(n_514) );
AND2x2_ASAP7_75t_L g725 ( .A(n_515), .B(n_650), .Y(n_725) );
INVx1_ASAP7_75t_L g515 ( .A(n_516), .Y(n_515) );
OAI22xp5_ASAP7_75t_L g664 ( .A1(n_516), .A2(n_623), .B1(n_665), .B2(n_667), .Y(n_664) );
OR2x2_ASAP7_75t_L g671 ( .A(n_516), .B(n_586), .Y(n_671) );
OR2x2_ASAP7_75t_L g695 ( .A(n_516), .B(n_696), .Y(n_695) );
NOR2xp33_ASAP7_75t_L g708 ( .A(n_516), .B(n_615), .Y(n_708) );
AND2x2_ASAP7_75t_L g601 ( .A(n_517), .B(n_602), .Y(n_601) );
AOI21xp5_ASAP7_75t_L g688 ( .A1(n_517), .A2(n_674), .B(n_689), .Y(n_688) );
AOI32xp33_ASAP7_75t_L g709 ( .A1(n_517), .A2(n_599), .A3(n_710), .B1(n_712), .B2(n_713), .Y(n_709) );
OR2x2_ASAP7_75t_L g720 ( .A(n_517), .B(n_721), .Y(n_720) );
CKINVDCx16_ASAP7_75t_R g517 ( .A(n_518), .Y(n_517) );
OR2x2_ASAP7_75t_L g588 ( .A(n_518), .B(n_589), .Y(n_588) );
NAND2xp5_ASAP7_75t_L g667 ( .A(n_518), .B(n_602), .Y(n_667) );
BUFx3_ASAP7_75t_L g518 ( .A(n_519), .Y(n_518) );
INVx4_ASAP7_75t_L g559 ( .A(n_519), .Y(n_559) );
AND2x2_ASAP7_75t_L g625 ( .A(n_519), .B(n_590), .Y(n_625) );
AND3x2_ASAP7_75t_L g634 ( .A(n_519), .B(n_530), .C(n_635), .Y(n_634) );
INVx1_ASAP7_75t_L g529 ( .A(n_530), .Y(n_529) );
AND2x2_ASAP7_75t_L g560 ( .A(n_531), .B(n_561), .Y(n_560) );
HB1xp67_ASAP7_75t_L g615 ( .A(n_531), .Y(n_615) );
NAND2xp5_ASAP7_75t_L g696 ( .A(n_531), .B(n_559), .Y(n_696) );
NAND2xp5_ASAP7_75t_L g532 ( .A(n_533), .B(n_534), .Y(n_532) );
AND2x2_ASAP7_75t_L g555 ( .A(n_533), .B(n_556), .Y(n_555) );
AND2x2_ASAP7_75t_L g595 ( .A(n_533), .B(n_596), .Y(n_595) );
AND2x2_ASAP7_75t_L g613 ( .A(n_533), .B(n_545), .Y(n_613) );
AND2x2_ASAP7_75t_L g631 ( .A(n_533), .B(n_535), .Y(n_631) );
OR2x2_ASAP7_75t_L g645 ( .A(n_533), .B(n_646), .Y(n_645) );
AND2x2_ASAP7_75t_L g691 ( .A(n_533), .B(n_619), .Y(n_691) );
NAND2xp5_ASAP7_75t_L g569 ( .A(n_534), .B(n_570), .Y(n_569) );
AND2x2_ASAP7_75t_L g534 ( .A(n_535), .B(n_545), .Y(n_534) );
AND2x2_ASAP7_75t_L g592 ( .A(n_535), .B(n_570), .Y(n_592) );
OR2x2_ASAP7_75t_L g646 ( .A(n_535), .B(n_570), .Y(n_646) );
AND2x2_ASAP7_75t_L g699 ( .A(n_535), .B(n_556), .Y(n_699) );
INVx2_ASAP7_75t_SL g535 ( .A(n_536), .Y(n_535) );
BUFx2_ASAP7_75t_L g597 ( .A(n_536), .Y(n_597) );
AND2x2_ASAP7_75t_L g619 ( .A(n_536), .B(n_545), .Y(n_619) );
INVx2_ASAP7_75t_L g556 ( .A(n_545), .Y(n_556) );
INVx1_ASAP7_75t_L g576 ( .A(n_545), .Y(n_576) );
AOI211xp5_ASAP7_75t_L g554 ( .A1(n_555), .A2(n_557), .B(n_562), .C(n_574), .Y(n_554) );
NAND2xp5_ASAP7_75t_L g665 ( .A(n_555), .B(n_666), .Y(n_665) );
INVx1_ASAP7_75t_L g718 ( .A(n_555), .Y(n_718) );
AND2x2_ASAP7_75t_L g596 ( .A(n_556), .B(n_597), .Y(n_596) );
AND2x2_ASAP7_75t_L g557 ( .A(n_558), .B(n_560), .Y(n_557) );
NAND2xp5_ASAP7_75t_L g568 ( .A(n_559), .B(n_560), .Y(n_568) );
INVx1_ASAP7_75t_L g653 ( .A(n_559), .Y(n_653) );
NAND2xp5_ASAP7_75t_L g677 ( .A(n_559), .B(n_580), .Y(n_677) );
AND2x2_ASAP7_75t_L g693 ( .A(n_559), .B(n_607), .Y(n_693) );
NAND2xp5_ASAP7_75t_SL g675 ( .A(n_560), .B(n_676), .Y(n_675) );
INVx2_ASAP7_75t_L g584 ( .A(n_561), .Y(n_584) );
OAI22xp5_ASAP7_75t_L g562 ( .A1(n_563), .A2(n_568), .B1(n_569), .B2(n_572), .Y(n_562) );
INVx1_ASAP7_75t_L g563 ( .A(n_564), .Y(n_563) );
NOR2xp33_ASAP7_75t_L g564 ( .A(n_565), .B(n_567), .Y(n_564) );
NOR2xp33_ASAP7_75t_L g717 ( .A(n_565), .B(n_718), .Y(n_717) );
INVx1_ASAP7_75t_L g565 ( .A(n_566), .Y(n_565) );
NAND2xp5_ASAP7_75t_L g612 ( .A(n_566), .B(n_613), .Y(n_612) );
AND2x2_ASAP7_75t_L g591 ( .A(n_567), .B(n_592), .Y(n_591) );
AOI221xp5_ASAP7_75t_SL g656 ( .A1(n_567), .A2(n_609), .B1(n_657), .B2(n_662), .C(n_664), .Y(n_656) );
NAND2xp5_ASAP7_75t_L g663 ( .A(n_567), .B(n_630), .Y(n_663) );
INVx1_ASAP7_75t_L g723 ( .A(n_569), .Y(n_723) );
BUFx3_ASAP7_75t_L g630 ( .A(n_570), .Y(n_630) );
INVx1_ASAP7_75t_L g572 ( .A(n_573), .Y(n_572) );
AOI21xp33_ASAP7_75t_SL g574 ( .A1(n_575), .A2(n_577), .B(n_578), .Y(n_574) );
INVx1_ASAP7_75t_L g639 ( .A(n_576), .Y(n_639) );
NAND2xp5_ASAP7_75t_L g683 ( .A(n_576), .B(n_630), .Y(n_683) );
INVx1_ASAP7_75t_L g640 ( .A(n_577), .Y(n_640) );
NAND2xp5_ASAP7_75t_SL g641 ( .A(n_577), .B(n_630), .Y(n_641) );
INVxp67_ASAP7_75t_L g661 ( .A(n_579), .Y(n_661) );
AND2x2_ASAP7_75t_L g602 ( .A(n_580), .B(n_603), .Y(n_602) );
O2A1O1Ixp33_ASAP7_75t_L g581 ( .A1(n_582), .A2(n_587), .B(n_591), .C(n_593), .Y(n_581) );
INVx1_ASAP7_75t_L g582 ( .A(n_583), .Y(n_582) );
NAND2xp5_ASAP7_75t_L g583 ( .A(n_584), .B(n_585), .Y(n_583) );
INVx1_ASAP7_75t_SL g616 ( .A(n_584), .Y(n_616) );
NAND2xp5_ASAP7_75t_L g627 ( .A(n_585), .B(n_616), .Y(n_627) );
NAND2xp5_ASAP7_75t_L g658 ( .A(n_585), .B(n_607), .Y(n_658) );
INVx2_ASAP7_75t_SL g585 ( .A(n_586), .Y(n_585) );
INVx1_ASAP7_75t_L g587 ( .A(n_588), .Y(n_587) );
OAI22xp5_ASAP7_75t_L g593 ( .A1(n_588), .A2(n_594), .B1(n_598), .B2(n_600), .Y(n_593) );
INVx1_ASAP7_75t_SL g589 ( .A(n_590), .Y(n_589) );
AND2x2_ASAP7_75t_L g609 ( .A(n_590), .B(n_610), .Y(n_609) );
AND2x2_ASAP7_75t_L g654 ( .A(n_590), .B(n_655), .Y(n_654) );
OAI21xp33_ASAP7_75t_L g657 ( .A1(n_592), .A2(n_658), .B(n_659), .Y(n_657) );
INVx1_ASAP7_75t_SL g594 ( .A(n_595), .Y(n_594) );
AOI221xp5_ASAP7_75t_L g604 ( .A1(n_596), .A2(n_605), .B1(n_608), .B2(n_609), .C(n_611), .Y(n_604) );
NAND2xp5_ASAP7_75t_L g673 ( .A(n_596), .B(n_630), .Y(n_673) );
NAND2xp5_ASAP7_75t_L g679 ( .A(n_596), .B(n_680), .Y(n_679) );
INVx1_ASAP7_75t_L g598 ( .A(n_599), .Y(n_598) );
INVx1_ASAP7_75t_L g600 ( .A(n_601), .Y(n_600) );
INVx1_ASAP7_75t_L g712 ( .A(n_602), .Y(n_712) );
INVxp67_ASAP7_75t_L g635 ( .A(n_603), .Y(n_635) );
INVx1_ASAP7_75t_L g642 ( .A(n_605), .Y(n_642) );
AND2x2_ASAP7_75t_L g605 ( .A(n_606), .B(n_607), .Y(n_605) );
AND2x2_ASAP7_75t_L g681 ( .A(n_606), .B(n_610), .Y(n_681) );
INVx1_ASAP7_75t_L g655 ( .A(n_610), .Y(n_655) );
NAND2xp5_ASAP7_75t_SL g685 ( .A(n_610), .B(n_625), .Y(n_685) );
OAI32xp33_ASAP7_75t_L g611 ( .A1(n_612), .A2(n_614), .A3(n_616), .B1(n_617), .B2(n_618), .Y(n_611) );
INVx1_ASAP7_75t_L g614 ( .A(n_615), .Y(n_614) );
INVx2_ASAP7_75t_SL g624 ( .A(n_619), .Y(n_624) );
NAND2xp5_ASAP7_75t_L g668 ( .A(n_619), .B(n_651), .Y(n_668) );
NAND2xp5_ASAP7_75t_L g711 ( .A(n_619), .B(n_680), .Y(n_711) );
NAND2x1p5_ASAP7_75t_L g719 ( .A(n_619), .B(n_630), .Y(n_719) );
NAND5xp2_ASAP7_75t_L g620 ( .A(n_621), .B(n_643), .C(n_656), .D(n_668), .E(n_669), .Y(n_620) );
AOI221xp5_ASAP7_75t_L g621 ( .A1(n_622), .A2(n_625), .B1(n_626), .B2(n_628), .C(n_632), .Y(n_621) );
NOR2xp33_ASAP7_75t_L g622 ( .A(n_623), .B(n_624), .Y(n_622) );
INVx1_ASAP7_75t_L g626 ( .A(n_627), .Y(n_626) );
NAND2xp33_ASAP7_75t_SL g647 ( .A(n_627), .B(n_648), .Y(n_647) );
INVx1_ASAP7_75t_L g628 ( .A(n_629), .Y(n_628) );
NAND2xp5_ASAP7_75t_L g629 ( .A(n_630), .B(n_631), .Y(n_629) );
NAND2xp5_ASAP7_75t_L g698 ( .A(n_630), .B(n_699), .Y(n_698) );
AOI22xp33_ASAP7_75t_L g643 ( .A1(n_631), .A2(n_644), .B1(n_647), .B2(n_651), .Y(n_643) );
INVx2_ASAP7_75t_SL g633 ( .A(n_634), .Y(n_633) );
OAI211xp5_ASAP7_75t_SL g638 ( .A1(n_634), .A2(n_639), .B(n_640), .C(n_641), .Y(n_638) );
INVx1_ASAP7_75t_L g636 ( .A(n_637), .Y(n_636) );
INVx1_ASAP7_75t_L g644 ( .A(n_645), .Y(n_644) );
INVx1_ASAP7_75t_SL g666 ( .A(n_646), .Y(n_666) );
INVx1_ASAP7_75t_SL g648 ( .A(n_649), .Y(n_648) );
INVx1_ASAP7_75t_SL g651 ( .A(n_652), .Y(n_651) );
NAND2xp5_ASAP7_75t_L g652 ( .A(n_653), .B(n_654), .Y(n_652) );
NAND2xp5_ASAP7_75t_L g714 ( .A(n_655), .B(n_704), .Y(n_714) );
OR2x2_ASAP7_75t_L g659 ( .A(n_660), .B(n_661), .Y(n_659) );
INVx1_ASAP7_75t_L g662 ( .A(n_663), .Y(n_662) );
AOI222xp33_ASAP7_75t_L g669 ( .A1(n_670), .A2(n_672), .B1(n_674), .B2(n_678), .C1(n_681), .C2(n_682), .Y(n_669) );
INVx1_ASAP7_75t_L g670 ( .A(n_671), .Y(n_670) );
INVx1_ASAP7_75t_L g672 ( .A(n_673), .Y(n_672) );
INVx1_ASAP7_75t_L g674 ( .A(n_675), .Y(n_674) );
INVx1_ASAP7_75t_L g676 ( .A(n_677), .Y(n_676) );
INVx1_ASAP7_75t_L g678 ( .A(n_679), .Y(n_678) );
INVx1_ASAP7_75t_L g682 ( .A(n_683), .Y(n_682) );
OAI221xp5_ASAP7_75t_L g684 ( .A1(n_685), .A2(n_686), .B1(n_688), .B2(n_690), .C(n_692), .Y(n_684) );
INVx1_ASAP7_75t_SL g690 ( .A(n_691), .Y(n_690) );
OAI21xp33_ASAP7_75t_L g692 ( .A1(n_693), .A2(n_694), .B(n_697), .Y(n_692) );
INVx2_ASAP7_75t_L g694 ( .A(n_695), .Y(n_694) );
INVx1_ASAP7_75t_L g704 ( .A(n_696), .Y(n_704) );
INVx1_ASAP7_75t_L g697 ( .A(n_698), .Y(n_697) );
OAI221xp5_ASAP7_75t_L g700 ( .A1(n_701), .A2(n_703), .B1(n_705), .B2(n_707), .C(n_709), .Y(n_700) );
INVx1_ASAP7_75t_L g701 ( .A(n_702), .Y(n_701) );
INVx1_ASAP7_75t_SL g705 ( .A(n_706), .Y(n_705) );
INVxp67_ASAP7_75t_L g707 ( .A(n_708), .Y(n_707) );
INVx1_ASAP7_75t_L g710 ( .A(n_711), .Y(n_710) );
INVx1_ASAP7_75t_L g713 ( .A(n_714), .Y(n_713) );
A2O1A1Ixp33_ASAP7_75t_L g715 ( .A1(n_716), .A2(n_719), .B(n_720), .C(n_722), .Y(n_715) );
INVxp67_ASAP7_75t_L g716 ( .A(n_717), .Y(n_716) );
OAI21xp33_ASAP7_75t_L g722 ( .A1(n_723), .A2(n_724), .B(n_725), .Y(n_722) );
INVx2_ASAP7_75t_L g726 ( .A(n_727), .Y(n_726) );
INVx1_ASAP7_75t_L g727 ( .A(n_728), .Y(n_727) );
OAI22xp5_ASAP7_75t_L g731 ( .A1(n_728), .A2(n_732), .B1(n_733), .B2(n_734), .Y(n_731) );
INVx1_ASAP7_75t_SL g735 ( .A(n_736), .Y(n_735) );
INVx2_ASAP7_75t_L g736 ( .A(n_737), .Y(n_736) );
INVx2_ASAP7_75t_SL g738 ( .A(n_739), .Y(n_738) );
endmodule