module fake_jpeg_19674_n_175 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_175);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_175;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_21;
wire n_57;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_24;
wire n_44;
wire n_143;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_161;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_36;
wire n_62;
wire n_167;
wire n_174;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

HB1xp67_ASAP7_75t_L g15 ( 
.A(n_4),
.Y(n_15)
);

BUFx16f_ASAP7_75t_L g16 ( 
.A(n_4),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_0),
.Y(n_17)
);

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_8),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_12),
.Y(n_19)
);

BUFx12_ASAP7_75t_L g20 ( 
.A(n_14),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_1),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_10),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_2),
.Y(n_23)
);

INVx5_ASAP7_75t_L g24 ( 
.A(n_10),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_0),
.Y(n_25)
);

INVx3_ASAP7_75t_L g26 ( 
.A(n_13),
.Y(n_26)
);

BUFx5_ASAP7_75t_L g27 ( 
.A(n_11),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_11),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_9),
.Y(n_29)
);

INVxp67_ASAP7_75t_L g30 ( 
.A(n_8),
.Y(n_30)
);

INVx3_ASAP7_75t_L g31 ( 
.A(n_20),
.Y(n_31)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_31),
.B(n_34),
.Y(n_48)
);

BUFx3_ASAP7_75t_L g32 ( 
.A(n_16),
.Y(n_32)
);

BUFx3_ASAP7_75t_L g55 ( 
.A(n_32),
.Y(n_55)
);

BUFx12f_ASAP7_75t_L g33 ( 
.A(n_18),
.Y(n_33)
);

INVx5_ASAP7_75t_L g54 ( 
.A(n_33),
.Y(n_54)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_17),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_17),
.Y(n_35)
);

NAND2xp5_ASAP7_75t_SL g51 ( 
.A(n_35),
.B(n_36),
.Y(n_51)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_15),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g37 ( 
.A(n_16),
.B(n_20),
.Y(n_37)
);

OR2x2_ASAP7_75t_L g52 ( 
.A(n_37),
.B(n_40),
.Y(n_52)
);

INVx4_ASAP7_75t_L g38 ( 
.A(n_27),
.Y(n_38)
);

INVx3_ASAP7_75t_L g53 ( 
.A(n_38),
.Y(n_53)
);

INVx5_ASAP7_75t_L g39 ( 
.A(n_18),
.Y(n_39)
);

INVx6_ASAP7_75t_L g43 ( 
.A(n_39),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g40 ( 
.A(n_16),
.B(n_0),
.Y(n_40)
);

AOI22xp33_ASAP7_75t_SL g41 ( 
.A1(n_38),
.A2(n_24),
.B1(n_26),
.B2(n_25),
.Y(n_41)
);

AOI22xp5_ASAP7_75t_SL g58 ( 
.A1(n_41),
.A2(n_44),
.B1(n_39),
.B2(n_24),
.Y(n_58)
);

AND2x2_ASAP7_75t_L g42 ( 
.A(n_37),
.B(n_16),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_SL g75 ( 
.A(n_42),
.B(n_21),
.Y(n_75)
);

AOI22xp33_ASAP7_75t_SL g44 ( 
.A1(n_38),
.A2(n_24),
.B1(n_26),
.B2(n_25),
.Y(n_44)
);

OR2x4_ASAP7_75t_L g45 ( 
.A(n_34),
.B(n_23),
.Y(n_45)
);

AND2x2_ASAP7_75t_L g72 ( 
.A(n_45),
.B(n_23),
.Y(n_72)
);

INVx11_ASAP7_75t_L g46 ( 
.A(n_33),
.Y(n_46)
);

INVx4_ASAP7_75t_L g74 ( 
.A(n_46),
.Y(n_74)
);

BUFx5_ASAP7_75t_L g47 ( 
.A(n_32),
.Y(n_47)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_47),
.Y(n_60)
);

BUFx12_ASAP7_75t_L g49 ( 
.A(n_32),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_49),
.B(n_54),
.Y(n_56)
);

HB1xp67_ASAP7_75t_L g50 ( 
.A(n_39),
.Y(n_50)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_50),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_56),
.B(n_75),
.Y(n_89)
);

BUFx2_ASAP7_75t_L g57 ( 
.A(n_46),
.Y(n_57)
);

INVx2_ASAP7_75t_L g92 ( 
.A(n_57),
.Y(n_92)
);

OAI22xp5_ASAP7_75t_L g79 ( 
.A1(n_58),
.A2(n_61),
.B1(n_22),
.B2(n_53),
.Y(n_79)
);

CKINVDCx16_ASAP7_75t_R g59 ( 
.A(n_55),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_SL g83 ( 
.A(n_59),
.B(n_66),
.Y(n_83)
);

OAI22xp5_ASAP7_75t_SL g61 ( 
.A1(n_52),
.A2(n_36),
.B1(n_35),
.B2(n_40),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_L g62 ( 
.A(n_51),
.B(n_33),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_L g81 ( 
.A(n_62),
.B(n_69),
.Y(n_81)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_54),
.Y(n_63)
);

BUFx2_ASAP7_75t_L g95 ( 
.A(n_63),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_48),
.B(n_19),
.Y(n_64)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_64),
.Y(n_85)
);

OAI21xp33_ASAP7_75t_SL g65 ( 
.A1(n_52),
.A2(n_20),
.B(n_15),
.Y(n_65)
);

NAND3xp33_ASAP7_75t_L g77 ( 
.A(n_65),
.B(n_69),
.C(n_62),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_45),
.B(n_21),
.Y(n_66)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_50),
.Y(n_68)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_68),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_L g69 ( 
.A(n_51),
.B(n_52),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_48),
.B(n_45),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_SL g96 ( 
.A(n_70),
.B(n_71),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_42),
.B(n_19),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_L g88 ( 
.A(n_72),
.B(n_73),
.Y(n_88)
);

OAI32xp33_ASAP7_75t_L g73 ( 
.A1(n_42),
.A2(n_22),
.A3(n_20),
.B1(n_30),
.B2(n_27),
.Y(n_73)
);

MAJIxp5_ASAP7_75t_L g76 ( 
.A(n_53),
.B(n_33),
.C(n_31),
.Y(n_76)
);

XNOR2xp5_ASAP7_75t_L g78 ( 
.A(n_76),
.B(n_46),
.Y(n_78)
);

OAI21xp5_ASAP7_75t_L g111 ( 
.A1(n_77),
.A2(n_28),
.B(n_29),
.Y(n_111)
);

AND2x2_ASAP7_75t_L g108 ( 
.A(n_78),
.B(n_79),
.Y(n_108)
);

XNOR2xp5_ASAP7_75t_L g80 ( 
.A(n_61),
.B(n_49),
.Y(n_80)
);

MAJIxp5_ASAP7_75t_L g102 ( 
.A(n_80),
.B(n_60),
.C(n_59),
.Y(n_102)
);

CKINVDCx20_ASAP7_75t_R g82 ( 
.A(n_67),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_SL g114 ( 
.A(n_82),
.B(n_91),
.Y(n_114)
);

AOI21xp5_ASAP7_75t_L g84 ( 
.A1(n_72),
.A2(n_49),
.B(n_54),
.Y(n_84)
);

OAI21xp5_ASAP7_75t_SL g107 ( 
.A1(n_84),
.A2(n_90),
.B(n_93),
.Y(n_107)
);

OAI32xp33_ASAP7_75t_L g87 ( 
.A1(n_66),
.A2(n_28),
.A3(n_18),
.B1(n_29),
.B2(n_43),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_L g97 ( 
.A(n_87),
.B(n_58),
.Y(n_97)
);

AND2x2_ASAP7_75t_L g90 ( 
.A(n_76),
.B(n_73),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_75),
.B(n_49),
.Y(n_91)
);

AND2x2_ASAP7_75t_L g93 ( 
.A(n_72),
.B(n_43),
.Y(n_93)
);

INVx2_ASAP7_75t_L g94 ( 
.A(n_57),
.Y(n_94)
);

CKINVDCx20_ASAP7_75t_R g101 ( 
.A(n_94),
.Y(n_101)
);

OAI22xp5_ASAP7_75t_L g116 ( 
.A1(n_97),
.A2(n_100),
.B1(n_88),
.B2(n_81),
.Y(n_116)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_86),
.Y(n_98)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_98),
.Y(n_127)
);

HAxp5_ASAP7_75t_SL g99 ( 
.A(n_84),
.B(n_68),
.CON(n_99),
.SN(n_99)
);

NOR3xp33_ASAP7_75t_L g118 ( 
.A(n_99),
.B(n_111),
.C(n_93),
.Y(n_118)
);

OAI22xp33_ASAP7_75t_SL g100 ( 
.A1(n_87),
.A2(n_43),
.B1(n_67),
.B2(n_74),
.Y(n_100)
);

XNOR2xp5_ASAP7_75t_L g119 ( 
.A(n_102),
.B(n_80),
.Y(n_119)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_95),
.Y(n_103)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_103),
.Y(n_123)
);

INVxp67_ASAP7_75t_L g104 ( 
.A(n_89),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_SL g117 ( 
.A(n_104),
.B(n_112),
.Y(n_117)
);

AOI32xp33_ASAP7_75t_L g105 ( 
.A1(n_90),
.A2(n_74),
.A3(n_60),
.B1(n_28),
.B2(n_57),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g120 ( 
.A(n_105),
.B(n_113),
.Y(n_120)
);

AO22x1_ASAP7_75t_L g106 ( 
.A1(n_88),
.A2(n_63),
.B1(n_55),
.B2(n_47),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_L g115 ( 
.A(n_106),
.B(n_109),
.Y(n_115)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_95),
.Y(n_109)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_78),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_L g125 ( 
.A(n_110),
.B(n_55),
.Y(n_125)
);

INVx1_ASAP7_75t_SL g112 ( 
.A(n_93),
.Y(n_112)
);

CKINVDCx20_ASAP7_75t_R g113 ( 
.A(n_85),
.Y(n_113)
);

AOI22xp5_ASAP7_75t_L g139 ( 
.A1(n_116),
.A2(n_121),
.B1(n_101),
.B2(n_109),
.Y(n_139)
);

INVxp67_ASAP7_75t_L g133 ( 
.A(n_118),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_L g132 ( 
.A(n_119),
.B(n_125),
.Y(n_132)
);

OAI22xp5_ASAP7_75t_L g121 ( 
.A1(n_97),
.A2(n_81),
.B1(n_90),
.B2(n_83),
.Y(n_121)
);

INVxp67_ASAP7_75t_L g122 ( 
.A(n_114),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_SL g131 ( 
.A(n_122),
.B(n_124),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_113),
.B(n_96),
.Y(n_124)
);

AOI21xp5_ASAP7_75t_L g126 ( 
.A1(n_107),
.A2(n_94),
.B(n_92),
.Y(n_126)
);

CKINVDCx16_ASAP7_75t_R g142 ( 
.A(n_126),
.Y(n_142)
);

XNOR2xp5_ASAP7_75t_L g128 ( 
.A(n_110),
.B(n_92),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_L g134 ( 
.A(n_128),
.B(n_129),
.Y(n_134)
);

OR2x2_ASAP7_75t_L g129 ( 
.A(n_112),
.B(n_29),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_L g130 ( 
.A(n_98),
.B(n_63),
.Y(n_130)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_130),
.Y(n_136)
);

OAI321xp33_ASAP7_75t_L g135 ( 
.A1(n_115),
.A2(n_108),
.A3(n_111),
.B1(n_106),
.B2(n_107),
.C(n_104),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_SL g147 ( 
.A(n_135),
.B(n_139),
.Y(n_147)
);

OAI22xp5_ASAP7_75t_L g137 ( 
.A1(n_120),
.A2(n_108),
.B1(n_106),
.B2(n_102),
.Y(n_137)
);

AOI22xp5_ASAP7_75t_L g145 ( 
.A1(n_137),
.A2(n_140),
.B1(n_141),
.B2(n_122),
.Y(n_145)
);

AO21x1_ASAP7_75t_L g138 ( 
.A1(n_115),
.A2(n_108),
.B(n_101),
.Y(n_138)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_138),
.Y(n_143)
);

AOI22xp5_ASAP7_75t_L g140 ( 
.A1(n_117),
.A2(n_103),
.B1(n_14),
.B2(n_13),
.Y(n_140)
);

AOI22xp5_ASAP7_75t_L g141 ( 
.A1(n_119),
.A2(n_12),
.B1(n_2),
.B2(n_3),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_SL g144 ( 
.A(n_131),
.B(n_141),
.Y(n_144)
);

NOR2xp33_ASAP7_75t_SL g152 ( 
.A(n_144),
.B(n_146),
.Y(n_152)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_145),
.Y(n_153)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_136),
.Y(n_146)
);

MAJIxp5_ASAP7_75t_L g148 ( 
.A(n_132),
.B(n_128),
.C(n_125),
.Y(n_148)
);

MAJIxp5_ASAP7_75t_L g158 ( 
.A(n_148),
.B(n_149),
.C(n_151),
.Y(n_158)
);

XNOR2xp5_ASAP7_75t_L g149 ( 
.A(n_139),
.B(n_126),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_SL g150 ( 
.A(n_136),
.B(n_127),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_SL g157 ( 
.A(n_150),
.B(n_134),
.Y(n_157)
);

XOR2xp5_ASAP7_75t_L g151 ( 
.A(n_132),
.B(n_129),
.Y(n_151)
);

OAI22xp5_ASAP7_75t_SL g154 ( 
.A1(n_147),
.A2(n_142),
.B1(n_138),
.B2(n_133),
.Y(n_154)
);

AOI22xp5_ASAP7_75t_L g159 ( 
.A1(n_154),
.A2(n_149),
.B1(n_134),
.B2(n_151),
.Y(n_159)
);

OAI21xp5_ASAP7_75t_SL g155 ( 
.A1(n_143),
.A2(n_133),
.B(n_140),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_L g162 ( 
.A(n_155),
.B(n_156),
.Y(n_162)
);

HB1xp67_ASAP7_75t_L g156 ( 
.A(n_148),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_SL g161 ( 
.A(n_157),
.B(n_123),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_SL g166 ( 
.A(n_159),
.B(n_164),
.Y(n_166)
);

BUFx24_ASAP7_75t_SL g160 ( 
.A(n_152),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_L g165 ( 
.A(n_160),
.B(n_161),
.Y(n_165)
);

AOI22xp5_ASAP7_75t_SL g163 ( 
.A1(n_153),
.A2(n_123),
.B1(n_2),
.B2(n_3),
.Y(n_163)
);

AOI22xp5_ASAP7_75t_SL g167 ( 
.A1(n_163),
.A2(n_158),
.B1(n_154),
.B2(n_5),
.Y(n_167)
);

MAJIxp5_ASAP7_75t_L g164 ( 
.A(n_158),
.B(n_1),
.C(n_3),
.Y(n_164)
);

MAJIxp5_ASAP7_75t_L g171 ( 
.A(n_167),
.B(n_6),
.C(n_7),
.Y(n_171)
);

OAI221xp5_ASAP7_75t_L g168 ( 
.A1(n_162),
.A2(n_1),
.B1(n_4),
.B2(n_5),
.C(n_6),
.Y(n_168)
);

AOI21xp5_ASAP7_75t_L g169 ( 
.A1(n_168),
.A2(n_5),
.B(n_6),
.Y(n_169)
);

OAI21xp5_ASAP7_75t_L g173 ( 
.A1(n_169),
.A2(n_171),
.B(n_7),
.Y(n_173)
);

BUFx24_ASAP7_75t_SL g170 ( 
.A(n_165),
.Y(n_170)
);

NOR4xp25_ASAP7_75t_L g172 ( 
.A(n_170),
.B(n_166),
.C(n_8),
.D(n_9),
.Y(n_172)
);

OAI21xp5_ASAP7_75t_L g174 ( 
.A1(n_172),
.A2(n_173),
.B(n_7),
.Y(n_174)
);

XNOR2xp5_ASAP7_75t_L g175 ( 
.A(n_174),
.B(n_9),
.Y(n_175)
);


endmodule