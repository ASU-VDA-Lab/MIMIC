module fake_jpeg_14188_n_562 (n_13, n_1, n_10, n_6, n_14, n_18, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_562);

input n_13;
input n_1;
input n_10;
input n_6;
input n_14;
input n_18;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_562;

wire n_529;
wire n_390;
wire n_552;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_525;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_519;
wire n_276;
wire n_143;
wire n_431;
wire n_102;
wire n_549;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_172;
wire n_547;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_513;
wire n_283;
wire n_107;
wire n_490;
wire n_517;
wire n_415;
wire n_479;
wire n_543;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_542;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_559;
wire n_48;
wire n_465;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_221;
wire n_256;
wire n_454;
wire n_540;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_508;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_544;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_530;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_557;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_298;
wire n_106;
wire n_545;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_474;
wire n_539;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_511;
wire n_486;
wire n_305;
wire n_161;
wire n_441;
wire n_555;
wire n_342;
wire n_101;
wire n_226;
wire n_509;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_560;
wire n_190;
wire n_510;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_536;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_537;
wire n_110;
wire n_531;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_554;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_523;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_533;
wire n_296;
wire n_384;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_491;
wire n_24;
wire n_526;
wire n_467;
wire n_269;
wire n_546;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_473;
wire n_45;
wire n_520;
wire n_476;
wire n_337;
wire n_317;
wire n_145;
wire n_20;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_481;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_522;
wire n_333;
wire n_518;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_302;
wire n_216;
wire n_528;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_199;
wire n_260;
wire n_550;
wire n_413;
wire n_275;
wire n_494;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_551;
wire n_36;
wire n_62;
wire n_492;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_515;
wire n_347;
wire n_521;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_538;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_534;
wire n_472;
wire n_279;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_484;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_469;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_553;
wire n_257;
wire n_61;
wire n_173;
wire n_561;
wire n_244;
wire n_232;
wire n_527;
wire n_482;
wire n_58;
wire n_41;
wire n_266;
wire n_548;
wire n_72;
wire n_512;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_516;
wire n_183;
wire n_409;
wire n_532;
wire n_249;
wire n_412;
wire n_217;
wire n_471;
wire n_541;
wire n_53;
wire n_372;
wire n_558;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_535;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_556;
wire n_524;
wire n_402;
wire n_504;
wire n_438;
wire n_475;
wire n_247;
wire n_157;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_514;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

INVx1_ASAP7_75t_L g19 ( 
.A(n_6),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_14),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_7),
.Y(n_21)
);

BUFx4f_ASAP7_75t_L g22 ( 
.A(n_7),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_16),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_9),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_18),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_9),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_6),
.Y(n_27)
);

INVx11_ASAP7_75t_L g28 ( 
.A(n_11),
.Y(n_28)
);

BUFx5_ASAP7_75t_L g29 ( 
.A(n_14),
.Y(n_29)
);

INVx2_ASAP7_75t_L g30 ( 
.A(n_15),
.Y(n_30)
);

BUFx3_ASAP7_75t_L g31 ( 
.A(n_10),
.Y(n_31)
);

INVx2_ASAP7_75t_L g32 ( 
.A(n_11),
.Y(n_32)
);

BUFx8_ASAP7_75t_L g33 ( 
.A(n_9),
.Y(n_33)
);

INVx1_ASAP7_75t_SL g34 ( 
.A(n_1),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_2),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g36 ( 
.A(n_10),
.B(n_8),
.Y(n_36)
);

BUFx10_ASAP7_75t_L g37 ( 
.A(n_17),
.Y(n_37)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_16),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_2),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_4),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_18),
.Y(n_41)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_1),
.Y(n_42)
);

BUFx12f_ASAP7_75t_L g43 ( 
.A(n_7),
.Y(n_43)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_3),
.Y(n_44)
);

BUFx10_ASAP7_75t_L g45 ( 
.A(n_16),
.Y(n_45)
);

BUFx12f_ASAP7_75t_L g46 ( 
.A(n_13),
.Y(n_46)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_17),
.Y(n_47)
);

OR2x2_ASAP7_75t_L g48 ( 
.A(n_18),
.B(n_12),
.Y(n_48)
);

INVx6_ASAP7_75t_L g49 ( 
.A(n_15),
.Y(n_49)
);

BUFx12_ASAP7_75t_L g50 ( 
.A(n_13),
.Y(n_50)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_4),
.Y(n_51)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_4),
.Y(n_52)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_11),
.Y(n_53)
);

INVx3_ASAP7_75t_L g54 ( 
.A(n_33),
.Y(n_54)
);

INVx3_ASAP7_75t_L g123 ( 
.A(n_54),
.Y(n_123)
);

CKINVDCx20_ASAP7_75t_R g55 ( 
.A(n_50),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g155 ( 
.A(n_55),
.B(n_62),
.Y(n_155)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_53),
.Y(n_56)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_56),
.Y(n_119)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_30),
.Y(n_57)
);

INVx2_ASAP7_75t_L g111 ( 
.A(n_57),
.Y(n_111)
);

BUFx12_ASAP7_75t_L g58 ( 
.A(n_37),
.Y(n_58)
);

BUFx4f_ASAP7_75t_SL g173 ( 
.A(n_58),
.Y(n_173)
);

INVx11_ASAP7_75t_L g59 ( 
.A(n_28),
.Y(n_59)
);

BUFx10_ASAP7_75t_L g136 ( 
.A(n_59),
.Y(n_136)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_53),
.Y(n_60)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_60),
.Y(n_150)
);

BUFx3_ASAP7_75t_L g61 ( 
.A(n_43),
.Y(n_61)
);

BUFx3_ASAP7_75t_L g126 ( 
.A(n_61),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_48),
.B(n_8),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_39),
.Y(n_63)
);

BUFx6f_ASAP7_75t_L g110 ( 
.A(n_63),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_SL g64 ( 
.A(n_36),
.B(n_8),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g161 ( 
.A(n_64),
.B(n_77),
.Y(n_161)
);

INVx8_ASAP7_75t_L g65 ( 
.A(n_29),
.Y(n_65)
);

INVx5_ASAP7_75t_L g125 ( 
.A(n_65),
.Y(n_125)
);

INVx6_ASAP7_75t_L g66 ( 
.A(n_39),
.Y(n_66)
);

INVx6_ASAP7_75t_L g116 ( 
.A(n_66),
.Y(n_116)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_39),
.Y(n_67)
);

BUFx6f_ASAP7_75t_L g151 ( 
.A(n_67),
.Y(n_151)
);

BUFx16f_ASAP7_75t_L g68 ( 
.A(n_43),
.Y(n_68)
);

BUFx12f_ASAP7_75t_L g117 ( 
.A(n_68),
.Y(n_117)
);

INVx4_ASAP7_75t_L g69 ( 
.A(n_29),
.Y(n_69)
);

INVx4_ASAP7_75t_L g113 ( 
.A(n_69),
.Y(n_113)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_19),
.Y(n_70)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_70),
.Y(n_165)
);

INVx2_ASAP7_75t_L g71 ( 
.A(n_30),
.Y(n_71)
);

INVx2_ASAP7_75t_L g114 ( 
.A(n_71),
.Y(n_114)
);

INVx3_ASAP7_75t_L g72 ( 
.A(n_33),
.Y(n_72)
);

INVx3_ASAP7_75t_L g127 ( 
.A(n_72),
.Y(n_127)
);

BUFx6f_ASAP7_75t_L g73 ( 
.A(n_40),
.Y(n_73)
);

BUFx6f_ASAP7_75t_L g164 ( 
.A(n_73),
.Y(n_164)
);

BUFx6f_ASAP7_75t_L g74 ( 
.A(n_40),
.Y(n_74)
);

INVx6_ASAP7_75t_L g132 ( 
.A(n_74),
.Y(n_132)
);

INVx6_ASAP7_75t_L g75 ( 
.A(n_40),
.Y(n_75)
);

INVx6_ASAP7_75t_L g137 ( 
.A(n_75),
.Y(n_137)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_19),
.Y(n_76)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_76),
.Y(n_175)
);

OR2x2_ASAP7_75t_L g77 ( 
.A(n_48),
.B(n_6),
.Y(n_77)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_21),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g170 ( 
.A(n_78),
.B(n_87),
.Y(n_170)
);

INVx6_ASAP7_75t_SL g79 ( 
.A(n_37),
.Y(n_79)
);

NAND2x1_ASAP7_75t_SL g121 ( 
.A(n_79),
.B(n_107),
.Y(n_121)
);

INVx8_ASAP7_75t_L g80 ( 
.A(n_28),
.Y(n_80)
);

INVx5_ASAP7_75t_L g135 ( 
.A(n_80),
.Y(n_135)
);

INVx8_ASAP7_75t_L g81 ( 
.A(n_28),
.Y(n_81)
);

INVx5_ASAP7_75t_L g148 ( 
.A(n_81),
.Y(n_148)
);

BUFx6f_ASAP7_75t_L g82 ( 
.A(n_22),
.Y(n_82)
);

INVx8_ASAP7_75t_L g156 ( 
.A(n_82),
.Y(n_156)
);

INVx2_ASAP7_75t_L g83 ( 
.A(n_32),
.Y(n_83)
);

INVx2_ASAP7_75t_L g118 ( 
.A(n_83),
.Y(n_118)
);

INVx6_ASAP7_75t_L g84 ( 
.A(n_23),
.Y(n_84)
);

INVx3_ASAP7_75t_SL g120 ( 
.A(n_84),
.Y(n_120)
);

INVx2_ASAP7_75t_SL g85 ( 
.A(n_43),
.Y(n_85)
);

HB1xp67_ASAP7_75t_L g166 ( 
.A(n_85),
.Y(n_166)
);

BUFx6f_ASAP7_75t_L g86 ( 
.A(n_22),
.Y(n_86)
);

BUFx2_ASAP7_75t_L g143 ( 
.A(n_86),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_SL g87 ( 
.A(n_36),
.B(n_10),
.Y(n_87)
);

INVx2_ASAP7_75t_L g88 ( 
.A(n_32),
.Y(n_88)
);

INVx2_ASAP7_75t_L g129 ( 
.A(n_88),
.Y(n_129)
);

INVx2_ASAP7_75t_L g89 ( 
.A(n_22),
.Y(n_89)
);

INVx2_ASAP7_75t_L g139 ( 
.A(n_89),
.Y(n_139)
);

INVx2_ASAP7_75t_L g90 ( 
.A(n_22),
.Y(n_90)
);

INVx2_ASAP7_75t_L g141 ( 
.A(n_90),
.Y(n_141)
);

INVx11_ASAP7_75t_L g91 ( 
.A(n_37),
.Y(n_91)
);

CKINVDCx16_ASAP7_75t_R g115 ( 
.A(n_91),
.Y(n_115)
);

INVx2_ASAP7_75t_L g92 ( 
.A(n_35),
.Y(n_92)
);

INVx2_ASAP7_75t_L g149 ( 
.A(n_92),
.Y(n_149)
);

CKINVDCx20_ASAP7_75t_R g93 ( 
.A(n_50),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_L g130 ( 
.A(n_93),
.B(n_101),
.Y(n_130)
);

INVx2_ASAP7_75t_L g94 ( 
.A(n_35),
.Y(n_94)
);

INVx2_ASAP7_75t_L g159 ( 
.A(n_94),
.Y(n_159)
);

INVx2_ASAP7_75t_L g95 ( 
.A(n_42),
.Y(n_95)
);

INVx2_ASAP7_75t_L g162 ( 
.A(n_95),
.Y(n_162)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_21),
.Y(n_96)
);

INVx2_ASAP7_75t_SL g144 ( 
.A(n_96),
.Y(n_144)
);

INVx2_ASAP7_75t_L g97 ( 
.A(n_42),
.Y(n_97)
);

INVx2_ASAP7_75t_L g167 ( 
.A(n_97),
.Y(n_167)
);

INVx8_ASAP7_75t_L g98 ( 
.A(n_37),
.Y(n_98)
);

INVx3_ASAP7_75t_L g131 ( 
.A(n_98),
.Y(n_131)
);

BUFx6f_ASAP7_75t_L g99 ( 
.A(n_23),
.Y(n_99)
);

BUFx12f_ASAP7_75t_L g133 ( 
.A(n_99),
.Y(n_133)
);

BUFx6f_ASAP7_75t_L g100 ( 
.A(n_23),
.Y(n_100)
);

BUFx12f_ASAP7_75t_L g146 ( 
.A(n_100),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_L g101 ( 
.A(n_48),
.B(n_27),
.Y(n_101)
);

BUFx6f_ASAP7_75t_L g102 ( 
.A(n_25),
.Y(n_102)
);

BUFx12f_ASAP7_75t_L g147 ( 
.A(n_102),
.Y(n_147)
);

HB1xp67_ASAP7_75t_L g103 ( 
.A(n_37),
.Y(n_103)
);

CKINVDCx16_ASAP7_75t_R g158 ( 
.A(n_103),
.Y(n_158)
);

INVx4_ASAP7_75t_L g104 ( 
.A(n_43),
.Y(n_104)
);

INVx4_ASAP7_75t_L g122 ( 
.A(n_104),
.Y(n_122)
);

INVx3_ASAP7_75t_L g105 ( 
.A(n_33),
.Y(n_105)
);

INVx3_ASAP7_75t_L g140 ( 
.A(n_105),
.Y(n_140)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_38),
.Y(n_106)
);

INVx2_ASAP7_75t_SL g157 ( 
.A(n_106),
.Y(n_157)
);

CKINVDCx5p33_ASAP7_75t_R g107 ( 
.A(n_45),
.Y(n_107)
);

BUFx6f_ASAP7_75t_L g108 ( 
.A(n_25),
.Y(n_108)
);

INVx3_ASAP7_75t_L g142 ( 
.A(n_108),
.Y(n_142)
);

INVxp67_ASAP7_75t_L g109 ( 
.A(n_103),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_L g178 ( 
.A(n_109),
.B(n_168),
.Y(n_178)
);

AOI22xp5_ASAP7_75t_L g112 ( 
.A1(n_84),
.A2(n_49),
.B1(n_25),
.B2(n_38),
.Y(n_112)
);

OAI22xp5_ASAP7_75t_L g195 ( 
.A1(n_112),
.A2(n_134),
.B1(n_154),
.B2(n_73),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_SL g124 ( 
.A(n_62),
.B(n_26),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_SL g213 ( 
.A(n_124),
.B(n_128),
.Y(n_213)
);

NAND2xp5_ASAP7_75t_SL g128 ( 
.A(n_77),
.B(n_26),
.Y(n_128)
);

AOI22xp33_ASAP7_75t_L g134 ( 
.A1(n_99),
.A2(n_49),
.B1(n_34),
.B2(n_45),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_SL g138 ( 
.A(n_85),
.B(n_27),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_L g236 ( 
.A(n_138),
.B(n_160),
.Y(n_236)
);

INVx3_ASAP7_75t_L g145 ( 
.A(n_68),
.Y(n_145)
);

INVx1_ASAP7_75t_SL g231 ( 
.A(n_145),
.Y(n_231)
);

AOI22xp33_ASAP7_75t_SL g152 ( 
.A1(n_65),
.A2(n_34),
.B1(n_31),
.B2(n_45),
.Y(n_152)
);

AOI22xp33_ASAP7_75t_SL g192 ( 
.A1(n_152),
.A2(n_45),
.B1(n_46),
.B2(n_67),
.Y(n_192)
);

INVx4_ASAP7_75t_L g153 ( 
.A(n_61),
.Y(n_153)
);

BUFx2_ASAP7_75t_L g232 ( 
.A(n_153),
.Y(n_232)
);

AOI22xp33_ASAP7_75t_L g154 ( 
.A1(n_100),
.A2(n_49),
.B1(n_34),
.B2(n_45),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_SL g160 ( 
.A(n_66),
.B(n_20),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_L g163 ( 
.A(n_82),
.B(n_20),
.Y(n_163)
);

AND2x2_ASAP7_75t_L g184 ( 
.A(n_163),
.B(n_174),
.Y(n_184)
);

INVxp67_ASAP7_75t_L g168 ( 
.A(n_98),
.Y(n_168)
);

CKINVDCx20_ASAP7_75t_R g169 ( 
.A(n_58),
.Y(n_169)
);

NOR2xp33_ASAP7_75t_L g185 ( 
.A(n_169),
.B(n_46),
.Y(n_185)
);

INVx2_ASAP7_75t_L g171 ( 
.A(n_86),
.Y(n_171)
);

INVx2_ASAP7_75t_L g190 ( 
.A(n_171),
.Y(n_190)
);

INVx4_ASAP7_75t_L g172 ( 
.A(n_80),
.Y(n_172)
);

INVx4_ASAP7_75t_L g197 ( 
.A(n_172),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_L g174 ( 
.A(n_75),
.B(n_24),
.Y(n_174)
);

AOI22xp5_ASAP7_75t_L g176 ( 
.A1(n_111),
.A2(n_108),
.B1(n_102),
.B2(n_74),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_L g268 ( 
.A(n_176),
.B(n_137),
.Y(n_268)
);

INVx3_ASAP7_75t_L g177 ( 
.A(n_133),
.Y(n_177)
);

BUFx2_ASAP7_75t_L g243 ( 
.A(n_177),
.Y(n_243)
);

CKINVDCx14_ASAP7_75t_R g179 ( 
.A(n_121),
.Y(n_179)
);

NOR2xp33_ASAP7_75t_L g248 ( 
.A(n_179),
.B(n_210),
.Y(n_248)
);

BUFx6f_ASAP7_75t_L g180 ( 
.A(n_110),
.Y(n_180)
);

BUFx6f_ASAP7_75t_L g290 ( 
.A(n_180),
.Y(n_290)
);

INVx3_ASAP7_75t_L g181 ( 
.A(n_133),
.Y(n_181)
);

INVx3_ASAP7_75t_L g281 ( 
.A(n_181),
.Y(n_281)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_119),
.Y(n_182)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_182),
.Y(n_242)
);

INVx3_ASAP7_75t_L g183 ( 
.A(n_146),
.Y(n_183)
);

INVx3_ASAP7_75t_L g286 ( 
.A(n_183),
.Y(n_286)
);

CKINVDCx16_ASAP7_75t_R g241 ( 
.A(n_185),
.Y(n_241)
);

MAJIxp5_ASAP7_75t_L g186 ( 
.A(n_130),
.B(n_47),
.C(n_41),
.Y(n_186)
);

XOR2xp5_ASAP7_75t_L g247 ( 
.A(n_186),
.B(n_199),
.Y(n_247)
);

BUFx3_ASAP7_75t_L g187 ( 
.A(n_117),
.Y(n_187)
);

BUFx3_ASAP7_75t_L g245 ( 
.A(n_187),
.Y(n_245)
);

AND2x2_ASAP7_75t_L g188 ( 
.A(n_170),
.B(n_33),
.Y(n_188)
);

AND2x2_ASAP7_75t_L g249 ( 
.A(n_188),
.B(n_222),
.Y(n_249)
);

INVx6_ASAP7_75t_SL g189 ( 
.A(n_121),
.Y(n_189)
);

CKINVDCx20_ASAP7_75t_R g244 ( 
.A(n_189),
.Y(n_244)
);

NOR2xp33_ASAP7_75t_L g191 ( 
.A(n_155),
.B(n_41),
.Y(n_191)
);

NOR2xp33_ASAP7_75t_SL g240 ( 
.A(n_191),
.B(n_203),
.Y(n_240)
);

INVxp67_ASAP7_75t_L g250 ( 
.A(n_192),
.Y(n_250)
);

INVx6_ASAP7_75t_L g193 ( 
.A(n_132),
.Y(n_193)
);

INVx6_ASAP7_75t_L g267 ( 
.A(n_193),
.Y(n_267)
);

BUFx6f_ASAP7_75t_L g194 ( 
.A(n_151),
.Y(n_194)
);

INVx8_ASAP7_75t_L g257 ( 
.A(n_194),
.Y(n_257)
);

AOI22xp5_ASAP7_75t_L g251 ( 
.A1(n_195),
.A2(n_205),
.B1(n_207),
.B2(n_214),
.Y(n_251)
);

INVx13_ASAP7_75t_L g196 ( 
.A(n_117),
.Y(n_196)
);

INVxp67_ASAP7_75t_L g270 ( 
.A(n_196),
.Y(n_270)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_150),
.Y(n_198)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_198),
.Y(n_252)
);

MAJIxp5_ASAP7_75t_L g199 ( 
.A(n_165),
.B(n_47),
.C(n_24),
.Y(n_199)
);

CKINVDCx20_ASAP7_75t_R g200 ( 
.A(n_166),
.Y(n_200)
);

NAND2xp5_ASAP7_75t_L g279 ( 
.A(n_200),
.B(n_204),
.Y(n_279)
);

INVx6_ASAP7_75t_L g201 ( 
.A(n_164),
.Y(n_201)
);

INVx8_ASAP7_75t_L g287 ( 
.A(n_201),
.Y(n_287)
);

BUFx5_ASAP7_75t_L g202 ( 
.A(n_136),
.Y(n_202)
);

INVx3_ASAP7_75t_L g293 ( 
.A(n_202),
.Y(n_293)
);

NOR2xp33_ASAP7_75t_L g203 ( 
.A(n_155),
.B(n_46),
.Y(n_203)
);

NOR2xp33_ASAP7_75t_L g204 ( 
.A(n_128),
.B(n_46),
.Y(n_204)
);

OAI22xp33_ASAP7_75t_L g205 ( 
.A1(n_134),
.A2(n_63),
.B1(n_31),
.B2(n_51),
.Y(n_205)
);

CKINVDCx20_ASAP7_75t_R g206 ( 
.A(n_166),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_L g291 ( 
.A(n_206),
.B(n_209),
.Y(n_291)
);

OAI22xp33_ASAP7_75t_SL g207 ( 
.A1(n_152),
.A2(n_31),
.B1(n_51),
.B2(n_44),
.Y(n_207)
);

INVx2_ASAP7_75t_L g208 ( 
.A(n_139),
.Y(n_208)
);

INVx2_ASAP7_75t_L g263 ( 
.A(n_208),
.Y(n_263)
);

CKINVDCx20_ASAP7_75t_R g209 ( 
.A(n_138),
.Y(n_209)
);

CKINVDCx20_ASAP7_75t_R g210 ( 
.A(n_144),
.Y(n_210)
);

INVx4_ASAP7_75t_L g211 ( 
.A(n_146),
.Y(n_211)
);

HB1xp67_ASAP7_75t_L g255 ( 
.A(n_211),
.Y(n_255)
);

INVx4_ASAP7_75t_L g212 ( 
.A(n_147),
.Y(n_212)
);

INVx2_ASAP7_75t_L g285 ( 
.A(n_212),
.Y(n_285)
);

AOI22xp33_ASAP7_75t_L g214 ( 
.A1(n_149),
.A2(n_167),
.B1(n_162),
.B2(n_159),
.Y(n_214)
);

NOR2xp33_ASAP7_75t_L g215 ( 
.A(n_124),
.B(n_44),
.Y(n_215)
);

NAND2xp5_ASAP7_75t_SL g269 ( 
.A(n_215),
.B(n_218),
.Y(n_269)
);

CKINVDCx12_ASAP7_75t_R g216 ( 
.A(n_173),
.Y(n_216)
);

INVxp67_ASAP7_75t_L g273 ( 
.A(n_216),
.Y(n_273)
);

AO22x1_ASAP7_75t_SL g217 ( 
.A1(n_114),
.A2(n_81),
.B1(n_50),
.B2(n_52),
.Y(n_217)
);

NAND2xp5_ASAP7_75t_L g295 ( 
.A(n_217),
.B(n_235),
.Y(n_295)
);

NOR2xp33_ASAP7_75t_L g218 ( 
.A(n_170),
.B(n_52),
.Y(n_218)
);

INVx2_ASAP7_75t_L g219 ( 
.A(n_141),
.Y(n_219)
);

INVx2_ASAP7_75t_L g288 ( 
.A(n_219),
.Y(n_288)
);

BUFx3_ASAP7_75t_L g220 ( 
.A(n_126),
.Y(n_220)
);

INVx2_ASAP7_75t_L g294 ( 
.A(n_220),
.Y(n_294)
);

OAI22xp33_ASAP7_75t_SL g221 ( 
.A1(n_142),
.A2(n_50),
.B1(n_12),
.B2(n_13),
.Y(n_221)
);

AOI22xp5_ASAP7_75t_L g262 ( 
.A1(n_221),
.A2(n_127),
.B1(n_140),
.B2(n_148),
.Y(n_262)
);

AND2x2_ASAP7_75t_L g222 ( 
.A(n_161),
.B(n_5),
.Y(n_222)
);

INVx2_ASAP7_75t_L g223 ( 
.A(n_175),
.Y(n_223)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_223),
.Y(n_264)
);

INVx11_ASAP7_75t_L g224 ( 
.A(n_136),
.Y(n_224)
);

INVxp67_ASAP7_75t_L g289 ( 
.A(n_224),
.Y(n_289)
);

AND2x2_ASAP7_75t_L g225 ( 
.A(n_161),
.B(n_5),
.Y(n_225)
);

AND2x2_ASAP7_75t_L g260 ( 
.A(n_225),
.B(n_228),
.Y(n_260)
);

INVx4_ASAP7_75t_L g226 ( 
.A(n_147),
.Y(n_226)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_226),
.Y(n_265)
);

INVx4_ASAP7_75t_L g227 ( 
.A(n_131),
.Y(n_227)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_227),
.Y(n_277)
);

INVx3_ASAP7_75t_L g228 ( 
.A(n_156),
.Y(n_228)
);

BUFx2_ASAP7_75t_SL g229 ( 
.A(n_123),
.Y(n_229)
);

CKINVDCx20_ASAP7_75t_R g246 ( 
.A(n_229),
.Y(n_246)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_144),
.Y(n_230)
);

NOR2xp33_ASAP7_75t_L g253 ( 
.A(n_230),
.B(n_237),
.Y(n_253)
);

NOR2xp33_ASAP7_75t_L g233 ( 
.A(n_157),
.B(n_160),
.Y(n_233)
);

NAND2xp5_ASAP7_75t_SL g284 ( 
.A(n_233),
.B(n_15),
.Y(n_284)
);

BUFx6f_ASAP7_75t_L g234 ( 
.A(n_116),
.Y(n_234)
);

AOI22xp33_ASAP7_75t_SL g258 ( 
.A1(n_234),
.A2(n_235),
.B1(n_120),
.B2(n_143),
.Y(n_258)
);

AOI22xp33_ASAP7_75t_SL g235 ( 
.A1(n_125),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_235)
);

AND2x2_ASAP7_75t_L g237 ( 
.A(n_118),
.B(n_5),
.Y(n_237)
);

INVx2_ASAP7_75t_L g238 ( 
.A(n_157),
.Y(n_238)
);

NOR2xp33_ASAP7_75t_L g266 ( 
.A(n_238),
.B(n_239),
.Y(n_266)
);

CKINVDCx20_ASAP7_75t_R g239 ( 
.A(n_158),
.Y(n_239)
);

CKINVDCx20_ASAP7_75t_R g254 ( 
.A(n_178),
.Y(n_254)
);

NOR2xp33_ASAP7_75t_L g299 ( 
.A(n_254),
.B(n_272),
.Y(n_299)
);

AND2x4_ASAP7_75t_SL g256 ( 
.A(n_236),
.B(n_129),
.Y(n_256)
);

AND2x2_ASAP7_75t_L g298 ( 
.A(n_256),
.B(n_268),
.Y(n_298)
);

INVxp67_ASAP7_75t_L g321 ( 
.A(n_258),
.Y(n_321)
);

AOI32xp33_ASAP7_75t_L g259 ( 
.A1(n_188),
.A2(n_113),
.A3(n_154),
.B1(n_115),
.B2(n_122),
.Y(n_259)
);

OR2x2_ASAP7_75t_L g305 ( 
.A(n_259),
.B(n_197),
.Y(n_305)
);

AOI22xp33_ASAP7_75t_L g261 ( 
.A1(n_217),
.A2(n_205),
.B1(n_184),
.B2(n_207),
.Y(n_261)
);

OAI22xp5_ASAP7_75t_L g341 ( 
.A1(n_261),
.A2(n_262),
.B1(n_271),
.B2(n_278),
.Y(n_341)
);

AOI22xp33_ASAP7_75t_L g271 ( 
.A1(n_217),
.A2(n_115),
.B1(n_158),
.B2(n_135),
.Y(n_271)
);

CKINVDCx20_ASAP7_75t_R g272 ( 
.A(n_214),
.Y(n_272)
);

CKINVDCx20_ASAP7_75t_R g274 ( 
.A(n_231),
.Y(n_274)
);

NOR2xp33_ASAP7_75t_L g302 ( 
.A(n_274),
.B(n_231),
.Y(n_302)
);

NAND2xp5_ASAP7_75t_L g275 ( 
.A(n_184),
.B(n_0),
.Y(n_275)
);

NAND2xp5_ASAP7_75t_L g300 ( 
.A(n_275),
.B(n_280),
.Y(n_300)
);

NOR2xp33_ASAP7_75t_L g276 ( 
.A(n_213),
.B(n_173),
.Y(n_276)
);

NAND2xp5_ASAP7_75t_SL g323 ( 
.A(n_276),
.B(n_284),
.Y(n_323)
);

AOI22xp5_ASAP7_75t_L g278 ( 
.A1(n_221),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_278)
);

NAND2xp5_ASAP7_75t_L g280 ( 
.A(n_237),
.B(n_222),
.Y(n_280)
);

AOI22xp5_ASAP7_75t_L g282 ( 
.A1(n_192),
.A2(n_0),
.B1(n_3),
.B2(n_4),
.Y(n_282)
);

OAI22xp5_ASAP7_75t_SL g335 ( 
.A1(n_282),
.A2(n_180),
.B1(n_194),
.B2(n_193),
.Y(n_335)
);

AOI22xp33_ASAP7_75t_SL g283 ( 
.A1(n_227),
.A2(n_3),
.B1(n_12),
.B2(n_14),
.Y(n_283)
);

INVxp67_ASAP7_75t_L g331 ( 
.A(n_283),
.Y(n_331)
);

OAI21xp5_ASAP7_75t_L g292 ( 
.A1(n_225),
.A2(n_3),
.B(n_17),
.Y(n_292)
);

AOI21xp5_ASAP7_75t_L g307 ( 
.A1(n_292),
.A2(n_232),
.B(n_224),
.Y(n_307)
);

AND2x2_ASAP7_75t_L g330 ( 
.A(n_295),
.B(n_202),
.Y(n_330)
);

CKINVDCx20_ASAP7_75t_R g296 ( 
.A(n_291),
.Y(n_296)
);

NOR2xp33_ASAP7_75t_L g353 ( 
.A(n_296),
.B(n_307),
.Y(n_353)
);

INVx13_ASAP7_75t_L g297 ( 
.A(n_273),
.Y(n_297)
);

INVxp67_ASAP7_75t_L g348 ( 
.A(n_297),
.Y(n_348)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_263),
.Y(n_301)
);

INVx1_ASAP7_75t_L g345 ( 
.A(n_301),
.Y(n_345)
);

NAND2xp5_ASAP7_75t_SL g350 ( 
.A(n_302),
.B(n_309),
.Y(n_350)
);

INVx2_ASAP7_75t_L g303 ( 
.A(n_287),
.Y(n_303)
);

INVx2_ASAP7_75t_L g382 ( 
.A(n_303),
.Y(n_382)
);

NOR2xp33_ASAP7_75t_SL g304 ( 
.A(n_280),
.B(n_197),
.Y(n_304)
);

NOR2xp33_ASAP7_75t_SL g377 ( 
.A(n_304),
.B(n_306),
.Y(n_377)
);

OAI21xp5_ASAP7_75t_L g351 ( 
.A1(n_305),
.A2(n_249),
.B(n_260),
.Y(n_351)
);

NOR2xp33_ASAP7_75t_L g306 ( 
.A(n_240),
.B(n_232),
.Y(n_306)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_263),
.Y(n_308)
);

INVx1_ASAP7_75t_L g347 ( 
.A(n_308),
.Y(n_347)
);

NOR2xp33_ASAP7_75t_L g309 ( 
.A(n_279),
.B(n_187),
.Y(n_309)
);

NAND2xp5_ASAP7_75t_L g310 ( 
.A(n_256),
.B(n_190),
.Y(n_310)
);

NAND2xp5_ASAP7_75t_L g352 ( 
.A(n_310),
.B(n_339),
.Y(n_352)
);

INVx2_ASAP7_75t_L g311 ( 
.A(n_287),
.Y(n_311)
);

INVx1_ASAP7_75t_L g386 ( 
.A(n_311),
.Y(n_386)
);

INVx13_ASAP7_75t_L g312 ( 
.A(n_273),
.Y(n_312)
);

CKINVDCx20_ASAP7_75t_R g373 ( 
.A(n_312),
.Y(n_373)
);

CKINVDCx20_ASAP7_75t_R g313 ( 
.A(n_255),
.Y(n_313)
);

NOR2xp33_ASAP7_75t_L g366 ( 
.A(n_313),
.B(n_314),
.Y(n_366)
);

CKINVDCx20_ASAP7_75t_R g314 ( 
.A(n_266),
.Y(n_314)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_288),
.Y(n_315)
);

INVx1_ASAP7_75t_L g354 ( 
.A(n_315),
.Y(n_354)
);

NOR2xp33_ASAP7_75t_L g316 ( 
.A(n_241),
.B(n_220),
.Y(n_316)
);

NAND2xp5_ASAP7_75t_SL g365 ( 
.A(n_316),
.B(n_327),
.Y(n_365)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_288),
.Y(n_317)
);

INVx1_ASAP7_75t_L g356 ( 
.A(n_317),
.Y(n_356)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_277),
.Y(n_318)
);

INVx1_ASAP7_75t_L g357 ( 
.A(n_318),
.Y(n_357)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_242),
.Y(n_319)
);

INVx1_ASAP7_75t_L g371 ( 
.A(n_319),
.Y(n_371)
);

INVx13_ASAP7_75t_L g320 ( 
.A(n_270),
.Y(n_320)
);

CKINVDCx20_ASAP7_75t_R g383 ( 
.A(n_320),
.Y(n_383)
);

INVx3_ASAP7_75t_L g322 ( 
.A(n_257),
.Y(n_322)
);

INVx1_ASAP7_75t_L g360 ( 
.A(n_322),
.Y(n_360)
);

MAJIxp5_ASAP7_75t_L g324 ( 
.A(n_256),
.B(n_247),
.C(n_249),
.Y(n_324)
);

MAJIxp5_ASAP7_75t_L g349 ( 
.A(n_324),
.B(n_326),
.C(n_249),
.Y(n_349)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_252),
.Y(n_325)
);

INVx1_ASAP7_75t_L g372 ( 
.A(n_325),
.Y(n_372)
);

MAJIxp5_ASAP7_75t_L g326 ( 
.A(n_247),
.B(n_228),
.C(n_177),
.Y(n_326)
);

NOR2xp33_ASAP7_75t_L g327 ( 
.A(n_269),
.B(n_244),
.Y(n_327)
);

NAND2xp5_ASAP7_75t_SL g328 ( 
.A(n_275),
.B(n_253),
.Y(n_328)
);

NAND2xp5_ASAP7_75t_SL g381 ( 
.A(n_328),
.B(n_334),
.Y(n_381)
);

AND2x6_ASAP7_75t_L g329 ( 
.A(n_248),
.B(n_250),
.Y(n_329)
);

NOR2xp33_ASAP7_75t_L g374 ( 
.A(n_329),
.B(n_337),
.Y(n_374)
);

AOI22xp5_ASAP7_75t_SL g361 ( 
.A1(n_330),
.A2(n_340),
.B1(n_343),
.B2(n_246),
.Y(n_361)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_264),
.Y(n_332)
);

INVx1_ASAP7_75t_L g378 ( 
.A(n_332),
.Y(n_378)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_267),
.Y(n_333)
);

INVx1_ASAP7_75t_L g380 ( 
.A(n_333),
.Y(n_380)
);

NOR2xp33_ASAP7_75t_L g334 ( 
.A(n_260),
.B(n_234),
.Y(n_334)
);

AOI22xp5_ASAP7_75t_L g375 ( 
.A1(n_335),
.A2(n_342),
.B1(n_289),
.B2(n_257),
.Y(n_375)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_267),
.Y(n_336)
);

INVx1_ASAP7_75t_L g363 ( 
.A(n_336),
.Y(n_363)
);

INVxp67_ASAP7_75t_L g337 ( 
.A(n_243),
.Y(n_337)
);

INVx13_ASAP7_75t_L g338 ( 
.A(n_270),
.Y(n_338)
);

INVx1_ASAP7_75t_L g367 ( 
.A(n_338),
.Y(n_367)
);

NAND2xp5_ASAP7_75t_L g339 ( 
.A(n_295),
.B(n_201),
.Y(n_339)
);

CKINVDCx14_ASAP7_75t_R g340 ( 
.A(n_260),
.Y(n_340)
);

OAI22xp5_ASAP7_75t_SL g342 ( 
.A1(n_251),
.A2(n_181),
.B1(n_183),
.B2(n_211),
.Y(n_342)
);

AOI22xp33_ASAP7_75t_L g343 ( 
.A1(n_251),
.A2(n_212),
.B1(n_226),
.B2(n_196),
.Y(n_343)
);

BUFx3_ASAP7_75t_L g344 ( 
.A(n_293),
.Y(n_344)
);

INVx1_ASAP7_75t_L g376 ( 
.A(n_344),
.Y(n_376)
);

AOI21xp5_ASAP7_75t_L g346 ( 
.A1(n_330),
.A2(n_250),
.B(n_282),
.Y(n_346)
);

A2O1A1Ixp33_ASAP7_75t_SL g411 ( 
.A1(n_346),
.A2(n_307),
.B(n_329),
.C(n_321),
.Y(n_411)
);

MAJIxp5_ASAP7_75t_L g390 ( 
.A(n_349),
.B(n_355),
.C(n_359),
.Y(n_390)
);

AO21x1_ASAP7_75t_L g416 ( 
.A1(n_351),
.A2(n_370),
.B(n_331),
.Y(n_416)
);

MAJIxp5_ASAP7_75t_L g355 ( 
.A(n_324),
.B(n_265),
.C(n_294),
.Y(n_355)
);

NAND2xp5_ASAP7_75t_L g358 ( 
.A(n_296),
.B(n_314),
.Y(n_358)
);

NAND2xp5_ASAP7_75t_L g391 ( 
.A(n_358),
.B(n_361),
.Y(n_391)
);

XNOR2xp5_ASAP7_75t_L g359 ( 
.A(n_326),
.B(n_292),
.Y(n_359)
);

NAND2xp5_ASAP7_75t_L g362 ( 
.A(n_298),
.B(n_278),
.Y(n_362)
);

NAND2xp5_ASAP7_75t_L g407 ( 
.A(n_362),
.B(n_364),
.Y(n_407)
);

NAND2xp5_ASAP7_75t_L g364 ( 
.A(n_298),
.B(n_262),
.Y(n_364)
);

XNOR2xp5_ASAP7_75t_L g368 ( 
.A(n_300),
.B(n_298),
.Y(n_368)
);

MAJIxp5_ASAP7_75t_L g419 ( 
.A(n_368),
.B(n_369),
.C(n_379),
.Y(n_419)
);

XNOR2xp5_ASAP7_75t_L g369 ( 
.A(n_300),
.B(n_286),
.Y(n_369)
);

OAI21xp5_ASAP7_75t_L g370 ( 
.A1(n_330),
.A2(n_294),
.B(n_268),
.Y(n_370)
);

OAI22xp5_ASAP7_75t_L g404 ( 
.A1(n_375),
.A2(n_384),
.B1(n_318),
.B2(n_336),
.Y(n_404)
);

MAJIxp5_ASAP7_75t_L g379 ( 
.A(n_305),
.B(n_286),
.C(n_281),
.Y(n_379)
);

AOI22xp5_ASAP7_75t_L g384 ( 
.A1(n_341),
.A2(n_290),
.B1(n_281),
.B2(n_243),
.Y(n_384)
);

OAI22xp5_ASAP7_75t_SL g385 ( 
.A1(n_339),
.A2(n_290),
.B1(n_289),
.B2(n_285),
.Y(n_385)
);

AOI22xp5_ASAP7_75t_L g392 ( 
.A1(n_385),
.A2(n_335),
.B1(n_342),
.B2(n_341),
.Y(n_392)
);

INVx2_ASAP7_75t_L g387 ( 
.A(n_382),
.Y(n_387)
);

INVx1_ASAP7_75t_L g440 ( 
.A(n_387),
.Y(n_440)
);

NAND2xp5_ASAP7_75t_SL g388 ( 
.A(n_358),
.B(n_299),
.Y(n_388)
);

CKINVDCx14_ASAP7_75t_R g439 ( 
.A(n_388),
.Y(n_439)
);

INVx1_ASAP7_75t_L g389 ( 
.A(n_366),
.Y(n_389)
);

INVx1_ASAP7_75t_L g423 ( 
.A(n_389),
.Y(n_423)
);

AND2x2_ASAP7_75t_L g426 ( 
.A(n_392),
.B(n_422),
.Y(n_426)
);

AOI22xp33_ASAP7_75t_L g393 ( 
.A1(n_385),
.A2(n_321),
.B1(n_331),
.B2(n_313),
.Y(n_393)
);

INVxp67_ASAP7_75t_L g441 ( 
.A(n_393),
.Y(n_441)
);

CKINVDCx20_ASAP7_75t_R g394 ( 
.A(n_365),
.Y(n_394)
);

NAND2xp5_ASAP7_75t_SL g427 ( 
.A(n_394),
.B(n_397),
.Y(n_427)
);

INVx3_ASAP7_75t_L g395 ( 
.A(n_376),
.Y(n_395)
);

INVx1_ASAP7_75t_L g431 ( 
.A(n_395),
.Y(n_431)
);

INVx1_ASAP7_75t_L g396 ( 
.A(n_357),
.Y(n_396)
);

INVx1_ASAP7_75t_L g442 ( 
.A(n_396),
.Y(n_442)
);

NOR2xp33_ASAP7_75t_L g397 ( 
.A(n_377),
.B(n_323),
.Y(n_397)
);

CKINVDCx20_ASAP7_75t_R g398 ( 
.A(n_350),
.Y(n_398)
);

NOR2xp33_ASAP7_75t_L g453 ( 
.A(n_398),
.B(n_405),
.Y(n_453)
);

INVx1_ASAP7_75t_L g399 ( 
.A(n_371),
.Y(n_399)
);

INVx1_ASAP7_75t_L g446 ( 
.A(n_399),
.Y(n_446)
);

INVx1_ASAP7_75t_L g400 ( 
.A(n_372),
.Y(n_400)
);

INVx1_ASAP7_75t_L g450 ( 
.A(n_400),
.Y(n_450)
);

AOI22xp5_ASAP7_75t_L g401 ( 
.A1(n_379),
.A2(n_351),
.B1(n_362),
.B2(n_364),
.Y(n_401)
);

OAI22xp5_ASAP7_75t_SL g424 ( 
.A1(n_401),
.A2(n_353),
.B1(n_346),
.B2(n_361),
.Y(n_424)
);

XNOR2xp5_ASAP7_75t_L g402 ( 
.A(n_349),
.B(n_310),
.Y(n_402)
);

MAJIxp5_ASAP7_75t_L g432 ( 
.A(n_402),
.B(n_414),
.C(n_355),
.Y(n_432)
);

INVx13_ASAP7_75t_L g403 ( 
.A(n_348),
.Y(n_403)
);

INVxp67_ASAP7_75t_L g445 ( 
.A(n_403),
.Y(n_445)
);

AOI22xp5_ASAP7_75t_L g429 ( 
.A1(n_404),
.A2(n_380),
.B1(n_363),
.B2(n_352),
.Y(n_429)
);

NOR2xp33_ASAP7_75t_SL g405 ( 
.A(n_381),
.B(n_304),
.Y(n_405)
);

INVx13_ASAP7_75t_L g406 ( 
.A(n_348),
.Y(n_406)
);

INVxp67_ASAP7_75t_L g451 ( 
.A(n_406),
.Y(n_451)
);

INVx1_ASAP7_75t_L g408 ( 
.A(n_378),
.Y(n_408)
);

INVx1_ASAP7_75t_L g452 ( 
.A(n_408),
.Y(n_452)
);

HB1xp67_ASAP7_75t_L g409 ( 
.A(n_376),
.Y(n_409)
);

CKINVDCx16_ASAP7_75t_R g447 ( 
.A(n_409),
.Y(n_447)
);

NAND2xp5_ASAP7_75t_L g410 ( 
.A(n_369),
.B(n_333),
.Y(n_410)
);

NAND2xp5_ASAP7_75t_L g434 ( 
.A(n_410),
.B(n_412),
.Y(n_434)
);

NAND2x1_ASAP7_75t_L g443 ( 
.A(n_411),
.B(n_413),
.Y(n_443)
);

INVx1_ASAP7_75t_L g412 ( 
.A(n_345),
.Y(n_412)
);

AND2x2_ASAP7_75t_L g413 ( 
.A(n_370),
.B(n_311),
.Y(n_413)
);

XNOR2xp5_ASAP7_75t_L g414 ( 
.A(n_368),
.B(n_325),
.Y(n_414)
);

NOR2xp33_ASAP7_75t_L g415 ( 
.A(n_373),
.B(n_319),
.Y(n_415)
);

CKINVDCx20_ASAP7_75t_R g425 ( 
.A(n_415),
.Y(n_425)
);

AOI21xp5_ASAP7_75t_L g430 ( 
.A1(n_416),
.A2(n_374),
.B(n_352),
.Y(n_430)
);

INVx13_ASAP7_75t_L g417 ( 
.A(n_367),
.Y(n_417)
);

CKINVDCx20_ASAP7_75t_R g428 ( 
.A(n_417),
.Y(n_428)
);

OAI22xp5_ASAP7_75t_L g418 ( 
.A1(n_384),
.A2(n_322),
.B1(n_303),
.B2(n_332),
.Y(n_418)
);

NAND2xp5_ASAP7_75t_L g435 ( 
.A(n_418),
.B(n_420),
.Y(n_435)
);

INVx1_ASAP7_75t_L g420 ( 
.A(n_347),
.Y(n_420)
);

CKINVDCx20_ASAP7_75t_R g421 ( 
.A(n_383),
.Y(n_421)
);

NOR3xp33_ASAP7_75t_SL g448 ( 
.A(n_421),
.B(n_399),
.C(n_400),
.Y(n_448)
);

INVx1_ASAP7_75t_L g422 ( 
.A(n_354),
.Y(n_422)
);

AOI22xp5_ASAP7_75t_L g456 ( 
.A1(n_424),
.A2(n_413),
.B1(n_411),
.B2(n_407),
.Y(n_456)
);

OAI22xp5_ASAP7_75t_L g475 ( 
.A1(n_429),
.A2(n_444),
.B1(n_392),
.B2(n_408),
.Y(n_475)
);

CKINVDCx16_ASAP7_75t_R g477 ( 
.A(n_430),
.Y(n_477)
);

XOR2xp5_ASAP7_75t_L g466 ( 
.A(n_432),
.B(n_438),
.Y(n_466)
);

MAJIxp5_ASAP7_75t_L g433 ( 
.A(n_390),
.B(n_359),
.C(n_356),
.Y(n_433)
);

MAJIxp5_ASAP7_75t_L g459 ( 
.A(n_433),
.B(n_436),
.C(n_454),
.Y(n_459)
);

MAJIxp5_ASAP7_75t_L g436 ( 
.A(n_390),
.B(n_363),
.C(n_360),
.Y(n_436)
);

AOI21xp5_ASAP7_75t_L g437 ( 
.A1(n_391),
.A2(n_375),
.B(n_367),
.Y(n_437)
);

NOR2xp33_ASAP7_75t_L g476 ( 
.A(n_437),
.B(n_449),
.Y(n_476)
);

XOR2xp5_ASAP7_75t_L g438 ( 
.A(n_419),
.B(n_360),
.Y(n_438)
);

AOI22xp5_ASAP7_75t_SL g444 ( 
.A1(n_391),
.A2(n_386),
.B1(n_382),
.B2(n_344),
.Y(n_444)
);

CKINVDCx20_ASAP7_75t_R g455 ( 
.A(n_448),
.Y(n_455)
);

AOI21xp5_ASAP7_75t_L g449 ( 
.A1(n_416),
.A2(n_337),
.B(n_386),
.Y(n_449)
);

XNOR2xp5_ASAP7_75t_L g454 ( 
.A(n_402),
.B(n_308),
.Y(n_454)
);

INVxp67_ASAP7_75t_L g501 ( 
.A(n_456),
.Y(n_501)
);

NAND2xp5_ASAP7_75t_L g457 ( 
.A(n_434),
.B(n_410),
.Y(n_457)
);

INVx1_ASAP7_75t_L g482 ( 
.A(n_457),
.Y(n_482)
);

INVx1_ASAP7_75t_L g458 ( 
.A(n_434),
.Y(n_458)
);

INVx1_ASAP7_75t_L g483 ( 
.A(n_458),
.Y(n_483)
);

INVx1_ASAP7_75t_L g460 ( 
.A(n_435),
.Y(n_460)
);

INVx1_ASAP7_75t_L g486 ( 
.A(n_460),
.Y(n_486)
);

INVx1_ASAP7_75t_L g461 ( 
.A(n_435),
.Y(n_461)
);

INVx1_ASAP7_75t_L g491 ( 
.A(n_461),
.Y(n_491)
);

NAND2xp5_ASAP7_75t_SL g462 ( 
.A(n_425),
.B(n_419),
.Y(n_462)
);

NAND2xp5_ASAP7_75t_SL g489 ( 
.A(n_462),
.B(n_471),
.Y(n_489)
);

INVx1_ASAP7_75t_L g463 ( 
.A(n_448),
.Y(n_463)
);

INVx1_ASAP7_75t_L g497 ( 
.A(n_463),
.Y(n_497)
);

INVx1_ASAP7_75t_L g464 ( 
.A(n_446),
.Y(n_464)
);

INVx1_ASAP7_75t_L g499 ( 
.A(n_464),
.Y(n_499)
);

NAND2xp5_ASAP7_75t_L g465 ( 
.A(n_429),
.B(n_414),
.Y(n_465)
);

INVx1_ASAP7_75t_L g500 ( 
.A(n_465),
.Y(n_500)
);

AOI22xp5_ASAP7_75t_L g467 ( 
.A1(n_426),
.A2(n_413),
.B1(n_407),
.B2(n_411),
.Y(n_467)
);

HB1xp67_ASAP7_75t_L g484 ( 
.A(n_467),
.Y(n_484)
);

INVx1_ASAP7_75t_L g468 ( 
.A(n_450),
.Y(n_468)
);

NOR2xp33_ASAP7_75t_L g488 ( 
.A(n_468),
.B(n_469),
.Y(n_488)
);

INVx1_ASAP7_75t_L g469 ( 
.A(n_452),
.Y(n_469)
);

AOI22xp5_ASAP7_75t_L g470 ( 
.A1(n_426),
.A2(n_441),
.B1(n_424),
.B2(n_443),
.Y(n_470)
);

BUFx3_ASAP7_75t_L g493 ( 
.A(n_470),
.Y(n_493)
);

CKINVDCx20_ASAP7_75t_R g471 ( 
.A(n_453),
.Y(n_471)
);

HB1xp67_ASAP7_75t_L g472 ( 
.A(n_423),
.Y(n_472)
);

AOI22xp5_ASAP7_75t_L g492 ( 
.A1(n_472),
.A2(n_473),
.B1(n_475),
.B2(n_479),
.Y(n_492)
);

INVx1_ASAP7_75t_L g473 ( 
.A(n_442),
.Y(n_473)
);

NAND2xp5_ASAP7_75t_L g474 ( 
.A(n_445),
.B(n_395),
.Y(n_474)
);

XNOR2xp5_ASAP7_75t_L g496 ( 
.A(n_474),
.B(n_431),
.Y(n_496)
);

NAND2xp5_ASAP7_75t_SL g478 ( 
.A(n_427),
.B(n_401),
.Y(n_478)
);

OAI21xp5_ASAP7_75t_SL g498 ( 
.A1(n_478),
.A2(n_480),
.B(n_447),
.Y(n_498)
);

OAI22xp5_ASAP7_75t_L g479 ( 
.A1(n_439),
.A2(n_411),
.B1(n_387),
.B2(n_417),
.Y(n_479)
);

NOR2xp33_ASAP7_75t_SL g480 ( 
.A(n_436),
.B(n_312),
.Y(n_480)
);

INVx1_ASAP7_75t_L g481 ( 
.A(n_426),
.Y(n_481)
);

AOI22xp5_ASAP7_75t_L g503 ( 
.A1(n_481),
.A2(n_451),
.B1(n_445),
.B2(n_443),
.Y(n_503)
);

MAJIxp5_ASAP7_75t_L g485 ( 
.A(n_459),
.B(n_438),
.C(n_433),
.Y(n_485)
);

NAND2xp5_ASAP7_75t_L g504 ( 
.A(n_485),
.B(n_487),
.Y(n_504)
);

MAJIxp5_ASAP7_75t_L g487 ( 
.A(n_459),
.B(n_466),
.C(n_432),
.Y(n_487)
);

MAJIxp5_ASAP7_75t_L g490 ( 
.A(n_466),
.B(n_454),
.C(n_430),
.Y(n_490)
);

NAND2xp5_ASAP7_75t_SL g519 ( 
.A(n_490),
.B(n_494),
.Y(n_519)
);

MAJIxp5_ASAP7_75t_L g494 ( 
.A(n_477),
.B(n_449),
.C(n_444),
.Y(n_494)
);

XOR2xp5_ASAP7_75t_L g495 ( 
.A(n_456),
.B(n_437),
.Y(n_495)
);

XNOR2xp5_ASAP7_75t_L g513 ( 
.A(n_495),
.B(n_476),
.Y(n_513)
);

INVx1_ASAP7_75t_L g518 ( 
.A(n_496),
.Y(n_518)
);

INVxp67_ASAP7_75t_L g510 ( 
.A(n_498),
.Y(n_510)
);

MAJIxp5_ASAP7_75t_L g502 ( 
.A(n_465),
.B(n_443),
.C(n_441),
.Y(n_502)
);

MAJIxp5_ASAP7_75t_L g512 ( 
.A(n_502),
.B(n_474),
.C(n_481),
.Y(n_512)
);

INVxp67_ASAP7_75t_L g514 ( 
.A(n_503),
.Y(n_514)
);

NOR2xp33_ASAP7_75t_L g505 ( 
.A(n_489),
.B(n_455),
.Y(n_505)
);

NAND2xp5_ASAP7_75t_L g533 ( 
.A(n_505),
.B(n_516),
.Y(n_533)
);

NOR2xp33_ASAP7_75t_SL g506 ( 
.A(n_497),
.B(n_463),
.Y(n_506)
);

INVx1_ASAP7_75t_L g522 ( 
.A(n_506),
.Y(n_522)
);

XOR2xp5_ASAP7_75t_L g507 ( 
.A(n_490),
.B(n_470),
.Y(n_507)
);

XNOR2xp5_ASAP7_75t_L g523 ( 
.A(n_507),
.B(n_511),
.Y(n_523)
);

BUFx12_ASAP7_75t_L g508 ( 
.A(n_495),
.Y(n_508)
);

INVx13_ASAP7_75t_L g529 ( 
.A(n_508),
.Y(n_529)
);

AOI22xp5_ASAP7_75t_L g509 ( 
.A1(n_500),
.A2(n_461),
.B1(n_460),
.B2(n_458),
.Y(n_509)
);

OAI22xp5_ASAP7_75t_L g527 ( 
.A1(n_509),
.A2(n_520),
.B1(n_521),
.B2(n_483),
.Y(n_527)
);

XOR2xp5_ASAP7_75t_L g511 ( 
.A(n_502),
.B(n_467),
.Y(n_511)
);

NAND2xp5_ASAP7_75t_L g535 ( 
.A(n_512),
.B(n_517),
.Y(n_535)
);

XNOR2xp5_ASAP7_75t_SL g531 ( 
.A(n_513),
.B(n_515),
.Y(n_531)
);

XNOR2xp5_ASAP7_75t_SL g515 ( 
.A(n_503),
.B(n_457),
.Y(n_515)
);

MAJIxp5_ASAP7_75t_L g516 ( 
.A(n_487),
.B(n_451),
.C(n_428),
.Y(n_516)
);

CKINVDCx20_ASAP7_75t_R g517 ( 
.A(n_488),
.Y(n_517)
);

AOI22xp5_ASAP7_75t_L g520 ( 
.A1(n_501),
.A2(n_482),
.B1(n_486),
.B2(n_491),
.Y(n_520)
);

AOI22xp5_ASAP7_75t_L g521 ( 
.A1(n_501),
.A2(n_464),
.B1(n_468),
.B2(n_469),
.Y(n_521)
);

OAI21xp5_ASAP7_75t_L g524 ( 
.A1(n_514),
.A2(n_484),
.B(n_493),
.Y(n_524)
);

OAI21xp5_ASAP7_75t_L g545 ( 
.A1(n_524),
.A2(n_525),
.B(n_406),
.Y(n_545)
);

AOI21xp5_ASAP7_75t_L g525 ( 
.A1(n_514),
.A2(n_494),
.B(n_510),
.Y(n_525)
);

INVx1_ASAP7_75t_L g526 ( 
.A(n_515),
.Y(n_526)
);

NAND2xp5_ASAP7_75t_L g544 ( 
.A(n_526),
.B(n_527),
.Y(n_544)
);

XOR2xp5_ASAP7_75t_L g528 ( 
.A(n_507),
.B(n_485),
.Y(n_528)
);

XNOR2xp5_ASAP7_75t_L g536 ( 
.A(n_528),
.B(n_519),
.Y(n_536)
);

INVx1_ASAP7_75t_L g530 ( 
.A(n_518),
.Y(n_530)
);

AOI22xp5_ASAP7_75t_L g539 ( 
.A1(n_530),
.A2(n_534),
.B1(n_508),
.B2(n_440),
.Y(n_539)
);

MAJIxp5_ASAP7_75t_L g532 ( 
.A(n_504),
.B(n_512),
.C(n_511),
.Y(n_532)
);

MAJIxp5_ASAP7_75t_L g542 ( 
.A(n_532),
.B(n_508),
.C(n_317),
.Y(n_542)
);

OAI22xp5_ASAP7_75t_SL g534 ( 
.A1(n_510),
.A2(n_493),
.B1(n_492),
.B2(n_499),
.Y(n_534)
);

MAJIxp5_ASAP7_75t_L g546 ( 
.A(n_536),
.B(n_542),
.C(n_543),
.Y(n_546)
);

NOR2xp33_ASAP7_75t_SL g537 ( 
.A(n_522),
.B(n_473),
.Y(n_537)
);

INVx1_ASAP7_75t_L g548 ( 
.A(n_537),
.Y(n_548)
);

NOR2x1_ASAP7_75t_L g538 ( 
.A(n_535),
.B(n_496),
.Y(n_538)
);

OAI21x1_ASAP7_75t_L g549 ( 
.A1(n_538),
.A2(n_540),
.B(n_525),
.Y(n_549)
);

NAND2xp33_ASAP7_75t_SL g550 ( 
.A(n_539),
.B(n_541),
.Y(n_550)
);

NOR2xp33_ASAP7_75t_L g540 ( 
.A(n_532),
.B(n_440),
.Y(n_540)
);

INVxp67_ASAP7_75t_L g541 ( 
.A(n_534),
.Y(n_541)
);

MAJIxp5_ASAP7_75t_L g543 ( 
.A(n_523),
.B(n_315),
.C(n_301),
.Y(n_543)
);

OAI22xp5_ASAP7_75t_L g551 ( 
.A1(n_545),
.A2(n_524),
.B1(n_529),
.B2(n_531),
.Y(n_551)
);

MAJIxp5_ASAP7_75t_L g547 ( 
.A(n_544),
.B(n_533),
.C(n_528),
.Y(n_547)
);

NOR2xp33_ASAP7_75t_L g552 ( 
.A(n_547),
.B(n_549),
.Y(n_552)
);

NOR2xp33_ASAP7_75t_L g553 ( 
.A(n_551),
.B(n_538),
.Y(n_553)
);

INVxp67_ASAP7_75t_L g556 ( 
.A(n_553),
.Y(n_556)
);

AND2x2_ASAP7_75t_L g554 ( 
.A(n_546),
.B(n_523),
.Y(n_554)
);

OAI21xp5_ASAP7_75t_SL g555 ( 
.A1(n_554),
.A2(n_550),
.B(n_541),
.Y(n_555)
);

AOI322xp5_ASAP7_75t_L g557 ( 
.A1(n_555),
.A2(n_552),
.A3(n_529),
.B1(n_550),
.B2(n_548),
.C1(n_543),
.C2(n_531),
.Y(n_557)
);

MAJIxp5_ASAP7_75t_L g558 ( 
.A(n_557),
.B(n_556),
.C(n_403),
.Y(n_558)
);

NAND2xp5_ASAP7_75t_SL g559 ( 
.A(n_558),
.B(n_245),
.Y(n_559)
);

NOR4xp25_ASAP7_75t_L g560 ( 
.A(n_559),
.B(n_297),
.C(n_320),
.D(n_338),
.Y(n_560)
);

XOR2xp5_ASAP7_75t_L g561 ( 
.A(n_560),
.B(n_245),
.Y(n_561)
);

MAJIxp5_ASAP7_75t_L g562 ( 
.A(n_561),
.B(n_293),
.C(n_285),
.Y(n_562)
);


endmodule