module real_aes_18052_n_103 (n_17, n_28, n_76, n_56, n_34, n_98, n_90, n_82, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_83, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_91, n_100, n_43, n_96, n_54, n_35, n_42, n_99, n_15, n_9, n_23, n_72, n_95, n_44, n_102, n_7, n_4, n_80, n_6, n_12, n_68, n_79, n_69, n_46, n_59, n_25, n_73, n_77, n_81, n_48, n_37, n_97, n_70, n_50, n_89, n_26, n_86, n_93, n_13, n_24, n_2, n_55, n_62, n_84, n_67, n_92, n_33, n_88, n_14, n_11, n_85, n_16, n_94, n_39, n_5, n_45, n_60, n_38, n_87, n_0, n_78, n_101, n_63, n_1, n_53, n_36, n_103);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_98;
input n_90;
input n_82;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_83;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_91;
input n_100;
input n_43;
input n_96;
input n_54;
input n_35;
input n_42;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_95;
input n_44;
input n_102;
input n_7;
input n_4;
input n_80;
input n_6;
input n_12;
input n_68;
input n_79;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_81;
input n_48;
input n_37;
input n_97;
input n_70;
input n_50;
input n_89;
input n_26;
input n_86;
input n_93;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_84;
input n_67;
input n_92;
input n_33;
input n_88;
input n_14;
input n_11;
input n_85;
input n_16;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_87;
input n_0;
input n_78;
input n_101;
input n_63;
input n_1;
input n_53;
input n_36;
output n_103;
wire n_480;
wire n_113;
wire n_476;
wire n_758;
wire n_887;
wire n_187;
wire n_436;
wire n_599;
wire n_684;
wire n_257;
wire n_390;
wire n_821;
wire n_830;
wire n_185;
wire n_285;
wire n_624;
wire n_618;
wire n_778;
wire n_800;
wire n_522;
wire n_838;
wire n_485;
wire n_822;
wire n_846;
wire n_222;
wire n_750;
wire n_631;
wire n_357;
wire n_287;
wire n_503;
wire n_635;
wire n_386;
wire n_673;
wire n_792;
wire n_518;
wire n_254;
wire n_207;
wire n_878;
wire n_665;
wire n_667;
wire n_577;
wire n_580;
wire n_469;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_759;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_718;
wire n_318;
wire n_841;
wire n_355;
wire n_239;
wire n_669;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_761;
wire n_742;
wire n_112;
wire n_364;
wire n_319;
wire n_421;
wire n_555;
wire n_329;
wire n_852;
wire n_766;
wire n_132;
wire n_857;
wire n_131;
wire n_144;
wire n_461;
wire n_242;
wire n_169;
wire n_571;
wire n_549;
wire n_376;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_752;
wire n_448;
wire n_545;
wire n_341;
wire n_556;
wire n_593;
wire n_232;
wire n_460;
wire n_773;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_865;
wire n_537;
wire n_320;
wire n_551;
wire n_666;
wire n_884;
wire n_560;
wire n_260;
wire n_660;
wire n_814;
wire n_886;
wire n_594;
wire n_856;
wire n_186;
wire n_767;
wire n_138;
wire n_696;
wire n_889;
wire n_704;
wire n_379;
wire n_374;
wire n_453;
wire n_647;
wire n_235;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_775;
wire n_161;
wire n_763;
wire n_189;
wire n_870;
wire n_271;
wire n_489;
wire n_548;
wire n_427;
wire n_678;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_519;
wire n_564;
wire n_638;
wire n_815;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_786;
wire n_512;
wire n_395;
wire n_332;
wire n_795;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_816;
wire n_116;
wire n_625;
wire n_289;
wire n_462;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_818;
wire n_716;
wire n_213;
wire n_883;
wire n_356;
wire n_478;
wire n_584;
wire n_408;
wire n_553;
wire n_184;
wire n_578;
wire n_372;
wire n_528;
wire n_202;
wire n_495;
wire n_370;
wire n_384;
wire n_744;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_824;
wire n_875;
wire n_467;
wire n_327;
wire n_774;
wire n_813;
wire n_106;
wire n_791;
wire n_559;
wire n_466;
wire n_636;
wire n_872;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_726;
wire n_517;
wire n_683;
wire n_780;
wire n_174;
wire n_840;
wire n_570;
wire n_675;
wire n_530;
wire n_835;
wire n_104;
wire n_535;
wire n_732;
wire n_834;
wire n_882;
wire n_784;
wire n_211;
wire n_281;
wire n_496;
wire n_693;
wire n_173;
wire n_468;
wire n_234;
wire n_755;
wire n_284;
wire n_153;
wire n_532;
wire n_316;
wire n_656;
wire n_746;
wire n_178;
wire n_409;
wire n_748;
wire n_781;
wire n_860;
wire n_523;
wire n_298;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_874;
wire n_796;
wire n_297;
wire n_801;
wire n_383;
wire n_529;
wire n_119;
wire n_310;
wire n_455;
wire n_504;
wire n_725;
wire n_164;
wire n_671;
wire n_231;
wire n_547;
wire n_659;
wire n_634;
wire n_682;
wire n_454;
wire n_122;
wire n_812;
wire n_782;
wire n_443;
wire n_565;
wire n_817;
wire n_760;
wire n_608;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_885;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_819;
wire n_267;
wire n_218;
wire n_737;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_828;
wire n_808;
wire n_770;
wire n_722;
wire n_867;
wire n_745;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_879;
wire n_331;
wire n_182;
wire n_363;
wire n_417;
wire n_449;
wire n_607;
wire n_754;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_142;
wire n_561;
wire n_876;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_783;
wire n_655;
wire n_654;
wire n_505;
wire n_434;
wire n_502;
wire n_527;
wire n_769;
wire n_600;
wire n_731;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_602;
wire n_402;
wire n_552;
wire n_617;
wire n_733;
wire n_171;
wire n_676;
wire n_658;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_146;
wire n_432;
wire n_880;
wire n_807;
wire n_226;
wire n_255;
wire n_286;
wire n_416;
wire n_790;
wire n_832;
wire n_410;
wire n_120;
wire n_799;
wire n_805;
wire n_751;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_859;
wire n_695;
wire n_685;
wire n_881;
wire n_165;
wire n_361;
wire n_632;
wire n_246;
wire n_176;
wire n_768;
wire n_412;
wire n_163;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_777;
wire n_488;
wire n_501;
wire n_251;
wire n_642;
wire n_613;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_702;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_734;
wire n_110;
wire n_848;
wire n_392;
wire n_562;
wire n_150;
wire n_147;
wire n_288;
wire n_404;
wire n_598;
wire n_713;
wire n_728;
wire n_735;
wire n_756;
wire n_334;
wire n_274;
wire n_160;
wire n_569;
wire n_303;
wire n_563;
wire n_785;
wire n_188;
wire n_269;
wire n_430;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_853;
wire n_810;
wire n_843;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_193;
wire n_397;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_649;
wire n_663;
wire n_749;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_707;
wire n_622;
wire n_470;
wire n_851;
wire n_133;
wire n_494;
wire n_711;
wire n_864;
wire n_377;
wire n_273;
wire n_723;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_845;
wire n_850;
wire n_265;
wire n_354;
wire n_720;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_730;
wire n_643;
wire n_747;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_847;
wire n_779;
wire n_148;
wire n_481;
wire n_498;
wire n_691;
wire n_765;
wire n_826;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_233;
wire n_831;
wire n_487;
wire n_290;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_155;
wire n_243;
wire n_692;
wire n_544;
wire n_268;
wire n_789;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_738;
wire n_701;
wire n_309;
wire n_344;
wire n_107;
wire n_229;
wire n_827;
wire n_809;
wire n_482;
wire n_520;
wire n_633;
wire n_679;
wire n_149;
wire n_472;
wire n_866;
wire n_452;
wire n_190;
wire n_787;
wire n_262;
wire n_630;
wire n_806;
wire n_689;
wire n_820;
wire n_715;
wire n_134;
wire n_349;
wire n_336;
wire n_420;
wire n_612;
wire n_858;
wire n_873;
wire n_195;
wire n_438;
wire n_764;
wire n_794;
wire n_300;
wire n_252;
wire n_283;
wire n_314;
wire n_753;
wire n_741;
wire n_249;
wire n_623;
wire n_446;
wire n_721;
wire n_221;
wire n_681;
wire n_156;
wire n_359;
wire n_456;
wire n_717;
wire n_312;
wire n_183;
wire n_266;
wire n_712;
wire n_205;
wire n_433;
wire n_516;
wire n_177;
wire n_335;
wire n_313;
wire n_627;
wire n_739;
wire n_140;
wire n_521;
wire n_418;
wire n_422;
wire n_771;
wire n_524;
wire n_219;
wire n_861;
wire n_705;
wire n_180;
wire n_212;
wire n_210;
wire n_575;
wire n_325;
wire n_762;
wire n_338;
wire n_479;
wire n_442;
wire n_825;
wire n_740;
wire n_371;
wire n_698;
wire n_166;
wire n_541;
wire n_224;
wire n_839;
wire n_151;
wire n_546;
wire n_587;
wire n_639;
wire n_811;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_863;
wire n_724;
wire n_440;
wire n_525;
wire n_644;
wire n_674;
wire n_152;
wire n_198;
wire n_836;
wire n_888;
wire n_793;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_833;
wire n_414;
wire n_757;
wire n_123;
wire n_279;
wire n_686;
wire n_776;
wire n_803;
wire n_543;
wire n_497;
wire n_514;
wire n_507;
wire n_270;
wire n_614;
wire n_305;
wire n_586;
wire n_772;
wire n_450;
wire n_788;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_465;
wire n_473;
wire n_719;
wire n_566;
wire n_837;
wire n_871;
wire n_474;
wire n_829;
wire n_170;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_168;
wire n_175;
wire n_241;
wire n_687;
wire n_729;
wire n_844;
wire n_646;
wire n_650;
wire n_710;
wire n_105;
wire n_743;
wire n_823;
wire n_294;
wire n_393;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_307;
wire n_500;
wire n_601;
wire n_661;
wire n_463;
wire n_396;
wire n_804;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_854;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_877;
wire n_802;
wire n_868;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_842;
wire n_259;
wire n_143;
wire n_849;
wire n_192;
wire n_475;
wire n_554;
wire n_264;
wire n_855;
wire n_798;
wire n_237;
wire n_668;
wire n_797;
wire n_862;
wire n_869;
CKINVDCx5p33_ASAP7_75t_R g265 ( .A(n_0), .Y(n_265) );
AND2x4_ASAP7_75t_L g885 ( .A(n_1), .B(n_886), .Y(n_885) );
INVx1_ASAP7_75t_L g108 ( .A(n_2), .Y(n_108) );
NOR2xp33_ASAP7_75t_L g835 ( .A(n_2), .B(n_109), .Y(n_835) );
NAND2xp5_ASAP7_75t_L g838 ( .A(n_3), .B(n_839), .Y(n_838) );
INVx1_ASAP7_75t_L g861 ( .A(n_4), .Y(n_861) );
NAND2xp5_ASAP7_75t_L g873 ( .A(n_4), .B(n_874), .Y(n_873) );
BUFx3_ASAP7_75t_L g191 ( .A(n_5), .Y(n_191) );
INVx1_ASAP7_75t_L g886 ( .A(n_6), .Y(n_886) );
NAND2xp5_ASAP7_75t_L g169 ( .A(n_7), .B(n_170), .Y(n_169) );
OR2x2_ASAP7_75t_L g118 ( .A(n_8), .B(n_23), .Y(n_118) );
BUFx2_ASAP7_75t_L g881 ( .A(n_8), .Y(n_881) );
BUFx6f_ASAP7_75t_L g141 ( .A(n_9), .Y(n_141) );
NAND2xp5_ASAP7_75t_SL g208 ( .A(n_10), .B(n_148), .Y(n_208) );
NAND2xp5_ASAP7_75t_SL g563 ( .A(n_11), .B(n_148), .Y(n_563) );
NAND2xp5_ASAP7_75t_L g209 ( .A(n_12), .B(n_210), .Y(n_209) );
AOI22xp33_ASAP7_75t_L g234 ( .A1(n_13), .A2(n_83), .B1(n_143), .B2(n_148), .Y(n_234) );
OAI21x1_ASAP7_75t_L g136 ( .A1(n_14), .A2(n_37), .B(n_137), .Y(n_136) );
NAND2xp5_ASAP7_75t_L g546 ( .A(n_15), .B(n_547), .Y(n_546) );
NAND2xp5_ASAP7_75t_L g199 ( .A(n_16), .B(n_200), .Y(n_199) );
OAI22xp5_ASAP7_75t_SL g831 ( .A1(n_17), .A2(n_60), .B1(n_832), .B2(n_833), .Y(n_831) );
INVx1_ASAP7_75t_L g833 ( .A(n_17), .Y(n_833) );
CKINVDCx5p33_ASAP7_75t_R g582 ( .A(n_18), .Y(n_582) );
AO32x1_ASAP7_75t_L g231 ( .A1(n_19), .A2(n_135), .A3(n_180), .B1(n_227), .B2(n_232), .Y(n_231) );
AO32x2_ASAP7_75t_L g270 ( .A1(n_19), .A2(n_135), .A3(n_180), .B1(n_227), .B2(n_232), .Y(n_270) );
NAND2xp5_ASAP7_75t_SL g545 ( .A(n_20), .B(n_532), .Y(n_545) );
NAND2xp5_ASAP7_75t_L g555 ( .A(n_21), .B(n_180), .Y(n_555) );
CKINVDCx5p33_ASAP7_75t_R g518 ( .A(n_22), .Y(n_518) );
HB1xp67_ASAP7_75t_L g879 ( .A(n_23), .Y(n_879) );
AOI22xp33_ASAP7_75t_L g239 ( .A1(n_24), .A2(n_43), .B1(n_188), .B2(n_200), .Y(n_239) );
NAND2xp5_ASAP7_75t_L g220 ( .A(n_25), .B(n_172), .Y(n_220) );
AOI22xp5_ASAP7_75t_L g233 ( .A1(n_26), .A2(n_91), .B1(n_143), .B2(n_173), .Y(n_233) );
CKINVDCx5p33_ASAP7_75t_R g585 ( .A(n_27), .Y(n_585) );
NAND2xp5_ASAP7_75t_SL g224 ( .A(n_28), .B(n_142), .Y(n_224) );
AOI22xp33_ASAP7_75t_L g237 ( .A1(n_29), .A2(n_65), .B1(n_173), .B2(n_238), .Y(n_237) );
AOI22xp5_ASAP7_75t_L g869 ( .A1(n_30), .A2(n_57), .B1(n_870), .B2(n_871), .Y(n_869) );
INVx1_ASAP7_75t_L g870 ( .A(n_30), .Y(n_870) );
NAND2xp5_ASAP7_75t_SL g508 ( .A(n_31), .B(n_148), .Y(n_508) );
INVx2_ASAP7_75t_L g113 ( .A(n_32), .Y(n_113) );
NAND2xp5_ASAP7_75t_L g542 ( .A(n_33), .B(n_150), .Y(n_542) );
BUFx3_ASAP7_75t_L g116 ( .A(n_34), .Y(n_116) );
INVx1_ASAP7_75t_L g854 ( .A(n_34), .Y(n_854) );
NAND2xp5_ASAP7_75t_L g225 ( .A(n_35), .B(n_226), .Y(n_225) );
NAND2xp5_ASAP7_75t_L g548 ( .A(n_36), .B(n_549), .Y(n_548) );
AND2x2_ASAP7_75t_L g587 ( .A(n_38), .B(n_549), .Y(n_587) );
CKINVDCx5p33_ASAP7_75t_R g260 ( .A(n_39), .Y(n_260) );
NAND2xp5_ASAP7_75t_L g607 ( .A(n_40), .B(n_140), .Y(n_607) );
NAND2xp5_ASAP7_75t_SL g570 ( .A(n_41), .B(n_532), .Y(n_570) );
CKINVDCx5p33_ASAP7_75t_R g156 ( .A(n_42), .Y(n_156) );
NAND2xp5_ASAP7_75t_L g522 ( .A(n_44), .B(n_523), .Y(n_522) );
AOI22xp5_ASAP7_75t_L g139 ( .A1(n_45), .A2(n_78), .B1(n_140), .B2(n_142), .Y(n_139) );
NAND2xp5_ASAP7_75t_L g573 ( .A(n_46), .B(n_238), .Y(n_573) );
A2O1A1Ixp33_ASAP7_75t_L g580 ( .A1(n_47), .A2(n_201), .B(n_263), .C(n_581), .Y(n_580) );
AOI22xp33_ASAP7_75t_L g186 ( .A1(n_48), .A2(n_80), .B1(n_143), .B2(n_148), .Y(n_186) );
INVx1_ASAP7_75t_L g137 ( .A(n_49), .Y(n_137) );
AND2x4_ASAP7_75t_L g153 ( .A(n_50), .B(n_154), .Y(n_153) );
AOI22xp33_ASAP7_75t_L g534 ( .A1(n_51), .A2(n_52), .B1(n_173), .B2(n_188), .Y(n_534) );
NAND2xp5_ASAP7_75t_L g524 ( .A(n_53), .B(n_180), .Y(n_524) );
NAND2xp5_ASAP7_75t_L g609 ( .A(n_54), .B(n_549), .Y(n_609) );
CKINVDCx5p33_ASAP7_75t_R g586 ( .A(n_55), .Y(n_586) );
NAND2xp5_ASAP7_75t_SL g512 ( .A(n_56), .B(n_173), .Y(n_512) );
INVxp67_ASAP7_75t_SL g871 ( .A(n_57), .Y(n_871) );
NAND2xp5_ASAP7_75t_L g168 ( .A(n_58), .B(n_143), .Y(n_168) );
INVx1_ASAP7_75t_L g154 ( .A(n_59), .Y(n_154) );
CKINVDCx5p33_ASAP7_75t_R g832 ( .A(n_60), .Y(n_832) );
CKINVDCx5p33_ASAP7_75t_R g848 ( .A(n_61), .Y(n_848) );
NAND2xp5_ASAP7_75t_L g179 ( .A(n_62), .B(n_180), .Y(n_179) );
A2O1A1Ixp33_ASAP7_75t_L g262 ( .A1(n_63), .A2(n_222), .B(n_263), .C(n_264), .Y(n_262) );
NAND3xp33_ASAP7_75t_L g177 ( .A(n_64), .B(n_143), .C(n_175), .Y(n_177) );
CKINVDCx5p33_ASAP7_75t_R g538 ( .A(n_66), .Y(n_538) );
NAND2xp5_ASAP7_75t_L g513 ( .A(n_67), .B(n_180), .Y(n_513) );
AND2x2_ASAP7_75t_L g267 ( .A(n_68), .B(n_268), .Y(n_267) );
CKINVDCx5p33_ASAP7_75t_R g241 ( .A(n_69), .Y(n_241) );
NAND2xp5_ASAP7_75t_L g569 ( .A(n_70), .B(n_511), .Y(n_569) );
NAND3xp33_ASAP7_75t_L g543 ( .A(n_71), .B(n_150), .C(n_200), .Y(n_543) );
AOI22xp33_ASAP7_75t_L g147 ( .A1(n_72), .A2(n_95), .B1(n_140), .B2(n_148), .Y(n_147) );
INVx2_ASAP7_75t_L g146 ( .A(n_73), .Y(n_146) );
NAND2xp5_ASAP7_75t_L g203 ( .A(n_74), .B(n_204), .Y(n_203) );
NAND2xp5_ASAP7_75t_L g558 ( .A(n_75), .B(n_511), .Y(n_558) );
NAND2xp5_ASAP7_75t_SL g521 ( .A(n_76), .B(n_148), .Y(n_521) );
NAND2xp5_ASAP7_75t_SL g604 ( .A(n_77), .B(n_145), .Y(n_604) );
CKINVDCx5p33_ASAP7_75t_R g259 ( .A(n_79), .Y(n_259) );
NAND2xp5_ASAP7_75t_L g561 ( .A(n_81), .B(n_204), .Y(n_561) );
AOI22xp33_ASAP7_75t_L g530 ( .A1(n_82), .A2(n_90), .B1(n_531), .B2(n_532), .Y(n_530) );
NAND2xp5_ASAP7_75t_L g519 ( .A(n_84), .B(n_148), .Y(n_519) );
NAND2xp5_ASAP7_75t_L g174 ( .A(n_85), .B(n_175), .Y(n_174) );
NAND2xp33_ASAP7_75t_SL g608 ( .A(n_86), .B(n_170), .Y(n_608) );
NAND2xp5_ASAP7_75t_L g507 ( .A(n_87), .B(n_198), .Y(n_507) );
AOI22xp33_ASAP7_75t_L g187 ( .A1(n_88), .A2(n_102), .B1(n_173), .B2(n_188), .Y(n_187) );
NAND2xp5_ASAP7_75t_SL g219 ( .A(n_89), .B(n_142), .Y(n_219) );
INVx1_ASAP7_75t_L g124 ( .A(n_92), .Y(n_124) );
NOR2xp33_ASAP7_75t_L g852 ( .A(n_92), .B(n_853), .Y(n_852) );
AOI22xp5_ASAP7_75t_L g103 ( .A1(n_93), .A2(n_104), .B1(n_875), .B2(n_887), .Y(n_103) );
NAND2xp5_ASAP7_75t_L g228 ( .A(n_94), .B(n_210), .Y(n_228) );
NAND2xp33_ASAP7_75t_L g559 ( .A(n_96), .B(n_170), .Y(n_559) );
NAND2xp5_ASAP7_75t_L g574 ( .A(n_97), .B(n_549), .Y(n_574) );
NAND3xp33_ASAP7_75t_L g605 ( .A(n_98), .B(n_145), .C(n_170), .Y(n_605) );
NAND2xp5_ASAP7_75t_L g510 ( .A(n_99), .B(n_511), .Y(n_510) );
CKINVDCx5p33_ASAP7_75t_R g196 ( .A(n_100), .Y(n_196) );
NAND2xp5_ASAP7_75t_SL g572 ( .A(n_101), .B(n_532), .Y(n_572) );
OR2x6_ASAP7_75t_L g104 ( .A(n_105), .B(n_855), .Y(n_104) );
NAND2xp5_ASAP7_75t_L g105 ( .A(n_106), .B(n_834), .Y(n_105) );
NAND2xp5_ASAP7_75t_L g106 ( .A(n_107), .B(n_119), .Y(n_106) );
NOR2xp33_ASAP7_75t_L g107 ( .A(n_108), .B(n_109), .Y(n_107) );
BUFx4f_ASAP7_75t_L g109 ( .A(n_110), .Y(n_109) );
INVx6_ASAP7_75t_L g110 ( .A(n_111), .Y(n_110) );
AND2x6_ASAP7_75t_SL g111 ( .A(n_112), .B(n_114), .Y(n_111) );
INVx1_ASAP7_75t_L g112 ( .A(n_113), .Y(n_112) );
NOR2xp33_ASAP7_75t_L g842 ( .A(n_113), .B(n_843), .Y(n_842) );
INVx3_ASAP7_75t_L g859 ( .A(n_113), .Y(n_859) );
NAND2xp5_ASAP7_75t_L g114 ( .A(n_115), .B(n_117), .Y(n_114) );
INVx1_ASAP7_75t_L g115 ( .A(n_116), .Y(n_115) );
NOR2x1_ASAP7_75t_L g845 ( .A(n_116), .B(n_118), .Y(n_845) );
AND2x6_ASAP7_75t_SL g851 ( .A(n_117), .B(n_852), .Y(n_851) );
AND3x2_ASAP7_75t_L g865 ( .A(n_117), .B(n_866), .C(n_867), .Y(n_865) );
INVx1_ASAP7_75t_L g117 ( .A(n_118), .Y(n_117) );
INVx2_ASAP7_75t_L g836 ( .A(n_119), .Y(n_836) );
XOR2x2_ASAP7_75t_L g119 ( .A(n_120), .B(n_831), .Y(n_119) );
AOI21x1_ASAP7_75t_L g120 ( .A1(n_121), .A2(n_125), .B(n_496), .Y(n_120) );
AOI21xp5_ASAP7_75t_L g496 ( .A1(n_121), .A2(n_497), .B(n_770), .Y(n_496) );
INVx3_ASAP7_75t_L g121 ( .A(n_122), .Y(n_121) );
BUFx8_ASAP7_75t_SL g122 ( .A(n_123), .Y(n_122) );
AND2x2_ASAP7_75t_L g844 ( .A(n_123), .B(n_845), .Y(n_844) );
INVx2_ASAP7_75t_L g123 ( .A(n_124), .Y(n_123) );
BUFx2_ASAP7_75t_L g867 ( .A(n_124), .Y(n_867) );
XNOR2x1_ASAP7_75t_L g868 ( .A(n_125), .B(n_869), .Y(n_868) );
OR2x2_ASAP7_75t_L g125 ( .A(n_126), .B(n_384), .Y(n_125) );
NAND4xp25_ASAP7_75t_L g126 ( .A(n_127), .B(n_316), .C(n_343), .D(n_374), .Y(n_126) );
NOR2xp33_ASAP7_75t_L g127 ( .A(n_128), .B(n_282), .Y(n_127) );
OAI21xp33_ASAP7_75t_L g128 ( .A1(n_129), .A2(n_212), .B(n_242), .Y(n_128) );
OR2x2_ASAP7_75t_L g129 ( .A(n_130), .B(n_159), .Y(n_129) );
INVx2_ASAP7_75t_L g130 ( .A(n_131), .Y(n_130) );
OR2x2_ASAP7_75t_L g404 ( .A(n_131), .B(n_293), .Y(n_404) );
AND2x2_ASAP7_75t_L g411 ( .A(n_131), .B(n_412), .Y(n_411) );
INVx2_ASAP7_75t_SL g131 ( .A(n_132), .Y(n_131) );
OR2x2_ASAP7_75t_L g320 ( .A(n_132), .B(n_321), .Y(n_320) );
INVx2_ASAP7_75t_L g132 ( .A(n_133), .Y(n_132) );
AND2x2_ASAP7_75t_L g249 ( .A(n_133), .B(n_182), .Y(n_249) );
AND2x2_ASAP7_75t_L g277 ( .A(n_133), .B(n_278), .Y(n_277) );
INVx1_ASAP7_75t_L g286 ( .A(n_133), .Y(n_286) );
OR2x2_ASAP7_75t_L g294 ( .A(n_133), .B(n_246), .Y(n_294) );
OR2x2_ASAP7_75t_L g315 ( .A(n_133), .B(n_278), .Y(n_315) );
AND2x2_ASAP7_75t_L g324 ( .A(n_133), .B(n_192), .Y(n_324) );
INVx1_ASAP7_75t_L g397 ( .A(n_133), .Y(n_397) );
AND2x2_ASAP7_75t_L g400 ( .A(n_133), .B(n_401), .Y(n_400) );
AO31x2_ASAP7_75t_L g133 ( .A1(n_134), .A2(n_138), .A3(n_151), .B(n_155), .Y(n_133) );
AO31x2_ASAP7_75t_L g235 ( .A1(n_134), .A2(n_153), .A3(n_236), .B(n_240), .Y(n_235) );
BUFx3_ASAP7_75t_L g134 ( .A(n_135), .Y(n_134) );
INVx4_ASAP7_75t_L g180 ( .A(n_135), .Y(n_180) );
NOR2xp33_ASAP7_75t_L g189 ( .A(n_135), .B(n_190), .Y(n_189) );
INVx2_ASAP7_75t_L g193 ( .A(n_135), .Y(n_193) );
INVx2_ASAP7_75t_SL g216 ( .A(n_135), .Y(n_216) );
NOR2xp33_ASAP7_75t_L g240 ( .A(n_135), .B(n_241), .Y(n_240) );
AND2x4_ASAP7_75t_SL g564 ( .A(n_135), .B(n_178), .Y(n_564) );
INVx1_ASAP7_75t_SL g601 ( .A(n_135), .Y(n_601) );
BUFx6f_ASAP7_75t_L g135 ( .A(n_136), .Y(n_135) );
INVx2_ASAP7_75t_L g158 ( .A(n_136), .Y(n_158) );
OAI22xp5_ASAP7_75t_L g138 ( .A1(n_139), .A2(n_144), .B1(n_147), .B2(n_149), .Y(n_138) );
NOR2xp33_ASAP7_75t_L g264 ( .A(n_140), .B(n_265), .Y(n_264) );
INVx1_ASAP7_75t_L g140 ( .A(n_141), .Y(n_140) );
INVx2_ASAP7_75t_L g143 ( .A(n_141), .Y(n_143) );
BUFx6f_ASAP7_75t_L g148 ( .A(n_141), .Y(n_148) );
BUFx6f_ASAP7_75t_L g170 ( .A(n_141), .Y(n_170) );
BUFx6f_ASAP7_75t_L g173 ( .A(n_141), .Y(n_173) );
INVx1_ASAP7_75t_L g188 ( .A(n_141), .Y(n_188) );
INVx1_ASAP7_75t_L g198 ( .A(n_141), .Y(n_198) );
BUFx6f_ASAP7_75t_L g200 ( .A(n_141), .Y(n_200) );
INVx1_ASAP7_75t_L g263 ( .A(n_141), .Y(n_263) );
INVx3_ASAP7_75t_L g511 ( .A(n_141), .Y(n_511) );
INVx1_ASAP7_75t_L g533 ( .A(n_141), .Y(n_533) );
INVx2_ASAP7_75t_SL g142 ( .A(n_143), .Y(n_142) );
NOR2xp33_ASAP7_75t_L g581 ( .A(n_143), .B(n_582), .Y(n_581) );
INVx1_ASAP7_75t_SL g144 ( .A(n_145), .Y(n_144) );
INVx1_ASAP7_75t_L g261 ( .A(n_145), .Y(n_261) );
INVx1_ASAP7_75t_L g145 ( .A(n_146), .Y(n_145) );
BUFx8_ASAP7_75t_L g150 ( .A(n_146), .Y(n_150) );
INVx1_ASAP7_75t_L g176 ( .A(n_146), .Y(n_176) );
INVx2_ASAP7_75t_L g206 ( .A(n_146), .Y(n_206) );
INVx3_ASAP7_75t_L g226 ( .A(n_148), .Y(n_226) );
INVx1_ASAP7_75t_L g547 ( .A(n_148), .Y(n_547) );
OAI21xp5_ASAP7_75t_L g603 ( .A1(n_148), .A2(n_604), .B(n_605), .Y(n_603) );
OAI22xp5_ASAP7_75t_L g185 ( .A1(n_149), .A2(n_150), .B1(n_186), .B2(n_187), .Y(n_185) );
AOI21xp5_ASAP7_75t_L g223 ( .A1(n_149), .A2(n_224), .B(n_225), .Y(n_223) );
OAI22xp5_ASAP7_75t_L g236 ( .A1(n_149), .A2(n_221), .B1(n_237), .B2(n_239), .Y(n_236) );
OAI22xp5_ASAP7_75t_L g529 ( .A1(n_149), .A2(n_530), .B1(n_534), .B2(n_535), .Y(n_529) );
INVx6_ASAP7_75t_L g149 ( .A(n_150), .Y(n_149) );
AOI21xp5_ASAP7_75t_L g167 ( .A1(n_150), .A2(n_168), .B(n_169), .Y(n_167) );
OAI22xp5_ASAP7_75t_L g232 ( .A1(n_150), .A2(n_201), .B1(n_233), .B2(n_234), .Y(n_232) );
AOI21xp5_ASAP7_75t_L g509 ( .A1(n_150), .A2(n_510), .B(n_512), .Y(n_509) );
O2A1O1Ixp5_ASAP7_75t_L g517 ( .A1(n_150), .A2(n_197), .B(n_518), .C(n_519), .Y(n_517) );
INVx2_ASAP7_75t_SL g151 ( .A(n_152), .Y(n_151) );
INVx2_ASAP7_75t_SL g227 ( .A(n_152), .Y(n_227) );
INVx1_ASAP7_75t_L g152 ( .A(n_153), .Y(n_152) );
BUFx10_ASAP7_75t_L g178 ( .A(n_153), .Y(n_178) );
INVx1_ASAP7_75t_L g266 ( .A(n_153), .Y(n_266) );
BUFx10_ASAP7_75t_L g536 ( .A(n_153), .Y(n_536) );
NOR2xp33_ASAP7_75t_L g155 ( .A(n_156), .B(n_157), .Y(n_155) );
INVx2_ASAP7_75t_L g268 ( .A(n_157), .Y(n_268) );
NOR2xp33_ASAP7_75t_L g537 ( .A(n_157), .B(n_538), .Y(n_537) );
INVx2_ASAP7_75t_L g157 ( .A(n_158), .Y(n_157) );
INVx2_ASAP7_75t_L g165 ( .A(n_158), .Y(n_165) );
INVx2_ASAP7_75t_L g211 ( .A(n_158), .Y(n_211) );
NAND2xp5_ASAP7_75t_L g159 ( .A(n_160), .B(n_181), .Y(n_159) );
INVx2_ASAP7_75t_L g313 ( .A(n_160), .Y(n_313) );
INVx2_ASAP7_75t_L g160 ( .A(n_161), .Y(n_160) );
INVx1_ASAP7_75t_L g421 ( .A(n_161), .Y(n_421) );
INVx1_ASAP7_75t_L g161 ( .A(n_162), .Y(n_161) );
INVx1_ASAP7_75t_L g366 ( .A(n_162), .Y(n_366) );
INVx2_ASAP7_75t_L g162 ( .A(n_163), .Y(n_162) );
OR2x2_ASAP7_75t_L g293 ( .A(n_163), .B(n_279), .Y(n_293) );
OAI21x1_ASAP7_75t_L g163 ( .A1(n_164), .A2(n_166), .B(n_179), .Y(n_163) );
OAI21xp5_ASAP7_75t_L g247 ( .A1(n_164), .A2(n_166), .B(n_179), .Y(n_247) );
OAI21x1_ASAP7_75t_L g515 ( .A1(n_164), .A2(n_516), .B(n_524), .Y(n_515) );
OAI21xp33_ASAP7_75t_SL g566 ( .A1(n_164), .A2(n_567), .B(n_574), .Y(n_566) );
OAI21x1_ASAP7_75t_L g616 ( .A1(n_164), .A2(n_567), .B(n_574), .Y(n_616) );
OAI21xp5_ASAP7_75t_L g670 ( .A1(n_164), .A2(n_516), .B(n_524), .Y(n_670) );
INVx2_ASAP7_75t_L g164 ( .A(n_165), .Y(n_164) );
INVx2_ASAP7_75t_L g549 ( .A(n_165), .Y(n_549) );
OAI21x1_ASAP7_75t_L g166 ( .A1(n_167), .A2(n_171), .B(n_178), .Y(n_166) );
INVx2_ASAP7_75t_L g523 ( .A(n_170), .Y(n_523) );
OAI21xp5_ASAP7_75t_L g171 ( .A1(n_172), .A2(n_174), .B(n_177), .Y(n_171) );
INVx2_ASAP7_75t_L g172 ( .A(n_173), .Y(n_172) );
INVx2_ASAP7_75t_L g531 ( .A(n_173), .Y(n_531) );
OAI21xp5_ASAP7_75t_L g541 ( .A1(n_173), .A2(n_542), .B(n_543), .Y(n_541) );
OAI22xp33_ASAP7_75t_L g584 ( .A1(n_173), .A2(n_511), .B1(n_585), .B2(n_586), .Y(n_584) );
INVx1_ASAP7_75t_L g175 ( .A(n_176), .Y(n_175) );
BUFx4f_ASAP7_75t_L g201 ( .A(n_176), .Y(n_201) );
AOI31xp67_ASAP7_75t_L g183 ( .A1(n_178), .A2(n_184), .A3(n_185), .B(n_189), .Y(n_183) );
OAI21x1_ASAP7_75t_L g194 ( .A1(n_178), .A2(n_195), .B(n_202), .Y(n_194) );
OAI21x1_ASAP7_75t_L g505 ( .A1(n_178), .A2(n_506), .B(n_509), .Y(n_505) );
OAI21x1_ASAP7_75t_L g516 ( .A1(n_178), .A2(n_517), .B(n_520), .Y(n_516) );
OAI21x1_ASAP7_75t_L g540 ( .A1(n_178), .A2(n_541), .B(n_544), .Y(n_540) );
OAI21x1_ASAP7_75t_L g567 ( .A1(n_178), .A2(n_568), .B(n_571), .Y(n_567) );
OAI21x1_ASAP7_75t_L g602 ( .A1(n_178), .A2(n_603), .B(n_606), .Y(n_602) );
INVx2_ASAP7_75t_L g184 ( .A(n_180), .Y(n_184) );
HB1xp67_ASAP7_75t_L g475 ( .A(n_181), .Y(n_475) );
AND2x2_ASAP7_75t_L g181 ( .A(n_182), .B(n_192), .Y(n_181) );
INVx2_ASAP7_75t_L g287 ( .A(n_182), .Y(n_287) );
AND2x2_ASAP7_75t_L g325 ( .A(n_182), .B(n_247), .Y(n_325) );
INVx2_ASAP7_75t_L g182 ( .A(n_183), .Y(n_182) );
INVx1_ASAP7_75t_L g279 ( .A(n_183), .Y(n_279) );
INVx1_ASAP7_75t_L g207 ( .A(n_188), .Y(n_207) );
OAI22xp5_ASAP7_75t_L g258 ( .A1(n_188), .A2(n_200), .B1(n_259), .B2(n_260), .Y(n_258) );
CKINVDCx5p33_ASAP7_75t_R g190 ( .A(n_191), .Y(n_190) );
AND2x2_ASAP7_75t_L g281 ( .A(n_192), .B(n_247), .Y(n_281) );
INVx1_ASAP7_75t_L g367 ( .A(n_192), .Y(n_367) );
OA21x2_ASAP7_75t_L g192 ( .A1(n_193), .A2(n_194), .B(n_209), .Y(n_192) );
OA21x2_ASAP7_75t_L g246 ( .A1(n_193), .A2(n_194), .B(n_209), .Y(n_246) );
OAI21x1_ASAP7_75t_L g504 ( .A1(n_193), .A2(n_505), .B(n_513), .Y(n_504) );
OA21x2_ASAP7_75t_L g539 ( .A1(n_193), .A2(n_540), .B(n_548), .Y(n_539) );
OAI21x1_ASAP7_75t_L g629 ( .A1(n_193), .A2(n_505), .B(n_513), .Y(n_629) );
OAI21x1_ASAP7_75t_L g667 ( .A1(n_193), .A2(n_540), .B(n_548), .Y(n_667) );
O2A1O1Ixp5_ASAP7_75t_L g195 ( .A1(n_196), .A2(n_197), .B(n_199), .C(n_201), .Y(n_195) );
INVx2_ASAP7_75t_L g197 ( .A(n_198), .Y(n_197) );
INVx2_ASAP7_75t_L g238 ( .A(n_200), .Y(n_238) );
AOI21xp5_ASAP7_75t_L g506 ( .A1(n_201), .A2(n_507), .B(n_508), .Y(n_506) );
AOI21xp5_ASAP7_75t_L g557 ( .A1(n_201), .A2(n_558), .B(n_559), .Y(n_557) );
AOI21xp5_ASAP7_75t_L g568 ( .A1(n_201), .A2(n_569), .B(n_570), .Y(n_568) );
AOI21xp5_ASAP7_75t_L g606 ( .A1(n_201), .A2(n_607), .B(n_608), .Y(n_606) );
OAI22xp5_ASAP7_75t_L g202 ( .A1(n_203), .A2(n_205), .B1(n_207), .B2(n_208), .Y(n_202) );
AOI21xp5_ASAP7_75t_L g520 ( .A1(n_204), .A2(n_521), .B(n_522), .Y(n_520) );
INVx2_ASAP7_75t_SL g204 ( .A(n_205), .Y(n_204) );
OAI22xp5_ASAP7_75t_L g560 ( .A1(n_205), .A2(n_561), .B1(n_562), .B2(n_563), .Y(n_560) );
INVx2_ASAP7_75t_L g205 ( .A(n_206), .Y(n_205) );
BUFx3_ASAP7_75t_L g222 ( .A(n_206), .Y(n_222) );
INVx2_ASAP7_75t_L g255 ( .A(n_210), .Y(n_255) );
NOR2xp67_ASAP7_75t_SL g577 ( .A(n_210), .B(n_578), .Y(n_577) );
INVx2_ASAP7_75t_L g210 ( .A(n_211), .Y(n_210) );
AO31x2_ASAP7_75t_L g528 ( .A1(n_211), .A2(n_529), .A3(n_536), .B(n_537), .Y(n_528) );
O2A1O1Ixp33_ASAP7_75t_SL g425 ( .A1(n_212), .A2(n_426), .B(n_427), .C(n_429), .Y(n_425) );
OR2x2_ASAP7_75t_L g212 ( .A(n_213), .B(n_229), .Y(n_212) );
OR2x2_ASAP7_75t_L g373 ( .A(n_213), .B(n_357), .Y(n_373) );
INVxp67_ASAP7_75t_SL g435 ( .A(n_213), .Y(n_435) );
INVx2_ASAP7_75t_L g213 ( .A(n_214), .Y(n_213) );
AND2x2_ASAP7_75t_L g269 ( .A(n_214), .B(n_270), .Y(n_269) );
OR2x2_ASAP7_75t_L g301 ( .A(n_214), .B(n_273), .Y(n_301) );
INVx3_ASAP7_75t_L g303 ( .A(n_214), .Y(n_303) );
INVxp67_ASAP7_75t_L g311 ( .A(n_214), .Y(n_311) );
INVx1_ASAP7_75t_L g321 ( .A(n_214), .Y(n_321) );
BUFx2_ASAP7_75t_L g347 ( .A(n_214), .Y(n_347) );
OR2x2_ASAP7_75t_L g370 ( .A(n_214), .B(n_371), .Y(n_370) );
AND2x2_ASAP7_75t_L g409 ( .A(n_214), .B(n_371), .Y(n_409) );
NAND2xp5_ASAP7_75t_L g457 ( .A(n_214), .B(n_235), .Y(n_457) );
INVx1_ASAP7_75t_L g483 ( .A(n_214), .Y(n_483) );
BUFx6f_ASAP7_75t_L g214 ( .A(n_215), .Y(n_214) );
OAI21x1_ASAP7_75t_L g215 ( .A1(n_216), .A2(n_217), .B(n_228), .Y(n_215) );
OAI21x1_ASAP7_75t_L g217 ( .A1(n_218), .A2(n_223), .B(n_227), .Y(n_217) );
AOI21x1_ASAP7_75t_L g218 ( .A1(n_219), .A2(n_220), .B(n_221), .Y(n_218) );
AOI21xp5_ASAP7_75t_L g571 ( .A1(n_221), .A2(n_572), .B(n_573), .Y(n_571) );
INVx2_ASAP7_75t_L g221 ( .A(n_222), .Y(n_221) );
INVx2_ASAP7_75t_L g535 ( .A(n_222), .Y(n_535) );
NOR2xp33_ASAP7_75t_L g462 ( .A(n_229), .B(n_301), .Y(n_462) );
INVx2_ASAP7_75t_SL g229 ( .A(n_230), .Y(n_229) );
AND2x2_ASAP7_75t_L g302 ( .A(n_230), .B(n_303), .Y(n_302) );
AND2x2_ASAP7_75t_L g388 ( .A(n_230), .B(n_335), .Y(n_388) );
AND2x2_ASAP7_75t_L g405 ( .A(n_230), .B(n_334), .Y(n_405) );
AND2x2_ASAP7_75t_L g230 ( .A(n_231), .B(n_235), .Y(n_230) );
OR2x2_ASAP7_75t_L g357 ( .A(n_231), .B(n_235), .Y(n_357) );
INVx1_ASAP7_75t_L g424 ( .A(n_231), .Y(n_424) );
INVx1_ASAP7_75t_L g437 ( .A(n_231), .Y(n_437) );
INVx3_ASAP7_75t_L g272 ( .A(n_235), .Y(n_272) );
AND2x2_ASAP7_75t_L g327 ( .A(n_235), .B(n_253), .Y(n_327) );
AND2x2_ASAP7_75t_L g348 ( .A(n_235), .B(n_349), .Y(n_348) );
AOI22xp5_ASAP7_75t_L g242 ( .A1(n_243), .A2(n_250), .B1(n_271), .B2(n_274), .Y(n_242) );
AOI22xp5_ASAP7_75t_L g484 ( .A1(n_243), .A2(n_382), .B1(n_485), .B2(n_487), .Y(n_484) );
INVx3_ASAP7_75t_L g243 ( .A(n_244), .Y(n_243) );
OR2x2_ASAP7_75t_L g244 ( .A(n_245), .B(n_248), .Y(n_244) );
OR2x2_ASAP7_75t_L g396 ( .A(n_245), .B(n_397), .Y(n_396) );
INVx1_ASAP7_75t_L g430 ( .A(n_245), .Y(n_430) );
OR2x2_ASAP7_75t_L g245 ( .A(n_246), .B(n_247), .Y(n_245) );
BUFx2_ASAP7_75t_L g306 ( .A(n_246), .Y(n_306) );
INVx2_ASAP7_75t_SL g330 ( .A(n_246), .Y(n_330) );
AND2x2_ASAP7_75t_L g350 ( .A(n_246), .B(n_286), .Y(n_350) );
INVx1_ASAP7_75t_L g401 ( .A(n_246), .Y(n_401) );
INVx1_ASAP7_75t_L g390 ( .A(n_248), .Y(n_390) );
INVx2_ASAP7_75t_L g248 ( .A(n_249), .Y(n_248) );
AND2x4_ASAP7_75t_L g382 ( .A(n_249), .B(n_364), .Y(n_382) );
AO22x1_ASAP7_75t_L g470 ( .A1(n_250), .A2(n_323), .B1(n_471), .B2(n_472), .Y(n_470) );
AND2x2_ASAP7_75t_L g250 ( .A(n_251), .B(n_269), .Y(n_250) );
INVx1_ASAP7_75t_L g251 ( .A(n_252), .Y(n_251) );
HB1xp67_ASAP7_75t_L g252 ( .A(n_253), .Y(n_252) );
INVx1_ASAP7_75t_L g289 ( .A(n_253), .Y(n_289) );
INVx1_ASAP7_75t_L g298 ( .A(n_253), .Y(n_298) );
INVx1_ASAP7_75t_L g349 ( .A(n_253), .Y(n_349) );
INVx2_ASAP7_75t_L g253 ( .A(n_254), .Y(n_253) );
INVx1_ASAP7_75t_L g273 ( .A(n_254), .Y(n_273) );
AOI21x1_ASAP7_75t_L g254 ( .A1(n_255), .A2(n_256), .B(n_267), .Y(n_254) );
AOI21xp5_ASAP7_75t_L g256 ( .A1(n_257), .A2(n_262), .B(n_266), .Y(n_256) );
NAND2xp5_ASAP7_75t_SL g257 ( .A(n_258), .B(n_261), .Y(n_257) );
AOI21x1_ASAP7_75t_L g544 ( .A1(n_261), .A2(n_545), .B(n_546), .Y(n_544) );
INVx1_ASAP7_75t_L g562 ( .A(n_263), .Y(n_562) );
AND2x2_ASAP7_75t_L g469 ( .A(n_269), .B(n_379), .Y(n_469) );
AND2x4_ASAP7_75t_L g336 ( .A(n_270), .B(n_272), .Y(n_336) );
INVx1_ASAP7_75t_L g371 ( .A(n_270), .Y(n_371) );
INVx1_ASAP7_75t_L g445 ( .A(n_270), .Y(n_445) );
NAND2xp5_ASAP7_75t_L g310 ( .A(n_271), .B(n_311), .Y(n_310) );
NAND2xp5_ASAP7_75t_L g488 ( .A(n_271), .B(n_489), .Y(n_488) );
AND2x2_ASAP7_75t_L g271 ( .A(n_272), .B(n_273), .Y(n_271) );
AND2x4_ASAP7_75t_L g297 ( .A(n_272), .B(n_298), .Y(n_297) );
INVx1_ASAP7_75t_L g416 ( .A(n_272), .Y(n_416) );
INVx1_ASAP7_75t_L g335 ( .A(n_273), .Y(n_335) );
INVx1_ASAP7_75t_L g355 ( .A(n_273), .Y(n_355) );
OR2x2_ASAP7_75t_L g436 ( .A(n_273), .B(n_437), .Y(n_436) );
INVx2_ASAP7_75t_L g274 ( .A(n_275), .Y(n_274) );
OR2x2_ASAP7_75t_L g275 ( .A(n_276), .B(n_280), .Y(n_275) );
INVx1_ASAP7_75t_L g276 ( .A(n_277), .Y(n_276) );
AND2x2_ASAP7_75t_L g463 ( .A(n_277), .B(n_306), .Y(n_463) );
AND2x2_ASAP7_75t_L g471 ( .A(n_277), .B(n_313), .Y(n_471) );
INVx1_ASAP7_75t_L g278 ( .A(n_279), .Y(n_278) );
OR2x2_ASAP7_75t_L g413 ( .A(n_280), .B(n_363), .Y(n_413) );
INVx1_ASAP7_75t_L g280 ( .A(n_281), .Y(n_280) );
AND2x2_ASAP7_75t_L g284 ( .A(n_281), .B(n_285), .Y(n_284) );
INVx1_ASAP7_75t_SL g391 ( .A(n_281), .Y(n_391) );
OAI211xp5_ASAP7_75t_L g282 ( .A1(n_283), .A2(n_288), .B(n_290), .C(n_308), .Y(n_282) );
OAI322xp33_ASAP7_75t_L g328 ( .A1(n_283), .A2(n_320), .A3(n_329), .B1(n_332), .B2(n_337), .C1(n_340), .C2(n_342), .Y(n_328) );
INVx2_ASAP7_75t_L g283 ( .A(n_284), .Y(n_283) );
AND2x2_ASAP7_75t_L g338 ( .A(n_285), .B(n_339), .Y(n_338) );
INVx2_ASAP7_75t_L g394 ( .A(n_285), .Y(n_394) );
AND2x2_ASAP7_75t_L g285 ( .A(n_286), .B(n_287), .Y(n_285) );
INVx1_ASAP7_75t_L g363 ( .A(n_287), .Y(n_363) );
AND2x2_ASAP7_75t_L g402 ( .A(n_287), .B(n_366), .Y(n_402) );
INVx1_ASAP7_75t_L g495 ( .A(n_287), .Y(n_495) );
INVx1_ASAP7_75t_L g473 ( .A(n_288), .Y(n_473) );
OAI211xp5_ASAP7_75t_L g493 ( .A1(n_288), .A2(n_372), .B(n_415), .C(n_494), .Y(n_493) );
INVx1_ASAP7_75t_L g288 ( .A(n_289), .Y(n_288) );
AOI22xp5_ASAP7_75t_L g290 ( .A1(n_291), .A2(n_295), .B1(n_302), .B2(n_304), .Y(n_290) );
OAI21xp5_ASAP7_75t_L g368 ( .A1(n_291), .A2(n_369), .B(n_372), .Y(n_368) );
INVx1_ASAP7_75t_L g291 ( .A(n_292), .Y(n_291) );
OR2x2_ASAP7_75t_L g292 ( .A(n_293), .B(n_294), .Y(n_292) );
INVx2_ASAP7_75t_L g307 ( .A(n_293), .Y(n_307) );
INVx1_ASAP7_75t_L g331 ( .A(n_293), .Y(n_331) );
INVx1_ASAP7_75t_L g412 ( .A(n_293), .Y(n_412) );
INVx1_ASAP7_75t_L g441 ( .A(n_294), .Y(n_441) );
NAND2xp5_ASAP7_75t_L g295 ( .A(n_296), .B(n_299), .Y(n_295) );
HB1xp67_ASAP7_75t_L g492 ( .A(n_296), .Y(n_492) );
INVx2_ASAP7_75t_L g296 ( .A(n_297), .Y(n_296) );
NAND2x1p5_ASAP7_75t_L g428 ( .A(n_297), .B(n_409), .Y(n_428) );
INVx1_ASAP7_75t_L g379 ( .A(n_298), .Y(n_379) );
INVx1_ASAP7_75t_L g299 ( .A(n_300), .Y(n_299) );
NAND2x1_ASAP7_75t_SL g340 ( .A(n_300), .B(n_341), .Y(n_340) );
INVx3_ASAP7_75t_L g300 ( .A(n_301), .Y(n_300) );
NOR2xp33_ASAP7_75t_L g360 ( .A(n_301), .B(n_336), .Y(n_360) );
AND2x2_ASAP7_75t_L g423 ( .A(n_303), .B(n_424), .Y(n_423) );
AND2x2_ASAP7_75t_L g304 ( .A(n_305), .B(n_307), .Y(n_304) );
INVx1_ASAP7_75t_L g305 ( .A(n_306), .Y(n_305) );
AND2x2_ASAP7_75t_L g322 ( .A(n_306), .B(n_307), .Y(n_322) );
NAND2xp5_ASAP7_75t_L g308 ( .A(n_309), .B(n_312), .Y(n_308) );
INVx1_ASAP7_75t_L g309 ( .A(n_310), .Y(n_309) );
AND2x2_ASAP7_75t_L g476 ( .A(n_311), .B(n_333), .Y(n_476) );
INVx1_ASAP7_75t_L g489 ( .A(n_311), .Y(n_489) );
AND2x2_ASAP7_75t_L g312 ( .A(n_313), .B(n_314), .Y(n_312) );
INVx1_ASAP7_75t_L g393 ( .A(n_313), .Y(n_393) );
NAND2xp5_ASAP7_75t_L g383 ( .A(n_314), .B(n_339), .Y(n_383) );
INVx1_ASAP7_75t_L g426 ( .A(n_314), .Y(n_426) );
INVx1_ASAP7_75t_L g314 ( .A(n_315), .Y(n_314) );
INVx1_ASAP7_75t_L g353 ( .A(n_315), .Y(n_353) );
OR2x2_ASAP7_75t_L g482 ( .A(n_315), .B(n_483), .Y(n_482) );
O2A1O1Ixp5_ASAP7_75t_L g316 ( .A1(n_317), .A2(n_323), .B(n_326), .C(n_328), .Y(n_316) );
INVxp67_ASAP7_75t_SL g317 ( .A(n_318), .Y(n_317) );
NAND2xp5_ASAP7_75t_SL g318 ( .A(n_319), .B(n_322), .Y(n_318) );
INVx1_ASAP7_75t_L g319 ( .A(n_320), .Y(n_319) );
AND2x2_ASAP7_75t_L g415 ( .A(n_321), .B(n_416), .Y(n_415) );
INVx2_ASAP7_75t_L g460 ( .A(n_322), .Y(n_460) );
INVx2_ASAP7_75t_L g453 ( .A(n_323), .Y(n_453) );
AND2x2_ASAP7_75t_L g323 ( .A(n_324), .B(n_325), .Y(n_323) );
AOI21xp5_ASAP7_75t_L g374 ( .A1(n_324), .A2(n_375), .B(n_380), .Y(n_374) );
AND2x2_ASAP7_75t_L g440 ( .A(n_325), .B(n_441), .Y(n_440) );
BUFx2_ASAP7_75t_L g326 ( .A(n_327), .Y(n_326) );
AND2x2_ASAP7_75t_L g408 ( .A(n_327), .B(n_409), .Y(n_408) );
AND2x4_ASAP7_75t_L g422 ( .A(n_327), .B(n_423), .Y(n_422) );
NAND2xp5_ASAP7_75t_L g449 ( .A(n_327), .B(n_450), .Y(n_449) );
NAND2xp5_ASAP7_75t_L g329 ( .A(n_330), .B(n_331), .Y(n_329) );
INVx2_ASAP7_75t_L g339 ( .A(n_330), .Y(n_339) );
NAND2xp5_ASAP7_75t_L g352 ( .A(n_330), .B(n_353), .Y(n_352) );
HB1xp67_ASAP7_75t_L g478 ( .A(n_330), .Y(n_478) );
AOI21xp33_ASAP7_75t_L g380 ( .A1(n_332), .A2(n_381), .B(n_383), .Y(n_380) );
INVx2_ASAP7_75t_L g332 ( .A(n_333), .Y(n_332) );
AND2x2_ASAP7_75t_L g333 ( .A(n_334), .B(n_336), .Y(n_333) );
INVx1_ASAP7_75t_L g334 ( .A(n_335), .Y(n_334) );
INVx3_ASAP7_75t_L g342 ( .A(n_336), .Y(n_342) );
AND2x4_ASAP7_75t_L g467 ( .A(n_336), .B(n_355), .Y(n_467) );
INVx2_ASAP7_75t_SL g337 ( .A(n_338), .Y(n_337) );
INVx2_ASAP7_75t_L g341 ( .A(n_342), .Y(n_341) );
AOI221xp5_ASAP7_75t_L g343 ( .A1(n_344), .A2(n_350), .B1(n_351), .B2(n_354), .C(n_358), .Y(n_343) );
INVx1_ASAP7_75t_L g344 ( .A(n_345), .Y(n_344) );
HB1xp67_ASAP7_75t_L g345 ( .A(n_346), .Y(n_345) );
INVx1_ASAP7_75t_L g464 ( .A(n_346), .Y(n_464) );
NAND2xp5_ASAP7_75t_L g346 ( .A(n_347), .B(n_348), .Y(n_346) );
BUFx2_ASAP7_75t_L g377 ( .A(n_347), .Y(n_377) );
INVx1_ASAP7_75t_L g351 ( .A(n_352), .Y(n_351) );
AND2x2_ASAP7_75t_L g354 ( .A(n_355), .B(n_356), .Y(n_354) );
OR2x2_ASAP7_75t_L g486 ( .A(n_355), .B(n_370), .Y(n_486) );
AND2x4_ASAP7_75t_L g378 ( .A(n_356), .B(n_379), .Y(n_378) );
INVx2_ASAP7_75t_L g356 ( .A(n_357), .Y(n_356) );
OAI21xp5_ASAP7_75t_SL g358 ( .A1(n_359), .A2(n_361), .B(n_368), .Y(n_358) );
INVxp67_ASAP7_75t_L g359 ( .A(n_360), .Y(n_359) );
INVx1_ASAP7_75t_L g361 ( .A(n_362), .Y(n_361) );
AND2x2_ASAP7_75t_L g362 ( .A(n_363), .B(n_364), .Y(n_362) );
AND2x2_ASAP7_75t_L g447 ( .A(n_364), .B(n_397), .Y(n_447) );
INVx2_ASAP7_75t_L g364 ( .A(n_365), .Y(n_364) );
NAND2x1p5_ASAP7_75t_L g365 ( .A(n_366), .B(n_367), .Y(n_365) );
INVx2_ASAP7_75t_L g369 ( .A(n_370), .Y(n_369) );
INVx2_ASAP7_75t_L g372 ( .A(n_373), .Y(n_372) );
INVx1_ASAP7_75t_L g375 ( .A(n_376), .Y(n_375) );
NAND2xp5_ASAP7_75t_L g376 ( .A(n_377), .B(n_378), .Y(n_376) );
INVx1_ASAP7_75t_L g459 ( .A(n_378), .Y(n_459) );
INVx1_ASAP7_75t_L g381 ( .A(n_382), .Y(n_381) );
NAND2xp5_ASAP7_75t_L g468 ( .A(n_382), .B(n_469), .Y(n_468) );
NAND3xp33_ASAP7_75t_SL g384 ( .A(n_385), .B(n_431), .C(n_474), .Y(n_384) );
NOR3xp33_ASAP7_75t_L g385 ( .A(n_386), .B(n_406), .C(n_425), .Y(n_385) );
OAI21xp5_ASAP7_75t_SL g386 ( .A1(n_387), .A2(n_389), .B(n_398), .Y(n_386) );
INVx2_ASAP7_75t_L g387 ( .A(n_388), .Y(n_387) );
AOI211x1_ASAP7_75t_SL g389 ( .A1(n_390), .A2(n_391), .B(n_392), .C(n_395), .Y(n_389) );
OAI322xp33_ASAP7_75t_L g432 ( .A1(n_390), .A2(n_433), .A3(n_438), .B1(n_439), .B2(n_442), .C1(n_446), .C2(n_448), .Y(n_432) );
NOR2xp67_ASAP7_75t_L g392 ( .A(n_393), .B(n_394), .Y(n_392) );
O2A1O1Ixp5_ASAP7_75t_SL g490 ( .A1(n_393), .A2(n_491), .B(n_492), .C(n_493), .Y(n_490) );
INVx3_ASAP7_75t_L g395 ( .A(n_396), .Y(n_395) );
NAND2xp5_ASAP7_75t_L g420 ( .A(n_397), .B(n_421), .Y(n_420) );
OAI21xp5_ASAP7_75t_L g398 ( .A1(n_399), .A2(n_403), .B(n_405), .Y(n_398) );
AOI22xp5_ASAP7_75t_L g461 ( .A1(n_399), .A2(n_462), .B1(n_463), .B2(n_464), .Y(n_461) );
AND2x4_ASAP7_75t_L g399 ( .A(n_400), .B(n_402), .Y(n_399) );
INVx1_ASAP7_75t_L g403 ( .A(n_404), .Y(n_403) );
OAI221xp5_ASAP7_75t_L g406 ( .A1(n_407), .A2(n_410), .B1(n_413), .B2(n_414), .C(n_417), .Y(n_406) );
INVx1_ASAP7_75t_L g407 ( .A(n_408), .Y(n_407) );
INVx1_ASAP7_75t_L g410 ( .A(n_411), .Y(n_410) );
INVx1_ASAP7_75t_L g414 ( .A(n_415), .Y(n_414) );
NAND2xp5_ASAP7_75t_L g417 ( .A(n_418), .B(n_422), .Y(n_417) );
INVx1_ASAP7_75t_L g418 ( .A(n_419), .Y(n_418) );
HB1xp67_ASAP7_75t_L g419 ( .A(n_420), .Y(n_419) );
INVx2_ASAP7_75t_L g451 ( .A(n_424), .Y(n_451) );
INVx1_ASAP7_75t_L g458 ( .A(n_424), .Y(n_458) );
HB1xp67_ASAP7_75t_L g427 ( .A(n_428), .Y(n_427) );
INVx1_ASAP7_75t_L g429 ( .A(n_430), .Y(n_429) );
INVx1_ASAP7_75t_L g438 ( .A(n_430), .Y(n_438) );
NOR4xp25_ASAP7_75t_L g431 ( .A(n_432), .B(n_452), .C(n_465), .D(n_470), .Y(n_431) );
INVx1_ASAP7_75t_L g433 ( .A(n_434), .Y(n_433) );
NOR2x1p5_ASAP7_75t_L g434 ( .A(n_435), .B(n_436), .Y(n_434) );
INVx2_ASAP7_75t_L g439 ( .A(n_440), .Y(n_439) );
INVx1_ASAP7_75t_L g442 ( .A(n_443), .Y(n_442) );
INVx2_ASAP7_75t_L g443 ( .A(n_444), .Y(n_443) );
INVx1_ASAP7_75t_L g444 ( .A(n_445), .Y(n_444) );
INVx2_ASAP7_75t_L g446 ( .A(n_447), .Y(n_446) );
HB1xp67_ASAP7_75t_L g448 ( .A(n_449), .Y(n_448) );
INVx2_ASAP7_75t_L g450 ( .A(n_451), .Y(n_450) );
NOR2xp33_ASAP7_75t_L g472 ( .A(n_451), .B(n_473), .Y(n_472) );
OAI221xp5_ASAP7_75t_L g452 ( .A1(n_453), .A2(n_454), .B1(n_459), .B2(n_460), .C(n_461), .Y(n_452) );
OAI21xp33_ASAP7_75t_L g465 ( .A1(n_453), .A2(n_466), .B(n_468), .Y(n_465) );
INVxp67_ASAP7_75t_L g454 ( .A(n_455), .Y(n_454) );
INVx2_ASAP7_75t_L g455 ( .A(n_456), .Y(n_455) );
OR2x2_ASAP7_75t_L g456 ( .A(n_457), .B(n_458), .Y(n_456) );
INVx1_ASAP7_75t_L g466 ( .A(n_467), .Y(n_466) );
INVx1_ASAP7_75t_L g481 ( .A(n_473), .Y(n_481) );
AOI211xp5_ASAP7_75t_L g474 ( .A1(n_475), .A2(n_476), .B(n_477), .C(n_490), .Y(n_474) );
OAI21xp5_ASAP7_75t_SL g477 ( .A1(n_478), .A2(n_479), .B(n_484), .Y(n_477) );
INVx1_ASAP7_75t_L g479 ( .A(n_480), .Y(n_479) );
NOR2x1_ASAP7_75t_L g480 ( .A(n_481), .B(n_482), .Y(n_480) );
HB1xp67_ASAP7_75t_L g491 ( .A(n_482), .Y(n_491) );
INVx1_ASAP7_75t_L g485 ( .A(n_486), .Y(n_485) );
INVx1_ASAP7_75t_L g487 ( .A(n_488), .Y(n_487) );
INVx1_ASAP7_75t_L g494 ( .A(n_495), .Y(n_494) );
NOR2x1_ASAP7_75t_L g497 ( .A(n_498), .B(n_700), .Y(n_497) );
NAND3xp33_ASAP7_75t_L g498 ( .A(n_499), .B(n_630), .C(n_676), .Y(n_498) );
AOI221x1_ASAP7_75t_L g499 ( .A1(n_500), .A2(n_550), .B1(n_588), .B2(n_591), .C(n_610), .Y(n_499) );
INVx1_ASAP7_75t_L g500 ( .A(n_501), .Y(n_500) );
NAND2xp5_ASAP7_75t_L g501 ( .A(n_502), .B(n_525), .Y(n_501) );
AND2x2_ASAP7_75t_L g589 ( .A(n_502), .B(n_590), .Y(n_589) );
INVx1_ASAP7_75t_L g728 ( .A(n_502), .Y(n_728) );
NAND2xp5_ASAP7_75t_L g829 ( .A(n_502), .B(n_692), .Y(n_829) );
AND2x2_ASAP7_75t_L g502 ( .A(n_503), .B(n_514), .Y(n_502) );
INVx1_ASAP7_75t_L g691 ( .A(n_503), .Y(n_691) );
INVx1_ASAP7_75t_L g503 ( .A(n_504), .Y(n_503) );
AND2x2_ASAP7_75t_L g634 ( .A(n_504), .B(n_635), .Y(n_634) );
AND2x2_ASAP7_75t_L g671 ( .A(n_504), .B(n_528), .Y(n_671) );
OR2x2_ASAP7_75t_L g727 ( .A(n_504), .B(n_528), .Y(n_727) );
INVx1_ASAP7_75t_L g626 ( .A(n_514), .Y(n_626) );
BUFx3_ASAP7_75t_L g648 ( .A(n_514), .Y(n_648) );
INVxp67_ASAP7_75t_SL g680 ( .A(n_514), .Y(n_680) );
AND2x2_ASAP7_75t_L g726 ( .A(n_514), .B(n_667), .Y(n_726) );
AND2x2_ASAP7_75t_L g743 ( .A(n_514), .B(n_539), .Y(n_743) );
INVx1_ASAP7_75t_L g790 ( .A(n_514), .Y(n_790) );
INVxp67_ASAP7_75t_SL g798 ( .A(n_514), .Y(n_798) );
INVx3_ASAP7_75t_L g514 ( .A(n_515), .Y(n_514) );
INVx1_ASAP7_75t_L g525 ( .A(n_526), .Y(n_525) );
INVx1_ASAP7_75t_L g526 ( .A(n_527), .Y(n_526) );
INVx2_ASAP7_75t_L g590 ( .A(n_527), .Y(n_590) );
OR2x2_ASAP7_75t_L g793 ( .A(n_527), .B(n_683), .Y(n_793) );
HB1xp67_ASAP7_75t_L g825 ( .A(n_527), .Y(n_825) );
OR2x2_ASAP7_75t_L g527 ( .A(n_528), .B(n_539), .Y(n_527) );
AND2x2_ASAP7_75t_L g627 ( .A(n_528), .B(n_628), .Y(n_627) );
INVx1_ASAP7_75t_L g635 ( .A(n_528), .Y(n_635) );
NAND2xp5_ASAP7_75t_L g647 ( .A(n_528), .B(n_539), .Y(n_647) );
AND2x2_ASAP7_75t_L g692 ( .A(n_528), .B(n_667), .Y(n_692) );
HB1xp67_ASAP7_75t_L g719 ( .A(n_528), .Y(n_719) );
INVx2_ASAP7_75t_L g532 ( .A(n_533), .Y(n_532) );
NAND2xp5_ASAP7_75t_L g583 ( .A(n_535), .B(n_584), .Y(n_583) );
INVx2_ASAP7_75t_L g578 ( .A(n_536), .Y(n_578) );
AND2x2_ASAP7_75t_L g669 ( .A(n_539), .B(n_670), .Y(n_669) );
NAND2x1p5_ASAP7_75t_L g802 ( .A(n_550), .B(n_621), .Y(n_802) );
AND2x2_ASAP7_75t_L g550 ( .A(n_551), .B(n_565), .Y(n_550) );
BUFx2_ASAP7_75t_L g762 ( .A(n_551), .Y(n_762) );
INVx1_ASAP7_75t_L g551 ( .A(n_552), .Y(n_551) );
AND2x2_ASAP7_75t_L g613 ( .A(n_552), .B(n_614), .Y(n_613) );
NAND2xp5_ASAP7_75t_SL g714 ( .A(n_552), .B(n_652), .Y(n_714) );
AND2x2_ASAP7_75t_L g758 ( .A(n_552), .B(n_618), .Y(n_758) );
INVx2_ASAP7_75t_L g552 ( .A(n_553), .Y(n_552) );
OR2x2_ASAP7_75t_L g597 ( .A(n_553), .B(n_598), .Y(n_597) );
NAND2x1_ASAP7_75t_L g643 ( .A(n_553), .B(n_644), .Y(n_643) );
AND2x2_ASAP7_75t_L g822 ( .A(n_553), .B(n_652), .Y(n_822) );
INVx4_ASAP7_75t_L g553 ( .A(n_554), .Y(n_553) );
BUFx2_ASAP7_75t_L g637 ( .A(n_554), .Y(n_637) );
INVx1_ASAP7_75t_L g660 ( .A(n_554), .Y(n_660) );
AND2x2_ASAP7_75t_L g675 ( .A(n_554), .B(n_645), .Y(n_675) );
OR2x2_ASAP7_75t_L g736 ( .A(n_554), .B(n_623), .Y(n_736) );
AND2x4_ASAP7_75t_L g554 ( .A(n_555), .B(n_556), .Y(n_554) );
OAI21x1_ASAP7_75t_L g556 ( .A1(n_557), .A2(n_560), .B(n_564), .Y(n_556) );
AND2x2_ASAP7_75t_L g732 ( .A(n_565), .B(n_659), .Y(n_732) );
NAND2xp5_ASAP7_75t_L g785 ( .A(n_565), .B(n_688), .Y(n_785) );
AND2x2_ASAP7_75t_L g565 ( .A(n_566), .B(n_575), .Y(n_565) );
BUFx2_ASAP7_75t_L g765 ( .A(n_566), .Y(n_765) );
AND2x2_ASAP7_75t_L g722 ( .A(n_575), .B(n_645), .Y(n_722) );
INVx1_ASAP7_75t_L g575 ( .A(n_576), .Y(n_575) );
INVx2_ASAP7_75t_L g595 ( .A(n_576), .Y(n_595) );
AND2x2_ASAP7_75t_L g639 ( .A(n_576), .B(n_600), .Y(n_639) );
AOI21x1_ASAP7_75t_L g576 ( .A1(n_577), .A2(n_579), .B(n_587), .Y(n_576) );
NAND2xp5_ASAP7_75t_L g579 ( .A(n_580), .B(n_583), .Y(n_579) );
HB1xp67_ASAP7_75t_L g588 ( .A(n_589), .Y(n_588) );
INVx1_ASAP7_75t_L g654 ( .A(n_590), .Y(n_654) );
AND2x4_ASAP7_75t_L g817 ( .A(n_590), .B(n_818), .Y(n_817) );
INVx1_ASAP7_75t_L g591 ( .A(n_592), .Y(n_591) );
INVx2_ASAP7_75t_L g592 ( .A(n_593), .Y(n_592) );
AND2x2_ASAP7_75t_L g593 ( .A(n_594), .B(n_596), .Y(n_593) );
NAND2xp5_ASAP7_75t_L g619 ( .A(n_594), .B(n_620), .Y(n_619) );
INVx2_ASAP7_75t_L g658 ( .A(n_594), .Y(n_658) );
AND2x2_ASAP7_75t_L g707 ( .A(n_594), .B(n_675), .Y(n_707) );
INVx2_ASAP7_75t_L g594 ( .A(n_595), .Y(n_594) );
AND2x2_ASAP7_75t_L g617 ( .A(n_595), .B(n_618), .Y(n_617) );
INVx2_ASAP7_75t_L g652 ( .A(n_595), .Y(n_652) );
INVx1_ASAP7_75t_L g696 ( .A(n_595), .Y(n_696) );
INVx1_ASAP7_75t_SL g596 ( .A(n_597), .Y(n_596) );
INVx1_ASAP7_75t_L g653 ( .A(n_597), .Y(n_653) );
OR2x2_ASAP7_75t_L g720 ( .A(n_597), .B(n_721), .Y(n_720) );
OAI21xp33_ASAP7_75t_L g806 ( .A1(n_597), .A2(n_651), .B(n_736), .Y(n_806) );
INVx1_ASAP7_75t_L g598 ( .A(n_599), .Y(n_598) );
INVx2_ASAP7_75t_L g618 ( .A(n_599), .Y(n_618) );
AND2x2_ASAP7_75t_L g659 ( .A(n_599), .B(n_660), .Y(n_659) );
HB1xp67_ASAP7_75t_L g688 ( .A(n_599), .Y(n_688) );
INVx2_ASAP7_75t_L g599 ( .A(n_600), .Y(n_599) );
INVx1_ASAP7_75t_L g623 ( .A(n_600), .Y(n_623) );
OAI21x1_ASAP7_75t_L g600 ( .A1(n_601), .A2(n_602), .B(n_609), .Y(n_600) );
AOI21xp5_ASAP7_75t_L g610 ( .A1(n_611), .A2(n_619), .B(n_624), .Y(n_610) );
INVx3_ASAP7_75t_L g611 ( .A(n_612), .Y(n_611) );
AOI22xp5_ASAP7_75t_L g827 ( .A1(n_612), .A2(n_690), .B1(n_828), .B2(n_830), .Y(n_827) );
AND2x4_ASAP7_75t_L g612 ( .A(n_613), .B(n_617), .Y(n_612) );
O2A1O1Ixp33_ASAP7_75t_L g676 ( .A1(n_613), .A2(n_639), .B(n_677), .C(n_685), .Y(n_676) );
INVx1_ASAP7_75t_L g787 ( .A(n_613), .Y(n_787) );
AND2x2_ASAP7_75t_L g638 ( .A(n_614), .B(n_639), .Y(n_638) );
AND2x2_ASAP7_75t_L g651 ( .A(n_614), .B(n_652), .Y(n_651) );
INVx2_ASAP7_75t_L g614 ( .A(n_615), .Y(n_614) );
AND2x2_ASAP7_75t_L g745 ( .A(n_615), .B(n_623), .Y(n_745) );
INVx1_ASAP7_75t_L g615 ( .A(n_616), .Y(n_615) );
INVx2_ASAP7_75t_L g645 ( .A(n_616), .Y(n_645) );
AND2x2_ASAP7_75t_L g807 ( .A(n_618), .B(n_722), .Y(n_807) );
INVx1_ASAP7_75t_L g620 ( .A(n_621), .Y(n_620) );
BUFx2_ASAP7_75t_L g621 ( .A(n_622), .Y(n_621) );
INVxp67_ASAP7_75t_L g622 ( .A(n_623), .Y(n_622) );
HB1xp67_ASAP7_75t_L g673 ( .A(n_623), .Y(n_673) );
OR2x2_ASAP7_75t_L g705 ( .A(n_623), .B(n_706), .Y(n_705) );
INVx1_ASAP7_75t_L g624 ( .A(n_625), .Y(n_624) );
AND2x2_ASAP7_75t_L g625 ( .A(n_626), .B(n_627), .Y(n_625) );
INVx1_ASAP7_75t_L g716 ( .A(n_626), .Y(n_716) );
AND2x4_ASAP7_75t_L g729 ( .A(n_626), .B(n_665), .Y(n_729) );
BUFx2_ASAP7_75t_L g663 ( .A(n_628), .Y(n_663) );
INVx1_ASAP7_75t_L g628 ( .A(n_629), .Y(n_628) );
BUFx3_ASAP7_75t_L g684 ( .A(n_629), .Y(n_684) );
AOI211xp5_ASAP7_75t_L g630 ( .A1(n_631), .A2(n_636), .B(n_640), .C(n_655), .Y(n_630) );
INVx1_ASAP7_75t_L g631 ( .A(n_632), .Y(n_631) );
INVx1_ASAP7_75t_L g632 ( .A(n_633), .Y(n_632) );
HB1xp67_ASAP7_75t_L g633 ( .A(n_634), .Y(n_633) );
AND2x2_ASAP7_75t_L g801 ( .A(n_634), .B(n_783), .Y(n_801) );
NAND2xp5_ASAP7_75t_L g810 ( .A(n_634), .B(n_789), .Y(n_810) );
AND2x4_ASAP7_75t_L g665 ( .A(n_635), .B(n_666), .Y(n_665) );
AND2x4_ASAP7_75t_L g636 ( .A(n_637), .B(n_638), .Y(n_636) );
INVx2_ASAP7_75t_L g642 ( .A(n_639), .Y(n_642) );
OAI22xp5_ASAP7_75t_L g640 ( .A1(n_641), .A2(n_646), .B1(n_649), .B2(n_654), .Y(n_640) );
INVx1_ASAP7_75t_L g702 ( .A(n_641), .Y(n_702) );
OAI32xp33_ASAP7_75t_L g754 ( .A1(n_641), .A2(n_733), .A3(n_755), .B1(n_757), .B2(n_759), .Y(n_754) );
OAI22xp33_ASAP7_75t_L g815 ( .A1(n_641), .A2(n_793), .B1(n_816), .B2(n_819), .Y(n_815) );
OR2x6_ASAP7_75t_L g641 ( .A(n_642), .B(n_643), .Y(n_641) );
INVx1_ASAP7_75t_L g763 ( .A(n_642), .Y(n_763) );
INVx1_ASAP7_75t_SL g713 ( .A(n_644), .Y(n_713) );
NAND2xp5_ASAP7_75t_L g757 ( .A(n_644), .B(n_758), .Y(n_757) );
INVx2_ASAP7_75t_L g644 ( .A(n_645), .Y(n_644) );
OR2x2_ASAP7_75t_L g646 ( .A(n_647), .B(n_648), .Y(n_646) );
NAND2xp5_ASAP7_75t_L g699 ( .A(n_648), .B(n_692), .Y(n_699) );
NAND2xp5_ASAP7_75t_L g752 ( .A(n_648), .B(n_753), .Y(n_752) );
INVx1_ASAP7_75t_L g649 ( .A(n_650), .Y(n_649) );
A2O1A1O1Ixp25_ASAP7_75t_L g778 ( .A1(n_650), .A2(n_755), .B(n_779), .C(n_782), .D(n_784), .Y(n_778) );
AND2x2_ASAP7_75t_L g650 ( .A(n_651), .B(n_653), .Y(n_650) );
OAI22xp33_ASAP7_75t_L g655 ( .A1(n_656), .A2(n_661), .B1(n_668), .B2(n_672), .Y(n_655) );
INVx1_ASAP7_75t_L g656 ( .A(n_657), .Y(n_656) );
AND2x2_ASAP7_75t_L g657 ( .A(n_658), .B(n_659), .Y(n_657) );
AND2x2_ASAP7_75t_L g767 ( .A(n_659), .B(n_722), .Y(n_767) );
AND2x2_ASAP7_75t_L g782 ( .A(n_659), .B(n_783), .Y(n_782) );
INVx1_ASAP7_75t_L g811 ( .A(n_659), .Y(n_811) );
OR2x2_ASAP7_75t_L g661 ( .A(n_662), .B(n_664), .Y(n_661) );
AND2x2_ASAP7_75t_L g738 ( .A(n_662), .B(n_726), .Y(n_738) );
INVx2_ASAP7_75t_L g662 ( .A(n_663), .Y(n_662) );
AND2x2_ASAP7_75t_L g739 ( .A(n_663), .B(n_740), .Y(n_739) );
INVx2_ASAP7_75t_L g664 ( .A(n_665), .Y(n_664) );
AND2x4_ASAP7_75t_L g681 ( .A(n_665), .B(n_682), .Y(n_681) );
NOR2xp67_ASAP7_75t_L g753 ( .A(n_666), .B(n_684), .Y(n_753) );
INVx1_ASAP7_75t_L g666 ( .A(n_667), .Y(n_666) );
INVx1_ASAP7_75t_L g734 ( .A(n_667), .Y(n_734) );
AND2x2_ASAP7_75t_L g740 ( .A(n_667), .B(n_670), .Y(n_740) );
AND2x2_ASAP7_75t_L g799 ( .A(n_667), .B(n_684), .Y(n_799) );
NAND2xp5_ASAP7_75t_L g668 ( .A(n_669), .B(n_671), .Y(n_668) );
NAND2xp5_ASAP7_75t_L g776 ( .A(n_669), .B(n_777), .Y(n_776) );
INVx1_ASAP7_75t_L g706 ( .A(n_670), .Y(n_706) );
INVx1_ASAP7_75t_L g709 ( .A(n_671), .Y(n_709) );
AND2x2_ASAP7_75t_L g742 ( .A(n_671), .B(n_743), .Y(n_742) );
NAND2xp5_ASAP7_75t_L g786 ( .A(n_671), .B(n_734), .Y(n_786) );
NAND2xp5_ASAP7_75t_L g788 ( .A(n_671), .B(n_789), .Y(n_788) );
OR2x2_ASAP7_75t_L g672 ( .A(n_673), .B(n_674), .Y(n_672) );
INVx1_ASAP7_75t_L g674 ( .A(n_675), .Y(n_674) );
AND2x2_ASAP7_75t_L g687 ( .A(n_675), .B(n_688), .Y(n_687) );
AND2x2_ASAP7_75t_L g694 ( .A(n_675), .B(n_695), .Y(n_694) );
INVx1_ASAP7_75t_L g677 ( .A(n_678), .Y(n_677) );
NAND2x1_ASAP7_75t_L g678 ( .A(n_679), .B(n_681), .Y(n_678) );
NOR3x1_ASAP7_75t_L g824 ( .A(n_679), .B(n_825), .C(n_826), .Y(n_824) );
BUFx2_ASAP7_75t_L g679 ( .A(n_680), .Y(n_679) );
AND2x2_ASAP7_75t_L g769 ( .A(n_680), .B(n_692), .Y(n_769) );
INVx2_ASAP7_75t_L g774 ( .A(n_681), .Y(n_774) );
INVx2_ASAP7_75t_L g682 ( .A(n_683), .Y(n_682) );
AND2x2_ASAP7_75t_L g804 ( .A(n_683), .B(n_692), .Y(n_804) );
HB1xp67_ASAP7_75t_L g826 ( .A(n_683), .Y(n_826) );
INVx3_ASAP7_75t_L g683 ( .A(n_684), .Y(n_683) );
OAI22xp5_ASAP7_75t_L g685 ( .A1(n_686), .A2(n_689), .B1(n_693), .B2(n_697), .Y(n_685) );
INVx3_ASAP7_75t_L g686 ( .A(n_687), .Y(n_686) );
INVx2_ASAP7_75t_L g689 ( .A(n_690), .Y(n_689) );
AND2x2_ASAP7_75t_L g690 ( .A(n_691), .B(n_692), .Y(n_690) );
HB1xp67_ASAP7_75t_L g756 ( .A(n_691), .Y(n_756) );
INVx1_ASAP7_75t_L g818 ( .A(n_691), .Y(n_818) );
INVx1_ASAP7_75t_L g693 ( .A(n_694), .Y(n_693) );
NAND3xp33_ASAP7_75t_L g791 ( .A(n_694), .B(n_704), .C(n_792), .Y(n_791) );
OR2x2_ASAP7_75t_L g819 ( .A(n_695), .B(n_811), .Y(n_819) );
INVx1_ASAP7_75t_L g695 ( .A(n_696), .Y(n_695) );
HB1xp67_ASAP7_75t_L g781 ( .A(n_696), .Y(n_781) );
INVxp67_ASAP7_75t_L g697 ( .A(n_698), .Y(n_697) );
INVx1_ASAP7_75t_L g698 ( .A(n_699), .Y(n_698) );
NAND3xp33_ASAP7_75t_L g700 ( .A(n_701), .B(n_710), .C(n_746), .Y(n_700) );
OAI21xp33_ASAP7_75t_L g701 ( .A1(n_702), .A2(n_703), .B(n_708), .Y(n_701) );
AND2x2_ASAP7_75t_L g703 ( .A(n_704), .B(n_707), .Y(n_703) );
INVx1_ASAP7_75t_L g704 ( .A(n_705), .Y(n_704) );
INVx1_ASAP7_75t_L g783 ( .A(n_706), .Y(n_783) );
AOI22xp5_ASAP7_75t_L g772 ( .A1(n_707), .A2(n_749), .B1(n_773), .B2(n_775), .Y(n_772) );
INVx1_ASAP7_75t_L g708 ( .A(n_709), .Y(n_708) );
NOR2xp33_ASAP7_75t_L g710 ( .A(n_711), .B(n_730), .Y(n_710) );
OAI22xp33_ASAP7_75t_L g711 ( .A1(n_712), .A2(n_715), .B1(n_720), .B2(n_723), .Y(n_711) );
OR2x2_ASAP7_75t_L g712 ( .A(n_713), .B(n_714), .Y(n_712) );
NAND2xp5_ASAP7_75t_L g715 ( .A(n_716), .B(n_717), .Y(n_715) );
INVx1_ASAP7_75t_L g717 ( .A(n_718), .Y(n_717) );
INVx1_ASAP7_75t_L g718 ( .A(n_719), .Y(n_718) );
OR2x2_ASAP7_75t_L g735 ( .A(n_721), .B(n_736), .Y(n_735) );
INVx1_ASAP7_75t_L g749 ( .A(n_721), .Y(n_749) );
INVx2_ASAP7_75t_L g721 ( .A(n_722), .Y(n_721) );
NOR2xp67_ASAP7_75t_L g723 ( .A(n_724), .B(n_729), .Y(n_723) );
NAND3xp33_ASAP7_75t_L g724 ( .A(n_725), .B(n_727), .C(n_728), .Y(n_724) );
INVx2_ASAP7_75t_SL g725 ( .A(n_726), .Y(n_725) );
INVx1_ASAP7_75t_L g777 ( .A(n_727), .Y(n_777) );
INVx1_ASAP7_75t_L g814 ( .A(n_727), .Y(n_814) );
OAI222xp33_ASAP7_75t_L g730 ( .A1(n_731), .A2(n_733), .B1(n_735), .B2(n_737), .C1(n_741), .C2(n_744), .Y(n_730) );
INVx2_ASAP7_75t_L g731 ( .A(n_732), .Y(n_731) );
INVx2_ASAP7_75t_L g733 ( .A(n_734), .Y(n_733) );
AOI211xp5_ASAP7_75t_L g746 ( .A1(n_736), .A2(n_747), .B(n_754), .C(n_760), .Y(n_746) );
NOR2xp33_ASAP7_75t_SL g737 ( .A(n_738), .B(n_739), .Y(n_737) );
INVx2_ASAP7_75t_L g759 ( .A(n_739), .Y(n_759) );
INVx2_ASAP7_75t_L g741 ( .A(n_742), .Y(n_741) );
AOI21xp5_ASAP7_75t_L g805 ( .A1(n_744), .A2(n_806), .B(n_807), .Y(n_805) );
INVx1_ASAP7_75t_L g744 ( .A(n_745), .Y(n_744) );
NOR2xp33_ASAP7_75t_L g747 ( .A(n_748), .B(n_750), .Y(n_747) );
INVx1_ASAP7_75t_L g748 ( .A(n_749), .Y(n_748) );
INVx1_ASAP7_75t_L g750 ( .A(n_751), .Y(n_750) );
INVx1_ASAP7_75t_L g751 ( .A(n_752), .Y(n_751) );
INVx1_ASAP7_75t_L g755 ( .A(n_756), .Y(n_755) );
AND2x2_ASAP7_75t_L g830 ( .A(n_758), .B(n_781), .Y(n_830) );
AOI21xp33_ASAP7_75t_L g760 ( .A1(n_761), .A2(n_766), .B(n_768), .Y(n_760) );
NAND3x2_ASAP7_75t_L g761 ( .A(n_762), .B(n_763), .C(n_764), .Y(n_761) );
INVx2_ASAP7_75t_L g764 ( .A(n_765), .Y(n_764) );
AO21x1_ASAP7_75t_L g808 ( .A1(n_765), .A2(n_809), .B(n_815), .Y(n_808) );
INVx1_ASAP7_75t_L g766 ( .A(n_767), .Y(n_766) );
INVxp67_ASAP7_75t_SL g768 ( .A(n_769), .Y(n_768) );
NOR4xp75_ASAP7_75t_L g770 ( .A(n_771), .B(n_794), .C(n_808), .D(n_820), .Y(n_770) );
NAND3x1_ASAP7_75t_L g771 ( .A(n_772), .B(n_778), .C(n_791), .Y(n_771) );
INVx2_ASAP7_75t_L g773 ( .A(n_774), .Y(n_773) );
INVx1_ASAP7_75t_L g775 ( .A(n_776), .Y(n_775) );
INVx1_ASAP7_75t_L g779 ( .A(n_780), .Y(n_779) );
INVx1_ASAP7_75t_L g780 ( .A(n_781), .Y(n_780) );
INVx1_ASAP7_75t_L g812 ( .A(n_782), .Y(n_812) );
OAI22xp33_ASAP7_75t_SL g784 ( .A1(n_785), .A2(n_786), .B1(n_787), .B2(n_788), .Y(n_784) );
INVx1_ASAP7_75t_L g789 ( .A(n_790), .Y(n_789) );
OR2x2_ASAP7_75t_L g800 ( .A(n_792), .B(n_801), .Y(n_800) );
INVx2_ASAP7_75t_L g792 ( .A(n_793), .Y(n_792) );
OAI22xp5_ASAP7_75t_L g794 ( .A1(n_795), .A2(n_802), .B1(n_803), .B2(n_805), .Y(n_794) );
NOR2x1_ASAP7_75t_L g795 ( .A(n_796), .B(n_800), .Y(n_795) );
BUFx2_ASAP7_75t_L g796 ( .A(n_797), .Y(n_796) );
AND2x4_ASAP7_75t_L g797 ( .A(n_798), .B(n_799), .Y(n_797) );
INVx2_ASAP7_75t_L g803 ( .A(n_804), .Y(n_803) );
OAI22xp5_ASAP7_75t_L g809 ( .A1(n_810), .A2(n_811), .B1(n_812), .B2(n_813), .Y(n_809) );
INVx1_ASAP7_75t_L g813 ( .A(n_814), .Y(n_813) );
INVx1_ASAP7_75t_L g816 ( .A(n_817), .Y(n_816) );
OAI21xp33_ASAP7_75t_SL g820 ( .A1(n_821), .A2(n_823), .B(n_827), .Y(n_820) );
INVx1_ASAP7_75t_L g821 ( .A(n_822), .Y(n_821) );
INVx2_ASAP7_75t_L g823 ( .A(n_824), .Y(n_823) );
INVx1_ASAP7_75t_L g828 ( .A(n_829), .Y(n_828) );
AOI21xp5_ASAP7_75t_L g834 ( .A1(n_835), .A2(n_836), .B(n_837), .Y(n_834) );
NAND2xp5_ASAP7_75t_SL g837 ( .A(n_838), .B(n_846), .Y(n_837) );
INVx1_ASAP7_75t_L g839 ( .A(n_840), .Y(n_839) );
INVx2_ASAP7_75t_L g840 ( .A(n_841), .Y(n_840) );
BUFx10_ASAP7_75t_L g841 ( .A(n_842), .Y(n_841) );
INVx1_ASAP7_75t_L g843 ( .A(n_844), .Y(n_843) );
OAI21xp5_ASAP7_75t_L g872 ( .A1(n_846), .A2(n_868), .B(n_873), .Y(n_872) );
INVx1_ASAP7_75t_L g846 ( .A(n_847), .Y(n_846) );
NOR2xp33_ASAP7_75t_L g847 ( .A(n_848), .B(n_849), .Y(n_847) );
BUFx12f_ASAP7_75t_L g849 ( .A(n_850), .Y(n_849) );
INVx4_ASAP7_75t_L g850 ( .A(n_851), .Y(n_850) );
CKINVDCx5p33_ASAP7_75t_R g874 ( .A(n_851), .Y(n_874) );
INVx1_ASAP7_75t_L g853 ( .A(n_854), .Y(n_853) );
HB1xp67_ASAP7_75t_L g866 ( .A(n_854), .Y(n_866) );
NOR2xp67_ASAP7_75t_L g855 ( .A(n_856), .B(n_860), .Y(n_855) );
INVx1_ASAP7_75t_L g856 ( .A(n_857), .Y(n_856) );
BUFx2_ASAP7_75t_L g857 ( .A(n_858), .Y(n_857) );
INVx2_ASAP7_75t_L g858 ( .A(n_859), .Y(n_858) );
AOI21x1_ASAP7_75t_L g860 ( .A1(n_861), .A2(n_862), .B(n_872), .Y(n_860) );
INVx1_ASAP7_75t_L g862 ( .A(n_863), .Y(n_862) );
NAND2xp5_ASAP7_75t_L g863 ( .A(n_864), .B(n_868), .Y(n_863) );
INVx4_ASAP7_75t_L g864 ( .A(n_865), .Y(n_864) );
NAND2xp5_ASAP7_75t_L g882 ( .A(n_866), .B(n_883), .Y(n_882) );
NAND2xp5_ASAP7_75t_L g884 ( .A(n_867), .B(n_885), .Y(n_884) );
INVx3_ASAP7_75t_SL g875 ( .A(n_876), .Y(n_875) );
OR2x6_ASAP7_75t_L g876 ( .A(n_877), .B(n_882), .Y(n_876) );
OR2x6_ASAP7_75t_L g889 ( .A(n_877), .B(n_882), .Y(n_889) );
INVx1_ASAP7_75t_L g877 ( .A(n_878), .Y(n_877) );
NOR2x1p5_ASAP7_75t_L g878 ( .A(n_879), .B(n_880), .Y(n_878) );
INVx1_ASAP7_75t_L g880 ( .A(n_881), .Y(n_880) );
INVx1_ASAP7_75t_L g883 ( .A(n_884), .Y(n_883) );
INVx1_ASAP7_75t_L g887 ( .A(n_888), .Y(n_887) );
INVx1_ASAP7_75t_L g888 ( .A(n_889), .Y(n_888) );
endmodule