module fake_jpeg_12547_n_266 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_266);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_266;

wire n_159;
wire n_117;
wire n_253;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_84;
wire n_59;
wire n_98;
wire n_252;
wire n_251;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_223;
wire n_234;
wire n_171;
wire n_263;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_44;
wire n_24;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_121;
wire n_99;
wire n_130;
wire n_102;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_262;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_216;
wire n_217;
wire n_264;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_48;
wire n_35;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_265;
wire n_176;
wire n_199;
wire n_112;
wire n_260;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_258;
wire n_96;

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_15),
.Y(n_16)
);

BUFx6f_ASAP7_75t_L g17 ( 
.A(n_15),
.Y(n_17)
);

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_1),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_14),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_12),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_1),
.Y(n_21)
);

INVx3_ASAP7_75t_L g22 ( 
.A(n_7),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_3),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_13),
.Y(n_24)
);

INVx6_ASAP7_75t_L g25 ( 
.A(n_9),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_13),
.Y(n_26)
);

BUFx12_ASAP7_75t_L g27 ( 
.A(n_3),
.Y(n_27)
);

BUFx10_ASAP7_75t_L g28 ( 
.A(n_11),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_2),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_8),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_2),
.Y(n_31)
);

INVx8_ASAP7_75t_L g32 ( 
.A(n_8),
.Y(n_32)
);

CKINVDCx16_ASAP7_75t_R g33 ( 
.A(n_8),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_4),
.Y(n_34)
);

INVx6_ASAP7_75t_L g35 ( 
.A(n_10),
.Y(n_35)
);

BUFx12f_ASAP7_75t_L g36 ( 
.A(n_13),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_2),
.Y(n_37)
);

INVx13_ASAP7_75t_L g38 ( 
.A(n_7),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_10),
.Y(n_39)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_3),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_11),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_6),
.Y(n_42)
);

BUFx3_ASAP7_75t_L g43 ( 
.A(n_36),
.Y(n_43)
);

BUFx12f_ASAP7_75t_L g126 ( 
.A(n_43),
.Y(n_126)
);

BUFx12f_ASAP7_75t_L g44 ( 
.A(n_28),
.Y(n_44)
);

INVx5_ASAP7_75t_L g92 ( 
.A(n_44),
.Y(n_92)
);

BUFx3_ASAP7_75t_L g45 ( 
.A(n_36),
.Y(n_45)
);

INVx5_ASAP7_75t_L g122 ( 
.A(n_45),
.Y(n_122)
);

INVx2_ASAP7_75t_L g46 ( 
.A(n_36),
.Y(n_46)
);

INVx2_ASAP7_75t_L g123 ( 
.A(n_46),
.Y(n_123)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_18),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g101 ( 
.A(n_47),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_16),
.B(n_41),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_SL g87 ( 
.A(n_48),
.B(n_66),
.Y(n_87)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_18),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g111 ( 
.A(n_49),
.Y(n_111)
);

BUFx3_ASAP7_75t_L g50 ( 
.A(n_36),
.Y(n_50)
);

INVx4_ASAP7_75t_L g90 ( 
.A(n_50),
.Y(n_90)
);

INVx5_ASAP7_75t_L g51 ( 
.A(n_32),
.Y(n_51)
);

INVx3_ASAP7_75t_L g94 ( 
.A(n_51),
.Y(n_94)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_18),
.Y(n_52)
);

INVx6_ASAP7_75t_L g91 ( 
.A(n_52),
.Y(n_91)
);

BUFx5_ASAP7_75t_L g53 ( 
.A(n_28),
.Y(n_53)
);

BUFx8_ASAP7_75t_L g103 ( 
.A(n_53),
.Y(n_103)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_21),
.Y(n_54)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_54),
.Y(n_128)
);

BUFx12f_ASAP7_75t_L g55 ( 
.A(n_28),
.Y(n_55)
);

INVx3_ASAP7_75t_L g102 ( 
.A(n_55),
.Y(n_102)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_21),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_56),
.B(n_61),
.Y(n_99)
);

BUFx12f_ASAP7_75t_L g57 ( 
.A(n_28),
.Y(n_57)
);

INVx3_ASAP7_75t_L g113 ( 
.A(n_57),
.Y(n_113)
);

INVx2_ASAP7_75t_SL g58 ( 
.A(n_22),
.Y(n_58)
);

AND2x2_ASAP7_75t_L g88 ( 
.A(n_58),
.B(n_64),
.Y(n_88)
);

BUFx12f_ASAP7_75t_L g59 ( 
.A(n_23),
.Y(n_59)
);

INVx3_ASAP7_75t_L g117 ( 
.A(n_59),
.Y(n_117)
);

INVx4_ASAP7_75t_L g60 ( 
.A(n_22),
.Y(n_60)
);

INVx2_ASAP7_75t_L g124 ( 
.A(n_60),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_SL g61 ( 
.A(n_16),
.B(n_14),
.Y(n_61)
);

INVx8_ASAP7_75t_L g62 ( 
.A(n_23),
.Y(n_62)
);

INVx6_ASAP7_75t_L g93 ( 
.A(n_62),
.Y(n_93)
);

BUFx24_ASAP7_75t_L g63 ( 
.A(n_38),
.Y(n_63)
);

INVx11_ASAP7_75t_L g118 ( 
.A(n_63),
.Y(n_118)
);

AOI21xp33_ASAP7_75t_L g64 ( 
.A1(n_20),
.A2(n_0),
.B(n_1),
.Y(n_64)
);

INVx2_ASAP7_75t_L g65 ( 
.A(n_35),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_L g96 ( 
.A(n_65),
.B(n_68),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_20),
.B(n_0),
.Y(n_66)
);

INVx8_ASAP7_75t_L g67 ( 
.A(n_23),
.Y(n_67)
);

INVx6_ASAP7_75t_L g115 ( 
.A(n_67),
.Y(n_115)
);

INVx2_ASAP7_75t_L g68 ( 
.A(n_35),
.Y(n_68)
);

BUFx12f_ASAP7_75t_L g69 ( 
.A(n_26),
.Y(n_69)
);

INVx6_ASAP7_75t_L g121 ( 
.A(n_69),
.Y(n_121)
);

CKINVDCx20_ASAP7_75t_R g70 ( 
.A(n_27),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_70),
.B(n_71),
.Y(n_105)
);

BUFx12f_ASAP7_75t_L g71 ( 
.A(n_26),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_29),
.B(n_0),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_SL g89 ( 
.A(n_72),
.B(n_73),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_29),
.B(n_4),
.Y(n_73)
);

BUFx6f_ASAP7_75t_L g74 ( 
.A(n_26),
.Y(n_74)
);

INVx8_ASAP7_75t_L g129 ( 
.A(n_74),
.Y(n_129)
);

INVx11_ASAP7_75t_L g75 ( 
.A(n_38),
.Y(n_75)
);

CKINVDCx20_ASAP7_75t_R g86 ( 
.A(n_75),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_L g76 ( 
.A(n_30),
.B(n_42),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_L g100 ( 
.A(n_76),
.B(n_77),
.Y(n_100)
);

BUFx6f_ASAP7_75t_L g77 ( 
.A(n_31),
.Y(n_77)
);

INVx2_ASAP7_75t_L g78 ( 
.A(n_35),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_L g104 ( 
.A(n_78),
.B(n_80),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_30),
.B(n_41),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_SL g98 ( 
.A(n_79),
.B(n_84),
.Y(n_98)
);

BUFx6f_ASAP7_75t_L g80 ( 
.A(n_31),
.Y(n_80)
);

INVx2_ASAP7_75t_L g81 ( 
.A(n_31),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g110 ( 
.A(n_81),
.B(n_82),
.Y(n_110)
);

BUFx6f_ASAP7_75t_L g82 ( 
.A(n_39),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_L g83 ( 
.A(n_37),
.B(n_4),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g120 ( 
.A(n_83),
.B(n_33),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_37),
.B(n_5),
.Y(n_84)
);

OAI22xp5_ASAP7_75t_SL g85 ( 
.A1(n_47),
.A2(n_19),
.B1(n_17),
.B2(n_25),
.Y(n_85)
);

AOI22xp33_ASAP7_75t_L g142 ( 
.A1(n_85),
.A2(n_82),
.B1(n_80),
.B2(n_77),
.Y(n_142)
);

AOI22xp33_ASAP7_75t_SL g95 ( 
.A1(n_63),
.A2(n_32),
.B1(n_25),
.B2(n_39),
.Y(n_95)
);

AOI21xp5_ASAP7_75t_L g135 ( 
.A1(n_95),
.A2(n_97),
.B(n_62),
.Y(n_135)
);

AOI22xp33_ASAP7_75t_SL g97 ( 
.A1(n_63),
.A2(n_32),
.B1(n_39),
.B2(n_19),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g106 ( 
.A(n_44),
.B(n_42),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_SL g139 ( 
.A(n_106),
.B(n_107),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_44),
.B(n_34),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_55),
.B(n_40),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_L g148 ( 
.A(n_108),
.B(n_109),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_SL g109 ( 
.A(n_58),
.B(n_34),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_SL g112 ( 
.A(n_43),
.B(n_40),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_L g150 ( 
.A(n_112),
.B(n_114),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_L g114 ( 
.A(n_55),
.B(n_24),
.Y(n_114)
);

AOI22xp33_ASAP7_75t_L g116 ( 
.A1(n_49),
.A2(n_33),
.B1(n_19),
.B2(n_17),
.Y(n_116)
);

OAI22xp5_ASAP7_75t_L g145 ( 
.A1(n_116),
.A2(n_127),
.B1(n_67),
.B2(n_74),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_L g119 ( 
.A(n_57),
.B(n_24),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_L g154 ( 
.A(n_119),
.B(n_120),
.Y(n_154)
);

NOR2xp33_ASAP7_75t_L g125 ( 
.A(n_57),
.B(n_17),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_L g159 ( 
.A(n_125),
.B(n_5),
.Y(n_159)
);

AOI22xp33_ASAP7_75t_L g127 ( 
.A1(n_52),
.A2(n_38),
.B1(n_27),
.B2(n_7),
.Y(n_127)
);

BUFx6f_ASAP7_75t_L g130 ( 
.A(n_101),
.Y(n_130)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_130),
.Y(n_168)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_128),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_L g169 ( 
.A(n_131),
.B(n_133),
.Y(n_169)
);

AND2x2_ASAP7_75t_L g132 ( 
.A(n_100),
.B(n_71),
.Y(n_132)
);

INVxp67_ASAP7_75t_L g177 ( 
.A(n_132),
.Y(n_177)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_105),
.Y(n_133)
);

INVx3_ASAP7_75t_L g134 ( 
.A(n_118),
.Y(n_134)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_134),
.Y(n_180)
);

AOI22xp33_ASAP7_75t_SL g173 ( 
.A1(n_135),
.A2(n_161),
.B1(n_166),
.B2(n_129),
.Y(n_173)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_123),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_L g178 ( 
.A(n_136),
.B(n_137),
.Y(n_178)
);

INVxp67_ASAP7_75t_L g137 ( 
.A(n_118),
.Y(n_137)
);

INVx3_ASAP7_75t_L g138 ( 
.A(n_121),
.Y(n_138)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_138),
.Y(n_181)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_124),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_L g182 ( 
.A(n_140),
.B(n_143),
.Y(n_182)
);

HB1xp67_ASAP7_75t_L g141 ( 
.A(n_90),
.Y(n_141)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_141),
.Y(n_185)
);

OAI22xp5_ASAP7_75t_L g179 ( 
.A1(n_142),
.A2(n_115),
.B1(n_121),
.B2(n_92),
.Y(n_179)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_94),
.Y(n_143)
);

INVx2_ASAP7_75t_L g144 ( 
.A(n_91),
.Y(n_144)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_144),
.Y(n_191)
);

AOI22xp5_ASAP7_75t_L g175 ( 
.A1(n_145),
.A2(n_158),
.B1(n_163),
.B2(n_111),
.Y(n_175)
);

INVxp67_ASAP7_75t_L g146 ( 
.A(n_95),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_L g193 ( 
.A(n_146),
.B(n_151),
.Y(n_193)
);

AOI32xp33_ASAP7_75t_L g147 ( 
.A1(n_88),
.A2(n_71),
.A3(n_69),
.B1(n_59),
.B2(n_10),
.Y(n_147)
);

AOI32xp33_ASAP7_75t_L g171 ( 
.A1(n_147),
.A2(n_126),
.A3(n_103),
.B1(n_122),
.B2(n_129),
.Y(n_171)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_96),
.Y(n_149)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_149),
.Y(n_192)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_117),
.Y(n_151)
);

A2O1A1Ixp33_ASAP7_75t_L g152 ( 
.A1(n_88),
.A2(n_5),
.B(n_6),
.C(n_9),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_SL g183 ( 
.A(n_152),
.B(n_157),
.Y(n_183)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_117),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_L g172 ( 
.A(n_153),
.B(n_155),
.Y(n_172)
);

INVx6_ASAP7_75t_L g155 ( 
.A(n_91),
.Y(n_155)
);

AND2x2_ASAP7_75t_SL g156 ( 
.A(n_104),
.B(n_69),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_SL g176 ( 
.A(n_156),
.B(n_132),
.Y(n_176)
);

NAND2xp33_ASAP7_75t_L g157 ( 
.A(n_89),
.B(n_27),
.Y(n_157)
);

OAI22xp5_ASAP7_75t_SL g158 ( 
.A1(n_116),
.A2(n_59),
.B1(n_27),
.B2(n_9),
.Y(n_158)
);

NAND3xp33_ASAP7_75t_L g174 ( 
.A(n_159),
.B(n_162),
.C(n_99),
.Y(n_174)
);

INVx2_ASAP7_75t_L g160 ( 
.A(n_101),
.Y(n_160)
);

NOR2xp33_ASAP7_75t_L g190 ( 
.A(n_160),
.B(n_165),
.Y(n_190)
);

AOI22xp33_ASAP7_75t_SL g161 ( 
.A1(n_93),
.A2(n_115),
.B1(n_90),
.B2(n_122),
.Y(n_161)
);

INVxp67_ASAP7_75t_L g162 ( 
.A(n_97),
.Y(n_162)
);

OAI22xp5_ASAP7_75t_SL g163 ( 
.A1(n_110),
.A2(n_6),
.B1(n_11),
.B2(n_12),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_L g164 ( 
.A(n_98),
.B(n_12),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_L g187 ( 
.A(n_164),
.B(n_167),
.Y(n_187)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_93),
.Y(n_165)
);

INVx2_ASAP7_75t_L g166 ( 
.A(n_111),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_L g167 ( 
.A(n_87),
.B(n_86),
.Y(n_167)
);

OR2x2_ASAP7_75t_L g170 ( 
.A(n_149),
.B(n_127),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_L g207 ( 
.A(n_170),
.B(n_192),
.Y(n_207)
);

OAI22xp5_ASAP7_75t_L g210 ( 
.A1(n_171),
.A2(n_175),
.B1(n_189),
.B2(n_170),
.Y(n_210)
);

INVxp67_ASAP7_75t_L g208 ( 
.A(n_173),
.Y(n_208)
);

NOR2xp33_ASAP7_75t_L g199 ( 
.A(n_174),
.B(n_130),
.Y(n_199)
);

NOR2xp67_ASAP7_75t_SL g198 ( 
.A(n_176),
.B(n_138),
.Y(n_198)
);

AOI22xp5_ASAP7_75t_L g213 ( 
.A1(n_179),
.A2(n_186),
.B1(n_194),
.B2(n_180),
.Y(n_213)
);

NAND2xp5_ASAP7_75t_SL g184 ( 
.A(n_167),
.B(n_113),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_SL g202 ( 
.A(n_184),
.B(n_195),
.Y(n_202)
);

OAI22xp5_ASAP7_75t_L g186 ( 
.A1(n_162),
.A2(n_102),
.B1(n_113),
.B2(n_92),
.Y(n_186)
);

NOR2xp33_ASAP7_75t_SL g188 ( 
.A(n_154),
.B(n_126),
.Y(n_188)
);

NOR2xp33_ASAP7_75t_SL g203 ( 
.A(n_188),
.B(n_160),
.Y(n_203)
);

AOI22xp33_ASAP7_75t_L g189 ( 
.A1(n_146),
.A2(n_103),
.B1(n_126),
.B2(n_158),
.Y(n_189)
);

OAI22xp5_ASAP7_75t_SL g194 ( 
.A1(n_135),
.A2(n_103),
.B1(n_148),
.B2(n_156),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_SL g195 ( 
.A(n_132),
.B(n_150),
.Y(n_195)
);

O2A1O1Ixp33_ASAP7_75t_L g196 ( 
.A1(n_193),
.A2(n_152),
.B(n_156),
.C(n_137),
.Y(n_196)
);

OAI21xp5_ASAP7_75t_L g219 ( 
.A1(n_196),
.A2(n_178),
.B(n_169),
.Y(n_219)
);

A2O1A1O1Ixp25_ASAP7_75t_L g197 ( 
.A1(n_176),
.A2(n_139),
.B(n_164),
.C(n_163),
.D(n_134),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_L g221 ( 
.A(n_197),
.B(n_200),
.Y(n_221)
);

NOR2xp33_ASAP7_75t_L g217 ( 
.A(n_198),
.B(n_199),
.Y(n_217)
);

XOR2xp5_ASAP7_75t_L g200 ( 
.A(n_195),
.B(n_144),
.Y(n_200)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_190),
.Y(n_201)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_201),
.Y(n_218)
);

NOR2xp33_ASAP7_75t_L g229 ( 
.A(n_203),
.B(n_204),
.Y(n_229)
);

MAJIxp5_ASAP7_75t_L g204 ( 
.A(n_177),
.B(n_166),
.C(n_155),
.Y(n_204)
);

INVx2_ASAP7_75t_L g205 ( 
.A(n_191),
.Y(n_205)
);

NAND2xp5_ASAP7_75t_L g225 ( 
.A(n_205),
.B(n_207),
.Y(n_225)
);

AOI22xp33_ASAP7_75t_L g206 ( 
.A1(n_194),
.A2(n_193),
.B1(n_192),
.B2(n_170),
.Y(n_206)
);

CKINVDCx20_ASAP7_75t_R g220 ( 
.A(n_206),
.Y(n_220)
);

NAND2xp5_ASAP7_75t_L g209 ( 
.A(n_187),
.B(n_184),
.Y(n_209)
);

NAND2xp5_ASAP7_75t_L g227 ( 
.A(n_209),
.B(n_211),
.Y(n_227)
);

AOI22xp5_ASAP7_75t_L g223 ( 
.A1(n_210),
.A2(n_216),
.B1(n_185),
.B2(n_180),
.Y(n_223)
);

OA22x2_ASAP7_75t_L g211 ( 
.A1(n_175),
.A2(n_171),
.B1(n_179),
.B2(n_181),
.Y(n_211)
);

AOI22xp33_ASAP7_75t_L g212 ( 
.A1(n_181),
.A2(n_186),
.B1(n_182),
.B2(n_168),
.Y(n_212)
);

CKINVDCx20_ASAP7_75t_R g222 ( 
.A(n_212),
.Y(n_222)
);

OAI22xp5_ASAP7_75t_SL g228 ( 
.A1(n_213),
.A2(n_214),
.B1(n_168),
.B2(n_207),
.Y(n_228)
);

AOI22xp5_ASAP7_75t_L g214 ( 
.A1(n_183),
.A2(n_187),
.B1(n_188),
.B2(n_191),
.Y(n_214)
);

NOR2xp33_ASAP7_75t_L g215 ( 
.A(n_169),
.B(n_183),
.Y(n_215)
);

CKINVDCx20_ASAP7_75t_R g226 ( 
.A(n_215),
.Y(n_226)
);

NAND2xp5_ASAP7_75t_L g216 ( 
.A(n_172),
.B(n_182),
.Y(n_216)
);

NOR2xp33_ASAP7_75t_L g238 ( 
.A(n_219),
.B(n_226),
.Y(n_238)
);

OAI22xp5_ASAP7_75t_SL g240 ( 
.A1(n_223),
.A2(n_230),
.B1(n_220),
.B2(n_222),
.Y(n_240)
);

AOI21xp5_ASAP7_75t_L g224 ( 
.A1(n_208),
.A2(n_178),
.B(n_185),
.Y(n_224)
);

OA21x2_ASAP7_75t_L g233 ( 
.A1(n_224),
.A2(n_217),
.B(n_230),
.Y(n_233)
);

AOI22xp5_ASAP7_75t_L g232 ( 
.A1(n_228),
.A2(n_196),
.B1(n_201),
.B2(n_211),
.Y(n_232)
);

AOI22xp5_ASAP7_75t_L g230 ( 
.A1(n_211),
.A2(n_208),
.B1(n_200),
.B2(n_209),
.Y(n_230)
);

MAJIxp5_ASAP7_75t_L g231 ( 
.A(n_221),
.B(n_202),
.C(n_214),
.Y(n_231)
);

MAJIxp5_ASAP7_75t_L g246 ( 
.A(n_231),
.B(n_234),
.C(n_235),
.Y(n_246)
);

OAI22xp5_ASAP7_75t_L g243 ( 
.A1(n_232),
.A2(n_236),
.B1(n_241),
.B2(n_223),
.Y(n_243)
);

NOR2xp33_ASAP7_75t_SL g245 ( 
.A(n_233),
.B(n_238),
.Y(n_245)
);

OAI322xp33_ASAP7_75t_L g234 ( 
.A1(n_221),
.A2(n_203),
.A3(n_216),
.B1(n_198),
.B2(n_197),
.C1(n_211),
.C2(n_204),
.Y(n_234)
);

MAJIxp5_ASAP7_75t_L g235 ( 
.A(n_230),
.B(n_213),
.C(n_205),
.Y(n_235)
);

AOI22xp5_ASAP7_75t_L g236 ( 
.A1(n_228),
.A2(n_220),
.B1(n_227),
.B2(n_222),
.Y(n_236)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_225),
.Y(n_237)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_237),
.Y(n_242)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_225),
.Y(n_239)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_239),
.Y(n_247)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_240),
.Y(n_248)
);

AOI22xp5_ASAP7_75t_L g241 ( 
.A1(n_227),
.A2(n_219),
.B1(n_226),
.B2(n_223),
.Y(n_241)
);

XNOR2x1_ASAP7_75t_L g253 ( 
.A(n_243),
.B(n_240),
.Y(n_253)
);

CKINVDCx16_ASAP7_75t_R g244 ( 
.A(n_241),
.Y(n_244)
);

NOR2xp33_ASAP7_75t_SL g250 ( 
.A(n_244),
.B(n_233),
.Y(n_250)
);

OAI21xp5_ASAP7_75t_SL g249 ( 
.A1(n_246),
.A2(n_217),
.B(n_233),
.Y(n_249)
);

AOI21xp5_ASAP7_75t_L g256 ( 
.A1(n_249),
.A2(n_252),
.B(n_219),
.Y(n_256)
);

NOR2xp33_ASAP7_75t_L g255 ( 
.A(n_250),
.B(n_253),
.Y(n_255)
);

OAI22xp5_ASAP7_75t_SL g251 ( 
.A1(n_245),
.A2(n_232),
.B1(n_236),
.B2(n_235),
.Y(n_251)
);

NAND2xp5_ASAP7_75t_L g254 ( 
.A(n_251),
.B(n_248),
.Y(n_254)
);

OAI21xp5_ASAP7_75t_SL g252 ( 
.A1(n_246),
.A2(n_224),
.B(n_218),
.Y(n_252)
);

AOI22xp5_ASAP7_75t_SL g260 ( 
.A1(n_254),
.A2(n_234),
.B1(n_242),
.B2(n_247),
.Y(n_260)
);

OAI21xp5_ASAP7_75t_L g258 ( 
.A1(n_256),
.A2(n_245),
.B(n_231),
.Y(n_258)
);

NOR2xp33_ASAP7_75t_L g257 ( 
.A(n_253),
.B(n_218),
.Y(n_257)
);

MAJIxp5_ASAP7_75t_L g259 ( 
.A(n_257),
.B(n_248),
.C(n_242),
.Y(n_259)
);

NAND2xp5_ASAP7_75t_L g261 ( 
.A(n_258),
.B(n_259),
.Y(n_261)
);

MAJIxp5_ASAP7_75t_L g262 ( 
.A(n_260),
.B(n_247),
.C(n_229),
.Y(n_262)
);

OAI21xp5_ASAP7_75t_L g263 ( 
.A1(n_262),
.A2(n_229),
.B(n_255),
.Y(n_263)
);

NAND2xp5_ASAP7_75t_L g265 ( 
.A(n_263),
.B(n_264),
.Y(n_265)
);

NAND2xp5_ASAP7_75t_L g264 ( 
.A(n_261),
.B(n_237),
.Y(n_264)
);

NAND2xp5_ASAP7_75t_SL g266 ( 
.A(n_265),
.B(n_239),
.Y(n_266)
);


endmodule