module fake_jpeg_28849_n_285 (n_13, n_11, n_14, n_17, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_285);

input n_13;
input n_11;
input n_14;
input n_17;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_285;

wire n_159;
wire n_117;
wire n_253;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_251;
wire n_252;
wire n_273;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_279;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_278;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_281;
wire n_31;
wire n_155;
wire n_207;
wire n_277;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_57;
wire n_21;
wire n_223;
wire n_234;
wire n_284;
wire n_272;
wire n_280;
wire n_171;
wire n_263;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_267;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_274;
wire n_186;
wire n_44;
wire n_24;
wire n_276;
wire n_143;
wire n_202;
wire n_25;
wire n_269;
wire n_122;
wire n_75;
wire n_246;
wire n_37;
wire n_233;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_266;
wire n_34;
wire n_283;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_262;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_271;
wire n_217;
wire n_216;
wire n_264;
wire n_184;
wire n_53;
wire n_268;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_192;
wire n_156;
wire n_115;
wire n_123;
wire n_265;
wire n_176;
wire n_199;
wire n_112;
wire n_260;
wire n_270;
wire n_222;
wire n_95;
wire n_275;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_140;
wire n_82;
wire n_128;
wire n_118;
wire n_258;
wire n_282;
wire n_96;

INVx6_ASAP7_75t_SL g18 ( 
.A(n_12),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_7),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_2),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_7),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_1),
.Y(n_22)
);

INVx6_ASAP7_75t_L g23 ( 
.A(n_16),
.Y(n_23)
);

BUFx12f_ASAP7_75t_L g24 ( 
.A(n_12),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_6),
.Y(n_25)
);

INVx6_ASAP7_75t_L g26 ( 
.A(n_13),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_13),
.Y(n_27)
);

BUFx8_ASAP7_75t_L g28 ( 
.A(n_17),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_14),
.Y(n_29)
);

BUFx12f_ASAP7_75t_L g30 ( 
.A(n_0),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_1),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_8),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_8),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_17),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_8),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_16),
.Y(n_36)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_12),
.Y(n_37)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_11),
.Y(n_38)
);

BUFx12f_ASAP7_75t_L g39 ( 
.A(n_35),
.Y(n_39)
);

CKINVDCx6p67_ASAP7_75t_R g83 ( 
.A(n_39),
.Y(n_83)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_35),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_40),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_SL g41 ( 
.A(n_34),
.B(n_36),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_41),
.B(n_42),
.Y(n_71)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_28),
.Y(n_42)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_20),
.Y(n_43)
);

INVx2_ASAP7_75t_L g54 ( 
.A(n_43),
.Y(n_54)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_20),
.Y(n_44)
);

INVx2_ASAP7_75t_L g55 ( 
.A(n_44),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g45 ( 
.A(n_28),
.B(n_0),
.Y(n_45)
);

OR2x2_ASAP7_75t_L g70 ( 
.A(n_45),
.B(n_47),
.Y(n_70)
);

BUFx3_ASAP7_75t_L g46 ( 
.A(n_35),
.Y(n_46)
);

INVx4_ASAP7_75t_L g67 ( 
.A(n_46),
.Y(n_67)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_28),
.Y(n_47)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_20),
.Y(n_48)
);

INVx2_ASAP7_75t_L g68 ( 
.A(n_48),
.Y(n_68)
);

INVx2_ASAP7_75t_L g49 ( 
.A(n_35),
.Y(n_49)
);

INVx2_ASAP7_75t_L g75 ( 
.A(n_49),
.Y(n_75)
);

INVx2_ASAP7_75t_SL g50 ( 
.A(n_18),
.Y(n_50)
);

INVxp33_ASAP7_75t_L g73 ( 
.A(n_50),
.Y(n_73)
);

INVx2_ASAP7_75t_SL g51 ( 
.A(n_18),
.Y(n_51)
);

INVxp67_ASAP7_75t_L g61 ( 
.A(n_51),
.Y(n_61)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_27),
.Y(n_52)
);

INVx2_ASAP7_75t_L g84 ( 
.A(n_52),
.Y(n_84)
);

AOI22xp33_ASAP7_75t_L g53 ( 
.A1(n_45),
.A2(n_26),
.B1(n_37),
.B2(n_33),
.Y(n_53)
);

AOI22xp33_ASAP7_75t_L g99 ( 
.A1(n_53),
.A2(n_81),
.B1(n_39),
.B2(n_3),
.Y(n_99)
);

OAI22xp5_ASAP7_75t_SL g56 ( 
.A1(n_49),
.A2(n_26),
.B1(n_23),
.B2(n_30),
.Y(n_56)
);

AND2x2_ASAP7_75t_L g114 ( 
.A(n_56),
.B(n_62),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_SL g57 ( 
.A(n_41),
.B(n_34),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_SL g111 ( 
.A(n_57),
.B(n_65),
.Y(n_111)
);

AOI22xp33_ASAP7_75t_SL g58 ( 
.A1(n_42),
.A2(n_18),
.B1(n_24),
.B2(n_30),
.Y(n_58)
);

AOI22xp33_ASAP7_75t_SL g96 ( 
.A1(n_58),
.A2(n_59),
.B1(n_77),
.B2(n_85),
.Y(n_96)
);

AOI22xp33_ASAP7_75t_SL g59 ( 
.A1(n_47),
.A2(n_24),
.B1(n_30),
.B2(n_26),
.Y(n_59)
);

AOI22xp5_ASAP7_75t_SL g60 ( 
.A1(n_50),
.A2(n_21),
.B1(n_32),
.B2(n_31),
.Y(n_60)
);

AOI21xp5_ASAP7_75t_L g122 ( 
.A1(n_60),
.A2(n_82),
.B(n_4),
.Y(n_122)
);

OAI22xp5_ASAP7_75t_SL g62 ( 
.A1(n_49),
.A2(n_23),
.B1(n_30),
.B2(n_24),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_L g63 ( 
.A(n_44),
.B(n_21),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_SL g101 ( 
.A(n_63),
.B(n_2),
.Y(n_101)
);

BUFx3_ASAP7_75t_L g64 ( 
.A(n_46),
.Y(n_64)
);

INVx1_ASAP7_75t_SL g118 ( 
.A(n_64),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_SL g65 ( 
.A(n_48),
.B(n_36),
.Y(n_65)
);

OAI22xp5_ASAP7_75t_SL g66 ( 
.A1(n_40),
.A2(n_23),
.B1(n_30),
.B2(n_24),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_L g93 ( 
.A(n_66),
.B(n_80),
.Y(n_93)
);

BUFx6f_ASAP7_75t_L g72 ( 
.A(n_40),
.Y(n_72)
);

BUFx6f_ASAP7_75t_L g91 ( 
.A(n_72),
.Y(n_91)
);

INVx3_ASAP7_75t_L g74 ( 
.A(n_46),
.Y(n_74)
);

INVx3_ASAP7_75t_L g119 ( 
.A(n_74),
.Y(n_119)
);

NAND2xp67_ASAP7_75t_SL g76 ( 
.A(n_50),
.B(n_28),
.Y(n_76)
);

OR2x2_ASAP7_75t_L g105 ( 
.A(n_76),
.B(n_78),
.Y(n_105)
);

AOI22xp33_ASAP7_75t_SL g77 ( 
.A1(n_50),
.A2(n_24),
.B1(n_30),
.B2(n_33),
.Y(n_77)
);

AND2x2_ASAP7_75t_L g78 ( 
.A(n_43),
.B(n_28),
.Y(n_78)
);

OA22x2_ASAP7_75t_L g79 ( 
.A1(n_43),
.A2(n_38),
.B1(n_37),
.B2(n_33),
.Y(n_79)
);

O2A1O1Ixp33_ASAP7_75t_SL g116 ( 
.A1(n_79),
.A2(n_3),
.B(n_4),
.C(n_5),
.Y(n_116)
);

OAI22xp5_ASAP7_75t_SL g80 ( 
.A1(n_40),
.A2(n_52),
.B1(n_39),
.B2(n_31),
.Y(n_80)
);

OAI22xp33_ASAP7_75t_SL g81 ( 
.A1(n_52),
.A2(n_38),
.B1(n_37),
.B2(n_27),
.Y(n_81)
);

AOI22xp5_ASAP7_75t_L g82 ( 
.A1(n_51),
.A2(n_27),
.B1(n_38),
.B2(n_29),
.Y(n_82)
);

AOI22xp33_ASAP7_75t_SL g85 ( 
.A1(n_51),
.A2(n_32),
.B1(n_29),
.B2(n_25),
.Y(n_85)
);

BUFx6f_ASAP7_75t_L g86 ( 
.A(n_39),
.Y(n_86)
);

BUFx6f_ASAP7_75t_L g109 ( 
.A(n_86),
.Y(n_109)
);

BUFx6f_ASAP7_75t_L g87 ( 
.A(n_39),
.Y(n_87)
);

INVx6_ASAP7_75t_L g108 ( 
.A(n_87),
.Y(n_108)
);

AOI22xp33_ASAP7_75t_SL g88 ( 
.A1(n_51),
.A2(n_25),
.B1(n_22),
.B2(n_19),
.Y(n_88)
);

AOI22xp33_ASAP7_75t_SL g104 ( 
.A1(n_88),
.A2(n_39),
.B1(n_4),
.B2(n_5),
.Y(n_104)
);

BUFx12_ASAP7_75t_L g89 ( 
.A(n_83),
.Y(n_89)
);

INVxp67_ASAP7_75t_SL g126 ( 
.A(n_89),
.Y(n_126)
);

CKINVDCx14_ASAP7_75t_R g90 ( 
.A(n_76),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g130 ( 
.A(n_90),
.B(n_92),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_SL g92 ( 
.A(n_71),
.B(n_22),
.Y(n_92)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_54),
.Y(n_94)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_94),
.Y(n_139)
);

INVx8_ASAP7_75t_L g95 ( 
.A(n_67),
.Y(n_95)
);

BUFx6f_ASAP7_75t_L g132 ( 
.A(n_95),
.Y(n_132)
);

A2O1A1Ixp33_ASAP7_75t_L g97 ( 
.A1(n_70),
.A2(n_19),
.B(n_1),
.C(n_2),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_SL g133 ( 
.A(n_97),
.B(n_92),
.Y(n_133)
);

NOR2x1_ASAP7_75t_L g98 ( 
.A(n_82),
.B(n_0),
.Y(n_98)
);

OR2x2_ASAP7_75t_L g152 ( 
.A(n_98),
.B(n_99),
.Y(n_152)
);

BUFx16f_ASAP7_75t_L g100 ( 
.A(n_83),
.Y(n_100)
);

INVx6_ASAP7_75t_SL g142 ( 
.A(n_100),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_L g145 ( 
.A(n_101),
.B(n_102),
.Y(n_145)
);

INVxp67_ASAP7_75t_L g102 ( 
.A(n_78),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_SL g103 ( 
.A(n_70),
.B(n_68),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g151 ( 
.A(n_103),
.B(n_121),
.Y(n_151)
);

OAI21xp5_ASAP7_75t_SL g135 ( 
.A1(n_104),
.A2(n_120),
.B(n_122),
.Y(n_135)
);

CKINVDCx12_ASAP7_75t_R g106 ( 
.A(n_61),
.Y(n_106)
);

INVxp67_ASAP7_75t_L g124 ( 
.A(n_106),
.Y(n_124)
);

HB1xp67_ASAP7_75t_L g107 ( 
.A(n_55),
.Y(n_107)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_107),
.Y(n_147)
);

AOI22xp33_ASAP7_75t_SL g110 ( 
.A1(n_68),
.A2(n_84),
.B1(n_54),
.B2(n_74),
.Y(n_110)
);

INVxp67_ASAP7_75t_L g129 ( 
.A(n_110),
.Y(n_129)
);

XNOR2xp5_ASAP7_75t_L g112 ( 
.A(n_78),
.B(n_3),
.Y(n_112)
);

XOR2xp5_ASAP7_75t_L g137 ( 
.A(n_112),
.B(n_66),
.Y(n_137)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_84),
.Y(n_113)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_113),
.Y(n_148)
);

INVx8_ASAP7_75t_L g115 ( 
.A(n_67),
.Y(n_115)
);

INVx3_ASAP7_75t_L g143 ( 
.A(n_115),
.Y(n_143)
);

OAI22xp5_ASAP7_75t_SL g125 ( 
.A1(n_116),
.A2(n_79),
.B1(n_61),
.B2(n_69),
.Y(n_125)
);

AOI22xp33_ASAP7_75t_SL g117 ( 
.A1(n_64),
.A2(n_83),
.B1(n_79),
.B2(n_60),
.Y(n_117)
);

INVxp67_ASAP7_75t_L g131 ( 
.A(n_117),
.Y(n_131)
);

AOI22xp33_ASAP7_75t_SL g120 ( 
.A1(n_83),
.A2(n_79),
.B1(n_75),
.B2(n_69),
.Y(n_120)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_80),
.Y(n_121)
);

AND2x2_ASAP7_75t_SL g123 ( 
.A(n_121),
.B(n_75),
.Y(n_123)
);

CKINVDCx16_ASAP7_75t_R g159 ( 
.A(n_123),
.Y(n_159)
);

AOI22xp5_ASAP7_75t_SL g174 ( 
.A1(n_125),
.A2(n_95),
.B1(n_108),
.B2(n_109),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_112),
.B(n_72),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_L g156 ( 
.A(n_127),
.B(n_128),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_L g128 ( 
.A(n_122),
.B(n_56),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_SL g170 ( 
.A(n_133),
.B(n_14),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_L g134 ( 
.A(n_98),
.B(n_62),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_L g165 ( 
.A(n_134),
.B(n_136),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_L g136 ( 
.A(n_105),
.B(n_87),
.Y(n_136)
);

XOR2xp5_ASAP7_75t_L g153 ( 
.A(n_137),
.B(n_114),
.Y(n_153)
);

AOI22xp33_ASAP7_75t_L g138 ( 
.A1(n_114),
.A2(n_73),
.B1(n_86),
.B2(n_7),
.Y(n_138)
);

OAI22xp5_ASAP7_75t_SL g168 ( 
.A1(n_138),
.A2(n_146),
.B1(n_91),
.B2(n_97),
.Y(n_168)
);

OAI22xp5_ASAP7_75t_SL g140 ( 
.A1(n_93),
.A2(n_73),
.B1(n_6),
.B2(n_9),
.Y(n_140)
);

AOI22xp5_ASAP7_75t_L g167 ( 
.A1(n_140),
.A2(n_149),
.B1(n_11),
.B2(n_13),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_L g141 ( 
.A(n_105),
.B(n_5),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_L g178 ( 
.A(n_141),
.B(n_14),
.Y(n_178)
);

INVx2_ASAP7_75t_SL g144 ( 
.A(n_100),
.Y(n_144)
);

NOR2xp33_ASAP7_75t_L g160 ( 
.A(n_144),
.B(n_150),
.Y(n_160)
);

AOI22xp33_ASAP7_75t_L g146 ( 
.A1(n_114),
.A2(n_6),
.B1(n_9),
.B2(n_10),
.Y(n_146)
);

OAI22xp5_ASAP7_75t_SL g149 ( 
.A1(n_93),
.A2(n_9),
.B1(n_10),
.B2(n_11),
.Y(n_149)
);

NOR2xp33_ASAP7_75t_L g150 ( 
.A(n_111),
.B(n_10),
.Y(n_150)
);

XOR2xp5_ASAP7_75t_L g198 ( 
.A(n_153),
.B(n_169),
.Y(n_198)
);

NOR2xp33_ASAP7_75t_L g154 ( 
.A(n_130),
.B(n_151),
.Y(n_154)
);

NOR2xp33_ASAP7_75t_L g196 ( 
.A(n_154),
.B(n_162),
.Y(n_196)
);

NOR2x1_ASAP7_75t_L g155 ( 
.A(n_125),
.B(n_116),
.Y(n_155)
);

OAI21xp5_ASAP7_75t_L g192 ( 
.A1(n_155),
.A2(n_152),
.B(n_133),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_SL g157 ( 
.A(n_151),
.B(n_102),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_L g184 ( 
.A(n_157),
.B(n_166),
.Y(n_184)
);

AOI21xp5_ASAP7_75t_L g158 ( 
.A1(n_131),
.A2(n_96),
.B(n_118),
.Y(n_158)
);

AOI21xp5_ASAP7_75t_L g197 ( 
.A1(n_158),
.A2(n_163),
.B(n_144),
.Y(n_197)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_139),
.Y(n_161)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_161),
.Y(n_185)
);

INVxp67_ASAP7_75t_L g162 ( 
.A(n_136),
.Y(n_162)
);

AOI21xp5_ASAP7_75t_L g163 ( 
.A1(n_135),
.A2(n_118),
.B(n_100),
.Y(n_163)
);

CKINVDCx20_ASAP7_75t_R g164 ( 
.A(n_123),
.Y(n_164)
);

CKINVDCx20_ASAP7_75t_R g183 ( 
.A(n_164),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_SL g166 ( 
.A(n_137),
.B(n_113),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_L g205 ( 
.A(n_167),
.B(n_173),
.Y(n_205)
);

AOI22xp5_ASAP7_75t_L g188 ( 
.A1(n_168),
.A2(n_182),
.B1(n_140),
.B2(n_149),
.Y(n_188)
);

MAJx2_ASAP7_75t_L g169 ( 
.A(n_127),
.B(n_94),
.C(n_89),
.Y(n_169)
);

NOR2xp33_ASAP7_75t_SL g202 ( 
.A(n_170),
.B(n_145),
.Y(n_202)
);

NOR2xp33_ASAP7_75t_L g171 ( 
.A(n_130),
.B(n_89),
.Y(n_171)
);

NOR2xp33_ASAP7_75t_L g191 ( 
.A(n_171),
.B(n_177),
.Y(n_191)
);

AOI22xp5_ASAP7_75t_L g172 ( 
.A1(n_123),
.A2(n_119),
.B1(n_91),
.B2(n_115),
.Y(n_172)
);

OAI22xp5_ASAP7_75t_SL g194 ( 
.A1(n_172),
.A2(n_174),
.B1(n_144),
.B2(n_143),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_SL g173 ( 
.A(n_123),
.B(n_119),
.Y(n_173)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_139),
.Y(n_175)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_175),
.Y(n_190)
);

CKINVDCx20_ASAP7_75t_R g176 ( 
.A(n_126),
.Y(n_176)
);

CKINVDCx20_ASAP7_75t_R g200 ( 
.A(n_176),
.Y(n_200)
);

INVxp67_ASAP7_75t_L g177 ( 
.A(n_143),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_L g206 ( 
.A(n_178),
.B(n_15),
.Y(n_206)
);

HAxp5_ASAP7_75t_SL g179 ( 
.A(n_141),
.B(n_15),
.CON(n_179),
.SN(n_179)
);

INVxp67_ASAP7_75t_L g186 ( 
.A(n_179),
.Y(n_186)
);

AND2x2_ASAP7_75t_L g180 ( 
.A(n_134),
.B(n_108),
.Y(n_180)
);

INVx1_ASAP7_75t_SL g199 ( 
.A(n_180),
.Y(n_199)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_148),
.Y(n_181)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_181),
.Y(n_195)
);

OAI22xp5_ASAP7_75t_L g182 ( 
.A1(n_128),
.A2(n_15),
.B1(n_109),
.B2(n_152),
.Y(n_182)
);

CKINVDCx16_ASAP7_75t_R g187 ( 
.A(n_180),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_SL g219 ( 
.A(n_187),
.B(n_193),
.Y(n_219)
);

OAI22xp5_ASAP7_75t_SL g207 ( 
.A1(n_188),
.A2(n_189),
.B1(n_201),
.B2(n_203),
.Y(n_207)
);

AOI22xp5_ASAP7_75t_L g189 ( 
.A1(n_182),
.A2(n_129),
.B1(n_135),
.B2(n_152),
.Y(n_189)
);

AOI21xp5_ASAP7_75t_L g221 ( 
.A1(n_192),
.A2(n_197),
.B(n_173),
.Y(n_221)
);

CKINVDCx16_ASAP7_75t_R g193 ( 
.A(n_180),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_L g216 ( 
.A(n_194),
.B(n_206),
.Y(n_216)
);

OAI22xp5_ASAP7_75t_L g201 ( 
.A1(n_174),
.A2(n_145),
.B1(n_148),
.B2(n_147),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_SL g223 ( 
.A(n_202),
.B(n_170),
.Y(n_223)
);

OAI22xp5_ASAP7_75t_L g203 ( 
.A1(n_165),
.A2(n_147),
.B1(n_132),
.B2(n_142),
.Y(n_203)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_161),
.Y(n_204)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_204),
.Y(n_215)
);

INVx1_ASAP7_75t_SL g208 ( 
.A(n_203),
.Y(n_208)
);

NAND2xp5_ASAP7_75t_L g237 ( 
.A(n_208),
.B(n_223),
.Y(n_237)
);

OAI21xp5_ASAP7_75t_L g209 ( 
.A1(n_197),
.A2(n_163),
.B(n_158),
.Y(n_209)
);

OAI21xp5_ASAP7_75t_L g230 ( 
.A1(n_209),
.A2(n_214),
.B(n_221),
.Y(n_230)
);

MAJIxp5_ASAP7_75t_L g210 ( 
.A(n_198),
.B(n_153),
.C(n_166),
.Y(n_210)
);

MAJIxp5_ASAP7_75t_L g228 ( 
.A(n_210),
.B(n_224),
.C(n_157),
.Y(n_228)
);

CKINVDCx20_ASAP7_75t_R g211 ( 
.A(n_196),
.Y(n_211)
);

CKINVDCx20_ASAP7_75t_R g232 ( 
.A(n_211),
.Y(n_232)
);

CKINVDCx16_ASAP7_75t_R g212 ( 
.A(n_185),
.Y(n_212)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_212),
.Y(n_241)
);

NOR2xp33_ASAP7_75t_L g213 ( 
.A(n_202),
.B(n_160),
.Y(n_213)
);

OAI21xp33_ASAP7_75t_L g239 ( 
.A1(n_213),
.A2(n_226),
.B(n_178),
.Y(n_239)
);

OAI21xp5_ASAP7_75t_L g214 ( 
.A1(n_192),
.A2(n_165),
.B(n_156),
.Y(n_214)
);

XNOR2x1_ASAP7_75t_L g217 ( 
.A(n_198),
.B(n_156),
.Y(n_217)
);

XNOR2xp5_ASAP7_75t_L g238 ( 
.A(n_217),
.B(n_220),
.Y(n_238)
);

OAI22xp5_ASAP7_75t_SL g218 ( 
.A1(n_189),
.A2(n_159),
.B1(n_155),
.B2(n_164),
.Y(n_218)
);

AOI22xp5_ASAP7_75t_L g227 ( 
.A1(n_218),
.A2(n_222),
.B1(n_187),
.B2(n_193),
.Y(n_227)
);

XNOR2xp5_ASAP7_75t_L g220 ( 
.A(n_184),
.B(n_169),
.Y(n_220)
);

OAI22xp5_ASAP7_75t_SL g222 ( 
.A1(n_188),
.A2(n_159),
.B1(n_155),
.B2(n_172),
.Y(n_222)
);

XNOR2xp5_ASAP7_75t_L g224 ( 
.A(n_184),
.B(n_169),
.Y(n_224)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_185),
.Y(n_225)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_225),
.Y(n_233)
);

NOR2xp33_ASAP7_75t_L g226 ( 
.A(n_196),
.B(n_160),
.Y(n_226)
);

NAND2xp5_ASAP7_75t_L g245 ( 
.A(n_227),
.B(n_231),
.Y(n_245)
);

XNOR2xp5_ASAP7_75t_L g247 ( 
.A(n_228),
.B(n_229),
.Y(n_247)
);

MAJIxp5_ASAP7_75t_L g229 ( 
.A(n_210),
.B(n_183),
.C(n_199),
.Y(n_229)
);

OAI22xp5_ASAP7_75t_SL g231 ( 
.A1(n_208),
.A2(n_199),
.B1(n_205),
.B2(n_183),
.Y(n_231)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_215),
.Y(n_234)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_234),
.Y(n_243)
);

AOI22xp5_ASAP7_75t_SL g235 ( 
.A1(n_207),
.A2(n_201),
.B1(n_194),
.B2(n_168),
.Y(n_235)
);

INVxp67_ASAP7_75t_L g244 ( 
.A(n_235),
.Y(n_244)
);

OAI21xp5_ASAP7_75t_SL g236 ( 
.A1(n_221),
.A2(n_205),
.B(n_191),
.Y(n_236)
);

AOI21xp5_ASAP7_75t_L g242 ( 
.A1(n_236),
.A2(n_209),
.B(n_218),
.Y(n_242)
);

INVx13_ASAP7_75t_L g252 ( 
.A(n_239),
.Y(n_252)
);

OAI22xp5_ASAP7_75t_SL g240 ( 
.A1(n_216),
.A2(n_204),
.B1(n_190),
.B2(n_195),
.Y(n_240)
);

NAND2xp5_ASAP7_75t_L g250 ( 
.A(n_240),
.B(n_225),
.Y(n_250)
);

XNOR2xp5_ASAP7_75t_L g262 ( 
.A(n_242),
.B(n_246),
.Y(n_262)
);

OAI21xp5_ASAP7_75t_SL g246 ( 
.A1(n_237),
.A2(n_219),
.B(n_186),
.Y(n_246)
);

XNOR2xp5_ASAP7_75t_L g248 ( 
.A(n_228),
.B(n_217),
.Y(n_248)
);

MAJIxp5_ASAP7_75t_L g256 ( 
.A(n_248),
.B(n_249),
.C(n_247),
.Y(n_256)
);

MAJx2_ASAP7_75t_L g249 ( 
.A(n_229),
.B(n_224),
.C(n_220),
.Y(n_249)
);

MAJIxp5_ASAP7_75t_L g255 ( 
.A(n_249),
.B(n_238),
.C(n_211),
.Y(n_255)
);

NAND2xp5_ASAP7_75t_L g259 ( 
.A(n_250),
.B(n_251),
.Y(n_259)
);

OAI21xp5_ASAP7_75t_L g251 ( 
.A1(n_230),
.A2(n_227),
.B(n_237),
.Y(n_251)
);

OAI21xp5_ASAP7_75t_L g253 ( 
.A1(n_230),
.A2(n_214),
.B(n_216),
.Y(n_253)
);

NOR2xp33_ASAP7_75t_L g263 ( 
.A(n_253),
.B(n_254),
.Y(n_263)
);

BUFx2_ASAP7_75t_L g254 ( 
.A(n_241),
.Y(n_254)
);

NAND2xp5_ASAP7_75t_SL g266 ( 
.A(n_255),
.B(n_256),
.Y(n_266)
);

NOR2xp33_ASAP7_75t_SL g257 ( 
.A(n_247),
.B(n_232),
.Y(n_257)
);

NOR2xp33_ASAP7_75t_L g270 ( 
.A(n_257),
.B(n_258),
.Y(n_270)
);

MAJIxp5_ASAP7_75t_L g258 ( 
.A(n_248),
.B(n_238),
.C(n_236),
.Y(n_258)
);

MAJIxp5_ASAP7_75t_L g260 ( 
.A(n_251),
.B(n_242),
.C(n_253),
.Y(n_260)
);

NOR2xp33_ASAP7_75t_SL g264 ( 
.A(n_260),
.B(n_261),
.Y(n_264)
);

OAI22xp5_ASAP7_75t_L g261 ( 
.A1(n_244),
.A2(n_235),
.B1(n_234),
.B2(n_233),
.Y(n_261)
);

OAI22xp5_ASAP7_75t_SL g265 ( 
.A1(n_263),
.A2(n_244),
.B1(n_245),
.B2(n_207),
.Y(n_265)
);

AOI22xp5_ASAP7_75t_L g271 ( 
.A1(n_265),
.A2(n_222),
.B1(n_240),
.B2(n_259),
.Y(n_271)
);

NOR2xp33_ASAP7_75t_SL g267 ( 
.A(n_262),
.B(n_206),
.Y(n_267)
);

CKINVDCx14_ASAP7_75t_R g273 ( 
.A(n_267),
.Y(n_273)
);

OAI21xp5_ASAP7_75t_SL g268 ( 
.A1(n_263),
.A2(n_231),
.B(n_243),
.Y(n_268)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_268),
.Y(n_272)
);

NOR2xp67_ASAP7_75t_L g269 ( 
.A(n_256),
.B(n_252),
.Y(n_269)
);

NOR2xp33_ASAP7_75t_SL g275 ( 
.A(n_269),
.B(n_200),
.Y(n_275)
);

OAI22xp5_ASAP7_75t_SL g279 ( 
.A1(n_271),
.A2(n_265),
.B1(n_268),
.B2(n_200),
.Y(n_279)
);

OAI22xp5_ASAP7_75t_SL g274 ( 
.A1(n_264),
.A2(n_233),
.B1(n_252),
.B2(n_215),
.Y(n_274)
);

NAND2xp5_ASAP7_75t_L g276 ( 
.A(n_274),
.B(n_275),
.Y(n_276)
);

NAND2xp5_ASAP7_75t_L g277 ( 
.A(n_274),
.B(n_254),
.Y(n_277)
);

OAI22xp5_ASAP7_75t_L g281 ( 
.A1(n_277),
.A2(n_278),
.B1(n_175),
.B2(n_176),
.Y(n_281)
);

NAND2xp5_ASAP7_75t_L g278 ( 
.A(n_273),
.B(n_270),
.Y(n_278)
);

AOI322xp5_ASAP7_75t_L g280 ( 
.A1(n_279),
.A2(n_272),
.A3(n_271),
.B1(n_195),
.B2(n_190),
.C1(n_266),
.C2(n_181),
.Y(n_280)
);

AOI322xp5_ASAP7_75t_L g282 ( 
.A1(n_280),
.A2(n_281),
.A3(n_276),
.B1(n_279),
.B2(n_132),
.C1(n_124),
.C2(n_142),
.Y(n_282)
);

MAJIxp5_ASAP7_75t_L g283 ( 
.A(n_282),
.B(n_132),
.C(n_167),
.Y(n_283)
);

INVxp67_ASAP7_75t_L g284 ( 
.A(n_283),
.Y(n_284)
);

BUFx24_ASAP7_75t_SL g285 ( 
.A(n_284),
.Y(n_285)
);


endmodule