module fake_netlist_6_551_n_1750 (n_52, n_16, n_1, n_91, n_119, n_46, n_146, n_18, n_21, n_147, n_154, n_88, n_3, n_98, n_113, n_39, n_63, n_73, n_4, n_148, n_138, n_22, n_68, n_28, n_50, n_49, n_7, n_83, n_5, n_101, n_144, n_127, n_125, n_153, n_77, n_149, n_152, n_106, n_92, n_145, n_42, n_133, n_96, n_8, n_90, n_24, n_105, n_131, n_54, n_132, n_102, n_0, n_87, n_32, n_66, n_85, n_99, n_78, n_84, n_130, n_100, n_129, n_13, n_121, n_11, n_137, n_17, n_23, n_142, n_20, n_143, n_2, n_19, n_47, n_62, n_29, n_75, n_109, n_150, n_122, n_45, n_34, n_140, n_70, n_120, n_37, n_15, n_67, n_33, n_82, n_27, n_38, n_110, n_151, n_61, n_112, n_81, n_59, n_76, n_36, n_26, n_124, n_55, n_126, n_94, n_97, n_108, n_58, n_116, n_64, n_117, n_118, n_48, n_65, n_25, n_40, n_93, n_80, n_141, n_135, n_139, n_41, n_134, n_114, n_86, n_104, n_95, n_9, n_107, n_10, n_71, n_74, n_6, n_14, n_123, n_136, n_72, n_89, n_103, n_111, n_60, n_35, n_115, n_12, n_69, n_128, n_30, n_79, n_43, n_31, n_57, n_53, n_51, n_44, n_56, n_1750);

input n_52;
input n_16;
input n_1;
input n_91;
input n_119;
input n_46;
input n_146;
input n_18;
input n_21;
input n_147;
input n_154;
input n_88;
input n_3;
input n_98;
input n_113;
input n_39;
input n_63;
input n_73;
input n_4;
input n_148;
input n_138;
input n_22;
input n_68;
input n_28;
input n_50;
input n_49;
input n_7;
input n_83;
input n_5;
input n_101;
input n_144;
input n_127;
input n_125;
input n_153;
input n_77;
input n_149;
input n_152;
input n_106;
input n_92;
input n_145;
input n_42;
input n_133;
input n_96;
input n_8;
input n_90;
input n_24;
input n_105;
input n_131;
input n_54;
input n_132;
input n_102;
input n_0;
input n_87;
input n_32;
input n_66;
input n_85;
input n_99;
input n_78;
input n_84;
input n_130;
input n_100;
input n_129;
input n_13;
input n_121;
input n_11;
input n_137;
input n_17;
input n_23;
input n_142;
input n_20;
input n_143;
input n_2;
input n_19;
input n_47;
input n_62;
input n_29;
input n_75;
input n_109;
input n_150;
input n_122;
input n_45;
input n_34;
input n_140;
input n_70;
input n_120;
input n_37;
input n_15;
input n_67;
input n_33;
input n_82;
input n_27;
input n_38;
input n_110;
input n_151;
input n_61;
input n_112;
input n_81;
input n_59;
input n_76;
input n_36;
input n_26;
input n_124;
input n_55;
input n_126;
input n_94;
input n_97;
input n_108;
input n_58;
input n_116;
input n_64;
input n_117;
input n_118;
input n_48;
input n_65;
input n_25;
input n_40;
input n_93;
input n_80;
input n_141;
input n_135;
input n_139;
input n_41;
input n_134;
input n_114;
input n_86;
input n_104;
input n_95;
input n_9;
input n_107;
input n_10;
input n_71;
input n_74;
input n_6;
input n_14;
input n_123;
input n_136;
input n_72;
input n_89;
input n_103;
input n_111;
input n_60;
input n_35;
input n_115;
input n_12;
input n_69;
input n_128;
input n_30;
input n_79;
input n_43;
input n_31;
input n_57;
input n_53;
input n_51;
input n_44;
input n_56;

output n_1750;

wire n_992;
wire n_1671;
wire n_801;
wire n_1613;
wire n_1234;
wire n_1458;
wire n_1199;
wire n_1674;
wire n_741;
wire n_1027;
wire n_1351;
wire n_625;
wire n_1189;
wire n_223;
wire n_1212;
wire n_226;
wire n_208;
wire n_726;
wire n_212;
wire n_700;
wire n_1307;
wire n_1038;
wire n_578;
wire n_1581;
wire n_1003;
wire n_365;
wire n_168;
wire n_1237;
wire n_1061;
wire n_1357;
wire n_783;
wire n_1738;
wire n_798;
wire n_188;
wire n_1575;
wire n_509;
wire n_1342;
wire n_245;
wire n_1209;
wire n_1348;
wire n_1387;
wire n_677;
wire n_1708;
wire n_805;
wire n_1151;
wire n_396;
wire n_1739;
wire n_350;
wire n_1380;
wire n_442;
wire n_480;
wire n_1402;
wire n_1688;
wire n_1691;
wire n_1009;
wire n_1743;
wire n_1160;
wire n_883;
wire n_1238;
wire n_1724;
wire n_1032;
wire n_1247;
wire n_1547;
wire n_1553;
wire n_893;
wire n_1099;
wire n_1264;
wire n_1192;
wire n_471;
wire n_424;
wire n_1700;
wire n_1555;
wire n_1415;
wire n_1370;
wire n_369;
wire n_287;
wire n_415;
wire n_830;
wire n_230;
wire n_461;
wire n_873;
wire n_383;
wire n_1285;
wire n_1371;
wire n_200;
wire n_447;
wire n_1172;
wire n_852;
wire n_229;
wire n_1590;
wire n_1532;
wire n_1393;
wire n_1517;
wire n_1704;
wire n_1078;
wire n_250;
wire n_544;
wire n_1711;
wire n_1140;
wire n_1444;
wire n_1670;
wire n_1603;
wire n_1579;
wire n_1263;
wire n_836;
wire n_375;
wire n_522;
wire n_1261;
wire n_945;
wire n_1649;
wire n_1511;
wire n_1143;
wire n_1422;
wire n_1232;
wire n_1572;
wire n_616;
wire n_658;
wire n_1119;
wire n_428;
wire n_1433;
wire n_1620;
wire n_1735;
wire n_1541;
wire n_1300;
wire n_641;
wire n_822;
wire n_693;
wire n_1313;
wire n_1056;
wire n_758;
wire n_516;
wire n_1455;
wire n_1163;
wire n_1180;
wire n_943;
wire n_1550;
wire n_491;
wire n_1591;
wire n_772;
wire n_1344;
wire n_666;
wire n_371;
wire n_940;
wire n_770;
wire n_567;
wire n_405;
wire n_213;
wire n_538;
wire n_1106;
wire n_886;
wire n_1471;
wire n_343;
wire n_953;
wire n_1094;
wire n_1345;
wire n_494;
wire n_539;
wire n_493;
wire n_155;
wire n_454;
wire n_1421;
wire n_638;
wire n_1404;
wire n_1211;
wire n_381;
wire n_887;
wire n_1660;
wire n_1280;
wire n_713;
wire n_1400;
wire n_1467;
wire n_976;
wire n_224;
wire n_1445;
wire n_1526;
wire n_1560;
wire n_734;
wire n_1088;
wire n_196;
wire n_1231;
wire n_917;
wire n_574;
wire n_907;
wire n_1446;
wire n_659;
wire n_407;
wire n_913;
wire n_1658;
wire n_808;
wire n_867;
wire n_1230;
wire n_473;
wire n_1193;
wire n_1054;
wire n_559;
wire n_1333;
wire n_1648;
wire n_163;
wire n_1644;
wire n_1558;
wire n_1732;
wire n_281;
wire n_551;
wire n_699;
wire n_564;
wire n_451;
wire n_824;
wire n_279;
wire n_686;
wire n_757;
wire n_594;
wire n_1641;
wire n_577;
wire n_166;
wire n_619;
wire n_1367;
wire n_1336;
wire n_521;
wire n_572;
wire n_395;
wire n_813;
wire n_1481;
wire n_323;
wire n_606;
wire n_1441;
wire n_818;
wire n_1123;
wire n_1309;
wire n_513;
wire n_645;
wire n_1381;
wire n_331;
wire n_1699;
wire n_916;
wire n_483;
wire n_608;
wire n_261;
wire n_630;
wire n_541;
wire n_512;
wire n_433;
wire n_792;
wire n_476;
wire n_1328;
wire n_219;
wire n_264;
wire n_263;
wire n_1162;
wire n_860;
wire n_1530;
wire n_788;
wire n_939;
wire n_1543;
wire n_821;
wire n_938;
wire n_1302;
wire n_1068;
wire n_1599;
wire n_329;
wire n_982;
wire n_549;
wire n_1075;
wire n_408;
wire n_932;
wire n_237;
wire n_1697;
wire n_243;
wire n_979;
wire n_905;
wire n_1680;
wire n_175;
wire n_322;
wire n_993;
wire n_689;
wire n_354;
wire n_1330;
wire n_1413;
wire n_1605;
wire n_1278;
wire n_547;
wire n_558;
wire n_1064;
wire n_1396;
wire n_634;
wire n_966;
wire n_764;
wire n_1663;
wire n_692;
wire n_733;
wire n_1233;
wire n_1289;
wire n_487;
wire n_241;
wire n_1107;
wire n_1014;
wire n_1290;
wire n_1703;
wire n_882;
wire n_1354;
wire n_586;
wire n_423;
wire n_1701;
wire n_318;
wire n_1111;
wire n_1713;
wire n_715;
wire n_1251;
wire n_1265;
wire n_1726;
wire n_530;
wire n_1563;
wire n_277;
wire n_618;
wire n_1297;
wire n_1662;
wire n_1312;
wire n_199;
wire n_1167;
wire n_1359;
wire n_674;
wire n_871;
wire n_922;
wire n_268;
wire n_1335;
wire n_210;
wire n_1069;
wire n_1664;
wire n_1722;
wire n_612;
wire n_178;
wire n_247;
wire n_1165;
wire n_355;
wire n_702;
wire n_347;
wire n_1175;
wire n_328;
wire n_1386;
wire n_429;
wire n_1747;
wire n_1012;
wire n_195;
wire n_780;
wire n_675;
wire n_903;
wire n_1540;
wire n_1504;
wire n_286;
wire n_254;
wire n_1655;
wire n_242;
wire n_928;
wire n_835;
wire n_1214;
wire n_690;
wire n_850;
wire n_1654;
wire n_816;
wire n_1157;
wire n_1462;
wire n_1188;
wire n_877;
wire n_604;
wire n_825;
wire n_728;
wire n_1063;
wire n_1588;
wire n_267;
wire n_1124;
wire n_1624;
wire n_515;
wire n_598;
wire n_696;
wire n_1515;
wire n_961;
wire n_437;
wire n_1082;
wire n_1317;
wire n_593;
wire n_514;
wire n_687;
wire n_697;
wire n_890;
wire n_637;
wire n_295;
wire n_701;
wire n_950;
wire n_388;
wire n_190;
wire n_484;
wire n_1709;
wire n_170;
wire n_891;
wire n_1412;
wire n_949;
wire n_1630;
wire n_678;
wire n_283;
wire n_507;
wire n_968;
wire n_909;
wire n_1369;
wire n_881;
wire n_1008;
wire n_760;
wire n_1546;
wire n_590;
wire n_362;
wire n_161;
wire n_462;
wire n_1052;
wire n_1033;
wire n_1296;
wire n_304;
wire n_694;
wire n_1294;
wire n_1420;
wire n_1634;
wire n_595;
wire n_627;
wire n_297;
wire n_524;
wire n_1465;
wire n_342;
wire n_1044;
wire n_1712;
wire n_1391;
wire n_449;
wire n_1523;
wire n_1208;
wire n_1164;
wire n_1295;
wire n_1627;
wire n_1072;
wire n_1527;
wire n_1495;
wire n_1438;
wire n_495;
wire n_815;
wire n_1100;
wire n_585;
wire n_1487;
wire n_840;
wire n_874;
wire n_1128;
wire n_382;
wire n_673;
wire n_1071;
wire n_1067;
wire n_1565;
wire n_1493;
wire n_898;
wire n_255;
wire n_284;
wire n_865;
wire n_925;
wire n_1101;
wire n_1026;
wire n_289;
wire n_1364;
wire n_615;
wire n_1249;
wire n_1293;
wire n_1127;
wire n_1512;
wire n_1451;
wire n_320;
wire n_639;
wire n_963;
wire n_794;
wire n_727;
wire n_894;
wire n_685;
wire n_353;
wire n_605;
wire n_1514;
wire n_826;
wire n_1646;
wire n_872;
wire n_1139;
wire n_1714;
wire n_718;
wire n_1018;
wire n_1521;
wire n_1366;
wire n_542;
wire n_847;
wire n_644;
wire n_682;
wire n_851;
wire n_305;
wire n_996;
wire n_532;
wire n_173;
wire n_1308;
wire n_1376;
wire n_1513;
wire n_413;
wire n_791;
wire n_510;
wire n_837;
wire n_1488;
wire n_948;
wire n_704;
wire n_977;
wire n_1005;
wire n_536;
wire n_622;
wire n_1469;
wire n_581;
wire n_765;
wire n_432;
wire n_987;
wire n_1492;
wire n_1340;
wire n_631;
wire n_720;
wire n_842;
wire n_1707;
wire n_1432;
wire n_156;
wire n_843;
wire n_656;
wire n_989;
wire n_1277;
wire n_797;
wire n_1473;
wire n_1723;
wire n_1246;
wire n_899;
wire n_189;
wire n_738;
wire n_1304;
wire n_1035;
wire n_294;
wire n_499;
wire n_1426;
wire n_705;
wire n_1004;
wire n_1176;
wire n_1529;
wire n_1022;
wire n_614;
wire n_529;
wire n_425;
wire n_684;
wire n_1431;
wire n_1615;
wire n_1474;
wire n_1571;
wire n_1577;
wire n_1181;
wire n_486;
wire n_947;
wire n_1117;
wire n_1087;
wire n_1448;
wire n_648;
wire n_657;
wire n_1049;
wire n_1666;
wire n_1505;
wire n_803;
wire n_290;
wire n_1717;
wire n_926;
wire n_927;
wire n_919;
wire n_1698;
wire n_478;
wire n_929;
wire n_1228;
wire n_417;
wire n_446;
wire n_1568;
wire n_1490;
wire n_777;
wire n_1299;
wire n_272;
wire n_526;
wire n_1183;
wire n_1436;
wire n_1384;
wire n_293;
wire n_458;
wire n_1070;
wire n_998;
wire n_717;
wire n_1665;
wire n_1383;
wire n_1178;
wire n_1424;
wire n_1073;
wire n_1000;
wire n_796;
wire n_252;
wire n_1195;
wire n_1626;
wire n_1507;
wire n_184;
wire n_552;
wire n_1358;
wire n_1388;
wire n_216;
wire n_912;
wire n_1519;
wire n_745;
wire n_1284;
wire n_1604;
wire n_1142;
wire n_716;
wire n_1475;
wire n_623;
wire n_1048;
wire n_1201;
wire n_1398;
wire n_884;
wire n_1395;
wire n_731;
wire n_1502;
wire n_1659;
wire n_755;
wire n_931;
wire n_1021;
wire n_474;
wire n_527;
wire n_683;
wire n_811;
wire n_1207;
wire n_312;
wire n_1368;
wire n_1418;
wire n_958;
wire n_292;
wire n_1250;
wire n_1137;
wire n_880;
wire n_889;
wire n_1478;
wire n_589;
wire n_1310;
wire n_819;
wire n_1363;
wire n_1334;
wire n_767;
wire n_1314;
wire n_600;
wire n_964;
wire n_831;
wire n_477;
wire n_954;
wire n_864;
wire n_1110;
wire n_1410;
wire n_399;
wire n_1440;
wire n_1382;
wire n_1534;
wire n_1564;
wire n_1736;
wire n_211;
wire n_1483;
wire n_1372;
wire n_231;
wire n_1457;
wire n_505;
wire n_1719;
wire n_319;
wire n_1339;
wire n_537;
wire n_1427;
wire n_311;
wire n_1466;
wire n_403;
wire n_1080;
wire n_723;
wire n_596;
wire n_546;
wire n_562;
wire n_1141;
wire n_1268;
wire n_386;
wire n_1220;
wire n_556;
wire n_162;
wire n_1602;
wire n_1136;
wire n_1125;
wire n_970;
wire n_642;
wire n_995;
wire n_276;
wire n_1159;
wire n_1092;
wire n_441;
wire n_221;
wire n_1060;
wire n_444;
wire n_1252;
wire n_1223;
wire n_303;
wire n_511;
wire n_193;
wire n_1286;
wire n_1053;
wire n_416;
wire n_1681;
wire n_520;
wire n_418;
wire n_1093;
wire n_1533;
wire n_1597;
wire n_266;
wire n_296;
wire n_775;
wire n_651;
wire n_1153;
wire n_439;
wire n_1618;
wire n_217;
wire n_518;
wire n_1531;
wire n_1185;
wire n_453;
wire n_215;
wire n_1745;
wire n_914;
wire n_759;
wire n_426;
wire n_317;
wire n_1653;
wire n_1679;
wire n_1625;
wire n_1453;
wire n_488;
wire n_497;
wire n_773;
wire n_920;
wire n_1374;
wire n_1315;
wire n_1647;
wire n_1224;
wire n_1614;
wire n_1459;
wire n_1135;
wire n_1169;
wire n_1179;
wire n_401;
wire n_324;
wire n_1617;
wire n_335;
wire n_1470;
wire n_463;
wire n_1243;
wire n_848;
wire n_301;
wire n_274;
wire n_1096;
wire n_1091;
wire n_1580;
wire n_1425;
wire n_1281;
wire n_1267;
wire n_983;
wire n_427;
wire n_1520;
wire n_496;
wire n_906;
wire n_1390;
wire n_688;
wire n_1077;
wire n_1733;
wire n_1419;
wire n_351;
wire n_259;
wire n_1731;
wire n_177;
wire n_1636;
wire n_1437;
wire n_1645;
wire n_385;
wire n_1687;
wire n_1439;
wire n_1323;
wire n_858;
wire n_1331;
wire n_613;
wire n_736;
wire n_501;
wire n_956;
wire n_960;
wire n_663;
wire n_856;
wire n_379;
wire n_778;
wire n_1668;
wire n_1134;
wire n_410;
wire n_1129;
wire n_554;
wire n_602;
wire n_1696;
wire n_1594;
wire n_664;
wire n_171;
wire n_169;
wire n_1429;
wire n_1610;
wire n_435;
wire n_793;
wire n_326;
wire n_587;
wire n_1593;
wire n_580;
wire n_762;
wire n_1030;
wire n_1202;
wire n_465;
wire n_1635;
wire n_1079;
wire n_341;
wire n_1744;
wire n_828;
wire n_607;
wire n_316;
wire n_419;
wire n_1551;
wire n_1103;
wire n_1203;
wire n_820;
wire n_951;
wire n_725;
wire n_952;
wire n_999;
wire n_358;
wire n_1254;
wire n_160;
wire n_186;
wire n_368;
wire n_575;
wire n_994;
wire n_1508;
wire n_732;
wire n_974;
wire n_392;
wire n_724;
wire n_1020;
wire n_1042;
wire n_628;
wire n_1273;
wire n_1434;
wire n_1573;
wire n_1728;
wire n_557;
wire n_349;
wire n_617;
wire n_845;
wire n_807;
wire n_1036;
wire n_1138;
wire n_1661;
wire n_1275;
wire n_485;
wire n_1549;
wire n_443;
wire n_1510;
wire n_892;
wire n_768;
wire n_421;
wire n_1468;
wire n_238;
wire n_1095;
wire n_1595;
wire n_202;
wire n_1718;
wire n_1749;
wire n_1683;
wire n_597;
wire n_280;
wire n_1270;
wire n_1187;
wire n_610;
wire n_1403;
wire n_1669;
wire n_1024;
wire n_198;
wire n_179;
wire n_248;
wire n_517;
wire n_1667;
wire n_667;
wire n_1206;
wire n_621;
wire n_1037;
wire n_1397;
wire n_1279;
wire n_1115;
wire n_750;
wire n_901;
wire n_1499;
wire n_468;
wire n_923;
wire n_504;
wire n_1409;
wire n_1639;
wire n_1623;
wire n_183;
wire n_1015;
wire n_1503;
wire n_466;
wire n_1057;
wire n_603;
wire n_991;
wire n_1657;
wire n_235;
wire n_1126;
wire n_340;
wire n_710;
wire n_1108;
wire n_1182;
wire n_1298;
wire n_1611;
wire n_785;
wire n_746;
wire n_609;
wire n_1601;
wire n_1686;
wire n_167;
wire n_1356;
wire n_1589;
wire n_1740;
wire n_1497;
wire n_1168;
wire n_1216;
wire n_1320;
wire n_1430;
wire n_1316;
wire n_1287;
wire n_1452;
wire n_1622;
wire n_1586;
wire n_302;
wire n_1694;
wire n_380;
wire n_1535;
wire n_1596;
wire n_1190;
wire n_1734;
wire n_397;
wire n_1262;
wire n_218;
wire n_1213;
wire n_1350;
wire n_1673;
wire n_1715;
wire n_172;
wire n_1443;
wire n_1272;
wire n_239;
wire n_782;
wire n_1539;
wire n_490;
wire n_220;
wire n_809;
wire n_1043;
wire n_1608;
wire n_986;
wire n_1472;
wire n_1081;
wire n_402;
wire n_352;
wire n_1692;
wire n_800;
wire n_1084;
wire n_1171;
wire n_460;
wire n_1361;
wire n_1491;
wire n_662;
wire n_374;
wire n_1152;
wire n_1705;
wire n_450;
wire n_1684;
wire n_921;
wire n_1346;
wire n_711;
wire n_1642;
wire n_579;
wire n_1352;
wire n_937;
wire n_1682;
wire n_370;
wire n_1695;
wire n_650;
wire n_1046;
wire n_1145;
wire n_330;
wire n_1121;
wire n_1102;
wire n_972;
wire n_1405;
wire n_258;
wire n_1406;
wire n_456;
wire n_1332;
wire n_260;
wire n_313;
wire n_624;
wire n_962;
wire n_1041;
wire n_565;
wire n_356;
wire n_1569;
wire n_936;
wire n_1288;
wire n_1186;
wire n_1062;
wire n_885;
wire n_896;
wire n_654;
wire n_411;
wire n_1222;
wire n_599;
wire n_776;
wire n_321;
wire n_227;
wire n_1720;
wire n_204;
wire n_482;
wire n_934;
wire n_1637;
wire n_1407;
wire n_420;
wire n_1341;
wire n_394;
wire n_1456;
wire n_1489;
wire n_164;
wire n_942;
wire n_1524;
wire n_543;
wire n_1496;
wire n_1271;
wire n_1545;
wire n_1355;
wire n_1225;
wire n_1544;
wire n_1485;
wire n_325;
wire n_1640;
wire n_804;
wire n_464;
wire n_533;
wire n_806;
wire n_879;
wire n_959;
wire n_584;
wire n_244;
wire n_1343;
wire n_1522;
wire n_548;
wire n_282;
wire n_1676;
wire n_833;
wire n_1567;
wire n_523;
wire n_1319;
wire n_707;
wire n_345;
wire n_799;
wire n_1548;
wire n_1155;
wire n_273;
wire n_1633;
wire n_787;
wire n_1416;
wire n_1528;
wire n_1146;
wire n_159;
wire n_1086;
wire n_1066;
wire n_157;
wire n_1282;
wire n_550;
wire n_275;
wire n_652;
wire n_560;
wire n_1484;
wire n_1321;
wire n_1241;
wire n_1672;
wire n_569;
wire n_737;
wire n_1318;
wire n_1235;
wire n_1229;
wire n_306;
wire n_1292;
wire n_1373;
wire n_346;
wire n_1029;
wire n_1447;
wire n_790;
wire n_1706;
wire n_1498;
wire n_1210;
wire n_299;
wire n_1248;
wire n_1556;
wire n_902;
wire n_333;
wire n_1047;
wire n_1385;
wire n_431;
wire n_459;
wire n_1269;
wire n_502;
wire n_672;
wire n_1257;
wire n_285;
wire n_1375;
wire n_655;
wire n_706;
wire n_1045;
wire n_1650;
wire n_786;
wire n_1236;
wire n_1559;
wire n_1725;
wire n_834;
wire n_743;
wire n_766;
wire n_430;
wire n_1741;
wire n_1325;
wire n_1002;
wire n_1746;
wire n_545;
wire n_489;
wire n_1727;
wire n_251;
wire n_1019;
wire n_636;
wire n_729;
wire n_876;
wire n_774;
wire n_1337;
wire n_660;
wire n_438;
wire n_1477;
wire n_1360;
wire n_1200;
wire n_479;
wire n_1607;
wire n_1353;
wire n_1454;
wire n_869;
wire n_1154;
wire n_1113;
wire n_1600;
wire n_646;
wire n_528;
wire n_391;
wire n_1098;
wire n_1329;
wire n_817;
wire n_262;
wire n_187;
wire n_897;
wire n_846;
wire n_841;
wire n_1476;
wire n_1001;
wire n_508;
wire n_1050;
wire n_1411;
wire n_1463;
wire n_1177;
wire n_332;
wire n_1150;
wire n_1742;
wire n_1562;
wire n_1690;
wire n_398;
wire n_1191;
wire n_566;
wire n_1023;
wire n_1076;
wire n_1118;
wire n_194;
wire n_1007;
wire n_1378;
wire n_855;
wire n_1592;
wire n_1631;
wire n_591;
wire n_1377;
wire n_256;
wire n_853;
wire n_440;
wire n_695;
wire n_1542;
wire n_875;
wire n_209;
wire n_367;
wire n_680;
wire n_1678;
wire n_661;
wire n_1716;
wire n_278;
wire n_1256;
wire n_671;
wire n_933;
wire n_740;
wire n_703;
wire n_978;
wire n_384;
wire n_1291;
wire n_1217;
wire n_751;
wire n_749;
wire n_310;
wire n_1628;
wire n_1324;
wire n_1399;
wire n_1435;
wire n_969;
wire n_988;
wire n_1065;
wire n_1401;
wire n_1255;
wire n_568;
wire n_1516;
wire n_1536;
wire n_180;
wire n_1204;
wire n_823;
wire n_1132;
wire n_643;
wire n_233;
wire n_698;
wire n_1074;
wire n_1394;
wire n_1327;
wire n_1326;
wire n_739;
wire n_400;
wire n_955;
wire n_337;
wire n_1379;
wire n_214;
wire n_246;
wire n_1338;
wire n_1097;
wire n_935;
wire n_781;
wire n_789;
wire n_1554;
wire n_1130;
wire n_181;
wire n_182;
wire n_573;
wire n_769;
wire n_676;
wire n_327;
wire n_1120;
wire n_832;
wire n_1583;
wire n_1730;
wire n_555;
wire n_389;
wire n_814;
wire n_1643;
wire n_1729;
wire n_669;
wire n_176;
wire n_300;
wire n_222;
wire n_747;
wire n_1389;
wire n_1105;
wire n_721;
wire n_1461;
wire n_742;
wire n_691;
wire n_535;
wire n_372;
wire n_314;
wire n_1408;
wire n_378;
wire n_1196;
wire n_377;
wire n_1598;
wire n_863;
wire n_601;
wire n_338;
wire n_1283;
wire n_918;
wire n_748;
wire n_506;
wire n_1114;
wire n_763;
wire n_1147;
wire n_360;
wire n_1506;
wire n_1652;
wire n_957;
wire n_895;
wire n_866;
wire n_1227;
wire n_191;
wire n_387;
wire n_452;
wire n_744;
wire n_971;
wire n_946;
wire n_344;
wire n_761;
wire n_1303;
wire n_1205;
wire n_1258;
wire n_1392;
wire n_174;
wire n_1173;
wire n_525;
wire n_1677;
wire n_1116;
wire n_611;
wire n_1702;
wire n_1570;
wire n_1219;
wire n_1689;
wire n_1174;
wire n_1016;
wire n_1347;
wire n_795;
wire n_1501;
wire n_1221;
wire n_1245;
wire n_838;
wire n_647;
wire n_197;
wire n_844;
wire n_448;
wire n_1017;
wire n_1083;
wire n_445;
wire n_1561;
wire n_930;
wire n_888;
wire n_1112;
wire n_234;
wire n_910;
wire n_1656;
wire n_1721;
wire n_1460;
wire n_911;
wire n_1464;
wire n_236;
wire n_653;
wire n_1737;
wire n_1414;
wire n_908;
wire n_752;
wire n_944;
wire n_576;
wire n_1028;
wire n_472;
wire n_270;
wire n_414;
wire n_563;
wire n_1011;
wire n_1566;
wire n_1215;
wire n_839;
wire n_708;
wire n_668;
wire n_626;
wire n_990;
wire n_1500;
wire n_779;
wire n_1537;
wire n_1104;
wire n_854;
wire n_1058;
wire n_498;
wire n_1122;
wire n_870;
wire n_904;
wire n_1253;
wire n_709;
wire n_1266;
wire n_366;
wire n_1509;
wire n_1693;
wire n_1109;
wire n_185;
wire n_712;
wire n_348;
wire n_1276;
wire n_376;
wire n_390;
wire n_1148;
wire n_334;
wire n_1161;
wire n_1085;
wire n_232;
wire n_1239;
wire n_771;
wire n_1584;
wire n_470;
wire n_475;
wire n_924;
wire n_298;
wire n_1582;
wire n_492;
wire n_1149;
wire n_265;
wire n_1184;
wire n_228;
wire n_719;
wire n_1525;
wire n_455;
wire n_1585;
wire n_363;
wire n_1090;
wire n_592;
wire n_1518;
wire n_829;
wire n_1156;
wire n_1362;
wire n_393;
wire n_984;
wire n_503;
wire n_1450;
wire n_1638;
wire n_868;
wire n_570;
wire n_859;
wire n_406;
wire n_735;
wire n_878;
wire n_620;
wire n_519;
wire n_307;
wire n_469;
wire n_1218;
wire n_500;
wire n_1482;
wire n_981;
wire n_714;
wire n_1349;
wire n_291;
wire n_1144;
wire n_357;
wire n_985;
wire n_481;
wire n_997;
wire n_1710;
wire n_1301;
wire n_802;
wire n_561;
wire n_980;
wire n_1306;
wire n_1651;
wire n_1198;
wire n_1609;
wire n_436;
wire n_409;
wire n_1244;
wire n_1685;
wire n_1574;
wire n_240;
wire n_756;
wire n_1619;
wire n_1606;
wire n_810;
wire n_1133;
wire n_635;
wire n_1194;
wire n_1051;
wire n_253;
wire n_1552;
wire n_583;
wire n_249;
wire n_201;
wire n_1039;
wire n_1442;
wire n_1034;
wire n_1480;
wire n_1158;
wire n_754;
wire n_941;
wire n_975;
wire n_1031;
wire n_1305;
wire n_553;
wire n_849;
wire n_753;
wire n_467;
wire n_269;
wire n_359;
wire n_973;
wire n_1479;
wire n_1055;
wire n_1675;
wire n_582;
wire n_861;
wire n_857;
wire n_967;
wire n_571;
wire n_404;
wire n_271;
wire n_158;
wire n_206;
wire n_679;
wire n_633;
wire n_1170;
wire n_665;
wire n_1629;
wire n_588;
wire n_225;
wire n_1260;
wire n_308;
wire n_309;
wire n_1010;
wire n_1040;
wire n_915;
wire n_632;
wire n_1166;
wire n_812;
wire n_1131;
wire n_534;
wire n_1578;
wire n_1006;
wire n_373;
wire n_1632;
wire n_257;
wire n_1557;
wire n_730;
wire n_1311;
wire n_1494;
wire n_670;
wire n_203;
wire n_207;
wire n_1089;
wire n_1587;
wire n_1365;
wire n_1417;
wire n_205;
wire n_1242;
wire n_681;
wire n_1226;
wire n_1274;
wire n_1486;
wire n_412;
wire n_640;
wire n_1322;
wire n_965;
wire n_1428;
wire n_1616;
wire n_1576;
wire n_339;
wire n_784;
wire n_315;
wire n_434;
wire n_288;
wire n_1059;
wire n_1197;
wire n_422;
wire n_722;
wire n_862;
wire n_165;
wire n_540;
wire n_1423;
wire n_457;
wire n_364;
wire n_629;
wire n_1621;
wire n_1748;
wire n_900;
wire n_1449;
wire n_531;
wire n_827;
wire n_361;
wire n_1025;
wire n_336;
wire n_1013;
wire n_1259;
wire n_192;
wire n_1538;
wire n_649;
wire n_1612;
wire n_1240;

CKINVDCx5p33_ASAP7_75t_R g155 ( 
.A(n_82),
.Y(n_155)
);

CKINVDCx5p33_ASAP7_75t_R g156 ( 
.A(n_35),
.Y(n_156)
);

CKINVDCx5p33_ASAP7_75t_R g157 ( 
.A(n_107),
.Y(n_157)
);

INVx2_ASAP7_75t_SL g158 ( 
.A(n_29),
.Y(n_158)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_26),
.Y(n_159)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_39),
.Y(n_160)
);

CKINVDCx5p33_ASAP7_75t_R g161 ( 
.A(n_151),
.Y(n_161)
);

CKINVDCx5p33_ASAP7_75t_R g162 ( 
.A(n_9),
.Y(n_162)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_55),
.Y(n_163)
);

CKINVDCx5p33_ASAP7_75t_R g164 ( 
.A(n_120),
.Y(n_164)
);

CKINVDCx5p33_ASAP7_75t_R g165 ( 
.A(n_39),
.Y(n_165)
);

CKINVDCx5p33_ASAP7_75t_R g166 ( 
.A(n_9),
.Y(n_166)
);

CKINVDCx5p33_ASAP7_75t_R g167 ( 
.A(n_141),
.Y(n_167)
);

CKINVDCx5p33_ASAP7_75t_R g168 ( 
.A(n_45),
.Y(n_168)
);

CKINVDCx5p33_ASAP7_75t_R g169 ( 
.A(n_57),
.Y(n_169)
);

INVx2_ASAP7_75t_L g170 ( 
.A(n_25),
.Y(n_170)
);

CKINVDCx20_ASAP7_75t_R g171 ( 
.A(n_100),
.Y(n_171)
);

CKINVDCx20_ASAP7_75t_R g172 ( 
.A(n_64),
.Y(n_172)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_22),
.Y(n_173)
);

CKINVDCx20_ASAP7_75t_R g174 ( 
.A(n_57),
.Y(n_174)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_153),
.Y(n_175)
);

CKINVDCx5p33_ASAP7_75t_R g176 ( 
.A(n_142),
.Y(n_176)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_71),
.Y(n_177)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_18),
.Y(n_178)
);

CKINVDCx5p33_ASAP7_75t_R g179 ( 
.A(n_14),
.Y(n_179)
);

CKINVDCx5p33_ASAP7_75t_R g180 ( 
.A(n_132),
.Y(n_180)
);

CKINVDCx5p33_ASAP7_75t_R g181 ( 
.A(n_146),
.Y(n_181)
);

CKINVDCx5p33_ASAP7_75t_R g182 ( 
.A(n_111),
.Y(n_182)
);

CKINVDCx5p33_ASAP7_75t_R g183 ( 
.A(n_93),
.Y(n_183)
);

CKINVDCx5p33_ASAP7_75t_R g184 ( 
.A(n_68),
.Y(n_184)
);

CKINVDCx5p33_ASAP7_75t_R g185 ( 
.A(n_86),
.Y(n_185)
);

INVx1_ASAP7_75t_SL g186 ( 
.A(n_16),
.Y(n_186)
);

CKINVDCx5p33_ASAP7_75t_R g187 ( 
.A(n_38),
.Y(n_187)
);

INVx2_ASAP7_75t_L g188 ( 
.A(n_80),
.Y(n_188)
);

CKINVDCx5p33_ASAP7_75t_R g189 ( 
.A(n_1),
.Y(n_189)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_53),
.Y(n_190)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_26),
.Y(n_191)
);

CKINVDCx5p33_ASAP7_75t_R g192 ( 
.A(n_0),
.Y(n_192)
);

CKINVDCx5p33_ASAP7_75t_R g193 ( 
.A(n_122),
.Y(n_193)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_134),
.Y(n_194)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_102),
.Y(n_195)
);

INVx2_ASAP7_75t_L g196 ( 
.A(n_91),
.Y(n_196)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_118),
.Y(n_197)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_88),
.Y(n_198)
);

CKINVDCx14_ASAP7_75t_R g199 ( 
.A(n_25),
.Y(n_199)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_50),
.Y(n_200)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_112),
.Y(n_201)
);

CKINVDCx5p33_ASAP7_75t_R g202 ( 
.A(n_116),
.Y(n_202)
);

BUFx5_ASAP7_75t_L g203 ( 
.A(n_32),
.Y(n_203)
);

CKINVDCx20_ASAP7_75t_R g204 ( 
.A(n_0),
.Y(n_204)
);

CKINVDCx5p33_ASAP7_75t_R g205 ( 
.A(n_124),
.Y(n_205)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_136),
.Y(n_206)
);

BUFx10_ASAP7_75t_L g207 ( 
.A(n_42),
.Y(n_207)
);

CKINVDCx5p33_ASAP7_75t_R g208 ( 
.A(n_117),
.Y(n_208)
);

CKINVDCx5p33_ASAP7_75t_R g209 ( 
.A(n_123),
.Y(n_209)
);

CKINVDCx20_ASAP7_75t_R g210 ( 
.A(n_97),
.Y(n_210)
);

HB1xp67_ASAP7_75t_L g211 ( 
.A(n_121),
.Y(n_211)
);

CKINVDCx5p33_ASAP7_75t_R g212 ( 
.A(n_23),
.Y(n_212)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_33),
.Y(n_213)
);

CKINVDCx5p33_ASAP7_75t_R g214 ( 
.A(n_5),
.Y(n_214)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_67),
.Y(n_215)
);

CKINVDCx5p33_ASAP7_75t_R g216 ( 
.A(n_24),
.Y(n_216)
);

BUFx8_ASAP7_75t_SL g217 ( 
.A(n_16),
.Y(n_217)
);

CKINVDCx5p33_ASAP7_75t_R g218 ( 
.A(n_30),
.Y(n_218)
);

CKINVDCx5p33_ASAP7_75t_R g219 ( 
.A(n_8),
.Y(n_219)
);

CKINVDCx5p33_ASAP7_75t_R g220 ( 
.A(n_40),
.Y(n_220)
);

CKINVDCx5p33_ASAP7_75t_R g221 ( 
.A(n_110),
.Y(n_221)
);

BUFx3_ASAP7_75t_L g222 ( 
.A(n_19),
.Y(n_222)
);

CKINVDCx5p33_ASAP7_75t_R g223 ( 
.A(n_144),
.Y(n_223)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_128),
.Y(n_224)
);

CKINVDCx5p33_ASAP7_75t_R g225 ( 
.A(n_53),
.Y(n_225)
);

CKINVDCx5p33_ASAP7_75t_R g226 ( 
.A(n_131),
.Y(n_226)
);

CKINVDCx5p33_ASAP7_75t_R g227 ( 
.A(n_1),
.Y(n_227)
);

CKINVDCx20_ASAP7_75t_R g228 ( 
.A(n_55),
.Y(n_228)
);

CKINVDCx20_ASAP7_75t_R g229 ( 
.A(n_139),
.Y(n_229)
);

CKINVDCx5p33_ASAP7_75t_R g230 ( 
.A(n_149),
.Y(n_230)
);

CKINVDCx5p33_ASAP7_75t_R g231 ( 
.A(n_119),
.Y(n_231)
);

BUFx5_ASAP7_75t_L g232 ( 
.A(n_14),
.Y(n_232)
);

BUFx6f_ASAP7_75t_L g233 ( 
.A(n_114),
.Y(n_233)
);

CKINVDCx5p33_ASAP7_75t_R g234 ( 
.A(n_109),
.Y(n_234)
);

INVx1_ASAP7_75t_SL g235 ( 
.A(n_83),
.Y(n_235)
);

BUFx6f_ASAP7_75t_L g236 ( 
.A(n_72),
.Y(n_236)
);

CKINVDCx5p33_ASAP7_75t_R g237 ( 
.A(n_42),
.Y(n_237)
);

INVx3_ASAP7_75t_L g238 ( 
.A(n_22),
.Y(n_238)
);

INVx2_ASAP7_75t_L g239 ( 
.A(n_150),
.Y(n_239)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_17),
.Y(n_240)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_74),
.Y(n_241)
);

CKINVDCx5p33_ASAP7_75t_R g242 ( 
.A(n_47),
.Y(n_242)
);

CKINVDCx5p33_ASAP7_75t_R g243 ( 
.A(n_63),
.Y(n_243)
);

CKINVDCx16_ASAP7_75t_R g244 ( 
.A(n_17),
.Y(n_244)
);

CKINVDCx5p33_ASAP7_75t_R g245 ( 
.A(n_50),
.Y(n_245)
);

CKINVDCx5p33_ASAP7_75t_R g246 ( 
.A(n_49),
.Y(n_246)
);

CKINVDCx20_ASAP7_75t_R g247 ( 
.A(n_133),
.Y(n_247)
);

CKINVDCx20_ASAP7_75t_R g248 ( 
.A(n_62),
.Y(n_248)
);

CKINVDCx5p33_ASAP7_75t_R g249 ( 
.A(n_138),
.Y(n_249)
);

INVx2_ASAP7_75t_SL g250 ( 
.A(n_5),
.Y(n_250)
);

CKINVDCx5p33_ASAP7_75t_R g251 ( 
.A(n_3),
.Y(n_251)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_34),
.Y(n_252)
);

CKINVDCx14_ASAP7_75t_R g253 ( 
.A(n_13),
.Y(n_253)
);

CKINVDCx14_ASAP7_75t_R g254 ( 
.A(n_94),
.Y(n_254)
);

CKINVDCx20_ASAP7_75t_R g255 ( 
.A(n_20),
.Y(n_255)
);

CKINVDCx5p33_ASAP7_75t_R g256 ( 
.A(n_28),
.Y(n_256)
);

BUFx6f_ASAP7_75t_L g257 ( 
.A(n_147),
.Y(n_257)
);

BUFx3_ASAP7_75t_L g258 ( 
.A(n_103),
.Y(n_258)
);

CKINVDCx20_ASAP7_75t_R g259 ( 
.A(n_44),
.Y(n_259)
);

CKINVDCx5p33_ASAP7_75t_R g260 ( 
.A(n_84),
.Y(n_260)
);

CKINVDCx5p33_ASAP7_75t_R g261 ( 
.A(n_75),
.Y(n_261)
);

CKINVDCx5p33_ASAP7_75t_R g262 ( 
.A(n_99),
.Y(n_262)
);

CKINVDCx5p33_ASAP7_75t_R g263 ( 
.A(n_64),
.Y(n_263)
);

CKINVDCx5p33_ASAP7_75t_R g264 ( 
.A(n_40),
.Y(n_264)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_89),
.Y(n_265)
);

CKINVDCx5p33_ASAP7_75t_R g266 ( 
.A(n_98),
.Y(n_266)
);

CKINVDCx5p33_ASAP7_75t_R g267 ( 
.A(n_113),
.Y(n_267)
);

CKINVDCx5p33_ASAP7_75t_R g268 ( 
.A(n_41),
.Y(n_268)
);

CKINVDCx5p33_ASAP7_75t_R g269 ( 
.A(n_106),
.Y(n_269)
);

BUFx2_ASAP7_75t_L g270 ( 
.A(n_108),
.Y(n_270)
);

CKINVDCx5p33_ASAP7_75t_R g271 ( 
.A(n_6),
.Y(n_271)
);

CKINVDCx5p33_ASAP7_75t_R g272 ( 
.A(n_61),
.Y(n_272)
);

BUFx6f_ASAP7_75t_L g273 ( 
.A(n_69),
.Y(n_273)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_101),
.Y(n_274)
);

CKINVDCx20_ASAP7_75t_R g275 ( 
.A(n_87),
.Y(n_275)
);

BUFx5_ASAP7_75t_L g276 ( 
.A(n_92),
.Y(n_276)
);

CKINVDCx5p33_ASAP7_75t_R g277 ( 
.A(n_135),
.Y(n_277)
);

CKINVDCx5p33_ASAP7_75t_R g278 ( 
.A(n_54),
.Y(n_278)
);

HB1xp67_ASAP7_75t_L g279 ( 
.A(n_59),
.Y(n_279)
);

CKINVDCx5p33_ASAP7_75t_R g280 ( 
.A(n_152),
.Y(n_280)
);

CKINVDCx5p33_ASAP7_75t_R g281 ( 
.A(n_19),
.Y(n_281)
);

CKINVDCx5p33_ASAP7_75t_R g282 ( 
.A(n_4),
.Y(n_282)
);

CKINVDCx5p33_ASAP7_75t_R g283 ( 
.A(n_58),
.Y(n_283)
);

CKINVDCx5p33_ASAP7_75t_R g284 ( 
.A(n_4),
.Y(n_284)
);

CKINVDCx5p33_ASAP7_75t_R g285 ( 
.A(n_54),
.Y(n_285)
);

CKINVDCx20_ASAP7_75t_R g286 ( 
.A(n_7),
.Y(n_286)
);

CKINVDCx5p33_ASAP7_75t_R g287 ( 
.A(n_130),
.Y(n_287)
);

CKINVDCx5p33_ASAP7_75t_R g288 ( 
.A(n_105),
.Y(n_288)
);

CKINVDCx5p33_ASAP7_75t_R g289 ( 
.A(n_127),
.Y(n_289)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_32),
.Y(n_290)
);

CKINVDCx5p33_ASAP7_75t_R g291 ( 
.A(n_35),
.Y(n_291)
);

INVxp67_ASAP7_75t_L g292 ( 
.A(n_7),
.Y(n_292)
);

CKINVDCx16_ASAP7_75t_R g293 ( 
.A(n_33),
.Y(n_293)
);

CKINVDCx5p33_ASAP7_75t_R g294 ( 
.A(n_65),
.Y(n_294)
);

CKINVDCx5p33_ASAP7_75t_R g295 ( 
.A(n_76),
.Y(n_295)
);

CKINVDCx5p33_ASAP7_75t_R g296 ( 
.A(n_125),
.Y(n_296)
);

CKINVDCx5p33_ASAP7_75t_R g297 ( 
.A(n_95),
.Y(n_297)
);

CKINVDCx5p33_ASAP7_75t_R g298 ( 
.A(n_145),
.Y(n_298)
);

CKINVDCx5p33_ASAP7_75t_R g299 ( 
.A(n_129),
.Y(n_299)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_52),
.Y(n_300)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_73),
.Y(n_301)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_154),
.Y(n_302)
);

CKINVDCx5p33_ASAP7_75t_R g303 ( 
.A(n_137),
.Y(n_303)
);

CKINVDCx5p33_ASAP7_75t_R g304 ( 
.A(n_13),
.Y(n_304)
);

CKINVDCx5p33_ASAP7_75t_R g305 ( 
.A(n_70),
.Y(n_305)
);

CKINVDCx5p33_ASAP7_75t_R g306 ( 
.A(n_148),
.Y(n_306)
);

INVx2_ASAP7_75t_SL g307 ( 
.A(n_62),
.Y(n_307)
);

CKINVDCx5p33_ASAP7_75t_R g308 ( 
.A(n_217),
.Y(n_308)
);

INVxp67_ASAP7_75t_L g309 ( 
.A(n_279),
.Y(n_309)
);

CKINVDCx5p33_ASAP7_75t_R g310 ( 
.A(n_183),
.Y(n_310)
);

NOR2xp33_ASAP7_75t_L g311 ( 
.A(n_270),
.B(n_2),
.Y(n_311)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_203),
.Y(n_312)
);

INVxp67_ASAP7_75t_L g313 ( 
.A(n_207),
.Y(n_313)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_203),
.Y(n_314)
);

CKINVDCx16_ASAP7_75t_R g315 ( 
.A(n_199),
.Y(n_315)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_203),
.Y(n_316)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_203),
.Y(n_317)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_203),
.Y(n_318)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_203),
.Y(n_319)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_203),
.Y(n_320)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_203),
.Y(n_321)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_232),
.Y(n_322)
);

CKINVDCx5p33_ASAP7_75t_R g323 ( 
.A(n_184),
.Y(n_323)
);

CKINVDCx5p33_ASAP7_75t_R g324 ( 
.A(n_185),
.Y(n_324)
);

CKINVDCx5p33_ASAP7_75t_R g325 ( 
.A(n_193),
.Y(n_325)
);

NOR2xp33_ASAP7_75t_L g326 ( 
.A(n_211),
.B(n_2),
.Y(n_326)
);

NOR2xp67_ASAP7_75t_L g327 ( 
.A(n_238),
.B(n_3),
.Y(n_327)
);

INVx2_ASAP7_75t_L g328 ( 
.A(n_232),
.Y(n_328)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_232),
.Y(n_329)
);

NOR2x1_ASAP7_75t_L g330 ( 
.A(n_258),
.B(n_6),
.Y(n_330)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_232),
.Y(n_331)
);

NAND2xp5_ASAP7_75t_L g332 ( 
.A(n_253),
.B(n_8),
.Y(n_332)
);

CKINVDCx5p33_ASAP7_75t_R g333 ( 
.A(n_202),
.Y(n_333)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_232),
.Y(n_334)
);

CKINVDCx20_ASAP7_75t_R g335 ( 
.A(n_171),
.Y(n_335)
);

INVxp67_ASAP7_75t_SL g336 ( 
.A(n_238),
.Y(n_336)
);

CKINVDCx5p33_ASAP7_75t_R g337 ( 
.A(n_205),
.Y(n_337)
);

INVx1_ASAP7_75t_L g338 ( 
.A(n_232),
.Y(n_338)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_232),
.Y(n_339)
);

CKINVDCx5p33_ASAP7_75t_R g340 ( 
.A(n_208),
.Y(n_340)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_232),
.Y(n_341)
);

INVxp67_ASAP7_75t_SL g342 ( 
.A(n_238),
.Y(n_342)
);

CKINVDCx20_ASAP7_75t_R g343 ( 
.A(n_210),
.Y(n_343)
);

OR2x2_ASAP7_75t_L g344 ( 
.A(n_159),
.B(n_10),
.Y(n_344)
);

INVx1_ASAP7_75t_L g345 ( 
.A(n_170),
.Y(n_345)
);

INVx1_ASAP7_75t_L g346 ( 
.A(n_170),
.Y(n_346)
);

INVx1_ASAP7_75t_L g347 ( 
.A(n_222),
.Y(n_347)
);

INVx1_ASAP7_75t_L g348 ( 
.A(n_222),
.Y(n_348)
);

INVx1_ASAP7_75t_L g349 ( 
.A(n_160),
.Y(n_349)
);

NOR2xp67_ASAP7_75t_L g350 ( 
.A(n_307),
.B(n_10),
.Y(n_350)
);

INVxp67_ASAP7_75t_SL g351 ( 
.A(n_258),
.Y(n_351)
);

INVx1_ASAP7_75t_L g352 ( 
.A(n_163),
.Y(n_352)
);

CKINVDCx20_ASAP7_75t_R g353 ( 
.A(n_229),
.Y(n_353)
);

CKINVDCx16_ASAP7_75t_R g354 ( 
.A(n_244),
.Y(n_354)
);

INVx1_ASAP7_75t_L g355 ( 
.A(n_173),
.Y(n_355)
);

CKINVDCx5p33_ASAP7_75t_R g356 ( 
.A(n_209),
.Y(n_356)
);

CKINVDCx20_ASAP7_75t_R g357 ( 
.A(n_247),
.Y(n_357)
);

CKINVDCx5p33_ASAP7_75t_R g358 ( 
.A(n_221),
.Y(n_358)
);

INVx1_ASAP7_75t_L g359 ( 
.A(n_178),
.Y(n_359)
);

INVx1_ASAP7_75t_L g360 ( 
.A(n_190),
.Y(n_360)
);

INVx1_ASAP7_75t_L g361 ( 
.A(n_191),
.Y(n_361)
);

CKINVDCx20_ASAP7_75t_R g362 ( 
.A(n_275),
.Y(n_362)
);

INVx1_ASAP7_75t_L g363 ( 
.A(n_200),
.Y(n_363)
);

INVxp67_ASAP7_75t_SL g364 ( 
.A(n_175),
.Y(n_364)
);

INVx1_ASAP7_75t_L g365 ( 
.A(n_213),
.Y(n_365)
);

INVx1_ASAP7_75t_L g366 ( 
.A(n_240),
.Y(n_366)
);

CKINVDCx20_ASAP7_75t_R g367 ( 
.A(n_254),
.Y(n_367)
);

CKINVDCx5p33_ASAP7_75t_R g368 ( 
.A(n_223),
.Y(n_368)
);

INVx1_ASAP7_75t_L g369 ( 
.A(n_252),
.Y(n_369)
);

INVx1_ASAP7_75t_L g370 ( 
.A(n_290),
.Y(n_370)
);

INVx1_ASAP7_75t_L g371 ( 
.A(n_300),
.Y(n_371)
);

INVxp67_ASAP7_75t_L g372 ( 
.A(n_207),
.Y(n_372)
);

CKINVDCx5p33_ASAP7_75t_R g373 ( 
.A(n_226),
.Y(n_373)
);

INVxp67_ASAP7_75t_SL g374 ( 
.A(n_177),
.Y(n_374)
);

NAND2xp5_ASAP7_75t_L g375 ( 
.A(n_158),
.B(n_11),
.Y(n_375)
);

AND2x2_ASAP7_75t_L g376 ( 
.A(n_158),
.B(n_11),
.Y(n_376)
);

CKINVDCx5p33_ASAP7_75t_R g377 ( 
.A(n_230),
.Y(n_377)
);

INVx1_ASAP7_75t_L g378 ( 
.A(n_250),
.Y(n_378)
);

HB1xp67_ASAP7_75t_L g379 ( 
.A(n_293),
.Y(n_379)
);

INVxp67_ASAP7_75t_SL g380 ( 
.A(n_194),
.Y(n_380)
);

CKINVDCx5p33_ASAP7_75t_R g381 ( 
.A(n_231),
.Y(n_381)
);

CKINVDCx20_ASAP7_75t_R g382 ( 
.A(n_234),
.Y(n_382)
);

CKINVDCx5p33_ASAP7_75t_R g383 ( 
.A(n_249),
.Y(n_383)
);

BUFx2_ASAP7_75t_L g384 ( 
.A(n_379),
.Y(n_384)
);

INVx1_ASAP7_75t_L g385 ( 
.A(n_328),
.Y(n_385)
);

AND2x4_ASAP7_75t_L g386 ( 
.A(n_327),
.B(n_188),
.Y(n_386)
);

NAND2xp5_ASAP7_75t_L g387 ( 
.A(n_336),
.B(n_155),
.Y(n_387)
);

INVx1_ASAP7_75t_L g388 ( 
.A(n_312),
.Y(n_388)
);

INVx1_ASAP7_75t_L g389 ( 
.A(n_312),
.Y(n_389)
);

AND2x2_ASAP7_75t_L g390 ( 
.A(n_342),
.B(n_364),
.Y(n_390)
);

NAND2xp5_ASAP7_75t_L g391 ( 
.A(n_374),
.B(n_155),
.Y(n_391)
);

AND2x2_ASAP7_75t_L g392 ( 
.A(n_380),
.B(n_351),
.Y(n_392)
);

NAND2xp5_ASAP7_75t_L g393 ( 
.A(n_314),
.B(n_157),
.Y(n_393)
);

INVx2_ASAP7_75t_L g394 ( 
.A(n_328),
.Y(n_394)
);

INVx2_ASAP7_75t_L g395 ( 
.A(n_328),
.Y(n_395)
);

OAI22xp33_ASAP7_75t_L g396 ( 
.A1(n_354),
.A2(n_204),
.B1(n_286),
.B2(n_259),
.Y(n_396)
);

INVx2_ASAP7_75t_L g397 ( 
.A(n_314),
.Y(n_397)
);

INVx1_ASAP7_75t_L g398 ( 
.A(n_316),
.Y(n_398)
);

INVxp67_ASAP7_75t_L g399 ( 
.A(n_347),
.Y(n_399)
);

BUFx6f_ASAP7_75t_L g400 ( 
.A(n_316),
.Y(n_400)
);

INVx2_ASAP7_75t_L g401 ( 
.A(n_317),
.Y(n_401)
);

INVx2_ASAP7_75t_L g402 ( 
.A(n_317),
.Y(n_402)
);

INVx2_ASAP7_75t_L g403 ( 
.A(n_318),
.Y(n_403)
);

AND2x2_ASAP7_75t_SL g404 ( 
.A(n_376),
.B(n_188),
.Y(n_404)
);

INVx1_ASAP7_75t_L g405 ( 
.A(n_318),
.Y(n_405)
);

NAND2xp5_ASAP7_75t_L g406 ( 
.A(n_319),
.B(n_157),
.Y(n_406)
);

INVx2_ASAP7_75t_L g407 ( 
.A(n_319),
.Y(n_407)
);

AND2x2_ASAP7_75t_L g408 ( 
.A(n_376),
.B(n_196),
.Y(n_408)
);

INVx2_ASAP7_75t_L g409 ( 
.A(n_320),
.Y(n_409)
);

INVxp67_ASAP7_75t_L g410 ( 
.A(n_347),
.Y(n_410)
);

CKINVDCx20_ASAP7_75t_R g411 ( 
.A(n_335),
.Y(n_411)
);

NAND2xp5_ASAP7_75t_L g412 ( 
.A(n_320),
.B(n_161),
.Y(n_412)
);

NAND2xp5_ASAP7_75t_L g413 ( 
.A(n_321),
.B(n_161),
.Y(n_413)
);

INVx1_ASAP7_75t_L g414 ( 
.A(n_321),
.Y(n_414)
);

INVxp67_ASAP7_75t_SL g415 ( 
.A(n_348),
.Y(n_415)
);

INVx2_ASAP7_75t_L g416 ( 
.A(n_322),
.Y(n_416)
);

BUFx6f_ASAP7_75t_L g417 ( 
.A(n_322),
.Y(n_417)
);

INVx2_ASAP7_75t_L g418 ( 
.A(n_329),
.Y(n_418)
);

INVx3_ASAP7_75t_L g419 ( 
.A(n_329),
.Y(n_419)
);

BUFx6f_ASAP7_75t_L g420 ( 
.A(n_331),
.Y(n_420)
);

INVx1_ASAP7_75t_L g421 ( 
.A(n_331),
.Y(n_421)
);

AND2x4_ASAP7_75t_L g422 ( 
.A(n_327),
.B(n_196),
.Y(n_422)
);

AND2x4_ASAP7_75t_L g423 ( 
.A(n_334),
.B(n_239),
.Y(n_423)
);

AND2x4_ASAP7_75t_L g424 ( 
.A(n_334),
.B(n_239),
.Y(n_424)
);

AND2x2_ASAP7_75t_L g425 ( 
.A(n_348),
.B(n_338),
.Y(n_425)
);

AND2x2_ASAP7_75t_L g426 ( 
.A(n_338),
.B(n_250),
.Y(n_426)
);

INVx1_ASAP7_75t_L g427 ( 
.A(n_339),
.Y(n_427)
);

OR2x6_ASAP7_75t_L g428 ( 
.A(n_330),
.B(n_307),
.Y(n_428)
);

INVx1_ASAP7_75t_L g429 ( 
.A(n_339),
.Y(n_429)
);

BUFx6f_ASAP7_75t_L g430 ( 
.A(n_341),
.Y(n_430)
);

BUFx6f_ASAP7_75t_L g431 ( 
.A(n_341),
.Y(n_431)
);

AND2x4_ASAP7_75t_L g432 ( 
.A(n_330),
.B(n_233),
.Y(n_432)
);

INVx1_ASAP7_75t_L g433 ( 
.A(n_349),
.Y(n_433)
);

INVx2_ASAP7_75t_L g434 ( 
.A(n_345),
.Y(n_434)
);

INVx1_ASAP7_75t_L g435 ( 
.A(n_349),
.Y(n_435)
);

INVx2_ASAP7_75t_L g436 ( 
.A(n_345),
.Y(n_436)
);

INVx1_ASAP7_75t_L g437 ( 
.A(n_352),
.Y(n_437)
);

INVx2_ASAP7_75t_L g438 ( 
.A(n_346),
.Y(n_438)
);

INVx1_ASAP7_75t_L g439 ( 
.A(n_352),
.Y(n_439)
);

NOR2xp33_ASAP7_75t_SL g440 ( 
.A(n_315),
.B(n_207),
.Y(n_440)
);

NAND2xp33_ASAP7_75t_L g441 ( 
.A(n_332),
.B(n_233),
.Y(n_441)
);

BUFx2_ASAP7_75t_L g442 ( 
.A(n_313),
.Y(n_442)
);

INVx6_ASAP7_75t_L g443 ( 
.A(n_344),
.Y(n_443)
);

INVx1_ASAP7_75t_L g444 ( 
.A(n_355),
.Y(n_444)
);

AND2x4_ASAP7_75t_L g445 ( 
.A(n_350),
.B(n_233),
.Y(n_445)
);

BUFx8_ASAP7_75t_L g446 ( 
.A(n_344),
.Y(n_446)
);

INVx1_ASAP7_75t_L g447 ( 
.A(n_346),
.Y(n_447)
);

INVx1_ASAP7_75t_L g448 ( 
.A(n_355),
.Y(n_448)
);

BUFx2_ASAP7_75t_L g449 ( 
.A(n_372),
.Y(n_449)
);

NAND2xp5_ASAP7_75t_L g450 ( 
.A(n_378),
.B(n_164),
.Y(n_450)
);

AND3x1_ASAP7_75t_L g451 ( 
.A(n_326),
.B(n_197),
.C(n_195),
.Y(n_451)
);

INVx1_ASAP7_75t_L g452 ( 
.A(n_359),
.Y(n_452)
);

INVx2_ASAP7_75t_SL g453 ( 
.A(n_443),
.Y(n_453)
);

INVx2_ASAP7_75t_L g454 ( 
.A(n_394),
.Y(n_454)
);

NAND2xp5_ASAP7_75t_L g455 ( 
.A(n_404),
.B(n_310),
.Y(n_455)
);

INVx1_ASAP7_75t_L g456 ( 
.A(n_388),
.Y(n_456)
);

AND2x2_ASAP7_75t_SL g457 ( 
.A(n_404),
.B(n_311),
.Y(n_457)
);

INVx4_ASAP7_75t_L g458 ( 
.A(n_400),
.Y(n_458)
);

NOR2xp33_ASAP7_75t_L g459 ( 
.A(n_387),
.B(n_323),
.Y(n_459)
);

BUFx3_ASAP7_75t_L g460 ( 
.A(n_425),
.Y(n_460)
);

NAND2xp5_ASAP7_75t_L g461 ( 
.A(n_404),
.B(n_324),
.Y(n_461)
);

CKINVDCx20_ASAP7_75t_R g462 ( 
.A(n_411),
.Y(n_462)
);

INVx1_ASAP7_75t_SL g463 ( 
.A(n_411),
.Y(n_463)
);

INVx2_ASAP7_75t_L g464 ( 
.A(n_394),
.Y(n_464)
);

INVx1_ASAP7_75t_L g465 ( 
.A(n_388),
.Y(n_465)
);

INVx1_ASAP7_75t_L g466 ( 
.A(n_389),
.Y(n_466)
);

AND2x2_ASAP7_75t_SL g467 ( 
.A(n_404),
.B(n_233),
.Y(n_467)
);

OAI22xp33_ASAP7_75t_L g468 ( 
.A1(n_440),
.A2(n_315),
.B1(n_375),
.B2(n_186),
.Y(n_468)
);

NAND2xp5_ASAP7_75t_SL g469 ( 
.A(n_440),
.B(n_325),
.Y(n_469)
);

CKINVDCx5p33_ASAP7_75t_R g470 ( 
.A(n_442),
.Y(n_470)
);

INVx3_ASAP7_75t_L g471 ( 
.A(n_400),
.Y(n_471)
);

NAND2xp5_ASAP7_75t_L g472 ( 
.A(n_392),
.B(n_333),
.Y(n_472)
);

INVx1_ASAP7_75t_L g473 ( 
.A(n_389),
.Y(n_473)
);

NAND2xp33_ASAP7_75t_SL g474 ( 
.A(n_442),
.B(n_367),
.Y(n_474)
);

INVx1_ASAP7_75t_L g475 ( 
.A(n_398),
.Y(n_475)
);

AOI22xp33_ASAP7_75t_L g476 ( 
.A1(n_443),
.A2(n_375),
.B1(n_350),
.B2(n_309),
.Y(n_476)
);

INVx1_ASAP7_75t_L g477 ( 
.A(n_398),
.Y(n_477)
);

INVx3_ASAP7_75t_L g478 ( 
.A(n_400),
.Y(n_478)
);

AND2x2_ASAP7_75t_L g479 ( 
.A(n_426),
.B(n_378),
.Y(n_479)
);

INVx4_ASAP7_75t_L g480 ( 
.A(n_400),
.Y(n_480)
);

NAND2xp5_ASAP7_75t_L g481 ( 
.A(n_392),
.B(n_337),
.Y(n_481)
);

NOR2xp33_ASAP7_75t_L g482 ( 
.A(n_387),
.B(n_340),
.Y(n_482)
);

NAND2xp5_ASAP7_75t_L g483 ( 
.A(n_392),
.B(n_356),
.Y(n_483)
);

INVx3_ASAP7_75t_L g484 ( 
.A(n_400),
.Y(n_484)
);

INVx3_ASAP7_75t_L g485 ( 
.A(n_400),
.Y(n_485)
);

NAND2xp5_ASAP7_75t_L g486 ( 
.A(n_408),
.B(n_358),
.Y(n_486)
);

BUFx6f_ASAP7_75t_L g487 ( 
.A(n_400),
.Y(n_487)
);

OR2x6_ASAP7_75t_L g488 ( 
.A(n_428),
.B(n_198),
.Y(n_488)
);

NOR2xp33_ASAP7_75t_L g489 ( 
.A(n_443),
.B(n_368),
.Y(n_489)
);

BUFx10_ASAP7_75t_L g490 ( 
.A(n_443),
.Y(n_490)
);

INVx5_ASAP7_75t_L g491 ( 
.A(n_400),
.Y(n_491)
);

AOI22xp33_ASAP7_75t_L g492 ( 
.A1(n_443),
.A2(n_233),
.B1(n_273),
.B2(n_236),
.Y(n_492)
);

BUFx2_ASAP7_75t_L g493 ( 
.A(n_384),
.Y(n_493)
);

AND2x2_ASAP7_75t_L g494 ( 
.A(n_426),
.B(n_425),
.Y(n_494)
);

INVx2_ASAP7_75t_L g495 ( 
.A(n_394),
.Y(n_495)
);

NAND2x1p5_ASAP7_75t_L g496 ( 
.A(n_432),
.B(n_201),
.Y(n_496)
);

INVx1_ASAP7_75t_L g497 ( 
.A(n_405),
.Y(n_497)
);

INVx3_ASAP7_75t_L g498 ( 
.A(n_417),
.Y(n_498)
);

INVx4_ASAP7_75t_L g499 ( 
.A(n_417),
.Y(n_499)
);

NOR2xp33_ASAP7_75t_L g500 ( 
.A(n_443),
.B(n_373),
.Y(n_500)
);

INVx3_ASAP7_75t_L g501 ( 
.A(n_417),
.Y(n_501)
);

INVx1_ASAP7_75t_L g502 ( 
.A(n_405),
.Y(n_502)
);

INVx2_ASAP7_75t_L g503 ( 
.A(n_394),
.Y(n_503)
);

INVx1_ASAP7_75t_L g504 ( 
.A(n_427),
.Y(n_504)
);

NOR2xp33_ASAP7_75t_SL g505 ( 
.A(n_396),
.B(n_308),
.Y(n_505)
);

AND2x2_ASAP7_75t_L g506 ( 
.A(n_426),
.B(n_425),
.Y(n_506)
);

INVx1_ASAP7_75t_L g507 ( 
.A(n_427),
.Y(n_507)
);

OAI22xp33_ASAP7_75t_L g508 ( 
.A1(n_428),
.A2(n_354),
.B1(n_245),
.B2(n_227),
.Y(n_508)
);

INVx1_ASAP7_75t_L g509 ( 
.A(n_429),
.Y(n_509)
);

NAND2xp5_ASAP7_75t_L g510 ( 
.A(n_408),
.B(n_377),
.Y(n_510)
);

NAND2xp5_ASAP7_75t_SL g511 ( 
.A(n_391),
.B(n_381),
.Y(n_511)
);

NAND2xp5_ASAP7_75t_SL g512 ( 
.A(n_391),
.B(n_383),
.Y(n_512)
);

AND2x4_ASAP7_75t_L g513 ( 
.A(n_432),
.B(n_386),
.Y(n_513)
);

INVx2_ASAP7_75t_L g514 ( 
.A(n_395),
.Y(n_514)
);

INVx2_ASAP7_75t_L g515 ( 
.A(n_395),
.Y(n_515)
);

INVx2_ASAP7_75t_SL g516 ( 
.A(n_443),
.Y(n_516)
);

INVx1_ASAP7_75t_L g517 ( 
.A(n_429),
.Y(n_517)
);

OAI21xp5_ASAP7_75t_L g518 ( 
.A1(n_408),
.A2(n_382),
.B(n_215),
.Y(n_518)
);

INVx1_ASAP7_75t_L g519 ( 
.A(n_414),
.Y(n_519)
);

NOR2xp33_ASAP7_75t_L g520 ( 
.A(n_390),
.B(n_343),
.Y(n_520)
);

INVx1_ASAP7_75t_L g521 ( 
.A(n_414),
.Y(n_521)
);

INVx1_ASAP7_75t_L g522 ( 
.A(n_414),
.Y(n_522)
);

NAND2xp5_ASAP7_75t_L g523 ( 
.A(n_390),
.B(n_235),
.Y(n_523)
);

INVx3_ASAP7_75t_L g524 ( 
.A(n_417),
.Y(n_524)
);

NAND2xp5_ASAP7_75t_L g525 ( 
.A(n_390),
.B(n_393),
.Y(n_525)
);

INVx1_ASAP7_75t_L g526 ( 
.A(n_421),
.Y(n_526)
);

INVx3_ASAP7_75t_L g527 ( 
.A(n_417),
.Y(n_527)
);

BUFx3_ASAP7_75t_L g528 ( 
.A(n_423),
.Y(n_528)
);

INVx1_ASAP7_75t_L g529 ( 
.A(n_421),
.Y(n_529)
);

OR2x6_ASAP7_75t_L g530 ( 
.A(n_428),
.B(n_206),
.Y(n_530)
);

INVx2_ASAP7_75t_L g531 ( 
.A(n_395),
.Y(n_531)
);

INVx4_ASAP7_75t_L g532 ( 
.A(n_417),
.Y(n_532)
);

AOI22xp5_ASAP7_75t_L g533 ( 
.A1(n_451),
.A2(n_255),
.B1(n_174),
.B2(n_172),
.Y(n_533)
);

NAND2xp5_ASAP7_75t_SL g534 ( 
.A(n_451),
.B(n_164),
.Y(n_534)
);

INVx2_ASAP7_75t_L g535 ( 
.A(n_395),
.Y(n_535)
);

INVx1_ASAP7_75t_SL g536 ( 
.A(n_384),
.Y(n_536)
);

INVx2_ASAP7_75t_L g537 ( 
.A(n_397),
.Y(n_537)
);

INVx1_ASAP7_75t_L g538 ( 
.A(n_421),
.Y(n_538)
);

OR2x6_ASAP7_75t_L g539 ( 
.A(n_428),
.B(n_224),
.Y(n_539)
);

NOR2xp33_ASAP7_75t_L g540 ( 
.A(n_442),
.B(n_353),
.Y(n_540)
);

INVx2_ASAP7_75t_L g541 ( 
.A(n_397),
.Y(n_541)
);

INVx2_ASAP7_75t_L g542 ( 
.A(n_397),
.Y(n_542)
);

NAND2xp5_ASAP7_75t_SL g543 ( 
.A(n_446),
.B(n_167),
.Y(n_543)
);

INVx5_ASAP7_75t_L g544 ( 
.A(n_417),
.Y(n_544)
);

INVxp33_ASAP7_75t_SL g545 ( 
.A(n_449),
.Y(n_545)
);

OR2x2_ASAP7_75t_L g546 ( 
.A(n_393),
.B(n_359),
.Y(n_546)
);

INVx5_ASAP7_75t_L g547 ( 
.A(n_417),
.Y(n_547)
);

INVx2_ASAP7_75t_L g548 ( 
.A(n_397),
.Y(n_548)
);

NAND2xp5_ASAP7_75t_L g549 ( 
.A(n_406),
.B(n_412),
.Y(n_549)
);

INVx2_ASAP7_75t_SL g550 ( 
.A(n_386),
.Y(n_550)
);

INVx1_ASAP7_75t_L g551 ( 
.A(n_419),
.Y(n_551)
);

INVx3_ASAP7_75t_L g552 ( 
.A(n_420),
.Y(n_552)
);

AOI22xp5_ASAP7_75t_L g553 ( 
.A1(n_428),
.A2(n_248),
.B1(n_228),
.B2(n_168),
.Y(n_553)
);

INVx2_ASAP7_75t_L g554 ( 
.A(n_401),
.Y(n_554)
);

INVx1_ASAP7_75t_L g555 ( 
.A(n_419),
.Y(n_555)
);

OR2x2_ASAP7_75t_L g556 ( 
.A(n_406),
.B(n_360),
.Y(n_556)
);

CKINVDCx20_ASAP7_75t_R g557 ( 
.A(n_384),
.Y(n_557)
);

INVx2_ASAP7_75t_SL g558 ( 
.A(n_386),
.Y(n_558)
);

NAND2xp5_ASAP7_75t_L g559 ( 
.A(n_412),
.B(n_260),
.Y(n_559)
);

NAND2xp5_ASAP7_75t_SL g560 ( 
.A(n_446),
.B(n_167),
.Y(n_560)
);

INVx2_ASAP7_75t_L g561 ( 
.A(n_401),
.Y(n_561)
);

INVx2_ASAP7_75t_L g562 ( 
.A(n_401),
.Y(n_562)
);

INVxp67_ASAP7_75t_SL g563 ( 
.A(n_419),
.Y(n_563)
);

AND2x4_ASAP7_75t_L g564 ( 
.A(n_432),
.B(n_386),
.Y(n_564)
);

AND2x4_ASAP7_75t_L g565 ( 
.A(n_432),
.B(n_241),
.Y(n_565)
);

AOI21x1_ASAP7_75t_L g566 ( 
.A1(n_423),
.A2(n_274),
.B(n_265),
.Y(n_566)
);

INVx5_ASAP7_75t_L g567 ( 
.A(n_420),
.Y(n_567)
);

BUFx6f_ASAP7_75t_L g568 ( 
.A(n_420),
.Y(n_568)
);

INVx1_ASAP7_75t_L g569 ( 
.A(n_419),
.Y(n_569)
);

NAND2xp5_ASAP7_75t_L g570 ( 
.A(n_413),
.B(n_445),
.Y(n_570)
);

INVx3_ASAP7_75t_L g571 ( 
.A(n_420),
.Y(n_571)
);

NOR2xp33_ASAP7_75t_L g572 ( 
.A(n_449),
.B(n_357),
.Y(n_572)
);

INVx1_ASAP7_75t_L g573 ( 
.A(n_419),
.Y(n_573)
);

BUFx3_ASAP7_75t_L g574 ( 
.A(n_423),
.Y(n_574)
);

INVx1_ASAP7_75t_L g575 ( 
.A(n_401),
.Y(n_575)
);

AND2x2_ASAP7_75t_L g576 ( 
.A(n_415),
.B(n_360),
.Y(n_576)
);

NAND2xp5_ASAP7_75t_SL g577 ( 
.A(n_446),
.B(n_176),
.Y(n_577)
);

OR2x2_ASAP7_75t_L g578 ( 
.A(n_413),
.B(n_361),
.Y(n_578)
);

NAND2xp5_ASAP7_75t_SL g579 ( 
.A(n_446),
.B(n_449),
.Y(n_579)
);

INVx2_ASAP7_75t_L g580 ( 
.A(n_402),
.Y(n_580)
);

INVx1_ASAP7_75t_L g581 ( 
.A(n_402),
.Y(n_581)
);

INVx2_ASAP7_75t_SL g582 ( 
.A(n_386),
.Y(n_582)
);

AOI22xp33_ASAP7_75t_L g583 ( 
.A1(n_386),
.A2(n_236),
.B1(n_257),
.B2(n_273),
.Y(n_583)
);

INVxp33_ASAP7_75t_SL g584 ( 
.A(n_450),
.Y(n_584)
);

AOI22xp33_ASAP7_75t_L g585 ( 
.A1(n_422),
.A2(n_236),
.B1(n_257),
.B2(n_273),
.Y(n_585)
);

INVx2_ASAP7_75t_SL g586 ( 
.A(n_422),
.Y(n_586)
);

INVx3_ASAP7_75t_L g587 ( 
.A(n_420),
.Y(n_587)
);

NAND2xp5_ASAP7_75t_SL g588 ( 
.A(n_446),
.B(n_176),
.Y(n_588)
);

INVx1_ASAP7_75t_L g589 ( 
.A(n_402),
.Y(n_589)
);

OR2x2_ASAP7_75t_L g590 ( 
.A(n_450),
.B(n_361),
.Y(n_590)
);

NOR2xp33_ASAP7_75t_L g591 ( 
.A(n_415),
.B(n_362),
.Y(n_591)
);

INVx5_ASAP7_75t_L g592 ( 
.A(n_420),
.Y(n_592)
);

NAND2xp5_ASAP7_75t_L g593 ( 
.A(n_445),
.B(n_261),
.Y(n_593)
);

OAI21xp33_ASAP7_75t_SL g594 ( 
.A1(n_428),
.A2(n_363),
.B(n_370),
.Y(n_594)
);

NAND2xp5_ASAP7_75t_L g595 ( 
.A(n_445),
.B(n_262),
.Y(n_595)
);

BUFx10_ASAP7_75t_L g596 ( 
.A(n_432),
.Y(n_596)
);

INVx1_ASAP7_75t_L g597 ( 
.A(n_402),
.Y(n_597)
);

INVx1_ASAP7_75t_SL g598 ( 
.A(n_428),
.Y(n_598)
);

BUFx2_ASAP7_75t_L g599 ( 
.A(n_446),
.Y(n_599)
);

NAND2xp5_ASAP7_75t_SL g600 ( 
.A(n_396),
.B(n_180),
.Y(n_600)
);

INVx2_ASAP7_75t_L g601 ( 
.A(n_403),
.Y(n_601)
);

O2A1O1Ixp33_ASAP7_75t_L g602 ( 
.A1(n_525),
.A2(n_441),
.B(n_410),
.C(n_399),
.Y(n_602)
);

NAND2xp5_ASAP7_75t_SL g603 ( 
.A(n_467),
.B(n_432),
.Y(n_603)
);

NOR2xp33_ASAP7_75t_L g604 ( 
.A(n_584),
.B(n_399),
.Y(n_604)
);

AND2x4_ASAP7_75t_L g605 ( 
.A(n_460),
.B(n_410),
.Y(n_605)
);

INVxp67_ASAP7_75t_L g606 ( 
.A(n_540),
.Y(n_606)
);

NAND2xp5_ASAP7_75t_L g607 ( 
.A(n_549),
.B(n_422),
.Y(n_607)
);

NAND2xp5_ASAP7_75t_SL g608 ( 
.A(n_467),
.B(n_422),
.Y(n_608)
);

OAI22xp33_ASAP7_75t_L g609 ( 
.A1(n_546),
.A2(n_292),
.B1(n_301),
.B2(n_302),
.Y(n_609)
);

INVxp67_ASAP7_75t_L g610 ( 
.A(n_572),
.Y(n_610)
);

INVx4_ASAP7_75t_L g611 ( 
.A(n_513),
.Y(n_611)
);

CKINVDCx16_ASAP7_75t_R g612 ( 
.A(n_462),
.Y(n_612)
);

NOR2xp33_ASAP7_75t_L g613 ( 
.A(n_584),
.B(n_180),
.Y(n_613)
);

OR2x2_ASAP7_75t_L g614 ( 
.A(n_536),
.B(n_433),
.Y(n_614)
);

NAND2xp5_ASAP7_75t_SL g615 ( 
.A(n_467),
.B(n_422),
.Y(n_615)
);

NAND2xp5_ASAP7_75t_SL g616 ( 
.A(n_513),
.B(n_422),
.Y(n_616)
);

NAND2xp5_ASAP7_75t_L g617 ( 
.A(n_459),
.B(n_445),
.Y(n_617)
);

NAND2xp5_ASAP7_75t_L g618 ( 
.A(n_482),
.B(n_457),
.Y(n_618)
);

NAND2xp5_ASAP7_75t_L g619 ( 
.A(n_457),
.B(n_445),
.Y(n_619)
);

NAND2xp5_ASAP7_75t_SL g620 ( 
.A(n_513),
.B(n_445),
.Y(n_620)
);

INVx1_ASAP7_75t_L g621 ( 
.A(n_460),
.Y(n_621)
);

INVxp67_ASAP7_75t_L g622 ( 
.A(n_493),
.Y(n_622)
);

NAND2xp5_ASAP7_75t_L g623 ( 
.A(n_457),
.B(n_441),
.Y(n_623)
);

NAND2xp5_ASAP7_75t_L g624 ( 
.A(n_550),
.B(n_423),
.Y(n_624)
);

INVx2_ASAP7_75t_L g625 ( 
.A(n_454),
.Y(n_625)
);

AOI22xp5_ASAP7_75t_L g626 ( 
.A1(n_455),
.A2(n_423),
.B1(n_424),
.B2(n_266),
.Y(n_626)
);

INVx1_ASAP7_75t_SL g627 ( 
.A(n_557),
.Y(n_627)
);

NAND2xp5_ASAP7_75t_SL g628 ( 
.A(n_513),
.B(n_564),
.Y(n_628)
);

NAND2xp5_ASAP7_75t_SL g629 ( 
.A(n_564),
.B(n_596),
.Y(n_629)
);

INVxp67_ASAP7_75t_L g630 ( 
.A(n_493),
.Y(n_630)
);

BUFx6f_ASAP7_75t_SL g631 ( 
.A(n_488),
.Y(n_631)
);

INVx2_ASAP7_75t_L g632 ( 
.A(n_519),
.Y(n_632)
);

INVx2_ASAP7_75t_L g633 ( 
.A(n_519),
.Y(n_633)
);

INVx2_ASAP7_75t_L g634 ( 
.A(n_521),
.Y(n_634)
);

INVxp67_ASAP7_75t_L g635 ( 
.A(n_520),
.Y(n_635)
);

INVx1_ASAP7_75t_L g636 ( 
.A(n_528),
.Y(n_636)
);

INVxp67_ASAP7_75t_L g637 ( 
.A(n_591),
.Y(n_637)
);

INVx1_ASAP7_75t_L g638 ( 
.A(n_528),
.Y(n_638)
);

NAND2xp5_ASAP7_75t_L g639 ( 
.A(n_550),
.B(n_423),
.Y(n_639)
);

AOI22xp33_ASAP7_75t_L g640 ( 
.A1(n_494),
.A2(n_424),
.B1(n_448),
.B2(n_452),
.Y(n_640)
);

OAI22xp5_ASAP7_75t_L g641 ( 
.A1(n_461),
.A2(n_424),
.B1(n_181),
.B2(n_295),
.Y(n_641)
);

NAND2xp33_ASAP7_75t_L g642 ( 
.A(n_453),
.B(n_276),
.Y(n_642)
);

NOR2xp33_ASAP7_75t_L g643 ( 
.A(n_472),
.B(n_181),
.Y(n_643)
);

BUFx6f_ASAP7_75t_L g644 ( 
.A(n_574),
.Y(n_644)
);

AO22x2_ASAP7_75t_L g645 ( 
.A1(n_579),
.A2(n_363),
.B1(n_365),
.B2(n_366),
.Y(n_645)
);

NAND2xp5_ASAP7_75t_L g646 ( 
.A(n_558),
.B(n_424),
.Y(n_646)
);

INVx2_ASAP7_75t_L g647 ( 
.A(n_521),
.Y(n_647)
);

INVx1_ASAP7_75t_L g648 ( 
.A(n_574),
.Y(n_648)
);

INVx8_ASAP7_75t_L g649 ( 
.A(n_488),
.Y(n_649)
);

NAND2xp5_ASAP7_75t_L g650 ( 
.A(n_558),
.B(n_424),
.Y(n_650)
);

AOI22xp33_ASAP7_75t_L g651 ( 
.A1(n_494),
.A2(n_424),
.B1(n_448),
.B2(n_452),
.Y(n_651)
);

NAND2xp5_ASAP7_75t_L g652 ( 
.A(n_582),
.B(n_420),
.Y(n_652)
);

OAI22xp33_ASAP7_75t_L g653 ( 
.A1(n_546),
.A2(n_433),
.B1(n_435),
.B2(n_437),
.Y(n_653)
);

NOR2xp33_ASAP7_75t_L g654 ( 
.A(n_481),
.B(n_483),
.Y(n_654)
);

NAND2xp5_ASAP7_75t_L g655 ( 
.A(n_582),
.B(n_420),
.Y(n_655)
);

NAND2xp5_ASAP7_75t_L g656 ( 
.A(n_586),
.B(n_430),
.Y(n_656)
);

AND2x6_ASAP7_75t_SL g657 ( 
.A(n_488),
.B(n_365),
.Y(n_657)
);

NAND2xp5_ASAP7_75t_L g658 ( 
.A(n_586),
.B(n_430),
.Y(n_658)
);

INVx2_ASAP7_75t_L g659 ( 
.A(n_522),
.Y(n_659)
);

AND2x2_ASAP7_75t_L g660 ( 
.A(n_576),
.B(n_518),
.Y(n_660)
);

NAND2xp5_ASAP7_75t_L g661 ( 
.A(n_506),
.B(n_430),
.Y(n_661)
);

NOR3xp33_ASAP7_75t_L g662 ( 
.A(n_468),
.B(n_435),
.C(n_437),
.Y(n_662)
);

INVx2_ASAP7_75t_SL g663 ( 
.A(n_590),
.Y(n_663)
);

A2O1A1Ixp33_ASAP7_75t_L g664 ( 
.A1(n_570),
.A2(n_407),
.B(n_409),
.C(n_416),
.Y(n_664)
);

NAND2xp5_ASAP7_75t_L g665 ( 
.A(n_506),
.B(n_430),
.Y(n_665)
);

OR2x6_ASAP7_75t_L g666 ( 
.A(n_488),
.B(n_366),
.Y(n_666)
);

INVx1_ASAP7_75t_L g667 ( 
.A(n_456),
.Y(n_667)
);

NAND2xp5_ASAP7_75t_L g668 ( 
.A(n_489),
.B(n_430),
.Y(n_668)
);

INVx1_ASAP7_75t_L g669 ( 
.A(n_456),
.Y(n_669)
);

INVx1_ASAP7_75t_L g670 ( 
.A(n_465),
.Y(n_670)
);

INVx1_ASAP7_75t_L g671 ( 
.A(n_465),
.Y(n_671)
);

NAND2xp5_ASAP7_75t_L g672 ( 
.A(n_500),
.B(n_430),
.Y(n_672)
);

O2A1O1Ixp5_ASAP7_75t_L g673 ( 
.A1(n_565),
.A2(n_403),
.B(n_407),
.C(n_409),
.Y(n_673)
);

OAI22xp33_ASAP7_75t_L g674 ( 
.A1(n_556),
.A2(n_439),
.B1(n_444),
.B2(n_156),
.Y(n_674)
);

NAND2xp5_ASAP7_75t_SL g675 ( 
.A(n_564),
.B(n_596),
.Y(n_675)
);

INVx1_ASAP7_75t_L g676 ( 
.A(n_466),
.Y(n_676)
);

INVx2_ASAP7_75t_SL g677 ( 
.A(n_590),
.Y(n_677)
);

NAND3xp33_ASAP7_75t_L g678 ( 
.A(n_476),
.B(n_219),
.C(n_187),
.Y(n_678)
);

INVx1_ASAP7_75t_L g679 ( 
.A(n_466),
.Y(n_679)
);

BUFx6f_ASAP7_75t_L g680 ( 
.A(n_564),
.Y(n_680)
);

NAND2xp5_ASAP7_75t_SL g681 ( 
.A(n_596),
.B(n_430),
.Y(n_681)
);

INVx1_ASAP7_75t_L g682 ( 
.A(n_473),
.Y(n_682)
);

NAND2x1_ASAP7_75t_L g683 ( 
.A(n_453),
.B(n_403),
.Y(n_683)
);

INVx2_ASAP7_75t_L g684 ( 
.A(n_522),
.Y(n_684)
);

BUFx6f_ASAP7_75t_L g685 ( 
.A(n_596),
.Y(n_685)
);

NAND2xp5_ASAP7_75t_L g686 ( 
.A(n_559),
.B(n_430),
.Y(n_686)
);

AND2x2_ASAP7_75t_L g687 ( 
.A(n_576),
.B(n_439),
.Y(n_687)
);

INVx1_ASAP7_75t_L g688 ( 
.A(n_473),
.Y(n_688)
);

NAND2xp5_ASAP7_75t_L g689 ( 
.A(n_475),
.B(n_431),
.Y(n_689)
);

NOR2xp33_ASAP7_75t_L g690 ( 
.A(n_486),
.B(n_182),
.Y(n_690)
);

AND2x2_ASAP7_75t_L g691 ( 
.A(n_556),
.B(n_444),
.Y(n_691)
);

INVx1_ASAP7_75t_L g692 ( 
.A(n_475),
.Y(n_692)
);

NAND2xp5_ASAP7_75t_L g693 ( 
.A(n_477),
.B(n_431),
.Y(n_693)
);

NAND2xp5_ASAP7_75t_SL g694 ( 
.A(n_490),
.B(n_431),
.Y(n_694)
);

INVx2_ASAP7_75t_L g695 ( 
.A(n_526),
.Y(n_695)
);

NAND3xp33_ASAP7_75t_L g696 ( 
.A(n_523),
.B(n_218),
.C(n_189),
.Y(n_696)
);

NAND2xp5_ASAP7_75t_L g697 ( 
.A(n_477),
.B(n_431),
.Y(n_697)
);

AOI22xp5_ASAP7_75t_L g698 ( 
.A1(n_598),
.A2(n_267),
.B1(n_269),
.B2(n_277),
.Y(n_698)
);

NAND2xp5_ASAP7_75t_SL g699 ( 
.A(n_490),
.B(n_431),
.Y(n_699)
);

NOR2xp33_ASAP7_75t_L g700 ( 
.A(n_510),
.B(n_182),
.Y(n_700)
);

NAND2xp5_ASAP7_75t_L g701 ( 
.A(n_497),
.B(n_431),
.Y(n_701)
);

INVx2_ASAP7_75t_L g702 ( 
.A(n_454),
.Y(n_702)
);

INVx2_ASAP7_75t_L g703 ( 
.A(n_526),
.Y(n_703)
);

INVx4_ASAP7_75t_L g704 ( 
.A(n_490),
.Y(n_704)
);

NOR2xp33_ASAP7_75t_L g705 ( 
.A(n_578),
.B(n_289),
.Y(n_705)
);

INVx2_ASAP7_75t_L g706 ( 
.A(n_464),
.Y(n_706)
);

NAND2xp5_ASAP7_75t_L g707 ( 
.A(n_497),
.B(n_431),
.Y(n_707)
);

NAND2xp5_ASAP7_75t_SL g708 ( 
.A(n_490),
.B(n_431),
.Y(n_708)
);

BUFx6f_ASAP7_75t_L g709 ( 
.A(n_516),
.Y(n_709)
);

INVx2_ASAP7_75t_L g710 ( 
.A(n_529),
.Y(n_710)
);

INVx8_ASAP7_75t_L g711 ( 
.A(n_488),
.Y(n_711)
);

NAND2xp5_ASAP7_75t_L g712 ( 
.A(n_502),
.B(n_504),
.Y(n_712)
);

BUFx6f_ASAP7_75t_L g713 ( 
.A(n_516),
.Y(n_713)
);

INVx2_ASAP7_75t_L g714 ( 
.A(n_529),
.Y(n_714)
);

NAND2xp5_ASAP7_75t_L g715 ( 
.A(n_502),
.B(n_403),
.Y(n_715)
);

INVx2_ASAP7_75t_L g716 ( 
.A(n_538),
.Y(n_716)
);

INVx1_ASAP7_75t_L g717 ( 
.A(n_504),
.Y(n_717)
);

NAND2xp5_ASAP7_75t_SL g718 ( 
.A(n_578),
.B(n_236),
.Y(n_718)
);

NAND2xp5_ASAP7_75t_L g719 ( 
.A(n_507),
.B(n_407),
.Y(n_719)
);

NOR2xp33_ASAP7_75t_SL g720 ( 
.A(n_545),
.B(n_289),
.Y(n_720)
);

NAND2xp5_ASAP7_75t_SL g721 ( 
.A(n_565),
.B(n_236),
.Y(n_721)
);

AND2x2_ASAP7_75t_L g722 ( 
.A(n_479),
.B(n_448),
.Y(n_722)
);

NAND2xp5_ASAP7_75t_SL g723 ( 
.A(n_565),
.B(n_257),
.Y(n_723)
);

OAI22xp5_ASAP7_75t_L g724 ( 
.A1(n_492),
.A2(n_296),
.B1(n_306),
.B2(n_305),
.Y(n_724)
);

NAND2xp5_ASAP7_75t_L g725 ( 
.A(n_507),
.B(n_407),
.Y(n_725)
);

NAND2xp5_ASAP7_75t_L g726 ( 
.A(n_509),
.B(n_409),
.Y(n_726)
);

NAND2xp5_ASAP7_75t_L g727 ( 
.A(n_509),
.B(n_409),
.Y(n_727)
);

AOI22xp5_ASAP7_75t_L g728 ( 
.A1(n_534),
.A2(n_280),
.B1(n_287),
.B2(n_288),
.Y(n_728)
);

AOI22xp33_ASAP7_75t_L g729 ( 
.A1(n_583),
.A2(n_452),
.B1(n_273),
.B2(n_257),
.Y(n_729)
);

XOR2x2_ASAP7_75t_L g730 ( 
.A(n_533),
.B(n_553),
.Y(n_730)
);

NOR2xp33_ASAP7_75t_L g731 ( 
.A(n_511),
.B(n_294),
.Y(n_731)
);

NAND2xp5_ASAP7_75t_L g732 ( 
.A(n_517),
.B(n_416),
.Y(n_732)
);

INVx2_ASAP7_75t_L g733 ( 
.A(n_538),
.Y(n_733)
);

INVx1_ASAP7_75t_L g734 ( 
.A(n_517),
.Y(n_734)
);

NAND2xp5_ASAP7_75t_SL g735 ( 
.A(n_565),
.B(n_257),
.Y(n_735)
);

AND2x6_ASAP7_75t_L g736 ( 
.A(n_551),
.B(n_273),
.Y(n_736)
);

NAND2xp5_ASAP7_75t_SL g737 ( 
.A(n_594),
.B(n_416),
.Y(n_737)
);

NAND2xp5_ASAP7_75t_L g738 ( 
.A(n_563),
.B(n_416),
.Y(n_738)
);

NOR2xp67_ASAP7_75t_L g739 ( 
.A(n_594),
.B(n_447),
.Y(n_739)
);

NAND2xp5_ASAP7_75t_L g740 ( 
.A(n_551),
.B(n_418),
.Y(n_740)
);

NAND2xp5_ASAP7_75t_L g741 ( 
.A(n_555),
.B(n_418),
.Y(n_741)
);

NAND2xp5_ASAP7_75t_SL g742 ( 
.A(n_496),
.B(n_418),
.Y(n_742)
);

INVx2_ASAP7_75t_L g743 ( 
.A(n_464),
.Y(n_743)
);

AND2x6_ASAP7_75t_SL g744 ( 
.A(n_530),
.B(n_369),
.Y(n_744)
);

INVx1_ASAP7_75t_L g745 ( 
.A(n_555),
.Y(n_745)
);

NAND2xp5_ASAP7_75t_L g746 ( 
.A(n_569),
.B(n_573),
.Y(n_746)
);

INVxp67_ASAP7_75t_SL g747 ( 
.A(n_487),
.Y(n_747)
);

OR2x6_ASAP7_75t_L g748 ( 
.A(n_530),
.B(n_369),
.Y(n_748)
);

HB1xp67_ASAP7_75t_L g749 ( 
.A(n_470),
.Y(n_749)
);

AOI22xp33_ASAP7_75t_L g750 ( 
.A1(n_585),
.A2(n_276),
.B1(n_418),
.B2(n_447),
.Y(n_750)
);

INVx1_ASAP7_75t_L g751 ( 
.A(n_569),
.Y(n_751)
);

NAND2xp5_ASAP7_75t_L g752 ( 
.A(n_573),
.B(n_385),
.Y(n_752)
);

INVx1_ASAP7_75t_L g753 ( 
.A(n_479),
.Y(n_753)
);

INVx2_ASAP7_75t_L g754 ( 
.A(n_537),
.Y(n_754)
);

INVx1_ASAP7_75t_L g755 ( 
.A(n_575),
.Y(n_755)
);

NOR2xp33_ASAP7_75t_L g756 ( 
.A(n_512),
.B(n_294),
.Y(n_756)
);

INVx2_ASAP7_75t_L g757 ( 
.A(n_495),
.Y(n_757)
);

INVx1_ASAP7_75t_L g758 ( 
.A(n_575),
.Y(n_758)
);

INVx1_ASAP7_75t_L g759 ( 
.A(n_581),
.Y(n_759)
);

OR2x2_ASAP7_75t_L g760 ( 
.A(n_463),
.B(n_470),
.Y(n_760)
);

NAND2xp5_ASAP7_75t_L g761 ( 
.A(n_593),
.B(n_595),
.Y(n_761)
);

AND2x2_ASAP7_75t_L g762 ( 
.A(n_533),
.B(n_370),
.Y(n_762)
);

NAND2xp5_ASAP7_75t_L g763 ( 
.A(n_496),
.B(n_385),
.Y(n_763)
);

INVx2_ASAP7_75t_L g764 ( 
.A(n_537),
.Y(n_764)
);

NAND2xp5_ASAP7_75t_L g765 ( 
.A(n_496),
.B(n_385),
.Y(n_765)
);

NAND2xp5_ASAP7_75t_L g766 ( 
.A(n_471),
.B(n_434),
.Y(n_766)
);

INVx1_ASAP7_75t_L g767 ( 
.A(n_581),
.Y(n_767)
);

INVx2_ASAP7_75t_L g768 ( 
.A(n_495),
.Y(n_768)
);

NAND2xp5_ASAP7_75t_SL g769 ( 
.A(n_508),
.B(n_276),
.Y(n_769)
);

OR2x2_ASAP7_75t_L g770 ( 
.A(n_600),
.B(n_371),
.Y(n_770)
);

NAND2xp5_ASAP7_75t_L g771 ( 
.A(n_471),
.B(n_434),
.Y(n_771)
);

INVx1_ASAP7_75t_L g772 ( 
.A(n_589),
.Y(n_772)
);

BUFx6f_ASAP7_75t_L g773 ( 
.A(n_487),
.Y(n_773)
);

HB1xp67_ASAP7_75t_L g774 ( 
.A(n_622),
.Y(n_774)
);

BUFx2_ASAP7_75t_L g775 ( 
.A(n_630),
.Y(n_775)
);

INVx2_ASAP7_75t_L g776 ( 
.A(n_632),
.Y(n_776)
);

AOI21xp5_ASAP7_75t_L g777 ( 
.A1(n_704),
.A2(n_480),
.B(n_458),
.Y(n_777)
);

INVx2_ASAP7_75t_SL g778 ( 
.A(n_614),
.Y(n_778)
);

NAND2xp5_ASAP7_75t_L g779 ( 
.A(n_654),
.B(n_545),
.Y(n_779)
);

AOI21xp5_ASAP7_75t_L g780 ( 
.A1(n_704),
.A2(n_480),
.B(n_458),
.Y(n_780)
);

NOR2xp33_ASAP7_75t_L g781 ( 
.A(n_637),
.B(n_553),
.Y(n_781)
);

NAND2xp5_ASAP7_75t_L g782 ( 
.A(n_654),
.B(n_530),
.Y(n_782)
);

AOI22xp5_ASAP7_75t_L g783 ( 
.A1(n_618),
.A2(n_539),
.B1(n_530),
.B2(n_469),
.Y(n_783)
);

O2A1O1Ixp33_ASAP7_75t_L g784 ( 
.A1(n_718),
.A2(n_588),
.B(n_560),
.C(n_543),
.Y(n_784)
);

AOI21xp5_ASAP7_75t_L g785 ( 
.A1(n_617),
.A2(n_480),
.B(n_458),
.Y(n_785)
);

NAND2xp5_ASAP7_75t_L g786 ( 
.A(n_660),
.B(n_607),
.Y(n_786)
);

AOI21xp5_ASAP7_75t_L g787 ( 
.A1(n_668),
.A2(n_532),
.B(n_499),
.Y(n_787)
);

NOR2xp33_ASAP7_75t_L g788 ( 
.A(n_635),
.B(n_505),
.Y(n_788)
);

O2A1O1Ixp5_ASAP7_75t_L g789 ( 
.A1(n_718),
.A2(n_577),
.B(n_566),
.C(n_524),
.Y(n_789)
);

INVx2_ASAP7_75t_L g790 ( 
.A(n_632),
.Y(n_790)
);

NAND2xp5_ASAP7_75t_SL g791 ( 
.A(n_680),
.B(n_599),
.Y(n_791)
);

O2A1O1Ixp33_ASAP7_75t_SL g792 ( 
.A1(n_769),
.A2(n_589),
.B(n_597),
.C(n_601),
.Y(n_792)
);

O2A1O1Ixp33_ASAP7_75t_L g793 ( 
.A1(n_663),
.A2(n_530),
.B(n_539),
.C(n_597),
.Y(n_793)
);

INVx2_ASAP7_75t_L g794 ( 
.A(n_633),
.Y(n_794)
);

INVx2_ASAP7_75t_L g795 ( 
.A(n_633),
.Y(n_795)
);

AOI21xp5_ASAP7_75t_L g796 ( 
.A1(n_672),
.A2(n_532),
.B(n_499),
.Y(n_796)
);

BUFx4f_ASAP7_75t_L g797 ( 
.A(n_649),
.Y(n_797)
);

NOR2xp33_ASAP7_75t_SL g798 ( 
.A(n_749),
.B(n_627),
.Y(n_798)
);

NAND2xp5_ASAP7_75t_L g799 ( 
.A(n_687),
.B(n_539),
.Y(n_799)
);

AOI22xp5_ASAP7_75t_L g800 ( 
.A1(n_619),
.A2(n_539),
.B1(n_474),
.B2(n_599),
.Y(n_800)
);

NAND2xp5_ASAP7_75t_L g801 ( 
.A(n_691),
.B(n_539),
.Y(n_801)
);

OAI21xp5_ASAP7_75t_L g802 ( 
.A1(n_673),
.A2(n_601),
.B(n_541),
.Y(n_802)
);

NAND2x1_ASAP7_75t_L g803 ( 
.A(n_685),
.B(n_471),
.Y(n_803)
);

AOI21x1_ASAP7_75t_L g804 ( 
.A1(n_742),
.A2(n_566),
.B(n_542),
.Y(n_804)
);

OAI22xp5_ASAP7_75t_L g805 ( 
.A1(n_623),
.A2(n_478),
.B1(n_587),
.B2(n_484),
.Y(n_805)
);

OAI21xp5_ASAP7_75t_L g806 ( 
.A1(n_603),
.A2(n_542),
.B(n_541),
.Y(n_806)
);

AOI21xp5_ASAP7_75t_L g807 ( 
.A1(n_616),
.A2(n_532),
.B(n_499),
.Y(n_807)
);

OAI22xp5_ASAP7_75t_L g808 ( 
.A1(n_603),
.A2(n_478),
.B1(n_587),
.B2(n_484),
.Y(n_808)
);

INVx2_ASAP7_75t_L g809 ( 
.A(n_634),
.Y(n_809)
);

BUFx4f_ASAP7_75t_L g810 ( 
.A(n_649),
.Y(n_810)
);

AOI21xp5_ASAP7_75t_L g811 ( 
.A1(n_616),
.A2(n_487),
.B(n_568),
.Y(n_811)
);

AOI21xp5_ASAP7_75t_L g812 ( 
.A1(n_620),
.A2(n_487),
.B(n_568),
.Y(n_812)
);

AOI21xp5_ASAP7_75t_L g813 ( 
.A1(n_620),
.A2(n_699),
.B(n_694),
.Y(n_813)
);

NAND2xp5_ASAP7_75t_L g814 ( 
.A(n_643),
.B(n_478),
.Y(n_814)
);

AOI21xp5_ASAP7_75t_L g815 ( 
.A1(n_694),
.A2(n_487),
.B(n_568),
.Y(n_815)
);

AOI21xp5_ASAP7_75t_L g816 ( 
.A1(n_699),
.A2(n_568),
.B(n_587),
.Y(n_816)
);

NOR2x1_ASAP7_75t_L g817 ( 
.A(n_604),
.B(n_484),
.Y(n_817)
);

NAND2xp5_ASAP7_75t_SL g818 ( 
.A(n_680),
.B(n_485),
.Y(n_818)
);

OR2x2_ASAP7_75t_L g819 ( 
.A(n_760),
.B(n_371),
.Y(n_819)
);

OAI22xp5_ASAP7_75t_L g820 ( 
.A1(n_608),
.A2(n_485),
.B1(n_498),
.B2(n_571),
.Y(n_820)
);

INVx2_ASAP7_75t_SL g821 ( 
.A(n_770),
.Y(n_821)
);

NOR2x1p5_ASAP7_75t_SL g822 ( 
.A(n_754),
.B(n_764),
.Y(n_822)
);

AOI21xp5_ASAP7_75t_L g823 ( 
.A1(n_708),
.A2(n_568),
.B(n_498),
.Y(n_823)
);

AOI21xp5_ASAP7_75t_L g824 ( 
.A1(n_708),
.A2(n_501),
.B(n_498),
.Y(n_824)
);

NAND2xp5_ASAP7_75t_L g825 ( 
.A(n_643),
.B(n_485),
.Y(n_825)
);

AND2x2_ASAP7_75t_L g826 ( 
.A(n_677),
.B(n_156),
.Y(n_826)
);

AND2x4_ASAP7_75t_L g827 ( 
.A(n_621),
.B(n_447),
.Y(n_827)
);

OAI21xp5_ASAP7_75t_L g828 ( 
.A1(n_661),
.A2(n_548),
.B(n_580),
.Y(n_828)
);

INVx2_ASAP7_75t_L g829 ( 
.A(n_634),
.Y(n_829)
);

INVx2_ASAP7_75t_L g830 ( 
.A(n_647),
.Y(n_830)
);

A2O1A1Ixp33_ASAP7_75t_L g831 ( 
.A1(n_705),
.A2(n_729),
.B(n_604),
.C(n_731),
.Y(n_831)
);

AOI22xp5_ASAP7_75t_L g832 ( 
.A1(n_628),
.A2(n_501),
.B1(n_524),
.B2(n_571),
.Y(n_832)
);

AOI21xp5_ASAP7_75t_L g833 ( 
.A1(n_608),
.A2(n_552),
.B(n_527),
.Y(n_833)
);

INVx1_ASAP7_75t_L g834 ( 
.A(n_647),
.Y(n_834)
);

AOI21xp5_ASAP7_75t_L g835 ( 
.A1(n_615),
.A2(n_552),
.B(n_527),
.Y(n_835)
);

OAI21xp5_ASAP7_75t_L g836 ( 
.A1(n_665),
.A2(n_548),
.B(n_580),
.Y(n_836)
);

AOI21xp5_ASAP7_75t_L g837 ( 
.A1(n_615),
.A2(n_552),
.B(n_571),
.Y(n_837)
);

INVx3_ASAP7_75t_L g838 ( 
.A(n_611),
.Y(n_838)
);

OAI21xp5_ASAP7_75t_L g839 ( 
.A1(n_664),
.A2(n_562),
.B(n_561),
.Y(n_839)
);

HB1xp67_ASAP7_75t_L g840 ( 
.A(n_605),
.Y(n_840)
);

AOI21xp5_ASAP7_75t_L g841 ( 
.A1(n_624),
.A2(n_524),
.B(n_527),
.Y(n_841)
);

INVx1_ASAP7_75t_L g842 ( 
.A(n_659),
.Y(n_842)
);

AOI21xp5_ASAP7_75t_L g843 ( 
.A1(n_639),
.A2(n_501),
.B(n_567),
.Y(n_843)
);

NOR2x1_ASAP7_75t_L g844 ( 
.A(n_696),
.B(n_554),
.Y(n_844)
);

A2O1A1Ixp33_ASAP7_75t_L g845 ( 
.A1(n_705),
.A2(n_179),
.B(n_168),
.C(n_166),
.Y(n_845)
);

INVx2_ASAP7_75t_L g846 ( 
.A(n_659),
.Y(n_846)
);

OAI22xp5_ASAP7_75t_L g847 ( 
.A1(n_626),
.A2(n_295),
.B1(n_299),
.B2(n_305),
.Y(n_847)
);

INVx2_ASAP7_75t_L g848 ( 
.A(n_684),
.Y(n_848)
);

BUFx6f_ASAP7_75t_L g849 ( 
.A(n_680),
.Y(n_849)
);

AOI21xp5_ASAP7_75t_L g850 ( 
.A1(n_646),
.A2(n_592),
.B(n_567),
.Y(n_850)
);

AOI21xp5_ASAP7_75t_L g851 ( 
.A1(n_650),
.A2(n_592),
.B(n_567),
.Y(n_851)
);

INVx2_ASAP7_75t_L g852 ( 
.A(n_684),
.Y(n_852)
);

O2A1O1Ixp5_ASAP7_75t_L g853 ( 
.A1(n_737),
.A2(n_769),
.B(n_742),
.C(n_712),
.Y(n_853)
);

NAND2xp5_ASAP7_75t_L g854 ( 
.A(n_722),
.B(n_554),
.Y(n_854)
);

HB1xp67_ASAP7_75t_L g855 ( 
.A(n_605),
.Y(n_855)
);

AOI21xp5_ASAP7_75t_L g856 ( 
.A1(n_681),
.A2(n_592),
.B(n_567),
.Y(n_856)
);

NAND2xp5_ASAP7_75t_L g857 ( 
.A(n_690),
.B(n_561),
.Y(n_857)
);

OAI21xp5_ASAP7_75t_L g858 ( 
.A1(n_737),
.A2(n_562),
.B(n_514),
.Y(n_858)
);

NOR2x1p5_ASAP7_75t_L g859 ( 
.A(n_762),
.B(n_162),
.Y(n_859)
);

INVx3_ASAP7_75t_L g860 ( 
.A(n_611),
.Y(n_860)
);

OAI21xp5_ASAP7_75t_L g861 ( 
.A1(n_761),
.A2(n_503),
.B(n_514),
.Y(n_861)
);

AOI21xp5_ASAP7_75t_L g862 ( 
.A1(n_681),
.A2(n_592),
.B(n_567),
.Y(n_862)
);

AOI21xp5_ASAP7_75t_L g863 ( 
.A1(n_686),
.A2(n_675),
.B(n_629),
.Y(n_863)
);

AOI21xp5_ASAP7_75t_L g864 ( 
.A1(n_629),
.A2(n_592),
.B(n_567),
.Y(n_864)
);

AOI21xp5_ASAP7_75t_L g865 ( 
.A1(n_675),
.A2(n_592),
.B(n_547),
.Y(n_865)
);

AOI21x1_ASAP7_75t_L g866 ( 
.A1(n_683),
.A2(n_503),
.B(n_535),
.Y(n_866)
);

NOR3xp33_ASAP7_75t_L g867 ( 
.A(n_606),
.B(n_296),
.C(n_297),
.Y(n_867)
);

NAND2xp5_ASAP7_75t_L g868 ( 
.A(n_690),
.B(n_515),
.Y(n_868)
);

NAND2xp5_ASAP7_75t_L g869 ( 
.A(n_700),
.B(n_515),
.Y(n_869)
);

CKINVDCx6p67_ASAP7_75t_R g870 ( 
.A(n_612),
.Y(n_870)
);

AOI21xp5_ASAP7_75t_L g871 ( 
.A1(n_652),
.A2(n_547),
.B(n_544),
.Y(n_871)
);

BUFx4f_ASAP7_75t_L g872 ( 
.A(n_649),
.Y(n_872)
);

INVx2_ASAP7_75t_L g873 ( 
.A(n_695),
.Y(n_873)
);

INVx1_ASAP7_75t_L g874 ( 
.A(n_695),
.Y(n_874)
);

AOI22xp5_ASAP7_75t_L g875 ( 
.A1(n_628),
.A2(n_303),
.B1(n_297),
.B2(n_298),
.Y(n_875)
);

O2A1O1Ixp33_ASAP7_75t_L g876 ( 
.A1(n_653),
.A2(n_535),
.B(n_531),
.C(n_434),
.Y(n_876)
);

AND2x2_ASAP7_75t_L g877 ( 
.A(n_613),
.B(n_162),
.Y(n_877)
);

NAND2xp5_ASAP7_75t_SL g878 ( 
.A(n_680),
.B(n_531),
.Y(n_878)
);

NAND2xp5_ASAP7_75t_L g879 ( 
.A(n_700),
.B(n_298),
.Y(n_879)
);

AOI22xp33_ASAP7_75t_L g880 ( 
.A1(n_730),
.A2(n_276),
.B1(n_166),
.B2(n_169),
.Y(n_880)
);

AOI22xp5_ASAP7_75t_L g881 ( 
.A1(n_636),
.A2(n_299),
.B1(n_303),
.B2(n_306),
.Y(n_881)
);

AOI21xp5_ASAP7_75t_L g882 ( 
.A1(n_655),
.A2(n_547),
.B(n_544),
.Y(n_882)
);

NOR2xp33_ASAP7_75t_L g883 ( 
.A(n_610),
.B(n_192),
.Y(n_883)
);

NOR2xp33_ASAP7_75t_L g884 ( 
.A(n_613),
.B(n_212),
.Y(n_884)
);

AOI21xp5_ASAP7_75t_L g885 ( 
.A1(n_656),
.A2(n_547),
.B(n_544),
.Y(n_885)
);

NAND2xp5_ASAP7_75t_L g886 ( 
.A(n_667),
.B(n_434),
.Y(n_886)
);

CKINVDCx10_ASAP7_75t_R g887 ( 
.A(n_631),
.Y(n_887)
);

A2O1A1Ixp33_ASAP7_75t_L g888 ( 
.A1(n_729),
.A2(n_165),
.B(n_169),
.C(n_179),
.Y(n_888)
);

OAI21xp5_ASAP7_75t_L g889 ( 
.A1(n_739),
.A2(n_547),
.B(n_544),
.Y(n_889)
);

NOR3xp33_ASAP7_75t_L g890 ( 
.A(n_731),
.B(n_268),
.C(n_264),
.Y(n_890)
);

NAND2xp5_ASAP7_75t_L g891 ( 
.A(n_669),
.B(n_436),
.Y(n_891)
);

BUFx6f_ASAP7_75t_L g892 ( 
.A(n_773),
.Y(n_892)
);

NAND2xp5_ASAP7_75t_L g893 ( 
.A(n_670),
.B(n_436),
.Y(n_893)
);

INVx1_ASAP7_75t_L g894 ( 
.A(n_703),
.Y(n_894)
);

AOI21xp5_ASAP7_75t_L g895 ( 
.A1(n_658),
.A2(n_547),
.B(n_544),
.Y(n_895)
);

A2O1A1Ixp33_ASAP7_75t_L g896 ( 
.A1(n_756),
.A2(n_165),
.B(n_291),
.C(n_304),
.Y(n_896)
);

INVx1_ASAP7_75t_L g897 ( 
.A(n_703),
.Y(n_897)
);

INVx1_ASAP7_75t_L g898 ( 
.A(n_710),
.Y(n_898)
);

NAND2xp5_ASAP7_75t_SL g899 ( 
.A(n_685),
.B(n_276),
.Y(n_899)
);

AOI21xp5_ASAP7_75t_L g900 ( 
.A1(n_763),
.A2(n_544),
.B(n_491),
.Y(n_900)
);

NAND2xp5_ASAP7_75t_SL g901 ( 
.A(n_685),
.B(n_276),
.Y(n_901)
);

AOI21xp5_ASAP7_75t_L g902 ( 
.A1(n_765),
.A2(n_491),
.B(n_438),
.Y(n_902)
);

INVx2_ASAP7_75t_L g903 ( 
.A(n_710),
.Y(n_903)
);

OAI21xp5_ASAP7_75t_L g904 ( 
.A1(n_746),
.A2(n_491),
.B(n_438),
.Y(n_904)
);

NAND2xp5_ASAP7_75t_L g905 ( 
.A(n_671),
.B(n_436),
.Y(n_905)
);

NAND2xp5_ASAP7_75t_L g906 ( 
.A(n_676),
.B(n_436),
.Y(n_906)
);

AOI22xp5_ASAP7_75t_L g907 ( 
.A1(n_638),
.A2(n_276),
.B1(n_438),
.B2(n_214),
.Y(n_907)
);

NOR2xp33_ASAP7_75t_L g908 ( 
.A(n_720),
.B(n_216),
.Y(n_908)
);

NAND2xp5_ASAP7_75t_L g909 ( 
.A(n_679),
.B(n_438),
.Y(n_909)
);

AOI21xp5_ASAP7_75t_L g910 ( 
.A1(n_747),
.A2(n_491),
.B(n_272),
.Y(n_910)
);

NAND2xp5_ASAP7_75t_L g911 ( 
.A(n_682),
.B(n_491),
.Y(n_911)
);

NAND2xp5_ASAP7_75t_L g912 ( 
.A(n_688),
.B(n_491),
.Y(n_912)
);

INVx4_ASAP7_75t_L g913 ( 
.A(n_644),
.Y(n_913)
);

INVx2_ASAP7_75t_L g914 ( 
.A(n_714),
.Y(n_914)
);

OAI21xp5_ASAP7_75t_L g915 ( 
.A1(n_740),
.A2(n_271),
.B(n_225),
.Y(n_915)
);

NAND2xp5_ASAP7_75t_L g916 ( 
.A(n_692),
.B(n_276),
.Y(n_916)
);

OAI22xp5_ASAP7_75t_L g917 ( 
.A1(n_640),
.A2(n_237),
.B1(n_220),
.B2(n_285),
.Y(n_917)
);

AOI21x1_ASAP7_75t_L g918 ( 
.A1(n_715),
.A2(n_143),
.B(n_77),
.Y(n_918)
);

OAI22xp5_ASAP7_75t_L g919 ( 
.A1(n_640),
.A2(n_242),
.B1(n_243),
.B2(n_284),
.Y(n_919)
);

OAI22xp5_ASAP7_75t_L g920 ( 
.A1(n_651),
.A2(n_278),
.B1(n_251),
.B2(n_283),
.Y(n_920)
);

O2A1O1Ixp33_ASAP7_75t_L g921 ( 
.A1(n_753),
.A2(n_304),
.B(n_291),
.C(n_282),
.Y(n_921)
);

NOR2xp67_ASAP7_75t_L g922 ( 
.A(n_756),
.B(n_104),
.Y(n_922)
);

A2O1A1Ixp33_ASAP7_75t_L g923 ( 
.A1(n_602),
.A2(n_281),
.B(n_263),
.C(n_256),
.Y(n_923)
);

CKINVDCx20_ASAP7_75t_R g924 ( 
.A(n_698),
.Y(n_924)
);

NAND2xp5_ASAP7_75t_L g925 ( 
.A(n_717),
.B(n_246),
.Y(n_925)
);

INVx4_ASAP7_75t_L g926 ( 
.A(n_644),
.Y(n_926)
);

AOI21xp5_ASAP7_75t_L g927 ( 
.A1(n_738),
.A2(n_140),
.B(n_126),
.Y(n_927)
);

BUFx3_ASAP7_75t_L g928 ( 
.A(n_644),
.Y(n_928)
);

BUFx3_ASAP7_75t_L g929 ( 
.A(n_644),
.Y(n_929)
);

OAI21xp33_ASAP7_75t_L g930 ( 
.A1(n_662),
.A2(n_12),
.B(n_15),
.Y(n_930)
);

AND2x2_ASAP7_75t_L g931 ( 
.A(n_734),
.B(n_651),
.Y(n_931)
);

INVx2_ASAP7_75t_L g932 ( 
.A(n_714),
.Y(n_932)
);

INVx2_ASAP7_75t_L g933 ( 
.A(n_716),
.Y(n_933)
);

INVx2_ASAP7_75t_L g934 ( 
.A(n_716),
.Y(n_934)
);

NAND2xp5_ASAP7_75t_SL g935 ( 
.A(n_685),
.B(n_115),
.Y(n_935)
);

O2A1O1Ixp33_ASAP7_75t_L g936 ( 
.A1(n_641),
.A2(n_12),
.B(n_15),
.C(n_18),
.Y(n_936)
);

BUFx2_ASAP7_75t_L g937 ( 
.A(n_645),
.Y(n_937)
);

AOI21xp5_ASAP7_75t_L g938 ( 
.A1(n_773),
.A2(n_96),
.B(n_90),
.Y(n_938)
);

NAND2xp5_ASAP7_75t_SL g939 ( 
.A(n_733),
.B(n_85),
.Y(n_939)
);

OAI21xp5_ASAP7_75t_L g940 ( 
.A1(n_741),
.A2(n_81),
.B(n_79),
.Y(n_940)
);

NAND2xp33_ASAP7_75t_L g941 ( 
.A(n_709),
.B(n_713),
.Y(n_941)
);

NAND2xp5_ASAP7_75t_L g942 ( 
.A(n_733),
.B(n_20),
.Y(n_942)
);

NAND2xp5_ASAP7_75t_L g943 ( 
.A(n_648),
.B(n_21),
.Y(n_943)
);

NOR2xp33_ASAP7_75t_L g944 ( 
.A(n_674),
.B(n_678),
.Y(n_944)
);

AND2x2_ASAP7_75t_SL g945 ( 
.A(n_750),
.B(n_709),
.Y(n_945)
);

BUFx6f_ASAP7_75t_L g946 ( 
.A(n_773),
.Y(n_946)
);

CKINVDCx10_ASAP7_75t_R g947 ( 
.A(n_631),
.Y(n_947)
);

OAI21xp5_ASAP7_75t_L g948 ( 
.A1(n_689),
.A2(n_78),
.B(n_66),
.Y(n_948)
);

NAND2xp5_ASAP7_75t_L g949 ( 
.A(n_745),
.B(n_751),
.Y(n_949)
);

NOR2xp33_ASAP7_75t_L g950 ( 
.A(n_609),
.B(n_21),
.Y(n_950)
);

NOR2xp33_ASAP7_75t_L g951 ( 
.A(n_728),
.B(n_23),
.Y(n_951)
);

AND2x2_ASAP7_75t_L g952 ( 
.A(n_666),
.B(n_24),
.Y(n_952)
);

AOI22xp5_ASAP7_75t_L g953 ( 
.A1(n_645),
.A2(n_27),
.B1(n_28),
.B2(n_29),
.Y(n_953)
);

NAND2xp5_ASAP7_75t_L g954 ( 
.A(n_709),
.B(n_27),
.Y(n_954)
);

OAI21xp5_ASAP7_75t_L g955 ( 
.A1(n_693),
.A2(n_30),
.B(n_31),
.Y(n_955)
);

OAI21xp5_ASAP7_75t_L g956 ( 
.A1(n_697),
.A2(n_31),
.B(n_34),
.Y(n_956)
);

AOI21xp5_ASAP7_75t_L g957 ( 
.A1(n_773),
.A2(n_36),
.B(n_37),
.Y(n_957)
);

NAND2xp5_ASAP7_75t_L g958 ( 
.A(n_709),
.B(n_36),
.Y(n_958)
);

CKINVDCx6p67_ASAP7_75t_R g959 ( 
.A(n_666),
.Y(n_959)
);

NAND2xp33_ASAP7_75t_L g960 ( 
.A(n_713),
.B(n_37),
.Y(n_960)
);

O2A1O1Ixp33_ASAP7_75t_L g961 ( 
.A1(n_721),
.A2(n_38),
.B(n_41),
.C(n_43),
.Y(n_961)
);

AND2x2_ASAP7_75t_SL g962 ( 
.A(n_750),
.B(n_43),
.Y(n_962)
);

A2O1A1Ixp33_ASAP7_75t_L g963 ( 
.A1(n_711),
.A2(n_772),
.B(n_767),
.C(n_759),
.Y(n_963)
);

AOI21xp5_ASAP7_75t_L g964 ( 
.A1(n_642),
.A2(n_44),
.B(n_45),
.Y(n_964)
);

OAI22xp5_ASAP7_75t_L g965 ( 
.A1(n_831),
.A2(n_713),
.B1(n_645),
.B2(n_711),
.Y(n_965)
);

INVx3_ASAP7_75t_L g966 ( 
.A(n_849),
.Y(n_966)
);

NAND2xp5_ASAP7_75t_L g967 ( 
.A(n_779),
.B(n_713),
.Y(n_967)
);

NAND2xp5_ASAP7_75t_L g968 ( 
.A(n_884),
.B(n_732),
.Y(n_968)
);

NAND2xp5_ASAP7_75t_L g969 ( 
.A(n_884),
.B(n_719),
.Y(n_969)
);

NAND3xp33_ASAP7_75t_L g970 ( 
.A(n_908),
.B(n_724),
.C(n_666),
.Y(n_970)
);

OAI21xp5_ASAP7_75t_L g971 ( 
.A1(n_853),
.A2(n_727),
.B(n_725),
.Y(n_971)
);

O2A1O1Ixp33_ASAP7_75t_L g972 ( 
.A1(n_831),
.A2(n_723),
.B(n_721),
.C(n_735),
.Y(n_972)
);

NAND2x1p5_ASAP7_75t_L g973 ( 
.A(n_849),
.B(n_755),
.Y(n_973)
);

NAND2xp5_ASAP7_75t_L g974 ( 
.A(n_786),
.B(n_726),
.Y(n_974)
);

BUFx6f_ASAP7_75t_L g975 ( 
.A(n_892),
.Y(n_975)
);

NOR2xp67_ASAP7_75t_SL g976 ( 
.A(n_838),
.B(n_735),
.Y(n_976)
);

NAND3xp33_ASAP7_75t_SL g977 ( 
.A(n_890),
.B(n_723),
.C(n_701),
.Y(n_977)
);

OAI22xp5_ASAP7_75t_L g978 ( 
.A1(n_782),
.A2(n_711),
.B1(n_748),
.B2(n_758),
.Y(n_978)
);

NAND2xp5_ASAP7_75t_L g979 ( 
.A(n_931),
.B(n_752),
.Y(n_979)
);

NOR2xp33_ASAP7_75t_L g980 ( 
.A(n_788),
.B(n_657),
.Y(n_980)
);

NOR2xp33_ASAP7_75t_L g981 ( 
.A(n_788),
.B(n_744),
.Y(n_981)
);

OAI22xp5_ASAP7_75t_L g982 ( 
.A1(n_945),
.A2(n_748),
.B1(n_707),
.B2(n_764),
.Y(n_982)
);

NAND2xp5_ASAP7_75t_L g983 ( 
.A(n_877),
.B(n_754),
.Y(n_983)
);

NAND2xp5_ASAP7_75t_L g984 ( 
.A(n_879),
.B(n_743),
.Y(n_984)
);

BUFx2_ASAP7_75t_L g985 ( 
.A(n_775),
.Y(n_985)
);

HB1xp67_ASAP7_75t_L g986 ( 
.A(n_774),
.Y(n_986)
);

NAND2xp5_ASAP7_75t_L g987 ( 
.A(n_944),
.B(n_625),
.Y(n_987)
);

INVx2_ASAP7_75t_SL g988 ( 
.A(n_778),
.Y(n_988)
);

INVx3_ASAP7_75t_L g989 ( 
.A(n_849),
.Y(n_989)
);

AOI21xp5_ASAP7_75t_L g990 ( 
.A1(n_941),
.A2(n_785),
.B(n_863),
.Y(n_990)
);

O2A1O1Ixp33_ASAP7_75t_L g991 ( 
.A1(n_951),
.A2(n_748),
.B(n_766),
.C(n_771),
.Y(n_991)
);

NAND2xp5_ASAP7_75t_L g992 ( 
.A(n_944),
.B(n_768),
.Y(n_992)
);

O2A1O1Ixp5_ASAP7_75t_L g993 ( 
.A1(n_899),
.A2(n_757),
.B(n_706),
.C(n_702),
.Y(n_993)
);

AOI22xp33_ASAP7_75t_L g994 ( 
.A1(n_962),
.A2(n_736),
.B1(n_47),
.B2(n_48),
.Y(n_994)
);

AOI21xp5_ASAP7_75t_L g995 ( 
.A1(n_813),
.A2(n_736),
.B(n_48),
.Y(n_995)
);

NAND2xp5_ASAP7_75t_L g996 ( 
.A(n_883),
.B(n_736),
.Y(n_996)
);

NOR2xp33_ASAP7_75t_L g997 ( 
.A(n_781),
.B(n_46),
.Y(n_997)
);

INVx3_ASAP7_75t_L g998 ( 
.A(n_849),
.Y(n_998)
);

AOI21xp5_ASAP7_75t_L g999 ( 
.A1(n_787),
.A2(n_736),
.B(n_49),
.Y(n_999)
);

AOI22xp33_ASAP7_75t_SL g1000 ( 
.A1(n_781),
.A2(n_736),
.B1(n_51),
.B2(n_52),
.Y(n_1000)
);

NOR2xp33_ASAP7_75t_L g1001 ( 
.A(n_883),
.B(n_46),
.Y(n_1001)
);

INVx2_ASAP7_75t_L g1002 ( 
.A(n_790),
.Y(n_1002)
);

OAI22xp5_ASAP7_75t_L g1003 ( 
.A1(n_945),
.A2(n_51),
.B1(n_56),
.B2(n_58),
.Y(n_1003)
);

NOR2xp33_ASAP7_75t_L g1004 ( 
.A(n_821),
.B(n_56),
.Y(n_1004)
);

NAND2xp5_ASAP7_75t_L g1005 ( 
.A(n_801),
.B(n_59),
.Y(n_1005)
);

AOI21xp5_ASAP7_75t_L g1006 ( 
.A1(n_796),
.A2(n_60),
.B(n_61),
.Y(n_1006)
);

INVxp67_ASAP7_75t_L g1007 ( 
.A(n_774),
.Y(n_1007)
);

INVx2_ASAP7_75t_SL g1008 ( 
.A(n_819),
.Y(n_1008)
);

NAND2xp5_ASAP7_75t_L g1009 ( 
.A(n_827),
.B(n_60),
.Y(n_1009)
);

OAI21xp33_ASAP7_75t_SL g1010 ( 
.A1(n_962),
.A2(n_63),
.B(n_922),
.Y(n_1010)
);

INVx5_ASAP7_75t_L g1011 ( 
.A(n_892),
.Y(n_1011)
);

A2O1A1Ixp33_ASAP7_75t_L g1012 ( 
.A1(n_951),
.A2(n_784),
.B(n_908),
.C(n_783),
.Y(n_1012)
);

BUFx2_ASAP7_75t_L g1013 ( 
.A(n_840),
.Y(n_1013)
);

NAND2xp5_ASAP7_75t_SL g1014 ( 
.A(n_799),
.B(n_800),
.Y(n_1014)
);

INVx2_ASAP7_75t_L g1015 ( 
.A(n_794),
.Y(n_1015)
);

A2O1A1Ixp33_ASAP7_75t_L g1016 ( 
.A1(n_793),
.A2(n_930),
.B(n_950),
.C(n_956),
.Y(n_1016)
);

INVx2_ASAP7_75t_L g1017 ( 
.A(n_794),
.Y(n_1017)
);

INVx3_ASAP7_75t_L g1018 ( 
.A(n_838),
.Y(n_1018)
);

AOI21xp5_ASAP7_75t_L g1019 ( 
.A1(n_807),
.A2(n_777),
.B(n_780),
.Y(n_1019)
);

AOI22xp33_ASAP7_75t_L g1020 ( 
.A1(n_955),
.A2(n_880),
.B1(n_950),
.B2(n_937),
.Y(n_1020)
);

AOI21xp5_ASAP7_75t_L g1021 ( 
.A1(n_889),
.A2(n_825),
.B(n_814),
.Y(n_1021)
);

INVx1_ASAP7_75t_L g1022 ( 
.A(n_809),
.Y(n_1022)
);

INVx1_ASAP7_75t_L g1023 ( 
.A(n_809),
.Y(n_1023)
);

INVxp67_ASAP7_75t_SL g1024 ( 
.A(n_892),
.Y(n_1024)
);

NAND2xp5_ASAP7_75t_SL g1025 ( 
.A(n_860),
.B(n_829),
.Y(n_1025)
);

INVx2_ASAP7_75t_SL g1026 ( 
.A(n_859),
.Y(n_1026)
);

AND2x2_ASAP7_75t_L g1027 ( 
.A(n_826),
.B(n_840),
.Y(n_1027)
);

NAND2xp5_ASAP7_75t_SL g1028 ( 
.A(n_860),
.B(n_830),
.Y(n_1028)
);

NAND2xp5_ASAP7_75t_SL g1029 ( 
.A(n_830),
.B(n_846),
.Y(n_1029)
);

NAND2xp5_ASAP7_75t_SL g1030 ( 
.A(n_846),
.B(n_848),
.Y(n_1030)
);

OAI21x1_ASAP7_75t_L g1031 ( 
.A1(n_804),
.A2(n_802),
.B(n_839),
.Y(n_1031)
);

NAND2xp5_ASAP7_75t_L g1032 ( 
.A(n_827),
.B(n_857),
.Y(n_1032)
);

NAND2x1p5_ASAP7_75t_L g1033 ( 
.A(n_913),
.B(n_926),
.Y(n_1033)
);

BUFx2_ASAP7_75t_L g1034 ( 
.A(n_855),
.Y(n_1034)
);

INVx2_ASAP7_75t_L g1035 ( 
.A(n_848),
.Y(n_1035)
);

INVx2_ASAP7_75t_L g1036 ( 
.A(n_873),
.Y(n_1036)
);

NAND2xp5_ASAP7_75t_L g1037 ( 
.A(n_854),
.B(n_868),
.Y(n_1037)
);

AO22x1_ASAP7_75t_L g1038 ( 
.A1(n_952),
.A2(n_867),
.B1(n_855),
.B2(n_948),
.Y(n_1038)
);

OAI21x1_ASAP7_75t_L g1039 ( 
.A1(n_858),
.A2(n_841),
.B(n_866),
.Y(n_1039)
);

AOI21xp5_ASAP7_75t_L g1040 ( 
.A1(n_904),
.A2(n_869),
.B(n_812),
.Y(n_1040)
);

INVx2_ASAP7_75t_L g1041 ( 
.A(n_873),
.Y(n_1041)
);

O2A1O1Ixp5_ASAP7_75t_L g1042 ( 
.A1(n_899),
.A2(n_901),
.B(n_923),
.C(n_791),
.Y(n_1042)
);

NOR2xp33_ASAP7_75t_L g1043 ( 
.A(n_798),
.B(n_924),
.Y(n_1043)
);

O2A1O1Ixp33_ASAP7_75t_L g1044 ( 
.A1(n_896),
.A2(n_845),
.B(n_936),
.C(n_923),
.Y(n_1044)
);

INVx1_ASAP7_75t_L g1045 ( 
.A(n_903),
.Y(n_1045)
);

INVx3_ASAP7_75t_SL g1046 ( 
.A(n_870),
.Y(n_1046)
);

NOR2xp33_ASAP7_75t_R g1047 ( 
.A(n_797),
.B(n_810),
.Y(n_1047)
);

NAND2xp5_ASAP7_75t_L g1048 ( 
.A(n_817),
.B(n_903),
.Y(n_1048)
);

INVx2_ASAP7_75t_L g1049 ( 
.A(n_932),
.Y(n_1049)
);

AOI21xp5_ASAP7_75t_L g1050 ( 
.A1(n_811),
.A2(n_861),
.B(n_833),
.Y(n_1050)
);

O2A1O1Ixp33_ASAP7_75t_L g1051 ( 
.A1(n_896),
.A2(n_845),
.B(n_943),
.C(n_921),
.Y(n_1051)
);

A2O1A1Ixp33_ASAP7_75t_L g1052 ( 
.A1(n_953),
.A2(n_880),
.B(n_940),
.C(n_961),
.Y(n_1052)
);

HB1xp67_ASAP7_75t_L g1053 ( 
.A(n_954),
.Y(n_1053)
);

NOR2xp33_ASAP7_75t_L g1054 ( 
.A(n_925),
.B(n_949),
.Y(n_1054)
);

NAND2xp5_ASAP7_75t_L g1055 ( 
.A(n_932),
.B(n_934),
.Y(n_1055)
);

NAND2xp5_ASAP7_75t_SL g1056 ( 
.A(n_934),
.B(n_795),
.Y(n_1056)
);

A2O1A1Ixp33_ASAP7_75t_SL g1057 ( 
.A1(n_828),
.A2(n_836),
.B(n_942),
.C(n_958),
.Y(n_1057)
);

INVxp67_ASAP7_75t_L g1058 ( 
.A(n_917),
.Y(n_1058)
);

INVx1_ASAP7_75t_L g1059 ( 
.A(n_834),
.Y(n_1059)
);

BUFx6f_ASAP7_75t_L g1060 ( 
.A(n_892),
.Y(n_1060)
);

NAND2xp5_ASAP7_75t_L g1061 ( 
.A(n_842),
.B(n_874),
.Y(n_1061)
);

NAND2xp5_ASAP7_75t_SL g1062 ( 
.A(n_852),
.B(n_914),
.Y(n_1062)
);

BUFx12f_ASAP7_75t_L g1063 ( 
.A(n_913),
.Y(n_1063)
);

AOI22xp5_ASAP7_75t_L g1064 ( 
.A1(n_844),
.A2(n_960),
.B1(n_935),
.B2(n_791),
.Y(n_1064)
);

OAI22xp5_ASAP7_75t_SL g1065 ( 
.A1(n_919),
.A2(n_920),
.B1(n_875),
.B2(n_887),
.Y(n_1065)
);

NAND2xp5_ASAP7_75t_L g1066 ( 
.A(n_894),
.B(n_897),
.Y(n_1066)
);

CKINVDCx20_ASAP7_75t_R g1067 ( 
.A(n_959),
.Y(n_1067)
);

INVx2_ASAP7_75t_L g1068 ( 
.A(n_933),
.Y(n_1068)
);

NAND2xp5_ASAP7_75t_L g1069 ( 
.A(n_898),
.B(n_915),
.Y(n_1069)
);

HB1xp67_ASAP7_75t_L g1070 ( 
.A(n_928),
.Y(n_1070)
);

O2A1O1Ixp33_ASAP7_75t_SL g1071 ( 
.A1(n_963),
.A2(n_939),
.B(n_888),
.C(n_935),
.Y(n_1071)
);

NOR2xp33_ASAP7_75t_L g1072 ( 
.A(n_881),
.B(n_847),
.Y(n_1072)
);

AOI21xp5_ASAP7_75t_L g1073 ( 
.A1(n_835),
.A2(n_837),
.B(n_815),
.Y(n_1073)
);

OR2x2_ASAP7_75t_L g1074 ( 
.A(n_916),
.B(n_928),
.Y(n_1074)
);

INVx1_ASAP7_75t_L g1075 ( 
.A(n_886),
.Y(n_1075)
);

INVx4_ASAP7_75t_L g1076 ( 
.A(n_946),
.Y(n_1076)
);

NAND2xp5_ASAP7_75t_L g1077 ( 
.A(n_888),
.B(n_929),
.Y(n_1077)
);

AOI21xp5_ASAP7_75t_L g1078 ( 
.A1(n_818),
.A2(n_820),
.B(n_808),
.Y(n_1078)
);

AOI21xp5_ASAP7_75t_L g1079 ( 
.A1(n_818),
.A2(n_806),
.B(n_823),
.Y(n_1079)
);

NAND2xp5_ASAP7_75t_L g1080 ( 
.A(n_929),
.B(n_926),
.Y(n_1080)
);

INVx3_ASAP7_75t_L g1081 ( 
.A(n_946),
.Y(n_1081)
);

A2O1A1Ixp33_ASAP7_75t_L g1082 ( 
.A1(n_964),
.A2(n_957),
.B(n_963),
.C(n_789),
.Y(n_1082)
);

NOR2x1_ASAP7_75t_L g1083 ( 
.A(n_939),
.B(n_901),
.Y(n_1083)
);

BUFx2_ASAP7_75t_L g1084 ( 
.A(n_946),
.Y(n_1084)
);

BUFx12f_ASAP7_75t_L g1085 ( 
.A(n_946),
.Y(n_1085)
);

HB1xp67_ASAP7_75t_L g1086 ( 
.A(n_797),
.Y(n_1086)
);

O2A1O1Ixp33_ASAP7_75t_L g1087 ( 
.A1(n_792),
.A2(n_805),
.B(n_905),
.C(n_909),
.Y(n_1087)
);

CKINVDCx5p33_ASAP7_75t_R g1088 ( 
.A(n_947),
.Y(n_1088)
);

NOR3xp33_ASAP7_75t_SL g1089 ( 
.A(n_938),
.B(n_927),
.C(n_878),
.Y(n_1089)
);

A2O1A1Ixp33_ASAP7_75t_L g1090 ( 
.A1(n_822),
.A2(n_907),
.B(n_876),
.C(n_810),
.Y(n_1090)
);

AOI22xp33_ASAP7_75t_L g1091 ( 
.A1(n_891),
.A2(n_906),
.B1(n_893),
.B2(n_878),
.Y(n_1091)
);

AND2x2_ASAP7_75t_L g1092 ( 
.A(n_872),
.B(n_832),
.Y(n_1092)
);

NOR2xp33_ASAP7_75t_L g1093 ( 
.A(n_872),
.B(n_912),
.Y(n_1093)
);

NOR2xp33_ASAP7_75t_L g1094 ( 
.A(n_911),
.B(n_792),
.Y(n_1094)
);

OAI22xp5_ASAP7_75t_L g1095 ( 
.A1(n_803),
.A2(n_824),
.B1(n_816),
.B2(n_843),
.Y(n_1095)
);

INVx3_ASAP7_75t_L g1096 ( 
.A(n_918),
.Y(n_1096)
);

OAI22xp33_ASAP7_75t_L g1097 ( 
.A1(n_910),
.A2(n_902),
.B1(n_864),
.B2(n_865),
.Y(n_1097)
);

AOI21xp5_ASAP7_75t_L g1098 ( 
.A1(n_850),
.A2(n_851),
.B(n_900),
.Y(n_1098)
);

INVx2_ASAP7_75t_L g1099 ( 
.A(n_871),
.Y(n_1099)
);

AND2x2_ASAP7_75t_L g1100 ( 
.A(n_856),
.B(n_862),
.Y(n_1100)
);

NAND2xp5_ASAP7_75t_SL g1101 ( 
.A(n_882),
.B(n_885),
.Y(n_1101)
);

AO21x1_ASAP7_75t_L g1102 ( 
.A1(n_895),
.A2(n_618),
.B(n_955),
.Y(n_1102)
);

AO32x2_ASAP7_75t_L g1103 ( 
.A1(n_805),
.A2(n_641),
.A3(n_808),
.B1(n_820),
.B2(n_677),
.Y(n_1103)
);

INVx1_ASAP7_75t_L g1104 ( 
.A(n_776),
.Y(n_1104)
);

OAI22xp5_ASAP7_75t_SL g1105 ( 
.A1(n_924),
.A2(n_462),
.B1(n_411),
.B2(n_781),
.Y(n_1105)
);

NAND2xp5_ASAP7_75t_L g1106 ( 
.A(n_779),
.B(n_654),
.Y(n_1106)
);

INVx3_ASAP7_75t_SL g1107 ( 
.A(n_870),
.Y(n_1107)
);

INVx2_ASAP7_75t_L g1108 ( 
.A(n_776),
.Y(n_1108)
);

NAND2xp5_ASAP7_75t_L g1109 ( 
.A(n_779),
.B(n_654),
.Y(n_1109)
);

AO21x1_ASAP7_75t_L g1110 ( 
.A1(n_1001),
.A2(n_1044),
.B(n_1014),
.Y(n_1110)
);

INVx1_ASAP7_75t_SL g1111 ( 
.A(n_985),
.Y(n_1111)
);

INVx1_ASAP7_75t_L g1112 ( 
.A(n_1059),
.Y(n_1112)
);

NOR2xp33_ASAP7_75t_SL g1113 ( 
.A(n_997),
.B(n_1001),
.Y(n_1113)
);

AO31x2_ASAP7_75t_L g1114 ( 
.A1(n_1102),
.A2(n_1082),
.A3(n_1012),
.B(n_965),
.Y(n_1114)
);

AO22x2_ASAP7_75t_L g1115 ( 
.A1(n_1003),
.A2(n_970),
.B1(n_1014),
.B2(n_978),
.Y(n_1115)
);

NAND3xp33_ASAP7_75t_L g1116 ( 
.A(n_997),
.B(n_1072),
.C(n_1106),
.Y(n_1116)
);

OAI21x1_ASAP7_75t_L g1117 ( 
.A1(n_1098),
.A2(n_1039),
.B(n_990),
.Y(n_1117)
);

OAI21xp5_ASAP7_75t_L g1118 ( 
.A1(n_1078),
.A2(n_1109),
.B(n_1052),
.Y(n_1118)
);

AO21x2_ASAP7_75t_L g1119 ( 
.A1(n_1050),
.A2(n_1082),
.B(n_1101),
.Y(n_1119)
);

OAI21x1_ASAP7_75t_L g1120 ( 
.A1(n_1073),
.A2(n_1079),
.B(n_1095),
.Y(n_1120)
);

AOI21xp5_ASAP7_75t_L g1121 ( 
.A1(n_1040),
.A2(n_974),
.B(n_968),
.Y(n_1121)
);

O2A1O1Ixp33_ASAP7_75t_SL g1122 ( 
.A1(n_1052),
.A2(n_1016),
.B(n_1090),
.C(n_969),
.Y(n_1122)
);

NAND2xp5_ASAP7_75t_L g1123 ( 
.A(n_1054),
.B(n_979),
.Y(n_1123)
);

O2A1O1Ixp33_ASAP7_75t_SL g1124 ( 
.A1(n_1058),
.A2(n_1072),
.B(n_1077),
.C(n_996),
.Y(n_1124)
);

AOI21xp5_ASAP7_75t_L g1125 ( 
.A1(n_1057),
.A2(n_1037),
.B(n_971),
.Y(n_1125)
);

AOI21xp5_ASAP7_75t_L g1126 ( 
.A1(n_1057),
.A2(n_1069),
.B(n_972),
.Y(n_1126)
);

AOI21xp5_ASAP7_75t_L g1127 ( 
.A1(n_1054),
.A2(n_991),
.B(n_1087),
.Y(n_1127)
);

OAI21x1_ASAP7_75t_L g1128 ( 
.A1(n_1031),
.A2(n_993),
.B(n_1099),
.Y(n_1128)
);

NAND2xp5_ASAP7_75t_L g1129 ( 
.A(n_1032),
.B(n_1020),
.Y(n_1129)
);

AOI22xp33_ASAP7_75t_L g1130 ( 
.A1(n_1065),
.A2(n_1020),
.B1(n_980),
.B2(n_981),
.Y(n_1130)
);

OAI22xp33_ASAP7_75t_L g1131 ( 
.A1(n_1008),
.A2(n_981),
.B1(n_980),
.B2(n_1043),
.Y(n_1131)
);

AOI21xp5_ASAP7_75t_L g1132 ( 
.A1(n_987),
.A2(n_992),
.B(n_967),
.Y(n_1132)
);

BUFx2_ASAP7_75t_L g1133 ( 
.A(n_986),
.Y(n_1133)
);

OAI21xp5_ASAP7_75t_L g1134 ( 
.A1(n_1042),
.A2(n_1010),
.B(n_1094),
.Y(n_1134)
);

AOI21xp5_ASAP7_75t_L g1135 ( 
.A1(n_1097),
.A2(n_984),
.B(n_1071),
.Y(n_1135)
);

AOI21xp5_ASAP7_75t_L g1136 ( 
.A1(n_1071),
.A2(n_1099),
.B(n_1094),
.Y(n_1136)
);

AOI221xp5_ASAP7_75t_L g1137 ( 
.A1(n_1051),
.A2(n_994),
.B1(n_1004),
.B2(n_1105),
.C(n_1043),
.Y(n_1137)
);

AO31x2_ASAP7_75t_L g1138 ( 
.A1(n_982),
.A2(n_995),
.A3(n_999),
.B(n_1006),
.Y(n_1138)
);

AOI21xp5_ASAP7_75t_L g1139 ( 
.A1(n_1100),
.A2(n_1083),
.B(n_983),
.Y(n_1139)
);

AOI22xp5_ASAP7_75t_L g1140 ( 
.A1(n_1027),
.A2(n_1026),
.B1(n_1092),
.B2(n_1053),
.Y(n_1140)
);

NAND2xp5_ASAP7_75t_L g1141 ( 
.A(n_1075),
.B(n_1002),
.Y(n_1141)
);

BUFx2_ASAP7_75t_L g1142 ( 
.A(n_1013),
.Y(n_1142)
);

AOI221x1_ASAP7_75t_L g1143 ( 
.A1(n_1005),
.A2(n_977),
.B1(n_1096),
.B2(n_1093),
.C(n_1004),
.Y(n_1143)
);

OAI21x1_ASAP7_75t_L g1144 ( 
.A1(n_1096),
.A2(n_1048),
.B(n_1030),
.Y(n_1144)
);

NAND2xp5_ASAP7_75t_SL g1145 ( 
.A(n_1007),
.B(n_988),
.Y(n_1145)
);

NOR2xp67_ASAP7_75t_SL g1146 ( 
.A(n_1063),
.B(n_1011),
.Y(n_1146)
);

CKINVDCx20_ASAP7_75t_R g1147 ( 
.A(n_1046),
.Y(n_1147)
);

INVx4_ASAP7_75t_L g1148 ( 
.A(n_1085),
.Y(n_1148)
);

CKINVDCx11_ASAP7_75t_R g1149 ( 
.A(n_1046),
.Y(n_1149)
);

AO32x2_ASAP7_75t_L g1150 ( 
.A1(n_1076),
.A2(n_1103),
.A3(n_994),
.B1(n_1038),
.B2(n_1064),
.Y(n_1150)
);

AO31x2_ASAP7_75t_L g1151 ( 
.A1(n_1093),
.A2(n_1108),
.A3(n_1015),
.B(n_1049),
.Y(n_1151)
);

INVx2_ASAP7_75t_SL g1152 ( 
.A(n_1034),
.Y(n_1152)
);

OR2x2_ASAP7_75t_L g1153 ( 
.A(n_1009),
.B(n_1070),
.Y(n_1153)
);

A2O1A1Ixp33_ASAP7_75t_L g1154 ( 
.A1(n_1089),
.A2(n_1074),
.B(n_976),
.C(n_1066),
.Y(n_1154)
);

AOI21xp5_ASAP7_75t_L g1155 ( 
.A1(n_1025),
.A2(n_1028),
.B(n_1091),
.Y(n_1155)
);

OAI21x1_ASAP7_75t_L g1156 ( 
.A1(n_1029),
.A2(n_1030),
.B(n_1028),
.Y(n_1156)
);

BUFx2_ASAP7_75t_L g1157 ( 
.A(n_1084),
.Y(n_1157)
);

OAI21xp5_ASAP7_75t_L g1158 ( 
.A1(n_1091),
.A2(n_1029),
.B(n_1056),
.Y(n_1158)
);

AOI21xp33_ASAP7_75t_L g1159 ( 
.A1(n_1061),
.A2(n_1000),
.B(n_1045),
.Y(n_1159)
);

HB1xp67_ASAP7_75t_L g1160 ( 
.A(n_966),
.Y(n_1160)
);

BUFx12f_ASAP7_75t_L g1161 ( 
.A(n_1088),
.Y(n_1161)
);

OAI21x1_ASAP7_75t_L g1162 ( 
.A1(n_1025),
.A2(n_1055),
.B(n_1056),
.Y(n_1162)
);

O2A1O1Ixp33_ASAP7_75t_L g1163 ( 
.A1(n_1086),
.A2(n_1062),
.B(n_1068),
.C(n_1107),
.Y(n_1163)
);

AND2x2_ASAP7_75t_L g1164 ( 
.A(n_1068),
.B(n_1107),
.Y(n_1164)
);

O2A1O1Ixp5_ASAP7_75t_L g1165 ( 
.A1(n_1062),
.A2(n_1080),
.B(n_1018),
.C(n_1023),
.Y(n_1165)
);

OAI21x1_ASAP7_75t_L g1166 ( 
.A1(n_973),
.A2(n_1035),
.B(n_1049),
.Y(n_1166)
);

NAND2xp5_ASAP7_75t_L g1167 ( 
.A(n_1017),
.B(n_1035),
.Y(n_1167)
);

OAI21xp5_ASAP7_75t_L g1168 ( 
.A1(n_1017),
.A2(n_1041),
.B(n_1036),
.Y(n_1168)
);

AOI221xp5_ASAP7_75t_L g1169 ( 
.A1(n_1022),
.A2(n_1104),
.B1(n_1047),
.B2(n_1067),
.C(n_1036),
.Y(n_1169)
);

OR2x2_ASAP7_75t_L g1170 ( 
.A(n_966),
.B(n_989),
.Y(n_1170)
);

AND2x4_ASAP7_75t_L g1171 ( 
.A(n_989),
.B(n_998),
.Y(n_1171)
);

A2O1A1Ixp33_ASAP7_75t_L g1172 ( 
.A1(n_998),
.A2(n_1024),
.B(n_1081),
.C(n_1011),
.Y(n_1172)
);

AND2x4_ASAP7_75t_L g1173 ( 
.A(n_1011),
.B(n_1076),
.Y(n_1173)
);

INVx1_ASAP7_75t_L g1174 ( 
.A(n_1081),
.Y(n_1174)
);

AO31x2_ASAP7_75t_L g1175 ( 
.A1(n_1103),
.A2(n_1011),
.A3(n_975),
.B(n_1060),
.Y(n_1175)
);

OA21x2_ASAP7_75t_L g1176 ( 
.A1(n_1103),
.A2(n_975),
.B(n_1060),
.Y(n_1176)
);

AOI221x1_ASAP7_75t_L g1177 ( 
.A1(n_1103),
.A2(n_975),
.B1(n_1060),
.B2(n_1047),
.C(n_1033),
.Y(n_1177)
);

AO32x2_ASAP7_75t_L g1178 ( 
.A1(n_1060),
.A2(n_965),
.A3(n_1003),
.B1(n_978),
.B2(n_982),
.Y(n_1178)
);

OAI21x1_ASAP7_75t_L g1179 ( 
.A1(n_1019),
.A2(n_1098),
.B(n_1039),
.Y(n_1179)
);

NAND3xp33_ASAP7_75t_L g1180 ( 
.A(n_1001),
.B(n_884),
.C(n_1012),
.Y(n_1180)
);

AO31x2_ASAP7_75t_L g1181 ( 
.A1(n_1102),
.A2(n_1082),
.A3(n_1012),
.B(n_965),
.Y(n_1181)
);

NAND2xp5_ASAP7_75t_L g1182 ( 
.A(n_1106),
.B(n_1109),
.Y(n_1182)
);

INVx1_ASAP7_75t_L g1183 ( 
.A(n_1059),
.Y(n_1183)
);

A2O1A1Ixp33_ASAP7_75t_L g1184 ( 
.A1(n_1012),
.A2(n_831),
.B(n_1001),
.C(n_1072),
.Y(n_1184)
);

NOR2x1_ASAP7_75t_SL g1185 ( 
.A(n_1011),
.B(n_685),
.Y(n_1185)
);

INVx1_ASAP7_75t_L g1186 ( 
.A(n_1059),
.Y(n_1186)
);

NAND2xp5_ASAP7_75t_SL g1187 ( 
.A(n_1106),
.B(n_779),
.Y(n_1187)
);

AOI22xp33_ASAP7_75t_L g1188 ( 
.A1(n_997),
.A2(n_1072),
.B1(n_730),
.B2(n_1001),
.Y(n_1188)
);

NOR2xp33_ASAP7_75t_L g1189 ( 
.A(n_1106),
.B(n_637),
.Y(n_1189)
);

AND2x4_ASAP7_75t_L g1190 ( 
.A(n_1086),
.B(n_1027),
.Y(n_1190)
);

INVx2_ASAP7_75t_SL g1191 ( 
.A(n_985),
.Y(n_1191)
);

NAND2xp5_ASAP7_75t_L g1192 ( 
.A(n_1106),
.B(n_1109),
.Y(n_1192)
);

O2A1O1Ixp33_ASAP7_75t_L g1193 ( 
.A1(n_1001),
.A2(n_1012),
.B(n_997),
.C(n_884),
.Y(n_1193)
);

INVx5_ASAP7_75t_L g1194 ( 
.A(n_975),
.Y(n_1194)
);

OAI21xp5_ASAP7_75t_L g1195 ( 
.A1(n_1012),
.A2(n_831),
.B(n_618),
.Y(n_1195)
);

AND2x2_ASAP7_75t_L g1196 ( 
.A(n_1027),
.B(n_877),
.Y(n_1196)
);

OAI21x1_ASAP7_75t_L g1197 ( 
.A1(n_1019),
.A2(n_1098),
.B(n_1039),
.Y(n_1197)
);

OAI22xp5_ASAP7_75t_L g1198 ( 
.A1(n_1020),
.A2(n_994),
.B1(n_1109),
.B2(n_1106),
.Y(n_1198)
);

INVx1_ASAP7_75t_SL g1199 ( 
.A(n_985),
.Y(n_1199)
);

OAI22xp5_ASAP7_75t_L g1200 ( 
.A1(n_1020),
.A2(n_994),
.B1(n_1109),
.B2(n_1106),
.Y(n_1200)
);

O2A1O1Ixp33_ASAP7_75t_L g1201 ( 
.A1(n_1001),
.A2(n_1012),
.B(n_997),
.C(n_884),
.Y(n_1201)
);

AND2x4_ASAP7_75t_L g1202 ( 
.A(n_1086),
.B(n_1027),
.Y(n_1202)
);

AO32x1_ASAP7_75t_L g1203 ( 
.A1(n_1003),
.A2(n_965),
.A3(n_978),
.B1(n_1095),
.B2(n_982),
.Y(n_1203)
);

O2A1O1Ixp33_ASAP7_75t_SL g1204 ( 
.A1(n_1012),
.A2(n_831),
.B(n_1052),
.C(n_1016),
.Y(n_1204)
);

A2O1A1Ixp33_ASAP7_75t_L g1205 ( 
.A1(n_1012),
.A2(n_831),
.B(n_1001),
.C(n_1072),
.Y(n_1205)
);

O2A1O1Ixp33_ASAP7_75t_L g1206 ( 
.A1(n_1001),
.A2(n_1012),
.B(n_997),
.C(n_884),
.Y(n_1206)
);

NOR2xp33_ASAP7_75t_L g1207 ( 
.A(n_1106),
.B(n_637),
.Y(n_1207)
);

NOR2xp33_ASAP7_75t_L g1208 ( 
.A(n_1106),
.B(n_637),
.Y(n_1208)
);

AOI221xp5_ASAP7_75t_L g1209 ( 
.A1(n_997),
.A2(n_880),
.B1(n_781),
.B2(n_396),
.C(n_1001),
.Y(n_1209)
);

AND2x2_ASAP7_75t_L g1210 ( 
.A(n_1027),
.B(n_877),
.Y(n_1210)
);

OAI21x1_ASAP7_75t_L g1211 ( 
.A1(n_1019),
.A2(n_1098),
.B(n_1039),
.Y(n_1211)
);

INVx1_ASAP7_75t_L g1212 ( 
.A(n_1059),
.Y(n_1212)
);

AOI221x1_ASAP7_75t_L g1213 ( 
.A1(n_1012),
.A2(n_1052),
.B1(n_997),
.B2(n_1001),
.C(n_1016),
.Y(n_1213)
);

AOI21xp5_ASAP7_75t_L g1214 ( 
.A1(n_990),
.A2(n_704),
.B(n_941),
.Y(n_1214)
);

CKINVDCx5p33_ASAP7_75t_R g1215 ( 
.A(n_1088),
.Y(n_1215)
);

OAI21x1_ASAP7_75t_L g1216 ( 
.A1(n_1019),
.A2(n_1098),
.B(n_1039),
.Y(n_1216)
);

AOI31xp67_ASAP7_75t_L g1217 ( 
.A1(n_1101),
.A2(n_1099),
.A3(n_1014),
.B(n_1064),
.Y(n_1217)
);

OAI22xp5_ASAP7_75t_R g1218 ( 
.A1(n_1088),
.A2(n_545),
.B1(n_730),
.B2(n_870),
.Y(n_1218)
);

NAND2xp5_ASAP7_75t_L g1219 ( 
.A(n_1106),
.B(n_1109),
.Y(n_1219)
);

AO31x2_ASAP7_75t_L g1220 ( 
.A1(n_1102),
.A2(n_1082),
.A3(n_1012),
.B(n_965),
.Y(n_1220)
);

AOI21xp5_ASAP7_75t_L g1221 ( 
.A1(n_990),
.A2(n_704),
.B(n_941),
.Y(n_1221)
);

OR2x2_ASAP7_75t_L g1222 ( 
.A(n_1106),
.B(n_463),
.Y(n_1222)
);

AOI21xp5_ASAP7_75t_L g1223 ( 
.A1(n_990),
.A2(n_704),
.B(n_941),
.Y(n_1223)
);

CKINVDCx6p67_ASAP7_75t_R g1224 ( 
.A(n_1046),
.Y(n_1224)
);

BUFx2_ASAP7_75t_L g1225 ( 
.A(n_985),
.Y(n_1225)
);

AOI21xp5_ASAP7_75t_L g1226 ( 
.A1(n_990),
.A2(n_704),
.B(n_941),
.Y(n_1226)
);

AO31x2_ASAP7_75t_L g1227 ( 
.A1(n_1102),
.A2(n_1082),
.A3(n_1012),
.B(n_965),
.Y(n_1227)
);

INVx1_ASAP7_75t_SL g1228 ( 
.A(n_985),
.Y(n_1228)
);

AOI21xp5_ASAP7_75t_SL g1229 ( 
.A1(n_1012),
.A2(n_704),
.B(n_685),
.Y(n_1229)
);

NAND2xp5_ASAP7_75t_L g1230 ( 
.A(n_1106),
.B(n_1109),
.Y(n_1230)
);

INVx3_ASAP7_75t_SL g1231 ( 
.A(n_1046),
.Y(n_1231)
);

AO31x2_ASAP7_75t_L g1232 ( 
.A1(n_1102),
.A2(n_1082),
.A3(n_1012),
.B(n_965),
.Y(n_1232)
);

O2A1O1Ixp33_ASAP7_75t_SL g1233 ( 
.A1(n_1012),
.A2(n_831),
.B(n_1052),
.C(n_1016),
.Y(n_1233)
);

NOR2xp33_ASAP7_75t_L g1234 ( 
.A(n_1106),
.B(n_637),
.Y(n_1234)
);

INVx4_ASAP7_75t_L g1235 ( 
.A(n_1085),
.Y(n_1235)
);

NAND2xp5_ASAP7_75t_L g1236 ( 
.A(n_1106),
.B(n_1109),
.Y(n_1236)
);

AOI21x1_ASAP7_75t_L g1237 ( 
.A1(n_1014),
.A2(n_1101),
.B(n_1021),
.Y(n_1237)
);

AOI21xp5_ASAP7_75t_L g1238 ( 
.A1(n_990),
.A2(n_704),
.B(n_941),
.Y(n_1238)
);

INVx4_ASAP7_75t_L g1239 ( 
.A(n_1085),
.Y(n_1239)
);

INVx1_ASAP7_75t_L g1240 ( 
.A(n_1112),
.Y(n_1240)
);

BUFx2_ASAP7_75t_L g1241 ( 
.A(n_1225),
.Y(n_1241)
);

INVx1_ASAP7_75t_L g1242 ( 
.A(n_1183),
.Y(n_1242)
);

INVx1_ASAP7_75t_L g1243 ( 
.A(n_1186),
.Y(n_1243)
);

OAI22xp33_ASAP7_75t_L g1244 ( 
.A1(n_1113),
.A2(n_1209),
.B1(n_1116),
.B2(n_1180),
.Y(n_1244)
);

INVx1_ASAP7_75t_SL g1245 ( 
.A(n_1111),
.Y(n_1245)
);

INVx1_ASAP7_75t_SL g1246 ( 
.A(n_1111),
.Y(n_1246)
);

AOI22xp33_ASAP7_75t_L g1247 ( 
.A1(n_1188),
.A2(n_1113),
.B1(n_1116),
.B2(n_1180),
.Y(n_1247)
);

BUFx8_ASAP7_75t_SL g1248 ( 
.A(n_1161),
.Y(n_1248)
);

CKINVDCx5p33_ASAP7_75t_R g1249 ( 
.A(n_1215),
.Y(n_1249)
);

NAND2xp5_ASAP7_75t_L g1250 ( 
.A(n_1189),
.B(n_1207),
.Y(n_1250)
);

INVx1_ASAP7_75t_L g1251 ( 
.A(n_1212),
.Y(n_1251)
);

AOI22xp33_ASAP7_75t_L g1252 ( 
.A1(n_1137),
.A2(n_1130),
.B1(n_1110),
.B2(n_1200),
.Y(n_1252)
);

NAND2x1p5_ASAP7_75t_L g1253 ( 
.A(n_1194),
.B(n_1146),
.Y(n_1253)
);

BUFx12f_ASAP7_75t_L g1254 ( 
.A(n_1149),
.Y(n_1254)
);

OAI22xp33_ASAP7_75t_R g1255 ( 
.A1(n_1208),
.A2(n_1234),
.B1(n_1222),
.B2(n_1218),
.Y(n_1255)
);

AOI22xp33_ASAP7_75t_L g1256 ( 
.A1(n_1198),
.A2(n_1200),
.B1(n_1118),
.B2(n_1187),
.Y(n_1256)
);

BUFx2_ASAP7_75t_L g1257 ( 
.A(n_1190),
.Y(n_1257)
);

OAI21xp5_ASAP7_75t_SL g1258 ( 
.A1(n_1193),
.A2(n_1201),
.B(n_1206),
.Y(n_1258)
);

BUFx12f_ASAP7_75t_L g1259 ( 
.A(n_1148),
.Y(n_1259)
);

INVx4_ASAP7_75t_L g1260 ( 
.A(n_1194),
.Y(n_1260)
);

AOI22xp33_ASAP7_75t_SL g1261 ( 
.A1(n_1198),
.A2(n_1115),
.B1(n_1195),
.B2(n_1118),
.Y(n_1261)
);

INVx6_ASAP7_75t_L g1262 ( 
.A(n_1194),
.Y(n_1262)
);

CKINVDCx6p67_ASAP7_75t_R g1263 ( 
.A(n_1231),
.Y(n_1263)
);

AOI22xp33_ASAP7_75t_L g1264 ( 
.A1(n_1195),
.A2(n_1115),
.B1(n_1123),
.B2(n_1230),
.Y(n_1264)
);

AOI22xp33_ASAP7_75t_L g1265 ( 
.A1(n_1123),
.A2(n_1219),
.B1(n_1182),
.B2(n_1236),
.Y(n_1265)
);

AOI21xp5_ASAP7_75t_L g1266 ( 
.A1(n_1136),
.A2(n_1121),
.B(n_1229),
.Y(n_1266)
);

CKINVDCx11_ASAP7_75t_R g1267 ( 
.A(n_1147),
.Y(n_1267)
);

AOI22xp33_ASAP7_75t_L g1268 ( 
.A1(n_1182),
.A2(n_1192),
.B1(n_1230),
.B2(n_1236),
.Y(n_1268)
);

NAND2x1p5_ASAP7_75t_L g1269 ( 
.A(n_1194),
.B(n_1173),
.Y(n_1269)
);

BUFx12f_ASAP7_75t_L g1270 ( 
.A(n_1148),
.Y(n_1270)
);

CKINVDCx20_ASAP7_75t_R g1271 ( 
.A(n_1224),
.Y(n_1271)
);

BUFx6f_ASAP7_75t_L g1272 ( 
.A(n_1173),
.Y(n_1272)
);

AOI22xp33_ASAP7_75t_L g1273 ( 
.A1(n_1192),
.A2(n_1219),
.B1(n_1129),
.B2(n_1127),
.Y(n_1273)
);

INVx6_ASAP7_75t_L g1274 ( 
.A(n_1235),
.Y(n_1274)
);

BUFx6f_ASAP7_75t_L g1275 ( 
.A(n_1171),
.Y(n_1275)
);

AOI22xp33_ASAP7_75t_SL g1276 ( 
.A1(n_1196),
.A2(n_1210),
.B1(n_1134),
.B2(n_1129),
.Y(n_1276)
);

AOI22xp33_ASAP7_75t_SL g1277 ( 
.A1(n_1134),
.A2(n_1190),
.B1(n_1202),
.B2(n_1213),
.Y(n_1277)
);

CKINVDCx11_ASAP7_75t_R g1278 ( 
.A(n_1199),
.Y(n_1278)
);

INVx6_ASAP7_75t_L g1279 ( 
.A(n_1235),
.Y(n_1279)
);

INVx3_ASAP7_75t_SL g1280 ( 
.A(n_1239),
.Y(n_1280)
);

AOI22xp33_ASAP7_75t_SL g1281 ( 
.A1(n_1202),
.A2(n_1164),
.B1(n_1205),
.B2(n_1184),
.Y(n_1281)
);

AOI22xp33_ASAP7_75t_L g1282 ( 
.A1(n_1131),
.A2(n_1159),
.B1(n_1140),
.B2(n_1169),
.Y(n_1282)
);

CKINVDCx6p67_ASAP7_75t_R g1283 ( 
.A(n_1239),
.Y(n_1283)
);

CKINVDCx5p33_ASAP7_75t_R g1284 ( 
.A(n_1199),
.Y(n_1284)
);

CKINVDCx11_ASAP7_75t_R g1285 ( 
.A(n_1228),
.Y(n_1285)
);

INVx6_ASAP7_75t_L g1286 ( 
.A(n_1170),
.Y(n_1286)
);

CKINVDCx5p33_ASAP7_75t_R g1287 ( 
.A(n_1133),
.Y(n_1287)
);

AOI22xp33_ASAP7_75t_SL g1288 ( 
.A1(n_1153),
.A2(n_1185),
.B1(n_1142),
.B2(n_1233),
.Y(n_1288)
);

NAND2xp5_ASAP7_75t_L g1289 ( 
.A(n_1132),
.B(n_1141),
.Y(n_1289)
);

AOI22xp33_ASAP7_75t_L g1290 ( 
.A1(n_1159),
.A2(n_1135),
.B1(n_1126),
.B2(n_1125),
.Y(n_1290)
);

OR2x2_ASAP7_75t_L g1291 ( 
.A(n_1152),
.B(n_1191),
.Y(n_1291)
);

CKINVDCx20_ASAP7_75t_R g1292 ( 
.A(n_1157),
.Y(n_1292)
);

AOI22xp33_ASAP7_75t_L g1293 ( 
.A1(n_1119),
.A2(n_1204),
.B1(n_1158),
.B2(n_1141),
.Y(n_1293)
);

AOI22xp33_ASAP7_75t_SL g1294 ( 
.A1(n_1119),
.A2(n_1122),
.B1(n_1176),
.B2(n_1150),
.Y(n_1294)
);

BUFx3_ASAP7_75t_L g1295 ( 
.A(n_1160),
.Y(n_1295)
);

AOI22xp33_ASAP7_75t_L g1296 ( 
.A1(n_1158),
.A2(n_1139),
.B1(n_1155),
.B2(n_1145),
.Y(n_1296)
);

INVx1_ASAP7_75t_L g1297 ( 
.A(n_1167),
.Y(n_1297)
);

OAI22xp5_ASAP7_75t_L g1298 ( 
.A1(n_1154),
.A2(n_1163),
.B1(n_1172),
.B2(n_1174),
.Y(n_1298)
);

AOI22xp33_ASAP7_75t_L g1299 ( 
.A1(n_1176),
.A2(n_1168),
.B1(n_1167),
.B2(n_1162),
.Y(n_1299)
);

AOI22xp33_ASAP7_75t_L g1300 ( 
.A1(n_1168),
.A2(n_1156),
.B1(n_1120),
.B2(n_1150),
.Y(n_1300)
);

AOI22xp33_ASAP7_75t_L g1301 ( 
.A1(n_1150),
.A2(n_1144),
.B1(n_1203),
.B2(n_1166),
.Y(n_1301)
);

INVx1_ASAP7_75t_L g1302 ( 
.A(n_1151),
.Y(n_1302)
);

BUFx4f_ASAP7_75t_SL g1303 ( 
.A(n_1124),
.Y(n_1303)
);

INVx6_ASAP7_75t_L g1304 ( 
.A(n_1165),
.Y(n_1304)
);

INVx6_ASAP7_75t_L g1305 ( 
.A(n_1143),
.Y(n_1305)
);

AOI22xp33_ASAP7_75t_L g1306 ( 
.A1(n_1203),
.A2(n_1128),
.B1(n_1226),
.B2(n_1223),
.Y(n_1306)
);

INVx6_ASAP7_75t_L g1307 ( 
.A(n_1217),
.Y(n_1307)
);

BUFx8_ASAP7_75t_L g1308 ( 
.A(n_1178),
.Y(n_1308)
);

OAI22xp33_ASAP7_75t_L g1309 ( 
.A1(n_1177),
.A2(n_1237),
.B1(n_1238),
.B2(n_1221),
.Y(n_1309)
);

AOI22xp33_ASAP7_75t_L g1310 ( 
.A1(n_1203),
.A2(n_1214),
.B1(n_1178),
.B2(n_1232),
.Y(n_1310)
);

INVx1_ASAP7_75t_L g1311 ( 
.A(n_1175),
.Y(n_1311)
);

OAI22xp33_ASAP7_75t_L g1312 ( 
.A1(n_1178),
.A2(n_1114),
.B1(n_1227),
.B2(n_1220),
.Y(n_1312)
);

CKINVDCx11_ASAP7_75t_R g1313 ( 
.A(n_1114),
.Y(n_1313)
);

AOI22xp33_ASAP7_75t_SL g1314 ( 
.A1(n_1114),
.A2(n_1232),
.B1(n_1227),
.B2(n_1220),
.Y(n_1314)
);

AND2x2_ASAP7_75t_L g1315 ( 
.A(n_1181),
.B(n_1232),
.Y(n_1315)
);

CKINVDCx11_ASAP7_75t_R g1316 ( 
.A(n_1181),
.Y(n_1316)
);

BUFx4f_ASAP7_75t_SL g1317 ( 
.A(n_1181),
.Y(n_1317)
);

AOI22xp33_ASAP7_75t_SL g1318 ( 
.A1(n_1220),
.A2(n_1227),
.B1(n_1117),
.B2(n_1179),
.Y(n_1318)
);

NAND2xp5_ASAP7_75t_L g1319 ( 
.A(n_1175),
.B(n_1138),
.Y(n_1319)
);

INVx2_ASAP7_75t_L g1320 ( 
.A(n_1138),
.Y(n_1320)
);

INVx4_ASAP7_75t_L g1321 ( 
.A(n_1138),
.Y(n_1321)
);

INVx1_ASAP7_75t_L g1322 ( 
.A(n_1197),
.Y(n_1322)
);

NAND2x1p5_ASAP7_75t_L g1323 ( 
.A(n_1211),
.B(n_1216),
.Y(n_1323)
);

AOI21xp5_ASAP7_75t_SL g1324 ( 
.A1(n_1193),
.A2(n_1206),
.B(n_1201),
.Y(n_1324)
);

OAI22xp5_ASAP7_75t_SL g1325 ( 
.A1(n_1188),
.A2(n_1130),
.B1(n_1065),
.B2(n_997),
.Y(n_1325)
);

NAND2xp5_ASAP7_75t_L g1326 ( 
.A(n_1189),
.B(n_1106),
.Y(n_1326)
);

HB1xp67_ASAP7_75t_L g1327 ( 
.A(n_1133),
.Y(n_1327)
);

INVx4_ASAP7_75t_L g1328 ( 
.A(n_1194),
.Y(n_1328)
);

AOI22xp33_ASAP7_75t_L g1329 ( 
.A1(n_1188),
.A2(n_1209),
.B1(n_1113),
.B2(n_1116),
.Y(n_1329)
);

BUFx4_ASAP7_75t_R g1330 ( 
.A(n_1185),
.Y(n_1330)
);

OAI22xp5_ASAP7_75t_L g1331 ( 
.A1(n_1188),
.A2(n_1130),
.B1(n_1116),
.B2(n_1180),
.Y(n_1331)
);

CKINVDCx20_ASAP7_75t_R g1332 ( 
.A(n_1215),
.Y(n_1332)
);

AOI22xp33_ASAP7_75t_L g1333 ( 
.A1(n_1188),
.A2(n_1209),
.B1(n_1113),
.B2(n_1116),
.Y(n_1333)
);

NAND2xp5_ASAP7_75t_L g1334 ( 
.A(n_1189),
.B(n_1106),
.Y(n_1334)
);

BUFx3_ASAP7_75t_L g1335 ( 
.A(n_1225),
.Y(n_1335)
);

AOI22xp33_ASAP7_75t_L g1336 ( 
.A1(n_1188),
.A2(n_1209),
.B1(n_1113),
.B2(n_1116),
.Y(n_1336)
);

OAI21xp5_ASAP7_75t_SL g1337 ( 
.A1(n_1188),
.A2(n_1209),
.B(n_1130),
.Y(n_1337)
);

NAND2x1p5_ASAP7_75t_L g1338 ( 
.A(n_1194),
.B(n_1011),
.Y(n_1338)
);

AOI22xp33_ASAP7_75t_L g1339 ( 
.A1(n_1188),
.A2(n_1209),
.B1(n_1113),
.B2(n_1116),
.Y(n_1339)
);

AOI22xp33_ASAP7_75t_L g1340 ( 
.A1(n_1188),
.A2(n_1209),
.B1(n_1113),
.B2(n_1116),
.Y(n_1340)
);

BUFx3_ASAP7_75t_L g1341 ( 
.A(n_1225),
.Y(n_1341)
);

OAI22xp5_ASAP7_75t_L g1342 ( 
.A1(n_1188),
.A2(n_1130),
.B1(n_1116),
.B2(n_1180),
.Y(n_1342)
);

BUFx12f_ASAP7_75t_L g1343 ( 
.A(n_1149),
.Y(n_1343)
);

AOI22xp33_ASAP7_75t_L g1344 ( 
.A1(n_1188),
.A2(n_1209),
.B1(n_1113),
.B2(n_1116),
.Y(n_1344)
);

BUFx10_ASAP7_75t_L g1345 ( 
.A(n_1215),
.Y(n_1345)
);

BUFx10_ASAP7_75t_L g1346 ( 
.A(n_1215),
.Y(n_1346)
);

INVx6_ASAP7_75t_L g1347 ( 
.A(n_1194),
.Y(n_1347)
);

CKINVDCx20_ASAP7_75t_R g1348 ( 
.A(n_1215),
.Y(n_1348)
);

INVx1_ASAP7_75t_L g1349 ( 
.A(n_1112),
.Y(n_1349)
);

BUFx3_ASAP7_75t_L g1350 ( 
.A(n_1225),
.Y(n_1350)
);

AOI22xp33_ASAP7_75t_L g1351 ( 
.A1(n_1188),
.A2(n_1209),
.B1(n_1113),
.B2(n_1116),
.Y(n_1351)
);

BUFx2_ASAP7_75t_SL g1352 ( 
.A(n_1147),
.Y(n_1352)
);

AOI22xp33_ASAP7_75t_L g1353 ( 
.A1(n_1188),
.A2(n_1209),
.B1(n_1113),
.B2(n_1116),
.Y(n_1353)
);

INVx1_ASAP7_75t_L g1354 ( 
.A(n_1302),
.Y(n_1354)
);

INVx5_ASAP7_75t_L g1355 ( 
.A(n_1307),
.Y(n_1355)
);

INVx1_ASAP7_75t_L g1356 ( 
.A(n_1311),
.Y(n_1356)
);

BUFx2_ASAP7_75t_L g1357 ( 
.A(n_1308),
.Y(n_1357)
);

INVx1_ASAP7_75t_L g1358 ( 
.A(n_1319),
.Y(n_1358)
);

INVxp67_ASAP7_75t_L g1359 ( 
.A(n_1327),
.Y(n_1359)
);

HB1xp67_ASAP7_75t_L g1360 ( 
.A(n_1320),
.Y(n_1360)
);

INVx1_ASAP7_75t_L g1361 ( 
.A(n_1315),
.Y(n_1361)
);

INVx1_ASAP7_75t_L g1362 ( 
.A(n_1289),
.Y(n_1362)
);

BUFx3_ASAP7_75t_L g1363 ( 
.A(n_1286),
.Y(n_1363)
);

AND2x2_ASAP7_75t_L g1364 ( 
.A(n_1261),
.B(n_1264),
.Y(n_1364)
);

OAI21x1_ASAP7_75t_L g1365 ( 
.A1(n_1266),
.A2(n_1323),
.B(n_1306),
.Y(n_1365)
);

AND2x2_ASAP7_75t_L g1366 ( 
.A(n_1264),
.B(n_1314),
.Y(n_1366)
);

INVx1_ASAP7_75t_L g1367 ( 
.A(n_1312),
.Y(n_1367)
);

INVx1_ASAP7_75t_L g1368 ( 
.A(n_1317),
.Y(n_1368)
);

BUFx3_ASAP7_75t_L g1369 ( 
.A(n_1286),
.Y(n_1369)
);

OAI21xp5_ASAP7_75t_L g1370 ( 
.A1(n_1324),
.A2(n_1258),
.B(n_1244),
.Y(n_1370)
);

INVx1_ASAP7_75t_L g1371 ( 
.A(n_1321),
.Y(n_1371)
);

INVx2_ASAP7_75t_L g1372 ( 
.A(n_1322),
.Y(n_1372)
);

OAI21x1_ASAP7_75t_L g1373 ( 
.A1(n_1323),
.A2(n_1306),
.B(n_1300),
.Y(n_1373)
);

INVx5_ASAP7_75t_L g1374 ( 
.A(n_1304),
.Y(n_1374)
);

OAI22xp5_ASAP7_75t_L g1375 ( 
.A1(n_1329),
.A2(n_1353),
.B1(n_1351),
.B2(n_1344),
.Y(n_1375)
);

INVx1_ASAP7_75t_SL g1376 ( 
.A(n_1245),
.Y(n_1376)
);

OAI21xp5_ASAP7_75t_L g1377 ( 
.A1(n_1331),
.A2(n_1342),
.B(n_1351),
.Y(n_1377)
);

INVx1_ASAP7_75t_L g1378 ( 
.A(n_1294),
.Y(n_1378)
);

AO21x2_ASAP7_75t_L g1379 ( 
.A1(n_1309),
.A2(n_1298),
.B(n_1349),
.Y(n_1379)
);

OR2x2_ASAP7_75t_L g1380 ( 
.A(n_1256),
.B(n_1273),
.Y(n_1380)
);

BUFx2_ASAP7_75t_L g1381 ( 
.A(n_1308),
.Y(n_1381)
);

AOI22xp5_ASAP7_75t_L g1382 ( 
.A1(n_1325),
.A2(n_1337),
.B1(n_1329),
.B2(n_1344),
.Y(n_1382)
);

INVx1_ASAP7_75t_L g1383 ( 
.A(n_1240),
.Y(n_1383)
);

INVx1_ASAP7_75t_L g1384 ( 
.A(n_1242),
.Y(n_1384)
);

AND2x2_ASAP7_75t_L g1385 ( 
.A(n_1256),
.B(n_1313),
.Y(n_1385)
);

BUFx2_ASAP7_75t_L g1386 ( 
.A(n_1304),
.Y(n_1386)
);

INVx1_ASAP7_75t_L g1387 ( 
.A(n_1243),
.Y(n_1387)
);

INVx1_ASAP7_75t_SL g1388 ( 
.A(n_1246),
.Y(n_1388)
);

BUFx2_ASAP7_75t_SL g1389 ( 
.A(n_1295),
.Y(n_1389)
);

NAND2xp5_ASAP7_75t_L g1390 ( 
.A(n_1273),
.B(n_1265),
.Y(n_1390)
);

INVx1_ASAP7_75t_L g1391 ( 
.A(n_1251),
.Y(n_1391)
);

OAI21xp5_ASAP7_75t_L g1392 ( 
.A1(n_1333),
.A2(n_1353),
.B(n_1339),
.Y(n_1392)
);

AND2x2_ASAP7_75t_L g1393 ( 
.A(n_1316),
.B(n_1247),
.Y(n_1393)
);

AND2x2_ASAP7_75t_L g1394 ( 
.A(n_1247),
.B(n_1276),
.Y(n_1394)
);

OAI21x1_ASAP7_75t_L g1395 ( 
.A1(n_1300),
.A2(n_1299),
.B(n_1301),
.Y(n_1395)
);

NOR2xp33_ASAP7_75t_L g1396 ( 
.A(n_1250),
.B(n_1326),
.Y(n_1396)
);

OAI21x1_ASAP7_75t_L g1397 ( 
.A1(n_1299),
.A2(n_1301),
.B(n_1310),
.Y(n_1397)
);

HB1xp67_ASAP7_75t_L g1398 ( 
.A(n_1304),
.Y(n_1398)
);

NAND2xp5_ASAP7_75t_L g1399 ( 
.A(n_1265),
.B(n_1268),
.Y(n_1399)
);

AND2x2_ASAP7_75t_L g1400 ( 
.A(n_1252),
.B(n_1310),
.Y(n_1400)
);

OR2x2_ASAP7_75t_L g1401 ( 
.A(n_1252),
.B(n_1293),
.Y(n_1401)
);

BUFx3_ASAP7_75t_L g1402 ( 
.A(n_1262),
.Y(n_1402)
);

AND2x2_ASAP7_75t_L g1403 ( 
.A(n_1290),
.B(n_1277),
.Y(n_1403)
);

INVx3_ASAP7_75t_L g1404 ( 
.A(n_1305),
.Y(n_1404)
);

INVx1_ASAP7_75t_SL g1405 ( 
.A(n_1241),
.Y(n_1405)
);

BUFx2_ASAP7_75t_L g1406 ( 
.A(n_1303),
.Y(n_1406)
);

OAI21x1_ASAP7_75t_L g1407 ( 
.A1(n_1290),
.A2(n_1293),
.B(n_1296),
.Y(n_1407)
);

NOR2x1_ASAP7_75t_SL g1408 ( 
.A(n_1260),
.B(n_1328),
.Y(n_1408)
);

AND2x2_ASAP7_75t_L g1409 ( 
.A(n_1296),
.B(n_1268),
.Y(n_1409)
);

INVx4_ASAP7_75t_L g1410 ( 
.A(n_1330),
.Y(n_1410)
);

INVx1_ASAP7_75t_L g1411 ( 
.A(n_1297),
.Y(n_1411)
);

INVx1_ASAP7_75t_L g1412 ( 
.A(n_1318),
.Y(n_1412)
);

BUFx2_ASAP7_75t_L g1413 ( 
.A(n_1335),
.Y(n_1413)
);

OA21x2_ASAP7_75t_L g1414 ( 
.A1(n_1333),
.A2(n_1336),
.B(n_1339),
.Y(n_1414)
);

NAND2xp5_ASAP7_75t_L g1415 ( 
.A(n_1334),
.B(n_1336),
.Y(n_1415)
);

INVx1_ASAP7_75t_L g1416 ( 
.A(n_1281),
.Y(n_1416)
);

OAI22xp5_ASAP7_75t_L g1417 ( 
.A1(n_1340),
.A2(n_1282),
.B1(n_1288),
.B2(n_1284),
.Y(n_1417)
);

BUFx2_ASAP7_75t_L g1418 ( 
.A(n_1341),
.Y(n_1418)
);

INVx1_ASAP7_75t_L g1419 ( 
.A(n_1262),
.Y(n_1419)
);

OAI22xp5_ASAP7_75t_L g1420 ( 
.A1(n_1382),
.A2(n_1340),
.B1(n_1282),
.B2(n_1287),
.Y(n_1420)
);

AND2x2_ASAP7_75t_L g1421 ( 
.A(n_1361),
.B(n_1257),
.Y(n_1421)
);

OAI21xp5_ASAP7_75t_L g1422 ( 
.A1(n_1370),
.A2(n_1253),
.B(n_1292),
.Y(n_1422)
);

NAND2xp5_ASAP7_75t_L g1423 ( 
.A(n_1396),
.B(n_1350),
.Y(n_1423)
);

AND2x2_ASAP7_75t_L g1424 ( 
.A(n_1413),
.B(n_1350),
.Y(n_1424)
);

BUFx12f_ASAP7_75t_L g1425 ( 
.A(n_1406),
.Y(n_1425)
);

AND2x6_ASAP7_75t_L g1426 ( 
.A(n_1362),
.B(n_1330),
.Y(n_1426)
);

OAI21xp5_ASAP7_75t_L g1427 ( 
.A1(n_1370),
.A2(n_1291),
.B(n_1269),
.Y(n_1427)
);

OAI21x1_ASAP7_75t_SL g1428 ( 
.A1(n_1377),
.A2(n_1255),
.B(n_1254),
.Y(n_1428)
);

OAI221xp5_ASAP7_75t_L g1429 ( 
.A1(n_1382),
.A2(n_1280),
.B1(n_1352),
.B2(n_1274),
.C(n_1279),
.Y(n_1429)
);

INVxp67_ASAP7_75t_L g1430 ( 
.A(n_1376),
.Y(n_1430)
);

O2A1O1Ixp5_ASAP7_75t_SL g1431 ( 
.A1(n_1377),
.A2(n_1278),
.B(n_1285),
.C(n_1274),
.Y(n_1431)
);

OAI22xp5_ASAP7_75t_L g1432 ( 
.A1(n_1375),
.A2(n_1274),
.B1(n_1279),
.B2(n_1280),
.Y(n_1432)
);

AND2x2_ASAP7_75t_L g1433 ( 
.A(n_1397),
.B(n_1275),
.Y(n_1433)
);

OR2x6_ASAP7_75t_L g1434 ( 
.A(n_1410),
.B(n_1347),
.Y(n_1434)
);

AND2x2_ASAP7_75t_L g1435 ( 
.A(n_1397),
.B(n_1275),
.Y(n_1435)
);

OAI21x1_ASAP7_75t_L g1436 ( 
.A1(n_1365),
.A2(n_1338),
.B(n_1269),
.Y(n_1436)
);

NAND2xp5_ASAP7_75t_L g1437 ( 
.A(n_1415),
.B(n_1272),
.Y(n_1437)
);

AOI221xp5_ASAP7_75t_L g1438 ( 
.A1(n_1375),
.A2(n_1271),
.B1(n_1249),
.B2(n_1332),
.C(n_1348),
.Y(n_1438)
);

HB1xp67_ASAP7_75t_L g1439 ( 
.A(n_1360),
.Y(n_1439)
);

NOR2xp67_ASAP7_75t_L g1440 ( 
.A(n_1398),
.B(n_1359),
.Y(n_1440)
);

AND2x4_ASAP7_75t_L g1441 ( 
.A(n_1374),
.B(n_1368),
.Y(n_1441)
);

AND2x4_ASAP7_75t_L g1442 ( 
.A(n_1374),
.B(n_1279),
.Y(n_1442)
);

NAND2xp33_ASAP7_75t_L g1443 ( 
.A(n_1392),
.B(n_1283),
.Y(n_1443)
);

AOI21xp5_ASAP7_75t_L g1444 ( 
.A1(n_1374),
.A2(n_1347),
.B(n_1270),
.Y(n_1444)
);

AND2x2_ASAP7_75t_L g1445 ( 
.A(n_1418),
.B(n_1346),
.Y(n_1445)
);

AOI221xp5_ASAP7_75t_L g1446 ( 
.A1(n_1392),
.A2(n_1263),
.B1(n_1259),
.B2(n_1270),
.C(n_1267),
.Y(n_1446)
);

AND2x2_ASAP7_75t_L g1447 ( 
.A(n_1397),
.B(n_1378),
.Y(n_1447)
);

NAND2xp5_ASAP7_75t_L g1448 ( 
.A(n_1359),
.B(n_1345),
.Y(n_1448)
);

A2O1A1Ixp33_ASAP7_75t_L g1449 ( 
.A1(n_1417),
.A2(n_1259),
.B(n_1254),
.C(n_1343),
.Y(n_1449)
);

OR2x2_ASAP7_75t_L g1450 ( 
.A(n_1383),
.B(n_1345),
.Y(n_1450)
);

AO32x1_ASAP7_75t_L g1451 ( 
.A1(n_1417),
.A2(n_1248),
.A3(n_1343),
.B1(n_1346),
.B2(n_1378),
.Y(n_1451)
);

OAI211xp5_ASAP7_75t_L g1452 ( 
.A1(n_1414),
.A2(n_1364),
.B(n_1416),
.C(n_1394),
.Y(n_1452)
);

A2O1A1Ixp33_ASAP7_75t_L g1453 ( 
.A1(n_1403),
.A2(n_1364),
.B(n_1394),
.C(n_1416),
.Y(n_1453)
);

A2O1A1Ixp33_ASAP7_75t_L g1454 ( 
.A1(n_1403),
.A2(n_1385),
.B(n_1380),
.C(n_1407),
.Y(n_1454)
);

OAI21x1_ASAP7_75t_L g1455 ( 
.A1(n_1365),
.A2(n_1373),
.B(n_1407),
.Y(n_1455)
);

OAI211xp5_ASAP7_75t_L g1456 ( 
.A1(n_1414),
.A2(n_1393),
.B(n_1399),
.C(n_1390),
.Y(n_1456)
);

O2A1O1Ixp33_ASAP7_75t_SL g1457 ( 
.A1(n_1380),
.A2(n_1401),
.B(n_1399),
.C(n_1390),
.Y(n_1457)
);

AND2x2_ASAP7_75t_L g1458 ( 
.A(n_1366),
.B(n_1367),
.Y(n_1458)
);

INVx2_ASAP7_75t_L g1459 ( 
.A(n_1372),
.Y(n_1459)
);

O2A1O1Ixp5_ASAP7_75t_L g1460 ( 
.A1(n_1410),
.A2(n_1409),
.B(n_1401),
.C(n_1404),
.Y(n_1460)
);

OR2x2_ASAP7_75t_L g1461 ( 
.A(n_1384),
.B(n_1387),
.Y(n_1461)
);

NOR2x1_ASAP7_75t_SL g1462 ( 
.A(n_1374),
.B(n_1379),
.Y(n_1462)
);

NAND2xp5_ASAP7_75t_L g1463 ( 
.A(n_1376),
.B(n_1388),
.Y(n_1463)
);

BUFx12f_ASAP7_75t_L g1464 ( 
.A(n_1406),
.Y(n_1464)
);

NAND2xp5_ASAP7_75t_L g1465 ( 
.A(n_1388),
.B(n_1405),
.Y(n_1465)
);

OAI21xp5_ASAP7_75t_L g1466 ( 
.A1(n_1414),
.A2(n_1407),
.B(n_1409),
.Y(n_1466)
);

AND2x4_ASAP7_75t_L g1467 ( 
.A(n_1404),
.B(n_1387),
.Y(n_1467)
);

NOR2xp33_ASAP7_75t_L g1468 ( 
.A(n_1398),
.B(n_1386),
.Y(n_1468)
);

AO32x2_ASAP7_75t_L g1469 ( 
.A1(n_1410),
.A2(n_1358),
.A3(n_1395),
.B1(n_1356),
.B2(n_1412),
.Y(n_1469)
);

AND2x2_ASAP7_75t_L g1470 ( 
.A(n_1418),
.B(n_1363),
.Y(n_1470)
);

NAND2xp5_ASAP7_75t_L g1471 ( 
.A(n_1405),
.B(n_1411),
.Y(n_1471)
);

AOI221xp5_ASAP7_75t_L g1472 ( 
.A1(n_1393),
.A2(n_1385),
.B1(n_1400),
.B2(n_1412),
.C(n_1379),
.Y(n_1472)
);

AOI22xp33_ASAP7_75t_L g1473 ( 
.A1(n_1420),
.A2(n_1414),
.B1(n_1400),
.B2(n_1379),
.Y(n_1473)
);

BUFx6f_ASAP7_75t_L g1474 ( 
.A(n_1455),
.Y(n_1474)
);

NOR2xp33_ASAP7_75t_L g1475 ( 
.A(n_1452),
.B(n_1386),
.Y(n_1475)
);

AND2x2_ASAP7_75t_L g1476 ( 
.A(n_1447),
.B(n_1395),
.Y(n_1476)
);

AOI22xp33_ASAP7_75t_L g1477 ( 
.A1(n_1428),
.A2(n_1414),
.B1(n_1379),
.B2(n_1357),
.Y(n_1477)
);

HB1xp67_ASAP7_75t_L g1478 ( 
.A(n_1439),
.Y(n_1478)
);

AND2x4_ASAP7_75t_L g1479 ( 
.A(n_1433),
.B(n_1355),
.Y(n_1479)
);

INVxp67_ASAP7_75t_L g1480 ( 
.A(n_1447),
.Y(n_1480)
);

AND2x2_ASAP7_75t_L g1481 ( 
.A(n_1469),
.B(n_1395),
.Y(n_1481)
);

AND2x2_ASAP7_75t_L g1482 ( 
.A(n_1469),
.B(n_1373),
.Y(n_1482)
);

INVxp67_ASAP7_75t_L g1483 ( 
.A(n_1461),
.Y(n_1483)
);

BUFx2_ASAP7_75t_L g1484 ( 
.A(n_1435),
.Y(n_1484)
);

OR2x2_ASAP7_75t_L g1485 ( 
.A(n_1466),
.B(n_1356),
.Y(n_1485)
);

AOI22xp33_ASAP7_75t_L g1486 ( 
.A1(n_1443),
.A2(n_1381),
.B1(n_1357),
.B2(n_1410),
.Y(n_1486)
);

INVxp67_ASAP7_75t_SL g1487 ( 
.A(n_1439),
.Y(n_1487)
);

INVx1_ASAP7_75t_L g1488 ( 
.A(n_1459),
.Y(n_1488)
);

INVx1_ASAP7_75t_L g1489 ( 
.A(n_1459),
.Y(n_1489)
);

NOR2x1p5_ASAP7_75t_L g1490 ( 
.A(n_1425),
.B(n_1369),
.Y(n_1490)
);

INVx1_ASAP7_75t_L g1491 ( 
.A(n_1471),
.Y(n_1491)
);

NOR2x1_ASAP7_75t_L g1492 ( 
.A(n_1440),
.B(n_1389),
.Y(n_1492)
);

AND2x2_ASAP7_75t_L g1493 ( 
.A(n_1469),
.B(n_1373),
.Y(n_1493)
);

INVx2_ASAP7_75t_L g1494 ( 
.A(n_1469),
.Y(n_1494)
);

AND2x2_ASAP7_75t_L g1495 ( 
.A(n_1455),
.B(n_1462),
.Y(n_1495)
);

INVx2_ASAP7_75t_L g1496 ( 
.A(n_1467),
.Y(n_1496)
);

INVx1_ASAP7_75t_L g1497 ( 
.A(n_1467),
.Y(n_1497)
);

NAND2xp5_ASAP7_75t_L g1498 ( 
.A(n_1458),
.B(n_1454),
.Y(n_1498)
);

INVx1_ASAP7_75t_SL g1499 ( 
.A(n_1450),
.Y(n_1499)
);

NAND2xp5_ASAP7_75t_L g1500 ( 
.A(n_1458),
.B(n_1391),
.Y(n_1500)
);

NAND2xp5_ASAP7_75t_L g1501 ( 
.A(n_1454),
.B(n_1391),
.Y(n_1501)
);

HB1xp67_ASAP7_75t_L g1502 ( 
.A(n_1478),
.Y(n_1502)
);

AND2x2_ASAP7_75t_L g1503 ( 
.A(n_1476),
.B(n_1460),
.Y(n_1503)
);

HB1xp67_ASAP7_75t_L g1504 ( 
.A(n_1478),
.Y(n_1504)
);

AO22x1_ASAP7_75t_L g1505 ( 
.A1(n_1492),
.A2(n_1426),
.B1(n_1422),
.B2(n_1381),
.Y(n_1505)
);

OR2x2_ASAP7_75t_L g1506 ( 
.A(n_1494),
.B(n_1465),
.Y(n_1506)
);

AOI22xp33_ASAP7_75t_L g1507 ( 
.A1(n_1473),
.A2(n_1472),
.B1(n_1443),
.B2(n_1438),
.Y(n_1507)
);

NAND2xp5_ASAP7_75t_L g1508 ( 
.A(n_1491),
.B(n_1456),
.Y(n_1508)
);

NAND2xp5_ASAP7_75t_L g1509 ( 
.A(n_1491),
.B(n_1430),
.Y(n_1509)
);

NAND2x1p5_ASAP7_75t_SL g1510 ( 
.A(n_1492),
.B(n_1451),
.Y(n_1510)
);

AND2x2_ASAP7_75t_L g1511 ( 
.A(n_1476),
.B(n_1470),
.Y(n_1511)
);

OR2x2_ASAP7_75t_L g1512 ( 
.A(n_1494),
.B(n_1463),
.Y(n_1512)
);

AOI22xp33_ASAP7_75t_L g1513 ( 
.A1(n_1473),
.A2(n_1446),
.B1(n_1475),
.B2(n_1498),
.Y(n_1513)
);

INVxp67_ASAP7_75t_SL g1514 ( 
.A(n_1501),
.Y(n_1514)
);

AND2x2_ASAP7_75t_L g1515 ( 
.A(n_1476),
.B(n_1421),
.Y(n_1515)
);

AND2x4_ASAP7_75t_L g1516 ( 
.A(n_1479),
.B(n_1436),
.Y(n_1516)
);

INVx1_ASAP7_75t_L g1517 ( 
.A(n_1487),
.Y(n_1517)
);

INVx2_ASAP7_75t_L g1518 ( 
.A(n_1494),
.Y(n_1518)
);

AND2x2_ASAP7_75t_L g1519 ( 
.A(n_1481),
.B(n_1484),
.Y(n_1519)
);

HB1xp67_ASAP7_75t_L g1520 ( 
.A(n_1480),
.Y(n_1520)
);

AND2x2_ASAP7_75t_L g1521 ( 
.A(n_1481),
.B(n_1371),
.Y(n_1521)
);

AND2x2_ASAP7_75t_L g1522 ( 
.A(n_1481),
.B(n_1371),
.Y(n_1522)
);

INVx1_ASAP7_75t_L g1523 ( 
.A(n_1487),
.Y(n_1523)
);

INVx3_ASAP7_75t_L g1524 ( 
.A(n_1474),
.Y(n_1524)
);

INVx1_ASAP7_75t_L g1525 ( 
.A(n_1488),
.Y(n_1525)
);

OR2x2_ASAP7_75t_L g1526 ( 
.A(n_1494),
.B(n_1354),
.Y(n_1526)
);

HB1xp67_ASAP7_75t_L g1527 ( 
.A(n_1480),
.Y(n_1527)
);

NAND2xp5_ASAP7_75t_L g1528 ( 
.A(n_1483),
.B(n_1457),
.Y(n_1528)
);

AOI22xp33_ASAP7_75t_L g1529 ( 
.A1(n_1475),
.A2(n_1498),
.B1(n_1429),
.B2(n_1477),
.Y(n_1529)
);

NOR2xp33_ASAP7_75t_L g1530 ( 
.A(n_1499),
.B(n_1448),
.Y(n_1530)
);

INVx1_ASAP7_75t_L g1531 ( 
.A(n_1488),
.Y(n_1531)
);

OR2x6_ASAP7_75t_L g1532 ( 
.A(n_1479),
.B(n_1436),
.Y(n_1532)
);

AOI22xp33_ASAP7_75t_L g1533 ( 
.A1(n_1477),
.A2(n_1432),
.B1(n_1426),
.B2(n_1437),
.Y(n_1533)
);

HB1xp67_ASAP7_75t_L g1534 ( 
.A(n_1489),
.Y(n_1534)
);

AND2x2_ASAP7_75t_L g1535 ( 
.A(n_1484),
.B(n_1424),
.Y(n_1535)
);

INVx1_ASAP7_75t_SL g1536 ( 
.A(n_1499),
.Y(n_1536)
);

NAND2xp5_ASAP7_75t_L g1537 ( 
.A(n_1514),
.B(n_1483),
.Y(n_1537)
);

AND2x2_ASAP7_75t_L g1538 ( 
.A(n_1519),
.B(n_1482),
.Y(n_1538)
);

NAND2xp5_ASAP7_75t_L g1539 ( 
.A(n_1514),
.B(n_1501),
.Y(n_1539)
);

AND2x2_ASAP7_75t_L g1540 ( 
.A(n_1519),
.B(n_1482),
.Y(n_1540)
);

INVx1_ASAP7_75t_L g1541 ( 
.A(n_1525),
.Y(n_1541)
);

INVx2_ASAP7_75t_L g1542 ( 
.A(n_1518),
.Y(n_1542)
);

AND2x2_ASAP7_75t_L g1543 ( 
.A(n_1519),
.B(n_1482),
.Y(n_1543)
);

INVx1_ASAP7_75t_L g1544 ( 
.A(n_1525),
.Y(n_1544)
);

AND2x2_ASAP7_75t_L g1545 ( 
.A(n_1503),
.B(n_1493),
.Y(n_1545)
);

INVx2_ASAP7_75t_L g1546 ( 
.A(n_1518),
.Y(n_1546)
);

INVx1_ASAP7_75t_SL g1547 ( 
.A(n_1536),
.Y(n_1547)
);

AOI22xp33_ASAP7_75t_L g1548 ( 
.A1(n_1507),
.A2(n_1426),
.B1(n_1427),
.B2(n_1486),
.Y(n_1548)
);

AND2x2_ASAP7_75t_L g1549 ( 
.A(n_1503),
.B(n_1493),
.Y(n_1549)
);

AND2x2_ASAP7_75t_L g1550 ( 
.A(n_1503),
.B(n_1493),
.Y(n_1550)
);

NAND2x1p5_ASAP7_75t_L g1551 ( 
.A(n_1524),
.B(n_1495),
.Y(n_1551)
);

INVx1_ASAP7_75t_L g1552 ( 
.A(n_1534),
.Y(n_1552)
);

AND2x4_ASAP7_75t_SL g1553 ( 
.A(n_1535),
.B(n_1434),
.Y(n_1553)
);

NAND2xp5_ASAP7_75t_L g1554 ( 
.A(n_1508),
.B(n_1500),
.Y(n_1554)
);

NAND2xp5_ASAP7_75t_L g1555 ( 
.A(n_1508),
.B(n_1500),
.Y(n_1555)
);

AND2x4_ASAP7_75t_L g1556 ( 
.A(n_1532),
.B(n_1495),
.Y(n_1556)
);

AND2x4_ASAP7_75t_L g1557 ( 
.A(n_1532),
.B(n_1495),
.Y(n_1557)
);

INVx2_ASAP7_75t_L g1558 ( 
.A(n_1518),
.Y(n_1558)
);

OR2x2_ASAP7_75t_L g1559 ( 
.A(n_1518),
.B(n_1485),
.Y(n_1559)
);

INVx1_ASAP7_75t_SL g1560 ( 
.A(n_1536),
.Y(n_1560)
);

NAND3xp33_ASAP7_75t_L g1561 ( 
.A(n_1513),
.B(n_1449),
.C(n_1431),
.Y(n_1561)
);

HB1xp67_ASAP7_75t_L g1562 ( 
.A(n_1502),
.Y(n_1562)
);

AND2x2_ASAP7_75t_L g1563 ( 
.A(n_1521),
.B(n_1484),
.Y(n_1563)
);

INVx1_ASAP7_75t_L g1564 ( 
.A(n_1534),
.Y(n_1564)
);

AND2x2_ASAP7_75t_L g1565 ( 
.A(n_1521),
.B(n_1496),
.Y(n_1565)
);

AND2x2_ASAP7_75t_L g1566 ( 
.A(n_1521),
.B(n_1496),
.Y(n_1566)
);

OR2x2_ASAP7_75t_L g1567 ( 
.A(n_1526),
.B(n_1485),
.Y(n_1567)
);

NOR2xp33_ASAP7_75t_L g1568 ( 
.A(n_1530),
.B(n_1449),
.Y(n_1568)
);

INVx1_ASAP7_75t_L g1569 ( 
.A(n_1526),
.Y(n_1569)
);

AND2x2_ASAP7_75t_L g1570 ( 
.A(n_1522),
.B(n_1496),
.Y(n_1570)
);

INVx1_ASAP7_75t_L g1571 ( 
.A(n_1526),
.Y(n_1571)
);

INVxp67_ASAP7_75t_SL g1572 ( 
.A(n_1528),
.Y(n_1572)
);

OR2x2_ASAP7_75t_L g1573 ( 
.A(n_1512),
.B(n_1485),
.Y(n_1573)
);

BUFx2_ASAP7_75t_L g1574 ( 
.A(n_1532),
.Y(n_1574)
);

INVx2_ASAP7_75t_L g1575 ( 
.A(n_1542),
.Y(n_1575)
);

AND2x2_ASAP7_75t_L g1576 ( 
.A(n_1563),
.B(n_1515),
.Y(n_1576)
);

INVx1_ASAP7_75t_L g1577 ( 
.A(n_1541),
.Y(n_1577)
);

NAND2xp5_ASAP7_75t_L g1578 ( 
.A(n_1554),
.B(n_1528),
.Y(n_1578)
);

OR2x2_ASAP7_75t_L g1579 ( 
.A(n_1539),
.B(n_1506),
.Y(n_1579)
);

NOR2xp33_ASAP7_75t_L g1580 ( 
.A(n_1568),
.B(n_1561),
.Y(n_1580)
);

INVx2_ASAP7_75t_SL g1581 ( 
.A(n_1553),
.Y(n_1581)
);

AND2x2_ASAP7_75t_L g1582 ( 
.A(n_1563),
.B(n_1574),
.Y(n_1582)
);

INVx1_ASAP7_75t_L g1583 ( 
.A(n_1541),
.Y(n_1583)
);

OR2x2_ASAP7_75t_L g1584 ( 
.A(n_1539),
.B(n_1506),
.Y(n_1584)
);

NAND2xp5_ASAP7_75t_L g1585 ( 
.A(n_1554),
.B(n_1513),
.Y(n_1585)
);

AND2x2_ASAP7_75t_L g1586 ( 
.A(n_1563),
.B(n_1515),
.Y(n_1586)
);

HB1xp67_ASAP7_75t_L g1587 ( 
.A(n_1547),
.Y(n_1587)
);

INVx1_ASAP7_75t_SL g1588 ( 
.A(n_1547),
.Y(n_1588)
);

HB1xp67_ASAP7_75t_L g1589 ( 
.A(n_1560),
.Y(n_1589)
);

NAND2xp5_ASAP7_75t_L g1590 ( 
.A(n_1555),
.B(n_1530),
.Y(n_1590)
);

AND2x2_ASAP7_75t_L g1591 ( 
.A(n_1574),
.B(n_1515),
.Y(n_1591)
);

INVx1_ASAP7_75t_L g1592 ( 
.A(n_1544),
.Y(n_1592)
);

AO21x1_ASAP7_75t_L g1593 ( 
.A1(n_1568),
.A2(n_1572),
.B(n_1562),
.Y(n_1593)
);

INVx1_ASAP7_75t_L g1594 ( 
.A(n_1544),
.Y(n_1594)
);

NAND3xp33_ASAP7_75t_SL g1595 ( 
.A(n_1561),
.B(n_1507),
.C(n_1529),
.Y(n_1595)
);

INVxp67_ASAP7_75t_L g1596 ( 
.A(n_1560),
.Y(n_1596)
);

NOR2xp33_ASAP7_75t_SL g1597 ( 
.A(n_1572),
.B(n_1425),
.Y(n_1597)
);

INVx2_ASAP7_75t_SL g1598 ( 
.A(n_1553),
.Y(n_1598)
);

O2A1O1Ixp5_ASAP7_75t_L g1599 ( 
.A1(n_1537),
.A2(n_1505),
.B(n_1516),
.C(n_1509),
.Y(n_1599)
);

NAND2xp5_ASAP7_75t_L g1600 ( 
.A(n_1555),
.B(n_1529),
.Y(n_1600)
);

OR2x2_ASAP7_75t_L g1601 ( 
.A(n_1537),
.B(n_1506),
.Y(n_1601)
);

HB1xp67_ASAP7_75t_L g1602 ( 
.A(n_1562),
.Y(n_1602)
);

AND2x2_ASAP7_75t_L g1603 ( 
.A(n_1574),
.B(n_1511),
.Y(n_1603)
);

NOR2xp33_ASAP7_75t_L g1604 ( 
.A(n_1553),
.B(n_1464),
.Y(n_1604)
);

NAND2xp5_ASAP7_75t_L g1605 ( 
.A(n_1573),
.B(n_1509),
.Y(n_1605)
);

INVx1_ASAP7_75t_L g1606 ( 
.A(n_1552),
.Y(n_1606)
);

INVx2_ASAP7_75t_L g1607 ( 
.A(n_1542),
.Y(n_1607)
);

NAND2xp5_ASAP7_75t_L g1608 ( 
.A(n_1573),
.B(n_1511),
.Y(n_1608)
);

NAND2xp5_ASAP7_75t_L g1609 ( 
.A(n_1573),
.B(n_1511),
.Y(n_1609)
);

INVx1_ASAP7_75t_L g1610 ( 
.A(n_1552),
.Y(n_1610)
);

INVxp67_ASAP7_75t_L g1611 ( 
.A(n_1567),
.Y(n_1611)
);

NOR2xp33_ASAP7_75t_R g1612 ( 
.A(n_1548),
.B(n_1464),
.Y(n_1612)
);

OR2x2_ASAP7_75t_L g1613 ( 
.A(n_1567),
.B(n_1512),
.Y(n_1613)
);

INVx1_ASAP7_75t_L g1614 ( 
.A(n_1564),
.Y(n_1614)
);

NAND2xp33_ASAP7_75t_L g1615 ( 
.A(n_1548),
.B(n_1490),
.Y(n_1615)
);

INVx1_ASAP7_75t_L g1616 ( 
.A(n_1564),
.Y(n_1616)
);

NAND2xp5_ASAP7_75t_L g1617 ( 
.A(n_1585),
.B(n_1512),
.Y(n_1617)
);

AND2x2_ASAP7_75t_L g1618 ( 
.A(n_1581),
.B(n_1545),
.Y(n_1618)
);

NAND2xp5_ASAP7_75t_L g1619 ( 
.A(n_1600),
.B(n_1545),
.Y(n_1619)
);

INVx1_ASAP7_75t_L g1620 ( 
.A(n_1577),
.Y(n_1620)
);

INVx1_ASAP7_75t_L g1621 ( 
.A(n_1602),
.Y(n_1621)
);

INVxp67_ASAP7_75t_L g1622 ( 
.A(n_1587),
.Y(n_1622)
);

INVx1_ASAP7_75t_SL g1623 ( 
.A(n_1588),
.Y(n_1623)
);

INVx2_ASAP7_75t_L g1624 ( 
.A(n_1575),
.Y(n_1624)
);

OAI21xp5_ASAP7_75t_L g1625 ( 
.A1(n_1595),
.A2(n_1453),
.B(n_1533),
.Y(n_1625)
);

NOR2xp33_ASAP7_75t_L g1626 ( 
.A(n_1580),
.B(n_1445),
.Y(n_1626)
);

OR2x2_ASAP7_75t_L g1627 ( 
.A(n_1588),
.B(n_1567),
.Y(n_1627)
);

INVx1_ASAP7_75t_L g1628 ( 
.A(n_1577),
.Y(n_1628)
);

NAND2xp5_ASAP7_75t_L g1629 ( 
.A(n_1590),
.B(n_1545),
.Y(n_1629)
);

INVx1_ASAP7_75t_L g1630 ( 
.A(n_1583),
.Y(n_1630)
);

NOR2xp33_ASAP7_75t_L g1631 ( 
.A(n_1604),
.B(n_1423),
.Y(n_1631)
);

OR2x2_ASAP7_75t_L g1632 ( 
.A(n_1605),
.B(n_1559),
.Y(n_1632)
);

AND2x2_ASAP7_75t_L g1633 ( 
.A(n_1581),
.B(n_1549),
.Y(n_1633)
);

OR2x2_ASAP7_75t_L g1634 ( 
.A(n_1589),
.B(n_1578),
.Y(n_1634)
);

INVx1_ASAP7_75t_SL g1635 ( 
.A(n_1597),
.Y(n_1635)
);

AOI211x1_ASAP7_75t_L g1636 ( 
.A1(n_1593),
.A2(n_1505),
.B(n_1549),
.C(n_1550),
.Y(n_1636)
);

INVx1_ASAP7_75t_L g1637 ( 
.A(n_1583),
.Y(n_1637)
);

NAND2xp5_ASAP7_75t_L g1638 ( 
.A(n_1596),
.B(n_1611),
.Y(n_1638)
);

INVx1_ASAP7_75t_L g1639 ( 
.A(n_1592),
.Y(n_1639)
);

AND2x2_ASAP7_75t_L g1640 ( 
.A(n_1598),
.B(n_1549),
.Y(n_1640)
);

NAND4xp25_ASAP7_75t_L g1641 ( 
.A(n_1599),
.B(n_1533),
.C(n_1453),
.D(n_1486),
.Y(n_1641)
);

INVx2_ASAP7_75t_L g1642 ( 
.A(n_1575),
.Y(n_1642)
);

NAND2xp5_ASAP7_75t_L g1643 ( 
.A(n_1608),
.B(n_1609),
.Y(n_1643)
);

NAND2xp5_ASAP7_75t_L g1644 ( 
.A(n_1598),
.B(n_1550),
.Y(n_1644)
);

INVx1_ASAP7_75t_L g1645 ( 
.A(n_1592),
.Y(n_1645)
);

OR2x2_ASAP7_75t_L g1646 ( 
.A(n_1601),
.B(n_1559),
.Y(n_1646)
);

INVx2_ASAP7_75t_L g1647 ( 
.A(n_1607),
.Y(n_1647)
);

NOR2xp33_ASAP7_75t_L g1648 ( 
.A(n_1597),
.B(n_1553),
.Y(n_1648)
);

INVx2_ASAP7_75t_L g1649 ( 
.A(n_1607),
.Y(n_1649)
);

NOR2xp33_ASAP7_75t_L g1650 ( 
.A(n_1615),
.B(n_1497),
.Y(n_1650)
);

NOR2xp33_ASAP7_75t_L g1651 ( 
.A(n_1601),
.B(n_1497),
.Y(n_1651)
);

INVx1_ASAP7_75t_L g1652 ( 
.A(n_1620),
.Y(n_1652)
);

INVx1_ASAP7_75t_L g1653 ( 
.A(n_1620),
.Y(n_1653)
);

AOI22xp5_ASAP7_75t_L g1654 ( 
.A1(n_1641),
.A2(n_1593),
.B1(n_1505),
.B2(n_1582),
.Y(n_1654)
);

INVx1_ASAP7_75t_L g1655 ( 
.A(n_1628),
.Y(n_1655)
);

INVx1_ASAP7_75t_L g1656 ( 
.A(n_1628),
.Y(n_1656)
);

AOI221xp5_ASAP7_75t_L g1657 ( 
.A1(n_1636),
.A2(n_1612),
.B1(n_1582),
.B2(n_1616),
.C(n_1614),
.Y(n_1657)
);

AOI21xp33_ASAP7_75t_L g1658 ( 
.A1(n_1635),
.A2(n_1610),
.B(n_1606),
.Y(n_1658)
);

OAI21xp5_ASAP7_75t_L g1659 ( 
.A1(n_1625),
.A2(n_1610),
.B(n_1606),
.Y(n_1659)
);

OAI22xp5_ASAP7_75t_L g1660 ( 
.A1(n_1623),
.A2(n_1648),
.B1(n_1622),
.B2(n_1619),
.Y(n_1660)
);

AOI22xp5_ASAP7_75t_L g1661 ( 
.A1(n_1650),
.A2(n_1603),
.B1(n_1614),
.B2(n_1616),
.Y(n_1661)
);

INVxp67_ASAP7_75t_L g1662 ( 
.A(n_1626),
.Y(n_1662)
);

AND2x2_ASAP7_75t_L g1663 ( 
.A(n_1618),
.B(n_1576),
.Y(n_1663)
);

NOR2xp33_ASAP7_75t_L g1664 ( 
.A(n_1638),
.B(n_1579),
.Y(n_1664)
);

XNOR2x1_ASAP7_75t_L g1665 ( 
.A(n_1634),
.B(n_1490),
.Y(n_1665)
);

OAI322xp33_ASAP7_75t_L g1666 ( 
.A1(n_1634),
.A2(n_1584),
.A3(n_1579),
.B1(n_1613),
.B2(n_1594),
.C1(n_1559),
.C2(n_1551),
.Y(n_1666)
);

OAI21xp5_ASAP7_75t_L g1667 ( 
.A1(n_1621),
.A2(n_1594),
.B(n_1603),
.Y(n_1667)
);

INVx1_ASAP7_75t_L g1668 ( 
.A(n_1630),
.Y(n_1668)
);

INVx1_ASAP7_75t_L g1669 ( 
.A(n_1630),
.Y(n_1669)
);

AND2x2_ASAP7_75t_L g1670 ( 
.A(n_1618),
.B(n_1576),
.Y(n_1670)
);

AND2x2_ASAP7_75t_L g1671 ( 
.A(n_1633),
.B(n_1586),
.Y(n_1671)
);

AOI222xp33_ASAP7_75t_L g1672 ( 
.A1(n_1617),
.A2(n_1550),
.B1(n_1591),
.B2(n_1586),
.C1(n_1540),
.C2(n_1538),
.Y(n_1672)
);

AND2x2_ASAP7_75t_L g1673 ( 
.A(n_1633),
.B(n_1591),
.Y(n_1673)
);

INVx1_ASAP7_75t_L g1674 ( 
.A(n_1637),
.Y(n_1674)
);

NAND2x1_ASAP7_75t_SL g1675 ( 
.A(n_1640),
.B(n_1556),
.Y(n_1675)
);

INVxp67_ASAP7_75t_L g1676 ( 
.A(n_1631),
.Y(n_1676)
);

NAND2x1_ASAP7_75t_L g1677 ( 
.A(n_1673),
.B(n_1640),
.Y(n_1677)
);

AOI22xp5_ASAP7_75t_L g1678 ( 
.A1(n_1654),
.A2(n_1644),
.B1(n_1629),
.B2(n_1651),
.Y(n_1678)
);

NOR2x1_ASAP7_75t_L g1679 ( 
.A(n_1659),
.B(n_1637),
.Y(n_1679)
);

INVx2_ASAP7_75t_SL g1680 ( 
.A(n_1675),
.Y(n_1680)
);

NAND3xp33_ASAP7_75t_SL g1681 ( 
.A(n_1657),
.B(n_1660),
.C(n_1667),
.Y(n_1681)
);

AOI22xp33_ASAP7_75t_L g1682 ( 
.A1(n_1664),
.A2(n_1643),
.B1(n_1632),
.B2(n_1627),
.Y(n_1682)
);

INVx1_ASAP7_75t_L g1683 ( 
.A(n_1652),
.Y(n_1683)
);

AOI32xp33_ASAP7_75t_L g1684 ( 
.A1(n_1665),
.A2(n_1627),
.A3(n_1645),
.B1(n_1639),
.B2(n_1557),
.Y(n_1684)
);

NOR3xp33_ASAP7_75t_L g1685 ( 
.A(n_1658),
.B(n_1645),
.C(n_1639),
.Y(n_1685)
);

INVx1_ASAP7_75t_L g1686 ( 
.A(n_1653),
.Y(n_1686)
);

XOR2x2_ASAP7_75t_L g1687 ( 
.A(n_1665),
.B(n_1444),
.Y(n_1687)
);

NOR2xp33_ASAP7_75t_L g1688 ( 
.A(n_1662),
.B(n_1632),
.Y(n_1688)
);

O2A1O1Ixp5_ASAP7_75t_L g1689 ( 
.A1(n_1666),
.A2(n_1646),
.B(n_1647),
.C(n_1649),
.Y(n_1689)
);

OAI33xp33_ASAP7_75t_L g1690 ( 
.A1(n_1655),
.A2(n_1646),
.A3(n_1642),
.B1(n_1649),
.B2(n_1647),
.B3(n_1624),
.Y(n_1690)
);

AND2x2_ASAP7_75t_L g1691 ( 
.A(n_1673),
.B(n_1565),
.Y(n_1691)
);

OAI22xp5_ASAP7_75t_L g1692 ( 
.A1(n_1676),
.A2(n_1584),
.B1(n_1551),
.B2(n_1451),
.Y(n_1692)
);

AOI21xp33_ASAP7_75t_SL g1693 ( 
.A1(n_1664),
.A2(n_1510),
.B(n_1551),
.Y(n_1693)
);

NAND2xp5_ASAP7_75t_SL g1694 ( 
.A(n_1661),
.B(n_1613),
.Y(n_1694)
);

OR2x2_ASAP7_75t_L g1695 ( 
.A(n_1663),
.B(n_1624),
.Y(n_1695)
);

NAND2xp5_ASAP7_75t_L g1696 ( 
.A(n_1688),
.B(n_1663),
.Y(n_1696)
);

XOR2x2_ASAP7_75t_L g1697 ( 
.A(n_1681),
.B(n_1670),
.Y(n_1697)
);

NOR2xp33_ASAP7_75t_L g1698 ( 
.A(n_1678),
.B(n_1694),
.Y(n_1698)
);

AOI21xp5_ASAP7_75t_L g1699 ( 
.A1(n_1679),
.A2(n_1668),
.B(n_1656),
.Y(n_1699)
);

OR2x2_ASAP7_75t_L g1700 ( 
.A(n_1695),
.B(n_1670),
.Y(n_1700)
);

NAND2xp5_ASAP7_75t_SL g1701 ( 
.A(n_1680),
.B(n_1672),
.Y(n_1701)
);

INVxp67_ASAP7_75t_L g1702 ( 
.A(n_1677),
.Y(n_1702)
);

OAI21xp5_ASAP7_75t_SL g1703 ( 
.A1(n_1684),
.A2(n_1671),
.B(n_1669),
.Y(n_1703)
);

AOI21xp5_ASAP7_75t_SL g1704 ( 
.A1(n_1692),
.A2(n_1674),
.B(n_1671),
.Y(n_1704)
);

OAI22xp5_ASAP7_75t_L g1705 ( 
.A1(n_1682),
.A2(n_1551),
.B1(n_1556),
.B2(n_1557),
.Y(n_1705)
);

AOI322xp5_ASAP7_75t_L g1706 ( 
.A1(n_1685),
.A2(n_1540),
.A3(n_1543),
.B1(n_1538),
.B2(n_1556),
.C1(n_1557),
.C2(n_1520),
.Y(n_1706)
);

NAND3xp33_ASAP7_75t_L g1707 ( 
.A(n_1698),
.B(n_1689),
.C(n_1686),
.Y(n_1707)
);

AND2x2_ASAP7_75t_L g1708 ( 
.A(n_1702),
.B(n_1687),
.Y(n_1708)
);

INVx1_ASAP7_75t_L g1709 ( 
.A(n_1700),
.Y(n_1709)
);

INVxp67_ASAP7_75t_L g1710 ( 
.A(n_1696),
.Y(n_1710)
);

OAI22xp5_ASAP7_75t_L g1711 ( 
.A1(n_1701),
.A2(n_1692),
.B1(n_1693),
.B2(n_1691),
.Y(n_1711)
);

NOR2xp33_ASAP7_75t_L g1712 ( 
.A(n_1703),
.B(n_1690),
.Y(n_1712)
);

NAND4xp25_ASAP7_75t_L g1713 ( 
.A(n_1699),
.B(n_1683),
.C(n_1642),
.D(n_1557),
.Y(n_1713)
);

NAND4xp75_ASAP7_75t_L g1714 ( 
.A(n_1697),
.B(n_1538),
.C(n_1540),
.D(n_1543),
.Y(n_1714)
);

NAND2xp5_ASAP7_75t_L g1715 ( 
.A(n_1704),
.B(n_1569),
.Y(n_1715)
);

NAND2xp5_ASAP7_75t_L g1716 ( 
.A(n_1706),
.B(n_1569),
.Y(n_1716)
);

OAI22xp5_ASAP7_75t_L g1717 ( 
.A1(n_1705),
.A2(n_1551),
.B1(n_1556),
.B2(n_1557),
.Y(n_1717)
);

AOI22xp5_ASAP7_75t_L g1718 ( 
.A1(n_1712),
.A2(n_1557),
.B1(n_1556),
.B2(n_1532),
.Y(n_1718)
);

AOI221xp5_ASAP7_75t_L g1719 ( 
.A1(n_1707),
.A2(n_1510),
.B1(n_1457),
.B2(n_1556),
.C(n_1524),
.Y(n_1719)
);

AOI221xp5_ASAP7_75t_L g1720 ( 
.A1(n_1711),
.A2(n_1510),
.B1(n_1524),
.B2(n_1523),
.C(n_1517),
.Y(n_1720)
);

NAND4xp75_ASAP7_75t_L g1721 ( 
.A(n_1709),
.B(n_1543),
.C(n_1523),
.D(n_1517),
.Y(n_1721)
);

NAND2xp5_ASAP7_75t_L g1722 ( 
.A(n_1708),
.B(n_1569),
.Y(n_1722)
);

NOR2x1_ASAP7_75t_L g1723 ( 
.A(n_1714),
.B(n_1542),
.Y(n_1723)
);

AOI21xp33_ASAP7_75t_SL g1724 ( 
.A1(n_1722),
.A2(n_1710),
.B(n_1715),
.Y(n_1724)
);

NAND2xp5_ASAP7_75t_L g1725 ( 
.A(n_1718),
.B(n_1713),
.Y(n_1725)
);

OAI221xp5_ASAP7_75t_L g1726 ( 
.A1(n_1720),
.A2(n_1716),
.B1(n_1717),
.B2(n_1524),
.C(n_1571),
.Y(n_1726)
);

OAI22xp5_ASAP7_75t_L g1727 ( 
.A1(n_1719),
.A2(n_1571),
.B1(n_1524),
.B2(n_1542),
.Y(n_1727)
);

HB1xp67_ASAP7_75t_L g1728 ( 
.A(n_1723),
.Y(n_1728)
);

AOI22xp33_ASAP7_75t_L g1729 ( 
.A1(n_1721),
.A2(n_1474),
.B1(n_1441),
.B2(n_1532),
.Y(n_1729)
);

NAND2xp5_ASAP7_75t_L g1730 ( 
.A(n_1724),
.B(n_1571),
.Y(n_1730)
);

INVx2_ASAP7_75t_L g1731 ( 
.A(n_1728),
.Y(n_1731)
);

NOR2xp33_ASAP7_75t_L g1732 ( 
.A(n_1725),
.B(n_1546),
.Y(n_1732)
);

NOR2xp33_ASAP7_75t_L g1733 ( 
.A(n_1726),
.B(n_1546),
.Y(n_1733)
);

NAND2xp5_ASAP7_75t_L g1734 ( 
.A(n_1727),
.B(n_1546),
.Y(n_1734)
);

AOI22x1_ASAP7_75t_L g1735 ( 
.A1(n_1731),
.A2(n_1729),
.B1(n_1546),
.B2(n_1558),
.Y(n_1735)
);

O2A1O1Ixp33_ASAP7_75t_L g1736 ( 
.A1(n_1730),
.A2(n_1558),
.B(n_1504),
.C(n_1502),
.Y(n_1736)
);

NOR2x1p5_ASAP7_75t_L g1737 ( 
.A(n_1734),
.B(n_1402),
.Y(n_1737)
);

OAI222xp33_ASAP7_75t_L g1738 ( 
.A1(n_1735),
.A2(n_1733),
.B1(n_1732),
.B2(n_1532),
.C1(n_1558),
.C2(n_1504),
.Y(n_1738)
);

AOI22x1_ASAP7_75t_L g1739 ( 
.A1(n_1738),
.A2(n_1737),
.B1(n_1736),
.B2(n_1558),
.Y(n_1739)
);

OAI22xp5_ASAP7_75t_L g1740 ( 
.A1(n_1739),
.A2(n_1520),
.B1(n_1527),
.B2(n_1532),
.Y(n_1740)
);

OAI22xp5_ASAP7_75t_SL g1741 ( 
.A1(n_1739),
.A2(n_1389),
.B1(n_1434),
.B2(n_1402),
.Y(n_1741)
);

AOI22x1_ASAP7_75t_L g1742 ( 
.A1(n_1741),
.A2(n_1527),
.B1(n_1442),
.B2(n_1419),
.Y(n_1742)
);

INVx1_ASAP7_75t_L g1743 ( 
.A(n_1740),
.Y(n_1743)
);

AOI22xp5_ASAP7_75t_L g1744 ( 
.A1(n_1743),
.A2(n_1570),
.B1(n_1566),
.B2(n_1565),
.Y(n_1744)
);

INVx1_ASAP7_75t_L g1745 ( 
.A(n_1742),
.Y(n_1745)
);

AOI21xp5_ASAP7_75t_L g1746 ( 
.A1(n_1745),
.A2(n_1451),
.B(n_1408),
.Y(n_1746)
);

OAI22xp5_ASAP7_75t_L g1747 ( 
.A1(n_1746),
.A2(n_1744),
.B1(n_1570),
.B2(n_1566),
.Y(n_1747)
);

INVx1_ASAP7_75t_L g1748 ( 
.A(n_1747),
.Y(n_1748)
);

OAI221xp5_ASAP7_75t_L g1749 ( 
.A1(n_1748),
.A2(n_1402),
.B1(n_1419),
.B2(n_1468),
.C(n_1531),
.Y(n_1749)
);

AOI211xp5_ASAP7_75t_L g1750 ( 
.A1(n_1749),
.A2(n_1442),
.B(n_1516),
.C(n_1468),
.Y(n_1750)
);


endmodule