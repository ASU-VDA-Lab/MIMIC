module fake_jpeg_12784_n_531 (n_13, n_11, n_14, n_17, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_531);

input n_13;
input n_11;
input n_14;
input n_17;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_531;

wire n_529;
wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_525;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_519;
wire n_276;
wire n_143;
wire n_431;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_513;
wire n_283;
wire n_107;
wire n_490;
wire n_517;
wire n_415;
wire n_479;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_48;
wire n_465;
wire n_200;
wire n_265;
wire n_192;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_221;
wire n_256;
wire n_454;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_508;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_530;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_474;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_511;
wire n_305;
wire n_161;
wire n_441;
wire n_342;
wire n_101;
wire n_226;
wire n_509;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_510;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_523;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_296;
wire n_384;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_491;
wire n_24;
wire n_526;
wire n_467;
wire n_269;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_473;
wire n_45;
wire n_520;
wire n_476;
wire n_337;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_344;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_481;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_522;
wire n_333;
wire n_518;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_302;
wire n_216;
wire n_528;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_199;
wire n_260;
wire n_413;
wire n_275;
wire n_494;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_492;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_515;
wire n_347;
wire n_521;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_472;
wire n_279;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_484;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_469;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_527;
wire n_482;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_512;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_516;
wire n_183;
wire n_409;
wire n_249;
wire n_412;
wire n_217;
wire n_471;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_524;
wire n_402;
wire n_504;
wire n_438;
wire n_475;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_514;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_10),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_15),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_13),
.Y(n_20)
);

BUFx4f_ASAP7_75t_L g21 ( 
.A(n_3),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_11),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_17),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_17),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_15),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_0),
.Y(n_26)
);

CKINVDCx16_ASAP7_75t_R g27 ( 
.A(n_13),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_12),
.Y(n_28)
);

INVx2_ASAP7_75t_SL g29 ( 
.A(n_1),
.Y(n_29)
);

BUFx3_ASAP7_75t_L g30 ( 
.A(n_16),
.Y(n_30)
);

BUFx16f_ASAP7_75t_L g31 ( 
.A(n_13),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_6),
.Y(n_32)
);

BUFx3_ASAP7_75t_L g33 ( 
.A(n_9),
.Y(n_33)
);

BUFx10_ASAP7_75t_L g34 ( 
.A(n_12),
.Y(n_34)
);

BUFx3_ASAP7_75t_L g35 ( 
.A(n_11),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_15),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_6),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_11),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_14),
.Y(n_39)
);

INVx11_ASAP7_75t_SL g40 ( 
.A(n_2),
.Y(n_40)
);

INVx8_ASAP7_75t_L g41 ( 
.A(n_5),
.Y(n_41)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_4),
.Y(n_42)
);

BUFx5_ASAP7_75t_L g43 ( 
.A(n_14),
.Y(n_43)
);

INVx11_ASAP7_75t_L g44 ( 
.A(n_16),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_7),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_8),
.Y(n_46)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_11),
.Y(n_47)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_10),
.Y(n_48)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_5),
.Y(n_49)
);

BUFx12f_ASAP7_75t_L g50 ( 
.A(n_16),
.Y(n_50)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_3),
.Y(n_51)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_12),
.Y(n_52)
);

BUFx12f_ASAP7_75t_L g53 ( 
.A(n_5),
.Y(n_53)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_4),
.Y(n_54)
);

BUFx12f_ASAP7_75t_L g55 ( 
.A(n_0),
.Y(n_55)
);

BUFx5_ASAP7_75t_L g56 ( 
.A(n_8),
.Y(n_56)
);

CKINVDCx20_ASAP7_75t_R g57 ( 
.A(n_4),
.Y(n_57)
);

CKINVDCx20_ASAP7_75t_R g58 ( 
.A(n_4),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_SL g59 ( 
.A(n_19),
.B(n_17),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_L g148 ( 
.A(n_59),
.B(n_61),
.Y(n_148)
);

BUFx3_ASAP7_75t_L g60 ( 
.A(n_56),
.Y(n_60)
);

INVx5_ASAP7_75t_L g123 ( 
.A(n_60),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_SL g61 ( 
.A(n_19),
.B(n_14),
.Y(n_61)
);

BUFx3_ASAP7_75t_L g62 ( 
.A(n_56),
.Y(n_62)
);

INVx5_ASAP7_75t_L g158 ( 
.A(n_62),
.Y(n_158)
);

INVx5_ASAP7_75t_SL g63 ( 
.A(n_34),
.Y(n_63)
);

INVx1_ASAP7_75t_SL g134 ( 
.A(n_63),
.Y(n_134)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_36),
.Y(n_64)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_64),
.Y(n_124)
);

OR2x2_ASAP7_75t_L g65 ( 
.A(n_36),
.B(n_0),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g137 ( 
.A(n_65),
.B(n_82),
.Y(n_137)
);

INVx3_ASAP7_75t_L g66 ( 
.A(n_43),
.Y(n_66)
);

INVx3_ASAP7_75t_L g175 ( 
.A(n_66),
.Y(n_175)
);

INVx11_ASAP7_75t_L g67 ( 
.A(n_34),
.Y(n_67)
);

INVx8_ASAP7_75t_L g193 ( 
.A(n_67),
.Y(n_193)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_22),
.Y(n_68)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_68),
.Y(n_131)
);

INVx3_ASAP7_75t_L g69 ( 
.A(n_31),
.Y(n_69)
);

INVx3_ASAP7_75t_L g200 ( 
.A(n_69),
.Y(n_200)
);

INVx3_ASAP7_75t_L g70 ( 
.A(n_43),
.Y(n_70)
);

INVx2_ASAP7_75t_SL g190 ( 
.A(n_70),
.Y(n_190)
);

NAND2xp5_ASAP7_75t_L g71 ( 
.A(n_24),
.B(n_0),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_L g169 ( 
.A(n_71),
.B(n_81),
.Y(n_169)
);

INVx11_ASAP7_75t_L g72 ( 
.A(n_34),
.Y(n_72)
);

INVx5_ASAP7_75t_L g160 ( 
.A(n_72),
.Y(n_160)
);

INVx2_ASAP7_75t_L g73 ( 
.A(n_21),
.Y(n_73)
);

INVx2_ASAP7_75t_L g142 ( 
.A(n_73),
.Y(n_142)
);

BUFx6f_ASAP7_75t_L g74 ( 
.A(n_38),
.Y(n_74)
);

BUFx6f_ASAP7_75t_L g133 ( 
.A(n_74),
.Y(n_133)
);

INVx6_ASAP7_75t_L g75 ( 
.A(n_38),
.Y(n_75)
);

BUFx6f_ASAP7_75t_L g157 ( 
.A(n_75),
.Y(n_157)
);

INVx8_ASAP7_75t_L g76 ( 
.A(n_56),
.Y(n_76)
);

INVx5_ASAP7_75t_L g167 ( 
.A(n_76),
.Y(n_167)
);

INVx3_ASAP7_75t_L g77 ( 
.A(n_31),
.Y(n_77)
);

INVx4_ASAP7_75t_L g144 ( 
.A(n_77),
.Y(n_144)
);

BUFx6f_ASAP7_75t_L g78 ( 
.A(n_38),
.Y(n_78)
);

BUFx6f_ASAP7_75t_L g165 ( 
.A(n_78),
.Y(n_165)
);

AND2x2_ASAP7_75t_L g79 ( 
.A(n_50),
.B(n_1),
.Y(n_79)
);

AND2x2_ASAP7_75t_L g125 ( 
.A(n_79),
.B(n_89),
.Y(n_125)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_22),
.Y(n_80)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_80),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_L g81 ( 
.A(n_24),
.B(n_13),
.Y(n_81)
);

CKINVDCx20_ASAP7_75t_R g82 ( 
.A(n_44),
.Y(n_82)
);

INVx2_ASAP7_75t_L g83 ( 
.A(n_21),
.Y(n_83)
);

INVx2_ASAP7_75t_L g154 ( 
.A(n_83),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_L g84 ( 
.A(n_25),
.B(n_1),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g188 ( 
.A(n_84),
.B(n_85),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_L g85 ( 
.A(n_25),
.B(n_1),
.Y(n_85)
);

INVx3_ASAP7_75t_L g86 ( 
.A(n_43),
.Y(n_86)
);

INVx4_ASAP7_75t_L g173 ( 
.A(n_86),
.Y(n_173)
);

BUFx5_ASAP7_75t_L g87 ( 
.A(n_44),
.Y(n_87)
);

BUFx4f_ASAP7_75t_SL g174 ( 
.A(n_87),
.Y(n_174)
);

BUFx6f_ASAP7_75t_L g88 ( 
.A(n_38),
.Y(n_88)
);

BUFx6f_ASAP7_75t_L g185 ( 
.A(n_88),
.Y(n_185)
);

AND2x2_ASAP7_75t_L g89 ( 
.A(n_50),
.B(n_30),
.Y(n_89)
);

CKINVDCx20_ASAP7_75t_R g90 ( 
.A(n_44),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g150 ( 
.A(n_90),
.B(n_94),
.Y(n_150)
);

INVx6_ASAP7_75t_L g91 ( 
.A(n_45),
.Y(n_91)
);

INVx6_ASAP7_75t_L g136 ( 
.A(n_91),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_39),
.B(n_2),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_SL g128 ( 
.A(n_92),
.B(n_113),
.Y(n_128)
);

BUFx6f_ASAP7_75t_L g93 ( 
.A(n_45),
.Y(n_93)
);

INVx6_ASAP7_75t_L g143 ( 
.A(n_93),
.Y(n_143)
);

CKINVDCx20_ASAP7_75t_R g94 ( 
.A(n_34),
.Y(n_94)
);

BUFx12f_ASAP7_75t_L g95 ( 
.A(n_33),
.Y(n_95)
);

INVx5_ASAP7_75t_L g178 ( 
.A(n_95),
.Y(n_178)
);

BUFx6f_ASAP7_75t_L g96 ( 
.A(n_45),
.Y(n_96)
);

INVx6_ASAP7_75t_L g182 ( 
.A(n_96),
.Y(n_182)
);

INVx3_ASAP7_75t_L g97 ( 
.A(n_31),
.Y(n_97)
);

BUFx2_ASAP7_75t_L g130 ( 
.A(n_97),
.Y(n_130)
);

BUFx4f_ASAP7_75t_SL g98 ( 
.A(n_34),
.Y(n_98)
);

BUFx4f_ASAP7_75t_SL g177 ( 
.A(n_98),
.Y(n_177)
);

INVx3_ASAP7_75t_L g99 ( 
.A(n_31),
.Y(n_99)
);

BUFx2_ASAP7_75t_L g138 ( 
.A(n_99),
.Y(n_138)
);

BUFx6f_ASAP7_75t_L g100 ( 
.A(n_21),
.Y(n_100)
);

BUFx2_ASAP7_75t_L g187 ( 
.A(n_100),
.Y(n_187)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_28),
.Y(n_101)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_101),
.Y(n_151)
);

INVx2_ASAP7_75t_L g102 ( 
.A(n_21),
.Y(n_102)
);

INVx2_ASAP7_75t_L g164 ( 
.A(n_102),
.Y(n_164)
);

INVx8_ASAP7_75t_L g103 ( 
.A(n_23),
.Y(n_103)
);

INVx5_ASAP7_75t_L g199 ( 
.A(n_103),
.Y(n_199)
);

INVx2_ASAP7_75t_L g104 ( 
.A(n_50),
.Y(n_104)
);

INVx2_ASAP7_75t_L g170 ( 
.A(n_104),
.Y(n_170)
);

BUFx3_ASAP7_75t_L g105 ( 
.A(n_53),
.Y(n_105)
);

INVx5_ASAP7_75t_L g192 ( 
.A(n_105),
.Y(n_192)
);

INVx4_ASAP7_75t_L g106 ( 
.A(n_53),
.Y(n_106)
);

INVx2_ASAP7_75t_L g180 ( 
.A(n_106),
.Y(n_180)
);

INVx8_ASAP7_75t_L g107 ( 
.A(n_23),
.Y(n_107)
);

INVx2_ASAP7_75t_L g186 ( 
.A(n_107),
.Y(n_186)
);

INVx3_ASAP7_75t_L g108 ( 
.A(n_50),
.Y(n_108)
);

INVx2_ASAP7_75t_L g189 ( 
.A(n_108),
.Y(n_189)
);

OR2x2_ASAP7_75t_SL g109 ( 
.A(n_27),
.B(n_12),
.Y(n_109)
);

OR2x2_ASAP7_75t_L g147 ( 
.A(n_109),
.B(n_42),
.Y(n_147)
);

INVx11_ASAP7_75t_SL g110 ( 
.A(n_40),
.Y(n_110)
);

BUFx4f_ASAP7_75t_SL g172 ( 
.A(n_110),
.Y(n_172)
);

BUFx6f_ASAP7_75t_L g111 ( 
.A(n_41),
.Y(n_111)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_111),
.Y(n_152)
);

BUFx3_ASAP7_75t_L g112 ( 
.A(n_53),
.Y(n_112)
);

AND2x2_ASAP7_75t_L g126 ( 
.A(n_112),
.B(n_115),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_L g113 ( 
.A(n_39),
.B(n_2),
.Y(n_113)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_28),
.Y(n_114)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_114),
.Y(n_184)
);

INVx3_ASAP7_75t_L g115 ( 
.A(n_50),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_L g116 ( 
.A(n_30),
.B(n_2),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_SL g163 ( 
.A(n_116),
.B(n_20),
.Y(n_163)
);

BUFx4f_ASAP7_75t_SL g117 ( 
.A(n_40),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_L g155 ( 
.A(n_117),
.B(n_118),
.Y(n_155)
);

CKINVDCx20_ASAP7_75t_R g118 ( 
.A(n_30),
.Y(n_118)
);

INVx3_ASAP7_75t_SL g119 ( 
.A(n_41),
.Y(n_119)
);

AND2x2_ASAP7_75t_L g127 ( 
.A(n_119),
.B(n_120),
.Y(n_127)
);

INVx2_ASAP7_75t_L g120 ( 
.A(n_53),
.Y(n_120)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_42),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_L g166 ( 
.A(n_121),
.B(n_18),
.Y(n_166)
);

BUFx8_ASAP7_75t_L g122 ( 
.A(n_27),
.Y(n_122)
);

AND2x2_ASAP7_75t_L g132 ( 
.A(n_122),
.B(n_55),
.Y(n_132)
);

AOI22xp5_ASAP7_75t_L g129 ( 
.A1(n_79),
.A2(n_23),
.B1(n_41),
.B2(n_33),
.Y(n_129)
);

OAI22xp5_ASAP7_75t_L g233 ( 
.A1(n_129),
.A2(n_135),
.B1(n_140),
.B2(n_141),
.Y(n_233)
);

AND2x2_ASAP7_75t_L g201 ( 
.A(n_132),
.B(n_162),
.Y(n_201)
);

AOI22xp33_ASAP7_75t_SL g135 ( 
.A1(n_119),
.A2(n_29),
.B1(n_35),
.B2(n_33),
.Y(n_135)
);

OAI22xp5_ASAP7_75t_SL g139 ( 
.A1(n_65),
.A2(n_35),
.B1(n_58),
.B2(n_47),
.Y(n_139)
);

AOI22xp5_ASAP7_75t_SL g244 ( 
.A1(n_139),
.A2(n_153),
.B1(n_176),
.B2(n_148),
.Y(n_244)
);

AOI22xp33_ASAP7_75t_SL g140 ( 
.A1(n_63),
.A2(n_29),
.B1(n_35),
.B2(n_53),
.Y(n_140)
);

AOI22xp33_ASAP7_75t_SL g141 ( 
.A1(n_76),
.A2(n_29),
.B1(n_55),
.B2(n_49),
.Y(n_141)
);

AOI22xp33_ASAP7_75t_SL g145 ( 
.A1(n_60),
.A2(n_29),
.B1(n_55),
.B2(n_49),
.Y(n_145)
);

OAI22xp5_ASAP7_75t_L g256 ( 
.A1(n_145),
.A2(n_146),
.B1(n_156),
.B2(n_159),
.Y(n_256)
);

AOI22xp33_ASAP7_75t_SL g146 ( 
.A1(n_62),
.A2(n_111),
.B1(n_109),
.B2(n_107),
.Y(n_146)
);

OR2x2_ASAP7_75t_SL g215 ( 
.A(n_147),
.B(n_128),
.Y(n_215)
);

OAI22xp5_ASAP7_75t_SL g153 ( 
.A1(n_91),
.A2(n_32),
.B1(n_57),
.B2(n_52),
.Y(n_153)
);

AOI22xp33_ASAP7_75t_L g156 ( 
.A1(n_93),
.A2(n_54),
.B1(n_48),
.B2(n_58),
.Y(n_156)
);

AOI22xp33_ASAP7_75t_L g159 ( 
.A1(n_96),
.A2(n_54),
.B1(n_48),
.B2(n_57),
.Y(n_159)
);

AOI22xp33_ASAP7_75t_L g161 ( 
.A1(n_75),
.A2(n_20),
.B1(n_52),
.B2(n_51),
.Y(n_161)
);

OAI22xp5_ASAP7_75t_SL g239 ( 
.A1(n_161),
.A2(n_9),
.B1(n_10),
.B2(n_181),
.Y(n_239)
);

AND2x2_ASAP7_75t_SL g162 ( 
.A(n_122),
.B(n_55),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_SL g202 ( 
.A(n_163),
.B(n_195),
.Y(n_202)
);

NOR2xp33_ASAP7_75t_L g231 ( 
.A(n_166),
.B(n_198),
.Y(n_231)
);

AOI21xp5_ASAP7_75t_L g168 ( 
.A1(n_89),
.A2(n_18),
.B(n_51),
.Y(n_168)
);

MAJIxp5_ASAP7_75t_L g206 ( 
.A(n_168),
.B(n_179),
.C(n_117),
.Y(n_206)
);

NOR2xp33_ASAP7_75t_L g171 ( 
.A(n_69),
.B(n_46),
.Y(n_171)
);

NOR2xp33_ASAP7_75t_SL g229 ( 
.A(n_171),
.B(n_194),
.Y(n_229)
);

AND2x2_ASAP7_75t_SL g176 ( 
.A(n_122),
.B(n_55),
.Y(n_176)
);

AND2x2_ASAP7_75t_L g258 ( 
.A(n_176),
.B(n_123),
.Y(n_258)
);

MAJIxp5_ASAP7_75t_L g179 ( 
.A(n_115),
.B(n_47),
.C(n_46),
.Y(n_179)
);

AOI22xp33_ASAP7_75t_SL g181 ( 
.A1(n_103),
.A2(n_37),
.B1(n_32),
.B2(n_26),
.Y(n_181)
);

AOI22xp33_ASAP7_75t_SL g216 ( 
.A1(n_181),
.A2(n_183),
.B1(n_191),
.B2(n_95),
.Y(n_216)
);

AOI22xp33_ASAP7_75t_SL g183 ( 
.A1(n_77),
.A2(n_37),
.B1(n_26),
.B2(n_6),
.Y(n_183)
);

AOI22xp33_ASAP7_75t_SL g191 ( 
.A1(n_67),
.A2(n_72),
.B1(n_106),
.B2(n_112),
.Y(n_191)
);

CKINVDCx20_ASAP7_75t_R g194 ( 
.A(n_110),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_L g195 ( 
.A(n_100),
.B(n_3),
.Y(n_195)
);

AND2x2_ASAP7_75t_L g196 ( 
.A(n_105),
.B(n_10),
.Y(n_196)
);

CKINVDCx14_ASAP7_75t_R g217 ( 
.A(n_196),
.Y(n_217)
);

NOR2xp33_ASAP7_75t_L g197 ( 
.A(n_98),
.B(n_3),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_SL g213 ( 
.A(n_197),
.B(n_5),
.Y(n_213)
);

CKINVDCx20_ASAP7_75t_R g198 ( 
.A(n_117),
.Y(n_198)
);

INVx2_ASAP7_75t_L g203 ( 
.A(n_142),
.Y(n_203)
);

INVx2_ASAP7_75t_L g282 ( 
.A(n_203),
.Y(n_282)
);

INVx4_ASAP7_75t_L g204 ( 
.A(n_178),
.Y(n_204)
);

BUFx2_ASAP7_75t_L g290 ( 
.A(n_204),
.Y(n_290)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_154),
.Y(n_205)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_205),
.Y(n_280)
);

AND2x2_ASAP7_75t_L g300 ( 
.A(n_206),
.B(n_220),
.Y(n_300)
);

AOI22xp33_ASAP7_75t_L g207 ( 
.A1(n_161),
.A2(n_156),
.B1(n_159),
.B2(n_88),
.Y(n_207)
);

OAI22xp5_ASAP7_75t_SL g273 ( 
.A1(n_207),
.A2(n_250),
.B1(n_165),
.B2(n_185),
.Y(n_273)
);

INVx2_ASAP7_75t_SL g208 ( 
.A(n_199),
.Y(n_208)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_208),
.Y(n_281)
);

CKINVDCx20_ASAP7_75t_R g209 ( 
.A(n_150),
.Y(n_209)
);

NOR2xp33_ASAP7_75t_L g271 ( 
.A(n_209),
.B(n_213),
.Y(n_271)
);

NAND2xp5_ASAP7_75t_L g210 ( 
.A(n_169),
.B(n_188),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_L g277 ( 
.A(n_210),
.B(n_236),
.Y(n_277)
);

CKINVDCx16_ASAP7_75t_R g211 ( 
.A(n_162),
.Y(n_211)
);

NOR2xp33_ASAP7_75t_L g268 ( 
.A(n_211),
.B(n_215),
.Y(n_268)
);

BUFx6f_ASAP7_75t_L g212 ( 
.A(n_133),
.Y(n_212)
);

BUFx6f_ASAP7_75t_L g270 ( 
.A(n_212),
.Y(n_270)
);

INVx2_ASAP7_75t_L g214 ( 
.A(n_164),
.Y(n_214)
);

INVx2_ASAP7_75t_L g294 ( 
.A(n_214),
.Y(n_294)
);

INVxp67_ASAP7_75t_L g291 ( 
.A(n_216),
.Y(n_291)
);

BUFx3_ASAP7_75t_L g218 ( 
.A(n_130),
.Y(n_218)
);

INVx3_ASAP7_75t_L g297 ( 
.A(n_218),
.Y(n_297)
);

INVx4_ASAP7_75t_L g219 ( 
.A(n_178),
.Y(n_219)
);

BUFx2_ASAP7_75t_L g306 ( 
.A(n_219),
.Y(n_306)
);

INVx1_ASAP7_75t_SL g220 ( 
.A(n_134),
.Y(n_220)
);

AOI22xp33_ASAP7_75t_SL g221 ( 
.A1(n_134),
.A2(n_95),
.B1(n_78),
.B2(n_74),
.Y(n_221)
);

INVxp67_ASAP7_75t_L g301 ( 
.A(n_221),
.Y(n_301)
);

MAJIxp5_ASAP7_75t_L g222 ( 
.A(n_125),
.B(n_98),
.C(n_7),
.Y(n_222)
);

MAJIxp5_ASAP7_75t_L g283 ( 
.A(n_222),
.B(n_241),
.C(n_253),
.Y(n_283)
);

AOI22xp33_ASAP7_75t_SL g223 ( 
.A1(n_146),
.A2(n_6),
.B1(n_7),
.B2(n_8),
.Y(n_223)
);

INVxp67_ASAP7_75t_L g305 ( 
.A(n_223),
.Y(n_305)
);

INVx2_ASAP7_75t_L g224 ( 
.A(n_136),
.Y(n_224)
);

INVx2_ASAP7_75t_L g308 ( 
.A(n_224),
.Y(n_308)
);

INVx2_ASAP7_75t_L g225 ( 
.A(n_136),
.Y(n_225)
);

INVx2_ASAP7_75t_L g316 ( 
.A(n_225),
.Y(n_316)
);

INVx2_ASAP7_75t_L g226 ( 
.A(n_170),
.Y(n_226)
);

HB1xp67_ASAP7_75t_L g278 ( 
.A(n_226),
.Y(n_278)
);

INVx6_ASAP7_75t_L g227 ( 
.A(n_143),
.Y(n_227)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_227),
.Y(n_287)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_131),
.Y(n_228)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_228),
.Y(n_289)
);

HB1xp67_ASAP7_75t_L g230 ( 
.A(n_180),
.Y(n_230)
);

CKINVDCx16_ASAP7_75t_R g295 ( 
.A(n_230),
.Y(n_295)
);

NOR2xp33_ASAP7_75t_L g232 ( 
.A(n_137),
.B(n_124),
.Y(n_232)
);

NOR2xp33_ASAP7_75t_L g275 ( 
.A(n_232),
.B(n_234),
.Y(n_275)
);

NOR2xp33_ASAP7_75t_L g234 ( 
.A(n_149),
.B(n_7),
.Y(n_234)
);

INVxp67_ASAP7_75t_L g235 ( 
.A(n_132),
.Y(n_235)
);

NOR2xp33_ASAP7_75t_L g299 ( 
.A(n_235),
.B(n_245),
.Y(n_299)
);

NAND2xp5_ASAP7_75t_L g236 ( 
.A(n_147),
.B(n_8),
.Y(n_236)
);

BUFx3_ASAP7_75t_L g237 ( 
.A(n_130),
.Y(n_237)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_237),
.Y(n_293)
);

INVx3_ASAP7_75t_L g238 ( 
.A(n_199),
.Y(n_238)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_238),
.Y(n_298)
);

AOI22xp5_ASAP7_75t_L g274 ( 
.A1(n_239),
.A2(n_193),
.B1(n_160),
.B2(n_177),
.Y(n_274)
);

BUFx3_ASAP7_75t_L g240 ( 
.A(n_138),
.Y(n_240)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_240),
.Y(n_314)
);

MAJIxp5_ASAP7_75t_L g241 ( 
.A(n_125),
.B(n_9),
.C(n_151),
.Y(n_241)
);

NAND2xp5_ASAP7_75t_L g242 ( 
.A(n_184),
.B(n_9),
.Y(n_242)
);

NAND2xp5_ASAP7_75t_SL g313 ( 
.A(n_242),
.B(n_249),
.Y(n_313)
);

INVx2_ASAP7_75t_L g243 ( 
.A(n_157),
.Y(n_243)
);

AND2x2_ASAP7_75t_L g309 ( 
.A(n_243),
.B(n_248),
.Y(n_309)
);

OAI22xp33_ASAP7_75t_SL g269 ( 
.A1(n_244),
.A2(n_141),
.B1(n_191),
.B2(n_165),
.Y(n_269)
);

CKINVDCx16_ASAP7_75t_R g245 ( 
.A(n_155),
.Y(n_245)
);

CKINVDCx20_ASAP7_75t_R g246 ( 
.A(n_127),
.Y(n_246)
);

NOR2xp33_ASAP7_75t_L g302 ( 
.A(n_246),
.B(n_251),
.Y(n_302)
);

AOI22xp5_ASAP7_75t_SL g247 ( 
.A1(n_196),
.A2(n_152),
.B1(n_127),
.B2(n_126),
.Y(n_247)
);

OAI21xp5_ASAP7_75t_L g272 ( 
.A1(n_247),
.A2(n_263),
.B(n_265),
.Y(n_272)
);

INVx3_ASAP7_75t_L g248 ( 
.A(n_144),
.Y(n_248)
);

NAND2xp5_ASAP7_75t_L g249 ( 
.A(n_189),
.B(n_186),
.Y(n_249)
);

AOI22xp33_ASAP7_75t_L g250 ( 
.A1(n_143),
.A2(n_182),
.B1(n_187),
.B2(n_133),
.Y(n_250)
);

INVxp67_ASAP7_75t_L g251 ( 
.A(n_126),
.Y(n_251)
);

INVx2_ASAP7_75t_L g252 ( 
.A(n_157),
.Y(n_252)
);

AND2x2_ASAP7_75t_L g312 ( 
.A(n_252),
.B(n_258),
.Y(n_312)
);

MAJIxp5_ASAP7_75t_L g253 ( 
.A(n_200),
.B(n_135),
.C(n_140),
.Y(n_253)
);

NOR2xp33_ASAP7_75t_L g254 ( 
.A(n_138),
.B(n_190),
.Y(n_254)
);

NOR2xp33_ASAP7_75t_L g317 ( 
.A(n_254),
.B(n_259),
.Y(n_317)
);

NAND2xp5_ASAP7_75t_L g255 ( 
.A(n_182),
.B(n_144),
.Y(n_255)
);

MAJIxp5_ASAP7_75t_L g304 ( 
.A(n_255),
.B(n_257),
.C(n_260),
.Y(n_304)
);

NAND2xp5_ASAP7_75t_L g257 ( 
.A(n_173),
.B(n_183),
.Y(n_257)
);

NAND2xp5_ASAP7_75t_SL g259 ( 
.A(n_190),
.B(n_173),
.Y(n_259)
);

NAND2xp5_ASAP7_75t_L g260 ( 
.A(n_175),
.B(n_185),
.Y(n_260)
);

CKINVDCx20_ASAP7_75t_R g261 ( 
.A(n_172),
.Y(n_261)
);

CKINVDCx20_ASAP7_75t_R g284 ( 
.A(n_261),
.Y(n_284)
);

AOI22xp33_ASAP7_75t_SL g262 ( 
.A1(n_123),
.A2(n_158),
.B1(n_167),
.B2(n_145),
.Y(n_262)
);

AOI22xp33_ASAP7_75t_SL g279 ( 
.A1(n_262),
.A2(n_174),
.B1(n_193),
.B2(n_251),
.Y(n_279)
);

AND2x2_ASAP7_75t_SL g263 ( 
.A(n_158),
.B(n_192),
.Y(n_263)
);

INVx4_ASAP7_75t_L g264 ( 
.A(n_192),
.Y(n_264)
);

CKINVDCx20_ASAP7_75t_R g285 ( 
.A(n_264),
.Y(n_285)
);

AND2x2_ASAP7_75t_L g265 ( 
.A(n_160),
.B(n_187),
.Y(n_265)
);

MAJx2_ASAP7_75t_L g266 ( 
.A(n_177),
.B(n_167),
.C(n_174),
.Y(n_266)
);

AOI21xp5_ASAP7_75t_L g276 ( 
.A1(n_266),
.A2(n_177),
.B(n_174),
.Y(n_276)
);

CKINVDCx20_ASAP7_75t_R g267 ( 
.A(n_172),
.Y(n_267)
);

CKINVDCx20_ASAP7_75t_R g286 ( 
.A(n_267),
.Y(n_286)
);

AOI22xp5_ASAP7_75t_SL g357 ( 
.A1(n_269),
.A2(n_303),
.B1(n_319),
.B2(n_273),
.Y(n_357)
);

AOI22xp33_ASAP7_75t_SL g336 ( 
.A1(n_273),
.A2(n_279),
.B1(n_315),
.B2(n_318),
.Y(n_336)
);

OAI22xp5_ASAP7_75t_L g351 ( 
.A1(n_274),
.A2(n_288),
.B1(n_305),
.B2(n_299),
.Y(n_351)
);

OAI21xp5_ASAP7_75t_SL g356 ( 
.A1(n_276),
.A2(n_312),
.B(n_281),
.Y(n_356)
);

AOI22xp5_ASAP7_75t_L g288 ( 
.A1(n_256),
.A2(n_233),
.B1(n_239),
.B2(n_257),
.Y(n_288)
);

AOI21xp5_ASAP7_75t_L g292 ( 
.A1(n_253),
.A2(n_258),
.B(n_201),
.Y(n_292)
);

AOI21xp5_ASAP7_75t_L g345 ( 
.A1(n_292),
.A2(n_276),
.B(n_283),
.Y(n_345)
);

AO22x1_ASAP7_75t_SL g296 ( 
.A1(n_244),
.A2(n_220),
.B1(n_266),
.B2(n_247),
.Y(n_296)
);

AO22x1_ASAP7_75t_SL g333 ( 
.A1(n_296),
.A2(n_263),
.B1(n_226),
.B2(n_214),
.Y(n_333)
);

OAI22xp33_ASAP7_75t_SL g303 ( 
.A1(n_206),
.A2(n_235),
.B1(n_215),
.B2(n_222),
.Y(n_303)
);

AOI22xp33_ASAP7_75t_SL g307 ( 
.A1(n_236),
.A2(n_238),
.B1(n_208),
.B2(n_229),
.Y(n_307)
);

INVxp67_ASAP7_75t_L g320 ( 
.A(n_307),
.Y(n_320)
);

CKINVDCx20_ASAP7_75t_R g310 ( 
.A(n_249),
.Y(n_310)
);

NOR2xp33_ASAP7_75t_L g327 ( 
.A(n_310),
.B(n_201),
.Y(n_327)
);

AOI22xp33_ASAP7_75t_SL g311 ( 
.A1(n_208),
.A2(n_264),
.B1(n_260),
.B2(n_255),
.Y(n_311)
);

INVxp67_ASAP7_75t_L g348 ( 
.A(n_311),
.Y(n_348)
);

AOI22xp33_ASAP7_75t_SL g315 ( 
.A1(n_248),
.A2(n_219),
.B1(n_204),
.B2(n_228),
.Y(n_315)
);

AOI22xp33_ASAP7_75t_SL g318 ( 
.A1(n_205),
.A2(n_218),
.B1(n_240),
.B2(n_237),
.Y(n_318)
);

AOI22xp33_ASAP7_75t_SL g319 ( 
.A1(n_224),
.A2(n_225),
.B1(n_263),
.B2(n_252),
.Y(n_319)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_289),
.Y(n_321)
);

INVx1_ASAP7_75t_L g387 ( 
.A(n_321),
.Y(n_387)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_289),
.Y(n_322)
);

INVx1_ASAP7_75t_L g390 ( 
.A(n_322),
.Y(n_390)
);

INVxp33_ASAP7_75t_L g323 ( 
.A(n_309),
.Y(n_323)
);

INVxp67_ASAP7_75t_SL g377 ( 
.A(n_323),
.Y(n_377)
);

MAJIxp5_ASAP7_75t_L g324 ( 
.A(n_300),
.B(n_201),
.C(n_258),
.Y(n_324)
);

MAJIxp5_ASAP7_75t_L g362 ( 
.A(n_324),
.B(n_344),
.C(n_346),
.Y(n_362)
);

OAI22xp5_ASAP7_75t_SL g325 ( 
.A1(n_288),
.A2(n_210),
.B1(n_242),
.B2(n_202),
.Y(n_325)
);

AOI22xp5_ASAP7_75t_L g378 ( 
.A1(n_325),
.A2(n_347),
.B1(n_350),
.B2(n_351),
.Y(n_378)
);

CKINVDCx20_ASAP7_75t_R g326 ( 
.A(n_278),
.Y(n_326)
);

NAND2xp5_ASAP7_75t_L g373 ( 
.A(n_326),
.B(n_328),
.Y(n_373)
);

NAND2xp5_ASAP7_75t_SL g383 ( 
.A(n_327),
.B(n_334),
.Y(n_383)
);

NAND2xp5_ASAP7_75t_L g328 ( 
.A(n_310),
.B(n_241),
.Y(n_328)
);

NAND2xp5_ASAP7_75t_L g329 ( 
.A(n_313),
.B(n_217),
.Y(n_329)
);

NAND2xp5_ASAP7_75t_L g379 ( 
.A(n_329),
.B(n_331),
.Y(n_379)
);

NOR2xp33_ASAP7_75t_L g330 ( 
.A(n_275),
.B(n_231),
.Y(n_330)
);

NOR2xp33_ASAP7_75t_SL g386 ( 
.A(n_330),
.B(n_337),
.Y(n_386)
);

CKINVDCx20_ASAP7_75t_R g331 ( 
.A(n_309),
.Y(n_331)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_280),
.Y(n_332)
);

INVx2_ASAP7_75t_L g363 ( 
.A(n_332),
.Y(n_363)
);

XNOR2x1_ASAP7_75t_L g391 ( 
.A(n_333),
.B(n_343),
.Y(n_391)
);

NAND2xp5_ASAP7_75t_L g334 ( 
.A(n_313),
.B(n_203),
.Y(n_334)
);

NAND2xp5_ASAP7_75t_L g335 ( 
.A(n_304),
.B(n_243),
.Y(n_335)
);

XNOR2xp5_ASAP7_75t_L g371 ( 
.A(n_335),
.B(n_342),
.Y(n_371)
);

NAND2xp5_ASAP7_75t_SL g337 ( 
.A(n_277),
.B(n_265),
.Y(n_337)
);

AND2x2_ASAP7_75t_L g338 ( 
.A(n_312),
.B(n_265),
.Y(n_338)
);

AND2x2_ASAP7_75t_L g370 ( 
.A(n_338),
.B(n_353),
.Y(n_370)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_280),
.Y(n_339)
);

INVx2_ASAP7_75t_L g388 ( 
.A(n_339),
.Y(n_388)
);

NOR2xp33_ASAP7_75t_SL g340 ( 
.A(n_277),
.B(n_227),
.Y(n_340)
);

CKINVDCx14_ASAP7_75t_R g374 ( 
.A(n_340),
.Y(n_374)
);

CKINVDCx20_ASAP7_75t_R g341 ( 
.A(n_309),
.Y(n_341)
);

CKINVDCx20_ASAP7_75t_R g361 ( 
.A(n_341),
.Y(n_361)
);

NAND2xp5_ASAP7_75t_L g342 ( 
.A(n_304),
.B(n_212),
.Y(n_342)
);

XNOR2xp5_ASAP7_75t_L g343 ( 
.A(n_300),
.B(n_292),
.Y(n_343)
);

XOR2xp5_ASAP7_75t_L g344 ( 
.A(n_300),
.B(n_283),
.Y(n_344)
);

OAI21xp5_ASAP7_75t_SL g359 ( 
.A1(n_345),
.A2(n_349),
.B(n_357),
.Y(n_359)
);

MAJIxp5_ASAP7_75t_L g346 ( 
.A(n_296),
.B(n_268),
.C(n_302),
.Y(n_346)
);

OAI22xp33_ASAP7_75t_SL g347 ( 
.A1(n_291),
.A2(n_274),
.B1(n_301),
.B2(n_296),
.Y(n_347)
);

AOI21xp33_ASAP7_75t_L g349 ( 
.A1(n_272),
.A2(n_296),
.B(n_268),
.Y(n_349)
);

OAI22xp5_ASAP7_75t_SL g350 ( 
.A1(n_291),
.A2(n_272),
.B1(n_301),
.B2(n_305),
.Y(n_350)
);

NAND2xp5_ASAP7_75t_SL g352 ( 
.A(n_317),
.B(n_271),
.Y(n_352)
);

XOR2xp5_ASAP7_75t_L g367 ( 
.A(n_352),
.B(n_287),
.Y(n_367)
);

INVx1_ASAP7_75t_L g353 ( 
.A(n_281),
.Y(n_353)
);

NOR2xp33_ASAP7_75t_SL g354 ( 
.A(n_284),
.B(n_286),
.Y(n_354)
);

CKINVDCx16_ASAP7_75t_R g372 ( 
.A(n_354),
.Y(n_372)
);

OAI21xp5_ASAP7_75t_L g355 ( 
.A1(n_284),
.A2(n_286),
.B(n_312),
.Y(n_355)
);

OAI21xp5_ASAP7_75t_L g360 ( 
.A1(n_355),
.A2(n_358),
.B(n_285),
.Y(n_360)
);

AOI21xp5_ASAP7_75t_L g364 ( 
.A1(n_356),
.A2(n_298),
.B(n_293),
.Y(n_364)
);

NOR2xp33_ASAP7_75t_L g358 ( 
.A(n_285),
.B(n_295),
.Y(n_358)
);

INVxp67_ASAP7_75t_L g394 ( 
.A(n_360),
.Y(n_394)
);

OAI21xp5_ASAP7_75t_SL g418 ( 
.A1(n_364),
.A2(n_376),
.B(n_381),
.Y(n_418)
);

OAI21xp5_ASAP7_75t_L g365 ( 
.A1(n_355),
.A2(n_298),
.B(n_314),
.Y(n_365)
);

AOI21xp5_ASAP7_75t_L g396 ( 
.A1(n_365),
.A2(n_368),
.B(n_369),
.Y(n_396)
);

OAI22xp5_ASAP7_75t_L g366 ( 
.A1(n_357),
.A2(n_287),
.B1(n_270),
.B2(n_316),
.Y(n_366)
);

AOI22xp5_ASAP7_75t_L g392 ( 
.A1(n_366),
.A2(n_321),
.B1(n_322),
.B2(n_341),
.Y(n_392)
);

XOR2xp5_ASAP7_75t_L g400 ( 
.A(n_367),
.B(n_343),
.Y(n_400)
);

OAI21xp5_ASAP7_75t_L g368 ( 
.A1(n_320),
.A2(n_293),
.B(n_314),
.Y(n_368)
);

OAI21xp5_ASAP7_75t_L g369 ( 
.A1(n_356),
.A2(n_290),
.B(n_306),
.Y(n_369)
);

CKINVDCx20_ASAP7_75t_R g375 ( 
.A(n_354),
.Y(n_375)
);

NOR2xp33_ASAP7_75t_L g401 ( 
.A(n_375),
.B(n_340),
.Y(n_401)
);

OAI21xp5_ASAP7_75t_L g376 ( 
.A1(n_348),
.A2(n_290),
.B(n_306),
.Y(n_376)
);

AOI22xp5_ASAP7_75t_L g380 ( 
.A1(n_351),
.A2(n_316),
.B1(n_308),
.B2(n_270),
.Y(n_380)
);

OAI22xp5_ASAP7_75t_SL g410 ( 
.A1(n_380),
.A2(n_384),
.B1(n_353),
.B2(n_339),
.Y(n_410)
);

AOI21xp5_ASAP7_75t_L g381 ( 
.A1(n_345),
.A2(n_290),
.B(n_306),
.Y(n_381)
);

XOR2xp5_ASAP7_75t_L g382 ( 
.A(n_344),
.B(n_295),
.Y(n_382)
);

MAJIxp5_ASAP7_75t_L g408 ( 
.A(n_382),
.B(n_337),
.C(n_327),
.Y(n_408)
);

AOI22xp5_ASAP7_75t_L g384 ( 
.A1(n_347),
.A2(n_308),
.B1(n_270),
.B2(n_294),
.Y(n_384)
);

AOI21xp5_ASAP7_75t_L g385 ( 
.A1(n_349),
.A2(n_297),
.B(n_282),
.Y(n_385)
);

AND2x2_ASAP7_75t_L g399 ( 
.A(n_385),
.B(n_389),
.Y(n_399)
);

AND2x2_ASAP7_75t_L g389 ( 
.A(n_338),
.B(n_282),
.Y(n_389)
);

OAI22xp5_ASAP7_75t_L g423 ( 
.A1(n_392),
.A2(n_402),
.B1(n_406),
.B2(n_415),
.Y(n_423)
);

NAND2xp5_ASAP7_75t_L g393 ( 
.A(n_375),
.B(n_334),
.Y(n_393)
);

INVx1_ASAP7_75t_L g422 ( 
.A(n_393),
.Y(n_422)
);

INVx1_ASAP7_75t_L g395 ( 
.A(n_363),
.Y(n_395)
);

INVx1_ASAP7_75t_L g425 ( 
.A(n_395),
.Y(n_425)
);

OAI22xp5_ASAP7_75t_L g397 ( 
.A1(n_378),
.A2(n_342),
.B1(n_335),
.B2(n_336),
.Y(n_397)
);

AOI22xp5_ASAP7_75t_L g426 ( 
.A1(n_397),
.A2(n_403),
.B1(n_373),
.B2(n_367),
.Y(n_426)
);

CKINVDCx14_ASAP7_75t_R g398 ( 
.A(n_379),
.Y(n_398)
);

NAND2xp5_ASAP7_75t_L g436 ( 
.A(n_398),
.B(n_401),
.Y(n_436)
);

XNOR2xp5_ASAP7_75t_SL g430 ( 
.A(n_400),
.B(n_407),
.Y(n_430)
);

AOI22xp5_ASAP7_75t_SL g402 ( 
.A1(n_374),
.A2(n_350),
.B1(n_346),
.B2(n_324),
.Y(n_402)
);

OAI22xp5_ASAP7_75t_L g403 ( 
.A1(n_378),
.A2(n_373),
.B1(n_372),
.B2(n_380),
.Y(n_403)
);

INVx1_ASAP7_75t_L g404 ( 
.A(n_363),
.Y(n_404)
);

INVx1_ASAP7_75t_L g439 ( 
.A(n_404),
.Y(n_439)
);

CKINVDCx20_ASAP7_75t_R g405 ( 
.A(n_372),
.Y(n_405)
);

NOR2xp33_ASAP7_75t_L g424 ( 
.A(n_405),
.B(n_412),
.Y(n_424)
);

AOI22xp5_ASAP7_75t_L g406 ( 
.A1(n_366),
.A2(n_325),
.B1(n_333),
.B2(n_328),
.Y(n_406)
);

XOR2xp5_ASAP7_75t_L g407 ( 
.A(n_362),
.B(n_329),
.Y(n_407)
);

XNOR2xp5_ASAP7_75t_L g420 ( 
.A(n_408),
.B(n_362),
.Y(n_420)
);

NOR2xp33_ASAP7_75t_L g409 ( 
.A(n_386),
.B(n_352),
.Y(n_409)
);

INVx1_ASAP7_75t_L g441 ( 
.A(n_409),
.Y(n_441)
);

INVx1_ASAP7_75t_L g427 ( 
.A(n_410),
.Y(n_427)
);

OR2x2_ASAP7_75t_L g411 ( 
.A(n_379),
.B(n_333),
.Y(n_411)
);

INVx1_ASAP7_75t_L g431 ( 
.A(n_411),
.Y(n_431)
);

CKINVDCx20_ASAP7_75t_R g412 ( 
.A(n_370),
.Y(n_412)
);

NOR2xp33_ASAP7_75t_SL g413 ( 
.A(n_386),
.B(n_330),
.Y(n_413)
);

NAND2xp5_ASAP7_75t_SL g440 ( 
.A(n_413),
.B(n_409),
.Y(n_440)
);

INVx1_ASAP7_75t_L g414 ( 
.A(n_388),
.Y(n_414)
);

INVxp67_ASAP7_75t_L g429 ( 
.A(n_414),
.Y(n_429)
);

AOI22xp5_ASAP7_75t_SL g415 ( 
.A1(n_361),
.A2(n_338),
.B1(n_336),
.B2(n_331),
.Y(n_415)
);

AOI22xp33_ASAP7_75t_L g416 ( 
.A1(n_361),
.A2(n_338),
.B1(n_333),
.B2(n_358),
.Y(n_416)
);

OAI22xp5_ASAP7_75t_SL g421 ( 
.A1(n_416),
.A2(n_360),
.B1(n_385),
.B2(n_364),
.Y(n_421)
);

CKINVDCx20_ASAP7_75t_R g417 ( 
.A(n_370),
.Y(n_417)
);

NOR2xp33_ASAP7_75t_L g432 ( 
.A(n_417),
.B(n_419),
.Y(n_432)
);

INVx1_ASAP7_75t_L g419 ( 
.A(n_388),
.Y(n_419)
);

MAJIxp5_ASAP7_75t_L g446 ( 
.A(n_420),
.B(n_400),
.C(n_371),
.Y(n_446)
);

AOI22xp5_ASAP7_75t_L g451 ( 
.A1(n_421),
.A2(n_433),
.B1(n_434),
.B2(n_397),
.Y(n_451)
);

INVx1_ASAP7_75t_L g454 ( 
.A(n_426),
.Y(n_454)
);

XNOR2x1_ASAP7_75t_L g428 ( 
.A(n_402),
.B(n_382),
.Y(n_428)
);

XOR2xp5_ASAP7_75t_L g447 ( 
.A(n_428),
.B(n_437),
.Y(n_447)
);

OAI22xp5_ASAP7_75t_SL g433 ( 
.A1(n_406),
.A2(n_384),
.B1(n_359),
.B2(n_383),
.Y(n_433)
);

OAI22xp5_ASAP7_75t_SL g434 ( 
.A1(n_411),
.A2(n_359),
.B1(n_383),
.B2(n_391),
.Y(n_434)
);

NOR3xp33_ASAP7_75t_SL g435 ( 
.A(n_393),
.B(n_405),
.C(n_413),
.Y(n_435)
);

NOR2xp33_ASAP7_75t_L g450 ( 
.A(n_435),
.B(n_442),
.Y(n_450)
);

XNOR2xp5_ASAP7_75t_L g437 ( 
.A(n_407),
.B(n_408),
.Y(n_437)
);

OAI21xp5_ASAP7_75t_L g438 ( 
.A1(n_396),
.A2(n_365),
.B(n_381),
.Y(n_438)
);

OAI21xp5_ASAP7_75t_L g455 ( 
.A1(n_438),
.A2(n_443),
.B(n_444),
.Y(n_455)
);

NOR2xp33_ASAP7_75t_SL g445 ( 
.A(n_440),
.B(n_417),
.Y(n_445)
);

CKINVDCx20_ASAP7_75t_R g442 ( 
.A(n_401),
.Y(n_442)
);

AOI22xp5_ASAP7_75t_SL g443 ( 
.A1(n_394),
.A2(n_370),
.B1(n_389),
.B2(n_391),
.Y(n_443)
);

AOI21xp5_ASAP7_75t_L g444 ( 
.A1(n_418),
.A2(n_368),
.B(n_369),
.Y(n_444)
);

INVx1_ASAP7_75t_L g475 ( 
.A(n_445),
.Y(n_475)
);

NAND2xp5_ASAP7_75t_SL g467 ( 
.A(n_446),
.B(n_452),
.Y(n_467)
);

NOR2xp33_ASAP7_75t_L g448 ( 
.A(n_436),
.B(n_398),
.Y(n_448)
);

INVx1_ASAP7_75t_L g478 ( 
.A(n_448),
.Y(n_478)
);

NAND2xp5_ASAP7_75t_L g449 ( 
.A(n_436),
.B(n_403),
.Y(n_449)
);

INVx1_ASAP7_75t_L g481 ( 
.A(n_449),
.Y(n_481)
);

OAI22xp5_ASAP7_75t_SL g466 ( 
.A1(n_451),
.A2(n_456),
.B1(n_458),
.B2(n_443),
.Y(n_466)
);

NOR2xp33_ASAP7_75t_L g452 ( 
.A(n_441),
.B(n_426),
.Y(n_452)
);

CKINVDCx20_ASAP7_75t_R g453 ( 
.A(n_424),
.Y(n_453)
);

NAND2xp5_ASAP7_75t_L g476 ( 
.A(n_453),
.B(n_460),
.Y(n_476)
);

AOI22xp5_ASAP7_75t_L g456 ( 
.A1(n_433),
.A2(n_399),
.B1(n_410),
.B2(n_412),
.Y(n_456)
);

NAND2xp5_ASAP7_75t_L g457 ( 
.A(n_429),
.B(n_392),
.Y(n_457)
);

INVx1_ASAP7_75t_L g482 ( 
.A(n_457),
.Y(n_482)
);

AOI22xp5_ASAP7_75t_SL g458 ( 
.A1(n_421),
.A2(n_423),
.B1(n_399),
.B2(n_427),
.Y(n_458)
);

XOR2xp5_ASAP7_75t_L g459 ( 
.A(n_430),
.B(n_371),
.Y(n_459)
);

XOR2xp5_ASAP7_75t_L g471 ( 
.A(n_459),
.B(n_462),
.Y(n_471)
);

NAND2xp5_ASAP7_75t_L g460 ( 
.A(n_429),
.B(n_395),
.Y(n_460)
);

INVx1_ASAP7_75t_L g461 ( 
.A(n_432),
.Y(n_461)
);

NAND2xp5_ASAP7_75t_L g480 ( 
.A(n_461),
.B(n_463),
.Y(n_480)
);

XOR2xp5_ASAP7_75t_L g462 ( 
.A(n_430),
.B(n_415),
.Y(n_462)
);

INVx1_ASAP7_75t_L g463 ( 
.A(n_431),
.Y(n_463)
);

NOR2xp33_ASAP7_75t_L g464 ( 
.A(n_437),
.B(n_326),
.Y(n_464)
);

NOR2xp33_ASAP7_75t_L g469 ( 
.A(n_464),
.B(n_420),
.Y(n_469)
);

NAND2xp5_ASAP7_75t_L g465 ( 
.A(n_431),
.B(n_419),
.Y(n_465)
);

NOR2xp67_ASAP7_75t_R g474 ( 
.A(n_465),
.B(n_411),
.Y(n_474)
);

AOI22xp33_ASAP7_75t_SL g486 ( 
.A1(n_466),
.A2(n_454),
.B1(n_449),
.B2(n_457),
.Y(n_486)
);

AOI22xp5_ASAP7_75t_L g468 ( 
.A1(n_454),
.A2(n_427),
.B1(n_434),
.B2(n_422),
.Y(n_468)
);

OAI22xp33_ASAP7_75t_SL g495 ( 
.A1(n_468),
.A2(n_474),
.B1(n_456),
.B2(n_463),
.Y(n_495)
);

HB1xp67_ASAP7_75t_L g488 ( 
.A(n_469),
.Y(n_488)
);

A2O1A1O1Ixp25_ASAP7_75t_L g470 ( 
.A1(n_448),
.A2(n_422),
.B(n_438),
.C(n_435),
.D(n_418),
.Y(n_470)
);

NAND2xp5_ASAP7_75t_L g490 ( 
.A(n_470),
.B(n_455),
.Y(n_490)
);

NOR2xp33_ASAP7_75t_L g472 ( 
.A(n_453),
.B(n_416),
.Y(n_472)
);

INVx1_ASAP7_75t_L g494 ( 
.A(n_472),
.Y(n_494)
);

NOR2xp33_ASAP7_75t_L g473 ( 
.A(n_445),
.B(n_461),
.Y(n_473)
);

CKINVDCx16_ASAP7_75t_R g493 ( 
.A(n_473),
.Y(n_493)
);

XNOR2xp5_ASAP7_75t_SL g477 ( 
.A(n_462),
.B(n_428),
.Y(n_477)
);

XNOR2xp5_ASAP7_75t_L g484 ( 
.A(n_477),
.B(n_479),
.Y(n_484)
);

XOR2xp5_ASAP7_75t_L g479 ( 
.A(n_459),
.B(n_444),
.Y(n_479)
);

NOR2xp33_ASAP7_75t_L g483 ( 
.A(n_467),
.B(n_450),
.Y(n_483)
);

NOR2xp33_ASAP7_75t_SL g505 ( 
.A(n_483),
.B(n_387),
.Y(n_505)
);

AOI21xp5_ASAP7_75t_L g485 ( 
.A1(n_475),
.A2(n_455),
.B(n_458),
.Y(n_485)
);

OAI21xp5_ASAP7_75t_L g501 ( 
.A1(n_485),
.A2(n_486),
.B(n_470),
.Y(n_501)
);

INVx1_ASAP7_75t_L g487 ( 
.A(n_476),
.Y(n_487)
);

NAND2xp5_ASAP7_75t_L g506 ( 
.A(n_487),
.B(n_492),
.Y(n_506)
);

MAJIxp5_ASAP7_75t_L g489 ( 
.A(n_471),
.B(n_446),
.C(n_447),
.Y(n_489)
);

NAND2xp5_ASAP7_75t_L g500 ( 
.A(n_489),
.B(n_491),
.Y(n_500)
);

AOI21xp5_ASAP7_75t_L g502 ( 
.A1(n_490),
.A2(n_399),
.B(n_396),
.Y(n_502)
);

MAJIxp5_ASAP7_75t_L g491 ( 
.A(n_471),
.B(n_447),
.C(n_451),
.Y(n_491)
);

NAND2xp5_ASAP7_75t_L g492 ( 
.A(n_478),
.B(n_476),
.Y(n_492)
);

AOI22xp5_ASAP7_75t_L g496 ( 
.A1(n_495),
.A2(n_466),
.B1(n_482),
.B2(n_481),
.Y(n_496)
);

INVx1_ASAP7_75t_L g515 ( 
.A(n_496),
.Y(n_515)
);

NAND2xp5_ASAP7_75t_SL g497 ( 
.A(n_493),
.B(n_480),
.Y(n_497)
);

NAND2xp5_ASAP7_75t_L g508 ( 
.A(n_497),
.B(n_498),
.Y(n_508)
);

MAJIxp5_ASAP7_75t_L g498 ( 
.A(n_491),
.B(n_479),
.C(n_468),
.Y(n_498)
);

NOR2xp33_ASAP7_75t_L g499 ( 
.A(n_488),
.B(n_480),
.Y(n_499)
);

NAND2xp5_ASAP7_75t_SL g514 ( 
.A(n_499),
.B(n_505),
.Y(n_514)
);

AND2x2_ASAP7_75t_L g510 ( 
.A(n_501),
.B(n_502),
.Y(n_510)
);

AOI22xp5_ASAP7_75t_L g503 ( 
.A1(n_494),
.A2(n_439),
.B1(n_425),
.B2(n_465),
.Y(n_503)
);

OAI22xp5_ASAP7_75t_SL g513 ( 
.A1(n_503),
.A2(n_504),
.B1(n_377),
.B2(n_390),
.Y(n_513)
);

AOI22xp33_ASAP7_75t_SL g504 ( 
.A1(n_487),
.A2(n_474),
.B1(n_460),
.B2(n_414),
.Y(n_504)
);

MAJIxp5_ASAP7_75t_L g507 ( 
.A(n_498),
.B(n_489),
.C(n_485),
.Y(n_507)
);

NAND2xp5_ASAP7_75t_L g517 ( 
.A(n_507),
.B(n_509),
.Y(n_517)
);

AOI22xp5_ASAP7_75t_SL g509 ( 
.A1(n_506),
.A2(n_490),
.B1(n_492),
.B2(n_399),
.Y(n_509)
);

AOI22xp5_ASAP7_75t_SL g511 ( 
.A1(n_501),
.A2(n_477),
.B1(n_484),
.B2(n_404),
.Y(n_511)
);

XNOR2xp5_ASAP7_75t_L g516 ( 
.A(n_511),
.B(n_504),
.Y(n_516)
);

XNOR2xp5_ASAP7_75t_L g512 ( 
.A(n_500),
.B(n_484),
.Y(n_512)
);

NOR2xp33_ASAP7_75t_SL g519 ( 
.A(n_512),
.B(n_496),
.Y(n_519)
);

INVx1_ASAP7_75t_L g518 ( 
.A(n_513),
.Y(n_518)
);

OR2x2_ASAP7_75t_L g523 ( 
.A(n_516),
.B(n_519),
.Y(n_523)
);

OAI21xp5_ASAP7_75t_L g520 ( 
.A1(n_508),
.A2(n_389),
.B(n_387),
.Y(n_520)
);

AOI21xp5_ASAP7_75t_L g524 ( 
.A1(n_520),
.A2(n_510),
.B(n_511),
.Y(n_524)
);

INVx1_ASAP7_75t_L g521 ( 
.A(n_514),
.Y(n_521)
);

NAND2xp5_ASAP7_75t_L g522 ( 
.A(n_521),
.B(n_507),
.Y(n_522)
);

NOR2xp33_ASAP7_75t_L g527 ( 
.A(n_522),
.B(n_524),
.Y(n_527)
);

NAND2xp5_ASAP7_75t_L g525 ( 
.A(n_518),
.B(n_515),
.Y(n_525)
);

AOI321xp33_ASAP7_75t_L g526 ( 
.A1(n_525),
.A2(n_517),
.A3(n_390),
.B1(n_516),
.B2(n_510),
.C(n_332),
.Y(n_526)
);

MAJIxp5_ASAP7_75t_L g528 ( 
.A(n_526),
.B(n_523),
.C(n_376),
.Y(n_528)
);

OAI21x1_ASAP7_75t_L g529 ( 
.A1(n_528),
.A2(n_527),
.B(n_297),
.Y(n_529)
);

NAND2xp5_ASAP7_75t_L g530 ( 
.A(n_529),
.B(n_294),
.Y(n_530)
);

BUFx24_ASAP7_75t_SL g531 ( 
.A(n_530),
.Y(n_531)
);


endmodule