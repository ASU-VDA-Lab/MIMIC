module real_jpeg_832_n_6 (n_5, n_4, n_0, n_1, n_2, n_3, n_6);

input n_5;
input n_4;
input n_0;
input n_1;
input n_2;
input n_3;

output n_6;

wire n_17;
wire n_43;
wire n_8;
wire n_37;
wire n_21;
wire n_35;
wire n_33;
wire n_38;
wire n_29;
wire n_49;
wire n_10;
wire n_31;
wire n_9;
wire n_12;
wire n_24;
wire n_34;
wire n_44;
wire n_28;
wire n_46;
wire n_23;
wire n_47;
wire n_14;
wire n_11;
wire n_45;
wire n_25;
wire n_42;
wire n_7;
wire n_22;
wire n_18;
wire n_40;
wire n_36;
wire n_39;
wire n_41;
wire n_27;
wire n_26;
wire n_20;
wire n_19;
wire n_48;
wire n_32;
wire n_30;
wire n_16;
wire n_15;
wire n_13;

NAND2xp5_ASAP7_75t_SL g8 ( 
.A(n_0),
.B(n_5),
.Y(n_8)
);

INVx1_ASAP7_75t_SL g12 ( 
.A(n_0),
.Y(n_12)
);

NAND2xp5_ASAP7_75t_L g36 ( 
.A(n_0),
.B(n_30),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g43 ( 
.A(n_0),
.B(n_44),
.Y(n_43)
);

NAND2xp5_ASAP7_75t_L g48 ( 
.A(n_0),
.B(n_49),
.Y(n_48)
);

OR2x4_ASAP7_75t_L g13 ( 
.A(n_1),
.B(n_14),
.Y(n_13)
);

AND2x2_ASAP7_75t_SL g30 ( 
.A(n_1),
.B(n_31),
.Y(n_30)
);

INVx1_ASAP7_75t_SL g41 ( 
.A(n_1),
.Y(n_41)
);

OA22x2_ASAP7_75t_L g16 ( 
.A1(n_2),
.A2(n_17),
.B1(n_18),
.B2(n_19),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_2),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_3),
.Y(n_22)
);

INVx1_ASAP7_75t_L g14 ( 
.A(n_4),
.Y(n_14)
);

OR2x2_ASAP7_75t_L g44 ( 
.A(n_4),
.B(n_41),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g21 ( 
.A(n_5),
.B(n_22),
.Y(n_21)
);

NAND2x1_ASAP7_75t_SL g23 ( 
.A(n_5),
.B(n_22),
.Y(n_23)
);

NAND2xp5_ASAP7_75t_L g42 ( 
.A(n_5),
.B(n_43),
.Y(n_42)
);

INVx1_ASAP7_75t_L g6 ( 
.A(n_7),
.Y(n_6)
);

AOI211xp5_ASAP7_75t_L g7 ( 
.A1(n_8),
.A2(n_9),
.B(n_25),
.C(n_47),
.Y(n_7)
);

NAND2xp5_ASAP7_75t_L g9 ( 
.A(n_10),
.B(n_15),
.Y(n_9)
);

CKINVDCx16_ASAP7_75t_R g10 ( 
.A(n_11),
.Y(n_10)
);

NOR2xp33_ASAP7_75t_L g11 ( 
.A(n_12),
.B(n_13),
.Y(n_11)
);

NAND2xp5_ASAP7_75t_L g29 ( 
.A(n_12),
.B(n_30),
.Y(n_29)
);

NAND2xp5_ASAP7_75t_L g39 ( 
.A(n_12),
.B(n_40),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_SL g46 ( 
.A(n_12),
.B(n_27),
.Y(n_46)
);

INVx1_ASAP7_75t_SL g24 ( 
.A(n_13),
.Y(n_24)
);

CKINVDCx16_ASAP7_75t_R g31 ( 
.A(n_14),
.Y(n_31)
);

AND2x2_ASAP7_75t_SL g40 ( 
.A(n_14),
.B(n_41),
.Y(n_40)
);

NAND2xp5_ASAP7_75t_SL g15 ( 
.A(n_16),
.B(n_24),
.Y(n_15)
);

NOR2xp33_ASAP7_75t_L g47 ( 
.A(n_16),
.B(n_48),
.Y(n_47)
);

OA21x2_ASAP7_75t_L g27 ( 
.A1(n_17),
.A2(n_21),
.B(n_23),
.Y(n_27)
);

OA21x2_ASAP7_75t_L g33 ( 
.A1(n_17),
.A2(n_20),
.B(n_34),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_19),
.Y(n_18)
);

AND2x2_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_23),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_21),
.Y(n_20)
);

CKINVDCx16_ASAP7_75t_R g34 ( 
.A(n_23),
.Y(n_34)
);

NAND4xp25_ASAP7_75t_L g25 ( 
.A(n_26),
.B(n_37),
.C(n_42),
.D(n_45),
.Y(n_25)
);

AOI22xp5_ASAP7_75t_L g26 ( 
.A1(n_27),
.A2(n_28),
.B1(n_32),
.B2(n_35),
.Y(n_26)
);

CKINVDCx16_ASAP7_75t_R g28 ( 
.A(n_29),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_33),
.Y(n_32)
);

NAND2xp5_ASAP7_75t_L g37 ( 
.A(n_33),
.B(n_38),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_36),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_39),
.Y(n_38)
);

NAND2xp5_ASAP7_75t_L g45 ( 
.A(n_40),
.B(n_46),
.Y(n_45)
);

INVx1_ASAP7_75t_SL g49 ( 
.A(n_44),
.Y(n_49)
);


endmodule