module fake_jpeg_24372_n_139 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_139);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_139;

wire n_117;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_73;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_29;
wire n_103;
wire n_50;
wire n_15;
wire n_124;
wire n_21;
wire n_57;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_30;
wire n_106;
wire n_111;
wire n_24;
wire n_44;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_78;
wire n_18;
wire n_20;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_97;
wire n_135;
wire n_36;
wire n_62;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_96;

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_2),
.Y(n_15)
);

BUFx12f_ASAP7_75t_L g16 ( 
.A(n_9),
.Y(n_16)
);

INVx5_ASAP7_75t_L g17 ( 
.A(n_3),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_5),
.Y(n_18)
);

BUFx12_ASAP7_75t_L g19 ( 
.A(n_14),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_0),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_3),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_9),
.Y(n_22)
);

INVx11_ASAP7_75t_L g23 ( 
.A(n_13),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_3),
.Y(n_24)
);

INVx2_ASAP7_75t_L g25 ( 
.A(n_14),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_10),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_12),
.Y(n_27)
);

INVx2_ASAP7_75t_L g28 ( 
.A(n_10),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_8),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_0),
.Y(n_30)
);

CKINVDCx9p33_ASAP7_75t_R g31 ( 
.A(n_23),
.Y(n_31)
);

INVx1_ASAP7_75t_SL g43 ( 
.A(n_31),
.Y(n_43)
);

INVx6_ASAP7_75t_SL g32 ( 
.A(n_16),
.Y(n_32)
);

NOR2xp33_ASAP7_75t_L g47 ( 
.A(n_32),
.B(n_36),
.Y(n_47)
);

OR2x2_ASAP7_75t_L g33 ( 
.A(n_15),
.B(n_0),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_33),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_L g34 ( 
.A(n_18),
.B(n_1),
.Y(n_34)
);

NAND2xp5_ASAP7_75t_L g54 ( 
.A(n_34),
.B(n_37),
.Y(n_54)
);

BUFx12f_ASAP7_75t_L g35 ( 
.A(n_16),
.Y(n_35)
);

CKINVDCx16_ASAP7_75t_R g49 ( 
.A(n_35),
.Y(n_49)
);

INVx3_ASAP7_75t_L g36 ( 
.A(n_23),
.Y(n_36)
);

NAND2xp5_ASAP7_75t_L g37 ( 
.A(n_18),
.B(n_24),
.Y(n_37)
);

INVx6_ASAP7_75t_SL g38 ( 
.A(n_16),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_38),
.B(n_19),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_SL g39 ( 
.A(n_20),
.B(n_1),
.Y(n_39)
);

NAND2xp5_ASAP7_75t_L g57 ( 
.A(n_39),
.B(n_29),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g40 ( 
.A(n_19),
.B(n_1),
.Y(n_40)
);

A2O1A1Ixp33_ASAP7_75t_L g46 ( 
.A1(n_40),
.A2(n_42),
.B(n_27),
.C(n_21),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_16),
.Y(n_41)
);

INVx4_ASAP7_75t_L g48 ( 
.A(n_41),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g42 ( 
.A(n_19),
.B(n_2),
.Y(n_42)
);

CKINVDCx14_ASAP7_75t_R g44 ( 
.A(n_40),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_44),
.B(n_46),
.Y(n_66)
);

OAI22xp5_ASAP7_75t_L g45 ( 
.A1(n_36),
.A2(n_28),
.B1(n_25),
.B2(n_17),
.Y(n_45)
);

OAI22xp5_ASAP7_75t_SL g67 ( 
.A1(n_45),
.A2(n_59),
.B1(n_26),
.B2(n_27),
.Y(n_67)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_37),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_L g61 ( 
.A(n_50),
.B(n_51),
.Y(n_61)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_34),
.Y(n_51)
);

AOI21xp33_ASAP7_75t_L g53 ( 
.A1(n_42),
.A2(n_22),
.B(n_30),
.Y(n_53)
);

AND2x2_ASAP7_75t_L g62 ( 
.A(n_53),
.B(n_57),
.Y(n_62)
);

BUFx12f_ASAP7_75t_L g55 ( 
.A(n_35),
.Y(n_55)
);

INVxp67_ASAP7_75t_L g63 ( 
.A(n_55),
.Y(n_63)
);

INVx4_ASAP7_75t_L g56 ( 
.A(n_35),
.Y(n_56)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_56),
.Y(n_70)
);

BUFx12f_ASAP7_75t_L g58 ( 
.A(n_35),
.Y(n_58)
);

INVxp67_ASAP7_75t_L g64 ( 
.A(n_58),
.Y(n_64)
);

OAI22xp5_ASAP7_75t_SL g59 ( 
.A1(n_35),
.A2(n_15),
.B1(n_30),
.B2(n_24),
.Y(n_59)
);

INVxp67_ASAP7_75t_L g71 ( 
.A(n_60),
.Y(n_71)
);

CKINVDCx20_ASAP7_75t_R g65 ( 
.A(n_59),
.Y(n_65)
);

CKINVDCx20_ASAP7_75t_R g92 ( 
.A(n_65),
.Y(n_92)
);

AND2x2_ASAP7_75t_L g83 ( 
.A(n_67),
.B(n_46),
.Y(n_83)
);

XNOR2xp5_ASAP7_75t_L g68 ( 
.A(n_54),
.B(n_38),
.Y(n_68)
);

MAJIxp5_ASAP7_75t_L g86 ( 
.A(n_68),
.B(n_73),
.C(n_58),
.Y(n_86)
);

CKINVDCx20_ASAP7_75t_R g69 ( 
.A(n_55),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_69),
.B(n_74),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_L g72 ( 
.A(n_54),
.B(n_33),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_L g81 ( 
.A(n_72),
.B(n_78),
.Y(n_81)
);

XNOR2xp5_ASAP7_75t_L g73 ( 
.A(n_57),
.B(n_38),
.Y(n_73)
);

INVxp67_ASAP7_75t_L g74 ( 
.A(n_47),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_56),
.B(n_32),
.Y(n_75)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_75),
.Y(n_82)
);

A2O1A1Ixp33_ASAP7_75t_SL g76 ( 
.A1(n_45),
.A2(n_41),
.B(n_4),
.C(n_6),
.Y(n_76)
);

OA22x2_ASAP7_75t_L g88 ( 
.A1(n_76),
.A2(n_58),
.B1(n_55),
.B2(n_43),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_49),
.B(n_2),
.Y(n_77)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_77),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g78 ( 
.A(n_52),
.B(n_41),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_L g79 ( 
.A(n_52),
.B(n_41),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_L g87 ( 
.A(n_79),
.B(n_80),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_L g80 ( 
.A(n_49),
.B(n_6),
.Y(n_80)
);

HB1xp67_ASAP7_75t_L g85 ( 
.A(n_70),
.Y(n_85)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_85),
.Y(n_101)
);

XNOR2xp5_ASAP7_75t_L g102 ( 
.A(n_86),
.B(n_73),
.Y(n_102)
);

MAJIxp5_ASAP7_75t_L g89 ( 
.A(n_68),
.B(n_58),
.C(n_55),
.Y(n_89)
);

MAJIxp5_ASAP7_75t_L g100 ( 
.A(n_89),
.B(n_86),
.C(n_93),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_L g91 ( 
.A(n_72),
.B(n_79),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_91),
.B(n_97),
.Y(n_99)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_78),
.Y(n_93)
);

CKINVDCx20_ASAP7_75t_R g94 ( 
.A(n_80),
.Y(n_94)
);

CKINVDCx20_ASAP7_75t_R g98 ( 
.A(n_94),
.Y(n_98)
);

INVx2_ASAP7_75t_L g95 ( 
.A(n_63),
.Y(n_95)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_95),
.Y(n_107)
);

BUFx3_ASAP7_75t_L g96 ( 
.A(n_63),
.Y(n_96)
);

CKINVDCx20_ASAP7_75t_R g109 ( 
.A(n_96),
.Y(n_109)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_61),
.Y(n_97)
);

MAJIxp5_ASAP7_75t_L g112 ( 
.A(n_100),
.B(n_87),
.C(n_97),
.Y(n_112)
);

XNOR2xp5_ASAP7_75t_L g113 ( 
.A(n_102),
.B(n_87),
.Y(n_113)
);

AOI22xp5_ASAP7_75t_L g103 ( 
.A1(n_89),
.A2(n_67),
.B1(n_66),
.B2(n_76),
.Y(n_103)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_81),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_SL g119 ( 
.A(n_104),
.B(n_105),
.Y(n_119)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_81),
.Y(n_105)
);

AO22x1_ASAP7_75t_L g106 ( 
.A1(n_88),
.A2(n_76),
.B1(n_62),
.B2(n_48),
.Y(n_106)
);

OAI21xp5_ASAP7_75t_L g118 ( 
.A1(n_106),
.A2(n_110),
.B(n_103),
.Y(n_118)
);

OAI22xp5_ASAP7_75t_SL g108 ( 
.A1(n_92),
.A2(n_76),
.B1(n_62),
.B2(n_71),
.Y(n_108)
);

AOI21xp5_ASAP7_75t_L g110 ( 
.A1(n_91),
.A2(n_64),
.B(n_74),
.Y(n_110)
);

XNOR2xp5_ASAP7_75t_SL g111 ( 
.A(n_102),
.B(n_83),
.Y(n_111)
);

MAJIxp5_ASAP7_75t_L g125 ( 
.A(n_111),
.B(n_112),
.C(n_113),
.Y(n_125)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_99),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g123 ( 
.A(n_114),
.B(n_116),
.Y(n_123)
);

MAJIxp5_ASAP7_75t_L g115 ( 
.A(n_100),
.B(n_90),
.C(n_82),
.Y(n_115)
);

MAJIxp5_ASAP7_75t_L g127 ( 
.A(n_115),
.B(n_121),
.C(n_107),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_SL g116 ( 
.A(n_98),
.B(n_82),
.Y(n_116)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_99),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_L g126 ( 
.A(n_117),
.B(n_120),
.Y(n_126)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_110),
.Y(n_120)
);

MAJIxp5_ASAP7_75t_L g121 ( 
.A(n_104),
.B(n_83),
.C(n_96),
.Y(n_121)
);

INVxp33_ASAP7_75t_L g122 ( 
.A(n_119),
.Y(n_122)
);

INVxp67_ASAP7_75t_L g128 ( 
.A(n_122),
.Y(n_128)
);

OAI21xp33_ASAP7_75t_L g124 ( 
.A1(n_118),
.A2(n_105),
.B(n_108),
.Y(n_124)
);

INVx5_ASAP7_75t_L g129 ( 
.A(n_122),
.Y(n_129)
);

AND2x2_ASAP7_75t_L g130 ( 
.A(n_123),
.B(n_124),
.Y(n_130)
);

AOI21xp5_ASAP7_75t_L g133 ( 
.A1(n_130),
.A2(n_101),
.B(n_64),
.Y(n_133)
);

AOI322xp5_ASAP7_75t_L g131 ( 
.A1(n_130),
.A2(n_126),
.A3(n_127),
.B1(n_125),
.B2(n_112),
.C1(n_109),
.C2(n_84),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_SL g136 ( 
.A(n_131),
.B(n_132),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_SL g132 ( 
.A(n_129),
.B(n_101),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_L g135 ( 
.A(n_133),
.B(n_134),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_SL g134 ( 
.A(n_128),
.B(n_11),
.Y(n_134)
);

AOI21xp5_ASAP7_75t_SL g137 ( 
.A1(n_135),
.A2(n_6),
.B(n_7),
.Y(n_137)
);

OAI33xp33_ASAP7_75t_L g138 ( 
.A1(n_137),
.A2(n_7),
.A3(n_43),
.B1(n_136),
.B2(n_134),
.B3(n_106),
.Y(n_138)
);

XOR2xp5_ASAP7_75t_L g139 ( 
.A(n_138),
.B(n_7),
.Y(n_139)
);


endmodule