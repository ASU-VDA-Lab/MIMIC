module fake_netlist_5_434_n_1938 (n_137, n_168, n_164, n_191, n_91, n_82, n_122, n_194, n_142, n_176, n_10, n_140, n_24, n_124, n_86, n_136, n_146, n_182, n_143, n_83, n_132, n_61, n_90, n_127, n_75, n_101, n_180, n_184, n_65, n_78, n_74, n_144, n_114, n_57, n_96, n_37, n_189, n_165, n_111, n_108, n_129, n_31, n_13, n_66, n_98, n_177, n_60, n_155, n_152, n_197, n_16, n_43, n_107, n_0, n_58, n_9, n_69, n_18, n_116, n_195, n_42, n_22, n_1, n_45, n_117, n_46, n_21, n_94, n_113, n_38, n_123, n_139, n_105, n_80, n_4, n_179, n_125, n_35, n_167, n_128, n_73, n_17, n_92, n_19, n_149, n_120, n_135, n_30, n_156, n_5, n_33, n_126, n_14, n_84, n_23, n_130, n_157, n_29, n_79, n_193, n_131, n_151, n_47, n_173, n_192, n_25, n_53, n_160, n_198, n_188, n_190, n_8, n_158, n_44, n_40, n_34, n_100, n_62, n_138, n_148, n_71, n_154, n_109, n_112, n_85, n_159, n_163, n_95, n_119, n_183, n_185, n_175, n_169, n_59, n_26, n_133, n_55, n_196, n_99, n_2, n_181, n_3, n_49, n_20, n_6, n_39, n_54, n_147, n_178, n_12, n_67, n_121, n_36, n_76, n_200, n_87, n_150, n_162, n_27, n_170, n_64, n_77, n_102, n_106, n_161, n_81, n_118, n_28, n_89, n_70, n_115, n_68, n_93, n_72, n_174, n_186, n_199, n_134, n_187, n_32, n_41, n_104, n_172, n_103, n_56, n_51, n_63, n_97, n_141, n_166, n_11, n_171, n_153, n_7, n_15, n_145, n_48, n_50, n_52, n_88, n_110, n_1938);

input n_137;
input n_168;
input n_164;
input n_191;
input n_91;
input n_82;
input n_122;
input n_194;
input n_142;
input n_176;
input n_10;
input n_140;
input n_24;
input n_124;
input n_86;
input n_136;
input n_146;
input n_182;
input n_143;
input n_83;
input n_132;
input n_61;
input n_90;
input n_127;
input n_75;
input n_101;
input n_180;
input n_184;
input n_65;
input n_78;
input n_74;
input n_144;
input n_114;
input n_57;
input n_96;
input n_37;
input n_189;
input n_165;
input n_111;
input n_108;
input n_129;
input n_31;
input n_13;
input n_66;
input n_98;
input n_177;
input n_60;
input n_155;
input n_152;
input n_197;
input n_16;
input n_43;
input n_107;
input n_0;
input n_58;
input n_9;
input n_69;
input n_18;
input n_116;
input n_195;
input n_42;
input n_22;
input n_1;
input n_45;
input n_117;
input n_46;
input n_21;
input n_94;
input n_113;
input n_38;
input n_123;
input n_139;
input n_105;
input n_80;
input n_4;
input n_179;
input n_125;
input n_35;
input n_167;
input n_128;
input n_73;
input n_17;
input n_92;
input n_19;
input n_149;
input n_120;
input n_135;
input n_30;
input n_156;
input n_5;
input n_33;
input n_126;
input n_14;
input n_84;
input n_23;
input n_130;
input n_157;
input n_29;
input n_79;
input n_193;
input n_131;
input n_151;
input n_47;
input n_173;
input n_192;
input n_25;
input n_53;
input n_160;
input n_198;
input n_188;
input n_190;
input n_8;
input n_158;
input n_44;
input n_40;
input n_34;
input n_100;
input n_62;
input n_138;
input n_148;
input n_71;
input n_154;
input n_109;
input n_112;
input n_85;
input n_159;
input n_163;
input n_95;
input n_119;
input n_183;
input n_185;
input n_175;
input n_169;
input n_59;
input n_26;
input n_133;
input n_55;
input n_196;
input n_99;
input n_2;
input n_181;
input n_3;
input n_49;
input n_20;
input n_6;
input n_39;
input n_54;
input n_147;
input n_178;
input n_12;
input n_67;
input n_121;
input n_36;
input n_76;
input n_200;
input n_87;
input n_150;
input n_162;
input n_27;
input n_170;
input n_64;
input n_77;
input n_102;
input n_106;
input n_161;
input n_81;
input n_118;
input n_28;
input n_89;
input n_70;
input n_115;
input n_68;
input n_93;
input n_72;
input n_174;
input n_186;
input n_199;
input n_134;
input n_187;
input n_32;
input n_41;
input n_104;
input n_172;
input n_103;
input n_56;
input n_51;
input n_63;
input n_97;
input n_141;
input n_166;
input n_11;
input n_171;
input n_153;
input n_7;
input n_15;
input n_145;
input n_48;
input n_50;
input n_52;
input n_88;
input n_110;

output n_1938;

wire n_924;
wire n_1263;
wire n_977;
wire n_1378;
wire n_611;
wire n_1126;
wire n_1423;
wire n_1729;
wire n_1166;
wire n_1751;
wire n_469;
wire n_1508;
wire n_785;
wire n_549;
wire n_532;
wire n_1161;
wire n_1859;
wire n_1677;
wire n_1150;
wire n_226;
wire n_1780;
wire n_1488;
wire n_667;
wire n_790;
wire n_1055;
wire n_1501;
wire n_880;
wire n_544;
wire n_1007;
wire n_552;
wire n_1528;
wire n_1370;
wire n_1292;
wire n_1198;
wire n_1360;
wire n_1099;
wire n_956;
wire n_564;
wire n_423;
wire n_1738;
wire n_1021;
wire n_551;
wire n_1323;
wire n_1466;
wire n_688;
wire n_1695;
wire n_1353;
wire n_800;
wire n_1347;
wire n_1535;
wire n_1789;
wire n_1666;
wire n_671;
wire n_819;
wire n_1451;
wire n_1022;
wire n_915;
wire n_1545;
wire n_864;
wire n_859;
wire n_951;
wire n_1264;
wire n_447;
wire n_247;
wire n_1494;
wire n_292;
wire n_625;
wire n_854;
wire n_1799;
wire n_1462;
wire n_1580;
wire n_674;
wire n_417;
wire n_1806;
wire n_516;
wire n_933;
wire n_1152;
wire n_497;
wire n_1869;
wire n_1607;
wire n_1563;
wire n_606;
wire n_275;
wire n_877;
wire n_1696;
wire n_755;
wire n_1118;
wire n_1686;
wire n_947;
wire n_1285;
wire n_373;
wire n_307;
wire n_1860;
wire n_1359;
wire n_530;
wire n_1107;
wire n_1728;
wire n_556;
wire n_1230;
wire n_668;
wire n_375;
wire n_301;
wire n_1896;
wire n_929;
wire n_1124;
wire n_1818;
wire n_902;
wire n_1576;
wire n_1104;
wire n_1294;
wire n_659;
wire n_1705;
wire n_1257;
wire n_1182;
wire n_579;
wire n_1698;
wire n_1261;
wire n_938;
wire n_1098;
wire n_320;
wire n_1154;
wire n_1242;
wire n_1135;
wire n_406;
wire n_519;
wire n_1016;
wire n_1243;
wire n_546;
wire n_1280;
wire n_1845;
wire n_281;
wire n_240;
wire n_291;
wire n_231;
wire n_257;
wire n_731;
wire n_371;
wire n_1483;
wire n_1314;
wire n_1512;
wire n_709;
wire n_1490;
wire n_317;
wire n_1236;
wire n_1633;
wire n_569;
wire n_1778;
wire n_227;
wire n_920;
wire n_1289;
wire n_1517;
wire n_335;
wire n_1669;
wire n_370;
wire n_976;
wire n_343;
wire n_1449;
wire n_308;
wire n_1566;
wire n_297;
wire n_1078;
wire n_1670;
wire n_775;
wire n_219;
wire n_600;
wire n_1484;
wire n_1374;
wire n_1328;
wire n_223;
wire n_264;
wire n_1877;
wire n_1831;
wire n_1598;
wire n_1723;
wire n_955;
wire n_1850;
wire n_339;
wire n_1146;
wire n_882;
wire n_243;
wire n_1036;
wire n_1097;
wire n_1749;
wire n_347;
wire n_550;
wire n_696;
wire n_897;
wire n_215;
wire n_350;
wire n_798;
wire n_646;
wire n_1428;
wire n_436;
wire n_1394;
wire n_1414;
wire n_1216;
wire n_290;
wire n_580;
wire n_1040;
wire n_1872;
wire n_1852;
wire n_578;
wire n_926;
wire n_344;
wire n_1218;
wire n_1931;
wire n_422;
wire n_475;
wire n_777;
wire n_1070;
wire n_1547;
wire n_1030;
wire n_1755;
wire n_415;
wire n_1071;
wire n_485;
wire n_1165;
wire n_1267;
wire n_1561;
wire n_496;
wire n_1801;
wire n_1391;
wire n_958;
wire n_1034;
wire n_670;
wire n_1513;
wire n_1600;
wire n_521;
wire n_663;
wire n_845;
wire n_1862;
wire n_673;
wire n_837;
wire n_1239;
wire n_528;
wire n_1796;
wire n_680;
wire n_1473;
wire n_1587;
wire n_395;
wire n_553;
wire n_901;
wire n_813;
wire n_1521;
wire n_1284;
wire n_1590;
wire n_214;
wire n_1748;
wire n_1672;
wire n_675;
wire n_888;
wire n_1880;
wire n_1167;
wire n_1626;
wire n_637;
wire n_1384;
wire n_1556;
wire n_446;
wire n_1863;
wire n_1064;
wire n_858;
wire n_923;
wire n_691;
wire n_1151;
wire n_881;
wire n_1405;
wire n_1706;
wire n_468;
wire n_213;
wire n_342;
wire n_464;
wire n_363;
wire n_1582;
wire n_1069;
wire n_1784;
wire n_1075;
wire n_1836;
wire n_1450;
wire n_1322;
wire n_1471;
wire n_1750;
wire n_1459;
wire n_460;
wire n_889;
wire n_973;
wire n_1700;
wire n_477;
wire n_571;
wire n_1585;
wire n_461;
wire n_1599;
wire n_1211;
wire n_1197;
wire n_1523;
wire n_907;
wire n_1447;
wire n_1377;
wire n_989;
wire n_1039;
wire n_228;
wire n_283;
wire n_1403;
wire n_488;
wire n_736;
wire n_892;
wire n_1000;
wire n_1202;
wire n_1278;
wire n_1002;
wire n_1463;
wire n_1581;
wire n_310;
wire n_593;
wire n_748;
wire n_586;
wire n_1058;
wire n_1667;
wire n_838;
wire n_332;
wire n_1053;
wire n_1224;
wire n_349;
wire n_1926;
wire n_1248;
wire n_230;
wire n_1331;
wire n_953;
wire n_279;
wire n_1014;
wire n_1241;
wire n_289;
wire n_963;
wire n_1052;
wire n_954;
wire n_627;
wire n_1385;
wire n_440;
wire n_793;
wire n_478;
wire n_1819;
wire n_476;
wire n_1527;
wire n_534;
wire n_1882;
wire n_884;
wire n_345;
wire n_944;
wire n_1754;
wire n_1623;
wire n_1854;
wire n_1565;
wire n_1809;
wire n_1856;
wire n_647;
wire n_237;
wire n_407;
wire n_1072;
wire n_832;
wire n_857;
wire n_207;
wire n_561;
wire n_1319;
wire n_1825;
wire n_1883;
wire n_1906;
wire n_1712;
wire n_1387;
wire n_1532;
wire n_1027;
wire n_971;
wire n_1156;
wire n_326;
wire n_794;
wire n_404;
wire n_686;
wire n_847;
wire n_1393;
wire n_596;
wire n_1775;
wire n_1368;
wire n_558;
wire n_702;
wire n_1276;
wire n_822;
wire n_1412;
wire n_1709;
wire n_728;
wire n_266;
wire n_1162;
wire n_272;
wire n_1538;
wire n_1838;
wire n_1199;
wire n_1847;
wire n_1779;
wire n_352;
wire n_1884;
wire n_1038;
wire n_520;
wire n_1369;
wire n_409;
wire n_1841;
wire n_1660;
wire n_887;
wire n_1905;
wire n_300;
wire n_809;
wire n_870;
wire n_931;
wire n_599;
wire n_1711;
wire n_1662;
wire n_1891;
wire n_1481;
wire n_434;
wire n_1544;
wire n_868;
wire n_639;
wire n_914;
wire n_411;
wire n_414;
wire n_1629;
wire n_1293;
wire n_965;
wire n_1876;
wire n_1743;
wire n_935;
wire n_1175;
wire n_817;
wire n_360;
wire n_1479;
wire n_1810;
wire n_1888;
wire n_759;
wire n_1892;
wire n_806;
wire n_1766;
wire n_1477;
wire n_324;
wire n_1635;
wire n_1571;
wire n_1189;
wire n_1259;
wire n_1690;
wire n_706;
wire n_746;
wire n_1649;
wire n_747;
wire n_784;
wire n_1733;
wire n_1244;
wire n_431;
wire n_1194;
wire n_1925;
wire n_1815;
wire n_615;
wire n_851;
wire n_1759;
wire n_843;
wire n_1788;
wire n_523;
wire n_913;
wire n_1537;
wire n_705;
wire n_865;
wire n_678;
wire n_697;
wire n_1222;
wire n_1679;
wire n_776;
wire n_1798;
wire n_1790;
wire n_1415;
wire n_367;
wire n_452;
wire n_525;
wire n_1260;
wire n_1746;
wire n_1647;
wire n_1829;
wire n_1464;
wire n_649;
wire n_547;
wire n_1444;
wire n_1191;
wire n_1674;
wire n_1833;
wire n_1830;
wire n_1710;
wire n_284;
wire n_1128;
wire n_1734;
wire n_744;
wire n_629;
wire n_590;
wire n_1308;
wire n_1767;
wire n_254;
wire n_1680;
wire n_1233;
wire n_1615;
wire n_1529;
wire n_526;
wire n_1916;
wire n_293;
wire n_677;
wire n_372;
wire n_244;
wire n_1333;
wire n_1121;
wire n_433;
wire n_604;
wire n_314;
wire n_368;
wire n_949;
wire n_1443;
wire n_1008;
wire n_946;
wire n_1539;
wire n_1001;
wire n_1503;
wire n_498;
wire n_1468;
wire n_1559;
wire n_1765;
wire n_1866;
wire n_689;
wire n_738;
wire n_1624;
wire n_640;
wire n_1510;
wire n_252;
wire n_624;
wire n_1380;
wire n_1744;
wire n_1617;
wire n_295;
wire n_1010;
wire n_1231;
wire n_739;
wire n_1279;
wire n_1406;
wire n_1195;
wire n_1837;
wire n_1839;
wire n_610;
wire n_1760;
wire n_936;
wire n_568;
wire n_1500;
wire n_1090;
wire n_757;
wire n_633;
wire n_439;
wire n_1832;
wire n_259;
wire n_448;
wire n_1851;
wire n_758;
wire n_999;
wire n_1933;
wire n_1656;
wire n_1158;
wire n_1509;
wire n_1874;
wire n_563;
wire n_1145;
wire n_878;
wire n_524;
wire n_204;
wire n_394;
wire n_1678;
wire n_1049;
wire n_1153;
wire n_741;
wire n_1639;
wire n_1306;
wire n_1068;
wire n_1871;
wire n_331;
wire n_906;
wire n_1163;
wire n_1207;
wire n_919;
wire n_908;
wire n_724;
wire n_1781;
wire n_658;
wire n_1740;
wire n_1362;
wire n_1586;
wire n_456;
wire n_959;
wire n_535;
wire n_940;
wire n_1445;
wire n_1492;
wire n_1923;
wire n_1773;
wire n_592;
wire n_1169;
wire n_1596;
wire n_1692;
wire n_1017;
wire n_978;
wire n_1434;
wire n_1054;
wire n_1474;
wire n_1665;
wire n_1269;
wire n_1095;
wire n_1828;
wire n_1614;
wire n_267;
wire n_514;
wire n_457;
wire n_1079;
wire n_1045;
wire n_1208;
wire n_603;
wire n_1431;
wire n_484;
wire n_1593;
wire n_1033;
wire n_442;
wire n_636;
wire n_660;
wire n_1640;
wire n_1732;
wire n_1009;
wire n_1148;
wire n_750;
wire n_742;
wire n_995;
wire n_454;
wire n_1609;
wire n_374;
wire n_396;
wire n_1887;
wire n_1383;
wire n_1073;
wire n_255;
wire n_662;
wire n_459;
wire n_218;
wire n_962;
wire n_1215;
wire n_1171;
wire n_1578;
wire n_723;
wire n_1920;
wire n_1065;
wire n_1592;
wire n_1336;
wire n_1721;
wire n_1758;
wire n_1574;
wire n_473;
wire n_1921;
wire n_1309;
wire n_1878;
wire n_1426;
wire n_1043;
wire n_355;
wire n_486;
wire n_1800;
wire n_1548;
wire n_614;
wire n_337;
wire n_1421;
wire n_1286;
wire n_1177;
wire n_1355;
wire n_974;
wire n_727;
wire n_1159;
wire n_957;
wire n_773;
wire n_208;
wire n_743;
wire n_299;
wire n_303;
wire n_296;
wire n_613;
wire n_1119;
wire n_1240;
wire n_1820;
wire n_829;
wire n_1612;
wire n_1416;
wire n_1724;
wire n_361;
wire n_700;
wire n_1237;
wire n_573;
wire n_1420;
wire n_1132;
wire n_388;
wire n_1366;
wire n_1300;
wire n_1127;
wire n_761;
wire n_1785;
wire n_1568;
wire n_1006;
wire n_329;
wire n_274;
wire n_1270;
wire n_1664;
wire n_1486;
wire n_582;
wire n_1332;
wire n_1390;
wire n_1870;
wire n_309;
wire n_512;
wire n_1591;
wire n_322;
wire n_1682;
wire n_1249;
wire n_652;
wire n_1111;
wire n_1365;
wire n_1927;
wire n_1349;
wire n_1093;
wire n_288;
wire n_1031;
wire n_263;
wire n_609;
wire n_1041;
wire n_1265;
wire n_1909;
wire n_224;
wire n_1562;
wire n_383;
wire n_834;
wire n_765;
wire n_893;
wire n_1015;
wire n_1140;
wire n_891;
wire n_1651;
wire n_239;
wire n_630;
wire n_1902;
wire n_1913;
wire n_504;
wire n_1823;
wire n_511;
wire n_874;
wire n_358;
wire n_1101;
wire n_1106;
wire n_1456;
wire n_1875;
wire n_1304;
wire n_1324;
wire n_987;
wire n_1846;
wire n_261;
wire n_1885;
wire n_1455;
wire n_767;
wire n_993;
wire n_1903;
wire n_1407;
wire n_1551;
wire n_545;
wire n_441;
wire n_860;
wire n_450;
wire n_1805;
wire n_1816;
wire n_429;
wire n_948;
wire n_1217;
wire n_628;
wire n_365;
wire n_1849;
wire n_729;
wire n_1131;
wire n_1084;
wire n_970;
wire n_1935;
wire n_911;
wire n_1430;
wire n_513;
wire n_1094;
wire n_1354;
wire n_560;
wire n_1534;
wire n_340;
wire n_1351;
wire n_1044;
wire n_1205;
wire n_346;
wire n_1209;
wire n_1552;
wire n_495;
wire n_602;
wire n_574;
wire n_1435;
wire n_879;
wire n_623;
wire n_405;
wire n_824;
wire n_359;
wire n_1645;
wire n_490;
wire n_1327;
wire n_996;
wire n_921;
wire n_1684;
wire n_233;
wire n_1717;
wire n_572;
wire n_366;
wire n_815;
wire n_1795;
wire n_1821;
wire n_327;
wire n_1381;
wire n_1611;
wire n_1037;
wire n_1080;
wire n_1274;
wire n_1316;
wire n_1708;
wire n_426;
wire n_1438;
wire n_1082;
wire n_1840;
wire n_589;
wire n_716;
wire n_1630;
wire n_562;
wire n_1436;
wire n_1691;
wire n_952;
wire n_1229;
wire n_391;
wire n_701;
wire n_1437;
wire n_1023;
wire n_645;
wire n_539;
wire n_803;
wire n_1092;
wire n_238;
wire n_1776;
wire n_531;
wire n_1757;
wire n_890;
wire n_1897;
wire n_764;
wire n_1919;
wire n_1056;
wire n_1424;
wire n_960;
wire n_1893;
wire n_222;
wire n_1290;
wire n_1123;
wire n_1467;
wire n_1047;
wire n_634;
wire n_1252;
wire n_348;
wire n_1382;
wire n_1029;
wire n_925;
wire n_1206;
wire n_424;
wire n_1311;
wire n_1519;
wire n_256;
wire n_950;
wire n_1553;
wire n_1811;
wire n_380;
wire n_419;
wire n_1346;
wire n_444;
wire n_1299;
wire n_1808;
wire n_1060;
wire n_1141;
wire n_316;
wire n_389;
wire n_418;
wire n_248;
wire n_912;
wire n_315;
wire n_968;
wire n_451;
wire n_619;
wire n_408;
wire n_1386;
wire n_1699;
wire n_376;
wire n_967;
wire n_1442;
wire n_1139;
wire n_515;
wire n_351;
wire n_885;
wire n_397;
wire n_1432;
wire n_1357;
wire n_483;
wire n_683;
wire n_1632;
wire n_1057;
wire n_1051;
wire n_1085;
wire n_1066;
wire n_721;
wire n_1157;
wire n_841;
wire n_1050;
wire n_802;
wire n_1608;
wire n_983;
wire n_1844;
wire n_280;
wire n_1305;
wire n_873;
wire n_1826;
wire n_378;
wire n_1112;
wire n_762;
wire n_1283;
wire n_1644;
wire n_690;
wire n_583;
wire n_302;
wire n_1343;
wire n_1203;
wire n_1631;
wire n_821;
wire n_1763;
wire n_1768;
wire n_321;
wire n_1179;
wire n_621;
wire n_753;
wire n_455;
wire n_1048;
wire n_1719;
wire n_1288;
wire n_212;
wire n_385;
wire n_507;
wire n_1560;
wire n_1605;
wire n_330;
wire n_1228;
wire n_972;
wire n_692;
wire n_820;
wire n_1200;
wire n_1911;
wire n_1301;
wire n_1363;
wire n_1668;
wire n_1185;
wire n_991;
wire n_828;
wire n_779;
wire n_576;
wire n_1143;
wire n_1579;
wire n_1329;
wire n_1312;
wire n_1439;
wire n_804;
wire n_537;
wire n_1688;
wire n_945;
wire n_492;
wire n_1504;
wire n_943;
wire n_341;
wire n_250;
wire n_992;
wire n_1932;
wire n_543;
wire n_260;
wire n_842;
wire n_650;
wire n_984;
wire n_694;
wire n_286;
wire n_1643;
wire n_883;
wire n_470;
wire n_449;
wire n_325;
wire n_1594;
wire n_1214;
wire n_1342;
wire n_1400;
wire n_900;
wire n_856;
wire n_1793;
wire n_918;
wire n_942;
wire n_1804;
wire n_1147;
wire n_1557;
wire n_1610;
wire n_1077;
wire n_1422;
wire n_540;
wire n_618;
wire n_896;
wire n_323;
wire n_356;
wire n_894;
wire n_1636;
wire n_1730;
wire n_831;
wire n_964;
wire n_1373;
wire n_1350;
wire n_1511;
wire n_1865;
wire n_1470;
wire n_1096;
wire n_234;
wire n_1575;
wire n_1697;
wire n_1735;
wire n_833;
wire n_1646;
wire n_225;
wire n_1307;
wire n_1881;
wire n_988;
wire n_814;
wire n_1549;
wire n_1934;
wire n_1201;
wire n_1114;
wire n_655;
wire n_1616;
wire n_1446;
wire n_669;
wire n_472;
wire n_1458;
wire n_1176;
wire n_1472;
wire n_1807;
wire n_387;
wire n_1149;
wire n_398;
wire n_1671;
wire n_635;
wire n_763;
wire n_1020;
wire n_1062;
wire n_211;
wire n_1824;
wire n_1917;
wire n_1219;
wire n_1204;
wire n_1814;
wire n_1035;
wire n_287;
wire n_555;
wire n_783;
wire n_1848;
wire n_1928;
wire n_1188;
wire n_1722;
wire n_661;
wire n_1802;
wire n_849;
wire n_584;
wire n_681;
wire n_336;
wire n_1638;
wire n_1786;
wire n_430;
wire n_510;
wire n_216;
wire n_311;
wire n_830;
wire n_1296;
wire n_1413;
wire n_801;
wire n_241;
wire n_875;
wire n_357;
wire n_1110;
wire n_1655;
wire n_445;
wire n_749;
wire n_1895;
wire n_1134;
wire n_1358;
wire n_717;
wire n_939;
wire n_482;
wire n_1088;
wire n_588;
wire n_1173;
wire n_789;
wire n_1232;
wire n_1603;
wire n_734;
wire n_638;
wire n_866;
wire n_969;
wire n_1401;
wire n_1019;
wire n_1105;
wire n_249;
wire n_304;
wire n_1338;
wire n_577;
wire n_1522;
wire n_1687;
wire n_1637;
wire n_1419;
wire n_338;
wire n_1653;
wire n_693;
wire n_1506;
wire n_836;
wire n_990;
wire n_1886;
wire n_1389;
wire n_1894;
wire n_975;
wire n_1908;
wire n_1256;
wire n_1702;
wire n_567;
wire n_1465;
wire n_778;
wire n_1122;
wire n_306;
wire n_458;
wire n_770;
wire n_1375;
wire n_1102;
wire n_1843;
wire n_711;
wire n_1499;
wire n_1187;
wire n_1441;
wire n_1392;
wire n_1597;
wire n_1929;
wire n_1164;
wire n_1659;
wire n_1834;
wire n_489;
wire n_1174;
wire n_1371;
wire n_617;
wire n_1303;
wire n_1572;
wire n_876;
wire n_1516;
wire n_1190;
wire n_1736;
wire n_1685;
wire n_601;
wire n_917;
wire n_1714;
wire n_966;
wire n_253;
wire n_1116;
wire n_1661;
wire n_1212;
wire n_1541;
wire n_206;
wire n_217;
wire n_726;
wire n_982;
wire n_1573;
wire n_1453;
wire n_1731;
wire n_818;
wire n_861;
wire n_1713;
wire n_1183;
wire n_1658;
wire n_899;
wire n_1253;
wire n_210;
wire n_1737;
wire n_1904;
wire n_774;
wire n_1628;
wire n_1335;
wire n_1514;
wire n_1777;
wire n_1059;
wire n_1345;
wire n_1133;
wire n_1771;
wire n_1912;
wire n_1899;
wire n_557;
wire n_1410;
wire n_1005;
wire n_607;
wire n_1003;
wire n_679;
wire n_710;
wire n_527;
wire n_1168;
wire n_707;
wire n_937;
wire n_1427;
wire n_393;
wire n_487;
wire n_1584;
wire n_665;
wire n_1835;
wire n_1726;
wire n_1440;
wire n_421;
wire n_1853;
wire n_1356;
wire n_1787;
wire n_910;
wire n_1657;
wire n_768;
wire n_1475;
wire n_1302;
wire n_1774;
wire n_1725;
wire n_205;
wire n_1136;
wire n_1313;
wire n_1491;
wire n_754;
wire n_1496;
wire n_1125;
wire n_410;
wire n_708;
wire n_529;
wire n_1812;
wire n_735;
wire n_232;
wire n_1915;
wire n_1109;
wire n_895;
wire n_1310;
wire n_1803;
wire n_202;
wire n_427;
wire n_1399;
wire n_1543;
wire n_791;
wire n_732;
wire n_1533;
wire n_808;
wire n_797;
wire n_1025;
wire n_1930;
wire n_500;
wire n_1067;
wire n_1720;
wire n_435;
wire n_766;
wire n_1457;
wire n_541;
wire n_538;
wire n_1117;
wire n_799;
wire n_687;
wire n_715;
wire n_1742;
wire n_1480;
wire n_1482;
wire n_1213;
wire n_1266;
wire n_536;
wire n_872;
wire n_594;
wire n_1291;
wire n_1297;
wire n_1753;
wire n_1782;
wire n_1155;
wire n_1418;
wire n_1524;
wire n_1689;
wire n_1485;
wire n_1011;
wire n_1184;
wire n_985;
wire n_1855;
wire n_869;
wire n_810;
wire n_416;
wire n_827;
wire n_401;
wire n_1703;
wire n_1352;
wire n_626;
wire n_1650;
wire n_1144;
wire n_1137;
wire n_1570;
wire n_1170;
wire n_305;
wire n_676;
wire n_294;
wire n_318;
wire n_653;
wire n_642;
wire n_1602;
wire n_855;
wire n_1178;
wire n_1461;
wire n_850;
wire n_684;
wire n_268;
wire n_664;
wire n_503;
wire n_235;
wire n_1372;
wire n_605;
wire n_1273;
wire n_1822;
wire n_353;
wire n_620;
wire n_643;
wire n_916;
wire n_1081;
wire n_493;
wire n_1235;
wire n_703;
wire n_698;
wire n_980;
wire n_1115;
wire n_1282;
wire n_1318;
wire n_1783;
wire n_780;
wire n_998;
wire n_1454;
wire n_467;
wire n_1227;
wire n_1531;
wire n_840;
wire n_1334;
wire n_1907;
wire n_501;
wire n_823;
wire n_245;
wire n_725;
wire n_1388;
wire n_1417;
wire n_1295;
wire n_672;
wire n_1898;
wire n_581;
wire n_382;
wire n_554;
wire n_1625;
wire n_898;
wire n_1762;
wire n_1013;
wire n_1452;
wire n_718;
wire n_265;
wire n_1120;
wire n_719;
wire n_443;
wire n_1791;
wire n_1890;
wire n_1747;
wire n_714;
wire n_1683;
wire n_1817;
wire n_909;
wire n_1530;
wire n_1497;
wire n_997;
wire n_932;
wire n_612;
wire n_1409;
wire n_788;
wire n_1326;
wire n_1268;
wire n_559;
wire n_825;
wire n_508;
wire n_506;
wire n_1320;
wire n_1663;
wire n_737;
wire n_1718;
wire n_986;
wire n_509;
wire n_1317;
wire n_1518;
wire n_1715;
wire n_1281;
wire n_1192;
wire n_1024;
wire n_1063;
wire n_1889;
wire n_209;
wire n_1792;
wire n_1564;
wire n_1868;
wire n_1613;
wire n_733;
wire n_1489;
wire n_1922;
wire n_1376;
wire n_941;
wire n_981;
wire n_1569;
wire n_867;
wire n_587;
wire n_792;
wire n_756;
wire n_1429;
wire n_399;
wire n_1238;
wire n_548;
wire n_812;
wire n_298;
wire n_518;
wire n_505;
wire n_1772;
wire n_282;
wire n_752;
wire n_905;
wire n_1476;
wire n_1108;
wire n_782;
wire n_1100;
wire n_1861;
wire n_1395;
wire n_862;
wire n_1425;
wire n_760;
wire n_1901;
wire n_1900;
wire n_1620;
wire n_381;
wire n_220;
wire n_390;
wire n_1330;
wire n_1867;
wire n_481;
wire n_1675;
wire n_1924;
wire n_1727;
wire n_1554;
wire n_1745;
wire n_769;
wire n_1046;
wire n_271;
wire n_934;
wire n_1618;
wire n_826;
wire n_1813;
wire n_886;
wire n_1221;
wire n_654;
wire n_1172;
wire n_379;
wire n_428;
wire n_1341;
wire n_570;
wire n_1641;
wire n_1361;
wire n_1707;
wire n_853;
wire n_377;
wire n_751;
wire n_786;
wire n_1083;
wire n_1142;
wire n_1129;
wire n_392;
wire n_704;
wire n_787;
wire n_1770;
wire n_961;
wire n_1756;
wire n_771;
wire n_276;
wire n_1716;
wire n_1225;
wire n_1520;
wire n_522;
wire n_1287;
wire n_1262;
wire n_400;
wire n_930;
wire n_1873;
wire n_1411;
wire n_221;
wire n_622;
wire n_1577;
wire n_1087;
wire n_386;
wire n_994;
wire n_1701;
wire n_848;
wire n_1550;
wire n_1498;
wire n_1223;
wire n_1272;
wire n_682;
wire n_1567;
wire n_1247;
wire n_922;
wire n_816;
wire n_1648;
wire n_591;
wire n_1536;
wire n_1857;
wire n_1344;
wire n_313;
wire n_631;
wire n_479;
wire n_1246;
wire n_1339;
wire n_1478;
wire n_1797;
wire n_432;
wire n_1769;
wire n_839;
wire n_1210;
wire n_1364;
wire n_328;
wire n_1250;
wire n_369;
wire n_1842;
wire n_871;
wire n_598;
wire n_685;
wire n_928;
wire n_608;
wire n_1367;
wire n_1460;
wire n_772;
wire n_1555;
wire n_499;
wire n_1589;
wire n_517;
wire n_402;
wire n_413;
wire n_1086;
wire n_796;
wire n_1858;
wire n_1619;
wire n_236;
wire n_1502;
wire n_1469;
wire n_1012;
wire n_1396;
wire n_1348;
wire n_903;
wire n_1525;
wire n_1752;
wire n_740;
wire n_203;
wire n_384;
wire n_1404;
wire n_1794;
wire n_1315;
wire n_277;
wire n_1061;
wire n_1910;
wire n_333;
wire n_1298;
wire n_1652;
wire n_462;
wire n_1193;
wire n_1676;
wire n_1255;
wire n_258;
wire n_1113;
wire n_1226;
wire n_722;
wire n_1277;
wire n_844;
wire n_201;
wire n_471;
wire n_852;
wire n_1487;
wire n_1864;
wire n_1028;
wire n_1601;
wire n_781;
wire n_474;
wire n_542;
wire n_463;
wire n_1546;
wire n_595;
wire n_502;
wire n_466;
wire n_420;
wire n_1337;
wire n_1495;
wire n_632;
wire n_699;
wire n_979;
wire n_1515;
wire n_1627;
wire n_1245;
wire n_846;
wire n_1673;
wire n_465;
wire n_362;
wire n_1321;
wire n_273;
wire n_1937;
wire n_585;
wire n_1739;
wire n_270;
wire n_616;
wire n_1914;
wire n_745;
wire n_1654;
wire n_1103;
wire n_648;
wire n_1379;
wire n_312;
wire n_1076;
wire n_1091;
wire n_1408;
wire n_494;
wire n_1761;
wire n_641;
wire n_730;
wire n_1325;
wire n_1595;
wire n_354;
wire n_575;
wire n_480;
wire n_425;
wire n_795;
wire n_695;
wire n_656;
wire n_1606;
wire n_1220;
wire n_1694;
wire n_1540;
wire n_229;
wire n_1936;
wire n_437;
wire n_1642;
wire n_403;
wire n_453;
wire n_1130;
wire n_720;
wire n_1918;
wire n_1526;
wire n_863;
wire n_805;
wire n_1604;
wire n_1275;
wire n_1764;
wire n_712;
wire n_246;
wire n_1583;
wire n_1042;
wire n_1402;
wire n_269;
wire n_285;
wire n_412;
wire n_1493;
wire n_657;
wire n_644;
wire n_1741;
wire n_1160;
wire n_1397;
wire n_491;
wire n_1258;
wire n_1074;
wire n_1621;
wire n_251;
wire n_566;
wire n_565;
wire n_1448;
wire n_1507;
wire n_1398;
wire n_1879;
wire n_597;
wire n_1181;
wire n_1505;
wire n_1634;
wire n_1196;
wire n_651;
wire n_1340;
wire n_334;
wire n_811;
wire n_1558;
wire n_807;
wire n_835;
wire n_666;
wire n_262;
wire n_1433;
wire n_1704;
wire n_1254;
wire n_1026;
wire n_1234;
wire n_319;
wire n_364;
wire n_1138;
wire n_927;
wire n_1089;
wire n_1004;
wire n_1186;
wire n_1032;
wire n_242;
wire n_1681;
wire n_1018;
wire n_1693;
wire n_438;
wire n_713;
wire n_904;
wire n_1588;
wire n_1622;
wire n_1180;
wire n_1827;
wire n_1271;
wire n_533;
wire n_1542;
wire n_1251;
wire n_278;

INVx1_ASAP7_75t_L g201 ( 
.A(n_31),
.Y(n_201)
);

CKINVDCx5p33_ASAP7_75t_R g202 ( 
.A(n_5),
.Y(n_202)
);

CKINVDCx5p33_ASAP7_75t_R g203 ( 
.A(n_176),
.Y(n_203)
);

CKINVDCx5p33_ASAP7_75t_R g204 ( 
.A(n_93),
.Y(n_204)
);

CKINVDCx5p33_ASAP7_75t_R g205 ( 
.A(n_139),
.Y(n_205)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_52),
.Y(n_206)
);

BUFx10_ASAP7_75t_L g207 ( 
.A(n_65),
.Y(n_207)
);

CKINVDCx20_ASAP7_75t_R g208 ( 
.A(n_43),
.Y(n_208)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_148),
.Y(n_209)
);

BUFx6f_ASAP7_75t_L g210 ( 
.A(n_17),
.Y(n_210)
);

CKINVDCx5p33_ASAP7_75t_R g211 ( 
.A(n_75),
.Y(n_211)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_42),
.Y(n_212)
);

CKINVDCx5p33_ASAP7_75t_R g213 ( 
.A(n_135),
.Y(n_213)
);

CKINVDCx5p33_ASAP7_75t_R g214 ( 
.A(n_140),
.Y(n_214)
);

CKINVDCx5p33_ASAP7_75t_R g215 ( 
.A(n_54),
.Y(n_215)
);

CKINVDCx5p33_ASAP7_75t_R g216 ( 
.A(n_142),
.Y(n_216)
);

BUFx3_ASAP7_75t_L g217 ( 
.A(n_161),
.Y(n_217)
);

CKINVDCx5p33_ASAP7_75t_R g218 ( 
.A(n_178),
.Y(n_218)
);

CKINVDCx5p33_ASAP7_75t_R g219 ( 
.A(n_8),
.Y(n_219)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_134),
.Y(n_220)
);

BUFx2_ASAP7_75t_L g221 ( 
.A(n_98),
.Y(n_221)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_153),
.Y(n_222)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_5),
.Y(n_223)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_124),
.Y(n_224)
);

CKINVDCx20_ASAP7_75t_R g225 ( 
.A(n_193),
.Y(n_225)
);

CKINVDCx5p33_ASAP7_75t_R g226 ( 
.A(n_17),
.Y(n_226)
);

CKINVDCx5p33_ASAP7_75t_R g227 ( 
.A(n_184),
.Y(n_227)
);

BUFx6f_ASAP7_75t_L g228 ( 
.A(n_188),
.Y(n_228)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_159),
.Y(n_229)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_152),
.Y(n_230)
);

BUFx3_ASAP7_75t_L g231 ( 
.A(n_14),
.Y(n_231)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_137),
.Y(n_232)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_187),
.Y(n_233)
);

CKINVDCx5p33_ASAP7_75t_R g234 ( 
.A(n_106),
.Y(n_234)
);

CKINVDCx5p33_ASAP7_75t_R g235 ( 
.A(n_27),
.Y(n_235)
);

CKINVDCx20_ASAP7_75t_R g236 ( 
.A(n_44),
.Y(n_236)
);

CKINVDCx5p33_ASAP7_75t_R g237 ( 
.A(n_121),
.Y(n_237)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_118),
.Y(n_238)
);

CKINVDCx5p33_ASAP7_75t_R g239 ( 
.A(n_100),
.Y(n_239)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_70),
.Y(n_240)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_130),
.Y(n_241)
);

INVxp33_ASAP7_75t_R g242 ( 
.A(n_13),
.Y(n_242)
);

CKINVDCx5p33_ASAP7_75t_R g243 ( 
.A(n_198),
.Y(n_243)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_81),
.Y(n_244)
);

CKINVDCx5p33_ASAP7_75t_R g245 ( 
.A(n_63),
.Y(n_245)
);

CKINVDCx5p33_ASAP7_75t_R g246 ( 
.A(n_92),
.Y(n_246)
);

CKINVDCx5p33_ASAP7_75t_R g247 ( 
.A(n_122),
.Y(n_247)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_136),
.Y(n_248)
);

INVx1_ASAP7_75t_SL g249 ( 
.A(n_115),
.Y(n_249)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_119),
.Y(n_250)
);

CKINVDCx5p33_ASAP7_75t_R g251 ( 
.A(n_23),
.Y(n_251)
);

CKINVDCx20_ASAP7_75t_R g252 ( 
.A(n_156),
.Y(n_252)
);

CKINVDCx5p33_ASAP7_75t_R g253 ( 
.A(n_46),
.Y(n_253)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_50),
.Y(n_254)
);

CKINVDCx5p33_ASAP7_75t_R g255 ( 
.A(n_62),
.Y(n_255)
);

CKINVDCx20_ASAP7_75t_R g256 ( 
.A(n_99),
.Y(n_256)
);

BUFx6f_ASAP7_75t_L g257 ( 
.A(n_149),
.Y(n_257)
);

BUFx10_ASAP7_75t_L g258 ( 
.A(n_12),
.Y(n_258)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_24),
.Y(n_259)
);

BUFx3_ASAP7_75t_L g260 ( 
.A(n_78),
.Y(n_260)
);

CKINVDCx5p33_ASAP7_75t_R g261 ( 
.A(n_175),
.Y(n_261)
);

CKINVDCx5p33_ASAP7_75t_R g262 ( 
.A(n_40),
.Y(n_262)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_172),
.Y(n_263)
);

CKINVDCx16_ASAP7_75t_R g264 ( 
.A(n_47),
.Y(n_264)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_123),
.Y(n_265)
);

CKINVDCx5p33_ASAP7_75t_R g266 ( 
.A(n_18),
.Y(n_266)
);

CKINVDCx5p33_ASAP7_75t_R g267 ( 
.A(n_104),
.Y(n_267)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_33),
.Y(n_268)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_90),
.Y(n_269)
);

CKINVDCx5p33_ASAP7_75t_R g270 ( 
.A(n_66),
.Y(n_270)
);

CKINVDCx5p33_ASAP7_75t_R g271 ( 
.A(n_27),
.Y(n_271)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_52),
.Y(n_272)
);

BUFx3_ASAP7_75t_L g273 ( 
.A(n_189),
.Y(n_273)
);

CKINVDCx5p33_ASAP7_75t_R g274 ( 
.A(n_62),
.Y(n_274)
);

CKINVDCx5p33_ASAP7_75t_R g275 ( 
.A(n_186),
.Y(n_275)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_117),
.Y(n_276)
);

CKINVDCx5p33_ASAP7_75t_R g277 ( 
.A(n_197),
.Y(n_277)
);

INVx2_ASAP7_75t_L g278 ( 
.A(n_108),
.Y(n_278)
);

CKINVDCx5p33_ASAP7_75t_R g279 ( 
.A(n_132),
.Y(n_279)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_77),
.Y(n_280)
);

CKINVDCx20_ASAP7_75t_R g281 ( 
.A(n_170),
.Y(n_281)
);

CKINVDCx5p33_ASAP7_75t_R g282 ( 
.A(n_191),
.Y(n_282)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_20),
.Y(n_283)
);

CKINVDCx5p33_ASAP7_75t_R g284 ( 
.A(n_110),
.Y(n_284)
);

CKINVDCx5p33_ASAP7_75t_R g285 ( 
.A(n_25),
.Y(n_285)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_15),
.Y(n_286)
);

CKINVDCx5p33_ASAP7_75t_R g287 ( 
.A(n_73),
.Y(n_287)
);

CKINVDCx5p33_ASAP7_75t_R g288 ( 
.A(n_8),
.Y(n_288)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_0),
.Y(n_289)
);

CKINVDCx5p33_ASAP7_75t_R g290 ( 
.A(n_19),
.Y(n_290)
);

CKINVDCx5p33_ASAP7_75t_R g291 ( 
.A(n_138),
.Y(n_291)
);

BUFx6f_ASAP7_75t_L g292 ( 
.A(n_80),
.Y(n_292)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_60),
.Y(n_293)
);

INVx2_ASAP7_75t_L g294 ( 
.A(n_96),
.Y(n_294)
);

CKINVDCx12_ASAP7_75t_R g295 ( 
.A(n_22),
.Y(n_295)
);

CKINVDCx5p33_ASAP7_75t_R g296 ( 
.A(n_127),
.Y(n_296)
);

CKINVDCx20_ASAP7_75t_R g297 ( 
.A(n_171),
.Y(n_297)
);

CKINVDCx5p33_ASAP7_75t_R g298 ( 
.A(n_38),
.Y(n_298)
);

INVx2_ASAP7_75t_L g299 ( 
.A(n_146),
.Y(n_299)
);

CKINVDCx5p33_ASAP7_75t_R g300 ( 
.A(n_95),
.Y(n_300)
);

CKINVDCx5p33_ASAP7_75t_R g301 ( 
.A(n_35),
.Y(n_301)
);

CKINVDCx20_ASAP7_75t_R g302 ( 
.A(n_154),
.Y(n_302)
);

CKINVDCx20_ASAP7_75t_R g303 ( 
.A(n_84),
.Y(n_303)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_164),
.Y(n_304)
);

INVx2_ASAP7_75t_L g305 ( 
.A(n_50),
.Y(n_305)
);

CKINVDCx20_ASAP7_75t_R g306 ( 
.A(n_199),
.Y(n_306)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_85),
.Y(n_307)
);

CKINVDCx5p33_ASAP7_75t_R g308 ( 
.A(n_20),
.Y(n_308)
);

CKINVDCx20_ASAP7_75t_R g309 ( 
.A(n_194),
.Y(n_309)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_141),
.Y(n_310)
);

CKINVDCx5p33_ASAP7_75t_R g311 ( 
.A(n_30),
.Y(n_311)
);

CKINVDCx5p33_ASAP7_75t_R g312 ( 
.A(n_64),
.Y(n_312)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_47),
.Y(n_313)
);

CKINVDCx20_ASAP7_75t_R g314 ( 
.A(n_59),
.Y(n_314)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_177),
.Y(n_315)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_112),
.Y(n_316)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_12),
.Y(n_317)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_6),
.Y(n_318)
);

CKINVDCx5p33_ASAP7_75t_R g319 ( 
.A(n_91),
.Y(n_319)
);

CKINVDCx5p33_ASAP7_75t_R g320 ( 
.A(n_35),
.Y(n_320)
);

CKINVDCx20_ASAP7_75t_R g321 ( 
.A(n_94),
.Y(n_321)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_46),
.Y(n_322)
);

CKINVDCx20_ASAP7_75t_R g323 ( 
.A(n_174),
.Y(n_323)
);

CKINVDCx5p33_ASAP7_75t_R g324 ( 
.A(n_30),
.Y(n_324)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_200),
.Y(n_325)
);

CKINVDCx14_ASAP7_75t_R g326 ( 
.A(n_150),
.Y(n_326)
);

CKINVDCx5p33_ASAP7_75t_R g327 ( 
.A(n_155),
.Y(n_327)
);

CKINVDCx5p33_ASAP7_75t_R g328 ( 
.A(n_87),
.Y(n_328)
);

CKINVDCx5p33_ASAP7_75t_R g329 ( 
.A(n_107),
.Y(n_329)
);

CKINVDCx5p33_ASAP7_75t_R g330 ( 
.A(n_165),
.Y(n_330)
);

CKINVDCx5p33_ASAP7_75t_R g331 ( 
.A(n_59),
.Y(n_331)
);

CKINVDCx5p33_ASAP7_75t_R g332 ( 
.A(n_42),
.Y(n_332)
);

CKINVDCx20_ASAP7_75t_R g333 ( 
.A(n_160),
.Y(n_333)
);

BUFx10_ASAP7_75t_L g334 ( 
.A(n_45),
.Y(n_334)
);

CKINVDCx5p33_ASAP7_75t_R g335 ( 
.A(n_61),
.Y(n_335)
);

CKINVDCx5p33_ASAP7_75t_R g336 ( 
.A(n_79),
.Y(n_336)
);

BUFx3_ASAP7_75t_L g337 ( 
.A(n_61),
.Y(n_337)
);

CKINVDCx5p33_ASAP7_75t_R g338 ( 
.A(n_38),
.Y(n_338)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_76),
.Y(n_339)
);

CKINVDCx5p33_ASAP7_75t_R g340 ( 
.A(n_39),
.Y(n_340)
);

CKINVDCx5p33_ASAP7_75t_R g341 ( 
.A(n_39),
.Y(n_341)
);

INVx1_ASAP7_75t_L g342 ( 
.A(n_26),
.Y(n_342)
);

CKINVDCx5p33_ASAP7_75t_R g343 ( 
.A(n_69),
.Y(n_343)
);

BUFx2_ASAP7_75t_L g344 ( 
.A(n_41),
.Y(n_344)
);

INVx2_ASAP7_75t_SL g345 ( 
.A(n_101),
.Y(n_345)
);

CKINVDCx5p33_ASAP7_75t_R g346 ( 
.A(n_10),
.Y(n_346)
);

CKINVDCx5p33_ASAP7_75t_R g347 ( 
.A(n_168),
.Y(n_347)
);

INVx1_ASAP7_75t_L g348 ( 
.A(n_33),
.Y(n_348)
);

CKINVDCx5p33_ASAP7_75t_R g349 ( 
.A(n_26),
.Y(n_349)
);

CKINVDCx5p33_ASAP7_75t_R g350 ( 
.A(n_40),
.Y(n_350)
);

INVx1_ASAP7_75t_L g351 ( 
.A(n_71),
.Y(n_351)
);

CKINVDCx5p33_ASAP7_75t_R g352 ( 
.A(n_180),
.Y(n_352)
);

BUFx10_ASAP7_75t_L g353 ( 
.A(n_128),
.Y(n_353)
);

CKINVDCx5p33_ASAP7_75t_R g354 ( 
.A(n_72),
.Y(n_354)
);

CKINVDCx5p33_ASAP7_75t_R g355 ( 
.A(n_157),
.Y(n_355)
);

CKINVDCx5p33_ASAP7_75t_R g356 ( 
.A(n_133),
.Y(n_356)
);

CKINVDCx5p33_ASAP7_75t_R g357 ( 
.A(n_0),
.Y(n_357)
);

BUFx10_ASAP7_75t_L g358 ( 
.A(n_55),
.Y(n_358)
);

CKINVDCx5p33_ASAP7_75t_R g359 ( 
.A(n_24),
.Y(n_359)
);

INVx1_ASAP7_75t_L g360 ( 
.A(n_67),
.Y(n_360)
);

CKINVDCx5p33_ASAP7_75t_R g361 ( 
.A(n_9),
.Y(n_361)
);

CKINVDCx5p33_ASAP7_75t_R g362 ( 
.A(n_162),
.Y(n_362)
);

CKINVDCx5p33_ASAP7_75t_R g363 ( 
.A(n_125),
.Y(n_363)
);

CKINVDCx5p33_ASAP7_75t_R g364 ( 
.A(n_21),
.Y(n_364)
);

CKINVDCx5p33_ASAP7_75t_R g365 ( 
.A(n_34),
.Y(n_365)
);

CKINVDCx5p33_ASAP7_75t_R g366 ( 
.A(n_145),
.Y(n_366)
);

CKINVDCx20_ASAP7_75t_R g367 ( 
.A(n_53),
.Y(n_367)
);

CKINVDCx5p33_ASAP7_75t_R g368 ( 
.A(n_163),
.Y(n_368)
);

CKINVDCx5p33_ASAP7_75t_R g369 ( 
.A(n_54),
.Y(n_369)
);

CKINVDCx5p33_ASAP7_75t_R g370 ( 
.A(n_88),
.Y(n_370)
);

INVx2_ASAP7_75t_L g371 ( 
.A(n_143),
.Y(n_371)
);

CKINVDCx5p33_ASAP7_75t_R g372 ( 
.A(n_102),
.Y(n_372)
);

INVx1_ASAP7_75t_L g373 ( 
.A(n_181),
.Y(n_373)
);

CKINVDCx5p33_ASAP7_75t_R g374 ( 
.A(n_4),
.Y(n_374)
);

INVx1_ASAP7_75t_L g375 ( 
.A(n_185),
.Y(n_375)
);

CKINVDCx5p33_ASAP7_75t_R g376 ( 
.A(n_14),
.Y(n_376)
);

INVx1_ASAP7_75t_L g377 ( 
.A(n_147),
.Y(n_377)
);

INVx1_ASAP7_75t_L g378 ( 
.A(n_25),
.Y(n_378)
);

BUFx2_ASAP7_75t_L g379 ( 
.A(n_89),
.Y(n_379)
);

INVx3_ASAP7_75t_L g380 ( 
.A(n_179),
.Y(n_380)
);

CKINVDCx5p33_ASAP7_75t_R g381 ( 
.A(n_97),
.Y(n_381)
);

INVx2_ASAP7_75t_L g382 ( 
.A(n_45),
.Y(n_382)
);

CKINVDCx5p33_ASAP7_75t_R g383 ( 
.A(n_167),
.Y(n_383)
);

CKINVDCx5p33_ASAP7_75t_R g384 ( 
.A(n_196),
.Y(n_384)
);

CKINVDCx5p33_ASAP7_75t_R g385 ( 
.A(n_18),
.Y(n_385)
);

INVx3_ASAP7_75t_L g386 ( 
.A(n_83),
.Y(n_386)
);

CKINVDCx5p33_ASAP7_75t_R g387 ( 
.A(n_129),
.Y(n_387)
);

INVx1_ASAP7_75t_L g388 ( 
.A(n_36),
.Y(n_388)
);

INVx1_ASAP7_75t_L g389 ( 
.A(n_37),
.Y(n_389)
);

INVx1_ASAP7_75t_L g390 ( 
.A(n_48),
.Y(n_390)
);

CKINVDCx5p33_ASAP7_75t_R g391 ( 
.A(n_32),
.Y(n_391)
);

CKINVDCx5p33_ASAP7_75t_R g392 ( 
.A(n_43),
.Y(n_392)
);

INVx2_ASAP7_75t_SL g393 ( 
.A(n_44),
.Y(n_393)
);

INVx1_ASAP7_75t_L g394 ( 
.A(n_173),
.Y(n_394)
);

INVx2_ASAP7_75t_L g395 ( 
.A(n_22),
.Y(n_395)
);

INVx1_ASAP7_75t_L g396 ( 
.A(n_34),
.Y(n_396)
);

CKINVDCx5p33_ASAP7_75t_R g397 ( 
.A(n_166),
.Y(n_397)
);

CKINVDCx5p33_ASAP7_75t_R g398 ( 
.A(n_109),
.Y(n_398)
);

CKINVDCx5p33_ASAP7_75t_R g399 ( 
.A(n_86),
.Y(n_399)
);

CKINVDCx5p33_ASAP7_75t_R g400 ( 
.A(n_7),
.Y(n_400)
);

INVx2_ASAP7_75t_SL g401 ( 
.A(n_28),
.Y(n_401)
);

CKINVDCx5p33_ASAP7_75t_R g402 ( 
.A(n_264),
.Y(n_402)
);

INVx1_ASAP7_75t_L g403 ( 
.A(n_210),
.Y(n_403)
);

CKINVDCx5p33_ASAP7_75t_R g404 ( 
.A(n_251),
.Y(n_404)
);

CKINVDCx5p33_ASAP7_75t_R g405 ( 
.A(n_253),
.Y(n_405)
);

CKINVDCx20_ASAP7_75t_R g406 ( 
.A(n_225),
.Y(n_406)
);

CKINVDCx5p33_ASAP7_75t_R g407 ( 
.A(n_255),
.Y(n_407)
);

CKINVDCx20_ASAP7_75t_R g408 ( 
.A(n_252),
.Y(n_408)
);

CKINVDCx20_ASAP7_75t_R g409 ( 
.A(n_256),
.Y(n_409)
);

BUFx3_ASAP7_75t_L g410 ( 
.A(n_217),
.Y(n_410)
);

CKINVDCx5p33_ASAP7_75t_R g411 ( 
.A(n_262),
.Y(n_411)
);

HB1xp67_ASAP7_75t_L g412 ( 
.A(n_295),
.Y(n_412)
);

NOR2xp33_ASAP7_75t_L g413 ( 
.A(n_221),
.B(n_1),
.Y(n_413)
);

INVx1_ASAP7_75t_L g414 ( 
.A(n_231),
.Y(n_414)
);

HB1xp67_ASAP7_75t_L g415 ( 
.A(n_344),
.Y(n_415)
);

INVxp67_ASAP7_75t_L g416 ( 
.A(n_258),
.Y(n_416)
);

INVx1_ASAP7_75t_L g417 ( 
.A(n_231),
.Y(n_417)
);

INVx1_ASAP7_75t_L g418 ( 
.A(n_337),
.Y(n_418)
);

INVx1_ASAP7_75t_L g419 ( 
.A(n_337),
.Y(n_419)
);

INVx3_ASAP7_75t_L g420 ( 
.A(n_210),
.Y(n_420)
);

CKINVDCx20_ASAP7_75t_R g421 ( 
.A(n_281),
.Y(n_421)
);

INVx1_ASAP7_75t_L g422 ( 
.A(n_210),
.Y(n_422)
);

INVx1_ASAP7_75t_L g423 ( 
.A(n_210),
.Y(n_423)
);

INVxp33_ASAP7_75t_SL g424 ( 
.A(n_202),
.Y(n_424)
);

NOR2xp67_ASAP7_75t_L g425 ( 
.A(n_380),
.B(n_1),
.Y(n_425)
);

INVxp33_ASAP7_75t_SL g426 ( 
.A(n_202),
.Y(n_426)
);

INVx2_ASAP7_75t_L g427 ( 
.A(n_210),
.Y(n_427)
);

CKINVDCx5p33_ASAP7_75t_R g428 ( 
.A(n_266),
.Y(n_428)
);

CKINVDCx5p33_ASAP7_75t_R g429 ( 
.A(n_271),
.Y(n_429)
);

CKINVDCx20_ASAP7_75t_R g430 ( 
.A(n_297),
.Y(n_430)
);

CKINVDCx5p33_ASAP7_75t_R g431 ( 
.A(n_274),
.Y(n_431)
);

BUFx6f_ASAP7_75t_SL g432 ( 
.A(n_207),
.Y(n_432)
);

CKINVDCx20_ASAP7_75t_R g433 ( 
.A(n_302),
.Y(n_433)
);

CKINVDCx20_ASAP7_75t_R g434 ( 
.A(n_303),
.Y(n_434)
);

CKINVDCx20_ASAP7_75t_R g435 ( 
.A(n_306),
.Y(n_435)
);

CKINVDCx5p33_ASAP7_75t_R g436 ( 
.A(n_288),
.Y(n_436)
);

INVx1_ASAP7_75t_L g437 ( 
.A(n_201),
.Y(n_437)
);

NAND2xp5_ASAP7_75t_L g438 ( 
.A(n_345),
.B(n_2),
.Y(n_438)
);

INVx1_ASAP7_75t_L g439 ( 
.A(n_206),
.Y(n_439)
);

INVx1_ASAP7_75t_L g440 ( 
.A(n_212),
.Y(n_440)
);

INVxp67_ASAP7_75t_L g441 ( 
.A(n_258),
.Y(n_441)
);

INVx1_ASAP7_75t_L g442 ( 
.A(n_223),
.Y(n_442)
);

CKINVDCx5p33_ASAP7_75t_R g443 ( 
.A(n_290),
.Y(n_443)
);

HB1xp67_ASAP7_75t_L g444 ( 
.A(n_215),
.Y(n_444)
);

INVx1_ASAP7_75t_L g445 ( 
.A(n_254),
.Y(n_445)
);

CKINVDCx5p33_ASAP7_75t_R g446 ( 
.A(n_298),
.Y(n_446)
);

INVx1_ASAP7_75t_L g447 ( 
.A(n_259),
.Y(n_447)
);

INVx1_ASAP7_75t_L g448 ( 
.A(n_268),
.Y(n_448)
);

CKINVDCx16_ASAP7_75t_R g449 ( 
.A(n_326),
.Y(n_449)
);

INVx1_ASAP7_75t_L g450 ( 
.A(n_272),
.Y(n_450)
);

INVx1_ASAP7_75t_L g451 ( 
.A(n_283),
.Y(n_451)
);

INVxp67_ASAP7_75t_SL g452 ( 
.A(n_379),
.Y(n_452)
);

INVx1_ASAP7_75t_L g453 ( 
.A(n_305),
.Y(n_453)
);

INVx1_ASAP7_75t_L g454 ( 
.A(n_286),
.Y(n_454)
);

INVx1_ASAP7_75t_L g455 ( 
.A(n_289),
.Y(n_455)
);

INVx1_ASAP7_75t_L g456 ( 
.A(n_293),
.Y(n_456)
);

CKINVDCx5p33_ASAP7_75t_R g457 ( 
.A(n_301),
.Y(n_457)
);

AND2x2_ASAP7_75t_L g458 ( 
.A(n_401),
.B(n_2),
.Y(n_458)
);

INVxp67_ASAP7_75t_SL g459 ( 
.A(n_217),
.Y(n_459)
);

CKINVDCx20_ASAP7_75t_R g460 ( 
.A(n_309),
.Y(n_460)
);

CKINVDCx5p33_ASAP7_75t_R g461 ( 
.A(n_308),
.Y(n_461)
);

INVx1_ASAP7_75t_L g462 ( 
.A(n_313),
.Y(n_462)
);

INVx1_ASAP7_75t_L g463 ( 
.A(n_317),
.Y(n_463)
);

CKINVDCx5p33_ASAP7_75t_R g464 ( 
.A(n_311),
.Y(n_464)
);

BUFx3_ASAP7_75t_L g465 ( 
.A(n_260),
.Y(n_465)
);

INVx1_ASAP7_75t_L g466 ( 
.A(n_305),
.Y(n_466)
);

INVx1_ASAP7_75t_L g467 ( 
.A(n_318),
.Y(n_467)
);

CKINVDCx5p33_ASAP7_75t_R g468 ( 
.A(n_320),
.Y(n_468)
);

INVx1_ASAP7_75t_L g469 ( 
.A(n_322),
.Y(n_469)
);

INVx1_ASAP7_75t_L g470 ( 
.A(n_342),
.Y(n_470)
);

INVx1_ASAP7_75t_L g471 ( 
.A(n_348),
.Y(n_471)
);

INVx1_ASAP7_75t_L g472 ( 
.A(n_378),
.Y(n_472)
);

CKINVDCx5p33_ASAP7_75t_R g473 ( 
.A(n_324),
.Y(n_473)
);

CKINVDCx20_ASAP7_75t_R g474 ( 
.A(n_321),
.Y(n_474)
);

CKINVDCx5p33_ASAP7_75t_R g475 ( 
.A(n_331),
.Y(n_475)
);

INVx1_ASAP7_75t_L g476 ( 
.A(n_388),
.Y(n_476)
);

XNOR2xp5_ASAP7_75t_L g477 ( 
.A(n_208),
.B(n_3),
.Y(n_477)
);

NOR2xp33_ASAP7_75t_L g478 ( 
.A(n_345),
.B(n_3),
.Y(n_478)
);

INVx1_ASAP7_75t_L g479 ( 
.A(n_389),
.Y(n_479)
);

OR2x2_ASAP7_75t_L g480 ( 
.A(n_390),
.B(n_4),
.Y(n_480)
);

CKINVDCx5p33_ASAP7_75t_R g481 ( 
.A(n_332),
.Y(n_481)
);

INVx1_ASAP7_75t_L g482 ( 
.A(n_396),
.Y(n_482)
);

INVxp67_ASAP7_75t_SL g483 ( 
.A(n_260),
.Y(n_483)
);

INVx1_ASAP7_75t_L g484 ( 
.A(n_273),
.Y(n_484)
);

INVx1_ASAP7_75t_L g485 ( 
.A(n_273),
.Y(n_485)
);

INVx1_ASAP7_75t_L g486 ( 
.A(n_209),
.Y(n_486)
);

CKINVDCx5p33_ASAP7_75t_R g487 ( 
.A(n_335),
.Y(n_487)
);

INVx1_ASAP7_75t_L g488 ( 
.A(n_220),
.Y(n_488)
);

INVxp67_ASAP7_75t_L g489 ( 
.A(n_258),
.Y(n_489)
);

CKINVDCx20_ASAP7_75t_R g490 ( 
.A(n_323),
.Y(n_490)
);

CKINVDCx20_ASAP7_75t_R g491 ( 
.A(n_333),
.Y(n_491)
);

INVx1_ASAP7_75t_L g492 ( 
.A(n_222),
.Y(n_492)
);

CKINVDCx20_ASAP7_75t_R g493 ( 
.A(n_243),
.Y(n_493)
);

NOR2xp33_ASAP7_75t_L g494 ( 
.A(n_380),
.B(n_6),
.Y(n_494)
);

INVx1_ASAP7_75t_L g495 ( 
.A(n_224),
.Y(n_495)
);

INVx1_ASAP7_75t_L g496 ( 
.A(n_229),
.Y(n_496)
);

INVx1_ASAP7_75t_L g497 ( 
.A(n_230),
.Y(n_497)
);

INVx1_ASAP7_75t_L g498 ( 
.A(n_232),
.Y(n_498)
);

CKINVDCx5p33_ASAP7_75t_R g499 ( 
.A(n_338),
.Y(n_499)
);

INVx1_ASAP7_75t_L g500 ( 
.A(n_382),
.Y(n_500)
);

INVxp67_ASAP7_75t_L g501 ( 
.A(n_334),
.Y(n_501)
);

CKINVDCx16_ASAP7_75t_R g502 ( 
.A(n_334),
.Y(n_502)
);

CKINVDCx20_ASAP7_75t_R g503 ( 
.A(n_245),
.Y(n_503)
);

INVx1_ASAP7_75t_L g504 ( 
.A(n_233),
.Y(n_504)
);

INVx3_ASAP7_75t_L g505 ( 
.A(n_420),
.Y(n_505)
);

AND2x2_ASAP7_75t_L g506 ( 
.A(n_484),
.B(n_380),
.Y(n_506)
);

INVx3_ASAP7_75t_L g507 ( 
.A(n_420),
.Y(n_507)
);

INVx1_ASAP7_75t_L g508 ( 
.A(n_403),
.Y(n_508)
);

INVx1_ASAP7_75t_L g509 ( 
.A(n_403),
.Y(n_509)
);

BUFx6f_ASAP7_75t_L g510 ( 
.A(n_427),
.Y(n_510)
);

INVx2_ASAP7_75t_L g511 ( 
.A(n_427),
.Y(n_511)
);

INVx1_ASAP7_75t_L g512 ( 
.A(n_422),
.Y(n_512)
);

CKINVDCx20_ASAP7_75t_R g513 ( 
.A(n_406),
.Y(n_513)
);

INVx1_ASAP7_75t_L g514 ( 
.A(n_422),
.Y(n_514)
);

OA21x2_ASAP7_75t_L g515 ( 
.A1(n_423),
.A2(n_395),
.B(n_382),
.Y(n_515)
);

AND2x2_ASAP7_75t_L g516 ( 
.A(n_485),
.B(n_386),
.Y(n_516)
);

INVx1_ASAP7_75t_L g517 ( 
.A(n_423),
.Y(n_517)
);

CKINVDCx5p33_ASAP7_75t_R g518 ( 
.A(n_493),
.Y(n_518)
);

INVx1_ASAP7_75t_L g519 ( 
.A(n_420),
.Y(n_519)
);

INVx1_ASAP7_75t_L g520 ( 
.A(n_453),
.Y(n_520)
);

INVx1_ASAP7_75t_L g521 ( 
.A(n_453),
.Y(n_521)
);

NOR2xp33_ASAP7_75t_L g522 ( 
.A(n_452),
.B(n_249),
.Y(n_522)
);

BUFx6f_ASAP7_75t_L g523 ( 
.A(n_466),
.Y(n_523)
);

HB1xp67_ASAP7_75t_L g524 ( 
.A(n_444),
.Y(n_524)
);

INVx2_ASAP7_75t_L g525 ( 
.A(n_466),
.Y(n_525)
);

INVx1_ASAP7_75t_L g526 ( 
.A(n_500),
.Y(n_526)
);

INVxp67_ASAP7_75t_L g527 ( 
.A(n_415),
.Y(n_527)
);

INVx1_ASAP7_75t_L g528 ( 
.A(n_500),
.Y(n_528)
);

AND2x6_ASAP7_75t_L g529 ( 
.A(n_458),
.B(n_386),
.Y(n_529)
);

INVx2_ASAP7_75t_L g530 ( 
.A(n_486),
.Y(n_530)
);

INVx1_ASAP7_75t_L g531 ( 
.A(n_437),
.Y(n_531)
);

INVx1_ASAP7_75t_L g532 ( 
.A(n_439),
.Y(n_532)
);

NAND2xp5_ASAP7_75t_L g533 ( 
.A(n_494),
.B(n_203),
.Y(n_533)
);

INVx4_ASAP7_75t_L g534 ( 
.A(n_410),
.Y(n_534)
);

INVx1_ASAP7_75t_L g535 ( 
.A(n_440),
.Y(n_535)
);

BUFx6f_ASAP7_75t_L g536 ( 
.A(n_488),
.Y(n_536)
);

INVx1_ASAP7_75t_L g537 ( 
.A(n_442),
.Y(n_537)
);

CKINVDCx5p33_ASAP7_75t_R g538 ( 
.A(n_503),
.Y(n_538)
);

BUFx2_ASAP7_75t_L g539 ( 
.A(n_402),
.Y(n_539)
);

HB1xp67_ASAP7_75t_L g540 ( 
.A(n_410),
.Y(n_540)
);

CKINVDCx5p33_ASAP7_75t_R g541 ( 
.A(n_404),
.Y(n_541)
);

NAND2xp5_ASAP7_75t_L g542 ( 
.A(n_492),
.B(n_203),
.Y(n_542)
);

INVx2_ASAP7_75t_L g543 ( 
.A(n_495),
.Y(n_543)
);

INVx1_ASAP7_75t_L g544 ( 
.A(n_445),
.Y(n_544)
);

CKINVDCx5p33_ASAP7_75t_R g545 ( 
.A(n_404),
.Y(n_545)
);

CKINVDCx5p33_ASAP7_75t_R g546 ( 
.A(n_405),
.Y(n_546)
);

INVx2_ASAP7_75t_L g547 ( 
.A(n_504),
.Y(n_547)
);

CKINVDCx20_ASAP7_75t_R g548 ( 
.A(n_408),
.Y(n_548)
);

INVx1_ASAP7_75t_L g549 ( 
.A(n_447),
.Y(n_549)
);

CKINVDCx20_ASAP7_75t_R g550 ( 
.A(n_409),
.Y(n_550)
);

INVx1_ASAP7_75t_L g551 ( 
.A(n_448),
.Y(n_551)
);

INVx1_ASAP7_75t_L g552 ( 
.A(n_450),
.Y(n_552)
);

INVx1_ASAP7_75t_L g553 ( 
.A(n_451),
.Y(n_553)
);

CKINVDCx5p33_ASAP7_75t_R g554 ( 
.A(n_405),
.Y(n_554)
);

INVx2_ASAP7_75t_L g555 ( 
.A(n_496),
.Y(n_555)
);

CKINVDCx5p33_ASAP7_75t_R g556 ( 
.A(n_407),
.Y(n_556)
);

CKINVDCx20_ASAP7_75t_R g557 ( 
.A(n_421),
.Y(n_557)
);

NAND2xp5_ASAP7_75t_L g558 ( 
.A(n_497),
.B(n_204),
.Y(n_558)
);

INVx1_ASAP7_75t_L g559 ( 
.A(n_454),
.Y(n_559)
);

INVx2_ASAP7_75t_L g560 ( 
.A(n_498),
.Y(n_560)
);

INVx2_ASAP7_75t_L g561 ( 
.A(n_455),
.Y(n_561)
);

CKINVDCx5p33_ASAP7_75t_R g562 ( 
.A(n_407),
.Y(n_562)
);

INVx3_ASAP7_75t_L g563 ( 
.A(n_456),
.Y(n_563)
);

BUFx3_ASAP7_75t_L g564 ( 
.A(n_465),
.Y(n_564)
);

INVx1_ASAP7_75t_L g565 ( 
.A(n_462),
.Y(n_565)
);

INVx3_ASAP7_75t_L g566 ( 
.A(n_463),
.Y(n_566)
);

CKINVDCx5p33_ASAP7_75t_R g567 ( 
.A(n_411),
.Y(n_567)
);

NOR2xp33_ASAP7_75t_L g568 ( 
.A(n_438),
.B(n_386),
.Y(n_568)
);

CKINVDCx20_ASAP7_75t_R g569 ( 
.A(n_430),
.Y(n_569)
);

INVx3_ASAP7_75t_L g570 ( 
.A(n_467),
.Y(n_570)
);

BUFx10_ASAP7_75t_L g571 ( 
.A(n_432),
.Y(n_571)
);

INVx1_ASAP7_75t_L g572 ( 
.A(n_469),
.Y(n_572)
);

INVx1_ASAP7_75t_L g573 ( 
.A(n_470),
.Y(n_573)
);

INVx2_ASAP7_75t_L g574 ( 
.A(n_471),
.Y(n_574)
);

INVx1_ASAP7_75t_L g575 ( 
.A(n_472),
.Y(n_575)
);

INVx1_ASAP7_75t_L g576 ( 
.A(n_476),
.Y(n_576)
);

AND2x4_ASAP7_75t_L g577 ( 
.A(n_425),
.B(n_278),
.Y(n_577)
);

INVx2_ASAP7_75t_L g578 ( 
.A(n_479),
.Y(n_578)
);

CKINVDCx20_ASAP7_75t_R g579 ( 
.A(n_433),
.Y(n_579)
);

CKINVDCx5p33_ASAP7_75t_R g580 ( 
.A(n_411),
.Y(n_580)
);

CKINVDCx5p33_ASAP7_75t_R g581 ( 
.A(n_428),
.Y(n_581)
);

BUFx6f_ASAP7_75t_L g582 ( 
.A(n_482),
.Y(n_582)
);

INVx1_ASAP7_75t_SL g583 ( 
.A(n_428),
.Y(n_583)
);

AND2x2_ASAP7_75t_L g584 ( 
.A(n_459),
.B(n_278),
.Y(n_584)
);

INVx2_ASAP7_75t_L g585 ( 
.A(n_465),
.Y(n_585)
);

INVx2_ASAP7_75t_L g586 ( 
.A(n_414),
.Y(n_586)
);

BUFx4f_ASAP7_75t_L g587 ( 
.A(n_515),
.Y(n_587)
);

INVx1_ASAP7_75t_L g588 ( 
.A(n_585),
.Y(n_588)
);

NAND2xp5_ASAP7_75t_SL g589 ( 
.A(n_568),
.B(n_294),
.Y(n_589)
);

INVx2_ASAP7_75t_L g590 ( 
.A(n_511),
.Y(n_590)
);

INVx2_ASAP7_75t_L g591 ( 
.A(n_511),
.Y(n_591)
);

AOI22xp33_ASAP7_75t_L g592 ( 
.A1(n_568),
.A2(n_458),
.B1(n_478),
.B2(n_413),
.Y(n_592)
);

NOR2xp33_ASAP7_75t_L g593 ( 
.A(n_522),
.B(n_449),
.Y(n_593)
);

INVxp67_ASAP7_75t_L g594 ( 
.A(n_540),
.Y(n_594)
);

NOR2xp33_ASAP7_75t_L g595 ( 
.A(n_534),
.B(n_424),
.Y(n_595)
);

INVx1_ASAP7_75t_L g596 ( 
.A(n_585),
.Y(n_596)
);

BUFx3_ASAP7_75t_L g597 ( 
.A(n_564),
.Y(n_597)
);

INVx1_ASAP7_75t_L g598 ( 
.A(n_531),
.Y(n_598)
);

INVx1_ASAP7_75t_L g599 ( 
.A(n_531),
.Y(n_599)
);

NAND2xp33_ASAP7_75t_L g600 ( 
.A(n_529),
.B(n_228),
.Y(n_600)
);

INVx2_ASAP7_75t_L g601 ( 
.A(n_511),
.Y(n_601)
);

NAND2xp5_ASAP7_75t_L g602 ( 
.A(n_533),
.B(n_483),
.Y(n_602)
);

INVx2_ASAP7_75t_L g603 ( 
.A(n_508),
.Y(n_603)
);

INVx2_ASAP7_75t_L g604 ( 
.A(n_508),
.Y(n_604)
);

INVx1_ASAP7_75t_L g605 ( 
.A(n_532),
.Y(n_605)
);

BUFx10_ASAP7_75t_L g606 ( 
.A(n_541),
.Y(n_606)
);

INVx1_ASAP7_75t_L g607 ( 
.A(n_532),
.Y(n_607)
);

OAI22xp33_ASAP7_75t_SL g608 ( 
.A1(n_533),
.A2(n_480),
.B1(n_558),
.B2(n_542),
.Y(n_608)
);

NOR2xp33_ASAP7_75t_L g609 ( 
.A(n_534),
.B(n_424),
.Y(n_609)
);

INVx3_ASAP7_75t_L g610 ( 
.A(n_510),
.Y(n_610)
);

NOR3xp33_ASAP7_75t_L g611 ( 
.A(n_527),
.B(n_502),
.C(n_441),
.Y(n_611)
);

NAND2xp5_ASAP7_75t_L g612 ( 
.A(n_584),
.B(n_577),
.Y(n_612)
);

INVx1_ASAP7_75t_L g613 ( 
.A(n_535),
.Y(n_613)
);

BUFx6f_ASAP7_75t_L g614 ( 
.A(n_515),
.Y(n_614)
);

NAND2xp5_ASAP7_75t_L g615 ( 
.A(n_584),
.B(n_429),
.Y(n_615)
);

NOR2xp33_ASAP7_75t_L g616 ( 
.A(n_534),
.B(n_426),
.Y(n_616)
);

OR2x2_ASAP7_75t_L g617 ( 
.A(n_527),
.B(n_429),
.Y(n_617)
);

INVx1_ASAP7_75t_L g618 ( 
.A(n_535),
.Y(n_618)
);

NAND2xp5_ASAP7_75t_L g619 ( 
.A(n_584),
.B(n_431),
.Y(n_619)
);

NAND2xp5_ASAP7_75t_L g620 ( 
.A(n_577),
.B(n_431),
.Y(n_620)
);

NAND2xp33_ASAP7_75t_SL g621 ( 
.A(n_540),
.B(n_393),
.Y(n_621)
);

NOR2xp33_ASAP7_75t_L g622 ( 
.A(n_534),
.B(n_426),
.Y(n_622)
);

INVx1_ASAP7_75t_L g623 ( 
.A(n_537),
.Y(n_623)
);

NAND2xp5_ASAP7_75t_SL g624 ( 
.A(n_577),
.B(n_294),
.Y(n_624)
);

INVx1_ASAP7_75t_L g625 ( 
.A(n_537),
.Y(n_625)
);

AND2x2_ASAP7_75t_L g626 ( 
.A(n_506),
.B(n_417),
.Y(n_626)
);

NAND2xp5_ASAP7_75t_L g627 ( 
.A(n_577),
.B(n_436),
.Y(n_627)
);

OR2x6_ASAP7_75t_L g628 ( 
.A(n_564),
.B(n_480),
.Y(n_628)
);

OR2x6_ASAP7_75t_L g629 ( 
.A(n_564),
.B(n_393),
.Y(n_629)
);

INVx2_ASAP7_75t_L g630 ( 
.A(n_509),
.Y(n_630)
);

INVx2_ASAP7_75t_L g631 ( 
.A(n_509),
.Y(n_631)
);

NAND2xp5_ASAP7_75t_SL g632 ( 
.A(n_583),
.B(n_299),
.Y(n_632)
);

NAND3xp33_ASAP7_75t_SL g633 ( 
.A(n_583),
.B(n_402),
.C(n_436),
.Y(n_633)
);

INVx2_ASAP7_75t_L g634 ( 
.A(n_512),
.Y(n_634)
);

BUFx3_ASAP7_75t_L g635 ( 
.A(n_515),
.Y(n_635)
);

INVx4_ASAP7_75t_L g636 ( 
.A(n_529),
.Y(n_636)
);

BUFx10_ASAP7_75t_L g637 ( 
.A(n_545),
.Y(n_637)
);

INVx1_ASAP7_75t_SL g638 ( 
.A(n_539),
.Y(n_638)
);

NAND3xp33_ASAP7_75t_L g639 ( 
.A(n_542),
.B(n_446),
.C(n_443),
.Y(n_639)
);

INVx2_ASAP7_75t_SL g640 ( 
.A(n_524),
.Y(n_640)
);

INVxp67_ASAP7_75t_L g641 ( 
.A(n_524),
.Y(n_641)
);

NAND2xp5_ASAP7_75t_L g642 ( 
.A(n_529),
.B(n_443),
.Y(n_642)
);

BUFx2_ASAP7_75t_L g643 ( 
.A(n_539),
.Y(n_643)
);

INVx2_ASAP7_75t_L g644 ( 
.A(n_512),
.Y(n_644)
);

INVx4_ASAP7_75t_L g645 ( 
.A(n_529),
.Y(n_645)
);

OR2x2_ASAP7_75t_L g646 ( 
.A(n_558),
.B(n_446),
.Y(n_646)
);

INVx1_ASAP7_75t_L g647 ( 
.A(n_544),
.Y(n_647)
);

INVx1_ASAP7_75t_SL g648 ( 
.A(n_513),
.Y(n_648)
);

INVx2_ASAP7_75t_L g649 ( 
.A(n_514),
.Y(n_649)
);

AND2x4_ASAP7_75t_L g650 ( 
.A(n_506),
.B(n_418),
.Y(n_650)
);

INVx2_ASAP7_75t_L g651 ( 
.A(n_514),
.Y(n_651)
);

INVx2_ASAP7_75t_L g652 ( 
.A(n_517),
.Y(n_652)
);

INVx2_ASAP7_75t_L g653 ( 
.A(n_517),
.Y(n_653)
);

INVx3_ASAP7_75t_L g654 ( 
.A(n_510),
.Y(n_654)
);

AND2x4_ASAP7_75t_L g655 ( 
.A(n_506),
.B(n_419),
.Y(n_655)
);

NOR2xp33_ASAP7_75t_SL g656 ( 
.A(n_546),
.B(n_434),
.Y(n_656)
);

NAND2xp5_ASAP7_75t_SL g657 ( 
.A(n_582),
.B(n_299),
.Y(n_657)
);

BUFx3_ASAP7_75t_L g658 ( 
.A(n_515),
.Y(n_658)
);

INVx3_ASAP7_75t_L g659 ( 
.A(n_510),
.Y(n_659)
);

BUFx3_ASAP7_75t_L g660 ( 
.A(n_515),
.Y(n_660)
);

INVx5_ASAP7_75t_L g661 ( 
.A(n_529),
.Y(n_661)
);

INVx3_ASAP7_75t_L g662 ( 
.A(n_510),
.Y(n_662)
);

INVx2_ASAP7_75t_L g663 ( 
.A(n_523),
.Y(n_663)
);

AND2x6_ASAP7_75t_L g664 ( 
.A(n_516),
.B(n_371),
.Y(n_664)
);

INVx1_ASAP7_75t_L g665 ( 
.A(n_544),
.Y(n_665)
);

NAND2xp33_ASAP7_75t_L g666 ( 
.A(n_529),
.B(n_228),
.Y(n_666)
);

BUFx6f_ASAP7_75t_L g667 ( 
.A(n_536),
.Y(n_667)
);

INVx1_ASAP7_75t_L g668 ( 
.A(n_549),
.Y(n_668)
);

NAND2xp5_ASAP7_75t_SL g669 ( 
.A(n_582),
.B(n_371),
.Y(n_669)
);

INVx1_ASAP7_75t_L g670 ( 
.A(n_549),
.Y(n_670)
);

NOR2xp33_ASAP7_75t_L g671 ( 
.A(n_554),
.B(n_457),
.Y(n_671)
);

BUFx6f_ASAP7_75t_L g672 ( 
.A(n_536),
.Y(n_672)
);

BUFx3_ASAP7_75t_L g673 ( 
.A(n_505),
.Y(n_673)
);

INVx2_ASAP7_75t_L g674 ( 
.A(n_523),
.Y(n_674)
);

INVx1_ASAP7_75t_L g675 ( 
.A(n_551),
.Y(n_675)
);

AND2x2_ASAP7_75t_L g676 ( 
.A(n_571),
.B(n_457),
.Y(n_676)
);

CKINVDCx5p33_ASAP7_75t_R g677 ( 
.A(n_518),
.Y(n_677)
);

INVx3_ASAP7_75t_L g678 ( 
.A(n_510),
.Y(n_678)
);

OAI21xp33_ASAP7_75t_L g679 ( 
.A1(n_552),
.A2(n_464),
.B(n_461),
.Y(n_679)
);

NOR2xp33_ASAP7_75t_L g680 ( 
.A(n_556),
.B(n_461),
.Y(n_680)
);

AND2x2_ASAP7_75t_L g681 ( 
.A(n_516),
.B(n_464),
.Y(n_681)
);

NAND2xp5_ASAP7_75t_L g682 ( 
.A(n_529),
.B(n_505),
.Y(n_682)
);

INVx2_ASAP7_75t_L g683 ( 
.A(n_523),
.Y(n_683)
);

OR2x2_ASAP7_75t_L g684 ( 
.A(n_516),
.B(n_468),
.Y(n_684)
);

INVx3_ASAP7_75t_L g685 ( 
.A(n_510),
.Y(n_685)
);

INVx2_ASAP7_75t_L g686 ( 
.A(n_523),
.Y(n_686)
);

BUFx6f_ASAP7_75t_L g687 ( 
.A(n_536),
.Y(n_687)
);

OAI22xp5_ASAP7_75t_L g688 ( 
.A1(n_562),
.A2(n_475),
.B1(n_499),
.B2(n_468),
.Y(n_688)
);

INVx2_ASAP7_75t_SL g689 ( 
.A(n_586),
.Y(n_689)
);

NAND2xp33_ASAP7_75t_L g690 ( 
.A(n_529),
.B(n_228),
.Y(n_690)
);

AO22x2_ASAP7_75t_L g691 ( 
.A1(n_586),
.A2(n_401),
.B1(n_395),
.B2(n_238),
.Y(n_691)
);

BUFx2_ASAP7_75t_L g692 ( 
.A(n_567),
.Y(n_692)
);

INVx2_ASAP7_75t_L g693 ( 
.A(n_523),
.Y(n_693)
);

NOR2xp33_ASAP7_75t_L g694 ( 
.A(n_580),
.B(n_473),
.Y(n_694)
);

INVx2_ASAP7_75t_L g695 ( 
.A(n_523),
.Y(n_695)
);

INVx2_ASAP7_75t_L g696 ( 
.A(n_523),
.Y(n_696)
);

INVx2_ASAP7_75t_L g697 ( 
.A(n_519),
.Y(n_697)
);

INVx6_ASAP7_75t_L g698 ( 
.A(n_571),
.Y(n_698)
);

INVx1_ASAP7_75t_L g699 ( 
.A(n_552),
.Y(n_699)
);

BUFx3_ASAP7_75t_L g700 ( 
.A(n_505),
.Y(n_700)
);

CKINVDCx20_ASAP7_75t_R g701 ( 
.A(n_548),
.Y(n_701)
);

AOI22xp33_ASAP7_75t_L g702 ( 
.A1(n_563),
.A2(n_292),
.B1(n_257),
.B2(n_228),
.Y(n_702)
);

INVx1_ASAP7_75t_L g703 ( 
.A(n_553),
.Y(n_703)
);

NOR2x1p5_ASAP7_75t_L g704 ( 
.A(n_581),
.B(n_473),
.Y(n_704)
);

INVx1_ASAP7_75t_SL g705 ( 
.A(n_550),
.Y(n_705)
);

AND2x6_ASAP7_75t_L g706 ( 
.A(n_563),
.B(n_228),
.Y(n_706)
);

CKINVDCx20_ASAP7_75t_R g707 ( 
.A(n_557),
.Y(n_707)
);

NAND2xp5_ASAP7_75t_SL g708 ( 
.A(n_582),
.B(n_257),
.Y(n_708)
);

AND2x2_ASAP7_75t_L g709 ( 
.A(n_586),
.B(n_475),
.Y(n_709)
);

BUFx6f_ASAP7_75t_L g710 ( 
.A(n_536),
.Y(n_710)
);

AND2x4_ASAP7_75t_L g711 ( 
.A(n_559),
.B(n_240),
.Y(n_711)
);

OR2x2_ASAP7_75t_L g712 ( 
.A(n_563),
.B(n_481),
.Y(n_712)
);

NAND2xp5_ASAP7_75t_SL g713 ( 
.A(n_582),
.B(n_257),
.Y(n_713)
);

NOR2xp33_ASAP7_75t_L g714 ( 
.A(n_563),
.B(n_481),
.Y(n_714)
);

INVxp67_ASAP7_75t_SL g715 ( 
.A(n_507),
.Y(n_715)
);

NOR2xp33_ASAP7_75t_L g716 ( 
.A(n_566),
.B(n_487),
.Y(n_716)
);

NAND2xp5_ASAP7_75t_SL g717 ( 
.A(n_582),
.B(n_257),
.Y(n_717)
);

INVxp67_ASAP7_75t_SL g718 ( 
.A(n_507),
.Y(n_718)
);

CKINVDCx6p67_ASAP7_75t_R g719 ( 
.A(n_571),
.Y(n_719)
);

NAND3xp33_ASAP7_75t_L g720 ( 
.A(n_565),
.B(n_499),
.C(n_487),
.Y(n_720)
);

INVx2_ASAP7_75t_L g721 ( 
.A(n_519),
.Y(n_721)
);

INVx2_ASAP7_75t_L g722 ( 
.A(n_507),
.Y(n_722)
);

INVx1_ASAP7_75t_L g723 ( 
.A(n_565),
.Y(n_723)
);

CKINVDCx20_ASAP7_75t_R g724 ( 
.A(n_569),
.Y(n_724)
);

NAND2xp5_ASAP7_75t_L g725 ( 
.A(n_507),
.B(n_246),
.Y(n_725)
);

NOR2xp33_ASAP7_75t_L g726 ( 
.A(n_566),
.B(n_432),
.Y(n_726)
);

INVx2_ASAP7_75t_L g727 ( 
.A(n_510),
.Y(n_727)
);

NAND2xp5_ASAP7_75t_SL g728 ( 
.A(n_582),
.B(n_257),
.Y(n_728)
);

INVx2_ASAP7_75t_L g729 ( 
.A(n_525),
.Y(n_729)
);

AND2x2_ASAP7_75t_L g730 ( 
.A(n_571),
.B(n_501),
.Y(n_730)
);

INVx3_ASAP7_75t_L g731 ( 
.A(n_536),
.Y(n_731)
);

BUFx10_ASAP7_75t_L g732 ( 
.A(n_538),
.Y(n_732)
);

OR2x2_ASAP7_75t_L g733 ( 
.A(n_566),
.B(n_416),
.Y(n_733)
);

CKINVDCx20_ASAP7_75t_R g734 ( 
.A(n_579),
.Y(n_734)
);

NAND2xp5_ASAP7_75t_L g735 ( 
.A(n_602),
.B(n_536),
.Y(n_735)
);

INVx1_ASAP7_75t_L g736 ( 
.A(n_598),
.Y(n_736)
);

NAND2xp5_ASAP7_75t_L g737 ( 
.A(n_612),
.B(n_536),
.Y(n_737)
);

INVx1_ASAP7_75t_L g738 ( 
.A(n_599),
.Y(n_738)
);

NAND2xp5_ASAP7_75t_L g739 ( 
.A(n_714),
.B(n_566),
.Y(n_739)
);

INVx1_ASAP7_75t_L g740 ( 
.A(n_605),
.Y(n_740)
);

NAND2xp5_ASAP7_75t_L g741 ( 
.A(n_716),
.B(n_570),
.Y(n_741)
);

AOI22xp33_ASAP7_75t_L g742 ( 
.A1(n_589),
.A2(n_570),
.B1(n_582),
.B2(n_304),
.Y(n_742)
);

AOI22xp5_ASAP7_75t_L g743 ( 
.A1(n_608),
.A2(n_435),
.B1(n_460),
.B2(n_474),
.Y(n_743)
);

INVxp67_ASAP7_75t_L g744 ( 
.A(n_617),
.Y(n_744)
);

NAND2xp5_ASAP7_75t_SL g745 ( 
.A(n_661),
.B(n_292),
.Y(n_745)
);

OAI22xp33_ASAP7_75t_L g746 ( 
.A1(n_615),
.A2(n_490),
.B1(n_491),
.B2(n_276),
.Y(n_746)
);

INVx2_ASAP7_75t_L g747 ( 
.A(n_603),
.Y(n_747)
);

O2A1O1Ixp33_ASAP7_75t_L g748 ( 
.A1(n_589),
.A2(n_573),
.B(n_576),
.C(n_575),
.Y(n_748)
);

NAND2xp5_ASAP7_75t_SL g749 ( 
.A(n_661),
.B(n_292),
.Y(n_749)
);

OAI22x1_ASAP7_75t_L g750 ( 
.A1(n_640),
.A2(n_477),
.B1(n_489),
.B2(n_242),
.Y(n_750)
);

NAND2xp5_ASAP7_75t_SL g751 ( 
.A(n_661),
.B(n_292),
.Y(n_751)
);

NAND2xp5_ASAP7_75t_L g752 ( 
.A(n_689),
.B(n_570),
.Y(n_752)
);

NAND2xp5_ASAP7_75t_L g753 ( 
.A(n_689),
.B(n_570),
.Y(n_753)
);

NAND2xp5_ASAP7_75t_SL g754 ( 
.A(n_661),
.B(n_292),
.Y(n_754)
);

INVx2_ASAP7_75t_SL g755 ( 
.A(n_684),
.Y(n_755)
);

A2O1A1Ixp33_ASAP7_75t_L g756 ( 
.A1(n_592),
.A2(n_573),
.B(n_576),
.C(n_575),
.Y(n_756)
);

NAND2xp5_ASAP7_75t_L g757 ( 
.A(n_614),
.B(n_530),
.Y(n_757)
);

INVx1_ASAP7_75t_L g758 ( 
.A(n_607),
.Y(n_758)
);

NAND2xp5_ASAP7_75t_L g759 ( 
.A(n_614),
.B(n_530),
.Y(n_759)
);

NAND2xp5_ASAP7_75t_SL g760 ( 
.A(n_661),
.B(n_241),
.Y(n_760)
);

NAND2xp5_ASAP7_75t_L g761 ( 
.A(n_614),
.B(n_530),
.Y(n_761)
);

NAND2xp5_ASAP7_75t_L g762 ( 
.A(n_614),
.B(n_543),
.Y(n_762)
);

INVx2_ASAP7_75t_L g763 ( 
.A(n_603),
.Y(n_763)
);

INVx2_ASAP7_75t_L g764 ( 
.A(n_604),
.Y(n_764)
);

INVxp67_ASAP7_75t_L g765 ( 
.A(n_640),
.Y(n_765)
);

NAND2xp5_ASAP7_75t_L g766 ( 
.A(n_715),
.B(n_543),
.Y(n_766)
);

BUFx6f_ASAP7_75t_L g767 ( 
.A(n_635),
.Y(n_767)
);

CKINVDCx5p33_ASAP7_75t_R g768 ( 
.A(n_677),
.Y(n_768)
);

NAND2xp5_ASAP7_75t_L g769 ( 
.A(n_718),
.B(n_543),
.Y(n_769)
);

OAI22xp5_ASAP7_75t_L g770 ( 
.A1(n_642),
.A2(n_280),
.B1(n_269),
.B2(n_265),
.Y(n_770)
);

INVx2_ASAP7_75t_L g771 ( 
.A(n_604),
.Y(n_771)
);

INVx1_ASAP7_75t_L g772 ( 
.A(n_613),
.Y(n_772)
);

AOI22xp33_ASAP7_75t_L g773 ( 
.A1(n_664),
.A2(n_307),
.B1(n_310),
.B2(n_315),
.Y(n_773)
);

INVx2_ASAP7_75t_L g774 ( 
.A(n_630),
.Y(n_774)
);

AND2x2_ASAP7_75t_L g775 ( 
.A(n_681),
.B(n_412),
.Y(n_775)
);

O2A1O1Ixp33_ASAP7_75t_L g776 ( 
.A1(n_619),
.A2(n_632),
.B(n_624),
.C(n_627),
.Y(n_776)
);

INVxp67_ASAP7_75t_L g777 ( 
.A(n_643),
.Y(n_777)
);

AOI221xp5_ASAP7_75t_L g778 ( 
.A1(n_632),
.A2(n_477),
.B1(n_285),
.B2(n_365),
.C(n_346),
.Y(n_778)
);

INVxp67_ASAP7_75t_L g779 ( 
.A(n_646),
.Y(n_779)
);

NOR2xp33_ASAP7_75t_L g780 ( 
.A(n_593),
.B(n_432),
.Y(n_780)
);

NAND2xp5_ASAP7_75t_SL g781 ( 
.A(n_636),
.B(n_244),
.Y(n_781)
);

NAND2xp5_ASAP7_75t_SL g782 ( 
.A(n_636),
.B(n_248),
.Y(n_782)
);

NOR2xp33_ASAP7_75t_L g783 ( 
.A(n_594),
.B(n_712),
.Y(n_783)
);

INVx1_ASAP7_75t_L g784 ( 
.A(n_618),
.Y(n_784)
);

NAND2xp5_ASAP7_75t_L g785 ( 
.A(n_709),
.B(n_547),
.Y(n_785)
);

AOI22xp5_ASAP7_75t_L g786 ( 
.A1(n_681),
.A2(n_284),
.B1(n_247),
.B2(n_261),
.Y(n_786)
);

AND2x2_ASAP7_75t_L g787 ( 
.A(n_709),
.B(n_572),
.Y(n_787)
);

NAND2xp5_ASAP7_75t_L g788 ( 
.A(n_623),
.B(n_547),
.Y(n_788)
);

INVx2_ASAP7_75t_L g789 ( 
.A(n_630),
.Y(n_789)
);

BUFx2_ASAP7_75t_L g790 ( 
.A(n_701),
.Y(n_790)
);

INVx2_ASAP7_75t_L g791 ( 
.A(n_631),
.Y(n_791)
);

NAND2xp5_ASAP7_75t_SL g792 ( 
.A(n_636),
.B(n_250),
.Y(n_792)
);

NOR2xp67_ASAP7_75t_L g793 ( 
.A(n_720),
.B(n_572),
.Y(n_793)
);

NOR2xp33_ASAP7_75t_L g794 ( 
.A(n_620),
.B(n_204),
.Y(n_794)
);

INVx2_ASAP7_75t_SL g795 ( 
.A(n_733),
.Y(n_795)
);

BUFx3_ASAP7_75t_L g796 ( 
.A(n_597),
.Y(n_796)
);

BUFx3_ASAP7_75t_L g797 ( 
.A(n_597),
.Y(n_797)
);

NAND2xp5_ASAP7_75t_L g798 ( 
.A(n_625),
.B(n_547),
.Y(n_798)
);

INVxp67_ASAP7_75t_L g799 ( 
.A(n_671),
.Y(n_799)
);

INVx1_ASAP7_75t_SL g800 ( 
.A(n_638),
.Y(n_800)
);

NOR2xp33_ASAP7_75t_L g801 ( 
.A(n_679),
.B(n_205),
.Y(n_801)
);

AOI22xp5_ASAP7_75t_L g802 ( 
.A1(n_595),
.A2(n_287),
.B1(n_267),
.B2(n_270),
.Y(n_802)
);

AOI21xp5_ASAP7_75t_L g803 ( 
.A1(n_587),
.A2(n_560),
.B(n_555),
.Y(n_803)
);

INVx2_ASAP7_75t_L g804 ( 
.A(n_631),
.Y(n_804)
);

INVx2_ASAP7_75t_L g805 ( 
.A(n_634),
.Y(n_805)
);

NAND2xp5_ASAP7_75t_SL g806 ( 
.A(n_645),
.B(n_263),
.Y(n_806)
);

NAND2xp5_ASAP7_75t_L g807 ( 
.A(n_647),
.B(n_560),
.Y(n_807)
);

NAND2xp5_ASAP7_75t_L g808 ( 
.A(n_665),
.B(n_316),
.Y(n_808)
);

NAND2xp5_ASAP7_75t_SL g809 ( 
.A(n_645),
.B(n_325),
.Y(n_809)
);

INVx2_ASAP7_75t_L g810 ( 
.A(n_634),
.Y(n_810)
);

OAI221xp5_ASAP7_75t_L g811 ( 
.A1(n_668),
.A2(n_578),
.B1(n_574),
.B2(n_561),
.C(n_377),
.Y(n_811)
);

NAND2xp5_ASAP7_75t_SL g812 ( 
.A(n_645),
.B(n_339),
.Y(n_812)
);

INVx2_ASAP7_75t_L g813 ( 
.A(n_644),
.Y(n_813)
);

AOI21xp5_ASAP7_75t_L g814 ( 
.A1(n_587),
.A2(n_574),
.B(n_561),
.Y(n_814)
);

INVx2_ASAP7_75t_L g815 ( 
.A(n_644),
.Y(n_815)
);

INVx1_ASAP7_75t_L g816 ( 
.A(n_670),
.Y(n_816)
);

NAND2xp5_ASAP7_75t_L g817 ( 
.A(n_675),
.B(n_351),
.Y(n_817)
);

INVx2_ASAP7_75t_L g818 ( 
.A(n_649),
.Y(n_818)
);

NOR2xp33_ASAP7_75t_SL g819 ( 
.A(n_719),
.B(n_236),
.Y(n_819)
);

INVx2_ASAP7_75t_SL g820 ( 
.A(n_626),
.Y(n_820)
);

INVxp67_ASAP7_75t_L g821 ( 
.A(n_680),
.Y(n_821)
);

AND2x2_ASAP7_75t_SL g822 ( 
.A(n_600),
.B(n_360),
.Y(n_822)
);

NAND2xp5_ASAP7_75t_L g823 ( 
.A(n_699),
.B(n_373),
.Y(n_823)
);

AOI22xp33_ASAP7_75t_L g824 ( 
.A1(n_664),
.A2(n_394),
.B1(n_375),
.B2(n_561),
.Y(n_824)
);

NAND2xp5_ASAP7_75t_SL g825 ( 
.A(n_682),
.B(n_275),
.Y(n_825)
);

NAND2xp33_ASAP7_75t_L g826 ( 
.A(n_664),
.B(n_205),
.Y(n_826)
);

NAND2xp5_ASAP7_75t_L g827 ( 
.A(n_703),
.B(n_574),
.Y(n_827)
);

NAND2xp5_ASAP7_75t_L g828 ( 
.A(n_723),
.B(n_578),
.Y(n_828)
);

NAND2xp5_ASAP7_75t_SL g829 ( 
.A(n_635),
.B(n_658),
.Y(n_829)
);

INVx2_ASAP7_75t_SL g830 ( 
.A(n_628),
.Y(n_830)
);

INVx3_ASAP7_75t_L g831 ( 
.A(n_673),
.Y(n_831)
);

OAI22xp33_ASAP7_75t_L g832 ( 
.A1(n_628),
.A2(n_314),
.B1(n_367),
.B2(n_215),
.Y(n_832)
);

O2A1O1Ixp33_ASAP7_75t_L g833 ( 
.A1(n_600),
.A2(n_578),
.B(n_528),
.C(n_526),
.Y(n_833)
);

INVx2_ASAP7_75t_L g834 ( 
.A(n_649),
.Y(n_834)
);

NAND2xp5_ASAP7_75t_L g835 ( 
.A(n_658),
.B(n_525),
.Y(n_835)
);

INVx5_ASAP7_75t_L g836 ( 
.A(n_667),
.Y(n_836)
);

OAI22xp5_ASAP7_75t_L g837 ( 
.A1(n_660),
.A2(n_237),
.B1(n_239),
.B2(n_399),
.Y(n_837)
);

NOR2xp33_ASAP7_75t_L g838 ( 
.A(n_688),
.B(n_211),
.Y(n_838)
);

INVx3_ASAP7_75t_L g839 ( 
.A(n_673),
.Y(n_839)
);

INVx3_ASAP7_75t_L g840 ( 
.A(n_700),
.Y(n_840)
);

INVx4_ASAP7_75t_L g841 ( 
.A(n_660),
.Y(n_841)
);

NAND2xp5_ASAP7_75t_L g842 ( 
.A(n_588),
.B(n_596),
.Y(n_842)
);

INVx3_ASAP7_75t_L g843 ( 
.A(n_700),
.Y(n_843)
);

INVx2_ASAP7_75t_L g844 ( 
.A(n_651),
.Y(n_844)
);

O2A1O1Ixp5_ASAP7_75t_L g845 ( 
.A1(n_657),
.A2(n_669),
.B(n_725),
.C(n_713),
.Y(n_845)
);

NOR2xp33_ASAP7_75t_L g846 ( 
.A(n_639),
.B(n_211),
.Y(n_846)
);

INVx2_ASAP7_75t_L g847 ( 
.A(n_651),
.Y(n_847)
);

NAND2xp5_ASAP7_75t_L g848 ( 
.A(n_726),
.B(n_525),
.Y(n_848)
);

INVx1_ASAP7_75t_L g849 ( 
.A(n_722),
.Y(n_849)
);

OR2x2_ASAP7_75t_L g850 ( 
.A(n_641),
.B(n_219),
.Y(n_850)
);

AOI22xp33_ASAP7_75t_L g851 ( 
.A1(n_664),
.A2(n_207),
.B1(n_353),
.B2(n_521),
.Y(n_851)
);

INVx2_ASAP7_75t_L g852 ( 
.A(n_652),
.Y(n_852)
);

AND2x6_ASAP7_75t_SL g853 ( 
.A(n_694),
.B(n_334),
.Y(n_853)
);

AOI22xp33_ASAP7_75t_L g854 ( 
.A1(n_664),
.A2(n_207),
.B1(n_353),
.B2(n_521),
.Y(n_854)
);

HB1xp67_ASAP7_75t_L g855 ( 
.A(n_628),
.Y(n_855)
);

NAND2xp5_ASAP7_75t_L g856 ( 
.A(n_650),
.B(n_520),
.Y(n_856)
);

NAND2xp5_ASAP7_75t_SL g857 ( 
.A(n_722),
.B(n_277),
.Y(n_857)
);

OAI221xp5_ASAP7_75t_L g858 ( 
.A1(n_621),
.A2(n_628),
.B1(n_609),
.B2(n_622),
.C(n_616),
.Y(n_858)
);

NAND2xp5_ASAP7_75t_L g859 ( 
.A(n_650),
.B(n_520),
.Y(n_859)
);

NAND2xp5_ASAP7_75t_L g860 ( 
.A(n_650),
.B(n_526),
.Y(n_860)
);

NAND2xp5_ASAP7_75t_L g861 ( 
.A(n_655),
.B(n_528),
.Y(n_861)
);

NOR2xp67_ASAP7_75t_L g862 ( 
.A(n_633),
.B(n_279),
.Y(n_862)
);

NAND2xp5_ASAP7_75t_L g863 ( 
.A(n_655),
.B(n_282),
.Y(n_863)
);

INVx2_ASAP7_75t_L g864 ( 
.A(n_652),
.Y(n_864)
);

NAND2xp5_ASAP7_75t_SL g865 ( 
.A(n_655),
.B(n_291),
.Y(n_865)
);

NAND2xp5_ASAP7_75t_SL g866 ( 
.A(n_653),
.B(n_296),
.Y(n_866)
);

AOI22xp33_ASAP7_75t_L g867 ( 
.A1(n_664),
.A2(n_353),
.B1(n_400),
.B2(n_235),
.Y(n_867)
);

INVxp67_ASAP7_75t_L g868 ( 
.A(n_656),
.Y(n_868)
);

AOI22xp33_ASAP7_75t_L g869 ( 
.A1(n_711),
.A2(n_219),
.B1(n_365),
.B2(n_364),
.Y(n_869)
);

NOR2xp33_ASAP7_75t_L g870 ( 
.A(n_730),
.B(n_213),
.Y(n_870)
);

AND2x6_ASAP7_75t_SL g871 ( 
.A(n_629),
.B(n_358),
.Y(n_871)
);

BUFx3_ASAP7_75t_L g872 ( 
.A(n_698),
.Y(n_872)
);

INVx2_ASAP7_75t_SL g873 ( 
.A(n_711),
.Y(n_873)
);

NAND2xp5_ASAP7_75t_SL g874 ( 
.A(n_653),
.B(n_300),
.Y(n_874)
);

NAND2xp5_ASAP7_75t_L g875 ( 
.A(n_697),
.B(n_721),
.Y(n_875)
);

AOI22xp33_ASAP7_75t_L g876 ( 
.A1(n_711),
.A2(n_666),
.B1(n_690),
.B2(n_721),
.Y(n_876)
);

NAND2xp5_ASAP7_75t_L g877 ( 
.A(n_697),
.B(n_610),
.Y(n_877)
);

NAND2xp5_ASAP7_75t_L g878 ( 
.A(n_610),
.B(n_312),
.Y(n_878)
);

AOI22xp5_ASAP7_75t_L g879 ( 
.A1(n_704),
.A2(n_621),
.B1(n_666),
.B2(n_690),
.Y(n_879)
);

INVx1_ASAP7_75t_L g880 ( 
.A(n_729),
.Y(n_880)
);

INVx2_ASAP7_75t_L g881 ( 
.A(n_729),
.Y(n_881)
);

INVx1_ASAP7_75t_L g882 ( 
.A(n_590),
.Y(n_882)
);

INVx1_ASAP7_75t_L g883 ( 
.A(n_590),
.Y(n_883)
);

OAI22xp5_ASAP7_75t_L g884 ( 
.A1(n_698),
.A2(n_216),
.B1(n_399),
.B2(n_398),
.Y(n_884)
);

NAND2xp5_ASAP7_75t_L g885 ( 
.A(n_610),
.B(n_319),
.Y(n_885)
);

NOR3xp33_ASAP7_75t_L g886 ( 
.A(n_611),
.B(n_340),
.C(n_392),
.Y(n_886)
);

NAND2xp5_ASAP7_75t_L g887 ( 
.A(n_654),
.B(n_659),
.Y(n_887)
);

INVxp67_ASAP7_75t_L g888 ( 
.A(n_692),
.Y(n_888)
);

OAI22xp33_ASAP7_75t_L g889 ( 
.A1(n_629),
.A2(n_400),
.B1(n_226),
.B2(n_235),
.Y(n_889)
);

NOR2xp33_ASAP7_75t_L g890 ( 
.A(n_676),
.B(n_213),
.Y(n_890)
);

NOR2xp33_ASAP7_75t_L g891 ( 
.A(n_629),
.B(n_214),
.Y(n_891)
);

NAND2xp5_ASAP7_75t_SL g892 ( 
.A(n_663),
.B(n_327),
.Y(n_892)
);

NAND2xp5_ASAP7_75t_SL g893 ( 
.A(n_663),
.B(n_328),
.Y(n_893)
);

NAND2xp5_ASAP7_75t_L g894 ( 
.A(n_654),
.B(n_329),
.Y(n_894)
);

OR2x2_ASAP7_75t_L g895 ( 
.A(n_648),
.B(n_226),
.Y(n_895)
);

INVx8_ASAP7_75t_L g896 ( 
.A(n_629),
.Y(n_896)
);

INVx1_ASAP7_75t_L g897 ( 
.A(n_591),
.Y(n_897)
);

AOI22xp5_ASAP7_75t_L g898 ( 
.A1(n_691),
.A2(n_330),
.B1(n_397),
.B2(n_336),
.Y(n_898)
);

NAND2xp5_ASAP7_75t_L g899 ( 
.A(n_654),
.B(n_343),
.Y(n_899)
);

OAI21xp5_ASAP7_75t_L g900 ( 
.A1(n_757),
.A2(n_727),
.B(n_674),
.Y(n_900)
);

AOI21xp5_ASAP7_75t_L g901 ( 
.A1(n_829),
.A2(n_708),
.B(n_717),
.Y(n_901)
);

OAI22xp5_ASAP7_75t_L g902 ( 
.A1(n_858),
.A2(n_698),
.B1(n_702),
.B2(n_719),
.Y(n_902)
);

AOI21xp5_ASAP7_75t_L g903 ( 
.A1(n_829),
.A2(n_708),
.B(n_717),
.Y(n_903)
);

AOI21xp5_ASAP7_75t_L g904 ( 
.A1(n_759),
.A2(n_728),
.B(n_693),
.Y(n_904)
);

NOR2xp33_ASAP7_75t_L g905 ( 
.A(n_799),
.B(n_705),
.Y(n_905)
);

AOI21xp5_ASAP7_75t_L g906 ( 
.A1(n_761),
.A2(n_728),
.B(n_686),
.Y(n_906)
);

O2A1O1Ixp33_ASAP7_75t_SL g907 ( 
.A1(n_781),
.A2(n_782),
.B(n_806),
.C(n_792),
.Y(n_907)
);

NOR2xp33_ASAP7_75t_L g908 ( 
.A(n_821),
.B(n_677),
.Y(n_908)
);

AOI21xp5_ASAP7_75t_L g909 ( 
.A1(n_762),
.A2(n_683),
.B(n_674),
.Y(n_909)
);

NAND2xp5_ASAP7_75t_L g910 ( 
.A(n_785),
.B(n_659),
.Y(n_910)
);

O2A1O1Ixp33_ASAP7_75t_L g911 ( 
.A1(n_756),
.A2(n_601),
.B(n_591),
.C(n_683),
.Y(n_911)
);

NAND2xp5_ASAP7_75t_L g912 ( 
.A(n_787),
.B(n_659),
.Y(n_912)
);

AOI21xp5_ASAP7_75t_L g913 ( 
.A1(n_835),
.A2(n_686),
.B(n_693),
.Y(n_913)
);

NOR3xp33_ASAP7_75t_L g914 ( 
.A(n_746),
.B(n_237),
.C(n_398),
.Y(n_914)
);

AND2x4_ASAP7_75t_L g915 ( 
.A(n_796),
.B(n_797),
.Y(n_915)
);

AND2x2_ASAP7_75t_L g916 ( 
.A(n_765),
.B(n_779),
.Y(n_916)
);

AND2x2_ASAP7_75t_L g917 ( 
.A(n_800),
.B(n_606),
.Y(n_917)
);

AOI21xp5_ASAP7_75t_L g918 ( 
.A1(n_737),
.A2(n_696),
.B(n_695),
.Y(n_918)
);

INVx1_ASAP7_75t_L g919 ( 
.A(n_747),
.Y(n_919)
);

AOI21xp5_ASAP7_75t_L g920 ( 
.A1(n_735),
.A2(n_731),
.B(n_678),
.Y(n_920)
);

AOI21xp5_ASAP7_75t_L g921 ( 
.A1(n_781),
.A2(n_687),
.B(n_672),
.Y(n_921)
);

BUFx4f_ASAP7_75t_L g922 ( 
.A(n_896),
.Y(n_922)
);

NOR2x1_ASAP7_75t_R g923 ( 
.A(n_768),
.B(n_285),
.Y(n_923)
);

NAND2xp5_ASAP7_75t_SL g924 ( 
.A(n_767),
.B(n_606),
.Y(n_924)
);

INVx1_ASAP7_75t_L g925 ( 
.A(n_747),
.Y(n_925)
);

AOI21xp5_ASAP7_75t_L g926 ( 
.A1(n_782),
.A2(n_687),
.B(n_672),
.Y(n_926)
);

NAND2xp5_ASAP7_75t_L g927 ( 
.A(n_783),
.B(n_662),
.Y(n_927)
);

AOI21xp5_ASAP7_75t_L g928 ( 
.A1(n_792),
.A2(n_809),
.B(n_806),
.Y(n_928)
);

AO21x1_ASAP7_75t_L g929 ( 
.A1(n_770),
.A2(n_601),
.B(n_691),
.Y(n_929)
);

NOR2xp33_ASAP7_75t_L g930 ( 
.A(n_744),
.B(n_606),
.Y(n_930)
);

A2O1A1Ixp33_ASAP7_75t_L g931 ( 
.A1(n_776),
.A2(n_801),
.B(n_846),
.C(n_794),
.Y(n_931)
);

AOI21xp5_ASAP7_75t_L g932 ( 
.A1(n_809),
.A2(n_812),
.B(n_741),
.Y(n_932)
);

AOI22xp5_ASAP7_75t_L g933 ( 
.A1(n_873),
.A2(n_731),
.B1(n_691),
.B2(n_637),
.Y(n_933)
);

AOI21xp5_ASAP7_75t_L g934 ( 
.A1(n_812),
.A2(n_687),
.B(n_667),
.Y(n_934)
);

NAND2xp5_ASAP7_75t_L g935 ( 
.A(n_795),
.B(n_678),
.Y(n_935)
);

NAND2xp5_ASAP7_75t_L g936 ( 
.A(n_739),
.B(n_678),
.Y(n_936)
);

BUFx12f_ASAP7_75t_L g937 ( 
.A(n_871),
.Y(n_937)
);

NAND2xp5_ASAP7_75t_SL g938 ( 
.A(n_767),
.B(n_637),
.Y(n_938)
);

O2A1O1Ixp5_ASAP7_75t_L g939 ( 
.A1(n_825),
.A2(n_685),
.B(n_706),
.C(n_710),
.Y(n_939)
);

AOI21xp5_ASAP7_75t_L g940 ( 
.A1(n_803),
.A2(n_814),
.B(n_887),
.Y(n_940)
);

AOI21xp5_ASAP7_75t_L g941 ( 
.A1(n_836),
.A2(n_841),
.B(n_877),
.Y(n_941)
);

AOI21xp5_ASAP7_75t_L g942 ( 
.A1(n_836),
.A2(n_841),
.B(n_848),
.Y(n_942)
);

OR2x6_ASAP7_75t_L g943 ( 
.A(n_896),
.B(n_732),
.Y(n_943)
);

AOI21xp5_ASAP7_75t_L g944 ( 
.A1(n_836),
.A2(n_672),
.B(n_710),
.Y(n_944)
);

NAND3xp33_ASAP7_75t_SL g945 ( 
.A(n_778),
.B(n_734),
.C(n_701),
.Y(n_945)
);

O2A1O1Ixp33_ASAP7_75t_L g946 ( 
.A1(n_756),
.A2(n_685),
.B(n_724),
.C(n_707),
.Y(n_946)
);

INVx1_ASAP7_75t_SL g947 ( 
.A(n_790),
.Y(n_947)
);

NAND2xp5_ASAP7_75t_L g948 ( 
.A(n_873),
.B(n_685),
.Y(n_948)
);

NAND2x1_ASAP7_75t_L g949 ( 
.A(n_767),
.B(n_667),
.Y(n_949)
);

NOR2xp33_ASAP7_75t_L g950 ( 
.A(n_777),
.B(n_637),
.Y(n_950)
);

OAI22xp5_ASAP7_75t_L g951 ( 
.A1(n_841),
.A2(n_366),
.B1(n_216),
.B2(n_218),
.Y(n_951)
);

A2O1A1Ixp33_ASAP7_75t_L g952 ( 
.A1(n_870),
.A2(n_366),
.B(n_218),
.C(n_227),
.Y(n_952)
);

INVx2_ASAP7_75t_L g953 ( 
.A(n_763),
.Y(n_953)
);

AND2x2_ASAP7_75t_L g954 ( 
.A(n_775),
.B(n_732),
.Y(n_954)
);

INVx4_ASAP7_75t_L g955 ( 
.A(n_767),
.Y(n_955)
);

NOR2xp67_ASAP7_75t_L g956 ( 
.A(n_888),
.B(n_368),
.Y(n_956)
);

NAND2xp5_ASAP7_75t_SL g957 ( 
.A(n_820),
.B(n_732),
.Y(n_957)
);

AOI21x1_ASAP7_75t_L g958 ( 
.A1(n_875),
.A2(n_672),
.B(n_710),
.Y(n_958)
);

AOI21xp5_ASAP7_75t_L g959 ( 
.A1(n_876),
.A2(n_710),
.B(n_667),
.Y(n_959)
);

AOI21xp5_ASAP7_75t_L g960 ( 
.A1(n_836),
.A2(n_687),
.B(n_372),
.Y(n_960)
);

NAND2xp5_ASAP7_75t_L g961 ( 
.A(n_736),
.B(n_738),
.Y(n_961)
);

INVx1_ASAP7_75t_L g962 ( 
.A(n_763),
.Y(n_962)
);

OAI22xp5_ASAP7_75t_L g963 ( 
.A1(n_879),
.A2(n_362),
.B1(n_227),
.B2(n_234),
.Y(n_963)
);

NAND2xp5_ASAP7_75t_L g964 ( 
.A(n_740),
.B(n_370),
.Y(n_964)
);

NAND2xp5_ASAP7_75t_L g965 ( 
.A(n_758),
.B(n_387),
.Y(n_965)
);

AND2x2_ASAP7_75t_L g966 ( 
.A(n_755),
.B(n_707),
.Y(n_966)
);

AOI21xp5_ASAP7_75t_L g967 ( 
.A1(n_836),
.A2(n_214),
.B(n_234),
.Y(n_967)
);

AOI21xp5_ASAP7_75t_L g968 ( 
.A1(n_878),
.A2(n_894),
.B(n_885),
.Y(n_968)
);

NAND2xp5_ASAP7_75t_L g969 ( 
.A(n_772),
.B(n_784),
.Y(n_969)
);

NAND3xp33_ASAP7_75t_SL g970 ( 
.A(n_838),
.B(n_734),
.C(n_724),
.Y(n_970)
);

INVx3_ASAP7_75t_L g971 ( 
.A(n_831),
.Y(n_971)
);

NAND2xp5_ASAP7_75t_SL g972 ( 
.A(n_890),
.B(n_239),
.Y(n_972)
);

AOI21xp5_ASAP7_75t_L g973 ( 
.A1(n_899),
.A2(n_381),
.B(n_347),
.Y(n_973)
);

INVx1_ASAP7_75t_L g974 ( 
.A(n_764),
.Y(n_974)
);

AND2x2_ASAP7_75t_L g975 ( 
.A(n_868),
.B(n_358),
.Y(n_975)
);

OAI21xp5_ASAP7_75t_L g976 ( 
.A1(n_845),
.A2(n_706),
.B(n_347),
.Y(n_976)
);

AOI21x1_ASAP7_75t_L g977 ( 
.A1(n_745),
.A2(n_706),
.B(n_384),
.Y(n_977)
);

AOI21xp5_ASAP7_75t_L g978 ( 
.A1(n_766),
.A2(n_362),
.B(n_352),
.Y(n_978)
);

NAND2xp5_ASAP7_75t_L g979 ( 
.A(n_816),
.B(n_352),
.Y(n_979)
);

OAI321xp33_ASAP7_75t_L g980 ( 
.A1(n_832),
.A2(n_358),
.A3(n_346),
.B1(n_349),
.B2(n_350),
.C(n_357),
.Y(n_980)
);

AND2x2_ASAP7_75t_L g981 ( 
.A(n_850),
.B(n_349),
.Y(n_981)
);

AOI22xp33_ASAP7_75t_L g982 ( 
.A1(n_822),
.A2(n_706),
.B1(n_354),
.B2(n_355),
.Y(n_982)
);

NOR2xp33_ASAP7_75t_L g983 ( 
.A(n_895),
.B(n_780),
.Y(n_983)
);

OAI22xp5_ASAP7_75t_L g984 ( 
.A1(n_831),
.A2(n_356),
.B1(n_355),
.B2(n_363),
.Y(n_984)
);

HB1xp67_ASAP7_75t_L g985 ( 
.A(n_855),
.Y(n_985)
);

AND2x2_ASAP7_75t_L g986 ( 
.A(n_768),
.B(n_350),
.Y(n_986)
);

AOI21xp5_ASAP7_75t_L g987 ( 
.A1(n_752),
.A2(n_354),
.B(n_356),
.Y(n_987)
);

AOI21xp5_ASAP7_75t_L g988 ( 
.A1(n_753),
.A2(n_363),
.B(n_381),
.Y(n_988)
);

NAND2xp5_ASAP7_75t_L g989 ( 
.A(n_856),
.B(n_383),
.Y(n_989)
);

NAND2xp5_ASAP7_75t_L g990 ( 
.A(n_859),
.B(n_383),
.Y(n_990)
);

AOI21xp5_ASAP7_75t_L g991 ( 
.A1(n_769),
.A2(n_384),
.B(n_391),
.Y(n_991)
);

AND2x2_ASAP7_75t_L g992 ( 
.A(n_869),
.B(n_364),
.Y(n_992)
);

AOI22xp33_ASAP7_75t_L g993 ( 
.A1(n_822),
.A2(n_706),
.B1(n_385),
.B2(n_376),
.Y(n_993)
);

A2O1A1Ixp33_ASAP7_75t_L g994 ( 
.A1(n_748),
.A2(n_374),
.B(n_369),
.C(n_341),
.Y(n_994)
);

A2O1A1Ixp33_ASAP7_75t_L g995 ( 
.A1(n_860),
.A2(n_361),
.B(n_359),
.C(n_357),
.Y(n_995)
);

NOR2xp33_ASAP7_75t_L g996 ( 
.A(n_786),
.B(n_361),
.Y(n_996)
);

O2A1O1Ixp33_ASAP7_75t_L g997 ( 
.A1(n_837),
.A2(n_359),
.B(n_9),
.C(n_10),
.Y(n_997)
);

AND2x2_ASAP7_75t_L g998 ( 
.A(n_891),
.B(n_7),
.Y(n_998)
);

AO21x1_ASAP7_75t_L g999 ( 
.A1(n_892),
.A2(n_11),
.B(n_13),
.Y(n_999)
);

NOR2xp33_ASAP7_75t_L g1000 ( 
.A(n_796),
.B(n_11),
.Y(n_1000)
);

NAND2xp5_ASAP7_75t_L g1001 ( 
.A(n_861),
.B(n_15),
.Y(n_1001)
);

NAND2xp5_ASAP7_75t_L g1002 ( 
.A(n_771),
.B(n_774),
.Y(n_1002)
);

NAND2xp5_ASAP7_75t_SL g1003 ( 
.A(n_793),
.B(n_68),
.Y(n_1003)
);

BUFx6f_ASAP7_75t_L g1004 ( 
.A(n_797),
.Y(n_1004)
);

OAI21xp5_ASAP7_75t_L g1005 ( 
.A1(n_771),
.A2(n_74),
.B(n_192),
.Y(n_1005)
);

NAND2xp5_ASAP7_75t_L g1006 ( 
.A(n_774),
.B(n_16),
.Y(n_1006)
);

INVxp67_ASAP7_75t_L g1007 ( 
.A(n_865),
.Y(n_1007)
);

OAI21xp5_ASAP7_75t_L g1008 ( 
.A1(n_789),
.A2(n_195),
.B(n_190),
.Y(n_1008)
);

OAI22xp5_ASAP7_75t_L g1009 ( 
.A1(n_831),
.A2(n_183),
.B1(n_182),
.B2(n_169),
.Y(n_1009)
);

AND2x2_ASAP7_75t_L g1010 ( 
.A(n_862),
.B(n_16),
.Y(n_1010)
);

BUFx6f_ASAP7_75t_L g1011 ( 
.A(n_872),
.Y(n_1011)
);

AOI22xp5_ASAP7_75t_L g1012 ( 
.A1(n_857),
.A2(n_158),
.B1(n_151),
.B2(n_144),
.Y(n_1012)
);

AOI21xp5_ASAP7_75t_L g1013 ( 
.A1(n_788),
.A2(n_131),
.B(n_126),
.Y(n_1013)
);

AOI21xp5_ASAP7_75t_L g1014 ( 
.A1(n_798),
.A2(n_120),
.B(n_116),
.Y(n_1014)
);

OAI22xp5_ASAP7_75t_L g1015 ( 
.A1(n_839),
.A2(n_114),
.B1(n_113),
.B2(n_111),
.Y(n_1015)
);

AOI21xp5_ASAP7_75t_L g1016 ( 
.A1(n_807),
.A2(n_828),
.B(n_827),
.Y(n_1016)
);

NOR2xp33_ASAP7_75t_R g1017 ( 
.A(n_819),
.B(n_105),
.Y(n_1017)
);

AOI21xp5_ASAP7_75t_L g1018 ( 
.A1(n_842),
.A2(n_103),
.B(n_82),
.Y(n_1018)
);

AOI21xp5_ASAP7_75t_L g1019 ( 
.A1(n_892),
.A2(n_19),
.B(n_21),
.Y(n_1019)
);

AOI221xp5_ASAP7_75t_L g1020 ( 
.A1(n_889),
.A2(n_23),
.B1(n_28),
.B2(n_29),
.C(n_31),
.Y(n_1020)
);

AOI21xp5_ASAP7_75t_L g1021 ( 
.A1(n_893),
.A2(n_29),
.B(n_32),
.Y(n_1021)
);

A2O1A1Ixp33_ASAP7_75t_L g1022 ( 
.A1(n_898),
.A2(n_36),
.B(n_37),
.C(n_41),
.Y(n_1022)
);

OAI21xp5_ASAP7_75t_L g1023 ( 
.A1(n_791),
.A2(n_48),
.B(n_49),
.Y(n_1023)
);

BUFx12f_ASAP7_75t_L g1024 ( 
.A(n_853),
.Y(n_1024)
);

INVx3_ASAP7_75t_L g1025 ( 
.A(n_839),
.Y(n_1025)
);

AOI21xp5_ASAP7_75t_L g1026 ( 
.A1(n_893),
.A2(n_49),
.B(n_51),
.Y(n_1026)
);

INVxp67_ASAP7_75t_L g1027 ( 
.A(n_865),
.Y(n_1027)
);

BUFx2_ASAP7_75t_L g1028 ( 
.A(n_830),
.Y(n_1028)
);

INVx3_ASAP7_75t_L g1029 ( 
.A(n_839),
.Y(n_1029)
);

NAND2xp5_ASAP7_75t_L g1030 ( 
.A(n_791),
.B(n_51),
.Y(n_1030)
);

O2A1O1Ixp33_ASAP7_75t_L g1031 ( 
.A1(n_866),
.A2(n_53),
.B(n_55),
.C(n_56),
.Y(n_1031)
);

INVx2_ASAP7_75t_L g1032 ( 
.A(n_804),
.Y(n_1032)
);

AOI21xp5_ASAP7_75t_L g1033 ( 
.A1(n_857),
.A2(n_56),
.B(n_57),
.Y(n_1033)
);

NAND2xp5_ASAP7_75t_SL g1034 ( 
.A(n_872),
.B(n_57),
.Y(n_1034)
);

NOR2xp33_ASAP7_75t_L g1035 ( 
.A(n_863),
.B(n_58),
.Y(n_1035)
);

NOR2xp33_ASAP7_75t_SL g1036 ( 
.A(n_896),
.B(n_58),
.Y(n_1036)
);

AOI21xp5_ASAP7_75t_L g1037 ( 
.A1(n_804),
.A2(n_60),
.B(n_852),
.Y(n_1037)
);

AOI21x1_ASAP7_75t_L g1038 ( 
.A1(n_749),
.A2(n_754),
.B(n_751),
.Y(n_1038)
);

AOI21xp5_ASAP7_75t_L g1039 ( 
.A1(n_840),
.A2(n_843),
.B(n_826),
.Y(n_1039)
);

AND2x2_ASAP7_75t_L g1040 ( 
.A(n_743),
.B(n_886),
.Y(n_1040)
);

NOR2x1_ASAP7_75t_L g1041 ( 
.A(n_840),
.B(n_843),
.Y(n_1041)
);

AOI21x1_ASAP7_75t_L g1042 ( 
.A1(n_749),
.A2(n_754),
.B(n_751),
.Y(n_1042)
);

NAND2xp5_ASAP7_75t_SL g1043 ( 
.A(n_802),
.B(n_867),
.Y(n_1043)
);

AOI21xp5_ASAP7_75t_L g1044 ( 
.A1(n_840),
.A2(n_843),
.B(n_826),
.Y(n_1044)
);

AOI21xp5_ASAP7_75t_L g1045 ( 
.A1(n_760),
.A2(n_849),
.B(n_815),
.Y(n_1045)
);

AOI21xp5_ASAP7_75t_L g1046 ( 
.A1(n_805),
.A2(n_834),
.B(n_844),
.Y(n_1046)
);

AOI21xp5_ASAP7_75t_L g1047 ( 
.A1(n_810),
.A2(n_847),
.B(n_818),
.Y(n_1047)
);

INVx3_ASAP7_75t_L g1048 ( 
.A(n_810),
.Y(n_1048)
);

NAND2xp5_ASAP7_75t_L g1049 ( 
.A(n_813),
.B(n_864),
.Y(n_1049)
);

AND2x2_ASAP7_75t_L g1050 ( 
.A(n_750),
.B(n_874),
.Y(n_1050)
);

OAI22xp5_ASAP7_75t_L g1051 ( 
.A1(n_851),
.A2(n_854),
.B1(n_824),
.B2(n_773),
.Y(n_1051)
);

NAND2xp5_ASAP7_75t_L g1052 ( 
.A(n_815),
.B(n_852),
.Y(n_1052)
);

NOR2xp33_ASAP7_75t_L g1053 ( 
.A(n_884),
.B(n_823),
.Y(n_1053)
);

AOI21xp5_ASAP7_75t_L g1054 ( 
.A1(n_818),
.A2(n_864),
.B(n_847),
.Y(n_1054)
);

NOR2xp33_ASAP7_75t_L g1055 ( 
.A(n_808),
.B(n_817),
.Y(n_1055)
);

OAI21xp5_ASAP7_75t_L g1056 ( 
.A1(n_881),
.A2(n_880),
.B(n_897),
.Y(n_1056)
);

AOI21xp5_ASAP7_75t_L g1057 ( 
.A1(n_881),
.A2(n_882),
.B(n_883),
.Y(n_1057)
);

NAND2xp5_ASAP7_75t_L g1058 ( 
.A(n_742),
.B(n_833),
.Y(n_1058)
);

AOI21xp5_ASAP7_75t_L g1059 ( 
.A1(n_896),
.A2(n_587),
.B(n_757),
.Y(n_1059)
);

AOI21x1_ASAP7_75t_L g1060 ( 
.A1(n_811),
.A2(n_825),
.B(n_642),
.Y(n_1060)
);

NAND2xp5_ASAP7_75t_L g1061 ( 
.A(n_785),
.B(n_602),
.Y(n_1061)
);

AOI21xp5_ASAP7_75t_L g1062 ( 
.A1(n_757),
.A2(n_587),
.B(n_759),
.Y(n_1062)
);

INVx4_ASAP7_75t_L g1063 ( 
.A(n_767),
.Y(n_1063)
);

A2O1A1Ixp33_ASAP7_75t_L g1064 ( 
.A1(n_776),
.A2(n_801),
.B(n_846),
.C(n_592),
.Y(n_1064)
);

NAND2xp5_ASAP7_75t_L g1065 ( 
.A(n_785),
.B(n_602),
.Y(n_1065)
);

OAI22xp5_ASAP7_75t_L g1066 ( 
.A1(n_858),
.A2(n_829),
.B1(n_841),
.B2(n_592),
.Y(n_1066)
);

NOR2xp33_ASAP7_75t_L g1067 ( 
.A(n_799),
.B(n_821),
.Y(n_1067)
);

INVx5_ASAP7_75t_L g1068 ( 
.A(n_767),
.Y(n_1068)
);

BUFx6f_ASAP7_75t_L g1069 ( 
.A(n_767),
.Y(n_1069)
);

NOR2xp67_ASAP7_75t_L g1070 ( 
.A(n_888),
.B(n_720),
.Y(n_1070)
);

NOR2xp33_ASAP7_75t_L g1071 ( 
.A(n_799),
.B(n_821),
.Y(n_1071)
);

NAND2xp5_ASAP7_75t_SL g1072 ( 
.A(n_767),
.B(n_787),
.Y(n_1072)
);

AOI21xp5_ASAP7_75t_L g1073 ( 
.A1(n_829),
.A2(n_587),
.B(n_757),
.Y(n_1073)
);

NAND2xp5_ASAP7_75t_L g1074 ( 
.A(n_785),
.B(n_602),
.Y(n_1074)
);

BUFx6f_ASAP7_75t_L g1075 ( 
.A(n_767),
.Y(n_1075)
);

NAND2xp5_ASAP7_75t_L g1076 ( 
.A(n_785),
.B(n_602),
.Y(n_1076)
);

NAND2x1p5_ASAP7_75t_L g1077 ( 
.A(n_1068),
.B(n_955),
.Y(n_1077)
);

AOI21xp5_ASAP7_75t_L g1078 ( 
.A1(n_940),
.A2(n_1044),
.B(n_1039),
.Y(n_1078)
);

OAI21xp33_ASAP7_75t_L g1079 ( 
.A1(n_996),
.A2(n_992),
.B(n_983),
.Y(n_1079)
);

NAND2xp5_ASAP7_75t_L g1080 ( 
.A(n_1061),
.B(n_1065),
.Y(n_1080)
);

AOI21xp5_ASAP7_75t_L g1081 ( 
.A1(n_1062),
.A2(n_1068),
.B(n_932),
.Y(n_1081)
);

BUFx4f_ASAP7_75t_L g1082 ( 
.A(n_943),
.Y(n_1082)
);

NAND2xp5_ASAP7_75t_L g1083 ( 
.A(n_1074),
.B(n_1076),
.Y(n_1083)
);

INVx1_ASAP7_75t_L g1084 ( 
.A(n_919),
.Y(n_1084)
);

NAND2xp5_ASAP7_75t_SL g1085 ( 
.A(n_954),
.B(n_1067),
.Y(n_1085)
);

NOR2x1_ASAP7_75t_L g1086 ( 
.A(n_917),
.B(n_955),
.Y(n_1086)
);

AOI21xp5_ASAP7_75t_L g1087 ( 
.A1(n_1068),
.A2(n_928),
.B(n_907),
.Y(n_1087)
);

HB1xp67_ASAP7_75t_L g1088 ( 
.A(n_985),
.Y(n_1088)
);

NAND2xp5_ASAP7_75t_L g1089 ( 
.A(n_1055),
.B(n_1064),
.Y(n_1089)
);

AO31x2_ASAP7_75t_L g1090 ( 
.A1(n_929),
.A2(n_931),
.A3(n_1066),
.B(n_999),
.Y(n_1090)
);

BUFx6f_ASAP7_75t_L g1091 ( 
.A(n_1069),
.Y(n_1091)
);

NAND2xp5_ASAP7_75t_L g1092 ( 
.A(n_1071),
.B(n_912),
.Y(n_1092)
);

INVx2_ASAP7_75t_L g1093 ( 
.A(n_1048),
.Y(n_1093)
);

OAI21xp5_ASAP7_75t_L g1094 ( 
.A1(n_1073),
.A2(n_906),
.B(n_904),
.Y(n_1094)
);

O2A1O1Ixp33_ASAP7_75t_L g1095 ( 
.A1(n_1022),
.A2(n_997),
.B(n_980),
.C(n_1043),
.Y(n_1095)
);

AOI21xp5_ASAP7_75t_L g1096 ( 
.A1(n_1068),
.A2(n_959),
.B(n_1073),
.Y(n_1096)
);

NAND2x1p5_ASAP7_75t_L g1097 ( 
.A(n_1063),
.B(n_1069),
.Y(n_1097)
);

OAI21x1_ASAP7_75t_SL g1098 ( 
.A1(n_946),
.A2(n_1023),
.B(n_1008),
.Y(n_1098)
);

INVx4_ASAP7_75t_L g1099 ( 
.A(n_1069),
.Y(n_1099)
);

NOR2xp33_ASAP7_75t_L g1100 ( 
.A(n_908),
.B(n_905),
.Y(n_1100)
);

INVx1_ASAP7_75t_L g1101 ( 
.A(n_925),
.Y(n_1101)
);

BUFx6f_ASAP7_75t_L g1102 ( 
.A(n_1075),
.Y(n_1102)
);

OAI21xp5_ASAP7_75t_L g1103 ( 
.A1(n_904),
.A2(n_906),
.B(n_913),
.Y(n_1103)
);

BUFx2_ASAP7_75t_L g1104 ( 
.A(n_966),
.Y(n_1104)
);

AOI21xp5_ASAP7_75t_L g1105 ( 
.A1(n_959),
.A2(n_968),
.B(n_1059),
.Y(n_1105)
);

AOI21xp5_ASAP7_75t_L g1106 ( 
.A1(n_1016),
.A2(n_910),
.B(n_936),
.Y(n_1106)
);

BUFx2_ASAP7_75t_L g1107 ( 
.A(n_947),
.Y(n_1107)
);

OAI21xp5_ASAP7_75t_L g1108 ( 
.A1(n_913),
.A2(n_909),
.B(n_903),
.Y(n_1108)
);

OAI21xp5_ASAP7_75t_L g1109 ( 
.A1(n_909),
.A2(n_903),
.B(n_901),
.Y(n_1109)
);

INVx3_ASAP7_75t_L g1110 ( 
.A(n_1075),
.Y(n_1110)
);

AOI21xp5_ASAP7_75t_L g1111 ( 
.A1(n_942),
.A2(n_901),
.B(n_1058),
.Y(n_1111)
);

OAI21x1_ASAP7_75t_SL g1112 ( 
.A1(n_1005),
.A2(n_1033),
.B(n_1021),
.Y(n_1112)
);

OAI21xp5_ASAP7_75t_L g1113 ( 
.A1(n_918),
.A2(n_911),
.B(n_939),
.Y(n_1113)
);

AOI21xp5_ASAP7_75t_L g1114 ( 
.A1(n_900),
.A2(n_1072),
.B(n_941),
.Y(n_1114)
);

BUFx2_ASAP7_75t_L g1115 ( 
.A(n_915),
.Y(n_1115)
);

AOI21xp5_ASAP7_75t_L g1116 ( 
.A1(n_1041),
.A2(n_949),
.B(n_920),
.Y(n_1116)
);

OAI21x1_ASAP7_75t_L g1117 ( 
.A1(n_1046),
.A2(n_1047),
.B(n_1054),
.Y(n_1117)
);

OAI22x1_ASAP7_75t_L g1118 ( 
.A1(n_1040),
.A2(n_1007),
.B1(n_1027),
.B2(n_933),
.Y(n_1118)
);

AO31x2_ASAP7_75t_L g1119 ( 
.A1(n_1037),
.A2(n_994),
.A3(n_1051),
.B(n_1035),
.Y(n_1119)
);

OAI21xp5_ASAP7_75t_L g1120 ( 
.A1(n_1002),
.A2(n_1049),
.B(n_1052),
.Y(n_1120)
);

OAI21xp5_ASAP7_75t_L g1121 ( 
.A1(n_1053),
.A2(n_1001),
.B(n_1045),
.Y(n_1121)
);

OAI21x1_ASAP7_75t_L g1122 ( 
.A1(n_921),
.A2(n_934),
.B(n_926),
.Y(n_1122)
);

AOI21xp5_ASAP7_75t_L g1123 ( 
.A1(n_948),
.A2(n_1056),
.B(n_971),
.Y(n_1123)
);

NAND2xp5_ASAP7_75t_L g1124 ( 
.A(n_961),
.B(n_969),
.Y(n_1124)
);

OAI21xp5_ASAP7_75t_L g1125 ( 
.A1(n_1057),
.A2(n_976),
.B(n_1060),
.Y(n_1125)
);

NAND2xp5_ASAP7_75t_L g1126 ( 
.A(n_927),
.B(n_971),
.Y(n_1126)
);

AO31x2_ASAP7_75t_L g1127 ( 
.A1(n_1037),
.A2(n_1006),
.A3(n_1030),
.B(n_902),
.Y(n_1127)
);

NAND2xp5_ASAP7_75t_L g1128 ( 
.A(n_1025),
.B(n_1029),
.Y(n_1128)
);

INVx1_ASAP7_75t_L g1129 ( 
.A(n_962),
.Y(n_1129)
);

NAND2xp5_ASAP7_75t_SL g1130 ( 
.A(n_1004),
.B(n_915),
.Y(n_1130)
);

NAND2xp5_ASAP7_75t_L g1131 ( 
.A(n_1048),
.B(n_974),
.Y(n_1131)
);

OAI21x1_ASAP7_75t_L g1132 ( 
.A1(n_1038),
.A2(n_1042),
.B(n_944),
.Y(n_1132)
);

BUFx2_ASAP7_75t_L g1133 ( 
.A(n_916),
.Y(n_1133)
);

AOI21xp5_ASAP7_75t_L g1134 ( 
.A1(n_1063),
.A2(n_1075),
.B(n_935),
.Y(n_1134)
);

NAND2xp5_ASAP7_75t_L g1135 ( 
.A(n_989),
.B(n_990),
.Y(n_1135)
);

OR2x2_ASAP7_75t_L g1136 ( 
.A(n_945),
.B(n_970),
.Y(n_1136)
);

A2O1A1Ixp33_ASAP7_75t_L g1137 ( 
.A1(n_998),
.A2(n_914),
.B(n_952),
.C(n_991),
.Y(n_1137)
);

O2A1O1Ixp5_ASAP7_75t_L g1138 ( 
.A1(n_972),
.A2(n_1003),
.B(n_977),
.C(n_987),
.Y(n_1138)
);

AND2x2_ASAP7_75t_L g1139 ( 
.A(n_981),
.B(n_986),
.Y(n_1139)
);

CKINVDCx5p33_ASAP7_75t_R g1140 ( 
.A(n_943),
.Y(n_1140)
);

BUFx2_ASAP7_75t_L g1141 ( 
.A(n_1004),
.Y(n_1141)
);

NOR2x1_ASAP7_75t_L g1142 ( 
.A(n_930),
.B(n_950),
.Y(n_1142)
);

NAND2xp5_ASAP7_75t_L g1143 ( 
.A(n_953),
.B(n_1032),
.Y(n_1143)
);

AND2x2_ASAP7_75t_SL g1144 ( 
.A(n_1036),
.B(n_922),
.Y(n_1144)
);

OAI21x1_ASAP7_75t_L g1145 ( 
.A1(n_1013),
.A2(n_1014),
.B(n_1018),
.Y(n_1145)
);

NAND2xp5_ASAP7_75t_L g1146 ( 
.A(n_1010),
.B(n_1050),
.Y(n_1146)
);

OAI21x1_ASAP7_75t_L g1147 ( 
.A1(n_1013),
.A2(n_1014),
.B(n_1018),
.Y(n_1147)
);

AOI21xp5_ASAP7_75t_L g1148 ( 
.A1(n_922),
.A2(n_965),
.B(n_964),
.Y(n_1148)
);

A2O1A1Ixp33_ASAP7_75t_L g1149 ( 
.A1(n_991),
.A2(n_1033),
.B(n_1026),
.C(n_1019),
.Y(n_1149)
);

OAI21x1_ASAP7_75t_L g1150 ( 
.A1(n_960),
.A2(n_1009),
.B(n_1015),
.Y(n_1150)
);

AO21x1_ASAP7_75t_L g1151 ( 
.A1(n_1031),
.A2(n_1019),
.B(n_1021),
.Y(n_1151)
);

NAND2xp5_ASAP7_75t_L g1152 ( 
.A(n_975),
.B(n_979),
.Y(n_1152)
);

OAI21x1_ASAP7_75t_L g1153 ( 
.A1(n_924),
.A2(n_938),
.B(n_987),
.Y(n_1153)
);

AOI21xp5_ASAP7_75t_L g1154 ( 
.A1(n_957),
.A2(n_973),
.B(n_1034),
.Y(n_1154)
);

AOI21xp5_ASAP7_75t_L g1155 ( 
.A1(n_1011),
.A2(n_1004),
.B(n_1012),
.Y(n_1155)
);

INVx5_ASAP7_75t_L g1156 ( 
.A(n_1011),
.Y(n_1156)
);

AOI21xp5_ASAP7_75t_L g1157 ( 
.A1(n_1011),
.A2(n_1070),
.B(n_988),
.Y(n_1157)
);

AO21x1_ASAP7_75t_L g1158 ( 
.A1(n_1026),
.A2(n_988),
.B(n_1000),
.Y(n_1158)
);

BUFx2_ASAP7_75t_L g1159 ( 
.A(n_1028),
.Y(n_1159)
);

AOI21xp5_ASAP7_75t_L g1160 ( 
.A1(n_978),
.A2(n_967),
.B(n_956),
.Y(n_1160)
);

NAND2xp5_ASAP7_75t_L g1161 ( 
.A(n_995),
.B(n_963),
.Y(n_1161)
);

OAI21xp5_ASAP7_75t_L g1162 ( 
.A1(n_993),
.A2(n_982),
.B(n_1020),
.Y(n_1162)
);

NAND2xp5_ASAP7_75t_L g1163 ( 
.A(n_951),
.B(n_984),
.Y(n_1163)
);

AO31x2_ASAP7_75t_L g1164 ( 
.A1(n_1020),
.A2(n_1017),
.A3(n_943),
.B(n_923),
.Y(n_1164)
);

OAI21xp5_ASAP7_75t_L g1165 ( 
.A1(n_937),
.A2(n_1064),
.B(n_1073),
.Y(n_1165)
);

NAND2x1p5_ASAP7_75t_L g1166 ( 
.A(n_1024),
.B(n_1068),
.Y(n_1166)
);

A2O1A1Ixp33_ASAP7_75t_L g1167 ( 
.A1(n_1064),
.A2(n_931),
.B(n_1035),
.C(n_1053),
.Y(n_1167)
);

NAND3xp33_ASAP7_75t_SL g1168 ( 
.A(n_914),
.B(n_583),
.C(n_545),
.Y(n_1168)
);

NAND2xp5_ASAP7_75t_L g1169 ( 
.A(n_1061),
.B(n_1065),
.Y(n_1169)
);

A2O1A1Ixp33_ASAP7_75t_L g1170 ( 
.A1(n_1064),
.A2(n_931),
.B(n_1035),
.C(n_1053),
.Y(n_1170)
);

INVx3_ASAP7_75t_L g1171 ( 
.A(n_1069),
.Y(n_1171)
);

BUFx3_ASAP7_75t_L g1172 ( 
.A(n_917),
.Y(n_1172)
);

HB1xp67_ASAP7_75t_L g1173 ( 
.A(n_985),
.Y(n_1173)
);

OAI21x1_ASAP7_75t_L g1174 ( 
.A1(n_909),
.A2(n_913),
.B(n_918),
.Y(n_1174)
);

NAND2xp33_ASAP7_75t_SL g1175 ( 
.A(n_1017),
.B(n_768),
.Y(n_1175)
);

NOR2xp33_ASAP7_75t_L g1176 ( 
.A(n_1067),
.B(n_1071),
.Y(n_1176)
);

OAI21xp5_ASAP7_75t_L g1177 ( 
.A1(n_1064),
.A2(n_1073),
.B(n_1062),
.Y(n_1177)
);

NAND2xp5_ASAP7_75t_L g1178 ( 
.A(n_1061),
.B(n_1065),
.Y(n_1178)
);

NAND2xp5_ASAP7_75t_SL g1179 ( 
.A(n_954),
.B(n_800),
.Y(n_1179)
);

AND2x2_ASAP7_75t_L g1180 ( 
.A(n_954),
.B(n_779),
.Y(n_1180)
);

BUFx6f_ASAP7_75t_L g1181 ( 
.A(n_1069),
.Y(n_1181)
);

NAND2xp5_ASAP7_75t_L g1182 ( 
.A(n_1061),
.B(n_1065),
.Y(n_1182)
);

NAND2x1p5_ASAP7_75t_L g1183 ( 
.A(n_1068),
.B(n_955),
.Y(n_1183)
);

AO21x1_ASAP7_75t_L g1184 ( 
.A1(n_1066),
.A2(n_1043),
.B(n_1023),
.Y(n_1184)
);

OAI21x1_ASAP7_75t_L g1185 ( 
.A1(n_909),
.A2(n_913),
.B(n_918),
.Y(n_1185)
);

OAI21xp5_ASAP7_75t_L g1186 ( 
.A1(n_1064),
.A2(n_1073),
.B(n_1062),
.Y(n_1186)
);

CKINVDCx5p33_ASAP7_75t_R g1187 ( 
.A(n_947),
.Y(n_1187)
);

OAI21x1_ASAP7_75t_L g1188 ( 
.A1(n_909),
.A2(n_913),
.B(n_918),
.Y(n_1188)
);

NAND2xp5_ASAP7_75t_L g1189 ( 
.A(n_1061),
.B(n_1065),
.Y(n_1189)
);

INVx6_ASAP7_75t_L g1190 ( 
.A(n_917),
.Y(n_1190)
);

INVx1_ASAP7_75t_L g1191 ( 
.A(n_919),
.Y(n_1191)
);

AO31x2_ASAP7_75t_L g1192 ( 
.A1(n_1064),
.A2(n_929),
.A3(n_931),
.B(n_1066),
.Y(n_1192)
);

OAI21x1_ASAP7_75t_L g1193 ( 
.A1(n_909),
.A2(n_913),
.B(n_918),
.Y(n_1193)
);

OAI221xp5_ASAP7_75t_L g1194 ( 
.A1(n_996),
.A2(n_778),
.B1(n_779),
.B2(n_522),
.C(n_593),
.Y(n_1194)
);

INVx2_ASAP7_75t_L g1195 ( 
.A(n_1048),
.Y(n_1195)
);

NAND2xp5_ASAP7_75t_L g1196 ( 
.A(n_1061),
.B(n_1065),
.Y(n_1196)
);

OAI21x1_ASAP7_75t_L g1197 ( 
.A1(n_909),
.A2(n_913),
.B(n_918),
.Y(n_1197)
);

AND2x4_ASAP7_75t_L g1198 ( 
.A(n_915),
.B(n_1004),
.Y(n_1198)
);

NAND2xp5_ASAP7_75t_SL g1199 ( 
.A(n_954),
.B(n_800),
.Y(n_1199)
);

INVx5_ASAP7_75t_L g1200 ( 
.A(n_1069),
.Y(n_1200)
);

OAI21x1_ASAP7_75t_L g1201 ( 
.A1(n_909),
.A2(n_913),
.B(n_918),
.Y(n_1201)
);

OAI21x1_ASAP7_75t_L g1202 ( 
.A1(n_909),
.A2(n_913),
.B(n_918),
.Y(n_1202)
);

NAND2xp5_ASAP7_75t_SL g1203 ( 
.A(n_954),
.B(n_800),
.Y(n_1203)
);

INVx2_ASAP7_75t_SL g1204 ( 
.A(n_916),
.Y(n_1204)
);

OAI21x1_ASAP7_75t_L g1205 ( 
.A1(n_909),
.A2(n_913),
.B(n_918),
.Y(n_1205)
);

OAI21x1_ASAP7_75t_L g1206 ( 
.A1(n_909),
.A2(n_913),
.B(n_918),
.Y(n_1206)
);

AOI21x1_ASAP7_75t_L g1207 ( 
.A1(n_1039),
.A2(n_1044),
.B(n_958),
.Y(n_1207)
);

INVx3_ASAP7_75t_L g1208 ( 
.A(n_1069),
.Y(n_1208)
);

O2A1O1Ixp5_ASAP7_75t_L g1209 ( 
.A1(n_931),
.A2(n_1064),
.B(n_1043),
.C(n_1053),
.Y(n_1209)
);

OAI21x1_ASAP7_75t_L g1210 ( 
.A1(n_909),
.A2(n_913),
.B(n_918),
.Y(n_1210)
);

AOI21x1_ASAP7_75t_L g1211 ( 
.A1(n_1039),
.A2(n_1044),
.B(n_958),
.Y(n_1211)
);

OAI21x1_ASAP7_75t_L g1212 ( 
.A1(n_909),
.A2(n_913),
.B(n_918),
.Y(n_1212)
);

BUFx12f_ASAP7_75t_L g1213 ( 
.A(n_943),
.Y(n_1213)
);

AOI211x1_ASAP7_75t_L g1214 ( 
.A1(n_1023),
.A2(n_999),
.B(n_1033),
.C(n_929),
.Y(n_1214)
);

AND2x2_ASAP7_75t_L g1215 ( 
.A(n_954),
.B(n_779),
.Y(n_1215)
);

NAND2x1_ASAP7_75t_L g1216 ( 
.A(n_955),
.B(n_767),
.Y(n_1216)
);

INVx1_ASAP7_75t_L g1217 ( 
.A(n_919),
.Y(n_1217)
);

NAND2xp33_ASAP7_75t_L g1218 ( 
.A(n_931),
.B(n_1064),
.Y(n_1218)
);

OAI22xp5_ASAP7_75t_L g1219 ( 
.A1(n_1064),
.A2(n_931),
.B1(n_592),
.B2(n_1061),
.Y(n_1219)
);

INVx1_ASAP7_75t_L g1220 ( 
.A(n_919),
.Y(n_1220)
);

AO31x2_ASAP7_75t_L g1221 ( 
.A1(n_1064),
.A2(n_929),
.A3(n_931),
.B(n_1066),
.Y(n_1221)
);

NAND2xp5_ASAP7_75t_SL g1222 ( 
.A(n_954),
.B(n_800),
.Y(n_1222)
);

NOR2x1_ASAP7_75t_SL g1223 ( 
.A(n_1068),
.B(n_1069),
.Y(n_1223)
);

AND3x2_ASAP7_75t_L g1224 ( 
.A(n_1036),
.B(n_1020),
.C(n_819),
.Y(n_1224)
);

AND2x4_ASAP7_75t_L g1225 ( 
.A(n_1198),
.B(n_1141),
.Y(n_1225)
);

BUFx6f_ASAP7_75t_L g1226 ( 
.A(n_1156),
.Y(n_1226)
);

INVx5_ASAP7_75t_L g1227 ( 
.A(n_1091),
.Y(n_1227)
);

INVx2_ASAP7_75t_L g1228 ( 
.A(n_1084),
.Y(n_1228)
);

OAI22xp5_ASAP7_75t_L g1229 ( 
.A1(n_1080),
.A2(n_1083),
.B1(n_1178),
.B2(n_1169),
.Y(n_1229)
);

INVx2_ASAP7_75t_L g1230 ( 
.A(n_1101),
.Y(n_1230)
);

AOI22xp5_ASAP7_75t_L g1231 ( 
.A1(n_1079),
.A2(n_1194),
.B1(n_1100),
.B2(n_1176),
.Y(n_1231)
);

INVx2_ASAP7_75t_SL g1232 ( 
.A(n_1190),
.Y(n_1232)
);

INVx2_ASAP7_75t_L g1233 ( 
.A(n_1129),
.Y(n_1233)
);

INVx1_ASAP7_75t_L g1234 ( 
.A(n_1191),
.Y(n_1234)
);

HB1xp67_ASAP7_75t_L g1235 ( 
.A(n_1107),
.Y(n_1235)
);

OAI21x1_ASAP7_75t_SL g1236 ( 
.A1(n_1165),
.A2(n_1148),
.B(n_1098),
.Y(n_1236)
);

NOR2x1_ASAP7_75t_SL g1237 ( 
.A(n_1200),
.B(n_1156),
.Y(n_1237)
);

NAND2xp5_ASAP7_75t_L g1238 ( 
.A(n_1182),
.B(n_1189),
.Y(n_1238)
);

INVx3_ASAP7_75t_L g1239 ( 
.A(n_1077),
.Y(n_1239)
);

OA21x2_ASAP7_75t_L g1240 ( 
.A1(n_1125),
.A2(n_1113),
.B(n_1108),
.Y(n_1240)
);

AND2x4_ASAP7_75t_L g1241 ( 
.A(n_1198),
.B(n_1130),
.Y(n_1241)
);

AOI22xp5_ASAP7_75t_L g1242 ( 
.A1(n_1189),
.A2(n_1196),
.B1(n_1162),
.B2(n_1139),
.Y(n_1242)
);

INVx2_ASAP7_75t_L g1243 ( 
.A(n_1217),
.Y(n_1243)
);

INVx2_ASAP7_75t_L g1244 ( 
.A(n_1220),
.Y(n_1244)
);

HB1xp67_ASAP7_75t_L g1245 ( 
.A(n_1133),
.Y(n_1245)
);

NAND3xp33_ASAP7_75t_L g1246 ( 
.A(n_1167),
.B(n_1170),
.C(n_1209),
.Y(n_1246)
);

BUFx2_ASAP7_75t_L g1247 ( 
.A(n_1187),
.Y(n_1247)
);

A2O1A1Ixp33_ASAP7_75t_L g1248 ( 
.A1(n_1089),
.A2(n_1095),
.B(n_1162),
.C(n_1165),
.Y(n_1248)
);

NAND2xp5_ASAP7_75t_L g1249 ( 
.A(n_1124),
.B(n_1092),
.Y(n_1249)
);

BUFx12f_ASAP7_75t_L g1250 ( 
.A(n_1213),
.Y(n_1250)
);

CKINVDCx20_ASAP7_75t_R g1251 ( 
.A(n_1175),
.Y(n_1251)
);

BUFx12f_ASAP7_75t_L g1252 ( 
.A(n_1140),
.Y(n_1252)
);

CKINVDCx8_ASAP7_75t_R g1253 ( 
.A(n_1156),
.Y(n_1253)
);

OAI21xp5_ASAP7_75t_L g1254 ( 
.A1(n_1089),
.A2(n_1219),
.B(n_1218),
.Y(n_1254)
);

INVx1_ASAP7_75t_L g1255 ( 
.A(n_1143),
.Y(n_1255)
);

AND2x2_ASAP7_75t_L g1256 ( 
.A(n_1180),
.B(n_1215),
.Y(n_1256)
);

INVx5_ASAP7_75t_L g1257 ( 
.A(n_1091),
.Y(n_1257)
);

NAND3xp33_ASAP7_75t_L g1258 ( 
.A(n_1219),
.B(n_1149),
.C(n_1224),
.Y(n_1258)
);

NAND2xp5_ASAP7_75t_L g1259 ( 
.A(n_1092),
.B(n_1135),
.Y(n_1259)
);

AOI22xp33_ASAP7_75t_SL g1260 ( 
.A1(n_1144),
.A2(n_1136),
.B1(n_1190),
.B2(n_1172),
.Y(n_1260)
);

OR2x2_ASAP7_75t_L g1261 ( 
.A(n_1104),
.B(n_1152),
.Y(n_1261)
);

INVx2_ASAP7_75t_SL g1262 ( 
.A(n_1159),
.Y(n_1262)
);

A2O1A1Ixp33_ASAP7_75t_L g1263 ( 
.A1(n_1137),
.A2(n_1161),
.B(n_1146),
.C(n_1163),
.Y(n_1263)
);

NAND2xp5_ASAP7_75t_L g1264 ( 
.A(n_1085),
.B(n_1204),
.Y(n_1264)
);

NOR2xp33_ASAP7_75t_L g1265 ( 
.A(n_1142),
.B(n_1179),
.Y(n_1265)
);

AND2x2_ASAP7_75t_L g1266 ( 
.A(n_1115),
.B(n_1199),
.Y(n_1266)
);

AND2x2_ASAP7_75t_L g1267 ( 
.A(n_1203),
.B(n_1222),
.Y(n_1267)
);

AOI22xp5_ASAP7_75t_L g1268 ( 
.A1(n_1118),
.A2(n_1184),
.B1(n_1168),
.B2(n_1146),
.Y(n_1268)
);

AOI22xp33_ASAP7_75t_L g1269 ( 
.A1(n_1158),
.A2(n_1151),
.B1(n_1112),
.B2(n_1086),
.Y(n_1269)
);

BUFx8_ASAP7_75t_SL g1270 ( 
.A(n_1082),
.Y(n_1270)
);

BUFx12f_ASAP7_75t_L g1271 ( 
.A(n_1166),
.Y(n_1271)
);

HB1xp67_ASAP7_75t_L g1272 ( 
.A(n_1088),
.Y(n_1272)
);

INVx5_ASAP7_75t_L g1273 ( 
.A(n_1091),
.Y(n_1273)
);

AOI22xp33_ASAP7_75t_L g1274 ( 
.A1(n_1121),
.A2(n_1157),
.B1(n_1195),
.B2(n_1093),
.Y(n_1274)
);

AO21x1_ASAP7_75t_L g1275 ( 
.A1(n_1121),
.A2(n_1087),
.B(n_1096),
.Y(n_1275)
);

CKINVDCx5p33_ASAP7_75t_R g1276 ( 
.A(n_1173),
.Y(n_1276)
);

AND2x4_ASAP7_75t_L g1277 ( 
.A(n_1156),
.B(n_1099),
.Y(n_1277)
);

INVx2_ASAP7_75t_SL g1278 ( 
.A(n_1166),
.Y(n_1278)
);

AOI21xp33_ASAP7_75t_L g1279 ( 
.A1(n_1177),
.A2(n_1186),
.B(n_1109),
.Y(n_1279)
);

BUFx2_ASAP7_75t_L g1280 ( 
.A(n_1102),
.Y(n_1280)
);

OAI22xp5_ASAP7_75t_L g1281 ( 
.A1(n_1214),
.A2(n_1082),
.B1(n_1131),
.B2(n_1155),
.Y(n_1281)
);

NAND2xp5_ASAP7_75t_L g1282 ( 
.A(n_1192),
.B(n_1221),
.Y(n_1282)
);

BUFx3_ASAP7_75t_L g1283 ( 
.A(n_1102),
.Y(n_1283)
);

NAND2xp5_ASAP7_75t_L g1284 ( 
.A(n_1192),
.B(n_1221),
.Y(n_1284)
);

AOI21xp33_ASAP7_75t_L g1285 ( 
.A1(n_1177),
.A2(n_1186),
.B(n_1109),
.Y(n_1285)
);

CKINVDCx20_ASAP7_75t_R g1286 ( 
.A(n_1102),
.Y(n_1286)
);

A2O1A1Ixp33_ASAP7_75t_L g1287 ( 
.A1(n_1154),
.A2(n_1138),
.B(n_1147),
.C(n_1145),
.Y(n_1287)
);

AOI21xp5_ASAP7_75t_L g1288 ( 
.A1(n_1106),
.A2(n_1105),
.B(n_1111),
.Y(n_1288)
);

BUFx6f_ASAP7_75t_L g1289 ( 
.A(n_1181),
.Y(n_1289)
);

INVx4_ASAP7_75t_L g1290 ( 
.A(n_1200),
.Y(n_1290)
);

BUFx6f_ASAP7_75t_L g1291 ( 
.A(n_1181),
.Y(n_1291)
);

NOR2xp33_ASAP7_75t_L g1292 ( 
.A(n_1128),
.B(n_1126),
.Y(n_1292)
);

NOR2xp33_ASAP7_75t_SL g1293 ( 
.A(n_1200),
.B(n_1099),
.Y(n_1293)
);

OAI22xp5_ASAP7_75t_L g1294 ( 
.A1(n_1126),
.A2(n_1200),
.B1(n_1120),
.B2(n_1113),
.Y(n_1294)
);

NAND2xp5_ASAP7_75t_L g1295 ( 
.A(n_1192),
.B(n_1221),
.Y(n_1295)
);

OAI21xp33_ASAP7_75t_L g1296 ( 
.A1(n_1120),
.A2(n_1125),
.B(n_1108),
.Y(n_1296)
);

BUFx3_ASAP7_75t_L g1297 ( 
.A(n_1110),
.Y(n_1297)
);

OAI22xp5_ASAP7_75t_L g1298 ( 
.A1(n_1077),
.A2(n_1183),
.B1(n_1097),
.B2(n_1123),
.Y(n_1298)
);

AOI21xp33_ASAP7_75t_SL g1299 ( 
.A1(n_1153),
.A2(n_1208),
.B(n_1171),
.Y(n_1299)
);

CKINVDCx11_ASAP7_75t_R g1300 ( 
.A(n_1164),
.Y(n_1300)
);

AND2x2_ASAP7_75t_L g1301 ( 
.A(n_1164),
.B(n_1208),
.Y(n_1301)
);

AND2x2_ASAP7_75t_L g1302 ( 
.A(n_1164),
.B(n_1119),
.Y(n_1302)
);

INVx1_ASAP7_75t_SL g1303 ( 
.A(n_1216),
.Y(n_1303)
);

BUFx3_ASAP7_75t_L g1304 ( 
.A(n_1119),
.Y(n_1304)
);

INVx1_ASAP7_75t_SL g1305 ( 
.A(n_1134),
.Y(n_1305)
);

BUFx6f_ASAP7_75t_L g1306 ( 
.A(n_1132),
.Y(n_1306)
);

OR2x2_ASAP7_75t_L g1307 ( 
.A(n_1090),
.B(n_1127),
.Y(n_1307)
);

INVx4_ASAP7_75t_L g1308 ( 
.A(n_1223),
.Y(n_1308)
);

INVx2_ASAP7_75t_SL g1309 ( 
.A(n_1127),
.Y(n_1309)
);

NAND2xp5_ASAP7_75t_L g1310 ( 
.A(n_1127),
.B(n_1114),
.Y(n_1310)
);

INVx1_ASAP7_75t_L g1311 ( 
.A(n_1174),
.Y(n_1311)
);

HB1xp67_ASAP7_75t_L g1312 ( 
.A(n_1094),
.Y(n_1312)
);

CKINVDCx16_ASAP7_75t_R g1313 ( 
.A(n_1103),
.Y(n_1313)
);

INVx1_ASAP7_75t_L g1314 ( 
.A(n_1185),
.Y(n_1314)
);

CKINVDCx20_ASAP7_75t_R g1315 ( 
.A(n_1160),
.Y(n_1315)
);

AOI21xp5_ASAP7_75t_L g1316 ( 
.A1(n_1081),
.A2(n_1116),
.B(n_1117),
.Y(n_1316)
);

NAND2xp5_ASAP7_75t_L g1317 ( 
.A(n_1188),
.B(n_1205),
.Y(n_1317)
);

NAND2xp5_ASAP7_75t_L g1318 ( 
.A(n_1193),
.B(n_1202),
.Y(n_1318)
);

AOI21xp5_ASAP7_75t_L g1319 ( 
.A1(n_1150),
.A2(n_1206),
.B(n_1212),
.Y(n_1319)
);

NOR3xp33_ASAP7_75t_L g1320 ( 
.A(n_1197),
.B(n_1201),
.C(n_1210),
.Y(n_1320)
);

BUFx6f_ASAP7_75t_L g1321 ( 
.A(n_1122),
.Y(n_1321)
);

NAND2xp5_ASAP7_75t_L g1322 ( 
.A(n_1080),
.B(n_1083),
.Y(n_1322)
);

INVx2_ASAP7_75t_SL g1323 ( 
.A(n_1190),
.Y(n_1323)
);

AND2x2_ASAP7_75t_L g1324 ( 
.A(n_1139),
.B(n_1180),
.Y(n_1324)
);

AOI21xp5_ASAP7_75t_L g1325 ( 
.A1(n_1080),
.A2(n_1083),
.B(n_1078),
.Y(n_1325)
);

BUFx6f_ASAP7_75t_L g1326 ( 
.A(n_1156),
.Y(n_1326)
);

OR2x6_ASAP7_75t_L g1327 ( 
.A(n_1190),
.B(n_1213),
.Y(n_1327)
);

NAND2xp5_ASAP7_75t_L g1328 ( 
.A(n_1080),
.B(n_1083),
.Y(n_1328)
);

OAI21xp5_ASAP7_75t_L g1329 ( 
.A1(n_1209),
.A2(n_1170),
.B(n_1167),
.Y(n_1329)
);

INVx2_ASAP7_75t_L g1330 ( 
.A(n_1084),
.Y(n_1330)
);

NAND2xp5_ASAP7_75t_L g1331 ( 
.A(n_1080),
.B(n_1083),
.Y(n_1331)
);

INVx1_ASAP7_75t_L g1332 ( 
.A(n_1084),
.Y(n_1332)
);

NAND2xp5_ASAP7_75t_L g1333 ( 
.A(n_1080),
.B(n_1083),
.Y(n_1333)
);

AND2x4_ASAP7_75t_L g1334 ( 
.A(n_1198),
.B(n_915),
.Y(n_1334)
);

INVx4_ASAP7_75t_L g1335 ( 
.A(n_1156),
.Y(n_1335)
);

CKINVDCx5p33_ASAP7_75t_R g1336 ( 
.A(n_1187),
.Y(n_1336)
);

AOI22xp33_ASAP7_75t_L g1337 ( 
.A1(n_1079),
.A2(n_945),
.B1(n_1194),
.B2(n_996),
.Y(n_1337)
);

OAI22xp5_ASAP7_75t_L g1338 ( 
.A1(n_1080),
.A2(n_1083),
.B1(n_1178),
.B2(n_1169),
.Y(n_1338)
);

NAND2xp5_ASAP7_75t_L g1339 ( 
.A(n_1080),
.B(n_1083),
.Y(n_1339)
);

NAND2xp5_ASAP7_75t_L g1340 ( 
.A(n_1080),
.B(n_1083),
.Y(n_1340)
);

AND2x6_ASAP7_75t_L g1341 ( 
.A(n_1089),
.B(n_1069),
.Y(n_1341)
);

INVx5_ASAP7_75t_L g1342 ( 
.A(n_1091),
.Y(n_1342)
);

BUFx6f_ASAP7_75t_L g1343 ( 
.A(n_1156),
.Y(n_1343)
);

NOR2xp33_ASAP7_75t_SL g1344 ( 
.A(n_1144),
.B(n_1036),
.Y(n_1344)
);

AOI21xp5_ASAP7_75t_L g1345 ( 
.A1(n_1080),
.A2(n_1083),
.B(n_1078),
.Y(n_1345)
);

BUFx6f_ASAP7_75t_L g1346 ( 
.A(n_1156),
.Y(n_1346)
);

NAND2xp5_ASAP7_75t_L g1347 ( 
.A(n_1080),
.B(n_1083),
.Y(n_1347)
);

INVx3_ASAP7_75t_L g1348 ( 
.A(n_1077),
.Y(n_1348)
);

HB1xp67_ASAP7_75t_L g1349 ( 
.A(n_1107),
.Y(n_1349)
);

NAND2xp5_ASAP7_75t_SL g1350 ( 
.A(n_1100),
.B(n_1176),
.Y(n_1350)
);

O2A1O1Ixp33_ASAP7_75t_L g1351 ( 
.A1(n_1194),
.A2(n_1079),
.B(n_1100),
.C(n_1167),
.Y(n_1351)
);

AND2x4_ASAP7_75t_L g1352 ( 
.A(n_1198),
.B(n_915),
.Y(n_1352)
);

NAND2xp5_ASAP7_75t_L g1353 ( 
.A(n_1080),
.B(n_1083),
.Y(n_1353)
);

NAND2xp5_ASAP7_75t_L g1354 ( 
.A(n_1080),
.B(n_1083),
.Y(n_1354)
);

NAND2xp5_ASAP7_75t_L g1355 ( 
.A(n_1080),
.B(n_1083),
.Y(n_1355)
);

CKINVDCx5p33_ASAP7_75t_R g1356 ( 
.A(n_1187),
.Y(n_1356)
);

AND2x4_ASAP7_75t_L g1357 ( 
.A(n_1198),
.B(n_915),
.Y(n_1357)
);

NOR2xp67_ASAP7_75t_L g1358 ( 
.A(n_1187),
.B(n_888),
.Y(n_1358)
);

AOI21xp5_ASAP7_75t_L g1359 ( 
.A1(n_1080),
.A2(n_1083),
.B(n_1078),
.Y(n_1359)
);

AND2x4_ASAP7_75t_L g1360 ( 
.A(n_1198),
.B(n_915),
.Y(n_1360)
);

OAI22xp5_ASAP7_75t_L g1361 ( 
.A1(n_1080),
.A2(n_1083),
.B1(n_1178),
.B2(n_1169),
.Y(n_1361)
);

A2O1A1Ixp33_ASAP7_75t_L g1362 ( 
.A1(n_1079),
.A2(n_1167),
.B(n_1170),
.C(n_1064),
.Y(n_1362)
);

BUFx2_ASAP7_75t_R g1363 ( 
.A(n_1336),
.Y(n_1363)
);

AND2x2_ASAP7_75t_L g1364 ( 
.A(n_1242),
.B(n_1238),
.Y(n_1364)
);

BUFx2_ASAP7_75t_L g1365 ( 
.A(n_1301),
.Y(n_1365)
);

OAI21xp5_ASAP7_75t_L g1366 ( 
.A1(n_1231),
.A2(n_1351),
.B(n_1263),
.Y(n_1366)
);

INVx1_ASAP7_75t_L g1367 ( 
.A(n_1228),
.Y(n_1367)
);

INVx1_ASAP7_75t_L g1368 ( 
.A(n_1230),
.Y(n_1368)
);

AOI22xp33_ASAP7_75t_SL g1369 ( 
.A1(n_1344),
.A2(n_1313),
.B1(n_1258),
.B2(n_1246),
.Y(n_1369)
);

AO21x2_ASAP7_75t_L g1370 ( 
.A1(n_1320),
.A2(n_1319),
.B(n_1287),
.Y(n_1370)
);

AND2x4_ASAP7_75t_L g1371 ( 
.A(n_1241),
.B(n_1334),
.Y(n_1371)
);

BUFx4f_ASAP7_75t_SL g1372 ( 
.A(n_1286),
.Y(n_1372)
);

AOI22xp5_ASAP7_75t_L g1373 ( 
.A1(n_1337),
.A2(n_1231),
.B1(n_1344),
.B2(n_1350),
.Y(n_1373)
);

OR2x2_ASAP7_75t_L g1374 ( 
.A(n_1312),
.B(n_1282),
.Y(n_1374)
);

NAND2xp5_ASAP7_75t_L g1375 ( 
.A(n_1322),
.B(n_1328),
.Y(n_1375)
);

INVx1_ASAP7_75t_L g1376 ( 
.A(n_1233),
.Y(n_1376)
);

AND2x4_ASAP7_75t_L g1377 ( 
.A(n_1241),
.B(n_1334),
.Y(n_1377)
);

NAND2x1p5_ASAP7_75t_L g1378 ( 
.A(n_1304),
.B(n_1305),
.Y(n_1378)
);

AOI22xp33_ASAP7_75t_SL g1379 ( 
.A1(n_1258),
.A2(n_1246),
.B1(n_1329),
.B2(n_1315),
.Y(n_1379)
);

INVx1_ASAP7_75t_L g1380 ( 
.A(n_1243),
.Y(n_1380)
);

AND2x2_ASAP7_75t_L g1381 ( 
.A(n_1229),
.B(n_1338),
.Y(n_1381)
);

AOI22xp33_ASAP7_75t_L g1382 ( 
.A1(n_1300),
.A2(n_1329),
.B1(n_1254),
.B2(n_1265),
.Y(n_1382)
);

INVx1_ASAP7_75t_L g1383 ( 
.A(n_1244),
.Y(n_1383)
);

OR2x2_ASAP7_75t_L g1384 ( 
.A(n_1284),
.B(n_1295),
.Y(n_1384)
);

INVx1_ASAP7_75t_L g1385 ( 
.A(n_1330),
.Y(n_1385)
);

INVx1_ASAP7_75t_L g1386 ( 
.A(n_1234),
.Y(n_1386)
);

AND2x4_ASAP7_75t_L g1387 ( 
.A(n_1352),
.B(n_1357),
.Y(n_1387)
);

INVx1_ASAP7_75t_SL g1388 ( 
.A(n_1276),
.Y(n_1388)
);

INVx2_ASAP7_75t_L g1389 ( 
.A(n_1255),
.Y(n_1389)
);

INVx1_ASAP7_75t_L g1390 ( 
.A(n_1307),
.Y(n_1390)
);

OAI22xp33_ASAP7_75t_L g1391 ( 
.A1(n_1331),
.A2(n_1355),
.B1(n_1347),
.B2(n_1353),
.Y(n_1391)
);

AND2x2_ASAP7_75t_L g1392 ( 
.A(n_1338),
.B(n_1361),
.Y(n_1392)
);

AOI22xp33_ASAP7_75t_L g1393 ( 
.A1(n_1254),
.A2(n_1361),
.B1(n_1302),
.B2(n_1267),
.Y(n_1393)
);

INVx1_ASAP7_75t_L g1394 ( 
.A(n_1309),
.Y(n_1394)
);

HB1xp67_ASAP7_75t_L g1395 ( 
.A(n_1235),
.Y(n_1395)
);

AOI22xp33_ASAP7_75t_L g1396 ( 
.A1(n_1260),
.A2(n_1285),
.B1(n_1279),
.B2(n_1259),
.Y(n_1396)
);

INVx1_ASAP7_75t_L g1397 ( 
.A(n_1310),
.Y(n_1397)
);

NAND2x1p5_ASAP7_75t_L g1398 ( 
.A(n_1305),
.B(n_1240),
.Y(n_1398)
);

INVx1_ASAP7_75t_L g1399 ( 
.A(n_1311),
.Y(n_1399)
);

BUFx2_ASAP7_75t_L g1400 ( 
.A(n_1341),
.Y(n_1400)
);

BUFx3_ASAP7_75t_L g1401 ( 
.A(n_1253),
.Y(n_1401)
);

AOI21x1_ASAP7_75t_L g1402 ( 
.A1(n_1317),
.A2(n_1318),
.B(n_1316),
.Y(n_1402)
);

BUFx3_ASAP7_75t_L g1403 ( 
.A(n_1247),
.Y(n_1403)
);

INVx3_ASAP7_75t_L g1404 ( 
.A(n_1341),
.Y(n_1404)
);

AND2x2_ASAP7_75t_L g1405 ( 
.A(n_1333),
.B(n_1339),
.Y(n_1405)
);

BUFx6f_ASAP7_75t_L g1406 ( 
.A(n_1226),
.Y(n_1406)
);

AOI22xp33_ASAP7_75t_L g1407 ( 
.A1(n_1279),
.A2(n_1285),
.B1(n_1324),
.B2(n_1340),
.Y(n_1407)
);

INVx1_ASAP7_75t_L g1408 ( 
.A(n_1314),
.Y(n_1408)
);

INVx2_ASAP7_75t_L g1409 ( 
.A(n_1332),
.Y(n_1409)
);

NAND2xp5_ASAP7_75t_L g1410 ( 
.A(n_1354),
.B(n_1249),
.Y(n_1410)
);

AOI22xp33_ASAP7_75t_L g1411 ( 
.A1(n_1268),
.A2(n_1236),
.B1(n_1266),
.B2(n_1256),
.Y(n_1411)
);

OA21x2_ASAP7_75t_L g1412 ( 
.A1(n_1296),
.A2(n_1275),
.B(n_1248),
.Y(n_1412)
);

INVx1_ASAP7_75t_SL g1413 ( 
.A(n_1349),
.Y(n_1413)
);

HB1xp67_ASAP7_75t_L g1414 ( 
.A(n_1245),
.Y(n_1414)
);

BUFx3_ASAP7_75t_L g1415 ( 
.A(n_1225),
.Y(n_1415)
);

NAND2xp5_ASAP7_75t_L g1416 ( 
.A(n_1261),
.B(n_1362),
.Y(n_1416)
);

CKINVDCx11_ASAP7_75t_R g1417 ( 
.A(n_1250),
.Y(n_1417)
);

HB1xp67_ASAP7_75t_L g1418 ( 
.A(n_1272),
.Y(n_1418)
);

HB1xp67_ASAP7_75t_L g1419 ( 
.A(n_1262),
.Y(n_1419)
);

AND2x2_ASAP7_75t_L g1420 ( 
.A(n_1292),
.B(n_1268),
.Y(n_1420)
);

INVx1_ASAP7_75t_L g1421 ( 
.A(n_1264),
.Y(n_1421)
);

OA21x2_ASAP7_75t_L g1422 ( 
.A1(n_1296),
.A2(n_1269),
.B(n_1359),
.Y(n_1422)
);

HB1xp67_ASAP7_75t_L g1423 ( 
.A(n_1225),
.Y(n_1423)
);

INVx3_ASAP7_75t_L g1424 ( 
.A(n_1341),
.Y(n_1424)
);

INVx1_ASAP7_75t_L g1425 ( 
.A(n_1294),
.Y(n_1425)
);

INVx3_ASAP7_75t_L g1426 ( 
.A(n_1341),
.Y(n_1426)
);

INVx5_ASAP7_75t_L g1427 ( 
.A(n_1326),
.Y(n_1427)
);

AO22x1_ASAP7_75t_L g1428 ( 
.A1(n_1278),
.A2(n_1281),
.B1(n_1308),
.B2(n_1303),
.Y(n_1428)
);

BUFx2_ASAP7_75t_L g1429 ( 
.A(n_1281),
.Y(n_1429)
);

CKINVDCx20_ASAP7_75t_R g1430 ( 
.A(n_1270),
.Y(n_1430)
);

INVx1_ASAP7_75t_SL g1431 ( 
.A(n_1356),
.Y(n_1431)
);

INVx8_ASAP7_75t_L g1432 ( 
.A(n_1227),
.Y(n_1432)
);

INVx1_ASAP7_75t_L g1433 ( 
.A(n_1289),
.Y(n_1433)
);

INVx2_ASAP7_75t_SL g1434 ( 
.A(n_1227),
.Y(n_1434)
);

INVx1_ASAP7_75t_L g1435 ( 
.A(n_1289),
.Y(n_1435)
);

INVx1_ASAP7_75t_L g1436 ( 
.A(n_1291),
.Y(n_1436)
);

INVx1_ASAP7_75t_L g1437 ( 
.A(n_1294),
.Y(n_1437)
);

HB1xp67_ASAP7_75t_L g1438 ( 
.A(n_1352),
.Y(n_1438)
);

AOI22xp33_ASAP7_75t_L g1439 ( 
.A1(n_1357),
.A2(n_1360),
.B1(n_1252),
.B2(n_1251),
.Y(n_1439)
);

OAI22xp33_ASAP7_75t_L g1440 ( 
.A1(n_1358),
.A2(n_1327),
.B1(n_1293),
.B2(n_1323),
.Y(n_1440)
);

INVx1_ASAP7_75t_L g1441 ( 
.A(n_1291),
.Y(n_1441)
);

CKINVDCx12_ASAP7_75t_R g1442 ( 
.A(n_1327),
.Y(n_1442)
);

INVx1_ASAP7_75t_L g1443 ( 
.A(n_1306),
.Y(n_1443)
);

AND2x2_ASAP7_75t_L g1444 ( 
.A(n_1274),
.B(n_1345),
.Y(n_1444)
);

INVx1_ASAP7_75t_L g1445 ( 
.A(n_1306),
.Y(n_1445)
);

INVx1_ASAP7_75t_L g1446 ( 
.A(n_1299),
.Y(n_1446)
);

BUFx8_ASAP7_75t_SL g1447 ( 
.A(n_1327),
.Y(n_1447)
);

INVx2_ASAP7_75t_SL g1448 ( 
.A(n_1227),
.Y(n_1448)
);

BUFx4f_ASAP7_75t_SL g1449 ( 
.A(n_1271),
.Y(n_1449)
);

AOI22xp33_ASAP7_75t_L g1450 ( 
.A1(n_1325),
.A2(n_1232),
.B1(n_1298),
.B2(n_1239),
.Y(n_1450)
);

OAI21x1_ASAP7_75t_L g1451 ( 
.A1(n_1298),
.A2(n_1348),
.B(n_1239),
.Y(n_1451)
);

AND2x2_ASAP7_75t_L g1452 ( 
.A(n_1348),
.B(n_1280),
.Y(n_1452)
);

OA21x2_ASAP7_75t_L g1453 ( 
.A1(n_1321),
.A2(n_1303),
.B(n_1277),
.Y(n_1453)
);

AND2x2_ASAP7_75t_L g1454 ( 
.A(n_1308),
.B(n_1277),
.Y(n_1454)
);

BUFx2_ASAP7_75t_L g1455 ( 
.A(n_1291),
.Y(n_1455)
);

AOI222xp33_ASAP7_75t_L g1456 ( 
.A1(n_1297),
.A2(n_1293),
.B1(n_1283),
.B2(n_1237),
.C1(n_1335),
.C2(n_1346),
.Y(n_1456)
);

AOI22xp33_ASAP7_75t_L g1457 ( 
.A1(n_1321),
.A2(n_1346),
.B1(n_1326),
.B2(n_1343),
.Y(n_1457)
);

BUFx6f_ASAP7_75t_L g1458 ( 
.A(n_1326),
.Y(n_1458)
);

AOI22xp33_ASAP7_75t_L g1459 ( 
.A1(n_1343),
.A2(n_1346),
.B1(n_1290),
.B2(n_1273),
.Y(n_1459)
);

AOI22xp33_ASAP7_75t_L g1460 ( 
.A1(n_1290),
.A2(n_1257),
.B1(n_1273),
.B2(n_1342),
.Y(n_1460)
);

INVx2_ASAP7_75t_L g1461 ( 
.A(n_1342),
.Y(n_1461)
);

AND2x2_ASAP7_75t_L g1462 ( 
.A(n_1257),
.B(n_1273),
.Y(n_1462)
);

AO21x2_ASAP7_75t_L g1463 ( 
.A1(n_1257),
.A2(n_1320),
.B(n_1319),
.Y(n_1463)
);

INVx2_ASAP7_75t_L g1464 ( 
.A(n_1342),
.Y(n_1464)
);

OR2x2_ASAP7_75t_L g1465 ( 
.A(n_1313),
.B(n_1312),
.Y(n_1465)
);

OR2x2_ASAP7_75t_L g1466 ( 
.A(n_1313),
.B(n_1312),
.Y(n_1466)
);

INVx1_ASAP7_75t_L g1467 ( 
.A(n_1228),
.Y(n_1467)
);

OAI22xp33_ASAP7_75t_R g1468 ( 
.A1(n_1261),
.A2(n_1100),
.B1(n_1176),
.B2(n_413),
.Y(n_1468)
);

CKINVDCx11_ASAP7_75t_R g1469 ( 
.A(n_1286),
.Y(n_1469)
);

BUFx3_ASAP7_75t_L g1470 ( 
.A(n_1286),
.Y(n_1470)
);

CKINVDCx5p33_ASAP7_75t_R g1471 ( 
.A(n_1336),
.Y(n_1471)
);

BUFx2_ASAP7_75t_L g1472 ( 
.A(n_1301),
.Y(n_1472)
);

HB1xp67_ASAP7_75t_L g1473 ( 
.A(n_1235),
.Y(n_1473)
);

BUFx3_ASAP7_75t_L g1474 ( 
.A(n_1286),
.Y(n_1474)
);

AO21x1_ASAP7_75t_L g1475 ( 
.A1(n_1351),
.A2(n_1219),
.B(n_1218),
.Y(n_1475)
);

OAI22xp5_ASAP7_75t_L g1476 ( 
.A1(n_1322),
.A2(n_1100),
.B1(n_1331),
.B2(n_1328),
.Y(n_1476)
);

OA21x2_ASAP7_75t_L g1477 ( 
.A1(n_1288),
.A2(n_1319),
.B(n_1186),
.Y(n_1477)
);

CKINVDCx11_ASAP7_75t_R g1478 ( 
.A(n_1286),
.Y(n_1478)
);

BUFx2_ASAP7_75t_L g1479 ( 
.A(n_1301),
.Y(n_1479)
);

OAI22xp33_ASAP7_75t_L g1480 ( 
.A1(n_1344),
.A2(n_1231),
.B1(n_1194),
.B2(n_819),
.Y(n_1480)
);

BUFx3_ASAP7_75t_L g1481 ( 
.A(n_1286),
.Y(n_1481)
);

AOI21x1_ASAP7_75t_L g1482 ( 
.A1(n_1319),
.A2(n_1211),
.B(n_1207),
.Y(n_1482)
);

AOI22xp33_ASAP7_75t_SL g1483 ( 
.A1(n_1344),
.A2(n_819),
.B1(n_1100),
.B2(n_1036),
.Y(n_1483)
);

INVx1_ASAP7_75t_L g1484 ( 
.A(n_1228),
.Y(n_1484)
);

INVx1_ASAP7_75t_L g1485 ( 
.A(n_1228),
.Y(n_1485)
);

INVx3_ASAP7_75t_L g1486 ( 
.A(n_1341),
.Y(n_1486)
);

HB1xp67_ASAP7_75t_SL g1487 ( 
.A(n_1363),
.Y(n_1487)
);

NAND3xp33_ASAP7_75t_L g1488 ( 
.A(n_1483),
.B(n_1373),
.C(n_1366),
.Y(n_1488)
);

HB1xp67_ASAP7_75t_L g1489 ( 
.A(n_1418),
.Y(n_1489)
);

AOI21x1_ASAP7_75t_L g1490 ( 
.A1(n_1482),
.A2(n_1428),
.B(n_1402),
.Y(n_1490)
);

AND2x4_ASAP7_75t_L g1491 ( 
.A(n_1451),
.B(n_1443),
.Y(n_1491)
);

HB1xp67_ASAP7_75t_L g1492 ( 
.A(n_1414),
.Y(n_1492)
);

HB1xp67_ASAP7_75t_L g1493 ( 
.A(n_1395),
.Y(n_1493)
);

INVx2_ASAP7_75t_SL g1494 ( 
.A(n_1453),
.Y(n_1494)
);

BUFx3_ASAP7_75t_L g1495 ( 
.A(n_1400),
.Y(n_1495)
);

HB1xp67_ASAP7_75t_L g1496 ( 
.A(n_1473),
.Y(n_1496)
);

AND2x2_ASAP7_75t_L g1497 ( 
.A(n_1381),
.B(n_1392),
.Y(n_1497)
);

HB1xp67_ASAP7_75t_L g1498 ( 
.A(n_1465),
.Y(n_1498)
);

NAND2x1p5_ASAP7_75t_L g1499 ( 
.A(n_1451),
.B(n_1400),
.Y(n_1499)
);

AND2x2_ASAP7_75t_L g1500 ( 
.A(n_1381),
.B(n_1392),
.Y(n_1500)
);

HB1xp67_ASAP7_75t_L g1501 ( 
.A(n_1465),
.Y(n_1501)
);

INVx2_ASAP7_75t_SL g1502 ( 
.A(n_1453),
.Y(n_1502)
);

AND2x4_ASAP7_75t_L g1503 ( 
.A(n_1443),
.B(n_1445),
.Y(n_1503)
);

NAND2xp5_ASAP7_75t_L g1504 ( 
.A(n_1405),
.B(n_1476),
.Y(n_1504)
);

BUFx2_ASAP7_75t_L g1505 ( 
.A(n_1378),
.Y(n_1505)
);

BUFx2_ASAP7_75t_L g1506 ( 
.A(n_1378),
.Y(n_1506)
);

HB1xp67_ASAP7_75t_L g1507 ( 
.A(n_1466),
.Y(n_1507)
);

AND2x2_ASAP7_75t_L g1508 ( 
.A(n_1365),
.B(n_1472),
.Y(n_1508)
);

INVx1_ASAP7_75t_L g1509 ( 
.A(n_1399),
.Y(n_1509)
);

BUFx2_ASAP7_75t_L g1510 ( 
.A(n_1378),
.Y(n_1510)
);

AOI21x1_ASAP7_75t_L g1511 ( 
.A1(n_1428),
.A2(n_1446),
.B(n_1444),
.Y(n_1511)
);

INVx2_ASAP7_75t_SL g1512 ( 
.A(n_1453),
.Y(n_1512)
);

INVx1_ASAP7_75t_L g1513 ( 
.A(n_1408),
.Y(n_1513)
);

HB1xp67_ASAP7_75t_L g1514 ( 
.A(n_1466),
.Y(n_1514)
);

OR2x2_ASAP7_75t_L g1515 ( 
.A(n_1374),
.B(n_1397),
.Y(n_1515)
);

INVx2_ASAP7_75t_SL g1516 ( 
.A(n_1453),
.Y(n_1516)
);

NOR2x1_ASAP7_75t_L g1517 ( 
.A(n_1391),
.B(n_1446),
.Y(n_1517)
);

NAND2xp5_ASAP7_75t_L g1518 ( 
.A(n_1405),
.B(n_1375),
.Y(n_1518)
);

OA21x2_ASAP7_75t_L g1519 ( 
.A1(n_1429),
.A2(n_1425),
.B(n_1437),
.Y(n_1519)
);

HB1xp67_ASAP7_75t_L g1520 ( 
.A(n_1413),
.Y(n_1520)
);

OR2x6_ASAP7_75t_L g1521 ( 
.A(n_1398),
.B(n_1444),
.Y(n_1521)
);

AND2x2_ASAP7_75t_L g1522 ( 
.A(n_1365),
.B(n_1472),
.Y(n_1522)
);

OR2x6_ASAP7_75t_L g1523 ( 
.A(n_1398),
.B(n_1429),
.Y(n_1523)
);

INVx1_ASAP7_75t_L g1524 ( 
.A(n_1390),
.Y(n_1524)
);

BUFx2_ASAP7_75t_L g1525 ( 
.A(n_1479),
.Y(n_1525)
);

INVx1_ASAP7_75t_L g1526 ( 
.A(n_1390),
.Y(n_1526)
);

INVx1_ASAP7_75t_L g1527 ( 
.A(n_1394),
.Y(n_1527)
);

BUFx2_ASAP7_75t_L g1528 ( 
.A(n_1479),
.Y(n_1528)
);

AO21x1_ASAP7_75t_L g1529 ( 
.A1(n_1480),
.A2(n_1420),
.B(n_1437),
.Y(n_1529)
);

NAND2xp5_ASAP7_75t_L g1530 ( 
.A(n_1410),
.B(n_1421),
.Y(n_1530)
);

BUFx2_ASAP7_75t_L g1531 ( 
.A(n_1398),
.Y(n_1531)
);

NAND2xp5_ASAP7_75t_L g1532 ( 
.A(n_1416),
.B(n_1407),
.Y(n_1532)
);

INVx1_ASAP7_75t_L g1533 ( 
.A(n_1374),
.Y(n_1533)
);

OR2x6_ASAP7_75t_L g1534 ( 
.A(n_1475),
.B(n_1422),
.Y(n_1534)
);

INVx1_ASAP7_75t_L g1535 ( 
.A(n_1384),
.Y(n_1535)
);

AO21x2_ASAP7_75t_L g1536 ( 
.A1(n_1370),
.A2(n_1463),
.B(n_1475),
.Y(n_1536)
);

INVx1_ASAP7_75t_L g1537 ( 
.A(n_1384),
.Y(n_1537)
);

AND2x2_ASAP7_75t_L g1538 ( 
.A(n_1420),
.B(n_1364),
.Y(n_1538)
);

AND2x2_ASAP7_75t_L g1539 ( 
.A(n_1364),
.B(n_1393),
.Y(n_1539)
);

INVx5_ASAP7_75t_L g1540 ( 
.A(n_1404),
.Y(n_1540)
);

HB1xp67_ASAP7_75t_L g1541 ( 
.A(n_1389),
.Y(n_1541)
);

OR2x2_ASAP7_75t_L g1542 ( 
.A(n_1412),
.B(n_1411),
.Y(n_1542)
);

AND2x2_ASAP7_75t_L g1543 ( 
.A(n_1412),
.B(n_1409),
.Y(n_1543)
);

INVx1_ASAP7_75t_L g1544 ( 
.A(n_1412),
.Y(n_1544)
);

CKINVDCx5p33_ASAP7_75t_R g1545 ( 
.A(n_1471),
.Y(n_1545)
);

INVx3_ASAP7_75t_L g1546 ( 
.A(n_1404),
.Y(n_1546)
);

INVx1_ASAP7_75t_L g1547 ( 
.A(n_1386),
.Y(n_1547)
);

BUFx3_ASAP7_75t_L g1548 ( 
.A(n_1403),
.Y(n_1548)
);

INVx1_ASAP7_75t_L g1549 ( 
.A(n_1422),
.Y(n_1549)
);

INVx3_ASAP7_75t_L g1550 ( 
.A(n_1424),
.Y(n_1550)
);

CKINVDCx5p33_ASAP7_75t_R g1551 ( 
.A(n_1471),
.Y(n_1551)
);

INVx3_ASAP7_75t_L g1552 ( 
.A(n_1424),
.Y(n_1552)
);

AOI22xp33_ASAP7_75t_L g1553 ( 
.A1(n_1379),
.A2(n_1468),
.B1(n_1369),
.B2(n_1382),
.Y(n_1553)
);

INVx2_ASAP7_75t_L g1554 ( 
.A(n_1367),
.Y(n_1554)
);

AOI222xp33_ASAP7_75t_L g1555 ( 
.A1(n_1468),
.A2(n_1396),
.B1(n_1439),
.B2(n_1372),
.C1(n_1440),
.C2(n_1388),
.Y(n_1555)
);

AND2x2_ASAP7_75t_L g1556 ( 
.A(n_1368),
.B(n_1385),
.Y(n_1556)
);

INVx3_ASAP7_75t_L g1557 ( 
.A(n_1426),
.Y(n_1557)
);

AND2x2_ASAP7_75t_L g1558 ( 
.A(n_1376),
.B(n_1467),
.Y(n_1558)
);

INVx2_ASAP7_75t_L g1559 ( 
.A(n_1380),
.Y(n_1559)
);

AND2x2_ASAP7_75t_L g1560 ( 
.A(n_1383),
.B(n_1485),
.Y(n_1560)
);

OAI21xp5_ASAP7_75t_L g1561 ( 
.A1(n_1450),
.A2(n_1419),
.B(n_1484),
.Y(n_1561)
);

HB1xp67_ASAP7_75t_L g1562 ( 
.A(n_1498),
.Y(n_1562)
);

OR2x2_ASAP7_75t_L g1563 ( 
.A(n_1521),
.B(n_1477),
.Y(n_1563)
);

AND2x4_ASAP7_75t_L g1564 ( 
.A(n_1491),
.B(n_1486),
.Y(n_1564)
);

AND2x2_ASAP7_75t_L g1565 ( 
.A(n_1538),
.B(n_1477),
.Y(n_1565)
);

AND2x4_ASAP7_75t_L g1566 ( 
.A(n_1491),
.B(n_1486),
.Y(n_1566)
);

AND2x4_ASAP7_75t_L g1567 ( 
.A(n_1491),
.B(n_1486),
.Y(n_1567)
);

NAND2xp5_ASAP7_75t_L g1568 ( 
.A(n_1518),
.B(n_1452),
.Y(n_1568)
);

INVx2_ASAP7_75t_L g1569 ( 
.A(n_1509),
.Y(n_1569)
);

HB1xp67_ASAP7_75t_L g1570 ( 
.A(n_1501),
.Y(n_1570)
);

INVx2_ASAP7_75t_L g1571 ( 
.A(n_1513),
.Y(n_1571)
);

BUFx2_ASAP7_75t_L g1572 ( 
.A(n_1505),
.Y(n_1572)
);

OAI22xp5_ASAP7_75t_L g1573 ( 
.A1(n_1553),
.A2(n_1401),
.B1(n_1459),
.B2(n_1457),
.Y(n_1573)
);

OAI222xp33_ASAP7_75t_L g1574 ( 
.A1(n_1532),
.A2(n_1438),
.B1(n_1423),
.B2(n_1452),
.C1(n_1371),
.C2(n_1377),
.Y(n_1574)
);

OR2x2_ASAP7_75t_L g1575 ( 
.A(n_1521),
.B(n_1533),
.Y(n_1575)
);

BUFx2_ASAP7_75t_L g1576 ( 
.A(n_1505),
.Y(n_1576)
);

BUFx2_ASAP7_75t_L g1577 ( 
.A(n_1506),
.Y(n_1577)
);

AND2x2_ASAP7_75t_L g1578 ( 
.A(n_1535),
.B(n_1371),
.Y(n_1578)
);

AND2x2_ASAP7_75t_L g1579 ( 
.A(n_1537),
.B(n_1371),
.Y(n_1579)
);

AND2x4_ASAP7_75t_L g1580 ( 
.A(n_1521),
.B(n_1454),
.Y(n_1580)
);

HB1xp67_ASAP7_75t_L g1581 ( 
.A(n_1507),
.Y(n_1581)
);

NAND2xp5_ASAP7_75t_L g1582 ( 
.A(n_1504),
.B(n_1481),
.Y(n_1582)
);

AOI222xp33_ASAP7_75t_L g1583 ( 
.A1(n_1488),
.A2(n_1417),
.B1(n_1470),
.B2(n_1481),
.C1(n_1474),
.C2(n_1478),
.Y(n_1583)
);

INVxp33_ASAP7_75t_L g1584 ( 
.A(n_1520),
.Y(n_1584)
);

INVx2_ASAP7_75t_L g1585 ( 
.A(n_1543),
.Y(n_1585)
);

NAND2xp5_ASAP7_75t_L g1586 ( 
.A(n_1514),
.B(n_1474),
.Y(n_1586)
);

INVx1_ASAP7_75t_SL g1587 ( 
.A(n_1525),
.Y(n_1587)
);

BUFx2_ASAP7_75t_L g1588 ( 
.A(n_1510),
.Y(n_1588)
);

AOI22xp33_ASAP7_75t_L g1589 ( 
.A1(n_1529),
.A2(n_1377),
.B1(n_1470),
.B2(n_1387),
.Y(n_1589)
);

NAND2xp5_ASAP7_75t_L g1590 ( 
.A(n_1530),
.B(n_1415),
.Y(n_1590)
);

AOI211xp5_ASAP7_75t_L g1591 ( 
.A1(n_1529),
.A2(n_1431),
.B(n_1387),
.C(n_1401),
.Y(n_1591)
);

NAND2xp5_ASAP7_75t_L g1592 ( 
.A(n_1489),
.B(n_1492),
.Y(n_1592)
);

NAND2xp5_ASAP7_75t_L g1593 ( 
.A(n_1493),
.B(n_1415),
.Y(n_1593)
);

BUFx6f_ASAP7_75t_L g1594 ( 
.A(n_1499),
.Y(n_1594)
);

AND2x2_ASAP7_75t_L g1595 ( 
.A(n_1521),
.B(n_1433),
.Y(n_1595)
);

AND2x2_ASAP7_75t_L g1596 ( 
.A(n_1521),
.B(n_1436),
.Y(n_1596)
);

AND2x4_ASAP7_75t_L g1597 ( 
.A(n_1503),
.B(n_1454),
.Y(n_1597)
);

NAND2xp5_ASAP7_75t_L g1598 ( 
.A(n_1496),
.B(n_1455),
.Y(n_1598)
);

NOR2xp33_ASAP7_75t_SL g1599 ( 
.A(n_1517),
.B(n_1447),
.Y(n_1599)
);

BUFx2_ASAP7_75t_L g1600 ( 
.A(n_1531),
.Y(n_1600)
);

AND2x2_ASAP7_75t_L g1601 ( 
.A(n_1508),
.B(n_1441),
.Y(n_1601)
);

AND2x2_ASAP7_75t_L g1602 ( 
.A(n_1508),
.B(n_1435),
.Y(n_1602)
);

INVx2_ASAP7_75t_L g1603 ( 
.A(n_1544),
.Y(n_1603)
);

NAND3xp33_ASAP7_75t_L g1604 ( 
.A(n_1517),
.B(n_1456),
.C(n_1469),
.Y(n_1604)
);

AND2x2_ASAP7_75t_L g1605 ( 
.A(n_1522),
.B(n_1461),
.Y(n_1605)
);

INVx1_ASAP7_75t_L g1606 ( 
.A(n_1527),
.Y(n_1606)
);

INVx4_ASAP7_75t_L g1607 ( 
.A(n_1540),
.Y(n_1607)
);

AND2x2_ASAP7_75t_L g1608 ( 
.A(n_1522),
.B(n_1461),
.Y(n_1608)
);

INVx1_ASAP7_75t_L g1609 ( 
.A(n_1527),
.Y(n_1609)
);

AOI21xp33_ASAP7_75t_SL g1610 ( 
.A1(n_1583),
.A2(n_1555),
.B(n_1545),
.Y(n_1610)
);

NOR2xp33_ASAP7_75t_L g1611 ( 
.A(n_1584),
.B(n_1548),
.Y(n_1611)
);

AOI22xp33_ASAP7_75t_L g1612 ( 
.A1(n_1604),
.A2(n_1539),
.B1(n_1523),
.B2(n_1542),
.Y(n_1612)
);

NAND2xp5_ASAP7_75t_L g1613 ( 
.A(n_1562),
.B(n_1539),
.Y(n_1613)
);

NAND2xp5_ASAP7_75t_L g1614 ( 
.A(n_1587),
.B(n_1519),
.Y(n_1614)
);

NAND2xp5_ASAP7_75t_L g1615 ( 
.A(n_1587),
.B(n_1519),
.Y(n_1615)
);

AND2x2_ASAP7_75t_L g1616 ( 
.A(n_1565),
.B(n_1523),
.Y(n_1616)
);

NAND2xp5_ASAP7_75t_L g1617 ( 
.A(n_1570),
.B(n_1519),
.Y(n_1617)
);

NAND2xp5_ASAP7_75t_L g1618 ( 
.A(n_1581),
.B(n_1592),
.Y(n_1618)
);

NAND2xp5_ASAP7_75t_L g1619 ( 
.A(n_1606),
.B(n_1519),
.Y(n_1619)
);

AND2x2_ASAP7_75t_L g1620 ( 
.A(n_1565),
.B(n_1523),
.Y(n_1620)
);

NAND2xp5_ASAP7_75t_L g1621 ( 
.A(n_1606),
.B(n_1515),
.Y(n_1621)
);

NAND2xp5_ASAP7_75t_L g1622 ( 
.A(n_1609),
.B(n_1515),
.Y(n_1622)
);

NAND2xp5_ASAP7_75t_L g1623 ( 
.A(n_1609),
.B(n_1524),
.Y(n_1623)
);

NAND2xp5_ASAP7_75t_L g1624 ( 
.A(n_1569),
.B(n_1524),
.Y(n_1624)
);

NAND2xp5_ASAP7_75t_SL g1625 ( 
.A(n_1599),
.B(n_1561),
.Y(n_1625)
);

NAND2xp5_ASAP7_75t_L g1626 ( 
.A(n_1569),
.B(n_1526),
.Y(n_1626)
);

OAI221xp5_ASAP7_75t_SL g1627 ( 
.A1(n_1591),
.A2(n_1542),
.B1(n_1534),
.B2(n_1525),
.C(n_1528),
.Y(n_1627)
);

INVx1_ASAP7_75t_L g1628 ( 
.A(n_1569),
.Y(n_1628)
);

NAND2xp5_ASAP7_75t_L g1629 ( 
.A(n_1571),
.B(n_1526),
.Y(n_1629)
);

NAND3xp33_ASAP7_75t_L g1630 ( 
.A(n_1599),
.B(n_1559),
.C(n_1554),
.Y(n_1630)
);

AOI22xp33_ASAP7_75t_L g1631 ( 
.A1(n_1604),
.A2(n_1528),
.B1(n_1495),
.B2(n_1478),
.Y(n_1631)
);

NAND4xp25_ASAP7_75t_L g1632 ( 
.A(n_1583),
.B(n_1560),
.C(n_1558),
.D(n_1556),
.Y(n_1632)
);

AND2x2_ASAP7_75t_L g1633 ( 
.A(n_1585),
.B(n_1494),
.Y(n_1633)
);

OAI21xp5_ASAP7_75t_SL g1634 ( 
.A1(n_1589),
.A2(n_1511),
.B(n_1497),
.Y(n_1634)
);

AND2x2_ASAP7_75t_L g1635 ( 
.A(n_1575),
.B(n_1595),
.Y(n_1635)
);

AND2x2_ASAP7_75t_L g1636 ( 
.A(n_1595),
.B(n_1502),
.Y(n_1636)
);

NAND4xp25_ASAP7_75t_L g1637 ( 
.A(n_1591),
.B(n_1560),
.C(n_1558),
.D(n_1556),
.Y(n_1637)
);

AND2x2_ASAP7_75t_L g1638 ( 
.A(n_1596),
.B(n_1512),
.Y(n_1638)
);

AND2x2_ASAP7_75t_L g1639 ( 
.A(n_1596),
.B(n_1605),
.Y(n_1639)
);

AOI22xp33_ASAP7_75t_L g1640 ( 
.A1(n_1573),
.A2(n_1495),
.B1(n_1469),
.B2(n_1447),
.Y(n_1640)
);

AOI22xp33_ASAP7_75t_L g1641 ( 
.A1(n_1582),
.A2(n_1495),
.B1(n_1497),
.B2(n_1500),
.Y(n_1641)
);

AND2x2_ASAP7_75t_L g1642 ( 
.A(n_1605),
.B(n_1512),
.Y(n_1642)
);

NAND3xp33_ASAP7_75t_L g1643 ( 
.A(n_1586),
.B(n_1598),
.C(n_1590),
.Y(n_1643)
);

OAI21xp5_ASAP7_75t_SL g1644 ( 
.A1(n_1574),
.A2(n_1511),
.B(n_1500),
.Y(n_1644)
);

AND2x2_ASAP7_75t_L g1645 ( 
.A(n_1608),
.B(n_1516),
.Y(n_1645)
);

AND2x2_ASAP7_75t_L g1646 ( 
.A(n_1608),
.B(n_1516),
.Y(n_1646)
);

AND2x2_ASAP7_75t_L g1647 ( 
.A(n_1600),
.B(n_1534),
.Y(n_1647)
);

OAI21xp5_ASAP7_75t_SL g1648 ( 
.A1(n_1580),
.A2(n_1487),
.B(n_1499),
.Y(n_1648)
);

AND2x2_ASAP7_75t_L g1649 ( 
.A(n_1564),
.B(n_1534),
.Y(n_1649)
);

NAND2xp5_ASAP7_75t_L g1650 ( 
.A(n_1568),
.B(n_1541),
.Y(n_1650)
);

AND2x2_ASAP7_75t_L g1651 ( 
.A(n_1564),
.B(n_1534),
.Y(n_1651)
);

AOI22xp33_ASAP7_75t_L g1652 ( 
.A1(n_1580),
.A2(n_1417),
.B1(n_1552),
.B2(n_1557),
.Y(n_1652)
);

AND2x2_ASAP7_75t_L g1653 ( 
.A(n_1564),
.B(n_1536),
.Y(n_1653)
);

AND2x2_ASAP7_75t_L g1654 ( 
.A(n_1564),
.B(n_1536),
.Y(n_1654)
);

NAND2xp5_ASAP7_75t_L g1655 ( 
.A(n_1578),
.B(n_1547),
.Y(n_1655)
);

NAND2xp5_ASAP7_75t_SL g1656 ( 
.A(n_1580),
.B(n_1551),
.Y(n_1656)
);

AND2x2_ASAP7_75t_L g1657 ( 
.A(n_1566),
.B(n_1567),
.Y(n_1657)
);

AOI22xp33_ASAP7_75t_L g1658 ( 
.A1(n_1580),
.A2(n_1550),
.B1(n_1546),
.B2(n_1557),
.Y(n_1658)
);

AND2x2_ASAP7_75t_SL g1659 ( 
.A(n_1607),
.B(n_1549),
.Y(n_1659)
);

AND2x4_ASAP7_75t_SL g1660 ( 
.A(n_1657),
.B(n_1607),
.Y(n_1660)
);

OR2x2_ASAP7_75t_L g1661 ( 
.A(n_1617),
.B(n_1572),
.Y(n_1661)
);

INVx2_ASAP7_75t_L g1662 ( 
.A(n_1628),
.Y(n_1662)
);

INVx1_ASAP7_75t_L g1663 ( 
.A(n_1628),
.Y(n_1663)
);

BUFx2_ASAP7_75t_L g1664 ( 
.A(n_1659),
.Y(n_1664)
);

OR2x2_ASAP7_75t_L g1665 ( 
.A(n_1617),
.B(n_1576),
.Y(n_1665)
);

NAND2xp5_ASAP7_75t_L g1666 ( 
.A(n_1643),
.B(n_1601),
.Y(n_1666)
);

AND2x2_ASAP7_75t_L g1667 ( 
.A(n_1635),
.B(n_1576),
.Y(n_1667)
);

INVx1_ASAP7_75t_L g1668 ( 
.A(n_1624),
.Y(n_1668)
);

NAND2xp5_ASAP7_75t_L g1669 ( 
.A(n_1643),
.B(n_1618),
.Y(n_1669)
);

BUFx2_ASAP7_75t_L g1670 ( 
.A(n_1659),
.Y(n_1670)
);

NAND2x1_ASAP7_75t_L g1671 ( 
.A(n_1614),
.B(n_1607),
.Y(n_1671)
);

INVx1_ASAP7_75t_L g1672 ( 
.A(n_1624),
.Y(n_1672)
);

INVx1_ASAP7_75t_L g1673 ( 
.A(n_1626),
.Y(n_1673)
);

NAND2xp5_ASAP7_75t_L g1674 ( 
.A(n_1613),
.B(n_1601),
.Y(n_1674)
);

OR2x2_ASAP7_75t_L g1675 ( 
.A(n_1614),
.B(n_1577),
.Y(n_1675)
);

OR2x2_ASAP7_75t_L g1676 ( 
.A(n_1615),
.B(n_1588),
.Y(n_1676)
);

INVx1_ASAP7_75t_L g1677 ( 
.A(n_1626),
.Y(n_1677)
);

INVx1_ASAP7_75t_L g1678 ( 
.A(n_1629),
.Y(n_1678)
);

NAND2xp5_ASAP7_75t_L g1679 ( 
.A(n_1650),
.B(n_1602),
.Y(n_1679)
);

HB1xp67_ASAP7_75t_L g1680 ( 
.A(n_1615),
.Y(n_1680)
);

AND2x2_ASAP7_75t_L g1681 ( 
.A(n_1639),
.B(n_1566),
.Y(n_1681)
);

NAND2xp5_ASAP7_75t_L g1682 ( 
.A(n_1655),
.B(n_1579),
.Y(n_1682)
);

BUFx2_ASAP7_75t_SL g1683 ( 
.A(n_1656),
.Y(n_1683)
);

OR2x2_ASAP7_75t_L g1684 ( 
.A(n_1633),
.B(n_1563),
.Y(n_1684)
);

AND2x2_ASAP7_75t_L g1685 ( 
.A(n_1649),
.B(n_1566),
.Y(n_1685)
);

OR2x2_ASAP7_75t_L g1686 ( 
.A(n_1619),
.B(n_1563),
.Y(n_1686)
);

NAND2xp5_ASAP7_75t_L g1687 ( 
.A(n_1621),
.B(n_1622),
.Y(n_1687)
);

INVx1_ASAP7_75t_L g1688 ( 
.A(n_1619),
.Y(n_1688)
);

INVx2_ASAP7_75t_L g1689 ( 
.A(n_1653),
.Y(n_1689)
);

INVx1_ASAP7_75t_L g1690 ( 
.A(n_1623),
.Y(n_1690)
);

INVx1_ASAP7_75t_L g1691 ( 
.A(n_1623),
.Y(n_1691)
);

AOI22xp33_ASAP7_75t_L g1692 ( 
.A1(n_1632),
.A2(n_1625),
.B1(n_1612),
.B2(n_1631),
.Y(n_1692)
);

AND2x2_ASAP7_75t_L g1693 ( 
.A(n_1649),
.B(n_1566),
.Y(n_1693)
);

AND2x4_ASAP7_75t_L g1694 ( 
.A(n_1651),
.B(n_1594),
.Y(n_1694)
);

AND2x2_ASAP7_75t_L g1695 ( 
.A(n_1651),
.B(n_1567),
.Y(n_1695)
);

INVxp67_ASAP7_75t_L g1696 ( 
.A(n_1611),
.Y(n_1696)
);

INVx3_ASAP7_75t_L g1697 ( 
.A(n_1653),
.Y(n_1697)
);

NOR2xp67_ASAP7_75t_L g1698 ( 
.A(n_1637),
.B(n_1607),
.Y(n_1698)
);

INVx2_ASAP7_75t_L g1699 ( 
.A(n_1662),
.Y(n_1699)
);

BUFx6f_ASAP7_75t_L g1700 ( 
.A(n_1671),
.Y(n_1700)
);

AND2x2_ASAP7_75t_L g1701 ( 
.A(n_1664),
.B(n_1654),
.Y(n_1701)
);

INVx1_ASAP7_75t_L g1702 ( 
.A(n_1663),
.Y(n_1702)
);

NOR2xp33_ASAP7_75t_L g1703 ( 
.A(n_1696),
.B(n_1610),
.Y(n_1703)
);

INVx1_ASAP7_75t_L g1704 ( 
.A(n_1663),
.Y(n_1704)
);

INVx1_ASAP7_75t_L g1705 ( 
.A(n_1662),
.Y(n_1705)
);

NAND2xp5_ASAP7_75t_L g1706 ( 
.A(n_1669),
.B(n_1636),
.Y(n_1706)
);

AND2x2_ASAP7_75t_L g1707 ( 
.A(n_1664),
.B(n_1654),
.Y(n_1707)
);

NAND2xp5_ASAP7_75t_L g1708 ( 
.A(n_1666),
.B(n_1636),
.Y(n_1708)
);

NAND2xp5_ASAP7_75t_L g1709 ( 
.A(n_1687),
.B(n_1638),
.Y(n_1709)
);

NAND2xp5_ASAP7_75t_L g1710 ( 
.A(n_1679),
.B(n_1638),
.Y(n_1710)
);

OR2x2_ASAP7_75t_L g1711 ( 
.A(n_1661),
.B(n_1621),
.Y(n_1711)
);

INVx2_ASAP7_75t_SL g1712 ( 
.A(n_1660),
.Y(n_1712)
);

INVx1_ASAP7_75t_L g1713 ( 
.A(n_1668),
.Y(n_1713)
);

OR2x2_ASAP7_75t_L g1714 ( 
.A(n_1661),
.B(n_1622),
.Y(n_1714)
);

INVx2_ASAP7_75t_L g1715 ( 
.A(n_1684),
.Y(n_1715)
);

INVx1_ASAP7_75t_L g1716 ( 
.A(n_1668),
.Y(n_1716)
);

OR2x2_ASAP7_75t_L g1717 ( 
.A(n_1665),
.B(n_1642),
.Y(n_1717)
);

OR2x2_ASAP7_75t_L g1718 ( 
.A(n_1665),
.B(n_1642),
.Y(n_1718)
);

INVx2_ASAP7_75t_L g1719 ( 
.A(n_1689),
.Y(n_1719)
);

AND2x2_ASAP7_75t_L g1720 ( 
.A(n_1670),
.B(n_1659),
.Y(n_1720)
);

AND2x2_ASAP7_75t_L g1721 ( 
.A(n_1670),
.B(n_1616),
.Y(n_1721)
);

INVx1_ASAP7_75t_L g1722 ( 
.A(n_1672),
.Y(n_1722)
);

AOI21x1_ASAP7_75t_L g1723 ( 
.A1(n_1671),
.A2(n_1490),
.B(n_1603),
.Y(n_1723)
);

NOR2x1p5_ASAP7_75t_L g1724 ( 
.A(n_1697),
.B(n_1632),
.Y(n_1724)
);

AND2x2_ASAP7_75t_SL g1725 ( 
.A(n_1692),
.B(n_1640),
.Y(n_1725)
);

INVx1_ASAP7_75t_L g1726 ( 
.A(n_1672),
.Y(n_1726)
);

NAND2xp5_ASAP7_75t_L g1727 ( 
.A(n_1690),
.B(n_1691),
.Y(n_1727)
);

AND2x2_ASAP7_75t_L g1728 ( 
.A(n_1685),
.B(n_1616),
.Y(n_1728)
);

OR2x2_ASAP7_75t_L g1729 ( 
.A(n_1686),
.B(n_1645),
.Y(n_1729)
);

AND2x4_ASAP7_75t_L g1730 ( 
.A(n_1660),
.B(n_1620),
.Y(n_1730)
);

INVx1_ASAP7_75t_L g1731 ( 
.A(n_1673),
.Y(n_1731)
);

INVx2_ASAP7_75t_L g1732 ( 
.A(n_1689),
.Y(n_1732)
);

NAND2xp5_ASAP7_75t_L g1733 ( 
.A(n_1690),
.B(n_1645),
.Y(n_1733)
);

INVx2_ASAP7_75t_L g1734 ( 
.A(n_1689),
.Y(n_1734)
);

AND2x2_ASAP7_75t_L g1735 ( 
.A(n_1685),
.B(n_1620),
.Y(n_1735)
);

INVx2_ASAP7_75t_L g1736 ( 
.A(n_1684),
.Y(n_1736)
);

INVx1_ASAP7_75t_L g1737 ( 
.A(n_1673),
.Y(n_1737)
);

NAND2xp5_ASAP7_75t_L g1738 ( 
.A(n_1691),
.B(n_1646),
.Y(n_1738)
);

INVx1_ASAP7_75t_L g1739 ( 
.A(n_1677),
.Y(n_1739)
);

NOR2xp33_ASAP7_75t_L g1740 ( 
.A(n_1674),
.B(n_1610),
.Y(n_1740)
);

AND2x2_ASAP7_75t_L g1741 ( 
.A(n_1693),
.B(n_1647),
.Y(n_1741)
);

INVx1_ASAP7_75t_L g1742 ( 
.A(n_1677),
.Y(n_1742)
);

INVx2_ASAP7_75t_L g1743 ( 
.A(n_1699),
.Y(n_1743)
);

OR2x2_ASAP7_75t_L g1744 ( 
.A(n_1736),
.B(n_1686),
.Y(n_1744)
);

AOI22xp5_ASAP7_75t_L g1745 ( 
.A1(n_1725),
.A2(n_1698),
.B1(n_1683),
.B2(n_1644),
.Y(n_1745)
);

HB1xp67_ASAP7_75t_L g1746 ( 
.A(n_1724),
.Y(n_1746)
);

AND2x2_ASAP7_75t_L g1747 ( 
.A(n_1720),
.B(n_1697),
.Y(n_1747)
);

AND2x2_ASAP7_75t_L g1748 ( 
.A(n_1720),
.B(n_1697),
.Y(n_1748)
);

OR2x2_ASAP7_75t_L g1749 ( 
.A(n_1736),
.B(n_1688),
.Y(n_1749)
);

INVx1_ASAP7_75t_L g1750 ( 
.A(n_1702),
.Y(n_1750)
);

INVx2_ASAP7_75t_SL g1751 ( 
.A(n_1712),
.Y(n_1751)
);

AND2x2_ASAP7_75t_L g1752 ( 
.A(n_1712),
.B(n_1697),
.Y(n_1752)
);

INVxp67_ASAP7_75t_SL g1753 ( 
.A(n_1724),
.Y(n_1753)
);

INVx1_ASAP7_75t_SL g1754 ( 
.A(n_1706),
.Y(n_1754)
);

NOR2xp33_ASAP7_75t_L g1755 ( 
.A(n_1703),
.B(n_1430),
.Y(n_1755)
);

OR2x2_ASAP7_75t_L g1756 ( 
.A(n_1715),
.B(n_1688),
.Y(n_1756)
);

BUFx2_ASAP7_75t_L g1757 ( 
.A(n_1700),
.Y(n_1757)
);

INVx1_ASAP7_75t_L g1758 ( 
.A(n_1702),
.Y(n_1758)
);

AND2x2_ASAP7_75t_L g1759 ( 
.A(n_1701),
.B(n_1693),
.Y(n_1759)
);

HB1xp67_ASAP7_75t_L g1760 ( 
.A(n_1727),
.Y(n_1760)
);

INVx2_ASAP7_75t_SL g1761 ( 
.A(n_1700),
.Y(n_1761)
);

INVx1_ASAP7_75t_L g1762 ( 
.A(n_1704),
.Y(n_1762)
);

AND2x2_ASAP7_75t_L g1763 ( 
.A(n_1701),
.B(n_1695),
.Y(n_1763)
);

OR2x2_ASAP7_75t_L g1764 ( 
.A(n_1715),
.B(n_1711),
.Y(n_1764)
);

NAND2xp5_ASAP7_75t_L g1765 ( 
.A(n_1740),
.B(n_1680),
.Y(n_1765)
);

AOI22xp5_ASAP7_75t_L g1766 ( 
.A1(n_1725),
.A2(n_1698),
.B1(n_1683),
.B2(n_1644),
.Y(n_1766)
);

INVx1_ASAP7_75t_L g1767 ( 
.A(n_1704),
.Y(n_1767)
);

NAND2x1p5_ASAP7_75t_L g1768 ( 
.A(n_1700),
.B(n_1594),
.Y(n_1768)
);

NAND2xp5_ASAP7_75t_L g1769 ( 
.A(n_1725),
.B(n_1678),
.Y(n_1769)
);

OR2x2_ASAP7_75t_L g1770 ( 
.A(n_1715),
.B(n_1675),
.Y(n_1770)
);

AND2x2_ASAP7_75t_L g1771 ( 
.A(n_1707),
.B(n_1695),
.Y(n_1771)
);

INVx2_ASAP7_75t_L g1772 ( 
.A(n_1699),
.Y(n_1772)
);

INVxp67_ASAP7_75t_L g1773 ( 
.A(n_1708),
.Y(n_1773)
);

NAND2xp5_ASAP7_75t_SL g1774 ( 
.A(n_1700),
.B(n_1630),
.Y(n_1774)
);

OR2x2_ASAP7_75t_L g1775 ( 
.A(n_1711),
.B(n_1675),
.Y(n_1775)
);

NOR2xp33_ASAP7_75t_L g1776 ( 
.A(n_1710),
.B(n_1430),
.Y(n_1776)
);

AND2x2_ASAP7_75t_L g1777 ( 
.A(n_1707),
.B(n_1660),
.Y(n_1777)
);

AND2x2_ASAP7_75t_L g1778 ( 
.A(n_1730),
.B(n_1681),
.Y(n_1778)
);

AND2x2_ASAP7_75t_L g1779 ( 
.A(n_1730),
.B(n_1681),
.Y(n_1779)
);

OR2x2_ASAP7_75t_L g1780 ( 
.A(n_1714),
.B(n_1676),
.Y(n_1780)
);

INVx2_ASAP7_75t_L g1781 ( 
.A(n_1699),
.Y(n_1781)
);

NOR2xp33_ASAP7_75t_L g1782 ( 
.A(n_1709),
.B(n_1682),
.Y(n_1782)
);

NAND2xp5_ASAP7_75t_L g1783 ( 
.A(n_1733),
.B(n_1678),
.Y(n_1783)
);

NAND2xp5_ASAP7_75t_L g1784 ( 
.A(n_1738),
.B(n_1721),
.Y(n_1784)
);

INVx1_ASAP7_75t_L g1785 ( 
.A(n_1713),
.Y(n_1785)
);

AND2x4_ASAP7_75t_L g1786 ( 
.A(n_1730),
.B(n_1694),
.Y(n_1786)
);

INVx2_ASAP7_75t_L g1787 ( 
.A(n_1719),
.Y(n_1787)
);

INVx1_ASAP7_75t_L g1788 ( 
.A(n_1713),
.Y(n_1788)
);

AOI22xp33_ASAP7_75t_L g1789 ( 
.A1(n_1746),
.A2(n_1700),
.B1(n_1637),
.B2(n_1652),
.Y(n_1789)
);

NOR2xp33_ASAP7_75t_L g1790 ( 
.A(n_1755),
.B(n_1728),
.Y(n_1790)
);

OR2x2_ASAP7_75t_L g1791 ( 
.A(n_1769),
.B(n_1714),
.Y(n_1791)
);

BUFx3_ASAP7_75t_L g1792 ( 
.A(n_1757),
.Y(n_1792)
);

INVxp67_ASAP7_75t_L g1793 ( 
.A(n_1753),
.Y(n_1793)
);

OR2x2_ASAP7_75t_L g1794 ( 
.A(n_1764),
.B(n_1729),
.Y(n_1794)
);

AND2x2_ASAP7_75t_L g1795 ( 
.A(n_1778),
.B(n_1730),
.Y(n_1795)
);

AND2x2_ASAP7_75t_L g1796 ( 
.A(n_1778),
.B(n_1721),
.Y(n_1796)
);

INVx1_ASAP7_75t_L g1797 ( 
.A(n_1750),
.Y(n_1797)
);

INVx1_ASAP7_75t_L g1798 ( 
.A(n_1750),
.Y(n_1798)
);

INVx1_ASAP7_75t_SL g1799 ( 
.A(n_1757),
.Y(n_1799)
);

INVx1_ASAP7_75t_SL g1800 ( 
.A(n_1751),
.Y(n_1800)
);

INVx1_ASAP7_75t_L g1801 ( 
.A(n_1758),
.Y(n_1801)
);

AND2x4_ASAP7_75t_SL g1802 ( 
.A(n_1786),
.B(n_1667),
.Y(n_1802)
);

NAND2xp5_ASAP7_75t_L g1803 ( 
.A(n_1754),
.B(n_1741),
.Y(n_1803)
);

INVx3_ASAP7_75t_SL g1804 ( 
.A(n_1774),
.Y(n_1804)
);

OR2x2_ASAP7_75t_L g1805 ( 
.A(n_1764),
.B(n_1729),
.Y(n_1805)
);

INVx2_ASAP7_75t_L g1806 ( 
.A(n_1747),
.Y(n_1806)
);

OAI22xp5_ASAP7_75t_L g1807 ( 
.A1(n_1745),
.A2(n_1627),
.B1(n_1648),
.B2(n_1634),
.Y(n_1807)
);

AOI22xp33_ASAP7_75t_L g1808 ( 
.A1(n_1765),
.A2(n_1630),
.B1(n_1694),
.B2(n_1597),
.Y(n_1808)
);

INVx1_ASAP7_75t_L g1809 ( 
.A(n_1758),
.Y(n_1809)
);

NAND2xp5_ASAP7_75t_L g1810 ( 
.A(n_1782),
.B(n_1741),
.Y(n_1810)
);

INVx2_ASAP7_75t_SL g1811 ( 
.A(n_1786),
.Y(n_1811)
);

INVx1_ASAP7_75t_SL g1812 ( 
.A(n_1751),
.Y(n_1812)
);

NOR2xp33_ASAP7_75t_L g1813 ( 
.A(n_1776),
.B(n_1728),
.Y(n_1813)
);

NAND2xp5_ASAP7_75t_L g1814 ( 
.A(n_1773),
.B(n_1735),
.Y(n_1814)
);

AND2x2_ASAP7_75t_L g1815 ( 
.A(n_1779),
.B(n_1735),
.Y(n_1815)
);

AND2x2_ASAP7_75t_L g1816 ( 
.A(n_1779),
.B(n_1719),
.Y(n_1816)
);

OR2x2_ASAP7_75t_L g1817 ( 
.A(n_1775),
.B(n_1717),
.Y(n_1817)
);

NAND2x1_ASAP7_75t_L g1818 ( 
.A(n_1786),
.B(n_1716),
.Y(n_1818)
);

AND2x2_ASAP7_75t_L g1819 ( 
.A(n_1777),
.B(n_1732),
.Y(n_1819)
);

NAND2xp5_ASAP7_75t_L g1820 ( 
.A(n_1760),
.B(n_1717),
.Y(n_1820)
);

AND2x2_ASAP7_75t_L g1821 ( 
.A(n_1777),
.B(n_1732),
.Y(n_1821)
);

NAND2xp5_ASAP7_75t_L g1822 ( 
.A(n_1784),
.B(n_1759),
.Y(n_1822)
);

INVx1_ASAP7_75t_SL g1823 ( 
.A(n_1752),
.Y(n_1823)
);

HB1xp67_ASAP7_75t_L g1824 ( 
.A(n_1785),
.Y(n_1824)
);

INVx1_ASAP7_75t_L g1825 ( 
.A(n_1762),
.Y(n_1825)
);

INVx2_ASAP7_75t_L g1826 ( 
.A(n_1747),
.Y(n_1826)
);

OAI211xp5_ASAP7_75t_SL g1827 ( 
.A1(n_1793),
.A2(n_1789),
.B(n_1799),
.C(n_1807),
.Y(n_1827)
);

NAND2xp5_ASAP7_75t_L g1828 ( 
.A(n_1804),
.B(n_1759),
.Y(n_1828)
);

AOI22xp33_ASAP7_75t_SL g1829 ( 
.A1(n_1802),
.A2(n_1790),
.B1(n_1813),
.B2(n_1795),
.Y(n_1829)
);

INVx1_ASAP7_75t_L g1830 ( 
.A(n_1824),
.Y(n_1830)
);

XOR2x2_ASAP7_75t_L g1831 ( 
.A(n_1804),
.B(n_1766),
.Y(n_1831)
);

INVx2_ASAP7_75t_L g1832 ( 
.A(n_1792),
.Y(n_1832)
);

OAI221xp5_ASAP7_75t_L g1833 ( 
.A1(n_1804),
.A2(n_1761),
.B1(n_1634),
.B2(n_1768),
.C(n_1770),
.Y(n_1833)
);

OAI21xp33_ASAP7_75t_L g1834 ( 
.A1(n_1800),
.A2(n_1770),
.B(n_1744),
.Y(n_1834)
);

INVx1_ASAP7_75t_L g1835 ( 
.A(n_1797),
.Y(n_1835)
);

INVx1_ASAP7_75t_L g1836 ( 
.A(n_1797),
.Y(n_1836)
);

HB1xp67_ASAP7_75t_L g1837 ( 
.A(n_1792),
.Y(n_1837)
);

INVx1_ASAP7_75t_L g1838 ( 
.A(n_1798),
.Y(n_1838)
);

NAND2xp5_ASAP7_75t_L g1839 ( 
.A(n_1812),
.B(n_1763),
.Y(n_1839)
);

AOI21xp33_ASAP7_75t_SL g1840 ( 
.A1(n_1811),
.A2(n_1761),
.B(n_1768),
.Y(n_1840)
);

NAND3xp33_ASAP7_75t_SL g1841 ( 
.A(n_1823),
.B(n_1768),
.C(n_1775),
.Y(n_1841)
);

NAND2xp5_ASAP7_75t_L g1842 ( 
.A(n_1796),
.B(n_1763),
.Y(n_1842)
);

INVxp67_ASAP7_75t_L g1843 ( 
.A(n_1811),
.Y(n_1843)
);

NAND2xp5_ASAP7_75t_L g1844 ( 
.A(n_1796),
.B(n_1771),
.Y(n_1844)
);

INVx1_ASAP7_75t_L g1845 ( 
.A(n_1798),
.Y(n_1845)
);

NAND2xp5_ASAP7_75t_L g1846 ( 
.A(n_1810),
.B(n_1771),
.Y(n_1846)
);

NAND2xp5_ASAP7_75t_L g1847 ( 
.A(n_1815),
.B(n_1783),
.Y(n_1847)
);

NAND2xp5_ASAP7_75t_L g1848 ( 
.A(n_1815),
.B(n_1748),
.Y(n_1848)
);

OAI22xp5_ASAP7_75t_L g1849 ( 
.A1(n_1808),
.A2(n_1648),
.B1(n_1748),
.B2(n_1780),
.Y(n_1849)
);

INVx1_ASAP7_75t_L g1850 ( 
.A(n_1801),
.Y(n_1850)
);

INVxp67_ASAP7_75t_L g1851 ( 
.A(n_1806),
.Y(n_1851)
);

O2A1O1Ixp5_ASAP7_75t_L g1852 ( 
.A1(n_1818),
.A2(n_1785),
.B(n_1788),
.C(n_1752),
.Y(n_1852)
);

INVx1_ASAP7_75t_L g1853 ( 
.A(n_1801),
.Y(n_1853)
);

NOR3xp33_ASAP7_75t_L g1854 ( 
.A(n_1791),
.B(n_1818),
.C(n_1820),
.Y(n_1854)
);

INVx2_ASAP7_75t_SL g1855 ( 
.A(n_1837),
.Y(n_1855)
);

INVx1_ASAP7_75t_L g1856 ( 
.A(n_1837),
.Y(n_1856)
);

INVx1_ASAP7_75t_L g1857 ( 
.A(n_1835),
.Y(n_1857)
);

AND2x2_ASAP7_75t_L g1858 ( 
.A(n_1829),
.B(n_1795),
.Y(n_1858)
);

NOR2xp33_ASAP7_75t_L g1859 ( 
.A(n_1827),
.B(n_1822),
.Y(n_1859)
);

INVx1_ASAP7_75t_L g1860 ( 
.A(n_1836),
.Y(n_1860)
);

INVx2_ASAP7_75t_L g1861 ( 
.A(n_1832),
.Y(n_1861)
);

NAND2xp5_ASAP7_75t_L g1862 ( 
.A(n_1830),
.B(n_1832),
.Y(n_1862)
);

AOI21xp5_ASAP7_75t_L g1863 ( 
.A1(n_1831),
.A2(n_1803),
.B(n_1814),
.Y(n_1863)
);

AOI221xp5_ASAP7_75t_L g1864 ( 
.A1(n_1854),
.A2(n_1826),
.B1(n_1806),
.B2(n_1809),
.C(n_1825),
.Y(n_1864)
);

NAND2xp5_ASAP7_75t_L g1865 ( 
.A(n_1851),
.B(n_1791),
.Y(n_1865)
);

NAND2xp5_ASAP7_75t_L g1866 ( 
.A(n_1843),
.B(n_1826),
.Y(n_1866)
);

NAND2x1p5_ASAP7_75t_L g1867 ( 
.A(n_1828),
.B(n_1427),
.Y(n_1867)
);

NOR2xp33_ASAP7_75t_L g1868 ( 
.A(n_1834),
.B(n_1817),
.Y(n_1868)
);

AOI22xp5_ASAP7_75t_L g1869 ( 
.A1(n_1831),
.A2(n_1802),
.B1(n_1821),
.B2(n_1819),
.Y(n_1869)
);

NAND2xp5_ASAP7_75t_L g1870 ( 
.A(n_1839),
.B(n_1819),
.Y(n_1870)
);

NAND2xp5_ASAP7_75t_L g1871 ( 
.A(n_1854),
.B(n_1821),
.Y(n_1871)
);

AND2x2_ASAP7_75t_L g1872 ( 
.A(n_1842),
.B(n_1816),
.Y(n_1872)
);

NAND2xp5_ASAP7_75t_L g1873 ( 
.A(n_1838),
.B(n_1825),
.Y(n_1873)
);

NOR2xp33_ASAP7_75t_L g1874 ( 
.A(n_1846),
.B(n_1817),
.Y(n_1874)
);

AND2x2_ASAP7_75t_L g1875 ( 
.A(n_1844),
.B(n_1816),
.Y(n_1875)
);

NOR3xp33_ASAP7_75t_L g1876 ( 
.A(n_1862),
.B(n_1841),
.C(n_1833),
.Y(n_1876)
);

INVx1_ASAP7_75t_L g1877 ( 
.A(n_1855),
.Y(n_1877)
);

NOR2x1_ASAP7_75t_L g1878 ( 
.A(n_1856),
.B(n_1845),
.Y(n_1878)
);

OAI211xp5_ASAP7_75t_L g1879 ( 
.A1(n_1871),
.A2(n_1840),
.B(n_1853),
.C(n_1850),
.Y(n_1879)
);

NOR2xp67_ASAP7_75t_SL g1880 ( 
.A(n_1861),
.B(n_1794),
.Y(n_1880)
);

NAND2xp5_ASAP7_75t_L g1881 ( 
.A(n_1868),
.B(n_1848),
.Y(n_1881)
);

NAND2xp5_ASAP7_75t_L g1882 ( 
.A(n_1863),
.B(n_1847),
.Y(n_1882)
);

NOR2x1_ASAP7_75t_L g1883 ( 
.A(n_1862),
.B(n_1809),
.Y(n_1883)
);

AOI211xp5_ASAP7_75t_L g1884 ( 
.A1(n_1859),
.A2(n_1849),
.B(n_1794),
.C(n_1805),
.Y(n_1884)
);

OAI221xp5_ASAP7_75t_L g1885 ( 
.A1(n_1869),
.A2(n_1852),
.B1(n_1805),
.B2(n_1744),
.C(n_1780),
.Y(n_1885)
);

OAI221xp5_ASAP7_75t_L g1886 ( 
.A1(n_1874),
.A2(n_1762),
.B1(n_1767),
.B2(n_1756),
.C(n_1749),
.Y(n_1886)
);

NOR2x1_ASAP7_75t_L g1887 ( 
.A(n_1857),
.B(n_1743),
.Y(n_1887)
);

OR2x6_ASAP7_75t_L g1888 ( 
.A(n_1865),
.B(n_1866),
.Y(n_1888)
);

NOR4xp25_ASAP7_75t_L g1889 ( 
.A(n_1879),
.B(n_1860),
.C(n_1864),
.D(n_1873),
.Y(n_1889)
);

AND3x4_ASAP7_75t_L g1890 ( 
.A(n_1876),
.B(n_1858),
.C(n_1870),
.Y(n_1890)
);

NOR2xp33_ASAP7_75t_L g1891 ( 
.A(n_1882),
.B(n_1865),
.Y(n_1891)
);

OAI211xp5_ASAP7_75t_L g1892 ( 
.A1(n_1878),
.A2(n_1884),
.B(n_1885),
.C(n_1883),
.Y(n_1892)
);

INVx1_ASAP7_75t_L g1893 ( 
.A(n_1877),
.Y(n_1893)
);

AND2x2_ASAP7_75t_L g1894 ( 
.A(n_1888),
.B(n_1872),
.Y(n_1894)
);

NOR3xp33_ASAP7_75t_L g1895 ( 
.A(n_1881),
.B(n_1873),
.C(n_1875),
.Y(n_1895)
);

AND2x4_ASAP7_75t_L g1896 ( 
.A(n_1888),
.B(n_1787),
.Y(n_1896)
);

NOR3xp33_ASAP7_75t_L g1897 ( 
.A(n_1886),
.B(n_1867),
.C(n_1772),
.Y(n_1897)
);

INVx2_ASAP7_75t_SL g1898 ( 
.A(n_1887),
.Y(n_1898)
);

NAND2xp5_ASAP7_75t_L g1899 ( 
.A(n_1880),
.B(n_1867),
.Y(n_1899)
);

OAI21x1_ASAP7_75t_L g1900 ( 
.A1(n_1878),
.A2(n_1772),
.B(n_1743),
.Y(n_1900)
);

NAND4xp25_ASAP7_75t_SL g1901 ( 
.A(n_1892),
.B(n_1895),
.C(n_1894),
.D(n_1899),
.Y(n_1901)
);

NAND4xp25_ASAP7_75t_L g1902 ( 
.A(n_1891),
.B(n_1756),
.C(n_1641),
.D(n_1749),
.Y(n_1902)
);

INVx1_ASAP7_75t_L g1903 ( 
.A(n_1898),
.Y(n_1903)
);

NAND2xp5_ASAP7_75t_L g1904 ( 
.A(n_1889),
.B(n_1787),
.Y(n_1904)
);

NOR2x1_ASAP7_75t_L g1905 ( 
.A(n_1893),
.B(n_1781),
.Y(n_1905)
);

NOR3xp33_ASAP7_75t_L g1906 ( 
.A(n_1897),
.B(n_1449),
.C(n_1781),
.Y(n_1906)
);

NOR3xp33_ASAP7_75t_L g1907 ( 
.A(n_1896),
.B(n_1593),
.C(n_1442),
.Y(n_1907)
);

AOI221xp5_ASAP7_75t_L g1908 ( 
.A1(n_1896),
.A2(n_1742),
.B1(n_1739),
.B2(n_1737),
.C(n_1716),
.Y(n_1908)
);

INVxp67_ASAP7_75t_SL g1909 ( 
.A(n_1904),
.Y(n_1909)
);

INVx1_ASAP7_75t_L g1910 ( 
.A(n_1903),
.Y(n_1910)
);

INVx1_ASAP7_75t_L g1911 ( 
.A(n_1905),
.Y(n_1911)
);

INVx1_ASAP7_75t_L g1912 ( 
.A(n_1902),
.Y(n_1912)
);

INVx1_ASAP7_75t_L g1913 ( 
.A(n_1906),
.Y(n_1913)
);

INVx2_ASAP7_75t_L g1914 ( 
.A(n_1901),
.Y(n_1914)
);

INVx1_ASAP7_75t_L g1915 ( 
.A(n_1907),
.Y(n_1915)
);

NOR2x1_ASAP7_75t_L g1916 ( 
.A(n_1908),
.B(n_1890),
.Y(n_1916)
);

NAND4xp25_ASAP7_75t_L g1917 ( 
.A(n_1916),
.B(n_1900),
.C(n_1442),
.D(n_1460),
.Y(n_1917)
);

NAND4xp75_ASAP7_75t_L g1918 ( 
.A(n_1910),
.B(n_1462),
.C(n_1448),
.D(n_1434),
.Y(n_1918)
);

AND3x2_ASAP7_75t_L g1919 ( 
.A(n_1909),
.B(n_1911),
.C(n_1914),
.Y(n_1919)
);

AND2x2_ASAP7_75t_L g1920 ( 
.A(n_1912),
.B(n_1718),
.Y(n_1920)
);

NOR3xp33_ASAP7_75t_L g1921 ( 
.A(n_1913),
.B(n_1448),
.C(n_1434),
.Y(n_1921)
);

AOI211xp5_ASAP7_75t_L g1922 ( 
.A1(n_1909),
.A2(n_1462),
.B(n_1739),
.C(n_1737),
.Y(n_1922)
);

INVx1_ASAP7_75t_L g1923 ( 
.A(n_1919),
.Y(n_1923)
);

INVx1_ASAP7_75t_L g1924 ( 
.A(n_1920),
.Y(n_1924)
);

INVx1_ASAP7_75t_L g1925 ( 
.A(n_1917),
.Y(n_1925)
);

INVx1_ASAP7_75t_L g1926 ( 
.A(n_1922),
.Y(n_1926)
);

AOI22xp5_ASAP7_75t_L g1927 ( 
.A1(n_1924),
.A2(n_1915),
.B1(n_1921),
.B2(n_1918),
.Y(n_1927)
);

INVx1_ASAP7_75t_L g1928 ( 
.A(n_1923),
.Y(n_1928)
);

INVx1_ASAP7_75t_L g1929 ( 
.A(n_1928),
.Y(n_1929)
);

AOI211x1_ASAP7_75t_L g1930 ( 
.A1(n_1929),
.A2(n_1926),
.B(n_1925),
.C(n_1927),
.Y(n_1930)
);

AOI22xp33_ASAP7_75t_L g1931 ( 
.A1(n_1929),
.A2(n_1742),
.B1(n_1722),
.B2(n_1731),
.Y(n_1931)
);

AO22x2_ASAP7_75t_L g1932 ( 
.A1(n_1930),
.A2(n_1722),
.B1(n_1731),
.B2(n_1726),
.Y(n_1932)
);

INVx2_ASAP7_75t_L g1933 ( 
.A(n_1931),
.Y(n_1933)
);

OAI22xp5_ASAP7_75t_L g1934 ( 
.A1(n_1933),
.A2(n_1726),
.B1(n_1734),
.B2(n_1718),
.Y(n_1934)
);

NAND2xp5_ASAP7_75t_SL g1935 ( 
.A(n_1934),
.B(n_1932),
.Y(n_1935)
);

AOI22xp33_ASAP7_75t_L g1936 ( 
.A1(n_1935),
.A2(n_1432),
.B1(n_1734),
.B2(n_1705),
.Y(n_1936)
);

OAI221xp5_ASAP7_75t_R g1937 ( 
.A1(n_1936),
.A2(n_1432),
.B1(n_1658),
.B2(n_1723),
.C(n_1705),
.Y(n_1937)
);

AOI211xp5_ASAP7_75t_L g1938 ( 
.A1(n_1937),
.A2(n_1464),
.B(n_1458),
.C(n_1406),
.Y(n_1938)
);


endmodule