module real_jpeg_5060_n_16 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_3, n_10, n_9, n_16);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_16;

wire n_384;
wire n_37;
wire n_430;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_460;
wire n_300;
wire n_415;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_446;
wire n_199;
wire n_95;
wire n_441;
wire n_238;
wire n_67;
wire n_350;
wire n_235;
wire n_107;
wire n_369;
wire n_376;
wire n_354;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_355;
wire n_123;
wire n_463;
wire n_425;
wire n_455;
wire n_462;
wire n_50;
wire n_409;
wire n_186;
wire n_137;
wire n_72;
wire n_440;
wire n_171;
wire n_151;
wire n_272;
wire n_461;
wire n_198;
wire n_203;
wire n_23;
wire n_362;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_326;
wire n_339;
wire n_80;
wire n_30;
wire n_328;
wire n_149;
wire n_332;
wire n_366;
wire n_456;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_353;
wire n_453;
wire n_230;
wire n_417;
wire n_428;
wire n_216;
wire n_128;
wire n_202;
wire n_367;
wire n_127;
wire n_356;
wire n_365;
wire n_423;
wire n_464;
wire n_36;
wire n_102;
wire n_81;
wire n_101;
wire n_422;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_348;
wire n_252;
wire n_363;
wire n_310;
wire n_345;
wire n_78;
wire n_83;
wire n_288;
wire n_221;
wire n_393;
wire n_104;
wire n_153;
wire n_443;
wire n_337;
wire n_131;
wire n_439;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_378;
wire n_200;
wire n_432;
wire n_465;
wire n_335;
wire n_214;
wire n_113;
wire n_251;
wire n_459;
wire n_139;
wire n_33;
wire n_175;
wire n_338;
wire n_156;
wire n_387;
wire n_434;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_390;
wire n_77;
wire n_399;
wire n_372;
wire n_219;
wire n_122;
wire n_19;
wire n_262;
wire n_334;
wire n_17;
wire n_383;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_426;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_371;
wire n_410;
wire n_421;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_382;
wire n_411;
wire n_20;
wire n_278;
wire n_314;
wire n_103;
wire n_232;
wire n_448;
wire n_212;
wire n_284;
wire n_402;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_452;
wire n_213;
wire n_25;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_407;
wire n_419;
wire n_386;
wire n_341;
wire n_331;
wire n_49;
wire n_68;
wire n_395;
wire n_146;
wire n_323;
wire n_215;
wire n_176;
wire n_166;
wire n_286;
wire n_312;
wire n_325;
wire n_307;
wire n_316;
wire n_161;
wire n_207;
wire n_431;
wire n_420;
wire n_357;
wire n_237;
wire n_445;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_380;
wire n_414;
wire n_140;
wire n_126;
wire n_342;
wire n_120;
wire n_155;
wire n_412;
wire n_405;
wire n_319;
wire n_93;
wire n_242;
wire n_142;
wire n_397;
wire n_76;
wire n_403;
wire n_79;
wire n_282;
wire n_147;
wire n_359;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_449;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_18;
wire n_145;
wire n_266;
wire n_377;
wire n_109;
wire n_391;
wire n_427;
wire n_401;
wire n_148;
wire n_373;
wire n_396;
wire n_392;
wire n_196;
wire n_375;
wire n_330;
wire n_298;
wire n_333;
wire n_450;
wire n_152;
wire n_270;
wire n_159;
wire n_429;
wire n_347;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_336;
wire n_258;
wire n_458;
wire n_150;
wire n_41;
wire n_74;
wire n_404;
wire n_158;
wire n_204;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_413;
wire n_75;
wire n_346;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_457;
wire n_119;
wire n_283;
wire n_181;
wire n_358;
wire n_256;
wire n_273;
wire n_253;
wire n_54;
wire n_168;
wire n_38;
wire n_442;
wire n_385;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_349;
wire n_418;
wire n_343;
wire n_292;
wire n_64;
wire n_291;
wire n_236;
wire n_370;
wire n_276;
wire n_374;
wire n_287;
wire n_400;
wire n_174;
wire n_388;
wire n_255;
wire n_243;
wire n_299;
wire n_352;
wire n_56;
wire n_293;
wire n_275;
wire n_381;
wire n_227;
wire n_229;
wire n_454;
wire n_379;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_444;
wire n_360;
wire n_398;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_451;
wire n_45;
wire n_437;
wire n_268;
wire n_42;
wire n_313;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_416;
wire n_143;
wire n_351;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_406;
wire n_303;
wire n_321;
wire n_100;
wire n_368;
wire n_51;
wire n_205;
wire n_361;
wire n_261;
wire n_86;
wire n_324;
wire n_70;
wire n_435;
wire n_32;
wire n_228;
wire n_389;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_438;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_394;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_436;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_424;
wire n_133;
wire n_257;
wire n_447;
wire n_344;
wire n_210;
wire n_206;
wire n_408;
wire n_85;
wire n_96;
wire n_308;
wire n_433;
wire n_364;

INVx8_ASAP7_75t_L g78 ( 
.A(n_0),
.Y(n_78)
);

AOI22xp5_ASAP7_75t_L g100 ( 
.A1(n_1),
.A2(n_93),
.B1(n_101),
.B2(n_102),
.Y(n_100)
);

CKINVDCx20_ASAP7_75t_R g102 ( 
.A(n_1),
.Y(n_102)
);

AOI22xp5_ASAP7_75t_L g137 ( 
.A1(n_1),
.A2(n_102),
.B1(n_138),
.B2(n_140),
.Y(n_137)
);

AOI22xp5_ASAP7_75t_SL g215 ( 
.A1(n_1),
.A2(n_60),
.B1(n_102),
.B2(n_216),
.Y(n_215)
);

OAI22xp5_ASAP7_75t_SL g279 ( 
.A1(n_1),
.A2(n_102),
.B1(n_280),
.B2(n_282),
.Y(n_279)
);

AOI22xp5_ASAP7_75t_L g128 ( 
.A1(n_2),
.A2(n_28),
.B1(n_129),
.B2(n_130),
.Y(n_128)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_2),
.Y(n_129)
);

AOI22xp5_ASAP7_75t_L g175 ( 
.A1(n_2),
.A2(n_129),
.B1(n_176),
.B2(n_178),
.Y(n_175)
);

OAI22xp5_ASAP7_75t_L g342 ( 
.A1(n_2),
.A2(n_129),
.B1(n_343),
.B2(n_346),
.Y(n_342)
);

AOI22xp33_ASAP7_75t_L g359 ( 
.A1(n_2),
.A2(n_129),
.B1(n_192),
.B2(n_360),
.Y(n_359)
);

INVx2_ASAP7_75t_L g52 ( 
.A(n_3),
.Y(n_52)
);

BUFx3_ASAP7_75t_L g61 ( 
.A(n_3),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g190 ( 
.A(n_3),
.Y(n_190)
);

OAI22xp5_ASAP7_75t_SL g92 ( 
.A1(n_4),
.A2(n_93),
.B1(n_96),
.B2(n_97),
.Y(n_92)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_4),
.Y(n_96)
);

AOI22xp33_ASAP7_75t_L g232 ( 
.A1(n_4),
.A2(n_96),
.B1(n_233),
.B2(n_235),
.Y(n_232)
);

AOI22xp33_ASAP7_75t_SL g349 ( 
.A1(n_4),
.A2(n_96),
.B1(n_350),
.B2(n_352),
.Y(n_349)
);

OAI22xp5_ASAP7_75t_L g412 ( 
.A1(n_4),
.A2(n_96),
.B1(n_413),
.B2(n_414),
.Y(n_412)
);

AOI22xp5_ASAP7_75t_L g67 ( 
.A1(n_5),
.A2(n_59),
.B1(n_68),
.B2(n_69),
.Y(n_67)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_5),
.Y(n_68)
);

OAI22xp5_ASAP7_75t_L g206 ( 
.A1(n_5),
.A2(n_68),
.B1(n_207),
.B2(n_208),
.Y(n_206)
);

OAI22xp5_ASAP7_75t_L g294 ( 
.A1(n_5),
.A2(n_68),
.B1(n_94),
.B2(n_295),
.Y(n_294)
);

INVx6_ASAP7_75t_L g81 ( 
.A(n_6),
.Y(n_81)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_7),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_7),
.Y(n_66)
);

INVx8_ASAP7_75t_L g220 ( 
.A(n_7),
.Y(n_220)
);

BUFx6f_ASAP7_75t_L g374 ( 
.A(n_7),
.Y(n_374)
);

OAI22xp5_ASAP7_75t_SL g57 ( 
.A1(n_8),
.A2(n_58),
.B1(n_62),
.B2(n_63),
.Y(n_57)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_8),
.Y(n_62)
);

AOI22xp33_ASAP7_75t_L g196 ( 
.A1(n_8),
.A2(n_62),
.B1(n_140),
.B2(n_197),
.Y(n_196)
);

AOI22xp33_ASAP7_75t_L g272 ( 
.A1(n_8),
.A2(n_62),
.B1(n_177),
.B2(n_273),
.Y(n_272)
);

AOI22xp33_ASAP7_75t_SL g457 ( 
.A1(n_8),
.A2(n_62),
.B1(n_112),
.B2(n_458),
.Y(n_457)
);

OAI22xp5_ASAP7_75t_SL g104 ( 
.A1(n_9),
.A2(n_30),
.B1(n_105),
.B2(n_108),
.Y(n_104)
);

CKINVDCx20_ASAP7_75t_R g108 ( 
.A(n_9),
.Y(n_108)
);

OAI22xp5_ASAP7_75t_L g249 ( 
.A1(n_9),
.A2(n_108),
.B1(n_229),
.B2(n_250),
.Y(n_249)
);

OAI22xp5_ASAP7_75t_L g334 ( 
.A1(n_9),
.A2(n_108),
.B1(n_140),
.B2(n_335),
.Y(n_334)
);

AOI22xp5_ASAP7_75t_L g369 ( 
.A1(n_9),
.A2(n_108),
.B1(n_370),
.B2(n_372),
.Y(n_369)
);

INVx3_ASAP7_75t_L g34 ( 
.A(n_10),
.Y(n_34)
);

BUFx5_ASAP7_75t_L g115 ( 
.A(n_10),
.Y(n_115)
);

INVx3_ASAP7_75t_L g119 ( 
.A(n_10),
.Y(n_119)
);

BUFx6f_ASAP7_75t_L g124 ( 
.A(n_10),
.Y(n_124)
);

INVx8_ASAP7_75t_L g27 ( 
.A(n_11),
.Y(n_27)
);

INVx6_ASAP7_75t_L g30 ( 
.A(n_12),
.Y(n_30)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_12),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g107 ( 
.A(n_12),
.Y(n_107)
);

INVx3_ASAP7_75t_L g113 ( 
.A(n_12),
.Y(n_113)
);

BUFx6f_ASAP7_75t_L g117 ( 
.A(n_12),
.Y(n_117)
);

BUFx6f_ASAP7_75t_L g132 ( 
.A(n_12),
.Y(n_132)
);

BUFx6f_ASAP7_75t_L g234 ( 
.A(n_12),
.Y(n_234)
);

INVx2_ASAP7_75t_L g281 ( 
.A(n_12),
.Y(n_281)
);

INVx2_ASAP7_75t_L g148 ( 
.A(n_13),
.Y(n_148)
);

INVx3_ASAP7_75t_L g151 ( 
.A(n_13),
.Y(n_151)
);

BUFx3_ASAP7_75t_L g157 ( 
.A(n_13),
.Y(n_157)
);

OAI22xp33_ASAP7_75t_SL g164 ( 
.A1(n_14),
.A2(n_165),
.B1(n_168),
.B2(n_169),
.Y(n_164)
);

CKINVDCx20_ASAP7_75t_R g168 ( 
.A(n_14),
.Y(n_168)
);

AOI22xp33_ASAP7_75t_L g187 ( 
.A1(n_14),
.A2(n_168),
.B1(n_188),
.B2(n_191),
.Y(n_187)
);

OAI22xp5_ASAP7_75t_SL g227 ( 
.A1(n_14),
.A2(n_88),
.B1(n_168),
.B2(n_228),
.Y(n_227)
);

AOI22xp33_ASAP7_75t_L g305 ( 
.A1(n_14),
.A2(n_30),
.B1(n_117),
.B2(n_168),
.Y(n_305)
);

NOR2xp33_ASAP7_75t_L g42 ( 
.A(n_15),
.B(n_43),
.Y(n_42)
);

AOI21xp5_ASAP7_75t_L g172 ( 
.A1(n_15),
.A2(n_42),
.B(n_116),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_L g246 ( 
.A(n_15),
.B(n_133),
.Y(n_246)
);

MAJIxp5_ASAP7_75t_L g318 ( 
.A(n_15),
.B(n_319),
.C(n_323),
.Y(n_318)
);

OAI22xp33_ASAP7_75t_L g328 ( 
.A1(n_15),
.A2(n_329),
.B1(n_330),
.B2(n_333),
.Y(n_328)
);

CKINVDCx20_ASAP7_75t_R g329 ( 
.A(n_15),
.Y(n_329)
);

NAND2xp5_ASAP7_75t_L g340 ( 
.A(n_15),
.B(n_226),
.Y(n_340)
);

OAI22xp5_ASAP7_75t_SL g376 ( 
.A1(n_15),
.A2(n_47),
.B1(n_369),
.B2(n_377),
.Y(n_376)
);

XNOR2xp5_ASAP7_75t_L g16 ( 
.A(n_17),
.B(n_443),
.Y(n_16)
);

OA21x2_ASAP7_75t_L g17 ( 
.A1(n_18),
.A2(n_307),
.B(n_437),
.Y(n_17)
);

NAND3xp33_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_254),
.C(n_287),
.Y(n_18)
);

NOR2xp33_ASAP7_75t_SL g19 ( 
.A(n_20),
.B(n_238),
.Y(n_19)
);

OAI21xp5_ASAP7_75t_L g438 ( 
.A1(n_20),
.A2(n_439),
.B(n_440),
.Y(n_438)
);

NOR2xp33_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_199),
.Y(n_20)
);

NAND2xp5_ASAP7_75t_L g440 ( 
.A(n_21),
.B(n_199),
.Y(n_440)
);

MAJIxp5_ASAP7_75t_L g21 ( 
.A(n_22),
.B(n_135),
.C(n_183),
.Y(n_21)
);

XOR2xp5_ASAP7_75t_L g252 ( 
.A(n_22),
.B(n_253),
.Y(n_252)
);

XOR2xp5_ASAP7_75t_L g22 ( 
.A(n_23),
.B(n_72),
.Y(n_22)
);

MAJIxp5_ASAP7_75t_L g200 ( 
.A(n_23),
.B(n_73),
.C(n_103),
.Y(n_200)
);

NAND2xp5_ASAP7_75t_L g23 ( 
.A(n_24),
.B(n_46),
.Y(n_23)
);

XNOR2xp5_ASAP7_75t_L g241 ( 
.A(n_24),
.B(n_46),
.Y(n_241)
);

OAI32xp33_ASAP7_75t_L g24 ( 
.A1(n_25),
.A2(n_28),
.A3(n_31),
.B1(n_35),
.B2(n_41),
.Y(n_24)
);

INVx4_ASAP7_75t_L g25 ( 
.A(n_26),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_27),
.Y(n_26)
);

INVx6_ASAP7_75t_L g38 ( 
.A(n_27),
.Y(n_38)
);

INVx3_ASAP7_75t_L g89 ( 
.A(n_27),
.Y(n_89)
);

BUFx6f_ASAP7_75t_L g95 ( 
.A(n_27),
.Y(n_95)
);

BUFx5_ASAP7_75t_L g122 ( 
.A(n_27),
.Y(n_122)
);

INVx2_ASAP7_75t_L g230 ( 
.A(n_27),
.Y(n_230)
);

INVx1_ASAP7_75t_SL g28 ( 
.A(n_29),
.Y(n_28)
);

INVx8_ASAP7_75t_L g29 ( 
.A(n_30),
.Y(n_29)
);

INVx2_ASAP7_75t_L g459 ( 
.A(n_30),
.Y(n_459)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_32),
.Y(n_31)
);

INVx6_ASAP7_75t_L g32 ( 
.A(n_33),
.Y(n_32)
);

OAI22xp5_ASAP7_75t_L g120 ( 
.A1(n_33),
.A2(n_121),
.B1(n_123),
.B2(n_125),
.Y(n_120)
);

INVx5_ASAP7_75t_L g33 ( 
.A(n_34),
.Y(n_33)
);

INVx3_ASAP7_75t_L g40 ( 
.A(n_34),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_SL g35 ( 
.A(n_36),
.B(n_39),
.Y(n_35)
);

INVx2_ASAP7_75t_L g36 ( 
.A(n_37),
.Y(n_36)
);

OAI22xp5_ASAP7_75t_SL g87 ( 
.A1(n_37),
.A2(n_88),
.B1(n_90),
.B2(n_91),
.Y(n_87)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_38),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g177 ( 
.A(n_38),
.Y(n_177)
);

BUFx6f_ASAP7_75t_L g180 ( 
.A(n_38),
.Y(n_180)
);

BUFx6f_ASAP7_75t_L g274 ( 
.A(n_38),
.Y(n_274)
);

BUFx6f_ASAP7_75t_L g399 ( 
.A(n_38),
.Y(n_399)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_40),
.Y(n_39)
);

INVxp33_ASAP7_75t_L g41 ( 
.A(n_42),
.Y(n_41)
);

INVx3_ASAP7_75t_L g43 ( 
.A(n_44),
.Y(n_43)
);

INVx2_ASAP7_75t_L g44 ( 
.A(n_45),
.Y(n_44)
);

INVx2_ASAP7_75t_L g235 ( 
.A(n_45),
.Y(n_235)
);

OAI22xp5_ASAP7_75t_L g46 ( 
.A1(n_47),
.A2(n_56),
.B1(n_65),
.B2(n_67),
.Y(n_46)
);

OAI21xp5_ASAP7_75t_L g184 ( 
.A1(n_47),
.A2(n_67),
.B(n_185),
.Y(n_184)
);

NOR2xp33_ASAP7_75t_L g212 ( 
.A(n_47),
.B(n_187),
.Y(n_212)
);

AOI21xp5_ASAP7_75t_L g261 ( 
.A1(n_47),
.A2(n_215),
.B(n_262),
.Y(n_261)
);

OAI21xp5_ASAP7_75t_L g348 ( 
.A1(n_47),
.A2(n_213),
.B(n_349),
.Y(n_348)
);

INVxp67_ASAP7_75t_L g361 ( 
.A(n_47),
.Y(n_361)
);

OAI22xp5_ASAP7_75t_SL g368 ( 
.A1(n_47),
.A2(n_359),
.B1(n_369),
.B2(n_373),
.Y(n_368)
);

OAI21xp5_ASAP7_75t_L g407 ( 
.A1(n_47),
.A2(n_185),
.B(n_215),
.Y(n_407)
);

OR2x2_ASAP7_75t_L g47 ( 
.A(n_48),
.B(n_53),
.Y(n_47)
);

INVx1_ASAP7_75t_L g360 ( 
.A(n_48),
.Y(n_360)
);

INVx6_ASAP7_75t_L g48 ( 
.A(n_49),
.Y(n_48)
);

INVx4_ASAP7_75t_L g49 ( 
.A(n_50),
.Y(n_49)
);

INVx4_ASAP7_75t_L g371 ( 
.A(n_50),
.Y(n_371)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_51),
.Y(n_50)
);

BUFx3_ASAP7_75t_L g51 ( 
.A(n_52),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g71 ( 
.A(n_52),
.Y(n_71)
);

BUFx6f_ASAP7_75t_L g351 ( 
.A(n_52),
.Y(n_351)
);

NAND2xp5_ASAP7_75t_L g185 ( 
.A(n_53),
.B(n_186),
.Y(n_185)
);

AOI21xp5_ASAP7_75t_L g244 ( 
.A1(n_53),
.A2(n_57),
.B(n_212),
.Y(n_244)
);

INVx3_ASAP7_75t_SL g53 ( 
.A(n_54),
.Y(n_53)
);

INVx4_ASAP7_75t_L g54 ( 
.A(n_55),
.Y(n_54)
);

INVx1_ASAP7_75t_L g381 ( 
.A(n_55),
.Y(n_381)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_57),
.Y(n_56)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_59),
.Y(n_58)
);

INVx8_ASAP7_75t_L g59 ( 
.A(n_60),
.Y(n_59)
);

BUFx2_ASAP7_75t_L g64 ( 
.A(n_60),
.Y(n_64)
);

AOI22xp5_ASAP7_75t_L g154 ( 
.A1(n_60),
.A2(n_155),
.B1(n_158),
.B2(n_160),
.Y(n_154)
);

BUFx8_ASAP7_75t_L g60 ( 
.A(n_61),
.Y(n_60)
);

BUFx3_ASAP7_75t_L g159 ( 
.A(n_61),
.Y(n_159)
);

BUFx5_ASAP7_75t_L g354 ( 
.A(n_61),
.Y(n_354)
);

INVx2_ASAP7_75t_L g385 ( 
.A(n_61),
.Y(n_385)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_64),
.Y(n_63)
);

INVx3_ASAP7_75t_L g65 ( 
.A(n_66),
.Y(n_65)
);

INVx1_ASAP7_75t_SL g69 ( 
.A(n_70),
.Y(n_69)
);

BUFx6f_ASAP7_75t_L g70 ( 
.A(n_71),
.Y(n_70)
);

INVx2_ASAP7_75t_L g193 ( 
.A(n_71),
.Y(n_193)
);

INVx5_ASAP7_75t_L g326 ( 
.A(n_71),
.Y(n_326)
);

XOR2xp5_ASAP7_75t_L g72 ( 
.A(n_73),
.B(n_103),
.Y(n_72)
);

AOI21xp5_ASAP7_75t_L g73 ( 
.A1(n_74),
.A2(n_92),
.B(n_99),
.Y(n_73)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_74),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_SL g275 ( 
.A(n_74),
.B(n_227),
.Y(n_275)
);

AOI22xp5_ASAP7_75t_L g292 ( 
.A1(n_74),
.A2(n_226),
.B1(n_293),
.B2(n_294),
.Y(n_292)
);

AOI22xp5_ASAP7_75t_L g409 ( 
.A1(n_74),
.A2(n_226),
.B1(n_249),
.B2(n_410),
.Y(n_409)
);

AOI21xp5_ASAP7_75t_L g452 ( 
.A1(n_74),
.A2(n_294),
.B(n_453),
.Y(n_452)
);

AND2x2_ASAP7_75t_L g74 ( 
.A(n_75),
.B(n_87),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_75),
.B(n_100),
.Y(n_99)
);

OAI22xp5_ASAP7_75t_L g174 ( 
.A1(n_75),
.A2(n_175),
.B1(n_181),
.B2(n_182),
.Y(n_174)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_75),
.Y(n_226)
);

OAI22xp5_ASAP7_75t_SL g247 ( 
.A1(n_75),
.A2(n_175),
.B1(n_181),
.B2(n_248),
.Y(n_247)
);

OAI21xp5_ASAP7_75t_L g271 ( 
.A1(n_75),
.A2(n_272),
.B(n_275),
.Y(n_271)
);

OA22x2_ASAP7_75t_L g75 ( 
.A1(n_76),
.A2(n_79),
.B1(n_82),
.B2(n_84),
.Y(n_75)
);

INVx3_ASAP7_75t_L g76 ( 
.A(n_77),
.Y(n_76)
);

INVx2_ASAP7_75t_L g167 ( 
.A(n_77),
.Y(n_167)
);

BUFx3_ASAP7_75t_L g77 ( 
.A(n_78),
.Y(n_77)
);

INVx11_ASAP7_75t_L g83 ( 
.A(n_78),
.Y(n_83)
);

INVx3_ASAP7_75t_L g145 ( 
.A(n_78),
.Y(n_145)
);

BUFx3_ASAP7_75t_L g153 ( 
.A(n_78),
.Y(n_153)
);

BUFx6f_ASAP7_75t_L g333 ( 
.A(n_78),
.Y(n_333)
);

INVx3_ASAP7_75t_L g345 ( 
.A(n_78),
.Y(n_345)
);

BUFx5_ASAP7_75t_L g346 ( 
.A(n_78),
.Y(n_346)
);

INVx2_ASAP7_75t_L g406 ( 
.A(n_78),
.Y(n_406)
);

INVx4_ASAP7_75t_L g79 ( 
.A(n_80),
.Y(n_79)
);

INVx3_ASAP7_75t_L g80 ( 
.A(n_81),
.Y(n_80)
);

INVx3_ASAP7_75t_L g86 ( 
.A(n_81),
.Y(n_86)
);

BUFx3_ASAP7_75t_L g91 ( 
.A(n_81),
.Y(n_91)
);

INVx3_ASAP7_75t_L g402 ( 
.A(n_81),
.Y(n_402)
);

INVx4_ASAP7_75t_L g140 ( 
.A(n_82),
.Y(n_140)
);

INVx5_ASAP7_75t_L g336 ( 
.A(n_82),
.Y(n_336)
);

INVx5_ASAP7_75t_L g82 ( 
.A(n_83),
.Y(n_82)
);

BUFx6f_ASAP7_75t_L g139 ( 
.A(n_83),
.Y(n_139)
);

BUFx6f_ASAP7_75t_L g170 ( 
.A(n_83),
.Y(n_170)
);

BUFx6f_ASAP7_75t_L g198 ( 
.A(n_83),
.Y(n_198)
);

INVx6_ASAP7_75t_L g317 ( 
.A(n_83),
.Y(n_317)
);

INVx6_ASAP7_75t_L g332 ( 
.A(n_83),
.Y(n_332)
);

BUFx6f_ASAP7_75t_L g415 ( 
.A(n_83),
.Y(n_415)
);

INVx3_ASAP7_75t_L g84 ( 
.A(n_85),
.Y(n_84)
);

INVx4_ASAP7_75t_L g85 ( 
.A(n_86),
.Y(n_85)
);

BUFx6f_ASAP7_75t_L g90 ( 
.A(n_86),
.Y(n_90)
);

INVx4_ASAP7_75t_L g88 ( 
.A(n_89),
.Y(n_88)
);

INVx4_ASAP7_75t_L g101 ( 
.A(n_89),
.Y(n_101)
);

INVx6_ASAP7_75t_L g396 ( 
.A(n_91),
.Y(n_396)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_92),
.Y(n_182)
);

INVx5_ASAP7_75t_L g93 ( 
.A(n_94),
.Y(n_93)
);

BUFx6f_ASAP7_75t_L g94 ( 
.A(n_95),
.Y(n_94)
);

INVx4_ASAP7_75t_L g98 ( 
.A(n_95),
.Y(n_98)
);

INVx3_ASAP7_75t_L g126 ( 
.A(n_95),
.Y(n_126)
);

INVx3_ASAP7_75t_L g97 ( 
.A(n_98),
.Y(n_97)
);

OAI21xp5_ASAP7_75t_L g224 ( 
.A1(n_100),
.A2(n_181),
.B(n_225),
.Y(n_224)
);

AOI22xp5_ASAP7_75t_L g103 ( 
.A1(n_104),
.A2(n_109),
.B1(n_127),
.B2(n_133),
.Y(n_103)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_104),
.Y(n_173)
);

INVx3_ASAP7_75t_L g105 ( 
.A(n_106),
.Y(n_105)
);

INVx8_ASAP7_75t_L g106 ( 
.A(n_107),
.Y(n_106)
);

AOI21xp5_ASAP7_75t_L g303 ( 
.A1(n_109),
.A2(n_279),
.B(n_304),
.Y(n_303)
);

NAND2xp5_ASAP7_75t_L g460 ( 
.A(n_109),
.B(n_461),
.Y(n_460)
);

INVx1_ASAP7_75t_SL g109 ( 
.A(n_110),
.Y(n_109)
);

OAI22xp5_ASAP7_75t_L g171 ( 
.A1(n_110),
.A2(n_134),
.B1(n_172),
.B2(n_173),
.Y(n_171)
);

OAI22xp5_ASAP7_75t_SL g231 ( 
.A1(n_110),
.A2(n_128),
.B1(n_134),
.B2(n_232),
.Y(n_231)
);

OAI21xp5_ASAP7_75t_SL g277 ( 
.A1(n_110),
.A2(n_232),
.B(n_278),
.Y(n_277)
);

OR2x2_ASAP7_75t_L g110 ( 
.A(n_111),
.B(n_120),
.Y(n_110)
);

AOI22xp33_ASAP7_75t_L g111 ( 
.A1(n_112),
.A2(n_114),
.B1(n_116),
.B2(n_118),
.Y(n_111)
);

INVx6_ASAP7_75t_L g112 ( 
.A(n_113),
.Y(n_112)
);

INVx6_ASAP7_75t_L g114 ( 
.A(n_115),
.Y(n_114)
);

INVx4_ASAP7_75t_L g116 ( 
.A(n_117),
.Y(n_116)
);

INVx3_ASAP7_75t_L g118 ( 
.A(n_119),
.Y(n_118)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_120),
.Y(n_134)
);

INVx5_ASAP7_75t_L g121 ( 
.A(n_122),
.Y(n_121)
);

INVx4_ASAP7_75t_L g123 ( 
.A(n_124),
.Y(n_123)
);

INVx4_ASAP7_75t_L g125 ( 
.A(n_126),
.Y(n_125)
);

INVxp67_ASAP7_75t_L g127 ( 
.A(n_128),
.Y(n_127)
);

INVx8_ASAP7_75t_L g130 ( 
.A(n_131),
.Y(n_130)
);

INVx8_ASAP7_75t_L g131 ( 
.A(n_132),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g278 ( 
.A(n_133),
.B(n_279),
.Y(n_278)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_134),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_L g304 ( 
.A(n_134),
.B(n_305),
.Y(n_304)
);

OAI21xp5_ASAP7_75t_L g456 ( 
.A1(n_134),
.A2(n_457),
.B(n_460),
.Y(n_456)
);

XNOR2xp5_ASAP7_75t_L g253 ( 
.A(n_135),
.B(n_183),
.Y(n_253)
);

MAJIxp5_ASAP7_75t_L g135 ( 
.A(n_136),
.B(n_171),
.C(n_174),
.Y(n_135)
);

FAx1_ASAP7_75t_SL g240 ( 
.A(n_136),
.B(n_171),
.CI(n_174),
.CON(n_240),
.SN(n_240)
);

OAI21xp5_ASAP7_75t_L g136 ( 
.A1(n_137),
.A2(n_141),
.B(n_161),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_L g297 ( 
.A(n_137),
.B(n_163),
.Y(n_297)
);

AOI21xp5_ASAP7_75t_L g451 ( 
.A1(n_137),
.A2(n_141),
.B(n_163),
.Y(n_451)
);

INVx2_ASAP7_75t_L g207 ( 
.A(n_138),
.Y(n_207)
);

INVx11_ASAP7_75t_L g138 ( 
.A(n_139),
.Y(n_138)
);

INVx3_ASAP7_75t_L g208 ( 
.A(n_140),
.Y(n_208)
);

OAI22xp5_ASAP7_75t_SL g194 ( 
.A1(n_141),
.A2(n_163),
.B1(n_195),
.B2(n_196),
.Y(n_194)
);

OAI21xp5_ASAP7_75t_L g265 ( 
.A1(n_141),
.A2(n_161),
.B(n_266),
.Y(n_265)
);

NOR2xp33_ASAP7_75t_SL g298 ( 
.A(n_141),
.B(n_195),
.Y(n_298)
);

OAI21xp5_ASAP7_75t_SL g426 ( 
.A1(n_141),
.A2(n_427),
.B(n_428),
.Y(n_426)
);

INVx2_ASAP7_75t_L g141 ( 
.A(n_142),
.Y(n_141)
);

AOI22xp5_ASAP7_75t_L g204 ( 
.A1(n_142),
.A2(n_162),
.B1(n_205),
.B2(n_206),
.Y(n_204)
);

AOI22xp5_ASAP7_75t_L g327 ( 
.A1(n_142),
.A2(n_162),
.B1(n_328),
.B2(n_334),
.Y(n_327)
);

AOI22xp5_ASAP7_75t_L g341 ( 
.A1(n_142),
.A2(n_162),
.B1(n_334),
.B2(n_342),
.Y(n_341)
);

AOI22xp5_ASAP7_75t_L g411 ( 
.A1(n_142),
.A2(n_162),
.B1(n_342),
.B2(n_412),
.Y(n_411)
);

AND2x2_ASAP7_75t_L g142 ( 
.A(n_143),
.B(n_154),
.Y(n_142)
);

OAI22xp33_ASAP7_75t_L g143 ( 
.A1(n_144),
.A2(n_146),
.B1(n_149),
.B2(n_152),
.Y(n_143)
);

INVx4_ASAP7_75t_L g144 ( 
.A(n_145),
.Y(n_144)
);

INVx3_ASAP7_75t_L g146 ( 
.A(n_147),
.Y(n_146)
);

BUFx6f_ASAP7_75t_L g147 ( 
.A(n_148),
.Y(n_147)
);

BUFx5_ASAP7_75t_L g160 ( 
.A(n_148),
.Y(n_160)
);

INVx4_ASAP7_75t_L g149 ( 
.A(n_150),
.Y(n_149)
);

INVx4_ASAP7_75t_L g150 ( 
.A(n_151),
.Y(n_150)
);

INVx5_ASAP7_75t_L g322 ( 
.A(n_151),
.Y(n_322)
);

INVx3_ASAP7_75t_L g152 ( 
.A(n_153),
.Y(n_152)
);

BUFx3_ASAP7_75t_L g163 ( 
.A(n_154),
.Y(n_163)
);

INVx2_ASAP7_75t_L g155 ( 
.A(n_156),
.Y(n_155)
);

INVx3_ASAP7_75t_L g156 ( 
.A(n_157),
.Y(n_156)
);

INVx5_ASAP7_75t_L g158 ( 
.A(n_159),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_L g161 ( 
.A(n_162),
.B(n_164),
.Y(n_161)
);

INVx2_ASAP7_75t_SL g162 ( 
.A(n_163),
.Y(n_162)
);

NOR2xp33_ASAP7_75t_L g367 ( 
.A(n_163),
.B(n_329),
.Y(n_367)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_164),
.Y(n_195)
);

INVx2_ASAP7_75t_L g165 ( 
.A(n_166),
.Y(n_165)
);

INVx2_ASAP7_75t_L g166 ( 
.A(n_167),
.Y(n_166)
);

INVx4_ASAP7_75t_L g169 ( 
.A(n_170),
.Y(n_169)
);

INVx2_ASAP7_75t_L g395 ( 
.A(n_170),
.Y(n_395)
);

INVx6_ASAP7_75t_L g295 ( 
.A(n_176),
.Y(n_295)
);

INVx6_ASAP7_75t_L g176 ( 
.A(n_177),
.Y(n_176)
);

INVx2_ASAP7_75t_L g178 ( 
.A(n_179),
.Y(n_178)
);

INVx4_ASAP7_75t_L g179 ( 
.A(n_180),
.Y(n_179)
);

INVx3_ASAP7_75t_L g251 ( 
.A(n_180),
.Y(n_251)
);

XNOR2xp5_ASAP7_75t_L g183 ( 
.A(n_184),
.B(n_194),
.Y(n_183)
);

AND2x2_ASAP7_75t_L g237 ( 
.A(n_184),
.B(n_194),
.Y(n_237)
);

INVxp67_ASAP7_75t_L g186 ( 
.A(n_187),
.Y(n_186)
);

INVx3_ASAP7_75t_L g188 ( 
.A(n_189),
.Y(n_188)
);

BUFx6f_ASAP7_75t_L g189 ( 
.A(n_190),
.Y(n_189)
);

INVx2_ASAP7_75t_L g218 ( 
.A(n_190),
.Y(n_218)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_192),
.Y(n_191)
);

INVx4_ASAP7_75t_L g192 ( 
.A(n_193),
.Y(n_192)
);

INVxp67_ASAP7_75t_L g205 ( 
.A(n_196),
.Y(n_205)
);

INVx4_ASAP7_75t_L g197 ( 
.A(n_198),
.Y(n_197)
);

XNOR2xp5_ASAP7_75t_L g199 ( 
.A(n_200),
.B(n_201),
.Y(n_199)
);

MAJIxp5_ASAP7_75t_L g286 ( 
.A(n_200),
.B(n_202),
.C(n_221),
.Y(n_286)
);

XNOR2xp5_ASAP7_75t_L g201 ( 
.A(n_202),
.B(n_221),
.Y(n_201)
);

OAI22xp5_ASAP7_75t_SL g202 ( 
.A1(n_203),
.A2(n_204),
.B1(n_209),
.B2(n_210),
.Y(n_202)
);

NAND2xp5_ASAP7_75t_L g269 ( 
.A(n_203),
.B(n_210),
.Y(n_269)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_204),
.Y(n_203)
);

INVxp67_ASAP7_75t_L g266 ( 
.A(n_206),
.Y(n_266)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_210),
.Y(n_209)
);

NAND2xp5_ASAP7_75t_L g210 ( 
.A(n_211),
.B(n_213),
.Y(n_210)
);

INVxp67_ASAP7_75t_L g211 ( 
.A(n_212),
.Y(n_211)
);

NAND2xp5_ASAP7_75t_SL g213 ( 
.A(n_214),
.B(n_219),
.Y(n_213)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_215),
.Y(n_214)
);

INVx2_ASAP7_75t_L g216 ( 
.A(n_217),
.Y(n_216)
);

INVx6_ASAP7_75t_L g217 ( 
.A(n_218),
.Y(n_217)
);

INVx2_ASAP7_75t_L g219 ( 
.A(n_220),
.Y(n_219)
);

BUFx6f_ASAP7_75t_L g264 ( 
.A(n_220),
.Y(n_264)
);

XNOR2xp5_ASAP7_75t_L g221 ( 
.A(n_222),
.B(n_237),
.Y(n_221)
);

AOI22xp5_ASAP7_75t_SL g222 ( 
.A1(n_223),
.A2(n_224),
.B1(n_231),
.B2(n_236),
.Y(n_222)
);

MAJIxp5_ASAP7_75t_L g256 ( 
.A(n_223),
.B(n_236),
.C(n_257),
.Y(n_256)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_224),
.Y(n_223)
);

INVxp67_ASAP7_75t_L g453 ( 
.A(n_225),
.Y(n_453)
);

NAND2xp5_ASAP7_75t_L g225 ( 
.A(n_226),
.B(n_227),
.Y(n_225)
);

INVx2_ASAP7_75t_L g228 ( 
.A(n_229),
.Y(n_228)
);

OAI32xp33_ASAP7_75t_L g393 ( 
.A1(n_229),
.A2(n_394),
.A3(n_396),
.B1(n_397),
.B2(n_400),
.Y(n_393)
);

INVx6_ASAP7_75t_L g229 ( 
.A(n_230),
.Y(n_229)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_231),
.Y(n_236)
);

INVx2_ASAP7_75t_L g233 ( 
.A(n_234),
.Y(n_233)
);

INVx4_ASAP7_75t_L g282 ( 
.A(n_235),
.Y(n_282)
);

INVxp67_ASAP7_75t_L g257 ( 
.A(n_237),
.Y(n_257)
);

NOR2xp33_ASAP7_75t_L g238 ( 
.A(n_239),
.B(n_252),
.Y(n_238)
);

NAND2xp5_ASAP7_75t_L g439 ( 
.A(n_239),
.B(n_252),
.Y(n_439)
);

MAJIxp5_ASAP7_75t_L g239 ( 
.A(n_240),
.B(n_241),
.C(n_242),
.Y(n_239)
);

XNOR2xp5_ASAP7_75t_L g434 ( 
.A(n_240),
.B(n_435),
.Y(n_434)
);

BUFx24_ASAP7_75t_SL g466 ( 
.A(n_240),
.Y(n_466)
);

XNOR2xp5_ASAP7_75t_L g435 ( 
.A(n_241),
.B(n_242),
.Y(n_435)
);

MAJIxp5_ASAP7_75t_L g242 ( 
.A(n_243),
.B(n_245),
.C(n_247),
.Y(n_242)
);

OAI22xp5_ASAP7_75t_SL g422 ( 
.A1(n_243),
.A2(n_244),
.B1(n_245),
.B2(n_246),
.Y(n_422)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_244),
.Y(n_243)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_246),
.Y(n_245)
);

XNOR2xp5_ASAP7_75t_SL g421 ( 
.A(n_247),
.B(n_422),
.Y(n_421)
);

INVxp67_ASAP7_75t_L g248 ( 
.A(n_249),
.Y(n_248)
);

INVx5_ASAP7_75t_L g250 ( 
.A(n_251),
.Y(n_250)
);

A2O1A1O1Ixp25_ASAP7_75t_L g437 ( 
.A1(n_254),
.A2(n_287),
.B(n_438),
.C(n_441),
.D(n_442),
.Y(n_437)
);

NAND2xp5_ASAP7_75t_SL g254 ( 
.A(n_255),
.B(n_286),
.Y(n_254)
);

NOR2xp33_ASAP7_75t_L g441 ( 
.A(n_255),
.B(n_286),
.Y(n_441)
);

XOR2xp5_ASAP7_75t_L g255 ( 
.A(n_256),
.B(n_258),
.Y(n_255)
);

MAJIxp5_ASAP7_75t_L g288 ( 
.A(n_256),
.B(n_259),
.C(n_285),
.Y(n_288)
);

AOI22xp5_ASAP7_75t_L g258 ( 
.A1(n_259),
.A2(n_268),
.B1(n_284),
.B2(n_285),
.Y(n_258)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_259),
.Y(n_284)
);

OAI22xp5_ASAP7_75t_L g259 ( 
.A1(n_260),
.A2(n_261),
.B1(n_265),
.B2(n_267),
.Y(n_259)
);

AOI22xp5_ASAP7_75t_L g302 ( 
.A1(n_260),
.A2(n_261),
.B1(n_303),
.B2(n_306),
.Y(n_302)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_261),
.Y(n_260)
);

NAND2xp5_ASAP7_75t_L g301 ( 
.A(n_261),
.B(n_265),
.Y(n_301)
);

AOI21xp33_ASAP7_75t_L g463 ( 
.A1(n_261),
.A2(n_301),
.B(n_303),
.Y(n_463)
);

INVx1_ASAP7_75t_L g363 ( 
.A(n_262),
.Y(n_363)
);

INVx2_ASAP7_75t_L g262 ( 
.A(n_263),
.Y(n_262)
);

INVx8_ASAP7_75t_L g263 ( 
.A(n_264),
.Y(n_263)
);

INVxp67_ASAP7_75t_L g267 ( 
.A(n_265),
.Y(n_267)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_268),
.Y(n_285)
);

XOR2xp5_ASAP7_75t_L g268 ( 
.A(n_269),
.B(n_270),
.Y(n_268)
);

MAJIxp5_ASAP7_75t_L g290 ( 
.A(n_269),
.B(n_276),
.C(n_283),
.Y(n_290)
);

OAI22xp5_ASAP7_75t_SL g270 ( 
.A1(n_271),
.A2(n_276),
.B1(n_277),
.B2(n_283),
.Y(n_270)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_271),
.Y(n_283)
);

INVxp67_ASAP7_75t_L g293 ( 
.A(n_272),
.Y(n_293)
);

INVx3_ASAP7_75t_L g273 ( 
.A(n_274),
.Y(n_273)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_277),
.Y(n_276)
);

INVx3_ASAP7_75t_L g280 ( 
.A(n_281),
.Y(n_280)
);

NAND2xp5_ASAP7_75t_L g287 ( 
.A(n_288),
.B(n_289),
.Y(n_287)
);

NOR2xp33_ASAP7_75t_L g442 ( 
.A(n_288),
.B(n_289),
.Y(n_442)
);

BUFx24_ASAP7_75t_SL g467 ( 
.A(n_289),
.Y(n_467)
);

FAx1_ASAP7_75t_SL g289 ( 
.A(n_290),
.B(n_291),
.CI(n_300),
.CON(n_289),
.SN(n_289)
);

MAJIxp5_ASAP7_75t_L g446 ( 
.A(n_290),
.B(n_291),
.C(n_300),
.Y(n_446)
);

OAI21xp5_ASAP7_75t_L g291 ( 
.A1(n_292),
.A2(n_296),
.B(n_299),
.Y(n_291)
);

NAND2xp5_ASAP7_75t_SL g299 ( 
.A(n_292),
.B(n_296),
.Y(n_299)
);

OAI21xp33_ASAP7_75t_SL g410 ( 
.A1(n_295),
.A2(n_329),
.B(n_397),
.Y(n_410)
);

NOR2xp33_ASAP7_75t_L g296 ( 
.A(n_297),
.B(n_298),
.Y(n_296)
);

INVxp67_ASAP7_75t_L g428 ( 
.A(n_297),
.Y(n_428)
);

FAx1_ASAP7_75t_SL g447 ( 
.A(n_299),
.B(n_448),
.CI(n_463),
.CON(n_447),
.SN(n_447)
);

XOR2xp5_ASAP7_75t_L g300 ( 
.A(n_301),
.B(n_302),
.Y(n_300)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_303),
.Y(n_306)
);

INVxp67_ASAP7_75t_L g461 ( 
.A(n_305),
.Y(n_461)
);

AOI21xp5_ASAP7_75t_L g307 ( 
.A1(n_308),
.A2(n_432),
.B(n_436),
.Y(n_307)
);

OAI21xp5_ASAP7_75t_SL g308 ( 
.A1(n_309),
.A2(n_417),
.B(n_431),
.Y(n_308)
);

AOI21xp5_ASAP7_75t_L g309 ( 
.A1(n_310),
.A2(n_389),
.B(n_416),
.Y(n_309)
);

OAI21xp5_ASAP7_75t_SL g310 ( 
.A1(n_311),
.A2(n_355),
.B(n_388),
.Y(n_310)
);

NOR2xp33_ASAP7_75t_L g311 ( 
.A(n_312),
.B(n_337),
.Y(n_311)
);

NAND2xp5_ASAP7_75t_L g388 ( 
.A(n_312),
.B(n_337),
.Y(n_388)
);

NOR2xp33_ASAP7_75t_L g312 ( 
.A(n_313),
.B(n_327),
.Y(n_312)
);

XNOR2xp5_ASAP7_75t_L g364 ( 
.A(n_313),
.B(n_327),
.Y(n_364)
);

NAND2xp5_ASAP7_75t_L g313 ( 
.A(n_314),
.B(n_318),
.Y(n_313)
);

INVx2_ASAP7_75t_L g314 ( 
.A(n_315),
.Y(n_314)
);

INVx2_ASAP7_75t_L g315 ( 
.A(n_316),
.Y(n_315)
);

INVx2_ASAP7_75t_L g316 ( 
.A(n_317),
.Y(n_316)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_320),
.Y(n_319)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_321),
.Y(n_320)
);

BUFx6f_ASAP7_75t_L g321 ( 
.A(n_322),
.Y(n_321)
);

INVx2_ASAP7_75t_L g323 ( 
.A(n_324),
.Y(n_323)
);

INVx3_ASAP7_75t_L g324 ( 
.A(n_325),
.Y(n_324)
);

BUFx6f_ASAP7_75t_L g325 ( 
.A(n_326),
.Y(n_325)
);

NOR2xp33_ASAP7_75t_L g380 ( 
.A(n_329),
.B(n_381),
.Y(n_380)
);

NAND2xp5_ASAP7_75t_L g397 ( 
.A(n_329),
.B(n_398),
.Y(n_397)
);

BUFx2_ASAP7_75t_L g330 ( 
.A(n_331),
.Y(n_330)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_332),
.Y(n_331)
);

INVx2_ASAP7_75t_L g335 ( 
.A(n_336),
.Y(n_335)
);

XNOR2xp5_ASAP7_75t_L g337 ( 
.A(n_338),
.B(n_348),
.Y(n_337)
);

AOI22xp5_ASAP7_75t_L g338 ( 
.A1(n_339),
.A2(n_340),
.B1(n_341),
.B2(n_347),
.Y(n_338)
);

MAJIxp5_ASAP7_75t_L g390 ( 
.A(n_339),
.B(n_347),
.C(n_348),
.Y(n_390)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_340),
.Y(n_339)
);

INVx1_ASAP7_75t_SL g347 ( 
.A(n_341),
.Y(n_347)
);

INVx4_ASAP7_75t_SL g343 ( 
.A(n_344),
.Y(n_343)
);

INVx2_ASAP7_75t_L g344 ( 
.A(n_345),
.Y(n_344)
);

INVxp67_ASAP7_75t_L g362 ( 
.A(n_349),
.Y(n_362)
);

HB1xp67_ASAP7_75t_L g350 ( 
.A(n_351),
.Y(n_350)
);

INVx8_ASAP7_75t_L g372 ( 
.A(n_351),
.Y(n_372)
);

CKINVDCx14_ASAP7_75t_R g352 ( 
.A(n_353),
.Y(n_352)
);

INVx2_ASAP7_75t_L g353 ( 
.A(n_354),
.Y(n_353)
);

AOI21xp5_ASAP7_75t_L g355 ( 
.A1(n_356),
.A2(n_365),
.B(n_387),
.Y(n_355)
);

NAND2xp5_ASAP7_75t_L g356 ( 
.A(n_357),
.B(n_364),
.Y(n_356)
);

NOR2xp33_ASAP7_75t_L g387 ( 
.A(n_357),
.B(n_364),
.Y(n_387)
);

AOI22xp5_ASAP7_75t_SL g357 ( 
.A1(n_358),
.A2(n_361),
.B1(n_362),
.B2(n_363),
.Y(n_357)
);

INVxp67_ASAP7_75t_L g358 ( 
.A(n_359),
.Y(n_358)
);

OAI21xp5_ASAP7_75t_SL g365 ( 
.A1(n_366),
.A2(n_375),
.B(n_386),
.Y(n_365)
);

NOR2xp33_ASAP7_75t_L g366 ( 
.A(n_367),
.B(n_368),
.Y(n_366)
);

NAND2xp5_ASAP7_75t_SL g386 ( 
.A(n_367),
.B(n_368),
.Y(n_386)
);

INVx2_ASAP7_75t_L g370 ( 
.A(n_371),
.Y(n_370)
);

INVx4_ASAP7_75t_L g378 ( 
.A(n_373),
.Y(n_378)
);

INVx4_ASAP7_75t_L g373 ( 
.A(n_374),
.Y(n_373)
);

NAND2xp5_ASAP7_75t_SL g375 ( 
.A(n_376),
.B(n_379),
.Y(n_375)
);

INVx1_ASAP7_75t_SL g377 ( 
.A(n_378),
.Y(n_377)
);

NOR2xp33_ASAP7_75t_SL g379 ( 
.A(n_380),
.B(n_382),
.Y(n_379)
);

INVx1_ASAP7_75t_L g382 ( 
.A(n_383),
.Y(n_382)
);

BUFx3_ASAP7_75t_L g383 ( 
.A(n_384),
.Y(n_383)
);

INVx1_ASAP7_75t_L g384 ( 
.A(n_385),
.Y(n_384)
);

NAND2xp5_ASAP7_75t_L g389 ( 
.A(n_390),
.B(n_391),
.Y(n_389)
);

NOR2xp33_ASAP7_75t_L g416 ( 
.A(n_390),
.B(n_391),
.Y(n_416)
);

XNOR2xp5_ASAP7_75t_L g391 ( 
.A(n_392),
.B(n_408),
.Y(n_391)
);

MAJIxp5_ASAP7_75t_L g418 ( 
.A(n_392),
.B(n_409),
.C(n_411),
.Y(n_418)
);

XNOR2xp5_ASAP7_75t_SL g392 ( 
.A(n_393),
.B(n_407),
.Y(n_392)
);

NAND2xp5_ASAP7_75t_L g425 ( 
.A(n_393),
.B(n_407),
.Y(n_425)
);

INVx1_ASAP7_75t_L g394 ( 
.A(n_395),
.Y(n_394)
);

BUFx6f_ASAP7_75t_L g398 ( 
.A(n_399),
.Y(n_398)
);

NOR2xp33_ASAP7_75t_L g400 ( 
.A(n_401),
.B(n_403),
.Y(n_400)
);

INVx6_ASAP7_75t_L g401 ( 
.A(n_402),
.Y(n_401)
);

INVx1_ASAP7_75t_L g403 ( 
.A(n_404),
.Y(n_403)
);

INVx2_ASAP7_75t_L g404 ( 
.A(n_405),
.Y(n_404)
);

INVx4_ASAP7_75t_L g413 ( 
.A(n_405),
.Y(n_413)
);

INVx4_ASAP7_75t_L g405 ( 
.A(n_406),
.Y(n_405)
);

XNOR2xp5_ASAP7_75t_L g408 ( 
.A(n_409),
.B(n_411),
.Y(n_408)
);

INVxp67_ASAP7_75t_L g427 ( 
.A(n_412),
.Y(n_427)
);

INVx2_ASAP7_75t_L g414 ( 
.A(n_415),
.Y(n_414)
);

NOR2xp33_ASAP7_75t_L g417 ( 
.A(n_418),
.B(n_419),
.Y(n_417)
);

NAND2xp5_ASAP7_75t_SL g431 ( 
.A(n_418),
.B(n_419),
.Y(n_431)
);

OAI22xp5_ASAP7_75t_SL g419 ( 
.A1(n_420),
.A2(n_421),
.B1(n_423),
.B2(n_424),
.Y(n_419)
);

MAJIxp5_ASAP7_75t_L g433 ( 
.A(n_420),
.B(n_426),
.C(n_429),
.Y(n_433)
);

INVx1_ASAP7_75t_L g420 ( 
.A(n_421),
.Y(n_420)
);

INVx1_ASAP7_75t_L g423 ( 
.A(n_424),
.Y(n_423)
);

OAI22xp5_ASAP7_75t_SL g424 ( 
.A1(n_425),
.A2(n_426),
.B1(n_429),
.B2(n_430),
.Y(n_424)
);

INVx1_ASAP7_75t_L g429 ( 
.A(n_425),
.Y(n_429)
);

INVx1_ASAP7_75t_L g430 ( 
.A(n_426),
.Y(n_430)
);

NAND2xp5_ASAP7_75t_L g432 ( 
.A(n_433),
.B(n_434),
.Y(n_432)
);

NOR2xp33_ASAP7_75t_L g436 ( 
.A(n_433),
.B(n_434),
.Y(n_436)
);

NAND2xp5_ASAP7_75t_L g443 ( 
.A(n_444),
.B(n_464),
.Y(n_443)
);

INVxp67_ASAP7_75t_L g444 ( 
.A(n_445),
.Y(n_444)
);

AND2x2_ASAP7_75t_L g445 ( 
.A(n_446),
.B(n_447),
.Y(n_445)
);

NOR2xp33_ASAP7_75t_L g465 ( 
.A(n_446),
.B(n_447),
.Y(n_465)
);

BUFx24_ASAP7_75t_SL g469 ( 
.A(n_447),
.Y(n_469)
);

OAI22xp5_ASAP7_75t_SL g448 ( 
.A1(n_449),
.A2(n_450),
.B1(n_456),
.B2(n_462),
.Y(n_448)
);

INVx1_ASAP7_75t_L g449 ( 
.A(n_450),
.Y(n_449)
);

AOI22xp5_ASAP7_75t_L g450 ( 
.A1(n_451),
.A2(n_452),
.B1(n_454),
.B2(n_455),
.Y(n_450)
);

INVx1_ASAP7_75t_L g455 ( 
.A(n_451),
.Y(n_455)
);

INVx1_ASAP7_75t_L g454 ( 
.A(n_452),
.Y(n_454)
);

INVx1_ASAP7_75t_L g462 ( 
.A(n_456),
.Y(n_462)
);

INVx2_ASAP7_75t_L g458 ( 
.A(n_459),
.Y(n_458)
);

INVx1_ASAP7_75t_L g464 ( 
.A(n_465),
.Y(n_464)
);


endmodule