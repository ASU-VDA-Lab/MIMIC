module fake_jpeg_2328_n_660 (n_13, n_1, n_10, n_6, n_14, n_19, n_18, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_660);

input n_13;
input n_1;
input n_10;
input n_6;
input n_14;
input n_19;
input n_18;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_660;

wire n_529;
wire n_595;
wire n_390;
wire n_552;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_252;
wire n_182;
wire n_525;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_586;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_657;
wire n_27;
wire n_365;
wire n_179;
wire n_620;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_611;
wire n_44;
wire n_355;
wire n_519;
wire n_276;
wire n_143;
wire n_431;
wire n_102;
wire n_549;
wire n_196;
wire n_66;
wire n_374;
wire n_566;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_597;
wire n_172;
wire n_547;
wire n_345;
wire n_591;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_513;
wire n_283;
wire n_107;
wire n_490;
wire n_635;
wire n_517;
wire n_629;
wire n_479;
wire n_415;
wire n_543;
wire n_357;
wire n_89;
wire n_131;
wire n_607;
wire n_294;
wire n_230;
wire n_643;
wire n_170;
wire n_602;
wire n_313;
wire n_542;
wire n_574;
wire n_264;
wire n_647;
wire n_437;
wire n_93;
wire n_227;
wire n_559;
wire n_641;
wire n_48;
wire n_465;
wire n_638;
wire n_200;
wire n_582;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_623;
wire n_579;
wire n_416;
wire n_256;
wire n_221;
wire n_454;
wire n_540;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_637;
wire n_370;
wire n_410;
wire n_571;
wire n_82;
wire n_155;
wire n_508;
wire n_309;
wire n_624;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_606;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_569;
wire n_596;
wire n_400;
wire n_646;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_544;
wire n_31;
wire n_277;
wire n_255;
wire n_605;
wire n_601;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_393;
wire n_349;
wire n_234;
wire n_530;
wire n_634;
wire n_23;
wire n_69;
wire n_658;
wire n_195;
wire n_450;
wire n_557;
wire n_408;
wire n_80;
wire n_562;
wire n_204;
wire n_639;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_645;
wire n_298;
wire n_106;
wire n_545;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_584;
wire n_254;
wire n_608;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_622;
wire n_463;
wire n_92;
wire n_332;
wire n_640;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_653;
wire n_474;
wire n_539;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_626;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_575;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_511;
wire n_305;
wire n_161;
wire n_441;
wire n_555;
wire n_342;
wire n_642;
wire n_101;
wire n_226;
wire n_509;
wire n_644;
wire n_149;
wire n_87;
wire n_46;
wire n_578;
wire n_656;
wire n_589;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_614;
wire n_97;
wire n_649;
wire n_573;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_610;
wire n_174;
wire n_198;
wire n_422;
wire n_560;
wire n_190;
wire n_510;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_536;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_537;
wire n_110;
wire n_594;
wire n_590;
wire n_531;
wire n_76;
wire n_278;
wire n_343;
wire n_577;
wire n_26;
wire n_88;
wire n_397;
wire n_592;
wire n_363;
wire n_570;
wire n_238;
wire n_598;
wire n_615;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_554;
wire n_301;
wire n_609;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_648;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_523;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_533;
wire n_612;
wire n_296;
wire n_384;
wire n_588;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_585;
wire n_491;
wire n_24;
wire n_526;
wire n_467;
wire n_269;
wire n_572;
wire n_546;
wire n_287;
wire n_219;
wire n_452;
wire n_631;
wire n_433;
wire n_636;
wire n_77;
wire n_473;
wire n_45;
wire n_520;
wire n_476;
wire n_337;
wire n_317;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_650;
wire n_218;
wire n_63;
wire n_652;
wire n_599;
wire n_239;
wire n_243;
wire n_481;
wire n_628;
wire n_619;
wire n_348;
wire n_587;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_583;
wire n_522;
wire n_333;
wire n_518;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_565;
wire n_302;
wire n_216;
wire n_528;
wire n_184;
wire n_655;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_199;
wire n_260;
wire n_550;
wire n_413;
wire n_275;
wire n_494;
wire n_604;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_551;
wire n_36;
wire n_62;
wire n_600;
wire n_492;
wire n_603;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_567;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_515;
wire n_347;
wire n_521;
wire n_424;
wire n_55;
wire n_358;
wire n_312;
wire n_47;
wire n_538;
wire n_625;
wire n_147;
wire n_449;
wire n_627;
wire n_98;
wire n_251;
wire n_534;
wire n_472;
wire n_279;
wire n_593;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_618;
wire n_356;
wire n_119;
wire n_484;
wire n_568;
wire n_83;
wire n_395;
wire n_659;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_576;
wire n_469;
wire n_111;
wire n_197;
wire n_396;
wire n_375;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_553;
wire n_257;
wire n_61;
wire n_173;
wire n_561;
wire n_244;
wire n_232;
wire n_527;
wire n_482;
wire n_58;
wire n_41;
wire n_613;
wire n_630;
wire n_266;
wire n_548;
wire n_72;
wire n_512;
wire n_654;
wire n_445;
wire n_443;
wire n_617;
wire n_215;
wire n_212;
wire n_516;
wire n_183;
wire n_409;
wire n_532;
wire n_249;
wire n_412;
wire n_581;
wire n_217;
wire n_471;
wire n_580;
wire n_541;
wire n_53;
wire n_372;
wire n_558;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_535;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_556;
wire n_524;
wire n_402;
wire n_563;
wire n_504;
wire n_438;
wire n_475;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_633;
wire n_112;
wire n_632;
wire n_616;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_514;
wire n_651;
wire n_564;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_621;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

INVx1_ASAP7_75t_L g20 ( 
.A(n_10),
.Y(n_20)
);

INVx13_ASAP7_75t_L g21 ( 
.A(n_18),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_12),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_2),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_15),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_16),
.Y(n_25)
);

BUFx10_ASAP7_75t_L g26 ( 
.A(n_8),
.Y(n_26)
);

INVx4_ASAP7_75t_L g27 ( 
.A(n_17),
.Y(n_27)
);

BUFx16f_ASAP7_75t_L g28 ( 
.A(n_19),
.Y(n_28)
);

BUFx12f_ASAP7_75t_L g29 ( 
.A(n_11),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_5),
.Y(n_30)
);

INVx2_ASAP7_75t_L g31 ( 
.A(n_2),
.Y(n_31)
);

INVx5_ASAP7_75t_L g32 ( 
.A(n_17),
.Y(n_32)
);

INVx2_ASAP7_75t_L g33 ( 
.A(n_9),
.Y(n_33)
);

BUFx5_ASAP7_75t_L g34 ( 
.A(n_15),
.Y(n_34)
);

INVx2_ASAP7_75t_L g35 ( 
.A(n_12),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_9),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_15),
.Y(n_37)
);

BUFx3_ASAP7_75t_L g38 ( 
.A(n_9),
.Y(n_38)
);

INVx2_ASAP7_75t_L g39 ( 
.A(n_14),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_5),
.Y(n_40)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_5),
.Y(n_41)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_2),
.Y(n_42)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_17),
.Y(n_43)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_5),
.Y(n_44)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_7),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_0),
.Y(n_46)
);

BUFx16f_ASAP7_75t_L g47 ( 
.A(n_6),
.Y(n_47)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_14),
.Y(n_48)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_15),
.Y(n_49)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_17),
.Y(n_50)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_18),
.Y(n_51)
);

BUFx3_ASAP7_75t_L g52 ( 
.A(n_13),
.Y(n_52)
);

BUFx12f_ASAP7_75t_L g53 ( 
.A(n_12),
.Y(n_53)
);

INVx2_ASAP7_75t_L g54 ( 
.A(n_6),
.Y(n_54)
);

BUFx12_ASAP7_75t_L g55 ( 
.A(n_10),
.Y(n_55)
);

INVx6_ASAP7_75t_SL g56 ( 
.A(n_13),
.Y(n_56)
);

CKINVDCx20_ASAP7_75t_R g57 ( 
.A(n_19),
.Y(n_57)
);

CKINVDCx20_ASAP7_75t_R g58 ( 
.A(n_2),
.Y(n_58)
);

BUFx12f_ASAP7_75t_L g59 ( 
.A(n_11),
.Y(n_59)
);

BUFx3_ASAP7_75t_L g60 ( 
.A(n_32),
.Y(n_60)
);

BUFx3_ASAP7_75t_L g180 ( 
.A(n_60),
.Y(n_180)
);

INVx4_ASAP7_75t_SL g61 ( 
.A(n_56),
.Y(n_61)
);

INVx5_ASAP7_75t_SL g183 ( 
.A(n_61),
.Y(n_183)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_25),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g136 ( 
.A(n_62),
.Y(n_136)
);

INVx1_ASAP7_75t_SL g63 ( 
.A(n_21),
.Y(n_63)
);

AND2x2_ASAP7_75t_L g215 ( 
.A(n_63),
.B(n_80),
.Y(n_215)
);

INVx2_ASAP7_75t_L g64 ( 
.A(n_31),
.Y(n_64)
);

INVx2_ASAP7_75t_L g138 ( 
.A(n_64),
.Y(n_138)
);

INVx4_ASAP7_75t_L g65 ( 
.A(n_34),
.Y(n_65)
);

INVx2_ASAP7_75t_SL g148 ( 
.A(n_65),
.Y(n_148)
);

INVx4_ASAP7_75t_L g66 ( 
.A(n_34),
.Y(n_66)
);

INVx2_ASAP7_75t_SL g153 ( 
.A(n_66),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_L g67 ( 
.A(n_35),
.B(n_19),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_L g170 ( 
.A(n_67),
.B(n_88),
.Y(n_170)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_25),
.Y(n_68)
);

BUFx6f_ASAP7_75t_L g185 ( 
.A(n_68),
.Y(n_185)
);

BUFx3_ASAP7_75t_L g69 ( 
.A(n_32),
.Y(n_69)
);

BUFx2_ASAP7_75t_L g217 ( 
.A(n_69),
.Y(n_217)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_31),
.Y(n_70)
);

INVx2_ASAP7_75t_L g149 ( 
.A(n_70),
.Y(n_149)
);

BUFx6f_ASAP7_75t_L g71 ( 
.A(n_25),
.Y(n_71)
);

BUFx6f_ASAP7_75t_L g186 ( 
.A(n_71),
.Y(n_186)
);

BUFx6f_ASAP7_75t_L g72 ( 
.A(n_25),
.Y(n_72)
);

BUFx6f_ASAP7_75t_L g194 ( 
.A(n_72),
.Y(n_194)
);

BUFx6f_ASAP7_75t_L g73 ( 
.A(n_30),
.Y(n_73)
);

BUFx6f_ASAP7_75t_L g210 ( 
.A(n_73),
.Y(n_210)
);

INVx3_ASAP7_75t_L g74 ( 
.A(n_27),
.Y(n_74)
);

INVx4_ASAP7_75t_SL g144 ( 
.A(n_74),
.Y(n_144)
);

INVx5_ASAP7_75t_L g75 ( 
.A(n_56),
.Y(n_75)
);

BUFx2_ASAP7_75t_L g225 ( 
.A(n_75),
.Y(n_225)
);

INVx3_ASAP7_75t_L g76 ( 
.A(n_27),
.Y(n_76)
);

INVx2_ASAP7_75t_SL g158 ( 
.A(n_76),
.Y(n_158)
);

INVx8_ASAP7_75t_L g77 ( 
.A(n_56),
.Y(n_77)
);

INVx5_ASAP7_75t_L g141 ( 
.A(n_77),
.Y(n_141)
);

INVx2_ASAP7_75t_L g78 ( 
.A(n_31),
.Y(n_78)
);

INVx2_ASAP7_75t_L g154 ( 
.A(n_78),
.Y(n_154)
);

BUFx6f_ASAP7_75t_L g79 ( 
.A(n_30),
.Y(n_79)
);

BUFx6f_ASAP7_75t_L g219 ( 
.A(n_79),
.Y(n_219)
);

HAxp5_ASAP7_75t_SL g80 ( 
.A(n_28),
.B(n_0),
.CON(n_80),
.SN(n_80)
);

BUFx6f_ASAP7_75t_L g81 ( 
.A(n_30),
.Y(n_81)
);

INVx6_ASAP7_75t_L g152 ( 
.A(n_81),
.Y(n_152)
);

BUFx6f_ASAP7_75t_L g82 ( 
.A(n_30),
.Y(n_82)
);

INVx6_ASAP7_75t_L g195 ( 
.A(n_82),
.Y(n_195)
);

BUFx6f_ASAP7_75t_L g83 ( 
.A(n_46),
.Y(n_83)
);

INVx6_ASAP7_75t_L g196 ( 
.A(n_83),
.Y(n_196)
);

BUFx3_ASAP7_75t_L g84 ( 
.A(n_32),
.Y(n_84)
);

INVx5_ASAP7_75t_L g164 ( 
.A(n_84),
.Y(n_164)
);

INVx11_ASAP7_75t_L g85 ( 
.A(n_29),
.Y(n_85)
);

INVx11_ASAP7_75t_L g221 ( 
.A(n_85),
.Y(n_221)
);

INVx6_ASAP7_75t_L g86 ( 
.A(n_46),
.Y(n_86)
);

INVx8_ASAP7_75t_L g145 ( 
.A(n_86),
.Y(n_145)
);

BUFx6f_ASAP7_75t_L g87 ( 
.A(n_46),
.Y(n_87)
);

INVx8_ASAP7_75t_L g218 ( 
.A(n_87),
.Y(n_218)
);

NAND2xp5_ASAP7_75t_L g88 ( 
.A(n_35),
.B(n_19),
.Y(n_88)
);

BUFx6f_ASAP7_75t_L g89 ( 
.A(n_46),
.Y(n_89)
);

INVx3_ASAP7_75t_L g165 ( 
.A(n_89),
.Y(n_165)
);

INVx2_ASAP7_75t_L g90 ( 
.A(n_33),
.Y(n_90)
);

INVx2_ASAP7_75t_L g157 ( 
.A(n_90),
.Y(n_157)
);

INVx8_ASAP7_75t_L g91 ( 
.A(n_28),
.Y(n_91)
);

INVx3_ASAP7_75t_L g212 ( 
.A(n_91),
.Y(n_212)
);

BUFx3_ASAP7_75t_L g92 ( 
.A(n_38),
.Y(n_92)
);

INVx4_ASAP7_75t_L g206 ( 
.A(n_92),
.Y(n_206)
);

BUFx6f_ASAP7_75t_L g93 ( 
.A(n_38),
.Y(n_93)
);

INVx4_ASAP7_75t_L g211 ( 
.A(n_93),
.Y(n_211)
);

INVx3_ASAP7_75t_L g94 ( 
.A(n_27),
.Y(n_94)
);

INVx3_ASAP7_75t_L g146 ( 
.A(n_94),
.Y(n_146)
);

BUFx6f_ASAP7_75t_L g95 ( 
.A(n_38),
.Y(n_95)
);

INVx4_ASAP7_75t_L g214 ( 
.A(n_95),
.Y(n_214)
);

BUFx3_ASAP7_75t_L g96 ( 
.A(n_52),
.Y(n_96)
);

INVx4_ASAP7_75t_L g216 ( 
.A(n_96),
.Y(n_216)
);

INVx2_ASAP7_75t_L g97 ( 
.A(n_33),
.Y(n_97)
);

INVx2_ASAP7_75t_L g162 ( 
.A(n_97),
.Y(n_162)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_33),
.Y(n_98)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_98),
.Y(n_139)
);

BUFx10_ASAP7_75t_L g99 ( 
.A(n_28),
.Y(n_99)
);

CKINVDCx16_ASAP7_75t_R g143 ( 
.A(n_99),
.Y(n_143)
);

BUFx12f_ASAP7_75t_L g100 ( 
.A(n_55),
.Y(n_100)
);

INVx3_ASAP7_75t_L g150 ( 
.A(n_100),
.Y(n_150)
);

INVx2_ASAP7_75t_L g101 ( 
.A(n_39),
.Y(n_101)
);

INVx2_ASAP7_75t_L g177 ( 
.A(n_101),
.Y(n_177)
);

BUFx6f_ASAP7_75t_L g102 ( 
.A(n_52),
.Y(n_102)
);

INVx2_ASAP7_75t_L g182 ( 
.A(n_102),
.Y(n_182)
);

INVx2_ASAP7_75t_L g103 ( 
.A(n_39),
.Y(n_103)
);

INVx2_ASAP7_75t_L g191 ( 
.A(n_103),
.Y(n_191)
);

BUFx6f_ASAP7_75t_L g104 ( 
.A(n_52),
.Y(n_104)
);

INVx2_ASAP7_75t_L g199 ( 
.A(n_104),
.Y(n_199)
);

INVx3_ASAP7_75t_L g105 ( 
.A(n_28),
.Y(n_105)
);

INVx3_ASAP7_75t_L g160 ( 
.A(n_105),
.Y(n_160)
);

INVx8_ASAP7_75t_L g106 ( 
.A(n_47),
.Y(n_106)
);

INVx3_ASAP7_75t_L g161 ( 
.A(n_106),
.Y(n_161)
);

INVx8_ASAP7_75t_L g107 ( 
.A(n_29),
.Y(n_107)
);

INVx3_ASAP7_75t_L g169 ( 
.A(n_107),
.Y(n_169)
);

BUFx6f_ASAP7_75t_L g108 ( 
.A(n_39),
.Y(n_108)
);

INVx2_ASAP7_75t_L g201 ( 
.A(n_108),
.Y(n_201)
);

BUFx6f_ASAP7_75t_L g109 ( 
.A(n_54),
.Y(n_109)
);

INVx2_ASAP7_75t_L g207 ( 
.A(n_109),
.Y(n_207)
);

BUFx5_ASAP7_75t_L g110 ( 
.A(n_47),
.Y(n_110)
);

INVx5_ASAP7_75t_SL g213 ( 
.A(n_110),
.Y(n_213)
);

BUFx5_ASAP7_75t_L g111 ( 
.A(n_47),
.Y(n_111)
);

CKINVDCx16_ASAP7_75t_R g159 ( 
.A(n_111),
.Y(n_159)
);

INVx3_ASAP7_75t_L g112 ( 
.A(n_47),
.Y(n_112)
);

INVx3_ASAP7_75t_L g184 ( 
.A(n_112),
.Y(n_184)
);

BUFx12f_ASAP7_75t_L g113 ( 
.A(n_55),
.Y(n_113)
);

INVx3_ASAP7_75t_L g200 ( 
.A(n_113),
.Y(n_200)
);

INVx3_ASAP7_75t_L g114 ( 
.A(n_29),
.Y(n_114)
);

INVx3_ASAP7_75t_L g203 ( 
.A(n_114),
.Y(n_203)
);

INVx2_ASAP7_75t_L g115 ( 
.A(n_54),
.Y(n_115)
);

INVx2_ASAP7_75t_L g209 ( 
.A(n_115),
.Y(n_209)
);

INVx11_ASAP7_75t_L g116 ( 
.A(n_29),
.Y(n_116)
);

INVx3_ASAP7_75t_L g208 ( 
.A(n_116),
.Y(n_208)
);

INVx2_ASAP7_75t_L g117 ( 
.A(n_54),
.Y(n_117)
);

INVx2_ASAP7_75t_L g223 ( 
.A(n_117),
.Y(n_223)
);

BUFx6f_ASAP7_75t_L g118 ( 
.A(n_59),
.Y(n_118)
);

INVx3_ASAP7_75t_L g222 ( 
.A(n_118),
.Y(n_222)
);

BUFx6f_ASAP7_75t_L g119 ( 
.A(n_59),
.Y(n_119)
);

HB1xp67_ASAP7_75t_L g135 ( 
.A(n_119),
.Y(n_135)
);

BUFx6f_ASAP7_75t_L g120 ( 
.A(n_59),
.Y(n_120)
);

HB1xp67_ASAP7_75t_L g198 ( 
.A(n_120),
.Y(n_198)
);

AOI22xp5_ASAP7_75t_L g121 ( 
.A1(n_22),
.A2(n_9),
.B1(n_16),
.B2(n_14),
.Y(n_121)
);

OAI22xp5_ASAP7_75t_SL g179 ( 
.A1(n_121),
.A2(n_37),
.B1(n_48),
.B2(n_42),
.Y(n_179)
);

BUFx6f_ASAP7_75t_L g122 ( 
.A(n_59),
.Y(n_122)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_122),
.Y(n_147)
);

BUFx6f_ASAP7_75t_L g123 ( 
.A(n_59),
.Y(n_123)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_123),
.Y(n_155)
);

BUFx6f_ASAP7_75t_L g124 ( 
.A(n_29),
.Y(n_124)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_124),
.Y(n_156)
);

INVx3_ASAP7_75t_L g125 ( 
.A(n_53),
.Y(n_125)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_125),
.Y(n_163)
);

BUFx12_ASAP7_75t_L g126 ( 
.A(n_21),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_L g132 ( 
.A(n_126),
.B(n_43),
.Y(n_132)
);

BUFx6f_ASAP7_75t_L g127 ( 
.A(n_53),
.Y(n_127)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_127),
.Y(n_166)
);

INVx6_ASAP7_75t_L g128 ( 
.A(n_53),
.Y(n_128)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_128),
.Y(n_171)
);

BUFx6f_ASAP7_75t_L g129 ( 
.A(n_53),
.Y(n_129)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_129),
.Y(n_173)
);

INVx3_ASAP7_75t_SL g130 ( 
.A(n_26),
.Y(n_130)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_130),
.Y(n_188)
);

BUFx6f_ASAP7_75t_L g131 ( 
.A(n_53),
.Y(n_131)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_131),
.Y(n_202)
);

CKINVDCx16_ASAP7_75t_R g230 ( 
.A(n_132),
.Y(n_230)
);

AOI22xp33_ASAP7_75t_SL g133 ( 
.A1(n_61),
.A2(n_58),
.B1(n_50),
.B2(n_49),
.Y(n_133)
);

OA22x2_ASAP7_75t_L g241 ( 
.A1(n_133),
.A2(n_142),
.B1(n_178),
.B2(n_181),
.Y(n_241)
);

NOR2xp33_ASAP7_75t_L g134 ( 
.A(n_77),
.B(n_91),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_SL g236 ( 
.A(n_134),
.B(n_137),
.Y(n_236)
);

NOR2xp33_ASAP7_75t_L g137 ( 
.A(n_106),
.B(n_22),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_SL g140 ( 
.A(n_130),
.B(n_44),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_SL g260 ( 
.A(n_140),
.B(n_174),
.Y(n_260)
);

AOI22xp5_ASAP7_75t_SL g142 ( 
.A1(n_93),
.A2(n_44),
.B1(n_57),
.B2(n_51),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_L g151 ( 
.A(n_100),
.B(n_36),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_L g229 ( 
.A(n_151),
.B(n_168),
.Y(n_229)
);

AOI22xp33_ASAP7_75t_L g167 ( 
.A1(n_83),
.A2(n_58),
.B1(n_23),
.B2(n_42),
.Y(n_167)
);

OAI22xp5_ASAP7_75t_L g231 ( 
.A1(n_167),
.A2(n_172),
.B1(n_197),
.B2(n_204),
.Y(n_231)
);

NOR2xp33_ASAP7_75t_L g168 ( 
.A(n_113),
.B(n_57),
.Y(n_168)
);

OAI22xp5_ASAP7_75t_L g172 ( 
.A1(n_62),
.A2(n_36),
.B1(n_51),
.B2(n_37),
.Y(n_172)
);

NOR2xp33_ASAP7_75t_SL g174 ( 
.A(n_118),
.B(n_40),
.Y(n_174)
);

NOR2xp33_ASAP7_75t_SL g175 ( 
.A(n_131),
.B(n_40),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_SL g263 ( 
.A(n_175),
.B(n_4),
.Y(n_263)
);

NAND2xp5_ASAP7_75t_L g176 ( 
.A(n_108),
.B(n_20),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_L g243 ( 
.A(n_176),
.B(n_187),
.Y(n_243)
);

AOI22xp33_ASAP7_75t_SL g178 ( 
.A1(n_80),
.A2(n_20),
.B1(n_50),
.B2(n_49),
.Y(n_178)
);

AOI22xp5_ASAP7_75t_SL g275 ( 
.A1(n_179),
.A2(n_0),
.B1(n_1),
.B2(n_3),
.Y(n_275)
);

AOI22xp33_ASAP7_75t_SL g181 ( 
.A1(n_95),
.A2(n_41),
.B1(n_24),
.B2(n_45),
.Y(n_181)
);

NOR2xp33_ASAP7_75t_L g187 ( 
.A(n_119),
.B(n_48),
.Y(n_187)
);

AOI22xp33_ASAP7_75t_SL g189 ( 
.A1(n_102),
.A2(n_45),
.B1(n_43),
.B2(n_41),
.Y(n_189)
);

OA22x2_ASAP7_75t_L g250 ( 
.A1(n_189),
.A2(n_192),
.B1(n_193),
.B2(n_220),
.Y(n_250)
);

NAND2xp5_ASAP7_75t_L g190 ( 
.A(n_109),
.B(n_24),
.Y(n_190)
);

NAND2xp5_ASAP7_75t_L g259 ( 
.A(n_190),
.B(n_205),
.Y(n_259)
);

AOI22xp33_ASAP7_75t_SL g192 ( 
.A1(n_104),
.A2(n_23),
.B1(n_26),
.B2(n_21),
.Y(n_192)
);

AOI22xp5_ASAP7_75t_SL g193 ( 
.A1(n_120),
.A2(n_26),
.B1(n_34),
.B2(n_55),
.Y(n_193)
);

AOI22xp33_ASAP7_75t_L g197 ( 
.A1(n_87),
.A2(n_26),
.B1(n_1),
.B2(n_2),
.Y(n_197)
);

AOI22xp33_ASAP7_75t_L g204 ( 
.A1(n_89),
.A2(n_26),
.B1(n_1),
.B2(n_3),
.Y(n_204)
);

NAND2xp5_ASAP7_75t_L g205 ( 
.A(n_68),
.B(n_11),
.Y(n_205)
);

AOI22xp33_ASAP7_75t_SL g220 ( 
.A1(n_122),
.A2(n_26),
.B1(n_55),
.B2(n_11),
.Y(n_220)
);

AOI22xp33_ASAP7_75t_SL g224 ( 
.A1(n_123),
.A2(n_55),
.B1(n_10),
.B2(n_12),
.Y(n_224)
);

OA22x2_ASAP7_75t_L g258 ( 
.A1(n_224),
.A2(n_6),
.B1(n_13),
.B2(n_8),
.Y(n_258)
);

INVx8_ASAP7_75t_L g226 ( 
.A(n_136),
.Y(n_226)
);

INVx5_ASAP7_75t_L g355 ( 
.A(n_226),
.Y(n_355)
);

BUFx6f_ASAP7_75t_L g227 ( 
.A(n_136),
.Y(n_227)
);

BUFx6f_ASAP7_75t_L g334 ( 
.A(n_227),
.Y(n_334)
);

INVx4_ASAP7_75t_L g228 ( 
.A(n_164),
.Y(n_228)
);

INVx3_ASAP7_75t_L g320 ( 
.A(n_228),
.Y(n_320)
);

OAI22xp5_ASAP7_75t_L g232 ( 
.A1(n_170),
.A2(n_81),
.B1(n_72),
.B2(n_73),
.Y(n_232)
);

OAI22xp5_ASAP7_75t_L g315 ( 
.A1(n_232),
.A2(n_255),
.B1(n_257),
.B2(n_272),
.Y(n_315)
);

BUFx3_ASAP7_75t_L g233 ( 
.A(n_212),
.Y(n_233)
);

BUFx3_ASAP7_75t_L g307 ( 
.A(n_233),
.Y(n_307)
);

BUFx6f_ASAP7_75t_L g234 ( 
.A(n_185),
.Y(n_234)
);

BUFx6f_ASAP7_75t_L g349 ( 
.A(n_234),
.Y(n_349)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_139),
.Y(n_235)
);

INVx2_ASAP7_75t_SL g340 ( 
.A(n_235),
.Y(n_340)
);

BUFx12f_ASAP7_75t_L g237 ( 
.A(n_212),
.Y(n_237)
);

HB1xp67_ASAP7_75t_L g322 ( 
.A(n_237),
.Y(n_322)
);

AND2x2_ASAP7_75t_SL g238 ( 
.A(n_215),
.B(n_157),
.Y(n_238)
);

CKINVDCx14_ASAP7_75t_R g306 ( 
.A(n_238),
.Y(n_306)
);

INVx5_ASAP7_75t_L g239 ( 
.A(n_141),
.Y(n_239)
);

INVx2_ASAP7_75t_L g308 ( 
.A(n_239),
.Y(n_308)
);

INVx4_ASAP7_75t_L g240 ( 
.A(n_164),
.Y(n_240)
);

INVx2_ASAP7_75t_L g316 ( 
.A(n_240),
.Y(n_316)
);

INVx2_ASAP7_75t_L g242 ( 
.A(n_171),
.Y(n_242)
);

INVxp67_ASAP7_75t_L g337 ( 
.A(n_242),
.Y(n_337)
);

AOI22xp33_ASAP7_75t_SL g244 ( 
.A1(n_215),
.A2(n_129),
.B1(n_127),
.B2(n_124),
.Y(n_244)
);

AOI22xp33_ASAP7_75t_SL g359 ( 
.A1(n_244),
.A2(n_248),
.B1(n_258),
.B2(n_297),
.Y(n_359)
);

OAI32xp33_ASAP7_75t_L g245 ( 
.A1(n_162),
.A2(n_99),
.A3(n_82),
.B1(n_79),
.B2(n_71),
.Y(n_245)
);

AND2x2_ASAP7_75t_L g313 ( 
.A(n_245),
.B(n_279),
.Y(n_313)
);

INVx2_ASAP7_75t_L g246 ( 
.A(n_158),
.Y(n_246)
);

INVxp67_ASAP7_75t_L g348 ( 
.A(n_246),
.Y(n_348)
);

INVx2_ASAP7_75t_L g247 ( 
.A(n_158),
.Y(n_247)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_247),
.Y(n_312)
);

AOI22xp33_ASAP7_75t_SL g248 ( 
.A1(n_217),
.A2(n_99),
.B1(n_126),
.B2(n_10),
.Y(n_248)
);

INVx5_ASAP7_75t_L g249 ( 
.A(n_141),
.Y(n_249)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_249),
.Y(n_314)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_225),
.Y(n_251)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_251),
.Y(n_325)
);

OAI22xp5_ASAP7_75t_SL g252 ( 
.A1(n_197),
.A2(n_0),
.B1(n_1),
.B2(n_3),
.Y(n_252)
);

AOI22xp5_ASAP7_75t_L g331 ( 
.A1(n_252),
.A2(n_264),
.B1(n_277),
.B2(n_284),
.Y(n_331)
);

NOR2xp33_ASAP7_75t_L g253 ( 
.A(n_183),
.B(n_7),
.Y(n_253)
);

NOR2xp33_ASAP7_75t_SL g360 ( 
.A(n_253),
.B(n_261),
.Y(n_360)
);

INVx2_ASAP7_75t_L g254 ( 
.A(n_201),
.Y(n_254)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_254),
.Y(n_326)
);

AOI22xp33_ASAP7_75t_L g255 ( 
.A1(n_167),
.A2(n_7),
.B1(n_16),
.B2(n_14),
.Y(n_255)
);

INVx2_ASAP7_75t_L g256 ( 
.A(n_207),
.Y(n_256)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_256),
.Y(n_330)
);

AOI22xp33_ASAP7_75t_L g257 ( 
.A1(n_165),
.A2(n_7),
.B1(n_16),
.B2(n_13),
.Y(n_257)
);

NAND2xp5_ASAP7_75t_L g261 ( 
.A(n_177),
.B(n_4),
.Y(n_261)
);

BUFx6f_ASAP7_75t_L g262 ( 
.A(n_185),
.Y(n_262)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_262),
.Y(n_332)
);

OAI21xp33_ASAP7_75t_L g362 ( 
.A1(n_263),
.A2(n_288),
.B(n_298),
.Y(n_362)
);

OAI22xp5_ASAP7_75t_SL g264 ( 
.A1(n_204),
.A2(n_0),
.B1(n_1),
.B2(n_3),
.Y(n_264)
);

INVx2_ASAP7_75t_L g265 ( 
.A(n_147),
.Y(n_265)
);

INVx1_ASAP7_75t_L g343 ( 
.A(n_265),
.Y(n_343)
);

CKINVDCx20_ASAP7_75t_R g266 ( 
.A(n_225),
.Y(n_266)
);

NAND2xp5_ASAP7_75t_SL g335 ( 
.A(n_266),
.B(n_278),
.Y(n_335)
);

BUFx6f_ASAP7_75t_L g267 ( 
.A(n_186),
.Y(n_267)
);

INVx1_ASAP7_75t_L g344 ( 
.A(n_267),
.Y(n_344)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_188),
.Y(n_268)
);

INVx1_ASAP7_75t_L g346 ( 
.A(n_268),
.Y(n_346)
);

INVx3_ASAP7_75t_L g269 ( 
.A(n_161),
.Y(n_269)
);

INVx1_ASAP7_75t_L g356 ( 
.A(n_269),
.Y(n_356)
);

NOR2xp33_ASAP7_75t_L g270 ( 
.A(n_183),
.B(n_4),
.Y(n_270)
);

NOR2xp33_ASAP7_75t_L g317 ( 
.A(n_270),
.B(n_281),
.Y(n_317)
);

INVx13_ASAP7_75t_L g271 ( 
.A(n_213),
.Y(n_271)
);

CKINVDCx14_ASAP7_75t_R g327 ( 
.A(n_271),
.Y(n_327)
);

AOI22xp33_ASAP7_75t_L g272 ( 
.A1(n_165),
.A2(n_4),
.B1(n_6),
.B2(n_8),
.Y(n_272)
);

INVx13_ASAP7_75t_L g273 ( 
.A(n_213),
.Y(n_273)
);

BUFx5_ASAP7_75t_L g309 ( 
.A(n_273),
.Y(n_309)
);

BUFx6f_ASAP7_75t_L g274 ( 
.A(n_186),
.Y(n_274)
);

INVx1_ASAP7_75t_L g361 ( 
.A(n_274),
.Y(n_361)
);

OAI22xp5_ASAP7_75t_L g336 ( 
.A1(n_275),
.A2(n_280),
.B1(n_159),
.B2(n_180),
.Y(n_336)
);

INVx2_ASAP7_75t_L g276 ( 
.A(n_155),
.Y(n_276)
);

INVx1_ASAP7_75t_L g366 ( 
.A(n_276),
.Y(n_366)
);

OAI22xp5_ASAP7_75t_SL g277 ( 
.A1(n_178),
.A2(n_3),
.B1(n_8),
.B2(n_18),
.Y(n_277)
);

NAND2xp5_ASAP7_75t_L g278 ( 
.A(n_191),
.B(n_18),
.Y(n_278)
);

INVx2_ASAP7_75t_L g279 ( 
.A(n_182),
.Y(n_279)
);

OAI22xp5_ASAP7_75t_L g280 ( 
.A1(n_133),
.A2(n_189),
.B1(n_181),
.B2(n_192),
.Y(n_280)
);

INVx3_ASAP7_75t_L g281 ( 
.A(n_156),
.Y(n_281)
);

INVx6_ASAP7_75t_L g282 ( 
.A(n_194),
.Y(n_282)
);

CKINVDCx20_ASAP7_75t_R g342 ( 
.A(n_282),
.Y(n_342)
);

INVx2_ASAP7_75t_L g283 ( 
.A(n_166),
.Y(n_283)
);

NOR2xp33_ASAP7_75t_L g318 ( 
.A(n_283),
.B(n_287),
.Y(n_318)
);

OAI22xp33_ASAP7_75t_L g284 ( 
.A1(n_220),
.A2(n_196),
.B1(n_224),
.B2(n_195),
.Y(n_284)
);

NAND2xp5_ASAP7_75t_L g285 ( 
.A(n_209),
.B(n_223),
.Y(n_285)
);

NAND2xp5_ASAP7_75t_SL g363 ( 
.A(n_285),
.B(n_286),
.Y(n_363)
);

CKINVDCx20_ASAP7_75t_R g286 ( 
.A(n_135),
.Y(n_286)
);

INVx2_ASAP7_75t_L g287 ( 
.A(n_173),
.Y(n_287)
);

NAND2xp5_ASAP7_75t_L g288 ( 
.A(n_138),
.B(n_154),
.Y(n_288)
);

INVx3_ASAP7_75t_L g289 ( 
.A(n_202),
.Y(n_289)
);

NOR2xp33_ASAP7_75t_L g324 ( 
.A(n_289),
.B(n_291),
.Y(n_324)
);

BUFx6f_ASAP7_75t_L g290 ( 
.A(n_194),
.Y(n_290)
);

CKINVDCx20_ASAP7_75t_R g352 ( 
.A(n_290),
.Y(n_352)
);

INVx6_ASAP7_75t_L g291 ( 
.A(n_210),
.Y(n_291)
);

OAI22xp5_ASAP7_75t_SL g292 ( 
.A1(n_149),
.A2(n_199),
.B1(n_196),
.B2(n_145),
.Y(n_292)
);

AO21x2_ASAP7_75t_L g338 ( 
.A1(n_292),
.A2(n_300),
.B(n_264),
.Y(n_338)
);

NOR2xp33_ASAP7_75t_L g293 ( 
.A(n_160),
.B(n_184),
.Y(n_293)
);

NOR2xp33_ASAP7_75t_L g345 ( 
.A(n_293),
.B(n_294),
.Y(n_345)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_163),
.Y(n_294)
);

INVxp33_ASAP7_75t_L g295 ( 
.A(n_198),
.Y(n_295)
);

NOR2xp33_ASAP7_75t_L g365 ( 
.A(n_295),
.B(n_296),
.Y(n_365)
);

INVx2_ASAP7_75t_L g296 ( 
.A(n_146),
.Y(n_296)
);

INVx2_ASAP7_75t_L g297 ( 
.A(n_203),
.Y(n_297)
);

NOR2xp33_ASAP7_75t_L g298 ( 
.A(n_143),
.B(n_148),
.Y(n_298)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_144),
.Y(n_299)
);

NAND2xp5_ASAP7_75t_L g311 ( 
.A(n_299),
.B(n_301),
.Y(n_311)
);

NAND2xp33_ASAP7_75t_SL g300 ( 
.A(n_217),
.B(n_216),
.Y(n_300)
);

AOI21xp5_ASAP7_75t_L g310 ( 
.A1(n_300),
.A2(n_248),
.B(n_244),
.Y(n_310)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_144),
.Y(n_301)
);

INVx2_ASAP7_75t_L g302 ( 
.A(n_206),
.Y(n_302)
);

NAND2xp5_ASAP7_75t_L g364 ( 
.A(n_302),
.B(n_303),
.Y(n_364)
);

INVx2_ASAP7_75t_L g303 ( 
.A(n_206),
.Y(n_303)
);

CKINVDCx20_ASAP7_75t_R g304 ( 
.A(n_152),
.Y(n_304)
);

NAND2xp5_ASAP7_75t_L g329 ( 
.A(n_304),
.B(n_305),
.Y(n_329)
);

INVx2_ASAP7_75t_L g305 ( 
.A(n_216),
.Y(n_305)
);

OR2x2_ASAP7_75t_L g395 ( 
.A(n_310),
.B(n_323),
.Y(n_395)
);

OAI22xp33_ASAP7_75t_SL g319 ( 
.A1(n_275),
.A2(n_214),
.B1(n_211),
.B2(n_222),
.Y(n_319)
);

AOI22xp33_ASAP7_75t_L g373 ( 
.A1(n_319),
.A2(n_239),
.B1(n_249),
.B2(n_273),
.Y(n_373)
);

OAI22xp5_ASAP7_75t_SL g321 ( 
.A1(n_259),
.A2(n_145),
.B1(n_195),
.B2(n_152),
.Y(n_321)
);

AOI22xp5_ASAP7_75t_L g367 ( 
.A1(n_321),
.A2(n_341),
.B1(n_351),
.B2(n_295),
.Y(n_367)
);

OA22x2_ASAP7_75t_L g323 ( 
.A1(n_245),
.A2(n_214),
.B1(n_211),
.B2(n_153),
.Y(n_323)
);

AND2x2_ASAP7_75t_L g375 ( 
.A(n_323),
.B(n_328),
.Y(n_375)
);

AND2x2_ASAP7_75t_SL g328 ( 
.A(n_243),
.B(n_148),
.Y(n_328)
);

AOI22xp33_ASAP7_75t_L g333 ( 
.A1(n_231),
.A2(n_210),
.B1(n_219),
.B2(n_153),
.Y(n_333)
);

OAI22xp33_ASAP7_75t_SL g393 ( 
.A1(n_333),
.A2(n_237),
.B1(n_338),
.B2(n_310),
.Y(n_393)
);

AND2x2_ASAP7_75t_L g376 ( 
.A(n_336),
.B(n_258),
.Y(n_376)
);

BUFx2_ASAP7_75t_L g398 ( 
.A(n_338),
.Y(n_398)
);

NAND2xp5_ASAP7_75t_L g339 ( 
.A(n_260),
.B(n_219),
.Y(n_339)
);

NAND2xp5_ASAP7_75t_L g386 ( 
.A(n_339),
.B(n_358),
.Y(n_386)
);

OAI22xp5_ASAP7_75t_SL g341 ( 
.A1(n_238),
.A2(n_218),
.B1(n_169),
.B2(n_180),
.Y(n_341)
);

XNOR2xp5_ASAP7_75t_L g347 ( 
.A(n_238),
.B(n_150),
.Y(n_347)
);

MAJIxp5_ASAP7_75t_L g371 ( 
.A(n_347),
.B(n_350),
.C(n_353),
.Y(n_371)
);

MAJIxp5_ASAP7_75t_L g350 ( 
.A(n_230),
.B(n_200),
.C(n_208),
.Y(n_350)
);

OAI22xp5_ASAP7_75t_SL g351 ( 
.A1(n_250),
.A2(n_241),
.B1(n_284),
.B2(n_252),
.Y(n_351)
);

MAJIxp5_ASAP7_75t_L g353 ( 
.A(n_229),
.B(n_218),
.C(n_221),
.Y(n_353)
);

XOR2xp5_ASAP7_75t_L g354 ( 
.A(n_236),
.B(n_221),
.Y(n_354)
);

MAJIxp5_ASAP7_75t_L g390 ( 
.A(n_354),
.B(n_302),
.C(n_303),
.Y(n_390)
);

AOI22xp5_ASAP7_75t_SL g357 ( 
.A1(n_277),
.A2(n_241),
.B1(n_250),
.B2(n_292),
.Y(n_357)
);

OAI21xp5_ASAP7_75t_SL g400 ( 
.A1(n_357),
.A2(n_359),
.B(n_323),
.Y(n_400)
);

NAND2xp5_ASAP7_75t_L g358 ( 
.A(n_241),
.B(n_256),
.Y(n_358)
);

OAI22xp5_ASAP7_75t_L g453 ( 
.A1(n_367),
.A2(n_369),
.B1(n_380),
.B2(n_384),
.Y(n_453)
);

XNOR2xp5_ASAP7_75t_L g368 ( 
.A(n_347),
.B(n_250),
.Y(n_368)
);

XOR2xp5_ASAP7_75t_L g423 ( 
.A(n_368),
.B(n_414),
.Y(n_423)
);

OAI22xp5_ASAP7_75t_L g369 ( 
.A1(n_357),
.A2(n_282),
.B1(n_291),
.B2(n_226),
.Y(n_369)
);

INVxp67_ASAP7_75t_L g370 ( 
.A(n_365),
.Y(n_370)
);

NOR2xp33_ASAP7_75t_L g426 ( 
.A(n_370),
.B(n_378),
.Y(n_426)
);

INVx1_ASAP7_75t_L g372 ( 
.A(n_329),
.Y(n_372)
);

INVx1_ASAP7_75t_L g416 ( 
.A(n_372),
.Y(n_416)
);

INVxp67_ASAP7_75t_L g436 ( 
.A(n_373),
.Y(n_436)
);

NOR2xp33_ASAP7_75t_L g374 ( 
.A(n_362),
.B(n_269),
.Y(n_374)
);

INVxp67_ASAP7_75t_L g439 ( 
.A(n_374),
.Y(n_439)
);

CKINVDCx14_ASAP7_75t_R g420 ( 
.A(n_376),
.Y(n_420)
);

OAI22xp5_ASAP7_75t_SL g377 ( 
.A1(n_358),
.A2(n_279),
.B1(n_254),
.B2(n_267),
.Y(n_377)
);

NAND2xp5_ASAP7_75t_L g415 ( 
.A(n_377),
.B(n_391),
.Y(n_415)
);

INVxp33_ASAP7_75t_L g378 ( 
.A(n_311),
.Y(n_378)
);

INVx1_ASAP7_75t_L g379 ( 
.A(n_329),
.Y(n_379)
);

INVx1_ASAP7_75t_L g427 ( 
.A(n_379),
.Y(n_427)
);

AOI22xp5_ASAP7_75t_L g380 ( 
.A1(n_313),
.A2(n_351),
.B1(n_331),
.B2(n_338),
.Y(n_380)
);

INVx1_ASAP7_75t_L g381 ( 
.A(n_340),
.Y(n_381)
);

INVx1_ASAP7_75t_L g428 ( 
.A(n_381),
.Y(n_428)
);

CKINVDCx20_ASAP7_75t_R g382 ( 
.A(n_327),
.Y(n_382)
);

NOR2xp33_ASAP7_75t_L g433 ( 
.A(n_382),
.B(n_409),
.Y(n_433)
);

INVx1_ASAP7_75t_L g383 ( 
.A(n_340),
.Y(n_383)
);

INVx1_ASAP7_75t_L g430 ( 
.A(n_383),
.Y(n_430)
);

AOI22xp5_ASAP7_75t_L g384 ( 
.A1(n_313),
.A2(n_281),
.B1(n_289),
.B2(n_290),
.Y(n_384)
);

AOI22xp5_ASAP7_75t_L g385 ( 
.A1(n_313),
.A2(n_227),
.B1(n_274),
.B2(n_262),
.Y(n_385)
);

OAI22xp5_ASAP7_75t_L g454 ( 
.A1(n_385),
.A2(n_387),
.B1(n_394),
.B2(n_411),
.Y(n_454)
);

AOI22xp5_ASAP7_75t_L g387 ( 
.A1(n_331),
.A2(n_234),
.B1(n_258),
.B2(n_305),
.Y(n_387)
);

INVx1_ASAP7_75t_L g388 ( 
.A(n_340),
.Y(n_388)
);

INVx1_ASAP7_75t_L g431 ( 
.A(n_388),
.Y(n_431)
);

INVx1_ASAP7_75t_L g389 ( 
.A(n_364),
.Y(n_389)
);

INVx1_ASAP7_75t_L g440 ( 
.A(n_389),
.Y(n_440)
);

XNOR2xp5_ASAP7_75t_SL g422 ( 
.A(n_390),
.B(n_330),
.Y(n_422)
);

OAI22xp5_ASAP7_75t_SL g391 ( 
.A1(n_338),
.A2(n_233),
.B1(n_228),
.B2(n_240),
.Y(n_391)
);

XOR2xp5_ASAP7_75t_L g392 ( 
.A(n_354),
.B(n_271),
.Y(n_392)
);

XNOR2xp5_ASAP7_75t_L g446 ( 
.A(n_392),
.B(n_407),
.Y(n_446)
);

INVx1_ASAP7_75t_L g443 ( 
.A(n_393),
.Y(n_443)
);

AOI22xp5_ASAP7_75t_L g394 ( 
.A1(n_338),
.A2(n_237),
.B1(n_315),
.B2(n_306),
.Y(n_394)
);

OAI21xp5_ASAP7_75t_SL g447 ( 
.A1(n_395),
.A2(n_400),
.B(n_404),
.Y(n_447)
);

NOR2xp33_ASAP7_75t_L g396 ( 
.A(n_345),
.B(n_339),
.Y(n_396)
);

INVxp67_ASAP7_75t_L g445 ( 
.A(n_396),
.Y(n_445)
);

NAND2xp5_ASAP7_75t_L g397 ( 
.A(n_363),
.B(n_335),
.Y(n_397)
);

NAND2xp5_ASAP7_75t_L g441 ( 
.A(n_397),
.B(n_399),
.Y(n_441)
);

NAND2xp5_ASAP7_75t_L g399 ( 
.A(n_353),
.B(n_317),
.Y(n_399)
);

NAND2xp5_ASAP7_75t_L g401 ( 
.A(n_328),
.B(n_360),
.Y(n_401)
);

NAND2xp5_ASAP7_75t_L g448 ( 
.A(n_401),
.B(n_326),
.Y(n_448)
);

NAND2xp5_ASAP7_75t_SL g402 ( 
.A(n_360),
.B(n_311),
.Y(n_402)
);

NAND2xp5_ASAP7_75t_SL g418 ( 
.A(n_402),
.B(n_408),
.Y(n_418)
);

AOI21xp5_ASAP7_75t_L g403 ( 
.A1(n_341),
.A2(n_350),
.B(n_364),
.Y(n_403)
);

OAI21xp5_ASAP7_75t_L g417 ( 
.A1(n_403),
.A2(n_314),
.B(n_316),
.Y(n_417)
);

AOI21xp5_ASAP7_75t_SL g404 ( 
.A1(n_328),
.A2(n_323),
.B(n_318),
.Y(n_404)
);

INVx2_ASAP7_75t_L g405 ( 
.A(n_309),
.Y(n_405)
);

INVx2_ASAP7_75t_L g452 ( 
.A(n_405),
.Y(n_452)
);

INVx1_ASAP7_75t_L g406 ( 
.A(n_325),
.Y(n_406)
);

INVx1_ASAP7_75t_SL g434 ( 
.A(n_406),
.Y(n_434)
);

MAJIxp5_ASAP7_75t_L g407 ( 
.A(n_346),
.B(n_312),
.C(n_343),
.Y(n_407)
);

NAND2xp5_ASAP7_75t_SL g408 ( 
.A(n_346),
.B(n_325),
.Y(n_408)
);

NAND2xp5_ASAP7_75t_SL g409 ( 
.A(n_312),
.B(n_356),
.Y(n_409)
);

AOI22xp33_ASAP7_75t_SL g410 ( 
.A1(n_352),
.A2(n_342),
.B1(n_356),
.B2(n_314),
.Y(n_410)
);

AOI22xp33_ASAP7_75t_SL g438 ( 
.A1(n_410),
.A2(n_308),
.B1(n_320),
.B2(n_355),
.Y(n_438)
);

OAI22xp5_ASAP7_75t_L g411 ( 
.A1(n_342),
.A2(n_321),
.B1(n_352),
.B2(n_324),
.Y(n_411)
);

INVx1_ASAP7_75t_L g412 ( 
.A(n_326),
.Y(n_412)
);

INVx1_ASAP7_75t_SL g450 ( 
.A(n_412),
.Y(n_450)
);

INVxp67_ASAP7_75t_L g413 ( 
.A(n_322),
.Y(n_413)
);

NOR2xp33_ASAP7_75t_L g444 ( 
.A(n_413),
.B(n_316),
.Y(n_444)
);

XNOR2xp5_ASAP7_75t_L g414 ( 
.A(n_343),
.B(n_366),
.Y(n_414)
);

XNOR2x1_ASAP7_75t_L g476 ( 
.A(n_417),
.B(n_422),
.Y(n_476)
);

OAI21xp5_ASAP7_75t_L g419 ( 
.A1(n_404),
.A2(n_348),
.B(n_366),
.Y(n_419)
);

OAI21xp5_ASAP7_75t_SL g477 ( 
.A1(n_419),
.A2(n_432),
.B(n_438),
.Y(n_477)
);

OA21x2_ASAP7_75t_SL g421 ( 
.A1(n_401),
.A2(n_399),
.B(n_386),
.Y(n_421)
);

OAI21xp5_ASAP7_75t_L g487 ( 
.A1(n_421),
.A2(n_451),
.B(n_307),
.Y(n_487)
);

CKINVDCx16_ASAP7_75t_R g424 ( 
.A(n_407),
.Y(n_424)
);

INVx1_ASAP7_75t_L g463 ( 
.A(n_424),
.Y(n_463)
);

OAI22xp5_ASAP7_75t_SL g425 ( 
.A1(n_380),
.A2(n_332),
.B1(n_344),
.B2(n_361),
.Y(n_425)
);

AOI22xp5_ASAP7_75t_L g458 ( 
.A1(n_425),
.A2(n_449),
.B1(n_383),
.B2(n_381),
.Y(n_458)
);

OA21x2_ASAP7_75t_L g429 ( 
.A1(n_395),
.A2(n_308),
.B(n_320),
.Y(n_429)
);

AND2x2_ASAP7_75t_L g468 ( 
.A(n_429),
.B(n_442),
.Y(n_468)
);

OAI21xp5_ASAP7_75t_L g432 ( 
.A1(n_395),
.A2(n_348),
.B(n_337),
.Y(n_432)
);

XOR2xp5_ASAP7_75t_L g435 ( 
.A(n_371),
.B(n_330),
.Y(n_435)
);

MAJIxp5_ASAP7_75t_L g464 ( 
.A(n_435),
.B(n_368),
.C(n_390),
.Y(n_464)
);

CKINVDCx20_ASAP7_75t_R g437 ( 
.A(n_413),
.Y(n_437)
);

CKINVDCx14_ASAP7_75t_R g466 ( 
.A(n_437),
.Y(n_466)
);

CKINVDCx20_ASAP7_75t_R g442 ( 
.A(n_370),
.Y(n_442)
);

NAND2xp5_ASAP7_75t_L g456 ( 
.A(n_444),
.B(n_448),
.Y(n_456)
);

OAI22xp5_ASAP7_75t_SL g449 ( 
.A1(n_386),
.A2(n_361),
.B1(n_332),
.B2(n_344),
.Y(n_449)
);

OAI21xp5_ASAP7_75t_SL g451 ( 
.A1(n_400),
.A2(n_337),
.B(n_355),
.Y(n_451)
);

INVx1_ASAP7_75t_SL g455 ( 
.A(n_419),
.Y(n_455)
);

NAND2xp5_ASAP7_75t_L g500 ( 
.A(n_455),
.B(n_459),
.Y(n_500)
);

OAI22xp5_ASAP7_75t_L g457 ( 
.A1(n_443),
.A2(n_397),
.B1(n_387),
.B2(n_394),
.Y(n_457)
);

OAI22xp5_ASAP7_75t_L g505 ( 
.A1(n_457),
.A2(n_465),
.B1(n_482),
.B2(n_484),
.Y(n_505)
);

INVx1_ASAP7_75t_L g494 ( 
.A(n_458),
.Y(n_494)
);

CKINVDCx20_ASAP7_75t_R g459 ( 
.A(n_433),
.Y(n_459)
);

XOR2xp5_ASAP7_75t_L g460 ( 
.A(n_435),
.B(n_371),
.Y(n_460)
);

MAJIxp5_ASAP7_75t_L g520 ( 
.A(n_460),
.B(n_464),
.C(n_483),
.Y(n_520)
);

OAI32xp33_ASAP7_75t_L g461 ( 
.A1(n_416),
.A2(n_375),
.A3(n_379),
.B1(n_372),
.B2(n_389),
.Y(n_461)
);

NAND2xp5_ASAP7_75t_L g503 ( 
.A(n_461),
.B(n_473),
.Y(n_503)
);

XNOR2xp5_ASAP7_75t_SL g462 ( 
.A(n_423),
.B(n_392),
.Y(n_462)
);

XNOR2xp5_ASAP7_75t_SL g522 ( 
.A(n_462),
.B(n_486),
.Y(n_522)
);

AOI22xp5_ASAP7_75t_L g465 ( 
.A1(n_443),
.A2(n_398),
.B1(n_375),
.B2(n_369),
.Y(n_465)
);

NAND2xp5_ASAP7_75t_L g467 ( 
.A(n_416),
.B(n_414),
.Y(n_467)
);

INVx1_ASAP7_75t_L g508 ( 
.A(n_467),
.Y(n_508)
);

INVx1_ASAP7_75t_L g469 ( 
.A(n_428),
.Y(n_469)
);

INVx1_ASAP7_75t_L g492 ( 
.A(n_469),
.Y(n_492)
);

OAI22xp5_ASAP7_75t_SL g470 ( 
.A1(n_420),
.A2(n_398),
.B1(n_367),
.B2(n_375),
.Y(n_470)
);

AOI22xp5_ASAP7_75t_L g495 ( 
.A1(n_470),
.A2(n_420),
.B1(n_429),
.B2(n_432),
.Y(n_495)
);

NAND2xp5_ASAP7_75t_SL g471 ( 
.A(n_418),
.B(n_382),
.Y(n_471)
);

NAND2xp5_ASAP7_75t_SL g498 ( 
.A(n_471),
.B(n_485),
.Y(n_498)
);

NAND2xp5_ASAP7_75t_L g472 ( 
.A(n_427),
.B(n_403),
.Y(n_472)
);

INVx1_ASAP7_75t_L g509 ( 
.A(n_472),
.Y(n_509)
);

CKINVDCx20_ASAP7_75t_R g473 ( 
.A(n_433),
.Y(n_473)
);

INVx1_ASAP7_75t_L g474 ( 
.A(n_428),
.Y(n_474)
);

INVx1_ASAP7_75t_L g493 ( 
.A(n_474),
.Y(n_493)
);

CKINVDCx20_ASAP7_75t_R g475 ( 
.A(n_444),
.Y(n_475)
);

NAND2xp5_ASAP7_75t_L g524 ( 
.A(n_475),
.B(n_479),
.Y(n_524)
);

NAND2xp5_ASAP7_75t_L g478 ( 
.A(n_427),
.B(n_411),
.Y(n_478)
);

INVx1_ASAP7_75t_L g510 ( 
.A(n_478),
.Y(n_510)
);

CKINVDCx20_ASAP7_75t_R g479 ( 
.A(n_426),
.Y(n_479)
);

BUFx2_ASAP7_75t_L g480 ( 
.A(n_452),
.Y(n_480)
);

INVx2_ASAP7_75t_L g502 ( 
.A(n_480),
.Y(n_502)
);

INVx1_ASAP7_75t_L g481 ( 
.A(n_430),
.Y(n_481)
);

INVx1_ASAP7_75t_L g501 ( 
.A(n_481),
.Y(n_501)
);

AOI22xp5_ASAP7_75t_L g482 ( 
.A1(n_454),
.A2(n_398),
.B1(n_391),
.B2(n_376),
.Y(n_482)
);

XOR2xp5_ASAP7_75t_L g483 ( 
.A(n_435),
.B(n_406),
.Y(n_483)
);

OAI22xp5_ASAP7_75t_L g484 ( 
.A1(n_453),
.A2(n_385),
.B1(n_376),
.B2(n_384),
.Y(n_484)
);

NAND2xp5_ASAP7_75t_SL g485 ( 
.A(n_418),
.B(n_412),
.Y(n_485)
);

A2O1A1O1Ixp25_ASAP7_75t_L g486 ( 
.A1(n_441),
.A2(n_388),
.B(n_377),
.C(n_405),
.D(n_309),
.Y(n_486)
);

CKINVDCx16_ASAP7_75t_R g504 ( 
.A(n_487),
.Y(n_504)
);

INVx1_ASAP7_75t_L g488 ( 
.A(n_430),
.Y(n_488)
);

INVx1_ASAP7_75t_L g516 ( 
.A(n_488),
.Y(n_516)
);

AOI21xp33_ASAP7_75t_L g489 ( 
.A1(n_439),
.A2(n_307),
.B(n_334),
.Y(n_489)
);

NOR2xp33_ASAP7_75t_L g496 ( 
.A(n_489),
.B(n_477),
.Y(n_496)
);

OAI22xp5_ASAP7_75t_L g490 ( 
.A1(n_453),
.A2(n_334),
.B1(n_349),
.B2(n_445),
.Y(n_490)
);

OAI22xp5_ASAP7_75t_L g518 ( 
.A1(n_490),
.A2(n_436),
.B1(n_437),
.B2(n_434),
.Y(n_518)
);

XNOR2xp5_ASAP7_75t_L g491 ( 
.A(n_421),
.B(n_349),
.Y(n_491)
);

XOR2xp5_ASAP7_75t_L g517 ( 
.A(n_491),
.B(n_446),
.Y(n_517)
);

OAI22xp5_ASAP7_75t_L g548 ( 
.A1(n_495),
.A2(n_514),
.B1(n_518),
.B2(n_448),
.Y(n_548)
);

INVxp67_ASAP7_75t_L g528 ( 
.A(n_496),
.Y(n_528)
);

XNOR2xp5_ASAP7_75t_L g497 ( 
.A(n_460),
.B(n_446),
.Y(n_497)
);

XOR2xp5_ASAP7_75t_L g536 ( 
.A(n_497),
.B(n_511),
.Y(n_536)
);

OAI22xp5_ASAP7_75t_SL g499 ( 
.A1(n_482),
.A2(n_441),
.B1(n_440),
.B2(n_415),
.Y(n_499)
);

AOI22xp5_ASAP7_75t_L g530 ( 
.A1(n_499),
.A2(n_513),
.B1(n_472),
.B2(n_417),
.Y(n_530)
);

CKINVDCx20_ASAP7_75t_R g506 ( 
.A(n_466),
.Y(n_506)
);

NAND2xp5_ASAP7_75t_L g529 ( 
.A(n_506),
.B(n_507),
.Y(n_529)
);

NOR2xp33_ASAP7_75t_L g507 ( 
.A(n_459),
.B(n_442),
.Y(n_507)
);

XNOR2xp5_ASAP7_75t_L g511 ( 
.A(n_464),
.B(n_446),
.Y(n_511)
);

BUFx3_ASAP7_75t_L g512 ( 
.A(n_480),
.Y(n_512)
);

INVx3_ASAP7_75t_L g541 ( 
.A(n_512),
.Y(n_541)
);

OAI22xp5_ASAP7_75t_SL g513 ( 
.A1(n_478),
.A2(n_440),
.B1(n_415),
.B2(n_447),
.Y(n_513)
);

AOI22xp5_ASAP7_75t_L g514 ( 
.A1(n_470),
.A2(n_454),
.B1(n_429),
.B2(n_425),
.Y(n_514)
);

INVx2_ASAP7_75t_L g515 ( 
.A(n_480),
.Y(n_515)
);

INVx1_ASAP7_75t_SL g556 ( 
.A(n_515),
.Y(n_556)
);

XOR2xp5_ASAP7_75t_L g551 ( 
.A(n_517),
.B(n_523),
.Y(n_551)
);

INVx1_ASAP7_75t_L g519 ( 
.A(n_469),
.Y(n_519)
);

INVx1_ASAP7_75t_L g532 ( 
.A(n_519),
.Y(n_532)
);

NOR2xp33_ASAP7_75t_L g521 ( 
.A(n_473),
.B(n_424),
.Y(n_521)
);

NAND2xp5_ASAP7_75t_L g542 ( 
.A(n_521),
.B(n_456),
.Y(n_542)
);

XNOR2xp5_ASAP7_75t_L g523 ( 
.A(n_483),
.B(n_422),
.Y(n_523)
);

XNOR2xp5_ASAP7_75t_SL g525 ( 
.A(n_462),
.B(n_423),
.Y(n_525)
);

XNOR2xp5_ASAP7_75t_SL g544 ( 
.A(n_525),
.B(n_476),
.Y(n_544)
);

INVx1_ASAP7_75t_L g526 ( 
.A(n_474),
.Y(n_526)
);

INVx1_ASAP7_75t_L g534 ( 
.A(n_526),
.Y(n_534)
);

OAI22xp5_ASAP7_75t_SL g527 ( 
.A1(n_514),
.A2(n_468),
.B1(n_455),
.B2(n_487),
.Y(n_527)
);

AOI22xp5_ASAP7_75t_L g565 ( 
.A1(n_527),
.A2(n_531),
.B1(n_538),
.B2(n_548),
.Y(n_565)
);

OAI22xp5_ASAP7_75t_L g566 ( 
.A1(n_530),
.A2(n_539),
.B1(n_522),
.B2(n_526),
.Y(n_566)
);

OAI22xp5_ASAP7_75t_SL g531 ( 
.A1(n_503),
.A2(n_468),
.B1(n_465),
.B2(n_479),
.Y(n_531)
);

MAJIxp5_ASAP7_75t_L g533 ( 
.A(n_520),
.B(n_463),
.C(n_422),
.Y(n_533)
);

MAJIxp5_ASAP7_75t_L g582 ( 
.A(n_533),
.B(n_540),
.C(n_434),
.Y(n_582)
);

AND2x2_ASAP7_75t_L g535 ( 
.A(n_494),
.B(n_468),
.Y(n_535)
);

INVx1_ASAP7_75t_L g571 ( 
.A(n_535),
.Y(n_571)
);

OR2x2_ASAP7_75t_L g537 ( 
.A(n_500),
.B(n_426),
.Y(n_537)
);

INVx1_ASAP7_75t_L g579 ( 
.A(n_537),
.Y(n_579)
);

OAI22xp5_ASAP7_75t_SL g538 ( 
.A1(n_503),
.A2(n_475),
.B1(n_456),
.B2(n_458),
.Y(n_538)
);

AOI22xp5_ASAP7_75t_L g539 ( 
.A1(n_505),
.A2(n_429),
.B1(n_491),
.B2(n_463),
.Y(n_539)
);

MAJIxp5_ASAP7_75t_L g540 ( 
.A(n_520),
.B(n_476),
.C(n_423),
.Y(n_540)
);

NAND2xp5_ASAP7_75t_SL g563 ( 
.A(n_542),
.B(n_546),
.Y(n_563)
);

NAND2xp5_ASAP7_75t_L g543 ( 
.A(n_498),
.B(n_461),
.Y(n_543)
);

NOR2xp33_ASAP7_75t_SL g576 ( 
.A(n_543),
.B(n_545),
.Y(n_576)
);

XNOR2xp5_ASAP7_75t_SL g568 ( 
.A(n_544),
.B(n_523),
.Y(n_568)
);

NOR2xp33_ASAP7_75t_L g545 ( 
.A(n_508),
.B(n_524),
.Y(n_545)
);

NAND2xp5_ASAP7_75t_L g546 ( 
.A(n_524),
.B(n_452),
.Y(n_546)
);

XNOR2xp5_ASAP7_75t_L g547 ( 
.A(n_511),
.B(n_447),
.Y(n_547)
);

XNOR2xp5_ASAP7_75t_L g560 ( 
.A(n_547),
.B(n_552),
.Y(n_560)
);

NOR2x1_ASAP7_75t_R g549 ( 
.A(n_513),
.B(n_477),
.Y(n_549)
);

INVx1_ASAP7_75t_L g572 ( 
.A(n_549),
.Y(n_572)
);

NOR2xp33_ASAP7_75t_L g550 ( 
.A(n_508),
.B(n_431),
.Y(n_550)
);

NAND2xp5_ASAP7_75t_SL g575 ( 
.A(n_550),
.B(n_554),
.Y(n_575)
);

XNOR2xp5_ASAP7_75t_L g552 ( 
.A(n_497),
.B(n_467),
.Y(n_552)
);

XOR2xp5_ASAP7_75t_L g553 ( 
.A(n_525),
.B(n_451),
.Y(n_553)
);

XOR2xp5_ASAP7_75t_L g561 ( 
.A(n_553),
.B(n_555),
.Y(n_561)
);

NAND2xp5_ASAP7_75t_SL g554 ( 
.A(n_500),
.B(n_431),
.Y(n_554)
);

XOR2xp5_ASAP7_75t_L g555 ( 
.A(n_517),
.B(n_481),
.Y(n_555)
);

CKINVDCx20_ASAP7_75t_R g557 ( 
.A(n_499),
.Y(n_557)
);

NAND2xp5_ASAP7_75t_SL g581 ( 
.A(n_557),
.B(n_547),
.Y(n_581)
);

OAI22xp5_ASAP7_75t_SL g558 ( 
.A1(n_539),
.A2(n_510),
.B1(n_494),
.B2(n_495),
.Y(n_558)
);

AOI22xp5_ASAP7_75t_L g584 ( 
.A1(n_558),
.A2(n_559),
.B1(n_566),
.B2(n_527),
.Y(n_584)
);

OAI22xp5_ASAP7_75t_SL g559 ( 
.A1(n_530),
.A2(n_510),
.B1(n_504),
.B2(n_509),
.Y(n_559)
);

NOR2xp33_ASAP7_75t_L g562 ( 
.A(n_528),
.B(n_509),
.Y(n_562)
);

NAND2xp5_ASAP7_75t_L g590 ( 
.A(n_562),
.B(n_578),
.Y(n_590)
);

NAND2xp5_ASAP7_75t_L g564 ( 
.A(n_538),
.B(n_488),
.Y(n_564)
);

INVx1_ASAP7_75t_L g596 ( 
.A(n_564),
.Y(n_596)
);

XNOR2xp5_ASAP7_75t_L g567 ( 
.A(n_533),
.B(n_536),
.Y(n_567)
);

XNOR2xp5_ASAP7_75t_L g585 ( 
.A(n_567),
.B(n_569),
.Y(n_585)
);

XOR2xp5_ASAP7_75t_L g593 ( 
.A(n_568),
.B(n_544),
.Y(n_593)
);

XNOR2xp5_ASAP7_75t_L g569 ( 
.A(n_536),
.B(n_522),
.Y(n_569)
);

NAND2xp5_ASAP7_75t_L g570 ( 
.A(n_529),
.B(n_519),
.Y(n_570)
);

CKINVDCx20_ASAP7_75t_R g597 ( 
.A(n_570),
.Y(n_597)
);

AOI22xp5_ASAP7_75t_L g573 ( 
.A1(n_531),
.A2(n_493),
.B1(n_501),
.B2(n_516),
.Y(n_573)
);

OAI22xp5_ASAP7_75t_SL g589 ( 
.A1(n_573),
.A2(n_534),
.B1(n_532),
.B2(n_556),
.Y(n_589)
);

OAI21xp5_ASAP7_75t_L g574 ( 
.A1(n_535),
.A2(n_486),
.B(n_492),
.Y(n_574)
);

INVxp33_ASAP7_75t_L g583 ( 
.A(n_574),
.Y(n_583)
);

OAI21xp5_ASAP7_75t_L g577 ( 
.A1(n_535),
.A2(n_438),
.B(n_449),
.Y(n_577)
);

AOI21xp5_ASAP7_75t_L g600 ( 
.A1(n_577),
.A2(n_502),
.B(n_515),
.Y(n_600)
);

HB1xp67_ASAP7_75t_L g578 ( 
.A(n_541),
.Y(n_578)
);

CKINVDCx20_ASAP7_75t_R g580 ( 
.A(n_537),
.Y(n_580)
);

NAND2xp5_ASAP7_75t_L g601 ( 
.A(n_580),
.B(n_450),
.Y(n_601)
);

OAI21x1_ASAP7_75t_L g586 ( 
.A1(n_581),
.A2(n_555),
.B(n_551),
.Y(n_586)
);

XNOR2xp5_ASAP7_75t_L g588 ( 
.A(n_582),
.B(n_551),
.Y(n_588)
);

XNOR2x1_ASAP7_75t_L g612 ( 
.A(n_584),
.B(n_593),
.Y(n_612)
);

AOI31xp33_ASAP7_75t_L g607 ( 
.A1(n_586),
.A2(n_579),
.A3(n_572),
.B(n_577),
.Y(n_607)
);

BUFx4f_ASAP7_75t_SL g587 ( 
.A(n_571),
.Y(n_587)
);

INVx1_ASAP7_75t_L g610 ( 
.A(n_587),
.Y(n_610)
);

XNOR2xp5_ASAP7_75t_L g611 ( 
.A(n_588),
.B(n_592),
.Y(n_611)
);

INVx1_ASAP7_75t_L g613 ( 
.A(n_589),
.Y(n_613)
);

MAJIxp5_ASAP7_75t_L g591 ( 
.A(n_582),
.B(n_540),
.C(n_552),
.Y(n_591)
);

NAND2xp5_ASAP7_75t_L g614 ( 
.A(n_591),
.B(n_594),
.Y(n_614)
);

XNOR2xp5_ASAP7_75t_L g592 ( 
.A(n_560),
.B(n_553),
.Y(n_592)
);

MAJIxp5_ASAP7_75t_L g594 ( 
.A(n_567),
.B(n_549),
.C(n_528),
.Y(n_594)
);

OAI22xp5_ASAP7_75t_SL g595 ( 
.A1(n_565),
.A2(n_556),
.B1(n_541),
.B2(n_502),
.Y(n_595)
);

NAND2xp5_ASAP7_75t_SL g604 ( 
.A(n_595),
.B(n_599),
.Y(n_604)
);

NOR2xp33_ASAP7_75t_L g598 ( 
.A(n_576),
.B(n_512),
.Y(n_598)
);

INVx1_ASAP7_75t_L g617 ( 
.A(n_598),
.Y(n_617)
);

MAJIxp5_ASAP7_75t_L g599 ( 
.A(n_560),
.B(n_450),
.C(n_434),
.Y(n_599)
);

MAJx2_ASAP7_75t_L g615 ( 
.A(n_600),
.B(n_559),
.C(n_564),
.Y(n_615)
);

INVx1_ASAP7_75t_L g619 ( 
.A(n_601),
.Y(n_619)
);

NAND2xp5_ASAP7_75t_SL g602 ( 
.A(n_575),
.B(n_450),
.Y(n_602)
);

OAI21xp5_ASAP7_75t_SL g606 ( 
.A1(n_602),
.A2(n_570),
.B(n_563),
.Y(n_606)
);

AOI21xp5_ASAP7_75t_L g603 ( 
.A1(n_583),
.A2(n_574),
.B(n_572),
.Y(n_603)
);

OR2x2_ASAP7_75t_L g621 ( 
.A(n_603),
.B(n_615),
.Y(n_621)
);

MAJIxp5_ASAP7_75t_L g605 ( 
.A(n_588),
.B(n_571),
.C(n_561),
.Y(n_605)
);

NAND2xp5_ASAP7_75t_L g632 ( 
.A(n_605),
.B(n_608),
.Y(n_632)
);

NAND2xp5_ASAP7_75t_SL g623 ( 
.A(n_606),
.B(n_618),
.Y(n_623)
);

OAI21xp5_ASAP7_75t_L g631 ( 
.A1(n_607),
.A2(n_587),
.B(n_593),
.Y(n_631)
);

AND2x2_ASAP7_75t_L g608 ( 
.A(n_600),
.B(n_565),
.Y(n_608)
);

MAJIxp5_ASAP7_75t_L g609 ( 
.A(n_591),
.B(n_561),
.C(n_569),
.Y(n_609)
);

NAND2xp5_ASAP7_75t_L g633 ( 
.A(n_609),
.B(n_616),
.Y(n_633)
);

MAJIxp5_ASAP7_75t_L g616 ( 
.A(n_585),
.B(n_558),
.C(n_573),
.Y(n_616)
);

XNOR2xp5_ASAP7_75t_L g618 ( 
.A(n_594),
.B(n_568),
.Y(n_618)
);

NOR2xp67_ASAP7_75t_SL g620 ( 
.A(n_614),
.B(n_585),
.Y(n_620)
);

AOI21xp5_ASAP7_75t_L g638 ( 
.A1(n_620),
.A2(n_618),
.B(n_612),
.Y(n_638)
);

XNOR2xp5_ASAP7_75t_L g622 ( 
.A(n_611),
.B(n_590),
.Y(n_622)
);

NAND2xp5_ASAP7_75t_SL g640 ( 
.A(n_622),
.B(n_624),
.Y(n_640)
);

MAJIxp5_ASAP7_75t_L g624 ( 
.A(n_611),
.B(n_584),
.C(n_599),
.Y(n_624)
);

XNOR2xp5_ASAP7_75t_L g625 ( 
.A(n_605),
.B(n_592),
.Y(n_625)
);

NOR2xp33_ASAP7_75t_SL g642 ( 
.A(n_625),
.B(n_626),
.Y(n_642)
);

NAND2xp5_ASAP7_75t_SL g626 ( 
.A(n_617),
.B(n_597),
.Y(n_626)
);

NOR2xp33_ASAP7_75t_SL g627 ( 
.A(n_609),
.B(n_583),
.Y(n_627)
);

NOR2xp33_ASAP7_75t_L g641 ( 
.A(n_627),
.B(n_612),
.Y(n_641)
);

BUFx6f_ASAP7_75t_L g628 ( 
.A(n_610),
.Y(n_628)
);

INVx1_ASAP7_75t_L g635 ( 
.A(n_628),
.Y(n_635)
);

XOR2xp5_ASAP7_75t_L g629 ( 
.A(n_616),
.B(n_595),
.Y(n_629)
);

AND2x2_ASAP7_75t_L g639 ( 
.A(n_629),
.B(n_630),
.Y(n_639)
);

MAJIxp5_ASAP7_75t_L g630 ( 
.A(n_604),
.B(n_596),
.C(n_589),
.Y(n_630)
);

MAJIxp5_ASAP7_75t_L g634 ( 
.A(n_630),
.B(n_608),
.C(n_615),
.Y(n_634)
);

AOI22xp5_ASAP7_75t_L g643 ( 
.A1(n_631),
.A2(n_587),
.B1(n_621),
.B2(n_628),
.Y(n_643)
);

INVxp33_ASAP7_75t_L g646 ( 
.A(n_634),
.Y(n_646)
);

MAJIxp5_ASAP7_75t_L g636 ( 
.A(n_629),
.B(n_608),
.C(n_613),
.Y(n_636)
);

NAND2xp5_ASAP7_75t_SL g649 ( 
.A(n_636),
.B(n_639),
.Y(n_649)
);

OAI21xp5_ASAP7_75t_SL g637 ( 
.A1(n_623),
.A2(n_603),
.B(n_619),
.Y(n_637)
);

OAI21xp5_ASAP7_75t_L g644 ( 
.A1(n_637),
.A2(n_638),
.B(n_643),
.Y(n_644)
);

NOR2xp33_ASAP7_75t_SL g648 ( 
.A(n_641),
.B(n_621),
.Y(n_648)
);

MAJIxp5_ASAP7_75t_L g645 ( 
.A(n_640),
.B(n_633),
.C(n_632),
.Y(n_645)
);

OR2x2_ASAP7_75t_L g654 ( 
.A(n_645),
.B(n_647),
.Y(n_654)
);

XOR2xp5_ASAP7_75t_L g647 ( 
.A(n_634),
.B(n_624),
.Y(n_647)
);

INVxp33_ASAP7_75t_SL g651 ( 
.A(n_648),
.Y(n_651)
);

XOR2xp5_ASAP7_75t_L g650 ( 
.A(n_639),
.B(n_636),
.Y(n_650)
);

NOR2xp67_ASAP7_75t_SL g652 ( 
.A(n_650),
.B(n_642),
.Y(n_652)
);

MAJIxp5_ASAP7_75t_L g656 ( 
.A(n_652),
.B(n_651),
.C(n_646),
.Y(n_656)
);

NOR2xp33_ASAP7_75t_SL g653 ( 
.A(n_644),
.B(n_635),
.Y(n_653)
);

NOR3xp33_ASAP7_75t_L g655 ( 
.A(n_653),
.B(n_649),
.C(n_650),
.Y(n_655)
);

INVxp67_ASAP7_75t_L g657 ( 
.A(n_655),
.Y(n_657)
);

NOR3xp33_ASAP7_75t_L g658 ( 
.A(n_657),
.B(n_656),
.C(n_654),
.Y(n_658)
);

XOR2xp5_ASAP7_75t_L g659 ( 
.A(n_658),
.B(n_646),
.Y(n_659)
);

BUFx24_ASAP7_75t_SL g660 ( 
.A(n_659),
.Y(n_660)
);


endmodule