module fake_netlist_5_2450_n_138 (n_54, n_29, n_16, n_43, n_0, n_12, n_9, n_47, n_58, n_36, n_25, n_53, n_18, n_27, n_42, n_22, n_1, n_8, n_45, n_10, n_24, n_28, n_46, n_21, n_44, n_40, n_34, n_38, n_4, n_32, n_35, n_41, n_56, n_51, n_11, n_17, n_19, n_57, n_7, n_37, n_59, n_15, n_26, n_30, n_20, n_5, n_33, n_55, n_14, n_48, n_2, n_31, n_23, n_13, n_50, n_3, n_49, n_52, n_6, n_39, n_138);

input n_54;
input n_29;
input n_16;
input n_43;
input n_0;
input n_12;
input n_9;
input n_47;
input n_58;
input n_36;
input n_25;
input n_53;
input n_18;
input n_27;
input n_42;
input n_22;
input n_1;
input n_8;
input n_45;
input n_10;
input n_24;
input n_28;
input n_46;
input n_21;
input n_44;
input n_40;
input n_34;
input n_38;
input n_4;
input n_32;
input n_35;
input n_41;
input n_56;
input n_51;
input n_11;
input n_17;
input n_19;
input n_57;
input n_7;
input n_37;
input n_59;
input n_15;
input n_26;
input n_30;
input n_20;
input n_5;
input n_33;
input n_55;
input n_14;
input n_48;
input n_2;
input n_31;
input n_23;
input n_13;
input n_50;
input n_3;
input n_49;
input n_52;
input n_6;
input n_39;

output n_138;

wire n_137;
wire n_91;
wire n_82;
wire n_122;
wire n_124;
wire n_86;
wire n_136;
wire n_83;
wire n_132;
wire n_61;
wire n_90;
wire n_127;
wire n_75;
wire n_101;
wire n_78;
wire n_65;
wire n_74;
wire n_114;
wire n_96;
wire n_111;
wire n_108;
wire n_129;
wire n_66;
wire n_98;
wire n_60;
wire n_107;
wire n_69;
wire n_116;
wire n_117;
wire n_94;
wire n_113;
wire n_123;
wire n_105;
wire n_80;
wire n_125;
wire n_128;
wire n_73;
wire n_92;
wire n_120;
wire n_135;
wire n_126;
wire n_84;
wire n_130;
wire n_79;
wire n_131;
wire n_100;
wire n_62;
wire n_71;
wire n_109;
wire n_112;
wire n_85;
wire n_95;
wire n_119;
wire n_133;
wire n_99;
wire n_67;
wire n_121;
wire n_76;
wire n_87;
wire n_64;
wire n_77;
wire n_106;
wire n_102;
wire n_81;
wire n_118;
wire n_89;
wire n_70;
wire n_115;
wire n_68;
wire n_93;
wire n_72;
wire n_134;
wire n_104;
wire n_103;
wire n_63;
wire n_97;
wire n_88;
wire n_110;

INVx1_ASAP7_75t_L g60 ( 
.A(n_23),
.Y(n_60)
);

OAI22xp5_ASAP7_75t_SL g61 ( 
.A1(n_19),
.A2(n_57),
.B1(n_36),
.B2(n_12),
.Y(n_61)
);

AND2x2_ASAP7_75t_L g62 ( 
.A(n_52),
.B(n_44),
.Y(n_62)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_27),
.Y(n_63)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_2),
.Y(n_64)
);

OAI22xp5_ASAP7_75t_L g65 ( 
.A1(n_28),
.A2(n_13),
.B1(n_31),
.B2(n_11),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_L g66 ( 
.A(n_17),
.B(n_9),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_L g67 ( 
.A(n_8),
.B(n_46),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_L g68 ( 
.A(n_59),
.B(n_5),
.Y(n_68)
);

INVx3_ASAP7_75t_L g69 ( 
.A(n_45),
.Y(n_69)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_30),
.Y(n_70)
);

INVx6_ASAP7_75t_L g71 ( 
.A(n_53),
.Y(n_71)
);

INVx2_ASAP7_75t_L g72 ( 
.A(n_21),
.Y(n_72)
);

AND2x2_ASAP7_75t_L g73 ( 
.A(n_25),
.B(n_40),
.Y(n_73)
);

INVx4_ASAP7_75t_L g74 ( 
.A(n_33),
.Y(n_74)
);

INVx4_ASAP7_75t_L g75 ( 
.A(n_54),
.Y(n_75)
);

BUFx3_ASAP7_75t_L g76 ( 
.A(n_39),
.Y(n_76)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_20),
.Y(n_77)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_3),
.Y(n_78)
);

CKINVDCx20_ASAP7_75t_R g79 ( 
.A(n_15),
.Y(n_79)
);

OAI22xp5_ASAP7_75t_L g80 ( 
.A1(n_51),
.A2(n_29),
.B1(n_48),
.B2(n_49),
.Y(n_80)
);

INVx2_ASAP7_75t_L g81 ( 
.A(n_58),
.Y(n_81)
);

AND2x4_ASAP7_75t_L g82 ( 
.A(n_50),
.B(n_7),
.Y(n_82)
);

BUFx6f_ASAP7_75t_L g83 ( 
.A(n_47),
.Y(n_83)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_42),
.Y(n_84)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_55),
.Y(n_85)
);

AND2x4_ASAP7_75t_L g86 ( 
.A(n_22),
.B(n_56),
.Y(n_86)
);

CKINVDCx5p33_ASAP7_75t_R g87 ( 
.A(n_6),
.Y(n_87)
);

HB1xp67_ASAP7_75t_L g88 ( 
.A(n_24),
.Y(n_88)
);

INVx3_ASAP7_75t_L g89 ( 
.A(n_43),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_SL g90 ( 
.A(n_88),
.B(n_89),
.Y(n_90)
);

AOI22xp33_ASAP7_75t_L g91 ( 
.A1(n_69),
.A2(n_0),
.B1(n_1),
.B2(n_4),
.Y(n_91)
);

INVx2_ASAP7_75t_SL g92 ( 
.A(n_71),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_60),
.B(n_10),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_L g94 ( 
.A(n_70),
.B(n_14),
.Y(n_94)
);

NAND3xp33_ASAP7_75t_L g95 ( 
.A(n_74),
.B(n_16),
.C(n_18),
.Y(n_95)
);

BUFx3_ASAP7_75t_L g96 ( 
.A(n_76),
.Y(n_96)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_63),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g98 ( 
.A(n_72),
.B(n_26),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_SL g99 ( 
.A(n_83),
.B(n_32),
.Y(n_99)
);

INVx2_ASAP7_75t_L g100 ( 
.A(n_64),
.Y(n_100)
);

BUFx6f_ASAP7_75t_L g101 ( 
.A(n_83),
.Y(n_101)
);

INVx2_ASAP7_75t_L g102 ( 
.A(n_77),
.Y(n_102)
);

BUFx8_ASAP7_75t_L g103 ( 
.A(n_62),
.Y(n_103)
);

AND2x4_ASAP7_75t_L g104 ( 
.A(n_78),
.B(n_34),
.Y(n_104)
);

OAI22xp33_ASAP7_75t_L g105 ( 
.A1(n_84),
.A2(n_35),
.B1(n_37),
.B2(n_38),
.Y(n_105)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_85),
.Y(n_106)
);

INVx4_ASAP7_75t_L g107 ( 
.A(n_96),
.Y(n_107)
);

OR2x6_ASAP7_75t_L g108 ( 
.A(n_92),
.B(n_61),
.Y(n_108)
);

OAI21x1_ASAP7_75t_L g109 ( 
.A1(n_94),
.A2(n_68),
.B(n_66),
.Y(n_109)
);

OAI21xp5_ASAP7_75t_L g110 ( 
.A1(n_90),
.A2(n_73),
.B(n_86),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_L g111 ( 
.A(n_104),
.B(n_81),
.Y(n_111)
);

OAI21xp5_ASAP7_75t_L g112 ( 
.A1(n_97),
.A2(n_106),
.B(n_93),
.Y(n_112)
);

OA22x2_ASAP7_75t_L g113 ( 
.A1(n_100),
.A2(n_87),
.B1(n_82),
.B2(n_75),
.Y(n_113)
);

AOI221xp5_ASAP7_75t_SL g114 ( 
.A1(n_102),
.A2(n_98),
.B1(n_105),
.B2(n_91),
.C(n_99),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g115 ( 
.A(n_101),
.B(n_67),
.Y(n_115)
);

AOI21xp33_ASAP7_75t_L g116 ( 
.A1(n_103),
.A2(n_80),
.B(n_65),
.Y(n_116)
);

AO21x2_ASAP7_75t_L g117 ( 
.A1(n_95),
.A2(n_79),
.B(n_41),
.Y(n_117)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_115),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_L g119 ( 
.A(n_111),
.B(n_110),
.Y(n_119)
);

INVx2_ASAP7_75t_L g120 ( 
.A(n_107),
.Y(n_120)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_113),
.Y(n_121)
);

BUFx2_ASAP7_75t_L g122 ( 
.A(n_108),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_L g123 ( 
.A(n_119),
.B(n_114),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_L g124 ( 
.A(n_118),
.B(n_112),
.Y(n_124)
);

INVx2_ASAP7_75t_L g125 ( 
.A(n_121),
.Y(n_125)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_120),
.Y(n_126)
);

INVx2_ASAP7_75t_L g127 ( 
.A(n_122),
.Y(n_127)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_125),
.Y(n_128)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_126),
.Y(n_129)
);

AOI22xp5_ASAP7_75t_L g130 ( 
.A1(n_123),
.A2(n_109),
.B1(n_117),
.B2(n_116),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_SL g131 ( 
.A(n_129),
.B(n_127),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_L g132 ( 
.A(n_131),
.B(n_124),
.Y(n_132)
);

INVx1_ASAP7_75t_SL g133 ( 
.A(n_132),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_L g134 ( 
.A(n_133),
.B(n_128),
.Y(n_134)
);

HB1xp67_ASAP7_75t_L g135 ( 
.A(n_133),
.Y(n_135)
);

HB1xp67_ASAP7_75t_L g136 ( 
.A(n_135),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_L g137 ( 
.A(n_136),
.B(n_134),
.Y(n_137)
);

AOI21xp5_ASAP7_75t_L g138 ( 
.A1(n_137),
.A2(n_130),
.B(n_108),
.Y(n_138)
);


endmodule