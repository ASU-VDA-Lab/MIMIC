module fake_jpeg_25049_n_226 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_226);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_226;

wire n_159;
wire n_117;
wire n_144;
wire n_225;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_57;
wire n_21;
wire n_223;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_24;
wire n_44;
wire n_143;
wire n_202;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_131;
wire n_56;
wire n_212;
wire n_211;
wire n_183;
wire n_79;
wire n_170;
wire n_162;
wire n_132;
wire n_133;
wire n_67;
wire n_216;
wire n_217;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

INVx1_ASAP7_75t_L g16 ( 
.A(n_15),
.Y(n_16)
);

BUFx12_ASAP7_75t_L g17 ( 
.A(n_5),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_14),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_5),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_2),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_11),
.Y(n_21)
);

BUFx12_ASAP7_75t_L g22 ( 
.A(n_13),
.Y(n_22)
);

BUFx12_ASAP7_75t_L g23 ( 
.A(n_9),
.Y(n_23)
);

INVx2_ASAP7_75t_L g24 ( 
.A(n_9),
.Y(n_24)
);

BUFx12f_ASAP7_75t_L g25 ( 
.A(n_4),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_15),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_6),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_6),
.Y(n_28)
);

INVx4_ASAP7_75t_L g29 ( 
.A(n_13),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_1),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_5),
.Y(n_31)
);

BUFx8_ASAP7_75t_L g32 ( 
.A(n_12),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_2),
.Y(n_33)
);

INVx2_ASAP7_75t_L g34 ( 
.A(n_24),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_34),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_25),
.Y(n_35)
);

INVx4_ASAP7_75t_L g54 ( 
.A(n_35),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_25),
.Y(n_36)
);

INVx4_ASAP7_75t_L g62 ( 
.A(n_36),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g37 ( 
.A(n_25),
.B(n_0),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_37),
.B(n_39),
.Y(n_66)
);

BUFx16f_ASAP7_75t_L g38 ( 
.A(n_17),
.Y(n_38)
);

INVx5_ASAP7_75t_L g49 ( 
.A(n_38),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_L g39 ( 
.A(n_24),
.B(n_0),
.Y(n_39)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_30),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_40),
.B(n_45),
.Y(n_55)
);

INVx2_ASAP7_75t_L g41 ( 
.A(n_25),
.Y(n_41)
);

BUFx2_ASAP7_75t_SL g59 ( 
.A(n_41),
.Y(n_59)
);

INVx4_ASAP7_75t_L g42 ( 
.A(n_25),
.Y(n_42)
);

HB1xp67_ASAP7_75t_L g67 ( 
.A(n_42),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_SL g43 ( 
.A(n_30),
.B(n_31),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_SL g48 ( 
.A(n_43),
.B(n_26),
.Y(n_48)
);

INVx2_ASAP7_75t_L g44 ( 
.A(n_20),
.Y(n_44)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_44),
.Y(n_52)
);

INVx3_ASAP7_75t_L g45 ( 
.A(n_20),
.Y(n_45)
);

MAJIxp5_ASAP7_75t_L g47 ( 
.A(n_39),
.B(n_29),
.C(n_20),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_47),
.B(n_48),
.Y(n_71)
);

INVxp67_ASAP7_75t_L g50 ( 
.A(n_37),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_50),
.B(n_51),
.Y(n_77)
);

INVx3_ASAP7_75t_L g51 ( 
.A(n_35),
.Y(n_51)
);

MAJIxp5_ASAP7_75t_L g53 ( 
.A(n_41),
.B(n_29),
.C(n_27),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_L g70 ( 
.A(n_53),
.B(n_63),
.Y(n_70)
);

INVx11_ASAP7_75t_L g56 ( 
.A(n_35),
.Y(n_56)
);

INVx8_ASAP7_75t_L g82 ( 
.A(n_56),
.Y(n_82)
);

AOI22xp33_ASAP7_75t_L g57 ( 
.A1(n_45),
.A2(n_29),
.B1(n_31),
.B2(n_19),
.Y(n_57)
);

OAI22xp5_ASAP7_75t_L g88 ( 
.A1(n_57),
.A2(n_32),
.B1(n_23),
.B2(n_17),
.Y(n_88)
);

INVx3_ASAP7_75t_L g58 ( 
.A(n_36),
.Y(n_58)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_58),
.Y(n_89)
);

AOI22xp33_ASAP7_75t_SL g60 ( 
.A1(n_44),
.A2(n_18),
.B1(n_26),
.B2(n_19),
.Y(n_60)
);

CKINVDCx14_ASAP7_75t_R g80 ( 
.A(n_60),
.Y(n_80)
);

OR2x2_ASAP7_75t_L g61 ( 
.A(n_34),
.B(n_18),
.Y(n_61)
);

CKINVDCx16_ASAP7_75t_R g73 ( 
.A(n_61),
.Y(n_73)
);

MAJIxp5_ASAP7_75t_L g63 ( 
.A(n_42),
.B(n_28),
.C(n_27),
.Y(n_63)
);

NOR2x1_ASAP7_75t_L g64 ( 
.A(n_43),
.B(n_32),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_L g75 ( 
.A(n_64),
.B(n_68),
.Y(n_75)
);

AOI22xp33_ASAP7_75t_SL g65 ( 
.A1(n_40),
.A2(n_33),
.B1(n_16),
.B2(n_32),
.Y(n_65)
);

OAI22xp5_ASAP7_75t_SL g81 ( 
.A1(n_65),
.A2(n_16),
.B1(n_32),
.B2(n_17),
.Y(n_81)
);

OR2x2_ASAP7_75t_L g68 ( 
.A(n_36),
.B(n_28),
.Y(n_68)
);

INVxp33_ASAP7_75t_L g69 ( 
.A(n_59),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_69),
.B(n_76),
.Y(n_90)
);

CKINVDCx20_ASAP7_75t_R g72 ( 
.A(n_67),
.Y(n_72)
);

CKINVDCx20_ASAP7_75t_R g110 ( 
.A(n_72),
.Y(n_110)
);

AOI22xp5_ASAP7_75t_L g74 ( 
.A1(n_52),
.A2(n_33),
.B1(n_21),
.B2(n_28),
.Y(n_74)
);

OAI22xp5_ASAP7_75t_SL g109 ( 
.A1(n_74),
.A2(n_51),
.B1(n_54),
.B2(n_62),
.Y(n_109)
);

CKINVDCx20_ASAP7_75t_R g76 ( 
.A(n_46),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_L g78 ( 
.A(n_66),
.B(n_27),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_L g94 ( 
.A(n_78),
.B(n_84),
.Y(n_94)
);

INVx2_ASAP7_75t_L g79 ( 
.A(n_46),
.Y(n_79)
);

INVx2_ASAP7_75t_L g98 ( 
.A(n_79),
.Y(n_98)
);

CKINVDCx14_ASAP7_75t_R g92 ( 
.A(n_81),
.Y(n_92)
);

INVx2_ASAP7_75t_L g83 ( 
.A(n_46),
.Y(n_83)
);

INVx2_ASAP7_75t_L g101 ( 
.A(n_83),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_L g84 ( 
.A(n_66),
.B(n_21),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g85 ( 
.A(n_47),
.B(n_21),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_L g103 ( 
.A(n_85),
.B(n_61),
.Y(n_103)
);

AOI22xp33_ASAP7_75t_L g86 ( 
.A1(n_53),
.A2(n_63),
.B1(n_68),
.B2(n_52),
.Y(n_86)
);

OAI22xp5_ASAP7_75t_L g99 ( 
.A1(n_86),
.A2(n_50),
.B1(n_68),
.B2(n_64),
.Y(n_99)
);

INVx3_ASAP7_75t_L g87 ( 
.A(n_56),
.Y(n_87)
);

BUFx6f_ASAP7_75t_L g97 ( 
.A(n_87),
.Y(n_97)
);

OAI22xp33_ASAP7_75t_SL g91 ( 
.A1(n_88),
.A2(n_62),
.B1(n_54),
.B2(n_58),
.Y(n_91)
);

AOI22xp5_ASAP7_75t_L g127 ( 
.A1(n_91),
.A2(n_99),
.B1(n_109),
.B2(n_83),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_77),
.B(n_55),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_SL g116 ( 
.A(n_93),
.B(n_95),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_77),
.B(n_48),
.Y(n_95)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_82),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_SL g131 ( 
.A(n_96),
.B(n_100),
.Y(n_131)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_82),
.Y(n_100)
);

INVx2_ASAP7_75t_L g102 ( 
.A(n_79),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_L g122 ( 
.A(n_102),
.B(n_106),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_L g125 ( 
.A(n_103),
.B(n_111),
.Y(n_125)
);

OAI21xp5_ASAP7_75t_SL g104 ( 
.A1(n_75),
.A2(n_61),
.B(n_64),
.Y(n_104)
);

OAI21xp5_ASAP7_75t_L g117 ( 
.A1(n_104),
.A2(n_75),
.B(n_73),
.Y(n_117)
);

MAJIxp5_ASAP7_75t_L g105 ( 
.A(n_85),
.B(n_70),
.C(n_71),
.Y(n_105)
);

MAJx2_ASAP7_75t_L g120 ( 
.A(n_105),
.B(n_73),
.C(n_84),
.Y(n_120)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_82),
.Y(n_106)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_74),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_L g132 ( 
.A(n_107),
.B(n_112),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_71),
.B(n_12),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_SL g133 ( 
.A(n_108),
.B(n_14),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_SL g111 ( 
.A(n_78),
.B(n_22),
.Y(n_111)
);

CKINVDCx16_ASAP7_75t_R g112 ( 
.A(n_88),
.Y(n_112)
);

AOI22xp33_ASAP7_75t_SL g113 ( 
.A1(n_110),
.A2(n_80),
.B1(n_72),
.B2(n_49),
.Y(n_113)
);

OAI22xp5_ASAP7_75t_L g140 ( 
.A1(n_113),
.A2(n_127),
.B1(n_96),
.B2(n_101),
.Y(n_140)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_90),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g142 ( 
.A(n_114),
.B(n_115),
.Y(n_142)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_109),
.Y(n_115)
);

XOR2xp5_ASAP7_75t_L g134 ( 
.A(n_117),
.B(n_121),
.Y(n_134)
);

AOI22x1_ASAP7_75t_L g118 ( 
.A1(n_92),
.A2(n_80),
.B1(n_86),
.B2(n_81),
.Y(n_118)
);

OA22x2_ASAP7_75t_L g137 ( 
.A1(n_118),
.A2(n_104),
.B1(n_107),
.B2(n_111),
.Y(n_137)
);

AND2x2_ASAP7_75t_L g119 ( 
.A(n_99),
.B(n_70),
.Y(n_119)
);

OAI21xp5_ASAP7_75t_SL g141 ( 
.A1(n_119),
.A2(n_38),
.B(n_32),
.Y(n_141)
);

MAJIxp5_ASAP7_75t_L g149 ( 
.A(n_120),
.B(n_23),
.C(n_17),
.Y(n_149)
);

XNOR2xp5_ASAP7_75t_SL g121 ( 
.A(n_105),
.B(n_74),
.Y(n_121)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_110),
.Y(n_123)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_123),
.Y(n_143)
);

BUFx2_ASAP7_75t_L g124 ( 
.A(n_97),
.Y(n_124)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_124),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_L g126 ( 
.A(n_94),
.B(n_76),
.Y(n_126)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_126),
.Y(n_135)
);

OAI22xp5_ASAP7_75t_L g128 ( 
.A1(n_112),
.A2(n_89),
.B1(n_87),
.B2(n_49),
.Y(n_128)
);

AOI22xp5_ASAP7_75t_L g146 ( 
.A1(n_128),
.A2(n_102),
.B1(n_101),
.B2(n_98),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_L g129 ( 
.A(n_94),
.B(n_89),
.Y(n_129)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_129),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_L g130 ( 
.A(n_103),
.B(n_87),
.Y(n_130)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_130),
.Y(n_138)
);

INVx1_ASAP7_75t_SL g147 ( 
.A(n_133),
.Y(n_147)
);

CKINVDCx14_ASAP7_75t_R g154 ( 
.A(n_137),
.Y(n_154)
);

AOI21xp5_ASAP7_75t_L g139 ( 
.A1(n_119),
.A2(n_106),
.B(n_100),
.Y(n_139)
);

OAI21xp5_ASAP7_75t_SL g155 ( 
.A1(n_139),
.A2(n_140),
.B(n_141),
.Y(n_155)
);

AOI21xp5_ASAP7_75t_L g144 ( 
.A1(n_119),
.A2(n_97),
.B(n_1),
.Y(n_144)
);

OAI21xp5_ASAP7_75t_L g160 ( 
.A1(n_144),
.A2(n_153),
.B(n_129),
.Y(n_160)
);

OAI22xp5_ASAP7_75t_L g168 ( 
.A1(n_146),
.A2(n_38),
.B1(n_23),
.B2(n_17),
.Y(n_168)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_122),
.Y(n_148)
);

NOR2xp33_ASAP7_75t_L g162 ( 
.A(n_148),
.B(n_150),
.Y(n_162)
);

MAJIxp5_ASAP7_75t_L g157 ( 
.A(n_149),
.B(n_151),
.C(n_120),
.Y(n_157)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_131),
.Y(n_150)
);

MAJIxp5_ASAP7_75t_L g151 ( 
.A(n_121),
.B(n_98),
.C(n_97),
.Y(n_151)
);

OAI22xp5_ASAP7_75t_SL g152 ( 
.A1(n_118),
.A2(n_115),
.B1(n_132),
.B2(n_127),
.Y(n_152)
);

AOI22xp5_ASAP7_75t_L g165 ( 
.A1(n_152),
.A2(n_126),
.B1(n_125),
.B2(n_124),
.Y(n_165)
);

AOI22xp5_ASAP7_75t_SL g153 ( 
.A1(n_118),
.A2(n_114),
.B1(n_123),
.B2(n_117),
.Y(n_153)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_142),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_L g177 ( 
.A(n_156),
.B(n_159),
.Y(n_177)
);

MAJIxp5_ASAP7_75t_L g173 ( 
.A(n_157),
.B(n_158),
.C(n_149),
.Y(n_173)
);

MAJIxp5_ASAP7_75t_L g158 ( 
.A(n_151),
.B(n_130),
.C(n_125),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_L g159 ( 
.A(n_135),
.B(n_136),
.Y(n_159)
);

OAI22xp5_ASAP7_75t_L g176 ( 
.A1(n_160),
.A2(n_165),
.B1(n_137),
.B2(n_141),
.Y(n_176)
);

NOR2xp33_ASAP7_75t_SL g161 ( 
.A(n_142),
.B(n_116),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_SL g175 ( 
.A(n_161),
.B(n_164),
.Y(n_175)
);

CKINVDCx20_ASAP7_75t_R g163 ( 
.A(n_143),
.Y(n_163)
);

CKINVDCx20_ASAP7_75t_R g186 ( 
.A(n_163),
.Y(n_186)
);

CKINVDCx16_ASAP7_75t_R g164 ( 
.A(n_146),
.Y(n_164)
);

CKINVDCx20_ASAP7_75t_R g166 ( 
.A(n_143),
.Y(n_166)
);

NOR2xp33_ASAP7_75t_L g181 ( 
.A(n_166),
.B(n_167),
.Y(n_181)
);

CKINVDCx20_ASAP7_75t_R g167 ( 
.A(n_139),
.Y(n_167)
);

AOI22xp5_ASAP7_75t_L g182 ( 
.A1(n_168),
.A2(n_170),
.B1(n_23),
.B2(n_147),
.Y(n_182)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_152),
.Y(n_169)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_169),
.Y(n_179)
);

OAI22xp5_ASAP7_75t_SL g170 ( 
.A1(n_153),
.A2(n_23),
.B1(n_22),
.B2(n_38),
.Y(n_170)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_144),
.Y(n_171)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_171),
.Y(n_183)
);

XOR2xp5_ASAP7_75t_L g172 ( 
.A(n_157),
.B(n_134),
.Y(n_172)
);

XNOR2xp5_ASAP7_75t_L g191 ( 
.A(n_172),
.B(n_159),
.Y(n_191)
);

MAJIxp5_ASAP7_75t_L g192 ( 
.A(n_173),
.B(n_174),
.C(n_178),
.Y(n_192)
);

MAJIxp5_ASAP7_75t_L g174 ( 
.A(n_158),
.B(n_134),
.C(n_138),
.Y(n_174)
);

AOI22xp5_ASAP7_75t_L g190 ( 
.A1(n_176),
.A2(n_169),
.B1(n_171),
.B2(n_155),
.Y(n_190)
);

MAJIxp5_ASAP7_75t_L g178 ( 
.A(n_156),
.B(n_137),
.C(n_145),
.Y(n_178)
);

AOI22xp5_ASAP7_75t_SL g180 ( 
.A1(n_170),
.A2(n_137),
.B1(n_145),
.B2(n_147),
.Y(n_180)
);

OAI22xp5_ASAP7_75t_SL g188 ( 
.A1(n_180),
.A2(n_182),
.B1(n_154),
.B2(n_160),
.Y(n_188)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_162),
.Y(n_184)
);

NOR2xp33_ASAP7_75t_L g193 ( 
.A(n_184),
.B(n_161),
.Y(n_193)
);

MAJIxp5_ASAP7_75t_L g185 ( 
.A(n_165),
.B(n_22),
.C(n_1),
.Y(n_185)
);

MAJIxp5_ASAP7_75t_L g194 ( 
.A(n_185),
.B(n_155),
.C(n_168),
.Y(n_194)
);

A2O1A1Ixp33_ASAP7_75t_SL g187 ( 
.A1(n_178),
.A2(n_167),
.B(n_166),
.C(n_163),
.Y(n_187)
);

OAI21xp5_ASAP7_75t_SL g198 ( 
.A1(n_187),
.A2(n_196),
.B(n_180),
.Y(n_198)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_188),
.Y(n_199)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_177),
.Y(n_189)
);

NOR2xp33_ASAP7_75t_L g201 ( 
.A(n_189),
.B(n_190),
.Y(n_201)
);

MAJIxp5_ASAP7_75t_L g202 ( 
.A(n_191),
.B(n_194),
.C(n_22),
.Y(n_202)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_193),
.Y(n_205)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_181),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_L g204 ( 
.A(n_195),
.B(n_3),
.Y(n_204)
);

AOI21xp5_ASAP7_75t_L g196 ( 
.A1(n_175),
.A2(n_0),
.B(n_2),
.Y(n_196)
);

NOR2xp33_ASAP7_75t_L g197 ( 
.A(n_186),
.B(n_3),
.Y(n_197)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_197),
.Y(n_206)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_198),
.Y(n_207)
);

AOI322xp5_ASAP7_75t_L g200 ( 
.A1(n_194),
.A2(n_174),
.A3(n_173),
.B1(n_185),
.B2(n_183),
.C1(n_179),
.C2(n_172),
.Y(n_200)
);

OAI21xp5_ASAP7_75t_L g212 ( 
.A1(n_200),
.A2(n_202),
.B(n_203),
.Y(n_212)
);

A2O1A1Ixp33_ASAP7_75t_L g203 ( 
.A1(n_187),
.A2(n_3),
.B(n_4),
.C(n_6),
.Y(n_203)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_204),
.Y(n_213)
);

AOI21xp5_ASAP7_75t_L g208 ( 
.A1(n_201),
.A2(n_187),
.B(n_191),
.Y(n_208)
);

OAI321xp33_ASAP7_75t_L g216 ( 
.A1(n_208),
.A2(n_209),
.A3(n_203),
.B1(n_7),
.B2(n_8),
.C(n_9),
.Y(n_216)
);

AOI22xp33_ASAP7_75t_SL g209 ( 
.A1(n_199),
.A2(n_187),
.B1(n_192),
.B2(n_8),
.Y(n_209)
);

INVxp67_ASAP7_75t_L g210 ( 
.A(n_204),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_L g217 ( 
.A(n_210),
.B(n_211),
.Y(n_217)
);

NAND2xp5_ASAP7_75t_L g211 ( 
.A(n_205),
.B(n_206),
.Y(n_211)
);

MAJIxp5_ASAP7_75t_L g214 ( 
.A(n_212),
.B(n_192),
.C(n_202),
.Y(n_214)
);

OAI21xp5_ASAP7_75t_L g221 ( 
.A1(n_214),
.A2(n_8),
.B(n_10),
.Y(n_221)
);

XOR2xp5_ASAP7_75t_L g215 ( 
.A(n_207),
.B(n_198),
.Y(n_215)
);

MAJx2_ASAP7_75t_L g220 ( 
.A(n_215),
.B(n_218),
.C(n_7),
.Y(n_220)
);

AOI21xp5_ASAP7_75t_SL g219 ( 
.A1(n_216),
.A2(n_4),
.B(n_7),
.Y(n_219)
);

XNOR2xp5_ASAP7_75t_L g218 ( 
.A(n_213),
.B(n_209),
.Y(n_218)
);

INVxp67_ASAP7_75t_L g222 ( 
.A(n_219),
.Y(n_222)
);

A2O1A1Ixp33_ASAP7_75t_L g223 ( 
.A1(n_220),
.A2(n_221),
.B(n_217),
.C(n_11),
.Y(n_223)
);

AO21x1_ASAP7_75t_SL g224 ( 
.A1(n_223),
.A2(n_215),
.B(n_10),
.Y(n_224)
);

MAJIxp5_ASAP7_75t_L g225 ( 
.A(n_224),
.B(n_222),
.C(n_10),
.Y(n_225)
);

XOR2xp5_ASAP7_75t_L g226 ( 
.A(n_225),
.B(n_11),
.Y(n_226)
);


endmodule