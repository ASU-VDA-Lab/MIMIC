module fake_jpeg_8874_n_229 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_229);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_229;

wire n_159;
wire n_117;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_84;
wire n_59;
wire n_98;
wire n_178;
wire n_228;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_223;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_44;
wire n_24;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_131;
wire n_56;
wire n_212;
wire n_211;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_216;
wire n_217;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

BUFx5_ASAP7_75t_L g16 ( 
.A(n_6),
.Y(n_16)
);

INVx2_ASAP7_75t_L g17 ( 
.A(n_3),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_9),
.Y(n_18)
);

INVx2_ASAP7_75t_L g19 ( 
.A(n_15),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_12),
.Y(n_20)
);

BUFx12f_ASAP7_75t_L g21 ( 
.A(n_9),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_9),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_3),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_10),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_8),
.Y(n_25)
);

BUFx3_ASAP7_75t_L g26 ( 
.A(n_3),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_14),
.Y(n_27)
);

BUFx5_ASAP7_75t_L g28 ( 
.A(n_6),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_14),
.Y(n_29)
);

BUFx3_ASAP7_75t_L g30 ( 
.A(n_15),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_2),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_6),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_4),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_21),
.Y(n_34)
);

INVx3_ASAP7_75t_L g61 ( 
.A(n_34),
.Y(n_61)
);

INVx2_ASAP7_75t_L g35 ( 
.A(n_16),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_35),
.B(n_37),
.Y(n_50)
);

INVx8_ASAP7_75t_L g36 ( 
.A(n_16),
.Y(n_36)
);

INVx3_ASAP7_75t_SL g64 ( 
.A(n_36),
.Y(n_64)
);

INVx4_ASAP7_75t_SL g37 ( 
.A(n_22),
.Y(n_37)
);

INVx6_ASAP7_75t_L g38 ( 
.A(n_22),
.Y(n_38)
);

INVx8_ASAP7_75t_L g47 ( 
.A(n_38),
.Y(n_47)
);

INVx3_ASAP7_75t_L g39 ( 
.A(n_22),
.Y(n_39)
);

INVx4_ASAP7_75t_L g51 ( 
.A(n_39),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_21),
.Y(n_40)
);

INVx3_ASAP7_75t_L g62 ( 
.A(n_40),
.Y(n_62)
);

INVx8_ASAP7_75t_L g41 ( 
.A(n_28),
.Y(n_41)
);

AOI22xp33_ASAP7_75t_SL g49 ( 
.A1(n_41),
.A2(n_19),
.B1(n_17),
.B2(n_28),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_21),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_42),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g43 ( 
.A(n_19),
.B(n_0),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_SL g52 ( 
.A(n_43),
.B(n_45),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_21),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_44),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g45 ( 
.A(n_27),
.B(n_0),
.Y(n_45)
);

AOI22xp5_ASAP7_75t_SL g46 ( 
.A1(n_38),
.A2(n_18),
.B1(n_32),
.B2(n_23),
.Y(n_46)
);

OAI22xp5_ASAP7_75t_SL g73 ( 
.A1(n_46),
.A2(n_56),
.B1(n_58),
.B2(n_59),
.Y(n_73)
);

INVxp67_ASAP7_75t_L g75 ( 
.A(n_49),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_L g53 ( 
.A(n_43),
.B(n_17),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_L g71 ( 
.A(n_53),
.B(n_29),
.Y(n_71)
);

BUFx3_ASAP7_75t_L g54 ( 
.A(n_34),
.Y(n_54)
);

INVx3_ASAP7_75t_L g88 ( 
.A(n_54),
.Y(n_88)
);

AO22x1_ASAP7_75t_SL g55 ( 
.A1(n_38),
.A2(n_39),
.B1(n_37),
.B2(n_40),
.Y(n_55)
);

AOI22xp5_ASAP7_75t_L g83 ( 
.A1(n_55),
.A2(n_44),
.B1(n_42),
.B2(n_26),
.Y(n_83)
);

OAI22xp5_ASAP7_75t_L g56 ( 
.A1(n_37),
.A2(n_18),
.B1(n_32),
.B2(n_25),
.Y(n_56)
);

AOI22xp33_ASAP7_75t_SL g57 ( 
.A1(n_36),
.A2(n_20),
.B1(n_31),
.B2(n_33),
.Y(n_57)
);

INVxp67_ASAP7_75t_L g81 ( 
.A(n_57),
.Y(n_81)
);

AOI22xp33_ASAP7_75t_L g58 ( 
.A1(n_36),
.A2(n_23),
.B1(n_24),
.B2(n_25),
.Y(n_58)
);

AOI22xp33_ASAP7_75t_SL g59 ( 
.A1(n_41),
.A2(n_20),
.B1(n_31),
.B2(n_33),
.Y(n_59)
);

INVx2_ASAP7_75t_L g63 ( 
.A(n_34),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_63),
.B(n_35),
.Y(n_68)
);

INVx4_ASAP7_75t_L g65 ( 
.A(n_40),
.Y(n_65)
);

INVx1_ASAP7_75t_SL g76 ( 
.A(n_65),
.Y(n_76)
);

CKINVDCx20_ASAP7_75t_R g66 ( 
.A(n_42),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_SL g84 ( 
.A(n_66),
.B(n_1),
.Y(n_84)
);

AOI22xp5_ASAP7_75t_SL g67 ( 
.A1(n_41),
.A2(n_24),
.B1(n_29),
.B2(n_27),
.Y(n_67)
);

OAI22xp5_ASAP7_75t_SL g78 ( 
.A1(n_67),
.A2(n_30),
.B1(n_26),
.B2(n_4),
.Y(n_78)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_68),
.Y(n_94)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_56),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_69),
.B(n_70),
.Y(n_93)
);

INVx4_ASAP7_75t_L g70 ( 
.A(n_65),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_SL g104 ( 
.A(n_71),
.B(n_82),
.Y(n_104)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_50),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_72),
.B(n_74),
.Y(n_96)
);

INVx2_ASAP7_75t_L g74 ( 
.A(n_64),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_52),
.B(n_0),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_77),
.B(n_79),
.Y(n_99)
);

AOI22xp5_ASAP7_75t_L g108 ( 
.A1(n_78),
.A2(n_83),
.B1(n_87),
.B2(n_51),
.Y(n_108)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_50),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_L g80 ( 
.A(n_53),
.B(n_44),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_L g98 ( 
.A(n_80),
.B(n_90),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_SL g82 ( 
.A(n_52),
.B(n_67),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_84),
.B(n_85),
.Y(n_103)
);

INVx2_ASAP7_75t_L g85 ( 
.A(n_64),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_66),
.B(n_46),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g112 ( 
.A(n_86),
.B(n_89),
.Y(n_112)
);

OAI22xp5_ASAP7_75t_SL g87 ( 
.A1(n_55),
.A2(n_26),
.B1(n_30),
.B2(n_4),
.Y(n_87)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_55),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g90 ( 
.A(n_55),
.B(n_1),
.Y(n_90)
);

HB1xp67_ASAP7_75t_L g91 ( 
.A(n_76),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g126 ( 
.A(n_91),
.B(n_101),
.Y(n_126)
);

INVxp67_ASAP7_75t_L g92 ( 
.A(n_83),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_SL g117 ( 
.A(n_92),
.B(n_102),
.Y(n_117)
);

AOI22xp5_ASAP7_75t_SL g95 ( 
.A1(n_75),
.A2(n_64),
.B1(n_47),
.B2(n_62),
.Y(n_95)
);

OAI22xp5_ASAP7_75t_L g124 ( 
.A1(n_95),
.A2(n_107),
.B1(n_108),
.B2(n_70),
.Y(n_124)
);

MAJIxp5_ASAP7_75t_L g97 ( 
.A(n_80),
.B(n_47),
.C(n_63),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g118 ( 
.A(n_97),
.B(n_100),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_L g100 ( 
.A(n_71),
.B(n_60),
.Y(n_100)
);

HB1xp67_ASAP7_75t_L g101 ( 
.A(n_76),
.Y(n_101)
);

CKINVDCx16_ASAP7_75t_R g102 ( 
.A(n_90),
.Y(n_102)
);

AOI21xp5_ASAP7_75t_L g105 ( 
.A1(n_81),
.A2(n_75),
.B(n_89),
.Y(n_105)
);

AOI21xp5_ASAP7_75t_L g133 ( 
.A1(n_105),
.A2(n_2),
.B(n_5),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_L g106 ( 
.A(n_72),
.B(n_60),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_L g129 ( 
.A(n_106),
.B(n_111),
.Y(n_129)
);

AOI22xp33_ASAP7_75t_SL g107 ( 
.A1(n_69),
.A2(n_47),
.B1(n_51),
.B2(n_61),
.Y(n_107)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_87),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_L g130 ( 
.A(n_109),
.B(n_110),
.Y(n_130)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_74),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_SL g111 ( 
.A(n_79),
.B(n_65),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_L g113 ( 
.A(n_85),
.B(n_62),
.Y(n_113)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_113),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_L g114 ( 
.A(n_73),
.B(n_61),
.Y(n_114)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_114),
.Y(n_121)
);

CKINVDCx20_ASAP7_75t_R g115 ( 
.A(n_106),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_SL g154 ( 
.A(n_115),
.B(n_120),
.Y(n_154)
);

OAI22xp5_ASAP7_75t_SL g119 ( 
.A1(n_109),
.A2(n_81),
.B1(n_73),
.B2(n_78),
.Y(n_119)
);

OAI22xp5_ASAP7_75t_SL g137 ( 
.A1(n_119),
.A2(n_131),
.B1(n_95),
.B2(n_112),
.Y(n_137)
);

CKINVDCx20_ASAP7_75t_R g120 ( 
.A(n_99),
.Y(n_120)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_113),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_L g148 ( 
.A(n_122),
.B(n_123),
.Y(n_148)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_96),
.Y(n_123)
);

A2O1A1Ixp33_ASAP7_75t_SL g141 ( 
.A1(n_124),
.A2(n_133),
.B(n_112),
.C(n_93),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_SL g125 ( 
.A(n_99),
.B(n_13),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_L g151 ( 
.A(n_125),
.B(n_134),
.Y(n_151)
);

OAI22xp5_ASAP7_75t_L g127 ( 
.A1(n_108),
.A2(n_88),
.B1(n_60),
.B2(n_48),
.Y(n_127)
);

O2A1O1Ixp33_ASAP7_75t_L g144 ( 
.A1(n_127),
.A2(n_128),
.B(n_110),
.C(n_100),
.Y(n_144)
);

OAI22xp5_ASAP7_75t_L g128 ( 
.A1(n_114),
.A2(n_88),
.B1(n_48),
.B2(n_54),
.Y(n_128)
);

AOI22xp5_ASAP7_75t_L g131 ( 
.A1(n_102),
.A2(n_48),
.B1(n_54),
.B2(n_5),
.Y(n_131)
);

AOI22xp5_ASAP7_75t_SL g132 ( 
.A1(n_105),
.A2(n_1),
.B1(n_2),
.B2(n_5),
.Y(n_132)
);

INVxp67_ASAP7_75t_L g140 ( 
.A(n_132),
.Y(n_140)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_96),
.Y(n_134)
);

CKINVDCx20_ASAP7_75t_R g135 ( 
.A(n_93),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_L g145 ( 
.A(n_135),
.B(n_136),
.Y(n_145)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_111),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_SL g167 ( 
.A(n_137),
.B(n_144),
.Y(n_167)
);

HB1xp67_ASAP7_75t_L g138 ( 
.A(n_126),
.Y(n_138)
);

INVxp67_ASAP7_75t_SL g159 ( 
.A(n_138),
.Y(n_159)
);

XNOR2xp5_ASAP7_75t_L g139 ( 
.A(n_118),
.B(n_98),
.Y(n_139)
);

MAJIxp5_ASAP7_75t_L g168 ( 
.A(n_139),
.B(n_143),
.C(n_152),
.Y(n_168)
);

AOI21xp5_ASAP7_75t_SL g163 ( 
.A1(n_141),
.A2(n_135),
.B(n_122),
.Y(n_163)
);

INVx2_ASAP7_75t_L g142 ( 
.A(n_131),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_L g170 ( 
.A(n_142),
.B(n_146),
.Y(n_170)
);

MAJIxp5_ASAP7_75t_L g143 ( 
.A(n_118),
.B(n_97),
.C(n_98),
.Y(n_143)
);

CKINVDCx20_ASAP7_75t_R g146 ( 
.A(n_130),
.Y(n_146)
);

CKINVDCx20_ASAP7_75t_R g147 ( 
.A(n_129),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_SL g158 ( 
.A(n_147),
.B(n_150),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_L g149 ( 
.A(n_129),
.B(n_104),
.Y(n_149)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_149),
.Y(n_161)
);

CKINVDCx14_ASAP7_75t_R g150 ( 
.A(n_117),
.Y(n_150)
);

MAJIxp5_ASAP7_75t_L g152 ( 
.A(n_115),
.B(n_136),
.C(n_121),
.Y(n_152)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_123),
.Y(n_153)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_153),
.Y(n_172)
);

INVxp67_ASAP7_75t_L g155 ( 
.A(n_132),
.Y(n_155)
);

INVxp67_ASAP7_75t_L g165 ( 
.A(n_155),
.Y(n_165)
);

CKINVDCx20_ASAP7_75t_R g156 ( 
.A(n_133),
.Y(n_156)
);

NOR2xp33_ASAP7_75t_SL g160 ( 
.A(n_156),
.B(n_121),
.Y(n_160)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_134),
.Y(n_157)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_157),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_SL g184 ( 
.A(n_160),
.B(n_162),
.Y(n_184)
);

BUFx6f_ASAP7_75t_L g162 ( 
.A(n_148),
.Y(n_162)
);

XNOR2xp5_ASAP7_75t_L g178 ( 
.A(n_163),
.B(n_137),
.Y(n_178)
);

AND2x2_ASAP7_75t_L g164 ( 
.A(n_152),
.B(n_116),
.Y(n_164)
);

AOI21xp5_ASAP7_75t_L g185 ( 
.A1(n_164),
.A2(n_116),
.B(n_141),
.Y(n_185)
);

MAJIxp5_ASAP7_75t_L g166 ( 
.A(n_143),
.B(n_120),
.C(n_104),
.Y(n_166)
);

MAJIxp5_ASAP7_75t_L g183 ( 
.A(n_166),
.B(n_169),
.C(n_171),
.Y(n_183)
);

XNOR2xp5_ASAP7_75t_SL g169 ( 
.A(n_139),
.B(n_119),
.Y(n_169)
);

MAJIxp5_ASAP7_75t_L g171 ( 
.A(n_149),
.B(n_145),
.C(n_154),
.Y(n_171)
);

XNOR2xp5_ASAP7_75t_L g173 ( 
.A(n_145),
.B(n_103),
.Y(n_173)
);

MAJIxp5_ASAP7_75t_L g189 ( 
.A(n_173),
.B(n_101),
.C(n_91),
.Y(n_189)
);

CKINVDCx20_ASAP7_75t_R g174 ( 
.A(n_151),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_L g179 ( 
.A(n_174),
.B(n_153),
.Y(n_179)
);

NOR2xp33_ASAP7_75t_L g176 ( 
.A(n_159),
.B(n_157),
.Y(n_176)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_176),
.Y(n_192)
);

OAI22xp5_ASAP7_75t_SL g177 ( 
.A1(n_167),
.A2(n_155),
.B1(n_140),
.B2(n_141),
.Y(n_177)
);

AOI22xp5_ASAP7_75t_L g193 ( 
.A1(n_177),
.A2(n_169),
.B1(n_164),
.B2(n_168),
.Y(n_193)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_178),
.Y(n_199)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_179),
.Y(n_196)
);

INVx2_ASAP7_75t_L g180 ( 
.A(n_159),
.Y(n_180)
);

CKINVDCx20_ASAP7_75t_R g194 ( 
.A(n_180),
.Y(n_194)
);

OAI22xp5_ASAP7_75t_L g181 ( 
.A1(n_170),
.A2(n_142),
.B1(n_140),
.B2(n_141),
.Y(n_181)
);

OAI22xp5_ASAP7_75t_L g191 ( 
.A1(n_181),
.A2(n_185),
.B1(n_186),
.B2(n_190),
.Y(n_191)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_158),
.Y(n_182)
);

NOR2xp33_ASAP7_75t_SL g201 ( 
.A(n_182),
.B(n_188),
.Y(n_201)
);

AOI22xp5_ASAP7_75t_L g186 ( 
.A1(n_165),
.A2(n_144),
.B1(n_103),
.B2(n_94),
.Y(n_186)
);

INVxp67_ASAP7_75t_L g187 ( 
.A(n_163),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_L g197 ( 
.A(n_187),
.B(n_188),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_L g188 ( 
.A(n_161),
.B(n_94),
.Y(n_188)
);

MAJIxp5_ASAP7_75t_L g195 ( 
.A(n_189),
.B(n_168),
.C(n_162),
.Y(n_195)
);

OAI22xp5_ASAP7_75t_L g190 ( 
.A1(n_165),
.A2(n_175),
.B1(n_172),
.B2(n_171),
.Y(n_190)
);

OAI22xp5_ASAP7_75t_SL g208 ( 
.A1(n_193),
.A2(n_198),
.B1(n_186),
.B2(n_8),
.Y(n_208)
);

MAJIxp5_ASAP7_75t_L g202 ( 
.A(n_195),
.B(n_183),
.C(n_189),
.Y(n_202)
);

AOI22xp5_ASAP7_75t_SL g198 ( 
.A1(n_187),
.A2(n_7),
.B1(n_8),
.B2(n_10),
.Y(n_198)
);

INVx3_ASAP7_75t_L g200 ( 
.A(n_180),
.Y(n_200)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_200),
.Y(n_206)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_201),
.Y(n_207)
);

NAND2xp5_ASAP7_75t_L g214 ( 
.A(n_202),
.B(n_205),
.Y(n_214)
);

NAND2xp5_ASAP7_75t_L g203 ( 
.A(n_192),
.B(n_184),
.Y(n_203)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_203),
.Y(n_212)
);

AOI22xp5_ASAP7_75t_L g204 ( 
.A1(n_199),
.A2(n_177),
.B1(n_178),
.B2(n_185),
.Y(n_204)
);

OAI22xp5_ASAP7_75t_SL g213 ( 
.A1(n_204),
.A2(n_196),
.B1(n_194),
.B2(n_200),
.Y(n_213)
);

MAJIxp5_ASAP7_75t_L g205 ( 
.A(n_195),
.B(n_193),
.C(n_183),
.Y(n_205)
);

A2O1A1Ixp33_ASAP7_75t_SL g211 ( 
.A1(n_208),
.A2(n_191),
.B(n_198),
.C(n_196),
.Y(n_211)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_197),
.Y(n_209)
);

NOR2xp33_ASAP7_75t_L g210 ( 
.A(n_209),
.B(n_197),
.Y(n_210)
);

NOR2xp33_ASAP7_75t_L g217 ( 
.A(n_210),
.B(n_213),
.Y(n_217)
);

AO21x1_ASAP7_75t_L g220 ( 
.A1(n_211),
.A2(n_215),
.B(n_7),
.Y(n_220)
);

NAND2xp5_ASAP7_75t_L g215 ( 
.A(n_207),
.B(n_7),
.Y(n_215)
);

AO21x1_ASAP7_75t_L g216 ( 
.A1(n_208),
.A2(n_13),
.B(n_10),
.Y(n_216)
);

NOR2xp33_ASAP7_75t_L g221 ( 
.A(n_216),
.B(n_11),
.Y(n_221)
);

OAI22xp5_ASAP7_75t_SL g218 ( 
.A1(n_214),
.A2(n_204),
.B1(n_202),
.B2(n_205),
.Y(n_218)
);

NAND2xp5_ASAP7_75t_L g223 ( 
.A(n_218),
.B(n_219),
.Y(n_223)
);

OAI22xp5_ASAP7_75t_SL g219 ( 
.A1(n_212),
.A2(n_206),
.B1(n_11),
.B2(n_12),
.Y(n_219)
);

XOR2xp5_ASAP7_75t_L g224 ( 
.A(n_220),
.B(n_11),
.Y(n_224)
);

OAI21xp5_ASAP7_75t_L g222 ( 
.A1(n_221),
.A2(n_215),
.B(n_211),
.Y(n_222)
);

XOR2xp5_ASAP7_75t_L g225 ( 
.A(n_222),
.B(n_219),
.Y(n_225)
);

AND2x2_ASAP7_75t_L g226 ( 
.A(n_224),
.B(n_12),
.Y(n_226)
);

MAJIxp5_ASAP7_75t_L g227 ( 
.A(n_225),
.B(n_226),
.C(n_223),
.Y(n_227)
);

AOI21xp5_ASAP7_75t_SL g228 ( 
.A1(n_227),
.A2(n_217),
.B(n_218),
.Y(n_228)
);

XOR2xp5_ASAP7_75t_L g229 ( 
.A(n_228),
.B(n_220),
.Y(n_229)
);


endmodule