module fake_netlist_6_29_n_2039 (n_52, n_16, n_1, n_91, n_119, n_46, n_146, n_163, n_18, n_21, n_193, n_147, n_154, n_191, n_88, n_3, n_98, n_113, n_39, n_63, n_73, n_4, n_148, n_199, n_138, n_22, n_161, n_208, n_68, n_166, n_28, n_184, n_50, n_158, n_49, n_7, n_83, n_206, n_5, n_101, n_167, n_144, n_174, n_127, n_125, n_153, n_168, n_178, n_77, n_156, n_149, n_152, n_106, n_92, n_145, n_42, n_133, n_96, n_8, n_90, n_160, n_24, n_105, n_131, n_54, n_132, n_188, n_102, n_186, n_204, n_0, n_87, n_195, n_189, n_32, n_66, n_85, n_99, n_78, n_84, n_130, n_164, n_100, n_129, n_13, n_121, n_197, n_11, n_137, n_17, n_23, n_203, n_142, n_20, n_143, n_207, n_2, n_180, n_19, n_47, n_62, n_29, n_155, n_75, n_109, n_150, n_122, n_45, n_205, n_34, n_140, n_70, n_120, n_37, n_15, n_67, n_33, n_82, n_27, n_38, n_110, n_151, n_61, n_112, n_172, n_81, n_59, n_181, n_76, n_36, n_182, n_26, n_124, n_55, n_126, n_202, n_94, n_97, n_108, n_58, n_116, n_64, n_117, n_118, n_175, n_48, n_65, n_25, n_40, n_93, n_80, n_141, n_135, n_196, n_200, n_165, n_139, n_41, n_134, n_177, n_176, n_114, n_86, n_198, n_104, n_95, n_179, n_9, n_107, n_10, n_71, n_74, n_6, n_190, n_14, n_123, n_136, n_72, n_187, n_89, n_173, n_201, n_103, n_111, n_60, n_159, n_157, n_162, n_170, n_185, n_35, n_183, n_115, n_12, n_69, n_128, n_30, n_79, n_43, n_194, n_171, n_31, n_192, n_57, n_169, n_53, n_51, n_44, n_56, n_2039);

input n_52;
input n_16;
input n_1;
input n_91;
input n_119;
input n_46;
input n_146;
input n_163;
input n_18;
input n_21;
input n_193;
input n_147;
input n_154;
input n_191;
input n_88;
input n_3;
input n_98;
input n_113;
input n_39;
input n_63;
input n_73;
input n_4;
input n_148;
input n_199;
input n_138;
input n_22;
input n_161;
input n_208;
input n_68;
input n_166;
input n_28;
input n_184;
input n_50;
input n_158;
input n_49;
input n_7;
input n_83;
input n_206;
input n_5;
input n_101;
input n_167;
input n_144;
input n_174;
input n_127;
input n_125;
input n_153;
input n_168;
input n_178;
input n_77;
input n_156;
input n_149;
input n_152;
input n_106;
input n_92;
input n_145;
input n_42;
input n_133;
input n_96;
input n_8;
input n_90;
input n_160;
input n_24;
input n_105;
input n_131;
input n_54;
input n_132;
input n_188;
input n_102;
input n_186;
input n_204;
input n_0;
input n_87;
input n_195;
input n_189;
input n_32;
input n_66;
input n_85;
input n_99;
input n_78;
input n_84;
input n_130;
input n_164;
input n_100;
input n_129;
input n_13;
input n_121;
input n_197;
input n_11;
input n_137;
input n_17;
input n_23;
input n_203;
input n_142;
input n_20;
input n_143;
input n_207;
input n_2;
input n_180;
input n_19;
input n_47;
input n_62;
input n_29;
input n_155;
input n_75;
input n_109;
input n_150;
input n_122;
input n_45;
input n_205;
input n_34;
input n_140;
input n_70;
input n_120;
input n_37;
input n_15;
input n_67;
input n_33;
input n_82;
input n_27;
input n_38;
input n_110;
input n_151;
input n_61;
input n_112;
input n_172;
input n_81;
input n_59;
input n_181;
input n_76;
input n_36;
input n_182;
input n_26;
input n_124;
input n_55;
input n_126;
input n_202;
input n_94;
input n_97;
input n_108;
input n_58;
input n_116;
input n_64;
input n_117;
input n_118;
input n_175;
input n_48;
input n_65;
input n_25;
input n_40;
input n_93;
input n_80;
input n_141;
input n_135;
input n_196;
input n_200;
input n_165;
input n_139;
input n_41;
input n_134;
input n_177;
input n_176;
input n_114;
input n_86;
input n_198;
input n_104;
input n_95;
input n_179;
input n_9;
input n_107;
input n_10;
input n_71;
input n_74;
input n_6;
input n_190;
input n_14;
input n_123;
input n_136;
input n_72;
input n_187;
input n_89;
input n_173;
input n_201;
input n_103;
input n_111;
input n_60;
input n_159;
input n_157;
input n_162;
input n_170;
input n_185;
input n_35;
input n_183;
input n_115;
input n_12;
input n_69;
input n_128;
input n_30;
input n_79;
input n_43;
input n_194;
input n_171;
input n_31;
input n_192;
input n_57;
input n_169;
input n_53;
input n_51;
input n_44;
input n_56;

output n_2039;

wire n_992;
wire n_1671;
wire n_801;
wire n_1613;
wire n_1234;
wire n_1458;
wire n_1199;
wire n_1674;
wire n_741;
wire n_1027;
wire n_1351;
wire n_625;
wire n_1189;
wire n_223;
wire n_1212;
wire n_226;
wire n_726;
wire n_212;
wire n_700;
wire n_1307;
wire n_2003;
wire n_1038;
wire n_578;
wire n_1581;
wire n_1003;
wire n_365;
wire n_1237;
wire n_1061;
wire n_1357;
wire n_1853;
wire n_783;
wire n_1738;
wire n_798;
wire n_1575;
wire n_1854;
wire n_1923;
wire n_509;
wire n_1342;
wire n_245;
wire n_1209;
wire n_1348;
wire n_1387;
wire n_677;
wire n_1708;
wire n_805;
wire n_1151;
wire n_396;
wire n_1739;
wire n_350;
wire n_1380;
wire n_442;
wire n_480;
wire n_1402;
wire n_1688;
wire n_1691;
wire n_1975;
wire n_1009;
wire n_1743;
wire n_1930;
wire n_1160;
wire n_883;
wire n_1238;
wire n_1991;
wire n_1724;
wire n_1032;
wire n_1247;
wire n_1547;
wire n_1553;
wire n_893;
wire n_1099;
wire n_1264;
wire n_1192;
wire n_471;
wire n_1844;
wire n_424;
wire n_1700;
wire n_1555;
wire n_1415;
wire n_1370;
wire n_1786;
wire n_369;
wire n_287;
wire n_415;
wire n_830;
wire n_230;
wire n_461;
wire n_873;
wire n_383;
wire n_1285;
wire n_1371;
wire n_1985;
wire n_447;
wire n_1803;
wire n_1172;
wire n_852;
wire n_229;
wire n_1590;
wire n_1532;
wire n_1393;
wire n_1517;
wire n_1867;
wire n_1704;
wire n_1078;
wire n_250;
wire n_544;
wire n_1711;
wire n_1140;
wire n_1444;
wire n_1670;
wire n_1603;
wire n_1579;
wire n_1263;
wire n_2019;
wire n_836;
wire n_375;
wire n_522;
wire n_1261;
wire n_945;
wire n_1649;
wire n_2018;
wire n_1903;
wire n_1511;
wire n_1143;
wire n_1422;
wire n_1232;
wire n_1772;
wire n_1572;
wire n_658;
wire n_616;
wire n_1874;
wire n_1119;
wire n_2013;
wire n_428;
wire n_1433;
wire n_1902;
wire n_1842;
wire n_1620;
wire n_1954;
wire n_1735;
wire n_1541;
wire n_1300;
wire n_641;
wire n_822;
wire n_693;
wire n_1313;
wire n_1056;
wire n_758;
wire n_516;
wire n_1455;
wire n_1163;
wire n_1180;
wire n_943;
wire n_1798;
wire n_1550;
wire n_491;
wire n_1591;
wire n_772;
wire n_1344;
wire n_666;
wire n_371;
wire n_940;
wire n_770;
wire n_567;
wire n_1781;
wire n_1971;
wire n_405;
wire n_213;
wire n_538;
wire n_2004;
wire n_1106;
wire n_886;
wire n_1471;
wire n_343;
wire n_953;
wire n_1094;
wire n_1345;
wire n_1820;
wire n_494;
wire n_539;
wire n_493;
wire n_454;
wire n_1421;
wire n_1936;
wire n_638;
wire n_1404;
wire n_1211;
wire n_381;
wire n_887;
wire n_1660;
wire n_1961;
wire n_1280;
wire n_713;
wire n_1400;
wire n_1467;
wire n_976;
wire n_224;
wire n_1445;
wire n_1526;
wire n_1560;
wire n_734;
wire n_1088;
wire n_1894;
wire n_1231;
wire n_1978;
wire n_917;
wire n_574;
wire n_907;
wire n_1446;
wire n_659;
wire n_1815;
wire n_407;
wire n_913;
wire n_1658;
wire n_808;
wire n_867;
wire n_1230;
wire n_473;
wire n_1193;
wire n_1967;
wire n_1054;
wire n_559;
wire n_1333;
wire n_1648;
wire n_1911;
wire n_1956;
wire n_1644;
wire n_2011;
wire n_1558;
wire n_1732;
wire n_281;
wire n_551;
wire n_699;
wire n_1986;
wire n_564;
wire n_451;
wire n_824;
wire n_279;
wire n_686;
wire n_757;
wire n_594;
wire n_1641;
wire n_1918;
wire n_577;
wire n_1843;
wire n_619;
wire n_1367;
wire n_1336;
wire n_521;
wire n_572;
wire n_395;
wire n_813;
wire n_1909;
wire n_1481;
wire n_323;
wire n_606;
wire n_1441;
wire n_818;
wire n_1123;
wire n_1309;
wire n_513;
wire n_645;
wire n_1381;
wire n_331;
wire n_1699;
wire n_916;
wire n_483;
wire n_1970;
wire n_608;
wire n_261;
wire n_630;
wire n_541;
wire n_512;
wire n_433;
wire n_792;
wire n_476;
wire n_1328;
wire n_1957;
wire n_219;
wire n_1907;
wire n_264;
wire n_263;
wire n_1162;
wire n_860;
wire n_1530;
wire n_788;
wire n_939;
wire n_1543;
wire n_821;
wire n_938;
wire n_1302;
wire n_1068;
wire n_1599;
wire n_329;
wire n_982;
wire n_549;
wire n_1762;
wire n_1910;
wire n_1075;
wire n_408;
wire n_932;
wire n_237;
wire n_1876;
wire n_1895;
wire n_1697;
wire n_243;
wire n_979;
wire n_1873;
wire n_905;
wire n_1866;
wire n_1680;
wire n_322;
wire n_993;
wire n_689;
wire n_2031;
wire n_354;
wire n_1330;
wire n_1413;
wire n_1605;
wire n_1988;
wire n_1278;
wire n_547;
wire n_558;
wire n_1064;
wire n_1396;
wire n_634;
wire n_966;
wire n_764;
wire n_1663;
wire n_2009;
wire n_692;
wire n_733;
wire n_1793;
wire n_1233;
wire n_1289;
wire n_487;
wire n_241;
wire n_1107;
wire n_1014;
wire n_1290;
wire n_1703;
wire n_882;
wire n_1354;
wire n_586;
wire n_423;
wire n_1865;
wire n_1875;
wire n_1701;
wire n_318;
wire n_1111;
wire n_1713;
wire n_715;
wire n_1251;
wire n_1265;
wire n_1726;
wire n_1950;
wire n_530;
wire n_1563;
wire n_1912;
wire n_277;
wire n_1982;
wire n_618;
wire n_1297;
wire n_1662;
wire n_1312;
wire n_1167;
wire n_1359;
wire n_674;
wire n_871;
wire n_922;
wire n_268;
wire n_1335;
wire n_1760;
wire n_1927;
wire n_210;
wire n_2028;
wire n_1069;
wire n_1664;
wire n_1722;
wire n_612;
wire n_247;
wire n_1165;
wire n_355;
wire n_702;
wire n_347;
wire n_2008;
wire n_1926;
wire n_1175;
wire n_328;
wire n_1386;
wire n_1896;
wire n_429;
wire n_1747;
wire n_1012;
wire n_780;
wire n_675;
wire n_903;
wire n_1540;
wire n_1977;
wire n_1802;
wire n_1504;
wire n_286;
wire n_254;
wire n_1655;
wire n_242;
wire n_835;
wire n_928;
wire n_1214;
wire n_690;
wire n_850;
wire n_1801;
wire n_1886;
wire n_1654;
wire n_816;
wire n_1157;
wire n_1750;
wire n_1462;
wire n_1188;
wire n_1752;
wire n_877;
wire n_1813;
wire n_604;
wire n_825;
wire n_728;
wire n_1063;
wire n_1588;
wire n_267;
wire n_1124;
wire n_1624;
wire n_515;
wire n_1965;
wire n_598;
wire n_696;
wire n_1515;
wire n_961;
wire n_437;
wire n_1082;
wire n_1317;
wire n_593;
wire n_514;
wire n_687;
wire n_697;
wire n_890;
wire n_637;
wire n_295;
wire n_701;
wire n_950;
wire n_388;
wire n_484;
wire n_2036;
wire n_1709;
wire n_1825;
wire n_1796;
wire n_1757;
wire n_1792;
wire n_891;
wire n_1412;
wire n_949;
wire n_1630;
wire n_678;
wire n_283;
wire n_1987;
wire n_507;
wire n_968;
wire n_909;
wire n_1369;
wire n_881;
wire n_1008;
wire n_760;
wire n_1546;
wire n_590;
wire n_362;
wire n_462;
wire n_1033;
wire n_1052;
wire n_1296;
wire n_1990;
wire n_304;
wire n_694;
wire n_1294;
wire n_1420;
wire n_1634;
wire n_297;
wire n_595;
wire n_627;
wire n_1767;
wire n_1779;
wire n_524;
wire n_1465;
wire n_342;
wire n_1858;
wire n_1044;
wire n_1712;
wire n_1391;
wire n_449;
wire n_1523;
wire n_1208;
wire n_1164;
wire n_1295;
wire n_1627;
wire n_1072;
wire n_1527;
wire n_1495;
wire n_1438;
wire n_495;
wire n_815;
wire n_1100;
wire n_585;
wire n_1487;
wire n_840;
wire n_874;
wire n_1756;
wire n_1128;
wire n_673;
wire n_382;
wire n_1969;
wire n_1071;
wire n_1067;
wire n_1565;
wire n_1493;
wire n_1968;
wire n_898;
wire n_255;
wire n_284;
wire n_1952;
wire n_865;
wire n_925;
wire n_1932;
wire n_1101;
wire n_1026;
wire n_1880;
wire n_289;
wire n_1364;
wire n_615;
wire n_1249;
wire n_1293;
wire n_1127;
wire n_1512;
wire n_1451;
wire n_320;
wire n_639;
wire n_963;
wire n_794;
wire n_727;
wire n_894;
wire n_1839;
wire n_685;
wire n_1765;
wire n_353;
wire n_605;
wire n_1514;
wire n_1863;
wire n_826;
wire n_1646;
wire n_872;
wire n_1139;
wire n_1714;
wire n_718;
wire n_1018;
wire n_1521;
wire n_1366;
wire n_542;
wire n_847;
wire n_644;
wire n_682;
wire n_851;
wire n_305;
wire n_996;
wire n_532;
wire n_1308;
wire n_1376;
wire n_1513;
wire n_413;
wire n_791;
wire n_1913;
wire n_510;
wire n_837;
wire n_1488;
wire n_1808;
wire n_948;
wire n_704;
wire n_977;
wire n_1005;
wire n_1947;
wire n_536;
wire n_1788;
wire n_1999;
wire n_622;
wire n_1469;
wire n_1838;
wire n_1835;
wire n_1766;
wire n_1776;
wire n_1959;
wire n_2002;
wire n_581;
wire n_765;
wire n_432;
wire n_987;
wire n_1492;
wire n_1340;
wire n_1771;
wire n_631;
wire n_720;
wire n_842;
wire n_1707;
wire n_1432;
wire n_843;
wire n_656;
wire n_989;
wire n_1277;
wire n_797;
wire n_1473;
wire n_1723;
wire n_1246;
wire n_1878;
wire n_899;
wire n_738;
wire n_2012;
wire n_1304;
wire n_1035;
wire n_294;
wire n_499;
wire n_1426;
wire n_705;
wire n_1004;
wire n_1176;
wire n_1529;
wire n_1022;
wire n_614;
wire n_529;
wire n_425;
wire n_684;
wire n_1431;
wire n_1615;
wire n_1474;
wire n_1571;
wire n_1809;
wire n_1577;
wire n_1181;
wire n_1822;
wire n_486;
wire n_947;
wire n_1117;
wire n_1087;
wire n_1448;
wire n_1992;
wire n_648;
wire n_657;
wire n_1049;
wire n_1666;
wire n_1505;
wire n_803;
wire n_290;
wire n_1717;
wire n_926;
wire n_1817;
wire n_927;
wire n_1849;
wire n_919;
wire n_1698;
wire n_478;
wire n_929;
wire n_1228;
wire n_417;
wire n_446;
wire n_1568;
wire n_1490;
wire n_777;
wire n_1299;
wire n_272;
wire n_526;
wire n_1183;
wire n_1436;
wire n_1384;
wire n_293;
wire n_458;
wire n_1070;
wire n_998;
wire n_717;
wire n_1665;
wire n_1383;
wire n_1178;
wire n_1424;
wire n_1073;
wire n_1000;
wire n_796;
wire n_252;
wire n_1195;
wire n_1626;
wire n_1507;
wire n_552;
wire n_1358;
wire n_1811;
wire n_1388;
wire n_216;
wire n_912;
wire n_1857;
wire n_1519;
wire n_745;
wire n_1284;
wire n_1604;
wire n_1142;
wire n_716;
wire n_1475;
wire n_623;
wire n_1048;
wire n_1201;
wire n_1398;
wire n_884;
wire n_1774;
wire n_1395;
wire n_731;
wire n_1502;
wire n_1659;
wire n_1955;
wire n_755;
wire n_931;
wire n_1021;
wire n_527;
wire n_474;
wire n_683;
wire n_811;
wire n_1207;
wire n_312;
wire n_1791;
wire n_1368;
wire n_1418;
wire n_958;
wire n_292;
wire n_1250;
wire n_1137;
wire n_1897;
wire n_880;
wire n_889;
wire n_1478;
wire n_589;
wire n_1310;
wire n_819;
wire n_1363;
wire n_1334;
wire n_1942;
wire n_1966;
wire n_767;
wire n_1314;
wire n_600;
wire n_964;
wire n_831;
wire n_1837;
wire n_477;
wire n_954;
wire n_864;
wire n_1110;
wire n_1410;
wire n_399;
wire n_1440;
wire n_1382;
wire n_1534;
wire n_1564;
wire n_1736;
wire n_211;
wire n_1483;
wire n_1834;
wire n_1372;
wire n_231;
wire n_1457;
wire n_505;
wire n_1719;
wire n_319;
wire n_1339;
wire n_1787;
wire n_537;
wire n_1993;
wire n_1427;
wire n_311;
wire n_1466;
wire n_403;
wire n_1919;
wire n_1080;
wire n_723;
wire n_1877;
wire n_596;
wire n_546;
wire n_562;
wire n_1141;
wire n_1268;
wire n_386;
wire n_1939;
wire n_2030;
wire n_1769;
wire n_1220;
wire n_1893;
wire n_556;
wire n_1755;
wire n_1602;
wire n_1136;
wire n_2025;
wire n_1125;
wire n_970;
wire n_1980;
wire n_642;
wire n_995;
wire n_276;
wire n_1159;
wire n_1092;
wire n_441;
wire n_221;
wire n_1060;
wire n_1951;
wire n_444;
wire n_1252;
wire n_1784;
wire n_1223;
wire n_303;
wire n_511;
wire n_1286;
wire n_1773;
wire n_1775;
wire n_1053;
wire n_416;
wire n_1681;
wire n_520;
wire n_418;
wire n_1093;
wire n_1783;
wire n_1533;
wire n_1597;
wire n_266;
wire n_296;
wire n_775;
wire n_651;
wire n_1153;
wire n_439;
wire n_1618;
wire n_217;
wire n_518;
wire n_1531;
wire n_1185;
wire n_453;
wire n_215;
wire n_1745;
wire n_914;
wire n_759;
wire n_1831;
wire n_426;
wire n_317;
wire n_1653;
wire n_1679;
wire n_1625;
wire n_1453;
wire n_488;
wire n_497;
wire n_773;
wire n_1901;
wire n_920;
wire n_1374;
wire n_1315;
wire n_1647;
wire n_1224;
wire n_1614;
wire n_1459;
wire n_1892;
wire n_1933;
wire n_1135;
wire n_1169;
wire n_1179;
wire n_401;
wire n_324;
wire n_1617;
wire n_335;
wire n_1470;
wire n_463;
wire n_1243;
wire n_848;
wire n_301;
wire n_274;
wire n_1096;
wire n_1091;
wire n_1917;
wire n_2000;
wire n_1580;
wire n_1425;
wire n_1881;
wire n_1267;
wire n_1281;
wire n_1806;
wire n_983;
wire n_2023;
wire n_427;
wire n_1520;
wire n_496;
wire n_906;
wire n_1390;
wire n_688;
wire n_1077;
wire n_1733;
wire n_1419;
wire n_351;
wire n_259;
wire n_1731;
wire n_1855;
wire n_1636;
wire n_1437;
wire n_1645;
wire n_1832;
wire n_385;
wire n_1687;
wire n_1439;
wire n_1323;
wire n_858;
wire n_1331;
wire n_613;
wire n_736;
wire n_501;
wire n_956;
wire n_960;
wire n_663;
wire n_856;
wire n_379;
wire n_778;
wire n_1668;
wire n_1134;
wire n_410;
wire n_1129;
wire n_554;
wire n_602;
wire n_1696;
wire n_1995;
wire n_1594;
wire n_664;
wire n_1869;
wire n_1764;
wire n_1429;
wire n_1610;
wire n_1889;
wire n_435;
wire n_1905;
wire n_2016;
wire n_793;
wire n_326;
wire n_587;
wire n_1593;
wire n_580;
wire n_762;
wire n_1030;
wire n_1202;
wire n_1937;
wire n_465;
wire n_1790;
wire n_1778;
wire n_1635;
wire n_1079;
wire n_341;
wire n_1744;
wire n_828;
wire n_607;
wire n_316;
wire n_419;
wire n_1551;
wire n_1103;
wire n_1203;
wire n_820;
wire n_951;
wire n_725;
wire n_952;
wire n_999;
wire n_358;
wire n_1254;
wire n_368;
wire n_575;
wire n_994;
wire n_1508;
wire n_732;
wire n_974;
wire n_392;
wire n_724;
wire n_1934;
wire n_1020;
wire n_1042;
wire n_628;
wire n_1273;
wire n_1434;
wire n_1573;
wire n_1728;
wire n_557;
wire n_1871;
wire n_349;
wire n_617;
wire n_845;
wire n_807;
wire n_1036;
wire n_1138;
wire n_1661;
wire n_1275;
wire n_485;
wire n_1549;
wire n_443;
wire n_1510;
wire n_892;
wire n_768;
wire n_421;
wire n_1468;
wire n_1859;
wire n_238;
wire n_1095;
wire n_2024;
wire n_1595;
wire n_1718;
wire n_1749;
wire n_1683;
wire n_1916;
wire n_597;
wire n_280;
wire n_1270;
wire n_1187;
wire n_610;
wire n_1403;
wire n_1669;
wire n_1852;
wire n_1024;
wire n_1768;
wire n_1847;
wire n_248;
wire n_517;
wire n_1667;
wire n_667;
wire n_1206;
wire n_621;
wire n_1037;
wire n_1397;
wire n_1279;
wire n_1115;
wire n_750;
wire n_901;
wire n_1499;
wire n_468;
wire n_923;
wire n_504;
wire n_1409;
wire n_1841;
wire n_1639;
wire n_1623;
wire n_1015;
wire n_1503;
wire n_466;
wire n_1057;
wire n_603;
wire n_991;
wire n_1657;
wire n_235;
wire n_1126;
wire n_1997;
wire n_340;
wire n_710;
wire n_1108;
wire n_1818;
wire n_1182;
wire n_1298;
wire n_1611;
wire n_785;
wire n_746;
wire n_609;
wire n_1601;
wire n_1960;
wire n_1686;
wire n_1356;
wire n_1589;
wire n_1740;
wire n_1497;
wire n_1168;
wire n_1216;
wire n_1943;
wire n_1320;
wire n_1430;
wire n_1316;
wire n_1287;
wire n_1452;
wire n_1622;
wire n_1586;
wire n_302;
wire n_1694;
wire n_380;
wire n_1535;
wire n_1596;
wire n_1190;
wire n_1734;
wire n_397;
wire n_1983;
wire n_1938;
wire n_1262;
wire n_218;
wire n_1891;
wire n_1213;
wire n_1350;
wire n_1673;
wire n_1715;
wire n_1443;
wire n_1272;
wire n_239;
wire n_2037;
wire n_782;
wire n_1539;
wire n_490;
wire n_220;
wire n_809;
wire n_1043;
wire n_1797;
wire n_1608;
wire n_986;
wire n_1472;
wire n_1081;
wire n_402;
wire n_1870;
wire n_352;
wire n_1692;
wire n_800;
wire n_1084;
wire n_1171;
wire n_460;
wire n_1827;
wire n_1361;
wire n_1864;
wire n_2006;
wire n_1491;
wire n_662;
wire n_374;
wire n_1152;
wire n_1840;
wire n_1705;
wire n_450;
wire n_1684;
wire n_921;
wire n_1346;
wire n_711;
wire n_1642;
wire n_579;
wire n_1352;
wire n_937;
wire n_1682;
wire n_2017;
wire n_370;
wire n_1695;
wire n_1828;
wire n_650;
wire n_1046;
wire n_1940;
wire n_1979;
wire n_1145;
wire n_330;
wire n_1121;
wire n_1102;
wire n_1963;
wire n_972;
wire n_1405;
wire n_258;
wire n_1406;
wire n_456;
wire n_1332;
wire n_260;
wire n_313;
wire n_624;
wire n_962;
wire n_1041;
wire n_565;
wire n_356;
wire n_1569;
wire n_936;
wire n_1883;
wire n_1288;
wire n_1186;
wire n_1062;
wire n_885;
wire n_896;
wire n_654;
wire n_411;
wire n_1222;
wire n_599;
wire n_776;
wire n_321;
wire n_1823;
wire n_227;
wire n_1974;
wire n_1720;
wire n_482;
wire n_934;
wire n_1637;
wire n_1407;
wire n_1795;
wire n_420;
wire n_1341;
wire n_394;
wire n_1456;
wire n_1845;
wire n_1489;
wire n_942;
wire n_1524;
wire n_543;
wire n_1964;
wire n_1920;
wire n_1496;
wire n_1271;
wire n_1545;
wire n_2007;
wire n_1946;
wire n_1355;
wire n_1225;
wire n_1544;
wire n_1485;
wire n_325;
wire n_1640;
wire n_804;
wire n_464;
wire n_1846;
wire n_533;
wire n_806;
wire n_879;
wire n_959;
wire n_584;
wire n_244;
wire n_1343;
wire n_1522;
wire n_548;
wire n_1782;
wire n_282;
wire n_1676;
wire n_833;
wire n_1830;
wire n_1567;
wire n_523;
wire n_1319;
wire n_707;
wire n_345;
wire n_1900;
wire n_799;
wire n_1548;
wire n_1155;
wire n_273;
wire n_1633;
wire n_787;
wire n_1416;
wire n_1528;
wire n_1146;
wire n_2021;
wire n_1086;
wire n_1066;
wire n_1948;
wire n_2026;
wire n_1282;
wire n_550;
wire n_275;
wire n_652;
wire n_560;
wire n_1906;
wire n_1484;
wire n_1241;
wire n_1321;
wire n_1672;
wire n_569;
wire n_1758;
wire n_1925;
wire n_737;
wire n_1318;
wire n_1914;
wire n_1235;
wire n_1229;
wire n_306;
wire n_1292;
wire n_1373;
wire n_346;
wire n_1029;
wire n_1447;
wire n_790;
wire n_1706;
wire n_1498;
wire n_1210;
wire n_299;
wire n_1248;
wire n_1556;
wire n_902;
wire n_333;
wire n_1047;
wire n_1984;
wire n_1385;
wire n_431;
wire n_459;
wire n_1269;
wire n_1931;
wire n_502;
wire n_672;
wire n_1257;
wire n_1751;
wire n_285;
wire n_1375;
wire n_1941;
wire n_655;
wire n_706;
wire n_1045;
wire n_1650;
wire n_786;
wire n_1794;
wire n_1236;
wire n_1962;
wire n_1559;
wire n_1725;
wire n_1928;
wire n_1872;
wire n_834;
wire n_743;
wire n_766;
wire n_430;
wire n_1746;
wire n_1325;
wire n_1002;
wire n_1741;
wire n_1949;
wire n_545;
wire n_489;
wire n_1804;
wire n_1727;
wire n_251;
wire n_1019;
wire n_636;
wire n_729;
wire n_876;
wire n_774;
wire n_1337;
wire n_660;
wire n_438;
wire n_1477;
wire n_1360;
wire n_1860;
wire n_1904;
wire n_1200;
wire n_479;
wire n_1607;
wire n_1353;
wire n_1777;
wire n_1908;
wire n_1454;
wire n_869;
wire n_1154;
wire n_1113;
wire n_1600;
wire n_646;
wire n_528;
wire n_391;
wire n_1098;
wire n_1329;
wire n_817;
wire n_262;
wire n_897;
wire n_846;
wire n_841;
wire n_1476;
wire n_1001;
wire n_508;
wire n_1800;
wire n_1050;
wire n_1411;
wire n_1463;
wire n_1177;
wire n_332;
wire n_1150;
wire n_1742;
wire n_1562;
wire n_1690;
wire n_398;
wire n_1191;
wire n_1826;
wire n_566;
wire n_1023;
wire n_1882;
wire n_1076;
wire n_1118;
wire n_1007;
wire n_1807;
wire n_1929;
wire n_1378;
wire n_855;
wire n_1592;
wire n_1759;
wire n_1814;
wire n_1631;
wire n_591;
wire n_1377;
wire n_1879;
wire n_256;
wire n_853;
wire n_440;
wire n_695;
wire n_1542;
wire n_875;
wire n_209;
wire n_367;
wire n_680;
wire n_1678;
wire n_661;
wire n_1716;
wire n_278;
wire n_1256;
wire n_671;
wire n_1953;
wire n_933;
wire n_740;
wire n_703;
wire n_978;
wire n_384;
wire n_1976;
wire n_1291;
wire n_1217;
wire n_751;
wire n_749;
wire n_1824;
wire n_310;
wire n_1628;
wire n_1324;
wire n_1399;
wire n_1435;
wire n_969;
wire n_988;
wire n_1065;
wire n_1401;
wire n_1255;
wire n_568;
wire n_1516;
wire n_1536;
wire n_2029;
wire n_1204;
wire n_823;
wire n_1132;
wire n_643;
wire n_233;
wire n_698;
wire n_1074;
wire n_1394;
wire n_1327;
wire n_1326;
wire n_739;
wire n_400;
wire n_955;
wire n_337;
wire n_1379;
wire n_214;
wire n_246;
wire n_1338;
wire n_1097;
wire n_935;
wire n_781;
wire n_789;
wire n_1554;
wire n_1130;
wire n_1810;
wire n_573;
wire n_769;
wire n_676;
wire n_327;
wire n_1120;
wire n_832;
wire n_1583;
wire n_1730;
wire n_555;
wire n_389;
wire n_814;
wire n_1643;
wire n_2020;
wire n_1729;
wire n_669;
wire n_300;
wire n_222;
wire n_2005;
wire n_747;
wire n_1389;
wire n_1105;
wire n_721;
wire n_1461;
wire n_742;
wire n_535;
wire n_691;
wire n_372;
wire n_314;
wire n_1408;
wire n_378;
wire n_1196;
wire n_377;
wire n_1598;
wire n_863;
wire n_601;
wire n_338;
wire n_1283;
wire n_918;
wire n_748;
wire n_506;
wire n_1114;
wire n_1785;
wire n_763;
wire n_1147;
wire n_1848;
wire n_360;
wire n_1754;
wire n_1506;
wire n_1652;
wire n_1812;
wire n_957;
wire n_1994;
wire n_895;
wire n_866;
wire n_1227;
wire n_387;
wire n_452;
wire n_744;
wire n_971;
wire n_946;
wire n_344;
wire n_761;
wire n_1303;
wire n_1205;
wire n_1258;
wire n_1392;
wire n_1173;
wire n_1924;
wire n_525;
wire n_1677;
wire n_1116;
wire n_611;
wire n_1570;
wire n_1702;
wire n_1219;
wire n_1780;
wire n_1689;
wire n_1174;
wire n_1944;
wire n_1016;
wire n_1347;
wire n_795;
wire n_1501;
wire n_1221;
wire n_1245;
wire n_838;
wire n_647;
wire n_844;
wire n_448;
wire n_1017;
wire n_1083;
wire n_445;
wire n_1561;
wire n_930;
wire n_888;
wire n_1112;
wire n_234;
wire n_2022;
wire n_1945;
wire n_910;
wire n_1656;
wire n_1721;
wire n_1460;
wire n_911;
wire n_1464;
wire n_653;
wire n_236;
wire n_1737;
wire n_1414;
wire n_752;
wire n_908;
wire n_944;
wire n_2034;
wire n_576;
wire n_1028;
wire n_472;
wire n_270;
wire n_414;
wire n_1922;
wire n_563;
wire n_2032;
wire n_1011;
wire n_1566;
wire n_1215;
wire n_839;
wire n_708;
wire n_1973;
wire n_668;
wire n_626;
wire n_990;
wire n_1500;
wire n_779;
wire n_1537;
wire n_1821;
wire n_1104;
wire n_854;
wire n_1058;
wire n_498;
wire n_1122;
wire n_870;
wire n_904;
wire n_1253;
wire n_709;
wire n_1266;
wire n_366;
wire n_1509;
wire n_1693;
wire n_1109;
wire n_712;
wire n_348;
wire n_1276;
wire n_376;
wire n_2015;
wire n_390;
wire n_1148;
wire n_334;
wire n_1989;
wire n_1161;
wire n_1085;
wire n_232;
wire n_2014;
wire n_1239;
wire n_771;
wire n_1584;
wire n_470;
wire n_475;
wire n_924;
wire n_298;
wire n_1582;
wire n_492;
wire n_1149;
wire n_265;
wire n_1184;
wire n_228;
wire n_719;
wire n_1972;
wire n_1525;
wire n_455;
wire n_1585;
wire n_1851;
wire n_363;
wire n_1799;
wire n_1090;
wire n_592;
wire n_1816;
wire n_1518;
wire n_829;
wire n_1156;
wire n_1362;
wire n_393;
wire n_984;
wire n_1829;
wire n_503;
wire n_2035;
wire n_1450;
wire n_1638;
wire n_868;
wire n_570;
wire n_859;
wire n_2033;
wire n_406;
wire n_735;
wire n_1789;
wire n_1770;
wire n_878;
wire n_620;
wire n_519;
wire n_307;
wire n_469;
wire n_1218;
wire n_500;
wire n_1482;
wire n_981;
wire n_714;
wire n_1349;
wire n_291;
wire n_1144;
wire n_357;
wire n_985;
wire n_481;
wire n_997;
wire n_1710;
wire n_1301;
wire n_802;
wire n_561;
wire n_980;
wire n_1306;
wire n_2010;
wire n_1651;
wire n_1198;
wire n_1609;
wire n_436;
wire n_409;
wire n_1244;
wire n_1685;
wire n_1763;
wire n_1998;
wire n_1574;
wire n_240;
wire n_756;
wire n_1619;
wire n_1981;
wire n_1606;
wire n_810;
wire n_1133;
wire n_635;
wire n_1194;
wire n_1051;
wire n_253;
wire n_1552;
wire n_583;
wire n_1996;
wire n_249;
wire n_1039;
wire n_1442;
wire n_1034;
wire n_1480;
wire n_1158;
wire n_754;
wire n_941;
wire n_975;
wire n_1031;
wire n_1305;
wire n_553;
wire n_849;
wire n_753;
wire n_1753;
wire n_467;
wire n_269;
wire n_359;
wire n_973;
wire n_1921;
wire n_1479;
wire n_1055;
wire n_1675;
wire n_582;
wire n_861;
wire n_857;
wire n_967;
wire n_571;
wire n_271;
wire n_404;
wire n_2001;
wire n_1884;
wire n_679;
wire n_633;
wire n_1170;
wire n_665;
wire n_1629;
wire n_588;
wire n_225;
wire n_1260;
wire n_308;
wire n_309;
wire n_1819;
wire n_1010;
wire n_1040;
wire n_915;
wire n_632;
wire n_1166;
wire n_2038;
wire n_812;
wire n_1131;
wire n_1761;
wire n_534;
wire n_1578;
wire n_1006;
wire n_1861;
wire n_373;
wire n_1632;
wire n_1890;
wire n_1805;
wire n_257;
wire n_1557;
wire n_1888;
wire n_1833;
wire n_730;
wire n_1311;
wire n_1494;
wire n_670;
wire n_1850;
wire n_1898;
wire n_1868;
wire n_1089;
wire n_1887;
wire n_1587;
wire n_1365;
wire n_1417;
wire n_1242;
wire n_1836;
wire n_681;
wire n_1226;
wire n_1274;
wire n_1486;
wire n_412;
wire n_640;
wire n_1322;
wire n_965;
wire n_1899;
wire n_1428;
wire n_1616;
wire n_1576;
wire n_1862;
wire n_1856;
wire n_1958;
wire n_339;
wire n_784;
wire n_434;
wire n_315;
wire n_288;
wire n_1059;
wire n_1197;
wire n_422;
wire n_722;
wire n_862;
wire n_540;
wire n_1423;
wire n_1935;
wire n_2027;
wire n_457;
wire n_364;
wire n_1915;
wire n_629;
wire n_1621;
wire n_1748;
wire n_900;
wire n_1449;
wire n_531;
wire n_827;
wire n_361;
wire n_1025;
wire n_336;
wire n_1885;
wire n_1013;
wire n_1259;
wire n_1538;
wire n_649;
wire n_1612;
wire n_1240;

CKINVDCx20_ASAP7_75t_R g209 ( 
.A(n_144),
.Y(n_209)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_155),
.Y(n_210)
);

BUFx6f_ASAP7_75t_L g211 ( 
.A(n_93),
.Y(n_211)
);

INVx1_ASAP7_75t_SL g212 ( 
.A(n_85),
.Y(n_212)
);

INVx2_ASAP7_75t_L g213 ( 
.A(n_171),
.Y(n_213)
);

CKINVDCx5p33_ASAP7_75t_R g214 ( 
.A(n_195),
.Y(n_214)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_60),
.Y(n_215)
);

CKINVDCx5p33_ASAP7_75t_R g216 ( 
.A(n_161),
.Y(n_216)
);

CKINVDCx5p33_ASAP7_75t_R g217 ( 
.A(n_2),
.Y(n_217)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_122),
.Y(n_218)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_110),
.Y(n_219)
);

CKINVDCx5p33_ASAP7_75t_R g220 ( 
.A(n_64),
.Y(n_220)
);

CKINVDCx5p33_ASAP7_75t_R g221 ( 
.A(n_174),
.Y(n_221)
);

BUFx2_ASAP7_75t_L g222 ( 
.A(n_125),
.Y(n_222)
);

CKINVDCx5p33_ASAP7_75t_R g223 ( 
.A(n_37),
.Y(n_223)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_118),
.Y(n_224)
);

CKINVDCx20_ASAP7_75t_R g225 ( 
.A(n_90),
.Y(n_225)
);

CKINVDCx5p33_ASAP7_75t_R g226 ( 
.A(n_136),
.Y(n_226)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_192),
.Y(n_227)
);

CKINVDCx20_ASAP7_75t_R g228 ( 
.A(n_121),
.Y(n_228)
);

CKINVDCx20_ASAP7_75t_R g229 ( 
.A(n_162),
.Y(n_229)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_166),
.Y(n_230)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_164),
.Y(n_231)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_176),
.Y(n_232)
);

CKINVDCx5p33_ASAP7_75t_R g233 ( 
.A(n_32),
.Y(n_233)
);

HB1xp67_ASAP7_75t_L g234 ( 
.A(n_18),
.Y(n_234)
);

INVx1_ASAP7_75t_SL g235 ( 
.A(n_135),
.Y(n_235)
);

CKINVDCx5p33_ASAP7_75t_R g236 ( 
.A(n_177),
.Y(n_236)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_37),
.Y(n_237)
);

CKINVDCx5p33_ASAP7_75t_R g238 ( 
.A(n_191),
.Y(n_238)
);

CKINVDCx5p33_ASAP7_75t_R g239 ( 
.A(n_69),
.Y(n_239)
);

CKINVDCx5p33_ASAP7_75t_R g240 ( 
.A(n_36),
.Y(n_240)
);

CKINVDCx5p33_ASAP7_75t_R g241 ( 
.A(n_63),
.Y(n_241)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_103),
.Y(n_242)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_25),
.Y(n_243)
);

CKINVDCx5p33_ASAP7_75t_R g244 ( 
.A(n_205),
.Y(n_244)
);

CKINVDCx5p33_ASAP7_75t_R g245 ( 
.A(n_147),
.Y(n_245)
);

CKINVDCx5p33_ASAP7_75t_R g246 ( 
.A(n_87),
.Y(n_246)
);

CKINVDCx5p33_ASAP7_75t_R g247 ( 
.A(n_9),
.Y(n_247)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_82),
.Y(n_248)
);

CKINVDCx5p33_ASAP7_75t_R g249 ( 
.A(n_17),
.Y(n_249)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_20),
.Y(n_250)
);

CKINVDCx5p33_ASAP7_75t_R g251 ( 
.A(n_95),
.Y(n_251)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_46),
.Y(n_252)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_178),
.Y(n_253)
);

CKINVDCx5p33_ASAP7_75t_R g254 ( 
.A(n_30),
.Y(n_254)
);

CKINVDCx5p33_ASAP7_75t_R g255 ( 
.A(n_153),
.Y(n_255)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_156),
.Y(n_256)
);

INVx2_ASAP7_75t_SL g257 ( 
.A(n_45),
.Y(n_257)
);

CKINVDCx5p33_ASAP7_75t_R g258 ( 
.A(n_165),
.Y(n_258)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_113),
.Y(n_259)
);

CKINVDCx5p33_ASAP7_75t_R g260 ( 
.A(n_132),
.Y(n_260)
);

CKINVDCx5p33_ASAP7_75t_R g261 ( 
.A(n_49),
.Y(n_261)
);

CKINVDCx5p33_ASAP7_75t_R g262 ( 
.A(n_199),
.Y(n_262)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_111),
.Y(n_263)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_127),
.Y(n_264)
);

CKINVDCx5p33_ASAP7_75t_R g265 ( 
.A(n_1),
.Y(n_265)
);

CKINVDCx5p33_ASAP7_75t_R g266 ( 
.A(n_148),
.Y(n_266)
);

CKINVDCx5p33_ASAP7_75t_R g267 ( 
.A(n_32),
.Y(n_267)
);

CKINVDCx20_ASAP7_75t_R g268 ( 
.A(n_193),
.Y(n_268)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_52),
.Y(n_269)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_65),
.Y(n_270)
);

CKINVDCx5p33_ASAP7_75t_R g271 ( 
.A(n_124),
.Y(n_271)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_170),
.Y(n_272)
);

CKINVDCx5p33_ASAP7_75t_R g273 ( 
.A(n_99),
.Y(n_273)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_38),
.Y(n_274)
);

CKINVDCx5p33_ASAP7_75t_R g275 ( 
.A(n_183),
.Y(n_275)
);

INVx1_ASAP7_75t_SL g276 ( 
.A(n_68),
.Y(n_276)
);

CKINVDCx5p33_ASAP7_75t_R g277 ( 
.A(n_123),
.Y(n_277)
);

CKINVDCx5p33_ASAP7_75t_R g278 ( 
.A(n_31),
.Y(n_278)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_190),
.Y(n_279)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_60),
.Y(n_280)
);

INVx1_ASAP7_75t_SL g281 ( 
.A(n_35),
.Y(n_281)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_181),
.Y(n_282)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_62),
.Y(n_283)
);

CKINVDCx20_ASAP7_75t_R g284 ( 
.A(n_128),
.Y(n_284)
);

CKINVDCx5p33_ASAP7_75t_R g285 ( 
.A(n_185),
.Y(n_285)
);

CKINVDCx20_ASAP7_75t_R g286 ( 
.A(n_204),
.Y(n_286)
);

CKINVDCx5p33_ASAP7_75t_R g287 ( 
.A(n_12),
.Y(n_287)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_13),
.Y(n_288)
);

BUFx2_ASAP7_75t_L g289 ( 
.A(n_34),
.Y(n_289)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_142),
.Y(n_290)
);

BUFx10_ASAP7_75t_L g291 ( 
.A(n_96),
.Y(n_291)
);

BUFx10_ASAP7_75t_L g292 ( 
.A(n_198),
.Y(n_292)
);

CKINVDCx5p33_ASAP7_75t_R g293 ( 
.A(n_158),
.Y(n_293)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_149),
.Y(n_294)
);

CKINVDCx5p33_ASAP7_75t_R g295 ( 
.A(n_68),
.Y(n_295)
);

INVx1_ASAP7_75t_SL g296 ( 
.A(n_88),
.Y(n_296)
);

BUFx3_ASAP7_75t_L g297 ( 
.A(n_43),
.Y(n_297)
);

CKINVDCx5p33_ASAP7_75t_R g298 ( 
.A(n_10),
.Y(n_298)
);

CKINVDCx5p33_ASAP7_75t_R g299 ( 
.A(n_151),
.Y(n_299)
);

CKINVDCx5p33_ASAP7_75t_R g300 ( 
.A(n_27),
.Y(n_300)
);

CKINVDCx5p33_ASAP7_75t_R g301 ( 
.A(n_196),
.Y(n_301)
);

CKINVDCx5p33_ASAP7_75t_R g302 ( 
.A(n_168),
.Y(n_302)
);

BUFx6f_ASAP7_75t_L g303 ( 
.A(n_6),
.Y(n_303)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_42),
.Y(n_304)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_72),
.Y(n_305)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_30),
.Y(n_306)
);

INVx2_ASAP7_75t_L g307 ( 
.A(n_65),
.Y(n_307)
);

INVx2_ASAP7_75t_L g308 ( 
.A(n_10),
.Y(n_308)
);

CKINVDCx20_ASAP7_75t_R g309 ( 
.A(n_38),
.Y(n_309)
);

CKINVDCx5p33_ASAP7_75t_R g310 ( 
.A(n_73),
.Y(n_310)
);

BUFx3_ASAP7_75t_L g311 ( 
.A(n_115),
.Y(n_311)
);

CKINVDCx5p33_ASAP7_75t_R g312 ( 
.A(n_152),
.Y(n_312)
);

CKINVDCx5p33_ASAP7_75t_R g313 ( 
.A(n_3),
.Y(n_313)
);

CKINVDCx5p33_ASAP7_75t_R g314 ( 
.A(n_77),
.Y(n_314)
);

INVx2_ASAP7_75t_L g315 ( 
.A(n_58),
.Y(n_315)
);

CKINVDCx5p33_ASAP7_75t_R g316 ( 
.A(n_89),
.Y(n_316)
);

CKINVDCx5p33_ASAP7_75t_R g317 ( 
.A(n_131),
.Y(n_317)
);

CKINVDCx14_ASAP7_75t_R g318 ( 
.A(n_25),
.Y(n_318)
);

BUFx3_ASAP7_75t_L g319 ( 
.A(n_117),
.Y(n_319)
);

CKINVDCx5p33_ASAP7_75t_R g320 ( 
.A(n_104),
.Y(n_320)
);

CKINVDCx5p33_ASAP7_75t_R g321 ( 
.A(n_1),
.Y(n_321)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_100),
.Y(n_322)
);

CKINVDCx5p33_ASAP7_75t_R g323 ( 
.A(n_180),
.Y(n_323)
);

CKINVDCx20_ASAP7_75t_R g324 ( 
.A(n_173),
.Y(n_324)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_36),
.Y(n_325)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_167),
.Y(n_326)
);

CKINVDCx5p33_ASAP7_75t_R g327 ( 
.A(n_78),
.Y(n_327)
);

CKINVDCx5p33_ASAP7_75t_R g328 ( 
.A(n_50),
.Y(n_328)
);

CKINVDCx16_ASAP7_75t_R g329 ( 
.A(n_163),
.Y(n_329)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_53),
.Y(n_330)
);

CKINVDCx5p33_ASAP7_75t_R g331 ( 
.A(n_57),
.Y(n_331)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_39),
.Y(n_332)
);

CKINVDCx5p33_ASAP7_75t_R g333 ( 
.A(n_140),
.Y(n_333)
);

CKINVDCx5p33_ASAP7_75t_R g334 ( 
.A(n_17),
.Y(n_334)
);

CKINVDCx5p33_ASAP7_75t_R g335 ( 
.A(n_75),
.Y(n_335)
);

CKINVDCx20_ASAP7_75t_R g336 ( 
.A(n_45),
.Y(n_336)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_52),
.Y(n_337)
);

INVx1_ASAP7_75t_L g338 ( 
.A(n_3),
.Y(n_338)
);

CKINVDCx5p33_ASAP7_75t_R g339 ( 
.A(n_33),
.Y(n_339)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_58),
.Y(n_340)
);

INVxp67_ASAP7_75t_L g341 ( 
.A(n_105),
.Y(n_341)
);

CKINVDCx5p33_ASAP7_75t_R g342 ( 
.A(n_130),
.Y(n_342)
);

CKINVDCx5p33_ASAP7_75t_R g343 ( 
.A(n_202),
.Y(n_343)
);

BUFx10_ASAP7_75t_L g344 ( 
.A(n_143),
.Y(n_344)
);

CKINVDCx5p33_ASAP7_75t_R g345 ( 
.A(n_79),
.Y(n_345)
);

CKINVDCx5p33_ASAP7_75t_R g346 ( 
.A(n_35),
.Y(n_346)
);

INVx1_ASAP7_75t_L g347 ( 
.A(n_108),
.Y(n_347)
);

CKINVDCx5p33_ASAP7_75t_R g348 ( 
.A(n_8),
.Y(n_348)
);

INVx1_ASAP7_75t_SL g349 ( 
.A(n_137),
.Y(n_349)
);

INVx1_ASAP7_75t_SL g350 ( 
.A(n_201),
.Y(n_350)
);

INVx1_ASAP7_75t_L g351 ( 
.A(n_24),
.Y(n_351)
);

INVx1_ASAP7_75t_L g352 ( 
.A(n_7),
.Y(n_352)
);

INVxp67_ASAP7_75t_SL g353 ( 
.A(n_169),
.Y(n_353)
);

CKINVDCx5p33_ASAP7_75t_R g354 ( 
.A(n_146),
.Y(n_354)
);

CKINVDCx5p33_ASAP7_75t_R g355 ( 
.A(n_187),
.Y(n_355)
);

CKINVDCx5p33_ASAP7_75t_R g356 ( 
.A(n_67),
.Y(n_356)
);

INVx1_ASAP7_75t_L g357 ( 
.A(n_9),
.Y(n_357)
);

INVx1_ASAP7_75t_L g358 ( 
.A(n_24),
.Y(n_358)
);

INVx1_ASAP7_75t_L g359 ( 
.A(n_81),
.Y(n_359)
);

CKINVDCx5p33_ASAP7_75t_R g360 ( 
.A(n_139),
.Y(n_360)
);

INVx1_ASAP7_75t_L g361 ( 
.A(n_94),
.Y(n_361)
);

CKINVDCx5p33_ASAP7_75t_R g362 ( 
.A(n_112),
.Y(n_362)
);

CKINVDCx5p33_ASAP7_75t_R g363 ( 
.A(n_84),
.Y(n_363)
);

INVx1_ASAP7_75t_SL g364 ( 
.A(n_29),
.Y(n_364)
);

INVx1_ASAP7_75t_SL g365 ( 
.A(n_80),
.Y(n_365)
);

HB1xp67_ASAP7_75t_L g366 ( 
.A(n_59),
.Y(n_366)
);

CKINVDCx5p33_ASAP7_75t_R g367 ( 
.A(n_189),
.Y(n_367)
);

BUFx3_ASAP7_75t_L g368 ( 
.A(n_114),
.Y(n_368)
);

INVx1_ASAP7_75t_L g369 ( 
.A(n_70),
.Y(n_369)
);

INVx1_ASAP7_75t_SL g370 ( 
.A(n_83),
.Y(n_370)
);

INVx1_ASAP7_75t_L g371 ( 
.A(n_48),
.Y(n_371)
);

BUFx5_ASAP7_75t_L g372 ( 
.A(n_11),
.Y(n_372)
);

CKINVDCx5p33_ASAP7_75t_R g373 ( 
.A(n_119),
.Y(n_373)
);

CKINVDCx5p33_ASAP7_75t_R g374 ( 
.A(n_39),
.Y(n_374)
);

INVx1_ASAP7_75t_L g375 ( 
.A(n_34),
.Y(n_375)
);

INVx1_ASAP7_75t_L g376 ( 
.A(n_150),
.Y(n_376)
);

INVx1_ASAP7_75t_L g377 ( 
.A(n_109),
.Y(n_377)
);

CKINVDCx5p33_ASAP7_75t_R g378 ( 
.A(n_120),
.Y(n_378)
);

INVxp67_ASAP7_75t_L g379 ( 
.A(n_67),
.Y(n_379)
);

BUFx10_ASAP7_75t_L g380 ( 
.A(n_76),
.Y(n_380)
);

CKINVDCx5p33_ASAP7_75t_R g381 ( 
.A(n_42),
.Y(n_381)
);

CKINVDCx5p33_ASAP7_75t_R g382 ( 
.A(n_47),
.Y(n_382)
);

INVx1_ASAP7_75t_L g383 ( 
.A(n_179),
.Y(n_383)
);

CKINVDCx16_ASAP7_75t_R g384 ( 
.A(n_54),
.Y(n_384)
);

CKINVDCx5p33_ASAP7_75t_R g385 ( 
.A(n_203),
.Y(n_385)
);

CKINVDCx20_ASAP7_75t_R g386 ( 
.A(n_7),
.Y(n_386)
);

CKINVDCx5p33_ASAP7_75t_R g387 ( 
.A(n_126),
.Y(n_387)
);

INVx1_ASAP7_75t_L g388 ( 
.A(n_14),
.Y(n_388)
);

CKINVDCx5p33_ASAP7_75t_R g389 ( 
.A(n_141),
.Y(n_389)
);

INVx1_ASAP7_75t_L g390 ( 
.A(n_194),
.Y(n_390)
);

INVx1_ASAP7_75t_L g391 ( 
.A(n_207),
.Y(n_391)
);

CKINVDCx5p33_ASAP7_75t_R g392 ( 
.A(n_102),
.Y(n_392)
);

INVx1_ASAP7_75t_L g393 ( 
.A(n_4),
.Y(n_393)
);

CKINVDCx5p33_ASAP7_75t_R g394 ( 
.A(n_86),
.Y(n_394)
);

CKINVDCx16_ASAP7_75t_R g395 ( 
.A(n_188),
.Y(n_395)
);

INVx1_ASAP7_75t_L g396 ( 
.A(n_106),
.Y(n_396)
);

INVx1_ASAP7_75t_L g397 ( 
.A(n_27),
.Y(n_397)
);

CKINVDCx5p33_ASAP7_75t_R g398 ( 
.A(n_71),
.Y(n_398)
);

BUFx10_ASAP7_75t_L g399 ( 
.A(n_107),
.Y(n_399)
);

CKINVDCx5p33_ASAP7_75t_R g400 ( 
.A(n_21),
.Y(n_400)
);

CKINVDCx5p33_ASAP7_75t_R g401 ( 
.A(n_44),
.Y(n_401)
);

CKINVDCx5p33_ASAP7_75t_R g402 ( 
.A(n_63),
.Y(n_402)
);

INVxp67_ASAP7_75t_L g403 ( 
.A(n_26),
.Y(n_403)
);

INVx1_ASAP7_75t_L g404 ( 
.A(n_15),
.Y(n_404)
);

INVx1_ASAP7_75t_L g405 ( 
.A(n_56),
.Y(n_405)
);

CKINVDCx5p33_ASAP7_75t_R g406 ( 
.A(n_47),
.Y(n_406)
);

BUFx3_ASAP7_75t_L g407 ( 
.A(n_59),
.Y(n_407)
);

INVx1_ASAP7_75t_L g408 ( 
.A(n_172),
.Y(n_408)
);

CKINVDCx5p33_ASAP7_75t_R g409 ( 
.A(n_51),
.Y(n_409)
);

INVx1_ASAP7_75t_L g410 ( 
.A(n_44),
.Y(n_410)
);

CKINVDCx5p33_ASAP7_75t_R g411 ( 
.A(n_160),
.Y(n_411)
);

INVx1_ASAP7_75t_L g412 ( 
.A(n_12),
.Y(n_412)
);

INVx2_ASAP7_75t_SL g413 ( 
.A(n_21),
.Y(n_413)
);

INVx1_ASAP7_75t_L g414 ( 
.A(n_33),
.Y(n_414)
);

BUFx5_ASAP7_75t_L g415 ( 
.A(n_0),
.Y(n_415)
);

INVx1_ASAP7_75t_L g416 ( 
.A(n_15),
.Y(n_416)
);

INVx1_ASAP7_75t_L g417 ( 
.A(n_372),
.Y(n_417)
);

CKINVDCx20_ASAP7_75t_R g418 ( 
.A(n_209),
.Y(n_418)
);

CKINVDCx5p33_ASAP7_75t_R g419 ( 
.A(n_318),
.Y(n_419)
);

BUFx6f_ASAP7_75t_SL g420 ( 
.A(n_291),
.Y(n_420)
);

INVx1_ASAP7_75t_L g421 ( 
.A(n_372),
.Y(n_421)
);

CKINVDCx5p33_ASAP7_75t_R g422 ( 
.A(n_384),
.Y(n_422)
);

CKINVDCx20_ASAP7_75t_R g423 ( 
.A(n_225),
.Y(n_423)
);

NOR2xp67_ASAP7_75t_L g424 ( 
.A(n_379),
.B(n_0),
.Y(n_424)
);

INVx1_ASAP7_75t_L g425 ( 
.A(n_372),
.Y(n_425)
);

CKINVDCx5p33_ASAP7_75t_R g426 ( 
.A(n_254),
.Y(n_426)
);

BUFx2_ASAP7_75t_L g427 ( 
.A(n_289),
.Y(n_427)
);

NOR2xp33_ASAP7_75t_L g428 ( 
.A(n_222),
.B(n_2),
.Y(n_428)
);

CKINVDCx5p33_ASAP7_75t_R g429 ( 
.A(n_261),
.Y(n_429)
);

INVx1_ASAP7_75t_L g430 ( 
.A(n_372),
.Y(n_430)
);

CKINVDCx5p33_ASAP7_75t_R g431 ( 
.A(n_265),
.Y(n_431)
);

CKINVDCx5p33_ASAP7_75t_R g432 ( 
.A(n_267),
.Y(n_432)
);

CKINVDCx5p33_ASAP7_75t_R g433 ( 
.A(n_278),
.Y(n_433)
);

INVx1_ASAP7_75t_L g434 ( 
.A(n_372),
.Y(n_434)
);

CKINVDCx16_ASAP7_75t_R g435 ( 
.A(n_329),
.Y(n_435)
);

CKINVDCx5p33_ASAP7_75t_R g436 ( 
.A(n_287),
.Y(n_436)
);

CKINVDCx20_ASAP7_75t_R g437 ( 
.A(n_228),
.Y(n_437)
);

CKINVDCx16_ASAP7_75t_R g438 ( 
.A(n_395),
.Y(n_438)
);

INVx1_ASAP7_75t_L g439 ( 
.A(n_372),
.Y(n_439)
);

CKINVDCx5p33_ASAP7_75t_R g440 ( 
.A(n_255),
.Y(n_440)
);

NOR2xp33_ASAP7_75t_L g441 ( 
.A(n_341),
.B(n_4),
.Y(n_441)
);

INVx1_ASAP7_75t_L g442 ( 
.A(n_372),
.Y(n_442)
);

INVx1_ASAP7_75t_L g443 ( 
.A(n_372),
.Y(n_443)
);

INVx1_ASAP7_75t_L g444 ( 
.A(n_415),
.Y(n_444)
);

INVx1_ASAP7_75t_L g445 ( 
.A(n_415),
.Y(n_445)
);

CKINVDCx5p33_ASAP7_75t_R g446 ( 
.A(n_295),
.Y(n_446)
);

CKINVDCx5p33_ASAP7_75t_R g447 ( 
.A(n_258),
.Y(n_447)
);

INVx1_ASAP7_75t_L g448 ( 
.A(n_415),
.Y(n_448)
);

INVx1_ASAP7_75t_L g449 ( 
.A(n_415),
.Y(n_449)
);

INVx1_ASAP7_75t_L g450 ( 
.A(n_415),
.Y(n_450)
);

INVx1_ASAP7_75t_L g451 ( 
.A(n_415),
.Y(n_451)
);

CKINVDCx5p33_ASAP7_75t_R g452 ( 
.A(n_260),
.Y(n_452)
);

CKINVDCx20_ASAP7_75t_R g453 ( 
.A(n_229),
.Y(n_453)
);

CKINVDCx20_ASAP7_75t_R g454 ( 
.A(n_268),
.Y(n_454)
);

INVx1_ASAP7_75t_L g455 ( 
.A(n_415),
.Y(n_455)
);

CKINVDCx20_ASAP7_75t_R g456 ( 
.A(n_284),
.Y(n_456)
);

INVx1_ASAP7_75t_L g457 ( 
.A(n_415),
.Y(n_457)
);

CKINVDCx5p33_ASAP7_75t_R g458 ( 
.A(n_262),
.Y(n_458)
);

INVx1_ASAP7_75t_L g459 ( 
.A(n_297),
.Y(n_459)
);

NAND2xp5_ASAP7_75t_L g460 ( 
.A(n_213),
.B(n_5),
.Y(n_460)
);

INVx2_ASAP7_75t_L g461 ( 
.A(n_303),
.Y(n_461)
);

CKINVDCx20_ASAP7_75t_R g462 ( 
.A(n_286),
.Y(n_462)
);

BUFx6f_ASAP7_75t_L g463 ( 
.A(n_211),
.Y(n_463)
);

BUFx6f_ASAP7_75t_L g464 ( 
.A(n_211),
.Y(n_464)
);

INVx1_ASAP7_75t_L g465 ( 
.A(n_297),
.Y(n_465)
);

INVx1_ASAP7_75t_L g466 ( 
.A(n_407),
.Y(n_466)
);

NOR2xp33_ASAP7_75t_L g467 ( 
.A(n_213),
.B(n_5),
.Y(n_467)
);

INVx1_ASAP7_75t_L g468 ( 
.A(n_407),
.Y(n_468)
);

INVx1_ASAP7_75t_L g469 ( 
.A(n_303),
.Y(n_469)
);

CKINVDCx20_ASAP7_75t_R g470 ( 
.A(n_324),
.Y(n_470)
);

CKINVDCx20_ASAP7_75t_R g471 ( 
.A(n_266),
.Y(n_471)
);

INVxp67_ASAP7_75t_SL g472 ( 
.A(n_311),
.Y(n_472)
);

CKINVDCx5p33_ASAP7_75t_R g473 ( 
.A(n_271),
.Y(n_473)
);

HB1xp67_ASAP7_75t_L g474 ( 
.A(n_234),
.Y(n_474)
);

HB1xp67_ASAP7_75t_L g475 ( 
.A(n_366),
.Y(n_475)
);

CKINVDCx20_ASAP7_75t_R g476 ( 
.A(n_273),
.Y(n_476)
);

INVx1_ASAP7_75t_L g477 ( 
.A(n_303),
.Y(n_477)
);

CKINVDCx5p33_ASAP7_75t_R g478 ( 
.A(n_300),
.Y(n_478)
);

INVx1_ASAP7_75t_L g479 ( 
.A(n_303),
.Y(n_479)
);

CKINVDCx20_ASAP7_75t_R g480 ( 
.A(n_275),
.Y(n_480)
);

INVx1_ASAP7_75t_L g481 ( 
.A(n_303),
.Y(n_481)
);

CKINVDCx5p33_ASAP7_75t_R g482 ( 
.A(n_321),
.Y(n_482)
);

CKINVDCx20_ASAP7_75t_R g483 ( 
.A(n_277),
.Y(n_483)
);

CKINVDCx20_ASAP7_75t_R g484 ( 
.A(n_285),
.Y(n_484)
);

INVx1_ASAP7_75t_L g485 ( 
.A(n_215),
.Y(n_485)
);

INVx1_ASAP7_75t_L g486 ( 
.A(n_237),
.Y(n_486)
);

CKINVDCx5p33_ASAP7_75t_R g487 ( 
.A(n_328),
.Y(n_487)
);

NOR2xp33_ASAP7_75t_L g488 ( 
.A(n_212),
.B(n_6),
.Y(n_488)
);

BUFx6f_ASAP7_75t_SL g489 ( 
.A(n_291),
.Y(n_489)
);

CKINVDCx5p33_ASAP7_75t_R g490 ( 
.A(n_331),
.Y(n_490)
);

BUFx3_ASAP7_75t_L g491 ( 
.A(n_311),
.Y(n_491)
);

INVxp67_ASAP7_75t_L g492 ( 
.A(n_243),
.Y(n_492)
);

CKINVDCx5p33_ASAP7_75t_R g493 ( 
.A(n_334),
.Y(n_493)
);

CKINVDCx16_ASAP7_75t_R g494 ( 
.A(n_291),
.Y(n_494)
);

INVx1_ASAP7_75t_L g495 ( 
.A(n_250),
.Y(n_495)
);

INVx1_ASAP7_75t_L g496 ( 
.A(n_252),
.Y(n_496)
);

NOR2xp67_ASAP7_75t_L g497 ( 
.A(n_403),
.B(n_8),
.Y(n_497)
);

CKINVDCx20_ASAP7_75t_R g498 ( 
.A(n_293),
.Y(n_498)
);

CKINVDCx5p33_ASAP7_75t_R g499 ( 
.A(n_339),
.Y(n_499)
);

HB1xp67_ASAP7_75t_L g500 ( 
.A(n_217),
.Y(n_500)
);

NOR2xp33_ASAP7_75t_L g501 ( 
.A(n_235),
.B(n_11),
.Y(n_501)
);

INVxp67_ASAP7_75t_SL g502 ( 
.A(n_319),
.Y(n_502)
);

CKINVDCx20_ASAP7_75t_R g503 ( 
.A(n_299),
.Y(n_503)
);

INVx1_ASAP7_75t_L g504 ( 
.A(n_269),
.Y(n_504)
);

CKINVDCx5p33_ASAP7_75t_R g505 ( 
.A(n_346),
.Y(n_505)
);

NAND2xp5_ASAP7_75t_L g506 ( 
.A(n_319),
.B(n_13),
.Y(n_506)
);

CKINVDCx20_ASAP7_75t_R g507 ( 
.A(n_301),
.Y(n_507)
);

CKINVDCx5p33_ASAP7_75t_R g508 ( 
.A(n_348),
.Y(n_508)
);

INVx3_ASAP7_75t_L g509 ( 
.A(n_368),
.Y(n_509)
);

INVx1_ASAP7_75t_L g510 ( 
.A(n_270),
.Y(n_510)
);

INVx1_ASAP7_75t_L g511 ( 
.A(n_274),
.Y(n_511)
);

CKINVDCx5p33_ASAP7_75t_R g512 ( 
.A(n_217),
.Y(n_512)
);

CKINVDCx5p33_ASAP7_75t_R g513 ( 
.A(n_220),
.Y(n_513)
);

CKINVDCx20_ASAP7_75t_R g514 ( 
.A(n_302),
.Y(n_514)
);

HB1xp67_ASAP7_75t_L g515 ( 
.A(n_220),
.Y(n_515)
);

CKINVDCx5p33_ASAP7_75t_R g516 ( 
.A(n_223),
.Y(n_516)
);

NAND2xp33_ASAP7_75t_R g517 ( 
.A(n_214),
.B(n_14),
.Y(n_517)
);

NOR2xp33_ASAP7_75t_L g518 ( 
.A(n_296),
.B(n_16),
.Y(n_518)
);

CKINVDCx5p33_ASAP7_75t_R g519 ( 
.A(n_223),
.Y(n_519)
);

INVx1_ASAP7_75t_L g520 ( 
.A(n_280),
.Y(n_520)
);

CKINVDCx5p33_ASAP7_75t_R g521 ( 
.A(n_233),
.Y(n_521)
);

CKINVDCx20_ASAP7_75t_R g522 ( 
.A(n_310),
.Y(n_522)
);

INVx1_ASAP7_75t_L g523 ( 
.A(n_283),
.Y(n_523)
);

CKINVDCx5p33_ASAP7_75t_R g524 ( 
.A(n_233),
.Y(n_524)
);

INVx2_ASAP7_75t_L g525 ( 
.A(n_461),
.Y(n_525)
);

NOR2x1_ASAP7_75t_L g526 ( 
.A(n_460),
.B(n_368),
.Y(n_526)
);

CKINVDCx5p33_ASAP7_75t_R g527 ( 
.A(n_440),
.Y(n_527)
);

CKINVDCx5p33_ASAP7_75t_R g528 ( 
.A(n_447),
.Y(n_528)
);

CKINVDCx5p33_ASAP7_75t_R g529 ( 
.A(n_452),
.Y(n_529)
);

AND2x2_ASAP7_75t_L g530 ( 
.A(n_472),
.B(n_257),
.Y(n_530)
);

INVx2_ASAP7_75t_L g531 ( 
.A(n_461),
.Y(n_531)
);

INVx2_ASAP7_75t_L g532 ( 
.A(n_469),
.Y(n_532)
);

BUFx3_ASAP7_75t_L g533 ( 
.A(n_491),
.Y(n_533)
);

CKINVDCx5p33_ASAP7_75t_R g534 ( 
.A(n_458),
.Y(n_534)
);

INVx3_ASAP7_75t_L g535 ( 
.A(n_463),
.Y(n_535)
);

INVx5_ASAP7_75t_L g536 ( 
.A(n_463),
.Y(n_536)
);

CKINVDCx5p33_ASAP7_75t_R g537 ( 
.A(n_473),
.Y(n_537)
);

NAND2xp5_ASAP7_75t_L g538 ( 
.A(n_502),
.B(n_210),
.Y(n_538)
);

CKINVDCx5p33_ASAP7_75t_R g539 ( 
.A(n_471),
.Y(n_539)
);

INVx1_ASAP7_75t_L g540 ( 
.A(n_477),
.Y(n_540)
);

BUFx6f_ASAP7_75t_L g541 ( 
.A(n_463),
.Y(n_541)
);

AND2x2_ASAP7_75t_L g542 ( 
.A(n_491),
.B(n_257),
.Y(n_542)
);

BUFx8_ASAP7_75t_L g543 ( 
.A(n_420),
.Y(n_543)
);

INVx1_ASAP7_75t_L g544 ( 
.A(n_479),
.Y(n_544)
);

AND2x2_ASAP7_75t_L g545 ( 
.A(n_459),
.B(n_413),
.Y(n_545)
);

NOR2xp33_ASAP7_75t_SL g546 ( 
.A(n_435),
.B(n_292),
.Y(n_546)
);

INVx2_ASAP7_75t_L g547 ( 
.A(n_463),
.Y(n_547)
);

CKINVDCx20_ASAP7_75t_R g548 ( 
.A(n_418),
.Y(n_548)
);

NOR2xp33_ASAP7_75t_SL g549 ( 
.A(n_438),
.B(n_292),
.Y(n_549)
);

INVx1_ASAP7_75t_L g550 ( 
.A(n_481),
.Y(n_550)
);

CKINVDCx5p33_ASAP7_75t_R g551 ( 
.A(n_476),
.Y(n_551)
);

AND2x4_ASAP7_75t_L g552 ( 
.A(n_509),
.B(n_218),
.Y(n_552)
);

NAND2xp5_ASAP7_75t_L g553 ( 
.A(n_509),
.B(n_219),
.Y(n_553)
);

INVx1_ASAP7_75t_L g554 ( 
.A(n_417),
.Y(n_554)
);

HB1xp67_ASAP7_75t_L g555 ( 
.A(n_422),
.Y(n_555)
);

AND2x4_ASAP7_75t_SL g556 ( 
.A(n_480),
.B(n_292),
.Y(n_556)
);

NOR2xp33_ASAP7_75t_R g557 ( 
.A(n_483),
.B(n_312),
.Y(n_557)
);

AND2x2_ASAP7_75t_L g558 ( 
.A(n_465),
.B(n_413),
.Y(n_558)
);

INVx1_ASAP7_75t_L g559 ( 
.A(n_421),
.Y(n_559)
);

CKINVDCx5p33_ASAP7_75t_R g560 ( 
.A(n_484),
.Y(n_560)
);

INVx1_ASAP7_75t_L g561 ( 
.A(n_425),
.Y(n_561)
);

NAND2xp5_ASAP7_75t_L g562 ( 
.A(n_509),
.B(n_224),
.Y(n_562)
);

INVx1_ASAP7_75t_L g563 ( 
.A(n_430),
.Y(n_563)
);

BUFx6f_ASAP7_75t_L g564 ( 
.A(n_463),
.Y(n_564)
);

CKINVDCx5p33_ASAP7_75t_R g565 ( 
.A(n_498),
.Y(n_565)
);

INVx1_ASAP7_75t_L g566 ( 
.A(n_434),
.Y(n_566)
);

CKINVDCx16_ASAP7_75t_R g567 ( 
.A(n_494),
.Y(n_567)
);

INVx2_ASAP7_75t_L g568 ( 
.A(n_464),
.Y(n_568)
);

CKINVDCx20_ASAP7_75t_R g569 ( 
.A(n_423),
.Y(n_569)
);

INVx1_ASAP7_75t_L g570 ( 
.A(n_439),
.Y(n_570)
);

NAND2xp5_ASAP7_75t_L g571 ( 
.A(n_466),
.B(n_227),
.Y(n_571)
);

CKINVDCx5p33_ASAP7_75t_R g572 ( 
.A(n_503),
.Y(n_572)
);

INVx1_ASAP7_75t_L g573 ( 
.A(n_442),
.Y(n_573)
);

CKINVDCx20_ASAP7_75t_R g574 ( 
.A(n_437),
.Y(n_574)
);

INVx2_ASAP7_75t_L g575 ( 
.A(n_464),
.Y(n_575)
);

NAND2xp5_ASAP7_75t_SL g576 ( 
.A(n_419),
.B(n_344),
.Y(n_576)
);

CKINVDCx5p33_ASAP7_75t_R g577 ( 
.A(n_507),
.Y(n_577)
);

CKINVDCx5p33_ASAP7_75t_R g578 ( 
.A(n_514),
.Y(n_578)
);

CKINVDCx5p33_ASAP7_75t_R g579 ( 
.A(n_522),
.Y(n_579)
);

AND2x4_ASAP7_75t_L g580 ( 
.A(n_443),
.B(n_230),
.Y(n_580)
);

INVx1_ASAP7_75t_L g581 ( 
.A(n_444),
.Y(n_581)
);

NAND2xp5_ASAP7_75t_L g582 ( 
.A(n_468),
.B(n_445),
.Y(n_582)
);

NAND2xp5_ASAP7_75t_L g583 ( 
.A(n_448),
.B(n_231),
.Y(n_583)
);

INVx1_ASAP7_75t_L g584 ( 
.A(n_449),
.Y(n_584)
);

CKINVDCx5p33_ASAP7_75t_R g585 ( 
.A(n_426),
.Y(n_585)
);

BUFx3_ASAP7_75t_L g586 ( 
.A(n_464),
.Y(n_586)
);

INVx1_ASAP7_75t_L g587 ( 
.A(n_450),
.Y(n_587)
);

INVx1_ASAP7_75t_L g588 ( 
.A(n_451),
.Y(n_588)
);

INVx1_ASAP7_75t_L g589 ( 
.A(n_455),
.Y(n_589)
);

OAI22xp5_ASAP7_75t_SL g590 ( 
.A1(n_453),
.A2(n_386),
.B1(n_336),
.B2(n_309),
.Y(n_590)
);

CKINVDCx5p33_ASAP7_75t_R g591 ( 
.A(n_426),
.Y(n_591)
);

CKINVDCx5p33_ASAP7_75t_R g592 ( 
.A(n_429),
.Y(n_592)
);

INVx2_ASAP7_75t_L g593 ( 
.A(n_464),
.Y(n_593)
);

BUFx6f_ASAP7_75t_L g594 ( 
.A(n_464),
.Y(n_594)
);

INVx1_ASAP7_75t_L g595 ( 
.A(n_457),
.Y(n_595)
);

NOR2xp33_ASAP7_75t_R g596 ( 
.A(n_429),
.B(n_314),
.Y(n_596)
);

AND2x2_ASAP7_75t_L g597 ( 
.A(n_485),
.B(n_307),
.Y(n_597)
);

INVx1_ASAP7_75t_L g598 ( 
.A(n_486),
.Y(n_598)
);

INVx1_ASAP7_75t_L g599 ( 
.A(n_495),
.Y(n_599)
);

INVx3_ASAP7_75t_L g600 ( 
.A(n_496),
.Y(n_600)
);

CKINVDCx5p33_ASAP7_75t_R g601 ( 
.A(n_431),
.Y(n_601)
);

NOR2xp33_ASAP7_75t_L g602 ( 
.A(n_419),
.B(n_349),
.Y(n_602)
);

CKINVDCx20_ASAP7_75t_R g603 ( 
.A(n_454),
.Y(n_603)
);

NAND2xp5_ASAP7_75t_L g604 ( 
.A(n_431),
.B(n_232),
.Y(n_604)
);

INVx2_ASAP7_75t_L g605 ( 
.A(n_504),
.Y(n_605)
);

AND3x1_ASAP7_75t_L g606 ( 
.A(n_428),
.B(n_308),
.C(n_307),
.Y(n_606)
);

INVx1_ASAP7_75t_L g607 ( 
.A(n_510),
.Y(n_607)
);

INVx1_ASAP7_75t_L g608 ( 
.A(n_511),
.Y(n_608)
);

BUFx2_ASAP7_75t_L g609 ( 
.A(n_422),
.Y(n_609)
);

CKINVDCx5p33_ASAP7_75t_R g610 ( 
.A(n_432),
.Y(n_610)
);

BUFx3_ASAP7_75t_L g611 ( 
.A(n_533),
.Y(n_611)
);

BUFx2_ASAP7_75t_L g612 ( 
.A(n_533),
.Y(n_612)
);

INVx2_ASAP7_75t_L g613 ( 
.A(n_531),
.Y(n_613)
);

INVx2_ASAP7_75t_L g614 ( 
.A(n_531),
.Y(n_614)
);

NOR2xp33_ASAP7_75t_L g615 ( 
.A(n_602),
.B(n_432),
.Y(n_615)
);

INVx4_ASAP7_75t_L g616 ( 
.A(n_541),
.Y(n_616)
);

INVx1_ASAP7_75t_L g617 ( 
.A(n_554),
.Y(n_617)
);

NAND2xp5_ASAP7_75t_L g618 ( 
.A(n_530),
.B(n_433),
.Y(n_618)
);

INVx1_ASAP7_75t_L g619 ( 
.A(n_554),
.Y(n_619)
);

AOI22xp5_ASAP7_75t_L g620 ( 
.A1(n_606),
.A2(n_501),
.B1(n_518),
.B2(n_488),
.Y(n_620)
);

INVxp67_ASAP7_75t_SL g621 ( 
.A(n_533),
.Y(n_621)
);

BUFx6f_ASAP7_75t_L g622 ( 
.A(n_541),
.Y(n_622)
);

NOR2xp33_ASAP7_75t_L g623 ( 
.A(n_604),
.B(n_433),
.Y(n_623)
);

INVx3_ASAP7_75t_L g624 ( 
.A(n_541),
.Y(n_624)
);

NAND2xp5_ASAP7_75t_SL g625 ( 
.A(n_596),
.B(n_436),
.Y(n_625)
);

BUFx3_ASAP7_75t_L g626 ( 
.A(n_580),
.Y(n_626)
);

INVx3_ASAP7_75t_L g627 ( 
.A(n_541),
.Y(n_627)
);

BUFx3_ASAP7_75t_L g628 ( 
.A(n_580),
.Y(n_628)
);

NOR2xp33_ASAP7_75t_L g629 ( 
.A(n_527),
.B(n_436),
.Y(n_629)
);

NAND2xp5_ASAP7_75t_L g630 ( 
.A(n_530),
.B(n_446),
.Y(n_630)
);

NAND2xp5_ASAP7_75t_L g631 ( 
.A(n_559),
.B(n_446),
.Y(n_631)
);

INVx1_ASAP7_75t_L g632 ( 
.A(n_559),
.Y(n_632)
);

INVx1_ASAP7_75t_SL g633 ( 
.A(n_609),
.Y(n_633)
);

AND2x2_ASAP7_75t_SL g634 ( 
.A(n_556),
.B(n_546),
.Y(n_634)
);

NAND2xp5_ASAP7_75t_L g635 ( 
.A(n_561),
.B(n_478),
.Y(n_635)
);

INVx2_ASAP7_75t_SL g636 ( 
.A(n_542),
.Y(n_636)
);

INVx1_ASAP7_75t_L g637 ( 
.A(n_561),
.Y(n_637)
);

NOR2xp33_ASAP7_75t_L g638 ( 
.A(n_528),
.B(n_478),
.Y(n_638)
);

NAND2xp5_ASAP7_75t_L g639 ( 
.A(n_563),
.B(n_482),
.Y(n_639)
);

NAND2xp5_ASAP7_75t_L g640 ( 
.A(n_563),
.B(n_482),
.Y(n_640)
);

NAND2xp5_ASAP7_75t_L g641 ( 
.A(n_566),
.B(n_487),
.Y(n_641)
);

NAND2xp5_ASAP7_75t_L g642 ( 
.A(n_566),
.B(n_487),
.Y(n_642)
);

NAND2xp5_ASAP7_75t_SL g643 ( 
.A(n_549),
.B(n_490),
.Y(n_643)
);

AND2x6_ASAP7_75t_L g644 ( 
.A(n_580),
.B(n_211),
.Y(n_644)
);

INVx2_ASAP7_75t_L g645 ( 
.A(n_525),
.Y(n_645)
);

INVx2_ASAP7_75t_SL g646 ( 
.A(n_542),
.Y(n_646)
);

NOR2xp33_ASAP7_75t_SL g647 ( 
.A(n_567),
.B(n_456),
.Y(n_647)
);

INVx1_ASAP7_75t_L g648 ( 
.A(n_570),
.Y(n_648)
);

AOI22xp33_ASAP7_75t_L g649 ( 
.A1(n_580),
.A2(n_467),
.B1(n_427),
.B2(n_441),
.Y(n_649)
);

INVx3_ASAP7_75t_L g650 ( 
.A(n_541),
.Y(n_650)
);

AND2x2_ASAP7_75t_L g651 ( 
.A(n_545),
.B(n_500),
.Y(n_651)
);

NAND2xp5_ASAP7_75t_SL g652 ( 
.A(n_529),
.B(n_490),
.Y(n_652)
);

INVx2_ASAP7_75t_L g653 ( 
.A(n_525),
.Y(n_653)
);

NAND2xp5_ASAP7_75t_SL g654 ( 
.A(n_534),
.B(n_493),
.Y(n_654)
);

NAND2xp5_ASAP7_75t_SL g655 ( 
.A(n_537),
.B(n_493),
.Y(n_655)
);

NAND2xp5_ASAP7_75t_SL g656 ( 
.A(n_557),
.B(n_499),
.Y(n_656)
);

INVx1_ASAP7_75t_L g657 ( 
.A(n_570),
.Y(n_657)
);

INVx1_ASAP7_75t_L g658 ( 
.A(n_573),
.Y(n_658)
);

CKINVDCx5p33_ASAP7_75t_R g659 ( 
.A(n_539),
.Y(n_659)
);

INVx3_ASAP7_75t_L g660 ( 
.A(n_541),
.Y(n_660)
);

INVx4_ASAP7_75t_L g661 ( 
.A(n_564),
.Y(n_661)
);

INVx6_ASAP7_75t_L g662 ( 
.A(n_552),
.Y(n_662)
);

NOR2xp33_ASAP7_75t_L g663 ( 
.A(n_576),
.B(n_499),
.Y(n_663)
);

AND2x4_ASAP7_75t_L g664 ( 
.A(n_552),
.B(n_526),
.Y(n_664)
);

CKINVDCx5p33_ASAP7_75t_R g665 ( 
.A(n_551),
.Y(n_665)
);

INVx3_ASAP7_75t_L g666 ( 
.A(n_564),
.Y(n_666)
);

AOI22xp33_ASAP7_75t_L g667 ( 
.A1(n_526),
.A2(n_506),
.B1(n_308),
.B2(n_315),
.Y(n_667)
);

INVx4_ASAP7_75t_L g668 ( 
.A(n_564),
.Y(n_668)
);

NAND2xp5_ASAP7_75t_SL g669 ( 
.A(n_543),
.B(n_505),
.Y(n_669)
);

NAND2xp5_ASAP7_75t_L g670 ( 
.A(n_573),
.B(n_505),
.Y(n_670)
);

BUFx2_ASAP7_75t_L g671 ( 
.A(n_609),
.Y(n_671)
);

NAND2xp5_ASAP7_75t_SL g672 ( 
.A(n_543),
.B(n_508),
.Y(n_672)
);

NAND2xp5_ASAP7_75t_L g673 ( 
.A(n_581),
.B(n_508),
.Y(n_673)
);

AND2x6_ASAP7_75t_L g674 ( 
.A(n_552),
.B(n_211),
.Y(n_674)
);

AND2x2_ASAP7_75t_L g675 ( 
.A(n_545),
.B(n_515),
.Y(n_675)
);

INVx2_ASAP7_75t_L g676 ( 
.A(n_532),
.Y(n_676)
);

INVx2_ASAP7_75t_L g677 ( 
.A(n_532),
.Y(n_677)
);

OAI22xp33_ASAP7_75t_L g678 ( 
.A1(n_538),
.A2(n_517),
.B1(n_281),
.B2(n_276),
.Y(n_678)
);

NOR2xp33_ASAP7_75t_L g679 ( 
.A(n_585),
.B(n_512),
.Y(n_679)
);

BUFx6f_ASAP7_75t_L g680 ( 
.A(n_564),
.Y(n_680)
);

OR2x2_ASAP7_75t_L g681 ( 
.A(n_567),
.B(n_512),
.Y(n_681)
);

INVx1_ASAP7_75t_L g682 ( 
.A(n_581),
.Y(n_682)
);

NAND2xp5_ASAP7_75t_L g683 ( 
.A(n_584),
.B(n_350),
.Y(n_683)
);

NAND2xp5_ASAP7_75t_SL g684 ( 
.A(n_543),
.B(n_513),
.Y(n_684)
);

INVx1_ASAP7_75t_L g685 ( 
.A(n_584),
.Y(n_685)
);

INVx5_ASAP7_75t_L g686 ( 
.A(n_564),
.Y(n_686)
);

AOI22xp33_ASAP7_75t_L g687 ( 
.A1(n_552),
.A2(n_588),
.B1(n_589),
.B2(n_587),
.Y(n_687)
);

INVx1_ASAP7_75t_SL g688 ( 
.A(n_548),
.Y(n_688)
);

NAND2xp5_ASAP7_75t_L g689 ( 
.A(n_587),
.B(n_588),
.Y(n_689)
);

BUFx2_ASAP7_75t_L g690 ( 
.A(n_591),
.Y(n_690)
);

INVx1_ASAP7_75t_L g691 ( 
.A(n_589),
.Y(n_691)
);

INVx3_ASAP7_75t_L g692 ( 
.A(n_564),
.Y(n_692)
);

AOI22xp33_ASAP7_75t_L g693 ( 
.A1(n_595),
.A2(n_315),
.B1(n_474),
.B2(n_475),
.Y(n_693)
);

AOI22xp33_ASAP7_75t_L g694 ( 
.A1(n_595),
.A2(n_330),
.B1(n_375),
.B2(n_304),
.Y(n_694)
);

OR2x2_ASAP7_75t_L g695 ( 
.A(n_555),
.B(n_513),
.Y(n_695)
);

INVx1_ASAP7_75t_L g696 ( 
.A(n_600),
.Y(n_696)
);

INVx1_ASAP7_75t_SL g697 ( 
.A(n_569),
.Y(n_697)
);

INVx1_ASAP7_75t_L g698 ( 
.A(n_600),
.Y(n_698)
);

INVx1_ASAP7_75t_L g699 ( 
.A(n_598),
.Y(n_699)
);

AND2x4_ASAP7_75t_L g700 ( 
.A(n_597),
.B(n_520),
.Y(n_700)
);

NAND2xp5_ASAP7_75t_L g701 ( 
.A(n_535),
.B(n_365),
.Y(n_701)
);

BUFx4f_ASAP7_75t_L g702 ( 
.A(n_600),
.Y(n_702)
);

BUFx3_ASAP7_75t_L g703 ( 
.A(n_586),
.Y(n_703)
);

NOR2xp33_ASAP7_75t_L g704 ( 
.A(n_592),
.B(n_516),
.Y(n_704)
);

NOR2x1p5_ASAP7_75t_L g705 ( 
.A(n_601),
.B(n_516),
.Y(n_705)
);

INVx2_ASAP7_75t_L g706 ( 
.A(n_540),
.Y(n_706)
);

INVx4_ASAP7_75t_L g707 ( 
.A(n_594),
.Y(n_707)
);

BUFx3_ASAP7_75t_L g708 ( 
.A(n_586),
.Y(n_708)
);

AND2x4_ASAP7_75t_L g709 ( 
.A(n_597),
.B(n_523),
.Y(n_709)
);

OR2x2_ASAP7_75t_L g710 ( 
.A(n_582),
.B(n_519),
.Y(n_710)
);

BUFx8_ASAP7_75t_SL g711 ( 
.A(n_574),
.Y(n_711)
);

INVx1_ASAP7_75t_L g712 ( 
.A(n_600),
.Y(n_712)
);

INVx1_ASAP7_75t_L g713 ( 
.A(n_540),
.Y(n_713)
);

NOR2xp33_ASAP7_75t_L g714 ( 
.A(n_610),
.B(n_519),
.Y(n_714)
);

NAND2xp5_ASAP7_75t_SL g715 ( 
.A(n_543),
.B(n_521),
.Y(n_715)
);

BUFx2_ASAP7_75t_L g716 ( 
.A(n_560),
.Y(n_716)
);

INVx1_ASAP7_75t_L g717 ( 
.A(n_598),
.Y(n_717)
);

INVx1_ASAP7_75t_L g718 ( 
.A(n_599),
.Y(n_718)
);

OR2x2_ASAP7_75t_L g719 ( 
.A(n_558),
.B(n_521),
.Y(n_719)
);

INVx2_ASAP7_75t_L g720 ( 
.A(n_544),
.Y(n_720)
);

AND2x4_ASAP7_75t_L g721 ( 
.A(n_558),
.B(n_242),
.Y(n_721)
);

BUFx6f_ASAP7_75t_L g722 ( 
.A(n_594),
.Y(n_722)
);

NAND2xp5_ASAP7_75t_SL g723 ( 
.A(n_556),
.B(n_524),
.Y(n_723)
);

AND2x2_ASAP7_75t_L g724 ( 
.A(n_599),
.B(n_607),
.Y(n_724)
);

AND2x6_ASAP7_75t_L g725 ( 
.A(n_553),
.B(n_211),
.Y(n_725)
);

NAND2xp5_ASAP7_75t_L g726 ( 
.A(n_535),
.B(n_370),
.Y(n_726)
);

BUFx3_ASAP7_75t_L g727 ( 
.A(n_586),
.Y(n_727)
);

NAND2xp5_ASAP7_75t_L g728 ( 
.A(n_535),
.B(n_316),
.Y(n_728)
);

HB1xp67_ASAP7_75t_L g729 ( 
.A(n_607),
.Y(n_729)
);

NAND2xp5_ASAP7_75t_SL g730 ( 
.A(n_556),
.B(n_524),
.Y(n_730)
);

NOR2xp33_ASAP7_75t_L g731 ( 
.A(n_571),
.B(n_420),
.Y(n_731)
);

INVx1_ASAP7_75t_L g732 ( 
.A(n_544),
.Y(n_732)
);

OR2x6_ASAP7_75t_L g733 ( 
.A(n_608),
.B(n_424),
.Y(n_733)
);

NAND2xp5_ASAP7_75t_SL g734 ( 
.A(n_608),
.B(n_344),
.Y(n_734)
);

INVx2_ASAP7_75t_L g735 ( 
.A(n_550),
.Y(n_735)
);

INVx1_ASAP7_75t_L g736 ( 
.A(n_550),
.Y(n_736)
);

NAND2xp5_ASAP7_75t_L g737 ( 
.A(n_535),
.B(n_317),
.Y(n_737)
);

BUFx10_ASAP7_75t_L g738 ( 
.A(n_565),
.Y(n_738)
);

NAND2xp5_ASAP7_75t_L g739 ( 
.A(n_583),
.B(n_320),
.Y(n_739)
);

AOI22xp33_ASAP7_75t_L g740 ( 
.A1(n_562),
.A2(n_388),
.B1(n_306),
.B2(n_325),
.Y(n_740)
);

INVx2_ASAP7_75t_L g741 ( 
.A(n_547),
.Y(n_741)
);

INVx2_ASAP7_75t_SL g742 ( 
.A(n_605),
.Y(n_742)
);

INVx1_ASAP7_75t_L g743 ( 
.A(n_605),
.Y(n_743)
);

INVx1_ASAP7_75t_L g744 ( 
.A(n_547),
.Y(n_744)
);

AOI22xp33_ASAP7_75t_L g745 ( 
.A1(n_547),
.A2(n_288),
.B1(n_416),
.B2(n_414),
.Y(n_745)
);

AOI22xp33_ASAP7_75t_L g746 ( 
.A1(n_568),
.A2(n_393),
.B1(n_337),
.B2(n_338),
.Y(n_746)
);

INVx1_ASAP7_75t_L g747 ( 
.A(n_568),
.Y(n_747)
);

INVx1_ASAP7_75t_L g748 ( 
.A(n_568),
.Y(n_748)
);

BUFx2_ASAP7_75t_L g749 ( 
.A(n_572),
.Y(n_749)
);

BUFx3_ASAP7_75t_L g750 ( 
.A(n_594),
.Y(n_750)
);

INVx2_ASAP7_75t_L g751 ( 
.A(n_575),
.Y(n_751)
);

INVx1_ASAP7_75t_L g752 ( 
.A(n_575),
.Y(n_752)
);

AND2x2_ASAP7_75t_L g753 ( 
.A(n_593),
.B(n_492),
.Y(n_753)
);

OR2x2_ASAP7_75t_L g754 ( 
.A(n_590),
.B(n_364),
.Y(n_754)
);

CKINVDCx20_ASAP7_75t_R g755 ( 
.A(n_603),
.Y(n_755)
);

BUFx3_ASAP7_75t_L g756 ( 
.A(n_594),
.Y(n_756)
);

AND2x2_ASAP7_75t_L g757 ( 
.A(n_593),
.B(n_497),
.Y(n_757)
);

NOR2xp33_ASAP7_75t_L g758 ( 
.A(n_593),
.B(n_420),
.Y(n_758)
);

NOR2xp33_ASAP7_75t_L g759 ( 
.A(n_577),
.B(n_489),
.Y(n_759)
);

INVx4_ASAP7_75t_L g760 ( 
.A(n_594),
.Y(n_760)
);

INVx2_ASAP7_75t_SL g761 ( 
.A(n_578),
.Y(n_761)
);

NOR2x1p5_ASAP7_75t_L g762 ( 
.A(n_681),
.B(n_579),
.Y(n_762)
);

NOR2xp33_ASAP7_75t_SL g763 ( 
.A(n_634),
.B(n_629),
.Y(n_763)
);

NAND2xp5_ASAP7_75t_L g764 ( 
.A(n_636),
.B(n_353),
.Y(n_764)
);

INVx2_ASAP7_75t_L g765 ( 
.A(n_645),
.Y(n_765)
);

NAND2xp5_ASAP7_75t_SL g766 ( 
.A(n_664),
.B(n_248),
.Y(n_766)
);

NAND2xp5_ASAP7_75t_SL g767 ( 
.A(n_664),
.B(n_253),
.Y(n_767)
);

INVxp67_ASAP7_75t_L g768 ( 
.A(n_671),
.Y(n_768)
);

OAI22xp33_ASAP7_75t_L g769 ( 
.A1(n_620),
.A2(n_754),
.B1(n_646),
.B2(n_636),
.Y(n_769)
);

AOI22xp33_ASAP7_75t_L g770 ( 
.A1(n_617),
.A2(n_340),
.B1(n_332),
.B2(n_351),
.Y(n_770)
);

INVxp67_ASAP7_75t_L g771 ( 
.A(n_671),
.Y(n_771)
);

INVx1_ASAP7_75t_L g772 ( 
.A(n_724),
.Y(n_772)
);

NOR2xp33_ASAP7_75t_L g773 ( 
.A(n_618),
.B(n_214),
.Y(n_773)
);

NAND3xp33_ASAP7_75t_L g774 ( 
.A(n_615),
.B(n_221),
.C(n_216),
.Y(n_774)
);

INVx1_ASAP7_75t_L g775 ( 
.A(n_724),
.Y(n_775)
);

NAND2xp5_ASAP7_75t_SL g776 ( 
.A(n_664),
.B(n_256),
.Y(n_776)
);

BUFx3_ASAP7_75t_L g777 ( 
.A(n_611),
.Y(n_777)
);

AND2x6_ASAP7_75t_SL g778 ( 
.A(n_679),
.B(n_704),
.Y(n_778)
);

INVx1_ASAP7_75t_L g779 ( 
.A(n_699),
.Y(n_779)
);

INVx2_ASAP7_75t_L g780 ( 
.A(n_613),
.Y(n_780)
);

NAND2xp5_ASAP7_75t_L g781 ( 
.A(n_646),
.B(n_259),
.Y(n_781)
);

NAND2xp5_ASAP7_75t_L g782 ( 
.A(n_623),
.B(n_263),
.Y(n_782)
);

NOR2xp33_ASAP7_75t_R g783 ( 
.A(n_659),
.B(n_462),
.Y(n_783)
);

NOR2xp33_ASAP7_75t_L g784 ( 
.A(n_630),
.B(n_216),
.Y(n_784)
);

INVxp67_ASAP7_75t_L g785 ( 
.A(n_719),
.Y(n_785)
);

AOI22xp5_ASAP7_75t_L g786 ( 
.A1(n_663),
.A2(n_470),
.B1(n_333),
.B2(n_327),
.Y(n_786)
);

AOI22xp5_ASAP7_75t_L g787 ( 
.A1(n_631),
.A2(n_323),
.B1(n_335),
.B2(n_355),
.Y(n_787)
);

AND2x2_ASAP7_75t_L g788 ( 
.A(n_651),
.B(n_240),
.Y(n_788)
);

NAND2xp5_ASAP7_75t_SL g789 ( 
.A(n_626),
.B(n_264),
.Y(n_789)
);

NOR2xp33_ASAP7_75t_L g790 ( 
.A(n_710),
.B(n_635),
.Y(n_790)
);

INVx2_ASAP7_75t_SL g791 ( 
.A(n_700),
.Y(n_791)
);

INVx1_ASAP7_75t_L g792 ( 
.A(n_717),
.Y(n_792)
);

NAND2xp5_ASAP7_75t_SL g793 ( 
.A(n_626),
.B(n_272),
.Y(n_793)
);

INVx1_ASAP7_75t_L g794 ( 
.A(n_718),
.Y(n_794)
);

NAND2xp5_ASAP7_75t_L g795 ( 
.A(n_617),
.B(n_619),
.Y(n_795)
);

NAND2xp5_ASAP7_75t_L g796 ( 
.A(n_619),
.B(n_279),
.Y(n_796)
);

NAND2xp5_ASAP7_75t_SL g797 ( 
.A(n_628),
.B(n_282),
.Y(n_797)
);

AOI22xp5_ASAP7_75t_L g798 ( 
.A1(n_639),
.A2(n_342),
.B1(n_354),
.B2(n_345),
.Y(n_798)
);

INVx1_ASAP7_75t_L g799 ( 
.A(n_628),
.Y(n_799)
);

INVx4_ASAP7_75t_L g800 ( 
.A(n_662),
.Y(n_800)
);

NAND2xp5_ASAP7_75t_SL g801 ( 
.A(n_696),
.B(n_290),
.Y(n_801)
);

NAND2xp5_ASAP7_75t_L g802 ( 
.A(n_632),
.B(n_294),
.Y(n_802)
);

NOR2xp33_ASAP7_75t_L g803 ( 
.A(n_710),
.B(n_221),
.Y(n_803)
);

INVxp33_ASAP7_75t_L g804 ( 
.A(n_711),
.Y(n_804)
);

NAND2xp5_ASAP7_75t_L g805 ( 
.A(n_632),
.B(n_305),
.Y(n_805)
);

INVx2_ASAP7_75t_L g806 ( 
.A(n_614),
.Y(n_806)
);

INVx2_ASAP7_75t_L g807 ( 
.A(n_614),
.Y(n_807)
);

INVx2_ASAP7_75t_L g808 ( 
.A(n_706),
.Y(n_808)
);

AOI22xp5_ASAP7_75t_L g809 ( 
.A1(n_640),
.A2(n_343),
.B1(n_362),
.B2(n_363),
.Y(n_809)
);

NAND2xp5_ASAP7_75t_SL g810 ( 
.A(n_696),
.B(n_322),
.Y(n_810)
);

AND2x4_ASAP7_75t_L g811 ( 
.A(n_611),
.B(n_621),
.Y(n_811)
);

INVx2_ASAP7_75t_L g812 ( 
.A(n_653),
.Y(n_812)
);

BUFx6f_ASAP7_75t_L g813 ( 
.A(n_703),
.Y(n_813)
);

NAND2xp5_ASAP7_75t_L g814 ( 
.A(n_648),
.B(n_326),
.Y(n_814)
);

NAND2xp5_ASAP7_75t_L g815 ( 
.A(n_648),
.B(n_347),
.Y(n_815)
);

NAND2xp5_ASAP7_75t_SL g816 ( 
.A(n_698),
.B(n_359),
.Y(n_816)
);

NAND2xp5_ASAP7_75t_L g817 ( 
.A(n_685),
.B(n_361),
.Y(n_817)
);

NAND2xp5_ASAP7_75t_L g818 ( 
.A(n_685),
.B(n_369),
.Y(n_818)
);

NAND2xp5_ASAP7_75t_L g819 ( 
.A(n_691),
.B(n_376),
.Y(n_819)
);

NOR2xp67_ASAP7_75t_L g820 ( 
.A(n_638),
.B(n_226),
.Y(n_820)
);

INVx1_ASAP7_75t_L g821 ( 
.A(n_713),
.Y(n_821)
);

NOR2x1p5_ASAP7_75t_L g822 ( 
.A(n_681),
.B(n_240),
.Y(n_822)
);

INVx2_ASAP7_75t_L g823 ( 
.A(n_676),
.Y(n_823)
);

NAND2xp5_ASAP7_75t_SL g824 ( 
.A(n_698),
.B(n_712),
.Y(n_824)
);

NAND2xp33_ASAP7_75t_L g825 ( 
.A(n_644),
.B(n_226),
.Y(n_825)
);

NAND2xp5_ASAP7_75t_SL g826 ( 
.A(n_712),
.B(n_687),
.Y(n_826)
);

NOR2xp33_ASAP7_75t_L g827 ( 
.A(n_641),
.B(n_236),
.Y(n_827)
);

HB1xp67_ASAP7_75t_L g828 ( 
.A(n_612),
.Y(n_828)
);

NAND2xp5_ASAP7_75t_SL g829 ( 
.A(n_702),
.B(n_377),
.Y(n_829)
);

NAND2xp5_ASAP7_75t_L g830 ( 
.A(n_691),
.B(n_637),
.Y(n_830)
);

INVx2_ASAP7_75t_L g831 ( 
.A(n_706),
.Y(n_831)
);

INVx4_ASAP7_75t_L g832 ( 
.A(n_662),
.Y(n_832)
);

NAND2xp5_ASAP7_75t_L g833 ( 
.A(n_657),
.B(n_383),
.Y(n_833)
);

OAI22xp33_ASAP7_75t_L g834 ( 
.A1(n_754),
.A2(n_371),
.B1(n_358),
.B2(n_357),
.Y(n_834)
);

NAND2xp5_ASAP7_75t_SL g835 ( 
.A(n_702),
.B(n_390),
.Y(n_835)
);

O2A1O1Ixp5_ASAP7_75t_L g836 ( 
.A1(n_658),
.A2(n_396),
.B(n_391),
.C(n_408),
.Y(n_836)
);

INVx2_ASAP7_75t_L g837 ( 
.A(n_720),
.Y(n_837)
);

AOI22xp33_ASAP7_75t_L g838 ( 
.A1(n_667),
.A2(n_352),
.B1(n_397),
.B2(n_404),
.Y(n_838)
);

HB1xp67_ASAP7_75t_L g839 ( 
.A(n_612),
.Y(n_839)
);

NOR2xp33_ASAP7_75t_L g840 ( 
.A(n_642),
.B(n_236),
.Y(n_840)
);

NAND2xp5_ASAP7_75t_SL g841 ( 
.A(n_702),
.B(n_238),
.Y(n_841)
);

NOR2xp33_ASAP7_75t_L g842 ( 
.A(n_670),
.B(n_238),
.Y(n_842)
);

INVx1_ASAP7_75t_L g843 ( 
.A(n_732),
.Y(n_843)
);

INVxp67_ASAP7_75t_L g844 ( 
.A(n_719),
.Y(n_844)
);

OR2x2_ASAP7_75t_L g845 ( 
.A(n_695),
.B(n_590),
.Y(n_845)
);

BUFx3_ASAP7_75t_L g846 ( 
.A(n_662),
.Y(n_846)
);

NOR2xp67_ASAP7_75t_SL g847 ( 
.A(n_662),
.B(n_536),
.Y(n_847)
);

NOR2x1p5_ASAP7_75t_L g848 ( 
.A(n_695),
.B(n_241),
.Y(n_848)
);

OAI21xp5_ASAP7_75t_L g849 ( 
.A1(n_689),
.A2(n_239),
.B(n_378),
.Y(n_849)
);

AOI22xp5_ASAP7_75t_L g850 ( 
.A1(n_673),
.A2(n_721),
.B1(n_651),
.B2(n_675),
.Y(n_850)
);

AO22x1_ASAP7_75t_L g851 ( 
.A1(n_675),
.A2(n_406),
.B1(n_356),
.B2(n_313),
.Y(n_851)
);

OR2x6_ASAP7_75t_L g852 ( 
.A(n_761),
.B(n_716),
.Y(n_852)
);

INVx3_ASAP7_75t_L g853 ( 
.A(n_703),
.Y(n_853)
);

NOR2xp33_ASAP7_75t_L g854 ( 
.A(n_729),
.B(n_239),
.Y(n_854)
);

INVx2_ASAP7_75t_SL g855 ( 
.A(n_700),
.Y(n_855)
);

NAND2xp5_ASAP7_75t_L g856 ( 
.A(n_682),
.B(n_594),
.Y(n_856)
);

NOR2x1_ASAP7_75t_L g857 ( 
.A(n_656),
.B(n_405),
.Y(n_857)
);

INVx2_ASAP7_75t_SL g858 ( 
.A(n_700),
.Y(n_858)
);

AND2x2_ASAP7_75t_SL g859 ( 
.A(n_634),
.B(n_649),
.Y(n_859)
);

BUFx3_ASAP7_75t_L g860 ( 
.A(n_708),
.Y(n_860)
);

NAND2xp5_ASAP7_75t_L g861 ( 
.A(n_739),
.B(n_244),
.Y(n_861)
);

BUFx8_ASAP7_75t_L g862 ( 
.A(n_716),
.Y(n_862)
);

INVx2_ASAP7_75t_L g863 ( 
.A(n_720),
.Y(n_863)
);

INVx1_ASAP7_75t_L g864 ( 
.A(n_736),
.Y(n_864)
);

NAND2xp5_ASAP7_75t_SL g865 ( 
.A(n_678),
.B(n_244),
.Y(n_865)
);

NAND2xp5_ASAP7_75t_SL g866 ( 
.A(n_683),
.B(n_245),
.Y(n_866)
);

INVxp67_ASAP7_75t_L g867 ( 
.A(n_714),
.Y(n_867)
);

AOI22xp5_ASAP7_75t_L g868 ( 
.A1(n_721),
.A2(n_733),
.B1(n_643),
.B2(n_709),
.Y(n_868)
);

NAND2xp5_ASAP7_75t_L g869 ( 
.A(n_757),
.B(n_245),
.Y(n_869)
);

NAND2xp5_ASAP7_75t_L g870 ( 
.A(n_757),
.B(n_246),
.Y(n_870)
);

BUFx6f_ASAP7_75t_L g871 ( 
.A(n_708),
.Y(n_871)
);

INVx2_ASAP7_75t_SL g872 ( 
.A(n_709),
.Y(n_872)
);

AOI22xp33_ASAP7_75t_L g873 ( 
.A1(n_721),
.A2(n_410),
.B1(n_412),
.B2(n_241),
.Y(n_873)
);

INVx2_ASAP7_75t_L g874 ( 
.A(n_676),
.Y(n_874)
);

AND2x2_ASAP7_75t_L g875 ( 
.A(n_633),
.B(n_247),
.Y(n_875)
);

INVx1_ASAP7_75t_L g876 ( 
.A(n_736),
.Y(n_876)
);

NAND2xp5_ASAP7_75t_L g877 ( 
.A(n_742),
.B(n_246),
.Y(n_877)
);

NOR2xp33_ASAP7_75t_L g878 ( 
.A(n_625),
.B(n_251),
.Y(n_878)
);

BUFx8_ASAP7_75t_L g879 ( 
.A(n_749),
.Y(n_879)
);

INVx1_ASAP7_75t_L g880 ( 
.A(n_742),
.Y(n_880)
);

NAND2xp5_ASAP7_75t_L g881 ( 
.A(n_753),
.B(n_251),
.Y(n_881)
);

INVx1_ASAP7_75t_L g882 ( 
.A(n_743),
.Y(n_882)
);

A2O1A1Ixp33_ASAP7_75t_L g883 ( 
.A1(n_709),
.A2(n_381),
.B(n_313),
.C(n_298),
.Y(n_883)
);

NOR3xp33_ASAP7_75t_L g884 ( 
.A(n_723),
.B(n_382),
.C(n_298),
.Y(n_884)
);

BUFx3_ASAP7_75t_L g885 ( 
.A(n_727),
.Y(n_885)
);

OAI22xp5_ASAP7_75t_L g886 ( 
.A1(n_733),
.A2(n_385),
.B1(n_360),
.B2(n_411),
.Y(n_886)
);

INVx1_ASAP7_75t_L g887 ( 
.A(n_735),
.Y(n_887)
);

AOI22xp5_ASAP7_75t_SL g888 ( 
.A1(n_659),
.A2(n_382),
.B1(n_249),
.B2(n_247),
.Y(n_888)
);

INVx2_ASAP7_75t_L g889 ( 
.A(n_677),
.Y(n_889)
);

INVx2_ASAP7_75t_SL g890 ( 
.A(n_753),
.Y(n_890)
);

INVx8_ASAP7_75t_L g891 ( 
.A(n_733),
.Y(n_891)
);

NAND2xp5_ASAP7_75t_L g892 ( 
.A(n_701),
.B(n_360),
.Y(n_892)
);

INVx1_ASAP7_75t_L g893 ( 
.A(n_735),
.Y(n_893)
);

AND2x4_ASAP7_75t_L g894 ( 
.A(n_727),
.B(n_362),
.Y(n_894)
);

NAND2xp5_ASAP7_75t_L g895 ( 
.A(n_726),
.B(n_363),
.Y(n_895)
);

INVx1_ASAP7_75t_L g896 ( 
.A(n_677),
.Y(n_896)
);

NAND2xp5_ASAP7_75t_L g897 ( 
.A(n_731),
.B(n_367),
.Y(n_897)
);

NAND2xp5_ASAP7_75t_L g898 ( 
.A(n_728),
.B(n_367),
.Y(n_898)
);

BUFx6f_ASAP7_75t_L g899 ( 
.A(n_750),
.Y(n_899)
);

NAND2xp5_ASAP7_75t_SL g900 ( 
.A(n_737),
.B(n_373),
.Y(n_900)
);

NAND2xp5_ASAP7_75t_L g901 ( 
.A(n_624),
.B(n_373),
.Y(n_901)
);

NAND2xp5_ASAP7_75t_L g902 ( 
.A(n_624),
.B(n_378),
.Y(n_902)
);

BUFx3_ASAP7_75t_L g903 ( 
.A(n_711),
.Y(n_903)
);

INVx2_ASAP7_75t_L g904 ( 
.A(n_741),
.Y(n_904)
);

INVx4_ASAP7_75t_L g905 ( 
.A(n_622),
.Y(n_905)
);

INVx1_ASAP7_75t_L g906 ( 
.A(n_747),
.Y(n_906)
);

INVx2_ASAP7_75t_L g907 ( 
.A(n_741),
.Y(n_907)
);

NOR2x1p5_ASAP7_75t_L g908 ( 
.A(n_665),
.B(n_249),
.Y(n_908)
);

NAND2xp5_ASAP7_75t_L g909 ( 
.A(n_624),
.B(n_385),
.Y(n_909)
);

INVx2_ASAP7_75t_L g910 ( 
.A(n_751),
.Y(n_910)
);

INVx1_ASAP7_75t_L g911 ( 
.A(n_747),
.Y(n_911)
);

NAND2xp33_ASAP7_75t_L g912 ( 
.A(n_644),
.B(n_387),
.Y(n_912)
);

NAND2xp5_ASAP7_75t_L g913 ( 
.A(n_627),
.B(n_387),
.Y(n_913)
);

INVx2_ASAP7_75t_SL g914 ( 
.A(n_733),
.Y(n_914)
);

O2A1O1Ixp5_ASAP7_75t_L g915 ( 
.A1(n_627),
.A2(n_489),
.B(n_344),
.C(n_380),
.Y(n_915)
);

INVx1_ASAP7_75t_L g916 ( 
.A(n_744),
.Y(n_916)
);

NAND2xp5_ASAP7_75t_L g917 ( 
.A(n_627),
.B(n_389),
.Y(n_917)
);

AOI22xp33_ASAP7_75t_L g918 ( 
.A1(n_674),
.A2(n_356),
.B1(n_374),
.B2(n_381),
.Y(n_918)
);

INVx2_ASAP7_75t_L g919 ( 
.A(n_748),
.Y(n_919)
);

AND2x4_ASAP7_75t_L g920 ( 
.A(n_734),
.B(n_389),
.Y(n_920)
);

NAND2xp5_ASAP7_75t_L g921 ( 
.A(n_650),
.B(n_392),
.Y(n_921)
);

BUFx6f_ASAP7_75t_L g922 ( 
.A(n_750),
.Y(n_922)
);

NAND2xp5_ASAP7_75t_SL g923 ( 
.A(n_752),
.B(n_392),
.Y(n_923)
);

NAND2xp5_ASAP7_75t_L g924 ( 
.A(n_650),
.B(n_394),
.Y(n_924)
);

AND2x6_ASAP7_75t_L g925 ( 
.A(n_772),
.B(n_758),
.Y(n_925)
);

HB1xp67_ASAP7_75t_L g926 ( 
.A(n_828),
.Y(n_926)
);

AND2x2_ASAP7_75t_L g927 ( 
.A(n_788),
.B(n_690),
.Y(n_927)
);

CKINVDCx5p33_ASAP7_75t_R g928 ( 
.A(n_783),
.Y(n_928)
);

AOI21xp5_ASAP7_75t_L g929 ( 
.A1(n_800),
.A2(n_668),
.B(n_760),
.Y(n_929)
);

AND2x2_ASAP7_75t_L g930 ( 
.A(n_790),
.B(n_690),
.Y(n_930)
);

OAI21xp33_ASAP7_75t_L g931 ( 
.A1(n_803),
.A2(n_693),
.B(n_647),
.Y(n_931)
);

NAND2xp5_ASAP7_75t_SL g932 ( 
.A(n_790),
.B(n_761),
.Y(n_932)
);

AOI21x1_ASAP7_75t_L g933 ( 
.A1(n_824),
.A2(n_655),
.B(n_652),
.Y(n_933)
);

NAND2xp5_ASAP7_75t_L g934 ( 
.A(n_890),
.B(n_650),
.Y(n_934)
);

AOI21xp5_ASAP7_75t_L g935 ( 
.A1(n_800),
.A2(n_760),
.B(n_661),
.Y(n_935)
);

OAI22xp5_ASAP7_75t_L g936 ( 
.A1(n_859),
.A2(n_740),
.B1(n_694),
.B2(n_746),
.Y(n_936)
);

NOR2xp33_ASAP7_75t_L g937 ( 
.A(n_867),
.B(n_654),
.Y(n_937)
);

NAND2xp5_ASAP7_75t_L g938 ( 
.A(n_782),
.B(n_827),
.Y(n_938)
);

BUFx6f_ASAP7_75t_L g939 ( 
.A(n_813),
.Y(n_939)
);

NAND2xp5_ASAP7_75t_SL g940 ( 
.A(n_850),
.B(n_665),
.Y(n_940)
);

NAND3xp33_ASAP7_75t_SL g941 ( 
.A(n_786),
.B(n_763),
.C(n_884),
.Y(n_941)
);

AOI21xp5_ASAP7_75t_L g942 ( 
.A1(n_832),
.A2(n_760),
.B(n_668),
.Y(n_942)
);

BUFx4f_ASAP7_75t_L g943 ( 
.A(n_852),
.Y(n_943)
);

AOI21xp5_ASAP7_75t_L g944 ( 
.A1(n_832),
.A2(n_707),
.B(n_661),
.Y(n_944)
);

NAND2xp5_ASAP7_75t_L g945 ( 
.A(n_775),
.B(n_660),
.Y(n_945)
);

AOI21xp5_ASAP7_75t_L g946 ( 
.A1(n_905),
.A2(n_707),
.B(n_661),
.Y(n_946)
);

INVx5_ASAP7_75t_L g947 ( 
.A(n_899),
.Y(n_947)
);

NOR2xp33_ASAP7_75t_L g948 ( 
.A(n_768),
.B(n_688),
.Y(n_948)
);

NAND2xp33_ASAP7_75t_L g949 ( 
.A(n_813),
.B(n_871),
.Y(n_949)
);

O2A1O1Ixp33_ASAP7_75t_L g950 ( 
.A1(n_769),
.A2(n_730),
.B(n_669),
.C(n_672),
.Y(n_950)
);

OR2x6_ASAP7_75t_SL g951 ( 
.A(n_845),
.B(n_374),
.Y(n_951)
);

INVx1_ASAP7_75t_L g952 ( 
.A(n_808),
.Y(n_952)
);

INVx2_ASAP7_75t_L g953 ( 
.A(n_780),
.Y(n_953)
);

NAND2xp5_ASAP7_75t_L g954 ( 
.A(n_827),
.B(n_660),
.Y(n_954)
);

NAND2xp5_ASAP7_75t_L g955 ( 
.A(n_840),
.B(n_660),
.Y(n_955)
);

AOI21xp5_ASAP7_75t_L g956 ( 
.A1(n_905),
.A2(n_668),
.B(n_707),
.Y(n_956)
);

AOI21xp5_ASAP7_75t_L g957 ( 
.A1(n_826),
.A2(n_616),
.B(n_680),
.Y(n_957)
);

BUFx6f_ASAP7_75t_L g958 ( 
.A(n_813),
.Y(n_958)
);

NAND2xp5_ASAP7_75t_L g959 ( 
.A(n_840),
.B(n_666),
.Y(n_959)
);

OAI22xp5_ASAP7_75t_L g960 ( 
.A1(n_859),
.A2(n_745),
.B1(n_705),
.B2(n_684),
.Y(n_960)
);

AOI21xp5_ASAP7_75t_L g961 ( 
.A1(n_826),
.A2(n_616),
.B(n_680),
.Y(n_961)
);

AOI22xp33_ASAP7_75t_SL g962 ( 
.A1(n_803),
.A2(n_749),
.B1(n_489),
.B2(n_738),
.Y(n_962)
);

OAI22xp5_ASAP7_75t_L g963 ( 
.A1(n_873),
.A2(n_715),
.B1(n_400),
.B2(n_401),
.Y(n_963)
);

NAND2xp5_ASAP7_75t_L g964 ( 
.A(n_842),
.B(n_666),
.Y(n_964)
);

AOI21xp5_ASAP7_75t_L g965 ( 
.A1(n_795),
.A2(n_616),
.B(n_680),
.Y(n_965)
);

OAI21xp5_ASAP7_75t_L g966 ( 
.A1(n_824),
.A2(n_666),
.B(n_692),
.Y(n_966)
);

AOI21xp5_ASAP7_75t_L g967 ( 
.A1(n_830),
.A2(n_722),
.B(n_622),
.Y(n_967)
);

AOI22xp5_ASAP7_75t_L g968 ( 
.A1(n_842),
.A2(n_759),
.B1(n_674),
.B2(n_644),
.Y(n_968)
);

OAI21xp5_ASAP7_75t_L g969 ( 
.A1(n_769),
.A2(n_692),
.B(n_644),
.Y(n_969)
);

INVx3_ASAP7_75t_L g970 ( 
.A(n_846),
.Y(n_970)
);

AOI21xp5_ASAP7_75t_L g971 ( 
.A1(n_811),
.A2(n_622),
.B(n_680),
.Y(n_971)
);

AOI21xp5_ASAP7_75t_L g972 ( 
.A1(n_811),
.A2(n_622),
.B(n_680),
.Y(n_972)
);

NAND2xp5_ASAP7_75t_L g973 ( 
.A(n_821),
.B(n_756),
.Y(n_973)
);

OAI21xp5_ASAP7_75t_L g974 ( 
.A1(n_766),
.A2(n_644),
.B(n_674),
.Y(n_974)
);

OAI21xp5_ASAP7_75t_L g975 ( 
.A1(n_766),
.A2(n_644),
.B(n_674),
.Y(n_975)
);

INVx4_ASAP7_75t_L g976 ( 
.A(n_813),
.Y(n_976)
);

BUFx6f_ASAP7_75t_L g977 ( 
.A(n_871),
.Y(n_977)
);

O2A1O1Ixp33_ASAP7_75t_L g978 ( 
.A1(n_849),
.A2(n_883),
.B(n_865),
.C(n_767),
.Y(n_978)
);

A2O1A1Ixp33_ASAP7_75t_L g979 ( 
.A1(n_773),
.A2(n_411),
.B(n_394),
.C(n_398),
.Y(n_979)
);

AOI21xp5_ASAP7_75t_L g980 ( 
.A1(n_776),
.A2(n_722),
.B(n_536),
.Y(n_980)
);

NOR2xp67_ASAP7_75t_L g981 ( 
.A(n_774),
.B(n_398),
.Y(n_981)
);

OAI21x1_ASAP7_75t_L g982 ( 
.A1(n_904),
.A2(n_674),
.B(n_722),
.Y(n_982)
);

AOI21xp5_ASAP7_75t_L g983 ( 
.A1(n_776),
.A2(n_722),
.B(n_536),
.Y(n_983)
);

AND2x2_ASAP7_75t_L g984 ( 
.A(n_875),
.B(n_738),
.Y(n_984)
);

AOI21xp5_ASAP7_75t_L g985 ( 
.A1(n_853),
.A2(n_536),
.B(n_686),
.Y(n_985)
);

AOI21xp5_ASAP7_75t_L g986 ( 
.A1(n_853),
.A2(n_536),
.B(n_686),
.Y(n_986)
);

BUFx3_ASAP7_75t_L g987 ( 
.A(n_862),
.Y(n_987)
);

AOI21xp5_ASAP7_75t_L g988 ( 
.A1(n_901),
.A2(n_686),
.B(n_697),
.Y(n_988)
);

AO21x2_ASAP7_75t_L g989 ( 
.A1(n_829),
.A2(n_725),
.B(n_674),
.Y(n_989)
);

NOR2xp33_ASAP7_75t_L g990 ( 
.A(n_771),
.B(n_755),
.Y(n_990)
);

BUFx12f_ASAP7_75t_L g991 ( 
.A(n_862),
.Y(n_991)
);

O2A1O1Ixp33_ASAP7_75t_L g992 ( 
.A1(n_883),
.A2(n_755),
.B(n_380),
.C(n_399),
.Y(n_992)
);

NOR2xp33_ASAP7_75t_L g993 ( 
.A(n_785),
.B(n_738),
.Y(n_993)
);

OAI21xp5_ASAP7_75t_L g994 ( 
.A1(n_843),
.A2(n_725),
.B(n_686),
.Y(n_994)
);

AND2x2_ASAP7_75t_L g995 ( 
.A(n_844),
.B(n_400),
.Y(n_995)
);

NOR2xp33_ASAP7_75t_L g996 ( 
.A(n_839),
.B(n_401),
.Y(n_996)
);

INVx4_ASAP7_75t_L g997 ( 
.A(n_871),
.Y(n_997)
);

AO21x1_ASAP7_75t_L g998 ( 
.A1(n_829),
.A2(n_725),
.B(n_399),
.Y(n_998)
);

AOI21xp5_ASAP7_75t_L g999 ( 
.A1(n_902),
.A2(n_686),
.B(n_725),
.Y(n_999)
);

AOI21xp5_ASAP7_75t_L g1000 ( 
.A1(n_909),
.A2(n_725),
.B(n_409),
.Y(n_1000)
);

NAND2xp5_ASAP7_75t_SL g1001 ( 
.A(n_791),
.B(n_399),
.Y(n_1001)
);

BUFx3_ASAP7_75t_L g1002 ( 
.A(n_879),
.Y(n_1002)
);

NAND2xp5_ASAP7_75t_L g1003 ( 
.A(n_864),
.B(n_725),
.Y(n_1003)
);

NOR2xp33_ASAP7_75t_L g1004 ( 
.A(n_773),
.B(n_409),
.Y(n_1004)
);

AOI21xp5_ASAP7_75t_L g1005 ( 
.A1(n_913),
.A2(n_406),
.B(n_402),
.Y(n_1005)
);

NAND2xp5_ASAP7_75t_L g1006 ( 
.A(n_876),
.B(n_402),
.Y(n_1006)
);

AOI21x1_ASAP7_75t_L g1007 ( 
.A1(n_856),
.A2(n_380),
.B(n_208),
.Y(n_1007)
);

OAI21xp5_ASAP7_75t_L g1008 ( 
.A1(n_831),
.A2(n_206),
.B(n_200),
.Y(n_1008)
);

NAND2xp5_ASAP7_75t_L g1009 ( 
.A(n_784),
.B(n_16),
.Y(n_1009)
);

NAND2xp5_ASAP7_75t_L g1010 ( 
.A(n_784),
.B(n_18),
.Y(n_1010)
);

NAND2xp5_ASAP7_75t_L g1011 ( 
.A(n_880),
.B(n_19),
.Y(n_1011)
);

INVx1_ASAP7_75t_L g1012 ( 
.A(n_837),
.Y(n_1012)
);

NOR2xp33_ASAP7_75t_L g1013 ( 
.A(n_878),
.B(n_19),
.Y(n_1013)
);

BUFx12f_ASAP7_75t_L g1014 ( 
.A(n_879),
.Y(n_1014)
);

OAI22xp5_ASAP7_75t_L g1015 ( 
.A1(n_873),
.A2(n_20),
.B1(n_22),
.B2(n_23),
.Y(n_1015)
);

NAND2xp5_ASAP7_75t_L g1016 ( 
.A(n_764),
.B(n_22),
.Y(n_1016)
);

NAND2xp5_ASAP7_75t_SL g1017 ( 
.A(n_855),
.B(n_197),
.Y(n_1017)
);

AOI21xp5_ASAP7_75t_L g1018 ( 
.A1(n_917),
.A2(n_186),
.B(n_184),
.Y(n_1018)
);

NAND2xp5_ASAP7_75t_L g1019 ( 
.A(n_779),
.B(n_23),
.Y(n_1019)
);

NAND2x1p5_ASAP7_75t_L g1020 ( 
.A(n_846),
.B(n_182),
.Y(n_1020)
);

NAND2xp5_ASAP7_75t_L g1021 ( 
.A(n_837),
.B(n_175),
.Y(n_1021)
);

AOI22xp5_ASAP7_75t_L g1022 ( 
.A1(n_799),
.A2(n_858),
.B1(n_872),
.B2(n_868),
.Y(n_1022)
);

NAND2xp5_ASAP7_75t_L g1023 ( 
.A(n_863),
.B(n_116),
.Y(n_1023)
);

NAND2xp5_ASAP7_75t_L g1024 ( 
.A(n_863),
.B(n_159),
.Y(n_1024)
);

NOR2xp33_ASAP7_75t_SL g1025 ( 
.A(n_903),
.B(n_157),
.Y(n_1025)
);

AND2x2_ASAP7_75t_L g1026 ( 
.A(n_854),
.B(n_26),
.Y(n_1026)
);

OAI21xp5_ASAP7_75t_L g1027 ( 
.A1(n_780),
.A2(n_154),
.B(n_145),
.Y(n_1027)
);

NAND2xp5_ASAP7_75t_SL g1028 ( 
.A(n_820),
.B(n_138),
.Y(n_1028)
);

NAND2xp5_ASAP7_75t_L g1029 ( 
.A(n_792),
.B(n_28),
.Y(n_1029)
);

AND2x4_ASAP7_75t_L g1030 ( 
.A(n_777),
.B(n_134),
.Y(n_1030)
);

AOI21xp5_ASAP7_75t_L g1031 ( 
.A1(n_921),
.A2(n_133),
.B(n_129),
.Y(n_1031)
);

INVx1_ASAP7_75t_L g1032 ( 
.A(n_887),
.Y(n_1032)
);

NAND2xp5_ASAP7_75t_L g1033 ( 
.A(n_893),
.B(n_101),
.Y(n_1033)
);

NAND2xp5_ASAP7_75t_SL g1034 ( 
.A(n_861),
.B(n_98),
.Y(n_1034)
);

INVx1_ASAP7_75t_L g1035 ( 
.A(n_896),
.Y(n_1035)
);

NAND2xp5_ASAP7_75t_L g1036 ( 
.A(n_794),
.B(n_40),
.Y(n_1036)
);

NAND2xp5_ASAP7_75t_L g1037 ( 
.A(n_892),
.B(n_40),
.Y(n_1037)
);

NAND2xp5_ASAP7_75t_L g1038 ( 
.A(n_895),
.B(n_41),
.Y(n_1038)
);

AOI21xp5_ASAP7_75t_L g1039 ( 
.A1(n_924),
.A2(n_97),
.B(n_92),
.Y(n_1039)
);

AOI21xp5_ASAP7_75t_L g1040 ( 
.A1(n_835),
.A2(n_91),
.B(n_74),
.Y(n_1040)
);

NOR2xp33_ASAP7_75t_L g1041 ( 
.A(n_878),
.B(n_41),
.Y(n_1041)
);

AOI221xp5_ASAP7_75t_L g1042 ( 
.A1(n_834),
.A2(n_43),
.B1(n_46),
.B2(n_48),
.C(n_49),
.Y(n_1042)
);

AOI21xp5_ASAP7_75t_L g1043 ( 
.A1(n_898),
.A2(n_50),
.B(n_51),
.Y(n_1043)
);

OAI22xp5_ASAP7_75t_L g1044 ( 
.A1(n_838),
.A2(n_53),
.B1(n_54),
.B2(n_55),
.Y(n_1044)
);

NAND2xp5_ASAP7_75t_L g1045 ( 
.A(n_881),
.B(n_869),
.Y(n_1045)
);

AOI21xp5_ASAP7_75t_L g1046 ( 
.A1(n_789),
.A2(n_55),
.B(n_56),
.Y(n_1046)
);

AND2x2_ASAP7_75t_L g1047 ( 
.A(n_854),
.B(n_57),
.Y(n_1047)
);

NAND2xp5_ASAP7_75t_L g1048 ( 
.A(n_870),
.B(n_61),
.Y(n_1048)
);

INVx3_ASAP7_75t_L g1049 ( 
.A(n_899),
.Y(n_1049)
);

INVx1_ASAP7_75t_L g1050 ( 
.A(n_906),
.Y(n_1050)
);

AND2x2_ASAP7_75t_L g1051 ( 
.A(n_852),
.B(n_66),
.Y(n_1051)
);

NAND2xp5_ASAP7_75t_L g1052 ( 
.A(n_781),
.B(n_66),
.Y(n_1052)
);

INVx3_ASAP7_75t_L g1053 ( 
.A(n_899),
.Y(n_1053)
);

NAND2xp5_ASAP7_75t_L g1054 ( 
.A(n_882),
.B(n_897),
.Y(n_1054)
);

O2A1O1Ixp5_ASAP7_75t_L g1055 ( 
.A1(n_900),
.A2(n_797),
.B(n_793),
.C(n_841),
.Y(n_1055)
);

AND2x2_ASAP7_75t_L g1056 ( 
.A(n_852),
.B(n_894),
.Y(n_1056)
);

NAND2xp5_ASAP7_75t_L g1057 ( 
.A(n_806),
.B(n_807),
.Y(n_1057)
);

OAI22xp5_ASAP7_75t_L g1058 ( 
.A1(n_838),
.A2(n_918),
.B1(n_770),
.B2(n_834),
.Y(n_1058)
);

INVx2_ASAP7_75t_L g1059 ( 
.A(n_806),
.Y(n_1059)
);

BUFx4f_ASAP7_75t_L g1060 ( 
.A(n_891),
.Y(n_1060)
);

NOR2x1_ASAP7_75t_L g1061 ( 
.A(n_762),
.B(n_777),
.Y(n_1061)
);

BUFx6f_ASAP7_75t_L g1062 ( 
.A(n_871),
.Y(n_1062)
);

NAND2xp5_ASAP7_75t_L g1063 ( 
.A(n_796),
.B(n_818),
.Y(n_1063)
);

OAI21xp33_ASAP7_75t_L g1064 ( 
.A1(n_809),
.A2(n_770),
.B(n_857),
.Y(n_1064)
);

AND2x2_ASAP7_75t_L g1065 ( 
.A(n_894),
.B(n_920),
.Y(n_1065)
);

BUFx6f_ASAP7_75t_L g1066 ( 
.A(n_899),
.Y(n_1066)
);

OAI21xp5_ASAP7_75t_L g1067 ( 
.A1(n_807),
.A2(n_814),
.B(n_802),
.Y(n_1067)
);

INVx1_ASAP7_75t_L g1068 ( 
.A(n_911),
.Y(n_1068)
);

BUFx6f_ASAP7_75t_L g1069 ( 
.A(n_922),
.Y(n_1069)
);

NAND3xp33_ASAP7_75t_L g1070 ( 
.A(n_866),
.B(n_798),
.C(n_787),
.Y(n_1070)
);

NAND2xp5_ASAP7_75t_L g1071 ( 
.A(n_805),
.B(n_819),
.Y(n_1071)
);

NAND2xp5_ASAP7_75t_SL g1072 ( 
.A(n_920),
.B(n_914),
.Y(n_1072)
);

OAI21x1_ASAP7_75t_L g1073 ( 
.A1(n_904),
.A2(n_907),
.B(n_910),
.Y(n_1073)
);

INVx1_ASAP7_75t_L g1074 ( 
.A(n_823),
.Y(n_1074)
);

INVx1_ASAP7_75t_L g1075 ( 
.A(n_874),
.Y(n_1075)
);

AND2x2_ASAP7_75t_L g1076 ( 
.A(n_866),
.B(n_783),
.Y(n_1076)
);

NAND2xp33_ASAP7_75t_L g1077 ( 
.A(n_922),
.B(n_891),
.Y(n_1077)
);

NOR2xp33_ASAP7_75t_L g1078 ( 
.A(n_778),
.B(n_886),
.Y(n_1078)
);

AOI21xp5_ASAP7_75t_L g1079 ( 
.A1(n_889),
.A2(n_922),
.B(n_900),
.Y(n_1079)
);

INVx1_ASAP7_75t_L g1080 ( 
.A(n_919),
.Y(n_1080)
);

NAND2xp5_ASAP7_75t_SL g1081 ( 
.A(n_860),
.B(n_885),
.Y(n_1081)
);

A2O1A1Ixp33_ASAP7_75t_L g1082 ( 
.A1(n_918),
.A2(n_817),
.B(n_815),
.C(n_916),
.Y(n_1082)
);

NAND2xp5_ASAP7_75t_L g1083 ( 
.A(n_877),
.B(n_860),
.Y(n_1083)
);

NAND2xp5_ASAP7_75t_L g1084 ( 
.A(n_885),
.B(n_833),
.Y(n_1084)
);

INVxp67_ASAP7_75t_L g1085 ( 
.A(n_848),
.Y(n_1085)
);

NAND2xp5_ASAP7_75t_SL g1086 ( 
.A(n_922),
.B(n_891),
.Y(n_1086)
);

INVx1_ASAP7_75t_L g1087 ( 
.A(n_919),
.Y(n_1087)
);

AOI221xp5_ASAP7_75t_L g1088 ( 
.A1(n_851),
.A2(n_923),
.B1(n_915),
.B2(n_816),
.C(n_810),
.Y(n_1088)
);

OAI21xp5_ASAP7_75t_L g1089 ( 
.A1(n_907),
.A2(n_810),
.B(n_816),
.Y(n_1089)
);

INVx2_ASAP7_75t_L g1090 ( 
.A(n_765),
.Y(n_1090)
);

INVx2_ASAP7_75t_L g1091 ( 
.A(n_812),
.Y(n_1091)
);

NAND2xp5_ASAP7_75t_L g1092 ( 
.A(n_923),
.B(n_801),
.Y(n_1092)
);

NAND2xp5_ASAP7_75t_L g1093 ( 
.A(n_847),
.B(n_822),
.Y(n_1093)
);

A2O1A1Ixp33_ASAP7_75t_L g1094 ( 
.A1(n_836),
.A2(n_825),
.B(n_912),
.C(n_888),
.Y(n_1094)
);

INVx3_ASAP7_75t_L g1095 ( 
.A(n_903),
.Y(n_1095)
);

OA22x2_ASAP7_75t_L g1096 ( 
.A1(n_908),
.A2(n_850),
.B1(n_620),
.B2(n_844),
.Y(n_1096)
);

AOI22xp5_ASAP7_75t_L g1097 ( 
.A1(n_804),
.A2(n_790),
.B1(n_859),
.B2(n_664),
.Y(n_1097)
);

NOR2xp33_ASAP7_75t_L g1098 ( 
.A(n_867),
.B(n_790),
.Y(n_1098)
);

AOI21xp5_ASAP7_75t_L g1099 ( 
.A1(n_800),
.A2(n_702),
.B(n_832),
.Y(n_1099)
);

BUFx4f_ASAP7_75t_L g1100 ( 
.A(n_852),
.Y(n_1100)
);

NAND2xp5_ASAP7_75t_SL g1101 ( 
.A(n_790),
.B(n_850),
.Y(n_1101)
);

NOR2xp33_ASAP7_75t_SL g1102 ( 
.A(n_862),
.B(n_659),
.Y(n_1102)
);

AOI21xp5_ASAP7_75t_L g1103 ( 
.A1(n_1099),
.A2(n_1071),
.B(n_1063),
.Y(n_1103)
);

NAND2xp5_ASAP7_75t_L g1104 ( 
.A(n_938),
.B(n_1098),
.Y(n_1104)
);

NOR2xp33_ASAP7_75t_L g1105 ( 
.A(n_930),
.B(n_937),
.Y(n_1105)
);

NAND2xp5_ASAP7_75t_L g1106 ( 
.A(n_1045),
.B(n_1101),
.Y(n_1106)
);

OR2x2_ASAP7_75t_L g1107 ( 
.A(n_927),
.B(n_926),
.Y(n_1107)
);

AOI21xp5_ASAP7_75t_L g1108 ( 
.A1(n_949),
.A2(n_972),
.B(n_971),
.Y(n_1108)
);

NAND2xp5_ASAP7_75t_SL g1109 ( 
.A(n_1097),
.B(n_984),
.Y(n_1109)
);

NAND2xp5_ASAP7_75t_L g1110 ( 
.A(n_1054),
.B(n_1004),
.Y(n_1110)
);

OAI21x1_ASAP7_75t_L g1111 ( 
.A1(n_982),
.A2(n_1073),
.B(n_961),
.Y(n_1111)
);

AOI21x1_ASAP7_75t_SL g1112 ( 
.A1(n_1009),
.A2(n_1010),
.B(n_1048),
.Y(n_1112)
);

O2A1O1Ixp33_ASAP7_75t_L g1113 ( 
.A1(n_1013),
.A2(n_1041),
.B(n_1058),
.C(n_1015),
.Y(n_1113)
);

NOR2x1_ASAP7_75t_SL g1114 ( 
.A(n_947),
.B(n_1066),
.Y(n_1114)
);

AOI21xp5_ASAP7_75t_SL g1115 ( 
.A1(n_1058),
.A2(n_1008),
.B(n_1027),
.Y(n_1115)
);

AOI21xp5_ASAP7_75t_L g1116 ( 
.A1(n_954),
.A2(n_959),
.B(n_955),
.Y(n_1116)
);

OAI22x1_ASAP7_75t_L g1117 ( 
.A1(n_1078),
.A2(n_940),
.B1(n_932),
.B2(n_1072),
.Y(n_1117)
);

AOI21xp33_ASAP7_75t_L g1118 ( 
.A1(n_978),
.A2(n_1096),
.B(n_1070),
.Y(n_1118)
);

OA22x2_ASAP7_75t_L g1119 ( 
.A1(n_931),
.A2(n_963),
.B1(n_1015),
.B2(n_1044),
.Y(n_1119)
);

OAI21x1_ASAP7_75t_L g1120 ( 
.A1(n_957),
.A2(n_1079),
.B(n_965),
.Y(n_1120)
);

OAI21x1_ASAP7_75t_L g1121 ( 
.A1(n_946),
.A2(n_956),
.B(n_966),
.Y(n_1121)
);

OAI21xp5_ASAP7_75t_L g1122 ( 
.A1(n_1082),
.A2(n_1055),
.B(n_969),
.Y(n_1122)
);

INVx2_ASAP7_75t_L g1123 ( 
.A(n_953),
.Y(n_1123)
);

OAI21x1_ASAP7_75t_SL g1124 ( 
.A1(n_1008),
.A2(n_1027),
.B(n_969),
.Y(n_1124)
);

INVx1_ASAP7_75t_L g1125 ( 
.A(n_1080),
.Y(n_1125)
);

OAI21x1_ASAP7_75t_L g1126 ( 
.A1(n_966),
.A2(n_967),
.B(n_935),
.Y(n_1126)
);

OAI22xp5_ASAP7_75t_L g1127 ( 
.A1(n_936),
.A2(n_1047),
.B1(n_1026),
.B2(n_1096),
.Y(n_1127)
);

OAI21x1_ASAP7_75t_L g1128 ( 
.A1(n_929),
.A2(n_944),
.B(n_942),
.Y(n_1128)
);

NAND2xp5_ASAP7_75t_L g1129 ( 
.A(n_1050),
.B(n_1068),
.Y(n_1129)
);

NOR2x1_ASAP7_75t_SL g1130 ( 
.A(n_947),
.B(n_1066),
.Y(n_1130)
);

AO31x2_ASAP7_75t_L g1131 ( 
.A1(n_998),
.A2(n_1094),
.A3(n_964),
.B(n_1033),
.Y(n_1131)
);

INVx4_ASAP7_75t_L g1132 ( 
.A(n_939),
.Y(n_1132)
);

AOI21xp5_ASAP7_75t_L g1133 ( 
.A1(n_947),
.A2(n_1067),
.B(n_1084),
.Y(n_1133)
);

O2A1O1Ixp5_ASAP7_75t_L g1134 ( 
.A1(n_1037),
.A2(n_1038),
.B(n_988),
.C(n_1052),
.Y(n_1134)
);

NOR2xp33_ASAP7_75t_L g1135 ( 
.A(n_948),
.B(n_993),
.Y(n_1135)
);

NAND3xp33_ASAP7_75t_L g1136 ( 
.A(n_990),
.B(n_963),
.C(n_996),
.Y(n_1136)
);

INVx1_ASAP7_75t_L g1137 ( 
.A(n_1087),
.Y(n_1137)
);

INVx3_ASAP7_75t_L g1138 ( 
.A(n_1066),
.Y(n_1138)
);

BUFx6f_ASAP7_75t_L g1139 ( 
.A(n_939),
.Y(n_1139)
);

NAND2xp5_ASAP7_75t_L g1140 ( 
.A(n_1083),
.B(n_1092),
.Y(n_1140)
);

INVx1_ASAP7_75t_L g1141 ( 
.A(n_952),
.Y(n_1141)
);

BUFx6f_ASAP7_75t_L g1142 ( 
.A(n_939),
.Y(n_1142)
);

AND2x2_ASAP7_75t_L g1143 ( 
.A(n_995),
.B(n_1065),
.Y(n_1143)
);

OAI21xp5_ASAP7_75t_L g1144 ( 
.A1(n_1067),
.A2(n_1057),
.B(n_1089),
.Y(n_1144)
);

CKINVDCx5p33_ASAP7_75t_R g1145 ( 
.A(n_928),
.Y(n_1145)
);

OAI21x1_ASAP7_75t_L g1146 ( 
.A1(n_1089),
.A2(n_999),
.B(n_1024),
.Y(n_1146)
);

BUFx6f_ASAP7_75t_L g1147 ( 
.A(n_958),
.Y(n_1147)
);

AND2x4_ASAP7_75t_L g1148 ( 
.A(n_1061),
.B(n_1081),
.Y(n_1148)
);

AOI21x1_ASAP7_75t_L g1149 ( 
.A1(n_1021),
.A2(n_1023),
.B(n_1024),
.Y(n_1149)
);

CKINVDCx5p33_ASAP7_75t_R g1150 ( 
.A(n_991),
.Y(n_1150)
);

NOR2xp33_ASAP7_75t_L g1151 ( 
.A(n_941),
.B(n_1076),
.Y(n_1151)
);

O2A1O1Ixp5_ASAP7_75t_L g1152 ( 
.A1(n_994),
.A2(n_1034),
.B(n_1016),
.C(n_1028),
.Y(n_1152)
);

AO31x2_ASAP7_75t_L g1153 ( 
.A1(n_1033),
.A2(n_1021),
.A3(n_1023),
.B(n_979),
.Y(n_1153)
);

A2O1A1Ixp33_ASAP7_75t_L g1154 ( 
.A1(n_1064),
.A2(n_950),
.B(n_1088),
.C(n_1022),
.Y(n_1154)
);

OAI21xp5_ASAP7_75t_L g1155 ( 
.A1(n_945),
.A2(n_936),
.B(n_1012),
.Y(n_1155)
);

BUFx6f_ASAP7_75t_SL g1156 ( 
.A(n_987),
.Y(n_1156)
);

OAI21x1_ASAP7_75t_L g1157 ( 
.A1(n_985),
.A2(n_986),
.B(n_994),
.Y(n_1157)
);

AO31x2_ASAP7_75t_L g1158 ( 
.A1(n_960),
.A2(n_1029),
.A3(n_1036),
.B(n_1019),
.Y(n_1158)
);

NAND2xp5_ASAP7_75t_SL g1159 ( 
.A(n_960),
.B(n_1030),
.Y(n_1159)
);

BUFx6f_ASAP7_75t_L g1160 ( 
.A(n_958),
.Y(n_1160)
);

OAI21xp33_ASAP7_75t_L g1161 ( 
.A1(n_1006),
.A2(n_1005),
.B(n_962),
.Y(n_1161)
);

AOI21x1_ASAP7_75t_SL g1162 ( 
.A1(n_1093),
.A2(n_1011),
.B(n_1003),
.Y(n_1162)
);

AOI211x1_ASAP7_75t_L g1163 ( 
.A1(n_1044),
.A2(n_1043),
.B(n_933),
.C(n_1046),
.Y(n_1163)
);

OAI21x1_ASAP7_75t_L g1164 ( 
.A1(n_973),
.A2(n_983),
.B(n_980),
.Y(n_1164)
);

INVx1_ASAP7_75t_L g1165 ( 
.A(n_1059),
.Y(n_1165)
);

AO31x2_ASAP7_75t_L g1166 ( 
.A1(n_1000),
.A2(n_1018),
.A3(n_1031),
.B(n_1039),
.Y(n_1166)
);

BUFx2_ASAP7_75t_L g1167 ( 
.A(n_1056),
.Y(n_1167)
);

OAI22xp5_ASAP7_75t_L g1168 ( 
.A1(n_1030),
.A2(n_1042),
.B1(n_1100),
.B2(n_943),
.Y(n_1168)
);

AND3x4_ASAP7_75t_L g1169 ( 
.A(n_1002),
.B(n_981),
.C(n_951),
.Y(n_1169)
);

A2O1A1Ixp33_ASAP7_75t_L g1170 ( 
.A1(n_992),
.A2(n_1032),
.B(n_968),
.C(n_1035),
.Y(n_1170)
);

NAND2xp5_ASAP7_75t_L g1171 ( 
.A(n_970),
.B(n_925),
.Y(n_1171)
);

AOI21xp5_ASAP7_75t_L g1172 ( 
.A1(n_947),
.A2(n_970),
.B(n_1077),
.Y(n_1172)
);

OR2x2_ASAP7_75t_L g1173 ( 
.A(n_1095),
.B(n_1085),
.Y(n_1173)
);

NAND2xp5_ASAP7_75t_L g1174 ( 
.A(n_925),
.B(n_1090),
.Y(n_1174)
);

OAI21xp5_ASAP7_75t_L g1175 ( 
.A1(n_974),
.A2(n_975),
.B(n_1075),
.Y(n_1175)
);

OAI21xp33_ASAP7_75t_L g1176 ( 
.A1(n_1102),
.A2(n_1051),
.B(n_1001),
.Y(n_1176)
);

OAI21xp5_ASAP7_75t_L g1177 ( 
.A1(n_974),
.A2(n_975),
.B(n_1074),
.Y(n_1177)
);

BUFx6f_ASAP7_75t_L g1178 ( 
.A(n_958),
.Y(n_1178)
);

AOI21x1_ASAP7_75t_L g1179 ( 
.A1(n_934),
.A2(n_1007),
.B(n_1017),
.Y(n_1179)
);

CKINVDCx5p33_ASAP7_75t_R g1180 ( 
.A(n_1014),
.Y(n_1180)
);

NAND2xp5_ASAP7_75t_L g1181 ( 
.A(n_925),
.B(n_1091),
.Y(n_1181)
);

NAND2x1p5_ASAP7_75t_L g1182 ( 
.A(n_976),
.B(n_997),
.Y(n_1182)
);

OAI21x1_ASAP7_75t_SL g1183 ( 
.A1(n_1040),
.A2(n_976),
.B(n_997),
.Y(n_1183)
);

AOI21xp5_ASAP7_75t_L g1184 ( 
.A1(n_1049),
.A2(n_1053),
.B(n_1086),
.Y(n_1184)
);

NAND2xp5_ASAP7_75t_L g1185 ( 
.A(n_925),
.B(n_977),
.Y(n_1185)
);

OAI21x1_ASAP7_75t_L g1186 ( 
.A1(n_1020),
.A2(n_1095),
.B(n_989),
.Y(n_1186)
);

AOI21xp5_ASAP7_75t_L g1187 ( 
.A1(n_1069),
.A2(n_1062),
.B(n_977),
.Y(n_1187)
);

OAI21x1_ASAP7_75t_L g1188 ( 
.A1(n_1020),
.A2(n_989),
.B(n_925),
.Y(n_1188)
);

HB1xp67_ASAP7_75t_L g1189 ( 
.A(n_977),
.Y(n_1189)
);

OAI22xp5_ASAP7_75t_L g1190 ( 
.A1(n_943),
.A2(n_1100),
.B1(n_1060),
.B2(n_1062),
.Y(n_1190)
);

NAND2xp5_ASAP7_75t_L g1191 ( 
.A(n_1069),
.B(n_1025),
.Y(n_1191)
);

AOI21xp33_ASAP7_75t_L g1192 ( 
.A1(n_1069),
.A2(n_1060),
.B(n_1004),
.Y(n_1192)
);

AOI21x1_ASAP7_75t_L g1193 ( 
.A1(n_954),
.A2(n_959),
.B(n_955),
.Y(n_1193)
);

OAI21x1_ASAP7_75t_L g1194 ( 
.A1(n_982),
.A2(n_1073),
.B(n_961),
.Y(n_1194)
);

NAND2xp5_ASAP7_75t_L g1195 ( 
.A(n_938),
.B(n_1098),
.Y(n_1195)
);

NAND2xp5_ASAP7_75t_L g1196 ( 
.A(n_938),
.B(n_1098),
.Y(n_1196)
);

OAI21xp5_ASAP7_75t_L g1197 ( 
.A1(n_978),
.A2(n_1101),
.B(n_1082),
.Y(n_1197)
);

OAI21xp5_ASAP7_75t_L g1198 ( 
.A1(n_978),
.A2(n_1101),
.B(n_1082),
.Y(n_1198)
);

INVx2_ASAP7_75t_L g1199 ( 
.A(n_953),
.Y(n_1199)
);

OAI21x1_ASAP7_75t_SL g1200 ( 
.A1(n_1008),
.A2(n_1027),
.B(n_969),
.Y(n_1200)
);

AOI21xp5_ASAP7_75t_L g1201 ( 
.A1(n_1099),
.A2(n_702),
.B(n_800),
.Y(n_1201)
);

INVx6_ASAP7_75t_L g1202 ( 
.A(n_939),
.Y(n_1202)
);

OAI21xp5_ASAP7_75t_L g1203 ( 
.A1(n_978),
.A2(n_1101),
.B(n_1082),
.Y(n_1203)
);

AND2x6_ASAP7_75t_L g1204 ( 
.A(n_1030),
.B(n_1065),
.Y(n_1204)
);

AOI221xp5_ASAP7_75t_SL g1205 ( 
.A1(n_1058),
.A2(n_769),
.B1(n_1041),
.B2(n_1013),
.C(n_883),
.Y(n_1205)
);

OAI21xp5_ASAP7_75t_L g1206 ( 
.A1(n_978),
.A2(n_1101),
.B(n_1082),
.Y(n_1206)
);

INVx1_ASAP7_75t_L g1207 ( 
.A(n_1080),
.Y(n_1207)
);

AOI21xp33_ASAP7_75t_L g1208 ( 
.A1(n_1004),
.A2(n_938),
.B(n_1013),
.Y(n_1208)
);

INVx1_ASAP7_75t_L g1209 ( 
.A(n_1080),
.Y(n_1209)
);

INVx2_ASAP7_75t_L g1210 ( 
.A(n_953),
.Y(n_1210)
);

NAND2xp5_ASAP7_75t_L g1211 ( 
.A(n_938),
.B(n_1098),
.Y(n_1211)
);

HB1xp67_ASAP7_75t_L g1212 ( 
.A(n_926),
.Y(n_1212)
);

NAND2xp5_ASAP7_75t_SL g1213 ( 
.A(n_937),
.B(n_763),
.Y(n_1213)
);

OAI21x1_ASAP7_75t_L g1214 ( 
.A1(n_982),
.A2(n_1073),
.B(n_961),
.Y(n_1214)
);

CKINVDCx5p33_ASAP7_75t_R g1215 ( 
.A(n_928),
.Y(n_1215)
);

BUFx2_ASAP7_75t_L g1216 ( 
.A(n_926),
.Y(n_1216)
);

INVxp67_ASAP7_75t_L g1217 ( 
.A(n_926),
.Y(n_1217)
);

NAND2xp5_ASAP7_75t_L g1218 ( 
.A(n_938),
.B(n_1098),
.Y(n_1218)
);

AOI21xp5_ASAP7_75t_L g1219 ( 
.A1(n_1099),
.A2(n_702),
.B(n_800),
.Y(n_1219)
);

NAND2xp33_ASAP7_75t_L g1220 ( 
.A(n_1009),
.B(n_1010),
.Y(n_1220)
);

AND2x2_ASAP7_75t_L g1221 ( 
.A(n_930),
.B(n_927),
.Y(n_1221)
);

AOI21xp33_ASAP7_75t_L g1222 ( 
.A1(n_1004),
.A2(n_938),
.B(n_1013),
.Y(n_1222)
);

OAI21x1_ASAP7_75t_SL g1223 ( 
.A1(n_1008),
.A2(n_1027),
.B(n_969),
.Y(n_1223)
);

AND2x2_ASAP7_75t_L g1224 ( 
.A(n_930),
.B(n_927),
.Y(n_1224)
);

OAI21x1_ASAP7_75t_L g1225 ( 
.A1(n_982),
.A2(n_1073),
.B(n_961),
.Y(n_1225)
);

AOI21x1_ASAP7_75t_L g1226 ( 
.A1(n_954),
.A2(n_959),
.B(n_955),
.Y(n_1226)
);

INVxp67_ASAP7_75t_L g1227 ( 
.A(n_926),
.Y(n_1227)
);

INVx2_ASAP7_75t_L g1228 ( 
.A(n_953),
.Y(n_1228)
);

OAI21x1_ASAP7_75t_L g1229 ( 
.A1(n_982),
.A2(n_1073),
.B(n_961),
.Y(n_1229)
);

A2O1A1Ixp33_ASAP7_75t_L g1230 ( 
.A1(n_1013),
.A2(n_1041),
.B(n_1004),
.C(n_978),
.Y(n_1230)
);

OAI21xp5_ASAP7_75t_L g1231 ( 
.A1(n_978),
.A2(n_1101),
.B(n_1082),
.Y(n_1231)
);

NAND2xp5_ASAP7_75t_L g1232 ( 
.A(n_938),
.B(n_1098),
.Y(n_1232)
);

INVx3_ASAP7_75t_L g1233 ( 
.A(n_1066),
.Y(n_1233)
);

A2O1A1Ixp33_ASAP7_75t_L g1234 ( 
.A1(n_1013),
.A2(n_1041),
.B(n_1004),
.C(n_978),
.Y(n_1234)
);

OAI21x1_ASAP7_75t_L g1235 ( 
.A1(n_982),
.A2(n_1073),
.B(n_961),
.Y(n_1235)
);

BUFx2_ASAP7_75t_L g1236 ( 
.A(n_926),
.Y(n_1236)
);

AOI21xp5_ASAP7_75t_L g1237 ( 
.A1(n_1099),
.A2(n_702),
.B(n_800),
.Y(n_1237)
);

AOI221xp5_ASAP7_75t_SL g1238 ( 
.A1(n_1058),
.A2(n_769),
.B1(n_1041),
.B2(n_1013),
.C(n_883),
.Y(n_1238)
);

CKINVDCx5p33_ASAP7_75t_R g1239 ( 
.A(n_928),
.Y(n_1239)
);

OAI21x1_ASAP7_75t_L g1240 ( 
.A1(n_982),
.A2(n_1073),
.B(n_961),
.Y(n_1240)
);

AND2x2_ASAP7_75t_L g1241 ( 
.A(n_930),
.B(n_927),
.Y(n_1241)
);

INVx1_ASAP7_75t_L g1242 ( 
.A(n_1080),
.Y(n_1242)
);

OAI21x1_ASAP7_75t_L g1243 ( 
.A1(n_982),
.A2(n_1073),
.B(n_961),
.Y(n_1243)
);

INVx3_ASAP7_75t_L g1244 ( 
.A(n_1066),
.Y(n_1244)
);

AOI21xp5_ASAP7_75t_L g1245 ( 
.A1(n_1099),
.A2(n_702),
.B(n_800),
.Y(n_1245)
);

AOI21xp5_ASAP7_75t_L g1246 ( 
.A1(n_1099),
.A2(n_702),
.B(n_800),
.Y(n_1246)
);

NOR2xp67_ASAP7_75t_L g1247 ( 
.A(n_928),
.B(n_761),
.Y(n_1247)
);

OAI21x1_ASAP7_75t_L g1248 ( 
.A1(n_982),
.A2(n_1073),
.B(n_961),
.Y(n_1248)
);

OAI21x1_ASAP7_75t_L g1249 ( 
.A1(n_982),
.A2(n_1073),
.B(n_961),
.Y(n_1249)
);

AOI21xp5_ASAP7_75t_L g1250 ( 
.A1(n_1099),
.A2(n_702),
.B(n_800),
.Y(n_1250)
);

AOI21x1_ASAP7_75t_L g1251 ( 
.A1(n_954),
.A2(n_959),
.B(n_955),
.Y(n_1251)
);

BUFx3_ASAP7_75t_L g1252 ( 
.A(n_1095),
.Y(n_1252)
);

OAI21xp5_ASAP7_75t_L g1253 ( 
.A1(n_978),
.A2(n_1101),
.B(n_1082),
.Y(n_1253)
);

AOI21xp5_ASAP7_75t_L g1254 ( 
.A1(n_1099),
.A2(n_702),
.B(n_800),
.Y(n_1254)
);

AOI21xp5_ASAP7_75t_L g1255 ( 
.A1(n_1099),
.A2(n_702),
.B(n_800),
.Y(n_1255)
);

AO31x2_ASAP7_75t_L g1256 ( 
.A1(n_998),
.A2(n_1041),
.A3(n_1013),
.B(n_1082),
.Y(n_1256)
);

OAI21x1_ASAP7_75t_L g1257 ( 
.A1(n_982),
.A2(n_1073),
.B(n_961),
.Y(n_1257)
);

INVx1_ASAP7_75t_L g1258 ( 
.A(n_1080),
.Y(n_1258)
);

AND2x4_ASAP7_75t_L g1259 ( 
.A(n_1148),
.B(n_1143),
.Y(n_1259)
);

INVx2_ASAP7_75t_L g1260 ( 
.A(n_1123),
.Y(n_1260)
);

INVx3_ASAP7_75t_L g1261 ( 
.A(n_1182),
.Y(n_1261)
);

NAND2xp5_ASAP7_75t_L g1262 ( 
.A(n_1104),
.B(n_1195),
.Y(n_1262)
);

AND2x2_ASAP7_75t_L g1263 ( 
.A(n_1221),
.B(n_1224),
.Y(n_1263)
);

AOI21xp5_ASAP7_75t_L g1264 ( 
.A1(n_1103),
.A2(n_1108),
.B(n_1115),
.Y(n_1264)
);

INVx1_ASAP7_75t_L g1265 ( 
.A(n_1129),
.Y(n_1265)
);

NOR2x1_ASAP7_75t_SL g1266 ( 
.A(n_1159),
.B(n_1190),
.Y(n_1266)
);

INVx1_ASAP7_75t_SL g1267 ( 
.A(n_1107),
.Y(n_1267)
);

AOI21xp5_ASAP7_75t_L g1268 ( 
.A1(n_1116),
.A2(n_1198),
.B(n_1197),
.Y(n_1268)
);

NAND2xp5_ASAP7_75t_L g1269 ( 
.A(n_1104),
.B(n_1195),
.Y(n_1269)
);

NAND2xp5_ASAP7_75t_SL g1270 ( 
.A(n_1135),
.B(n_1110),
.Y(n_1270)
);

AOI21xp5_ASAP7_75t_L g1271 ( 
.A1(n_1197),
.A2(n_1203),
.B(n_1198),
.Y(n_1271)
);

AOI21xp5_ASAP7_75t_L g1272 ( 
.A1(n_1203),
.A2(n_1231),
.B(n_1206),
.Y(n_1272)
);

A2O1A1Ixp33_ASAP7_75t_L g1273 ( 
.A1(n_1230),
.A2(n_1234),
.B(n_1113),
.C(n_1222),
.Y(n_1273)
);

AOI22xp5_ASAP7_75t_L g1274 ( 
.A1(n_1136),
.A2(n_1105),
.B1(n_1205),
.B2(n_1238),
.Y(n_1274)
);

AOI21xp5_ASAP7_75t_L g1275 ( 
.A1(n_1206),
.A2(n_1253),
.B(n_1231),
.Y(n_1275)
);

AND2x4_ASAP7_75t_L g1276 ( 
.A(n_1148),
.B(n_1252),
.Y(n_1276)
);

OAI22xp5_ASAP7_75t_L g1277 ( 
.A1(n_1196),
.A2(n_1232),
.B1(n_1211),
.B2(n_1218),
.Y(n_1277)
);

INVx2_ASAP7_75t_SL g1278 ( 
.A(n_1216),
.Y(n_1278)
);

OAI22xp33_ASAP7_75t_L g1279 ( 
.A1(n_1110),
.A2(n_1232),
.B1(n_1196),
.B2(n_1211),
.Y(n_1279)
);

OAI22xp5_ASAP7_75t_L g1280 ( 
.A1(n_1218),
.A2(n_1119),
.B1(n_1154),
.B2(n_1208),
.Y(n_1280)
);

AND2x4_ASAP7_75t_L g1281 ( 
.A(n_1167),
.B(n_1204),
.Y(n_1281)
);

NAND2xp5_ASAP7_75t_L g1282 ( 
.A(n_1106),
.B(n_1208),
.Y(n_1282)
);

INVx2_ASAP7_75t_L g1283 ( 
.A(n_1199),
.Y(n_1283)
);

BUFx6f_ASAP7_75t_L g1284 ( 
.A(n_1139),
.Y(n_1284)
);

HB1xp67_ASAP7_75t_L g1285 ( 
.A(n_1212),
.Y(n_1285)
);

NAND2xp5_ASAP7_75t_L g1286 ( 
.A(n_1106),
.B(n_1222),
.Y(n_1286)
);

BUFx6f_ASAP7_75t_L g1287 ( 
.A(n_1139),
.Y(n_1287)
);

BUFx3_ASAP7_75t_L g1288 ( 
.A(n_1236),
.Y(n_1288)
);

A2O1A1Ixp33_ASAP7_75t_L g1289 ( 
.A1(n_1118),
.A2(n_1151),
.B(n_1161),
.C(n_1127),
.Y(n_1289)
);

INVx1_ASAP7_75t_L g1290 ( 
.A(n_1141),
.Y(n_1290)
);

INVxp67_ASAP7_75t_SL g1291 ( 
.A(n_1114),
.Y(n_1291)
);

BUFx4f_ASAP7_75t_L g1292 ( 
.A(n_1204),
.Y(n_1292)
);

BUFx2_ASAP7_75t_L g1293 ( 
.A(n_1217),
.Y(n_1293)
);

NAND3xp33_ASAP7_75t_L g1294 ( 
.A(n_1220),
.B(n_1118),
.C(n_1127),
.Y(n_1294)
);

AND2x2_ASAP7_75t_L g1295 ( 
.A(n_1241),
.B(n_1213),
.Y(n_1295)
);

OAI22xp5_ASAP7_75t_L g1296 ( 
.A1(n_1119),
.A2(n_1109),
.B1(n_1140),
.B2(n_1168),
.Y(n_1296)
);

BUFx6f_ASAP7_75t_L g1297 ( 
.A(n_1139),
.Y(n_1297)
);

AND2x4_ASAP7_75t_L g1298 ( 
.A(n_1204),
.B(n_1173),
.Y(n_1298)
);

INVx3_ASAP7_75t_SL g1299 ( 
.A(n_1150),
.Y(n_1299)
);

OAI221xp5_ASAP7_75t_L g1300 ( 
.A1(n_1176),
.A2(n_1168),
.B1(n_1253),
.B2(n_1247),
.C(n_1227),
.Y(n_1300)
);

CKINVDCx8_ASAP7_75t_R g1301 ( 
.A(n_1180),
.Y(n_1301)
);

BUFx10_ASAP7_75t_L g1302 ( 
.A(n_1156),
.Y(n_1302)
);

BUFx2_ASAP7_75t_L g1303 ( 
.A(n_1189),
.Y(n_1303)
);

AND2x2_ASAP7_75t_L g1304 ( 
.A(n_1140),
.B(n_1117),
.Y(n_1304)
);

AND2x4_ASAP7_75t_L g1305 ( 
.A(n_1204),
.B(n_1191),
.Y(n_1305)
);

AOI21xp5_ASAP7_75t_SL g1306 ( 
.A1(n_1130),
.A2(n_1170),
.B(n_1144),
.Y(n_1306)
);

AOI21xp5_ASAP7_75t_L g1307 ( 
.A1(n_1201),
.A2(n_1250),
.B(n_1255),
.Y(n_1307)
);

AND2x4_ASAP7_75t_L g1308 ( 
.A(n_1204),
.B(n_1191),
.Y(n_1308)
);

AOI21xp5_ASAP7_75t_L g1309 ( 
.A1(n_1219),
.A2(n_1246),
.B(n_1245),
.Y(n_1309)
);

OR2x6_ASAP7_75t_L g1310 ( 
.A(n_1190),
.B(n_1182),
.Y(n_1310)
);

HB1xp67_ASAP7_75t_L g1311 ( 
.A(n_1142),
.Y(n_1311)
);

AND2x2_ASAP7_75t_L g1312 ( 
.A(n_1145),
.B(n_1215),
.Y(n_1312)
);

INVxp67_ASAP7_75t_L g1313 ( 
.A(n_1239),
.Y(n_1313)
);

INVx2_ASAP7_75t_SL g1314 ( 
.A(n_1202),
.Y(n_1314)
);

NAND2xp5_ASAP7_75t_L g1315 ( 
.A(n_1155),
.B(n_1192),
.Y(n_1315)
);

BUFx2_ASAP7_75t_L g1316 ( 
.A(n_1142),
.Y(n_1316)
);

OAI21xp5_ASAP7_75t_L g1317 ( 
.A1(n_1122),
.A2(n_1144),
.B(n_1155),
.Y(n_1317)
);

AOI21xp5_ASAP7_75t_L g1318 ( 
.A1(n_1237),
.A2(n_1254),
.B(n_1122),
.Y(n_1318)
);

BUFx2_ASAP7_75t_L g1319 ( 
.A(n_1142),
.Y(n_1319)
);

INVx1_ASAP7_75t_SL g1320 ( 
.A(n_1202),
.Y(n_1320)
);

NOR2xp67_ASAP7_75t_SL g1321 ( 
.A(n_1147),
.B(n_1160),
.Y(n_1321)
);

NAND2xp5_ASAP7_75t_L g1322 ( 
.A(n_1192),
.B(n_1158),
.Y(n_1322)
);

BUFx6f_ASAP7_75t_L g1323 ( 
.A(n_1147),
.Y(n_1323)
);

NAND2x1p5_ASAP7_75t_L g1324 ( 
.A(n_1132),
.B(n_1147),
.Y(n_1324)
);

A2O1A1Ixp33_ASAP7_75t_L g1325 ( 
.A1(n_1152),
.A2(n_1134),
.B(n_1133),
.C(n_1174),
.Y(n_1325)
);

BUFx10_ASAP7_75t_L g1326 ( 
.A(n_1156),
.Y(n_1326)
);

OAI22xp33_ASAP7_75t_SL g1327 ( 
.A1(n_1125),
.A2(n_1258),
.B1(n_1209),
.B2(n_1207),
.Y(n_1327)
);

O2A1O1Ixp5_ASAP7_75t_L g1328 ( 
.A1(n_1193),
.A2(n_1251),
.B(n_1226),
.C(n_1149),
.Y(n_1328)
);

AND2x2_ASAP7_75t_L g1329 ( 
.A(n_1137),
.B(n_1242),
.Y(n_1329)
);

INVx3_ASAP7_75t_SL g1330 ( 
.A(n_1202),
.Y(n_1330)
);

AND2x4_ASAP7_75t_L g1331 ( 
.A(n_1132),
.B(n_1244),
.Y(n_1331)
);

AND2x2_ASAP7_75t_SL g1332 ( 
.A(n_1185),
.B(n_1171),
.Y(n_1332)
);

NAND2xp33_ASAP7_75t_L g1333 ( 
.A(n_1160),
.B(n_1178),
.Y(n_1333)
);

INVx1_ASAP7_75t_SL g1334 ( 
.A(n_1160),
.Y(n_1334)
);

AOI21xp5_ASAP7_75t_L g1335 ( 
.A1(n_1124),
.A2(n_1223),
.B(n_1200),
.Y(n_1335)
);

CKINVDCx20_ASAP7_75t_R g1336 ( 
.A(n_1178),
.Y(n_1336)
);

INVx2_ASAP7_75t_L g1337 ( 
.A(n_1210),
.Y(n_1337)
);

INVx1_ASAP7_75t_L g1338 ( 
.A(n_1165),
.Y(n_1338)
);

AND2x2_ASAP7_75t_L g1339 ( 
.A(n_1228),
.B(n_1158),
.Y(n_1339)
);

OAI22xp5_ASAP7_75t_L g1340 ( 
.A1(n_1163),
.A2(n_1177),
.B1(n_1175),
.B2(n_1172),
.Y(n_1340)
);

AND2x4_ASAP7_75t_L g1341 ( 
.A(n_1138),
.B(n_1233),
.Y(n_1341)
);

BUFx6f_ASAP7_75t_L g1342 ( 
.A(n_1138),
.Y(n_1342)
);

INVxp67_ASAP7_75t_L g1343 ( 
.A(n_1233),
.Y(n_1343)
);

HB1xp67_ASAP7_75t_L g1344 ( 
.A(n_1158),
.Y(n_1344)
);

AND2x4_ASAP7_75t_L g1345 ( 
.A(n_1171),
.B(n_1186),
.Y(n_1345)
);

AND2x2_ASAP7_75t_L g1346 ( 
.A(n_1256),
.B(n_1175),
.Y(n_1346)
);

AOI21xp5_ASAP7_75t_L g1347 ( 
.A1(n_1128),
.A2(n_1120),
.B(n_1121),
.Y(n_1347)
);

NAND2xp5_ASAP7_75t_L g1348 ( 
.A(n_1256),
.B(n_1181),
.Y(n_1348)
);

NAND2xp5_ASAP7_75t_L g1349 ( 
.A(n_1256),
.B(n_1174),
.Y(n_1349)
);

INVx3_ASAP7_75t_L g1350 ( 
.A(n_1188),
.Y(n_1350)
);

OAI22xp5_ASAP7_75t_L g1351 ( 
.A1(n_1177),
.A2(n_1169),
.B1(n_1187),
.B2(n_1184),
.Y(n_1351)
);

HB1xp67_ASAP7_75t_L g1352 ( 
.A(n_1153),
.Y(n_1352)
);

OR2x6_ASAP7_75t_L g1353 ( 
.A(n_1183),
.B(n_1126),
.Y(n_1353)
);

OAI22xp5_ASAP7_75t_L g1354 ( 
.A1(n_1179),
.A2(n_1112),
.B1(n_1162),
.B2(n_1153),
.Y(n_1354)
);

BUFx3_ASAP7_75t_L g1355 ( 
.A(n_1164),
.Y(n_1355)
);

AND2x2_ASAP7_75t_L g1356 ( 
.A(n_1153),
.B(n_1131),
.Y(n_1356)
);

INVx2_ASAP7_75t_L g1357 ( 
.A(n_1111),
.Y(n_1357)
);

NOR2xp67_ASAP7_75t_L g1358 ( 
.A(n_1131),
.B(n_1166),
.Y(n_1358)
);

HB1xp67_ASAP7_75t_L g1359 ( 
.A(n_1131),
.Y(n_1359)
);

O2A1O1Ixp33_ASAP7_75t_SL g1360 ( 
.A1(n_1166),
.A2(n_1157),
.B(n_1146),
.C(n_1214),
.Y(n_1360)
);

INVx1_ASAP7_75t_SL g1361 ( 
.A(n_1225),
.Y(n_1361)
);

OAI22xp5_ASAP7_75t_L g1362 ( 
.A1(n_1166),
.A2(n_1229),
.B1(n_1235),
.B2(n_1240),
.Y(n_1362)
);

NAND2xp5_ASAP7_75t_L g1363 ( 
.A(n_1243),
.B(n_1248),
.Y(n_1363)
);

NOR2xp33_ASAP7_75t_SL g1364 ( 
.A(n_1249),
.B(n_1257),
.Y(n_1364)
);

INVx4_ASAP7_75t_L g1365 ( 
.A(n_1139),
.Y(n_1365)
);

NOR2xp33_ASAP7_75t_L g1366 ( 
.A(n_1105),
.B(n_1135),
.Y(n_1366)
);

INVx3_ASAP7_75t_L g1367 ( 
.A(n_1182),
.Y(n_1367)
);

INVx2_ASAP7_75t_L g1368 ( 
.A(n_1123),
.Y(n_1368)
);

OAI22xp5_ASAP7_75t_L g1369 ( 
.A1(n_1230),
.A2(n_1234),
.B1(n_1195),
.B2(n_1196),
.Y(n_1369)
);

AO21x1_ASAP7_75t_L g1370 ( 
.A1(n_1113),
.A2(n_1222),
.B(n_1208),
.Y(n_1370)
);

AND2x4_ASAP7_75t_L g1371 ( 
.A(n_1148),
.B(n_1143),
.Y(n_1371)
);

INVx1_ASAP7_75t_L g1372 ( 
.A(n_1129),
.Y(n_1372)
);

AND2x2_ASAP7_75t_L g1373 ( 
.A(n_1221),
.B(n_1224),
.Y(n_1373)
);

INVx2_ASAP7_75t_L g1374 ( 
.A(n_1123),
.Y(n_1374)
);

CKINVDCx20_ASAP7_75t_R g1375 ( 
.A(n_1145),
.Y(n_1375)
);

HB1xp67_ASAP7_75t_L g1376 ( 
.A(n_1212),
.Y(n_1376)
);

BUFx12f_ASAP7_75t_L g1377 ( 
.A(n_1150),
.Y(n_1377)
);

INVx2_ASAP7_75t_L g1378 ( 
.A(n_1123),
.Y(n_1378)
);

INVx2_ASAP7_75t_L g1379 ( 
.A(n_1123),
.Y(n_1379)
);

NAND2xp5_ASAP7_75t_L g1380 ( 
.A(n_1104),
.B(n_1195),
.Y(n_1380)
);

OAI22xp5_ASAP7_75t_L g1381 ( 
.A1(n_1230),
.A2(n_1234),
.B1(n_1110),
.B2(n_1195),
.Y(n_1381)
);

INVxp67_ASAP7_75t_L g1382 ( 
.A(n_1212),
.Y(n_1382)
);

AOI21xp5_ASAP7_75t_L g1383 ( 
.A1(n_1103),
.A2(n_702),
.B(n_1108),
.Y(n_1383)
);

OAI21x1_ASAP7_75t_L g1384 ( 
.A1(n_1111),
.A2(n_1214),
.B(n_1194),
.Y(n_1384)
);

BUFx2_ASAP7_75t_L g1385 ( 
.A(n_1216),
.Y(n_1385)
);

CKINVDCx20_ASAP7_75t_R g1386 ( 
.A(n_1145),
.Y(n_1386)
);

INVx1_ASAP7_75t_L g1387 ( 
.A(n_1129),
.Y(n_1387)
);

NOR2xp33_ASAP7_75t_L g1388 ( 
.A(n_1105),
.B(n_1135),
.Y(n_1388)
);

INVx2_ASAP7_75t_SL g1389 ( 
.A(n_1216),
.Y(n_1389)
);

OR2x6_ASAP7_75t_L g1390 ( 
.A(n_1191),
.B(n_1190),
.Y(n_1390)
);

OR2x6_ASAP7_75t_L g1391 ( 
.A(n_1191),
.B(n_1190),
.Y(n_1391)
);

OAI22xp5_ASAP7_75t_L g1392 ( 
.A1(n_1230),
.A2(n_1234),
.B1(n_1195),
.B2(n_1196),
.Y(n_1392)
);

NAND2xp5_ASAP7_75t_SL g1393 ( 
.A(n_1135),
.B(n_930),
.Y(n_1393)
);

BUFx6f_ASAP7_75t_SL g1394 ( 
.A(n_1252),
.Y(n_1394)
);

OR2x6_ASAP7_75t_L g1395 ( 
.A(n_1191),
.B(n_1190),
.Y(n_1395)
);

BUFx6f_ASAP7_75t_L g1396 ( 
.A(n_1139),
.Y(n_1396)
);

AND2x4_ASAP7_75t_L g1397 ( 
.A(n_1148),
.B(n_1143),
.Y(n_1397)
);

NOR2xp33_ASAP7_75t_L g1398 ( 
.A(n_1105),
.B(n_1135),
.Y(n_1398)
);

NAND2xp5_ASAP7_75t_L g1399 ( 
.A(n_1104),
.B(n_1195),
.Y(n_1399)
);

NOR2xp33_ASAP7_75t_SL g1400 ( 
.A(n_1230),
.B(n_1058),
.Y(n_1400)
);

AOI21xp5_ASAP7_75t_L g1401 ( 
.A1(n_1103),
.A2(n_702),
.B(n_1108),
.Y(n_1401)
);

BUFx12f_ASAP7_75t_L g1402 ( 
.A(n_1150),
.Y(n_1402)
);

INVx3_ASAP7_75t_L g1403 ( 
.A(n_1182),
.Y(n_1403)
);

INVx1_ASAP7_75t_SL g1404 ( 
.A(n_1107),
.Y(n_1404)
);

OR2x6_ASAP7_75t_L g1405 ( 
.A(n_1191),
.B(n_1190),
.Y(n_1405)
);

NAND2xp5_ASAP7_75t_SL g1406 ( 
.A(n_1135),
.B(n_930),
.Y(n_1406)
);

BUFx4f_ASAP7_75t_L g1407 ( 
.A(n_1204),
.Y(n_1407)
);

AOI21xp5_ASAP7_75t_L g1408 ( 
.A1(n_1103),
.A2(n_702),
.B(n_1108),
.Y(n_1408)
);

AND2x4_ASAP7_75t_L g1409 ( 
.A(n_1148),
.B(n_1143),
.Y(n_1409)
);

NOR2xp33_ASAP7_75t_L g1410 ( 
.A(n_1105),
.B(n_1135),
.Y(n_1410)
);

AND2x4_ASAP7_75t_L g1411 ( 
.A(n_1148),
.B(n_1143),
.Y(n_1411)
);

AND2x4_ASAP7_75t_L g1412 ( 
.A(n_1148),
.B(n_1143),
.Y(n_1412)
);

AOI21xp5_ASAP7_75t_L g1413 ( 
.A1(n_1103),
.A2(n_702),
.B(n_1108),
.Y(n_1413)
);

NAND2xp5_ASAP7_75t_L g1414 ( 
.A(n_1104),
.B(n_1195),
.Y(n_1414)
);

O2A1O1Ixp33_ASAP7_75t_L g1415 ( 
.A1(n_1208),
.A2(n_1222),
.B(n_1234),
.C(n_1230),
.Y(n_1415)
);

BUFx6f_ASAP7_75t_L g1416 ( 
.A(n_1139),
.Y(n_1416)
);

NAND2xp5_ASAP7_75t_L g1417 ( 
.A(n_1104),
.B(n_1195),
.Y(n_1417)
);

OR2x2_ASAP7_75t_L g1418 ( 
.A(n_1107),
.B(n_1221),
.Y(n_1418)
);

AOI22xp33_ASAP7_75t_L g1419 ( 
.A1(n_1366),
.A2(n_1388),
.B1(n_1410),
.B2(n_1398),
.Y(n_1419)
);

NAND2xp5_ASAP7_75t_L g1420 ( 
.A(n_1270),
.B(n_1279),
.Y(n_1420)
);

INVx2_ASAP7_75t_SL g1421 ( 
.A(n_1288),
.Y(n_1421)
);

INVx1_ASAP7_75t_SL g1422 ( 
.A(n_1267),
.Y(n_1422)
);

OAI22xp33_ASAP7_75t_L g1423 ( 
.A1(n_1400),
.A2(n_1300),
.B1(n_1417),
.B2(n_1414),
.Y(n_1423)
);

BUFx2_ASAP7_75t_L g1424 ( 
.A(n_1390),
.Y(n_1424)
);

INVx3_ASAP7_75t_L g1425 ( 
.A(n_1292),
.Y(n_1425)
);

AND2x2_ASAP7_75t_L g1426 ( 
.A(n_1274),
.B(n_1265),
.Y(n_1426)
);

OAI22xp5_ASAP7_75t_L g1427 ( 
.A1(n_1262),
.A2(n_1399),
.B1(n_1269),
.B2(n_1380),
.Y(n_1427)
);

OAI21x1_ASAP7_75t_L g1428 ( 
.A1(n_1384),
.A2(n_1309),
.B(n_1307),
.Y(n_1428)
);

AOI22xp33_ASAP7_75t_L g1429 ( 
.A1(n_1400),
.A2(n_1370),
.B1(n_1381),
.B2(n_1392),
.Y(n_1429)
);

BUFx3_ASAP7_75t_L g1430 ( 
.A(n_1336),
.Y(n_1430)
);

AOI22xp33_ASAP7_75t_L g1431 ( 
.A1(n_1369),
.A2(n_1392),
.B1(n_1295),
.B2(n_1296),
.Y(n_1431)
);

BUFx2_ASAP7_75t_R g1432 ( 
.A(n_1301),
.Y(n_1432)
);

INVx6_ASAP7_75t_L g1433 ( 
.A(n_1365),
.Y(n_1433)
);

NAND2x1p5_ASAP7_75t_L g1434 ( 
.A(n_1292),
.B(n_1407),
.Y(n_1434)
);

INVx2_ASAP7_75t_L g1435 ( 
.A(n_1290),
.Y(n_1435)
);

BUFx2_ASAP7_75t_SL g1436 ( 
.A(n_1375),
.Y(n_1436)
);

CKINVDCx11_ASAP7_75t_R g1437 ( 
.A(n_1299),
.Y(n_1437)
);

AOI22xp33_ASAP7_75t_L g1438 ( 
.A1(n_1369),
.A2(n_1280),
.B1(n_1393),
.B2(n_1406),
.Y(n_1438)
);

NAND2x1p5_ASAP7_75t_L g1439 ( 
.A(n_1407),
.B(n_1261),
.Y(n_1439)
);

BUFx2_ASAP7_75t_R g1440 ( 
.A(n_1330),
.Y(n_1440)
);

INVx1_ASAP7_75t_L g1441 ( 
.A(n_1338),
.Y(n_1441)
);

INVx1_ASAP7_75t_L g1442 ( 
.A(n_1260),
.Y(n_1442)
);

BUFx2_ASAP7_75t_SL g1443 ( 
.A(n_1386),
.Y(n_1443)
);

CKINVDCx20_ASAP7_75t_R g1444 ( 
.A(n_1377),
.Y(n_1444)
);

INVx1_ASAP7_75t_L g1445 ( 
.A(n_1283),
.Y(n_1445)
);

OA21x2_ASAP7_75t_L g1446 ( 
.A1(n_1328),
.A2(n_1268),
.B(n_1325),
.Y(n_1446)
);

OAI21x1_ASAP7_75t_L g1447 ( 
.A1(n_1347),
.A2(n_1401),
.B(n_1383),
.Y(n_1447)
);

HB1xp67_ASAP7_75t_L g1448 ( 
.A(n_1267),
.Y(n_1448)
);

INVx1_ASAP7_75t_L g1449 ( 
.A(n_1337),
.Y(n_1449)
);

INVx1_ASAP7_75t_L g1450 ( 
.A(n_1368),
.Y(n_1450)
);

AOI22xp33_ASAP7_75t_L g1451 ( 
.A1(n_1280),
.A2(n_1391),
.B1(n_1390),
.B2(n_1395),
.Y(n_1451)
);

INVx1_ASAP7_75t_L g1452 ( 
.A(n_1374),
.Y(n_1452)
);

AND2x2_ASAP7_75t_L g1453 ( 
.A(n_1274),
.B(n_1372),
.Y(n_1453)
);

BUFx12f_ASAP7_75t_L g1454 ( 
.A(n_1302),
.Y(n_1454)
);

AOI22xp5_ASAP7_75t_L g1455 ( 
.A1(n_1259),
.A2(n_1397),
.B1(n_1409),
.B2(n_1412),
.Y(n_1455)
);

CKINVDCx11_ASAP7_75t_R g1456 ( 
.A(n_1402),
.Y(n_1456)
);

INVx1_ASAP7_75t_L g1457 ( 
.A(n_1378),
.Y(n_1457)
);

CKINVDCx6p67_ASAP7_75t_R g1458 ( 
.A(n_1394),
.Y(n_1458)
);

INVx2_ASAP7_75t_L g1459 ( 
.A(n_1387),
.Y(n_1459)
);

AND2x2_ASAP7_75t_L g1460 ( 
.A(n_1282),
.B(n_1286),
.Y(n_1460)
);

CKINVDCx8_ASAP7_75t_R g1461 ( 
.A(n_1385),
.Y(n_1461)
);

INVx1_ASAP7_75t_L g1462 ( 
.A(n_1379),
.Y(n_1462)
);

INVx2_ASAP7_75t_L g1463 ( 
.A(n_1339),
.Y(n_1463)
);

HB1xp67_ASAP7_75t_L g1464 ( 
.A(n_1404),
.Y(n_1464)
);

AOI21xp5_ASAP7_75t_L g1465 ( 
.A1(n_1264),
.A2(n_1413),
.B(n_1408),
.Y(n_1465)
);

NAND2xp5_ASAP7_75t_L g1466 ( 
.A(n_1277),
.B(n_1263),
.Y(n_1466)
);

INVxp67_ASAP7_75t_SL g1467 ( 
.A(n_1285),
.Y(n_1467)
);

AOI22xp33_ASAP7_75t_L g1468 ( 
.A1(n_1390),
.A2(n_1391),
.B1(n_1395),
.B2(n_1405),
.Y(n_1468)
);

OAI21x1_ASAP7_75t_L g1469 ( 
.A1(n_1318),
.A2(n_1362),
.B(n_1363),
.Y(n_1469)
);

AND2x2_ASAP7_75t_L g1470 ( 
.A(n_1304),
.B(n_1273),
.Y(n_1470)
);

BUFx2_ASAP7_75t_L g1471 ( 
.A(n_1391),
.Y(n_1471)
);

INVx3_ASAP7_75t_L g1472 ( 
.A(n_1345),
.Y(n_1472)
);

BUFx12f_ASAP7_75t_L g1473 ( 
.A(n_1302),
.Y(n_1473)
);

CKINVDCx11_ASAP7_75t_R g1474 ( 
.A(n_1326),
.Y(n_1474)
);

AND2x2_ASAP7_75t_L g1475 ( 
.A(n_1315),
.B(n_1346),
.Y(n_1475)
);

BUFx12f_ASAP7_75t_L g1476 ( 
.A(n_1326),
.Y(n_1476)
);

BUFx3_ASAP7_75t_L g1477 ( 
.A(n_1276),
.Y(n_1477)
);

HB1xp67_ASAP7_75t_L g1478 ( 
.A(n_1404),
.Y(n_1478)
);

OAI21xp5_ASAP7_75t_SL g1479 ( 
.A1(n_1415),
.A2(n_1289),
.B(n_1294),
.Y(n_1479)
);

OA21x2_ASAP7_75t_L g1480 ( 
.A1(n_1271),
.A2(n_1275),
.B(n_1272),
.Y(n_1480)
);

OAI22xp5_ASAP7_75t_L g1481 ( 
.A1(n_1277),
.A2(n_1405),
.B1(n_1395),
.B2(n_1418),
.Y(n_1481)
);

INVx6_ASAP7_75t_L g1482 ( 
.A(n_1365),
.Y(n_1482)
);

OR2x6_ASAP7_75t_L g1483 ( 
.A(n_1310),
.B(n_1306),
.Y(n_1483)
);

BUFx6f_ASAP7_75t_L g1484 ( 
.A(n_1284),
.Y(n_1484)
);

CKINVDCx11_ASAP7_75t_R g1485 ( 
.A(n_1293),
.Y(n_1485)
);

INVx1_ASAP7_75t_L g1486 ( 
.A(n_1327),
.Y(n_1486)
);

INVx1_ASAP7_75t_L g1487 ( 
.A(n_1327),
.Y(n_1487)
);

INVx1_ASAP7_75t_L g1488 ( 
.A(n_1259),
.Y(n_1488)
);

BUFx2_ASAP7_75t_L g1489 ( 
.A(n_1405),
.Y(n_1489)
);

OR2x2_ASAP7_75t_L g1490 ( 
.A(n_1348),
.B(n_1349),
.Y(n_1490)
);

BUFx6f_ASAP7_75t_L g1491 ( 
.A(n_1284),
.Y(n_1491)
);

INVx1_ASAP7_75t_L g1492 ( 
.A(n_1371),
.Y(n_1492)
);

OR2x6_ASAP7_75t_L g1493 ( 
.A(n_1310),
.B(n_1335),
.Y(n_1493)
);

BUFx6f_ASAP7_75t_L g1494 ( 
.A(n_1284),
.Y(n_1494)
);

NOR2xp33_ASAP7_75t_L g1495 ( 
.A(n_1373),
.B(n_1371),
.Y(n_1495)
);

OAI22xp33_ASAP7_75t_L g1496 ( 
.A1(n_1294),
.A2(n_1310),
.B1(n_1278),
.B2(n_1389),
.Y(n_1496)
);

INVx1_ASAP7_75t_L g1497 ( 
.A(n_1397),
.Y(n_1497)
);

AOI22xp33_ASAP7_75t_L g1498 ( 
.A1(n_1409),
.A2(n_1412),
.B1(n_1411),
.B2(n_1317),
.Y(n_1498)
);

AO21x2_ASAP7_75t_L g1499 ( 
.A1(n_1358),
.A2(n_1354),
.B(n_1360),
.Y(n_1499)
);

AND2x4_ASAP7_75t_L g1500 ( 
.A(n_1281),
.B(n_1308),
.Y(n_1500)
);

AOI22xp33_ASAP7_75t_SL g1501 ( 
.A1(n_1266),
.A2(n_1411),
.B1(n_1317),
.B2(n_1281),
.Y(n_1501)
);

HB1xp67_ASAP7_75t_L g1502 ( 
.A(n_1376),
.Y(n_1502)
);

OAI22xp5_ASAP7_75t_L g1503 ( 
.A1(n_1382),
.A2(n_1332),
.B1(n_1322),
.B2(n_1298),
.Y(n_1503)
);

OAI21xp5_ASAP7_75t_L g1504 ( 
.A1(n_1351),
.A2(n_1340),
.B(n_1358),
.Y(n_1504)
);

BUFx10_ASAP7_75t_L g1505 ( 
.A(n_1394),
.Y(n_1505)
);

AOI21x1_ASAP7_75t_L g1506 ( 
.A1(n_1340),
.A2(n_1351),
.B(n_1357),
.Y(n_1506)
);

INVx1_ASAP7_75t_L g1507 ( 
.A(n_1344),
.Y(n_1507)
);

INVx1_ASAP7_75t_L g1508 ( 
.A(n_1311),
.Y(n_1508)
);

BUFx6f_ASAP7_75t_L g1509 ( 
.A(n_1287),
.Y(n_1509)
);

INVx1_ASAP7_75t_SL g1510 ( 
.A(n_1312),
.Y(n_1510)
);

INVx3_ASAP7_75t_L g1511 ( 
.A(n_1308),
.Y(n_1511)
);

AOI22xp33_ASAP7_75t_L g1512 ( 
.A1(n_1298),
.A2(n_1303),
.B1(n_1352),
.B2(n_1356),
.Y(n_1512)
);

AOI22xp33_ASAP7_75t_L g1513 ( 
.A1(n_1359),
.A2(n_1313),
.B1(n_1403),
.B2(n_1367),
.Y(n_1513)
);

AOI21x1_ASAP7_75t_L g1514 ( 
.A1(n_1353),
.A2(n_1321),
.B(n_1316),
.Y(n_1514)
);

BUFx2_ASAP7_75t_R g1515 ( 
.A(n_1319),
.Y(n_1515)
);

OAI22xp5_ASAP7_75t_L g1516 ( 
.A1(n_1291),
.A2(n_1343),
.B1(n_1320),
.B2(n_1367),
.Y(n_1516)
);

INVx1_ASAP7_75t_L g1517 ( 
.A(n_1341),
.Y(n_1517)
);

OAI21xp5_ASAP7_75t_L g1518 ( 
.A1(n_1353),
.A2(n_1361),
.B(n_1355),
.Y(n_1518)
);

HB1xp67_ASAP7_75t_L g1519 ( 
.A(n_1320),
.Y(n_1519)
);

CKINVDCx11_ASAP7_75t_R g1520 ( 
.A(n_1287),
.Y(n_1520)
);

OR2x2_ASAP7_75t_L g1521 ( 
.A(n_1353),
.B(n_1361),
.Y(n_1521)
);

HB1xp67_ASAP7_75t_SL g1522 ( 
.A(n_1287),
.Y(n_1522)
);

AOI22xp5_ASAP7_75t_L g1523 ( 
.A1(n_1314),
.A2(n_1331),
.B1(n_1334),
.B2(n_1333),
.Y(n_1523)
);

CKINVDCx11_ASAP7_75t_R g1524 ( 
.A(n_1297),
.Y(n_1524)
);

INVx1_ASAP7_75t_L g1525 ( 
.A(n_1342),
.Y(n_1525)
);

INVx2_ASAP7_75t_L g1526 ( 
.A(n_1350),
.Y(n_1526)
);

INVx1_ASAP7_75t_L g1527 ( 
.A(n_1342),
.Y(n_1527)
);

INVx1_ASAP7_75t_SL g1528 ( 
.A(n_1334),
.Y(n_1528)
);

OAI22xp33_ASAP7_75t_L g1529 ( 
.A1(n_1324),
.A2(n_1297),
.B1(n_1323),
.B2(n_1396),
.Y(n_1529)
);

AOI21x1_ASAP7_75t_L g1530 ( 
.A1(n_1364),
.A2(n_1297),
.B(n_1323),
.Y(n_1530)
);

INVx1_ASAP7_75t_L g1531 ( 
.A(n_1396),
.Y(n_1531)
);

OAI21x1_ASAP7_75t_SL g1532 ( 
.A1(n_1364),
.A2(n_1396),
.B(n_1416),
.Y(n_1532)
);

NAND2x1p5_ASAP7_75t_L g1533 ( 
.A(n_1416),
.B(n_1292),
.Y(n_1533)
);

AO21x1_ASAP7_75t_SL g1534 ( 
.A1(n_1416),
.A2(n_1322),
.B(n_1348),
.Y(n_1534)
);

INVx1_ASAP7_75t_L g1535 ( 
.A(n_1329),
.Y(n_1535)
);

BUFx6f_ASAP7_75t_L g1536 ( 
.A(n_1284),
.Y(n_1536)
);

AOI22xp33_ASAP7_75t_L g1537 ( 
.A1(n_1366),
.A2(n_859),
.B1(n_1136),
.B2(n_1388),
.Y(n_1537)
);

INVx1_ASAP7_75t_L g1538 ( 
.A(n_1329),
.Y(n_1538)
);

AOI22xp5_ASAP7_75t_L g1539 ( 
.A1(n_1366),
.A2(n_1398),
.B1(n_1410),
.B2(n_1388),
.Y(n_1539)
);

BUFx3_ASAP7_75t_L g1540 ( 
.A(n_1336),
.Y(n_1540)
);

INVx1_ASAP7_75t_L g1541 ( 
.A(n_1329),
.Y(n_1541)
);

OAI22xp33_ASAP7_75t_L g1542 ( 
.A1(n_1400),
.A2(n_763),
.B1(n_546),
.B2(n_549),
.Y(n_1542)
);

AND2x4_ASAP7_75t_L g1543 ( 
.A(n_1281),
.B(n_1305),
.Y(n_1543)
);

AND2x4_ASAP7_75t_L g1544 ( 
.A(n_1281),
.B(n_1305),
.Y(n_1544)
);

AOI22xp33_ASAP7_75t_L g1545 ( 
.A1(n_1366),
.A2(n_859),
.B1(n_1136),
.B2(n_1388),
.Y(n_1545)
);

INVx1_ASAP7_75t_L g1546 ( 
.A(n_1329),
.Y(n_1546)
);

INVx1_ASAP7_75t_L g1547 ( 
.A(n_1329),
.Y(n_1547)
);

AO21x1_ASAP7_75t_SL g1548 ( 
.A1(n_1322),
.A2(n_1349),
.B(n_1348),
.Y(n_1548)
);

BUFx10_ASAP7_75t_L g1549 ( 
.A(n_1394),
.Y(n_1549)
);

INVx2_ASAP7_75t_SL g1550 ( 
.A(n_1288),
.Y(n_1550)
);

INVx2_ASAP7_75t_L g1551 ( 
.A(n_1329),
.Y(n_1551)
);

AND2x2_ASAP7_75t_L g1552 ( 
.A(n_1274),
.B(n_1265),
.Y(n_1552)
);

NOR2xp33_ASAP7_75t_L g1553 ( 
.A(n_1366),
.B(n_1388),
.Y(n_1553)
);

BUFx10_ASAP7_75t_L g1554 ( 
.A(n_1394),
.Y(n_1554)
);

CKINVDCx11_ASAP7_75t_R g1555 ( 
.A(n_1301),
.Y(n_1555)
);

AOI22xp33_ASAP7_75t_L g1556 ( 
.A1(n_1366),
.A2(n_859),
.B1(n_1136),
.B2(n_1388),
.Y(n_1556)
);

AOI22xp33_ASAP7_75t_L g1557 ( 
.A1(n_1366),
.A2(n_859),
.B1(n_1136),
.B2(n_1388),
.Y(n_1557)
);

BUFx2_ASAP7_75t_R g1558 ( 
.A(n_1301),
.Y(n_1558)
);

OAI22xp33_ASAP7_75t_L g1559 ( 
.A1(n_1400),
.A2(n_763),
.B1(n_546),
.B2(n_549),
.Y(n_1559)
);

BUFx3_ASAP7_75t_L g1560 ( 
.A(n_1336),
.Y(n_1560)
);

NAND2xp5_ASAP7_75t_L g1561 ( 
.A(n_1366),
.B(n_1388),
.Y(n_1561)
);

NAND2xp5_ASAP7_75t_L g1562 ( 
.A(n_1366),
.B(n_1388),
.Y(n_1562)
);

INVx2_ASAP7_75t_L g1563 ( 
.A(n_1329),
.Y(n_1563)
);

INVx1_ASAP7_75t_L g1564 ( 
.A(n_1329),
.Y(n_1564)
);

CKINVDCx20_ASAP7_75t_R g1565 ( 
.A(n_1375),
.Y(n_1565)
);

BUFx8_ASAP7_75t_SL g1566 ( 
.A(n_1377),
.Y(n_1566)
);

OA21x2_ASAP7_75t_L g1567 ( 
.A1(n_1504),
.A2(n_1465),
.B(n_1447),
.Y(n_1567)
);

HB1xp67_ASAP7_75t_L g1568 ( 
.A(n_1448),
.Y(n_1568)
);

BUFx12f_ASAP7_75t_L g1569 ( 
.A(n_1555),
.Y(n_1569)
);

NAND2xp5_ASAP7_75t_L g1570 ( 
.A(n_1460),
.B(n_1553),
.Y(n_1570)
);

NAND2xp5_ASAP7_75t_L g1571 ( 
.A(n_1460),
.B(n_1553),
.Y(n_1571)
);

CKINVDCx14_ASAP7_75t_R g1572 ( 
.A(n_1555),
.Y(n_1572)
);

OAI21x1_ASAP7_75t_L g1573 ( 
.A1(n_1447),
.A2(n_1428),
.B(n_1469),
.Y(n_1573)
);

AND2x2_ASAP7_75t_L g1574 ( 
.A(n_1475),
.B(n_1463),
.Y(n_1574)
);

INVx1_ASAP7_75t_L g1575 ( 
.A(n_1507),
.Y(n_1575)
);

NAND2xp5_ASAP7_75t_L g1576 ( 
.A(n_1427),
.B(n_1539),
.Y(n_1576)
);

AND2x2_ASAP7_75t_L g1577 ( 
.A(n_1475),
.B(n_1470),
.Y(n_1577)
);

INVx1_ASAP7_75t_L g1578 ( 
.A(n_1486),
.Y(n_1578)
);

NAND2xp5_ASAP7_75t_L g1579 ( 
.A(n_1419),
.B(n_1561),
.Y(n_1579)
);

OAI21xp5_ASAP7_75t_L g1580 ( 
.A1(n_1542),
.A2(n_1559),
.B(n_1479),
.Y(n_1580)
);

NOR2xp33_ASAP7_75t_L g1581 ( 
.A(n_1562),
.B(n_1495),
.Y(n_1581)
);

INVx1_ASAP7_75t_L g1582 ( 
.A(n_1487),
.Y(n_1582)
);

INVx1_ASAP7_75t_L g1583 ( 
.A(n_1521),
.Y(n_1583)
);

AND2x2_ASAP7_75t_L g1584 ( 
.A(n_1470),
.B(n_1548),
.Y(n_1584)
);

INVx5_ASAP7_75t_SL g1585 ( 
.A(n_1483),
.Y(n_1585)
);

NOR2xp33_ASAP7_75t_L g1586 ( 
.A(n_1495),
.B(n_1510),
.Y(n_1586)
);

INVxp67_ASAP7_75t_L g1587 ( 
.A(n_1464),
.Y(n_1587)
);

HB1xp67_ASAP7_75t_L g1588 ( 
.A(n_1478),
.Y(n_1588)
);

OR2x2_ASAP7_75t_L g1589 ( 
.A(n_1490),
.B(n_1466),
.Y(n_1589)
);

INVx1_ASAP7_75t_L g1590 ( 
.A(n_1521),
.Y(n_1590)
);

AND2x2_ASAP7_75t_L g1591 ( 
.A(n_1490),
.B(n_1426),
.Y(n_1591)
);

AOI21x1_ASAP7_75t_L g1592 ( 
.A1(n_1530),
.A2(n_1506),
.B(n_1514),
.Y(n_1592)
);

OAI21xp5_ASAP7_75t_L g1593 ( 
.A1(n_1537),
.A2(n_1556),
.B(n_1545),
.Y(n_1593)
);

AND2x2_ASAP7_75t_L g1594 ( 
.A(n_1426),
.B(n_1453),
.Y(n_1594)
);

AOI21x1_ASAP7_75t_L g1595 ( 
.A1(n_1420),
.A2(n_1446),
.B(n_1483),
.Y(n_1595)
);

AOI21x1_ASAP7_75t_L g1596 ( 
.A1(n_1446),
.A2(n_1483),
.B(n_1516),
.Y(n_1596)
);

INVx1_ASAP7_75t_L g1597 ( 
.A(n_1435),
.Y(n_1597)
);

INVx2_ASAP7_75t_SL g1598 ( 
.A(n_1435),
.Y(n_1598)
);

INVx1_ASAP7_75t_L g1599 ( 
.A(n_1441),
.Y(n_1599)
);

AND2x2_ASAP7_75t_L g1600 ( 
.A(n_1453),
.B(n_1552),
.Y(n_1600)
);

BUFx6f_ASAP7_75t_L g1601 ( 
.A(n_1434),
.Y(n_1601)
);

AO21x2_ASAP7_75t_L g1602 ( 
.A1(n_1499),
.A2(n_1518),
.B(n_1526),
.Y(n_1602)
);

BUFx2_ASAP7_75t_SL g1603 ( 
.A(n_1461),
.Y(n_1603)
);

INVx1_ASAP7_75t_L g1604 ( 
.A(n_1459),
.Y(n_1604)
);

OR2x2_ASAP7_75t_L g1605 ( 
.A(n_1424),
.B(n_1471),
.Y(n_1605)
);

BUFx6f_ASAP7_75t_L g1606 ( 
.A(n_1434),
.Y(n_1606)
);

NAND2x1_ASAP7_75t_L g1607 ( 
.A(n_1483),
.B(n_1493),
.Y(n_1607)
);

AND2x4_ASAP7_75t_L g1608 ( 
.A(n_1511),
.B(n_1500),
.Y(n_1608)
);

AND2x4_ASAP7_75t_L g1609 ( 
.A(n_1500),
.B(n_1543),
.Y(n_1609)
);

BUFx2_ASAP7_75t_L g1610 ( 
.A(n_1424),
.Y(n_1610)
);

INVxp67_ASAP7_75t_L g1611 ( 
.A(n_1502),
.Y(n_1611)
);

INVxp67_ASAP7_75t_L g1612 ( 
.A(n_1519),
.Y(n_1612)
);

INVx1_ASAP7_75t_L g1613 ( 
.A(n_1472),
.Y(n_1613)
);

BUFx12f_ASAP7_75t_L g1614 ( 
.A(n_1456),
.Y(n_1614)
);

AND2x2_ASAP7_75t_L g1615 ( 
.A(n_1552),
.B(n_1451),
.Y(n_1615)
);

INVx1_ASAP7_75t_L g1616 ( 
.A(n_1472),
.Y(n_1616)
);

AO21x2_ASAP7_75t_L g1617 ( 
.A1(n_1499),
.A2(n_1532),
.B(n_1423),
.Y(n_1617)
);

AOI21x1_ASAP7_75t_L g1618 ( 
.A1(n_1446),
.A2(n_1493),
.B(n_1480),
.Y(n_1618)
);

BUFx2_ASAP7_75t_L g1619 ( 
.A(n_1471),
.Y(n_1619)
);

INVx1_ASAP7_75t_L g1620 ( 
.A(n_1493),
.Y(n_1620)
);

INVx1_ASAP7_75t_L g1621 ( 
.A(n_1493),
.Y(n_1621)
);

BUFx2_ASAP7_75t_L g1622 ( 
.A(n_1489),
.Y(n_1622)
);

INVx1_ASAP7_75t_L g1623 ( 
.A(n_1489),
.Y(n_1623)
);

NOR2xp33_ASAP7_75t_L g1624 ( 
.A(n_1488),
.B(n_1492),
.Y(n_1624)
);

BUFx12f_ASAP7_75t_L g1625 ( 
.A(n_1456),
.Y(n_1625)
);

INVx3_ASAP7_75t_L g1626 ( 
.A(n_1500),
.Y(n_1626)
);

INVxp67_ASAP7_75t_L g1627 ( 
.A(n_1422),
.Y(n_1627)
);

NAND2xp5_ASAP7_75t_L g1628 ( 
.A(n_1557),
.B(n_1551),
.Y(n_1628)
);

AND2x2_ASAP7_75t_L g1629 ( 
.A(n_1563),
.B(n_1429),
.Y(n_1629)
);

INVx1_ASAP7_75t_L g1630 ( 
.A(n_1481),
.Y(n_1630)
);

INVx2_ASAP7_75t_SL g1631 ( 
.A(n_1433),
.Y(n_1631)
);

INVx1_ASAP7_75t_L g1632 ( 
.A(n_1442),
.Y(n_1632)
);

AOI21x1_ASAP7_75t_L g1633 ( 
.A1(n_1503),
.A2(n_1449),
.B(n_1445),
.Y(n_1633)
);

INVx2_ASAP7_75t_L g1634 ( 
.A(n_1450),
.Y(n_1634)
);

AND2x4_ASAP7_75t_L g1635 ( 
.A(n_1543),
.B(n_1544),
.Y(n_1635)
);

OR2x2_ASAP7_75t_L g1636 ( 
.A(n_1431),
.B(n_1438),
.Y(n_1636)
);

INVx2_ASAP7_75t_L g1637 ( 
.A(n_1452),
.Y(n_1637)
);

AO21x2_ASAP7_75t_L g1638 ( 
.A1(n_1496),
.A2(n_1529),
.B(n_1457),
.Y(n_1638)
);

HB1xp67_ASAP7_75t_L g1639 ( 
.A(n_1467),
.Y(n_1639)
);

INVx1_ASAP7_75t_L g1640 ( 
.A(n_1462),
.Y(n_1640)
);

OAI21x1_ASAP7_75t_L g1641 ( 
.A1(n_1425),
.A2(n_1439),
.B(n_1468),
.Y(n_1641)
);

INVx1_ASAP7_75t_L g1642 ( 
.A(n_1535),
.Y(n_1642)
);

INVx1_ASAP7_75t_L g1643 ( 
.A(n_1538),
.Y(n_1643)
);

INVx1_ASAP7_75t_SL g1644 ( 
.A(n_1485),
.Y(n_1644)
);

INVx2_ASAP7_75t_L g1645 ( 
.A(n_1541),
.Y(n_1645)
);

OA21x2_ASAP7_75t_L g1646 ( 
.A1(n_1512),
.A2(n_1513),
.B(n_1498),
.Y(n_1646)
);

INVx2_ASAP7_75t_SL g1647 ( 
.A(n_1433),
.Y(n_1647)
);

AO21x2_ASAP7_75t_L g1648 ( 
.A1(n_1546),
.A2(n_1564),
.B(n_1547),
.Y(n_1648)
);

INVx1_ASAP7_75t_L g1649 ( 
.A(n_1501),
.Y(n_1649)
);

OR2x2_ASAP7_75t_L g1650 ( 
.A(n_1497),
.B(n_1508),
.Y(n_1650)
);

INVx3_ASAP7_75t_L g1651 ( 
.A(n_1543),
.Y(n_1651)
);

INVx1_ASAP7_75t_L g1652 ( 
.A(n_1531),
.Y(n_1652)
);

HB1xp67_ASAP7_75t_L g1653 ( 
.A(n_1528),
.Y(n_1653)
);

AND2x2_ASAP7_75t_L g1654 ( 
.A(n_1534),
.B(n_1544),
.Y(n_1654)
);

INVx2_ASAP7_75t_L g1655 ( 
.A(n_1544),
.Y(n_1655)
);

NOR2xp33_ASAP7_75t_L g1656 ( 
.A(n_1485),
.B(n_1565),
.Y(n_1656)
);

BUFx6f_ASAP7_75t_L g1657 ( 
.A(n_1439),
.Y(n_1657)
);

HB1xp67_ASAP7_75t_L g1658 ( 
.A(n_1461),
.Y(n_1658)
);

INVx2_ASAP7_75t_SL g1659 ( 
.A(n_1433),
.Y(n_1659)
);

AND2x2_ASAP7_75t_L g1660 ( 
.A(n_1578),
.B(n_1582),
.Y(n_1660)
);

AND2x2_ASAP7_75t_L g1661 ( 
.A(n_1578),
.B(n_1582),
.Y(n_1661)
);

AND2x2_ASAP7_75t_L g1662 ( 
.A(n_1574),
.B(n_1525),
.Y(n_1662)
);

NAND2xp5_ASAP7_75t_L g1663 ( 
.A(n_1591),
.B(n_1523),
.Y(n_1663)
);

AND2x2_ASAP7_75t_L g1664 ( 
.A(n_1583),
.B(n_1527),
.Y(n_1664)
);

NAND2x1_ASAP7_75t_L g1665 ( 
.A(n_1620),
.B(n_1482),
.Y(n_1665)
);

AND2x4_ASAP7_75t_L g1666 ( 
.A(n_1621),
.B(n_1477),
.Y(n_1666)
);

AND2x2_ASAP7_75t_L g1667 ( 
.A(n_1583),
.B(n_1517),
.Y(n_1667)
);

AOI21xp33_ASAP7_75t_SL g1668 ( 
.A1(n_1576),
.A2(n_1421),
.B(n_1550),
.Y(n_1668)
);

OAI22xp33_ASAP7_75t_L g1669 ( 
.A1(n_1580),
.A2(n_1455),
.B1(n_1430),
.B2(n_1560),
.Y(n_1669)
);

NAND4xp25_ASAP7_75t_L g1670 ( 
.A(n_1579),
.B(n_1581),
.C(n_1593),
.D(n_1570),
.Y(n_1670)
);

NAND3xp33_ASAP7_75t_L g1671 ( 
.A(n_1636),
.B(n_1474),
.C(n_1421),
.Y(n_1671)
);

BUFx2_ASAP7_75t_SL g1672 ( 
.A(n_1631),
.Y(n_1672)
);

OAI221xp5_ASAP7_75t_L g1673 ( 
.A1(n_1636),
.A2(n_1550),
.B1(n_1477),
.B2(n_1430),
.C(n_1560),
.Y(n_1673)
);

NOR2x1_ASAP7_75t_SL g1674 ( 
.A(n_1617),
.B(n_1595),
.Y(n_1674)
);

AND2x2_ASAP7_75t_L g1675 ( 
.A(n_1590),
.B(n_1540),
.Y(n_1675)
);

AND2x2_ASAP7_75t_L g1676 ( 
.A(n_1590),
.B(n_1540),
.Y(n_1676)
);

AND2x2_ASAP7_75t_L g1677 ( 
.A(n_1577),
.B(n_1494),
.Y(n_1677)
);

HB1xp67_ASAP7_75t_L g1678 ( 
.A(n_1648),
.Y(n_1678)
);

NAND2xp5_ASAP7_75t_L g1679 ( 
.A(n_1591),
.B(n_1494),
.Y(n_1679)
);

NAND2xp5_ASAP7_75t_L g1680 ( 
.A(n_1589),
.B(n_1491),
.Y(n_1680)
);

BUFx6f_ASAP7_75t_L g1681 ( 
.A(n_1607),
.Y(n_1681)
);

HB1xp67_ASAP7_75t_L g1682 ( 
.A(n_1648),
.Y(n_1682)
);

NAND2xp5_ASAP7_75t_L g1683 ( 
.A(n_1589),
.B(n_1484),
.Y(n_1683)
);

AOI22xp33_ASAP7_75t_L g1684 ( 
.A1(n_1571),
.A2(n_1437),
.B1(n_1443),
.B2(n_1436),
.Y(n_1684)
);

AND2x2_ASAP7_75t_L g1685 ( 
.A(n_1618),
.B(n_1509),
.Y(n_1685)
);

HB1xp67_ASAP7_75t_L g1686 ( 
.A(n_1648),
.Y(n_1686)
);

OR2x6_ASAP7_75t_L g1687 ( 
.A(n_1607),
.B(n_1533),
.Y(n_1687)
);

AND2x2_ASAP7_75t_L g1688 ( 
.A(n_1602),
.B(n_1509),
.Y(n_1688)
);

INVxp67_ASAP7_75t_SL g1689 ( 
.A(n_1575),
.Y(n_1689)
);

BUFx2_ASAP7_75t_L g1690 ( 
.A(n_1610),
.Y(n_1690)
);

AND2x2_ASAP7_75t_L g1691 ( 
.A(n_1602),
.B(n_1509),
.Y(n_1691)
);

AND2x2_ASAP7_75t_L g1692 ( 
.A(n_1602),
.B(n_1509),
.Y(n_1692)
);

HB1xp67_ASAP7_75t_L g1693 ( 
.A(n_1575),
.Y(n_1693)
);

NOR2x1_ASAP7_75t_SL g1694 ( 
.A(n_1617),
.B(n_1454),
.Y(n_1694)
);

NAND2xp5_ASAP7_75t_L g1695 ( 
.A(n_1594),
.B(n_1536),
.Y(n_1695)
);

OR2x2_ASAP7_75t_L g1696 ( 
.A(n_1623),
.B(n_1536),
.Y(n_1696)
);

AOI221xp5_ASAP7_75t_L g1697 ( 
.A1(n_1587),
.A2(n_1444),
.B1(n_1565),
.B2(n_1533),
.C(n_1440),
.Y(n_1697)
);

BUFx6f_ASAP7_75t_L g1698 ( 
.A(n_1595),
.Y(n_1698)
);

HB1xp67_ASAP7_75t_L g1699 ( 
.A(n_1619),
.Y(n_1699)
);

AND2x2_ASAP7_75t_L g1700 ( 
.A(n_1613),
.B(n_1458),
.Y(n_1700)
);

CKINVDCx5p33_ASAP7_75t_R g1701 ( 
.A(n_1569),
.Y(n_1701)
);

AND2x2_ASAP7_75t_L g1702 ( 
.A(n_1616),
.B(n_1458),
.Y(n_1702)
);

NAND2xp33_ASAP7_75t_SL g1703 ( 
.A(n_1701),
.B(n_1584),
.Y(n_1703)
);

NAND2xp5_ASAP7_75t_SL g1704 ( 
.A(n_1668),
.B(n_1669),
.Y(n_1704)
);

NAND3xp33_ASAP7_75t_L g1705 ( 
.A(n_1670),
.B(n_1639),
.C(n_1624),
.Y(n_1705)
);

NOR2xp33_ASAP7_75t_L g1706 ( 
.A(n_1670),
.B(n_1644),
.Y(n_1706)
);

NAND2xp5_ASAP7_75t_SL g1707 ( 
.A(n_1668),
.B(n_1657),
.Y(n_1707)
);

AND2x2_ASAP7_75t_L g1708 ( 
.A(n_1660),
.B(n_1600),
.Y(n_1708)
);

NAND2xp5_ASAP7_75t_SL g1709 ( 
.A(n_1669),
.B(n_1657),
.Y(n_1709)
);

AND2x2_ASAP7_75t_L g1710 ( 
.A(n_1660),
.B(n_1619),
.Y(n_1710)
);

NAND2xp5_ASAP7_75t_L g1711 ( 
.A(n_1680),
.B(n_1568),
.Y(n_1711)
);

NAND2xp5_ASAP7_75t_L g1712 ( 
.A(n_1683),
.B(n_1588),
.Y(n_1712)
);

OR2x2_ASAP7_75t_L g1713 ( 
.A(n_1699),
.B(n_1690),
.Y(n_1713)
);

OAI22xp5_ASAP7_75t_L g1714 ( 
.A1(n_1671),
.A2(n_1603),
.B1(n_1649),
.B2(n_1515),
.Y(n_1714)
);

AOI211xp5_ASAP7_75t_SL g1715 ( 
.A1(n_1673),
.A2(n_1649),
.B(n_1630),
.C(n_1628),
.Y(n_1715)
);

NAND2xp5_ASAP7_75t_L g1716 ( 
.A(n_1675),
.B(n_1630),
.Y(n_1716)
);

AND2x2_ASAP7_75t_L g1717 ( 
.A(n_1661),
.B(n_1622),
.Y(n_1717)
);

AND2x2_ASAP7_75t_L g1718 ( 
.A(n_1661),
.B(n_1615),
.Y(n_1718)
);

AND2x2_ASAP7_75t_L g1719 ( 
.A(n_1661),
.B(n_1615),
.Y(n_1719)
);

AND2x2_ASAP7_75t_L g1720 ( 
.A(n_1688),
.B(n_1617),
.Y(n_1720)
);

NAND3xp33_ASAP7_75t_L g1721 ( 
.A(n_1671),
.B(n_1612),
.C(n_1627),
.Y(n_1721)
);

NAND2xp5_ASAP7_75t_L g1722 ( 
.A(n_1676),
.B(n_1611),
.Y(n_1722)
);

AND2x2_ASAP7_75t_SL g1723 ( 
.A(n_1698),
.B(n_1567),
.Y(n_1723)
);

AOI221xp5_ASAP7_75t_L g1724 ( 
.A1(n_1673),
.A2(n_1653),
.B1(n_1586),
.B2(n_1643),
.C(n_1642),
.Y(n_1724)
);

HB1xp67_ASAP7_75t_L g1725 ( 
.A(n_1699),
.Y(n_1725)
);

NAND2xp5_ASAP7_75t_L g1726 ( 
.A(n_1664),
.B(n_1599),
.Y(n_1726)
);

OAI22xp5_ASAP7_75t_L g1727 ( 
.A1(n_1684),
.A2(n_1603),
.B1(n_1658),
.B2(n_1585),
.Y(n_1727)
);

NAND2xp5_ASAP7_75t_L g1728 ( 
.A(n_1664),
.B(n_1605),
.Y(n_1728)
);

AND2x2_ASAP7_75t_L g1729 ( 
.A(n_1688),
.B(n_1616),
.Y(n_1729)
);

OAI21xp5_ASAP7_75t_SL g1730 ( 
.A1(n_1697),
.A2(n_1572),
.B(n_1656),
.Y(n_1730)
);

OAI21xp33_ASAP7_75t_L g1731 ( 
.A1(n_1684),
.A2(n_1663),
.B(n_1697),
.Y(n_1731)
);

OAI22xp5_ASAP7_75t_L g1732 ( 
.A1(n_1663),
.A2(n_1585),
.B1(n_1646),
.B2(n_1601),
.Y(n_1732)
);

AND2x2_ASAP7_75t_L g1733 ( 
.A(n_1691),
.B(n_1692),
.Y(n_1733)
);

AND2x2_ASAP7_75t_L g1734 ( 
.A(n_1691),
.B(n_1596),
.Y(n_1734)
);

NAND2xp5_ASAP7_75t_L g1735 ( 
.A(n_1679),
.B(n_1598),
.Y(n_1735)
);

NAND2xp5_ASAP7_75t_L g1736 ( 
.A(n_1679),
.B(n_1598),
.Y(n_1736)
);

NAND2xp5_ASAP7_75t_L g1737 ( 
.A(n_1667),
.B(n_1597),
.Y(n_1737)
);

AND2x2_ASAP7_75t_L g1738 ( 
.A(n_1691),
.B(n_1596),
.Y(n_1738)
);

OAI21xp5_ASAP7_75t_SL g1739 ( 
.A1(n_1700),
.A2(n_1654),
.B(n_1629),
.Y(n_1739)
);

AND2x2_ASAP7_75t_L g1740 ( 
.A(n_1692),
.B(n_1677),
.Y(n_1740)
);

NAND3xp33_ASAP7_75t_L g1741 ( 
.A(n_1700),
.B(n_1650),
.C(n_1640),
.Y(n_1741)
);

OAI22xp5_ASAP7_75t_L g1742 ( 
.A1(n_1700),
.A2(n_1585),
.B1(n_1646),
.B2(n_1606),
.Y(n_1742)
);

AOI221x1_ASAP7_75t_SL g1743 ( 
.A1(n_1695),
.A2(n_1642),
.B1(n_1643),
.B2(n_1652),
.C(n_1645),
.Y(n_1743)
);

NAND2xp5_ASAP7_75t_L g1744 ( 
.A(n_1667),
.B(n_1604),
.Y(n_1744)
);

NAND2xp5_ASAP7_75t_L g1745 ( 
.A(n_1667),
.B(n_1690),
.Y(n_1745)
);

OAI21xp5_ASAP7_75t_L g1746 ( 
.A1(n_1702),
.A2(n_1641),
.B(n_1633),
.Y(n_1746)
);

AOI22xp5_ASAP7_75t_L g1747 ( 
.A1(n_1702),
.A2(n_1646),
.B1(n_1629),
.B2(n_1638),
.Y(n_1747)
);

AND2x2_ASAP7_75t_L g1748 ( 
.A(n_1692),
.B(n_1567),
.Y(n_1748)
);

OAI221xp5_ASAP7_75t_L g1749 ( 
.A1(n_1665),
.A2(n_1655),
.B1(n_1626),
.B2(n_1651),
.C(n_1650),
.Y(n_1749)
);

NAND2xp5_ASAP7_75t_SL g1750 ( 
.A(n_1681),
.B(n_1657),
.Y(n_1750)
);

AOI22xp33_ASAP7_75t_L g1751 ( 
.A1(n_1666),
.A2(n_1608),
.B1(n_1655),
.B2(n_1646),
.Y(n_1751)
);

OA21x2_ASAP7_75t_L g1752 ( 
.A1(n_1678),
.A2(n_1573),
.B(n_1592),
.Y(n_1752)
);

NAND2xp5_ASAP7_75t_L g1753 ( 
.A(n_1662),
.B(n_1645),
.Y(n_1753)
);

AND2x2_ASAP7_75t_L g1754 ( 
.A(n_1677),
.B(n_1567),
.Y(n_1754)
);

OAI21xp5_ASAP7_75t_SL g1755 ( 
.A1(n_1702),
.A2(n_1654),
.B(n_1609),
.Y(n_1755)
);

NAND3xp33_ASAP7_75t_L g1756 ( 
.A(n_1682),
.B(n_1640),
.C(n_1632),
.Y(n_1756)
);

NAND4xp25_ASAP7_75t_L g1757 ( 
.A(n_1696),
.B(n_1632),
.C(n_1637),
.D(n_1634),
.Y(n_1757)
);

AND2x2_ASAP7_75t_L g1758 ( 
.A(n_1733),
.B(n_1685),
.Y(n_1758)
);

INVx1_ASAP7_75t_L g1759 ( 
.A(n_1725),
.Y(n_1759)
);

AND2x2_ASAP7_75t_L g1760 ( 
.A(n_1733),
.B(n_1685),
.Y(n_1760)
);

NAND2xp5_ASAP7_75t_L g1761 ( 
.A(n_1743),
.B(n_1689),
.Y(n_1761)
);

INVx3_ASAP7_75t_L g1762 ( 
.A(n_1754),
.Y(n_1762)
);

INVx1_ASAP7_75t_L g1763 ( 
.A(n_1713),
.Y(n_1763)
);

OR2x2_ASAP7_75t_L g1764 ( 
.A(n_1713),
.B(n_1682),
.Y(n_1764)
);

INVx1_ASAP7_75t_L g1765 ( 
.A(n_1756),
.Y(n_1765)
);

INVx2_ASAP7_75t_L g1766 ( 
.A(n_1754),
.Y(n_1766)
);

INVx1_ASAP7_75t_L g1767 ( 
.A(n_1756),
.Y(n_1767)
);

INVx1_ASAP7_75t_L g1768 ( 
.A(n_1729),
.Y(n_1768)
);

AND2x4_ASAP7_75t_L g1769 ( 
.A(n_1734),
.B(n_1681),
.Y(n_1769)
);

NAND2xp5_ASAP7_75t_L g1770 ( 
.A(n_1720),
.B(n_1689),
.Y(n_1770)
);

OR2x2_ASAP7_75t_L g1771 ( 
.A(n_1745),
.B(n_1686),
.Y(n_1771)
);

AND2x2_ASAP7_75t_L g1772 ( 
.A(n_1740),
.B(n_1685),
.Y(n_1772)
);

BUFx3_ASAP7_75t_L g1773 ( 
.A(n_1749),
.Y(n_1773)
);

OR2x2_ASAP7_75t_L g1774 ( 
.A(n_1728),
.B(n_1686),
.Y(n_1774)
);

AND2x4_ASAP7_75t_L g1775 ( 
.A(n_1734),
.B(n_1681),
.Y(n_1775)
);

INVx1_ASAP7_75t_SL g1776 ( 
.A(n_1729),
.Y(n_1776)
);

INVx2_ASAP7_75t_L g1777 ( 
.A(n_1748),
.Y(n_1777)
);

NAND2xp5_ASAP7_75t_L g1778 ( 
.A(n_1720),
.B(n_1693),
.Y(n_1778)
);

AND2x4_ASAP7_75t_L g1779 ( 
.A(n_1738),
.B(n_1681),
.Y(n_1779)
);

AND2x2_ASAP7_75t_L g1780 ( 
.A(n_1748),
.B(n_1674),
.Y(n_1780)
);

INVx1_ASAP7_75t_L g1781 ( 
.A(n_1726),
.Y(n_1781)
);

AND2x2_ASAP7_75t_L g1782 ( 
.A(n_1738),
.B(n_1674),
.Y(n_1782)
);

NAND2xp5_ASAP7_75t_L g1783 ( 
.A(n_1718),
.B(n_1719),
.Y(n_1783)
);

INVx5_ASAP7_75t_L g1784 ( 
.A(n_1710),
.Y(n_1784)
);

INVx1_ASAP7_75t_L g1785 ( 
.A(n_1710),
.Y(n_1785)
);

AOI22xp5_ASAP7_75t_L g1786 ( 
.A1(n_1731),
.A2(n_1638),
.B1(n_1585),
.B2(n_1635),
.Y(n_1786)
);

NAND2xp5_ASAP7_75t_L g1787 ( 
.A(n_1718),
.B(n_1719),
.Y(n_1787)
);

AND2x4_ASAP7_75t_L g1788 ( 
.A(n_1750),
.B(n_1681),
.Y(n_1788)
);

INVx1_ASAP7_75t_L g1789 ( 
.A(n_1717),
.Y(n_1789)
);

INVx1_ASAP7_75t_L g1790 ( 
.A(n_1737),
.Y(n_1790)
);

INVx2_ASAP7_75t_L g1791 ( 
.A(n_1752),
.Y(n_1791)
);

NAND2xp5_ASAP7_75t_L g1792 ( 
.A(n_1708),
.B(n_1693),
.Y(n_1792)
);

INVx2_ASAP7_75t_L g1793 ( 
.A(n_1752),
.Y(n_1793)
);

INVx1_ASAP7_75t_SL g1794 ( 
.A(n_1707),
.Y(n_1794)
);

AND2x2_ASAP7_75t_L g1795 ( 
.A(n_1723),
.B(n_1698),
.Y(n_1795)
);

INVx1_ASAP7_75t_L g1796 ( 
.A(n_1744),
.Y(n_1796)
);

INVx1_ASAP7_75t_L g1797 ( 
.A(n_1763),
.Y(n_1797)
);

INVx1_ASAP7_75t_L g1798 ( 
.A(n_1763),
.Y(n_1798)
);

INVx2_ASAP7_75t_L g1799 ( 
.A(n_1777),
.Y(n_1799)
);

OR2x6_ASAP7_75t_L g1800 ( 
.A(n_1773),
.B(n_1687),
.Y(n_1800)
);

AND2x2_ASAP7_75t_L g1801 ( 
.A(n_1769),
.B(n_1708),
.Y(n_1801)
);

HB1xp67_ASAP7_75t_L g1802 ( 
.A(n_1759),
.Y(n_1802)
);

INVx1_ASAP7_75t_L g1803 ( 
.A(n_1768),
.Y(n_1803)
);

NAND2xp5_ASAP7_75t_SL g1804 ( 
.A(n_1773),
.B(n_1705),
.Y(n_1804)
);

INVx1_ASAP7_75t_L g1805 ( 
.A(n_1768),
.Y(n_1805)
);

NAND3xp33_ASAP7_75t_L g1806 ( 
.A(n_1786),
.B(n_1704),
.C(n_1705),
.Y(n_1806)
);

INVx2_ASAP7_75t_L g1807 ( 
.A(n_1777),
.Y(n_1807)
);

AND2x2_ASAP7_75t_L g1808 ( 
.A(n_1769),
.B(n_1747),
.Y(n_1808)
);

INVxp67_ASAP7_75t_SL g1809 ( 
.A(n_1761),
.Y(n_1809)
);

INVx1_ASAP7_75t_L g1810 ( 
.A(n_1792),
.Y(n_1810)
);

NAND2xp5_ASAP7_75t_L g1811 ( 
.A(n_1781),
.B(n_1716),
.Y(n_1811)
);

AND2x2_ASAP7_75t_L g1812 ( 
.A(n_1769),
.B(n_1747),
.Y(n_1812)
);

OR2x2_ASAP7_75t_L g1813 ( 
.A(n_1770),
.B(n_1711),
.Y(n_1813)
);

AND2x2_ASAP7_75t_L g1814 ( 
.A(n_1769),
.B(n_1694),
.Y(n_1814)
);

AND2x2_ASAP7_75t_L g1815 ( 
.A(n_1775),
.B(n_1694),
.Y(n_1815)
);

NAND3xp33_ASAP7_75t_L g1816 ( 
.A(n_1786),
.B(n_1715),
.C(n_1721),
.Y(n_1816)
);

NAND2xp5_ASAP7_75t_L g1817 ( 
.A(n_1781),
.B(n_1712),
.Y(n_1817)
);

INVx2_ASAP7_75t_SL g1818 ( 
.A(n_1784),
.Y(n_1818)
);

INVx1_ASAP7_75t_L g1819 ( 
.A(n_1792),
.Y(n_1819)
);

AND2x2_ASAP7_75t_L g1820 ( 
.A(n_1775),
.B(n_1746),
.Y(n_1820)
);

OR2x2_ASAP7_75t_L g1821 ( 
.A(n_1770),
.B(n_1753),
.Y(n_1821)
);

INVx1_ASAP7_75t_L g1822 ( 
.A(n_1759),
.Y(n_1822)
);

INVx2_ASAP7_75t_L g1823 ( 
.A(n_1777),
.Y(n_1823)
);

OAI21xp33_ASAP7_75t_L g1824 ( 
.A1(n_1773),
.A2(n_1731),
.B(n_1739),
.Y(n_1824)
);

INVx2_ASAP7_75t_L g1825 ( 
.A(n_1766),
.Y(n_1825)
);

INVx1_ASAP7_75t_L g1826 ( 
.A(n_1764),
.Y(n_1826)
);

OR2x2_ASAP7_75t_L g1827 ( 
.A(n_1778),
.B(n_1735),
.Y(n_1827)
);

OR2x2_ASAP7_75t_L g1828 ( 
.A(n_1778),
.B(n_1736),
.Y(n_1828)
);

NAND2xp5_ASAP7_75t_SL g1829 ( 
.A(n_1794),
.B(n_1721),
.Y(n_1829)
);

NAND2x1p5_ASAP7_75t_L g1830 ( 
.A(n_1784),
.B(n_1681),
.Y(n_1830)
);

NAND3xp33_ASAP7_75t_L g1831 ( 
.A(n_1765),
.B(n_1724),
.C(n_1706),
.Y(n_1831)
);

INVx1_ASAP7_75t_L g1832 ( 
.A(n_1764),
.Y(n_1832)
);

INVx1_ASAP7_75t_L g1833 ( 
.A(n_1761),
.Y(n_1833)
);

AND2x2_ASAP7_75t_SL g1834 ( 
.A(n_1765),
.B(n_1723),
.Y(n_1834)
);

AND2x2_ASAP7_75t_L g1835 ( 
.A(n_1775),
.B(n_1723),
.Y(n_1835)
);

INVx1_ASAP7_75t_L g1836 ( 
.A(n_1785),
.Y(n_1836)
);

AND2x2_ASAP7_75t_L g1837 ( 
.A(n_1775),
.B(n_1755),
.Y(n_1837)
);

OR2x6_ASAP7_75t_L g1838 ( 
.A(n_1795),
.B(n_1687),
.Y(n_1838)
);

OR2x2_ASAP7_75t_L g1839 ( 
.A(n_1771),
.B(n_1722),
.Y(n_1839)
);

AND2x2_ASAP7_75t_L g1840 ( 
.A(n_1779),
.B(n_1755),
.Y(n_1840)
);

NOR2x1_ASAP7_75t_L g1841 ( 
.A(n_1767),
.B(n_1741),
.Y(n_1841)
);

NOR2xp33_ASAP7_75t_L g1842 ( 
.A(n_1831),
.B(n_1794),
.Y(n_1842)
);

AND2x4_ASAP7_75t_L g1843 ( 
.A(n_1837),
.B(n_1784),
.Y(n_1843)
);

OR2x2_ASAP7_75t_L g1844 ( 
.A(n_1813),
.B(n_1783),
.Y(n_1844)
);

NOR2xp33_ASAP7_75t_L g1845 ( 
.A(n_1824),
.B(n_1730),
.Y(n_1845)
);

INVx1_ASAP7_75t_SL g1846 ( 
.A(n_1829),
.Y(n_1846)
);

OR2x2_ASAP7_75t_L g1847 ( 
.A(n_1813),
.B(n_1783),
.Y(n_1847)
);

NOR2xp33_ASAP7_75t_L g1848 ( 
.A(n_1804),
.B(n_1614),
.Y(n_1848)
);

AND2x2_ASAP7_75t_L g1849 ( 
.A(n_1837),
.B(n_1779),
.Y(n_1849)
);

NAND2xp5_ASAP7_75t_L g1850 ( 
.A(n_1809),
.B(n_1790),
.Y(n_1850)
);

INVx2_ASAP7_75t_L g1851 ( 
.A(n_1799),
.Y(n_1851)
);

INVx1_ASAP7_75t_L g1852 ( 
.A(n_1802),
.Y(n_1852)
);

AND2x2_ASAP7_75t_L g1853 ( 
.A(n_1840),
.B(n_1779),
.Y(n_1853)
);

INVx2_ASAP7_75t_SL g1854 ( 
.A(n_1801),
.Y(n_1854)
);

INVx1_ASAP7_75t_L g1855 ( 
.A(n_1822),
.Y(n_1855)
);

NAND2xp5_ASAP7_75t_L g1856 ( 
.A(n_1833),
.B(n_1790),
.Y(n_1856)
);

AND2x4_ASAP7_75t_L g1857 ( 
.A(n_1840),
.B(n_1784),
.Y(n_1857)
);

INVx2_ASAP7_75t_SL g1858 ( 
.A(n_1801),
.Y(n_1858)
);

HB1xp67_ASAP7_75t_L g1859 ( 
.A(n_1841),
.Y(n_1859)
);

AND2x2_ASAP7_75t_L g1860 ( 
.A(n_1808),
.B(n_1779),
.Y(n_1860)
);

AND2x2_ASAP7_75t_SL g1861 ( 
.A(n_1834),
.B(n_1767),
.Y(n_1861)
);

NAND2xp5_ASAP7_75t_L g1862 ( 
.A(n_1833),
.B(n_1796),
.Y(n_1862)
);

INVx1_ASAP7_75t_L g1863 ( 
.A(n_1797),
.Y(n_1863)
);

OAI211xp5_ASAP7_75t_L g1864 ( 
.A1(n_1816),
.A2(n_1709),
.B(n_1739),
.C(n_1795),
.Y(n_1864)
);

AOI21xp33_ASAP7_75t_SL g1865 ( 
.A1(n_1806),
.A2(n_1714),
.B(n_1727),
.Y(n_1865)
);

NAND2xp5_ASAP7_75t_L g1866 ( 
.A(n_1810),
.B(n_1796),
.Y(n_1866)
);

INVx1_ASAP7_75t_L g1867 ( 
.A(n_1797),
.Y(n_1867)
);

AOI22xp5_ASAP7_75t_L g1868 ( 
.A1(n_1834),
.A2(n_1732),
.B1(n_1742),
.B2(n_1703),
.Y(n_1868)
);

NAND2xp5_ASAP7_75t_L g1869 ( 
.A(n_1810),
.B(n_1819),
.Y(n_1869)
);

NOR2xp33_ASAP7_75t_L g1870 ( 
.A(n_1817),
.B(n_1614),
.Y(n_1870)
);

INVx2_ASAP7_75t_L g1871 ( 
.A(n_1799),
.Y(n_1871)
);

INVx1_ASAP7_75t_L g1872 ( 
.A(n_1798),
.Y(n_1872)
);

INVx1_ASAP7_75t_L g1873 ( 
.A(n_1798),
.Y(n_1873)
);

OR2x2_ASAP7_75t_L g1874 ( 
.A(n_1839),
.B(n_1787),
.Y(n_1874)
);

AOI221xp5_ASAP7_75t_L g1875 ( 
.A1(n_1819),
.A2(n_1795),
.B1(n_1782),
.B2(n_1780),
.C(n_1741),
.Y(n_1875)
);

INVx1_ASAP7_75t_L g1876 ( 
.A(n_1836),
.Y(n_1876)
);

INVx1_ASAP7_75t_L g1877 ( 
.A(n_1836),
.Y(n_1877)
);

NOR3x1_ASAP7_75t_L g1878 ( 
.A(n_1818),
.B(n_1757),
.C(n_1771),
.Y(n_1878)
);

OR2x2_ASAP7_75t_L g1879 ( 
.A(n_1839),
.B(n_1787),
.Y(n_1879)
);

INVx1_ASAP7_75t_L g1880 ( 
.A(n_1803),
.Y(n_1880)
);

NAND2xp5_ASAP7_75t_L g1881 ( 
.A(n_1811),
.B(n_1758),
.Y(n_1881)
);

INVxp67_ASAP7_75t_L g1882 ( 
.A(n_1800),
.Y(n_1882)
);

HB1xp67_ASAP7_75t_L g1883 ( 
.A(n_1803),
.Y(n_1883)
);

INVx2_ASAP7_75t_L g1884 ( 
.A(n_1807),
.Y(n_1884)
);

INVx1_ASAP7_75t_L g1885 ( 
.A(n_1805),
.Y(n_1885)
);

INVx1_ASAP7_75t_L g1886 ( 
.A(n_1805),
.Y(n_1886)
);

INVx1_ASAP7_75t_L g1887 ( 
.A(n_1826),
.Y(n_1887)
);

INVx1_ASAP7_75t_L g1888 ( 
.A(n_1883),
.Y(n_1888)
);

HB1xp67_ASAP7_75t_L g1889 ( 
.A(n_1859),
.Y(n_1889)
);

OR2x2_ASAP7_75t_L g1890 ( 
.A(n_1844),
.B(n_1847),
.Y(n_1890)
);

INVx1_ASAP7_75t_L g1891 ( 
.A(n_1883),
.Y(n_1891)
);

INVx1_ASAP7_75t_L g1892 ( 
.A(n_1876),
.Y(n_1892)
);

CKINVDCx16_ASAP7_75t_R g1893 ( 
.A(n_1859),
.Y(n_1893)
);

INVxp67_ASAP7_75t_L g1894 ( 
.A(n_1842),
.Y(n_1894)
);

INVx1_ASAP7_75t_SL g1895 ( 
.A(n_1846),
.Y(n_1895)
);

INVx1_ASAP7_75t_SL g1896 ( 
.A(n_1861),
.Y(n_1896)
);

OAI22xp5_ASAP7_75t_L g1897 ( 
.A1(n_1861),
.A2(n_1800),
.B1(n_1784),
.B2(n_1838),
.Y(n_1897)
);

INVxp67_ASAP7_75t_SL g1898 ( 
.A(n_1842),
.Y(n_1898)
);

AND2x2_ASAP7_75t_L g1899 ( 
.A(n_1860),
.B(n_1808),
.Y(n_1899)
);

OR2x2_ASAP7_75t_L g1900 ( 
.A(n_1874),
.B(n_1826),
.Y(n_1900)
);

INVxp67_ASAP7_75t_L g1901 ( 
.A(n_1845),
.Y(n_1901)
);

INVx3_ASAP7_75t_L g1902 ( 
.A(n_1843),
.Y(n_1902)
);

INVx2_ASAP7_75t_L g1903 ( 
.A(n_1851),
.Y(n_1903)
);

INVx1_ASAP7_75t_L g1904 ( 
.A(n_1877),
.Y(n_1904)
);

NAND2xp5_ASAP7_75t_L g1905 ( 
.A(n_1865),
.B(n_1827),
.Y(n_1905)
);

INVx1_ASAP7_75t_SL g1906 ( 
.A(n_1848),
.Y(n_1906)
);

INVx4_ASAP7_75t_L g1907 ( 
.A(n_1843),
.Y(n_1907)
);

INVx1_ASAP7_75t_L g1908 ( 
.A(n_1880),
.Y(n_1908)
);

INVx1_ASAP7_75t_SL g1909 ( 
.A(n_1848),
.Y(n_1909)
);

AND2x2_ASAP7_75t_L g1910 ( 
.A(n_1849),
.B(n_1812),
.Y(n_1910)
);

NAND2xp5_ASAP7_75t_L g1911 ( 
.A(n_1845),
.B(n_1827),
.Y(n_1911)
);

INVx1_ASAP7_75t_L g1912 ( 
.A(n_1885),
.Y(n_1912)
);

AOI222xp33_ASAP7_75t_SL g1913 ( 
.A1(n_1852),
.A2(n_1832),
.B1(n_1776),
.B2(n_1762),
.C1(n_1825),
.C2(n_1823),
.Y(n_1913)
);

BUFx2_ASAP7_75t_L g1914 ( 
.A(n_1843),
.Y(n_1914)
);

INVx2_ASAP7_75t_L g1915 ( 
.A(n_1851),
.Y(n_1915)
);

NOR3xp33_ASAP7_75t_L g1916 ( 
.A(n_1864),
.B(n_1474),
.C(n_1818),
.Y(n_1916)
);

AND2x4_ASAP7_75t_SL g1917 ( 
.A(n_1857),
.B(n_1800),
.Y(n_1917)
);

AND2x2_ASAP7_75t_L g1918 ( 
.A(n_1853),
.B(n_1812),
.Y(n_1918)
);

AND2x2_ASAP7_75t_L g1919 ( 
.A(n_1857),
.B(n_1835),
.Y(n_1919)
);

AND2x2_ASAP7_75t_L g1920 ( 
.A(n_1857),
.B(n_1835),
.Y(n_1920)
);

INVx2_ASAP7_75t_L g1921 ( 
.A(n_1871),
.Y(n_1921)
);

NOR2xp33_ASAP7_75t_L g1922 ( 
.A(n_1870),
.B(n_1625),
.Y(n_1922)
);

OAI221xp5_ASAP7_75t_L g1923 ( 
.A1(n_1868),
.A2(n_1800),
.B1(n_1830),
.B2(n_1838),
.C(n_1820),
.Y(n_1923)
);

OAI221xp5_ASAP7_75t_L g1924 ( 
.A1(n_1875),
.A2(n_1830),
.B1(n_1838),
.B2(n_1820),
.C(n_1832),
.Y(n_1924)
);

AND2x2_ASAP7_75t_L g1925 ( 
.A(n_1878),
.B(n_1814),
.Y(n_1925)
);

INVx1_ASAP7_75t_SL g1926 ( 
.A(n_1870),
.Y(n_1926)
);

OAI221xp5_ASAP7_75t_L g1927 ( 
.A1(n_1894),
.A2(n_1882),
.B1(n_1850),
.B2(n_1830),
.C(n_1858),
.Y(n_1927)
);

AOI22xp5_ASAP7_75t_L g1928 ( 
.A1(n_1898),
.A2(n_1882),
.B1(n_1854),
.B2(n_1838),
.Y(n_1928)
);

AND2x2_ASAP7_75t_L g1929 ( 
.A(n_1919),
.B(n_1814),
.Y(n_1929)
);

AOI31xp33_ASAP7_75t_L g1930 ( 
.A1(n_1896),
.A2(n_1625),
.A3(n_1432),
.B(n_1558),
.Y(n_1930)
);

HB1xp67_ASAP7_75t_L g1931 ( 
.A(n_1889),
.Y(n_1931)
);

AND2x2_ASAP7_75t_L g1932 ( 
.A(n_1919),
.B(n_1815),
.Y(n_1932)
);

AOI22xp5_ASAP7_75t_L g1933 ( 
.A1(n_1913),
.A2(n_1862),
.B1(n_1856),
.B2(n_1887),
.Y(n_1933)
);

INVx1_ASAP7_75t_L g1934 ( 
.A(n_1888),
.Y(n_1934)
);

OAI22xp5_ASAP7_75t_L g1935 ( 
.A1(n_1893),
.A2(n_1905),
.B1(n_1916),
.B2(n_1924),
.Y(n_1935)
);

NAND2xp5_ASAP7_75t_SL g1936 ( 
.A(n_1893),
.B(n_1784),
.Y(n_1936)
);

NAND2xp5_ASAP7_75t_L g1937 ( 
.A(n_1895),
.B(n_1855),
.Y(n_1937)
);

O2A1O1Ixp33_ASAP7_75t_L g1938 ( 
.A1(n_1901),
.A2(n_1869),
.B(n_1867),
.C(n_1863),
.Y(n_1938)
);

NAND2xp5_ASAP7_75t_L g1939 ( 
.A(n_1911),
.B(n_1881),
.Y(n_1939)
);

NAND3x2_ASAP7_75t_L g1940 ( 
.A(n_1914),
.B(n_1879),
.C(n_1815),
.Y(n_1940)
);

INVx1_ASAP7_75t_L g1941 ( 
.A(n_1888),
.Y(n_1941)
);

NAND2xp5_ASAP7_75t_L g1942 ( 
.A(n_1926),
.B(n_1866),
.Y(n_1942)
);

AOI21xp33_ASAP7_75t_L g1943 ( 
.A1(n_1906),
.A2(n_1873),
.B(n_1872),
.Y(n_1943)
);

OAI21xp5_ASAP7_75t_SL g1944 ( 
.A1(n_1909),
.A2(n_1751),
.B(n_1782),
.Y(n_1944)
);

OAI21xp5_ASAP7_75t_L g1945 ( 
.A1(n_1923),
.A2(n_1886),
.B(n_1884),
.Y(n_1945)
);

AOI22xp5_ASAP7_75t_L g1946 ( 
.A1(n_1925),
.A2(n_1782),
.B1(n_1788),
.B2(n_1780),
.Y(n_1946)
);

INVx1_ASAP7_75t_L g1947 ( 
.A(n_1891),
.Y(n_1947)
);

AOI22xp5_ASAP7_75t_L g1948 ( 
.A1(n_1925),
.A2(n_1788),
.B1(n_1780),
.B2(n_1681),
.Y(n_1948)
);

INVx1_ASAP7_75t_L g1949 ( 
.A(n_1891),
.Y(n_1949)
);

NAND2xp5_ASAP7_75t_L g1950 ( 
.A(n_1926),
.B(n_1828),
.Y(n_1950)
);

NAND2xp5_ASAP7_75t_L g1951 ( 
.A(n_1914),
.B(n_1828),
.Y(n_1951)
);

INVx1_ASAP7_75t_L g1952 ( 
.A(n_1892),
.Y(n_1952)
);

OAI33xp33_ASAP7_75t_L g1953 ( 
.A1(n_1892),
.A2(n_1912),
.A3(n_1908),
.B1(n_1904),
.B2(n_1897),
.B3(n_1900),
.Y(n_1953)
);

OAI322xp33_ASAP7_75t_L g1954 ( 
.A1(n_1900),
.A2(n_1884),
.A3(n_1871),
.B1(n_1791),
.B2(n_1793),
.C1(n_1821),
.C2(n_1774),
.Y(n_1954)
);

O2A1O1Ixp33_ASAP7_75t_SL g1955 ( 
.A1(n_1922),
.A2(n_1902),
.B(n_1908),
.C(n_1912),
.Y(n_1955)
);

AND2x4_ASAP7_75t_L g1956 ( 
.A(n_1931),
.B(n_1907),
.Y(n_1956)
);

INVx1_ASAP7_75t_L g1957 ( 
.A(n_1931),
.Y(n_1957)
);

BUFx4f_ASAP7_75t_SL g1958 ( 
.A(n_1936),
.Y(n_1958)
);

NOR2xp33_ASAP7_75t_L g1959 ( 
.A(n_1930),
.B(n_1907),
.Y(n_1959)
);

NAND2xp5_ASAP7_75t_L g1960 ( 
.A(n_1942),
.B(n_1910),
.Y(n_1960)
);

AND2x2_ASAP7_75t_L g1961 ( 
.A(n_1929),
.B(n_1920),
.Y(n_1961)
);

INVx1_ASAP7_75t_L g1962 ( 
.A(n_1952),
.Y(n_1962)
);

INVx1_ASAP7_75t_SL g1963 ( 
.A(n_1950),
.Y(n_1963)
);

INVx1_ASAP7_75t_L g1964 ( 
.A(n_1934),
.Y(n_1964)
);

INVx2_ASAP7_75t_L g1965 ( 
.A(n_1936),
.Y(n_1965)
);

NAND2xp5_ASAP7_75t_L g1966 ( 
.A(n_1937),
.B(n_1910),
.Y(n_1966)
);

NOR2x1p5_ASAP7_75t_SL g1967 ( 
.A(n_1941),
.B(n_1947),
.Y(n_1967)
);

INVx1_ASAP7_75t_L g1968 ( 
.A(n_1949),
.Y(n_1968)
);

INVx1_ASAP7_75t_L g1969 ( 
.A(n_1951),
.Y(n_1969)
);

OR2x2_ASAP7_75t_L g1970 ( 
.A(n_1939),
.B(n_1890),
.Y(n_1970)
);

NAND2xp5_ASAP7_75t_L g1971 ( 
.A(n_1933),
.B(n_1918),
.Y(n_1971)
);

INVx1_ASAP7_75t_L g1972 ( 
.A(n_1938),
.Y(n_1972)
);

INVx2_ASAP7_75t_L g1973 ( 
.A(n_1932),
.Y(n_1973)
);

AND2x2_ASAP7_75t_L g1974 ( 
.A(n_1945),
.B(n_1920),
.Y(n_1974)
);

OAI21xp33_ASAP7_75t_L g1975 ( 
.A1(n_1928),
.A2(n_1917),
.B(n_1890),
.Y(n_1975)
);

NAND2xp5_ASAP7_75t_L g1976 ( 
.A(n_1943),
.B(n_1918),
.Y(n_1976)
);

NAND2xp5_ASAP7_75t_L g1977 ( 
.A(n_1955),
.B(n_1899),
.Y(n_1977)
);

AND2x4_ASAP7_75t_SL g1978 ( 
.A(n_1948),
.B(n_1907),
.Y(n_1978)
);

OR2x2_ASAP7_75t_L g1979 ( 
.A(n_1940),
.B(n_1902),
.Y(n_1979)
);

INVx1_ASAP7_75t_L g1980 ( 
.A(n_1957),
.Y(n_1980)
);

OAI21xp33_ASAP7_75t_SL g1981 ( 
.A1(n_1977),
.A2(n_1935),
.B(n_1907),
.Y(n_1981)
);

NAND2xp5_ASAP7_75t_L g1982 ( 
.A(n_1956),
.B(n_1899),
.Y(n_1982)
);

AOI22xp5_ASAP7_75t_SL g1983 ( 
.A1(n_1972),
.A2(n_1959),
.B1(n_1956),
.B2(n_1963),
.Y(n_1983)
);

AOI22xp33_ASAP7_75t_L g1984 ( 
.A1(n_1959),
.A2(n_1953),
.B1(n_1927),
.B2(n_1917),
.Y(n_1984)
);

AOI221xp5_ASAP7_75t_L g1985 ( 
.A1(n_1971),
.A2(n_1953),
.B1(n_1954),
.B2(n_1944),
.C(n_1902),
.Y(n_1985)
);

OAI22xp5_ASAP7_75t_L g1986 ( 
.A1(n_1958),
.A2(n_1946),
.B1(n_1917),
.B2(n_1902),
.Y(n_1986)
);

OR2x2_ASAP7_75t_L g1987 ( 
.A(n_1966),
.B(n_1960),
.Y(n_1987)
);

INVx1_ASAP7_75t_L g1988 ( 
.A(n_1956),
.Y(n_1988)
);

NAND3xp33_ASAP7_75t_L g1989 ( 
.A(n_1965),
.B(n_1904),
.C(n_1903),
.Y(n_1989)
);

OAI221xp5_ASAP7_75t_L g1990 ( 
.A1(n_1975),
.A2(n_1921),
.B1(n_1915),
.B2(n_1903),
.C(n_1784),
.Y(n_1990)
);

AOI221x1_ASAP7_75t_L g1991 ( 
.A1(n_1964),
.A2(n_1968),
.B1(n_1962),
.B2(n_1965),
.C(n_1969),
.Y(n_1991)
);

NAND3xp33_ASAP7_75t_L g1992 ( 
.A(n_1979),
.B(n_1915),
.C(n_1903),
.Y(n_1992)
);

NOR2xp33_ASAP7_75t_L g1993 ( 
.A(n_1981),
.B(n_1970),
.Y(n_1993)
);

AOI22xp5_ASAP7_75t_L g1994 ( 
.A1(n_1985),
.A2(n_1974),
.B1(n_1973),
.B2(n_1961),
.Y(n_1994)
);

NOR4xp25_ASAP7_75t_L g1995 ( 
.A(n_1988),
.B(n_1967),
.C(n_1976),
.D(n_1974),
.Y(n_1995)
);

NAND2xp5_ASAP7_75t_L g1996 ( 
.A(n_1983),
.B(n_1973),
.Y(n_1996)
);

NOR2x1p5_ASAP7_75t_L g1997 ( 
.A(n_1982),
.B(n_1569),
.Y(n_1997)
);

AND4x1_ASAP7_75t_L g1998 ( 
.A(n_1984),
.B(n_1961),
.C(n_1566),
.D(n_1958),
.Y(n_1998)
);

INVxp67_ASAP7_75t_L g1999 ( 
.A(n_1987),
.Y(n_1999)
);

AND5x1_ASAP7_75t_L g2000 ( 
.A(n_1986),
.B(n_1978),
.C(n_1921),
.D(n_1915),
.E(n_1566),
.Y(n_2000)
);

NOR2x1_ASAP7_75t_L g2001 ( 
.A(n_1989),
.B(n_1992),
.Y(n_2001)
);

NOR2xp33_ASAP7_75t_L g2002 ( 
.A(n_1980),
.B(n_1978),
.Y(n_2002)
);

AOI211xp5_ASAP7_75t_L g2003 ( 
.A1(n_1990),
.A2(n_1921),
.B(n_1437),
.C(n_1788),
.Y(n_2003)
);

NAND4xp25_ASAP7_75t_L g2004 ( 
.A(n_1994),
.B(n_1993),
.C(n_2002),
.D(n_2003),
.Y(n_2004)
);

AOI221xp5_ASAP7_75t_L g2005 ( 
.A1(n_1995),
.A2(n_1991),
.B1(n_1793),
.B2(n_1791),
.C(n_1788),
.Y(n_2005)
);

INVx1_ASAP7_75t_L g2006 ( 
.A(n_1996),
.Y(n_2006)
);

AOI211xp5_ASAP7_75t_L g2007 ( 
.A1(n_1999),
.A2(n_1554),
.B(n_1505),
.C(n_1549),
.Y(n_2007)
);

NAND2xp5_ASAP7_75t_SL g2008 ( 
.A(n_2001),
.B(n_1444),
.Y(n_2008)
);

NOR3xp33_ASAP7_75t_L g2009 ( 
.A(n_1998),
.B(n_1524),
.C(n_1520),
.Y(n_2009)
);

NOR3xp33_ASAP7_75t_SL g2010 ( 
.A(n_2000),
.B(n_1997),
.C(n_1454),
.Y(n_2010)
);

NAND2xp5_ASAP7_75t_L g2011 ( 
.A(n_2006),
.B(n_1821),
.Y(n_2011)
);

INVxp67_ASAP7_75t_L g2012 ( 
.A(n_2008),
.Y(n_2012)
);

INVx2_ASAP7_75t_L g2013 ( 
.A(n_2009),
.Y(n_2013)
);

NAND2xp5_ASAP7_75t_L g2014 ( 
.A(n_2004),
.B(n_2007),
.Y(n_2014)
);

INVx1_ASAP7_75t_L g2015 ( 
.A(n_2010),
.Y(n_2015)
);

NOR2x1_ASAP7_75t_L g2016 ( 
.A(n_2005),
.B(n_1473),
.Y(n_2016)
);

INVx1_ASAP7_75t_L g2017 ( 
.A(n_2006),
.Y(n_2017)
);

NOR2x1_ASAP7_75t_L g2018 ( 
.A(n_2017),
.B(n_1473),
.Y(n_2018)
);

NOR3x2_ASAP7_75t_L g2019 ( 
.A(n_2015),
.B(n_1476),
.C(n_1549),
.Y(n_2019)
);

NOR3xp33_ASAP7_75t_L g2020 ( 
.A(n_2013),
.B(n_1476),
.C(n_1554),
.Y(n_2020)
);

INVx2_ASAP7_75t_L g2021 ( 
.A(n_2012),
.Y(n_2021)
);

INVx1_ASAP7_75t_L g2022 ( 
.A(n_2011),
.Y(n_2022)
);

OAI221xp5_ASAP7_75t_L g2023 ( 
.A1(n_2016),
.A2(n_1825),
.B1(n_1823),
.B2(n_1807),
.C(n_1631),
.Y(n_2023)
);

NOR3xp33_ASAP7_75t_SL g2024 ( 
.A(n_2022),
.B(n_2014),
.C(n_1554),
.Y(n_2024)
);

BUFx2_ASAP7_75t_L g2025 ( 
.A(n_2018),
.Y(n_2025)
);

INVx2_ASAP7_75t_L g2026 ( 
.A(n_2019),
.Y(n_2026)
);

XNOR2xp5_ASAP7_75t_L g2027 ( 
.A(n_2021),
.B(n_1522),
.Y(n_2027)
);

XNOR2x1_ASAP7_75t_L g2028 ( 
.A(n_2027),
.B(n_2020),
.Y(n_2028)
);

INVx2_ASAP7_75t_L g2029 ( 
.A(n_2028),
.Y(n_2029)
);

AOI221x1_ASAP7_75t_L g2030 ( 
.A1(n_2029),
.A2(n_2026),
.B1(n_2024),
.B2(n_2025),
.C(n_2023),
.Y(n_2030)
);

OAI22xp5_ASAP7_75t_L g2031 ( 
.A1(n_2029),
.A2(n_2024),
.B1(n_1762),
.B2(n_1791),
.Y(n_2031)
);

NAND2xp5_ASAP7_75t_L g2032 ( 
.A(n_2030),
.B(n_1647),
.Y(n_2032)
);

OAI22xp5_ASAP7_75t_L g2033 ( 
.A1(n_2031),
.A2(n_1762),
.B1(n_1793),
.B2(n_1774),
.Y(n_2033)
);

AOI21xp33_ASAP7_75t_L g2034 ( 
.A1(n_2032),
.A2(n_1659),
.B(n_1647),
.Y(n_2034)
);

AOI222xp33_ASAP7_75t_L g2035 ( 
.A1(n_2033),
.A2(n_1520),
.B1(n_1524),
.B2(n_1760),
.C1(n_1758),
.C2(n_1772),
.Y(n_2035)
);

NAND3xp33_ASAP7_75t_L g2036 ( 
.A(n_2034),
.B(n_1659),
.C(n_1606),
.Y(n_2036)
);

INVx1_ASAP7_75t_L g2037 ( 
.A(n_2036),
.Y(n_2037)
);

AOI221xp5_ASAP7_75t_L g2038 ( 
.A1(n_2037),
.A2(n_2035),
.B1(n_1762),
.B2(n_1672),
.C(n_1789),
.Y(n_2038)
);

AOI211xp5_ASAP7_75t_L g2039 ( 
.A1(n_2038),
.A2(n_1601),
.B(n_1606),
.C(n_1657),
.Y(n_2039)
);


endmodule