module fake_jpeg_22515_n_4 (n_0, n_1, n_4);

input n_0;
input n_1;

output n_4;

wire n_3;
wire n_2;

CKINVDCx20_ASAP7_75t_R g2 ( 
.A(n_1),
.Y(n_2)
);

XNOR2xp5_ASAP7_75t_L g3 ( 
.A(n_0),
.B(n_1),
.Y(n_3)
);

AOI322xp5_ASAP7_75t_L g4 ( 
.A1(n_3),
.A2(n_0),
.A3(n_1),
.B1(n_2),
.B2(n_0),
.C1(n_1),
.C2(n_2),
.Y(n_4)
);


endmodule