module fake_jpeg_12320_n_114 (n_13, n_21, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_19, n_18, n_20, n_4, n_30, n_16, n_3, n_0, n_24, n_28, n_26, n_9, n_5, n_11, n_17, n_25, n_31, n_2, n_29, n_12, n_8, n_15, n_7, n_114);

input n_13;
input n_21;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_4;
input n_30;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_26;
input n_9;
input n_5;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_12;
input n_8;
input n_15;
input n_7;

output n_114;

wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_73;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_42;
wire n_49;
wire n_76;
wire n_38;
wire n_88;
wire n_74;
wire n_103;
wire n_50;
wire n_57;
wire n_69;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_109;
wire n_113;
wire n_106;
wire n_111;
wire n_44;
wire n_75;
wire n_37;
wire n_102;
wire n_99;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_56;
wire n_79;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_101;
wire n_48;
wire n_35;
wire n_87;
wire n_46;
wire n_86;
wire n_112;
wire n_95;
wire n_97;
wire n_36;
wire n_62;
wire n_43;
wire n_32;
wire n_100;
wire n_82;
wire n_96;

INVx1_ASAP7_75t_L g32 ( 
.A(n_21),
.Y(n_32)
);

INVx3_ASAP7_75t_L g33 ( 
.A(n_25),
.Y(n_33)
);

NAND2xp5_ASAP7_75t_L g34 ( 
.A(n_30),
.B(n_17),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_8),
.Y(n_35)
);

BUFx12_ASAP7_75t_L g36 ( 
.A(n_1),
.Y(n_36)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_3),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_26),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_19),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_5),
.Y(n_40)
);

BUFx12f_ASAP7_75t_L g41 ( 
.A(n_24),
.Y(n_41)
);

CKINVDCx14_ASAP7_75t_R g42 ( 
.A(n_29),
.Y(n_42)
);

BUFx12f_ASAP7_75t_L g43 ( 
.A(n_0),
.Y(n_43)
);

INVx13_ASAP7_75t_L g44 ( 
.A(n_4),
.Y(n_44)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_4),
.Y(n_45)
);

BUFx3_ASAP7_75t_L g46 ( 
.A(n_41),
.Y(n_46)
);

INVx5_ASAP7_75t_L g62 ( 
.A(n_46),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g47 ( 
.A(n_40),
.B(n_0),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_47),
.B(n_52),
.Y(n_56)
);

INVx5_ASAP7_75t_L g48 ( 
.A(n_41),
.Y(n_48)
);

INVx5_ASAP7_75t_L g67 ( 
.A(n_48),
.Y(n_67)
);

BUFx12f_ASAP7_75t_L g49 ( 
.A(n_35),
.Y(n_49)
);

INVx3_ASAP7_75t_L g66 ( 
.A(n_49),
.Y(n_66)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_37),
.Y(n_50)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_50),
.Y(n_61)
);

INVx2_ASAP7_75t_L g51 ( 
.A(n_43),
.Y(n_51)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_51),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_34),
.B(n_1),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_38),
.B(n_2),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g57 ( 
.A(n_53),
.B(n_42),
.Y(n_57)
);

INVx3_ASAP7_75t_L g54 ( 
.A(n_43),
.Y(n_54)
);

INVx6_ASAP7_75t_L g64 ( 
.A(n_54),
.Y(n_64)
);

AO21x1_ASAP7_75t_L g55 ( 
.A1(n_47),
.A2(n_45),
.B(n_42),
.Y(n_55)
);

AOI21xp5_ASAP7_75t_L g81 ( 
.A1(n_55),
.A2(n_60),
.B(n_6),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_57),
.B(n_59),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_52),
.B(n_49),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_L g71 ( 
.A(n_58),
.B(n_65),
.Y(n_71)
);

CKINVDCx16_ASAP7_75t_R g59 ( 
.A(n_48),
.Y(n_59)
);

AOI22xp5_ASAP7_75t_SL g60 ( 
.A1(n_51),
.A2(n_41),
.B1(n_44),
.B2(n_33),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_L g65 ( 
.A(n_52),
.B(n_39),
.Y(n_65)
);

CKINVDCx20_ASAP7_75t_R g68 ( 
.A(n_61),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_68),
.B(n_70),
.Y(n_85)
);

MAJIxp5_ASAP7_75t_L g69 ( 
.A(n_63),
.B(n_32),
.C(n_44),
.Y(n_69)
);

MAJIxp5_ASAP7_75t_L g92 ( 
.A(n_69),
.B(n_75),
.C(n_76),
.Y(n_92)
);

CKINVDCx20_ASAP7_75t_R g70 ( 
.A(n_66),
.Y(n_70)
);

CKINVDCx20_ASAP7_75t_R g73 ( 
.A(n_66),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_73),
.B(n_74),
.Y(n_88)
);

CKINVDCx20_ASAP7_75t_R g74 ( 
.A(n_64),
.Y(n_74)
);

MAJIxp5_ASAP7_75t_L g75 ( 
.A(n_56),
.B(n_36),
.C(n_15),
.Y(n_75)
);

MAJx2_ASAP7_75t_L g76 ( 
.A(n_55),
.B(n_14),
.C(n_31),
.Y(n_76)
);

INVxp67_ASAP7_75t_L g77 ( 
.A(n_62),
.Y(n_77)
);

HB1xp67_ASAP7_75t_L g84 ( 
.A(n_77),
.Y(n_84)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_67),
.Y(n_78)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_78),
.Y(n_83)
);

CKINVDCx20_ASAP7_75t_R g79 ( 
.A(n_67),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_79),
.B(n_22),
.Y(n_95)
);

BUFx12_ASAP7_75t_L g80 ( 
.A(n_59),
.Y(n_80)
);

CKINVDCx20_ASAP7_75t_R g82 ( 
.A(n_80),
.Y(n_82)
);

INVxp67_ASAP7_75t_L g89 ( 
.A(n_81),
.Y(n_89)
);

OR2x2_ASAP7_75t_L g86 ( 
.A(n_69),
.B(n_7),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_SL g100 ( 
.A(n_86),
.B(n_87),
.Y(n_100)
);

OAI22xp5_ASAP7_75t_SL g87 ( 
.A1(n_72),
.A2(n_9),
.B1(n_10),
.B2(n_11),
.Y(n_87)
);

XNOR2xp5_ASAP7_75t_SL g90 ( 
.A(n_71),
.B(n_12),
.Y(n_90)
);

MAJIxp5_ASAP7_75t_L g97 ( 
.A(n_90),
.B(n_94),
.C(n_23),
.Y(n_97)
);

OAI22xp5_ASAP7_75t_L g91 ( 
.A1(n_76),
.A2(n_13),
.B1(n_16),
.B2(n_18),
.Y(n_91)
);

AND2x2_ASAP7_75t_L g102 ( 
.A(n_91),
.B(n_95),
.Y(n_102)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_80),
.Y(n_93)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_93),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_SL g94 ( 
.A(n_71),
.B(n_20),
.Y(n_94)
);

XNOR2xp5_ASAP7_75t_L g106 ( 
.A(n_97),
.B(n_98),
.Y(n_106)
);

MAJIxp5_ASAP7_75t_L g98 ( 
.A(n_92),
.B(n_86),
.C(n_85),
.Y(n_98)
);

MAJIxp5_ASAP7_75t_L g99 ( 
.A(n_82),
.B(n_27),
.C(n_28),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_99),
.B(n_103),
.Y(n_105)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_88),
.Y(n_101)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_101),
.Y(n_107)
);

CKINVDCx20_ASAP7_75t_R g103 ( 
.A(n_84),
.Y(n_103)
);

OAI21xp5_ASAP7_75t_L g104 ( 
.A1(n_96),
.A2(n_89),
.B(n_83),
.Y(n_104)
);

XNOR2xp5_ASAP7_75t_L g108 ( 
.A(n_104),
.B(n_84),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_SL g110 ( 
.A(n_108),
.B(n_109),
.Y(n_110)
);

OAI21xp5_ASAP7_75t_SL g109 ( 
.A1(n_107),
.A2(n_100),
.B(n_102),
.Y(n_109)
);

XNOR2xp5_ASAP7_75t_L g111 ( 
.A(n_110),
.B(n_106),
.Y(n_111)
);

XNOR2xp5_ASAP7_75t_L g112 ( 
.A(n_111),
.B(n_105),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_SL g113 ( 
.A(n_112),
.B(n_105),
.Y(n_113)
);

XNOR2xp5_ASAP7_75t_L g114 ( 
.A(n_113),
.B(n_100),
.Y(n_114)
);


endmodule