module fake_netlist_1_1492_n_17 (n_1, n_2, n_0, n_17);
input n_1;
input n_2;
input n_0;
output n_17;
wire n_11;
wire n_13;
wire n_16;
wire n_12;
wire n_6;
wire n_4;
wire n_3;
wire n_9;
wire n_5;
wire n_14;
wire n_7;
wire n_15;
wire n_10;
wire n_8;
INVx2_ASAP7_75t_L g3 ( .A(n_2), .Y(n_3) );
INVx2_ASAP7_75t_L g4 ( .A(n_2), .Y(n_4) );
INVx5_ASAP7_75t_L g5 ( .A(n_2), .Y(n_5) );
INVx2_ASAP7_75t_SL g6 ( .A(n_5), .Y(n_6) );
AND2x4_ASAP7_75t_L g7 ( .A(n_5), .B(n_0), .Y(n_7) );
BUFx2_ASAP7_75t_L g8 ( .A(n_7), .Y(n_8) );
NAND2xp5_ASAP7_75t_L g9 ( .A(n_6), .B(n_3), .Y(n_9) );
OR2x2_ASAP7_75t_L g10 ( .A(n_9), .B(n_7), .Y(n_10) );
INVx1_ASAP7_75t_L g11 ( .A(n_8), .Y(n_11) );
INVxp67_ASAP7_75t_L g12 ( .A(n_10), .Y(n_12) );
OAI322xp33_ASAP7_75t_L g13 ( .A1(n_11), .A2(n_0), .A3(n_1), .B1(n_4), .B2(n_6), .C1(n_7), .C2(n_9), .Y(n_13) );
INVx1_ASAP7_75t_L g14 ( .A(n_13), .Y(n_14) );
NOR4xp25_ASAP7_75t_L g15 ( .A(n_12), .B(n_0), .C(n_1), .D(n_7), .Y(n_15) );
INVx1_ASAP7_75t_L g16 ( .A(n_14), .Y(n_16) );
OAI21xp5_ASAP7_75t_L g17 ( .A1(n_16), .A2(n_15), .B(n_14), .Y(n_17) );
endmodule