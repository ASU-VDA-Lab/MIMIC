module fake_netlist_6_1050_n_2086 (n_52, n_435, n_1, n_91, n_326, n_256, n_440, n_507, n_209, n_367, n_465, n_63, n_223, n_278, n_341, n_362, n_148, n_226, n_161, n_22, n_208, n_462, n_68, n_316, n_419, n_28, n_304, n_212, n_50, n_7, n_144, n_365, n_125, n_168, n_384, n_297, n_342, n_77, n_106, n_358, n_160, n_449, n_131, n_188, n_310, n_509, n_186, n_245, n_0, n_368, n_396, n_495, n_350, n_78, n_84, n_392, n_442, n_480, n_142, n_143, n_382, n_180, n_62, n_349, n_233, n_255, n_284, n_400, n_140, n_337, n_214, n_485, n_67, n_15, n_443, n_246, n_38, n_471, n_289, n_421, n_424, n_59, n_181, n_182, n_238, n_202, n_320, n_108, n_327, n_369, n_280, n_287, n_353, n_389, n_415, n_65, n_230, n_461, n_141, n_383, n_200, n_447, n_176, n_114, n_86, n_198, n_104, n_222, n_179, n_248, n_300, n_71, n_74, n_229, n_305, n_72, n_173, n_250, n_372, n_468, n_111, n_504, n_314, n_378, n_413, n_377, n_35, n_183, n_510, n_79, n_375, n_338, n_466, n_506, n_56, n_360, n_119, n_235, n_147, n_191, n_340, n_387, n_452, n_39, n_344, n_73, n_428, n_432, n_101, n_167, n_174, n_127, n_153, n_156, n_491, n_145, n_42, n_133, n_96, n_8, n_371, n_189, n_405, n_213, n_294, n_302, n_499, n_380, n_129, n_197, n_11, n_137, n_17, n_343, n_448, n_20, n_494, n_493, n_397, n_155, n_109, n_445, n_425, n_122, n_45, n_454, n_34, n_218, n_70, n_234, n_37, n_486, n_381, n_82, n_27, n_236, n_112, n_172, n_472, n_270, n_239, n_126, n_414, n_97, n_58, n_490, n_290, n_220, n_118, n_224, n_48, n_25, n_93, n_80, n_196, n_402, n_352, n_478, n_9, n_460, n_107, n_6, n_417, n_14, n_446, n_498, n_89, n_374, n_366, n_407, n_450, n_103, n_272, n_185, n_348, n_69, n_376, n_390, n_473, n_293, n_31, n_334, n_53, n_370, n_44, n_458, n_232, n_16, n_163, n_46, n_330, n_470, n_475, n_298, n_18, n_492, n_281, n_258, n_154, n_456, n_98, n_260, n_265, n_313, n_451, n_279, n_252, n_228, n_356, n_166, n_184, n_216, n_455, n_83, n_363, n_395, n_323, n_393, n_411, n_503, n_152, n_92, n_513, n_321, n_331, n_105, n_227, n_132, n_406, n_483, n_102, n_204, n_482, n_474, n_261, n_420, n_312, n_394, n_32, n_66, n_130, n_512, n_164, n_292, n_100, n_121, n_307, n_469, n_433, n_500, n_23, n_476, n_2, n_291, n_219, n_357, n_150, n_264, n_263, n_481, n_325, n_329, n_464, n_33, n_477, n_408, n_61, n_237, n_244, n_399, n_76, n_243, n_124, n_94, n_282, n_436, n_116, n_211, n_117, n_175, n_322, n_345, n_409, n_231, n_354, n_40, n_505, n_240, n_139, n_319, n_41, n_134, n_273, n_95, n_311, n_10, n_403, n_253, n_123, n_136, n_249, n_201, n_386, n_159, n_157, n_162, n_115, n_487, n_128, n_241, n_30, n_275, n_43, n_276, n_441, n_221, n_444, n_423, n_146, n_318, n_303, n_511, n_467, n_306, n_21, n_193, n_269, n_359, n_346, n_88, n_3, n_416, n_277, n_418, n_113, n_4, n_199, n_138, n_266, n_296, n_268, n_271, n_404, n_439, n_158, n_217, n_49, n_210, n_299, n_206, n_5, n_453, n_333, n_215, n_178, n_247, n_225, n_308, n_309, n_355, n_426, n_317, n_149, n_431, n_90, n_347, n_24, n_459, n_54, n_502, n_328, n_488, n_429, n_373, n_87, n_195, n_285, n_497, n_85, n_99, n_257, n_13, n_203, n_286, n_254, n_207, n_242, n_19, n_47, n_29, n_75, n_401, n_324, n_335, n_430, n_463, n_489, n_205, n_120, n_251, n_301, n_274, n_110, n_151, n_412, n_81, n_36, n_26, n_55, n_267, n_438, n_339, n_315, n_434, n_515, n_64, n_288, n_427, n_479, n_496, n_422, n_135, n_165, n_351, n_437, n_259, n_177, n_514, n_391, n_457, n_364, n_295, n_385, n_388, n_190, n_262, n_484, n_187, n_501, n_60, n_361, n_508, n_379, n_170, n_332, n_336, n_12, n_398, n_410, n_194, n_171, n_192, n_57, n_169, n_51, n_283, n_2086);

input n_52;
input n_435;
input n_1;
input n_91;
input n_326;
input n_256;
input n_440;
input n_507;
input n_209;
input n_367;
input n_465;
input n_63;
input n_223;
input n_278;
input n_341;
input n_362;
input n_148;
input n_226;
input n_161;
input n_22;
input n_208;
input n_462;
input n_68;
input n_316;
input n_419;
input n_28;
input n_304;
input n_212;
input n_50;
input n_7;
input n_144;
input n_365;
input n_125;
input n_168;
input n_384;
input n_297;
input n_342;
input n_77;
input n_106;
input n_358;
input n_160;
input n_449;
input n_131;
input n_188;
input n_310;
input n_509;
input n_186;
input n_245;
input n_0;
input n_368;
input n_396;
input n_495;
input n_350;
input n_78;
input n_84;
input n_392;
input n_442;
input n_480;
input n_142;
input n_143;
input n_382;
input n_180;
input n_62;
input n_349;
input n_233;
input n_255;
input n_284;
input n_400;
input n_140;
input n_337;
input n_214;
input n_485;
input n_67;
input n_15;
input n_443;
input n_246;
input n_38;
input n_471;
input n_289;
input n_421;
input n_424;
input n_59;
input n_181;
input n_182;
input n_238;
input n_202;
input n_320;
input n_108;
input n_327;
input n_369;
input n_280;
input n_287;
input n_353;
input n_389;
input n_415;
input n_65;
input n_230;
input n_461;
input n_141;
input n_383;
input n_200;
input n_447;
input n_176;
input n_114;
input n_86;
input n_198;
input n_104;
input n_222;
input n_179;
input n_248;
input n_300;
input n_71;
input n_74;
input n_229;
input n_305;
input n_72;
input n_173;
input n_250;
input n_372;
input n_468;
input n_111;
input n_504;
input n_314;
input n_378;
input n_413;
input n_377;
input n_35;
input n_183;
input n_510;
input n_79;
input n_375;
input n_338;
input n_466;
input n_506;
input n_56;
input n_360;
input n_119;
input n_235;
input n_147;
input n_191;
input n_340;
input n_387;
input n_452;
input n_39;
input n_344;
input n_73;
input n_428;
input n_432;
input n_101;
input n_167;
input n_174;
input n_127;
input n_153;
input n_156;
input n_491;
input n_145;
input n_42;
input n_133;
input n_96;
input n_8;
input n_371;
input n_189;
input n_405;
input n_213;
input n_294;
input n_302;
input n_499;
input n_380;
input n_129;
input n_197;
input n_11;
input n_137;
input n_17;
input n_343;
input n_448;
input n_20;
input n_494;
input n_493;
input n_397;
input n_155;
input n_109;
input n_445;
input n_425;
input n_122;
input n_45;
input n_454;
input n_34;
input n_218;
input n_70;
input n_234;
input n_37;
input n_486;
input n_381;
input n_82;
input n_27;
input n_236;
input n_112;
input n_172;
input n_472;
input n_270;
input n_239;
input n_126;
input n_414;
input n_97;
input n_58;
input n_490;
input n_290;
input n_220;
input n_118;
input n_224;
input n_48;
input n_25;
input n_93;
input n_80;
input n_196;
input n_402;
input n_352;
input n_478;
input n_9;
input n_460;
input n_107;
input n_6;
input n_417;
input n_14;
input n_446;
input n_498;
input n_89;
input n_374;
input n_366;
input n_407;
input n_450;
input n_103;
input n_272;
input n_185;
input n_348;
input n_69;
input n_376;
input n_390;
input n_473;
input n_293;
input n_31;
input n_334;
input n_53;
input n_370;
input n_44;
input n_458;
input n_232;
input n_16;
input n_163;
input n_46;
input n_330;
input n_470;
input n_475;
input n_298;
input n_18;
input n_492;
input n_281;
input n_258;
input n_154;
input n_456;
input n_98;
input n_260;
input n_265;
input n_313;
input n_451;
input n_279;
input n_252;
input n_228;
input n_356;
input n_166;
input n_184;
input n_216;
input n_455;
input n_83;
input n_363;
input n_395;
input n_323;
input n_393;
input n_411;
input n_503;
input n_152;
input n_92;
input n_513;
input n_321;
input n_331;
input n_105;
input n_227;
input n_132;
input n_406;
input n_483;
input n_102;
input n_204;
input n_482;
input n_474;
input n_261;
input n_420;
input n_312;
input n_394;
input n_32;
input n_66;
input n_130;
input n_512;
input n_164;
input n_292;
input n_100;
input n_121;
input n_307;
input n_469;
input n_433;
input n_500;
input n_23;
input n_476;
input n_2;
input n_291;
input n_219;
input n_357;
input n_150;
input n_264;
input n_263;
input n_481;
input n_325;
input n_329;
input n_464;
input n_33;
input n_477;
input n_408;
input n_61;
input n_237;
input n_244;
input n_399;
input n_76;
input n_243;
input n_124;
input n_94;
input n_282;
input n_436;
input n_116;
input n_211;
input n_117;
input n_175;
input n_322;
input n_345;
input n_409;
input n_231;
input n_354;
input n_40;
input n_505;
input n_240;
input n_139;
input n_319;
input n_41;
input n_134;
input n_273;
input n_95;
input n_311;
input n_10;
input n_403;
input n_253;
input n_123;
input n_136;
input n_249;
input n_201;
input n_386;
input n_159;
input n_157;
input n_162;
input n_115;
input n_487;
input n_128;
input n_241;
input n_30;
input n_275;
input n_43;
input n_276;
input n_441;
input n_221;
input n_444;
input n_423;
input n_146;
input n_318;
input n_303;
input n_511;
input n_467;
input n_306;
input n_21;
input n_193;
input n_269;
input n_359;
input n_346;
input n_88;
input n_3;
input n_416;
input n_277;
input n_418;
input n_113;
input n_4;
input n_199;
input n_138;
input n_266;
input n_296;
input n_268;
input n_271;
input n_404;
input n_439;
input n_158;
input n_217;
input n_49;
input n_210;
input n_299;
input n_206;
input n_5;
input n_453;
input n_333;
input n_215;
input n_178;
input n_247;
input n_225;
input n_308;
input n_309;
input n_355;
input n_426;
input n_317;
input n_149;
input n_431;
input n_90;
input n_347;
input n_24;
input n_459;
input n_54;
input n_502;
input n_328;
input n_488;
input n_429;
input n_373;
input n_87;
input n_195;
input n_285;
input n_497;
input n_85;
input n_99;
input n_257;
input n_13;
input n_203;
input n_286;
input n_254;
input n_207;
input n_242;
input n_19;
input n_47;
input n_29;
input n_75;
input n_401;
input n_324;
input n_335;
input n_430;
input n_463;
input n_489;
input n_205;
input n_120;
input n_251;
input n_301;
input n_274;
input n_110;
input n_151;
input n_412;
input n_81;
input n_36;
input n_26;
input n_55;
input n_267;
input n_438;
input n_339;
input n_315;
input n_434;
input n_515;
input n_64;
input n_288;
input n_427;
input n_479;
input n_496;
input n_422;
input n_135;
input n_165;
input n_351;
input n_437;
input n_259;
input n_177;
input n_514;
input n_391;
input n_457;
input n_364;
input n_295;
input n_385;
input n_388;
input n_190;
input n_262;
input n_484;
input n_187;
input n_501;
input n_60;
input n_361;
input n_508;
input n_379;
input n_170;
input n_332;
input n_336;
input n_12;
input n_398;
input n_410;
input n_194;
input n_171;
input n_192;
input n_57;
input n_169;
input n_51;
input n_283;

output n_2086;

wire n_992;
wire n_1671;
wire n_801;
wire n_1613;
wire n_1234;
wire n_1458;
wire n_1199;
wire n_1674;
wire n_741;
wire n_1027;
wire n_1351;
wire n_625;
wire n_1189;
wire n_1212;
wire n_726;
wire n_700;
wire n_1307;
wire n_2003;
wire n_1038;
wire n_578;
wire n_1581;
wire n_1003;
wire n_1237;
wire n_1061;
wire n_1357;
wire n_1853;
wire n_783;
wire n_1738;
wire n_798;
wire n_1575;
wire n_1854;
wire n_1923;
wire n_1342;
wire n_1209;
wire n_1348;
wire n_1387;
wire n_677;
wire n_1708;
wire n_805;
wire n_1151;
wire n_1739;
wire n_2051;
wire n_1380;
wire n_1402;
wire n_1691;
wire n_1688;
wire n_1975;
wire n_1009;
wire n_1743;
wire n_1930;
wire n_1160;
wire n_883;
wire n_1238;
wire n_1991;
wire n_1724;
wire n_1032;
wire n_1247;
wire n_1547;
wire n_1553;
wire n_893;
wire n_1099;
wire n_1264;
wire n_1192;
wire n_1844;
wire n_1700;
wire n_1555;
wire n_1415;
wire n_1370;
wire n_1786;
wire n_830;
wire n_873;
wire n_1371;
wire n_1285;
wire n_1985;
wire n_1803;
wire n_1172;
wire n_852;
wire n_1590;
wire n_1532;
wire n_1393;
wire n_1517;
wire n_1867;
wire n_1704;
wire n_1078;
wire n_544;
wire n_1711;
wire n_1140;
wire n_1444;
wire n_1670;
wire n_1603;
wire n_1579;
wire n_1263;
wire n_2019;
wire n_836;
wire n_2074;
wire n_522;
wire n_1261;
wire n_945;
wire n_1649;
wire n_2018;
wire n_1903;
wire n_1511;
wire n_1143;
wire n_1422;
wire n_1232;
wire n_1772;
wire n_1572;
wire n_616;
wire n_658;
wire n_1874;
wire n_1119;
wire n_2013;
wire n_1433;
wire n_1902;
wire n_1842;
wire n_1620;
wire n_2044;
wire n_1954;
wire n_1735;
wire n_1541;
wire n_1300;
wire n_641;
wire n_822;
wire n_693;
wire n_1313;
wire n_1056;
wire n_758;
wire n_516;
wire n_1455;
wire n_1163;
wire n_1180;
wire n_943;
wire n_1798;
wire n_1550;
wire n_1591;
wire n_772;
wire n_1344;
wire n_666;
wire n_940;
wire n_770;
wire n_567;
wire n_1781;
wire n_1971;
wire n_2058;
wire n_538;
wire n_2004;
wire n_1106;
wire n_886;
wire n_1471;
wire n_953;
wire n_1094;
wire n_1345;
wire n_1820;
wire n_539;
wire n_1421;
wire n_1936;
wire n_638;
wire n_1404;
wire n_1211;
wire n_887;
wire n_1660;
wire n_1961;
wire n_1280;
wire n_713;
wire n_1400;
wire n_1467;
wire n_976;
wire n_1445;
wire n_1560;
wire n_1526;
wire n_734;
wire n_1088;
wire n_1894;
wire n_1231;
wire n_1978;
wire n_2085;
wire n_917;
wire n_574;
wire n_907;
wire n_1446;
wire n_659;
wire n_1815;
wire n_913;
wire n_1658;
wire n_808;
wire n_867;
wire n_1230;
wire n_1193;
wire n_1967;
wire n_1054;
wire n_559;
wire n_1333;
wire n_1648;
wire n_1911;
wire n_1956;
wire n_1644;
wire n_2011;
wire n_1558;
wire n_1732;
wire n_551;
wire n_699;
wire n_1986;
wire n_564;
wire n_824;
wire n_686;
wire n_757;
wire n_594;
wire n_1641;
wire n_1918;
wire n_577;
wire n_1843;
wire n_619;
wire n_1367;
wire n_1336;
wire n_521;
wire n_572;
wire n_813;
wire n_1909;
wire n_2080;
wire n_1481;
wire n_606;
wire n_1441;
wire n_818;
wire n_1123;
wire n_1309;
wire n_645;
wire n_1381;
wire n_1699;
wire n_916;
wire n_1970;
wire n_608;
wire n_630;
wire n_2059;
wire n_541;
wire n_2073;
wire n_792;
wire n_1328;
wire n_1957;
wire n_1907;
wire n_1162;
wire n_860;
wire n_1530;
wire n_788;
wire n_939;
wire n_1543;
wire n_821;
wire n_938;
wire n_1302;
wire n_1068;
wire n_1599;
wire n_982;
wire n_549;
wire n_1762;
wire n_1910;
wire n_1075;
wire n_932;
wire n_1876;
wire n_1895;
wire n_1697;
wire n_979;
wire n_1873;
wire n_905;
wire n_1866;
wire n_1680;
wire n_993;
wire n_689;
wire n_2031;
wire n_1330;
wire n_1413;
wire n_1605;
wire n_1988;
wire n_1278;
wire n_547;
wire n_558;
wire n_1064;
wire n_1396;
wire n_634;
wire n_966;
wire n_764;
wire n_1663;
wire n_2009;
wire n_692;
wire n_733;
wire n_1793;
wire n_1233;
wire n_1289;
wire n_2068;
wire n_1107;
wire n_1014;
wire n_1290;
wire n_1703;
wire n_882;
wire n_2072;
wire n_1354;
wire n_586;
wire n_1865;
wire n_1875;
wire n_1701;
wire n_1111;
wire n_1713;
wire n_715;
wire n_1251;
wire n_1265;
wire n_1726;
wire n_1950;
wire n_530;
wire n_1563;
wire n_1912;
wire n_1982;
wire n_618;
wire n_1297;
wire n_1662;
wire n_1312;
wire n_1167;
wire n_1359;
wire n_674;
wire n_871;
wire n_922;
wire n_1335;
wire n_1760;
wire n_1927;
wire n_2028;
wire n_1069;
wire n_1722;
wire n_1664;
wire n_612;
wire n_1165;
wire n_702;
wire n_2008;
wire n_1926;
wire n_1175;
wire n_1386;
wire n_1896;
wire n_1747;
wire n_1012;
wire n_780;
wire n_675;
wire n_903;
wire n_1540;
wire n_1977;
wire n_1802;
wire n_1504;
wire n_1655;
wire n_835;
wire n_928;
wire n_1214;
wire n_850;
wire n_690;
wire n_1886;
wire n_1801;
wire n_1654;
wire n_816;
wire n_1157;
wire n_1750;
wire n_1462;
wire n_1188;
wire n_1752;
wire n_877;
wire n_1813;
wire n_604;
wire n_825;
wire n_728;
wire n_1063;
wire n_1588;
wire n_1124;
wire n_1624;
wire n_1965;
wire n_598;
wire n_696;
wire n_1515;
wire n_961;
wire n_1082;
wire n_1317;
wire n_593;
wire n_697;
wire n_687;
wire n_890;
wire n_637;
wire n_701;
wire n_950;
wire n_2036;
wire n_1709;
wire n_1825;
wire n_1757;
wire n_1796;
wire n_1792;
wire n_891;
wire n_2067;
wire n_2082;
wire n_1412;
wire n_949;
wire n_1630;
wire n_678;
wire n_2075;
wire n_1987;
wire n_968;
wire n_909;
wire n_1369;
wire n_881;
wire n_1008;
wire n_760;
wire n_1546;
wire n_590;
wire n_1033;
wire n_1052;
wire n_1296;
wire n_1990;
wire n_694;
wire n_1294;
wire n_1420;
wire n_1634;
wire n_2078;
wire n_627;
wire n_595;
wire n_1767;
wire n_1779;
wire n_524;
wire n_1465;
wire n_1858;
wire n_1044;
wire n_1712;
wire n_1391;
wire n_1523;
wire n_1208;
wire n_1164;
wire n_1295;
wire n_1627;
wire n_1072;
wire n_1527;
wire n_1495;
wire n_1438;
wire n_815;
wire n_1100;
wire n_585;
wire n_1487;
wire n_840;
wire n_874;
wire n_1756;
wire n_1128;
wire n_673;
wire n_1969;
wire n_1071;
wire n_1067;
wire n_1565;
wire n_1493;
wire n_1968;
wire n_898;
wire n_1952;
wire n_865;
wire n_925;
wire n_1932;
wire n_1101;
wire n_1026;
wire n_1880;
wire n_1364;
wire n_615;
wire n_1249;
wire n_1293;
wire n_1127;
wire n_1512;
wire n_1451;
wire n_963;
wire n_639;
wire n_794;
wire n_727;
wire n_894;
wire n_1839;
wire n_685;
wire n_1765;
wire n_605;
wire n_1514;
wire n_1863;
wire n_826;
wire n_1646;
wire n_872;
wire n_1139;
wire n_1714;
wire n_718;
wire n_1018;
wire n_1521;
wire n_1366;
wire n_542;
wire n_847;
wire n_851;
wire n_682;
wire n_644;
wire n_996;
wire n_532;
wire n_1308;
wire n_1376;
wire n_1513;
wire n_791;
wire n_1913;
wire n_837;
wire n_1488;
wire n_1808;
wire n_948;
wire n_704;
wire n_977;
wire n_1005;
wire n_1947;
wire n_536;
wire n_1788;
wire n_1999;
wire n_622;
wire n_1469;
wire n_2060;
wire n_1838;
wire n_1835;
wire n_1776;
wire n_1766;
wire n_1959;
wire n_2002;
wire n_581;
wire n_765;
wire n_987;
wire n_1492;
wire n_1340;
wire n_1771;
wire n_631;
wire n_720;
wire n_842;
wire n_1707;
wire n_1432;
wire n_843;
wire n_656;
wire n_989;
wire n_1277;
wire n_797;
wire n_1473;
wire n_1723;
wire n_1246;
wire n_1878;
wire n_899;
wire n_738;
wire n_2012;
wire n_1304;
wire n_1035;
wire n_1426;
wire n_705;
wire n_1004;
wire n_1176;
wire n_1529;
wire n_1022;
wire n_614;
wire n_529;
wire n_2069;
wire n_684;
wire n_1431;
wire n_1615;
wire n_1474;
wire n_1571;
wire n_1809;
wire n_1577;
wire n_1181;
wire n_1822;
wire n_947;
wire n_1117;
wire n_1087;
wire n_1448;
wire n_1992;
wire n_648;
wire n_657;
wire n_1049;
wire n_2057;
wire n_1666;
wire n_1505;
wire n_803;
wire n_1717;
wire n_926;
wire n_1817;
wire n_927;
wire n_1849;
wire n_919;
wire n_1698;
wire n_929;
wire n_1228;
wire n_1568;
wire n_1490;
wire n_777;
wire n_1299;
wire n_526;
wire n_1183;
wire n_1436;
wire n_1384;
wire n_1070;
wire n_998;
wire n_717;
wire n_1665;
wire n_1383;
wire n_1178;
wire n_1424;
wire n_1073;
wire n_1000;
wire n_796;
wire n_1195;
wire n_1626;
wire n_1507;
wire n_552;
wire n_1358;
wire n_1811;
wire n_1388;
wire n_912;
wire n_1857;
wire n_1519;
wire n_745;
wire n_1284;
wire n_1604;
wire n_1142;
wire n_716;
wire n_1475;
wire n_623;
wire n_1048;
wire n_1201;
wire n_1398;
wire n_884;
wire n_1774;
wire n_1395;
wire n_731;
wire n_1502;
wire n_1659;
wire n_1955;
wire n_755;
wire n_931;
wire n_1021;
wire n_527;
wire n_683;
wire n_811;
wire n_1207;
wire n_1791;
wire n_1368;
wire n_1418;
wire n_958;
wire n_1250;
wire n_1137;
wire n_1897;
wire n_2064;
wire n_880;
wire n_2053;
wire n_889;
wire n_1478;
wire n_589;
wire n_1310;
wire n_819;
wire n_1363;
wire n_1334;
wire n_1966;
wire n_1942;
wire n_767;
wire n_1314;
wire n_600;
wire n_964;
wire n_831;
wire n_1837;
wire n_954;
wire n_864;
wire n_1110;
wire n_1410;
wire n_1440;
wire n_2063;
wire n_1382;
wire n_1534;
wire n_1564;
wire n_1736;
wire n_1483;
wire n_1834;
wire n_1372;
wire n_1457;
wire n_1719;
wire n_1339;
wire n_1787;
wire n_537;
wire n_1993;
wire n_1427;
wire n_1466;
wire n_1919;
wire n_1080;
wire n_723;
wire n_1877;
wire n_596;
wire n_546;
wire n_562;
wire n_1141;
wire n_1268;
wire n_1939;
wire n_2030;
wire n_1769;
wire n_1220;
wire n_1893;
wire n_556;
wire n_1755;
wire n_1602;
wire n_1136;
wire n_2025;
wire n_1125;
wire n_970;
wire n_1980;
wire n_642;
wire n_995;
wire n_1159;
wire n_1092;
wire n_1060;
wire n_1951;
wire n_1252;
wire n_1784;
wire n_1223;
wire n_1286;
wire n_1773;
wire n_1775;
wire n_1053;
wire n_1681;
wire n_520;
wire n_1093;
wire n_1783;
wire n_1533;
wire n_1597;
wire n_775;
wire n_651;
wire n_1153;
wire n_1618;
wire n_518;
wire n_1531;
wire n_1185;
wire n_1745;
wire n_914;
wire n_759;
wire n_1831;
wire n_1653;
wire n_1679;
wire n_1625;
wire n_1453;
wire n_773;
wire n_1901;
wire n_920;
wire n_1374;
wire n_1315;
wire n_1647;
wire n_1224;
wire n_1614;
wire n_1459;
wire n_1892;
wire n_1933;
wire n_1135;
wire n_1179;
wire n_1169;
wire n_1617;
wire n_1470;
wire n_1243;
wire n_848;
wire n_1096;
wire n_1091;
wire n_1917;
wire n_2000;
wire n_1580;
wire n_1425;
wire n_1881;
wire n_1281;
wire n_1267;
wire n_1806;
wire n_983;
wire n_2023;
wire n_1520;
wire n_906;
wire n_1390;
wire n_688;
wire n_1077;
wire n_1733;
wire n_1419;
wire n_1731;
wire n_1855;
wire n_1636;
wire n_1437;
wire n_1645;
wire n_1832;
wire n_1687;
wire n_1439;
wire n_1323;
wire n_858;
wire n_2049;
wire n_1331;
wire n_736;
wire n_613;
wire n_956;
wire n_960;
wire n_663;
wire n_856;
wire n_778;
wire n_1668;
wire n_1134;
wire n_1129;
wire n_554;
wire n_602;
wire n_1696;
wire n_1995;
wire n_1594;
wire n_664;
wire n_1869;
wire n_1764;
wire n_1429;
wire n_1610;
wire n_1889;
wire n_1905;
wire n_2016;
wire n_793;
wire n_587;
wire n_1593;
wire n_580;
wire n_762;
wire n_1030;
wire n_1202;
wire n_1937;
wire n_1790;
wire n_1778;
wire n_1635;
wire n_1079;
wire n_1744;
wire n_828;
wire n_607;
wire n_1551;
wire n_1103;
wire n_1203;
wire n_820;
wire n_951;
wire n_952;
wire n_725;
wire n_999;
wire n_1254;
wire n_575;
wire n_994;
wire n_1508;
wire n_732;
wire n_974;
wire n_724;
wire n_1934;
wire n_1020;
wire n_1042;
wire n_628;
wire n_1273;
wire n_1434;
wire n_1573;
wire n_1728;
wire n_557;
wire n_1871;
wire n_617;
wire n_845;
wire n_807;
wire n_1036;
wire n_1138;
wire n_1661;
wire n_1275;
wire n_1549;
wire n_1510;
wire n_892;
wire n_768;
wire n_1468;
wire n_1859;
wire n_1095;
wire n_2024;
wire n_1595;
wire n_1718;
wire n_1749;
wire n_1683;
wire n_1916;
wire n_597;
wire n_1270;
wire n_1187;
wire n_610;
wire n_1403;
wire n_1669;
wire n_1852;
wire n_1024;
wire n_1768;
wire n_1847;
wire n_2052;
wire n_517;
wire n_1667;
wire n_667;
wire n_1206;
wire n_621;
wire n_1037;
wire n_1397;
wire n_1279;
wire n_1115;
wire n_750;
wire n_901;
wire n_1499;
wire n_923;
wire n_1409;
wire n_1841;
wire n_1639;
wire n_1623;
wire n_1015;
wire n_1503;
wire n_1057;
wire n_603;
wire n_991;
wire n_1657;
wire n_1126;
wire n_1997;
wire n_710;
wire n_1108;
wire n_1818;
wire n_1182;
wire n_1298;
wire n_1611;
wire n_785;
wire n_746;
wire n_609;
wire n_1601;
wire n_1960;
wire n_2061;
wire n_1686;
wire n_1356;
wire n_1589;
wire n_1740;
wire n_1497;
wire n_1168;
wire n_1216;
wire n_1943;
wire n_1320;
wire n_1430;
wire n_1316;
wire n_1287;
wire n_1452;
wire n_1622;
wire n_1586;
wire n_1694;
wire n_1535;
wire n_1596;
wire n_1190;
wire n_1734;
wire n_1983;
wire n_1938;
wire n_1262;
wire n_1891;
wire n_1213;
wire n_1350;
wire n_1673;
wire n_1715;
wire n_1443;
wire n_1272;
wire n_2037;
wire n_782;
wire n_1539;
wire n_809;
wire n_1043;
wire n_1797;
wire n_1608;
wire n_986;
wire n_1472;
wire n_2050;
wire n_1081;
wire n_1870;
wire n_1692;
wire n_800;
wire n_1084;
wire n_1171;
wire n_1827;
wire n_1361;
wire n_1864;
wire n_2006;
wire n_1491;
wire n_662;
wire n_1152;
wire n_1840;
wire n_1705;
wire n_1684;
wire n_921;
wire n_1346;
wire n_711;
wire n_1642;
wire n_579;
wire n_1352;
wire n_937;
wire n_1682;
wire n_2017;
wire n_1695;
wire n_1828;
wire n_2046;
wire n_650;
wire n_1046;
wire n_1940;
wire n_1979;
wire n_1145;
wire n_1121;
wire n_1102;
wire n_1963;
wire n_972;
wire n_1405;
wire n_1406;
wire n_1332;
wire n_624;
wire n_962;
wire n_1041;
wire n_565;
wire n_1569;
wire n_936;
wire n_1883;
wire n_1288;
wire n_1186;
wire n_1062;
wire n_885;
wire n_896;
wire n_2084;
wire n_654;
wire n_1222;
wire n_599;
wire n_776;
wire n_1823;
wire n_1974;
wire n_1720;
wire n_934;
wire n_1637;
wire n_1407;
wire n_1795;
wire n_1341;
wire n_1456;
wire n_1845;
wire n_1489;
wire n_942;
wire n_1524;
wire n_543;
wire n_1964;
wire n_1920;
wire n_1496;
wire n_1271;
wire n_1545;
wire n_2007;
wire n_2039;
wire n_1946;
wire n_1355;
wire n_1225;
wire n_1544;
wire n_1485;
wire n_1640;
wire n_804;
wire n_1846;
wire n_533;
wire n_806;
wire n_879;
wire n_959;
wire n_584;
wire n_1343;
wire n_1522;
wire n_548;
wire n_1782;
wire n_1676;
wire n_833;
wire n_1830;
wire n_1567;
wire n_523;
wire n_1319;
wire n_707;
wire n_1900;
wire n_799;
wire n_1548;
wire n_1155;
wire n_1633;
wire n_787;
wire n_1416;
wire n_1528;
wire n_1146;
wire n_2021;
wire n_1086;
wire n_1066;
wire n_1948;
wire n_2026;
wire n_1282;
wire n_550;
wire n_652;
wire n_560;
wire n_1906;
wire n_1484;
wire n_1241;
wire n_1321;
wire n_1672;
wire n_569;
wire n_1758;
wire n_1925;
wire n_737;
wire n_1318;
wire n_1914;
wire n_1235;
wire n_1229;
wire n_1373;
wire n_1292;
wire n_1029;
wire n_1447;
wire n_2056;
wire n_790;
wire n_1706;
wire n_1498;
wire n_1210;
wire n_1248;
wire n_1556;
wire n_902;
wire n_1047;
wire n_1984;
wire n_1385;
wire n_1269;
wire n_1931;
wire n_2083;
wire n_672;
wire n_1257;
wire n_1751;
wire n_1375;
wire n_1941;
wire n_655;
wire n_706;
wire n_1045;
wire n_1650;
wire n_786;
wire n_1794;
wire n_1236;
wire n_1962;
wire n_1559;
wire n_1725;
wire n_1928;
wire n_1872;
wire n_834;
wire n_743;
wire n_766;
wire n_1741;
wire n_1325;
wire n_1002;
wire n_1746;
wire n_1949;
wire n_545;
wire n_1804;
wire n_1727;
wire n_1019;
wire n_636;
wire n_2054;
wire n_729;
wire n_876;
wire n_774;
wire n_1337;
wire n_660;
wire n_2062;
wire n_2041;
wire n_1477;
wire n_1360;
wire n_1860;
wire n_1904;
wire n_1200;
wire n_2070;
wire n_1607;
wire n_1353;
wire n_1908;
wire n_1777;
wire n_1454;
wire n_869;
wire n_1154;
wire n_1113;
wire n_1600;
wire n_646;
wire n_528;
wire n_1098;
wire n_1329;
wire n_2045;
wire n_817;
wire n_897;
wire n_846;
wire n_2066;
wire n_841;
wire n_1476;
wire n_1001;
wire n_1800;
wire n_1050;
wire n_1411;
wire n_1463;
wire n_1177;
wire n_1150;
wire n_1742;
wire n_1562;
wire n_1690;
wire n_1191;
wire n_1826;
wire n_566;
wire n_1023;
wire n_1882;
wire n_1076;
wire n_1118;
wire n_1007;
wire n_1807;
wire n_1929;
wire n_1378;
wire n_855;
wire n_1592;
wire n_1759;
wire n_1814;
wire n_1631;
wire n_591;
wire n_1377;
wire n_1879;
wire n_853;
wire n_695;
wire n_1542;
wire n_875;
wire n_680;
wire n_1678;
wire n_661;
wire n_1716;
wire n_1256;
wire n_671;
wire n_1953;
wire n_933;
wire n_740;
wire n_703;
wire n_978;
wire n_1976;
wire n_1291;
wire n_1217;
wire n_751;
wire n_749;
wire n_1824;
wire n_1628;
wire n_1324;
wire n_1399;
wire n_1435;
wire n_969;
wire n_988;
wire n_1065;
wire n_1401;
wire n_1255;
wire n_568;
wire n_1516;
wire n_1536;
wire n_2029;
wire n_1204;
wire n_823;
wire n_1132;
wire n_643;
wire n_1074;
wire n_698;
wire n_1394;
wire n_1327;
wire n_1326;
wire n_739;
wire n_955;
wire n_1379;
wire n_1338;
wire n_1097;
wire n_935;
wire n_781;
wire n_789;
wire n_1554;
wire n_1130;
wire n_1810;
wire n_573;
wire n_769;
wire n_676;
wire n_1120;
wire n_832;
wire n_1583;
wire n_1730;
wire n_555;
wire n_814;
wire n_1643;
wire n_2020;
wire n_1729;
wire n_669;
wire n_2048;
wire n_2005;
wire n_747;
wire n_1389;
wire n_1105;
wire n_721;
wire n_1461;
wire n_742;
wire n_691;
wire n_535;
wire n_2076;
wire n_1408;
wire n_1196;
wire n_1598;
wire n_863;
wire n_601;
wire n_1283;
wire n_918;
wire n_748;
wire n_1114;
wire n_1848;
wire n_1147;
wire n_763;
wire n_1785;
wire n_1754;
wire n_1506;
wire n_1652;
wire n_1812;
wire n_957;
wire n_1994;
wire n_895;
wire n_866;
wire n_1227;
wire n_744;
wire n_971;
wire n_946;
wire n_761;
wire n_1303;
wire n_1205;
wire n_1258;
wire n_1392;
wire n_1173;
wire n_1924;
wire n_525;
wire n_1677;
wire n_1116;
wire n_611;
wire n_1570;
wire n_1702;
wire n_1219;
wire n_1780;
wire n_1689;
wire n_1174;
wire n_1944;
wire n_1016;
wire n_1347;
wire n_795;
wire n_1501;
wire n_1221;
wire n_1245;
wire n_838;
wire n_647;
wire n_844;
wire n_1017;
wire n_1083;
wire n_1561;
wire n_930;
wire n_888;
wire n_1112;
wire n_2081;
wire n_2022;
wire n_1945;
wire n_910;
wire n_1721;
wire n_1656;
wire n_1460;
wire n_911;
wire n_1464;
wire n_653;
wire n_1737;
wire n_1414;
wire n_908;
wire n_752;
wire n_944;
wire n_2034;
wire n_576;
wire n_1028;
wire n_1922;
wire n_563;
wire n_2032;
wire n_1011;
wire n_1566;
wire n_1215;
wire n_839;
wire n_708;
wire n_1973;
wire n_668;
wire n_626;
wire n_990;
wire n_1500;
wire n_779;
wire n_1537;
wire n_1821;
wire n_1104;
wire n_854;
wire n_1058;
wire n_1122;
wire n_870;
wire n_904;
wire n_1253;
wire n_709;
wire n_1266;
wire n_1509;
wire n_1693;
wire n_1109;
wire n_712;
wire n_1276;
wire n_2015;
wire n_1148;
wire n_1989;
wire n_1161;
wire n_1085;
wire n_2014;
wire n_2042;
wire n_1239;
wire n_771;
wire n_1584;
wire n_924;
wire n_1582;
wire n_1149;
wire n_1184;
wire n_719;
wire n_1972;
wire n_1525;
wire n_1585;
wire n_1851;
wire n_1799;
wire n_1090;
wire n_592;
wire n_1816;
wire n_1518;
wire n_829;
wire n_1156;
wire n_1362;
wire n_984;
wire n_1829;
wire n_2035;
wire n_1450;
wire n_1638;
wire n_868;
wire n_859;
wire n_570;
wire n_2033;
wire n_735;
wire n_1789;
wire n_1770;
wire n_878;
wire n_620;
wire n_519;
wire n_1218;
wire n_1482;
wire n_981;
wire n_714;
wire n_1349;
wire n_1144;
wire n_2071;
wire n_985;
wire n_997;
wire n_1710;
wire n_1301;
wire n_802;
wire n_561;
wire n_980;
wire n_1306;
wire n_2010;
wire n_1651;
wire n_1198;
wire n_2047;
wire n_1609;
wire n_1244;
wire n_1685;
wire n_1763;
wire n_1998;
wire n_1574;
wire n_756;
wire n_1619;
wire n_1981;
wire n_1606;
wire n_810;
wire n_1133;
wire n_635;
wire n_1194;
wire n_1051;
wire n_1552;
wire n_583;
wire n_1996;
wire n_1039;
wire n_1442;
wire n_1034;
wire n_2043;
wire n_1480;
wire n_1158;
wire n_754;
wire n_941;
wire n_975;
wire n_1031;
wire n_1305;
wire n_553;
wire n_849;
wire n_753;
wire n_1753;
wire n_973;
wire n_1921;
wire n_1479;
wire n_1055;
wire n_1675;
wire n_582;
wire n_2065;
wire n_861;
wire n_857;
wire n_967;
wire n_571;
wire n_2001;
wire n_1884;
wire n_2040;
wire n_679;
wire n_633;
wire n_1170;
wire n_665;
wire n_1629;
wire n_588;
wire n_1260;
wire n_1819;
wire n_2055;
wire n_1010;
wire n_1040;
wire n_915;
wire n_632;
wire n_1166;
wire n_2038;
wire n_812;
wire n_1131;
wire n_1761;
wire n_534;
wire n_1578;
wire n_1006;
wire n_1861;
wire n_1632;
wire n_1890;
wire n_1805;
wire n_1557;
wire n_1888;
wire n_1833;
wire n_730;
wire n_1311;
wire n_1494;
wire n_670;
wire n_1850;
wire n_1898;
wire n_1868;
wire n_2079;
wire n_1089;
wire n_1887;
wire n_1587;
wire n_1365;
wire n_1417;
wire n_1242;
wire n_1836;
wire n_681;
wire n_1226;
wire n_1274;
wire n_1486;
wire n_640;
wire n_1322;
wire n_965;
wire n_1899;
wire n_1428;
wire n_1616;
wire n_1576;
wire n_1856;
wire n_1862;
wire n_1958;
wire n_2077;
wire n_784;
wire n_1059;
wire n_1197;
wire n_722;
wire n_862;
wire n_540;
wire n_1423;
wire n_1935;
wire n_2027;
wire n_1915;
wire n_629;
wire n_1621;
wire n_1748;
wire n_900;
wire n_1449;
wire n_531;
wire n_827;
wire n_1025;
wire n_1885;
wire n_1013;
wire n_1259;
wire n_1538;
wire n_649;
wire n_1612;
wire n_1240;

INVx1_ASAP7_75t_L g516 ( 
.A(n_424),
.Y(n_516)
);

INVx1_ASAP7_75t_L g517 ( 
.A(n_476),
.Y(n_517)
);

BUFx6f_ASAP7_75t_L g518 ( 
.A(n_435),
.Y(n_518)
);

CKINVDCx20_ASAP7_75t_R g519 ( 
.A(n_36),
.Y(n_519)
);

CKINVDCx5p33_ASAP7_75t_R g520 ( 
.A(n_133),
.Y(n_520)
);

INVx4_ASAP7_75t_R g521 ( 
.A(n_414),
.Y(n_521)
);

CKINVDCx5p33_ASAP7_75t_R g522 ( 
.A(n_205),
.Y(n_522)
);

CKINVDCx5p33_ASAP7_75t_R g523 ( 
.A(n_211),
.Y(n_523)
);

CKINVDCx5p33_ASAP7_75t_R g524 ( 
.A(n_362),
.Y(n_524)
);

HB1xp67_ASAP7_75t_L g525 ( 
.A(n_467),
.Y(n_525)
);

INVx1_ASAP7_75t_L g526 ( 
.A(n_100),
.Y(n_526)
);

CKINVDCx5p33_ASAP7_75t_R g527 ( 
.A(n_290),
.Y(n_527)
);

CKINVDCx5p33_ASAP7_75t_R g528 ( 
.A(n_239),
.Y(n_528)
);

INVx1_ASAP7_75t_L g529 ( 
.A(n_330),
.Y(n_529)
);

CKINVDCx5p33_ASAP7_75t_R g530 ( 
.A(n_103),
.Y(n_530)
);

INVx1_ASAP7_75t_SL g531 ( 
.A(n_341),
.Y(n_531)
);

CKINVDCx5p33_ASAP7_75t_R g532 ( 
.A(n_286),
.Y(n_532)
);

CKINVDCx5p33_ASAP7_75t_R g533 ( 
.A(n_483),
.Y(n_533)
);

CKINVDCx5p33_ASAP7_75t_R g534 ( 
.A(n_10),
.Y(n_534)
);

CKINVDCx20_ASAP7_75t_R g535 ( 
.A(n_495),
.Y(n_535)
);

CKINVDCx5p33_ASAP7_75t_R g536 ( 
.A(n_127),
.Y(n_536)
);

INVx1_ASAP7_75t_L g537 ( 
.A(n_224),
.Y(n_537)
);

CKINVDCx5p33_ASAP7_75t_R g538 ( 
.A(n_413),
.Y(n_538)
);

CKINVDCx5p33_ASAP7_75t_R g539 ( 
.A(n_428),
.Y(n_539)
);

CKINVDCx5p33_ASAP7_75t_R g540 ( 
.A(n_318),
.Y(n_540)
);

CKINVDCx20_ASAP7_75t_R g541 ( 
.A(n_58),
.Y(n_541)
);

INVx1_ASAP7_75t_L g542 ( 
.A(n_453),
.Y(n_542)
);

CKINVDCx5p33_ASAP7_75t_R g543 ( 
.A(n_117),
.Y(n_543)
);

CKINVDCx16_ASAP7_75t_R g544 ( 
.A(n_249),
.Y(n_544)
);

CKINVDCx5p33_ASAP7_75t_R g545 ( 
.A(n_317),
.Y(n_545)
);

INVx1_ASAP7_75t_L g546 ( 
.A(n_443),
.Y(n_546)
);

CKINVDCx20_ASAP7_75t_R g547 ( 
.A(n_245),
.Y(n_547)
);

INVx1_ASAP7_75t_L g548 ( 
.A(n_416),
.Y(n_548)
);

INVx1_ASAP7_75t_L g549 ( 
.A(n_32),
.Y(n_549)
);

CKINVDCx5p33_ASAP7_75t_R g550 ( 
.A(n_331),
.Y(n_550)
);

CKINVDCx5p33_ASAP7_75t_R g551 ( 
.A(n_271),
.Y(n_551)
);

CKINVDCx5p33_ASAP7_75t_R g552 ( 
.A(n_125),
.Y(n_552)
);

INVx2_ASAP7_75t_L g553 ( 
.A(n_471),
.Y(n_553)
);

CKINVDCx5p33_ASAP7_75t_R g554 ( 
.A(n_512),
.Y(n_554)
);

BUFx10_ASAP7_75t_L g555 ( 
.A(n_445),
.Y(n_555)
);

BUFx6f_ASAP7_75t_L g556 ( 
.A(n_293),
.Y(n_556)
);

CKINVDCx5p33_ASAP7_75t_R g557 ( 
.A(n_491),
.Y(n_557)
);

INVx1_ASAP7_75t_L g558 ( 
.A(n_324),
.Y(n_558)
);

CKINVDCx5p33_ASAP7_75t_R g559 ( 
.A(n_400),
.Y(n_559)
);

INVx1_ASAP7_75t_L g560 ( 
.A(n_479),
.Y(n_560)
);

CKINVDCx20_ASAP7_75t_R g561 ( 
.A(n_48),
.Y(n_561)
);

CKINVDCx5p33_ASAP7_75t_R g562 ( 
.A(n_300),
.Y(n_562)
);

CKINVDCx5p33_ASAP7_75t_R g563 ( 
.A(n_460),
.Y(n_563)
);

CKINVDCx5p33_ASAP7_75t_R g564 ( 
.A(n_266),
.Y(n_564)
);

CKINVDCx5p33_ASAP7_75t_R g565 ( 
.A(n_310),
.Y(n_565)
);

CKINVDCx5p33_ASAP7_75t_R g566 ( 
.A(n_180),
.Y(n_566)
);

CKINVDCx5p33_ASAP7_75t_R g567 ( 
.A(n_179),
.Y(n_567)
);

CKINVDCx5p33_ASAP7_75t_R g568 ( 
.A(n_315),
.Y(n_568)
);

CKINVDCx5p33_ASAP7_75t_R g569 ( 
.A(n_130),
.Y(n_569)
);

CKINVDCx5p33_ASAP7_75t_R g570 ( 
.A(n_182),
.Y(n_570)
);

CKINVDCx16_ASAP7_75t_R g571 ( 
.A(n_143),
.Y(n_571)
);

CKINVDCx5p33_ASAP7_75t_R g572 ( 
.A(n_189),
.Y(n_572)
);

CKINVDCx20_ASAP7_75t_R g573 ( 
.A(n_110),
.Y(n_573)
);

HB1xp67_ASAP7_75t_L g574 ( 
.A(n_223),
.Y(n_574)
);

INVx2_ASAP7_75t_SL g575 ( 
.A(n_153),
.Y(n_575)
);

CKINVDCx5p33_ASAP7_75t_R g576 ( 
.A(n_141),
.Y(n_576)
);

CKINVDCx5p33_ASAP7_75t_R g577 ( 
.A(n_102),
.Y(n_577)
);

INVxp67_ASAP7_75t_L g578 ( 
.A(n_66),
.Y(n_578)
);

CKINVDCx5p33_ASAP7_75t_R g579 ( 
.A(n_11),
.Y(n_579)
);

HB1xp67_ASAP7_75t_L g580 ( 
.A(n_68),
.Y(n_580)
);

BUFx6f_ASAP7_75t_L g581 ( 
.A(n_252),
.Y(n_581)
);

CKINVDCx5p33_ASAP7_75t_R g582 ( 
.A(n_180),
.Y(n_582)
);

CKINVDCx5p33_ASAP7_75t_R g583 ( 
.A(n_3),
.Y(n_583)
);

INVx1_ASAP7_75t_L g584 ( 
.A(n_287),
.Y(n_584)
);

CKINVDCx5p33_ASAP7_75t_R g585 ( 
.A(n_0),
.Y(n_585)
);

CKINVDCx5p33_ASAP7_75t_R g586 ( 
.A(n_150),
.Y(n_586)
);

CKINVDCx5p33_ASAP7_75t_R g587 ( 
.A(n_276),
.Y(n_587)
);

CKINVDCx5p33_ASAP7_75t_R g588 ( 
.A(n_299),
.Y(n_588)
);

INVx1_ASAP7_75t_L g589 ( 
.A(n_70),
.Y(n_589)
);

INVx1_ASAP7_75t_L g590 ( 
.A(n_218),
.Y(n_590)
);

INVx1_ASAP7_75t_SL g591 ( 
.A(n_370),
.Y(n_591)
);

CKINVDCx5p33_ASAP7_75t_R g592 ( 
.A(n_228),
.Y(n_592)
);

INVx2_ASAP7_75t_SL g593 ( 
.A(n_68),
.Y(n_593)
);

INVx2_ASAP7_75t_SL g594 ( 
.A(n_289),
.Y(n_594)
);

CKINVDCx5p33_ASAP7_75t_R g595 ( 
.A(n_105),
.Y(n_595)
);

CKINVDCx5p33_ASAP7_75t_R g596 ( 
.A(n_178),
.Y(n_596)
);

CKINVDCx14_ASAP7_75t_R g597 ( 
.A(n_248),
.Y(n_597)
);

CKINVDCx5p33_ASAP7_75t_R g598 ( 
.A(n_160),
.Y(n_598)
);

CKINVDCx5p33_ASAP7_75t_R g599 ( 
.A(n_294),
.Y(n_599)
);

CKINVDCx20_ASAP7_75t_R g600 ( 
.A(n_58),
.Y(n_600)
);

INVx1_ASAP7_75t_L g601 ( 
.A(n_487),
.Y(n_601)
);

INVx1_ASAP7_75t_SL g602 ( 
.A(n_254),
.Y(n_602)
);

CKINVDCx5p33_ASAP7_75t_R g603 ( 
.A(n_264),
.Y(n_603)
);

INVx1_ASAP7_75t_L g604 ( 
.A(n_160),
.Y(n_604)
);

CKINVDCx5p33_ASAP7_75t_R g605 ( 
.A(n_234),
.Y(n_605)
);

CKINVDCx5p33_ASAP7_75t_R g606 ( 
.A(n_504),
.Y(n_606)
);

INVx1_ASAP7_75t_L g607 ( 
.A(n_235),
.Y(n_607)
);

CKINVDCx16_ASAP7_75t_R g608 ( 
.A(n_72),
.Y(n_608)
);

INVx1_ASAP7_75t_L g609 ( 
.A(n_44),
.Y(n_609)
);

BUFx3_ASAP7_75t_L g610 ( 
.A(n_472),
.Y(n_610)
);

INVx2_ASAP7_75t_L g611 ( 
.A(n_153),
.Y(n_611)
);

CKINVDCx5p33_ASAP7_75t_R g612 ( 
.A(n_88),
.Y(n_612)
);

BUFx6f_ASAP7_75t_L g613 ( 
.A(n_395),
.Y(n_613)
);

INVx1_ASAP7_75t_L g614 ( 
.A(n_387),
.Y(n_614)
);

CKINVDCx5p33_ASAP7_75t_R g615 ( 
.A(n_11),
.Y(n_615)
);

CKINVDCx20_ASAP7_75t_R g616 ( 
.A(n_219),
.Y(n_616)
);

INVx1_ASAP7_75t_L g617 ( 
.A(n_3),
.Y(n_617)
);

CKINVDCx16_ASAP7_75t_R g618 ( 
.A(n_345),
.Y(n_618)
);

CKINVDCx5p33_ASAP7_75t_R g619 ( 
.A(n_88),
.Y(n_619)
);

INVx2_ASAP7_75t_L g620 ( 
.A(n_368),
.Y(n_620)
);

CKINVDCx20_ASAP7_75t_R g621 ( 
.A(n_90),
.Y(n_621)
);

INVx2_ASAP7_75t_L g622 ( 
.A(n_237),
.Y(n_622)
);

INVx1_ASAP7_75t_L g623 ( 
.A(n_232),
.Y(n_623)
);

CKINVDCx5p33_ASAP7_75t_R g624 ( 
.A(n_173),
.Y(n_624)
);

CKINVDCx5p33_ASAP7_75t_R g625 ( 
.A(n_507),
.Y(n_625)
);

CKINVDCx20_ASAP7_75t_R g626 ( 
.A(n_326),
.Y(n_626)
);

INVx1_ASAP7_75t_L g627 ( 
.A(n_217),
.Y(n_627)
);

CKINVDCx5p33_ASAP7_75t_R g628 ( 
.A(n_386),
.Y(n_628)
);

CKINVDCx5p33_ASAP7_75t_R g629 ( 
.A(n_408),
.Y(n_629)
);

CKINVDCx5p33_ASAP7_75t_R g630 ( 
.A(n_403),
.Y(n_630)
);

CKINVDCx5p33_ASAP7_75t_R g631 ( 
.A(n_477),
.Y(n_631)
);

INVx1_ASAP7_75t_L g632 ( 
.A(n_351),
.Y(n_632)
);

INVx1_ASAP7_75t_L g633 ( 
.A(n_10),
.Y(n_633)
);

INVx1_ASAP7_75t_L g634 ( 
.A(n_340),
.Y(n_634)
);

CKINVDCx5p33_ASAP7_75t_R g635 ( 
.A(n_45),
.Y(n_635)
);

CKINVDCx5p33_ASAP7_75t_R g636 ( 
.A(n_364),
.Y(n_636)
);

INVx1_ASAP7_75t_L g637 ( 
.A(n_29),
.Y(n_637)
);

CKINVDCx5p33_ASAP7_75t_R g638 ( 
.A(n_394),
.Y(n_638)
);

CKINVDCx5p33_ASAP7_75t_R g639 ( 
.A(n_151),
.Y(n_639)
);

INVxp67_ASAP7_75t_L g640 ( 
.A(n_462),
.Y(n_640)
);

INVx2_ASAP7_75t_SL g641 ( 
.A(n_496),
.Y(n_641)
);

INVx1_ASAP7_75t_L g642 ( 
.A(n_473),
.Y(n_642)
);

CKINVDCx5p33_ASAP7_75t_R g643 ( 
.A(n_84),
.Y(n_643)
);

CKINVDCx5p33_ASAP7_75t_R g644 ( 
.A(n_105),
.Y(n_644)
);

CKINVDCx5p33_ASAP7_75t_R g645 ( 
.A(n_383),
.Y(n_645)
);

INVx1_ASAP7_75t_SL g646 ( 
.A(n_399),
.Y(n_646)
);

INVx1_ASAP7_75t_L g647 ( 
.A(n_470),
.Y(n_647)
);

CKINVDCx5p33_ASAP7_75t_R g648 ( 
.A(n_481),
.Y(n_648)
);

CKINVDCx5p33_ASAP7_75t_R g649 ( 
.A(n_148),
.Y(n_649)
);

INVx2_ASAP7_75t_L g650 ( 
.A(n_474),
.Y(n_650)
);

BUFx5_ASAP7_75t_L g651 ( 
.A(n_61),
.Y(n_651)
);

INVx1_ASAP7_75t_L g652 ( 
.A(n_159),
.Y(n_652)
);

CKINVDCx5p33_ASAP7_75t_R g653 ( 
.A(n_75),
.Y(n_653)
);

INVx2_ASAP7_75t_SL g654 ( 
.A(n_63),
.Y(n_654)
);

CKINVDCx20_ASAP7_75t_R g655 ( 
.A(n_307),
.Y(n_655)
);

INVx1_ASAP7_75t_L g656 ( 
.A(n_217),
.Y(n_656)
);

INVx1_ASAP7_75t_SL g657 ( 
.A(n_103),
.Y(n_657)
);

CKINVDCx5p33_ASAP7_75t_R g658 ( 
.A(n_380),
.Y(n_658)
);

CKINVDCx5p33_ASAP7_75t_R g659 ( 
.A(n_278),
.Y(n_659)
);

CKINVDCx5p33_ASAP7_75t_R g660 ( 
.A(n_221),
.Y(n_660)
);

INVx1_ASAP7_75t_L g661 ( 
.A(n_388),
.Y(n_661)
);

CKINVDCx5p33_ASAP7_75t_R g662 ( 
.A(n_291),
.Y(n_662)
);

CKINVDCx5p33_ASAP7_75t_R g663 ( 
.A(n_339),
.Y(n_663)
);

INVx1_ASAP7_75t_L g664 ( 
.A(n_44),
.Y(n_664)
);

INVx2_ASAP7_75t_L g665 ( 
.A(n_322),
.Y(n_665)
);

INVx1_ASAP7_75t_L g666 ( 
.A(n_410),
.Y(n_666)
);

CKINVDCx5p33_ASAP7_75t_R g667 ( 
.A(n_275),
.Y(n_667)
);

INVx1_ASAP7_75t_L g668 ( 
.A(n_75),
.Y(n_668)
);

CKINVDCx5p33_ASAP7_75t_R g669 ( 
.A(n_124),
.Y(n_669)
);

INVx1_ASAP7_75t_L g670 ( 
.A(n_49),
.Y(n_670)
);

CKINVDCx5p33_ASAP7_75t_R g671 ( 
.A(n_350),
.Y(n_671)
);

CKINVDCx5p33_ASAP7_75t_R g672 ( 
.A(n_280),
.Y(n_672)
);

INVx1_ASAP7_75t_L g673 ( 
.A(n_22),
.Y(n_673)
);

CKINVDCx5p33_ASAP7_75t_R g674 ( 
.A(n_301),
.Y(n_674)
);

INVx2_ASAP7_75t_SL g675 ( 
.A(n_267),
.Y(n_675)
);

CKINVDCx5p33_ASAP7_75t_R g676 ( 
.A(n_211),
.Y(n_676)
);

BUFx2_ASAP7_75t_L g677 ( 
.A(n_506),
.Y(n_677)
);

INVx1_ASAP7_75t_L g678 ( 
.A(n_285),
.Y(n_678)
);

INVx1_ASAP7_75t_SL g679 ( 
.A(n_270),
.Y(n_679)
);

INVx1_ASAP7_75t_L g680 ( 
.A(n_478),
.Y(n_680)
);

CKINVDCx20_ASAP7_75t_R g681 ( 
.A(n_16),
.Y(n_681)
);

CKINVDCx5p33_ASAP7_75t_R g682 ( 
.A(n_283),
.Y(n_682)
);

CKINVDCx14_ASAP7_75t_R g683 ( 
.A(n_89),
.Y(n_683)
);

INVx1_ASAP7_75t_L g684 ( 
.A(n_181),
.Y(n_684)
);

INVx1_ASAP7_75t_L g685 ( 
.A(n_335),
.Y(n_685)
);

INVx1_ASAP7_75t_L g686 ( 
.A(n_415),
.Y(n_686)
);

INVx1_ASAP7_75t_L g687 ( 
.A(n_509),
.Y(n_687)
);

INVx2_ASAP7_75t_SL g688 ( 
.A(n_247),
.Y(n_688)
);

CKINVDCx5p33_ASAP7_75t_R g689 ( 
.A(n_298),
.Y(n_689)
);

CKINVDCx5p33_ASAP7_75t_R g690 ( 
.A(n_288),
.Y(n_690)
);

INVx1_ASAP7_75t_L g691 ( 
.A(n_174),
.Y(n_691)
);

CKINVDCx5p33_ASAP7_75t_R g692 ( 
.A(n_323),
.Y(n_692)
);

INVx1_ASAP7_75t_L g693 ( 
.A(n_377),
.Y(n_693)
);

INVx2_ASAP7_75t_L g694 ( 
.A(n_47),
.Y(n_694)
);

CKINVDCx5p33_ASAP7_75t_R g695 ( 
.A(n_259),
.Y(n_695)
);

CKINVDCx5p33_ASAP7_75t_R g696 ( 
.A(n_216),
.Y(n_696)
);

INVxp67_ASAP7_75t_L g697 ( 
.A(n_34),
.Y(n_697)
);

CKINVDCx5p33_ASAP7_75t_R g698 ( 
.A(n_332),
.Y(n_698)
);

CKINVDCx5p33_ASAP7_75t_R g699 ( 
.A(n_57),
.Y(n_699)
);

INVx1_ASAP7_75t_L g700 ( 
.A(n_475),
.Y(n_700)
);

INVxp67_ASAP7_75t_L g701 ( 
.A(n_442),
.Y(n_701)
);

INVx1_ASAP7_75t_L g702 ( 
.A(n_108),
.Y(n_702)
);

INVx1_ASAP7_75t_L g703 ( 
.A(n_385),
.Y(n_703)
);

CKINVDCx5p33_ASAP7_75t_R g704 ( 
.A(n_292),
.Y(n_704)
);

CKINVDCx5p33_ASAP7_75t_R g705 ( 
.A(n_210),
.Y(n_705)
);

INVx1_ASAP7_75t_L g706 ( 
.A(n_82),
.Y(n_706)
);

INVx1_ASAP7_75t_L g707 ( 
.A(n_499),
.Y(n_707)
);

CKINVDCx20_ASAP7_75t_R g708 ( 
.A(n_52),
.Y(n_708)
);

CKINVDCx5p33_ASAP7_75t_R g709 ( 
.A(n_379),
.Y(n_709)
);

INVx1_ASAP7_75t_L g710 ( 
.A(n_308),
.Y(n_710)
);

INVx1_ASAP7_75t_L g711 ( 
.A(n_24),
.Y(n_711)
);

CKINVDCx5p33_ASAP7_75t_R g712 ( 
.A(n_213),
.Y(n_712)
);

CKINVDCx5p33_ASAP7_75t_R g713 ( 
.A(n_493),
.Y(n_713)
);

CKINVDCx5p33_ASAP7_75t_R g714 ( 
.A(n_480),
.Y(n_714)
);

CKINVDCx5p33_ASAP7_75t_R g715 ( 
.A(n_197),
.Y(n_715)
);

CKINVDCx20_ASAP7_75t_R g716 ( 
.A(n_167),
.Y(n_716)
);

INVx1_ASAP7_75t_L g717 ( 
.A(n_85),
.Y(n_717)
);

INVx1_ASAP7_75t_L g718 ( 
.A(n_210),
.Y(n_718)
);

CKINVDCx5p33_ASAP7_75t_R g719 ( 
.A(n_304),
.Y(n_719)
);

CKINVDCx5p33_ASAP7_75t_R g720 ( 
.A(n_436),
.Y(n_720)
);

INVx2_ASAP7_75t_L g721 ( 
.A(n_21),
.Y(n_721)
);

CKINVDCx5p33_ASAP7_75t_R g722 ( 
.A(n_117),
.Y(n_722)
);

CKINVDCx5p33_ASAP7_75t_R g723 ( 
.A(n_455),
.Y(n_723)
);

CKINVDCx5p33_ASAP7_75t_R g724 ( 
.A(n_220),
.Y(n_724)
);

CKINVDCx5p33_ASAP7_75t_R g725 ( 
.A(n_297),
.Y(n_725)
);

INVx1_ASAP7_75t_L g726 ( 
.A(n_261),
.Y(n_726)
);

CKINVDCx5p33_ASAP7_75t_R g727 ( 
.A(n_524),
.Y(n_727)
);

INVx1_ASAP7_75t_L g728 ( 
.A(n_651),
.Y(n_728)
);

BUFx6f_ASAP7_75t_L g729 ( 
.A(n_518),
.Y(n_729)
);

INVx1_ASAP7_75t_L g730 ( 
.A(n_651),
.Y(n_730)
);

INVx1_ASAP7_75t_L g731 ( 
.A(n_651),
.Y(n_731)
);

INVx1_ASAP7_75t_L g732 ( 
.A(n_651),
.Y(n_732)
);

CKINVDCx20_ASAP7_75t_R g733 ( 
.A(n_519),
.Y(n_733)
);

INVx1_ASAP7_75t_L g734 ( 
.A(n_651),
.Y(n_734)
);

INVxp67_ASAP7_75t_L g735 ( 
.A(n_580),
.Y(n_735)
);

INVx1_ASAP7_75t_L g736 ( 
.A(n_651),
.Y(n_736)
);

INVx1_ASAP7_75t_L g737 ( 
.A(n_651),
.Y(n_737)
);

CKINVDCx20_ASAP7_75t_R g738 ( 
.A(n_519),
.Y(n_738)
);

INVx1_ASAP7_75t_L g739 ( 
.A(n_526),
.Y(n_739)
);

CKINVDCx20_ASAP7_75t_R g740 ( 
.A(n_561),
.Y(n_740)
);

INVx1_ASAP7_75t_L g741 ( 
.A(n_549),
.Y(n_741)
);

INVx1_ASAP7_75t_L g742 ( 
.A(n_589),
.Y(n_742)
);

CKINVDCx20_ASAP7_75t_R g743 ( 
.A(n_561),
.Y(n_743)
);

INVxp67_ASAP7_75t_SL g744 ( 
.A(n_525),
.Y(n_744)
);

INVx1_ASAP7_75t_L g745 ( 
.A(n_590),
.Y(n_745)
);

INVx2_ASAP7_75t_L g746 ( 
.A(n_611),
.Y(n_746)
);

INVx1_ASAP7_75t_L g747 ( 
.A(n_604),
.Y(n_747)
);

INVx1_ASAP7_75t_L g748 ( 
.A(n_609),
.Y(n_748)
);

CKINVDCx20_ASAP7_75t_R g749 ( 
.A(n_573),
.Y(n_749)
);

INVx1_ASAP7_75t_L g750 ( 
.A(n_617),
.Y(n_750)
);

INVx1_ASAP7_75t_L g751 ( 
.A(n_627),
.Y(n_751)
);

CKINVDCx20_ASAP7_75t_R g752 ( 
.A(n_573),
.Y(n_752)
);

INVx1_ASAP7_75t_L g753 ( 
.A(n_633),
.Y(n_753)
);

INVx1_ASAP7_75t_L g754 ( 
.A(n_637),
.Y(n_754)
);

INVxp67_ASAP7_75t_SL g755 ( 
.A(n_574),
.Y(n_755)
);

INVx1_ASAP7_75t_L g756 ( 
.A(n_652),
.Y(n_756)
);

CKINVDCx5p33_ASAP7_75t_R g757 ( 
.A(n_527),
.Y(n_757)
);

CKINVDCx20_ASAP7_75t_R g758 ( 
.A(n_600),
.Y(n_758)
);

CKINVDCx20_ASAP7_75t_R g759 ( 
.A(n_600),
.Y(n_759)
);

INVx1_ASAP7_75t_L g760 ( 
.A(n_656),
.Y(n_760)
);

BUFx10_ASAP7_75t_L g761 ( 
.A(n_520),
.Y(n_761)
);

CKINVDCx5p33_ASAP7_75t_R g762 ( 
.A(n_528),
.Y(n_762)
);

HB1xp67_ASAP7_75t_L g763 ( 
.A(n_571),
.Y(n_763)
);

INVx2_ASAP7_75t_L g764 ( 
.A(n_611),
.Y(n_764)
);

INVx1_ASAP7_75t_L g765 ( 
.A(n_664),
.Y(n_765)
);

INVx3_ASAP7_75t_L g766 ( 
.A(n_694),
.Y(n_766)
);

CKINVDCx5p33_ASAP7_75t_R g767 ( 
.A(n_532),
.Y(n_767)
);

CKINVDCx5p33_ASAP7_75t_R g768 ( 
.A(n_533),
.Y(n_768)
);

INVx1_ASAP7_75t_L g769 ( 
.A(n_668),
.Y(n_769)
);

INVx1_ASAP7_75t_L g770 ( 
.A(n_670),
.Y(n_770)
);

INVx1_ASAP7_75t_L g771 ( 
.A(n_673),
.Y(n_771)
);

CKINVDCx5p33_ASAP7_75t_R g772 ( 
.A(n_538),
.Y(n_772)
);

CKINVDCx5p33_ASAP7_75t_R g773 ( 
.A(n_539),
.Y(n_773)
);

INVxp67_ASAP7_75t_SL g774 ( 
.A(n_677),
.Y(n_774)
);

INVx1_ASAP7_75t_L g775 ( 
.A(n_684),
.Y(n_775)
);

INVx1_ASAP7_75t_L g776 ( 
.A(n_691),
.Y(n_776)
);

INVxp33_ASAP7_75t_L g777 ( 
.A(n_694),
.Y(n_777)
);

INVx1_ASAP7_75t_L g778 ( 
.A(n_702),
.Y(n_778)
);

INVx1_ASAP7_75t_L g779 ( 
.A(n_706),
.Y(n_779)
);

INVx1_ASAP7_75t_L g780 ( 
.A(n_711),
.Y(n_780)
);

INVxp67_ASAP7_75t_L g781 ( 
.A(n_717),
.Y(n_781)
);

INVx2_ASAP7_75t_L g782 ( 
.A(n_721),
.Y(n_782)
);

INVxp33_ASAP7_75t_L g783 ( 
.A(n_721),
.Y(n_783)
);

INVx2_ASAP7_75t_L g784 ( 
.A(n_718),
.Y(n_784)
);

INVx1_ASAP7_75t_L g785 ( 
.A(n_610),
.Y(n_785)
);

INVx1_ASAP7_75t_L g786 ( 
.A(n_610),
.Y(n_786)
);

CKINVDCx5p33_ASAP7_75t_R g787 ( 
.A(n_540),
.Y(n_787)
);

CKINVDCx5p33_ASAP7_75t_R g788 ( 
.A(n_545),
.Y(n_788)
);

INVx1_ASAP7_75t_L g789 ( 
.A(n_516),
.Y(n_789)
);

INVx2_ASAP7_75t_L g790 ( 
.A(n_518),
.Y(n_790)
);

CKINVDCx20_ASAP7_75t_R g791 ( 
.A(n_616),
.Y(n_791)
);

INVx1_ASAP7_75t_L g792 ( 
.A(n_517),
.Y(n_792)
);

INVx1_ASAP7_75t_L g793 ( 
.A(n_529),
.Y(n_793)
);

BUFx3_ASAP7_75t_L g794 ( 
.A(n_555),
.Y(n_794)
);

INVxp33_ASAP7_75t_L g795 ( 
.A(n_553),
.Y(n_795)
);

INVxp67_ASAP7_75t_SL g796 ( 
.A(n_640),
.Y(n_796)
);

INVx1_ASAP7_75t_L g797 ( 
.A(n_537),
.Y(n_797)
);

INVx1_ASAP7_75t_L g798 ( 
.A(n_542),
.Y(n_798)
);

INVx1_ASAP7_75t_L g799 ( 
.A(n_546),
.Y(n_799)
);

INVx1_ASAP7_75t_L g800 ( 
.A(n_548),
.Y(n_800)
);

CKINVDCx5p33_ASAP7_75t_R g801 ( 
.A(n_550),
.Y(n_801)
);

INVx1_ASAP7_75t_L g802 ( 
.A(n_558),
.Y(n_802)
);

INVx1_ASAP7_75t_L g803 ( 
.A(n_560),
.Y(n_803)
);

INVx1_ASAP7_75t_L g804 ( 
.A(n_584),
.Y(n_804)
);

INVx1_ASAP7_75t_L g805 ( 
.A(n_601),
.Y(n_805)
);

INVx1_ASAP7_75t_L g806 ( 
.A(n_607),
.Y(n_806)
);

BUFx2_ASAP7_75t_L g807 ( 
.A(n_683),
.Y(n_807)
);

INVx1_ASAP7_75t_L g808 ( 
.A(n_614),
.Y(n_808)
);

INVx1_ASAP7_75t_L g809 ( 
.A(n_623),
.Y(n_809)
);

CKINVDCx16_ASAP7_75t_R g810 ( 
.A(n_608),
.Y(n_810)
);

CKINVDCx5p33_ASAP7_75t_R g811 ( 
.A(n_551),
.Y(n_811)
);

CKINVDCx5p33_ASAP7_75t_R g812 ( 
.A(n_554),
.Y(n_812)
);

CKINVDCx20_ASAP7_75t_R g813 ( 
.A(n_616),
.Y(n_813)
);

CKINVDCx5p33_ASAP7_75t_R g814 ( 
.A(n_557),
.Y(n_814)
);

INVx1_ASAP7_75t_L g815 ( 
.A(n_632),
.Y(n_815)
);

INVx1_ASAP7_75t_L g816 ( 
.A(n_634),
.Y(n_816)
);

INVx1_ASAP7_75t_L g817 ( 
.A(n_642),
.Y(n_817)
);

INVx1_ASAP7_75t_L g818 ( 
.A(n_647),
.Y(n_818)
);

CKINVDCx16_ASAP7_75t_R g819 ( 
.A(n_544),
.Y(n_819)
);

INVx1_ASAP7_75t_L g820 ( 
.A(n_790),
.Y(n_820)
);

INVx2_ASAP7_75t_L g821 ( 
.A(n_790),
.Y(n_821)
);

BUFx6f_ASAP7_75t_L g822 ( 
.A(n_729),
.Y(n_822)
);

CKINVDCx6p67_ASAP7_75t_R g823 ( 
.A(n_810),
.Y(n_823)
);

NAND2xp5_ASAP7_75t_SL g824 ( 
.A(n_819),
.B(n_807),
.Y(n_824)
);

NAND2xp5_ASAP7_75t_SL g825 ( 
.A(n_794),
.B(n_618),
.Y(n_825)
);

INVx1_ASAP7_75t_L g826 ( 
.A(n_746),
.Y(n_826)
);

INVx1_ASAP7_75t_L g827 ( 
.A(n_746),
.Y(n_827)
);

HB1xp67_ASAP7_75t_L g828 ( 
.A(n_763),
.Y(n_828)
);

INVx1_ASAP7_75t_L g829 ( 
.A(n_764),
.Y(n_829)
);

INVx2_ASAP7_75t_L g830 ( 
.A(n_729),
.Y(n_830)
);

NAND2x1_ASAP7_75t_L g831 ( 
.A(n_729),
.B(n_521),
.Y(n_831)
);

INVx1_ASAP7_75t_L g832 ( 
.A(n_764),
.Y(n_832)
);

BUFx6f_ASAP7_75t_L g833 ( 
.A(n_729),
.Y(n_833)
);

HB1xp67_ASAP7_75t_L g834 ( 
.A(n_794),
.Y(n_834)
);

CKINVDCx20_ASAP7_75t_R g835 ( 
.A(n_733),
.Y(n_835)
);

OAI22xp5_ASAP7_75t_L g836 ( 
.A1(n_774),
.A2(n_683),
.B1(n_755),
.B2(n_744),
.Y(n_836)
);

INVx1_ASAP7_75t_L g837 ( 
.A(n_782),
.Y(n_837)
);

INVx2_ASAP7_75t_L g838 ( 
.A(n_728),
.Y(n_838)
);

BUFx6f_ASAP7_75t_L g839 ( 
.A(n_782),
.Y(n_839)
);

INVx1_ASAP7_75t_L g840 ( 
.A(n_784),
.Y(n_840)
);

BUFx6f_ASAP7_75t_L g841 ( 
.A(n_730),
.Y(n_841)
);

AND2x2_ASAP7_75t_L g842 ( 
.A(n_795),
.B(n_597),
.Y(n_842)
);

INVx1_ASAP7_75t_L g843 ( 
.A(n_784),
.Y(n_843)
);

INVx2_ASAP7_75t_L g844 ( 
.A(n_731),
.Y(n_844)
);

INVx1_ASAP7_75t_L g845 ( 
.A(n_732),
.Y(n_845)
);

NOR2xp33_ASAP7_75t_SL g846 ( 
.A(n_761),
.B(n_655),
.Y(n_846)
);

BUFx2_ASAP7_75t_L g847 ( 
.A(n_727),
.Y(n_847)
);

INVx2_ASAP7_75t_L g848 ( 
.A(n_734),
.Y(n_848)
);

AND2x2_ASAP7_75t_L g849 ( 
.A(n_795),
.B(n_597),
.Y(n_849)
);

AND2x4_ASAP7_75t_L g850 ( 
.A(n_789),
.B(n_594),
.Y(n_850)
);

INVx3_ASAP7_75t_L g851 ( 
.A(n_736),
.Y(n_851)
);

INVx2_ASAP7_75t_L g852 ( 
.A(n_737),
.Y(n_852)
);

AND3x1_ASAP7_75t_L g853 ( 
.A(n_785),
.B(n_593),
.C(n_575),
.Y(n_853)
);

INVx3_ASAP7_75t_L g854 ( 
.A(n_766),
.Y(n_854)
);

INVx1_ASAP7_75t_L g855 ( 
.A(n_739),
.Y(n_855)
);

INVx1_ASAP7_75t_L g856 ( 
.A(n_741),
.Y(n_856)
);

NOR2xp33_ASAP7_75t_L g857 ( 
.A(n_757),
.B(n_531),
.Y(n_857)
);

INVx2_ASAP7_75t_L g858 ( 
.A(n_792),
.Y(n_858)
);

INVx2_ASAP7_75t_L g859 ( 
.A(n_793),
.Y(n_859)
);

AND2x2_ASAP7_75t_L g860 ( 
.A(n_786),
.B(n_654),
.Y(n_860)
);

INVx1_ASAP7_75t_L g861 ( 
.A(n_742),
.Y(n_861)
);

BUFx6f_ASAP7_75t_L g862 ( 
.A(n_797),
.Y(n_862)
);

INVx1_ASAP7_75t_L g863 ( 
.A(n_745),
.Y(n_863)
);

INVx2_ASAP7_75t_L g864 ( 
.A(n_798),
.Y(n_864)
);

OAI22xp5_ASAP7_75t_SL g865 ( 
.A1(n_733),
.A2(n_621),
.B1(n_681),
.B2(n_541),
.Y(n_865)
);

INVx4_ASAP7_75t_L g866 ( 
.A(n_766),
.Y(n_866)
);

INVx2_ASAP7_75t_L g867 ( 
.A(n_799),
.Y(n_867)
);

BUFx3_ASAP7_75t_L g868 ( 
.A(n_800),
.Y(n_868)
);

INVx1_ASAP7_75t_L g869 ( 
.A(n_747),
.Y(n_869)
);

INVx2_ASAP7_75t_L g870 ( 
.A(n_802),
.Y(n_870)
);

NAND2xp5_ASAP7_75t_L g871 ( 
.A(n_762),
.B(n_641),
.Y(n_871)
);

AND2x4_ASAP7_75t_L g872 ( 
.A(n_803),
.B(n_675),
.Y(n_872)
);

BUFx3_ASAP7_75t_L g873 ( 
.A(n_804),
.Y(n_873)
);

BUFx6f_ASAP7_75t_L g874 ( 
.A(n_805),
.Y(n_874)
);

INVx2_ASAP7_75t_L g875 ( 
.A(n_806),
.Y(n_875)
);

AND2x2_ASAP7_75t_L g876 ( 
.A(n_777),
.B(n_555),
.Y(n_876)
);

INVx2_ASAP7_75t_L g877 ( 
.A(n_808),
.Y(n_877)
);

CKINVDCx11_ASAP7_75t_R g878 ( 
.A(n_738),
.Y(n_878)
);

CKINVDCx20_ASAP7_75t_R g879 ( 
.A(n_738),
.Y(n_879)
);

INVx1_ASAP7_75t_L g880 ( 
.A(n_845),
.Y(n_880)
);

INVx1_ASAP7_75t_L g881 ( 
.A(n_845),
.Y(n_881)
);

INVx1_ASAP7_75t_L g882 ( 
.A(n_838),
.Y(n_882)
);

BUFx2_ASAP7_75t_L g883 ( 
.A(n_876),
.Y(n_883)
);

AND2x2_ASAP7_75t_L g884 ( 
.A(n_876),
.B(n_860),
.Y(n_884)
);

INVx1_ASAP7_75t_L g885 ( 
.A(n_838),
.Y(n_885)
);

INVx3_ASAP7_75t_L g886 ( 
.A(n_822),
.Y(n_886)
);

INVx1_ASAP7_75t_L g887 ( 
.A(n_848),
.Y(n_887)
);

INVx1_ASAP7_75t_L g888 ( 
.A(n_848),
.Y(n_888)
);

INVx1_ASAP7_75t_L g889 ( 
.A(n_852),
.Y(n_889)
);

HB1xp67_ASAP7_75t_L g890 ( 
.A(n_828),
.Y(n_890)
);

AOI22xp5_ASAP7_75t_SL g891 ( 
.A1(n_836),
.A2(n_681),
.B1(n_621),
.B2(n_708),
.Y(n_891)
);

INVx1_ASAP7_75t_L g892 ( 
.A(n_852),
.Y(n_892)
);

INVx2_ASAP7_75t_L g893 ( 
.A(n_821),
.Y(n_893)
);

HB1xp67_ASAP7_75t_L g894 ( 
.A(n_834),
.Y(n_894)
);

INVx1_ASAP7_75t_SL g895 ( 
.A(n_878),
.Y(n_895)
);

INVx2_ASAP7_75t_L g896 ( 
.A(n_821),
.Y(n_896)
);

NAND2xp33_ASAP7_75t_R g897 ( 
.A(n_847),
.B(n_767),
.Y(n_897)
);

BUFx6f_ASAP7_75t_L g898 ( 
.A(n_822),
.Y(n_898)
);

INVx1_ASAP7_75t_L g899 ( 
.A(n_844),
.Y(n_899)
);

NAND2xp5_ASAP7_75t_L g900 ( 
.A(n_842),
.B(n_768),
.Y(n_900)
);

NAND2xp5_ASAP7_75t_SL g901 ( 
.A(n_842),
.B(n_553),
.Y(n_901)
);

INVx1_ASAP7_75t_L g902 ( 
.A(n_844),
.Y(n_902)
);

INVx1_ASAP7_75t_L g903 ( 
.A(n_844),
.Y(n_903)
);

INVx3_ASAP7_75t_L g904 ( 
.A(n_822),
.Y(n_904)
);

HB1xp67_ASAP7_75t_L g905 ( 
.A(n_868),
.Y(n_905)
);

INVx1_ASAP7_75t_L g906 ( 
.A(n_841),
.Y(n_906)
);

INVx3_ASAP7_75t_L g907 ( 
.A(n_822),
.Y(n_907)
);

INVx2_ASAP7_75t_L g908 ( 
.A(n_839),
.Y(n_908)
);

NAND2xp5_ASAP7_75t_L g909 ( 
.A(n_849),
.B(n_772),
.Y(n_909)
);

BUFx6f_ASAP7_75t_L g910 ( 
.A(n_822),
.Y(n_910)
);

INVx2_ASAP7_75t_L g911 ( 
.A(n_839),
.Y(n_911)
);

INVx1_ASAP7_75t_L g912 ( 
.A(n_841),
.Y(n_912)
);

INVx2_ASAP7_75t_L g913 ( 
.A(n_839),
.Y(n_913)
);

CKINVDCx20_ASAP7_75t_R g914 ( 
.A(n_835),
.Y(n_914)
);

INVx1_ASAP7_75t_L g915 ( 
.A(n_841),
.Y(n_915)
);

INVx2_ASAP7_75t_L g916 ( 
.A(n_839),
.Y(n_916)
);

INVx2_ASAP7_75t_L g917 ( 
.A(n_839),
.Y(n_917)
);

AND2x4_ASAP7_75t_L g918 ( 
.A(n_868),
.B(n_748),
.Y(n_918)
);

HB1xp67_ASAP7_75t_L g919 ( 
.A(n_868),
.Y(n_919)
);

BUFx6f_ASAP7_75t_L g920 ( 
.A(n_833),
.Y(n_920)
);

NAND2xp5_ASAP7_75t_L g921 ( 
.A(n_849),
.B(n_773),
.Y(n_921)
);

INVx2_ASAP7_75t_L g922 ( 
.A(n_820),
.Y(n_922)
);

AND2x4_ASAP7_75t_L g923 ( 
.A(n_873),
.B(n_750),
.Y(n_923)
);

INVx3_ASAP7_75t_L g924 ( 
.A(n_833),
.Y(n_924)
);

BUFx6f_ASAP7_75t_L g925 ( 
.A(n_833),
.Y(n_925)
);

NAND2xp5_ASAP7_75t_L g926 ( 
.A(n_857),
.B(n_787),
.Y(n_926)
);

INVx1_ASAP7_75t_L g927 ( 
.A(n_841),
.Y(n_927)
);

INVx1_ASAP7_75t_L g928 ( 
.A(n_851),
.Y(n_928)
);

INVx2_ASAP7_75t_L g929 ( 
.A(n_820),
.Y(n_929)
);

BUFx2_ASAP7_75t_L g930 ( 
.A(n_853),
.Y(n_930)
);

INVx3_ASAP7_75t_L g931 ( 
.A(n_833),
.Y(n_931)
);

INVx1_ASAP7_75t_L g932 ( 
.A(n_851),
.Y(n_932)
);

HB1xp67_ASAP7_75t_L g933 ( 
.A(n_873),
.Y(n_933)
);

NAND2xp5_ASAP7_75t_L g934 ( 
.A(n_866),
.B(n_788),
.Y(n_934)
);

NAND2xp5_ASAP7_75t_SL g935 ( 
.A(n_871),
.B(n_620),
.Y(n_935)
);

BUFx6f_ASAP7_75t_L g936 ( 
.A(n_833),
.Y(n_936)
);

INVx1_ASAP7_75t_L g937 ( 
.A(n_851),
.Y(n_937)
);

OAI22xp33_ASAP7_75t_SL g938 ( 
.A1(n_825),
.A2(n_735),
.B1(n_796),
.B2(n_781),
.Y(n_938)
);

INVx1_ASAP7_75t_L g939 ( 
.A(n_851),
.Y(n_939)
);

INVx1_ASAP7_75t_L g940 ( 
.A(n_855),
.Y(n_940)
);

INVx1_ASAP7_75t_SL g941 ( 
.A(n_879),
.Y(n_941)
);

INVxp67_ASAP7_75t_L g942 ( 
.A(n_846),
.Y(n_942)
);

NAND2xp5_ASAP7_75t_SL g943 ( 
.A(n_850),
.B(n_620),
.Y(n_943)
);

INVx1_ASAP7_75t_L g944 ( 
.A(n_855),
.Y(n_944)
);

INVx1_ASAP7_75t_L g945 ( 
.A(n_856),
.Y(n_945)
);

INVx2_ASAP7_75t_L g946 ( 
.A(n_830),
.Y(n_946)
);

INVx1_ASAP7_75t_L g947 ( 
.A(n_856),
.Y(n_947)
);

INVx2_ASAP7_75t_L g948 ( 
.A(n_858),
.Y(n_948)
);

NAND2xp5_ASAP7_75t_L g949 ( 
.A(n_866),
.B(n_801),
.Y(n_949)
);

INVx1_ASAP7_75t_L g950 ( 
.A(n_861),
.Y(n_950)
);

NAND2xp5_ASAP7_75t_SL g951 ( 
.A(n_850),
.B(n_622),
.Y(n_951)
);

HB1xp67_ASAP7_75t_L g952 ( 
.A(n_873),
.Y(n_952)
);

BUFx2_ASAP7_75t_L g953 ( 
.A(n_853),
.Y(n_953)
);

INVx2_ASAP7_75t_L g954 ( 
.A(n_858),
.Y(n_954)
);

INVx1_ASAP7_75t_L g955 ( 
.A(n_861),
.Y(n_955)
);

INVx1_ASAP7_75t_L g956 ( 
.A(n_863),
.Y(n_956)
);

OAI22xp5_ASAP7_75t_SL g957 ( 
.A1(n_865),
.A2(n_716),
.B1(n_743),
.B2(n_740),
.Y(n_957)
);

INVx1_ASAP7_75t_L g958 ( 
.A(n_858),
.Y(n_958)
);

INVx1_ASAP7_75t_L g959 ( 
.A(n_863),
.Y(n_959)
);

NAND2xp5_ASAP7_75t_SL g960 ( 
.A(n_883),
.B(n_847),
.Y(n_960)
);

NAND2xp5_ASAP7_75t_L g961 ( 
.A(n_884),
.B(n_811),
.Y(n_961)
);

INVx1_ASAP7_75t_L g962 ( 
.A(n_940),
.Y(n_962)
);

INVx2_ASAP7_75t_L g963 ( 
.A(n_893),
.Y(n_963)
);

NOR2xp33_ASAP7_75t_L g964 ( 
.A(n_926),
.B(n_812),
.Y(n_964)
);

AND2x2_ASAP7_75t_L g965 ( 
.A(n_884),
.B(n_777),
.Y(n_965)
);

INVx1_ASAP7_75t_L g966 ( 
.A(n_944),
.Y(n_966)
);

A2O1A1Ixp33_ASAP7_75t_L g967 ( 
.A1(n_880),
.A2(n_872),
.B(n_850),
.C(n_622),
.Y(n_967)
);

INVx1_ASAP7_75t_L g968 ( 
.A(n_945),
.Y(n_968)
);

INVx1_ASAP7_75t_L g969 ( 
.A(n_947),
.Y(n_969)
);

INVx2_ASAP7_75t_L g970 ( 
.A(n_893),
.Y(n_970)
);

AOI22xp5_ASAP7_75t_L g971 ( 
.A1(n_883),
.A2(n_655),
.B1(n_850),
.B2(n_872),
.Y(n_971)
);

INVx2_ASAP7_75t_L g972 ( 
.A(n_896),
.Y(n_972)
);

NAND2xp5_ASAP7_75t_L g973 ( 
.A(n_881),
.B(n_814),
.Y(n_973)
);

NAND2xp5_ASAP7_75t_L g974 ( 
.A(n_934),
.B(n_866),
.Y(n_974)
);

NAND2xp33_ASAP7_75t_L g975 ( 
.A(n_949),
.B(n_900),
.Y(n_975)
);

NOR2xp67_ASAP7_75t_L g976 ( 
.A(n_889),
.B(n_866),
.Y(n_976)
);

INVx2_ASAP7_75t_L g977 ( 
.A(n_896),
.Y(n_977)
);

NAND2xp5_ASAP7_75t_L g978 ( 
.A(n_950),
.B(n_831),
.Y(n_978)
);

AO21x2_ASAP7_75t_L g979 ( 
.A1(n_901),
.A2(n_666),
.B(n_661),
.Y(n_979)
);

NAND2xp5_ASAP7_75t_L g980 ( 
.A(n_955),
.B(n_831),
.Y(n_980)
);

NAND2xp5_ASAP7_75t_L g981 ( 
.A(n_956),
.B(n_862),
.Y(n_981)
);

NOR2xp33_ASAP7_75t_L g982 ( 
.A(n_909),
.B(n_824),
.Y(n_982)
);

INVx1_ASAP7_75t_L g983 ( 
.A(n_959),
.Y(n_983)
);

NAND2xp5_ASAP7_75t_L g984 ( 
.A(n_921),
.B(n_862),
.Y(n_984)
);

BUFx3_ASAP7_75t_L g985 ( 
.A(n_914),
.Y(n_985)
);

BUFx5_ASAP7_75t_L g986 ( 
.A(n_928),
.Y(n_986)
);

NAND3xp33_ASAP7_75t_L g987 ( 
.A(n_935),
.B(n_860),
.C(n_872),
.Y(n_987)
);

OR2x6_ASAP7_75t_L g988 ( 
.A(n_890),
.B(n_865),
.Y(n_988)
);

NOR2xp33_ASAP7_75t_L g989 ( 
.A(n_905),
.B(n_761),
.Y(n_989)
);

NAND2xp5_ASAP7_75t_L g990 ( 
.A(n_901),
.B(n_862),
.Y(n_990)
);

INVx1_ASAP7_75t_L g991 ( 
.A(n_919),
.Y(n_991)
);

INVxp33_ASAP7_75t_L g992 ( 
.A(n_957),
.Y(n_992)
);

NOR2xp67_ASAP7_75t_L g993 ( 
.A(n_889),
.B(n_859),
.Y(n_993)
);

INVx1_ASAP7_75t_L g994 ( 
.A(n_933),
.Y(n_994)
);

NAND2xp5_ASAP7_75t_L g995 ( 
.A(n_935),
.B(n_862),
.Y(n_995)
);

NOR2xp33_ASAP7_75t_L g996 ( 
.A(n_952),
.B(n_823),
.Y(n_996)
);

OA21x2_ASAP7_75t_L g997 ( 
.A1(n_932),
.A2(n_815),
.B(n_809),
.Y(n_997)
);

INVx1_ASAP7_75t_L g998 ( 
.A(n_918),
.Y(n_998)
);

AND2x2_ASAP7_75t_SL g999 ( 
.A(n_930),
.B(n_650),
.Y(n_999)
);

INVxp67_ASAP7_75t_L g1000 ( 
.A(n_894),
.Y(n_1000)
);

NAND2xp5_ASAP7_75t_SL g1001 ( 
.A(n_938),
.B(n_872),
.Y(n_1001)
);

INVx2_ASAP7_75t_L g1002 ( 
.A(n_948),
.Y(n_1002)
);

INVxp67_ASAP7_75t_L g1003 ( 
.A(n_897),
.Y(n_1003)
);

INVx1_ASAP7_75t_SL g1004 ( 
.A(n_914),
.Y(n_1004)
);

NOR2xp67_ASAP7_75t_L g1005 ( 
.A(n_882),
.B(n_864),
.Y(n_1005)
);

AOI22xp5_ASAP7_75t_L g1006 ( 
.A1(n_930),
.A2(n_547),
.B1(n_626),
.B2(n_535),
.Y(n_1006)
);

BUFx6f_ASAP7_75t_L g1007 ( 
.A(n_918),
.Y(n_1007)
);

NAND2xp5_ASAP7_75t_SL g1008 ( 
.A(n_918),
.B(n_591),
.Y(n_1008)
);

BUFx6f_ASAP7_75t_L g1009 ( 
.A(n_923),
.Y(n_1009)
);

NAND2xp5_ASAP7_75t_SL g1010 ( 
.A(n_923),
.B(n_602),
.Y(n_1010)
);

INVx1_ASAP7_75t_L g1011 ( 
.A(n_948),
.Y(n_1011)
);

INVx2_ASAP7_75t_SL g1012 ( 
.A(n_943),
.Y(n_1012)
);

NAND2xp5_ASAP7_75t_L g1013 ( 
.A(n_937),
.B(n_874),
.Y(n_1013)
);

NAND3xp33_ASAP7_75t_L g1014 ( 
.A(n_943),
.B(n_817),
.C(n_816),
.Y(n_1014)
);

NAND2xp5_ASAP7_75t_L g1015 ( 
.A(n_939),
.B(n_862),
.Y(n_1015)
);

NAND2xp5_ASAP7_75t_SL g1016 ( 
.A(n_942),
.B(n_646),
.Y(n_1016)
);

NAND2xp5_ASAP7_75t_L g1017 ( 
.A(n_885),
.B(n_874),
.Y(n_1017)
);

INVx1_ASAP7_75t_L g1018 ( 
.A(n_954),
.Y(n_1018)
);

NAND2xp5_ASAP7_75t_L g1019 ( 
.A(n_887),
.B(n_874),
.Y(n_1019)
);

AOI22xp33_ASAP7_75t_L g1020 ( 
.A1(n_888),
.A2(n_665),
.B1(n_650),
.B2(n_678),
.Y(n_1020)
);

INVxp67_ASAP7_75t_SL g1021 ( 
.A(n_898),
.Y(n_1021)
);

AND2x2_ASAP7_75t_L g1022 ( 
.A(n_953),
.B(n_783),
.Y(n_1022)
);

INVx2_ASAP7_75t_L g1023 ( 
.A(n_922),
.Y(n_1023)
);

NOR2xp33_ASAP7_75t_L g1024 ( 
.A(n_941),
.B(n_891),
.Y(n_1024)
);

NAND2xp5_ASAP7_75t_L g1025 ( 
.A(n_892),
.B(n_874),
.Y(n_1025)
);

NOR3xp33_ASAP7_75t_L g1026 ( 
.A(n_895),
.B(n_697),
.C(n_578),
.Y(n_1026)
);

INVx1_ASAP7_75t_L g1027 ( 
.A(n_922),
.Y(n_1027)
);

NAND2xp5_ASAP7_75t_SL g1028 ( 
.A(n_958),
.B(n_679),
.Y(n_1028)
);

NAND2xp33_ASAP7_75t_L g1029 ( 
.A(n_908),
.B(n_559),
.Y(n_1029)
);

INVx2_ASAP7_75t_L g1030 ( 
.A(n_929),
.Y(n_1030)
);

NAND2xp33_ASAP7_75t_L g1031 ( 
.A(n_908),
.B(n_562),
.Y(n_1031)
);

BUFx6f_ASAP7_75t_L g1032 ( 
.A(n_898),
.Y(n_1032)
);

INVx2_ASAP7_75t_L g1033 ( 
.A(n_929),
.Y(n_1033)
);

AND2x2_ASAP7_75t_L g1034 ( 
.A(n_951),
.B(n_783),
.Y(n_1034)
);

NAND2xp5_ASAP7_75t_L g1035 ( 
.A(n_958),
.B(n_874),
.Y(n_1035)
);

NAND2xp5_ASAP7_75t_SL g1036 ( 
.A(n_951),
.B(n_563),
.Y(n_1036)
);

INVx2_ASAP7_75t_L g1037 ( 
.A(n_899),
.Y(n_1037)
);

BUFx6f_ASAP7_75t_L g1038 ( 
.A(n_898),
.Y(n_1038)
);

INVx1_ASAP7_75t_L g1039 ( 
.A(n_946),
.Y(n_1039)
);

INVx2_ASAP7_75t_L g1040 ( 
.A(n_899),
.Y(n_1040)
);

NOR2xp33_ASAP7_75t_L g1041 ( 
.A(n_906),
.B(n_740),
.Y(n_1041)
);

NAND2xp5_ASAP7_75t_L g1042 ( 
.A(n_912),
.B(n_915),
.Y(n_1042)
);

AND2x2_ASAP7_75t_L g1043 ( 
.A(n_946),
.B(n_869),
.Y(n_1043)
);

NAND2xp33_ASAP7_75t_L g1044 ( 
.A(n_911),
.B(n_564),
.Y(n_1044)
);

AND2x6_ASAP7_75t_L g1045 ( 
.A(n_911),
.B(n_665),
.Y(n_1045)
);

OR2x6_ASAP7_75t_L g1046 ( 
.A(n_913),
.B(n_869),
.Y(n_1046)
);

INVx2_ASAP7_75t_L g1047 ( 
.A(n_902),
.Y(n_1047)
);

NAND2xp5_ASAP7_75t_L g1048 ( 
.A(n_927),
.B(n_864),
.Y(n_1048)
);

INVx1_ASAP7_75t_L g1049 ( 
.A(n_903),
.Y(n_1049)
);

NOR2xp33_ASAP7_75t_L g1050 ( 
.A(n_913),
.B(n_743),
.Y(n_1050)
);

NAND2xp5_ASAP7_75t_L g1051 ( 
.A(n_916),
.B(n_867),
.Y(n_1051)
);

NOR2x1p5_ASAP7_75t_L g1052 ( 
.A(n_916),
.B(n_522),
.Y(n_1052)
);

NAND2xp5_ASAP7_75t_L g1053 ( 
.A(n_917),
.B(n_886),
.Y(n_1053)
);

NAND2xp5_ASAP7_75t_L g1054 ( 
.A(n_886),
.B(n_867),
.Y(n_1054)
);

INVx2_ASAP7_75t_L g1055 ( 
.A(n_886),
.Y(n_1055)
);

NOR2xp67_ASAP7_75t_L g1056 ( 
.A(n_904),
.B(n_870),
.Y(n_1056)
);

INVx1_ASAP7_75t_L g1057 ( 
.A(n_904),
.Y(n_1057)
);

INVx1_ASAP7_75t_L g1058 ( 
.A(n_907),
.Y(n_1058)
);

INVx1_ASAP7_75t_L g1059 ( 
.A(n_907),
.Y(n_1059)
);

NAND3xp33_ASAP7_75t_L g1060 ( 
.A(n_907),
.B(n_818),
.C(n_530),
.Y(n_1060)
);

NAND2xp33_ASAP7_75t_L g1061 ( 
.A(n_898),
.B(n_565),
.Y(n_1061)
);

INVx2_ASAP7_75t_L g1062 ( 
.A(n_924),
.Y(n_1062)
);

NAND2xp5_ASAP7_75t_L g1063 ( 
.A(n_924),
.B(n_870),
.Y(n_1063)
);

INVx8_ASAP7_75t_L g1064 ( 
.A(n_898),
.Y(n_1064)
);

BUFx5_ASAP7_75t_L g1065 ( 
.A(n_924),
.Y(n_1065)
);

NAND2xp5_ASAP7_75t_SL g1066 ( 
.A(n_910),
.B(n_568),
.Y(n_1066)
);

INVx2_ASAP7_75t_L g1067 ( 
.A(n_931),
.Y(n_1067)
);

INVx2_ASAP7_75t_L g1068 ( 
.A(n_931),
.Y(n_1068)
);

NAND2xp5_ASAP7_75t_L g1069 ( 
.A(n_910),
.B(n_875),
.Y(n_1069)
);

NAND2xp5_ASAP7_75t_L g1070 ( 
.A(n_910),
.B(n_875),
.Y(n_1070)
);

NOR2xp33_ASAP7_75t_L g1071 ( 
.A(n_910),
.B(n_749),
.Y(n_1071)
);

NAND2xp5_ASAP7_75t_L g1072 ( 
.A(n_910),
.B(n_877),
.Y(n_1072)
);

INVx2_ASAP7_75t_L g1073 ( 
.A(n_936),
.Y(n_1073)
);

BUFx2_ASAP7_75t_L g1074 ( 
.A(n_920),
.Y(n_1074)
);

INVxp67_ASAP7_75t_SL g1075 ( 
.A(n_920),
.Y(n_1075)
);

INVx2_ASAP7_75t_L g1076 ( 
.A(n_936),
.Y(n_1076)
);

NOR2xp33_ASAP7_75t_L g1077 ( 
.A(n_920),
.B(n_749),
.Y(n_1077)
);

AND2x2_ASAP7_75t_L g1078 ( 
.A(n_920),
.B(n_877),
.Y(n_1078)
);

AOI221xp5_ASAP7_75t_L g1079 ( 
.A1(n_920),
.A2(n_657),
.B1(n_534),
.B2(n_543),
.C(n_536),
.Y(n_1079)
);

NAND2xp33_ASAP7_75t_SL g1080 ( 
.A(n_925),
.B(n_579),
.Y(n_1080)
);

INVx2_ASAP7_75t_L g1081 ( 
.A(n_1023),
.Y(n_1081)
);

NAND2xp5_ASAP7_75t_L g1082 ( 
.A(n_964),
.B(n_925),
.Y(n_1082)
);

OAI22xp33_ASAP7_75t_SL g1083 ( 
.A1(n_971),
.A2(n_552),
.B1(n_566),
.B2(n_523),
.Y(n_1083)
);

NAND2x1p5_ASAP7_75t_L g1084 ( 
.A(n_1007),
.B(n_854),
.Y(n_1084)
);

AO22x2_ASAP7_75t_L g1085 ( 
.A1(n_1001),
.A2(n_752),
.B1(n_759),
.B2(n_758),
.Y(n_1085)
);

INVx1_ASAP7_75t_L g1086 ( 
.A(n_1043),
.Y(n_1086)
);

INVx1_ASAP7_75t_L g1087 ( 
.A(n_1049),
.Y(n_1087)
);

CKINVDCx20_ASAP7_75t_R g1088 ( 
.A(n_985),
.Y(n_1088)
);

OR2x6_ASAP7_75t_L g1089 ( 
.A(n_988),
.B(n_751),
.Y(n_1089)
);

INVx1_ASAP7_75t_L g1090 ( 
.A(n_1030),
.Y(n_1090)
);

NAND2xp5_ASAP7_75t_L g1091 ( 
.A(n_965),
.B(n_925),
.Y(n_1091)
);

INVx1_ASAP7_75t_L g1092 ( 
.A(n_1033),
.Y(n_1092)
);

AOI22xp5_ASAP7_75t_L g1093 ( 
.A1(n_982),
.A2(n_701),
.B1(n_688),
.B2(n_685),
.Y(n_1093)
);

AND2x2_ASAP7_75t_L g1094 ( 
.A(n_1022),
.B(n_752),
.Y(n_1094)
);

INVx1_ASAP7_75t_L g1095 ( 
.A(n_962),
.Y(n_1095)
);

CKINVDCx20_ASAP7_75t_R g1096 ( 
.A(n_1004),
.Y(n_1096)
);

INVx1_ASAP7_75t_L g1097 ( 
.A(n_966),
.Y(n_1097)
);

NOR2xp33_ASAP7_75t_L g1098 ( 
.A(n_1003),
.B(n_758),
.Y(n_1098)
);

AND2x2_ASAP7_75t_L g1099 ( 
.A(n_1034),
.B(n_989),
.Y(n_1099)
);

INVx1_ASAP7_75t_L g1100 ( 
.A(n_968),
.Y(n_1100)
);

AND2x6_ASAP7_75t_L g1101 ( 
.A(n_1007),
.B(n_1009),
.Y(n_1101)
);

INVx1_ASAP7_75t_L g1102 ( 
.A(n_969),
.Y(n_1102)
);

NOR2xp33_ASAP7_75t_L g1103 ( 
.A(n_961),
.B(n_759),
.Y(n_1103)
);

BUFx3_ASAP7_75t_L g1104 ( 
.A(n_991),
.Y(n_1104)
);

INVx1_ASAP7_75t_L g1105 ( 
.A(n_983),
.Y(n_1105)
);

NAND2x1p5_ASAP7_75t_L g1106 ( 
.A(n_1007),
.B(n_854),
.Y(n_1106)
);

AO22x2_ASAP7_75t_L g1107 ( 
.A1(n_999),
.A2(n_813),
.B1(n_791),
.B2(n_686),
.Y(n_1107)
);

NAND2xp5_ASAP7_75t_SL g1108 ( 
.A(n_1009),
.B(n_587),
.Y(n_1108)
);

AO22x2_ASAP7_75t_L g1109 ( 
.A1(n_960),
.A2(n_813),
.B1(n_791),
.B2(n_687),
.Y(n_1109)
);

INVx1_ASAP7_75t_L g1110 ( 
.A(n_998),
.Y(n_1110)
);

INVxp67_ASAP7_75t_L g1111 ( 
.A(n_1050),
.Y(n_1111)
);

AND2x4_ASAP7_75t_L g1112 ( 
.A(n_1052),
.B(n_753),
.Y(n_1112)
);

INVx1_ASAP7_75t_L g1113 ( 
.A(n_1048),
.Y(n_1113)
);

INVx1_ASAP7_75t_L g1114 ( 
.A(n_1051),
.Y(n_1114)
);

AO22x2_ASAP7_75t_L g1115 ( 
.A1(n_1006),
.A2(n_994),
.B1(n_992),
.B2(n_1026),
.Y(n_1115)
);

NOR2xp33_ASAP7_75t_L g1116 ( 
.A(n_1000),
.B(n_567),
.Y(n_1116)
);

CKINVDCx20_ASAP7_75t_R g1117 ( 
.A(n_1006),
.Y(n_1117)
);

INVx1_ASAP7_75t_L g1118 ( 
.A(n_1037),
.Y(n_1118)
);

INVx1_ASAP7_75t_L g1119 ( 
.A(n_1040),
.Y(n_1119)
);

BUFx2_ASAP7_75t_L g1120 ( 
.A(n_1009),
.Y(n_1120)
);

AND2x2_ASAP7_75t_L g1121 ( 
.A(n_971),
.B(n_854),
.Y(n_1121)
);

INVx1_ASAP7_75t_L g1122 ( 
.A(n_1047),
.Y(n_1122)
);

NAND2xp5_ASAP7_75t_L g1123 ( 
.A(n_1012),
.B(n_925),
.Y(n_1123)
);

AND2x2_ASAP7_75t_L g1124 ( 
.A(n_1071),
.B(n_854),
.Y(n_1124)
);

INVx1_ASAP7_75t_L g1125 ( 
.A(n_1039),
.Y(n_1125)
);

AND2x4_ASAP7_75t_L g1126 ( 
.A(n_1046),
.B(n_754),
.Y(n_1126)
);

INVx2_ASAP7_75t_L g1127 ( 
.A(n_963),
.Y(n_1127)
);

OR2x2_ASAP7_75t_SL g1128 ( 
.A(n_973),
.B(n_756),
.Y(n_1128)
);

AND2x4_ASAP7_75t_L g1129 ( 
.A(n_1077),
.B(n_760),
.Y(n_1129)
);

INVx2_ASAP7_75t_L g1130 ( 
.A(n_970),
.Y(n_1130)
);

AO22x2_ASAP7_75t_L g1131 ( 
.A1(n_987),
.A2(n_693),
.B1(n_700),
.B2(n_680),
.Y(n_1131)
);

AND2x2_ASAP7_75t_L g1132 ( 
.A(n_1041),
.B(n_996),
.Y(n_1132)
);

NAND2xp5_ASAP7_75t_L g1133 ( 
.A(n_984),
.B(n_936),
.Y(n_1133)
);

INVx1_ASAP7_75t_L g1134 ( 
.A(n_972),
.Y(n_1134)
);

INVx2_ASAP7_75t_L g1135 ( 
.A(n_977),
.Y(n_1135)
);

INVx2_ASAP7_75t_L g1136 ( 
.A(n_1002),
.Y(n_1136)
);

AND2x2_ASAP7_75t_L g1137 ( 
.A(n_1016),
.B(n_765),
.Y(n_1137)
);

INVx1_ASAP7_75t_L g1138 ( 
.A(n_1011),
.Y(n_1138)
);

INVx3_ASAP7_75t_L g1139 ( 
.A(n_1046),
.Y(n_1139)
);

INVx1_ASAP7_75t_L g1140 ( 
.A(n_1018),
.Y(n_1140)
);

AND2x4_ASAP7_75t_L g1141 ( 
.A(n_1046),
.B(n_1008),
.Y(n_1141)
);

AO22x2_ASAP7_75t_L g1142 ( 
.A1(n_988),
.A2(n_707),
.B1(n_710),
.B2(n_703),
.Y(n_1142)
);

INVx2_ASAP7_75t_SL g1143 ( 
.A(n_1010),
.Y(n_1143)
);

INVx1_ASAP7_75t_L g1144 ( 
.A(n_1054),
.Y(n_1144)
);

INVx1_ASAP7_75t_L g1145 ( 
.A(n_1063),
.Y(n_1145)
);

INVx1_ASAP7_75t_L g1146 ( 
.A(n_1078),
.Y(n_1146)
);

NAND2xp5_ASAP7_75t_L g1147 ( 
.A(n_975),
.B(n_936),
.Y(n_1147)
);

NAND2xp5_ASAP7_75t_L g1148 ( 
.A(n_993),
.B(n_936),
.Y(n_1148)
);

INVxp67_ASAP7_75t_L g1149 ( 
.A(n_1024),
.Y(n_1149)
);

INVx1_ASAP7_75t_L g1150 ( 
.A(n_1069),
.Y(n_1150)
);

INVx1_ASAP7_75t_L g1151 ( 
.A(n_1070),
.Y(n_1151)
);

AND2x4_ASAP7_75t_L g1152 ( 
.A(n_1005),
.B(n_769),
.Y(n_1152)
);

AND2x2_ASAP7_75t_L g1153 ( 
.A(n_1079),
.B(n_770),
.Y(n_1153)
);

INVx1_ASAP7_75t_L g1154 ( 
.A(n_1072),
.Y(n_1154)
);

NOR2x1p5_ASAP7_75t_L g1155 ( 
.A(n_978),
.B(n_569),
.Y(n_1155)
);

OAI221xp5_ASAP7_75t_L g1156 ( 
.A1(n_1014),
.A2(n_576),
.B1(n_577),
.B2(n_572),
.C(n_570),
.Y(n_1156)
);

CKINVDCx20_ASAP7_75t_R g1157 ( 
.A(n_1080),
.Y(n_1157)
);

NAND2xp5_ASAP7_75t_SL g1158 ( 
.A(n_980),
.B(n_588),
.Y(n_1158)
);

INVx1_ASAP7_75t_L g1159 ( 
.A(n_1057),
.Y(n_1159)
);

INVx1_ASAP7_75t_L g1160 ( 
.A(n_1058),
.Y(n_1160)
);

NAND2x1p5_ASAP7_75t_L g1161 ( 
.A(n_1074),
.B(n_826),
.Y(n_1161)
);

NAND2xp5_ASAP7_75t_L g1162 ( 
.A(n_993),
.B(n_726),
.Y(n_1162)
);

NAND2xp5_ASAP7_75t_L g1163 ( 
.A(n_974),
.B(n_826),
.Y(n_1163)
);

INVx1_ASAP7_75t_L g1164 ( 
.A(n_1059),
.Y(n_1164)
);

INVx2_ASAP7_75t_L g1165 ( 
.A(n_997),
.Y(n_1165)
);

INVx2_ASAP7_75t_SL g1166 ( 
.A(n_988),
.Y(n_1166)
);

INVx1_ASAP7_75t_L g1167 ( 
.A(n_1042),
.Y(n_1167)
);

INVx1_ASAP7_75t_L g1168 ( 
.A(n_981),
.Y(n_1168)
);

INVx1_ASAP7_75t_L g1169 ( 
.A(n_1055),
.Y(n_1169)
);

INVx3_ASAP7_75t_L g1170 ( 
.A(n_1062),
.Y(n_1170)
);

OAI22xp5_ASAP7_75t_L g1171 ( 
.A1(n_976),
.A2(n_599),
.B1(n_603),
.B2(n_592),
.Y(n_1171)
);

HB1xp67_ASAP7_75t_L g1172 ( 
.A(n_1014),
.Y(n_1172)
);

AND2x4_ASAP7_75t_L g1173 ( 
.A(n_1060),
.B(n_771),
.Y(n_1173)
);

INVx2_ASAP7_75t_L g1174 ( 
.A(n_1067),
.Y(n_1174)
);

AO22x2_ASAP7_75t_L g1175 ( 
.A1(n_1036),
.A2(n_776),
.B1(n_778),
.B2(n_775),
.Y(n_1175)
);

AO22x2_ASAP7_75t_L g1176 ( 
.A1(n_1028),
.A2(n_780),
.B1(n_779),
.B2(n_9),
.Y(n_1176)
);

AND2x2_ASAP7_75t_L g1177 ( 
.A(n_979),
.B(n_840),
.Y(n_1177)
);

NAND2xp5_ASAP7_75t_L g1178 ( 
.A(n_976),
.B(n_827),
.Y(n_1178)
);

NAND2xp5_ASAP7_75t_L g1179 ( 
.A(n_1021),
.B(n_827),
.Y(n_1179)
);

BUFx8_ASAP7_75t_L g1180 ( 
.A(n_1045),
.Y(n_1180)
);

BUFx8_ASAP7_75t_L g1181 ( 
.A(n_1045),
.Y(n_1181)
);

INVx3_ASAP7_75t_L g1182 ( 
.A(n_1068),
.Y(n_1182)
);

AND2x2_ASAP7_75t_L g1183 ( 
.A(n_979),
.B(n_843),
.Y(n_1183)
);

AO22x2_ASAP7_75t_L g1184 ( 
.A1(n_990),
.A2(n_2),
.B1(n_0),
.B2(n_1),
.Y(n_1184)
);

NAND2xp5_ASAP7_75t_L g1185 ( 
.A(n_1075),
.B(n_829),
.Y(n_1185)
);

AO22x2_ASAP7_75t_L g1186 ( 
.A1(n_995),
.A2(n_4),
.B1(n_1),
.B2(n_2),
.Y(n_1186)
);

INVx2_ASAP7_75t_SL g1187 ( 
.A(n_1045),
.Y(n_1187)
);

INVx1_ASAP7_75t_L g1188 ( 
.A(n_1017),
.Y(n_1188)
);

INVxp67_ASAP7_75t_SL g1189 ( 
.A(n_1032),
.Y(n_1189)
);

INVx1_ASAP7_75t_L g1190 ( 
.A(n_1019),
.Y(n_1190)
);

AO22x2_ASAP7_75t_L g1191 ( 
.A1(n_1073),
.A2(n_1076),
.B1(n_1066),
.B2(n_14),
.Y(n_1191)
);

INVx1_ASAP7_75t_SL g1192 ( 
.A(n_1025),
.Y(n_1192)
);

INVxp67_ASAP7_75t_L g1193 ( 
.A(n_1045),
.Y(n_1193)
);

INVx2_ASAP7_75t_L g1194 ( 
.A(n_986),
.Y(n_1194)
);

AND2x2_ASAP7_75t_L g1195 ( 
.A(n_967),
.B(n_840),
.Y(n_1195)
);

AO22x2_ASAP7_75t_L g1196 ( 
.A1(n_1053),
.A2(n_6),
.B1(n_4),
.B2(n_5),
.Y(n_1196)
);

AOI22xp5_ASAP7_75t_L g1197 ( 
.A1(n_1029),
.A2(n_606),
.B1(n_625),
.B2(n_605),
.Y(n_1197)
);

INVx1_ASAP7_75t_L g1198 ( 
.A(n_1035),
.Y(n_1198)
);

INVx1_ASAP7_75t_L g1199 ( 
.A(n_1013),
.Y(n_1199)
);

INVx1_ASAP7_75t_L g1200 ( 
.A(n_1015),
.Y(n_1200)
);

AO22x2_ASAP7_75t_L g1201 ( 
.A1(n_1020),
.A2(n_7),
.B1(n_5),
.B2(n_6),
.Y(n_1201)
);

INVx1_ASAP7_75t_L g1202 ( 
.A(n_1056),
.Y(n_1202)
);

AOI22xp5_ASAP7_75t_L g1203 ( 
.A1(n_1031),
.A2(n_629),
.B1(n_630),
.B2(n_628),
.Y(n_1203)
);

AO22x2_ASAP7_75t_L g1204 ( 
.A1(n_986),
.A2(n_9),
.B1(n_7),
.B2(n_8),
.Y(n_1204)
);

INVx1_ASAP7_75t_L g1205 ( 
.A(n_986),
.Y(n_1205)
);

BUFx8_ASAP7_75t_L g1206 ( 
.A(n_1032),
.Y(n_1206)
);

INVx1_ASAP7_75t_L g1207 ( 
.A(n_1032),
.Y(n_1207)
);

AO22x2_ASAP7_75t_L g1208 ( 
.A1(n_1044),
.A2(n_13),
.B1(n_8),
.B2(n_12),
.Y(n_1208)
);

NAND2x1p5_ASAP7_75t_L g1209 ( 
.A(n_1038),
.B(n_829),
.Y(n_1209)
);

INVx1_ASAP7_75t_L g1210 ( 
.A(n_1038),
.Y(n_1210)
);

OAI22xp5_ASAP7_75t_SL g1211 ( 
.A1(n_1061),
.A2(n_583),
.B1(n_585),
.B2(n_582),
.Y(n_1211)
);

NOR2xp33_ASAP7_75t_SL g1212 ( 
.A(n_1064),
.B(n_555),
.Y(n_1212)
);

NAND2xp33_ASAP7_75t_L g1213 ( 
.A(n_1065),
.B(n_631),
.Y(n_1213)
);

AO22x2_ASAP7_75t_L g1214 ( 
.A1(n_1065),
.A2(n_14),
.B1(n_12),
.B2(n_13),
.Y(n_1214)
);

INVx1_ASAP7_75t_L g1215 ( 
.A(n_1064),
.Y(n_1215)
);

AND2x2_ASAP7_75t_L g1216 ( 
.A(n_1064),
.B(n_586),
.Y(n_1216)
);

AO22x2_ASAP7_75t_L g1217 ( 
.A1(n_1001),
.A2(n_17),
.B1(n_15),
.B2(n_16),
.Y(n_1217)
);

AOI22xp5_ASAP7_75t_L g1218 ( 
.A1(n_982),
.A2(n_638),
.B1(n_645),
.B2(n_636),
.Y(n_1218)
);

NAND2x1p5_ASAP7_75t_L g1219 ( 
.A(n_1007),
.B(n_832),
.Y(n_1219)
);

AND2x4_ASAP7_75t_L g1220 ( 
.A(n_998),
.B(n_832),
.Y(n_1220)
);

NAND2xp5_ASAP7_75t_L g1221 ( 
.A(n_964),
.B(n_837),
.Y(n_1221)
);

INVx1_ASAP7_75t_L g1222 ( 
.A(n_1027),
.Y(n_1222)
);

AO22x2_ASAP7_75t_L g1223 ( 
.A1(n_1001),
.A2(n_18),
.B1(n_15),
.B2(n_17),
.Y(n_1223)
);

INVx1_ASAP7_75t_L g1224 ( 
.A(n_1027),
.Y(n_1224)
);

NAND2x1p5_ASAP7_75t_L g1225 ( 
.A(n_1007),
.B(n_837),
.Y(n_1225)
);

INVx1_ASAP7_75t_L g1226 ( 
.A(n_1027),
.Y(n_1226)
);

AOI22xp5_ASAP7_75t_L g1227 ( 
.A1(n_982),
.A2(n_658),
.B1(n_659),
.B2(n_648),
.Y(n_1227)
);

INVx1_ASAP7_75t_L g1228 ( 
.A(n_1027),
.Y(n_1228)
);

AND2x4_ASAP7_75t_L g1229 ( 
.A(n_985),
.B(n_595),
.Y(n_1229)
);

INVx1_ASAP7_75t_L g1230 ( 
.A(n_1027),
.Y(n_1230)
);

INVx1_ASAP7_75t_L g1231 ( 
.A(n_1027),
.Y(n_1231)
);

NAND2xp5_ASAP7_75t_L g1232 ( 
.A(n_964),
.B(n_660),
.Y(n_1232)
);

BUFx6f_ASAP7_75t_L g1233 ( 
.A(n_985),
.Y(n_1233)
);

HB1xp67_ASAP7_75t_L g1234 ( 
.A(n_965),
.Y(n_1234)
);

INVx1_ASAP7_75t_L g1235 ( 
.A(n_1027),
.Y(n_1235)
);

NAND2xp5_ASAP7_75t_L g1236 ( 
.A(n_964),
.B(n_662),
.Y(n_1236)
);

AND2x4_ASAP7_75t_L g1237 ( 
.A(n_998),
.B(n_222),
.Y(n_1237)
);

INVx2_ASAP7_75t_SL g1238 ( 
.A(n_1052),
.Y(n_1238)
);

INVx2_ASAP7_75t_L g1239 ( 
.A(n_1023),
.Y(n_1239)
);

AOI22xp5_ASAP7_75t_L g1240 ( 
.A1(n_982),
.A2(n_667),
.B1(n_671),
.B2(n_663),
.Y(n_1240)
);

INVx1_ASAP7_75t_L g1241 ( 
.A(n_1027),
.Y(n_1241)
);

NAND2x1p5_ASAP7_75t_L g1242 ( 
.A(n_1007),
.B(n_518),
.Y(n_1242)
);

CKINVDCx14_ASAP7_75t_R g1243 ( 
.A(n_985),
.Y(n_1243)
);

AO22x2_ASAP7_75t_L g1244 ( 
.A1(n_1001),
.A2(n_20),
.B1(n_18),
.B2(n_19),
.Y(n_1244)
);

AND2x4_ASAP7_75t_L g1245 ( 
.A(n_998),
.B(n_225),
.Y(n_1245)
);

NAND3xp33_ASAP7_75t_SL g1246 ( 
.A(n_1006),
.B(n_598),
.C(n_596),
.Y(n_1246)
);

INVx1_ASAP7_75t_L g1247 ( 
.A(n_1027),
.Y(n_1247)
);

INVx2_ASAP7_75t_L g1248 ( 
.A(n_1023),
.Y(n_1248)
);

NOR2xp67_ASAP7_75t_L g1249 ( 
.A(n_1003),
.B(n_672),
.Y(n_1249)
);

INVx1_ASAP7_75t_L g1250 ( 
.A(n_1027),
.Y(n_1250)
);

AO22x2_ASAP7_75t_L g1251 ( 
.A1(n_1001),
.A2(n_21),
.B1(n_19),
.B2(n_20),
.Y(n_1251)
);

INVx1_ASAP7_75t_L g1252 ( 
.A(n_1027),
.Y(n_1252)
);

NAND2xp5_ASAP7_75t_L g1253 ( 
.A(n_964),
.B(n_674),
.Y(n_1253)
);

AOI22xp33_ASAP7_75t_L g1254 ( 
.A1(n_1012),
.A2(n_556),
.B1(n_581),
.B2(n_518),
.Y(n_1254)
);

NAND2xp5_ASAP7_75t_L g1255 ( 
.A(n_1099),
.B(n_682),
.Y(n_1255)
);

INVx1_ASAP7_75t_L g1256 ( 
.A(n_1095),
.Y(n_1256)
);

NAND2xp5_ASAP7_75t_L g1257 ( 
.A(n_1086),
.B(n_689),
.Y(n_1257)
);

OAI321xp33_ASAP7_75t_L g1258 ( 
.A1(n_1093),
.A2(n_613),
.A3(n_581),
.B1(n_556),
.B2(n_615),
.C(n_612),
.Y(n_1258)
);

NAND2xp5_ASAP7_75t_L g1259 ( 
.A(n_1192),
.B(n_690),
.Y(n_1259)
);

INVx1_ASAP7_75t_L g1260 ( 
.A(n_1097),
.Y(n_1260)
);

OAI22x1_ASAP7_75t_L g1261 ( 
.A1(n_1103),
.A2(n_624),
.B1(n_635),
.B2(n_619),
.Y(n_1261)
);

INVx1_ASAP7_75t_L g1262 ( 
.A(n_1100),
.Y(n_1262)
);

AOI21x1_ASAP7_75t_L g1263 ( 
.A1(n_1082),
.A2(n_581),
.B(n_556),
.Y(n_1263)
);

NAND3xp33_ASAP7_75t_L g1264 ( 
.A(n_1098),
.B(n_643),
.C(n_639),
.Y(n_1264)
);

AO21x1_ASAP7_75t_L g1265 ( 
.A1(n_1147),
.A2(n_613),
.B(n_22),
.Y(n_1265)
);

AOI21xp5_ASAP7_75t_L g1266 ( 
.A1(n_1133),
.A2(n_613),
.B(n_692),
.Y(n_1266)
);

O2A1O1Ixp33_ASAP7_75t_L g1267 ( 
.A1(n_1111),
.A2(n_649),
.B(n_653),
.C(n_644),
.Y(n_1267)
);

NAND2xp5_ASAP7_75t_L g1268 ( 
.A(n_1113),
.B(n_695),
.Y(n_1268)
);

BUFx12f_ASAP7_75t_L g1269 ( 
.A(n_1233),
.Y(n_1269)
);

NOR2xp67_ASAP7_75t_L g1270 ( 
.A(n_1149),
.B(n_698),
.Y(n_1270)
);

AOI21xp5_ASAP7_75t_L g1271 ( 
.A1(n_1213),
.A2(n_613),
.B(n_704),
.Y(n_1271)
);

AND2x2_ASAP7_75t_L g1272 ( 
.A(n_1234),
.B(n_669),
.Y(n_1272)
);

AOI21xp5_ASAP7_75t_L g1273 ( 
.A1(n_1178),
.A2(n_713),
.B(n_709),
.Y(n_1273)
);

BUFx8_ASAP7_75t_L g1274 ( 
.A(n_1233),
.Y(n_1274)
);

AOI22xp33_ASAP7_75t_L g1275 ( 
.A1(n_1246),
.A2(n_719),
.B1(n_720),
.B2(n_714),
.Y(n_1275)
);

NAND2xp5_ASAP7_75t_L g1276 ( 
.A(n_1221),
.B(n_723),
.Y(n_1276)
);

AND2x2_ASAP7_75t_L g1277 ( 
.A(n_1132),
.B(n_676),
.Y(n_1277)
);

NAND2xp5_ASAP7_75t_SL g1278 ( 
.A(n_1141),
.B(n_724),
.Y(n_1278)
);

AOI22xp33_ASAP7_75t_L g1279 ( 
.A1(n_1153),
.A2(n_1131),
.B1(n_1121),
.B2(n_1172),
.Y(n_1279)
);

NAND2xp5_ASAP7_75t_SL g1280 ( 
.A(n_1141),
.B(n_725),
.Y(n_1280)
);

AND2x4_ASAP7_75t_L g1281 ( 
.A(n_1120),
.B(n_226),
.Y(n_1281)
);

NAND2xp5_ASAP7_75t_L g1282 ( 
.A(n_1232),
.B(n_696),
.Y(n_1282)
);

AND2x4_ASAP7_75t_SL g1283 ( 
.A(n_1088),
.B(n_227),
.Y(n_1283)
);

OAI22xp5_ASAP7_75t_L g1284 ( 
.A1(n_1236),
.A2(n_705),
.B1(n_712),
.B2(n_699),
.Y(n_1284)
);

NOR3xp33_ASAP7_75t_L g1285 ( 
.A(n_1083),
.B(n_722),
.C(n_715),
.Y(n_1285)
);

HB1xp67_ASAP7_75t_L g1286 ( 
.A(n_1104),
.Y(n_1286)
);

INVx1_ASAP7_75t_L g1287 ( 
.A(n_1102),
.Y(n_1287)
);

AOI21xp5_ASAP7_75t_L g1288 ( 
.A1(n_1148),
.A2(n_230),
.B(n_229),
.Y(n_1288)
);

AOI22xp5_ASAP7_75t_L g1289 ( 
.A1(n_1143),
.A2(n_233),
.B1(n_236),
.B2(n_231),
.Y(n_1289)
);

O2A1O1Ixp5_ASAP7_75t_SL g1290 ( 
.A1(n_1158),
.A2(n_25),
.B(n_23),
.C(n_24),
.Y(n_1290)
);

BUFx2_ASAP7_75t_L g1291 ( 
.A(n_1096),
.Y(n_1291)
);

AOI22xp5_ASAP7_75t_L g1292 ( 
.A1(n_1253),
.A2(n_240),
.B1(n_241),
.B2(n_238),
.Y(n_1292)
);

OAI22xp5_ASAP7_75t_L g1293 ( 
.A1(n_1146),
.A2(n_243),
.B1(n_244),
.B2(n_242),
.Y(n_1293)
);

AOI21xp5_ASAP7_75t_L g1294 ( 
.A1(n_1163),
.A2(n_250),
.B(n_246),
.Y(n_1294)
);

AOI21xp5_ASAP7_75t_L g1295 ( 
.A1(n_1091),
.A2(n_253),
.B(n_251),
.Y(n_1295)
);

NAND2xp5_ASAP7_75t_L g1296 ( 
.A(n_1114),
.B(n_1198),
.Y(n_1296)
);

AOI21xp5_ASAP7_75t_L g1297 ( 
.A1(n_1123),
.A2(n_256),
.B(n_255),
.Y(n_1297)
);

NOR2xp33_ASAP7_75t_L g1298 ( 
.A(n_1094),
.B(n_23),
.Y(n_1298)
);

NAND2xp5_ASAP7_75t_SL g1299 ( 
.A(n_1120),
.B(n_1139),
.Y(n_1299)
);

A2O1A1Ixp33_ASAP7_75t_L g1300 ( 
.A1(n_1105),
.A2(n_27),
.B(n_25),
.C(n_26),
.Y(n_1300)
);

NAND2xp5_ASAP7_75t_L g1301 ( 
.A(n_1168),
.B(n_1199),
.Y(n_1301)
);

NAND2xp5_ASAP7_75t_SL g1302 ( 
.A(n_1249),
.B(n_257),
.Y(n_1302)
);

INVx1_ASAP7_75t_L g1303 ( 
.A(n_1087),
.Y(n_1303)
);

BUFx2_ASAP7_75t_L g1304 ( 
.A(n_1206),
.Y(n_1304)
);

NAND2xp5_ASAP7_75t_L g1305 ( 
.A(n_1200),
.B(n_26),
.Y(n_1305)
);

NOR2xp33_ASAP7_75t_L g1306 ( 
.A(n_1116),
.B(n_27),
.Y(n_1306)
);

AOI21xp5_ASAP7_75t_L g1307 ( 
.A1(n_1194),
.A2(n_260),
.B(n_258),
.Y(n_1307)
);

INVx1_ASAP7_75t_L g1308 ( 
.A(n_1110),
.Y(n_1308)
);

NAND2xp5_ASAP7_75t_L g1309 ( 
.A(n_1188),
.B(n_28),
.Y(n_1309)
);

AOI21xp5_ASAP7_75t_L g1310 ( 
.A1(n_1150),
.A2(n_263),
.B(n_262),
.Y(n_1310)
);

AOI21xp5_ASAP7_75t_L g1311 ( 
.A1(n_1151),
.A2(n_268),
.B(n_265),
.Y(n_1311)
);

INVx1_ASAP7_75t_L g1312 ( 
.A(n_1138),
.Y(n_1312)
);

HB1xp67_ASAP7_75t_L g1313 ( 
.A(n_1126),
.Y(n_1313)
);

BUFx6f_ASAP7_75t_L g1314 ( 
.A(n_1101),
.Y(n_1314)
);

BUFx3_ASAP7_75t_L g1315 ( 
.A(n_1229),
.Y(n_1315)
);

NOR2xp33_ASAP7_75t_L g1316 ( 
.A(n_1117),
.B(n_28),
.Y(n_1316)
);

OAI22x1_ASAP7_75t_L g1317 ( 
.A1(n_1166),
.A2(n_31),
.B1(n_29),
.B2(n_30),
.Y(n_1317)
);

NAND2xp5_ASAP7_75t_L g1318 ( 
.A(n_1190),
.B(n_30),
.Y(n_1318)
);

AOI21xp5_ASAP7_75t_L g1319 ( 
.A1(n_1154),
.A2(n_272),
.B(n_269),
.Y(n_1319)
);

AOI21xp5_ASAP7_75t_L g1320 ( 
.A1(n_1179),
.A2(n_274),
.B(n_273),
.Y(n_1320)
);

NAND2xp5_ASAP7_75t_L g1321 ( 
.A(n_1144),
.B(n_31),
.Y(n_1321)
);

O2A1O1Ixp33_ASAP7_75t_L g1322 ( 
.A1(n_1156),
.A2(n_34),
.B(n_32),
.C(n_33),
.Y(n_1322)
);

A2O1A1Ixp33_ASAP7_75t_L g1323 ( 
.A1(n_1145),
.A2(n_36),
.B(n_33),
.C(n_35),
.Y(n_1323)
);

AOI21xp5_ASAP7_75t_L g1324 ( 
.A1(n_1185),
.A2(n_279),
.B(n_277),
.Y(n_1324)
);

OAI22xp5_ASAP7_75t_L g1325 ( 
.A1(n_1205),
.A2(n_282),
.B1(n_284),
.B2(n_281),
.Y(n_1325)
);

BUFx6f_ASAP7_75t_L g1326 ( 
.A(n_1101),
.Y(n_1326)
);

NOR2xp33_ASAP7_75t_L g1327 ( 
.A(n_1129),
.B(n_35),
.Y(n_1327)
);

NAND2xp5_ASAP7_75t_L g1328 ( 
.A(n_1124),
.B(n_37),
.Y(n_1328)
);

O2A1O1Ixp33_ASAP7_75t_L g1329 ( 
.A1(n_1238),
.A2(n_39),
.B(n_37),
.C(n_38),
.Y(n_1329)
);

BUFx6f_ASAP7_75t_L g1330 ( 
.A(n_1101),
.Y(n_1330)
);

A2O1A1Ixp33_ASAP7_75t_L g1331 ( 
.A1(n_1237),
.A2(n_40),
.B(n_38),
.C(n_39),
.Y(n_1331)
);

NAND3xp33_ASAP7_75t_L g1332 ( 
.A(n_1218),
.B(n_40),
.C(n_41),
.Y(n_1332)
);

A2O1A1Ixp33_ASAP7_75t_L g1333 ( 
.A1(n_1237),
.A2(n_43),
.B(n_41),
.C(n_42),
.Y(n_1333)
);

NAND2xp5_ASAP7_75t_L g1334 ( 
.A(n_1152),
.B(n_42),
.Y(n_1334)
);

NAND2xp5_ASAP7_75t_L g1335 ( 
.A(n_1152),
.B(n_43),
.Y(n_1335)
);

INVx1_ASAP7_75t_L g1336 ( 
.A(n_1140),
.Y(n_1336)
);

CKINVDCx5p33_ASAP7_75t_R g1337 ( 
.A(n_1243),
.Y(n_1337)
);

INVx1_ASAP7_75t_L g1338 ( 
.A(n_1125),
.Y(n_1338)
);

OA22x2_ASAP7_75t_L g1339 ( 
.A1(n_1089),
.A2(n_47),
.B1(n_45),
.B2(n_46),
.Y(n_1339)
);

NAND2xp5_ASAP7_75t_SL g1340 ( 
.A(n_1126),
.B(n_295),
.Y(n_1340)
);

OR2x6_ASAP7_75t_L g1341 ( 
.A(n_1089),
.B(n_46),
.Y(n_1341)
);

OAI22xp5_ASAP7_75t_L g1342 ( 
.A1(n_1222),
.A2(n_1224),
.B1(n_1228),
.B2(n_1226),
.Y(n_1342)
);

NAND2xp5_ASAP7_75t_SL g1343 ( 
.A(n_1245),
.B(n_296),
.Y(n_1343)
);

NAND2xp5_ASAP7_75t_SL g1344 ( 
.A(n_1245),
.B(n_302),
.Y(n_1344)
);

AND2x2_ASAP7_75t_SL g1345 ( 
.A(n_1212),
.B(n_48),
.Y(n_1345)
);

NOR2xp33_ASAP7_75t_L g1346 ( 
.A(n_1128),
.B(n_49),
.Y(n_1346)
);

NAND3xp33_ASAP7_75t_L g1347 ( 
.A(n_1227),
.B(n_50),
.C(n_51),
.Y(n_1347)
);

NAND2xp5_ASAP7_75t_L g1348 ( 
.A(n_1230),
.B(n_50),
.Y(n_1348)
);

NAND2xp5_ASAP7_75t_L g1349 ( 
.A(n_1231),
.B(n_51),
.Y(n_1349)
);

AOI21xp5_ASAP7_75t_L g1350 ( 
.A1(n_1189),
.A2(n_1108),
.B(n_1202),
.Y(n_1350)
);

HB1xp67_ASAP7_75t_L g1351 ( 
.A(n_1220),
.Y(n_1351)
);

NAND2xp5_ASAP7_75t_L g1352 ( 
.A(n_1235),
.B(n_52),
.Y(n_1352)
);

O2A1O1Ixp5_ASAP7_75t_L g1353 ( 
.A1(n_1162),
.A2(n_305),
.B(n_306),
.C(n_303),
.Y(n_1353)
);

NAND2xp5_ASAP7_75t_L g1354 ( 
.A(n_1241),
.B(n_53),
.Y(n_1354)
);

NAND2xp5_ASAP7_75t_L g1355 ( 
.A(n_1247),
.B(n_53),
.Y(n_1355)
);

AOI22xp5_ASAP7_75t_L g1356 ( 
.A1(n_1155),
.A2(n_311),
.B1(n_312),
.B2(n_309),
.Y(n_1356)
);

AOI21x1_ASAP7_75t_L g1357 ( 
.A1(n_1165),
.A2(n_314),
.B(n_313),
.Y(n_1357)
);

INVx4_ASAP7_75t_L g1358 ( 
.A(n_1220),
.Y(n_1358)
);

NAND2xp5_ASAP7_75t_L g1359 ( 
.A(n_1250),
.B(n_54),
.Y(n_1359)
);

HB1xp67_ASAP7_75t_L g1360 ( 
.A(n_1112),
.Y(n_1360)
);

NOR2x1p5_ASAP7_75t_SL g1361 ( 
.A(n_1174),
.B(n_316),
.Y(n_1361)
);

BUFx6f_ASAP7_75t_L g1362 ( 
.A(n_1207),
.Y(n_1362)
);

OAI22xp5_ASAP7_75t_L g1363 ( 
.A1(n_1252),
.A2(n_320),
.B1(n_321),
.B2(n_319),
.Y(n_1363)
);

NAND2xp5_ASAP7_75t_L g1364 ( 
.A(n_1175),
.B(n_54),
.Y(n_1364)
);

O2A1O1Ixp5_ASAP7_75t_L g1365 ( 
.A1(n_1195),
.A2(n_327),
.B(n_328),
.C(n_325),
.Y(n_1365)
);

O2A1O1Ixp33_ASAP7_75t_L g1366 ( 
.A1(n_1118),
.A2(n_57),
.B(n_55),
.C(n_56),
.Y(n_1366)
);

OR2x6_ASAP7_75t_SL g1367 ( 
.A(n_1119),
.B(n_55),
.Y(n_1367)
);

OAI22x1_ASAP7_75t_L g1368 ( 
.A1(n_1112),
.A2(n_1107),
.B1(n_1085),
.B2(n_1109),
.Y(n_1368)
);

INVx5_ASAP7_75t_L g1369 ( 
.A(n_1216),
.Y(n_1369)
);

AOI22xp5_ASAP7_75t_L g1370 ( 
.A1(n_1115),
.A2(n_333),
.B1(n_334),
.B2(n_329),
.Y(n_1370)
);

A2O1A1Ixp33_ASAP7_75t_L g1371 ( 
.A1(n_1122),
.A2(n_60),
.B(n_56),
.C(n_59),
.Y(n_1371)
);

INVxp67_ASAP7_75t_L g1372 ( 
.A(n_1137),
.Y(n_1372)
);

BUFx2_ASAP7_75t_L g1373 ( 
.A(n_1115),
.Y(n_1373)
);

NOR2xp33_ASAP7_75t_L g1374 ( 
.A(n_1240),
.B(n_59),
.Y(n_1374)
);

AOI21xp5_ASAP7_75t_L g1375 ( 
.A1(n_1177),
.A2(n_337),
.B(n_336),
.Y(n_1375)
);

INVx3_ASAP7_75t_L g1376 ( 
.A(n_1084),
.Y(n_1376)
);

OR2x2_ASAP7_75t_L g1377 ( 
.A(n_1090),
.B(n_60),
.Y(n_1377)
);

AOI21xp5_ASAP7_75t_L g1378 ( 
.A1(n_1183),
.A2(n_342),
.B(n_338),
.Y(n_1378)
);

BUFx4f_ASAP7_75t_L g1379 ( 
.A(n_1161),
.Y(n_1379)
);

AOI21xp5_ASAP7_75t_L g1380 ( 
.A1(n_1210),
.A2(n_344),
.B(n_343),
.Y(n_1380)
);

NAND2xp5_ASAP7_75t_SL g1381 ( 
.A(n_1173),
.B(n_346),
.Y(n_1381)
);

OAI21xp5_ASAP7_75t_L g1382 ( 
.A1(n_1193),
.A2(n_1092),
.B(n_1134),
.Y(n_1382)
);

INVx3_ASAP7_75t_L g1383 ( 
.A(n_1106),
.Y(n_1383)
);

INVx2_ASAP7_75t_SL g1384 ( 
.A(n_1173),
.Y(n_1384)
);

BUFx2_ASAP7_75t_L g1385 ( 
.A(n_1085),
.Y(n_1385)
);

AOI21xp5_ASAP7_75t_L g1386 ( 
.A1(n_1219),
.A2(n_348),
.B(n_347),
.Y(n_1386)
);

NAND2xp5_ASAP7_75t_L g1387 ( 
.A(n_1081),
.B(n_61),
.Y(n_1387)
);

NAND2xp5_ASAP7_75t_L g1388 ( 
.A(n_1239),
.B(n_62),
.Y(n_1388)
);

OAI22xp33_ASAP7_75t_L g1389 ( 
.A1(n_1157),
.A2(n_1160),
.B1(n_1164),
.B2(n_1159),
.Y(n_1389)
);

OAI21xp33_ASAP7_75t_L g1390 ( 
.A1(n_1107),
.A2(n_62),
.B(n_63),
.Y(n_1390)
);

BUFx2_ASAP7_75t_SL g1391 ( 
.A(n_1215),
.Y(n_1391)
);

HB1xp67_ASAP7_75t_L g1392 ( 
.A(n_1248),
.Y(n_1392)
);

AOI22x1_ASAP7_75t_L g1393 ( 
.A1(n_1131),
.A2(n_352),
.B1(n_353),
.B2(n_349),
.Y(n_1393)
);

O2A1O1Ixp33_ASAP7_75t_SL g1394 ( 
.A1(n_1187),
.A2(n_355),
.B(n_356),
.C(n_354),
.Y(n_1394)
);

AOI21xp5_ASAP7_75t_L g1395 ( 
.A1(n_1225),
.A2(n_358),
.B(n_357),
.Y(n_1395)
);

BUFx12f_ASAP7_75t_L g1396 ( 
.A(n_1180),
.Y(n_1396)
);

AOI21xp5_ASAP7_75t_L g1397 ( 
.A1(n_1127),
.A2(n_1135),
.B(n_1130),
.Y(n_1397)
);

AOI22xp5_ASAP7_75t_L g1398 ( 
.A1(n_1171),
.A2(n_360),
.B1(n_361),
.B2(n_359),
.Y(n_1398)
);

INVxp67_ASAP7_75t_L g1399 ( 
.A(n_1109),
.Y(n_1399)
);

NAND2xp5_ASAP7_75t_L g1400 ( 
.A(n_1136),
.B(n_64),
.Y(n_1400)
);

BUFx4f_ASAP7_75t_L g1401 ( 
.A(n_1242),
.Y(n_1401)
);

BUFx8_ASAP7_75t_L g1402 ( 
.A(n_1169),
.Y(n_1402)
);

NAND2xp5_ASAP7_75t_L g1403 ( 
.A(n_1170),
.B(n_65),
.Y(n_1403)
);

NOR2x1_ASAP7_75t_L g1404 ( 
.A(n_1182),
.B(n_363),
.Y(n_1404)
);

NOR2xp33_ASAP7_75t_L g1405 ( 
.A(n_1211),
.B(n_67),
.Y(n_1405)
);

OAI22xp5_ASAP7_75t_L g1406 ( 
.A1(n_1191),
.A2(n_366),
.B1(n_367),
.B2(n_365),
.Y(n_1406)
);

NOR2xp33_ASAP7_75t_L g1407 ( 
.A(n_1197),
.B(n_1203),
.Y(n_1407)
);

NAND2xp5_ASAP7_75t_L g1408 ( 
.A(n_1176),
.B(n_67),
.Y(n_1408)
);

NAND2xp5_ASAP7_75t_L g1409 ( 
.A(n_1176),
.B(n_1191),
.Y(n_1409)
);

O2A1O1Ixp5_ASAP7_75t_L g1410 ( 
.A1(n_1217),
.A2(n_371),
.B(n_372),
.C(n_369),
.Y(n_1410)
);

OAI21xp5_ASAP7_75t_L g1411 ( 
.A1(n_1254),
.A2(n_374),
.B(n_373),
.Y(n_1411)
);

OAI21xp5_ASAP7_75t_L g1412 ( 
.A1(n_1209),
.A2(n_376),
.B(n_375),
.Y(n_1412)
);

INVx4_ASAP7_75t_L g1413 ( 
.A(n_1223),
.Y(n_1413)
);

AOI21xp5_ASAP7_75t_L g1414 ( 
.A1(n_1201),
.A2(n_381),
.B(n_378),
.Y(n_1414)
);

O2A1O1Ixp5_ASAP7_75t_L g1415 ( 
.A1(n_1223),
.A2(n_384),
.B(n_389),
.C(n_382),
.Y(n_1415)
);

NAND2xp5_ASAP7_75t_L g1416 ( 
.A(n_1142),
.B(n_69),
.Y(n_1416)
);

AOI21xp5_ASAP7_75t_L g1417 ( 
.A1(n_1201),
.A2(n_1251),
.B(n_1244),
.Y(n_1417)
);

NAND2xp5_ASAP7_75t_SL g1418 ( 
.A(n_1181),
.B(n_390),
.Y(n_1418)
);

AOI21xp33_ASAP7_75t_L g1419 ( 
.A1(n_1244),
.A2(n_69),
.B(n_70),
.Y(n_1419)
);

NOR2xp33_ASAP7_75t_L g1420 ( 
.A(n_1142),
.B(n_71),
.Y(n_1420)
);

BUFx12f_ASAP7_75t_L g1421 ( 
.A(n_1208),
.Y(n_1421)
);

NAND2xp5_ASAP7_75t_SL g1422 ( 
.A(n_1251),
.B(n_391),
.Y(n_1422)
);

NAND2xp5_ASAP7_75t_L g1423 ( 
.A(n_1208),
.B(n_71),
.Y(n_1423)
);

NAND2xp5_ASAP7_75t_L g1424 ( 
.A(n_1204),
.B(n_72),
.Y(n_1424)
);

NAND2xp5_ASAP7_75t_L g1425 ( 
.A(n_1204),
.B(n_73),
.Y(n_1425)
);

BUFx2_ASAP7_75t_L g1426 ( 
.A(n_1196),
.Y(n_1426)
);

NOR2xp33_ASAP7_75t_L g1427 ( 
.A(n_1184),
.B(n_73),
.Y(n_1427)
);

NAND2xp5_ASAP7_75t_L g1428 ( 
.A(n_1186),
.B(n_74),
.Y(n_1428)
);

INVx1_ASAP7_75t_L g1429 ( 
.A(n_1214),
.Y(n_1429)
);

INVx5_ASAP7_75t_L g1430 ( 
.A(n_1214),
.Y(n_1430)
);

AOI21xp5_ASAP7_75t_L g1431 ( 
.A1(n_1186),
.A2(n_393),
.B(n_392),
.Y(n_1431)
);

NAND2xp5_ASAP7_75t_L g1432 ( 
.A(n_1184),
.B(n_74),
.Y(n_1432)
);

NAND2xp5_ASAP7_75t_L g1433 ( 
.A(n_1196),
.B(n_76),
.Y(n_1433)
);

AND2x2_ASAP7_75t_L g1434 ( 
.A(n_1234),
.B(n_76),
.Y(n_1434)
);

NAND2xp5_ASAP7_75t_L g1435 ( 
.A(n_1167),
.B(n_77),
.Y(n_1435)
);

INVx1_ASAP7_75t_L g1436 ( 
.A(n_1095),
.Y(n_1436)
);

NAND2xp5_ASAP7_75t_L g1437 ( 
.A(n_1296),
.B(n_1301),
.Y(n_1437)
);

INVx3_ASAP7_75t_L g1438 ( 
.A(n_1314),
.Y(n_1438)
);

AND2x2_ASAP7_75t_L g1439 ( 
.A(n_1277),
.B(n_78),
.Y(n_1439)
);

AND3x1_ASAP7_75t_SL g1440 ( 
.A(n_1256),
.B(n_78),
.C(n_79),
.Y(n_1440)
);

AND2x2_ASAP7_75t_L g1441 ( 
.A(n_1272),
.B(n_79),
.Y(n_1441)
);

NAND2xp5_ASAP7_75t_L g1442 ( 
.A(n_1279),
.B(n_80),
.Y(n_1442)
);

NAND2xp5_ASAP7_75t_L g1443 ( 
.A(n_1372),
.B(n_80),
.Y(n_1443)
);

NAND2xp5_ASAP7_75t_SL g1444 ( 
.A(n_1389),
.B(n_81),
.Y(n_1444)
);

INVx1_ASAP7_75t_L g1445 ( 
.A(n_1260),
.Y(n_1445)
);

BUFx8_ASAP7_75t_L g1446 ( 
.A(n_1304),
.Y(n_1446)
);

INVx3_ASAP7_75t_L g1447 ( 
.A(n_1314),
.Y(n_1447)
);

OAI21xp5_ASAP7_75t_L g1448 ( 
.A1(n_1407),
.A2(n_397),
.B(n_396),
.Y(n_1448)
);

NAND2xp5_ASAP7_75t_L g1449 ( 
.A(n_1282),
.B(n_81),
.Y(n_1449)
);

NOR2x1_ASAP7_75t_L g1450 ( 
.A(n_1302),
.B(n_398),
.Y(n_1450)
);

AND2x2_ASAP7_75t_L g1451 ( 
.A(n_1434),
.B(n_82),
.Y(n_1451)
);

INVx6_ASAP7_75t_L g1452 ( 
.A(n_1274),
.Y(n_1452)
);

CKINVDCx11_ASAP7_75t_R g1453 ( 
.A(n_1269),
.Y(n_1453)
);

BUFx12f_ASAP7_75t_L g1454 ( 
.A(n_1274),
.Y(n_1454)
);

INVx2_ASAP7_75t_L g1455 ( 
.A(n_1262),
.Y(n_1455)
);

INVx1_ASAP7_75t_L g1456 ( 
.A(n_1287),
.Y(n_1456)
);

CKINVDCx20_ASAP7_75t_R g1457 ( 
.A(n_1291),
.Y(n_1457)
);

CKINVDCx11_ASAP7_75t_R g1458 ( 
.A(n_1396),
.Y(n_1458)
);

BUFx2_ASAP7_75t_L g1459 ( 
.A(n_1286),
.Y(n_1459)
);

NAND2xp5_ASAP7_75t_L g1460 ( 
.A(n_1384),
.B(n_83),
.Y(n_1460)
);

NAND2xp5_ASAP7_75t_L g1461 ( 
.A(n_1276),
.B(n_1435),
.Y(n_1461)
);

AND2x2_ASAP7_75t_L g1462 ( 
.A(n_1298),
.B(n_1351),
.Y(n_1462)
);

BUFx2_ASAP7_75t_SL g1463 ( 
.A(n_1369),
.Y(n_1463)
);

NAND2xp5_ASAP7_75t_SL g1464 ( 
.A(n_1379),
.B(n_83),
.Y(n_1464)
);

NAND2xp5_ASAP7_75t_SL g1465 ( 
.A(n_1379),
.B(n_84),
.Y(n_1465)
);

HB1xp67_ASAP7_75t_L g1466 ( 
.A(n_1313),
.Y(n_1466)
);

NAND2xp5_ASAP7_75t_L g1467 ( 
.A(n_1268),
.B(n_86),
.Y(n_1467)
);

AOI22xp33_ASAP7_75t_L g1468 ( 
.A1(n_1374),
.A2(n_89),
.B1(n_86),
.B2(n_87),
.Y(n_1468)
);

INVx1_ASAP7_75t_L g1469 ( 
.A(n_1436),
.Y(n_1469)
);

AND2x2_ASAP7_75t_L g1470 ( 
.A(n_1316),
.B(n_87),
.Y(n_1470)
);

BUFx12f_ASAP7_75t_L g1471 ( 
.A(n_1337),
.Y(n_1471)
);

INVx1_ASAP7_75t_L g1472 ( 
.A(n_1303),
.Y(n_1472)
);

NAND2x1p5_ASAP7_75t_L g1473 ( 
.A(n_1314),
.B(n_401),
.Y(n_1473)
);

AND2x2_ASAP7_75t_L g1474 ( 
.A(n_1327),
.B(n_90),
.Y(n_1474)
);

INVx1_ASAP7_75t_L g1475 ( 
.A(n_1308),
.Y(n_1475)
);

NAND2xp5_ASAP7_75t_L g1476 ( 
.A(n_1255),
.B(n_1306),
.Y(n_1476)
);

INVx3_ASAP7_75t_L g1477 ( 
.A(n_1326),
.Y(n_1477)
);

INVx2_ASAP7_75t_L g1478 ( 
.A(n_1312),
.Y(n_1478)
);

BUFx3_ASAP7_75t_L g1479 ( 
.A(n_1315),
.Y(n_1479)
);

HB1xp67_ASAP7_75t_L g1480 ( 
.A(n_1360),
.Y(n_1480)
);

CKINVDCx5p33_ASAP7_75t_R g1481 ( 
.A(n_1402),
.Y(n_1481)
);

INVx1_ASAP7_75t_L g1482 ( 
.A(n_1336),
.Y(n_1482)
);

CKINVDCx5p33_ASAP7_75t_R g1483 ( 
.A(n_1402),
.Y(n_1483)
);

AND2x4_ASAP7_75t_L g1484 ( 
.A(n_1358),
.B(n_402),
.Y(n_1484)
);

NAND2xp5_ASAP7_75t_SL g1485 ( 
.A(n_1369),
.B(n_91),
.Y(n_1485)
);

AND2x2_ASAP7_75t_L g1486 ( 
.A(n_1373),
.B(n_91),
.Y(n_1486)
);

INVx3_ASAP7_75t_SL g1487 ( 
.A(n_1341),
.Y(n_1487)
);

BUFx3_ASAP7_75t_L g1488 ( 
.A(n_1369),
.Y(n_1488)
);

HB1xp67_ASAP7_75t_L g1489 ( 
.A(n_1392),
.Y(n_1489)
);

AOI22xp5_ASAP7_75t_L g1490 ( 
.A1(n_1405),
.A2(n_94),
.B1(n_92),
.B2(n_93),
.Y(n_1490)
);

NAND2xp5_ASAP7_75t_L g1491 ( 
.A(n_1259),
.B(n_92),
.Y(n_1491)
);

NAND2xp5_ASAP7_75t_SL g1492 ( 
.A(n_1345),
.B(n_93),
.Y(n_1492)
);

INVx1_ASAP7_75t_L g1493 ( 
.A(n_1338),
.Y(n_1493)
);

CKINVDCx5p33_ASAP7_75t_R g1494 ( 
.A(n_1283),
.Y(n_1494)
);

NAND2xp5_ASAP7_75t_L g1495 ( 
.A(n_1358),
.B(n_95),
.Y(n_1495)
);

NAND2xp5_ASAP7_75t_L g1496 ( 
.A(n_1321),
.B(n_95),
.Y(n_1496)
);

NAND2xp5_ASAP7_75t_L g1497 ( 
.A(n_1305),
.B(n_96),
.Y(n_1497)
);

NOR2xp33_ASAP7_75t_R g1498 ( 
.A(n_1326),
.B(n_1330),
.Y(n_1498)
);

AND2x4_ASAP7_75t_L g1499 ( 
.A(n_1281),
.B(n_515),
.Y(n_1499)
);

NAND2xp5_ASAP7_75t_L g1500 ( 
.A(n_1309),
.B(n_96),
.Y(n_1500)
);

AND2x2_ASAP7_75t_L g1501 ( 
.A(n_1346),
.B(n_97),
.Y(n_1501)
);

NAND2xp5_ASAP7_75t_L g1502 ( 
.A(n_1318),
.B(n_97),
.Y(n_1502)
);

AND2x2_ASAP7_75t_L g1503 ( 
.A(n_1385),
.B(n_98),
.Y(n_1503)
);

CKINVDCx5p33_ASAP7_75t_R g1504 ( 
.A(n_1341),
.Y(n_1504)
);

NOR2xp67_ASAP7_75t_SL g1505 ( 
.A(n_1326),
.B(n_98),
.Y(n_1505)
);

AOI22xp33_ASAP7_75t_L g1506 ( 
.A1(n_1413),
.A2(n_101),
.B1(n_99),
.B2(n_100),
.Y(n_1506)
);

INVx1_ASAP7_75t_L g1507 ( 
.A(n_1342),
.Y(n_1507)
);

CKINVDCx5p33_ASAP7_75t_R g1508 ( 
.A(n_1367),
.Y(n_1508)
);

AND2x2_ASAP7_75t_L g1509 ( 
.A(n_1426),
.B(n_99),
.Y(n_1509)
);

INVxp67_ASAP7_75t_L g1510 ( 
.A(n_1377),
.Y(n_1510)
);

INVx1_ASAP7_75t_L g1511 ( 
.A(n_1387),
.Y(n_1511)
);

INVx3_ASAP7_75t_L g1512 ( 
.A(n_1330),
.Y(n_1512)
);

INVx1_ASAP7_75t_L g1513 ( 
.A(n_1388),
.Y(n_1513)
);

A2O1A1Ixp33_ASAP7_75t_L g1514 ( 
.A1(n_1267),
.A2(n_1264),
.B(n_1411),
.C(n_1322),
.Y(n_1514)
);

NAND2xp5_ASAP7_75t_L g1515 ( 
.A(n_1281),
.B(n_101),
.Y(n_1515)
);

INVxp67_ASAP7_75t_SL g1516 ( 
.A(n_1362),
.Y(n_1516)
);

HB1xp67_ASAP7_75t_L g1517 ( 
.A(n_1362),
.Y(n_1517)
);

INVx2_ASAP7_75t_L g1518 ( 
.A(n_1362),
.Y(n_1518)
);

BUFx12f_ASAP7_75t_L g1519 ( 
.A(n_1330),
.Y(n_1519)
);

INVx1_ASAP7_75t_L g1520 ( 
.A(n_1400),
.Y(n_1520)
);

AOI22xp5_ASAP7_75t_L g1521 ( 
.A1(n_1390),
.A2(n_107),
.B1(n_104),
.B2(n_106),
.Y(n_1521)
);

BUFx8_ASAP7_75t_L g1522 ( 
.A(n_1421),
.Y(n_1522)
);

INVx1_ASAP7_75t_L g1523 ( 
.A(n_1348),
.Y(n_1523)
);

CKINVDCx20_ASAP7_75t_R g1524 ( 
.A(n_1418),
.Y(n_1524)
);

INVx1_ASAP7_75t_L g1525 ( 
.A(n_1349),
.Y(n_1525)
);

AND2x2_ASAP7_75t_L g1526 ( 
.A(n_1399),
.B(n_104),
.Y(n_1526)
);

NAND2xp5_ASAP7_75t_SL g1527 ( 
.A(n_1270),
.B(n_106),
.Y(n_1527)
);

CKINVDCx8_ASAP7_75t_R g1528 ( 
.A(n_1391),
.Y(n_1528)
);

CKINVDCx5p33_ASAP7_75t_R g1529 ( 
.A(n_1368),
.Y(n_1529)
);

AND2x2_ASAP7_75t_L g1530 ( 
.A(n_1339),
.B(n_1420),
.Y(n_1530)
);

INVx1_ASAP7_75t_L g1531 ( 
.A(n_1352),
.Y(n_1531)
);

CKINVDCx5p33_ASAP7_75t_R g1532 ( 
.A(n_1261),
.Y(n_1532)
);

INVx1_ASAP7_75t_L g1533 ( 
.A(n_1354),
.Y(n_1533)
);

INVx1_ASAP7_75t_L g1534 ( 
.A(n_1355),
.Y(n_1534)
);

INVx1_ASAP7_75t_L g1535 ( 
.A(n_1359),
.Y(n_1535)
);

BUFx2_ASAP7_75t_L g1536 ( 
.A(n_1334),
.Y(n_1536)
);

NAND2xp5_ASAP7_75t_L g1537 ( 
.A(n_1257),
.B(n_107),
.Y(n_1537)
);

NAND2xp5_ASAP7_75t_L g1538 ( 
.A(n_1328),
.B(n_108),
.Y(n_1538)
);

NAND2xp5_ASAP7_75t_L g1539 ( 
.A(n_1335),
.B(n_109),
.Y(n_1539)
);

AND2x2_ASAP7_75t_L g1540 ( 
.A(n_1416),
.B(n_109),
.Y(n_1540)
);

INVx1_ASAP7_75t_L g1541 ( 
.A(n_1403),
.Y(n_1541)
);

INVx2_ASAP7_75t_L g1542 ( 
.A(n_1376),
.Y(n_1542)
);

AND2x2_ASAP7_75t_SL g1543 ( 
.A(n_1413),
.B(n_110),
.Y(n_1543)
);

OAI22xp5_ASAP7_75t_SL g1544 ( 
.A1(n_1427),
.A2(n_1408),
.B1(n_1370),
.B2(n_1430),
.Y(n_1544)
);

AOI221xp5_ASAP7_75t_L g1545 ( 
.A1(n_1419),
.A2(n_111),
.B1(n_112),
.B2(n_113),
.C(n_114),
.Y(n_1545)
);

CKINVDCx16_ASAP7_75t_R g1546 ( 
.A(n_1356),
.Y(n_1546)
);

NAND2xp5_ASAP7_75t_SL g1547 ( 
.A(n_1430),
.B(n_1285),
.Y(n_1547)
);

CKINVDCx5p33_ASAP7_75t_R g1548 ( 
.A(n_1278),
.Y(n_1548)
);

INVx1_ASAP7_75t_L g1549 ( 
.A(n_1397),
.Y(n_1549)
);

NAND2xp5_ASAP7_75t_L g1550 ( 
.A(n_1409),
.B(n_111),
.Y(n_1550)
);

AOI22xp5_ASAP7_75t_L g1551 ( 
.A1(n_1332),
.A2(n_1347),
.B1(n_1422),
.B2(n_1423),
.Y(n_1551)
);

BUFx6f_ASAP7_75t_L g1552 ( 
.A(n_1299),
.Y(n_1552)
);

NAND2xp5_ASAP7_75t_L g1553 ( 
.A(n_1284),
.B(n_1417),
.Y(n_1553)
);

INVx1_ASAP7_75t_L g1554 ( 
.A(n_1429),
.Y(n_1554)
);

NAND2xp5_ASAP7_75t_L g1555 ( 
.A(n_1343),
.B(n_112),
.Y(n_1555)
);

INVx1_ASAP7_75t_L g1556 ( 
.A(n_1424),
.Y(n_1556)
);

AOI22xp33_ASAP7_75t_L g1557 ( 
.A1(n_1430),
.A2(n_115),
.B1(n_113),
.B2(n_114),
.Y(n_1557)
);

INVx3_ASAP7_75t_L g1558 ( 
.A(n_1376),
.Y(n_1558)
);

OR2x2_ASAP7_75t_L g1559 ( 
.A(n_1280),
.B(n_115),
.Y(n_1559)
);

AO22x1_ASAP7_75t_L g1560 ( 
.A1(n_1433),
.A2(n_119),
.B1(n_116),
.B2(n_118),
.Y(n_1560)
);

INVx1_ASAP7_75t_SL g1561 ( 
.A(n_1428),
.Y(n_1561)
);

AND3x1_ASAP7_75t_SL g1562 ( 
.A(n_1317),
.B(n_116),
.C(n_118),
.Y(n_1562)
);

INVx2_ASAP7_75t_L g1563 ( 
.A(n_1383),
.Y(n_1563)
);

AOI22xp33_ASAP7_75t_L g1564 ( 
.A1(n_1344),
.A2(n_121),
.B1(n_119),
.B2(n_120),
.Y(n_1564)
);

A2O1A1Ixp33_ASAP7_75t_L g1565 ( 
.A1(n_1414),
.A2(n_122),
.B(n_120),
.C(n_121),
.Y(n_1565)
);

NAND2xp5_ASAP7_75t_L g1566 ( 
.A(n_1364),
.B(n_122),
.Y(n_1566)
);

INVx4_ASAP7_75t_L g1567 ( 
.A(n_1383),
.Y(n_1567)
);

NAND2x1_ASAP7_75t_L g1568 ( 
.A(n_1404),
.B(n_404),
.Y(n_1568)
);

AND2x2_ASAP7_75t_L g1569 ( 
.A(n_1432),
.B(n_123),
.Y(n_1569)
);

AND3x1_ASAP7_75t_SL g1570 ( 
.A(n_1425),
.B(n_123),
.C(n_124),
.Y(n_1570)
);

INVx2_ASAP7_75t_L g1571 ( 
.A(n_1357),
.Y(n_1571)
);

NAND2xp5_ASAP7_75t_L g1572 ( 
.A(n_1382),
.B(n_125),
.Y(n_1572)
);

NOR2x1_ASAP7_75t_L g1573 ( 
.A(n_1381),
.B(n_405),
.Y(n_1573)
);

BUFx6f_ASAP7_75t_L g1574 ( 
.A(n_1401),
.Y(n_1574)
);

OAI22xp5_ASAP7_75t_SL g1575 ( 
.A1(n_1406),
.A2(n_1289),
.B1(n_1292),
.B2(n_1398),
.Y(n_1575)
);

OAI22xp5_ASAP7_75t_SL g1576 ( 
.A1(n_1412),
.A2(n_126),
.B1(n_127),
.B2(n_128),
.Y(n_1576)
);

INVx4_ASAP7_75t_L g1577 ( 
.A(n_1401),
.Y(n_1577)
);

INVx1_ASAP7_75t_L g1578 ( 
.A(n_1265),
.Y(n_1578)
);

A2O1A1Ixp33_ASAP7_75t_L g1579 ( 
.A1(n_1375),
.A2(n_126),
.B(n_128),
.C(n_129),
.Y(n_1579)
);

CKINVDCx5p33_ASAP7_75t_R g1580 ( 
.A(n_1293),
.Y(n_1580)
);

AOI22xp5_ASAP7_75t_L g1581 ( 
.A1(n_1340),
.A2(n_129),
.B1(n_130),
.B2(n_131),
.Y(n_1581)
);

NAND2xp5_ASAP7_75t_SL g1582 ( 
.A(n_1275),
.B(n_1350),
.Y(n_1582)
);

NAND2xp5_ASAP7_75t_L g1583 ( 
.A(n_1331),
.B(n_131),
.Y(n_1583)
);

AOI22x1_ASAP7_75t_L g1584 ( 
.A1(n_1431),
.A2(n_412),
.B1(n_513),
.B2(n_511),
.Y(n_1584)
);

INVx1_ASAP7_75t_L g1585 ( 
.A(n_1371),
.Y(n_1585)
);

OAI22xp5_ASAP7_75t_L g1586 ( 
.A1(n_1333),
.A2(n_132),
.B1(n_134),
.B2(n_135),
.Y(n_1586)
);

OAI22xp5_ASAP7_75t_L g1587 ( 
.A1(n_1273),
.A2(n_135),
.B1(n_136),
.B2(n_137),
.Y(n_1587)
);

INVx1_ASAP7_75t_L g1588 ( 
.A(n_1323),
.Y(n_1588)
);

HB1xp67_ASAP7_75t_L g1589 ( 
.A(n_1300),
.Y(n_1589)
);

AND3x1_ASAP7_75t_SL g1590 ( 
.A(n_1366),
.B(n_136),
.C(n_137),
.Y(n_1590)
);

BUFx6f_ASAP7_75t_L g1591 ( 
.A(n_1263),
.Y(n_1591)
);

INVx1_ASAP7_75t_L g1592 ( 
.A(n_1361),
.Y(n_1592)
);

AND2x2_ASAP7_75t_L g1593 ( 
.A(n_1329),
.B(n_138),
.Y(n_1593)
);

AND2x4_ASAP7_75t_L g1594 ( 
.A(n_1386),
.B(n_406),
.Y(n_1594)
);

CKINVDCx20_ASAP7_75t_R g1595 ( 
.A(n_1363),
.Y(n_1595)
);

OAI22xp5_ASAP7_75t_SL g1596 ( 
.A1(n_1325),
.A2(n_1258),
.B1(n_1415),
.B2(n_1410),
.Y(n_1596)
);

AND2x2_ASAP7_75t_L g1597 ( 
.A(n_1290),
.B(n_1310),
.Y(n_1597)
);

NOR2xp67_ASAP7_75t_L g1598 ( 
.A(n_1266),
.B(n_407),
.Y(n_1598)
);

CKINVDCx8_ASAP7_75t_R g1599 ( 
.A(n_1393),
.Y(n_1599)
);

INVx2_ASAP7_75t_L g1600 ( 
.A(n_1365),
.Y(n_1600)
);

INVx1_ASAP7_75t_L g1601 ( 
.A(n_1394),
.Y(n_1601)
);

OAI22xp5_ASAP7_75t_L g1602 ( 
.A1(n_1378),
.A2(n_138),
.B1(n_139),
.B2(n_140),
.Y(n_1602)
);

BUFx8_ASAP7_75t_L g1603 ( 
.A(n_1395),
.Y(n_1603)
);

A2O1A1Ixp33_ASAP7_75t_L g1604 ( 
.A1(n_1294),
.A2(n_1320),
.B(n_1324),
.C(n_1311),
.Y(n_1604)
);

NAND2xp5_ASAP7_75t_L g1605 ( 
.A(n_1271),
.B(n_139),
.Y(n_1605)
);

AND2x2_ASAP7_75t_L g1606 ( 
.A(n_1319),
.B(n_140),
.Y(n_1606)
);

AND2x4_ASAP7_75t_L g1607 ( 
.A(n_1295),
.B(n_514),
.Y(n_1607)
);

NOR2xp33_ASAP7_75t_L g1608 ( 
.A(n_1297),
.B(n_141),
.Y(n_1608)
);

CKINVDCx5p33_ASAP7_75t_R g1609 ( 
.A(n_1453),
.Y(n_1609)
);

INVx2_ASAP7_75t_L g1610 ( 
.A(n_1455),
.Y(n_1610)
);

NAND2xp5_ASAP7_75t_L g1611 ( 
.A(n_1437),
.B(n_1288),
.Y(n_1611)
);

BUFx2_ASAP7_75t_SL g1612 ( 
.A(n_1528),
.Y(n_1612)
);

BUFx2_ASAP7_75t_L g1613 ( 
.A(n_1459),
.Y(n_1613)
);

AOI21xp5_ASAP7_75t_L g1614 ( 
.A1(n_1604),
.A2(n_1582),
.B(n_1461),
.Y(n_1614)
);

AND2x6_ASAP7_75t_L g1615 ( 
.A(n_1573),
.B(n_1353),
.Y(n_1615)
);

NOR2xp33_ASAP7_75t_L g1616 ( 
.A(n_1476),
.B(n_1380),
.Y(n_1616)
);

INVx2_ASAP7_75t_SL g1617 ( 
.A(n_1452),
.Y(n_1617)
);

BUFx8_ASAP7_75t_SL g1618 ( 
.A(n_1454),
.Y(n_1618)
);

NOR2xp33_ASAP7_75t_L g1619 ( 
.A(n_1523),
.B(n_1307),
.Y(n_1619)
);

NAND2xp5_ASAP7_75t_L g1620 ( 
.A(n_1525),
.B(n_1531),
.Y(n_1620)
);

BUFx6f_ASAP7_75t_L g1621 ( 
.A(n_1574),
.Y(n_1621)
);

AOI21xp5_ASAP7_75t_L g1622 ( 
.A1(n_1575),
.A2(n_411),
.B(n_409),
.Y(n_1622)
);

BUFx6f_ASAP7_75t_L g1623 ( 
.A(n_1574),
.Y(n_1623)
);

INVx2_ASAP7_75t_L g1624 ( 
.A(n_1478),
.Y(n_1624)
);

INVx1_ASAP7_75t_L g1625 ( 
.A(n_1445),
.Y(n_1625)
);

NAND2x1p5_ASAP7_75t_L g1626 ( 
.A(n_1577),
.B(n_1488),
.Y(n_1626)
);

CKINVDCx5p33_ASAP7_75t_R g1627 ( 
.A(n_1458),
.Y(n_1627)
);

CKINVDCx5p33_ASAP7_75t_R g1628 ( 
.A(n_1471),
.Y(n_1628)
);

NOR2x1_ASAP7_75t_L g1629 ( 
.A(n_1463),
.B(n_417),
.Y(n_1629)
);

BUFx10_ASAP7_75t_L g1630 ( 
.A(n_1452),
.Y(n_1630)
);

INVx1_ASAP7_75t_SL g1631 ( 
.A(n_1457),
.Y(n_1631)
);

AND2x2_ASAP7_75t_L g1632 ( 
.A(n_1462),
.B(n_1530),
.Y(n_1632)
);

NOR2xp33_ASAP7_75t_SL g1633 ( 
.A(n_1577),
.B(n_418),
.Y(n_1633)
);

NAND2xp5_ASAP7_75t_L g1634 ( 
.A(n_1533),
.B(n_142),
.Y(n_1634)
);

AOI21xp5_ASAP7_75t_L g1635 ( 
.A1(n_1600),
.A2(n_420),
.B(n_419),
.Y(n_1635)
);

AND2x2_ASAP7_75t_L g1636 ( 
.A(n_1501),
.B(n_142),
.Y(n_1636)
);

BUFx3_ASAP7_75t_L g1637 ( 
.A(n_1479),
.Y(n_1637)
);

CKINVDCx20_ASAP7_75t_R g1638 ( 
.A(n_1446),
.Y(n_1638)
);

AOI21xp5_ASAP7_75t_L g1639 ( 
.A1(n_1514),
.A2(n_510),
.B(n_422),
.Y(n_1639)
);

BUFx2_ASAP7_75t_SL g1640 ( 
.A(n_1574),
.Y(n_1640)
);

NOR2xp33_ASAP7_75t_SL g1641 ( 
.A(n_1494),
.B(n_421),
.Y(n_1641)
);

INVx2_ASAP7_75t_L g1642 ( 
.A(n_1456),
.Y(n_1642)
);

CKINVDCx5p33_ASAP7_75t_R g1643 ( 
.A(n_1446),
.Y(n_1643)
);

CKINVDCx11_ASAP7_75t_R g1644 ( 
.A(n_1487),
.Y(n_1644)
);

AOI21xp5_ASAP7_75t_L g1645 ( 
.A1(n_1549),
.A2(n_425),
.B(n_423),
.Y(n_1645)
);

INVx2_ASAP7_75t_L g1646 ( 
.A(n_1469),
.Y(n_1646)
);

AOI21xp5_ASAP7_75t_L g1647 ( 
.A1(n_1596),
.A2(n_427),
.B(n_426),
.Y(n_1647)
);

BUFx6f_ASAP7_75t_L g1648 ( 
.A(n_1519),
.Y(n_1648)
);

INVxp67_ASAP7_75t_L g1649 ( 
.A(n_1489),
.Y(n_1649)
);

BUFx3_ASAP7_75t_L g1650 ( 
.A(n_1480),
.Y(n_1650)
);

AOI21xp5_ASAP7_75t_L g1651 ( 
.A1(n_1596),
.A2(n_430),
.B(n_429),
.Y(n_1651)
);

BUFx3_ASAP7_75t_L g1652 ( 
.A(n_1466),
.Y(n_1652)
);

BUFx3_ASAP7_75t_L g1653 ( 
.A(n_1438),
.Y(n_1653)
);

INVx1_ASAP7_75t_L g1654 ( 
.A(n_1472),
.Y(n_1654)
);

AOI21x1_ASAP7_75t_L g1655 ( 
.A1(n_1578),
.A2(n_1571),
.B(n_1597),
.Y(n_1655)
);

AO31x2_ASAP7_75t_L g1656 ( 
.A1(n_1601),
.A2(n_143),
.A3(n_144),
.B(n_145),
.Y(n_1656)
);

AOI21xp5_ASAP7_75t_L g1657 ( 
.A1(n_1448),
.A2(n_508),
.B(n_432),
.Y(n_1657)
);

NAND2xp5_ASAP7_75t_SL g1658 ( 
.A(n_1546),
.B(n_144),
.Y(n_1658)
);

CKINVDCx20_ASAP7_75t_R g1659 ( 
.A(n_1524),
.Y(n_1659)
);

AND2x4_ASAP7_75t_L g1660 ( 
.A(n_1499),
.B(n_431),
.Y(n_1660)
);

BUFx2_ASAP7_75t_L g1661 ( 
.A(n_1517),
.Y(n_1661)
);

INVx1_ASAP7_75t_L g1662 ( 
.A(n_1475),
.Y(n_1662)
);

NAND2xp5_ASAP7_75t_L g1663 ( 
.A(n_1534),
.B(n_145),
.Y(n_1663)
);

O2A1O1Ixp5_ASAP7_75t_SL g1664 ( 
.A1(n_1602),
.A2(n_146),
.B(n_147),
.C(n_148),
.Y(n_1664)
);

HB1xp67_ASAP7_75t_L g1665 ( 
.A(n_1510),
.Y(n_1665)
);

OR2x2_ASAP7_75t_L g1666 ( 
.A(n_1561),
.B(n_146),
.Y(n_1666)
);

BUFx2_ASAP7_75t_L g1667 ( 
.A(n_1498),
.Y(n_1667)
);

CKINVDCx20_ASAP7_75t_R g1668 ( 
.A(n_1548),
.Y(n_1668)
);

HB1xp67_ASAP7_75t_L g1669 ( 
.A(n_1518),
.Y(n_1669)
);

INVx1_ASAP7_75t_L g1670 ( 
.A(n_1482),
.Y(n_1670)
);

BUFx2_ASAP7_75t_L g1671 ( 
.A(n_1516),
.Y(n_1671)
);

OAI22xp5_ASAP7_75t_L g1672 ( 
.A1(n_1595),
.A2(n_147),
.B1(n_149),
.B2(n_150),
.Y(n_1672)
);

INVx1_ASAP7_75t_L g1673 ( 
.A(n_1493),
.Y(n_1673)
);

AND2x2_ASAP7_75t_L g1674 ( 
.A(n_1451),
.B(n_149),
.Y(n_1674)
);

INVx5_ASAP7_75t_L g1675 ( 
.A(n_1438),
.Y(n_1675)
);

AOI21xp5_ASAP7_75t_L g1676 ( 
.A1(n_1598),
.A2(n_1576),
.B(n_1607),
.Y(n_1676)
);

BUFx6f_ASAP7_75t_L g1677 ( 
.A(n_1552),
.Y(n_1677)
);

BUFx12f_ASAP7_75t_L g1678 ( 
.A(n_1481),
.Y(n_1678)
);

AND2x4_ASAP7_75t_L g1679 ( 
.A(n_1499),
.B(n_433),
.Y(n_1679)
);

OAI22xp5_ASAP7_75t_L g1680 ( 
.A1(n_1580),
.A2(n_152),
.B1(n_154),
.B2(n_155),
.Y(n_1680)
);

INVx4_ASAP7_75t_L g1681 ( 
.A(n_1447),
.Y(n_1681)
);

INVxp67_ASAP7_75t_L g1682 ( 
.A(n_1536),
.Y(n_1682)
);

AOI22xp5_ASAP7_75t_L g1683 ( 
.A1(n_1444),
.A2(n_152),
.B1(n_154),
.B2(n_155),
.Y(n_1683)
);

BUFx3_ASAP7_75t_L g1684 ( 
.A(n_1447),
.Y(n_1684)
);

NAND2xp5_ASAP7_75t_L g1685 ( 
.A(n_1535),
.B(n_156),
.Y(n_1685)
);

AOI21xp5_ASAP7_75t_L g1686 ( 
.A1(n_1598),
.A2(n_437),
.B(n_503),
.Y(n_1686)
);

AOI21xp5_ASAP7_75t_L g1687 ( 
.A1(n_1607),
.A2(n_1553),
.B(n_1513),
.Y(n_1687)
);

INVx3_ASAP7_75t_L g1688 ( 
.A(n_1552),
.Y(n_1688)
);

BUFx3_ASAP7_75t_L g1689 ( 
.A(n_1477),
.Y(n_1689)
);

INVx2_ASAP7_75t_SL g1690 ( 
.A(n_1477),
.Y(n_1690)
);

OAI21xp5_ASAP7_75t_L g1691 ( 
.A1(n_1608),
.A2(n_156),
.B(n_157),
.Y(n_1691)
);

AND2x2_ASAP7_75t_L g1692 ( 
.A(n_1569),
.B(n_157),
.Y(n_1692)
);

BUFx12f_ASAP7_75t_L g1693 ( 
.A(n_1483),
.Y(n_1693)
);

HB1xp67_ASAP7_75t_L g1694 ( 
.A(n_1552),
.Y(n_1694)
);

NAND2xp5_ASAP7_75t_L g1695 ( 
.A(n_1556),
.B(n_158),
.Y(n_1695)
);

INVx2_ASAP7_75t_L g1696 ( 
.A(n_1554),
.Y(n_1696)
);

NAND2x1p5_ASAP7_75t_L g1697 ( 
.A(n_1567),
.B(n_434),
.Y(n_1697)
);

NAND2x1p5_ASAP7_75t_L g1698 ( 
.A(n_1567),
.B(n_438),
.Y(n_1698)
);

AO21x2_ASAP7_75t_L g1699 ( 
.A1(n_1592),
.A2(n_439),
.B(n_502),
.Y(n_1699)
);

AOI21xp5_ASAP7_75t_L g1700 ( 
.A1(n_1511),
.A2(n_505),
.B(n_501),
.Y(n_1700)
);

INVx1_ASAP7_75t_L g1701 ( 
.A(n_1507),
.Y(n_1701)
);

NAND2xp5_ASAP7_75t_L g1702 ( 
.A(n_1520),
.B(n_1541),
.Y(n_1702)
);

OR2x2_ASAP7_75t_L g1703 ( 
.A(n_1538),
.B(n_158),
.Y(n_1703)
);

AND2x2_ASAP7_75t_L g1704 ( 
.A(n_1441),
.B(n_159),
.Y(n_1704)
);

NAND2xp5_ASAP7_75t_L g1705 ( 
.A(n_1442),
.B(n_161),
.Y(n_1705)
);

BUFx2_ASAP7_75t_L g1706 ( 
.A(n_1512),
.Y(n_1706)
);

NOR2xp33_ASAP7_75t_L g1707 ( 
.A(n_1449),
.B(n_440),
.Y(n_1707)
);

CKINVDCx16_ASAP7_75t_R g1708 ( 
.A(n_1470),
.Y(n_1708)
);

BUFx3_ASAP7_75t_L g1709 ( 
.A(n_1512),
.Y(n_1709)
);

AND2x4_ASAP7_75t_L g1710 ( 
.A(n_1558),
.B(n_441),
.Y(n_1710)
);

NAND2xp5_ASAP7_75t_L g1711 ( 
.A(n_1551),
.B(n_161),
.Y(n_1711)
);

NAND2xp5_ASAP7_75t_L g1712 ( 
.A(n_1551),
.B(n_162),
.Y(n_1712)
);

INVx1_ASAP7_75t_SL g1713 ( 
.A(n_1504),
.Y(n_1713)
);

BUFx3_ASAP7_75t_L g1714 ( 
.A(n_1522),
.Y(n_1714)
);

NOR2xp33_ASAP7_75t_L g1715 ( 
.A(n_1491),
.B(n_444),
.Y(n_1715)
);

INVx1_ASAP7_75t_SL g1716 ( 
.A(n_1486),
.Y(n_1716)
);

BUFx3_ASAP7_75t_L g1717 ( 
.A(n_1522),
.Y(n_1717)
);

OAI22xp33_ASAP7_75t_L g1718 ( 
.A1(n_1490),
.A2(n_1521),
.B1(n_1581),
.B2(n_1492),
.Y(n_1718)
);

INVx2_ASAP7_75t_SL g1719 ( 
.A(n_1542),
.Y(n_1719)
);

INVx3_ASAP7_75t_L g1720 ( 
.A(n_1558),
.Y(n_1720)
);

BUFx6f_ASAP7_75t_L g1721 ( 
.A(n_1484),
.Y(n_1721)
);

AND2x2_ASAP7_75t_SL g1722 ( 
.A(n_1543),
.B(n_162),
.Y(n_1722)
);

BUFx6f_ASAP7_75t_L g1723 ( 
.A(n_1484),
.Y(n_1723)
);

NAND3xp33_ASAP7_75t_L g1724 ( 
.A(n_1490),
.B(n_1468),
.C(n_1579),
.Y(n_1724)
);

AOI21xp5_ASAP7_75t_L g1725 ( 
.A1(n_1594),
.A2(n_1605),
.B(n_1547),
.Y(n_1725)
);

AND2x4_ASAP7_75t_L g1726 ( 
.A(n_1563),
.B(n_1515),
.Y(n_1726)
);

HB1xp67_ASAP7_75t_L g1727 ( 
.A(n_1460),
.Y(n_1727)
);

AOI22xp33_ASAP7_75t_SL g1728 ( 
.A1(n_1544),
.A2(n_163),
.B1(n_164),
.B2(n_165),
.Y(n_1728)
);

INVx3_ASAP7_75t_L g1729 ( 
.A(n_1603),
.Y(n_1729)
);

AND2x4_ASAP7_75t_L g1730 ( 
.A(n_1495),
.B(n_446),
.Y(n_1730)
);

INVx1_ASAP7_75t_L g1731 ( 
.A(n_1572),
.Y(n_1731)
);

INVx1_ASAP7_75t_L g1732 ( 
.A(n_1496),
.Y(n_1732)
);

INVx1_ASAP7_75t_SL g1733 ( 
.A(n_1509),
.Y(n_1733)
);

INVx3_ASAP7_75t_L g1734 ( 
.A(n_1603),
.Y(n_1734)
);

OR2x6_ASAP7_75t_SL g1735 ( 
.A(n_1532),
.B(n_165),
.Y(n_1735)
);

A2O1A1Ixp33_ASAP7_75t_L g1736 ( 
.A1(n_1467),
.A2(n_166),
.B(n_167),
.C(n_168),
.Y(n_1736)
);

AOI21xp5_ASAP7_75t_L g1737 ( 
.A1(n_1594),
.A2(n_447),
.B(n_498),
.Y(n_1737)
);

OAI21x1_ASAP7_75t_SL g1738 ( 
.A1(n_1583),
.A2(n_1550),
.B(n_1566),
.Y(n_1738)
);

INVx2_ASAP7_75t_L g1739 ( 
.A(n_1588),
.Y(n_1739)
);

HB1xp67_ASAP7_75t_L g1740 ( 
.A(n_1443),
.Y(n_1740)
);

OR2x2_ASAP7_75t_L g1741 ( 
.A(n_1497),
.B(n_166),
.Y(n_1741)
);

INVx1_ASAP7_75t_L g1742 ( 
.A(n_1500),
.Y(n_1742)
);

INVx1_ASAP7_75t_L g1743 ( 
.A(n_1502),
.Y(n_1743)
);

OAI22xp5_ASAP7_75t_L g1744 ( 
.A1(n_1529),
.A2(n_168),
.B1(n_169),
.B2(n_170),
.Y(n_1744)
);

AND2x4_ASAP7_75t_L g1745 ( 
.A(n_1573),
.B(n_448),
.Y(n_1745)
);

BUFx4f_ASAP7_75t_L g1746 ( 
.A(n_1473),
.Y(n_1746)
);

INVx1_ASAP7_75t_L g1747 ( 
.A(n_1555),
.Y(n_1747)
);

OAI22xp5_ASAP7_75t_L g1748 ( 
.A1(n_1521),
.A2(n_1589),
.B1(n_1599),
.B2(n_1581),
.Y(n_1748)
);

INVx1_ASAP7_75t_L g1749 ( 
.A(n_1537),
.Y(n_1749)
);

BUFx2_ASAP7_75t_L g1750 ( 
.A(n_1508),
.Y(n_1750)
);

BUFx3_ASAP7_75t_L g1751 ( 
.A(n_1439),
.Y(n_1751)
);

AOI21xp5_ASAP7_75t_L g1752 ( 
.A1(n_1585),
.A2(n_500),
.B(n_497),
.Y(n_1752)
);

NAND2xp5_ASAP7_75t_L g1753 ( 
.A(n_1540),
.B(n_169),
.Y(n_1753)
);

O2A1O1Ixp5_ASAP7_75t_L g1754 ( 
.A1(n_1647),
.A2(n_1565),
.B(n_1586),
.C(n_1560),
.Y(n_1754)
);

INVx1_ASAP7_75t_L g1755 ( 
.A(n_1696),
.Y(n_1755)
);

INVx3_ASAP7_75t_SL g1756 ( 
.A(n_1643),
.Y(n_1756)
);

INVx2_ASAP7_75t_L g1757 ( 
.A(n_1610),
.Y(n_1757)
);

INVx1_ASAP7_75t_L g1758 ( 
.A(n_1701),
.Y(n_1758)
);

AND2x4_ASAP7_75t_L g1759 ( 
.A(n_1671),
.B(n_1526),
.Y(n_1759)
);

INVxp67_ASAP7_75t_L g1760 ( 
.A(n_1665),
.Y(n_1760)
);

INVx2_ASAP7_75t_L g1761 ( 
.A(n_1624),
.Y(n_1761)
);

INVx2_ASAP7_75t_L g1762 ( 
.A(n_1642),
.Y(n_1762)
);

A2O1A1Ixp33_ASAP7_75t_L g1763 ( 
.A1(n_1676),
.A2(n_1539),
.B(n_1545),
.C(n_1564),
.Y(n_1763)
);

NAND2x1p5_ASAP7_75t_L g1764 ( 
.A(n_1675),
.B(n_1505),
.Y(n_1764)
);

O2A1O1Ixp33_ASAP7_75t_L g1765 ( 
.A1(n_1691),
.A2(n_1465),
.B(n_1464),
.C(n_1527),
.Y(n_1765)
);

NAND2xp5_ASAP7_75t_L g1766 ( 
.A(n_1731),
.B(n_1593),
.Y(n_1766)
);

AND2x2_ASAP7_75t_L g1767 ( 
.A(n_1632),
.B(n_1474),
.Y(n_1767)
);

NAND2x1p5_ASAP7_75t_L g1768 ( 
.A(n_1675),
.B(n_1729),
.Y(n_1768)
);

INVx1_ASAP7_75t_L g1769 ( 
.A(n_1625),
.Y(n_1769)
);

OAI211xp5_ASAP7_75t_L g1770 ( 
.A1(n_1728),
.A2(n_1506),
.B(n_1557),
.C(n_1559),
.Y(n_1770)
);

O2A1O1Ixp5_ASAP7_75t_L g1771 ( 
.A1(n_1651),
.A2(n_1587),
.B(n_1485),
.C(n_1606),
.Y(n_1771)
);

OR2x6_ASAP7_75t_SL g1772 ( 
.A(n_1609),
.B(n_1570),
.Y(n_1772)
);

OAI22xp5_ASAP7_75t_L g1773 ( 
.A1(n_1718),
.A2(n_1503),
.B1(n_1562),
.B2(n_1584),
.Y(n_1773)
);

AND2x4_ASAP7_75t_L g1774 ( 
.A(n_1734),
.B(n_1450),
.Y(n_1774)
);

HB1xp67_ASAP7_75t_L g1775 ( 
.A(n_1613),
.Y(n_1775)
);

AOI21xp5_ASAP7_75t_L g1776 ( 
.A1(n_1614),
.A2(n_1450),
.B(n_1568),
.Y(n_1776)
);

BUFx4f_ASAP7_75t_SL g1777 ( 
.A(n_1678),
.Y(n_1777)
);

OAI22xp5_ASAP7_75t_L g1778 ( 
.A1(n_1724),
.A2(n_1590),
.B1(n_1440),
.B2(n_1591),
.Y(n_1778)
);

NAND2xp5_ASAP7_75t_L g1779 ( 
.A(n_1687),
.B(n_1591),
.Y(n_1779)
);

INVx2_ASAP7_75t_L g1780 ( 
.A(n_1646),
.Y(n_1780)
);

A2O1A1Ixp33_ASAP7_75t_SL g1781 ( 
.A1(n_1616),
.A2(n_170),
.B(n_171),
.C(n_172),
.Y(n_1781)
);

AND2x4_ASAP7_75t_L g1782 ( 
.A(n_1721),
.B(n_449),
.Y(n_1782)
);

AND2x2_ASAP7_75t_L g1783 ( 
.A(n_1716),
.B(n_450),
.Y(n_1783)
);

OR2x6_ASAP7_75t_L g1784 ( 
.A(n_1725),
.B(n_451),
.Y(n_1784)
);

AND2x2_ASAP7_75t_L g1785 ( 
.A(n_1733),
.B(n_452),
.Y(n_1785)
);

AND2x4_ASAP7_75t_L g1786 ( 
.A(n_1721),
.B(n_454),
.Y(n_1786)
);

NAND2xp5_ASAP7_75t_L g1787 ( 
.A(n_1620),
.B(n_171),
.Y(n_1787)
);

INVxp33_ASAP7_75t_L g1788 ( 
.A(n_1694),
.Y(n_1788)
);

OAI22xp5_ASAP7_75t_SL g1789 ( 
.A1(n_1722),
.A2(n_172),
.B1(n_173),
.B2(n_174),
.Y(n_1789)
);

AOI21xp5_ASAP7_75t_L g1790 ( 
.A1(n_1611),
.A2(n_494),
.B(n_492),
.Y(n_1790)
);

INVx1_ASAP7_75t_L g1791 ( 
.A(n_1654),
.Y(n_1791)
);

OAI22xp5_ASAP7_75t_L g1792 ( 
.A1(n_1748),
.A2(n_175),
.B1(n_176),
.B2(n_177),
.Y(n_1792)
);

AND2x2_ASAP7_75t_L g1793 ( 
.A(n_1692),
.B(n_456),
.Y(n_1793)
);

OAI22xp5_ASAP7_75t_L g1794 ( 
.A1(n_1683),
.A2(n_175),
.B1(n_176),
.B2(n_177),
.Y(n_1794)
);

INVx1_ASAP7_75t_L g1795 ( 
.A(n_1662),
.Y(n_1795)
);

NAND2xp5_ASAP7_75t_L g1796 ( 
.A(n_1702),
.B(n_178),
.Y(n_1796)
);

INVx1_ASAP7_75t_L g1797 ( 
.A(n_1670),
.Y(n_1797)
);

O2A1O1Ixp33_ASAP7_75t_L g1798 ( 
.A1(n_1736),
.A2(n_1658),
.B(n_1712),
.C(n_1711),
.Y(n_1798)
);

A2O1A1Ixp33_ASAP7_75t_L g1799 ( 
.A1(n_1622),
.A2(n_1657),
.B(n_1715),
.C(n_1707),
.Y(n_1799)
);

AND2x2_ASAP7_75t_L g1800 ( 
.A(n_1636),
.B(n_457),
.Y(n_1800)
);

AND2x4_ASAP7_75t_L g1801 ( 
.A(n_1721),
.B(n_458),
.Y(n_1801)
);

AND2x4_ASAP7_75t_L g1802 ( 
.A(n_1723),
.B(n_459),
.Y(n_1802)
);

AND2x2_ASAP7_75t_L g1803 ( 
.A(n_1669),
.B(n_461),
.Y(n_1803)
);

NAND2xp5_ASAP7_75t_L g1804 ( 
.A(n_1749),
.B(n_1732),
.Y(n_1804)
);

AND2x2_ASAP7_75t_L g1805 ( 
.A(n_1674),
.B(n_463),
.Y(n_1805)
);

BUFx2_ASAP7_75t_L g1806 ( 
.A(n_1650),
.Y(n_1806)
);

INVx2_ASAP7_75t_L g1807 ( 
.A(n_1673),
.Y(n_1807)
);

HB1xp67_ASAP7_75t_L g1808 ( 
.A(n_1661),
.Y(n_1808)
);

NAND2x1p5_ASAP7_75t_L g1809 ( 
.A(n_1675),
.B(n_464),
.Y(n_1809)
);

AND2x2_ASAP7_75t_L g1810 ( 
.A(n_1726),
.B(n_465),
.Y(n_1810)
);

AND2x4_ASAP7_75t_L g1811 ( 
.A(n_1723),
.B(n_466),
.Y(n_1811)
);

BUFx3_ASAP7_75t_L g1812 ( 
.A(n_1637),
.Y(n_1812)
);

BUFx6f_ASAP7_75t_L g1813 ( 
.A(n_1621),
.Y(n_1813)
);

INVxp67_ASAP7_75t_SL g1814 ( 
.A(n_1649),
.Y(n_1814)
);

CKINVDCx5p33_ASAP7_75t_R g1815 ( 
.A(n_1618),
.Y(n_1815)
);

OR2x2_ASAP7_75t_L g1816 ( 
.A(n_1740),
.B(n_179),
.Y(n_1816)
);

AND2x2_ASAP7_75t_L g1817 ( 
.A(n_1726),
.B(n_468),
.Y(n_1817)
);

NAND2xp5_ASAP7_75t_L g1818 ( 
.A(n_1742),
.B(n_181),
.Y(n_1818)
);

HB1xp67_ASAP7_75t_L g1819 ( 
.A(n_1652),
.Y(n_1819)
);

HB1xp67_ASAP7_75t_L g1820 ( 
.A(n_1682),
.Y(n_1820)
);

AND2x4_ASAP7_75t_L g1821 ( 
.A(n_1723),
.B(n_469),
.Y(n_1821)
);

AND2x2_ASAP7_75t_L g1822 ( 
.A(n_1704),
.B(n_490),
.Y(n_1822)
);

INVx2_ASAP7_75t_L g1823 ( 
.A(n_1719),
.Y(n_1823)
);

NAND2xp5_ASAP7_75t_L g1824 ( 
.A(n_1743),
.B(n_182),
.Y(n_1824)
);

AND2x2_ASAP7_75t_L g1825 ( 
.A(n_1727),
.B(n_489),
.Y(n_1825)
);

A2O1A1Ixp33_ASAP7_75t_SL g1826 ( 
.A1(n_1619),
.A2(n_183),
.B(n_184),
.C(n_185),
.Y(n_1826)
);

BUFx2_ASAP7_75t_L g1827 ( 
.A(n_1677),
.Y(n_1827)
);

A2O1A1Ixp33_ASAP7_75t_L g1828 ( 
.A1(n_1639),
.A2(n_183),
.B(n_184),
.C(n_185),
.Y(n_1828)
);

AND2x2_ASAP7_75t_L g1829 ( 
.A(n_1751),
.B(n_488),
.Y(n_1829)
);

NOR2x2_ASAP7_75t_L g1830 ( 
.A(n_1739),
.B(n_186),
.Y(n_1830)
);

OR2x2_ASAP7_75t_L g1831 ( 
.A(n_1747),
.B(n_186),
.Y(n_1831)
);

AND2x2_ASAP7_75t_L g1832 ( 
.A(n_1708),
.B(n_486),
.Y(n_1832)
);

CKINVDCx14_ASAP7_75t_R g1833 ( 
.A(n_1627),
.Y(n_1833)
);

INVx3_ASAP7_75t_L g1834 ( 
.A(n_1681),
.Y(n_1834)
);

INVx1_ASAP7_75t_L g1835 ( 
.A(n_1656),
.Y(n_1835)
);

HB1xp67_ASAP7_75t_L g1836 ( 
.A(n_1706),
.Y(n_1836)
);

INVx2_ASAP7_75t_L g1837 ( 
.A(n_1720),
.Y(n_1837)
);

NAND2xp5_ASAP7_75t_L g1838 ( 
.A(n_1738),
.B(n_187),
.Y(n_1838)
);

OR2x2_ASAP7_75t_SL g1839 ( 
.A(n_1703),
.B(n_188),
.Y(n_1839)
);

OR2x2_ASAP7_75t_L g1840 ( 
.A(n_1741),
.B(n_190),
.Y(n_1840)
);

AND2x2_ASAP7_75t_L g1841 ( 
.A(n_1753),
.B(n_485),
.Y(n_1841)
);

OA21x2_ASAP7_75t_L g1842 ( 
.A1(n_1655),
.A2(n_190),
.B(n_191),
.Y(n_1842)
);

AND2x2_ASAP7_75t_L g1843 ( 
.A(n_1688),
.B(n_484),
.Y(n_1843)
);

INVx2_ASAP7_75t_L g1844 ( 
.A(n_1690),
.Y(n_1844)
);

AND2x2_ASAP7_75t_L g1845 ( 
.A(n_1705),
.B(n_482),
.Y(n_1845)
);

HB1xp67_ASAP7_75t_L g1846 ( 
.A(n_1677),
.Y(n_1846)
);

CKINVDCx20_ASAP7_75t_R g1847 ( 
.A(n_1638),
.Y(n_1847)
);

OAI22xp33_ASAP7_75t_L g1848 ( 
.A1(n_1773),
.A2(n_1735),
.B1(n_1633),
.B2(n_1672),
.Y(n_1848)
);

OAI21xp5_ASAP7_75t_L g1849 ( 
.A1(n_1799),
.A2(n_1737),
.B(n_1700),
.Y(n_1849)
);

INVx2_ASAP7_75t_L g1850 ( 
.A(n_1762),
.Y(n_1850)
);

INVx1_ASAP7_75t_L g1851 ( 
.A(n_1758),
.Y(n_1851)
);

INVx3_ASAP7_75t_L g1852 ( 
.A(n_1780),
.Y(n_1852)
);

BUFx6f_ASAP7_75t_L g1853 ( 
.A(n_1812),
.Y(n_1853)
);

AOI22xp33_ASAP7_75t_L g1854 ( 
.A1(n_1789),
.A2(n_1680),
.B1(n_1730),
.B2(n_1744),
.Y(n_1854)
);

INVx4_ASAP7_75t_L g1855 ( 
.A(n_1834),
.Y(n_1855)
);

OR2x2_ASAP7_75t_SL g1856 ( 
.A(n_1838),
.B(n_1819),
.Y(n_1856)
);

OAI22xp5_ASAP7_75t_L g1857 ( 
.A1(n_1789),
.A2(n_1746),
.B1(n_1659),
.B2(n_1667),
.Y(n_1857)
);

INVx1_ASAP7_75t_L g1858 ( 
.A(n_1769),
.Y(n_1858)
);

BUFx3_ASAP7_75t_L g1859 ( 
.A(n_1806),
.Y(n_1859)
);

INVx2_ASAP7_75t_L g1860 ( 
.A(n_1807),
.Y(n_1860)
);

OAI22xp33_ASAP7_75t_L g1861 ( 
.A1(n_1773),
.A2(n_1641),
.B1(n_1695),
.B2(n_1663),
.Y(n_1861)
);

AOI22xp33_ASAP7_75t_L g1862 ( 
.A1(n_1794),
.A2(n_1730),
.B1(n_1745),
.B2(n_1615),
.Y(n_1862)
);

NAND3xp33_ASAP7_75t_L g1863 ( 
.A(n_1828),
.B(n_1664),
.C(n_1634),
.Y(n_1863)
);

AOI21xp5_ASAP7_75t_L g1864 ( 
.A1(n_1776),
.A2(n_1635),
.B(n_1686),
.Y(n_1864)
);

INVx3_ASAP7_75t_SL g1865 ( 
.A(n_1815),
.Y(n_1865)
);

CKINVDCx5p33_ASAP7_75t_R g1866 ( 
.A(n_1847),
.Y(n_1866)
);

AND2x4_ASAP7_75t_L g1867 ( 
.A(n_1791),
.B(n_1677),
.Y(n_1867)
);

BUFx2_ASAP7_75t_L g1868 ( 
.A(n_1775),
.Y(n_1868)
);

NAND2xp5_ASAP7_75t_L g1869 ( 
.A(n_1766),
.B(n_1685),
.Y(n_1869)
);

AOI22xp5_ASAP7_75t_L g1870 ( 
.A1(n_1770),
.A2(n_1794),
.B1(n_1792),
.B2(n_1778),
.Y(n_1870)
);

INVx1_ASAP7_75t_L g1871 ( 
.A(n_1795),
.Y(n_1871)
);

INVx1_ASAP7_75t_L g1872 ( 
.A(n_1797),
.Y(n_1872)
);

AOI22xp33_ASAP7_75t_L g1873 ( 
.A1(n_1792),
.A2(n_1745),
.B1(n_1615),
.B2(n_1750),
.Y(n_1873)
);

BUFx3_ASAP7_75t_L g1874 ( 
.A(n_1827),
.Y(n_1874)
);

OAI22xp5_ASAP7_75t_L g1875 ( 
.A1(n_1772),
.A2(n_1660),
.B1(n_1679),
.B2(n_1668),
.Y(n_1875)
);

OAI21xp5_ASAP7_75t_SL g1876 ( 
.A1(n_1765),
.A2(n_1679),
.B(n_1629),
.Y(n_1876)
);

INVx2_ASAP7_75t_L g1877 ( 
.A(n_1755),
.Y(n_1877)
);

AOI22xp33_ASAP7_75t_L g1878 ( 
.A1(n_1778),
.A2(n_1615),
.B1(n_1717),
.B2(n_1714),
.Y(n_1878)
);

AOI22xp33_ASAP7_75t_SL g1879 ( 
.A1(n_1784),
.A2(n_1838),
.B1(n_1615),
.B2(n_1766),
.Y(n_1879)
);

AOI22xp33_ASAP7_75t_L g1880 ( 
.A1(n_1784),
.A2(n_1644),
.B1(n_1666),
.B2(n_1631),
.Y(n_1880)
);

INVx1_ASAP7_75t_SL g1881 ( 
.A(n_1767),
.Y(n_1881)
);

OAI22xp5_ASAP7_75t_L g1882 ( 
.A1(n_1763),
.A2(n_1612),
.B1(n_1626),
.B2(n_1713),
.Y(n_1882)
);

BUFx6f_ASAP7_75t_SL g1883 ( 
.A(n_1782),
.Y(n_1883)
);

AOI22xp33_ASAP7_75t_L g1884 ( 
.A1(n_1784),
.A2(n_1645),
.B1(n_1699),
.B2(n_1710),
.Y(n_1884)
);

INVx1_ASAP7_75t_SL g1885 ( 
.A(n_1808),
.Y(n_1885)
);

AOI22xp33_ASAP7_75t_SL g1886 ( 
.A1(n_1774),
.A2(n_1752),
.B1(n_1698),
.B2(n_1697),
.Y(n_1886)
);

CKINVDCx5p33_ASAP7_75t_R g1887 ( 
.A(n_1833),
.Y(n_1887)
);

HB1xp67_ASAP7_75t_L g1888 ( 
.A(n_1836),
.Y(n_1888)
);

INVx1_ASAP7_75t_L g1889 ( 
.A(n_1835),
.Y(n_1889)
);

AOI22xp33_ASAP7_75t_L g1890 ( 
.A1(n_1845),
.A2(n_1710),
.B1(n_1617),
.B2(n_1648),
.Y(n_1890)
);

BUFx5_ASAP7_75t_L g1891 ( 
.A(n_1774),
.Y(n_1891)
);

AOI22xp5_ASAP7_75t_L g1892 ( 
.A1(n_1759),
.A2(n_1640),
.B1(n_1648),
.B2(n_1621),
.Y(n_1892)
);

AOI22xp5_ASAP7_75t_L g1893 ( 
.A1(n_1759),
.A2(n_1648),
.B1(n_1623),
.B2(n_1621),
.Y(n_1893)
);

BUFx2_ASAP7_75t_L g1894 ( 
.A(n_1846),
.Y(n_1894)
);

CKINVDCx5p33_ASAP7_75t_R g1895 ( 
.A(n_1756),
.Y(n_1895)
);

INVx3_ASAP7_75t_L g1896 ( 
.A(n_1834),
.Y(n_1896)
);

AOI22xp33_ASAP7_75t_L g1897 ( 
.A1(n_1841),
.A2(n_1630),
.B1(n_1693),
.B2(n_1689),
.Y(n_1897)
);

OAI21xp33_ASAP7_75t_L g1898 ( 
.A1(n_1798),
.A2(n_1709),
.B(n_1684),
.Y(n_1898)
);

INVx2_ASAP7_75t_L g1899 ( 
.A(n_1757),
.Y(n_1899)
);

INVx3_ASAP7_75t_L g1900 ( 
.A(n_1768),
.Y(n_1900)
);

AOI22xp33_ASAP7_75t_L g1901 ( 
.A1(n_1832),
.A2(n_1630),
.B1(n_1653),
.B2(n_1623),
.Y(n_1901)
);

OAI22xp5_ASAP7_75t_L g1902 ( 
.A1(n_1839),
.A2(n_1623),
.B1(n_1681),
.B2(n_1628),
.Y(n_1902)
);

INVx1_ASAP7_75t_L g1903 ( 
.A(n_1851),
.Y(n_1903)
);

AND2x2_ASAP7_75t_L g1904 ( 
.A(n_1858),
.B(n_1842),
.Y(n_1904)
);

AND2x2_ASAP7_75t_L g1905 ( 
.A(n_1871),
.B(n_1842),
.Y(n_1905)
);

BUFx3_ASAP7_75t_L g1906 ( 
.A(n_1853),
.Y(n_1906)
);

NAND2xp33_ASAP7_75t_L g1907 ( 
.A(n_1870),
.B(n_1764),
.Y(n_1907)
);

AOI221x1_ASAP7_75t_SL g1908 ( 
.A1(n_1848),
.A2(n_1804),
.B1(n_1818),
.B2(n_1824),
.C(n_1796),
.Y(n_1908)
);

AO21x2_ASAP7_75t_L g1909 ( 
.A1(n_1849),
.A2(n_1779),
.B(n_1826),
.Y(n_1909)
);

A2O1A1Ixp33_ASAP7_75t_L g1910 ( 
.A1(n_1870),
.A2(n_1754),
.B(n_1771),
.C(n_1781),
.Y(n_1910)
);

AOI22xp33_ASAP7_75t_L g1911 ( 
.A1(n_1861),
.A2(n_1790),
.B1(n_1817),
.B2(n_1810),
.Y(n_1911)
);

INVx2_ASAP7_75t_L g1912 ( 
.A(n_1877),
.Y(n_1912)
);

AND2x2_ASAP7_75t_L g1913 ( 
.A(n_1872),
.B(n_1779),
.Y(n_1913)
);

CKINVDCx5p33_ASAP7_75t_R g1914 ( 
.A(n_1866),
.Y(n_1914)
);

OR2x2_ASAP7_75t_L g1915 ( 
.A(n_1856),
.B(n_1814),
.Y(n_1915)
);

OR2x2_ASAP7_75t_L g1916 ( 
.A(n_1888),
.B(n_1868),
.Y(n_1916)
);

INVx2_ASAP7_75t_L g1917 ( 
.A(n_1860),
.Y(n_1917)
);

INVx2_ASAP7_75t_L g1918 ( 
.A(n_1889),
.Y(n_1918)
);

NOR2x1_ASAP7_75t_SL g1919 ( 
.A(n_1876),
.B(n_1855),
.Y(n_1919)
);

AND2x2_ASAP7_75t_L g1920 ( 
.A(n_1891),
.B(n_1656),
.Y(n_1920)
);

INVx1_ASAP7_75t_L g1921 ( 
.A(n_1850),
.Y(n_1921)
);

CKINVDCx5p33_ASAP7_75t_R g1922 ( 
.A(n_1887),
.Y(n_1922)
);

BUFx4f_ASAP7_75t_SL g1923 ( 
.A(n_1865),
.Y(n_1923)
);

AO32x2_ASAP7_75t_L g1924 ( 
.A1(n_1902),
.A2(n_1830),
.A3(n_1760),
.B1(n_1656),
.B2(n_1820),
.Y(n_1924)
);

NAND2x1p5_ASAP7_75t_L g1925 ( 
.A(n_1855),
.B(n_1896),
.Y(n_1925)
);

INVx1_ASAP7_75t_L g1926 ( 
.A(n_1899),
.Y(n_1926)
);

HB1xp67_ASAP7_75t_L g1927 ( 
.A(n_1885),
.Y(n_1927)
);

OR2x2_ASAP7_75t_L g1928 ( 
.A(n_1881),
.B(n_1816),
.Y(n_1928)
);

AND2x2_ASAP7_75t_L g1929 ( 
.A(n_1891),
.B(n_1761),
.Y(n_1929)
);

OR2x2_ASAP7_75t_L g1930 ( 
.A(n_1894),
.B(n_1831),
.Y(n_1930)
);

AOI22xp33_ASAP7_75t_L g1931 ( 
.A1(n_1879),
.A2(n_1793),
.B1(n_1805),
.B2(n_1822),
.Y(n_1931)
);

CKINVDCx5p33_ASAP7_75t_R g1932 ( 
.A(n_1895),
.Y(n_1932)
);

INVx5_ASAP7_75t_SL g1933 ( 
.A(n_1853),
.Y(n_1933)
);

INVx2_ASAP7_75t_L g1934 ( 
.A(n_1918),
.Y(n_1934)
);

AOI22xp33_ASAP7_75t_SL g1935 ( 
.A1(n_1907),
.A2(n_1882),
.B1(n_1883),
.B2(n_1863),
.Y(n_1935)
);

AND2x2_ASAP7_75t_L g1936 ( 
.A(n_1916),
.B(n_1920),
.Y(n_1936)
);

INVx1_ASAP7_75t_L g1937 ( 
.A(n_1918),
.Y(n_1937)
);

INVx2_ASAP7_75t_L g1938 ( 
.A(n_1912),
.Y(n_1938)
);

INVx1_ASAP7_75t_L g1939 ( 
.A(n_1903),
.Y(n_1939)
);

AND2x4_ASAP7_75t_L g1940 ( 
.A(n_1929),
.B(n_1867),
.Y(n_1940)
);

NAND2xp5_ASAP7_75t_L g1941 ( 
.A(n_1913),
.B(n_1869),
.Y(n_1941)
);

HB1xp67_ASAP7_75t_L g1942 ( 
.A(n_1927),
.Y(n_1942)
);

AND2x2_ASAP7_75t_L g1943 ( 
.A(n_1916),
.B(n_1859),
.Y(n_1943)
);

HB1xp67_ASAP7_75t_L g1944 ( 
.A(n_1915),
.Y(n_1944)
);

INVx2_ASAP7_75t_L g1945 ( 
.A(n_1912),
.Y(n_1945)
);

INVx1_ASAP7_75t_L g1946 ( 
.A(n_1917),
.Y(n_1946)
);

INVx2_ASAP7_75t_L g1947 ( 
.A(n_1917),
.Y(n_1947)
);

AND2x2_ASAP7_75t_L g1948 ( 
.A(n_1920),
.B(n_1891),
.Y(n_1948)
);

NOR2xp67_ASAP7_75t_L g1949 ( 
.A(n_1915),
.B(n_1853),
.Y(n_1949)
);

AND2x2_ASAP7_75t_L g1950 ( 
.A(n_1913),
.B(n_1929),
.Y(n_1950)
);

INVx1_ASAP7_75t_L g1951 ( 
.A(n_1904),
.Y(n_1951)
);

INVx1_ASAP7_75t_L g1952 ( 
.A(n_1921),
.Y(n_1952)
);

OR2x2_ASAP7_75t_L g1953 ( 
.A(n_1930),
.B(n_1852),
.Y(n_1953)
);

AND2x2_ASAP7_75t_L g1954 ( 
.A(n_1904),
.B(n_1891),
.Y(n_1954)
);

INVx1_ASAP7_75t_L g1955 ( 
.A(n_1905),
.Y(n_1955)
);

A2O1A1Ixp33_ASAP7_75t_L g1956 ( 
.A1(n_1935),
.A2(n_1908),
.B(n_1910),
.C(n_1907),
.Y(n_1956)
);

INVx1_ASAP7_75t_L g1957 ( 
.A(n_1939),
.Y(n_1957)
);

AND2x2_ASAP7_75t_L g1958 ( 
.A(n_1936),
.B(n_1906),
.Y(n_1958)
);

INVx1_ASAP7_75t_L g1959 ( 
.A(n_1939),
.Y(n_1959)
);

INVx2_ASAP7_75t_L g1960 ( 
.A(n_1934),
.Y(n_1960)
);

AOI21xp5_ASAP7_75t_L g1961 ( 
.A1(n_1949),
.A2(n_1919),
.B(n_1864),
.Y(n_1961)
);

INVx1_ASAP7_75t_L g1962 ( 
.A(n_1937),
.Y(n_1962)
);

AOI21xp5_ASAP7_75t_L g1963 ( 
.A1(n_1941),
.A2(n_1909),
.B(n_1911),
.Y(n_1963)
);

NAND2xp5_ASAP7_75t_L g1964 ( 
.A(n_1951),
.B(n_1926),
.Y(n_1964)
);

INVx1_ASAP7_75t_L g1965 ( 
.A(n_1957),
.Y(n_1965)
);

OR2x2_ASAP7_75t_L g1966 ( 
.A(n_1963),
.B(n_1944),
.Y(n_1966)
);

AND2x2_ASAP7_75t_L g1967 ( 
.A(n_1958),
.B(n_1936),
.Y(n_1967)
);

INVx2_ASAP7_75t_L g1968 ( 
.A(n_1960),
.Y(n_1968)
);

AND2x2_ASAP7_75t_L g1969 ( 
.A(n_1961),
.B(n_1954),
.Y(n_1969)
);

INVx1_ASAP7_75t_L g1970 ( 
.A(n_1959),
.Y(n_1970)
);

AND2x2_ASAP7_75t_L g1971 ( 
.A(n_1967),
.B(n_1940),
.Y(n_1971)
);

INVx1_ASAP7_75t_L g1972 ( 
.A(n_1965),
.Y(n_1972)
);

INVx2_ASAP7_75t_SL g1973 ( 
.A(n_1967),
.Y(n_1973)
);

OR2x2_ASAP7_75t_L g1974 ( 
.A(n_1966),
.B(n_1942),
.Y(n_1974)
);

INVx2_ASAP7_75t_L g1975 ( 
.A(n_1968),
.Y(n_1975)
);

OA21x2_ASAP7_75t_L g1976 ( 
.A1(n_1968),
.A2(n_1956),
.B(n_1962),
.Y(n_1976)
);

OR2x2_ASAP7_75t_L g1977 ( 
.A(n_1970),
.B(n_1953),
.Y(n_1977)
);

NAND2xp5_ASAP7_75t_SL g1978 ( 
.A(n_1969),
.B(n_1922),
.Y(n_1978)
);

INVx1_ASAP7_75t_L g1979 ( 
.A(n_1969),
.Y(n_1979)
);

INVx1_ASAP7_75t_L g1980 ( 
.A(n_1975),
.Y(n_1980)
);

INVx1_ASAP7_75t_L g1981 ( 
.A(n_1975),
.Y(n_1981)
);

INVx2_ASAP7_75t_L g1982 ( 
.A(n_1973),
.Y(n_1982)
);

OAI211xp5_ASAP7_75t_L g1983 ( 
.A1(n_1976),
.A2(n_1854),
.B(n_1880),
.C(n_1878),
.Y(n_1983)
);

OAI21xp5_ASAP7_75t_L g1984 ( 
.A1(n_1976),
.A2(n_1857),
.B(n_1875),
.Y(n_1984)
);

INVx2_ASAP7_75t_SL g1985 ( 
.A(n_1974),
.Y(n_1985)
);

INVx2_ASAP7_75t_L g1986 ( 
.A(n_1976),
.Y(n_1986)
);

AND2x2_ASAP7_75t_L g1987 ( 
.A(n_1971),
.B(n_1940),
.Y(n_1987)
);

AOI21xp33_ASAP7_75t_SL g1988 ( 
.A1(n_1978),
.A2(n_1922),
.B(n_1932),
.Y(n_1988)
);

INVx2_ASAP7_75t_L g1989 ( 
.A(n_1977),
.Y(n_1989)
);

OR2x2_ASAP7_75t_L g1990 ( 
.A(n_1979),
.B(n_1953),
.Y(n_1990)
);

INVx2_ASAP7_75t_L g1991 ( 
.A(n_1987),
.Y(n_1991)
);

OR2x2_ASAP7_75t_L g1992 ( 
.A(n_1985),
.B(n_1989),
.Y(n_1992)
);

INVx1_ASAP7_75t_L g1993 ( 
.A(n_1980),
.Y(n_1993)
);

INVx1_ASAP7_75t_L g1994 ( 
.A(n_1981),
.Y(n_1994)
);

AOI22xp33_ASAP7_75t_L g1995 ( 
.A1(n_1984),
.A2(n_1978),
.B1(n_1972),
.B2(n_1909),
.Y(n_1995)
);

INVx2_ASAP7_75t_L g1996 ( 
.A(n_1986),
.Y(n_1996)
);

INVx1_ASAP7_75t_L g1997 ( 
.A(n_1982),
.Y(n_1997)
);

INVxp67_ASAP7_75t_L g1998 ( 
.A(n_1986),
.Y(n_1998)
);

OAI21xp5_ASAP7_75t_L g1999 ( 
.A1(n_1995),
.A2(n_1984),
.B(n_1983),
.Y(n_1999)
);

O2A1O1Ixp33_ASAP7_75t_L g2000 ( 
.A1(n_1998),
.A2(n_1983),
.B(n_1988),
.C(n_1982),
.Y(n_2000)
);

INVx1_ASAP7_75t_L g2001 ( 
.A(n_1996),
.Y(n_2001)
);

INVxp67_ASAP7_75t_L g2002 ( 
.A(n_1992),
.Y(n_2002)
);

AOI22xp33_ASAP7_75t_SL g2003 ( 
.A1(n_1999),
.A2(n_1991),
.B1(n_2002),
.B2(n_1997),
.Y(n_2003)
);

INVx1_ASAP7_75t_SL g2004 ( 
.A(n_2001),
.Y(n_2004)
);

NAND2xp5_ASAP7_75t_L g2005 ( 
.A(n_2000),
.B(n_1998),
.Y(n_2005)
);

NAND2xp5_ASAP7_75t_L g2006 ( 
.A(n_2002),
.B(n_1993),
.Y(n_2006)
);

NAND3xp33_ASAP7_75t_L g2007 ( 
.A(n_2005),
.B(n_1994),
.C(n_1990),
.Y(n_2007)
);

INVx1_ASAP7_75t_L g2008 ( 
.A(n_2006),
.Y(n_2008)
);

NOR3xp33_ASAP7_75t_L g2009 ( 
.A(n_2003),
.B(n_1840),
.C(n_1824),
.Y(n_2009)
);

NAND3xp33_ASAP7_75t_L g2010 ( 
.A(n_2004),
.B(n_1787),
.C(n_1796),
.Y(n_2010)
);

AOI22xp5_ASAP7_75t_L g2011 ( 
.A1(n_2005),
.A2(n_1914),
.B1(n_1933),
.B2(n_1932),
.Y(n_2011)
);

NAND2xp5_ASAP7_75t_L g2012 ( 
.A(n_2009),
.B(n_1943),
.Y(n_2012)
);

INVx1_ASAP7_75t_L g2013 ( 
.A(n_2007),
.Y(n_2013)
);

OAI22xp5_ASAP7_75t_L g2014 ( 
.A1(n_2011),
.A2(n_1914),
.B1(n_1923),
.B2(n_1777),
.Y(n_2014)
);

OR2x2_ASAP7_75t_L g2015 ( 
.A(n_2008),
.B(n_1928),
.Y(n_2015)
);

AND2x2_ASAP7_75t_L g2016 ( 
.A(n_2010),
.B(n_1943),
.Y(n_2016)
);

NOR2xp33_ASAP7_75t_L g2017 ( 
.A(n_2007),
.B(n_1906),
.Y(n_2017)
);

INVx1_ASAP7_75t_L g2018 ( 
.A(n_2007),
.Y(n_2018)
);

NAND2xp5_ASAP7_75t_L g2019 ( 
.A(n_2009),
.B(n_1964),
.Y(n_2019)
);

NOR2xp33_ASAP7_75t_L g2020 ( 
.A(n_2007),
.B(n_1897),
.Y(n_2020)
);

NAND2xp5_ASAP7_75t_L g2021 ( 
.A(n_2009),
.B(n_1964),
.Y(n_2021)
);

AOI21xp33_ASAP7_75t_L g2022 ( 
.A1(n_2020),
.A2(n_1787),
.B(n_1788),
.Y(n_2022)
);

AOI221x1_ASAP7_75t_L g2023 ( 
.A1(n_2013),
.A2(n_2018),
.B1(n_2017),
.B2(n_2014),
.C(n_2012),
.Y(n_2023)
);

NAND4xp25_ASAP7_75t_L g2024 ( 
.A(n_2015),
.B(n_1901),
.C(n_1931),
.D(n_1890),
.Y(n_2024)
);

AOI211xp5_ASAP7_75t_L g2025 ( 
.A1(n_2016),
.A2(n_1783),
.B(n_1785),
.C(n_1829),
.Y(n_2025)
);

NAND2xp5_ASAP7_75t_L g2026 ( 
.A(n_2019),
.B(n_1952),
.Y(n_2026)
);

OAI221xp5_ASAP7_75t_L g2027 ( 
.A1(n_2021),
.A2(n_1898),
.B1(n_1873),
.B2(n_1862),
.C(n_1892),
.Y(n_2027)
);

OAI21xp5_ASAP7_75t_L g2028 ( 
.A1(n_2013),
.A2(n_1825),
.B(n_1800),
.Y(n_2028)
);

OAI21xp33_ASAP7_75t_L g2029 ( 
.A1(n_2020),
.A2(n_1892),
.B(n_1893),
.Y(n_2029)
);

NAND4xp25_ASAP7_75t_L g2030 ( 
.A(n_2017),
.B(n_1893),
.C(n_1886),
.D(n_1884),
.Y(n_2030)
);

OAI221xp5_ASAP7_75t_L g2031 ( 
.A1(n_2013),
.A2(n_1809),
.B1(n_1900),
.B2(n_1925),
.C(n_1844),
.Y(n_2031)
);

OAI211xp5_ASAP7_75t_L g2032 ( 
.A1(n_2013),
.A2(n_1803),
.B(n_193),
.C(n_194),
.Y(n_2032)
);

NAND2xp5_ASAP7_75t_L g2033 ( 
.A(n_2023),
.B(n_1946),
.Y(n_2033)
);

NOR3xp33_ASAP7_75t_L g2034 ( 
.A(n_2032),
.B(n_1843),
.C(n_1786),
.Y(n_2034)
);

NAND2xp5_ASAP7_75t_L g2035 ( 
.A(n_2025),
.B(n_1947),
.Y(n_2035)
);

NAND2xp5_ASAP7_75t_L g2036 ( 
.A(n_2028),
.B(n_1947),
.Y(n_2036)
);

INVx1_ASAP7_75t_SL g2037 ( 
.A(n_2026),
.Y(n_2037)
);

NAND3xp33_ASAP7_75t_L g2038 ( 
.A(n_2031),
.B(n_1782),
.C(n_1786),
.Y(n_2038)
);

NAND2xp5_ASAP7_75t_L g2039 ( 
.A(n_2029),
.B(n_1938),
.Y(n_2039)
);

NAND2xp5_ASAP7_75t_L g2040 ( 
.A(n_2022),
.B(n_1938),
.Y(n_2040)
);

NOR2x1_ASAP7_75t_L g2041 ( 
.A(n_2030),
.B(n_1801),
.Y(n_2041)
);

NAND2xp5_ASAP7_75t_L g2042 ( 
.A(n_2024),
.B(n_1945),
.Y(n_2042)
);

XOR2xp5_ASAP7_75t_L g2043 ( 
.A(n_2033),
.B(n_2041),
.Y(n_2043)
);

AND2x2_ASAP7_75t_SL g2044 ( 
.A(n_2042),
.B(n_1801),
.Y(n_2044)
);

NOR2x1p5_ASAP7_75t_L g2045 ( 
.A(n_2039),
.B(n_2038),
.Y(n_2045)
);

OR2x2_ASAP7_75t_L g2046 ( 
.A(n_2037),
.B(n_2027),
.Y(n_2046)
);

AND2x2_ASAP7_75t_L g2047 ( 
.A(n_2035),
.B(n_1950),
.Y(n_2047)
);

NAND4xp75_ASAP7_75t_L g2048 ( 
.A(n_2040),
.B(n_192),
.C(n_194),
.D(n_195),
.Y(n_2048)
);

NOR2x1_ASAP7_75t_L g2049 ( 
.A(n_2036),
.B(n_195),
.Y(n_2049)
);

AND2x4_ASAP7_75t_L g2050 ( 
.A(n_2045),
.B(n_2034),
.Y(n_2050)
);

NOR3xp33_ASAP7_75t_SL g2051 ( 
.A(n_2048),
.B(n_196),
.C(n_197),
.Y(n_2051)
);

AOI322xp5_ASAP7_75t_L g2052 ( 
.A1(n_2044),
.A2(n_1954),
.A3(n_1948),
.B1(n_1955),
.B2(n_1951),
.C1(n_1924),
.C2(n_1802),
.Y(n_2052)
);

OR2x2_ASAP7_75t_L g2053 ( 
.A(n_2046),
.B(n_1955),
.Y(n_2053)
);

NOR3xp33_ASAP7_75t_L g2054 ( 
.A(n_2049),
.B(n_1802),
.C(n_1811),
.Y(n_2054)
);

NAND3xp33_ASAP7_75t_L g2055 ( 
.A(n_2047),
.B(n_196),
.C(n_198),
.Y(n_2055)
);

AND2x4_ASAP7_75t_L g2056 ( 
.A(n_2043),
.B(n_1940),
.Y(n_2056)
);

INVx2_ASAP7_75t_L g2057 ( 
.A(n_2056),
.Y(n_2057)
);

INVx1_ASAP7_75t_L g2058 ( 
.A(n_2055),
.Y(n_2058)
);

NOR2xp33_ASAP7_75t_L g2059 ( 
.A(n_2050),
.B(n_198),
.Y(n_2059)
);

INVx1_ASAP7_75t_L g2060 ( 
.A(n_2051),
.Y(n_2060)
);

INVx2_ASAP7_75t_L g2061 ( 
.A(n_2053),
.Y(n_2061)
);

OAI22xp5_ASAP7_75t_SL g2062 ( 
.A1(n_2060),
.A2(n_2054),
.B1(n_1821),
.B2(n_1811),
.Y(n_2062)
);

AOI221xp5_ASAP7_75t_L g2063 ( 
.A1(n_2059),
.A2(n_2058),
.B1(n_2057),
.B2(n_2061),
.C(n_2052),
.Y(n_2063)
);

NAND2xp5_ASAP7_75t_L g2064 ( 
.A(n_2059),
.B(n_199),
.Y(n_2064)
);

OAI221xp5_ASAP7_75t_L g2065 ( 
.A1(n_2059),
.A2(n_1900),
.B1(n_1837),
.B2(n_1823),
.C(n_1925),
.Y(n_2065)
);

NAND3xp33_ASAP7_75t_SL g2066 ( 
.A(n_2063),
.B(n_199),
.C(n_200),
.Y(n_2066)
);

NOR3xp33_ASAP7_75t_L g2067 ( 
.A(n_2064),
.B(n_200),
.C(n_201),
.Y(n_2067)
);

AOI221xp5_ASAP7_75t_SL g2068 ( 
.A1(n_2062),
.A2(n_2065),
.B1(n_202),
.B2(n_203),
.C(n_204),
.Y(n_2068)
);

NAND2xp5_ASAP7_75t_L g2069 ( 
.A(n_2063),
.B(n_201),
.Y(n_2069)
);

OR3x1_ASAP7_75t_L g2070 ( 
.A(n_2063),
.B(n_202),
.C(n_203),
.Y(n_2070)
);

AND4x1_ASAP7_75t_L g2071 ( 
.A(n_2069),
.B(n_204),
.C(n_205),
.D(n_206),
.Y(n_2071)
);

INVx1_ASAP7_75t_L g2072 ( 
.A(n_2070),
.Y(n_2072)
);

AOI22xp33_ASAP7_75t_L g2073 ( 
.A1(n_2066),
.A2(n_1933),
.B1(n_1821),
.B2(n_1813),
.Y(n_2073)
);

AOI22xp5_ASAP7_75t_L g2074 ( 
.A1(n_2067),
.A2(n_1933),
.B1(n_1883),
.B2(n_1813),
.Y(n_2074)
);

NAND2xp5_ASAP7_75t_SL g2075 ( 
.A(n_2071),
.B(n_2068),
.Y(n_2075)
);

INVx1_ASAP7_75t_L g2076 ( 
.A(n_2072),
.Y(n_2076)
);

NAND2xp5_ASAP7_75t_L g2077 ( 
.A(n_2074),
.B(n_2073),
.Y(n_2077)
);

AOI22xp5_ASAP7_75t_L g2078 ( 
.A1(n_2076),
.A2(n_1933),
.B1(n_1813),
.B2(n_1948),
.Y(n_2078)
);

AOI22xp33_ASAP7_75t_L g2079 ( 
.A1(n_2075),
.A2(n_1909),
.B1(n_1874),
.B2(n_1945),
.Y(n_2079)
);

XNOR2xp5_ASAP7_75t_L g2080 ( 
.A(n_2077),
.B(n_206),
.Y(n_2080)
);

NAND2xp5_ASAP7_75t_L g2081 ( 
.A(n_2080),
.B(n_207),
.Y(n_2081)
);

NAND2xp5_ASAP7_75t_L g2082 ( 
.A(n_2078),
.B(n_207),
.Y(n_2082)
);

AOI21xp33_ASAP7_75t_L g2083 ( 
.A1(n_2081),
.A2(n_2079),
.B(n_209),
.Y(n_2083)
);

AO221x2_ASAP7_75t_L g2084 ( 
.A1(n_2083),
.A2(n_2082),
.B1(n_209),
.B2(n_212),
.C(n_213),
.Y(n_2084)
);

OAI22xp5_ASAP7_75t_L g2085 ( 
.A1(n_2084),
.A2(n_208),
.B1(n_212),
.B2(n_214),
.Y(n_2085)
);

AOI211xp5_ASAP7_75t_L g2086 ( 
.A1(n_2085),
.A2(n_208),
.B(n_214),
.C(n_215),
.Y(n_2086)
);


endmodule