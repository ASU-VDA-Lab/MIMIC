module fake_jpeg_19752_n_311 (n_3, n_2, n_1, n_0, n_10, n_4, n_8, n_9, n_6, n_5, n_7, n_311);

input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_311;

wire n_253;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_15;
wire n_141;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_13;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_11;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_14;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_18;
wire n_145;
wire n_20;
wire n_303;
wire n_259;
wire n_90;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_12;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_208;
wire n_308;
wire n_297;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

CKINVDCx20_ASAP7_75t_R g11 ( 
.A(n_0),
.Y(n_11)
);

BUFx6f_ASAP7_75t_L g12 ( 
.A(n_7),
.Y(n_12)
);

CKINVDCx20_ASAP7_75t_R g13 ( 
.A(n_6),
.Y(n_13)
);

INVx4_ASAP7_75t_L g14 ( 
.A(n_3),
.Y(n_14)
);

BUFx16f_ASAP7_75t_L g15 ( 
.A(n_4),
.Y(n_15)
);

INVx2_ASAP7_75t_L g16 ( 
.A(n_10),
.Y(n_16)
);

BUFx24_ASAP7_75t_L g17 ( 
.A(n_7),
.Y(n_17)
);

BUFx4f_ASAP7_75t_SL g18 ( 
.A(n_9),
.Y(n_18)
);

BUFx12_ASAP7_75t_L g19 ( 
.A(n_8),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_6),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_10),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_0),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_7),
.Y(n_23)
);

BUFx3_ASAP7_75t_L g24 ( 
.A(n_17),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_24),
.Y(n_42)
);

INVx5_ASAP7_75t_L g25 ( 
.A(n_17),
.Y(n_25)
);

INVx3_ASAP7_75t_L g36 ( 
.A(n_25),
.Y(n_36)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_18),
.Y(n_26)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_26),
.Y(n_40)
);

INVx2_ASAP7_75t_L g27 ( 
.A(n_22),
.Y(n_27)
);

INVx3_ASAP7_75t_L g38 ( 
.A(n_27),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_L g28 ( 
.A(n_16),
.B(n_13),
.Y(n_28)
);

NAND2xp5_ASAP7_75t_SL g43 ( 
.A(n_28),
.B(n_29),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g29 ( 
.A(n_16),
.B(n_10),
.Y(n_29)
);

NOR2xp33_ASAP7_75t_L g30 ( 
.A(n_16),
.B(n_10),
.Y(n_30)
);

NAND2xp5_ASAP7_75t_L g44 ( 
.A(n_30),
.B(n_33),
.Y(n_44)
);

BUFx3_ASAP7_75t_L g31 ( 
.A(n_17),
.Y(n_31)
);

INVx3_ASAP7_75t_L g39 ( 
.A(n_31),
.Y(n_39)
);

INVx4_ASAP7_75t_L g32 ( 
.A(n_14),
.Y(n_32)
);

INVx3_ASAP7_75t_L g41 ( 
.A(n_32),
.Y(n_41)
);

AND2x2_ASAP7_75t_L g33 ( 
.A(n_15),
.B(n_0),
.Y(n_33)
);

AOI22xp5_ASAP7_75t_L g34 ( 
.A1(n_16),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_34)
);

AOI22xp33_ASAP7_75t_SL g35 ( 
.A1(n_34),
.A2(n_17),
.B1(n_14),
.B2(n_11),
.Y(n_35)
);

AOI22xp5_ASAP7_75t_L g51 ( 
.A1(n_35),
.A2(n_37),
.B1(n_33),
.B2(n_26),
.Y(n_51)
);

AOI22xp33_ASAP7_75t_L g37 ( 
.A1(n_27),
.A2(n_14),
.B1(n_17),
.B2(n_11),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g45 ( 
.A(n_43),
.B(n_28),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_SL g75 ( 
.A(n_45),
.B(n_54),
.Y(n_75)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_40),
.Y(n_46)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_46),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_L g47 ( 
.A(n_44),
.B(n_43),
.Y(n_47)
);

NAND2xp5_ASAP7_75t_L g67 ( 
.A(n_47),
.B(n_53),
.Y(n_67)
);

INVx11_ASAP7_75t_L g48 ( 
.A(n_42),
.Y(n_48)
);

INVx3_ASAP7_75t_SL g65 ( 
.A(n_48),
.Y(n_65)
);

INVx3_ASAP7_75t_L g49 ( 
.A(n_41),
.Y(n_49)
);

INVx2_ASAP7_75t_L g69 ( 
.A(n_49),
.Y(n_69)
);

INVx11_ASAP7_75t_L g50 ( 
.A(n_42),
.Y(n_50)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_50),
.Y(n_78)
);

OAI22xp5_ASAP7_75t_L g62 ( 
.A1(n_51),
.A2(n_60),
.B1(n_25),
.B2(n_26),
.Y(n_62)
);

INVx4_ASAP7_75t_L g52 ( 
.A(n_42),
.Y(n_52)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_52),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_L g53 ( 
.A(n_44),
.B(n_33),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_44),
.B(n_28),
.Y(n_54)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_40),
.Y(n_55)
);

CKINVDCx20_ASAP7_75t_R g70 ( 
.A(n_55),
.Y(n_70)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_40),
.Y(n_56)
);

AND2x2_ASAP7_75t_SL g72 ( 
.A(n_56),
.B(n_59),
.Y(n_72)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_41),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_57),
.B(n_58),
.Y(n_63)
);

INVx4_ASAP7_75t_L g58 ( 
.A(n_42),
.Y(n_58)
);

AND2x2_ASAP7_75t_L g59 ( 
.A(n_35),
.B(n_33),
.Y(n_59)
);

AOI22xp33_ASAP7_75t_SL g60 ( 
.A1(n_36),
.A2(n_17),
.B1(n_25),
.B2(n_14),
.Y(n_60)
);

AOI22xp5_ASAP7_75t_L g81 ( 
.A1(n_62),
.A2(n_71),
.B1(n_74),
.B2(n_76),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_45),
.B(n_30),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_L g79 ( 
.A(n_64),
.B(n_47),
.Y(n_79)
);

INVxp67_ASAP7_75t_L g66 ( 
.A(n_60),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_66),
.B(n_36),
.Y(n_85)
);

INVx2_ASAP7_75t_R g68 ( 
.A(n_46),
.Y(n_68)
);

INVx1_ASAP7_75t_SL g83 ( 
.A(n_68),
.Y(n_83)
);

OAI22xp5_ASAP7_75t_SL g71 ( 
.A1(n_51),
.A2(n_27),
.B1(n_34),
.B2(n_38),
.Y(n_71)
);

OAI22xp5_ASAP7_75t_SL g74 ( 
.A1(n_51),
.A2(n_27),
.B1(n_34),
.B2(n_38),
.Y(n_74)
);

AOI22xp33_ASAP7_75t_L g76 ( 
.A1(n_59),
.A2(n_38),
.B1(n_32),
.B2(n_25),
.Y(n_76)
);

NAND2x1_ASAP7_75t_SL g77 ( 
.A(n_59),
.B(n_17),
.Y(n_77)
);

OAI21xp5_ASAP7_75t_L g84 ( 
.A1(n_77),
.A2(n_59),
.B(n_33),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g103 ( 
.A(n_79),
.B(n_90),
.Y(n_103)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_63),
.Y(n_80)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_80),
.Y(n_105)
);

OAI22xp5_ASAP7_75t_SL g82 ( 
.A1(n_71),
.A2(n_59),
.B1(n_47),
.B2(n_54),
.Y(n_82)
);

AOI22xp5_ASAP7_75t_L g106 ( 
.A1(n_82),
.A2(n_88),
.B1(n_74),
.B2(n_71),
.Y(n_106)
);

OAI21xp5_ASAP7_75t_L g100 ( 
.A1(n_84),
.A2(n_97),
.B(n_96),
.Y(n_100)
);

INVxp67_ASAP7_75t_L g101 ( 
.A(n_85),
.Y(n_101)
);

CKINVDCx20_ASAP7_75t_R g86 ( 
.A(n_61),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_86),
.B(n_89),
.Y(n_108)
);

INVx3_ASAP7_75t_L g87 ( 
.A(n_69),
.Y(n_87)
);

INVx2_ASAP7_75t_SL g109 ( 
.A(n_87),
.Y(n_109)
);

AOI22xp33_ASAP7_75t_L g88 ( 
.A1(n_68),
.A2(n_46),
.B1(n_56),
.B2(n_55),
.Y(n_88)
);

CKINVDCx20_ASAP7_75t_R g89 ( 
.A(n_61),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g90 ( 
.A(n_67),
.B(n_53),
.Y(n_90)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_63),
.Y(n_91)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_91),
.Y(n_107)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_73),
.Y(n_92)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_92),
.Y(n_114)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_73),
.Y(n_93)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_93),
.Y(n_117)
);

XNOR2xp5_ASAP7_75t_L g94 ( 
.A(n_67),
.B(n_53),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_SL g115 ( 
.A(n_94),
.B(n_96),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_75),
.B(n_56),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g113 ( 
.A(n_95),
.B(n_97),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_L g96 ( 
.A(n_67),
.B(n_55),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g97 ( 
.A(n_75),
.B(n_33),
.Y(n_97)
);

CKINVDCx20_ASAP7_75t_R g98 ( 
.A(n_92),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_SL g136 ( 
.A(n_98),
.B(n_99),
.Y(n_136)
);

CKINVDCx16_ASAP7_75t_R g99 ( 
.A(n_95),
.Y(n_99)
);

XNOR2xp5_ASAP7_75t_SL g122 ( 
.A(n_100),
.B(n_94),
.Y(n_122)
);

AOI22xp5_ASAP7_75t_SL g102 ( 
.A1(n_84),
.A2(n_62),
.B1(n_77),
.B2(n_76),
.Y(n_102)
);

OAI21xp5_ASAP7_75t_L g135 ( 
.A1(n_102),
.A2(n_78),
.B(n_29),
.Y(n_135)
);

OAI21xp5_ASAP7_75t_L g104 ( 
.A1(n_86),
.A2(n_68),
.B(n_72),
.Y(n_104)
);

AOI21xp5_ASAP7_75t_L g129 ( 
.A1(n_104),
.A2(n_83),
.B(n_70),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_L g148 ( 
.A(n_106),
.B(n_112),
.Y(n_148)
);

AOI21xp5_ASAP7_75t_SL g110 ( 
.A1(n_85),
.A2(n_68),
.B(n_72),
.Y(n_110)
);

OAI21xp5_ASAP7_75t_SL g138 ( 
.A1(n_110),
.A2(n_111),
.B(n_119),
.Y(n_138)
);

AOI21xp5_ASAP7_75t_L g111 ( 
.A1(n_82),
.A2(n_72),
.B(n_77),
.Y(n_111)
);

INVxp67_ASAP7_75t_L g112 ( 
.A(n_88),
.Y(n_112)
);

CKINVDCx20_ASAP7_75t_R g116 ( 
.A(n_93),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_L g153 ( 
.A(n_116),
.B(n_118),
.Y(n_153)
);

INVxp67_ASAP7_75t_L g118 ( 
.A(n_79),
.Y(n_118)
);

AOI21xp5_ASAP7_75t_L g119 ( 
.A1(n_80),
.A2(n_72),
.B(n_77),
.Y(n_119)
);

INVxp67_ASAP7_75t_L g120 ( 
.A(n_81),
.Y(n_120)
);

INVxp67_ASAP7_75t_L g123 ( 
.A(n_120),
.Y(n_123)
);

O2A1O1Ixp33_ASAP7_75t_L g121 ( 
.A1(n_89),
.A2(n_70),
.B(n_74),
.C(n_72),
.Y(n_121)
);

OAI21xp5_ASAP7_75t_SL g139 ( 
.A1(n_121),
.A2(n_37),
.B(n_31),
.Y(n_139)
);

XNOR2xp5_ASAP7_75t_L g162 ( 
.A(n_122),
.B(n_124),
.Y(n_162)
);

XNOR2xp5_ASAP7_75t_SL g124 ( 
.A(n_100),
.B(n_94),
.Y(n_124)
);

XOR2xp5_ASAP7_75t_L g160 ( 
.A(n_124),
.B(n_146),
.Y(n_160)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_108),
.Y(n_125)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_125),
.Y(n_161)
);

MAJIxp5_ASAP7_75t_L g126 ( 
.A(n_111),
.B(n_90),
.C(n_81),
.Y(n_126)
);

MAJIxp5_ASAP7_75t_L g154 ( 
.A(n_126),
.B(n_127),
.C(n_102),
.Y(n_154)
);

MAJIxp5_ASAP7_75t_L g127 ( 
.A(n_119),
.B(n_91),
.C(n_64),
.Y(n_127)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_108),
.Y(n_128)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_128),
.Y(n_163)
);

OAI21xp5_ASAP7_75t_L g182 ( 
.A1(n_129),
.A2(n_132),
.B(n_24),
.Y(n_182)
);

INVxp67_ASAP7_75t_L g130 ( 
.A(n_110),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_L g169 ( 
.A(n_130),
.B(n_134),
.Y(n_169)
);

AOI22xp5_ASAP7_75t_L g131 ( 
.A1(n_121),
.A2(n_83),
.B1(n_87),
.B2(n_78),
.Y(n_131)
);

OAI22xp5_ASAP7_75t_SL g174 ( 
.A1(n_131),
.A2(n_101),
.B1(n_109),
.B2(n_65),
.Y(n_174)
);

AOI21xp5_ASAP7_75t_L g132 ( 
.A1(n_104),
.A2(n_83),
.B(n_69),
.Y(n_132)
);

OAI22xp5_ASAP7_75t_L g133 ( 
.A1(n_99),
.A2(n_34),
.B1(n_78),
.B2(n_87),
.Y(n_133)
);

OAI22xp5_ASAP7_75t_L g171 ( 
.A1(n_133),
.A2(n_150),
.B1(n_98),
.B2(n_109),
.Y(n_171)
);

NOR2xp33_ASAP7_75t_SL g134 ( 
.A(n_113),
.B(n_29),
.Y(n_134)
);

AOI21xp5_ASAP7_75t_L g158 ( 
.A1(n_135),
.A2(n_104),
.B(n_136),
.Y(n_158)
);

CKINVDCx20_ASAP7_75t_R g137 ( 
.A(n_114),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_L g170 ( 
.A(n_137),
.B(n_141),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_L g156 ( 
.A(n_139),
.B(n_147),
.Y(n_156)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_114),
.Y(n_140)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_140),
.Y(n_165)
);

INVxp67_ASAP7_75t_L g141 ( 
.A(n_110),
.Y(n_141)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_117),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_L g179 ( 
.A(n_142),
.B(n_144),
.Y(n_179)
);

AOI22xp33_ASAP7_75t_L g143 ( 
.A1(n_105),
.A2(n_69),
.B1(n_65),
.B2(n_58),
.Y(n_143)
);

OAI22xp33_ASAP7_75t_SL g175 ( 
.A1(n_143),
.A2(n_109),
.B1(n_36),
.B2(n_39),
.Y(n_175)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_117),
.Y(n_144)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_105),
.Y(n_145)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_145),
.Y(n_181)
);

XOR2xp5_ASAP7_75t_L g146 ( 
.A(n_113),
.B(n_30),
.Y(n_146)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_107),
.Y(n_147)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_107),
.Y(n_149)
);

CKINVDCx20_ASAP7_75t_R g168 ( 
.A(n_149),
.Y(n_168)
);

OAI22xp5_ASAP7_75t_L g150 ( 
.A1(n_106),
.A2(n_65),
.B1(n_58),
.B2(n_52),
.Y(n_150)
);

BUFx24_ASAP7_75t_SL g151 ( 
.A(n_103),
.Y(n_151)
);

NOR2xp33_ASAP7_75t_L g166 ( 
.A(n_151),
.B(n_116),
.Y(n_166)
);

OAI22xp5_ASAP7_75t_SL g152 ( 
.A1(n_121),
.A2(n_65),
.B1(n_52),
.B2(n_57),
.Y(n_152)
);

AOI22xp5_ASAP7_75t_L g167 ( 
.A1(n_152),
.A2(n_147),
.B1(n_145),
.B2(n_123),
.Y(n_167)
);

XOR2xp5_ASAP7_75t_L g193 ( 
.A(n_154),
.B(n_162),
.Y(n_193)
);

CKINVDCx16_ASAP7_75t_R g155 ( 
.A(n_125),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_L g197 ( 
.A(n_155),
.B(n_166),
.Y(n_197)
);

MAJIxp5_ASAP7_75t_L g157 ( 
.A(n_127),
.B(n_102),
.C(n_115),
.Y(n_157)
);

MAJIxp5_ASAP7_75t_L g185 ( 
.A(n_157),
.B(n_177),
.C(n_132),
.Y(n_185)
);

XNOR2xp5_ASAP7_75t_L g201 ( 
.A(n_158),
.B(n_148),
.Y(n_201)
);

XOR2xp5_ASAP7_75t_SL g159 ( 
.A(n_138),
.B(n_103),
.Y(n_159)
);

AOI22xp5_ASAP7_75t_SL g207 ( 
.A1(n_159),
.A2(n_178),
.B1(n_32),
.B2(n_11),
.Y(n_207)
);

NAND4xp25_ASAP7_75t_SL g164 ( 
.A(n_128),
.B(n_19),
.C(n_49),
.D(n_57),
.Y(n_164)
);

CKINVDCx20_ASAP7_75t_R g187 ( 
.A(n_164),
.Y(n_187)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_167),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_L g202 ( 
.A(n_171),
.B(n_172),
.Y(n_202)
);

INVxp67_ASAP7_75t_L g172 ( 
.A(n_153),
.Y(n_172)
);

XNOR2xp5_ASAP7_75t_L g173 ( 
.A(n_122),
.B(n_115),
.Y(n_173)
);

XOR2xp5_ASAP7_75t_L g194 ( 
.A(n_173),
.B(n_180),
.Y(n_194)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_174),
.Y(n_189)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_175),
.Y(n_191)
);

AND2x2_ASAP7_75t_L g176 ( 
.A(n_131),
.B(n_31),
.Y(n_176)
);

OAI21xp5_ASAP7_75t_L g192 ( 
.A1(n_176),
.A2(n_182),
.B(n_139),
.Y(n_192)
);

MAJIxp5_ASAP7_75t_L g177 ( 
.A(n_126),
.B(n_49),
.C(n_39),
.Y(n_177)
);

XOR2x2_ASAP7_75t_L g178 ( 
.A(n_138),
.B(n_109),
.Y(n_178)
);

XOR2xp5_ASAP7_75t_L g180 ( 
.A(n_135),
.B(n_32),
.Y(n_180)
);

NOR2xp33_ASAP7_75t_L g184 ( 
.A(n_169),
.B(n_153),
.Y(n_184)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_184),
.Y(n_212)
);

XOR2xp5_ASAP7_75t_L g214 ( 
.A(n_185),
.B(n_204),
.Y(n_214)
);

AND2x6_ASAP7_75t_L g186 ( 
.A(n_178),
.B(n_130),
.Y(n_186)
);

OAI21xp5_ASAP7_75t_SL g211 ( 
.A1(n_186),
.A2(n_159),
.B(n_172),
.Y(n_211)
);

NOR3xp33_ASAP7_75t_L g188 ( 
.A(n_161),
.B(n_141),
.C(n_129),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_L g210 ( 
.A(n_188),
.B(n_196),
.Y(n_210)
);

MAJIxp5_ASAP7_75t_L g190 ( 
.A(n_157),
.B(n_146),
.C(n_140),
.Y(n_190)
);

MAJIxp5_ASAP7_75t_L g209 ( 
.A(n_190),
.B(n_195),
.C(n_206),
.Y(n_209)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_192),
.Y(n_216)
);

MAJIxp5_ASAP7_75t_L g195 ( 
.A(n_154),
.B(n_148),
.C(n_152),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_SL g196 ( 
.A(n_163),
.B(n_123),
.Y(n_196)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_179),
.Y(n_198)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_198),
.Y(n_221)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_170),
.Y(n_199)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_199),
.Y(n_224)
);

HB1xp67_ASAP7_75t_L g200 ( 
.A(n_164),
.Y(n_200)
);

INVxp33_ASAP7_75t_SL g220 ( 
.A(n_200),
.Y(n_220)
);

XNOR2xp5_ASAP7_75t_SL g208 ( 
.A(n_201),
.B(n_207),
.Y(n_208)
);

NOR2xp33_ASAP7_75t_L g203 ( 
.A(n_168),
.B(n_13),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_L g219 ( 
.A(n_203),
.B(n_205),
.Y(n_219)
);

XOR2xp5_ASAP7_75t_L g204 ( 
.A(n_162),
.B(n_19),
.Y(n_204)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_165),
.Y(n_205)
);

MAJIxp5_ASAP7_75t_L g206 ( 
.A(n_160),
.B(n_39),
.C(n_41),
.Y(n_206)
);

OAI21xp5_ASAP7_75t_SL g246 ( 
.A1(n_211),
.A2(n_19),
.B(n_48),
.Y(n_246)
);

XNOR2xp5_ASAP7_75t_L g213 ( 
.A(n_185),
.B(n_177),
.Y(n_213)
);

XNOR2xp5_ASAP7_75t_L g239 ( 
.A(n_213),
.B(n_19),
.Y(n_239)
);

AOI22xp5_ASAP7_75t_L g215 ( 
.A1(n_189),
.A2(n_174),
.B1(n_156),
.B2(n_176),
.Y(n_215)
);

OAI22xp5_ASAP7_75t_SL g234 ( 
.A1(n_215),
.A2(n_217),
.B1(n_192),
.B2(n_207),
.Y(n_234)
);

AOI22xp5_ASAP7_75t_L g217 ( 
.A1(n_183),
.A2(n_156),
.B1(n_176),
.B2(n_167),
.Y(n_217)
);

OAI22xp5_ASAP7_75t_SL g218 ( 
.A1(n_191),
.A2(n_158),
.B1(n_181),
.B2(n_182),
.Y(n_218)
);

AOI22xp5_ASAP7_75t_L g233 ( 
.A1(n_218),
.A2(n_228),
.B1(n_230),
.B2(n_187),
.Y(n_233)
);

MAJIxp5_ASAP7_75t_L g222 ( 
.A(n_190),
.B(n_160),
.C(n_173),
.Y(n_222)
);

NOR2xp33_ASAP7_75t_L g243 ( 
.A(n_222),
.B(n_225),
.Y(n_243)
);

XNOR2x2_ASAP7_75t_L g223 ( 
.A(n_186),
.B(n_180),
.Y(n_223)
);

XNOR2xp5_ASAP7_75t_SL g241 ( 
.A(n_223),
.B(n_19),
.Y(n_241)
);

MAJIxp5_ASAP7_75t_L g225 ( 
.A(n_206),
.B(n_193),
.C(n_195),
.Y(n_225)
);

MAJIxp5_ASAP7_75t_L g226 ( 
.A(n_193),
.B(n_15),
.C(n_22),
.Y(n_226)
);

XNOR2xp5_ASAP7_75t_L g231 ( 
.A(n_226),
.B(n_229),
.Y(n_231)
);

NAND2xp5_ASAP7_75t_L g227 ( 
.A(n_197),
.B(n_13),
.Y(n_227)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_227),
.Y(n_232)
);

OAI22xp5_ASAP7_75t_SL g228 ( 
.A1(n_202),
.A2(n_20),
.B1(n_21),
.B2(n_50),
.Y(n_228)
);

MAJIxp5_ASAP7_75t_L g229 ( 
.A(n_194),
.B(n_15),
.C(n_22),
.Y(n_229)
);

OAI22xp5_ASAP7_75t_SL g230 ( 
.A1(n_202),
.A2(n_20),
.B1(n_21),
.B2(n_50),
.Y(n_230)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_233),
.Y(n_260)
);

AOI22xp5_ASAP7_75t_L g254 ( 
.A1(n_234),
.A2(n_222),
.B1(n_9),
.B2(n_8),
.Y(n_254)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_219),
.Y(n_235)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_235),
.Y(n_261)
);

AOI22xp5_ASAP7_75t_L g236 ( 
.A1(n_212),
.A2(n_201),
.B1(n_194),
.B2(n_204),
.Y(n_236)
);

OAI22xp5_ASAP7_75t_SL g255 ( 
.A1(n_236),
.A2(n_240),
.B1(n_9),
.B2(n_8),
.Y(n_255)
);

XOR2xp5_ASAP7_75t_L g237 ( 
.A(n_214),
.B(n_19),
.Y(n_237)
);

XOR2xp5_ASAP7_75t_L g256 ( 
.A(n_237),
.B(n_239),
.Y(n_256)
);

INVx1_ASAP7_75t_SL g238 ( 
.A(n_220),
.Y(n_238)
);

NOR2xp33_ASAP7_75t_L g263 ( 
.A(n_238),
.B(n_242),
.Y(n_263)
);

AOI22xp5_ASAP7_75t_L g240 ( 
.A1(n_221),
.A2(n_210),
.B1(n_224),
.B2(n_223),
.Y(n_240)
);

AOI22xp33_ASAP7_75t_SL g257 ( 
.A1(n_241),
.A2(n_31),
.B1(n_24),
.B2(n_9),
.Y(n_257)
);

OAI22xp5_ASAP7_75t_SL g242 ( 
.A1(n_215),
.A2(n_21),
.B1(n_20),
.B2(n_48),
.Y(n_242)
);

XNOR2xp5_ASAP7_75t_L g244 ( 
.A(n_225),
.B(n_19),
.Y(n_244)
);

MAJIxp5_ASAP7_75t_L g250 ( 
.A(n_244),
.B(n_248),
.C(n_226),
.Y(n_250)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_220),
.Y(n_245)
);

CKINVDCx20_ASAP7_75t_R g262 ( 
.A(n_245),
.Y(n_262)
);

AOI21xp5_ASAP7_75t_L g249 ( 
.A1(n_246),
.A2(n_247),
.B(n_0),
.Y(n_249)
);

AND2x2_ASAP7_75t_L g247 ( 
.A(n_216),
.B(n_23),
.Y(n_247)
);

XNOR2xp5_ASAP7_75t_L g248 ( 
.A(n_213),
.B(n_15),
.Y(n_248)
);

CKINVDCx20_ASAP7_75t_R g271 ( 
.A(n_249),
.Y(n_271)
);

XOR2xp5_ASAP7_75t_L g267 ( 
.A(n_250),
.B(n_255),
.Y(n_267)
);

OA21x2_ASAP7_75t_L g251 ( 
.A1(n_241),
.A2(n_217),
.B(n_208),
.Y(n_251)
);

AOI22xp33_ASAP7_75t_SL g277 ( 
.A1(n_251),
.A2(n_18),
.B1(n_23),
.B2(n_12),
.Y(n_277)
);

OAI22xp5_ASAP7_75t_SL g252 ( 
.A1(n_238),
.A2(n_209),
.B1(n_229),
.B2(n_208),
.Y(n_252)
);

AOI22xp5_ASAP7_75t_L g274 ( 
.A1(n_252),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_274)
);

MAJIxp5_ASAP7_75t_L g253 ( 
.A(n_243),
.B(n_209),
.C(n_214),
.Y(n_253)
);

MAJIxp5_ASAP7_75t_L g270 ( 
.A(n_253),
.B(n_237),
.C(n_15),
.Y(n_270)
);

NAND2xp5_ASAP7_75t_SL g266 ( 
.A(n_254),
.B(n_258),
.Y(n_266)
);

XNOR2xp5_ASAP7_75t_SL g273 ( 
.A(n_257),
.B(n_24),
.Y(n_273)
);

INVxp67_ASAP7_75t_L g258 ( 
.A(n_247),
.Y(n_258)
);

AOI22xp5_ASAP7_75t_L g259 ( 
.A1(n_231),
.A2(n_8),
.B1(n_7),
.B2(n_6),
.Y(n_259)
);

NAND2xp5_ASAP7_75t_SL g268 ( 
.A(n_259),
.B(n_232),
.Y(n_268)
);

AOI21xp5_ASAP7_75t_L g264 ( 
.A1(n_262),
.A2(n_244),
.B(n_239),
.Y(n_264)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_264),
.Y(n_280)
);

CKINVDCx16_ASAP7_75t_R g265 ( 
.A(n_263),
.Y(n_265)
);

NAND2xp5_ASAP7_75t_L g286 ( 
.A(n_265),
.B(n_268),
.Y(n_286)
);

NAND2xp5_ASAP7_75t_SL g269 ( 
.A(n_260),
.B(n_248),
.Y(n_269)
);

NAND2xp5_ASAP7_75t_L g289 ( 
.A(n_269),
.B(n_270),
.Y(n_289)
);

AOI21xp5_ASAP7_75t_L g272 ( 
.A1(n_254),
.A2(n_6),
.B(n_2),
.Y(n_272)
);

OAI21xp5_ASAP7_75t_L g279 ( 
.A1(n_272),
.A2(n_251),
.B(n_2),
.Y(n_279)
);

MAJIxp5_ASAP7_75t_L g281 ( 
.A(n_273),
.B(n_256),
.C(n_12),
.Y(n_281)
);

NAND2xp5_ASAP7_75t_SL g287 ( 
.A(n_274),
.B(n_275),
.Y(n_287)
);

NOR2xp33_ASAP7_75t_SL g275 ( 
.A(n_253),
.B(n_15),
.Y(n_275)
);

NAND2xp5_ASAP7_75t_SL g276 ( 
.A(n_261),
.B(n_252),
.Y(n_276)
);

NOR2xp33_ASAP7_75t_L g282 ( 
.A(n_276),
.B(n_267),
.Y(n_282)
);

XOR2xp5_ASAP7_75t_SL g283 ( 
.A(n_277),
.B(n_18),
.Y(n_283)
);

AOI322xp5_ASAP7_75t_L g278 ( 
.A1(n_266),
.A2(n_258),
.A3(n_251),
.B1(n_250),
.B2(n_259),
.C1(n_256),
.C2(n_12),
.Y(n_278)
);

NAND2xp5_ASAP7_75t_L g296 ( 
.A(n_278),
.B(n_282),
.Y(n_296)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_279),
.Y(n_295)
);

XNOR2xp5_ASAP7_75t_SL g297 ( 
.A(n_281),
.B(n_283),
.Y(n_297)
);

MAJIxp5_ASAP7_75t_L g284 ( 
.A(n_267),
.B(n_22),
.C(n_12),
.Y(n_284)
);

OAI21xp5_ASAP7_75t_L g292 ( 
.A1(n_284),
.A2(n_285),
.B(n_288),
.Y(n_292)
);

MAJIxp5_ASAP7_75t_L g285 ( 
.A(n_270),
.B(n_271),
.C(n_273),
.Y(n_285)
);

NAND3xp33_ASAP7_75t_L g288 ( 
.A(n_277),
.B(n_1),
.C(n_2),
.Y(n_288)
);

AOI21x1_ASAP7_75t_L g290 ( 
.A1(n_286),
.A2(n_12),
.B(n_23),
.Y(n_290)
);

AOI21xp5_ASAP7_75t_L g302 ( 
.A1(n_290),
.A2(n_293),
.B(n_294),
.Y(n_302)
);

AOI21xp5_ASAP7_75t_L g291 ( 
.A1(n_280),
.A2(n_1),
.B(n_3),
.Y(n_291)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_291),
.Y(n_299)
);

NOR2xp67_ASAP7_75t_L g293 ( 
.A(n_283),
.B(n_23),
.Y(n_293)
);

NOR2x1_ASAP7_75t_L g294 ( 
.A(n_287),
.B(n_23),
.Y(n_294)
);

AOI21xp5_ASAP7_75t_L g298 ( 
.A1(n_289),
.A2(n_1),
.B(n_3),
.Y(n_298)
);

OAI21xp5_ASAP7_75t_L g301 ( 
.A1(n_298),
.A2(n_3),
.B(n_4),
.Y(n_301)
);

MAJIxp5_ASAP7_75t_L g300 ( 
.A(n_296),
.B(n_284),
.C(n_288),
.Y(n_300)
);

NAND2xp5_ASAP7_75t_SL g304 ( 
.A(n_300),
.B(n_297),
.Y(n_304)
);

MAJIxp5_ASAP7_75t_L g303 ( 
.A(n_301),
.B(n_295),
.C(n_292),
.Y(n_303)
);

AOI21xp5_ASAP7_75t_L g306 ( 
.A1(n_303),
.A2(n_304),
.B(n_305),
.Y(n_306)
);

OAI21xp5_ASAP7_75t_L g305 ( 
.A1(n_302),
.A2(n_18),
.B(n_22),
.Y(n_305)
);

AOI211xp5_ASAP7_75t_L g307 ( 
.A1(n_306),
.A2(n_299),
.B(n_18),
.C(n_5),
.Y(n_307)
);

OAI321xp33_ASAP7_75t_L g308 ( 
.A1(n_307),
.A2(n_4),
.A3(n_5),
.B1(n_18),
.B2(n_283),
.C(n_293),
.Y(n_308)
);

AOI21xp5_ASAP7_75t_L g309 ( 
.A1(n_308),
.A2(n_4),
.B(n_5),
.Y(n_309)
);

MAJIxp5_ASAP7_75t_L g310 ( 
.A(n_309),
.B(n_4),
.C(n_5),
.Y(n_310)
);

BUFx24_ASAP7_75t_SL g311 ( 
.A(n_310),
.Y(n_311)
);


endmodule