module fake_jpeg_7224_n_328 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_328);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_328;

wire n_253;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_7),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_12),
.Y(n_18)
);

BUFx5_ASAP7_75t_L g19 ( 
.A(n_1),
.Y(n_19)
);

INVx1_ASAP7_75t_SL g20 ( 
.A(n_16),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_3),
.Y(n_21)
);

BUFx12_ASAP7_75t_L g22 ( 
.A(n_12),
.Y(n_22)
);

BUFx12f_ASAP7_75t_L g23 ( 
.A(n_1),
.Y(n_23)
);

BUFx10_ASAP7_75t_L g24 ( 
.A(n_3),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_10),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_5),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_10),
.Y(n_27)
);

BUFx5_ASAP7_75t_L g28 ( 
.A(n_11),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_6),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_5),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_14),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_0),
.Y(n_32)
);

INVx3_ASAP7_75t_L g33 ( 
.A(n_13),
.Y(n_33)
);

BUFx12f_ASAP7_75t_L g34 ( 
.A(n_10),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_L g35 ( 
.A(n_20),
.B(n_34),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_SL g46 ( 
.A(n_35),
.B(n_44),
.Y(n_46)
);

INVx2_ASAP7_75t_L g36 ( 
.A(n_19),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_36),
.B(n_41),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_L g37 ( 
.A(n_23),
.B(n_0),
.Y(n_37)
);

NAND2xp5_ASAP7_75t_L g55 ( 
.A(n_37),
.B(n_23),
.Y(n_55)
);

INVx6_ASAP7_75t_L g38 ( 
.A(n_30),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g59 ( 
.A(n_38),
.Y(n_59)
);

INVx4_ASAP7_75t_L g39 ( 
.A(n_23),
.Y(n_39)
);

INVx4_ASAP7_75t_L g50 ( 
.A(n_39),
.Y(n_50)
);

BUFx24_ASAP7_75t_L g40 ( 
.A(n_19),
.Y(n_40)
);

BUFx10_ASAP7_75t_L g54 ( 
.A(n_40),
.Y(n_54)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_19),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_34),
.Y(n_42)
);

INVx3_ASAP7_75t_L g69 ( 
.A(n_42),
.Y(n_69)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_34),
.Y(n_43)
);

INVx3_ASAP7_75t_L g49 ( 
.A(n_43),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g44 ( 
.A(n_20),
.B(n_34),
.Y(n_44)
);

INVx2_ASAP7_75t_L g45 ( 
.A(n_42),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_45),
.B(n_51),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_SL g47 ( 
.A(n_37),
.B(n_25),
.Y(n_47)
);

NAND2xp5_ASAP7_75t_L g73 ( 
.A(n_47),
.B(n_61),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g51 ( 
.A(n_37),
.B(n_20),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_35),
.B(n_26),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_52),
.B(n_57),
.Y(n_83)
);

AOI22xp33_ASAP7_75t_L g53 ( 
.A1(n_38),
.A2(n_33),
.B1(n_18),
.B2(n_27),
.Y(n_53)
);

OAI22xp5_ASAP7_75t_L g78 ( 
.A1(n_53),
.A2(n_68),
.B1(n_29),
.B2(n_21),
.Y(n_78)
);

XNOR2xp5_ASAP7_75t_SL g80 ( 
.A(n_55),
.B(n_56),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_L g56 ( 
.A(n_35),
.B(n_23),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g57 ( 
.A(n_44),
.B(n_26),
.Y(n_57)
);

INVx5_ASAP7_75t_L g58 ( 
.A(n_42),
.Y(n_58)
);

INVx2_ASAP7_75t_L g91 ( 
.A(n_58),
.Y(n_91)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_42),
.Y(n_60)
);

INVxp67_ASAP7_75t_SL g95 ( 
.A(n_60),
.Y(n_95)
);

CKINVDCx16_ASAP7_75t_R g61 ( 
.A(n_44),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_39),
.B(n_26),
.Y(n_62)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_62),
.Y(n_90)
);

OAI22xp5_ASAP7_75t_L g63 ( 
.A1(n_38),
.A2(n_33),
.B1(n_28),
.B2(n_32),
.Y(n_63)
);

AOI22xp5_ASAP7_75t_L g72 ( 
.A1(n_63),
.A2(n_29),
.B1(n_18),
.B2(n_27),
.Y(n_72)
);

INVx2_ASAP7_75t_L g64 ( 
.A(n_42),
.Y(n_64)
);

INVx2_ASAP7_75t_SL g88 ( 
.A(n_64),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_39),
.B(n_25),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_L g76 ( 
.A(n_65),
.B(n_66),
.Y(n_76)
);

CKINVDCx16_ASAP7_75t_R g66 ( 
.A(n_40),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_39),
.B(n_25),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_L g94 ( 
.A(n_67),
.B(n_43),
.Y(n_94)
);

AOI22xp5_ASAP7_75t_L g68 ( 
.A1(n_38),
.A2(n_33),
.B1(n_28),
.B2(n_30),
.Y(n_68)
);

INVx5_ASAP7_75t_L g70 ( 
.A(n_43),
.Y(n_70)
);

AOI22xp33_ASAP7_75t_SL g87 ( 
.A1(n_70),
.A2(n_36),
.B1(n_40),
.B2(n_30),
.Y(n_87)
);

AND2x2_ASAP7_75t_L g71 ( 
.A(n_47),
.B(n_41),
.Y(n_71)
);

OAI21xp5_ASAP7_75t_SL g122 ( 
.A1(n_71),
.A2(n_77),
.B(n_34),
.Y(n_122)
);

OAI22xp33_ASAP7_75t_SL g103 ( 
.A1(n_72),
.A2(n_78),
.B1(n_87),
.B2(n_89),
.Y(n_103)
);

INVx3_ASAP7_75t_L g74 ( 
.A(n_45),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_74),
.B(n_92),
.Y(n_101)
);

AND2x2_ASAP7_75t_SL g75 ( 
.A(n_55),
.B(n_41),
.Y(n_75)
);

MAJIxp5_ASAP7_75t_L g96 ( 
.A(n_75),
.B(n_56),
.C(n_46),
.Y(n_96)
);

AND2x2_ASAP7_75t_L g77 ( 
.A(n_61),
.B(n_28),
.Y(n_77)
);

AOI22xp33_ASAP7_75t_L g79 ( 
.A1(n_51),
.A2(n_29),
.B1(n_18),
.B2(n_27),
.Y(n_79)
);

AOI22xp33_ASAP7_75t_L g102 ( 
.A1(n_79),
.A2(n_52),
.B1(n_21),
.B2(n_32),
.Y(n_102)
);

OA22x2_ASAP7_75t_L g82 ( 
.A1(n_59),
.A2(n_40),
.B1(n_43),
.B2(n_36),
.Y(n_82)
);

AOI22xp5_ASAP7_75t_L g116 ( 
.A1(n_82),
.A2(n_66),
.B1(n_70),
.B2(n_58),
.Y(n_116)
);

INVxp67_ASAP7_75t_L g84 ( 
.A(n_48),
.Y(n_84)
);

INVxp67_ASAP7_75t_L g111 ( 
.A(n_84),
.Y(n_111)
);

AOI22xp5_ASAP7_75t_SL g85 ( 
.A1(n_46),
.A2(n_31),
.B1(n_17),
.B2(n_21),
.Y(n_85)
);

INVxp67_ASAP7_75t_L g123 ( 
.A(n_85),
.Y(n_123)
);

BUFx3_ASAP7_75t_L g86 ( 
.A(n_54),
.Y(n_86)
);

CKINVDCx16_ASAP7_75t_R g105 ( 
.A(n_86),
.Y(n_105)
);

AOI22xp33_ASAP7_75t_SL g89 ( 
.A1(n_58),
.A2(n_17),
.B1(n_31),
.B2(n_32),
.Y(n_89)
);

INVx4_ASAP7_75t_L g92 ( 
.A(n_50),
.Y(n_92)
);

CKINVDCx16_ASAP7_75t_R g93 ( 
.A(n_62),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_93),
.B(n_94),
.Y(n_109)
);

XNOR2xp5_ASAP7_75t_L g128 ( 
.A(n_96),
.B(n_119),
.Y(n_128)
);

AO22x2_ASAP7_75t_SL g97 ( 
.A1(n_82),
.A2(n_59),
.B1(n_68),
.B2(n_63),
.Y(n_97)
);

OAI22xp5_ASAP7_75t_SL g141 ( 
.A1(n_97),
.A2(n_116),
.B1(n_118),
.B2(n_88),
.Y(n_141)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_82),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_SL g136 ( 
.A(n_98),
.B(n_100),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_SL g99 ( 
.A(n_71),
.B(n_57),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g130 ( 
.A(n_99),
.B(n_114),
.Y(n_130)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_82),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g132 ( 
.A(n_102),
.B(n_104),
.Y(n_132)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_82),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_SL g106 ( 
.A(n_83),
.B(n_67),
.Y(n_106)
);

NOR3xp33_ASAP7_75t_L g150 ( 
.A(n_106),
.B(n_77),
.C(n_90),
.Y(n_150)
);

CKINVDCx16_ASAP7_75t_R g107 ( 
.A(n_76),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_L g142 ( 
.A(n_107),
.B(n_108),
.Y(n_142)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_81),
.Y(n_108)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_81),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_L g144 ( 
.A(n_110),
.B(n_115),
.Y(n_144)
);

NOR2xp33_ASAP7_75t_L g112 ( 
.A(n_90),
.B(n_65),
.Y(n_112)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_112),
.Y(n_124)
);

OAI22xp33_ASAP7_75t_SL g113 ( 
.A1(n_93),
.A2(n_60),
.B1(n_64),
.B2(n_70),
.Y(n_113)
);

AOI22xp33_ASAP7_75t_L g138 ( 
.A1(n_113),
.A2(n_91),
.B1(n_88),
.B2(n_74),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_SL g114 ( 
.A(n_71),
.B(n_48),
.Y(n_114)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_94),
.Y(n_115)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_72),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_L g147 ( 
.A(n_117),
.B(n_121),
.Y(n_147)
);

AOI22xp5_ASAP7_75t_L g118 ( 
.A1(n_80),
.A2(n_69),
.B1(n_49),
.B2(n_50),
.Y(n_118)
);

XNOR2xp5_ASAP7_75t_L g119 ( 
.A(n_80),
.B(n_40),
.Y(n_119)
);

MAJIxp5_ASAP7_75t_L g120 ( 
.A(n_80),
.B(n_43),
.C(n_50),
.Y(n_120)
);

AND2x2_ASAP7_75t_L g134 ( 
.A(n_120),
.B(n_122),
.Y(n_134)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_83),
.Y(n_121)
);

CKINVDCx20_ASAP7_75t_R g125 ( 
.A(n_101),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_SL g172 ( 
.A(n_125),
.B(n_129),
.Y(n_172)
);

AOI22xp5_ASAP7_75t_L g126 ( 
.A1(n_97),
.A2(n_117),
.B1(n_98),
.B2(n_100),
.Y(n_126)
);

OAI22xp5_ASAP7_75t_SL g171 ( 
.A1(n_126),
.A2(n_151),
.B1(n_131),
.B2(n_148),
.Y(n_171)
);

XNOR2x1_ASAP7_75t_SL g127 ( 
.A(n_119),
.B(n_75),
.Y(n_127)
);

OAI21xp5_ASAP7_75t_L g160 ( 
.A1(n_127),
.A2(n_146),
.B(n_96),
.Y(n_160)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_101),
.Y(n_129)
);

INVx2_ASAP7_75t_SL g131 ( 
.A(n_97),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_L g152 ( 
.A(n_131),
.B(n_133),
.Y(n_152)
);

CKINVDCx16_ASAP7_75t_R g133 ( 
.A(n_112),
.Y(n_133)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_109),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_L g153 ( 
.A(n_135),
.B(n_138),
.Y(n_153)
);

A2O1A1Ixp33_ASAP7_75t_L g137 ( 
.A1(n_123),
.A2(n_73),
.B(n_71),
.C(n_75),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_L g158 ( 
.A(n_137),
.B(n_139),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_L g139 ( 
.A(n_114),
.B(n_75),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_L g140 ( 
.A(n_120),
.B(n_73),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_L g163 ( 
.A(n_140),
.B(n_143),
.Y(n_163)
);

NOR2xp33_ASAP7_75t_L g156 ( 
.A(n_141),
.B(n_148),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_L g143 ( 
.A(n_115),
.B(n_107),
.Y(n_143)
);

BUFx3_ASAP7_75t_L g145 ( 
.A(n_105),
.Y(n_145)
);

INVx13_ASAP7_75t_L g169 ( 
.A(n_145),
.Y(n_169)
);

AOI32xp33_ASAP7_75t_L g146 ( 
.A1(n_109),
.A2(n_76),
.A3(n_77),
.B1(n_85),
.B2(n_69),
.Y(n_146)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_118),
.Y(n_148)
);

BUFx12f_ASAP7_75t_L g149 ( 
.A(n_105),
.Y(n_149)
);

INVx4_ASAP7_75t_L g170 ( 
.A(n_149),
.Y(n_170)
);

NOR2xp33_ASAP7_75t_L g177 ( 
.A(n_150),
.B(n_22),
.Y(n_177)
);

AOI22xp5_ASAP7_75t_L g151 ( 
.A1(n_97),
.A2(n_78),
.B1(n_91),
.B2(n_77),
.Y(n_151)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_144),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_L g188 ( 
.A(n_154),
.B(n_162),
.Y(n_188)
);

AOI21xp5_ASAP7_75t_SL g155 ( 
.A1(n_135),
.A2(n_122),
.B(n_99),
.Y(n_155)
);

OAI21xp33_ASAP7_75t_SL g192 ( 
.A1(n_155),
.A2(n_159),
.B(n_177),
.Y(n_192)
);

HB1xp67_ASAP7_75t_L g157 ( 
.A(n_145),
.Y(n_157)
);

NOR2xp33_ASAP7_75t_L g200 ( 
.A(n_157),
.B(n_165),
.Y(n_200)
);

OAI22x1_ASAP7_75t_L g159 ( 
.A1(n_151),
.A2(n_103),
.B1(n_111),
.B2(n_108),
.Y(n_159)
);

XNOR2xp5_ASAP7_75t_SL g196 ( 
.A(n_160),
.B(n_128),
.Y(n_196)
);

BUFx6f_ASAP7_75t_L g161 ( 
.A(n_149),
.Y(n_161)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_161),
.Y(n_181)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_143),
.Y(n_162)
);

XOR2xp5_ASAP7_75t_L g164 ( 
.A(n_140),
.B(n_110),
.Y(n_164)
);

XOR2xp5_ASAP7_75t_L g198 ( 
.A(n_164),
.B(n_40),
.Y(n_198)
);

NAND3xp33_ASAP7_75t_L g165 ( 
.A(n_127),
.B(n_121),
.C(n_106),
.Y(n_165)
);

CKINVDCx20_ASAP7_75t_R g166 ( 
.A(n_149),
.Y(n_166)
);

NOR2xp33_ASAP7_75t_L g207 ( 
.A(n_166),
.B(n_173),
.Y(n_207)
);

OAI22xp5_ASAP7_75t_L g167 ( 
.A1(n_131),
.A2(n_104),
.B1(n_116),
.B2(n_102),
.Y(n_167)
);

OAI22xp5_ASAP7_75t_SL g206 ( 
.A1(n_167),
.A2(n_180),
.B1(n_153),
.B2(n_176),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_L g168 ( 
.A(n_139),
.B(n_23),
.Y(n_168)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_168),
.Y(n_195)
);

AOI22xp5_ASAP7_75t_L g182 ( 
.A1(n_171),
.A2(n_179),
.B1(n_180),
.B2(n_141),
.Y(n_182)
);

OR2x2_ASAP7_75t_L g173 ( 
.A(n_147),
.B(n_92),
.Y(n_173)
);

INVx2_ASAP7_75t_L g174 ( 
.A(n_149),
.Y(n_174)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_174),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_L g175 ( 
.A(n_130),
.B(n_23),
.Y(n_175)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_175),
.Y(n_186)
);

INVx1_ASAP7_75t_SL g176 ( 
.A(n_130),
.Y(n_176)
);

INVx1_ASAP7_75t_SL g193 ( 
.A(n_176),
.Y(n_193)
);

INVx2_ASAP7_75t_L g178 ( 
.A(n_129),
.Y(n_178)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_178),
.Y(n_189)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_142),
.Y(n_179)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_136),
.Y(n_180)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_182),
.Y(n_209)
);

AOI22xp5_ASAP7_75t_L g184 ( 
.A1(n_171),
.A2(n_132),
.B1(n_125),
.B2(n_126),
.Y(n_184)
);

OAI22xp5_ASAP7_75t_SL g218 ( 
.A1(n_184),
.A2(n_187),
.B1(n_191),
.B2(n_194),
.Y(n_218)
);

CKINVDCx20_ASAP7_75t_R g185 ( 
.A(n_172),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_SL g226 ( 
.A(n_185),
.B(n_190),
.Y(n_226)
);

AOI22xp5_ASAP7_75t_L g187 ( 
.A1(n_156),
.A2(n_124),
.B1(n_134),
.B2(n_137),
.Y(n_187)
);

INVxp67_ASAP7_75t_L g190 ( 
.A(n_152),
.Y(n_190)
);

AOI22xp5_ASAP7_75t_L g191 ( 
.A1(n_159),
.A2(n_124),
.B1(n_134),
.B2(n_92),
.Y(n_191)
);

AOI22xp5_ASAP7_75t_L g194 ( 
.A1(n_162),
.A2(n_134),
.B1(n_69),
.B2(n_128),
.Y(n_194)
);

XOR2xp5_ASAP7_75t_L g224 ( 
.A(n_196),
.B(n_202),
.Y(n_224)
);

CKINVDCx20_ASAP7_75t_R g197 ( 
.A(n_173),
.Y(n_197)
);

NOR2xp33_ASAP7_75t_SL g229 ( 
.A(n_197),
.B(n_205),
.Y(n_229)
);

MAJIxp5_ASAP7_75t_L g223 ( 
.A(n_198),
.B(n_199),
.C(n_201),
.Y(n_223)
);

XOR2xp5_ASAP7_75t_L g199 ( 
.A(n_160),
.B(n_40),
.Y(n_199)
);

XOR2xp5_ASAP7_75t_L g201 ( 
.A(n_164),
.B(n_95),
.Y(n_201)
);

XOR2xp5_ASAP7_75t_L g202 ( 
.A(n_163),
.B(n_95),
.Y(n_202)
);

AOI21xp5_ASAP7_75t_L g203 ( 
.A1(n_158),
.A2(n_86),
.B(n_54),
.Y(n_203)
);

OAI21xp5_ASAP7_75t_L g219 ( 
.A1(n_203),
.A2(n_166),
.B(n_154),
.Y(n_219)
);

XOR2xp5_ASAP7_75t_L g204 ( 
.A(n_163),
.B(n_54),
.Y(n_204)
);

XNOR2xp5_ASAP7_75t_L g211 ( 
.A(n_204),
.B(n_168),
.Y(n_211)
);

CKINVDCx20_ASAP7_75t_R g205 ( 
.A(n_169),
.Y(n_205)
);

AOI22xp5_ASAP7_75t_L g215 ( 
.A1(n_206),
.A2(n_155),
.B1(n_167),
.B2(n_179),
.Y(n_215)
);

NAND2xp5_ASAP7_75t_L g208 ( 
.A(n_193),
.B(n_175),
.Y(n_208)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_208),
.Y(n_241)
);

AOI22xp5_ASAP7_75t_SL g210 ( 
.A1(n_190),
.A2(n_192),
.B1(n_193),
.B2(n_186),
.Y(n_210)
);

OAI22xp5_ASAP7_75t_L g235 ( 
.A1(n_210),
.A2(n_215),
.B1(n_219),
.B2(n_203),
.Y(n_235)
);

MAJIxp5_ASAP7_75t_L g238 ( 
.A(n_211),
.B(n_228),
.C(n_231),
.Y(n_238)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_188),
.Y(n_212)
);

NAND2xp5_ASAP7_75t_L g234 ( 
.A(n_212),
.B(n_216),
.Y(n_234)
);

NAND2xp5_ASAP7_75t_L g213 ( 
.A(n_188),
.B(n_178),
.Y(n_213)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_213),
.Y(n_250)
);

NAND2xp5_ASAP7_75t_L g214 ( 
.A(n_206),
.B(n_158),
.Y(n_214)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_214),
.Y(n_252)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_207),
.Y(n_216)
);

NOR2xp33_ASAP7_75t_L g217 ( 
.A(n_181),
.B(n_174),
.Y(n_217)
);

NAND2xp5_ASAP7_75t_L g245 ( 
.A(n_217),
.B(n_220),
.Y(n_245)
);

CKINVDCx20_ASAP7_75t_R g220 ( 
.A(n_182),
.Y(n_220)
);

NAND2xp5_ASAP7_75t_L g221 ( 
.A(n_195),
.B(n_161),
.Y(n_221)
);

CKINVDCx20_ASAP7_75t_R g247 ( 
.A(n_221),
.Y(n_247)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_189),
.Y(n_222)
);

NOR2xp33_ASAP7_75t_L g233 ( 
.A(n_222),
.B(n_227),
.Y(n_233)
);

NAND2xp5_ASAP7_75t_L g225 ( 
.A(n_195),
.B(n_170),
.Y(n_225)
);

CKINVDCx16_ASAP7_75t_R g237 ( 
.A(n_225),
.Y(n_237)
);

NAND2xp5_ASAP7_75t_L g227 ( 
.A(n_202),
.B(n_170),
.Y(n_227)
);

XNOR2xp5_ASAP7_75t_L g228 ( 
.A(n_196),
.B(n_199),
.Y(n_228)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_191),
.Y(n_230)
);

NOR2xp33_ASAP7_75t_L g254 ( 
.A(n_230),
.B(n_232),
.Y(n_254)
);

XNOR2xp5_ASAP7_75t_L g231 ( 
.A(n_201),
.B(n_169),
.Y(n_231)
);

NAND2xp5_ASAP7_75t_L g232 ( 
.A(n_204),
.B(n_30),
.Y(n_232)
);

AOI21xp5_ASAP7_75t_L g256 ( 
.A1(n_235),
.A2(n_219),
.B(n_214),
.Y(n_256)
);

XNOR2xp5_ASAP7_75t_L g236 ( 
.A(n_231),
.B(n_194),
.Y(n_236)
);

XOR2xp5_ASAP7_75t_L g267 ( 
.A(n_236),
.B(n_240),
.Y(n_267)
);

AOI22xp5_ASAP7_75t_L g239 ( 
.A1(n_218),
.A2(n_200),
.B1(n_184),
.B2(n_183),
.Y(n_239)
);

AOI22xp33_ASAP7_75t_L g270 ( 
.A1(n_239),
.A2(n_244),
.B1(n_24),
.B2(n_22),
.Y(n_270)
);

XNOR2xp5_ASAP7_75t_L g240 ( 
.A(n_211),
.B(n_187),
.Y(n_240)
);

XNOR2xp5_ASAP7_75t_L g242 ( 
.A(n_223),
.B(n_198),
.Y(n_242)
);

XOR2xp5_ASAP7_75t_L g271 ( 
.A(n_242),
.B(n_246),
.Y(n_271)
);

AOI22xp5_ASAP7_75t_L g243 ( 
.A1(n_218),
.A2(n_49),
.B1(n_86),
.B2(n_88),
.Y(n_243)
);

AOI22xp5_ASAP7_75t_L g269 ( 
.A1(n_243),
.A2(n_250),
.B1(n_254),
.B2(n_253),
.Y(n_269)
);

AOI22xp5_ASAP7_75t_L g244 ( 
.A1(n_209),
.A2(n_34),
.B1(n_24),
.B2(n_54),
.Y(n_244)
);

XOR2xp5_ASAP7_75t_L g246 ( 
.A(n_224),
.B(n_54),
.Y(n_246)
);

XNOR2xp5_ASAP7_75t_L g248 ( 
.A(n_223),
.B(n_24),
.Y(n_248)
);

MAJIxp5_ASAP7_75t_L g260 ( 
.A(n_248),
.B(n_249),
.C(n_251),
.Y(n_260)
);

MAJIxp5_ASAP7_75t_L g249 ( 
.A(n_224),
.B(n_24),
.C(n_22),
.Y(n_249)
);

XOR2xp5_ASAP7_75t_L g251 ( 
.A(n_228),
.B(n_24),
.Y(n_251)
);

XOR2xp5_ASAP7_75t_L g253 ( 
.A(n_227),
.B(n_24),
.Y(n_253)
);

XNOR2xp5_ASAP7_75t_L g257 ( 
.A(n_253),
.B(n_213),
.Y(n_257)
);

NOR2xp33_ASAP7_75t_SL g255 ( 
.A(n_234),
.B(n_226),
.Y(n_255)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_255),
.Y(n_280)
);

OAI21xp5_ASAP7_75t_SL g275 ( 
.A1(n_256),
.A2(n_265),
.B(n_246),
.Y(n_275)
);

XNOR2xp5_ASAP7_75t_L g283 ( 
.A(n_257),
.B(n_269),
.Y(n_283)
);

NOR2xp33_ASAP7_75t_L g258 ( 
.A(n_252),
.B(n_229),
.Y(n_258)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_258),
.Y(n_284)
);

HB1xp67_ASAP7_75t_L g259 ( 
.A(n_237),
.Y(n_259)
);

NOR2xp33_ASAP7_75t_L g274 ( 
.A(n_259),
.B(n_268),
.Y(n_274)
);

XNOR2xp5_ASAP7_75t_L g261 ( 
.A(n_236),
.B(n_215),
.Y(n_261)
);

MAJIxp5_ASAP7_75t_L g273 ( 
.A(n_261),
.B(n_238),
.C(n_249),
.Y(n_273)
);

XNOR2xp5_ASAP7_75t_SL g262 ( 
.A(n_240),
.B(n_232),
.Y(n_262)
);

MAJx2_ASAP7_75t_L g281 ( 
.A(n_262),
.B(n_266),
.C(n_22),
.Y(n_281)
);

NOR2xp33_ASAP7_75t_SL g263 ( 
.A(n_233),
.B(n_210),
.Y(n_263)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_263),
.Y(n_286)
);

NOR2xp33_ASAP7_75t_L g264 ( 
.A(n_241),
.B(n_208),
.Y(n_264)
);

CKINVDCx14_ASAP7_75t_R g276 ( 
.A(n_264),
.Y(n_276)
);

AOI21xp5_ASAP7_75t_L g265 ( 
.A1(n_245),
.A2(n_221),
.B(n_225),
.Y(n_265)
);

XNOR2xp5_ASAP7_75t_SL g266 ( 
.A(n_242),
.B(n_248),
.Y(n_266)
);

NOR2xp33_ASAP7_75t_L g268 ( 
.A(n_247),
.B(n_22),
.Y(n_268)
);

HB1xp67_ASAP7_75t_L g279 ( 
.A(n_270),
.Y(n_279)
);

OAI21xp5_ASAP7_75t_L g272 ( 
.A1(n_243),
.A2(n_8),
.B(n_16),
.Y(n_272)
);

AOI21xp5_ASAP7_75t_L g285 ( 
.A1(n_272),
.A2(n_22),
.B(n_7),
.Y(n_285)
);

XNOR2xp5_ASAP7_75t_L g294 ( 
.A(n_273),
.B(n_6),
.Y(n_294)
);

AOI21xp5_ASAP7_75t_L g295 ( 
.A1(n_275),
.A2(n_287),
.B(n_15),
.Y(n_295)
);

AOI21xp5_ASAP7_75t_SL g277 ( 
.A1(n_272),
.A2(n_238),
.B(n_251),
.Y(n_277)
);

AOI21xp5_ASAP7_75t_SL g292 ( 
.A1(n_277),
.A2(n_260),
.B(n_271),
.Y(n_292)
);

MAJIxp5_ASAP7_75t_L g278 ( 
.A(n_267),
.B(n_8),
.C(n_16),
.Y(n_278)
);

MAJIxp5_ASAP7_75t_L g289 ( 
.A(n_278),
.B(n_282),
.C(n_269),
.Y(n_289)
);

AOI22xp5_ASAP7_75t_SL g299 ( 
.A1(n_281),
.A2(n_15),
.B1(n_12),
.B2(n_11),
.Y(n_299)
);

MAJIxp5_ASAP7_75t_L g282 ( 
.A(n_267),
.B(n_8),
.C(n_15),
.Y(n_282)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_285),
.Y(n_291)
);

OAI21xp5_ASAP7_75t_L g287 ( 
.A1(n_260),
.A2(n_7),
.B(n_14),
.Y(n_287)
);

AOI22xp5_ASAP7_75t_L g288 ( 
.A1(n_276),
.A2(n_262),
.B1(n_261),
.B2(n_266),
.Y(n_288)
);

OAI22xp5_ASAP7_75t_SL g305 ( 
.A1(n_288),
.A2(n_297),
.B1(n_299),
.B2(n_1),
.Y(n_305)
);

NAND2xp5_ASAP7_75t_L g301 ( 
.A(n_289),
.B(n_290),
.Y(n_301)
);

NAND2xp5_ASAP7_75t_SL g290 ( 
.A(n_280),
.B(n_257),
.Y(n_290)
);

AO21x1_ASAP7_75t_SL g304 ( 
.A1(n_292),
.A2(n_298),
.B(n_0),
.Y(n_304)
);

OAI22xp5_ASAP7_75t_SL g293 ( 
.A1(n_286),
.A2(n_271),
.B1(n_9),
.B2(n_11),
.Y(n_293)
);

INVxp67_ASAP7_75t_L g306 ( 
.A(n_293),
.Y(n_306)
);

XNOR2xp5_ASAP7_75t_L g308 ( 
.A(n_294),
.B(n_295),
.Y(n_308)
);

NOR2xp33_ASAP7_75t_L g296 ( 
.A(n_274),
.B(n_6),
.Y(n_296)
);

AOI21xp5_ASAP7_75t_L g307 ( 
.A1(n_296),
.A2(n_300),
.B(n_2),
.Y(n_307)
);

AOI22xp5_ASAP7_75t_L g297 ( 
.A1(n_284),
.A2(n_9),
.B1(n_14),
.B2(n_13),
.Y(n_297)
);

OAI21x1_ASAP7_75t_L g298 ( 
.A1(n_277),
.A2(n_5),
.B(n_13),
.Y(n_298)
);

MAJIxp5_ASAP7_75t_L g300 ( 
.A(n_273),
.B(n_0),
.C(n_1),
.Y(n_300)
);

AOI322xp5_ASAP7_75t_L g302 ( 
.A1(n_291),
.A2(n_283),
.A3(n_279),
.B1(n_281),
.B2(n_282),
.C1(n_278),
.C2(n_9),
.Y(n_302)
);

OR2x2_ASAP7_75t_L g311 ( 
.A(n_302),
.B(n_304),
.Y(n_311)
);

XOR2xp5_ASAP7_75t_L g303 ( 
.A(n_292),
.B(n_283),
.Y(n_303)
);

MAJIxp5_ASAP7_75t_L g315 ( 
.A(n_303),
.B(n_2),
.C(n_3),
.Y(n_315)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_305),
.Y(n_312)
);

NAND2xp5_ASAP7_75t_L g316 ( 
.A(n_307),
.B(n_309),
.Y(n_316)
);

XNOR2xp5_ASAP7_75t_L g309 ( 
.A(n_294),
.B(n_300),
.Y(n_309)
);

OAI22xp5_ASAP7_75t_SL g310 ( 
.A1(n_289),
.A2(n_2),
.B1(n_3),
.B2(n_4),
.Y(n_310)
);

NOR2xp33_ASAP7_75t_L g314 ( 
.A(n_310),
.B(n_2),
.Y(n_314)
);

NOR2xp33_ASAP7_75t_SL g313 ( 
.A(n_304),
.B(n_299),
.Y(n_313)
);

OAI21xp5_ASAP7_75t_L g321 ( 
.A1(n_313),
.A2(n_315),
.B(n_317),
.Y(n_321)
);

NOR2xp33_ASAP7_75t_SL g320 ( 
.A(n_314),
.B(n_4),
.Y(n_320)
);

MAJIxp5_ASAP7_75t_L g317 ( 
.A(n_301),
.B(n_4),
.C(n_303),
.Y(n_317)
);

AOI21xp5_ASAP7_75t_SL g318 ( 
.A1(n_306),
.A2(n_4),
.B(n_308),
.Y(n_318)
);

OAI21xp5_ASAP7_75t_SL g322 ( 
.A1(n_318),
.A2(n_313),
.B(n_312),
.Y(n_322)
);

NOR2xp67_ASAP7_75t_L g319 ( 
.A(n_311),
.B(n_306),
.Y(n_319)
);

OAI21xp5_ASAP7_75t_L g324 ( 
.A1(n_319),
.A2(n_320),
.B(n_323),
.Y(n_324)
);

INVxp67_ASAP7_75t_L g325 ( 
.A(n_322),
.Y(n_325)
);

INVxp67_ASAP7_75t_L g323 ( 
.A(n_316),
.Y(n_323)
);

NAND2xp5_ASAP7_75t_L g326 ( 
.A(n_325),
.B(n_321),
.Y(n_326)
);

BUFx24_ASAP7_75t_SL g327 ( 
.A(n_326),
.Y(n_327)
);

XOR2xp5_ASAP7_75t_L g328 ( 
.A(n_327),
.B(n_324),
.Y(n_328)
);


endmodule