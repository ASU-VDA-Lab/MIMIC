module real_jpeg_20227_n_16 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_3, n_10, n_9, n_16);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_16;

wire n_108;
wire n_54;
wire n_37;
wire n_168;
wire n_73;
wire n_35;
wire n_38;
wire n_29;
wire n_91;
wire n_49;
wire n_201;
wire n_114;
wire n_68;
wire n_146;
wire n_78;
wire n_83;
wire n_166;
wire n_176;
wire n_104;
wire n_153;
wire n_194;
wire n_161;
wire n_64;
wire n_177;
wire n_47;
wire n_131;
wire n_163;
wire n_22;
wire n_174;
wire n_87;
wire n_197;
wire n_40;
wire n_173;
wire n_105;
wire n_115;
wire n_98;
wire n_27;
wire n_56;
wire n_184;
wire n_48;
wire n_164;
wire n_200;
wire n_140;
wire n_126;
wire n_113;
wire n_120;
wire n_155;
wire n_199;
wire n_93;
wire n_141;
wire n_95;
wire n_65;
wire n_33;
wire n_139;
wire n_188;
wire n_142;
wire n_175;
wire n_76;
wire n_178;
wire n_67;
wire n_79;
wire n_107;
wire n_156;
wire n_147;
wire n_189;
wire n_170;
wire n_66;
wire n_136;
wire n_28;
wire n_44;
wire n_62;
wire n_162;
wire n_121;
wire n_106;
wire n_160;
wire n_172;
wire n_45;
wire n_112;
wire n_42;
wire n_18;
wire n_145;
wire n_77;
wire n_109;
wire n_39;
wire n_122;
wire n_94;
wire n_26;
wire n_19;
wire n_148;
wire n_118;
wire n_17;
wire n_123;
wire n_116;
wire n_21;
wire n_50;
wire n_143;
wire n_196;
wire n_69;
wire n_186;
wire n_31;
wire n_137;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_165;
wire n_134;
wire n_72;
wire n_159;
wire n_171;
wire n_151;
wire n_183;
wire n_198;
wire n_192;
wire n_100;
wire n_23;
wire n_51;
wire n_71;
wire n_90;
wire n_61;
wire n_195;
wire n_110;
wire n_117;
wire n_99;
wire n_193;
wire n_86;
wire n_150;
wire n_41;
wire n_74;
wire n_80;
wire n_32;
wire n_20;
wire n_70;
wire n_30;
wire n_158;
wire n_149;
wire n_144;
wire n_130;
wire n_103;
wire n_43;
wire n_57;
wire n_157;
wire n_84;
wire n_82;
wire n_111;
wire n_132;
wire n_185;
wire n_125;
wire n_55;
wire n_180;
wire n_58;
wire n_52;
wire n_191;
wire n_63;
wire n_124;
wire n_24;
wire n_92;
wire n_75;
wire n_97;
wire n_187;
wire n_34;
wire n_190;
wire n_60;
wire n_46;
wire n_88;
wire n_169;
wire n_59;
wire n_167;
wire n_202;
wire n_128;
wire n_179;
wire n_133;
wire n_138;
wire n_25;
wire n_53;
wire n_127;
wire n_119;
wire n_36;
wire n_81;
wire n_102;
wire n_85;
wire n_181;
wire n_101;
wire n_182;
wire n_96;
wire n_89;

OAI22xp5_ASAP7_75t_SL g53 ( 
.A1(n_0),
.A2(n_40),
.B1(n_41),
.B2(n_54),
.Y(n_53)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_0),
.Y(n_54)
);

AOI22xp5_ASAP7_75t_L g100 ( 
.A1(n_0),
.A2(n_54),
.B1(n_62),
.B2(n_63),
.Y(n_100)
);

OAI22xp5_ASAP7_75t_SL g165 ( 
.A1(n_0),
.A2(n_10),
.B1(n_28),
.B2(n_54),
.Y(n_165)
);

AOI22xp5_ASAP7_75t_SL g39 ( 
.A1(n_1),
.A2(n_40),
.B1(n_41),
.B2(n_42),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_1),
.Y(n_42)
);

AOI22xp33_ASAP7_75t_SL g87 ( 
.A1(n_1),
.A2(n_10),
.B1(n_28),
.B2(n_42),
.Y(n_87)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_2),
.Y(n_63)
);

CKINVDCx20_ASAP7_75t_R g74 ( 
.A(n_3),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_L g114 ( 
.A(n_3),
.B(n_78),
.Y(n_114)
);

AOI21xp33_ASAP7_75t_L g137 ( 
.A1(n_3),
.A2(n_10),
.B(n_14),
.Y(n_137)
);

AOI22xp33_ASAP7_75t_SL g140 ( 
.A1(n_3),
.A2(n_40),
.B1(n_41),
.B2(n_74),
.Y(n_140)
);

OAI22xp5_ASAP7_75t_L g148 ( 
.A1(n_3),
.A2(n_26),
.B1(n_33),
.B2(n_146),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_L g158 ( 
.A(n_3),
.B(n_118),
.Y(n_158)
);

NOR2xp33_ASAP7_75t_L g173 ( 
.A(n_3),
.B(n_62),
.Y(n_173)
);

AOI21xp33_ASAP7_75t_L g177 ( 
.A1(n_3),
.A2(n_62),
.B(n_173),
.Y(n_177)
);

AOI22xp33_ASAP7_75t_L g66 ( 
.A1(n_4),
.A2(n_62),
.B1(n_63),
.B2(n_67),
.Y(n_66)
);

CKINVDCx20_ASAP7_75t_R g67 ( 
.A(n_4),
.Y(n_67)
);

AOI22xp5_ASAP7_75t_SL g93 ( 
.A1(n_4),
.A2(n_67),
.B1(n_72),
.B2(n_81),
.Y(n_93)
);

AOI22xp33_ASAP7_75t_SL g130 ( 
.A1(n_4),
.A2(n_10),
.B1(n_28),
.B2(n_67),
.Y(n_130)
);

AOI22xp33_ASAP7_75t_SL g161 ( 
.A1(n_4),
.A2(n_40),
.B1(n_41),
.B2(n_67),
.Y(n_161)
);

INVx13_ASAP7_75t_L g76 ( 
.A(n_5),
.Y(n_76)
);

OAI22xp5_ASAP7_75t_L g78 ( 
.A1(n_5),
.A2(n_62),
.B1(n_63),
.B2(n_76),
.Y(n_78)
);

BUFx16f_ASAP7_75t_L g73 ( 
.A(n_6),
.Y(n_73)
);

OAI22xp5_ASAP7_75t_SL g79 ( 
.A1(n_7),
.A2(n_72),
.B1(n_80),
.B2(n_81),
.Y(n_79)
);

CKINVDCx20_ASAP7_75t_R g80 ( 
.A(n_7),
.Y(n_80)
);

AOI22xp33_ASAP7_75t_SL g117 ( 
.A1(n_7),
.A2(n_62),
.B1(n_63),
.B2(n_80),
.Y(n_117)
);

AOI22xp5_ASAP7_75t_SL g141 ( 
.A1(n_7),
.A2(n_40),
.B1(n_41),
.B2(n_80),
.Y(n_141)
);

AOI22xp5_ASAP7_75t_L g146 ( 
.A1(n_7),
.A2(n_10),
.B1(n_28),
.B2(n_80),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_L g27 ( 
.A(n_8),
.B(n_28),
.Y(n_27)
);

INVx8_ASAP7_75t_L g33 ( 
.A(n_8),
.Y(n_33)
);

INVx6_ASAP7_75t_L g111 ( 
.A(n_8),
.Y(n_111)
);

AOI22xp33_ASAP7_75t_SL g68 ( 
.A1(n_9),
.A2(n_62),
.B1(n_63),
.B2(n_69),
.Y(n_68)
);

CKINVDCx20_ASAP7_75t_R g69 ( 
.A(n_9),
.Y(n_69)
);

AOI22xp33_ASAP7_75t_SL g133 ( 
.A1(n_9),
.A2(n_10),
.B1(n_28),
.B2(n_69),
.Y(n_133)
);

AOI22xp33_ASAP7_75t_SL g180 ( 
.A1(n_9),
.A2(n_40),
.B1(n_41),
.B2(n_69),
.Y(n_180)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_10),
.Y(n_28)
);

AOI22xp33_ASAP7_75t_SL g29 ( 
.A1(n_10),
.A2(n_13),
.B1(n_28),
.B2(n_30),
.Y(n_29)
);

AOI22xp33_ASAP7_75t_L g34 ( 
.A1(n_10),
.A2(n_11),
.B1(n_28),
.B2(n_35),
.Y(n_34)
);

AOI22xp5_ASAP7_75t_SL g37 ( 
.A1(n_10),
.A2(n_14),
.B1(n_28),
.B2(n_38),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_11),
.Y(n_35)
);

OAI22xp33_ASAP7_75t_SL g44 ( 
.A1(n_11),
.A2(n_35),
.B1(n_40),
.B2(n_41),
.Y(n_44)
);

INVx13_ASAP7_75t_L g61 ( 
.A(n_12),
.Y(n_61)
);

CKINVDCx14_ASAP7_75t_R g30 ( 
.A(n_13),
.Y(n_30)
);

INVx11_ASAP7_75t_L g38 ( 
.A(n_14),
.Y(n_38)
);

A2O1A1Ixp33_ASAP7_75t_L g46 ( 
.A1(n_14),
.A2(n_37),
.B(n_40),
.C(n_47),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g47 ( 
.A(n_14),
.B(n_40),
.Y(n_47)
);

INVx11_ASAP7_75t_SL g40 ( 
.A(n_15),
.Y(n_40)
);

XNOR2xp5_ASAP7_75t_L g16 ( 
.A(n_17),
.B(n_122),
.Y(n_16)
);

NAND2xp5_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_120),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_19),
.Y(n_18)
);

AND2x2_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_102),
.Y(n_19)
);

NOR2xp33_ASAP7_75t_L g121 ( 
.A(n_20),
.B(n_102),
.Y(n_121)
);

OAI22xp5_ASAP7_75t_SL g20 ( 
.A1(n_21),
.A2(n_22),
.B1(n_82),
.B2(n_101),
.Y(n_20)
);

CKINVDCx14_ASAP7_75t_R g21 ( 
.A(n_22),
.Y(n_21)
);

XNOR2xp5_ASAP7_75t_SL g22 ( 
.A(n_23),
.B(n_49),
.Y(n_22)
);

OAI22xp5_ASAP7_75t_L g23 ( 
.A1(n_24),
.A2(n_25),
.B1(n_36),
.B2(n_48),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_25),
.Y(n_24)
);

OAI21xp5_ASAP7_75t_L g25 ( 
.A1(n_26),
.A2(n_29),
.B(n_31),
.Y(n_25)
);

OAI22xp5_ASAP7_75t_SL g86 ( 
.A1(n_26),
.A2(n_29),
.B1(n_33),
.B2(n_87),
.Y(n_86)
);

OAI22xp5_ASAP7_75t_SL g145 ( 
.A1(n_26),
.A2(n_111),
.B1(n_130),
.B2(n_146),
.Y(n_145)
);

OAI21xp5_ASAP7_75t_L g162 ( 
.A1(n_26),
.A2(n_133),
.B(n_163),
.Y(n_162)
);

CKINVDCx16_ASAP7_75t_R g26 ( 
.A(n_27),
.Y(n_26)
);

NAND2xp5_ASAP7_75t_SL g112 ( 
.A(n_27),
.B(n_113),
.Y(n_112)
);

AOI22xp5_ASAP7_75t_L g128 ( 
.A1(n_27),
.A2(n_129),
.B1(n_131),
.B2(n_132),
.Y(n_128)
);

AOI21xp5_ASAP7_75t_L g171 ( 
.A1(n_27),
.A2(n_32),
.B(n_165),
.Y(n_171)
);

NOR2xp33_ASAP7_75t_L g149 ( 
.A(n_28),
.B(n_150),
.Y(n_149)
);

INVxp67_ASAP7_75t_L g31 ( 
.A(n_32),
.Y(n_31)
);

NOR2xp33_ASAP7_75t_L g32 ( 
.A(n_33),
.B(n_34),
.Y(n_32)
);

INVx2_ASAP7_75t_L g131 ( 
.A(n_33),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_L g150 ( 
.A(n_33),
.B(n_74),
.Y(n_150)
);

CKINVDCx16_ASAP7_75t_R g113 ( 
.A(n_34),
.Y(n_113)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_36),
.Y(n_48)
);

OAI21xp5_ASAP7_75t_L g36 ( 
.A1(n_37),
.A2(n_39),
.B(n_43),
.Y(n_36)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_37),
.Y(n_56)
);

OAI22xp5_ASAP7_75t_SL g139 ( 
.A1(n_37),
.A2(n_46),
.B1(n_140),
.B2(n_141),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_L g144 ( 
.A(n_37),
.B(n_74),
.Y(n_144)
);

OAI22xp5_ASAP7_75t_SL g160 ( 
.A1(n_37),
.A2(n_46),
.B1(n_141),
.B2(n_161),
.Y(n_160)
);

OAI22xp5_ASAP7_75t_SL g179 ( 
.A1(n_37),
.A2(n_46),
.B1(n_161),
.B2(n_180),
.Y(n_179)
);

A2O1A1Ixp33_ASAP7_75t_L g136 ( 
.A1(n_38),
.A2(n_41),
.B(n_74),
.C(n_137),
.Y(n_136)
);

INVx11_ASAP7_75t_L g41 ( 
.A(n_40),
.Y(n_41)
);

AOI22xp5_ASAP7_75t_L g65 ( 
.A1(n_40),
.A2(n_41),
.B1(n_60),
.B2(n_61),
.Y(n_65)
);

AOI32xp33_ASAP7_75t_L g172 ( 
.A1(n_40),
.A2(n_61),
.A3(n_63),
.B1(n_173),
.B2(n_174),
.Y(n_172)
);

NAND2xp33_ASAP7_75t_SL g174 ( 
.A(n_41),
.B(n_60),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_L g43 ( 
.A(n_44),
.B(n_45),
.Y(n_43)
);

NAND2xp5_ASAP7_75t_SL g55 ( 
.A(n_44),
.B(n_56),
.Y(n_55)
);

INVxp67_ASAP7_75t_L g45 ( 
.A(n_46),
.Y(n_45)
);

OAI21xp5_ASAP7_75t_SL g51 ( 
.A1(n_46),
.A2(n_52),
.B(n_55),
.Y(n_51)
);

OAI21xp5_ASAP7_75t_SL g194 ( 
.A1(n_46),
.A2(n_180),
.B(n_195),
.Y(n_194)
);

MAJIxp5_ASAP7_75t_L g49 ( 
.A(n_50),
.B(n_57),
.C(n_70),
.Y(n_49)
);

AOI22xp5_ASAP7_75t_L g104 ( 
.A1(n_50),
.A2(n_51),
.B1(n_57),
.B2(n_58),
.Y(n_104)
);

CKINVDCx16_ASAP7_75t_R g50 ( 
.A(n_51),
.Y(n_50)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_53),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_SL g195 ( 
.A(n_53),
.B(n_56),
.Y(n_195)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_58),
.Y(n_57)
);

OAI22xp5_ASAP7_75t_SL g58 ( 
.A1(n_59),
.A2(n_65),
.B1(n_66),
.B2(n_68),
.Y(n_58)
);

CKINVDCx14_ASAP7_75t_R g97 ( 
.A(n_59),
.Y(n_97)
);

OAI22xp5_ASAP7_75t_SL g176 ( 
.A1(n_59),
.A2(n_65),
.B1(n_117),
.B2(n_177),
.Y(n_176)
);

A2O1A1Ixp33_ASAP7_75t_L g59 ( 
.A1(n_60),
.A2(n_62),
.B(n_64),
.C(n_65),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_60),
.B(n_62),
.Y(n_64)
);

INVx11_ASAP7_75t_L g60 ( 
.A(n_61),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_62),
.B(n_76),
.Y(n_85)
);

INVx8_ASAP7_75t_L g62 ( 
.A(n_63),
.Y(n_62)
);

OAI22xp5_ASAP7_75t_SL g84 ( 
.A1(n_63),
.A2(n_71),
.B1(n_77),
.B2(n_85),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_65),
.B(n_100),
.Y(n_99)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_65),
.Y(n_118)
);

CKINVDCx20_ASAP7_75t_R g119 ( 
.A(n_66),
.Y(n_119)
);

CKINVDCx20_ASAP7_75t_R g98 ( 
.A(n_68),
.Y(n_98)
);

XNOR2xp5_ASAP7_75t_SL g103 ( 
.A(n_70),
.B(n_104),
.Y(n_103)
);

AOI22xp5_ASAP7_75t_L g70 ( 
.A1(n_71),
.A2(n_75),
.B1(n_78),
.B2(n_79),
.Y(n_70)
);

HAxp5_ASAP7_75t_SL g71 ( 
.A(n_72),
.B(n_74),
.CON(n_71),
.SN(n_71)
);

O2A1O1Ixp33_ASAP7_75t_L g75 ( 
.A1(n_72),
.A2(n_76),
.B(n_77),
.C(n_78),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_L g77 ( 
.A(n_72),
.B(n_76),
.Y(n_77)
);

CKINVDCx20_ASAP7_75t_R g81 ( 
.A(n_72),
.Y(n_81)
);

BUFx2_ASAP7_75t_L g72 ( 
.A(n_73),
.Y(n_72)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_75),
.Y(n_91)
);

CKINVDCx20_ASAP7_75t_R g94 ( 
.A(n_78),
.Y(n_94)
);

CKINVDCx20_ASAP7_75t_R g92 ( 
.A(n_79),
.Y(n_92)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_82),
.Y(n_101)
);

XOR2xp5_ASAP7_75t_L g82 ( 
.A(n_83),
.B(n_88),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_L g83 ( 
.A(n_84),
.B(n_86),
.Y(n_83)
);

XOR2xp5_ASAP7_75t_L g106 ( 
.A(n_84),
.B(n_86),
.Y(n_106)
);

OAI21xp5_ASAP7_75t_L g110 ( 
.A1(n_87),
.A2(n_111),
.B(n_112),
.Y(n_110)
);

OAI22xp5_ASAP7_75t_SL g88 ( 
.A1(n_89),
.A2(n_90),
.B1(n_95),
.B2(n_96),
.Y(n_88)
);

CKINVDCx14_ASAP7_75t_R g89 ( 
.A(n_90),
.Y(n_89)
);

OAI22xp5_ASAP7_75t_SL g90 ( 
.A1(n_91),
.A2(n_92),
.B1(n_93),
.B2(n_94),
.Y(n_90)
);

CKINVDCx16_ASAP7_75t_R g95 ( 
.A(n_96),
.Y(n_95)
);

AOI21xp5_ASAP7_75t_L g96 ( 
.A1(n_97),
.A2(n_98),
.B(n_99),
.Y(n_96)
);

AOI22xp5_ASAP7_75t_L g115 ( 
.A1(n_97),
.A2(n_116),
.B1(n_118),
.B2(n_119),
.Y(n_115)
);

MAJIxp5_ASAP7_75t_L g102 ( 
.A(n_103),
.B(n_105),
.C(n_107),
.Y(n_102)
);

XOR2xp5_ASAP7_75t_L g200 ( 
.A(n_103),
.B(n_201),
.Y(n_200)
);

OAI22xp5_ASAP7_75t_L g201 ( 
.A1(n_105),
.A2(n_106),
.B1(n_107),
.B2(n_108),
.Y(n_201)
);

CKINVDCx20_ASAP7_75t_R g105 ( 
.A(n_106),
.Y(n_105)
);

CKINVDCx16_ASAP7_75t_R g107 ( 
.A(n_108),
.Y(n_107)
);

MAJIxp5_ASAP7_75t_L g108 ( 
.A(n_109),
.B(n_114),
.C(n_115),
.Y(n_108)
);

AOI22xp5_ASAP7_75t_L g190 ( 
.A1(n_109),
.A2(n_110),
.B1(n_114),
.B2(n_191),
.Y(n_190)
);

CKINVDCx20_ASAP7_75t_R g109 ( 
.A(n_110),
.Y(n_109)
);

INVx5_ASAP7_75t_L g164 ( 
.A(n_111),
.Y(n_164)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_114),
.Y(n_191)
);

XNOR2xp5_ASAP7_75t_SL g189 ( 
.A(n_115),
.B(n_190),
.Y(n_189)
);

CKINVDCx16_ASAP7_75t_R g116 ( 
.A(n_117),
.Y(n_116)
);

INVxp67_ASAP7_75t_L g120 ( 
.A(n_121),
.Y(n_120)
);

AOI21xp5_ASAP7_75t_L g122 ( 
.A1(n_123),
.A2(n_198),
.B(n_202),
.Y(n_122)
);

OAI21xp5_ASAP7_75t_SL g123 ( 
.A1(n_124),
.A2(n_185),
.B(n_197),
.Y(n_123)
);

AOI21xp5_ASAP7_75t_L g124 ( 
.A1(n_125),
.A2(n_167),
.B(n_184),
.Y(n_124)
);

OAI21xp5_ASAP7_75t_SL g125 ( 
.A1(n_126),
.A2(n_153),
.B(n_166),
.Y(n_125)
);

AOI21xp5_ASAP7_75t_L g126 ( 
.A1(n_127),
.A2(n_142),
.B(n_152),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_128),
.B(n_134),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_L g152 ( 
.A(n_128),
.B(n_134),
.Y(n_152)
);

CKINVDCx20_ASAP7_75t_R g129 ( 
.A(n_130),
.Y(n_129)
);

CKINVDCx20_ASAP7_75t_R g132 ( 
.A(n_133),
.Y(n_132)
);

AOI22xp5_ASAP7_75t_L g134 ( 
.A1(n_135),
.A2(n_136),
.B1(n_138),
.B2(n_139),
.Y(n_134)
);

CKINVDCx20_ASAP7_75t_R g135 ( 
.A(n_136),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_SL g154 ( 
.A(n_136),
.B(n_138),
.Y(n_154)
);

CKINVDCx20_ASAP7_75t_R g138 ( 
.A(n_139),
.Y(n_138)
);

OAI21xp5_ASAP7_75t_SL g142 ( 
.A1(n_143),
.A2(n_147),
.B(n_151),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_L g143 ( 
.A(n_144),
.B(n_145),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_L g151 ( 
.A(n_144),
.B(n_145),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_SL g147 ( 
.A(n_148),
.B(n_149),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_L g153 ( 
.A(n_154),
.B(n_155),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_SL g166 ( 
.A(n_154),
.B(n_155),
.Y(n_166)
);

XNOR2xp5_ASAP7_75t_L g155 ( 
.A(n_156),
.B(n_162),
.Y(n_155)
);

AOI22xp5_ASAP7_75t_L g156 ( 
.A1(n_157),
.A2(n_158),
.B1(n_159),
.B2(n_160),
.Y(n_156)
);

MAJIxp5_ASAP7_75t_L g168 ( 
.A(n_157),
.B(n_160),
.C(n_162),
.Y(n_168)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_158),
.Y(n_157)
);

CKINVDCx20_ASAP7_75t_R g159 ( 
.A(n_160),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_L g163 ( 
.A(n_164),
.B(n_165),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_L g167 ( 
.A(n_168),
.B(n_169),
.Y(n_167)
);

NOR2xp33_ASAP7_75t_L g184 ( 
.A(n_168),
.B(n_169),
.Y(n_184)
);

AOI22xp5_ASAP7_75t_L g169 ( 
.A1(n_170),
.A2(n_175),
.B1(n_182),
.B2(n_183),
.Y(n_169)
);

CKINVDCx20_ASAP7_75t_R g182 ( 
.A(n_170),
.Y(n_182)
);

XOR2xp5_ASAP7_75t_L g170 ( 
.A(n_171),
.B(n_172),
.Y(n_170)
);

NOR2xp33_ASAP7_75t_L g196 ( 
.A(n_171),
.B(n_172),
.Y(n_196)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_175),
.Y(n_183)
);

AOI22xp5_ASAP7_75t_L g175 ( 
.A1(n_176),
.A2(n_178),
.B1(n_179),
.B2(n_181),
.Y(n_175)
);

CKINVDCx20_ASAP7_75t_R g181 ( 
.A(n_176),
.Y(n_181)
);

MAJIxp5_ASAP7_75t_L g186 ( 
.A(n_178),
.B(n_181),
.C(n_182),
.Y(n_186)
);

CKINVDCx20_ASAP7_75t_R g178 ( 
.A(n_179),
.Y(n_178)
);

NOR2xp33_ASAP7_75t_L g185 ( 
.A(n_186),
.B(n_187),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_SL g197 ( 
.A(n_186),
.B(n_187),
.Y(n_197)
);

OAI22xp5_ASAP7_75t_SL g187 ( 
.A1(n_188),
.A2(n_189),
.B1(n_192),
.B2(n_193),
.Y(n_187)
);

MAJIxp5_ASAP7_75t_L g199 ( 
.A(n_188),
.B(n_194),
.C(n_196),
.Y(n_199)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_189),
.Y(n_188)
);

CKINVDCx20_ASAP7_75t_R g192 ( 
.A(n_193),
.Y(n_192)
);

XOR2x2_ASAP7_75t_SL g193 ( 
.A(n_194),
.B(n_196),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_L g198 ( 
.A(n_199),
.B(n_200),
.Y(n_198)
);

NOR2xp33_ASAP7_75t_SL g202 ( 
.A(n_199),
.B(n_200),
.Y(n_202)
);


endmodule