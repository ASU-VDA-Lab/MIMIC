module fake_jpeg_20031_n_190 (n_13, n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_190);

input n_13;
input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_190;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_14;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_84;
wire n_59;
wire n_98;
wire n_178;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_16;
wire n_49;
wire n_127;
wire n_76;
wire n_154;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_186;
wire n_44;
wire n_24;
wire n_143;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_177;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_161;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_176;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_189;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_120;
wire n_43;
wire n_32;
wire n_118;
wire n_140;
wire n_82;
wire n_128;
wire n_100;
wire n_96;

INVx6_ASAP7_75t_L g14 ( 
.A(n_7),
.Y(n_14)
);

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_7),
.Y(n_15)
);

CKINVDCx5p33_ASAP7_75t_R g16 ( 
.A(n_11),
.Y(n_16)
);

BUFx6f_ASAP7_75t_L g17 ( 
.A(n_5),
.Y(n_17)
);

INVxp67_ASAP7_75t_L g18 ( 
.A(n_0),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_4),
.Y(n_19)
);

BUFx3_ASAP7_75t_L g20 ( 
.A(n_10),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_7),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_0),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_9),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_4),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_9),
.Y(n_25)
);

BUFx12_ASAP7_75t_L g26 ( 
.A(n_2),
.Y(n_26)
);

BUFx4f_ASAP7_75t_L g27 ( 
.A(n_1),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_6),
.Y(n_28)
);

INVx11_ASAP7_75t_SL g29 ( 
.A(n_8),
.Y(n_29)
);

BUFx12f_ASAP7_75t_L g30 ( 
.A(n_0),
.Y(n_30)
);

INVx8_ASAP7_75t_L g31 ( 
.A(n_30),
.Y(n_31)
);

INVx8_ASAP7_75t_L g57 ( 
.A(n_31),
.Y(n_57)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_19),
.Y(n_32)
);

NOR2xp33_ASAP7_75t_L g47 ( 
.A(n_32),
.B(n_35),
.Y(n_47)
);

BUFx16f_ASAP7_75t_L g33 ( 
.A(n_16),
.Y(n_33)
);

INVx11_ASAP7_75t_L g60 ( 
.A(n_33),
.Y(n_60)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_27),
.Y(n_34)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_34),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g35 ( 
.A(n_26),
.B(n_1),
.Y(n_35)
);

BUFx3_ASAP7_75t_L g36 ( 
.A(n_30),
.Y(n_36)
);

INVx4_ASAP7_75t_L g64 ( 
.A(n_36),
.Y(n_64)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_27),
.Y(n_37)
);

INVx1_ASAP7_75t_SL g48 ( 
.A(n_37),
.Y(n_48)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_19),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_38),
.B(n_39),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g39 ( 
.A(n_26),
.B(n_1),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g40 ( 
.A(n_26),
.B(n_30),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_40),
.B(n_41),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g41 ( 
.A(n_30),
.B(n_2),
.Y(n_41)
);

INVx4_ASAP7_75t_L g42 ( 
.A(n_27),
.Y(n_42)
);

INVx3_ASAP7_75t_L g63 ( 
.A(n_42),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_SL g43 ( 
.A(n_16),
.B(n_15),
.Y(n_43)
);

OAI21xp5_ASAP7_75t_L g53 ( 
.A1(n_43),
.A2(n_18),
.B(n_22),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g44 ( 
.A(n_15),
.B(n_2),
.Y(n_44)
);

NAND2xp5_ASAP7_75t_L g62 ( 
.A(n_44),
.B(n_3),
.Y(n_62)
);

CKINVDCx16_ASAP7_75t_R g45 ( 
.A(n_21),
.Y(n_45)
);

INVx13_ASAP7_75t_L g59 ( 
.A(n_45),
.Y(n_59)
);

BUFx3_ASAP7_75t_L g46 ( 
.A(n_36),
.Y(n_46)
);

INVx4_ASAP7_75t_L g65 ( 
.A(n_46),
.Y(n_65)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_36),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g76 ( 
.A(n_49),
.Y(n_76)
);

INVx2_ASAP7_75t_L g50 ( 
.A(n_34),
.Y(n_50)
);

INVx6_ASAP7_75t_L g87 ( 
.A(n_50),
.Y(n_87)
);

AOI22xp33_ASAP7_75t_SL g51 ( 
.A1(n_42),
.A2(n_14),
.B1(n_29),
.B2(n_28),
.Y(n_51)
);

INVxp67_ASAP7_75t_L g70 ( 
.A(n_51),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_SL g75 ( 
.A(n_53),
.B(n_33),
.Y(n_75)
);

OAI22xp33_ASAP7_75t_SL g55 ( 
.A1(n_32),
.A2(n_14),
.B1(n_18),
.B2(n_21),
.Y(n_55)
);

OAI22xp5_ASAP7_75t_SL g74 ( 
.A1(n_55),
.A2(n_38),
.B1(n_45),
.B2(n_37),
.Y(n_74)
);

AOI22xp33_ASAP7_75t_SL g56 ( 
.A1(n_42),
.A2(n_28),
.B1(n_22),
.B2(n_23),
.Y(n_56)
);

CKINVDCx16_ASAP7_75t_R g86 ( 
.A(n_56),
.Y(n_86)
);

INVx6_ASAP7_75t_L g61 ( 
.A(n_31),
.Y(n_61)
);

INVx8_ASAP7_75t_L g78 ( 
.A(n_61),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_L g85 ( 
.A(n_62),
.B(n_58),
.Y(n_85)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_59),
.Y(n_66)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_66),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_47),
.B(n_43),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_SL g110 ( 
.A(n_67),
.B(n_81),
.Y(n_110)
);

INVx3_ASAP7_75t_L g68 ( 
.A(n_64),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_68),
.B(n_73),
.Y(n_94)
);

INVx2_ASAP7_75t_L g69 ( 
.A(n_63),
.Y(n_69)
);

INVx4_ASAP7_75t_L g102 ( 
.A(n_69),
.Y(n_102)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_59),
.Y(n_71)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_71),
.Y(n_98)
);

INVx2_ASAP7_75t_L g72 ( 
.A(n_63),
.Y(n_72)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_72),
.Y(n_111)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_59),
.Y(n_73)
);

OAI22xp33_ASAP7_75t_SL g112 ( 
.A1(n_74),
.A2(n_80),
.B1(n_20),
.B2(n_4),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_75),
.B(n_77),
.Y(n_99)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_54),
.Y(n_77)
);

O2A1O1Ixp33_ASAP7_75t_SL g79 ( 
.A1(n_53),
.A2(n_33),
.B(n_38),
.C(n_31),
.Y(n_79)
);

AO22x1_ASAP7_75t_SL g113 ( 
.A1(n_79),
.A2(n_3),
.B1(n_5),
.B2(n_6),
.Y(n_113)
);

AOI22xp33_ASAP7_75t_L g80 ( 
.A1(n_52),
.A2(n_37),
.B1(n_34),
.B2(n_41),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_47),
.B(n_44),
.Y(n_81)
);

BUFx8_ASAP7_75t_L g82 ( 
.A(n_60),
.Y(n_82)
);

INVx1_ASAP7_75t_SL g100 ( 
.A(n_82),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_52),
.B(n_39),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_83),
.B(n_84),
.Y(n_108)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_54),
.Y(n_84)
);

OR2x2_ASAP7_75t_L g115 ( 
.A(n_85),
.B(n_92),
.Y(n_115)
);

O2A1O1Ixp33_ASAP7_75t_L g88 ( 
.A1(n_58),
.A2(n_40),
.B(n_33),
.C(n_35),
.Y(n_88)
);

OAI22xp5_ASAP7_75t_SL g97 ( 
.A1(n_88),
.A2(n_93),
.B1(n_61),
.B2(n_57),
.Y(n_97)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_64),
.Y(n_89)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_89),
.Y(n_103)
);

INVx13_ASAP7_75t_L g90 ( 
.A(n_60),
.Y(n_90)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_90),
.Y(n_105)
);

AND2x2_ASAP7_75t_L g91 ( 
.A(n_50),
.B(n_31),
.Y(n_91)
);

AND2x2_ASAP7_75t_L g104 ( 
.A(n_91),
.B(n_61),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_SL g92 ( 
.A(n_62),
.B(n_25),
.Y(n_92)
);

OAI22xp5_ASAP7_75t_SL g93 ( 
.A1(n_48),
.A2(n_24),
.B1(n_17),
.B2(n_33),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_L g96 ( 
.A(n_88),
.B(n_48),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g116 ( 
.A(n_96),
.B(n_91),
.Y(n_116)
);

AOI22xp5_ASAP7_75t_L g121 ( 
.A1(n_97),
.A2(n_106),
.B1(n_109),
.B2(n_112),
.Y(n_121)
);

MAJx2_ASAP7_75t_L g101 ( 
.A(n_79),
.B(n_20),
.C(n_24),
.Y(n_101)
);

XNOR2xp5_ASAP7_75t_L g129 ( 
.A(n_101),
.B(n_97),
.Y(n_129)
);

OAI21xp5_ASAP7_75t_SL g119 ( 
.A1(n_104),
.A2(n_113),
.B(n_70),
.Y(n_119)
);

OAI22xp5_ASAP7_75t_SL g106 ( 
.A1(n_86),
.A2(n_57),
.B1(n_17),
.B2(n_49),
.Y(n_106)
);

HB1xp67_ASAP7_75t_L g107 ( 
.A(n_82),
.Y(n_107)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_107),
.Y(n_117)
);

OAI22xp5_ASAP7_75t_SL g109 ( 
.A1(n_70),
.A2(n_57),
.B1(n_49),
.B2(n_46),
.Y(n_109)
);

NOR2x1_ASAP7_75t_L g114 ( 
.A(n_74),
.B(n_3),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_SL g127 ( 
.A(n_114),
.B(n_115),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_L g141 ( 
.A(n_116),
.B(n_118),
.Y(n_141)
);

CKINVDCx20_ASAP7_75t_R g118 ( 
.A(n_111),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_SL g139 ( 
.A(n_119),
.B(n_120),
.Y(n_139)
);

CKINVDCx20_ASAP7_75t_R g120 ( 
.A(n_103),
.Y(n_120)
);

OAI22xp5_ASAP7_75t_SL g122 ( 
.A1(n_96),
.A2(n_87),
.B1(n_93),
.B2(n_69),
.Y(n_122)
);

INVxp67_ASAP7_75t_L g134 ( 
.A(n_122),
.Y(n_134)
);

OAI22xp5_ASAP7_75t_L g123 ( 
.A1(n_99),
.A2(n_87),
.B1(n_78),
.B2(n_72),
.Y(n_123)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_123),
.Y(n_136)
);

OAI21xp5_ASAP7_75t_L g124 ( 
.A1(n_101),
.A2(n_91),
.B(n_90),
.Y(n_124)
);

XNOR2xp5_ASAP7_75t_L g142 ( 
.A(n_124),
.B(n_129),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_L g125 ( 
.A(n_113),
.B(n_78),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_SL g143 ( 
.A(n_125),
.B(n_127),
.Y(n_143)
);

BUFx3_ASAP7_75t_L g126 ( 
.A(n_102),
.Y(n_126)
);

BUFx12f_ASAP7_75t_L g144 ( 
.A(n_126),
.Y(n_144)
);

MAJIxp5_ASAP7_75t_L g128 ( 
.A(n_108),
.B(n_68),
.C(n_65),
.Y(n_128)
);

MAJIxp5_ASAP7_75t_L g140 ( 
.A(n_128),
.B(n_94),
.C(n_109),
.Y(n_140)
);

BUFx6f_ASAP7_75t_L g130 ( 
.A(n_102),
.Y(n_130)
);

INVx6_ASAP7_75t_L g135 ( 
.A(n_130),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_SL g131 ( 
.A(n_110),
.B(n_12),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_L g133 ( 
.A(n_131),
.B(n_132),
.Y(n_133)
);

OAI22xp5_ASAP7_75t_SL g132 ( 
.A1(n_114),
.A2(n_113),
.B1(n_115),
.B2(n_104),
.Y(n_132)
);

XOR2xp5_ASAP7_75t_SL g137 ( 
.A(n_124),
.B(n_104),
.Y(n_137)
);

XOR2xp5_ASAP7_75t_L g150 ( 
.A(n_137),
.B(n_140),
.Y(n_150)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_117),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_L g149 ( 
.A(n_138),
.B(n_145),
.Y(n_149)
);

CKINVDCx20_ASAP7_75t_R g145 ( 
.A(n_117),
.Y(n_145)
);

A2O1A1O1Ixp25_ASAP7_75t_L g146 ( 
.A1(n_129),
.A2(n_106),
.B(n_98),
.C(n_95),
.D(n_103),
.Y(n_146)
);

AND2x2_ASAP7_75t_L g147 ( 
.A(n_146),
.B(n_121),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_SL g163 ( 
.A(n_147),
.B(n_157),
.Y(n_163)
);

OAI21xp5_ASAP7_75t_L g148 ( 
.A1(n_139),
.A2(n_119),
.B(n_116),
.Y(n_148)
);

INVxp67_ASAP7_75t_L g165 ( 
.A(n_148),
.Y(n_165)
);

OAI22xp5_ASAP7_75t_SL g151 ( 
.A1(n_134),
.A2(n_121),
.B1(n_125),
.B2(n_122),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_L g162 ( 
.A(n_151),
.B(n_155),
.Y(n_162)
);

NOR2xp33_ASAP7_75t_L g152 ( 
.A(n_133),
.B(n_128),
.Y(n_152)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_152),
.Y(n_160)
);

MAJIxp5_ASAP7_75t_L g153 ( 
.A(n_142),
.B(n_132),
.C(n_118),
.Y(n_153)
);

MAJIxp5_ASAP7_75t_L g164 ( 
.A(n_153),
.B(n_144),
.C(n_76),
.Y(n_164)
);

OAI22xp5_ASAP7_75t_SL g154 ( 
.A1(n_134),
.A2(n_136),
.B1(n_141),
.B2(n_143),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_L g168 ( 
.A(n_154),
.B(n_156),
.Y(n_168)
);

NOR2xp33_ASAP7_75t_SL g155 ( 
.A(n_142),
.B(n_11),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_SL g156 ( 
.A(n_140),
.B(n_12),
.Y(n_156)
);

NOR2xp33_ASAP7_75t_L g157 ( 
.A(n_144),
.B(n_126),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_L g158 ( 
.A(n_135),
.B(n_105),
.Y(n_158)
);

XNOR2xp5_ASAP7_75t_L g167 ( 
.A(n_158),
.B(n_159),
.Y(n_167)
);

OAI22xp5_ASAP7_75t_SL g159 ( 
.A1(n_137),
.A2(n_105),
.B1(n_65),
.B2(n_100),
.Y(n_159)
);

MAJIxp5_ASAP7_75t_L g161 ( 
.A(n_150),
.B(n_146),
.C(n_130),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_L g170 ( 
.A(n_161),
.B(n_166),
.Y(n_170)
);

MAJIxp5_ASAP7_75t_L g173 ( 
.A(n_164),
.B(n_159),
.C(n_154),
.Y(n_173)
);

MAJIxp5_ASAP7_75t_L g166 ( 
.A(n_150),
.B(n_144),
.C(n_76),
.Y(n_166)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_167),
.Y(n_169)
);

NOR2xp33_ASAP7_75t_L g177 ( 
.A(n_169),
.B(n_172),
.Y(n_177)
);

OAI22xp5_ASAP7_75t_SL g171 ( 
.A1(n_165),
.A2(n_151),
.B1(n_153),
.B2(n_147),
.Y(n_171)
);

AOI22xp5_ASAP7_75t_L g178 ( 
.A1(n_171),
.A2(n_175),
.B1(n_164),
.B2(n_135),
.Y(n_178)
);

AOI21xp5_ASAP7_75t_SL g172 ( 
.A1(n_163),
.A2(n_148),
.B(n_149),
.Y(n_172)
);

NOR2xp33_ASAP7_75t_SL g180 ( 
.A(n_173),
.B(n_174),
.Y(n_180)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_168),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_L g175 ( 
.A(n_160),
.B(n_162),
.Y(n_175)
);

OR2x2_ASAP7_75t_L g176 ( 
.A(n_172),
.B(n_165),
.Y(n_176)
);

NOR2xp33_ASAP7_75t_L g181 ( 
.A(n_176),
.B(n_178),
.Y(n_181)
);

AOI22xp33_ASAP7_75t_L g179 ( 
.A1(n_173),
.A2(n_100),
.B1(n_82),
.B2(n_6),
.Y(n_179)
);

AOI21x1_ASAP7_75t_SL g183 ( 
.A1(n_179),
.A2(n_171),
.B(n_5),
.Y(n_183)
);

NOR2xp67_ASAP7_75t_L g182 ( 
.A(n_176),
.B(n_177),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_L g184 ( 
.A(n_182),
.B(n_180),
.Y(n_184)
);

MAJIxp5_ASAP7_75t_L g185 ( 
.A(n_183),
.B(n_170),
.C(n_179),
.Y(n_185)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_184),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_L g187 ( 
.A(n_185),
.B(n_181),
.Y(n_187)
);

AOI22xp5_ASAP7_75t_SL g188 ( 
.A1(n_187),
.A2(n_13),
.B1(n_8),
.B2(n_10),
.Y(n_188)
);

XOR2xp5_ASAP7_75t_L g189 ( 
.A(n_188),
.B(n_186),
.Y(n_189)
);

XOR2xp5_ASAP7_75t_L g190 ( 
.A(n_189),
.B(n_13),
.Y(n_190)
);


endmodule