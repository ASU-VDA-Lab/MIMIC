module fake_netlist_6_4173_n_74 (n_16, n_1, n_9, n_8, n_18, n_10, n_21, n_6, n_15, n_3, n_14, n_0, n_4, n_13, n_11, n_17, n_12, n_20, n_7, n_2, n_5, n_19, n_74);

input n_16;
input n_1;
input n_9;
input n_8;
input n_18;
input n_10;
input n_21;
input n_6;
input n_15;
input n_3;
input n_14;
input n_0;
input n_4;
input n_13;
input n_11;
input n_17;
input n_12;
input n_20;
input n_7;
input n_2;
input n_5;
input n_19;

output n_74;

wire n_41;
wire n_52;
wire n_45;
wire n_46;
wire n_34;
wire n_42;
wire n_70;
wire n_24;
wire n_71;
wire n_37;
wire n_33;
wire n_54;
wire n_67;
wire n_27;
wire n_38;
wire n_72;
wire n_61;
wire n_39;
wire n_63;
wire n_60;
wire n_59;
wire n_73;
wire n_32;
wire n_66;
wire n_36;
wire n_22;
wire n_26;
wire n_68;
wire n_55;
wire n_35;
wire n_28;
wire n_23;
wire n_58;
wire n_69;
wire n_50;
wire n_49;
wire n_30;
wire n_64;
wire n_43;
wire n_47;
wire n_48;
wire n_29;
wire n_62;
wire n_31;
wire n_65;
wire n_40;
wire n_57;
wire n_25;
wire n_53;
wire n_51;
wire n_44;
wire n_56;

OAI21x1_ASAP7_75t_L g22 ( 
.A1(n_14),
.A2(n_19),
.B(n_9),
.Y(n_22)
);

OAI22xp5_ASAP7_75t_L g23 ( 
.A1(n_4),
.A2(n_6),
.B1(n_3),
.B2(n_11),
.Y(n_23)
);

NAND2xp5_ASAP7_75t_L g24 ( 
.A(n_21),
.B(n_8),
.Y(n_24)
);

INVx2_ASAP7_75t_L g25 ( 
.A(n_15),
.Y(n_25)
);

AND2x2_ASAP7_75t_L g26 ( 
.A(n_3),
.B(n_10),
.Y(n_26)
);

INVx3_ASAP7_75t_L g27 ( 
.A(n_16),
.Y(n_27)
);

OAI22x1_ASAP7_75t_SL g28 ( 
.A1(n_17),
.A2(n_5),
.B1(n_0),
.B2(n_4),
.Y(n_28)
);

NAND2xp5_ASAP7_75t_L g29 ( 
.A(n_1),
.B(n_7),
.Y(n_29)
);

AND2x2_ASAP7_75t_L g30 ( 
.A(n_18),
.B(n_1),
.Y(n_30)
);

NAND2xp5_ASAP7_75t_L g31 ( 
.A(n_0),
.B(n_13),
.Y(n_31)
);

INVx2_ASAP7_75t_L g32 ( 
.A(n_20),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_5),
.Y(n_33)
);

INVx5_ASAP7_75t_L g34 ( 
.A(n_12),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_2),
.Y(n_35)
);

INVx3_ASAP7_75t_L g36 ( 
.A(n_2),
.Y(n_36)
);

NAND2xp5_ASAP7_75t_L g37 ( 
.A(n_27),
.B(n_32),
.Y(n_37)
);

INVx3_ASAP7_75t_L g38 ( 
.A(n_35),
.Y(n_38)
);

NAND2xp5_ASAP7_75t_SL g39 ( 
.A(n_26),
.B(n_30),
.Y(n_39)
);

AOI221xp5_ASAP7_75t_L g40 ( 
.A1(n_36),
.A2(n_33),
.B1(n_28),
.B2(n_35),
.C(n_23),
.Y(n_40)
);

NAND2xp5_ASAP7_75t_SL g41 ( 
.A(n_26),
.B(n_30),
.Y(n_41)
);

INVx2_ASAP7_75t_L g42 ( 
.A(n_35),
.Y(n_42)
);

INVx2_ASAP7_75t_L g43 ( 
.A(n_35),
.Y(n_43)
);

INVx2_ASAP7_75t_L g44 ( 
.A(n_35),
.Y(n_44)
);

NAND2xp5_ASAP7_75t_SL g45 ( 
.A(n_36),
.B(n_27),
.Y(n_45)
);

NAND2xp5_ASAP7_75t_SL g46 ( 
.A(n_36),
.B(n_27),
.Y(n_46)
);

INVx2_ASAP7_75t_L g47 ( 
.A(n_42),
.Y(n_47)
);

BUFx4f_ASAP7_75t_SL g48 ( 
.A(n_45),
.Y(n_48)
);

AOI21xp33_ASAP7_75t_L g49 ( 
.A1(n_39),
.A2(n_31),
.B(n_29),
.Y(n_49)
);

INVxp67_ASAP7_75t_SL g50 ( 
.A(n_37),
.Y(n_50)
);

INVx2_ASAP7_75t_L g51 ( 
.A(n_47),
.Y(n_51)
);

INVx3_ASAP7_75t_L g52 ( 
.A(n_47),
.Y(n_52)
);

INVx2_ASAP7_75t_L g53 ( 
.A(n_48),
.Y(n_53)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_50),
.Y(n_54)
);

INVx2_ASAP7_75t_L g55 ( 
.A(n_49),
.Y(n_55)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_52),
.Y(n_56)
);

NOR2x1_ASAP7_75t_L g57 ( 
.A(n_55),
.B(n_24),
.Y(n_57)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_51),
.Y(n_58)
);

AND2x2_ASAP7_75t_L g59 ( 
.A(n_54),
.B(n_49),
.Y(n_59)
);

HB1xp67_ASAP7_75t_L g60 ( 
.A(n_54),
.Y(n_60)
);

OR2x2_ASAP7_75t_L g61 ( 
.A(n_59),
.B(n_53),
.Y(n_61)
);

OR2x2_ASAP7_75t_L g62 ( 
.A(n_60),
.B(n_33),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_SL g63 ( 
.A(n_57),
.B(n_40),
.Y(n_63)
);

O2A1O1Ixp33_ASAP7_75t_R g64 ( 
.A1(n_61),
.A2(n_58),
.B(n_25),
.C(n_32),
.Y(n_64)
);

NAND4xp25_ASAP7_75t_SL g65 ( 
.A(n_64),
.B(n_62),
.C(n_63),
.D(n_25),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_64),
.B(n_56),
.Y(n_66)
);

NOR2x1_ASAP7_75t_L g67 ( 
.A(n_65),
.B(n_46),
.Y(n_67)
);

NOR2xp67_ASAP7_75t_L g68 ( 
.A(n_66),
.B(n_34),
.Y(n_68)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_68),
.Y(n_69)
);

AOI221xp5_ASAP7_75t_L g70 ( 
.A1(n_67),
.A2(n_41),
.B1(n_34),
.B2(n_43),
.C(n_44),
.Y(n_70)
);

AOI21x1_ASAP7_75t_L g71 ( 
.A1(n_69),
.A2(n_22),
.B(n_38),
.Y(n_71)
);

OA22x2_ASAP7_75t_L g72 ( 
.A1(n_70),
.A2(n_22),
.B1(n_38),
.B2(n_34),
.Y(n_72)
);

OAI21x1_ASAP7_75t_L g73 ( 
.A1(n_71),
.A2(n_34),
.B(n_72),
.Y(n_73)
);

OR2x6_ASAP7_75t_L g74 ( 
.A(n_73),
.B(n_34),
.Y(n_74)
);


endmodule