module real_jpeg_15116_n_17 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_16, n_3, n_10, n_9, n_17);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_16;
input n_3;
input n_10;
input n_9;

output n_17;

wire n_384;
wire n_37;
wire n_430;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_300;
wire n_415;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_199;
wire n_95;
wire n_441;
wire n_238;
wire n_67;
wire n_350;
wire n_235;
wire n_107;
wire n_369;
wire n_376;
wire n_354;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_355;
wire n_123;
wire n_425;
wire n_50;
wire n_409;
wire n_186;
wire n_137;
wire n_72;
wire n_440;
wire n_171;
wire n_151;
wire n_272;
wire n_198;
wire n_203;
wire n_23;
wire n_362;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_326;
wire n_339;
wire n_80;
wire n_30;
wire n_328;
wire n_149;
wire n_366;
wire n_332;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_353;
wire n_230;
wire n_417;
wire n_428;
wire n_128;
wire n_202;
wire n_216;
wire n_367;
wire n_127;
wire n_365;
wire n_356;
wire n_423;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_422;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_348;
wire n_252;
wire n_363;
wire n_310;
wire n_345;
wire n_78;
wire n_83;
wire n_288;
wire n_221;
wire n_393;
wire n_104;
wire n_153;
wire n_443;
wire n_337;
wire n_131;
wire n_439;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_378;
wire n_200;
wire n_432;
wire n_335;
wire n_214;
wire n_113;
wire n_251;
wire n_139;
wire n_33;
wire n_175;
wire n_338;
wire n_156;
wire n_387;
wire n_434;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_390;
wire n_77;
wire n_399;
wire n_219;
wire n_372;
wire n_122;
wire n_19;
wire n_262;
wire n_334;
wire n_383;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_426;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_371;
wire n_410;
wire n_421;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_382;
wire n_411;
wire n_20;
wire n_278;
wire n_314;
wire n_103;
wire n_232;
wire n_212;
wire n_284;
wire n_402;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_213;
wire n_25;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_407;
wire n_419;
wire n_386;
wire n_341;
wire n_331;
wire n_49;
wire n_68;
wire n_395;
wire n_146;
wire n_286;
wire n_166;
wire n_176;
wire n_215;
wire n_323;
wire n_312;
wire n_325;
wire n_307;
wire n_316;
wire n_161;
wire n_207;
wire n_431;
wire n_420;
wire n_357;
wire n_237;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_380;
wire n_414;
wire n_140;
wire n_126;
wire n_342;
wire n_120;
wire n_155;
wire n_412;
wire n_405;
wire n_319;
wire n_93;
wire n_242;
wire n_142;
wire n_397;
wire n_76;
wire n_403;
wire n_79;
wire n_282;
wire n_147;
wire n_359;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_18;
wire n_145;
wire n_266;
wire n_377;
wire n_109;
wire n_391;
wire n_427;
wire n_401;
wire n_148;
wire n_373;
wire n_396;
wire n_392;
wire n_196;
wire n_375;
wire n_298;
wire n_330;
wire n_333;
wire n_152;
wire n_270;
wire n_159;
wire n_429;
wire n_347;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_336;
wire n_258;
wire n_150;
wire n_41;
wire n_74;
wire n_404;
wire n_204;
wire n_158;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_413;
wire n_75;
wire n_346;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_119;
wire n_283;
wire n_358;
wire n_181;
wire n_256;
wire n_253;
wire n_273;
wire n_54;
wire n_168;
wire n_38;
wire n_442;
wire n_385;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_349;
wire n_418;
wire n_292;
wire n_343;
wire n_64;
wire n_291;
wire n_236;
wire n_370;
wire n_276;
wire n_374;
wire n_287;
wire n_388;
wire n_174;
wire n_400;
wire n_255;
wire n_243;
wire n_299;
wire n_352;
wire n_56;
wire n_293;
wire n_275;
wire n_381;
wire n_227;
wire n_229;
wire n_379;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_360;
wire n_398;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_45;
wire n_437;
wire n_268;
wire n_42;
wire n_313;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_416;
wire n_143;
wire n_351;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_406;
wire n_303;
wire n_321;
wire n_100;
wire n_368;
wire n_51;
wire n_205;
wire n_361;
wire n_261;
wire n_86;
wire n_324;
wire n_70;
wire n_435;
wire n_32;
wire n_228;
wire n_389;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_438;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_394;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_436;
wire n_169;
wire n_88;
wire n_167;
wire n_295;
wire n_424;
wire n_133;
wire n_257;
wire n_344;
wire n_210;
wire n_206;
wire n_408;
wire n_85;
wire n_96;
wire n_308;
wire n_433;
wire n_364;

AOI22x1_ASAP7_75t_L g42 ( 
.A1(n_0),
.A2(n_6),
.B1(n_43),
.B2(n_47),
.Y(n_42)
);

NAND2xp5_ASAP7_75t_SL g118 ( 
.A(n_0),
.B(n_119),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_SL g130 ( 
.A(n_0),
.B(n_131),
.Y(n_130)
);

AND2x2_ASAP7_75t_L g207 ( 
.A(n_0),
.B(n_208),
.Y(n_207)
);

AOI31xp67_ASAP7_75t_L g247 ( 
.A1(n_0),
.A2(n_42),
.A3(n_248),
.B(n_252),
.Y(n_247)
);

NAND2xp5_ASAP7_75t_L g284 ( 
.A(n_0),
.B(n_285),
.Y(n_284)
);

NAND2xp5_ASAP7_75t_L g307 ( 
.A(n_0),
.B(n_308),
.Y(n_307)
);

AND2x2_ASAP7_75t_L g311 ( 
.A(n_0),
.B(n_312),
.Y(n_311)
);

NAND2xp5_ASAP7_75t_L g352 ( 
.A(n_0),
.B(n_353),
.Y(n_352)
);

AND2x2_ASAP7_75t_L g136 ( 
.A(n_1),
.B(n_137),
.Y(n_136)
);

INVx1_ASAP7_75t_SL g160 ( 
.A(n_1),
.Y(n_160)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_2),
.Y(n_63)
);

BUFx6f_ASAP7_75t_L g116 ( 
.A(n_2),
.Y(n_116)
);

BUFx3_ASAP7_75t_L g176 ( 
.A(n_2),
.Y(n_176)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_2),
.Y(n_212)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_3),
.Y(n_78)
);

BUFx5_ASAP7_75t_L g83 ( 
.A(n_3),
.Y(n_83)
);

BUFx6f_ASAP7_75t_L g101 ( 
.A(n_3),
.Y(n_101)
);

BUFx6f_ASAP7_75t_L g171 ( 
.A(n_3),
.Y(n_171)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_3),
.Y(n_217)
);

BUFx6f_ASAP7_75t_L g340 ( 
.A(n_3),
.Y(n_340)
);

NAND2xp5_ASAP7_75t_SL g72 ( 
.A(n_4),
.B(n_73),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_L g262 ( 
.A(n_4),
.B(n_263),
.Y(n_262)
);

NAND2xp5_ASAP7_75t_SL g280 ( 
.A(n_4),
.B(n_281),
.Y(n_280)
);

NAND2xp5_ASAP7_75t_L g303 ( 
.A(n_4),
.B(n_304),
.Y(n_303)
);

NAND2xp5_ASAP7_75t_L g348 ( 
.A(n_4),
.B(n_349),
.Y(n_348)
);

NAND2xp5_ASAP7_75t_SL g357 ( 
.A(n_4),
.B(n_358),
.Y(n_357)
);

NAND2xp5_ASAP7_75t_SL g365 ( 
.A(n_4),
.B(n_366),
.Y(n_365)
);

AND2x2_ASAP7_75t_L g75 ( 
.A(n_5),
.B(n_76),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_L g113 ( 
.A(n_5),
.B(n_114),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_SL g122 ( 
.A(n_5),
.B(n_123),
.Y(n_122)
);

AND2x2_ASAP7_75t_L g149 ( 
.A(n_5),
.B(n_150),
.Y(n_149)
);

CKINVDCx16_ASAP7_75t_R g202 ( 
.A(n_5),
.Y(n_202)
);

AND2x2_ASAP7_75t_L g259 ( 
.A(n_5),
.B(n_46),
.Y(n_259)
);

NAND2xp5_ASAP7_75t_L g423 ( 
.A(n_5),
.B(n_424),
.Y(n_423)
);

AND2x2_ASAP7_75t_L g32 ( 
.A(n_6),
.B(n_33),
.Y(n_32)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_6),
.B(n_100),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_SL g177 ( 
.A(n_6),
.B(n_178),
.Y(n_177)
);

CKINVDCx16_ASAP7_75t_R g253 ( 
.A(n_6),
.Y(n_253)
);

NAND2x1_ASAP7_75t_L g427 ( 
.A(n_6),
.B(n_428),
.Y(n_427)
);

INVx2_ASAP7_75t_L g40 ( 
.A(n_7),
.Y(n_40)
);

BUFx5_ASAP7_75t_L g46 ( 
.A(n_7),
.Y(n_46)
);

BUFx5_ASAP7_75t_L g205 ( 
.A(n_7),
.Y(n_205)
);

AND2x2_ASAP7_75t_L g64 ( 
.A(n_8),
.B(n_35),
.Y(n_64)
);

AND2x2_ASAP7_75t_L g80 ( 
.A(n_8),
.B(n_81),
.Y(n_80)
);

NAND2x1_ASAP7_75t_L g106 ( 
.A(n_8),
.B(n_107),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_L g173 ( 
.A(n_8),
.B(n_174),
.Y(n_173)
);

AND2x2_ASAP7_75t_SL g203 ( 
.A(n_8),
.B(n_204),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_SL g412 ( 
.A(n_8),
.B(n_413),
.Y(n_412)
);

INVx3_ASAP7_75t_L g71 ( 
.A(n_9),
.Y(n_71)
);

BUFx3_ASAP7_75t_L g108 ( 
.A(n_9),
.Y(n_108)
);

BUFx6f_ASAP7_75t_L g180 ( 
.A(n_9),
.Y(n_180)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_9),
.Y(n_222)
);

BUFx5_ASAP7_75t_L g286 ( 
.A(n_9),
.Y(n_286)
);

AND2x2_ASAP7_75t_L g58 ( 
.A(n_10),
.B(n_59),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_L g84 ( 
.A(n_10),
.B(n_85),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g110 ( 
.A(n_10),
.B(n_111),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_SL g153 ( 
.A(n_10),
.B(n_154),
.Y(n_153)
);

AND2x2_ASAP7_75t_L g218 ( 
.A(n_10),
.B(n_219),
.Y(n_218)
);

AND2x2_ASAP7_75t_L g317 ( 
.A(n_10),
.B(n_45),
.Y(n_317)
);

NAND2xp5_ASAP7_75t_L g319 ( 
.A(n_10),
.B(n_320),
.Y(n_319)
);

NAND2xp5_ASAP7_75t_L g334 ( 
.A(n_10),
.B(n_335),
.Y(n_334)
);

NAND2xp5_ASAP7_75t_SL g27 ( 
.A(n_11),
.B(n_28),
.Y(n_27)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_11),
.Y(n_55)
);

AND2x2_ASAP7_75t_L g68 ( 
.A(n_11),
.B(n_69),
.Y(n_68)
);

AND2x2_ASAP7_75t_L g95 ( 
.A(n_11),
.B(n_96),
.Y(n_95)
);

AND2x2_ASAP7_75t_L g127 ( 
.A(n_11),
.B(n_128),
.Y(n_127)
);

AND2x2_ASAP7_75t_L g213 ( 
.A(n_11),
.B(n_214),
.Y(n_213)
);

AND2x2_ASAP7_75t_L g258 ( 
.A(n_11),
.B(n_35),
.Y(n_258)
);

AND2x2_ASAP7_75t_L g321 ( 
.A(n_11),
.B(n_37),
.Y(n_321)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_12),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g121 ( 
.A(n_12),
.Y(n_121)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_13),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g251 ( 
.A(n_13),
.Y(n_251)
);

BUFx12f_ASAP7_75t_L g35 ( 
.A(n_14),
.Y(n_35)
);

INVx2_ASAP7_75t_L g142 ( 
.A(n_14),
.Y(n_142)
);

BUFx4f_ASAP7_75t_L g162 ( 
.A(n_14),
.Y(n_162)
);

BUFx6f_ASAP7_75t_L g316 ( 
.A(n_14),
.Y(n_316)
);

AND2x2_ASAP7_75t_L g36 ( 
.A(n_15),
.B(n_37),
.Y(n_36)
);

AND2x2_ASAP7_75t_L g139 ( 
.A(n_15),
.B(n_140),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_SL g168 ( 
.A(n_15),
.B(n_169),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_L g432 ( 
.A(n_15),
.B(n_107),
.Y(n_432)
);

INVx2_ASAP7_75t_L g30 ( 
.A(n_16),
.Y(n_30)
);

BUFx3_ASAP7_75t_L g74 ( 
.A(n_16),
.Y(n_74)
);

XNOR2xp5_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_400),
.Y(n_17)
);

OAI21xp5_ASAP7_75t_L g18 ( 
.A1(n_19),
.A2(n_230),
.B(n_399),
.Y(n_18)
);

AND2x2_ASAP7_75t_SL g19 ( 
.A(n_20),
.B(n_183),
.Y(n_19)
);

OR2x2_ASAP7_75t_L g399 ( 
.A(n_20),
.B(n_183),
.Y(n_399)
);

XNOR2xp5_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_102),
.Y(n_20)
);

INVx1_ASAP7_75t_L g404 ( 
.A(n_21),
.Y(n_404)
);

MAJIxp5_ASAP7_75t_L g21 ( 
.A(n_22),
.B(n_65),
.C(n_89),
.Y(n_21)
);

INVxp33_ASAP7_75t_SL g22 ( 
.A(n_23),
.Y(n_22)
);

XNOR2xp5_ASAP7_75t_L g186 ( 
.A(n_23),
.B(n_187),
.Y(n_186)
);

MAJIxp5_ASAP7_75t_L g23 ( 
.A(n_24),
.B(n_41),
.C(n_52),
.Y(n_23)
);

XNOR2xp5_ASAP7_75t_L g265 ( 
.A(n_24),
.B(n_266),
.Y(n_265)
);

XNOR2xp5_ASAP7_75t_L g24 ( 
.A(n_25),
.B(n_31),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_26),
.Y(n_25)
);

XNOR2xp5_ASAP7_75t_L g436 ( 
.A(n_26),
.B(n_149),
.Y(n_436)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_27),
.Y(n_26)
);

MAJIxp5_ASAP7_75t_L g92 ( 
.A(n_27),
.B(n_32),
.C(n_36),
.Y(n_92)
);

INVx4_ASAP7_75t_L g28 ( 
.A(n_29),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_30),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g134 ( 
.A(n_30),
.Y(n_134)
);

XNOR2xp5_ASAP7_75t_L g31 ( 
.A(n_32),
.B(n_36),
.Y(n_31)
);

INVx2_ASAP7_75t_L g33 ( 
.A(n_34),
.Y(n_33)
);

INVx2_ASAP7_75t_L g34 ( 
.A(n_35),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g201 ( 
.A(n_35),
.Y(n_201)
);

INVx2_ASAP7_75t_L g37 ( 
.A(n_38),
.Y(n_37)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_39),
.Y(n_38)
);

INVx2_ASAP7_75t_L g39 ( 
.A(n_40),
.Y(n_39)
);

INVx3_ASAP7_75t_L g137 ( 
.A(n_40),
.Y(n_137)
);

AOI22xp5_ASAP7_75t_SL g266 ( 
.A1(n_41),
.A2(n_42),
.B1(n_52),
.B2(n_267),
.Y(n_266)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_42),
.Y(n_41)
);

INVx4_ASAP7_75t_L g43 ( 
.A(n_44),
.Y(n_43)
);

INVx6_ASAP7_75t_L g44 ( 
.A(n_45),
.Y(n_44)
);

BUFx12f_ASAP7_75t_L g45 ( 
.A(n_46),
.Y(n_45)
);

INVx2_ASAP7_75t_L g47 ( 
.A(n_48),
.Y(n_47)
);

HB1xp67_ASAP7_75t_L g48 ( 
.A(n_49),
.Y(n_48)
);

INVx2_ASAP7_75t_SL g49 ( 
.A(n_50),
.Y(n_49)
);

BUFx5_ASAP7_75t_L g50 ( 
.A(n_51),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g88 ( 
.A(n_51),
.Y(n_88)
);

BUFx6f_ASAP7_75t_L g97 ( 
.A(n_51),
.Y(n_97)
);

INVx2_ASAP7_75t_L g152 ( 
.A(n_51),
.Y(n_152)
);

BUFx6f_ASAP7_75t_L g283 ( 
.A(n_51),
.Y(n_283)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_52),
.Y(n_267)
);

MAJx2_ASAP7_75t_L g52 ( 
.A(n_53),
.B(n_58),
.C(n_64),
.Y(n_52)
);

AOI22xp5_ASAP7_75t_L g156 ( 
.A1(n_53),
.A2(n_54),
.B1(n_157),
.B2(n_158),
.Y(n_156)
);

AOI22xp5_ASAP7_75t_L g196 ( 
.A1(n_53),
.A2(n_54),
.B1(n_64),
.B2(n_197),
.Y(n_196)
);

INVx1_ASAP7_75t_SL g53 ( 
.A(n_54),
.Y(n_53)
);

MAJx2_ASAP7_75t_L g437 ( 
.A(n_54),
.B(n_136),
.C(n_159),
.Y(n_437)
);

OR2x2_ASAP7_75t_L g54 ( 
.A(n_55),
.B(n_56),
.Y(n_54)
);

INVx4_ASAP7_75t_L g56 ( 
.A(n_57),
.Y(n_56)
);

INVx3_ASAP7_75t_L g112 ( 
.A(n_57),
.Y(n_112)
);

BUFx6f_ASAP7_75t_L g263 ( 
.A(n_57),
.Y(n_263)
);

XNOR2xp5_ASAP7_75t_L g195 ( 
.A(n_58),
.B(n_196),
.Y(n_195)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_60),
.Y(n_59)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_61),
.Y(n_60)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_62),
.Y(n_61)
);

INVx2_ASAP7_75t_L g128 ( 
.A(n_62),
.Y(n_128)
);

INVx2_ASAP7_75t_L g306 ( 
.A(n_62),
.Y(n_306)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_63),
.Y(n_62)
);

CKINVDCx20_ASAP7_75t_R g197 ( 
.A(n_64),
.Y(n_197)
);

HB1xp67_ASAP7_75t_L g65 ( 
.A(n_66),
.Y(n_65)
);

AOI22xp5_ASAP7_75t_SL g187 ( 
.A1(n_66),
.A2(n_90),
.B1(n_91),
.B2(n_188),
.Y(n_187)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_66),
.Y(n_188)
);

MAJIxp5_ASAP7_75t_L g66 ( 
.A(n_67),
.B(n_79),
.C(n_84),
.Y(n_66)
);

XOR2xp5_ASAP7_75t_SL g224 ( 
.A(n_67),
.B(n_225),
.Y(n_224)
);

MAJIxp5_ASAP7_75t_L g67 ( 
.A(n_68),
.B(n_72),
.C(n_75),
.Y(n_67)
);

AOI22xp5_ASAP7_75t_L g244 ( 
.A1(n_68),
.A2(n_75),
.B1(n_245),
.B2(n_246),
.Y(n_244)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_68),
.Y(n_245)
);

XNOR2xp5_ASAP7_75t_L g301 ( 
.A(n_68),
.B(n_302),
.Y(n_301)
);

BUFx3_ASAP7_75t_L g69 ( 
.A(n_70),
.Y(n_69)
);

BUFx6f_ASAP7_75t_L g349 ( 
.A(n_70),
.Y(n_349)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_71),
.Y(n_70)
);

INVx2_ASAP7_75t_L g125 ( 
.A(n_71),
.Y(n_125)
);

XOR2xp5_ASAP7_75t_L g243 ( 
.A(n_72),
.B(n_244),
.Y(n_243)
);

BUFx6f_ASAP7_75t_L g73 ( 
.A(n_74),
.Y(n_73)
);

BUFx6f_ASAP7_75t_L g154 ( 
.A(n_74),
.Y(n_154)
);

INVxp67_ASAP7_75t_L g246 ( 
.A(n_75),
.Y(n_246)
);

INVx8_ASAP7_75t_L g76 ( 
.A(n_77),
.Y(n_76)
);

INVx3_ASAP7_75t_L g308 ( 
.A(n_77),
.Y(n_308)
);

BUFx6f_ASAP7_75t_L g77 ( 
.A(n_78),
.Y(n_77)
);

AOI22xp5_ASAP7_75t_L g225 ( 
.A1(n_79),
.A2(n_80),
.B1(n_84),
.B2(n_226),
.Y(n_225)
);

INVx1_ASAP7_75t_SL g79 ( 
.A(n_80),
.Y(n_79)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_82),
.Y(n_81)
);

INVx2_ASAP7_75t_L g82 ( 
.A(n_83),
.Y(n_82)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_84),
.Y(n_226)
);

BUFx2_ASAP7_75t_L g85 ( 
.A(n_86),
.Y(n_85)
);

INVx2_ASAP7_75t_L g86 ( 
.A(n_87),
.Y(n_86)
);

INVx2_ASAP7_75t_L g87 ( 
.A(n_88),
.Y(n_87)
);

HB1xp67_ASAP7_75t_L g89 ( 
.A(n_90),
.Y(n_89)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_91),
.Y(n_90)
);

XNOR2xp5_ASAP7_75t_L g91 ( 
.A(n_92),
.B(n_93),
.Y(n_91)
);

MAJx2_ASAP7_75t_L g145 ( 
.A(n_92),
.B(n_94),
.C(n_99),
.Y(n_145)
);

AOI22xp5_ASAP7_75t_L g93 ( 
.A1(n_94),
.A2(n_95),
.B1(n_98),
.B2(n_99),
.Y(n_93)
);

AOI22xp5_ASAP7_75t_L g388 ( 
.A1(n_94),
.A2(n_95),
.B1(n_261),
.B2(n_262),
.Y(n_388)
);

INVx2_ASAP7_75t_SL g94 ( 
.A(n_95),
.Y(n_94)
);

HB1xp67_ASAP7_75t_L g260 ( 
.A(n_95),
.Y(n_260)
);

BUFx6f_ASAP7_75t_L g96 ( 
.A(n_97),
.Y(n_96)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_99),
.Y(n_98)
);

BUFx3_ASAP7_75t_L g100 ( 
.A(n_101),
.Y(n_100)
);

INVx8_ASAP7_75t_L g361 ( 
.A(n_101),
.Y(n_361)
);

AOI22xp5_ASAP7_75t_SL g102 ( 
.A1(n_103),
.A2(n_155),
.B1(n_181),
.B2(n_182),
.Y(n_102)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_103),
.Y(n_181)
);

XNOR2xp5_ASAP7_75t_L g103 ( 
.A(n_104),
.B(n_144),
.Y(n_103)
);

MAJIxp5_ASAP7_75t_SL g407 ( 
.A(n_104),
.B(n_145),
.C(n_408),
.Y(n_407)
);

MAJIxp5_ASAP7_75t_L g104 ( 
.A(n_105),
.B(n_117),
.C(n_129),
.Y(n_104)
);

XNOR2x2_ASAP7_75t_SL g189 ( 
.A(n_105),
.B(n_190),
.Y(n_189)
);

XOR2x1_ASAP7_75t_L g105 ( 
.A(n_106),
.B(n_109),
.Y(n_105)
);

MAJIxp5_ASAP7_75t_L g147 ( 
.A(n_106),
.B(n_110),
.C(n_113),
.Y(n_147)
);

BUFx6f_ASAP7_75t_L g107 ( 
.A(n_108),
.Y(n_107)
);

XNOR2xp5_ASAP7_75t_L g109 ( 
.A(n_110),
.B(n_113),
.Y(n_109)
);

INVx2_ASAP7_75t_L g111 ( 
.A(n_112),
.Y(n_111)
);

HB1xp67_ASAP7_75t_L g114 ( 
.A(n_115),
.Y(n_114)
);

BUFx6f_ASAP7_75t_L g115 ( 
.A(n_116),
.Y(n_115)
);

XNOR2xp5_ASAP7_75t_L g190 ( 
.A(n_117),
.B(n_129),
.Y(n_190)
);

MAJIxp5_ASAP7_75t_L g117 ( 
.A(n_118),
.B(n_122),
.C(n_126),
.Y(n_117)
);

AOI22xp5_ASAP7_75t_L g228 ( 
.A1(n_118),
.A2(n_126),
.B1(n_127),
.B2(n_229),
.Y(n_228)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_118),
.Y(n_229)
);

INVx2_ASAP7_75t_L g119 ( 
.A(n_120),
.Y(n_119)
);

INVx2_ASAP7_75t_L g120 ( 
.A(n_121),
.Y(n_120)
);

INVx3_ASAP7_75t_L g425 ( 
.A(n_121),
.Y(n_425)
);

XOR2xp5_ASAP7_75t_L g227 ( 
.A(n_122),
.B(n_228),
.Y(n_227)
);

INVx2_ASAP7_75t_L g123 ( 
.A(n_124),
.Y(n_123)
);

INVx5_ASAP7_75t_L g124 ( 
.A(n_125),
.Y(n_124)
);

MAJIxp5_ASAP7_75t_L g279 ( 
.A(n_126),
.B(n_280),
.C(n_284),
.Y(n_279)
);

AOI22xp5_ASAP7_75t_L g328 ( 
.A1(n_126),
.A2(n_127),
.B1(n_280),
.B2(n_329),
.Y(n_328)
);

INVx2_ASAP7_75t_SL g126 ( 
.A(n_127),
.Y(n_126)
);

XNOR2xp5_ASAP7_75t_L g129 ( 
.A(n_130),
.B(n_135),
.Y(n_129)
);

MAJIxp5_ASAP7_75t_L g165 ( 
.A(n_130),
.B(n_136),
.C(n_166),
.Y(n_165)
);

INVx3_ASAP7_75t_L g131 ( 
.A(n_132),
.Y(n_131)
);

INVx6_ASAP7_75t_L g132 ( 
.A(n_133),
.Y(n_132)
);

INVx8_ASAP7_75t_L g133 ( 
.A(n_134),
.Y(n_133)
);

AOI22xp5_ASAP7_75t_SL g135 ( 
.A1(n_136),
.A2(n_138),
.B1(n_139),
.B2(n_143),
.Y(n_135)
);

INVx1_ASAP7_75t_SL g143 ( 
.A(n_136),
.Y(n_143)
);

OAI22xp5_ASAP7_75t_SL g158 ( 
.A1(n_136),
.A2(n_143),
.B1(n_159),
.B2(n_163),
.Y(n_158)
);

BUFx3_ASAP7_75t_L g255 ( 
.A(n_137),
.Y(n_255)
);

INVx6_ASAP7_75t_L g354 ( 
.A(n_137),
.Y(n_354)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_139),
.Y(n_138)
);

HB1xp67_ASAP7_75t_L g166 ( 
.A(n_139),
.Y(n_166)
);

INVx2_ASAP7_75t_L g140 ( 
.A(n_141),
.Y(n_140)
);

BUFx6f_ASAP7_75t_L g141 ( 
.A(n_142),
.Y(n_141)
);

XNOR2xp5_ASAP7_75t_L g144 ( 
.A(n_145),
.B(n_146),
.Y(n_144)
);

HB1xp67_ASAP7_75t_L g408 ( 
.A(n_146),
.Y(n_408)
);

XNOR2xp5_ASAP7_75t_L g146 ( 
.A(n_147),
.B(n_148),
.Y(n_146)
);

MAJIxp5_ASAP7_75t_L g440 ( 
.A(n_147),
.B(n_153),
.C(n_441),
.Y(n_440)
);

XNOR2x1_ASAP7_75t_SL g148 ( 
.A(n_149),
.B(n_153),
.Y(n_148)
);

INVx1_ASAP7_75t_L g441 ( 
.A(n_149),
.Y(n_441)
);

INVx4_ASAP7_75t_L g150 ( 
.A(n_151),
.Y(n_150)
);

BUFx6f_ASAP7_75t_L g151 ( 
.A(n_152),
.Y(n_151)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_155),
.Y(n_182)
);

HB1xp67_ASAP7_75t_L g405 ( 
.A(n_155),
.Y(n_405)
);

XOR2xp5_ASAP7_75t_L g155 ( 
.A(n_156),
.B(n_164),
.Y(n_155)
);

MAJIxp5_ASAP7_75t_L g442 ( 
.A(n_156),
.B(n_165),
.C(n_167),
.Y(n_442)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_158),
.Y(n_157)
);

INVx1_ASAP7_75t_SL g163 ( 
.A(n_159),
.Y(n_163)
);

AOI22xp33_ASAP7_75t_L g414 ( 
.A1(n_159),
.A2(n_163),
.B1(n_415),
.B2(n_416),
.Y(n_414)
);

OR2x2_ASAP7_75t_L g159 ( 
.A(n_160),
.B(n_161),
.Y(n_159)
);

OR2x2_ASAP7_75t_L g416 ( 
.A(n_160),
.B(n_417),
.Y(n_416)
);

INVx2_ASAP7_75t_L g320 ( 
.A(n_161),
.Y(n_320)
);

INVx2_ASAP7_75t_L g161 ( 
.A(n_162),
.Y(n_161)
);

BUFx6f_ASAP7_75t_L g368 ( 
.A(n_162),
.Y(n_368)
);

XNOR2xp5_ASAP7_75t_L g164 ( 
.A(n_165),
.B(n_167),
.Y(n_164)
);

XNOR2xp5_ASAP7_75t_L g167 ( 
.A(n_168),
.B(n_172),
.Y(n_167)
);

MAJIxp5_ASAP7_75t_L g421 ( 
.A(n_168),
.B(n_173),
.C(n_177),
.Y(n_421)
);

INVx4_ASAP7_75t_L g169 ( 
.A(n_170),
.Y(n_169)
);

INVx6_ASAP7_75t_L g170 ( 
.A(n_171),
.Y(n_170)
);

XNOR2xp5_ASAP7_75t_L g172 ( 
.A(n_173),
.B(n_177),
.Y(n_172)
);

INVx2_ASAP7_75t_L g174 ( 
.A(n_175),
.Y(n_174)
);

INVx2_ASAP7_75t_L g175 ( 
.A(n_176),
.Y(n_175)
);

INVx2_ASAP7_75t_L g431 ( 
.A(n_176),
.Y(n_431)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_179),
.Y(n_178)
);

INVx6_ASAP7_75t_L g179 ( 
.A(n_180),
.Y(n_179)
);

MAJIxp5_ASAP7_75t_L g403 ( 
.A(n_181),
.B(n_404),
.C(n_405),
.Y(n_403)
);

MAJIxp5_ASAP7_75t_L g183 ( 
.A(n_184),
.B(n_189),
.C(n_191),
.Y(n_183)
);

HB1xp67_ASAP7_75t_L g184 ( 
.A(n_185),
.Y(n_184)
);

AOI22xp5_ASAP7_75t_SL g236 ( 
.A1(n_185),
.A2(n_186),
.B1(n_189),
.B2(n_237),
.Y(n_236)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_186),
.Y(n_185)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_189),
.Y(n_237)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_192),
.Y(n_191)
);

XNOR2xp5_ASAP7_75t_L g235 ( 
.A(n_192),
.B(n_236),
.Y(n_235)
);

MAJIxp5_ASAP7_75t_L g192 ( 
.A(n_193),
.B(n_223),
.C(n_227),
.Y(n_192)
);

XNOR2xp5_ASAP7_75t_L g240 ( 
.A(n_193),
.B(n_241),
.Y(n_240)
);

MAJIxp5_ASAP7_75t_L g193 ( 
.A(n_194),
.B(n_198),
.C(n_206),
.Y(n_193)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_195),
.Y(n_194)
);

XNOR2x1_ASAP7_75t_SL g289 ( 
.A(n_195),
.B(n_290),
.Y(n_289)
);

XNOR2x1_ASAP7_75t_L g290 ( 
.A(n_198),
.B(n_206),
.Y(n_290)
);

NAND2xp5_ASAP7_75t_L g198 ( 
.A(n_199),
.B(n_203),
.Y(n_198)
);

XOR2xp5_ASAP7_75t_L g288 ( 
.A(n_199),
.B(n_203),
.Y(n_288)
);

NOR2xp33_ASAP7_75t_L g199 ( 
.A(n_200),
.B(n_202),
.Y(n_199)
);

INVx2_ASAP7_75t_L g200 ( 
.A(n_201),
.Y(n_200)
);

BUFx3_ASAP7_75t_L g204 ( 
.A(n_205),
.Y(n_204)
);

MAJIxp5_ASAP7_75t_L g206 ( 
.A(n_207),
.B(n_213),
.C(n_218),
.Y(n_206)
);

AOI22xp5_ASAP7_75t_SL g275 ( 
.A1(n_207),
.A2(n_213),
.B1(n_276),
.B2(n_277),
.Y(n_275)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_207),
.Y(n_276)
);

INVx2_ASAP7_75t_L g208 ( 
.A(n_209),
.Y(n_208)
);

INVx2_ASAP7_75t_L g209 ( 
.A(n_210),
.Y(n_209)
);

INVx4_ASAP7_75t_L g210 ( 
.A(n_211),
.Y(n_210)
);

BUFx3_ASAP7_75t_L g211 ( 
.A(n_212),
.Y(n_211)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_213),
.Y(n_277)
);

OAI22xp5_ASAP7_75t_SL g346 ( 
.A1(n_213),
.A2(n_277),
.B1(n_347),
.B2(n_348),
.Y(n_346)
);

MAJIxp5_ASAP7_75t_L g375 ( 
.A(n_213),
.B(n_347),
.C(n_376),
.Y(n_375)
);

INVx2_ASAP7_75t_L g214 ( 
.A(n_215),
.Y(n_214)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_216),
.Y(n_215)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_217),
.Y(n_216)
);

BUFx3_ASAP7_75t_L g419 ( 
.A(n_217),
.Y(n_419)
);

XOR2x1_ASAP7_75t_SL g274 ( 
.A(n_218),
.B(n_275),
.Y(n_274)
);

INVx3_ASAP7_75t_L g219 ( 
.A(n_220),
.Y(n_219)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_221),
.Y(n_220)
);

INVx2_ASAP7_75t_L g221 ( 
.A(n_222),
.Y(n_221)
);

HB1xp67_ASAP7_75t_L g223 ( 
.A(n_224),
.Y(n_223)
);

XNOR2xp5_ASAP7_75t_L g241 ( 
.A(n_224),
.B(n_227),
.Y(n_241)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_231),
.Y(n_230)
);

HB1xp67_ASAP7_75t_L g231 ( 
.A(n_232),
.Y(n_231)
);

NAND2xp5_ASAP7_75t_L g232 ( 
.A(n_233),
.B(n_293),
.Y(n_232)
);

MAJIxp5_ASAP7_75t_L g233 ( 
.A(n_234),
.B(n_238),
.C(n_268),
.Y(n_233)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_235),
.Y(n_234)
);

NAND2xp5_ASAP7_75t_L g295 ( 
.A(n_235),
.B(n_239),
.Y(n_295)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_239),
.Y(n_238)
);

MAJIxp5_ASAP7_75t_L g239 ( 
.A(n_240),
.B(n_242),
.C(n_264),
.Y(n_239)
);

XOR2xp5_ASAP7_75t_L g291 ( 
.A(n_240),
.B(n_292),
.Y(n_291)
);

XNOR2xp5_ASAP7_75t_L g292 ( 
.A(n_242),
.B(n_265),
.Y(n_292)
);

MAJIxp5_ASAP7_75t_L g242 ( 
.A(n_243),
.B(n_247),
.C(n_256),
.Y(n_242)
);

XNOR2xp5_ASAP7_75t_L g271 ( 
.A(n_243),
.B(n_247),
.Y(n_271)
);

MAJIxp5_ASAP7_75t_L g326 ( 
.A(n_245),
.B(n_303),
.C(n_307),
.Y(n_326)
);

INVx6_ASAP7_75t_L g248 ( 
.A(n_249),
.Y(n_248)
);

INVx6_ASAP7_75t_L g249 ( 
.A(n_250),
.Y(n_249)
);

BUFx6f_ASAP7_75t_L g250 ( 
.A(n_251),
.Y(n_250)
);

NOR2xp33_ASAP7_75t_L g252 ( 
.A(n_253),
.B(n_254),
.Y(n_252)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_255),
.Y(n_254)
);

XOR2xp5_ASAP7_75t_L g270 ( 
.A(n_256),
.B(n_271),
.Y(n_270)
);

MAJIxp5_ASAP7_75t_L g256 ( 
.A(n_257),
.B(n_260),
.C(n_261),
.Y(n_256)
);

XNOR2xp5_ASAP7_75t_SL g387 ( 
.A(n_257),
.B(n_388),
.Y(n_387)
);

AND2x2_ASAP7_75t_L g257 ( 
.A(n_258),
.B(n_259),
.Y(n_257)
);

XNOR2x1_ASAP7_75t_SL g333 ( 
.A(n_258),
.B(n_259),
.Y(n_333)
);

CKINVDCx16_ASAP7_75t_R g351 ( 
.A(n_258),
.Y(n_351)
);

AOI22xp5_ASAP7_75t_L g362 ( 
.A1(n_258),
.A2(n_351),
.B1(n_352),
.B2(n_363),
.Y(n_362)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_262),
.Y(n_261)
);

HB1xp67_ASAP7_75t_L g264 ( 
.A(n_265),
.Y(n_264)
);

NOR2x1_ASAP7_75t_L g268 ( 
.A(n_269),
.B(n_291),
.Y(n_268)
);

NAND2xp5_ASAP7_75t_L g294 ( 
.A(n_269),
.B(n_291),
.Y(n_294)
);

MAJIxp5_ASAP7_75t_L g269 ( 
.A(n_270),
.B(n_272),
.C(n_289),
.Y(n_269)
);

XNOR2xp5_ASAP7_75t_L g396 ( 
.A(n_270),
.B(n_397),
.Y(n_396)
);

HB1xp67_ASAP7_75t_L g272 ( 
.A(n_273),
.Y(n_272)
);

XNOR2xp5_ASAP7_75t_L g397 ( 
.A(n_273),
.B(n_289),
.Y(n_397)
);

MAJIxp5_ASAP7_75t_L g273 ( 
.A(n_274),
.B(n_278),
.C(n_287),
.Y(n_273)
);

XOR2x1_ASAP7_75t_L g382 ( 
.A(n_274),
.B(n_383),
.Y(n_382)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_279),
.Y(n_278)
);

XNOR2xp5_ASAP7_75t_L g383 ( 
.A(n_279),
.B(n_288),
.Y(n_383)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_280),
.Y(n_329)
);

INVx2_ASAP7_75t_L g281 ( 
.A(n_282),
.Y(n_281)
);

INVx1_ASAP7_75t_L g413 ( 
.A(n_282),
.Y(n_413)
);

INVx2_ASAP7_75t_L g282 ( 
.A(n_283),
.Y(n_282)
);

XOR2x2_ASAP7_75t_L g327 ( 
.A(n_284),
.B(n_328),
.Y(n_327)
);

BUFx6f_ASAP7_75t_L g285 ( 
.A(n_286),
.Y(n_285)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_288),
.Y(n_287)
);

NAND3xp33_ASAP7_75t_L g293 ( 
.A(n_294),
.B(n_295),
.C(n_296),
.Y(n_293)
);

OAI21xp5_ASAP7_75t_SL g296 ( 
.A1(n_297),
.A2(n_394),
.B(n_398),
.Y(n_296)
);

AOI21xp5_ASAP7_75t_L g297 ( 
.A1(n_298),
.A2(n_379),
.B(n_393),
.Y(n_297)
);

OAI21x1_ASAP7_75t_L g298 ( 
.A1(n_299),
.A2(n_341),
.B(n_378),
.Y(n_298)
);

AND2x2_ASAP7_75t_L g299 ( 
.A(n_300),
.B(n_324),
.Y(n_299)
);

OR2x2_ASAP7_75t_L g378 ( 
.A(n_300),
.B(n_324),
.Y(n_378)
);

MAJIxp5_ASAP7_75t_L g300 ( 
.A(n_301),
.B(n_309),
.C(n_318),
.Y(n_300)
);

XOR2x1_ASAP7_75t_SL g372 ( 
.A(n_301),
.B(n_373),
.Y(n_372)
);

XNOR2xp5_ASAP7_75t_L g302 ( 
.A(n_303),
.B(n_307),
.Y(n_302)
);

INVx2_ASAP7_75t_L g304 ( 
.A(n_305),
.Y(n_304)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_306),
.Y(n_305)
);

AOI22xp5_ASAP7_75t_L g373 ( 
.A1(n_309),
.A2(n_310),
.B1(n_318),
.B2(n_374),
.Y(n_373)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_310),
.Y(n_309)
);

NAND2xp5_ASAP7_75t_L g310 ( 
.A(n_311),
.B(n_317),
.Y(n_310)
);

XNOR2xp5_ASAP7_75t_L g345 ( 
.A(n_311),
.B(n_317),
.Y(n_345)
);

INVx3_ASAP7_75t_L g312 ( 
.A(n_313),
.Y(n_312)
);

INVx2_ASAP7_75t_L g313 ( 
.A(n_314),
.Y(n_313)
);

INVx2_ASAP7_75t_L g314 ( 
.A(n_315),
.Y(n_314)
);

INVx3_ASAP7_75t_L g315 ( 
.A(n_316),
.Y(n_315)
);

INVx1_ASAP7_75t_L g374 ( 
.A(n_318),
.Y(n_374)
);

AO22x1_ASAP7_75t_SL g318 ( 
.A1(n_319),
.A2(n_321),
.B1(n_322),
.B2(n_323),
.Y(n_318)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_319),
.Y(n_322)
);

INVx1_ASAP7_75t_SL g323 ( 
.A(n_321),
.Y(n_323)
);

NAND2xp5_ASAP7_75t_L g331 ( 
.A(n_321),
.B(n_322),
.Y(n_331)
);

NOR2xp33_ASAP7_75t_L g364 ( 
.A(n_323),
.B(n_365),
.Y(n_364)
);

XOR2xp5_ASAP7_75t_L g324 ( 
.A(n_325),
.B(n_330),
.Y(n_324)
);

XNOR2xp5_ASAP7_75t_L g325 ( 
.A(n_326),
.B(n_327),
.Y(n_325)
);

MAJIxp5_ASAP7_75t_L g391 ( 
.A(n_326),
.B(n_327),
.C(n_392),
.Y(n_391)
);

HB1xp67_ASAP7_75t_L g392 ( 
.A(n_330),
.Y(n_392)
);

XOR2xp5_ASAP7_75t_L g330 ( 
.A(n_331),
.B(n_332),
.Y(n_330)
);

MAJx2_ASAP7_75t_L g390 ( 
.A(n_331),
.B(n_333),
.C(n_334),
.Y(n_390)
);

XNOR2xp5_ASAP7_75t_L g332 ( 
.A(n_333),
.B(n_334),
.Y(n_332)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_336),
.Y(n_335)
);

HB1xp67_ASAP7_75t_L g336 ( 
.A(n_337),
.Y(n_336)
);

INVx4_ASAP7_75t_L g337 ( 
.A(n_338),
.Y(n_337)
);

INVx3_ASAP7_75t_L g338 ( 
.A(n_339),
.Y(n_338)
);

INVx6_ASAP7_75t_L g339 ( 
.A(n_340),
.Y(n_339)
);

AOI21x1_ASAP7_75t_L g341 ( 
.A1(n_342),
.A2(n_371),
.B(n_377),
.Y(n_341)
);

OAI21x1_ASAP7_75t_SL g342 ( 
.A1(n_343),
.A2(n_355),
.B(n_370),
.Y(n_342)
);

NOR2xp67_ASAP7_75t_SL g343 ( 
.A(n_344),
.B(n_350),
.Y(n_343)
);

NAND2xp5_ASAP7_75t_L g370 ( 
.A(n_344),
.B(n_350),
.Y(n_370)
);

XNOR2xp5_ASAP7_75t_L g344 ( 
.A(n_345),
.B(n_346),
.Y(n_344)
);

INVx1_ASAP7_75t_L g376 ( 
.A(n_345),
.Y(n_376)
);

INVx1_ASAP7_75t_L g347 ( 
.A(n_348),
.Y(n_347)
);

NOR2xp33_ASAP7_75t_SL g350 ( 
.A(n_351),
.B(n_352),
.Y(n_350)
);

INVx1_ASAP7_75t_L g363 ( 
.A(n_352),
.Y(n_363)
);

INVx6_ASAP7_75t_L g353 ( 
.A(n_354),
.Y(n_353)
);

AOI21xp5_ASAP7_75t_L g355 ( 
.A1(n_356),
.A2(n_364),
.B(n_369),
.Y(n_355)
);

NAND2xp5_ASAP7_75t_L g356 ( 
.A(n_357),
.B(n_362),
.Y(n_356)
);

NOR2xp33_ASAP7_75t_L g369 ( 
.A(n_357),
.B(n_362),
.Y(n_369)
);

INVx1_ASAP7_75t_L g358 ( 
.A(n_359),
.Y(n_358)
);

INVx1_ASAP7_75t_L g359 ( 
.A(n_360),
.Y(n_359)
);

INVx2_ASAP7_75t_L g360 ( 
.A(n_361),
.Y(n_360)
);

INVx1_ASAP7_75t_SL g366 ( 
.A(n_367),
.Y(n_366)
);

INVx1_ASAP7_75t_L g367 ( 
.A(n_368),
.Y(n_367)
);

NAND2xp5_ASAP7_75t_SL g371 ( 
.A(n_372),
.B(n_375),
.Y(n_371)
);

NOR2xp67_ASAP7_75t_L g377 ( 
.A(n_372),
.B(n_375),
.Y(n_377)
);

NAND2xp5_ASAP7_75t_SL g379 ( 
.A(n_380),
.B(n_391),
.Y(n_379)
);

NOR2xp67_ASAP7_75t_L g393 ( 
.A(n_380),
.B(n_391),
.Y(n_393)
);

AOI22xp5_ASAP7_75t_L g380 ( 
.A1(n_381),
.A2(n_382),
.B1(n_384),
.B2(n_385),
.Y(n_380)
);

MAJIxp5_ASAP7_75t_L g395 ( 
.A(n_381),
.B(n_386),
.C(n_390),
.Y(n_395)
);

INVx1_ASAP7_75t_L g381 ( 
.A(n_382),
.Y(n_381)
);

INVx1_ASAP7_75t_L g384 ( 
.A(n_385),
.Y(n_384)
);

AOI22xp5_ASAP7_75t_L g385 ( 
.A1(n_386),
.A2(n_387),
.B1(n_389),
.B2(n_390),
.Y(n_385)
);

INVx1_ASAP7_75t_L g386 ( 
.A(n_387),
.Y(n_386)
);

INVx1_ASAP7_75t_L g389 ( 
.A(n_390),
.Y(n_389)
);

NOR2xp67_ASAP7_75t_L g394 ( 
.A(n_395),
.B(n_396),
.Y(n_394)
);

NAND2xp5_ASAP7_75t_L g398 ( 
.A(n_395),
.B(n_396),
.Y(n_398)
);

NOR2xp33_ASAP7_75t_L g400 ( 
.A(n_401),
.B(n_443),
.Y(n_400)
);

INVxp33_ASAP7_75t_L g401 ( 
.A(n_402),
.Y(n_401)
);

OR2x2_ASAP7_75t_L g402 ( 
.A(n_403),
.B(n_406),
.Y(n_402)
);

AND2x2_ASAP7_75t_L g443 ( 
.A(n_403),
.B(n_406),
.Y(n_443)
);

XOR2xp5_ASAP7_75t_L g406 ( 
.A(n_407),
.B(n_409),
.Y(n_406)
);

XNOR2x1_ASAP7_75t_L g409 ( 
.A(n_410),
.B(n_433),
.Y(n_409)
);

XNOR2xp5_ASAP7_75t_L g410 ( 
.A(n_411),
.B(n_420),
.Y(n_410)
);

XOR2xp5_ASAP7_75t_SL g411 ( 
.A(n_412),
.B(n_414),
.Y(n_411)
);

INVx1_ASAP7_75t_SL g415 ( 
.A(n_416),
.Y(n_415)
);

INVx3_ASAP7_75t_L g417 ( 
.A(n_418),
.Y(n_417)
);

INVx4_ASAP7_75t_L g418 ( 
.A(n_419),
.Y(n_418)
);

XNOR2xp5_ASAP7_75t_L g420 ( 
.A(n_421),
.B(n_422),
.Y(n_420)
);

XOR2xp5_ASAP7_75t_L g422 ( 
.A(n_423),
.B(n_426),
.Y(n_422)
);

INVx3_ASAP7_75t_L g424 ( 
.A(n_425),
.Y(n_424)
);

XNOR2xp5_ASAP7_75t_L g426 ( 
.A(n_427),
.B(n_432),
.Y(n_426)
);

INVx2_ASAP7_75t_L g428 ( 
.A(n_429),
.Y(n_428)
);

INVx2_ASAP7_75t_L g429 ( 
.A(n_430),
.Y(n_429)
);

INVx2_ASAP7_75t_L g430 ( 
.A(n_431),
.Y(n_430)
);

XNOR2x1_ASAP7_75t_L g433 ( 
.A(n_434),
.B(n_442),
.Y(n_433)
);

XNOR2xp5_ASAP7_75t_L g434 ( 
.A(n_435),
.B(n_440),
.Y(n_434)
);

AOI22xp5_ASAP7_75t_L g435 ( 
.A1(n_436),
.A2(n_437),
.B1(n_438),
.B2(n_439),
.Y(n_435)
);

INVx1_ASAP7_75t_L g438 ( 
.A(n_436),
.Y(n_438)
);

INVx1_ASAP7_75t_SL g439 ( 
.A(n_437),
.Y(n_439)
);


endmodule