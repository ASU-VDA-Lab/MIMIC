module real_jpeg_25514_n_5 (n_36, n_4, n_39, n_0, n_37, n_1, n_2, n_38, n_3, n_5);

input n_36;
input n_4;
input n_39;
input n_0;
input n_37;
input n_1;
input n_2;
input n_38;
input n_3;

output n_5;

wire n_17;
wire n_8;
wire n_21;
wire n_33;
wire n_29;
wire n_10;
wire n_31;
wire n_9;
wire n_12;
wire n_24;
wire n_6;
wire n_34;
wire n_28;
wire n_23;
wire n_11;
wire n_14;
wire n_25;
wire n_7;
wire n_22;
wire n_18;
wire n_26;
wire n_32;
wire n_20;
wire n_19;
wire n_27;
wire n_30;
wire n_16;
wire n_15;
wire n_13;

BUFx10_ASAP7_75t_L g12 ( 
.A(n_0),
.Y(n_12)
);

INVx6_ASAP7_75t_SL g27 ( 
.A(n_0),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_1),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g8 ( 
.A(n_2),
.Y(n_8)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_3),
.Y(n_19)
);

NOR2xp33_ASAP7_75t_L g31 ( 
.A(n_4),
.B(n_32),
.Y(n_31)
);

NAND2xp5_ASAP7_75t_SL g34 ( 
.A(n_4),
.B(n_32),
.Y(n_34)
);

XOR2xp5_ASAP7_75t_L g5 ( 
.A(n_6),
.B(n_16),
.Y(n_5)
);

NAND2xp5_ASAP7_75t_SL g6 ( 
.A(n_7),
.B(n_14),
.Y(n_6)
);

NAND2xp5_ASAP7_75t_L g7 ( 
.A(n_8),
.B(n_9),
.Y(n_7)
);

NOR2xp33_ASAP7_75t_SL g15 ( 
.A(n_8),
.B(n_9),
.Y(n_15)
);

OR2x2_ASAP7_75t_L g9 ( 
.A(n_10),
.B(n_13),
.Y(n_9)
);

CKINVDCx20_ASAP7_75t_R g10 ( 
.A(n_11),
.Y(n_10)
);

INVx1_ASAP7_75t_L g11 ( 
.A(n_12),
.Y(n_11)
);

NOR2xp33_ASAP7_75t_SL g21 ( 
.A(n_12),
.B(n_22),
.Y(n_21)
);

NOR2xp33_ASAP7_75t_SL g32 ( 
.A(n_12),
.B(n_33),
.Y(n_32)
);

INVxp67_ASAP7_75t_L g14 ( 
.A(n_15),
.Y(n_14)
);

OAI21xp5_ASAP7_75t_SL g16 ( 
.A1(n_17),
.A2(n_31),
.B(n_34),
.Y(n_16)
);

AOI21xp5_ASAP7_75t_L g17 ( 
.A1(n_18),
.A2(n_23),
.B(n_30),
.Y(n_17)
);

NAND2xp5_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_20),
.Y(n_18)
);

NOR2xp33_ASAP7_75t_SL g30 ( 
.A(n_19),
.B(n_20),
.Y(n_30)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_21),
.Y(n_20)
);

NOR2xp33_ASAP7_75t_SL g23 ( 
.A(n_24),
.B(n_29),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_25),
.Y(n_24)
);

NOR2xp33_ASAP7_75t_SL g25 ( 
.A(n_26),
.B(n_28),
.Y(n_25)
);

INVx8_ASAP7_75t_L g26 ( 
.A(n_27),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g13 ( 
.A(n_36),
.Y(n_13)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_37),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_38),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_39),
.Y(n_33)
);


endmodule