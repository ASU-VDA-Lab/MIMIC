module fake_jpeg_22102_n_319 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_319);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_319;

wire n_253;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVx3_ASAP7_75t_L g17 ( 
.A(n_2),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_15),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_4),
.Y(n_19)
);

INVx5_ASAP7_75t_L g20 ( 
.A(n_13),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_0),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_6),
.Y(n_22)
);

BUFx12f_ASAP7_75t_L g23 ( 
.A(n_5),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_11),
.Y(n_24)
);

BUFx12f_ASAP7_75t_L g25 ( 
.A(n_2),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_7),
.Y(n_26)
);

BUFx5_ASAP7_75t_L g27 ( 
.A(n_4),
.Y(n_27)
);

INVx2_ASAP7_75t_L g28 ( 
.A(n_13),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_5),
.Y(n_29)
);

BUFx12_ASAP7_75t_L g30 ( 
.A(n_11),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_9),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_10),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_1),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_11),
.Y(n_34)
);

INVx2_ASAP7_75t_L g35 ( 
.A(n_30),
.Y(n_35)
);

INVx6_ASAP7_75t_L g56 ( 
.A(n_35),
.Y(n_56)
);

INVx4_ASAP7_75t_L g36 ( 
.A(n_20),
.Y(n_36)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_36),
.Y(n_53)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_23),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_37),
.B(n_39),
.Y(n_50)
);

INVx2_ASAP7_75t_L g38 ( 
.A(n_30),
.Y(n_38)
);

INVx5_ASAP7_75t_L g61 ( 
.A(n_38),
.Y(n_61)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_23),
.Y(n_39)
);

INVx8_ASAP7_75t_L g40 ( 
.A(n_23),
.Y(n_40)
);

INVx2_ASAP7_75t_L g48 ( 
.A(n_40),
.Y(n_48)
);

BUFx4f_ASAP7_75t_SL g41 ( 
.A(n_23),
.Y(n_41)
);

BUFx10_ASAP7_75t_L g46 ( 
.A(n_41),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g42 ( 
.A(n_30),
.B(n_0),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_42),
.B(n_0),
.Y(n_52)
);

BUFx5_ASAP7_75t_L g43 ( 
.A(n_23),
.Y(n_43)
);

BUFx3_ASAP7_75t_L g45 ( 
.A(n_43),
.Y(n_45)
);

AOI22xp33_ASAP7_75t_SL g44 ( 
.A1(n_36),
.A2(n_20),
.B1(n_17),
.B2(n_28),
.Y(n_44)
);

AOI21xp5_ASAP7_75t_L g89 ( 
.A1(n_44),
.A2(n_49),
.B(n_64),
.Y(n_89)
);

OAI22xp5_ASAP7_75t_SL g47 ( 
.A1(n_36),
.A2(n_17),
.B1(n_28),
.B2(n_25),
.Y(n_47)
);

OAI22xp5_ASAP7_75t_L g77 ( 
.A1(n_47),
.A2(n_51),
.B1(n_54),
.B2(n_57),
.Y(n_77)
);

AOI22xp33_ASAP7_75t_SL g49 ( 
.A1(n_36),
.A2(n_20),
.B1(n_17),
.B2(n_28),
.Y(n_49)
);

AOI22xp33_ASAP7_75t_L g51 ( 
.A1(n_40),
.A2(n_25),
.B1(n_27),
.B2(n_42),
.Y(n_51)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_52),
.Y(n_87)
);

AOI22xp33_ASAP7_75t_L g54 ( 
.A1(n_40),
.A2(n_25),
.B1(n_27),
.B2(n_42),
.Y(n_54)
);

INVx4_ASAP7_75t_L g55 ( 
.A(n_41),
.Y(n_55)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_55),
.Y(n_93)
);

OAI22xp5_ASAP7_75t_L g57 ( 
.A1(n_40),
.A2(n_25),
.B1(n_27),
.B2(n_26),
.Y(n_57)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_41),
.Y(n_58)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_58),
.Y(n_94)
);

AOI22xp33_ASAP7_75t_L g59 ( 
.A1(n_40),
.A2(n_25),
.B1(n_26),
.B2(n_21),
.Y(n_59)
);

AOI22xp33_ASAP7_75t_L g73 ( 
.A1(n_59),
.A2(n_62),
.B1(n_22),
.B2(n_31),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_37),
.B(n_32),
.Y(n_60)
);

CKINVDCx20_ASAP7_75t_R g68 ( 
.A(n_60),
.Y(n_68)
);

OAI22xp5_ASAP7_75t_L g62 ( 
.A1(n_35),
.A2(n_26),
.B1(n_21),
.B2(n_22),
.Y(n_62)
);

OA22x2_ASAP7_75t_L g63 ( 
.A1(n_41),
.A2(n_19),
.B1(n_33),
.B2(n_24),
.Y(n_63)
);

AOI22xp33_ASAP7_75t_SL g84 ( 
.A1(n_63),
.A2(n_22),
.B1(n_29),
.B2(n_19),
.Y(n_84)
);

AOI22xp33_ASAP7_75t_SL g64 ( 
.A1(n_41),
.A2(n_32),
.B1(n_31),
.B2(n_21),
.Y(n_64)
);

MAJIxp5_ASAP7_75t_L g65 ( 
.A(n_41),
.B(n_29),
.C(n_34),
.Y(n_65)
);

AOI21xp5_ASAP7_75t_L g92 ( 
.A1(n_65),
.A2(n_52),
.B(n_64),
.Y(n_92)
);

INVx2_ASAP7_75t_SL g66 ( 
.A(n_43),
.Y(n_66)
);

INVx11_ASAP7_75t_L g82 ( 
.A(n_66),
.Y(n_82)
);

NOR4xp25_ASAP7_75t_SL g67 ( 
.A(n_63),
.B(n_43),
.C(n_16),
.D(n_15),
.Y(n_67)
);

OAI21xp5_ASAP7_75t_L g98 ( 
.A1(n_67),
.A2(n_65),
.B(n_63),
.Y(n_98)
);

INVx2_ASAP7_75t_L g69 ( 
.A(n_45),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g122 ( 
.A(n_69),
.B(n_70),
.Y(n_122)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_45),
.Y(n_70)
);

INVxp67_ASAP7_75t_L g71 ( 
.A(n_45),
.Y(n_71)
);

INVx1_ASAP7_75t_SL g106 ( 
.A(n_71),
.Y(n_106)
);

CKINVDCx20_ASAP7_75t_R g72 ( 
.A(n_60),
.Y(n_72)
);

CKINVDCx20_ASAP7_75t_R g97 ( 
.A(n_72),
.Y(n_97)
);

OAI22xp5_ASAP7_75t_L g101 ( 
.A1(n_73),
.A2(n_74),
.B1(n_79),
.B2(n_84),
.Y(n_101)
);

AOI22xp33_ASAP7_75t_L g74 ( 
.A1(n_63),
.A2(n_18),
.B1(n_24),
.B2(n_32),
.Y(n_74)
);

CKINVDCx20_ASAP7_75t_R g75 ( 
.A(n_62),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_SL g103 ( 
.A(n_75),
.B(n_47),
.Y(n_103)
);

BUFx6f_ASAP7_75t_L g76 ( 
.A(n_48),
.Y(n_76)
);

CKINVDCx16_ASAP7_75t_R g118 ( 
.A(n_76),
.Y(n_118)
);

INVx4_ASAP7_75t_L g78 ( 
.A(n_61),
.Y(n_78)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_78),
.Y(n_100)
);

AOI22xp33_ASAP7_75t_L g79 ( 
.A1(n_63),
.A2(n_18),
.B1(n_31),
.B2(n_34),
.Y(n_79)
);

INVx3_ASAP7_75t_L g80 ( 
.A(n_57),
.Y(n_80)
);

INVx5_ASAP7_75t_L g111 ( 
.A(n_80),
.Y(n_111)
);

INVx2_ASAP7_75t_L g81 ( 
.A(n_48),
.Y(n_81)
);

INVxp67_ASAP7_75t_L g113 ( 
.A(n_81),
.Y(n_113)
);

INVx4_ASAP7_75t_L g83 ( 
.A(n_61),
.Y(n_83)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_83),
.Y(n_107)
);

BUFx6f_ASAP7_75t_L g85 ( 
.A(n_56),
.Y(n_85)
);

INVx3_ASAP7_75t_L g115 ( 
.A(n_85),
.Y(n_115)
);

AOI22xp33_ASAP7_75t_SL g86 ( 
.A1(n_61),
.A2(n_38),
.B1(n_35),
.B2(n_33),
.Y(n_86)
);

AOI22xp5_ASAP7_75t_SL g112 ( 
.A1(n_86),
.A2(n_90),
.B1(n_66),
.B2(n_53),
.Y(n_112)
);

INVx2_ASAP7_75t_L g88 ( 
.A(n_56),
.Y(n_88)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_88),
.Y(n_109)
);

AOI22xp33_ASAP7_75t_SL g90 ( 
.A1(n_66),
.A2(n_38),
.B1(n_43),
.B2(n_39),
.Y(n_90)
);

HB1xp67_ASAP7_75t_L g91 ( 
.A(n_53),
.Y(n_91)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_91),
.Y(n_110)
);

MAJIxp5_ASAP7_75t_L g99 ( 
.A(n_92),
.B(n_47),
.C(n_58),
.Y(n_99)
);

NOR2x1_ASAP7_75t_L g95 ( 
.A(n_91),
.B(n_63),
.Y(n_95)
);

OAI21xp5_ASAP7_75t_L g150 ( 
.A1(n_95),
.A2(n_103),
.B(n_93),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_L g96 ( 
.A(n_92),
.B(n_65),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g124 ( 
.A(n_96),
.B(n_102),
.Y(n_124)
);

AOI21xp5_ASAP7_75t_SL g147 ( 
.A1(n_98),
.A2(n_101),
.B(n_117),
.Y(n_147)
);

XNOR2xp5_ASAP7_75t_L g143 ( 
.A(n_99),
.B(n_46),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_L g102 ( 
.A(n_87),
.B(n_68),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_L g104 ( 
.A(n_87),
.B(n_72),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_L g132 ( 
.A(n_104),
.B(n_94),
.Y(n_132)
);

OAI22xp5_ASAP7_75t_L g105 ( 
.A1(n_80),
.A2(n_44),
.B1(n_49),
.B2(n_51),
.Y(n_105)
);

OAI22xp5_ASAP7_75t_L g145 ( 
.A1(n_105),
.A2(n_112),
.B1(n_37),
.B2(n_69),
.Y(n_145)
);

OAI22xp5_ASAP7_75t_SL g108 ( 
.A1(n_75),
.A2(n_89),
.B1(n_77),
.B2(n_67),
.Y(n_108)
);

OAI22xp5_ASAP7_75t_SL g128 ( 
.A1(n_108),
.A2(n_117),
.B1(n_77),
.B2(n_68),
.Y(n_128)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_78),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_L g142 ( 
.A(n_114),
.B(n_116),
.Y(n_142)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_78),
.Y(n_116)
);

OA22x2_ASAP7_75t_L g117 ( 
.A1(n_89),
.A2(n_54),
.B1(n_46),
.B2(n_59),
.Y(n_117)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_83),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_SL g125 ( 
.A(n_119),
.B(n_120),
.Y(n_125)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_83),
.Y(n_120)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_81),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_L g130 ( 
.A(n_121),
.B(n_88),
.Y(n_130)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_122),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_L g162 ( 
.A(n_123),
.B(n_126),
.Y(n_162)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_122),
.Y(n_126)
);

CKINVDCx20_ASAP7_75t_R g127 ( 
.A(n_102),
.Y(n_127)
);

CKINVDCx20_ASAP7_75t_R g171 ( 
.A(n_127),
.Y(n_171)
);

AOI22xp5_ASAP7_75t_L g173 ( 
.A1(n_128),
.A2(n_134),
.B1(n_145),
.B2(n_114),
.Y(n_173)
);

AOI21xp5_ASAP7_75t_L g129 ( 
.A1(n_96),
.A2(n_94),
.B(n_55),
.Y(n_129)
);

OAI21xp5_ASAP7_75t_SL g154 ( 
.A1(n_129),
.A2(n_147),
.B(n_150),
.Y(n_154)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_130),
.Y(n_160)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_104),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_L g174 ( 
.A(n_131),
.B(n_133),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_L g155 ( 
.A(n_132),
.B(n_136),
.Y(n_155)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_103),
.Y(n_133)
);

OAI22xp5_ASAP7_75t_SL g134 ( 
.A1(n_111),
.A2(n_56),
.B1(n_55),
.B2(n_39),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_L g135 ( 
.A(n_100),
.B(n_70),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_L g164 ( 
.A(n_135),
.B(n_137),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_L g136 ( 
.A(n_97),
.B(n_50),
.Y(n_136)
);

INVxp67_ASAP7_75t_L g137 ( 
.A(n_112),
.Y(n_137)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_95),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_SL g179 ( 
.A(n_138),
.B(n_141),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_L g139 ( 
.A(n_97),
.B(n_98),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_L g156 ( 
.A(n_139),
.B(n_144),
.Y(n_156)
);

XOR2xp5_ASAP7_75t_L g140 ( 
.A(n_108),
.B(n_50),
.Y(n_140)
);

MAJIxp5_ASAP7_75t_L g153 ( 
.A(n_140),
.B(n_105),
.C(n_110),
.Y(n_153)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_95),
.Y(n_141)
);

XNOR2xp5_ASAP7_75t_L g180 ( 
.A(n_143),
.B(n_144),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_L g144 ( 
.A(n_99),
.B(n_76),
.Y(n_144)
);

XNOR2x1_ASAP7_75t_L g146 ( 
.A(n_117),
.B(n_46),
.Y(n_146)
);

MAJIxp5_ASAP7_75t_SL g175 ( 
.A(n_146),
.B(n_148),
.C(n_149),
.Y(n_175)
);

AND2x2_ASAP7_75t_L g148 ( 
.A(n_117),
.B(n_46),
.Y(n_148)
);

A2O1A1O1Ixp25_ASAP7_75t_L g149 ( 
.A1(n_101),
.A2(n_46),
.B(n_66),
.C(n_85),
.D(n_30),
.Y(n_149)
);

AOI22xp33_ASAP7_75t_L g151 ( 
.A1(n_111),
.A2(n_93),
.B1(n_82),
.B2(n_85),
.Y(n_151)
);

OAI22xp5_ASAP7_75t_L g176 ( 
.A1(n_151),
.A2(n_115),
.B1(n_107),
.B2(n_109),
.Y(n_176)
);

CKINVDCx20_ASAP7_75t_R g152 ( 
.A(n_113),
.Y(n_152)
);

CKINVDCx20_ASAP7_75t_R g172 ( 
.A(n_152),
.Y(n_172)
);

XNOR2xp5_ASAP7_75t_L g184 ( 
.A(n_153),
.B(n_170),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_L g157 ( 
.A(n_127),
.B(n_131),
.Y(n_157)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_157),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_L g158 ( 
.A(n_132),
.B(n_110),
.Y(n_158)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_158),
.Y(n_209)
);

NAND2xp5_ASAP7_75t_L g159 ( 
.A(n_124),
.B(n_133),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_L g187 ( 
.A(n_159),
.B(n_169),
.Y(n_187)
);

OAI22xp5_ASAP7_75t_SL g161 ( 
.A1(n_146),
.A2(n_139),
.B1(n_137),
.B2(n_138),
.Y(n_161)
);

AOI22xp5_ASAP7_75t_L g195 ( 
.A1(n_161),
.A2(n_176),
.B1(n_178),
.B2(n_134),
.Y(n_195)
);

XOR2xp5_ASAP7_75t_L g163 ( 
.A(n_140),
.B(n_117),
.Y(n_163)
);

MAJIxp5_ASAP7_75t_L g194 ( 
.A(n_163),
.B(n_181),
.C(n_182),
.Y(n_194)
);

AOI22xp33_ASAP7_75t_SL g165 ( 
.A1(n_152),
.A2(n_115),
.B1(n_120),
.B2(n_119),
.Y(n_165)
);

CKINVDCx14_ASAP7_75t_R g186 ( 
.A(n_165),
.Y(n_186)
);

NOR2xp33_ASAP7_75t_L g166 ( 
.A(n_142),
.B(n_100),
.Y(n_166)
);

CKINVDCx14_ASAP7_75t_R g204 ( 
.A(n_166),
.Y(n_204)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_142),
.Y(n_167)
);

NOR2xp33_ASAP7_75t_L g188 ( 
.A(n_167),
.B(n_168),
.Y(n_188)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_125),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_L g169 ( 
.A(n_124),
.B(n_121),
.Y(n_169)
);

OAI21xp5_ASAP7_75t_SL g170 ( 
.A1(n_129),
.A2(n_107),
.B(n_116),
.Y(n_170)
);

NOR2xp33_ASAP7_75t_L g205 ( 
.A(n_173),
.B(n_183),
.Y(n_205)
);

NAND2xp5_ASAP7_75t_L g177 ( 
.A(n_136),
.B(n_109),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_L g190 ( 
.A(n_177),
.B(n_123),
.Y(n_190)
);

OAI22xp5_ASAP7_75t_SL g178 ( 
.A1(n_141),
.A2(n_118),
.B1(n_82),
.B2(n_46),
.Y(n_178)
);

XNOR2xp5_ASAP7_75t_SL g197 ( 
.A(n_180),
.B(n_148),
.Y(n_197)
);

MAJIxp5_ASAP7_75t_L g181 ( 
.A(n_128),
.B(n_143),
.C(n_150),
.Y(n_181)
);

XOR2xp5_ASAP7_75t_L g182 ( 
.A(n_147),
.B(n_106),
.Y(n_182)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_125),
.Y(n_183)
);

CKINVDCx16_ASAP7_75t_R g185 ( 
.A(n_162),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_L g213 ( 
.A(n_185),
.B(n_196),
.Y(n_213)
);

INVx5_ASAP7_75t_L g189 ( 
.A(n_160),
.Y(n_189)
);

NOR2xp33_ASAP7_75t_L g217 ( 
.A(n_189),
.B(n_192),
.Y(n_217)
);

NAND2xp5_ASAP7_75t_L g221 ( 
.A(n_190),
.B(n_200),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_L g191 ( 
.A(n_155),
.B(n_126),
.Y(n_191)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_191),
.Y(n_211)
);

NOR3xp33_ASAP7_75t_L g192 ( 
.A(n_171),
.B(n_145),
.C(n_149),
.Y(n_192)
);

OAI21xp5_ASAP7_75t_L g214 ( 
.A1(n_195),
.A2(n_173),
.B(n_164),
.Y(n_214)
);

CKINVDCx16_ASAP7_75t_R g196 ( 
.A(n_162),
.Y(n_196)
);

MAJIxp5_ASAP7_75t_L g215 ( 
.A(n_197),
.B(n_198),
.C(n_199),
.Y(n_215)
);

MAJIxp5_ASAP7_75t_L g198 ( 
.A(n_156),
.B(n_148),
.C(n_106),
.Y(n_198)
);

MAJIxp5_ASAP7_75t_L g199 ( 
.A(n_156),
.B(n_118),
.C(n_76),
.Y(n_199)
);

INVx1_ASAP7_75t_SL g200 ( 
.A(n_179),
.Y(n_200)
);

NOR2xp33_ASAP7_75t_SL g201 ( 
.A(n_167),
.B(n_8),
.Y(n_201)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_201),
.Y(n_212)
);

CKINVDCx20_ASAP7_75t_R g202 ( 
.A(n_172),
.Y(n_202)
);

NAND2xp5_ASAP7_75t_L g230 ( 
.A(n_202),
.B(n_203),
.Y(n_230)
);

NOR3xp33_ASAP7_75t_SL g203 ( 
.A(n_179),
.B(n_171),
.C(n_175),
.Y(n_203)
);

INVx13_ASAP7_75t_L g206 ( 
.A(n_172),
.Y(n_206)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_206),
.Y(n_223)
);

A2O1A1O1Ixp25_ASAP7_75t_L g207 ( 
.A1(n_175),
.A2(n_30),
.B(n_8),
.C(n_9),
.D(n_16),
.Y(n_207)
);

XNOR2xp5_ASAP7_75t_SL g224 ( 
.A(n_207),
.B(n_178),
.Y(n_224)
);

AOI22xp5_ASAP7_75t_L g208 ( 
.A1(n_161),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_208)
);

AOI22xp5_ASAP7_75t_L g234 ( 
.A1(n_208),
.A2(n_176),
.B1(n_168),
.B2(n_183),
.Y(n_234)
);

MAJIxp5_ASAP7_75t_L g210 ( 
.A(n_181),
.B(n_1),
.C(n_2),
.Y(n_210)
);

MAJIxp5_ASAP7_75t_L g219 ( 
.A(n_210),
.B(n_153),
.C(n_163),
.Y(n_219)
);

AOI21xp5_ASAP7_75t_L g248 ( 
.A1(n_214),
.A2(n_228),
.B(n_174),
.Y(n_248)
);

AOI21xp5_ASAP7_75t_L g216 ( 
.A1(n_193),
.A2(n_154),
.B(n_170),
.Y(n_216)
);

OAI21xp5_ASAP7_75t_SL g250 ( 
.A1(n_216),
.A2(n_231),
.B(n_200),
.Y(n_250)
);

INVxp67_ASAP7_75t_L g218 ( 
.A(n_205),
.Y(n_218)
);

NAND2xp5_ASAP7_75t_L g239 ( 
.A(n_218),
.B(n_227),
.Y(n_239)
);

MAJIxp5_ASAP7_75t_L g240 ( 
.A(n_219),
.B(n_222),
.C(n_229),
.Y(n_240)
);

BUFx10_ASAP7_75t_L g220 ( 
.A(n_206),
.Y(n_220)
);

INVx13_ASAP7_75t_L g249 ( 
.A(n_220),
.Y(n_249)
);

MAJIxp5_ASAP7_75t_L g222 ( 
.A(n_194),
.B(n_182),
.C(n_180),
.Y(n_222)
);

AOI22xp5_ASAP7_75t_SL g247 ( 
.A1(n_224),
.A2(n_203),
.B1(n_191),
.B2(n_209),
.Y(n_247)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_188),
.Y(n_225)
);

NAND2xp5_ASAP7_75t_SL g244 ( 
.A(n_225),
.B(n_226),
.Y(n_244)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_190),
.Y(n_226)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_187),
.Y(n_227)
);

AND2x2_ASAP7_75t_L g228 ( 
.A(n_198),
.B(n_157),
.Y(n_228)
);

MAJIxp5_ASAP7_75t_L g229 ( 
.A(n_194),
.B(n_169),
.C(n_159),
.Y(n_229)
);

AOI21xp5_ASAP7_75t_L g231 ( 
.A1(n_193),
.A2(n_154),
.B(n_174),
.Y(n_231)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_187),
.Y(n_232)
);

NAND2xp5_ASAP7_75t_L g252 ( 
.A(n_232),
.B(n_158),
.Y(n_252)
);

INVx3_ASAP7_75t_L g233 ( 
.A(n_189),
.Y(n_233)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_233),
.Y(n_236)
);

OAI22xp5_ASAP7_75t_L g251 ( 
.A1(n_234),
.A2(n_195),
.B1(n_208),
.B2(n_186),
.Y(n_251)
);

XNOR2xp5_ASAP7_75t_L g235 ( 
.A(n_184),
.B(n_155),
.Y(n_235)
);

XNOR2xp5_ASAP7_75t_L g241 ( 
.A(n_235),
.B(n_197),
.Y(n_241)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_221),
.Y(n_237)
);

NAND2xp5_ASAP7_75t_L g268 ( 
.A(n_237),
.B(n_238),
.Y(n_268)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_221),
.Y(n_238)
);

XOR2xp5_ASAP7_75t_L g259 ( 
.A(n_241),
.B(n_246),
.Y(n_259)
);

CKINVDCx20_ASAP7_75t_R g242 ( 
.A(n_213),
.Y(n_242)
);

NOR2xp33_ASAP7_75t_L g267 ( 
.A(n_242),
.B(n_252),
.Y(n_267)
);

MAJIxp5_ASAP7_75t_L g243 ( 
.A(n_222),
.B(n_199),
.C(n_209),
.Y(n_243)
);

MAJIxp5_ASAP7_75t_L g261 ( 
.A(n_243),
.B(n_215),
.C(n_231),
.Y(n_261)
);

BUFx2_ASAP7_75t_L g245 ( 
.A(n_233),
.Y(n_245)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_245),
.Y(n_265)
);

XNOR2xp5_ASAP7_75t_L g246 ( 
.A(n_219),
.B(n_184),
.Y(n_246)
);

OAI22xp5_ASAP7_75t_SL g260 ( 
.A1(n_247),
.A2(n_250),
.B1(n_216),
.B2(n_230),
.Y(n_260)
);

XOR2xp5_ASAP7_75t_L g270 ( 
.A(n_248),
.B(n_224),
.Y(n_270)
);

AOI22xp5_ASAP7_75t_L g257 ( 
.A1(n_251),
.A2(n_255),
.B1(n_211),
.B2(n_228),
.Y(n_257)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_220),
.Y(n_253)
);

AOI22xp5_ASAP7_75t_SL g269 ( 
.A1(n_253),
.A2(n_254),
.B1(n_160),
.B2(n_220),
.Y(n_269)
);

AND2x2_ASAP7_75t_L g254 ( 
.A(n_230),
.B(n_202),
.Y(n_254)
);

OAI22xp5_ASAP7_75t_L g255 ( 
.A1(n_218),
.A2(n_204),
.B1(n_177),
.B2(n_210),
.Y(n_255)
);

OR2x2_ASAP7_75t_L g256 ( 
.A(n_254),
.B(n_217),
.Y(n_256)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_256),
.Y(n_280)
);

OAI22xp5_ASAP7_75t_L g279 ( 
.A1(n_257),
.A2(n_271),
.B1(n_238),
.B2(n_252),
.Y(n_279)
);

XNOR2xp5_ASAP7_75t_L g258 ( 
.A(n_240),
.B(n_229),
.Y(n_258)
);

XNOR2xp5_ASAP7_75t_L g272 ( 
.A(n_258),
.B(n_262),
.Y(n_272)
);

XOR2xp5_ASAP7_75t_L g284 ( 
.A(n_260),
.B(n_264),
.Y(n_284)
);

MAJIxp5_ASAP7_75t_L g277 ( 
.A(n_261),
.B(n_263),
.C(n_239),
.Y(n_277)
);

XNOR2xp5_ASAP7_75t_L g262 ( 
.A(n_240),
.B(n_215),
.Y(n_262)
);

MAJIxp5_ASAP7_75t_L g263 ( 
.A(n_243),
.B(n_223),
.C(n_214),
.Y(n_263)
);

XNOR2xp5_ASAP7_75t_SL g264 ( 
.A(n_248),
.B(n_247),
.Y(n_264)
);

XNOR2xp5_ASAP7_75t_L g266 ( 
.A(n_246),
.B(n_235),
.Y(n_266)
);

XNOR2xp5_ASAP7_75t_L g276 ( 
.A(n_266),
.B(n_239),
.Y(n_276)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_269),
.Y(n_281)
);

XOR2xp5_ASAP7_75t_L g285 ( 
.A(n_270),
.B(n_207),
.Y(n_285)
);

AOI22xp5_ASAP7_75t_L g271 ( 
.A1(n_237),
.A2(n_234),
.B1(n_228),
.B2(n_212),
.Y(n_271)
);

NAND2xp5_ASAP7_75t_L g273 ( 
.A(n_269),
.B(n_220),
.Y(n_273)
);

NAND2xp5_ASAP7_75t_L g287 ( 
.A(n_273),
.B(n_278),
.Y(n_287)
);

MAJx2_ASAP7_75t_L g274 ( 
.A(n_270),
.B(n_241),
.C(n_250),
.Y(n_274)
);

OAI21xp5_ASAP7_75t_SL g295 ( 
.A1(n_274),
.A2(n_275),
.B(n_236),
.Y(n_295)
);

AND2x6_ASAP7_75t_L g275 ( 
.A(n_256),
.B(n_254),
.Y(n_275)
);

XOR2xp5_ASAP7_75t_L g288 ( 
.A(n_276),
.B(n_285),
.Y(n_288)
);

MAJIxp5_ASAP7_75t_L g294 ( 
.A(n_277),
.B(n_259),
.C(n_253),
.Y(n_294)
);

BUFx10_ASAP7_75t_L g278 ( 
.A(n_265),
.Y(n_278)
);

NAND2xp5_ASAP7_75t_L g296 ( 
.A(n_279),
.B(n_282),
.Y(n_296)
);

NOR2xp33_ASAP7_75t_SL g282 ( 
.A(n_267),
.B(n_249),
.Y(n_282)
);

XNOR2xp5_ASAP7_75t_L g283 ( 
.A(n_259),
.B(n_244),
.Y(n_283)
);

NOR2xp33_ASAP7_75t_L g286 ( 
.A(n_283),
.B(n_272),
.Y(n_286)
);

NAND2xp5_ASAP7_75t_SL g302 ( 
.A(n_286),
.B(n_289),
.Y(n_302)
);

NOR2xp33_ASAP7_75t_SL g289 ( 
.A(n_277),
.B(n_263),
.Y(n_289)
);

OAI22xp5_ASAP7_75t_SL g290 ( 
.A1(n_280),
.A2(n_268),
.B1(n_261),
.B2(n_264),
.Y(n_290)
);

NAND2xp5_ASAP7_75t_L g301 ( 
.A(n_290),
.B(n_291),
.Y(n_301)
);

OAI21x1_ASAP7_75t_L g291 ( 
.A1(n_275),
.A2(n_274),
.B(n_284),
.Y(n_291)
);

HB1xp67_ASAP7_75t_L g292 ( 
.A(n_278),
.Y(n_292)
);

NAND2xp5_ASAP7_75t_L g306 ( 
.A(n_292),
.B(n_293),
.Y(n_306)
);

NOR2xp33_ASAP7_75t_L g293 ( 
.A(n_281),
.B(n_249),
.Y(n_293)
);

OAI21xp5_ASAP7_75t_SL g298 ( 
.A1(n_294),
.A2(n_295),
.B(n_287),
.Y(n_298)
);

BUFx24_ASAP7_75t_SL g297 ( 
.A(n_284),
.Y(n_297)
);

XNOR2xp5_ASAP7_75t_L g305 ( 
.A(n_297),
.B(n_8),
.Y(n_305)
);

AOI21xp5_ASAP7_75t_L g309 ( 
.A1(n_298),
.A2(n_300),
.B(n_303),
.Y(n_309)
);

OAI22xp5_ASAP7_75t_SL g299 ( 
.A1(n_296),
.A2(n_285),
.B1(n_236),
.B2(n_278),
.Y(n_299)
);

NOR2xp33_ASAP7_75t_L g307 ( 
.A(n_299),
.B(n_305),
.Y(n_307)
);

NOR2xp33_ASAP7_75t_L g300 ( 
.A(n_294),
.B(n_245),
.Y(n_300)
);

OAI21xp5_ASAP7_75t_SL g303 ( 
.A1(n_288),
.A2(n_9),
.B(n_15),
.Y(n_303)
);

BUFx2_ASAP7_75t_L g304 ( 
.A(n_288),
.Y(n_304)
);

AOI322xp5_ASAP7_75t_L g308 ( 
.A1(n_304),
.A2(n_14),
.A3(n_13),
.B1(n_12),
.B2(n_10),
.C1(n_16),
.C2(n_1),
.Y(n_308)
);

AOI322xp5_ASAP7_75t_L g316 ( 
.A1(n_308),
.A2(n_310),
.A3(n_311),
.B1(n_312),
.B2(n_313),
.C1(n_7),
.C2(n_307),
.Y(n_316)
);

OAI22xp5_ASAP7_75t_L g310 ( 
.A1(n_301),
.A2(n_14),
.B1(n_12),
.B2(n_10),
.Y(n_310)
);

AND2x2_ASAP7_75t_L g311 ( 
.A(n_304),
.B(n_12),
.Y(n_311)
);

AOI322xp5_ASAP7_75t_L g312 ( 
.A1(n_300),
.A2(n_14),
.A3(n_4),
.B1(n_5),
.B2(n_6),
.C1(n_7),
.C2(n_3),
.Y(n_312)
);

AOI322xp5_ASAP7_75t_L g313 ( 
.A1(n_302),
.A2(n_306),
.A3(n_4),
.B1(n_5),
.B2(n_6),
.C1(n_7),
.C2(n_3),
.Y(n_313)
);

OAI21xp5_ASAP7_75t_SL g314 ( 
.A1(n_309),
.A2(n_3),
.B(n_6),
.Y(n_314)
);

NAND2xp5_ASAP7_75t_L g317 ( 
.A(n_314),
.B(n_315),
.Y(n_317)
);

NAND2xp5_ASAP7_75t_L g315 ( 
.A(n_311),
.B(n_3),
.Y(n_315)
);

NOR2xp33_ASAP7_75t_L g318 ( 
.A(n_317),
.B(n_316),
.Y(n_318)
);

BUFx24_ASAP7_75t_SL g319 ( 
.A(n_318),
.Y(n_319)
);


endmodule