module real_jpeg_15835_n_14 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_2, n_13, n_6, n_7, n_3, n_10, n_9, n_14);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_2;
input n_13;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_14;

wire n_384;
wire n_37;
wire n_430;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_460;
wire n_300;
wire n_415;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_446;
wire n_199;
wire n_95;
wire n_441;
wire n_238;
wire n_67;
wire n_350;
wire n_235;
wire n_107;
wire n_369;
wire n_376;
wire n_354;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_355;
wire n_123;
wire n_463;
wire n_425;
wire n_455;
wire n_462;
wire n_50;
wire n_409;
wire n_186;
wire n_137;
wire n_72;
wire n_440;
wire n_171;
wire n_151;
wire n_272;
wire n_461;
wire n_198;
wire n_203;
wire n_23;
wire n_362;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_339;
wire n_326;
wire n_80;
wire n_30;
wire n_332;
wire n_149;
wire n_328;
wire n_366;
wire n_456;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_466;
wire n_353;
wire n_453;
wire n_230;
wire n_417;
wire n_428;
wire n_128;
wire n_202;
wire n_216;
wire n_367;
wire n_127;
wire n_365;
wire n_356;
wire n_423;
wire n_464;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_422;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_348;
wire n_252;
wire n_363;
wire n_310;
wire n_345;
wire n_78;
wire n_83;
wire n_288;
wire n_221;
wire n_393;
wire n_104;
wire n_153;
wire n_443;
wire n_337;
wire n_131;
wire n_439;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_378;
wire n_200;
wire n_432;
wire n_465;
wire n_335;
wire n_214;
wire n_113;
wire n_251;
wire n_459;
wire n_139;
wire n_33;
wire n_175;
wire n_338;
wire n_156;
wire n_387;
wire n_434;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_390;
wire n_77;
wire n_399;
wire n_219;
wire n_372;
wire n_122;
wire n_19;
wire n_262;
wire n_334;
wire n_17;
wire n_383;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_426;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_371;
wire n_410;
wire n_421;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_382;
wire n_411;
wire n_20;
wire n_314;
wire n_278;
wire n_103;
wire n_232;
wire n_448;
wire n_212;
wire n_284;
wire n_402;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_452;
wire n_213;
wire n_25;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_407;
wire n_419;
wire n_386;
wire n_341;
wire n_331;
wire n_49;
wire n_68;
wire n_395;
wire n_146;
wire n_286;
wire n_166;
wire n_176;
wire n_215;
wire n_323;
wire n_312;
wire n_325;
wire n_316;
wire n_307;
wire n_161;
wire n_207;
wire n_431;
wire n_420;
wire n_357;
wire n_237;
wire n_445;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_380;
wire n_414;
wire n_140;
wire n_126;
wire n_342;
wire n_120;
wire n_155;
wire n_412;
wire n_405;
wire n_319;
wire n_93;
wire n_242;
wire n_142;
wire n_397;
wire n_76;
wire n_403;
wire n_79;
wire n_282;
wire n_147;
wire n_359;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_449;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_145;
wire n_18;
wire n_266;
wire n_377;
wire n_109;
wire n_391;
wire n_427;
wire n_401;
wire n_148;
wire n_373;
wire n_396;
wire n_392;
wire n_375;
wire n_196;
wire n_298;
wire n_330;
wire n_450;
wire n_333;
wire n_152;
wire n_270;
wire n_159;
wire n_429;
wire n_347;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_336;
wire n_258;
wire n_458;
wire n_150;
wire n_41;
wire n_74;
wire n_404;
wire n_158;
wire n_204;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_413;
wire n_75;
wire n_346;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_457;
wire n_119;
wire n_283;
wire n_358;
wire n_181;
wire n_256;
wire n_253;
wire n_273;
wire n_16;
wire n_54;
wire n_168;
wire n_38;
wire n_442;
wire n_385;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_349;
wire n_418;
wire n_292;
wire n_343;
wire n_64;
wire n_291;
wire n_236;
wire n_370;
wire n_276;
wire n_374;
wire n_287;
wire n_388;
wire n_174;
wire n_400;
wire n_255;
wire n_243;
wire n_299;
wire n_352;
wire n_56;
wire n_293;
wire n_275;
wire n_381;
wire n_227;
wire n_229;
wire n_454;
wire n_379;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_444;
wire n_360;
wire n_398;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_451;
wire n_45;
wire n_437;
wire n_268;
wire n_42;
wire n_313;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_416;
wire n_143;
wire n_351;
wire n_467;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_406;
wire n_303;
wire n_321;
wire n_100;
wire n_368;
wire n_51;
wire n_205;
wire n_361;
wire n_261;
wire n_86;
wire n_324;
wire n_70;
wire n_435;
wire n_32;
wire n_228;
wire n_389;
wire n_15;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_438;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_394;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_436;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_424;
wire n_468;
wire n_133;
wire n_257;
wire n_447;
wire n_344;
wire n_210;
wire n_206;
wire n_408;
wire n_85;
wire n_96;
wire n_308;
wire n_433;
wire n_364;

AOI21xp5_ASAP7_75t_L g14 ( 
.A1(n_0),
.A2(n_15),
.B(n_467),
.Y(n_14)
);

NOR2xp33_ASAP7_75t_L g467 ( 
.A(n_0),
.B(n_468),
.Y(n_467)
);

INVx2_ASAP7_75t_L g45 ( 
.A(n_1),
.Y(n_45)
);

OAI22xp5_ASAP7_75t_SL g93 ( 
.A1(n_1),
.A2(n_45),
.B1(n_94),
.B2(n_98),
.Y(n_93)
);

AOI22xp5_ASAP7_75t_SL g357 ( 
.A1(n_1),
.A2(n_44),
.B1(n_358),
.B2(n_362),
.Y(n_357)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_2),
.Y(n_109)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_2),
.Y(n_117)
);

BUFx6f_ASAP7_75t_L g80 ( 
.A(n_3),
.Y(n_80)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_3),
.Y(n_83)
);

BUFx5_ASAP7_75t_L g86 ( 
.A(n_3),
.Y(n_86)
);

BUFx5_ASAP7_75t_L g90 ( 
.A(n_3),
.Y(n_90)
);

INVx4_ASAP7_75t_L g60 ( 
.A(n_4),
.Y(n_60)
);

OAI22xp5_ASAP7_75t_SL g186 ( 
.A1(n_4),
.A2(n_60),
.B1(n_187),
.B2(n_190),
.Y(n_186)
);

OAI22xp5_ASAP7_75t_SL g205 ( 
.A1(n_4),
.A2(n_60),
.B1(n_206),
.B2(n_209),
.Y(n_205)
);

AOI22xp5_ASAP7_75t_L g257 ( 
.A1(n_4),
.A2(n_60),
.B1(n_258),
.B2(n_260),
.Y(n_257)
);

AOI22xp5_ASAP7_75t_L g63 ( 
.A1(n_5),
.A2(n_50),
.B1(n_64),
.B2(n_65),
.Y(n_63)
);

INVx1_ASAP7_75t_SL g65 ( 
.A(n_5),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_SL g162 ( 
.A(n_5),
.B(n_132),
.Y(n_162)
);

AOI22xp5_ASAP7_75t_L g178 ( 
.A1(n_5),
.A2(n_65),
.B1(n_179),
.B2(n_181),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_L g197 ( 
.A(n_5),
.B(n_198),
.Y(n_197)
);

OAI22xp5_ASAP7_75t_SL g219 ( 
.A1(n_5),
.A2(n_65),
.B1(n_220),
.B2(n_222),
.Y(n_219)
);

NAND2xp5_ASAP7_75t_L g296 ( 
.A(n_5),
.B(n_126),
.Y(n_296)
);

NAND2xp5_ASAP7_75t_L g319 ( 
.A(n_5),
.B(n_320),
.Y(n_319)
);

NAND2xp5_ASAP7_75t_L g329 ( 
.A(n_5),
.B(n_291),
.Y(n_329)
);

BUFx5_ASAP7_75t_L g203 ( 
.A(n_6),
.Y(n_203)
);

BUFx5_ASAP7_75t_L g215 ( 
.A(n_6),
.Y(n_215)
);

INVx2_ASAP7_75t_L g246 ( 
.A(n_6),
.Y(n_246)
);

INVx3_ASAP7_75t_L g71 ( 
.A(n_7),
.Y(n_71)
);

BUFx3_ASAP7_75t_L g73 ( 
.A(n_7),
.Y(n_73)
);

BUFx6f_ASAP7_75t_L g88 ( 
.A(n_7),
.Y(n_88)
);

BUFx6f_ASAP7_75t_L g121 ( 
.A(n_7),
.Y(n_121)
);

INVx2_ASAP7_75t_L g123 ( 
.A(n_7),
.Y(n_123)
);

BUFx5_ASAP7_75t_L g259 ( 
.A(n_7),
.Y(n_259)
);

BUFx3_ASAP7_75t_L g380 ( 
.A(n_7),
.Y(n_380)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_8),
.Y(n_26)
);

BUFx5_ASAP7_75t_L g29 ( 
.A(n_8),
.Y(n_29)
);

INVx6_ASAP7_75t_L g39 ( 
.A(n_8),
.Y(n_39)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_8),
.Y(n_234)
);

CKINVDCx20_ASAP7_75t_R g468 ( 
.A(n_9),
.Y(n_468)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_10),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g102 ( 
.A(n_10),
.Y(n_102)
);

BUFx6f_ASAP7_75t_L g78 ( 
.A(n_11),
.Y(n_78)
);

BUFx12f_ASAP7_75t_L g208 ( 
.A(n_11),
.Y(n_208)
);

INVx2_ASAP7_75t_L g218 ( 
.A(n_11),
.Y(n_218)
);

BUFx4f_ASAP7_75t_L g369 ( 
.A(n_11),
.Y(n_369)
);

AOI22xp33_ASAP7_75t_SL g47 ( 
.A1(n_12),
.A2(n_48),
.B1(n_50),
.B2(n_53),
.Y(n_47)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_12),
.Y(n_53)
);

OAI22xp33_ASAP7_75t_SL g67 ( 
.A1(n_12),
.A2(n_53),
.B1(n_68),
.B2(n_72),
.Y(n_67)
);

OAI22xp5_ASAP7_75t_L g127 ( 
.A1(n_12),
.A2(n_53),
.B1(n_128),
.B2(n_130),
.Y(n_127)
);

AOI22xp5_ASAP7_75t_L g364 ( 
.A1(n_12),
.A2(n_53),
.B1(n_365),
.B2(n_370),
.Y(n_364)
);

INVx2_ASAP7_75t_L g24 ( 
.A(n_13),
.Y(n_24)
);

BUFx3_ASAP7_75t_L g31 ( 
.A(n_13),
.Y(n_31)
);

BUFx5_ASAP7_75t_L g52 ( 
.A(n_13),
.Y(n_52)
);

BUFx5_ASAP7_75t_L g62 ( 
.A(n_13),
.Y(n_62)
);

XNOR2xp5_ASAP7_75t_L g15 ( 
.A(n_16),
.B(n_145),
.Y(n_15)
);

NAND2xp5_ASAP7_75t_SL g16 ( 
.A(n_17),
.B(n_143),
.Y(n_16)
);

NAND2xp5_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_54),
.Y(n_17)
);

NOR2xp33_ASAP7_75t_L g144 ( 
.A(n_18),
.B(n_54),
.Y(n_144)
);

OAI22xp5_ASAP7_75t_SL g18 ( 
.A1(n_19),
.A2(n_32),
.B1(n_40),
.B2(n_47),
.Y(n_18)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_19),
.Y(n_139)
);

HB1xp67_ASAP7_75t_L g19 ( 
.A(n_20),
.Y(n_19)
);

OA22x2_ASAP7_75t_L g57 ( 
.A1(n_20),
.A2(n_32),
.B1(n_58),
.B2(n_63),
.Y(n_57)
);

OA22x2_ASAP7_75t_L g157 ( 
.A1(n_20),
.A2(n_32),
.B1(n_58),
.B2(n_63),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_SL g408 ( 
.A(n_20),
.B(n_32),
.Y(n_408)
);

OAI21x1_ASAP7_75t_L g20 ( 
.A1(n_21),
.A2(n_27),
.B(n_32),
.Y(n_20)
);

INVxp67_ASAP7_75t_L g240 ( 
.A(n_21),
.Y(n_240)
);

AND2x2_ASAP7_75t_L g21 ( 
.A(n_22),
.B(n_25),
.Y(n_21)
);

INVx6_ASAP7_75t_L g22 ( 
.A(n_23),
.Y(n_22)
);

INVx4_ASAP7_75t_L g49 ( 
.A(n_23),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_24),
.Y(n_23)
);

INVx6_ASAP7_75t_L g25 ( 
.A(n_26),
.Y(n_25)
);

NOR2xp33_ASAP7_75t_L g27 ( 
.A(n_28),
.B(n_30),
.Y(n_27)
);

INVx3_ASAP7_75t_L g28 ( 
.A(n_29),
.Y(n_28)
);

INVx4_ASAP7_75t_L g35 ( 
.A(n_29),
.Y(n_35)
);

BUFx2_ASAP7_75t_L g46 ( 
.A(n_30),
.Y(n_46)
);

INVx5_ASAP7_75t_L g64 ( 
.A(n_30),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_31),
.Y(n_30)
);

BUFx12f_ASAP7_75t_L g42 ( 
.A(n_31),
.Y(n_42)
);

OAI21xp5_ASAP7_75t_L g136 ( 
.A1(n_32),
.A2(n_40),
.B(n_137),
.Y(n_136)
);

INVxp67_ASAP7_75t_L g198 ( 
.A(n_32),
.Y(n_198)
);

OA22x2_ASAP7_75t_L g32 ( 
.A1(n_33),
.A2(n_35),
.B1(n_36),
.B2(n_38),
.Y(n_32)
);

INVx4_ASAP7_75t_L g97 ( 
.A(n_33),
.Y(n_97)
);

BUFx3_ASAP7_75t_L g191 ( 
.A(n_33),
.Y(n_191)
);

BUFx6f_ASAP7_75t_L g237 ( 
.A(n_33),
.Y(n_237)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_34),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_34),
.Y(n_37)
);

INVx2_ASAP7_75t_L g113 ( 
.A(n_34),
.Y(n_113)
);

BUFx6f_ASAP7_75t_L g135 ( 
.A(n_34),
.Y(n_135)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_36),
.Y(n_118)
);

INVx3_ASAP7_75t_L g36 ( 
.A(n_37),
.Y(n_36)
);

INVx4_ASAP7_75t_L g38 ( 
.A(n_39),
.Y(n_38)
);

AOI22xp33_ASAP7_75t_SL g40 ( 
.A1(n_41),
.A2(n_43),
.B1(n_44),
.B2(n_46),
.Y(n_40)
);

INVx3_ASAP7_75t_L g41 ( 
.A(n_42),
.Y(n_41)
);

OAI22xp33_ASAP7_75t_SL g376 ( 
.A1(n_43),
.A2(n_44),
.B1(n_377),
.B2(n_381),
.Y(n_376)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_44),
.Y(n_43)
);

BUFx2_ASAP7_75t_L g44 ( 
.A(n_45),
.Y(n_44)
);

AOI22xp5_ASAP7_75t_L g58 ( 
.A1(n_46),
.A2(n_59),
.B1(n_60),
.B2(n_61),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_L g228 ( 
.A(n_46),
.B(n_65),
.Y(n_228)
);

INVx3_ASAP7_75t_L g48 ( 
.A(n_49),
.Y(n_48)
);

INVx6_ASAP7_75t_L g50 ( 
.A(n_51),
.Y(n_50)
);

INVx4_ASAP7_75t_L g51 ( 
.A(n_52),
.Y(n_51)
);

MAJIxp5_ASAP7_75t_L g54 ( 
.A(n_55),
.B(n_136),
.C(n_140),
.Y(n_54)
);

FAx1_ASAP7_75t_SL g168 ( 
.A(n_55),
.B(n_136),
.CI(n_140),
.CON(n_168),
.SN(n_168)
);

MAJIxp5_ASAP7_75t_L g55 ( 
.A(n_56),
.B(n_66),
.C(n_92),
.Y(n_55)
);

HB1xp67_ASAP7_75t_L g56 ( 
.A(n_57),
.Y(n_56)
);

AOI22xp5_ASAP7_75t_L g150 ( 
.A1(n_57),
.A2(n_151),
.B1(n_152),
.B2(n_153),
.Y(n_150)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_57),
.Y(n_151)
);

OAI22xp5_ASAP7_75t_L g372 ( 
.A1(n_57),
.A2(n_151),
.B1(n_184),
.B2(n_185),
.Y(n_372)
);

MAJIxp5_ASAP7_75t_L g397 ( 
.A(n_57),
.B(n_355),
.C(n_398),
.Y(n_397)
);

MAJIxp5_ASAP7_75t_L g419 ( 
.A(n_57),
.B(n_254),
.C(n_420),
.Y(n_419)
);

OAI22xp5_ASAP7_75t_L g430 ( 
.A1(n_57),
.A2(n_151),
.B1(n_194),
.B2(n_255),
.Y(n_430)
);

INVx2_ASAP7_75t_L g59 ( 
.A(n_60),
.Y(n_59)
);

INVx8_ASAP7_75t_L g61 ( 
.A(n_62),
.Y(n_61)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_63),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_L g163 ( 
.A(n_65),
.B(n_164),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_SL g313 ( 
.A(n_65),
.B(n_314),
.Y(n_313)
);

XOR2xp5_ASAP7_75t_SL g153 ( 
.A(n_66),
.B(n_92),
.Y(n_153)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_66),
.Y(n_159)
);

XNOR2xp5_ASAP7_75t_L g453 ( 
.A(n_66),
.B(n_160),
.Y(n_453)
);

AND2x2_ASAP7_75t_L g66 ( 
.A(n_67),
.B(n_74),
.Y(n_66)
);

AOI22xp5_ASAP7_75t_SL g402 ( 
.A1(n_67),
.A2(n_290),
.B1(n_291),
.B2(n_376),
.Y(n_402)
);

BUFx3_ASAP7_75t_L g68 ( 
.A(n_69),
.Y(n_68)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_70),
.Y(n_69)
);

HB1xp67_ASAP7_75t_L g315 ( 
.A(n_70),
.Y(n_315)
);

BUFx3_ASAP7_75t_L g70 ( 
.A(n_71),
.Y(n_70)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_71),
.Y(n_91)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_71),
.Y(n_183)
);

INVx3_ASAP7_75t_L g260 ( 
.A(n_72),
.Y(n_260)
);

INVx5_ASAP7_75t_L g72 ( 
.A(n_73),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_L g74 ( 
.A(n_75),
.B(n_84),
.Y(n_74)
);

NAND2x1p5_ASAP7_75t_L g84 ( 
.A(n_75),
.B(n_85),
.Y(n_84)
);

AOI21xp5_ASAP7_75t_L g177 ( 
.A1(n_75),
.A2(n_84),
.B(n_178),
.Y(n_177)
);

OA22x2_ASAP7_75t_L g256 ( 
.A1(n_75),
.A2(n_84),
.B1(n_178),
.B2(n_257),
.Y(n_256)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_75),
.Y(n_291)
);

OAI21xp5_ASAP7_75t_SL g374 ( 
.A1(n_75),
.A2(n_375),
.B(n_384),
.Y(n_374)
);

OA22x2_ASAP7_75t_L g75 ( 
.A1(n_76),
.A2(n_79),
.B1(n_81),
.B2(n_82),
.Y(n_75)
);

INVx2_ASAP7_75t_L g76 ( 
.A(n_77),
.Y(n_76)
);

INVx2_ASAP7_75t_L g77 ( 
.A(n_78),
.Y(n_77)
);

INVx2_ASAP7_75t_L g81 ( 
.A(n_78),
.Y(n_81)
);

INVx3_ASAP7_75t_L g327 ( 
.A(n_78),
.Y(n_327)
);

INVx8_ASAP7_75t_L g79 ( 
.A(n_80),
.Y(n_79)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_82),
.Y(n_310)
);

INVx2_ASAP7_75t_L g82 ( 
.A(n_83),
.Y(n_82)
);

INVx2_ASAP7_75t_L g290 ( 
.A(n_84),
.Y(n_290)
);

OAI22xp5_ASAP7_75t_L g85 ( 
.A1(n_86),
.A2(n_87),
.B1(n_89),
.B2(n_91),
.Y(n_85)
);

INVx2_ASAP7_75t_L g87 ( 
.A(n_88),
.Y(n_87)
);

BUFx6f_ASAP7_75t_L g180 ( 
.A(n_88),
.Y(n_180)
);

INVx6_ASAP7_75t_L g275 ( 
.A(n_88),
.Y(n_275)
);

INVx2_ASAP7_75t_L g89 ( 
.A(n_90),
.Y(n_89)
);

AOI22xp5_ASAP7_75t_L g92 ( 
.A1(n_93),
.A2(n_103),
.B1(n_126),
.B2(n_127),
.Y(n_92)
);

AOI22xp5_ASAP7_75t_L g160 ( 
.A1(n_93),
.A2(n_103),
.B1(n_126),
.B2(n_161),
.Y(n_160)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_95),
.Y(n_94)
);

INVx2_ASAP7_75t_L g95 ( 
.A(n_96),
.Y(n_95)
);

INVx2_ASAP7_75t_L g96 ( 
.A(n_97),
.Y(n_96)
);

INVx1_ASAP7_75t_SL g98 ( 
.A(n_99),
.Y(n_98)
);

BUFx3_ASAP7_75t_L g99 ( 
.A(n_100),
.Y(n_99)
);

INVx2_ASAP7_75t_SL g100 ( 
.A(n_101),
.Y(n_100)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_102),
.Y(n_101)
);

BUFx6f_ASAP7_75t_L g129 ( 
.A(n_102),
.Y(n_129)
);

INVx3_ASAP7_75t_L g167 ( 
.A(n_102),
.Y(n_167)
);

INVx1_ASAP7_75t_SL g142 ( 
.A(n_103),
.Y(n_142)
);

AOI22x1_ASAP7_75t_L g185 ( 
.A1(n_103),
.A2(n_126),
.B1(n_161),
.B2(n_186),
.Y(n_185)
);

OAI21xp5_ASAP7_75t_L g395 ( 
.A1(n_103),
.A2(n_126),
.B(n_161),
.Y(n_395)
);

AND2x4_ASAP7_75t_L g103 ( 
.A(n_104),
.B(n_119),
.Y(n_103)
);

OAI22xp5_ASAP7_75t_L g104 ( 
.A1(n_105),
.A2(n_110),
.B1(n_114),
.B2(n_118),
.Y(n_104)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_106),
.Y(n_105)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_107),
.Y(n_106)
);

INVx2_ASAP7_75t_L g120 ( 
.A(n_107),
.Y(n_120)
);

INVx2_ASAP7_75t_L g107 ( 
.A(n_108),
.Y(n_107)
);

BUFx3_ASAP7_75t_L g108 ( 
.A(n_109),
.Y(n_108)
);

BUFx3_ASAP7_75t_L g125 ( 
.A(n_109),
.Y(n_125)
);

INVx2_ASAP7_75t_L g110 ( 
.A(n_111),
.Y(n_110)
);

INVx8_ASAP7_75t_L g111 ( 
.A(n_112),
.Y(n_111)
);

BUFx6f_ASAP7_75t_L g112 ( 
.A(n_113),
.Y(n_112)
);

BUFx6f_ASAP7_75t_L g189 ( 
.A(n_113),
.Y(n_189)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_115),
.Y(n_114)
);

INVx2_ASAP7_75t_L g268 ( 
.A(n_115),
.Y(n_268)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_116),
.Y(n_115)
);

BUFx6f_ASAP7_75t_L g116 ( 
.A(n_117),
.Y(n_116)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_119),
.Y(n_126)
);

NAND2xp33_ASAP7_75t_SL g141 ( 
.A(n_119),
.B(n_142),
.Y(n_141)
);

OA22x2_ASAP7_75t_L g194 ( 
.A1(n_119),
.A2(n_142),
.B1(n_195),
.B2(n_196),
.Y(n_194)
);

OA22x2_ASAP7_75t_SL g119 ( 
.A1(n_120),
.A2(n_121),
.B1(n_122),
.B2(n_124),
.Y(n_119)
);

BUFx3_ASAP7_75t_L g265 ( 
.A(n_121),
.Y(n_265)
);

BUFx12f_ASAP7_75t_L g304 ( 
.A(n_121),
.Y(n_304)
);

INVx4_ASAP7_75t_L g383 ( 
.A(n_121),
.Y(n_383)
);

BUFx6f_ASAP7_75t_L g122 ( 
.A(n_123),
.Y(n_122)
);

INVx4_ASAP7_75t_L g124 ( 
.A(n_125),
.Y(n_124)
);

NAND2xp33_ASAP7_75t_SL g140 ( 
.A(n_127),
.B(n_141),
.Y(n_140)
);

BUFx6f_ASAP7_75t_L g128 ( 
.A(n_129),
.Y(n_128)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_131),
.Y(n_130)
);

INVx2_ASAP7_75t_L g131 ( 
.A(n_132),
.Y(n_131)
);

INVx3_ASAP7_75t_L g132 ( 
.A(n_133),
.Y(n_132)
);

INVx2_ASAP7_75t_L g133 ( 
.A(n_134),
.Y(n_133)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_134),
.Y(n_264)
);

INVx2_ASAP7_75t_L g134 ( 
.A(n_135),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_L g137 ( 
.A(n_138),
.B(n_139),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_L g407 ( 
.A(n_138),
.B(n_408),
.Y(n_407)
);

INVxp67_ASAP7_75t_L g143 ( 
.A(n_144),
.Y(n_143)
);

OAI21xp5_ASAP7_75t_L g145 ( 
.A1(n_146),
.A2(n_169),
.B(n_465),
.Y(n_145)
);

INVxp67_ASAP7_75t_L g146 ( 
.A(n_147),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_SL g147 ( 
.A(n_148),
.B(n_168),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_L g466 ( 
.A(n_148),
.B(n_168),
.Y(n_466)
);

MAJIxp5_ASAP7_75t_L g148 ( 
.A(n_149),
.B(n_154),
.C(n_158),
.Y(n_148)
);

OAI22xp5_ASAP7_75t_SL g450 ( 
.A1(n_149),
.A2(n_150),
.B1(n_154),
.B2(n_155),
.Y(n_450)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_150),
.Y(n_149)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_153),
.Y(n_152)
);

MAJIxp5_ASAP7_75t_L g158 ( 
.A(n_154),
.B(n_159),
.C(n_160),
.Y(n_158)
);

XOR2x1_ASAP7_75t_SL g174 ( 
.A(n_154),
.B(n_175),
.Y(n_174)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_155),
.Y(n_154)
);

MAJIxp5_ASAP7_75t_L g388 ( 
.A(n_155),
.B(n_389),
.C(n_394),
.Y(n_388)
);

XNOR2xp5_ASAP7_75t_L g452 ( 
.A(n_155),
.B(n_453),
.Y(n_452)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_156),
.Y(n_155)
);

OAI22xp5_ASAP7_75t_SL g415 ( 
.A1(n_156),
.A2(n_157),
.B1(n_395),
.B2(n_416),
.Y(n_415)
);

MAJIxp5_ASAP7_75t_L g434 ( 
.A(n_156),
.B(n_177),
.C(n_184),
.Y(n_434)
);

INVx2_ASAP7_75t_L g156 ( 
.A(n_157),
.Y(n_156)
);

XOR2xp5_ASAP7_75t_L g449 ( 
.A(n_158),
.B(n_450),
.Y(n_449)
);

INVxp67_ASAP7_75t_SL g196 ( 
.A(n_161),
.Y(n_196)
);

NAND2xp5_ASAP7_75t_L g161 ( 
.A(n_162),
.B(n_163),
.Y(n_161)
);

OAI32xp33_ASAP7_75t_L g262 ( 
.A1(n_163),
.A2(n_263),
.A3(n_265),
.B1(n_266),
.B2(n_269),
.Y(n_262)
);

INVx2_ASAP7_75t_L g164 ( 
.A(n_165),
.Y(n_164)
);

INVx2_ASAP7_75t_L g165 ( 
.A(n_166),
.Y(n_165)
);

INVx2_ASAP7_75t_L g166 ( 
.A(n_167),
.Y(n_166)
);

BUFx24_ASAP7_75t_SL g469 ( 
.A(n_168),
.Y(n_469)
);

AOI21xp5_ASAP7_75t_L g169 ( 
.A1(n_170),
.A2(n_447),
.B(n_462),
.Y(n_169)
);

AO221x1_ASAP7_75t_L g170 ( 
.A1(n_171),
.A2(n_351),
.B1(n_440),
.B2(n_445),
.C(n_446),
.Y(n_170)
);

OAI21xp5_ASAP7_75t_L g171 ( 
.A1(n_172),
.A2(n_282),
.B(n_350),
.Y(n_171)
);

NOR2xp33_ASAP7_75t_L g172 ( 
.A(n_173),
.B(n_247),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_L g350 ( 
.A(n_173),
.B(n_247),
.Y(n_350)
);

XOR2xp5_ASAP7_75t_L g173 ( 
.A(n_174),
.B(n_192),
.Y(n_173)
);

MAJIxp5_ASAP7_75t_L g436 ( 
.A(n_174),
.B(n_193),
.C(n_225),
.Y(n_436)
);

OAI22xp5_ASAP7_75t_L g175 ( 
.A1(n_176),
.A2(n_177),
.B1(n_184),
.B2(n_185),
.Y(n_175)
);

INVxp67_ASAP7_75t_L g176 ( 
.A(n_177),
.Y(n_176)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_178),
.Y(n_289)
);

INVx4_ASAP7_75t_L g179 ( 
.A(n_180),
.Y(n_179)
);

INVx2_ASAP7_75t_L g181 ( 
.A(n_182),
.Y(n_181)
);

INVx2_ASAP7_75t_L g182 ( 
.A(n_183),
.Y(n_182)
);

AOI22xp5_ASAP7_75t_L g286 ( 
.A1(n_184),
.A2(n_185),
.B1(n_287),
.B2(n_288),
.Y(n_286)
);

HB1xp67_ASAP7_75t_L g344 ( 
.A(n_184),
.Y(n_344)
);

INVx2_ASAP7_75t_L g184 ( 
.A(n_185),
.Y(n_184)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_186),
.Y(n_195)
);

HB1xp67_ASAP7_75t_L g187 ( 
.A(n_188),
.Y(n_187)
);

INVx4_ASAP7_75t_L g188 ( 
.A(n_189),
.Y(n_188)
);

BUFx6f_ASAP7_75t_L g239 ( 
.A(n_189),
.Y(n_239)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_191),
.Y(n_190)
);

XOR2xp5_ASAP7_75t_L g192 ( 
.A(n_193),
.B(n_225),
.Y(n_192)
);

MAJIxp5_ASAP7_75t_L g193 ( 
.A(n_194),
.B(n_197),
.C(n_199),
.Y(n_193)
);

INVx3_ASAP7_75t_L g255 ( 
.A(n_194),
.Y(n_255)
);

AND2x2_ASAP7_75t_L g403 ( 
.A(n_194),
.B(n_402),
.Y(n_403)
);

AOI22xp5_ASAP7_75t_L g251 ( 
.A1(n_197),
.A2(n_199),
.B1(n_252),
.B2(n_253),
.Y(n_251)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_197),
.Y(n_252)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_199),
.Y(n_253)
);

NOR2xp67_ASAP7_75t_SL g317 ( 
.A(n_199),
.B(n_318),
.Y(n_317)
);

OA21x2_ASAP7_75t_L g199 ( 
.A1(n_200),
.A2(n_204),
.B(n_212),
.Y(n_199)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_201),
.Y(n_200)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_202),
.Y(n_201)
);

INVx3_ASAP7_75t_L g202 ( 
.A(n_203),
.Y(n_202)
);

INVxp67_ASAP7_75t_L g204 ( 
.A(n_205),
.Y(n_204)
);

AOI22xp5_ASAP7_75t_L g242 ( 
.A1(n_205),
.A2(n_213),
.B1(n_219),
.B2(n_243),
.Y(n_242)
);

INVx2_ASAP7_75t_L g206 ( 
.A(n_207),
.Y(n_206)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_208),
.Y(n_207)
);

INVx2_ASAP7_75t_L g211 ( 
.A(n_208),
.Y(n_211)
);

INVx5_ASAP7_75t_L g224 ( 
.A(n_208),
.Y(n_224)
);

INVx3_ASAP7_75t_L g308 ( 
.A(n_208),
.Y(n_308)
);

BUFx6f_ASAP7_75t_L g370 ( 
.A(n_208),
.Y(n_370)
);

INVx2_ASAP7_75t_L g209 ( 
.A(n_210),
.Y(n_209)
);

INVx2_ASAP7_75t_L g210 ( 
.A(n_211),
.Y(n_210)
);

OAI21xp5_ASAP7_75t_SL g391 ( 
.A1(n_212),
.A2(n_357),
.B(n_392),
.Y(n_391)
);

NAND2xp5_ASAP7_75t_L g212 ( 
.A(n_213),
.B(n_219),
.Y(n_212)
);

NOR2xp33_ASAP7_75t_L g278 ( 
.A(n_213),
.B(n_279),
.Y(n_278)
);

INVxp67_ASAP7_75t_L g363 ( 
.A(n_213),
.Y(n_363)
);

AND2x2_ASAP7_75t_L g213 ( 
.A(n_214),
.B(n_216),
.Y(n_213)
);

INVx2_ASAP7_75t_L g214 ( 
.A(n_215),
.Y(n_214)
);

BUFx12f_ASAP7_75t_L g393 ( 
.A(n_215),
.Y(n_393)
);

INVx4_ASAP7_75t_L g216 ( 
.A(n_217),
.Y(n_216)
);

BUFx6f_ASAP7_75t_L g221 ( 
.A(n_217),
.Y(n_221)
);

BUFx6f_ASAP7_75t_L g217 ( 
.A(n_218),
.Y(n_217)
);

INVxp33_ASAP7_75t_L g277 ( 
.A(n_219),
.Y(n_277)
);

INVx3_ASAP7_75t_L g220 ( 
.A(n_221),
.Y(n_220)
);

BUFx3_ASAP7_75t_L g312 ( 
.A(n_221),
.Y(n_312)
);

INVx2_ASAP7_75t_L g222 ( 
.A(n_223),
.Y(n_222)
);

INVx3_ASAP7_75t_L g223 ( 
.A(n_224),
.Y(n_223)
);

OAI22xp5_ASAP7_75t_L g225 ( 
.A1(n_226),
.A2(n_227),
.B1(n_241),
.B2(n_242),
.Y(n_225)
);

INVxp67_ASAP7_75t_L g226 ( 
.A(n_227),
.Y(n_226)
);

NAND2xp5_ASAP7_75t_L g420 ( 
.A(n_227),
.B(n_241),
.Y(n_420)
);

OAI22xp5_ASAP7_75t_L g227 ( 
.A1(n_228),
.A2(n_229),
.B1(n_238),
.B2(n_240),
.Y(n_227)
);

NOR2xp33_ASAP7_75t_L g229 ( 
.A(n_230),
.B(n_235),
.Y(n_229)
);

INVx2_ASAP7_75t_L g230 ( 
.A(n_231),
.Y(n_230)
);

INVx2_ASAP7_75t_L g231 ( 
.A(n_232),
.Y(n_231)
);

INVx2_ASAP7_75t_L g232 ( 
.A(n_233),
.Y(n_232)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_234),
.Y(n_233)
);

INVx2_ASAP7_75t_L g235 ( 
.A(n_236),
.Y(n_235)
);

BUFx3_ASAP7_75t_L g236 ( 
.A(n_237),
.Y(n_236)
);

INVx3_ASAP7_75t_L g238 ( 
.A(n_239),
.Y(n_238)
);

AOI22xp5_ASAP7_75t_L g334 ( 
.A1(n_241),
.A2(n_242),
.B1(n_335),
.B2(n_336),
.Y(n_334)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_242),
.Y(n_241)
);

HB1xp67_ASAP7_75t_L g295 ( 
.A(n_242),
.Y(n_295)
);

NAND2xp5_ASAP7_75t_L g328 ( 
.A(n_242),
.B(n_329),
.Y(n_328)
);

NOR2xp33_ASAP7_75t_L g330 ( 
.A(n_242),
.B(n_329),
.Y(n_330)
);

INVx2_ASAP7_75t_L g243 ( 
.A(n_244),
.Y(n_243)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_245),
.Y(n_244)
);

BUFx6f_ASAP7_75t_L g281 ( 
.A(n_245),
.Y(n_281)
);

INVx2_ASAP7_75t_L g245 ( 
.A(n_246),
.Y(n_245)
);

MAJIxp5_ASAP7_75t_L g247 ( 
.A(n_248),
.B(n_256),
.C(n_261),
.Y(n_247)
);

AOI22xp5_ASAP7_75t_L g345 ( 
.A1(n_248),
.A2(n_249),
.B1(n_346),
.B2(n_348),
.Y(n_345)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_249),
.Y(n_248)
);

OAI22xp5_ASAP7_75t_L g249 ( 
.A1(n_250),
.A2(n_251),
.B1(n_254),
.B2(n_255),
.Y(n_249)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_251),
.Y(n_250)
);

NOR2xp67_ASAP7_75t_SL g299 ( 
.A(n_253),
.B(n_300),
.Y(n_299)
);

NAND2xp5_ASAP7_75t_L g331 ( 
.A(n_253),
.B(n_300),
.Y(n_331)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_255),
.Y(n_254)
);

AOI21x1_ASAP7_75t_L g400 ( 
.A1(n_255),
.A2(n_401),
.B(n_403),
.Y(n_400)
);

MAJIxp5_ASAP7_75t_L g294 ( 
.A(n_256),
.B(n_295),
.C(n_296),
.Y(n_294)
);

OAI22xp5_ASAP7_75t_SL g336 ( 
.A1(n_256),
.A2(n_296),
.B1(n_337),
.B2(n_338),
.Y(n_336)
);

INVx2_ASAP7_75t_SL g337 ( 
.A(n_256),
.Y(n_337)
);

OAI22xp5_ASAP7_75t_L g346 ( 
.A1(n_256),
.A2(n_261),
.B1(n_337),
.B2(n_347),
.Y(n_346)
);

OAI22xp5_ASAP7_75t_L g417 ( 
.A1(n_256),
.A2(n_337),
.B1(n_356),
.B2(n_418),
.Y(n_417)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_257),
.Y(n_292)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_259),
.Y(n_258)
);

INVx1_ASAP7_75t_L g347 ( 
.A(n_261),
.Y(n_347)
);

NAND2xp5_ASAP7_75t_L g261 ( 
.A(n_262),
.B(n_276),
.Y(n_261)
);

XOR2xp5_ASAP7_75t_L g293 ( 
.A(n_262),
.B(n_276),
.Y(n_293)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_264),
.Y(n_263)
);

HB1xp67_ASAP7_75t_L g266 ( 
.A(n_267),
.Y(n_266)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_268),
.Y(n_267)
);

HB1xp67_ASAP7_75t_L g270 ( 
.A(n_268),
.Y(n_270)
);

NOR2xp33_ASAP7_75t_L g269 ( 
.A(n_270),
.B(n_271),
.Y(n_269)
);

INVx2_ASAP7_75t_L g271 ( 
.A(n_272),
.Y(n_271)
);

INVx2_ASAP7_75t_L g272 ( 
.A(n_273),
.Y(n_272)
);

INVx2_ASAP7_75t_L g273 ( 
.A(n_274),
.Y(n_273)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_275),
.Y(n_274)
);

NOR2xp33_ASAP7_75t_L g276 ( 
.A(n_277),
.B(n_278),
.Y(n_276)
);

NOR2xp67_ASAP7_75t_SL g386 ( 
.A(n_278),
.B(n_364),
.Y(n_386)
);

INVx2_ASAP7_75t_L g279 ( 
.A(n_280),
.Y(n_279)
);

INVx2_ASAP7_75t_L g280 ( 
.A(n_281),
.Y(n_280)
);

BUFx6f_ASAP7_75t_L g322 ( 
.A(n_281),
.Y(n_322)
);

INVx1_ASAP7_75t_L g371 ( 
.A(n_281),
.Y(n_371)
);

AOI21xp5_ASAP7_75t_L g282 ( 
.A1(n_283),
.A2(n_341),
.B(n_349),
.Y(n_282)
);

OAI21x1_ASAP7_75t_L g283 ( 
.A1(n_284),
.A2(n_297),
.B(n_340),
.Y(n_283)
);

NOR2xp33_ASAP7_75t_L g284 ( 
.A(n_285),
.B(n_294),
.Y(n_284)
);

NAND2xp5_ASAP7_75t_L g340 ( 
.A(n_285),
.B(n_294),
.Y(n_340)
);

XNOR2xp5_ASAP7_75t_L g285 ( 
.A(n_286),
.B(n_293),
.Y(n_285)
);

OAI22xp5_ASAP7_75t_SL g300 ( 
.A1(n_287),
.A2(n_288),
.B1(n_301),
.B2(n_302),
.Y(n_300)
);

OAI22xp5_ASAP7_75t_SL g431 ( 
.A1(n_287),
.A2(n_288),
.B1(n_391),
.B2(n_432),
.Y(n_431)
);

INVx1_ASAP7_75t_SL g287 ( 
.A(n_288),
.Y(n_287)
);

NAND2xp33_ASAP7_75t_R g333 ( 
.A(n_288),
.B(n_302),
.Y(n_333)
);

HB1xp67_ASAP7_75t_L g343 ( 
.A(n_288),
.Y(n_343)
);

AND2x2_ASAP7_75t_L g390 ( 
.A(n_288),
.B(n_391),
.Y(n_390)
);

AO22x2_ASAP7_75t_L g288 ( 
.A1(n_289),
.A2(n_290),
.B1(n_291),
.B2(n_292),
.Y(n_288)
);

NAND2xp5_ASAP7_75t_L g384 ( 
.A(n_289),
.B(n_290),
.Y(n_384)
);

MAJIxp5_ASAP7_75t_L g342 ( 
.A(n_293),
.B(n_343),
.C(n_344),
.Y(n_342)
);

INVx1_ASAP7_75t_L g338 ( 
.A(n_296),
.Y(n_338)
);

AOI21xp5_ASAP7_75t_L g297 ( 
.A1(n_298),
.A2(n_332),
.B(n_339),
.Y(n_297)
);

OAI21xp5_ASAP7_75t_SL g298 ( 
.A1(n_299),
.A2(n_316),
.B(n_331),
.Y(n_298)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_302),
.Y(n_301)
);

OAI32xp33_ASAP7_75t_L g302 ( 
.A1(n_303),
.A2(n_305),
.A3(n_309),
.B1(n_311),
.B2(n_313),
.Y(n_302)
);

INVx2_ASAP7_75t_L g303 ( 
.A(n_304),
.Y(n_303)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_306),
.Y(n_305)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_307),
.Y(n_306)
);

INVx3_ASAP7_75t_L g307 ( 
.A(n_308),
.Y(n_307)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_310),
.Y(n_309)
);

NOR2xp33_ASAP7_75t_L g311 ( 
.A(n_310),
.B(n_312),
.Y(n_311)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_315),
.Y(n_314)
);

AOI21xp5_ASAP7_75t_L g316 ( 
.A1(n_317),
.A2(n_328),
.B(n_330),
.Y(n_316)
);

NAND2xp5_ASAP7_75t_SL g318 ( 
.A(n_319),
.B(n_323),
.Y(n_318)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_321),
.Y(n_320)
);

INVx2_ASAP7_75t_L g321 ( 
.A(n_322),
.Y(n_321)
);

BUFx6f_ASAP7_75t_L g323 ( 
.A(n_324),
.Y(n_323)
);

INVx3_ASAP7_75t_L g324 ( 
.A(n_325),
.Y(n_324)
);

INVx2_ASAP7_75t_L g325 ( 
.A(n_326),
.Y(n_325)
);

BUFx2_ASAP7_75t_L g362 ( 
.A(n_326),
.Y(n_362)
);

INVx2_ASAP7_75t_L g326 ( 
.A(n_327),
.Y(n_326)
);

INVx2_ASAP7_75t_L g361 ( 
.A(n_327),
.Y(n_361)
);

NAND2xp5_ASAP7_75t_L g332 ( 
.A(n_333),
.B(n_334),
.Y(n_332)
);

NOR2xp33_ASAP7_75t_L g339 ( 
.A(n_333),
.B(n_334),
.Y(n_339)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_336),
.Y(n_335)
);

NAND2xp5_ASAP7_75t_SL g355 ( 
.A(n_337),
.B(n_356),
.Y(n_355)
);

NAND2xp5_ASAP7_75t_L g341 ( 
.A(n_342),
.B(n_345),
.Y(n_341)
);

NOR2x1_ASAP7_75t_L g349 ( 
.A(n_342),
.B(n_345),
.Y(n_349)
);

INVx1_ASAP7_75t_L g398 ( 
.A(n_344),
.Y(n_398)
);

INVx1_ASAP7_75t_L g348 ( 
.A(n_346),
.Y(n_348)
);

NOR3xp33_ASAP7_75t_SL g351 ( 
.A(n_352),
.B(n_410),
.C(n_423),
.Y(n_351)
);

INVx1_ASAP7_75t_L g445 ( 
.A(n_352),
.Y(n_445)
);

AND2x2_ASAP7_75t_L g352 ( 
.A(n_353),
.B(n_396),
.Y(n_352)
);

NOR2xp33_ASAP7_75t_L g446 ( 
.A(n_353),
.B(n_396),
.Y(n_446)
);

MAJIxp5_ASAP7_75t_L g353 ( 
.A(n_354),
.B(n_373),
.C(n_388),
.Y(n_353)
);

XOR2xp5_ASAP7_75t_L g422 ( 
.A(n_354),
.B(n_373),
.Y(n_422)
);

XNOR2x1_ASAP7_75t_L g354 ( 
.A(n_355),
.B(n_372),
.Y(n_354)
);

INVxp67_ASAP7_75t_L g418 ( 
.A(n_356),
.Y(n_418)
);

OAI22xp5_ASAP7_75t_SL g356 ( 
.A1(n_357),
.A2(n_363),
.B1(n_364),
.B2(n_371),
.Y(n_356)
);

INVx1_ASAP7_75t_L g358 ( 
.A(n_359),
.Y(n_358)
);

INVx3_ASAP7_75t_L g359 ( 
.A(n_360),
.Y(n_359)
);

INVx2_ASAP7_75t_L g360 ( 
.A(n_361),
.Y(n_360)
);

HB1xp67_ASAP7_75t_L g365 ( 
.A(n_366),
.Y(n_365)
);

INVx2_ASAP7_75t_L g366 ( 
.A(n_367),
.Y(n_366)
);

INVx2_ASAP7_75t_L g367 ( 
.A(n_368),
.Y(n_367)
);

INVx2_ASAP7_75t_L g368 ( 
.A(n_369),
.Y(n_368)
);

OAI22xp5_ASAP7_75t_SL g373 ( 
.A1(n_374),
.A2(n_385),
.B1(n_386),
.B2(n_387),
.Y(n_373)
);

INVxp67_ASAP7_75t_L g387 ( 
.A(n_374),
.Y(n_387)
);

NAND2xp5_ASAP7_75t_L g405 ( 
.A(n_374),
.B(n_386),
.Y(n_405)
);

INVx1_ASAP7_75t_L g375 ( 
.A(n_376),
.Y(n_375)
);

BUFx3_ASAP7_75t_L g377 ( 
.A(n_378),
.Y(n_377)
);

INVx2_ASAP7_75t_L g378 ( 
.A(n_379),
.Y(n_378)
);

INVx3_ASAP7_75t_L g379 ( 
.A(n_380),
.Y(n_379)
);

INVx2_ASAP7_75t_L g381 ( 
.A(n_382),
.Y(n_381)
);

INVx2_ASAP7_75t_L g382 ( 
.A(n_383),
.Y(n_382)
);

OAI22xp5_ASAP7_75t_L g406 ( 
.A1(n_385),
.A2(n_386),
.B1(n_407),
.B2(n_409),
.Y(n_406)
);

INVx1_ASAP7_75t_L g385 ( 
.A(n_386),
.Y(n_385)
);

AOI21xp33_ASAP7_75t_L g455 ( 
.A1(n_386),
.A2(n_405),
.B(n_407),
.Y(n_455)
);

XNOR2xp5_ASAP7_75t_L g421 ( 
.A(n_388),
.B(n_422),
.Y(n_421)
);

INVxp67_ASAP7_75t_L g389 ( 
.A(n_390),
.Y(n_389)
);

XNOR2x1_ASAP7_75t_L g414 ( 
.A(n_390),
.B(n_415),
.Y(n_414)
);

INVx1_ASAP7_75t_L g432 ( 
.A(n_391),
.Y(n_432)
);

INVx6_ASAP7_75t_L g392 ( 
.A(n_393),
.Y(n_392)
);

HB1xp67_ASAP7_75t_L g394 ( 
.A(n_395),
.Y(n_394)
);

INVx1_ASAP7_75t_L g416 ( 
.A(n_395),
.Y(n_416)
);

XNOR2xp5_ASAP7_75t_L g396 ( 
.A(n_397),
.B(n_399),
.Y(n_396)
);

INVx1_ASAP7_75t_L g461 ( 
.A(n_397),
.Y(n_461)
);

XOR2xp5_ASAP7_75t_L g399 ( 
.A(n_400),
.B(n_404),
.Y(n_399)
);

MAJIxp5_ASAP7_75t_L g460 ( 
.A(n_400),
.B(n_404),
.C(n_461),
.Y(n_460)
);

INVxp67_ASAP7_75t_L g401 ( 
.A(n_402),
.Y(n_401)
);

MAJIxp5_ASAP7_75t_L g451 ( 
.A(n_403),
.B(n_452),
.C(n_454),
.Y(n_451)
);

XOR2xp5_ASAP7_75t_L g458 ( 
.A(n_403),
.B(n_452),
.Y(n_458)
);

XOR2xp5_ASAP7_75t_L g404 ( 
.A(n_405),
.B(n_406),
.Y(n_404)
);

INVx1_ASAP7_75t_L g409 ( 
.A(n_407),
.Y(n_409)
);

A2O1A1Ixp33_ASAP7_75t_L g440 ( 
.A1(n_410),
.A2(n_441),
.B(n_442),
.C(n_444),
.Y(n_440)
);

AND2x2_ASAP7_75t_L g410 ( 
.A(n_411),
.B(n_421),
.Y(n_410)
);

OR2x2_ASAP7_75t_L g444 ( 
.A(n_411),
.B(n_421),
.Y(n_444)
);

MAJIxp5_ASAP7_75t_L g411 ( 
.A(n_412),
.B(n_417),
.C(n_419),
.Y(n_411)
);

HB1xp67_ASAP7_75t_L g412 ( 
.A(n_413),
.Y(n_412)
);

OAI22xp5_ASAP7_75t_L g426 ( 
.A1(n_413),
.A2(n_414),
.B1(n_417),
.B2(n_427),
.Y(n_426)
);

INVx2_ASAP7_75t_L g413 ( 
.A(n_414),
.Y(n_413)
);

INVx1_ASAP7_75t_L g427 ( 
.A(n_417),
.Y(n_427)
);

XNOR2xp5_ASAP7_75t_L g425 ( 
.A(n_419),
.B(n_426),
.Y(n_425)
);

XNOR2x1_ASAP7_75t_L g429 ( 
.A(n_420),
.B(n_430),
.Y(n_429)
);

NAND2xp5_ASAP7_75t_SL g423 ( 
.A(n_424),
.B(n_435),
.Y(n_423)
);

NAND2xp5_ASAP7_75t_L g442 ( 
.A(n_424),
.B(n_443),
.Y(n_442)
);

NAND2xp5_ASAP7_75t_SL g424 ( 
.A(n_425),
.B(n_428),
.Y(n_424)
);

OR2x2_ASAP7_75t_L g441 ( 
.A(n_425),
.B(n_428),
.Y(n_441)
);

MAJIxp5_ASAP7_75t_L g428 ( 
.A(n_429),
.B(n_431),
.C(n_433),
.Y(n_428)
);

XNOR2xp5_ASAP7_75t_L g437 ( 
.A(n_429),
.B(n_438),
.Y(n_437)
);

OAI22xp5_ASAP7_75t_SL g438 ( 
.A1(n_431),
.A2(n_433),
.B1(n_434),
.B2(n_439),
.Y(n_438)
);

INVx1_ASAP7_75t_L g439 ( 
.A(n_431),
.Y(n_439)
);

INVx1_ASAP7_75t_L g433 ( 
.A(n_434),
.Y(n_433)
);

NAND2xp5_ASAP7_75t_L g435 ( 
.A(n_436),
.B(n_437),
.Y(n_435)
);

NOR2x1_ASAP7_75t_L g443 ( 
.A(n_436),
.B(n_437),
.Y(n_443)
);

NOR2xp33_ASAP7_75t_L g447 ( 
.A(n_448),
.B(n_456),
.Y(n_447)
);

OAI21xp5_ASAP7_75t_L g462 ( 
.A1(n_448),
.A2(n_463),
.B(n_464),
.Y(n_462)
);

NOR2xp33_ASAP7_75t_L g448 ( 
.A(n_449),
.B(n_451),
.Y(n_448)
);

NAND2xp5_ASAP7_75t_L g464 ( 
.A(n_449),
.B(n_451),
.Y(n_464)
);

OAI22xp5_ASAP7_75t_SL g457 ( 
.A1(n_454),
.A2(n_455),
.B1(n_458),
.B2(n_459),
.Y(n_457)
);

INVx1_ASAP7_75t_L g454 ( 
.A(n_455),
.Y(n_454)
);

NOR2xp33_ASAP7_75t_SL g456 ( 
.A(n_457),
.B(n_460),
.Y(n_456)
);

NAND2xp5_ASAP7_75t_L g463 ( 
.A(n_457),
.B(n_460),
.Y(n_463)
);

INVx1_ASAP7_75t_L g459 ( 
.A(n_458),
.Y(n_459)
);

INVx1_ASAP7_75t_L g465 ( 
.A(n_466),
.Y(n_465)
);


endmodule