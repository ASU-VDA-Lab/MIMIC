module fake_aes_11668_n_39 (n_11, n_1, n_2, n_6, n_4, n_3, n_9, n_5, n_7, n_10, n_8, n_0, n_39);
input n_11;
input n_1;
input n_2;
input n_6;
input n_4;
input n_3;
input n_9;
input n_5;
input n_7;
input n_10;
input n_8;
input n_0;
output n_39;
wire n_20;
wire n_38;
wire n_36;
wire n_37;
wire n_34;
wire n_23;
wire n_28;
wire n_31;
wire n_22;
wire n_25;
wire n_16;
wire n_26;
wire n_13;
wire n_30;
wire n_33;
wire n_18;
wire n_32;
wire n_35;
wire n_12;
wire n_17;
wire n_14;
wire n_15;
wire n_24;
wire n_19;
wire n_21;
wire n_29;
wire n_27;
CKINVDCx5p33_ASAP7_75t_R g12 ( .A(n_10), .Y(n_12) );
CKINVDCx5p33_ASAP7_75t_R g13 ( .A(n_9), .Y(n_13) );
INVx1_ASAP7_75t_L g14 ( .A(n_5), .Y(n_14) );
INVx2_ASAP7_75t_L g15 ( .A(n_0), .Y(n_15) );
NAND2xp5_ASAP7_75t_L g16 ( .A(n_6), .B(n_11), .Y(n_16) );
BUFx6f_ASAP7_75t_L g17 ( .A(n_4), .Y(n_17) );
INVx1_ASAP7_75t_L g18 ( .A(n_15), .Y(n_18) );
INVx1_ASAP7_75t_L g19 ( .A(n_15), .Y(n_19) );
INVx2_ASAP7_75t_L g20 ( .A(n_17), .Y(n_20) );
AND2x4_ASAP7_75t_L g21 ( .A(n_14), .B(n_0), .Y(n_21) );
OAI21x1_ASAP7_75t_L g22 ( .A1(n_20), .A2(n_16), .B(n_12), .Y(n_22) );
AOI22xp33_ASAP7_75t_L g23 ( .A1(n_21), .A2(n_19), .B1(n_18), .B2(n_17), .Y(n_23) );
CKINVDCx5p33_ASAP7_75t_R g24 ( .A(n_23), .Y(n_24) );
HB1xp67_ASAP7_75t_L g25 ( .A(n_22), .Y(n_25) );
NAND2xp5_ASAP7_75t_L g26 ( .A(n_25), .B(n_21), .Y(n_26) );
NAND2xp5_ASAP7_75t_SL g27 ( .A(n_24), .B(n_12), .Y(n_27) );
INVx1_ASAP7_75t_L g28 ( .A(n_26), .Y(n_28) );
AND2x2_ASAP7_75t_L g29 ( .A(n_27), .B(n_25), .Y(n_29) );
AOI222xp33_ASAP7_75t_L g30 ( .A1(n_28), .A2(n_21), .B1(n_17), .B2(n_22), .C1(n_20), .C2(n_13), .Y(n_30) );
OAI322xp33_ASAP7_75t_SL g31 ( .A1(n_28), .A2(n_1), .A3(n_2), .B1(n_3), .B2(n_4), .C1(n_5), .C2(n_17), .Y(n_31) );
NAND2xp33_ASAP7_75t_SL g32 ( .A(n_29), .B(n_17), .Y(n_32) );
INVx2_ASAP7_75t_SL g33 ( .A(n_31), .Y(n_33) );
AND4x2_ASAP7_75t_L g34 ( .A(n_32), .B(n_1), .C(n_2), .D(n_3), .Y(n_34) );
AND4x2_ASAP7_75t_L g35 ( .A(n_30), .B(n_29), .C(n_7), .D(n_8), .Y(n_35) );
AND2x4_ASAP7_75t_L g36 ( .A(n_33), .B(n_34), .Y(n_36) );
BUFx2_ASAP7_75t_L g37 ( .A(n_35), .Y(n_37) );
INVx1_ASAP7_75t_L g38 ( .A(n_36), .Y(n_38) );
AOI22xp5_ASAP7_75t_L g39 ( .A1(n_38), .A2(n_36), .B1(n_37), .B2(n_33), .Y(n_39) );
endmodule