module fake_aes_2917_n_42 (n_1, n_2, n_6, n_4, n_3, n_9, n_5, n_7, n_10, n_8, n_0, n_42);
input n_1;
input n_2;
input n_6;
input n_4;
input n_3;
input n_9;
input n_5;
input n_7;
input n_10;
input n_8;
input n_0;
output n_42;
wire n_20;
wire n_38;
wire n_36;
wire n_37;
wire n_34;
wire n_28;
wire n_23;
wire n_31;
wire n_22;
wire n_11;
wire n_30;
wire n_16;
wire n_26;
wire n_13;
wire n_33;
wire n_25;
wire n_18;
wire n_32;
wire n_41;
wire n_35;
wire n_12;
wire n_17;
wire n_14;
wire n_15;
wire n_24;
wire n_19;
wire n_21;
wire n_29;
wire n_40;
wire n_27;
wire n_39;
BUFx6f_ASAP7_75t_L g11 ( .A(n_2), .Y(n_11) );
INVx2_ASAP7_75t_L g12 ( .A(n_4), .Y(n_12) );
CKINVDCx5p33_ASAP7_75t_R g13 ( .A(n_3), .Y(n_13) );
CKINVDCx5p33_ASAP7_75t_R g14 ( .A(n_4), .Y(n_14) );
CKINVDCx5p33_ASAP7_75t_R g15 ( .A(n_0), .Y(n_15) );
INVx1_ASAP7_75t_L g16 ( .A(n_8), .Y(n_16) );
INVx1_ASAP7_75t_L g17 ( .A(n_10), .Y(n_17) );
INVx1_ASAP7_75t_SL g18 ( .A(n_14), .Y(n_18) );
OR2x6_ASAP7_75t_L g19 ( .A(n_12), .B(n_0), .Y(n_19) );
INVx1_ASAP7_75t_L g20 ( .A(n_12), .Y(n_20) );
AO22x1_ASAP7_75t_L g21 ( .A1(n_14), .A2(n_1), .B1(n_2), .B2(n_3), .Y(n_21) );
BUFx3_ASAP7_75t_L g22 ( .A(n_16), .Y(n_22) );
INVx6_ASAP7_75t_L g23 ( .A(n_11), .Y(n_23) );
AOI221xp5_ASAP7_75t_L g24 ( .A1(n_18), .A2(n_15), .B1(n_13), .B2(n_11), .C(n_17), .Y(n_24) );
O2A1O1Ixp33_ASAP7_75t_L g25 ( .A1(n_20), .A2(n_11), .B(n_5), .C(n_6), .Y(n_25) );
OA21x2_ASAP7_75t_L g26 ( .A1(n_22), .A2(n_9), .B(n_11), .Y(n_26) );
OAI22xp5_ASAP7_75t_L g27 ( .A1(n_19), .A2(n_11), .B1(n_5), .B2(n_6), .Y(n_27) );
NOR2x1_ASAP7_75t_SL g28 ( .A(n_27), .B(n_19), .Y(n_28) );
HB1xp67_ASAP7_75t_L g29 ( .A(n_24), .Y(n_29) );
INVx2_ASAP7_75t_L g30 ( .A(n_26), .Y(n_30) );
INVxp67_ASAP7_75t_SL g31 ( .A(n_28), .Y(n_31) );
INVx1_ASAP7_75t_L g32 ( .A(n_30), .Y(n_32) );
NAND2xp5_ASAP7_75t_L g33 ( .A(n_31), .B(n_29), .Y(n_33) );
AOI21xp5_ASAP7_75t_L g34 ( .A1(n_32), .A2(n_29), .B(n_19), .Y(n_34) );
NOR2xp33_ASAP7_75t_SL g35 ( .A(n_33), .B(n_31), .Y(n_35) );
OAI221xp5_ASAP7_75t_L g36 ( .A1(n_34), .A2(n_19), .B1(n_22), .B2(n_25), .C(n_32), .Y(n_36) );
OR2x2_ASAP7_75t_L g37 ( .A(n_33), .B(n_21), .Y(n_37) );
OAI22xp5_ASAP7_75t_L g38 ( .A1(n_37), .A2(n_32), .B1(n_21), .B2(n_23), .Y(n_38) );
CKINVDCx5p33_ASAP7_75t_R g39 ( .A(n_35), .Y(n_39) );
OAI221xp5_ASAP7_75t_L g40 ( .A1(n_38), .A2(n_36), .B1(n_23), .B2(n_7), .C(n_1), .Y(n_40) );
INVx2_ASAP7_75t_L g41 ( .A(n_39), .Y(n_41) );
AOI22xp5_ASAP7_75t_L g42 ( .A1(n_40), .A2(n_7), .B1(n_23), .B2(n_41), .Y(n_42) );
endmodule