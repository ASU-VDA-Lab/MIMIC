module fake_jpeg_402_n_546 (n_13, n_1, n_10, n_6, n_14, n_18, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_546);

input n_13;
input n_1;
input n_10;
input n_6;
input n_14;
input n_18;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_546;

wire n_529;
wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_525;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_519;
wire n_276;
wire n_143;
wire n_431;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_513;
wire n_283;
wire n_107;
wire n_490;
wire n_517;
wire n_415;
wire n_479;
wire n_543;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_542;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_48;
wire n_465;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_256;
wire n_221;
wire n_454;
wire n_540;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_508;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_544;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_349;
wire n_21;
wire n_288;
wire n_393;
wire n_234;
wire n_530;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_298;
wire n_106;
wire n_545;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_474;
wire n_539;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_511;
wire n_305;
wire n_161;
wire n_441;
wire n_342;
wire n_101;
wire n_226;
wire n_509;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_510;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_536;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_537;
wire n_110;
wire n_531;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_523;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_533;
wire n_296;
wire n_384;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_491;
wire n_24;
wire n_526;
wire n_467;
wire n_269;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_473;
wire n_45;
wire n_520;
wire n_476;
wire n_337;
wire n_317;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_344;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_481;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_522;
wire n_333;
wire n_518;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_302;
wire n_216;
wire n_528;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_199;
wire n_260;
wire n_413;
wire n_275;
wire n_494;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_492;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_515;
wire n_347;
wire n_521;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_538;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_534;
wire n_472;
wire n_279;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_484;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_469;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_527;
wire n_482;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_512;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_516;
wire n_183;
wire n_409;
wire n_532;
wire n_249;
wire n_412;
wire n_217;
wire n_471;
wire n_541;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_535;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_524;
wire n_402;
wire n_504;
wire n_438;
wire n_475;
wire n_247;
wire n_157;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_514;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

NOR2xp33_ASAP7_75t_L g19 ( 
.A(n_16),
.B(n_4),
.Y(n_19)
);

INVx5_ASAP7_75t_L g20 ( 
.A(n_17),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_10),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_0),
.Y(n_22)
);

INVx11_ASAP7_75t_L g23 ( 
.A(n_2),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_15),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_6),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_0),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_10),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_4),
.Y(n_28)
);

INVx1_ASAP7_75t_SL g29 ( 
.A(n_11),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_3),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_5),
.Y(n_31)
);

BUFx3_ASAP7_75t_L g32 ( 
.A(n_18),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_13),
.Y(n_33)
);

INVx11_ASAP7_75t_L g34 ( 
.A(n_11),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_12),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_10),
.Y(n_36)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_11),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_12),
.Y(n_38)
);

INVx1_ASAP7_75t_SL g39 ( 
.A(n_4),
.Y(n_39)
);

BUFx3_ASAP7_75t_L g40 ( 
.A(n_9),
.Y(n_40)
);

BUFx3_ASAP7_75t_L g41 ( 
.A(n_14),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_7),
.Y(n_42)
);

BUFx12f_ASAP7_75t_L g43 ( 
.A(n_15),
.Y(n_43)
);

INVx2_ASAP7_75t_L g44 ( 
.A(n_8),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_15),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_2),
.Y(n_46)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_13),
.Y(n_47)
);

BUFx4f_ASAP7_75t_SL g48 ( 
.A(n_12),
.Y(n_48)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_8),
.Y(n_49)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_14),
.Y(n_50)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_14),
.Y(n_51)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_4),
.Y(n_52)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_0),
.Y(n_53)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_7),
.Y(n_54)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_9),
.Y(n_55)
);

CKINVDCx20_ASAP7_75t_R g56 ( 
.A(n_8),
.Y(n_56)
);

CKINVDCx20_ASAP7_75t_R g57 ( 
.A(n_5),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_SL g58 ( 
.A(n_19),
.B(n_18),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_L g147 ( 
.A(n_58),
.B(n_60),
.Y(n_147)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_21),
.Y(n_59)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_59),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_19),
.B(n_17),
.Y(n_60)
);

NOR3xp33_ASAP7_75t_L g61 ( 
.A(n_29),
.B(n_39),
.C(n_56),
.Y(n_61)
);

NAND3xp33_ASAP7_75t_L g128 ( 
.A(n_61),
.B(n_75),
.C(n_46),
.Y(n_128)
);

AOI22xp5_ASAP7_75t_L g62 ( 
.A1(n_33),
.A2(n_18),
.B1(n_17),
.B2(n_16),
.Y(n_62)
);

OAI22xp5_ASAP7_75t_L g185 ( 
.A1(n_62),
.A2(n_26),
.B1(n_53),
.B2(n_52),
.Y(n_185)
);

BUFx5_ASAP7_75t_L g63 ( 
.A(n_48),
.Y(n_63)
);

INVx2_ASAP7_75t_SL g198 ( 
.A(n_63),
.Y(n_198)
);

INVx6_ASAP7_75t_L g64 ( 
.A(n_25),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g162 ( 
.A(n_64),
.Y(n_162)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_33),
.Y(n_65)
);

BUFx6f_ASAP7_75t_L g166 ( 
.A(n_65),
.Y(n_166)
);

AND2x2_ASAP7_75t_L g66 ( 
.A(n_29),
.B(n_13),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g133 ( 
.A(n_66),
.B(n_74),
.Y(n_133)
);

INVx4_ASAP7_75t_L g67 ( 
.A(n_34),
.Y(n_67)
);

INVx3_ASAP7_75t_L g144 ( 
.A(n_67),
.Y(n_144)
);

INVx4_ASAP7_75t_SL g68 ( 
.A(n_43),
.Y(n_68)
);

CKINVDCx6p67_ASAP7_75t_R g172 ( 
.A(n_68),
.Y(n_172)
);

INVx11_ASAP7_75t_L g69 ( 
.A(n_43),
.Y(n_69)
);

INVx11_ASAP7_75t_L g141 ( 
.A(n_69),
.Y(n_141)
);

INVx5_ASAP7_75t_L g70 ( 
.A(n_20),
.Y(n_70)
);

INVx3_ASAP7_75t_L g152 ( 
.A(n_70),
.Y(n_152)
);

INVx2_ASAP7_75t_L g71 ( 
.A(n_44),
.Y(n_71)
);

INVx2_ASAP7_75t_L g143 ( 
.A(n_71),
.Y(n_143)
);

INVx5_ASAP7_75t_L g72 ( 
.A(n_20),
.Y(n_72)
);

INVx3_ASAP7_75t_L g187 ( 
.A(n_72),
.Y(n_187)
);

INVx2_ASAP7_75t_L g73 ( 
.A(n_44),
.Y(n_73)
);

INVx2_ASAP7_75t_L g168 ( 
.A(n_73),
.Y(n_168)
);

CKINVDCx20_ASAP7_75t_R g74 ( 
.A(n_20),
.Y(n_74)
);

CKINVDCx14_ASAP7_75t_R g75 ( 
.A(n_39),
.Y(n_75)
);

INVx11_ASAP7_75t_L g76 ( 
.A(n_43),
.Y(n_76)
);

INVx11_ASAP7_75t_L g161 ( 
.A(n_76),
.Y(n_161)
);

BUFx6f_ASAP7_75t_L g77 ( 
.A(n_33),
.Y(n_77)
);

BUFx6f_ASAP7_75t_L g174 ( 
.A(n_77),
.Y(n_174)
);

BUFx6f_ASAP7_75t_L g78 ( 
.A(n_33),
.Y(n_78)
);

BUFx6f_ASAP7_75t_L g188 ( 
.A(n_78),
.Y(n_188)
);

INVx3_ASAP7_75t_L g79 ( 
.A(n_43),
.Y(n_79)
);

INVx3_ASAP7_75t_L g206 ( 
.A(n_79),
.Y(n_206)
);

INVx11_ASAP7_75t_L g80 ( 
.A(n_43),
.Y(n_80)
);

INVx4_ASAP7_75t_L g126 ( 
.A(n_80),
.Y(n_126)
);

BUFx5_ASAP7_75t_L g81 ( 
.A(n_48),
.Y(n_81)
);

BUFx5_ASAP7_75t_L g201 ( 
.A(n_81),
.Y(n_201)
);

BUFx3_ASAP7_75t_L g82 ( 
.A(n_25),
.Y(n_82)
);

INVx5_ASAP7_75t_L g129 ( 
.A(n_82),
.Y(n_129)
);

INVx2_ASAP7_75t_L g83 ( 
.A(n_44),
.Y(n_83)
);

INVx2_ASAP7_75t_L g173 ( 
.A(n_83),
.Y(n_173)
);

BUFx6f_ASAP7_75t_L g84 ( 
.A(n_38),
.Y(n_84)
);

INVx6_ASAP7_75t_L g165 ( 
.A(n_84),
.Y(n_165)
);

INVx2_ASAP7_75t_L g85 ( 
.A(n_48),
.Y(n_85)
);

INVx2_ASAP7_75t_L g190 ( 
.A(n_85),
.Y(n_190)
);

BUFx6f_ASAP7_75t_L g86 ( 
.A(n_38),
.Y(n_86)
);

INVx8_ASAP7_75t_L g150 ( 
.A(n_86),
.Y(n_150)
);

BUFx6f_ASAP7_75t_L g87 ( 
.A(n_38),
.Y(n_87)
);

INVx5_ASAP7_75t_L g132 ( 
.A(n_87),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_L g88 ( 
.A(n_24),
.B(n_16),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_L g151 ( 
.A(n_88),
.B(n_90),
.Y(n_151)
);

BUFx6f_ASAP7_75t_L g89 ( 
.A(n_38),
.Y(n_89)
);

INVx5_ASAP7_75t_L g134 ( 
.A(n_89),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_L g90 ( 
.A(n_24),
.B(n_9),
.Y(n_90)
);

BUFx6f_ASAP7_75t_L g91 ( 
.A(n_25),
.Y(n_91)
);

INVx5_ASAP7_75t_L g164 ( 
.A(n_91),
.Y(n_164)
);

BUFx6f_ASAP7_75t_L g92 ( 
.A(n_25),
.Y(n_92)
);

INVx5_ASAP7_75t_L g170 ( 
.A(n_92),
.Y(n_170)
);

INVx3_ASAP7_75t_SL g93 ( 
.A(n_28),
.Y(n_93)
);

INVx2_ASAP7_75t_L g195 ( 
.A(n_93),
.Y(n_195)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_35),
.B(n_0),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_L g160 ( 
.A(n_94),
.B(n_121),
.Y(n_160)
);

BUFx5_ASAP7_75t_L g95 ( 
.A(n_48),
.Y(n_95)
);

INVx4_ASAP7_75t_L g136 ( 
.A(n_95),
.Y(n_136)
);

CKINVDCx9p33_ASAP7_75t_R g96 ( 
.A(n_48),
.Y(n_96)
);

BUFx12f_ASAP7_75t_L g155 ( 
.A(n_96),
.Y(n_155)
);

INVx11_ASAP7_75t_L g97 ( 
.A(n_23),
.Y(n_97)
);

INVx4_ASAP7_75t_L g142 ( 
.A(n_97),
.Y(n_142)
);

INVx3_ASAP7_75t_L g98 ( 
.A(n_32),
.Y(n_98)
);

INVx3_ASAP7_75t_L g135 ( 
.A(n_98),
.Y(n_135)
);

INVx3_ASAP7_75t_L g99 ( 
.A(n_32),
.Y(n_99)
);

INVx3_ASAP7_75t_L g158 ( 
.A(n_99),
.Y(n_158)
);

INVx5_ASAP7_75t_L g100 ( 
.A(n_32),
.Y(n_100)
);

INVx3_ASAP7_75t_L g163 ( 
.A(n_100),
.Y(n_163)
);

INVx8_ASAP7_75t_L g101 ( 
.A(n_28),
.Y(n_101)
);

INVx5_ASAP7_75t_L g194 ( 
.A(n_101),
.Y(n_194)
);

BUFx6f_ASAP7_75t_L g102 ( 
.A(n_28),
.Y(n_102)
);

BUFx12f_ASAP7_75t_L g167 ( 
.A(n_102),
.Y(n_167)
);

INVx2_ASAP7_75t_L g103 ( 
.A(n_22),
.Y(n_103)
);

INVx2_ASAP7_75t_L g196 ( 
.A(n_103),
.Y(n_196)
);

INVx2_ASAP7_75t_L g104 ( 
.A(n_22),
.Y(n_104)
);

INVx2_ASAP7_75t_L g197 ( 
.A(n_104),
.Y(n_197)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_21),
.Y(n_105)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_105),
.Y(n_138)
);

INVx5_ASAP7_75t_L g106 ( 
.A(n_40),
.Y(n_106)
);

INVx2_ASAP7_75t_L g202 ( 
.A(n_106),
.Y(n_202)
);

CKINVDCx16_ASAP7_75t_R g107 ( 
.A(n_28),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_L g148 ( 
.A(n_107),
.B(n_119),
.Y(n_148)
);

BUFx6f_ASAP7_75t_L g108 ( 
.A(n_40),
.Y(n_108)
);

BUFx12f_ASAP7_75t_L g181 ( 
.A(n_108),
.Y(n_181)
);

INVx4_ASAP7_75t_L g109 ( 
.A(n_34),
.Y(n_109)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_109),
.Y(n_146)
);

INVx3_ASAP7_75t_L g110 ( 
.A(n_40),
.Y(n_110)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_110),
.Y(n_203)
);

BUFx12f_ASAP7_75t_L g111 ( 
.A(n_34),
.Y(n_111)
);

BUFx12_ASAP7_75t_L g176 ( 
.A(n_111),
.Y(n_176)
);

HAxp5_ASAP7_75t_SL g112 ( 
.A(n_29),
.B(n_8),
.CON(n_112),
.SN(n_112)
);

AO22x1_ASAP7_75t_L g200 ( 
.A1(n_112),
.A2(n_114),
.B1(n_1),
.B2(n_2),
.Y(n_200)
);

BUFx12f_ASAP7_75t_L g113 ( 
.A(n_39),
.Y(n_113)
);

AND2x2_ASAP7_75t_L g145 ( 
.A(n_113),
.B(n_115),
.Y(n_145)
);

INVx8_ASAP7_75t_L g114 ( 
.A(n_23),
.Y(n_114)
);

INVx4_ASAP7_75t_L g115 ( 
.A(n_23),
.Y(n_115)
);

BUFx6f_ASAP7_75t_L g116 ( 
.A(n_41),
.Y(n_116)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_116),
.Y(n_207)
);

INVx6_ASAP7_75t_L g117 ( 
.A(n_41),
.Y(n_117)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_117),
.Y(n_208)
);

BUFx3_ASAP7_75t_L g118 ( 
.A(n_41),
.Y(n_118)
);

AND2x2_ASAP7_75t_L g178 ( 
.A(n_118),
.B(n_120),
.Y(n_178)
);

OR2x2_ASAP7_75t_L g119 ( 
.A(n_27),
.B(n_1),
.Y(n_119)
);

BUFx3_ASAP7_75t_L g120 ( 
.A(n_27),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_L g121 ( 
.A(n_35),
.B(n_45),
.Y(n_121)
);

BUFx6f_ASAP7_75t_L g122 ( 
.A(n_36),
.Y(n_122)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_122),
.Y(n_209)
);

BUFx6f_ASAP7_75t_L g123 ( 
.A(n_36),
.Y(n_123)
);

CKINVDCx20_ASAP7_75t_R g137 ( 
.A(n_123),
.Y(n_137)
);

INVx5_ASAP7_75t_L g124 ( 
.A(n_45),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_L g157 ( 
.A(n_124),
.B(n_125),
.Y(n_157)
);

INVx4_ASAP7_75t_L g125 ( 
.A(n_26),
.Y(n_125)
);

MAJIxp5_ASAP7_75t_L g127 ( 
.A(n_66),
.B(n_118),
.C(n_119),
.Y(n_127)
);

AND2x2_ASAP7_75t_L g257 ( 
.A(n_127),
.B(n_128),
.Y(n_257)
);

AOI22xp33_ASAP7_75t_SL g131 ( 
.A1(n_68),
.A2(n_113),
.B1(n_109),
.B2(n_111),
.Y(n_131)
);

OA22x2_ASAP7_75t_L g222 ( 
.A1(n_131),
.A2(n_139),
.B1(n_153),
.B2(n_171),
.Y(n_222)
);

AOI22xp33_ASAP7_75t_SL g139 ( 
.A1(n_113),
.A2(n_55),
.B1(n_51),
.B2(n_50),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_SL g140 ( 
.A(n_125),
.B(n_55),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_SL g223 ( 
.A(n_140),
.B(n_149),
.Y(n_223)
);

NOR2xp33_ASAP7_75t_SL g149 ( 
.A(n_120),
.B(n_51),
.Y(n_149)
);

AOI22xp33_ASAP7_75t_SL g153 ( 
.A1(n_111),
.A2(n_50),
.B1(n_47),
.B2(n_37),
.Y(n_153)
);

CKINVDCx20_ASAP7_75t_R g154 ( 
.A(n_122),
.Y(n_154)
);

NOR2xp33_ASAP7_75t_L g217 ( 
.A(n_154),
.B(n_156),
.Y(n_217)
);

CKINVDCx20_ASAP7_75t_R g156 ( 
.A(n_123),
.Y(n_156)
);

NOR2xp33_ASAP7_75t_SL g159 ( 
.A(n_108),
.B(n_37),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_SL g230 ( 
.A(n_159),
.B(n_155),
.Y(n_230)
);

NAND2xp5_ASAP7_75t_L g169 ( 
.A(n_61),
.B(n_47),
.Y(n_169)
);

NOR2xp33_ASAP7_75t_SL g250 ( 
.A(n_169),
.B(n_180),
.Y(n_250)
);

AOI22xp33_ASAP7_75t_SL g171 ( 
.A1(n_112),
.A2(n_31),
.B1(n_56),
.B2(n_54),
.Y(n_171)
);

CKINVDCx20_ASAP7_75t_R g175 ( 
.A(n_64),
.Y(n_175)
);

NOR2xp33_ASAP7_75t_L g221 ( 
.A(n_175),
.B(n_177),
.Y(n_221)
);

NOR2xp33_ASAP7_75t_L g177 ( 
.A(n_75),
.B(n_31),
.Y(n_177)
);

NOR2xp33_ASAP7_75t_L g179 ( 
.A(n_117),
.B(n_57),
.Y(n_179)
);

NOR2xp33_ASAP7_75t_L g235 ( 
.A(n_179),
.B(n_182),
.Y(n_235)
);

NAND2xp5_ASAP7_75t_L g180 ( 
.A(n_93),
.B(n_30),
.Y(n_180)
);

NOR2xp33_ASAP7_75t_L g182 ( 
.A(n_116),
.B(n_57),
.Y(n_182)
);

NOR2xp33_ASAP7_75t_L g183 ( 
.A(n_82),
.B(n_30),
.Y(n_183)
);

NOR2xp33_ASAP7_75t_L g255 ( 
.A(n_183),
.B(n_189),
.Y(n_255)
);

AND2x2_ASAP7_75t_SL g184 ( 
.A(n_65),
.B(n_1),
.Y(n_184)
);

CKINVDCx16_ASAP7_75t_R g239 ( 
.A(n_184),
.Y(n_239)
);

AOI22xp5_ASAP7_75t_L g216 ( 
.A1(n_185),
.A2(n_186),
.B1(n_199),
.B2(n_204),
.Y(n_216)
);

OAI22xp5_ASAP7_75t_L g186 ( 
.A1(n_77),
.A2(n_42),
.B1(n_53),
.B2(n_52),
.Y(n_186)
);

CKINVDCx20_ASAP7_75t_R g189 ( 
.A(n_78),
.Y(n_189)
);

AOI22xp33_ASAP7_75t_SL g191 ( 
.A1(n_114),
.A2(n_54),
.B1(n_49),
.B2(n_46),
.Y(n_191)
);

AOI22xp33_ASAP7_75t_SL g215 ( 
.A1(n_191),
.A2(n_193),
.B1(n_6),
.B2(n_7),
.Y(n_215)
);

NOR2xp33_ASAP7_75t_L g192 ( 
.A(n_101),
.B(n_49),
.Y(n_192)
);

NOR2xp33_ASAP7_75t_L g263 ( 
.A(n_192),
.B(n_205),
.Y(n_263)
);

AOI22xp33_ASAP7_75t_SL g193 ( 
.A1(n_91),
.A2(n_42),
.B1(n_2),
.B2(n_3),
.Y(n_193)
);

OAI22xp33_ASAP7_75t_SL g199 ( 
.A1(n_84),
.A2(n_89),
.B1(n_87),
.B2(n_86),
.Y(n_199)
);

INVx1_ASAP7_75t_SL g251 ( 
.A(n_200),
.Y(n_251)
);

OAI22xp33_ASAP7_75t_SL g204 ( 
.A1(n_92),
.A2(n_1),
.B1(n_3),
.B2(n_5),
.Y(n_204)
);

CKINVDCx20_ASAP7_75t_R g205 ( 
.A(n_102),
.Y(n_205)
);

NOR2xp33_ASAP7_75t_L g210 ( 
.A(n_60),
.B(n_3),
.Y(n_210)
);

NOR2xp33_ASAP7_75t_L g272 ( 
.A(n_210),
.B(n_211),
.Y(n_272)
);

NOR2xp33_ASAP7_75t_L g211 ( 
.A(n_60),
.B(n_5),
.Y(n_211)
);

AOI22xp33_ASAP7_75t_L g212 ( 
.A1(n_96),
.A2(n_6),
.B1(n_7),
.B2(n_91),
.Y(n_212)
);

OAI22xp5_ASAP7_75t_L g273 ( 
.A1(n_212),
.A2(n_166),
.B1(n_174),
.B2(n_188),
.Y(n_273)
);

BUFx12_ASAP7_75t_L g213 ( 
.A(n_172),
.Y(n_213)
);

INVxp67_ASAP7_75t_SL g311 ( 
.A(n_213),
.Y(n_311)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_209),
.Y(n_214)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_214),
.Y(n_288)
);

INVxp67_ASAP7_75t_L g292 ( 
.A(n_215),
.Y(n_292)
);

BUFx3_ASAP7_75t_L g218 ( 
.A(n_172),
.Y(n_218)
);

BUFx3_ASAP7_75t_L g317 ( 
.A(n_218),
.Y(n_317)
);

INVxp67_ASAP7_75t_L g219 ( 
.A(n_145),
.Y(n_219)
);

INVxp67_ASAP7_75t_L g297 ( 
.A(n_219),
.Y(n_297)
);

NAND2xp5_ASAP7_75t_L g220 ( 
.A(n_184),
.B(n_6),
.Y(n_220)
);

NAND2xp5_ASAP7_75t_L g289 ( 
.A(n_220),
.B(n_226),
.Y(n_289)
);

CKINVDCx20_ASAP7_75t_R g224 ( 
.A(n_172),
.Y(n_224)
);

NAND2xp5_ASAP7_75t_SL g299 ( 
.A(n_224),
.B(n_229),
.Y(n_299)
);

OAI22xp33_ASAP7_75t_SL g225 ( 
.A1(n_171),
.A2(n_148),
.B1(n_212),
.B2(n_191),
.Y(n_225)
);

AOI22xp5_ASAP7_75t_SL g306 ( 
.A1(n_225),
.A2(n_246),
.B1(n_285),
.B2(n_219),
.Y(n_306)
);

NAND2xp5_ASAP7_75t_L g226 ( 
.A(n_200),
.B(n_151),
.Y(n_226)
);

AOI22xp33_ASAP7_75t_L g227 ( 
.A1(n_199),
.A2(n_204),
.B1(n_197),
.B2(n_196),
.Y(n_227)
);

OAI22xp5_ASAP7_75t_L g307 ( 
.A1(n_227),
.A2(n_231),
.B1(n_265),
.B2(n_284),
.Y(n_307)
);

AOI22xp33_ASAP7_75t_SL g228 ( 
.A1(n_157),
.A2(n_155),
.B1(n_137),
.B2(n_145),
.Y(n_228)
);

INVxp67_ASAP7_75t_L g315 ( 
.A(n_228),
.Y(n_315)
);

CKINVDCx20_ASAP7_75t_R g229 ( 
.A(n_178),
.Y(n_229)
);

NAND3xp33_ASAP7_75t_L g328 ( 
.A(n_230),
.B(n_252),
.C(n_258),
.Y(n_328)
);

AOI22xp5_ASAP7_75t_L g231 ( 
.A1(n_128),
.A2(n_133),
.B1(n_168),
.B2(n_173),
.Y(n_231)
);

CKINVDCx16_ASAP7_75t_R g232 ( 
.A(n_178),
.Y(n_232)
);

NAND2xp5_ASAP7_75t_SL g310 ( 
.A(n_232),
.B(n_243),
.Y(n_310)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_195),
.Y(n_233)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_233),
.Y(n_295)
);

NAND2xp5_ASAP7_75t_L g234 ( 
.A(n_130),
.B(n_138),
.Y(n_234)
);

NAND2xp5_ASAP7_75t_L g293 ( 
.A(n_234),
.B(n_236),
.Y(n_293)
);

NAND2xp5_ASAP7_75t_L g236 ( 
.A(n_143),
.B(n_147),
.Y(n_236)
);

OAI22xp5_ASAP7_75t_SL g237 ( 
.A1(n_193),
.A2(n_153),
.B1(n_139),
.B2(n_162),
.Y(n_237)
);

AOI22xp5_ASAP7_75t_L g291 ( 
.A1(n_237),
.A2(n_273),
.B1(n_238),
.B2(n_258),
.Y(n_291)
);

INVxp67_ASAP7_75t_L g238 ( 
.A(n_131),
.Y(n_238)
);

INVxp67_ASAP7_75t_L g321 ( 
.A(n_238),
.Y(n_321)
);

AOI22xp33_ASAP7_75t_SL g240 ( 
.A1(n_155),
.A2(n_163),
.B1(n_158),
.B2(n_135),
.Y(n_240)
);

INVxp67_ASAP7_75t_L g322 ( 
.A(n_240),
.Y(n_322)
);

INVxp67_ASAP7_75t_L g241 ( 
.A(n_198),
.Y(n_241)
);

INVxp67_ASAP7_75t_L g324 ( 
.A(n_241),
.Y(n_324)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_208),
.Y(n_242)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_242),
.Y(n_303)
);

NAND2xp5_ASAP7_75t_L g243 ( 
.A(n_160),
.B(n_190),
.Y(n_243)
);

INVx2_ASAP7_75t_L g244 ( 
.A(n_207),
.Y(n_244)
);

INVx2_ASAP7_75t_L g245 ( 
.A(n_135),
.Y(n_245)
);

OAI22xp33_ASAP7_75t_SL g246 ( 
.A1(n_158),
.A2(n_162),
.B1(n_163),
.B2(n_203),
.Y(n_246)
);

AOI22xp33_ASAP7_75t_SL g247 ( 
.A1(n_198),
.A2(n_202),
.B1(n_187),
.B2(n_152),
.Y(n_247)
);

AOI22xp33_ASAP7_75t_SL g334 ( 
.A1(n_247),
.A2(n_269),
.B1(n_277),
.B2(n_281),
.Y(n_334)
);

INVx8_ASAP7_75t_L g248 ( 
.A(n_181),
.Y(n_248)
);

HB1xp67_ASAP7_75t_L g249 ( 
.A(n_206),
.Y(n_249)
);

BUFx2_ASAP7_75t_L g330 ( 
.A(n_249),
.Y(n_330)
);

CKINVDCx20_ASAP7_75t_R g252 ( 
.A(n_194),
.Y(n_252)
);

NAND2xp5_ASAP7_75t_L g253 ( 
.A(n_165),
.B(n_170),
.Y(n_253)
);

OAI32xp33_ASAP7_75t_L g316 ( 
.A1(n_253),
.A2(n_268),
.A3(n_278),
.B1(n_254),
.B2(n_220),
.Y(n_316)
);

INVx2_ASAP7_75t_L g254 ( 
.A(n_165),
.Y(n_254)
);

BUFx4f_ASAP7_75t_L g256 ( 
.A(n_136),
.Y(n_256)
);

INVx2_ASAP7_75t_SL g305 ( 
.A(n_256),
.Y(n_305)
);

A2O1A1Ixp33_ASAP7_75t_L g258 ( 
.A1(n_146),
.A2(n_176),
.B(n_201),
.C(n_136),
.Y(n_258)
);

INVx3_ASAP7_75t_L g259 ( 
.A(n_194),
.Y(n_259)
);

INVx3_ASAP7_75t_L g300 ( 
.A(n_259),
.Y(n_300)
);

AND2x2_ASAP7_75t_SL g260 ( 
.A(n_129),
.B(n_167),
.Y(n_260)
);

CKINVDCx16_ASAP7_75t_R g323 ( 
.A(n_260),
.Y(n_323)
);

NAND2xp5_ASAP7_75t_SL g261 ( 
.A(n_144),
.B(n_132),
.Y(n_261)
);

NOR2xp33_ASAP7_75t_L g287 ( 
.A(n_261),
.B(n_262),
.Y(n_287)
);

INVxp67_ASAP7_75t_L g262 ( 
.A(n_176),
.Y(n_262)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_164),
.Y(n_264)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_264),
.Y(n_304)
);

AOI22xp33_ASAP7_75t_L g265 ( 
.A1(n_164),
.A2(n_170),
.B1(n_132),
.B2(n_134),
.Y(n_265)
);

CKINVDCx20_ASAP7_75t_R g266 ( 
.A(n_134),
.Y(n_266)
);

NOR2xp33_ASAP7_75t_L g308 ( 
.A(n_266),
.B(n_275),
.Y(n_308)
);

INVx5_ASAP7_75t_L g267 ( 
.A(n_181),
.Y(n_267)
);

NAND2xp5_ASAP7_75t_L g268 ( 
.A(n_166),
.B(n_174),
.Y(n_268)
);

AOI22xp33_ASAP7_75t_SL g269 ( 
.A1(n_129),
.A2(n_181),
.B1(n_141),
.B2(n_161),
.Y(n_269)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_150),
.Y(n_270)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_270),
.Y(n_319)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_150),
.Y(n_271)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_271),
.Y(n_329)
);

CKINVDCx16_ASAP7_75t_R g274 ( 
.A(n_176),
.Y(n_274)
);

INVx11_ASAP7_75t_L g302 ( 
.A(n_274),
.Y(n_302)
);

INVxp67_ASAP7_75t_L g275 ( 
.A(n_141),
.Y(n_275)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_126),
.Y(n_276)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_276),
.Y(n_286)
);

INVx1_ASAP7_75t_SL g277 ( 
.A(n_126),
.Y(n_277)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_188),
.Y(n_278)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_278),
.Y(n_296)
);

INVx2_ASAP7_75t_L g279 ( 
.A(n_167),
.Y(n_279)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_279),
.Y(n_298)
);

INVxp67_ASAP7_75t_L g280 ( 
.A(n_161),
.Y(n_280)
);

NOR2xp33_ASAP7_75t_L g309 ( 
.A(n_280),
.B(n_282),
.Y(n_309)
);

AOI22xp33_ASAP7_75t_SL g281 ( 
.A1(n_167),
.A2(n_96),
.B1(n_23),
.B2(n_39),
.Y(n_281)
);

OR2x2_ASAP7_75t_L g282 ( 
.A(n_142),
.B(n_169),
.Y(n_282)
);

NOR2xp33_ASAP7_75t_L g283 ( 
.A(n_142),
.B(n_160),
.Y(n_283)
);

NOR2xp33_ASAP7_75t_L g326 ( 
.A(n_283),
.B(n_250),
.Y(n_326)
);

AOI22xp5_ASAP7_75t_L g284 ( 
.A1(n_204),
.A2(n_199),
.B1(n_185),
.B2(n_200),
.Y(n_284)
);

AOI22xp33_ASAP7_75t_SL g285 ( 
.A1(n_148),
.A2(n_96),
.B1(n_23),
.B2(n_39),
.Y(n_285)
);

CKINVDCx20_ASAP7_75t_R g290 ( 
.A(n_217),
.Y(n_290)
);

NAND2xp5_ASAP7_75t_SL g335 ( 
.A(n_290),
.B(n_294),
.Y(n_335)
);

AOI22xp5_ASAP7_75t_L g350 ( 
.A1(n_291),
.A2(n_323),
.B1(n_321),
.B2(n_315),
.Y(n_350)
);

CKINVDCx20_ASAP7_75t_R g294 ( 
.A(n_234),
.Y(n_294)
);

INVx8_ASAP7_75t_L g301 ( 
.A(n_224),
.Y(n_301)
);

INVx2_ASAP7_75t_L g351 ( 
.A(n_301),
.Y(n_351)
);

AND2x2_ASAP7_75t_L g371 ( 
.A(n_306),
.B(n_316),
.Y(n_371)
);

MAJx2_ASAP7_75t_L g312 ( 
.A(n_236),
.B(n_243),
.C(n_257),
.Y(n_312)
);

MAJIxp5_ASAP7_75t_L g358 ( 
.A(n_312),
.B(n_320),
.C(n_260),
.Y(n_358)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_214),
.Y(n_313)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_313),
.Y(n_340)
);

CKINVDCx20_ASAP7_75t_R g314 ( 
.A(n_263),
.Y(n_314)
);

NAND2xp5_ASAP7_75t_SL g337 ( 
.A(n_314),
.B(n_250),
.Y(n_337)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_244),
.Y(n_318)
);

INVx1_ASAP7_75t_L g348 ( 
.A(n_318),
.Y(n_348)
);

MAJIxp5_ASAP7_75t_L g320 ( 
.A(n_257),
.B(n_239),
.C(n_229),
.Y(n_320)
);

BUFx6f_ASAP7_75t_L g325 ( 
.A(n_213),
.Y(n_325)
);

BUFx6f_ASAP7_75t_L g336 ( 
.A(n_325),
.Y(n_336)
);

NOR2xp33_ASAP7_75t_L g360 ( 
.A(n_326),
.B(n_233),
.Y(n_360)
);

AOI22xp33_ASAP7_75t_L g327 ( 
.A1(n_273),
.A2(n_251),
.B1(n_216),
.B2(n_284),
.Y(n_327)
);

AOI22xp33_ASAP7_75t_SL g355 ( 
.A1(n_327),
.A2(n_253),
.B1(n_268),
.B2(n_252),
.Y(n_355)
);

AOI22xp5_ASAP7_75t_L g331 ( 
.A1(n_251),
.A2(n_216),
.B1(n_237),
.B2(n_226),
.Y(n_331)
);

OAI22xp5_ASAP7_75t_SL g369 ( 
.A1(n_331),
.A2(n_276),
.B1(n_256),
.B2(n_279),
.Y(n_369)
);

INVx5_ASAP7_75t_L g332 ( 
.A(n_218),
.Y(n_332)
);

BUFx6f_ASAP7_75t_L g338 ( 
.A(n_332),
.Y(n_338)
);

INVx6_ASAP7_75t_L g333 ( 
.A(n_248),
.Y(n_333)
);

INVx1_ASAP7_75t_L g352 ( 
.A(n_333),
.Y(n_352)
);

NOR2xp33_ASAP7_75t_SL g376 ( 
.A(n_337),
.B(n_360),
.Y(n_376)
);

AOI21xp5_ASAP7_75t_SL g339 ( 
.A1(n_309),
.A2(n_257),
.B(n_223),
.Y(n_339)
);

NOR2xp67_ASAP7_75t_SL g386 ( 
.A(n_339),
.B(n_368),
.Y(n_386)
);

MAJx2_ASAP7_75t_L g341 ( 
.A(n_312),
.B(n_231),
.C(n_239),
.Y(n_341)
);

MAJIxp5_ASAP7_75t_L g391 ( 
.A(n_341),
.B(n_353),
.C(n_358),
.Y(n_391)
);

NAND2xp5_ASAP7_75t_L g342 ( 
.A(n_293),
.B(n_235),
.Y(n_342)
);

NAND2xp5_ASAP7_75t_L g397 ( 
.A(n_342),
.B(n_359),
.Y(n_397)
);

CKINVDCx16_ASAP7_75t_R g343 ( 
.A(n_330),
.Y(n_343)
);

NOR2xp33_ASAP7_75t_L g384 ( 
.A(n_343),
.B(n_345),
.Y(n_384)
);

OAI21xp5_ASAP7_75t_SL g344 ( 
.A1(n_315),
.A2(n_282),
.B(n_221),
.Y(n_344)
);

INVxp67_ASAP7_75t_L g377 ( 
.A(n_344),
.Y(n_377)
);

INVxp67_ASAP7_75t_L g345 ( 
.A(n_311),
.Y(n_345)
);

CKINVDCx20_ASAP7_75t_R g346 ( 
.A(n_330),
.Y(n_346)
);

NOR2xp33_ASAP7_75t_L g388 ( 
.A(n_346),
.B(n_373),
.Y(n_388)
);

FAx1_ASAP7_75t_SL g347 ( 
.A(n_320),
.B(n_282),
.CI(n_272),
.CON(n_347),
.SN(n_347)
);

NOR2xp33_ASAP7_75t_SL g383 ( 
.A(n_347),
.B(n_349),
.Y(n_383)
);

NAND2xp5_ASAP7_75t_SL g349 ( 
.A(n_293),
.B(n_255),
.Y(n_349)
);

AOI22xp5_ASAP7_75t_L g404 ( 
.A1(n_350),
.A2(n_369),
.B1(n_305),
.B2(n_304),
.Y(n_404)
);

XOR2xp5_ASAP7_75t_L g353 ( 
.A(n_310),
.B(n_222),
.Y(n_353)
);

AOI21xp5_ASAP7_75t_L g354 ( 
.A1(n_321),
.A2(n_222),
.B(n_241),
.Y(n_354)
);

AND2x2_ASAP7_75t_L g385 ( 
.A(n_354),
.B(n_366),
.Y(n_385)
);

OAI22xp5_ASAP7_75t_SL g380 ( 
.A1(n_355),
.A2(n_292),
.B1(n_334),
.B2(n_322),
.Y(n_380)
);

CKINVDCx20_ASAP7_75t_R g356 ( 
.A(n_325),
.Y(n_356)
);

INVx13_ASAP7_75t_L g405 ( 
.A(n_356),
.Y(n_405)
);

AOI22xp33_ASAP7_75t_SL g357 ( 
.A1(n_322),
.A2(n_222),
.B1(n_266),
.B2(n_256),
.Y(n_357)
);

BUFx12_ASAP7_75t_L g407 ( 
.A(n_357),
.Y(n_407)
);

A2O1A1Ixp33_ASAP7_75t_L g359 ( 
.A1(n_289),
.A2(n_222),
.B(n_242),
.C(n_260),
.Y(n_359)
);

BUFx24_ASAP7_75t_L g361 ( 
.A(n_302),
.Y(n_361)
);

INVx1_ASAP7_75t_L g362 ( 
.A(n_288),
.Y(n_362)
);

INVx1_ASAP7_75t_L g389 ( 
.A(n_362),
.Y(n_389)
);

NAND2xp5_ASAP7_75t_SL g363 ( 
.A(n_289),
.B(n_245),
.Y(n_363)
);

NOR2xp33_ASAP7_75t_SL g400 ( 
.A(n_363),
.B(n_372),
.Y(n_400)
);

INVx1_ASAP7_75t_L g364 ( 
.A(n_288),
.Y(n_364)
);

INVx1_ASAP7_75t_L g390 ( 
.A(n_364),
.Y(n_390)
);

NAND2xp5_ASAP7_75t_L g365 ( 
.A(n_331),
.B(n_271),
.Y(n_365)
);

NOR2x1_ASAP7_75t_L g382 ( 
.A(n_365),
.B(n_370),
.Y(n_382)
);

AOI22xp5_ASAP7_75t_SL g366 ( 
.A1(n_292),
.A2(n_274),
.B1(n_259),
.B2(n_270),
.Y(n_366)
);

MAJIxp5_ASAP7_75t_L g367 ( 
.A(n_297),
.B(n_262),
.C(n_264),
.Y(n_367)
);

MAJIxp5_ASAP7_75t_L g406 ( 
.A(n_367),
.B(n_324),
.C(n_286),
.Y(n_406)
);

AOI21xp5_ASAP7_75t_L g368 ( 
.A1(n_291),
.A2(n_280),
.B(n_275),
.Y(n_368)
);

NAND2xp5_ASAP7_75t_L g370 ( 
.A(n_316),
.B(n_267),
.Y(n_370)
);

NOR2xp33_ASAP7_75t_L g372 ( 
.A(n_287),
.B(n_277),
.Y(n_372)
);

INVxp67_ASAP7_75t_L g373 ( 
.A(n_308),
.Y(n_373)
);

INVx1_ASAP7_75t_L g374 ( 
.A(n_296),
.Y(n_374)
);

INVx1_ASAP7_75t_L g392 ( 
.A(n_374),
.Y(n_392)
);

NOR2xp33_ASAP7_75t_L g375 ( 
.A(n_297),
.B(n_213),
.Y(n_375)
);

NOR2xp33_ASAP7_75t_L g396 ( 
.A(n_375),
.B(n_324),
.Y(n_396)
);

XOR2xp5_ASAP7_75t_L g378 ( 
.A(n_358),
.B(n_299),
.Y(n_378)
);

MAJIxp5_ASAP7_75t_L g411 ( 
.A(n_378),
.B(n_406),
.C(n_373),
.Y(n_411)
);

OAI22x1_ASAP7_75t_SL g379 ( 
.A1(n_350),
.A2(n_306),
.B1(n_328),
.B2(n_307),
.Y(n_379)
);

OA21x2_ASAP7_75t_L g423 ( 
.A1(n_379),
.A2(n_351),
.B(n_352),
.Y(n_423)
);

AOI22xp5_ASAP7_75t_SL g412 ( 
.A1(n_380),
.A2(n_371),
.B1(n_370),
.B2(n_369),
.Y(n_412)
);

AND2x6_ASAP7_75t_L g381 ( 
.A(n_347),
.B(n_302),
.Y(n_381)
);

NAND2xp5_ASAP7_75t_SL g408 ( 
.A(n_381),
.B(n_387),
.Y(n_408)
);

AND2x6_ASAP7_75t_L g387 ( 
.A(n_347),
.B(n_301),
.Y(n_387)
);

CKINVDCx20_ASAP7_75t_R g393 ( 
.A(n_335),
.Y(n_393)
);

NAND2xp5_ASAP7_75t_SL g414 ( 
.A(n_393),
.B(n_394),
.Y(n_414)
);

CKINVDCx20_ASAP7_75t_R g394 ( 
.A(n_345),
.Y(n_394)
);

INVx1_ASAP7_75t_L g395 ( 
.A(n_362),
.Y(n_395)
);

INVx1_ASAP7_75t_L g409 ( 
.A(n_395),
.Y(n_409)
);

NAND2xp5_ASAP7_75t_SL g434 ( 
.A(n_396),
.B(n_402),
.Y(n_434)
);

OAI22xp5_ASAP7_75t_SL g398 ( 
.A1(n_371),
.A2(n_303),
.B1(n_329),
.B2(n_319),
.Y(n_398)
);

AOI22xp5_ASAP7_75t_L g425 ( 
.A1(n_398),
.A2(n_401),
.B1(n_404),
.B2(n_374),
.Y(n_425)
);

INVx1_ASAP7_75t_L g399 ( 
.A(n_364),
.Y(n_399)
);

INVx1_ASAP7_75t_L g424 ( 
.A(n_399),
.Y(n_424)
);

OAI22xp5_ASAP7_75t_SL g401 ( 
.A1(n_371),
.A2(n_303),
.B1(n_329),
.B2(n_319),
.Y(n_401)
);

INVx1_ASAP7_75t_L g402 ( 
.A(n_340),
.Y(n_402)
);

CKINVDCx20_ASAP7_75t_R g403 ( 
.A(n_338),
.Y(n_403)
);

CKINVDCx20_ASAP7_75t_R g410 ( 
.A(n_403),
.Y(n_410)
);

MAJIxp5_ASAP7_75t_L g438 ( 
.A(n_411),
.B(n_418),
.C(n_420),
.Y(n_438)
);

OAI22xp5_ASAP7_75t_L g447 ( 
.A1(n_412),
.A2(n_417),
.B1(n_423),
.B2(n_425),
.Y(n_447)
);

CKINVDCx20_ASAP7_75t_R g413 ( 
.A(n_388),
.Y(n_413)
);

NAND2xp5_ASAP7_75t_L g448 ( 
.A(n_413),
.B(n_415),
.Y(n_448)
);

CKINVDCx16_ASAP7_75t_R g415 ( 
.A(n_384),
.Y(n_415)
);

OAI21xp5_ASAP7_75t_SL g416 ( 
.A1(n_377),
.A2(n_354),
.B(n_368),
.Y(n_416)
);

INVxp67_ASAP7_75t_L g459 ( 
.A(n_416),
.Y(n_459)
);

OAI22xp5_ASAP7_75t_L g417 ( 
.A1(n_397),
.A2(n_353),
.B1(n_365),
.B2(n_342),
.Y(n_417)
);

MAJIxp5_ASAP7_75t_L g418 ( 
.A(n_391),
.B(n_378),
.C(n_341),
.Y(n_418)
);

OAI21xp5_ASAP7_75t_L g419 ( 
.A1(n_377),
.A2(n_359),
.B(n_344),
.Y(n_419)
);

HB1xp67_ASAP7_75t_L g458 ( 
.A(n_419),
.Y(n_458)
);

MAJIxp5_ASAP7_75t_L g420 ( 
.A(n_391),
.B(n_339),
.C(n_367),
.Y(n_420)
);

XNOR2xp5_ASAP7_75t_L g421 ( 
.A(n_397),
.B(n_340),
.Y(n_421)
);

XOR2xp5_ASAP7_75t_L g450 ( 
.A(n_421),
.B(n_401),
.Y(n_450)
);

AOI21xp5_ASAP7_75t_L g422 ( 
.A1(n_385),
.A2(n_351),
.B(n_366),
.Y(n_422)
);

BUFx12f_ASAP7_75t_L g442 ( 
.A(n_422),
.Y(n_442)
);

FAx1_ASAP7_75t_SL g426 ( 
.A(n_383),
.B(n_361),
.CI(n_348),
.CON(n_426),
.SN(n_426)
);

NOR2xp33_ASAP7_75t_L g440 ( 
.A(n_426),
.B(n_428),
.Y(n_440)
);

MAJIxp5_ASAP7_75t_L g427 ( 
.A(n_406),
.B(n_295),
.C(n_298),
.Y(n_427)
);

MAJIxp5_ASAP7_75t_L g443 ( 
.A(n_427),
.B(n_386),
.C(n_402),
.Y(n_443)
);

AOI21xp5_ASAP7_75t_L g428 ( 
.A1(n_385),
.A2(n_356),
.B(n_361),
.Y(n_428)
);

NAND3xp33_ASAP7_75t_L g429 ( 
.A(n_393),
.B(n_348),
.C(n_295),
.Y(n_429)
);

NOR2xp33_ASAP7_75t_L g441 ( 
.A(n_429),
.B(n_431),
.Y(n_441)
);

OA21x2_ASAP7_75t_L g430 ( 
.A1(n_385),
.A2(n_352),
.B(n_361),
.Y(n_430)
);

AOI22xp5_ASAP7_75t_L g455 ( 
.A1(n_430),
.A2(n_432),
.B1(n_433),
.B2(n_395),
.Y(n_455)
);

CKINVDCx20_ASAP7_75t_R g431 ( 
.A(n_376),
.Y(n_431)
);

OAI22xp5_ASAP7_75t_SL g432 ( 
.A1(n_404),
.A2(n_338),
.B1(n_336),
.B2(n_300),
.Y(n_432)
);

OAI22xp5_ASAP7_75t_SL g433 ( 
.A1(n_382),
.A2(n_336),
.B1(n_300),
.B2(n_304),
.Y(n_433)
);

OAI22xp5_ASAP7_75t_L g435 ( 
.A1(n_382),
.A2(n_332),
.B1(n_333),
.B2(n_317),
.Y(n_435)
);

OAI22xp5_ASAP7_75t_L g452 ( 
.A1(n_435),
.A2(n_423),
.B1(n_422),
.B2(n_425),
.Y(n_452)
);

CKINVDCx20_ASAP7_75t_R g436 ( 
.A(n_400),
.Y(n_436)
);

NOR2xp33_ASAP7_75t_L g461 ( 
.A(n_436),
.B(n_392),
.Y(n_461)
);

NAND2xp5_ASAP7_75t_SL g437 ( 
.A(n_415),
.B(n_383),
.Y(n_437)
);

NOR2xp33_ASAP7_75t_SL g465 ( 
.A(n_437),
.B(n_461),
.Y(n_465)
);

CKINVDCx20_ASAP7_75t_R g439 ( 
.A(n_414),
.Y(n_439)
);

NOR2xp33_ASAP7_75t_L g469 ( 
.A(n_439),
.B(n_444),
.Y(n_469)
);

MAJIxp5_ASAP7_75t_L g474 ( 
.A(n_443),
.B(n_446),
.C(n_453),
.Y(n_474)
);

CKINVDCx20_ASAP7_75t_R g444 ( 
.A(n_434),
.Y(n_444)
);

XNOR2xp5_ASAP7_75t_L g445 ( 
.A(n_418),
.B(n_411),
.Y(n_445)
);

XOR2xp5_ASAP7_75t_L g466 ( 
.A(n_445),
.B(n_450),
.Y(n_466)
);

MAJIxp5_ASAP7_75t_L g446 ( 
.A(n_420),
.B(n_386),
.C(n_398),
.Y(n_446)
);

INVx1_ASAP7_75t_L g449 ( 
.A(n_409),
.Y(n_449)
);

INVx1_ASAP7_75t_L g464 ( 
.A(n_449),
.Y(n_464)
);

OAI22xp5_ASAP7_75t_SL g451 ( 
.A1(n_412),
.A2(n_387),
.B1(n_381),
.B2(n_379),
.Y(n_451)
);

AOI22xp5_ASAP7_75t_L g477 ( 
.A1(n_451),
.A2(n_452),
.B1(n_457),
.B2(n_430),
.Y(n_477)
);

MAJIxp5_ASAP7_75t_L g453 ( 
.A(n_427),
.B(n_394),
.C(n_399),
.Y(n_453)
);

XNOR2xp5_ASAP7_75t_L g454 ( 
.A(n_417),
.B(n_389),
.Y(n_454)
);

XOR2xp5_ASAP7_75t_L g482 ( 
.A(n_454),
.B(n_460),
.Y(n_482)
);

OAI22xp5_ASAP7_75t_L g476 ( 
.A1(n_455),
.A2(n_435),
.B1(n_430),
.B2(n_428),
.Y(n_476)
);

OAI22xp5_ASAP7_75t_L g456 ( 
.A1(n_436),
.A2(n_390),
.B1(n_389),
.B2(n_403),
.Y(n_456)
);

INVx1_ASAP7_75t_L g467 ( 
.A(n_456),
.Y(n_467)
);

OAI22xp5_ASAP7_75t_SL g457 ( 
.A1(n_408),
.A2(n_407),
.B1(n_390),
.B2(n_380),
.Y(n_457)
);

XNOR2xp5_ASAP7_75t_L g460 ( 
.A(n_421),
.B(n_419),
.Y(n_460)
);

XNOR2xp5_ASAP7_75t_SL g462 ( 
.A(n_416),
.B(n_392),
.Y(n_462)
);

NAND2xp5_ASAP7_75t_SL g463 ( 
.A(n_462),
.B(n_423),
.Y(n_463)
);

XNOR2xp5_ASAP7_75t_L g492 ( 
.A(n_463),
.B(n_478),
.Y(n_492)
);

NAND2xp5_ASAP7_75t_L g468 ( 
.A(n_448),
.B(n_413),
.Y(n_468)
);

INVx1_ASAP7_75t_L g485 ( 
.A(n_468),
.Y(n_485)
);

NAND2xp5_ASAP7_75t_L g470 ( 
.A(n_441),
.B(n_433),
.Y(n_470)
);

INVx1_ASAP7_75t_L g488 ( 
.A(n_470),
.Y(n_488)
);

INVx1_ASAP7_75t_L g471 ( 
.A(n_455),
.Y(n_471)
);

INVx1_ASAP7_75t_L g490 ( 
.A(n_471),
.Y(n_490)
);

NOR2xp33_ASAP7_75t_L g472 ( 
.A(n_453),
.B(n_431),
.Y(n_472)
);

INVx1_ASAP7_75t_L g493 ( 
.A(n_472),
.Y(n_493)
);

NOR2xp33_ASAP7_75t_SL g473 ( 
.A(n_460),
.B(n_410),
.Y(n_473)
);

OAI22xp5_ASAP7_75t_L g489 ( 
.A1(n_473),
.A2(n_476),
.B1(n_477),
.B2(n_479),
.Y(n_489)
);

INVx1_ASAP7_75t_L g475 ( 
.A(n_447),
.Y(n_475)
);

INVx1_ASAP7_75t_L g497 ( 
.A(n_475),
.Y(n_497)
);

NAND2xp5_ASAP7_75t_L g478 ( 
.A(n_454),
.B(n_410),
.Y(n_478)
);

AOI22xp5_ASAP7_75t_L g479 ( 
.A1(n_457),
.A2(n_432),
.B1(n_426),
.B2(n_407),
.Y(n_479)
);

NOR2xp33_ASAP7_75t_SL g480 ( 
.A(n_443),
.B(n_409),
.Y(n_480)
);

NOR2xp33_ASAP7_75t_L g486 ( 
.A(n_480),
.B(n_481),
.Y(n_486)
);

CKINVDCx20_ASAP7_75t_R g481 ( 
.A(n_440),
.Y(n_481)
);

OAI21xp5_ASAP7_75t_L g483 ( 
.A1(n_458),
.A2(n_426),
.B(n_424),
.Y(n_483)
);

O2A1O1Ixp33_ASAP7_75t_L g491 ( 
.A1(n_483),
.A2(n_459),
.B(n_462),
.C(n_450),
.Y(n_491)
);

MAJIxp5_ASAP7_75t_L g484 ( 
.A(n_474),
.B(n_445),
.C(n_438),
.Y(n_484)
);

MAJIxp5_ASAP7_75t_L g509 ( 
.A(n_484),
.B(n_467),
.C(n_475),
.Y(n_509)
);

XOR2xp5_ASAP7_75t_L g487 ( 
.A(n_466),
.B(n_446),
.Y(n_487)
);

MAJx2_ASAP7_75t_L g512 ( 
.A(n_487),
.B(n_494),
.C(n_495),
.Y(n_512)
);

OAI21xp5_ASAP7_75t_L g500 ( 
.A1(n_491),
.A2(n_463),
.B(n_483),
.Y(n_500)
);

XOR2xp5_ASAP7_75t_SL g494 ( 
.A(n_482),
.B(n_451),
.Y(n_494)
);

XOR2xp5_ASAP7_75t_L g495 ( 
.A(n_466),
.B(n_438),
.Y(n_495)
);

XOR2xp5_ASAP7_75t_L g496 ( 
.A(n_474),
.B(n_459),
.Y(n_496)
);

XOR2xp5_ASAP7_75t_L g501 ( 
.A(n_496),
.B(n_478),
.Y(n_501)
);

XNOR2xp5_ASAP7_75t_L g498 ( 
.A(n_482),
.B(n_424),
.Y(n_498)
);

NOR2xp33_ASAP7_75t_L g507 ( 
.A(n_498),
.B(n_499),
.Y(n_507)
);

XNOR2xp5_ASAP7_75t_L g499 ( 
.A(n_480),
.B(n_442),
.Y(n_499)
);

OR2x2_ASAP7_75t_L g513 ( 
.A(n_500),
.B(n_505),
.Y(n_513)
);

XNOR2xp5_ASAP7_75t_L g521 ( 
.A(n_501),
.B(n_498),
.Y(n_521)
);

INVx1_ASAP7_75t_L g502 ( 
.A(n_485),
.Y(n_502)
);

INVx1_ASAP7_75t_L g517 ( 
.A(n_502),
.Y(n_517)
);

NOR2xp67_ASAP7_75t_L g503 ( 
.A(n_493),
.B(n_465),
.Y(n_503)
);

NAND2xp5_ASAP7_75t_L g519 ( 
.A(n_503),
.B(n_504),
.Y(n_519)
);

INVx1_ASAP7_75t_L g504 ( 
.A(n_488),
.Y(n_504)
);

OAI21xp5_ASAP7_75t_L g505 ( 
.A1(n_491),
.A2(n_481),
.B(n_471),
.Y(n_505)
);

INVx1_ASAP7_75t_L g506 ( 
.A(n_486),
.Y(n_506)
);

NAND2xp5_ASAP7_75t_L g522 ( 
.A(n_506),
.B(n_509),
.Y(n_522)
);

OAI21xp5_ASAP7_75t_SL g508 ( 
.A1(n_489),
.A2(n_468),
.B(n_470),
.Y(n_508)
);

OAI21xp5_ASAP7_75t_L g514 ( 
.A1(n_508),
.A2(n_473),
.B(n_479),
.Y(n_514)
);

AOI22xp33_ASAP7_75t_SL g510 ( 
.A1(n_497),
.A2(n_476),
.B1(n_467),
.B2(n_442),
.Y(n_510)
);

INVxp67_ASAP7_75t_L g516 ( 
.A(n_510),
.Y(n_516)
);

INVx1_ASAP7_75t_L g511 ( 
.A(n_490),
.Y(n_511)
);

NOR2xp33_ASAP7_75t_L g520 ( 
.A(n_511),
.B(n_465),
.Y(n_520)
);

NAND2xp5_ASAP7_75t_L g529 ( 
.A(n_514),
.B(n_515),
.Y(n_529)
);

MAJIxp5_ASAP7_75t_L g515 ( 
.A(n_509),
.B(n_484),
.C(n_495),
.Y(n_515)
);

MAJIxp5_ASAP7_75t_L g518 ( 
.A(n_501),
.B(n_496),
.C(n_487),
.Y(n_518)
);

INVxp67_ASAP7_75t_SL g525 ( 
.A(n_518),
.Y(n_525)
);

NOR2xp33_ASAP7_75t_L g528 ( 
.A(n_520),
.B(n_523),
.Y(n_528)
);

XOR2xp5_ASAP7_75t_L g524 ( 
.A(n_521),
.B(n_500),
.Y(n_524)
);

NOR2xp33_ASAP7_75t_SL g523 ( 
.A(n_507),
.B(n_469),
.Y(n_523)
);

NOR2xp33_ASAP7_75t_L g533 ( 
.A(n_524),
.B(n_527),
.Y(n_533)
);

OAI21x1_ASAP7_75t_L g526 ( 
.A1(n_522),
.A2(n_505),
.B(n_477),
.Y(n_526)
);

NOR2xp67_ASAP7_75t_L g535 ( 
.A(n_526),
.B(n_513),
.Y(n_535)
);

MAJIxp5_ASAP7_75t_L g527 ( 
.A(n_515),
.B(n_512),
.C(n_510),
.Y(n_527)
);

AOI322xp5_ASAP7_75t_L g530 ( 
.A1(n_519),
.A2(n_407),
.A3(n_442),
.B1(n_464),
.B2(n_494),
.C1(n_405),
.C2(n_499),
.Y(n_530)
);

NOR2xp33_ASAP7_75t_L g534 ( 
.A(n_530),
.B(n_516),
.Y(n_534)
);

INVxp67_ASAP7_75t_L g531 ( 
.A(n_513),
.Y(n_531)
);

INVx1_ASAP7_75t_L g532 ( 
.A(n_531),
.Y(n_532)
);

INVxp67_ASAP7_75t_L g539 ( 
.A(n_534),
.Y(n_539)
);

MAJx2_ASAP7_75t_L g541 ( 
.A(n_535),
.B(n_536),
.C(n_524),
.Y(n_541)
);

AOI21xp5_ASAP7_75t_L g536 ( 
.A1(n_531),
.A2(n_516),
.B(n_492),
.Y(n_536)
);

NOR2xp33_ASAP7_75t_L g537 ( 
.A(n_529),
.B(n_517),
.Y(n_537)
);

NOR2xp33_ASAP7_75t_L g540 ( 
.A(n_537),
.B(n_525),
.Y(n_540)
);

FAx1_ASAP7_75t_SL g538 ( 
.A(n_532),
.B(n_518),
.CI(n_512),
.CON(n_538),
.SN(n_538)
);

OAI21xp5_ASAP7_75t_L g543 ( 
.A1(n_538),
.A2(n_536),
.B(n_539),
.Y(n_543)
);

AOI21x1_ASAP7_75t_L g542 ( 
.A1(n_540),
.A2(n_541),
.B(n_533),
.Y(n_542)
);

OAI21xp5_ASAP7_75t_L g544 ( 
.A1(n_542),
.A2(n_543),
.B(n_528),
.Y(n_544)
);

OAI21xp5_ASAP7_75t_L g545 ( 
.A1(n_544),
.A2(n_492),
.B(n_464),
.Y(n_545)
);

XNOR2xp5_ASAP7_75t_L g546 ( 
.A(n_545),
.B(n_405),
.Y(n_546)
);


endmodule