module real_jpeg_1538_n_29 (n_17, n_8, n_0, n_21, n_168, n_2, n_10, n_9, n_12, n_24, n_165, n_166, n_6, n_159, n_28, n_161, n_162, n_167, n_23, n_11, n_14, n_160, n_25, n_163, n_7, n_22, n_18, n_3, n_5, n_4, n_1, n_26, n_27, n_20, n_19, n_164, n_158, n_16, n_15, n_13, n_29);

input n_17;
input n_8;
input n_0;
input n_21;
input n_168;
input n_2;
input n_10;
input n_9;
input n_12;
input n_24;
input n_165;
input n_166;
input n_6;
input n_159;
input n_28;
input n_161;
input n_162;
input n_167;
input n_23;
input n_11;
input n_14;
input n_160;
input n_25;
input n_163;
input n_7;
input n_22;
input n_18;
input n_3;
input n_5;
input n_4;
input n_1;
input n_26;
input n_27;
input n_20;
input n_19;
input n_164;
input n_158;
input n_16;
input n_15;
input n_13;

output n_29;

wire n_108;
wire n_54;
wire n_37;
wire n_73;
wire n_35;
wire n_38;
wire n_91;
wire n_49;
wire n_114;
wire n_68;
wire n_146;
wire n_78;
wire n_83;
wire n_104;
wire n_153;
wire n_64;
wire n_47;
wire n_131;
wire n_87;
wire n_40;
wire n_105;
wire n_115;
wire n_98;
wire n_56;
wire n_48;
wire n_140;
wire n_126;
wire n_113;
wire n_120;
wire n_155;
wire n_93;
wire n_141;
wire n_95;
wire n_139;
wire n_33;
wire n_65;
wire n_142;
wire n_76;
wire n_67;
wire n_79;
wire n_107;
wire n_156;
wire n_147;
wire n_66;
wire n_136;
wire n_44;
wire n_62;
wire n_121;
wire n_106;
wire n_45;
wire n_112;
wire n_42;
wire n_145;
wire n_77;
wire n_109;
wire n_39;
wire n_122;
wire n_94;
wire n_148;
wire n_118;
wire n_123;
wire n_116;
wire n_50;
wire n_143;
wire n_69;
wire n_31;
wire n_137;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_134;
wire n_72;
wire n_151;
wire n_100;
wire n_51;
wire n_71;
wire n_90;
wire n_110;
wire n_61;
wire n_117;
wire n_99;
wire n_86;
wire n_150;
wire n_41;
wire n_70;
wire n_80;
wire n_32;
wire n_74;
wire n_30;
wire n_149;
wire n_144;
wire n_130;
wire n_103;
wire n_57;
wire n_43;
wire n_84;
wire n_82;
wire n_111;
wire n_132;
wire n_125;
wire n_55;
wire n_58;
wire n_52;
wire n_63;
wire n_124;
wire n_92;
wire n_75;
wire n_97;
wire n_34;
wire n_60;
wire n_46;
wire n_88;
wire n_59;
wire n_128;
wire n_133;
wire n_138;
wire n_53;
wire n_127;
wire n_119;
wire n_36;
wire n_81;
wire n_102;
wire n_85;
wire n_101;
wire n_96;
wire n_89;

CKINVDCx20_ASAP7_75t_R g151 ( 
.A(n_0),
.Y(n_151)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_1),
.Y(n_123)
);

AO22x1_ASAP7_75t_L g79 ( 
.A1(n_2),
.A2(n_80),
.B1(n_82),
.B2(n_93),
.Y(n_79)
);

CKINVDCx20_ASAP7_75t_R g92 ( 
.A(n_2),
.Y(n_92)
);

AND2x2_ASAP7_75t_L g84 ( 
.A(n_3),
.B(n_85),
.Y(n_84)
);

CKINVDCx20_ASAP7_75t_R g146 ( 
.A(n_4),
.Y(n_146)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_5),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g72 ( 
.A(n_6),
.Y(n_72)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_7),
.Y(n_67)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_8),
.Y(n_103)
);

OAI21xp5_ASAP7_75t_SL g83 ( 
.A1(n_9),
.A2(n_84),
.B(n_88),
.Y(n_83)
);

INVx3_ASAP7_75t_L g38 ( 
.A(n_10),
.Y(n_38)
);

BUFx16f_ASAP7_75t_L g87 ( 
.A(n_10),
.Y(n_87)
);

BUFx4f_ASAP7_75t_SL g90 ( 
.A(n_10),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g118 ( 
.A(n_11),
.B(n_119),
.Y(n_118)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_11),
.Y(n_134)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_12),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_L g142 ( 
.A(n_12),
.B(n_57),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_L g115 ( 
.A(n_13),
.B(n_116),
.Y(n_115)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_13),
.Y(n_130)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_14),
.Y(n_96)
);

CKINVDCx20_ASAP7_75t_R g154 ( 
.A(n_15),
.Y(n_154)
);

CKINVDCx20_ASAP7_75t_R g141 ( 
.A(n_16),
.Y(n_141)
);

CKINVDCx20_ASAP7_75t_R g120 ( 
.A(n_17),
.Y(n_120)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_18),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g65 ( 
.A(n_19),
.Y(n_65)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_20),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g114 ( 
.A(n_20),
.B(n_70),
.Y(n_114)
);

CKINVDCx20_ASAP7_75t_R g58 ( 
.A(n_21),
.Y(n_58)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_22),
.Y(n_138)
);

MAJIxp5_ASAP7_75t_L g76 ( 
.A(n_23),
.B(n_77),
.C(n_101),
.Y(n_76)
);

AOI22xp5_ASAP7_75t_SL g74 ( 
.A1(n_24),
.A2(n_75),
.B1(n_107),
.B2(n_110),
.Y(n_74)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_24),
.Y(n_108)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_25),
.Y(n_53)
);

MAJIxp5_ASAP7_75t_L g78 ( 
.A(n_26),
.B(n_79),
.C(n_94),
.Y(n_78)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_27),
.Y(n_52)
);

AOI22xp5_ASAP7_75t_L g30 ( 
.A1(n_28),
.A2(n_31),
.B1(n_32),
.B2(n_39),
.Y(n_30)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_28),
.Y(n_39)
);

AOI22xp5_ASAP7_75t_SL g41 ( 
.A1(n_28),
.A2(n_42),
.B1(n_148),
.B2(n_150),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g43 ( 
.A(n_28),
.B(n_44),
.Y(n_43)
);

NAND2xp5_ASAP7_75t_L g147 ( 
.A(n_28),
.B(n_44),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_L g152 ( 
.A(n_28),
.B(n_153),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_L g156 ( 
.A(n_28),
.B(n_153),
.Y(n_156)
);

XOR2xp5_ASAP7_75t_L g29 ( 
.A(n_30),
.B(n_40),
.Y(n_29)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_32),
.Y(n_31)
);

NOR2xp33_ASAP7_75t_L g32 ( 
.A(n_33),
.B(n_34),
.Y(n_32)
);

NOR2xp33_ASAP7_75t_L g150 ( 
.A(n_34),
.B(n_151),
.Y(n_150)
);

BUFx2_ASAP7_75t_L g155 ( 
.A(n_34),
.Y(n_155)
);

BUFx4f_ASAP7_75t_SL g34 ( 
.A(n_35),
.Y(n_34)
);

BUFx3_ASAP7_75t_L g46 ( 
.A(n_35),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g51 ( 
.A(n_35),
.B(n_52),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g145 ( 
.A(n_35),
.B(n_146),
.Y(n_145)
);

INVx13_ASAP7_75t_L g35 ( 
.A(n_36),
.Y(n_35)
);

INVx3_ASAP7_75t_L g59 ( 
.A(n_36),
.Y(n_59)
);

CKINVDCx6p67_ASAP7_75t_R g36 ( 
.A(n_37),
.Y(n_36)
);

BUFx10_ASAP7_75t_L g66 ( 
.A(n_37),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_37),
.B(n_81),
.Y(n_80)
);

INVx5_ASAP7_75t_L g37 ( 
.A(n_38),
.Y(n_37)
);

INVx8_ASAP7_75t_L g71 ( 
.A(n_38),
.Y(n_71)
);

INVx6_ASAP7_75t_SL g100 ( 
.A(n_38),
.Y(n_100)
);

INVx4_ASAP7_75t_SL g121 ( 
.A(n_38),
.Y(n_121)
);

MAJx2_ASAP7_75t_L g47 ( 
.A(n_39),
.B(n_48),
.C(n_144),
.Y(n_47)
);

NAND2xp5_ASAP7_75t_L g148 ( 
.A(n_39),
.B(n_149),
.Y(n_148)
);

OAI21xp5_ASAP7_75t_L g40 ( 
.A1(n_41),
.A2(n_152),
.B(n_156),
.Y(n_40)
);

OAI21xp5_ASAP7_75t_L g42 ( 
.A1(n_43),
.A2(n_47),
.B(n_147),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g44 ( 
.A(n_45),
.B(n_46),
.Y(n_44)
);

AOI21xp5_ASAP7_75t_L g48 ( 
.A1(n_49),
.A2(n_54),
.B(n_143),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_SL g49 ( 
.A(n_50),
.B(n_53),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g143 ( 
.A(n_50),
.B(n_53),
.Y(n_143)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_51),
.Y(n_50)
);

A2O1A1Ixp33_ASAP7_75t_L g54 ( 
.A1(n_55),
.A2(n_56),
.B(n_60),
.C(n_142),
.Y(n_54)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_57),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g57 ( 
.A(n_58),
.B(n_59),
.Y(n_57)
);

MAJx2_ASAP7_75t_L g60 ( 
.A(n_61),
.B(n_138),
.C(n_139),
.Y(n_60)
);

AOI21xp5_ASAP7_75t_L g61 ( 
.A1(n_62),
.A2(n_68),
.B(n_137),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_SL g62 ( 
.A(n_63),
.B(n_67),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g137 ( 
.A(n_63),
.B(n_67),
.Y(n_137)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_64),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_65),
.B(n_66),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g125 ( 
.A(n_66),
.B(n_126),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_L g140 ( 
.A(n_66),
.B(n_141),
.Y(n_140)
);

OAI221xp5_ASAP7_75t_L g68 ( 
.A1(n_69),
.A2(n_73),
.B1(n_74),
.B2(n_112),
.C(n_127),
.Y(n_68)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_70),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_SL g70 ( 
.A(n_71),
.B(n_72),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_71),
.B(n_106),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_71),
.B(n_111),
.Y(n_110)
);

MAJIxp5_ASAP7_75t_L g75 ( 
.A(n_76),
.B(n_103),
.C(n_104),
.Y(n_75)
);

MAJIxp5_ASAP7_75t_L g77 ( 
.A(n_78),
.B(n_96),
.C(n_97),
.Y(n_77)
);

NAND3xp33_ASAP7_75t_L g82 ( 
.A(n_83),
.B(n_91),
.C(n_92),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_L g93 ( 
.A(n_83),
.B(n_91),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_L g91 ( 
.A(n_84),
.B(n_88),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_86),
.B(n_87),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_87),
.B(n_95),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_87),
.B(n_102),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_SL g116 ( 
.A(n_87),
.B(n_117),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_89),
.B(n_90),
.Y(n_88)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_98),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_99),
.B(n_100),
.Y(n_98)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_105),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_L g107 ( 
.A(n_108),
.B(n_109),
.Y(n_107)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_110),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_SL g112 ( 
.A(n_113),
.B(n_122),
.Y(n_112)
);

AOI322xp5_ASAP7_75t_L g127 ( 
.A1(n_113),
.A2(n_128),
.A3(n_129),
.B1(n_132),
.B2(n_133),
.C1(n_136),
.C2(n_168),
.Y(n_127)
);

NOR3xp33_ASAP7_75t_SL g113 ( 
.A(n_114),
.B(n_115),
.C(n_118),
.Y(n_113)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_114),
.Y(n_132)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_116),
.Y(n_131)
);

INVxp67_ASAP7_75t_L g128 ( 
.A(n_118),
.Y(n_128)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_119),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_L g119 ( 
.A(n_120),
.B(n_121),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_L g122 ( 
.A(n_123),
.B(n_124),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_L g136 ( 
.A(n_123),
.B(n_124),
.Y(n_136)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_125),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_L g129 ( 
.A(n_130),
.B(n_131),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_L g133 ( 
.A(n_134),
.B(n_135),
.Y(n_133)
);

CKINVDCx16_ASAP7_75t_R g139 ( 
.A(n_140),
.Y(n_139)
);

CKINVDCx20_ASAP7_75t_R g144 ( 
.A(n_145),
.Y(n_144)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_150),
.Y(n_149)
);

NOR2xp33_ASAP7_75t_L g153 ( 
.A(n_154),
.B(n_155),
.Y(n_153)
);

CKINVDCx20_ASAP7_75t_R g81 ( 
.A(n_158),
.Y(n_81)
);

INVxp67_ASAP7_75t_L g86 ( 
.A(n_159),
.Y(n_86)
);

INVxp67_ASAP7_75t_L g89 ( 
.A(n_160),
.Y(n_89)
);

CKINVDCx20_ASAP7_75t_R g95 ( 
.A(n_161),
.Y(n_95)
);

CKINVDCx20_ASAP7_75t_R g99 ( 
.A(n_162),
.Y(n_99)
);

CKINVDCx20_ASAP7_75t_R g102 ( 
.A(n_163),
.Y(n_102)
);

CKINVDCx20_ASAP7_75t_R g106 ( 
.A(n_164),
.Y(n_106)
);

CKINVDCx20_ASAP7_75t_R g111 ( 
.A(n_165),
.Y(n_111)
);

CKINVDCx20_ASAP7_75t_R g117 ( 
.A(n_166),
.Y(n_117)
);

CKINVDCx20_ASAP7_75t_R g126 ( 
.A(n_167),
.Y(n_126)
);


endmodule