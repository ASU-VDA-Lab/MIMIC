module fake_jpeg_24761_n_332 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_332);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_332;

wire n_253;
wire n_330;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_15;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

BUFx6f_ASAP7_75t_L g15 ( 
.A(n_12),
.Y(n_15)
);

BUFx24_ASAP7_75t_L g16 ( 
.A(n_12),
.Y(n_16)
);

CKINVDCx14_ASAP7_75t_R g17 ( 
.A(n_8),
.Y(n_17)
);

BUFx5_ASAP7_75t_L g18 ( 
.A(n_8),
.Y(n_18)
);

BUFx5_ASAP7_75t_L g19 ( 
.A(n_12),
.Y(n_19)
);

BUFx3_ASAP7_75t_L g20 ( 
.A(n_5),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_13),
.Y(n_21)
);

INVx2_ASAP7_75t_L g22 ( 
.A(n_13),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_5),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_10),
.Y(n_24)
);

INVx8_ASAP7_75t_L g25 ( 
.A(n_6),
.Y(n_25)
);

BUFx16f_ASAP7_75t_L g26 ( 
.A(n_6),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_3),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_7),
.Y(n_28)
);

INVx5_ASAP7_75t_L g29 ( 
.A(n_2),
.Y(n_29)
);

INVx2_ASAP7_75t_L g30 ( 
.A(n_1),
.Y(n_30)
);

INVx8_ASAP7_75t_L g31 ( 
.A(n_23),
.Y(n_31)
);

INVx2_ASAP7_75t_L g43 ( 
.A(n_31),
.Y(n_43)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_16),
.Y(n_32)
);

NAND2xp5_ASAP7_75t_L g57 ( 
.A(n_32),
.B(n_26),
.Y(n_57)
);

INVx8_ASAP7_75t_L g33 ( 
.A(n_23),
.Y(n_33)
);

INVx2_ASAP7_75t_L g47 ( 
.A(n_33),
.Y(n_47)
);

INVx4_ASAP7_75t_SL g34 ( 
.A(n_16),
.Y(n_34)
);

CKINVDCx6p67_ASAP7_75t_R g53 ( 
.A(n_34),
.Y(n_53)
);

INVx3_ASAP7_75t_L g35 ( 
.A(n_16),
.Y(n_35)
);

INVx8_ASAP7_75t_L g51 ( 
.A(n_35),
.Y(n_51)
);

BUFx12f_ASAP7_75t_L g36 ( 
.A(n_16),
.Y(n_36)
);

BUFx12f_ASAP7_75t_L g44 ( 
.A(n_36),
.Y(n_44)
);

INVx11_ASAP7_75t_L g37 ( 
.A(n_30),
.Y(n_37)
);

INVx4_ASAP7_75t_L g52 ( 
.A(n_37),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_20),
.Y(n_38)
);

INVx6_ASAP7_75t_L g48 ( 
.A(n_38),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_20),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_39),
.Y(n_45)
);

INVx2_ASAP7_75t_L g40 ( 
.A(n_25),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g42 ( 
.A(n_40),
.B(n_30),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g41 ( 
.A(n_26),
.B(n_0),
.Y(n_41)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_41),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_SL g75 ( 
.A(n_42),
.B(n_61),
.Y(n_75)
);

INVx5_ASAP7_75t_L g46 ( 
.A(n_36),
.Y(n_46)
);

INVx4_ASAP7_75t_L g68 ( 
.A(n_46),
.Y(n_68)
);

INVx3_ASAP7_75t_L g49 ( 
.A(n_37),
.Y(n_49)
);

INVx5_ASAP7_75t_L g82 ( 
.A(n_49),
.Y(n_82)
);

INVx5_ASAP7_75t_L g54 ( 
.A(n_36),
.Y(n_54)
);

INVx4_ASAP7_75t_L g83 ( 
.A(n_54),
.Y(n_83)
);

INVx4_ASAP7_75t_L g55 ( 
.A(n_37),
.Y(n_55)
);

AOI22xp33_ASAP7_75t_SL g87 ( 
.A1(n_55),
.A2(n_34),
.B1(n_35),
.B2(n_36),
.Y(n_87)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_36),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_56),
.Y(n_66)
);

AND2x2_ASAP7_75t_L g79 ( 
.A(n_57),
.B(n_59),
.Y(n_79)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_36),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g88 ( 
.A(n_58),
.Y(n_88)
);

CKINVDCx14_ASAP7_75t_R g59 ( 
.A(n_41),
.Y(n_59)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_41),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_L g65 ( 
.A(n_60),
.B(n_62),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_35),
.B(n_26),
.Y(n_61)
);

CKINVDCx16_ASAP7_75t_R g62 ( 
.A(n_38),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_35),
.B(n_21),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_L g86 ( 
.A(n_63),
.B(n_32),
.Y(n_86)
);

INVx2_ASAP7_75t_L g64 ( 
.A(n_51),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_64),
.B(n_71),
.Y(n_99)
);

OA22x2_ASAP7_75t_L g67 ( 
.A1(n_53),
.A2(n_36),
.B1(n_34),
.B2(n_18),
.Y(n_67)
);

OAI22xp5_ASAP7_75t_L g106 ( 
.A1(n_67),
.A2(n_87),
.B1(n_54),
.B2(n_48),
.Y(n_106)
);

CKINVDCx9p33_ASAP7_75t_R g69 ( 
.A(n_53),
.Y(n_69)
);

INVx1_ASAP7_75t_SL g108 ( 
.A(n_69),
.Y(n_108)
);

BUFx2_ASAP7_75t_L g70 ( 
.A(n_53),
.Y(n_70)
);

CKINVDCx16_ASAP7_75t_R g114 ( 
.A(n_70),
.Y(n_114)
);

INVx2_ASAP7_75t_L g71 ( 
.A(n_51),
.Y(n_71)
);

A2O1A1Ixp33_ASAP7_75t_L g72 ( 
.A1(n_57),
.A2(n_17),
.B(n_21),
.C(n_38),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_SL g93 ( 
.A(n_72),
.B(n_80),
.Y(n_93)
);

INVx2_ASAP7_75t_L g73 ( 
.A(n_53),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_73),
.B(n_74),
.Y(n_101)
);

INVx3_ASAP7_75t_L g74 ( 
.A(n_45),
.Y(n_74)
);

BUFx12_ASAP7_75t_L g76 ( 
.A(n_44),
.Y(n_76)
);

INVx2_ASAP7_75t_L g91 ( 
.A(n_76),
.Y(n_91)
);

BUFx12f_ASAP7_75t_L g77 ( 
.A(n_44),
.Y(n_77)
);

INVxp67_ASAP7_75t_L g103 ( 
.A(n_77),
.Y(n_103)
);

INVx2_ASAP7_75t_L g78 ( 
.A(n_44),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_78),
.B(n_81),
.Y(n_107)
);

AND2x2_ASAP7_75t_L g80 ( 
.A(n_50),
.B(n_36),
.Y(n_80)
);

CKINVDCx12_ASAP7_75t_R g81 ( 
.A(n_44),
.Y(n_81)
);

INVx2_ASAP7_75t_L g84 ( 
.A(n_45),
.Y(n_84)
);

HB1xp67_ASAP7_75t_L g113 ( 
.A(n_84),
.Y(n_113)
);

INVx4_ASAP7_75t_L g85 ( 
.A(n_46),
.Y(n_85)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_85),
.Y(n_92)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_86),
.Y(n_94)
);

INVx3_ASAP7_75t_L g89 ( 
.A(n_77),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g116 ( 
.A(n_89),
.B(n_76),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_L g90 ( 
.A(n_79),
.B(n_80),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_L g118 ( 
.A(n_90),
.B(n_96),
.Y(n_118)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_65),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g125 ( 
.A(n_95),
.B(n_102),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_L g96 ( 
.A(n_79),
.B(n_60),
.Y(n_96)
);

INVx2_ASAP7_75t_L g97 ( 
.A(n_76),
.Y(n_97)
);

INVx6_ASAP7_75t_L g138 ( 
.A(n_97),
.Y(n_138)
);

OR2x2_ASAP7_75t_L g98 ( 
.A(n_67),
.B(n_34),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g119 ( 
.A(n_98),
.B(n_100),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_SL g100 ( 
.A(n_75),
.B(n_50),
.Y(n_100)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_70),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_L g104 ( 
.A(n_72),
.B(n_48),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_L g120 ( 
.A(n_104),
.B(n_105),
.Y(n_120)
);

OR2x2_ASAP7_75t_L g105 ( 
.A(n_67),
.B(n_34),
.Y(n_105)
);

INVxp67_ASAP7_75t_L g121 ( 
.A(n_106),
.Y(n_121)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_68),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_109),
.B(n_110),
.Y(n_128)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_68),
.Y(n_110)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_83),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_L g132 ( 
.A(n_111),
.B(n_82),
.Y(n_132)
);

MAJIxp5_ASAP7_75t_L g112 ( 
.A(n_77),
.B(n_32),
.C(n_18),
.Y(n_112)
);

XOR2xp5_ASAP7_75t_L g141 ( 
.A(n_112),
.B(n_19),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_SL g115 ( 
.A(n_95),
.B(n_40),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_L g143 ( 
.A(n_115),
.B(n_127),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_SL g163 ( 
.A(n_116),
.B(n_123),
.Y(n_163)
);

MAJx2_ASAP7_75t_L g117 ( 
.A(n_90),
.B(n_19),
.C(n_87),
.Y(n_117)
);

MAJx2_ASAP7_75t_L g165 ( 
.A(n_117),
.B(n_39),
.C(n_29),
.Y(n_165)
);

CKINVDCx20_ASAP7_75t_R g122 ( 
.A(n_99),
.Y(n_122)
);

CKINVDCx20_ASAP7_75t_R g148 ( 
.A(n_122),
.Y(n_148)
);

INVx1_ASAP7_75t_SL g123 ( 
.A(n_108),
.Y(n_123)
);

INVx5_ASAP7_75t_L g124 ( 
.A(n_113),
.Y(n_124)
);

AOI22xp33_ASAP7_75t_SL g147 ( 
.A1(n_124),
.A2(n_130),
.B1(n_139),
.B2(n_102),
.Y(n_147)
);

CKINVDCx20_ASAP7_75t_R g126 ( 
.A(n_99),
.Y(n_126)
);

CKINVDCx20_ASAP7_75t_R g157 ( 
.A(n_126),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_93),
.B(n_82),
.Y(n_127)
);

OAI22xp5_ASAP7_75t_L g129 ( 
.A1(n_104),
.A2(n_43),
.B1(n_47),
.B2(n_33),
.Y(n_129)
);

AOI22xp5_ASAP7_75t_L g153 ( 
.A1(n_129),
.A2(n_131),
.B1(n_31),
.B2(n_33),
.Y(n_153)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_101),
.Y(n_130)
);

OAI22xp5_ASAP7_75t_SL g131 ( 
.A1(n_93),
.A2(n_47),
.B1(n_43),
.B2(n_40),
.Y(n_131)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_132),
.Y(n_151)
);

INVxp67_ASAP7_75t_L g133 ( 
.A(n_107),
.Y(n_133)
);

INVxp33_ASAP7_75t_L g160 ( 
.A(n_133),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_L g134 ( 
.A(n_96),
.B(n_49),
.Y(n_134)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_134),
.Y(n_155)
);

AND2x6_ASAP7_75t_L g135 ( 
.A(n_98),
.B(n_10),
.Y(n_135)
);

XNOR2xp5_ASAP7_75t_L g146 ( 
.A(n_135),
.B(n_107),
.Y(n_146)
);

INVx3_ASAP7_75t_L g136 ( 
.A(n_114),
.Y(n_136)
);

INVx11_ASAP7_75t_L g145 ( 
.A(n_136),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_L g137 ( 
.A(n_100),
.B(n_38),
.Y(n_137)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_137),
.Y(n_158)
);

CKINVDCx16_ASAP7_75t_R g139 ( 
.A(n_101),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_L g140 ( 
.A(n_114),
.B(n_85),
.Y(n_140)
);

AOI22xp33_ASAP7_75t_L g164 ( 
.A1(n_140),
.A2(n_108),
.B1(n_55),
.B2(n_52),
.Y(n_164)
);

MAJIxp5_ASAP7_75t_L g144 ( 
.A(n_141),
.B(n_112),
.C(n_94),
.Y(n_144)
);

OAI22xp33_ASAP7_75t_L g142 ( 
.A1(n_121),
.A2(n_106),
.B1(n_83),
.B2(n_105),
.Y(n_142)
);

OAI22xp5_ASAP7_75t_SL g189 ( 
.A1(n_142),
.A2(n_156),
.B1(n_167),
.B2(n_139),
.Y(n_189)
);

XNOR2xp5_ASAP7_75t_L g172 ( 
.A(n_144),
.B(n_161),
.Y(n_172)
);

NOR2xp33_ASAP7_75t_L g174 ( 
.A(n_146),
.B(n_141),
.Y(n_174)
);

OAI22xp5_ASAP7_75t_L g186 ( 
.A1(n_147),
.A2(n_152),
.B1(n_153),
.B2(n_159),
.Y(n_186)
);

AOI22xp5_ASAP7_75t_SL g149 ( 
.A1(n_127),
.A2(n_105),
.B1(n_98),
.B2(n_94),
.Y(n_149)
);

OAI22xp5_ASAP7_75t_L g194 ( 
.A1(n_149),
.A2(n_164),
.B1(n_124),
.B2(n_69),
.Y(n_194)
);

AOI21xp5_ASAP7_75t_L g150 ( 
.A1(n_120),
.A2(n_111),
.B(n_110),
.Y(n_150)
);

OAI21xp5_ASAP7_75t_SL g173 ( 
.A1(n_150),
.A2(n_154),
.B(n_162),
.Y(n_173)
);

OAI22xp5_ASAP7_75t_L g152 ( 
.A1(n_120),
.A2(n_31),
.B1(n_33),
.B2(n_40),
.Y(n_152)
);

XOR2x2_ASAP7_75t_L g154 ( 
.A(n_117),
.B(n_37),
.Y(n_154)
);

OAI22xp5_ASAP7_75t_SL g156 ( 
.A1(n_119),
.A2(n_31),
.B1(n_33),
.B2(n_74),
.Y(n_156)
);

OAI22xp5_ASAP7_75t_L g159 ( 
.A1(n_134),
.A2(n_31),
.B1(n_22),
.B2(n_37),
.Y(n_159)
);

XNOR2xp5_ASAP7_75t_L g161 ( 
.A(n_118),
.B(n_38),
.Y(n_161)
);

AOI21xp5_ASAP7_75t_L g162 ( 
.A1(n_119),
.A2(n_109),
.B(n_92),
.Y(n_162)
);

OAI21xp5_ASAP7_75t_SL g180 ( 
.A1(n_165),
.A2(n_137),
.B(n_115),
.Y(n_180)
);

XNOR2xp5_ASAP7_75t_L g166 ( 
.A(n_118),
.B(n_39),
.Y(n_166)
);

XNOR2xp5_ASAP7_75t_L g179 ( 
.A(n_166),
.B(n_129),
.Y(n_179)
);

OAI22xp5_ASAP7_75t_SL g167 ( 
.A1(n_117),
.A2(n_52),
.B1(n_92),
.B2(n_22),
.Y(n_167)
);

AND2x2_ASAP7_75t_L g168 ( 
.A(n_167),
.B(n_131),
.Y(n_168)
);

OAI21xp5_ASAP7_75t_SL g217 ( 
.A1(n_168),
.A2(n_171),
.B(n_177),
.Y(n_217)
);

INVx4_ASAP7_75t_L g169 ( 
.A(n_145),
.Y(n_169)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_169),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_L g170 ( 
.A(n_155),
.B(n_122),
.Y(n_170)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_170),
.Y(n_205)
);

HAxp5_ASAP7_75t_SL g171 ( 
.A(n_154),
.B(n_126),
.CON(n_171),
.SN(n_171)
);

NOR2xp33_ASAP7_75t_L g197 ( 
.A(n_174),
.B(n_176),
.Y(n_197)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_150),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_L g201 ( 
.A(n_175),
.B(n_178),
.Y(n_201)
);

NOR2xp33_ASAP7_75t_SL g176 ( 
.A(n_148),
.B(n_125),
.Y(n_176)
);

AND2x6_ASAP7_75t_L g177 ( 
.A(n_146),
.B(n_135),
.Y(n_177)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_143),
.Y(n_178)
);

XNOR2xp5_ASAP7_75t_L g208 ( 
.A(n_179),
.B(n_39),
.Y(n_208)
);

XOR2xp5_ASAP7_75t_L g206 ( 
.A(n_180),
.B(n_185),
.Y(n_206)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_143),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_L g211 ( 
.A(n_181),
.B(n_191),
.Y(n_211)
);

INVx13_ASAP7_75t_L g182 ( 
.A(n_145),
.Y(n_182)
);

NOR2xp33_ASAP7_75t_L g213 ( 
.A(n_182),
.B(n_183),
.Y(n_213)
);

INVx13_ASAP7_75t_L g183 ( 
.A(n_160),
.Y(n_183)
);

INVx6_ASAP7_75t_L g184 ( 
.A(n_160),
.Y(n_184)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_184),
.Y(n_214)
);

XNOR2xp5_ASAP7_75t_L g185 ( 
.A(n_161),
.B(n_125),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_SL g187 ( 
.A(n_157),
.B(n_132),
.Y(n_187)
);

CKINVDCx16_ASAP7_75t_R g199 ( 
.A(n_187),
.Y(n_199)
);

NOR2xp33_ASAP7_75t_L g188 ( 
.A(n_166),
.B(n_138),
.Y(n_188)
);

INVxp67_ASAP7_75t_L g204 ( 
.A(n_188),
.Y(n_204)
);

AOI22xp5_ASAP7_75t_L g219 ( 
.A1(n_189),
.A2(n_194),
.B1(n_123),
.B2(n_25),
.Y(n_219)
);

NOR2xp33_ASAP7_75t_L g190 ( 
.A(n_162),
.B(n_138),
.Y(n_190)
);

INVxp67_ASAP7_75t_L g212 ( 
.A(n_190),
.Y(n_212)
);

INVx1_ASAP7_75t_SL g191 ( 
.A(n_163),
.Y(n_191)
);

OAI32xp33_ASAP7_75t_L g192 ( 
.A1(n_165),
.A2(n_130),
.A3(n_128),
.B1(n_39),
.B2(n_29),
.Y(n_192)
);

XOR2xp5_ASAP7_75t_L g215 ( 
.A(n_192),
.B(n_15),
.Y(n_215)
);

NAND2xp5_ASAP7_75t_SL g193 ( 
.A(n_151),
.B(n_128),
.Y(n_193)
);

CKINVDCx20_ASAP7_75t_R g207 ( 
.A(n_193),
.Y(n_207)
);

AOI21xp5_ASAP7_75t_L g195 ( 
.A1(n_175),
.A2(n_155),
.B(n_151),
.Y(n_195)
);

AOI21xp5_ASAP7_75t_L g232 ( 
.A1(n_195),
.A2(n_191),
.B(n_186),
.Y(n_232)
);

OAI22xp5_ASAP7_75t_SL g196 ( 
.A1(n_173),
.A2(n_149),
.B1(n_142),
.B2(n_158),
.Y(n_196)
);

AOI22xp5_ASAP7_75t_L g229 ( 
.A1(n_196),
.A2(n_218),
.B1(n_212),
.B2(n_205),
.Y(n_229)
);

OR2x2_ASAP7_75t_L g200 ( 
.A(n_183),
.B(n_156),
.Y(n_200)
);

NAND2xp5_ASAP7_75t_L g237 ( 
.A(n_200),
.B(n_56),
.Y(n_237)
);

MAJIxp5_ASAP7_75t_L g202 ( 
.A(n_172),
.B(n_144),
.C(n_158),
.Y(n_202)
);

MAJIxp5_ASAP7_75t_L g228 ( 
.A(n_202),
.B(n_185),
.C(n_179),
.Y(n_228)
);

NOR2x1_ASAP7_75t_L g203 ( 
.A(n_170),
.B(n_153),
.Y(n_203)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_203),
.Y(n_223)
);

XOR2xp5_ASAP7_75t_L g224 ( 
.A(n_208),
.B(n_172),
.Y(n_224)
);

CKINVDCx20_ASAP7_75t_R g209 ( 
.A(n_169),
.Y(n_209)
);

CKINVDCx20_ASAP7_75t_R g241 ( 
.A(n_209),
.Y(n_241)
);

OAI22xp5_ASAP7_75t_L g210 ( 
.A1(n_173),
.A2(n_138),
.B1(n_136),
.B2(n_89),
.Y(n_210)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_210),
.Y(n_225)
);

NAND2xp5_ASAP7_75t_SL g231 ( 
.A(n_215),
.B(n_168),
.Y(n_231)
);

NAND3xp33_ASAP7_75t_L g216 ( 
.A(n_177),
.B(n_14),
.C(n_13),
.Y(n_216)
);

NAND3xp33_ASAP7_75t_L g233 ( 
.A(n_216),
.B(n_11),
.C(n_14),
.Y(n_233)
);

XNOR2x1_ASAP7_75t_L g218 ( 
.A(n_171),
.B(n_103),
.Y(n_218)
);

XNOR2xp5_ASAP7_75t_SL g234 ( 
.A(n_218),
.B(n_58),
.Y(n_234)
);

OAI22xp5_ASAP7_75t_L g222 ( 
.A1(n_219),
.A2(n_203),
.B1(n_212),
.B2(n_220),
.Y(n_222)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_184),
.Y(n_220)
);

NAND2xp5_ASAP7_75t_L g226 ( 
.A(n_220),
.B(n_182),
.Y(n_226)
);

OAI22xp5_ASAP7_75t_SL g221 ( 
.A1(n_217),
.A2(n_178),
.B1(n_181),
.B2(n_180),
.Y(n_221)
);

AOI22xp5_ASAP7_75t_L g246 ( 
.A1(n_221),
.A2(n_222),
.B1(n_227),
.B2(n_240),
.Y(n_246)
);

XOR2xp5_ASAP7_75t_L g258 ( 
.A(n_224),
.B(n_235),
.Y(n_258)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_226),
.Y(n_245)
);

OAI22xp5_ASAP7_75t_SL g227 ( 
.A1(n_217),
.A2(n_189),
.B1(n_168),
.B2(n_192),
.Y(n_227)
);

MAJIxp5_ASAP7_75t_L g244 ( 
.A(n_228),
.B(n_238),
.C(n_196),
.Y(n_244)
);

OAI22xp5_ASAP7_75t_SL g248 ( 
.A1(n_229),
.A2(n_233),
.B1(n_219),
.B2(n_207),
.Y(n_248)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_211),
.Y(n_230)
);

NAND2xp5_ASAP7_75t_SL g260 ( 
.A(n_230),
.B(n_231),
.Y(n_260)
);

OAI21xp5_ASAP7_75t_L g243 ( 
.A1(n_232),
.A2(n_195),
.B(n_201),
.Y(n_243)
);

XNOR2xp5_ASAP7_75t_SL g249 ( 
.A(n_234),
.B(n_200),
.Y(n_249)
);

XNOR2xp5_ASAP7_75t_L g235 ( 
.A(n_206),
.B(n_97),
.Y(n_235)
);

XNOR2xp5_ASAP7_75t_L g236 ( 
.A(n_206),
.B(n_91),
.Y(n_236)
);

XNOR2xp5_ASAP7_75t_L g250 ( 
.A(n_236),
.B(n_208),
.Y(n_250)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_237),
.Y(n_256)
);

XOR2xp5_ASAP7_75t_L g238 ( 
.A(n_202),
.B(n_91),
.Y(n_238)
);

NAND2xp5_ASAP7_75t_L g239 ( 
.A(n_199),
.B(n_9),
.Y(n_239)
);

CKINVDCx14_ASAP7_75t_R g254 ( 
.A(n_239),
.Y(n_254)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_211),
.Y(n_240)
);

NAND2xp5_ASAP7_75t_SL g242 ( 
.A(n_204),
.B(n_9),
.Y(n_242)
);

CKINVDCx14_ASAP7_75t_R g261 ( 
.A(n_242),
.Y(n_261)
);

AOI21xp5_ASAP7_75t_L g272 ( 
.A1(n_243),
.A2(n_234),
.B(n_1),
.Y(n_272)
);

MAJIxp5_ASAP7_75t_L g274 ( 
.A(n_244),
.B(n_247),
.C(n_253),
.Y(n_274)
);

MAJIxp5_ASAP7_75t_L g247 ( 
.A(n_238),
.B(n_205),
.C(n_201),
.Y(n_247)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_248),
.Y(n_270)
);

XNOR2xp5_ASAP7_75t_L g263 ( 
.A(n_249),
.B(n_252),
.Y(n_263)
);

XNOR2xp5_ASAP7_75t_L g271 ( 
.A(n_250),
.B(n_251),
.Y(n_271)
);

XNOR2xp5_ASAP7_75t_SL g251 ( 
.A(n_221),
.B(n_197),
.Y(n_251)
);

XNOR2xp5_ASAP7_75t_L g252 ( 
.A(n_224),
.B(n_215),
.Y(n_252)
);

MAJIxp5_ASAP7_75t_L g253 ( 
.A(n_228),
.B(n_214),
.C(n_204),
.Y(n_253)
);

AOI22xp5_ASAP7_75t_L g255 ( 
.A1(n_225),
.A2(n_214),
.B1(n_198),
.B2(n_213),
.Y(n_255)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_255),
.Y(n_273)
);

AOI22xp5_ASAP7_75t_L g257 ( 
.A1(n_223),
.A2(n_24),
.B1(n_15),
.B2(n_28),
.Y(n_257)
);

NAND2xp5_ASAP7_75t_L g266 ( 
.A(n_257),
.B(n_262),
.Y(n_266)
);

AO22x1_ASAP7_75t_L g259 ( 
.A1(n_232),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_259)
);

AOI21xp5_ASAP7_75t_SL g275 ( 
.A1(n_259),
.A2(n_0),
.B(n_1),
.Y(n_275)
);

CKINVDCx16_ASAP7_75t_R g262 ( 
.A(n_237),
.Y(n_262)
);

AND2x2_ASAP7_75t_L g264 ( 
.A(n_252),
.B(n_227),
.Y(n_264)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_264),
.Y(n_290)
);

OA21x2_ASAP7_75t_SL g265 ( 
.A1(n_251),
.A2(n_236),
.B(n_235),
.Y(n_265)
);

AOI22xp5_ASAP7_75t_SL g283 ( 
.A1(n_265),
.A2(n_250),
.B1(n_258),
.B2(n_254),
.Y(n_283)
);

INVx1_ASAP7_75t_SL g267 ( 
.A(n_260),
.Y(n_267)
);

INVx4_ASAP7_75t_L g292 ( 
.A(n_267),
.Y(n_292)
);

XNOR2xp5_ASAP7_75t_L g268 ( 
.A(n_258),
.B(n_229),
.Y(n_268)
);

XNOR2xp5_ASAP7_75t_L g284 ( 
.A(n_268),
.B(n_24),
.Y(n_284)
);

NAND2xp5_ASAP7_75t_L g269 ( 
.A(n_261),
.B(n_241),
.Y(n_269)
);

NAND2xp5_ASAP7_75t_L g285 ( 
.A(n_269),
.B(n_275),
.Y(n_285)
);

XOR2xp5_ASAP7_75t_L g281 ( 
.A(n_272),
.B(n_249),
.Y(n_281)
);

NAND2xp5_ASAP7_75t_L g276 ( 
.A(n_245),
.B(n_9),
.Y(n_276)
);

NAND2xp5_ASAP7_75t_L g294 ( 
.A(n_276),
.B(n_278),
.Y(n_294)
);

MAJIxp5_ASAP7_75t_L g277 ( 
.A(n_253),
.B(n_88),
.C(n_66),
.Y(n_277)
);

MAJIxp5_ASAP7_75t_L g282 ( 
.A(n_277),
.B(n_256),
.C(n_244),
.Y(n_282)
);

AND2x2_ASAP7_75t_L g278 ( 
.A(n_247),
.B(n_243),
.Y(n_278)
);

CKINVDCx20_ASAP7_75t_R g279 ( 
.A(n_246),
.Y(n_279)
);

NOR2xp33_ASAP7_75t_SL g280 ( 
.A(n_279),
.B(n_259),
.Y(n_280)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_280),
.Y(n_297)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_281),
.Y(n_300)
);

MAJIxp5_ASAP7_75t_L g307 ( 
.A(n_282),
.B(n_286),
.C(n_289),
.Y(n_307)
);

XOR2xp5_ASAP7_75t_L g295 ( 
.A(n_283),
.B(n_284),
.Y(n_295)
);

MAJIxp5_ASAP7_75t_L g286 ( 
.A(n_274),
.B(n_88),
.C(n_66),
.Y(n_286)
);

NOR2xp33_ASAP7_75t_L g287 ( 
.A(n_267),
.B(n_14),
.Y(n_287)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_287),
.Y(n_302)
);

OAI22xp5_ASAP7_75t_L g288 ( 
.A1(n_270),
.A2(n_11),
.B1(n_10),
.B2(n_3),
.Y(n_288)
);

AOI22xp5_ASAP7_75t_L g304 ( 
.A1(n_288),
.A2(n_3),
.B1(n_4),
.B2(n_5),
.Y(n_304)
);

MAJIxp5_ASAP7_75t_L g289 ( 
.A(n_274),
.B(n_0),
.C(n_2),
.Y(n_289)
);

XOR2xp5_ASAP7_75t_L g291 ( 
.A(n_271),
.B(n_11),
.Y(n_291)
);

NAND2xp5_ASAP7_75t_L g298 ( 
.A(n_291),
.B(n_275),
.Y(n_298)
);

AOI22xp5_ASAP7_75t_SL g293 ( 
.A1(n_273),
.A2(n_264),
.B1(n_278),
.B2(n_266),
.Y(n_293)
);

NOR2xp33_ASAP7_75t_L g296 ( 
.A(n_293),
.B(n_277),
.Y(n_296)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_296),
.Y(n_310)
);

NAND2xp5_ASAP7_75t_L g314 ( 
.A(n_298),
.B(n_301),
.Y(n_314)
);

AOI21xp5_ASAP7_75t_L g299 ( 
.A1(n_290),
.A2(n_271),
.B(n_263),
.Y(n_299)
);

MAJIxp5_ASAP7_75t_L g309 ( 
.A(n_299),
.B(n_289),
.C(n_291),
.Y(n_309)
);

NAND2xp5_ASAP7_75t_L g301 ( 
.A(n_285),
.B(n_28),
.Y(n_301)
);

FAx1_ASAP7_75t_SL g303 ( 
.A(n_281),
.B(n_2),
.CI(n_3),
.CON(n_303),
.SN(n_303)
);

NAND2xp5_ASAP7_75t_L g316 ( 
.A(n_303),
.B(n_304),
.Y(n_316)
);

AOI22xp33_ASAP7_75t_SL g305 ( 
.A1(n_292),
.A2(n_4),
.B1(n_5),
.B2(n_6),
.Y(n_305)
);

AOI22xp5_ASAP7_75t_L g312 ( 
.A1(n_305),
.A2(n_302),
.B1(n_297),
.B2(n_300),
.Y(n_312)
);

NAND2xp5_ASAP7_75t_L g306 ( 
.A(n_294),
.B(n_292),
.Y(n_306)
);

NOR2xp33_ASAP7_75t_SL g315 ( 
.A(n_306),
.B(n_4),
.Y(n_315)
);

MAJIxp5_ASAP7_75t_L g308 ( 
.A(n_307),
.B(n_282),
.C(n_286),
.Y(n_308)
);

MAJIxp5_ASAP7_75t_L g321 ( 
.A(n_308),
.B(n_309),
.C(n_311),
.Y(n_321)
);

MAJIxp5_ASAP7_75t_L g311 ( 
.A(n_307),
.B(n_27),
.C(n_6),
.Y(n_311)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_312),
.Y(n_319)
);

XOR2xp5_ASAP7_75t_L g313 ( 
.A(n_295),
.B(n_27),
.Y(n_313)
);

MAJIxp5_ASAP7_75t_L g322 ( 
.A(n_313),
.B(n_295),
.C(n_305),
.Y(n_322)
);

NAND2xp5_ASAP7_75t_SL g320 ( 
.A(n_315),
.B(n_303),
.Y(n_320)
);

INVxp67_ASAP7_75t_L g317 ( 
.A(n_308),
.Y(n_317)
);

OAI21xp5_ASAP7_75t_SL g325 ( 
.A1(n_317),
.A2(n_322),
.B(n_323),
.Y(n_325)
);

NOR2xp33_ASAP7_75t_L g318 ( 
.A(n_310),
.B(n_304),
.Y(n_318)
);

NOR2xp33_ASAP7_75t_SL g326 ( 
.A(n_318),
.B(n_320),
.Y(n_326)
);

NOR2xp33_ASAP7_75t_L g323 ( 
.A(n_316),
.B(n_314),
.Y(n_323)
);

OAI21x1_ASAP7_75t_L g324 ( 
.A1(n_321),
.A2(n_313),
.B(n_7),
.Y(n_324)
);

MAJIxp5_ASAP7_75t_L g327 ( 
.A(n_324),
.B(n_319),
.C(n_7),
.Y(n_327)
);

NOR2xp67_ASAP7_75t_SL g328 ( 
.A(n_327),
.B(n_326),
.Y(n_328)
);

OAI21xp5_ASAP7_75t_L g329 ( 
.A1(n_328),
.A2(n_317),
.B(n_325),
.Y(n_329)
);

NAND2xp5_ASAP7_75t_SL g330 ( 
.A(n_329),
.B(n_4),
.Y(n_330)
);

XOR2xp5_ASAP7_75t_L g331 ( 
.A(n_330),
.B(n_7),
.Y(n_331)
);

AOI21xp5_ASAP7_75t_L g332 ( 
.A1(n_331),
.A2(n_8),
.B(n_302),
.Y(n_332)
);


endmodule