module fake_jpeg_2625_n_175 (n_13, n_21, n_33, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_40, n_19, n_18, n_20, n_35, n_41, n_4, n_34, n_30, n_39, n_42, n_16, n_3, n_0, n_24, n_28, n_38, n_26, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_12, n_32, n_8, n_15, n_7, n_175);

input n_13;
input n_21;
input n_33;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_42;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_175;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_59;
wire n_84;
wire n_98;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_155;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_57;
wire n_171;
wire n_119;
wire n_69;
wire n_83;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_168;
wire n_106;
wire n_111;
wire n_44;
wire n_143;
wire n_75;
wire n_122;
wire n_102;
wire n_121;
wire n_99;
wire n_130;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_91;
wire n_54;
wire n_93;
wire n_161;
wire n_138;
wire n_101;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_62;
wire n_167;
wire n_174;
wire n_120;
wire n_43;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

INVx1_ASAP7_75t_L g43 ( 
.A(n_39),
.Y(n_43)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_38),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_1),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_0),
.Y(n_46)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_15),
.Y(n_47)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_0),
.Y(n_48)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_36),
.Y(n_49)
);

INVx2_ASAP7_75t_L g50 ( 
.A(n_37),
.Y(n_50)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_12),
.Y(n_51)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_42),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_41),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_16),
.Y(n_54)
);

CKINVDCx20_ASAP7_75t_R g55 ( 
.A(n_27),
.Y(n_55)
);

BUFx10_ASAP7_75t_L g56 ( 
.A(n_28),
.Y(n_56)
);

INVx1_ASAP7_75t_SL g57 ( 
.A(n_22),
.Y(n_57)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_40),
.Y(n_58)
);

BUFx5_ASAP7_75t_L g59 ( 
.A(n_10),
.Y(n_59)
);

INVx11_ASAP7_75t_L g60 ( 
.A(n_56),
.Y(n_60)
);

INVx4_ASAP7_75t_L g72 ( 
.A(n_60),
.Y(n_72)
);

CKINVDCx20_ASAP7_75t_R g61 ( 
.A(n_49),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_61),
.B(n_62),
.Y(n_74)
);

OR2x2_ASAP7_75t_L g62 ( 
.A(n_47),
.B(n_1),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_53),
.Y(n_63)
);

INVx6_ASAP7_75t_L g69 ( 
.A(n_63),
.Y(n_69)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_53),
.Y(n_64)
);

INVx8_ASAP7_75t_L g68 ( 
.A(n_64),
.Y(n_68)
);

INVx6_ASAP7_75t_SL g65 ( 
.A(n_56),
.Y(n_65)
);

INVx3_ASAP7_75t_L g77 ( 
.A(n_65),
.Y(n_77)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_50),
.Y(n_66)
);

INVx2_ASAP7_75t_L g75 ( 
.A(n_66),
.Y(n_75)
);

AOI22xp33_ASAP7_75t_L g67 ( 
.A1(n_63),
.A2(n_45),
.B1(n_46),
.B2(n_47),
.Y(n_67)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_67),
.Y(n_81)
);

INVx3_ASAP7_75t_L g70 ( 
.A(n_65),
.Y(n_70)
);

INVx2_ASAP7_75t_L g94 ( 
.A(n_70),
.Y(n_94)
);

INVx3_ASAP7_75t_L g71 ( 
.A(n_65),
.Y(n_71)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_71),
.Y(n_83)
);

AOI22xp33_ASAP7_75t_SL g73 ( 
.A1(n_60),
.A2(n_50),
.B1(n_57),
.B2(n_59),
.Y(n_73)
);

CKINVDCx16_ASAP7_75t_R g82 ( 
.A(n_73),
.Y(n_82)
);

INVx2_ASAP7_75t_L g76 ( 
.A(n_66),
.Y(n_76)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_76),
.Y(n_93)
);

INVx4_ASAP7_75t_L g78 ( 
.A(n_60),
.Y(n_78)
);

BUFx6f_ASAP7_75t_L g84 ( 
.A(n_78),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_74),
.B(n_61),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_L g96 ( 
.A(n_79),
.B(n_80),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_70),
.B(n_62),
.Y(n_80)
);

MAJIxp5_ASAP7_75t_L g85 ( 
.A(n_75),
.B(n_43),
.C(n_58),
.Y(n_85)
);

MAJIxp5_ASAP7_75t_L g105 ( 
.A(n_85),
.B(n_57),
.C(n_48),
.Y(n_105)
);

NOR2x1_ASAP7_75t_L g86 ( 
.A(n_71),
.B(n_62),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g112 ( 
.A(n_86),
.B(n_92),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_L g87 ( 
.A(n_77),
.B(n_43),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_87),
.B(n_90),
.Y(n_99)
);

BUFx6f_ASAP7_75t_L g88 ( 
.A(n_69),
.Y(n_88)
);

INVx3_ASAP7_75t_L g102 ( 
.A(n_88),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_SL g89 ( 
.A(n_72),
.B(n_49),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_SL g114 ( 
.A(n_89),
.B(n_91),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g90 ( 
.A(n_69),
.B(n_58),
.Y(n_90)
);

CKINVDCx20_ASAP7_75t_R g91 ( 
.A(n_68),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_SL g92 ( 
.A(n_72),
.B(n_51),
.Y(n_92)
);

CKINVDCx16_ASAP7_75t_R g95 ( 
.A(n_78),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g100 ( 
.A(n_95),
.B(n_44),
.Y(n_100)
);

OAI22xp5_ASAP7_75t_SL g97 ( 
.A1(n_81),
.A2(n_73),
.B1(n_64),
.B2(n_63),
.Y(n_97)
);

AOI22xp5_ASAP7_75t_L g115 ( 
.A1(n_97),
.A2(n_98),
.B1(n_103),
.B2(n_88),
.Y(n_115)
);

OAI22xp33_ASAP7_75t_SL g98 ( 
.A1(n_82),
.A2(n_64),
.B1(n_63),
.B2(n_45),
.Y(n_98)
);

CKINVDCx14_ASAP7_75t_R g126 ( 
.A(n_100),
.Y(n_126)
);

AOI22xp5_ASAP7_75t_L g101 ( 
.A1(n_90),
.A2(n_64),
.B1(n_68),
.B2(n_46),
.Y(n_101)
);

OAI22xp5_ASAP7_75t_L g116 ( 
.A1(n_101),
.A2(n_106),
.B1(n_54),
.B2(n_84),
.Y(n_116)
);

OAI21xp33_ASAP7_75t_L g103 ( 
.A1(n_86),
.A2(n_55),
.B(n_52),
.Y(n_103)
);

OAI21xp5_ASAP7_75t_L g120 ( 
.A1(n_103),
.A2(n_3),
.B(n_4),
.Y(n_120)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_83),
.Y(n_104)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_104),
.Y(n_123)
);

XNOR2xp5_ASAP7_75t_L g118 ( 
.A(n_105),
.B(n_2),
.Y(n_118)
);

AOI22xp5_ASAP7_75t_L g106 ( 
.A1(n_87),
.A2(n_54),
.B1(n_56),
.B2(n_59),
.Y(n_106)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_83),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_L g124 ( 
.A(n_107),
.B(n_108),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_L g108 ( 
.A(n_85),
.B(n_2),
.Y(n_108)
);

INVxp67_ASAP7_75t_L g109 ( 
.A(n_93),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_L g125 ( 
.A(n_109),
.B(n_111),
.Y(n_125)
);

OR2x2_ASAP7_75t_SL g110 ( 
.A(n_93),
.B(n_56),
.Y(n_110)
);

OAI21xp5_ASAP7_75t_SL g130 ( 
.A1(n_110),
.A2(n_3),
.B(n_5),
.Y(n_130)
);

INVxp67_ASAP7_75t_L g111 ( 
.A(n_94),
.Y(n_111)
);

BUFx24_ASAP7_75t_SL g113 ( 
.A(n_94),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_L g133 ( 
.A(n_113),
.B(n_23),
.Y(n_133)
);

AOI22xp5_ASAP7_75t_L g135 ( 
.A1(n_115),
.A2(n_116),
.B1(n_131),
.B2(n_6),
.Y(n_135)
);

INVx4_ASAP7_75t_L g117 ( 
.A(n_102),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_L g136 ( 
.A(n_117),
.B(n_121),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_L g147 ( 
.A(n_118),
.B(n_128),
.Y(n_147)
);

AOI22xp5_ASAP7_75t_L g119 ( 
.A1(n_99),
.A2(n_84),
.B1(n_4),
.B2(n_5),
.Y(n_119)
);

OAI22xp5_ASAP7_75t_SL g137 ( 
.A1(n_119),
.A2(n_122),
.B1(n_7),
.B2(n_8),
.Y(n_137)
);

OAI21xp5_ASAP7_75t_SL g139 ( 
.A1(n_120),
.A2(n_124),
.B(n_129),
.Y(n_139)
);

INVxp67_ASAP7_75t_L g121 ( 
.A(n_114),
.Y(n_121)
);

AOI22xp33_ASAP7_75t_L g122 ( 
.A1(n_102),
.A2(n_109),
.B1(n_112),
.B2(n_111),
.Y(n_122)
);

XNOR2xp5_ASAP7_75t_L g127 ( 
.A(n_96),
.B(n_20),
.Y(n_127)
);

XNOR2xp5_ASAP7_75t_L g144 ( 
.A(n_127),
.B(n_129),
.Y(n_144)
);

CKINVDCx14_ASAP7_75t_R g128 ( 
.A(n_105),
.Y(n_128)
);

XNOR2xp5_ASAP7_75t_SL g129 ( 
.A(n_110),
.B(n_19),
.Y(n_129)
);

INVxp67_ASAP7_75t_L g148 ( 
.A(n_130),
.Y(n_148)
);

OAI22xp5_ASAP7_75t_SL g131 ( 
.A1(n_99),
.A2(n_6),
.B1(n_7),
.B2(n_8),
.Y(n_131)
);

INVxp67_ASAP7_75t_L g132 ( 
.A(n_114),
.Y(n_132)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_132),
.Y(n_145)
);

BUFx24_ASAP7_75t_SL g146 ( 
.A(n_133),
.Y(n_146)
);

CKINVDCx20_ASAP7_75t_R g134 ( 
.A(n_125),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_L g152 ( 
.A(n_134),
.B(n_137),
.Y(n_152)
);

HB1xp67_ASAP7_75t_L g155 ( 
.A(n_135),
.Y(n_155)
);

AOI22xp5_ASAP7_75t_L g138 ( 
.A1(n_121),
.A2(n_9),
.B1(n_10),
.B2(n_11),
.Y(n_138)
);

OAI22xp5_ASAP7_75t_SL g151 ( 
.A1(n_138),
.A2(n_141),
.B1(n_143),
.B2(n_29),
.Y(n_151)
);

AOI21x1_ASAP7_75t_L g156 ( 
.A1(n_139),
.A2(n_142),
.B(n_34),
.Y(n_156)
);

AOI22xp5_ASAP7_75t_L g140 ( 
.A1(n_132),
.A2(n_9),
.B1(n_11),
.B2(n_12),
.Y(n_140)
);

AOI22xp5_ASAP7_75t_L g149 ( 
.A1(n_140),
.A2(n_18),
.B1(n_21),
.B2(n_24),
.Y(n_149)
);

AOI22xp5_ASAP7_75t_L g141 ( 
.A1(n_123),
.A2(n_13),
.B1(n_14),
.B2(n_15),
.Y(n_141)
);

OAI21xp5_ASAP7_75t_L g142 ( 
.A1(n_122),
.A2(n_126),
.B(n_117),
.Y(n_142)
);

AOI22xp33_ASAP7_75t_L g143 ( 
.A1(n_127),
.A2(n_13),
.B1(n_14),
.B2(n_17),
.Y(n_143)
);

OAI22xp5_ASAP7_75t_SL g163 ( 
.A1(n_149),
.A2(n_150),
.B1(n_154),
.B2(n_148),
.Y(n_163)
);

AOI21xp5_ASAP7_75t_L g150 ( 
.A1(n_142),
.A2(n_25),
.B(n_26),
.Y(n_150)
);

AOI22xp5_ASAP7_75t_SL g161 ( 
.A1(n_151),
.A2(n_148),
.B1(n_138),
.B2(n_141),
.Y(n_161)
);

NOR2xp33_ASAP7_75t_L g153 ( 
.A(n_145),
.B(n_30),
.Y(n_153)
);

XNOR2xp5_ASAP7_75t_L g159 ( 
.A(n_153),
.B(n_156),
.Y(n_159)
);

AOI22xp5_ASAP7_75t_L g154 ( 
.A1(n_136),
.A2(n_31),
.B1(n_32),
.B2(n_33),
.Y(n_154)
);

CKINVDCx20_ASAP7_75t_R g157 ( 
.A(n_146),
.Y(n_157)
);

BUFx5_ASAP7_75t_L g160 ( 
.A(n_157),
.Y(n_160)
);

MAJIxp5_ASAP7_75t_L g158 ( 
.A(n_155),
.B(n_147),
.C(n_144),
.Y(n_158)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_158),
.Y(n_165)
);

OAI22xp5_ASAP7_75t_SL g164 ( 
.A1(n_161),
.A2(n_162),
.B1(n_163),
.B2(n_154),
.Y(n_164)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_152),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_L g168 ( 
.A(n_164),
.B(n_166),
.Y(n_168)
);

OAI21xp5_ASAP7_75t_L g166 ( 
.A1(n_158),
.A2(n_151),
.B(n_149),
.Y(n_166)
);

OAI21xp5_ASAP7_75t_SL g167 ( 
.A1(n_165),
.A2(n_159),
.B(n_160),
.Y(n_167)
);

BUFx6f_ASAP7_75t_L g169 ( 
.A(n_167),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_L g170 ( 
.A(n_169),
.B(n_168),
.Y(n_170)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_170),
.Y(n_171)
);

INVxp67_ASAP7_75t_L g172 ( 
.A(n_171),
.Y(n_172)
);

OAI21xp5_ASAP7_75t_L g173 ( 
.A1(n_172),
.A2(n_166),
.B(n_144),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_L g174 ( 
.A(n_173),
.B(n_160),
.Y(n_174)
);

XOR2xp5_ASAP7_75t_L g175 ( 
.A(n_174),
.B(n_35),
.Y(n_175)
);


endmodule