module fake_jpeg_10063_n_343 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_343);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_343;

wire n_253;
wire n_330;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_340;
wire n_291;
wire n_236;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

BUFx6f_ASAP7_75t_L g16 ( 
.A(n_9),
.Y(n_16)
);

BUFx5_ASAP7_75t_L g17 ( 
.A(n_10),
.Y(n_17)
);

INVx3_ASAP7_75t_L g18 ( 
.A(n_14),
.Y(n_18)
);

BUFx12f_ASAP7_75t_L g19 ( 
.A(n_4),
.Y(n_19)
);

INVx2_ASAP7_75t_SL g20 ( 
.A(n_1),
.Y(n_20)
);

BUFx12_ASAP7_75t_L g21 ( 
.A(n_6),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_14),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_12),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_14),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_9),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_13),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_2),
.Y(n_27)
);

BUFx16f_ASAP7_75t_L g28 ( 
.A(n_15),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_12),
.Y(n_29)
);

BUFx3_ASAP7_75t_L g30 ( 
.A(n_2),
.Y(n_30)
);

BUFx12f_ASAP7_75t_L g31 ( 
.A(n_1),
.Y(n_31)
);

BUFx12f_ASAP7_75t_L g32 ( 
.A(n_11),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_12),
.Y(n_33)
);

INVx2_ASAP7_75t_L g34 ( 
.A(n_5),
.Y(n_34)
);

BUFx3_ASAP7_75t_L g35 ( 
.A(n_7),
.Y(n_35)
);

INVx13_ASAP7_75t_L g36 ( 
.A(n_13),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g37 ( 
.A(n_22),
.B(n_26),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_37),
.B(n_39),
.Y(n_53)
);

INVx5_ASAP7_75t_L g38 ( 
.A(n_36),
.Y(n_38)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_38),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_L g39 ( 
.A(n_22),
.B(n_0),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_31),
.Y(n_40)
);

INVx6_ASAP7_75t_L g58 ( 
.A(n_40),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_31),
.Y(n_41)
);

INVx3_ASAP7_75t_L g67 ( 
.A(n_41),
.Y(n_67)
);

HB1xp67_ASAP7_75t_L g42 ( 
.A(n_21),
.Y(n_42)
);

INVx2_ASAP7_75t_L g59 ( 
.A(n_42),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_31),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_43),
.Y(n_52)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_28),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g57 ( 
.A(n_44),
.B(n_46),
.Y(n_57)
);

INVx2_ASAP7_75t_L g45 ( 
.A(n_28),
.Y(n_45)
);

HB1xp67_ASAP7_75t_L g63 ( 
.A(n_45),
.Y(n_63)
);

INVx2_ASAP7_75t_L g46 ( 
.A(n_28),
.Y(n_46)
);

INVx2_ASAP7_75t_L g47 ( 
.A(n_28),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_47),
.B(n_48),
.Y(n_61)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_17),
.Y(n_48)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_39),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_L g98 ( 
.A(n_49),
.B(n_51),
.Y(n_98)
);

INVx2_ASAP7_75t_SL g50 ( 
.A(n_38),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_50),
.B(n_19),
.Y(n_71)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_45),
.Y(n_51)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_46),
.Y(n_54)
);

AND2x2_ASAP7_75t_L g83 ( 
.A(n_54),
.B(n_60),
.Y(n_83)
);

AOI22xp33_ASAP7_75t_SL g55 ( 
.A1(n_47),
.A2(n_18),
.B1(n_34),
.B2(n_20),
.Y(n_55)
);

AOI22xp33_ASAP7_75t_SL g94 ( 
.A1(n_55),
.A2(n_65),
.B1(n_27),
.B2(n_16),
.Y(n_94)
);

AND2x2_ASAP7_75t_L g60 ( 
.A(n_44),
.B(n_36),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_48),
.B(n_25),
.Y(n_62)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_62),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_40),
.B(n_25),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_SL g76 ( 
.A(n_64),
.B(n_66),
.Y(n_76)
);

AOI22xp33_ASAP7_75t_SL g65 ( 
.A1(n_40),
.A2(n_18),
.B1(n_34),
.B2(n_20),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_41),
.B(n_24),
.Y(n_66)
);

INVx6_ASAP7_75t_L g68 ( 
.A(n_52),
.Y(n_68)
);

CKINVDCx20_ASAP7_75t_R g135 ( 
.A(n_68),
.Y(n_135)
);

INVx2_ASAP7_75t_L g69 ( 
.A(n_63),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_69),
.B(n_73),
.Y(n_110)
);

AO22x1_ASAP7_75t_L g70 ( 
.A1(n_60),
.A2(n_17),
.B1(n_20),
.B2(n_36),
.Y(n_70)
);

AND2x4_ASAP7_75t_L g111 ( 
.A(n_70),
.B(n_55),
.Y(n_111)
);

CKINVDCx16_ASAP7_75t_R g130 ( 
.A(n_71),
.Y(n_130)
);

AOI22xp5_ASAP7_75t_L g72 ( 
.A1(n_49),
.A2(n_24),
.B1(n_23),
.B2(n_29),
.Y(n_72)
);

OAI22xp5_ASAP7_75t_L g131 ( 
.A1(n_72),
.A2(n_87),
.B1(n_100),
.B2(n_33),
.Y(n_131)
);

INVx2_ASAP7_75t_L g73 ( 
.A(n_63),
.Y(n_73)
);

INVx2_ASAP7_75t_SL g74 ( 
.A(n_50),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g119 ( 
.A(n_74),
.B(n_75),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_62),
.B(n_29),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_61),
.B(n_23),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g120 ( 
.A(n_77),
.B(n_79),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_SL g78 ( 
.A(n_53),
.B(n_26),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_SL g115 ( 
.A(n_78),
.B(n_81),
.Y(n_115)
);

INVx3_ASAP7_75t_L g79 ( 
.A(n_52),
.Y(n_79)
);

BUFx6f_ASAP7_75t_L g80 ( 
.A(n_52),
.Y(n_80)
);

INVx3_ASAP7_75t_L g117 ( 
.A(n_80),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_SL g81 ( 
.A(n_53),
.B(n_21),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_61),
.B(n_66),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g122 ( 
.A(n_82),
.B(n_84),
.Y(n_122)
);

INVx3_ASAP7_75t_L g84 ( 
.A(n_52),
.Y(n_84)
);

AND2x2_ASAP7_75t_SL g85 ( 
.A(n_51),
.B(n_43),
.Y(n_85)
);

AND2x2_ASAP7_75t_L g125 ( 
.A(n_85),
.B(n_104),
.Y(n_125)
);

CKINVDCx20_ASAP7_75t_R g86 ( 
.A(n_64),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_86),
.B(n_88),
.Y(n_124)
);

AOI22xp33_ASAP7_75t_L g87 ( 
.A1(n_58),
.A2(n_27),
.B1(n_16),
.B2(n_33),
.Y(n_87)
);

CKINVDCx16_ASAP7_75t_R g88 ( 
.A(n_57),
.Y(n_88)
);

INVx4_ASAP7_75t_L g89 ( 
.A(n_67),
.Y(n_89)
);

INVx8_ASAP7_75t_L g126 ( 
.A(n_89),
.Y(n_126)
);

INVx3_ASAP7_75t_L g90 ( 
.A(n_50),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g133 ( 
.A(n_90),
.B(n_91),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_57),
.B(n_19),
.Y(n_91)
);

BUFx12f_ASAP7_75t_L g92 ( 
.A(n_50),
.Y(n_92)
);

INVxp67_ASAP7_75t_L g121 ( 
.A(n_92),
.Y(n_121)
);

INVx3_ASAP7_75t_L g93 ( 
.A(n_56),
.Y(n_93)
);

INVx2_ASAP7_75t_L g109 ( 
.A(n_93),
.Y(n_109)
);

OAI22xp33_ASAP7_75t_SL g127 ( 
.A1(n_94),
.A2(n_102),
.B1(n_105),
.B2(n_65),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_SL g95 ( 
.A(n_54),
.B(n_43),
.Y(n_95)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_95),
.Y(n_112)
);

INVx2_ASAP7_75t_L g96 ( 
.A(n_56),
.Y(n_96)
);

INVx2_ASAP7_75t_L g116 ( 
.A(n_96),
.Y(n_116)
);

INVx2_ASAP7_75t_L g99 ( 
.A(n_67),
.Y(n_99)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_99),
.Y(n_128)
);

AOI22xp33_ASAP7_75t_L g100 ( 
.A1(n_58),
.A2(n_27),
.B1(n_16),
.B2(n_33),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_SL g101 ( 
.A(n_60),
.B(n_41),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_L g106 ( 
.A(n_101),
.B(n_70),
.Y(n_106)
);

INVx2_ASAP7_75t_L g102 ( 
.A(n_67),
.Y(n_102)
);

INVx4_ASAP7_75t_L g103 ( 
.A(n_58),
.Y(n_103)
);

OAI22xp33_ASAP7_75t_L g134 ( 
.A1(n_103),
.A2(n_35),
.B1(n_30),
.B2(n_32),
.Y(n_134)
);

AND2x2_ASAP7_75t_L g104 ( 
.A(n_60),
.B(n_0),
.Y(n_104)
);

INVx2_ASAP7_75t_SL g105 ( 
.A(n_59),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_SL g148 ( 
.A(n_106),
.B(n_0),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_L g107 ( 
.A(n_98),
.B(n_59),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_L g154 ( 
.A(n_107),
.B(n_108),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_L g108 ( 
.A(n_83),
.B(n_31),
.Y(n_108)
);

OAI21xp5_ASAP7_75t_SL g140 ( 
.A1(n_111),
.A2(n_85),
.B(n_97),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_L g113 ( 
.A(n_83),
.B(n_31),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_L g156 ( 
.A(n_113),
.B(n_114),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_L g114 ( 
.A(n_83),
.B(n_32),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g118 ( 
.A(n_104),
.B(n_32),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_L g157 ( 
.A(n_118),
.B(n_123),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_L g123 ( 
.A(n_104),
.B(n_72),
.Y(n_123)
);

AOI22xp33_ASAP7_75t_L g137 ( 
.A1(n_127),
.A2(n_131),
.B1(n_134),
.B2(n_93),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_L g129 ( 
.A(n_76),
.B(n_32),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_L g164 ( 
.A(n_129),
.B(n_132),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_L g132 ( 
.A(n_85),
.B(n_32),
.Y(n_132)
);

BUFx2_ASAP7_75t_L g136 ( 
.A(n_126),
.Y(n_136)
);

CKINVDCx16_ASAP7_75t_R g175 ( 
.A(n_136),
.Y(n_175)
);

OAI22xp5_ASAP7_75t_L g181 ( 
.A1(n_137),
.A2(n_160),
.B1(n_161),
.B2(n_126),
.Y(n_181)
);

INVxp67_ASAP7_75t_L g138 ( 
.A(n_110),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_L g169 ( 
.A(n_138),
.B(n_141),
.Y(n_169)
);

NOR2xp33_ASAP7_75t_L g139 ( 
.A(n_109),
.B(n_105),
.Y(n_139)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_139),
.Y(n_171)
);

XNOR2xp5_ASAP7_75t_SL g173 ( 
.A(n_140),
.B(n_114),
.Y(n_173)
);

NOR2xp33_ASAP7_75t_SL g141 ( 
.A(n_115),
.B(n_11),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_L g142 ( 
.A(n_109),
.B(n_69),
.Y(n_142)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_142),
.Y(n_172)
);

O2A1O1Ixp33_ASAP7_75t_SL g143 ( 
.A1(n_111),
.A2(n_102),
.B(n_99),
.C(n_89),
.Y(n_143)
);

OAI21xp5_ASAP7_75t_SL g167 ( 
.A1(n_143),
.A2(n_132),
.B(n_106),
.Y(n_167)
);

NOR2xp33_ASAP7_75t_L g144 ( 
.A(n_120),
.B(n_73),
.Y(n_144)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_144),
.Y(n_178)
);

INVx2_ASAP7_75t_L g145 ( 
.A(n_116),
.Y(n_145)
);

AOI22xp33_ASAP7_75t_SL g196 ( 
.A1(n_145),
.A2(n_117),
.B1(n_135),
.B2(n_116),
.Y(n_196)
);

BUFx6f_ASAP7_75t_L g146 ( 
.A(n_117),
.Y(n_146)
);

BUFx6f_ASAP7_75t_L g186 ( 
.A(n_146),
.Y(n_186)
);

MAJIxp5_ASAP7_75t_L g147 ( 
.A(n_108),
.B(n_103),
.C(n_96),
.Y(n_147)
);

XNOR2xp5_ASAP7_75t_L g198 ( 
.A(n_147),
.B(n_165),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_L g187 ( 
.A(n_148),
.B(n_149),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_SL g149 ( 
.A(n_115),
.B(n_68),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_SL g150 ( 
.A(n_107),
.B(n_13),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_L g190 ( 
.A(n_150),
.B(n_151),
.Y(n_190)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_122),
.Y(n_151)
);

OAI22xp5_ASAP7_75t_SL g152 ( 
.A1(n_111),
.A2(n_84),
.B1(n_79),
.B2(n_90),
.Y(n_152)
);

AOI22xp5_ASAP7_75t_L g185 ( 
.A1(n_152),
.A2(n_135),
.B1(n_128),
.B2(n_131),
.Y(n_185)
);

NOR2xp33_ASAP7_75t_L g153 ( 
.A(n_112),
.B(n_74),
.Y(n_153)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_153),
.Y(n_184)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_124),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_L g168 ( 
.A(n_155),
.B(n_159),
.Y(n_168)
);

NOR3xp33_ASAP7_75t_L g158 ( 
.A(n_123),
.B(n_35),
.C(n_30),
.Y(n_158)
);

NAND3xp33_ASAP7_75t_L g197 ( 
.A(n_158),
.B(n_92),
.C(n_11),
.Y(n_197)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_133),
.Y(n_159)
);

AOI22xp33_ASAP7_75t_SL g160 ( 
.A1(n_111),
.A2(n_9),
.B1(n_15),
.B2(n_2),
.Y(n_160)
);

AOI22xp33_ASAP7_75t_SL g161 ( 
.A1(n_111),
.A2(n_10),
.B1(n_15),
.B2(n_3),
.Y(n_161)
);

BUFx2_ASAP7_75t_L g162 ( 
.A(n_126),
.Y(n_162)
);

CKINVDCx20_ASAP7_75t_R g188 ( 
.A(n_162),
.Y(n_188)
);

AND2x6_ASAP7_75t_L g163 ( 
.A(n_125),
.B(n_10),
.Y(n_163)
);

BUFx2_ASAP7_75t_L g170 ( 
.A(n_163),
.Y(n_170)
);

MAJIxp5_ASAP7_75t_L g165 ( 
.A(n_113),
.B(n_92),
.C(n_80),
.Y(n_165)
);

NAND2x1_ASAP7_75t_SL g166 ( 
.A(n_143),
.B(n_125),
.Y(n_166)
);

OAI21xp5_ASAP7_75t_SL g201 ( 
.A1(n_166),
.A2(n_177),
.B(n_179),
.Y(n_201)
);

AOI21xp5_ASAP7_75t_L g220 ( 
.A1(n_167),
.A2(n_176),
.B(n_182),
.Y(n_220)
);

XOR2xp5_ASAP7_75t_L g219 ( 
.A(n_173),
.B(n_199),
.Y(n_219)
);

NAND2xp5_ASAP7_75t_L g174 ( 
.A(n_154),
.B(n_129),
.Y(n_174)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_174),
.Y(n_200)
);

AND2x2_ASAP7_75t_L g176 ( 
.A(n_147),
.B(n_125),
.Y(n_176)
);

INVxp67_ASAP7_75t_L g177 ( 
.A(n_152),
.Y(n_177)
);

INVxp67_ASAP7_75t_L g179 ( 
.A(n_165),
.Y(n_179)
);

OAI21xp5_ASAP7_75t_L g180 ( 
.A1(n_157),
.A2(n_118),
.B(n_130),
.Y(n_180)
);

OAI21xp5_ASAP7_75t_L g230 ( 
.A1(n_180),
.A2(n_121),
.B(n_19),
.Y(n_230)
);

INVxp67_ASAP7_75t_L g222 ( 
.A(n_181),
.Y(n_222)
);

OAI21xp5_ASAP7_75t_SL g182 ( 
.A1(n_143),
.A2(n_130),
.B(n_112),
.Y(n_182)
);

INVxp33_ASAP7_75t_L g183 ( 
.A(n_136),
.Y(n_183)
);

NOR2xp33_ASAP7_75t_L g203 ( 
.A(n_183),
.B(n_191),
.Y(n_203)
);

OAI22xp5_ASAP7_75t_L g212 ( 
.A1(n_185),
.A2(n_138),
.B1(n_159),
.B2(n_151),
.Y(n_212)
);

INVxp67_ASAP7_75t_L g189 ( 
.A(n_136),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_L g204 ( 
.A(n_189),
.B(n_146),
.Y(n_204)
);

CKINVDCx20_ASAP7_75t_R g191 ( 
.A(n_162),
.Y(n_191)
);

INVx1_ASAP7_75t_SL g192 ( 
.A(n_164),
.Y(n_192)
);

NOR2xp33_ASAP7_75t_L g207 ( 
.A(n_192),
.B(n_193),
.Y(n_207)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_164),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_L g194 ( 
.A(n_154),
.B(n_119),
.Y(n_194)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_194),
.Y(n_205)
);

NAND2xp5_ASAP7_75t_L g195 ( 
.A(n_157),
.B(n_119),
.Y(n_195)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_195),
.Y(n_208)
);

INVxp67_ASAP7_75t_L g228 ( 
.A(n_196),
.Y(n_228)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_197),
.Y(n_211)
);

XNOR2xp5_ASAP7_75t_L g199 ( 
.A(n_140),
.B(n_156),
.Y(n_199)
);

CKINVDCx20_ASAP7_75t_R g202 ( 
.A(n_168),
.Y(n_202)
);

NAND2xp5_ASAP7_75t_L g233 ( 
.A(n_202),
.B(n_206),
.Y(n_233)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_204),
.Y(n_236)
);

CKINVDCx5p33_ASAP7_75t_R g206 ( 
.A(n_183),
.Y(n_206)
);

AND2x2_ASAP7_75t_L g209 ( 
.A(n_199),
.B(n_166),
.Y(n_209)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_209),
.Y(n_237)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_168),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_L g254 ( 
.A(n_210),
.B(n_217),
.Y(n_254)
);

NAND2xp5_ASAP7_75t_SL g251 ( 
.A(n_212),
.B(n_221),
.Y(n_251)
);

NAND2xp5_ASAP7_75t_L g213 ( 
.A(n_194),
.B(n_192),
.Y(n_213)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_213),
.Y(n_242)
);

NOR2xp33_ASAP7_75t_L g214 ( 
.A(n_188),
.B(n_184),
.Y(n_214)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_214),
.Y(n_243)
);

NAND2xp5_ASAP7_75t_L g215 ( 
.A(n_195),
.B(n_156),
.Y(n_215)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_215),
.Y(n_255)
);

AND2x2_ASAP7_75t_L g216 ( 
.A(n_198),
.B(n_163),
.Y(n_216)
);

AND2x2_ASAP7_75t_L g244 ( 
.A(n_216),
.B(n_226),
.Y(n_244)
);

CKINVDCx20_ASAP7_75t_R g217 ( 
.A(n_190),
.Y(n_217)
);

NAND2xp5_ASAP7_75t_L g218 ( 
.A(n_174),
.B(n_155),
.Y(n_218)
);

NAND2xp5_ASAP7_75t_L g240 ( 
.A(n_218),
.B(n_223),
.Y(n_240)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_169),
.Y(n_221)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_185),
.Y(n_223)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_187),
.Y(n_224)
);

NAND2xp5_ASAP7_75t_L g249 ( 
.A(n_224),
.B(n_227),
.Y(n_249)
);

INVx13_ASAP7_75t_L g225 ( 
.A(n_186),
.Y(n_225)
);

INVx3_ASAP7_75t_L g235 ( 
.A(n_225),
.Y(n_235)
);

AND2x2_ASAP7_75t_L g226 ( 
.A(n_198),
.B(n_128),
.Y(n_226)
);

NAND2xp5_ASAP7_75t_L g227 ( 
.A(n_182),
.B(n_141),
.Y(n_227)
);

NOR2xp33_ASAP7_75t_L g229 ( 
.A(n_171),
.B(n_145),
.Y(n_229)
);

NOR2xp33_ASAP7_75t_L g250 ( 
.A(n_229),
.B(n_19),
.Y(n_250)
);

MAJx2_ASAP7_75t_L g232 ( 
.A(n_230),
.B(n_180),
.C(n_167),
.Y(n_232)
);

AOI22xp5_ASAP7_75t_L g231 ( 
.A1(n_223),
.A2(n_177),
.B1(n_179),
.B2(n_170),
.Y(n_231)
);

OAI22xp5_ASAP7_75t_SL g256 ( 
.A1(n_231),
.A2(n_245),
.B1(n_228),
.B2(n_210),
.Y(n_256)
);

XNOR2xp5_ASAP7_75t_SL g266 ( 
.A(n_232),
.B(n_241),
.Y(n_266)
);

MAJIxp5_ASAP7_75t_L g234 ( 
.A(n_219),
.B(n_173),
.C(n_176),
.Y(n_234)
);

XNOR2xp5_ASAP7_75t_L g262 ( 
.A(n_234),
.B(n_246),
.Y(n_262)
);

INVx1_ASAP7_75t_SL g238 ( 
.A(n_204),
.Y(n_238)
);

NAND2xp5_ASAP7_75t_L g269 ( 
.A(n_238),
.B(n_205),
.Y(n_269)
);

CKINVDCx20_ASAP7_75t_R g239 ( 
.A(n_203),
.Y(n_239)
);

NOR2xp33_ASAP7_75t_SL g270 ( 
.A(n_239),
.B(n_253),
.Y(n_270)
);

MAJx2_ASAP7_75t_L g241 ( 
.A(n_219),
.B(n_176),
.C(n_170),
.Y(n_241)
);

AOI22xp5_ASAP7_75t_L g245 ( 
.A1(n_222),
.A2(n_189),
.B1(n_178),
.B2(n_175),
.Y(n_245)
);

XNOR2xp5_ASAP7_75t_L g246 ( 
.A(n_220),
.B(n_172),
.Y(n_246)
);

MAJIxp5_ASAP7_75t_L g247 ( 
.A(n_201),
.B(n_186),
.C(n_121),
.Y(n_247)
);

XNOR2xp5_ASAP7_75t_L g265 ( 
.A(n_247),
.B(n_201),
.Y(n_265)
);

OAI22xp5_ASAP7_75t_SL g248 ( 
.A1(n_222),
.A2(n_35),
.B1(n_30),
.B2(n_19),
.Y(n_248)
);

AOI22xp5_ASAP7_75t_L g258 ( 
.A1(n_248),
.A2(n_228),
.B1(n_237),
.B2(n_225),
.Y(n_258)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_250),
.Y(n_257)
);

NOR2xp33_ASAP7_75t_L g252 ( 
.A(n_224),
.B(n_21),
.Y(n_252)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_252),
.Y(n_261)
);

CKINVDCx20_ASAP7_75t_R g253 ( 
.A(n_206),
.Y(n_253)
);

AOI22xp5_ASAP7_75t_L g285 ( 
.A1(n_256),
.A2(n_259),
.B1(n_276),
.B2(n_242),
.Y(n_285)
);

OAI22xp5_ASAP7_75t_SL g283 ( 
.A1(n_258),
.A2(n_271),
.B1(n_272),
.B2(n_247),
.Y(n_283)
);

OAI22xp5_ASAP7_75t_SL g259 ( 
.A1(n_231),
.A2(n_205),
.B1(n_208),
.B2(n_213),
.Y(n_259)
);

OAI21xp5_ASAP7_75t_SL g260 ( 
.A1(n_233),
.A2(n_220),
.B(n_236),
.Y(n_260)
);

AOI21xp5_ASAP7_75t_L g293 ( 
.A1(n_260),
.A2(n_273),
.B(n_274),
.Y(n_293)
);

NOR2xp33_ASAP7_75t_L g263 ( 
.A(n_235),
.B(n_218),
.Y(n_263)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_263),
.Y(n_282)
);

NOR2xp33_ASAP7_75t_L g264 ( 
.A(n_235),
.B(n_207),
.Y(n_264)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_264),
.Y(n_286)
);

MAJIxp5_ASAP7_75t_L g287 ( 
.A(n_265),
.B(n_238),
.C(n_215),
.Y(n_287)
);

NOR2xp33_ASAP7_75t_L g267 ( 
.A(n_243),
.B(n_200),
.Y(n_267)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_267),
.Y(n_289)
);

NOR2xp33_ASAP7_75t_L g268 ( 
.A(n_255),
.B(n_200),
.Y(n_268)
);

NAND2xp5_ASAP7_75t_L g277 ( 
.A(n_268),
.B(n_275),
.Y(n_277)
);

INVxp67_ASAP7_75t_L g279 ( 
.A(n_269),
.Y(n_279)
);

OAI22xp5_ASAP7_75t_L g271 ( 
.A1(n_245),
.A2(n_227),
.B1(n_208),
.B2(n_216),
.Y(n_271)
);

OAI22xp5_ASAP7_75t_L g272 ( 
.A1(n_251),
.A2(n_216),
.B1(n_211),
.B2(n_230),
.Y(n_272)
);

INVxp67_ASAP7_75t_L g273 ( 
.A(n_240),
.Y(n_273)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_254),
.Y(n_274)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_240),
.Y(n_275)
);

CKINVDCx14_ASAP7_75t_R g276 ( 
.A(n_249),
.Y(n_276)
);

XNOR2x1_ASAP7_75t_L g278 ( 
.A(n_266),
.B(n_241),
.Y(n_278)
);

XNOR2x1_ASAP7_75t_L g298 ( 
.A(n_278),
.B(n_209),
.Y(n_298)
);

XOR2xp5_ASAP7_75t_L g280 ( 
.A(n_266),
.B(n_234),
.Y(n_280)
);

XOR2xp5_ASAP7_75t_L g300 ( 
.A(n_280),
.B(n_281),
.Y(n_300)
);

XOR2xp5_ASAP7_75t_L g281 ( 
.A(n_262),
.B(n_246),
.Y(n_281)
);

AOI22xp5_ASAP7_75t_L g299 ( 
.A1(n_283),
.A2(n_256),
.B1(n_273),
.B2(n_257),
.Y(n_299)
);

XNOR2xp5_ASAP7_75t_L g284 ( 
.A(n_265),
.B(n_249),
.Y(n_284)
);

NOR2xp33_ASAP7_75t_SL g303 ( 
.A(n_284),
.B(n_290),
.Y(n_303)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_285),
.Y(n_308)
);

XNOR2xp5_ASAP7_75t_L g297 ( 
.A(n_287),
.B(n_259),
.Y(n_297)
);

MAJIxp5_ASAP7_75t_L g288 ( 
.A(n_262),
.B(n_226),
.C(n_244),
.Y(n_288)
);

OAI21xp5_ASAP7_75t_L g309 ( 
.A1(n_288),
.A2(n_291),
.B(n_21),
.Y(n_309)
);

XNOR2xp5_ASAP7_75t_L g290 ( 
.A(n_258),
.B(n_248),
.Y(n_290)
);

MAJIxp5_ASAP7_75t_L g291 ( 
.A(n_260),
.B(n_226),
.C(n_244),
.Y(n_291)
);

OAI22xp5_ASAP7_75t_L g292 ( 
.A1(n_274),
.A2(n_232),
.B1(n_209),
.B2(n_3),
.Y(n_292)
);

NAND2xp5_ASAP7_75t_SL g295 ( 
.A(n_292),
.B(n_294),
.Y(n_295)
);

NOR2xp33_ASAP7_75t_SL g294 ( 
.A(n_261),
.B(n_6),
.Y(n_294)
);

NOR2xp33_ASAP7_75t_L g296 ( 
.A(n_286),
.B(n_270),
.Y(n_296)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_296),
.Y(n_312)
);

XNOR2xp5_ASAP7_75t_L g310 ( 
.A(n_297),
.B(n_309),
.Y(n_310)
);

OAI22xp5_ASAP7_75t_SL g313 ( 
.A1(n_298),
.A2(n_299),
.B1(n_307),
.B2(n_291),
.Y(n_313)
);

CKINVDCx20_ASAP7_75t_R g301 ( 
.A(n_277),
.Y(n_301)
);

NOR2xp33_ASAP7_75t_SL g319 ( 
.A(n_301),
.B(n_306),
.Y(n_319)
);

NAND2xp5_ASAP7_75t_L g302 ( 
.A(n_282),
.B(n_269),
.Y(n_302)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_302),
.Y(n_314)
);

OR2x2_ASAP7_75t_L g304 ( 
.A(n_279),
.B(n_5),
.Y(n_304)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_304),
.Y(n_315)
);

OAI21xp33_ASAP7_75t_L g305 ( 
.A1(n_278),
.A2(n_5),
.B(n_8),
.Y(n_305)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_305),
.Y(n_316)
);

NOR2xp33_ASAP7_75t_L g306 ( 
.A(n_289),
.B(n_6),
.Y(n_306)
);

CKINVDCx20_ASAP7_75t_R g307 ( 
.A(n_293),
.Y(n_307)
);

XNOR2xp5_ASAP7_75t_L g311 ( 
.A(n_297),
.B(n_287),
.Y(n_311)
);

AND2x2_ASAP7_75t_L g328 ( 
.A(n_311),
.B(n_317),
.Y(n_328)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_313),
.Y(n_324)
);

MAJIxp5_ASAP7_75t_L g317 ( 
.A(n_300),
.B(n_281),
.C(n_288),
.Y(n_317)
);

OAI22xp5_ASAP7_75t_SL g318 ( 
.A1(n_308),
.A2(n_279),
.B1(n_295),
.B2(n_298),
.Y(n_318)
);

NAND2xp5_ASAP7_75t_SL g322 ( 
.A(n_318),
.B(n_305),
.Y(n_322)
);

AOI22xp5_ASAP7_75t_L g320 ( 
.A1(n_303),
.A2(n_280),
.B1(n_1),
.B2(n_0),
.Y(n_320)
);

OAI22xp5_ASAP7_75t_SL g327 ( 
.A1(n_320),
.A2(n_4),
.B1(n_7),
.B2(n_8),
.Y(n_327)
);

NOR2xp33_ASAP7_75t_L g321 ( 
.A(n_319),
.B(n_304),
.Y(n_321)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_321),
.Y(n_330)
);

NAND2xp5_ASAP7_75t_L g332 ( 
.A(n_322),
.B(n_323),
.Y(n_332)
);

NAND2xp5_ASAP7_75t_L g323 ( 
.A(n_312),
.B(n_300),
.Y(n_323)
);

NAND2xp5_ASAP7_75t_SL g325 ( 
.A(n_314),
.B(n_3),
.Y(n_325)
);

OAI21xp5_ASAP7_75t_L g329 ( 
.A1(n_325),
.A2(n_316),
.B(n_4),
.Y(n_329)
);

NOR2xp33_ASAP7_75t_L g326 ( 
.A(n_315),
.B(n_311),
.Y(n_326)
);

NAND2xp5_ASAP7_75t_L g333 ( 
.A(n_326),
.B(n_327),
.Y(n_333)
);

CKINVDCx20_ASAP7_75t_R g336 ( 
.A(n_329),
.Y(n_336)
);

XOR2xp5_ASAP7_75t_L g331 ( 
.A(n_328),
.B(n_317),
.Y(n_331)
);

MAJIxp5_ASAP7_75t_L g334 ( 
.A(n_331),
.B(n_332),
.C(n_324),
.Y(n_334)
);

INVxp67_ASAP7_75t_L g337 ( 
.A(n_334),
.Y(n_337)
);

NOR2xp33_ASAP7_75t_L g335 ( 
.A(n_330),
.B(n_325),
.Y(n_335)
);

INVx1_ASAP7_75t_L g338 ( 
.A(n_337),
.Y(n_338)
);

OAI21xp5_ASAP7_75t_L g339 ( 
.A1(n_338),
.A2(n_333),
.B(n_335),
.Y(n_339)
);

NOR3xp33_ASAP7_75t_L g340 ( 
.A(n_339),
.B(n_336),
.C(n_331),
.Y(n_340)
);

OAI21xp5_ASAP7_75t_L g341 ( 
.A1(n_340),
.A2(n_320),
.B(n_310),
.Y(n_341)
);

O2A1O1Ixp33_ASAP7_75t_SL g342 ( 
.A1(n_341),
.A2(n_310),
.B(n_7),
.C(n_8),
.Y(n_342)
);

XNOR2xp5_ASAP7_75t_L g343 ( 
.A(n_342),
.B(n_1),
.Y(n_343)
);


endmodule