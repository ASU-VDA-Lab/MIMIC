module fake_jpeg_4657_n_339 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_339);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_339;

wire n_253;
wire n_330;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_13),
.Y(n_16)
);

BUFx12f_ASAP7_75t_L g17 ( 
.A(n_15),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_0),
.Y(n_18)
);

BUFx5_ASAP7_75t_L g19 ( 
.A(n_0),
.Y(n_19)
);

INVx6_ASAP7_75t_L g20 ( 
.A(n_12),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_6),
.Y(n_21)
);

INVx2_ASAP7_75t_L g22 ( 
.A(n_15),
.Y(n_22)
);

BUFx10_ASAP7_75t_L g23 ( 
.A(n_8),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_14),
.Y(n_24)
);

BUFx4f_ASAP7_75t_L g25 ( 
.A(n_9),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_14),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_4),
.Y(n_27)
);

INVx11_ASAP7_75t_L g28 ( 
.A(n_6),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_10),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_9),
.Y(n_30)
);

BUFx12f_ASAP7_75t_L g31 ( 
.A(n_6),
.Y(n_31)
);

INVx13_ASAP7_75t_L g32 ( 
.A(n_8),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_8),
.Y(n_33)
);

BUFx12f_ASAP7_75t_L g34 ( 
.A(n_19),
.Y(n_34)
);

INVx6_ASAP7_75t_L g72 ( 
.A(n_34),
.Y(n_72)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_23),
.Y(n_35)
);

NAND2xp5_ASAP7_75t_L g52 ( 
.A(n_35),
.B(n_37),
.Y(n_52)
);

INVx3_ASAP7_75t_L g36 ( 
.A(n_25),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_36),
.B(n_24),
.Y(n_73)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_23),
.Y(n_37)
);

NOR2xp67_ASAP7_75t_L g38 ( 
.A(n_19),
.B(n_25),
.Y(n_38)
);

AOI21xp33_ASAP7_75t_SL g71 ( 
.A1(n_38),
.A2(n_25),
.B(n_23),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g39 ( 
.A(n_32),
.B(n_22),
.Y(n_39)
);

NAND2xp5_ASAP7_75t_SL g65 ( 
.A(n_39),
.B(n_43),
.Y(n_65)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_26),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g57 ( 
.A(n_40),
.Y(n_57)
);

BUFx5_ASAP7_75t_L g41 ( 
.A(n_19),
.Y(n_41)
);

CKINVDCx14_ASAP7_75t_R g64 ( 
.A(n_41),
.Y(n_64)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_23),
.Y(n_42)
);

NAND2xp5_ASAP7_75t_L g60 ( 
.A(n_42),
.B(n_23),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g43 ( 
.A(n_32),
.B(n_15),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g44 ( 
.A(n_32),
.B(n_14),
.Y(n_44)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_44),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g45 ( 
.A(n_32),
.B(n_13),
.Y(n_45)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_45),
.Y(n_54)
);

OR2x2_ASAP7_75t_L g46 ( 
.A(n_38),
.B(n_18),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_46),
.B(n_53),
.Y(n_81)
);

AOI22xp5_ASAP7_75t_L g47 ( 
.A1(n_38),
.A2(n_20),
.B1(n_22),
.B2(n_28),
.Y(n_47)
);

OAI22xp5_ASAP7_75t_SL g92 ( 
.A1(n_47),
.A2(n_44),
.B1(n_16),
.B2(n_30),
.Y(n_92)
);

INVx2_ASAP7_75t_L g48 ( 
.A(n_41),
.Y(n_48)
);

INVx8_ASAP7_75t_L g94 ( 
.A(n_48),
.Y(n_94)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_41),
.Y(n_50)
);

BUFx3_ASAP7_75t_L g90 ( 
.A(n_50),
.Y(n_90)
);

BUFx8_ASAP7_75t_L g51 ( 
.A(n_41),
.Y(n_51)
);

CKINVDCx16_ASAP7_75t_R g77 ( 
.A(n_51),
.Y(n_77)
);

INVx3_ASAP7_75t_L g53 ( 
.A(n_36),
.Y(n_53)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_39),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_55),
.B(n_56),
.Y(n_83)
);

INVx4_ASAP7_75t_L g56 ( 
.A(n_36),
.Y(n_56)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_36),
.Y(n_58)
);

INVx6_ASAP7_75t_L g79 ( 
.A(n_58),
.Y(n_79)
);

INVx2_ASAP7_75t_L g59 ( 
.A(n_35),
.Y(n_59)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_59),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_60),
.B(n_66),
.Y(n_88)
);

AOI22xp33_ASAP7_75t_SL g61 ( 
.A1(n_35),
.A2(n_20),
.B1(n_22),
.B2(n_28),
.Y(n_61)
);

AOI21xp5_ASAP7_75t_L g74 ( 
.A1(n_61),
.A2(n_63),
.B(n_45),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_L g62 ( 
.A(n_43),
.B(n_27),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_L g75 ( 
.A(n_62),
.B(n_67),
.Y(n_75)
);

AOI22xp33_ASAP7_75t_SL g63 ( 
.A1(n_37),
.A2(n_20),
.B1(n_28),
.B2(n_33),
.Y(n_63)
);

INVx4_ASAP7_75t_L g66 ( 
.A(n_37),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_L g67 ( 
.A(n_43),
.B(n_27),
.Y(n_67)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_39),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_L g97 ( 
.A(n_68),
.B(n_70),
.Y(n_97)
);

OAI22xp5_ASAP7_75t_L g69 ( 
.A1(n_42),
.A2(n_20),
.B1(n_18),
.B2(n_33),
.Y(n_69)
);

AOI22xp5_ASAP7_75t_L g78 ( 
.A1(n_69),
.A2(n_33),
.B1(n_26),
.B2(n_40),
.Y(n_78)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_45),
.Y(n_70)
);

O2A1O1Ixp33_ASAP7_75t_L g96 ( 
.A1(n_71),
.A2(n_69),
.B(n_65),
.C(n_46),
.Y(n_96)
);

CKINVDCx16_ASAP7_75t_R g89 ( 
.A(n_73),
.Y(n_89)
);

AOI22xp5_ASAP7_75t_SL g119 ( 
.A1(n_74),
.A2(n_29),
.B1(n_25),
.B2(n_72),
.Y(n_119)
);

OAI22xp5_ASAP7_75t_L g76 ( 
.A1(n_47),
.A2(n_42),
.B1(n_40),
.B2(n_18),
.Y(n_76)
);

AOI22xp5_ASAP7_75t_L g115 ( 
.A1(n_76),
.A2(n_92),
.B1(n_96),
.B2(n_54),
.Y(n_115)
);

OAI22xp33_ASAP7_75t_SL g124 ( 
.A1(n_78),
.A2(n_84),
.B1(n_99),
.B2(n_29),
.Y(n_124)
);

INVx3_ASAP7_75t_L g80 ( 
.A(n_56),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_80),
.B(n_85),
.Y(n_101)
);

AOI22xp33_ASAP7_75t_L g84 ( 
.A1(n_55),
.A2(n_16),
.B1(n_30),
.B2(n_26),
.Y(n_84)
);

INVx2_ASAP7_75t_L g85 ( 
.A(n_66),
.Y(n_85)
);

INVx2_ASAP7_75t_SL g86 ( 
.A(n_58),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g112 ( 
.A(n_86),
.B(n_24),
.Y(n_112)
);

CKINVDCx20_ASAP7_75t_R g87 ( 
.A(n_57),
.Y(n_87)
);

CKINVDCx20_ASAP7_75t_R g126 ( 
.A(n_87),
.Y(n_126)
);

INVx5_ASAP7_75t_L g91 ( 
.A(n_53),
.Y(n_91)
);

INVxp33_ASAP7_75t_L g122 ( 
.A(n_91),
.Y(n_122)
);

INVx2_ASAP7_75t_L g93 ( 
.A(n_59),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g113 ( 
.A(n_93),
.B(n_24),
.Y(n_113)
);

INVxp67_ASAP7_75t_L g95 ( 
.A(n_60),
.Y(n_95)
);

INVxp67_ASAP7_75t_L g106 ( 
.A(n_95),
.Y(n_106)
);

BUFx12f_ASAP7_75t_L g98 ( 
.A(n_51),
.Y(n_98)
);

INVx8_ASAP7_75t_L g102 ( 
.A(n_98),
.Y(n_102)
);

AOI22xp33_ASAP7_75t_L g99 ( 
.A1(n_68),
.A2(n_29),
.B1(n_25),
.B2(n_24),
.Y(n_99)
);

OAI22xp5_ASAP7_75t_SL g100 ( 
.A1(n_81),
.A2(n_46),
.B1(n_52),
.B2(n_54),
.Y(n_100)
);

AOI22xp5_ASAP7_75t_L g132 ( 
.A1(n_100),
.A2(n_104),
.B1(n_89),
.B2(n_86),
.Y(n_132)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_78),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g149 ( 
.A(n_103),
.B(n_105),
.Y(n_149)
);

OAI22xp5_ASAP7_75t_SL g104 ( 
.A1(n_81),
.A2(n_52),
.B1(n_70),
.B2(n_49),
.Y(n_104)
);

CKINVDCx16_ASAP7_75t_R g105 ( 
.A(n_88),
.Y(n_105)
);

INVx2_ASAP7_75t_L g107 ( 
.A(n_91),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_L g136 ( 
.A(n_107),
.B(n_109),
.Y(n_136)
);

MAJIxp5_ASAP7_75t_L g108 ( 
.A(n_88),
.B(n_64),
.C(n_49),
.Y(n_108)
);

MAJIxp5_ASAP7_75t_L g129 ( 
.A(n_108),
.B(n_120),
.C(n_123),
.Y(n_129)
);

INVx2_ASAP7_75t_L g109 ( 
.A(n_90),
.Y(n_109)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_97),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_L g153 ( 
.A(n_110),
.B(n_111),
.Y(n_153)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_97),
.Y(n_111)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_112),
.Y(n_130)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_113),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_L g114 ( 
.A(n_87),
.B(n_57),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g146 ( 
.A(n_114),
.B(n_117),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_SL g140 ( 
.A(n_115),
.B(n_118),
.Y(n_140)
);

INVx4_ASAP7_75t_L g116 ( 
.A(n_90),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_L g152 ( 
.A(n_116),
.B(n_121),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_SL g117 ( 
.A(n_75),
.B(n_92),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_L g118 ( 
.A(n_75),
.B(n_67),
.Y(n_118)
);

OAI21xp5_ASAP7_75t_L g148 ( 
.A1(n_119),
.A2(n_23),
.B(n_51),
.Y(n_148)
);

XOR2xp5_ASAP7_75t_L g120 ( 
.A(n_76),
.B(n_62),
.Y(n_120)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_83),
.Y(n_121)
);

AND2x2_ASAP7_75t_SL g123 ( 
.A(n_96),
.B(n_34),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_SL g139 ( 
.A(n_124),
.B(n_125),
.Y(n_139)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_83),
.Y(n_125)
);

XNOR2xp5_ASAP7_75t_L g127 ( 
.A(n_96),
.B(n_74),
.Y(n_127)
);

XNOR2xp5_ASAP7_75t_L g155 ( 
.A(n_127),
.B(n_34),
.Y(n_155)
);

INVx2_ASAP7_75t_L g128 ( 
.A(n_90),
.Y(n_128)
);

AOI22xp33_ASAP7_75t_SL g150 ( 
.A1(n_128),
.A2(n_51),
.B1(n_98),
.B2(n_50),
.Y(n_150)
);

OAI22xp5_ASAP7_75t_L g131 ( 
.A1(n_123),
.A2(n_89),
.B1(n_79),
.B2(n_86),
.Y(n_131)
);

AOI22xp5_ASAP7_75t_L g169 ( 
.A1(n_131),
.A2(n_142),
.B1(n_148),
.B2(n_151),
.Y(n_169)
);

OAI22xp5_ASAP7_75t_L g181 ( 
.A1(n_132),
.A2(n_21),
.B1(n_17),
.B2(n_31),
.Y(n_181)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_101),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_L g184 ( 
.A(n_134),
.B(n_143),
.Y(n_184)
);

MAJIxp5_ASAP7_75t_L g135 ( 
.A(n_123),
.B(n_120),
.C(n_108),
.Y(n_135)
);

MAJIxp5_ASAP7_75t_L g166 ( 
.A(n_135),
.B(n_126),
.C(n_112),
.Y(n_166)
);

AOI22xp5_ASAP7_75t_L g137 ( 
.A1(n_103),
.A2(n_79),
.B1(n_93),
.B2(n_82),
.Y(n_137)
);

OAI22xp5_ASAP7_75t_SL g174 ( 
.A1(n_137),
.A2(n_138),
.B1(n_141),
.B2(n_147),
.Y(n_174)
);

AOI22xp5_ASAP7_75t_L g138 ( 
.A1(n_123),
.A2(n_79),
.B1(n_82),
.B2(n_85),
.Y(n_138)
);

AOI22xp5_ASAP7_75t_L g141 ( 
.A1(n_117),
.A2(n_48),
.B1(n_80),
.B2(n_94),
.Y(n_141)
);

OAI22xp5_ASAP7_75t_L g142 ( 
.A1(n_127),
.A2(n_72),
.B1(n_94),
.B2(n_77),
.Y(n_142)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_114),
.Y(n_143)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_104),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_L g157 ( 
.A(n_144),
.B(n_156),
.Y(n_157)
);

CKINVDCx20_ASAP7_75t_R g145 ( 
.A(n_126),
.Y(n_145)
);

CKINVDCx20_ASAP7_75t_R g158 ( 
.A(n_145),
.Y(n_158)
);

AOI22xp5_ASAP7_75t_L g147 ( 
.A1(n_100),
.A2(n_94),
.B1(n_44),
.B2(n_77),
.Y(n_147)
);

CKINVDCx20_ASAP7_75t_R g163 ( 
.A(n_150),
.Y(n_163)
);

OAI22xp5_ASAP7_75t_SL g151 ( 
.A1(n_115),
.A2(n_21),
.B1(n_34),
.B2(n_31),
.Y(n_151)
);

AOI22xp5_ASAP7_75t_L g154 ( 
.A1(n_105),
.A2(n_21),
.B1(n_31),
.B2(n_34),
.Y(n_154)
);

OAI22xp5_ASAP7_75t_SL g179 ( 
.A1(n_154),
.A2(n_102),
.B1(n_116),
.B2(n_98),
.Y(n_179)
);

XNOR2xp5_ASAP7_75t_L g175 ( 
.A(n_155),
.B(n_34),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_SL g156 ( 
.A(n_118),
.B(n_0),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_L g159 ( 
.A(n_146),
.B(n_111),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_L g189 ( 
.A(n_159),
.B(n_162),
.Y(n_189)
);

XOR2xp5_ASAP7_75t_SL g160 ( 
.A(n_155),
.B(n_110),
.Y(n_160)
);

XNOR2xp5_ASAP7_75t_L g201 ( 
.A(n_160),
.B(n_164),
.Y(n_201)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_153),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_SL g194 ( 
.A(n_161),
.B(n_167),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_L g162 ( 
.A(n_146),
.B(n_143),
.Y(n_162)
);

OAI32xp33_ASAP7_75t_L g164 ( 
.A1(n_140),
.A2(n_119),
.A3(n_125),
.B1(n_121),
.B2(n_106),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_L g165 ( 
.A(n_140),
.B(n_153),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_L g191 ( 
.A(n_165),
.B(n_166),
.Y(n_191)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_137),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_L g168 ( 
.A(n_144),
.B(n_34),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_L g208 ( 
.A(n_168),
.B(n_172),
.Y(n_208)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_152),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_SL g199 ( 
.A(n_170),
.B(n_178),
.Y(n_199)
);

AOI22xp5_ASAP7_75t_L g171 ( 
.A1(n_151),
.A2(n_107),
.B1(n_128),
.B2(n_109),
.Y(n_171)
);

OAI22xp5_ASAP7_75t_SL g195 ( 
.A1(n_171),
.A2(n_176),
.B1(n_154),
.B2(n_133),
.Y(n_195)
);

MAJIxp5_ASAP7_75t_L g172 ( 
.A(n_135),
.B(n_129),
.C(n_142),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_L g173 ( 
.A(n_145),
.B(n_34),
.Y(n_173)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_173),
.Y(n_204)
);

NOR2xp33_ASAP7_75t_L g209 ( 
.A(n_175),
.B(n_180),
.Y(n_209)
);

AOI22xp5_ASAP7_75t_L g176 ( 
.A1(n_131),
.A2(n_102),
.B1(n_122),
.B2(n_21),
.Y(n_176)
);

XOR2xp5_ASAP7_75t_L g177 ( 
.A(n_129),
.B(n_50),
.Y(n_177)
);

AOI21xp5_ASAP7_75t_L g196 ( 
.A1(n_177),
.A2(n_132),
.B(n_147),
.Y(n_196)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_141),
.Y(n_178)
);

AOI22xp5_ASAP7_75t_L g186 ( 
.A1(n_179),
.A2(n_181),
.B1(n_148),
.B2(n_130),
.Y(n_186)
);

MAJIxp5_ASAP7_75t_L g180 ( 
.A(n_138),
.B(n_98),
.C(n_102),
.Y(n_180)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_149),
.Y(n_182)
);

AOI22xp33_ASAP7_75t_L g192 ( 
.A1(n_182),
.A2(n_130),
.B1(n_133),
.B2(n_149),
.Y(n_192)
);

CKINVDCx20_ASAP7_75t_R g183 ( 
.A(n_136),
.Y(n_183)
);

NOR2xp33_ASAP7_75t_SL g185 ( 
.A(n_183),
.B(n_134),
.Y(n_185)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_185),
.Y(n_212)
);

OAI22xp5_ASAP7_75t_L g223 ( 
.A1(n_186),
.A2(n_192),
.B1(n_203),
.B2(n_206),
.Y(n_223)
);

CKINVDCx20_ASAP7_75t_R g187 ( 
.A(n_158),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_L g232 ( 
.A(n_187),
.B(n_190),
.Y(n_232)
);

INVx3_ASAP7_75t_L g188 ( 
.A(n_171),
.Y(n_188)
);

NOR2xp33_ASAP7_75t_L g226 ( 
.A(n_188),
.B(n_202),
.Y(n_226)
);

INVx1_ASAP7_75t_SL g190 ( 
.A(n_173),
.Y(n_190)
);

INVxp67_ASAP7_75t_L g193 ( 
.A(n_179),
.Y(n_193)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_193),
.Y(n_218)
);

AOI22xp5_ASAP7_75t_L g214 ( 
.A1(n_195),
.A2(n_200),
.B1(n_180),
.B2(n_163),
.Y(n_214)
);

MAJIxp5_ASAP7_75t_L g216 ( 
.A(n_196),
.B(n_166),
.C(n_159),
.Y(n_216)
);

INVxp67_ASAP7_75t_L g197 ( 
.A(n_176),
.Y(n_197)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_197),
.Y(n_219)
);

AOI322xp5_ASAP7_75t_L g198 ( 
.A1(n_160),
.A2(n_139),
.A3(n_156),
.B1(n_17),
.B2(n_31),
.C1(n_9),
.C2(n_12),
.Y(n_198)
);

XNOR2xp5_ASAP7_75t_L g224 ( 
.A(n_198),
.B(n_157),
.Y(n_224)
);

OAI22xp5_ASAP7_75t_L g200 ( 
.A1(n_178),
.A2(n_139),
.B1(n_17),
.B2(n_31),
.Y(n_200)
);

INVx2_ASAP7_75t_L g202 ( 
.A(n_170),
.Y(n_202)
);

AOI22xp5_ASAP7_75t_L g203 ( 
.A1(n_174),
.A2(n_169),
.B1(n_167),
.B2(n_165),
.Y(n_203)
);

CKINVDCx16_ASAP7_75t_R g205 ( 
.A(n_184),
.Y(n_205)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_205),
.Y(n_220)
);

AOI22xp5_ASAP7_75t_L g206 ( 
.A1(n_174),
.A2(n_31),
.B1(n_17),
.B2(n_2),
.Y(n_206)
);

NOR2xp33_ASAP7_75t_SL g207 ( 
.A(n_161),
.B(n_17),
.Y(n_207)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_207),
.Y(n_228)
);

AOI22xp5_ASAP7_75t_L g210 ( 
.A1(n_169),
.A2(n_17),
.B1(n_1),
.B2(n_2),
.Y(n_210)
);

OAI22xp5_ASAP7_75t_L g229 ( 
.A1(n_210),
.A2(n_12),
.B1(n_11),
.B2(n_10),
.Y(n_229)
);

CKINVDCx16_ASAP7_75t_R g211 ( 
.A(n_162),
.Y(n_211)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_211),
.Y(n_233)
);

XNOR2x1_ASAP7_75t_L g213 ( 
.A(n_201),
.B(n_177),
.Y(n_213)
);

XOR2xp5_ASAP7_75t_L g249 ( 
.A(n_213),
.B(n_215),
.Y(n_249)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_214),
.Y(n_242)
);

XOR2xp5_ASAP7_75t_L g215 ( 
.A(n_208),
.B(n_172),
.Y(n_215)
);

XOR2xp5_ASAP7_75t_L g251 ( 
.A(n_216),
.B(n_217),
.Y(n_251)
);

XOR2xp5_ASAP7_75t_L g217 ( 
.A(n_208),
.B(n_175),
.Y(n_217)
);

MAJIxp5_ASAP7_75t_L g221 ( 
.A(n_209),
.B(n_168),
.C(n_182),
.Y(n_221)
);

MAJIxp5_ASAP7_75t_L g238 ( 
.A(n_221),
.B(n_191),
.C(n_204),
.Y(n_238)
);

AOI22xp5_ASAP7_75t_SL g222 ( 
.A1(n_193),
.A2(n_163),
.B1(n_164),
.B2(n_157),
.Y(n_222)
);

INVxp67_ASAP7_75t_L g241 ( 
.A(n_222),
.Y(n_241)
);

NAND2xp5_ASAP7_75t_SL g260 ( 
.A(n_224),
.B(n_225),
.Y(n_260)
);

INVxp67_ASAP7_75t_L g225 ( 
.A(n_207),
.Y(n_225)
);

XOR2xp5_ASAP7_75t_L g227 ( 
.A(n_201),
.B(n_13),
.Y(n_227)
);

XOR2xp5_ASAP7_75t_L g255 ( 
.A(n_227),
.B(n_234),
.Y(n_255)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_229),
.Y(n_243)
);

OAI22xp5_ASAP7_75t_L g230 ( 
.A1(n_203),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_230)
);

CKINVDCx16_ASAP7_75t_R g258 ( 
.A(n_230),
.Y(n_258)
);

AOI22xp5_ASAP7_75t_SL g231 ( 
.A1(n_197),
.A2(n_188),
.B1(n_204),
.B2(n_187),
.Y(n_231)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_231),
.Y(n_245)
);

XOR2xp5_ASAP7_75t_L g234 ( 
.A(n_196),
.B(n_11),
.Y(n_234)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_189),
.Y(n_235)
);

NAND2xp5_ASAP7_75t_L g239 ( 
.A(n_235),
.B(n_236),
.Y(n_239)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_189),
.Y(n_236)
);

A2O1A1Ixp33_ASAP7_75t_SL g237 ( 
.A1(n_210),
.A2(n_1),
.B(n_2),
.C(n_3),
.Y(n_237)
);

AOI21xp5_ASAP7_75t_L g254 ( 
.A1(n_237),
.A2(n_195),
.B(n_3),
.Y(n_254)
);

MAJIxp5_ASAP7_75t_L g263 ( 
.A(n_238),
.B(n_240),
.C(n_246),
.Y(n_263)
);

MAJIxp5_ASAP7_75t_L g240 ( 
.A(n_215),
.B(n_191),
.C(n_186),
.Y(n_240)
);

AND2x2_ASAP7_75t_L g244 ( 
.A(n_234),
.B(n_190),
.Y(n_244)
);

OAI21xp5_ASAP7_75t_SL g275 ( 
.A1(n_244),
.A2(n_254),
.B(n_259),
.Y(n_275)
);

MAJIxp5_ASAP7_75t_L g246 ( 
.A(n_217),
.B(n_194),
.C(n_199),
.Y(n_246)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_232),
.Y(n_247)
);

NAND2xp5_ASAP7_75t_L g267 ( 
.A(n_247),
.B(n_250),
.Y(n_267)
);

XNOR2xp5_ASAP7_75t_L g248 ( 
.A(n_216),
.B(n_213),
.Y(n_248)
);

XNOR2xp5_ASAP7_75t_L g261 ( 
.A(n_248),
.B(n_227),
.Y(n_261)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_226),
.Y(n_250)
);

NAND2xp5_ASAP7_75t_L g252 ( 
.A(n_233),
.B(n_202),
.Y(n_252)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_252),
.Y(n_264)
);

NAND2xp5_ASAP7_75t_L g253 ( 
.A(n_228),
.B(n_206),
.Y(n_253)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_253),
.Y(n_274)
);

NAND2xp5_ASAP7_75t_L g256 ( 
.A(n_225),
.B(n_1),
.Y(n_256)
);

CKINVDCx20_ASAP7_75t_R g276 ( 
.A(n_256),
.Y(n_276)
);

NAND2xp5_ASAP7_75t_L g257 ( 
.A(n_231),
.B(n_3),
.Y(n_257)
);

CKINVDCx20_ASAP7_75t_R g277 ( 
.A(n_257),
.Y(n_277)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_223),
.Y(n_259)
);

XOR2xp5_ASAP7_75t_L g288 ( 
.A(n_261),
.B(n_265),
.Y(n_288)
);

OAI22xp33_ASAP7_75t_R g262 ( 
.A1(n_244),
.A2(n_237),
.B1(n_222),
.B2(n_221),
.Y(n_262)
);

OAI21x1_ASAP7_75t_L g290 ( 
.A1(n_262),
.A2(n_273),
.B(n_243),
.Y(n_290)
);

MAJx2_ASAP7_75t_L g265 ( 
.A(n_249),
.B(n_224),
.C(n_218),
.Y(n_265)
);

A2O1A1O1Ixp25_ASAP7_75t_L g266 ( 
.A1(n_241),
.A2(n_219),
.B(n_212),
.C(n_237),
.D(n_220),
.Y(n_266)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_266),
.Y(n_282)
);

OAI22xp5_ASAP7_75t_SL g268 ( 
.A1(n_241),
.A2(n_242),
.B1(n_245),
.B2(n_240),
.Y(n_268)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_268),
.Y(n_283)
);

AOI22xp5_ASAP7_75t_L g269 ( 
.A1(n_244),
.A2(n_237),
.B1(n_4),
.B2(n_5),
.Y(n_269)
);

OAI22xp5_ASAP7_75t_L g280 ( 
.A1(n_269),
.A2(n_271),
.B1(n_254),
.B2(n_258),
.Y(n_280)
);

MAJIxp5_ASAP7_75t_L g270 ( 
.A(n_251),
.B(n_3),
.C(n_4),
.Y(n_270)
);

MAJIxp5_ASAP7_75t_L g286 ( 
.A(n_270),
.B(n_279),
.C(n_255),
.Y(n_286)
);

AOI22xp5_ASAP7_75t_L g271 ( 
.A1(n_257),
.A2(n_4),
.B1(n_5),
.B2(n_6),
.Y(n_271)
);

CKINVDCx16_ASAP7_75t_R g272 ( 
.A(n_252),
.Y(n_272)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_272),
.Y(n_291)
);

OA21x2_ASAP7_75t_SL g273 ( 
.A1(n_255),
.A2(n_10),
.B(n_11),
.Y(n_273)
);

NOR3xp33_ASAP7_75t_SL g278 ( 
.A(n_260),
.B(n_5),
.C(n_7),
.Y(n_278)
);

AOI21xp33_ASAP7_75t_L g285 ( 
.A1(n_278),
.A2(n_253),
.B(n_256),
.Y(n_285)
);

XNOR2xp5_ASAP7_75t_L g279 ( 
.A(n_248),
.B(n_5),
.Y(n_279)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_280),
.Y(n_299)
);

CKINVDCx16_ASAP7_75t_R g281 ( 
.A(n_267),
.Y(n_281)
);

NAND2xp5_ASAP7_75t_L g298 ( 
.A(n_281),
.B(n_292),
.Y(n_298)
);

HB1xp67_ASAP7_75t_L g284 ( 
.A(n_264),
.Y(n_284)
);

NOR2xp33_ASAP7_75t_L g297 ( 
.A(n_284),
.B(n_286),
.Y(n_297)
);

OAI321xp33_ASAP7_75t_L g309 ( 
.A1(n_285),
.A2(n_290),
.A3(n_7),
.B1(n_261),
.B2(n_279),
.C(n_295),
.Y(n_309)
);

HB1xp67_ASAP7_75t_L g287 ( 
.A(n_274),
.Y(n_287)
);

NOR2xp33_ASAP7_75t_L g304 ( 
.A(n_287),
.B(n_277),
.Y(n_304)
);

MAJIxp5_ASAP7_75t_L g289 ( 
.A(n_263),
.B(n_251),
.C(n_238),
.Y(n_289)
);

MAJIxp5_ASAP7_75t_L g296 ( 
.A(n_289),
.B(n_263),
.C(n_249),
.Y(n_296)
);

CKINVDCx16_ASAP7_75t_R g292 ( 
.A(n_271),
.Y(n_292)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_269),
.Y(n_293)
);

NAND2xp5_ASAP7_75t_L g302 ( 
.A(n_293),
.B(n_295),
.Y(n_302)
);

NAND2xp5_ASAP7_75t_L g294 ( 
.A(n_276),
.B(n_239),
.Y(n_294)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_294),
.Y(n_303)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_266),
.Y(n_295)
);

XOR2xp5_ASAP7_75t_L g310 ( 
.A(n_296),
.B(n_300),
.Y(n_310)
);

XNOR2xp5_ASAP7_75t_L g300 ( 
.A(n_289),
.B(n_268),
.Y(n_300)
);

FAx1_ASAP7_75t_SL g301 ( 
.A(n_294),
.B(n_275),
.CI(n_239),
.CON(n_301),
.SN(n_301)
);

NAND2xp5_ASAP7_75t_L g319 ( 
.A(n_301),
.B(n_306),
.Y(n_319)
);

CKINVDCx16_ASAP7_75t_R g314 ( 
.A(n_304),
.Y(n_314)
);

NOR2xp33_ASAP7_75t_L g305 ( 
.A(n_282),
.B(n_278),
.Y(n_305)
);

CKINVDCx16_ASAP7_75t_R g318 ( 
.A(n_305),
.Y(n_318)
);

NOR2xp33_ASAP7_75t_L g306 ( 
.A(n_283),
.B(n_246),
.Y(n_306)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_291),
.Y(n_307)
);

NOR2xp33_ASAP7_75t_L g312 ( 
.A(n_307),
.B(n_291),
.Y(n_312)
);

OAI22xp5_ASAP7_75t_SL g308 ( 
.A1(n_283),
.A2(n_275),
.B1(n_265),
.B2(n_270),
.Y(n_308)
);

INVxp67_ASAP7_75t_L g320 ( 
.A(n_308),
.Y(n_320)
);

XNOR2xp5_ASAP7_75t_SL g315 ( 
.A(n_309),
.B(n_7),
.Y(n_315)
);

XNOR2xp5_ASAP7_75t_L g311 ( 
.A(n_300),
.B(n_286),
.Y(n_311)
);

NAND2xp5_ASAP7_75t_L g322 ( 
.A(n_311),
.B(n_308),
.Y(n_322)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_312),
.Y(n_324)
);

NOR2xp33_ASAP7_75t_L g313 ( 
.A(n_303),
.B(n_293),
.Y(n_313)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_313),
.Y(n_326)
);

MAJIxp5_ASAP7_75t_L g325 ( 
.A(n_315),
.B(n_302),
.C(n_299),
.Y(n_325)
);

OR2x2_ASAP7_75t_L g316 ( 
.A(n_297),
.B(n_288),
.Y(n_316)
);

AOI21xp5_ASAP7_75t_L g321 ( 
.A1(n_316),
.A2(n_317),
.B(n_319),
.Y(n_321)
);

OAI21xp5_ASAP7_75t_SL g317 ( 
.A1(n_296),
.A2(n_288),
.B(n_7),
.Y(n_317)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_321),
.Y(n_329)
);

MAJIxp5_ASAP7_75t_L g330 ( 
.A(n_322),
.B(n_323),
.C(n_327),
.Y(n_330)
);

NAND2xp5_ASAP7_75t_L g323 ( 
.A(n_314),
.B(n_298),
.Y(n_323)
);

NOR2xp33_ASAP7_75t_SL g331 ( 
.A(n_325),
.B(n_318),
.Y(n_331)
);

XNOR2x1_ASAP7_75t_L g327 ( 
.A(n_320),
.B(n_301),
.Y(n_327)
);

AOI21xp33_ASAP7_75t_L g328 ( 
.A1(n_312),
.A2(n_301),
.B(n_310),
.Y(n_328)
);

NOR2xp33_ASAP7_75t_L g333 ( 
.A(n_328),
.B(n_324),
.Y(n_333)
);

OAI21xp5_ASAP7_75t_L g335 ( 
.A1(n_331),
.A2(n_332),
.B(n_333),
.Y(n_335)
);

XNOR2xp5_ASAP7_75t_L g332 ( 
.A(n_327),
.B(n_313),
.Y(n_332)
);

CKINVDCx14_ASAP7_75t_R g334 ( 
.A(n_333),
.Y(n_334)
);

MAJIxp5_ASAP7_75t_L g336 ( 
.A(n_334),
.B(n_330),
.C(n_329),
.Y(n_336)
);

NAND2xp5_ASAP7_75t_SL g337 ( 
.A(n_336),
.B(n_335),
.Y(n_337)
);

NOR2xp33_ASAP7_75t_SL g338 ( 
.A(n_337),
.B(n_326),
.Y(n_338)
);

BUFx24_ASAP7_75t_SL g339 ( 
.A(n_338),
.Y(n_339)
);


endmodule