module fake_jpeg_1405_n_496 (n_13, n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_496);

input n_13;
input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_496;

wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_15;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_17;
wire n_431;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_490;
wire n_415;
wire n_479;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_48;
wire n_465;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_221;
wire n_256;
wire n_454;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_429;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_474;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_305;
wire n_161;
wire n_441;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_14;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_352;
wire n_350;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_389;
wire n_457;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_296;
wire n_384;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_491;
wire n_24;
wire n_467;
wire n_269;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_473;
wire n_45;
wire n_476;
wire n_337;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_481;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_199;
wire n_260;
wire n_413;
wire n_275;
wire n_494;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_492;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_472;
wire n_279;
wire n_154;
wire n_495;
wire n_205;
wire n_379;
wire n_114;
wire n_444;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_484;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_469;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_482;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_183;
wire n_409;
wire n_249;
wire n_412;
wire n_217;
wire n_471;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_402;
wire n_438;
wire n_475;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

BUFx6f_ASAP7_75t_L g14 ( 
.A(n_8),
.Y(n_14)
);

BUFx6f_ASAP7_75t_L g15 ( 
.A(n_3),
.Y(n_15)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_7),
.Y(n_16)
);

BUFx6f_ASAP7_75t_L g17 ( 
.A(n_13),
.Y(n_17)
);

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_8),
.Y(n_18)
);

INVx8_ASAP7_75t_L g19 ( 
.A(n_10),
.Y(n_19)
);

BUFx12_ASAP7_75t_L g20 ( 
.A(n_2),
.Y(n_20)
);

INVx4_ASAP7_75t_L g21 ( 
.A(n_4),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_8),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_4),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_2),
.Y(n_24)
);

INVx6_ASAP7_75t_L g25 ( 
.A(n_4),
.Y(n_25)
);

INVx2_ASAP7_75t_L g26 ( 
.A(n_0),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_11),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_7),
.Y(n_28)
);

BUFx5_ASAP7_75t_L g29 ( 
.A(n_13),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_10),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_7),
.Y(n_31)
);

INVx2_ASAP7_75t_L g32 ( 
.A(n_9),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_3),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_3),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_9),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_13),
.Y(n_36)
);

INVx5_ASAP7_75t_L g37 ( 
.A(n_13),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_0),
.Y(n_38)
);

INVx6_ASAP7_75t_L g39 ( 
.A(n_4),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_8),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_3),
.Y(n_41)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_10),
.Y(n_42)
);

INVx5_ASAP7_75t_L g43 ( 
.A(n_19),
.Y(n_43)
);

BUFx2_ASAP7_75t_L g130 ( 
.A(n_43),
.Y(n_130)
);

INVx2_ASAP7_75t_L g44 ( 
.A(n_26),
.Y(n_44)
);

INVx2_ASAP7_75t_L g98 ( 
.A(n_44),
.Y(n_98)
);

BUFx3_ASAP7_75t_L g45 ( 
.A(n_37),
.Y(n_45)
);

BUFx3_ASAP7_75t_L g106 ( 
.A(n_45),
.Y(n_106)
);

BUFx8_ASAP7_75t_L g46 ( 
.A(n_29),
.Y(n_46)
);

CKINVDCx14_ASAP7_75t_R g122 ( 
.A(n_46),
.Y(n_122)
);

BUFx2_ASAP7_75t_L g47 ( 
.A(n_19),
.Y(n_47)
);

CKINVDCx16_ASAP7_75t_R g126 ( 
.A(n_47),
.Y(n_126)
);

INVx3_ASAP7_75t_L g48 ( 
.A(n_21),
.Y(n_48)
);

INVx3_ASAP7_75t_L g127 ( 
.A(n_48),
.Y(n_127)
);

INVx2_ASAP7_75t_R g49 ( 
.A(n_21),
.Y(n_49)
);

AND2x2_ASAP7_75t_L g112 ( 
.A(n_49),
.B(n_50),
.Y(n_112)
);

INVx1_ASAP7_75t_SL g50 ( 
.A(n_21),
.Y(n_50)
);

INVx8_ASAP7_75t_L g51 ( 
.A(n_14),
.Y(n_51)
);

INVx5_ASAP7_75t_L g113 ( 
.A(n_51),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_36),
.B(n_12),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_L g108 ( 
.A(n_52),
.B(n_67),
.Y(n_108)
);

BUFx12f_ASAP7_75t_L g53 ( 
.A(n_20),
.Y(n_53)
);

INVx8_ASAP7_75t_L g103 ( 
.A(n_53),
.Y(n_103)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_17),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g99 ( 
.A(n_54),
.Y(n_99)
);

INVx4_ASAP7_75t_L g55 ( 
.A(n_29),
.Y(n_55)
);

INVx3_ASAP7_75t_L g143 ( 
.A(n_55),
.Y(n_143)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_17),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g118 ( 
.A(n_56),
.Y(n_118)
);

INVx3_ASAP7_75t_SL g57 ( 
.A(n_19),
.Y(n_57)
);

INVx2_ASAP7_75t_L g116 ( 
.A(n_57),
.Y(n_116)
);

INVx6_ASAP7_75t_L g58 ( 
.A(n_17),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g152 ( 
.A(n_58),
.Y(n_152)
);

INVx1_ASAP7_75t_SL g59 ( 
.A(n_26),
.Y(n_59)
);

AND2x2_ASAP7_75t_L g132 ( 
.A(n_59),
.B(n_96),
.Y(n_132)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_26),
.Y(n_60)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_60),
.Y(n_114)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_32),
.Y(n_61)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_61),
.Y(n_146)
);

BUFx12f_ASAP7_75t_L g62 ( 
.A(n_20),
.Y(n_62)
);

INVx8_ASAP7_75t_L g129 ( 
.A(n_62),
.Y(n_129)
);

INVx6_ASAP7_75t_L g63 ( 
.A(n_17),
.Y(n_63)
);

BUFx6f_ASAP7_75t_L g155 ( 
.A(n_63),
.Y(n_155)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_14),
.Y(n_64)
);

INVx6_ASAP7_75t_L g128 ( 
.A(n_64),
.Y(n_128)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_14),
.Y(n_65)
);

INVx8_ASAP7_75t_L g134 ( 
.A(n_65),
.Y(n_134)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_32),
.Y(n_66)
);

INVx2_ASAP7_75t_L g119 ( 
.A(n_66),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_L g67 ( 
.A(n_23),
.B(n_12),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_36),
.B(n_12),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_68),
.B(n_80),
.Y(n_97)
);

INVx2_ASAP7_75t_L g69 ( 
.A(n_32),
.Y(n_69)
);

INVx2_ASAP7_75t_L g124 ( 
.A(n_69),
.Y(n_124)
);

INVx4_ASAP7_75t_L g70 ( 
.A(n_29),
.Y(n_70)
);

INVx3_ASAP7_75t_L g145 ( 
.A(n_70),
.Y(n_145)
);

INVx4_ASAP7_75t_L g71 ( 
.A(n_19),
.Y(n_71)
);

INVx3_ASAP7_75t_L g148 ( 
.A(n_71),
.Y(n_148)
);

BUFx5_ASAP7_75t_L g72 ( 
.A(n_20),
.Y(n_72)
);

INVx4_ASAP7_75t_L g104 ( 
.A(n_72),
.Y(n_104)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_25),
.Y(n_73)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_73),
.Y(n_153)
);

BUFx6f_ASAP7_75t_L g74 ( 
.A(n_14),
.Y(n_74)
);

INVx5_ASAP7_75t_L g121 ( 
.A(n_74),
.Y(n_121)
);

INVx11_ASAP7_75t_L g75 ( 
.A(n_20),
.Y(n_75)
);

INVx4_ASAP7_75t_L g107 ( 
.A(n_75),
.Y(n_107)
);

INVx3_ASAP7_75t_L g76 ( 
.A(n_37),
.Y(n_76)
);

INVx3_ASAP7_75t_L g156 ( 
.A(n_76),
.Y(n_156)
);

BUFx3_ASAP7_75t_L g77 ( 
.A(n_37),
.Y(n_77)
);

INVx4_ASAP7_75t_L g131 ( 
.A(n_77),
.Y(n_131)
);

BUFx12_ASAP7_75t_L g78 ( 
.A(n_20),
.Y(n_78)
);

BUFx12_ASAP7_75t_L g111 ( 
.A(n_78),
.Y(n_111)
);

BUFx6f_ASAP7_75t_L g79 ( 
.A(n_15),
.Y(n_79)
);

INVx4_ASAP7_75t_L g136 ( 
.A(n_79),
.Y(n_136)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_25),
.Y(n_80)
);

INVx4_ASAP7_75t_L g81 ( 
.A(n_25),
.Y(n_81)
);

INVx4_ASAP7_75t_L g141 ( 
.A(n_81),
.Y(n_141)
);

CKINVDCx20_ASAP7_75t_R g82 ( 
.A(n_25),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_82),
.B(n_83),
.Y(n_100)
);

OR2x2_ASAP7_75t_L g83 ( 
.A(n_16),
.B(n_12),
.Y(n_83)
);

INVx8_ASAP7_75t_L g84 ( 
.A(n_15),
.Y(n_84)
);

INVx4_ASAP7_75t_L g142 ( 
.A(n_84),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_23),
.B(n_41),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_85),
.B(n_86),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_30),
.B(n_0),
.Y(n_86)
);

CKINVDCx20_ASAP7_75t_R g87 ( 
.A(n_39),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_87),
.B(n_92),
.Y(n_102)
);

INVx3_ASAP7_75t_L g88 ( 
.A(n_39),
.Y(n_88)
);

INVx4_ASAP7_75t_L g149 ( 
.A(n_88),
.Y(n_149)
);

INVx2_ASAP7_75t_L g89 ( 
.A(n_39),
.Y(n_89)
);

INVx2_ASAP7_75t_L g125 ( 
.A(n_89),
.Y(n_125)
);

INVx2_ASAP7_75t_L g90 ( 
.A(n_39),
.Y(n_90)
);

INVx2_ASAP7_75t_L g133 ( 
.A(n_90),
.Y(n_133)
);

INVx2_ASAP7_75t_L g91 ( 
.A(n_15),
.Y(n_91)
);

INVx2_ASAP7_75t_L g135 ( 
.A(n_91),
.Y(n_135)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_15),
.Y(n_92)
);

INVx2_ASAP7_75t_L g93 ( 
.A(n_18),
.Y(n_93)
);

INVx2_ASAP7_75t_L g140 ( 
.A(n_93),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_SL g94 ( 
.A(n_30),
.B(n_0),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_SL g109 ( 
.A(n_94),
.B(n_40),
.Y(n_109)
);

OR2x2_ASAP7_75t_L g95 ( 
.A(n_16),
.B(n_0),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_95),
.B(n_27),
.Y(n_117)
);

INVx4_ASAP7_75t_L g96 ( 
.A(n_18),
.Y(n_96)
);

OAI22xp5_ASAP7_75t_SL g105 ( 
.A1(n_58),
.A2(n_18),
.B1(n_35),
.B2(n_28),
.Y(n_105)
);

AOI22xp5_ASAP7_75t_L g184 ( 
.A1(n_105),
.A2(n_38),
.B1(n_34),
.B2(n_24),
.Y(n_184)
);

NOR2xp33_ASAP7_75t_SL g173 ( 
.A(n_109),
.B(n_110),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_SL g110 ( 
.A(n_83),
.B(n_41),
.Y(n_110)
);

CKINVDCx20_ASAP7_75t_R g115 ( 
.A(n_47),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_L g170 ( 
.A(n_115),
.B(n_117),
.Y(n_170)
);

CKINVDCx20_ASAP7_75t_R g120 ( 
.A(n_64),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_L g171 ( 
.A(n_120),
.B(n_138),
.Y(n_171)
);

OR2x4_ASAP7_75t_L g123 ( 
.A(n_49),
.B(n_95),
.Y(n_123)
);

AND2x4_ASAP7_75t_L g181 ( 
.A(n_123),
.B(n_24),
.Y(n_181)
);

AOI22xp5_ASAP7_75t_L g137 ( 
.A1(n_65),
.A2(n_18),
.B1(n_35),
.B2(n_28),
.Y(n_137)
);

OAI22xp5_ASAP7_75t_L g192 ( 
.A1(n_137),
.A2(n_151),
.B1(n_38),
.B2(n_22),
.Y(n_192)
);

NAND3xp33_ASAP7_75t_SL g138 ( 
.A(n_46),
.B(n_42),
.C(n_16),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_L g139 ( 
.A(n_59),
.B(n_40),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_L g179 ( 
.A(n_139),
.B(n_144),
.Y(n_179)
);

CKINVDCx20_ASAP7_75t_R g144 ( 
.A(n_74),
.Y(n_144)
);

NOR2xp33_ASAP7_75t_L g147 ( 
.A(n_53),
.B(n_27),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_L g186 ( 
.A(n_147),
.B(n_150),
.Y(n_186)
);

CKINVDCx20_ASAP7_75t_R g150 ( 
.A(n_79),
.Y(n_150)
);

AOI22xp33_ASAP7_75t_L g151 ( 
.A1(n_54),
.A2(n_35),
.B1(n_28),
.B2(n_27),
.Y(n_151)
);

NOR2xp33_ASAP7_75t_L g154 ( 
.A(n_53),
.B(n_38),
.Y(n_154)
);

NOR2xp33_ASAP7_75t_L g187 ( 
.A(n_154),
.B(n_62),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_SL g157 ( 
.A(n_108),
.B(n_100),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_SL g220 ( 
.A(n_157),
.B(n_124),
.Y(n_220)
);

AOI22xp33_ASAP7_75t_SL g158 ( 
.A1(n_123),
.A2(n_46),
.B1(n_71),
.B2(n_70),
.Y(n_158)
);

AOI22xp33_ASAP7_75t_SL g218 ( 
.A1(n_158),
.A2(n_168),
.B1(n_175),
.B2(n_189),
.Y(n_218)
);

INVx2_ASAP7_75t_L g159 ( 
.A(n_125),
.Y(n_159)
);

BUFx2_ASAP7_75t_L g210 ( 
.A(n_159),
.Y(n_210)
);

OAI22xp33_ASAP7_75t_SL g160 ( 
.A1(n_151),
.A2(n_55),
.B1(n_96),
.B2(n_77),
.Y(n_160)
);

AOI22xp33_ASAP7_75t_L g226 ( 
.A1(n_160),
.A2(n_75),
.B1(n_145),
.B2(n_143),
.Y(n_226)
);

INVx11_ASAP7_75t_L g161 ( 
.A(n_122),
.Y(n_161)
);

INVx4_ASAP7_75t_L g224 ( 
.A(n_161),
.Y(n_224)
);

INVx2_ASAP7_75t_L g162 ( 
.A(n_133),
.Y(n_162)
);

INVx2_ASAP7_75t_L g203 ( 
.A(n_162),
.Y(n_203)
);

BUFx10_ASAP7_75t_L g163 ( 
.A(n_111),
.Y(n_163)
);

INVx8_ASAP7_75t_L g227 ( 
.A(n_163),
.Y(n_227)
);

INVx3_ASAP7_75t_L g164 ( 
.A(n_116),
.Y(n_164)
);

INVx3_ASAP7_75t_L g208 ( 
.A(n_164),
.Y(n_208)
);

CKINVDCx12_ASAP7_75t_R g165 ( 
.A(n_112),
.Y(n_165)
);

INVx1_ASAP7_75t_SL g213 ( 
.A(n_165),
.Y(n_213)
);

INVx3_ASAP7_75t_L g166 ( 
.A(n_142),
.Y(n_166)
);

INVx3_ASAP7_75t_L g216 ( 
.A(n_166),
.Y(n_216)
);

BUFx6f_ASAP7_75t_L g167 ( 
.A(n_99),
.Y(n_167)
);

INVx3_ASAP7_75t_L g230 ( 
.A(n_167),
.Y(n_230)
);

AOI22xp33_ASAP7_75t_SL g168 ( 
.A1(n_112),
.A2(n_45),
.B1(n_31),
.B2(n_42),
.Y(n_168)
);

INVx5_ASAP7_75t_L g169 ( 
.A(n_103),
.Y(n_169)
);

HB1xp67_ASAP7_75t_L g222 ( 
.A(n_169),
.Y(n_222)
);

INVx2_ASAP7_75t_L g172 ( 
.A(n_135),
.Y(n_172)
);

INVx2_ASAP7_75t_L g207 ( 
.A(n_172),
.Y(n_207)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_114),
.Y(n_174)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_174),
.Y(n_201)
);

AOI22xp33_ASAP7_75t_SL g175 ( 
.A1(n_105),
.A2(n_31),
.B1(n_42),
.B2(n_22),
.Y(n_175)
);

INVx1_ASAP7_75t_SL g176 ( 
.A(n_132),
.Y(n_176)
);

AND2x2_ASAP7_75t_L g202 ( 
.A(n_176),
.B(n_177),
.Y(n_202)
);

OA22x2_ASAP7_75t_L g177 ( 
.A1(n_137),
.A2(n_81),
.B1(n_63),
.B2(n_56),
.Y(n_177)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_146),
.Y(n_178)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_178),
.Y(n_204)
);

INVx3_ASAP7_75t_L g180 ( 
.A(n_142),
.Y(n_180)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_180),
.Y(n_206)
);

AND2x2_ASAP7_75t_L g225 ( 
.A(n_181),
.B(n_183),
.Y(n_225)
);

INVx2_ASAP7_75t_L g182 ( 
.A(n_140),
.Y(n_182)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_182),
.Y(n_212)
);

INVx13_ASAP7_75t_L g183 ( 
.A(n_111),
.Y(n_183)
);

AOI22xp5_ASAP7_75t_L g211 ( 
.A1(n_184),
.A2(n_192),
.B1(n_31),
.B2(n_34),
.Y(n_211)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_153),
.Y(n_185)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_185),
.Y(n_217)
);

NOR2xp33_ASAP7_75t_L g214 ( 
.A(n_187),
.B(n_190),
.Y(n_214)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_132),
.Y(n_188)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_188),
.Y(n_219)
);

BUFx12f_ASAP7_75t_L g189 ( 
.A(n_103),
.Y(n_189)
);

NOR2xp33_ASAP7_75t_L g190 ( 
.A(n_101),
.B(n_62),
.Y(n_190)
);

AOI22xp5_ASAP7_75t_SL g191 ( 
.A1(n_97),
.A2(n_102),
.B1(n_57),
.B2(n_143),
.Y(n_191)
);

OR2x2_ASAP7_75t_L g209 ( 
.A(n_191),
.B(n_198),
.Y(n_209)
);

INVx3_ASAP7_75t_L g193 ( 
.A(n_113),
.Y(n_193)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_193),
.Y(n_231)
);

NOR2xp33_ASAP7_75t_L g194 ( 
.A(n_98),
.B(n_51),
.Y(n_194)
);

NOR2xp33_ASAP7_75t_L g229 ( 
.A(n_194),
.B(n_197),
.Y(n_229)
);

OAI22xp5_ASAP7_75t_L g195 ( 
.A1(n_128),
.A2(n_84),
.B1(n_28),
.B2(n_35),
.Y(n_195)
);

OAI22xp5_ASAP7_75t_L g215 ( 
.A1(n_195),
.A2(n_128),
.B1(n_118),
.B2(n_136),
.Y(n_215)
);

INVx3_ASAP7_75t_L g196 ( 
.A(n_113),
.Y(n_196)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_196),
.Y(n_233)
);

INVx2_ASAP7_75t_L g197 ( 
.A(n_141),
.Y(n_197)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_141),
.Y(n_198)
);

INVx13_ASAP7_75t_L g199 ( 
.A(n_111),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_L g205 ( 
.A(n_199),
.B(n_200),
.Y(n_205)
);

INVx6_ASAP7_75t_L g200 ( 
.A(n_99),
.Y(n_200)
);

AOI22xp5_ASAP7_75t_L g238 ( 
.A1(n_211),
.A2(n_215),
.B1(n_221),
.B2(n_223),
.Y(n_238)
);

NAND2xp5_ASAP7_75t_SL g240 ( 
.A(n_220),
.B(n_231),
.Y(n_240)
);

OAI22xp5_ASAP7_75t_L g221 ( 
.A1(n_192),
.A2(n_155),
.B1(n_152),
.B2(n_136),
.Y(n_221)
);

AOI22xp5_ASAP7_75t_L g223 ( 
.A1(n_181),
.A2(n_119),
.B1(n_155),
.B2(n_152),
.Y(n_223)
);

AOI22xp33_ASAP7_75t_SL g254 ( 
.A1(n_226),
.A2(n_228),
.B1(n_161),
.B2(n_186),
.Y(n_254)
);

AOI22xp33_ASAP7_75t_L g228 ( 
.A1(n_171),
.A2(n_127),
.B1(n_156),
.B2(n_121),
.Y(n_228)
);

NAND2xp5_ASAP7_75t_SL g232 ( 
.A(n_157),
.B(n_149),
.Y(n_232)
);

NAND2xp5_ASAP7_75t_L g256 ( 
.A(n_232),
.B(n_234),
.Y(n_256)
);

OAI21xp5_ASAP7_75t_L g234 ( 
.A1(n_181),
.A2(n_145),
.B(n_34),
.Y(n_234)
);

AND2x2_ASAP7_75t_L g242 ( 
.A(n_234),
.B(n_188),
.Y(n_242)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_201),
.Y(n_235)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_235),
.Y(n_262)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_201),
.Y(n_236)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_236),
.Y(n_284)
);

CKINVDCx20_ASAP7_75t_R g237 ( 
.A(n_210),
.Y(n_237)
);

NOR2xp33_ASAP7_75t_L g278 ( 
.A(n_237),
.B(n_253),
.Y(n_278)
);

AOI22xp5_ASAP7_75t_SL g239 ( 
.A1(n_202),
.A2(n_181),
.B1(n_165),
.B2(n_176),
.Y(n_239)
);

OAI21xp5_ASAP7_75t_SL g283 ( 
.A1(n_239),
.A2(n_242),
.B(n_206),
.Y(n_283)
);

NAND2xp5_ASAP7_75t_SL g273 ( 
.A(n_240),
.B(n_247),
.Y(n_273)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_204),
.Y(n_241)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_241),
.Y(n_287)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_204),
.Y(n_243)
);

INVxp67_ASAP7_75t_L g268 ( 
.A(n_243),
.Y(n_268)
);

CKINVDCx14_ASAP7_75t_R g244 ( 
.A(n_225),
.Y(n_244)
);

NAND2xp5_ASAP7_75t_SL g267 ( 
.A(n_244),
.B(n_258),
.Y(n_267)
);

MAJx2_ASAP7_75t_L g245 ( 
.A(n_232),
.B(n_191),
.C(n_178),
.Y(n_245)
);

FAx1_ASAP7_75t_SL g275 ( 
.A(n_245),
.B(n_213),
.CI(n_222),
.CON(n_275),
.SN(n_275)
);

BUFx6f_ASAP7_75t_L g246 ( 
.A(n_230),
.Y(n_246)
);

INVx4_ASAP7_75t_L g269 ( 
.A(n_246),
.Y(n_269)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_217),
.Y(n_247)
);

AOI22xp5_ASAP7_75t_L g248 ( 
.A1(n_202),
.A2(n_195),
.B1(n_184),
.B2(n_177),
.Y(n_248)
);

OAI22xp5_ASAP7_75t_L g280 ( 
.A1(n_248),
.A2(n_215),
.B1(n_205),
.B2(n_233),
.Y(n_280)
);

INVx3_ASAP7_75t_L g249 ( 
.A(n_230),
.Y(n_249)
);

INVx4_ASAP7_75t_L g274 ( 
.A(n_249),
.Y(n_274)
);

BUFx2_ASAP7_75t_L g250 ( 
.A(n_216),
.Y(n_250)
);

AOI22xp33_ASAP7_75t_SL g276 ( 
.A1(n_250),
.A2(n_254),
.B1(n_255),
.B2(n_257),
.Y(n_276)
);

NOR2xp33_ASAP7_75t_L g251 ( 
.A(n_214),
.B(n_170),
.Y(n_251)
);

CKINVDCx14_ASAP7_75t_R g270 ( 
.A(n_251),
.Y(n_270)
);

HB1xp67_ASAP7_75t_L g252 ( 
.A(n_208),
.Y(n_252)
);

CKINVDCx20_ASAP7_75t_R g265 ( 
.A(n_252),
.Y(n_265)
);

CKINVDCx20_ASAP7_75t_R g253 ( 
.A(n_210),
.Y(n_253)
);

BUFx6f_ASAP7_75t_L g255 ( 
.A(n_231),
.Y(n_255)
);

NAND2xp5_ASAP7_75t_L g263 ( 
.A(n_256),
.B(n_259),
.Y(n_263)
);

INVx2_ASAP7_75t_L g257 ( 
.A(n_217),
.Y(n_257)
);

NOR2xp33_ASAP7_75t_L g258 ( 
.A(n_220),
.B(n_179),
.Y(n_258)
);

CKINVDCx16_ASAP7_75t_R g259 ( 
.A(n_225),
.Y(n_259)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_212),
.Y(n_260)
);

NAND2xp5_ASAP7_75t_L g281 ( 
.A(n_260),
.B(n_261),
.Y(n_281)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_212),
.Y(n_261)
);

OAI221xp5_ASAP7_75t_L g264 ( 
.A1(n_256),
.A2(n_219),
.B1(n_218),
.B2(n_229),
.C(n_225),
.Y(n_264)
);

NAND2xp5_ASAP7_75t_SL g312 ( 
.A(n_264),
.B(n_224),
.Y(n_312)
);

AOI22xp5_ASAP7_75t_L g266 ( 
.A1(n_248),
.A2(n_202),
.B1(n_209),
.B2(n_221),
.Y(n_266)
);

OAI22xp5_ASAP7_75t_SL g293 ( 
.A1(n_266),
.A2(n_240),
.B1(n_235),
.B2(n_236),
.Y(n_293)
);

OAI22xp5_ASAP7_75t_SL g271 ( 
.A1(n_238),
.A2(n_209),
.B1(n_211),
.B2(n_223),
.Y(n_271)
);

AOI22xp5_ASAP7_75t_L g291 ( 
.A1(n_271),
.A2(n_272),
.B1(n_280),
.B2(n_282),
.Y(n_291)
);

OAI22xp5_ASAP7_75t_SL g272 ( 
.A1(n_238),
.A2(n_209),
.B1(n_219),
.B2(n_205),
.Y(n_272)
);

OR2x2_ASAP7_75t_L g305 ( 
.A(n_275),
.B(n_288),
.Y(n_305)
);

XNOR2xp5_ASAP7_75t_L g277 ( 
.A(n_239),
.B(n_213),
.Y(n_277)
);

XOR2xp5_ASAP7_75t_L g289 ( 
.A(n_277),
.B(n_279),
.Y(n_289)
);

XNOR2xp5_ASAP7_75t_L g279 ( 
.A(n_245),
.B(n_174),
.Y(n_279)
);

OAI22xp5_ASAP7_75t_SL g282 ( 
.A1(n_242),
.A2(n_177),
.B1(n_200),
.B2(n_233),
.Y(n_282)
);

CKINVDCx14_ASAP7_75t_R g304 ( 
.A(n_283),
.Y(n_304)
);

XNOR2xp5_ASAP7_75t_L g285 ( 
.A(n_245),
.B(n_185),
.Y(n_285)
);

XOR2xp5_ASAP7_75t_L g295 ( 
.A(n_285),
.B(n_286),
.Y(n_295)
);

XNOR2xp5_ASAP7_75t_L g286 ( 
.A(n_242),
.B(n_173),
.Y(n_286)
);

AOI21xp5_ASAP7_75t_L g288 ( 
.A1(n_259),
.A2(n_224),
.B(n_216),
.Y(n_288)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_281),
.Y(n_290)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_290),
.Y(n_319)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_281),
.Y(n_292)
);

INVx1_ASAP7_75t_L g342 ( 
.A(n_292),
.Y(n_342)
);

AOI22xp5_ASAP7_75t_L g333 ( 
.A1(n_293),
.A2(n_282),
.B1(n_264),
.B2(n_275),
.Y(n_333)
);

CKINVDCx12_ASAP7_75t_R g294 ( 
.A(n_265),
.Y(n_294)
);

BUFx5_ASAP7_75t_L g330 ( 
.A(n_294),
.Y(n_330)
);

INVx13_ASAP7_75t_L g296 ( 
.A(n_288),
.Y(n_296)
);

CKINVDCx14_ASAP7_75t_R g321 ( 
.A(n_296),
.Y(n_321)
);

INVx13_ASAP7_75t_L g297 ( 
.A(n_265),
.Y(n_297)
);

CKINVDCx14_ASAP7_75t_R g336 ( 
.A(n_297),
.Y(n_336)
);

NAND2xp5_ASAP7_75t_L g298 ( 
.A(n_273),
.B(n_257),
.Y(n_298)
);

NAND2xp5_ASAP7_75t_L g318 ( 
.A(n_298),
.B(n_309),
.Y(n_318)
);

CKINVDCx20_ASAP7_75t_R g299 ( 
.A(n_268),
.Y(n_299)
);

NOR2xp33_ASAP7_75t_L g320 ( 
.A(n_299),
.B(n_303),
.Y(n_320)
);

XNOR2xp5_ASAP7_75t_L g300 ( 
.A(n_279),
.B(n_241),
.Y(n_300)
);

XOR2xp5_ASAP7_75t_L g328 ( 
.A(n_300),
.B(n_286),
.Y(n_328)
);

AOI22xp5_ASAP7_75t_L g301 ( 
.A1(n_271),
.A2(n_243),
.B1(n_247),
.B2(n_237),
.Y(n_301)
);

OAI22xp5_ASAP7_75t_SL g324 ( 
.A1(n_301),
.A2(n_287),
.B1(n_284),
.B2(n_263),
.Y(n_324)
);

XOR2xp5_ASAP7_75t_L g302 ( 
.A(n_285),
.B(n_261),
.Y(n_302)
);

MAJIxp5_ASAP7_75t_L g325 ( 
.A(n_302),
.B(n_277),
.C(n_283),
.Y(n_325)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_262),
.Y(n_303)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_262),
.Y(n_306)
);

NOR2xp33_ASAP7_75t_L g331 ( 
.A(n_306),
.B(n_310),
.Y(n_331)
);

OAI22xp5_ASAP7_75t_L g307 ( 
.A1(n_266),
.A2(n_253),
.B1(n_260),
.B2(n_249),
.Y(n_307)
);

AOI22xp33_ASAP7_75t_L g340 ( 
.A1(n_307),
.A2(n_308),
.B1(n_314),
.B2(n_210),
.Y(n_340)
);

OAI22xp5_ASAP7_75t_L g308 ( 
.A1(n_280),
.A2(n_246),
.B1(n_255),
.B2(n_250),
.Y(n_308)
);

AND2x6_ASAP7_75t_L g309 ( 
.A(n_275),
.B(n_183),
.Y(n_309)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_284),
.Y(n_310)
);

NOR2xp33_ASAP7_75t_L g311 ( 
.A(n_270),
.B(n_173),
.Y(n_311)
);

NOR2xp33_ASAP7_75t_SL g327 ( 
.A(n_311),
.B(n_267),
.Y(n_327)
);

OAI21xp5_ASAP7_75t_L g343 ( 
.A1(n_312),
.A2(n_305),
.B(n_304),
.Y(n_343)
);

CKINVDCx20_ASAP7_75t_R g313 ( 
.A(n_268),
.Y(n_313)
);

NOR2xp33_ASAP7_75t_L g332 ( 
.A(n_313),
.B(n_287),
.Y(n_332)
);

OAI22xp5_ASAP7_75t_L g314 ( 
.A1(n_263),
.A2(n_246),
.B1(n_255),
.B2(n_250),
.Y(n_314)
);

NAND2xp5_ASAP7_75t_L g315 ( 
.A(n_273),
.B(n_206),
.Y(n_315)
);

NAND2xp5_ASAP7_75t_L g322 ( 
.A(n_315),
.B(n_278),
.Y(n_322)
);

INVx13_ASAP7_75t_L g316 ( 
.A(n_274),
.Y(n_316)
);

INVx3_ASAP7_75t_L g344 ( 
.A(n_316),
.Y(n_344)
);

INVxp67_ASAP7_75t_L g317 ( 
.A(n_293),
.Y(n_317)
);

NOR2xp33_ASAP7_75t_L g347 ( 
.A(n_317),
.B(n_323),
.Y(n_347)
);

INVx1_ASAP7_75t_L g355 ( 
.A(n_322),
.Y(n_355)
);

CKINVDCx20_ASAP7_75t_R g323 ( 
.A(n_314),
.Y(n_323)
);

AOI22xp5_ASAP7_75t_L g366 ( 
.A1(n_324),
.A2(n_316),
.B1(n_162),
.B2(n_159),
.Y(n_366)
);

XNOR2xp5_ASAP7_75t_L g350 ( 
.A(n_325),
.B(n_328),
.Y(n_350)
);

NAND2xp5_ASAP7_75t_L g326 ( 
.A(n_299),
.B(n_272),
.Y(n_326)
);

INVx1_ASAP7_75t_L g361 ( 
.A(n_326),
.Y(n_361)
);

NAND2xp5_ASAP7_75t_SL g346 ( 
.A(n_327),
.B(n_300),
.Y(n_346)
);

CKINVDCx20_ASAP7_75t_R g329 ( 
.A(n_298),
.Y(n_329)
);

NOR2xp33_ASAP7_75t_L g353 ( 
.A(n_329),
.B(n_337),
.Y(n_353)
);

INVx1_ASAP7_75t_L g367 ( 
.A(n_332),
.Y(n_367)
);

OAI22xp5_ASAP7_75t_SL g348 ( 
.A1(n_333),
.A2(n_305),
.B1(n_291),
.B2(n_326),
.Y(n_348)
);

AND2x2_ASAP7_75t_L g334 ( 
.A(n_307),
.B(n_274),
.Y(n_334)
);

INVx1_ASAP7_75t_SL g369 ( 
.A(n_334),
.Y(n_369)
);

NAND2xp5_ASAP7_75t_L g335 ( 
.A(n_313),
.B(n_269),
.Y(n_335)
);

INVx1_ASAP7_75t_L g371 ( 
.A(n_335),
.Y(n_371)
);

CKINVDCx20_ASAP7_75t_R g337 ( 
.A(n_315),
.Y(n_337)
);

NOR4xp25_ASAP7_75t_L g338 ( 
.A(n_290),
.B(n_276),
.C(n_207),
.D(n_203),
.Y(n_338)
);

AOI21xp33_ASAP7_75t_L g358 ( 
.A1(n_338),
.A2(n_339),
.B(n_341),
.Y(n_358)
);

NOR2xp33_ASAP7_75t_L g339 ( 
.A(n_292),
.B(n_269),
.Y(n_339)
);

OAI22xp5_ASAP7_75t_L g345 ( 
.A1(n_340),
.A2(n_308),
.B1(n_291),
.B2(n_301),
.Y(n_345)
);

NOR2xp33_ASAP7_75t_L g341 ( 
.A(n_303),
.B(n_208),
.Y(n_341)
);

OAI21xp5_ASAP7_75t_SL g349 ( 
.A1(n_343),
.A2(n_305),
.B(n_309),
.Y(n_349)
);

OAI22xp5_ASAP7_75t_L g375 ( 
.A1(n_345),
.A2(n_357),
.B1(n_363),
.B2(n_366),
.Y(n_375)
);

NAND2xp5_ASAP7_75t_L g383 ( 
.A(n_346),
.B(n_349),
.Y(n_383)
);

AOI22xp5_ASAP7_75t_SL g381 ( 
.A1(n_348),
.A2(n_321),
.B1(n_334),
.B2(n_338),
.Y(n_381)
);

XOR2x2_ASAP7_75t_SL g351 ( 
.A(n_324),
.B(n_289),
.Y(n_351)
);

XNOR2xp5_ASAP7_75t_L g372 ( 
.A(n_351),
.B(n_322),
.Y(n_372)
);

AOI21xp5_ASAP7_75t_L g352 ( 
.A1(n_343),
.A2(n_296),
.B(n_294),
.Y(n_352)
);

HB1xp67_ASAP7_75t_L g396 ( 
.A(n_352),
.Y(n_396)
);

MAJIxp5_ASAP7_75t_L g354 ( 
.A(n_325),
.B(n_302),
.C(n_295),
.Y(n_354)
);

MAJIxp5_ASAP7_75t_L g373 ( 
.A(n_354),
.B(n_360),
.C(n_362),
.Y(n_373)
);

NAND2xp5_ASAP7_75t_SL g356 ( 
.A(n_327),
.B(n_295),
.Y(n_356)
);

NAND2xp5_ASAP7_75t_L g384 ( 
.A(n_356),
.B(n_364),
.Y(n_384)
);

OAI22xp5_ASAP7_75t_L g357 ( 
.A1(n_337),
.A2(n_296),
.B1(n_289),
.B2(n_306),
.Y(n_357)
);

MAJx2_ASAP7_75t_L g359 ( 
.A(n_328),
.B(n_310),
.C(n_297),
.Y(n_359)
);

XNOR2xp5_ASAP7_75t_SL g388 ( 
.A(n_359),
.B(n_331),
.Y(n_388)
);

MAJIxp5_ASAP7_75t_L g360 ( 
.A(n_319),
.B(n_297),
.C(n_196),
.Y(n_360)
);

MAJIxp5_ASAP7_75t_L g362 ( 
.A(n_319),
.B(n_342),
.C(n_332),
.Y(n_362)
);

OAI22xp5_ASAP7_75t_L g363 ( 
.A1(n_342),
.A2(n_316),
.B1(n_227),
.B2(n_177),
.Y(n_363)
);

NAND2xp5_ASAP7_75t_SL g364 ( 
.A(n_318),
.B(n_203),
.Y(n_364)
);

NOR2xp33_ASAP7_75t_L g365 ( 
.A(n_318),
.B(n_207),
.Y(n_365)
);

NAND2xp5_ASAP7_75t_L g391 ( 
.A(n_365),
.B(n_344),
.Y(n_391)
);

XOR2xp5_ASAP7_75t_L g368 ( 
.A(n_333),
.B(n_199),
.Y(n_368)
);

XOR2xp5_ASAP7_75t_L g393 ( 
.A(n_368),
.B(n_198),
.Y(n_393)
);

AOI22xp5_ASAP7_75t_L g370 ( 
.A1(n_323),
.A2(n_227),
.B1(n_167),
.B2(n_193),
.Y(n_370)
);

OAI22xp5_ASAP7_75t_SL g374 ( 
.A1(n_370),
.A2(n_340),
.B1(n_336),
.B2(n_334),
.Y(n_374)
);

XNOR2xp5_ASAP7_75t_L g406 ( 
.A(n_372),
.B(n_376),
.Y(n_406)
);

INVx1_ASAP7_75t_L g417 ( 
.A(n_374),
.Y(n_417)
);

XNOR2xp5_ASAP7_75t_L g376 ( 
.A(n_351),
.B(n_320),
.Y(n_376)
);

NAND2xp5_ASAP7_75t_SL g377 ( 
.A(n_349),
.B(n_320),
.Y(n_377)
);

NAND3xp33_ASAP7_75t_L g403 ( 
.A(n_377),
.B(n_392),
.C(n_394),
.Y(n_403)
);

INVx1_ASAP7_75t_L g378 ( 
.A(n_353),
.Y(n_378)
);

INVx1_ASAP7_75t_L g402 ( 
.A(n_378),
.Y(n_402)
);

AOI22xp5_ASAP7_75t_L g379 ( 
.A1(n_345),
.A2(n_361),
.B1(n_348),
.B2(n_347),
.Y(n_379)
);

OAI22xp5_ASAP7_75t_L g398 ( 
.A1(n_379),
.A2(n_380),
.B1(n_381),
.B2(n_385),
.Y(n_398)
);

AOI22xp5_ASAP7_75t_L g380 ( 
.A1(n_361),
.A2(n_329),
.B1(n_334),
.B2(n_321),
.Y(n_380)
);

XNOR2xp5_ASAP7_75t_L g382 ( 
.A(n_350),
.B(n_339),
.Y(n_382)
);

XNOR2xp5_ASAP7_75t_L g409 ( 
.A(n_382),
.B(n_395),
.Y(n_409)
);

AOI22xp5_ASAP7_75t_L g385 ( 
.A1(n_367),
.A2(n_336),
.B1(n_335),
.B2(n_331),
.Y(n_385)
);

INVx1_ASAP7_75t_L g386 ( 
.A(n_362),
.Y(n_386)
);

INVx1_ASAP7_75t_L g414 ( 
.A(n_386),
.Y(n_414)
);

INVx1_ASAP7_75t_L g387 ( 
.A(n_367),
.Y(n_387)
);

HB1xp67_ASAP7_75t_L g404 ( 
.A(n_387),
.Y(n_404)
);

XOR2xp5_ASAP7_75t_L g401 ( 
.A(n_388),
.B(n_393),
.Y(n_401)
);

AOI22xp5_ASAP7_75t_SL g389 ( 
.A1(n_357),
.A2(n_344),
.B1(n_341),
.B2(n_330),
.Y(n_389)
);

OAI22xp5_ASAP7_75t_L g408 ( 
.A1(n_389),
.A2(n_368),
.B1(n_370),
.B2(n_358),
.Y(n_408)
);

MAJIxp5_ASAP7_75t_L g390 ( 
.A(n_354),
.B(n_330),
.C(n_344),
.Y(n_390)
);

MAJIxp5_ASAP7_75t_L g399 ( 
.A(n_390),
.B(n_359),
.C(n_360),
.Y(n_399)
);

NAND2xp5_ASAP7_75t_L g405 ( 
.A(n_391),
.B(n_366),
.Y(n_405)
);

NOR2xp33_ASAP7_75t_L g392 ( 
.A(n_355),
.B(n_227),
.Y(n_392)
);

CKINVDCx20_ASAP7_75t_R g394 ( 
.A(n_352),
.Y(n_394)
);

XOR2xp5_ASAP7_75t_L g395 ( 
.A(n_350),
.B(n_163),
.Y(n_395)
);

INVx1_ASAP7_75t_L g397 ( 
.A(n_355),
.Y(n_397)
);

HB1xp67_ASAP7_75t_L g413 ( 
.A(n_397),
.Y(n_413)
);

NAND2xp5_ASAP7_75t_SL g421 ( 
.A(n_399),
.B(n_400),
.Y(n_421)
);

MAJIxp5_ASAP7_75t_L g400 ( 
.A(n_373),
.B(n_369),
.C(n_371),
.Y(n_400)
);

INVx1_ASAP7_75t_L g422 ( 
.A(n_405),
.Y(n_422)
);

MAJIxp5_ASAP7_75t_L g407 ( 
.A(n_373),
.B(n_369),
.C(n_371),
.Y(n_407)
);

NAND2xp5_ASAP7_75t_SL g435 ( 
.A(n_407),
.B(n_416),
.Y(n_435)
);

AOI22xp5_ASAP7_75t_L g428 ( 
.A1(n_408),
.A2(n_411),
.B1(n_381),
.B2(n_134),
.Y(n_428)
);

NOR2xp33_ASAP7_75t_L g410 ( 
.A(n_382),
.B(n_363),
.Y(n_410)
);

NOR2xp67_ASAP7_75t_L g426 ( 
.A(n_410),
.B(n_418),
.Y(n_426)
);

AOI22xp5_ASAP7_75t_L g411 ( 
.A1(n_375),
.A2(n_167),
.B1(n_180),
.B2(n_166),
.Y(n_411)
);

INVxp67_ASAP7_75t_SL g412 ( 
.A(n_390),
.Y(n_412)
);

INVx1_ASAP7_75t_L g427 ( 
.A(n_412),
.Y(n_427)
);

NAND2xp5_ASAP7_75t_L g415 ( 
.A(n_385),
.B(n_182),
.Y(n_415)
);

AOI21xp5_ASAP7_75t_L g424 ( 
.A1(n_415),
.A2(n_393),
.B(n_395),
.Y(n_424)
);

CKINVDCx20_ASAP7_75t_R g416 ( 
.A(n_396),
.Y(n_416)
);

NOR2xp33_ASAP7_75t_L g418 ( 
.A(n_384),
.B(n_164),
.Y(n_418)
);

CKINVDCx20_ASAP7_75t_R g419 ( 
.A(n_380),
.Y(n_419)
);

NOR2xp33_ASAP7_75t_L g429 ( 
.A(n_419),
.B(n_169),
.Y(n_429)
);

MAJx2_ASAP7_75t_L g420 ( 
.A(n_406),
.B(n_376),
.C(n_372),
.Y(n_420)
);

XNOR2xp5_ASAP7_75t_L g446 ( 
.A(n_420),
.B(n_401),
.Y(n_446)
);

OAI21xp33_ASAP7_75t_L g423 ( 
.A1(n_398),
.A2(n_383),
.B(n_379),
.Y(n_423)
);

OAI21xp5_ASAP7_75t_L g439 ( 
.A1(n_423),
.A2(n_436),
.B(n_404),
.Y(n_439)
);

INVx1_ASAP7_75t_L g441 ( 
.A(n_424),
.Y(n_441)
);

AOI21xp5_ASAP7_75t_L g425 ( 
.A1(n_403),
.A2(n_389),
.B(n_388),
.Y(n_425)
);

AOI21xp5_ASAP7_75t_L g442 ( 
.A1(n_425),
.A2(n_433),
.B(n_402),
.Y(n_442)
);

AOI22xp5_ASAP7_75t_L g440 ( 
.A1(n_428),
.A2(n_417),
.B1(n_413),
.B2(n_411),
.Y(n_440)
);

INVx1_ASAP7_75t_L g444 ( 
.A(n_429),
.Y(n_444)
);

MAJIxp5_ASAP7_75t_L g430 ( 
.A(n_400),
.B(n_148),
.C(n_197),
.Y(n_430)
);

NAND2xp5_ASAP7_75t_L g443 ( 
.A(n_430),
.B(n_431),
.Y(n_443)
);

MAJIxp5_ASAP7_75t_L g431 ( 
.A(n_407),
.B(n_148),
.C(n_163),
.Y(n_431)
);

MAJIxp5_ASAP7_75t_L g432 ( 
.A(n_399),
.B(n_163),
.C(n_130),
.Y(n_432)
);

NAND2xp5_ASAP7_75t_L g450 ( 
.A(n_432),
.B(n_434),
.Y(n_450)
);

AOI21xp5_ASAP7_75t_L g433 ( 
.A1(n_414),
.A2(n_104),
.B(n_156),
.Y(n_433)
);

XNOR2xp5_ASAP7_75t_L g434 ( 
.A(n_406),
.B(n_130),
.Y(n_434)
);

AOI21xp5_ASAP7_75t_SL g436 ( 
.A1(n_417),
.A2(n_172),
.B(n_33),
.Y(n_436)
);

XOR2xp5_ASAP7_75t_L g437 ( 
.A(n_409),
.B(n_189),
.Y(n_437)
);

AND2x2_ASAP7_75t_L g454 ( 
.A(n_437),
.B(n_129),
.Y(n_454)
);

MAJIxp5_ASAP7_75t_L g438 ( 
.A(n_409),
.B(n_126),
.C(n_149),
.Y(n_438)
);

MAJIxp5_ASAP7_75t_L g447 ( 
.A(n_438),
.B(n_104),
.C(n_131),
.Y(n_447)
);

INVx1_ASAP7_75t_L g462 ( 
.A(n_439),
.Y(n_462)
);

AOI22xp5_ASAP7_75t_L g459 ( 
.A1(n_440),
.A2(n_451),
.B1(n_33),
.B2(n_431),
.Y(n_459)
);

XNOR2xp5_ASAP7_75t_L g461 ( 
.A(n_442),
.B(n_446),
.Y(n_461)
);

AOI22xp5_ASAP7_75t_L g445 ( 
.A1(n_423),
.A2(n_415),
.B1(n_405),
.B2(n_401),
.Y(n_445)
);

OAI22xp5_ASAP7_75t_L g463 ( 
.A1(n_445),
.A2(n_449),
.B1(n_453),
.B2(n_440),
.Y(n_463)
);

NAND2xp5_ASAP7_75t_L g455 ( 
.A(n_447),
.B(n_452),
.Y(n_455)
);

AOI21xp5_ASAP7_75t_L g448 ( 
.A1(n_421),
.A2(n_131),
.B(n_107),
.Y(n_448)
);

AOI21xp5_ASAP7_75t_L g456 ( 
.A1(n_448),
.A2(n_426),
.B(n_438),
.Y(n_456)
);

AOI22xp5_ASAP7_75t_L g449 ( 
.A1(n_435),
.A2(n_118),
.B1(n_134),
.B2(n_121),
.Y(n_449)
);

AOI211xp5_ASAP7_75t_L g451 ( 
.A1(n_427),
.A2(n_189),
.B(n_22),
.C(n_24),
.Y(n_451)
);

NOR2xp33_ASAP7_75t_SL g452 ( 
.A(n_430),
.B(n_127),
.Y(n_452)
);

AOI22xp5_ASAP7_75t_SL g453 ( 
.A1(n_422),
.A2(n_106),
.B1(n_107),
.B2(n_189),
.Y(n_453)
);

NAND2xp5_ASAP7_75t_L g465 ( 
.A(n_454),
.B(n_129),
.Y(n_465)
);

INVx1_ASAP7_75t_L g471 ( 
.A(n_456),
.Y(n_471)
);

NOR2xp33_ASAP7_75t_L g457 ( 
.A(n_444),
.B(n_420),
.Y(n_457)
);

INVx1_ASAP7_75t_L g472 ( 
.A(n_457),
.Y(n_472)
);

MAJIxp5_ASAP7_75t_L g458 ( 
.A(n_441),
.B(n_437),
.C(n_434),
.Y(n_458)
);

NAND2xp5_ASAP7_75t_SL g468 ( 
.A(n_458),
.B(n_464),
.Y(n_468)
);

INVx1_ASAP7_75t_L g477 ( 
.A(n_459),
.Y(n_477)
);

AOI21xp5_ASAP7_75t_L g460 ( 
.A1(n_439),
.A2(n_432),
.B(n_436),
.Y(n_460)
);

OAI21xp5_ASAP7_75t_SL g475 ( 
.A1(n_460),
.A2(n_466),
.B(n_455),
.Y(n_475)
);

NOR2xp33_ASAP7_75t_L g473 ( 
.A(n_463),
.B(n_465),
.Y(n_473)
);

NOR2xp33_ASAP7_75t_SL g464 ( 
.A(n_446),
.B(n_106),
.Y(n_464)
);

AOI21xp5_ASAP7_75t_SL g466 ( 
.A1(n_445),
.A2(n_33),
.B(n_78),
.Y(n_466)
);

MAJIxp5_ASAP7_75t_L g467 ( 
.A(n_443),
.B(n_78),
.C(n_20),
.Y(n_467)
);

MAJIxp5_ASAP7_75t_L g474 ( 
.A(n_467),
.B(n_1),
.C(n_2),
.Y(n_474)
);

NOR2xp67_ASAP7_75t_L g469 ( 
.A(n_461),
.B(n_454),
.Y(n_469)
);

OAI321xp33_ASAP7_75t_L g484 ( 
.A1(n_469),
.A2(n_470),
.A3(n_1),
.B1(n_3),
.B2(n_4),
.C(n_5),
.Y(n_484)
);

AOI322xp5_ASAP7_75t_L g470 ( 
.A1(n_462),
.A2(n_450),
.A3(n_453),
.B1(n_449),
.B2(n_447),
.C1(n_5),
.C2(n_6),
.Y(n_470)
);

INVx1_ASAP7_75t_L g479 ( 
.A(n_474),
.Y(n_479)
);

NOR2xp33_ASAP7_75t_L g482 ( 
.A(n_475),
.B(n_1),
.Y(n_482)
);

NOR2xp33_ASAP7_75t_L g476 ( 
.A(n_461),
.B(n_11),
.Y(n_476)
);

NAND2xp5_ASAP7_75t_SL g481 ( 
.A(n_476),
.B(n_1),
.Y(n_481)
);

OAI21xp5_ASAP7_75t_L g478 ( 
.A1(n_472),
.A2(n_466),
.B(n_458),
.Y(n_478)
);

AOI22x1_ASAP7_75t_L g488 ( 
.A1(n_478),
.A2(n_483),
.B1(n_5),
.B2(n_6),
.Y(n_488)
);

AOI21xp5_ASAP7_75t_L g480 ( 
.A1(n_471),
.A2(n_467),
.B(n_2),
.Y(n_480)
);

AOI22xp5_ASAP7_75t_L g485 ( 
.A1(n_480),
.A2(n_482),
.B1(n_484),
.B2(n_477),
.Y(n_485)
);

NOR2xp33_ASAP7_75t_SL g487 ( 
.A(n_481),
.B(n_5),
.Y(n_487)
);

OAI21xp5_ASAP7_75t_L g483 ( 
.A1(n_475),
.A2(n_1),
.B(n_2),
.Y(n_483)
);

OAI21xp5_ASAP7_75t_L g492 ( 
.A1(n_485),
.A2(n_486),
.B(n_488),
.Y(n_492)
);

AOI322xp5_ASAP7_75t_L g486 ( 
.A1(n_479),
.A2(n_473),
.A3(n_468),
.B1(n_474),
.B2(n_8),
.C1(n_9),
.C2(n_5),
.Y(n_486)
);

NOR3xp33_ASAP7_75t_L g491 ( 
.A(n_487),
.B(n_6),
.C(n_9),
.Y(n_491)
);

A2O1A1O1Ixp25_ASAP7_75t_L g489 ( 
.A1(n_478),
.A2(n_6),
.B(n_7),
.C(n_9),
.D(n_10),
.Y(n_489)
);

OAI21xp5_ASAP7_75t_SL g490 ( 
.A1(n_489),
.A2(n_11),
.B(n_7),
.Y(n_490)
);

OAI21xp5_ASAP7_75t_SL g493 ( 
.A1(n_490),
.A2(n_491),
.B(n_492),
.Y(n_493)
);

NAND2xp5_ASAP7_75t_L g494 ( 
.A(n_493),
.B(n_6),
.Y(n_494)
);

NAND2xp5_ASAP7_75t_L g495 ( 
.A(n_494),
.B(n_10),
.Y(n_495)
);

XOR2xp5_ASAP7_75t_L g496 ( 
.A(n_495),
.B(n_11),
.Y(n_496)
);


endmodule