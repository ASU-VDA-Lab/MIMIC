module fake_netlist_6_4716_n_109 (n_41, n_16, n_45, n_1, n_46, n_34, n_42, n_9, n_8, n_18, n_10, n_21, n_24, n_37, n_6, n_15, n_33, n_27, n_3, n_14, n_38, n_0, n_39, n_32, n_4, n_36, n_22, n_26, n_13, n_35, n_11, n_28, n_17, n_23, n_12, n_20, n_50, n_49, n_7, n_30, n_2, n_43, n_5, n_19, n_47, n_48, n_29, n_31, n_25, n_40, n_44, n_109);

input n_41;
input n_16;
input n_45;
input n_1;
input n_46;
input n_34;
input n_42;
input n_9;
input n_8;
input n_18;
input n_10;
input n_21;
input n_24;
input n_37;
input n_6;
input n_15;
input n_33;
input n_27;
input n_3;
input n_14;
input n_38;
input n_0;
input n_39;
input n_32;
input n_4;
input n_36;
input n_22;
input n_26;
input n_13;
input n_35;
input n_11;
input n_28;
input n_17;
input n_23;
input n_12;
input n_20;
input n_50;
input n_49;
input n_7;
input n_30;
input n_2;
input n_43;
input n_5;
input n_19;
input n_47;
input n_48;
input n_29;
input n_31;
input n_25;
input n_40;
input n_44;

output n_109;

wire n_52;
wire n_91;
wire n_88;
wire n_98;
wire n_63;
wire n_73;
wire n_68;
wire n_83;
wire n_101;
wire n_77;
wire n_106;
wire n_92;
wire n_96;
wire n_90;
wire n_105;
wire n_54;
wire n_102;
wire n_87;
wire n_85;
wire n_66;
wire n_99;
wire n_78;
wire n_84;
wire n_100;
wire n_62;
wire n_75;
wire n_70;
wire n_67;
wire n_82;
wire n_61;
wire n_81;
wire n_59;
wire n_76;
wire n_55;
wire n_94;
wire n_97;
wire n_108;
wire n_58;
wire n_64;
wire n_65;
wire n_93;
wire n_80;
wire n_86;
wire n_104;
wire n_95;
wire n_107;
wire n_71;
wire n_74;
wire n_72;
wire n_89;
wire n_103;
wire n_60;
wire n_69;
wire n_79;
wire n_57;
wire n_53;
wire n_51;
wire n_56;

OA21x2_ASAP7_75t_L g51 ( 
.A1(n_35),
.A2(n_18),
.B(n_8),
.Y(n_51)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_50),
.Y(n_52)
);

INVx2_ASAP7_75t_L g53 ( 
.A(n_21),
.Y(n_53)
);

HB1xp67_ASAP7_75t_L g54 ( 
.A(n_40),
.Y(n_54)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_24),
.Y(n_55)
);

HB1xp67_ASAP7_75t_L g56 ( 
.A(n_16),
.Y(n_56)
);

AND2x6_ASAP7_75t_L g57 ( 
.A(n_3),
.B(n_5),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_SL g58 ( 
.A(n_39),
.B(n_31),
.Y(n_58)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_4),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_L g60 ( 
.A(n_30),
.B(n_13),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_28),
.B(n_11),
.Y(n_61)
);

OAI21x1_ASAP7_75t_L g62 ( 
.A1(n_32),
.A2(n_26),
.B(n_2),
.Y(n_62)
);

HB1xp67_ASAP7_75t_L g63 ( 
.A(n_9),
.Y(n_63)
);

AND2x2_ASAP7_75t_L g64 ( 
.A(n_33),
.B(n_19),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_48),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_L g66 ( 
.A(n_38),
.B(n_1),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_L g67 ( 
.A(n_22),
.B(n_6),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_L g68 ( 
.A(n_46),
.B(n_25),
.Y(n_68)
);

AOI22xp5_ASAP7_75t_L g69 ( 
.A1(n_37),
.A2(n_49),
.B1(n_15),
.B2(n_0),
.Y(n_69)
);

BUFx6f_ASAP7_75t_L g70 ( 
.A(n_23),
.Y(n_70)
);

AND2x4_ASAP7_75t_L g71 ( 
.A(n_27),
.B(n_45),
.Y(n_71)
);

INVx2_ASAP7_75t_L g72 ( 
.A(n_29),
.Y(n_72)
);

BUFx6f_ASAP7_75t_L g73 ( 
.A(n_47),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_L g74 ( 
.A(n_7),
.B(n_34),
.Y(n_74)
);

BUFx6f_ASAP7_75t_L g75 ( 
.A(n_36),
.Y(n_75)
);

INVx2_ASAP7_75t_L g76 ( 
.A(n_52),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_L g77 ( 
.A(n_54),
.B(n_0),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_L g78 ( 
.A(n_56),
.B(n_10),
.Y(n_78)
);

NOR2xp67_ASAP7_75t_L g79 ( 
.A(n_63),
.B(n_12),
.Y(n_79)
);

NOR3xp33_ASAP7_75t_L g80 ( 
.A(n_58),
.B(n_14),
.C(n_17),
.Y(n_80)
);

AND2x2_ASAP7_75t_L g81 ( 
.A(n_53),
.B(n_20),
.Y(n_81)
);

BUFx6f_ASAP7_75t_L g82 ( 
.A(n_65),
.Y(n_82)
);

NAND3xp33_ASAP7_75t_L g83 ( 
.A(n_69),
.B(n_41),
.C(n_42),
.Y(n_83)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_55),
.Y(n_84)
);

BUFx2_ASAP7_75t_L g85 ( 
.A(n_59),
.Y(n_85)
);

AOI22xp5_ASAP7_75t_L g86 ( 
.A1(n_64),
.A2(n_43),
.B1(n_44),
.B2(n_57),
.Y(n_86)
);

AOI21xp5_ASAP7_75t_L g87 ( 
.A1(n_78),
.A2(n_67),
.B(n_74),
.Y(n_87)
);

AND2x2_ASAP7_75t_SL g88 ( 
.A(n_80),
.B(n_71),
.Y(n_88)
);

INVx1_ASAP7_75t_SL g89 ( 
.A(n_85),
.Y(n_89)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_82),
.Y(n_90)
);

NAND3xp33_ASAP7_75t_SL g91 ( 
.A(n_77),
.B(n_66),
.C(n_60),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_SL g92 ( 
.A(n_79),
.B(n_72),
.Y(n_92)
);

OAI21x1_ASAP7_75t_L g93 ( 
.A1(n_81),
.A2(n_62),
.B(n_68),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_L g94 ( 
.A(n_88),
.B(n_84),
.Y(n_94)
);

OR2x6_ASAP7_75t_L g95 ( 
.A(n_90),
.B(n_83),
.Y(n_95)
);

AND2x2_ASAP7_75t_L g96 ( 
.A(n_89),
.B(n_76),
.Y(n_96)
);

OAI21x1_ASAP7_75t_L g97 ( 
.A1(n_93),
.A2(n_86),
.B(n_51),
.Y(n_97)
);

OAI21x1_ASAP7_75t_L g98 ( 
.A1(n_87),
.A2(n_61),
.B(n_57),
.Y(n_98)
);

INVx2_ASAP7_75t_L g99 ( 
.A(n_96),
.Y(n_99)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_94),
.Y(n_100)
);

OR2x2_ASAP7_75t_L g101 ( 
.A(n_95),
.B(n_91),
.Y(n_101)
);

AND2x4_ASAP7_75t_L g102 ( 
.A(n_99),
.B(n_97),
.Y(n_102)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_102),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_L g104 ( 
.A(n_103),
.B(n_100),
.Y(n_104)
);

AND2x4_ASAP7_75t_L g105 ( 
.A(n_104),
.B(n_101),
.Y(n_105)
);

INVx3_ASAP7_75t_L g106 ( 
.A(n_105),
.Y(n_106)
);

OAI21xp33_ASAP7_75t_L g107 ( 
.A1(n_106),
.A2(n_92),
.B(n_98),
.Y(n_107)
);

AOI22xp33_ASAP7_75t_SL g108 ( 
.A1(n_107),
.A2(n_70),
.B1(n_73),
.B2(n_75),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_SL g109 ( 
.A(n_108),
.B(n_82),
.Y(n_109)
);


endmodule