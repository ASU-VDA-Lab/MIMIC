module fake_jpeg_4513_n_322 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_322);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_322;

wire n_253;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_15;
wire n_141;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

BUFx12_ASAP7_75t_L g15 ( 
.A(n_6),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_7),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_10),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_12),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_8),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_0),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_8),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_1),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_3),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_0),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_9),
.Y(n_25)
);

BUFx3_ASAP7_75t_L g26 ( 
.A(n_9),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_9),
.Y(n_27)
);

CKINVDCx16_ASAP7_75t_R g28 ( 
.A(n_10),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_2),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_4),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_4),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_4),
.Y(n_32)
);

CKINVDCx16_ASAP7_75t_R g33 ( 
.A(n_3),
.Y(n_33)
);

BUFx12_ASAP7_75t_L g34 ( 
.A(n_1),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_6),
.Y(n_35)
);

BUFx12f_ASAP7_75t_L g36 ( 
.A(n_1),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_11),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_2),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_22),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_SL g64 ( 
.A(n_39),
.B(n_42),
.Y(n_64)
);

INVx5_ASAP7_75t_L g40 ( 
.A(n_15),
.Y(n_40)
);

INVx5_ASAP7_75t_L g80 ( 
.A(n_40),
.Y(n_80)
);

INVx2_ASAP7_75t_L g41 ( 
.A(n_26),
.Y(n_41)
);

INVx8_ASAP7_75t_L g105 ( 
.A(n_41),
.Y(n_105)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_22),
.Y(n_42)
);

NAND2xp5_ASAP7_75t_L g43 ( 
.A(n_20),
.B(n_0),
.Y(n_43)
);

NAND2xp5_ASAP7_75t_L g76 ( 
.A(n_43),
.B(n_45),
.Y(n_76)
);

BUFx5_ASAP7_75t_L g44 ( 
.A(n_34),
.Y(n_44)
);

BUFx3_ASAP7_75t_L g93 ( 
.A(n_44),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_L g45 ( 
.A(n_20),
.B(n_0),
.Y(n_45)
);

INVx3_ASAP7_75t_L g46 ( 
.A(n_15),
.Y(n_46)
);

INVx5_ASAP7_75t_L g89 ( 
.A(n_46),
.Y(n_89)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_30),
.Y(n_47)
);

INVx6_ASAP7_75t_L g63 ( 
.A(n_47),
.Y(n_63)
);

INVx3_ASAP7_75t_L g48 ( 
.A(n_15),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_48),
.B(n_49),
.Y(n_81)
);

HB1xp67_ASAP7_75t_L g49 ( 
.A(n_30),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_17),
.B(n_8),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_SL g68 ( 
.A(n_50),
.B(n_58),
.Y(n_68)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_26),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_L g91 ( 
.A(n_51),
.B(n_56),
.Y(n_91)
);

INVx11_ASAP7_75t_L g52 ( 
.A(n_30),
.Y(n_52)
);

INVx6_ASAP7_75t_L g85 ( 
.A(n_52),
.Y(n_85)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_30),
.Y(n_53)
);

INVx6_ASAP7_75t_L g97 ( 
.A(n_53),
.Y(n_97)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_32),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g96 ( 
.A(n_54),
.Y(n_96)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_32),
.Y(n_55)
);

BUFx3_ASAP7_75t_L g99 ( 
.A(n_55),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_SL g56 ( 
.A(n_16),
.B(n_7),
.Y(n_56)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_26),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_L g92 ( 
.A(n_57),
.B(n_59),
.Y(n_92)
);

CKINVDCx20_ASAP7_75t_R g58 ( 
.A(n_24),
.Y(n_58)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_20),
.Y(n_59)
);

INVx3_ASAP7_75t_L g60 ( 
.A(n_15),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_60),
.B(n_32),
.Y(n_82)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_17),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_L g104 ( 
.A(n_61),
.B(n_62),
.Y(n_104)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_17),
.Y(n_62)
);

AOI22xp33_ASAP7_75t_SL g65 ( 
.A1(n_52),
.A2(n_33),
.B1(n_18),
.B2(n_28),
.Y(n_65)
);

AOI22xp33_ASAP7_75t_SL g126 ( 
.A1(n_65),
.A2(n_70),
.B1(n_71),
.B2(n_84),
.Y(n_126)
);

OAI22xp33_ASAP7_75t_SL g66 ( 
.A1(n_52),
.A2(n_38),
.B1(n_29),
.B2(n_24),
.Y(n_66)
);

OAI22xp33_ASAP7_75t_SL g133 ( 
.A1(n_66),
.A2(n_72),
.B1(n_101),
.B2(n_87),
.Y(n_133)
);

INVx4_ASAP7_75t_L g67 ( 
.A(n_40),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g119 ( 
.A(n_67),
.B(n_69),
.Y(n_119)
);

INVx2_ASAP7_75t_L g69 ( 
.A(n_44),
.Y(n_69)
);

AOI22xp33_ASAP7_75t_SL g70 ( 
.A1(n_46),
.A2(n_33),
.B1(n_18),
.B2(n_28),
.Y(n_70)
);

AOI22xp33_ASAP7_75t_SL g71 ( 
.A1(n_48),
.A2(n_18),
.B1(n_38),
.B2(n_29),
.Y(n_71)
);

OAI22xp5_ASAP7_75t_L g72 ( 
.A1(n_39),
.A2(n_16),
.B1(n_35),
.B2(n_31),
.Y(n_72)
);

OR2x2_ASAP7_75t_L g73 ( 
.A(n_42),
.B(n_37),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g139 ( 
.A(n_73),
.B(n_86),
.Y(n_139)
);

BUFx12f_ASAP7_75t_L g74 ( 
.A(n_60),
.Y(n_74)
);

CKINVDCx20_ASAP7_75t_R g121 ( 
.A(n_74),
.Y(n_121)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_43),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g131 ( 
.A(n_75),
.B(n_77),
.Y(n_131)
);

INVx4_ASAP7_75t_L g77 ( 
.A(n_49),
.Y(n_77)
);

INVx3_ASAP7_75t_L g78 ( 
.A(n_41),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g143 ( 
.A(n_78),
.B(n_100),
.Y(n_143)
);

INVx2_ASAP7_75t_L g79 ( 
.A(n_47),
.Y(n_79)
);

HB1xp67_ASAP7_75t_L g125 ( 
.A(n_79),
.Y(n_125)
);

INVxp33_ASAP7_75t_L g114 ( 
.A(n_82),
.Y(n_114)
);

OAI22xp33_ASAP7_75t_L g83 ( 
.A1(n_47),
.A2(n_32),
.B1(n_36),
.B2(n_35),
.Y(n_83)
);

OAI22xp5_ASAP7_75t_L g142 ( 
.A1(n_83),
.A2(n_87),
.B1(n_90),
.B2(n_34),
.Y(n_142)
);

AOI22xp33_ASAP7_75t_SL g84 ( 
.A1(n_51),
.A2(n_37),
.B1(n_19),
.B2(n_21),
.Y(n_84)
);

INVx3_ASAP7_75t_L g86 ( 
.A(n_53),
.Y(n_86)
);

AOI22xp33_ASAP7_75t_L g87 ( 
.A1(n_57),
.A2(n_19),
.B1(n_31),
.B2(n_21),
.Y(n_87)
);

INVx4_ASAP7_75t_L g88 ( 
.A(n_53),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g141 ( 
.A(n_88),
.B(n_98),
.Y(n_141)
);

AOI22xp33_ASAP7_75t_L g90 ( 
.A1(n_58),
.A2(n_23),
.B1(n_27),
.B2(n_25),
.Y(n_90)
);

BUFx12f_ASAP7_75t_L g94 ( 
.A(n_54),
.Y(n_94)
);

CKINVDCx20_ASAP7_75t_R g124 ( 
.A(n_94),
.Y(n_124)
);

INVx2_ASAP7_75t_L g95 ( 
.A(n_54),
.Y(n_95)
);

INVx3_ASAP7_75t_L g128 ( 
.A(n_95),
.Y(n_128)
);

INVx4_ASAP7_75t_L g98 ( 
.A(n_55),
.Y(n_98)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_45),
.Y(n_100)
);

OR2x2_ASAP7_75t_L g101 ( 
.A(n_56),
.B(n_62),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_SL g140 ( 
.A(n_101),
.B(n_106),
.Y(n_140)
);

CKINVDCx20_ASAP7_75t_R g102 ( 
.A(n_50),
.Y(n_102)
);

CKINVDCx20_ASAP7_75t_R g127 ( 
.A(n_102),
.Y(n_127)
);

INVx2_ASAP7_75t_L g103 ( 
.A(n_55),
.Y(n_103)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_103),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_L g106 ( 
.A(n_61),
.B(n_27),
.Y(n_106)
);

INVx2_ASAP7_75t_L g107 ( 
.A(n_59),
.Y(n_107)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_107),
.Y(n_118)
);

INVx3_ASAP7_75t_L g108 ( 
.A(n_40),
.Y(n_108)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_108),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_L g109 ( 
.A(n_43),
.B(n_25),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_L g115 ( 
.A(n_109),
.B(n_23),
.Y(n_115)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_43),
.Y(n_110)
);

INVx1_ASAP7_75t_SL g135 ( 
.A(n_110),
.Y(n_135)
);

INVx3_ASAP7_75t_L g111 ( 
.A(n_40),
.Y(n_111)
);

INVx4_ASAP7_75t_L g116 ( 
.A(n_111),
.Y(n_116)
);

AOI22x1_ASAP7_75t_L g112 ( 
.A1(n_83),
.A2(n_36),
.B1(n_34),
.B2(n_15),
.Y(n_112)
);

OAI22xp5_ASAP7_75t_SL g175 ( 
.A1(n_112),
.A2(n_122),
.B1(n_124),
.B2(n_128),
.Y(n_175)
);

NOR2xp33_ASAP7_75t_SL g149 ( 
.A(n_115),
.B(n_84),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_L g117 ( 
.A(n_76),
.B(n_36),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_L g145 ( 
.A(n_117),
.B(n_129),
.Y(n_145)
);

INVx2_ASAP7_75t_L g120 ( 
.A(n_99),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_L g155 ( 
.A(n_120),
.B(n_123),
.Y(n_155)
);

OA22x2_ASAP7_75t_L g122 ( 
.A1(n_80),
.A2(n_36),
.B1(n_34),
.B2(n_3),
.Y(n_122)
);

BUFx6f_ASAP7_75t_L g123 ( 
.A(n_89),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_L g129 ( 
.A(n_104),
.B(n_36),
.Y(n_129)
);

INVx2_ASAP7_75t_L g130 ( 
.A(n_99),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_L g132 ( 
.A(n_91),
.B(n_1),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_L g172 ( 
.A(n_132),
.B(n_138),
.Y(n_172)
);

AOI22xp33_ASAP7_75t_L g154 ( 
.A1(n_133),
.A2(n_66),
.B1(n_73),
.B2(n_34),
.Y(n_154)
);

AOI22xp33_ASAP7_75t_SL g134 ( 
.A1(n_63),
.A2(n_10),
.B1(n_14),
.B2(n_5),
.Y(n_134)
);

AOI22xp33_ASAP7_75t_SL g165 ( 
.A1(n_134),
.A2(n_12),
.B1(n_13),
.B2(n_14),
.Y(n_165)
);

AOI22xp33_ASAP7_75t_L g136 ( 
.A1(n_63),
.A2(n_11),
.B1(n_14),
.B2(n_5),
.Y(n_136)
);

OAI22xp5_ASAP7_75t_L g152 ( 
.A1(n_136),
.A2(n_90),
.B1(n_70),
.B2(n_68),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_L g138 ( 
.A(n_92),
.B(n_2),
.Y(n_138)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_142),
.Y(n_146)
);

AOI22xp5_ASAP7_75t_L g144 ( 
.A1(n_142),
.A2(n_97),
.B1(n_105),
.B2(n_85),
.Y(n_144)
);

OAI22xp5_ASAP7_75t_SL g202 ( 
.A1(n_144),
.A2(n_147),
.B1(n_116),
.B2(n_146),
.Y(n_202)
);

AOI22xp5_ASAP7_75t_L g147 ( 
.A1(n_117),
.A2(n_97),
.B1(n_105),
.B2(n_85),
.Y(n_147)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_143),
.Y(n_148)
);

NOR2xp33_ASAP7_75t_L g203 ( 
.A(n_148),
.B(n_150),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_SL g211 ( 
.A(n_149),
.B(n_166),
.Y(n_211)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_143),
.Y(n_150)
);

AOI21xp5_ASAP7_75t_L g151 ( 
.A1(n_126),
.A2(n_71),
.B(n_65),
.Y(n_151)
);

OAI21xp5_ASAP7_75t_SL g195 ( 
.A1(n_151),
.A2(n_157),
.B(n_167),
.Y(n_195)
);

AOI22xp33_ASAP7_75t_L g208 ( 
.A1(n_152),
.A2(n_158),
.B1(n_160),
.B2(n_150),
.Y(n_208)
);

MAJIxp5_ASAP7_75t_L g153 ( 
.A(n_129),
.B(n_81),
.C(n_64),
.Y(n_153)
);

MAJIxp5_ASAP7_75t_L g181 ( 
.A(n_153),
.B(n_172),
.C(n_170),
.Y(n_181)
);

OAI22xp5_ASAP7_75t_L g204 ( 
.A1(n_154),
.A2(n_156),
.B1(n_165),
.B2(n_151),
.Y(n_204)
);

AOI22xp33_ASAP7_75t_L g156 ( 
.A1(n_112),
.A2(n_96),
.B1(n_94),
.B2(n_74),
.Y(n_156)
);

AND2x2_ASAP7_75t_L g157 ( 
.A(n_135),
.B(n_94),
.Y(n_157)
);

OAI21xp5_ASAP7_75t_L g158 ( 
.A1(n_140),
.A2(n_2),
.B(n_3),
.Y(n_158)
);

AOI21xp5_ASAP7_75t_L g210 ( 
.A1(n_158),
.A2(n_178),
.B(n_159),
.Y(n_210)
);

NOR2xp33_ASAP7_75t_L g159 ( 
.A(n_140),
.B(n_5),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_SL g186 ( 
.A(n_159),
.B(n_162),
.Y(n_186)
);

OA22x2_ASAP7_75t_L g160 ( 
.A1(n_112),
.A2(n_96),
.B1(n_74),
.B2(n_93),
.Y(n_160)
);

AO22x1_ASAP7_75t_SL g197 ( 
.A1(n_160),
.A2(n_123),
.B1(n_116),
.B2(n_137),
.Y(n_197)
);

CKINVDCx20_ASAP7_75t_R g161 ( 
.A(n_131),
.Y(n_161)
);

CKINVDCx20_ASAP7_75t_R g180 ( 
.A(n_161),
.Y(n_180)
);

NOR2xp33_ASAP7_75t_L g162 ( 
.A(n_127),
.B(n_6),
.Y(n_162)
);

NOR2xp33_ASAP7_75t_SL g163 ( 
.A(n_127),
.B(n_7),
.Y(n_163)
);

NOR2xp33_ASAP7_75t_L g164 ( 
.A(n_138),
.B(n_11),
.Y(n_164)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_141),
.Y(n_166)
);

AND2x2_ASAP7_75t_L g167 ( 
.A(n_135),
.B(n_12),
.Y(n_167)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_141),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_L g184 ( 
.A(n_168),
.B(n_170),
.Y(n_184)
);

INVx1_ASAP7_75t_SL g169 ( 
.A(n_122),
.Y(n_169)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_169),
.Y(n_188)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_139),
.Y(n_170)
);

INVx1_ASAP7_75t_SL g171 ( 
.A(n_122),
.Y(n_171)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_171),
.Y(n_191)
);

AND2x2_ASAP7_75t_L g173 ( 
.A(n_132),
.B(n_13),
.Y(n_173)
);

AND2x2_ASAP7_75t_L g196 ( 
.A(n_173),
.B(n_175),
.Y(n_196)
);

NOR2xp33_ASAP7_75t_L g174 ( 
.A(n_114),
.B(n_121),
.Y(n_174)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_174),
.Y(n_192)
);

AND2x2_ASAP7_75t_L g176 ( 
.A(n_115),
.B(n_122),
.Y(n_176)
);

AND2x2_ASAP7_75t_L g199 ( 
.A(n_176),
.B(n_137),
.Y(n_199)
);

NOR2xp33_ASAP7_75t_L g177 ( 
.A(n_139),
.B(n_123),
.Y(n_177)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_177),
.Y(n_194)
);

OAI21x1_ASAP7_75t_SL g178 ( 
.A1(n_125),
.A2(n_128),
.B(n_113),
.Y(n_178)
);

AOI22xp5_ASAP7_75t_L g179 ( 
.A1(n_146),
.A2(n_113),
.B1(n_130),
.B2(n_120),
.Y(n_179)
);

OAI22xp5_ASAP7_75t_SL g231 ( 
.A1(n_179),
.A2(n_208),
.B1(n_169),
.B2(n_171),
.Y(n_231)
);

XNOR2xp5_ASAP7_75t_L g232 ( 
.A(n_181),
.B(n_152),
.Y(n_232)
);

CKINVDCx16_ASAP7_75t_R g182 ( 
.A(n_155),
.Y(n_182)
);

NOR2xp33_ASAP7_75t_L g214 ( 
.A(n_182),
.B(n_190),
.Y(n_214)
);

MAJIxp5_ASAP7_75t_L g183 ( 
.A(n_145),
.B(n_121),
.C(n_124),
.Y(n_183)
);

MAJIxp5_ASAP7_75t_L g213 ( 
.A(n_183),
.B(n_209),
.C(n_187),
.Y(n_213)
);

CKINVDCx20_ASAP7_75t_R g185 ( 
.A(n_178),
.Y(n_185)
);

CKINVDCx20_ASAP7_75t_R g221 ( 
.A(n_185),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_L g187 ( 
.A(n_145),
.B(n_118),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_L g212 ( 
.A(n_187),
.B(n_198),
.Y(n_212)
);

CKINVDCx20_ASAP7_75t_R g189 ( 
.A(n_161),
.Y(n_189)
);

CKINVDCx20_ASAP7_75t_R g219 ( 
.A(n_189),
.Y(n_219)
);

CKINVDCx20_ASAP7_75t_R g190 ( 
.A(n_162),
.Y(n_190)
);

OAI21xp5_ASAP7_75t_L g193 ( 
.A1(n_149),
.A2(n_119),
.B(n_118),
.Y(n_193)
);

AOI21xp5_ASAP7_75t_L g234 ( 
.A1(n_193),
.A2(n_167),
.B(n_173),
.Y(n_234)
);

OAI22xp33_ASAP7_75t_SL g230 ( 
.A1(n_197),
.A2(n_166),
.B1(n_168),
.B2(n_157),
.Y(n_230)
);

CKINVDCx20_ASAP7_75t_R g198 ( 
.A(n_177),
.Y(n_198)
);

AOI22xp5_ASAP7_75t_L g220 ( 
.A1(n_199),
.A2(n_202),
.B1(n_204),
.B2(n_175),
.Y(n_220)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_147),
.Y(n_200)
);

NAND2xp5_ASAP7_75t_L g216 ( 
.A(n_200),
.B(n_201),
.Y(n_216)
);

CKINVDCx20_ASAP7_75t_R g201 ( 
.A(n_163),
.Y(n_201)
);

CKINVDCx20_ASAP7_75t_R g205 ( 
.A(n_157),
.Y(n_205)
);

NAND2xp5_ASAP7_75t_L g227 ( 
.A(n_205),
.B(n_209),
.Y(n_227)
);

BUFx2_ASAP7_75t_L g206 ( 
.A(n_160),
.Y(n_206)
);

BUFx6f_ASAP7_75t_L g229 ( 
.A(n_206),
.Y(n_229)
);

CKINVDCx16_ASAP7_75t_R g207 ( 
.A(n_144),
.Y(n_207)
);

NOR2xp33_ASAP7_75t_SL g222 ( 
.A(n_207),
.B(n_176),
.Y(n_222)
);

NAND2xp5_ASAP7_75t_L g209 ( 
.A(n_172),
.B(n_176),
.Y(n_209)
);

OAI21xp5_ASAP7_75t_L g233 ( 
.A1(n_210),
.A2(n_164),
.B(n_167),
.Y(n_233)
);

MAJIxp5_ASAP7_75t_L g257 ( 
.A(n_213),
.B(n_190),
.C(n_186),
.Y(n_257)
);

CKINVDCx16_ASAP7_75t_R g215 ( 
.A(n_203),
.Y(n_215)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_215),
.Y(n_238)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_179),
.Y(n_217)
);

NAND2xp5_ASAP7_75t_L g249 ( 
.A(n_217),
.B(n_218),
.Y(n_249)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_184),
.Y(n_218)
);

OAI22xp5_ASAP7_75t_SL g255 ( 
.A1(n_220),
.A2(n_192),
.B1(n_210),
.B2(n_180),
.Y(n_255)
);

CKINVDCx14_ASAP7_75t_R g237 ( 
.A(n_222),
.Y(n_237)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_184),
.Y(n_223)
);

NAND2xp5_ASAP7_75t_L g251 ( 
.A(n_223),
.B(n_224),
.Y(n_251)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_183),
.Y(n_224)
);

OAI21xp5_ASAP7_75t_SL g225 ( 
.A1(n_211),
.A2(n_160),
.B(n_148),
.Y(n_225)
);

AOI21xp5_ASAP7_75t_L g256 ( 
.A1(n_225),
.A2(n_234),
.B(n_236),
.Y(n_256)
);

AOI22xp5_ASAP7_75t_L g226 ( 
.A1(n_202),
.A2(n_200),
.B1(n_196),
.B2(n_185),
.Y(n_226)
);

OAI22xp5_ASAP7_75t_L g244 ( 
.A1(n_226),
.A2(n_197),
.B1(n_188),
.B2(n_191),
.Y(n_244)
);

XOR2xp5_ASAP7_75t_L g228 ( 
.A(n_195),
.B(n_153),
.Y(n_228)
);

MAJIxp5_ASAP7_75t_L g242 ( 
.A(n_228),
.B(n_232),
.C(n_235),
.Y(n_242)
);

AO21x1_ASAP7_75t_L g240 ( 
.A1(n_230),
.A2(n_197),
.B(n_193),
.Y(n_240)
);

AOI22xp5_ASAP7_75t_L g248 ( 
.A1(n_231),
.A2(n_199),
.B1(n_196),
.B2(n_188),
.Y(n_248)
);

AOI21xp5_ASAP7_75t_SL g252 ( 
.A1(n_233),
.A2(n_199),
.B(n_196),
.Y(n_252)
);

XOR2xp5_ASAP7_75t_L g235 ( 
.A(n_195),
.B(n_173),
.Y(n_235)
);

OAI21xp5_ASAP7_75t_SL g236 ( 
.A1(n_198),
.A2(n_205),
.B(n_194),
.Y(n_236)
);

NAND3xp33_ASAP7_75t_L g239 ( 
.A(n_219),
.B(n_180),
.C(n_189),
.Y(n_239)
);

NOR2xp33_ASAP7_75t_L g260 ( 
.A(n_239),
.B(n_240),
.Y(n_260)
);

CKINVDCx20_ASAP7_75t_R g241 ( 
.A(n_214),
.Y(n_241)
);

NAND2xp5_ASAP7_75t_L g261 ( 
.A(n_241),
.B(n_243),
.Y(n_261)
);

CKINVDCx20_ASAP7_75t_R g243 ( 
.A(n_219),
.Y(n_243)
);

AOI22xp5_ASAP7_75t_L g262 ( 
.A1(n_244),
.A2(n_255),
.B1(n_231),
.B2(n_217),
.Y(n_262)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_212),
.Y(n_245)
);

NOR2xp33_ASAP7_75t_L g266 ( 
.A(n_245),
.B(n_246),
.Y(n_266)
);

CKINVDCx20_ASAP7_75t_R g246 ( 
.A(n_212),
.Y(n_246)
);

INVx2_ASAP7_75t_SL g247 ( 
.A(n_229),
.Y(n_247)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_247),
.Y(n_258)
);

OAI22xp5_ASAP7_75t_L g272 ( 
.A1(n_248),
.A2(n_252),
.B1(n_254),
.B2(n_234),
.Y(n_272)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_216),
.Y(n_250)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_250),
.Y(n_259)
);

MAJIxp5_ASAP7_75t_L g253 ( 
.A(n_224),
.B(n_181),
.C(n_194),
.Y(n_253)
);

MAJIxp5_ASAP7_75t_L g267 ( 
.A(n_253),
.B(n_257),
.C(n_213),
.Y(n_267)
);

AOI22xp5_ASAP7_75t_L g254 ( 
.A1(n_221),
.A2(n_191),
.B1(n_206),
.B2(n_192),
.Y(n_254)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_262),
.Y(n_276)
);

AOI22xp5_ASAP7_75t_L g263 ( 
.A1(n_255),
.A2(n_227),
.B1(n_220),
.B2(n_226),
.Y(n_263)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_263),
.Y(n_280)
);

INVx1_ASAP7_75t_SL g264 ( 
.A(n_247),
.Y(n_264)
);

NAND2xp5_ASAP7_75t_L g285 ( 
.A(n_264),
.B(n_268),
.Y(n_285)
);

AOI22xp5_ASAP7_75t_L g265 ( 
.A1(n_244),
.A2(n_227),
.B1(n_223),
.B2(n_218),
.Y(n_265)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_265),
.Y(n_284)
);

MAJIxp5_ASAP7_75t_L g274 ( 
.A(n_267),
.B(n_269),
.C(n_273),
.Y(n_274)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_249),
.Y(n_268)
);

MAJIxp5_ASAP7_75t_L g269 ( 
.A(n_242),
.B(n_228),
.C(n_235),
.Y(n_269)
);

AOI22xp5_ASAP7_75t_L g270 ( 
.A1(n_237),
.A2(n_216),
.B1(n_233),
.B2(n_236),
.Y(n_270)
);

CKINVDCx14_ASAP7_75t_R g283 ( 
.A(n_270),
.Y(n_283)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_249),
.Y(n_271)
);

NAND2xp5_ASAP7_75t_SL g287 ( 
.A(n_271),
.B(n_245),
.Y(n_287)
);

XNOR2xp5_ASAP7_75t_L g277 ( 
.A(n_272),
.B(n_256),
.Y(n_277)
);

XOR2xp5_ASAP7_75t_L g273 ( 
.A(n_242),
.B(n_232),
.Y(n_273)
);

NOR2xp33_ASAP7_75t_SL g275 ( 
.A(n_270),
.B(n_201),
.Y(n_275)
);

NAND2xp5_ASAP7_75t_SL g291 ( 
.A(n_275),
.B(n_260),
.Y(n_291)
);

XOR2xp5_ASAP7_75t_L g296 ( 
.A(n_277),
.B(n_282),
.Y(n_296)
);

MAJIxp5_ASAP7_75t_L g278 ( 
.A(n_273),
.B(n_253),
.C(n_252),
.Y(n_278)
);

MAJIxp5_ASAP7_75t_L g290 ( 
.A(n_278),
.B(n_279),
.C(n_251),
.Y(n_290)
);

MAJIxp5_ASAP7_75t_L g279 ( 
.A(n_269),
.B(n_251),
.C(n_257),
.Y(n_279)
);

NAND2xp5_ASAP7_75t_L g281 ( 
.A(n_261),
.B(n_250),
.Y(n_281)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_281),
.Y(n_288)
);

XNOR2xp5_ASAP7_75t_L g282 ( 
.A(n_267),
.B(n_256),
.Y(n_282)
);

BUFx12f_ASAP7_75t_SL g286 ( 
.A(n_261),
.Y(n_286)
);

AOI22xp5_ASAP7_75t_L g289 ( 
.A1(n_286),
.A2(n_259),
.B1(n_243),
.B2(n_266),
.Y(n_289)
);

NAND2xp5_ASAP7_75t_L g299 ( 
.A(n_287),
.B(n_246),
.Y(n_299)
);

XNOR2xp5_ASAP7_75t_SL g304 ( 
.A(n_289),
.B(n_281),
.Y(n_304)
);

MAJIxp5_ASAP7_75t_L g303 ( 
.A(n_290),
.B(n_293),
.C(n_295),
.Y(n_303)
);

NAND2xp5_ASAP7_75t_L g305 ( 
.A(n_291),
.B(n_294),
.Y(n_305)
);

BUFx24_ASAP7_75t_SL g292 ( 
.A(n_282),
.Y(n_292)
);

NOR2xp33_ASAP7_75t_L g300 ( 
.A(n_292),
.B(n_277),
.Y(n_300)
);

MAJIxp5_ASAP7_75t_L g293 ( 
.A(n_279),
.B(n_259),
.C(n_265),
.Y(n_293)
);

NOR2xp33_ASAP7_75t_L g294 ( 
.A(n_276),
.B(n_258),
.Y(n_294)
);

NAND2xp5_ASAP7_75t_SL g295 ( 
.A(n_280),
.B(n_238),
.Y(n_295)
);

OAI22xp5_ASAP7_75t_L g297 ( 
.A1(n_286),
.A2(n_262),
.B1(n_263),
.B2(n_248),
.Y(n_297)
);

NAND2xp5_ASAP7_75t_SL g301 ( 
.A(n_297),
.B(n_299),
.Y(n_301)
);

NOR2xp33_ASAP7_75t_L g298 ( 
.A(n_284),
.B(n_258),
.Y(n_298)
);

NAND2xp5_ASAP7_75t_L g307 ( 
.A(n_298),
.B(n_264),
.Y(n_307)
);

NOR2xp33_ASAP7_75t_SL g312 ( 
.A(n_300),
.B(n_296),
.Y(n_312)
);

XNOR2xp5_ASAP7_75t_L g302 ( 
.A(n_293),
.B(n_290),
.Y(n_302)
);

MAJIxp5_ASAP7_75t_L g310 ( 
.A(n_302),
.B(n_304),
.C(n_296),
.Y(n_310)
);

OR2x2_ASAP7_75t_L g306 ( 
.A(n_288),
.B(n_241),
.Y(n_306)
);

OR2x2_ASAP7_75t_L g308 ( 
.A(n_306),
.B(n_240),
.Y(n_308)
);

NAND2xp5_ASAP7_75t_L g311 ( 
.A(n_307),
.B(n_238),
.Y(n_311)
);

NAND2xp5_ASAP7_75t_SL g314 ( 
.A(n_308),
.B(n_309),
.Y(n_314)
);

OR2x2_ASAP7_75t_L g309 ( 
.A(n_301),
.B(n_240),
.Y(n_309)
);

NAND2xp5_ASAP7_75t_SL g316 ( 
.A(n_310),
.B(n_311),
.Y(n_316)
);

HB1xp67_ASAP7_75t_L g315 ( 
.A(n_312),
.Y(n_315)
);

OAI22xp5_ASAP7_75t_SL g313 ( 
.A1(n_301),
.A2(n_283),
.B1(n_278),
.B2(n_285),
.Y(n_313)
);

NAND2xp5_ASAP7_75t_L g317 ( 
.A(n_316),
.B(n_305),
.Y(n_317)
);

AOI322xp5_ASAP7_75t_L g319 ( 
.A1(n_317),
.A2(n_318),
.A3(n_315),
.B1(n_308),
.B2(n_274),
.C1(n_225),
.C2(n_254),
.Y(n_319)
);

AOI22xp5_ASAP7_75t_L g318 ( 
.A1(n_314),
.A2(n_313),
.B1(n_303),
.B2(n_309),
.Y(n_318)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_319),
.Y(n_320)
);

NAND2xp5_ASAP7_75t_L g321 ( 
.A(n_320),
.B(n_318),
.Y(n_321)
);

XOR2xp5_ASAP7_75t_L g322 ( 
.A(n_321),
.B(n_274),
.Y(n_322)
);


endmodule