module fake_jpeg_14478_n_54 (n_3, n_2, n_1, n_0, n_4, n_6, n_5, n_54);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_6;
input n_5;

output n_54;

wire n_13;
wire n_21;
wire n_53;
wire n_33;
wire n_45;
wire n_10;
wire n_23;
wire n_27;
wire n_22;
wire n_47;
wire n_51;
wire n_14;
wire n_40;
wire n_19;
wire n_18;
wire n_20;
wire n_35;
wire n_48;
wire n_52;
wire n_46;
wire n_41;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_16;
wire n_49;
wire n_24;
wire n_28;
wire n_44;
wire n_26;
wire n_38;
wire n_9;
wire n_36;
wire n_11;
wire n_17;
wire n_31;
wire n_25;
wire n_29;
wire n_37;
wire n_43;
wire n_50;
wire n_12;
wire n_32;
wire n_8;
wire n_15;
wire n_7;

INVx11_ASAP7_75t_SL g7 ( 
.A(n_2),
.Y(n_7)
);

INVx1_ASAP7_75t_L g8 ( 
.A(n_1),
.Y(n_8)
);

INVx1_ASAP7_75t_L g9 ( 
.A(n_3),
.Y(n_9)
);

INVx6_ASAP7_75t_L g10 ( 
.A(n_5),
.Y(n_10)
);

CKINVDCx20_ASAP7_75t_R g11 ( 
.A(n_4),
.Y(n_11)
);

BUFx10_ASAP7_75t_L g12 ( 
.A(n_1),
.Y(n_12)
);

INVx3_ASAP7_75t_L g13 ( 
.A(n_3),
.Y(n_13)
);

INVx1_ASAP7_75t_L g14 ( 
.A(n_5),
.Y(n_14)
);

NOR2xp33_ASAP7_75t_L g15 ( 
.A(n_4),
.B(n_2),
.Y(n_15)
);

INVx1_ASAP7_75t_SL g16 ( 
.A(n_6),
.Y(n_16)
);

OAI22xp5_ASAP7_75t_L g17 ( 
.A1(n_10),
.A2(n_0),
.B1(n_1),
.B2(n_6),
.Y(n_17)
);

NOR2xp33_ASAP7_75t_L g25 ( 
.A(n_17),
.B(n_18),
.Y(n_25)
);

OR2x2_ASAP7_75t_L g18 ( 
.A(n_8),
.B(n_0),
.Y(n_18)
);

INVx2_ASAP7_75t_L g19 ( 
.A(n_8),
.Y(n_19)
);

INVx2_ASAP7_75t_L g24 ( 
.A(n_19),
.Y(n_24)
);

NOR2xp33_ASAP7_75t_L g20 ( 
.A(n_16),
.B(n_0),
.Y(n_20)
);

NOR2xp33_ASAP7_75t_L g26 ( 
.A(n_20),
.B(n_21),
.Y(n_26)
);

NOR2xp33_ASAP7_75t_L g21 ( 
.A(n_16),
.B(n_15),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_9),
.Y(n_22)
);

NOR2xp33_ASAP7_75t_L g28 ( 
.A(n_22),
.B(n_23),
.Y(n_28)
);

HAxp5_ASAP7_75t_SL g23 ( 
.A(n_12),
.B(n_7),
.CON(n_23),
.SN(n_23)
);

BUFx3_ASAP7_75t_L g27 ( 
.A(n_19),
.Y(n_27)
);

BUFx12f_ASAP7_75t_L g38 ( 
.A(n_27),
.Y(n_38)
);

AOI22xp33_ASAP7_75t_L g29 ( 
.A1(n_22),
.A2(n_12),
.B1(n_13),
.B2(n_10),
.Y(n_29)
);

OAI22xp5_ASAP7_75t_L g35 ( 
.A1(n_29),
.A2(n_18),
.B1(n_12),
.B2(n_14),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g30 ( 
.A(n_21),
.B(n_11),
.Y(n_30)
);

AOI21xp5_ASAP7_75t_SL g33 ( 
.A1(n_30),
.A2(n_31),
.B(n_20),
.Y(n_33)
);

OAI21xp5_ASAP7_75t_L g31 ( 
.A1(n_18),
.A2(n_12),
.B(n_13),
.Y(n_31)
);

CKINVDCx14_ASAP7_75t_R g32 ( 
.A(n_28),
.Y(n_32)
);

OAI21xp5_ASAP7_75t_L g42 ( 
.A1(n_32),
.A2(n_33),
.B(n_37),
.Y(n_42)
);

INVx2_ASAP7_75t_L g34 ( 
.A(n_24),
.Y(n_34)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_34),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g41 ( 
.A(n_35),
.B(n_36),
.Y(n_41)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_24),
.Y(n_36)
);

OAI22xp5_ASAP7_75t_SL g37 ( 
.A1(n_25),
.A2(n_17),
.B1(n_9),
.B2(n_14),
.Y(n_37)
);

AOI21xp5_ASAP7_75t_L g39 ( 
.A1(n_32),
.A2(n_31),
.B(n_25),
.Y(n_39)
);

NAND2xp5_ASAP7_75t_SL g44 ( 
.A(n_39),
.B(n_28),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_40),
.Y(n_43)
);

NAND2xp5_ASAP7_75t_L g46 ( 
.A(n_43),
.B(n_45),
.Y(n_46)
);

MAJIxp5_ASAP7_75t_L g47 ( 
.A(n_44),
.B(n_42),
.C(n_30),
.Y(n_47)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_41),
.Y(n_45)
);

XNOR2xp5_ASAP7_75t_SL g49 ( 
.A(n_47),
.B(n_26),
.Y(n_49)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_46),
.Y(n_48)
);

HB1xp67_ASAP7_75t_L g50 ( 
.A(n_48),
.Y(n_50)
);

MAJIxp5_ASAP7_75t_L g51 ( 
.A(n_50),
.B(n_49),
.C(n_26),
.Y(n_51)
);

MAJIxp5_ASAP7_75t_L g52 ( 
.A(n_51),
.B(n_45),
.C(n_38),
.Y(n_52)
);

AOI21xp5_ASAP7_75t_L g53 ( 
.A1(n_52),
.A2(n_38),
.B(n_27),
.Y(n_53)
);

XOR2xp5_ASAP7_75t_L g54 ( 
.A(n_53),
.B(n_38),
.Y(n_54)
);


endmodule