module fake_jpeg_2460_n_114 (n_13, n_21, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_19, n_18, n_20, n_4, n_30, n_16, n_3, n_0, n_24, n_28, n_26, n_9, n_5, n_11, n_17, n_25, n_2, n_29, n_12, n_8, n_15, n_7, n_114);

input n_13;
input n_21;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_4;
input n_30;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_26;
input n_9;
input n_5;
input n_11;
input n_17;
input n_25;
input n_2;
input n_29;
input n_12;
input n_8;
input n_15;
input n_7;

output n_114;

wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_73;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_42;
wire n_49;
wire n_76;
wire n_38;
wire n_88;
wire n_74;
wire n_31;
wire n_103;
wire n_50;
wire n_57;
wire n_69;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_109;
wire n_113;
wire n_106;
wire n_111;
wire n_44;
wire n_75;
wire n_37;
wire n_102;
wire n_99;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_56;
wire n_79;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_101;
wire n_48;
wire n_35;
wire n_87;
wire n_46;
wire n_86;
wire n_112;
wire n_95;
wire n_97;
wire n_36;
wire n_62;
wire n_43;
wire n_32;
wire n_100;
wire n_82;
wire n_96;

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_22),
.Y(n_31)
);

BUFx2_ASAP7_75t_L g32 ( 
.A(n_10),
.Y(n_32)
);

INVx13_ASAP7_75t_L g33 ( 
.A(n_5),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_19),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_17),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_7),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_25),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_8),
.Y(n_38)
);

BUFx6f_ASAP7_75t_SL g39 ( 
.A(n_12),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_26),
.Y(n_40)
);

INVx3_ASAP7_75t_L g41 ( 
.A(n_1),
.Y(n_41)
);

BUFx3_ASAP7_75t_L g42 ( 
.A(n_13),
.Y(n_42)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_30),
.Y(n_43)
);

INVx3_ASAP7_75t_L g44 ( 
.A(n_41),
.Y(n_44)
);

INVx4_ASAP7_75t_L g54 ( 
.A(n_44),
.Y(n_54)
);

INVx2_ASAP7_75t_R g45 ( 
.A(n_33),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g57 ( 
.A(n_45),
.B(n_31),
.Y(n_57)
);

INVx3_ASAP7_75t_L g46 ( 
.A(n_41),
.Y(n_46)
);

BUFx12f_ASAP7_75t_L g59 ( 
.A(n_46),
.Y(n_59)
);

BUFx3_ASAP7_75t_L g47 ( 
.A(n_32),
.Y(n_47)
);

INVx5_ASAP7_75t_L g51 ( 
.A(n_47),
.Y(n_51)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_36),
.Y(n_48)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_48),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g49 ( 
.A(n_37),
.B(n_0),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_L g60 ( 
.A(n_49),
.B(n_38),
.Y(n_60)
);

INVx2_ASAP7_75t_L g50 ( 
.A(n_43),
.Y(n_50)
);

INVx2_ASAP7_75t_L g53 ( 
.A(n_50),
.Y(n_53)
);

INVx5_ASAP7_75t_L g52 ( 
.A(n_47),
.Y(n_52)
);

INVx4_ASAP7_75t_L g64 ( 
.A(n_52),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_SL g55 ( 
.A(n_46),
.B(n_31),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_55),
.B(n_56),
.Y(n_61)
);

AOI21xp5_ASAP7_75t_L g56 ( 
.A1(n_45),
.A2(n_32),
.B(n_43),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_57),
.B(n_60),
.Y(n_72)
);

AOI22xp5_ASAP7_75t_L g62 ( 
.A1(n_53),
.A2(n_39),
.B1(n_35),
.B2(n_34),
.Y(n_62)
);

OAI22xp5_ASAP7_75t_L g76 ( 
.A1(n_62),
.A2(n_67),
.B1(n_42),
.B2(n_15),
.Y(n_76)
);

INVx2_ASAP7_75t_L g63 ( 
.A(n_58),
.Y(n_63)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_63),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_L g65 ( 
.A(n_54),
.B(n_36),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_L g84 ( 
.A(n_65),
.B(n_16),
.Y(n_84)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_54),
.Y(n_66)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_66),
.Y(n_83)
);

AOI22xp5_ASAP7_75t_L g67 ( 
.A1(n_51),
.A2(n_39),
.B1(n_35),
.B2(n_34),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_L g68 ( 
.A(n_59),
.B(n_40),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_L g75 ( 
.A(n_68),
.B(n_42),
.Y(n_75)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_51),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_69),
.B(n_71),
.Y(n_79)
);

CKINVDCx20_ASAP7_75t_R g70 ( 
.A(n_52),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_SL g77 ( 
.A(n_70),
.B(n_64),
.Y(n_77)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_59),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_L g73 ( 
.A(n_61),
.B(n_59),
.Y(n_73)
);

XNOR2xp5_ASAP7_75t_L g92 ( 
.A(n_73),
.B(n_82),
.Y(n_92)
);

OR2x2_ASAP7_75t_L g74 ( 
.A(n_63),
.B(n_33),
.Y(n_74)
);

CKINVDCx14_ASAP7_75t_R g90 ( 
.A(n_74),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_75),
.B(n_77),
.Y(n_86)
);

AOI22xp5_ASAP7_75t_L g85 ( 
.A1(n_76),
.A2(n_67),
.B1(n_3),
.B2(n_4),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_72),
.B(n_0),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_SL g97 ( 
.A(n_80),
.B(n_81),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_64),
.B(n_1),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_62),
.B(n_2),
.Y(n_82)
);

MAJIxp5_ASAP7_75t_L g87 ( 
.A(n_84),
.B(n_18),
.C(n_29),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_85),
.B(n_87),
.Y(n_99)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_83),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_SL g98 ( 
.A(n_88),
.B(n_89),
.Y(n_98)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_79),
.Y(n_89)
);

MAJIxp5_ASAP7_75t_L g91 ( 
.A(n_73),
.B(n_14),
.C(n_28),
.Y(n_91)
);

MAJIxp5_ASAP7_75t_L g101 ( 
.A(n_91),
.B(n_96),
.C(n_20),
.Y(n_101)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_78),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_SL g104 ( 
.A(n_93),
.B(n_94),
.Y(n_104)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_74),
.Y(n_94)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_83),
.Y(n_95)
);

OAI21xp33_ASAP7_75t_L g100 ( 
.A1(n_95),
.A2(n_2),
.B(n_3),
.Y(n_100)
);

MAJIxp5_ASAP7_75t_L g96 ( 
.A(n_73),
.B(n_11),
.C(n_27),
.Y(n_96)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_100),
.Y(n_105)
);

MAJIxp5_ASAP7_75t_L g106 ( 
.A(n_101),
.B(n_102),
.C(n_103),
.Y(n_106)
);

A2O1A1O1Ixp25_ASAP7_75t_L g102 ( 
.A1(n_86),
.A2(n_9),
.B(n_24),
.C(n_23),
.D(n_21),
.Y(n_102)
);

MAJIxp5_ASAP7_75t_L g103 ( 
.A(n_86),
.B(n_92),
.C(n_90),
.Y(n_103)
);

MAJIxp5_ASAP7_75t_L g107 ( 
.A(n_98),
.B(n_90),
.C(n_97),
.Y(n_107)
);

OAI321xp33_ASAP7_75t_L g108 ( 
.A1(n_107),
.A2(n_98),
.A3(n_104),
.B1(n_99),
.B2(n_7),
.C(n_4),
.Y(n_108)
);

OAI21xp5_ASAP7_75t_SL g109 ( 
.A1(n_108),
.A2(n_105),
.B(n_6),
.Y(n_109)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_109),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_SL g111 ( 
.A(n_110),
.B(n_106),
.Y(n_111)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_111),
.Y(n_112)
);

CKINVDCx20_ASAP7_75t_R g113 ( 
.A(n_112),
.Y(n_113)
);

XOR2xp5_ASAP7_75t_L g114 ( 
.A(n_113),
.B(n_5),
.Y(n_114)
);


endmodule