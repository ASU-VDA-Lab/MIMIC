module fake_jpeg_2285_n_657 (n_13, n_1, n_10, n_6, n_14, n_19, n_18, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_657);

input n_13;
input n_1;
input n_10;
input n_6;
input n_14;
input n_19;
input n_18;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_657;

wire n_529;
wire n_595;
wire n_390;
wire n_552;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_252;
wire n_525;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_586;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_620;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_611;
wire n_44;
wire n_355;
wire n_519;
wire n_276;
wire n_143;
wire n_431;
wire n_102;
wire n_549;
wire n_196;
wire n_66;
wire n_374;
wire n_566;
wire n_142;
wire n_417;
wire n_362;
wire n_470;
wire n_597;
wire n_172;
wire n_547;
wire n_345;
wire n_591;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_513;
wire n_283;
wire n_107;
wire n_490;
wire n_635;
wire n_517;
wire n_629;
wire n_415;
wire n_479;
wire n_543;
wire n_357;
wire n_89;
wire n_131;
wire n_607;
wire n_294;
wire n_230;
wire n_643;
wire n_170;
wire n_602;
wire n_313;
wire n_542;
wire n_574;
wire n_264;
wire n_647;
wire n_437;
wire n_93;
wire n_227;
wire n_559;
wire n_641;
wire n_48;
wire n_465;
wire n_638;
wire n_200;
wire n_582;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_623;
wire n_579;
wire n_416;
wire n_221;
wire n_256;
wire n_454;
wire n_540;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_637;
wire n_370;
wire n_410;
wire n_571;
wire n_82;
wire n_155;
wire n_508;
wire n_309;
wire n_624;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_606;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_569;
wire n_596;
wire n_400;
wire n_646;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_544;
wire n_31;
wire n_277;
wire n_255;
wire n_605;
wire n_601;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_393;
wire n_349;
wire n_234;
wire n_530;
wire n_634;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_557;
wire n_408;
wire n_80;
wire n_562;
wire n_204;
wire n_639;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_645;
wire n_298;
wire n_106;
wire n_545;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_584;
wire n_254;
wire n_608;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_622;
wire n_463;
wire n_92;
wire n_332;
wire n_640;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_653;
wire n_474;
wire n_539;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_626;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_575;
wire n_268;
wire n_404;
wire n_91;
wire n_511;
wire n_486;
wire n_305;
wire n_161;
wire n_441;
wire n_555;
wire n_342;
wire n_642;
wire n_101;
wire n_226;
wire n_509;
wire n_644;
wire n_149;
wire n_87;
wire n_46;
wire n_578;
wire n_656;
wire n_589;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_614;
wire n_97;
wire n_649;
wire n_573;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_610;
wire n_174;
wire n_198;
wire n_422;
wire n_560;
wire n_190;
wire n_510;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_536;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_537;
wire n_110;
wire n_594;
wire n_590;
wire n_531;
wire n_76;
wire n_278;
wire n_343;
wire n_577;
wire n_26;
wire n_88;
wire n_397;
wire n_592;
wire n_363;
wire n_570;
wire n_238;
wire n_598;
wire n_615;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_554;
wire n_301;
wire n_609;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_648;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_523;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_533;
wire n_612;
wire n_296;
wire n_384;
wire n_588;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_585;
wire n_491;
wire n_24;
wire n_526;
wire n_467;
wire n_269;
wire n_572;
wire n_546;
wire n_287;
wire n_219;
wire n_452;
wire n_631;
wire n_433;
wire n_636;
wire n_77;
wire n_473;
wire n_45;
wire n_520;
wire n_476;
wire n_337;
wire n_317;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_344;
wire n_328;
wire n_650;
wire n_218;
wire n_63;
wire n_652;
wire n_599;
wire n_239;
wire n_243;
wire n_481;
wire n_628;
wire n_619;
wire n_348;
wire n_587;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_583;
wire n_522;
wire n_333;
wire n_518;
wire n_132;
wire n_133;
wire n_419;
wire n_378;
wire n_565;
wire n_302;
wire n_216;
wire n_528;
wire n_184;
wire n_655;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_260;
wire n_199;
wire n_550;
wire n_413;
wire n_275;
wire n_494;
wire n_604;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_551;
wire n_36;
wire n_62;
wire n_600;
wire n_492;
wire n_603;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_567;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_515;
wire n_347;
wire n_521;
wire n_424;
wire n_55;
wire n_358;
wire n_312;
wire n_47;
wire n_538;
wire n_625;
wire n_147;
wire n_449;
wire n_627;
wire n_98;
wire n_251;
wire n_534;
wire n_472;
wire n_279;
wire n_593;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_618;
wire n_356;
wire n_119;
wire n_484;
wire n_568;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_576;
wire n_469;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_553;
wire n_257;
wire n_61;
wire n_173;
wire n_561;
wire n_244;
wire n_232;
wire n_527;
wire n_482;
wire n_58;
wire n_41;
wire n_613;
wire n_630;
wire n_266;
wire n_548;
wire n_72;
wire n_512;
wire n_654;
wire n_445;
wire n_443;
wire n_617;
wire n_215;
wire n_212;
wire n_516;
wire n_183;
wire n_409;
wire n_532;
wire n_249;
wire n_412;
wire n_581;
wire n_217;
wire n_471;
wire n_580;
wire n_541;
wire n_53;
wire n_372;
wire n_558;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_535;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_556;
wire n_524;
wire n_402;
wire n_563;
wire n_504;
wire n_438;
wire n_475;
wire n_247;
wire n_157;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_633;
wire n_112;
wire n_632;
wire n_616;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_514;
wire n_651;
wire n_564;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_621;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

BUFx12f_ASAP7_75t_L g20 ( 
.A(n_13),
.Y(n_20)
);

BUFx12_ASAP7_75t_L g21 ( 
.A(n_14),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_0),
.Y(n_22)
);

BUFx12f_ASAP7_75t_L g23 ( 
.A(n_15),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_4),
.Y(n_24)
);

INVx2_ASAP7_75t_L g25 ( 
.A(n_19),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_3),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_0),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_8),
.Y(n_28)
);

BUFx3_ASAP7_75t_L g29 ( 
.A(n_18),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_7),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_5),
.Y(n_31)
);

BUFx16f_ASAP7_75t_L g32 ( 
.A(n_8),
.Y(n_32)
);

INVx2_ASAP7_75t_L g33 ( 
.A(n_6),
.Y(n_33)
);

BUFx4f_ASAP7_75t_L g34 ( 
.A(n_1),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_15),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_15),
.Y(n_36)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_19),
.Y(n_37)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_10),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_13),
.Y(n_39)
);

BUFx12f_ASAP7_75t_L g40 ( 
.A(n_4),
.Y(n_40)
);

INVx2_ASAP7_75t_L g41 ( 
.A(n_6),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_1),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_6),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_10),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_6),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_15),
.Y(n_46)
);

BUFx12_ASAP7_75t_L g47 ( 
.A(n_2),
.Y(n_47)
);

INVx1_ASAP7_75t_SL g48 ( 
.A(n_8),
.Y(n_48)
);

INVx1_ASAP7_75t_SL g49 ( 
.A(n_9),
.Y(n_49)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_16),
.Y(n_50)
);

INVxp67_ASAP7_75t_L g51 ( 
.A(n_16),
.Y(n_51)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_11),
.Y(n_52)
);

INVx3_ASAP7_75t_L g53 ( 
.A(n_18),
.Y(n_53)
);

INVx2_ASAP7_75t_L g54 ( 
.A(n_7),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_19),
.Y(n_55)
);

CKINVDCx20_ASAP7_75t_R g56 ( 
.A(n_16),
.Y(n_56)
);

BUFx8_ASAP7_75t_L g57 ( 
.A(n_2),
.Y(n_57)
);

CKINVDCx20_ASAP7_75t_R g58 ( 
.A(n_18),
.Y(n_58)
);

INVx6_ASAP7_75t_SL g59 ( 
.A(n_32),
.Y(n_59)
);

CKINVDCx6p67_ASAP7_75t_R g203 ( 
.A(n_59),
.Y(n_203)
);

INVx3_ASAP7_75t_L g60 ( 
.A(n_32),
.Y(n_60)
);

INVx2_ASAP7_75t_SL g181 ( 
.A(n_60),
.Y(n_181)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_25),
.Y(n_61)
);

INVx2_ASAP7_75t_L g143 ( 
.A(n_61),
.Y(n_143)
);

INVx8_ASAP7_75t_L g62 ( 
.A(n_40),
.Y(n_62)
);

INVx5_ASAP7_75t_L g144 ( 
.A(n_62),
.Y(n_144)
);

CKINVDCx20_ASAP7_75t_R g63 ( 
.A(n_32),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g164 ( 
.A(n_63),
.B(n_70),
.Y(n_164)
);

BUFx3_ASAP7_75t_L g64 ( 
.A(n_29),
.Y(n_64)
);

BUFx3_ASAP7_75t_L g201 ( 
.A(n_64),
.Y(n_201)
);

INVx2_ASAP7_75t_L g65 ( 
.A(n_25),
.Y(n_65)
);

INVx2_ASAP7_75t_L g151 ( 
.A(n_65),
.Y(n_151)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_30),
.Y(n_66)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_66),
.Y(n_157)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_30),
.Y(n_67)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_67),
.Y(n_183)
);

INVx2_ASAP7_75t_L g68 ( 
.A(n_33),
.Y(n_68)
);

INVx2_ASAP7_75t_L g158 ( 
.A(n_68),
.Y(n_158)
);

INVx4_ASAP7_75t_L g69 ( 
.A(n_32),
.Y(n_69)
);

INVx3_ASAP7_75t_L g140 ( 
.A(n_69),
.Y(n_140)
);

CKINVDCx20_ASAP7_75t_R g70 ( 
.A(n_51),
.Y(n_70)
);

BUFx6f_ASAP7_75t_L g71 ( 
.A(n_45),
.Y(n_71)
);

BUFx6f_ASAP7_75t_L g132 ( 
.A(n_71),
.Y(n_132)
);

BUFx12f_ASAP7_75t_L g72 ( 
.A(n_57),
.Y(n_72)
);

BUFx10_ASAP7_75t_L g197 ( 
.A(n_72),
.Y(n_197)
);

CKINVDCx20_ASAP7_75t_R g73 ( 
.A(n_45),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g166 ( 
.A(n_73),
.B(n_75),
.Y(n_166)
);

INVx4_ASAP7_75t_L g74 ( 
.A(n_40),
.Y(n_74)
);

INVx3_ASAP7_75t_L g150 ( 
.A(n_74),
.Y(n_150)
);

INVx6_ASAP7_75t_SL g75 ( 
.A(n_57),
.Y(n_75)
);

BUFx16f_ASAP7_75t_L g76 ( 
.A(n_57),
.Y(n_76)
);

BUFx3_ASAP7_75t_L g215 ( 
.A(n_76),
.Y(n_215)
);

BUFx6f_ASAP7_75t_L g77 ( 
.A(n_45),
.Y(n_77)
);

BUFx6f_ASAP7_75t_L g173 ( 
.A(n_77),
.Y(n_173)
);

INVx2_ASAP7_75t_L g78 ( 
.A(n_33),
.Y(n_78)
);

INVx2_ASAP7_75t_L g165 ( 
.A(n_78),
.Y(n_165)
);

BUFx8_ASAP7_75t_L g79 ( 
.A(n_57),
.Y(n_79)
);

BUFx2_ASAP7_75t_L g141 ( 
.A(n_79),
.Y(n_141)
);

BUFx6f_ASAP7_75t_L g80 ( 
.A(n_45),
.Y(n_80)
);

BUFx6f_ASAP7_75t_L g199 ( 
.A(n_80),
.Y(n_199)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_36),
.B(n_10),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g139 ( 
.A(n_81),
.B(n_83),
.Y(n_139)
);

BUFx6f_ASAP7_75t_L g82 ( 
.A(n_46),
.Y(n_82)
);

BUFx6f_ASAP7_75t_L g212 ( 
.A(n_82),
.Y(n_212)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_36),
.B(n_10),
.Y(n_83)
);

INVx2_ASAP7_75t_L g84 ( 
.A(n_41),
.Y(n_84)
);

INVx2_ASAP7_75t_L g191 ( 
.A(n_84),
.Y(n_191)
);

INVx2_ASAP7_75t_L g85 ( 
.A(n_41),
.Y(n_85)
);

INVx2_ASAP7_75t_L g198 ( 
.A(n_85),
.Y(n_198)
);

BUFx6f_ASAP7_75t_L g86 ( 
.A(n_46),
.Y(n_86)
);

BUFx6f_ASAP7_75t_L g217 ( 
.A(n_86),
.Y(n_217)
);

INVx3_ASAP7_75t_L g87 ( 
.A(n_40),
.Y(n_87)
);

INVx3_ASAP7_75t_L g188 ( 
.A(n_87),
.Y(n_188)
);

CKINVDCx20_ASAP7_75t_R g88 ( 
.A(n_46),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g170 ( 
.A(n_88),
.B(n_100),
.Y(n_170)
);

BUFx6f_ASAP7_75t_L g89 ( 
.A(n_46),
.Y(n_89)
);

BUFx6f_ASAP7_75t_L g227 ( 
.A(n_89),
.Y(n_227)
);

INVx2_ASAP7_75t_L g90 ( 
.A(n_54),
.Y(n_90)
);

INVx2_ASAP7_75t_L g207 ( 
.A(n_90),
.Y(n_207)
);

BUFx4f_ASAP7_75t_SL g91 ( 
.A(n_57),
.Y(n_91)
);

BUFx3_ASAP7_75t_L g218 ( 
.A(n_91),
.Y(n_218)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_37),
.Y(n_92)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_92),
.Y(n_185)
);

AOI22xp33_ASAP7_75t_SL g93 ( 
.A1(n_34),
.A2(n_9),
.B1(n_18),
.B2(n_17),
.Y(n_93)
);

OAI22xp5_ASAP7_75t_L g149 ( 
.A1(n_93),
.A2(n_49),
.B1(n_26),
.B2(n_42),
.Y(n_149)
);

INVx2_ASAP7_75t_L g94 ( 
.A(n_54),
.Y(n_94)
);

INVx2_ASAP7_75t_L g160 ( 
.A(n_94),
.Y(n_160)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_37),
.Y(n_95)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_95),
.Y(n_186)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_38),
.B(n_9),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g148 ( 
.A(n_96),
.B(n_115),
.Y(n_148)
);

NAND2xp33_ASAP7_75t_SL g97 ( 
.A(n_48),
.B(n_0),
.Y(n_97)
);

HAxp5_ASAP7_75t_SL g153 ( 
.A(n_97),
.B(n_0),
.CON(n_153),
.SN(n_153)
);

INVx2_ASAP7_75t_L g98 ( 
.A(n_34),
.Y(n_98)
);

INVx2_ASAP7_75t_L g205 ( 
.A(n_98),
.Y(n_205)
);

INVx3_ASAP7_75t_L g99 ( 
.A(n_40),
.Y(n_99)
);

INVx3_ASAP7_75t_L g228 ( 
.A(n_99),
.Y(n_228)
);

CKINVDCx20_ASAP7_75t_R g100 ( 
.A(n_35),
.Y(n_100)
);

INVx2_ASAP7_75t_L g101 ( 
.A(n_34),
.Y(n_101)
);

INVx2_ASAP7_75t_L g208 ( 
.A(n_101),
.Y(n_208)
);

INVx13_ASAP7_75t_L g102 ( 
.A(n_48),
.Y(n_102)
);

BUFx2_ASAP7_75t_L g163 ( 
.A(n_102),
.Y(n_163)
);

CKINVDCx20_ASAP7_75t_R g103 ( 
.A(n_35),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g175 ( 
.A(n_103),
.B(n_114),
.Y(n_175)
);

BUFx6f_ASAP7_75t_L g104 ( 
.A(n_35),
.Y(n_104)
);

INVx6_ASAP7_75t_L g136 ( 
.A(n_104),
.Y(n_136)
);

BUFx3_ASAP7_75t_L g105 ( 
.A(n_29),
.Y(n_105)
);

BUFx2_ASAP7_75t_L g194 ( 
.A(n_105),
.Y(n_194)
);

INVx2_ASAP7_75t_L g106 ( 
.A(n_34),
.Y(n_106)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_106),
.Y(n_190)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_38),
.Y(n_107)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_107),
.Y(n_193)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_50),
.Y(n_108)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_108),
.Y(n_219)
);

INVx3_ASAP7_75t_L g109 ( 
.A(n_40),
.Y(n_109)
);

INVx4_ASAP7_75t_L g137 ( 
.A(n_109),
.Y(n_137)
);

BUFx6f_ASAP7_75t_L g110 ( 
.A(n_43),
.Y(n_110)
);

INVx6_ASAP7_75t_L g154 ( 
.A(n_110),
.Y(n_154)
);

BUFx6f_ASAP7_75t_L g111 ( 
.A(n_43),
.Y(n_111)
);

INVx6_ASAP7_75t_L g172 ( 
.A(n_111),
.Y(n_172)
);

INVx3_ASAP7_75t_L g112 ( 
.A(n_29),
.Y(n_112)
);

INVx4_ASAP7_75t_L g161 ( 
.A(n_112),
.Y(n_161)
);

INVx2_ASAP7_75t_SL g113 ( 
.A(n_20),
.Y(n_113)
);

INVx4_ASAP7_75t_L g168 ( 
.A(n_113),
.Y(n_168)
);

CKINVDCx20_ASAP7_75t_R g114 ( 
.A(n_43),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_L g115 ( 
.A(n_50),
.B(n_9),
.Y(n_115)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_24),
.Y(n_116)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_116),
.Y(n_225)
);

INVx3_ASAP7_75t_L g117 ( 
.A(n_53),
.Y(n_117)
);

INVx4_ASAP7_75t_L g171 ( 
.A(n_117),
.Y(n_171)
);

NOR2xp33_ASAP7_75t_L g118 ( 
.A(n_28),
.B(n_58),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_L g156 ( 
.A(n_118),
.B(n_56),
.Y(n_156)
);

BUFx6f_ASAP7_75t_L g119 ( 
.A(n_44),
.Y(n_119)
);

INVx6_ASAP7_75t_L g176 ( 
.A(n_119),
.Y(n_176)
);

INVx3_ASAP7_75t_L g120 ( 
.A(n_53),
.Y(n_120)
);

INVx4_ASAP7_75t_L g178 ( 
.A(n_120),
.Y(n_178)
);

CKINVDCx20_ASAP7_75t_R g121 ( 
.A(n_44),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_L g177 ( 
.A(n_121),
.B(n_122),
.Y(n_177)
);

INVx3_ASAP7_75t_SL g122 ( 
.A(n_53),
.Y(n_122)
);

AND2x2_ASAP7_75t_L g134 ( 
.A(n_122),
.B(n_131),
.Y(n_134)
);

BUFx12f_ASAP7_75t_L g123 ( 
.A(n_21),
.Y(n_123)
);

INVx8_ASAP7_75t_L g133 ( 
.A(n_123),
.Y(n_133)
);

BUFx6f_ASAP7_75t_L g124 ( 
.A(n_44),
.Y(n_124)
);

INVx8_ASAP7_75t_L g142 ( 
.A(n_124),
.Y(n_142)
);

BUFx6f_ASAP7_75t_L g125 ( 
.A(n_55),
.Y(n_125)
);

INVx8_ASAP7_75t_L g174 ( 
.A(n_125),
.Y(n_174)
);

INVx3_ASAP7_75t_L g126 ( 
.A(n_20),
.Y(n_126)
);

INVx4_ASAP7_75t_L g222 ( 
.A(n_126),
.Y(n_222)
);

BUFx6f_ASAP7_75t_L g127 ( 
.A(n_55),
.Y(n_127)
);

INVx8_ASAP7_75t_L g195 ( 
.A(n_127),
.Y(n_195)
);

BUFx6f_ASAP7_75t_L g128 ( 
.A(n_55),
.Y(n_128)
);

INVx8_ASAP7_75t_L g216 ( 
.A(n_128),
.Y(n_216)
);

BUFx12f_ASAP7_75t_L g129 ( 
.A(n_21),
.Y(n_129)
);

INVx5_ASAP7_75t_L g189 ( 
.A(n_129),
.Y(n_189)
);

BUFx6f_ASAP7_75t_L g130 ( 
.A(n_20),
.Y(n_130)
);

INVx5_ASAP7_75t_L g210 ( 
.A(n_130),
.Y(n_210)
);

INVx4_ASAP7_75t_L g131 ( 
.A(n_20),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_SL g135 ( 
.A(n_117),
.B(n_58),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_SL g246 ( 
.A(n_135),
.B(n_145),
.Y(n_246)
);

AOI22xp33_ASAP7_75t_L g138 ( 
.A1(n_104),
.A2(n_22),
.B1(n_26),
.B2(n_27),
.Y(n_138)
);

OAI22xp5_ASAP7_75t_L g290 ( 
.A1(n_138),
.A2(n_159),
.B1(n_167),
.B2(n_179),
.Y(n_290)
);

CKINVDCx20_ASAP7_75t_R g145 ( 
.A(n_76),
.Y(n_145)
);

AOI22xp33_ASAP7_75t_SL g146 ( 
.A1(n_79),
.A2(n_49),
.B1(n_48),
.B2(n_20),
.Y(n_146)
);

OA22x2_ASAP7_75t_L g272 ( 
.A1(n_146),
.A2(n_147),
.B1(n_152),
.B2(n_180),
.Y(n_272)
);

AOI22xp33_ASAP7_75t_SL g147 ( 
.A1(n_79),
.A2(n_49),
.B1(n_23),
.B2(n_22),
.Y(n_147)
);

AOI22xp5_ASAP7_75t_L g241 ( 
.A1(n_149),
.A2(n_202),
.B1(n_77),
.B2(n_89),
.Y(n_241)
);

AOI22xp33_ASAP7_75t_SL g152 ( 
.A1(n_72),
.A2(n_23),
.B1(n_27),
.B2(n_42),
.Y(n_152)
);

OAI21xp33_ASAP7_75t_L g288 ( 
.A1(n_153),
.A2(n_224),
.B(n_180),
.Y(n_288)
);

NAND2xp5_ASAP7_75t_SL g155 ( 
.A(n_120),
.B(n_56),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_SL g249 ( 
.A(n_155),
.B(n_156),
.Y(n_249)
);

AOI22xp5_ASAP7_75t_L g159 ( 
.A1(n_110),
.A2(n_39),
.B1(n_31),
.B2(n_28),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_L g162 ( 
.A(n_87),
.B(n_52),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_L g243 ( 
.A(n_162),
.B(n_196),
.Y(n_243)
);

OAI22xp5_ASAP7_75t_L g167 ( 
.A1(n_111),
.A2(n_52),
.B1(n_39),
.B2(n_31),
.Y(n_167)
);

CKINVDCx20_ASAP7_75t_R g169 ( 
.A(n_76),
.Y(n_169)
);

NOR2xp33_ASAP7_75t_L g237 ( 
.A(n_169),
.B(n_184),
.Y(n_237)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_177),
.Y(n_250)
);

AOI22xp33_ASAP7_75t_L g179 ( 
.A1(n_119),
.A2(n_24),
.B1(n_23),
.B2(n_47),
.Y(n_179)
);

AOI22xp33_ASAP7_75t_SL g180 ( 
.A1(n_72),
.A2(n_23),
.B1(n_47),
.B2(n_21),
.Y(n_180)
);

AOI22xp33_ASAP7_75t_SL g182 ( 
.A1(n_113),
.A2(n_23),
.B1(n_47),
.B2(n_21),
.Y(n_182)
);

OAI22xp33_ASAP7_75t_L g254 ( 
.A1(n_182),
.A2(n_204),
.B1(n_221),
.B2(n_224),
.Y(n_254)
);

AND2x2_ASAP7_75t_L g184 ( 
.A(n_69),
.B(n_11),
.Y(n_184)
);

NOR2xp33_ASAP7_75t_SL g187 ( 
.A(n_60),
.B(n_11),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_SL g238 ( 
.A(n_187),
.B(n_192),
.Y(n_238)
);

NOR2xp33_ASAP7_75t_SL g192 ( 
.A(n_74),
.B(n_11),
.Y(n_192)
);

NOR2xp33_ASAP7_75t_L g196 ( 
.A(n_91),
.B(n_12),
.Y(n_196)
);

NOR2xp33_ASAP7_75t_L g200 ( 
.A(n_91),
.B(n_12),
.Y(n_200)
);

NAND2xp5_ASAP7_75t_L g245 ( 
.A(n_200),
.B(n_211),
.Y(n_245)
);

OAI22xp5_ASAP7_75t_SL g202 ( 
.A1(n_124),
.A2(n_21),
.B1(n_47),
.B2(n_12),
.Y(n_202)
);

AOI22xp33_ASAP7_75t_SL g204 ( 
.A1(n_112),
.A2(n_47),
.B1(n_8),
.B2(n_12),
.Y(n_204)
);

AND2x2_ASAP7_75t_L g206 ( 
.A(n_99),
.B(n_109),
.Y(n_206)
);

NOR2xp33_ASAP7_75t_L g267 ( 
.A(n_206),
.B(n_4),
.Y(n_267)
);

CKINVDCx14_ASAP7_75t_SL g209 ( 
.A(n_102),
.Y(n_209)
);

INVx11_ASAP7_75t_L g275 ( 
.A(n_209),
.Y(n_275)
);

NOR2xp33_ASAP7_75t_L g211 ( 
.A(n_123),
.B(n_7),
.Y(n_211)
);

NAND2xp5_ASAP7_75t_L g213 ( 
.A(n_126),
.B(n_7),
.Y(n_213)
);

NAND2xp5_ASAP7_75t_L g253 ( 
.A(n_213),
.B(n_214),
.Y(n_253)
);

NOR2xp33_ASAP7_75t_L g214 ( 
.A(n_123),
.B(n_19),
.Y(n_214)
);

NAND2xp5_ASAP7_75t_L g220 ( 
.A(n_97),
.B(n_131),
.Y(n_220)
);

NAND2xp5_ASAP7_75t_L g269 ( 
.A(n_220),
.B(n_226),
.Y(n_269)
);

AOI22xp33_ASAP7_75t_SL g221 ( 
.A1(n_64),
.A2(n_5),
.B1(n_16),
.B2(n_14),
.Y(n_221)
);

AOI22xp5_ASAP7_75t_SL g223 ( 
.A1(n_105),
.A2(n_17),
.B1(n_14),
.B2(n_13),
.Y(n_223)
);

OAI22xp33_ASAP7_75t_SL g240 ( 
.A1(n_223),
.A2(n_125),
.B1(n_128),
.B2(n_127),
.Y(n_240)
);

AOI22xp33_ASAP7_75t_SL g224 ( 
.A1(n_62),
.A2(n_17),
.B1(n_14),
.B2(n_13),
.Y(n_224)
);

NOR2xp33_ASAP7_75t_L g226 ( 
.A(n_129),
.B(n_17),
.Y(n_226)
);

INVx2_ASAP7_75t_L g229 ( 
.A(n_205),
.Y(n_229)
);

INVx2_ASAP7_75t_L g322 ( 
.A(n_229),
.Y(n_322)
);

INVx4_ASAP7_75t_SL g230 ( 
.A(n_203),
.Y(n_230)
);

NOR2xp33_ASAP7_75t_L g325 ( 
.A(n_230),
.B(n_262),
.Y(n_325)
);

INVx2_ASAP7_75t_L g231 ( 
.A(n_205),
.Y(n_231)
);

INVx2_ASAP7_75t_L g343 ( 
.A(n_231),
.Y(n_343)
);

INVx5_ASAP7_75t_L g232 ( 
.A(n_218),
.Y(n_232)
);

INVx4_ASAP7_75t_L g334 ( 
.A(n_232),
.Y(n_334)
);

BUFx6f_ASAP7_75t_L g233 ( 
.A(n_132),
.Y(n_233)
);

INVx2_ASAP7_75t_L g371 ( 
.A(n_233),
.Y(n_371)
);

NAND2xp5_ASAP7_75t_L g234 ( 
.A(n_139),
.B(n_0),
.Y(n_234)
);

NAND2xp5_ASAP7_75t_L g314 ( 
.A(n_234),
.B(n_239),
.Y(n_314)
);

BUFx3_ASAP7_75t_L g235 ( 
.A(n_215),
.Y(n_235)
);

HB1xp67_ASAP7_75t_L g329 ( 
.A(n_235),
.Y(n_329)
);

MAJIxp5_ASAP7_75t_L g236 ( 
.A(n_225),
.B(n_130),
.C(n_93),
.Y(n_236)
);

MAJIxp5_ASAP7_75t_L g370 ( 
.A(n_236),
.B(n_252),
.C(n_255),
.Y(n_370)
);

NAND2xp5_ASAP7_75t_L g239 ( 
.A(n_148),
.B(n_1),
.Y(n_239)
);

AOI22xp5_ASAP7_75t_L g317 ( 
.A1(n_240),
.A2(n_244),
.B1(n_285),
.B2(n_189),
.Y(n_317)
);

OA22x2_ASAP7_75t_L g367 ( 
.A1(n_241),
.A2(n_280),
.B1(n_266),
.B2(n_260),
.Y(n_367)
);

BUFx6f_ASAP7_75t_L g242 ( 
.A(n_132),
.Y(n_242)
);

INVxp67_ASAP7_75t_L g332 ( 
.A(n_242),
.Y(n_332)
);

OAI22xp33_ASAP7_75t_SL g244 ( 
.A1(n_159),
.A2(n_223),
.B1(n_175),
.B2(n_170),
.Y(n_244)
);

INVx2_ASAP7_75t_L g247 ( 
.A(n_208),
.Y(n_247)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_247),
.Y(n_312)
);

BUFx6f_ASAP7_75t_L g248 ( 
.A(n_173),
.Y(n_248)
);

INVxp67_ASAP7_75t_L g361 ( 
.A(n_248),
.Y(n_361)
);

HB1xp67_ASAP7_75t_L g251 ( 
.A(n_168),
.Y(n_251)
);

CKINVDCx16_ASAP7_75t_R g321 ( 
.A(n_251),
.Y(n_321)
);

AND2x2_ASAP7_75t_L g252 ( 
.A(n_134),
.B(n_129),
.Y(n_252)
);

AND2x2_ASAP7_75t_L g255 ( 
.A(n_134),
.B(n_1),
.Y(n_255)
);

AOI22xp5_ASAP7_75t_L g256 ( 
.A1(n_202),
.A2(n_86),
.B1(n_82),
.B2(n_80),
.Y(n_256)
);

OAI22xp5_ASAP7_75t_L g326 ( 
.A1(n_256),
.A2(n_260),
.B1(n_266),
.B2(n_280),
.Y(n_326)
);

AND2x2_ASAP7_75t_L g257 ( 
.A(n_206),
.B(n_1),
.Y(n_257)
);

XNOR2xp5_ASAP7_75t_L g340 ( 
.A(n_257),
.B(n_258),
.Y(n_340)
);

AND2x2_ASAP7_75t_L g258 ( 
.A(n_184),
.B(n_2),
.Y(n_258)
);

NAND2xp5_ASAP7_75t_SL g259 ( 
.A(n_157),
.B(n_71),
.Y(n_259)
);

NOR2xp33_ASAP7_75t_SL g333 ( 
.A(n_259),
.B(n_276),
.Y(n_333)
);

AOI22xp5_ASAP7_75t_L g260 ( 
.A1(n_160),
.A2(n_5),
.B1(n_3),
.B2(n_4),
.Y(n_260)
);

BUFx6f_ASAP7_75t_L g261 ( 
.A(n_173),
.Y(n_261)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_261),
.Y(n_320)
);

CKINVDCx16_ASAP7_75t_R g262 ( 
.A(n_203),
.Y(n_262)
);

NAND2xp5_ASAP7_75t_L g263 ( 
.A(n_183),
.B(n_2),
.Y(n_263)
);

NAND2xp5_ASAP7_75t_L g315 ( 
.A(n_263),
.B(n_268),
.Y(n_315)
);

CKINVDCx20_ASAP7_75t_R g264 ( 
.A(n_203),
.Y(n_264)
);

NAND3xp33_ASAP7_75t_L g360 ( 
.A(n_264),
.B(n_267),
.C(n_271),
.Y(n_360)
);

INVx3_ASAP7_75t_L g265 ( 
.A(n_215),
.Y(n_265)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_265),
.Y(n_323)
);

AOI22xp5_ASAP7_75t_L g266 ( 
.A1(n_160),
.A2(n_5),
.B1(n_3),
.B2(n_4),
.Y(n_266)
);

NAND2xp5_ASAP7_75t_L g268 ( 
.A(n_185),
.B(n_2),
.Y(n_268)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_186),
.Y(n_270)
);

NOR2xp33_ASAP7_75t_L g363 ( 
.A(n_270),
.B(n_279),
.Y(n_363)
);

CKINVDCx20_ASAP7_75t_R g271 ( 
.A(n_164),
.Y(n_271)
);

INVx2_ASAP7_75t_L g273 ( 
.A(n_208),
.Y(n_273)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_273),
.Y(n_336)
);

BUFx6f_ASAP7_75t_L g274 ( 
.A(n_199),
.Y(n_274)
);

INVx1_ASAP7_75t_L g342 ( 
.A(n_274),
.Y(n_342)
);

NAND2xp5_ASAP7_75t_L g276 ( 
.A(n_193),
.B(n_3),
.Y(n_276)
);

NOR2xp33_ASAP7_75t_L g277 ( 
.A(n_219),
.B(n_3),
.Y(n_277)
);

NOR2xp33_ASAP7_75t_L g331 ( 
.A(n_277),
.B(n_281),
.Y(n_331)
);

AND2x2_ASAP7_75t_L g278 ( 
.A(n_163),
.B(n_168),
.Y(n_278)
);

XNOR2xp5_ASAP7_75t_L g352 ( 
.A(n_278),
.B(n_287),
.Y(n_352)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_190),
.Y(n_279)
);

AOI22xp5_ASAP7_75t_L g280 ( 
.A1(n_143),
.A2(n_165),
.B1(n_207),
.B2(n_158),
.Y(n_280)
);

CKINVDCx16_ASAP7_75t_R g281 ( 
.A(n_163),
.Y(n_281)
);

CKINVDCx20_ASAP7_75t_R g282 ( 
.A(n_166),
.Y(n_282)
);

NOR2xp33_ASAP7_75t_L g356 ( 
.A(n_282),
.B(n_296),
.Y(n_356)
);

NAND2xp5_ASAP7_75t_L g283 ( 
.A(n_151),
.B(n_198),
.Y(n_283)
);

NAND2xp5_ASAP7_75t_L g337 ( 
.A(n_283),
.B(n_294),
.Y(n_337)
);

NAND2xp5_ASAP7_75t_SL g284 ( 
.A(n_191),
.B(n_181),
.Y(n_284)
);

NAND2xp5_ASAP7_75t_SL g328 ( 
.A(n_284),
.B(n_301),
.Y(n_328)
);

OAI22xp33_ASAP7_75t_SL g285 ( 
.A1(n_152),
.A2(n_147),
.B1(n_221),
.B2(n_146),
.Y(n_285)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_181),
.Y(n_286)
);

INVx1_ASAP7_75t_L g347 ( 
.A(n_286),
.Y(n_347)
);

AND2x2_ASAP7_75t_L g287 ( 
.A(n_171),
.B(n_178),
.Y(n_287)
);

OAI21xp5_ASAP7_75t_L g319 ( 
.A1(n_288),
.A2(n_133),
.B(n_216),
.Y(n_319)
);

INVx4_ASAP7_75t_L g289 ( 
.A(n_144),
.Y(n_289)
);

INVx1_ASAP7_75t_L g348 ( 
.A(n_289),
.Y(n_348)
);

A2O1A1Ixp33_ASAP7_75t_L g291 ( 
.A1(n_153),
.A2(n_182),
.B(n_197),
.C(n_218),
.Y(n_291)
);

A2O1A1Ixp33_ASAP7_75t_L g345 ( 
.A1(n_291),
.A2(n_305),
.B(n_236),
.C(n_306),
.Y(n_345)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_140),
.Y(n_292)
);

INVx1_ASAP7_75t_L g354 ( 
.A(n_292),
.Y(n_354)
);

INVx3_ASAP7_75t_L g293 ( 
.A(n_144),
.Y(n_293)
);

INVx1_ASAP7_75t_L g359 ( 
.A(n_293),
.Y(n_359)
);

NAND2xp5_ASAP7_75t_L g294 ( 
.A(n_228),
.B(n_188),
.Y(n_294)
);

INVx6_ASAP7_75t_L g295 ( 
.A(n_142),
.Y(n_295)
);

INVx1_ASAP7_75t_L g362 ( 
.A(n_295),
.Y(n_362)
);

NOR2xp33_ASAP7_75t_L g296 ( 
.A(n_140),
.B(n_228),
.Y(n_296)
);

INVx2_ASAP7_75t_L g297 ( 
.A(n_161),
.Y(n_297)
);

INVx1_ASAP7_75t_L g364 ( 
.A(n_297),
.Y(n_364)
);

BUFx6f_ASAP7_75t_L g298 ( 
.A(n_199),
.Y(n_298)
);

INVx1_ASAP7_75t_L g366 ( 
.A(n_298),
.Y(n_366)
);

NOR2xp33_ASAP7_75t_L g299 ( 
.A(n_188),
.B(n_150),
.Y(n_299)
);

NOR2xp33_ASAP7_75t_L g369 ( 
.A(n_299),
.B(n_302),
.Y(n_369)
);

NAND2xp5_ASAP7_75t_L g300 ( 
.A(n_150),
.B(n_137),
.Y(n_300)
);

NAND2xp5_ASAP7_75t_L g341 ( 
.A(n_300),
.B(n_308),
.Y(n_341)
);

NAND2xp5_ASAP7_75t_L g301 ( 
.A(n_137),
.B(n_222),
.Y(n_301)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_161),
.Y(n_302)
);

NOR2xp33_ASAP7_75t_L g303 ( 
.A(n_194),
.B(n_178),
.Y(n_303)
);

OR2x2_ASAP7_75t_L g318 ( 
.A(n_303),
.B(n_306),
.Y(n_318)
);

INVx3_ASAP7_75t_L g304 ( 
.A(n_222),
.Y(n_304)
);

CKINVDCx20_ASAP7_75t_R g316 ( 
.A(n_304),
.Y(n_316)
);

AOI32xp33_ASAP7_75t_L g305 ( 
.A1(n_171),
.A2(n_197),
.A3(n_204),
.B1(n_194),
.B2(n_141),
.Y(n_305)
);

NAND2xp33_ASAP7_75t_SL g306 ( 
.A(n_141),
.B(n_201),
.Y(n_306)
);

INVx6_ASAP7_75t_L g307 ( 
.A(n_142),
.Y(n_307)
);

CKINVDCx20_ASAP7_75t_R g324 ( 
.A(n_307),
.Y(n_324)
);

NAND2xp5_ASAP7_75t_L g308 ( 
.A(n_136),
.B(n_176),
.Y(n_308)
);

INVx3_ASAP7_75t_L g309 ( 
.A(n_210),
.Y(n_309)
);

CKINVDCx20_ASAP7_75t_R g349 ( 
.A(n_309),
.Y(n_349)
);

NAND2xp5_ASAP7_75t_L g310 ( 
.A(n_136),
.B(n_176),
.Y(n_310)
);

NAND2xp5_ASAP7_75t_L g346 ( 
.A(n_310),
.B(n_311),
.Y(n_346)
);

AOI22xp5_ASAP7_75t_L g311 ( 
.A1(n_227),
.A2(n_217),
.B1(n_212),
.B2(n_216),
.Y(n_311)
);

OAI22xp5_ASAP7_75t_SL g335 ( 
.A1(n_311),
.A2(n_154),
.B1(n_172),
.B2(n_174),
.Y(n_335)
);

AOI22xp33_ASAP7_75t_SL g313 ( 
.A1(n_290),
.A2(n_201),
.B1(n_189),
.B2(n_133),
.Y(n_313)
);

INVxp67_ASAP7_75t_L g378 ( 
.A(n_313),
.Y(n_378)
);

AND2x2_ASAP7_75t_L g416 ( 
.A(n_317),
.B(n_345),
.Y(n_416)
);

INVxp67_ASAP7_75t_L g383 ( 
.A(n_319),
.Y(n_383)
);

OAI22xp33_ASAP7_75t_SL g327 ( 
.A1(n_241),
.A2(n_227),
.B1(n_217),
.B2(n_212),
.Y(n_327)
);

AOI22xp5_ASAP7_75t_L g390 ( 
.A1(n_327),
.A2(n_335),
.B1(n_338),
.B2(n_339),
.Y(n_390)
);

AOI22xp5_ASAP7_75t_L g330 ( 
.A1(n_256),
.A2(n_174),
.B1(n_195),
.B2(n_210),
.Y(n_330)
);

OAI22xp5_ASAP7_75t_L g391 ( 
.A1(n_330),
.A2(n_355),
.B1(n_368),
.B2(n_293),
.Y(n_391)
);

OAI22xp5_ASAP7_75t_SL g338 ( 
.A1(n_269),
.A2(n_154),
.B1(n_172),
.B2(n_195),
.Y(n_338)
);

OAI22xp5_ASAP7_75t_SL g339 ( 
.A1(n_243),
.A2(n_263),
.B1(n_268),
.B2(n_308),
.Y(n_339)
);

OAI22xp5_ASAP7_75t_SL g344 ( 
.A1(n_310),
.A2(n_197),
.B1(n_253),
.B2(n_254),
.Y(n_344)
);

AOI22xp5_ASAP7_75t_L g406 ( 
.A1(n_344),
.A2(n_367),
.B1(n_338),
.B2(n_318),
.Y(n_406)
);

NAND2xp5_ASAP7_75t_L g380 ( 
.A(n_346),
.B(n_350),
.Y(n_380)
);

NAND2xp5_ASAP7_75t_L g350 ( 
.A(n_258),
.B(n_283),
.Y(n_350)
);

NAND2xp5_ASAP7_75t_L g351 ( 
.A(n_258),
.B(n_239),
.Y(n_351)
);

NAND2xp5_ASAP7_75t_L g387 ( 
.A(n_351),
.B(n_353),
.Y(n_387)
);

NAND2xp5_ASAP7_75t_L g353 ( 
.A(n_234),
.B(n_245),
.Y(n_353)
);

AOI22xp5_ASAP7_75t_L g355 ( 
.A1(n_288),
.A2(n_254),
.B1(n_291),
.B2(n_257),
.Y(n_355)
);

CKINVDCx20_ASAP7_75t_R g357 ( 
.A(n_278),
.Y(n_357)
);

NOR2xp33_ASAP7_75t_L g374 ( 
.A(n_357),
.B(n_372),
.Y(n_374)
);

NAND2xp5_ASAP7_75t_L g358 ( 
.A(n_294),
.B(n_257),
.Y(n_358)
);

NAND2xp5_ASAP7_75t_SL g384 ( 
.A(n_358),
.B(n_287),
.Y(n_384)
);

OR2x2_ASAP7_75t_L g365 ( 
.A(n_246),
.B(n_250),
.Y(n_365)
);

CKINVDCx16_ASAP7_75t_R g382 ( 
.A(n_365),
.Y(n_382)
);

AOI22xp5_ASAP7_75t_L g368 ( 
.A1(n_237),
.A2(n_255),
.B1(n_300),
.B2(n_272),
.Y(n_368)
);

CKINVDCx20_ASAP7_75t_R g372 ( 
.A(n_278),
.Y(n_372)
);

MAJIxp5_ASAP7_75t_L g373 ( 
.A(n_370),
.B(n_252),
.C(n_272),
.Y(n_373)
);

MAJIxp5_ASAP7_75t_L g426 ( 
.A(n_373),
.B(n_385),
.C(n_388),
.Y(n_426)
);

AOI21xp5_ASAP7_75t_L g375 ( 
.A1(n_319),
.A2(n_272),
.B(n_252),
.Y(n_375)
);

AOI21xp5_ASAP7_75t_L g456 ( 
.A1(n_375),
.A2(n_396),
.B(n_413),
.Y(n_456)
);

NOR2xp33_ASAP7_75t_L g376 ( 
.A(n_365),
.B(n_249),
.Y(n_376)
);

NOR2xp33_ASAP7_75t_SL g427 ( 
.A(n_376),
.B(n_377),
.Y(n_427)
);

NOR2xp33_ASAP7_75t_L g377 ( 
.A(n_365),
.B(n_238),
.Y(n_377)
);

OAI22xp5_ASAP7_75t_SL g379 ( 
.A1(n_368),
.A2(n_272),
.B1(n_255),
.B2(n_298),
.Y(n_379)
);

AOI22xp5_ASAP7_75t_L g421 ( 
.A1(n_379),
.A2(n_391),
.B1(n_398),
.B2(n_402),
.Y(n_421)
);

INVx4_ASAP7_75t_L g381 ( 
.A(n_371),
.Y(n_381)
);

INVx1_ASAP7_75t_L g422 ( 
.A(n_381),
.Y(n_422)
);

NAND2xp5_ASAP7_75t_SL g452 ( 
.A(n_384),
.B(n_321),
.Y(n_452)
);

XOR2xp5_ASAP7_75t_L g385 ( 
.A(n_370),
.B(n_287),
.Y(n_385)
);

OAI21xp5_ASAP7_75t_L g386 ( 
.A1(n_345),
.A2(n_265),
.B(n_297),
.Y(n_386)
);

OAI21xp5_ASAP7_75t_SL g429 ( 
.A1(n_386),
.A2(n_393),
.B(n_407),
.Y(n_429)
);

MAJIxp5_ASAP7_75t_L g388 ( 
.A(n_340),
.B(n_229),
.C(n_273),
.Y(n_388)
);

NOR2xp33_ASAP7_75t_L g389 ( 
.A(n_356),
.B(n_230),
.Y(n_389)
);

NOR2xp33_ASAP7_75t_SL g431 ( 
.A(n_389),
.B(n_397),
.Y(n_431)
);

OA21x2_ASAP7_75t_L g392 ( 
.A1(n_318),
.A2(n_304),
.B(n_289),
.Y(n_392)
);

NAND2xp5_ASAP7_75t_L g432 ( 
.A(n_392),
.B(n_403),
.Y(n_432)
);

OAI21xp5_ASAP7_75t_L g393 ( 
.A1(n_318),
.A2(n_235),
.B(n_231),
.Y(n_393)
);

INVx5_ASAP7_75t_L g394 ( 
.A(n_334),
.Y(n_394)
);

INVx1_ASAP7_75t_L g430 ( 
.A(n_394),
.Y(n_430)
);

BUFx3_ASAP7_75t_L g395 ( 
.A(n_334),
.Y(n_395)
);

INVx1_ASAP7_75t_L g434 ( 
.A(n_395),
.Y(n_434)
);

O2A1O1Ixp33_ASAP7_75t_L g396 ( 
.A1(n_326),
.A2(n_275),
.B(n_247),
.C(n_232),
.Y(n_396)
);

NAND2xp5_ASAP7_75t_SL g397 ( 
.A(n_315),
.B(n_307),
.Y(n_397)
);

OAI22xp5_ASAP7_75t_SL g398 ( 
.A1(n_355),
.A2(n_233),
.B1(n_242),
.B2(n_248),
.Y(n_398)
);

INVxp67_ASAP7_75t_L g399 ( 
.A(n_331),
.Y(n_399)
);

NOR2xp33_ASAP7_75t_L g439 ( 
.A(n_399),
.B(n_408),
.Y(n_439)
);

INVx1_ASAP7_75t_L g400 ( 
.A(n_347),
.Y(n_400)
);

INVx1_ASAP7_75t_L g442 ( 
.A(n_400),
.Y(n_442)
);

INVx1_ASAP7_75t_L g401 ( 
.A(n_347),
.Y(n_401)
);

INVx1_ASAP7_75t_L g445 ( 
.A(n_401),
.Y(n_445)
);

OAI22xp5_ASAP7_75t_SL g402 ( 
.A1(n_317),
.A2(n_261),
.B1(n_274),
.B2(n_295),
.Y(n_402)
);

NOR2xp33_ASAP7_75t_L g403 ( 
.A(n_333),
.B(n_309),
.Y(n_403)
);

INVx1_ASAP7_75t_L g404 ( 
.A(n_312),
.Y(n_404)
);

INVx1_ASAP7_75t_L g447 ( 
.A(n_404),
.Y(n_447)
);

OAI22xp5_ASAP7_75t_L g405 ( 
.A1(n_341),
.A2(n_275),
.B1(n_346),
.B2(n_326),
.Y(n_405)
);

AOI22xp5_ASAP7_75t_L g435 ( 
.A1(n_405),
.A2(n_406),
.B1(n_415),
.B2(n_359),
.Y(n_435)
);

OAI21xp5_ASAP7_75t_L g407 ( 
.A1(n_337),
.A2(n_328),
.B(n_341),
.Y(n_407)
);

FAx1_ASAP7_75t_SL g408 ( 
.A(n_339),
.B(n_344),
.CI(n_353),
.CON(n_408),
.SN(n_408)
);

NOR2xp33_ASAP7_75t_L g409 ( 
.A(n_333),
.B(n_369),
.Y(n_409)
);

NAND2xp5_ASAP7_75t_L g453 ( 
.A(n_409),
.B(n_343),
.Y(n_453)
);

INVx2_ASAP7_75t_L g410 ( 
.A(n_322),
.Y(n_410)
);

INVx1_ASAP7_75t_L g450 ( 
.A(n_410),
.Y(n_450)
);

XNOR2xp5_ASAP7_75t_L g411 ( 
.A(n_314),
.B(n_340),
.Y(n_411)
);

XNOR2xp5_ASAP7_75t_L g436 ( 
.A(n_411),
.B(n_354),
.Y(n_436)
);

MAJIxp5_ASAP7_75t_L g412 ( 
.A(n_358),
.B(n_350),
.C(n_337),
.Y(n_412)
);

MAJIxp5_ASAP7_75t_L g460 ( 
.A(n_412),
.B(n_417),
.C(n_419),
.Y(n_460)
);

AOI21xp5_ASAP7_75t_L g413 ( 
.A1(n_325),
.A2(n_372),
.B(n_357),
.Y(n_413)
);

INVx2_ASAP7_75t_L g414 ( 
.A(n_322),
.Y(n_414)
);

INVx1_ASAP7_75t_L g461 ( 
.A(n_414),
.Y(n_461)
);

OAI22xp5_ASAP7_75t_SL g415 ( 
.A1(n_315),
.A2(n_367),
.B1(n_328),
.B2(n_330),
.Y(n_415)
);

MAJIxp5_ASAP7_75t_L g417 ( 
.A(n_352),
.B(n_314),
.C(n_351),
.Y(n_417)
);

AOI22xp5_ASAP7_75t_L g418 ( 
.A1(n_367),
.A2(n_335),
.B1(n_352),
.B2(n_324),
.Y(n_418)
);

OAI22xp5_ASAP7_75t_L g424 ( 
.A1(n_418),
.A2(n_420),
.B1(n_367),
.B2(n_325),
.Y(n_424)
);

MAJIxp5_ASAP7_75t_L g419 ( 
.A(n_363),
.B(n_354),
.C(n_321),
.Y(n_419)
);

AOI22xp5_ASAP7_75t_L g420 ( 
.A1(n_367),
.A2(n_324),
.B1(n_360),
.B2(n_362),
.Y(n_420)
);

INVxp67_ASAP7_75t_L g423 ( 
.A(n_389),
.Y(n_423)
);

NOR2xp33_ASAP7_75t_L g473 ( 
.A(n_423),
.B(n_458),
.Y(n_473)
);

AND2x2_ASAP7_75t_L g463 ( 
.A(n_424),
.B(n_425),
.Y(n_463)
);

OAI22xp5_ASAP7_75t_SL g425 ( 
.A1(n_406),
.A2(n_362),
.B1(n_349),
.B2(n_363),
.Y(n_425)
);

OAI22xp5_ASAP7_75t_SL g428 ( 
.A1(n_418),
.A2(n_349),
.B1(n_320),
.B2(n_366),
.Y(n_428)
);

OAI22xp5_ASAP7_75t_SL g462 ( 
.A1(n_428),
.A2(n_435),
.B1(n_446),
.B2(n_448),
.Y(n_462)
);

OAI21xp5_ASAP7_75t_L g433 ( 
.A1(n_383),
.A2(n_316),
.B(n_323),
.Y(n_433)
);

OAI21xp5_ASAP7_75t_SL g480 ( 
.A1(n_433),
.A2(n_437),
.B(n_451),
.Y(n_480)
);

XNOR2xp5_ASAP7_75t_SL g482 ( 
.A(n_436),
.B(n_440),
.Y(n_482)
);

OAI21xp5_ASAP7_75t_L g437 ( 
.A1(n_413),
.A2(n_316),
.B(n_323),
.Y(n_437)
);

CKINVDCx20_ASAP7_75t_R g438 ( 
.A(n_394),
.Y(n_438)
);

CKINVDCx14_ASAP7_75t_R g467 ( 
.A(n_438),
.Y(n_467)
);

XNOR2xp5_ASAP7_75t_L g440 ( 
.A(n_411),
.B(n_359),
.Y(n_440)
);

OAI22xp5_ASAP7_75t_L g441 ( 
.A1(n_405),
.A2(n_342),
.B1(n_320),
.B2(n_366),
.Y(n_441)
);

OAI22xp5_ASAP7_75t_L g478 ( 
.A1(n_441),
.A2(n_444),
.B1(n_392),
.B2(n_401),
.Y(n_478)
);

XNOR2xp5_ASAP7_75t_L g443 ( 
.A(n_385),
.B(n_312),
.Y(n_443)
);

MAJIxp5_ASAP7_75t_L g489 ( 
.A(n_443),
.B(n_388),
.C(n_412),
.Y(n_489)
);

OAI22xp5_ASAP7_75t_L g444 ( 
.A1(n_420),
.A2(n_342),
.B1(n_371),
.B2(n_332),
.Y(n_444)
);

OAI22xp5_ASAP7_75t_SL g446 ( 
.A1(n_416),
.A2(n_348),
.B1(n_361),
.B2(n_336),
.Y(n_446)
);

OAI22xp5_ASAP7_75t_SL g448 ( 
.A1(n_416),
.A2(n_348),
.B1(n_336),
.B2(n_343),
.Y(n_448)
);

NOR2xp33_ASAP7_75t_L g449 ( 
.A(n_382),
.B(n_364),
.Y(n_449)
);

OR2x2_ASAP7_75t_L g487 ( 
.A(n_449),
.B(n_452),
.Y(n_487)
);

OAI21xp5_ASAP7_75t_L g451 ( 
.A1(n_375),
.A2(n_329),
.B(n_364),
.Y(n_451)
);

NAND2xp5_ASAP7_75t_SL g486 ( 
.A(n_453),
.B(n_459),
.Y(n_486)
);

NAND2xp5_ASAP7_75t_L g454 ( 
.A(n_380),
.B(n_387),
.Y(n_454)
);

INVx1_ASAP7_75t_L g465 ( 
.A(n_454),
.Y(n_465)
);

OAI21xp5_ASAP7_75t_SL g455 ( 
.A1(n_386),
.A2(n_416),
.B(n_393),
.Y(n_455)
);

OAI21xp5_ASAP7_75t_SL g483 ( 
.A1(n_455),
.A2(n_392),
.B(n_374),
.Y(n_483)
);

OAI22xp5_ASAP7_75t_SL g457 ( 
.A1(n_390),
.A2(n_380),
.B1(n_407),
.B2(n_397),
.Y(n_457)
);

OAI22xp5_ASAP7_75t_SL g477 ( 
.A1(n_457),
.A2(n_387),
.B1(n_390),
.B2(n_408),
.Y(n_477)
);

CKINVDCx20_ASAP7_75t_R g458 ( 
.A(n_394),
.Y(n_458)
);

NOR2xp33_ASAP7_75t_L g459 ( 
.A(n_382),
.B(n_419),
.Y(n_459)
);

OAI21xp5_ASAP7_75t_L g464 ( 
.A1(n_455),
.A2(n_392),
.B(n_374),
.Y(n_464)
);

OAI21xp5_ASAP7_75t_SL g517 ( 
.A1(n_464),
.A2(n_483),
.B(n_488),
.Y(n_517)
);

INVx1_ASAP7_75t_L g466 ( 
.A(n_442),
.Y(n_466)
);

INVx1_ASAP7_75t_L g507 ( 
.A(n_466),
.Y(n_507)
);

CKINVDCx20_ASAP7_75t_R g468 ( 
.A(n_453),
.Y(n_468)
);

NAND2xp5_ASAP7_75t_L g504 ( 
.A(n_468),
.B(n_469),
.Y(n_504)
);

CKINVDCx16_ASAP7_75t_R g469 ( 
.A(n_437),
.Y(n_469)
);

INVx1_ASAP7_75t_L g470 ( 
.A(n_442),
.Y(n_470)
);

INVx1_ASAP7_75t_L g515 ( 
.A(n_470),
.Y(n_515)
);

INVx1_ASAP7_75t_L g471 ( 
.A(n_445),
.Y(n_471)
);

INVx1_ASAP7_75t_L g527 ( 
.A(n_471),
.Y(n_527)
);

HB1xp67_ASAP7_75t_L g472 ( 
.A(n_434),
.Y(n_472)
);

INVx1_ASAP7_75t_L g529 ( 
.A(n_472),
.Y(n_529)
);

XNOR2xp5_ASAP7_75t_L g474 ( 
.A(n_460),
.B(n_417),
.Y(n_474)
);

XOR2xp5_ASAP7_75t_L g500 ( 
.A(n_474),
.B(n_494),
.Y(n_500)
);

INVx1_ASAP7_75t_L g475 ( 
.A(n_445),
.Y(n_475)
);

INVx1_ASAP7_75t_L g530 ( 
.A(n_475),
.Y(n_530)
);

INVx1_ASAP7_75t_L g476 ( 
.A(n_447),
.Y(n_476)
);

NAND2xp5_ASAP7_75t_L g525 ( 
.A(n_476),
.B(n_485),
.Y(n_525)
);

HB1xp67_ASAP7_75t_L g516 ( 
.A(n_477),
.Y(n_516)
);

NAND2xp5_ASAP7_75t_L g528 ( 
.A(n_478),
.B(n_481),
.Y(n_528)
);

INVx2_ASAP7_75t_L g479 ( 
.A(n_447),
.Y(n_479)
);

INVxp67_ASAP7_75t_L g509 ( 
.A(n_479),
.Y(n_509)
);

INVx2_ASAP7_75t_SL g481 ( 
.A(n_450),
.Y(n_481)
);

INVx2_ASAP7_75t_L g484 ( 
.A(n_450),
.Y(n_484)
);

INVxp67_ASAP7_75t_L g522 ( 
.A(n_484),
.Y(n_522)
);

INVx1_ASAP7_75t_L g485 ( 
.A(n_461),
.Y(n_485)
);

OAI21xp5_ASAP7_75t_L g488 ( 
.A1(n_429),
.A2(n_373),
.B(n_379),
.Y(n_488)
);

MAJIxp5_ASAP7_75t_L g501 ( 
.A(n_489),
.B(n_490),
.C(n_495),
.Y(n_501)
);

XOR2xp5_ASAP7_75t_L g490 ( 
.A(n_426),
.B(n_384),
.Y(n_490)
);

CKINVDCx20_ASAP7_75t_R g491 ( 
.A(n_431),
.Y(n_491)
);

NAND2xp5_ASAP7_75t_L g535 ( 
.A(n_491),
.B(n_492),
.Y(n_535)
);

INVx1_ASAP7_75t_L g492 ( 
.A(n_461),
.Y(n_492)
);

AOI21xp5_ASAP7_75t_L g493 ( 
.A1(n_456),
.A2(n_378),
.B(n_391),
.Y(n_493)
);

AOI21xp5_ASAP7_75t_L g521 ( 
.A1(n_493),
.A2(n_464),
.B(n_480),
.Y(n_521)
);

XNOR2xp5_ASAP7_75t_L g494 ( 
.A(n_460),
.B(n_403),
.Y(n_494)
);

XOR2xp5_ASAP7_75t_L g495 ( 
.A(n_426),
.B(n_415),
.Y(n_495)
);

INVx1_ASAP7_75t_L g496 ( 
.A(n_441),
.Y(n_496)
);

NOR2xp33_ASAP7_75t_L g534 ( 
.A(n_496),
.B(n_497),
.Y(n_534)
);

INVxp33_ASAP7_75t_SL g497 ( 
.A(n_431),
.Y(n_497)
);

OAI22xp5_ASAP7_75t_L g498 ( 
.A1(n_435),
.A2(n_408),
.B1(n_396),
.B2(n_402),
.Y(n_498)
);

AOI22xp5_ASAP7_75t_L g508 ( 
.A1(n_498),
.A2(n_424),
.B1(n_457),
.B2(n_425),
.Y(n_508)
);

CKINVDCx20_ASAP7_75t_R g499 ( 
.A(n_433),
.Y(n_499)
);

CKINVDCx14_ASAP7_75t_R g510 ( 
.A(n_499),
.Y(n_510)
);

XOR2xp5_ASAP7_75t_SL g502 ( 
.A(n_488),
.B(n_439),
.Y(n_502)
);

NOR2xp33_ASAP7_75t_L g540 ( 
.A(n_502),
.B(n_487),
.Y(n_540)
);

MAJIxp5_ASAP7_75t_L g503 ( 
.A(n_490),
.B(n_426),
.C(n_460),
.Y(n_503)
);

MAJIxp5_ASAP7_75t_L g541 ( 
.A(n_503),
.B(n_513),
.C(n_524),
.Y(n_541)
);

XOR2xp5_ASAP7_75t_L g505 ( 
.A(n_474),
.B(n_443),
.Y(n_505)
);

XOR2xp5_ASAP7_75t_L g543 ( 
.A(n_505),
.B(n_506),
.Y(n_543)
);

XNOR2x1_ASAP7_75t_L g506 ( 
.A(n_495),
.B(n_443),
.Y(n_506)
);

AOI22xp5_ASAP7_75t_L g536 ( 
.A1(n_508),
.A2(n_526),
.B1(n_532),
.B2(n_498),
.Y(n_536)
);

XNOR2x2_ASAP7_75t_L g511 ( 
.A(n_487),
.B(n_454),
.Y(n_511)
);

XNOR2xp5_ASAP7_75t_L g550 ( 
.A(n_511),
.B(n_480),
.Y(n_550)
);

NAND2xp5_ASAP7_75t_SL g512 ( 
.A(n_491),
.B(n_427),
.Y(n_512)
);

NOR2xp33_ASAP7_75t_SL g538 ( 
.A(n_512),
.B(n_519),
.Y(n_538)
);

MAJIxp5_ASAP7_75t_L g513 ( 
.A(n_489),
.B(n_440),
.C(n_459),
.Y(n_513)
);

OAI21xp5_ASAP7_75t_L g514 ( 
.A1(n_483),
.A2(n_429),
.B(n_456),
.Y(n_514)
);

OAI21xp5_ASAP7_75t_SL g537 ( 
.A1(n_514),
.A2(n_521),
.B(n_533),
.Y(n_537)
);

XNOR2xp5_ASAP7_75t_L g518 ( 
.A(n_494),
.B(n_436),
.Y(n_518)
);

XOR2xp5_ASAP7_75t_L g554 ( 
.A(n_518),
.B(n_520),
.Y(n_554)
);

BUFx24_ASAP7_75t_SL g519 ( 
.A(n_465),
.Y(n_519)
);

XNOR2xp5_ASAP7_75t_L g520 ( 
.A(n_482),
.B(n_439),
.Y(n_520)
);

XOR2xp5_ASAP7_75t_L g523 ( 
.A(n_482),
.B(n_452),
.Y(n_523)
);

XOR2xp5_ASAP7_75t_L g555 ( 
.A(n_523),
.B(n_476),
.Y(n_555)
);

MAJIxp5_ASAP7_75t_L g524 ( 
.A(n_486),
.B(n_451),
.C(n_449),
.Y(n_524)
);

AOI22xp5_ASAP7_75t_L g526 ( 
.A1(n_463),
.A2(n_428),
.B1(n_432),
.B2(n_421),
.Y(n_526)
);

MAJIxp5_ASAP7_75t_L g531 ( 
.A(n_465),
.B(n_446),
.C(n_448),
.Y(n_531)
);

MAJIxp5_ASAP7_75t_L g548 ( 
.A(n_531),
.B(n_496),
.C(n_462),
.Y(n_548)
);

OAI22xp5_ASAP7_75t_SL g532 ( 
.A1(n_463),
.A2(n_421),
.B1(n_432),
.B2(n_396),
.Y(n_532)
);

AOI22xp5_ASAP7_75t_SL g533 ( 
.A1(n_463),
.A2(n_444),
.B1(n_398),
.B2(n_427),
.Y(n_533)
);

OAI22xp5_ASAP7_75t_SL g574 ( 
.A1(n_536),
.A2(n_539),
.B1(n_549),
.B2(n_526),
.Y(n_574)
);

AOI22xp5_ASAP7_75t_L g539 ( 
.A1(n_528),
.A2(n_462),
.B1(n_493),
.B2(n_477),
.Y(n_539)
);

AOI22xp5_ASAP7_75t_SL g567 ( 
.A1(n_540),
.A2(n_504),
.B1(n_516),
.B2(n_511),
.Y(n_567)
);

INVx1_ASAP7_75t_L g542 ( 
.A(n_535),
.Y(n_542)
);

INVx1_ASAP7_75t_L g570 ( 
.A(n_542),
.Y(n_570)
);

NAND2xp5_ASAP7_75t_SL g544 ( 
.A(n_513),
.B(n_376),
.Y(n_544)
);

NOR2xp33_ASAP7_75t_SL g569 ( 
.A(n_544),
.B(n_545),
.Y(n_569)
);

NOR2xp33_ASAP7_75t_L g545 ( 
.A(n_534),
.B(n_377),
.Y(n_545)
);

NAND2xp5_ASAP7_75t_L g546 ( 
.A(n_522),
.B(n_473),
.Y(n_546)
);

INVx1_ASAP7_75t_L g575 ( 
.A(n_546),
.Y(n_575)
);

NAND2xp5_ASAP7_75t_L g547 ( 
.A(n_522),
.B(n_468),
.Y(n_547)
);

INVx1_ASAP7_75t_L g582 ( 
.A(n_547),
.Y(n_582)
);

XNOR2xp5_ASAP7_75t_L g583 ( 
.A(n_548),
.B(n_557),
.Y(n_583)
);

AOI22xp5_ASAP7_75t_L g549 ( 
.A1(n_528),
.A2(n_478),
.B1(n_499),
.B2(n_467),
.Y(n_549)
);

MAJx2_ASAP7_75t_L g573 ( 
.A(n_550),
.B(n_555),
.C(n_559),
.Y(n_573)
);

NAND2xp5_ASAP7_75t_SL g551 ( 
.A(n_500),
.B(n_409),
.Y(n_551)
);

NAND2xp5_ASAP7_75t_L g579 ( 
.A(n_551),
.B(n_553),
.Y(n_579)
);

MAJIxp5_ASAP7_75t_L g552 ( 
.A(n_501),
.B(n_466),
.C(n_470),
.Y(n_552)
);

MAJIxp5_ASAP7_75t_L g577 ( 
.A(n_552),
.B(n_560),
.C(n_524),
.Y(n_577)
);

NAND2xp5_ASAP7_75t_L g553 ( 
.A(n_509),
.B(n_535),
.Y(n_553)
);

INVx1_ASAP7_75t_L g556 ( 
.A(n_525),
.Y(n_556)
);

NAND2xp5_ASAP7_75t_L g578 ( 
.A(n_556),
.B(n_563),
.Y(n_578)
);

XNOR2xp5_ASAP7_75t_L g557 ( 
.A(n_500),
.B(n_475),
.Y(n_557)
);

OAI21xp5_ASAP7_75t_L g558 ( 
.A1(n_521),
.A2(n_481),
.B(n_492),
.Y(n_558)
);

OAI21xp5_ASAP7_75t_SL g572 ( 
.A1(n_558),
.A2(n_514),
.B(n_517),
.Y(n_572)
);

XOR2xp5_ASAP7_75t_L g559 ( 
.A(n_501),
.B(n_503),
.Y(n_559)
);

MAJIxp5_ASAP7_75t_L g560 ( 
.A(n_505),
.B(n_471),
.C(n_485),
.Y(n_560)
);

CKINVDCx20_ASAP7_75t_R g561 ( 
.A(n_510),
.Y(n_561)
);

NAND2xp5_ASAP7_75t_SL g566 ( 
.A(n_561),
.B(n_564),
.Y(n_566)
);

XNOR2xp5_ASAP7_75t_L g562 ( 
.A(n_518),
.B(n_479),
.Y(n_562)
);

XNOR2xp5_ASAP7_75t_L g588 ( 
.A(n_562),
.B(n_530),
.Y(n_588)
);

INVxp67_ASAP7_75t_L g563 ( 
.A(n_529),
.Y(n_563)
);

NAND2xp5_ASAP7_75t_SL g564 ( 
.A(n_502),
.B(n_400),
.Y(n_564)
);

INVx1_ASAP7_75t_L g565 ( 
.A(n_507),
.Y(n_565)
);

NAND2xp5_ASAP7_75t_L g581 ( 
.A(n_565),
.B(n_527),
.Y(n_581)
);

OAI22xp5_ASAP7_75t_L g604 ( 
.A1(n_567),
.A2(n_585),
.B1(n_580),
.B2(n_575),
.Y(n_604)
);

XOR2xp5_ASAP7_75t_L g568 ( 
.A(n_543),
.B(n_506),
.Y(n_568)
);

XOR2xp5_ASAP7_75t_L g602 ( 
.A(n_568),
.B(n_576),
.Y(n_602)
);

HB1xp67_ASAP7_75t_L g571 ( 
.A(n_562),
.Y(n_571)
);

INVx1_ASAP7_75t_L g590 ( 
.A(n_571),
.Y(n_590)
);

AOI21xp5_ASAP7_75t_SL g592 ( 
.A1(n_572),
.A2(n_537),
.B(n_558),
.Y(n_592)
);

AOI22xp5_ASAP7_75t_L g601 ( 
.A1(n_574),
.A2(n_539),
.B1(n_547),
.B2(n_553),
.Y(n_601)
);

XOR2xp5_ASAP7_75t_L g576 ( 
.A(n_543),
.B(n_517),
.Y(n_576)
);

XNOR2xp5_ASAP7_75t_L g593 ( 
.A(n_577),
.B(n_584),
.Y(n_593)
);

AOI21xp5_ASAP7_75t_L g580 ( 
.A1(n_537),
.A2(n_508),
.B(n_531),
.Y(n_580)
);

INVxp67_ASAP7_75t_L g589 ( 
.A(n_580),
.Y(n_589)
);

INVx1_ASAP7_75t_L g599 ( 
.A(n_581),
.Y(n_599)
);

XOR2xp5_ASAP7_75t_L g584 ( 
.A(n_557),
.B(n_559),
.Y(n_584)
);

AOI22xp5_ASAP7_75t_L g585 ( 
.A1(n_536),
.A2(n_532),
.B1(n_533),
.B2(n_509),
.Y(n_585)
);

MAJIxp5_ASAP7_75t_SL g586 ( 
.A(n_550),
.B(n_520),
.C(n_523),
.Y(n_586)
);

XNOR2xp5_ASAP7_75t_L g597 ( 
.A(n_586),
.B(n_588),
.Y(n_597)
);

BUFx12_ASAP7_75t_L g587 ( 
.A(n_560),
.Y(n_587)
);

NAND2xp5_ASAP7_75t_L g591 ( 
.A(n_587),
.B(n_552),
.Y(n_591)
);

NAND2xp5_ASAP7_75t_L g616 ( 
.A(n_591),
.B(n_595),
.Y(n_616)
);

XOR2xp5_ASAP7_75t_L g610 ( 
.A(n_592),
.B(n_572),
.Y(n_610)
);

NAND2xp5_ASAP7_75t_L g594 ( 
.A(n_566),
.B(n_563),
.Y(n_594)
);

INVx1_ASAP7_75t_L g621 ( 
.A(n_594),
.Y(n_621)
);

NAND3xp33_ASAP7_75t_L g595 ( 
.A(n_569),
.B(n_538),
.C(n_541),
.Y(n_595)
);

MAJIxp5_ASAP7_75t_L g596 ( 
.A(n_584),
.B(n_541),
.C(n_548),
.Y(n_596)
);

NAND2xp5_ASAP7_75t_SL g623 ( 
.A(n_596),
.B(n_598),
.Y(n_623)
);

MAJIxp5_ASAP7_75t_L g598 ( 
.A(n_577),
.B(n_554),
.C(n_555),
.Y(n_598)
);

MAJIxp5_ASAP7_75t_L g600 ( 
.A(n_583),
.B(n_554),
.C(n_549),
.Y(n_600)
);

XNOR2xp5_ASAP7_75t_L g613 ( 
.A(n_600),
.B(n_605),
.Y(n_613)
);

AOI22xp5_ASAP7_75t_L g608 ( 
.A1(n_601),
.A2(n_603),
.B1(n_604),
.B2(n_607),
.Y(n_608)
);

NOR2xp33_ASAP7_75t_L g603 ( 
.A(n_579),
.B(n_556),
.Y(n_603)
);

MAJIxp5_ASAP7_75t_L g605 ( 
.A(n_583),
.B(n_546),
.C(n_484),
.Y(n_605)
);

INVx1_ASAP7_75t_L g606 ( 
.A(n_578),
.Y(n_606)
);

NOR2xp33_ASAP7_75t_L g611 ( 
.A(n_606),
.B(n_582),
.Y(n_611)
);

NOR2xp33_ASAP7_75t_L g607 ( 
.A(n_578),
.B(n_434),
.Y(n_607)
);

MAJx2_ASAP7_75t_L g609 ( 
.A(n_600),
.B(n_573),
.C(n_576),
.Y(n_609)
);

NAND2xp5_ASAP7_75t_L g625 ( 
.A(n_609),
.B(n_611),
.Y(n_625)
);

OAI21xp5_ASAP7_75t_L g628 ( 
.A1(n_610),
.A2(n_622),
.B(n_592),
.Y(n_628)
);

XOR2xp5_ASAP7_75t_L g612 ( 
.A(n_602),
.B(n_573),
.Y(n_612)
);

AND2x2_ASAP7_75t_L g629 ( 
.A(n_612),
.B(n_615),
.Y(n_629)
);

NOR2xp33_ASAP7_75t_L g614 ( 
.A(n_605),
.B(n_589),
.Y(n_614)
);

NAND2xp5_ASAP7_75t_L g634 ( 
.A(n_614),
.B(n_617),
.Y(n_634)
);

XOR2xp5_ASAP7_75t_L g615 ( 
.A(n_602),
.B(n_568),
.Y(n_615)
);

XNOR2xp5_ASAP7_75t_L g617 ( 
.A(n_593),
.B(n_567),
.Y(n_617)
);

NOR2xp33_ASAP7_75t_L g618 ( 
.A(n_589),
.B(n_570),
.Y(n_618)
);

NOR2xp33_ASAP7_75t_SL g626 ( 
.A(n_618),
.B(n_515),
.Y(n_626)
);

MAJIxp5_ASAP7_75t_L g619 ( 
.A(n_596),
.B(n_588),
.C(n_574),
.Y(n_619)
);

NAND2xp5_ASAP7_75t_SL g630 ( 
.A(n_619),
.B(n_620),
.Y(n_630)
);

MAJIxp5_ASAP7_75t_L g620 ( 
.A(n_593),
.B(n_587),
.C(n_585),
.Y(n_620)
);

AOI21xp5_ASAP7_75t_SL g622 ( 
.A1(n_599),
.A2(n_581),
.B(n_565),
.Y(n_622)
);

MAJIxp5_ASAP7_75t_L g624 ( 
.A(n_620),
.B(n_598),
.C(n_590),
.Y(n_624)
);

NAND2xp5_ASAP7_75t_L g636 ( 
.A(n_624),
.B(n_627),
.Y(n_636)
);

NAND2xp5_ASAP7_75t_SL g637 ( 
.A(n_626),
.B(n_632),
.Y(n_637)
);

AOI21xp5_ASAP7_75t_L g627 ( 
.A1(n_616),
.A2(n_610),
.B(n_623),
.Y(n_627)
);

NAND2xp5_ASAP7_75t_L g638 ( 
.A(n_628),
.B(n_631),
.Y(n_638)
);

AOI21xp5_ASAP7_75t_L g631 ( 
.A1(n_621),
.A2(n_619),
.B(n_608),
.Y(n_631)
);

OAI21xp5_ASAP7_75t_SL g632 ( 
.A1(n_622),
.A2(n_601),
.B(n_587),
.Y(n_632)
);

OAI22xp5_ASAP7_75t_SL g633 ( 
.A1(n_609),
.A2(n_586),
.B1(n_597),
.B2(n_481),
.Y(n_633)
);

INVxp67_ASAP7_75t_L g639 ( 
.A(n_633),
.Y(n_639)
);

O2A1O1Ixp33_ASAP7_75t_L g635 ( 
.A1(n_612),
.A2(n_597),
.B(n_422),
.C(n_430),
.Y(n_635)
);

NAND2xp5_ASAP7_75t_L g641 ( 
.A(n_635),
.B(n_458),
.Y(n_641)
);

MAJIxp5_ASAP7_75t_L g640 ( 
.A(n_630),
.B(n_613),
.C(n_615),
.Y(n_640)
);

NAND2xp5_ASAP7_75t_SL g647 ( 
.A(n_640),
.B(n_642),
.Y(n_647)
);

INVxp67_ASAP7_75t_L g649 ( 
.A(n_641),
.Y(n_649)
);

NAND2xp5_ASAP7_75t_L g642 ( 
.A(n_634),
.B(n_430),
.Y(n_642)
);

NOR2xp33_ASAP7_75t_L g643 ( 
.A(n_624),
.B(n_438),
.Y(n_643)
);

NOR2xp33_ASAP7_75t_SL g645 ( 
.A(n_643),
.B(n_625),
.Y(n_645)
);

XOR2xp5_ASAP7_75t_L g644 ( 
.A(n_628),
.B(n_422),
.Y(n_644)
);

NOR2xp33_ASAP7_75t_L g648 ( 
.A(n_644),
.B(n_629),
.Y(n_648)
);

OAI21xp5_ASAP7_75t_L g652 ( 
.A1(n_645),
.A2(n_646),
.B(n_648),
.Y(n_652)
);

NAND4xp25_ASAP7_75t_L g646 ( 
.A(n_636),
.B(n_633),
.C(n_629),
.D(n_635),
.Y(n_646)
);

AOI21xp5_ASAP7_75t_L g650 ( 
.A1(n_647),
.A2(n_638),
.B(n_637),
.Y(n_650)
);

OAI321xp33_ASAP7_75t_L g654 ( 
.A1(n_650),
.A2(n_381),
.A3(n_395),
.B1(n_410),
.B2(n_414),
.C(n_652),
.Y(n_654)
);

MAJIxp5_ASAP7_75t_L g651 ( 
.A(n_649),
.B(n_639),
.C(n_644),
.Y(n_651)
);

MAJIxp5_ASAP7_75t_L g653 ( 
.A(n_651),
.B(n_639),
.C(n_404),
.Y(n_653)
);

MAJIxp5_ASAP7_75t_L g655 ( 
.A(n_653),
.B(n_654),
.C(n_381),
.Y(n_655)
);

NAND2xp5_ASAP7_75t_SL g656 ( 
.A(n_655),
.B(n_395),
.Y(n_656)
);

BUFx24_ASAP7_75t_SL g657 ( 
.A(n_656),
.Y(n_657)
);


endmodule