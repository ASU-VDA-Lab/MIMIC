module fake_jpeg_10673_n_36 (n_3, n_2, n_1, n_0, n_4, n_5, n_36);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_5;

output n_36;

wire n_13;
wire n_21;
wire n_33;
wire n_10;
wire n_23;
wire n_27;
wire n_6;
wire n_22;
wire n_14;
wire n_19;
wire n_18;
wire n_20;
wire n_35;
wire n_34;
wire n_30;
wire n_16;
wire n_24;
wire n_28;
wire n_26;
wire n_9;
wire n_11;
wire n_17;
wire n_25;
wire n_31;
wire n_29;
wire n_12;
wire n_32;
wire n_8;
wire n_15;
wire n_7;

NAND2xp5_ASAP7_75t_L g6 ( 
.A(n_1),
.B(n_2),
.Y(n_6)
);

CKINVDCx20_ASAP7_75t_R g7 ( 
.A(n_3),
.Y(n_7)
);

INVx1_ASAP7_75t_L g8 ( 
.A(n_4),
.Y(n_8)
);

BUFx6f_ASAP7_75t_L g9 ( 
.A(n_1),
.Y(n_9)
);

INVx8_ASAP7_75t_L g10 ( 
.A(n_5),
.Y(n_10)
);

INVx3_ASAP7_75t_L g11 ( 
.A(n_0),
.Y(n_11)
);

NAND2xp5_ASAP7_75t_L g12 ( 
.A(n_6),
.B(n_0),
.Y(n_12)
);

NAND2xp5_ASAP7_75t_L g22 ( 
.A(n_12),
.B(n_14),
.Y(n_22)
);

OAI22xp5_ASAP7_75t_L g13 ( 
.A1(n_11),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_13)
);

AOI22xp5_ASAP7_75t_L g18 ( 
.A1(n_13),
.A2(n_11),
.B1(n_10),
.B2(n_8),
.Y(n_18)
);

INVx1_ASAP7_75t_L g14 ( 
.A(n_6),
.Y(n_14)
);

NOR2xp33_ASAP7_75t_L g15 ( 
.A(n_6),
.B(n_2),
.Y(n_15)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_15),
.Y(n_19)
);

INVx13_ASAP7_75t_L g16 ( 
.A(n_10),
.Y(n_16)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_16),
.Y(n_20)
);

NAND2xp5_ASAP7_75t_SL g17 ( 
.A(n_7),
.B(n_3),
.Y(n_17)
);

NAND2xp5_ASAP7_75t_SL g21 ( 
.A(n_17),
.B(n_8),
.Y(n_21)
);

AOI22xp5_ASAP7_75t_L g23 ( 
.A1(n_18),
.A2(n_11),
.B1(n_10),
.B2(n_13),
.Y(n_23)
);

OAI21xp5_ASAP7_75t_SL g26 ( 
.A1(n_21),
.A2(n_17),
.B(n_14),
.Y(n_26)
);

XOR2xp5_ASAP7_75t_L g29 ( 
.A(n_23),
.B(n_24),
.Y(n_29)
);

XOR2xp5_ASAP7_75t_L g24 ( 
.A(n_22),
.B(n_12),
.Y(n_24)
);

INVxp67_ASAP7_75t_L g25 ( 
.A(n_20),
.Y(n_25)
);

AOI21xp5_ASAP7_75t_L g27 ( 
.A1(n_25),
.A2(n_26),
.B(n_22),
.Y(n_27)
);

NOR2xp33_ASAP7_75t_L g31 ( 
.A(n_27),
.B(n_19),
.Y(n_31)
);

AOI21xp5_ASAP7_75t_L g28 ( 
.A1(n_25),
.A2(n_18),
.B(n_7),
.Y(n_28)
);

XNOR2xp5_ASAP7_75t_L g30 ( 
.A(n_28),
.B(n_9),
.Y(n_30)
);

OAI21xp5_ASAP7_75t_L g32 ( 
.A1(n_30),
.A2(n_31),
.B(n_29),
.Y(n_32)
);

NAND2xp5_ASAP7_75t_L g34 ( 
.A(n_32),
.B(n_33),
.Y(n_34)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_30),
.Y(n_33)
);

OAI221xp5_ASAP7_75t_L g35 ( 
.A1(n_34),
.A2(n_16),
.B1(n_9),
.B2(n_5),
.C(n_4),
.Y(n_35)
);

AOI21xp5_ASAP7_75t_SL g36 ( 
.A1(n_35),
.A2(n_9),
.B(n_8),
.Y(n_36)
);


endmodule