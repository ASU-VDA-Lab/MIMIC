module fake_jpeg_3086_n_412 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_412);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_412;

wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_385;
wire n_228;
wire n_134;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_340;
wire n_381;
wire n_377;
wire n_291;
wire n_236;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_401;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_39;
wire n_371;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_305;
wire n_161;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_382;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_389;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_384;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_378;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_379;
wire n_114;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_409;
wire n_249;
wire n_217;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_391;
wire n_209;
wire n_22;
wire n_138;
wire n_402;
wire n_247;
wire n_157;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

BUFx8_ASAP7_75t_L g17 ( 
.A(n_3),
.Y(n_17)
);

BUFx12f_ASAP7_75t_L g18 ( 
.A(n_13),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_9),
.Y(n_19)
);

BUFx12f_ASAP7_75t_L g20 ( 
.A(n_4),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_6),
.Y(n_21)
);

BUFx12f_ASAP7_75t_L g22 ( 
.A(n_9),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_14),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_5),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_16),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_11),
.Y(n_26)
);

BUFx3_ASAP7_75t_L g27 ( 
.A(n_1),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_0),
.Y(n_28)
);

INVx2_ASAP7_75t_L g29 ( 
.A(n_2),
.Y(n_29)
);

BUFx16f_ASAP7_75t_L g30 ( 
.A(n_9),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_13),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_5),
.Y(n_32)
);

INVx8_ASAP7_75t_L g33 ( 
.A(n_3),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_6),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_16),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_16),
.Y(n_36)
);

BUFx3_ASAP7_75t_L g37 ( 
.A(n_5),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_14),
.Y(n_38)
);

INVx2_ASAP7_75t_L g39 ( 
.A(n_11),
.Y(n_39)
);

BUFx3_ASAP7_75t_L g40 ( 
.A(n_2),
.Y(n_40)
);

INVx3_ASAP7_75t_L g41 ( 
.A(n_12),
.Y(n_41)
);

BUFx10_ASAP7_75t_L g42 ( 
.A(n_12),
.Y(n_42)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_7),
.Y(n_43)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_0),
.Y(n_44)
);

INVx1_ASAP7_75t_SL g45 ( 
.A(n_14),
.Y(n_45)
);

CKINVDCx16_ASAP7_75t_R g46 ( 
.A(n_11),
.Y(n_46)
);

BUFx3_ASAP7_75t_L g47 ( 
.A(n_8),
.Y(n_47)
);

INVx3_ASAP7_75t_L g48 ( 
.A(n_7),
.Y(n_48)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_10),
.Y(n_49)
);

INVx2_ASAP7_75t_L g50 ( 
.A(n_0),
.Y(n_50)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_6),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_3),
.Y(n_52)
);

INVx2_ASAP7_75t_R g53 ( 
.A(n_0),
.Y(n_53)
);

INVx8_ASAP7_75t_L g54 ( 
.A(n_20),
.Y(n_54)
);

BUFx2_ASAP7_75t_L g115 ( 
.A(n_54),
.Y(n_115)
);

CKINVDCx20_ASAP7_75t_R g55 ( 
.A(n_30),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g119 ( 
.A(n_55),
.B(n_56),
.Y(n_119)
);

CKINVDCx20_ASAP7_75t_R g56 ( 
.A(n_30),
.Y(n_56)
);

INVx3_ASAP7_75t_SL g57 ( 
.A(n_17),
.Y(n_57)
);

BUFx2_ASAP7_75t_L g148 ( 
.A(n_57),
.Y(n_148)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_39),
.Y(n_58)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_58),
.Y(n_116)
);

INVx8_ASAP7_75t_L g59 ( 
.A(n_20),
.Y(n_59)
);

INVx3_ASAP7_75t_L g133 ( 
.A(n_59),
.Y(n_133)
);

CKINVDCx20_ASAP7_75t_R g60 ( 
.A(n_30),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g146 ( 
.A(n_60),
.B(n_70),
.Y(n_146)
);

INVx11_ASAP7_75t_L g61 ( 
.A(n_17),
.Y(n_61)
);

INVx4_ASAP7_75t_L g127 ( 
.A(n_61),
.Y(n_127)
);

INVx8_ASAP7_75t_L g62 ( 
.A(n_20),
.Y(n_62)
);

INVx3_ASAP7_75t_L g167 ( 
.A(n_62),
.Y(n_167)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_52),
.Y(n_63)
);

BUFx6f_ASAP7_75t_L g124 ( 
.A(n_63),
.Y(n_124)
);

INVx2_ASAP7_75t_L g64 ( 
.A(n_29),
.Y(n_64)
);

INVx2_ASAP7_75t_L g113 ( 
.A(n_64),
.Y(n_113)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_52),
.Y(n_65)
);

BUFx6f_ASAP7_75t_L g128 ( 
.A(n_65),
.Y(n_128)
);

INVx4_ASAP7_75t_L g66 ( 
.A(n_20),
.Y(n_66)
);

INVx2_ASAP7_75t_SL g134 ( 
.A(n_66),
.Y(n_134)
);

INVx4_ASAP7_75t_SL g67 ( 
.A(n_17),
.Y(n_67)
);

BUFx3_ASAP7_75t_L g157 ( 
.A(n_67),
.Y(n_157)
);

INVx2_ASAP7_75t_L g68 ( 
.A(n_29),
.Y(n_68)
);

INVx2_ASAP7_75t_L g139 ( 
.A(n_68),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_19),
.B(n_8),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_L g118 ( 
.A(n_69),
.B(n_75),
.Y(n_118)
);

CKINVDCx20_ASAP7_75t_R g70 ( 
.A(n_52),
.Y(n_70)
);

INVxp67_ASAP7_75t_L g71 ( 
.A(n_17),
.Y(n_71)
);

CKINVDCx6p67_ASAP7_75t_R g147 ( 
.A(n_71),
.Y(n_147)
);

BUFx12f_ASAP7_75t_L g72 ( 
.A(n_33),
.Y(n_72)
);

INVx4_ASAP7_75t_L g137 ( 
.A(n_72),
.Y(n_137)
);

INVx3_ASAP7_75t_L g73 ( 
.A(n_18),
.Y(n_73)
);

HB1xp67_ASAP7_75t_L g162 ( 
.A(n_73),
.Y(n_162)
);

BUFx6f_ASAP7_75t_L g74 ( 
.A(n_27),
.Y(n_74)
);

BUFx6f_ASAP7_75t_L g143 ( 
.A(n_74),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_L g75 ( 
.A(n_39),
.B(n_8),
.Y(n_75)
);

INVx8_ASAP7_75t_L g76 ( 
.A(n_18),
.Y(n_76)
);

INVx4_ASAP7_75t_L g156 ( 
.A(n_76),
.Y(n_156)
);

INVx3_ASAP7_75t_L g77 ( 
.A(n_18),
.Y(n_77)
);

BUFx12f_ASAP7_75t_L g140 ( 
.A(n_77),
.Y(n_140)
);

INVx2_ASAP7_75t_L g78 ( 
.A(n_50),
.Y(n_78)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_78),
.Y(n_158)
);

CKINVDCx20_ASAP7_75t_R g79 ( 
.A(n_19),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g154 ( 
.A(n_79),
.B(n_89),
.Y(n_154)
);

INVx3_ASAP7_75t_SL g80 ( 
.A(n_33),
.Y(n_80)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_80),
.Y(n_168)
);

INVx2_ASAP7_75t_L g81 ( 
.A(n_50),
.Y(n_81)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_81),
.Y(n_171)
);

BUFx5_ASAP7_75t_L g82 ( 
.A(n_53),
.Y(n_82)
);

BUFx5_ASAP7_75t_L g138 ( 
.A(n_82),
.Y(n_138)
);

INVx6_ASAP7_75t_L g83 ( 
.A(n_18),
.Y(n_83)
);

BUFx6f_ASAP7_75t_L g149 ( 
.A(n_83),
.Y(n_149)
);

BUFx6f_ASAP7_75t_L g84 ( 
.A(n_27),
.Y(n_84)
);

INVx6_ASAP7_75t_L g114 ( 
.A(n_84),
.Y(n_114)
);

BUFx6f_ASAP7_75t_L g85 ( 
.A(n_40),
.Y(n_85)
);

BUFx12f_ASAP7_75t_L g151 ( 
.A(n_85),
.Y(n_151)
);

BUFx12f_ASAP7_75t_SL g86 ( 
.A(n_22),
.Y(n_86)
);

AND2x2_ASAP7_75t_L g144 ( 
.A(n_86),
.B(n_87),
.Y(n_144)
);

BUFx3_ASAP7_75t_L g87 ( 
.A(n_40),
.Y(n_87)
);

BUFx6f_ASAP7_75t_L g88 ( 
.A(n_22),
.Y(n_88)
);

CKINVDCx16_ASAP7_75t_R g160 ( 
.A(n_88),
.Y(n_160)
);

INVx4_ASAP7_75t_L g89 ( 
.A(n_22),
.Y(n_89)
);

INVx5_ASAP7_75t_L g90 ( 
.A(n_22),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g155 ( 
.A(n_90),
.B(n_93),
.Y(n_155)
);

INVx6_ASAP7_75t_L g91 ( 
.A(n_37),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_L g122 ( 
.A(n_91),
.B(n_92),
.Y(n_122)
);

BUFx6f_ASAP7_75t_L g92 ( 
.A(n_37),
.Y(n_92)
);

INVx3_ASAP7_75t_L g93 ( 
.A(n_47),
.Y(n_93)
);

CKINVDCx20_ASAP7_75t_R g94 ( 
.A(n_21),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g159 ( 
.A(n_94),
.B(n_98),
.Y(n_159)
);

BUFx6f_ASAP7_75t_L g95 ( 
.A(n_47),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g129 ( 
.A(n_95),
.B(n_97),
.Y(n_129)
);

INVx5_ASAP7_75t_L g96 ( 
.A(n_41),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g173 ( 
.A(n_96),
.B(n_105),
.Y(n_173)
);

INVx2_ASAP7_75t_L g97 ( 
.A(n_41),
.Y(n_97)
);

CKINVDCx20_ASAP7_75t_R g98 ( 
.A(n_21),
.Y(n_98)
);

INVx3_ASAP7_75t_L g99 ( 
.A(n_48),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g163 ( 
.A(n_99),
.B(n_101),
.Y(n_163)
);

BUFx6f_ASAP7_75t_L g100 ( 
.A(n_48),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_L g130 ( 
.A(n_100),
.B(n_102),
.Y(n_130)
);

BUFx3_ASAP7_75t_L g101 ( 
.A(n_45),
.Y(n_101)
);

INVx2_ASAP7_75t_L g102 ( 
.A(n_28),
.Y(n_102)
);

INVx2_ASAP7_75t_L g103 ( 
.A(n_28),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_L g132 ( 
.A(n_103),
.B(n_104),
.Y(n_132)
);

BUFx6f_ASAP7_75t_L g104 ( 
.A(n_44),
.Y(n_104)
);

CKINVDCx20_ASAP7_75t_R g105 ( 
.A(n_23),
.Y(n_105)
);

CKINVDCx20_ASAP7_75t_R g106 ( 
.A(n_23),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_SL g131 ( 
.A(n_106),
.B(n_26),
.Y(n_131)
);

INVx2_ASAP7_75t_SL g107 ( 
.A(n_44),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_L g152 ( 
.A(n_107),
.B(n_108),
.Y(n_152)
);

BUFx10_ASAP7_75t_L g108 ( 
.A(n_42),
.Y(n_108)
);

INVx5_ASAP7_75t_L g109 ( 
.A(n_42),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_L g153 ( 
.A(n_109),
.B(n_1),
.Y(n_153)
);

AOI22xp33_ASAP7_75t_SL g110 ( 
.A1(n_67),
.A2(n_45),
.B1(n_53),
.B2(n_31),
.Y(n_110)
);

AOI22xp33_ASAP7_75t_SL g181 ( 
.A1(n_110),
.A2(n_111),
.B1(n_166),
.B2(n_169),
.Y(n_181)
);

AOI22xp33_ASAP7_75t_SL g111 ( 
.A1(n_71),
.A2(n_53),
.B1(n_31),
.B2(n_38),
.Y(n_111)
);

AO22x1_ASAP7_75t_SL g112 ( 
.A1(n_57),
.A2(n_42),
.B1(n_51),
.B2(n_32),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_L g176 ( 
.A(n_112),
.B(n_110),
.Y(n_176)
);

AOI22xp5_ASAP7_75t_SL g117 ( 
.A1(n_96),
.A2(n_46),
.B1(n_51),
.B2(n_32),
.Y(n_117)
);

OR2x2_ASAP7_75t_L g210 ( 
.A(n_117),
.B(n_123),
.Y(n_210)
);

O2A1O1Ixp33_ASAP7_75t_SL g120 ( 
.A1(n_107),
.A2(n_42),
.B(n_49),
.C(n_26),
.Y(n_120)
);

A2O1A1Ixp33_ASAP7_75t_L g184 ( 
.A1(n_120),
.A2(n_165),
.B(n_144),
.C(n_147),
.Y(n_184)
);

OAI22xp5_ASAP7_75t_L g121 ( 
.A1(n_100),
.A2(n_24),
.B1(n_38),
.B2(n_49),
.Y(n_121)
);

AOI22xp5_ASAP7_75t_L g192 ( 
.A1(n_121),
.A2(n_125),
.B1(n_126),
.B2(n_136),
.Y(n_192)
);

OA22x2_ASAP7_75t_L g123 ( 
.A1(n_91),
.A2(n_43),
.B1(n_36),
.B2(n_35),
.Y(n_123)
);

AOI22xp33_ASAP7_75t_L g125 ( 
.A1(n_63),
.A2(n_34),
.B1(n_43),
.B2(n_36),
.Y(n_125)
);

OAI22xp5_ASAP7_75t_L g126 ( 
.A1(n_65),
.A2(n_24),
.B1(n_35),
.B2(n_34),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_L g174 ( 
.A(n_131),
.B(n_159),
.Y(n_174)
);

AOI22xp5_ASAP7_75t_SL g135 ( 
.A1(n_109),
.A2(n_46),
.B1(n_25),
.B2(n_10),
.Y(n_135)
);

NOR2x1_ASAP7_75t_L g198 ( 
.A(n_135),
.B(n_141),
.Y(n_198)
);

AOI22xp33_ASAP7_75t_L g136 ( 
.A1(n_61),
.A2(n_25),
.B1(n_2),
.B2(n_3),
.Y(n_136)
);

AOI22xp5_ASAP7_75t_SL g141 ( 
.A1(n_80),
.A2(n_10),
.B1(n_13),
.B2(n_12),
.Y(n_141)
);

OAI22xp5_ASAP7_75t_SL g142 ( 
.A1(n_92),
.A2(n_7),
.B1(n_15),
.B2(n_4),
.Y(n_142)
);

AOI22xp5_ASAP7_75t_L g220 ( 
.A1(n_142),
.A2(n_145),
.B1(n_150),
.B2(n_164),
.Y(n_220)
);

OAI22xp5_ASAP7_75t_SL g145 ( 
.A1(n_95),
.A2(n_15),
.B1(n_2),
.B2(n_4),
.Y(n_145)
);

AOI22xp33_ASAP7_75t_L g150 ( 
.A1(n_104),
.A2(n_1),
.B1(n_4),
.B2(n_15),
.Y(n_150)
);

AND2x2_ASAP7_75t_L g188 ( 
.A(n_153),
.B(n_127),
.Y(n_188)
);

AOI22xp5_ASAP7_75t_SL g161 ( 
.A1(n_101),
.A2(n_87),
.B1(n_89),
.B2(n_84),
.Y(n_161)
);

OAI21xp5_ASAP7_75t_L g221 ( 
.A1(n_161),
.A2(n_172),
.B(n_170),
.Y(n_221)
);

AOI22xp33_ASAP7_75t_L g164 ( 
.A1(n_74),
.A2(n_1),
.B1(n_85),
.B2(n_88),
.Y(n_164)
);

A2O1A1Ixp33_ASAP7_75t_L g165 ( 
.A1(n_108),
.A2(n_66),
.B(n_59),
.C(n_62),
.Y(n_165)
);

OAI22xp5_ASAP7_75t_SL g166 ( 
.A1(n_83),
.A2(n_72),
.B1(n_76),
.B2(n_54),
.Y(n_166)
);

AOI22xp33_ASAP7_75t_SL g169 ( 
.A1(n_72),
.A2(n_67),
.B1(n_71),
.B2(n_61),
.Y(n_169)
);

AOI22xp33_ASAP7_75t_SL g170 ( 
.A1(n_108),
.A2(n_67),
.B1(n_71),
.B2(n_61),
.Y(n_170)
);

AOI22xp33_ASAP7_75t_SL g197 ( 
.A1(n_170),
.A2(n_172),
.B1(n_157),
.B2(n_127),
.Y(n_197)
);

AOI22xp33_ASAP7_75t_SL g172 ( 
.A1(n_67),
.A2(n_71),
.B1(n_61),
.B2(n_17),
.Y(n_172)
);

NOR2xp33_ASAP7_75t_SL g242 ( 
.A(n_174),
.B(n_183),
.Y(n_242)
);

INVx8_ASAP7_75t_L g175 ( 
.A(n_151),
.Y(n_175)
);

INVx5_ASAP7_75t_L g264 ( 
.A(n_175),
.Y(n_264)
);

AND2x2_ASAP7_75t_L g262 ( 
.A(n_176),
.B(n_200),
.Y(n_262)
);

CKINVDCx20_ASAP7_75t_R g177 ( 
.A(n_154),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_SL g232 ( 
.A(n_177),
.B(n_182),
.Y(n_232)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_146),
.Y(n_178)
);

INVx1_ASAP7_75t_SL g247 ( 
.A(n_178),
.Y(n_247)
);

NAND2xp5_ASAP7_75t_L g179 ( 
.A(n_132),
.B(n_130),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_L g228 ( 
.A(n_179),
.B(n_191),
.Y(n_228)
);

HB1xp67_ASAP7_75t_L g180 ( 
.A(n_168),
.Y(n_180)
);

INVx1_ASAP7_75t_SL g257 ( 
.A(n_180),
.Y(n_257)
);

CKINVDCx20_ASAP7_75t_R g182 ( 
.A(n_119),
.Y(n_182)
);

NOR2xp33_ASAP7_75t_L g183 ( 
.A(n_118),
.B(n_173),
.Y(n_183)
);

A2O1A1Ixp33_ASAP7_75t_SL g235 ( 
.A1(n_184),
.A2(n_197),
.B(n_210),
.C(n_189),
.Y(n_235)
);

INVxp67_ASAP7_75t_L g185 ( 
.A(n_147),
.Y(n_185)
);

INVxp33_ASAP7_75t_L g241 ( 
.A(n_185),
.Y(n_241)
);

INVxp67_ASAP7_75t_L g186 ( 
.A(n_147),
.Y(n_186)
);

INVxp67_ASAP7_75t_L g245 ( 
.A(n_186),
.Y(n_245)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_148),
.Y(n_187)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_187),
.Y(n_251)
);

NAND2xp5_ASAP7_75t_SL g252 ( 
.A(n_188),
.B(n_195),
.Y(n_252)
);

AND2x2_ASAP7_75t_L g189 ( 
.A(n_144),
.B(n_152),
.Y(n_189)
);

CKINVDCx16_ASAP7_75t_R g261 ( 
.A(n_189),
.Y(n_261)
);

BUFx6f_ASAP7_75t_L g190 ( 
.A(n_124),
.Y(n_190)
);

INVx8_ASAP7_75t_L g244 ( 
.A(n_190),
.Y(n_244)
);

NAND2xp5_ASAP7_75t_L g191 ( 
.A(n_129),
.B(n_158),
.Y(n_191)
);

INVx2_ASAP7_75t_L g193 ( 
.A(n_134),
.Y(n_193)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_193),
.Y(n_265)
);

AOI22xp33_ASAP7_75t_L g194 ( 
.A1(n_120),
.A2(n_116),
.B1(n_123),
.B2(n_112),
.Y(n_194)
);

OAI22xp33_ASAP7_75t_SL g239 ( 
.A1(n_194),
.A2(n_209),
.B1(n_211),
.B2(n_222),
.Y(n_239)
);

CKINVDCx16_ASAP7_75t_R g195 ( 
.A(n_148),
.Y(n_195)
);

NOR2xp33_ASAP7_75t_L g196 ( 
.A(n_155),
.B(n_171),
.Y(n_196)
);

NOR2xp33_ASAP7_75t_SL g253 ( 
.A(n_196),
.B(n_203),
.Y(n_253)
);

INVx4_ASAP7_75t_L g199 ( 
.A(n_156),
.Y(n_199)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_199),
.Y(n_269)
);

INVx2_ASAP7_75t_L g200 ( 
.A(n_134),
.Y(n_200)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_162),
.Y(n_201)
);

NOR2xp33_ASAP7_75t_L g238 ( 
.A(n_201),
.B(n_205),
.Y(n_238)
);

NAND2xp5_ASAP7_75t_L g202 ( 
.A(n_122),
.B(n_139),
.Y(n_202)
);

NAND2xp5_ASAP7_75t_L g236 ( 
.A(n_202),
.B(n_206),
.Y(n_236)
);

NOR2xp33_ASAP7_75t_L g203 ( 
.A(n_163),
.B(n_113),
.Y(n_203)
);

INVx13_ASAP7_75t_L g204 ( 
.A(n_157),
.Y(n_204)
);

BUFx24_ASAP7_75t_L g255 ( 
.A(n_204),
.Y(n_255)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_133),
.Y(n_205)
);

NAND2xp5_ASAP7_75t_L g206 ( 
.A(n_112),
.B(n_123),
.Y(n_206)
);

INVx3_ASAP7_75t_L g207 ( 
.A(n_156),
.Y(n_207)
);

AND2x2_ASAP7_75t_L g268 ( 
.A(n_207),
.B(n_215),
.Y(n_268)
);

NAND2xp5_ASAP7_75t_L g208 ( 
.A(n_111),
.B(n_150),
.Y(n_208)
);

NAND2xp5_ASAP7_75t_L g248 ( 
.A(n_208),
.B(n_214),
.Y(n_248)
);

AOI22xp33_ASAP7_75t_SL g209 ( 
.A1(n_165),
.A2(n_167),
.B1(n_133),
.B2(n_115),
.Y(n_209)
);

AOI22xp33_ASAP7_75t_L g211 ( 
.A1(n_125),
.A2(n_164),
.B1(n_124),
.B2(n_128),
.Y(n_211)
);

HB1xp67_ASAP7_75t_L g212 ( 
.A(n_167),
.Y(n_212)
);

CKINVDCx20_ASAP7_75t_R g233 ( 
.A(n_212),
.Y(n_233)
);

CKINVDCx20_ASAP7_75t_R g213 ( 
.A(n_115),
.Y(n_213)
);

NOR2xp33_ASAP7_75t_L g240 ( 
.A(n_213),
.B(n_216),
.Y(n_240)
);

NAND2xp5_ASAP7_75t_L g214 ( 
.A(n_141),
.B(n_114),
.Y(n_214)
);

INVx2_ASAP7_75t_L g215 ( 
.A(n_114),
.Y(n_215)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_137),
.Y(n_216)
);

NOR2xp33_ASAP7_75t_L g217 ( 
.A(n_140),
.B(n_137),
.Y(n_217)
);

NOR2xp33_ASAP7_75t_L g243 ( 
.A(n_217),
.B(n_227),
.Y(n_243)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_149),
.Y(n_218)
);

OR2x2_ASAP7_75t_L g256 ( 
.A(n_218),
.B(n_219),
.Y(n_256)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_149),
.Y(n_219)
);

AOI21xp5_ASAP7_75t_L g231 ( 
.A1(n_221),
.A2(n_181),
.B(n_210),
.Y(n_231)
);

AOI22xp33_ASAP7_75t_SL g222 ( 
.A1(n_151),
.A2(n_140),
.B1(n_169),
.B2(n_136),
.Y(n_222)
);

NAND2xp5_ASAP7_75t_L g223 ( 
.A(n_128),
.B(n_143),
.Y(n_223)
);

NAND2xp5_ASAP7_75t_L g258 ( 
.A(n_223),
.B(n_190),
.Y(n_258)
);

BUFx6f_ASAP7_75t_L g224 ( 
.A(n_143),
.Y(n_224)
);

CKINVDCx20_ASAP7_75t_R g254 ( 
.A(n_224),
.Y(n_254)
);

INVx5_ASAP7_75t_L g225 ( 
.A(n_151),
.Y(n_225)
);

CKINVDCx20_ASAP7_75t_R g266 ( 
.A(n_225),
.Y(n_266)
);

INVx3_ASAP7_75t_L g226 ( 
.A(n_140),
.Y(n_226)
);

CKINVDCx10_ASAP7_75t_R g267 ( 
.A(n_226),
.Y(n_267)
);

NAND2xp5_ASAP7_75t_SL g227 ( 
.A(n_160),
.B(n_138),
.Y(n_227)
);

OAI21xp5_ASAP7_75t_L g229 ( 
.A1(n_184),
.A2(n_138),
.B(n_176),
.Y(n_229)
);

AND2x2_ASAP7_75t_L g272 ( 
.A(n_229),
.B(n_230),
.Y(n_272)
);

MAJIxp5_ASAP7_75t_L g230 ( 
.A(n_189),
.B(n_191),
.C(n_202),
.Y(n_230)
);

INVxp67_ASAP7_75t_L g295 ( 
.A(n_231),
.Y(n_295)
);

AOI22xp33_ASAP7_75t_L g234 ( 
.A1(n_206),
.A2(n_208),
.B1(n_214),
.B2(n_221),
.Y(n_234)
);

OAI22xp5_ASAP7_75t_SL g277 ( 
.A1(n_234),
.A2(n_225),
.B1(n_175),
.B2(n_204),
.Y(n_277)
);

AOI22xp5_ASAP7_75t_SL g293 ( 
.A1(n_235),
.A2(n_261),
.B1(n_259),
.B2(n_243),
.Y(n_293)
);

AND2x6_ASAP7_75t_L g237 ( 
.A(n_198),
.B(n_179),
.Y(n_237)
);

NAND2xp5_ASAP7_75t_SL g276 ( 
.A(n_237),
.B(n_260),
.Y(n_276)
);

NOR2xp33_ASAP7_75t_L g246 ( 
.A(n_185),
.B(n_186),
.Y(n_246)
);

NOR2xp33_ASAP7_75t_SL g282 ( 
.A(n_246),
.B(n_249),
.Y(n_282)
);

MAJIxp5_ASAP7_75t_L g249 ( 
.A(n_188),
.B(n_207),
.C(n_223),
.Y(n_249)
);

MAJIxp5_ASAP7_75t_L g250 ( 
.A(n_188),
.B(n_198),
.C(n_199),
.Y(n_250)
);

NOR2xp33_ASAP7_75t_SL g287 ( 
.A(n_250),
.B(n_259),
.Y(n_287)
);

NAND2xp5_ASAP7_75t_L g274 ( 
.A(n_258),
.B(n_224),
.Y(n_274)
);

MAJIxp5_ASAP7_75t_SL g259 ( 
.A(n_220),
.B(n_192),
.C(n_218),
.Y(n_259)
);

MAJIxp5_ASAP7_75t_L g260 ( 
.A(n_193),
.B(n_200),
.C(n_187),
.Y(n_260)
);

NOR2xp33_ASAP7_75t_L g263 ( 
.A(n_226),
.B(n_215),
.Y(n_263)
);

NAND2xp5_ASAP7_75t_SL g284 ( 
.A(n_263),
.B(n_241),
.Y(n_284)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_251),
.Y(n_270)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_270),
.Y(n_321)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_251),
.Y(n_271)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_271),
.Y(n_324)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_256),
.Y(n_273)
);

NOR2xp33_ASAP7_75t_L g312 ( 
.A(n_273),
.B(n_278),
.Y(n_312)
);

NAND2xp5_ASAP7_75t_L g303 ( 
.A(n_274),
.B(n_281),
.Y(n_303)
);

AO22x1_ASAP7_75t_L g275 ( 
.A1(n_262),
.A2(n_192),
.B1(n_219),
.B2(n_220),
.Y(n_275)
);

OAI21xp5_ASAP7_75t_L g304 ( 
.A1(n_275),
.A2(n_235),
.B(n_233),
.Y(n_304)
);

INVxp67_ASAP7_75t_L g319 ( 
.A(n_277),
.Y(n_319)
);

CKINVDCx20_ASAP7_75t_R g278 ( 
.A(n_240),
.Y(n_278)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_256),
.Y(n_279)
);

NOR2xp33_ASAP7_75t_L g316 ( 
.A(n_279),
.B(n_280),
.Y(n_316)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_268),
.Y(n_280)
);

OAI22xp5_ASAP7_75t_SL g281 ( 
.A1(n_236),
.A2(n_248),
.B1(n_231),
.B2(n_229),
.Y(n_281)
);

INVx1_ASAP7_75t_SL g283 ( 
.A(n_267),
.Y(n_283)
);

NAND2xp5_ASAP7_75t_L g305 ( 
.A(n_283),
.B(n_288),
.Y(n_305)
);

INVxp33_ASAP7_75t_L g314 ( 
.A(n_284),
.Y(n_314)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_268),
.Y(n_285)
);

NAND2xp5_ASAP7_75t_SL g302 ( 
.A(n_285),
.B(n_286),
.Y(n_302)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_268),
.Y(n_286)
);

INVx1_ASAP7_75t_SL g288 ( 
.A(n_267),
.Y(n_288)
);

INVx1_ASAP7_75t_SL g289 ( 
.A(n_262),
.Y(n_289)
);

NAND2xp5_ASAP7_75t_L g307 ( 
.A(n_289),
.B(n_291),
.Y(n_307)
);

INVx5_ASAP7_75t_SL g290 ( 
.A(n_255),
.Y(n_290)
);

CKINVDCx16_ASAP7_75t_R g309 ( 
.A(n_290),
.Y(n_309)
);

CKINVDCx20_ASAP7_75t_R g291 ( 
.A(n_238),
.Y(n_291)
);

AOI22xp5_ASAP7_75t_L g292 ( 
.A1(n_248),
.A2(n_236),
.B1(n_239),
.B2(n_262),
.Y(n_292)
);

OAI22xp5_ASAP7_75t_L g308 ( 
.A1(n_292),
.A2(n_300),
.B1(n_260),
.B2(n_233),
.Y(n_308)
);

OAI21xp5_ASAP7_75t_SL g318 ( 
.A1(n_293),
.A2(n_301),
.B(n_245),
.Y(n_318)
);

NAND2xp5_ASAP7_75t_L g294 ( 
.A(n_228),
.B(n_230),
.Y(n_294)
);

NAND2xp5_ASAP7_75t_L g313 ( 
.A(n_294),
.B(n_296),
.Y(n_313)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_258),
.Y(n_296)
);

NAND2xp5_ASAP7_75t_L g297 ( 
.A(n_228),
.B(n_249),
.Y(n_297)
);

NAND2xp5_ASAP7_75t_L g320 ( 
.A(n_297),
.B(n_298),
.Y(n_320)
);

OAI22xp5_ASAP7_75t_SL g298 ( 
.A1(n_235),
.A2(n_237),
.B1(n_250),
.B2(n_252),
.Y(n_298)
);

NAND2xp5_ASAP7_75t_SL g299 ( 
.A(n_242),
.B(n_253),
.Y(n_299)
);

AOI221xp5_ASAP7_75t_L g315 ( 
.A1(n_299),
.A2(n_257),
.B1(n_245),
.B2(n_269),
.C(n_266),
.Y(n_315)
);

OAI22xp5_ASAP7_75t_SL g300 ( 
.A1(n_235),
.A2(n_254),
.B1(n_232),
.B2(n_247),
.Y(n_300)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_265),
.Y(n_301)
);

INVx1_ASAP7_75t_SL g342 ( 
.A(n_304),
.Y(n_342)
);

OAI21xp5_ASAP7_75t_L g306 ( 
.A1(n_295),
.A2(n_235),
.B(n_241),
.Y(n_306)
);

OAI21xp5_ASAP7_75t_SL g340 ( 
.A1(n_306),
.A2(n_318),
.B(n_280),
.Y(n_340)
);

NAND2xp5_ASAP7_75t_L g336 ( 
.A(n_308),
.B(n_311),
.Y(n_336)
);

MAJIxp5_ASAP7_75t_L g310 ( 
.A(n_272),
.B(n_265),
.C(n_269),
.Y(n_310)
);

MAJIxp5_ASAP7_75t_L g334 ( 
.A(n_310),
.B(n_317),
.C(n_272),
.Y(n_334)
);

OAI22xp5_ASAP7_75t_SL g311 ( 
.A1(n_292),
.A2(n_254),
.B1(n_247),
.B2(n_266),
.Y(n_311)
);

BUFx24_ASAP7_75t_SL g326 ( 
.A(n_315),
.Y(n_326)
);

XNOR2xp5_ASAP7_75t_L g317 ( 
.A(n_297),
.B(n_294),
.Y(n_317)
);

OAI22xp5_ASAP7_75t_SL g322 ( 
.A1(n_276),
.A2(n_244),
.B1(n_257),
.B2(n_264),
.Y(n_322)
);

NAND2xp5_ASAP7_75t_L g345 ( 
.A(n_322),
.B(n_277),
.Y(n_345)
);

OAI22xp5_ASAP7_75t_L g323 ( 
.A1(n_296),
.A2(n_244),
.B1(n_264),
.B2(n_255),
.Y(n_323)
);

AOI22xp33_ASAP7_75t_L g329 ( 
.A1(n_323),
.A2(n_319),
.B1(n_309),
.B2(n_288),
.Y(n_329)
);

AOI21xp5_ASAP7_75t_L g325 ( 
.A1(n_295),
.A2(n_255),
.B(n_281),
.Y(n_325)
);

AOI21xp5_ASAP7_75t_L g333 ( 
.A1(n_325),
.A2(n_289),
.B(n_300),
.Y(n_333)
);

XOR2xp5_ASAP7_75t_L g327 ( 
.A(n_317),
.B(n_272),
.Y(n_327)
);

MAJIxp5_ASAP7_75t_L g347 ( 
.A(n_327),
.B(n_341),
.C(n_310),
.Y(n_347)
);

NOR2xp33_ASAP7_75t_SL g328 ( 
.A(n_312),
.B(n_278),
.Y(n_328)
);

NOR2xp33_ASAP7_75t_L g361 ( 
.A(n_328),
.B(n_330),
.Y(n_361)
);

OAI22xp5_ASAP7_75t_SL g348 ( 
.A1(n_329),
.A2(n_335),
.B1(n_337),
.B2(n_343),
.Y(n_348)
);

NOR2xp33_ASAP7_75t_L g330 ( 
.A(n_317),
.B(n_291),
.Y(n_330)
);

NAND2xp5_ASAP7_75t_SL g331 ( 
.A(n_307),
.B(n_282),
.Y(n_331)
);

INVx1_ASAP7_75t_L g362 ( 
.A(n_331),
.Y(n_362)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_321),
.Y(n_332)
);

NAND2xp33_ASAP7_75t_SL g353 ( 
.A(n_332),
.B(n_333),
.Y(n_353)
);

XNOR2xp5_ASAP7_75t_L g346 ( 
.A(n_334),
.B(n_338),
.Y(n_346)
);

NOR2xp33_ASAP7_75t_L g335 ( 
.A(n_312),
.B(n_273),
.Y(n_335)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_321),
.Y(n_337)
);

OAI21xp33_ASAP7_75t_L g338 ( 
.A1(n_307),
.A2(n_287),
.B(n_298),
.Y(n_338)
);

MAJx2_ASAP7_75t_L g339 ( 
.A(n_320),
.B(n_293),
.C(n_279),
.Y(n_339)
);

XNOR2xp5_ASAP7_75t_L g358 ( 
.A(n_339),
.B(n_340),
.Y(n_358)
);

MAJIxp5_ASAP7_75t_L g341 ( 
.A(n_320),
.B(n_286),
.C(n_285),
.Y(n_341)
);

INVx1_ASAP7_75t_L g343 ( 
.A(n_324),
.Y(n_343)
);

INVx1_ASAP7_75t_L g344 ( 
.A(n_324),
.Y(n_344)
);

OAI22xp5_ASAP7_75t_SL g351 ( 
.A1(n_344),
.A2(n_345),
.B1(n_270),
.B2(n_271),
.Y(n_351)
);

XNOR2xp5_ASAP7_75t_L g365 ( 
.A(n_347),
.B(n_357),
.Y(n_365)
);

MAJIxp5_ASAP7_75t_L g349 ( 
.A(n_334),
.B(n_310),
.C(n_313),
.Y(n_349)
);

MAJIxp5_ASAP7_75t_L g363 ( 
.A(n_349),
.B(n_350),
.C(n_360),
.Y(n_363)
);

MAJIxp5_ASAP7_75t_L g350 ( 
.A(n_327),
.B(n_341),
.C(n_339),
.Y(n_350)
);

NAND2xp5_ASAP7_75t_L g371 ( 
.A(n_351),
.B(n_354),
.Y(n_371)
);

XNOR2x1_ASAP7_75t_L g352 ( 
.A(n_339),
.B(n_303),
.Y(n_352)
);

XOR2xp5_ASAP7_75t_L g372 ( 
.A(n_352),
.B(n_355),
.Y(n_372)
);

AOI22xp5_ASAP7_75t_L g354 ( 
.A1(n_336),
.A2(n_308),
.B1(n_322),
.B2(n_304),
.Y(n_354)
);

XOR2xp5_ASAP7_75t_L g355 ( 
.A(n_331),
.B(n_313),
.Y(n_355)
);

OA22x2_ASAP7_75t_L g356 ( 
.A1(n_342),
.A2(n_304),
.B1(n_314),
.B2(n_325),
.Y(n_356)
);

HB1xp67_ASAP7_75t_L g373 ( 
.A(n_356),
.Y(n_373)
);

XNOR2xp5_ASAP7_75t_SL g357 ( 
.A(n_326),
.B(n_303),
.Y(n_357)
);

OAI22xp5_ASAP7_75t_SL g359 ( 
.A1(n_345),
.A2(n_316),
.B1(n_302),
.B2(n_274),
.Y(n_359)
);

INVxp67_ASAP7_75t_L g364 ( 
.A(n_359),
.Y(n_364)
);

MAJIxp5_ASAP7_75t_L g360 ( 
.A(n_336),
.B(n_322),
.C(n_318),
.Y(n_360)
);

INVx1_ASAP7_75t_L g366 ( 
.A(n_362),
.Y(n_366)
);

INVx1_ASAP7_75t_L g376 ( 
.A(n_366),
.Y(n_376)
);

INVx1_ASAP7_75t_L g367 ( 
.A(n_348),
.Y(n_367)
);

NOR2xp33_ASAP7_75t_L g378 ( 
.A(n_367),
.B(n_374),
.Y(n_378)
);

MAJIxp5_ASAP7_75t_L g368 ( 
.A(n_347),
.B(n_302),
.C(n_342),
.Y(n_368)
);

MAJIxp5_ASAP7_75t_L g381 ( 
.A(n_368),
.B(n_350),
.C(n_346),
.Y(n_381)
);

NOR2xp33_ASAP7_75t_L g369 ( 
.A(n_361),
.B(n_328),
.Y(n_369)
);

NAND2xp5_ASAP7_75t_SL g380 ( 
.A(n_369),
.B(n_370),
.Y(n_380)
);

NAND2xp5_ASAP7_75t_L g370 ( 
.A(n_355),
.B(n_316),
.Y(n_370)
);

INVx1_ASAP7_75t_L g374 ( 
.A(n_353),
.Y(n_374)
);

INVx1_ASAP7_75t_L g375 ( 
.A(n_356),
.Y(n_375)
);

NOR2xp33_ASAP7_75t_L g382 ( 
.A(n_375),
.B(n_371),
.Y(n_382)
);

OAI21xp5_ASAP7_75t_SL g377 ( 
.A1(n_364),
.A2(n_333),
.B(n_354),
.Y(n_377)
);

NAND2xp5_ASAP7_75t_SL g389 ( 
.A(n_377),
.B(n_379),
.Y(n_389)
);

MAJIxp5_ASAP7_75t_L g379 ( 
.A(n_363),
.B(n_346),
.C(n_349),
.Y(n_379)
);

NOR2xp33_ASAP7_75t_L g386 ( 
.A(n_381),
.B(n_385),
.Y(n_386)
);

INVx1_ASAP7_75t_L g388 ( 
.A(n_382),
.Y(n_388)
);

MAJIxp5_ASAP7_75t_L g383 ( 
.A(n_363),
.B(n_360),
.C(n_358),
.Y(n_383)
);

MAJIxp5_ASAP7_75t_L g387 ( 
.A(n_383),
.B(n_384),
.C(n_365),
.Y(n_387)
);

XOR2xp5_ASAP7_75t_L g384 ( 
.A(n_368),
.B(n_358),
.Y(n_384)
);

OAI21xp5_ASAP7_75t_SL g385 ( 
.A1(n_364),
.A2(n_340),
.B(n_305),
.Y(n_385)
);

AND2x2_ASAP7_75t_L g399 ( 
.A(n_387),
.B(n_392),
.Y(n_399)
);

INVx1_ASAP7_75t_L g390 ( 
.A(n_376),
.Y(n_390)
);

INVx1_ASAP7_75t_L g396 ( 
.A(n_390),
.Y(n_396)
);

CKINVDCx5p33_ASAP7_75t_R g391 ( 
.A(n_378),
.Y(n_391)
);

NOR2xp33_ASAP7_75t_SL g395 ( 
.A(n_391),
.B(n_365),
.Y(n_395)
);

AOI22xp5_ASAP7_75t_L g392 ( 
.A1(n_380),
.A2(n_373),
.B1(n_371),
.B2(n_372),
.Y(n_392)
);

OAI22xp5_ASAP7_75t_SL g393 ( 
.A1(n_383),
.A2(n_356),
.B1(n_352),
.B2(n_306),
.Y(n_393)
);

XOR2xp5_ASAP7_75t_L g397 ( 
.A(n_393),
.B(n_372),
.Y(n_397)
);

AOI21xp5_ASAP7_75t_L g394 ( 
.A1(n_389),
.A2(n_381),
.B(n_384),
.Y(n_394)
);

AOI21xp5_ASAP7_75t_L g402 ( 
.A1(n_394),
.A2(n_395),
.B(n_398),
.Y(n_402)
);

NOR2xp33_ASAP7_75t_L g404 ( 
.A(n_397),
.B(n_387),
.Y(n_404)
);

OAI21xp5_ASAP7_75t_L g398 ( 
.A1(n_386),
.A2(n_311),
.B(n_306),
.Y(n_398)
);

HB1xp67_ASAP7_75t_L g400 ( 
.A(n_395),
.Y(n_400)
);

XNOR2xp5_ASAP7_75t_L g406 ( 
.A(n_400),
.B(n_401),
.Y(n_406)
);

NOR2xp33_ASAP7_75t_L g401 ( 
.A(n_399),
.B(n_388),
.Y(n_401)
);

NOR2xp33_ASAP7_75t_L g403 ( 
.A(n_396),
.B(n_391),
.Y(n_403)
);

OAI21xp5_ASAP7_75t_L g407 ( 
.A1(n_403),
.A2(n_390),
.B(n_392),
.Y(n_407)
);

INVxp67_ASAP7_75t_L g405 ( 
.A(n_404),
.Y(n_405)
);

OAI22xp5_ASAP7_75t_L g409 ( 
.A1(n_407),
.A2(n_315),
.B1(n_343),
.B2(n_344),
.Y(n_409)
);

FAx1_ASAP7_75t_SL g408 ( 
.A(n_406),
.B(n_393),
.CI(n_402),
.CON(n_408),
.SN(n_408)
);

NAND3xp33_ASAP7_75t_SL g410 ( 
.A(n_408),
.B(n_409),
.C(n_405),
.Y(n_410)
);

O2A1O1Ixp33_ASAP7_75t_SL g411 ( 
.A1(n_410),
.A2(n_408),
.B(n_357),
.C(n_337),
.Y(n_411)
);

XOR2xp5_ASAP7_75t_L g412 ( 
.A(n_411),
.B(n_408),
.Y(n_412)
);


endmodule