module fake_jpeg_8001_n_257 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_257);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_257;

wire n_159;
wire n_117;
wire n_253;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_84;
wire n_59;
wire n_98;
wire n_252;
wire n_251;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_223;
wire n_187;
wire n_57;
wire n_21;
wire n_234;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_24;
wire n_44;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_121;
wire n_99;
wire n_102;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_170;
wire n_162;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_216;
wire n_217;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

INVx1_ASAP7_75t_L g16 ( 
.A(n_3),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_7),
.Y(n_17)
);

INVx6_ASAP7_75t_L g18 ( 
.A(n_12),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_15),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_11),
.Y(n_20)
);

NOR2xp33_ASAP7_75t_L g21 ( 
.A(n_15),
.B(n_5),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_4),
.Y(n_22)
);

INVx1_ASAP7_75t_SL g23 ( 
.A(n_4),
.Y(n_23)
);

BUFx5_ASAP7_75t_L g24 ( 
.A(n_4),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_11),
.Y(n_25)
);

INVx1_ASAP7_75t_SL g26 ( 
.A(n_9),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_8),
.Y(n_27)
);

OR2x2_ASAP7_75t_L g28 ( 
.A(n_5),
.B(n_6),
.Y(n_28)
);

BUFx16f_ASAP7_75t_L g29 ( 
.A(n_12),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_10),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_10),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_2),
.Y(n_32)
);

INVx4_ASAP7_75t_L g33 ( 
.A(n_29),
.Y(n_33)
);

INVx1_ASAP7_75t_SL g54 ( 
.A(n_33),
.Y(n_54)
);

CKINVDCx16_ASAP7_75t_R g34 ( 
.A(n_24),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_L g45 ( 
.A(n_34),
.B(n_37),
.Y(n_45)
);

INVx2_ASAP7_75t_L g35 ( 
.A(n_29),
.Y(n_35)
);

HB1xp67_ASAP7_75t_L g59 ( 
.A(n_35),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_29),
.Y(n_36)
);

INVx6_ASAP7_75t_L g56 ( 
.A(n_36),
.Y(n_56)
);

INVx3_ASAP7_75t_L g37 ( 
.A(n_19),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_29),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_38),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_29),
.Y(n_39)
);

INVx2_ASAP7_75t_L g42 ( 
.A(n_39),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_24),
.Y(n_40)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_40),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g41 ( 
.A(n_28),
.B(n_15),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_41),
.B(n_28),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_L g43 ( 
.A(n_41),
.B(n_28),
.Y(n_43)
);

NAND2xp5_ASAP7_75t_L g74 ( 
.A(n_43),
.B(n_58),
.Y(n_74)
);

OR2x2_ASAP7_75t_L g44 ( 
.A(n_33),
.B(n_17),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_SL g62 ( 
.A(n_44),
.B(n_50),
.Y(n_62)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_37),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_47),
.B(n_52),
.Y(n_78)
);

AND2x2_ASAP7_75t_L g48 ( 
.A(n_35),
.B(n_24),
.Y(n_48)
);

AND2x2_ASAP7_75t_L g61 ( 
.A(n_48),
.B(n_53),
.Y(n_61)
);

AOI22xp5_ASAP7_75t_L g51 ( 
.A1(n_37),
.A2(n_18),
.B1(n_26),
.B2(n_23),
.Y(n_51)
);

OAI22xp5_ASAP7_75t_SL g80 ( 
.A1(n_51),
.A2(n_18),
.B1(n_23),
.B2(n_16),
.Y(n_80)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_35),
.Y(n_52)
);

NAND2xp33_ASAP7_75t_SL g53 ( 
.A(n_33),
.B(n_28),
.Y(n_53)
);

CKINVDCx20_ASAP7_75t_R g55 ( 
.A(n_36),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_SL g75 ( 
.A(n_55),
.B(n_57),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g57 ( 
.A(n_34),
.B(n_21),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_L g58 ( 
.A(n_36),
.B(n_26),
.Y(n_58)
);

BUFx5_ASAP7_75t_L g60 ( 
.A(n_54),
.Y(n_60)
);

INVx5_ASAP7_75t_L g100 ( 
.A(n_60),
.Y(n_100)
);

CKINVDCx14_ASAP7_75t_R g63 ( 
.A(n_45),
.Y(n_63)
);

AOI22xp33_ASAP7_75t_L g104 ( 
.A1(n_63),
.A2(n_56),
.B1(n_42),
.B2(n_20),
.Y(n_104)
);

INVxp67_ASAP7_75t_L g64 ( 
.A(n_45),
.Y(n_64)
);

INVxp67_ASAP7_75t_L g91 ( 
.A(n_64),
.Y(n_91)
);

CKINVDCx20_ASAP7_75t_R g65 ( 
.A(n_56),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_65),
.B(n_67),
.Y(n_92)
);

AOI22xp33_ASAP7_75t_SL g66 ( 
.A1(n_54),
.A2(n_18),
.B1(n_26),
.B2(n_23),
.Y(n_66)
);

AOI21xp5_ASAP7_75t_L g102 ( 
.A1(n_66),
.A2(n_84),
.B(n_87),
.Y(n_102)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_58),
.Y(n_67)
);

BUFx2_ASAP7_75t_SL g68 ( 
.A(n_49),
.Y(n_68)
);

BUFx2_ASAP7_75t_L g106 ( 
.A(n_68),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_SL g69 ( 
.A(n_43),
.B(n_50),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_L g109 ( 
.A(n_69),
.B(n_81),
.Y(n_109)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_51),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_70),
.B(n_71),
.Y(n_95)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_48),
.Y(n_71)
);

CKINVDCx16_ASAP7_75t_R g72 ( 
.A(n_48),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_72),
.B(n_73),
.Y(n_96)
);

INVxp67_ASAP7_75t_L g73 ( 
.A(n_57),
.Y(n_73)
);

BUFx6f_ASAP7_75t_L g76 ( 
.A(n_49),
.Y(n_76)
);

INVx3_ASAP7_75t_L g99 ( 
.A(n_76),
.Y(n_99)
);

OAI22xp5_ASAP7_75t_L g77 ( 
.A1(n_53),
.A2(n_18),
.B1(n_16),
.B2(n_25),
.Y(n_77)
);

OAI22xp5_ASAP7_75t_SL g114 ( 
.A1(n_77),
.A2(n_31),
.B1(n_27),
.B2(n_19),
.Y(n_114)
);

INVx2_ASAP7_75t_L g79 ( 
.A(n_59),
.Y(n_79)
);

CKINVDCx20_ASAP7_75t_R g101 ( 
.A(n_79),
.Y(n_101)
);

AOI22xp5_ASAP7_75t_L g111 ( 
.A1(n_80),
.A2(n_20),
.B1(n_22),
.B2(n_42),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_SL g81 ( 
.A(n_44),
.B(n_39),
.Y(n_81)
);

INVx2_ASAP7_75t_L g82 ( 
.A(n_59),
.Y(n_82)
);

CKINVDCx20_ASAP7_75t_R g108 ( 
.A(n_82),
.Y(n_108)
);

INVx13_ASAP7_75t_L g83 ( 
.A(n_54),
.Y(n_83)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_83),
.Y(n_89)
);

AOI22xp33_ASAP7_75t_SL g84 ( 
.A1(n_48),
.A2(n_16),
.B1(n_25),
.B2(n_30),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_SL g85 ( 
.A(n_44),
.B(n_21),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_L g110 ( 
.A(n_85),
.B(n_69),
.Y(n_110)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_47),
.Y(n_86)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_86),
.Y(n_93)
);

AOI22xp33_ASAP7_75t_SL g87 ( 
.A1(n_56),
.A2(n_25),
.B1(n_30),
.B2(n_17),
.Y(n_87)
);

AND2x2_ASAP7_75t_L g88 ( 
.A(n_52),
.B(n_0),
.Y(n_88)
);

MAJIxp5_ASAP7_75t_SL g103 ( 
.A(n_88),
.B(n_32),
.C(n_31),
.Y(n_103)
);

XNOR2xp5_ASAP7_75t_SL g90 ( 
.A(n_74),
.B(n_40),
.Y(n_90)
);

MAJx2_ASAP7_75t_L g121 ( 
.A(n_90),
.B(n_105),
.C(n_88),
.Y(n_121)
);

MAJIxp5_ASAP7_75t_L g94 ( 
.A(n_72),
.B(n_55),
.C(n_46),
.Y(n_94)
);

AND2x2_ASAP7_75t_L g140 ( 
.A(n_94),
.B(n_103),
.Y(n_140)
);

OAI21xp5_ASAP7_75t_L g97 ( 
.A1(n_81),
.A2(n_46),
.B(n_22),
.Y(n_97)
);

OAI21xp5_ASAP7_75t_L g135 ( 
.A1(n_97),
.A2(n_78),
.B(n_86),
.Y(n_135)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_78),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_98),
.B(n_104),
.Y(n_124)
);

XNOR2xp5_ASAP7_75t_SL g105 ( 
.A(n_74),
.B(n_40),
.Y(n_105)
);

AND2x2_ASAP7_75t_L g107 ( 
.A(n_71),
.B(n_0),
.Y(n_107)
);

AOI21xp5_ASAP7_75t_L g122 ( 
.A1(n_107),
.A2(n_88),
.B(n_75),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_L g126 ( 
.A(n_110),
.B(n_62),
.Y(n_126)
);

OAI22xp5_ASAP7_75t_SL g132 ( 
.A1(n_111),
.A2(n_113),
.B1(n_65),
.B2(n_83),
.Y(n_132)
);

O2A1O1Ixp33_ASAP7_75t_L g112 ( 
.A1(n_77),
.A2(n_40),
.B(n_36),
.C(n_39),
.Y(n_112)
);

AOI22xp5_ASAP7_75t_L g137 ( 
.A1(n_112),
.A2(n_114),
.B1(n_80),
.B2(n_68),
.Y(n_137)
);

OAI22xp5_ASAP7_75t_L g113 ( 
.A1(n_70),
.A2(n_67),
.B1(n_61),
.B2(n_63),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_L g115 ( 
.A(n_109),
.B(n_61),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_L g149 ( 
.A(n_115),
.B(n_120),
.Y(n_149)
);

CKINVDCx16_ASAP7_75t_R g116 ( 
.A(n_92),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_SL g162 ( 
.A(n_116),
.B(n_123),
.Y(n_162)
);

AOI22xp33_ASAP7_75t_SL g117 ( 
.A1(n_100),
.A2(n_98),
.B1(n_89),
.B2(n_83),
.Y(n_117)
);

OAI22xp5_ASAP7_75t_L g147 ( 
.A1(n_117),
.A2(n_137),
.B1(n_91),
.B2(n_99),
.Y(n_147)
);

INVx2_ASAP7_75t_L g118 ( 
.A(n_100),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_L g165 ( 
.A(n_118),
.B(n_125),
.Y(n_165)
);

A2O1A1Ixp33_ASAP7_75t_L g119 ( 
.A1(n_95),
.A2(n_61),
.B(n_62),
.C(n_85),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_SL g163 ( 
.A(n_119),
.B(n_126),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_L g120 ( 
.A(n_109),
.B(n_75),
.Y(n_120)
);

XNOR2xp5_ASAP7_75t_SL g154 ( 
.A(n_121),
.B(n_38),
.Y(n_154)
);

OAI21xp5_ASAP7_75t_L g143 ( 
.A1(n_122),
.A2(n_135),
.B(n_102),
.Y(n_143)
);

CKINVDCx16_ASAP7_75t_R g123 ( 
.A(n_106),
.Y(n_123)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_112),
.Y(n_125)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_93),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_L g156 ( 
.A(n_127),
.B(n_130),
.Y(n_156)
);

INVxp33_ASAP7_75t_L g128 ( 
.A(n_106),
.Y(n_128)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_128),
.Y(n_151)
);

BUFx3_ASAP7_75t_L g129 ( 
.A(n_106),
.Y(n_129)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_129),
.Y(n_152)
);

CKINVDCx20_ASAP7_75t_R g130 ( 
.A(n_97),
.Y(n_130)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_93),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g164 ( 
.A(n_131),
.B(n_134),
.Y(n_164)
);

AOI22xp5_ASAP7_75t_L g146 ( 
.A1(n_132),
.A2(n_91),
.B1(n_89),
.B2(n_105),
.Y(n_146)
);

INVx2_ASAP7_75t_L g133 ( 
.A(n_101),
.Y(n_133)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_133),
.Y(n_142)
);

INVxp67_ASAP7_75t_L g134 ( 
.A(n_96),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_L g136 ( 
.A(n_110),
.B(n_82),
.Y(n_136)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_136),
.Y(n_157)
);

AOI22xp5_ASAP7_75t_L g138 ( 
.A1(n_114),
.A2(n_79),
.B1(n_60),
.B2(n_19),
.Y(n_138)
);

OAI22xp5_ASAP7_75t_SL g145 ( 
.A1(n_138),
.A2(n_103),
.B1(n_111),
.B2(n_99),
.Y(n_145)
);

INVxp67_ASAP7_75t_L g139 ( 
.A(n_102),
.Y(n_139)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_139),
.Y(n_158)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_113),
.Y(n_141)
);

A2O1A1Ixp33_ASAP7_75t_SL g161 ( 
.A1(n_141),
.A2(n_32),
.B(n_31),
.C(n_27),
.Y(n_161)
);

OAI21xp5_ASAP7_75t_SL g175 ( 
.A1(n_143),
.A2(n_148),
.B(n_150),
.Y(n_175)
);

XOR2xp5_ASAP7_75t_L g144 ( 
.A(n_121),
.B(n_90),
.Y(n_144)
);

MAJIxp5_ASAP7_75t_L g180 ( 
.A(n_144),
.B(n_153),
.C(n_155),
.Y(n_180)
);

AOI22xp5_ASAP7_75t_L g173 ( 
.A1(n_145),
.A2(n_132),
.B1(n_167),
.B2(n_125),
.Y(n_173)
);

OAI22xp5_ASAP7_75t_L g184 ( 
.A1(n_146),
.A2(n_32),
.B1(n_27),
.B2(n_19),
.Y(n_184)
);

AOI221xp5_ASAP7_75t_L g187 ( 
.A1(n_147),
.A2(n_76),
.B1(n_2),
.B2(n_3),
.C(n_5),
.Y(n_187)
);

AOI21xp5_ASAP7_75t_L g148 ( 
.A1(n_139),
.A2(n_94),
.B(n_107),
.Y(n_148)
);

OAI21xp5_ASAP7_75t_L g150 ( 
.A1(n_130),
.A2(n_107),
.B(n_108),
.Y(n_150)
);

XOR2xp5_ASAP7_75t_L g153 ( 
.A(n_115),
.B(n_38),
.Y(n_153)
);

XNOR2xp5_ASAP7_75t_SL g181 ( 
.A(n_154),
.B(n_159),
.Y(n_181)
);

MAJIxp5_ASAP7_75t_L g155 ( 
.A(n_141),
.B(n_108),
.C(n_101),
.Y(n_155)
);

MAJIxp5_ASAP7_75t_L g159 ( 
.A(n_136),
.B(n_39),
.C(n_38),
.Y(n_159)
);

AOI21xp5_ASAP7_75t_L g160 ( 
.A1(n_140),
.A2(n_49),
.B(n_0),
.Y(n_160)
);

OAI21xp5_ASAP7_75t_L g171 ( 
.A1(n_160),
.A2(n_166),
.B(n_138),
.Y(n_171)
);

AOI22xp5_ASAP7_75t_SL g190 ( 
.A1(n_161),
.A2(n_1),
.B1(n_3),
.B2(n_6),
.Y(n_190)
);

OAI21xp5_ASAP7_75t_L g166 ( 
.A1(n_122),
.A2(n_32),
.B(n_31),
.Y(n_166)
);

XNOR2x1_ASAP7_75t_L g167 ( 
.A(n_140),
.B(n_27),
.Y(n_167)
);

OAI322xp33_ASAP7_75t_L g179 ( 
.A1(n_167),
.A2(n_120),
.A3(n_135),
.B1(n_131),
.B2(n_127),
.C1(n_137),
.C2(n_124),
.Y(n_179)
);

NOR2xp33_ASAP7_75t_SL g168 ( 
.A(n_119),
.B(n_10),
.Y(n_168)
);

OR2x2_ASAP7_75t_L g189 ( 
.A(n_168),
.B(n_1),
.Y(n_189)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_164),
.Y(n_169)
);

NOR2xp33_ASAP7_75t_L g198 ( 
.A(n_169),
.B(n_170),
.Y(n_198)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_164),
.Y(n_170)
);

XNOR2xp5_ASAP7_75t_L g205 ( 
.A(n_171),
.B(n_184),
.Y(n_205)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_165),
.Y(n_172)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_172),
.Y(n_193)
);

OAI22xp5_ASAP7_75t_SL g204 ( 
.A1(n_173),
.A2(n_185),
.B1(n_150),
.B2(n_161),
.Y(n_204)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_162),
.Y(n_174)
);

NOR2xp33_ASAP7_75t_SL g191 ( 
.A(n_174),
.B(n_176),
.Y(n_191)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_156),
.Y(n_176)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_156),
.Y(n_177)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_177),
.Y(n_203)
);

AOI21xp5_ASAP7_75t_L g178 ( 
.A1(n_158),
.A2(n_140),
.B(n_134),
.Y(n_178)
);

OAI22xp5_ASAP7_75t_L g192 ( 
.A1(n_178),
.A2(n_190),
.B1(n_160),
.B2(n_166),
.Y(n_192)
);

XNOR2xp5_ASAP7_75t_SL g208 ( 
.A(n_179),
.B(n_153),
.Y(n_208)
);

OAI22xp5_ASAP7_75t_SL g182 ( 
.A1(n_158),
.A2(n_133),
.B1(n_118),
.B2(n_129),
.Y(n_182)
);

AOI22xp5_ASAP7_75t_L g201 ( 
.A1(n_182),
.A2(n_187),
.B1(n_157),
.B2(n_161),
.Y(n_201)
);

INVxp67_ASAP7_75t_L g183 ( 
.A(n_155),
.Y(n_183)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_183),
.Y(n_194)
);

AOI22xp5_ASAP7_75t_L g185 ( 
.A1(n_145),
.A2(n_76),
.B1(n_0),
.B2(n_2),
.Y(n_185)
);

BUFx3_ASAP7_75t_L g186 ( 
.A(n_152),
.Y(n_186)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_186),
.Y(n_197)
);

CKINVDCx20_ASAP7_75t_R g188 ( 
.A(n_142),
.Y(n_188)
);

NOR4xp25_ASAP7_75t_L g200 ( 
.A(n_188),
.B(n_149),
.C(n_151),
.D(n_157),
.Y(n_200)
);

AOI21xp33_ASAP7_75t_L g196 ( 
.A1(n_189),
.A2(n_163),
.B(n_149),
.Y(n_196)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_192),
.Y(n_211)
);

XOR2xp5_ASAP7_75t_L g195 ( 
.A(n_180),
.B(n_144),
.Y(n_195)
);

MAJIxp5_ASAP7_75t_L g210 ( 
.A(n_195),
.B(n_181),
.C(n_175),
.Y(n_210)
);

NOR2xp33_ASAP7_75t_SL g213 ( 
.A(n_196),
.B(n_189),
.Y(n_213)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_182),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_L g214 ( 
.A(n_199),
.B(n_206),
.Y(n_214)
);

AND2x2_ASAP7_75t_L g218 ( 
.A(n_200),
.B(n_161),
.Y(n_218)
);

NOR2xp33_ASAP7_75t_L g221 ( 
.A(n_201),
.B(n_204),
.Y(n_221)
);

OAI22xp5_ASAP7_75t_L g202 ( 
.A1(n_185),
.A2(n_146),
.B1(n_143),
.B2(n_148),
.Y(n_202)
);

INVxp67_ASAP7_75t_L g212 ( 
.A(n_202),
.Y(n_212)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_169),
.Y(n_206)
);

OAI22xp5_ASAP7_75t_SL g207 ( 
.A1(n_173),
.A2(n_159),
.B1(n_142),
.B2(n_154),
.Y(n_207)
);

NAND2xp5_ASAP7_75t_SL g220 ( 
.A(n_207),
.B(n_205),
.Y(n_220)
);

XNOR2xp5_ASAP7_75t_L g219 ( 
.A(n_208),
.B(n_181),
.Y(n_219)
);

XNOR2xp5_ASAP7_75t_L g209 ( 
.A(n_208),
.B(n_180),
.Y(n_209)
);

XNOR2xp5_ASAP7_75t_L g229 ( 
.A(n_209),
.B(n_210),
.Y(n_229)
);

INVxp67_ASAP7_75t_L g222 ( 
.A(n_213),
.Y(n_222)
);

NAND2xp5_ASAP7_75t_L g215 ( 
.A(n_193),
.B(n_172),
.Y(n_215)
);

NAND2xp5_ASAP7_75t_L g231 ( 
.A(n_215),
.B(n_216),
.Y(n_231)
);

NAND2xp5_ASAP7_75t_L g216 ( 
.A(n_198),
.B(n_183),
.Y(n_216)
);

AOI22xp33_ASAP7_75t_SL g217 ( 
.A1(n_199),
.A2(n_190),
.B1(n_178),
.B2(n_161),
.Y(n_217)
);

OAI22xp5_ASAP7_75t_SL g223 ( 
.A1(n_217),
.A2(n_220),
.B1(n_201),
.B2(n_194),
.Y(n_223)
);

OR2x2_ASAP7_75t_L g227 ( 
.A(n_218),
.B(n_191),
.Y(n_227)
);

HB1xp67_ASAP7_75t_L g232 ( 
.A(n_219),
.Y(n_232)
);

XOR2xp5_ASAP7_75t_L g237 ( 
.A(n_223),
.B(n_195),
.Y(n_237)
);

INVxp67_ASAP7_75t_L g224 ( 
.A(n_214),
.Y(n_224)
);

NAND2xp5_ASAP7_75t_L g240 ( 
.A(n_224),
.B(n_227),
.Y(n_240)
);

AOI22xp33_ASAP7_75t_SL g225 ( 
.A1(n_211),
.A2(n_203),
.B1(n_206),
.B2(n_197),
.Y(n_225)
);

OAI22xp5_ASAP7_75t_L g234 ( 
.A1(n_225),
.A2(n_228),
.B1(n_197),
.B2(n_186),
.Y(n_234)
);

INVx6_ASAP7_75t_L g226 ( 
.A(n_218),
.Y(n_226)
);

NAND2xp5_ASAP7_75t_SL g238 ( 
.A(n_226),
.B(n_224),
.Y(n_238)
);

AOI22xp5_ASAP7_75t_L g228 ( 
.A1(n_212),
.A2(n_221),
.B1(n_204),
.B2(n_207),
.Y(n_228)
);

OAI22xp5_ASAP7_75t_L g230 ( 
.A1(n_212),
.A2(n_194),
.B1(n_171),
.B2(n_205),
.Y(n_230)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_230),
.Y(n_236)
);

AOI22xp5_ASAP7_75t_SL g233 ( 
.A1(n_226),
.A2(n_217),
.B1(n_175),
.B2(n_210),
.Y(n_233)
);

XNOR2xp5_ASAP7_75t_L g246 ( 
.A(n_233),
.B(n_7),
.Y(n_246)
);

AOI21xp5_ASAP7_75t_L g245 ( 
.A1(n_234),
.A2(n_238),
.B(n_6),
.Y(n_245)
);

NOR2xp33_ASAP7_75t_SL g235 ( 
.A(n_227),
.B(n_209),
.Y(n_235)
);

NAND2xp5_ASAP7_75t_L g241 ( 
.A(n_235),
.B(n_239),
.Y(n_241)
);

AND2x2_ASAP7_75t_L g244 ( 
.A(n_237),
.B(n_229),
.Y(n_244)
);

NOR2xp33_ASAP7_75t_L g239 ( 
.A(n_231),
.B(n_1),
.Y(n_239)
);

NAND2xp5_ASAP7_75t_L g242 ( 
.A(n_240),
.B(n_222),
.Y(n_242)
);

MAJIxp5_ASAP7_75t_L g250 ( 
.A(n_242),
.B(n_246),
.C(n_8),
.Y(n_250)
);

AOI21xp5_ASAP7_75t_SL g243 ( 
.A1(n_240),
.A2(n_225),
.B(n_232),
.Y(n_243)
);

OAI21xp5_ASAP7_75t_L g248 ( 
.A1(n_243),
.A2(n_245),
.B(n_7),
.Y(n_248)
);

A2O1A1O1Ixp25_ASAP7_75t_L g247 ( 
.A1(n_244),
.A2(n_233),
.B(n_237),
.C(n_236),
.D(n_11),
.Y(n_247)
);

AOI21xp5_ASAP7_75t_L g251 ( 
.A1(n_247),
.A2(n_248),
.B(n_249),
.Y(n_251)
);

AOI21x1_ASAP7_75t_SL g249 ( 
.A1(n_241),
.A2(n_14),
.B(n_9),
.Y(n_249)
);

NAND2xp5_ASAP7_75t_L g252 ( 
.A(n_250),
.B(n_8),
.Y(n_252)
);

AOI21xp5_ASAP7_75t_L g254 ( 
.A1(n_252),
.A2(n_253),
.B(n_12),
.Y(n_254)
);

NAND2xp5_ASAP7_75t_L g253 ( 
.A(n_250),
.B(n_9),
.Y(n_253)
);

AO21x1_ASAP7_75t_L g256 ( 
.A1(n_254),
.A2(n_255),
.B(n_13),
.Y(n_256)
);

OAI21xp5_ASAP7_75t_SL g255 ( 
.A1(n_251),
.A2(n_13),
.B(n_14),
.Y(n_255)
);

XOR2xp5_ASAP7_75t_L g257 ( 
.A(n_256),
.B(n_13),
.Y(n_257)
);


endmodule