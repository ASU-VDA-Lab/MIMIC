module fake_jpeg_23236_n_32 (n_3, n_2, n_1, n_0, n_4, n_5, n_32);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_5;

output n_32;

wire n_13;
wire n_21;
wire n_10;
wire n_23;
wire n_27;
wire n_6;
wire n_22;
wire n_14;
wire n_19;
wire n_18;
wire n_20;
wire n_30;
wire n_16;
wire n_24;
wire n_28;
wire n_26;
wire n_9;
wire n_11;
wire n_17;
wire n_25;
wire n_31;
wire n_29;
wire n_12;
wire n_8;
wire n_15;
wire n_7;

NOR2xp33_ASAP7_75t_SL g6 ( 
.A(n_5),
.B(n_4),
.Y(n_6)
);

INVx3_ASAP7_75t_L g7 ( 
.A(n_4),
.Y(n_7)
);

BUFx6f_ASAP7_75t_L g8 ( 
.A(n_0),
.Y(n_8)
);

INVx2_ASAP7_75t_L g9 ( 
.A(n_1),
.Y(n_9)
);

BUFx6f_ASAP7_75t_L g10 ( 
.A(n_2),
.Y(n_10)
);

INVx6_ASAP7_75t_L g11 ( 
.A(n_2),
.Y(n_11)
);

INVx6_ASAP7_75t_L g12 ( 
.A(n_3),
.Y(n_12)
);

NAND2xp5_ASAP7_75t_L g13 ( 
.A(n_10),
.B(n_0),
.Y(n_13)
);

XNOR2xp5_ASAP7_75t_L g19 ( 
.A(n_13),
.B(n_17),
.Y(n_19)
);

NAND2xp5_ASAP7_75t_L g14 ( 
.A(n_6),
.B(n_0),
.Y(n_14)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_14),
.Y(n_18)
);

NOR2xp33_ASAP7_75t_SL g15 ( 
.A(n_7),
.B(n_3),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_15),
.Y(n_20)
);

INVx3_ASAP7_75t_L g16 ( 
.A(n_11),
.Y(n_16)
);

INVx5_ASAP7_75t_L g21 ( 
.A(n_16),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g17 ( 
.A(n_11),
.Y(n_17)
);

INVx1_ASAP7_75t_SL g22 ( 
.A(n_21),
.Y(n_22)
);

OAI21xp5_ASAP7_75t_SL g25 ( 
.A1(n_22),
.A2(n_23),
.B(n_18),
.Y(n_25)
);

NOR2xp33_ASAP7_75t_L g23 ( 
.A(n_20),
.B(n_13),
.Y(n_23)
);

OAI22xp5_ASAP7_75t_L g24 ( 
.A1(n_18),
.A2(n_16),
.B1(n_12),
.B2(n_9),
.Y(n_24)
);

OAI22xp5_ASAP7_75t_SL g26 ( 
.A1(n_24),
.A2(n_12),
.B1(n_21),
.B2(n_10),
.Y(n_26)
);

FAx1_ASAP7_75t_SL g28 ( 
.A(n_25),
.B(n_19),
.CI(n_8),
.CON(n_28),
.SN(n_28)
);

AOI22xp5_ASAP7_75t_L g27 ( 
.A1(n_26),
.A2(n_22),
.B1(n_17),
.B2(n_8),
.Y(n_27)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_27),
.Y(n_29)
);

AOI21xp5_ASAP7_75t_SL g30 ( 
.A1(n_29),
.A2(n_28),
.B(n_19),
.Y(n_30)
);

O2A1O1Ixp33_ASAP7_75t_SL g31 ( 
.A1(n_30),
.A2(n_28),
.B(n_27),
.C(n_5),
.Y(n_31)
);

OAI221xp5_ASAP7_75t_L g32 ( 
.A1(n_31),
.A2(n_1),
.B1(n_28),
.B2(n_20),
.C(n_23),
.Y(n_32)
);


endmodule