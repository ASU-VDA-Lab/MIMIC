module fake_netlist_5_2058_n_2048 (n_137, n_168, n_164, n_191, n_91, n_82, n_122, n_142, n_176, n_10, n_140, n_24, n_124, n_86, n_136, n_146, n_182, n_143, n_83, n_132, n_61, n_90, n_127, n_75, n_101, n_180, n_184, n_65, n_78, n_74, n_144, n_114, n_57, n_96, n_37, n_189, n_165, n_111, n_108, n_129, n_31, n_13, n_66, n_98, n_177, n_60, n_155, n_152, n_16, n_43, n_107, n_0, n_58, n_9, n_69, n_18, n_116, n_42, n_22, n_1, n_45, n_117, n_46, n_21, n_94, n_113, n_38, n_123, n_139, n_105, n_80, n_4, n_179, n_125, n_35, n_167, n_128, n_73, n_17, n_92, n_19, n_149, n_120, n_135, n_30, n_156, n_5, n_33, n_126, n_14, n_84, n_23, n_130, n_157, n_29, n_79, n_131, n_151, n_47, n_173, n_192, n_25, n_53, n_160, n_188, n_190, n_8, n_158, n_44, n_40, n_34, n_100, n_62, n_138, n_148, n_71, n_154, n_109, n_112, n_85, n_159, n_163, n_95, n_119, n_183, n_185, n_175, n_169, n_59, n_26, n_133, n_55, n_99, n_2, n_181, n_3, n_49, n_20, n_6, n_39, n_54, n_147, n_178, n_12, n_67, n_121, n_36, n_76, n_87, n_150, n_162, n_27, n_170, n_64, n_77, n_102, n_106, n_161, n_81, n_118, n_28, n_89, n_70, n_115, n_68, n_93, n_72, n_174, n_186, n_134, n_187, n_32, n_41, n_104, n_172, n_103, n_56, n_51, n_63, n_97, n_141, n_166, n_11, n_171, n_153, n_7, n_15, n_145, n_48, n_50, n_52, n_88, n_110, n_2048);

input n_137;
input n_168;
input n_164;
input n_191;
input n_91;
input n_82;
input n_122;
input n_142;
input n_176;
input n_10;
input n_140;
input n_24;
input n_124;
input n_86;
input n_136;
input n_146;
input n_182;
input n_143;
input n_83;
input n_132;
input n_61;
input n_90;
input n_127;
input n_75;
input n_101;
input n_180;
input n_184;
input n_65;
input n_78;
input n_74;
input n_144;
input n_114;
input n_57;
input n_96;
input n_37;
input n_189;
input n_165;
input n_111;
input n_108;
input n_129;
input n_31;
input n_13;
input n_66;
input n_98;
input n_177;
input n_60;
input n_155;
input n_152;
input n_16;
input n_43;
input n_107;
input n_0;
input n_58;
input n_9;
input n_69;
input n_18;
input n_116;
input n_42;
input n_22;
input n_1;
input n_45;
input n_117;
input n_46;
input n_21;
input n_94;
input n_113;
input n_38;
input n_123;
input n_139;
input n_105;
input n_80;
input n_4;
input n_179;
input n_125;
input n_35;
input n_167;
input n_128;
input n_73;
input n_17;
input n_92;
input n_19;
input n_149;
input n_120;
input n_135;
input n_30;
input n_156;
input n_5;
input n_33;
input n_126;
input n_14;
input n_84;
input n_23;
input n_130;
input n_157;
input n_29;
input n_79;
input n_131;
input n_151;
input n_47;
input n_173;
input n_192;
input n_25;
input n_53;
input n_160;
input n_188;
input n_190;
input n_8;
input n_158;
input n_44;
input n_40;
input n_34;
input n_100;
input n_62;
input n_138;
input n_148;
input n_71;
input n_154;
input n_109;
input n_112;
input n_85;
input n_159;
input n_163;
input n_95;
input n_119;
input n_183;
input n_185;
input n_175;
input n_169;
input n_59;
input n_26;
input n_133;
input n_55;
input n_99;
input n_2;
input n_181;
input n_3;
input n_49;
input n_20;
input n_6;
input n_39;
input n_54;
input n_147;
input n_178;
input n_12;
input n_67;
input n_121;
input n_36;
input n_76;
input n_87;
input n_150;
input n_162;
input n_27;
input n_170;
input n_64;
input n_77;
input n_102;
input n_106;
input n_161;
input n_81;
input n_118;
input n_28;
input n_89;
input n_70;
input n_115;
input n_68;
input n_93;
input n_72;
input n_174;
input n_186;
input n_134;
input n_187;
input n_32;
input n_41;
input n_104;
input n_172;
input n_103;
input n_56;
input n_51;
input n_63;
input n_97;
input n_141;
input n_166;
input n_11;
input n_171;
input n_153;
input n_7;
input n_15;
input n_145;
input n_48;
input n_50;
input n_52;
input n_88;
input n_110;

output n_2048;

wire n_924;
wire n_1263;
wire n_977;
wire n_1378;
wire n_611;
wire n_1126;
wire n_1423;
wire n_1729;
wire n_1166;
wire n_1751;
wire n_469;
wire n_1508;
wire n_785;
wire n_549;
wire n_532;
wire n_1161;
wire n_1859;
wire n_1677;
wire n_1150;
wire n_226;
wire n_1780;
wire n_1488;
wire n_667;
wire n_790;
wire n_1055;
wire n_1501;
wire n_880;
wire n_544;
wire n_1007;
wire n_552;
wire n_1528;
wire n_1370;
wire n_1292;
wire n_1198;
wire n_1360;
wire n_1099;
wire n_956;
wire n_564;
wire n_423;
wire n_1738;
wire n_2021;
wire n_1021;
wire n_1960;
wire n_551;
wire n_1323;
wire n_1466;
wire n_688;
wire n_1695;
wire n_1353;
wire n_800;
wire n_1347;
wire n_1535;
wire n_1789;
wire n_1666;
wire n_671;
wire n_819;
wire n_1451;
wire n_1022;
wire n_915;
wire n_1545;
wire n_864;
wire n_859;
wire n_951;
wire n_1947;
wire n_1264;
wire n_447;
wire n_247;
wire n_2001;
wire n_1494;
wire n_292;
wire n_625;
wire n_854;
wire n_1462;
wire n_1799;
wire n_1580;
wire n_674;
wire n_417;
wire n_1939;
wire n_1806;
wire n_516;
wire n_933;
wire n_1152;
wire n_497;
wire n_1869;
wire n_1607;
wire n_1563;
wire n_606;
wire n_275;
wire n_2011;
wire n_877;
wire n_2024;
wire n_1696;
wire n_755;
wire n_1118;
wire n_1686;
wire n_947;
wire n_1285;
wire n_373;
wire n_307;
wire n_1860;
wire n_1359;
wire n_530;
wire n_1107;
wire n_1728;
wire n_556;
wire n_2031;
wire n_1230;
wire n_668;
wire n_375;
wire n_301;
wire n_1896;
wire n_929;
wire n_1124;
wire n_1818;
wire n_902;
wire n_1576;
wire n_1104;
wire n_1294;
wire n_659;
wire n_1705;
wire n_1257;
wire n_1182;
wire n_579;
wire n_1698;
wire n_1261;
wire n_938;
wire n_1098;
wire n_320;
wire n_1154;
wire n_1242;
wire n_1135;
wire n_406;
wire n_519;
wire n_1016;
wire n_1243;
wire n_546;
wire n_2047;
wire n_1280;
wire n_1845;
wire n_281;
wire n_240;
wire n_291;
wire n_231;
wire n_257;
wire n_731;
wire n_371;
wire n_1483;
wire n_1314;
wire n_1512;
wire n_709;
wire n_1490;
wire n_317;
wire n_1236;
wire n_1633;
wire n_569;
wire n_1778;
wire n_227;
wire n_920;
wire n_1289;
wire n_1517;
wire n_335;
wire n_1669;
wire n_370;
wire n_976;
wire n_1949;
wire n_343;
wire n_1449;
wire n_308;
wire n_1946;
wire n_1566;
wire n_2032;
wire n_297;
wire n_1078;
wire n_1670;
wire n_775;
wire n_219;
wire n_600;
wire n_1484;
wire n_1374;
wire n_1328;
wire n_223;
wire n_1948;
wire n_1984;
wire n_264;
wire n_1877;
wire n_1831;
wire n_1598;
wire n_1723;
wire n_955;
wire n_1850;
wire n_339;
wire n_1146;
wire n_882;
wire n_243;
wire n_1036;
wire n_1097;
wire n_1749;
wire n_347;
wire n_550;
wire n_696;
wire n_897;
wire n_215;
wire n_350;
wire n_196;
wire n_798;
wire n_646;
wire n_1428;
wire n_436;
wire n_1394;
wire n_1414;
wire n_1216;
wire n_290;
wire n_580;
wire n_1040;
wire n_1872;
wire n_1852;
wire n_578;
wire n_926;
wire n_344;
wire n_1218;
wire n_1931;
wire n_475;
wire n_422;
wire n_777;
wire n_1070;
wire n_1547;
wire n_1030;
wire n_1755;
wire n_415;
wire n_1071;
wire n_485;
wire n_1165;
wire n_1267;
wire n_1561;
wire n_496;
wire n_1801;
wire n_1391;
wire n_958;
wire n_1034;
wire n_670;
wire n_1513;
wire n_1600;
wire n_521;
wire n_845;
wire n_663;
wire n_1862;
wire n_673;
wire n_837;
wire n_1239;
wire n_528;
wire n_1796;
wire n_680;
wire n_1473;
wire n_1587;
wire n_395;
wire n_553;
wire n_901;
wire n_813;
wire n_1521;
wire n_1284;
wire n_1590;
wire n_214;
wire n_1748;
wire n_1672;
wire n_675;
wire n_888;
wire n_1880;
wire n_1167;
wire n_1626;
wire n_637;
wire n_1384;
wire n_1556;
wire n_446;
wire n_1863;
wire n_1064;
wire n_858;
wire n_923;
wire n_691;
wire n_1151;
wire n_881;
wire n_1405;
wire n_1706;
wire n_468;
wire n_213;
wire n_342;
wire n_464;
wire n_363;
wire n_1582;
wire n_197;
wire n_1069;
wire n_1784;
wire n_1075;
wire n_1836;
wire n_1450;
wire n_1322;
wire n_1471;
wire n_1986;
wire n_1750;
wire n_1459;
wire n_460;
wire n_889;
wire n_973;
wire n_1700;
wire n_477;
wire n_571;
wire n_1585;
wire n_461;
wire n_1971;
wire n_1599;
wire n_1211;
wire n_1197;
wire n_1523;
wire n_1950;
wire n_907;
wire n_1447;
wire n_1377;
wire n_989;
wire n_1039;
wire n_228;
wire n_283;
wire n_1403;
wire n_488;
wire n_736;
wire n_892;
wire n_1000;
wire n_1202;
wire n_1278;
wire n_1002;
wire n_1463;
wire n_1581;
wire n_310;
wire n_593;
wire n_748;
wire n_586;
wire n_1058;
wire n_1667;
wire n_838;
wire n_332;
wire n_1053;
wire n_1224;
wire n_349;
wire n_1926;
wire n_1248;
wire n_230;
wire n_1331;
wire n_953;
wire n_279;
wire n_1014;
wire n_1241;
wire n_289;
wire n_963;
wire n_1052;
wire n_954;
wire n_627;
wire n_1385;
wire n_440;
wire n_793;
wire n_478;
wire n_1819;
wire n_476;
wire n_1527;
wire n_2042;
wire n_534;
wire n_1882;
wire n_884;
wire n_345;
wire n_944;
wire n_1754;
wire n_1623;
wire n_1854;
wire n_1565;
wire n_1809;
wire n_1856;
wire n_647;
wire n_237;
wire n_407;
wire n_1072;
wire n_832;
wire n_857;
wire n_207;
wire n_561;
wire n_1319;
wire n_1825;
wire n_1951;
wire n_1883;
wire n_1906;
wire n_1712;
wire n_1387;
wire n_1532;
wire n_1027;
wire n_971;
wire n_1156;
wire n_326;
wire n_794;
wire n_404;
wire n_686;
wire n_847;
wire n_1393;
wire n_596;
wire n_1775;
wire n_2028;
wire n_1368;
wire n_558;
wire n_702;
wire n_1276;
wire n_822;
wire n_1412;
wire n_1709;
wire n_728;
wire n_266;
wire n_1162;
wire n_272;
wire n_1538;
wire n_1838;
wire n_1199;
wire n_1847;
wire n_1779;
wire n_352;
wire n_1884;
wire n_1038;
wire n_520;
wire n_1369;
wire n_409;
wire n_1841;
wire n_1660;
wire n_887;
wire n_1905;
wire n_300;
wire n_809;
wire n_870;
wire n_931;
wire n_599;
wire n_1711;
wire n_1662;
wire n_1891;
wire n_1481;
wire n_1942;
wire n_434;
wire n_1978;
wire n_1544;
wire n_868;
wire n_639;
wire n_914;
wire n_411;
wire n_414;
wire n_1629;
wire n_1293;
wire n_965;
wire n_1876;
wire n_1743;
wire n_935;
wire n_1175;
wire n_817;
wire n_360;
wire n_1479;
wire n_1810;
wire n_1888;
wire n_2009;
wire n_759;
wire n_1892;
wire n_806;
wire n_1997;
wire n_1766;
wire n_1477;
wire n_324;
wire n_1635;
wire n_1963;
wire n_1571;
wire n_1189;
wire n_1259;
wire n_1690;
wire n_706;
wire n_746;
wire n_1649;
wire n_747;
wire n_784;
wire n_1733;
wire n_1244;
wire n_431;
wire n_1194;
wire n_1925;
wire n_1815;
wire n_615;
wire n_851;
wire n_1759;
wire n_843;
wire n_1788;
wire n_523;
wire n_913;
wire n_1537;
wire n_705;
wire n_865;
wire n_678;
wire n_697;
wire n_1222;
wire n_1679;
wire n_776;
wire n_1798;
wire n_2022;
wire n_1790;
wire n_1415;
wire n_367;
wire n_452;
wire n_525;
wire n_1260;
wire n_1746;
wire n_1647;
wire n_1829;
wire n_1464;
wire n_649;
wire n_547;
wire n_1444;
wire n_1191;
wire n_1674;
wire n_1833;
wire n_1830;
wire n_1710;
wire n_284;
wire n_1128;
wire n_1734;
wire n_744;
wire n_629;
wire n_590;
wire n_1308;
wire n_1767;
wire n_254;
wire n_1680;
wire n_1233;
wire n_1615;
wire n_1529;
wire n_2005;
wire n_526;
wire n_1916;
wire n_372;
wire n_293;
wire n_677;
wire n_244;
wire n_1333;
wire n_1121;
wire n_433;
wire n_604;
wire n_368;
wire n_314;
wire n_2007;
wire n_949;
wire n_1443;
wire n_1008;
wire n_946;
wire n_1539;
wire n_1001;
wire n_1503;
wire n_498;
wire n_1468;
wire n_1559;
wire n_1765;
wire n_1866;
wire n_689;
wire n_738;
wire n_1624;
wire n_640;
wire n_1510;
wire n_252;
wire n_624;
wire n_1380;
wire n_1744;
wire n_1617;
wire n_295;
wire n_1010;
wire n_1994;
wire n_1231;
wire n_739;
wire n_1279;
wire n_1406;
wire n_1195;
wire n_1837;
wire n_1839;
wire n_610;
wire n_1760;
wire n_936;
wire n_568;
wire n_1500;
wire n_1090;
wire n_757;
wire n_633;
wire n_439;
wire n_1832;
wire n_259;
wire n_448;
wire n_1851;
wire n_758;
wire n_999;
wire n_2046;
wire n_1933;
wire n_1656;
wire n_1158;
wire n_2045;
wire n_1509;
wire n_1874;
wire n_2040;
wire n_563;
wire n_1987;
wire n_1145;
wire n_878;
wire n_524;
wire n_394;
wire n_204;
wire n_1678;
wire n_1049;
wire n_1153;
wire n_741;
wire n_1639;
wire n_1306;
wire n_1068;
wire n_1871;
wire n_1964;
wire n_331;
wire n_906;
wire n_1163;
wire n_2039;
wire n_1207;
wire n_919;
wire n_908;
wire n_724;
wire n_1781;
wire n_2035;
wire n_658;
wire n_1740;
wire n_1362;
wire n_1586;
wire n_456;
wire n_959;
wire n_535;
wire n_940;
wire n_1445;
wire n_1492;
wire n_1923;
wire n_1773;
wire n_592;
wire n_1169;
wire n_1596;
wire n_1692;
wire n_1017;
wire n_978;
wire n_1434;
wire n_1054;
wire n_1474;
wire n_1665;
wire n_1269;
wire n_1095;
wire n_1828;
wire n_1614;
wire n_267;
wire n_514;
wire n_457;
wire n_1079;
wire n_1045;
wire n_1208;
wire n_2038;
wire n_603;
wire n_1431;
wire n_484;
wire n_1593;
wire n_1033;
wire n_442;
wire n_636;
wire n_660;
wire n_1640;
wire n_1732;
wire n_1009;
wire n_1148;
wire n_750;
wire n_742;
wire n_2029;
wire n_995;
wire n_454;
wire n_1609;
wire n_374;
wire n_1989;
wire n_396;
wire n_1887;
wire n_1383;
wire n_1073;
wire n_255;
wire n_662;
wire n_459;
wire n_218;
wire n_962;
wire n_1215;
wire n_1171;
wire n_1578;
wire n_723;
wire n_1920;
wire n_1065;
wire n_1592;
wire n_1336;
wire n_1721;
wire n_1959;
wire n_1758;
wire n_1574;
wire n_473;
wire n_1921;
wire n_1309;
wire n_1878;
wire n_1426;
wire n_1043;
wire n_355;
wire n_486;
wire n_1800;
wire n_1548;
wire n_614;
wire n_337;
wire n_1421;
wire n_1286;
wire n_1177;
wire n_1355;
wire n_974;
wire n_727;
wire n_1159;
wire n_957;
wire n_773;
wire n_208;
wire n_743;
wire n_299;
wire n_303;
wire n_296;
wire n_613;
wire n_1119;
wire n_1240;
wire n_1820;
wire n_829;
wire n_1612;
wire n_1416;
wire n_1724;
wire n_361;
wire n_700;
wire n_1237;
wire n_573;
wire n_1420;
wire n_1132;
wire n_388;
wire n_1366;
wire n_1300;
wire n_1127;
wire n_761;
wire n_1785;
wire n_1568;
wire n_1006;
wire n_329;
wire n_274;
wire n_1270;
wire n_1664;
wire n_1486;
wire n_582;
wire n_1332;
wire n_1390;
wire n_2017;
wire n_1870;
wire n_309;
wire n_512;
wire n_1591;
wire n_2033;
wire n_322;
wire n_1682;
wire n_1980;
wire n_1249;
wire n_652;
wire n_1111;
wire n_1365;
wire n_1927;
wire n_1349;
wire n_1093;
wire n_288;
wire n_1031;
wire n_263;
wire n_609;
wire n_1041;
wire n_1265;
wire n_1909;
wire n_224;
wire n_1562;
wire n_383;
wire n_834;
wire n_765;
wire n_893;
wire n_1015;
wire n_1140;
wire n_891;
wire n_1651;
wire n_1965;
wire n_239;
wire n_630;
wire n_1902;
wire n_1941;
wire n_1913;
wire n_504;
wire n_1823;
wire n_511;
wire n_874;
wire n_358;
wire n_1101;
wire n_1106;
wire n_1456;
wire n_2015;
wire n_1875;
wire n_1982;
wire n_1304;
wire n_1324;
wire n_987;
wire n_1846;
wire n_261;
wire n_1885;
wire n_1455;
wire n_767;
wire n_993;
wire n_1903;
wire n_1407;
wire n_1551;
wire n_545;
wire n_441;
wire n_860;
wire n_450;
wire n_1805;
wire n_1816;
wire n_429;
wire n_948;
wire n_1217;
wire n_628;
wire n_365;
wire n_1849;
wire n_729;
wire n_1131;
wire n_1084;
wire n_1961;
wire n_970;
wire n_1935;
wire n_911;
wire n_1430;
wire n_513;
wire n_1094;
wire n_1354;
wire n_560;
wire n_1534;
wire n_340;
wire n_1351;
wire n_1044;
wire n_1205;
wire n_346;
wire n_1209;
wire n_1552;
wire n_495;
wire n_602;
wire n_574;
wire n_1435;
wire n_879;
wire n_623;
wire n_405;
wire n_824;
wire n_359;
wire n_1645;
wire n_490;
wire n_1327;
wire n_996;
wire n_921;
wire n_1684;
wire n_233;
wire n_1717;
wire n_572;
wire n_366;
wire n_815;
wire n_1795;
wire n_1821;
wire n_327;
wire n_1381;
wire n_1611;
wire n_1037;
wire n_1080;
wire n_1274;
wire n_1316;
wire n_1708;
wire n_426;
wire n_1438;
wire n_1082;
wire n_1840;
wire n_589;
wire n_716;
wire n_1630;
wire n_562;
wire n_1436;
wire n_1691;
wire n_952;
wire n_1229;
wire n_391;
wire n_701;
wire n_1437;
wire n_1023;
wire n_645;
wire n_539;
wire n_803;
wire n_1092;
wire n_238;
wire n_1776;
wire n_531;
wire n_1757;
wire n_890;
wire n_1897;
wire n_764;
wire n_1919;
wire n_1056;
wire n_1424;
wire n_960;
wire n_1893;
wire n_222;
wire n_1290;
wire n_1123;
wire n_1467;
wire n_1047;
wire n_634;
wire n_199;
wire n_1958;
wire n_1252;
wire n_348;
wire n_1382;
wire n_1029;
wire n_925;
wire n_1206;
wire n_424;
wire n_1311;
wire n_1519;
wire n_256;
wire n_950;
wire n_1553;
wire n_1811;
wire n_380;
wire n_419;
wire n_1346;
wire n_444;
wire n_1299;
wire n_1808;
wire n_1060;
wire n_1141;
wire n_316;
wire n_389;
wire n_418;
wire n_248;
wire n_912;
wire n_315;
wire n_968;
wire n_451;
wire n_619;
wire n_408;
wire n_1386;
wire n_1699;
wire n_376;
wire n_967;
wire n_1442;
wire n_1139;
wire n_515;
wire n_351;
wire n_885;
wire n_397;
wire n_1432;
wire n_1357;
wire n_483;
wire n_683;
wire n_1632;
wire n_1057;
wire n_1051;
wire n_1085;
wire n_1066;
wire n_721;
wire n_1157;
wire n_841;
wire n_1050;
wire n_802;
wire n_1954;
wire n_1608;
wire n_983;
wire n_1844;
wire n_280;
wire n_1305;
wire n_873;
wire n_1826;
wire n_378;
wire n_1112;
wire n_762;
wire n_1283;
wire n_1644;
wire n_690;
wire n_1974;
wire n_583;
wire n_302;
wire n_1343;
wire n_1203;
wire n_1631;
wire n_821;
wire n_1763;
wire n_1966;
wire n_1768;
wire n_321;
wire n_1179;
wire n_621;
wire n_753;
wire n_455;
wire n_1048;
wire n_1719;
wire n_1288;
wire n_212;
wire n_385;
wire n_507;
wire n_1560;
wire n_1605;
wire n_330;
wire n_1228;
wire n_972;
wire n_692;
wire n_2037;
wire n_1953;
wire n_1938;
wire n_820;
wire n_1200;
wire n_1911;
wire n_1301;
wire n_1363;
wire n_1668;
wire n_1185;
wire n_991;
wire n_828;
wire n_1967;
wire n_779;
wire n_576;
wire n_1143;
wire n_1579;
wire n_1329;
wire n_1312;
wire n_1439;
wire n_804;
wire n_537;
wire n_1688;
wire n_945;
wire n_492;
wire n_1504;
wire n_943;
wire n_341;
wire n_250;
wire n_992;
wire n_1932;
wire n_543;
wire n_260;
wire n_842;
wire n_650;
wire n_984;
wire n_694;
wire n_286;
wire n_1992;
wire n_1643;
wire n_883;
wire n_1983;
wire n_470;
wire n_449;
wire n_325;
wire n_1594;
wire n_1214;
wire n_1342;
wire n_1400;
wire n_900;
wire n_856;
wire n_1793;
wire n_1976;
wire n_918;
wire n_942;
wire n_1804;
wire n_1147;
wire n_1557;
wire n_1977;
wire n_1610;
wire n_1077;
wire n_1422;
wire n_540;
wire n_618;
wire n_896;
wire n_323;
wire n_195;
wire n_356;
wire n_894;
wire n_1636;
wire n_1730;
wire n_831;
wire n_964;
wire n_1373;
wire n_1350;
wire n_1511;
wire n_1865;
wire n_1470;
wire n_1096;
wire n_234;
wire n_1575;
wire n_1697;
wire n_1735;
wire n_833;
wire n_2020;
wire n_1646;
wire n_225;
wire n_1307;
wire n_1881;
wire n_988;
wire n_2043;
wire n_1940;
wire n_814;
wire n_1549;
wire n_1934;
wire n_1201;
wire n_1114;
wire n_655;
wire n_2025;
wire n_1616;
wire n_1446;
wire n_669;
wire n_472;
wire n_1458;
wire n_1176;
wire n_1472;
wire n_1807;
wire n_387;
wire n_1149;
wire n_398;
wire n_1671;
wire n_635;
wire n_763;
wire n_1020;
wire n_1062;
wire n_211;
wire n_1824;
wire n_1917;
wire n_1219;
wire n_1204;
wire n_1814;
wire n_1035;
wire n_287;
wire n_555;
wire n_783;
wire n_1848;
wire n_1928;
wire n_1188;
wire n_1722;
wire n_661;
wire n_1802;
wire n_849;
wire n_584;
wire n_681;
wire n_336;
wire n_1638;
wire n_1786;
wire n_430;
wire n_2002;
wire n_510;
wire n_216;
wire n_311;
wire n_830;
wire n_1296;
wire n_1413;
wire n_801;
wire n_241;
wire n_875;
wire n_357;
wire n_1110;
wire n_1655;
wire n_445;
wire n_749;
wire n_1895;
wire n_1134;
wire n_1358;
wire n_717;
wire n_939;
wire n_482;
wire n_1088;
wire n_588;
wire n_1173;
wire n_789;
wire n_1232;
wire n_1603;
wire n_734;
wire n_638;
wire n_866;
wire n_969;
wire n_1401;
wire n_1019;
wire n_1105;
wire n_249;
wire n_1998;
wire n_304;
wire n_1338;
wire n_577;
wire n_2016;
wire n_1522;
wire n_1687;
wire n_1637;
wire n_2034;
wire n_1419;
wire n_338;
wire n_1653;
wire n_693;
wire n_1506;
wire n_836;
wire n_990;
wire n_1886;
wire n_1389;
wire n_1894;
wire n_975;
wire n_1908;
wire n_1256;
wire n_1702;
wire n_567;
wire n_1465;
wire n_778;
wire n_1122;
wire n_306;
wire n_458;
wire n_770;
wire n_1375;
wire n_1102;
wire n_1843;
wire n_711;
wire n_1499;
wire n_1187;
wire n_1441;
wire n_1392;
wire n_1597;
wire n_1929;
wire n_1164;
wire n_1659;
wire n_1834;
wire n_489;
wire n_1174;
wire n_1371;
wire n_617;
wire n_1303;
wire n_1572;
wire n_1968;
wire n_876;
wire n_1516;
wire n_1190;
wire n_1736;
wire n_1685;
wire n_601;
wire n_917;
wire n_1714;
wire n_966;
wire n_253;
wire n_1116;
wire n_2000;
wire n_1661;
wire n_1212;
wire n_1541;
wire n_206;
wire n_217;
wire n_726;
wire n_982;
wire n_1573;
wire n_1453;
wire n_1731;
wire n_818;
wire n_1970;
wire n_861;
wire n_1713;
wire n_1183;
wire n_1658;
wire n_899;
wire n_1253;
wire n_210;
wire n_1737;
wire n_1904;
wire n_1993;
wire n_774;
wire n_1628;
wire n_1335;
wire n_1514;
wire n_1777;
wire n_1957;
wire n_1059;
wire n_1345;
wire n_1133;
wire n_1771;
wire n_1912;
wire n_1899;
wire n_557;
wire n_1410;
wire n_1005;
wire n_607;
wire n_1003;
wire n_679;
wire n_710;
wire n_527;
wire n_1168;
wire n_707;
wire n_937;
wire n_1427;
wire n_393;
wire n_487;
wire n_1584;
wire n_665;
wire n_1726;
wire n_1835;
wire n_1440;
wire n_421;
wire n_1988;
wire n_1853;
wire n_1356;
wire n_1787;
wire n_910;
wire n_1657;
wire n_768;
wire n_1475;
wire n_1302;
wire n_1774;
wire n_1725;
wire n_205;
wire n_1136;
wire n_1313;
wire n_1491;
wire n_754;
wire n_1496;
wire n_1125;
wire n_410;
wire n_708;
wire n_529;
wire n_1812;
wire n_735;
wire n_232;
wire n_1915;
wire n_1109;
wire n_895;
wire n_1310;
wire n_1803;
wire n_202;
wire n_427;
wire n_1399;
wire n_1543;
wire n_1991;
wire n_1979;
wire n_791;
wire n_732;
wire n_1533;
wire n_193;
wire n_808;
wire n_797;
wire n_1025;
wire n_1930;
wire n_1955;
wire n_500;
wire n_1067;
wire n_1720;
wire n_435;
wire n_2003;
wire n_766;
wire n_1457;
wire n_541;
wire n_538;
wire n_2008;
wire n_1117;
wire n_799;
wire n_687;
wire n_715;
wire n_1742;
wire n_1480;
wire n_1482;
wire n_1213;
wire n_1266;
wire n_536;
wire n_872;
wire n_2012;
wire n_594;
wire n_200;
wire n_1291;
wire n_1297;
wire n_1753;
wire n_1782;
wire n_1155;
wire n_1418;
wire n_1972;
wire n_1524;
wire n_1689;
wire n_1485;
wire n_1011;
wire n_1184;
wire n_985;
wire n_1855;
wire n_869;
wire n_810;
wire n_416;
wire n_827;
wire n_401;
wire n_1703;
wire n_1352;
wire n_626;
wire n_1650;
wire n_1144;
wire n_1137;
wire n_1570;
wire n_1170;
wire n_305;
wire n_2023;
wire n_676;
wire n_294;
wire n_318;
wire n_653;
wire n_642;
wire n_1602;
wire n_194;
wire n_855;
wire n_1178;
wire n_1461;
wire n_850;
wire n_684;
wire n_268;
wire n_664;
wire n_1999;
wire n_503;
wire n_235;
wire n_1372;
wire n_605;
wire n_1273;
wire n_1822;
wire n_353;
wire n_620;
wire n_643;
wire n_916;
wire n_1081;
wire n_493;
wire n_1235;
wire n_980;
wire n_703;
wire n_698;
wire n_1115;
wire n_1282;
wire n_1318;
wire n_1783;
wire n_780;
wire n_998;
wire n_1454;
wire n_467;
wire n_1227;
wire n_1531;
wire n_840;
wire n_1334;
wire n_1907;
wire n_501;
wire n_823;
wire n_245;
wire n_725;
wire n_1388;
wire n_1417;
wire n_1295;
wire n_672;
wire n_1985;
wire n_1898;
wire n_581;
wire n_382;
wire n_554;
wire n_1625;
wire n_898;
wire n_1762;
wire n_1013;
wire n_1452;
wire n_718;
wire n_265;
wire n_1120;
wire n_719;
wire n_443;
wire n_1791;
wire n_198;
wire n_1890;
wire n_1747;
wire n_714;
wire n_1683;
wire n_1817;
wire n_909;
wire n_1944;
wire n_1497;
wire n_1530;
wire n_997;
wire n_932;
wire n_612;
wire n_1409;
wire n_788;
wire n_1326;
wire n_1268;
wire n_559;
wire n_825;
wire n_1981;
wire n_508;
wire n_506;
wire n_1320;
wire n_1663;
wire n_737;
wire n_1718;
wire n_986;
wire n_509;
wire n_1317;
wire n_1518;
wire n_1715;
wire n_1281;
wire n_1952;
wire n_1192;
wire n_1024;
wire n_1063;
wire n_1889;
wire n_209;
wire n_1792;
wire n_1564;
wire n_1868;
wire n_1613;
wire n_733;
wire n_1489;
wire n_1922;
wire n_1376;
wire n_941;
wire n_981;
wire n_1569;
wire n_867;
wire n_587;
wire n_792;
wire n_756;
wire n_1429;
wire n_399;
wire n_1238;
wire n_548;
wire n_812;
wire n_298;
wire n_518;
wire n_505;
wire n_1772;
wire n_282;
wire n_752;
wire n_905;
wire n_1476;
wire n_1108;
wire n_782;
wire n_1100;
wire n_1861;
wire n_1395;
wire n_862;
wire n_1425;
wire n_760;
wire n_1901;
wire n_1900;
wire n_1620;
wire n_381;
wire n_220;
wire n_390;
wire n_1330;
wire n_1867;
wire n_1945;
wire n_481;
wire n_1675;
wire n_1924;
wire n_1727;
wire n_1554;
wire n_1745;
wire n_769;
wire n_2006;
wire n_1995;
wire n_1046;
wire n_271;
wire n_934;
wire n_1618;
wire n_826;
wire n_1813;
wire n_886;
wire n_2014;
wire n_1221;
wire n_654;
wire n_1172;
wire n_428;
wire n_379;
wire n_1341;
wire n_570;
wire n_1641;
wire n_1361;
wire n_1707;
wire n_853;
wire n_377;
wire n_751;
wire n_1973;
wire n_786;
wire n_1083;
wire n_1142;
wire n_1129;
wire n_392;
wire n_704;
wire n_787;
wire n_1770;
wire n_961;
wire n_1756;
wire n_771;
wire n_276;
wire n_1716;
wire n_1225;
wire n_1520;
wire n_522;
wire n_1287;
wire n_1262;
wire n_400;
wire n_930;
wire n_1873;
wire n_1411;
wire n_221;
wire n_622;
wire n_1962;
wire n_1577;
wire n_1087;
wire n_386;
wire n_994;
wire n_1701;
wire n_848;
wire n_1550;
wire n_1498;
wire n_1223;
wire n_1272;
wire n_682;
wire n_1567;
wire n_1247;
wire n_922;
wire n_816;
wire n_1648;
wire n_591;
wire n_1536;
wire n_1857;
wire n_1344;
wire n_2041;
wire n_313;
wire n_631;
wire n_479;
wire n_1246;
wire n_1339;
wire n_1478;
wire n_1797;
wire n_432;
wire n_1769;
wire n_839;
wire n_1210;
wire n_1364;
wire n_328;
wire n_1250;
wire n_369;
wire n_1842;
wire n_871;
wire n_685;
wire n_598;
wire n_928;
wire n_608;
wire n_1367;
wire n_1943;
wire n_1460;
wire n_772;
wire n_2018;
wire n_1555;
wire n_499;
wire n_1589;
wire n_517;
wire n_402;
wire n_413;
wire n_1086;
wire n_796;
wire n_1858;
wire n_1619;
wire n_236;
wire n_1502;
wire n_1469;
wire n_1012;
wire n_1396;
wire n_1348;
wire n_2030;
wire n_903;
wire n_1525;
wire n_1752;
wire n_740;
wire n_203;
wire n_384;
wire n_1404;
wire n_1794;
wire n_1315;
wire n_277;
wire n_1061;
wire n_1910;
wire n_333;
wire n_1298;
wire n_1652;
wire n_462;
wire n_1193;
wire n_1676;
wire n_1255;
wire n_258;
wire n_1113;
wire n_1226;
wire n_722;
wire n_1277;
wire n_844;
wire n_201;
wire n_471;
wire n_852;
wire n_1487;
wire n_1864;
wire n_1028;
wire n_1601;
wire n_781;
wire n_474;
wire n_542;
wire n_463;
wire n_1546;
wire n_595;
wire n_502;
wire n_466;
wire n_420;
wire n_1337;
wire n_1495;
wire n_632;
wire n_699;
wire n_979;
wire n_1515;
wire n_1627;
wire n_1245;
wire n_846;
wire n_1673;
wire n_465;
wire n_362;
wire n_1321;
wire n_1975;
wire n_273;
wire n_1937;
wire n_585;
wire n_1739;
wire n_270;
wire n_616;
wire n_1914;
wire n_745;
wire n_1654;
wire n_1103;
wire n_648;
wire n_1379;
wire n_312;
wire n_1076;
wire n_1091;
wire n_1408;
wire n_494;
wire n_1761;
wire n_641;
wire n_730;
wire n_2036;
wire n_1325;
wire n_1595;
wire n_354;
wire n_575;
wire n_480;
wire n_425;
wire n_795;
wire n_695;
wire n_656;
wire n_1606;
wire n_1220;
wire n_1694;
wire n_1540;
wire n_229;
wire n_1936;
wire n_1956;
wire n_437;
wire n_1642;
wire n_2027;
wire n_403;
wire n_453;
wire n_1130;
wire n_720;
wire n_1918;
wire n_1526;
wire n_863;
wire n_805;
wire n_1604;
wire n_1275;
wire n_1764;
wire n_712;
wire n_246;
wire n_1583;
wire n_1042;
wire n_1402;
wire n_269;
wire n_285;
wire n_412;
wire n_1493;
wire n_657;
wire n_644;
wire n_1741;
wire n_1160;
wire n_1397;
wire n_491;
wire n_1258;
wire n_1074;
wire n_2004;
wire n_1621;
wire n_251;
wire n_566;
wire n_565;
wire n_1448;
wire n_1507;
wire n_1398;
wire n_1879;
wire n_597;
wire n_1996;
wire n_1181;
wire n_1505;
wire n_1634;
wire n_1196;
wire n_2019;
wire n_651;
wire n_1340;
wire n_334;
wire n_811;
wire n_1558;
wire n_807;
wire n_835;
wire n_666;
wire n_262;
wire n_1433;
wire n_1704;
wire n_1254;
wire n_1026;
wire n_2026;
wire n_1969;
wire n_1234;
wire n_319;
wire n_364;
wire n_1138;
wire n_927;
wire n_1089;
wire n_2013;
wire n_1990;
wire n_2044;
wire n_1004;
wire n_1186;
wire n_242;
wire n_1032;
wire n_1681;
wire n_2010;
wire n_1018;
wire n_1693;
wire n_438;
wire n_713;
wire n_904;
wire n_1588;
wire n_1622;
wire n_1180;
wire n_1827;
wire n_1271;
wire n_533;
wire n_1542;
wire n_1251;
wire n_278;

INVx1_ASAP7_75t_L g193 ( 
.A(n_80),
.Y(n_193)
);

CKINVDCx5p33_ASAP7_75t_R g194 ( 
.A(n_147),
.Y(n_194)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_164),
.Y(n_195)
);

CKINVDCx5p33_ASAP7_75t_R g196 ( 
.A(n_43),
.Y(n_196)
);

INVx1_ASAP7_75t_SL g197 ( 
.A(n_100),
.Y(n_197)
);

CKINVDCx20_ASAP7_75t_R g198 ( 
.A(n_15),
.Y(n_198)
);

INVx2_ASAP7_75t_SL g199 ( 
.A(n_28),
.Y(n_199)
);

CKINVDCx5p33_ASAP7_75t_R g200 ( 
.A(n_7),
.Y(n_200)
);

CKINVDCx5p33_ASAP7_75t_R g201 ( 
.A(n_62),
.Y(n_201)
);

CKINVDCx5p33_ASAP7_75t_R g202 ( 
.A(n_8),
.Y(n_202)
);

CKINVDCx5p33_ASAP7_75t_R g203 ( 
.A(n_38),
.Y(n_203)
);

CKINVDCx5p33_ASAP7_75t_R g204 ( 
.A(n_69),
.Y(n_204)
);

CKINVDCx5p33_ASAP7_75t_R g205 ( 
.A(n_10),
.Y(n_205)
);

INVxp67_ASAP7_75t_L g206 ( 
.A(n_186),
.Y(n_206)
);

BUFx3_ASAP7_75t_L g207 ( 
.A(n_95),
.Y(n_207)
);

CKINVDCx5p33_ASAP7_75t_R g208 ( 
.A(n_136),
.Y(n_208)
);

CKINVDCx5p33_ASAP7_75t_R g209 ( 
.A(n_6),
.Y(n_209)
);

CKINVDCx5p33_ASAP7_75t_R g210 ( 
.A(n_179),
.Y(n_210)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_144),
.Y(n_211)
);

INVx1_ASAP7_75t_SL g212 ( 
.A(n_25),
.Y(n_212)
);

CKINVDCx5p33_ASAP7_75t_R g213 ( 
.A(n_54),
.Y(n_213)
);

CKINVDCx5p33_ASAP7_75t_R g214 ( 
.A(n_139),
.Y(n_214)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_97),
.Y(n_215)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_56),
.Y(n_216)
);

CKINVDCx20_ASAP7_75t_R g217 ( 
.A(n_86),
.Y(n_217)
);

CKINVDCx5p33_ASAP7_75t_R g218 ( 
.A(n_104),
.Y(n_218)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_84),
.Y(n_219)
);

CKINVDCx5p33_ASAP7_75t_R g220 ( 
.A(n_185),
.Y(n_220)
);

INVx1_ASAP7_75t_SL g221 ( 
.A(n_167),
.Y(n_221)
);

CKINVDCx5p33_ASAP7_75t_R g222 ( 
.A(n_156),
.Y(n_222)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_13),
.Y(n_223)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_85),
.Y(n_224)
);

INVx2_ASAP7_75t_SL g225 ( 
.A(n_159),
.Y(n_225)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_93),
.Y(n_226)
);

CKINVDCx5p33_ASAP7_75t_R g227 ( 
.A(n_162),
.Y(n_227)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_37),
.Y(n_228)
);

INVxp33_ASAP7_75t_SL g229 ( 
.A(n_103),
.Y(n_229)
);

CKINVDCx5p33_ASAP7_75t_R g230 ( 
.A(n_108),
.Y(n_230)
);

CKINVDCx5p33_ASAP7_75t_R g231 ( 
.A(n_68),
.Y(n_231)
);

CKINVDCx5p33_ASAP7_75t_R g232 ( 
.A(n_134),
.Y(n_232)
);

BUFx10_ASAP7_75t_L g233 ( 
.A(n_180),
.Y(n_233)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_20),
.Y(n_234)
);

CKINVDCx5p33_ASAP7_75t_R g235 ( 
.A(n_70),
.Y(n_235)
);

CKINVDCx5p33_ASAP7_75t_R g236 ( 
.A(n_25),
.Y(n_236)
);

CKINVDCx5p33_ASAP7_75t_R g237 ( 
.A(n_24),
.Y(n_237)
);

CKINVDCx5p33_ASAP7_75t_R g238 ( 
.A(n_110),
.Y(n_238)
);

CKINVDCx5p33_ASAP7_75t_R g239 ( 
.A(n_1),
.Y(n_239)
);

INVx2_ASAP7_75t_L g240 ( 
.A(n_172),
.Y(n_240)
);

CKINVDCx20_ASAP7_75t_R g241 ( 
.A(n_74),
.Y(n_241)
);

CKINVDCx5p33_ASAP7_75t_R g242 ( 
.A(n_99),
.Y(n_242)
);

CKINVDCx5p33_ASAP7_75t_R g243 ( 
.A(n_154),
.Y(n_243)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_5),
.Y(n_244)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_36),
.Y(n_245)
);

CKINVDCx5p33_ASAP7_75t_R g246 ( 
.A(n_8),
.Y(n_246)
);

CKINVDCx5p33_ASAP7_75t_R g247 ( 
.A(n_29),
.Y(n_247)
);

CKINVDCx5p33_ASAP7_75t_R g248 ( 
.A(n_61),
.Y(n_248)
);

INVx2_ASAP7_75t_L g249 ( 
.A(n_5),
.Y(n_249)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_46),
.Y(n_250)
);

CKINVDCx5p33_ASAP7_75t_R g251 ( 
.A(n_49),
.Y(n_251)
);

CKINVDCx5p33_ASAP7_75t_R g252 ( 
.A(n_133),
.Y(n_252)
);

CKINVDCx20_ASAP7_75t_R g253 ( 
.A(n_55),
.Y(n_253)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_168),
.Y(n_254)
);

CKINVDCx20_ASAP7_75t_R g255 ( 
.A(n_174),
.Y(n_255)
);

CKINVDCx5p33_ASAP7_75t_R g256 ( 
.A(n_40),
.Y(n_256)
);

CKINVDCx20_ASAP7_75t_R g257 ( 
.A(n_48),
.Y(n_257)
);

CKINVDCx5p33_ASAP7_75t_R g258 ( 
.A(n_96),
.Y(n_258)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_122),
.Y(n_259)
);

CKINVDCx5p33_ASAP7_75t_R g260 ( 
.A(n_10),
.Y(n_260)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_132),
.Y(n_261)
);

BUFx3_ASAP7_75t_L g262 ( 
.A(n_181),
.Y(n_262)
);

CKINVDCx5p33_ASAP7_75t_R g263 ( 
.A(n_115),
.Y(n_263)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_151),
.Y(n_264)
);

BUFx6f_ASAP7_75t_L g265 ( 
.A(n_119),
.Y(n_265)
);

CKINVDCx5p33_ASAP7_75t_R g266 ( 
.A(n_170),
.Y(n_266)
);

CKINVDCx5p33_ASAP7_75t_R g267 ( 
.A(n_42),
.Y(n_267)
);

BUFx3_ASAP7_75t_L g268 ( 
.A(n_163),
.Y(n_268)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_14),
.Y(n_269)
);

CKINVDCx5p33_ASAP7_75t_R g270 ( 
.A(n_55),
.Y(n_270)
);

HB1xp67_ASAP7_75t_L g271 ( 
.A(n_184),
.Y(n_271)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_37),
.Y(n_272)
);

CKINVDCx5p33_ASAP7_75t_R g273 ( 
.A(n_54),
.Y(n_273)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_43),
.Y(n_274)
);

BUFx2_ASAP7_75t_L g275 ( 
.A(n_106),
.Y(n_275)
);

CKINVDCx20_ASAP7_75t_R g276 ( 
.A(n_1),
.Y(n_276)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_140),
.Y(n_277)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_135),
.Y(n_278)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_44),
.Y(n_279)
);

CKINVDCx5p33_ASAP7_75t_R g280 ( 
.A(n_146),
.Y(n_280)
);

CKINVDCx5p33_ASAP7_75t_R g281 ( 
.A(n_130),
.Y(n_281)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_189),
.Y(n_282)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_176),
.Y(n_283)
);

CKINVDCx5p33_ASAP7_75t_R g284 ( 
.A(n_125),
.Y(n_284)
);

BUFx2_ASAP7_75t_SL g285 ( 
.A(n_145),
.Y(n_285)
);

CKINVDCx5p33_ASAP7_75t_R g286 ( 
.A(n_11),
.Y(n_286)
);

CKINVDCx20_ASAP7_75t_R g287 ( 
.A(n_129),
.Y(n_287)
);

CKINVDCx5p33_ASAP7_75t_R g288 ( 
.A(n_89),
.Y(n_288)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_35),
.Y(n_289)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_149),
.Y(n_290)
);

INVx2_ASAP7_75t_SL g291 ( 
.A(n_158),
.Y(n_291)
);

CKINVDCx5p33_ASAP7_75t_R g292 ( 
.A(n_68),
.Y(n_292)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_153),
.Y(n_293)
);

BUFx2_ASAP7_75t_L g294 ( 
.A(n_183),
.Y(n_294)
);

CKINVDCx5p33_ASAP7_75t_R g295 ( 
.A(n_35),
.Y(n_295)
);

HB1xp67_ASAP7_75t_L g296 ( 
.A(n_38),
.Y(n_296)
);

CKINVDCx5p33_ASAP7_75t_R g297 ( 
.A(n_31),
.Y(n_297)
);

CKINVDCx5p33_ASAP7_75t_R g298 ( 
.A(n_120),
.Y(n_298)
);

CKINVDCx5p33_ASAP7_75t_R g299 ( 
.A(n_138),
.Y(n_299)
);

CKINVDCx5p33_ASAP7_75t_R g300 ( 
.A(n_102),
.Y(n_300)
);

CKINVDCx20_ASAP7_75t_R g301 ( 
.A(n_82),
.Y(n_301)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_50),
.Y(n_302)
);

CKINVDCx5p33_ASAP7_75t_R g303 ( 
.A(n_150),
.Y(n_303)
);

CKINVDCx5p33_ASAP7_75t_R g304 ( 
.A(n_87),
.Y(n_304)
);

CKINVDCx5p33_ASAP7_75t_R g305 ( 
.A(n_141),
.Y(n_305)
);

CKINVDCx5p33_ASAP7_75t_R g306 ( 
.A(n_31),
.Y(n_306)
);

CKINVDCx5p33_ASAP7_75t_R g307 ( 
.A(n_4),
.Y(n_307)
);

CKINVDCx5p33_ASAP7_75t_R g308 ( 
.A(n_71),
.Y(n_308)
);

CKINVDCx5p33_ASAP7_75t_R g309 ( 
.A(n_190),
.Y(n_309)
);

CKINVDCx5p33_ASAP7_75t_R g310 ( 
.A(n_113),
.Y(n_310)
);

CKINVDCx5p33_ASAP7_75t_R g311 ( 
.A(n_7),
.Y(n_311)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_165),
.Y(n_312)
);

BUFx3_ASAP7_75t_L g313 ( 
.A(n_155),
.Y(n_313)
);

CKINVDCx5p33_ASAP7_75t_R g314 ( 
.A(n_45),
.Y(n_314)
);

BUFx6f_ASAP7_75t_L g315 ( 
.A(n_32),
.Y(n_315)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_26),
.Y(n_316)
);

BUFx6f_ASAP7_75t_L g317 ( 
.A(n_148),
.Y(n_317)
);

BUFx6f_ASAP7_75t_L g318 ( 
.A(n_175),
.Y(n_318)
);

INVx1_ASAP7_75t_SL g319 ( 
.A(n_45),
.Y(n_319)
);

CKINVDCx20_ASAP7_75t_R g320 ( 
.A(n_77),
.Y(n_320)
);

CKINVDCx5p33_ASAP7_75t_R g321 ( 
.A(n_91),
.Y(n_321)
);

CKINVDCx5p33_ASAP7_75t_R g322 ( 
.A(n_46),
.Y(n_322)
);

CKINVDCx5p33_ASAP7_75t_R g323 ( 
.A(n_30),
.Y(n_323)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_6),
.Y(n_324)
);

CKINVDCx5p33_ASAP7_75t_R g325 ( 
.A(n_40),
.Y(n_325)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_81),
.Y(n_326)
);

CKINVDCx20_ASAP7_75t_R g327 ( 
.A(n_101),
.Y(n_327)
);

CKINVDCx5p33_ASAP7_75t_R g328 ( 
.A(n_63),
.Y(n_328)
);

BUFx5_ASAP7_75t_L g329 ( 
.A(n_191),
.Y(n_329)
);

INVx2_ASAP7_75t_SL g330 ( 
.A(n_76),
.Y(n_330)
);

CKINVDCx5p33_ASAP7_75t_R g331 ( 
.A(n_13),
.Y(n_331)
);

CKINVDCx5p33_ASAP7_75t_R g332 ( 
.A(n_142),
.Y(n_332)
);

BUFx3_ASAP7_75t_L g333 ( 
.A(n_44),
.Y(n_333)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_36),
.Y(n_334)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_126),
.Y(n_335)
);

CKINVDCx5p33_ASAP7_75t_R g336 ( 
.A(n_105),
.Y(n_336)
);

CKINVDCx5p33_ASAP7_75t_R g337 ( 
.A(n_188),
.Y(n_337)
);

INVx1_ASAP7_75t_SL g338 ( 
.A(n_166),
.Y(n_338)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_17),
.Y(n_339)
);

BUFx10_ASAP7_75t_L g340 ( 
.A(n_98),
.Y(n_340)
);

CKINVDCx5p33_ASAP7_75t_R g341 ( 
.A(n_56),
.Y(n_341)
);

INVx1_ASAP7_75t_L g342 ( 
.A(n_15),
.Y(n_342)
);

CKINVDCx5p33_ASAP7_75t_R g343 ( 
.A(n_22),
.Y(n_343)
);

CKINVDCx5p33_ASAP7_75t_R g344 ( 
.A(n_26),
.Y(n_344)
);

INVx1_ASAP7_75t_L g345 ( 
.A(n_47),
.Y(n_345)
);

BUFx5_ASAP7_75t_L g346 ( 
.A(n_118),
.Y(n_346)
);

INVx2_ASAP7_75t_L g347 ( 
.A(n_0),
.Y(n_347)
);

CKINVDCx5p33_ASAP7_75t_R g348 ( 
.A(n_173),
.Y(n_348)
);

CKINVDCx5p33_ASAP7_75t_R g349 ( 
.A(n_29),
.Y(n_349)
);

INVx1_ASAP7_75t_L g350 ( 
.A(n_143),
.Y(n_350)
);

INVx1_ASAP7_75t_L g351 ( 
.A(n_39),
.Y(n_351)
);

INVx1_ASAP7_75t_L g352 ( 
.A(n_112),
.Y(n_352)
);

CKINVDCx5p33_ASAP7_75t_R g353 ( 
.A(n_27),
.Y(n_353)
);

BUFx3_ASAP7_75t_L g354 ( 
.A(n_72),
.Y(n_354)
);

BUFx10_ASAP7_75t_L g355 ( 
.A(n_78),
.Y(n_355)
);

CKINVDCx5p33_ASAP7_75t_R g356 ( 
.A(n_61),
.Y(n_356)
);

CKINVDCx20_ASAP7_75t_R g357 ( 
.A(n_24),
.Y(n_357)
);

INVx1_ASAP7_75t_L g358 ( 
.A(n_109),
.Y(n_358)
);

INVx1_ASAP7_75t_SL g359 ( 
.A(n_21),
.Y(n_359)
);

CKINVDCx5p33_ASAP7_75t_R g360 ( 
.A(n_19),
.Y(n_360)
);

BUFx10_ASAP7_75t_L g361 ( 
.A(n_47),
.Y(n_361)
);

CKINVDCx5p33_ASAP7_75t_R g362 ( 
.A(n_0),
.Y(n_362)
);

INVx1_ASAP7_75t_L g363 ( 
.A(n_60),
.Y(n_363)
);

CKINVDCx5p33_ASAP7_75t_R g364 ( 
.A(n_62),
.Y(n_364)
);

INVx1_ASAP7_75t_SL g365 ( 
.A(n_123),
.Y(n_365)
);

INVx1_ASAP7_75t_L g366 ( 
.A(n_94),
.Y(n_366)
);

CKINVDCx5p33_ASAP7_75t_R g367 ( 
.A(n_73),
.Y(n_367)
);

CKINVDCx5p33_ASAP7_75t_R g368 ( 
.A(n_65),
.Y(n_368)
);

INVx2_ASAP7_75t_L g369 ( 
.A(n_92),
.Y(n_369)
);

INVx4_ASAP7_75t_R g370 ( 
.A(n_111),
.Y(n_370)
);

INVx1_ASAP7_75t_L g371 ( 
.A(n_28),
.Y(n_371)
);

CKINVDCx20_ASAP7_75t_R g372 ( 
.A(n_11),
.Y(n_372)
);

CKINVDCx5p33_ASAP7_75t_R g373 ( 
.A(n_48),
.Y(n_373)
);

CKINVDCx20_ASAP7_75t_R g374 ( 
.A(n_117),
.Y(n_374)
);

CKINVDCx5p33_ASAP7_75t_R g375 ( 
.A(n_124),
.Y(n_375)
);

CKINVDCx5p33_ASAP7_75t_R g376 ( 
.A(n_2),
.Y(n_376)
);

CKINVDCx5p33_ASAP7_75t_R g377 ( 
.A(n_177),
.Y(n_377)
);

CKINVDCx20_ASAP7_75t_R g378 ( 
.A(n_60),
.Y(n_378)
);

CKINVDCx5p33_ASAP7_75t_R g379 ( 
.A(n_79),
.Y(n_379)
);

CKINVDCx5p33_ASAP7_75t_R g380 ( 
.A(n_127),
.Y(n_380)
);

INVx1_ASAP7_75t_L g381 ( 
.A(n_23),
.Y(n_381)
);

CKINVDCx5p33_ASAP7_75t_R g382 ( 
.A(n_116),
.Y(n_382)
);

CKINVDCx14_ASAP7_75t_R g383 ( 
.A(n_65),
.Y(n_383)
);

CKINVDCx5p33_ASAP7_75t_R g384 ( 
.A(n_2),
.Y(n_384)
);

CKINVDCx5p33_ASAP7_75t_R g385 ( 
.A(n_187),
.Y(n_385)
);

CKINVDCx5p33_ASAP7_75t_R g386 ( 
.A(n_66),
.Y(n_386)
);

INVx1_ASAP7_75t_L g387 ( 
.A(n_34),
.Y(n_387)
);

CKINVDCx14_ASAP7_75t_R g388 ( 
.A(n_32),
.Y(n_388)
);

CKINVDCx5p33_ASAP7_75t_R g389 ( 
.A(n_90),
.Y(n_389)
);

CKINVDCx20_ASAP7_75t_R g390 ( 
.A(n_27),
.Y(n_390)
);

CKINVDCx5p33_ASAP7_75t_R g391 ( 
.A(n_18),
.Y(n_391)
);

INVx1_ASAP7_75t_L g392 ( 
.A(n_315),
.Y(n_392)
);

INVx1_ASAP7_75t_L g393 ( 
.A(n_315),
.Y(n_393)
);

INVx1_ASAP7_75t_L g394 ( 
.A(n_315),
.Y(n_394)
);

INVx1_ASAP7_75t_L g395 ( 
.A(n_333),
.Y(n_395)
);

INVx1_ASAP7_75t_L g396 ( 
.A(n_333),
.Y(n_396)
);

INVx1_ASAP7_75t_L g397 ( 
.A(n_315),
.Y(n_397)
);

CKINVDCx20_ASAP7_75t_R g398 ( 
.A(n_217),
.Y(n_398)
);

CKINVDCx5p33_ASAP7_75t_R g399 ( 
.A(n_383),
.Y(n_399)
);

INVx1_ASAP7_75t_L g400 ( 
.A(n_315),
.Y(n_400)
);

INVxp33_ASAP7_75t_L g401 ( 
.A(n_296),
.Y(n_401)
);

INVx1_ASAP7_75t_L g402 ( 
.A(n_216),
.Y(n_402)
);

INVxp67_ASAP7_75t_SL g403 ( 
.A(n_271),
.Y(n_403)
);

INVx1_ASAP7_75t_L g404 ( 
.A(n_223),
.Y(n_404)
);

CKINVDCx5p33_ASAP7_75t_R g405 ( 
.A(n_388),
.Y(n_405)
);

INVxp67_ASAP7_75t_L g406 ( 
.A(n_361),
.Y(n_406)
);

INVx1_ASAP7_75t_L g407 ( 
.A(n_228),
.Y(n_407)
);

CKINVDCx5p33_ASAP7_75t_R g408 ( 
.A(n_231),
.Y(n_408)
);

CKINVDCx5p33_ASAP7_75t_R g409 ( 
.A(n_236),
.Y(n_409)
);

CKINVDCx20_ASAP7_75t_R g410 ( 
.A(n_241),
.Y(n_410)
);

INVx1_ASAP7_75t_L g411 ( 
.A(n_249),
.Y(n_411)
);

INVx1_ASAP7_75t_L g412 ( 
.A(n_249),
.Y(n_412)
);

INVx1_ASAP7_75t_L g413 ( 
.A(n_347),
.Y(n_413)
);

INVx1_ASAP7_75t_L g414 ( 
.A(n_347),
.Y(n_414)
);

INVx1_ASAP7_75t_L g415 ( 
.A(n_234),
.Y(n_415)
);

INVx1_ASAP7_75t_L g416 ( 
.A(n_244),
.Y(n_416)
);

BUFx3_ASAP7_75t_L g417 ( 
.A(n_207),
.Y(n_417)
);

CKINVDCx5p33_ASAP7_75t_R g418 ( 
.A(n_237),
.Y(n_418)
);

HB1xp67_ASAP7_75t_L g419 ( 
.A(n_196),
.Y(n_419)
);

INVx1_ASAP7_75t_L g420 ( 
.A(n_245),
.Y(n_420)
);

CKINVDCx5p33_ASAP7_75t_R g421 ( 
.A(n_239),
.Y(n_421)
);

CKINVDCx16_ASAP7_75t_R g422 ( 
.A(n_361),
.Y(n_422)
);

INVx1_ASAP7_75t_L g423 ( 
.A(n_250),
.Y(n_423)
);

CKINVDCx20_ASAP7_75t_R g424 ( 
.A(n_255),
.Y(n_424)
);

HB1xp67_ASAP7_75t_L g425 ( 
.A(n_196),
.Y(n_425)
);

INVxp33_ASAP7_75t_L g426 ( 
.A(n_269),
.Y(n_426)
);

INVx2_ASAP7_75t_L g427 ( 
.A(n_329),
.Y(n_427)
);

INVxp67_ASAP7_75t_L g428 ( 
.A(n_361),
.Y(n_428)
);

CKINVDCx5p33_ASAP7_75t_R g429 ( 
.A(n_246),
.Y(n_429)
);

CKINVDCx20_ASAP7_75t_R g430 ( 
.A(n_287),
.Y(n_430)
);

INVx1_ASAP7_75t_L g431 ( 
.A(n_272),
.Y(n_431)
);

INVx1_ASAP7_75t_L g432 ( 
.A(n_274),
.Y(n_432)
);

CKINVDCx20_ASAP7_75t_R g433 ( 
.A(n_301),
.Y(n_433)
);

INVx1_ASAP7_75t_L g434 ( 
.A(n_279),
.Y(n_434)
);

INVx2_ASAP7_75t_L g435 ( 
.A(n_329),
.Y(n_435)
);

INVx2_ASAP7_75t_L g436 ( 
.A(n_329),
.Y(n_436)
);

CKINVDCx5p33_ASAP7_75t_R g437 ( 
.A(n_247),
.Y(n_437)
);

INVx1_ASAP7_75t_L g438 ( 
.A(n_289),
.Y(n_438)
);

INVxp67_ASAP7_75t_SL g439 ( 
.A(n_275),
.Y(n_439)
);

CKINVDCx5p33_ASAP7_75t_R g440 ( 
.A(n_248),
.Y(n_440)
);

CKINVDCx5p33_ASAP7_75t_R g441 ( 
.A(n_251),
.Y(n_441)
);

HB1xp67_ASAP7_75t_L g442 ( 
.A(n_200),
.Y(n_442)
);

BUFx6f_ASAP7_75t_L g443 ( 
.A(n_265),
.Y(n_443)
);

INVx1_ASAP7_75t_L g444 ( 
.A(n_302),
.Y(n_444)
);

INVx1_ASAP7_75t_L g445 ( 
.A(n_316),
.Y(n_445)
);

INVx1_ASAP7_75t_L g446 ( 
.A(n_324),
.Y(n_446)
);

INVx1_ASAP7_75t_L g447 ( 
.A(n_334),
.Y(n_447)
);

INVx1_ASAP7_75t_L g448 ( 
.A(n_339),
.Y(n_448)
);

INVx1_ASAP7_75t_L g449 ( 
.A(n_342),
.Y(n_449)
);

INVx1_ASAP7_75t_L g450 ( 
.A(n_345),
.Y(n_450)
);

BUFx6f_ASAP7_75t_L g451 ( 
.A(n_265),
.Y(n_451)
);

INVx1_ASAP7_75t_L g452 ( 
.A(n_351),
.Y(n_452)
);

INVx1_ASAP7_75t_L g453 ( 
.A(n_363),
.Y(n_453)
);

BUFx6f_ASAP7_75t_L g454 ( 
.A(n_265),
.Y(n_454)
);

INVx1_ASAP7_75t_L g455 ( 
.A(n_371),
.Y(n_455)
);

CKINVDCx5p33_ASAP7_75t_R g456 ( 
.A(n_256),
.Y(n_456)
);

CKINVDCx20_ASAP7_75t_R g457 ( 
.A(n_320),
.Y(n_457)
);

INVxp33_ASAP7_75t_SL g458 ( 
.A(n_200),
.Y(n_458)
);

INVxp33_ASAP7_75t_SL g459 ( 
.A(n_201),
.Y(n_459)
);

INVxp67_ASAP7_75t_L g460 ( 
.A(n_381),
.Y(n_460)
);

INVx1_ASAP7_75t_L g461 ( 
.A(n_387),
.Y(n_461)
);

INVx1_ASAP7_75t_L g462 ( 
.A(n_207),
.Y(n_462)
);

INVx1_ASAP7_75t_L g463 ( 
.A(n_262),
.Y(n_463)
);

INVxp33_ASAP7_75t_SL g464 ( 
.A(n_201),
.Y(n_464)
);

CKINVDCx20_ASAP7_75t_R g465 ( 
.A(n_327),
.Y(n_465)
);

INVx1_ASAP7_75t_L g466 ( 
.A(n_262),
.Y(n_466)
);

INVx1_ASAP7_75t_L g467 ( 
.A(n_268),
.Y(n_467)
);

HB1xp67_ASAP7_75t_L g468 ( 
.A(n_202),
.Y(n_468)
);

CKINVDCx16_ASAP7_75t_R g469 ( 
.A(n_374),
.Y(n_469)
);

CKINVDCx20_ASAP7_75t_R g470 ( 
.A(n_230),
.Y(n_470)
);

INVx1_ASAP7_75t_L g471 ( 
.A(n_268),
.Y(n_471)
);

INVx1_ASAP7_75t_L g472 ( 
.A(n_313),
.Y(n_472)
);

INVxp33_ASAP7_75t_SL g473 ( 
.A(n_202),
.Y(n_473)
);

INVx1_ASAP7_75t_L g474 ( 
.A(n_313),
.Y(n_474)
);

INVx1_ASAP7_75t_L g475 ( 
.A(n_354),
.Y(n_475)
);

CKINVDCx16_ASAP7_75t_R g476 ( 
.A(n_233),
.Y(n_476)
);

CKINVDCx20_ASAP7_75t_R g477 ( 
.A(n_232),
.Y(n_477)
);

CKINVDCx5p33_ASAP7_75t_R g478 ( 
.A(n_260),
.Y(n_478)
);

INVx2_ASAP7_75t_L g479 ( 
.A(n_329),
.Y(n_479)
);

INVxp67_ASAP7_75t_SL g480 ( 
.A(n_294),
.Y(n_480)
);

INVxp67_ASAP7_75t_SL g481 ( 
.A(n_354),
.Y(n_481)
);

CKINVDCx5p33_ASAP7_75t_R g482 ( 
.A(n_267),
.Y(n_482)
);

CKINVDCx20_ASAP7_75t_R g483 ( 
.A(n_235),
.Y(n_483)
);

CKINVDCx20_ASAP7_75t_R g484 ( 
.A(n_238),
.Y(n_484)
);

INVxp67_ASAP7_75t_L g485 ( 
.A(n_203),
.Y(n_485)
);

INVx1_ASAP7_75t_L g486 ( 
.A(n_199),
.Y(n_486)
);

CKINVDCx5p33_ASAP7_75t_R g487 ( 
.A(n_270),
.Y(n_487)
);

CKINVDCx5p33_ASAP7_75t_R g488 ( 
.A(n_273),
.Y(n_488)
);

INVxp67_ASAP7_75t_SL g489 ( 
.A(n_206),
.Y(n_489)
);

CKINVDCx16_ASAP7_75t_R g490 ( 
.A(n_233),
.Y(n_490)
);

BUFx2_ASAP7_75t_L g491 ( 
.A(n_203),
.Y(n_491)
);

CKINVDCx20_ASAP7_75t_R g492 ( 
.A(n_242),
.Y(n_492)
);

CKINVDCx20_ASAP7_75t_R g493 ( 
.A(n_243),
.Y(n_493)
);

CKINVDCx16_ASAP7_75t_R g494 ( 
.A(n_233),
.Y(n_494)
);

CKINVDCx20_ASAP7_75t_R g495 ( 
.A(n_252),
.Y(n_495)
);

INVx1_ASAP7_75t_L g496 ( 
.A(n_199),
.Y(n_496)
);

INVx1_ASAP7_75t_L g497 ( 
.A(n_240),
.Y(n_497)
);

INVx2_ASAP7_75t_L g498 ( 
.A(n_329),
.Y(n_498)
);

NAND2xp5_ASAP7_75t_L g499 ( 
.A(n_462),
.B(n_225),
.Y(n_499)
);

INVx2_ASAP7_75t_L g500 ( 
.A(n_443),
.Y(n_500)
);

BUFx8_ASAP7_75t_L g501 ( 
.A(n_491),
.Y(n_501)
);

INVx1_ASAP7_75t_L g502 ( 
.A(n_392),
.Y(n_502)
);

NAND2xp5_ASAP7_75t_L g503 ( 
.A(n_463),
.B(n_225),
.Y(n_503)
);

CKINVDCx5p33_ASAP7_75t_R g504 ( 
.A(n_470),
.Y(n_504)
);

INVx5_ASAP7_75t_L g505 ( 
.A(n_443),
.Y(n_505)
);

NAND2xp5_ASAP7_75t_SL g506 ( 
.A(n_399),
.B(n_340),
.Y(n_506)
);

INVx2_ASAP7_75t_L g507 ( 
.A(n_443),
.Y(n_507)
);

CKINVDCx5p33_ASAP7_75t_R g508 ( 
.A(n_477),
.Y(n_508)
);

AND2x4_ASAP7_75t_L g509 ( 
.A(n_392),
.B(n_291),
.Y(n_509)
);

INVx2_ASAP7_75t_L g510 ( 
.A(n_443),
.Y(n_510)
);

BUFx8_ASAP7_75t_L g511 ( 
.A(n_491),
.Y(n_511)
);

HB1xp67_ASAP7_75t_L g512 ( 
.A(n_419),
.Y(n_512)
);

BUFx2_ASAP7_75t_L g513 ( 
.A(n_399),
.Y(n_513)
);

AND2x6_ASAP7_75t_L g514 ( 
.A(n_443),
.B(n_265),
.Y(n_514)
);

HB1xp67_ASAP7_75t_L g515 ( 
.A(n_425),
.Y(n_515)
);

AND2x2_ASAP7_75t_L g516 ( 
.A(n_481),
.B(n_340),
.Y(n_516)
);

NAND2xp5_ASAP7_75t_SL g517 ( 
.A(n_405),
.B(n_340),
.Y(n_517)
);

INVx3_ASAP7_75t_L g518 ( 
.A(n_451),
.Y(n_518)
);

AND2x2_ASAP7_75t_L g519 ( 
.A(n_466),
.B(n_291),
.Y(n_519)
);

INVx2_ASAP7_75t_L g520 ( 
.A(n_451),
.Y(n_520)
);

CKINVDCx5p33_ASAP7_75t_R g521 ( 
.A(n_483),
.Y(n_521)
);

INVx1_ASAP7_75t_L g522 ( 
.A(n_393),
.Y(n_522)
);

CKINVDCx5p33_ASAP7_75t_R g523 ( 
.A(n_484),
.Y(n_523)
);

INVx1_ASAP7_75t_L g524 ( 
.A(n_393),
.Y(n_524)
);

AND2x2_ASAP7_75t_L g525 ( 
.A(n_467),
.B(n_330),
.Y(n_525)
);

AND2x4_ASAP7_75t_L g526 ( 
.A(n_394),
.B(n_330),
.Y(n_526)
);

BUFx3_ASAP7_75t_L g527 ( 
.A(n_417),
.Y(n_527)
);

INVx1_ASAP7_75t_L g528 ( 
.A(n_394),
.Y(n_528)
);

INVx1_ASAP7_75t_L g529 ( 
.A(n_397),
.Y(n_529)
);

AND2x2_ASAP7_75t_L g530 ( 
.A(n_471),
.B(n_240),
.Y(n_530)
);

INVx2_ASAP7_75t_L g531 ( 
.A(n_451),
.Y(n_531)
);

INVx4_ASAP7_75t_L g532 ( 
.A(n_451),
.Y(n_532)
);

CKINVDCx5p33_ASAP7_75t_R g533 ( 
.A(n_492),
.Y(n_533)
);

CKINVDCx5p33_ASAP7_75t_R g534 ( 
.A(n_493),
.Y(n_534)
);

AND2x4_ASAP7_75t_L g535 ( 
.A(n_400),
.B(n_369),
.Y(n_535)
);

NAND2xp5_ASAP7_75t_L g536 ( 
.A(n_472),
.B(n_474),
.Y(n_536)
);

INVx2_ASAP7_75t_L g537 ( 
.A(n_451),
.Y(n_537)
);

NOR2xp33_ASAP7_75t_L g538 ( 
.A(n_439),
.B(n_229),
.Y(n_538)
);

AND2x4_ASAP7_75t_L g539 ( 
.A(n_475),
.B(n_369),
.Y(n_539)
);

INVx1_ASAP7_75t_L g540 ( 
.A(n_497),
.Y(n_540)
);

INVx1_ASAP7_75t_L g541 ( 
.A(n_415),
.Y(n_541)
);

INVx2_ASAP7_75t_L g542 ( 
.A(n_454),
.Y(n_542)
);

NOR2xp33_ASAP7_75t_R g543 ( 
.A(n_495),
.B(n_258),
.Y(n_543)
);

INVx2_ASAP7_75t_L g544 ( 
.A(n_454),
.Y(n_544)
);

AOI22xp5_ASAP7_75t_L g545 ( 
.A1(n_403),
.A2(n_276),
.B1(n_390),
.B2(n_253),
.Y(n_545)
);

INVx2_ASAP7_75t_L g546 ( 
.A(n_454),
.Y(n_546)
);

AND2x2_ASAP7_75t_L g547 ( 
.A(n_417),
.B(n_355),
.Y(n_547)
);

INVx3_ASAP7_75t_L g548 ( 
.A(n_454),
.Y(n_548)
);

NAND2xp5_ASAP7_75t_L g549 ( 
.A(n_395),
.B(n_396),
.Y(n_549)
);

INVxp67_ASAP7_75t_L g550 ( 
.A(n_442),
.Y(n_550)
);

INVx1_ASAP7_75t_L g551 ( 
.A(n_415),
.Y(n_551)
);

INVx1_ASAP7_75t_L g552 ( 
.A(n_416),
.Y(n_552)
);

INVx1_ASAP7_75t_L g553 ( 
.A(n_416),
.Y(n_553)
);

OAI22xp5_ASAP7_75t_L g554 ( 
.A1(n_401),
.A2(n_198),
.B1(n_372),
.B2(n_357),
.Y(n_554)
);

INVx1_ASAP7_75t_L g555 ( 
.A(n_420),
.Y(n_555)
);

INVx2_ASAP7_75t_L g556 ( 
.A(n_454),
.Y(n_556)
);

INVx2_ASAP7_75t_L g557 ( 
.A(n_427),
.Y(n_557)
);

OA21x2_ASAP7_75t_L g558 ( 
.A1(n_427),
.A2(n_195),
.B(n_193),
.Y(n_558)
);

INVx1_ASAP7_75t_L g559 ( 
.A(n_420),
.Y(n_559)
);

INVx2_ASAP7_75t_L g560 ( 
.A(n_435),
.Y(n_560)
);

AND2x4_ASAP7_75t_L g561 ( 
.A(n_435),
.B(n_211),
.Y(n_561)
);

BUFx6f_ASAP7_75t_L g562 ( 
.A(n_436),
.Y(n_562)
);

INVx1_ASAP7_75t_L g563 ( 
.A(n_423),
.Y(n_563)
);

CKINVDCx5p33_ASAP7_75t_R g564 ( 
.A(n_408),
.Y(n_564)
);

AND2x4_ASAP7_75t_L g565 ( 
.A(n_436),
.B(n_215),
.Y(n_565)
);

OAI22xp5_ASAP7_75t_L g566 ( 
.A1(n_458),
.A2(n_378),
.B1(n_257),
.B2(n_319),
.Y(n_566)
);

INVx2_ASAP7_75t_L g567 ( 
.A(n_479),
.Y(n_567)
);

INVx2_ASAP7_75t_L g568 ( 
.A(n_479),
.Y(n_568)
);

INVx1_ASAP7_75t_L g569 ( 
.A(n_423),
.Y(n_569)
);

INVx1_ASAP7_75t_L g570 ( 
.A(n_411),
.Y(n_570)
);

INVxp33_ASAP7_75t_L g571 ( 
.A(n_468),
.Y(n_571)
);

HB1xp67_ASAP7_75t_L g572 ( 
.A(n_485),
.Y(n_572)
);

INVx1_ASAP7_75t_L g573 ( 
.A(n_411),
.Y(n_573)
);

NAND2xp5_ASAP7_75t_L g574 ( 
.A(n_489),
.B(n_194),
.Y(n_574)
);

INVx1_ASAP7_75t_L g575 ( 
.A(n_412),
.Y(n_575)
);

INVx1_ASAP7_75t_L g576 ( 
.A(n_412),
.Y(n_576)
);

NAND2xp5_ASAP7_75t_L g577 ( 
.A(n_402),
.B(n_194),
.Y(n_577)
);

HB1xp67_ASAP7_75t_L g578 ( 
.A(n_408),
.Y(n_578)
);

NAND2xp5_ASAP7_75t_SL g579 ( 
.A(n_405),
.B(n_355),
.Y(n_579)
);

INVx1_ASAP7_75t_L g580 ( 
.A(n_413),
.Y(n_580)
);

INVx1_ASAP7_75t_L g581 ( 
.A(n_413),
.Y(n_581)
);

NAND2xp5_ASAP7_75t_SL g582 ( 
.A(n_476),
.B(n_355),
.Y(n_582)
);

INVx2_ASAP7_75t_L g583 ( 
.A(n_557),
.Y(n_583)
);

INVx2_ASAP7_75t_L g584 ( 
.A(n_557),
.Y(n_584)
);

AND2x2_ASAP7_75t_L g585 ( 
.A(n_530),
.B(n_480),
.Y(n_585)
);

INVx2_ASAP7_75t_L g586 ( 
.A(n_557),
.Y(n_586)
);

INVx1_ASAP7_75t_L g587 ( 
.A(n_560),
.Y(n_587)
);

INVx2_ASAP7_75t_L g588 ( 
.A(n_560),
.Y(n_588)
);

BUFx3_ASAP7_75t_L g589 ( 
.A(n_527),
.Y(n_589)
);

INVx2_ASAP7_75t_L g590 ( 
.A(n_560),
.Y(n_590)
);

NOR2xp33_ASAP7_75t_L g591 ( 
.A(n_538),
.B(n_458),
.Y(n_591)
);

AOI22xp5_ASAP7_75t_L g592 ( 
.A1(n_566),
.A2(n_464),
.B1(n_473),
.B2(n_459),
.Y(n_592)
);

INVx2_ASAP7_75t_L g593 ( 
.A(n_567),
.Y(n_593)
);

INVx1_ASAP7_75t_L g594 ( 
.A(n_567),
.Y(n_594)
);

NAND2xp5_ASAP7_75t_SL g595 ( 
.A(n_543),
.B(n_490),
.Y(n_595)
);

INVx1_ASAP7_75t_L g596 ( 
.A(n_567),
.Y(n_596)
);

INVx1_ASAP7_75t_L g597 ( 
.A(n_568),
.Y(n_597)
);

INVx2_ASAP7_75t_L g598 ( 
.A(n_568),
.Y(n_598)
);

INVx1_ASAP7_75t_L g599 ( 
.A(n_568),
.Y(n_599)
);

INVx1_ASAP7_75t_L g600 ( 
.A(n_502),
.Y(n_600)
);

NAND3xp33_ASAP7_75t_L g601 ( 
.A(n_530),
.B(n_460),
.C(n_407),
.Y(n_601)
);

AOI22xp33_ASAP7_75t_SL g602 ( 
.A1(n_566),
.A2(n_494),
.B1(n_422),
.B2(n_464),
.Y(n_602)
);

INVx2_ASAP7_75t_L g603 ( 
.A(n_562),
.Y(n_603)
);

INVx2_ASAP7_75t_L g604 ( 
.A(n_562),
.Y(n_604)
);

INVx3_ASAP7_75t_L g605 ( 
.A(n_562),
.Y(n_605)
);

AND2x2_ASAP7_75t_L g606 ( 
.A(n_530),
.B(n_414),
.Y(n_606)
);

INVxp33_ASAP7_75t_SL g607 ( 
.A(n_504),
.Y(n_607)
);

INVx1_ASAP7_75t_L g608 ( 
.A(n_502),
.Y(n_608)
);

NAND2xp5_ASAP7_75t_L g609 ( 
.A(n_561),
.B(n_498),
.Y(n_609)
);

INVx1_ASAP7_75t_SL g610 ( 
.A(n_547),
.Y(n_610)
);

INVx2_ASAP7_75t_L g611 ( 
.A(n_562),
.Y(n_611)
);

INVx3_ASAP7_75t_L g612 ( 
.A(n_562),
.Y(n_612)
);

INVx3_ASAP7_75t_L g613 ( 
.A(n_562),
.Y(n_613)
);

INVx3_ASAP7_75t_L g614 ( 
.A(n_532),
.Y(n_614)
);

INVx1_ASAP7_75t_L g615 ( 
.A(n_522),
.Y(n_615)
);

INVx4_ASAP7_75t_L g616 ( 
.A(n_514),
.Y(n_616)
);

AOI22xp33_ASAP7_75t_L g617 ( 
.A1(n_539),
.A2(n_459),
.B1(n_473),
.B2(n_229),
.Y(n_617)
);

INVx5_ASAP7_75t_L g618 ( 
.A(n_514),
.Y(n_618)
);

INVx2_ASAP7_75t_L g619 ( 
.A(n_500),
.Y(n_619)
);

INVx1_ASAP7_75t_L g620 ( 
.A(n_522),
.Y(n_620)
);

NAND2xp5_ASAP7_75t_SL g621 ( 
.A(n_574),
.B(n_409),
.Y(n_621)
);

NAND3xp33_ASAP7_75t_SL g622 ( 
.A(n_545),
.B(n_359),
.C(n_212),
.Y(n_622)
);

BUFx3_ASAP7_75t_L g623 ( 
.A(n_527),
.Y(n_623)
);

INVx1_ASAP7_75t_L g624 ( 
.A(n_524),
.Y(n_624)
);

AND3x2_ASAP7_75t_L g625 ( 
.A(n_513),
.B(n_428),
.C(n_406),
.Y(n_625)
);

INVx1_ASAP7_75t_L g626 ( 
.A(n_524),
.Y(n_626)
);

NAND2xp33_ASAP7_75t_SL g627 ( 
.A(n_571),
.B(n_409),
.Y(n_627)
);

INVx2_ASAP7_75t_L g628 ( 
.A(n_500),
.Y(n_628)
);

BUFx10_ASAP7_75t_L g629 ( 
.A(n_564),
.Y(n_629)
);

INVx2_ASAP7_75t_L g630 ( 
.A(n_500),
.Y(n_630)
);

INVx1_ASAP7_75t_L g631 ( 
.A(n_528),
.Y(n_631)
);

INVx2_ASAP7_75t_L g632 ( 
.A(n_507),
.Y(n_632)
);

NOR2xp33_ASAP7_75t_L g633 ( 
.A(n_574),
.B(n_418),
.Y(n_633)
);

INVx2_ASAP7_75t_L g634 ( 
.A(n_507),
.Y(n_634)
);

INVx3_ASAP7_75t_L g635 ( 
.A(n_532),
.Y(n_635)
);

INVx2_ASAP7_75t_L g636 ( 
.A(n_507),
.Y(n_636)
);

INVx1_ASAP7_75t_L g637 ( 
.A(n_528),
.Y(n_637)
);

INVx3_ASAP7_75t_L g638 ( 
.A(n_532),
.Y(n_638)
);

INVx1_ASAP7_75t_L g639 ( 
.A(n_529),
.Y(n_639)
);

INVx2_ASAP7_75t_L g640 ( 
.A(n_510),
.Y(n_640)
);

INVx1_ASAP7_75t_L g641 ( 
.A(n_529),
.Y(n_641)
);

INVx2_ASAP7_75t_L g642 ( 
.A(n_510),
.Y(n_642)
);

INVx1_ASAP7_75t_L g643 ( 
.A(n_535),
.Y(n_643)
);

INVx2_ASAP7_75t_L g644 ( 
.A(n_510),
.Y(n_644)
);

INVx1_ASAP7_75t_L g645 ( 
.A(n_535),
.Y(n_645)
);

INVx2_ASAP7_75t_L g646 ( 
.A(n_520),
.Y(n_646)
);

INVx2_ASAP7_75t_L g647 ( 
.A(n_520),
.Y(n_647)
);

BUFx6f_ASAP7_75t_L g648 ( 
.A(n_505),
.Y(n_648)
);

INVx1_ASAP7_75t_L g649 ( 
.A(n_535),
.Y(n_649)
);

INVx1_ASAP7_75t_L g650 ( 
.A(n_535),
.Y(n_650)
);

INVx1_ASAP7_75t_L g651 ( 
.A(n_561),
.Y(n_651)
);

AND2x2_ASAP7_75t_L g652 ( 
.A(n_519),
.B(n_414),
.Y(n_652)
);

BUFx3_ASAP7_75t_L g653 ( 
.A(n_527),
.Y(n_653)
);

INVx3_ASAP7_75t_L g654 ( 
.A(n_532),
.Y(n_654)
);

INVx3_ASAP7_75t_L g655 ( 
.A(n_518),
.Y(n_655)
);

INVx4_ASAP7_75t_L g656 ( 
.A(n_514),
.Y(n_656)
);

INVx2_ASAP7_75t_L g657 ( 
.A(n_520),
.Y(n_657)
);

INVx1_ASAP7_75t_L g658 ( 
.A(n_561),
.Y(n_658)
);

AND2x2_ASAP7_75t_L g659 ( 
.A(n_519),
.B(n_486),
.Y(n_659)
);

NAND2xp5_ASAP7_75t_SL g660 ( 
.A(n_516),
.B(n_418),
.Y(n_660)
);

NAND2xp33_ASAP7_75t_SL g661 ( 
.A(n_582),
.B(n_421),
.Y(n_661)
);

INVx2_ASAP7_75t_L g662 ( 
.A(n_531),
.Y(n_662)
);

INVx2_ASAP7_75t_L g663 ( 
.A(n_531),
.Y(n_663)
);

NAND2xp5_ASAP7_75t_L g664 ( 
.A(n_561),
.B(n_498),
.Y(n_664)
);

INVx1_ASAP7_75t_L g665 ( 
.A(n_565),
.Y(n_665)
);

NAND2xp5_ASAP7_75t_L g666 ( 
.A(n_565),
.B(n_329),
.Y(n_666)
);

NAND2xp5_ASAP7_75t_L g667 ( 
.A(n_565),
.B(n_329),
.Y(n_667)
);

INVx2_ASAP7_75t_L g668 ( 
.A(n_531),
.Y(n_668)
);

NAND2xp5_ASAP7_75t_SL g669 ( 
.A(n_516),
.B(n_421),
.Y(n_669)
);

INVx1_ASAP7_75t_L g670 ( 
.A(n_565),
.Y(n_670)
);

INVx1_ASAP7_75t_L g671 ( 
.A(n_558),
.Y(n_671)
);

INVx2_ASAP7_75t_L g672 ( 
.A(n_537),
.Y(n_672)
);

INVx2_ASAP7_75t_L g673 ( 
.A(n_537),
.Y(n_673)
);

OAI22xp5_ASAP7_75t_L g674 ( 
.A1(n_545),
.A2(n_209),
.B1(n_213),
.B2(n_205),
.Y(n_674)
);

BUFx6f_ASAP7_75t_L g675 ( 
.A(n_505),
.Y(n_675)
);

INVx1_ASAP7_75t_L g676 ( 
.A(n_558),
.Y(n_676)
);

INVx2_ASAP7_75t_L g677 ( 
.A(n_537),
.Y(n_677)
);

AND2x2_ASAP7_75t_L g678 ( 
.A(n_525),
.B(n_496),
.Y(n_678)
);

INVx1_ASAP7_75t_L g679 ( 
.A(n_558),
.Y(n_679)
);

INVx1_ASAP7_75t_L g680 ( 
.A(n_558),
.Y(n_680)
);

NAND2xp5_ASAP7_75t_SL g681 ( 
.A(n_547),
.B(n_429),
.Y(n_681)
);

BUFx10_ASAP7_75t_L g682 ( 
.A(n_578),
.Y(n_682)
);

NAND2xp5_ASAP7_75t_SL g683 ( 
.A(n_572),
.B(n_429),
.Y(n_683)
);

INVx2_ASAP7_75t_L g684 ( 
.A(n_542),
.Y(n_684)
);

INVx1_ASAP7_75t_L g685 ( 
.A(n_558),
.Y(n_685)
);

INVx2_ASAP7_75t_L g686 ( 
.A(n_542),
.Y(n_686)
);

AND2x2_ASAP7_75t_L g687 ( 
.A(n_525),
.B(n_496),
.Y(n_687)
);

INVx1_ASAP7_75t_L g688 ( 
.A(n_541),
.Y(n_688)
);

NAND2xp33_ASAP7_75t_SL g689 ( 
.A(n_572),
.B(n_437),
.Y(n_689)
);

NOR2xp33_ASAP7_75t_L g690 ( 
.A(n_550),
.B(n_437),
.Y(n_690)
);

INVx1_ASAP7_75t_L g691 ( 
.A(n_541),
.Y(n_691)
);

CKINVDCx5p33_ASAP7_75t_R g692 ( 
.A(n_508),
.Y(n_692)
);

INVx3_ASAP7_75t_L g693 ( 
.A(n_518),
.Y(n_693)
);

INVx1_ASAP7_75t_L g694 ( 
.A(n_551),
.Y(n_694)
);

AND2x2_ASAP7_75t_L g695 ( 
.A(n_525),
.B(n_404),
.Y(n_695)
);

OR2x6_ASAP7_75t_L g696 ( 
.A(n_536),
.B(n_285),
.Y(n_696)
);

AND3x2_ASAP7_75t_L g697 ( 
.A(n_513),
.B(n_224),
.C(n_219),
.Y(n_697)
);

INVx2_ASAP7_75t_L g698 ( 
.A(n_542),
.Y(n_698)
);

INVx1_ASAP7_75t_L g699 ( 
.A(n_551),
.Y(n_699)
);

INVx1_ASAP7_75t_L g700 ( 
.A(n_552),
.Y(n_700)
);

INVx1_ASAP7_75t_L g701 ( 
.A(n_552),
.Y(n_701)
);

INVx2_ASAP7_75t_SL g702 ( 
.A(n_512),
.Y(n_702)
);

INVx2_ASAP7_75t_L g703 ( 
.A(n_544),
.Y(n_703)
);

BUFx2_ASAP7_75t_L g704 ( 
.A(n_512),
.Y(n_704)
);

BUFx3_ASAP7_75t_L g705 ( 
.A(n_518),
.Y(n_705)
);

INVx4_ASAP7_75t_L g706 ( 
.A(n_514),
.Y(n_706)
);

NAND3xp33_ASAP7_75t_L g707 ( 
.A(n_499),
.B(n_432),
.C(n_431),
.Y(n_707)
);

AND2x2_ASAP7_75t_L g708 ( 
.A(n_539),
.B(n_434),
.Y(n_708)
);

NAND3xp33_ASAP7_75t_L g709 ( 
.A(n_499),
.B(n_444),
.C(n_438),
.Y(n_709)
);

INVx2_ASAP7_75t_L g710 ( 
.A(n_544),
.Y(n_710)
);

OR2x2_ASAP7_75t_L g711 ( 
.A(n_515),
.B(n_469),
.Y(n_711)
);

CKINVDCx16_ASAP7_75t_R g712 ( 
.A(n_578),
.Y(n_712)
);

INVx1_ASAP7_75t_L g713 ( 
.A(n_553),
.Y(n_713)
);

INVx2_ASAP7_75t_SL g714 ( 
.A(n_515),
.Y(n_714)
);

CKINVDCx6p67_ASAP7_75t_R g715 ( 
.A(n_506),
.Y(n_715)
);

INVx4_ASAP7_75t_L g716 ( 
.A(n_514),
.Y(n_716)
);

INVx2_ASAP7_75t_L g717 ( 
.A(n_544),
.Y(n_717)
);

AND2x2_ASAP7_75t_L g718 ( 
.A(n_539),
.B(n_445),
.Y(n_718)
);

NOR2xp33_ASAP7_75t_L g719 ( 
.A(n_550),
.B(n_440),
.Y(n_719)
);

INVx2_ASAP7_75t_L g720 ( 
.A(n_546),
.Y(n_720)
);

INVx2_ASAP7_75t_L g721 ( 
.A(n_546),
.Y(n_721)
);

NAND2xp5_ASAP7_75t_L g722 ( 
.A(n_509),
.B(n_329),
.Y(n_722)
);

NAND2xp5_ASAP7_75t_L g723 ( 
.A(n_509),
.B(n_346),
.Y(n_723)
);

INVx2_ASAP7_75t_L g724 ( 
.A(n_546),
.Y(n_724)
);

INVx2_ASAP7_75t_L g725 ( 
.A(n_556),
.Y(n_725)
);

INVx2_ASAP7_75t_L g726 ( 
.A(n_556),
.Y(n_726)
);

INVx2_ASAP7_75t_L g727 ( 
.A(n_556),
.Y(n_727)
);

INVx1_ASAP7_75t_L g728 ( 
.A(n_553),
.Y(n_728)
);

BUFx6f_ASAP7_75t_L g729 ( 
.A(n_505),
.Y(n_729)
);

INVx1_ASAP7_75t_L g730 ( 
.A(n_555),
.Y(n_730)
);

INVx1_ASAP7_75t_L g731 ( 
.A(n_555),
.Y(n_731)
);

INVx2_ASAP7_75t_L g732 ( 
.A(n_518),
.Y(n_732)
);

AND2x2_ASAP7_75t_SL g733 ( 
.A(n_509),
.B(n_265),
.Y(n_733)
);

INVxp67_ASAP7_75t_SL g734 ( 
.A(n_548),
.Y(n_734)
);

AOI22xp5_ASAP7_75t_L g735 ( 
.A1(n_591),
.A2(n_633),
.B1(n_610),
.B2(n_621),
.Y(n_735)
);

NAND2xp5_ASAP7_75t_SL g736 ( 
.A(n_610),
.B(n_501),
.Y(n_736)
);

NAND2xp5_ASAP7_75t_L g737 ( 
.A(n_733),
.B(n_509),
.Y(n_737)
);

INVx1_ASAP7_75t_L g738 ( 
.A(n_688),
.Y(n_738)
);

NOR2xp67_ASAP7_75t_L g739 ( 
.A(n_595),
.B(n_521),
.Y(n_739)
);

INVx1_ASAP7_75t_L g740 ( 
.A(n_688),
.Y(n_740)
);

NAND2xp5_ASAP7_75t_L g741 ( 
.A(n_733),
.B(n_691),
.Y(n_741)
);

AOI21xp5_ASAP7_75t_L g742 ( 
.A1(n_609),
.A2(n_536),
.B(n_505),
.Y(n_742)
);

INVx1_ASAP7_75t_L g743 ( 
.A(n_691),
.Y(n_743)
);

INVx3_ASAP7_75t_L g744 ( 
.A(n_705),
.Y(n_744)
);

AND2x2_ASAP7_75t_L g745 ( 
.A(n_702),
.B(n_440),
.Y(n_745)
);

NOR2xp33_ASAP7_75t_L g746 ( 
.A(n_690),
.B(n_517),
.Y(n_746)
);

NAND2xp5_ASAP7_75t_SL g747 ( 
.A(n_733),
.B(n_317),
.Y(n_747)
);

NOR2xp33_ASAP7_75t_L g748 ( 
.A(n_719),
.B(n_579),
.Y(n_748)
);

OAI221xp5_ASAP7_75t_L g749 ( 
.A1(n_601),
.A2(n_503),
.B1(n_577),
.B2(n_549),
.C(n_563),
.Y(n_749)
);

NAND2xp5_ASAP7_75t_L g750 ( 
.A(n_694),
.B(n_526),
.Y(n_750)
);

NAND2xp5_ASAP7_75t_L g751 ( 
.A(n_694),
.B(n_526),
.Y(n_751)
);

NOR2xp33_ASAP7_75t_L g752 ( 
.A(n_660),
.B(n_441),
.Y(n_752)
);

NAND2xp5_ASAP7_75t_L g753 ( 
.A(n_699),
.B(n_526),
.Y(n_753)
);

NAND2xp5_ASAP7_75t_SL g754 ( 
.A(n_616),
.B(n_317),
.Y(n_754)
);

INVx2_ASAP7_75t_SL g755 ( 
.A(n_695),
.Y(n_755)
);

AND2x2_ASAP7_75t_L g756 ( 
.A(n_702),
.B(n_441),
.Y(n_756)
);

NAND2xp5_ASAP7_75t_L g757 ( 
.A(n_699),
.B(n_526),
.Y(n_757)
);

INVx2_ASAP7_75t_L g758 ( 
.A(n_583),
.Y(n_758)
);

NOR3xp33_ASAP7_75t_L g759 ( 
.A(n_622),
.B(n_554),
.C(n_712),
.Y(n_759)
);

NOR2xp33_ASAP7_75t_SL g760 ( 
.A(n_607),
.B(n_523),
.Y(n_760)
);

NAND2xp5_ASAP7_75t_SL g761 ( 
.A(n_616),
.B(n_317),
.Y(n_761)
);

INVx2_ASAP7_75t_L g762 ( 
.A(n_583),
.Y(n_762)
);

NAND2xp5_ASAP7_75t_SL g763 ( 
.A(n_616),
.B(n_317),
.Y(n_763)
);

NOR2xp33_ASAP7_75t_L g764 ( 
.A(n_669),
.B(n_456),
.Y(n_764)
);

NAND2xp5_ASAP7_75t_L g765 ( 
.A(n_700),
.B(n_539),
.Y(n_765)
);

NAND2xp5_ASAP7_75t_L g766 ( 
.A(n_700),
.B(n_577),
.Y(n_766)
);

INVxp33_ASAP7_75t_L g767 ( 
.A(n_704),
.Y(n_767)
);

NAND3xp33_ASAP7_75t_L g768 ( 
.A(n_617),
.B(n_478),
.C(n_456),
.Y(n_768)
);

INVxp67_ASAP7_75t_SL g769 ( 
.A(n_614),
.Y(n_769)
);

NAND2xp5_ASAP7_75t_SL g770 ( 
.A(n_616),
.B(n_317),
.Y(n_770)
);

INVx3_ASAP7_75t_L g771 ( 
.A(n_705),
.Y(n_771)
);

INVx1_ASAP7_75t_L g772 ( 
.A(n_701),
.Y(n_772)
);

INVx1_ASAP7_75t_L g773 ( 
.A(n_713),
.Y(n_773)
);

INVx1_ASAP7_75t_L g774 ( 
.A(n_713),
.Y(n_774)
);

AND2x4_ASAP7_75t_L g775 ( 
.A(n_589),
.B(n_559),
.Y(n_775)
);

BUFx3_ASAP7_75t_L g776 ( 
.A(n_589),
.Y(n_776)
);

NAND2xp5_ASAP7_75t_L g777 ( 
.A(n_728),
.B(n_478),
.Y(n_777)
);

NAND2xp5_ASAP7_75t_L g778 ( 
.A(n_728),
.B(n_482),
.Y(n_778)
);

NAND2xp5_ASAP7_75t_L g779 ( 
.A(n_730),
.B(n_482),
.Y(n_779)
);

NAND2xp5_ASAP7_75t_SL g780 ( 
.A(n_585),
.B(n_714),
.Y(n_780)
);

INVx2_ASAP7_75t_L g781 ( 
.A(n_583),
.Y(n_781)
);

INVx3_ASAP7_75t_L g782 ( 
.A(n_705),
.Y(n_782)
);

NAND2xp5_ASAP7_75t_L g783 ( 
.A(n_730),
.B(n_487),
.Y(n_783)
);

BUFx6f_ASAP7_75t_L g784 ( 
.A(n_589),
.Y(n_784)
);

OAI22xp33_ASAP7_75t_L g785 ( 
.A1(n_592),
.A2(n_503),
.B1(n_554),
.B2(n_426),
.Y(n_785)
);

NAND2xp5_ASAP7_75t_SL g786 ( 
.A(n_585),
.B(n_501),
.Y(n_786)
);

NAND2xp5_ASAP7_75t_L g787 ( 
.A(n_731),
.B(n_487),
.Y(n_787)
);

OR2x6_ASAP7_75t_L g788 ( 
.A(n_714),
.B(n_704),
.Y(n_788)
);

AOI22xp5_ASAP7_75t_L g789 ( 
.A1(n_643),
.A2(n_410),
.B1(n_424),
.B2(n_398),
.Y(n_789)
);

AND2x2_ASAP7_75t_SL g790 ( 
.A(n_712),
.B(n_318),
.Y(n_790)
);

AOI22xp5_ASAP7_75t_L g791 ( 
.A1(n_643),
.A2(n_433),
.B1(n_457),
.B2(n_430),
.Y(n_791)
);

NAND2xp5_ASAP7_75t_L g792 ( 
.A(n_671),
.B(n_676),
.Y(n_792)
);

INVx2_ASAP7_75t_L g793 ( 
.A(n_584),
.Y(n_793)
);

AOI22xp5_ASAP7_75t_L g794 ( 
.A1(n_645),
.A2(n_465),
.B1(n_488),
.B2(n_338),
.Y(n_794)
);

NAND2xp5_ASAP7_75t_L g795 ( 
.A(n_671),
.B(n_488),
.Y(n_795)
);

NAND2xp5_ASAP7_75t_SL g796 ( 
.A(n_695),
.B(n_501),
.Y(n_796)
);

NAND2xp5_ASAP7_75t_SL g797 ( 
.A(n_656),
.B(n_318),
.Y(n_797)
);

INVx8_ASAP7_75t_L g798 ( 
.A(n_696),
.Y(n_798)
);

INVx2_ASAP7_75t_L g799 ( 
.A(n_584),
.Y(n_799)
);

NAND2xp5_ASAP7_75t_L g800 ( 
.A(n_676),
.B(n_679),
.Y(n_800)
);

INVx1_ASAP7_75t_L g801 ( 
.A(n_645),
.Y(n_801)
);

NAND2xp5_ASAP7_75t_SL g802 ( 
.A(n_656),
.B(n_706),
.Y(n_802)
);

INVx2_ASAP7_75t_L g803 ( 
.A(n_584),
.Y(n_803)
);

NAND2xp5_ASAP7_75t_L g804 ( 
.A(n_679),
.B(n_680),
.Y(n_804)
);

INVx2_ASAP7_75t_L g805 ( 
.A(n_586),
.Y(n_805)
);

NAND2xp5_ASAP7_75t_L g806 ( 
.A(n_680),
.B(n_548),
.Y(n_806)
);

NAND2xp5_ASAP7_75t_L g807 ( 
.A(n_685),
.B(n_548),
.Y(n_807)
);

NAND3xp33_ASAP7_75t_L g808 ( 
.A(n_592),
.B(n_511),
.C(n_501),
.Y(n_808)
);

INVx2_ASAP7_75t_L g809 ( 
.A(n_586),
.Y(n_809)
);

NOR2xp33_ASAP7_75t_SL g810 ( 
.A(n_629),
.B(n_533),
.Y(n_810)
);

INVx1_ASAP7_75t_L g811 ( 
.A(n_649),
.Y(n_811)
);

INVx2_ASAP7_75t_SL g812 ( 
.A(n_606),
.Y(n_812)
);

NOR2xp33_ASAP7_75t_L g813 ( 
.A(n_681),
.B(n_549),
.Y(n_813)
);

INVx1_ASAP7_75t_L g814 ( 
.A(n_649),
.Y(n_814)
);

NAND2xp33_ASAP7_75t_SL g815 ( 
.A(n_711),
.B(n_205),
.Y(n_815)
);

INVx2_ASAP7_75t_L g816 ( 
.A(n_586),
.Y(n_816)
);

BUFx3_ASAP7_75t_L g817 ( 
.A(n_623),
.Y(n_817)
);

BUFx6f_ASAP7_75t_SL g818 ( 
.A(n_629),
.Y(n_818)
);

INVx2_ASAP7_75t_L g819 ( 
.A(n_588),
.Y(n_819)
);

INVxp33_ASAP7_75t_L g820 ( 
.A(n_711),
.Y(n_820)
);

INVx2_ASAP7_75t_L g821 ( 
.A(n_588),
.Y(n_821)
);

NAND2xp5_ASAP7_75t_SL g822 ( 
.A(n_656),
.B(n_318),
.Y(n_822)
);

NOR2xp33_ASAP7_75t_L g823 ( 
.A(n_683),
.B(n_197),
.Y(n_823)
);

NOR3xp33_ASAP7_75t_L g824 ( 
.A(n_622),
.B(n_534),
.C(n_365),
.Y(n_824)
);

OR2x2_ASAP7_75t_L g825 ( 
.A(n_689),
.B(n_559),
.Y(n_825)
);

INVx2_ASAP7_75t_L g826 ( 
.A(n_588),
.Y(n_826)
);

NAND2xp5_ASAP7_75t_SL g827 ( 
.A(n_656),
.B(n_318),
.Y(n_827)
);

OAI22xp5_ASAP7_75t_L g828 ( 
.A1(n_651),
.A2(n_665),
.B1(n_670),
.B2(n_658),
.Y(n_828)
);

INVx1_ASAP7_75t_L g829 ( 
.A(n_650),
.Y(n_829)
);

INVx2_ASAP7_75t_L g830 ( 
.A(n_590),
.Y(n_830)
);

AOI22xp5_ASAP7_75t_L g831 ( 
.A1(n_650),
.A2(n_221),
.B1(n_337),
.B2(n_284),
.Y(n_831)
);

NAND2xp5_ASAP7_75t_L g832 ( 
.A(n_685),
.B(n_548),
.Y(n_832)
);

INVx8_ASAP7_75t_L g833 ( 
.A(n_696),
.Y(n_833)
);

NAND2xp5_ASAP7_75t_SL g834 ( 
.A(n_706),
.B(n_318),
.Y(n_834)
);

NAND2xp5_ASAP7_75t_L g835 ( 
.A(n_665),
.B(n_540),
.Y(n_835)
);

NOR2xp33_ASAP7_75t_L g836 ( 
.A(n_623),
.B(n_204),
.Y(n_836)
);

AOI22xp33_ASAP7_75t_L g837 ( 
.A1(n_606),
.A2(n_346),
.B1(n_226),
.B2(n_254),
.Y(n_837)
);

INVx1_ASAP7_75t_L g838 ( 
.A(n_670),
.Y(n_838)
);

NOR3xp33_ASAP7_75t_L g839 ( 
.A(n_627),
.B(n_447),
.C(n_446),
.Y(n_839)
);

INVx1_ASAP7_75t_L g840 ( 
.A(n_639),
.Y(n_840)
);

INVx1_ASAP7_75t_L g841 ( 
.A(n_639),
.Y(n_841)
);

NOR2xp33_ASAP7_75t_L g842 ( 
.A(n_623),
.B(n_204),
.Y(n_842)
);

NAND2xp5_ASAP7_75t_SL g843 ( 
.A(n_706),
.B(n_346),
.Y(n_843)
);

NOR2xp33_ASAP7_75t_L g844 ( 
.A(n_653),
.B(n_208),
.Y(n_844)
);

NOR2xp33_ASAP7_75t_L g845 ( 
.A(n_653),
.B(n_208),
.Y(n_845)
);

NOR2xp33_ASAP7_75t_SL g846 ( 
.A(n_629),
.B(n_511),
.Y(n_846)
);

NOR2xp33_ASAP7_75t_L g847 ( 
.A(n_653),
.B(n_210),
.Y(n_847)
);

NAND2xp5_ASAP7_75t_L g848 ( 
.A(n_600),
.B(n_540),
.Y(n_848)
);

NOR2xp33_ASAP7_75t_L g849 ( 
.A(n_696),
.B(n_210),
.Y(n_849)
);

NOR2xp33_ASAP7_75t_L g850 ( 
.A(n_696),
.B(n_214),
.Y(n_850)
);

NOR2xp33_ASAP7_75t_SL g851 ( 
.A(n_629),
.B(n_511),
.Y(n_851)
);

NAND2xp5_ASAP7_75t_SL g852 ( 
.A(n_706),
.B(n_346),
.Y(n_852)
);

INVx4_ASAP7_75t_L g853 ( 
.A(n_618),
.Y(n_853)
);

INVx2_ASAP7_75t_L g854 ( 
.A(n_590),
.Y(n_854)
);

INVx1_ASAP7_75t_L g855 ( 
.A(n_641),
.Y(n_855)
);

BUFx3_ASAP7_75t_L g856 ( 
.A(n_708),
.Y(n_856)
);

NAND2xp5_ASAP7_75t_SL g857 ( 
.A(n_716),
.B(n_346),
.Y(n_857)
);

AOI22xp33_ASAP7_75t_SL g858 ( 
.A1(n_674),
.A2(n_511),
.B1(n_362),
.B2(n_360),
.Y(n_858)
);

NAND2x1_ASAP7_75t_L g859 ( 
.A(n_716),
.B(n_614),
.Y(n_859)
);

INVx1_ASAP7_75t_L g860 ( 
.A(n_641),
.Y(n_860)
);

AND2x2_ASAP7_75t_SL g861 ( 
.A(n_722),
.B(n_259),
.Y(n_861)
);

NOR2xp33_ASAP7_75t_L g862 ( 
.A(n_696),
.B(n_214),
.Y(n_862)
);

OR2x6_ASAP7_75t_L g863 ( 
.A(n_659),
.B(n_448),
.Y(n_863)
);

AOI22xp5_ASAP7_75t_L g864 ( 
.A1(n_661),
.A2(n_336),
.B1(n_266),
.B2(n_263),
.Y(n_864)
);

INVx2_ASAP7_75t_L g865 ( 
.A(n_590),
.Y(n_865)
);

INVx3_ASAP7_75t_L g866 ( 
.A(n_655),
.Y(n_866)
);

NAND2xp5_ASAP7_75t_L g867 ( 
.A(n_600),
.B(n_608),
.Y(n_867)
);

AOI22xp33_ASAP7_75t_L g868 ( 
.A1(n_652),
.A2(n_346),
.B1(n_264),
.B2(n_277),
.Y(n_868)
);

NAND2xp33_ASAP7_75t_L g869 ( 
.A(n_608),
.B(n_615),
.Y(n_869)
);

NAND2xp5_ASAP7_75t_L g870 ( 
.A(n_615),
.B(n_261),
.Y(n_870)
);

NOR2xp33_ASAP7_75t_L g871 ( 
.A(n_620),
.B(n_218),
.Y(n_871)
);

AOI22xp33_ASAP7_75t_L g872 ( 
.A1(n_652),
.A2(n_346),
.B1(n_278),
.B2(n_335),
.Y(n_872)
);

OAI22xp5_ASAP7_75t_SL g873 ( 
.A1(n_602),
.A2(n_213),
.B1(n_209),
.B2(n_360),
.Y(n_873)
);

NAND2xp5_ASAP7_75t_L g874 ( 
.A(n_620),
.B(n_282),
.Y(n_874)
);

AND2x2_ASAP7_75t_L g875 ( 
.A(n_659),
.B(n_569),
.Y(n_875)
);

NAND2xp5_ASAP7_75t_SL g876 ( 
.A(n_716),
.B(n_283),
.Y(n_876)
);

INVx2_ASAP7_75t_L g877 ( 
.A(n_593),
.Y(n_877)
);

NAND2xp5_ASAP7_75t_L g878 ( 
.A(n_624),
.B(n_290),
.Y(n_878)
);

INVx8_ASAP7_75t_L g879 ( 
.A(n_692),
.Y(n_879)
);

AOI22xp5_ASAP7_75t_L g880 ( 
.A1(n_715),
.A2(n_300),
.B1(n_280),
.B2(n_281),
.Y(n_880)
);

NAND2xp5_ASAP7_75t_L g881 ( 
.A(n_624),
.B(n_626),
.Y(n_881)
);

AND2x2_ASAP7_75t_SL g882 ( 
.A(n_722),
.B(n_293),
.Y(n_882)
);

NAND2xp5_ASAP7_75t_L g883 ( 
.A(n_626),
.B(n_312),
.Y(n_883)
);

NAND2xp5_ASAP7_75t_L g884 ( 
.A(n_631),
.B(n_326),
.Y(n_884)
);

O2A1O1Ixp33_ASAP7_75t_L g885 ( 
.A1(n_678),
.A2(n_450),
.B(n_449),
.C(n_452),
.Y(n_885)
);

NOR3xp33_ASAP7_75t_L g886 ( 
.A(n_674),
.B(n_455),
.C(n_453),
.Y(n_886)
);

AOI22xp5_ASAP7_75t_L g887 ( 
.A1(n_715),
.A2(n_718),
.B1(n_708),
.B2(n_687),
.Y(n_887)
);

HB1xp67_ASAP7_75t_L g888 ( 
.A(n_678),
.Y(n_888)
);

NAND2xp5_ASAP7_75t_L g889 ( 
.A(n_637),
.B(n_350),
.Y(n_889)
);

NAND2xp5_ASAP7_75t_L g890 ( 
.A(n_734),
.B(n_352),
.Y(n_890)
);

NAND2xp5_ASAP7_75t_SL g891 ( 
.A(n_609),
.B(n_358),
.Y(n_891)
);

CKINVDCx5p33_ASAP7_75t_R g892 ( 
.A(n_715),
.Y(n_892)
);

INVx1_ASAP7_75t_L g893 ( 
.A(n_718),
.Y(n_893)
);

OR2x2_ASAP7_75t_L g894 ( 
.A(n_687),
.B(n_461),
.Y(n_894)
);

NAND2xp5_ASAP7_75t_L g895 ( 
.A(n_664),
.B(n_366),
.Y(n_895)
);

NAND3xp33_ASAP7_75t_SL g896 ( 
.A(n_707),
.B(n_362),
.C(n_364),
.Y(n_896)
);

INVx2_ASAP7_75t_L g897 ( 
.A(n_593),
.Y(n_897)
);

INVx2_ASAP7_75t_L g898 ( 
.A(n_838),
.Y(n_898)
);

INVx3_ASAP7_75t_L g899 ( 
.A(n_784),
.Y(n_899)
);

AND2x6_ASAP7_75t_L g900 ( 
.A(n_792),
.B(n_723),
.Y(n_900)
);

NOR2xp33_ASAP7_75t_L g901 ( 
.A(n_735),
.B(n_682),
.Y(n_901)
);

AOI21xp5_ASAP7_75t_L g902 ( 
.A1(n_802),
.A2(n_635),
.B(n_614),
.Y(n_902)
);

INVx1_ASAP7_75t_L g903 ( 
.A(n_801),
.Y(n_903)
);

BUFx3_ASAP7_75t_L g904 ( 
.A(n_879),
.Y(n_904)
);

AND2x4_ASAP7_75t_L g905 ( 
.A(n_856),
.B(n_697),
.Y(n_905)
);

INVx2_ASAP7_75t_L g906 ( 
.A(n_811),
.Y(n_906)
);

A2O1A1Ixp33_ASAP7_75t_L g907 ( 
.A1(n_746),
.A2(n_723),
.B(n_709),
.C(n_707),
.Y(n_907)
);

NOR2xp33_ASAP7_75t_L g908 ( 
.A(n_746),
.B(n_682),
.Y(n_908)
);

AOI21xp5_ASAP7_75t_L g909 ( 
.A1(n_802),
.A2(n_635),
.B(n_614),
.Y(n_909)
);

AND2x4_ASAP7_75t_L g910 ( 
.A(n_856),
.B(n_709),
.Y(n_910)
);

INVx1_ASAP7_75t_L g911 ( 
.A(n_814),
.Y(n_911)
);

INVx2_ASAP7_75t_SL g912 ( 
.A(n_788),
.Y(n_912)
);

BUFx4f_ASAP7_75t_L g913 ( 
.A(n_879),
.Y(n_913)
);

INVx2_ASAP7_75t_L g914 ( 
.A(n_866),
.Y(n_914)
);

NAND2xp5_ASAP7_75t_L g915 ( 
.A(n_766),
.B(n_664),
.Y(n_915)
);

INVx3_ASAP7_75t_L g916 ( 
.A(n_784),
.Y(n_916)
);

NOR2xp33_ASAP7_75t_SL g917 ( 
.A(n_760),
.B(n_682),
.Y(n_917)
);

INVx1_ASAP7_75t_L g918 ( 
.A(n_829),
.Y(n_918)
);

INVx2_ASAP7_75t_L g919 ( 
.A(n_866),
.Y(n_919)
);

NAND2xp5_ASAP7_75t_L g920 ( 
.A(n_769),
.B(n_635),
.Y(n_920)
);

INVx1_ASAP7_75t_L g921 ( 
.A(n_738),
.Y(n_921)
);

NAND2xp5_ASAP7_75t_SL g922 ( 
.A(n_861),
.B(n_682),
.Y(n_922)
);

NAND2xp5_ASAP7_75t_L g923 ( 
.A(n_795),
.B(n_635),
.Y(n_923)
);

NAND2xp5_ASAP7_75t_L g924 ( 
.A(n_840),
.B(n_638),
.Y(n_924)
);

NAND2xp5_ASAP7_75t_L g925 ( 
.A(n_841),
.B(n_638),
.Y(n_925)
);

BUFx6f_ASAP7_75t_L g926 ( 
.A(n_784),
.Y(n_926)
);

OR2x6_ASAP7_75t_L g927 ( 
.A(n_879),
.B(n_666),
.Y(n_927)
);

BUFx2_ASAP7_75t_L g928 ( 
.A(n_788),
.Y(n_928)
);

NAND2xp5_ASAP7_75t_L g929 ( 
.A(n_855),
.B(n_638),
.Y(n_929)
);

INVx1_ASAP7_75t_L g930 ( 
.A(n_740),
.Y(n_930)
);

INVxp67_ASAP7_75t_L g931 ( 
.A(n_745),
.Y(n_931)
);

HB1xp67_ASAP7_75t_L g932 ( 
.A(n_788),
.Y(n_932)
);

BUFx3_ASAP7_75t_L g933 ( 
.A(n_776),
.Y(n_933)
);

NOR2xp33_ASAP7_75t_L g934 ( 
.A(n_748),
.B(n_625),
.Y(n_934)
);

BUFx4f_ASAP7_75t_L g935 ( 
.A(n_798),
.Y(n_935)
);

NAND2x1p5_ASAP7_75t_L g936 ( 
.A(n_776),
.B(n_618),
.Y(n_936)
);

INVx2_ASAP7_75t_L g937 ( 
.A(n_758),
.Y(n_937)
);

INVx1_ASAP7_75t_L g938 ( 
.A(n_743),
.Y(n_938)
);

HB1xp67_ASAP7_75t_L g939 ( 
.A(n_888),
.Y(n_939)
);

NAND2xp5_ASAP7_75t_SL g940 ( 
.A(n_861),
.B(n_638),
.Y(n_940)
);

INVx2_ASAP7_75t_SL g941 ( 
.A(n_894),
.Y(n_941)
);

NAND2xp5_ASAP7_75t_SL g942 ( 
.A(n_882),
.B(n_654),
.Y(n_942)
);

BUFx3_ASAP7_75t_L g943 ( 
.A(n_817),
.Y(n_943)
);

INVx1_ASAP7_75t_L g944 ( 
.A(n_772),
.Y(n_944)
);

HB1xp67_ASAP7_75t_L g945 ( 
.A(n_888),
.Y(n_945)
);

NAND2xp5_ASAP7_75t_L g946 ( 
.A(n_860),
.B(n_654),
.Y(n_946)
);

AND2x6_ASAP7_75t_SL g947 ( 
.A(n_748),
.B(n_570),
.Y(n_947)
);

AOI22xp33_ASAP7_75t_L g948 ( 
.A1(n_882),
.A2(n_666),
.B1(n_667),
.B2(n_597),
.Y(n_948)
);

AOI21xp5_ASAP7_75t_L g949 ( 
.A1(n_859),
.A2(n_654),
.B(n_667),
.Y(n_949)
);

NAND2xp5_ASAP7_75t_SL g950 ( 
.A(n_790),
.B(n_654),
.Y(n_950)
);

BUFx2_ASAP7_75t_SL g951 ( 
.A(n_818),
.Y(n_951)
);

NAND2xp5_ASAP7_75t_SL g952 ( 
.A(n_790),
.B(n_618),
.Y(n_952)
);

INVx2_ASAP7_75t_L g953 ( 
.A(n_762),
.Y(n_953)
);

NAND2xp5_ASAP7_75t_SL g954 ( 
.A(n_741),
.B(n_618),
.Y(n_954)
);

INVx1_ASAP7_75t_L g955 ( 
.A(n_773),
.Y(n_955)
);

INVx2_ASAP7_75t_SL g956 ( 
.A(n_863),
.Y(n_956)
);

BUFx3_ASAP7_75t_L g957 ( 
.A(n_817),
.Y(n_957)
);

CKINVDCx20_ASAP7_75t_R g958 ( 
.A(n_789),
.Y(n_958)
);

NAND2xp5_ASAP7_75t_L g959 ( 
.A(n_774),
.B(n_655),
.Y(n_959)
);

AND2x4_ASAP7_75t_L g960 ( 
.A(n_755),
.B(n_570),
.Y(n_960)
);

NAND2xp5_ASAP7_75t_SL g961 ( 
.A(n_887),
.B(n_618),
.Y(n_961)
);

INVx2_ASAP7_75t_SL g962 ( 
.A(n_863),
.Y(n_962)
);

INVx2_ASAP7_75t_L g963 ( 
.A(n_781),
.Y(n_963)
);

OAI22xp5_ASAP7_75t_L g964 ( 
.A1(n_737),
.A2(n_693),
.B1(n_655),
.B2(n_604),
.Y(n_964)
);

OR2x2_ASAP7_75t_L g965 ( 
.A(n_780),
.B(n_767),
.Y(n_965)
);

INVx1_ASAP7_75t_L g966 ( 
.A(n_812),
.Y(n_966)
);

BUFx2_ASAP7_75t_L g967 ( 
.A(n_791),
.Y(n_967)
);

NAND2xp5_ASAP7_75t_L g968 ( 
.A(n_867),
.B(n_693),
.Y(n_968)
);

NAND2xp5_ASAP7_75t_L g969 ( 
.A(n_881),
.B(n_693),
.Y(n_969)
);

AOI22xp33_ASAP7_75t_L g970 ( 
.A1(n_837),
.A2(n_587),
.B1(n_594),
.B2(n_596),
.Y(n_970)
);

INVx6_ASAP7_75t_L g971 ( 
.A(n_775),
.Y(n_971)
);

NAND2xp5_ASAP7_75t_L g972 ( 
.A(n_875),
.B(n_693),
.Y(n_972)
);

BUFx8_ASAP7_75t_SL g973 ( 
.A(n_818),
.Y(n_973)
);

INVx1_ASAP7_75t_L g974 ( 
.A(n_893),
.Y(n_974)
);

BUFx12f_ASAP7_75t_L g975 ( 
.A(n_892),
.Y(n_975)
);

BUFx6f_ASAP7_75t_L g976 ( 
.A(n_744),
.Y(n_976)
);

BUFx3_ASAP7_75t_L g977 ( 
.A(n_775),
.Y(n_977)
);

NAND2xp5_ASAP7_75t_SL g978 ( 
.A(n_750),
.B(n_618),
.Y(n_978)
);

NAND2xp5_ASAP7_75t_L g979 ( 
.A(n_800),
.B(n_603),
.Y(n_979)
);

BUFx3_ASAP7_75t_L g980 ( 
.A(n_798),
.Y(n_980)
);

HB1xp67_ASAP7_75t_L g981 ( 
.A(n_863),
.Y(n_981)
);

BUFx6f_ASAP7_75t_L g982 ( 
.A(n_771),
.Y(n_982)
);

NAND2xp5_ASAP7_75t_L g983 ( 
.A(n_804),
.B(n_603),
.Y(n_983)
);

NAND2xp5_ASAP7_75t_L g984 ( 
.A(n_813),
.B(n_603),
.Y(n_984)
);

INVx3_ASAP7_75t_SL g985 ( 
.A(n_736),
.Y(n_985)
);

NAND2xp5_ASAP7_75t_SL g986 ( 
.A(n_751),
.B(n_753),
.Y(n_986)
);

NAND2xp5_ASAP7_75t_SL g987 ( 
.A(n_757),
.B(n_604),
.Y(n_987)
);

OR2x2_ASAP7_75t_SL g988 ( 
.A(n_808),
.B(n_573),
.Y(n_988)
);

A2O1A1Ixp33_ASAP7_75t_L g989 ( 
.A1(n_823),
.A2(n_384),
.B(n_364),
.C(n_368),
.Y(n_989)
);

AND2x4_ASAP7_75t_L g990 ( 
.A(n_839),
.B(n_573),
.Y(n_990)
);

INVx2_ASAP7_75t_SL g991 ( 
.A(n_756),
.Y(n_991)
);

NAND2xp5_ASAP7_75t_L g992 ( 
.A(n_813),
.B(n_604),
.Y(n_992)
);

NOR2xp33_ASAP7_75t_L g993 ( 
.A(n_777),
.B(n_605),
.Y(n_993)
);

INVx6_ASAP7_75t_L g994 ( 
.A(n_798),
.Y(n_994)
);

INVx2_ASAP7_75t_L g995 ( 
.A(n_793),
.Y(n_995)
);

INVx2_ASAP7_75t_SL g996 ( 
.A(n_825),
.Y(n_996)
);

A2O1A1Ixp33_ASAP7_75t_L g997 ( 
.A1(n_823),
.A2(n_368),
.B(n_373),
.C(n_376),
.Y(n_997)
);

INVx5_ASAP7_75t_L g998 ( 
.A(n_853),
.Y(n_998)
);

NOR2xp33_ASAP7_75t_L g999 ( 
.A(n_778),
.B(n_605),
.Y(n_999)
);

INVx1_ASAP7_75t_L g1000 ( 
.A(n_835),
.Y(n_1000)
);

INVx1_ASAP7_75t_L g1001 ( 
.A(n_848),
.Y(n_1001)
);

INVx1_ASAP7_75t_L g1002 ( 
.A(n_765),
.Y(n_1002)
);

AOI22xp33_ASAP7_75t_L g1003 ( 
.A1(n_837),
.A2(n_587),
.B1(n_594),
.B2(n_596),
.Y(n_1003)
);

OR2x2_ASAP7_75t_L g1004 ( 
.A(n_820),
.B(n_779),
.Y(n_1004)
);

AND2x2_ASAP7_75t_L g1005 ( 
.A(n_752),
.B(n_575),
.Y(n_1005)
);

AND2x4_ASAP7_75t_L g1006 ( 
.A(n_786),
.B(n_796),
.Y(n_1006)
);

NAND2xp5_ASAP7_75t_L g1007 ( 
.A(n_871),
.B(n_611),
.Y(n_1007)
);

INVx1_ASAP7_75t_L g1008 ( 
.A(n_828),
.Y(n_1008)
);

INVx1_ASAP7_75t_L g1009 ( 
.A(n_869),
.Y(n_1009)
);

NAND2xp5_ASAP7_75t_SL g1010 ( 
.A(n_783),
.B(n_787),
.Y(n_1010)
);

NAND2xp5_ASAP7_75t_L g1011 ( 
.A(n_871),
.B(n_611),
.Y(n_1011)
);

NAND2xp5_ASAP7_75t_L g1012 ( 
.A(n_836),
.B(n_611),
.Y(n_1012)
);

AOI22xp5_ASAP7_75t_L g1013 ( 
.A1(n_752),
.A2(n_605),
.B1(n_612),
.B2(n_613),
.Y(n_1013)
);

INVx1_ASAP7_75t_L g1014 ( 
.A(n_799),
.Y(n_1014)
);

NOR2xp33_ASAP7_75t_L g1015 ( 
.A(n_764),
.B(n_605),
.Y(n_1015)
);

NAND2xp5_ASAP7_75t_SL g1016 ( 
.A(n_853),
.B(n_612),
.Y(n_1016)
);

OAI21xp5_ASAP7_75t_L g1017 ( 
.A1(n_806),
.A2(n_832),
.B(n_807),
.Y(n_1017)
);

INVx2_ASAP7_75t_L g1018 ( 
.A(n_803),
.Y(n_1018)
);

INVx2_ASAP7_75t_L g1019 ( 
.A(n_805),
.Y(n_1019)
);

AND2x2_ASAP7_75t_L g1020 ( 
.A(n_764),
.B(n_794),
.Y(n_1020)
);

INVx1_ASAP7_75t_L g1021 ( 
.A(n_809),
.Y(n_1021)
);

INVx2_ASAP7_75t_SL g1022 ( 
.A(n_870),
.Y(n_1022)
);

NOR2xp33_ASAP7_75t_R g1023 ( 
.A(n_810),
.B(n_220),
.Y(n_1023)
);

O2A1O1Ixp33_ASAP7_75t_L g1024 ( 
.A1(n_749),
.A2(n_597),
.B(n_599),
.C(n_598),
.Y(n_1024)
);

BUFx6f_ASAP7_75t_L g1025 ( 
.A(n_771),
.Y(n_1025)
);

INVx1_ASAP7_75t_L g1026 ( 
.A(n_816),
.Y(n_1026)
);

BUFx4f_ASAP7_75t_L g1027 ( 
.A(n_833),
.Y(n_1027)
);

INVxp67_ASAP7_75t_L g1028 ( 
.A(n_815),
.Y(n_1028)
);

AOI22xp33_ASAP7_75t_L g1029 ( 
.A1(n_868),
.A2(n_872),
.B1(n_747),
.B2(n_873),
.Y(n_1029)
);

NAND2xp5_ASAP7_75t_SL g1030 ( 
.A(n_782),
.B(n_612),
.Y(n_1030)
);

BUFx4f_ASAP7_75t_L g1031 ( 
.A(n_833),
.Y(n_1031)
);

NOR2x1_ASAP7_75t_L g1032 ( 
.A(n_739),
.B(n_768),
.Y(n_1032)
);

AOI22xp33_ASAP7_75t_L g1033 ( 
.A1(n_868),
.A2(n_599),
.B1(n_593),
.B2(n_598),
.Y(n_1033)
);

CKINVDCx20_ASAP7_75t_R g1034 ( 
.A(n_880),
.Y(n_1034)
);

CKINVDCx5p33_ASAP7_75t_R g1035 ( 
.A(n_864),
.Y(n_1035)
);

INVx2_ASAP7_75t_L g1036 ( 
.A(n_819),
.Y(n_1036)
);

INVx2_ASAP7_75t_L g1037 ( 
.A(n_821),
.Y(n_1037)
);

NAND2xp5_ASAP7_75t_SL g1038 ( 
.A(n_782),
.B(n_612),
.Y(n_1038)
);

AOI22xp33_ASAP7_75t_L g1039 ( 
.A1(n_872),
.A2(n_747),
.B1(n_896),
.B2(n_785),
.Y(n_1039)
);

NAND2xp5_ASAP7_75t_SL g1040 ( 
.A(n_895),
.B(n_613),
.Y(n_1040)
);

NOR2xp33_ASAP7_75t_L g1041 ( 
.A(n_785),
.B(n_613),
.Y(n_1041)
);

HB1xp67_ASAP7_75t_L g1042 ( 
.A(n_890),
.Y(n_1042)
);

INVx4_ASAP7_75t_L g1043 ( 
.A(n_833),
.Y(n_1043)
);

INVx2_ASAP7_75t_L g1044 ( 
.A(n_826),
.Y(n_1044)
);

INVx1_ASAP7_75t_L g1045 ( 
.A(n_830),
.Y(n_1045)
);

NAND2xp5_ASAP7_75t_L g1046 ( 
.A(n_836),
.B(n_613),
.Y(n_1046)
);

INVx1_ASAP7_75t_L g1047 ( 
.A(n_854),
.Y(n_1047)
);

INVx1_ASAP7_75t_L g1048 ( 
.A(n_865),
.Y(n_1048)
);

AOI22xp33_ASAP7_75t_L g1049 ( 
.A1(n_886),
.A2(n_598),
.B1(n_384),
.B2(n_376),
.Y(n_1049)
);

CKINVDCx5p33_ASAP7_75t_R g1050 ( 
.A(n_858),
.Y(n_1050)
);

HB1xp67_ASAP7_75t_L g1051 ( 
.A(n_842),
.Y(n_1051)
);

AND2x2_ASAP7_75t_L g1052 ( 
.A(n_824),
.B(n_575),
.Y(n_1052)
);

NAND2xp5_ASAP7_75t_L g1053 ( 
.A(n_842),
.B(n_732),
.Y(n_1053)
);

AND2x6_ASAP7_75t_SL g1054 ( 
.A(n_849),
.B(n_850),
.Y(n_1054)
);

BUFx3_ASAP7_75t_L g1055 ( 
.A(n_844),
.Y(n_1055)
);

AOI22xp5_ASAP7_75t_L g1056 ( 
.A1(n_849),
.A2(n_732),
.B1(n_309),
.B2(n_310),
.Y(n_1056)
);

INVx1_ASAP7_75t_L g1057 ( 
.A(n_877),
.Y(n_1057)
);

INVx1_ASAP7_75t_L g1058 ( 
.A(n_897),
.Y(n_1058)
);

INVx2_ASAP7_75t_L g1059 ( 
.A(n_874),
.Y(n_1059)
);

INVx2_ASAP7_75t_L g1060 ( 
.A(n_878),
.Y(n_1060)
);

AOI22xp33_ASAP7_75t_L g1061 ( 
.A1(n_850),
.A2(n_386),
.B1(n_373),
.B2(n_726),
.Y(n_1061)
);

AND2x2_ASAP7_75t_L g1062 ( 
.A(n_862),
.B(n_576),
.Y(n_1062)
);

OR2x4_ASAP7_75t_L g1063 ( 
.A(n_862),
.B(n_576),
.Y(n_1063)
);

INVx3_ASAP7_75t_L g1064 ( 
.A(n_883),
.Y(n_1064)
);

AOI22xp33_ASAP7_75t_L g1065 ( 
.A1(n_891),
.A2(n_386),
.B1(n_727),
.B2(n_726),
.Y(n_1065)
);

INVx3_ASAP7_75t_L g1066 ( 
.A(n_884),
.Y(n_1066)
);

AOI22xp33_ASAP7_75t_L g1067 ( 
.A1(n_891),
.A2(n_634),
.B1(n_727),
.B2(n_726),
.Y(n_1067)
);

BUFx3_ASAP7_75t_L g1068 ( 
.A(n_845),
.Y(n_1068)
);

INVx1_ASAP7_75t_L g1069 ( 
.A(n_889),
.Y(n_1069)
);

NAND2xp5_ASAP7_75t_SL g1070 ( 
.A(n_742),
.B(n_732),
.Y(n_1070)
);

INVx1_ASAP7_75t_L g1071 ( 
.A(n_885),
.Y(n_1071)
);

INVx5_ASAP7_75t_L g1072 ( 
.A(n_754),
.Y(n_1072)
);

INVx1_ASAP7_75t_L g1073 ( 
.A(n_847),
.Y(n_1073)
);

INVx1_ASAP7_75t_L g1074 ( 
.A(n_847),
.Y(n_1074)
);

INVx1_ASAP7_75t_SL g1075 ( 
.A(n_846),
.Y(n_1075)
);

AOI22xp33_ASAP7_75t_L g1076 ( 
.A1(n_876),
.A2(n_634),
.B1(n_727),
.B2(n_725),
.Y(n_1076)
);

AND3x2_ASAP7_75t_SL g1077 ( 
.A(n_851),
.B(n_3),
.C(n_4),
.Y(n_1077)
);

NAND2xp5_ASAP7_75t_L g1078 ( 
.A(n_831),
.B(n_619),
.Y(n_1078)
);

INVx4_ASAP7_75t_L g1079 ( 
.A(n_926),
.Y(n_1079)
);

INVx2_ASAP7_75t_L g1080 ( 
.A(n_898),
.Y(n_1080)
);

AOI21xp5_ASAP7_75t_L g1081 ( 
.A1(n_902),
.A2(n_876),
.B(n_761),
.Y(n_1081)
);

BUFx6f_ASAP7_75t_L g1082 ( 
.A(n_926),
.Y(n_1082)
);

NOR2xp33_ASAP7_75t_R g1083 ( 
.A(n_913),
.B(n_220),
.Y(n_1083)
);

BUFx6f_ASAP7_75t_L g1084 ( 
.A(n_926),
.Y(n_1084)
);

AOI21xp5_ASAP7_75t_L g1085 ( 
.A1(n_909),
.A2(n_761),
.B(n_754),
.Y(n_1085)
);

AOI21xp5_ASAP7_75t_L g1086 ( 
.A1(n_998),
.A2(n_770),
.B(n_763),
.Y(n_1086)
);

NAND2xp5_ASAP7_75t_L g1087 ( 
.A(n_1001),
.B(n_763),
.Y(n_1087)
);

AO22x1_ASAP7_75t_L g1088 ( 
.A1(n_908),
.A2(n_314),
.B1(n_322),
.B2(n_325),
.Y(n_1088)
);

INVx2_ASAP7_75t_L g1089 ( 
.A(n_898),
.Y(n_1089)
);

O2A1O1Ixp33_ASAP7_75t_L g1090 ( 
.A1(n_989),
.A2(n_834),
.B(n_797),
.C(n_822),
.Y(n_1090)
);

BUFx2_ASAP7_75t_L g1091 ( 
.A(n_932),
.Y(n_1091)
);

NAND2xp5_ASAP7_75t_L g1092 ( 
.A(n_915),
.B(n_827),
.Y(n_1092)
);

BUFx6f_ASAP7_75t_L g1093 ( 
.A(n_926),
.Y(n_1093)
);

OAI22xp5_ASAP7_75t_SL g1094 ( 
.A1(n_958),
.A2(n_307),
.B1(n_286),
.B2(n_292),
.Y(n_1094)
);

NOR2xp33_ASAP7_75t_L g1095 ( 
.A(n_908),
.B(n_834),
.Y(n_1095)
);

AOI21xp5_ASAP7_75t_L g1096 ( 
.A1(n_998),
.A2(n_852),
.B(n_843),
.Y(n_1096)
);

AOI21xp5_ASAP7_75t_L g1097 ( 
.A1(n_920),
.A2(n_852),
.B(n_843),
.Y(n_1097)
);

INVx2_ASAP7_75t_L g1098 ( 
.A(n_906),
.Y(n_1098)
);

BUFx6f_ASAP7_75t_L g1099 ( 
.A(n_933),
.Y(n_1099)
);

INVx3_ASAP7_75t_L g1100 ( 
.A(n_976),
.Y(n_1100)
);

INVx3_ASAP7_75t_L g1101 ( 
.A(n_976),
.Y(n_1101)
);

AND2x4_ASAP7_75t_L g1102 ( 
.A(n_980),
.B(n_857),
.Y(n_1102)
);

AOI22xp5_ASAP7_75t_L g1103 ( 
.A1(n_1020),
.A2(n_857),
.B1(n_305),
.B2(n_348),
.Y(n_1103)
);

HB1xp67_ASAP7_75t_L g1104 ( 
.A(n_939),
.Y(n_1104)
);

O2A1O1Ixp33_ASAP7_75t_L g1105 ( 
.A1(n_989),
.A2(n_668),
.B(n_663),
.C(n_662),
.Y(n_1105)
);

NAND2xp5_ASAP7_75t_L g1106 ( 
.A(n_1000),
.B(n_619),
.Y(n_1106)
);

INVx2_ASAP7_75t_L g1107 ( 
.A(n_995),
.Y(n_1107)
);

CKINVDCx5p33_ASAP7_75t_R g1108 ( 
.A(n_973),
.Y(n_1108)
);

NOR2xp33_ASAP7_75t_L g1109 ( 
.A(n_1051),
.B(n_295),
.Y(n_1109)
);

INVx1_ASAP7_75t_L g1110 ( 
.A(n_903),
.Y(n_1110)
);

O2A1O1Ixp33_ASAP7_75t_L g1111 ( 
.A1(n_997),
.A2(n_672),
.B(n_668),
.C(n_663),
.Y(n_1111)
);

INVx1_ASAP7_75t_L g1112 ( 
.A(n_911),
.Y(n_1112)
);

AOI21xp5_ASAP7_75t_L g1113 ( 
.A1(n_923),
.A2(n_949),
.B(n_986),
.Y(n_1113)
);

NOR3xp33_ASAP7_75t_SL g1114 ( 
.A(n_1050),
.B(n_306),
.C(n_297),
.Y(n_1114)
);

HB1xp67_ASAP7_75t_L g1115 ( 
.A(n_939),
.Y(n_1115)
);

NAND2xp5_ASAP7_75t_SL g1116 ( 
.A(n_1055),
.B(n_222),
.Y(n_1116)
);

AOI22xp5_ASAP7_75t_L g1117 ( 
.A1(n_901),
.A2(n_304),
.B1(n_303),
.B2(n_299),
.Y(n_1117)
);

OAI22xp5_ASAP7_75t_L g1118 ( 
.A1(n_1029),
.A2(n_391),
.B1(n_311),
.B2(n_323),
.Y(n_1118)
);

BUFx4f_ASAP7_75t_L g1119 ( 
.A(n_985),
.Y(n_1119)
);

INVx4_ASAP7_75t_L g1120 ( 
.A(n_994),
.Y(n_1120)
);

NAND2xp5_ASAP7_75t_L g1121 ( 
.A(n_1002),
.B(n_628),
.Y(n_1121)
);

INVx1_ASAP7_75t_L g1122 ( 
.A(n_918),
.Y(n_1122)
);

AOI21xp5_ASAP7_75t_L g1123 ( 
.A1(n_986),
.A2(n_505),
.B(n_729),
.Y(n_1123)
);

INVx2_ASAP7_75t_L g1124 ( 
.A(n_995),
.Y(n_1124)
);

NOR2xp33_ASAP7_75t_L g1125 ( 
.A(n_1051),
.B(n_328),
.Y(n_1125)
);

AOI22xp33_ASAP7_75t_L g1126 ( 
.A1(n_1039),
.A2(n_222),
.B1(n_377),
.B2(n_379),
.Y(n_1126)
);

NOR2xp33_ASAP7_75t_L g1127 ( 
.A(n_1010),
.B(n_331),
.Y(n_1127)
);

INVx3_ASAP7_75t_L g1128 ( 
.A(n_976),
.Y(n_1128)
);

INVx2_ASAP7_75t_L g1129 ( 
.A(n_1019),
.Y(n_1129)
);

NOR2xp33_ASAP7_75t_L g1130 ( 
.A(n_1010),
.B(n_341),
.Y(n_1130)
);

INVx1_ASAP7_75t_L g1131 ( 
.A(n_921),
.Y(n_1131)
);

NAND2xp5_ASAP7_75t_SL g1132 ( 
.A(n_1055),
.B(n_227),
.Y(n_1132)
);

AO32x2_ASAP7_75t_L g1133 ( 
.A1(n_964),
.A2(n_3),
.A3(n_9),
.B1(n_12),
.B2(n_14),
.Y(n_1133)
);

A2O1A1Ixp33_ASAP7_75t_L g1134 ( 
.A1(n_901),
.A2(n_630),
.B(n_725),
.C(n_724),
.Y(n_1134)
);

BUFx12f_ASAP7_75t_L g1135 ( 
.A(n_928),
.Y(n_1135)
);

A2O1A1Ixp33_ASAP7_75t_L g1136 ( 
.A1(n_1041),
.A2(n_647),
.B(n_724),
.C(n_721),
.Y(n_1136)
);

NOR2xp33_ASAP7_75t_L g1137 ( 
.A(n_1073),
.B(n_343),
.Y(n_1137)
);

INVx1_ASAP7_75t_L g1138 ( 
.A(n_930),
.Y(n_1138)
);

INVx1_ASAP7_75t_L g1139 ( 
.A(n_938),
.Y(n_1139)
);

NOR2xp33_ASAP7_75t_L g1140 ( 
.A(n_1074),
.B(n_344),
.Y(n_1140)
);

INVx1_ASAP7_75t_L g1141 ( 
.A(n_944),
.Y(n_1141)
);

OAI22xp5_ASAP7_75t_L g1142 ( 
.A1(n_1029),
.A2(n_349),
.B1(n_353),
.B2(n_356),
.Y(n_1142)
);

O2A1O1Ixp5_ASAP7_75t_L g1143 ( 
.A1(n_1015),
.A2(n_632),
.B(n_721),
.C(n_720),
.Y(n_1143)
);

INVx2_ASAP7_75t_L g1144 ( 
.A(n_1019),
.Y(n_1144)
);

AOI22xp33_ASAP7_75t_L g1145 ( 
.A1(n_1039),
.A2(n_227),
.B1(n_298),
.B2(n_367),
.Y(n_1145)
);

BUFx12f_ASAP7_75t_L g1146 ( 
.A(n_975),
.Y(n_1146)
);

NOR2xp33_ASAP7_75t_L g1147 ( 
.A(n_1004),
.B(n_298),
.Y(n_1147)
);

AOI21xp5_ASAP7_75t_L g1148 ( 
.A1(n_940),
.A2(n_942),
.B(n_1046),
.Y(n_1148)
);

NOR2xp33_ASAP7_75t_SL g1149 ( 
.A(n_913),
.B(n_367),
.Y(n_1149)
);

NOR2xp33_ASAP7_75t_L g1150 ( 
.A(n_1068),
.B(n_375),
.Y(n_1150)
);

NAND2xp5_ASAP7_75t_SL g1151 ( 
.A(n_1068),
.B(n_375),
.Y(n_1151)
);

BUFx6f_ASAP7_75t_L g1152 ( 
.A(n_933),
.Y(n_1152)
);

NAND2xp5_ASAP7_75t_SL g1153 ( 
.A(n_917),
.B(n_377),
.Y(n_1153)
);

INVx2_ASAP7_75t_SL g1154 ( 
.A(n_991),
.Y(n_1154)
);

NOR2xp33_ASAP7_75t_SL g1155 ( 
.A(n_1035),
.B(n_379),
.Y(n_1155)
);

NOR2xp33_ASAP7_75t_L g1156 ( 
.A(n_996),
.B(n_380),
.Y(n_1156)
);

OAI22xp5_ASAP7_75t_L g1157 ( 
.A1(n_1041),
.A2(n_385),
.B1(n_382),
.B2(n_380),
.Y(n_1157)
);

A2O1A1Ixp33_ASAP7_75t_SL g1158 ( 
.A1(n_934),
.A2(n_640),
.B(n_721),
.C(n_720),
.Y(n_1158)
);

BUFx2_ASAP7_75t_L g1159 ( 
.A(n_932),
.Y(n_1159)
);

CKINVDCx16_ASAP7_75t_R g1160 ( 
.A(n_904),
.Y(n_1160)
);

INVx2_ASAP7_75t_L g1161 ( 
.A(n_937),
.Y(n_1161)
);

INVx2_ASAP7_75t_L g1162 ( 
.A(n_953),
.Y(n_1162)
);

BUFx6f_ASAP7_75t_L g1163 ( 
.A(n_943),
.Y(n_1163)
);

OAI21xp5_ASAP7_75t_L g1164 ( 
.A1(n_1017),
.A2(n_640),
.B(n_720),
.Y(n_1164)
);

CKINVDCx5p33_ASAP7_75t_R g1165 ( 
.A(n_904),
.Y(n_1165)
);

A2O1A1Ixp33_ASAP7_75t_L g1166 ( 
.A1(n_907),
.A2(n_686),
.B(n_673),
.C(n_677),
.Y(n_1166)
);

NAND2xp5_ASAP7_75t_SL g1167 ( 
.A(n_941),
.B(n_382),
.Y(n_1167)
);

OAI22xp5_ASAP7_75t_L g1168 ( 
.A1(n_1008),
.A2(n_385),
.B1(n_389),
.B2(n_581),
.Y(n_1168)
);

HB1xp67_ASAP7_75t_L g1169 ( 
.A(n_945),
.Y(n_1169)
);

INVx3_ASAP7_75t_SL g1170 ( 
.A(n_985),
.Y(n_1170)
);

AOI21xp5_ASAP7_75t_L g1171 ( 
.A1(n_1012),
.A2(n_729),
.B(n_648),
.Y(n_1171)
);

INVx3_ASAP7_75t_L g1172 ( 
.A(n_976),
.Y(n_1172)
);

NOR3xp33_ASAP7_75t_SL g1173 ( 
.A(n_934),
.B(n_389),
.C(n_308),
.Y(n_1173)
);

INVx1_ASAP7_75t_L g1174 ( 
.A(n_955),
.Y(n_1174)
);

OAI22xp5_ASAP7_75t_L g1175 ( 
.A1(n_907),
.A2(n_580),
.B1(n_703),
.B2(n_630),
.Y(n_1175)
);

NAND2xp5_ASAP7_75t_SL g1176 ( 
.A(n_931),
.B(n_288),
.Y(n_1176)
);

AOI21xp5_ASAP7_75t_L g1177 ( 
.A1(n_984),
.A2(n_729),
.B(n_648),
.Y(n_1177)
);

AND2x2_ASAP7_75t_L g1178 ( 
.A(n_1005),
.B(n_321),
.Y(n_1178)
);

AND2x4_ASAP7_75t_L g1179 ( 
.A(n_980),
.B(n_632),
.Y(n_1179)
);

NAND2xp5_ASAP7_75t_L g1180 ( 
.A(n_1069),
.B(n_634),
.Y(n_1180)
);

NAND2xp5_ASAP7_75t_L g1181 ( 
.A(n_1059),
.B(n_636),
.Y(n_1181)
);

NAND2xp5_ASAP7_75t_SL g1182 ( 
.A(n_977),
.B(n_332),
.Y(n_1182)
);

BUFx2_ASAP7_75t_L g1183 ( 
.A(n_981),
.Y(n_1183)
);

BUFx2_ASAP7_75t_L g1184 ( 
.A(n_981),
.Y(n_1184)
);

BUFx6f_ASAP7_75t_L g1185 ( 
.A(n_943),
.Y(n_1185)
);

INVx2_ASAP7_75t_L g1186 ( 
.A(n_963),
.Y(n_1186)
);

NAND2xp5_ASAP7_75t_L g1187 ( 
.A(n_1060),
.B(n_1042),
.Y(n_1187)
);

NAND2xp5_ASAP7_75t_L g1188 ( 
.A(n_1042),
.B(n_1062),
.Y(n_1188)
);

NAND2xp5_ASAP7_75t_L g1189 ( 
.A(n_1022),
.B(n_636),
.Y(n_1189)
);

O2A1O1Ixp33_ASAP7_75t_L g1190 ( 
.A1(n_997),
.A2(n_668),
.B(n_636),
.C(n_640),
.Y(n_1190)
);

INVx5_ASAP7_75t_L g1191 ( 
.A(n_982),
.Y(n_1191)
);

INVx1_ASAP7_75t_L g1192 ( 
.A(n_974),
.Y(n_1192)
);

AOI21xp5_ASAP7_75t_L g1193 ( 
.A1(n_992),
.A2(n_729),
.B(n_648),
.Y(n_1193)
);

INVx5_ASAP7_75t_L g1194 ( 
.A(n_982),
.Y(n_1194)
);

INVx2_ASAP7_75t_L g1195 ( 
.A(n_1018),
.Y(n_1195)
);

INVx2_ASAP7_75t_L g1196 ( 
.A(n_1036),
.Y(n_1196)
);

INVx2_ASAP7_75t_L g1197 ( 
.A(n_1037),
.Y(n_1197)
);

OR2x6_ASAP7_75t_SL g1198 ( 
.A(n_965),
.B(n_642),
.Y(n_1198)
);

AOI22xp5_ASAP7_75t_L g1199 ( 
.A1(n_1006),
.A2(n_717),
.B1(n_710),
.B2(n_703),
.Y(n_1199)
);

OAI21xp5_ASAP7_75t_L g1200 ( 
.A1(n_948),
.A2(n_717),
.B(n_710),
.Y(n_1200)
);

NOR2xp33_ASAP7_75t_L g1201 ( 
.A(n_967),
.B(n_644),
.Y(n_1201)
);

OAI22xp5_ASAP7_75t_L g1202 ( 
.A1(n_1063),
.A2(n_717),
.B1(n_703),
.B2(n_698),
.Y(n_1202)
);

AOI22xp33_ASAP7_75t_L g1203 ( 
.A1(n_910),
.A2(n_698),
.B1(n_686),
.B2(n_684),
.Y(n_1203)
);

INVx2_ASAP7_75t_L g1204 ( 
.A(n_1044),
.Y(n_1204)
);

HB1xp67_ASAP7_75t_L g1205 ( 
.A(n_945),
.Y(n_1205)
);

CKINVDCx10_ASAP7_75t_R g1206 ( 
.A(n_927),
.Y(n_1206)
);

NAND2xp5_ASAP7_75t_L g1207 ( 
.A(n_1015),
.B(n_644),
.Y(n_1207)
);

INVx1_ASAP7_75t_L g1208 ( 
.A(n_960),
.Y(n_1208)
);

INVx1_ASAP7_75t_L g1209 ( 
.A(n_960),
.Y(n_1209)
);

NAND2xp5_ASAP7_75t_SL g1210 ( 
.A(n_977),
.B(n_644),
.Y(n_1210)
);

AOI21xp5_ASAP7_75t_L g1211 ( 
.A1(n_979),
.A2(n_648),
.B(n_675),
.Y(n_1211)
);

NAND3xp33_ASAP7_75t_SL g1212 ( 
.A(n_1023),
.B(n_1034),
.C(n_1075),
.Y(n_1212)
);

NOR2xp33_ASAP7_75t_L g1213 ( 
.A(n_947),
.B(n_646),
.Y(n_1213)
);

AOI22xp33_ASAP7_75t_L g1214 ( 
.A1(n_910),
.A2(n_1071),
.B1(n_1052),
.B2(n_990),
.Y(n_1214)
);

AOI22xp33_ASAP7_75t_L g1215 ( 
.A1(n_990),
.A2(n_684),
.B1(n_677),
.B2(n_646),
.Y(n_1215)
);

AND2x2_ASAP7_75t_L g1216 ( 
.A(n_966),
.B(n_647),
.Y(n_1216)
);

NOR2xp33_ASAP7_75t_L g1217 ( 
.A(n_1063),
.B(n_647),
.Y(n_1217)
);

INVxp67_ASAP7_75t_L g1218 ( 
.A(n_912),
.Y(n_1218)
);

INVx1_ASAP7_75t_L g1219 ( 
.A(n_1014),
.Y(n_1219)
);

INVx1_ASAP7_75t_L g1220 ( 
.A(n_1021),
.Y(n_1220)
);

NAND2xp5_ASAP7_75t_L g1221 ( 
.A(n_1064),
.B(n_657),
.Y(n_1221)
);

NAND2xp5_ASAP7_75t_L g1222 ( 
.A(n_1064),
.B(n_657),
.Y(n_1222)
);

NAND2xp5_ASAP7_75t_L g1223 ( 
.A(n_1066),
.B(n_657),
.Y(n_1223)
);

OAI22xp5_ASAP7_75t_L g1224 ( 
.A1(n_1072),
.A2(n_662),
.B1(n_663),
.B2(n_672),
.Y(n_1224)
);

OAI22xp5_ASAP7_75t_L g1225 ( 
.A1(n_1072),
.A2(n_662),
.B1(n_672),
.B2(n_673),
.Y(n_1225)
);

INVx8_ASAP7_75t_L g1226 ( 
.A(n_1191),
.Y(n_1226)
);

OAI21x1_ASAP7_75t_L g1227 ( 
.A1(n_1113),
.A2(n_1070),
.B(n_987),
.Y(n_1227)
);

OAI21x1_ASAP7_75t_L g1228 ( 
.A1(n_1085),
.A2(n_1070),
.B(n_987),
.Y(n_1228)
);

INVx2_ASAP7_75t_SL g1229 ( 
.A(n_1119),
.Y(n_1229)
);

NAND2xp5_ASAP7_75t_L g1230 ( 
.A(n_1188),
.B(n_1187),
.Y(n_1230)
);

BUFx4f_ASAP7_75t_L g1231 ( 
.A(n_1146),
.Y(n_1231)
);

NAND2x1_ASAP7_75t_L g1232 ( 
.A(n_1120),
.B(n_982),
.Y(n_1232)
);

AOI21xp5_ASAP7_75t_L g1233 ( 
.A1(n_1092),
.A2(n_1053),
.B(n_1011),
.Y(n_1233)
);

OAI21xp5_ASAP7_75t_L g1234 ( 
.A1(n_1148),
.A2(n_1007),
.B(n_1040),
.Y(n_1234)
);

NOR2xp33_ASAP7_75t_L g1235 ( 
.A(n_1155),
.B(n_1054),
.Y(n_1235)
);

NOR2xp33_ASAP7_75t_L g1236 ( 
.A(n_1155),
.B(n_1028),
.Y(n_1236)
);

AND2x4_ASAP7_75t_L g1237 ( 
.A(n_1120),
.B(n_1099),
.Y(n_1237)
);

AO31x2_ASAP7_75t_L g1238 ( 
.A1(n_1224),
.A2(n_999),
.A3(n_993),
.B(n_1009),
.Y(n_1238)
);

HB1xp67_ASAP7_75t_L g1239 ( 
.A(n_1104),
.Y(n_1239)
);

INVx1_ASAP7_75t_L g1240 ( 
.A(n_1110),
.Y(n_1240)
);

AO31x2_ASAP7_75t_L g1241 ( 
.A1(n_1224),
.A2(n_999),
.A3(n_993),
.B(n_1078),
.Y(n_1241)
);

INVx2_ASAP7_75t_L g1242 ( 
.A(n_1080),
.Y(n_1242)
);

INVx5_ASAP7_75t_L g1243 ( 
.A(n_1082),
.Y(n_1243)
);

INVx1_ASAP7_75t_L g1244 ( 
.A(n_1112),
.Y(n_1244)
);

OAI21x1_ASAP7_75t_L g1245 ( 
.A1(n_1081),
.A2(n_1040),
.B(n_1024),
.Y(n_1245)
);

AOI21xp5_ASAP7_75t_L g1246 ( 
.A1(n_1092),
.A2(n_950),
.B(n_968),
.Y(n_1246)
);

A2O1A1Ixp33_ASAP7_75t_L g1247 ( 
.A1(n_1095),
.A2(n_1127),
.B(n_1130),
.C(n_1090),
.Y(n_1247)
);

INVx1_ASAP7_75t_L g1248 ( 
.A(n_1122),
.Y(n_1248)
);

NAND2xp5_ASAP7_75t_L g1249 ( 
.A(n_1187),
.B(n_1066),
.Y(n_1249)
);

OAI21x1_ASAP7_75t_L g1250 ( 
.A1(n_1143),
.A2(n_983),
.B(n_1038),
.Y(n_1250)
);

AO31x2_ASAP7_75t_L g1251 ( 
.A1(n_1225),
.A2(n_969),
.A3(n_924),
.B(n_925),
.Y(n_1251)
);

INVxp67_ASAP7_75t_L g1252 ( 
.A(n_1115),
.Y(n_1252)
);

OAI21x1_ASAP7_75t_L g1253 ( 
.A1(n_1164),
.A2(n_1038),
.B(n_1030),
.Y(n_1253)
);

AND2x2_ASAP7_75t_L g1254 ( 
.A(n_1178),
.B(n_956),
.Y(n_1254)
);

NAND2xp5_ASAP7_75t_L g1255 ( 
.A(n_1214),
.B(n_1208),
.Y(n_1255)
);

BUFx3_ASAP7_75t_L g1256 ( 
.A(n_1135),
.Y(n_1256)
);

AND2x4_ASAP7_75t_L g1257 ( 
.A(n_1099),
.B(n_957),
.Y(n_1257)
);

NAND2xp5_ASAP7_75t_L g1258 ( 
.A(n_1209),
.B(n_1137),
.Y(n_1258)
);

OAI22x1_ASAP7_75t_L g1259 ( 
.A1(n_1170),
.A2(n_922),
.B1(n_1159),
.B2(n_1091),
.Y(n_1259)
);

INVx1_ASAP7_75t_L g1260 ( 
.A(n_1131),
.Y(n_1260)
);

CKINVDCx6p67_ASAP7_75t_R g1261 ( 
.A(n_1160),
.Y(n_1261)
);

AOI21xp5_ASAP7_75t_L g1262 ( 
.A1(n_1097),
.A2(n_950),
.B(n_1072),
.Y(n_1262)
);

NOR2xp67_ASAP7_75t_SL g1263 ( 
.A(n_1108),
.B(n_951),
.Y(n_1263)
);

CKINVDCx11_ASAP7_75t_R g1264 ( 
.A(n_1099),
.Y(n_1264)
);

A2O1A1Ixp33_ASAP7_75t_L g1265 ( 
.A1(n_1217),
.A2(n_1032),
.B(n_962),
.C(n_1056),
.Y(n_1265)
);

NOR2xp33_ASAP7_75t_L g1266 ( 
.A(n_1150),
.B(n_957),
.Y(n_1266)
);

AO31x2_ASAP7_75t_L g1267 ( 
.A1(n_1225),
.A2(n_929),
.A3(n_946),
.B(n_959),
.Y(n_1267)
);

OAI21xp5_ASAP7_75t_SL g1268 ( 
.A1(n_1126),
.A2(n_1049),
.B(n_1061),
.Y(n_1268)
);

NOR2xp33_ASAP7_75t_R g1269 ( 
.A(n_1165),
.B(n_935),
.Y(n_1269)
);

AND3x2_ASAP7_75t_L g1270 ( 
.A(n_1149),
.B(n_905),
.C(n_1077),
.Y(n_1270)
);

INVx5_ASAP7_75t_L g1271 ( 
.A(n_1082),
.Y(n_1271)
);

O2A1O1Ixp33_ASAP7_75t_L g1272 ( 
.A1(n_1118),
.A2(n_952),
.B(n_927),
.C(n_1049),
.Y(n_1272)
);

OAI22x1_ASAP7_75t_L g1273 ( 
.A1(n_1183),
.A2(n_1077),
.B1(n_905),
.B2(n_1043),
.Y(n_1273)
);

OAI22xp5_ASAP7_75t_L g1274 ( 
.A1(n_1145),
.A2(n_1072),
.B1(n_948),
.B2(n_971),
.Y(n_1274)
);

NAND2xp5_ASAP7_75t_L g1275 ( 
.A(n_1140),
.B(n_972),
.Y(n_1275)
);

OAI21x1_ASAP7_75t_L g1276 ( 
.A1(n_1177),
.A2(n_1067),
.B(n_1076),
.Y(n_1276)
);

OAI22x1_ASAP7_75t_L g1277 ( 
.A1(n_1184),
.A2(n_988),
.B1(n_952),
.B2(n_1023),
.Y(n_1277)
);

O2A1O1Ixp5_ASAP7_75t_SL g1278 ( 
.A1(n_1175),
.A2(n_954),
.B(n_1045),
.C(n_1026),
.Y(n_1278)
);

AOI221x1_ASAP7_75t_L g1279 ( 
.A1(n_1118),
.A2(n_1142),
.B1(n_1157),
.B2(n_1175),
.C(n_1207),
.Y(n_1279)
);

NAND2xp5_ASAP7_75t_L g1280 ( 
.A(n_1147),
.B(n_900),
.Y(n_1280)
);

INVx1_ASAP7_75t_L g1281 ( 
.A(n_1138),
.Y(n_1281)
);

NAND3xp33_ASAP7_75t_SL g1282 ( 
.A(n_1117),
.B(n_1061),
.C(n_1065),
.Y(n_1282)
);

AOI221x1_ASAP7_75t_L g1283 ( 
.A1(n_1142),
.A2(n_1047),
.B1(n_1048),
.B2(n_1057),
.C(n_1058),
.Y(n_1283)
);

NAND3x1_ASAP7_75t_L g1284 ( 
.A(n_1213),
.B(n_899),
.C(n_916),
.Y(n_1284)
);

OAI22xp5_ASAP7_75t_L g1285 ( 
.A1(n_1087),
.A2(n_971),
.B1(n_1003),
.B2(n_970),
.Y(n_1285)
);

INVx1_ASAP7_75t_L g1286 ( 
.A(n_1139),
.Y(n_1286)
);

OR2x2_ASAP7_75t_L g1287 ( 
.A(n_1169),
.B(n_1205),
.Y(n_1287)
);

AND2x4_ASAP7_75t_L g1288 ( 
.A(n_1152),
.B(n_927),
.Y(n_1288)
);

AND2x2_ASAP7_75t_L g1289 ( 
.A(n_1109),
.B(n_971),
.Y(n_1289)
);

NAND2xp5_ASAP7_75t_L g1290 ( 
.A(n_1201),
.B(n_900),
.Y(n_1290)
);

OAI22xp5_ASAP7_75t_L g1291 ( 
.A1(n_1103),
.A2(n_935),
.B1(n_1031),
.B2(n_1027),
.Y(n_1291)
);

NAND2xp5_ASAP7_75t_L g1292 ( 
.A(n_1125),
.B(n_900),
.Y(n_1292)
);

NAND2xp5_ASAP7_75t_L g1293 ( 
.A(n_1192),
.B(n_900),
.Y(n_1293)
);

OAI22x1_ASAP7_75t_L g1294 ( 
.A1(n_1116),
.A2(n_1013),
.B1(n_954),
.B2(n_961),
.Y(n_1294)
);

AOI21xp5_ASAP7_75t_L g1295 ( 
.A1(n_1096),
.A2(n_978),
.B(n_961),
.Y(n_1295)
);

INVx1_ASAP7_75t_L g1296 ( 
.A(n_1141),
.Y(n_1296)
);

AO31x2_ASAP7_75t_L g1297 ( 
.A1(n_1134),
.A2(n_919),
.A3(n_914),
.B(n_673),
.Y(n_1297)
);

INVx2_ASAP7_75t_L g1298 ( 
.A(n_1089),
.Y(n_1298)
);

OAI21x1_ASAP7_75t_L g1299 ( 
.A1(n_1193),
.A2(n_1200),
.B(n_1171),
.Y(n_1299)
);

AND2x2_ASAP7_75t_L g1300 ( 
.A(n_1114),
.B(n_1156),
.Y(n_1300)
);

AO22x2_ASAP7_75t_L g1301 ( 
.A1(n_1157),
.A2(n_1133),
.B1(n_1212),
.B2(n_1153),
.Y(n_1301)
);

INVxp67_ASAP7_75t_SL g1302 ( 
.A(n_1082),
.Y(n_1302)
);

AOI21xp5_ASAP7_75t_SL g1303 ( 
.A1(n_1102),
.A2(n_1025),
.B(n_982),
.Y(n_1303)
);

INVx1_ASAP7_75t_L g1304 ( 
.A(n_1174),
.Y(n_1304)
);

AND2x2_ASAP7_75t_L g1305 ( 
.A(n_1154),
.B(n_1216),
.Y(n_1305)
);

AOI21xp5_ASAP7_75t_L g1306 ( 
.A1(n_1086),
.A2(n_1016),
.B(n_1025),
.Y(n_1306)
);

OR2x2_ASAP7_75t_L g1307 ( 
.A(n_1132),
.B(n_916),
.Y(n_1307)
);

NAND2xp5_ASAP7_75t_SL g1308 ( 
.A(n_1152),
.B(n_936),
.Y(n_1308)
);

INVx2_ASAP7_75t_L g1309 ( 
.A(n_1098),
.Y(n_1309)
);

OAI21xp5_ASAP7_75t_L g1310 ( 
.A1(n_1166),
.A2(n_1003),
.B(n_970),
.Y(n_1310)
);

AO21x2_ASAP7_75t_L g1311 ( 
.A1(n_1158),
.A2(n_1033),
.B(n_936),
.Y(n_1311)
);

AOI22xp5_ASAP7_75t_L g1312 ( 
.A1(n_1094),
.A2(n_994),
.B1(n_514),
.B2(n_370),
.Y(n_1312)
);

NAND2xp5_ASAP7_75t_L g1313 ( 
.A(n_1088),
.B(n_9),
.Y(n_1313)
);

INVx1_ASAP7_75t_L g1314 ( 
.A(n_1107),
.Y(n_1314)
);

INVx2_ASAP7_75t_L g1315 ( 
.A(n_1124),
.Y(n_1315)
);

OAI21xp5_ASAP7_75t_L g1316 ( 
.A1(n_1136),
.A2(n_514),
.B(n_83),
.Y(n_1316)
);

HB1xp67_ASAP7_75t_L g1317 ( 
.A(n_1152),
.Y(n_1317)
);

OAI21x1_ASAP7_75t_L g1318 ( 
.A1(n_1123),
.A2(n_75),
.B(n_88),
.Y(n_1318)
);

NAND2xp5_ASAP7_75t_L g1319 ( 
.A(n_1219),
.B(n_12),
.Y(n_1319)
);

INVx1_ASAP7_75t_L g1320 ( 
.A(n_1129),
.Y(n_1320)
);

INVx3_ASAP7_75t_SL g1321 ( 
.A(n_1163),
.Y(n_1321)
);

O2A1O1Ixp33_ASAP7_75t_L g1322 ( 
.A1(n_1151),
.A2(n_16),
.B(n_17),
.C(n_18),
.Y(n_1322)
);

OAI21x1_ASAP7_75t_L g1323 ( 
.A1(n_1211),
.A2(n_114),
.B(n_107),
.Y(n_1323)
);

AOI21xp5_ASAP7_75t_L g1324 ( 
.A1(n_1121),
.A2(n_675),
.B(n_648),
.Y(n_1324)
);

INVx2_ASAP7_75t_L g1325 ( 
.A(n_1144),
.Y(n_1325)
);

A2O1A1Ixp33_ASAP7_75t_L g1326 ( 
.A1(n_1173),
.A2(n_16),
.B(n_19),
.C(n_20),
.Y(n_1326)
);

NOR2xp67_ASAP7_75t_L g1327 ( 
.A(n_1191),
.B(n_1194),
.Y(n_1327)
);

INVxp67_ASAP7_75t_SL g1328 ( 
.A(n_1084),
.Y(n_1328)
);

NAND2xp5_ASAP7_75t_L g1329 ( 
.A(n_1220),
.B(n_21),
.Y(n_1329)
);

AO31x2_ASAP7_75t_L g1330 ( 
.A1(n_1202),
.A2(n_1121),
.A3(n_1221),
.B(n_1180),
.Y(n_1330)
);

INVx2_ASAP7_75t_L g1331 ( 
.A(n_1161),
.Y(n_1331)
);

A2O1A1Ixp33_ASAP7_75t_L g1332 ( 
.A1(n_1105),
.A2(n_22),
.B(n_23),
.C(n_30),
.Y(n_1332)
);

AOI21xp5_ASAP7_75t_L g1333 ( 
.A1(n_1106),
.A2(n_675),
.B(n_514),
.Y(n_1333)
);

BUFx2_ASAP7_75t_L g1334 ( 
.A(n_1163),
.Y(n_1334)
);

AO21x2_ASAP7_75t_L g1335 ( 
.A1(n_1202),
.A2(n_128),
.B(n_192),
.Y(n_1335)
);

A2O1A1Ixp33_ASAP7_75t_L g1336 ( 
.A1(n_1111),
.A2(n_33),
.B(n_34),
.C(n_39),
.Y(n_1336)
);

INVx3_ASAP7_75t_L g1337 ( 
.A(n_1191),
.Y(n_1337)
);

NAND3xp33_ASAP7_75t_L g1338 ( 
.A(n_1149),
.B(n_33),
.C(n_41),
.Y(n_1338)
);

INVx1_ASAP7_75t_L g1339 ( 
.A(n_1162),
.Y(n_1339)
);

INVx1_ASAP7_75t_L g1340 ( 
.A(n_1186),
.Y(n_1340)
);

NAND2xp33_ASAP7_75t_R g1341 ( 
.A(n_1083),
.B(n_131),
.Y(n_1341)
);

AO21x1_ASAP7_75t_L g1342 ( 
.A1(n_1190),
.A2(n_42),
.B(n_49),
.Y(n_1342)
);

NAND2x1p5_ASAP7_75t_L g1343 ( 
.A(n_1191),
.B(n_1194),
.Y(n_1343)
);

OAI21x1_ASAP7_75t_L g1344 ( 
.A1(n_1221),
.A2(n_137),
.B(n_182),
.Y(n_1344)
);

NAND3xp33_ASAP7_75t_SL g1345 ( 
.A(n_1167),
.B(n_51),
.C(n_52),
.Y(n_1345)
);

AND2x4_ASAP7_75t_L g1346 ( 
.A(n_1163),
.B(n_121),
.Y(n_1346)
);

NAND2xp5_ASAP7_75t_L g1347 ( 
.A(n_1181),
.B(n_52),
.Y(n_1347)
);

O2A1O1Ixp5_ASAP7_75t_SL g1348 ( 
.A1(n_1168),
.A2(n_53),
.B(n_57),
.C(n_58),
.Y(n_1348)
);

NAND2xp5_ASAP7_75t_L g1349 ( 
.A(n_1181),
.B(n_53),
.Y(n_1349)
);

OAI21x1_ASAP7_75t_L g1350 ( 
.A1(n_1222),
.A2(n_152),
.B(n_171),
.Y(n_1350)
);

NOR2xp33_ASAP7_75t_L g1351 ( 
.A(n_1176),
.B(n_57),
.Y(n_1351)
);

AOI21xp5_ASAP7_75t_SL g1352 ( 
.A1(n_1084),
.A2(n_178),
.B(n_169),
.Y(n_1352)
);

O2A1O1Ixp5_ASAP7_75t_L g1353 ( 
.A1(n_1182),
.A2(n_58),
.B(n_59),
.C(n_63),
.Y(n_1353)
);

BUFx6f_ASAP7_75t_L g1354 ( 
.A(n_1185),
.Y(n_1354)
);

INVx2_ASAP7_75t_SL g1355 ( 
.A(n_1185),
.Y(n_1355)
);

AOI22xp5_ASAP7_75t_L g1356 ( 
.A1(n_1168),
.A2(n_59),
.B1(n_64),
.B2(n_66),
.Y(n_1356)
);

OAI21x1_ASAP7_75t_L g1357 ( 
.A1(n_1223),
.A2(n_157),
.B(n_160),
.Y(n_1357)
);

INVx1_ASAP7_75t_L g1358 ( 
.A(n_1195),
.Y(n_1358)
);

INVxp67_ASAP7_75t_L g1359 ( 
.A(n_1198),
.Y(n_1359)
);

OAI21xp33_ASAP7_75t_L g1360 ( 
.A1(n_1218),
.A2(n_64),
.B(n_67),
.Y(n_1360)
);

INVx6_ASAP7_75t_L g1361 ( 
.A(n_1194),
.Y(n_1361)
);

AND2x6_ASAP7_75t_L g1362 ( 
.A(n_1084),
.B(n_161),
.Y(n_1362)
);

BUFx6f_ASAP7_75t_L g1363 ( 
.A(n_1093),
.Y(n_1363)
);

AOI21xp5_ASAP7_75t_L g1364 ( 
.A1(n_1194),
.A2(n_67),
.B(n_1189),
.Y(n_1364)
);

OAI21x1_ASAP7_75t_L g1365 ( 
.A1(n_1199),
.A2(n_1203),
.B(n_1215),
.Y(n_1365)
);

AND2x2_ASAP7_75t_L g1366 ( 
.A(n_1196),
.B(n_1197),
.Y(n_1366)
);

OAI21x1_ASAP7_75t_L g1367 ( 
.A1(n_1210),
.A2(n_1128),
.B(n_1172),
.Y(n_1367)
);

OAI21xp5_ASAP7_75t_L g1368 ( 
.A1(n_1204),
.A2(n_1128),
.B(n_1100),
.Y(n_1368)
);

INVx2_ASAP7_75t_L g1369 ( 
.A(n_1100),
.Y(n_1369)
);

INVx1_ASAP7_75t_L g1370 ( 
.A(n_1093),
.Y(n_1370)
);

OR2x2_ASAP7_75t_L g1371 ( 
.A(n_1179),
.B(n_1101),
.Y(n_1371)
);

AO21x1_ASAP7_75t_L g1372 ( 
.A1(n_1079),
.A2(n_1133),
.B(n_1093),
.Y(n_1372)
);

AO21x2_ASAP7_75t_L g1373 ( 
.A1(n_1133),
.A2(n_1079),
.B(n_1206),
.Y(n_1373)
);

OR2x6_ASAP7_75t_L g1374 ( 
.A(n_1120),
.B(n_904),
.Y(n_1374)
);

BUFx12f_ASAP7_75t_L g1375 ( 
.A(n_1146),
.Y(n_1375)
);

AOI21xp5_ASAP7_75t_L g1376 ( 
.A1(n_1113),
.A2(n_909),
.B(n_902),
.Y(n_1376)
);

OAI22xp33_ASAP7_75t_L g1377 ( 
.A1(n_1155),
.A2(n_712),
.B1(n_735),
.B2(n_1050),
.Y(n_1377)
);

OAI21xp5_ASAP7_75t_L g1378 ( 
.A1(n_1148),
.A2(n_1095),
.B(n_907),
.Y(n_1378)
);

BUFx6f_ASAP7_75t_L g1379 ( 
.A(n_1099),
.Y(n_1379)
);

BUFx6f_ASAP7_75t_L g1380 ( 
.A(n_1226),
.Y(n_1380)
);

OA21x2_ASAP7_75t_L g1381 ( 
.A1(n_1299),
.A2(n_1283),
.B(n_1378),
.Y(n_1381)
);

NAND2x1p5_ASAP7_75t_L g1382 ( 
.A(n_1327),
.B(n_1337),
.Y(n_1382)
);

INVx2_ASAP7_75t_L g1383 ( 
.A(n_1315),
.Y(n_1383)
);

AND2x4_ASAP7_75t_L g1384 ( 
.A(n_1288),
.B(n_1371),
.Y(n_1384)
);

OAI21xp5_ASAP7_75t_L g1385 ( 
.A1(n_1247),
.A2(n_1275),
.B(n_1282),
.Y(n_1385)
);

INVx1_ASAP7_75t_L g1386 ( 
.A(n_1240),
.Y(n_1386)
);

AND2x2_ASAP7_75t_L g1387 ( 
.A(n_1305),
.B(n_1289),
.Y(n_1387)
);

INVx2_ASAP7_75t_SL g1388 ( 
.A(n_1354),
.Y(n_1388)
);

OAI21x1_ASAP7_75t_L g1389 ( 
.A1(n_1245),
.A2(n_1295),
.B(n_1306),
.Y(n_1389)
);

OAI21x1_ASAP7_75t_L g1390 ( 
.A1(n_1250),
.A2(n_1323),
.B(n_1324),
.Y(n_1390)
);

AND2x2_ASAP7_75t_L g1391 ( 
.A(n_1254),
.B(n_1366),
.Y(n_1391)
);

OAI21x1_ASAP7_75t_L g1392 ( 
.A1(n_1262),
.A2(n_1276),
.B(n_1318),
.Y(n_1392)
);

OAI21x1_ASAP7_75t_L g1393 ( 
.A1(n_1234),
.A2(n_1278),
.B(n_1253),
.Y(n_1393)
);

AOI22xp33_ASAP7_75t_L g1394 ( 
.A1(n_1360),
.A2(n_1356),
.B1(n_1338),
.B2(n_1345),
.Y(n_1394)
);

INVx2_ASAP7_75t_L g1395 ( 
.A(n_1325),
.Y(n_1395)
);

BUFx2_ASAP7_75t_L g1396 ( 
.A(n_1257),
.Y(n_1396)
);

INVx2_ASAP7_75t_L g1397 ( 
.A(n_1242),
.Y(n_1397)
);

NOR2xp33_ASAP7_75t_L g1398 ( 
.A(n_1377),
.B(n_1268),
.Y(n_1398)
);

NAND2x1p5_ASAP7_75t_L g1399 ( 
.A(n_1327),
.B(n_1337),
.Y(n_1399)
);

NAND2x1p5_ASAP7_75t_L g1400 ( 
.A(n_1243),
.B(n_1271),
.Y(n_1400)
);

OR2x2_ASAP7_75t_L g1401 ( 
.A(n_1287),
.B(n_1230),
.Y(n_1401)
);

AND2x4_ASAP7_75t_L g1402 ( 
.A(n_1288),
.B(n_1369),
.Y(n_1402)
);

CKINVDCx5p33_ASAP7_75t_R g1403 ( 
.A(n_1264),
.Y(n_1403)
);

AND2x2_ASAP7_75t_L g1404 ( 
.A(n_1266),
.B(n_1258),
.Y(n_1404)
);

OAI21x1_ASAP7_75t_L g1405 ( 
.A1(n_1344),
.A2(n_1357),
.B(n_1350),
.Y(n_1405)
);

AOI22xp33_ASAP7_75t_L g1406 ( 
.A1(n_1360),
.A2(n_1356),
.B1(n_1338),
.B2(n_1313),
.Y(n_1406)
);

BUFx6f_ASAP7_75t_L g1407 ( 
.A(n_1226),
.Y(n_1407)
);

OAI21x1_ASAP7_75t_L g1408 ( 
.A1(n_1233),
.A2(n_1378),
.B(n_1246),
.Y(n_1408)
);

INVx1_ASAP7_75t_L g1409 ( 
.A(n_1244),
.Y(n_1409)
);

BUFx6f_ASAP7_75t_L g1410 ( 
.A(n_1226),
.Y(n_1410)
);

INVx1_ASAP7_75t_L g1411 ( 
.A(n_1248),
.Y(n_1411)
);

INVx2_ASAP7_75t_L g1412 ( 
.A(n_1298),
.Y(n_1412)
);

INVx1_ASAP7_75t_L g1413 ( 
.A(n_1260),
.Y(n_1413)
);

AND2x2_ASAP7_75t_L g1414 ( 
.A(n_1300),
.B(n_1359),
.Y(n_1414)
);

CKINVDCx11_ASAP7_75t_R g1415 ( 
.A(n_1375),
.Y(n_1415)
);

AOI22xp33_ASAP7_75t_L g1416 ( 
.A1(n_1351),
.A2(n_1235),
.B1(n_1301),
.B2(n_1270),
.Y(n_1416)
);

OR2x2_ASAP7_75t_L g1417 ( 
.A(n_1239),
.B(n_1249),
.Y(n_1417)
);

INVx2_ASAP7_75t_L g1418 ( 
.A(n_1309),
.Y(n_1418)
);

NAND2xp5_ASAP7_75t_L g1419 ( 
.A(n_1268),
.B(n_1236),
.Y(n_1419)
);

CKINVDCx6p67_ASAP7_75t_R g1420 ( 
.A(n_1321),
.Y(n_1420)
);

AOI21x1_ASAP7_75t_L g1421 ( 
.A1(n_1280),
.A2(n_1292),
.B(n_1294),
.Y(n_1421)
);

INVx2_ASAP7_75t_L g1422 ( 
.A(n_1314),
.Y(n_1422)
);

INVx1_ASAP7_75t_L g1423 ( 
.A(n_1281),
.Y(n_1423)
);

OA21x2_ASAP7_75t_L g1424 ( 
.A1(n_1279),
.A2(n_1316),
.B(n_1372),
.Y(n_1424)
);

INVx2_ASAP7_75t_L g1425 ( 
.A(n_1320),
.Y(n_1425)
);

AOI222xp33_ASAP7_75t_SL g1426 ( 
.A1(n_1252),
.A2(n_1286),
.B1(n_1296),
.B2(n_1304),
.C1(n_1339),
.C2(n_1358),
.Y(n_1426)
);

AOI22xp33_ASAP7_75t_L g1427 ( 
.A1(n_1301),
.A2(n_1373),
.B1(n_1342),
.B2(n_1255),
.Y(n_1427)
);

OAI21x1_ASAP7_75t_L g1428 ( 
.A1(n_1333),
.A2(n_1368),
.B(n_1367),
.Y(n_1428)
);

OA21x2_ASAP7_75t_L g1429 ( 
.A1(n_1310),
.A2(n_1290),
.B(n_1336),
.Y(n_1429)
);

OA21x2_ASAP7_75t_L g1430 ( 
.A1(n_1310),
.A2(n_1332),
.B(n_1365),
.Y(n_1430)
);

INVx2_ASAP7_75t_L g1431 ( 
.A(n_1297),
.Y(n_1431)
);

INVx1_ASAP7_75t_L g1432 ( 
.A(n_1340),
.Y(n_1432)
);

INVx3_ASAP7_75t_L g1433 ( 
.A(n_1361),
.Y(n_1433)
);

AO22x2_ASAP7_75t_L g1434 ( 
.A1(n_1274),
.A2(n_1285),
.B1(n_1373),
.B2(n_1291),
.Y(n_1434)
);

INVx1_ASAP7_75t_L g1435 ( 
.A(n_1331),
.Y(n_1435)
);

OAI21x1_ASAP7_75t_L g1436 ( 
.A1(n_1368),
.A2(n_1284),
.B(n_1364),
.Y(n_1436)
);

AND2x4_ASAP7_75t_L g1437 ( 
.A(n_1257),
.B(n_1237),
.Y(n_1437)
);

O2A1O1Ixp33_ASAP7_75t_L g1438 ( 
.A1(n_1326),
.A2(n_1322),
.B(n_1265),
.C(n_1272),
.Y(n_1438)
);

OAI22xp5_ASAP7_75t_L g1439 ( 
.A1(n_1274),
.A2(n_1307),
.B1(n_1285),
.B2(n_1229),
.Y(n_1439)
);

INVx1_ASAP7_75t_L g1440 ( 
.A(n_1319),
.Y(n_1440)
);

OAI21xp5_ASAP7_75t_L g1441 ( 
.A1(n_1353),
.A2(n_1347),
.B(n_1349),
.Y(n_1441)
);

INVx1_ASAP7_75t_L g1442 ( 
.A(n_1329),
.Y(n_1442)
);

AND2x2_ASAP7_75t_L g1443 ( 
.A(n_1317),
.B(n_1346),
.Y(n_1443)
);

INVx2_ASAP7_75t_L g1444 ( 
.A(n_1297),
.Y(n_1444)
);

AOI21xp5_ASAP7_75t_L g1445 ( 
.A1(n_1303),
.A2(n_1308),
.B(n_1311),
.Y(n_1445)
);

AND2x4_ASAP7_75t_L g1446 ( 
.A(n_1237),
.B(n_1346),
.Y(n_1446)
);

INVx1_ASAP7_75t_L g1447 ( 
.A(n_1370),
.Y(n_1447)
);

INVx2_ASAP7_75t_SL g1448 ( 
.A(n_1354),
.Y(n_1448)
);

OAI21xp5_ASAP7_75t_L g1449 ( 
.A1(n_1348),
.A2(n_1312),
.B(n_1328),
.Y(n_1449)
);

INVx3_ASAP7_75t_L g1450 ( 
.A(n_1361),
.Y(n_1450)
);

NAND2xp33_ASAP7_75t_R g1451 ( 
.A(n_1269),
.B(n_1334),
.Y(n_1451)
);

OAI21x1_ASAP7_75t_L g1452 ( 
.A1(n_1343),
.A2(n_1232),
.B(n_1352),
.Y(n_1452)
);

OAI21x1_ASAP7_75t_L g1453 ( 
.A1(n_1312),
.A2(n_1297),
.B(n_1302),
.Y(n_1453)
);

NOR2xp33_ASAP7_75t_L g1454 ( 
.A(n_1354),
.B(n_1379),
.Y(n_1454)
);

OAI21x1_ASAP7_75t_L g1455 ( 
.A1(n_1267),
.A2(n_1251),
.B(n_1311),
.Y(n_1455)
);

NOR2x1_ASAP7_75t_SL g1456 ( 
.A(n_1374),
.B(n_1335),
.Y(n_1456)
);

OA21x2_ASAP7_75t_L g1457 ( 
.A1(n_1238),
.A2(n_1241),
.B(n_1251),
.Y(n_1457)
);

OAI21x1_ASAP7_75t_L g1458 ( 
.A1(n_1267),
.A2(n_1330),
.B(n_1241),
.Y(n_1458)
);

A2O1A1Ixp33_ASAP7_75t_L g1459 ( 
.A1(n_1341),
.A2(n_1355),
.B(n_1277),
.C(n_1263),
.Y(n_1459)
);

AOI22xp5_ASAP7_75t_L g1460 ( 
.A1(n_1259),
.A2(n_1273),
.B1(n_1261),
.B2(n_1256),
.Y(n_1460)
);

AOI22xp33_ASAP7_75t_L g1461 ( 
.A1(n_1362),
.A2(n_1231),
.B1(n_1374),
.B2(n_1379),
.Y(n_1461)
);

HB1xp67_ASAP7_75t_L g1462 ( 
.A(n_1330),
.Y(n_1462)
);

INVx2_ASAP7_75t_L g1463 ( 
.A(n_1330),
.Y(n_1463)
);

AO31x2_ASAP7_75t_L g1464 ( 
.A1(n_1238),
.A2(n_1267),
.A3(n_1362),
.B(n_1271),
.Y(n_1464)
);

OAI21x1_ASAP7_75t_L g1465 ( 
.A1(n_1362),
.A2(n_1243),
.B(n_1363),
.Y(n_1465)
);

NAND2x1p5_ASAP7_75t_L g1466 ( 
.A(n_1363),
.B(n_1231),
.Y(n_1466)
);

INVx1_ASAP7_75t_L g1467 ( 
.A(n_1362),
.Y(n_1467)
);

INVx4_ASAP7_75t_L g1468 ( 
.A(n_1226),
.Y(n_1468)
);

INVx1_ASAP7_75t_L g1469 ( 
.A(n_1240),
.Y(n_1469)
);

NAND2x1p5_ASAP7_75t_L g1470 ( 
.A(n_1327),
.B(n_1120),
.Y(n_1470)
);

OAI21x1_ASAP7_75t_L g1471 ( 
.A1(n_1227),
.A2(n_1376),
.B(n_1228),
.Y(n_1471)
);

OAI21x1_ASAP7_75t_SL g1472 ( 
.A1(n_1342),
.A2(n_1272),
.B(n_1293),
.Y(n_1472)
);

OR2x2_ASAP7_75t_L g1473 ( 
.A(n_1287),
.B(n_1230),
.Y(n_1473)
);

NOR2xp33_ASAP7_75t_L g1474 ( 
.A(n_1247),
.B(n_908),
.Y(n_1474)
);

NAND2x1p5_ASAP7_75t_L g1475 ( 
.A(n_1327),
.B(n_1120),
.Y(n_1475)
);

AND2x2_ASAP7_75t_L g1476 ( 
.A(n_1305),
.B(n_1289),
.Y(n_1476)
);

OR2x2_ASAP7_75t_L g1477 ( 
.A(n_1287),
.B(n_1230),
.Y(n_1477)
);

AND2x4_ASAP7_75t_L g1478 ( 
.A(n_1288),
.B(n_1371),
.Y(n_1478)
);

AOI21xp5_ASAP7_75t_L g1479 ( 
.A1(n_1247),
.A2(n_1233),
.B(n_1378),
.Y(n_1479)
);

BUFx3_ASAP7_75t_L g1480 ( 
.A(n_1321),
.Y(n_1480)
);

NOR2xp33_ASAP7_75t_L g1481 ( 
.A(n_1247),
.B(n_908),
.Y(n_1481)
);

AND2x2_ASAP7_75t_L g1482 ( 
.A(n_1305),
.B(n_1289),
.Y(n_1482)
);

NAND2x1p5_ASAP7_75t_L g1483 ( 
.A(n_1327),
.B(n_1120),
.Y(n_1483)
);

NAND2xp5_ASAP7_75t_L g1484 ( 
.A(n_1230),
.B(n_1275),
.Y(n_1484)
);

AOI22xp33_ASAP7_75t_L g1485 ( 
.A1(n_1282),
.A2(n_1020),
.B1(n_1360),
.B2(n_759),
.Y(n_1485)
);

BUFx12f_ASAP7_75t_L g1486 ( 
.A(n_1264),
.Y(n_1486)
);

OAI21x1_ASAP7_75t_L g1487 ( 
.A1(n_1227),
.A2(n_1376),
.B(n_1228),
.Y(n_1487)
);

OAI22xp5_ASAP7_75t_L g1488 ( 
.A1(n_1247),
.A2(n_908),
.B1(n_748),
.B2(n_746),
.Y(n_1488)
);

OAI21x1_ASAP7_75t_SL g1489 ( 
.A1(n_1342),
.A2(n_1272),
.B(n_1293),
.Y(n_1489)
);

INVx1_ASAP7_75t_L g1490 ( 
.A(n_1240),
.Y(n_1490)
);

O2A1O1Ixp33_ASAP7_75t_L g1491 ( 
.A1(n_1247),
.A2(n_748),
.B(n_746),
.C(n_908),
.Y(n_1491)
);

A2O1A1Ixp33_ASAP7_75t_L g1492 ( 
.A1(n_1247),
.A2(n_1095),
.B(n_1268),
.C(n_1310),
.Y(n_1492)
);

O2A1O1Ixp33_ASAP7_75t_L g1493 ( 
.A1(n_1247),
.A2(n_748),
.B(n_746),
.C(n_908),
.Y(n_1493)
);

OAI21x1_ASAP7_75t_L g1494 ( 
.A1(n_1227),
.A2(n_1376),
.B(n_1228),
.Y(n_1494)
);

NAND2xp5_ASAP7_75t_L g1495 ( 
.A(n_1230),
.B(n_1275),
.Y(n_1495)
);

INVx1_ASAP7_75t_L g1496 ( 
.A(n_1240),
.Y(n_1496)
);

OAI21xp5_ASAP7_75t_L g1497 ( 
.A1(n_1247),
.A2(n_748),
.B(n_746),
.Y(n_1497)
);

CKINVDCx6p67_ASAP7_75t_R g1498 ( 
.A(n_1321),
.Y(n_1498)
);

OAI21x1_ASAP7_75t_L g1499 ( 
.A1(n_1227),
.A2(n_1376),
.B(n_1228),
.Y(n_1499)
);

AND2x2_ASAP7_75t_L g1500 ( 
.A(n_1305),
.B(n_1289),
.Y(n_1500)
);

NOR2xp33_ASAP7_75t_L g1501 ( 
.A(n_1247),
.B(n_908),
.Y(n_1501)
);

AOI22xp33_ASAP7_75t_SL g1502 ( 
.A1(n_1235),
.A2(n_1020),
.B1(n_1155),
.B2(n_851),
.Y(n_1502)
);

INVx1_ASAP7_75t_L g1503 ( 
.A(n_1240),
.Y(n_1503)
);

INVx1_ASAP7_75t_L g1504 ( 
.A(n_1240),
.Y(n_1504)
);

INVx1_ASAP7_75t_L g1505 ( 
.A(n_1240),
.Y(n_1505)
);

INVx1_ASAP7_75t_L g1506 ( 
.A(n_1240),
.Y(n_1506)
);

BUFx3_ASAP7_75t_L g1507 ( 
.A(n_1321),
.Y(n_1507)
);

AOI22xp33_ASAP7_75t_L g1508 ( 
.A1(n_1282),
.A2(n_1020),
.B1(n_1360),
.B2(n_759),
.Y(n_1508)
);

OAI21x1_ASAP7_75t_L g1509 ( 
.A1(n_1227),
.A2(n_1376),
.B(n_1228),
.Y(n_1509)
);

A2O1A1Ixp33_ASAP7_75t_L g1510 ( 
.A1(n_1247),
.A2(n_1095),
.B(n_1268),
.C(n_1310),
.Y(n_1510)
);

BUFx3_ASAP7_75t_L g1511 ( 
.A(n_1321),
.Y(n_1511)
);

INVx2_ASAP7_75t_L g1512 ( 
.A(n_1315),
.Y(n_1512)
);

INVx2_ASAP7_75t_L g1513 ( 
.A(n_1315),
.Y(n_1513)
);

NAND2xp5_ASAP7_75t_L g1514 ( 
.A(n_1230),
.B(n_1275),
.Y(n_1514)
);

OR2x2_ASAP7_75t_L g1515 ( 
.A(n_1287),
.B(n_1230),
.Y(n_1515)
);

AOI21xp5_ASAP7_75t_L g1516 ( 
.A1(n_1247),
.A2(n_1233),
.B(n_1378),
.Y(n_1516)
);

INVx1_ASAP7_75t_SL g1517 ( 
.A(n_1287),
.Y(n_1517)
);

AOI221xp5_ASAP7_75t_L g1518 ( 
.A1(n_1268),
.A2(n_746),
.B1(n_748),
.B2(n_785),
.C(n_591),
.Y(n_1518)
);

OAI21x1_ASAP7_75t_L g1519 ( 
.A1(n_1227),
.A2(n_1376),
.B(n_1228),
.Y(n_1519)
);

NOR2xp33_ASAP7_75t_L g1520 ( 
.A(n_1247),
.B(n_908),
.Y(n_1520)
);

OAI21xp5_ASAP7_75t_L g1521 ( 
.A1(n_1247),
.A2(n_748),
.B(n_746),
.Y(n_1521)
);

INVx2_ASAP7_75t_L g1522 ( 
.A(n_1315),
.Y(n_1522)
);

AO31x2_ASAP7_75t_L g1523 ( 
.A1(n_1247),
.A2(n_1372),
.A3(n_1342),
.B(n_1283),
.Y(n_1523)
);

AO21x1_ASAP7_75t_L g1524 ( 
.A1(n_1268),
.A2(n_1095),
.B(n_908),
.Y(n_1524)
);

INVx2_ASAP7_75t_L g1525 ( 
.A(n_1315),
.Y(n_1525)
);

OAI21x1_ASAP7_75t_L g1526 ( 
.A1(n_1227),
.A2(n_1376),
.B(n_1228),
.Y(n_1526)
);

AND2x2_ASAP7_75t_L g1527 ( 
.A(n_1305),
.B(n_1289),
.Y(n_1527)
);

INVx3_ASAP7_75t_L g1528 ( 
.A(n_1226),
.Y(n_1528)
);

NOR2xp33_ASAP7_75t_L g1529 ( 
.A(n_1247),
.B(n_908),
.Y(n_1529)
);

AO21x2_ASAP7_75t_L g1530 ( 
.A1(n_1247),
.A2(n_1378),
.B(n_1376),
.Y(n_1530)
);

OAI21xp5_ASAP7_75t_L g1531 ( 
.A1(n_1247),
.A2(n_748),
.B(n_746),
.Y(n_1531)
);

CKINVDCx5p33_ASAP7_75t_R g1532 ( 
.A(n_1264),
.Y(n_1532)
);

AOI22xp33_ASAP7_75t_L g1533 ( 
.A1(n_1282),
.A2(n_1020),
.B1(n_1360),
.B2(n_759),
.Y(n_1533)
);

INVx3_ASAP7_75t_L g1534 ( 
.A(n_1226),
.Y(n_1534)
);

OAI21x1_ASAP7_75t_L g1535 ( 
.A1(n_1227),
.A2(n_1376),
.B(n_1228),
.Y(n_1535)
);

AO31x2_ASAP7_75t_L g1536 ( 
.A1(n_1247),
.A2(n_1372),
.A3(n_1342),
.B(n_1283),
.Y(n_1536)
);

INVx3_ASAP7_75t_L g1537 ( 
.A(n_1226),
.Y(n_1537)
);

INVx1_ASAP7_75t_L g1538 ( 
.A(n_1240),
.Y(n_1538)
);

INVx1_ASAP7_75t_L g1539 ( 
.A(n_1240),
.Y(n_1539)
);

CKINVDCx5p33_ASAP7_75t_R g1540 ( 
.A(n_1264),
.Y(n_1540)
);

O2A1O1Ixp33_ASAP7_75t_L g1541 ( 
.A1(n_1247),
.A2(n_748),
.B(n_746),
.C(n_908),
.Y(n_1541)
);

OAI22xp5_ASAP7_75t_L g1542 ( 
.A1(n_1518),
.A2(n_1502),
.B1(n_1416),
.B2(n_1394),
.Y(n_1542)
);

O2A1O1Ixp5_ASAP7_75t_L g1543 ( 
.A1(n_1497),
.A2(n_1531),
.B(n_1521),
.C(n_1488),
.Y(n_1543)
);

AOI21xp5_ASAP7_75t_SL g1544 ( 
.A1(n_1491),
.A2(n_1541),
.B(n_1493),
.Y(n_1544)
);

INVx2_ASAP7_75t_L g1545 ( 
.A(n_1383),
.Y(n_1545)
);

CKINVDCx20_ASAP7_75t_R g1546 ( 
.A(n_1415),
.Y(n_1546)
);

HB1xp67_ASAP7_75t_L g1547 ( 
.A(n_1462),
.Y(n_1547)
);

OA21x2_ASAP7_75t_L g1548 ( 
.A1(n_1455),
.A2(n_1458),
.B(n_1393),
.Y(n_1548)
);

AND2x2_ASAP7_75t_L g1549 ( 
.A(n_1387),
.B(n_1476),
.Y(n_1549)
);

OAI22xp5_ASAP7_75t_L g1550 ( 
.A1(n_1416),
.A2(n_1394),
.B1(n_1533),
.B2(n_1485),
.Y(n_1550)
);

NAND2xp5_ASAP7_75t_L g1551 ( 
.A(n_1484),
.B(n_1495),
.Y(n_1551)
);

OAI22xp5_ASAP7_75t_L g1552 ( 
.A1(n_1485),
.A2(n_1508),
.B1(n_1533),
.B2(n_1406),
.Y(n_1552)
);

AND2x4_ASAP7_75t_SL g1553 ( 
.A(n_1420),
.B(n_1498),
.Y(n_1553)
);

OAI22xp5_ASAP7_75t_L g1554 ( 
.A1(n_1508),
.A2(n_1406),
.B1(n_1501),
.B2(n_1520),
.Y(n_1554)
);

AND2x2_ASAP7_75t_L g1555 ( 
.A(n_1482),
.B(n_1500),
.Y(n_1555)
);

NAND2xp5_ASAP7_75t_L g1556 ( 
.A(n_1514),
.B(n_1404),
.Y(n_1556)
);

AOI21xp5_ASAP7_75t_SL g1557 ( 
.A1(n_1474),
.A2(n_1501),
.B(n_1481),
.Y(n_1557)
);

INVx1_ASAP7_75t_L g1558 ( 
.A(n_1386),
.Y(n_1558)
);

OR2x2_ASAP7_75t_L g1559 ( 
.A(n_1401),
.B(n_1473),
.Y(n_1559)
);

AOI221xp5_ASAP7_75t_L g1560 ( 
.A1(n_1474),
.A2(n_1529),
.B1(n_1520),
.B2(n_1481),
.C(n_1510),
.Y(n_1560)
);

AND2x4_ASAP7_75t_L g1561 ( 
.A(n_1384),
.B(n_1478),
.Y(n_1561)
);

OAI22xp5_ASAP7_75t_L g1562 ( 
.A1(n_1529),
.A2(n_1419),
.B1(n_1398),
.B2(n_1492),
.Y(n_1562)
);

BUFx2_ASAP7_75t_L g1563 ( 
.A(n_1396),
.Y(n_1563)
);

OAI22xp5_ASAP7_75t_L g1564 ( 
.A1(n_1398),
.A2(n_1492),
.B1(n_1510),
.B2(n_1460),
.Y(n_1564)
);

AOI21xp5_ASAP7_75t_L g1565 ( 
.A1(n_1530),
.A2(n_1385),
.B(n_1408),
.Y(n_1565)
);

OAI22xp5_ASAP7_75t_L g1566 ( 
.A1(n_1461),
.A2(n_1440),
.B1(n_1442),
.B2(n_1459),
.Y(n_1566)
);

OAI22xp5_ASAP7_75t_SL g1567 ( 
.A1(n_1486),
.A2(n_1540),
.B1(n_1403),
.B2(n_1532),
.Y(n_1567)
);

O2A1O1Ixp5_ASAP7_75t_L g1568 ( 
.A1(n_1524),
.A2(n_1441),
.B(n_1421),
.C(n_1449),
.Y(n_1568)
);

BUFx2_ASAP7_75t_L g1569 ( 
.A(n_1437),
.Y(n_1569)
);

OA21x2_ASAP7_75t_L g1570 ( 
.A1(n_1392),
.A2(n_1390),
.B(n_1389),
.Y(n_1570)
);

OR2x2_ASAP7_75t_L g1571 ( 
.A(n_1477),
.B(n_1515),
.Y(n_1571)
);

O2A1O1Ixp5_ASAP7_75t_L g1572 ( 
.A1(n_1445),
.A2(n_1463),
.B(n_1459),
.C(n_1439),
.Y(n_1572)
);

AND2x2_ASAP7_75t_L g1573 ( 
.A(n_1527),
.B(n_1391),
.Y(n_1573)
);

A2O1A1Ixp33_ASAP7_75t_L g1574 ( 
.A1(n_1438),
.A2(n_1436),
.B(n_1408),
.C(n_1427),
.Y(n_1574)
);

INVx1_ASAP7_75t_L g1575 ( 
.A(n_1409),
.Y(n_1575)
);

OAI22xp5_ASAP7_75t_L g1576 ( 
.A1(n_1461),
.A2(n_1467),
.B1(n_1427),
.B2(n_1414),
.Y(n_1576)
);

HB1xp67_ASAP7_75t_L g1577 ( 
.A(n_1464),
.Y(n_1577)
);

INVx1_ASAP7_75t_L g1578 ( 
.A(n_1411),
.Y(n_1578)
);

OR2x2_ASAP7_75t_L g1579 ( 
.A(n_1517),
.B(n_1417),
.Y(n_1579)
);

INVx1_ASAP7_75t_L g1580 ( 
.A(n_1413),
.Y(n_1580)
);

NAND2xp5_ASAP7_75t_L g1581 ( 
.A(n_1384),
.B(n_1478),
.Y(n_1581)
);

NAND2xp5_ASAP7_75t_L g1582 ( 
.A(n_1384),
.B(n_1478),
.Y(n_1582)
);

AND2x2_ASAP7_75t_L g1583 ( 
.A(n_1443),
.B(n_1437),
.Y(n_1583)
);

AOI221xp5_ASAP7_75t_L g1584 ( 
.A1(n_1434),
.A2(n_1489),
.B1(n_1472),
.B2(n_1538),
.C(n_1496),
.Y(n_1584)
);

OAI22xp5_ASAP7_75t_L g1585 ( 
.A1(n_1434),
.A2(n_1466),
.B1(n_1507),
.B2(n_1511),
.Y(n_1585)
);

HB1xp67_ASAP7_75t_L g1586 ( 
.A(n_1464),
.Y(n_1586)
);

BUFx3_ASAP7_75t_L g1587 ( 
.A(n_1480),
.Y(n_1587)
);

OR2x2_ASAP7_75t_L g1588 ( 
.A(n_1423),
.B(n_1469),
.Y(n_1588)
);

AND2x2_ASAP7_75t_SL g1589 ( 
.A(n_1424),
.B(n_1446),
.Y(n_1589)
);

OAI22xp5_ASAP7_75t_L g1590 ( 
.A1(n_1434),
.A2(n_1466),
.B1(n_1507),
.B2(n_1480),
.Y(n_1590)
);

HB1xp67_ASAP7_75t_L g1591 ( 
.A(n_1464),
.Y(n_1591)
);

AOI221x1_ASAP7_75t_SL g1592 ( 
.A1(n_1490),
.A2(n_1503),
.B1(n_1539),
.B2(n_1504),
.C(n_1505),
.Y(n_1592)
);

O2A1O1Ixp5_ASAP7_75t_L g1593 ( 
.A1(n_1431),
.A2(n_1444),
.B(n_1425),
.C(n_1422),
.Y(n_1593)
);

AND2x2_ASAP7_75t_L g1594 ( 
.A(n_1402),
.B(n_1383),
.Y(n_1594)
);

NAND2x1p5_ASAP7_75t_L g1595 ( 
.A(n_1465),
.B(n_1452),
.Y(n_1595)
);

AOI211xp5_ASAP7_75t_L g1596 ( 
.A1(n_1506),
.A2(n_1432),
.B(n_1511),
.C(n_1454),
.Y(n_1596)
);

AND2x2_ASAP7_75t_L g1597 ( 
.A(n_1395),
.B(n_1418),
.Y(n_1597)
);

NAND2xp5_ASAP7_75t_L g1598 ( 
.A(n_1435),
.B(n_1412),
.Y(n_1598)
);

OR2x2_ASAP7_75t_L g1599 ( 
.A(n_1422),
.B(n_1425),
.Y(n_1599)
);

INVx1_ASAP7_75t_SL g1600 ( 
.A(n_1403),
.Y(n_1600)
);

AND2x2_ASAP7_75t_SL g1601 ( 
.A(n_1430),
.B(n_1381),
.Y(n_1601)
);

BUFx10_ASAP7_75t_L g1602 ( 
.A(n_1532),
.Y(n_1602)
);

AND2x2_ASAP7_75t_L g1603 ( 
.A(n_1397),
.B(n_1525),
.Y(n_1603)
);

INVx1_ASAP7_75t_L g1604 ( 
.A(n_1397),
.Y(n_1604)
);

BUFx3_ASAP7_75t_L g1605 ( 
.A(n_1486),
.Y(n_1605)
);

AND2x2_ASAP7_75t_L g1606 ( 
.A(n_1418),
.B(n_1525),
.Y(n_1606)
);

OAI22xp5_ASAP7_75t_L g1607 ( 
.A1(n_1433),
.A2(n_1450),
.B1(n_1540),
.B2(n_1483),
.Y(n_1607)
);

INVx1_ASAP7_75t_L g1608 ( 
.A(n_1512),
.Y(n_1608)
);

AND2x2_ASAP7_75t_L g1609 ( 
.A(n_1513),
.B(n_1522),
.Y(n_1609)
);

AND2x2_ASAP7_75t_L g1610 ( 
.A(n_1513),
.B(n_1522),
.Y(n_1610)
);

A2O1A1Ixp33_ASAP7_75t_L g1611 ( 
.A1(n_1465),
.A2(n_1453),
.B(n_1450),
.C(n_1433),
.Y(n_1611)
);

CKINVDCx5p33_ASAP7_75t_R g1612 ( 
.A(n_1415),
.Y(n_1612)
);

NAND2x1p5_ASAP7_75t_L g1613 ( 
.A(n_1468),
.B(n_1537),
.Y(n_1613)
);

INVx2_ASAP7_75t_L g1614 ( 
.A(n_1447),
.Y(n_1614)
);

INVxp33_ASAP7_75t_L g1615 ( 
.A(n_1400),
.Y(n_1615)
);

AND2x4_ASAP7_75t_L g1616 ( 
.A(n_1528),
.B(n_1537),
.Y(n_1616)
);

BUFx2_ASAP7_75t_L g1617 ( 
.A(n_1388),
.Y(n_1617)
);

INVx2_ASAP7_75t_L g1618 ( 
.A(n_1382),
.Y(n_1618)
);

A2O1A1Ixp33_ASAP7_75t_L g1619 ( 
.A1(n_1405),
.A2(n_1428),
.B(n_1534),
.C(n_1448),
.Y(n_1619)
);

INVx3_ASAP7_75t_L g1620 ( 
.A(n_1380),
.Y(n_1620)
);

O2A1O1Ixp5_ASAP7_75t_L g1621 ( 
.A1(n_1444),
.A2(n_1536),
.B(n_1523),
.C(n_1430),
.Y(n_1621)
);

OR2x6_ASAP7_75t_L g1622 ( 
.A(n_1429),
.B(n_1430),
.Y(n_1622)
);

OA21x2_ASAP7_75t_L g1623 ( 
.A1(n_1471),
.A2(n_1509),
.B(n_1535),
.Y(n_1623)
);

O2A1O1Ixp5_ASAP7_75t_L g1624 ( 
.A1(n_1536),
.A2(n_1523),
.B(n_1426),
.C(n_1456),
.Y(n_1624)
);

AOI21x1_ASAP7_75t_SL g1625 ( 
.A1(n_1523),
.A2(n_1536),
.B(n_1429),
.Y(n_1625)
);

NAND2xp5_ASAP7_75t_L g1626 ( 
.A(n_1523),
.B(n_1536),
.Y(n_1626)
);

HB1xp67_ASAP7_75t_L g1627 ( 
.A(n_1457),
.Y(n_1627)
);

NAND2xp5_ASAP7_75t_L g1628 ( 
.A(n_1382),
.B(n_1399),
.Y(n_1628)
);

OA21x2_ASAP7_75t_L g1629 ( 
.A1(n_1471),
.A2(n_1526),
.B(n_1519),
.Y(n_1629)
);

NAND2xp5_ASAP7_75t_L g1630 ( 
.A(n_1399),
.B(n_1407),
.Y(n_1630)
);

OA21x2_ASAP7_75t_L g1631 ( 
.A1(n_1487),
.A2(n_1499),
.B(n_1494),
.Y(n_1631)
);

INVx2_ASAP7_75t_L g1632 ( 
.A(n_1470),
.Y(n_1632)
);

CKINVDCx5p33_ASAP7_75t_R g1633 ( 
.A(n_1451),
.Y(n_1633)
);

AND2x2_ASAP7_75t_L g1634 ( 
.A(n_1407),
.B(n_1410),
.Y(n_1634)
);

INVx2_ASAP7_75t_L g1635 ( 
.A(n_1475),
.Y(n_1635)
);

OAI22xp5_ASAP7_75t_L g1636 ( 
.A1(n_1475),
.A2(n_1483),
.B1(n_1410),
.B2(n_1407),
.Y(n_1636)
);

AND2x2_ASAP7_75t_L g1637 ( 
.A(n_1410),
.B(n_1457),
.Y(n_1637)
);

INVx1_ASAP7_75t_SL g1638 ( 
.A(n_1451),
.Y(n_1638)
);

INVxp67_ASAP7_75t_L g1639 ( 
.A(n_1426),
.Y(n_1639)
);

O2A1O1Ixp33_ASAP7_75t_L g1640 ( 
.A1(n_1488),
.A2(n_1521),
.B(n_1531),
.C(n_1497),
.Y(n_1640)
);

A2O1A1Ixp33_ASAP7_75t_L g1641 ( 
.A1(n_1518),
.A2(n_1493),
.B(n_1541),
.C(n_1491),
.Y(n_1641)
);

AND2x2_ASAP7_75t_L g1642 ( 
.A(n_1387),
.B(n_1476),
.Y(n_1642)
);

HB1xp67_ASAP7_75t_L g1643 ( 
.A(n_1462),
.Y(n_1643)
);

INVx1_ASAP7_75t_L g1644 ( 
.A(n_1386),
.Y(n_1644)
);

AND2x2_ASAP7_75t_L g1645 ( 
.A(n_1387),
.B(n_1476),
.Y(n_1645)
);

OAI22xp5_ASAP7_75t_L g1646 ( 
.A1(n_1518),
.A2(n_1502),
.B1(n_1416),
.B2(n_1394),
.Y(n_1646)
);

OAI22xp5_ASAP7_75t_L g1647 ( 
.A1(n_1518),
.A2(n_1502),
.B1(n_1416),
.B2(n_1394),
.Y(n_1647)
);

O2A1O1Ixp33_ASAP7_75t_L g1648 ( 
.A1(n_1488),
.A2(n_1521),
.B(n_1531),
.C(n_1497),
.Y(n_1648)
);

INVx1_ASAP7_75t_L g1649 ( 
.A(n_1386),
.Y(n_1649)
);

AND2x4_ASAP7_75t_L g1650 ( 
.A(n_1384),
.B(n_1478),
.Y(n_1650)
);

AND2x4_ASAP7_75t_L g1651 ( 
.A(n_1384),
.B(n_1478),
.Y(n_1651)
);

AND2x2_ASAP7_75t_L g1652 ( 
.A(n_1387),
.B(n_1476),
.Y(n_1652)
);

OAI22x1_ASAP7_75t_L g1653 ( 
.A1(n_1460),
.A2(n_1398),
.B1(n_1481),
.B2(n_1474),
.Y(n_1653)
);

AND2x2_ASAP7_75t_L g1654 ( 
.A(n_1387),
.B(n_1476),
.Y(n_1654)
);

INVx1_ASAP7_75t_L g1655 ( 
.A(n_1386),
.Y(n_1655)
);

OR2x2_ASAP7_75t_L g1656 ( 
.A(n_1401),
.B(n_1473),
.Y(n_1656)
);

BUFx4f_ASAP7_75t_SL g1657 ( 
.A(n_1486),
.Y(n_1657)
);

NOR2xp67_ASAP7_75t_R g1658 ( 
.A(n_1486),
.B(n_1467),
.Y(n_1658)
);

BUFx6f_ASAP7_75t_L g1659 ( 
.A(n_1480),
.Y(n_1659)
);

O2A1O1Ixp33_ASAP7_75t_L g1660 ( 
.A1(n_1488),
.A2(n_1521),
.B(n_1531),
.C(n_1497),
.Y(n_1660)
);

NOR2xp67_ASAP7_75t_L g1661 ( 
.A(n_1433),
.B(n_1229),
.Y(n_1661)
);

AOI21xp5_ASAP7_75t_L g1662 ( 
.A1(n_1479),
.A2(n_1516),
.B(n_1247),
.Y(n_1662)
);

O2A1O1Ixp5_ASAP7_75t_L g1663 ( 
.A1(n_1497),
.A2(n_1521),
.B(n_1531),
.C(n_1488),
.Y(n_1663)
);

O2A1O1Ixp33_ASAP7_75t_L g1664 ( 
.A1(n_1488),
.A2(n_1521),
.B(n_1531),
.C(n_1497),
.Y(n_1664)
);

CKINVDCx5p33_ASAP7_75t_R g1665 ( 
.A(n_1415),
.Y(n_1665)
);

AND2x2_ASAP7_75t_L g1666 ( 
.A(n_1589),
.B(n_1637),
.Y(n_1666)
);

INVx3_ASAP7_75t_L g1667 ( 
.A(n_1595),
.Y(n_1667)
);

INVx3_ASAP7_75t_L g1668 ( 
.A(n_1595),
.Y(n_1668)
);

INVx2_ASAP7_75t_L g1669 ( 
.A(n_1593),
.Y(n_1669)
);

NAND2xp5_ASAP7_75t_L g1670 ( 
.A(n_1559),
.B(n_1571),
.Y(n_1670)
);

NAND2xp5_ASAP7_75t_L g1671 ( 
.A(n_1656),
.B(n_1551),
.Y(n_1671)
);

OR2x2_ASAP7_75t_L g1672 ( 
.A(n_1626),
.B(n_1547),
.Y(n_1672)
);

AND2x2_ASAP7_75t_L g1673 ( 
.A(n_1601),
.B(n_1558),
.Y(n_1673)
);

INVx3_ASAP7_75t_L g1674 ( 
.A(n_1548),
.Y(n_1674)
);

AND2x4_ASAP7_75t_L g1675 ( 
.A(n_1619),
.B(n_1622),
.Y(n_1675)
);

INVx2_ASAP7_75t_SL g1676 ( 
.A(n_1588),
.Y(n_1676)
);

INVx3_ASAP7_75t_L g1677 ( 
.A(n_1548),
.Y(n_1677)
);

OR2x2_ASAP7_75t_L g1678 ( 
.A(n_1547),
.B(n_1643),
.Y(n_1678)
);

AOI22xp5_ASAP7_75t_L g1679 ( 
.A1(n_1542),
.A2(n_1647),
.B1(n_1646),
.B2(n_1550),
.Y(n_1679)
);

OR2x6_ASAP7_75t_L g1680 ( 
.A(n_1662),
.B(n_1565),
.Y(n_1680)
);

AND2x2_ASAP7_75t_L g1681 ( 
.A(n_1575),
.B(n_1578),
.Y(n_1681)
);

NAND2xp5_ASAP7_75t_L g1682 ( 
.A(n_1556),
.B(n_1560),
.Y(n_1682)
);

AND2x2_ASAP7_75t_L g1683 ( 
.A(n_1580),
.B(n_1644),
.Y(n_1683)
);

INVx2_ASAP7_75t_L g1684 ( 
.A(n_1622),
.Y(n_1684)
);

AOI22xp33_ASAP7_75t_L g1685 ( 
.A1(n_1554),
.A2(n_1552),
.B1(n_1560),
.B2(n_1562),
.Y(n_1685)
);

NOR2xp33_ASAP7_75t_L g1686 ( 
.A(n_1638),
.B(n_1633),
.Y(n_1686)
);

AND2x2_ASAP7_75t_L g1687 ( 
.A(n_1649),
.B(n_1655),
.Y(n_1687)
);

NAND2xp5_ASAP7_75t_L g1688 ( 
.A(n_1579),
.B(n_1557),
.Y(n_1688)
);

AND2x2_ASAP7_75t_L g1689 ( 
.A(n_1653),
.B(n_1594),
.Y(n_1689)
);

INVxp33_ASAP7_75t_L g1690 ( 
.A(n_1549),
.Y(n_1690)
);

INVx1_ASAP7_75t_L g1691 ( 
.A(n_1627),
.Y(n_1691)
);

INVx1_ASAP7_75t_L g1692 ( 
.A(n_1627),
.Y(n_1692)
);

INVx1_ASAP7_75t_L g1693 ( 
.A(n_1599),
.Y(n_1693)
);

INVx1_ASAP7_75t_L g1694 ( 
.A(n_1604),
.Y(n_1694)
);

CKINVDCx5p33_ASAP7_75t_R g1695 ( 
.A(n_1612),
.Y(n_1695)
);

INVx2_ASAP7_75t_SL g1696 ( 
.A(n_1614),
.Y(n_1696)
);

OR2x6_ASAP7_75t_L g1697 ( 
.A(n_1662),
.B(n_1565),
.Y(n_1697)
);

INVx1_ASAP7_75t_L g1698 ( 
.A(n_1608),
.Y(n_1698)
);

INVxp67_ASAP7_75t_SL g1699 ( 
.A(n_1598),
.Y(n_1699)
);

INVx4_ASAP7_75t_L g1700 ( 
.A(n_1659),
.Y(n_1700)
);

INVx1_ASAP7_75t_L g1701 ( 
.A(n_1577),
.Y(n_1701)
);

AND2x2_ASAP7_75t_L g1702 ( 
.A(n_1574),
.B(n_1577),
.Y(n_1702)
);

INVx1_ASAP7_75t_L g1703 ( 
.A(n_1586),
.Y(n_1703)
);

AND2x2_ASAP7_75t_L g1704 ( 
.A(n_1586),
.B(n_1591),
.Y(n_1704)
);

BUFx2_ASAP7_75t_L g1705 ( 
.A(n_1591),
.Y(n_1705)
);

INVx1_ASAP7_75t_L g1706 ( 
.A(n_1545),
.Y(n_1706)
);

AND2x2_ASAP7_75t_L g1707 ( 
.A(n_1564),
.B(n_1597),
.Y(n_1707)
);

AND2x2_ASAP7_75t_L g1708 ( 
.A(n_1603),
.B(n_1606),
.Y(n_1708)
);

OAI211xp5_ASAP7_75t_L g1709 ( 
.A1(n_1544),
.A2(n_1639),
.B(n_1641),
.C(n_1640),
.Y(n_1709)
);

INVx1_ASAP7_75t_L g1710 ( 
.A(n_1621),
.Y(n_1710)
);

HB1xp67_ASAP7_75t_L g1711 ( 
.A(n_1592),
.Y(n_1711)
);

INVx2_ASAP7_75t_SL g1712 ( 
.A(n_1659),
.Y(n_1712)
);

INVx2_ASAP7_75t_L g1713 ( 
.A(n_1621),
.Y(n_1713)
);

INVx2_ASAP7_75t_SL g1714 ( 
.A(n_1659),
.Y(n_1714)
);

BUFx3_ASAP7_75t_L g1715 ( 
.A(n_1613),
.Y(n_1715)
);

AO21x2_ASAP7_75t_L g1716 ( 
.A1(n_1640),
.A2(n_1664),
.B(n_1648),
.Y(n_1716)
);

AO21x2_ASAP7_75t_L g1717 ( 
.A1(n_1648),
.A2(n_1664),
.B(n_1660),
.Y(n_1717)
);

BUFx2_ASAP7_75t_L g1718 ( 
.A(n_1611),
.Y(n_1718)
);

INVx2_ASAP7_75t_L g1719 ( 
.A(n_1570),
.Y(n_1719)
);

NAND2xp5_ASAP7_75t_L g1720 ( 
.A(n_1609),
.B(n_1610),
.Y(n_1720)
);

INVxp67_ASAP7_75t_L g1721 ( 
.A(n_1555),
.Y(n_1721)
);

NAND2xp5_ASAP7_75t_L g1722 ( 
.A(n_1639),
.B(n_1581),
.Y(n_1722)
);

INVx1_ASAP7_75t_L g1723 ( 
.A(n_1572),
.Y(n_1723)
);

AO21x2_ASAP7_75t_L g1724 ( 
.A1(n_1660),
.A2(n_1576),
.B(n_1566),
.Y(n_1724)
);

AND2x4_ASAP7_75t_L g1725 ( 
.A(n_1561),
.B(n_1650),
.Y(n_1725)
);

INVx1_ASAP7_75t_L g1726 ( 
.A(n_1572),
.Y(n_1726)
);

INVx1_ASAP7_75t_L g1727 ( 
.A(n_1624),
.Y(n_1727)
);

INVx1_ASAP7_75t_L g1728 ( 
.A(n_1624),
.Y(n_1728)
);

AND2x2_ASAP7_75t_L g1729 ( 
.A(n_1584),
.B(n_1652),
.Y(n_1729)
);

INVx1_ASAP7_75t_L g1730 ( 
.A(n_1568),
.Y(n_1730)
);

INVx1_ASAP7_75t_L g1731 ( 
.A(n_1568),
.Y(n_1731)
);

OR2x2_ASAP7_75t_L g1732 ( 
.A(n_1585),
.B(n_1590),
.Y(n_1732)
);

INVx1_ASAP7_75t_L g1733 ( 
.A(n_1584),
.Y(n_1733)
);

OA21x2_ASAP7_75t_L g1734 ( 
.A1(n_1543),
.A2(n_1663),
.B(n_1625),
.Y(n_1734)
);

NAND2xp5_ASAP7_75t_L g1735 ( 
.A(n_1582),
.B(n_1573),
.Y(n_1735)
);

OA21x2_ASAP7_75t_L g1736 ( 
.A1(n_1543),
.A2(n_1663),
.B(n_1628),
.Y(n_1736)
);

OR2x2_ASAP7_75t_L g1737 ( 
.A(n_1563),
.B(n_1569),
.Y(n_1737)
);

BUFx2_ASAP7_75t_SL g1738 ( 
.A(n_1587),
.Y(n_1738)
);

NAND3xp33_ASAP7_75t_L g1739 ( 
.A(n_1709),
.B(n_1596),
.C(n_1607),
.Y(n_1739)
);

INVx2_ASAP7_75t_L g1740 ( 
.A(n_1719),
.Y(n_1740)
);

AND2x2_ASAP7_75t_L g1741 ( 
.A(n_1680),
.B(n_1631),
.Y(n_1741)
);

OAI22xp33_ASAP7_75t_L g1742 ( 
.A1(n_1679),
.A2(n_1657),
.B1(n_1615),
.B2(n_1605),
.Y(n_1742)
);

OR2x2_ASAP7_75t_L g1743 ( 
.A(n_1710),
.B(n_1623),
.Y(n_1743)
);

OR2x2_ASAP7_75t_L g1744 ( 
.A(n_1710),
.B(n_1629),
.Y(n_1744)
);

AND2x2_ASAP7_75t_L g1745 ( 
.A(n_1680),
.B(n_1631),
.Y(n_1745)
);

INVx1_ASAP7_75t_L g1746 ( 
.A(n_1691),
.Y(n_1746)
);

NAND2xp5_ASAP7_75t_SL g1747 ( 
.A(n_1679),
.B(n_1651),
.Y(n_1747)
);

NAND2xp5_ASAP7_75t_L g1748 ( 
.A(n_1699),
.B(n_1645),
.Y(n_1748)
);

OAI22xp5_ASAP7_75t_L g1749 ( 
.A1(n_1685),
.A2(n_1657),
.B1(n_1654),
.B2(n_1642),
.Y(n_1749)
);

HB1xp67_ASAP7_75t_L g1750 ( 
.A(n_1691),
.Y(n_1750)
);

AND2x2_ASAP7_75t_L g1751 ( 
.A(n_1680),
.B(n_1650),
.Y(n_1751)
);

OR2x2_ASAP7_75t_L g1752 ( 
.A(n_1672),
.B(n_1618),
.Y(n_1752)
);

OR2x2_ASAP7_75t_L g1753 ( 
.A(n_1672),
.B(n_1617),
.Y(n_1753)
);

OR2x2_ASAP7_75t_L g1754 ( 
.A(n_1692),
.B(n_1630),
.Y(n_1754)
);

NAND2xp5_ASAP7_75t_L g1755 ( 
.A(n_1716),
.B(n_1632),
.Y(n_1755)
);

AND2x2_ASAP7_75t_L g1756 ( 
.A(n_1697),
.B(n_1583),
.Y(n_1756)
);

INVx1_ASAP7_75t_L g1757 ( 
.A(n_1692),
.Y(n_1757)
);

INVx1_ASAP7_75t_SL g1758 ( 
.A(n_1688),
.Y(n_1758)
);

NAND2xp5_ASAP7_75t_L g1759 ( 
.A(n_1716),
.B(n_1635),
.Y(n_1759)
);

NAND2xp5_ASAP7_75t_L g1760 ( 
.A(n_1716),
.B(n_1658),
.Y(n_1760)
);

AND2x2_ASAP7_75t_L g1761 ( 
.A(n_1673),
.B(n_1634),
.Y(n_1761)
);

INVx1_ASAP7_75t_L g1762 ( 
.A(n_1694),
.Y(n_1762)
);

NAND2xp5_ASAP7_75t_L g1763 ( 
.A(n_1717),
.B(n_1620),
.Y(n_1763)
);

INVxp67_ASAP7_75t_SL g1764 ( 
.A(n_1669),
.Y(n_1764)
);

AND2x4_ASAP7_75t_SL g1765 ( 
.A(n_1675),
.B(n_1616),
.Y(n_1765)
);

AND2x2_ASAP7_75t_L g1766 ( 
.A(n_1684),
.B(n_1702),
.Y(n_1766)
);

OAI221xp5_ASAP7_75t_L g1767 ( 
.A1(n_1733),
.A2(n_1661),
.B1(n_1600),
.B2(n_1567),
.C(n_1636),
.Y(n_1767)
);

INVxp67_ASAP7_75t_L g1768 ( 
.A(n_1711),
.Y(n_1768)
);

AND2x2_ASAP7_75t_L g1769 ( 
.A(n_1702),
.B(n_1666),
.Y(n_1769)
);

INVx4_ASAP7_75t_SL g1770 ( 
.A(n_1675),
.Y(n_1770)
);

HB1xp67_ASAP7_75t_L g1771 ( 
.A(n_1705),
.Y(n_1771)
);

NAND2xp5_ASAP7_75t_L g1772 ( 
.A(n_1717),
.B(n_1676),
.Y(n_1772)
);

NAND2xp5_ASAP7_75t_L g1773 ( 
.A(n_1758),
.B(n_1670),
.Y(n_1773)
);

OAI22xp33_ASAP7_75t_L g1774 ( 
.A1(n_1739),
.A2(n_1732),
.B1(n_1733),
.B2(n_1718),
.Y(n_1774)
);

NOR4xp25_ASAP7_75t_SL g1775 ( 
.A(n_1767),
.B(n_1718),
.C(n_1731),
.D(n_1730),
.Y(n_1775)
);

AND4x1_ASAP7_75t_L g1776 ( 
.A(n_1739),
.B(n_1686),
.C(n_1760),
.D(n_1731),
.Y(n_1776)
);

OAI221xp5_ASAP7_75t_L g1777 ( 
.A1(n_1768),
.A2(n_1682),
.B1(n_1722),
.B2(n_1732),
.C(n_1671),
.Y(n_1777)
);

AOI22xp33_ASAP7_75t_L g1778 ( 
.A1(n_1768),
.A2(n_1724),
.B1(n_1717),
.B2(n_1727),
.Y(n_1778)
);

OAI211xp5_ASAP7_75t_SL g1779 ( 
.A1(n_1758),
.A2(n_1767),
.B(n_1772),
.C(n_1747),
.Y(n_1779)
);

NAND4xp25_ASAP7_75t_L g1780 ( 
.A(n_1755),
.B(n_1728),
.C(n_1727),
.D(n_1729),
.Y(n_1780)
);

INVx1_ASAP7_75t_L g1781 ( 
.A(n_1746),
.Y(n_1781)
);

AO21x1_ASAP7_75t_SL g1782 ( 
.A1(n_1760),
.A2(n_1728),
.B(n_1723),
.Y(n_1782)
);

AND2x2_ASAP7_75t_L g1783 ( 
.A(n_1769),
.B(n_1666),
.Y(n_1783)
);

AOI221xp5_ASAP7_75t_L g1784 ( 
.A1(n_1749),
.A2(n_1772),
.B1(n_1717),
.B2(n_1742),
.C(n_1729),
.Y(n_1784)
);

NAND3xp33_ASAP7_75t_L g1785 ( 
.A(n_1759),
.B(n_1763),
.C(n_1736),
.Y(n_1785)
);

NAND2xp5_ASAP7_75t_L g1786 ( 
.A(n_1748),
.B(n_1676),
.Y(n_1786)
);

OR2x2_ASAP7_75t_L g1787 ( 
.A(n_1752),
.B(n_1693),
.Y(n_1787)
);

INVx2_ASAP7_75t_L g1788 ( 
.A(n_1740),
.Y(n_1788)
);

AOI22xp33_ASAP7_75t_L g1789 ( 
.A1(n_1749),
.A2(n_1724),
.B1(n_1723),
.B2(n_1726),
.Y(n_1789)
);

OR2x2_ASAP7_75t_L g1790 ( 
.A(n_1752),
.B(n_1693),
.Y(n_1790)
);

NOR3xp33_ASAP7_75t_SL g1791 ( 
.A(n_1742),
.B(n_1665),
.C(n_1695),
.Y(n_1791)
);

AND2x2_ASAP7_75t_SL g1792 ( 
.A(n_1765),
.B(n_1675),
.Y(n_1792)
);

AND2x4_ASAP7_75t_L g1793 ( 
.A(n_1770),
.B(n_1675),
.Y(n_1793)
);

BUFx2_ASAP7_75t_SL g1794 ( 
.A(n_1761),
.Y(n_1794)
);

AND2x2_ASAP7_75t_L g1795 ( 
.A(n_1769),
.B(n_1689),
.Y(n_1795)
);

AOI221xp5_ASAP7_75t_L g1796 ( 
.A1(n_1759),
.A2(n_1726),
.B1(n_1724),
.B2(n_1690),
.C(n_1721),
.Y(n_1796)
);

NAND3xp33_ASAP7_75t_L g1797 ( 
.A(n_1763),
.B(n_1736),
.C(n_1689),
.Y(n_1797)
);

INVx1_ASAP7_75t_L g1798 ( 
.A(n_1746),
.Y(n_1798)
);

OAI22xp5_ASAP7_75t_L g1799 ( 
.A1(n_1748),
.A2(n_1738),
.B1(n_1737),
.B2(n_1707),
.Y(n_1799)
);

OAI31xp33_ASAP7_75t_SL g1800 ( 
.A1(n_1769),
.A2(n_1707),
.A3(n_1725),
.B(n_1724),
.Y(n_1800)
);

INVx4_ASAP7_75t_L g1801 ( 
.A(n_1770),
.Y(n_1801)
);

AOI222xp33_ASAP7_75t_L g1802 ( 
.A1(n_1756),
.A2(n_1735),
.B1(n_1553),
.B2(n_1546),
.C1(n_1683),
.C2(n_1681),
.Y(n_1802)
);

AND2x2_ASAP7_75t_L g1803 ( 
.A(n_1766),
.B(n_1704),
.Y(n_1803)
);

AOI221xp5_ASAP7_75t_L g1804 ( 
.A1(n_1764),
.A2(n_1681),
.B1(n_1683),
.B2(n_1687),
.C(n_1696),
.Y(n_1804)
);

AOI22xp33_ASAP7_75t_L g1805 ( 
.A1(n_1753),
.A2(n_1736),
.B1(n_1734),
.B2(n_1737),
.Y(n_1805)
);

AOI221xp5_ASAP7_75t_L g1806 ( 
.A1(n_1764),
.A2(n_1687),
.B1(n_1696),
.B2(n_1698),
.C(n_1706),
.Y(n_1806)
);

OAI221xp5_ASAP7_75t_L g1807 ( 
.A1(n_1753),
.A2(n_1738),
.B1(n_1712),
.B2(n_1714),
.C(n_1715),
.Y(n_1807)
);

OAI221xp5_ASAP7_75t_L g1808 ( 
.A1(n_1753),
.A2(n_1712),
.B1(n_1714),
.B2(n_1715),
.C(n_1700),
.Y(n_1808)
);

AOI322xp5_ASAP7_75t_L g1809 ( 
.A1(n_1766),
.A2(n_1704),
.A3(n_1713),
.B1(n_1705),
.B2(n_1708),
.C1(n_1703),
.C2(n_1701),
.Y(n_1809)
);

NAND2xp5_ASAP7_75t_L g1810 ( 
.A(n_1754),
.B(n_1708),
.Y(n_1810)
);

AOI22xp33_ASAP7_75t_L g1811 ( 
.A1(n_1756),
.A2(n_1734),
.B1(n_1725),
.B2(n_1602),
.Y(n_1811)
);

BUFx3_ASAP7_75t_L g1812 ( 
.A(n_1754),
.Y(n_1812)
);

NAND2xp5_ASAP7_75t_L g1813 ( 
.A(n_1754),
.B(n_1720),
.Y(n_1813)
);

NAND4xp25_ASAP7_75t_L g1814 ( 
.A(n_1752),
.B(n_1698),
.C(n_1678),
.D(n_1701),
.Y(n_1814)
);

OAI221xp5_ASAP7_75t_L g1815 ( 
.A1(n_1751),
.A2(n_1715),
.B1(n_1700),
.B2(n_1667),
.C(n_1668),
.Y(n_1815)
);

INVx1_ASAP7_75t_L g1816 ( 
.A(n_1757),
.Y(n_1816)
);

HB1xp67_ASAP7_75t_L g1817 ( 
.A(n_1771),
.Y(n_1817)
);

NOR2xp33_ASAP7_75t_R g1818 ( 
.A(n_1762),
.B(n_1602),
.Y(n_1818)
);

BUFx2_ASAP7_75t_L g1819 ( 
.A(n_1801),
.Y(n_1819)
);

INVx1_ASAP7_75t_L g1820 ( 
.A(n_1781),
.Y(n_1820)
);

INVx1_ASAP7_75t_L g1821 ( 
.A(n_1798),
.Y(n_1821)
);

BUFx3_ASAP7_75t_L g1822 ( 
.A(n_1801),
.Y(n_1822)
);

NAND2xp5_ASAP7_75t_L g1823 ( 
.A(n_1800),
.B(n_1750),
.Y(n_1823)
);

INVx1_ASAP7_75t_L g1824 ( 
.A(n_1816),
.Y(n_1824)
);

OAI21xp5_ASAP7_75t_L g1825 ( 
.A1(n_1784),
.A2(n_1734),
.B(n_1741),
.Y(n_1825)
);

BUFx2_ASAP7_75t_L g1826 ( 
.A(n_1801),
.Y(n_1826)
);

OAI21xp5_ASAP7_75t_L g1827 ( 
.A1(n_1776),
.A2(n_1734),
.B(n_1741),
.Y(n_1827)
);

NAND2xp5_ASAP7_75t_L g1828 ( 
.A(n_1796),
.B(n_1750),
.Y(n_1828)
);

INVx2_ASAP7_75t_L g1829 ( 
.A(n_1788),
.Y(n_1829)
);

INVx2_ASAP7_75t_L g1830 ( 
.A(n_1788),
.Y(n_1830)
);

NAND3xp33_ASAP7_75t_L g1831 ( 
.A(n_1778),
.B(n_1713),
.C(n_1744),
.Y(n_1831)
);

OAI21xp5_ASAP7_75t_L g1832 ( 
.A1(n_1778),
.A2(n_1741),
.B(n_1745),
.Y(n_1832)
);

INVxp67_ASAP7_75t_SL g1833 ( 
.A(n_1817),
.Y(n_1833)
);

OAI21x1_ASAP7_75t_L g1834 ( 
.A1(n_1805),
.A2(n_1674),
.B(n_1677),
.Y(n_1834)
);

OR2x2_ASAP7_75t_L g1835 ( 
.A(n_1785),
.B(n_1743),
.Y(n_1835)
);

AND2x2_ASAP7_75t_L g1836 ( 
.A(n_1794),
.B(n_1745),
.Y(n_1836)
);

INVx1_ASAP7_75t_SL g1837 ( 
.A(n_1818),
.Y(n_1837)
);

AND2x2_ASAP7_75t_L g1838 ( 
.A(n_1783),
.B(n_1745),
.Y(n_1838)
);

HB1xp67_ASAP7_75t_L g1839 ( 
.A(n_1812),
.Y(n_1839)
);

CKINVDCx5p33_ASAP7_75t_R g1840 ( 
.A(n_1818),
.Y(n_1840)
);

INVx3_ASAP7_75t_L g1841 ( 
.A(n_1793),
.Y(n_1841)
);

INVxp33_ASAP7_75t_L g1842 ( 
.A(n_1791),
.Y(n_1842)
);

INVx2_ASAP7_75t_L g1843 ( 
.A(n_1812),
.Y(n_1843)
);

AND2x4_ASAP7_75t_L g1844 ( 
.A(n_1793),
.B(n_1770),
.Y(n_1844)
);

NAND3xp33_ASAP7_75t_L g1845 ( 
.A(n_1775),
.B(n_1713),
.C(n_1743),
.Y(n_1845)
);

INVx4_ASAP7_75t_L g1846 ( 
.A(n_1793),
.Y(n_1846)
);

INVx2_ASAP7_75t_SL g1847 ( 
.A(n_1792),
.Y(n_1847)
);

INVx2_ASAP7_75t_L g1848 ( 
.A(n_1803),
.Y(n_1848)
);

HB1xp67_ASAP7_75t_L g1849 ( 
.A(n_1814),
.Y(n_1849)
);

NAND2xp5_ASAP7_75t_L g1850 ( 
.A(n_1797),
.B(n_1757),
.Y(n_1850)
);

NAND2xp67_ASAP7_75t_L g1851 ( 
.A(n_1843),
.B(n_1773),
.Y(n_1851)
);

NAND4xp25_ASAP7_75t_L g1852 ( 
.A(n_1825),
.B(n_1789),
.C(n_1779),
.D(n_1777),
.Y(n_1852)
);

INVx2_ASAP7_75t_L g1853 ( 
.A(n_1829),
.Y(n_1853)
);

INVx2_ASAP7_75t_L g1854 ( 
.A(n_1829),
.Y(n_1854)
);

NOR2xp67_ASAP7_75t_L g1855 ( 
.A(n_1847),
.B(n_1780),
.Y(n_1855)
);

NAND4xp25_ASAP7_75t_SL g1856 ( 
.A(n_1825),
.B(n_1802),
.C(n_1789),
.D(n_1809),
.Y(n_1856)
);

INVx1_ASAP7_75t_L g1857 ( 
.A(n_1820),
.Y(n_1857)
);

INVx2_ASAP7_75t_L g1858 ( 
.A(n_1829),
.Y(n_1858)
);

AND2x2_ASAP7_75t_L g1859 ( 
.A(n_1844),
.B(n_1795),
.Y(n_1859)
);

AND2x4_ASAP7_75t_L g1860 ( 
.A(n_1844),
.B(n_1770),
.Y(n_1860)
);

INVx1_ASAP7_75t_L g1861 ( 
.A(n_1820),
.Y(n_1861)
);

AND2x2_ASAP7_75t_L g1862 ( 
.A(n_1844),
.B(n_1782),
.Y(n_1862)
);

INVx2_ASAP7_75t_L g1863 ( 
.A(n_1829),
.Y(n_1863)
);

NAND2x1p5_ASAP7_75t_L g1864 ( 
.A(n_1822),
.B(n_1792),
.Y(n_1864)
);

INVx1_ASAP7_75t_L g1865 ( 
.A(n_1820),
.Y(n_1865)
);

INVx3_ASAP7_75t_L g1866 ( 
.A(n_1844),
.Y(n_1866)
);

OR2x2_ASAP7_75t_L g1867 ( 
.A(n_1850),
.B(n_1810),
.Y(n_1867)
);

OR2x2_ASAP7_75t_L g1868 ( 
.A(n_1850),
.B(n_1787),
.Y(n_1868)
);

INVx2_ASAP7_75t_L g1869 ( 
.A(n_1829),
.Y(n_1869)
);

NAND2xp5_ASAP7_75t_L g1870 ( 
.A(n_1849),
.B(n_1774),
.Y(n_1870)
);

AND2x2_ASAP7_75t_L g1871 ( 
.A(n_1844),
.B(n_1803),
.Y(n_1871)
);

INVx1_ASAP7_75t_L g1872 ( 
.A(n_1821),
.Y(n_1872)
);

AND2x2_ASAP7_75t_L g1873 ( 
.A(n_1844),
.B(n_1846),
.Y(n_1873)
);

INVx1_ASAP7_75t_L g1874 ( 
.A(n_1821),
.Y(n_1874)
);

OR2x2_ASAP7_75t_L g1875 ( 
.A(n_1850),
.B(n_1790),
.Y(n_1875)
);

NAND3xp33_ASAP7_75t_L g1876 ( 
.A(n_1825),
.B(n_1805),
.C(n_1811),
.Y(n_1876)
);

OAI31xp33_ASAP7_75t_L g1877 ( 
.A1(n_1849),
.A2(n_1842),
.A3(n_1831),
.B(n_1823),
.Y(n_1877)
);

NAND2xp5_ASAP7_75t_L g1878 ( 
.A(n_1843),
.B(n_1804),
.Y(n_1878)
);

NAND2xp5_ASAP7_75t_L g1879 ( 
.A(n_1843),
.B(n_1799),
.Y(n_1879)
);

INVx2_ASAP7_75t_SL g1880 ( 
.A(n_1844),
.Y(n_1880)
);

NAND2xp5_ASAP7_75t_L g1881 ( 
.A(n_1843),
.B(n_1766),
.Y(n_1881)
);

NOR2x1_ASAP7_75t_L g1882 ( 
.A(n_1837),
.B(n_1822),
.Y(n_1882)
);

OR2x2_ASAP7_75t_L g1883 ( 
.A(n_1828),
.B(n_1813),
.Y(n_1883)
);

BUFx3_ASAP7_75t_L g1884 ( 
.A(n_1840),
.Y(n_1884)
);

NOR3xp33_ASAP7_75t_L g1885 ( 
.A(n_1832),
.B(n_1831),
.C(n_1828),
.Y(n_1885)
);

INVxp67_ASAP7_75t_L g1886 ( 
.A(n_1839),
.Y(n_1886)
);

INVx2_ASAP7_75t_L g1887 ( 
.A(n_1830),
.Y(n_1887)
);

AND2x2_ASAP7_75t_L g1888 ( 
.A(n_1846),
.B(n_1770),
.Y(n_1888)
);

AND2x2_ASAP7_75t_L g1889 ( 
.A(n_1846),
.B(n_1847),
.Y(n_1889)
);

INVx1_ASAP7_75t_L g1890 ( 
.A(n_1821),
.Y(n_1890)
);

AOI31xp33_ASAP7_75t_L g1891 ( 
.A1(n_1842),
.A2(n_1811),
.A3(n_1807),
.B(n_1808),
.Y(n_1891)
);

OR2x2_ASAP7_75t_L g1892 ( 
.A(n_1828),
.B(n_1786),
.Y(n_1892)
);

INVx1_ASAP7_75t_L g1893 ( 
.A(n_1824),
.Y(n_1893)
);

NAND3xp33_ASAP7_75t_L g1894 ( 
.A(n_1831),
.B(n_1806),
.C(n_1815),
.Y(n_1894)
);

AND2x2_ASAP7_75t_L g1895 ( 
.A(n_1846),
.B(n_1770),
.Y(n_1895)
);

INVx1_ASAP7_75t_L g1896 ( 
.A(n_1824),
.Y(n_1896)
);

INVx1_ASAP7_75t_L g1897 ( 
.A(n_1861),
.Y(n_1897)
);

INVx1_ASAP7_75t_L g1898 ( 
.A(n_1861),
.Y(n_1898)
);

NAND2xp5_ASAP7_75t_L g1899 ( 
.A(n_1870),
.B(n_1837),
.Y(n_1899)
);

AND2x2_ASAP7_75t_L g1900 ( 
.A(n_1864),
.B(n_1862),
.Y(n_1900)
);

INVx1_ASAP7_75t_SL g1901 ( 
.A(n_1884),
.Y(n_1901)
);

OAI22xp33_ASAP7_75t_L g1902 ( 
.A1(n_1852),
.A2(n_1823),
.B1(n_1837),
.B2(n_1832),
.Y(n_1902)
);

INVx1_ASAP7_75t_L g1903 ( 
.A(n_1865),
.Y(n_1903)
);

AND2x4_ASAP7_75t_L g1904 ( 
.A(n_1882),
.B(n_1847),
.Y(n_1904)
);

INVx2_ASAP7_75t_L g1905 ( 
.A(n_1853),
.Y(n_1905)
);

NAND2xp5_ASAP7_75t_L g1906 ( 
.A(n_1877),
.B(n_1839),
.Y(n_1906)
);

NOR2xp33_ASAP7_75t_L g1907 ( 
.A(n_1884),
.B(n_1840),
.Y(n_1907)
);

AND2x2_ASAP7_75t_L g1908 ( 
.A(n_1864),
.B(n_1862),
.Y(n_1908)
);

NAND2x1_ASAP7_75t_L g1909 ( 
.A(n_1860),
.B(n_1846),
.Y(n_1909)
);

NAND2xp5_ASAP7_75t_L g1910 ( 
.A(n_1886),
.B(n_1823),
.Y(n_1910)
);

NAND2xp5_ASAP7_75t_L g1911 ( 
.A(n_1885),
.B(n_1838),
.Y(n_1911)
);

INVx1_ASAP7_75t_L g1912 ( 
.A(n_1865),
.Y(n_1912)
);

INVx1_ASAP7_75t_SL g1913 ( 
.A(n_1864),
.Y(n_1913)
);

INVx1_ASAP7_75t_L g1914 ( 
.A(n_1872),
.Y(n_1914)
);

NOR2x1_ASAP7_75t_L g1915 ( 
.A(n_1894),
.B(n_1822),
.Y(n_1915)
);

INVxp67_ASAP7_75t_L g1916 ( 
.A(n_1878),
.Y(n_1916)
);

INVx1_ASAP7_75t_L g1917 ( 
.A(n_1872),
.Y(n_1917)
);

INVx1_ASAP7_75t_L g1918 ( 
.A(n_1874),
.Y(n_1918)
);

NAND2xp5_ASAP7_75t_L g1919 ( 
.A(n_1851),
.B(n_1838),
.Y(n_1919)
);

NAND2xp5_ASAP7_75t_L g1920 ( 
.A(n_1851),
.B(n_1838),
.Y(n_1920)
);

AND2x2_ASAP7_75t_L g1921 ( 
.A(n_1860),
.B(n_1847),
.Y(n_1921)
);

O2A1O1Ixp33_ASAP7_75t_L g1922 ( 
.A1(n_1891),
.A2(n_1832),
.B(n_1827),
.C(n_1835),
.Y(n_1922)
);

HB1xp67_ASAP7_75t_L g1923 ( 
.A(n_1874),
.Y(n_1923)
);

INVx2_ASAP7_75t_L g1924 ( 
.A(n_1853),
.Y(n_1924)
);

AND2x2_ASAP7_75t_L g1925 ( 
.A(n_1860),
.B(n_1819),
.Y(n_1925)
);

NAND2xp5_ASAP7_75t_L g1926 ( 
.A(n_1883),
.B(n_1838),
.Y(n_1926)
);

AND2x2_ASAP7_75t_L g1927 ( 
.A(n_1866),
.B(n_1819),
.Y(n_1927)
);

NOR2xp33_ASAP7_75t_L g1928 ( 
.A(n_1856),
.B(n_1846),
.Y(n_1928)
);

OR2x2_ASAP7_75t_L g1929 ( 
.A(n_1868),
.B(n_1835),
.Y(n_1929)
);

INVx1_ASAP7_75t_SL g1930 ( 
.A(n_1889),
.Y(n_1930)
);

OR2x2_ASAP7_75t_L g1931 ( 
.A(n_1868),
.B(n_1835),
.Y(n_1931)
);

OR2x2_ASAP7_75t_L g1932 ( 
.A(n_1875),
.B(n_1835),
.Y(n_1932)
);

NAND2xp5_ASAP7_75t_L g1933 ( 
.A(n_1883),
.B(n_1848),
.Y(n_1933)
);

AOI22xp33_ASAP7_75t_L g1934 ( 
.A1(n_1902),
.A2(n_1876),
.B1(n_1855),
.B2(n_1892),
.Y(n_1934)
);

NOR2x1_ASAP7_75t_L g1935 ( 
.A(n_1915),
.B(n_1822),
.Y(n_1935)
);

OR2x2_ASAP7_75t_L g1936 ( 
.A(n_1910),
.B(n_1892),
.Y(n_1936)
);

AND2x2_ASAP7_75t_L g1937 ( 
.A(n_1900),
.B(n_1866),
.Y(n_1937)
);

INVx1_ASAP7_75t_L g1938 ( 
.A(n_1923),
.Y(n_1938)
);

NOR2x1_ASAP7_75t_L g1939 ( 
.A(n_1901),
.B(n_1822),
.Y(n_1939)
);

HB1xp67_ASAP7_75t_L g1940 ( 
.A(n_1904),
.Y(n_1940)
);

INVx1_ASAP7_75t_L g1941 ( 
.A(n_1897),
.Y(n_1941)
);

AOI22xp33_ASAP7_75t_L g1942 ( 
.A1(n_1928),
.A2(n_1906),
.B1(n_1916),
.B2(n_1911),
.Y(n_1942)
);

INVx2_ASAP7_75t_L g1943 ( 
.A(n_1904),
.Y(n_1943)
);

NAND2xp5_ASAP7_75t_SL g1944 ( 
.A(n_1922),
.B(n_1819),
.Y(n_1944)
);

AND2x4_ASAP7_75t_L g1945 ( 
.A(n_1904),
.B(n_1880),
.Y(n_1945)
);

OR2x2_ASAP7_75t_L g1946 ( 
.A(n_1926),
.B(n_1867),
.Y(n_1946)
);

INVx2_ASAP7_75t_L g1947 ( 
.A(n_1927),
.Y(n_1947)
);

INVx1_ASAP7_75t_SL g1948 ( 
.A(n_1900),
.Y(n_1948)
);

NAND2xp5_ASAP7_75t_L g1949 ( 
.A(n_1899),
.B(n_1879),
.Y(n_1949)
);

INVxp67_ASAP7_75t_L g1950 ( 
.A(n_1907),
.Y(n_1950)
);

OR2x2_ASAP7_75t_L g1951 ( 
.A(n_1929),
.B(n_1931),
.Y(n_1951)
);

AND2x2_ASAP7_75t_L g1952 ( 
.A(n_1908),
.B(n_1866),
.Y(n_1952)
);

INVx1_ASAP7_75t_L g1953 ( 
.A(n_1897),
.Y(n_1953)
);

NAND2xp5_ASAP7_75t_L g1954 ( 
.A(n_1930),
.B(n_1867),
.Y(n_1954)
);

INVx1_ASAP7_75t_L g1955 ( 
.A(n_1903),
.Y(n_1955)
);

INVx1_ASAP7_75t_L g1956 ( 
.A(n_1903),
.Y(n_1956)
);

INVx1_ASAP7_75t_SL g1957 ( 
.A(n_1908),
.Y(n_1957)
);

CKINVDCx16_ASAP7_75t_R g1958 ( 
.A(n_1925),
.Y(n_1958)
);

INVx1_ASAP7_75t_L g1959 ( 
.A(n_1918),
.Y(n_1959)
);

HB1xp67_ASAP7_75t_L g1960 ( 
.A(n_1927),
.Y(n_1960)
);

BUFx2_ASAP7_75t_L g1961 ( 
.A(n_1925),
.Y(n_1961)
);

AOI221xp5_ASAP7_75t_L g1962 ( 
.A1(n_1944),
.A2(n_1913),
.B1(n_1919),
.B2(n_1920),
.C(n_1933),
.Y(n_1962)
);

NAND2xp5_ASAP7_75t_L g1963 ( 
.A(n_1938),
.B(n_1898),
.Y(n_1963)
);

INVx1_ASAP7_75t_L g1964 ( 
.A(n_1951),
.Y(n_1964)
);

NOR3xp33_ASAP7_75t_L g1965 ( 
.A(n_1950),
.B(n_1921),
.C(n_1909),
.Y(n_1965)
);

AOI21xp5_ASAP7_75t_L g1966 ( 
.A1(n_1935),
.A2(n_1909),
.B(n_1932),
.Y(n_1966)
);

AND2x2_ASAP7_75t_L g1967 ( 
.A(n_1958),
.B(n_1921),
.Y(n_1967)
);

NAND2xp5_ASAP7_75t_L g1968 ( 
.A(n_1938),
.B(n_1912),
.Y(n_1968)
);

OR2x2_ASAP7_75t_L g1969 ( 
.A(n_1951),
.B(n_1929),
.Y(n_1969)
);

AOI21xp5_ASAP7_75t_L g1970 ( 
.A1(n_1934),
.A2(n_1932),
.B(n_1931),
.Y(n_1970)
);

OR2x2_ASAP7_75t_L g1971 ( 
.A(n_1936),
.B(n_1875),
.Y(n_1971)
);

INVx1_ASAP7_75t_L g1972 ( 
.A(n_1941),
.Y(n_1972)
);

INVx1_ASAP7_75t_L g1973 ( 
.A(n_1941),
.Y(n_1973)
);

AOI22xp33_ASAP7_75t_L g1974 ( 
.A1(n_1942),
.A2(n_1880),
.B1(n_1873),
.B2(n_1827),
.Y(n_1974)
);

OAI21xp33_ASAP7_75t_SL g1975 ( 
.A1(n_1939),
.A2(n_1873),
.B(n_1889),
.Y(n_1975)
);

AOI22xp5_ASAP7_75t_L g1976 ( 
.A1(n_1958),
.A2(n_1888),
.B1(n_1895),
.B2(n_1827),
.Y(n_1976)
);

NOR2xp33_ASAP7_75t_L g1977 ( 
.A(n_1949),
.B(n_1846),
.Y(n_1977)
);

INVx1_ASAP7_75t_L g1978 ( 
.A(n_1953),
.Y(n_1978)
);

INVx1_ASAP7_75t_L g1979 ( 
.A(n_1953),
.Y(n_1979)
);

OR2x2_ASAP7_75t_L g1980 ( 
.A(n_1936),
.B(n_1881),
.Y(n_1980)
);

OAI32xp33_ASAP7_75t_L g1981 ( 
.A1(n_1948),
.A2(n_1845),
.A3(n_1918),
.B1(n_1917),
.B2(n_1914),
.Y(n_1981)
);

AOI322xp5_ASAP7_75t_L g1982 ( 
.A1(n_1940),
.A2(n_1833),
.A3(n_1871),
.B1(n_1859),
.B2(n_1848),
.C1(n_1836),
.C2(n_1888),
.Y(n_1982)
);

NOR3xp33_ASAP7_75t_L g1983 ( 
.A(n_1957),
.B(n_1826),
.C(n_1924),
.Y(n_1983)
);

AND2x2_ASAP7_75t_L g1984 ( 
.A(n_1967),
.B(n_1961),
.Y(n_1984)
);

AND2x4_ASAP7_75t_L g1985 ( 
.A(n_1964),
.B(n_1961),
.Y(n_1985)
);

INVx1_ASAP7_75t_L g1986 ( 
.A(n_1969),
.Y(n_1986)
);

INVx2_ASAP7_75t_L g1987 ( 
.A(n_1971),
.Y(n_1987)
);

AND2x2_ASAP7_75t_L g1988 ( 
.A(n_1965),
.B(n_1960),
.Y(n_1988)
);

NAND2xp5_ASAP7_75t_L g1989 ( 
.A(n_1970),
.B(n_1943),
.Y(n_1989)
);

AND2x2_ASAP7_75t_L g1990 ( 
.A(n_1983),
.B(n_1937),
.Y(n_1990)
);

AND2x2_ASAP7_75t_L g1991 ( 
.A(n_1977),
.B(n_1937),
.Y(n_1991)
);

OAI222xp33_ASAP7_75t_L g1992 ( 
.A1(n_1974),
.A2(n_1954),
.B1(n_1946),
.B2(n_1952),
.C1(n_1945),
.C2(n_1943),
.Y(n_1992)
);

INVx1_ASAP7_75t_L g1993 ( 
.A(n_1972),
.Y(n_1993)
);

NAND2xp5_ASAP7_75t_L g1994 ( 
.A(n_1962),
.B(n_1947),
.Y(n_1994)
);

OR2x2_ASAP7_75t_L g1995 ( 
.A(n_1980),
.B(n_1946),
.Y(n_1995)
);

BUFx2_ASAP7_75t_L g1996 ( 
.A(n_1975),
.Y(n_1996)
);

AND2x2_ASAP7_75t_L g1997 ( 
.A(n_1982),
.B(n_1952),
.Y(n_1997)
);

NAND2xp5_ASAP7_75t_L g1998 ( 
.A(n_1966),
.B(n_1947),
.Y(n_1998)
);

NOR3xp33_ASAP7_75t_L g1999 ( 
.A(n_1989),
.B(n_1968),
.C(n_1963),
.Y(n_1999)
);

NOR3x1_ASAP7_75t_L g2000 ( 
.A(n_1994),
.B(n_1968),
.C(n_1963),
.Y(n_2000)
);

AOI21xp5_ASAP7_75t_L g2001 ( 
.A1(n_1992),
.A2(n_1981),
.B(n_1978),
.Y(n_2001)
);

AOI31xp33_ASAP7_75t_L g2002 ( 
.A1(n_1984),
.A2(n_1979),
.A3(n_1973),
.B(n_1976),
.Y(n_2002)
);

OAI221xp5_ASAP7_75t_L g2003 ( 
.A1(n_1996),
.A2(n_1826),
.B1(n_1956),
.B2(n_1955),
.C(n_1959),
.Y(n_2003)
);

AOI21xp5_ASAP7_75t_L g2004 ( 
.A1(n_1996),
.A2(n_1945),
.B(n_1956),
.Y(n_2004)
);

AOI21xp5_ASAP7_75t_L g2005 ( 
.A1(n_1998),
.A2(n_1945),
.B(n_1955),
.Y(n_2005)
);

OAI32xp33_ASAP7_75t_L g2006 ( 
.A1(n_1997),
.A2(n_1959),
.A3(n_1845),
.B1(n_1841),
.B2(n_1905),
.Y(n_2006)
);

NAND2xp5_ASAP7_75t_L g2007 ( 
.A(n_1984),
.B(n_1871),
.Y(n_2007)
);

OAI221xp5_ASAP7_75t_L g2008 ( 
.A1(n_1986),
.A2(n_1987),
.B1(n_1995),
.B2(n_1997),
.C(n_1988),
.Y(n_2008)
);

INVx1_ASAP7_75t_SL g2009 ( 
.A(n_1985),
.Y(n_2009)
);

NAND2xp5_ASAP7_75t_L g2010 ( 
.A(n_1985),
.B(n_1859),
.Y(n_2010)
);

INVx1_ASAP7_75t_L g2011 ( 
.A(n_2009),
.Y(n_2011)
);

INVx2_ASAP7_75t_SL g2012 ( 
.A(n_2010),
.Y(n_2012)
);

AOI221xp5_ASAP7_75t_L g2013 ( 
.A1(n_2002),
.A2(n_1988),
.B1(n_1990),
.B2(n_1986),
.C(n_1985),
.Y(n_2013)
);

OAI21xp33_ASAP7_75t_L g2014 ( 
.A1(n_2007),
.A2(n_1990),
.B(n_1991),
.Y(n_2014)
);

AOI322xp5_ASAP7_75t_L g2015 ( 
.A1(n_1999),
.A2(n_1987),
.A3(n_1993),
.B1(n_1991),
.B2(n_1833),
.C1(n_1826),
.C2(n_1896),
.Y(n_2015)
);

INVx1_ASAP7_75t_L g2016 ( 
.A(n_2004),
.Y(n_2016)
);

AOI21xp5_ASAP7_75t_L g2017 ( 
.A1(n_2001),
.A2(n_1995),
.B(n_1924),
.Y(n_2017)
);

NAND2xp5_ASAP7_75t_L g2018 ( 
.A(n_2013),
.B(n_2005),
.Y(n_2018)
);

NAND2xp5_ASAP7_75t_L g2019 ( 
.A(n_2011),
.B(n_2000),
.Y(n_2019)
);

INVx1_ASAP7_75t_SL g2020 ( 
.A(n_2016),
.Y(n_2020)
);

AND2x2_ASAP7_75t_L g2021 ( 
.A(n_2012),
.B(n_2006),
.Y(n_2021)
);

INVx1_ASAP7_75t_L g2022 ( 
.A(n_2014),
.Y(n_2022)
);

INVx1_ASAP7_75t_L g2023 ( 
.A(n_2017),
.Y(n_2023)
);

INVx1_ASAP7_75t_L g2024 ( 
.A(n_2015),
.Y(n_2024)
);

NAND2xp5_ASAP7_75t_L g2025 ( 
.A(n_2013),
.B(n_2008),
.Y(n_2025)
);

NOR2x1_ASAP7_75t_L g2026 ( 
.A(n_2023),
.B(n_2003),
.Y(n_2026)
);

NOR2x1_ASAP7_75t_L g2027 ( 
.A(n_2019),
.B(n_1905),
.Y(n_2027)
);

OAI21xp5_ASAP7_75t_L g2028 ( 
.A1(n_2025),
.A2(n_1834),
.B(n_1895),
.Y(n_2028)
);

INVx1_ASAP7_75t_L g2029 ( 
.A(n_2021),
.Y(n_2029)
);

NOR2xp33_ASAP7_75t_R g2030 ( 
.A(n_2022),
.B(n_1841),
.Y(n_2030)
);

NAND2xp5_ASAP7_75t_L g2031 ( 
.A(n_2021),
.B(n_1857),
.Y(n_2031)
);

INVx3_ASAP7_75t_L g2032 ( 
.A(n_2029),
.Y(n_2032)
);

INVx1_ASAP7_75t_L g2033 ( 
.A(n_2031),
.Y(n_2033)
);

NAND4xp75_ASAP7_75t_L g2034 ( 
.A(n_2026),
.B(n_2018),
.C(n_2024),
.D(n_2020),
.Y(n_2034)
);

INVx4_ASAP7_75t_L g2035 ( 
.A(n_2032),
.Y(n_2035)
);

AOI322xp5_ASAP7_75t_L g2036 ( 
.A1(n_2035),
.A2(n_2027),
.A3(n_2032),
.B1(n_2033),
.B2(n_2034),
.C1(n_2030),
.C2(n_2028),
.Y(n_2036)
);

AND2x4_ASAP7_75t_SL g2037 ( 
.A(n_2036),
.B(n_1841),
.Y(n_2037)
);

HB1xp67_ASAP7_75t_L g2038 ( 
.A(n_2036),
.Y(n_2038)
);

BUFx2_ASAP7_75t_L g2039 ( 
.A(n_2038),
.Y(n_2039)
);

OAI21x1_ASAP7_75t_L g2040 ( 
.A1(n_2037),
.A2(n_1858),
.B(n_1854),
.Y(n_2040)
);

INVx1_ASAP7_75t_L g2041 ( 
.A(n_2039),
.Y(n_2041)
);

INVx1_ASAP7_75t_L g2042 ( 
.A(n_2040),
.Y(n_2042)
);

OAI22xp5_ASAP7_75t_L g2043 ( 
.A1(n_2041),
.A2(n_2040),
.B1(n_1854),
.B2(n_1858),
.Y(n_2043)
);

AOI21xp5_ASAP7_75t_SL g2044 ( 
.A1(n_2043),
.A2(n_2042),
.B(n_1890),
.Y(n_2044)
);

NAND2xp5_ASAP7_75t_L g2045 ( 
.A(n_2044),
.B(n_1890),
.Y(n_2045)
);

AOI22xp33_ASAP7_75t_L g2046 ( 
.A1(n_2045),
.A2(n_1863),
.B1(n_1887),
.B2(n_1869),
.Y(n_2046)
);

AOI22xp5_ASAP7_75t_L g2047 ( 
.A1(n_2046),
.A2(n_1887),
.B1(n_1869),
.B2(n_1863),
.Y(n_2047)
);

AOI211xp5_ASAP7_75t_L g2048 ( 
.A1(n_2047),
.A2(n_1896),
.B(n_1893),
.C(n_1845),
.Y(n_2048)
);


endmodule