module fake_jpeg_31011_n_152 (n_13, n_21, n_33, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_40, n_19, n_18, n_20, n_35, n_41, n_4, n_34, n_30, n_39, n_42, n_16, n_3, n_0, n_24, n_28, n_38, n_26, n_44, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_43, n_12, n_32, n_8, n_15, n_7, n_152);

input n_13;
input n_21;
input n_33;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_42;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_44;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_43;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_152;

wire n_117;
wire n_144;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_147;
wire n_73;
wire n_84;
wire n_59;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_49;
wire n_76;
wire n_127;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_103;
wire n_50;
wire n_150;
wire n_124;
wire n_141;
wire n_57;
wire n_119;
wire n_69;
wire n_83;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_106;
wire n_111;
wire n_143;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_78;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_91;
wire n_54;
wire n_93;
wire n_138;
wire n_101;
wire n_48;
wire n_149;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_135;
wire n_62;
wire n_120;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

INVx1_ASAP7_75t_L g45 ( 
.A(n_31),
.Y(n_45)
);

INVx6_ASAP7_75t_L g46 ( 
.A(n_5),
.Y(n_46)
);

BUFx12f_ASAP7_75t_L g47 ( 
.A(n_3),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_40),
.Y(n_48)
);

INVx3_ASAP7_75t_L g49 ( 
.A(n_6),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_39),
.Y(n_50)
);

BUFx12f_ASAP7_75t_L g51 ( 
.A(n_11),
.Y(n_51)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_23),
.Y(n_52)
);

BUFx5_ASAP7_75t_L g53 ( 
.A(n_32),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_5),
.Y(n_54)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_21),
.Y(n_55)
);

BUFx12f_ASAP7_75t_L g56 ( 
.A(n_37),
.Y(n_56)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_16),
.Y(n_57)
);

CKINVDCx20_ASAP7_75t_R g58 ( 
.A(n_28),
.Y(n_58)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_38),
.Y(n_59)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_27),
.Y(n_60)
);

CKINVDCx20_ASAP7_75t_R g61 ( 
.A(n_11),
.Y(n_61)
);

BUFx12f_ASAP7_75t_L g62 ( 
.A(n_8),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_48),
.Y(n_63)
);

INVx5_ASAP7_75t_L g77 ( 
.A(n_63),
.Y(n_77)
);

BUFx12f_ASAP7_75t_L g64 ( 
.A(n_54),
.Y(n_64)
);

CKINVDCx14_ASAP7_75t_R g79 ( 
.A(n_64),
.Y(n_79)
);

INVx5_ASAP7_75t_L g65 ( 
.A(n_53),
.Y(n_65)
);

BUFx3_ASAP7_75t_L g74 ( 
.A(n_65),
.Y(n_74)
);

AND2x2_ASAP7_75t_SL g66 ( 
.A(n_46),
.B(n_19),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_66),
.B(n_67),
.Y(n_72)
);

AOI21xp33_ASAP7_75t_SL g67 ( 
.A1(n_56),
.A2(n_47),
.B(n_51),
.Y(n_67)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_48),
.Y(n_68)
);

HB1xp67_ASAP7_75t_L g81 ( 
.A(n_68),
.Y(n_81)
);

CKINVDCx20_ASAP7_75t_R g69 ( 
.A(n_61),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_L g76 ( 
.A(n_69),
.B(n_50),
.Y(n_76)
);

INVx8_ASAP7_75t_L g70 ( 
.A(n_46),
.Y(n_70)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_70),
.Y(n_73)
);

INVx5_ASAP7_75t_L g71 ( 
.A(n_54),
.Y(n_71)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_71),
.Y(n_80)
);

CKINVDCx20_ASAP7_75t_R g75 ( 
.A(n_66),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_SL g90 ( 
.A(n_75),
.B(n_47),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_76),
.B(n_78),
.Y(n_86)
);

INVxp67_ASAP7_75t_L g78 ( 
.A(n_64),
.Y(n_78)
);

AOI22xp33_ASAP7_75t_L g82 ( 
.A1(n_63),
.A2(n_47),
.B1(n_49),
.B2(n_56),
.Y(n_82)
);

AOI22xp5_ASAP7_75t_L g88 ( 
.A1(n_82),
.A2(n_83),
.B1(n_84),
.B2(n_78),
.Y(n_88)
);

OA22x2_ASAP7_75t_L g83 ( 
.A1(n_70),
.A2(n_56),
.B1(n_60),
.B2(n_59),
.Y(n_83)
);

OAI22xp5_ASAP7_75t_L g84 ( 
.A1(n_68),
.A2(n_52),
.B1(n_58),
.B2(n_57),
.Y(n_84)
);

CKINVDCx12_ASAP7_75t_R g85 ( 
.A(n_67),
.Y(n_85)
);

CKINVDCx16_ASAP7_75t_R g100 ( 
.A(n_85),
.Y(n_100)
);

AND2x2_ASAP7_75t_L g87 ( 
.A(n_72),
.B(n_55),
.Y(n_87)
);

OAI21xp5_ASAP7_75t_SL g111 ( 
.A1(n_87),
.A2(n_92),
.B(n_101),
.Y(n_111)
);

OAI22xp5_ASAP7_75t_L g113 ( 
.A1(n_88),
.A2(n_2),
.B1(n_4),
.B2(n_6),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_83),
.B(n_45),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g112 ( 
.A(n_89),
.B(n_90),
.Y(n_112)
);

OAI22xp33_ASAP7_75t_L g91 ( 
.A1(n_73),
.A2(n_62),
.B1(n_51),
.B2(n_22),
.Y(n_91)
);

AOI22xp5_ASAP7_75t_L g107 ( 
.A1(n_91),
.A2(n_2),
.B1(n_3),
.B2(n_4),
.Y(n_107)
);

AND2x2_ASAP7_75t_L g92 ( 
.A(n_83),
.B(n_62),
.Y(n_92)
);

INVxp67_ASAP7_75t_L g93 ( 
.A(n_82),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g119 ( 
.A(n_93),
.B(n_95),
.Y(n_119)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_81),
.Y(n_94)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_94),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_79),
.B(n_0),
.Y(n_95)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_80),
.Y(n_96)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_96),
.Y(n_115)
);

INVx2_ASAP7_75t_SL g97 ( 
.A(n_74),
.Y(n_97)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_97),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_74),
.B(n_0),
.Y(n_98)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_98),
.Y(n_121)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_77),
.Y(n_99)
);

INVx2_ASAP7_75t_L g106 ( 
.A(n_99),
.Y(n_106)
);

AND2x2_ASAP7_75t_L g101 ( 
.A(n_77),
.B(n_1),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_75),
.B(n_1),
.Y(n_102)
);

CKINVDCx20_ASAP7_75t_R g109 ( 
.A(n_102),
.Y(n_109)
);

AND2x6_ASAP7_75t_L g103 ( 
.A(n_87),
.B(n_20),
.Y(n_103)
);

FAx1_ASAP7_75t_SL g128 ( 
.A(n_103),
.B(n_104),
.CI(n_108),
.CON(n_128),
.SN(n_128)
);

XOR2x2_ASAP7_75t_SL g104 ( 
.A(n_92),
.B(n_24),
.Y(n_104)
);

AOI22xp5_ASAP7_75t_L g132 ( 
.A1(n_107),
.A2(n_113),
.B1(n_117),
.B2(n_7),
.Y(n_132)
);

AND2x6_ASAP7_75t_L g108 ( 
.A(n_100),
.B(n_25),
.Y(n_108)
);

CKINVDCx20_ASAP7_75t_R g110 ( 
.A(n_86),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_L g123 ( 
.A(n_110),
.B(n_114),
.Y(n_123)
);

CKINVDCx20_ASAP7_75t_R g114 ( 
.A(n_101),
.Y(n_114)
);

OAI22xp5_ASAP7_75t_SL g117 ( 
.A1(n_88),
.A2(n_7),
.B1(n_8),
.B2(n_9),
.Y(n_117)
);

CKINVDCx20_ASAP7_75t_R g118 ( 
.A(n_94),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_L g136 ( 
.A(n_118),
.B(n_122),
.Y(n_136)
);

AOI21xp33_ASAP7_75t_L g120 ( 
.A1(n_91),
.A2(n_29),
.B(n_44),
.Y(n_120)
);

OAI21xp5_ASAP7_75t_SL g124 ( 
.A1(n_120),
.A2(n_93),
.B(n_9),
.Y(n_124)
);

CKINVDCx20_ASAP7_75t_R g122 ( 
.A(n_97),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_L g140 ( 
.A(n_124),
.B(n_125),
.Y(n_140)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_115),
.Y(n_125)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_105),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_L g141 ( 
.A(n_126),
.B(n_130),
.Y(n_141)
);

MAJIxp5_ASAP7_75t_L g127 ( 
.A(n_111),
.B(n_30),
.C(n_43),
.Y(n_127)
);

MAJIxp5_ASAP7_75t_L g138 ( 
.A(n_127),
.B(n_129),
.C(n_133),
.Y(n_138)
);

MAJIxp5_ASAP7_75t_L g129 ( 
.A(n_112),
.B(n_26),
.C(n_42),
.Y(n_129)
);

CKINVDCx20_ASAP7_75t_R g130 ( 
.A(n_119),
.Y(n_130)
);

CKINVDCx20_ASAP7_75t_R g131 ( 
.A(n_106),
.Y(n_131)
);

OAI21xp5_ASAP7_75t_SL g139 ( 
.A1(n_131),
.A2(n_134),
.B(n_121),
.Y(n_139)
);

XNOR2xp5_ASAP7_75t_L g137 ( 
.A(n_132),
.B(n_135),
.Y(n_137)
);

MAJIxp5_ASAP7_75t_L g133 ( 
.A(n_104),
.B(n_18),
.C(n_12),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_SL g134 ( 
.A(n_109),
.B(n_10),
.Y(n_134)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_116),
.Y(n_135)
);

NOR3xp33_ASAP7_75t_SL g144 ( 
.A(n_139),
.B(n_120),
.C(n_128),
.Y(n_144)
);

MAJIxp5_ASAP7_75t_L g142 ( 
.A(n_123),
.B(n_103),
.C(n_108),
.Y(n_142)
);

MAJIxp5_ASAP7_75t_L g145 ( 
.A(n_142),
.B(n_127),
.C(n_133),
.Y(n_145)
);

AOI22xp5_ASAP7_75t_L g143 ( 
.A1(n_137),
.A2(n_132),
.B1(n_107),
.B2(n_136),
.Y(n_143)
);

OAI22xp5_ASAP7_75t_SL g146 ( 
.A1(n_143),
.A2(n_144),
.B1(n_140),
.B2(n_141),
.Y(n_146)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_145),
.Y(n_147)
);

AOI322xp5_ASAP7_75t_L g148 ( 
.A1(n_146),
.A2(n_128),
.A3(n_129),
.B1(n_14),
.B2(n_15),
.C1(n_17),
.C2(n_33),
.Y(n_148)
);

OAI21xp5_ASAP7_75t_SL g149 ( 
.A1(n_148),
.A2(n_138),
.B(n_147),
.Y(n_149)
);

MAJIxp5_ASAP7_75t_L g150 ( 
.A(n_149),
.B(n_13),
.C(n_34),
.Y(n_150)
);

OAI21xp5_ASAP7_75t_SL g151 ( 
.A1(n_150),
.A2(n_35),
.B(n_36),
.Y(n_151)
);

XNOR2xp5_ASAP7_75t_L g152 ( 
.A(n_151),
.B(n_41),
.Y(n_152)
);


endmodule