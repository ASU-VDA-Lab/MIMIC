module fake_jpeg_20366_n_115 (n_3, n_2, n_1, n_0, n_4, n_8, n_6, n_5, n_7, n_115);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_8;
input n_6;
input n_5;
input n_7;

output n_115;

wire n_10;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_114;
wire n_74;
wire n_31;
wire n_29;
wire n_103;
wire n_50;
wire n_15;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_109;
wire n_113;
wire n_30;
wire n_106;
wire n_111;
wire n_24;
wire n_44;
wire n_17;
wire n_25;
wire n_75;
wire n_37;
wire n_102;
wire n_99;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_18;
wire n_20;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_11;
wire n_56;
wire n_79;
wire n_12;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_22;
wire n_101;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_112;
wire n_95;
wire n_97;
wire n_9;
wire n_36;
wire n_62;
wire n_43;
wire n_32;
wire n_100;
wire n_82;
wire n_96;

INVxp67_ASAP7_75t_L g9 ( 
.A(n_5),
.Y(n_9)
);

CKINVDCx20_ASAP7_75t_R g10 ( 
.A(n_4),
.Y(n_10)
);

CKINVDCx20_ASAP7_75t_R g11 ( 
.A(n_1),
.Y(n_11)
);

CKINVDCx20_ASAP7_75t_R g12 ( 
.A(n_6),
.Y(n_12)
);

INVx1_ASAP7_75t_L g13 ( 
.A(n_7),
.Y(n_13)
);

INVx2_ASAP7_75t_L g14 ( 
.A(n_3),
.Y(n_14)
);

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_3),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_6),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_0),
.Y(n_17)
);

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_14),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_18),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_14),
.Y(n_19)
);

INVx5_ASAP7_75t_L g26 ( 
.A(n_19),
.Y(n_26)
);

BUFx4f_ASAP7_75t_L g20 ( 
.A(n_14),
.Y(n_20)
);

BUFx8_ASAP7_75t_L g27 ( 
.A(n_20),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_17),
.Y(n_21)
);

NAND2xp5_ASAP7_75t_L g30 ( 
.A(n_21),
.B(n_23),
.Y(n_30)
);

INVx6_ASAP7_75t_L g22 ( 
.A(n_17),
.Y(n_22)
);

AND2x2_ASAP7_75t_L g25 ( 
.A(n_22),
.B(n_24),
.Y(n_25)
);

BUFx12f_ASAP7_75t_L g23 ( 
.A(n_9),
.Y(n_23)
);

MAJIxp5_ASAP7_75t_L g24 ( 
.A(n_11),
.B(n_0),
.C(n_1),
.Y(n_24)
);

OAI22xp33_ASAP7_75t_SL g28 ( 
.A1(n_22),
.A2(n_16),
.B1(n_15),
.B2(n_11),
.Y(n_28)
);

AOI22xp5_ASAP7_75t_L g35 ( 
.A1(n_28),
.A2(n_31),
.B1(n_12),
.B2(n_10),
.Y(n_35)
);

OAI22xp33_ASAP7_75t_SL g31 ( 
.A1(n_18),
.A2(n_16),
.B1(n_15),
.B2(n_12),
.Y(n_31)
);

HAxp5_ASAP7_75t_SL g32 ( 
.A(n_24),
.B(n_12),
.CON(n_32),
.SN(n_32)
);

OR2x2_ASAP7_75t_L g39 ( 
.A(n_32),
.B(n_10),
.Y(n_39)
);

AOI21xp5_ASAP7_75t_L g33 ( 
.A1(n_20),
.A2(n_0),
.B(n_13),
.Y(n_33)
);

INVxp67_ASAP7_75t_L g36 ( 
.A(n_33),
.Y(n_36)
);

NAND2xp5_ASAP7_75t_L g34 ( 
.A(n_25),
.B(n_20),
.Y(n_34)
);

NAND2xp5_ASAP7_75t_SL g47 ( 
.A(n_34),
.B(n_35),
.Y(n_47)
);

INVx4_ASAP7_75t_L g37 ( 
.A(n_29),
.Y(n_37)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_37),
.Y(n_46)
);

INVx4_ASAP7_75t_L g38 ( 
.A(n_29),
.Y(n_38)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_38),
.Y(n_54)
);

AND2x2_ASAP7_75t_L g53 ( 
.A(n_39),
.B(n_21),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_SL g40 ( 
.A(n_25),
.B(n_19),
.Y(n_40)
);

NAND2xp5_ASAP7_75t_SL g51 ( 
.A(n_40),
.B(n_41),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_SL g41 ( 
.A(n_25),
.B(n_32),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_30),
.Y(n_42)
);

MAJIxp5_ASAP7_75t_SL g44 ( 
.A(n_42),
.B(n_13),
.C(n_27),
.Y(n_44)
);

AOI22xp33_ASAP7_75t_L g43 ( 
.A1(n_33),
.A2(n_17),
.B1(n_13),
.B2(n_10),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_43),
.B(n_26),
.Y(n_48)
);

AND2x2_ASAP7_75t_L g58 ( 
.A(n_44),
.B(n_48),
.Y(n_58)
);

INVx2_ASAP7_75t_L g45 ( 
.A(n_37),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_45),
.B(n_49),
.Y(n_59)
);

CKINVDCx16_ASAP7_75t_R g49 ( 
.A(n_39),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_42),
.B(n_23),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_L g56 ( 
.A(n_50),
.B(n_52),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_41),
.B(n_23),
.Y(n_52)
);

OAI21xp5_ASAP7_75t_SL g63 ( 
.A1(n_53),
.A2(n_47),
.B(n_44),
.Y(n_63)
);

CKINVDCx20_ASAP7_75t_R g55 ( 
.A(n_46),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_SL g69 ( 
.A(n_55),
.B(n_65),
.Y(n_69)
);

OAI21xp5_ASAP7_75t_L g57 ( 
.A1(n_49),
.A2(n_36),
.B(n_39),
.Y(n_57)
);

OAI21xp5_ASAP7_75t_L g72 ( 
.A1(n_57),
.A2(n_62),
.B(n_63),
.Y(n_72)
);

XOR2xp5_ASAP7_75t_L g60 ( 
.A(n_51),
.B(n_34),
.Y(n_60)
);

XOR2xp5_ASAP7_75t_L g71 ( 
.A(n_60),
.B(n_27),
.Y(n_71)
);

INVx13_ASAP7_75t_L g61 ( 
.A(n_45),
.Y(n_61)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_61),
.Y(n_75)
);

OAI21xp5_ASAP7_75t_L g62 ( 
.A1(n_53),
.A2(n_40),
.B(n_43),
.Y(n_62)
);

XNOR2x2_ASAP7_75t_L g64 ( 
.A(n_53),
.B(n_35),
.Y(n_64)
);

A2O1A1O1Ixp25_ASAP7_75t_L g66 ( 
.A1(n_64),
.A2(n_26),
.B(n_27),
.C(n_37),
.D(n_38),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_SL g65 ( 
.A(n_46),
.B(n_35),
.Y(n_65)
);

OAI21xp5_ASAP7_75t_SL g84 ( 
.A1(n_66),
.A2(n_70),
.B(n_2),
.Y(n_84)
);

INVx2_ASAP7_75t_SL g67 ( 
.A(n_61),
.Y(n_67)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_67),
.Y(n_77)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_59),
.Y(n_68)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_68),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_SL g70 ( 
.A(n_56),
.B(n_60),
.Y(n_70)
);

XOR2xp5_ASAP7_75t_L g81 ( 
.A(n_71),
.B(n_54),
.Y(n_81)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_64),
.Y(n_73)
);

CKINVDCx20_ASAP7_75t_R g80 ( 
.A(n_73),
.Y(n_80)
);

OR2x2_ASAP7_75t_L g74 ( 
.A(n_58),
.B(n_38),
.Y(n_74)
);

OAI22xp5_ASAP7_75t_L g78 ( 
.A1(n_74),
.A2(n_76),
.B1(n_58),
.B2(n_54),
.Y(n_78)
);

OAI22xp5_ASAP7_75t_L g76 ( 
.A1(n_62),
.A2(n_57),
.B1(n_58),
.B2(n_63),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_SL g88 ( 
.A(n_78),
.B(n_79),
.Y(n_88)
);

NAND3xp33_ASAP7_75t_L g79 ( 
.A(n_68),
.B(n_5),
.C(n_1),
.Y(n_79)
);

XOR2xp5_ASAP7_75t_L g90 ( 
.A(n_81),
.B(n_83),
.Y(n_90)
);

OAI21xp33_ASAP7_75t_L g83 ( 
.A1(n_73),
.A2(n_0),
.B(n_2),
.Y(n_83)
);

MAJIxp5_ASAP7_75t_L g92 ( 
.A(n_84),
.B(n_72),
.C(n_71),
.Y(n_92)
);

OAI32xp33_ASAP7_75t_L g85 ( 
.A1(n_69),
.A2(n_2),
.A3(n_3),
.B1(n_4),
.B2(n_5),
.Y(n_85)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_85),
.Y(n_86)
);

INVx13_ASAP7_75t_L g87 ( 
.A(n_77),
.Y(n_87)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_87),
.Y(n_97)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_82),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g93 ( 
.A(n_89),
.B(n_91),
.Y(n_93)
);

NOR2x1_ASAP7_75t_L g91 ( 
.A(n_80),
.B(n_74),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_92),
.B(n_81),
.Y(n_94)
);

OAI21xp5_ASAP7_75t_SL g100 ( 
.A1(n_94),
.A2(n_88),
.B(n_89),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_87),
.B(n_75),
.Y(n_95)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_95),
.Y(n_101)
);

XOR2xp5_ASAP7_75t_L g96 ( 
.A(n_90),
.B(n_72),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_96),
.B(n_90),
.Y(n_99)
);

OAI22xp5_ASAP7_75t_L g98 ( 
.A1(n_86),
.A2(n_85),
.B1(n_66),
.B2(n_83),
.Y(n_98)
);

INVxp67_ASAP7_75t_L g102 ( 
.A(n_98),
.Y(n_102)
);

XOR2xp5_ASAP7_75t_L g107 ( 
.A(n_99),
.B(n_100),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_97),
.B(n_87),
.Y(n_103)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_103),
.Y(n_104)
);

OAI21x1_ASAP7_75t_L g105 ( 
.A1(n_101),
.A2(n_88),
.B(n_91),
.Y(n_105)
);

AO21x1_ASAP7_75t_SL g108 ( 
.A1(n_105),
.A2(n_91),
.B(n_93),
.Y(n_108)
);

AOI21xp5_ASAP7_75t_SL g106 ( 
.A1(n_102),
.A2(n_93),
.B(n_86),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_106),
.B(n_90),
.Y(n_109)
);

AOI22xp5_ASAP7_75t_L g111 ( 
.A1(n_108),
.A2(n_109),
.B1(n_102),
.B2(n_92),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_104),
.B(n_67),
.Y(n_110)
);

XNOR2xp5_ASAP7_75t_L g112 ( 
.A(n_110),
.B(n_107),
.Y(n_112)
);

AOI322xp5_ASAP7_75t_L g113 ( 
.A1(n_111),
.A2(n_112),
.A3(n_96),
.B1(n_6),
.B2(n_7),
.C1(n_8),
.C2(n_4),
.Y(n_113)
);

MAJIxp5_ASAP7_75t_L g114 ( 
.A(n_113),
.B(n_7),
.C(n_8),
.Y(n_114)
);

XNOR2xp5_ASAP7_75t_L g115 ( 
.A(n_114),
.B(n_8),
.Y(n_115)
);


endmodule