module fake_jpeg_12399_n_196 (n_13, n_21, n_53, n_33, n_54, n_1, n_45, n_10, n_23, n_27, n_6, n_22, n_47, n_51, n_14, n_40, n_19, n_18, n_20, n_35, n_48, n_52, n_46, n_41, n_4, n_34, n_30, n_39, n_42, n_16, n_49, n_3, n_0, n_24, n_28, n_38, n_26, n_44, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_43, n_50, n_12, n_32, n_8, n_15, n_7, n_196);

input n_13;
input n_21;
input n_53;
input n_33;
input n_54;
input n_1;
input n_45;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_47;
input n_51;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_48;
input n_52;
input n_46;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_42;
input n_16;
input n_49;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_44;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_43;
input n_50;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_196;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_64;
wire n_55;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_84;
wire n_59;
wire n_98;
wire n_178;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_127;
wire n_76;
wire n_154;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_155;
wire n_103;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_57;
wire n_171;
wire n_119;
wire n_69;
wire n_195;
wire n_83;
wire n_179;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_168;
wire n_106;
wire n_111;
wire n_186;
wire n_143;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_177;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_145;
wire n_108;
wire n_68;
wire n_94;
wire n_58;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_184;
wire n_91;
wire n_93;
wire n_161;
wire n_138;
wire n_101;
wire n_149;
wire n_157;
wire n_87;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_189;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_120;
wire n_190;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

CKINVDCx20_ASAP7_75t_R g55 ( 
.A(n_47),
.Y(n_55)
);

CKINVDCx20_ASAP7_75t_R g56 ( 
.A(n_34),
.Y(n_56)
);

INVx13_ASAP7_75t_L g57 ( 
.A(n_51),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_24),
.Y(n_58)
);

INVx6_ASAP7_75t_L g59 ( 
.A(n_29),
.Y(n_59)
);

CKINVDCx20_ASAP7_75t_R g60 ( 
.A(n_46),
.Y(n_60)
);

INVx1_ASAP7_75t_SL g61 ( 
.A(n_43),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_32),
.Y(n_62)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_38),
.Y(n_63)
);

INVx6_ASAP7_75t_L g64 ( 
.A(n_0),
.Y(n_64)
);

CKINVDCx16_ASAP7_75t_R g65 ( 
.A(n_3),
.Y(n_65)
);

BUFx3_ASAP7_75t_L g66 ( 
.A(n_18),
.Y(n_66)
);

CKINVDCx20_ASAP7_75t_R g67 ( 
.A(n_41),
.Y(n_67)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_14),
.Y(n_68)
);

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_0),
.Y(n_69)
);

BUFx3_ASAP7_75t_L g70 ( 
.A(n_9),
.Y(n_70)
);

BUFx4f_ASAP7_75t_L g71 ( 
.A(n_1),
.Y(n_71)
);

INVx8_ASAP7_75t_L g72 ( 
.A(n_44),
.Y(n_72)
);

INVx4_ASAP7_75t_L g73 ( 
.A(n_3),
.Y(n_73)
);

CKINVDCx20_ASAP7_75t_R g74 ( 
.A(n_5),
.Y(n_74)
);

CKINVDCx20_ASAP7_75t_R g75 ( 
.A(n_31),
.Y(n_75)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_27),
.Y(n_76)
);

INVx3_ASAP7_75t_L g77 ( 
.A(n_40),
.Y(n_77)
);

CKINVDCx20_ASAP7_75t_R g78 ( 
.A(n_5),
.Y(n_78)
);

BUFx6f_ASAP7_75t_L g79 ( 
.A(n_26),
.Y(n_79)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_2),
.Y(n_80)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_19),
.Y(n_81)
);

BUFx6f_ASAP7_75t_L g82 ( 
.A(n_48),
.Y(n_82)
);

CKINVDCx20_ASAP7_75t_R g83 ( 
.A(n_28),
.Y(n_83)
);

INVx2_ASAP7_75t_L g84 ( 
.A(n_71),
.Y(n_84)
);

INVx2_ASAP7_75t_L g97 ( 
.A(n_84),
.Y(n_97)
);

BUFx6f_ASAP7_75t_L g85 ( 
.A(n_58),
.Y(n_85)
);

BUFx6f_ASAP7_75t_L g99 ( 
.A(n_85),
.Y(n_99)
);

BUFx6f_ASAP7_75t_L g86 ( 
.A(n_58),
.Y(n_86)
);

BUFx6f_ASAP7_75t_L g104 ( 
.A(n_86),
.Y(n_104)
);

INVx6_ASAP7_75t_SL g87 ( 
.A(n_57),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_87),
.B(n_65),
.Y(n_105)
);

INVx2_ASAP7_75t_L g88 ( 
.A(n_71),
.Y(n_88)
);

INVx2_ASAP7_75t_L g107 ( 
.A(n_88),
.Y(n_107)
);

INVx8_ASAP7_75t_L g89 ( 
.A(n_62),
.Y(n_89)
);

BUFx2_ASAP7_75t_L g106 ( 
.A(n_89),
.Y(n_106)
);

INVx8_ASAP7_75t_L g90 ( 
.A(n_62),
.Y(n_90)
);

INVx2_ASAP7_75t_L g109 ( 
.A(n_90),
.Y(n_109)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_80),
.Y(n_91)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_91),
.Y(n_96)
);

BUFx24_ASAP7_75t_L g92 ( 
.A(n_57),
.Y(n_92)
);

AND2x2_ASAP7_75t_L g95 ( 
.A(n_92),
.B(n_61),
.Y(n_95)
);

INVx8_ASAP7_75t_L g93 ( 
.A(n_79),
.Y(n_93)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_93),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_SL g94 ( 
.A(n_87),
.B(n_78),
.Y(n_94)
);

AND2x2_ASAP7_75t_L g124 ( 
.A(n_94),
.B(n_95),
.Y(n_124)
);

OAI22xp33_ASAP7_75t_SL g98 ( 
.A1(n_85),
.A2(n_82),
.B1(n_79),
.B2(n_69),
.Y(n_98)
);

AOI22xp5_ASAP7_75t_SL g120 ( 
.A1(n_98),
.A2(n_86),
.B1(n_69),
.B2(n_64),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_L g101 ( 
.A(n_92),
.B(n_74),
.Y(n_101)
);

A2O1A1Ixp33_ASAP7_75t_L g126 ( 
.A1(n_101),
.A2(n_102),
.B(n_103),
.C(n_68),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_L g102 ( 
.A(n_92),
.B(n_83),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_L g103 ( 
.A(n_89),
.B(n_75),
.Y(n_103)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_105),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_90),
.B(n_55),
.Y(n_108)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_108),
.Y(n_116)
);

CKINVDCx20_ASAP7_75t_R g110 ( 
.A(n_95),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_L g140 ( 
.A(n_110),
.B(n_111),
.Y(n_140)
);

CKINVDCx20_ASAP7_75t_R g111 ( 
.A(n_96),
.Y(n_111)
);

INVx2_ASAP7_75t_L g112 ( 
.A(n_97),
.Y(n_112)
);

INVx2_ASAP7_75t_L g141 ( 
.A(n_112),
.Y(n_141)
);

INVx2_ASAP7_75t_SL g113 ( 
.A(n_100),
.Y(n_113)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_113),
.Y(n_134)
);

CKINVDCx20_ASAP7_75t_R g115 ( 
.A(n_106),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_L g145 ( 
.A(n_115),
.B(n_118),
.Y(n_145)
);

BUFx2_ASAP7_75t_L g117 ( 
.A(n_109),
.Y(n_117)
);

INVx1_ASAP7_75t_SL g131 ( 
.A(n_117),
.Y(n_131)
);

CKINVDCx20_ASAP7_75t_R g118 ( 
.A(n_106),
.Y(n_118)
);

INVx6_ASAP7_75t_L g119 ( 
.A(n_99),
.Y(n_119)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_119),
.Y(n_137)
);

OAI22xp5_ASAP7_75t_L g132 ( 
.A1(n_120),
.A2(n_122),
.B1(n_72),
.B2(n_77),
.Y(n_132)
);

OR2x2_ASAP7_75t_L g121 ( 
.A(n_107),
.B(n_73),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_SL g136 ( 
.A(n_121),
.B(n_126),
.Y(n_136)
);

AOI22xp33_ASAP7_75t_L g122 ( 
.A1(n_98),
.A2(n_93),
.B1(n_65),
.B2(n_70),
.Y(n_122)
);

BUFx4f_ASAP7_75t_SL g123 ( 
.A(n_99),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_L g139 ( 
.A(n_123),
.B(n_128),
.Y(n_139)
);

INVx4_ASAP7_75t_L g125 ( 
.A(n_104),
.Y(n_125)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_125),
.Y(n_142)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_104),
.Y(n_127)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_127),
.Y(n_146)
);

CKINVDCx20_ASAP7_75t_R g128 ( 
.A(n_102),
.Y(n_128)
);

AOI22xp33_ASAP7_75t_SL g129 ( 
.A1(n_106),
.A2(n_72),
.B1(n_66),
.B2(n_59),
.Y(n_129)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_96),
.Y(n_130)
);

CKINVDCx16_ASAP7_75t_R g151 ( 
.A(n_130),
.Y(n_151)
);

AOI22xp5_ASAP7_75t_L g157 ( 
.A1(n_132),
.A2(n_143),
.B1(n_45),
.B2(n_20),
.Y(n_157)
);

AOI22xp33_ASAP7_75t_SL g133 ( 
.A1(n_129),
.A2(n_81),
.B1(n_76),
.B2(n_63),
.Y(n_133)
);

INVxp67_ASAP7_75t_L g166 ( 
.A(n_133),
.Y(n_166)
);

CKINVDCx20_ASAP7_75t_R g135 ( 
.A(n_113),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_L g154 ( 
.A(n_135),
.B(n_148),
.Y(n_154)
);

AOI22xp33_ASAP7_75t_SL g138 ( 
.A1(n_117),
.A2(n_67),
.B1(n_60),
.B2(n_56),
.Y(n_138)
);

OAI22xp33_ASAP7_75t_SL g143 ( 
.A1(n_122),
.A2(n_22),
.B1(n_53),
.B2(n_52),
.Y(n_143)
);

CKINVDCx16_ASAP7_75t_R g144 ( 
.A(n_124),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_SL g162 ( 
.A(n_144),
.B(n_10),
.Y(n_162)
);

AOI22xp5_ASAP7_75t_SL g147 ( 
.A1(n_124),
.A2(n_1),
.B1(n_2),
.B2(n_4),
.Y(n_147)
);

OAI22xp5_ASAP7_75t_SL g161 ( 
.A1(n_147),
.A2(n_10),
.B1(n_11),
.B2(n_12),
.Y(n_161)
);

CKINVDCx20_ASAP7_75t_R g148 ( 
.A(n_123),
.Y(n_148)
);

MAJIxp5_ASAP7_75t_L g149 ( 
.A(n_114),
.B(n_23),
.C(n_50),
.Y(n_149)
);

MAJIxp5_ASAP7_75t_L g155 ( 
.A(n_149),
.B(n_25),
.C(n_49),
.Y(n_155)
);

AOI22xp33_ASAP7_75t_SL g150 ( 
.A1(n_116),
.A2(n_6),
.B1(n_7),
.B2(n_8),
.Y(n_150)
);

CKINVDCx20_ASAP7_75t_R g152 ( 
.A(n_145),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_L g169 ( 
.A(n_152),
.B(n_153),
.Y(n_169)
);

NOR2xp33_ASAP7_75t_L g153 ( 
.A(n_140),
.B(n_8),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_L g177 ( 
.A(n_155),
.B(n_159),
.Y(n_177)
);

MAJIxp5_ASAP7_75t_L g156 ( 
.A(n_139),
.B(n_54),
.C(n_21),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_SL g171 ( 
.A(n_156),
.B(n_165),
.Y(n_171)
);

OAI22xp5_ASAP7_75t_L g168 ( 
.A1(n_157),
.A2(n_150),
.B1(n_138),
.B2(n_133),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_L g158 ( 
.A(n_136),
.B(n_9),
.Y(n_158)
);

OR2x2_ASAP7_75t_L g174 ( 
.A(n_158),
.B(n_161),
.Y(n_174)
);

INVx13_ASAP7_75t_L g159 ( 
.A(n_131),
.Y(n_159)
);

INVxp33_ASAP7_75t_L g160 ( 
.A(n_131),
.Y(n_160)
);

OAI21xp5_ASAP7_75t_L g175 ( 
.A1(n_160),
.A2(n_164),
.B(n_167),
.Y(n_175)
);

OAI21xp5_ASAP7_75t_SL g173 ( 
.A1(n_162),
.A2(n_13),
.B(n_15),
.Y(n_173)
);

BUFx2_ASAP7_75t_L g163 ( 
.A(n_137),
.Y(n_163)
);

BUFx6f_ASAP7_75t_L g172 ( 
.A(n_163),
.Y(n_172)
);

NOR2xp33_ASAP7_75t_SL g164 ( 
.A(n_151),
.B(n_11),
.Y(n_164)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_146),
.Y(n_165)
);

CKINVDCx20_ASAP7_75t_R g167 ( 
.A(n_141),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_L g183 ( 
.A(n_168),
.B(n_170),
.Y(n_183)
);

AOI22xp5_ASAP7_75t_L g170 ( 
.A1(n_166),
.A2(n_143),
.B1(n_134),
.B2(n_142),
.Y(n_170)
);

XNOR2xp5_ASAP7_75t_L g180 ( 
.A(n_173),
.B(n_156),
.Y(n_180)
);

OAI21xp5_ASAP7_75t_L g176 ( 
.A1(n_166),
.A2(n_16),
.B(n_17),
.Y(n_176)
);

AOI21xp5_ASAP7_75t_L g182 ( 
.A1(n_176),
.A2(n_178),
.B(n_155),
.Y(n_182)
);

AOI21xp5_ASAP7_75t_L g178 ( 
.A1(n_154),
.A2(n_30),
.B(n_33),
.Y(n_178)
);

XOR2xp5_ASAP7_75t_L g179 ( 
.A(n_177),
.B(n_171),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_SL g187 ( 
.A(n_179),
.B(n_180),
.Y(n_187)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_172),
.Y(n_181)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_181),
.Y(n_186)
);

CKINVDCx20_ASAP7_75t_R g185 ( 
.A(n_182),
.Y(n_185)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_175),
.Y(n_184)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_186),
.Y(n_188)
);

OA21x2_ASAP7_75t_L g189 ( 
.A1(n_188),
.A2(n_184),
.B(n_169),
.Y(n_189)
);

MAJIxp5_ASAP7_75t_L g190 ( 
.A(n_189),
.B(n_185),
.C(n_174),
.Y(n_190)
);

XNOR2xp5_ASAP7_75t_L g191 ( 
.A(n_190),
.B(n_179),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_SL g192 ( 
.A(n_191),
.B(n_187),
.Y(n_192)
);

AOI21xp5_ASAP7_75t_L g193 ( 
.A1(n_192),
.A2(n_177),
.B(n_171),
.Y(n_193)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_193),
.Y(n_194)
);

AOI321xp33_ASAP7_75t_L g195 ( 
.A1(n_194),
.A2(n_183),
.A3(n_36),
.B1(n_37),
.B2(n_39),
.C(n_42),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_L g196 ( 
.A(n_195),
.B(n_35),
.Y(n_196)
);


endmodule