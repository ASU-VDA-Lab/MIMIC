module real_jpeg_11620_n_20 (n_17, n_8, n_0, n_2, n_10, n_9, n_12, n_6, n_11, n_14, n_7, n_18, n_3, n_5, n_4, n_1, n_19, n_16, n_15, n_13, n_20);

input n_17;
input n_8;
input n_0;
input n_2;
input n_10;
input n_9;
input n_12;
input n_6;
input n_11;
input n_14;
input n_7;
input n_18;
input n_3;
input n_5;
input n_4;
input n_1;
input n_19;
input n_16;
input n_15;
input n_13;

output n_20;

wire n_37;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_300;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_199;
wire n_95;
wire n_238;
wire n_67;
wire n_235;
wire n_107;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_123;
wire n_50;
wire n_186;
wire n_137;
wire n_72;
wire n_171;
wire n_151;
wire n_272;
wire n_198;
wire n_203;
wire n_23;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_326;
wire n_339;
wire n_80;
wire n_30;
wire n_328;
wire n_149;
wire n_332;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_230;
wire n_128;
wire n_202;
wire n_216;
wire n_127;
wire n_36;
wire n_102;
wire n_81;
wire n_101;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_252;
wire n_310;
wire n_78;
wire n_83;
wire n_288;
wire n_221;
wire n_104;
wire n_153;
wire n_337;
wire n_131;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_200;
wire n_335;
wire n_214;
wire n_113;
wire n_251;
wire n_139;
wire n_33;
wire n_338;
wire n_175;
wire n_156;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_77;
wire n_219;
wire n_122;
wire n_262;
wire n_334;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_314;
wire n_278;
wire n_103;
wire n_232;
wire n_212;
wire n_284;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_213;
wire n_25;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_341;
wire n_331;
wire n_49;
wire n_68;
wire n_146;
wire n_286;
wire n_215;
wire n_176;
wire n_166;
wire n_323;
wire n_312;
wire n_325;
wire n_307;
wire n_316;
wire n_161;
wire n_207;
wire n_237;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_140;
wire n_126;
wire n_120;
wire n_155;
wire n_319;
wire n_93;
wire n_242;
wire n_142;
wire n_76;
wire n_79;
wire n_282;
wire n_147;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_145;
wire n_266;
wire n_109;
wire n_148;
wire n_196;
wire n_298;
wire n_330;
wire n_333;
wire n_152;
wire n_270;
wire n_159;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_336;
wire n_258;
wire n_150;
wire n_41;
wire n_74;
wire n_158;
wire n_204;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_75;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_119;
wire n_283;
wire n_181;
wire n_256;
wire n_253;
wire n_273;
wire n_54;
wire n_168;
wire n_38;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_292;
wire n_64;
wire n_291;
wire n_236;
wire n_276;
wire n_287;
wire n_174;
wire n_255;
wire n_243;
wire n_299;
wire n_56;
wire n_293;
wire n_275;
wire n_227;
wire n_229;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_45;
wire n_268;
wire n_42;
wire n_313;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_143;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_303;
wire n_321;
wire n_100;
wire n_51;
wire n_205;
wire n_261;
wire n_86;
wire n_324;
wire n_70;
wire n_32;
wire n_228;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_133;
wire n_257;
wire n_210;
wire n_206;
wire n_85;
wire n_96;
wire n_308;

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_0),
.Y(n_47)
);

CKINVDCx20_ASAP7_75t_R g180 ( 
.A(n_1),
.Y(n_180)
);

AOI21xp33_ASAP7_75t_L g200 ( 
.A1(n_1),
.A2(n_65),
.B(n_201),
.Y(n_200)
);

NAND2xp5_ASAP7_75t_L g216 ( 
.A(n_1),
.B(n_191),
.Y(n_216)
);

NOR2xp33_ASAP7_75t_L g239 ( 
.A(n_1),
.B(n_63),
.Y(n_239)
);

OAI22xp33_ASAP7_75t_L g253 ( 
.A1(n_1),
.A2(n_46),
.B1(n_48),
.B2(n_180),
.Y(n_253)
);

O2A1O1Ixp33_ASAP7_75t_L g255 ( 
.A1(n_1),
.A2(n_48),
.B(n_51),
.C(n_256),
.Y(n_255)
);

NAND2xp5_ASAP7_75t_SL g259 ( 
.A(n_1),
.B(n_85),
.Y(n_259)
);

NAND2xp5_ASAP7_75t_L g277 ( 
.A(n_1),
.B(n_38),
.Y(n_277)
);

NAND2xp5_ASAP7_75t_L g280 ( 
.A(n_1),
.B(n_56),
.Y(n_280)
);

AOI21xp33_ASAP7_75t_L g289 ( 
.A1(n_1),
.A2(n_63),
.B(n_239),
.Y(n_289)
);

OAI22xp5_ASAP7_75t_L g54 ( 
.A1(n_2),
.A2(n_46),
.B1(n_48),
.B2(n_55),
.Y(n_54)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_2),
.Y(n_55)
);

AOI22xp33_ASAP7_75t_L g98 ( 
.A1(n_2),
.A2(n_55),
.B1(n_60),
.B2(n_63),
.Y(n_98)
);

AOI22xp33_ASAP7_75t_L g116 ( 
.A1(n_2),
.A2(n_34),
.B1(n_41),
.B2(n_55),
.Y(n_116)
);

OAI22xp5_ASAP7_75t_L g322 ( 
.A1(n_2),
.A2(n_55),
.B1(n_65),
.B2(n_66),
.Y(n_322)
);

BUFx12f_ASAP7_75t_L g60 ( 
.A(n_3),
.Y(n_60)
);

AOI22xp33_ASAP7_75t_SL g76 ( 
.A1(n_4),
.A2(n_60),
.B1(n_63),
.B2(n_77),
.Y(n_76)
);

CKINVDCx20_ASAP7_75t_R g77 ( 
.A(n_4),
.Y(n_77)
);

AOI22xp33_ASAP7_75t_SL g91 ( 
.A1(n_4),
.A2(n_65),
.B1(n_66),
.B2(n_77),
.Y(n_91)
);

AOI22xp33_ASAP7_75t_L g120 ( 
.A1(n_4),
.A2(n_46),
.B1(n_48),
.B2(n_77),
.Y(n_120)
);

OAI22xp5_ASAP7_75t_L g176 ( 
.A1(n_4),
.A2(n_34),
.B1(n_41),
.B2(n_77),
.Y(n_176)
);

BUFx8_ASAP7_75t_L g62 ( 
.A(n_5),
.Y(n_62)
);

INVx11_ASAP7_75t_L g36 ( 
.A(n_6),
.Y(n_36)
);

OAI22xp5_ASAP7_75t_L g44 ( 
.A1(n_7),
.A2(n_45),
.B1(n_46),
.B2(n_48),
.Y(n_44)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_7),
.Y(n_45)
);

OAI22xp5_ASAP7_75t_L g84 ( 
.A1(n_7),
.A2(n_45),
.B1(n_60),
.B2(n_63),
.Y(n_84)
);

AOI22xp33_ASAP7_75t_SL g138 ( 
.A1(n_7),
.A2(n_45),
.B1(n_65),
.B2(n_66),
.Y(n_138)
);

OAI22xp5_ASAP7_75t_L g152 ( 
.A1(n_7),
.A2(n_34),
.B1(n_41),
.B2(n_45),
.Y(n_152)
);

BUFx12_ASAP7_75t_L g67 ( 
.A(n_8),
.Y(n_67)
);

BUFx12_ASAP7_75t_L g81 ( 
.A(n_9),
.Y(n_81)
);

OAI22xp5_ASAP7_75t_L g39 ( 
.A1(n_10),
.A2(n_34),
.B1(n_40),
.B2(n_41),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_10),
.Y(n_40)
);

OAI22xp5_ASAP7_75t_SL g87 ( 
.A1(n_10),
.A2(n_40),
.B1(n_46),
.B2(n_48),
.Y(n_87)
);

AOI22xp33_ASAP7_75t_SL g136 ( 
.A1(n_10),
.A2(n_40),
.B1(n_60),
.B2(n_63),
.Y(n_136)
);

OAI22xp5_ASAP7_75t_SL g329 ( 
.A1(n_10),
.A2(n_40),
.B1(n_65),
.B2(n_66),
.Y(n_329)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_11),
.Y(n_341)
);

AOI22xp33_ASAP7_75t_SL g160 ( 
.A1(n_12),
.A2(n_65),
.B1(n_66),
.B2(n_161),
.Y(n_160)
);

CKINVDCx20_ASAP7_75t_R g161 ( 
.A(n_12),
.Y(n_161)
);

AOI22xp33_ASAP7_75t_SL g204 ( 
.A1(n_12),
.A2(n_60),
.B1(n_63),
.B2(n_161),
.Y(n_204)
);

OAI22xp5_ASAP7_75t_L g261 ( 
.A1(n_12),
.A2(n_46),
.B1(n_48),
.B2(n_161),
.Y(n_261)
);

OAI22xp33_ASAP7_75t_SL g268 ( 
.A1(n_12),
.A2(n_34),
.B1(n_41),
.B2(n_161),
.Y(n_268)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_13),
.Y(n_38)
);

BUFx16f_ASAP7_75t_L g51 ( 
.A(n_14),
.Y(n_51)
);

AOI22xp33_ASAP7_75t_L g187 ( 
.A1(n_15),
.A2(n_65),
.B1(n_66),
.B2(n_188),
.Y(n_187)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_15),
.Y(n_188)
);

AOI22xp33_ASAP7_75t_SL g214 ( 
.A1(n_15),
.A2(n_60),
.B1(n_63),
.B2(n_188),
.Y(n_214)
);

OAI22xp5_ASAP7_75t_L g254 ( 
.A1(n_15),
.A2(n_46),
.B1(n_48),
.B2(n_188),
.Y(n_254)
);

OAI22xp33_ASAP7_75t_SL g275 ( 
.A1(n_15),
.A2(n_34),
.B1(n_41),
.B2(n_188),
.Y(n_275)
);

AOI22xp33_ASAP7_75t_SL g68 ( 
.A1(n_16),
.A2(n_65),
.B1(n_66),
.B2(n_69),
.Y(n_68)
);

CKINVDCx20_ASAP7_75t_R g69 ( 
.A(n_16),
.Y(n_69)
);

AOI22xp33_ASAP7_75t_SL g158 ( 
.A1(n_16),
.A2(n_60),
.B1(n_63),
.B2(n_69),
.Y(n_158)
);

OAI22xp5_ASAP7_75t_L g206 ( 
.A1(n_16),
.A2(n_46),
.B1(n_48),
.B2(n_69),
.Y(n_206)
);

OAI22xp5_ASAP7_75t_SL g242 ( 
.A1(n_16),
.A2(n_34),
.B1(n_41),
.B2(n_69),
.Y(n_242)
);

AOI22xp33_ASAP7_75t_SL g124 ( 
.A1(n_17),
.A2(n_65),
.B1(n_66),
.B2(n_125),
.Y(n_124)
);

CKINVDCx20_ASAP7_75t_R g125 ( 
.A(n_17),
.Y(n_125)
);

AOI22xp33_ASAP7_75t_SL g183 ( 
.A1(n_17),
.A2(n_60),
.B1(n_63),
.B2(n_125),
.Y(n_183)
);

AOI22xp33_ASAP7_75t_SL g233 ( 
.A1(n_17),
.A2(n_46),
.B1(n_48),
.B2(n_125),
.Y(n_233)
);

OAI22xp5_ASAP7_75t_SL g263 ( 
.A1(n_17),
.A2(n_34),
.B1(n_41),
.B2(n_125),
.Y(n_263)
);

AOI22xp33_ASAP7_75t_SL g70 ( 
.A1(n_18),
.A2(n_65),
.B1(n_66),
.B2(n_71),
.Y(n_70)
);

CKINVDCx20_ASAP7_75t_R g71 ( 
.A(n_18),
.Y(n_71)
);

AOI22xp33_ASAP7_75t_SL g122 ( 
.A1(n_18),
.A2(n_60),
.B1(n_63),
.B2(n_71),
.Y(n_122)
);

OAI22xp5_ASAP7_75t_L g155 ( 
.A1(n_18),
.A2(n_46),
.B1(n_48),
.B2(n_71),
.Y(n_155)
);

OAI22xp5_ASAP7_75t_L g218 ( 
.A1(n_18),
.A2(n_34),
.B1(n_41),
.B2(n_71),
.Y(n_218)
);

AOI21xp5_ASAP7_75t_L g20 ( 
.A1(n_19),
.A2(n_21),
.B(n_340),
.Y(n_20)
);

NOR2xp33_ASAP7_75t_L g340 ( 
.A(n_19),
.B(n_341),
.Y(n_340)
);

AOI21xp33_ASAP7_75t_L g21 ( 
.A1(n_22),
.A2(n_335),
.B(n_338),
.Y(n_21)
);

OAI21xp5_ASAP7_75t_L g22 ( 
.A1(n_23),
.A2(n_327),
.B(n_331),
.Y(n_22)
);

AOI21xp5_ASAP7_75t_L g23 ( 
.A1(n_24),
.A2(n_314),
.B(n_326),
.Y(n_23)
);

AO21x1_ASAP7_75t_L g24 ( 
.A1(n_25),
.A2(n_139),
.B(n_311),
.Y(n_24)
);

NOR2xp33_ASAP7_75t_L g25 ( 
.A(n_26),
.B(n_126),
.Y(n_25)
);

NOR2xp33_ASAP7_75t_SL g26 ( 
.A(n_27),
.B(n_102),
.Y(n_26)
);

NAND2xp5_ASAP7_75t_L g312 ( 
.A(n_27),
.B(n_102),
.Y(n_312)
);

XOR2xp5_ASAP7_75t_L g27 ( 
.A(n_28),
.B(n_72),
.Y(n_27)
);

MAJIxp5_ASAP7_75t_L g127 ( 
.A(n_28),
.B(n_88),
.C(n_100),
.Y(n_127)
);

OAI21xp5_ASAP7_75t_L g28 ( 
.A1(n_29),
.A2(n_32),
.B(n_57),
.Y(n_28)
);

OAI22xp5_ASAP7_75t_L g104 ( 
.A1(n_29),
.A2(n_30),
.B1(n_105),
.B2(n_106),
.Y(n_104)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_30),
.Y(n_29)
);

NAND2xp5_ASAP7_75t_L g30 ( 
.A(n_31),
.B(n_42),
.Y(n_30)
);

AOI22xp5_ASAP7_75t_L g106 ( 
.A1(n_31),
.A2(n_32),
.B1(n_57),
.B2(n_107),
.Y(n_106)
);

AOI22xp5_ASAP7_75t_L g145 ( 
.A1(n_31),
.A2(n_32),
.B1(n_42),
.B2(n_43),
.Y(n_145)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_32),
.Y(n_31)
);

OAI21xp5_ASAP7_75t_SL g32 ( 
.A1(n_33),
.A2(n_38),
.B(n_39),
.Y(n_32)
);

AOI22xp5_ASAP7_75t_L g114 ( 
.A1(n_33),
.A2(n_38),
.B1(n_39),
.B2(n_115),
.Y(n_114)
);

CKINVDCx20_ASAP7_75t_R g150 ( 
.A(n_33),
.Y(n_150)
);

AOI22xp5_ASAP7_75t_L g175 ( 
.A1(n_33),
.A2(n_38),
.B1(n_152),
.B2(n_176),
.Y(n_175)
);

AOI22xp5_ASAP7_75t_L g217 ( 
.A1(n_33),
.A2(n_38),
.B1(n_176),
.B2(n_218),
.Y(n_217)
);

AOI22xp5_ASAP7_75t_L g241 ( 
.A1(n_33),
.A2(n_38),
.B1(n_218),
.B2(n_242),
.Y(n_241)
);

AOI22xp5_ASAP7_75t_SL g262 ( 
.A1(n_33),
.A2(n_38),
.B1(n_242),
.B2(n_263),
.Y(n_262)
);

AOI22xp5_ASAP7_75t_SL g274 ( 
.A1(n_33),
.A2(n_38),
.B1(n_180),
.B2(n_275),
.Y(n_274)
);

AOI22xp33_ASAP7_75t_L g279 ( 
.A1(n_33),
.A2(n_38),
.B1(n_268),
.B2(n_275),
.Y(n_279)
);

AND2x2_ASAP7_75t_L g33 ( 
.A(n_34),
.B(n_37),
.Y(n_33)
);

INVx11_ASAP7_75t_L g41 ( 
.A(n_34),
.Y(n_41)
);

OA22x2_ASAP7_75t_L g53 ( 
.A1(n_34),
.A2(n_41),
.B1(n_51),
.B2(n_52),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_SL g276 ( 
.A(n_34),
.B(n_277),
.Y(n_276)
);

BUFx12f_ASAP7_75t_L g34 ( 
.A(n_35),
.Y(n_34)
);

INVx8_ASAP7_75t_L g35 ( 
.A(n_36),
.Y(n_35)
);

OAI22xp5_ASAP7_75t_L g149 ( 
.A1(n_37),
.A2(n_116),
.B1(n_150),
.B2(n_151),
.Y(n_149)
);

OAI22xp5_ASAP7_75t_SL g266 ( 
.A1(n_37),
.A2(n_150),
.B1(n_267),
.B2(n_269),
.Y(n_266)
);

INVx2_ASAP7_75t_L g37 ( 
.A(n_38),
.Y(n_37)
);

OAI21xp33_ASAP7_75t_L g256 ( 
.A1(n_41),
.A2(n_52),
.B(n_180),
.Y(n_256)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_43),
.Y(n_42)
);

AOI22xp5_ASAP7_75t_L g43 ( 
.A1(n_44),
.A2(n_49),
.B1(n_54),
.B2(n_56),
.Y(n_43)
);

AOI22xp5_ASAP7_75t_L g118 ( 
.A1(n_44),
.A2(n_49),
.B1(n_56),
.B2(n_119),
.Y(n_118)
);

INVx4_ASAP7_75t_L g48 ( 
.A(n_46),
.Y(n_48)
);

OAI22xp33_ASAP7_75t_L g50 ( 
.A1(n_46),
.A2(n_48),
.B1(n_51),
.B2(n_52),
.Y(n_50)
);

OA22x2_ASAP7_75t_L g83 ( 
.A1(n_46),
.A2(n_48),
.B1(n_81),
.B2(n_82),
.Y(n_83)
);

OAI32xp33_ASAP7_75t_L g237 ( 
.A1(n_46),
.A2(n_63),
.A3(n_81),
.B1(n_238),
.B2(n_240),
.Y(n_237)
);

BUFx12f_ASAP7_75t_L g46 ( 
.A(n_47),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g240 ( 
.A(n_48),
.B(n_82),
.Y(n_240)
);

AOI22xp5_ASAP7_75t_L g86 ( 
.A1(n_49),
.A2(n_54),
.B1(n_56),
.B2(n_87),
.Y(n_86)
);

OAI21xp5_ASAP7_75t_L g94 ( 
.A1(n_49),
.A2(n_56),
.B(n_87),
.Y(n_94)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_49),
.Y(n_156)
);

AOI22xp5_ASAP7_75t_L g205 ( 
.A1(n_49),
.A2(n_56),
.B1(n_155),
.B2(n_206),
.Y(n_205)
);

AOI22xp5_ASAP7_75t_L g231 ( 
.A1(n_49),
.A2(n_56),
.B1(n_206),
.B2(n_232),
.Y(n_231)
);

AOI22xp5_ASAP7_75t_L g252 ( 
.A1(n_49),
.A2(n_56),
.B1(n_253),
.B2(n_254),
.Y(n_252)
);

AOI22xp5_ASAP7_75t_L g260 ( 
.A1(n_49),
.A2(n_56),
.B1(n_254),
.B2(n_261),
.Y(n_260)
);

AND2x2_ASAP7_75t_L g49 ( 
.A(n_50),
.B(n_53),
.Y(n_49)
);

INVx6_ASAP7_75t_L g52 ( 
.A(n_51),
.Y(n_52)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_53),
.Y(n_56)
);

OAI22xp5_ASAP7_75t_L g153 ( 
.A1(n_53),
.A2(n_120),
.B1(n_154),
.B2(n_156),
.Y(n_153)
);

OAI22xp5_ASAP7_75t_SL g290 ( 
.A1(n_53),
.A2(n_156),
.B1(n_233),
.B2(n_291),
.Y(n_290)
);

CKINVDCx14_ASAP7_75t_R g107 ( 
.A(n_57),
.Y(n_107)
);

OAI22xp5_ASAP7_75t_SL g57 ( 
.A1(n_58),
.A2(n_59),
.B1(n_68),
.B2(n_70),
.Y(n_57)
);

OAI22xp5_ASAP7_75t_L g90 ( 
.A1(n_58),
.A2(n_59),
.B1(n_70),
.B2(n_91),
.Y(n_90)
);

OAI22xp5_ASAP7_75t_SL g123 ( 
.A1(n_58),
.A2(n_59),
.B1(n_68),
.B2(n_124),
.Y(n_123)
);

OAI22xp5_ASAP7_75t_SL g137 ( 
.A1(n_58),
.A2(n_59),
.B1(n_91),
.B2(n_138),
.Y(n_137)
);

OAI22xp5_ASAP7_75t_SL g159 ( 
.A1(n_58),
.A2(n_59),
.B1(n_124),
.B2(n_160),
.Y(n_159)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_58),
.Y(n_189)
);

OAI22xp5_ASAP7_75t_SL g199 ( 
.A1(n_58),
.A2(n_59),
.B1(n_187),
.B2(n_200),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_SL g58 ( 
.A(n_59),
.B(n_64),
.Y(n_58)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_59),
.Y(n_191)
);

OA22x2_ASAP7_75t_L g59 ( 
.A1(n_60),
.A2(n_61),
.B1(n_62),
.B2(n_63),
.Y(n_59)
);

INVx8_ASAP7_75t_L g63 ( 
.A(n_60),
.Y(n_63)
);

OAI22xp5_ASAP7_75t_SL g80 ( 
.A1(n_60),
.A2(n_63),
.B1(n_81),
.B2(n_82),
.Y(n_80)
);

OAI32xp33_ASAP7_75t_L g177 ( 
.A1(n_60),
.A2(n_62),
.A3(n_65),
.B1(n_178),
.B2(n_179),
.Y(n_177)
);

OAI22xp5_ASAP7_75t_SL g64 ( 
.A1(n_61),
.A2(n_62),
.B1(n_65),
.B2(n_66),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g178 ( 
.A(n_61),
.B(n_63),
.Y(n_178)
);

INVx11_ASAP7_75t_L g61 ( 
.A(n_62),
.Y(n_61)
);

INVx6_ASAP7_75t_L g65 ( 
.A(n_66),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_SL g179 ( 
.A(n_66),
.B(n_180),
.Y(n_179)
);

BUFx16f_ASAP7_75t_L g66 ( 
.A(n_67),
.Y(n_66)
);

AOI22xp5_ASAP7_75t_L g72 ( 
.A1(n_73),
.A2(n_88),
.B1(n_100),
.B2(n_101),
.Y(n_72)
);

CKINVDCx20_ASAP7_75t_R g100 ( 
.A(n_73),
.Y(n_100)
);

OAI21xp33_ASAP7_75t_L g109 ( 
.A1(n_73),
.A2(n_74),
.B(n_86),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_SL g73 ( 
.A(n_74),
.B(n_86),
.Y(n_73)
);

AOI22xp5_ASAP7_75t_L g74 ( 
.A1(n_75),
.A2(n_78),
.B1(n_84),
.B2(n_85),
.Y(n_74)
);

INVxp67_ASAP7_75t_L g75 ( 
.A(n_76),
.Y(n_75)
);

OAI22xp5_ASAP7_75t_SL g121 ( 
.A1(n_76),
.A2(n_79),
.B1(n_83),
.B2(n_122),
.Y(n_121)
);

AOI22xp5_ASAP7_75t_L g96 ( 
.A1(n_78),
.A2(n_84),
.B1(n_85),
.B2(n_97),
.Y(n_96)
);

AOI22xp5_ASAP7_75t_L g181 ( 
.A1(n_78),
.A2(n_85),
.B1(n_182),
.B2(n_184),
.Y(n_181)
);

AOI22xp5_ASAP7_75t_L g212 ( 
.A1(n_78),
.A2(n_85),
.B1(n_213),
.B2(n_215),
.Y(n_212)
);

OAI21xp5_ASAP7_75t_SL g318 ( 
.A1(n_78),
.A2(n_85),
.B(n_319),
.Y(n_318)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_79),
.Y(n_78)
);

OAI22xp5_ASAP7_75t_SL g135 ( 
.A1(n_79),
.A2(n_83),
.B1(n_98),
.B2(n_136),
.Y(n_135)
);

OAI22xp5_ASAP7_75t_SL g157 ( 
.A1(n_79),
.A2(n_83),
.B1(n_122),
.B2(n_158),
.Y(n_157)
);

OAI22xp5_ASAP7_75t_SL g203 ( 
.A1(n_79),
.A2(n_83),
.B1(n_183),
.B2(n_204),
.Y(n_203)
);

OAI22xp5_ASAP7_75t_SL g288 ( 
.A1(n_79),
.A2(n_83),
.B1(n_214),
.B2(n_289),
.Y(n_288)
);

NAND2xp5_ASAP7_75t_L g79 ( 
.A(n_80),
.B(n_83),
.Y(n_79)
);

INVx8_ASAP7_75t_L g82 ( 
.A(n_81),
.Y(n_82)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_83),
.Y(n_85)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_88),
.Y(n_101)
);

AOI22xp5_ASAP7_75t_L g88 ( 
.A1(n_89),
.A2(n_90),
.B1(n_92),
.B2(n_93),
.Y(n_88)
);

AOI22xp5_ASAP7_75t_SL g130 ( 
.A1(n_89),
.A2(n_90),
.B1(n_131),
.B2(n_132),
.Y(n_130)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_90),
.Y(n_89)
);

MAJIxp5_ASAP7_75t_L g129 ( 
.A(n_90),
.B(n_94),
.C(n_96),
.Y(n_129)
);

MAJIxp5_ASAP7_75t_L g315 ( 
.A(n_90),
.B(n_129),
.C(n_132),
.Y(n_315)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_93),
.Y(n_92)
);

OAI22xp5_ASAP7_75t_SL g93 ( 
.A1(n_94),
.A2(n_95),
.B1(n_96),
.B2(n_99),
.Y(n_93)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_94),
.Y(n_99)
);

AOI22xp5_ASAP7_75t_L g133 ( 
.A1(n_94),
.A2(n_99),
.B1(n_134),
.B2(n_135),
.Y(n_133)
);

MAJIxp5_ASAP7_75t_L g325 ( 
.A(n_94),
.B(n_135),
.C(n_137),
.Y(n_325)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_96),
.Y(n_95)
);

CKINVDCx14_ASAP7_75t_R g97 ( 
.A(n_98),
.Y(n_97)
);

MAJIxp5_ASAP7_75t_L g102 ( 
.A(n_103),
.B(n_108),
.C(n_110),
.Y(n_102)
);

AOI22xp5_ASAP7_75t_L g163 ( 
.A1(n_103),
.A2(n_104),
.B1(n_108),
.B2(n_109),
.Y(n_163)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_104),
.Y(n_103)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_106),
.Y(n_105)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_109),
.Y(n_108)
);

XOR2xp5_ASAP7_75t_L g162 ( 
.A(n_110),
.B(n_163),
.Y(n_162)
);

MAJIxp5_ASAP7_75t_L g110 ( 
.A(n_111),
.B(n_121),
.C(n_123),
.Y(n_110)
);

AOI22xp5_ASAP7_75t_L g142 ( 
.A1(n_111),
.A2(n_112),
.B1(n_143),
.B2(n_144),
.Y(n_142)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_112),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_L g112 ( 
.A(n_113),
.B(n_117),
.Y(n_112)
);

OAI22xp5_ASAP7_75t_SL g171 ( 
.A1(n_113),
.A2(n_114),
.B1(n_117),
.B2(n_118),
.Y(n_171)
);

CKINVDCx14_ASAP7_75t_R g113 ( 
.A(n_114),
.Y(n_113)
);

INVxp67_ASAP7_75t_L g115 ( 
.A(n_116),
.Y(n_115)
);

CKINVDCx14_ASAP7_75t_R g117 ( 
.A(n_118),
.Y(n_117)
);

INVxp67_ASAP7_75t_L g119 ( 
.A(n_120),
.Y(n_119)
);

XOR2xp5_ASAP7_75t_L g144 ( 
.A(n_121),
.B(n_123),
.Y(n_144)
);

OAI21xp5_ASAP7_75t_L g311 ( 
.A1(n_126),
.A2(n_312),
.B(n_313),
.Y(n_311)
);

NOR2xp33_ASAP7_75t_L g126 ( 
.A(n_127),
.B(n_128),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_L g313 ( 
.A(n_127),
.B(n_128),
.Y(n_313)
);

XNOR2xp5_ASAP7_75t_L g128 ( 
.A(n_129),
.B(n_130),
.Y(n_128)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_132),
.Y(n_131)
);

XNOR2xp5_ASAP7_75t_L g132 ( 
.A(n_133),
.B(n_137),
.Y(n_132)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_135),
.Y(n_134)
);

CKINVDCx16_ASAP7_75t_R g319 ( 
.A(n_136),
.Y(n_319)
);

CKINVDCx20_ASAP7_75t_R g321 ( 
.A(n_138),
.Y(n_321)
);

OAI21xp5_ASAP7_75t_L g139 ( 
.A1(n_140),
.A2(n_164),
.B(n_310),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_L g140 ( 
.A(n_141),
.B(n_162),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_L g310 ( 
.A(n_141),
.B(n_162),
.Y(n_310)
);

MAJIxp5_ASAP7_75t_L g141 ( 
.A(n_142),
.B(n_145),
.C(n_146),
.Y(n_141)
);

XNOR2xp5_ASAP7_75t_L g193 ( 
.A(n_142),
.B(n_145),
.Y(n_193)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_144),
.Y(n_143)
);

XNOR2xp5_ASAP7_75t_L g192 ( 
.A(n_146),
.B(n_193),
.Y(n_192)
);

MAJIxp5_ASAP7_75t_L g146 ( 
.A(n_147),
.B(n_157),
.C(n_159),
.Y(n_146)
);

AOI22xp5_ASAP7_75t_L g168 ( 
.A1(n_147),
.A2(n_148),
.B1(n_169),
.B2(n_170),
.Y(n_168)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_148),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_L g148 ( 
.A(n_149),
.B(n_153),
.Y(n_148)
);

XNOR2xp5_ASAP7_75t_L g222 ( 
.A(n_149),
.B(n_153),
.Y(n_222)
);

CKINVDCx16_ASAP7_75t_R g151 ( 
.A(n_152),
.Y(n_151)
);

CKINVDCx16_ASAP7_75t_R g154 ( 
.A(n_155),
.Y(n_154)
);

XOR2xp5_ASAP7_75t_L g170 ( 
.A(n_157),
.B(n_159),
.Y(n_170)
);

INVxp67_ASAP7_75t_L g184 ( 
.A(n_158),
.Y(n_184)
);

INVxp67_ASAP7_75t_L g190 ( 
.A(n_160),
.Y(n_190)
);

AOI21xp5_ASAP7_75t_SL g164 ( 
.A1(n_165),
.A2(n_194),
.B(n_309),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_L g165 ( 
.A(n_166),
.B(n_192),
.Y(n_165)
);

NOR2xp33_ASAP7_75t_L g309 ( 
.A(n_166),
.B(n_192),
.Y(n_309)
);

MAJIxp5_ASAP7_75t_L g166 ( 
.A(n_167),
.B(n_171),
.C(n_172),
.Y(n_166)
);

AOI22xp5_ASAP7_75t_L g306 ( 
.A1(n_167),
.A2(n_168),
.B1(n_171),
.B2(n_307),
.Y(n_306)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_168),
.Y(n_167)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_170),
.Y(n_169)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_171),
.Y(n_307)
);

XNOR2xp5_ASAP7_75t_L g305 ( 
.A(n_172),
.B(n_306),
.Y(n_305)
);

MAJIxp5_ASAP7_75t_L g172 ( 
.A(n_173),
.B(n_181),
.C(n_185),
.Y(n_172)
);

XOR2xp5_ASAP7_75t_L g223 ( 
.A(n_173),
.B(n_224),
.Y(n_223)
);

NAND2xp5_ASAP7_75t_SL g173 ( 
.A(n_174),
.B(n_177),
.Y(n_173)
);

OAI22xp5_ASAP7_75t_SL g209 ( 
.A1(n_174),
.A2(n_175),
.B1(n_177),
.B2(n_210),
.Y(n_209)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_175),
.Y(n_174)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_177),
.Y(n_210)
);

INVxp67_ASAP7_75t_L g201 ( 
.A(n_179),
.Y(n_201)
);

XOR2xp5_ASAP7_75t_L g224 ( 
.A(n_181),
.B(n_185),
.Y(n_224)
);

INVxp67_ASAP7_75t_L g182 ( 
.A(n_183),
.Y(n_182)
);

AOI22xp5_ASAP7_75t_L g185 ( 
.A1(n_186),
.A2(n_189),
.B1(n_190),
.B2(n_191),
.Y(n_185)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_187),
.Y(n_186)
);

AOI22xp5_ASAP7_75t_L g320 ( 
.A1(n_189),
.A2(n_191),
.B1(n_321),
.B2(n_322),
.Y(n_320)
);

AOI22xp5_ASAP7_75t_SL g328 ( 
.A1(n_189),
.A2(n_191),
.B1(n_322),
.B2(n_329),
.Y(n_328)
);

OAI21xp5_ASAP7_75t_L g337 ( 
.A1(n_189),
.A2(n_191),
.B(n_329),
.Y(n_337)
);

A2O1A1Ixp33_ASAP7_75t_SL g194 ( 
.A1(n_195),
.A2(n_225),
.B(n_303),
.C(n_308),
.Y(n_194)
);

OR2x2_ASAP7_75t_L g195 ( 
.A(n_196),
.B(n_219),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_L g302 ( 
.A(n_196),
.B(n_219),
.Y(n_302)
);

MAJIxp5_ASAP7_75t_L g196 ( 
.A(n_197),
.B(n_209),
.C(n_211),
.Y(n_196)
);

OAI22xp5_ASAP7_75t_SL g243 ( 
.A1(n_197),
.A2(n_198),
.B1(n_244),
.B2(n_245),
.Y(n_243)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_198),
.Y(n_197)
);

XOR2xp5_ASAP7_75t_L g198 ( 
.A(n_199),
.B(n_202),
.Y(n_198)
);

MAJIxp5_ASAP7_75t_L g221 ( 
.A(n_199),
.B(n_203),
.C(n_208),
.Y(n_221)
);

AOI22xp5_ASAP7_75t_L g202 ( 
.A1(n_203),
.A2(n_205),
.B1(n_207),
.B2(n_208),
.Y(n_202)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_203),
.Y(n_207)
);

INVxp67_ASAP7_75t_L g215 ( 
.A(n_204),
.Y(n_215)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_205),
.Y(n_208)
);

XNOR2xp5_ASAP7_75t_SL g244 ( 
.A(n_209),
.B(n_211),
.Y(n_244)
);

MAJIxp5_ASAP7_75t_L g211 ( 
.A(n_212),
.B(n_216),
.C(n_217),
.Y(n_211)
);

XNOR2xp5_ASAP7_75t_SL g229 ( 
.A(n_212),
.B(n_230),
.Y(n_229)
);

INVxp67_ASAP7_75t_L g213 ( 
.A(n_214),
.Y(n_213)
);

XNOR2xp5_ASAP7_75t_L g230 ( 
.A(n_216),
.B(n_217),
.Y(n_230)
);

XNOR2xp5_ASAP7_75t_L g219 ( 
.A(n_220),
.B(n_223),
.Y(n_219)
);

XNOR2xp5_ASAP7_75t_L g220 ( 
.A(n_221),
.B(n_222),
.Y(n_220)
);

MAJIxp5_ASAP7_75t_L g304 ( 
.A(n_221),
.B(n_222),
.C(n_223),
.Y(n_304)
);

NAND2xp5_ASAP7_75t_SL g225 ( 
.A(n_226),
.B(n_302),
.Y(n_225)
);

OAI21xp5_ASAP7_75t_L g226 ( 
.A1(n_227),
.A2(n_246),
.B(n_301),
.Y(n_226)
);

NOR2xp33_ASAP7_75t_L g227 ( 
.A(n_228),
.B(n_243),
.Y(n_227)
);

NAND2xp5_ASAP7_75t_SL g301 ( 
.A(n_228),
.B(n_243),
.Y(n_301)
);

MAJIxp5_ASAP7_75t_L g228 ( 
.A(n_229),
.B(n_231),
.C(n_234),
.Y(n_228)
);

XOR2xp5_ASAP7_75t_L g297 ( 
.A(n_229),
.B(n_298),
.Y(n_297)
);

OAI22xp5_ASAP7_75t_L g298 ( 
.A1(n_231),
.A2(n_234),
.B1(n_235),
.B2(n_299),
.Y(n_298)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_231),
.Y(n_299)
);

INVxp67_ASAP7_75t_L g232 ( 
.A(n_233),
.Y(n_232)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_235),
.Y(n_234)
);

NOR2xp33_ASAP7_75t_L g235 ( 
.A(n_236),
.B(n_241),
.Y(n_235)
);

OAI22xp5_ASAP7_75t_SL g292 ( 
.A1(n_236),
.A2(n_237),
.B1(n_241),
.B2(n_293),
.Y(n_292)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_237),
.Y(n_236)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_239),
.Y(n_238)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_241),
.Y(n_293)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_244),
.Y(n_245)
);

AOI21xp5_ASAP7_75t_L g246 ( 
.A1(n_247),
.A2(n_295),
.B(n_300),
.Y(n_246)
);

OAI21xp5_ASAP7_75t_SL g247 ( 
.A1(n_248),
.A2(n_284),
.B(n_294),
.Y(n_247)
);

AOI21xp5_ASAP7_75t_L g248 ( 
.A1(n_249),
.A2(n_264),
.B(n_283),
.Y(n_248)
);

NAND2xp5_ASAP7_75t_L g249 ( 
.A(n_250),
.B(n_257),
.Y(n_249)
);

NOR2xp33_ASAP7_75t_SL g283 ( 
.A(n_250),
.B(n_257),
.Y(n_283)
);

NAND2xp5_ASAP7_75t_SL g250 ( 
.A(n_251),
.B(n_255),
.Y(n_250)
);

OAI22xp5_ASAP7_75t_SL g270 ( 
.A1(n_251),
.A2(n_252),
.B1(n_255),
.B2(n_271),
.Y(n_270)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_252),
.Y(n_251)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_255),
.Y(n_271)
);

XNOR2xp5_ASAP7_75t_L g257 ( 
.A(n_258),
.B(n_262),
.Y(n_257)
);

XNOR2xp5_ASAP7_75t_L g258 ( 
.A(n_259),
.B(n_260),
.Y(n_258)
);

MAJIxp5_ASAP7_75t_L g285 ( 
.A(n_259),
.B(n_260),
.C(n_262),
.Y(n_285)
);

INVxp67_ASAP7_75t_L g291 ( 
.A(n_261),
.Y(n_291)
);

CKINVDCx14_ASAP7_75t_R g269 ( 
.A(n_263),
.Y(n_269)
);

OAI21xp5_ASAP7_75t_SL g264 ( 
.A1(n_265),
.A2(n_272),
.B(n_282),
.Y(n_264)
);

NOR2xp33_ASAP7_75t_L g265 ( 
.A(n_266),
.B(n_270),
.Y(n_265)
);

NAND2xp5_ASAP7_75t_SL g282 ( 
.A(n_266),
.B(n_270),
.Y(n_282)
);

INVxp67_ASAP7_75t_L g267 ( 
.A(n_268),
.Y(n_267)
);

AOI21xp5_ASAP7_75t_L g272 ( 
.A1(n_273),
.A2(n_278),
.B(n_281),
.Y(n_272)
);

NOR2xp33_ASAP7_75t_SL g273 ( 
.A(n_274),
.B(n_276),
.Y(n_273)
);

NAND2xp5_ASAP7_75t_L g278 ( 
.A(n_279),
.B(n_280),
.Y(n_278)
);

NOR2xp33_ASAP7_75t_SL g281 ( 
.A(n_279),
.B(n_280),
.Y(n_281)
);

NOR2xp33_ASAP7_75t_L g284 ( 
.A(n_285),
.B(n_286),
.Y(n_284)
);

NAND2xp5_ASAP7_75t_SL g294 ( 
.A(n_285),
.B(n_286),
.Y(n_294)
);

XNOR2xp5_ASAP7_75t_L g286 ( 
.A(n_287),
.B(n_292),
.Y(n_286)
);

XNOR2xp5_ASAP7_75t_L g287 ( 
.A(n_288),
.B(n_290),
.Y(n_287)
);

MAJIxp5_ASAP7_75t_L g296 ( 
.A(n_288),
.B(n_290),
.C(n_292),
.Y(n_296)
);

NAND2xp5_ASAP7_75t_L g295 ( 
.A(n_296),
.B(n_297),
.Y(n_295)
);

NOR2xp33_ASAP7_75t_SL g300 ( 
.A(n_296),
.B(n_297),
.Y(n_300)
);

NOR2xp33_ASAP7_75t_L g303 ( 
.A(n_304),
.B(n_305),
.Y(n_303)
);

NAND2xp5_ASAP7_75t_L g308 ( 
.A(n_304),
.B(n_305),
.Y(n_308)
);

NAND2xp5_ASAP7_75t_SL g314 ( 
.A(n_315),
.B(n_316),
.Y(n_314)
);

NOR2xp33_ASAP7_75t_L g326 ( 
.A(n_315),
.B(n_316),
.Y(n_326)
);

XNOR2xp5_ASAP7_75t_L g316 ( 
.A(n_317),
.B(n_325),
.Y(n_316)
);

AOI22xp5_ASAP7_75t_L g317 ( 
.A1(n_318),
.A2(n_320),
.B1(n_323),
.B2(n_324),
.Y(n_317)
);

CKINVDCx20_ASAP7_75t_R g323 ( 
.A(n_318),
.Y(n_323)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_320),
.Y(n_324)
);

MAJIxp5_ASAP7_75t_L g330 ( 
.A(n_320),
.B(n_323),
.C(n_325),
.Y(n_330)
);

NOR2xp33_ASAP7_75t_L g327 ( 
.A(n_328),
.B(n_330),
.Y(n_327)
);

CKINVDCx20_ASAP7_75t_R g333 ( 
.A(n_328),
.Y(n_333)
);

NAND2xp5_ASAP7_75t_L g335 ( 
.A(n_328),
.B(n_336),
.Y(n_335)
);

CKINVDCx14_ASAP7_75t_R g334 ( 
.A(n_330),
.Y(n_334)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_332),
.Y(n_331)
);

NOR2xp33_ASAP7_75t_L g332 ( 
.A(n_333),
.B(n_334),
.Y(n_332)
);

NAND2xp5_ASAP7_75t_L g339 ( 
.A(n_333),
.B(n_337),
.Y(n_339)
);

CKINVDCx20_ASAP7_75t_R g336 ( 
.A(n_337),
.Y(n_336)
);

CKINVDCx20_ASAP7_75t_R g338 ( 
.A(n_339),
.Y(n_338)
);


endmodule