module fake_jpeg_12758_n_627 (n_13, n_1, n_10, n_6, n_14, n_18, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_627);

input n_13;
input n_1;
input n_10;
input n_6;
input n_14;
input n_18;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_627;

wire n_529;
wire n_595;
wire n_390;
wire n_552;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_252;
wire n_19;
wire n_182;
wire n_525;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_586;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_620;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_611;
wire n_44;
wire n_355;
wire n_519;
wire n_276;
wire n_143;
wire n_431;
wire n_102;
wire n_549;
wire n_196;
wire n_66;
wire n_374;
wire n_566;
wire n_142;
wire n_417;
wire n_362;
wire n_470;
wire n_597;
wire n_172;
wire n_547;
wire n_345;
wire n_591;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_513;
wire n_283;
wire n_107;
wire n_490;
wire n_517;
wire n_415;
wire n_479;
wire n_543;
wire n_357;
wire n_89;
wire n_131;
wire n_607;
wire n_294;
wire n_230;
wire n_170;
wire n_602;
wire n_313;
wire n_542;
wire n_574;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_559;
wire n_48;
wire n_465;
wire n_200;
wire n_582;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_623;
wire n_579;
wire n_416;
wire n_221;
wire n_256;
wire n_454;
wire n_540;
wire n_292;
wire n_213;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_571;
wire n_82;
wire n_155;
wire n_508;
wire n_309;
wire n_624;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_606;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_569;
wire n_596;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_544;
wire n_31;
wire n_277;
wire n_255;
wire n_605;
wire n_601;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_393;
wire n_349;
wire n_234;
wire n_530;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_557;
wire n_408;
wire n_80;
wire n_562;
wire n_204;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_298;
wire n_106;
wire n_545;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_584;
wire n_254;
wire n_608;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_622;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_474;
wire n_539;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_626;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_575;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_511;
wire n_305;
wire n_161;
wire n_441;
wire n_555;
wire n_342;
wire n_101;
wire n_226;
wire n_509;
wire n_149;
wire n_87;
wire n_46;
wire n_578;
wire n_589;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_614;
wire n_97;
wire n_573;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_610;
wire n_174;
wire n_198;
wire n_422;
wire n_560;
wire n_190;
wire n_510;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_536;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_537;
wire n_110;
wire n_594;
wire n_590;
wire n_531;
wire n_76;
wire n_278;
wire n_343;
wire n_577;
wire n_26;
wire n_88;
wire n_397;
wire n_592;
wire n_363;
wire n_570;
wire n_238;
wire n_598;
wire n_615;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_554;
wire n_301;
wire n_609;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_523;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_533;
wire n_612;
wire n_296;
wire n_384;
wire n_588;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_585;
wire n_491;
wire n_24;
wire n_526;
wire n_467;
wire n_269;
wire n_572;
wire n_546;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_473;
wire n_45;
wire n_520;
wire n_476;
wire n_337;
wire n_317;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_344;
wire n_328;
wire n_218;
wire n_63;
wire n_599;
wire n_239;
wire n_243;
wire n_481;
wire n_619;
wire n_348;
wire n_587;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_583;
wire n_522;
wire n_333;
wire n_518;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_565;
wire n_302;
wire n_216;
wire n_528;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_199;
wire n_260;
wire n_550;
wire n_413;
wire n_275;
wire n_494;
wire n_604;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_551;
wire n_36;
wire n_62;
wire n_600;
wire n_492;
wire n_603;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_567;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_515;
wire n_347;
wire n_521;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_538;
wire n_625;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_534;
wire n_472;
wire n_279;
wire n_593;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_618;
wire n_356;
wire n_119;
wire n_484;
wire n_568;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_576;
wire n_469;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_553;
wire n_257;
wire n_61;
wire n_173;
wire n_561;
wire n_244;
wire n_232;
wire n_527;
wire n_482;
wire n_58;
wire n_41;
wire n_613;
wire n_266;
wire n_548;
wire n_72;
wire n_512;
wire n_445;
wire n_443;
wire n_617;
wire n_215;
wire n_212;
wire n_516;
wire n_183;
wire n_409;
wire n_532;
wire n_249;
wire n_412;
wire n_581;
wire n_217;
wire n_471;
wire n_580;
wire n_541;
wire n_53;
wire n_372;
wire n_558;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_535;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_556;
wire n_524;
wire n_402;
wire n_563;
wire n_504;
wire n_438;
wire n_475;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_616;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_514;
wire n_564;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_621;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

BUFx12f_ASAP7_75t_L g19 ( 
.A(n_2),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_18),
.Y(n_20)
);

BUFx5_ASAP7_75t_L g21 ( 
.A(n_1),
.Y(n_21)
);

INVx6_ASAP7_75t_L g22 ( 
.A(n_9),
.Y(n_22)
);

BUFx5_ASAP7_75t_L g23 ( 
.A(n_9),
.Y(n_23)
);

INVx4_ASAP7_75t_L g24 ( 
.A(n_14),
.Y(n_24)
);

BUFx4f_ASAP7_75t_L g25 ( 
.A(n_13),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_15),
.Y(n_26)
);

HB1xp67_ASAP7_75t_L g27 ( 
.A(n_8),
.Y(n_27)
);

BUFx12_ASAP7_75t_L g28 ( 
.A(n_12),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_10),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_0),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_18),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_4),
.Y(n_32)
);

INVx2_ASAP7_75t_L g33 ( 
.A(n_0),
.Y(n_33)
);

INVx8_ASAP7_75t_L g34 ( 
.A(n_2),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_0),
.Y(n_35)
);

INVx2_ASAP7_75t_L g36 ( 
.A(n_14),
.Y(n_36)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_1),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_11),
.Y(n_38)
);

INVx8_ASAP7_75t_L g39 ( 
.A(n_7),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_7),
.Y(n_40)
);

INVx5_ASAP7_75t_L g41 ( 
.A(n_3),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_0),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_9),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_2),
.Y(n_44)
);

BUFx12f_ASAP7_75t_L g45 ( 
.A(n_2),
.Y(n_45)
);

INVx3_ASAP7_75t_L g46 ( 
.A(n_18),
.Y(n_46)
);

INVx8_ASAP7_75t_L g47 ( 
.A(n_14),
.Y(n_47)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_8),
.Y(n_48)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_1),
.Y(n_49)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_7),
.Y(n_50)
);

INVx6_ASAP7_75t_L g51 ( 
.A(n_13),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_17),
.Y(n_52)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_13),
.Y(n_53)
);

INVx2_ASAP7_75t_L g54 ( 
.A(n_14),
.Y(n_54)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_11),
.Y(n_55)
);

CKINVDCx20_ASAP7_75t_R g56 ( 
.A(n_0),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_2),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_1),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_SL g59 ( 
.A(n_27),
.B(n_10),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_L g130 ( 
.A(n_59),
.B(n_108),
.Y(n_130)
);

INVx4_ASAP7_75t_L g60 ( 
.A(n_19),
.Y(n_60)
);

INVx3_ASAP7_75t_L g135 ( 
.A(n_60),
.Y(n_135)
);

INVx2_ASAP7_75t_SL g61 ( 
.A(n_19),
.Y(n_61)
);

BUFx3_ASAP7_75t_L g150 ( 
.A(n_61),
.Y(n_150)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_30),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g149 ( 
.A(n_62),
.Y(n_149)
);

BUFx3_ASAP7_75t_L g63 ( 
.A(n_23),
.Y(n_63)
);

BUFx12f_ASAP7_75t_L g177 ( 
.A(n_63),
.Y(n_177)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_20),
.Y(n_64)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_64),
.Y(n_172)
);

INVx11_ASAP7_75t_L g65 ( 
.A(n_21),
.Y(n_65)
);

INVx11_ASAP7_75t_L g154 ( 
.A(n_65),
.Y(n_154)
);

INVx4_ASAP7_75t_L g66 ( 
.A(n_19),
.Y(n_66)
);

INVx3_ASAP7_75t_L g137 ( 
.A(n_66),
.Y(n_137)
);

INVx5_ASAP7_75t_L g67 ( 
.A(n_24),
.Y(n_67)
);

BUFx2_ASAP7_75t_L g140 ( 
.A(n_67),
.Y(n_140)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_20),
.Y(n_68)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_68),
.Y(n_185)
);

INVx2_ASAP7_75t_L g69 ( 
.A(n_33),
.Y(n_69)
);

INVx2_ASAP7_75t_L g134 ( 
.A(n_69),
.Y(n_134)
);

INVx3_ASAP7_75t_L g70 ( 
.A(n_24),
.Y(n_70)
);

INVx3_ASAP7_75t_L g156 ( 
.A(n_70),
.Y(n_156)
);

INVx2_ASAP7_75t_L g71 ( 
.A(n_33),
.Y(n_71)
);

INVx2_ASAP7_75t_L g139 ( 
.A(n_71),
.Y(n_139)
);

INVx8_ASAP7_75t_L g72 ( 
.A(n_23),
.Y(n_72)
);

INVx5_ASAP7_75t_L g209 ( 
.A(n_72),
.Y(n_209)
);

INVx8_ASAP7_75t_L g73 ( 
.A(n_21),
.Y(n_73)
);

BUFx6f_ASAP7_75t_L g159 ( 
.A(n_73),
.Y(n_159)
);

INVx2_ASAP7_75t_L g74 ( 
.A(n_36),
.Y(n_74)
);

INVx2_ASAP7_75t_L g144 ( 
.A(n_74),
.Y(n_144)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_26),
.B(n_10),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_SL g169 ( 
.A(n_75),
.B(n_118),
.Y(n_169)
);

INVx3_ASAP7_75t_L g76 ( 
.A(n_19),
.Y(n_76)
);

INVx3_ASAP7_75t_L g160 ( 
.A(n_76),
.Y(n_160)
);

INVx3_ASAP7_75t_L g77 ( 
.A(n_45),
.Y(n_77)
);

INVx3_ASAP7_75t_L g162 ( 
.A(n_77),
.Y(n_162)
);

BUFx6f_ASAP7_75t_L g78 ( 
.A(n_30),
.Y(n_78)
);

BUFx6f_ASAP7_75t_L g179 ( 
.A(n_78),
.Y(n_179)
);

INVx2_ASAP7_75t_L g79 ( 
.A(n_36),
.Y(n_79)
);

INVx2_ASAP7_75t_L g145 ( 
.A(n_79),
.Y(n_145)
);

INVx3_ASAP7_75t_L g80 ( 
.A(n_45),
.Y(n_80)
);

INVx3_ASAP7_75t_L g165 ( 
.A(n_80),
.Y(n_165)
);

AOI22xp5_ASAP7_75t_L g81 ( 
.A1(n_54),
.A2(n_10),
.B1(n_17),
.B2(n_16),
.Y(n_81)
);

OAI22xp33_ASAP7_75t_SL g206 ( 
.A1(n_81),
.A2(n_12),
.B1(n_17),
.B2(n_5),
.Y(n_206)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_31),
.Y(n_82)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_82),
.Y(n_186)
);

BUFx6f_ASAP7_75t_L g83 ( 
.A(n_30),
.Y(n_83)
);

BUFx6f_ASAP7_75t_L g192 ( 
.A(n_83),
.Y(n_192)
);

INVx8_ASAP7_75t_L g84 ( 
.A(n_40),
.Y(n_84)
);

BUFx6f_ASAP7_75t_L g211 ( 
.A(n_84),
.Y(n_211)
);

INVx11_ASAP7_75t_L g85 ( 
.A(n_34),
.Y(n_85)
);

INVx5_ASAP7_75t_SL g153 ( 
.A(n_85),
.Y(n_153)
);

INVx2_ASAP7_75t_L g86 ( 
.A(n_54),
.Y(n_86)
);

INVx2_ASAP7_75t_L g148 ( 
.A(n_86),
.Y(n_148)
);

BUFx6f_ASAP7_75t_L g87 ( 
.A(n_32),
.Y(n_87)
);

BUFx6f_ASAP7_75t_L g214 ( 
.A(n_87),
.Y(n_214)
);

BUFx6f_ASAP7_75t_L g88 ( 
.A(n_32),
.Y(n_88)
);

BUFx6f_ASAP7_75t_L g217 ( 
.A(n_88),
.Y(n_217)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_31),
.Y(n_89)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_89),
.Y(n_199)
);

INVx11_ASAP7_75t_L g90 ( 
.A(n_34),
.Y(n_90)
);

INVx3_ASAP7_75t_SL g143 ( 
.A(n_90),
.Y(n_143)
);

BUFx6f_ASAP7_75t_L g91 ( 
.A(n_32),
.Y(n_91)
);

INVx6_ASAP7_75t_L g152 ( 
.A(n_91),
.Y(n_152)
);

BUFx12f_ASAP7_75t_SL g92 ( 
.A(n_41),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g155 ( 
.A(n_92),
.B(n_103),
.Y(n_155)
);

BUFx6f_ASAP7_75t_L g93 ( 
.A(n_42),
.Y(n_93)
);

INVx6_ASAP7_75t_L g163 ( 
.A(n_93),
.Y(n_163)
);

BUFx6f_ASAP7_75t_L g94 ( 
.A(n_42),
.Y(n_94)
);

INVx6_ASAP7_75t_L g191 ( 
.A(n_94),
.Y(n_191)
);

INVx2_ASAP7_75t_L g95 ( 
.A(n_25),
.Y(n_95)
);

INVx2_ASAP7_75t_L g175 ( 
.A(n_95),
.Y(n_175)
);

INVx3_ASAP7_75t_L g96 ( 
.A(n_45),
.Y(n_96)
);

INVx3_ASAP7_75t_L g166 ( 
.A(n_96),
.Y(n_166)
);

INVx2_ASAP7_75t_L g97 ( 
.A(n_25),
.Y(n_97)
);

INVx2_ASAP7_75t_L g176 ( 
.A(n_97),
.Y(n_176)
);

BUFx6f_ASAP7_75t_L g98 ( 
.A(n_42),
.Y(n_98)
);

INVx6_ASAP7_75t_L g202 ( 
.A(n_98),
.Y(n_202)
);

BUFx6f_ASAP7_75t_L g99 ( 
.A(n_44),
.Y(n_99)
);

BUFx3_ASAP7_75t_L g174 ( 
.A(n_99),
.Y(n_174)
);

INVx2_ASAP7_75t_L g100 ( 
.A(n_25),
.Y(n_100)
);

INVx2_ASAP7_75t_L g178 ( 
.A(n_100),
.Y(n_178)
);

BUFx6f_ASAP7_75t_L g101 ( 
.A(n_44),
.Y(n_101)
);

BUFx3_ASAP7_75t_L g193 ( 
.A(n_101),
.Y(n_193)
);

BUFx6f_ASAP7_75t_L g102 ( 
.A(n_44),
.Y(n_102)
);

INVx4_ASAP7_75t_L g151 ( 
.A(n_102),
.Y(n_151)
);

CKINVDCx20_ASAP7_75t_R g103 ( 
.A(n_28),
.Y(n_103)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_48),
.Y(n_104)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_104),
.Y(n_216)
);

BUFx6f_ASAP7_75t_L g105 ( 
.A(n_57),
.Y(n_105)
);

INVx4_ASAP7_75t_L g182 ( 
.A(n_105),
.Y(n_182)
);

BUFx12f_ASAP7_75t_L g106 ( 
.A(n_40),
.Y(n_106)
);

INVx4_ASAP7_75t_L g138 ( 
.A(n_106),
.Y(n_138)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_48),
.Y(n_107)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_107),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_L g108 ( 
.A(n_26),
.B(n_18),
.Y(n_108)
);

INVx2_ASAP7_75t_L g109 ( 
.A(n_25),
.Y(n_109)
);

INVx2_ASAP7_75t_L g201 ( 
.A(n_109),
.Y(n_201)
);

INVx2_ASAP7_75t_L g110 ( 
.A(n_46),
.Y(n_110)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_110),
.Y(n_222)
);

INVx2_ASAP7_75t_L g111 ( 
.A(n_46),
.Y(n_111)
);

HB1xp67_ASAP7_75t_L g195 ( 
.A(n_111),
.Y(n_195)
);

BUFx3_ASAP7_75t_L g112 ( 
.A(n_45),
.Y(n_112)
);

INVx4_ASAP7_75t_L g142 ( 
.A(n_112),
.Y(n_142)
);

INVx11_ASAP7_75t_L g113 ( 
.A(n_34),
.Y(n_113)
);

INVxp67_ASAP7_75t_L g132 ( 
.A(n_113),
.Y(n_132)
);

BUFx2_ASAP7_75t_L g114 ( 
.A(n_39),
.Y(n_114)
);

INVx4_ASAP7_75t_L g146 ( 
.A(n_114),
.Y(n_146)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_50),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_L g157 ( 
.A(n_115),
.B(n_53),
.Y(n_157)
);

BUFx6f_ASAP7_75t_L g116 ( 
.A(n_57),
.Y(n_116)
);

INVx3_ASAP7_75t_L g184 ( 
.A(n_116),
.Y(n_184)
);

BUFx6f_ASAP7_75t_L g117 ( 
.A(n_57),
.Y(n_117)
);

INVx3_ASAP7_75t_L g188 ( 
.A(n_117),
.Y(n_188)
);

NOR2xp33_ASAP7_75t_L g118 ( 
.A(n_29),
.B(n_9),
.Y(n_118)
);

BUFx6f_ASAP7_75t_L g119 ( 
.A(n_58),
.Y(n_119)
);

INVx3_ASAP7_75t_L g189 ( 
.A(n_119),
.Y(n_189)
);

BUFx5_ASAP7_75t_L g120 ( 
.A(n_40),
.Y(n_120)
);

INVx4_ASAP7_75t_L g161 ( 
.A(n_120),
.Y(n_161)
);

BUFx6f_ASAP7_75t_L g121 ( 
.A(n_58),
.Y(n_121)
);

INVx3_ASAP7_75t_L g194 ( 
.A(n_121),
.Y(n_194)
);

INVx4_ASAP7_75t_L g122 ( 
.A(n_41),
.Y(n_122)
);

INVx3_ASAP7_75t_L g198 ( 
.A(n_122),
.Y(n_198)
);

BUFx6f_ASAP7_75t_L g123 ( 
.A(n_58),
.Y(n_123)
);

INVx3_ASAP7_75t_L g213 ( 
.A(n_123),
.Y(n_213)
);

BUFx3_ASAP7_75t_L g124 ( 
.A(n_43),
.Y(n_124)
);

INVx4_ASAP7_75t_L g168 ( 
.A(n_124),
.Y(n_168)
);

INVx2_ASAP7_75t_L g125 ( 
.A(n_50),
.Y(n_125)
);

HB1xp67_ASAP7_75t_L g200 ( 
.A(n_125),
.Y(n_200)
);

BUFx3_ASAP7_75t_L g126 ( 
.A(n_43),
.Y(n_126)
);

INVx4_ASAP7_75t_L g204 ( 
.A(n_126),
.Y(n_204)
);

INVx3_ASAP7_75t_L g127 ( 
.A(n_39),
.Y(n_127)
);

INVx4_ASAP7_75t_L g207 ( 
.A(n_127),
.Y(n_207)
);

INVx11_ASAP7_75t_L g128 ( 
.A(n_39),
.Y(n_128)
);

INVx4_ASAP7_75t_L g212 ( 
.A(n_128),
.Y(n_212)
);

NOR2xp33_ASAP7_75t_L g129 ( 
.A(n_29),
.B(n_8),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_SL g197 ( 
.A(n_129),
.B(n_11),
.Y(n_197)
);

AOI22xp5_ASAP7_75t_L g131 ( 
.A1(n_62),
.A2(n_22),
.B1(n_51),
.B2(n_52),
.Y(n_131)
);

OA22x2_ASAP7_75t_L g228 ( 
.A1(n_131),
.A2(n_164),
.B1(n_196),
.B2(n_206),
.Y(n_228)
);

NAND2xp5_ASAP7_75t_L g133 ( 
.A(n_61),
.B(n_38),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_L g253 ( 
.A(n_133),
.B(n_147),
.Y(n_253)
);

AOI22xp33_ASAP7_75t_SL g136 ( 
.A1(n_72),
.A2(n_47),
.B1(n_22),
.B2(n_51),
.Y(n_136)
);

AOI21xp5_ASAP7_75t_L g275 ( 
.A1(n_136),
.A2(n_141),
.B(n_173),
.Y(n_275)
);

AOI22xp33_ASAP7_75t_SL g141 ( 
.A1(n_73),
.A2(n_47),
.B1(n_51),
.B2(n_52),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_L g147 ( 
.A(n_60),
.B(n_38),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_L g262 ( 
.A(n_157),
.B(n_181),
.Y(n_262)
);

AND2x2_ASAP7_75t_L g158 ( 
.A(n_66),
.B(n_55),
.Y(n_158)
);

CKINVDCx14_ASAP7_75t_R g281 ( 
.A(n_158),
.Y(n_281)
);

AOI22xp5_ASAP7_75t_L g164 ( 
.A1(n_78),
.A2(n_52),
.B1(n_43),
.B2(n_47),
.Y(n_164)
);

NOR2xp33_ASAP7_75t_SL g167 ( 
.A(n_112),
.B(n_56),
.Y(n_167)
);

NOR2xp33_ASAP7_75t_SL g227 ( 
.A(n_167),
.B(n_170),
.Y(n_227)
);

NOR2xp33_ASAP7_75t_L g170 ( 
.A(n_63),
.B(n_55),
.Y(n_170)
);

NOR2xp33_ASAP7_75t_L g171 ( 
.A(n_122),
.B(n_53),
.Y(n_171)
);

NOR2xp33_ASAP7_75t_SL g284 ( 
.A(n_171),
.B(n_180),
.Y(n_284)
);

AOI22xp33_ASAP7_75t_SL g173 ( 
.A1(n_114),
.A2(n_37),
.B1(n_49),
.B2(n_56),
.Y(n_173)
);

CKINVDCx20_ASAP7_75t_R g180 ( 
.A(n_85),
.Y(n_180)
);

OR2x2_ASAP7_75t_L g181 ( 
.A(n_65),
.B(n_37),
.Y(n_181)
);

AOI22xp33_ASAP7_75t_SL g183 ( 
.A1(n_84),
.A2(n_49),
.B1(n_35),
.B2(n_12),
.Y(n_183)
);

AOI21xp5_ASAP7_75t_L g277 ( 
.A1(n_183),
.A2(n_219),
.B(n_220),
.Y(n_277)
);

OAI21xp33_ASAP7_75t_L g187 ( 
.A1(n_90),
.A2(n_35),
.B(n_11),
.Y(n_187)
);

OAI21xp33_ASAP7_75t_L g259 ( 
.A1(n_187),
.A2(n_5),
.B(n_6),
.Y(n_259)
);

CKINVDCx20_ASAP7_75t_R g190 ( 
.A(n_113),
.Y(n_190)
);

NOR2xp33_ASAP7_75t_L g265 ( 
.A(n_190),
.B(n_205),
.Y(n_265)
);

AOI22xp33_ASAP7_75t_L g196 ( 
.A1(n_83),
.A2(n_1),
.B1(n_3),
.B2(n_4),
.Y(n_196)
);

NAND2xp5_ASAP7_75t_L g276 ( 
.A(n_197),
.B(n_203),
.Y(n_276)
);

NAND2xp5_ASAP7_75t_L g203 ( 
.A(n_87),
.B(n_12),
.Y(n_203)
);

CKINVDCx20_ASAP7_75t_R g205 ( 
.A(n_128),
.Y(n_205)
);

NOR2xp33_ASAP7_75t_L g208 ( 
.A(n_106),
.B(n_8),
.Y(n_208)
);

NAND2xp5_ASAP7_75t_SL g229 ( 
.A(n_208),
.B(n_3),
.Y(n_229)
);

INVx6_ASAP7_75t_SL g210 ( 
.A(n_106),
.Y(n_210)
);

CKINVDCx16_ASAP7_75t_R g301 ( 
.A(n_210),
.Y(n_301)
);

OR2x2_ASAP7_75t_L g215 ( 
.A(n_124),
.B(n_28),
.Y(n_215)
);

NOR2xp33_ASAP7_75t_L g266 ( 
.A(n_215),
.B(n_6),
.Y(n_266)
);

AND2x2_ASAP7_75t_L g218 ( 
.A(n_126),
.B(n_13),
.Y(n_218)
);

AND2x2_ASAP7_75t_L g224 ( 
.A(n_218),
.B(n_3),
.Y(n_224)
);

AOI22xp33_ASAP7_75t_SL g219 ( 
.A1(n_88),
.A2(n_7),
.B1(n_17),
.B2(n_5),
.Y(n_219)
);

AOI22xp33_ASAP7_75t_SL g220 ( 
.A1(n_91),
.A2(n_5),
.B1(n_6),
.B2(n_15),
.Y(n_220)
);

INVx4_ASAP7_75t_L g223 ( 
.A(n_146),
.Y(n_223)
);

INVx4_ASAP7_75t_L g342 ( 
.A(n_223),
.Y(n_342)
);

XNOR2x1_ASAP7_75t_L g311 ( 
.A(n_224),
.B(n_289),
.Y(n_311)
);

INVx6_ASAP7_75t_L g225 ( 
.A(n_149),
.Y(n_225)
);

BUFx6f_ASAP7_75t_L g357 ( 
.A(n_225),
.Y(n_357)
);

INVx3_ASAP7_75t_L g226 ( 
.A(n_150),
.Y(n_226)
);

BUFx2_ASAP7_75t_L g303 ( 
.A(n_226),
.Y(n_303)
);

NOR2xp33_ASAP7_75t_L g318 ( 
.A(n_229),
.B(n_235),
.Y(n_318)
);

INVx3_ASAP7_75t_L g230 ( 
.A(n_150),
.Y(n_230)
);

INVx3_ASAP7_75t_L g316 ( 
.A(n_230),
.Y(n_316)
);

INVx2_ASAP7_75t_SL g231 ( 
.A(n_135),
.Y(n_231)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_231),
.Y(n_313)
);

BUFx3_ASAP7_75t_L g232 ( 
.A(n_177),
.Y(n_232)
);

INVxp67_ASAP7_75t_SL g333 ( 
.A(n_232),
.Y(n_333)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_172),
.Y(n_233)
);

INVx1_ASAP7_75t_SL g302 ( 
.A(n_233),
.Y(n_302)
);

INVx2_ASAP7_75t_L g234 ( 
.A(n_175),
.Y(n_234)
);

INVx2_ASAP7_75t_L g319 ( 
.A(n_234),
.Y(n_319)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_185),
.Y(n_235)
);

AOI22xp33_ASAP7_75t_L g236 ( 
.A1(n_200),
.A2(n_98),
.B1(n_121),
.B2(n_119),
.Y(n_236)
);

OAI22xp5_ASAP7_75t_L g354 ( 
.A1(n_236),
.A2(n_292),
.B1(n_297),
.B2(n_301),
.Y(n_354)
);

BUFx3_ASAP7_75t_L g237 ( 
.A(n_177),
.Y(n_237)
);

INVx5_ASAP7_75t_L g348 ( 
.A(n_237),
.Y(n_348)
);

MAJIxp5_ASAP7_75t_L g238 ( 
.A(n_186),
.B(n_94),
.C(n_117),
.Y(n_238)
);

MAJIxp5_ASAP7_75t_L g346 ( 
.A(n_238),
.B(n_290),
.C(n_214),
.Y(n_346)
);

INVx3_ASAP7_75t_L g239 ( 
.A(n_211),
.Y(n_239)
);

INVx3_ASAP7_75t_L g358 ( 
.A(n_239),
.Y(n_358)
);

INVx2_ASAP7_75t_L g240 ( 
.A(n_176),
.Y(n_240)
);

INVx2_ASAP7_75t_L g339 ( 
.A(n_240),
.Y(n_339)
);

INVx3_ASAP7_75t_L g241 ( 
.A(n_211),
.Y(n_241)
);

INVx2_ASAP7_75t_L g351 ( 
.A(n_241),
.Y(n_351)
);

BUFx12_ASAP7_75t_L g242 ( 
.A(n_153),
.Y(n_242)
);

BUFx4f_ASAP7_75t_SL g343 ( 
.A(n_242),
.Y(n_343)
);

AO22x1_ASAP7_75t_SL g243 ( 
.A1(n_196),
.A2(n_145),
.B1(n_144),
.B2(n_148),
.Y(n_243)
);

NAND2xp5_ASAP7_75t_L g323 ( 
.A(n_243),
.B(n_299),
.Y(n_323)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_199),
.Y(n_244)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_244),
.Y(n_327)
);

CKINVDCx20_ASAP7_75t_R g245 ( 
.A(n_200),
.Y(n_245)
);

NOR2xp33_ASAP7_75t_L g305 ( 
.A(n_245),
.B(n_247),
.Y(n_305)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_216),
.Y(n_246)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_246),
.Y(n_332)
);

CKINVDCx20_ASAP7_75t_R g247 ( 
.A(n_195),
.Y(n_247)
);

NAND2xp5_ASAP7_75t_SL g248 ( 
.A(n_130),
.B(n_93),
.Y(n_248)
);

NOR2xp33_ASAP7_75t_SL g309 ( 
.A(n_248),
.B(n_279),
.Y(n_309)
);

INVx1_ASAP7_75t_SL g249 ( 
.A(n_177),
.Y(n_249)
);

AND2x2_ASAP7_75t_L g304 ( 
.A(n_249),
.B(n_251),
.Y(n_304)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_221),
.Y(n_250)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_250),
.Y(n_335)
);

AND2x4_ASAP7_75t_SL g251 ( 
.A(n_134),
.B(n_116),
.Y(n_251)
);

AOI22xp33_ASAP7_75t_SL g252 ( 
.A1(n_143),
.A2(n_123),
.B1(n_105),
.B2(n_102),
.Y(n_252)
);

INVxp67_ASAP7_75t_L g308 ( 
.A(n_252),
.Y(n_308)
);

BUFx2_ASAP7_75t_SL g254 ( 
.A(n_153),
.Y(n_254)
);

INVxp67_ASAP7_75t_L g322 ( 
.A(n_254),
.Y(n_322)
);

AOI22xp33_ASAP7_75t_SL g255 ( 
.A1(n_143),
.A2(n_101),
.B1(n_99),
.B2(n_28),
.Y(n_255)
);

AOI22xp33_ASAP7_75t_SL g349 ( 
.A1(n_255),
.A2(n_270),
.B1(n_273),
.B2(n_288),
.Y(n_349)
);

INVx2_ASAP7_75t_L g256 ( 
.A(n_178),
.Y(n_256)
);

INVx1_ASAP7_75t_L g353 ( 
.A(n_256),
.Y(n_353)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_195),
.Y(n_257)
);

NOR2xp33_ASAP7_75t_L g310 ( 
.A(n_257),
.B(n_258),
.Y(n_310)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_201),
.Y(n_258)
);

AND2x2_ASAP7_75t_L g306 ( 
.A(n_259),
.B(n_266),
.Y(n_306)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_222),
.Y(n_260)
);

NOR2xp33_ASAP7_75t_L g320 ( 
.A(n_260),
.B(n_261),
.Y(n_320)
);

CKINVDCx20_ASAP7_75t_R g261 ( 
.A(n_158),
.Y(n_261)
);

BUFx3_ASAP7_75t_L g263 ( 
.A(n_140),
.Y(n_263)
);

INVx8_ASAP7_75t_L g345 ( 
.A(n_263),
.Y(n_345)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_139),
.Y(n_264)
);

NOR2xp33_ASAP7_75t_L g324 ( 
.A(n_264),
.B(n_269),
.Y(n_324)
);

INVx1_ASAP7_75t_SL g267 ( 
.A(n_140),
.Y(n_267)
);

CKINVDCx16_ASAP7_75t_R g331 ( 
.A(n_267),
.Y(n_331)
);

NAND2xp67_ASAP7_75t_SL g268 ( 
.A(n_169),
.B(n_6),
.Y(n_268)
);

CKINVDCx14_ASAP7_75t_R g317 ( 
.A(n_268),
.Y(n_317)
);

INVx2_ASAP7_75t_L g269 ( 
.A(n_137),
.Y(n_269)
);

AOI22xp33_ASAP7_75t_SL g270 ( 
.A1(n_209),
.A2(n_28),
.B1(n_15),
.B2(n_16),
.Y(n_270)
);

INVx2_ASAP7_75t_L g271 ( 
.A(n_184),
.Y(n_271)
);

NOR2xp33_ASAP7_75t_L g325 ( 
.A(n_271),
.B(n_272),
.Y(n_325)
);

INVx2_ASAP7_75t_L g272 ( 
.A(n_188),
.Y(n_272)
);

BUFx6f_ASAP7_75t_L g273 ( 
.A(n_149),
.Y(n_273)
);

AOI22x1_ASAP7_75t_L g274 ( 
.A1(n_218),
.A2(n_187),
.B1(n_215),
.B2(n_141),
.Y(n_274)
);

AOI21xp5_ASAP7_75t_L g315 ( 
.A1(n_274),
.A2(n_132),
.B(n_182),
.Y(n_315)
);

BUFx2_ASAP7_75t_L g278 ( 
.A(n_159),
.Y(n_278)
);

CKINVDCx16_ASAP7_75t_R g341 ( 
.A(n_278),
.Y(n_341)
);

NAND2xp5_ASAP7_75t_L g279 ( 
.A(n_155),
.B(n_15),
.Y(n_279)
);

NAND2xp5_ASAP7_75t_L g280 ( 
.A(n_181),
.B(n_16),
.Y(n_280)
);

NOR2xp33_ASAP7_75t_SL g321 ( 
.A(n_280),
.B(n_291),
.Y(n_321)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_156),
.Y(n_282)
);

NOR2xp33_ASAP7_75t_L g329 ( 
.A(n_282),
.B(n_283),
.Y(n_329)
);

INVx5_ASAP7_75t_L g283 ( 
.A(n_159),
.Y(n_283)
);

INVxp67_ASAP7_75t_L g285 ( 
.A(n_173),
.Y(n_285)
);

NOR2xp33_ASAP7_75t_L g334 ( 
.A(n_285),
.B(n_287),
.Y(n_334)
);

INVx3_ASAP7_75t_L g286 ( 
.A(n_168),
.Y(n_286)
);

CKINVDCx20_ASAP7_75t_R g340 ( 
.A(n_286),
.Y(n_340)
);

INVx3_ASAP7_75t_L g287 ( 
.A(n_204),
.Y(n_287)
);

INVx1_ASAP7_75t_SL g288 ( 
.A(n_160),
.Y(n_288)
);

AND2x2_ASAP7_75t_L g289 ( 
.A(n_198),
.B(n_3),
.Y(n_289)
);

AND2x2_ASAP7_75t_L g290 ( 
.A(n_207),
.B(n_4),
.Y(n_290)
);

NOR2xp33_ASAP7_75t_L g291 ( 
.A(n_162),
.B(n_16),
.Y(n_291)
);

AOI22xp33_ASAP7_75t_L g292 ( 
.A1(n_189),
.A2(n_4),
.B1(n_194),
.B2(n_213),
.Y(n_292)
);

AOI22xp33_ASAP7_75t_SL g293 ( 
.A1(n_142),
.A2(n_4),
.B1(n_166),
.B2(n_165),
.Y(n_293)
);

AOI22xp33_ASAP7_75t_SL g352 ( 
.A1(n_293),
.A2(n_295),
.B1(n_296),
.B2(n_298),
.Y(n_352)
);

NOR2xp33_ASAP7_75t_L g294 ( 
.A(n_138),
.B(n_161),
.Y(n_294)
);

BUFx24_ASAP7_75t_SL g326 ( 
.A(n_294),
.Y(n_326)
);

INVx2_ASAP7_75t_L g295 ( 
.A(n_151),
.Y(n_295)
);

INVx2_ASAP7_75t_L g296 ( 
.A(n_151),
.Y(n_296)
);

AOI22xp33_ASAP7_75t_L g297 ( 
.A1(n_182),
.A2(n_202),
.B1(n_152),
.B2(n_191),
.Y(n_297)
);

BUFx3_ASAP7_75t_L g298 ( 
.A(n_174),
.Y(n_298)
);

INVx11_ASAP7_75t_L g299 ( 
.A(n_154),
.Y(n_299)
);

INVx3_ASAP7_75t_L g300 ( 
.A(n_174),
.Y(n_300)
);

NAND2xp5_ASAP7_75t_L g355 ( 
.A(n_300),
.B(n_267),
.Y(n_355)
);

OAI21xp5_ASAP7_75t_L g307 ( 
.A1(n_285),
.A2(n_183),
.B(n_219),
.Y(n_307)
);

OAI21xp5_ASAP7_75t_L g362 ( 
.A1(n_307),
.A2(n_337),
.B(n_344),
.Y(n_362)
);

XOR2xp5_ASAP7_75t_L g312 ( 
.A(n_253),
.B(n_206),
.Y(n_312)
);

AND2x2_ASAP7_75t_L g376 ( 
.A(n_312),
.B(n_315),
.Y(n_376)
);

OAI22xp5_ASAP7_75t_SL g314 ( 
.A1(n_275),
.A2(n_136),
.B1(n_220),
.B2(n_152),
.Y(n_314)
);

AOI22xp5_ASAP7_75t_L g365 ( 
.A1(n_314),
.A2(n_336),
.B1(n_308),
.B2(n_307),
.Y(n_365)
);

AOI22xp5_ASAP7_75t_L g328 ( 
.A1(n_228),
.A2(n_163),
.B1(n_191),
.B2(n_202),
.Y(n_328)
);

OAI22xp5_ASAP7_75t_SL g361 ( 
.A1(n_328),
.A2(n_330),
.B1(n_308),
.B2(n_323),
.Y(n_361)
);

AOI22xp5_ASAP7_75t_L g330 ( 
.A1(n_228),
.A2(n_163),
.B1(n_217),
.B2(n_179),
.Y(n_330)
);

OAI22xp5_ASAP7_75t_SL g336 ( 
.A1(n_275),
.A2(n_179),
.B1(n_192),
.B2(n_214),
.Y(n_336)
);

OAI21xp5_ASAP7_75t_SL g337 ( 
.A1(n_277),
.A2(n_281),
.B(n_274),
.Y(n_337)
);

XNOR2xp5_ASAP7_75t_SL g338 ( 
.A(n_276),
.B(n_132),
.Y(n_338)
);

NAND2xp5_ASAP7_75t_SL g381 ( 
.A(n_338),
.B(n_288),
.Y(n_381)
);

OAI21xp5_ASAP7_75t_L g344 ( 
.A1(n_262),
.A2(n_193),
.B(n_192),
.Y(n_344)
);

AND2x2_ASAP7_75t_L g383 ( 
.A(n_346),
.B(n_347),
.Y(n_383)
);

MAJIxp5_ASAP7_75t_L g347 ( 
.A(n_238),
.B(n_217),
.C(n_212),
.Y(n_347)
);

AOI21xp5_ASAP7_75t_L g350 ( 
.A1(n_277),
.A2(n_193),
.B(n_265),
.Y(n_350)
);

INVxp67_ASAP7_75t_L g396 ( 
.A(n_350),
.Y(n_396)
);

AND2x2_ASAP7_75t_L g406 ( 
.A(n_354),
.B(n_360),
.Y(n_406)
);

INVx1_ASAP7_75t_L g369 ( 
.A(n_355),
.Y(n_369)
);

NAND2xp5_ASAP7_75t_L g356 ( 
.A(n_224),
.B(n_290),
.Y(n_356)
);

NAND2xp5_ASAP7_75t_L g366 ( 
.A(n_356),
.B(n_359),
.Y(n_366)
);

NAND2xp5_ASAP7_75t_L g359 ( 
.A(n_224),
.B(n_290),
.Y(n_359)
);

MAJIxp5_ASAP7_75t_L g360 ( 
.A(n_251),
.B(n_256),
.C(n_234),
.Y(n_360)
);

AOI22xp33_ASAP7_75t_L g443 ( 
.A1(n_361),
.A2(n_341),
.B1(n_316),
.B2(n_342),
.Y(n_443)
);

NOR2xp33_ASAP7_75t_L g363 ( 
.A(n_309),
.B(n_284),
.Y(n_363)
);

NOR2xp33_ASAP7_75t_SL g427 ( 
.A(n_363),
.B(n_375),
.Y(n_427)
);

OAI22xp5_ASAP7_75t_SL g364 ( 
.A1(n_330),
.A2(n_328),
.B1(n_315),
.B2(n_323),
.Y(n_364)
);

AOI22xp5_ASAP7_75t_L g423 ( 
.A1(n_364),
.A2(n_374),
.B1(n_382),
.B2(n_322),
.Y(n_423)
);

OAI22xp5_ASAP7_75t_L g442 ( 
.A1(n_365),
.A2(n_368),
.B1(n_371),
.B2(n_395),
.Y(n_442)
);

CKINVDCx20_ASAP7_75t_R g367 ( 
.A(n_305),
.Y(n_367)
);

NOR2xp33_ASAP7_75t_L g414 ( 
.A(n_367),
.B(n_377),
.Y(n_414)
);

AOI22xp5_ASAP7_75t_L g368 ( 
.A1(n_314),
.A2(n_228),
.B1(n_243),
.B2(n_259),
.Y(n_368)
);

NAND2xp5_ASAP7_75t_L g370 ( 
.A(n_346),
.B(n_312),
.Y(n_370)
);

NAND2xp5_ASAP7_75t_L g411 ( 
.A(n_370),
.B(n_373),
.Y(n_411)
);

AOI22xp5_ASAP7_75t_L g371 ( 
.A1(n_336),
.A2(n_228),
.B1(n_243),
.B2(n_251),
.Y(n_371)
);

INVx2_ASAP7_75t_L g372 ( 
.A(n_351),
.Y(n_372)
);

INVx2_ASAP7_75t_L g433 ( 
.A(n_372),
.Y(n_433)
);

A2O1A1Ixp33_ASAP7_75t_L g373 ( 
.A1(n_337),
.A2(n_268),
.B(n_289),
.C(n_227),
.Y(n_373)
);

OAI22xp5_ASAP7_75t_SL g374 ( 
.A1(n_350),
.A2(n_241),
.B1(n_239),
.B2(n_272),
.Y(n_374)
);

NOR2xp33_ASAP7_75t_SL g375 ( 
.A(n_318),
.B(n_289),
.Y(n_375)
);

CKINVDCx20_ASAP7_75t_R g377 ( 
.A(n_310),
.Y(n_377)
);

NAND2xp5_ASAP7_75t_L g378 ( 
.A(n_338),
.B(n_240),
.Y(n_378)
);

NAND2xp5_ASAP7_75t_SL g410 ( 
.A(n_378),
.B(n_384),
.Y(n_410)
);

INVx1_ASAP7_75t_L g379 ( 
.A(n_313),
.Y(n_379)
);

INVx1_ASAP7_75t_L g409 ( 
.A(n_379),
.Y(n_409)
);

INVx2_ASAP7_75t_L g380 ( 
.A(n_351),
.Y(n_380)
);

INVx1_ASAP7_75t_L g424 ( 
.A(n_380),
.Y(n_424)
);

XNOR2xp5_ASAP7_75t_L g441 ( 
.A(n_381),
.B(n_393),
.Y(n_441)
);

OAI22xp5_ASAP7_75t_SL g382 ( 
.A1(n_347),
.A2(n_271),
.B1(n_225),
.B2(n_278),
.Y(n_382)
);

NOR2xp33_ASAP7_75t_L g384 ( 
.A(n_309),
.B(n_269),
.Y(n_384)
);

NOR2xp33_ASAP7_75t_L g385 ( 
.A(n_320),
.B(n_231),
.Y(n_385)
);

NAND2xp5_ASAP7_75t_SL g426 ( 
.A(n_385),
.B(n_389),
.Y(n_426)
);

NOR2x1p5_ASAP7_75t_L g386 ( 
.A(n_304),
.B(n_242),
.Y(n_386)
);

CKINVDCx14_ASAP7_75t_R g420 ( 
.A(n_386),
.Y(n_420)
);

AO22x1_ASAP7_75t_SL g387 ( 
.A1(n_304),
.A2(n_296),
.B1(n_295),
.B2(n_299),
.Y(n_387)
);

INVx1_ASAP7_75t_L g434 ( 
.A(n_387),
.Y(n_434)
);

BUFx24_ASAP7_75t_SL g388 ( 
.A(n_326),
.Y(n_388)
);

INVxp67_ASAP7_75t_L g408 ( 
.A(n_388),
.Y(n_408)
);

NAND2xp5_ASAP7_75t_SL g389 ( 
.A(n_356),
.B(n_359),
.Y(n_389)
);

HB1xp67_ASAP7_75t_L g390 ( 
.A(n_358),
.Y(n_390)
);

CKINVDCx20_ASAP7_75t_R g416 ( 
.A(n_390),
.Y(n_416)
);

NOR2xp33_ASAP7_75t_L g391 ( 
.A(n_321),
.B(n_302),
.Y(n_391)
);

NOR2xp33_ASAP7_75t_L g430 ( 
.A(n_391),
.B(n_398),
.Y(n_430)
);

HB1xp67_ASAP7_75t_L g392 ( 
.A(n_358),
.Y(n_392)
);

CKINVDCx20_ASAP7_75t_R g431 ( 
.A(n_392),
.Y(n_431)
);

NAND2xp5_ASAP7_75t_L g393 ( 
.A(n_318),
.B(n_360),
.Y(n_393)
);

INVx2_ASAP7_75t_L g394 ( 
.A(n_319),
.Y(n_394)
);

INVx1_ASAP7_75t_L g435 ( 
.A(n_394),
.Y(n_435)
);

AOI22xp5_ASAP7_75t_L g395 ( 
.A1(n_354),
.A2(n_283),
.B1(n_273),
.B2(n_300),
.Y(n_395)
);

INVx1_ASAP7_75t_L g397 ( 
.A(n_313),
.Y(n_397)
);

INVx1_ASAP7_75t_L g438 ( 
.A(n_397),
.Y(n_438)
);

CKINVDCx20_ASAP7_75t_R g398 ( 
.A(n_329),
.Y(n_398)
);

INVx13_ASAP7_75t_L g399 ( 
.A(n_343),
.Y(n_399)
);

INVx3_ASAP7_75t_SL g425 ( 
.A(n_399),
.Y(n_425)
);

NAND2xp5_ASAP7_75t_L g400 ( 
.A(n_344),
.B(n_287),
.Y(n_400)
);

XOR2xp5_ASAP7_75t_L g417 ( 
.A(n_400),
.B(n_376),
.Y(n_417)
);

NOR2xp33_ASAP7_75t_SL g401 ( 
.A(n_321),
.B(n_286),
.Y(n_401)
);

CKINVDCx16_ASAP7_75t_R g412 ( 
.A(n_401),
.Y(n_412)
);

INVxp67_ASAP7_75t_L g402 ( 
.A(n_324),
.Y(n_402)
);

CKINVDCx20_ASAP7_75t_R g432 ( 
.A(n_402),
.Y(n_432)
);

NOR2xp33_ASAP7_75t_L g403 ( 
.A(n_302),
.B(n_223),
.Y(n_403)
);

OAI21xp5_ASAP7_75t_L g429 ( 
.A1(n_403),
.A2(n_404),
.B(n_303),
.Y(n_429)
);

NOR2xp33_ASAP7_75t_L g404 ( 
.A(n_327),
.B(n_263),
.Y(n_404)
);

INVx1_ASAP7_75t_L g405 ( 
.A(n_355),
.Y(n_405)
);

CKINVDCx20_ASAP7_75t_R g444 ( 
.A(n_405),
.Y(n_444)
);

OAI22xp5_ASAP7_75t_SL g407 ( 
.A1(n_368),
.A2(n_334),
.B1(n_349),
.B2(n_352),
.Y(n_407)
);

AOI22xp5_ASAP7_75t_L g455 ( 
.A1(n_407),
.A2(n_415),
.B1(n_421),
.B2(n_436),
.Y(n_455)
);

OAI32xp33_ASAP7_75t_L g413 ( 
.A1(n_378),
.A2(n_317),
.A3(n_325),
.B1(n_332),
.B2(n_327),
.Y(n_413)
);

NAND2xp5_ASAP7_75t_L g456 ( 
.A(n_413),
.B(n_428),
.Y(n_456)
);

OAI22xp5_ASAP7_75t_SL g415 ( 
.A1(n_365),
.A2(n_304),
.B1(n_311),
.B2(n_335),
.Y(n_415)
);

XOR2xp5_ASAP7_75t_L g462 ( 
.A(n_417),
.B(n_406),
.Y(n_462)
);

AOI32xp33_ASAP7_75t_L g418 ( 
.A1(n_362),
.A2(n_306),
.A3(n_311),
.B1(n_340),
.B2(n_322),
.Y(n_418)
);

OAI21xp5_ASAP7_75t_SL g451 ( 
.A1(n_418),
.A2(n_422),
.B(n_381),
.Y(n_451)
);

XOR2xp5_ASAP7_75t_L g419 ( 
.A(n_370),
.B(n_306),
.Y(n_419)
);

MAJIxp5_ASAP7_75t_L g447 ( 
.A(n_419),
.B(n_383),
.C(n_393),
.Y(n_447)
);

OAI22xp5_ASAP7_75t_SL g421 ( 
.A1(n_371),
.A2(n_335),
.B1(n_332),
.B2(n_306),
.Y(n_421)
);

XOR2xp5_ASAP7_75t_SL g422 ( 
.A(n_376),
.B(n_343),
.Y(n_422)
);

OAI22xp5_ASAP7_75t_L g466 ( 
.A1(n_423),
.A2(n_443),
.B1(n_403),
.B2(n_404),
.Y(n_466)
);

OAI32xp33_ASAP7_75t_L g428 ( 
.A1(n_366),
.A2(n_353),
.A3(n_319),
.B1(n_339),
.B2(n_303),
.Y(n_428)
);

NAND2xp5_ASAP7_75t_L g465 ( 
.A(n_429),
.B(n_387),
.Y(n_465)
);

OAI22xp5_ASAP7_75t_SL g436 ( 
.A1(n_362),
.A2(n_357),
.B1(n_340),
.B2(n_331),
.Y(n_436)
);

AOI21xp5_ASAP7_75t_L g437 ( 
.A1(n_396),
.A2(n_348),
.B(n_303),
.Y(n_437)
);

AOI21xp5_ASAP7_75t_L g453 ( 
.A1(n_437),
.A2(n_400),
.B(n_387),
.Y(n_453)
);

OAI22xp5_ASAP7_75t_SL g439 ( 
.A1(n_369),
.A2(n_357),
.B1(n_331),
.B2(n_353),
.Y(n_439)
);

AOI22xp5_ASAP7_75t_L g458 ( 
.A1(n_439),
.A2(n_440),
.B1(n_361),
.B2(n_397),
.Y(n_458)
);

OAI22xp5_ASAP7_75t_SL g440 ( 
.A1(n_369),
.A2(n_357),
.B1(n_341),
.B2(n_339),
.Y(n_440)
);

INVx1_ASAP7_75t_L g445 ( 
.A(n_409),
.Y(n_445)
);

INVx1_ASAP7_75t_L g491 ( 
.A(n_445),
.Y(n_491)
);

INVx1_ASAP7_75t_L g446 ( 
.A(n_409),
.Y(n_446)
);

INVx1_ASAP7_75t_L g511 ( 
.A(n_446),
.Y(n_511)
);

MAJIxp5_ASAP7_75t_L g482 ( 
.A(n_447),
.B(n_449),
.C(n_454),
.Y(n_482)
);

INVx1_ASAP7_75t_L g448 ( 
.A(n_438),
.Y(n_448)
);

INVx1_ASAP7_75t_L g503 ( 
.A(n_448),
.Y(n_503)
);

XNOR2xp5_ASAP7_75t_L g449 ( 
.A(n_441),
.B(n_383),
.Y(n_449)
);

OAI22xp5_ASAP7_75t_SL g450 ( 
.A1(n_434),
.A2(n_405),
.B1(n_376),
.B2(n_364),
.Y(n_450)
);

AOI22xp5_ASAP7_75t_L g493 ( 
.A1(n_450),
.A2(n_463),
.B1(n_466),
.B2(n_469),
.Y(n_493)
);

OAI21xp5_ASAP7_75t_L g508 ( 
.A1(n_451),
.A2(n_453),
.B(n_460),
.Y(n_508)
);

NOR2xp33_ASAP7_75t_L g452 ( 
.A(n_427),
.B(n_367),
.Y(n_452)
);

NOR2xp33_ASAP7_75t_SL g485 ( 
.A(n_452),
.B(n_457),
.Y(n_485)
);

MAJIxp5_ASAP7_75t_L g454 ( 
.A(n_419),
.B(n_383),
.C(n_366),
.Y(n_454)
);

NOR2xp33_ASAP7_75t_L g457 ( 
.A(n_427),
.B(n_377),
.Y(n_457)
);

OAI22xp5_ASAP7_75t_L g487 ( 
.A1(n_458),
.A2(n_473),
.B1(n_476),
.B2(n_432),
.Y(n_487)
);

MAJIxp5_ASAP7_75t_L g459 ( 
.A(n_441),
.B(n_417),
.C(n_422),
.Y(n_459)
);

MAJIxp5_ASAP7_75t_L g488 ( 
.A(n_459),
.B(n_461),
.C(n_462),
.Y(n_488)
);

AOI21xp5_ASAP7_75t_L g460 ( 
.A1(n_437),
.A2(n_406),
.B(n_373),
.Y(n_460)
);

XNOR2xp5_ASAP7_75t_L g461 ( 
.A(n_411),
.B(n_389),
.Y(n_461)
);

OAI22xp5_ASAP7_75t_SL g463 ( 
.A1(n_434),
.A2(n_406),
.B1(n_395),
.B2(n_384),
.Y(n_463)
);

INVx1_ASAP7_75t_L g464 ( 
.A(n_438),
.Y(n_464)
);

INVx1_ASAP7_75t_L g490 ( 
.A(n_464),
.Y(n_490)
);

CKINVDCx14_ASAP7_75t_R g496 ( 
.A(n_465),
.Y(n_496)
);

AOI21x1_ASAP7_75t_SL g467 ( 
.A1(n_411),
.A2(n_373),
.B(n_387),
.Y(n_467)
);

INVx1_ASAP7_75t_L g497 ( 
.A(n_467),
.Y(n_497)
);

AOI21xp5_ASAP7_75t_L g468 ( 
.A1(n_422),
.A2(n_399),
.B(n_398),
.Y(n_468)
);

NAND2xp5_ASAP7_75t_L g484 ( 
.A(n_468),
.B(n_471),
.Y(n_484)
);

OAI22x1_ASAP7_75t_SL g469 ( 
.A1(n_423),
.A2(n_374),
.B1(n_379),
.B2(n_401),
.Y(n_469)
);

INVx1_ASAP7_75t_L g470 ( 
.A(n_414),
.Y(n_470)
);

NOR2xp33_ASAP7_75t_SL g489 ( 
.A(n_470),
.B(n_474),
.Y(n_489)
);

INVx1_ASAP7_75t_L g471 ( 
.A(n_428),
.Y(n_471)
);

XNOR2xp5_ASAP7_75t_L g472 ( 
.A(n_426),
.B(n_391),
.Y(n_472)
);

MAJIxp5_ASAP7_75t_L g492 ( 
.A(n_472),
.B(n_477),
.C(n_421),
.Y(n_492)
);

AOI22xp5_ASAP7_75t_L g473 ( 
.A1(n_442),
.A2(n_382),
.B1(n_375),
.B2(n_392),
.Y(n_473)
);

NOR2xp33_ASAP7_75t_L g474 ( 
.A(n_432),
.B(n_363),
.Y(n_474)
);

XNOR2xp5_ASAP7_75t_SL g475 ( 
.A(n_426),
.B(n_385),
.Y(n_475)
);

XOR2xp5_ASAP7_75t_L g501 ( 
.A(n_475),
.B(n_439),
.Y(n_501)
);

NAND2xp5_ASAP7_75t_SL g476 ( 
.A(n_414),
.B(n_390),
.Y(n_476)
);

MAJIxp5_ASAP7_75t_L g477 ( 
.A(n_415),
.B(n_386),
.C(n_333),
.Y(n_477)
);

OAI21xp5_ASAP7_75t_L g478 ( 
.A1(n_420),
.A2(n_386),
.B(n_399),
.Y(n_478)
);

NAND2xp5_ASAP7_75t_L g494 ( 
.A(n_478),
.B(n_479),
.Y(n_494)
);

INVx1_ASAP7_75t_L g479 ( 
.A(n_435),
.Y(n_479)
);

OAI22xp5_ASAP7_75t_SL g480 ( 
.A1(n_455),
.A2(n_444),
.B1(n_442),
.B2(n_412),
.Y(n_480)
);

AOI22xp5_ASAP7_75t_L g518 ( 
.A1(n_480),
.A2(n_486),
.B1(n_487),
.B2(n_500),
.Y(n_518)
);

XNOR2xp5_ASAP7_75t_L g481 ( 
.A(n_449),
.B(n_410),
.Y(n_481)
);

XOR2xp5_ASAP7_75t_L g524 ( 
.A(n_481),
.B(n_483),
.Y(n_524)
);

XNOR2xp5_ASAP7_75t_L g483 ( 
.A(n_454),
.B(n_410),
.Y(n_483)
);

OAI22xp5_ASAP7_75t_SL g486 ( 
.A1(n_455),
.A2(n_444),
.B1(n_412),
.B2(n_443),
.Y(n_486)
);

XOR2xp5_ASAP7_75t_L g527 ( 
.A(n_492),
.B(n_495),
.Y(n_527)
);

XNOR2xp5_ASAP7_75t_L g495 ( 
.A(n_447),
.B(n_430),
.Y(n_495)
);

AOI22xp5_ASAP7_75t_L g498 ( 
.A1(n_471),
.A2(n_407),
.B1(n_436),
.B2(n_420),
.Y(n_498)
);

OAI22xp5_ASAP7_75t_SL g521 ( 
.A1(n_498),
.A2(n_478),
.B1(n_479),
.B2(n_425),
.Y(n_521)
);

NAND2xp5_ASAP7_75t_L g499 ( 
.A(n_472),
.B(n_430),
.Y(n_499)
);

INVx1_ASAP7_75t_L g515 ( 
.A(n_499),
.Y(n_515)
);

OAI22xp5_ASAP7_75t_SL g500 ( 
.A1(n_473),
.A2(n_418),
.B1(n_413),
.B2(n_429),
.Y(n_500)
);

XNOR2xp5_ASAP7_75t_SL g530 ( 
.A(n_501),
.B(n_343),
.Y(n_530)
);

OAI22xp5_ASAP7_75t_L g502 ( 
.A1(n_458),
.A2(n_431),
.B1(n_416),
.B2(n_425),
.Y(n_502)
);

INVx1_ASAP7_75t_L g522 ( 
.A(n_502),
.Y(n_522)
);

MAJIxp5_ASAP7_75t_L g504 ( 
.A(n_462),
.B(n_431),
.C(n_416),
.Y(n_504)
);

MAJIxp5_ASAP7_75t_L g520 ( 
.A(n_504),
.B(n_506),
.C(n_510),
.Y(n_520)
);

OAI22xp5_ASAP7_75t_L g505 ( 
.A1(n_456),
.A2(n_425),
.B1(n_424),
.B2(n_435),
.Y(n_505)
);

INVx1_ASAP7_75t_L g525 ( 
.A(n_505),
.Y(n_525)
);

MAJIxp5_ASAP7_75t_L g506 ( 
.A(n_459),
.B(n_451),
.C(n_477),
.Y(n_506)
);

XOR2xp5_ASAP7_75t_L g507 ( 
.A(n_461),
.B(n_440),
.Y(n_507)
);

XOR2xp5_ASAP7_75t_L g533 ( 
.A(n_507),
.B(n_343),
.Y(n_533)
);

NAND2xp5_ASAP7_75t_L g509 ( 
.A(n_445),
.B(n_464),
.Y(n_509)
);

INVx1_ASAP7_75t_L g532 ( 
.A(n_509),
.Y(n_532)
);

MAJIxp5_ASAP7_75t_L g510 ( 
.A(n_475),
.B(n_468),
.C(n_450),
.Y(n_510)
);

XNOR2xp5_ASAP7_75t_L g512 ( 
.A(n_488),
.B(n_460),
.Y(n_512)
);

XNOR2xp5_ASAP7_75t_L g549 ( 
.A(n_512),
.B(n_501),
.Y(n_549)
);

CKINVDCx16_ASAP7_75t_R g513 ( 
.A(n_509),
.Y(n_513)
);

NAND2xp5_ASAP7_75t_L g553 ( 
.A(n_513),
.B(n_514),
.Y(n_553)
);

NOR2xp33_ASAP7_75t_L g514 ( 
.A(n_485),
.B(n_456),
.Y(n_514)
);

NAND2xp5_ASAP7_75t_L g516 ( 
.A(n_480),
.B(n_446),
.Y(n_516)
);

INVx1_ASAP7_75t_L g556 ( 
.A(n_516),
.Y(n_556)
);

AOI22xp5_ASAP7_75t_SL g517 ( 
.A1(n_500),
.A2(n_463),
.B1(n_465),
.B2(n_467),
.Y(n_517)
);

OAI22xp5_ASAP7_75t_SL g551 ( 
.A1(n_517),
.A2(n_519),
.B1(n_528),
.B2(n_498),
.Y(n_551)
);

AOI22xp5_ASAP7_75t_L g519 ( 
.A1(n_486),
.A2(n_469),
.B1(n_453),
.B2(n_448),
.Y(n_519)
);

AOI22xp5_ASAP7_75t_L g558 ( 
.A1(n_521),
.A2(n_539),
.B1(n_490),
.B2(n_511),
.Y(n_558)
);

MAJIxp5_ASAP7_75t_L g523 ( 
.A(n_482),
.B(n_424),
.C(n_316),
.Y(n_523)
);

MAJIxp5_ASAP7_75t_L g546 ( 
.A(n_523),
.B(n_535),
.C(n_536),
.Y(n_546)
);

NAND2xp5_ASAP7_75t_L g526 ( 
.A(n_496),
.B(n_433),
.Y(n_526)
);

INVx1_ASAP7_75t_L g557 ( 
.A(n_526),
.Y(n_557)
);

AOI22xp5_ASAP7_75t_SL g528 ( 
.A1(n_510),
.A2(n_433),
.B1(n_386),
.B2(n_348),
.Y(n_528)
);

HB1xp67_ASAP7_75t_L g529 ( 
.A(n_499),
.Y(n_529)
);

CKINVDCx14_ASAP7_75t_R g554 ( 
.A(n_529),
.Y(n_554)
);

XNOR2xp5_ASAP7_75t_SL g548 ( 
.A(n_530),
.B(n_533),
.Y(n_548)
);

OAI21xp5_ASAP7_75t_SL g531 ( 
.A1(n_484),
.A2(n_372),
.B(n_380),
.Y(n_531)
);

NOR2xp33_ASAP7_75t_L g540 ( 
.A(n_531),
.B(n_534),
.Y(n_540)
);

INVx1_ASAP7_75t_L g534 ( 
.A(n_489),
.Y(n_534)
);

MAJIxp5_ASAP7_75t_L g535 ( 
.A(n_482),
.B(n_394),
.C(n_249),
.Y(n_535)
);

MAJIxp5_ASAP7_75t_L g536 ( 
.A(n_488),
.B(n_226),
.C(n_230),
.Y(n_536)
);

AO22x1_ASAP7_75t_L g537 ( 
.A1(n_508),
.A2(n_342),
.B1(n_242),
.B2(n_345),
.Y(n_537)
);

A2O1A1Ixp33_ASAP7_75t_SL g542 ( 
.A1(n_537),
.A2(n_497),
.B(n_494),
.C(n_508),
.Y(n_542)
);

MAJIxp5_ASAP7_75t_L g538 ( 
.A(n_504),
.B(n_345),
.C(n_298),
.Y(n_538)
);

MAJIxp5_ASAP7_75t_L g559 ( 
.A(n_538),
.B(n_536),
.C(n_523),
.Y(n_559)
);

CKINVDCx20_ASAP7_75t_R g539 ( 
.A(n_494),
.Y(n_539)
);

XOR2xp5_ASAP7_75t_L g541 ( 
.A(n_512),
.B(n_492),
.Y(n_541)
);

XOR2xp5_ASAP7_75t_L g561 ( 
.A(n_541),
.B(n_547),
.Y(n_561)
);

OAI22xp5_ASAP7_75t_L g564 ( 
.A1(n_542),
.A2(n_519),
.B1(n_517),
.B2(n_518),
.Y(n_564)
);

MAJIxp5_ASAP7_75t_L g543 ( 
.A(n_527),
.B(n_506),
.C(n_495),
.Y(n_543)
);

NOR2xp33_ASAP7_75t_L g563 ( 
.A(n_543),
.B(n_545),
.Y(n_563)
);

FAx1_ASAP7_75t_L g544 ( 
.A(n_521),
.B(n_497),
.CI(n_484),
.CON(n_544),
.SN(n_544)
);

NAND2xp5_ASAP7_75t_L g565 ( 
.A(n_544),
.B(n_516),
.Y(n_565)
);

BUFx24_ASAP7_75t_SL g545 ( 
.A(n_527),
.Y(n_545)
);

XOR2xp5_ASAP7_75t_L g547 ( 
.A(n_520),
.B(n_483),
.Y(n_547)
);

XOR2xp5_ASAP7_75t_L g566 ( 
.A(n_549),
.B(n_550),
.Y(n_566)
);

XOR2xp5_ASAP7_75t_L g550 ( 
.A(n_520),
.B(n_524),
.Y(n_550)
);

XOR2xp5_ASAP7_75t_L g568 ( 
.A(n_551),
.B(n_555),
.Y(n_568)
);

XNOR2xp5_ASAP7_75t_L g552 ( 
.A(n_524),
.B(n_481),
.Y(n_552)
);

MAJIxp5_ASAP7_75t_L g571 ( 
.A(n_552),
.B(n_559),
.C(n_560),
.Y(n_571)
);

XOR2xp5_ASAP7_75t_L g555 ( 
.A(n_530),
.B(n_507),
.Y(n_555)
);

INVx1_ASAP7_75t_L g562 ( 
.A(n_558),
.Y(n_562)
);

MAJIxp5_ASAP7_75t_L g560 ( 
.A(n_535),
.B(n_493),
.C(n_503),
.Y(n_560)
);

XOR2xp5_ASAP7_75t_L g590 ( 
.A(n_564),
.B(n_542),
.Y(n_590)
);

NAND2xp5_ASAP7_75t_L g579 ( 
.A(n_565),
.B(n_569),
.Y(n_579)
);

AOI21xp5_ASAP7_75t_L g567 ( 
.A1(n_540),
.A2(n_525),
.B(n_531),
.Y(n_567)
);

AOI21xp5_ASAP7_75t_L g589 ( 
.A1(n_567),
.A2(n_542),
.B(n_408),
.Y(n_589)
);

CKINVDCx20_ASAP7_75t_R g569 ( 
.A(n_553),
.Y(n_569)
);

NOR2xp33_ASAP7_75t_SL g570 ( 
.A(n_557),
.B(n_515),
.Y(n_570)
);

NOR2xp33_ASAP7_75t_SL g580 ( 
.A(n_570),
.B(n_578),
.Y(n_580)
);

XOR2xp5_ASAP7_75t_L g572 ( 
.A(n_541),
.B(n_533),
.Y(n_572)
);

XNOR2xp5_ASAP7_75t_L g582 ( 
.A(n_572),
.B(n_575),
.Y(n_582)
);

INVx11_ASAP7_75t_L g573 ( 
.A(n_554),
.Y(n_573)
);

NAND2xp5_ASAP7_75t_L g593 ( 
.A(n_573),
.B(n_574),
.Y(n_593)
);

MAJIxp5_ASAP7_75t_L g574 ( 
.A(n_547),
.B(n_538),
.C(n_522),
.Y(n_574)
);

OAI22xp5_ASAP7_75t_L g575 ( 
.A1(n_556),
.A2(n_518),
.B1(n_493),
.B2(n_532),
.Y(n_575)
);

MAJIxp5_ASAP7_75t_L g576 ( 
.A(n_559),
.B(n_528),
.C(n_526),
.Y(n_576)
);

MAJIxp5_ASAP7_75t_L g581 ( 
.A(n_576),
.B(n_546),
.C(n_550),
.Y(n_581)
);

OAI22xp5_ASAP7_75t_SL g577 ( 
.A1(n_544),
.A2(n_537),
.B1(n_490),
.B2(n_491),
.Y(n_577)
);

XNOR2xp5_ASAP7_75t_L g584 ( 
.A(n_577),
.B(n_548),
.Y(n_584)
);

NOR2xp33_ASAP7_75t_SL g578 ( 
.A(n_555),
.B(n_537),
.Y(n_578)
);

XNOR2xp5_ASAP7_75t_L g597 ( 
.A(n_581),
.B(n_589),
.Y(n_597)
);

MAJIxp5_ASAP7_75t_L g583 ( 
.A(n_561),
.B(n_546),
.C(n_548),
.Y(n_583)
);

NAND2xp5_ASAP7_75t_L g599 ( 
.A(n_583),
.B(n_585),
.Y(n_599)
);

XNOR2x1_ASAP7_75t_L g600 ( 
.A(n_584),
.B(n_590),
.Y(n_600)
);

XNOR2xp5_ASAP7_75t_L g585 ( 
.A(n_571),
.B(n_544),
.Y(n_585)
);

NOR2xp33_ASAP7_75t_L g586 ( 
.A(n_569),
.B(n_345),
.Y(n_586)
);

NAND2xp5_ASAP7_75t_L g601 ( 
.A(n_586),
.B(n_587),
.Y(n_601)
);

OAI22xp5_ASAP7_75t_SL g587 ( 
.A1(n_562),
.A2(n_542),
.B1(n_237),
.B2(n_232),
.Y(n_587)
);

NOR2xp33_ASAP7_75t_L g588 ( 
.A(n_563),
.B(n_570),
.Y(n_588)
);

NOR2xp33_ASAP7_75t_L g596 ( 
.A(n_588),
.B(n_591),
.Y(n_596)
);

NOR2xp33_ASAP7_75t_L g591 ( 
.A(n_571),
.B(n_574),
.Y(n_591)
);

NOR2xp33_ASAP7_75t_L g592 ( 
.A(n_576),
.B(n_562),
.Y(n_592)
);

NOR2xp33_ASAP7_75t_L g604 ( 
.A(n_592),
.B(n_566),
.Y(n_604)
);

OAI21xp5_ASAP7_75t_SL g594 ( 
.A1(n_579),
.A2(n_565),
.B(n_567),
.Y(n_594)
);

AOI21xp5_ASAP7_75t_L g609 ( 
.A1(n_594),
.A2(n_598),
.B(n_584),
.Y(n_609)
);

XOR2xp5_ASAP7_75t_L g595 ( 
.A(n_582),
.B(n_564),
.Y(n_595)
);

XOR2xp5_ASAP7_75t_L g610 ( 
.A(n_595),
.B(n_587),
.Y(n_610)
);

NOR2xp67_ASAP7_75t_L g598 ( 
.A(n_585),
.B(n_573),
.Y(n_598)
);

OAI22xp5_ASAP7_75t_L g602 ( 
.A1(n_580),
.A2(n_575),
.B1(n_577),
.B2(n_578),
.Y(n_602)
);

AOI22xp5_ASAP7_75t_L g611 ( 
.A1(n_602),
.A2(n_605),
.B1(n_568),
.B2(n_583),
.Y(n_611)
);

MAJIxp5_ASAP7_75t_L g603 ( 
.A(n_581),
.B(n_561),
.C(n_566),
.Y(n_603)
);

NAND2xp5_ASAP7_75t_L g607 ( 
.A(n_603),
.B(n_604),
.Y(n_607)
);

OAI22xp5_ASAP7_75t_SL g605 ( 
.A1(n_590),
.A2(n_568),
.B1(n_572),
.B2(n_593),
.Y(n_605)
);

NOR2xp67_ASAP7_75t_L g606 ( 
.A(n_597),
.B(n_603),
.Y(n_606)
);

OAI21xp5_ASAP7_75t_L g616 ( 
.A1(n_606),
.A2(n_609),
.B(n_612),
.Y(n_616)
);

NAND2xp5_ASAP7_75t_L g608 ( 
.A(n_596),
.B(n_582),
.Y(n_608)
);

NOR2xp33_ASAP7_75t_SL g615 ( 
.A(n_608),
.B(n_613),
.Y(n_615)
);

XNOR2xp5_ASAP7_75t_L g614 ( 
.A(n_610),
.B(n_611),
.Y(n_614)
);

INVxp67_ASAP7_75t_SL g612 ( 
.A(n_597),
.Y(n_612)
);

XNOR2xp5_ASAP7_75t_L g613 ( 
.A(n_599),
.B(n_600),
.Y(n_613)
);

NOR2xp33_ASAP7_75t_L g617 ( 
.A(n_607),
.B(n_594),
.Y(n_617)
);

NAND2xp5_ASAP7_75t_L g619 ( 
.A(n_617),
.B(n_618),
.Y(n_619)
);

NOR2xp33_ASAP7_75t_L g618 ( 
.A(n_612),
.B(n_595),
.Y(n_618)
);

NAND2xp5_ASAP7_75t_L g620 ( 
.A(n_616),
.B(n_601),
.Y(n_620)
);

NAND2xp5_ASAP7_75t_L g622 ( 
.A(n_620),
.B(n_621),
.Y(n_622)
);

INVxp67_ASAP7_75t_L g621 ( 
.A(n_615),
.Y(n_621)
);

NAND2xp5_ASAP7_75t_L g623 ( 
.A(n_619),
.B(n_614),
.Y(n_623)
);

NAND2xp5_ASAP7_75t_L g624 ( 
.A(n_623),
.B(n_614),
.Y(n_624)
);

BUFx24_ASAP7_75t_SL g625 ( 
.A(n_624),
.Y(n_625)
);

MAJIxp5_ASAP7_75t_L g626 ( 
.A(n_625),
.B(n_622),
.C(n_610),
.Y(n_626)
);

MAJIxp5_ASAP7_75t_L g627 ( 
.A(n_626),
.B(n_600),
.C(n_605),
.Y(n_627)
);


endmodule