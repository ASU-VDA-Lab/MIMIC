module fake_jpeg_527_n_221 (n_13, n_21, n_53, n_33, n_1, n_45, n_10, n_23, n_27, n_6, n_22, n_47, n_51, n_14, n_40, n_19, n_18, n_20, n_35, n_48, n_52, n_46, n_41, n_4, n_34, n_30, n_39, n_42, n_16, n_49, n_3, n_0, n_24, n_28, n_38, n_26, n_44, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_43, n_50, n_12, n_32, n_8, n_15, n_7, n_221);

input n_13;
input n_21;
input n_53;
input n_33;
input n_1;
input n_45;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_47;
input n_51;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_48;
input n_52;
input n_46;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_42;
input n_16;
input n_49;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_44;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_43;
input n_50;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_221;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_64;
wire n_55;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_84;
wire n_59;
wire n_98;
wire n_178;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_155;
wire n_207;
wire n_103;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_57;
wire n_171;
wire n_119;
wire n_69;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_143;
wire n_202;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_145;
wire n_108;
wire n_68;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_131;
wire n_56;
wire n_212;
wire n_211;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_216;
wire n_217;
wire n_184;
wire n_91;
wire n_93;
wire n_54;
wire n_161;
wire n_209;
wire n_208;
wire n_138;
wire n_101;
wire n_210;
wire n_149;
wire n_157;
wire n_87;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_46),
.Y(n_54)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_48),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_38),
.Y(n_56)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_3),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_44),
.Y(n_58)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_39),
.Y(n_59)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_8),
.Y(n_60)
);

INVx1_ASAP7_75t_SL g61 ( 
.A(n_31),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_47),
.Y(n_62)
);

CKINVDCx20_ASAP7_75t_R g63 ( 
.A(n_51),
.Y(n_63)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_18),
.Y(n_64)
);

BUFx2_ASAP7_75t_L g65 ( 
.A(n_36),
.Y(n_65)
);

INVx6_ASAP7_75t_SL g66 ( 
.A(n_25),
.Y(n_66)
);

CKINVDCx20_ASAP7_75t_R g67 ( 
.A(n_23),
.Y(n_67)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_17),
.Y(n_68)
);

BUFx12f_ASAP7_75t_L g69 ( 
.A(n_4),
.Y(n_69)
);

INVx11_ASAP7_75t_L g70 ( 
.A(n_19),
.Y(n_70)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_28),
.Y(n_71)
);

CKINVDCx20_ASAP7_75t_R g72 ( 
.A(n_33),
.Y(n_72)
);

INVx3_ASAP7_75t_L g73 ( 
.A(n_41),
.Y(n_73)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_22),
.Y(n_74)
);

BUFx6f_ASAP7_75t_L g75 ( 
.A(n_18),
.Y(n_75)
);

INVx8_ASAP7_75t_SL g76 ( 
.A(n_6),
.Y(n_76)
);

CKINVDCx20_ASAP7_75t_R g77 ( 
.A(n_40),
.Y(n_77)
);

INVx2_ASAP7_75t_L g78 ( 
.A(n_10),
.Y(n_78)
);

CKINVDCx20_ASAP7_75t_R g79 ( 
.A(n_34),
.Y(n_79)
);

CKINVDCx20_ASAP7_75t_R g80 ( 
.A(n_76),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_80),
.B(n_82),
.Y(n_92)
);

BUFx3_ASAP7_75t_L g81 ( 
.A(n_66),
.Y(n_81)
);

BUFx3_ASAP7_75t_L g95 ( 
.A(n_81),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_SL g82 ( 
.A(n_78),
.B(n_53),
.Y(n_82)
);

MAJIxp5_ASAP7_75t_L g83 ( 
.A(n_78),
.B(n_52),
.C(n_50),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_83),
.B(n_86),
.Y(n_93)
);

BUFx10_ASAP7_75t_L g84 ( 
.A(n_69),
.Y(n_84)
);

INVx4_ASAP7_75t_L g100 ( 
.A(n_84),
.Y(n_100)
);

INVx2_ASAP7_75t_L g85 ( 
.A(n_69),
.Y(n_85)
);

INVx2_ASAP7_75t_L g89 ( 
.A(n_85),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_SL g86 ( 
.A(n_57),
.B(n_60),
.Y(n_86)
);

BUFx5_ASAP7_75t_L g87 ( 
.A(n_66),
.Y(n_87)
);

INVx3_ASAP7_75t_L g88 ( 
.A(n_87),
.Y(n_88)
);

INVx6_ASAP7_75t_L g90 ( 
.A(n_81),
.Y(n_90)
);

BUFx2_ASAP7_75t_L g116 ( 
.A(n_90),
.Y(n_116)
);

OAI22xp5_ASAP7_75t_SL g91 ( 
.A1(n_82),
.A2(n_68),
.B1(n_75),
.B2(n_64),
.Y(n_91)
);

AOI22xp5_ASAP7_75t_L g112 ( 
.A1(n_91),
.A2(n_56),
.B1(n_58),
.B2(n_73),
.Y(n_112)
);

CKINVDCx20_ASAP7_75t_R g94 ( 
.A(n_86),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_SL g105 ( 
.A(n_94),
.B(n_57),
.Y(n_105)
);

BUFx6f_ASAP7_75t_L g96 ( 
.A(n_85),
.Y(n_96)
);

INVx5_ASAP7_75t_L g110 ( 
.A(n_96),
.Y(n_110)
);

AOI22xp5_ASAP7_75t_L g97 ( 
.A1(n_85),
.A2(n_64),
.B1(n_75),
.B2(n_68),
.Y(n_97)
);

OAI22xp5_ASAP7_75t_L g106 ( 
.A1(n_97),
.A2(n_99),
.B1(n_83),
.B2(n_70),
.Y(n_106)
);

AOI22xp33_ASAP7_75t_SL g98 ( 
.A1(n_80),
.A2(n_69),
.B1(n_70),
.B2(n_60),
.Y(n_98)
);

AOI22xp33_ASAP7_75t_SL g118 ( 
.A1(n_98),
.A2(n_61),
.B1(n_84),
.B2(n_81),
.Y(n_118)
);

OAI22xp5_ASAP7_75t_L g99 ( 
.A1(n_83),
.A2(n_58),
.B1(n_62),
.B2(n_56),
.Y(n_99)
);

INVx2_ASAP7_75t_L g101 ( 
.A(n_96),
.Y(n_101)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_101),
.Y(n_121)
);

INVx11_ASAP7_75t_L g102 ( 
.A(n_100),
.Y(n_102)
);

INVx3_ASAP7_75t_L g131 ( 
.A(n_102),
.Y(n_131)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_100),
.Y(n_103)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_103),
.Y(n_125)
);

CKINVDCx20_ASAP7_75t_R g104 ( 
.A(n_90),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_L g123 ( 
.A(n_104),
.B(n_107),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_SL g140 ( 
.A(n_105),
.B(n_113),
.Y(n_140)
);

AND2x2_ASAP7_75t_L g133 ( 
.A(n_106),
.B(n_112),
.Y(n_133)
);

OAI22xp5_ASAP7_75t_L g107 ( 
.A1(n_97),
.A2(n_65),
.B1(n_73),
.B2(n_62),
.Y(n_107)
);

OAI22xp33_ASAP7_75t_SL g108 ( 
.A1(n_93),
.A2(n_80),
.B1(n_65),
.B2(n_67),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_SL g122 ( 
.A(n_108),
.B(n_109),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_SL g109 ( 
.A(n_94),
.B(n_79),
.Y(n_109)
);

INVx2_ASAP7_75t_L g111 ( 
.A(n_89),
.Y(n_111)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_111),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_SL g113 ( 
.A(n_92),
.B(n_79),
.Y(n_113)
);

INVx3_ASAP7_75t_L g114 ( 
.A(n_88),
.Y(n_114)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_114),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_SL g115 ( 
.A(n_91),
.B(n_55),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_115),
.B(n_119),
.Y(n_127)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_89),
.Y(n_117)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_117),
.Y(n_137)
);

AOI21xp5_ASAP7_75t_L g141 ( 
.A1(n_118),
.A2(n_84),
.B(n_61),
.Y(n_141)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_88),
.Y(n_119)
);

MAJIxp5_ASAP7_75t_L g120 ( 
.A(n_117),
.B(n_99),
.C(n_71),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_L g151 ( 
.A(n_120),
.B(n_128),
.Y(n_151)
);

AND2x6_ASAP7_75t_L g124 ( 
.A(n_112),
.B(n_27),
.Y(n_124)
);

AOI21xp33_ASAP7_75t_L g157 ( 
.A1(n_124),
.A2(n_126),
.B(n_141),
.Y(n_157)
);

XNOR2xp5_ASAP7_75t_SL g126 ( 
.A(n_119),
.B(n_111),
.Y(n_126)
);

MAJIxp5_ASAP7_75t_L g128 ( 
.A(n_114),
.B(n_55),
.C(n_59),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_L g130 ( 
.A(n_104),
.B(n_67),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_L g149 ( 
.A(n_130),
.B(n_134),
.Y(n_149)
);

NOR2xp33_ASAP7_75t_L g134 ( 
.A(n_116),
.B(n_71),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_L g135 ( 
.A(n_101),
.B(n_74),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_L g150 ( 
.A(n_135),
.B(n_138),
.Y(n_150)
);

AND2x2_ASAP7_75t_L g136 ( 
.A(n_103),
.B(n_95),
.Y(n_136)
);

INVxp67_ASAP7_75t_SL g154 ( 
.A(n_136),
.Y(n_154)
);

NOR2xp33_ASAP7_75t_L g138 ( 
.A(n_116),
.B(n_59),
.Y(n_138)
);

OR2x2_ASAP7_75t_L g139 ( 
.A(n_102),
.B(n_95),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_SL g143 ( 
.A(n_139),
.B(n_110),
.Y(n_143)
);

AO21x2_ASAP7_75t_L g142 ( 
.A1(n_123),
.A2(n_110),
.B(n_74),
.Y(n_142)
);

INVxp67_ASAP7_75t_SL g173 ( 
.A(n_142),
.Y(n_173)
);

OR2x2_ASAP7_75t_L g166 ( 
.A(n_143),
.B(n_147),
.Y(n_166)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_137),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_L g171 ( 
.A(n_144),
.B(n_146),
.Y(n_171)
);

AOI21xp5_ASAP7_75t_L g145 ( 
.A1(n_139),
.A2(n_77),
.B(n_72),
.Y(n_145)
);

CKINVDCx16_ASAP7_75t_R g184 ( 
.A(n_145),
.Y(n_184)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_125),
.Y(n_146)
);

AOI22xp5_ASAP7_75t_SL g147 ( 
.A1(n_133),
.A2(n_127),
.B1(n_122),
.B2(n_141),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_SL g148 ( 
.A(n_140),
.B(n_63),
.Y(n_148)
);

NOR2xp33_ASAP7_75t_SL g174 ( 
.A(n_148),
.B(n_155),
.Y(n_174)
);

INVx2_ASAP7_75t_L g152 ( 
.A(n_129),
.Y(n_152)
);

INVx2_ASAP7_75t_L g167 ( 
.A(n_152),
.Y(n_167)
);

AO21x1_ASAP7_75t_SL g153 ( 
.A1(n_126),
.A2(n_87),
.B(n_84),
.Y(n_153)
);

AOI22xp5_ASAP7_75t_L g180 ( 
.A1(n_153),
.A2(n_156),
.B1(n_159),
.B2(n_12),
.Y(n_180)
);

NOR2xp33_ASAP7_75t_L g155 ( 
.A(n_128),
.B(n_54),
.Y(n_155)
);

O2A1O1Ixp33_ASAP7_75t_SL g156 ( 
.A1(n_133),
.A2(n_84),
.B(n_87),
.C(n_49),
.Y(n_156)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_121),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_L g182 ( 
.A(n_158),
.B(n_160),
.Y(n_182)
);

OAI22xp5_ASAP7_75t_SL g159 ( 
.A1(n_135),
.A2(n_84),
.B1(n_1),
.B2(n_2),
.Y(n_159)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_132),
.Y(n_160)
);

INVxp67_ASAP7_75t_L g161 ( 
.A(n_136),
.Y(n_161)
);

NOR2xp33_ASAP7_75t_L g178 ( 
.A(n_161),
.B(n_142),
.Y(n_178)
);

AOI22xp5_ASAP7_75t_L g162 ( 
.A1(n_120),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_162)
);

OAI22xp5_ASAP7_75t_L g172 ( 
.A1(n_162),
.A2(n_163),
.B1(n_164),
.B2(n_7),
.Y(n_172)
);

AOI22xp5_ASAP7_75t_L g163 ( 
.A1(n_124),
.A2(n_0),
.B1(n_3),
.B2(n_4),
.Y(n_163)
);

AOI22xp5_ASAP7_75t_L g164 ( 
.A1(n_131),
.A2(n_45),
.B1(n_43),
.B2(n_42),
.Y(n_164)
);

OAI21xp5_ASAP7_75t_L g165 ( 
.A1(n_131),
.A2(n_5),
.B(n_6),
.Y(n_165)
);

XNOR2xp5_ASAP7_75t_L g169 ( 
.A(n_165),
.B(n_5),
.Y(n_169)
);

MAJIxp5_ASAP7_75t_L g168 ( 
.A(n_151),
.B(n_37),
.C(n_35),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_SL g194 ( 
.A(n_168),
.B(n_172),
.Y(n_194)
);

NOR2xp33_ASAP7_75t_L g185 ( 
.A(n_169),
.B(n_177),
.Y(n_185)
);

OAI22xp5_ASAP7_75t_SL g170 ( 
.A1(n_147),
.A2(n_7),
.B1(n_8),
.B2(n_9),
.Y(n_170)
);

AOI22xp5_ASAP7_75t_L g189 ( 
.A1(n_170),
.A2(n_175),
.B1(n_176),
.B2(n_13),
.Y(n_189)
);

OAI22xp5_ASAP7_75t_SL g175 ( 
.A1(n_142),
.A2(n_157),
.B1(n_150),
.B2(n_154),
.Y(n_175)
);

OAI22xp5_ASAP7_75t_SL g176 ( 
.A1(n_142),
.A2(n_9),
.B1(n_10),
.B2(n_11),
.Y(n_176)
);

XNOR2xp5_ASAP7_75t_L g177 ( 
.A(n_154),
.B(n_161),
.Y(n_177)
);

NOR2xp33_ASAP7_75t_L g186 ( 
.A(n_178),
.B(n_179),
.Y(n_186)
);

NOR2xp33_ASAP7_75t_SL g179 ( 
.A(n_149),
.B(n_11),
.Y(n_179)
);

OAI22xp5_ASAP7_75t_L g193 ( 
.A1(n_180),
.A2(n_181),
.B1(n_15),
.B2(n_16),
.Y(n_193)
);

AOI22xp5_ASAP7_75t_L g181 ( 
.A1(n_153),
.A2(n_12),
.B1(n_13),
.B2(n_14),
.Y(n_181)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_165),
.Y(n_183)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_183),
.Y(n_187)
);

AOI21xp5_ASAP7_75t_L g188 ( 
.A1(n_166),
.A2(n_156),
.B(n_164),
.Y(n_188)
);

NAND2xp33_ASAP7_75t_SL g198 ( 
.A(n_188),
.B(n_181),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_L g196 ( 
.A(n_189),
.B(n_191),
.Y(n_196)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_182),
.Y(n_190)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_190),
.Y(n_202)
);

NAND2xp5_ASAP7_75t_L g191 ( 
.A(n_177),
.B(n_32),
.Y(n_191)
);

NOR2xp33_ASAP7_75t_L g192 ( 
.A(n_174),
.B(n_14),
.Y(n_192)
);

XNOR2xp5_ASAP7_75t_L g203 ( 
.A(n_192),
.B(n_26),
.Y(n_203)
);

AOI22xp5_ASAP7_75t_L g200 ( 
.A1(n_193),
.A2(n_195),
.B1(n_169),
.B2(n_194),
.Y(n_200)
);

OAI22xp5_ASAP7_75t_L g195 ( 
.A1(n_173),
.A2(n_15),
.B1(n_16),
.B2(n_17),
.Y(n_195)
);

MAJIxp5_ASAP7_75t_L g197 ( 
.A(n_187),
.B(n_166),
.C(n_168),
.Y(n_197)
);

MAJIxp5_ASAP7_75t_L g207 ( 
.A(n_197),
.B(n_204),
.C(n_199),
.Y(n_207)
);

NAND2xp5_ASAP7_75t_SL g205 ( 
.A(n_198),
.B(n_200),
.Y(n_205)
);

XOR2x1_ASAP7_75t_SL g199 ( 
.A(n_188),
.B(n_184),
.Y(n_199)
);

MAJIxp5_ASAP7_75t_L g208 ( 
.A(n_199),
.B(n_201),
.C(n_203),
.Y(n_208)
);

MAJIxp5_ASAP7_75t_L g201 ( 
.A(n_191),
.B(n_171),
.C(n_167),
.Y(n_201)
);

CKINVDCx20_ASAP7_75t_R g204 ( 
.A(n_186),
.Y(n_204)
);

XOR2xp5_ASAP7_75t_L g206 ( 
.A(n_197),
.B(n_185),
.Y(n_206)
);

NOR2xp33_ASAP7_75t_L g211 ( 
.A(n_206),
.B(n_207),
.Y(n_211)
);

FAx1_ASAP7_75t_SL g209 ( 
.A(n_198),
.B(n_189),
.CI(n_173),
.CON(n_209),
.SN(n_209)
);

OAI22xp5_ASAP7_75t_SL g212 ( 
.A1(n_209),
.A2(n_24),
.B1(n_30),
.B2(n_21),
.Y(n_212)
);

AOI22xp5_ASAP7_75t_L g210 ( 
.A1(n_205),
.A2(n_202),
.B1(n_196),
.B2(n_29),
.Y(n_210)
);

MAJIxp5_ASAP7_75t_L g213 ( 
.A(n_210),
.B(n_212),
.C(n_208),
.Y(n_213)
);

NOR2xp33_ASAP7_75t_SL g215 ( 
.A(n_213),
.B(n_214),
.Y(n_215)
);

NOR2x1_ASAP7_75t_L g214 ( 
.A(n_211),
.B(n_207),
.Y(n_214)
);

OAI21xp5_ASAP7_75t_SL g216 ( 
.A1(n_215),
.A2(n_210),
.B(n_212),
.Y(n_216)
);

INVxp67_ASAP7_75t_L g217 ( 
.A(n_216),
.Y(n_217)
);

CKINVDCx20_ASAP7_75t_R g218 ( 
.A(n_217),
.Y(n_218)
);

MAJIxp5_ASAP7_75t_L g219 ( 
.A(n_218),
.B(n_206),
.C(n_209),
.Y(n_219)
);

XNOR2xp5_ASAP7_75t_L g220 ( 
.A(n_219),
.B(n_19),
.Y(n_220)
);

AOI22xp5_ASAP7_75t_L g221 ( 
.A1(n_220),
.A2(n_20),
.B1(n_21),
.B2(n_212),
.Y(n_221)
);


endmodule