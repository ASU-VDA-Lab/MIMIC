module fake_jpeg_21964_n_32 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_32);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_32;

wire n_21;
wire n_23;
wire n_27;
wire n_22;
wire n_19;
wire n_20;
wire n_18;
wire n_30;
wire n_16;
wire n_24;
wire n_28;
wire n_26;
wire n_17;
wire n_25;
wire n_31;
wire n_29;

BUFx4f_ASAP7_75t_SL g16 ( 
.A(n_12),
.Y(n_16)
);

BUFx6f_ASAP7_75t_L g17 ( 
.A(n_9),
.Y(n_17)
);

INVx5_ASAP7_75t_L g18 ( 
.A(n_14),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_5),
.Y(n_19)
);

INVx2_ASAP7_75t_L g20 ( 
.A(n_16),
.Y(n_20)
);

MAJIxp5_ASAP7_75t_L g26 ( 
.A(n_20),
.B(n_15),
.C(n_2),
.Y(n_26)
);

BUFx10_ASAP7_75t_L g21 ( 
.A(n_18),
.Y(n_21)
);

AO21x1_ASAP7_75t_L g25 ( 
.A1(n_21),
.A2(n_23),
.B(n_19),
.Y(n_25)
);

AOI21xp5_ASAP7_75t_L g22 ( 
.A1(n_19),
.A2(n_7),
.B(n_1),
.Y(n_22)
);

XNOR2xp5_ASAP7_75t_L g24 ( 
.A(n_22),
.B(n_8),
.Y(n_24)
);

BUFx3_ASAP7_75t_L g23 ( 
.A(n_17),
.Y(n_23)
);

MAJIxp5_ASAP7_75t_SL g28 ( 
.A(n_24),
.B(n_25),
.C(n_26),
.Y(n_28)
);

OAI22xp5_ASAP7_75t_SL g27 ( 
.A1(n_22),
.A2(n_3),
.B1(n_4),
.B2(n_6),
.Y(n_27)
);

FAx1_ASAP7_75t_L g29 ( 
.A(n_27),
.B(n_10),
.CI(n_11),
.CON(n_29),
.SN(n_29)
);

AOI21xp5_ASAP7_75t_SL g30 ( 
.A1(n_29),
.A2(n_13),
.B(n_0),
.Y(n_30)
);

NOR2xp33_ASAP7_75t_SL g31 ( 
.A(n_30),
.B(n_28),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_31),
.Y(n_32)
);


endmodule