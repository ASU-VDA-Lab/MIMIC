module real_aes_18286_n_376 (n_76, n_113, n_187, n_90, n_257, n_65, n_74, n_185, n_285, n_30, n_222, n_61, n_20, n_287, n_357, n_64, n_254, n_207, n_10, n_83, n_181, n_362, n_124, n_191, n_209, n_299, n_322, n_328, n_19, n_40, n_318, n_355, n_239, n_100, n_54, n_112, n_319, n_364, n_35, n_42, n_329, n_132, n_131, n_144, n_169, n_242, n_308, n_172, n_341, n_232, n_6, n_69, n_317, n_353, n_321, n_73, n_320, n_77, n_260, n_37, n_97, n_186, n_138, n_374, n_26, n_235, n_245, n_161, n_189, n_271, n_2, n_145, n_227, n_92, n_330, n_332, n_292, n_116, n_94, n_289, n_280, n_333, n_213, n_356, n_184, n_28, n_372, n_202, n_56, n_370, n_34, n_98, n_121, n_352, n_125, n_216, n_82, n_327, n_47, n_106, n_32, n_263, n_230, n_51, n_248, n_301, n_27, n_343, n_369, n_174, n_18, n_104, n_211, n_281, n_173, n_234, n_284, n_153, n_316, n_75, n_178, n_298, n_49, n_43, n_297, n_9, n_119, n_310, n_164, n_231, n_44, n_102, n_122, n_141, n_128, n_111, n_167, n_80, n_179, n_12, n_68, n_129, n_345, n_304, n_311, n_324, n_25, n_278, n_236, n_367, n_267, n_218, n_48, n_204, n_339, n_89, n_277, n_331, n_93, n_182, n_363, n_323, n_199, n_350, n_142, n_223, n_67, n_368, n_250, n_85, n_45, n_5, n_244, n_118, n_139, n_87, n_171, n_78, n_146, n_17, n_226, n_255, n_286, n_120, n_261, n_238, n_360, n_58, n_165, n_361, n_246, n_176, n_163, n_29, n_52, n_251, n_220, n_197, n_296, n_3, n_41, n_256, n_71, n_302, n_351, n_126, n_200, n_115, n_96, n_110, n_150, n_147, n_288, n_23, n_334, n_274, n_160, n_303, n_95, n_188, n_269, n_201, n_306, n_158, n_4, n_366, n_346, n_193, n_293, n_162, n_358, n_275, n_214, n_46, n_109, n_59, n_203, n_81, n_133, n_273, n_114, n_276, n_295, n_265, n_354, n_154, n_127, n_326, n_24, n_217, n_55, n_62, n_291, n_148, n_88, n_159, n_11, n_108, n_373, n_60, n_233, n_290, n_365, n_155, n_243, n_268, n_136, n_157, n_282, n_101, n_309, n_344, n_229, n_107, n_33, n_53, n_36, n_149, n_190, n_262, n_134, n_349, n_336, n_195, n_300, n_252, n_283, n_314, n_249, n_221, n_156, n_359, n_57, n_66, n_21, n_31, n_8, n_312, n_183, n_266, n_205, n_335, n_177, n_313, n_22, n_140, n_219, n_180, n_212, n_210, n_325, n_338, n_371, n_103, n_166, n_224, n_151, n_130, n_253, n_99, n_15, n_72, n_152, n_198, n_7, n_228, n_272, n_196, n_347, n_315, n_123, n_279, n_79, n_270, n_305, n_117, n_208, n_215, n_135, n_70, n_50, n_170, n_86, n_375, n_340, n_13, n_168, n_175, n_241, n_105, n_84, n_294, n_258, n_206, n_307, n_342, n_348, n_14, n_194, n_137, n_225, n_16, n_39, n_337, n_247, n_240, n_38, n_259, n_143, n_192, n_0, n_264, n_63, n_1, n_237, n_91, n_376);
input n_76;
input n_113;
input n_187;
input n_90;
input n_257;
input n_65;
input n_74;
input n_185;
input n_285;
input n_30;
input n_222;
input n_61;
input n_20;
input n_287;
input n_357;
input n_64;
input n_254;
input n_207;
input n_10;
input n_83;
input n_181;
input n_362;
input n_124;
input n_191;
input n_209;
input n_299;
input n_322;
input n_328;
input n_19;
input n_40;
input n_318;
input n_355;
input n_239;
input n_100;
input n_54;
input n_112;
input n_319;
input n_364;
input n_35;
input n_42;
input n_329;
input n_132;
input n_131;
input n_144;
input n_169;
input n_242;
input n_308;
input n_172;
input n_341;
input n_232;
input n_6;
input n_69;
input n_317;
input n_353;
input n_321;
input n_73;
input n_320;
input n_77;
input n_260;
input n_37;
input n_97;
input n_186;
input n_138;
input n_374;
input n_26;
input n_235;
input n_245;
input n_161;
input n_189;
input n_271;
input n_2;
input n_145;
input n_227;
input n_92;
input n_330;
input n_332;
input n_292;
input n_116;
input n_94;
input n_289;
input n_280;
input n_333;
input n_213;
input n_356;
input n_184;
input n_28;
input n_372;
input n_202;
input n_56;
input n_370;
input n_34;
input n_98;
input n_121;
input n_352;
input n_125;
input n_216;
input n_82;
input n_327;
input n_47;
input n_106;
input n_32;
input n_263;
input n_230;
input n_51;
input n_248;
input n_301;
input n_27;
input n_343;
input n_369;
input n_174;
input n_18;
input n_104;
input n_211;
input n_281;
input n_173;
input n_234;
input n_284;
input n_153;
input n_316;
input n_75;
input n_178;
input n_298;
input n_49;
input n_43;
input n_297;
input n_9;
input n_119;
input n_310;
input n_164;
input n_231;
input n_44;
input n_102;
input n_122;
input n_141;
input n_128;
input n_111;
input n_167;
input n_80;
input n_179;
input n_12;
input n_68;
input n_129;
input n_345;
input n_304;
input n_311;
input n_324;
input n_25;
input n_278;
input n_236;
input n_367;
input n_267;
input n_218;
input n_48;
input n_204;
input n_339;
input n_89;
input n_277;
input n_331;
input n_93;
input n_182;
input n_363;
input n_323;
input n_199;
input n_350;
input n_142;
input n_223;
input n_67;
input n_368;
input n_250;
input n_85;
input n_45;
input n_5;
input n_244;
input n_118;
input n_139;
input n_87;
input n_171;
input n_78;
input n_146;
input n_17;
input n_226;
input n_255;
input n_286;
input n_120;
input n_261;
input n_238;
input n_360;
input n_58;
input n_165;
input n_361;
input n_246;
input n_176;
input n_163;
input n_29;
input n_52;
input n_251;
input n_220;
input n_197;
input n_296;
input n_3;
input n_41;
input n_256;
input n_71;
input n_302;
input n_351;
input n_126;
input n_200;
input n_115;
input n_96;
input n_110;
input n_150;
input n_147;
input n_288;
input n_23;
input n_334;
input n_274;
input n_160;
input n_303;
input n_95;
input n_188;
input n_269;
input n_201;
input n_306;
input n_158;
input n_4;
input n_366;
input n_346;
input n_193;
input n_293;
input n_162;
input n_358;
input n_275;
input n_214;
input n_46;
input n_109;
input n_59;
input n_203;
input n_81;
input n_133;
input n_273;
input n_114;
input n_276;
input n_295;
input n_265;
input n_354;
input n_154;
input n_127;
input n_326;
input n_24;
input n_217;
input n_55;
input n_62;
input n_291;
input n_148;
input n_88;
input n_159;
input n_11;
input n_108;
input n_373;
input n_60;
input n_233;
input n_290;
input n_365;
input n_155;
input n_243;
input n_268;
input n_136;
input n_157;
input n_282;
input n_101;
input n_309;
input n_344;
input n_229;
input n_107;
input n_33;
input n_53;
input n_36;
input n_149;
input n_190;
input n_262;
input n_134;
input n_349;
input n_336;
input n_195;
input n_300;
input n_252;
input n_283;
input n_314;
input n_249;
input n_221;
input n_156;
input n_359;
input n_57;
input n_66;
input n_21;
input n_31;
input n_8;
input n_312;
input n_183;
input n_266;
input n_205;
input n_335;
input n_177;
input n_313;
input n_22;
input n_140;
input n_219;
input n_180;
input n_212;
input n_210;
input n_325;
input n_338;
input n_371;
input n_103;
input n_166;
input n_224;
input n_151;
input n_130;
input n_253;
input n_99;
input n_15;
input n_72;
input n_152;
input n_198;
input n_7;
input n_228;
input n_272;
input n_196;
input n_347;
input n_315;
input n_123;
input n_279;
input n_79;
input n_270;
input n_305;
input n_117;
input n_208;
input n_215;
input n_135;
input n_70;
input n_50;
input n_170;
input n_86;
input n_375;
input n_340;
input n_13;
input n_168;
input n_175;
input n_241;
input n_105;
input n_84;
input n_294;
input n_258;
input n_206;
input n_307;
input n_342;
input n_348;
input n_14;
input n_194;
input n_137;
input n_225;
input n_16;
input n_39;
input n_337;
input n_247;
input n_240;
input n_38;
input n_259;
input n_143;
input n_192;
input n_0;
input n_264;
input n_63;
input n_1;
input n_237;
input n_91;
output n_376;
wire n_476;
wire n_599;
wire n_887;
wire n_1279;
wire n_1314;
wire n_830;
wire n_1371;
wire n_624;
wire n_618;
wire n_1797;
wire n_933;
wire n_485;
wire n_822;
wire n_1641;
wire n_750;
wire n_503;
wire n_1781;
wire n_1762;
wire n_1591;
wire n_1903;
wire n_469;
wire n_1310;
wire n_1376;
wire n_592;
wire n_1621;
wire n_1729;
wire n_1929;
wire n_1737;
wire n_761;
wire n_421;
wire n_919;
wire n_1217;
wire n_1888;
wire n_1423;
wire n_571;
wire n_549;
wire n_1034;
wire n_1328;
wire n_1219;
wire n_952;
wire n_1166;
wire n_752;
wire n_448;
wire n_556;
wire n_593;
wire n_989;
wire n_431;
wire n_1044;
wire n_1730;
wire n_1744;
wire n_963;
wire n_551;
wire n_884;
wire n_814;
wire n_944;
wire n_1936;
wire n_1283;
wire n_983;
wire n_955;
wire n_975;
wire n_941;
wire n_1313;
wire n_1873;
wire n_1835;
wire n_1871;
wire n_1468;
wire n_1713;
wire n_1967;
wire n_1920;
wire n_870;
wire n_1248;
wire n_1602;
wire n_548;
wire n_1859;
wire n_572;
wire n_815;
wire n_1140;
wire n_1520;
wire n_1453;
wire n_786;
wire n_512;
wire n_395;
wire n_795;
wire n_1379;
wire n_400;
wire n_1597;
wire n_1845;
wire n_1415;
wire n_1160;
wire n_1849;
wire n_1287;
wire n_883;
wire n_478;
wire n_1575;
wire n_1687;
wire n_553;
wire n_1805;
wire n_1367;
wire n_744;
wire n_1325;
wire n_1382;
wire n_1441;
wire n_875;
wire n_1199;
wire n_951;
wire n_1225;
wire n_1543;
wire n_791;
wire n_976;
wire n_636;
wire n_906;
wire n_477;
wire n_1833;
wire n_1477;
wire n_1944;
wire n_1893;
wire n_595;
wire n_1960;
wire n_1282;
wire n_683;
wire n_840;
wire n_570;
wire n_675;
wire n_835;
wire n_732;
wire n_784;
wire n_962;
wire n_1599;
wire n_1959;
wire n_755;
wire n_409;
wire n_781;
wire n_576;
wire n_1688;
wire n_956;
wire n_1242;
wire n_1537;
wire n_874;
wire n_796;
wire n_1126;
wire n_383;
wire n_1607;
wire n_455;
wire n_1771;
wire n_1809;
wire n_682;
wire n_1745;
wire n_1820;
wire n_812;
wire n_782;
wire n_817;
wire n_1883;
wire n_608;
wire n_760;
wire n_534;
wire n_1454;
wire n_708;
wire n_1020;
wire n_885;
wire n_950;
wire n_381;
wire n_1196;
wire n_1013;
wire n_1905;
wire n_808;
wire n_1639;
wire n_1224;
wire n_1872;
wire n_1694;
wire n_688;
wire n_1042;
wire n_1588;
wire n_1317;
wire n_417;
wire n_690;
wire n_1419;
wire n_499;
wire n_1142;
wire n_1731;
wire n_1589;
wire n_947;
wire n_970;
wire n_1677;
wire n_1149;
wire n_527;
wire n_1676;
wire n_1342;
wire n_1440;
wire n_1966;
wire n_552;
wire n_1346;
wire n_1383;
wire n_1890;
wire n_1675;
wire n_1954;
wire n_590;
wire n_1293;
wire n_1880;
wire n_432;
wire n_1882;
wire n_1131;
wire n_1008;
wire n_1491;
wire n_1865;
wire n_805;
wire n_1600;
wire n_619;
wire n_1095;
wire n_1284;
wire n_1583;
wire n_1250;
wire n_1465;
wire n_859;
wire n_1486;
wire n_1304;
wire n_685;
wire n_1080;
wire n_917;
wire n_1247;
wire n_488;
wire n_501;
wire n_1380;
wire n_1658;
wire n_1866;
wire n_954;
wire n_702;
wire n_1874;
wire n_1007;
wire n_1906;
wire n_898;
wire n_1926;
wire n_562;
wire n_1897;
wire n_1022;
wire n_1502;
wire n_404;
wire n_1073;
wire n_1632;
wire n_728;
wire n_1301;
wire n_1201;
wire n_997;
wire n_1105;
wire n_1768;
wire n_1243;
wire n_1846;
wire n_1003;
wire n_749;
wire n_1870;
wire n_914;
wire n_1837;
wire n_1286;
wire n_494;
wire n_1661;
wire n_927;
wire n_723;
wire n_972;
wire n_1351;
wire n_1813;
wire n_1628;
wire n_1587;
wire n_1821;
wire n_1570;
wire n_1209;
wire n_411;
wire n_498;
wire n_1397;
wire n_765;
wire n_1554;
wire n_648;
wire n_1487;
wire n_939;
wire n_1825;
wire n_1615;
wire n_1763;
wire n_928;
wire n_1384;
wire n_789;
wire n_1515;
wire n_738;
wire n_1387;
wire n_922;
wire n_1956;
wire n_1048;
wire n_1422;
wire n_787;
wire n_1214;
wire n_806;
wire n_1940;
wire n_715;
wire n_1714;
wire n_420;
wire n_1666;
wire n_1490;
wire n_1258;
wire n_873;
wire n_438;
wire n_1814;
wire n_446;
wire n_1281;
wire n_1559;
wire n_1510;
wire n_1495;
wire n_1727;
wire n_712;
wire n_1921;
wire n_422;
wire n_861;
wire n_1574;
wire n_479;
wire n_825;
wire n_541;
wire n_839;
wire n_811;
wire n_558;
wire n_1742;
wire n_724;
wire n_1648;
wire n_1914;
wire n_440;
wire n_1945;
wire n_1231;
wire n_1305;
wire n_1161;
wire n_686;
wire n_1299;
wire n_949;
wire n_586;
wire n_1508;
wire n_1421;
wire n_788;
wire n_441;
wire n_1045;
wire n_1339;
wire n_1793;
wire n_837;
wire n_1349;
wire n_1708;
wire n_1445;
wire n_1631;
wire n_829;
wire n_1030;
wire n_1348;
wire n_1391;
wire n_597;
wire n_1036;
wire n_687;
wire n_1751;
wire n_1765;
wire n_1538;
wire n_652;
wire n_500;
wire n_804;
wire n_1173;
wire n_854;
wire n_1787;
wire n_424;
wire n_877;
wire n_802;
wire n_1876;
wire n_1488;
wire n_1572;
wire n_1514;
wire n_480;
wire n_1652;
wire n_684;
wire n_1178;
wire n_1531;
wire n_821;
wire n_1657;
wire n_1616;
wire n_1828;
wire n_1860;
wire n_1563;
wire n_1018;
wire n_980;
wire n_1233;
wire n_1106;
wire n_1205;
wire n_838;
wire n_1561;
wire n_635;
wire n_792;
wire n_1542;
wire n_1392;
wire n_665;
wire n_667;
wire n_991;
wire n_1712;
wire n_1556;
wire n_580;
wire n_1004;
wire n_1370;
wire n_1417;
wire n_1703;
wire n_1717;
wire n_1723;
wire n_1951;
wire n_979;
wire n_445;
wire n_596;
wire n_1740;
wire n_1197;
wire n_657;
wire n_1260;
wire n_1606;
wire n_1129;
wire n_1760;
wire n_1285;
wire n_742;
wire n_1014;
wire n_1385;
wire n_1629;
wire n_1618;
wire n_461;
wire n_1770;
wire n_1047;
wire n_1016;
wire n_1545;
wire n_694;
wire n_1350;
wire n_894;
wire n_1750;
wire n_1852;
wire n_545;
wire n_1459;
wire n_1530;
wire n_401;
wire n_538;
wire n_1830;
wire n_1594;
wire n_1864;
wire n_537;
wire n_1767;
wire n_1651;
wire n_560;
wire n_1094;
wire n_1776;
wire n_1719;
wire n_1220;
wire n_696;
wire n_1147;
wire n_1425;
wire n_1613;
wire n_1504;
wire n_704;
wire n_453;
wire n_647;
wire n_399;
wire n_1499;
wire n_700;
wire n_948;
wire n_677;
wire n_1269;
wire n_378;
wire n_591;
wire n_1635;
wire n_1518;
wire n_1702;
wire n_1366;
wire n_678;
wire n_415;
wire n_1400;
wire n_564;
wire n_638;
wire n_1361;
wire n_510;
wire n_1358;
wire n_1577;
wire n_1839;
wire n_1642;
wire n_1406;
wire n_550;
wire n_966;
wire n_1881;
wire n_1568;
wire n_1368;
wire n_994;
wire n_384;
wire n_1479;
wire n_1612;
wire n_1128;
wire n_1098;
wire n_824;
wire n_1238;
wire n_1611;
wire n_992;
wire n_813;
wire n_981;
wire n_1338;
wire n_1884;
wire n_1182;
wire n_872;
wire n_1401;
wire n_1946;
wire n_1086;
wire n_1070;
wire n_1189;
wire n_1665;
wire n_535;
wire n_882;
wire n_1210;
wire n_1741;
wire n_1456;
wire n_1879;
wire n_746;
wire n_1614;
wire n_656;
wire n_1148;
wire n_860;
wire n_748;
wire n_1261;
wire n_1062;
wire n_1439;
wire n_651;
wire n_1585;
wire n_1500;
wire n_801;
wire n_1271;
wire n_1653;
wire n_529;
wire n_504;
wire n_973;
wire n_1364;
wire n_1853;
wire n_659;
wire n_634;
wire n_903;
wire n_1668;
wire n_565;
wire n_925;
wire n_1389;
wire n_1393;
wire n_1930;
wire n_457;
wire n_1121;
wire n_1059;
wire n_493;
wire n_1362;
wire n_610;
wire n_1035;
wire n_620;
wire n_722;
wire n_1174;
wire n_1193;
wire n_1553;
wire n_754;
wire n_508;
wire n_1141;
wire n_1769;
wire n_1812;
wire n_1112;
wire n_1485;
wire n_1408;
wire n_1680;
wire n_428;
wire n_783;
wire n_1107;
wire n_1564;
wire n_505;
wire n_600;
wire n_731;
wire n_964;
wire n_605;
wire n_1516;
wire n_1386;
wire n_406;
wire n_1493;
wire n_1579;
wire n_1854;
wire n_617;
wire n_1404;
wire n_402;
wire n_602;
wire n_733;
wire n_658;
wire n_676;
wire n_1856;
wire n_531;
wire n_1848;
wire n_1031;
wire n_1394;
wire n_807;
wire n_1011;
wire n_416;
wire n_1567;
wire n_1569;
wire n_895;
wire n_799;
wire n_490;
wire n_391;
wire n_695;
wire n_1181;
wire n_881;
wire n_1626;
wire n_645;
wire n_1145;
wire n_1529;
wire n_557;
wire n_1681;
wire n_1620;
wire n_777;
wire n_985;
wire n_1659;
wire n_910;
wire n_642;
wire n_613;
wire n_1773;
wire n_1125;
wire n_1347;
wire n_1655;
wire n_1766;
wire n_1522;
wire n_1163;
wire n_1278;
wire n_734;
wire n_1623;
wire n_1907;
wire n_735;
wire n_1179;
wire n_569;
wire n_1171;
wire n_785;
wire n_1203;
wire n_1716;
wire n_1232;
wire n_471;
wire n_1857;
wire n_853;
wire n_810;
wire n_1136;
wire n_699;
wire n_1580;
wire n_1000;
wire n_1187;
wire n_649;
wire n_1234;
wire n_1915;
wire n_622;
wire n_1634;
wire n_1353;
wire n_1002;
wire n_1165;
wire n_1551;
wire n_1667;
wire n_1058;
wire n_1216;
wire n_662;
wire n_1862;
wire n_1965;
wire n_850;
wire n_720;
wire n_1026;
wire n_1756;
wire n_1803;
wire n_492;
wire n_407;
wire n_419;
wire n_1023;
wire n_730;
wire n_1699;
wire n_1794;
wire n_1748;
wire n_643;
wire n_1403;
wire n_486;
wire n_779;
wire n_481;
wire n_691;
wire n_589;
wire n_526;
wire n_1513;
wire n_1194;
wire n_389;
wire n_1609;
wire n_1462;
wire n_701;
wire n_1934;
wire n_809;
wire n_1532;
wire n_679;
wire n_520;
wire n_926;
wire n_1643;
wire n_942;
wire n_1374;
wire n_1120;
wire n_1497;
wire n_1548;
wire n_1784;
wire n_1526;
wire n_689;
wire n_1483;
wire n_946;
wire n_753;
wire n_1409;
wire n_1188;
wire n_623;
wire n_1474;
wire n_1032;
wire n_1431;
wire n_721;
wire n_1806;
wire n_1829;
wire n_1133;
wire n_1775;
wire n_1593;
wire n_739;
wire n_1322;
wire n_1525;
wire n_1732;
wire n_1162;
wire n_1463;
wire n_1524;
wire n_762;
wire n_1298;
wire n_442;
wire n_1633;
wire n_740;
wire n_1686;
wire n_1357;
wire n_639;
wire n_1186;
wire n_1365;
wire n_1807;
wire n_459;
wire n_1172;
wire n_998;
wire n_1689;
wire n_1625;
wire n_1910;
wire n_1395;
wire n_1276;
wire n_836;
wire n_1733;
wire n_1957;
wire n_1184;
wire n_583;
wire n_414;
wire n_1336;
wire n_776;
wire n_1138;
wire n_890;
wire n_1306;
wire n_1961;
wire n_1413;
wire n_1783;
wire n_1759;
wire n_1266;
wire n_497;
wire n_911;
wire n_1904;
wire n_450;
wire n_1578;
wire n_473;
wire n_1779;
wire n_967;
wire n_1709;
wire n_474;
wire n_1159;
wire n_1908;
wire n_1315;
wire n_1055;
wire n_611;
wire n_380;
wire n_1576;
wire n_844;
wire n_1840;
wire n_968;
wire n_710;
wire n_1040;
wire n_1102;
wire n_661;
wire n_1185;
wire n_447;
wire n_1795;
wire n_403;
wire n_1039;
wire n_1119;
wire n_574;
wire n_1069;
wire n_1451;
wire n_842;
wire n_1788;
wire n_1938;
wire n_798;
wire n_1700;
wire n_668;
wire n_862;
wire n_869;
wire n_1816;
wire n_1952;
wire n_1811;
wire n_1066;
wire n_1917;
wire n_1377;
wire n_800;
wire n_1175;
wire n_778;
wire n_1170;
wire n_522;
wire n_1475;
wire n_1928;
wire n_943;
wire n_977;
wire n_905;
wire n_386;
wire n_878;
wire n_1734;
wire n_1333;
wire n_577;
wire n_1610;
wire n_759;
wire n_1235;
wire n_900;
wire n_841;
wire n_1724;
wire n_1218;
wire n_736;
wire n_1706;
wire n_766;
wire n_852;
wire n_1268;
wire n_1113;
wire n_1695;
wire n_1089;
wire n_1122;
wire n_908;
wire n_1123;
wire n_923;
wire n_1302;
wire n_1289;
wire n_937;
wire n_1442;
wire n_773;
wire n_1446;
wire n_1778;
wire n_865;
wire n_1644;
wire n_1736;
wire n_1932;
wire n_1707;
wire n_594;
wire n_856;
wire n_1146;
wire n_1685;
wire n_1810;
wire n_1435;
wire n_1800;
wire n_932;
wire n_958;
wire n_1755;
wire n_775;
wire n_763;
wire n_1093;
wire n_427;
wire n_1540;
wire n_519;
wire n_1878;
wire n_1116;
wire n_709;
wire n_1834;
wire n_388;
wire n_1913;
wire n_1899;
wire n_816;
wire n_1470;
wire n_625;
wire n_953;
wire n_1565;
wire n_1953;
wire n_1373;
wire n_1558;
wire n_716;
wire n_1683;
wire n_584;
wire n_896;
wire n_1817;
wire n_1722;
wire n_528;
wire n_1638;
wire n_1078;
wire n_495;
wire n_1072;
wire n_1663;
wire n_935;
wire n_1505;
wire n_467;
wire n_1213;
wire n_1053;
wire n_515;
wire n_1019;
wire n_680;
wire n_1180;
wire n_904;
wire n_920;
wire n_1117;
wire n_1923;
wire n_1168;
wire n_1598;
wire n_1309;
wire n_909;
wire n_523;
wire n_996;
wire n_439;
wire n_506;
wire n_606;
wire n_513;
wire n_1850;
wire n_1332;
wire n_1927;
wire n_1411;
wire n_1263;
wire n_1922;
wire n_1115;
wire n_725;
wire n_960;
wire n_671;
wire n_1084;
wire n_1726;
wire n_1827;
wire n_1656;
wire n_454;
wire n_1303;
wire n_1471;
wire n_443;
wire n_1949;
wire n_1029;
wire n_1207;
wire n_1555;
wire n_1962;
wire n_664;
wire n_1017;
wire n_1942;
wire n_581;
wire n_936;
wire n_1215;
wire n_582;
wire n_641;
wire n_1738;
wire n_940;
wire n_745;
wire n_1608;
wire n_1167;
wire n_1939;
wire n_1327;
wire n_609;
wire n_1743;
wire n_1752;
wire n_1792;
wire n_1006;
wire n_1869;
wire n_1259;
wire n_561;
wire n_437;
wire n_1560;
wire n_405;
wire n_1223;
wire n_621;
wire n_1012;
wire n_1241;
wire n_1671;
wire n_1414;
wire n_502;
wire n_769;
wire n_434;
wire n_1455;
wire n_1212;
wire n_1054;
wire n_1669;
wire n_1308;
wire n_1050;
wire n_426;
wire n_1550;
wire n_1134;
wire n_1895;
wire n_1670;
wire n_1941;
wire n_1319;
wire n_1363;
wire n_616;
wire n_880;
wire n_1103;
wire n_1274;
wire n_832;
wire n_1321;
wire n_1429;
wire n_1660;
wire n_1060;
wire n_1154;
wire n_1786;
wire n_632;
wire n_1344;
wire n_1450;
wire n_1603;
wire n_1720;
wire n_714;
wire n_1331;
wire n_1222;
wire n_1041;
wire n_1764;
wire n_1512;
wire n_957;
wire n_1255;
wire n_995;
wire n_1124;
wire n_1335;
wire n_1405;
wire n_1948;
wire n_912;
wire n_464;
wire n_1227;
wire n_1509;
wire n_945;
wire n_392;
wire n_563;
wire n_891;
wire n_568;
wire n_1586;
wire n_413;
wire n_1157;
wire n_902;
wire n_1749;
wire n_1158;
wire n_1886;
wire n_1079;
wire n_1330;
wire n_1033;
wire n_1464;
wire n_1028;
wire n_1832;
wire n_727;
wire n_1083;
wire n_397;
wire n_1056;
wire n_1592;
wire n_1605;
wire n_1802;
wire n_1855;
wire n_663;
wire n_588;
wire n_1682;
wire n_1698;
wire n_1448;
wire n_707;
wire n_915;
wire n_1774;
wire n_1785;
wire n_1001;
wire n_1418;
wire n_711;
wire n_864;
wire n_1782;
wire n_1169;
wire n_377;
wire n_1139;
wire n_1482;
wire n_1798;
wire n_1038;
wire n_1085;
wire n_845;
wire n_1838;
wire n_1673;
wire n_1619;
wire n_1127;
wire n_1718;
wire n_484;
wire n_893;
wire n_1068;
wire n_747;
wire n_1672;
wire n_1753;
wire n_1244;
wire n_1581;
wire n_1863;
wire n_697;
wire n_978;
wire n_847;
wire n_1452;
wire n_826;
wire n_628;
wire n_487;
wire n_831;
wire n_1772;
wire n_653;
wire n_1725;
wire n_692;
wire n_1433;
wire n_1051;
wire n_1696;
wire n_1355;
wire n_1494;
wire n_1517;
wire n_827;
wire n_472;
wire n_866;
wire n_452;
wire n_630;
wire n_820;
wire n_1208;
wire n_612;
wire n_1426;
wire n_858;
wire n_764;
wire n_741;
wire n_1090;
wire n_456;
wire n_1469;
wire n_1164;
wire n_433;
wire n_627;
wire n_1693;
wire n_1791;
wire n_418;
wire n_771;
wire n_1378;
wire n_524;
wire n_1496;
wire n_705;
wire n_1191;
wire n_1206;
wire n_1824;
wire n_1933;
wire n_1270;
wire n_1566;
wire n_1399;
wire n_546;
wire n_1010;
wire n_1375;
wire n_1015;
wire n_1761;
wire n_863;
wire n_525;
wire n_1226;
wire n_1617;
wire n_1790;
wire n_644;
wire n_1150;
wire n_1861;
wire n_1341;
wire n_833;
wire n_1229;
wire n_1690;
wire n_929;
wire n_1143;
wire n_1190;
wire n_1728;
wire n_543;
wire n_1710;
wire n_585;
wire n_1343;
wire n_719;
wire n_465;
wire n_1457;
wire n_1604;
wire n_1156;
wire n_988;
wire n_1757;
wire n_1466;
wire n_921;
wire n_1396;
wire n_1799;
wire n_1931;
wire n_640;
wire n_1176;
wire n_1691;
wire n_1721;
wire n_1511;
wire n_1151;
wire n_1501;
wire n_1254;
wire n_1458;
wire n_646;
wire n_650;
wire n_1211;
wire n_743;
wire n_823;
wire n_393;
wire n_1804;
wire n_1480;
wire n_1101;
wire n_1076;
wire n_1251;
wire n_1434;
wire n_1461;
wire n_1449;
wire n_1715;
wire n_1407;
wire n_1104;
wire n_1964;
wire n_849;
wire n_1061;
wire n_554;
wire n_1153;
wire n_1337;
wire n_797;
wire n_1704;
wire n_1844;
wire n_1177;
wire n_758;
wire n_436;
wire n_390;
wire n_1096;
wire n_1316;
wire n_1590;
wire n_1937;
wire n_1420;
wire n_1552;
wire n_1544;
wire n_1571;
wire n_1092;
wire n_1841;
wire n_846;
wire n_631;
wire n_673;
wire n_1410;
wire n_1067;
wire n_518;
wire n_1192;
wire n_1292;
wire n_1478;
wire n_1507;
wire n_1240;
wire n_1789;
wire n_987;
wire n_1596;
wire n_1065;
wire n_1064;
wire n_540;
wire n_1075;
wire n_1822;
wire n_718;
wire n_1955;
wire n_669;
wire n_1091;
wire n_423;
wire n_1969;
wire n_1221;
wire n_458;
wire n_1200;
wire n_444;
wire n_1777;
wire n_555;
wire n_1295;
wire n_974;
wire n_1329;
wire n_857;
wire n_1424;
wire n_1819;
wire n_1887;
wire n_1674;
wire n_491;
wire n_1294;
wire n_1902;
wire n_1110;
wire n_1137;
wire n_1533;
wire n_1889;
wire n_460;
wire n_1679;
wire n_1595;
wire n_1735;
wire n_666;
wire n_660;
wire n_1359;
wire n_886;
wire n_1896;
wire n_767;
wire n_889;
wire n_1398;
wire n_1911;
wire n_379;
wire n_1847;
wire n_1432;
wire n_1021;
wire n_1297;
wire n_1046;
wire n_1109;
wire n_961;
wire n_1447;
wire n_489;
wire n_1912;
wire n_1622;
wire n_1381;
wire n_1582;
wire n_1747;
wire n_573;
wire n_1654;
wire n_1099;
wire n_626;
wire n_539;
wire n_1919;
wire n_462;
wire n_615;
wire n_1118;
wire n_990;
wire n_1108;
wire n_670;
wire n_818;
wire n_918;
wire n_1272;
wire n_1541;
wire n_408;
wire n_1754;
wire n_892;
wire n_578;
wire n_938;
wire n_774;
wire n_466;
wire n_1584;
wire n_559;
wire n_1277;
wire n_1049;
wire n_1950;
wire n_984;
wire n_726;
wire n_517;
wire n_931;
wire n_780;
wire n_1851;
wire n_530;
wire n_834;
wire n_693;
wire n_496;
wire n_1257;
wire n_1082;
wire n_1360;
wire n_468;
wire n_1916;
wire n_532;
wire n_1025;
wire n_1875;
wire n_1826;
wire n_1836;
wire n_1909;
wire n_924;
wire n_1264;
wire n_1858;
wire n_1527;
wire n_1245;
wire n_1152;
wire n_1539;
wire n_1901;
wire n_1081;
wire n_547;
wire n_1324;
wire n_1198;
wire n_1678;
wire n_1943;
wire n_1307;
wire n_993;
wire n_819;
wire n_737;
wire n_1489;
wire n_1637;
wire n_1318;
wire n_1290;
wire n_1063;
wire n_1135;
wire n_828;
wire n_770;
wire n_867;
wire n_398;
wire n_1100;
wire n_1519;
wire n_425;
wire n_1650;
wire n_879;
wire n_1640;
wire n_449;
wire n_1340;
wire n_1562;
wire n_607;
wire n_629;
wire n_706;
wire n_901;
wire n_876;
wire n_1443;
wire n_1818;
wire n_655;
wire n_654;
wire n_1521;
wire n_672;
wire n_567;
wire n_916;
wire n_1354;
wire n_1780;
wire n_1547;
wire n_1823;
wire n_1867;
wire n_1334;
wire n_1291;
wire n_1437;
wire n_1473;
wire n_986;
wire n_451;
wire n_1037;
wire n_1891;
wire n_1267;
wire n_790;
wire n_1262;
wire n_1843;
wire n_410;
wire n_1684;
wire n_1444;
wire n_751;
wire n_999;
wire n_913;
wire n_1237;
wire n_1506;
wire n_1885;
wire n_1356;
wire n_1646;
wire n_768;
wire n_412;
wire n_542;
wire n_1256;
wire n_1427;
wire n_1077;
wire n_1111;
wire n_1503;
wire n_1249;
wire n_1416;
wire n_387;
wire n_1239;
wire n_1796;
wire n_1662;
wire n_1963;
wire n_1958;
wire n_969;
wire n_1535;
wire n_1009;
wire n_1202;
wire n_1498;
wire n_1925;
wire n_1801;
wire n_1549;
wire n_604;
wire n_848;
wire n_756;
wire n_713;
wire n_598;
wire n_1968;
wire n_1252;
wire n_1647;
wire n_430;
wire n_1132;
wire n_1947;
wire n_1649;
wire n_1275;
wire n_843;
wire n_579;
wire n_533;
wire n_1472;
wire n_385;
wire n_536;
wire n_470;
wire n_851;
wire n_1155;
wire n_934;
wire n_1636;
wire n_1027;
wire n_965;
wire n_1894;
wire n_1296;
wire n_382;
wire n_1484;
wire n_1043;
wire n_435;
wire n_511;
wire n_1808;
wire n_1492;
wire n_1467;
wire n_509;
wire n_1204;
wire n_930;
wire n_1265;
wire n_1057;
wire n_1481;
wire n_907;
wire n_1430;
wire n_1758;
wire n_1005;
wire n_1312;
wire n_1697;
wire n_1877;
wire n_1900;
wire n_899;
wire n_637;
wire n_544;
wire n_1476;
wire n_1087;
wire n_1842;
wire n_1536;
wire n_1746;
wire n_1898;
wire n_1711;
wire n_482;
wire n_633;
wire n_1892;
wire n_971;
wire n_1052;
wire n_1071;
wire n_1311;
wire n_1601;
wire n_1438;
wire n_1273;
wire n_959;
wire n_1573;
wire n_1130;
wire n_1918;
wire n_794;
wire n_1228;
wire n_681;
wire n_982;
wire n_717;
wire n_1624;
wire n_1253;
wire n_1183;
wire n_1831;
wire n_516;
wire n_1460;
wire n_521;
wire n_1195;
wire n_575;
wire n_1300;
wire n_1372;
wire n_698;
wire n_1345;
wire n_587;
wire n_1701;
wire n_1664;
wire n_1428;
wire n_1246;
wire n_1074;
wire n_674;
wire n_888;
wire n_1546;
wire n_1436;
wire n_793;
wire n_1390;
wire n_1815;
wire n_1924;
wire n_1412;
wire n_1868;
wire n_757;
wire n_1534;
wire n_803;
wire n_514;
wire n_507;
wire n_1557;
wire n_614;
wire n_772;
wire n_1114;
wire n_566;
wire n_871;
wire n_1739;
wire n_1088;
wire n_1230;
wire n_1326;
wire n_1402;
wire n_1388;
wire n_483;
wire n_1630;
wire n_394;
wire n_729;
wire n_1280;
wire n_1323;
wire n_1352;
wire n_1097;
wire n_703;
wire n_1369;
wire n_601;
wire n_463;
wire n_396;
wire n_1236;
wire n_1523;
wire n_1528;
wire n_603;
wire n_1692;
wire n_1288;
wire n_868;
wire n_1705;
wire n_1024;
wire n_1144;
wire n_1627;
wire n_475;
wire n_897;
wire n_1320;
wire n_855;
wire n_1935;
wire n_1645;
wire n_429;
INVx1_ASAP7_75t_L g1624 ( .A(n_0), .Y(n_1624) );
AOI22xp33_ASAP7_75t_L g1717 ( .A1(n_1), .A2(n_106), .B1(n_1674), .B2(n_1677), .Y(n_1717) );
INVx1_ASAP7_75t_L g389 ( .A(n_2), .Y(n_389) );
NOR2xp33_ASAP7_75t_L g470 ( .A(n_2), .B(n_399), .Y(n_470) );
AND2x2_ASAP7_75t_L g907 ( .A(n_2), .B(n_551), .Y(n_907) );
AND2x2_ASAP7_75t_L g964 ( .A(n_2), .B(n_272), .Y(n_964) );
INVx1_ASAP7_75t_L g871 ( .A(n_3), .Y(n_871) );
INVx1_ASAP7_75t_L g689 ( .A(n_4), .Y(n_689) );
OAI22xp5_ASAP7_75t_L g1625 ( .A1(n_5), .A2(n_283), .B1(n_1626), .B2(n_1627), .Y(n_1625) );
OAI211xp5_ASAP7_75t_L g1629 ( .A1(n_5), .A2(n_1630), .B(n_1632), .C(n_1638), .Y(n_1629) );
INVx1_ASAP7_75t_L g1289 ( .A(n_6), .Y(n_1289) );
INVx1_ASAP7_75t_L g1395 ( .A(n_7), .Y(n_1395) );
OAI22xp5_ASAP7_75t_L g1477 ( .A1(n_8), .A2(n_159), .B1(n_555), .B2(n_1478), .Y(n_1477) );
OAI22xp5_ASAP7_75t_L g1490 ( .A1(n_8), .A2(n_159), .B1(n_512), .B2(n_803), .Y(n_1490) );
OAI22xp5_ASAP7_75t_L g1907 ( .A1(n_9), .A2(n_290), .B1(n_1026), .B2(n_1442), .Y(n_1907) );
OAI22xp33_ASAP7_75t_L g1914 ( .A1(n_9), .A2(n_290), .B1(n_512), .B2(n_1067), .Y(n_1914) );
OAI22xp33_ASAP7_75t_L g1934 ( .A1(n_10), .A2(n_305), .B1(n_763), .B2(n_1935), .Y(n_1934) );
OAI22xp33_ASAP7_75t_L g1941 ( .A1(n_10), .A2(n_305), .B1(n_705), .B2(n_1942), .Y(n_1941) );
OAI22xp33_ASAP7_75t_L g1479 ( .A1(n_11), .A2(n_298), .B1(n_391), .B2(n_548), .Y(n_1479) );
OAI22xp33_ASAP7_75t_L g1485 ( .A1(n_11), .A2(n_298), .B1(n_534), .B2(n_630), .Y(n_1485) );
OAI211xp5_ASAP7_75t_L g685 ( .A1(n_12), .A2(n_518), .B(n_686), .C(n_687), .Y(n_685) );
INVx1_ASAP7_75t_L g702 ( .A(n_12), .Y(n_702) );
INVx1_ASAP7_75t_L g717 ( .A(n_13), .Y(n_717) );
AOI22xp33_ASAP7_75t_L g1587 ( .A1(n_14), .A2(n_79), .B1(n_742), .B2(n_1296), .Y(n_1587) );
AOI22xp33_ASAP7_75t_L g1600 ( .A1(n_14), .A2(n_240), .B1(n_1356), .B2(n_1368), .Y(n_1600) );
AOI22xp33_ASAP7_75t_L g1285 ( .A1(n_15), .A2(n_83), .B1(n_1286), .B2(n_1287), .Y(n_1285) );
AOI221xp5_ASAP7_75t_L g1307 ( .A1(n_15), .A2(n_25), .B1(n_954), .B2(n_1308), .C(n_1310), .Y(n_1307) );
INVx1_ASAP7_75t_L g418 ( .A(n_16), .Y(n_418) );
OAI22xp5_ASAP7_75t_L g752 ( .A1(n_17), .A2(n_50), .B1(n_682), .B2(n_753), .Y(n_752) );
OAI22xp5_ASAP7_75t_L g768 ( .A1(n_17), .A2(n_50), .B1(n_548), .B2(n_769), .Y(n_768) );
AOI22xp33_ASAP7_75t_L g1615 ( .A1(n_18), .A2(n_320), .B1(n_742), .B2(n_1270), .Y(n_1615) );
AOI22xp33_ASAP7_75t_L g1642 ( .A1(n_18), .A2(n_367), .B1(n_954), .B2(n_1643), .Y(n_1642) );
AOI22xp33_ASAP7_75t_L g1174 ( .A1(n_19), .A2(n_31), .B1(n_1141), .B2(n_1175), .Y(n_1174) );
INVx1_ASAP7_75t_L g1216 ( .A(n_19), .Y(n_1216) );
OAI211xp5_ASAP7_75t_L g1543 ( .A1(n_20), .A2(n_619), .B(n_757), .C(n_1544), .Y(n_1543) );
INVx1_ASAP7_75t_L g1551 ( .A(n_20), .Y(n_1551) );
INVx1_ASAP7_75t_L g1425 ( .A(n_21), .Y(n_1425) );
OAI211xp5_ASAP7_75t_L g1430 ( .A1(n_21), .A2(n_757), .B(n_1431), .C(n_1432), .Y(n_1430) );
INVx1_ASAP7_75t_L g1341 ( .A(n_22), .Y(n_1341) );
OAI22xp33_ASAP7_75t_L g628 ( .A1(n_23), .A2(n_179), .B1(n_629), .B2(n_630), .Y(n_628) );
OAI22xp33_ASAP7_75t_L g633 ( .A1(n_23), .A2(n_179), .B1(n_391), .B2(n_634), .Y(n_633) );
INVx1_ASAP7_75t_L g1398 ( .A(n_24), .Y(n_1398) );
AOI22xp33_ASAP7_75t_SL g1298 ( .A1(n_25), .A2(n_255), .B1(n_1175), .B2(n_1299), .Y(n_1298) );
INVx1_ASAP7_75t_L g1905 ( .A(n_26), .Y(n_1905) );
INVx1_ASAP7_75t_L g1530 ( .A(n_27), .Y(n_1530) );
INVx2_ASAP7_75t_L g416 ( .A(n_28), .Y(n_416) );
INVx1_ASAP7_75t_L g1880 ( .A(n_29), .Y(n_1880) );
OAI211xp5_ASAP7_75t_L g1903 ( .A1(n_30), .A2(n_792), .B(n_1253), .C(n_1904), .Y(n_1903) );
INVx1_ASAP7_75t_L g1913 ( .A(n_30), .Y(n_1913) );
AOI221xp5_ASAP7_75t_L g1195 ( .A1(n_31), .A2(n_49), .B1(n_1196), .B2(n_1198), .C(n_1199), .Y(n_1195) );
INVx1_ASAP7_75t_L g1956 ( .A(n_32), .Y(n_1956) );
INVx1_ASAP7_75t_L g1293 ( .A(n_33), .Y(n_1293) );
INVx1_ASAP7_75t_L g457 ( .A(n_34), .Y(n_457) );
OAI22xp5_ASAP7_75t_L g880 ( .A1(n_35), .A2(n_312), .B1(n_534), .B2(n_626), .Y(n_880) );
OAI22xp5_ASAP7_75t_L g888 ( .A1(n_35), .A2(n_343), .B1(n_555), .B2(n_558), .Y(n_888) );
INVx1_ASAP7_75t_L g1569 ( .A(n_36), .Y(n_1569) );
INVx1_ASAP7_75t_L g1406 ( .A(n_37), .Y(n_1406) );
OA222x2_ASAP7_75t_L g1077 ( .A1(n_38), .A2(n_90), .B1(n_266), .B2(n_1078), .C1(n_1082), .C2(n_1086), .Y(n_1077) );
INVx1_ASAP7_75t_L g1139 ( .A(n_38), .Y(n_1139) );
HB1xp67_ASAP7_75t_L g384 ( .A(n_39), .Y(n_384) );
AND2x2_ASAP7_75t_L g1668 ( .A(n_39), .B(n_382), .Y(n_1668) );
INVx1_ASAP7_75t_L g1889 ( .A(n_40), .Y(n_1889) );
INVx1_ASAP7_75t_L g1459 ( .A(n_41), .Y(n_1459) );
AOI22xp33_ASAP7_75t_L g1238 ( .A1(n_42), .A2(n_348), .B1(n_955), .B2(n_1239), .Y(n_1238) );
INVxp67_ASAP7_75t_SL g1258 ( .A(n_42), .Y(n_1258) );
AOI22xp33_ASAP7_75t_L g1176 ( .A1(n_43), .A2(n_234), .B1(n_742), .B2(n_998), .Y(n_1176) );
INVx1_ASAP7_75t_L g1201 ( .A(n_43), .Y(n_1201) );
INVx1_ASAP7_75t_L g718 ( .A(n_44), .Y(n_718) );
OAI22xp5_ASAP7_75t_L g1344 ( .A1(n_45), .A2(n_295), .B1(n_547), .B2(n_548), .Y(n_1344) );
OAI22xp5_ASAP7_75t_L g1349 ( .A1(n_45), .A2(n_202), .B1(n_534), .B2(n_763), .Y(n_1349) );
XNOR2xp5_ASAP7_75t_L g1519 ( .A(n_46), .B(n_1520), .Y(n_1519) );
AOI22xp33_ASAP7_75t_L g1716 ( .A1(n_46), .A2(n_87), .B1(n_1667), .B2(n_1671), .Y(n_1716) );
OAI22xp33_ASAP7_75t_L g1928 ( .A1(n_47), .A2(n_201), .B1(n_684), .B2(n_1060), .Y(n_1928) );
OAI22xp33_ASAP7_75t_L g1943 ( .A1(n_47), .A2(n_201), .B1(n_391), .B2(n_800), .Y(n_1943) );
INVx1_ASAP7_75t_L g1030 ( .A(n_48), .Y(n_1030) );
AOI22xp33_ASAP7_75t_SL g1181 ( .A1(n_49), .A2(n_339), .B1(n_1175), .B2(n_1182), .Y(n_1181) );
INVxp67_ASAP7_75t_SL g1292 ( .A(n_51), .Y(n_1292) );
OAI22xp5_ASAP7_75t_L g1315 ( .A1(n_51), .A2(n_190), .B1(n_679), .B2(n_1316), .Y(n_1315) );
AOI22xp33_ASAP7_75t_SL g1352 ( .A1(n_52), .A2(n_135), .B1(n_1353), .B2(n_1354), .Y(n_1352) );
AOI22xp33_ASAP7_75t_SL g1380 ( .A1(n_52), .A2(n_271), .B1(n_1260), .B2(n_1375), .Y(n_1380) );
INVx1_ASAP7_75t_L g645 ( .A(n_53), .Y(n_645) );
INVx1_ASAP7_75t_L g447 ( .A(n_54), .Y(n_447) );
INVx1_ASAP7_75t_L g1036 ( .A(n_55), .Y(n_1036) );
INVx1_ASAP7_75t_L g596 ( .A(n_56), .Y(n_596) );
OAI211xp5_ASAP7_75t_L g789 ( .A1(n_57), .A2(n_790), .B(n_792), .C(n_793), .Y(n_789) );
INVx1_ASAP7_75t_L g807 ( .A(n_57), .Y(n_807) );
CKINVDCx5p33_ASAP7_75t_R g1106 ( .A(n_58), .Y(n_1106) );
INVx1_ASAP7_75t_L g1303 ( .A(n_59), .Y(n_1303) );
INVx1_ASAP7_75t_L g864 ( .A(n_60), .Y(n_864) );
INVx1_ASAP7_75t_L g623 ( .A(n_61), .Y(n_623) );
AOI22xp33_ASAP7_75t_SL g1244 ( .A1(n_62), .A2(n_282), .B1(n_955), .B2(n_1245), .Y(n_1244) );
AOI22xp33_ASAP7_75t_L g1259 ( .A1(n_62), .A2(n_259), .B1(n_1130), .B2(n_1260), .Y(n_1259) );
OAI22xp33_ASAP7_75t_L g691 ( .A1(n_63), .A2(n_150), .B1(n_509), .B2(n_692), .Y(n_691) );
OAI22xp5_ASAP7_75t_L g703 ( .A1(n_63), .A2(n_150), .B1(n_704), .B2(n_705), .Y(n_703) );
CKINVDCx5p33_ASAP7_75t_R g1291 ( .A(n_64), .Y(n_1291) );
INVx1_ASAP7_75t_L g1326 ( .A(n_65), .Y(n_1326) );
BUFx6f_ASAP7_75t_L g396 ( .A(n_66), .Y(n_396) );
AOI22xp33_ASAP7_75t_L g1177 ( .A1(n_67), .A2(n_80), .B1(n_1178), .B2(n_1180), .Y(n_1177) );
INVx1_ASAP7_75t_L g1200 ( .A(n_67), .Y(n_1200) );
INVx1_ASAP7_75t_L g592 ( .A(n_68), .Y(n_592) );
INVx1_ASAP7_75t_L g821 ( .A(n_69), .Y(n_821) );
OAI22xp33_ASAP7_75t_SL g1234 ( .A1(n_70), .A2(n_268), .B1(n_494), .B2(n_1105), .Y(n_1234) );
INVx1_ASAP7_75t_L g1274 ( .A(n_70), .Y(n_1274) );
XNOR2xp5_ASAP7_75t_L g405 ( .A(n_71), .B(n_406), .Y(n_405) );
INVx1_ASAP7_75t_L g1462 ( .A(n_72), .Y(n_1462) );
INVx1_ASAP7_75t_L g1495 ( .A(n_73), .Y(n_1495) );
AOI21xp33_ASAP7_75t_L g967 ( .A1(n_74), .A2(n_968), .B(n_969), .Y(n_967) );
AOI221xp5_ASAP7_75t_L g1004 ( .A1(n_74), .A2(n_292), .B1(n_998), .B2(n_1005), .C(n_1007), .Y(n_1004) );
CKINVDCx5p33_ASAP7_75t_R g1166 ( .A(n_75), .Y(n_1166) );
AOI22xp5_ASAP7_75t_L g1692 ( .A1(n_76), .A2(n_122), .B1(n_1667), .B2(n_1671), .Y(n_1692) );
AOI22xp5_ASAP7_75t_L g1682 ( .A1(n_77), .A2(n_276), .B1(n_1667), .B2(n_1671), .Y(n_1682) );
OAI222xp33_ASAP7_75t_L g900 ( .A1(n_78), .A2(n_88), .B1(n_95), .B2(n_901), .C1(n_915), .C2(n_924), .Y(n_900) );
AOI22xp33_ASAP7_75t_SL g1597 ( .A1(n_79), .A2(n_114), .B1(n_1363), .B2(n_1598), .Y(n_1597) );
INVx1_ASAP7_75t_L g1220 ( .A(n_80), .Y(n_1220) );
INVx1_ASAP7_75t_L g532 ( .A(n_81), .Y(n_532) );
OAI211xp5_ASAP7_75t_L g563 ( .A1(n_81), .A2(n_564), .B(n_568), .C(n_573), .Y(n_563) );
OAI22xp33_ASAP7_75t_L g1606 ( .A1(n_82), .A2(n_327), .B1(n_910), .B2(n_1607), .Y(n_1606) );
INVx1_ASAP7_75t_L g1633 ( .A(n_82), .Y(n_1633) );
INVx1_ASAP7_75t_L g1325 ( .A(n_83), .Y(n_1325) );
INVx1_ASAP7_75t_L g868 ( .A(n_84), .Y(n_868) );
OAI22xp33_ASAP7_75t_L g1025 ( .A1(n_85), .A2(n_89), .B1(n_781), .B2(n_1026), .Y(n_1025) );
OAI22xp33_ASAP7_75t_L g1066 ( .A1(n_85), .A2(n_89), .B1(n_512), .B2(n_1067), .Y(n_1066) );
CKINVDCx5p33_ASAP7_75t_R g939 ( .A(n_86), .Y(n_939) );
OAI221xp5_ASAP7_75t_L g1123 ( .A1(n_90), .A2(n_215), .B1(n_1124), .B2(n_1126), .C(n_1128), .Y(n_1123) );
OAI22xp5_ASAP7_75t_L g1209 ( .A1(n_91), .A2(n_324), .B1(n_478), .B2(n_679), .Y(n_1209) );
INVx1_ASAP7_75t_L g1222 ( .A(n_91), .Y(n_1222) );
INVx1_ASAP7_75t_L g1096 ( .A(n_92), .Y(n_1096) );
AOI22xp33_ASAP7_75t_L g1157 ( .A1(n_92), .A2(n_146), .B1(n_999), .B2(n_1158), .Y(n_1157) );
INVx1_ASAP7_75t_L g1045 ( .A(n_93), .Y(n_1045) );
XOR2x2_ASAP7_75t_L g1434 ( .A(n_94), .B(n_1435), .Y(n_1434) );
AOI22xp33_ASAP7_75t_L g1704 ( .A1(n_94), .A2(n_263), .B1(n_1667), .B2(n_1671), .Y(n_1704) );
OAI22xp5_ASAP7_75t_L g983 ( .A1(n_95), .A2(n_371), .B1(n_984), .B2(n_988), .Y(n_983) );
INVx1_ASAP7_75t_L g1957 ( .A(n_96), .Y(n_1957) );
AOI22xp5_ASAP7_75t_L g1686 ( .A1(n_97), .A2(n_270), .B1(n_1674), .B2(n_1677), .Y(n_1686) );
AOI22xp5_ASAP7_75t_L g1687 ( .A1(n_98), .A2(n_115), .B1(n_1667), .B2(n_1688), .Y(n_1687) );
INVx1_ASAP7_75t_L g1568 ( .A(n_99), .Y(n_1568) );
AO22x1_ASAP7_75t_L g1710 ( .A1(n_100), .A2(n_277), .B1(n_1674), .B2(n_1677), .Y(n_1710) );
AOI22xp33_ASAP7_75t_SL g1589 ( .A1(n_101), .A2(n_188), .B1(n_1175), .B2(n_1373), .Y(n_1589) );
AOI22xp33_ASAP7_75t_L g1594 ( .A1(n_101), .A2(n_247), .B1(n_1356), .B2(n_1595), .Y(n_1594) );
INVx1_ASAP7_75t_L g1439 ( .A(n_102), .Y(n_1439) );
XOR2x2_ASAP7_75t_L g849 ( .A(n_103), .B(n_850), .Y(n_849) );
AOI22xp33_ASAP7_75t_L g971 ( .A1(n_104), .A2(n_177), .B1(n_972), .B2(n_974), .Y(n_971) );
INVx1_ASAP7_75t_L g1001 ( .A(n_104), .Y(n_1001) );
INVx1_ASAP7_75t_L g442 ( .A(n_105), .Y(n_442) );
XNOR2xp5_ASAP7_75t_L g640 ( .A(n_107), .B(n_641), .Y(n_640) );
CKINVDCx5p33_ASAP7_75t_R g1302 ( .A(n_108), .Y(n_1302) );
AOI22xp33_ASAP7_75t_SL g1616 ( .A1(n_109), .A2(n_275), .B1(n_1158), .B2(n_1265), .Y(n_1616) );
AOI221xp5_ASAP7_75t_L g1639 ( .A1(n_109), .A2(n_329), .B1(n_1342), .B2(n_1640), .C(n_1641), .Y(n_1639) );
AOI22xp33_ASAP7_75t_L g1295 ( .A1(n_110), .A2(n_344), .B1(n_1178), .B2(n_1296), .Y(n_1295) );
AOI221xp5_ASAP7_75t_L g1322 ( .A1(n_110), .A2(n_230), .B1(n_955), .B2(n_1198), .C(n_1323), .Y(n_1322) );
OAI211xp5_ASAP7_75t_L g1480 ( .A1(n_111), .A2(n_790), .B(n_792), .C(n_1481), .Y(n_1480) );
INVx1_ASAP7_75t_L g1489 ( .A(n_111), .Y(n_1489) );
INVx1_ASAP7_75t_L g652 ( .A(n_112), .Y(n_652) );
INVx1_ASAP7_75t_L g593 ( .A(n_113), .Y(n_593) );
AOI22xp33_ASAP7_75t_L g1586 ( .A1(n_114), .A2(n_240), .B1(n_742), .B2(n_1296), .Y(n_1586) );
INVx1_ASAP7_75t_L g1224 ( .A(n_115), .Y(n_1224) );
OAI22xp5_ASAP7_75t_L g1023 ( .A1(n_116), .A2(n_158), .B1(n_548), .B2(n_1024), .Y(n_1023) );
OAI22xp5_ASAP7_75t_L g1059 ( .A1(n_116), .A2(n_158), .B1(n_1060), .B2(n_1062), .Y(n_1059) );
OAI22xp33_ASAP7_75t_L g1420 ( .A1(n_117), .A2(n_121), .B1(n_634), .B2(n_771), .Y(n_1420) );
OAI22xp33_ASAP7_75t_L g1428 ( .A1(n_117), .A2(n_121), .B1(n_537), .B2(n_1060), .Y(n_1428) );
OAI22xp5_ASAP7_75t_L g1547 ( .A1(n_118), .A2(n_199), .B1(n_512), .B2(n_684), .Y(n_1547) );
OAI22xp5_ASAP7_75t_L g1552 ( .A1(n_118), .A2(n_239), .B1(n_704), .B2(n_1553), .Y(n_1552) );
INVx1_ASAP7_75t_L g382 ( .A(n_119), .Y(n_382) );
INVx1_ASAP7_75t_L g434 ( .A(n_120), .Y(n_434) );
INVx1_ASAP7_75t_L g1527 ( .A(n_123), .Y(n_1527) );
AO221x2_ASAP7_75t_L g1777 ( .A1(n_124), .A2(n_359), .B1(n_1674), .B2(n_1677), .C(n_1778), .Y(n_1777) );
INVx1_ASAP7_75t_L g854 ( .A(n_125), .Y(n_854) );
OAI211xp5_ASAP7_75t_L g1437 ( .A1(n_126), .A2(n_792), .B(n_1253), .C(n_1438), .Y(n_1437) );
INVx1_ASAP7_75t_L g1449 ( .A(n_126), .Y(n_1449) );
OAI22xp5_ASAP7_75t_L g796 ( .A1(n_127), .A2(n_373), .B1(n_555), .B2(n_797), .Y(n_796) );
OAI22xp5_ASAP7_75t_L g802 ( .A1(n_127), .A2(n_133), .B1(n_534), .B2(n_803), .Y(n_802) );
INVx1_ASAP7_75t_L g1883 ( .A(n_128), .Y(n_1883) );
INVx1_ASAP7_75t_L g1483 ( .A(n_129), .Y(n_1483) );
OAI211xp5_ASAP7_75t_L g1486 ( .A1(n_129), .A2(n_518), .B(n_1487), .C(n_1488), .Y(n_1486) );
XOR2xp5_ASAP7_75t_L g1924 ( .A(n_130), .B(n_1925), .Y(n_1924) );
OAI22xp5_ASAP7_75t_L g1233 ( .A1(n_131), .A2(n_164), .B1(n_719), .B2(n_1097), .Y(n_1233) );
NOR2xp33_ASAP7_75t_L g1278 ( .A(n_131), .B(n_803), .Y(n_1278) );
CKINVDCx5p33_ASAP7_75t_R g1191 ( .A(n_132), .Y(n_1191) );
OAI22xp33_ASAP7_75t_L g799 ( .A1(n_133), .A2(n_342), .B1(n_391), .B2(n_800), .Y(n_799) );
INVx1_ASAP7_75t_L g1465 ( .A(n_134), .Y(n_1465) );
AOI22xp33_ASAP7_75t_L g1370 ( .A1(n_135), .A2(n_250), .B1(n_1371), .B2(n_1373), .Y(n_1370) );
OAI22xp5_ASAP7_75t_L g1426 ( .A1(n_136), .A2(n_315), .B1(n_704), .B2(n_797), .Y(n_1426) );
OAI22xp5_ASAP7_75t_L g1429 ( .A1(n_136), .A2(n_315), .B1(n_692), .B2(n_1067), .Y(n_1429) );
AOI22xp33_ASAP7_75t_L g1613 ( .A1(n_137), .A2(n_367), .B1(n_742), .B2(n_1614), .Y(n_1613) );
AOI21xp33_ASAP7_75t_L g1651 ( .A1(n_137), .A2(n_1652), .B(n_1653), .Y(n_1651) );
INVx1_ASAP7_75t_L g1953 ( .A(n_138), .Y(n_1953) );
INVx1_ASAP7_75t_L g1424 ( .A(n_139), .Y(n_1424) );
OAI22xp5_ASAP7_75t_L g885 ( .A1(n_140), .A2(n_343), .B1(n_512), .B2(n_809), .Y(n_885) );
OAI22xp33_ASAP7_75t_L g887 ( .A1(n_140), .A2(n_312), .B1(n_391), .B2(n_634), .Y(n_887) );
INVx1_ASAP7_75t_L g1388 ( .A(n_141), .Y(n_1388) );
INVx1_ASAP7_75t_L g595 ( .A(n_142), .Y(n_595) );
INVx1_ASAP7_75t_L g1566 ( .A(n_143), .Y(n_1566) );
INVx1_ASAP7_75t_L g761 ( .A(n_144), .Y(n_761) );
OAI211xp5_ASAP7_75t_L g772 ( .A1(n_144), .A2(n_773), .B(n_774), .C(n_778), .Y(n_772) );
OAI211xp5_ASAP7_75t_L g618 ( .A1(n_145), .A2(n_518), .B(n_619), .C(n_622), .Y(n_618) );
INVx1_ASAP7_75t_L g638 ( .A(n_145), .Y(n_638) );
AOI22xp33_ASAP7_75t_L g1107 ( .A1(n_146), .A2(n_197), .B1(n_986), .B2(n_1108), .Y(n_1107) );
OAI22xp33_ASAP7_75t_L g1908 ( .A1(n_147), .A2(n_347), .B1(n_548), .B2(n_1024), .Y(n_1908) );
OAI22xp5_ASAP7_75t_L g1910 ( .A1(n_147), .A2(n_347), .B1(n_536), .B2(n_1062), .Y(n_1910) );
OAI22xp5_ASAP7_75t_L g1441 ( .A1(n_148), .A2(n_355), .B1(n_704), .B2(n_1442), .Y(n_1441) );
OAI22xp5_ASAP7_75t_L g1445 ( .A1(n_148), .A2(n_355), .B1(n_764), .B2(n_803), .Y(n_1445) );
INVx1_ASAP7_75t_L g606 ( .A(n_149), .Y(n_606) );
OAI22xp5_ASAP7_75t_L g1113 ( .A1(n_151), .A2(n_215), .B1(n_1114), .B2(n_1117), .Y(n_1113) );
INVx1_ASAP7_75t_L g1140 ( .A(n_151), .Y(n_1140) );
INVx1_ASAP7_75t_L g725 ( .A(n_152), .Y(n_725) );
OAI22xp33_ASAP7_75t_L g1443 ( .A1(n_153), .A2(n_204), .B1(n_634), .B2(n_771), .Y(n_1443) );
OAI22xp33_ASAP7_75t_L g1450 ( .A1(n_153), .A2(n_204), .B1(n_536), .B2(n_537), .Y(n_1450) );
AO22x1_ASAP7_75t_L g1673 ( .A1(n_154), .A2(n_363), .B1(n_1674), .B2(n_1677), .Y(n_1673) );
INVx1_ASAP7_75t_L g1039 ( .A(n_155), .Y(n_1039) );
INVx1_ASAP7_75t_L g1534 ( .A(n_156), .Y(n_1534) );
INVx1_ASAP7_75t_L g1620 ( .A(n_157), .Y(n_1620) );
OAI221xp5_ASAP7_75t_L g1645 ( .A1(n_157), .A2(n_217), .B1(n_1646), .B2(n_1647), .C(n_1649), .Y(n_1645) );
OAI221xp5_ASAP7_75t_L g1248 ( .A1(n_160), .A2(n_350), .B1(n_1249), .B2(n_1252), .C(n_1253), .Y(n_1248) );
INVx1_ASAP7_75t_L g1271 ( .A(n_160), .Y(n_1271) );
INVx1_ASAP7_75t_L g1236 ( .A(n_161), .Y(n_1236) );
AOI22xp33_ASAP7_75t_L g1264 ( .A1(n_161), .A2(n_282), .B1(n_1130), .B2(n_1265), .Y(n_1264) );
INVx1_ASAP7_75t_L g666 ( .A(n_162), .Y(n_666) );
CKINVDCx5p33_ASAP7_75t_R g1241 ( .A(n_163), .Y(n_1241) );
INVx1_ASAP7_75t_L g1273 ( .A(n_164), .Y(n_1273) );
INVx1_ASAP7_75t_L g659 ( .A(n_165), .Y(n_659) );
INVx1_ASAP7_75t_L g1339 ( .A(n_166), .Y(n_1339) );
OAI211xp5_ASAP7_75t_L g1347 ( .A1(n_166), .A2(n_518), .B(n_805), .C(n_1348), .Y(n_1347) );
INVx1_ASAP7_75t_L g1933 ( .A(n_167), .Y(n_1933) );
OAI211xp5_ASAP7_75t_L g1938 ( .A1(n_167), .A2(n_566), .B(n_697), .C(n_1939), .Y(n_1938) );
OAI211xp5_ASAP7_75t_L g881 ( .A1(n_168), .A2(n_757), .B(n_805), .C(n_882), .Y(n_881) );
INVx1_ASAP7_75t_L g894 ( .A(n_168), .Y(n_894) );
INVx1_ASAP7_75t_L g1546 ( .A(n_169), .Y(n_1546) );
OAI211xp5_ASAP7_75t_SL g1549 ( .A1(n_169), .A2(n_792), .B(n_890), .C(n_1550), .Y(n_1549) );
OAI22xp33_ASAP7_75t_L g533 ( .A1(n_170), .A2(n_278), .B1(n_534), .B2(n_537), .Y(n_533) );
OAI22xp5_ASAP7_75t_L g546 ( .A1(n_170), .A2(n_278), .B1(n_547), .B2(n_548), .Y(n_546) );
INVx1_ASAP7_75t_L g1402 ( .A(n_171), .Y(n_1402) );
OAI22xp5_ASAP7_75t_L g1542 ( .A1(n_172), .A2(n_239), .B1(n_534), .B2(n_626), .Y(n_1542) );
OAI22xp33_ASAP7_75t_L g1554 ( .A1(n_172), .A2(n_199), .B1(n_391), .B2(n_634), .Y(n_1554) );
INVx1_ASAP7_75t_L g1482 ( .A(n_173), .Y(n_1482) );
INVx1_ASAP7_75t_L g426 ( .A(n_174), .Y(n_426) );
INVx1_ASAP7_75t_L g1951 ( .A(n_175), .Y(n_1951) );
INVx1_ASAP7_75t_L g451 ( .A(n_176), .Y(n_451) );
INVxp67_ASAP7_75t_SL g1008 ( .A(n_177), .Y(n_1008) );
INVx1_ASAP7_75t_L g601 ( .A(n_178), .Y(n_601) );
INVx1_ASAP7_75t_L g661 ( .A(n_180), .Y(n_661) );
OAI22xp33_ASAP7_75t_L g681 ( .A1(n_181), .A2(n_358), .B1(n_682), .B2(n_684), .Y(n_681) );
OAI22xp33_ASAP7_75t_L g695 ( .A1(n_181), .A2(n_358), .B1(n_391), .B2(n_634), .Y(n_695) );
OAI22xp33_ASAP7_75t_L g508 ( .A1(n_182), .A2(n_212), .B1(n_509), .B2(n_512), .Y(n_508) );
OAI22xp33_ASAP7_75t_L g554 ( .A1(n_182), .A2(n_212), .B1(n_555), .B2(n_558), .Y(n_554) );
OAI211xp5_ASAP7_75t_L g1421 ( .A1(n_183), .A2(n_773), .B(n_1422), .C(n_1423), .Y(n_1421) );
INVx1_ASAP7_75t_L g1433 ( .A(n_183), .Y(n_1433) );
XNOR2xp5_ASAP7_75t_L g1560 ( .A(n_184), .B(n_1561), .Y(n_1560) );
AO22x1_ASAP7_75t_L g1708 ( .A1(n_184), .A2(n_364), .B1(n_1667), .B2(n_1709), .Y(n_1708) );
CKINVDCx16_ASAP7_75t_R g1779 ( .A(n_185), .Y(n_1779) );
INVx1_ASAP7_75t_L g647 ( .A(n_186), .Y(n_647) );
INVx1_ASAP7_75t_L g1954 ( .A(n_187), .Y(n_1954) );
AOI22xp33_ASAP7_75t_SL g1599 ( .A1(n_188), .A2(n_326), .B1(n_1357), .B2(n_1598), .Y(n_1599) );
XOR2x2_ASAP7_75t_L g709 ( .A(n_189), .B(n_710), .Y(n_709) );
INVxp67_ASAP7_75t_SL g1305 ( .A(n_190), .Y(n_1305) );
CKINVDCx5p33_ASAP7_75t_R g1102 ( .A(n_191), .Y(n_1102) );
INVx1_ASAP7_75t_L g760 ( .A(n_192), .Y(n_760) );
INVx1_ASAP7_75t_L g730 ( .A(n_193), .Y(n_730) );
INVx1_ASAP7_75t_L g1227 ( .A(n_194), .Y(n_1227) );
INVx1_ASAP7_75t_L g816 ( .A(n_195), .Y(n_816) );
INVx1_ASAP7_75t_L g1571 ( .A(n_196), .Y(n_1571) );
OAI22xp5_ASAP7_75t_L g1576 ( .A1(n_196), .A2(n_318), .B1(n_1577), .B2(n_1578), .Y(n_1576) );
INVx1_ASAP7_75t_L g1153 ( .A(n_197), .Y(n_1153) );
INVx1_ASAP7_75t_L g794 ( .A(n_198), .Y(n_794) );
INVx1_ASAP7_75t_L g1461 ( .A(n_200), .Y(n_1461) );
INVx1_ASAP7_75t_L g1337 ( .A(n_202), .Y(n_1337) );
INVx1_ASAP7_75t_L g1440 ( .A(n_203), .Y(n_1440) );
OAI211xp5_ASAP7_75t_L g1446 ( .A1(n_203), .A2(n_757), .B(n_1447), .C(n_1448), .Y(n_1446) );
INVx1_ASAP7_75t_L g1906 ( .A(n_205), .Y(n_1906) );
OAI211xp5_ASAP7_75t_L g1911 ( .A1(n_205), .A2(n_427), .B(n_518), .C(n_1912), .Y(n_1911) );
OAI22xp33_ASAP7_75t_L g625 ( .A1(n_206), .A2(n_360), .B1(n_512), .B2(n_626), .Y(n_625) );
OAI22xp33_ASAP7_75t_L g635 ( .A1(n_206), .A2(n_360), .B1(n_555), .B2(n_558), .Y(n_635) );
INVx1_ASAP7_75t_L g1948 ( .A(n_207), .Y(n_1948) );
INVx1_ASAP7_75t_L g966 ( .A(n_208), .Y(n_966) );
AOI221x1_ASAP7_75t_SL g997 ( .A1(n_208), .A2(n_285), .B1(n_436), .B2(n_998), .C(n_1000), .Y(n_997) );
INVx1_ASAP7_75t_L g1394 ( .A(n_209), .Y(n_1394) );
AOI221x1_ASAP7_75t_SL g1088 ( .A1(n_210), .A2(n_280), .B1(n_1089), .B2(n_1093), .C(n_1095), .Y(n_1088) );
AOI21xp33_ASAP7_75t_L g1155 ( .A1(n_210), .A2(n_600), .B(n_1156), .Y(n_1155) );
AOI21xp33_ASAP7_75t_L g979 ( .A1(n_211), .A2(n_980), .B(n_981), .Y(n_979) );
INVx1_ASAP7_75t_L g1009 ( .A(n_211), .Y(n_1009) );
INVx2_ASAP7_75t_L g1670 ( .A(n_213), .Y(n_1670) );
AND2x2_ASAP7_75t_L g1672 ( .A(n_213), .B(n_321), .Y(n_1672) );
AND2x2_ASAP7_75t_L g1678 ( .A(n_213), .B(n_1676), .Y(n_1678) );
INVx1_ASAP7_75t_L g822 ( .A(n_214), .Y(n_822) );
OAI22xp33_ASAP7_75t_L g762 ( .A1(n_216), .A2(n_279), .B1(n_763), .B2(n_764), .Y(n_762) );
OAI22xp33_ASAP7_75t_L g780 ( .A1(n_216), .A2(n_279), .B1(n_704), .B2(n_781), .Y(n_780) );
INVx1_ASAP7_75t_L g1618 ( .A(n_217), .Y(n_1618) );
INVx1_ASAP7_75t_L g826 ( .A(n_218), .Y(n_826) );
INVx1_ASAP7_75t_L g1343 ( .A(n_219), .Y(n_1343) );
INVx1_ASAP7_75t_L g1021 ( .A(n_220), .Y(n_1021) );
INVx1_ASAP7_75t_L g1932 ( .A(n_221), .Y(n_1932) );
INVx1_ASAP7_75t_L g883 ( .A(n_222), .Y(n_883) );
CKINVDCx5p33_ASAP7_75t_R g1098 ( .A(n_223), .Y(n_1098) );
INVx1_ASAP7_75t_L g833 ( .A(n_224), .Y(n_833) );
AOI22xp33_ASAP7_75t_L g1355 ( .A1(n_225), .A2(n_357), .B1(n_1356), .B2(n_1357), .Y(n_1355) );
AOI22xp33_ASAP7_75t_L g1377 ( .A1(n_225), .A2(n_229), .B1(n_1378), .B2(n_1379), .Y(n_1377) );
INVx1_ASAP7_75t_L g1881 ( .A(n_226), .Y(n_1881) );
OAI211xp5_ASAP7_75t_L g1019 ( .A1(n_227), .A2(n_568), .B(n_610), .C(n_1020), .Y(n_1019) );
INVx1_ASAP7_75t_L g1065 ( .A(n_227), .Y(n_1065) );
XOR2x2_ASAP7_75t_L g1473 ( .A(n_228), .B(n_1474), .Y(n_1473) );
AOI22xp33_ASAP7_75t_SL g1367 ( .A1(n_229), .A2(n_352), .B1(n_1356), .B2(n_1368), .Y(n_1367) );
AOI22xp33_ASAP7_75t_L g1284 ( .A1(n_230), .A2(n_330), .B1(n_436), .B2(n_1180), .Y(n_1284) );
XNOR2xp5_ASAP7_75t_L g786 ( .A(n_231), .B(n_787), .Y(n_786) );
INVx1_ASAP7_75t_L g722 ( .A(n_232), .Y(n_722) );
INVx1_ASAP7_75t_L g872 ( .A(n_233), .Y(n_872) );
INVx1_ASAP7_75t_L g1218 ( .A(n_234), .Y(n_1218) );
INVx1_ASAP7_75t_L g723 ( .A(n_235), .Y(n_723) );
INVx2_ASAP7_75t_L g415 ( .A(n_236), .Y(n_415) );
INVx1_ASAP7_75t_L g464 ( .A(n_236), .Y(n_464) );
NAND2xp5_ASAP7_75t_L g914 ( .A(n_236), .B(n_416), .Y(n_914) );
INVx1_ASAP7_75t_L g655 ( .A(n_237), .Y(n_655) );
INVx1_ASAP7_75t_L g1407 ( .A(n_238), .Y(n_1407) );
XNOR2xp5_ASAP7_75t_L g1601 ( .A(n_241), .B(n_1602), .Y(n_1601) );
INVx1_ASAP7_75t_L g1545 ( .A(n_242), .Y(n_1545) );
INVx1_ASAP7_75t_L g898 ( .A(n_243), .Y(n_898) );
INVx1_ASAP7_75t_L g834 ( .A(n_244), .Y(n_834) );
INVx1_ASAP7_75t_L g1399 ( .A(n_245), .Y(n_1399) );
INVx1_ASAP7_75t_L g1533 ( .A(n_246), .Y(n_1533) );
AOI22xp33_ASAP7_75t_SL g1583 ( .A1(n_247), .A2(n_326), .B1(n_1299), .B2(n_1584), .Y(n_1583) );
BUFx3_ASAP7_75t_L g423 ( .A(n_248), .Y(n_423) );
AOI22xp33_ASAP7_75t_L g1705 ( .A1(n_249), .A2(n_253), .B1(n_1674), .B2(n_1677), .Y(n_1705) );
AOI22xp33_ASAP7_75t_SL g1361 ( .A1(n_250), .A2(n_271), .B1(n_1362), .B2(n_1363), .Y(n_1361) );
INVx1_ASAP7_75t_L g732 ( .A(n_251), .Y(n_732) );
INVx1_ASAP7_75t_L g624 ( .A(n_252), .Y(n_624) );
OAI211xp5_ASAP7_75t_L g636 ( .A1(n_252), .A2(n_564), .B(n_568), .C(n_637), .Y(n_636) );
OAI22xp5_ASAP7_75t_SL g946 ( .A1(n_254), .A2(n_302), .B1(n_947), .B2(n_949), .Y(n_946) );
CKINVDCx5p33_ASAP7_75t_R g960 ( .A(n_254), .Y(n_960) );
INVx1_ASAP7_75t_L g1324 ( .A(n_255), .Y(n_1324) );
AOI22xp33_ASAP7_75t_L g1610 ( .A1(n_256), .A2(n_329), .B1(n_1299), .B2(n_1611), .Y(n_1610) );
AOI22xp33_ASAP7_75t_L g1654 ( .A1(n_256), .A2(n_275), .B1(n_954), .B2(n_1198), .Y(n_1654) );
INVx1_ASAP7_75t_L g1455 ( .A(n_257), .Y(n_1455) );
INVx1_ASAP7_75t_L g1947 ( .A(n_258), .Y(n_1947) );
AOI21xp33_ASAP7_75t_L g1237 ( .A1(n_259), .A2(n_980), .B(n_981), .Y(n_1237) );
INVx1_ASAP7_75t_L g858 ( .A(n_260), .Y(n_858) );
INVx1_ASAP7_75t_L g1035 ( .A(n_261), .Y(n_1035) );
INVx1_ASAP7_75t_L g1498 ( .A(n_262), .Y(n_1498) );
INVx1_ASAP7_75t_L g1950 ( .A(n_264), .Y(n_1950) );
INVx1_ASAP7_75t_L g1531 ( .A(n_265), .Y(n_1531) );
INVx1_ASAP7_75t_L g1129 ( .A(n_266), .Y(n_1129) );
INVx1_ASAP7_75t_L g456 ( .A(n_267), .Y(n_456) );
INVx1_ASAP7_75t_L g1277 ( .A(n_268), .Y(n_1277) );
INVx1_ASAP7_75t_L g814 ( .A(n_269), .Y(n_814) );
BUFx3_ASAP7_75t_L g399 ( .A(n_272), .Y(n_399) );
INVx1_ASAP7_75t_L g551 ( .A(n_272), .Y(n_551) );
CKINVDCx20_ASAP7_75t_R g1781 ( .A(n_273), .Y(n_1781) );
AOI22xp5_ASAP7_75t_L g1681 ( .A1(n_274), .A2(n_294), .B1(n_1674), .B2(n_1677), .Y(n_1681) );
INVx1_ASAP7_75t_L g1152 ( .A(n_280), .Y(n_1152) );
INVx1_ASAP7_75t_L g1524 ( .A(n_281), .Y(n_1524) );
INVx1_ASAP7_75t_L g1075 ( .A(n_284), .Y(n_1075) );
AOI22xp33_ASAP7_75t_L g982 ( .A1(n_285), .A2(n_292), .B1(n_972), .B2(n_974), .Y(n_982) );
INVx1_ASAP7_75t_L g1525 ( .A(n_286), .Y(n_1525) );
INVx1_ASAP7_75t_L g1504 ( .A(n_287), .Y(n_1504) );
INVx1_ASAP7_75t_L g1022 ( .A(n_288), .Y(n_1022) );
OAI211xp5_ASAP7_75t_L g1063 ( .A1(n_288), .A2(n_518), .B(n_604), .C(n_1064), .Y(n_1063) );
INVx1_ASAP7_75t_L g855 ( .A(n_289), .Y(n_855) );
INVx1_ASAP7_75t_L g1893 ( .A(n_291), .Y(n_1893) );
INVx1_ASAP7_75t_L g1458 ( .A(n_293), .Y(n_1458) );
OAI22xp5_ASAP7_75t_L g1346 ( .A1(n_295), .A2(n_375), .B1(n_753), .B2(n_764), .Y(n_1346) );
INVx1_ASAP7_75t_L g1040 ( .A(n_296), .Y(n_1040) );
INVx1_ASAP7_75t_L g1503 ( .A(n_297), .Y(n_1503) );
CKINVDCx5p33_ASAP7_75t_R g1193 ( .A(n_299), .Y(n_1193) );
AOI22xp5_ASAP7_75t_L g1691 ( .A1(n_300), .A2(n_369), .B1(n_1674), .B2(n_1677), .Y(n_1691) );
AO22x1_ASAP7_75t_L g1666 ( .A1(n_301), .A2(n_307), .B1(n_1667), .B2(n_1671), .Y(n_1666) );
INVx1_ASAP7_75t_L g953 ( .A(n_302), .Y(n_953) );
INVx1_ASAP7_75t_L g1500 ( .A(n_303), .Y(n_1500) );
INVx1_ASAP7_75t_L g425 ( .A(n_304), .Y(n_425) );
INVx1_ASAP7_75t_L g431 ( .A(n_304), .Y(n_431) );
INVx1_ASAP7_75t_L g690 ( .A(n_306), .Y(n_690) );
OAI211xp5_ASAP7_75t_L g696 ( .A1(n_306), .A2(n_564), .B(n_697), .C(n_698), .Y(n_696) );
INVx1_ASAP7_75t_L g1887 ( .A(n_308), .Y(n_1887) );
INVx1_ASAP7_75t_L g598 ( .A(n_309), .Y(n_598) );
INVx1_ASAP7_75t_L g1507 ( .A(n_310), .Y(n_1507) );
INVx1_ASAP7_75t_L g857 ( .A(n_311), .Y(n_857) );
INVx1_ASAP7_75t_L g977 ( .A(n_313), .Y(n_977) );
INVx1_ASAP7_75t_L g528 ( .A(n_314), .Y(n_528) );
INVx1_ASAP7_75t_L g727 ( .A(n_316), .Y(n_727) );
AOI22xp5_ASAP7_75t_L g1015 ( .A1(n_317), .A2(n_1016), .B1(n_1017), .B2(n_1068), .Y(n_1015) );
INVxp67_ASAP7_75t_SL g1068 ( .A(n_317), .Y(n_1068) );
INVx1_ASAP7_75t_L g1572 ( .A(n_318), .Y(n_1572) );
CKINVDCx5p33_ASAP7_75t_R g1186 ( .A(n_319), .Y(n_1186) );
INVxp67_ASAP7_75t_SL g1650 ( .A(n_320), .Y(n_1650) );
AND2x2_ASAP7_75t_L g1669 ( .A(n_321), .B(n_1670), .Y(n_1669) );
INVx1_ASAP7_75t_L g1676 ( .A(n_321), .Y(n_1676) );
OAI211xp5_ASAP7_75t_SL g514 ( .A1(n_322), .A2(n_515), .B(n_518), .C(n_522), .Y(n_514) );
INVx1_ASAP7_75t_L g582 ( .A(n_322), .Y(n_582) );
INVx1_ASAP7_75t_L g1573 ( .A(n_323), .Y(n_1573) );
INVx1_ASAP7_75t_L g1170 ( .A(n_324), .Y(n_1170) );
OAI211xp5_ASAP7_75t_L g754 ( .A1(n_325), .A2(n_755), .B(n_757), .C(n_758), .Y(n_754) );
INVx1_ASAP7_75t_L g779 ( .A(n_325), .Y(n_779) );
INVx1_ASAP7_75t_L g1635 ( .A(n_327), .Y(n_1635) );
INVx1_ASAP7_75t_L g1454 ( .A(n_328), .Y(n_1454) );
INVx1_ASAP7_75t_L g1312 ( .A(n_330), .Y(n_1312) );
INVx1_ASAP7_75t_L g828 ( .A(n_331), .Y(n_828) );
INVx1_ASAP7_75t_L g795 ( .A(n_332), .Y(n_795) );
OAI211xp5_ASAP7_75t_L g804 ( .A1(n_332), .A2(n_757), .B(n_805), .C(n_806), .Y(n_804) );
INVx1_ASAP7_75t_L g1247 ( .A(n_333), .Y(n_1247) );
INVx1_ASAP7_75t_L g665 ( .A(n_334), .Y(n_665) );
INVx1_ASAP7_75t_L g1885 ( .A(n_335), .Y(n_1885) );
INVx1_ASAP7_75t_L g1506 ( .A(n_336), .Y(n_1506) );
INVx1_ASAP7_75t_L g1528 ( .A(n_337), .Y(n_1528) );
OAI22xp5_ASAP7_75t_L g1329 ( .A1(n_338), .A2(n_1330), .B1(n_1381), .B2(n_1382), .Y(n_1329) );
INVxp67_ASAP7_75t_SL g1382 ( .A(n_338), .Y(n_1382) );
AOI211xp5_ASAP7_75t_SL g1213 ( .A1(n_339), .A2(n_1214), .B(n_1215), .C(n_1217), .Y(n_1213) );
INVx1_ASAP7_75t_L g1404 ( .A(n_340), .Y(n_1404) );
AOI21xp5_ASAP7_75t_SL g1242 ( .A1(n_341), .A2(n_980), .B(n_1243), .Y(n_1242) );
INVx1_ASAP7_75t_L g1257 ( .A(n_341), .Y(n_1257) );
OAI22xp5_ASAP7_75t_L g808 ( .A1(n_342), .A2(n_373), .B1(n_512), .B2(n_809), .Y(n_808) );
INVx1_ASAP7_75t_L g1311 ( .A(n_344), .Y(n_1311) );
XNOR2xp5_ASAP7_75t_L g587 ( .A(n_345), .B(n_588), .Y(n_587) );
INVx1_ASAP7_75t_L g603 ( .A(n_346), .Y(n_603) );
INVxp67_ASAP7_75t_L g1263 ( .A(n_348), .Y(n_1263) );
OAI211xp5_ASAP7_75t_L g1929 ( .A1(n_349), .A2(n_757), .B(n_1930), .C(n_1931), .Y(n_1929) );
INVx1_ASAP7_75t_L g1940 ( .A(n_349), .Y(n_1940) );
INVxp67_ASAP7_75t_SL g1276 ( .A(n_350), .Y(n_1276) );
BUFx6f_ASAP7_75t_L g395 ( .A(n_351), .Y(n_395) );
AOI22xp33_ASAP7_75t_SL g1374 ( .A1(n_352), .A2(n_357), .B1(n_1296), .B2(n_1375), .Y(n_1374) );
INVx1_ASAP7_75t_L g1033 ( .A(n_353), .Y(n_1033) );
INVx1_ASAP7_75t_L g1046 ( .A(n_354), .Y(n_1046) );
CKINVDCx5p33_ASAP7_75t_R g1120 ( .A(n_356), .Y(n_1120) );
INVx1_ASAP7_75t_L g1565 ( .A(n_361), .Y(n_1565) );
INVx1_ASAP7_75t_L g1464 ( .A(n_362), .Y(n_1464) );
INVx1_ASAP7_75t_L g1501 ( .A(n_365), .Y(n_1501) );
INVx1_ASAP7_75t_L g884 ( .A(n_366), .Y(n_884) );
OAI211xp5_ASAP7_75t_L g889 ( .A1(n_366), .A2(n_568), .B(n_890), .C(n_892), .Y(n_889) );
INVx1_ASAP7_75t_L g413 ( .A(n_368), .Y(n_413) );
INVx1_ASAP7_75t_L g463 ( .A(n_368), .Y(n_463) );
INVx2_ASAP7_75t_L g469 ( .A(n_368), .Y(n_469) );
XOR2x2_ASAP7_75t_L g1875 ( .A(n_369), .B(n_1876), .Y(n_1875) );
AOI22xp33_ASAP7_75t_L g1919 ( .A1(n_369), .A2(n_1920), .B1(n_1923), .B2(n_1964), .Y(n_1919) );
CKINVDCx5p33_ASAP7_75t_R g1121 ( .A(n_370), .Y(n_1121) );
INVx1_ASAP7_75t_L g945 ( .A(n_371), .Y(n_945) );
INVx1_ASAP7_75t_L g1894 ( .A(n_372), .Y(n_1894) );
CKINVDCx5p33_ASAP7_75t_R g1172 ( .A(n_374), .Y(n_1172) );
INVx1_ASAP7_75t_L g1335 ( .A(n_375), .Y(n_1335) );
AOI21xp5_ASAP7_75t_L g376 ( .A1(n_377), .A2(n_400), .B(n_1658), .Y(n_376) );
INVx2_ASAP7_75t_L g377 ( .A(n_378), .Y(n_377) );
OR2x2_ASAP7_75t_L g378 ( .A(n_379), .B(n_385), .Y(n_378) );
NOR2xp33_ASAP7_75t_L g1918 ( .A(n_379), .B(n_388), .Y(n_1918) );
INVx1_ASAP7_75t_L g379 ( .A(n_380), .Y(n_379) );
NOR2xp33_ASAP7_75t_L g380 ( .A(n_381), .B(n_383), .Y(n_380) );
NOR2xp33_ASAP7_75t_L g1922 ( .A(n_381), .B(n_384), .Y(n_1922) );
INVx1_ASAP7_75t_L g1967 ( .A(n_381), .Y(n_1967) );
HB1xp67_ASAP7_75t_L g381 ( .A(n_382), .Y(n_381) );
INVx1_ASAP7_75t_L g383 ( .A(n_384), .Y(n_383) );
NOR2xp33_ASAP7_75t_L g1969 ( .A(n_384), .B(n_1967), .Y(n_1969) );
INVx1_ASAP7_75t_L g385 ( .A(n_386), .Y(n_385) );
NAND2xp5_ASAP7_75t_L g386 ( .A(n_387), .B(n_390), .Y(n_386) );
INVx1_ASAP7_75t_L g387 ( .A(n_388), .Y(n_387) );
AND2x4_ASAP7_75t_L g584 ( .A(n_388), .B(n_585), .Y(n_584) );
INVx1_ASAP7_75t_L g388 ( .A(n_389), .Y(n_388) );
AND2x4_ASAP7_75t_L g497 ( .A(n_389), .B(n_399), .Y(n_497) );
AND2x4_ASAP7_75t_L g970 ( .A(n_389), .B(n_398), .Y(n_970) );
INVxp67_ASAP7_75t_SL g547 ( .A(n_390), .Y(n_547) );
INVx1_ASAP7_75t_L g1024 ( .A(n_390), .Y(n_1024) );
AOI22xp33_ASAP7_75t_L g1567 ( .A1(n_390), .A2(n_549), .B1(n_1568), .B2(n_1569), .Y(n_1567) );
AND2x4_ASAP7_75t_SL g1917 ( .A(n_390), .B(n_1918), .Y(n_1917) );
INVx3_ASAP7_75t_L g390 ( .A(n_391), .Y(n_390) );
OR2x6_ASAP7_75t_L g391 ( .A(n_392), .B(n_397), .Y(n_391) );
INVx1_ASAP7_75t_L g504 ( .A(n_392), .Y(n_504) );
OR2x6_ASAP7_75t_L g557 ( .A(n_392), .B(n_550), .Y(n_557) );
BUFx4f_ASAP7_75t_L g669 ( .A(n_392), .Y(n_669) );
INVx2_ASAP7_75t_L g392 ( .A(n_393), .Y(n_392) );
BUFx4f_ASAP7_75t_L g474 ( .A(n_393), .Y(n_474) );
INVx3_ASAP7_75t_L g679 ( .A(n_393), .Y(n_679) );
INVx3_ASAP7_75t_L g393 ( .A(n_394), .Y(n_393) );
OR2x2_ASAP7_75t_L g394 ( .A(n_395), .B(n_396), .Y(n_394) );
INVx2_ASAP7_75t_L g480 ( .A(n_395), .Y(n_480) );
INVx2_ASAP7_75t_L g487 ( .A(n_395), .Y(n_487) );
NAND2x1_ASAP7_75t_L g491 ( .A(n_395), .B(n_396), .Y(n_491) );
AND2x2_ASAP7_75t_L g552 ( .A(n_395), .B(n_553), .Y(n_552) );
AND2x2_ASAP7_75t_L g572 ( .A(n_395), .B(n_396), .Y(n_572) );
INVx1_ASAP7_75t_L g581 ( .A(n_395), .Y(n_581) );
NAND2xp5_ASAP7_75t_L g479 ( .A(n_396), .B(n_480), .Y(n_479) );
OR2x2_ASAP7_75t_L g486 ( .A(n_396), .B(n_487), .Y(n_486) );
INVx2_ASAP7_75t_L g553 ( .A(n_396), .Y(n_553) );
BUFx2_ASAP7_75t_L g576 ( .A(n_396), .Y(n_576) );
INVx1_ASAP7_75t_L g909 ( .A(n_396), .Y(n_909) );
AND2x2_ASAP7_75t_L g975 ( .A(n_396), .B(n_480), .Y(n_975) );
OR2x6_ASAP7_75t_L g771 ( .A(n_397), .B(n_679), .Y(n_771) );
INVxp67_ASAP7_75t_L g397 ( .A(n_398), .Y(n_397) );
INVx1_ASAP7_75t_L g570 ( .A(n_398), .Y(n_570) );
INVx2_ASAP7_75t_L g398 ( .A(n_399), .Y(n_398) );
BUFx2_ASAP7_75t_L g562 ( .A(n_399), .Y(n_562) );
AND2x4_ASAP7_75t_L g579 ( .A(n_399), .B(n_580), .Y(n_579) );
XNOR2xp5_ASAP7_75t_L g400 ( .A(n_401), .B(n_844), .Y(n_400) );
XNOR2xp5_ASAP7_75t_L g401 ( .A(n_402), .B(n_784), .Y(n_401) );
HB1xp67_ASAP7_75t_L g402 ( .A(n_403), .Y(n_402) );
XNOR2xp5_ASAP7_75t_L g403 ( .A(n_404), .B(n_639), .Y(n_403) );
XOR2xp5_ASAP7_75t_L g404 ( .A(n_405), .B(n_587), .Y(n_404) );
AND3x1_ASAP7_75t_L g406 ( .A(n_407), .B(n_507), .C(n_545), .Y(n_406) );
NOR2xp33_ASAP7_75t_L g407 ( .A(n_408), .B(n_465), .Y(n_407) );
OAI33xp33_ASAP7_75t_L g408 ( .A1(n_409), .A2(n_417), .A3(n_433), .B1(n_446), .B2(n_455), .B3(n_458), .Y(n_408) );
OAI33xp33_ASAP7_75t_L g590 ( .A1(n_409), .A2(n_458), .A3(n_591), .B1(n_594), .B2(n_597), .B3(n_602), .Y(n_590) );
OAI33xp33_ASAP7_75t_L g835 ( .A1(n_409), .A2(n_458), .A3(n_836), .B1(n_838), .B2(n_839), .B3(n_841), .Y(n_835) );
OAI33xp33_ASAP7_75t_L g1508 ( .A1(n_409), .A2(n_458), .A3(n_1509), .B1(n_1512), .B2(n_1513), .B3(n_1516), .Y(n_1508) );
OAI33xp33_ASAP7_75t_L g1535 ( .A1(n_409), .A2(n_1266), .A3(n_1536), .B1(n_1537), .B2(n_1539), .B3(n_1540), .Y(n_1535) );
BUFx4f_ASAP7_75t_L g409 ( .A(n_410), .Y(n_409) );
BUFx4f_ASAP7_75t_L g657 ( .A(n_410), .Y(n_657) );
BUFx8_ASAP7_75t_L g735 ( .A(n_410), .Y(n_735) );
BUFx2_ASAP7_75t_L g1392 ( .A(n_410), .Y(n_1392) );
OR2x2_ASAP7_75t_L g410 ( .A(n_411), .B(n_414), .Y(n_410) );
INVx1_ASAP7_75t_L g499 ( .A(n_411), .Y(n_499) );
HB1xp67_ASAP7_75t_L g544 ( .A(n_411), .Y(n_544) );
OR2x2_ASAP7_75t_L g913 ( .A(n_411), .B(n_914), .Y(n_913) );
AND2x2_ASAP7_75t_SL g1417 ( .A(n_411), .B(n_497), .Y(n_1417) );
INVx2_ASAP7_75t_L g411 ( .A(n_412), .Y(n_411) );
BUFx2_ASAP7_75t_L g586 ( .A(n_412), .Y(n_586) );
INVx1_ASAP7_75t_L g412 ( .A(n_413), .Y(n_412) );
BUFx2_ASAP7_75t_L g1156 ( .A(n_414), .Y(n_1156) );
NAND2xp33_ASAP7_75t_SL g414 ( .A(n_415), .B(n_416), .Y(n_414) );
HB1xp67_ASAP7_75t_L g542 ( .A(n_415), .Y(n_542) );
INVx1_ASAP7_75t_L g929 ( .A(n_415), .Y(n_929) );
AND3x4_ASAP7_75t_L g1011 ( .A(n_415), .B(n_526), .C(n_995), .Y(n_1011) );
INVx3_ASAP7_75t_L g461 ( .A(n_416), .Y(n_461) );
BUFx3_ASAP7_75t_L g526 ( .A(n_416), .Y(n_526) );
OAI22xp33_ASAP7_75t_L g417 ( .A1(n_418), .A2(n_419), .B1(n_426), .B2(n_427), .Y(n_417) );
OAI22xp33_ASAP7_75t_L g471 ( .A1(n_418), .A2(n_456), .B1(n_472), .B2(n_475), .Y(n_471) );
OAI22xp33_ASAP7_75t_L g455 ( .A1(n_419), .A2(n_427), .B1(n_456), .B2(n_457), .Y(n_455) );
OAI22xp33_ASAP7_75t_L g591 ( .A1(n_419), .A2(n_427), .B1(n_592), .B2(n_593), .Y(n_591) );
OAI22xp33_ASAP7_75t_L g602 ( .A1(n_419), .A2(n_603), .B1(n_604), .B2(n_606), .Y(n_602) );
OAI22xp33_ASAP7_75t_L g1959 ( .A1(n_419), .A2(n_1947), .B1(n_1953), .B2(n_1960), .Y(n_1959) );
OAI22xp33_ASAP7_75t_L g1963 ( .A1(n_419), .A2(n_1003), .B1(n_1948), .B2(n_1954), .Y(n_1963) );
INVx2_ASAP7_75t_L g419 ( .A(n_420), .Y(n_419) );
INVx1_ASAP7_75t_L g420 ( .A(n_421), .Y(n_420) );
BUFx3_ASAP7_75t_L g421 ( .A(n_422), .Y(n_421) );
OR2x4_ASAP7_75t_L g510 ( .A(n_422), .B(n_511), .Y(n_510) );
OR2x4_ASAP7_75t_L g536 ( .A(n_422), .B(n_461), .Y(n_536) );
INVx2_ASAP7_75t_L g654 ( .A(n_422), .Y(n_654) );
BUFx3_ASAP7_75t_L g660 ( .A(n_422), .Y(n_660) );
BUFx4f_ASAP7_75t_L g843 ( .A(n_422), .Y(n_843) );
OR2x2_ASAP7_75t_L g422 ( .A(n_423), .B(n_424), .Y(n_422) );
BUFx6f_ASAP7_75t_L g432 ( .A(n_423), .Y(n_432) );
INVx2_ASAP7_75t_L g441 ( .A(n_423), .Y(n_441) );
NAND2xp5_ASAP7_75t_L g445 ( .A(n_423), .B(n_431), .Y(n_445) );
AND2x4_ASAP7_75t_L g520 ( .A(n_423), .B(n_521), .Y(n_520) );
INVx1_ASAP7_75t_L g927 ( .A(n_424), .Y(n_927) );
INVx1_ASAP7_75t_L g424 ( .A(n_425), .Y(n_424) );
INVxp67_ASAP7_75t_L g440 ( .A(n_425), .Y(n_440) );
OAI22xp33_ASAP7_75t_L g492 ( .A1(n_426), .A2(n_457), .B1(n_488), .B2(n_493), .Y(n_492) );
OAI22xp33_ASAP7_75t_L g841 ( .A1(n_427), .A2(n_816), .B1(n_828), .B2(n_842), .Y(n_841) );
OAI22xp33_ASAP7_75t_L g853 ( .A1(n_427), .A2(n_842), .B1(n_854), .B2(n_855), .Y(n_853) );
OAI22xp33_ASAP7_75t_L g1516 ( .A1(n_427), .A2(n_1498), .B1(n_1504), .B2(n_1517), .Y(n_1516) );
OAI22xp33_ASAP7_75t_L g1536 ( .A1(n_427), .A2(n_837), .B1(n_1524), .B2(n_1530), .Y(n_1536) );
OAI22xp33_ASAP7_75t_L g1892 ( .A1(n_427), .A2(n_1510), .B1(n_1893), .B2(n_1894), .Y(n_1892) );
BUFx6f_ASAP7_75t_L g427 ( .A(n_428), .Y(n_427) );
INVx2_ASAP7_75t_L g605 ( .A(n_428), .Y(n_605) );
OAI22xp33_ASAP7_75t_L g1470 ( .A1(n_428), .A2(n_653), .B1(n_1455), .B2(n_1462), .Y(n_1470) );
BUFx3_ASAP7_75t_L g428 ( .A(n_429), .Y(n_428) );
BUFx2_ASAP7_75t_L g517 ( .A(n_429), .Y(n_517) );
BUFx6f_ASAP7_75t_L g739 ( .A(n_429), .Y(n_739) );
NAND2x1p5_ASAP7_75t_L g429 ( .A(n_430), .B(n_432), .Y(n_429) );
BUFx2_ASAP7_75t_L g531 ( .A(n_430), .Y(n_531) );
INVx1_ASAP7_75t_L g430 ( .A(n_431), .Y(n_430) );
INVx2_ASAP7_75t_L g521 ( .A(n_431), .Y(n_521) );
BUFx2_ASAP7_75t_L g527 ( .A(n_432), .Y(n_527) );
INVx2_ASAP7_75t_L g936 ( .A(n_432), .Y(n_936) );
AND2x4_ASAP7_75t_L g999 ( .A(n_432), .B(n_944), .Y(n_999) );
OAI22xp5_ASAP7_75t_L g433 ( .A1(n_434), .A2(n_435), .B1(n_442), .B2(n_443), .Y(n_433) );
OAI22xp5_ASAP7_75t_L g481 ( .A1(n_434), .A2(n_447), .B1(n_482), .B2(n_488), .Y(n_481) );
OAI22xp5_ASAP7_75t_L g594 ( .A1(n_435), .A2(n_443), .B1(n_595), .B2(n_596), .Y(n_594) );
OAI22xp5_ASAP7_75t_L g1034 ( .A1(n_435), .A2(n_1035), .B1(n_1036), .B2(n_1037), .Y(n_1034) );
OAI22xp5_ASAP7_75t_L g1539 ( .A1(n_435), .A2(n_859), .B1(n_1528), .B2(n_1534), .Y(n_1539) );
INVx2_ASAP7_75t_L g435 ( .A(n_436), .Y(n_435) );
INVx1_ASAP7_75t_L g646 ( .A(n_436), .Y(n_646) );
INVx8_ASAP7_75t_L g436 ( .A(n_437), .Y(n_436) );
BUFx3_ASAP7_75t_L g664 ( .A(n_437), .Y(n_664) );
OAI22xp5_ASAP7_75t_L g1962 ( .A1(n_437), .A2(n_648), .B1(n_1951), .B2(n_1957), .Y(n_1962) );
INVx5_ASAP7_75t_L g437 ( .A(n_438), .Y(n_437) );
INVx3_ASAP7_75t_L g450 ( .A(n_438), .Y(n_450) );
INVx2_ASAP7_75t_SL g1179 ( .A(n_438), .Y(n_1179) );
AOI22xp33_ASAP7_75t_L g1272 ( .A1(n_438), .A2(n_1175), .B1(n_1273), .B2(n_1274), .Y(n_1272) );
HB1xp67_ASAP7_75t_L g1515 ( .A(n_438), .Y(n_1515) );
INVx2_ASAP7_75t_SL g1538 ( .A(n_438), .Y(n_1538) );
BUFx6f_ASAP7_75t_L g438 ( .A(n_439), .Y(n_438) );
BUFx6f_ASAP7_75t_L g539 ( .A(n_439), .Y(n_539) );
BUFx8_ASAP7_75t_L g600 ( .A(n_439), .Y(n_600) );
INVx2_ASAP7_75t_L g863 ( .A(n_439), .Y(n_863) );
AND2x4_ASAP7_75t_L g439 ( .A(n_440), .B(n_441), .Y(n_439) );
AND2x4_ASAP7_75t_L g926 ( .A(n_441), .B(n_927), .Y(n_926) );
OAI22xp5_ASAP7_75t_L g500 ( .A1(n_442), .A2(n_451), .B1(n_501), .B2(n_505), .Y(n_500) );
OAI22xp5_ASAP7_75t_L g663 ( .A1(n_443), .A2(n_664), .B1(n_665), .B2(n_666), .Y(n_663) );
OAI22xp5_ASAP7_75t_L g838 ( .A1(n_443), .A2(n_599), .B1(n_821), .B2(n_833), .Y(n_838) );
OAI22xp5_ASAP7_75t_L g1537 ( .A1(n_443), .A2(n_1527), .B1(n_1533), .B2(n_1538), .Y(n_1537) );
BUFx3_ASAP7_75t_L g443 ( .A(n_444), .Y(n_443) );
OR2x6_ASAP7_75t_L g513 ( .A(n_444), .B(n_461), .Y(n_513) );
INVx1_ASAP7_75t_L g650 ( .A(n_444), .Y(n_650) );
BUFx2_ASAP7_75t_L g444 ( .A(n_445), .Y(n_444) );
INVx1_ASAP7_75t_L g454 ( .A(n_445), .Y(n_454) );
OAI22xp5_ASAP7_75t_L g446 ( .A1(n_447), .A2(n_448), .B1(n_451), .B2(n_452), .Y(n_446) );
OAI22xp33_ASAP7_75t_SL g856 ( .A1(n_448), .A2(n_857), .B1(n_858), .B2(n_859), .Y(n_856) );
INVx2_ASAP7_75t_L g448 ( .A(n_449), .Y(n_448) );
AOI22xp33_ASAP7_75t_L g1136 ( .A1(n_449), .A2(n_1120), .B1(n_1121), .B2(n_1137), .Y(n_1136) );
INVx2_ASAP7_75t_L g449 ( .A(n_450), .Y(n_449) );
OAI22xp5_ASAP7_75t_L g597 ( .A1(n_452), .A2(n_598), .B1(n_599), .B2(n_601), .Y(n_597) );
OAI22xp5_ASAP7_75t_L g869 ( .A1(n_452), .A2(n_870), .B1(n_871), .B2(n_872), .Y(n_869) );
INVx3_ASAP7_75t_L g452 ( .A(n_453), .Y(n_452) );
INVx3_ASAP7_75t_L g743 ( .A(n_453), .Y(n_743) );
CKINVDCx8_ASAP7_75t_R g750 ( .A(n_453), .Y(n_750) );
INVx3_ASAP7_75t_L g1037 ( .A(n_453), .Y(n_1037) );
INVx1_ASAP7_75t_L g1400 ( .A(n_453), .Y(n_1400) );
BUFx6f_ASAP7_75t_L g453 ( .A(n_454), .Y(n_453) );
INVx1_ASAP7_75t_L g948 ( .A(n_454), .Y(n_948) );
OAI33xp33_ASAP7_75t_L g852 ( .A1(n_458), .A2(n_656), .A3(n_853), .B1(n_856), .B2(n_860), .B3(n_869), .Y(n_852) );
INVx2_ASAP7_75t_L g458 ( .A(n_459), .Y(n_458) );
CKINVDCx5p33_ASAP7_75t_R g662 ( .A(n_459), .Y(n_662) );
AOI221xp5_ASAP7_75t_L g996 ( .A1(n_459), .A2(n_997), .B1(n_1004), .B2(n_1010), .C(n_1012), .Y(n_996) );
INVx2_ASAP7_75t_L g1266 ( .A(n_459), .Y(n_1266) );
NAND3xp33_ASAP7_75t_L g1376 ( .A(n_459), .B(n_1377), .C(n_1380), .Y(n_1376) );
INVx3_ASAP7_75t_L g459 ( .A(n_460), .Y(n_459) );
INVx3_ASAP7_75t_L g1043 ( .A(n_460), .Y(n_1043) );
NAND3x1_ASAP7_75t_L g460 ( .A(n_461), .B(n_462), .C(n_464), .Y(n_460) );
INVx1_ASAP7_75t_L g511 ( .A(n_461), .Y(n_511) );
AND2x4_ASAP7_75t_L g519 ( .A(n_461), .B(n_520), .Y(n_519) );
NAND2x1p5_ASAP7_75t_L g747 ( .A(n_461), .B(n_464), .Y(n_747) );
AND2x4_ASAP7_75t_L g928 ( .A(n_461), .B(n_929), .Y(n_928) );
INVx1_ASAP7_75t_L g462 ( .A(n_463), .Y(n_462) );
INVx1_ASAP7_75t_L g938 ( .A(n_463), .Y(n_938) );
NAND2xp5_ASAP7_75t_L g1085 ( .A(n_463), .B(n_907), .Y(n_1085) );
OAI33xp33_ASAP7_75t_L g465 ( .A1(n_466), .A2(n_471), .A3(n_481), .B1(n_492), .B2(n_495), .B3(n_500), .Y(n_465) );
OAI33xp33_ASAP7_75t_L g607 ( .A1(n_466), .A2(n_495), .A3(n_608), .B1(n_609), .B2(n_611), .B3(n_615), .Y(n_607) );
INVx1_ASAP7_75t_L g466 ( .A(n_467), .Y(n_466) );
INVx1_ASAP7_75t_L g671 ( .A(n_467), .Y(n_671) );
INVx4_ASAP7_75t_L g715 ( .A(n_467), .Y(n_715) );
INVx2_ASAP7_75t_L g874 ( .A(n_467), .Y(n_874) );
INVx2_ASAP7_75t_L g1456 ( .A(n_467), .Y(n_1456) );
INVx2_ASAP7_75t_L g1593 ( .A(n_467), .Y(n_1593) );
AND2x4_ASAP7_75t_L g467 ( .A(n_468), .B(n_470), .Y(n_467) );
OR2x6_ASAP7_75t_L g746 ( .A(n_468), .B(n_747), .Y(n_746) );
INVx1_ASAP7_75t_L g1160 ( .A(n_468), .Y(n_1160) );
BUFx2_ASAP7_75t_L g468 ( .A(n_469), .Y(n_468) );
INVx2_ASAP7_75t_L g995 ( .A(n_469), .Y(n_995) );
NAND2xp5_ASAP7_75t_L g1112 ( .A(n_469), .B(n_964), .Y(n_1112) );
OAI22xp33_ASAP7_75t_L g608 ( .A1(n_472), .A2(n_475), .B1(n_592), .B2(n_603), .Y(n_608) );
INVx2_ASAP7_75t_L g472 ( .A(n_473), .Y(n_472) );
INVx3_ASAP7_75t_L g731 ( .A(n_473), .Y(n_731) );
INVx2_ASAP7_75t_SL g815 ( .A(n_473), .Y(n_815) );
BUFx6f_ASAP7_75t_L g473 ( .A(n_474), .Y(n_473) );
INVx3_ASAP7_75t_L g1051 ( .A(n_474), .Y(n_1051) );
INVx4_ASAP7_75t_L g1219 ( .A(n_474), .Y(n_1219) );
OAI22xp5_ASAP7_75t_L g677 ( .A1(n_475), .A2(n_647), .B1(n_666), .B2(n_678), .Y(n_677) );
INVx6_ASAP7_75t_L g475 ( .A(n_476), .Y(n_475) );
INVx5_ASAP7_75t_L g616 ( .A(n_476), .Y(n_616) );
BUFx6f_ASAP7_75t_L g476 ( .A(n_477), .Y(n_476) );
INVx1_ASAP7_75t_L g506 ( .A(n_477), .Y(n_506) );
INVx1_ASAP7_75t_L g670 ( .A(n_477), .Y(n_670) );
INVx2_ASAP7_75t_L g720 ( .A(n_477), .Y(n_720) );
INVx2_ASAP7_75t_L g733 ( .A(n_477), .Y(n_733) );
INVx2_ASAP7_75t_SL g819 ( .A(n_477), .Y(n_819) );
INVx4_ASAP7_75t_L g1054 ( .A(n_477), .Y(n_1054) );
INVx2_ASAP7_75t_L g1316 ( .A(n_477), .Y(n_1316) );
INVx8_ASAP7_75t_L g477 ( .A(n_478), .Y(n_477) );
OR2x2_ASAP7_75t_L g561 ( .A(n_478), .B(n_562), .Y(n_561) );
BUFx2_ASAP7_75t_L g1415 ( .A(n_478), .Y(n_1415) );
BUFx6f_ASAP7_75t_L g478 ( .A(n_479), .Y(n_478) );
INVx1_ASAP7_75t_L g482 ( .A(n_483), .Y(n_482) );
INVx1_ASAP7_75t_L g483 ( .A(n_484), .Y(n_483) );
OAI22xp5_ASAP7_75t_L g1055 ( .A1(n_484), .A2(n_773), .B1(n_1035), .B2(n_1039), .Y(n_1055) );
OAI22xp5_ASAP7_75t_L g1056 ( .A1(n_484), .A2(n_773), .B1(n_1033), .B2(n_1046), .Y(n_1056) );
OAI221xp5_ASAP7_75t_L g1310 ( .A1(n_484), .A2(n_970), .B1(n_978), .B2(n_1311), .C(n_1312), .Y(n_1310) );
OAI22xp5_ASAP7_75t_L g1499 ( .A1(n_484), .A2(n_773), .B1(n_1500), .B2(n_1501), .Y(n_1499) );
OAI22xp5_ASAP7_75t_L g1502 ( .A1(n_484), .A2(n_488), .B1(n_1503), .B2(n_1504), .Y(n_1502) );
OAI22xp5_ASAP7_75t_L g1898 ( .A1(n_484), .A2(n_1883), .B1(n_1887), .B2(n_1899), .Y(n_1898) );
INVx2_ASAP7_75t_L g484 ( .A(n_485), .Y(n_484) );
INVx2_ASAP7_75t_L g1202 ( .A(n_485), .Y(n_1202) );
INVx2_ASAP7_75t_L g485 ( .A(n_486), .Y(n_485) );
BUFx3_ASAP7_75t_L g494 ( .A(n_486), .Y(n_494) );
BUFx2_ASAP7_75t_L g614 ( .A(n_486), .Y(n_614) );
INVx1_ASAP7_75t_L g1104 ( .A(n_486), .Y(n_1104) );
BUFx2_ASAP7_75t_L g1411 ( .A(n_486), .Y(n_1411) );
AND2x2_ASAP7_75t_L g908 ( .A(n_487), .B(n_909), .Y(n_908) );
HB1xp67_ASAP7_75t_L g962 ( .A(n_487), .Y(n_962) );
OAI22xp5_ASAP7_75t_L g611 ( .A1(n_488), .A2(n_593), .B1(n_606), .B2(n_612), .Y(n_611) );
OAI22xp5_ASAP7_75t_L g672 ( .A1(n_488), .A2(n_645), .B1(n_665), .B2(n_673), .Y(n_672) );
OAI22xp5_ASAP7_75t_L g721 ( .A1(n_488), .A2(n_673), .B1(n_722), .B2(n_723), .Y(n_721) );
OAI22xp5_ASAP7_75t_L g1529 ( .A1(n_488), .A2(n_824), .B1(n_1530), .B2(n_1531), .Y(n_1529) );
INVx5_ASAP7_75t_L g488 ( .A(n_489), .Y(n_488) );
INVx2_ASAP7_75t_SL g489 ( .A(n_490), .Y(n_489) );
BUFx2_ASAP7_75t_SL g676 ( .A(n_490), .Y(n_676) );
BUFx3_ASAP7_75t_L g891 ( .A(n_490), .Y(n_891) );
OR2x2_ASAP7_75t_L g1086 ( .A(n_490), .B(n_1085), .Y(n_1086) );
NAND2xp5_ASAP7_75t_L g1211 ( .A(n_490), .B(n_1212), .Y(n_1211) );
NAND2xp5_ASAP7_75t_L g1318 ( .A(n_490), .B(n_1319), .Y(n_1318) );
BUFx3_ASAP7_75t_L g490 ( .A(n_491), .Y(n_490) );
BUFx6f_ASAP7_75t_L g567 ( .A(n_491), .Y(n_567) );
HB1xp67_ASAP7_75t_L g493 ( .A(n_494), .Y(n_493) );
OAI22xp5_ASAP7_75t_L g609 ( .A1(n_494), .A2(n_595), .B1(n_598), .B2(n_610), .Y(n_609) );
INVx2_ASAP7_75t_L g825 ( .A(n_494), .Y(n_825) );
OAI21xp33_ASAP7_75t_L g1215 ( .A1(n_494), .A2(n_497), .B(n_1216), .Y(n_1215) );
OAI221xp5_ASAP7_75t_L g1323 ( .A1(n_494), .A2(n_497), .B1(n_567), .B2(n_1324), .C(n_1325), .Y(n_1323) );
OAI33xp33_ASAP7_75t_L g667 ( .A1(n_495), .A2(n_668), .A3(n_671), .B1(n_672), .B2(n_674), .B3(n_677), .Y(n_667) );
OAI33xp33_ASAP7_75t_L g873 ( .A1(n_495), .A2(n_874), .A3(n_875), .B1(n_876), .B2(n_877), .B3(n_878), .Y(n_873) );
INVx2_ASAP7_75t_L g495 ( .A(n_496), .Y(n_495) );
CKINVDCx5p33_ASAP7_75t_R g728 ( .A(n_496), .Y(n_728) );
NAND3xp33_ASAP7_75t_L g1360 ( .A(n_496), .B(n_1361), .C(n_1367), .Y(n_1360) );
AOI33xp33_ASAP7_75t_L g1590 ( .A1(n_496), .A2(n_1591), .A3(n_1594), .B1(n_1597), .B2(n_1599), .B3(n_1600), .Y(n_1590) );
AND2x4_ASAP7_75t_L g496 ( .A(n_497), .B(n_498), .Y(n_496) );
NAND2xp5_ASAP7_75t_L g831 ( .A(n_497), .B(n_498), .Y(n_831) );
INVx4_ASAP7_75t_L g981 ( .A(n_497), .Y(n_981) );
INVx1_ASAP7_75t_SL g1641 ( .A(n_497), .Y(n_1641) );
INVx1_ASAP7_75t_L g498 ( .A(n_499), .Y(n_498) );
OAI22xp33_ASAP7_75t_L g615 ( .A1(n_501), .A2(n_596), .B1(n_601), .B2(n_616), .Y(n_615) );
OAI22xp33_ASAP7_75t_L g878 ( .A1(n_501), .A2(n_790), .B1(n_858), .B2(n_868), .Y(n_878) );
INVx1_ASAP7_75t_L g501 ( .A(n_502), .Y(n_501) );
INVx1_ASAP7_75t_L g502 ( .A(n_503), .Y(n_502) );
INVx1_ASAP7_75t_L g503 ( .A(n_504), .Y(n_503) );
OAI22xp5_ASAP7_75t_L g832 ( .A1(n_505), .A2(n_815), .B1(n_833), .B2(n_834), .Y(n_832) );
OAI22xp5_ASAP7_75t_L g1532 ( .A1(n_505), .A2(n_815), .B1(n_1533), .B2(n_1534), .Y(n_1532) );
BUFx3_ASAP7_75t_L g505 ( .A(n_506), .Y(n_505) );
OAI31xp33_ASAP7_75t_L g507 ( .A1(n_508), .A2(n_514), .A3(n_533), .B(n_540), .Y(n_507) );
BUFx2_ASAP7_75t_L g509 ( .A(n_510), .Y(n_509) );
INVx2_ASAP7_75t_SL g627 ( .A(n_510), .Y(n_627) );
BUFx3_ASAP7_75t_L g763 ( .A(n_510), .Y(n_763) );
BUFx2_ASAP7_75t_L g803 ( .A(n_510), .Y(n_803) );
AND2x4_ASAP7_75t_L g538 ( .A(n_511), .B(n_539), .Y(n_538) );
BUFx3_ASAP7_75t_L g512 ( .A(n_513), .Y(n_512) );
INVx1_ASAP7_75t_L g693 ( .A(n_513), .Y(n_693) );
INVx2_ASAP7_75t_L g765 ( .A(n_513), .Y(n_765) );
INVx1_ASAP7_75t_L g1936 ( .A(n_513), .Y(n_1936) );
INVxp67_ASAP7_75t_L g515 ( .A(n_516), .Y(n_515) );
INVx1_ASAP7_75t_L g745 ( .A(n_516), .Y(n_745) );
INVx1_ASAP7_75t_L g1396 ( .A(n_516), .Y(n_1396) );
INVx1_ASAP7_75t_L g516 ( .A(n_517), .Y(n_516) );
INVx1_ASAP7_75t_L g621 ( .A(n_517), .Y(n_621) );
CKINVDCx8_ASAP7_75t_R g518 ( .A(n_519), .Y(n_518) );
CKINVDCx8_ASAP7_75t_R g757 ( .A(n_519), .Y(n_757) );
OAI31xp33_ASAP7_75t_L g1267 ( .A1(n_519), .A2(n_1268), .A3(n_1278), .B(n_1279), .Y(n_1267) );
AOI211xp5_ASAP7_75t_L g1575 ( .A1(n_519), .A2(n_1287), .B(n_1573), .C(n_1576), .Y(n_1575) );
BUFx2_ASAP7_75t_L g1013 ( .A(n_520), .Y(n_1013) );
BUFx3_ASAP7_75t_L g1132 ( .A(n_520), .Y(n_1132) );
BUFx2_ASAP7_75t_L g1141 ( .A(n_520), .Y(n_1141) );
INVx2_ASAP7_75t_L g1183 ( .A(n_520), .Y(n_1183) );
BUFx2_ASAP7_75t_L g1265 ( .A(n_520), .Y(n_1265) );
BUFx2_ASAP7_75t_L g1299 ( .A(n_520), .Y(n_1299) );
INVx1_ASAP7_75t_L g944 ( .A(n_521), .Y(n_944) );
AOI22xp33_ASAP7_75t_L g522 ( .A1(n_523), .A2(n_528), .B1(n_529), .B2(n_532), .Y(n_522) );
AOI22xp33_ASAP7_75t_L g622 ( .A1(n_523), .A2(n_529), .B1(n_623), .B2(n_624), .Y(n_622) );
AOI22xp33_ASAP7_75t_L g1064 ( .A1(n_523), .A2(n_529), .B1(n_1021), .B2(n_1065), .Y(n_1064) );
AOI22xp33_ASAP7_75t_L g1348 ( .A1(n_523), .A2(n_529), .B1(n_1341), .B2(n_1343), .Y(n_1348) );
AOI22xp33_ASAP7_75t_L g1488 ( .A1(n_523), .A2(n_529), .B1(n_1482), .B2(n_1489), .Y(n_1488) );
AOI22xp33_ASAP7_75t_L g1912 ( .A1(n_523), .A2(n_529), .B1(n_1905), .B2(n_1913), .Y(n_1912) );
BUFx3_ASAP7_75t_L g523 ( .A(n_524), .Y(n_523) );
BUFx3_ASAP7_75t_L g688 ( .A(n_524), .Y(n_688) );
AND2x2_ASAP7_75t_L g524 ( .A(n_525), .B(n_527), .Y(n_524) );
AND2x4_ASAP7_75t_L g530 ( .A(n_525), .B(n_531), .Y(n_530) );
AND2x4_ASAP7_75t_L g759 ( .A(n_525), .B(n_527), .Y(n_759) );
A2O1A1Ixp33_ASAP7_75t_L g1268 ( .A1(n_525), .A2(n_1269), .B(n_1272), .C(n_1275), .Y(n_1268) );
INVx3_ASAP7_75t_L g525 ( .A(n_526), .Y(n_525) );
AOI22xp33_ASAP7_75t_L g573 ( .A1(n_528), .A2(n_574), .B1(n_577), .B2(n_582), .Y(n_573) );
AOI22xp33_ASAP7_75t_L g687 ( .A1(n_529), .A2(n_688), .B1(n_689), .B2(n_690), .Y(n_687) );
BUFx6f_ASAP7_75t_L g529 ( .A(n_530), .Y(n_529) );
AOI22xp33_ASAP7_75t_L g758 ( .A1(n_530), .A2(n_759), .B1(n_760), .B2(n_761), .Y(n_758) );
AOI22xp33_ASAP7_75t_L g806 ( .A1(n_530), .A2(n_759), .B1(n_794), .B2(n_807), .Y(n_806) );
AOI22xp33_ASAP7_75t_L g882 ( .A1(n_530), .A2(n_759), .B1(n_883), .B2(n_884), .Y(n_882) );
AOI22xp5_ASAP7_75t_L g1275 ( .A1(n_530), .A2(n_759), .B1(n_1276), .B2(n_1277), .Y(n_1275) );
AOI22xp33_ASAP7_75t_SL g1432 ( .A1(n_530), .A2(n_759), .B1(n_1424), .B2(n_1433), .Y(n_1432) );
AOI22xp33_ASAP7_75t_L g1448 ( .A1(n_530), .A2(n_759), .B1(n_1439), .B2(n_1449), .Y(n_1448) );
AOI22xp33_ASAP7_75t_L g1544 ( .A1(n_530), .A2(n_759), .B1(n_1545), .B2(n_1546), .Y(n_1544) );
INVx1_ASAP7_75t_L g1578 ( .A(n_530), .Y(n_1578) );
AOI22xp33_ASAP7_75t_SL g1931 ( .A1(n_530), .A2(n_688), .B1(n_1932), .B2(n_1933), .Y(n_1931) );
INVx2_ASAP7_75t_L g534 ( .A(n_535), .Y(n_534) );
AOI22xp33_ASAP7_75t_L g1581 ( .A1(n_535), .A2(n_538), .B1(n_1568), .B2(n_1569), .Y(n_1581) );
INVx2_ASAP7_75t_SL g535 ( .A(n_536), .Y(n_535) );
HB1xp67_ASAP7_75t_L g629 ( .A(n_536), .Y(n_629) );
INVx1_ASAP7_75t_L g683 ( .A(n_536), .Y(n_683) );
INVx2_ASAP7_75t_SL g1061 ( .A(n_536), .Y(n_1061) );
INVx1_ASAP7_75t_L g537 ( .A(n_538), .Y(n_537) );
INVx1_ASAP7_75t_L g630 ( .A(n_538), .Y(n_630) );
INVx2_ASAP7_75t_L g684 ( .A(n_538), .Y(n_684) );
INVxp67_ASAP7_75t_L g753 ( .A(n_538), .Y(n_753) );
INVx1_ASAP7_75t_L g809 ( .A(n_538), .Y(n_809) );
INVx2_ASAP7_75t_L g1062 ( .A(n_538), .Y(n_1062) );
BUFx6f_ASAP7_75t_L g742 ( .A(n_539), .Y(n_742) );
INVx2_ASAP7_75t_L g749 ( .A(n_539), .Y(n_749) );
BUFx6f_ASAP7_75t_L g1151 ( .A(n_539), .Y(n_1151) );
INVx2_ASAP7_75t_L g1884 ( .A(n_539), .Y(n_1884) );
OAI31xp33_ASAP7_75t_L g680 ( .A1(n_540), .A2(n_681), .A3(n_685), .B(n_691), .Y(n_680) );
AND2x2_ASAP7_75t_L g540 ( .A(n_541), .B(n_543), .Y(n_540) );
AND2x4_ASAP7_75t_L g631 ( .A(n_541), .B(n_543), .Y(n_631) );
AND2x2_ASAP7_75t_L g766 ( .A(n_541), .B(n_543), .Y(n_766) );
AND2x2_ASAP7_75t_SL g810 ( .A(n_541), .B(n_543), .Y(n_810) );
AND2x2_ASAP7_75t_L g1279 ( .A(n_541), .B(n_543), .Y(n_1279) );
INVx1_ASAP7_75t_SL g541 ( .A(n_542), .Y(n_541) );
INVx1_ASAP7_75t_L g543 ( .A(n_544), .Y(n_543) );
OAI31xp33_ASAP7_75t_SL g545 ( .A1(n_546), .A2(n_554), .A3(n_563), .B(n_583), .Y(n_545) );
INVx3_ASAP7_75t_SL g548 ( .A(n_549), .Y(n_548) );
CKINVDCx16_ASAP7_75t_R g634 ( .A(n_549), .Y(n_634) );
INVx4_ASAP7_75t_L g800 ( .A(n_549), .Y(n_800) );
AND2x4_ASAP7_75t_L g549 ( .A(n_550), .B(n_552), .Y(n_549) );
HB1xp67_ASAP7_75t_L g550 ( .A(n_551), .Y(n_550) );
BUFx6f_ASAP7_75t_L g923 ( .A(n_552), .Y(n_923) );
BUFx3_ASAP7_75t_L g968 ( .A(n_552), .Y(n_968) );
INVx2_ASAP7_75t_L g1092 ( .A(n_552), .Y(n_1092) );
INVx1_ASAP7_75t_L g555 ( .A(n_556), .Y(n_555) );
INVx1_ASAP7_75t_L g556 ( .A(n_557), .Y(n_556) );
BUFx6f_ASAP7_75t_L g704 ( .A(n_557), .Y(n_704) );
HB1xp67_ASAP7_75t_L g1026 ( .A(n_557), .Y(n_1026) );
BUFx2_ASAP7_75t_L g1942 ( .A(n_557), .Y(n_1942) );
INVx1_ASAP7_75t_L g558 ( .A(n_559), .Y(n_558) );
INVx2_ASAP7_75t_SL g559 ( .A(n_560), .Y(n_559) );
HB1xp67_ASAP7_75t_L g1553 ( .A(n_560), .Y(n_1553) );
BUFx2_ASAP7_75t_L g560 ( .A(n_561), .Y(n_560) );
INVx2_ASAP7_75t_L g706 ( .A(n_561), .Y(n_706) );
INVx1_ASAP7_75t_L g798 ( .A(n_561), .Y(n_798) );
AND2x4_ASAP7_75t_L g575 ( .A(n_562), .B(n_576), .Y(n_575) );
AND2x2_ASAP7_75t_L g699 ( .A(n_562), .B(n_576), .Y(n_699) );
AND2x2_ASAP7_75t_L g1334 ( .A(n_562), .B(n_955), .Y(n_1334) );
INVx1_ASAP7_75t_L g564 ( .A(n_565), .Y(n_564) );
INVx1_ASAP7_75t_L g565 ( .A(n_566), .Y(n_565) );
OAI22xp5_ASAP7_75t_L g724 ( .A1(n_566), .A2(n_725), .B1(n_726), .B2(n_727), .Y(n_724) );
OAI22xp5_ASAP7_75t_L g1410 ( .A1(n_566), .A2(n_1398), .B1(n_1402), .B2(n_1411), .Y(n_1410) );
OAI22xp5_ASAP7_75t_L g1949 ( .A1(n_566), .A2(n_824), .B1(n_1950), .B2(n_1951), .Y(n_1949) );
BUFx4f_ASAP7_75t_L g566 ( .A(n_567), .Y(n_566) );
BUFx4f_ASAP7_75t_L g610 ( .A(n_567), .Y(n_610) );
BUFx4f_ASAP7_75t_L g773 ( .A(n_567), .Y(n_773) );
INVx4_ASAP7_75t_L g791 ( .A(n_567), .Y(n_791) );
BUFx4f_ASAP7_75t_L g1105 ( .A(n_567), .Y(n_1105) );
OR2x6_ASAP7_75t_L g1109 ( .A(n_567), .B(n_1110), .Y(n_1109) );
BUFx6f_ASAP7_75t_L g1253 ( .A(n_567), .Y(n_1253) );
INVx1_ASAP7_75t_L g568 ( .A(n_569), .Y(n_568) );
INVx1_ASAP7_75t_L g697 ( .A(n_569), .Y(n_697) );
INVx3_ASAP7_75t_L g792 ( .A(n_569), .Y(n_792) );
AND2x2_ASAP7_75t_L g569 ( .A(n_570), .B(n_571), .Y(n_569) );
AND2x2_ASAP7_75t_L g775 ( .A(n_570), .B(n_776), .Y(n_775) );
AND2x4_ASAP7_75t_SL g991 ( .A(n_571), .B(n_907), .Y(n_991) );
BUFx6f_ASAP7_75t_L g1094 ( .A(n_571), .Y(n_1094) );
BUFx3_ASAP7_75t_L g1214 ( .A(n_571), .Y(n_1214) );
BUFx3_ASAP7_75t_L g1342 ( .A(n_571), .Y(n_1342) );
AND2x6_ASAP7_75t_L g1644 ( .A(n_571), .B(n_964), .Y(n_1644) );
BUFx6f_ASAP7_75t_L g571 ( .A(n_572), .Y(n_571) );
INVx1_ASAP7_75t_L g777 ( .A(n_572), .Y(n_777) );
AOI22xp33_ASAP7_75t_L g637 ( .A1(n_574), .A2(n_577), .B1(n_623), .B2(n_638), .Y(n_637) );
AOI22xp33_ASAP7_75t_L g793 ( .A1(n_574), .A2(n_700), .B1(n_794), .B2(n_795), .Y(n_793) );
AOI22xp33_ASAP7_75t_L g892 ( .A1(n_574), .A2(n_883), .B1(n_893), .B2(n_894), .Y(n_892) );
AOI22xp33_ASAP7_75t_L g1020 ( .A1(n_574), .A2(n_893), .B1(n_1021), .B2(n_1022), .Y(n_1020) );
AOI22xp33_ASAP7_75t_L g1481 ( .A1(n_574), .A2(n_893), .B1(n_1482), .B2(n_1483), .Y(n_1481) );
AOI22xp33_ASAP7_75t_L g1550 ( .A1(n_574), .A2(n_893), .B1(n_1545), .B2(n_1551), .Y(n_1550) );
BUFx3_ASAP7_75t_L g574 ( .A(n_575), .Y(n_574) );
AOI22xp33_ASAP7_75t_L g778 ( .A1(n_575), .A2(n_579), .B1(n_760), .B2(n_779), .Y(n_778) );
AOI22xp33_ASAP7_75t_L g1438 ( .A1(n_575), .A2(n_579), .B1(n_1439), .B2(n_1440), .Y(n_1438) );
AOI222xp33_ASAP7_75t_L g1570 ( .A1(n_575), .A2(n_1214), .B1(n_1340), .B2(n_1571), .C1(n_1572), .C2(n_1573), .Y(n_1570) );
AOI22xp33_ASAP7_75t_L g1904 ( .A1(n_575), .A2(n_1340), .B1(n_1905), .B2(n_1906), .Y(n_1904) );
BUFx2_ASAP7_75t_L g959 ( .A(n_576), .Y(n_959) );
INVx1_ASAP7_75t_L g1116 ( .A(n_576), .Y(n_1116) );
AOI22xp33_ASAP7_75t_L g1212 ( .A1(n_576), .A2(n_961), .B1(n_1166), .B2(n_1191), .Y(n_1212) );
INVx1_ASAP7_75t_L g1251 ( .A(n_576), .Y(n_1251) );
AOI22xp33_ASAP7_75t_L g1939 ( .A1(n_577), .A2(n_699), .B1(n_1932), .B2(n_1940), .Y(n_1939) );
INVx2_ASAP7_75t_L g577 ( .A(n_578), .Y(n_577) );
INVx2_ASAP7_75t_L g1340 ( .A(n_578), .Y(n_1340) );
INVx2_ASAP7_75t_L g578 ( .A(n_579), .Y(n_578) );
INVx2_ASAP7_75t_L g701 ( .A(n_579), .Y(n_701) );
BUFx3_ASAP7_75t_L g893 ( .A(n_579), .Y(n_893) );
NAND2xp5_ASAP7_75t_L g1118 ( .A(n_580), .B(n_964), .Y(n_1118) );
INVx1_ASAP7_75t_L g580 ( .A(n_581), .Y(n_580) );
OAI31xp33_ASAP7_75t_L g632 ( .A1(n_583), .A2(n_633), .A3(n_635), .B(n_636), .Y(n_632) );
OAI31xp33_ASAP7_75t_L g886 ( .A1(n_583), .A2(n_887), .A3(n_888), .B(n_889), .Y(n_886) );
OAI31xp33_ASAP7_75t_L g1436 ( .A1(n_583), .A2(n_1437), .A3(n_1441), .B(n_1443), .Y(n_1436) );
OAI31xp33_ASAP7_75t_L g1548 ( .A1(n_583), .A2(n_1549), .A3(n_1552), .B(n_1554), .Y(n_1548) );
OAI31xp33_ASAP7_75t_L g1937 ( .A1(n_583), .A2(n_1938), .A3(n_1941), .B(n_1943), .Y(n_1937) );
BUFx2_ASAP7_75t_SL g583 ( .A(n_584), .Y(n_583) );
BUFx3_ASAP7_75t_L g707 ( .A(n_584), .Y(n_707) );
BUFx2_ASAP7_75t_L g782 ( .A(n_584), .Y(n_782) );
OAI31xp33_ASAP7_75t_L g1018 ( .A1(n_584), .A2(n_1019), .A3(n_1023), .B(n_1025), .Y(n_1018) );
INVx1_ASAP7_75t_L g1475 ( .A(n_584), .Y(n_1475) );
AOI22xp5_ASAP7_75t_L g1562 ( .A1(n_584), .A2(n_631), .B1(n_1563), .B2(n_1574), .Y(n_1562) );
INVx1_ASAP7_75t_L g585 ( .A(n_586), .Y(n_585) );
INVx1_ASAP7_75t_L g905 ( .A(n_586), .Y(n_905) );
INVxp67_ASAP7_75t_L g930 ( .A(n_586), .Y(n_930) );
OR2x2_ASAP7_75t_L g1117 ( .A(n_586), .B(n_1118), .Y(n_1117) );
AND3x1_ASAP7_75t_L g588 ( .A(n_589), .B(n_617), .C(n_632), .Y(n_588) );
NOR2xp33_ASAP7_75t_L g589 ( .A(n_590), .B(n_607), .Y(n_589) );
INVx3_ASAP7_75t_L g599 ( .A(n_600), .Y(n_599) );
INVx3_ASAP7_75t_L g840 ( .A(n_600), .Y(n_840) );
INVx2_ASAP7_75t_SL g1006 ( .A(n_600), .Y(n_1006) );
AND2x4_ASAP7_75t_L g1187 ( .A(n_600), .B(n_1169), .Y(n_1187) );
INVx2_ASAP7_75t_SL g1403 ( .A(n_600), .Y(n_1403) );
OAI22xp5_ASAP7_75t_L g651 ( .A1(n_604), .A2(n_652), .B1(n_653), .B2(n_655), .Y(n_651) );
OAI22xp33_ASAP7_75t_L g658 ( .A1(n_604), .A2(n_659), .B1(n_660), .B2(n_661), .Y(n_658) );
OAI22xp33_ASAP7_75t_L g836 ( .A1(n_604), .A2(n_814), .B1(n_826), .B2(n_837), .Y(n_836) );
OAI22xp5_ASAP7_75t_L g1044 ( .A1(n_604), .A2(n_1031), .B1(n_1045), .B2(n_1046), .Y(n_1044) );
OAI22xp33_ASAP7_75t_L g1509 ( .A1(n_604), .A2(n_1495), .B1(n_1503), .B2(n_1510), .Y(n_1509) );
INVx2_ASAP7_75t_L g604 ( .A(n_605), .Y(n_604) );
INVx1_ASAP7_75t_L g1431 ( .A(n_605), .Y(n_1431) );
OAI22xp5_ASAP7_75t_L g876 ( .A1(n_610), .A2(n_612), .B1(n_857), .B2(n_864), .Y(n_876) );
OAI22xp5_ASAP7_75t_L g1526 ( .A1(n_610), .A2(n_612), .B1(n_1527), .B2(n_1528), .Y(n_1526) );
OAI22xp5_ASAP7_75t_L g820 ( .A1(n_612), .A2(n_773), .B1(n_821), .B2(n_822), .Y(n_820) );
INVx2_ASAP7_75t_L g612 ( .A(n_613), .Y(n_612) );
INVx4_ASAP7_75t_L g673 ( .A(n_613), .Y(n_673) );
INVx2_ASAP7_75t_L g675 ( .A(n_613), .Y(n_675) );
INVx2_ASAP7_75t_L g726 ( .A(n_613), .Y(n_726) );
INVx4_ASAP7_75t_L g613 ( .A(n_614), .Y(n_613) );
OAI22xp33_ASAP7_75t_L g1463 ( .A1(n_616), .A2(n_669), .B1(n_1464), .B2(n_1465), .Y(n_1463) );
OAI22xp5_ASAP7_75t_L g1955 ( .A1(n_616), .A2(n_669), .B1(n_1956), .B2(n_1957), .Y(n_1955) );
OAI31xp33_ASAP7_75t_L g617 ( .A1(n_618), .A2(n_625), .A3(n_628), .B(n_631), .Y(n_617) );
HB1xp67_ASAP7_75t_L g619 ( .A(n_620), .Y(n_619) );
INVxp67_ASAP7_75t_SL g620 ( .A(n_621), .Y(n_620) );
INVx1_ASAP7_75t_L g686 ( .A(n_621), .Y(n_686) );
INVxp67_ASAP7_75t_SL g1408 ( .A(n_621), .Y(n_1408) );
INVx2_ASAP7_75t_L g626 ( .A(n_627), .Y(n_626) );
INVx1_ASAP7_75t_L g1067 ( .A(n_627), .Y(n_1067) );
OAI31xp33_ASAP7_75t_L g1345 ( .A1(n_631), .A2(n_1346), .A3(n_1347), .B(n_1349), .Y(n_1345) );
CKINVDCx14_ASAP7_75t_R g1491 ( .A(n_631), .Y(n_1491) );
OAI31xp33_ASAP7_75t_L g1541 ( .A1(n_631), .A2(n_1542), .A3(n_1543), .B(n_1547), .Y(n_1541) );
OAI31xp33_ASAP7_75t_L g1927 ( .A1(n_631), .A2(n_1928), .A3(n_1929), .B(n_1934), .Y(n_1927) );
OA22x2_ASAP7_75t_L g639 ( .A1(n_640), .A2(n_708), .B1(n_709), .B2(n_783), .Y(n_639) );
INVx1_ASAP7_75t_L g783 ( .A(n_640), .Y(n_783) );
NAND3xp33_ASAP7_75t_L g641 ( .A(n_642), .B(n_680), .C(n_694), .Y(n_641) );
NOR2xp33_ASAP7_75t_L g642 ( .A(n_643), .B(n_667), .Y(n_642) );
OAI33xp33_ASAP7_75t_L g643 ( .A1(n_644), .A2(n_651), .A3(n_656), .B1(n_658), .B2(n_662), .B3(n_663), .Y(n_643) );
OAI22xp33_ASAP7_75t_SL g644 ( .A1(n_645), .A2(n_646), .B1(n_647), .B2(n_648), .Y(n_644) );
OAI22xp5_ASAP7_75t_L g1961 ( .A1(n_648), .A2(n_1150), .B1(n_1950), .B2(n_1956), .Y(n_1961) );
INVx3_ASAP7_75t_L g648 ( .A(n_649), .Y(n_648) );
BUFx2_ASAP7_75t_L g649 ( .A(n_650), .Y(n_649) );
INVx1_ASAP7_75t_L g859 ( .A(n_650), .Y(n_859) );
OAI22xp33_ASAP7_75t_L g668 ( .A1(n_652), .A2(n_659), .B1(n_669), .B2(n_670), .Y(n_668) );
OAI22xp33_ASAP7_75t_L g736 ( .A1(n_653), .A2(n_717), .B1(n_725), .B2(n_737), .Y(n_736) );
OAI22xp33_ASAP7_75t_L g744 ( .A1(n_653), .A2(n_718), .B1(n_727), .B2(n_745), .Y(n_744) );
BUFx4f_ASAP7_75t_SL g1002 ( .A(n_653), .Y(n_1002) );
OAI22xp33_ASAP7_75t_L g1467 ( .A1(n_653), .A2(n_755), .B1(n_1454), .B2(n_1461), .Y(n_1467) );
INVx3_ASAP7_75t_L g653 ( .A(n_654), .Y(n_653) );
INVx2_ASAP7_75t_SL g837 ( .A(n_654), .Y(n_837) );
OAI22xp5_ASAP7_75t_L g674 ( .A1(n_655), .A2(n_661), .B1(n_675), .B2(n_676), .Y(n_674) );
OAI33xp33_ASAP7_75t_L g1028 ( .A1(n_656), .A2(n_1029), .A3(n_1034), .B1(n_1038), .B2(n_1041), .B3(n_1044), .Y(n_1028) );
OAI22xp33_ASAP7_75t_L g1254 ( .A1(n_656), .A2(n_1255), .B1(n_1261), .B2(n_1266), .Y(n_1254) );
BUFx3_ASAP7_75t_L g656 ( .A(n_657), .Y(n_656) );
OAI221xp5_ASAP7_75t_L g1146 ( .A1(n_660), .A2(n_1098), .B1(n_1106), .B2(n_1147), .C(n_1148), .Y(n_1146) );
OAI22xp33_ASAP7_75t_L g1405 ( .A1(n_660), .A2(n_1406), .B1(n_1407), .B2(n_1408), .Y(n_1405) );
OAI22xp33_ASAP7_75t_L g716 ( .A1(n_669), .A2(n_717), .B1(n_718), .B2(n_719), .Y(n_716) );
OAI22xp5_ASAP7_75t_L g1414 ( .A1(n_669), .A2(n_1399), .B1(n_1404), .B2(n_1415), .Y(n_1414) );
OAI33xp33_ASAP7_75t_L g812 ( .A1(n_671), .A2(n_813), .A3(n_820), .B1(n_823), .B2(n_829), .B3(n_832), .Y(n_812) );
OAI33xp33_ASAP7_75t_L g1047 ( .A1(n_671), .A2(n_829), .A3(n_1048), .B1(n_1055), .B2(n_1056), .B3(n_1057), .Y(n_1047) );
INVx1_ASAP7_75t_L g1099 ( .A(n_671), .Y(n_1099) );
OAI22xp5_ASAP7_75t_L g1418 ( .A1(n_673), .A2(n_827), .B1(n_1395), .B2(n_1407), .Y(n_1418) );
OAI22xp5_ASAP7_75t_L g1460 ( .A1(n_673), .A2(n_827), .B1(n_1461), .B2(n_1462), .Y(n_1460) );
OAI22xp5_ASAP7_75t_L g1952 ( .A1(n_673), .A2(n_1105), .B1(n_1953), .B2(n_1954), .Y(n_1952) );
OAI22xp33_ASAP7_75t_L g1946 ( .A1(n_678), .A2(n_733), .B1(n_1947), .B2(n_1948), .Y(n_1946) );
BUFx3_ASAP7_75t_L g678 ( .A(n_679), .Y(n_678) );
BUFx3_ASAP7_75t_L g1097 ( .A(n_679), .Y(n_1097) );
BUFx6f_ASAP7_75t_L g1413 ( .A(n_679), .Y(n_1413) );
INVx1_ASAP7_75t_L g682 ( .A(n_683), .Y(n_682) );
AOI22xp33_ASAP7_75t_L g698 ( .A1(n_689), .A2(n_699), .B1(n_700), .B2(n_702), .Y(n_698) );
INVx1_ASAP7_75t_L g692 ( .A(n_693), .Y(n_692) );
OAI31xp33_ASAP7_75t_L g694 ( .A1(n_695), .A2(n_696), .A3(n_703), .B(n_707), .Y(n_694) );
AOI222xp33_ASAP7_75t_L g1338 ( .A1(n_699), .A2(n_1339), .B1(n_1340), .B2(n_1341), .C1(n_1342), .C2(n_1343), .Y(n_1338) );
AOI22xp33_ASAP7_75t_L g1423 ( .A1(n_699), .A2(n_1340), .B1(n_1424), .B2(n_1425), .Y(n_1423) );
INVx2_ASAP7_75t_L g700 ( .A(n_701), .Y(n_700) );
INVx1_ASAP7_75t_L g705 ( .A(n_706), .Y(n_705) );
INVx1_ASAP7_75t_L g781 ( .A(n_706), .Y(n_781) );
INVx2_ASAP7_75t_L g1442 ( .A(n_706), .Y(n_1442) );
OAI31xp33_ASAP7_75t_L g788 ( .A1(n_707), .A2(n_789), .A3(n_796), .B(n_799), .Y(n_788) );
OAI31xp33_ASAP7_75t_L g1902 ( .A1(n_707), .A2(n_1903), .A3(n_1907), .B(n_1908), .Y(n_1902) );
INVx2_ASAP7_75t_SL g708 ( .A(n_709), .Y(n_708) );
NAND3xp33_ASAP7_75t_L g710 ( .A(n_711), .B(n_751), .C(n_767), .Y(n_710) );
NOR2xp33_ASAP7_75t_L g711 ( .A(n_712), .B(n_734), .Y(n_711) );
OAI33xp33_ASAP7_75t_L g712 ( .A1(n_713), .A2(n_716), .A3(n_721), .B1(n_724), .B2(n_728), .B3(n_729), .Y(n_712) );
OAI33xp33_ASAP7_75t_L g1945 ( .A1(n_713), .A2(n_728), .A3(n_1946), .B1(n_1949), .B2(n_1952), .B3(n_1955), .Y(n_1945) );
INVx1_ASAP7_75t_L g713 ( .A(n_714), .Y(n_713) );
INVx2_ASAP7_75t_SL g714 ( .A(n_715), .Y(n_714) );
INVx2_ASAP7_75t_SL g1359 ( .A(n_715), .Y(n_1359) );
OAI33xp33_ASAP7_75t_L g1522 ( .A1(n_715), .A2(n_831), .A3(n_1523), .B1(n_1526), .B2(n_1529), .B3(n_1532), .Y(n_1522) );
OAI22xp5_ASAP7_75t_L g1095 ( .A1(n_719), .A2(n_1096), .B1(n_1097), .B2(n_1098), .Y(n_1095) );
BUFx6f_ASAP7_75t_L g719 ( .A(n_720), .Y(n_719) );
OAI22xp5_ASAP7_75t_L g740 ( .A1(n_722), .A2(n_730), .B1(n_741), .B2(n_743), .Y(n_740) );
OAI22xp5_ASAP7_75t_L g748 ( .A1(n_723), .A2(n_732), .B1(n_749), .B2(n_750), .Y(n_748) );
OAI21xp5_ASAP7_75t_L g1100 ( .A1(n_728), .A2(n_1101), .B(n_1109), .Y(n_1100) );
OAI22xp5_ASAP7_75t_L g729 ( .A1(n_730), .A2(n_731), .B1(n_732), .B2(n_733), .Y(n_729) );
OAI33xp33_ASAP7_75t_L g734 ( .A1(n_735), .A2(n_736), .A3(n_740), .B1(n_744), .B2(n_746), .B3(n_748), .Y(n_734) );
OAI33xp33_ASAP7_75t_L g1958 ( .A1(n_735), .A2(n_1890), .A3(n_1959), .B1(n_1961), .B2(n_1962), .B3(n_1963), .Y(n_1958) );
INVx1_ASAP7_75t_L g737 ( .A(n_738), .Y(n_737) );
INVx2_ASAP7_75t_L g1003 ( .A(n_738), .Y(n_1003) );
INVx2_ASAP7_75t_L g1147 ( .A(n_738), .Y(n_1147) );
INVx1_ASAP7_75t_L g1487 ( .A(n_738), .Y(n_1487) );
INVx1_ASAP7_75t_L g1960 ( .A(n_738), .Y(n_1960) );
INVx4_ASAP7_75t_L g738 ( .A(n_739), .Y(n_738) );
INVx3_ASAP7_75t_L g756 ( .A(n_739), .Y(n_756) );
BUFx6f_ASAP7_75t_L g867 ( .A(n_739), .Y(n_867) );
OR2x2_ASAP7_75t_L g949 ( .A(n_739), .B(n_913), .Y(n_949) );
INVx1_ASAP7_75t_L g741 ( .A(n_742), .Y(n_741) );
OAI22xp5_ASAP7_75t_L g839 ( .A1(n_743), .A2(n_822), .B1(n_834), .B2(n_840), .Y(n_839) );
OAI22xp5_ASAP7_75t_L g1401 ( .A1(n_743), .A2(n_1402), .B1(n_1403), .B2(n_1404), .Y(n_1401) );
OAI22xp5_ASAP7_75t_L g1469 ( .A1(n_743), .A2(n_1403), .B1(n_1459), .B2(n_1465), .Y(n_1469) );
OAI22xp5_ASAP7_75t_L g1513 ( .A1(n_743), .A2(n_1501), .B1(n_1507), .B2(n_1514), .Y(n_1513) );
INVx1_ASAP7_75t_L g1184 ( .A(n_746), .Y(n_1184) );
OAI33xp33_ASAP7_75t_L g1391 ( .A1(n_746), .A2(n_1392), .A3(n_1393), .B1(n_1397), .B2(n_1401), .B3(n_1405), .Y(n_1391) );
OAI33xp33_ASAP7_75t_L g1466 ( .A1(n_746), .A2(n_1392), .A3(n_1467), .B1(n_1468), .B2(n_1469), .B3(n_1470), .Y(n_1466) );
INVx3_ASAP7_75t_L g1148 ( .A(n_747), .Y(n_1148) );
OAI22xp5_ASAP7_75t_L g1149 ( .A1(n_750), .A2(n_1150), .B1(n_1152), .B2(n_1153), .Y(n_1149) );
OAI221xp5_ASAP7_75t_L g1255 ( .A1(n_750), .A2(n_1256), .B1(n_1257), .B2(n_1258), .C(n_1259), .Y(n_1255) );
OAI221xp5_ASAP7_75t_L g1261 ( .A1(n_750), .A2(n_1241), .B1(n_1262), .B2(n_1263), .C(n_1264), .Y(n_1261) );
OAI31xp33_ASAP7_75t_L g751 ( .A1(n_752), .A2(n_754), .A3(n_762), .B(n_766), .Y(n_751) );
OAI22xp5_ASAP7_75t_L g1007 ( .A1(n_755), .A2(n_843), .B1(n_1008), .B2(n_1009), .Y(n_1007) );
OAI211xp5_ASAP7_75t_L g1154 ( .A1(n_755), .A2(n_1102), .B(n_1155), .C(n_1157), .Y(n_1154) );
HB1xp67_ASAP7_75t_L g1930 ( .A(n_755), .Y(n_1930) );
INVx2_ASAP7_75t_L g755 ( .A(n_756), .Y(n_755) );
INVx2_ASAP7_75t_L g805 ( .A(n_756), .Y(n_805) );
INVx1_ASAP7_75t_L g1577 ( .A(n_759), .Y(n_1577) );
INVx1_ASAP7_75t_L g1580 ( .A(n_763), .Y(n_1580) );
INVx2_ASAP7_75t_L g764 ( .A(n_765), .Y(n_764) );
AOI22xp33_ASAP7_75t_L g1579 ( .A1(n_765), .A2(n_1565), .B1(n_1566), .B2(n_1580), .Y(n_1579) );
OAI31xp33_ASAP7_75t_SL g1427 ( .A1(n_766), .A2(n_1428), .A3(n_1429), .B(n_1430), .Y(n_1427) );
OAI31xp33_ASAP7_75t_L g1444 ( .A1(n_766), .A2(n_1445), .A3(n_1446), .B(n_1450), .Y(n_1444) );
OAI31xp33_ASAP7_75t_SL g767 ( .A1(n_768), .A2(n_772), .A3(n_780), .B(n_782), .Y(n_767) );
INVx1_ASAP7_75t_L g769 ( .A(n_770), .Y(n_769) );
INVx1_ASAP7_75t_L g770 ( .A(n_771), .Y(n_770) );
OAI22xp5_ASAP7_75t_L g1900 ( .A1(n_773), .A2(n_824), .B1(n_1881), .B2(n_1894), .Y(n_1900) );
INVx2_ASAP7_75t_L g774 ( .A(n_775), .Y(n_774) );
INVx2_ASAP7_75t_L g1422 ( .A(n_775), .Y(n_1422) );
INVx1_ASAP7_75t_L g1358 ( .A(n_776), .Y(n_1358) );
INVx1_ASAP7_75t_L g776 ( .A(n_777), .Y(n_776) );
BUFx2_ASAP7_75t_L g1366 ( .A(n_777), .Y(n_1366) );
OAI21xp5_ASAP7_75t_L g1331 ( .A1(n_782), .A2(n_1332), .B(n_1344), .Y(n_1331) );
OAI31xp33_ASAP7_75t_L g1419 ( .A1(n_782), .A2(n_1420), .A3(n_1421), .B(n_1426), .Y(n_1419) );
BUFx3_ASAP7_75t_L g784 ( .A(n_785), .Y(n_784) );
INVx1_ASAP7_75t_L g785 ( .A(n_786), .Y(n_785) );
NAND3xp33_ASAP7_75t_SL g787 ( .A(n_788), .B(n_801), .C(n_811), .Y(n_787) );
OAI211xp5_ASAP7_75t_L g965 ( .A1(n_790), .A2(n_966), .B(n_967), .C(n_971), .Y(n_965) );
INVx1_ASAP7_75t_L g790 ( .A(n_791), .Y(n_790) );
INVx2_ASAP7_75t_L g827 ( .A(n_791), .Y(n_827) );
INVx1_ASAP7_75t_L g957 ( .A(n_791), .Y(n_957) );
INVx2_ASAP7_75t_L g978 ( .A(n_791), .Y(n_978) );
NAND3xp33_ASAP7_75t_L g1332 ( .A(n_792), .B(n_1333), .C(n_1338), .Y(n_1332) );
NAND4xp25_ASAP7_75t_L g1563 ( .A(n_792), .B(n_1564), .C(n_1567), .D(n_1570), .Y(n_1563) );
INVx2_ASAP7_75t_L g1336 ( .A(n_797), .Y(n_1336) );
INVx2_ASAP7_75t_L g797 ( .A(n_798), .Y(n_797) );
AOI22xp33_ASAP7_75t_L g1564 ( .A1(n_798), .A2(n_1334), .B1(n_1565), .B2(n_1566), .Y(n_1564) );
OAI31xp33_ASAP7_75t_SL g801 ( .A1(n_802), .A2(n_804), .A3(n_808), .B(n_810), .Y(n_801) );
OAI22xp33_ASAP7_75t_L g1540 ( .A1(n_805), .A2(n_837), .B1(n_1525), .B2(n_1531), .Y(n_1540) );
OAI31xp33_ASAP7_75t_SL g879 ( .A1(n_810), .A2(n_880), .A3(n_881), .B(n_885), .Y(n_879) );
OAI31xp33_ASAP7_75t_L g1058 ( .A1(n_810), .A2(n_1059), .A3(n_1063), .B(n_1066), .Y(n_1058) );
BUFx2_ASAP7_75t_L g1915 ( .A(n_810), .Y(n_1915) );
NOR2xp33_ASAP7_75t_SL g811 ( .A(n_812), .B(n_835), .Y(n_811) );
OAI22xp5_ASAP7_75t_L g813 ( .A1(n_814), .A2(n_815), .B1(n_816), .B2(n_817), .Y(n_813) );
OAI22xp5_ASAP7_75t_L g875 ( .A1(n_815), .A2(n_817), .B1(n_854), .B2(n_871), .Y(n_875) );
OAI22xp5_ASAP7_75t_L g1523 ( .A1(n_815), .A2(n_817), .B1(n_1524), .B2(n_1525), .Y(n_1523) );
OAI22xp5_ASAP7_75t_L g877 ( .A1(n_817), .A2(n_824), .B1(n_855), .B2(n_872), .Y(n_877) );
INVx1_ASAP7_75t_L g817 ( .A(n_818), .Y(n_817) );
INVx1_ASAP7_75t_L g818 ( .A(n_819), .Y(n_818) );
OAI22xp5_ASAP7_75t_L g823 ( .A1(n_824), .A2(n_826), .B1(n_827), .B2(n_828), .Y(n_823) );
INVx3_ASAP7_75t_L g824 ( .A(n_825), .Y(n_824) );
OAI211xp5_ASAP7_75t_SL g1649 ( .A1(n_827), .A2(n_1650), .B(n_1651), .C(n_1654), .Y(n_1649) );
HB1xp67_ASAP7_75t_L g1899 ( .A(n_827), .Y(n_1899) );
OAI33xp33_ASAP7_75t_L g1493 ( .A1(n_829), .A2(n_1456), .A3(n_1494), .B1(n_1499), .B2(n_1502), .B3(n_1505), .Y(n_1493) );
OAI33xp33_ASAP7_75t_L g1895 ( .A1(n_829), .A2(n_1456), .A3(n_1896), .B1(n_1898), .B2(n_1900), .B3(n_1901), .Y(n_1895) );
INVx2_ASAP7_75t_L g829 ( .A(n_830), .Y(n_829) );
INVx1_ASAP7_75t_L g830 ( .A(n_831), .Y(n_830) );
OR2x6_ASAP7_75t_L g910 ( .A(n_837), .B(n_911), .Y(n_910) );
INVx2_ASAP7_75t_SL g1032 ( .A(n_837), .Y(n_1032) );
OAI22xp5_ASAP7_75t_L g1038 ( .A1(n_840), .A2(n_1037), .B1(n_1039), .B2(n_1040), .Y(n_1038) );
INVx1_ASAP7_75t_L g1378 ( .A(n_840), .Y(n_1378) );
HB1xp67_ASAP7_75t_L g842 ( .A(n_843), .Y(n_842) );
HB1xp67_ASAP7_75t_L g870 ( .A(n_843), .Y(n_870) );
INVx1_ASAP7_75t_L g1511 ( .A(n_843), .Y(n_1511) );
OAI22xp5_ASAP7_75t_L g844 ( .A1(n_845), .A2(n_846), .B1(n_1557), .B2(n_1657), .Y(n_844) );
INVx1_ASAP7_75t_L g845 ( .A(n_846), .Y(n_845) );
XNOR2x1_ASAP7_75t_L g846 ( .A(n_847), .B(n_1383), .Y(n_846) );
XNOR2x1_ASAP7_75t_L g847 ( .A(n_848), .B(n_1070), .Y(n_847) );
XNOR2xp5_ASAP7_75t_L g848 ( .A(n_849), .B(n_895), .Y(n_848) );
NAND3xp33_ASAP7_75t_L g850 ( .A(n_851), .B(n_879), .C(n_886), .Y(n_850) );
NOR2xp33_ASAP7_75t_SL g851 ( .A(n_852), .B(n_873), .Y(n_851) );
OAI22xp5_ASAP7_75t_L g860 ( .A1(n_861), .A2(n_864), .B1(n_865), .B2(n_868), .Y(n_860) );
OAI22xp5_ASAP7_75t_L g1512 ( .A1(n_861), .A2(n_1037), .B1(n_1500), .B2(n_1506), .Y(n_1512) );
INVx1_ASAP7_75t_L g861 ( .A(n_862), .Y(n_861) );
INVx1_ASAP7_75t_L g862 ( .A(n_863), .Y(n_862) );
INVx3_ASAP7_75t_L g919 ( .A(n_863), .Y(n_919) );
BUFx2_ASAP7_75t_L g1372 ( .A(n_863), .Y(n_1372) );
OAI22xp5_ASAP7_75t_L g1029 ( .A1(n_865), .A2(n_1030), .B1(n_1031), .B2(n_1033), .Y(n_1029) );
INVx2_ASAP7_75t_SL g865 ( .A(n_866), .Y(n_865) );
INVx1_ASAP7_75t_L g866 ( .A(n_867), .Y(n_866) );
OAI22xp33_ASAP7_75t_L g1879 ( .A1(n_867), .A2(n_1510), .B1(n_1880), .B2(n_1881), .Y(n_1879) );
OAI33xp33_ASAP7_75t_L g1409 ( .A1(n_874), .A2(n_1410), .A3(n_1412), .B1(n_1414), .B2(n_1416), .B3(n_1418), .Y(n_1409) );
BUFx2_ASAP7_75t_L g890 ( .A(n_891), .Y(n_890) );
INVx2_ASAP7_75t_L g895 ( .A(n_896), .Y(n_895) );
AO22x2_ASAP7_75t_L g896 ( .A1(n_897), .A2(n_1014), .B1(n_1015), .B2(n_1069), .Y(n_896) );
INVx1_ASAP7_75t_SL g1069 ( .A(n_897), .Y(n_1069) );
XNOR2x1_ASAP7_75t_L g897 ( .A(n_898), .B(n_899), .Y(n_897) );
NOR2x1_ASAP7_75t_L g899 ( .A(n_900), .B(n_931), .Y(n_899) );
INVxp67_ASAP7_75t_L g901 ( .A(n_902), .Y(n_901) );
NAND2xp5_ASAP7_75t_L g902 ( .A(n_903), .B(n_910), .Y(n_902) );
INVx3_ASAP7_75t_L g903 ( .A(n_904), .Y(n_903) );
AOI22xp5_ASAP7_75t_L g1119 ( .A1(n_904), .A2(n_921), .B1(n_1120), .B2(n_1121), .Y(n_1119) );
AND2x4_ASAP7_75t_L g904 ( .A(n_905), .B(n_906), .Y(n_904) );
AND2x4_ASAP7_75t_L g921 ( .A(n_905), .B(n_922), .Y(n_921) );
BUFx6f_ASAP7_75t_L g1634 ( .A(n_906), .Y(n_1634) );
AND2x2_ASAP7_75t_L g906 ( .A(n_907), .B(n_908), .Y(n_906) );
AND2x2_ASAP7_75t_L g922 ( .A(n_907), .B(n_923), .Y(n_922) );
AND2x2_ASAP7_75t_L g985 ( .A(n_907), .B(n_986), .Y(n_985) );
BUFx2_ASAP7_75t_L g1205 ( .A(n_907), .Y(n_1205) );
AND2x4_ASAP7_75t_L g1631 ( .A(n_907), .B(n_1239), .Y(n_1631) );
AND2x4_ASAP7_75t_L g1637 ( .A(n_907), .B(n_923), .Y(n_1637) );
BUFx6f_ASAP7_75t_L g955 ( .A(n_908), .Y(n_955) );
INVx3_ASAP7_75t_L g973 ( .A(n_908), .Y(n_973) );
NAND2xp5_ASAP7_75t_L g1081 ( .A(n_908), .B(n_964), .Y(n_1081) );
INVxp67_ASAP7_75t_L g911 ( .A(n_912), .Y(n_911) );
AND2x2_ASAP7_75t_L g918 ( .A(n_912), .B(n_919), .Y(n_918) );
INVx1_ASAP7_75t_L g912 ( .A(n_913), .Y(n_912) );
OR2x2_ASAP7_75t_L g947 ( .A(n_913), .B(n_948), .Y(n_947) );
INVx1_ASAP7_75t_L g1169 ( .A(n_913), .Y(n_1169) );
INVx1_ASAP7_75t_L g1144 ( .A(n_914), .Y(n_1144) );
INVx1_ASAP7_75t_L g915 ( .A(n_916), .Y(n_915) );
NAND2x1_ASAP7_75t_L g916 ( .A(n_917), .B(n_920), .Y(n_916) );
INVx2_ASAP7_75t_SL g917 ( .A(n_918), .Y(n_917) );
INVx2_ASAP7_75t_L g1262 ( .A(n_919), .Y(n_1262) );
INVx2_ASAP7_75t_L g920 ( .A(n_921), .Y(n_920) );
BUFx6f_ASAP7_75t_L g980 ( .A(n_923), .Y(n_980) );
INVx2_ASAP7_75t_L g1208 ( .A(n_923), .Y(n_1208) );
INVx5_ASAP7_75t_L g1223 ( .A(n_924), .Y(n_1223) );
OR2x6_ASAP7_75t_L g924 ( .A(n_925), .B(n_930), .Y(n_924) );
OR2x2_ASAP7_75t_L g1627 ( .A(n_925), .B(n_930), .Y(n_1627) );
NAND2x1p5_ASAP7_75t_L g925 ( .A(n_926), .B(n_928), .Y(n_925) );
INVx8_ASAP7_75t_L g1131 ( .A(n_926), .Y(n_1131) );
HB1xp67_ASAP7_75t_L g1137 ( .A(n_926), .Y(n_1137) );
BUFx3_ASAP7_75t_L g1286 ( .A(n_926), .Y(n_1286) );
BUFx3_ASAP7_75t_L g1585 ( .A(n_926), .Y(n_1585) );
AND2x4_ASAP7_75t_L g937 ( .A(n_928), .B(n_938), .Y(n_937) );
AND2x6_ASAP7_75t_L g1125 ( .A(n_928), .B(n_935), .Y(n_1125) );
AND2x2_ASAP7_75t_L g1127 ( .A(n_928), .B(n_943), .Y(n_1127) );
INVx1_ASAP7_75t_L g1134 ( .A(n_928), .Y(n_1134) );
NAND3xp33_ASAP7_75t_SL g931 ( .A(n_932), .B(n_950), .C(n_996), .Y(n_931) );
AOI221xp5_ASAP7_75t_L g932 ( .A1(n_933), .A2(n_939), .B1(n_940), .B2(n_945), .C(n_946), .Y(n_932) );
INVx2_ASAP7_75t_L g933 ( .A(n_934), .Y(n_933) );
NAND2x1_ASAP7_75t_L g934 ( .A(n_935), .B(n_937), .Y(n_934) );
AND2x4_ASAP7_75t_SL g1190 ( .A(n_935), .B(n_937), .Y(n_1190) );
AND2x2_ASAP7_75t_L g1619 ( .A(n_935), .B(n_937), .Y(n_1619) );
INVx3_ASAP7_75t_L g935 ( .A(n_936), .Y(n_935) );
AND2x4_ASAP7_75t_L g940 ( .A(n_937), .B(n_941), .Y(n_940) );
AND2x4_ASAP7_75t_L g1012 ( .A(n_937), .B(n_1013), .Y(n_1012) );
AND2x4_ASAP7_75t_SL g1192 ( .A(n_937), .B(n_941), .Y(n_1192) );
OR2x2_ASAP7_75t_L g1080 ( .A(n_938), .B(n_1081), .Y(n_1080) );
AOI22xp33_ASAP7_75t_L g958 ( .A1(n_939), .A2(n_959), .B1(n_960), .B2(n_961), .Y(n_958) );
AOI22xp33_ASAP7_75t_L g1617 ( .A1(n_940), .A2(n_1618), .B1(n_1619), .B2(n_1620), .Y(n_1617) );
INVx2_ASAP7_75t_L g941 ( .A(n_942), .Y(n_941) );
INVx1_ASAP7_75t_L g942 ( .A(n_943), .Y(n_942) );
INVx1_ASAP7_75t_L g943 ( .A(n_944), .Y(n_943) );
INVx1_ASAP7_75t_L g1171 ( .A(n_947), .Y(n_1171) );
AND2x4_ASAP7_75t_L g1623 ( .A(n_947), .B(n_1080), .Y(n_1623) );
BUFx3_ASAP7_75t_L g1888 ( .A(n_948), .Y(n_1888) );
INVx2_ASAP7_75t_L g1165 ( .A(n_949), .Y(n_1165) );
AND2x4_ASAP7_75t_L g1626 ( .A(n_949), .B(n_1117), .Y(n_1626) );
OAI21xp5_ASAP7_75t_L g950 ( .A1(n_951), .A2(n_983), .B(n_992), .Y(n_950) );
NAND3xp33_ASAP7_75t_L g951 ( .A(n_952), .B(n_965), .C(n_976), .Y(n_951) );
A2O1A1Ixp33_ASAP7_75t_L g952 ( .A1(n_953), .A2(n_954), .B(n_956), .C(n_963), .Y(n_952) );
A2O1A1Ixp33_ASAP7_75t_SL g1246 ( .A1(n_954), .A2(n_963), .B(n_1247), .C(n_1248), .Y(n_1246) );
BUFx6f_ASAP7_75t_L g954 ( .A(n_955), .Y(n_954) );
INVx3_ASAP7_75t_L g1197 ( .A(n_955), .Y(n_1197) );
A2O1A1Ixp33_ASAP7_75t_L g1210 ( .A1(n_955), .A2(n_963), .B(n_1172), .C(n_1211), .Y(n_1210) );
A2O1A1Ixp33_ASAP7_75t_L g1317 ( .A1(n_955), .A2(n_1293), .B(n_1318), .C(n_1320), .Y(n_1317) );
NAND2xp5_ASAP7_75t_SL g956 ( .A(n_957), .B(n_958), .Y(n_956) );
OAI22xp5_ASAP7_75t_SL g1457 ( .A1(n_957), .A2(n_1411), .B1(n_1458), .B2(n_1459), .Y(n_1457) );
AOI22xp5_ASAP7_75t_L g1319 ( .A1(n_959), .A2(n_961), .B1(n_1291), .B2(n_1302), .Y(n_1319) );
INVx1_ASAP7_75t_L g1252 ( .A(n_961), .Y(n_1252) );
INVx1_ASAP7_75t_L g961 ( .A(n_962), .Y(n_961) );
HB1xp67_ASAP7_75t_L g963 ( .A(n_964), .Y(n_963) );
INVx1_ASAP7_75t_L g1321 ( .A(n_964), .Y(n_1321) );
BUFx2_ASAP7_75t_L g1353 ( .A(n_968), .Y(n_1353) );
HB1xp67_ASAP7_75t_L g1640 ( .A(n_968), .Y(n_1640) );
INVx2_ASAP7_75t_L g969 ( .A(n_970), .Y(n_969) );
OAI221xp5_ASAP7_75t_L g1199 ( .A1(n_970), .A2(n_978), .B1(n_1200), .B2(n_1201), .C(n_1202), .Y(n_1199) );
INVx1_ASAP7_75t_L g1243 ( .A(n_970), .Y(n_1243) );
INVx3_ASAP7_75t_L g1653 ( .A(n_970), .Y(n_1653) );
INVx1_ASAP7_75t_L g972 ( .A(n_973), .Y(n_972) );
INVx2_ASAP7_75t_L g1108 ( .A(n_973), .Y(n_1108) );
INVx1_ASAP7_75t_L g1356 ( .A(n_973), .Y(n_1356) );
BUFx3_ASAP7_75t_L g1354 ( .A(n_974), .Y(n_1354) );
INVx1_ASAP7_75t_SL g1596 ( .A(n_974), .Y(n_1596) );
BUFx3_ASAP7_75t_L g974 ( .A(n_975), .Y(n_974) );
INVx2_ASAP7_75t_L g987 ( .A(n_975), .Y(n_987) );
BUFx3_ASAP7_75t_L g1198 ( .A(n_975), .Y(n_1198) );
BUFx6f_ASAP7_75t_L g1239 ( .A(n_975), .Y(n_1239) );
OAI211xp5_ASAP7_75t_L g976 ( .A1(n_977), .A2(n_978), .B(n_979), .C(n_982), .Y(n_976) );
OAI22xp5_ASAP7_75t_L g1000 ( .A1(n_977), .A2(n_1001), .B1(n_1002), .B2(n_1003), .Y(n_1000) );
BUFx3_ASAP7_75t_L g1598 ( .A(n_980), .Y(n_1598) );
INVx2_ASAP7_75t_L g984 ( .A(n_985), .Y(n_984) );
AND2x4_ASAP7_75t_L g1083 ( .A(n_986), .B(n_1084), .Y(n_1083) );
INVx3_ASAP7_75t_L g986 ( .A(n_987), .Y(n_986) );
INVx1_ASAP7_75t_L g1245 ( .A(n_987), .Y(n_1245) );
INVx2_ASAP7_75t_L g988 ( .A(n_989), .Y(n_988) );
INVx2_ASAP7_75t_L g1646 ( .A(n_989), .Y(n_1646) );
INVx4_ASAP7_75t_L g989 ( .A(n_990), .Y(n_989) );
INVx2_ASAP7_75t_L g990 ( .A(n_991), .Y(n_990) );
HB1xp67_ASAP7_75t_L g992 ( .A(n_993), .Y(n_992) );
INVx1_ASAP7_75t_L g1656 ( .A(n_993), .Y(n_1656) );
BUFx2_ASAP7_75t_L g993 ( .A(n_994), .Y(n_993) );
OAI31xp33_ASAP7_75t_L g1194 ( .A1(n_994), .A2(n_1195), .A3(n_1203), .B(n_1213), .Y(n_1194) );
HB1xp67_ASAP7_75t_L g1230 ( .A(n_994), .Y(n_1230) );
OAI31xp33_ASAP7_75t_L g1306 ( .A1(n_994), .A2(n_1307), .A3(n_1313), .B(n_1322), .Y(n_1306) );
INVx1_ASAP7_75t_L g994 ( .A(n_995), .Y(n_994) );
AOI22xp33_ASAP7_75t_L g1138 ( .A1(n_998), .A2(n_1139), .B1(n_1140), .B2(n_1141), .Y(n_1138) );
BUFx3_ASAP7_75t_L g998 ( .A(n_999), .Y(n_998) );
BUFx3_ASAP7_75t_L g1180 ( .A(n_999), .Y(n_1180) );
BUFx12f_ASAP7_75t_L g1270 ( .A(n_999), .Y(n_1270) );
INVx5_ASAP7_75t_L g1297 ( .A(n_999), .Y(n_1297) );
OAI22xp33_ASAP7_75t_L g1393 ( .A1(n_1002), .A2(n_1394), .B1(n_1395), .B2(n_1396), .Y(n_1393) );
INVx1_ASAP7_75t_L g1005 ( .A(n_1006), .Y(n_1005) );
NAND3xp33_ASAP7_75t_L g1369 ( .A(n_1010), .B(n_1370), .C(n_1374), .Y(n_1369) );
AOI33xp33_ASAP7_75t_L g1582 ( .A1(n_1010), .A2(n_1583), .A3(n_1586), .B1(n_1587), .B2(n_1588), .B3(n_1589), .Y(n_1582) );
BUFx3_ASAP7_75t_L g1010 ( .A(n_1011), .Y(n_1010) );
AOI33xp33_ASAP7_75t_L g1173 ( .A1(n_1011), .A2(n_1174), .A3(n_1176), .B1(n_1177), .B2(n_1181), .B3(n_1184), .Y(n_1173) );
NAND3xp33_ASAP7_75t_L g1283 ( .A(n_1011), .B(n_1284), .C(n_1285), .Y(n_1283) );
AOI33xp33_ASAP7_75t_L g1609 ( .A1(n_1011), .A2(n_1184), .A3(n_1610), .B1(n_1613), .B2(n_1615), .B3(n_1616), .Y(n_1609) );
AOI221xp5_ASAP7_75t_L g1189 ( .A1(n_1012), .A2(n_1190), .B1(n_1191), .B2(n_1192), .C(n_1193), .Y(n_1189) );
AOI221xp5_ASAP7_75t_L g1301 ( .A1(n_1012), .A2(n_1190), .B1(n_1192), .B2(n_1302), .C(n_1303), .Y(n_1301) );
INVx3_ASAP7_75t_L g1605 ( .A(n_1012), .Y(n_1605) );
INVx1_ASAP7_75t_L g1014 ( .A(n_1015), .Y(n_1014) );
INVx1_ASAP7_75t_L g1016 ( .A(n_1017), .Y(n_1016) );
NAND3xp33_ASAP7_75t_L g1017 ( .A(n_1018), .B(n_1027), .C(n_1058), .Y(n_1017) );
NOR2xp33_ASAP7_75t_SL g1027 ( .A(n_1028), .B(n_1047), .Y(n_1027) );
OAI22xp5_ASAP7_75t_L g1048 ( .A1(n_1030), .A2(n_1045), .B1(n_1049), .B2(n_1052), .Y(n_1048) );
INVx1_ASAP7_75t_L g1031 ( .A(n_1032), .Y(n_1031) );
INVx1_ASAP7_75t_L g1517 ( .A(n_1032), .Y(n_1517) );
OAI22xp5_ASAP7_75t_L g1057 ( .A1(n_1036), .A2(n_1040), .B1(n_1049), .B2(n_1052), .Y(n_1057) );
OAI22xp5_ASAP7_75t_L g1882 ( .A1(n_1037), .A2(n_1883), .B1(n_1884), .B2(n_1885), .Y(n_1882) );
INVx1_ASAP7_75t_L g1041 ( .A(n_1042), .Y(n_1041) );
BUFx2_ASAP7_75t_L g1042 ( .A(n_1043), .Y(n_1042) );
BUFx2_ASAP7_75t_L g1588 ( .A(n_1043), .Y(n_1588) );
BUFx2_ASAP7_75t_L g1891 ( .A(n_1043), .Y(n_1891) );
INVx2_ASAP7_75t_L g1049 ( .A(n_1050), .Y(n_1049) );
INVx2_ASAP7_75t_SL g1050 ( .A(n_1051), .Y(n_1050) );
OAI22xp5_ASAP7_75t_L g1494 ( .A1(n_1052), .A2(n_1495), .B1(n_1496), .B2(n_1498), .Y(n_1494) );
OAI22xp5_ASAP7_75t_L g1505 ( .A1(n_1052), .A2(n_1496), .B1(n_1506), .B2(n_1507), .Y(n_1505) );
OAI22xp5_ASAP7_75t_L g1901 ( .A1(n_1052), .A2(n_1496), .B1(n_1885), .B2(n_1889), .Y(n_1901) );
INVx2_ASAP7_75t_L g1052 ( .A(n_1053), .Y(n_1052) );
INVx2_ASAP7_75t_L g1053 ( .A(n_1054), .Y(n_1053) );
OAI22xp5_ASAP7_75t_L g1217 ( .A1(n_1054), .A2(n_1218), .B1(n_1219), .B2(n_1220), .Y(n_1217) );
OAI22xp33_ASAP7_75t_L g1412 ( .A1(n_1054), .A2(n_1394), .B1(n_1406), .B2(n_1413), .Y(n_1412) );
OAI22xp33_ASAP7_75t_L g1453 ( .A1(n_1054), .A2(n_1413), .B1(n_1454), .B2(n_1455), .Y(n_1453) );
HB1xp67_ASAP7_75t_L g1897 ( .A(n_1054), .Y(n_1897) );
INVx2_ASAP7_75t_SL g1060 ( .A(n_1061), .Y(n_1060) );
XNOR2x1_ASAP7_75t_L g1070 ( .A(n_1071), .B(n_1328), .Y(n_1070) );
OA22x2_ASAP7_75t_L g1071 ( .A1(n_1072), .A2(n_1073), .B1(n_1225), .B2(n_1327), .Y(n_1071) );
INVx1_ASAP7_75t_L g1072 ( .A(n_1073), .Y(n_1072) );
XOR2xp5_ASAP7_75t_L g1073 ( .A(n_1074), .B(n_1161), .Y(n_1073) );
XNOR2x1_ASAP7_75t_L g1074 ( .A(n_1075), .B(n_1076), .Y(n_1074) );
NAND4xp75_ASAP7_75t_L g1076 ( .A(n_1077), .B(n_1087), .C(n_1119), .D(n_1122), .Y(n_1076) );
INVx1_ASAP7_75t_L g1078 ( .A(n_1079), .Y(n_1078) );
INVx1_ASAP7_75t_L g1079 ( .A(n_1080), .Y(n_1079) );
INVx1_ASAP7_75t_L g1082 ( .A(n_1083), .Y(n_1082) );
INVx1_ASAP7_75t_L g1084 ( .A(n_1085), .Y(n_1084) );
AOI211x1_ASAP7_75t_L g1087 ( .A1(n_1088), .A2(n_1099), .B(n_1100), .C(n_1113), .Y(n_1087) );
INVx2_ASAP7_75t_L g1089 ( .A(n_1090), .Y(n_1089) );
INVx2_ASAP7_75t_L g1090 ( .A(n_1091), .Y(n_1090) );
HB1xp67_ASAP7_75t_L g1362 ( .A(n_1091), .Y(n_1362) );
INVx2_ASAP7_75t_L g1091 ( .A(n_1092), .Y(n_1091) );
INVx2_ASAP7_75t_L g1652 ( .A(n_1092), .Y(n_1652) );
BUFx2_ASAP7_75t_L g1093 ( .A(n_1094), .Y(n_1093) );
AOI221xp5_ASAP7_75t_L g1206 ( .A1(n_1094), .A2(n_1186), .B1(n_1193), .B2(n_1207), .C(n_1209), .Y(n_1206) );
AOI221xp5_ASAP7_75t_L g1314 ( .A1(n_1094), .A2(n_1207), .B1(n_1289), .B2(n_1303), .C(n_1315), .Y(n_1314) );
INVx1_ASAP7_75t_L g1497 ( .A(n_1097), .Y(n_1497) );
OAI221xp5_ASAP7_75t_L g1101 ( .A1(n_1102), .A2(n_1103), .B1(n_1105), .B2(n_1106), .C(n_1107), .Y(n_1101) );
INVx2_ASAP7_75t_L g1103 ( .A(n_1104), .Y(n_1103) );
OAI211xp5_ASAP7_75t_SL g1235 ( .A1(n_1105), .A2(n_1236), .B(n_1237), .C(n_1238), .Y(n_1235) );
OAI211xp5_ASAP7_75t_SL g1240 ( .A1(n_1105), .A2(n_1241), .B(n_1242), .C(n_1244), .Y(n_1240) );
INVx1_ASAP7_75t_L g1110 ( .A(n_1111), .Y(n_1110) );
NAND2x2_ASAP7_75t_L g1114 ( .A(n_1111), .B(n_1115), .Y(n_1114) );
INVx2_ASAP7_75t_L g1111 ( .A(n_1112), .Y(n_1111) );
INVx2_ASAP7_75t_SL g1115 ( .A(n_1116), .Y(n_1115) );
OAI31xp67_ASAP7_75t_L g1122 ( .A1(n_1123), .A2(n_1135), .A3(n_1145), .B(n_1159), .Y(n_1122) );
INVx4_ASAP7_75t_L g1124 ( .A(n_1125), .Y(n_1124) );
INVx2_ASAP7_75t_L g1126 ( .A(n_1127), .Y(n_1126) );
A2O1A1Ixp33_ASAP7_75t_L g1128 ( .A1(n_1129), .A2(n_1130), .B(n_1132), .C(n_1133), .Y(n_1128) );
CKINVDCx5p33_ASAP7_75t_R g1130 ( .A(n_1131), .Y(n_1130) );
INVx3_ASAP7_75t_L g1158 ( .A(n_1131), .Y(n_1158) );
INVx2_ASAP7_75t_L g1168 ( .A(n_1131), .Y(n_1168) );
INVx8_ASAP7_75t_L g1175 ( .A(n_1131), .Y(n_1175) );
AOI22xp33_ASAP7_75t_L g1269 ( .A1(n_1132), .A2(n_1247), .B1(n_1270), .B2(n_1271), .Y(n_1269) );
INVx1_ASAP7_75t_L g1133 ( .A(n_1134), .Y(n_1133) );
AOI21xp33_ASAP7_75t_L g1135 ( .A1(n_1136), .A2(n_1138), .B(n_1142), .Y(n_1135) );
INVx1_ASAP7_75t_L g1142 ( .A(n_1143), .Y(n_1142) );
HB1xp67_ASAP7_75t_L g1143 ( .A(n_1144), .Y(n_1143) );
OAI21xp5_ASAP7_75t_SL g1145 ( .A1(n_1146), .A2(n_1149), .B(n_1154), .Y(n_1145) );
HB1xp67_ASAP7_75t_L g1447 ( .A(n_1147), .Y(n_1447) );
INVx2_ASAP7_75t_L g1150 ( .A(n_1151), .Y(n_1150) );
INVx2_ASAP7_75t_SL g1256 ( .A(n_1151), .Y(n_1256) );
BUFx2_ASAP7_75t_L g1159 ( .A(n_1160), .Y(n_1159) );
XNOR2x1_ASAP7_75t_L g1161 ( .A(n_1162), .B(n_1224), .Y(n_1161) );
OR2x2_ASAP7_75t_L g1162 ( .A(n_1163), .B(n_1188), .Y(n_1162) );
NAND3xp33_ASAP7_75t_L g1163 ( .A(n_1164), .B(n_1173), .C(n_1185), .Y(n_1163) );
AOI222xp33_ASAP7_75t_L g1164 ( .A1(n_1165), .A2(n_1166), .B1(n_1167), .B2(n_1170), .C1(n_1171), .C2(n_1172), .Y(n_1164) );
AOI222xp33_ASAP7_75t_L g1290 ( .A1(n_1165), .A2(n_1167), .B1(n_1171), .B2(n_1291), .C1(n_1292), .C2(n_1293), .Y(n_1290) );
AND2x4_ASAP7_75t_L g1167 ( .A(n_1168), .B(n_1169), .Y(n_1167) );
INVx2_ASAP7_75t_L g1178 ( .A(n_1179), .Y(n_1178) );
INVx1_ASAP7_75t_L g1182 ( .A(n_1183), .Y(n_1182) );
INVx2_ASAP7_75t_L g1260 ( .A(n_1183), .Y(n_1260) );
INVx1_ASAP7_75t_L g1287 ( .A(n_1183), .Y(n_1287) );
NAND3xp33_ASAP7_75t_L g1294 ( .A(n_1184), .B(n_1295), .C(n_1298), .Y(n_1294) );
NAND2xp5_ASAP7_75t_L g1185 ( .A(n_1186), .B(n_1187), .Y(n_1185) );
NAND2xp5_ASAP7_75t_L g1288 ( .A(n_1187), .B(n_1289), .Y(n_1288) );
INVx2_ASAP7_75t_L g1607 ( .A(n_1187), .Y(n_1607) );
NAND3xp33_ASAP7_75t_SL g1188 ( .A(n_1189), .B(n_1194), .C(n_1221), .Y(n_1188) );
INVx1_ASAP7_75t_L g1196 ( .A(n_1197), .Y(n_1196) );
OAI21xp33_ASAP7_75t_L g1203 ( .A1(n_1204), .A2(n_1206), .B(n_1210), .Y(n_1203) );
OAI21xp5_ASAP7_75t_SL g1313 ( .A1(n_1204), .A2(n_1314), .B(n_1317), .Y(n_1313) );
INVxp67_ASAP7_75t_L g1204 ( .A(n_1205), .Y(n_1204) );
OAI21xp5_ASAP7_75t_L g1232 ( .A1(n_1205), .A2(n_1233), .B(n_1234), .Y(n_1232) );
INVx2_ASAP7_75t_L g1207 ( .A(n_1208), .Y(n_1207) );
NAND2xp5_ASAP7_75t_L g1221 ( .A(n_1222), .B(n_1223), .Y(n_1221) );
NAND2xp5_ASAP7_75t_L g1304 ( .A(n_1223), .B(n_1305), .Y(n_1304) );
XNOR2xp5_ASAP7_75t_L g1225 ( .A(n_1226), .B(n_1280), .Y(n_1225) );
XOR2xp5_ASAP7_75t_L g1327 ( .A(n_1226), .B(n_1280), .Y(n_1327) );
XNOR2x1_ASAP7_75t_L g1226 ( .A(n_1227), .B(n_1228), .Y(n_1226) );
AND2x2_ASAP7_75t_L g1228 ( .A(n_1229), .B(n_1267), .Y(n_1228) );
AOI21xp5_ASAP7_75t_L g1229 ( .A1(n_1230), .A2(n_1231), .B(n_1254), .Y(n_1229) );
NAND4xp25_ASAP7_75t_L g1231 ( .A(n_1232), .B(n_1235), .C(n_1240), .D(n_1246), .Y(n_1231) );
INVx1_ASAP7_75t_L g1309 ( .A(n_1239), .Y(n_1309) );
BUFx2_ASAP7_75t_L g1368 ( .A(n_1239), .Y(n_1368) );
HB1xp67_ASAP7_75t_L g1643 ( .A(n_1239), .Y(n_1643) );
INVx1_ASAP7_75t_L g1249 ( .A(n_1250), .Y(n_1249) );
INVx1_ASAP7_75t_L g1250 ( .A(n_1251), .Y(n_1250) );
NOR2x1_ASAP7_75t_L g1648 ( .A(n_1251), .B(n_1321), .Y(n_1648) );
HB1xp67_ASAP7_75t_L g1373 ( .A(n_1265), .Y(n_1373) );
XNOR2x1_ASAP7_75t_L g1280 ( .A(n_1281), .B(n_1326), .Y(n_1280) );
OR2x2_ASAP7_75t_L g1281 ( .A(n_1282), .B(n_1300), .Y(n_1281) );
NAND4xp25_ASAP7_75t_SL g1282 ( .A(n_1283), .B(n_1288), .C(n_1290), .D(n_1294), .Y(n_1282) );
BUFx3_ASAP7_75t_L g1375 ( .A(n_1286), .Y(n_1375) );
INVx1_ASAP7_75t_L g1612 ( .A(n_1286), .Y(n_1612) );
INVx2_ASAP7_75t_L g1296 ( .A(n_1297), .Y(n_1296) );
INVx1_ASAP7_75t_L g1379 ( .A(n_1297), .Y(n_1379) );
INVx2_ASAP7_75t_R g1614 ( .A(n_1297), .Y(n_1614) );
NAND3xp33_ASAP7_75t_SL g1300 ( .A(n_1301), .B(n_1304), .C(n_1306), .Y(n_1300) );
INVx1_ASAP7_75t_L g1308 ( .A(n_1309), .Y(n_1308) );
INVx1_ASAP7_75t_L g1320 ( .A(n_1321), .Y(n_1320) );
INVx2_ASAP7_75t_L g1328 ( .A(n_1329), .Y(n_1328) );
INVx1_ASAP7_75t_L g1381 ( .A(n_1330), .Y(n_1381) );
NAND3xp33_ASAP7_75t_L g1330 ( .A(n_1331), .B(n_1345), .C(n_1350), .Y(n_1330) );
AOI22xp5_ASAP7_75t_L g1333 ( .A1(n_1334), .A2(n_1335), .B1(n_1336), .B2(n_1337), .Y(n_1333) );
INVx2_ASAP7_75t_L g1478 ( .A(n_1336), .Y(n_1478) );
AND4x1_ASAP7_75t_L g1350 ( .A(n_1351), .B(n_1360), .C(n_1369), .D(n_1376), .Y(n_1350) );
NAND3xp33_ASAP7_75t_L g1351 ( .A(n_1352), .B(n_1355), .C(n_1359), .Y(n_1351) );
INVx2_ASAP7_75t_L g1357 ( .A(n_1358), .Y(n_1357) );
INVx1_ASAP7_75t_L g1363 ( .A(n_1364), .Y(n_1363) );
INVx1_ASAP7_75t_L g1364 ( .A(n_1365), .Y(n_1364) );
INVx2_ASAP7_75t_L g1365 ( .A(n_1366), .Y(n_1365) );
INVx2_ASAP7_75t_L g1371 ( .A(n_1372), .Y(n_1371) );
OAI22xp5_ASAP7_75t_L g1397 ( .A1(n_1372), .A2(n_1398), .B1(n_1399), .B2(n_1400), .Y(n_1397) );
OAI22xp5_ASAP7_75t_L g1468 ( .A1(n_1372), .A2(n_1400), .B1(n_1458), .B2(n_1464), .Y(n_1468) );
OAI22xp5_ASAP7_75t_L g1886 ( .A1(n_1372), .A2(n_1887), .B1(n_1888), .B2(n_1889), .Y(n_1886) );
XNOR2xp5_ASAP7_75t_L g1383 ( .A(n_1384), .B(n_1472), .Y(n_1383) );
AOI22xp5_ASAP7_75t_L g1384 ( .A1(n_1385), .A2(n_1386), .B1(n_1434), .B2(n_1471), .Y(n_1384) );
INVx1_ASAP7_75t_L g1385 ( .A(n_1386), .Y(n_1385) );
HB1xp67_ASAP7_75t_L g1386 ( .A(n_1387), .Y(n_1386) );
XNOR2xp5_ASAP7_75t_L g1387 ( .A(n_1388), .B(n_1389), .Y(n_1387) );
AND3x1_ASAP7_75t_L g1389 ( .A(n_1390), .B(n_1419), .C(n_1427), .Y(n_1389) );
NOR2xp33_ASAP7_75t_SL g1390 ( .A(n_1391), .B(n_1409), .Y(n_1390) );
OAI33xp33_ASAP7_75t_L g1878 ( .A1(n_1392), .A2(n_1879), .A3(n_1882), .B1(n_1886), .B2(n_1890), .B3(n_1892), .Y(n_1878) );
OAI33xp33_ASAP7_75t_L g1452 ( .A1(n_1416), .A2(n_1453), .A3(n_1456), .B1(n_1457), .B2(n_1460), .B3(n_1463), .Y(n_1452) );
INVx2_ASAP7_75t_L g1416 ( .A(n_1417), .Y(n_1416) );
INVx1_ASAP7_75t_L g1471 ( .A(n_1434), .Y(n_1471) );
NAND3xp33_ASAP7_75t_L g1435 ( .A(n_1436), .B(n_1444), .C(n_1451), .Y(n_1435) );
NOR2xp33_ASAP7_75t_SL g1451 ( .A(n_1452), .B(n_1466), .Y(n_1451) );
OAI22xp5_ASAP7_75t_L g1472 ( .A1(n_1473), .A2(n_1518), .B1(n_1555), .B2(n_1556), .Y(n_1472) );
INVx1_ASAP7_75t_L g1555 ( .A(n_1473), .Y(n_1555) );
OAI221xp5_ASAP7_75t_L g1474 ( .A1(n_1475), .A2(n_1476), .B1(n_1484), .B2(n_1491), .C(n_1492), .Y(n_1474) );
NOR3xp33_ASAP7_75t_L g1476 ( .A(n_1477), .B(n_1479), .C(n_1480), .Y(n_1476) );
NOR3xp33_ASAP7_75t_L g1484 ( .A(n_1485), .B(n_1486), .C(n_1490), .Y(n_1484) );
NOR2xp33_ASAP7_75t_L g1492 ( .A(n_1493), .B(n_1508), .Y(n_1492) );
OAI22xp5_ASAP7_75t_SL g1896 ( .A1(n_1496), .A2(n_1880), .B1(n_1893), .B2(n_1897), .Y(n_1896) );
INVx2_ASAP7_75t_L g1496 ( .A(n_1497), .Y(n_1496) );
INVx2_ASAP7_75t_L g1510 ( .A(n_1511), .Y(n_1510) );
INVx1_ASAP7_75t_L g1514 ( .A(n_1515), .Y(n_1514) );
INVx1_ASAP7_75t_L g1556 ( .A(n_1518), .Y(n_1556) );
BUFx2_ASAP7_75t_L g1518 ( .A(n_1519), .Y(n_1518) );
NAND3xp33_ASAP7_75t_L g1520 ( .A(n_1521), .B(n_1541), .C(n_1548), .Y(n_1520) );
NOR2xp33_ASAP7_75t_L g1521 ( .A(n_1522), .B(n_1535), .Y(n_1521) );
INVx1_ASAP7_75t_L g1657 ( .A(n_1557), .Y(n_1657) );
INVx1_ASAP7_75t_L g1557 ( .A(n_1558), .Y(n_1557) );
INVx1_ASAP7_75t_L g1558 ( .A(n_1559), .Y(n_1558) );
XNOR2x1_ASAP7_75t_L g1559 ( .A(n_1560), .B(n_1601), .Y(n_1559) );
NAND3x1_ASAP7_75t_L g1561 ( .A(n_1562), .B(n_1582), .C(n_1590), .Y(n_1561) );
NAND3xp33_ASAP7_75t_L g1574 ( .A(n_1575), .B(n_1579), .C(n_1581), .Y(n_1574) );
BUFx2_ASAP7_75t_L g1584 ( .A(n_1585), .Y(n_1584) );
INVx1_ASAP7_75t_L g1591 ( .A(n_1592), .Y(n_1591) );
BUFx6f_ASAP7_75t_L g1592 ( .A(n_1593), .Y(n_1592) );
INVx1_ASAP7_75t_SL g1595 ( .A(n_1596), .Y(n_1595) );
AND3x1_ASAP7_75t_L g1602 ( .A(n_1603), .B(n_1621), .C(n_1628), .Y(n_1602) );
NOR3xp33_ASAP7_75t_L g1603 ( .A(n_1604), .B(n_1606), .C(n_1608), .Y(n_1603) );
INVx2_ASAP7_75t_SL g1604 ( .A(n_1605), .Y(n_1604) );
NAND2xp5_ASAP7_75t_SL g1608 ( .A(n_1609), .B(n_1617), .Y(n_1608) );
INVx1_ASAP7_75t_L g1611 ( .A(n_1612), .Y(n_1611) );
AOI21xp33_ASAP7_75t_L g1621 ( .A1(n_1622), .A2(n_1624), .B(n_1625), .Y(n_1621) );
INVx8_ASAP7_75t_L g1622 ( .A(n_1623), .Y(n_1622) );
OAI21xp5_ASAP7_75t_SL g1628 ( .A1(n_1629), .A2(n_1645), .B(n_1655), .Y(n_1628) );
INVx3_ASAP7_75t_L g1630 ( .A(n_1631), .Y(n_1630) );
AOI22xp33_ASAP7_75t_L g1632 ( .A1(n_1633), .A2(n_1634), .B1(n_1635), .B2(n_1636), .Y(n_1632) );
BUFx6f_ASAP7_75t_L g1636 ( .A(n_1637), .Y(n_1636) );
AOI21xp5_ASAP7_75t_L g1638 ( .A1(n_1639), .A2(n_1642), .B(n_1644), .Y(n_1638) );
INVx2_ASAP7_75t_L g1647 ( .A(n_1648), .Y(n_1647) );
INVx1_ASAP7_75t_L g1655 ( .A(n_1656), .Y(n_1655) );
OAI221xp5_ASAP7_75t_L g1658 ( .A1(n_1659), .A2(n_1872), .B1(n_1875), .B2(n_1916), .C(n_1919), .Y(n_1658) );
AOI21xp5_ASAP7_75t_L g1659 ( .A1(n_1660), .A2(n_1783), .B(n_1842), .Y(n_1659) );
NAND5xp2_ASAP7_75t_L g1660 ( .A(n_1661), .B(n_1726), .C(n_1746), .D(n_1759), .E(n_1769), .Y(n_1660) );
O2A1O1Ixp33_ASAP7_75t_L g1661 ( .A1(n_1662), .A2(n_1693), .B(n_1700), .C(n_1711), .Y(n_1661) );
INVx1_ASAP7_75t_L g1730 ( .A(n_1662), .Y(n_1730) );
AND2x2_ASAP7_75t_L g1662 ( .A(n_1663), .B(n_1683), .Y(n_1662) );
AND2x2_ASAP7_75t_L g1719 ( .A(n_1663), .B(n_1690), .Y(n_1719) );
AND2x2_ASAP7_75t_L g1758 ( .A(n_1663), .B(n_1685), .Y(n_1758) );
AND2x2_ASAP7_75t_L g1787 ( .A(n_1663), .B(n_1684), .Y(n_1787) );
NAND2xp5_ASAP7_75t_L g1795 ( .A(n_1663), .B(n_1796), .Y(n_1795) );
NAND2xp5_ASAP7_75t_L g1831 ( .A(n_1663), .B(n_1697), .Y(n_1831) );
INVx1_ASAP7_75t_L g1854 ( .A(n_1663), .Y(n_1854) );
AND2x2_ASAP7_75t_L g1663 ( .A(n_1664), .B(n_1679), .Y(n_1663) );
AND2x2_ASAP7_75t_L g1724 ( .A(n_1664), .B(n_1725), .Y(n_1724) );
NAND2xp5_ASAP7_75t_L g1737 ( .A(n_1664), .B(n_1684), .Y(n_1737) );
AND2x2_ASAP7_75t_L g1745 ( .A(n_1664), .B(n_1680), .Y(n_1745) );
AND3x1_ASAP7_75t_L g1819 ( .A(n_1664), .B(n_1680), .C(n_1684), .Y(n_1819) );
OR2x2_ASAP7_75t_L g1860 ( .A(n_1664), .B(n_1725), .Y(n_1860) );
INVx2_ASAP7_75t_L g1664 ( .A(n_1665), .Y(n_1664) );
AND2x2_ASAP7_75t_L g1699 ( .A(n_1665), .B(n_1679), .Y(n_1699) );
AND2x2_ASAP7_75t_L g1750 ( .A(n_1665), .B(n_1680), .Y(n_1750) );
OR2x2_ASAP7_75t_L g1665 ( .A(n_1666), .B(n_1673), .Y(n_1665) );
INVx2_ASAP7_75t_L g1780 ( .A(n_1667), .Y(n_1780) );
AND2x6_ASAP7_75t_L g1667 ( .A(n_1668), .B(n_1669), .Y(n_1667) );
AND2x2_ASAP7_75t_L g1671 ( .A(n_1668), .B(n_1672), .Y(n_1671) );
AND2x4_ASAP7_75t_L g1674 ( .A(n_1668), .B(n_1675), .Y(n_1674) );
AND2x6_ASAP7_75t_L g1677 ( .A(n_1668), .B(n_1678), .Y(n_1677) );
AND2x2_ASAP7_75t_L g1688 ( .A(n_1668), .B(n_1672), .Y(n_1688) );
AND2x2_ASAP7_75t_L g1709 ( .A(n_1668), .B(n_1672), .Y(n_1709) );
AND2x2_ASAP7_75t_L g1675 ( .A(n_1670), .B(n_1676), .Y(n_1675) );
INVxp67_ASAP7_75t_L g1782 ( .A(n_1671), .Y(n_1782) );
INVx2_ASAP7_75t_L g1874 ( .A(n_1677), .Y(n_1874) );
HB1xp67_ASAP7_75t_L g1966 ( .A(n_1678), .Y(n_1966) );
AND2x2_ASAP7_75t_L g1822 ( .A(n_1679), .B(n_1725), .Y(n_1822) );
INVx1_ASAP7_75t_L g1679 ( .A(n_1680), .Y(n_1679) );
OR2x2_ASAP7_75t_L g1755 ( .A(n_1680), .B(n_1725), .Y(n_1755) );
AND2x2_ASAP7_75t_L g1816 ( .A(n_1680), .B(n_1725), .Y(n_1816) );
AND2x2_ASAP7_75t_L g1680 ( .A(n_1681), .B(n_1682), .Y(n_1680) );
AND2x2_ASAP7_75t_L g1744 ( .A(n_1683), .B(n_1745), .Y(n_1744) );
NAND2xp5_ASAP7_75t_L g1830 ( .A(n_1683), .B(n_1750), .Y(n_1830) );
INVx1_ASAP7_75t_L g1857 ( .A(n_1683), .Y(n_1857) );
AND2x2_ASAP7_75t_L g1683 ( .A(n_1684), .B(n_1689), .Y(n_1683) );
AND2x2_ASAP7_75t_L g1765 ( .A(n_1684), .B(n_1699), .Y(n_1765) );
OR2x2_ASAP7_75t_L g1767 ( .A(n_1684), .B(n_1768), .Y(n_1767) );
INVx2_ASAP7_75t_L g1684 ( .A(n_1685), .Y(n_1684) );
AND2x2_ASAP7_75t_L g1698 ( .A(n_1685), .B(n_1699), .Y(n_1698) );
OAI322xp33_ASAP7_75t_L g1711 ( .A1(n_1685), .A2(n_1707), .A3(n_1712), .B1(n_1718), .B2(n_1720), .C1(n_1722), .C2(n_1723), .Y(n_1711) );
BUFx2_ASAP7_75t_L g1725 ( .A(n_1685), .Y(n_1725) );
OR2x2_ASAP7_75t_L g1748 ( .A(n_1685), .B(n_1749), .Y(n_1748) );
AOI321xp33_ASAP7_75t_L g1769 ( .A1(n_1685), .A2(n_1770), .A3(n_1771), .B1(n_1772), .B2(n_1774), .C(n_1776), .Y(n_1769) );
AND2x2_ASAP7_75t_L g1807 ( .A(n_1685), .B(n_1750), .Y(n_1807) );
OR2x2_ASAP7_75t_L g1868 ( .A(n_1685), .B(n_1802), .Y(n_1868) );
AND2x2_ASAP7_75t_L g1685 ( .A(n_1686), .B(n_1687), .Y(n_1685) );
NAND2xp5_ASAP7_75t_L g1764 ( .A(n_1689), .B(n_1701), .Y(n_1764) );
NAND2xp5_ASAP7_75t_L g1768 ( .A(n_1689), .B(n_1750), .Y(n_1768) );
NOR2xp33_ASAP7_75t_L g1774 ( .A(n_1689), .B(n_1775), .Y(n_1774) );
AND2x2_ASAP7_75t_L g1817 ( .A(n_1689), .B(n_1741), .Y(n_1817) );
NAND2xp5_ASAP7_75t_L g1841 ( .A(n_1689), .B(n_1699), .Y(n_1841) );
OAI21xp33_ASAP7_75t_L g1862 ( .A1(n_1689), .A2(n_1841), .B(n_1863), .Y(n_1862) );
INVx2_ASAP7_75t_L g1689 ( .A(n_1690), .Y(n_1689) );
INVx1_ASAP7_75t_L g1697 ( .A(n_1690), .Y(n_1697) );
AND2x2_ASAP7_75t_L g1736 ( .A(n_1690), .B(n_1703), .Y(n_1736) );
AND2x2_ASAP7_75t_L g1771 ( .A(n_1690), .B(n_1707), .Y(n_1771) );
AND2x2_ASAP7_75t_L g1794 ( .A(n_1690), .B(n_1725), .Y(n_1794) );
NAND2xp5_ASAP7_75t_L g1802 ( .A(n_1690), .B(n_1750), .Y(n_1802) );
NAND2xp5_ASAP7_75t_L g1850 ( .A(n_1690), .B(n_1715), .Y(n_1850) );
AND2x2_ASAP7_75t_L g1690 ( .A(n_1691), .B(n_1692), .Y(n_1690) );
INVx1_ASAP7_75t_L g1693 ( .A(n_1694), .Y(n_1693) );
NAND2xp5_ASAP7_75t_L g1694 ( .A(n_1695), .B(n_1698), .Y(n_1694) );
NAND2xp5_ASAP7_75t_L g1824 ( .A(n_1695), .B(n_1760), .Y(n_1824) );
INVx1_ASAP7_75t_L g1695 ( .A(n_1696), .Y(n_1695) );
NAND2xp5_ASAP7_75t_L g1712 ( .A(n_1696), .B(n_1713), .Y(n_1712) );
NOR2xp33_ASAP7_75t_L g1754 ( .A(n_1696), .B(n_1755), .Y(n_1754) );
NAND2xp5_ASAP7_75t_L g1786 ( .A(n_1696), .B(n_1787), .Y(n_1786) );
AND2x2_ASAP7_75t_L g1818 ( .A(n_1696), .B(n_1819), .Y(n_1818) );
AND2x2_ASAP7_75t_L g1826 ( .A(n_1696), .B(n_1765), .Y(n_1826) );
INVx2_ASAP7_75t_L g1696 ( .A(n_1697), .Y(n_1696) );
AND2x2_ASAP7_75t_L g1796 ( .A(n_1697), .B(n_1713), .Y(n_1796) );
O2A1O1Ixp33_ASAP7_75t_L g1870 ( .A1(n_1697), .A2(n_1839), .B(n_1840), .C(n_1871), .Y(n_1870) );
INVx1_ASAP7_75t_L g1871 ( .A(n_1698), .Y(n_1871) );
OR2x2_ASAP7_75t_L g1770 ( .A(n_1699), .B(n_1745), .Y(n_1770) );
INVx1_ASAP7_75t_L g1840 ( .A(n_1699), .Y(n_1840) );
AND2x2_ASAP7_75t_L g1700 ( .A(n_1701), .B(n_1706), .Y(n_1700) );
NAND2xp5_ASAP7_75t_L g1773 ( .A(n_1701), .B(n_1707), .Y(n_1773) );
INVx2_ASAP7_75t_L g1791 ( .A(n_1701), .Y(n_1791) );
A2O1A1O1Ixp25_ASAP7_75t_L g1836 ( .A1(n_1701), .A2(n_1715), .B(n_1793), .C(n_1837), .D(n_1838), .Y(n_1836) );
OR2x2_ASAP7_75t_L g1851 ( .A(n_1701), .B(n_1852), .Y(n_1851) );
INVx2_ASAP7_75t_L g1701 ( .A(n_1702), .Y(n_1701) );
AND2x2_ASAP7_75t_L g1721 ( .A(n_1702), .B(n_1706), .Y(n_1721) );
AND2x2_ASAP7_75t_L g1729 ( .A(n_1702), .B(n_1715), .Y(n_1729) );
INVx1_ASAP7_75t_L g1702 ( .A(n_1703), .Y(n_1702) );
OR2x2_ASAP7_75t_L g1714 ( .A(n_1703), .B(n_1715), .Y(n_1714) );
AND2x2_ASAP7_75t_L g1741 ( .A(n_1703), .B(n_1742), .Y(n_1741) );
AND2x2_ASAP7_75t_L g1829 ( .A(n_1703), .B(n_1715), .Y(n_1829) );
AND2x2_ASAP7_75t_L g1703 ( .A(n_1704), .B(n_1705), .Y(n_1703) );
NAND2xp5_ASAP7_75t_L g1722 ( .A(n_1706), .B(n_1713), .Y(n_1722) );
NOR2xp33_ASAP7_75t_L g1753 ( .A(n_1706), .B(n_1714), .Y(n_1753) );
AND2x2_ASAP7_75t_L g1788 ( .A(n_1706), .B(n_1741), .Y(n_1788) );
AND2x2_ASAP7_75t_L g1798 ( .A(n_1706), .B(n_1715), .Y(n_1798) );
OR2x2_ASAP7_75t_L g1809 ( .A(n_1706), .B(n_1715), .Y(n_1809) );
CKINVDCx6p67_ASAP7_75t_R g1706 ( .A(n_1707), .Y(n_1706) );
OR2x2_ASAP7_75t_L g1752 ( .A(n_1707), .B(n_1715), .Y(n_1752) );
AND2x2_ASAP7_75t_L g1760 ( .A(n_1707), .B(n_1715), .Y(n_1760) );
NAND2xp5_ASAP7_75t_L g1833 ( .A(n_1707), .B(n_1834), .Y(n_1833) );
CKINVDCx5p33_ASAP7_75t_R g1855 ( .A(n_1707), .Y(n_1855) );
OR2x2_ASAP7_75t_L g1858 ( .A(n_1707), .B(n_1728), .Y(n_1858) );
OR2x6_ASAP7_75t_L g1707 ( .A(n_1708), .B(n_1710), .Y(n_1707) );
OR2x2_ASAP7_75t_L g1811 ( .A(n_1708), .B(n_1710), .Y(n_1811) );
INVx1_ASAP7_75t_L g1844 ( .A(n_1712), .Y(n_1844) );
NAND2xp5_ASAP7_75t_L g1738 ( .A(n_1713), .B(n_1719), .Y(n_1738) );
INVx2_ASAP7_75t_L g1713 ( .A(n_1714), .Y(n_1713) );
INVx3_ASAP7_75t_L g1733 ( .A(n_1715), .Y(n_1733) );
INVx1_ASAP7_75t_L g1742 ( .A(n_1715), .Y(n_1742) );
AOI22xp5_ASAP7_75t_L g1759 ( .A1(n_1715), .A2(n_1760), .B1(n_1761), .B2(n_1766), .Y(n_1759) );
AND2x4_ASAP7_75t_L g1715 ( .A(n_1716), .B(n_1717), .Y(n_1715) );
INVxp67_ASAP7_75t_L g1718 ( .A(n_1719), .Y(n_1718) );
INVx1_ASAP7_75t_L g1720 ( .A(n_1721), .Y(n_1720) );
NAND2xp5_ASAP7_75t_L g1757 ( .A(n_1721), .B(n_1758), .Y(n_1757) );
INVx1_ASAP7_75t_L g1869 ( .A(n_1722), .Y(n_1869) );
CKINVDCx14_ASAP7_75t_R g1723 ( .A(n_1724), .Y(n_1723) );
AND2x2_ASAP7_75t_L g1799 ( .A(n_1725), .B(n_1745), .Y(n_1799) );
NOR2xp33_ASAP7_75t_L g1726 ( .A(n_1727), .B(n_1739), .Y(n_1726) );
OAI211xp5_ASAP7_75t_L g1727 ( .A1(n_1728), .A2(n_1730), .B(n_1731), .C(n_1738), .Y(n_1727) );
AOI21xp33_ASAP7_75t_L g1800 ( .A1(n_1728), .A2(n_1801), .B(n_1802), .Y(n_1800) );
CKINVDCx6p67_ASAP7_75t_R g1728 ( .A(n_1729), .Y(n_1728) );
AOI21xp33_ASAP7_75t_L g1864 ( .A1(n_1730), .A2(n_1805), .B(n_1865), .Y(n_1864) );
NAND2xp5_ASAP7_75t_L g1731 ( .A(n_1732), .B(n_1734), .Y(n_1731) );
CKINVDCx14_ASAP7_75t_R g1732 ( .A(n_1733), .Y(n_1732) );
AOI221xp5_ASAP7_75t_L g1866 ( .A1(n_1734), .A2(n_1760), .B1(n_1867), .B2(n_1869), .C(n_1870), .Y(n_1866) );
NOR2xp33_ASAP7_75t_L g1734 ( .A(n_1735), .B(n_1737), .Y(n_1734) );
CKINVDCx14_ASAP7_75t_R g1735 ( .A(n_1736), .Y(n_1735) );
INVx1_ASAP7_75t_L g1834 ( .A(n_1737), .Y(n_1834) );
NOR2xp33_ASAP7_75t_L g1739 ( .A(n_1740), .B(n_1743), .Y(n_1739) );
AOI21xp5_ASAP7_75t_L g1845 ( .A1(n_1740), .A2(n_1846), .B(n_1847), .Y(n_1845) );
INVx1_ASAP7_75t_L g1740 ( .A(n_1741), .Y(n_1740) );
INVx1_ASAP7_75t_L g1743 ( .A(n_1744), .Y(n_1743) );
INVx1_ASAP7_75t_L g1775 ( .A(n_1745), .Y(n_1775) );
AOI221xp5_ASAP7_75t_L g1746 ( .A1(n_1747), .A2(n_1751), .B1(n_1753), .B2(n_1754), .C(n_1756), .Y(n_1746) );
INVx1_ASAP7_75t_L g1747 ( .A(n_1748), .Y(n_1747) );
NAND2xp5_ASAP7_75t_L g1820 ( .A(n_1748), .B(n_1821), .Y(n_1820) );
INVx1_ASAP7_75t_L g1749 ( .A(n_1750), .Y(n_1749) );
AND2x2_ASAP7_75t_L g1793 ( .A(n_1750), .B(n_1794), .Y(n_1793) );
INVx1_ASAP7_75t_L g1751 ( .A(n_1752), .Y(n_1751) );
NAND2xp5_ASAP7_75t_L g1801 ( .A(n_1752), .B(n_1758), .Y(n_1801) );
OAI221xp5_ASAP7_75t_L g1838 ( .A1(n_1752), .A2(n_1776), .B1(n_1839), .B2(n_1840), .C(n_1841), .Y(n_1838) );
AOI221xp5_ASAP7_75t_L g1848 ( .A1(n_1753), .A2(n_1787), .B1(n_1849), .B2(n_1855), .C(n_1856), .Y(n_1848) );
INVx1_ASAP7_75t_L g1756 ( .A(n_1757), .Y(n_1756) );
AOI222xp33_ASAP7_75t_L g1812 ( .A1(n_1760), .A2(n_1813), .B1(n_1817), .B2(n_1818), .C1(n_1820), .C2(n_1823), .Y(n_1812) );
NAND2xp5_ASAP7_75t_L g1839 ( .A(n_1760), .B(n_1791), .Y(n_1839) );
INVx1_ASAP7_75t_L g1761 ( .A(n_1762), .Y(n_1761) );
NOR2xp33_ASAP7_75t_L g1810 ( .A(n_1762), .B(n_1811), .Y(n_1810) );
NAND2xp5_ASAP7_75t_L g1762 ( .A(n_1763), .B(n_1765), .Y(n_1762) );
OAI21xp33_ASAP7_75t_L g1797 ( .A1(n_1763), .A2(n_1798), .B(n_1799), .Y(n_1797) );
INVx1_ASAP7_75t_L g1763 ( .A(n_1764), .Y(n_1763) );
INVx1_ASAP7_75t_L g1814 ( .A(n_1765), .Y(n_1814) );
INVx1_ASAP7_75t_L g1766 ( .A(n_1767), .Y(n_1766) );
AOI211xp5_ASAP7_75t_SL g1856 ( .A1(n_1768), .A2(n_1857), .B(n_1858), .C(n_1859), .Y(n_1856) );
INVx1_ASAP7_75t_L g1772 ( .A(n_1773), .Y(n_1772) );
OAI22xp5_ASAP7_75t_L g1827 ( .A1(n_1773), .A2(n_1828), .B1(n_1830), .B2(n_1831), .Y(n_1827) );
INVx2_ASAP7_75t_SL g1776 ( .A(n_1777), .Y(n_1776) );
OAI22xp5_ASAP7_75t_SL g1778 ( .A1(n_1779), .A2(n_1780), .B1(n_1781), .B2(n_1782), .Y(n_1778) );
NAND5xp2_ASAP7_75t_L g1783 ( .A(n_1784), .B(n_1803), .C(n_1812), .D(n_1825), .E(n_1836), .Y(n_1783) );
AOI211xp5_ASAP7_75t_L g1784 ( .A1(n_1785), .A2(n_1788), .B(n_1789), .C(n_1800), .Y(n_1784) );
INVx1_ASAP7_75t_L g1785 ( .A(n_1786), .Y(n_1785) );
AOI221xp5_ASAP7_75t_L g1861 ( .A1(n_1788), .A2(n_1818), .B1(n_1829), .B2(n_1862), .C(n_1864), .Y(n_1861) );
OAI211xp5_ASAP7_75t_L g1789 ( .A1(n_1790), .A2(n_1792), .B(n_1795), .C(n_1797), .Y(n_1789) );
NAND2xp5_ASAP7_75t_L g1805 ( .A(n_1790), .B(n_1806), .Y(n_1805) );
INVx2_ASAP7_75t_L g1790 ( .A(n_1791), .Y(n_1790) );
INVx1_ASAP7_75t_L g1792 ( .A(n_1793), .Y(n_1792) );
INVx1_ASAP7_75t_L g1853 ( .A(n_1794), .Y(n_1853) );
INVx1_ASAP7_75t_L g1835 ( .A(n_1796), .Y(n_1835) );
INVx1_ASAP7_75t_L g1865 ( .A(n_1798), .Y(n_1865) );
INVx1_ASAP7_75t_L g1863 ( .A(n_1799), .Y(n_1863) );
INVxp67_ASAP7_75t_SL g1837 ( .A(n_1801), .Y(n_1837) );
INVx1_ASAP7_75t_L g1806 ( .A(n_1802), .Y(n_1806) );
O2A1O1Ixp33_ASAP7_75t_SL g1803 ( .A1(n_1804), .A2(n_1807), .B(n_1808), .C(n_1810), .Y(n_1803) );
INVxp67_ASAP7_75t_SL g1804 ( .A(n_1805), .Y(n_1804) );
INVx1_ASAP7_75t_L g1847 ( .A(n_1807), .Y(n_1847) );
INVx1_ASAP7_75t_L g1808 ( .A(n_1809), .Y(n_1808) );
AOI211xp5_ASAP7_75t_L g1825 ( .A1(n_1811), .A2(n_1826), .B(n_1827), .C(n_1832), .Y(n_1825) );
A2O1A1Ixp33_ASAP7_75t_L g1843 ( .A1(n_1811), .A2(n_1816), .B(n_1844), .C(n_1845), .Y(n_1843) );
NAND2xp5_ASAP7_75t_SL g1813 ( .A(n_1814), .B(n_1815), .Y(n_1813) );
INVx1_ASAP7_75t_L g1815 ( .A(n_1816), .Y(n_1815) );
AOI21xp33_ASAP7_75t_L g1832 ( .A1(n_1821), .A2(n_1833), .B(n_1835), .Y(n_1832) );
OAI21xp33_ASAP7_75t_L g1849 ( .A1(n_1821), .A2(n_1850), .B(n_1851), .Y(n_1849) );
INVx1_ASAP7_75t_L g1821 ( .A(n_1822), .Y(n_1821) );
INVxp67_ASAP7_75t_SL g1823 ( .A(n_1824), .Y(n_1823) );
INVx1_ASAP7_75t_L g1846 ( .A(n_1826), .Y(n_1846) );
INVx2_ASAP7_75t_L g1828 ( .A(n_1829), .Y(n_1828) );
NAND4xp25_ASAP7_75t_L g1842 ( .A(n_1843), .B(n_1848), .C(n_1861), .D(n_1866), .Y(n_1842) );
OR2x2_ASAP7_75t_L g1852 ( .A(n_1853), .B(n_1854), .Y(n_1852) );
INVx1_ASAP7_75t_L g1859 ( .A(n_1860), .Y(n_1859) );
INVx1_ASAP7_75t_L g1867 ( .A(n_1868), .Y(n_1867) );
CKINVDCx20_ASAP7_75t_R g1872 ( .A(n_1873), .Y(n_1872) );
CKINVDCx20_ASAP7_75t_R g1873 ( .A(n_1874), .Y(n_1873) );
NAND3xp33_ASAP7_75t_L g1876 ( .A(n_1877), .B(n_1902), .C(n_1909), .Y(n_1876) );
NOR2xp33_ASAP7_75t_L g1877 ( .A(n_1878), .B(n_1895), .Y(n_1877) );
INVx1_ASAP7_75t_L g1890 ( .A(n_1891), .Y(n_1890) );
OAI31xp33_ASAP7_75t_L g1909 ( .A1(n_1910), .A2(n_1911), .A3(n_1914), .B(n_1915), .Y(n_1909) );
INVx3_ASAP7_75t_L g1916 ( .A(n_1917), .Y(n_1916) );
HB1xp67_ASAP7_75t_L g1920 ( .A(n_1921), .Y(n_1920) );
BUFx3_ASAP7_75t_L g1921 ( .A(n_1922), .Y(n_1921) );
INVxp33_ASAP7_75t_L g1923 ( .A(n_1924), .Y(n_1923) );
HB1xp67_ASAP7_75t_L g1925 ( .A(n_1926), .Y(n_1925) );
NAND3xp33_ASAP7_75t_L g1926 ( .A(n_1927), .B(n_1937), .C(n_1944), .Y(n_1926) );
INVx1_ASAP7_75t_L g1935 ( .A(n_1936), .Y(n_1935) );
NOR2xp33_ASAP7_75t_L g1944 ( .A(n_1945), .B(n_1958), .Y(n_1944) );
HB1xp67_ASAP7_75t_L g1964 ( .A(n_1965), .Y(n_1964) );
OAI21xp5_ASAP7_75t_L g1965 ( .A1(n_1966), .A2(n_1967), .B(n_1968), .Y(n_1965) );
INVx1_ASAP7_75t_L g1968 ( .A(n_1969), .Y(n_1968) );
endmodule