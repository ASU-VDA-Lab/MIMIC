module fake_jpeg_11056_n_648 (n_13, n_1, n_10, n_6, n_14, n_18, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_648);

input n_13;
input n_1;
input n_10;
input n_6;
input n_14;
input n_18;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_648;

wire n_529;
wire n_595;
wire n_390;
wire n_552;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_252;
wire n_19;
wire n_182;
wire n_525;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_586;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_620;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_611;
wire n_44;
wire n_355;
wire n_519;
wire n_276;
wire n_143;
wire n_431;
wire n_102;
wire n_549;
wire n_196;
wire n_66;
wire n_374;
wire n_566;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_597;
wire n_172;
wire n_547;
wire n_345;
wire n_591;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_513;
wire n_283;
wire n_107;
wire n_490;
wire n_635;
wire n_517;
wire n_629;
wire n_415;
wire n_479;
wire n_543;
wire n_357;
wire n_89;
wire n_131;
wire n_607;
wire n_294;
wire n_230;
wire n_643;
wire n_170;
wire n_602;
wire n_313;
wire n_542;
wire n_574;
wire n_264;
wire n_647;
wire n_437;
wire n_93;
wire n_227;
wire n_559;
wire n_641;
wire n_48;
wire n_465;
wire n_638;
wire n_200;
wire n_582;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_623;
wire n_579;
wire n_416;
wire n_221;
wire n_256;
wire n_454;
wire n_540;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_637;
wire n_370;
wire n_410;
wire n_571;
wire n_82;
wire n_155;
wire n_508;
wire n_309;
wire n_624;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_606;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_569;
wire n_596;
wire n_400;
wire n_646;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_544;
wire n_31;
wire n_277;
wire n_255;
wire n_605;
wire n_601;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_530;
wire n_634;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_557;
wire n_408;
wire n_80;
wire n_562;
wire n_204;
wire n_639;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_645;
wire n_298;
wire n_106;
wire n_545;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_584;
wire n_254;
wire n_608;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_622;
wire n_463;
wire n_92;
wire n_332;
wire n_640;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_474;
wire n_539;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_626;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_575;
wire n_268;
wire n_404;
wire n_91;
wire n_511;
wire n_486;
wire n_305;
wire n_161;
wire n_441;
wire n_555;
wire n_342;
wire n_642;
wire n_101;
wire n_226;
wire n_509;
wire n_644;
wire n_149;
wire n_87;
wire n_46;
wire n_578;
wire n_589;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_614;
wire n_97;
wire n_573;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_610;
wire n_174;
wire n_198;
wire n_422;
wire n_560;
wire n_190;
wire n_510;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_536;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_537;
wire n_110;
wire n_594;
wire n_590;
wire n_531;
wire n_76;
wire n_278;
wire n_343;
wire n_577;
wire n_26;
wire n_88;
wire n_397;
wire n_592;
wire n_363;
wire n_570;
wire n_238;
wire n_598;
wire n_615;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_554;
wire n_301;
wire n_609;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_523;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_533;
wire n_612;
wire n_384;
wire n_296;
wire n_588;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_585;
wire n_491;
wire n_24;
wire n_526;
wire n_467;
wire n_269;
wire n_572;
wire n_546;
wire n_287;
wire n_219;
wire n_452;
wire n_631;
wire n_433;
wire n_636;
wire n_77;
wire n_473;
wire n_45;
wire n_520;
wire n_476;
wire n_337;
wire n_317;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_344;
wire n_328;
wire n_218;
wire n_63;
wire n_599;
wire n_239;
wire n_243;
wire n_481;
wire n_628;
wire n_619;
wire n_348;
wire n_587;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_583;
wire n_522;
wire n_333;
wire n_518;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_565;
wire n_302;
wire n_216;
wire n_528;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_199;
wire n_260;
wire n_550;
wire n_413;
wire n_275;
wire n_494;
wire n_604;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_551;
wire n_36;
wire n_62;
wire n_600;
wire n_492;
wire n_603;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_567;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_515;
wire n_347;
wire n_521;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_538;
wire n_625;
wire n_147;
wire n_449;
wire n_627;
wire n_98;
wire n_251;
wire n_534;
wire n_472;
wire n_279;
wire n_593;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_618;
wire n_356;
wire n_119;
wire n_484;
wire n_568;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_576;
wire n_469;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_553;
wire n_257;
wire n_61;
wire n_173;
wire n_561;
wire n_244;
wire n_232;
wire n_527;
wire n_482;
wire n_58;
wire n_41;
wire n_613;
wire n_630;
wire n_266;
wire n_548;
wire n_72;
wire n_512;
wire n_445;
wire n_443;
wire n_617;
wire n_215;
wire n_212;
wire n_516;
wire n_183;
wire n_409;
wire n_532;
wire n_249;
wire n_412;
wire n_581;
wire n_217;
wire n_471;
wire n_580;
wire n_541;
wire n_53;
wire n_372;
wire n_558;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_535;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_556;
wire n_524;
wire n_402;
wire n_563;
wire n_504;
wire n_438;
wire n_475;
wire n_247;
wire n_157;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_633;
wire n_112;
wire n_632;
wire n_616;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_514;
wire n_564;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_621;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_6),
.Y(n_19)
);

INVx8_ASAP7_75t_L g20 ( 
.A(n_18),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_0),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_11),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_17),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_0),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_11),
.Y(n_25)
);

NOR2xp33_ASAP7_75t_L g26 ( 
.A(n_3),
.B(n_18),
.Y(n_26)
);

INVx11_ASAP7_75t_L g27 ( 
.A(n_5),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_5),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_8),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_18),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_15),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_16),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_18),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_17),
.Y(n_34)
);

BUFx12f_ASAP7_75t_L g35 ( 
.A(n_0),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_0),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_15),
.Y(n_37)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_4),
.Y(n_38)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_5),
.Y(n_39)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_9),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_15),
.Y(n_41)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_4),
.Y(n_42)
);

BUFx12f_ASAP7_75t_L g43 ( 
.A(n_14),
.Y(n_43)
);

BUFx12_ASAP7_75t_L g44 ( 
.A(n_12),
.Y(n_44)
);

BUFx12f_ASAP7_75t_L g45 ( 
.A(n_17),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_10),
.Y(n_46)
);

BUFx4f_ASAP7_75t_L g47 ( 
.A(n_13),
.Y(n_47)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_11),
.Y(n_48)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_14),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_2),
.Y(n_50)
);

OR2x2_ASAP7_75t_L g51 ( 
.A(n_6),
.B(n_5),
.Y(n_51)
);

BUFx2_ASAP7_75t_L g52 ( 
.A(n_6),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_6),
.Y(n_53)
);

INVxp67_ASAP7_75t_L g54 ( 
.A(n_8),
.Y(n_54)
);

BUFx16f_ASAP7_75t_L g55 ( 
.A(n_13),
.Y(n_55)
);

BUFx5_ASAP7_75t_L g56 ( 
.A(n_7),
.Y(n_56)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_1),
.Y(n_57)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_14),
.Y(n_58)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_9),
.Y(n_59)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_13),
.Y(n_60)
);

BUFx5_ASAP7_75t_L g61 ( 
.A(n_17),
.Y(n_61)
);

CKINVDCx20_ASAP7_75t_R g62 ( 
.A(n_9),
.Y(n_62)
);

BUFx3_ASAP7_75t_L g63 ( 
.A(n_56),
.Y(n_63)
);

INVx5_ASAP7_75t_L g150 ( 
.A(n_63),
.Y(n_150)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_38),
.Y(n_64)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_64),
.Y(n_133)
);

INVx3_ASAP7_75t_L g65 ( 
.A(n_55),
.Y(n_65)
);

INVx3_ASAP7_75t_L g134 ( 
.A(n_65),
.Y(n_134)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_47),
.Y(n_66)
);

INVx2_ASAP7_75t_L g131 ( 
.A(n_66),
.Y(n_131)
);

INVx3_ASAP7_75t_L g67 ( 
.A(n_55),
.Y(n_67)
);

INVx3_ASAP7_75t_L g151 ( 
.A(n_67),
.Y(n_151)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_19),
.Y(n_68)
);

BUFx6f_ASAP7_75t_L g132 ( 
.A(n_68),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_SL g69 ( 
.A(n_26),
.B(n_1),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_L g164 ( 
.A(n_69),
.B(n_71),
.Y(n_164)
);

BUFx6f_ASAP7_75t_L g70 ( 
.A(n_19),
.Y(n_70)
);

BUFx6f_ASAP7_75t_L g138 ( 
.A(n_70),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_SL g71 ( 
.A(n_26),
.B(n_1),
.Y(n_71)
);

BUFx6f_ASAP7_75t_L g72 ( 
.A(n_19),
.Y(n_72)
);

BUFx6f_ASAP7_75t_L g158 ( 
.A(n_72),
.Y(n_158)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_38),
.Y(n_73)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_73),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_51),
.B(n_54),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_SL g170 ( 
.A(n_74),
.B(n_107),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_L g75 ( 
.A(n_51),
.B(n_1),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_L g177 ( 
.A(n_75),
.B(n_116),
.Y(n_177)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_39),
.Y(n_76)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_76),
.Y(n_153)
);

INVx2_ASAP7_75t_L g77 ( 
.A(n_47),
.Y(n_77)
);

INVx2_ASAP7_75t_L g136 ( 
.A(n_77),
.Y(n_136)
);

INVx11_ASAP7_75t_L g78 ( 
.A(n_27),
.Y(n_78)
);

INVx11_ASAP7_75t_L g145 ( 
.A(n_78),
.Y(n_145)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_39),
.Y(n_79)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_79),
.Y(n_155)
);

BUFx12f_ASAP7_75t_L g80 ( 
.A(n_56),
.Y(n_80)
);

INVx5_ASAP7_75t_L g187 ( 
.A(n_80),
.Y(n_187)
);

INVx3_ASAP7_75t_L g81 ( 
.A(n_55),
.Y(n_81)
);

INVx3_ASAP7_75t_L g174 ( 
.A(n_81),
.Y(n_174)
);

INVx11_ASAP7_75t_L g82 ( 
.A(n_27),
.Y(n_82)
);

BUFx2_ASAP7_75t_L g208 ( 
.A(n_82),
.Y(n_208)
);

INVx2_ASAP7_75t_SL g83 ( 
.A(n_56),
.Y(n_83)
);

INVx13_ASAP7_75t_L g165 ( 
.A(n_83),
.Y(n_165)
);

OR2x2_ASAP7_75t_L g84 ( 
.A(n_40),
.B(n_42),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g139 ( 
.A(n_84),
.B(n_99),
.Y(n_139)
);

INVx6_ASAP7_75t_L g85 ( 
.A(n_19),
.Y(n_85)
);

BUFx6f_ASAP7_75t_L g160 ( 
.A(n_85),
.Y(n_160)
);

INVx4_ASAP7_75t_L g86 ( 
.A(n_35),
.Y(n_86)
);

INVx3_ASAP7_75t_L g179 ( 
.A(n_86),
.Y(n_179)
);

BUFx3_ASAP7_75t_L g87 ( 
.A(n_61),
.Y(n_87)
);

INVx4_ASAP7_75t_L g135 ( 
.A(n_87),
.Y(n_135)
);

BUFx6f_ASAP7_75t_L g88 ( 
.A(n_32),
.Y(n_88)
);

BUFx6f_ASAP7_75t_L g161 ( 
.A(n_88),
.Y(n_161)
);

INVx3_ASAP7_75t_L g89 ( 
.A(n_55),
.Y(n_89)
);

INVx3_ASAP7_75t_L g188 ( 
.A(n_89),
.Y(n_188)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_40),
.Y(n_90)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_90),
.Y(n_159)
);

INVx2_ASAP7_75t_L g91 ( 
.A(n_47),
.Y(n_91)
);

INVx2_ASAP7_75t_L g143 ( 
.A(n_91),
.Y(n_143)
);

BUFx3_ASAP7_75t_L g92 ( 
.A(n_61),
.Y(n_92)
);

INVx4_ASAP7_75t_L g144 ( 
.A(n_92),
.Y(n_144)
);

INVx4_ASAP7_75t_SL g93 ( 
.A(n_27),
.Y(n_93)
);

INVx2_ASAP7_75t_SL g210 ( 
.A(n_93),
.Y(n_210)
);

BUFx6f_ASAP7_75t_L g94 ( 
.A(n_32),
.Y(n_94)
);

BUFx6f_ASAP7_75t_L g168 ( 
.A(n_94),
.Y(n_168)
);

BUFx3_ASAP7_75t_L g95 ( 
.A(n_61),
.Y(n_95)
);

INVx4_ASAP7_75t_L g148 ( 
.A(n_95),
.Y(n_148)
);

INVx3_ASAP7_75t_L g96 ( 
.A(n_55),
.Y(n_96)
);

INVx3_ASAP7_75t_L g190 ( 
.A(n_96),
.Y(n_190)
);

BUFx6f_ASAP7_75t_L g97 ( 
.A(n_32),
.Y(n_97)
);

INVx6_ASAP7_75t_L g178 ( 
.A(n_97),
.Y(n_178)
);

BUFx6f_ASAP7_75t_L g98 ( 
.A(n_32),
.Y(n_98)
);

INVx6_ASAP7_75t_L g181 ( 
.A(n_98),
.Y(n_181)
);

CKINVDCx16_ASAP7_75t_R g99 ( 
.A(n_44),
.Y(n_99)
);

BUFx6f_ASAP7_75t_L g100 ( 
.A(n_50),
.Y(n_100)
);

INVx6_ASAP7_75t_L g202 ( 
.A(n_100),
.Y(n_202)
);

INVx3_ASAP7_75t_SL g101 ( 
.A(n_20),
.Y(n_101)
);

INVx2_ASAP7_75t_L g146 ( 
.A(n_101),
.Y(n_146)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_42),
.Y(n_102)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_102),
.Y(n_172)
);

INVx11_ASAP7_75t_L g103 ( 
.A(n_44),
.Y(n_103)
);

INVx4_ASAP7_75t_L g156 ( 
.A(n_103),
.Y(n_156)
);

BUFx6f_ASAP7_75t_L g104 ( 
.A(n_50),
.Y(n_104)
);

INVx3_ASAP7_75t_SL g176 ( 
.A(n_104),
.Y(n_176)
);

INVx3_ASAP7_75t_L g105 ( 
.A(n_35),
.Y(n_105)
);

INVx3_ASAP7_75t_L g191 ( 
.A(n_105),
.Y(n_191)
);

BUFx3_ASAP7_75t_L g106 ( 
.A(n_35),
.Y(n_106)
);

INVx4_ASAP7_75t_L g171 ( 
.A(n_106),
.Y(n_171)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_51),
.B(n_2),
.Y(n_107)
);

BUFx24_ASAP7_75t_L g108 ( 
.A(n_44),
.Y(n_108)
);

INVx4_ASAP7_75t_L g197 ( 
.A(n_108),
.Y(n_197)
);

BUFx6f_ASAP7_75t_L g109 ( 
.A(n_50),
.Y(n_109)
);

INVx4_ASAP7_75t_L g198 ( 
.A(n_109),
.Y(n_198)
);

INVx3_ASAP7_75t_L g110 ( 
.A(n_35),
.Y(n_110)
);

INVx3_ASAP7_75t_L g205 ( 
.A(n_110),
.Y(n_205)
);

BUFx6f_ASAP7_75t_L g111 ( 
.A(n_50),
.Y(n_111)
);

INVx2_ASAP7_75t_L g154 ( 
.A(n_111),
.Y(n_154)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_49),
.Y(n_112)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_112),
.Y(n_173)
);

INVx3_ASAP7_75t_L g113 ( 
.A(n_35),
.Y(n_113)
);

INVx2_ASAP7_75t_L g157 ( 
.A(n_113),
.Y(n_157)
);

INVx2_ASAP7_75t_L g114 ( 
.A(n_47),
.Y(n_114)
);

INVx2_ASAP7_75t_L g169 ( 
.A(n_114),
.Y(n_169)
);

BUFx12_ASAP7_75t_L g115 ( 
.A(n_44),
.Y(n_115)
);

CKINVDCx20_ASAP7_75t_R g182 ( 
.A(n_115),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_L g116 ( 
.A(n_51),
.B(n_16),
.Y(n_116)
);

BUFx6f_ASAP7_75t_L g117 ( 
.A(n_53),
.Y(n_117)
);

INVx2_ASAP7_75t_L g183 ( 
.A(n_117),
.Y(n_183)
);

INVx3_ASAP7_75t_L g118 ( 
.A(n_43),
.Y(n_118)
);

INVx2_ASAP7_75t_L g185 ( 
.A(n_118),
.Y(n_185)
);

BUFx6f_ASAP7_75t_L g119 ( 
.A(n_53),
.Y(n_119)
);

INVx2_ASAP7_75t_L g186 ( 
.A(n_119),
.Y(n_186)
);

INVx13_ASAP7_75t_L g120 ( 
.A(n_44),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_L g152 ( 
.A(n_120),
.B(n_121),
.Y(n_152)
);

BUFx12_ASAP7_75t_L g121 ( 
.A(n_43),
.Y(n_121)
);

INVx3_ASAP7_75t_L g122 ( 
.A(n_43),
.Y(n_122)
);

INVx2_ASAP7_75t_L g189 ( 
.A(n_122),
.Y(n_189)
);

INVx5_ASAP7_75t_L g123 ( 
.A(n_20),
.Y(n_123)
);

INVx2_ASAP7_75t_L g199 ( 
.A(n_123),
.Y(n_199)
);

INVx2_ASAP7_75t_L g124 ( 
.A(n_47),
.Y(n_124)
);

INVx2_ASAP7_75t_L g200 ( 
.A(n_124),
.Y(n_200)
);

INVx6_ASAP7_75t_L g125 ( 
.A(n_53),
.Y(n_125)
);

INVx2_ASAP7_75t_L g209 ( 
.A(n_125),
.Y(n_209)
);

INVx8_ASAP7_75t_L g126 ( 
.A(n_53),
.Y(n_126)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_126),
.Y(n_175)
);

INVx6_ASAP7_75t_L g127 ( 
.A(n_20),
.Y(n_127)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_127),
.Y(n_184)
);

CKINVDCx16_ASAP7_75t_R g128 ( 
.A(n_43),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_L g192 ( 
.A(n_128),
.B(n_129),
.Y(n_192)
);

NOR2xp33_ASAP7_75t_SL g129 ( 
.A(n_21),
.B(n_2),
.Y(n_129)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_49),
.Y(n_130)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_130),
.Y(n_194)
);

AOI22xp33_ASAP7_75t_SL g137 ( 
.A1(n_101),
.A2(n_52),
.B1(n_43),
.B2(n_45),
.Y(n_137)
);

AOI21xp5_ASAP7_75t_L g235 ( 
.A1(n_137),
.A2(n_142),
.B(n_147),
.Y(n_235)
);

OAI22xp5_ASAP7_75t_L g141 ( 
.A1(n_107),
.A2(n_62),
.B1(n_29),
.B2(n_30),
.Y(n_141)
);

AOI22xp5_ASAP7_75t_L g260 ( 
.A1(n_141),
.A2(n_180),
.B1(n_196),
.B2(n_204),
.Y(n_260)
);

AOI22xp33_ASAP7_75t_SL g142 ( 
.A1(n_83),
.A2(n_52),
.B1(n_45),
.B2(n_25),
.Y(n_142)
);

AOI22xp33_ASAP7_75t_SL g147 ( 
.A1(n_127),
.A2(n_52),
.B1(n_45),
.B2(n_25),
.Y(n_147)
);

AND2x2_ASAP7_75t_L g149 ( 
.A(n_74),
.B(n_45),
.Y(n_149)
);

OAI21xp5_ASAP7_75t_SL g286 ( 
.A1(n_149),
.A2(n_167),
.B(n_33),
.Y(n_286)
);

MAJIxp5_ASAP7_75t_L g162 ( 
.A(n_84),
.B(n_60),
.C(n_59),
.Y(n_162)
);

MAJIxp5_ASAP7_75t_L g226 ( 
.A(n_162),
.B(n_29),
.C(n_22),
.Y(n_226)
);

AOI22xp33_ASAP7_75t_L g163 ( 
.A1(n_85),
.A2(n_52),
.B1(n_25),
.B2(n_28),
.Y(n_163)
);

OAI22xp5_ASAP7_75t_SL g263 ( 
.A1(n_163),
.A2(n_166),
.B1(n_142),
.B2(n_176),
.Y(n_263)
);

AOI22xp33_ASAP7_75t_L g166 ( 
.A1(n_125),
.A2(n_28),
.B1(n_31),
.B2(n_59),
.Y(n_166)
);

AND2x2_ASAP7_75t_L g167 ( 
.A(n_86),
.B(n_45),
.Y(n_167)
);

OAI22xp5_ASAP7_75t_L g180 ( 
.A1(n_68),
.A2(n_24),
.B1(n_48),
.B2(n_46),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_SL g193 ( 
.A(n_106),
.B(n_24),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_L g248 ( 
.A(n_193),
.B(n_201),
.Y(n_248)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_126),
.Y(n_195)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_195),
.Y(n_217)
);

OAI22xp33_ASAP7_75t_SL g196 ( 
.A1(n_70),
.A2(n_31),
.B1(n_28),
.B2(n_57),
.Y(n_196)
);

NAND2xp5_ASAP7_75t_SL g201 ( 
.A(n_80),
.B(n_23),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_L g203 ( 
.A(n_72),
.B(n_23),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_L g250 ( 
.A(n_203),
.B(n_207),
.Y(n_250)
);

OAI22xp5_ASAP7_75t_SL g204 ( 
.A1(n_88),
.A2(n_94),
.B1(n_119),
.B2(n_117),
.Y(n_204)
);

OAI22xp5_ASAP7_75t_L g206 ( 
.A1(n_97),
.A2(n_22),
.B1(n_48),
.B2(n_46),
.Y(n_206)
);

AOI22xp5_ASAP7_75t_SL g215 ( 
.A1(n_206),
.A2(n_212),
.B1(n_108),
.B2(n_34),
.Y(n_215)
);

NAND2xp5_ASAP7_75t_L g207 ( 
.A(n_98),
.B(n_21),
.Y(n_207)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_100),
.Y(n_211)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_211),
.Y(n_218)
);

AOI22xp33_ASAP7_75t_SL g212 ( 
.A1(n_63),
.A2(n_31),
.B1(n_58),
.B2(n_57),
.Y(n_212)
);

NAND2xp5_ASAP7_75t_SL g213 ( 
.A(n_80),
.B(n_62),
.Y(n_213)
);

NAND2xp5_ASAP7_75t_L g290 ( 
.A(n_213),
.B(n_214),
.Y(n_290)
);

NAND2xp5_ASAP7_75t_L g214 ( 
.A(n_104),
.B(n_34),
.Y(n_214)
);

OAI22xp5_ASAP7_75t_L g307 ( 
.A1(n_215),
.A2(n_289),
.B1(n_187),
.B2(n_150),
.Y(n_307)
);

INVx4_ASAP7_75t_L g216 ( 
.A(n_134),
.Y(n_216)
);

INVx3_ASAP7_75t_L g352 ( 
.A(n_216),
.Y(n_352)
);

INVx1_ASAP7_75t_SL g219 ( 
.A(n_146),
.Y(n_219)
);

INVx1_ASAP7_75t_SL g295 ( 
.A(n_219),
.Y(n_295)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_133),
.Y(n_220)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_220),
.Y(n_291)
);

NOR2xp33_ASAP7_75t_L g221 ( 
.A(n_192),
.B(n_58),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_SL g318 ( 
.A(n_221),
.B(n_224),
.Y(n_318)
);

HB1xp67_ASAP7_75t_L g222 ( 
.A(n_210),
.Y(n_222)
);

HB1xp67_ASAP7_75t_L g345 ( 
.A(n_222),
.Y(n_345)
);

INVx5_ASAP7_75t_L g223 ( 
.A(n_135),
.Y(n_223)
);

HB1xp67_ASAP7_75t_L g351 ( 
.A(n_223),
.Y(n_351)
);

NOR2xp33_ASAP7_75t_L g224 ( 
.A(n_139),
.B(n_60),
.Y(n_224)
);

INVx2_ASAP7_75t_SL g225 ( 
.A(n_151),
.Y(n_225)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_225),
.Y(n_293)
);

NOR2xp33_ASAP7_75t_L g301 ( 
.A(n_226),
.B(n_229),
.Y(n_301)
);

INVx4_ASAP7_75t_L g227 ( 
.A(n_174),
.Y(n_227)
);

INVx2_ASAP7_75t_L g308 ( 
.A(n_227),
.Y(n_308)
);

BUFx2_ASAP7_75t_SL g228 ( 
.A(n_165),
.Y(n_228)
);

INVxp67_ASAP7_75t_L g303 ( 
.A(n_228),
.Y(n_303)
);

CKINVDCx20_ASAP7_75t_R g229 ( 
.A(n_152),
.Y(n_229)
);

OAI22xp33_ASAP7_75t_SL g230 ( 
.A1(n_147),
.A2(n_111),
.B1(n_109),
.B2(n_92),
.Y(n_230)
);

AOI22xp5_ASAP7_75t_L g347 ( 
.A1(n_230),
.A2(n_252),
.B1(n_263),
.B2(n_273),
.Y(n_347)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_140),
.Y(n_231)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_231),
.Y(n_296)
);

INVx4_ASAP7_75t_L g232 ( 
.A(n_188),
.Y(n_232)
);

INVx2_ASAP7_75t_L g314 ( 
.A(n_232),
.Y(n_314)
);

INVx2_ASAP7_75t_L g233 ( 
.A(n_131),
.Y(n_233)
);

INVx2_ASAP7_75t_L g317 ( 
.A(n_233),
.Y(n_317)
);

INVx4_ASAP7_75t_L g234 ( 
.A(n_190),
.Y(n_234)
);

INVx2_ASAP7_75t_L g321 ( 
.A(n_234),
.Y(n_321)
);

BUFx6f_ASAP7_75t_L g236 ( 
.A(n_132),
.Y(n_236)
);

INVx6_ASAP7_75t_L g311 ( 
.A(n_236),
.Y(n_311)
);

INVx2_ASAP7_75t_L g237 ( 
.A(n_136),
.Y(n_237)
);

INVx2_ASAP7_75t_L g329 ( 
.A(n_237),
.Y(n_329)
);

NOR2xp33_ASAP7_75t_L g238 ( 
.A(n_170),
.B(n_41),
.Y(n_238)
);

NAND2xp5_ASAP7_75t_SL g334 ( 
.A(n_238),
.B(n_242),
.Y(n_334)
);

BUFx3_ASAP7_75t_L g239 ( 
.A(n_210),
.Y(n_239)
);

BUFx3_ASAP7_75t_L g346 ( 
.A(n_239),
.Y(n_346)
);

INVx2_ASAP7_75t_L g240 ( 
.A(n_143),
.Y(n_240)
);

INVx2_ASAP7_75t_L g330 ( 
.A(n_240),
.Y(n_330)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_153),
.Y(n_241)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_241),
.Y(n_300)
);

NOR2xp33_ASAP7_75t_SL g242 ( 
.A(n_164),
.B(n_37),
.Y(n_242)
);

INVxp67_ASAP7_75t_L g243 ( 
.A(n_212),
.Y(n_243)
);

NOR2xp33_ASAP7_75t_L g306 ( 
.A(n_243),
.B(n_246),
.Y(n_306)
);

INVx4_ASAP7_75t_L g244 ( 
.A(n_171),
.Y(n_244)
);

INVx2_ASAP7_75t_L g339 ( 
.A(n_244),
.Y(n_339)
);

INVx2_ASAP7_75t_L g245 ( 
.A(n_169),
.Y(n_245)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_245),
.Y(n_304)
);

CKINVDCx20_ASAP7_75t_R g246 ( 
.A(n_166),
.Y(n_246)
);

INVx3_ASAP7_75t_L g247 ( 
.A(n_175),
.Y(n_247)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_247),
.Y(n_326)
);

INVxp67_ASAP7_75t_L g249 ( 
.A(n_167),
.Y(n_249)
);

NOR2xp33_ASAP7_75t_L g320 ( 
.A(n_249),
.B(n_254),
.Y(n_320)
);

INVx2_ASAP7_75t_L g251 ( 
.A(n_200),
.Y(n_251)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_251),
.Y(n_336)
);

OAI22xp33_ASAP7_75t_SL g252 ( 
.A1(n_137),
.A2(n_87),
.B1(n_95),
.B2(n_120),
.Y(n_252)
);

INVx3_ASAP7_75t_L g253 ( 
.A(n_171),
.Y(n_253)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_253),
.Y(n_337)
);

NOR2xp33_ASAP7_75t_L g254 ( 
.A(n_155),
.B(n_41),
.Y(n_254)
);

INVx2_ASAP7_75t_L g255 ( 
.A(n_209),
.Y(n_255)
);

INVx1_ASAP7_75t_L g348 ( 
.A(n_255),
.Y(n_348)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_159),
.Y(n_256)
);

NOR2xp33_ASAP7_75t_L g343 ( 
.A(n_256),
.B(n_257),
.Y(n_343)
);

CKINVDCx20_ASAP7_75t_R g257 ( 
.A(n_163),
.Y(n_257)
);

INVx11_ASAP7_75t_L g258 ( 
.A(n_145),
.Y(n_258)
);

INVx8_ASAP7_75t_L g292 ( 
.A(n_258),
.Y(n_292)
);

BUFx6f_ASAP7_75t_L g259 ( 
.A(n_132),
.Y(n_259)
);

AOI22xp33_ASAP7_75t_SL g316 ( 
.A1(n_259),
.A2(n_275),
.B1(n_277),
.B2(n_279),
.Y(n_316)
);

INVx3_ASAP7_75t_L g261 ( 
.A(n_199),
.Y(n_261)
);

AND2x2_ASAP7_75t_L g322 ( 
.A(n_261),
.B(n_265),
.Y(n_322)
);

CKINVDCx14_ASAP7_75t_R g262 ( 
.A(n_165),
.Y(n_262)
);

OR2x2_ASAP7_75t_L g342 ( 
.A(n_262),
.B(n_267),
.Y(n_342)
);

CKINVDCx20_ASAP7_75t_R g264 ( 
.A(n_172),
.Y(n_264)
);

CKINVDCx20_ASAP7_75t_R g309 ( 
.A(n_264),
.Y(n_309)
);

NOR2xp33_ASAP7_75t_L g265 ( 
.A(n_173),
.B(n_37),
.Y(n_265)
);

INVx2_ASAP7_75t_L g266 ( 
.A(n_154),
.Y(n_266)
);

AND2x2_ASAP7_75t_L g335 ( 
.A(n_266),
.B(n_268),
.Y(n_335)
);

CKINVDCx5p33_ASAP7_75t_R g267 ( 
.A(n_197),
.Y(n_267)
);

INVx5_ASAP7_75t_L g268 ( 
.A(n_135),
.Y(n_268)
);

AND2x2_ASAP7_75t_L g269 ( 
.A(n_149),
.B(n_93),
.Y(n_269)
);

MAJIxp5_ASAP7_75t_L g299 ( 
.A(n_269),
.B(n_270),
.C(n_274),
.Y(n_299)
);

AND2x2_ASAP7_75t_L g270 ( 
.A(n_194),
.B(n_2),
.Y(n_270)
);

INVx2_ASAP7_75t_L g271 ( 
.A(n_183),
.Y(n_271)
);

CKINVDCx20_ASAP7_75t_R g324 ( 
.A(n_271),
.Y(n_324)
);

INVxp67_ASAP7_75t_L g272 ( 
.A(n_184),
.Y(n_272)
);

CKINVDCx20_ASAP7_75t_R g333 ( 
.A(n_272),
.Y(n_333)
);

OAI22xp5_ASAP7_75t_SL g273 ( 
.A1(n_177),
.A2(n_36),
.B1(n_33),
.B2(n_30),
.Y(n_273)
);

AND2x2_ASAP7_75t_L g274 ( 
.A(n_157),
.B(n_3),
.Y(n_274)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_185),
.Y(n_275)
);

CKINVDCx16_ASAP7_75t_R g276 ( 
.A(n_145),
.Y(n_276)
);

NAND2xp5_ASAP7_75t_L g294 ( 
.A(n_276),
.B(n_280),
.Y(n_294)
);

INVx5_ASAP7_75t_L g277 ( 
.A(n_144),
.Y(n_277)
);

MAJIxp5_ASAP7_75t_L g278 ( 
.A(n_189),
.B(n_121),
.C(n_115),
.Y(n_278)
);

XNOR2xp5_ASAP7_75t_L g327 ( 
.A(n_278),
.B(n_168),
.Y(n_327)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_179),
.Y(n_279)
);

CKINVDCx20_ASAP7_75t_R g280 ( 
.A(n_182),
.Y(n_280)
);

NOR2xp33_ASAP7_75t_L g281 ( 
.A(n_144),
.B(n_36),
.Y(n_281)
);

NAND2xp5_ASAP7_75t_L g297 ( 
.A(n_281),
.B(n_288),
.Y(n_297)
);

BUFx12f_ASAP7_75t_L g282 ( 
.A(n_138),
.Y(n_282)
);

AOI22xp33_ASAP7_75t_SL g328 ( 
.A1(n_282),
.A2(n_283),
.B1(n_284),
.B2(n_285),
.Y(n_328)
);

INVx2_ASAP7_75t_L g283 ( 
.A(n_186),
.Y(n_283)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_191),
.Y(n_284)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_205),
.Y(n_285)
);

AND2x2_ASAP7_75t_SL g305 ( 
.A(n_286),
.B(n_197),
.Y(n_305)
);

INVx2_ASAP7_75t_L g287 ( 
.A(n_160),
.Y(n_287)
);

AOI22xp33_ASAP7_75t_SL g332 ( 
.A1(n_287),
.A2(n_158),
.B1(n_208),
.B2(n_156),
.Y(n_332)
);

CKINVDCx20_ASAP7_75t_R g288 ( 
.A(n_176),
.Y(n_288)
);

AOI22xp33_ASAP7_75t_L g289 ( 
.A1(n_196),
.A2(n_3),
.B1(n_4),
.B2(n_7),
.Y(n_289)
);

NAND2xp5_ASAP7_75t_L g298 ( 
.A(n_250),
.B(n_198),
.Y(n_298)
);

NAND2xp5_ASAP7_75t_L g365 ( 
.A(n_298),
.B(n_310),
.Y(n_365)
);

OAI22xp5_ASAP7_75t_SL g302 ( 
.A1(n_260),
.A2(n_243),
.B1(n_235),
.B2(n_215),
.Y(n_302)
);

AOI22xp5_ASAP7_75t_L g362 ( 
.A1(n_302),
.A2(n_307),
.B1(n_313),
.B2(n_315),
.Y(n_362)
);

OAI21xp33_ASAP7_75t_L g382 ( 
.A1(n_305),
.A2(n_232),
.B(n_216),
.Y(n_382)
);

NAND2xp5_ASAP7_75t_L g310 ( 
.A(n_270),
.B(n_198),
.Y(n_310)
);

XOR2xp5_ASAP7_75t_L g312 ( 
.A(n_290),
.B(n_148),
.Y(n_312)
);

MAJIxp5_ASAP7_75t_L g377 ( 
.A(n_312),
.B(n_225),
.C(n_240),
.Y(n_377)
);

OAI22xp5_ASAP7_75t_SL g313 ( 
.A1(n_260),
.A2(n_160),
.B1(n_202),
.B2(n_181),
.Y(n_313)
);

OAI22xp5_ASAP7_75t_SL g315 ( 
.A1(n_235),
.A2(n_178),
.B1(n_202),
.B2(n_181),
.Y(n_315)
);

NAND2xp5_ASAP7_75t_L g319 ( 
.A(n_270),
.B(n_148),
.Y(n_319)
);

NAND2xp5_ASAP7_75t_L g389 ( 
.A(n_319),
.B(n_349),
.Y(n_389)
);

OAI21xp5_ASAP7_75t_SL g323 ( 
.A1(n_269),
.A2(n_156),
.B(n_4),
.Y(n_323)
);

AOI21xp5_ASAP7_75t_L g368 ( 
.A1(n_323),
.A2(n_341),
.B(n_223),
.Y(n_368)
);

OAI22xp5_ASAP7_75t_L g325 ( 
.A1(n_248),
.A2(n_178),
.B1(n_168),
.B2(n_161),
.Y(n_325)
);

AOI22xp5_ASAP7_75t_L g364 ( 
.A1(n_325),
.A2(n_331),
.B1(n_338),
.B2(n_219),
.Y(n_364)
);

XNOR2xp5_ASAP7_75t_L g383 ( 
.A(n_327),
.B(n_253),
.Y(n_383)
);

OAI22xp5_ASAP7_75t_L g331 ( 
.A1(n_249),
.A2(n_161),
.B1(n_158),
.B2(n_138),
.Y(n_331)
);

INVxp67_ASAP7_75t_L g363 ( 
.A(n_332),
.Y(n_363)
);

OAI22xp5_ASAP7_75t_SL g338 ( 
.A1(n_263),
.A2(n_208),
.B1(n_7),
.B2(n_8),
.Y(n_338)
);

AOI22xp33_ASAP7_75t_L g340 ( 
.A1(n_273),
.A2(n_3),
.B1(n_7),
.B2(n_8),
.Y(n_340)
);

OAI22xp5_ASAP7_75t_L g391 ( 
.A1(n_340),
.A2(n_12),
.B1(n_16),
.B2(n_341),
.Y(n_391)
);

AOI21xp5_ASAP7_75t_L g341 ( 
.A1(n_269),
.A2(n_9),
.B(n_10),
.Y(n_341)
);

A2O1A1Ixp33_ASAP7_75t_L g344 ( 
.A1(n_226),
.A2(n_10),
.B(n_11),
.C(n_12),
.Y(n_344)
);

NOR2x1_ASAP7_75t_L g381 ( 
.A(n_344),
.B(n_350),
.Y(n_381)
);

NAND2xp5_ASAP7_75t_L g349 ( 
.A(n_274),
.B(n_233),
.Y(n_349)
);

AOI32xp33_ASAP7_75t_L g350 ( 
.A1(n_267),
.A2(n_10),
.A3(n_12),
.B1(n_13),
.B2(n_14),
.Y(n_350)
);

OAI21xp33_ASAP7_75t_SL g353 ( 
.A1(n_319),
.A2(n_268),
.B(n_277),
.Y(n_353)
);

OAI21xp5_ASAP7_75t_SL g440 ( 
.A1(n_353),
.A2(n_368),
.B(n_398),
.Y(n_440)
);

OAI22xp5_ASAP7_75t_L g354 ( 
.A1(n_347),
.A2(n_278),
.B1(n_287),
.B2(n_259),
.Y(n_354)
);

AOI22xp5_ASAP7_75t_L g403 ( 
.A1(n_354),
.A2(n_372),
.B1(n_374),
.B2(n_387),
.Y(n_403)
);

INVx1_ASAP7_75t_L g355 ( 
.A(n_304),
.Y(n_355)
);

INVx1_ASAP7_75t_L g408 ( 
.A(n_355),
.Y(n_408)
);

INVx1_ASAP7_75t_L g356 ( 
.A(n_304),
.Y(n_356)
);

INVx1_ASAP7_75t_L g411 ( 
.A(n_356),
.Y(n_411)
);

FAx1_ASAP7_75t_SL g357 ( 
.A(n_299),
.B(n_274),
.CI(n_258),
.CON(n_357),
.SN(n_357)
);

NOR2xp33_ASAP7_75t_SL g414 ( 
.A(n_357),
.B(n_375),
.Y(n_414)
);

INVx1_ASAP7_75t_L g358 ( 
.A(n_291),
.Y(n_358)
);

INVx1_ASAP7_75t_L g413 ( 
.A(n_358),
.Y(n_413)
);

NOR2xp33_ASAP7_75t_L g359 ( 
.A(n_309),
.B(n_318),
.Y(n_359)
);

NAND2xp5_ASAP7_75t_SL g406 ( 
.A(n_359),
.B(n_360),
.Y(n_406)
);

NAND2xp5_ASAP7_75t_SL g360 ( 
.A(n_309),
.B(n_217),
.Y(n_360)
);

NOR2xp33_ASAP7_75t_L g361 ( 
.A(n_297),
.B(n_239),
.Y(n_361)
);

NAND2xp5_ASAP7_75t_SL g429 ( 
.A(n_361),
.B(n_366),
.Y(n_429)
);

AND2x2_ASAP7_75t_L g435 ( 
.A(n_364),
.B(n_382),
.Y(n_435)
);

CKINVDCx16_ASAP7_75t_R g366 ( 
.A(n_294),
.Y(n_366)
);

AOI22xp5_ASAP7_75t_L g367 ( 
.A1(n_302),
.A2(n_313),
.B1(n_315),
.B2(n_338),
.Y(n_367)
);

OAI22xp5_ASAP7_75t_L g431 ( 
.A1(n_367),
.A2(n_385),
.B1(n_388),
.B2(n_397),
.Y(n_431)
);

INVx1_ASAP7_75t_L g369 ( 
.A(n_291),
.Y(n_369)
);

INVx1_ASAP7_75t_L g417 ( 
.A(n_369),
.Y(n_417)
);

CKINVDCx16_ASAP7_75t_R g370 ( 
.A(n_294),
.Y(n_370)
);

NAND2xp5_ASAP7_75t_SL g436 ( 
.A(n_370),
.B(n_384),
.Y(n_436)
);

CKINVDCx6p67_ASAP7_75t_R g371 ( 
.A(n_303),
.Y(n_371)
);

INVx4_ASAP7_75t_L g425 ( 
.A(n_371),
.Y(n_425)
);

OAI22xp5_ASAP7_75t_L g372 ( 
.A1(n_347),
.A2(n_236),
.B1(n_271),
.B2(n_266),
.Y(n_372)
);

INVx1_ASAP7_75t_L g373 ( 
.A(n_296),
.Y(n_373)
);

INVx1_ASAP7_75t_L g421 ( 
.A(n_373),
.Y(n_421)
);

OAI22xp5_ASAP7_75t_SL g374 ( 
.A1(n_306),
.A2(n_283),
.B1(n_218),
.B2(n_261),
.Y(n_374)
);

FAx1_ASAP7_75t_SL g375 ( 
.A(n_299),
.B(n_272),
.CI(n_237),
.CON(n_375),
.SN(n_375)
);

INVx2_ASAP7_75t_SL g376 ( 
.A(n_335),
.Y(n_376)
);

INVx2_ASAP7_75t_L g412 ( 
.A(n_376),
.Y(n_412)
);

MAJIxp5_ASAP7_75t_L g426 ( 
.A(n_377),
.B(n_380),
.C(n_383),
.Y(n_426)
);

INVx1_ASAP7_75t_L g378 ( 
.A(n_296),
.Y(n_378)
);

INVx1_ASAP7_75t_L g430 ( 
.A(n_378),
.Y(n_430)
);

INVx1_ASAP7_75t_L g379 ( 
.A(n_300),
.Y(n_379)
);

INVx1_ASAP7_75t_L g434 ( 
.A(n_379),
.Y(n_434)
);

MAJIxp5_ASAP7_75t_L g380 ( 
.A(n_312),
.B(n_245),
.C(n_247),
.Y(n_380)
);

CKINVDCx16_ASAP7_75t_R g384 ( 
.A(n_335),
.Y(n_384)
);

AOI22xp5_ASAP7_75t_L g385 ( 
.A1(n_298),
.A2(n_310),
.B1(n_349),
.B2(n_305),
.Y(n_385)
);

NOR2xp33_ASAP7_75t_L g386 ( 
.A(n_297),
.B(n_227),
.Y(n_386)
);

INVxp67_ASAP7_75t_L g402 ( 
.A(n_386),
.Y(n_402)
);

OAI22xp5_ASAP7_75t_SL g387 ( 
.A1(n_343),
.A2(n_234),
.B1(n_282),
.B2(n_244),
.Y(n_387)
);

AOI22xp33_ASAP7_75t_L g388 ( 
.A1(n_322),
.A2(n_282),
.B1(n_15),
.B2(n_16),
.Y(n_388)
);

INVx1_ASAP7_75t_L g390 ( 
.A(n_300),
.Y(n_390)
);

INVx1_ASAP7_75t_L g441 ( 
.A(n_390),
.Y(n_441)
);

AOI22xp5_ASAP7_75t_L g404 ( 
.A1(n_391),
.A2(n_394),
.B1(n_295),
.B2(n_303),
.Y(n_404)
);

NOR2xp33_ASAP7_75t_L g392 ( 
.A(n_301),
.B(n_320),
.Y(n_392)
);

CKINVDCx16_ASAP7_75t_R g427 ( 
.A(n_392),
.Y(n_427)
);

MAJIxp5_ASAP7_75t_L g393 ( 
.A(n_327),
.B(n_305),
.C(n_322),
.Y(n_393)
);

NAND2xp5_ASAP7_75t_L g410 ( 
.A(n_393),
.B(n_396),
.Y(n_410)
);

OAI22xp5_ASAP7_75t_L g394 ( 
.A1(n_342),
.A2(n_333),
.B1(n_316),
.B2(n_295),
.Y(n_394)
);

CKINVDCx16_ASAP7_75t_R g395 ( 
.A(n_335),
.Y(n_395)
);

INVx1_ASAP7_75t_SL g401 ( 
.A(n_395),
.Y(n_401)
);

NAND2xp5_ASAP7_75t_L g396 ( 
.A(n_322),
.B(n_333),
.Y(n_396)
);

AOI22xp5_ASAP7_75t_L g397 ( 
.A1(n_293),
.A2(n_324),
.B1(n_344),
.B2(n_336),
.Y(n_397)
);

CKINVDCx14_ASAP7_75t_R g398 ( 
.A(n_342),
.Y(n_398)
);

MAJIxp5_ASAP7_75t_L g399 ( 
.A(n_323),
.B(n_336),
.C(n_345),
.Y(n_399)
);

NAND2xp5_ASAP7_75t_L g415 ( 
.A(n_399),
.B(n_400),
.Y(n_415)
);

MAJIxp5_ASAP7_75t_L g400 ( 
.A(n_348),
.B(n_326),
.C(n_337),
.Y(n_400)
);

NAND2xp5_ASAP7_75t_L g471 ( 
.A(n_404),
.B(n_407),
.Y(n_471)
);

CKINVDCx20_ASAP7_75t_R g405 ( 
.A(n_400),
.Y(n_405)
);

NOR2xp33_ASAP7_75t_L g453 ( 
.A(n_405),
.B(n_422),
.Y(n_453)
);

OAI32xp33_ASAP7_75t_L g407 ( 
.A1(n_365),
.A2(n_334),
.A3(n_293),
.B1(n_337),
.B2(n_326),
.Y(n_407)
);

OAI22x1_ASAP7_75t_SL g409 ( 
.A1(n_362),
.A2(n_328),
.B1(n_352),
.B2(n_314),
.Y(n_409)
);

NAND2xp5_ASAP7_75t_L g476 ( 
.A(n_409),
.B(n_416),
.Y(n_476)
);

OAI32xp33_ASAP7_75t_L g416 ( 
.A1(n_365),
.A2(n_292),
.A3(n_348),
.B1(n_308),
.B2(n_314),
.Y(n_416)
);

AOI21xp5_ASAP7_75t_L g418 ( 
.A1(n_363),
.A2(n_352),
.B(n_308),
.Y(n_418)
);

AOI21xp5_ASAP7_75t_L g465 ( 
.A1(n_418),
.A2(n_432),
.B(n_371),
.Y(n_465)
);

OAI21xp5_ASAP7_75t_L g419 ( 
.A1(n_396),
.A2(n_324),
.B(n_321),
.Y(n_419)
);

OAI21xp5_ASAP7_75t_L g445 ( 
.A1(n_419),
.A2(n_368),
.B(n_356),
.Y(n_445)
);

AOI22xp5_ASAP7_75t_L g420 ( 
.A1(n_354),
.A2(n_311),
.B1(n_321),
.B2(n_317),
.Y(n_420)
);

OAI22xp5_ASAP7_75t_SL g442 ( 
.A1(n_420),
.A2(n_424),
.B1(n_364),
.B2(n_355),
.Y(n_442)
);

CKINVDCx20_ASAP7_75t_R g422 ( 
.A(n_387),
.Y(n_422)
);

CKINVDCx20_ASAP7_75t_R g423 ( 
.A(n_374),
.Y(n_423)
);

NOR2xp33_ASAP7_75t_L g462 ( 
.A(n_423),
.B(n_433),
.Y(n_462)
);

AOI22xp5_ASAP7_75t_L g424 ( 
.A1(n_372),
.A2(n_311),
.B1(n_330),
.B2(n_317),
.Y(n_424)
);

BUFx5_ASAP7_75t_L g428 ( 
.A(n_371),
.Y(n_428)
);

INVx2_ASAP7_75t_L g444 ( 
.A(n_428),
.Y(n_444)
);

AOI21xp5_ASAP7_75t_L g432 ( 
.A1(n_363),
.A2(n_351),
.B(n_339),
.Y(n_432)
);

NAND2xp5_ASAP7_75t_L g433 ( 
.A(n_389),
.B(n_329),
.Y(n_433)
);

NAND2xp5_ASAP7_75t_L g437 ( 
.A(n_389),
.B(n_329),
.Y(n_437)
);

NOR2xp33_ASAP7_75t_L g474 ( 
.A(n_437),
.B(n_379),
.Y(n_474)
);

AND2x2_ASAP7_75t_L g438 ( 
.A(n_376),
.B(n_292),
.Y(n_438)
);

OAI21xp5_ASAP7_75t_SL g452 ( 
.A1(n_438),
.A2(n_439),
.B(n_339),
.Y(n_452)
);

AND2x2_ASAP7_75t_L g439 ( 
.A(n_376),
.B(n_330),
.Y(n_439)
);

INVx1_ASAP7_75t_L g509 ( 
.A(n_442),
.Y(n_509)
);

OAI22xp5_ASAP7_75t_SL g443 ( 
.A1(n_403),
.A2(n_367),
.B1(n_362),
.B2(n_385),
.Y(n_443)
);

AOI22xp5_ASAP7_75t_L g490 ( 
.A1(n_443),
.A2(n_451),
.B1(n_431),
.B2(n_409),
.Y(n_490)
);

INVxp67_ASAP7_75t_L g507 ( 
.A(n_445),
.Y(n_507)
);

XOR2xp5_ASAP7_75t_L g446 ( 
.A(n_426),
.B(n_383),
.Y(n_446)
);

MAJIxp5_ASAP7_75t_L g482 ( 
.A(n_446),
.B(n_455),
.C(n_459),
.Y(n_482)
);

CKINVDCx20_ASAP7_75t_R g447 ( 
.A(n_429),
.Y(n_447)
);

NAND2xp5_ASAP7_75t_L g495 ( 
.A(n_447),
.B(n_452),
.Y(n_495)
);

OA21x2_ASAP7_75t_L g448 ( 
.A1(n_435),
.A2(n_397),
.B(n_394),
.Y(n_448)
);

OAI21xp5_ASAP7_75t_SL g501 ( 
.A1(n_448),
.A2(n_465),
.B(n_468),
.Y(n_501)
);

XNOR2xp5_ASAP7_75t_SL g449 ( 
.A(n_426),
.B(n_393),
.Y(n_449)
);

XOR2xp5_ASAP7_75t_L g479 ( 
.A(n_449),
.B(n_407),
.Y(n_479)
);

INVx1_ASAP7_75t_L g450 ( 
.A(n_413),
.Y(n_450)
);

INVx1_ASAP7_75t_SL g506 ( 
.A(n_450),
.Y(n_506)
);

OAI22xp5_ASAP7_75t_SL g451 ( 
.A1(n_403),
.A2(n_377),
.B1(n_380),
.B2(n_399),
.Y(n_451)
);

OR2x2_ASAP7_75t_L g454 ( 
.A(n_440),
.B(n_414),
.Y(n_454)
);

CKINVDCx20_ASAP7_75t_R g485 ( 
.A(n_454),
.Y(n_485)
);

MAJIxp5_ASAP7_75t_L g455 ( 
.A(n_410),
.B(n_375),
.C(n_357),
.Y(n_455)
);

CKINVDCx20_ASAP7_75t_R g456 ( 
.A(n_433),
.Y(n_456)
);

NAND2xp5_ASAP7_75t_L g502 ( 
.A(n_456),
.B(n_458),
.Y(n_502)
);

NAND3xp33_ASAP7_75t_L g457 ( 
.A(n_406),
.B(n_375),
.C(n_390),
.Y(n_457)
);

NOR2xp33_ASAP7_75t_L g494 ( 
.A(n_457),
.B(n_472),
.Y(n_494)
);

INVx1_ASAP7_75t_L g458 ( 
.A(n_413),
.Y(n_458)
);

XOR2xp5_ASAP7_75t_L g459 ( 
.A(n_410),
.B(n_357),
.Y(n_459)
);

NOR2xp33_ASAP7_75t_SL g460 ( 
.A(n_427),
.B(n_402),
.Y(n_460)
);

NOR2xp33_ASAP7_75t_SL g508 ( 
.A(n_460),
.B(n_475),
.Y(n_508)
);

INVx1_ASAP7_75t_L g461 ( 
.A(n_417),
.Y(n_461)
);

NAND2xp5_ASAP7_75t_L g504 ( 
.A(n_461),
.B(n_466),
.Y(n_504)
);

OAI21xp5_ASAP7_75t_SL g463 ( 
.A1(n_435),
.A2(n_381),
.B(n_371),
.Y(n_463)
);

AOI21xp5_ASAP7_75t_L g483 ( 
.A1(n_463),
.A2(n_435),
.B(n_414),
.Y(n_483)
);

MAJIxp5_ASAP7_75t_L g464 ( 
.A(n_415),
.B(n_373),
.C(n_358),
.Y(n_464)
);

MAJIxp5_ASAP7_75t_L g484 ( 
.A(n_464),
.B(n_470),
.C(n_477),
.Y(n_484)
);

CKINVDCx20_ASAP7_75t_R g466 ( 
.A(n_437),
.Y(n_466)
);

NOR2xp33_ASAP7_75t_L g467 ( 
.A(n_436),
.B(n_369),
.Y(n_467)
);

NAND2xp5_ASAP7_75t_SL g486 ( 
.A(n_467),
.B(n_469),
.Y(n_486)
);

AOI21xp5_ASAP7_75t_L g468 ( 
.A1(n_440),
.A2(n_381),
.B(n_378),
.Y(n_468)
);

CKINVDCx16_ASAP7_75t_R g469 ( 
.A(n_419),
.Y(n_469)
);

MAJIxp5_ASAP7_75t_L g470 ( 
.A(n_415),
.B(n_405),
.C(n_401),
.Y(n_470)
);

INVx1_ASAP7_75t_L g472 ( 
.A(n_417),
.Y(n_472)
);

INVx1_ASAP7_75t_L g473 ( 
.A(n_421),
.Y(n_473)
);

NAND2xp5_ASAP7_75t_SL g488 ( 
.A(n_473),
.B(n_441),
.Y(n_488)
);

CKINVDCx14_ASAP7_75t_R g503 ( 
.A(n_474),
.Y(n_503)
);

NOR2xp33_ASAP7_75t_L g475 ( 
.A(n_421),
.B(n_346),
.Y(n_475)
);

XNOR2xp5_ASAP7_75t_L g477 ( 
.A(n_401),
.B(n_346),
.Y(n_477)
);

CKINVDCx20_ASAP7_75t_R g478 ( 
.A(n_439),
.Y(n_478)
);

CKINVDCx20_ASAP7_75t_R g489 ( 
.A(n_478),
.Y(n_489)
);

XNOR2xp5_ASAP7_75t_SL g521 ( 
.A(n_479),
.B(n_471),
.Y(n_521)
);

INVx3_ASAP7_75t_L g480 ( 
.A(n_444),
.Y(n_480)
);

INVx1_ASAP7_75t_L g523 ( 
.A(n_480),
.Y(n_523)
);

OAI22xp5_ASAP7_75t_L g481 ( 
.A1(n_453),
.A2(n_422),
.B1(n_404),
.B2(n_423),
.Y(n_481)
);

AOI22xp5_ASAP7_75t_L g522 ( 
.A1(n_481),
.A2(n_491),
.B1(n_493),
.B2(n_499),
.Y(n_522)
);

AOI21xp5_ASAP7_75t_L g531 ( 
.A1(n_483),
.A2(n_445),
.B(n_463),
.Y(n_531)
);

XOR2xp5_ASAP7_75t_L g487 ( 
.A(n_446),
.B(n_402),
.Y(n_487)
);

XOR2xp5_ASAP7_75t_L g514 ( 
.A(n_487),
.B(n_497),
.Y(n_514)
);

INVx1_ASAP7_75t_L g524 ( 
.A(n_488),
.Y(n_524)
);

OAI22xp5_ASAP7_75t_SL g519 ( 
.A1(n_490),
.A2(n_492),
.B1(n_511),
.B2(n_465),
.Y(n_519)
);

OAI22xp5_ASAP7_75t_SL g491 ( 
.A1(n_453),
.A2(n_431),
.B1(n_420),
.B2(n_432),
.Y(n_491)
);

AOI22xp5_ASAP7_75t_L g492 ( 
.A1(n_443),
.A2(n_412),
.B1(n_425),
.B2(n_441),
.Y(n_492)
);

OAI22xp5_ASAP7_75t_L g493 ( 
.A1(n_462),
.A2(n_412),
.B1(n_418),
.B2(n_424),
.Y(n_493)
);

CKINVDCx16_ASAP7_75t_R g496 ( 
.A(n_475),
.Y(n_496)
);

NAND2xp5_ASAP7_75t_L g539 ( 
.A(n_496),
.B(n_485),
.Y(n_539)
);

XOR2xp5_ASAP7_75t_L g497 ( 
.A(n_449),
.B(n_416),
.Y(n_497)
);

XOR2xp5_ASAP7_75t_L g498 ( 
.A(n_459),
.B(n_439),
.Y(n_498)
);

MAJIxp5_ASAP7_75t_L g515 ( 
.A(n_498),
.B(n_500),
.C(n_512),
.Y(n_515)
);

OAI22xp5_ASAP7_75t_SL g499 ( 
.A1(n_476),
.A2(n_430),
.B1(n_434),
.B2(n_408),
.Y(n_499)
);

MAJIxp5_ASAP7_75t_L g500 ( 
.A(n_470),
.B(n_438),
.C(n_430),
.Y(n_500)
);

AO21x1_ASAP7_75t_L g505 ( 
.A1(n_476),
.A2(n_438),
.B(n_411),
.Y(n_505)
);

INVxp67_ASAP7_75t_L g520 ( 
.A(n_505),
.Y(n_520)
);

NAND2xp5_ASAP7_75t_SL g510 ( 
.A(n_447),
.B(n_434),
.Y(n_510)
);

CKINVDCx14_ASAP7_75t_R g536 ( 
.A(n_510),
.Y(n_536)
);

AOI22xp5_ASAP7_75t_L g511 ( 
.A1(n_448),
.A2(n_425),
.B1(n_411),
.B2(n_408),
.Y(n_511)
);

MAJIxp5_ASAP7_75t_L g512 ( 
.A(n_464),
.B(n_455),
.C(n_451),
.Y(n_512)
);

INVx1_ASAP7_75t_L g513 ( 
.A(n_502),
.Y(n_513)
);

INVx1_ASAP7_75t_L g545 ( 
.A(n_513),
.Y(n_545)
);

MAJIxp5_ASAP7_75t_L g516 ( 
.A(n_487),
.B(n_469),
.C(n_468),
.Y(n_516)
);

MAJIxp5_ASAP7_75t_L g554 ( 
.A(n_516),
.B(n_532),
.C(n_535),
.Y(n_554)
);

INVx1_ASAP7_75t_L g517 ( 
.A(n_502),
.Y(n_517)
);

INVx1_ASAP7_75t_L g564 ( 
.A(n_517),
.Y(n_564)
);

CKINVDCx20_ASAP7_75t_R g518 ( 
.A(n_504),
.Y(n_518)
);

NAND2xp5_ASAP7_75t_SL g546 ( 
.A(n_518),
.B(n_525),
.Y(n_546)
);

AOI22xp5_ASAP7_75t_L g544 ( 
.A1(n_519),
.A2(n_499),
.B1(n_491),
.B2(n_481),
.Y(n_544)
);

XOR2xp5_ASAP7_75t_L g558 ( 
.A(n_521),
.B(n_541),
.Y(n_558)
);

NOR2xp33_ASAP7_75t_SL g525 ( 
.A(n_494),
.B(n_460),
.Y(n_525)
);

CKINVDCx20_ASAP7_75t_R g526 ( 
.A(n_504),
.Y(n_526)
);

NOR2xp33_ASAP7_75t_SL g559 ( 
.A(n_526),
.B(n_533),
.Y(n_559)
);

INVx1_ASAP7_75t_L g527 ( 
.A(n_506),
.Y(n_527)
);

INVx1_ASAP7_75t_L g565 ( 
.A(n_527),
.Y(n_565)
);

INVx1_ASAP7_75t_L g528 ( 
.A(n_506),
.Y(n_528)
);

INVx1_ASAP7_75t_SL g563 ( 
.A(n_528),
.Y(n_563)
);

INVx1_ASAP7_75t_L g529 ( 
.A(n_495),
.Y(n_529)
);

NAND2xp5_ASAP7_75t_L g547 ( 
.A(n_529),
.B(n_530),
.Y(n_547)
);

INVx1_ASAP7_75t_L g530 ( 
.A(n_495),
.Y(n_530)
);

OAI21xp5_ASAP7_75t_L g551 ( 
.A1(n_531),
.A2(n_537),
.B(n_501),
.Y(n_551)
);

MAJIxp5_ASAP7_75t_L g532 ( 
.A(n_484),
.B(n_454),
.C(n_477),
.Y(n_532)
);

NOR2xp67_ASAP7_75t_SL g533 ( 
.A(n_500),
.B(n_448),
.Y(n_533)
);

CKINVDCx20_ASAP7_75t_R g534 ( 
.A(n_486),
.Y(n_534)
);

NAND2xp5_ASAP7_75t_L g549 ( 
.A(n_534),
.B(n_539),
.Y(n_549)
);

MAJIxp5_ASAP7_75t_L g535 ( 
.A(n_484),
.B(n_454),
.C(n_448),
.Y(n_535)
);

AOI21xp5_ASAP7_75t_L g537 ( 
.A1(n_501),
.A2(n_471),
.B(n_462),
.Y(n_537)
);

MAJIxp5_ASAP7_75t_L g538 ( 
.A(n_512),
.B(n_478),
.C(n_466),
.Y(n_538)
);

MAJIxp5_ASAP7_75t_L g557 ( 
.A(n_538),
.B(n_498),
.C(n_497),
.Y(n_557)
);

INVx1_ASAP7_75t_L g540 ( 
.A(n_508),
.Y(n_540)
);

HB1xp67_ASAP7_75t_L g553 ( 
.A(n_540),
.Y(n_553)
);

XNOR2xp5_ASAP7_75t_L g541 ( 
.A(n_479),
.B(n_474),
.Y(n_541)
);

XNOR2xp5_ASAP7_75t_L g542 ( 
.A(n_482),
.B(n_452),
.Y(n_542)
);

XOR2xp5_ASAP7_75t_L g566 ( 
.A(n_542),
.B(n_514),
.Y(n_566)
);

INVx1_ASAP7_75t_L g543 ( 
.A(n_508),
.Y(n_543)
);

NAND2xp5_ASAP7_75t_L g562 ( 
.A(n_543),
.B(n_503),
.Y(n_562)
);

OAI22xp5_ASAP7_75t_SL g571 ( 
.A1(n_544),
.A2(n_522),
.B1(n_517),
.B2(n_509),
.Y(n_571)
);

OAI21xp33_ASAP7_75t_L g548 ( 
.A1(n_524),
.A2(n_485),
.B(n_489),
.Y(n_548)
);

INVx1_ASAP7_75t_L g572 ( 
.A(n_548),
.Y(n_572)
);

CKINVDCx16_ASAP7_75t_R g550 ( 
.A(n_539),
.Y(n_550)
);

NAND2xp5_ASAP7_75t_L g589 ( 
.A(n_550),
.B(n_555),
.Y(n_589)
);

XNOR2xp5_ASAP7_75t_L g576 ( 
.A(n_551),
.B(n_557),
.Y(n_576)
);

NOR3xp33_ASAP7_75t_SL g552 ( 
.A(n_529),
.B(n_530),
.C(n_536),
.Y(n_552)
);

OAI22xp5_ASAP7_75t_L g574 ( 
.A1(n_552),
.A2(n_520),
.B1(n_505),
.B2(n_507),
.Y(n_574)
);

CKINVDCx16_ASAP7_75t_R g555 ( 
.A(n_537),
.Y(n_555)
);

NAND2xp5_ASAP7_75t_SL g556 ( 
.A(n_513),
.B(n_496),
.Y(n_556)
);

INVx1_ASAP7_75t_L g581 ( 
.A(n_556),
.Y(n_581)
);

OAI22xp5_ASAP7_75t_L g560 ( 
.A1(n_522),
.A2(n_490),
.B1(n_511),
.B2(n_505),
.Y(n_560)
);

INVx1_ASAP7_75t_L g586 ( 
.A(n_560),
.Y(n_586)
);

FAx1_ASAP7_75t_SL g561 ( 
.A(n_535),
.B(n_482),
.CI(n_483),
.CON(n_561),
.SN(n_561)
);

NOR2xp33_ASAP7_75t_L g573 ( 
.A(n_561),
.B(n_516),
.Y(n_573)
);

CKINVDCx20_ASAP7_75t_R g579 ( 
.A(n_562),
.Y(n_579)
);

XOR2xp5_ASAP7_75t_L g585 ( 
.A(n_566),
.B(n_521),
.Y(n_585)
);

NAND2xp5_ASAP7_75t_L g567 ( 
.A(n_527),
.B(n_489),
.Y(n_567)
);

INVx1_ASAP7_75t_L g582 ( 
.A(n_567),
.Y(n_582)
);

NAND2xp5_ASAP7_75t_L g568 ( 
.A(n_528),
.B(n_456),
.Y(n_568)
);

INVx1_ASAP7_75t_L g584 ( 
.A(n_568),
.Y(n_584)
);

HB1xp67_ASAP7_75t_L g569 ( 
.A(n_553),
.Y(n_569)
);

INVx1_ASAP7_75t_L g594 ( 
.A(n_569),
.Y(n_594)
);

MAJIxp5_ASAP7_75t_L g570 ( 
.A(n_554),
.B(n_538),
.C(n_515),
.Y(n_570)
);

NAND2xp5_ASAP7_75t_L g606 ( 
.A(n_570),
.B(n_575),
.Y(n_606)
);

AOI22xp5_ASAP7_75t_L g592 ( 
.A1(n_571),
.A2(n_588),
.B1(n_560),
.B2(n_509),
.Y(n_592)
);

INVxp67_ASAP7_75t_L g602 ( 
.A(n_573),
.Y(n_602)
);

INVx1_ASAP7_75t_L g597 ( 
.A(n_574),
.Y(n_597)
);

MAJIxp5_ASAP7_75t_L g575 ( 
.A(n_554),
.B(n_515),
.C(n_557),
.Y(n_575)
);

NOR2xp33_ASAP7_75t_L g577 ( 
.A(n_559),
.B(n_523),
.Y(n_577)
);

INVx1_ASAP7_75t_L g599 ( 
.A(n_577),
.Y(n_599)
);

XNOR2xp5_ASAP7_75t_L g578 ( 
.A(n_558),
.B(n_532),
.Y(n_578)
);

NOR2xp67_ASAP7_75t_SL g590 ( 
.A(n_578),
.B(n_583),
.Y(n_590)
);

NOR2xp33_ASAP7_75t_L g580 ( 
.A(n_559),
.B(n_541),
.Y(n_580)
);

CKINVDCx20_ASAP7_75t_R g593 ( 
.A(n_580),
.Y(n_593)
);

MAJIxp5_ASAP7_75t_L g583 ( 
.A(n_566),
.B(n_542),
.C(n_514),
.Y(n_583)
);

XNOR2xp5_ASAP7_75t_L g604 ( 
.A(n_585),
.B(n_549),
.Y(n_604)
);

MAJIxp5_ASAP7_75t_L g587 ( 
.A(n_558),
.B(n_507),
.C(n_519),
.Y(n_587)
);

MAJIxp5_ASAP7_75t_L g598 ( 
.A(n_587),
.B(n_551),
.C(n_567),
.Y(n_598)
);

OAI22xp5_ASAP7_75t_SL g588 ( 
.A1(n_544),
.A2(n_555),
.B1(n_550),
.B2(n_520),
.Y(n_588)
);

AND2x2_ASAP7_75t_L g591 ( 
.A(n_576),
.B(n_549),
.Y(n_591)
);

INVxp67_ASAP7_75t_L g618 ( 
.A(n_591),
.Y(n_618)
);

INVxp67_ASAP7_75t_L g620 ( 
.A(n_592),
.Y(n_620)
);

NOR2xp33_ASAP7_75t_L g595 ( 
.A(n_572),
.B(n_546),
.Y(n_595)
);

NAND2xp5_ASAP7_75t_L g611 ( 
.A(n_595),
.B(n_600),
.Y(n_611)
);

AOI22xp5_ASAP7_75t_L g596 ( 
.A1(n_586),
.A2(n_588),
.B1(n_571),
.B2(n_584),
.Y(n_596)
);

OAI22xp5_ASAP7_75t_SL g608 ( 
.A1(n_596),
.A2(n_587),
.B1(n_589),
.B2(n_531),
.Y(n_608)
);

NAND2xp5_ASAP7_75t_SL g610 ( 
.A(n_598),
.B(n_604),
.Y(n_610)
);

OAI22xp5_ASAP7_75t_L g600 ( 
.A1(n_586),
.A2(n_579),
.B1(n_582),
.B2(n_562),
.Y(n_600)
);

MAJIxp5_ASAP7_75t_L g601 ( 
.A(n_570),
.B(n_563),
.C(n_547),
.Y(n_601)
);

NAND2xp5_ASAP7_75t_L g619 ( 
.A(n_601),
.B(n_603),
.Y(n_619)
);

MAJIxp5_ASAP7_75t_L g603 ( 
.A(n_575),
.B(n_563),
.C(n_547),
.Y(n_603)
);

MAJIxp5_ASAP7_75t_L g605 ( 
.A(n_576),
.B(n_564),
.C(n_545),
.Y(n_605)
);

MAJIxp5_ASAP7_75t_L g614 ( 
.A(n_605),
.B(n_565),
.C(n_578),
.Y(n_614)
);

OAI22xp5_ASAP7_75t_SL g607 ( 
.A1(n_581),
.A2(n_564),
.B1(n_545),
.B2(n_556),
.Y(n_607)
);

AOI22xp5_ASAP7_75t_L g616 ( 
.A1(n_607),
.A2(n_493),
.B1(n_458),
.B2(n_450),
.Y(n_616)
);

INVx1_ASAP7_75t_L g626 ( 
.A(n_608),
.Y(n_626)
);

OAI21xp5_ASAP7_75t_L g609 ( 
.A1(n_597),
.A2(n_589),
.B(n_568),
.Y(n_609)
);

AOI21xp5_ASAP7_75t_L g623 ( 
.A1(n_609),
.A2(n_598),
.B(n_601),
.Y(n_623)
);

OR2x2_ASAP7_75t_L g612 ( 
.A(n_605),
.B(n_552),
.Y(n_612)
);

A2O1A1Ixp33_ASAP7_75t_L g625 ( 
.A1(n_612),
.A2(n_603),
.B(n_606),
.C(n_604),
.Y(n_625)
);

OAI22xp5_ASAP7_75t_SL g613 ( 
.A1(n_599),
.A2(n_565),
.B1(n_492),
.B2(n_561),
.Y(n_613)
);

OR2x2_ASAP7_75t_L g631 ( 
.A(n_613),
.B(n_614),
.Y(n_631)
);

NOR2xp33_ASAP7_75t_SL g615 ( 
.A(n_602),
.B(n_583),
.Y(n_615)
);

NOR2xp33_ASAP7_75t_L g622 ( 
.A(n_615),
.B(n_617),
.Y(n_622)
);

NAND2xp5_ASAP7_75t_SL g630 ( 
.A(n_616),
.B(n_621),
.Y(n_630)
);

NOR2xp33_ASAP7_75t_SL g617 ( 
.A(n_602),
.B(n_472),
.Y(n_617)
);

AOI22xp5_ASAP7_75t_L g621 ( 
.A1(n_591),
.A2(n_561),
.B1(n_585),
.B2(n_442),
.Y(n_621)
);

AOI21xp5_ASAP7_75t_L g633 ( 
.A1(n_623),
.A2(n_625),
.B(n_628),
.Y(n_633)
);

INVxp67_ASAP7_75t_L g624 ( 
.A(n_610),
.Y(n_624)
);

NAND2xp5_ASAP7_75t_L g634 ( 
.A(n_624),
.B(n_627),
.Y(n_634)
);

BUFx2_ASAP7_75t_L g627 ( 
.A(n_619),
.Y(n_627)
);

OAI21xp5_ASAP7_75t_SL g628 ( 
.A1(n_612),
.A2(n_590),
.B(n_593),
.Y(n_628)
);

OAI21xp5_ASAP7_75t_SL g629 ( 
.A1(n_611),
.A2(n_596),
.B(n_594),
.Y(n_629)
);

NAND2xp5_ASAP7_75t_L g635 ( 
.A(n_629),
.B(n_618),
.Y(n_635)
);

OAI21xp5_ASAP7_75t_SL g632 ( 
.A1(n_626),
.A2(n_618),
.B(n_614),
.Y(n_632)
);

MAJIxp5_ASAP7_75t_L g641 ( 
.A(n_632),
.B(n_630),
.C(n_592),
.Y(n_641)
);

AO21x1_ASAP7_75t_L g642 ( 
.A1(n_635),
.A2(n_637),
.B(n_638),
.Y(n_642)
);

NAND2xp5_ASAP7_75t_L g636 ( 
.A(n_622),
.B(n_620),
.Y(n_636)
);

INVxp67_ASAP7_75t_SL g639 ( 
.A(n_636),
.Y(n_639)
);

NOR2xp33_ASAP7_75t_SL g637 ( 
.A(n_622),
.B(n_609),
.Y(n_637)
);

NAND2xp5_ASAP7_75t_L g638 ( 
.A(n_631),
.B(n_620),
.Y(n_638)
);

OAI31xp33_ASAP7_75t_L g640 ( 
.A1(n_633),
.A2(n_630),
.A3(n_621),
.B(n_616),
.Y(n_640)
);

OAI21xp5_ASAP7_75t_L g644 ( 
.A1(n_640),
.A2(n_639),
.B(n_642),
.Y(n_644)
);

AOI22xp5_ASAP7_75t_L g643 ( 
.A1(n_641),
.A2(n_634),
.B1(n_633),
.B2(n_480),
.Y(n_643)
);

NAND3xp33_ASAP7_75t_L g645 ( 
.A(n_643),
.B(n_644),
.C(n_461),
.Y(n_645)
);

OR2x2_ASAP7_75t_L g646 ( 
.A(n_645),
.B(n_444),
.Y(n_646)
);

NAND2xp5_ASAP7_75t_SL g647 ( 
.A(n_646),
.B(n_428),
.Y(n_647)
);

AND2x2_ASAP7_75t_L g648 ( 
.A(n_647),
.B(n_473),
.Y(n_648)
);


endmodule