module fake_jpeg_3551_n_449 (n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_449);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_449;

wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_385;
wire n_228;
wire n_134;
wire n_428;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_377;
wire n_291;
wire n_236;
wire n_15;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_17;
wire n_431;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_415;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_13;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_429;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_305;
wire n_161;
wire n_441;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_382;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_14;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_389;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_384;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_433;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_413;
wire n_275;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_379;
wire n_114;
wire n_444;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_183;
wire n_409;
wire n_249;
wire n_412;
wire n_217;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_391;
wire n_209;
wire n_22;
wire n_138;
wire n_402;
wire n_438;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

BUFx5_ASAP7_75t_L g13 ( 
.A(n_7),
.Y(n_13)
);

BUFx12f_ASAP7_75t_L g14 ( 
.A(n_5),
.Y(n_14)
);

INVx1_ASAP7_75t_L g15 ( 
.A(n_7),
.Y(n_15)
);

BUFx6f_ASAP7_75t_L g16 ( 
.A(n_12),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_9),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_1),
.Y(n_18)
);

INVx1_ASAP7_75t_SL g19 ( 
.A(n_4),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_5),
.Y(n_20)
);

INVx3_ASAP7_75t_L g21 ( 
.A(n_8),
.Y(n_21)
);

BUFx12f_ASAP7_75t_L g22 ( 
.A(n_11),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_4),
.Y(n_23)
);

BUFx12f_ASAP7_75t_L g24 ( 
.A(n_12),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_12),
.Y(n_25)
);

BUFx24_ASAP7_75t_L g26 ( 
.A(n_7),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_3),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_6),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_6),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_7),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_12),
.Y(n_31)
);

BUFx12_ASAP7_75t_L g32 ( 
.A(n_3),
.Y(n_32)
);

INVxp33_ASAP7_75t_L g33 ( 
.A(n_2),
.Y(n_33)
);

INVx6_ASAP7_75t_L g34 ( 
.A(n_4),
.Y(n_34)
);

BUFx3_ASAP7_75t_L g35 ( 
.A(n_3),
.Y(n_35)
);

INVx6_ASAP7_75t_L g36 ( 
.A(n_0),
.Y(n_36)
);

INVx11_ASAP7_75t_L g37 ( 
.A(n_2),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_9),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_2),
.Y(n_39)
);

BUFx12f_ASAP7_75t_L g40 ( 
.A(n_0),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_1),
.Y(n_41)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_3),
.Y(n_42)
);

BUFx5_ASAP7_75t_L g43 ( 
.A(n_5),
.Y(n_43)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_8),
.Y(n_44)
);

BUFx12f_ASAP7_75t_L g45 ( 
.A(n_32),
.Y(n_45)
);

INVx1_ASAP7_75t_SL g131 ( 
.A(n_45),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g46 ( 
.A(n_21),
.B(n_0),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_L g115 ( 
.A(n_46),
.B(n_49),
.Y(n_115)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_34),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_47),
.B(n_59),
.Y(n_101)
);

BUFx5_ASAP7_75t_L g48 ( 
.A(n_26),
.Y(n_48)
);

BUFx5_ASAP7_75t_L g109 ( 
.A(n_48),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_L g49 ( 
.A(n_21),
.B(n_0),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_16),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g103 ( 
.A(n_50),
.Y(n_103)
);

BUFx3_ASAP7_75t_L g51 ( 
.A(n_35),
.Y(n_51)
);

BUFx3_ASAP7_75t_L g128 ( 
.A(n_51),
.Y(n_128)
);

INVx6_ASAP7_75t_L g52 ( 
.A(n_16),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g105 ( 
.A(n_52),
.Y(n_105)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_16),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g142 ( 
.A(n_53),
.Y(n_142)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_23),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g149 ( 
.A(n_54),
.Y(n_149)
);

BUFx10_ASAP7_75t_L g55 ( 
.A(n_24),
.Y(n_55)
);

INVx2_ASAP7_75t_SL g125 ( 
.A(n_55),
.Y(n_125)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_23),
.Y(n_56)
);

INVx6_ASAP7_75t_L g132 ( 
.A(n_56),
.Y(n_132)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_23),
.Y(n_57)
);

INVx8_ASAP7_75t_L g117 ( 
.A(n_57),
.Y(n_117)
);

INVx4_ASAP7_75t_L g58 ( 
.A(n_40),
.Y(n_58)
);

INVx3_ASAP7_75t_L g136 ( 
.A(n_58),
.Y(n_136)
);

CKINVDCx20_ASAP7_75t_R g59 ( 
.A(n_34),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_30),
.Y(n_60)
);

INVx2_ASAP7_75t_L g108 ( 
.A(n_60),
.Y(n_108)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_30),
.Y(n_61)
);

INVx2_ASAP7_75t_L g112 ( 
.A(n_61),
.Y(n_112)
);

AND2x2_ASAP7_75t_SL g62 ( 
.A(n_40),
.B(n_0),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g118 ( 
.A(n_62),
.B(n_69),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_L g63 ( 
.A(n_33),
.B(n_11),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_L g135 ( 
.A(n_63),
.B(n_65),
.Y(n_135)
);

INVx11_ASAP7_75t_L g64 ( 
.A(n_40),
.Y(n_64)
);

INVx4_ASAP7_75t_L g98 ( 
.A(n_64),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g65 ( 
.A(n_36),
.B(n_1),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_15),
.B(n_1),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_SL g133 ( 
.A(n_66),
.B(n_70),
.Y(n_133)
);

BUFx12f_ASAP7_75t_L g67 ( 
.A(n_32),
.Y(n_67)
);

INVx4_ASAP7_75t_L g107 ( 
.A(n_67),
.Y(n_107)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_30),
.Y(n_68)
);

INVx2_ASAP7_75t_L g114 ( 
.A(n_68),
.Y(n_114)
);

CKINVDCx20_ASAP7_75t_R g69 ( 
.A(n_34),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_15),
.B(n_2),
.Y(n_70)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_17),
.Y(n_71)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_71),
.Y(n_102)
);

BUFx6f_ASAP7_75t_L g72 ( 
.A(n_41),
.Y(n_72)
);

INVx2_ASAP7_75t_L g124 ( 
.A(n_72),
.Y(n_124)
);

NAND2xp33_ASAP7_75t_SL g73 ( 
.A(n_19),
.B(n_4),
.Y(n_73)
);

NAND3xp33_ASAP7_75t_L g111 ( 
.A(n_73),
.B(n_27),
.C(n_39),
.Y(n_111)
);

BUFx10_ASAP7_75t_L g74 ( 
.A(n_24),
.Y(n_74)
);

BUFx2_ASAP7_75t_SL g140 ( 
.A(n_74),
.Y(n_140)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_17),
.Y(n_75)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_75),
.Y(n_126)
);

CKINVDCx16_ASAP7_75t_R g76 ( 
.A(n_26),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g120 ( 
.A(n_76),
.B(n_77),
.Y(n_120)
);

CKINVDCx20_ASAP7_75t_R g77 ( 
.A(n_36),
.Y(n_77)
);

BUFx6f_ASAP7_75t_L g78 ( 
.A(n_41),
.Y(n_78)
);

INVx2_ASAP7_75t_L g127 ( 
.A(n_78),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_18),
.B(n_5),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g137 ( 
.A(n_79),
.B(n_85),
.Y(n_137)
);

BUFx6f_ASAP7_75t_L g80 ( 
.A(n_41),
.Y(n_80)
);

INVx4_ASAP7_75t_L g119 ( 
.A(n_80),
.Y(n_119)
);

INVx11_ASAP7_75t_L g81 ( 
.A(n_40),
.Y(n_81)
);

INVx4_ASAP7_75t_L g121 ( 
.A(n_81),
.Y(n_121)
);

INVx11_ASAP7_75t_L g82 ( 
.A(n_40),
.Y(n_82)
);

INVx2_ASAP7_75t_L g104 ( 
.A(n_82),
.Y(n_104)
);

INVx11_ASAP7_75t_L g83 ( 
.A(n_24),
.Y(n_83)
);

INVx2_ASAP7_75t_L g123 ( 
.A(n_83),
.Y(n_123)
);

BUFx5_ASAP7_75t_L g84 ( 
.A(n_26),
.Y(n_84)
);

INVx2_ASAP7_75t_L g145 ( 
.A(n_84),
.Y(n_145)
);

CKINVDCx20_ASAP7_75t_R g85 ( 
.A(n_36),
.Y(n_85)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_18),
.Y(n_86)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_86),
.Y(n_138)
);

BUFx3_ASAP7_75t_L g87 ( 
.A(n_35),
.Y(n_87)
);

INVx2_ASAP7_75t_L g146 ( 
.A(n_87),
.Y(n_146)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_20),
.Y(n_88)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_88),
.Y(n_141)
);

INVx11_ASAP7_75t_L g89 ( 
.A(n_24),
.Y(n_89)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_89),
.Y(n_150)
);

INVx2_ASAP7_75t_L g90 ( 
.A(n_24),
.Y(n_90)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_90),
.Y(n_152)
);

CKINVDCx20_ASAP7_75t_R g91 ( 
.A(n_32),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g147 ( 
.A(n_91),
.B(n_96),
.Y(n_147)
);

INVx8_ASAP7_75t_L g92 ( 
.A(n_14),
.Y(n_92)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_92),
.Y(n_153)
);

INVx3_ASAP7_75t_L g93 ( 
.A(n_14),
.Y(n_93)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_93),
.Y(n_154)
);

INVx2_ASAP7_75t_L g94 ( 
.A(n_14),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_SL g139 ( 
.A(n_94),
.B(n_97),
.Y(n_139)
);

BUFx2_ASAP7_75t_L g95 ( 
.A(n_35),
.Y(n_95)
);

CKINVDCx20_ASAP7_75t_R g116 ( 
.A(n_95),
.Y(n_116)
);

INVx8_ASAP7_75t_L g96 ( 
.A(n_14),
.Y(n_96)
);

INVx3_ASAP7_75t_L g97 ( 
.A(n_22),
.Y(n_97)
);

AOI22xp5_ASAP7_75t_L g99 ( 
.A1(n_65),
.A2(n_19),
.B1(n_42),
.B2(n_31),
.Y(n_99)
);

OAI22xp5_ASAP7_75t_SL g190 ( 
.A1(n_99),
.A2(n_129),
.B1(n_143),
.B2(n_13),
.Y(n_190)
);

OAI22xp5_ASAP7_75t_L g100 ( 
.A1(n_46),
.A2(n_49),
.B1(n_52),
.B2(n_72),
.Y(n_100)
);

OAI22xp5_ASAP7_75t_L g166 ( 
.A1(n_100),
.A2(n_106),
.B1(n_113),
.B2(n_134),
.Y(n_166)
);

AOI22xp33_ASAP7_75t_L g106 ( 
.A1(n_50),
.A2(n_27),
.B1(n_39),
.B2(n_38),
.Y(n_106)
);

AOI22xp33_ASAP7_75t_SL g110 ( 
.A1(n_64),
.A2(n_19),
.B1(n_37),
.B2(n_22),
.Y(n_110)
);

OA22x2_ASAP7_75t_L g195 ( 
.A1(n_110),
.A2(n_122),
.B1(n_130),
.B2(n_144),
.Y(n_195)
);

AND2x2_ASAP7_75t_L g159 ( 
.A(n_111),
.B(n_62),
.Y(n_159)
);

AOI22xp33_ASAP7_75t_L g113 ( 
.A1(n_53),
.A2(n_28),
.B1(n_29),
.B2(n_38),
.Y(n_113)
);

AOI22xp33_ASAP7_75t_SL g122 ( 
.A1(n_81),
.A2(n_37),
.B1(n_22),
.B2(n_44),
.Y(n_122)
);

AOI22xp5_ASAP7_75t_L g129 ( 
.A1(n_54),
.A2(n_44),
.B1(n_42),
.B2(n_31),
.Y(n_129)
);

AOI22xp5_ASAP7_75t_SL g130 ( 
.A1(n_94),
.A2(n_97),
.B1(n_93),
.B2(n_95),
.Y(n_130)
);

OAI22xp33_ASAP7_75t_L g134 ( 
.A1(n_56),
.A2(n_37),
.B1(n_25),
.B2(n_20),
.Y(n_134)
);

AOI22xp33_ASAP7_75t_L g143 ( 
.A1(n_57),
.A2(n_29),
.B1(n_28),
.B2(n_25),
.Y(n_143)
);

AOI22xp33_ASAP7_75t_SL g144 ( 
.A1(n_82),
.A2(n_22),
.B1(n_26),
.B2(n_43),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_SL g148 ( 
.A(n_73),
.B(n_6),
.Y(n_148)
);

NOR2xp33_ASAP7_75t_SL g174 ( 
.A(n_148),
.B(n_151),
.Y(n_174)
);

NOR2xp33_ASAP7_75t_L g151 ( 
.A(n_45),
.B(n_6),
.Y(n_151)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_102),
.Y(n_155)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_155),
.Y(n_204)
);

BUFx6f_ASAP7_75t_L g156 ( 
.A(n_103),
.Y(n_156)
);

BUFx6f_ASAP7_75t_L g225 ( 
.A(n_156),
.Y(n_225)
);

BUFx6f_ASAP7_75t_L g157 ( 
.A(n_103),
.Y(n_157)
);

INVx6_ASAP7_75t_L g223 ( 
.A(n_157),
.Y(n_223)
);

CKINVDCx16_ASAP7_75t_R g158 ( 
.A(n_120),
.Y(n_158)
);

NOR2xp33_ASAP7_75t_L g209 ( 
.A(n_158),
.B(n_170),
.Y(n_209)
);

NOR2xp33_ASAP7_75t_SL g212 ( 
.A(n_159),
.B(n_168),
.Y(n_212)
);

INVx4_ASAP7_75t_L g160 ( 
.A(n_125),
.Y(n_160)
);

INVx4_ASAP7_75t_L g205 ( 
.A(n_160),
.Y(n_205)
);

NAND2xp5_ASAP7_75t_L g161 ( 
.A(n_115),
.B(n_62),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_L g230 ( 
.A(n_161),
.B(n_172),
.Y(n_230)
);

O2A1O1Ixp33_ASAP7_75t_L g162 ( 
.A1(n_118),
.A2(n_48),
.B(n_84),
.C(n_51),
.Y(n_162)
);

AOI21xp5_ASAP7_75t_L g206 ( 
.A1(n_162),
.A2(n_110),
.B(n_122),
.Y(n_206)
);

AO22x2_ASAP7_75t_L g163 ( 
.A1(n_146),
.A2(n_58),
.B1(n_90),
.B2(n_55),
.Y(n_163)
);

AND2x2_ASAP7_75t_L g214 ( 
.A(n_163),
.B(n_167),
.Y(n_214)
);

INVx2_ASAP7_75t_SL g164 ( 
.A(n_125),
.Y(n_164)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_164),
.Y(n_218)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_126),
.Y(n_165)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_165),
.Y(n_220)
);

AND2x2_ASAP7_75t_L g167 ( 
.A(n_139),
.B(n_99),
.Y(n_167)
);

NOR2xp33_ASAP7_75t_L g168 ( 
.A(n_133),
.B(n_87),
.Y(n_168)
);

AOI22xp33_ASAP7_75t_SL g169 ( 
.A1(n_116),
.A2(n_89),
.B1(n_83),
.B2(n_137),
.Y(n_169)
);

AOI22xp33_ASAP7_75t_SL g222 ( 
.A1(n_169),
.A2(n_179),
.B1(n_196),
.B2(n_197),
.Y(n_222)
);

NOR2xp33_ASAP7_75t_L g170 ( 
.A(n_138),
.B(n_96),
.Y(n_170)
);

NOR2xp33_ASAP7_75t_L g171 ( 
.A(n_141),
.B(n_101),
.Y(n_171)
);

NOR2xp33_ASAP7_75t_L g211 ( 
.A(n_171),
.B(n_173),
.Y(n_211)
);

NAND2xp5_ASAP7_75t_L g172 ( 
.A(n_135),
.B(n_78),
.Y(n_172)
);

NOR2xp33_ASAP7_75t_L g173 ( 
.A(n_147),
.B(n_92),
.Y(n_173)
);

INVxp33_ASAP7_75t_L g175 ( 
.A(n_130),
.Y(n_175)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_175),
.Y(n_224)
);

INVx2_ASAP7_75t_L g176 ( 
.A(n_108),
.Y(n_176)
);

INVx2_ASAP7_75t_L g201 ( 
.A(n_176),
.Y(n_201)
);

BUFx3_ASAP7_75t_L g177 ( 
.A(n_131),
.Y(n_177)
);

INVx3_ASAP7_75t_L g213 ( 
.A(n_177),
.Y(n_213)
);

NOR2xp33_ASAP7_75t_L g178 ( 
.A(n_154),
.B(n_45),
.Y(n_178)
);

NOR2xp33_ASAP7_75t_L g216 ( 
.A(n_178),
.B(n_183),
.Y(n_216)
);

AOI22xp33_ASAP7_75t_SL g179 ( 
.A1(n_131),
.A2(n_67),
.B1(n_68),
.B2(n_80),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_L g180 ( 
.A(n_152),
.B(n_61),
.Y(n_180)
);

MAJIxp5_ASAP7_75t_L g199 ( 
.A(n_180),
.B(n_181),
.C(n_182),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_L g181 ( 
.A(n_108),
.B(n_60),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_L g182 ( 
.A(n_112),
.B(n_67),
.Y(n_182)
);

CKINVDCx16_ASAP7_75t_R g183 ( 
.A(n_140),
.Y(n_183)
);

INVx2_ASAP7_75t_L g184 ( 
.A(n_112),
.Y(n_184)
);

INVx2_ASAP7_75t_L g208 ( 
.A(n_184),
.Y(n_208)
);

INVx8_ASAP7_75t_L g185 ( 
.A(n_142),
.Y(n_185)
);

INVx3_ASAP7_75t_L g229 ( 
.A(n_185),
.Y(n_229)
);

CKINVDCx20_ASAP7_75t_R g186 ( 
.A(n_105),
.Y(n_186)
);

NOR2xp33_ASAP7_75t_L g219 ( 
.A(n_186),
.B(n_189),
.Y(n_219)
);

INVx2_ASAP7_75t_L g187 ( 
.A(n_114),
.Y(n_187)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_187),
.Y(n_231)
);

NAND2xp5_ASAP7_75t_L g188 ( 
.A(n_114),
.B(n_8),
.Y(n_188)
);

MAJIxp5_ASAP7_75t_L g210 ( 
.A(n_188),
.B(n_194),
.C(n_150),
.Y(n_210)
);

BUFx12f_ASAP7_75t_L g189 ( 
.A(n_136),
.Y(n_189)
);

AOI22xp5_ASAP7_75t_L g202 ( 
.A1(n_190),
.A2(n_134),
.B1(n_127),
.B2(n_119),
.Y(n_202)
);

INVxp67_ASAP7_75t_L g191 ( 
.A(n_145),
.Y(n_191)
);

NOR2xp33_ASAP7_75t_L g227 ( 
.A(n_191),
.B(n_193),
.Y(n_227)
);

INVx5_ASAP7_75t_L g192 ( 
.A(n_128),
.Y(n_192)
);

CKINVDCx20_ASAP7_75t_R g228 ( 
.A(n_192),
.Y(n_228)
);

INVxp67_ASAP7_75t_L g193 ( 
.A(n_136),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_L g194 ( 
.A(n_124),
.B(n_8),
.Y(n_194)
);

AOI22xp33_ASAP7_75t_SL g196 ( 
.A1(n_144),
.A2(n_43),
.B1(n_13),
.B2(n_74),
.Y(n_196)
);

BUFx6f_ASAP7_75t_SL g197 ( 
.A(n_104),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_SL g198 ( 
.A(n_153),
.B(n_9),
.Y(n_198)
);

OR2x2_ASAP7_75t_L g215 ( 
.A(n_198),
.B(n_121),
.Y(n_215)
);

OAI22xp5_ASAP7_75t_SL g200 ( 
.A1(n_167),
.A2(n_129),
.B1(n_124),
.B2(n_127),
.Y(n_200)
);

AOI22xp5_ASAP7_75t_L g248 ( 
.A1(n_200),
.A2(n_176),
.B1(n_187),
.B2(n_184),
.Y(n_248)
);

OAI22xp5_ASAP7_75t_L g250 ( 
.A1(n_202),
.A2(n_207),
.B1(n_217),
.B2(n_221),
.Y(n_250)
);

FAx1_ASAP7_75t_SL g203 ( 
.A(n_161),
.B(n_74),
.CI(n_55),
.CON(n_203),
.SN(n_203)
);

NOR2xp33_ASAP7_75t_SL g242 ( 
.A(n_203),
.B(n_215),
.Y(n_242)
);

INVx1_ASAP7_75t_SL g253 ( 
.A(n_206),
.Y(n_253)
);

AOI22xp5_ASAP7_75t_L g207 ( 
.A1(n_166),
.A2(n_105),
.B1(n_119),
.B2(n_142),
.Y(n_207)
);

NAND2xp5_ASAP7_75t_L g237 ( 
.A(n_210),
.B(n_174),
.Y(n_237)
);

OAI22xp5_ASAP7_75t_L g217 ( 
.A1(n_172),
.A2(n_167),
.B1(n_188),
.B2(n_194),
.Y(n_217)
);

AOI22xp33_ASAP7_75t_L g221 ( 
.A1(n_175),
.A2(n_149),
.B1(n_123),
.B2(n_98),
.Y(n_221)
);

MAJIxp5_ASAP7_75t_L g226 ( 
.A(n_159),
.B(n_107),
.C(n_128),
.Y(n_226)
);

XNOR2xp5_ASAP7_75t_L g245 ( 
.A(n_226),
.B(n_163),
.Y(n_245)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_218),
.Y(n_232)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_232),
.Y(n_265)
);

CKINVDCx20_ASAP7_75t_R g233 ( 
.A(n_219),
.Y(n_233)
);

NOR2xp33_ASAP7_75t_L g271 ( 
.A(n_233),
.B(n_246),
.Y(n_271)
);

OAI22xp5_ASAP7_75t_L g234 ( 
.A1(n_207),
.A2(n_214),
.B1(n_217),
.B2(n_202),
.Y(n_234)
);

AOI22xp5_ASAP7_75t_SL g264 ( 
.A1(n_234),
.A2(n_258),
.B1(n_200),
.B2(n_228),
.Y(n_264)
);

INVx2_ASAP7_75t_SL g235 ( 
.A(n_218),
.Y(n_235)
);

INVx1_ASAP7_75t_SL g274 ( 
.A(n_235),
.Y(n_274)
);

AO21x1_ASAP7_75t_L g236 ( 
.A1(n_214),
.A2(n_159),
.B(n_162),
.Y(n_236)
);

OAI21xp5_ASAP7_75t_SL g270 ( 
.A1(n_236),
.A2(n_241),
.B(n_243),
.Y(n_270)
);

NAND2xp5_ASAP7_75t_SL g281 ( 
.A(n_237),
.B(n_244),
.Y(n_281)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_231),
.Y(n_238)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_238),
.Y(n_268)
);

INVx5_ASAP7_75t_L g239 ( 
.A(n_223),
.Y(n_239)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_239),
.Y(n_269)
);

AOI21xp5_ASAP7_75t_L g240 ( 
.A1(n_206),
.A2(n_195),
.B(n_164),
.Y(n_240)
);

AOI21xp5_ASAP7_75t_L g262 ( 
.A1(n_240),
.A2(n_222),
.B(n_203),
.Y(n_262)
);

OAI21xp5_ASAP7_75t_L g241 ( 
.A1(n_214),
.A2(n_190),
.B(n_182),
.Y(n_241)
);

AOI22xp5_ASAP7_75t_SL g243 ( 
.A1(n_212),
.A2(n_195),
.B1(n_192),
.B2(n_180),
.Y(n_243)
);

NOR2xp33_ASAP7_75t_SL g244 ( 
.A(n_230),
.B(n_181),
.Y(n_244)
);

MAJIxp5_ASAP7_75t_L g266 ( 
.A(n_245),
.B(n_251),
.C(n_255),
.Y(n_266)
);

OR2x2_ASAP7_75t_L g246 ( 
.A(n_212),
.B(n_195),
.Y(n_246)
);

CKINVDCx20_ASAP7_75t_R g247 ( 
.A(n_227),
.Y(n_247)
);

NAND2xp5_ASAP7_75t_L g263 ( 
.A(n_247),
.B(n_256),
.Y(n_263)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_248),
.Y(n_279)
);

AOI22xp33_ASAP7_75t_L g249 ( 
.A1(n_224),
.A2(n_163),
.B1(n_195),
.B2(n_149),
.Y(n_249)
);

INVxp67_ASAP7_75t_L g277 ( 
.A(n_249),
.Y(n_277)
);

XOR2xp5_ASAP7_75t_L g251 ( 
.A(n_230),
.B(n_163),
.Y(n_251)
);

INVx2_ASAP7_75t_L g252 ( 
.A(n_201),
.Y(n_252)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_252),
.Y(n_280)
);

BUFx5_ASAP7_75t_L g254 ( 
.A(n_201),
.Y(n_254)
);

CKINVDCx16_ASAP7_75t_R g276 ( 
.A(n_254),
.Y(n_276)
);

XNOR2xp5_ASAP7_75t_SL g255 ( 
.A(n_210),
.B(n_109),
.Y(n_255)
);

NAND2xp5_ASAP7_75t_L g256 ( 
.A(n_199),
.B(n_191),
.Y(n_256)
);

HB1xp67_ASAP7_75t_L g257 ( 
.A(n_205),
.Y(n_257)
);

CKINVDCx20_ASAP7_75t_R g267 ( 
.A(n_257),
.Y(n_267)
);

OAI22xp5_ASAP7_75t_SL g258 ( 
.A1(n_224),
.A2(n_132),
.B1(n_117),
.B2(n_157),
.Y(n_258)
);

CKINVDCx20_ASAP7_75t_R g259 ( 
.A(n_211),
.Y(n_259)
);

NAND2xp5_ASAP7_75t_L g275 ( 
.A(n_259),
.B(n_209),
.Y(n_275)
);

NAND2xp5_ASAP7_75t_L g260 ( 
.A(n_256),
.B(n_199),
.Y(n_260)
);

NAND2xp5_ASAP7_75t_L g291 ( 
.A(n_260),
.B(n_261),
.Y(n_291)
);

NAND2xp5_ASAP7_75t_L g261 ( 
.A(n_244),
.B(n_203),
.Y(n_261)
);

OAI21xp5_ASAP7_75t_L g287 ( 
.A1(n_262),
.A2(n_273),
.B(n_240),
.Y(n_287)
);

OAI22xp5_ASAP7_75t_SL g302 ( 
.A1(n_264),
.A2(n_235),
.B1(n_248),
.B2(n_232),
.Y(n_302)
);

MAJIxp5_ASAP7_75t_L g272 ( 
.A(n_255),
.B(n_226),
.C(n_204),
.Y(n_272)
);

MAJIxp5_ASAP7_75t_L g289 ( 
.A(n_272),
.B(n_245),
.C(n_246),
.Y(n_289)
);

AOI21xp5_ASAP7_75t_L g273 ( 
.A1(n_253),
.A2(n_228),
.B(n_213),
.Y(n_273)
);

CKINVDCx14_ASAP7_75t_R g300 ( 
.A(n_275),
.Y(n_300)
);

CKINVDCx20_ASAP7_75t_R g278 ( 
.A(n_239),
.Y(n_278)
);

INVx11_ASAP7_75t_L g296 ( 
.A(n_278),
.Y(n_296)
);

CKINVDCx16_ASAP7_75t_R g282 ( 
.A(n_236),
.Y(n_282)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_282),
.Y(n_293)
);

OAI22xp5_ASAP7_75t_SL g283 ( 
.A1(n_253),
.A2(n_215),
.B1(n_132),
.B2(n_204),
.Y(n_283)
);

NAND2xp5_ASAP7_75t_L g298 ( 
.A(n_283),
.B(n_284),
.Y(n_298)
);

FAx1_ASAP7_75t_SL g284 ( 
.A(n_241),
.B(n_216),
.CI(n_220),
.CON(n_284),
.SN(n_284)
);

NAND2xp5_ASAP7_75t_L g285 ( 
.A(n_251),
.B(n_220),
.Y(n_285)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_285),
.Y(n_304)
);

INVx2_ASAP7_75t_L g286 ( 
.A(n_265),
.Y(n_286)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_286),
.Y(n_322)
);

AOI21xp5_ASAP7_75t_L g313 ( 
.A1(n_287),
.A2(n_310),
.B(n_262),
.Y(n_313)
);

AOI22xp33_ASAP7_75t_SL g288 ( 
.A1(n_277),
.A2(n_258),
.B1(n_233),
.B2(n_250),
.Y(n_288)
);

AOI21xp33_ASAP7_75t_L g329 ( 
.A1(n_288),
.A2(n_270),
.B(n_279),
.Y(n_329)
);

MAJIxp5_ASAP7_75t_L g320 ( 
.A(n_289),
.B(n_292),
.C(n_294),
.Y(n_320)
);

INVx1_ASAP7_75t_SL g290 ( 
.A(n_273),
.Y(n_290)
);

NAND2xp5_ASAP7_75t_L g317 ( 
.A(n_290),
.B(n_301),
.Y(n_317)
);

XOR2xp5_ASAP7_75t_L g292 ( 
.A(n_266),
.B(n_237),
.Y(n_292)
);

MAJIxp5_ASAP7_75t_L g294 ( 
.A(n_266),
.B(n_247),
.C(n_243),
.Y(n_294)
);

AOI22xp5_ASAP7_75t_SL g295 ( 
.A1(n_282),
.A2(n_242),
.B1(n_234),
.B2(n_259),
.Y(n_295)
);

OAI22xp5_ASAP7_75t_SL g328 ( 
.A1(n_295),
.A2(n_261),
.B1(n_284),
.B2(n_270),
.Y(n_328)
);

XOR2xp5_ASAP7_75t_L g297 ( 
.A(n_266),
.B(n_242),
.Y(n_297)
);

MAJIxp5_ASAP7_75t_L g326 ( 
.A(n_297),
.B(n_299),
.C(n_305),
.Y(n_326)
);

XOR2xp5_ASAP7_75t_L g299 ( 
.A(n_260),
.B(n_236),
.Y(n_299)
);

INVx1_ASAP7_75t_SL g301 ( 
.A(n_273),
.Y(n_301)
);

AOI22xp5_ASAP7_75t_L g324 ( 
.A1(n_302),
.A2(n_283),
.B1(n_279),
.B2(n_285),
.Y(n_324)
);

CKINVDCx20_ASAP7_75t_R g303 ( 
.A(n_275),
.Y(n_303)
);

NAND2xp5_ASAP7_75t_L g319 ( 
.A(n_303),
.B(n_306),
.Y(n_319)
);

MAJIxp5_ASAP7_75t_L g305 ( 
.A(n_272),
.B(n_238),
.C(n_235),
.Y(n_305)
);

CKINVDCx20_ASAP7_75t_R g306 ( 
.A(n_267),
.Y(n_306)
);

MAJIxp5_ASAP7_75t_L g307 ( 
.A(n_272),
.B(n_231),
.C(n_107),
.Y(n_307)
);

MAJIxp5_ASAP7_75t_L g334 ( 
.A(n_307),
.B(n_268),
.C(n_280),
.Y(n_334)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_265),
.Y(n_308)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_308),
.Y(n_327)
);

NOR2xp33_ASAP7_75t_SL g309 ( 
.A(n_281),
.B(n_252),
.Y(n_309)
);

NOR2xp33_ASAP7_75t_L g315 ( 
.A(n_309),
.B(n_311),
.Y(n_315)
);

AOI21x1_ASAP7_75t_L g310 ( 
.A1(n_270),
.A2(n_262),
.B(n_271),
.Y(n_310)
);

NOR2xp33_ASAP7_75t_L g311 ( 
.A(n_263),
.B(n_205),
.Y(n_311)
);

XNOR2xp5_ASAP7_75t_L g312 ( 
.A(n_292),
.B(n_260),
.Y(n_312)
);

XOR2xp5_ASAP7_75t_L g357 ( 
.A(n_312),
.B(n_314),
.Y(n_357)
);

INVxp33_ASAP7_75t_L g344 ( 
.A(n_313),
.Y(n_344)
);

XOR2xp5_ASAP7_75t_L g314 ( 
.A(n_289),
.B(n_263),
.Y(n_314)
);

XOR2xp5_ASAP7_75t_L g316 ( 
.A(n_297),
.B(n_271),
.Y(n_316)
);

MAJIxp5_ASAP7_75t_L g338 ( 
.A(n_316),
.B(n_325),
.C(n_334),
.Y(n_338)
);

NOR2xp33_ASAP7_75t_L g318 ( 
.A(n_303),
.B(n_281),
.Y(n_318)
);

NOR2xp33_ASAP7_75t_SL g345 ( 
.A(n_318),
.B(n_323),
.Y(n_345)
);

NAND2xp5_ASAP7_75t_L g321 ( 
.A(n_300),
.B(n_267),
.Y(n_321)
);

NAND2xp5_ASAP7_75t_L g337 ( 
.A(n_321),
.B(n_330),
.Y(n_337)
);

NOR2xp33_ASAP7_75t_L g323 ( 
.A(n_291),
.B(n_269),
.Y(n_323)
);

OAI22xp5_ASAP7_75t_SL g349 ( 
.A1(n_324),
.A2(n_329),
.B1(n_293),
.B2(n_287),
.Y(n_349)
);

XOR2xp5_ASAP7_75t_L g325 ( 
.A(n_299),
.B(n_285),
.Y(n_325)
);

AOI22xp5_ASAP7_75t_L g354 ( 
.A1(n_328),
.A2(n_283),
.B1(n_284),
.B2(n_274),
.Y(n_354)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_286),
.Y(n_330)
);

NAND2xp5_ASAP7_75t_L g331 ( 
.A(n_306),
.B(n_304),
.Y(n_331)
);

NAND2xp5_ASAP7_75t_L g343 ( 
.A(n_331),
.B(n_332),
.Y(n_343)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_308),
.Y(n_332)
);

XNOR2xp5_ASAP7_75t_SL g333 ( 
.A(n_291),
.B(n_304),
.Y(n_333)
);

XNOR2xp5_ASAP7_75t_SL g340 ( 
.A(n_333),
.B(n_294),
.Y(n_340)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_302),
.Y(n_335)
);

NOR2xp33_ASAP7_75t_L g342 ( 
.A(n_335),
.B(n_298),
.Y(n_342)
);

MAJIxp5_ASAP7_75t_L g336 ( 
.A(n_305),
.B(n_261),
.C(n_284),
.Y(n_336)
);

MAJIxp5_ASAP7_75t_L g341 ( 
.A(n_336),
.B(n_307),
.C(n_295),
.Y(n_341)
);

NAND2xp5_ASAP7_75t_SL g339 ( 
.A(n_314),
.B(n_312),
.Y(n_339)
);

NOR2xp33_ASAP7_75t_SL g366 ( 
.A(n_339),
.B(n_351),
.Y(n_366)
);

XNOR2xp5_ASAP7_75t_SL g367 ( 
.A(n_340),
.B(n_317),
.Y(n_367)
);

NAND2xp5_ASAP7_75t_SL g363 ( 
.A(n_341),
.B(n_348),
.Y(n_363)
);

INVx1_ASAP7_75t_L g361 ( 
.A(n_342),
.Y(n_361)
);

MAJIxp5_ASAP7_75t_L g346 ( 
.A(n_326),
.B(n_310),
.C(n_298),
.Y(n_346)
);

MAJIxp5_ASAP7_75t_L g369 ( 
.A(n_346),
.B(n_347),
.C(n_353),
.Y(n_369)
);

MAJIxp5_ASAP7_75t_L g347 ( 
.A(n_326),
.B(n_320),
.C(n_334),
.Y(n_347)
);

CKINVDCx14_ASAP7_75t_R g348 ( 
.A(n_315),
.Y(n_348)
);

AOI22xp5_ASAP7_75t_L g370 ( 
.A1(n_349),
.A2(n_327),
.B1(n_322),
.B2(n_276),
.Y(n_370)
);

XNOR2xp5_ASAP7_75t_L g350 ( 
.A(n_316),
.B(n_293),
.Y(n_350)
);

XOR2xp5_ASAP7_75t_L g368 ( 
.A(n_350),
.B(n_358),
.Y(n_368)
);

NOR2xp33_ASAP7_75t_L g351 ( 
.A(n_336),
.B(n_328),
.Y(n_351)
);

CKINVDCx16_ASAP7_75t_R g352 ( 
.A(n_319),
.Y(n_352)
);

NAND2xp5_ASAP7_75t_SL g378 ( 
.A(n_352),
.B(n_355),
.Y(n_378)
);

MAJIxp5_ASAP7_75t_L g353 ( 
.A(n_320),
.B(n_301),
.C(n_290),
.Y(n_353)
);

NOR2xp33_ASAP7_75t_L g360 ( 
.A(n_354),
.B(n_331),
.Y(n_360)
);

OAI22xp5_ASAP7_75t_SL g355 ( 
.A1(n_324),
.A2(n_264),
.B1(n_274),
.B2(n_268),
.Y(n_355)
);

MAJIxp5_ASAP7_75t_L g356 ( 
.A(n_325),
.B(n_274),
.C(n_278),
.Y(n_356)
);

MAJIxp5_ASAP7_75t_L g377 ( 
.A(n_356),
.B(n_213),
.C(n_208),
.Y(n_377)
);

XNOR2xp5_ASAP7_75t_L g358 ( 
.A(n_333),
.B(n_264),
.Y(n_358)
);

NOR2xp33_ASAP7_75t_L g359 ( 
.A(n_319),
.B(n_269),
.Y(n_359)
);

NOR2xp33_ASAP7_75t_SL g379 ( 
.A(n_359),
.B(n_208),
.Y(n_379)
);

INVxp67_ASAP7_75t_L g388 ( 
.A(n_360),
.Y(n_388)
);

OAI21xp5_ASAP7_75t_SL g362 ( 
.A1(n_344),
.A2(n_313),
.B(n_317),
.Y(n_362)
);

NAND2xp5_ASAP7_75t_SL g389 ( 
.A(n_362),
.B(n_377),
.Y(n_389)
);

NOR2xp33_ASAP7_75t_L g364 ( 
.A(n_345),
.B(n_321),
.Y(n_364)
);

INVx1_ASAP7_75t_L g380 ( 
.A(n_364),
.Y(n_380)
);

INVx1_ASAP7_75t_L g365 ( 
.A(n_343),
.Y(n_365)
);

INVx1_ASAP7_75t_L g385 ( 
.A(n_365),
.Y(n_385)
);

MAJIxp5_ASAP7_75t_L g386 ( 
.A(n_367),
.B(n_371),
.C(n_372),
.Y(n_386)
);

AOI22xp5_ASAP7_75t_L g390 ( 
.A1(n_370),
.A2(n_379),
.B1(n_354),
.B2(n_350),
.Y(n_390)
);

XOR2xp5_ASAP7_75t_L g371 ( 
.A(n_338),
.B(n_280),
.Y(n_371)
);

XOR2xp5_ASAP7_75t_L g372 ( 
.A(n_338),
.B(n_296),
.Y(n_372)
);

AOI21xp5_ASAP7_75t_L g373 ( 
.A1(n_344),
.A2(n_296),
.B(n_276),
.Y(n_373)
);

HB1xp67_ASAP7_75t_L g384 ( 
.A(n_373),
.Y(n_384)
);

NOR2xp33_ASAP7_75t_L g374 ( 
.A(n_347),
.B(n_229),
.Y(n_374)
);

INVx1_ASAP7_75t_L g387 ( 
.A(n_374),
.Y(n_387)
);

NOR2xp33_ASAP7_75t_L g375 ( 
.A(n_357),
.B(n_229),
.Y(n_375)
);

INVx1_ASAP7_75t_L g393 ( 
.A(n_375),
.Y(n_393)
);

INVx1_ASAP7_75t_L g376 ( 
.A(n_337),
.Y(n_376)
);

INVx1_ASAP7_75t_L g396 ( 
.A(n_376),
.Y(n_396)
);

MAJIxp5_ASAP7_75t_L g381 ( 
.A(n_371),
.B(n_357),
.C(n_356),
.Y(n_381)
);

NAND2xp5_ASAP7_75t_L g407 ( 
.A(n_381),
.B(n_382),
.Y(n_407)
);

MAJIxp5_ASAP7_75t_L g382 ( 
.A(n_372),
.B(n_369),
.C(n_377),
.Y(n_382)
);

MAJIxp5_ASAP7_75t_L g383 ( 
.A(n_369),
.B(n_341),
.C(n_353),
.Y(n_383)
);

NAND2xp5_ASAP7_75t_SL g406 ( 
.A(n_383),
.B(n_392),
.Y(n_406)
);

INVx1_ASAP7_75t_L g398 ( 
.A(n_390),
.Y(n_398)
);

NOR2xp33_ASAP7_75t_L g391 ( 
.A(n_366),
.B(n_346),
.Y(n_391)
);

INVx1_ASAP7_75t_L g399 ( 
.A(n_391),
.Y(n_399)
);

MAJIxp5_ASAP7_75t_L g392 ( 
.A(n_363),
.B(n_340),
.C(n_358),
.Y(n_392)
);

BUFx3_ASAP7_75t_L g394 ( 
.A(n_376),
.Y(n_394)
);

CKINVDCx20_ASAP7_75t_R g400 ( 
.A(n_394),
.Y(n_400)
);

MAJIxp5_ASAP7_75t_L g395 ( 
.A(n_368),
.B(n_367),
.C(n_362),
.Y(n_395)
);

XNOR2xp5_ASAP7_75t_L g408 ( 
.A(n_395),
.B(n_225),
.Y(n_408)
);

INVxp67_ASAP7_75t_L g397 ( 
.A(n_384),
.Y(n_397)
);

INVx1_ASAP7_75t_L g419 ( 
.A(n_397),
.Y(n_419)
);

OAI21xp5_ASAP7_75t_L g401 ( 
.A1(n_382),
.A2(n_378),
.B(n_361),
.Y(n_401)
);

OR2x2_ASAP7_75t_L g423 ( 
.A(n_401),
.B(n_177),
.Y(n_423)
);

AOI22xp5_ASAP7_75t_L g402 ( 
.A1(n_380),
.A2(n_361),
.B1(n_365),
.B2(n_370),
.Y(n_402)
);

NAND2xp5_ASAP7_75t_L g414 ( 
.A(n_402),
.B(n_404),
.Y(n_414)
);

XOR2xp5_ASAP7_75t_L g403 ( 
.A(n_381),
.B(n_368),
.Y(n_403)
);

XOR2xp5_ASAP7_75t_L g415 ( 
.A(n_403),
.B(n_410),
.Y(n_415)
);

MAJIxp5_ASAP7_75t_L g404 ( 
.A(n_383),
.B(n_373),
.C(n_225),
.Y(n_404)
);

MAJIxp5_ASAP7_75t_L g405 ( 
.A(n_386),
.B(n_225),
.C(n_156),
.Y(n_405)
);

NAND2xp5_ASAP7_75t_L g417 ( 
.A(n_405),
.B(n_408),
.Y(n_417)
);

MAJIxp5_ASAP7_75t_L g409 ( 
.A(n_389),
.B(n_193),
.C(n_164),
.Y(n_409)
);

NOR2xp33_ASAP7_75t_L g412 ( 
.A(n_409),
.B(n_411),
.Y(n_412)
);

XOR2xp5_ASAP7_75t_L g410 ( 
.A(n_395),
.B(n_254),
.Y(n_410)
);

MAJIxp5_ASAP7_75t_L g411 ( 
.A(n_387),
.B(n_121),
.C(n_98),
.Y(n_411)
);

NOR2xp33_ASAP7_75t_SL g413 ( 
.A(n_407),
.B(n_396),
.Y(n_413)
);

NAND2xp5_ASAP7_75t_L g426 ( 
.A(n_413),
.B(n_420),
.Y(n_426)
);

AOI21xp5_ASAP7_75t_L g416 ( 
.A1(n_397),
.A2(n_388),
.B(n_385),
.Y(n_416)
);

AOI21xp5_ASAP7_75t_L g433 ( 
.A1(n_416),
.A2(n_421),
.B(n_423),
.Y(n_433)
);

AOI22xp5_ASAP7_75t_L g418 ( 
.A1(n_398),
.A2(n_388),
.B1(n_394),
.B2(n_393),
.Y(n_418)
);

AOI22xp5_ASAP7_75t_L g431 ( 
.A1(n_418),
.A2(n_117),
.B1(n_197),
.B2(n_189),
.Y(n_431)
);

NOR2xp33_ASAP7_75t_SL g420 ( 
.A(n_406),
.B(n_160),
.Y(n_420)
);

OAI21xp5_ASAP7_75t_SL g421 ( 
.A1(n_400),
.A2(n_109),
.B(n_223),
.Y(n_421)
);

INVx1_ASAP7_75t_L g422 ( 
.A(n_404),
.Y(n_422)
);

NAND2xp5_ASAP7_75t_L g428 ( 
.A(n_422),
.B(n_424),
.Y(n_428)
);

NOR2xp33_ASAP7_75t_L g424 ( 
.A(n_399),
.B(n_185),
.Y(n_424)
);

MAJIxp5_ASAP7_75t_L g425 ( 
.A(n_414),
.B(n_403),
.C(n_410),
.Y(n_425)
);

OR2x2_ASAP7_75t_L g440 ( 
.A(n_425),
.B(n_429),
.Y(n_440)
);

AND2x2_ASAP7_75t_L g427 ( 
.A(n_415),
.B(n_405),
.Y(n_427)
);

AO21x1_ASAP7_75t_L g438 ( 
.A1(n_427),
.A2(n_430),
.B(n_417),
.Y(n_438)
);

XNOR2xp5_ASAP7_75t_L g429 ( 
.A(n_415),
.B(n_409),
.Y(n_429)
);

NOR2xp33_ASAP7_75t_L g430 ( 
.A(n_419),
.B(n_411),
.Y(n_430)
);

NAND2xp5_ASAP7_75t_L g436 ( 
.A(n_431),
.B(n_421),
.Y(n_436)
);

OAI21xp5_ASAP7_75t_SL g432 ( 
.A1(n_416),
.A2(n_423),
.B(n_418),
.Y(n_432)
);

AOI21xp5_ASAP7_75t_L g439 ( 
.A1(n_432),
.A2(n_434),
.B(n_11),
.Y(n_439)
);

AOI21xp5_ASAP7_75t_L g434 ( 
.A1(n_412),
.A2(n_189),
.B(n_32),
.Y(n_434)
);

INVxp33_ASAP7_75t_L g435 ( 
.A(n_428),
.Y(n_435)
);

AOI21xp5_ASAP7_75t_L g444 ( 
.A1(n_435),
.A2(n_437),
.B(n_9),
.Y(n_444)
);

INVx1_ASAP7_75t_L g443 ( 
.A(n_436),
.Y(n_443)
);

CKINVDCx14_ASAP7_75t_R g437 ( 
.A(n_430),
.Y(n_437)
);

OAI21xp33_ASAP7_75t_L g442 ( 
.A1(n_438),
.A2(n_439),
.B(n_433),
.Y(n_442)
);

MAJIxp5_ASAP7_75t_L g441 ( 
.A(n_440),
.B(n_427),
.C(n_426),
.Y(n_441)
);

NAND2xp5_ASAP7_75t_L g445 ( 
.A(n_441),
.B(n_442),
.Y(n_445)
);

AO21x1_ASAP7_75t_L g446 ( 
.A1(n_444),
.A2(n_10),
.B(n_11),
.Y(n_446)
);

MAJIxp5_ASAP7_75t_L g447 ( 
.A(n_446),
.B(n_443),
.C(n_10),
.Y(n_447)
);

MAJIxp5_ASAP7_75t_L g448 ( 
.A(n_447),
.B(n_445),
.C(n_10),
.Y(n_448)
);

XNOR2xp5_ASAP7_75t_L g449 ( 
.A(n_448),
.B(n_10),
.Y(n_449)
);


endmodule