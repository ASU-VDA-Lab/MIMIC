module fake_jpeg_9115_n_250 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_250);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_250;

wire n_159;
wire n_117;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_57;
wire n_21;
wire n_223;
wire n_234;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_24;
wire n_44;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_170;
wire n_162;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_216;
wire n_217;
wire n_184;
wire n_53;
wire n_33;
wire n_91;
wire n_93;
wire n_54;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_5),
.Y(n_15)
);

BUFx6f_ASAP7_75t_L g16 ( 
.A(n_10),
.Y(n_16)
);

BUFx5_ASAP7_75t_L g17 ( 
.A(n_8),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_1),
.Y(n_18)
);

INVx5_ASAP7_75t_L g19 ( 
.A(n_9),
.Y(n_19)
);

INVx2_ASAP7_75t_L g20 ( 
.A(n_14),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_9),
.Y(n_21)
);

NOR2xp33_ASAP7_75t_L g22 ( 
.A(n_13),
.B(n_12),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_8),
.Y(n_23)
);

INVx6_ASAP7_75t_L g24 ( 
.A(n_1),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_5),
.Y(n_25)
);

BUFx12f_ASAP7_75t_L g26 ( 
.A(n_11),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_4),
.Y(n_27)
);

BUFx12f_ASAP7_75t_L g28 ( 
.A(n_5),
.Y(n_28)
);

INVx11_ASAP7_75t_L g29 ( 
.A(n_10),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_3),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_8),
.Y(n_31)
);

INVx2_ASAP7_75t_L g32 ( 
.A(n_29),
.Y(n_32)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_32),
.B(n_38),
.Y(n_50)
);

INVx5_ASAP7_75t_L g33 ( 
.A(n_19),
.Y(n_33)
);

INVx2_ASAP7_75t_L g53 ( 
.A(n_33),
.Y(n_53)
);

AND2x2_ASAP7_75t_SL g34 ( 
.A(n_17),
.B(n_0),
.Y(n_34)
);

AND2x2_ASAP7_75t_L g45 ( 
.A(n_34),
.B(n_37),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g35 ( 
.A(n_22),
.B(n_14),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_SL g64 ( 
.A(n_35),
.B(n_12),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_28),
.Y(n_36)
);

INVx6_ASAP7_75t_L g58 ( 
.A(n_36),
.Y(n_58)
);

AOI21xp33_ASAP7_75t_L g37 ( 
.A1(n_22),
.A2(n_0),
.B(n_1),
.Y(n_37)
);

INVx3_ASAP7_75t_L g38 ( 
.A(n_16),
.Y(n_38)
);

BUFx5_ASAP7_75t_L g39 ( 
.A(n_17),
.Y(n_39)
);

BUFx5_ASAP7_75t_L g65 ( 
.A(n_39),
.Y(n_65)
);

INVx2_ASAP7_75t_L g40 ( 
.A(n_29),
.Y(n_40)
);

INVx8_ASAP7_75t_L g47 ( 
.A(n_40),
.Y(n_47)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_17),
.Y(n_41)
);

NAND2xp5_ASAP7_75t_SL g54 ( 
.A(n_41),
.B(n_42),
.Y(n_54)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_31),
.Y(n_42)
);

NAND2xp5_ASAP7_75t_L g43 ( 
.A(n_34),
.B(n_20),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_43),
.B(n_49),
.Y(n_66)
);

OAI22xp5_ASAP7_75t_L g44 ( 
.A1(n_38),
.A2(n_20),
.B1(n_24),
.B2(n_19),
.Y(n_44)
);

OAI22xp5_ASAP7_75t_SL g77 ( 
.A1(n_44),
.A2(n_48),
.B1(n_52),
.B2(n_59),
.Y(n_77)
);

AOI22xp33_ASAP7_75t_SL g46 ( 
.A1(n_33),
.A2(n_24),
.B1(n_20),
.B2(n_19),
.Y(n_46)
);

AOI22xp33_ASAP7_75t_SL g69 ( 
.A1(n_46),
.A2(n_56),
.B1(n_32),
.B2(n_27),
.Y(n_69)
);

AOI22xp33_ASAP7_75t_L g48 ( 
.A1(n_38),
.A2(n_24),
.B1(n_29),
.B2(n_25),
.Y(n_48)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_34),
.Y(n_49)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_42),
.Y(n_51)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_51),
.Y(n_78)
);

OAI22xp33_ASAP7_75t_SL g52 ( 
.A1(n_33),
.A2(n_24),
.B1(n_25),
.B2(n_31),
.Y(n_52)
);

INVx3_ASAP7_75t_L g55 ( 
.A(n_36),
.Y(n_55)
);

INVx4_ASAP7_75t_L g82 ( 
.A(n_55),
.Y(n_82)
);

AOI22xp33_ASAP7_75t_SL g56 ( 
.A1(n_40),
.A2(n_31),
.B1(n_25),
.B2(n_23),
.Y(n_56)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_34),
.Y(n_57)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_57),
.Y(n_80)
);

AOI22xp5_ASAP7_75t_L g59 ( 
.A1(n_32),
.A2(n_16),
.B1(n_23),
.B2(n_21),
.Y(n_59)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_34),
.Y(n_60)
);

AND2x2_ASAP7_75t_L g73 ( 
.A(n_60),
.B(n_63),
.Y(n_73)
);

OAI22xp5_ASAP7_75t_SL g61 ( 
.A1(n_37),
.A2(n_30),
.B1(n_18),
.B2(n_27),
.Y(n_61)
);

OAI22xp5_ASAP7_75t_SL g84 ( 
.A1(n_61),
.A2(n_15),
.B1(n_26),
.B2(n_28),
.Y(n_84)
);

BUFx2_ASAP7_75t_L g62 ( 
.A(n_39),
.Y(n_62)
);

CKINVDCx16_ASAP7_75t_R g68 ( 
.A(n_62),
.Y(n_68)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_39),
.Y(n_63)
);

CKINVDCx20_ASAP7_75t_R g81 ( 
.A(n_64),
.Y(n_81)
);

AOI21xp33_ASAP7_75t_L g67 ( 
.A1(n_45),
.A2(n_35),
.B(n_18),
.Y(n_67)
);

MAJIxp5_ASAP7_75t_L g88 ( 
.A(n_67),
.B(n_70),
.C(n_61),
.Y(n_88)
);

AOI21xp5_ASAP7_75t_L g99 ( 
.A1(n_69),
.A2(n_75),
.B(n_56),
.Y(n_99)
);

MAJIxp5_ASAP7_75t_L g70 ( 
.A(n_57),
.B(n_41),
.C(n_36),
.Y(n_70)
);

BUFx2_ASAP7_75t_L g71 ( 
.A(n_65),
.Y(n_71)
);

CKINVDCx20_ASAP7_75t_R g87 ( 
.A(n_71),
.Y(n_87)
);

INVxp67_ASAP7_75t_L g72 ( 
.A(n_65),
.Y(n_72)
);

INVx4_ASAP7_75t_SL g97 ( 
.A(n_72),
.Y(n_97)
);

OA22x2_ASAP7_75t_L g74 ( 
.A1(n_49),
.A2(n_36),
.B1(n_28),
.B2(n_26),
.Y(n_74)
);

OAI22xp5_ASAP7_75t_SL g106 ( 
.A1(n_74),
.A2(n_79),
.B1(n_83),
.B2(n_48),
.Y(n_106)
);

AND2x2_ASAP7_75t_L g75 ( 
.A(n_60),
.B(n_0),
.Y(n_75)
);

NAND2xp33_ASAP7_75t_SL g76 ( 
.A(n_43),
.B(n_0),
.Y(n_76)
);

OR2x2_ASAP7_75t_SL g89 ( 
.A(n_76),
.B(n_51),
.Y(n_89)
);

AOI22xp33_ASAP7_75t_L g79 ( 
.A1(n_53),
.A2(n_16),
.B1(n_21),
.B2(n_30),
.Y(n_79)
);

OAI22xp5_ASAP7_75t_L g83 ( 
.A1(n_46),
.A2(n_16),
.B1(n_15),
.B2(n_26),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_SL g105 ( 
.A(n_84),
.B(n_52),
.Y(n_105)
);

INVx13_ASAP7_75t_L g85 ( 
.A(n_65),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_85),
.B(n_86),
.Y(n_92)
);

INVx13_ASAP7_75t_L g86 ( 
.A(n_62),
.Y(n_86)
);

AND2x2_ASAP7_75t_L g131 ( 
.A(n_88),
.B(n_105),
.Y(n_131)
);

OAI21xp33_ASAP7_75t_L g122 ( 
.A1(n_89),
.A2(n_75),
.B(n_73),
.Y(n_122)
);

INVxp67_ASAP7_75t_L g90 ( 
.A(n_69),
.Y(n_90)
);

INVxp67_ASAP7_75t_L g120 ( 
.A(n_90),
.Y(n_120)
);

INVx3_ASAP7_75t_L g91 ( 
.A(n_86),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_91),
.B(n_93),
.Y(n_128)
);

INVx13_ASAP7_75t_L g93 ( 
.A(n_71),
.Y(n_93)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_74),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_SL g114 ( 
.A(n_94),
.B(n_101),
.Y(n_114)
);

INVx2_ASAP7_75t_L g95 ( 
.A(n_82),
.Y(n_95)
);

CKINVDCx20_ASAP7_75t_R g119 ( 
.A(n_95),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_78),
.B(n_54),
.Y(n_96)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_96),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_78),
.B(n_54),
.Y(n_98)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_98),
.Y(n_117)
);

OAI21xp5_ASAP7_75t_SL g112 ( 
.A1(n_99),
.A2(n_102),
.B(n_84),
.Y(n_112)
);

BUFx12f_ASAP7_75t_L g100 ( 
.A(n_71),
.Y(n_100)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_100),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_81),
.B(n_64),
.Y(n_101)
);

AND2x6_ASAP7_75t_L g102 ( 
.A(n_67),
.B(n_45),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_L g103 ( 
.A(n_66),
.B(n_45),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_L g110 ( 
.A(n_103),
.B(n_107),
.Y(n_110)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_74),
.Y(n_104)
);

AOI22xp33_ASAP7_75t_SL g123 ( 
.A1(n_104),
.A2(n_108),
.B1(n_82),
.B2(n_47),
.Y(n_123)
);

AOI22xp5_ASAP7_75t_L g113 ( 
.A1(n_106),
.A2(n_109),
.B1(n_77),
.B2(n_53),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_SL g107 ( 
.A(n_75),
.B(n_45),
.Y(n_107)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_74),
.Y(n_108)
);

OAI22xp5_ASAP7_75t_SL g109 ( 
.A1(n_70),
.A2(n_59),
.B1(n_50),
.B2(n_47),
.Y(n_109)
);

OAI22xp5_ASAP7_75t_SL g111 ( 
.A1(n_94),
.A2(n_70),
.B1(n_80),
.B2(n_77),
.Y(n_111)
);

AOI22xp5_ASAP7_75t_L g132 ( 
.A1(n_111),
.A2(n_107),
.B1(n_102),
.B2(n_89),
.Y(n_132)
);

AOI21xp5_ASAP7_75t_L g153 ( 
.A1(n_112),
.A2(n_123),
.B(n_129),
.Y(n_153)
);

OAI22xp5_ASAP7_75t_SL g140 ( 
.A1(n_113),
.A2(n_121),
.B1(n_126),
.B2(n_127),
.Y(n_140)
);

MAJIxp5_ASAP7_75t_L g116 ( 
.A(n_88),
.B(n_66),
.C(n_80),
.Y(n_116)
);

MAJIxp5_ASAP7_75t_L g146 ( 
.A(n_116),
.B(n_118),
.C(n_92),
.Y(n_146)
);

MAJIxp5_ASAP7_75t_L g118 ( 
.A(n_103),
.B(n_73),
.C(n_74),
.Y(n_118)
);

AOI22xp5_ASAP7_75t_L g121 ( 
.A1(n_106),
.A2(n_74),
.B1(n_76),
.B2(n_83),
.Y(n_121)
);

OAI21xp5_ASAP7_75t_L g133 ( 
.A1(n_122),
.A2(n_125),
.B(n_114),
.Y(n_133)
);

AOI21xp5_ASAP7_75t_L g125 ( 
.A1(n_104),
.A2(n_73),
.B(n_75),
.Y(n_125)
);

OAI21xp5_ASAP7_75t_SL g134 ( 
.A1(n_125),
.A2(n_114),
.B(n_110),
.Y(n_134)
);

AOI22xp5_ASAP7_75t_L g126 ( 
.A1(n_109),
.A2(n_73),
.B1(n_47),
.B2(n_50),
.Y(n_126)
);

AOI22xp5_ASAP7_75t_L g127 ( 
.A1(n_108),
.A2(n_58),
.B1(n_55),
.B2(n_82),
.Y(n_127)
);

A2O1A1Ixp33_ASAP7_75t_SL g129 ( 
.A1(n_99),
.A2(n_44),
.B(n_63),
.C(n_71),
.Y(n_129)
);

AOI22xp5_ASAP7_75t_L g130 ( 
.A1(n_105),
.A2(n_58),
.B1(n_55),
.B2(n_81),
.Y(n_130)
);

OAI22xp5_ASAP7_75t_SL g141 ( 
.A1(n_130),
.A2(n_96),
.B1(n_79),
.B2(n_58),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_L g170 ( 
.A(n_132),
.B(n_135),
.Y(n_170)
);

OAI21xp5_ASAP7_75t_SL g165 ( 
.A1(n_133),
.A2(n_134),
.B(n_138),
.Y(n_165)
);

INVx13_ASAP7_75t_L g135 ( 
.A(n_128),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_SL g136 ( 
.A(n_115),
.B(n_101),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_SL g168 ( 
.A(n_136),
.B(n_137),
.Y(n_168)
);

NOR2xp33_ASAP7_75t_L g137 ( 
.A(n_115),
.B(n_87),
.Y(n_137)
);

AND2x2_ASAP7_75t_L g138 ( 
.A(n_118),
.B(n_85),
.Y(n_138)
);

XNOR2xp5_ASAP7_75t_L g139 ( 
.A(n_116),
.B(n_98),
.Y(n_139)
);

MAJIxp5_ASAP7_75t_L g156 ( 
.A(n_139),
.B(n_146),
.C(n_126),
.Y(n_156)
);

AOI22xp5_ASAP7_75t_L g158 ( 
.A1(n_141),
.A2(n_145),
.B1(n_144),
.B2(n_140),
.Y(n_158)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_128),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_SL g169 ( 
.A(n_142),
.B(n_143),
.Y(n_169)
);

CKINVDCx14_ASAP7_75t_R g143 ( 
.A(n_130),
.Y(n_143)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_127),
.Y(n_144)
);

NOR2xp33_ASAP7_75t_L g173 ( 
.A(n_144),
.B(n_148),
.Y(n_173)
);

OAI22xp5_ASAP7_75t_SL g145 ( 
.A1(n_113),
.A2(n_87),
.B1(n_97),
.B2(n_68),
.Y(n_145)
);

OAI22xp5_ASAP7_75t_L g147 ( 
.A1(n_123),
.A2(n_95),
.B1(n_85),
.B2(n_97),
.Y(n_147)
);

OAI22xp5_ASAP7_75t_L g160 ( 
.A1(n_147),
.A2(n_149),
.B1(n_93),
.B2(n_86),
.Y(n_160)
);

CKINVDCx20_ASAP7_75t_R g148 ( 
.A(n_119),
.Y(n_148)
);

OAI22xp5_ASAP7_75t_L g149 ( 
.A1(n_121),
.A2(n_97),
.B1(n_68),
.B2(n_93),
.Y(n_149)
);

INVx2_ASAP7_75t_L g150 ( 
.A(n_119),
.Y(n_150)
);

CKINVDCx20_ASAP7_75t_R g162 ( 
.A(n_150),
.Y(n_162)
);

NOR2xp33_ASAP7_75t_SL g151 ( 
.A(n_117),
.B(n_12),
.Y(n_151)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_151),
.Y(n_166)
);

NOR2xp33_ASAP7_75t_L g152 ( 
.A(n_124),
.B(n_100),
.Y(n_152)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_152),
.Y(n_167)
);

INVx6_ASAP7_75t_L g154 ( 
.A(n_124),
.Y(n_154)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_154),
.Y(n_175)
);

NAND3xp33_ASAP7_75t_SL g155 ( 
.A(n_153),
.B(n_110),
.C(n_112),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_L g190 ( 
.A(n_155),
.B(n_161),
.Y(n_190)
);

MAJIxp5_ASAP7_75t_L g181 ( 
.A(n_156),
.B(n_157),
.C(n_163),
.Y(n_181)
);

XOR2xp5_ASAP7_75t_L g157 ( 
.A(n_132),
.B(n_131),
.Y(n_157)
);

OAI22xp5_ASAP7_75t_L g179 ( 
.A1(n_158),
.A2(n_160),
.B1(n_150),
.B2(n_148),
.Y(n_179)
);

AOI22xp5_ASAP7_75t_L g159 ( 
.A1(n_140),
.A2(n_111),
.B1(n_129),
.B2(n_120),
.Y(n_159)
);

OAI22xp5_ASAP7_75t_SL g178 ( 
.A1(n_159),
.A2(n_164),
.B1(n_129),
.B2(n_149),
.Y(n_178)
);

NAND3xp33_ASAP7_75t_L g161 ( 
.A(n_136),
.B(n_117),
.C(n_131),
.Y(n_161)
);

MAJIxp5_ASAP7_75t_L g163 ( 
.A(n_146),
.B(n_139),
.C(n_134),
.Y(n_163)
);

AOI22xp5_ASAP7_75t_L g164 ( 
.A1(n_145),
.A2(n_129),
.B1(n_131),
.B2(n_91),
.Y(n_164)
);

OAI221xp5_ASAP7_75t_L g171 ( 
.A1(n_133),
.A2(n_129),
.B1(n_62),
.B2(n_28),
.C(n_26),
.Y(n_171)
);

CKINVDCx20_ASAP7_75t_R g177 ( 
.A(n_171),
.Y(n_177)
);

INVx4_ASAP7_75t_L g172 ( 
.A(n_154),
.Y(n_172)
);

CKINVDCx20_ASAP7_75t_R g180 ( 
.A(n_172),
.Y(n_180)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_137),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_L g191 ( 
.A(n_174),
.B(n_100),
.Y(n_191)
);

AOI22xp5_ASAP7_75t_L g176 ( 
.A1(n_170),
.A2(n_153),
.B1(n_141),
.B2(n_129),
.Y(n_176)
);

OAI22xp5_ASAP7_75t_SL g194 ( 
.A1(n_176),
.A2(n_192),
.B1(n_193),
.B2(n_175),
.Y(n_194)
);

AOI22xp5_ASAP7_75t_L g197 ( 
.A1(n_178),
.A2(n_188),
.B1(n_177),
.B2(n_183),
.Y(n_197)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_179),
.Y(n_208)
);

MAJIxp5_ASAP7_75t_L g182 ( 
.A(n_163),
.B(n_138),
.C(n_142),
.Y(n_182)
);

XOR2xp5_ASAP7_75t_L g200 ( 
.A(n_182),
.B(n_186),
.Y(n_200)
);

XNOR2x2_ASAP7_75t_L g183 ( 
.A(n_171),
.B(n_138),
.Y(n_183)
);

AOI21xp5_ASAP7_75t_L g202 ( 
.A1(n_183),
.A2(n_184),
.B(n_167),
.Y(n_202)
);

AOI21xp5_ASAP7_75t_L g184 ( 
.A1(n_165),
.A2(n_173),
.B(n_174),
.Y(n_184)
);

OAI22xp5_ASAP7_75t_L g185 ( 
.A1(n_158),
.A2(n_135),
.B1(n_147),
.B2(n_154),
.Y(n_185)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_185),
.Y(n_198)
);

XOR2xp5_ASAP7_75t_L g186 ( 
.A(n_157),
.B(n_135),
.Y(n_186)
);

CKINVDCx16_ASAP7_75t_R g187 ( 
.A(n_169),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_SL g195 ( 
.A(n_187),
.B(n_189),
.Y(n_195)
);

INVxp67_ASAP7_75t_L g188 ( 
.A(n_164),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_L g199 ( 
.A(n_188),
.B(n_191),
.Y(n_199)
);

OAI22xp5_ASAP7_75t_L g189 ( 
.A1(n_159),
.A2(n_151),
.B1(n_100),
.B2(n_3),
.Y(n_189)
);

AOI22xp5_ASAP7_75t_L g192 ( 
.A1(n_168),
.A2(n_28),
.B1(n_26),
.B2(n_3),
.Y(n_192)
);

AOI22xp5_ASAP7_75t_L g193 ( 
.A1(n_168),
.A2(n_175),
.B1(n_162),
.B2(n_172),
.Y(n_193)
);

CKINVDCx14_ASAP7_75t_R g220 ( 
.A(n_194),
.Y(n_220)
);

NOR2xp33_ASAP7_75t_SL g196 ( 
.A(n_190),
.B(n_166),
.Y(n_196)
);

NAND2xp5_ASAP7_75t_SL g214 ( 
.A(n_196),
.B(n_206),
.Y(n_214)
);

OAI22xp5_ASAP7_75t_SL g218 ( 
.A1(n_197),
.A2(n_201),
.B1(n_205),
.B2(n_191),
.Y(n_218)
);

AOI22xp5_ASAP7_75t_L g201 ( 
.A1(n_178),
.A2(n_162),
.B1(n_167),
.B2(n_165),
.Y(n_201)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_202),
.Y(n_212)
);

INVx2_ASAP7_75t_SL g203 ( 
.A(n_180),
.Y(n_203)
);

AOI22xp33_ASAP7_75t_SL g209 ( 
.A1(n_203),
.A2(n_204),
.B1(n_207),
.B2(n_184),
.Y(n_209)
);

AOI21xp5_ASAP7_75t_L g204 ( 
.A1(n_177),
.A2(n_183),
.B(n_185),
.Y(n_204)
);

OAI22xp5_ASAP7_75t_SL g205 ( 
.A1(n_176),
.A2(n_156),
.B1(n_166),
.B2(n_3),
.Y(n_205)
);

NOR2xp33_ASAP7_75t_L g206 ( 
.A(n_180),
.B(n_26),
.Y(n_206)
);

BUFx2_ASAP7_75t_L g207 ( 
.A(n_193),
.Y(n_207)
);

OAI22xp5_ASAP7_75t_SL g222 ( 
.A1(n_209),
.A2(n_197),
.B1(n_208),
.B2(n_203),
.Y(n_222)
);

AOI21xp5_ASAP7_75t_L g210 ( 
.A1(n_199),
.A2(n_198),
.B(n_190),
.Y(n_210)
);

MAJIxp5_ASAP7_75t_L g224 ( 
.A(n_210),
.B(n_211),
.C(n_215),
.Y(n_224)
);

XNOR2xp5_ASAP7_75t_L g211 ( 
.A(n_202),
.B(n_181),
.Y(n_211)
);

MAJIxp5_ASAP7_75t_L g213 ( 
.A(n_200),
.B(n_181),
.C(n_182),
.Y(n_213)
);

MAJIxp5_ASAP7_75t_L g229 ( 
.A(n_213),
.B(n_219),
.C(n_11),
.Y(n_229)
);

XNOR2xp5_ASAP7_75t_L g215 ( 
.A(n_201),
.B(n_186),
.Y(n_215)
);

MAJIxp5_ASAP7_75t_L g216 ( 
.A(n_200),
.B(n_199),
.C(n_205),
.Y(n_216)
);

MAJIxp5_ASAP7_75t_L g226 ( 
.A(n_216),
.B(n_213),
.C(n_215),
.Y(n_226)
);

XOR2xp5_ASAP7_75t_SL g217 ( 
.A(n_204),
.B(n_192),
.Y(n_217)
);

XOR2xp5_ASAP7_75t_L g221 ( 
.A(n_217),
.B(n_218),
.Y(n_221)
);

MAJIxp5_ASAP7_75t_L g219 ( 
.A(n_194),
.B(n_28),
.C(n_2),
.Y(n_219)
);

AOI22xp5_ASAP7_75t_SL g232 ( 
.A1(n_222),
.A2(n_223),
.B1(n_220),
.B2(n_2),
.Y(n_232)
);

AOI22xp33_ASAP7_75t_SL g223 ( 
.A1(n_212),
.A2(n_203),
.B1(n_207),
.B2(n_195),
.Y(n_223)
);

AND2x2_ASAP7_75t_L g225 ( 
.A(n_216),
.B(n_14),
.Y(n_225)
);

OR2x2_ASAP7_75t_L g233 ( 
.A(n_225),
.B(n_10),
.Y(n_233)
);

XNOR2xp5_ASAP7_75t_L g235 ( 
.A(n_226),
.B(n_228),
.Y(n_235)
);

MAJIxp5_ASAP7_75t_L g227 ( 
.A(n_211),
.B(n_13),
.C(n_11),
.Y(n_227)
);

NAND2xp5_ASAP7_75t_L g236 ( 
.A(n_227),
.B(n_1),
.Y(n_236)
);

XOR2xp5_ASAP7_75t_L g228 ( 
.A(n_218),
.B(n_13),
.Y(n_228)
);

OAI21xp5_ASAP7_75t_L g230 ( 
.A1(n_229),
.A2(n_214),
.B(n_217),
.Y(n_230)
);

NAND2xp5_ASAP7_75t_L g240 ( 
.A(n_230),
.B(n_231),
.Y(n_240)
);

NOR2xp33_ASAP7_75t_L g231 ( 
.A(n_228),
.B(n_219),
.Y(n_231)
);

OAI21xp5_ASAP7_75t_L g241 ( 
.A1(n_232),
.A2(n_234),
.B(n_236),
.Y(n_241)
);

AO22x1_ASAP7_75t_L g239 ( 
.A1(n_233),
.A2(n_223),
.B1(n_4),
.B2(n_5),
.Y(n_239)
);

NOR2xp33_ASAP7_75t_L g234 ( 
.A(n_221),
.B(n_9),
.Y(n_234)
);

AND2x2_ASAP7_75t_L g237 ( 
.A(n_235),
.B(n_224),
.Y(n_237)
);

NAND2xp5_ASAP7_75t_L g242 ( 
.A(n_237),
.B(n_238),
.Y(n_242)
);

HB1xp67_ASAP7_75t_L g238 ( 
.A(n_232),
.Y(n_238)
);

AOI22xp33_ASAP7_75t_L g244 ( 
.A1(n_239),
.A2(n_233),
.B1(n_4),
.B2(n_6),
.Y(n_244)
);

MAJIxp5_ASAP7_75t_L g243 ( 
.A(n_240),
.B(n_221),
.C(n_225),
.Y(n_243)
);

NAND2xp5_ASAP7_75t_L g247 ( 
.A(n_243),
.B(n_6),
.Y(n_247)
);

AOI332xp33_ASAP7_75t_L g246 ( 
.A1(n_244),
.A2(n_245),
.A3(n_2),
.B1(n_6),
.B2(n_7),
.B3(n_233),
.C1(n_217),
.C2(n_239),
.Y(n_246)
);

FAx1_ASAP7_75t_SL g245 ( 
.A(n_241),
.B(n_2),
.CI(n_4),
.CON(n_245),
.SN(n_245)
);

MAJIxp5_ASAP7_75t_L g248 ( 
.A(n_246),
.B(n_247),
.C(n_243),
.Y(n_248)
);

O2A1O1Ixp33_ASAP7_75t_SL g249 ( 
.A1(n_248),
.A2(n_242),
.B(n_245),
.C(n_6),
.Y(n_249)
);

XNOR2xp5_ASAP7_75t_L g250 ( 
.A(n_249),
.B(n_245),
.Y(n_250)
);


endmodule