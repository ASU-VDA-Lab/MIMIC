module fake_jpeg_12916_n_387 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_387);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_387;

wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_385;
wire n_228;
wire n_134;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_340;
wire n_381;
wire n_377;
wire n_291;
wire n_236;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_370;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_39;
wire n_371;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_382;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_352;
wire n_350;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_384;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_360;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_378;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_379;
wire n_114;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_356;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_375;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_247;
wire n_157;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVx1_ASAP7_75t_L g17 ( 
.A(n_16),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_5),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_4),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_16),
.Y(n_20)
);

BUFx3_ASAP7_75t_L g21 ( 
.A(n_4),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_4),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_3),
.Y(n_23)
);

BUFx6f_ASAP7_75t_SL g24 ( 
.A(n_16),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_7),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_15),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_0),
.Y(n_27)
);

BUFx10_ASAP7_75t_L g28 ( 
.A(n_12),
.Y(n_28)
);

INVx3_ASAP7_75t_L g29 ( 
.A(n_14),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_10),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_8),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_13),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_14),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_0),
.Y(n_34)
);

INVx1_ASAP7_75t_SL g35 ( 
.A(n_12),
.Y(n_35)
);

BUFx5_ASAP7_75t_L g36 ( 
.A(n_2),
.Y(n_36)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_7),
.Y(n_37)
);

INVx2_ASAP7_75t_L g38 ( 
.A(n_5),
.Y(n_38)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_7),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_8),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_5),
.Y(n_41)
);

INVx4_ASAP7_75t_L g42 ( 
.A(n_8),
.Y(n_42)
);

INVx4_ASAP7_75t_L g43 ( 
.A(n_0),
.Y(n_43)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_6),
.Y(n_44)
);

INVx4_ASAP7_75t_L g45 ( 
.A(n_11),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_15),
.Y(n_46)
);

INVx2_ASAP7_75t_L g47 ( 
.A(n_10),
.Y(n_47)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_10),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_12),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_11),
.Y(n_50)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_14),
.Y(n_51)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_15),
.Y(n_52)
);

INVx8_ASAP7_75t_L g53 ( 
.A(n_13),
.Y(n_53)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_3),
.Y(n_54)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_13),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_19),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g130 ( 
.A(n_56),
.Y(n_130)
);

INVxp67_ASAP7_75t_L g57 ( 
.A(n_17),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g144 ( 
.A(n_57),
.B(n_76),
.Y(n_144)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_18),
.B(n_3),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_SL g161 ( 
.A(n_58),
.B(n_59),
.Y(n_161)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_18),
.B(n_6),
.Y(n_59)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_38),
.Y(n_60)
);

INVx2_ASAP7_75t_L g114 ( 
.A(n_60),
.Y(n_114)
);

INVx5_ASAP7_75t_L g61 ( 
.A(n_43),
.Y(n_61)
);

INVx4_ASAP7_75t_L g115 ( 
.A(n_61),
.Y(n_115)
);

INVx8_ASAP7_75t_L g62 ( 
.A(n_36),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g175 ( 
.A(n_62),
.Y(n_175)
);

INVx3_ASAP7_75t_L g63 ( 
.A(n_42),
.Y(n_63)
);

HB1xp67_ASAP7_75t_L g147 ( 
.A(n_63),
.Y(n_147)
);

INVx11_ASAP7_75t_L g64 ( 
.A(n_24),
.Y(n_64)
);

INVx11_ASAP7_75t_L g122 ( 
.A(n_64),
.Y(n_122)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_19),
.Y(n_65)
);

INVx4_ASAP7_75t_L g151 ( 
.A(n_65),
.Y(n_151)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_38),
.Y(n_66)
);

INVx2_ASAP7_75t_L g128 ( 
.A(n_66),
.Y(n_128)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_55),
.Y(n_67)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_67),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_20),
.B(n_6),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_SL g123 ( 
.A(n_68),
.B(n_71),
.Y(n_123)
);

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_19),
.Y(n_69)
);

INVx4_ASAP7_75t_L g160 ( 
.A(n_69),
.Y(n_160)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_17),
.Y(n_70)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_70),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_20),
.B(n_9),
.Y(n_71)
);

INVx8_ASAP7_75t_L g72 ( 
.A(n_36),
.Y(n_72)
);

INVx3_ASAP7_75t_L g113 ( 
.A(n_72),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_22),
.B(n_9),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_SL g136 ( 
.A(n_73),
.B(n_99),
.Y(n_136)
);

BUFx10_ASAP7_75t_L g74 ( 
.A(n_24),
.Y(n_74)
);

CKINVDCx16_ASAP7_75t_R g127 ( 
.A(n_74),
.Y(n_127)
);

INVx2_ASAP7_75t_SL g75 ( 
.A(n_28),
.Y(n_75)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_75),
.Y(n_145)
);

CKINVDCx20_ASAP7_75t_R g76 ( 
.A(n_28),
.Y(n_76)
);

INVx8_ASAP7_75t_L g77 ( 
.A(n_28),
.Y(n_77)
);

INVx3_ASAP7_75t_L g143 ( 
.A(n_77),
.Y(n_143)
);

INVx11_ASAP7_75t_L g78 ( 
.A(n_28),
.Y(n_78)
);

INVx11_ASAP7_75t_L g150 ( 
.A(n_78),
.Y(n_150)
);

AND2x2_ASAP7_75t_L g79 ( 
.A(n_35),
.B(n_9),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g148 ( 
.A(n_79),
.B(n_82),
.Y(n_148)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_26),
.Y(n_80)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_80),
.Y(n_157)
);

BUFx5_ASAP7_75t_L g81 ( 
.A(n_28),
.Y(n_81)
);

INVx3_ASAP7_75t_L g163 ( 
.A(n_81),
.Y(n_163)
);

CKINVDCx20_ASAP7_75t_R g82 ( 
.A(n_22),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_SL g83 ( 
.A(n_23),
.B(n_11),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g156 ( 
.A(n_83),
.B(n_93),
.Y(n_156)
);

INVx3_ASAP7_75t_L g84 ( 
.A(n_42),
.Y(n_84)
);

INVx3_ASAP7_75t_L g169 ( 
.A(n_84),
.Y(n_169)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_55),
.Y(n_85)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_85),
.Y(n_158)
);

INVx6_ASAP7_75t_SL g86 ( 
.A(n_35),
.Y(n_86)
);

CKINVDCx12_ASAP7_75t_R g119 ( 
.A(n_86),
.Y(n_119)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_54),
.Y(n_87)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_87),
.Y(n_172)
);

BUFx12f_ASAP7_75t_L g88 ( 
.A(n_21),
.Y(n_88)
);

BUFx12_ASAP7_75t_L g174 ( 
.A(n_88),
.Y(n_174)
);

BUFx8_ASAP7_75t_L g89 ( 
.A(n_53),
.Y(n_89)
);

AND2x2_ASAP7_75t_L g167 ( 
.A(n_89),
.B(n_95),
.Y(n_167)
);

INVx4_ASAP7_75t_L g90 ( 
.A(n_43),
.Y(n_90)
);

INVx2_ASAP7_75t_L g131 ( 
.A(n_90),
.Y(n_131)
);

INVx3_ASAP7_75t_L g91 ( 
.A(n_45),
.Y(n_91)
);

INVx2_ASAP7_75t_L g134 ( 
.A(n_91),
.Y(n_134)
);

BUFx3_ASAP7_75t_L g92 ( 
.A(n_21),
.Y(n_92)
);

INVx2_ASAP7_75t_L g135 ( 
.A(n_92),
.Y(n_135)
);

BUFx12f_ASAP7_75t_L g93 ( 
.A(n_21),
.Y(n_93)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_54),
.Y(n_94)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_94),
.Y(n_176)
);

BUFx5_ASAP7_75t_L g95 ( 
.A(n_30),
.Y(n_95)
);

INVx3_ASAP7_75t_L g96 ( 
.A(n_45),
.Y(n_96)
);

INVx2_ASAP7_75t_L g152 ( 
.A(n_96),
.Y(n_152)
);

INVx4_ASAP7_75t_L g97 ( 
.A(n_29),
.Y(n_97)
);

INVx2_ASAP7_75t_L g153 ( 
.A(n_97),
.Y(n_153)
);

BUFx12f_ASAP7_75t_L g98 ( 
.A(n_30),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g166 ( 
.A(n_98),
.B(n_101),
.Y(n_166)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_23),
.B(n_0),
.Y(n_99)
);

INVx2_ASAP7_75t_L g100 ( 
.A(n_47),
.Y(n_100)
);

INVx2_ASAP7_75t_L g154 ( 
.A(n_100),
.Y(n_154)
);

BUFx12f_ASAP7_75t_L g101 ( 
.A(n_30),
.Y(n_101)
);

INVx3_ASAP7_75t_L g102 ( 
.A(n_29),
.Y(n_102)
);

INVx2_ASAP7_75t_L g173 ( 
.A(n_102),
.Y(n_173)
);

INVx2_ASAP7_75t_L g103 ( 
.A(n_47),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g170 ( 
.A(n_103),
.B(n_104),
.Y(n_170)
);

INVx2_ASAP7_75t_L g104 ( 
.A(n_40),
.Y(n_104)
);

AND2x2_ASAP7_75t_L g105 ( 
.A(n_53),
.B(n_1),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g177 ( 
.A(n_105),
.B(n_106),
.Y(n_177)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_26),
.Y(n_106)
);

BUFx6f_ASAP7_75t_L g107 ( 
.A(n_40),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_L g117 ( 
.A(n_107),
.B(n_49),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_SL g108 ( 
.A(n_25),
.B(n_1),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_SL g162 ( 
.A(n_108),
.B(n_109),
.Y(n_162)
);

CKINVDCx20_ASAP7_75t_R g109 ( 
.A(n_25),
.Y(n_109)
);

INVx8_ASAP7_75t_L g110 ( 
.A(n_40),
.Y(n_110)
);

AOI22xp33_ASAP7_75t_SL g118 ( 
.A1(n_110),
.A2(n_112),
.B1(n_53),
.B2(n_49),
.Y(n_118)
);

CKINVDCx20_ASAP7_75t_R g111 ( 
.A(n_31),
.Y(n_111)
);

CKINVDCx20_ASAP7_75t_R g129 ( 
.A(n_111),
.Y(n_129)
);

INVx8_ASAP7_75t_L g112 ( 
.A(n_49),
.Y(n_112)
);

OAI21xp5_ASAP7_75t_SL g116 ( 
.A1(n_105),
.A2(n_37),
.B(n_51),
.Y(n_116)
);

XNOR2xp5_ASAP7_75t_L g194 ( 
.A(n_116),
.B(n_2),
.Y(n_194)
);

AND2x2_ASAP7_75t_L g201 ( 
.A(n_117),
.B(n_149),
.Y(n_201)
);

INVx5_ASAP7_75t_L g225 ( 
.A(n_118),
.Y(n_225)
);

CKINVDCx12_ASAP7_75t_R g121 ( 
.A(n_79),
.Y(n_121)
);

NAND3xp33_ASAP7_75t_L g216 ( 
.A(n_121),
.B(n_119),
.C(n_149),
.Y(n_216)
);

OAI22xp5_ASAP7_75t_L g124 ( 
.A1(n_56),
.A2(n_52),
.B1(n_50),
.B2(n_48),
.Y(n_124)
);

AOI22xp5_ASAP7_75t_L g223 ( 
.A1(n_124),
.A2(n_133),
.B1(n_168),
.B2(n_127),
.Y(n_223)
);

AOI22xp33_ASAP7_75t_SL g125 ( 
.A1(n_97),
.A2(n_39),
.B1(n_51),
.B2(n_37),
.Y(n_125)
);

AOI22xp33_ASAP7_75t_SL g186 ( 
.A1(n_125),
.A2(n_138),
.B1(n_171),
.B2(n_88),
.Y(n_186)
);

CKINVDCx20_ASAP7_75t_R g132 ( 
.A(n_64),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_L g180 ( 
.A(n_132),
.B(n_137),
.Y(n_180)
);

OAI22xp5_ASAP7_75t_SL g133 ( 
.A1(n_65),
.A2(n_39),
.B1(n_32),
.B2(n_52),
.Y(n_133)
);

CKINVDCx20_ASAP7_75t_R g137 ( 
.A(n_78),
.Y(n_137)
);

AOI22xp33_ASAP7_75t_SL g138 ( 
.A1(n_84),
.A2(n_32),
.B1(n_48),
.B2(n_46),
.Y(n_138)
);

AOI22xp33_ASAP7_75t_L g139 ( 
.A1(n_69),
.A2(n_34),
.B1(n_27),
.B2(n_50),
.Y(n_139)
);

OAI22xp5_ASAP7_75t_L g178 ( 
.A1(n_139),
.A2(n_77),
.B1(n_72),
.B2(n_89),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_L g140 ( 
.A(n_57),
.B(n_34),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_L g181 ( 
.A(n_140),
.B(n_142),
.Y(n_181)
);

CKINVDCx20_ASAP7_75t_R g141 ( 
.A(n_74),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_L g187 ( 
.A(n_141),
.B(n_146),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_L g142 ( 
.A(n_90),
.B(n_27),
.Y(n_142)
);

CKINVDCx20_ASAP7_75t_R g146 ( 
.A(n_74),
.Y(n_146)
);

AND2x2_ASAP7_75t_SL g149 ( 
.A(n_61),
.B(n_1),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_L g155 ( 
.A(n_110),
.B(n_31),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_L g217 ( 
.A(n_155),
.B(n_159),
.Y(n_217)
);

NAND2xp5_ASAP7_75t_L g159 ( 
.A(n_112),
.B(n_33),
.Y(n_159)
);

CKINVDCx20_ASAP7_75t_R g164 ( 
.A(n_75),
.Y(n_164)
);

NOR2xp33_ASAP7_75t_L g188 ( 
.A(n_164),
.B(n_88),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_L g165 ( 
.A(n_107),
.B(n_33),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_L g229 ( 
.A(n_165),
.B(n_167),
.Y(n_229)
);

OAI22xp33_ASAP7_75t_SL g168 ( 
.A1(n_92),
.A2(n_41),
.B1(n_44),
.B2(n_46),
.Y(n_168)
);

AOI22xp33_ASAP7_75t_SL g171 ( 
.A1(n_62),
.A2(n_41),
.B1(n_44),
.B2(n_1),
.Y(n_171)
);

AOI22xp5_ASAP7_75t_L g250 ( 
.A1(n_178),
.A2(n_196),
.B1(n_220),
.B2(n_232),
.Y(n_250)
);

BUFx6f_ASAP7_75t_L g179 ( 
.A(n_130),
.Y(n_179)
);

INVx5_ASAP7_75t_L g238 ( 
.A(n_179),
.Y(n_238)
);

CKINVDCx20_ASAP7_75t_R g182 ( 
.A(n_129),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_L g266 ( 
.A(n_182),
.B(n_199),
.Y(n_266)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_120),
.Y(n_183)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_183),
.Y(n_240)
);

INVx2_ASAP7_75t_L g184 ( 
.A(n_135),
.Y(n_184)
);

INVx2_ASAP7_75t_L g237 ( 
.A(n_184),
.Y(n_237)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_126),
.Y(n_185)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_185),
.Y(n_248)
);

INVxp67_ASAP7_75t_L g239 ( 
.A(n_186),
.Y(n_239)
);

NOR2xp33_ASAP7_75t_L g236 ( 
.A(n_188),
.B(n_210),
.Y(n_236)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_155),
.Y(n_189)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_189),
.Y(n_249)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_159),
.Y(n_190)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_190),
.Y(n_252)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_157),
.Y(n_191)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_191),
.Y(n_254)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_158),
.Y(n_192)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_192),
.Y(n_260)
);

NAND2xp5_ASAP7_75t_SL g193 ( 
.A(n_162),
.B(n_93),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_SL g243 ( 
.A(n_193),
.B(n_197),
.Y(n_243)
);

XOR2xp5_ASAP7_75t_L g264 ( 
.A(n_194),
.B(n_174),
.Y(n_264)
);

INVx2_ASAP7_75t_SL g195 ( 
.A(n_145),
.Y(n_195)
);

INVx2_ASAP7_75t_L g244 ( 
.A(n_195),
.Y(n_244)
);

OAI22xp5_ASAP7_75t_SL g196 ( 
.A1(n_117),
.A2(n_98),
.B1(n_101),
.B2(n_93),
.Y(n_196)
);

NAND2xp5_ASAP7_75t_SL g197 ( 
.A(n_148),
.B(n_89),
.Y(n_197)
);

INVx2_ASAP7_75t_L g198 ( 
.A(n_135),
.Y(n_198)
);

INVx3_ASAP7_75t_L g246 ( 
.A(n_198),
.Y(n_246)
);

NOR2xp33_ASAP7_75t_L g199 ( 
.A(n_123),
.B(n_98),
.Y(n_199)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_172),
.Y(n_200)
);

INVxp67_ASAP7_75t_L g251 ( 
.A(n_200),
.Y(n_251)
);

NOR2xp33_ASAP7_75t_L g202 ( 
.A(n_136),
.B(n_101),
.Y(n_202)
);

NAND2xp5_ASAP7_75t_SL g245 ( 
.A(n_202),
.B(n_205),
.Y(n_245)
);

AND2x2_ASAP7_75t_L g203 ( 
.A(n_149),
.B(n_2),
.Y(n_203)
);

MAJIxp5_ASAP7_75t_L g255 ( 
.A(n_203),
.B(n_206),
.C(n_222),
.Y(n_255)
);

BUFx6f_ASAP7_75t_L g204 ( 
.A(n_130),
.Y(n_204)
);

INVx5_ASAP7_75t_L g267 ( 
.A(n_204),
.Y(n_267)
);

NAND2xp5_ASAP7_75t_SL g205 ( 
.A(n_177),
.B(n_2),
.Y(n_205)
);

OAI21xp5_ASAP7_75t_SL g206 ( 
.A1(n_142),
.A2(n_140),
.B(n_165),
.Y(n_206)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_176),
.Y(n_207)
);

INVxp67_ASAP7_75t_L g262 ( 
.A(n_207),
.Y(n_262)
);

NAND2xp5_ASAP7_75t_SL g208 ( 
.A(n_161),
.B(n_156),
.Y(n_208)
);

NAND2xp5_ASAP7_75t_SL g247 ( 
.A(n_208),
.B(n_209),
.Y(n_247)
);

NOR2xp33_ASAP7_75t_L g209 ( 
.A(n_144),
.B(n_116),
.Y(n_209)
);

NAND2xp5_ASAP7_75t_SL g210 ( 
.A(n_170),
.B(n_154),
.Y(n_210)
);

NOR2xp33_ASAP7_75t_L g211 ( 
.A(n_147),
.B(n_114),
.Y(n_211)
);

NOR2xp33_ASAP7_75t_L g242 ( 
.A(n_211),
.B(n_213),
.Y(n_242)
);

BUFx2_ASAP7_75t_L g212 ( 
.A(n_175),
.Y(n_212)
);

INVx3_ASAP7_75t_L g269 ( 
.A(n_212),
.Y(n_269)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_134),
.Y(n_213)
);

NOR2xp33_ASAP7_75t_L g214 ( 
.A(n_114),
.B(n_154),
.Y(n_214)
);

NOR2xp33_ASAP7_75t_L g258 ( 
.A(n_214),
.B(n_216),
.Y(n_258)
);

INVx6_ASAP7_75t_L g215 ( 
.A(n_151),
.Y(n_215)
);

BUFx5_ASAP7_75t_L g234 ( 
.A(n_215),
.Y(n_234)
);

BUFx2_ASAP7_75t_L g218 ( 
.A(n_175),
.Y(n_218)
);

NOR2xp33_ASAP7_75t_L g263 ( 
.A(n_218),
.B(n_221),
.Y(n_263)
);

BUFx2_ASAP7_75t_SL g219 ( 
.A(n_163),
.Y(n_219)
);

AOI22xp33_ASAP7_75t_SL g253 ( 
.A1(n_219),
.A2(n_228),
.B1(n_231),
.B2(n_163),
.Y(n_253)
);

OAI22xp33_ASAP7_75t_SL g220 ( 
.A1(n_151),
.A2(n_160),
.B1(n_173),
.B2(n_133),
.Y(n_220)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_134),
.Y(n_221)
);

XOR2xp5_ASAP7_75t_L g222 ( 
.A(n_128),
.B(n_166),
.Y(n_222)
);

OAI22xp5_ASAP7_75t_L g261 ( 
.A1(n_223),
.A2(n_174),
.B1(n_190),
.B2(n_217),
.Y(n_261)
);

INVx3_ASAP7_75t_L g224 ( 
.A(n_115),
.Y(n_224)
);

NOR2xp33_ASAP7_75t_L g271 ( 
.A(n_224),
.B(n_226),
.Y(n_271)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_152),
.Y(n_226)
);

AND2x2_ASAP7_75t_L g227 ( 
.A(n_128),
.B(n_152),
.Y(n_227)
);

MAJIxp5_ASAP7_75t_L g259 ( 
.A(n_227),
.B(n_167),
.C(n_143),
.Y(n_259)
);

BUFx6f_ASAP7_75t_L g228 ( 
.A(n_160),
.Y(n_228)
);

NAND2xp5_ASAP7_75t_L g233 ( 
.A(n_229),
.B(n_230),
.Y(n_233)
);

NAND2xp5_ASAP7_75t_L g230 ( 
.A(n_173),
.B(n_131),
.Y(n_230)
);

BUFx5_ASAP7_75t_L g231 ( 
.A(n_122),
.Y(n_231)
);

OAI22xp5_ASAP7_75t_L g232 ( 
.A1(n_113),
.A2(n_153),
.B1(n_169),
.B2(n_131),
.Y(n_232)
);

OA22x2_ASAP7_75t_L g235 ( 
.A1(n_223),
.A2(n_113),
.B1(n_150),
.B2(n_153),
.Y(n_235)
);

OA21x2_ASAP7_75t_L g301 ( 
.A1(n_235),
.A2(n_250),
.B(n_237),
.Y(n_301)
);

NAND2xp5_ASAP7_75t_L g241 ( 
.A(n_217),
.B(n_169),
.Y(n_241)
);

NAND2xp5_ASAP7_75t_L g278 ( 
.A(n_241),
.B(n_268),
.Y(n_278)
);

INVxp67_ASAP7_75t_L g283 ( 
.A(n_253),
.Y(n_283)
);

OAI21xp5_ASAP7_75t_L g256 ( 
.A1(n_206),
.A2(n_167),
.B(n_150),
.Y(n_256)
);

AOI21xp5_ASAP7_75t_L g289 ( 
.A1(n_256),
.A2(n_268),
.B(n_241),
.Y(n_289)
);

OAI22xp33_ASAP7_75t_SL g257 ( 
.A1(n_189),
.A2(n_143),
.B1(n_115),
.B2(n_122),
.Y(n_257)
);

AOI22xp5_ASAP7_75t_L g282 ( 
.A1(n_257),
.A2(n_261),
.B1(n_215),
.B2(n_228),
.Y(n_282)
);

XNOR2xp5_ASAP7_75t_L g304 ( 
.A(n_259),
.B(n_264),
.Y(n_304)
);

AOI22xp5_ASAP7_75t_L g265 ( 
.A1(n_225),
.A2(n_201),
.B1(n_229),
.B2(n_196),
.Y(n_265)
);

OAI22xp5_ASAP7_75t_L g280 ( 
.A1(n_265),
.A2(n_272),
.B1(n_212),
.B2(n_218),
.Y(n_280)
);

NAND2xp5_ASAP7_75t_L g268 ( 
.A(n_181),
.B(n_174),
.Y(n_268)
);

A2O1A1O1Ixp25_ASAP7_75t_L g270 ( 
.A1(n_181),
.A2(n_201),
.B(n_203),
.C(n_222),
.D(n_180),
.Y(n_270)
);

OAI21xp5_ASAP7_75t_SL g274 ( 
.A1(n_270),
.A2(n_187),
.B(n_230),
.Y(n_274)
);

AOI22xp33_ASAP7_75t_L g272 ( 
.A1(n_201),
.A2(n_225),
.B1(n_227),
.B2(n_200),
.Y(n_272)
);

NAND2xp5_ASAP7_75t_L g273 ( 
.A(n_203),
.B(n_194),
.Y(n_273)
);

NAND2xp5_ASAP7_75t_L g290 ( 
.A(n_273),
.B(n_233),
.Y(n_290)
);

A2O1A1O1Ixp25_ASAP7_75t_L g310 ( 
.A1(n_274),
.A2(n_299),
.B(n_246),
.C(n_234),
.D(n_238),
.Y(n_310)
);

XOR2x2_ASAP7_75t_L g275 ( 
.A(n_255),
.B(n_264),
.Y(n_275)
);

XNOR2xp5_ASAP7_75t_L g318 ( 
.A(n_275),
.B(n_290),
.Y(n_318)
);

MAJIxp5_ASAP7_75t_L g276 ( 
.A(n_255),
.B(n_227),
.C(n_195),
.Y(n_276)
);

MAJIxp5_ASAP7_75t_L g316 ( 
.A(n_276),
.B(n_291),
.C(n_298),
.Y(n_316)
);

A2O1A1Ixp33_ASAP7_75t_L g277 ( 
.A1(n_233),
.A2(n_184),
.B(n_198),
.C(n_224),
.Y(n_277)
);

NAND2xp5_ASAP7_75t_L g315 ( 
.A(n_277),
.B(n_280),
.Y(n_315)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_244),
.Y(n_279)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_279),
.Y(n_307)
);

CKINVDCx20_ASAP7_75t_R g281 ( 
.A(n_263),
.Y(n_281)
);

NOR2xp33_ASAP7_75t_L g305 ( 
.A(n_281),
.B(n_285),
.Y(n_305)
);

INVx1_ASAP7_75t_SL g306 ( 
.A(n_282),
.Y(n_306)
);

OAI22xp5_ASAP7_75t_SL g284 ( 
.A1(n_265),
.A2(n_179),
.B1(n_204),
.B2(n_231),
.Y(n_284)
);

OAI22xp5_ASAP7_75t_SL g313 ( 
.A1(n_284),
.A2(n_286),
.B1(n_238),
.B2(n_267),
.Y(n_313)
);

CKINVDCx20_ASAP7_75t_R g285 ( 
.A(n_271),
.Y(n_285)
);

AOI22xp33_ASAP7_75t_L g286 ( 
.A1(n_239),
.A2(n_235),
.B1(n_252),
.B2(n_249),
.Y(n_286)
);

NOR2xp33_ASAP7_75t_L g287 ( 
.A(n_247),
.B(n_266),
.Y(n_287)
);

NAND2xp5_ASAP7_75t_SL g309 ( 
.A(n_287),
.B(n_288),
.Y(n_309)
);

INVxp67_ASAP7_75t_L g288 ( 
.A(n_236),
.Y(n_288)
);

A2O1A1Ixp33_ASAP7_75t_SL g321 ( 
.A1(n_289),
.A2(n_300),
.B(n_301),
.C(n_280),
.Y(n_321)
);

XOR2xp5_ASAP7_75t_L g291 ( 
.A(n_273),
.B(n_270),
.Y(n_291)
);

INVx1_ASAP7_75t_SL g292 ( 
.A(n_244),
.Y(n_292)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_292),
.Y(n_314)
);

OR2x2_ASAP7_75t_L g293 ( 
.A(n_259),
.B(n_256),
.Y(n_293)
);

OAI21xp5_ASAP7_75t_L g308 ( 
.A1(n_293),
.A2(n_296),
.B(n_303),
.Y(n_308)
);

NOR2xp33_ASAP7_75t_L g294 ( 
.A(n_243),
.B(n_245),
.Y(n_294)
);

NAND2xp5_ASAP7_75t_SL g311 ( 
.A(n_294),
.B(n_297),
.Y(n_311)
);

CKINVDCx20_ASAP7_75t_R g295 ( 
.A(n_242),
.Y(n_295)
);

NOR2xp33_ASAP7_75t_L g312 ( 
.A(n_295),
.B(n_302),
.Y(n_312)
);

OR2x2_ASAP7_75t_L g296 ( 
.A(n_250),
.B(n_235),
.Y(n_296)
);

NOR2xp33_ASAP7_75t_L g297 ( 
.A(n_251),
.B(n_248),
.Y(n_297)
);

MAJIxp5_ASAP7_75t_L g298 ( 
.A(n_258),
.B(n_240),
.C(n_260),
.Y(n_298)
);

NAND2xp5_ASAP7_75t_L g299 ( 
.A(n_251),
.B(n_235),
.Y(n_299)
);

INVx13_ASAP7_75t_L g300 ( 
.A(n_269),
.Y(n_300)
);

OAI32xp33_ASAP7_75t_L g302 ( 
.A1(n_254),
.A2(n_239),
.A3(n_237),
.B1(n_262),
.B2(n_269),
.Y(n_302)
);

OAI21xp5_ASAP7_75t_SL g303 ( 
.A1(n_262),
.A2(n_246),
.B(n_234),
.Y(n_303)
);

NAND2xp5_ASAP7_75t_SL g333 ( 
.A(n_310),
.B(n_317),
.Y(n_333)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_313),
.Y(n_335)
);

NOR2xp33_ASAP7_75t_L g317 ( 
.A(n_295),
.B(n_267),
.Y(n_317)
);

MAJIxp5_ASAP7_75t_L g319 ( 
.A(n_275),
.B(n_304),
.C(n_291),
.Y(n_319)
);

MAJIxp5_ASAP7_75t_L g328 ( 
.A(n_319),
.B(n_326),
.C(n_293),
.Y(n_328)
);

NOR2xp33_ASAP7_75t_L g320 ( 
.A(n_285),
.B(n_281),
.Y(n_320)
);

NAND2xp5_ASAP7_75t_SL g339 ( 
.A(n_320),
.B(n_324),
.Y(n_339)
);

A2O1A1Ixp33_ASAP7_75t_SL g342 ( 
.A1(n_321),
.A2(n_301),
.B(n_300),
.C(n_292),
.Y(n_342)
);

OAI32xp33_ASAP7_75t_L g322 ( 
.A1(n_278),
.A2(n_299),
.A3(n_290),
.B1(n_277),
.B2(n_287),
.Y(n_322)
);

NOR2xp33_ASAP7_75t_L g330 ( 
.A(n_322),
.B(n_325),
.Y(n_330)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_279),
.Y(n_323)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_323),
.Y(n_336)
);

NOR2xp33_ASAP7_75t_L g324 ( 
.A(n_298),
.B(n_274),
.Y(n_324)
);

BUFx6f_ASAP7_75t_L g325 ( 
.A(n_300),
.Y(n_325)
);

XOR2xp5_ASAP7_75t_L g326 ( 
.A(n_275),
.B(n_304),
.Y(n_326)
);

NOR2x1_ASAP7_75t_L g327 ( 
.A(n_308),
.B(n_315),
.Y(n_327)
);

NOR2xp33_ASAP7_75t_L g350 ( 
.A(n_327),
.B(n_329),
.Y(n_350)
);

MAJIxp5_ASAP7_75t_L g343 ( 
.A(n_328),
.B(n_340),
.C(n_341),
.Y(n_343)
);

OAI21xp5_ASAP7_75t_L g329 ( 
.A1(n_308),
.A2(n_293),
.B(n_289),
.Y(n_329)
);

AOI21xp5_ASAP7_75t_L g331 ( 
.A1(n_312),
.A2(n_283),
.B(n_303),
.Y(n_331)
);

NOR2xp33_ASAP7_75t_L g351 ( 
.A(n_331),
.B(n_334),
.Y(n_351)
);

NOR2xp33_ASAP7_75t_L g332 ( 
.A(n_311),
.B(n_278),
.Y(n_332)
);

NOR2xp33_ASAP7_75t_SL g345 ( 
.A(n_332),
.B(n_337),
.Y(n_345)
);

CKINVDCx20_ASAP7_75t_R g334 ( 
.A(n_305),
.Y(n_334)
);

NOR2xp33_ASAP7_75t_L g337 ( 
.A(n_309),
.B(n_297),
.Y(n_337)
);

OAI322xp33_ASAP7_75t_L g338 ( 
.A1(n_326),
.A2(n_276),
.A3(n_302),
.B1(n_301),
.B2(n_282),
.C1(n_296),
.C2(n_284),
.Y(n_338)
);

XNOR2xp5_ASAP7_75t_SL g352 ( 
.A(n_338),
.B(n_310),
.Y(n_352)
);

MAJIxp5_ASAP7_75t_L g340 ( 
.A(n_319),
.B(n_316),
.C(n_318),
.Y(n_340)
);

XOR2xp5_ASAP7_75t_L g341 ( 
.A(n_318),
.B(n_296),
.Y(n_341)
);

AOI22xp5_ASAP7_75t_L g348 ( 
.A1(n_342),
.A2(n_301),
.B1(n_315),
.B2(n_321),
.Y(n_348)
);

CKINVDCx20_ASAP7_75t_R g344 ( 
.A(n_334),
.Y(n_344)
);

NAND2xp5_ASAP7_75t_L g364 ( 
.A(n_344),
.B(n_347),
.Y(n_364)
);

MAJIxp5_ASAP7_75t_L g346 ( 
.A(n_328),
.B(n_316),
.C(n_321),
.Y(n_346)
);

MAJIxp5_ASAP7_75t_L g359 ( 
.A(n_346),
.B(n_354),
.C(n_329),
.Y(n_359)
);

BUFx2_ASAP7_75t_L g347 ( 
.A(n_335),
.Y(n_347)
);

OAI21xp5_ASAP7_75t_SL g362 ( 
.A1(n_348),
.A2(n_327),
.B(n_342),
.Y(n_362)
);

AOI22xp5_ASAP7_75t_L g349 ( 
.A1(n_335),
.A2(n_306),
.B1(n_313),
.B2(n_321),
.Y(n_349)
);

AND2x2_ASAP7_75t_L g356 ( 
.A(n_349),
.B(n_342),
.Y(n_356)
);

NAND2xp5_ASAP7_75t_SL g355 ( 
.A(n_352),
.B(n_341),
.Y(n_355)
);

INVx2_ASAP7_75t_L g353 ( 
.A(n_336),
.Y(n_353)
);

INVx1_ASAP7_75t_L g358 ( 
.A(n_353),
.Y(n_358)
);

XNOR2xp5_ASAP7_75t_L g354 ( 
.A(n_340),
.B(n_322),
.Y(n_354)
);

XOR2xp5_ASAP7_75t_L g366 ( 
.A(n_355),
.B(n_362),
.Y(n_366)
);

NAND2xp5_ASAP7_75t_L g369 ( 
.A(n_356),
.B(n_357),
.Y(n_369)
);

AOI21xp5_ASAP7_75t_L g357 ( 
.A1(n_350),
.A2(n_330),
.B(n_333),
.Y(n_357)
);

MAJIxp5_ASAP7_75t_L g365 ( 
.A(n_359),
.B(n_361),
.C(n_343),
.Y(n_365)
);

NAND2xp5_ASAP7_75t_SL g360 ( 
.A(n_351),
.B(n_339),
.Y(n_360)
);

NOR2xp33_ASAP7_75t_SL g371 ( 
.A(n_360),
.B(n_345),
.Y(n_371)
);

MAJIxp5_ASAP7_75t_L g361 ( 
.A(n_343),
.B(n_339),
.C(n_333),
.Y(n_361)
);

INVx1_ASAP7_75t_L g363 ( 
.A(n_353),
.Y(n_363)
);

OR2x2_ASAP7_75t_L g367 ( 
.A(n_363),
.B(n_325),
.Y(n_367)
);

XNOR2xp5_ASAP7_75t_L g374 ( 
.A(n_365),
.B(n_368),
.Y(n_374)
);

NAND2xp5_ASAP7_75t_L g372 ( 
.A(n_367),
.B(n_370),
.Y(n_372)
);

MAJIxp5_ASAP7_75t_L g368 ( 
.A(n_361),
.B(n_346),
.C(n_354),
.Y(n_368)
);

MAJIxp5_ASAP7_75t_L g370 ( 
.A(n_359),
.B(n_352),
.C(n_331),
.Y(n_370)
);

OAI21xp5_ASAP7_75t_L g373 ( 
.A1(n_371),
.A2(n_357),
.B(n_364),
.Y(n_373)
);

NAND2xp5_ASAP7_75t_SL g378 ( 
.A(n_373),
.B(n_375),
.Y(n_378)
);

NAND2xp5_ASAP7_75t_L g375 ( 
.A(n_369),
.B(n_358),
.Y(n_375)
);

NAND2xp33_ASAP7_75t_SL g376 ( 
.A(n_366),
.B(n_348),
.Y(n_376)
);

AOI21xp5_ASAP7_75t_L g380 ( 
.A1(n_376),
.A2(n_362),
.B(n_356),
.Y(n_380)
);

XNOR2xp5_ASAP7_75t_L g377 ( 
.A(n_374),
.B(n_327),
.Y(n_377)
);

NAND2xp5_ASAP7_75t_L g383 ( 
.A(n_377),
.B(n_379),
.Y(n_383)
);

NOR2xp33_ASAP7_75t_L g379 ( 
.A(n_372),
.B(n_371),
.Y(n_379)
);

OAI21x1_ASAP7_75t_L g381 ( 
.A1(n_380),
.A2(n_376),
.B(n_342),
.Y(n_381)
);

OAI221xp5_ASAP7_75t_L g385 ( 
.A1(n_381),
.A2(n_382),
.B1(n_349),
.B2(n_314),
.C(n_307),
.Y(n_385)
);

A2O1A1O1Ixp25_ASAP7_75t_L g382 ( 
.A1(n_378),
.A2(n_342),
.B(n_336),
.C(n_347),
.D(n_323),
.Y(n_382)
);

BUFx24_ASAP7_75t_SL g384 ( 
.A(n_383),
.Y(n_384)
);

OAI21xp5_ASAP7_75t_L g386 ( 
.A1(n_384),
.A2(n_385),
.B(n_314),
.Y(n_386)
);

XOR2xp5_ASAP7_75t_L g387 ( 
.A(n_386),
.B(n_306),
.Y(n_387)
);


endmodule