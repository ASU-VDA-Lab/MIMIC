module fake_ariane_455_n_908 (n_83, n_8, n_56, n_60, n_170, n_190, n_160, n_64, n_179, n_180, n_119, n_124, n_167, n_90, n_195, n_38, n_47, n_110, n_153, n_18, n_197, n_86, n_75, n_89, n_67, n_176, n_149, n_34, n_158, n_172, n_69, n_95, n_175, n_92, n_143, n_183, n_150, n_98, n_74, n_113, n_114, n_33, n_19, n_40, n_181, n_152, n_120, n_169, n_106, n_12, n_53, n_173, n_111, n_21, n_115, n_133, n_66, n_71, n_24, n_7, n_109, n_96, n_156, n_49, n_20, n_174, n_100, n_17, n_50, n_187, n_132, n_62, n_147, n_51, n_166, n_76, n_103, n_79, n_26, n_3, n_46, n_0, n_84, n_36, n_199, n_91, n_159, n_107, n_189, n_72, n_105, n_128, n_44, n_30, n_82, n_178, n_31, n_42, n_57, n_131, n_70, n_10, n_117, n_139, n_165, n_85, n_130, n_144, n_6, n_48, n_94, n_101, n_4, n_134, n_188, n_185, n_2, n_32, n_37, n_58, n_65, n_123, n_9, n_138, n_112, n_45, n_162, n_11, n_129, n_126, n_137, n_122, n_198, n_148, n_164, n_52, n_157, n_184, n_177, n_135, n_73, n_77, n_171, n_15, n_118, n_93, n_121, n_23, n_61, n_108, n_102, n_182, n_196, n_125, n_22, n_168, n_43, n_1, n_81, n_87, n_13, n_27, n_29, n_41, n_140, n_55, n_191, n_151, n_136, n_192, n_28, n_80, n_146, n_194, n_97, n_154, n_142, n_161, n_14, n_163, n_88, n_186, n_141, n_68, n_116, n_104, n_145, n_78, n_193, n_39, n_59, n_63, n_99, n_16, n_5, n_155, n_127, n_35, n_54, n_25, n_908);

input n_83;
input n_8;
input n_56;
input n_60;
input n_170;
input n_190;
input n_160;
input n_64;
input n_179;
input n_180;
input n_119;
input n_124;
input n_167;
input n_90;
input n_195;
input n_38;
input n_47;
input n_110;
input n_153;
input n_18;
input n_197;
input n_86;
input n_75;
input n_89;
input n_67;
input n_176;
input n_149;
input n_34;
input n_158;
input n_172;
input n_69;
input n_95;
input n_175;
input n_92;
input n_143;
input n_183;
input n_150;
input n_98;
input n_74;
input n_113;
input n_114;
input n_33;
input n_19;
input n_40;
input n_181;
input n_152;
input n_120;
input n_169;
input n_106;
input n_12;
input n_53;
input n_173;
input n_111;
input n_21;
input n_115;
input n_133;
input n_66;
input n_71;
input n_24;
input n_7;
input n_109;
input n_96;
input n_156;
input n_49;
input n_20;
input n_174;
input n_100;
input n_17;
input n_50;
input n_187;
input n_132;
input n_62;
input n_147;
input n_51;
input n_166;
input n_76;
input n_103;
input n_79;
input n_26;
input n_3;
input n_46;
input n_0;
input n_84;
input n_36;
input n_199;
input n_91;
input n_159;
input n_107;
input n_189;
input n_72;
input n_105;
input n_128;
input n_44;
input n_30;
input n_82;
input n_178;
input n_31;
input n_42;
input n_57;
input n_131;
input n_70;
input n_10;
input n_117;
input n_139;
input n_165;
input n_85;
input n_130;
input n_144;
input n_6;
input n_48;
input n_94;
input n_101;
input n_4;
input n_134;
input n_188;
input n_185;
input n_2;
input n_32;
input n_37;
input n_58;
input n_65;
input n_123;
input n_9;
input n_138;
input n_112;
input n_45;
input n_162;
input n_11;
input n_129;
input n_126;
input n_137;
input n_122;
input n_198;
input n_148;
input n_164;
input n_52;
input n_157;
input n_184;
input n_177;
input n_135;
input n_73;
input n_77;
input n_171;
input n_15;
input n_118;
input n_93;
input n_121;
input n_23;
input n_61;
input n_108;
input n_102;
input n_182;
input n_196;
input n_125;
input n_22;
input n_168;
input n_43;
input n_1;
input n_81;
input n_87;
input n_13;
input n_27;
input n_29;
input n_41;
input n_140;
input n_55;
input n_191;
input n_151;
input n_136;
input n_192;
input n_28;
input n_80;
input n_146;
input n_194;
input n_97;
input n_154;
input n_142;
input n_161;
input n_14;
input n_163;
input n_88;
input n_186;
input n_141;
input n_68;
input n_116;
input n_104;
input n_145;
input n_78;
input n_193;
input n_39;
input n_59;
input n_63;
input n_99;
input n_16;
input n_5;
input n_155;
input n_127;
input n_35;
input n_54;
input n_25;

output n_908;

wire n_295;
wire n_356;
wire n_556;
wire n_698;
wire n_695;
wire n_730;
wire n_386;
wire n_307;
wire n_516;
wire n_589;
wire n_332;
wire n_581;
wire n_294;
wire n_646;
wire n_640;
wire n_463;
wire n_830;
wire n_691;
wire n_404;
wire n_678;
wire n_651;
wire n_347;
wire n_423;
wire n_469;
wire n_479;
wire n_726;
wire n_603;
wire n_878;
wire n_373;
wire n_299;
wire n_836;
wire n_541;
wire n_499;
wire n_789;
wire n_788;
wire n_850;
wire n_771;
wire n_564;
wire n_610;
wire n_205;
wire n_752;
wire n_341;
wire n_245;
wire n_421;
wire n_549;
wire n_522;
wire n_319;
wire n_591;
wire n_760;
wire n_690;
wire n_906;
wire n_416;
wire n_283;
wire n_525;
wire n_806;
wire n_367;
wire n_713;
wire n_649;
wire n_598;
wire n_345;
wire n_374;
wire n_318;
wire n_817;
wire n_244;
wire n_643;
wire n_679;
wire n_226;
wire n_781;
wire n_220;
wire n_261;
wire n_682;
wire n_663;
wire n_370;
wire n_706;
wire n_717;
wire n_819;
wire n_286;
wire n_443;
wire n_586;
wire n_864;
wire n_686;
wire n_605;
wire n_776;
wire n_424;
wire n_528;
wire n_584;
wire n_387;
wire n_406;
wire n_826;
wire n_524;
wire n_634;
wire n_391;
wire n_349;
wire n_756;
wire n_466;
wire n_346;
wire n_214;
wire n_764;
wire n_348;
wire n_552;
wire n_462;
wire n_607;
wire n_670;
wire n_897;
wire n_410;
wire n_379;
wire n_445;
wire n_515;
wire n_807;
wire n_765;
wire n_264;
wire n_891;
wire n_737;
wire n_885;
wire n_232;
wire n_441;
wire n_568;
wire n_385;
wire n_637;
wire n_327;
wire n_766;
wire n_372;
wire n_377;
wire n_396;
wire n_802;
wire n_631;
wire n_399;
wire n_554;
wire n_520;
wire n_870;
wire n_714;
wire n_279;
wire n_905;
wire n_702;
wire n_207;
wire n_857;
wire n_790;
wire n_898;
wire n_363;
wire n_720;
wire n_354;
wire n_813;
wire n_725;
wire n_419;
wire n_230;
wire n_270;
wire n_633;
wire n_900;
wire n_883;
wire n_338;
wire n_285;
wire n_473;
wire n_801;
wire n_202;
wire n_733;
wire n_761;
wire n_818;
wire n_500;
wire n_665;
wire n_336;
wire n_731;
wire n_779;
wire n_754;
wire n_871;
wire n_315;
wire n_903;
wire n_594;
wire n_311;
wire n_239;
wire n_402;
wire n_272;
wire n_829;
wire n_668;
wire n_339;
wire n_758;
wire n_738;
wire n_833;
wire n_672;
wire n_487;
wire n_740;
wire n_879;
wire n_422;
wire n_648;
wire n_784;
wire n_269;
wire n_597;
wire n_816;
wire n_855;
wire n_259;
wire n_835;
wire n_808;
wire n_446;
wire n_553;
wire n_753;
wire n_566;
wire n_814;
wire n_578;
wire n_701;
wire n_625;
wire n_405;
wire n_557;
wire n_858;
wire n_242;
wire n_645;
wire n_309;
wire n_331;
wire n_320;
wire n_559;
wire n_401;
wire n_485;
wire n_267;
wire n_495;
wire n_504;
wire n_647;
wire n_483;
wire n_335;
wire n_435;
wire n_350;
wire n_291;
wire n_822;
wire n_381;
wire n_344;
wire n_795;
wire n_426;
wire n_433;
wire n_481;
wire n_600;
wire n_721;
wire n_840;
wire n_398;
wire n_210;
wire n_200;
wire n_529;
wire n_502;
wire n_253;
wire n_561;
wire n_770;
wire n_821;
wire n_218;
wire n_839;
wire n_271;
wire n_465;
wire n_507;
wire n_486;
wire n_901;
wire n_759;
wire n_247;
wire n_569;
wire n_567;
wire n_825;
wire n_732;
wire n_369;
wire n_240;
wire n_224;
wire n_787;
wire n_894;
wire n_547;
wire n_420;
wire n_562;
wire n_518;
wire n_439;
wire n_604;
wire n_677;
wire n_614;
wire n_222;
wire n_478;
wire n_703;
wire n_748;
wire n_786;
wire n_510;
wire n_831;
wire n_256;
wire n_868;
wire n_326;
wire n_681;
wire n_778;
wire n_227;
wire n_874;
wire n_323;
wire n_550;
wire n_635;
wire n_707;
wire n_330;
wire n_400;
wire n_689;
wire n_694;
wire n_884;
wire n_282;
wire n_328;
wire n_368;
wire n_699;
wire n_590;
wire n_727;
wire n_277;
wire n_248;
wire n_301;
wire n_467;
wire n_432;
wire n_545;
wire n_536;
wire n_644;
wire n_293;
wire n_823;
wire n_620;
wire n_228;
wire n_325;
wire n_276;
wire n_688;
wire n_859;
wire n_636;
wire n_427;
wire n_587;
wire n_497;
wire n_693;
wire n_863;
wire n_303;
wire n_671;
wire n_442;
wire n_777;
wire n_206;
wire n_352;
wire n_538;
wire n_899;
wire n_576;
wire n_843;
wire n_511;
wire n_611;
wire n_238;
wire n_365;
wire n_455;
wire n_429;
wire n_654;
wire n_588;
wire n_638;
wire n_334;
wire n_729;
wire n_887;
wire n_661;
wire n_488;
wire n_775;
wire n_667;
wire n_300;
wire n_533;
wire n_904;
wire n_505;
wire n_869;
wire n_846;
wire n_390;
wire n_498;
wire n_501;
wire n_438;
wire n_314;
wire n_684;
wire n_440;
wire n_627;
wire n_273;
wire n_305;
wire n_539;
wire n_312;
wire n_233;
wire n_728;
wire n_388;
wire n_333;
wire n_449;
wire n_612;
wire n_413;
wire n_392;
wire n_376;
wire n_512;
wire n_715;
wire n_889;
wire n_579;
wire n_844;
wire n_459;
wire n_685;
wire n_221;
wire n_321;
wire n_361;
wire n_458;
wire n_383;
wire n_623;
wire n_838;
wire n_237;
wire n_780;
wire n_861;
wire n_711;
wire n_877;
wire n_453;
wire n_734;
wire n_491;
wire n_810;
wire n_723;
wire n_616;
wire n_617;
wire n_658;
wire n_630;
wire n_705;
wire n_570;
wire n_260;
wire n_362;
wire n_543;
wire n_310;
wire n_709;
wire n_236;
wire n_601;
wire n_683;
wire n_565;
wire n_281;
wire n_628;
wire n_809;
wire n_461;
wire n_209;
wire n_262;
wire n_490;
wire n_743;
wire n_225;
wire n_907;
wire n_235;
wire n_881;
wire n_660;
wire n_464;
wire n_735;
wire n_575;
wire n_546;
wire n_297;
wire n_662;
wire n_641;
wire n_503;
wire n_700;
wire n_527;
wire n_290;
wire n_747;
wire n_741;
wire n_772;
wire n_847;
wire n_371;
wire n_845;
wire n_888;
wire n_639;
wire n_217;
wire n_452;
wire n_673;
wire n_676;
wire n_551;
wire n_308;
wire n_708;
wire n_417;
wire n_201;
wire n_572;
wire n_343;
wire n_865;
wire n_414;
wire n_571;
wire n_680;
wire n_287;
wire n_302;
wire n_380;
wire n_582;
wire n_284;
wire n_448;
wire n_593;
wire n_755;
wire n_710;
wire n_860;
wire n_249;
wire n_534;
wire n_355;
wire n_212;
wire n_444;
wire n_609;
wire n_278;
wire n_851;
wire n_255;
wire n_560;
wire n_450;
wire n_890;
wire n_257;
wire n_842;
wire n_652;
wire n_451;
wire n_613;
wire n_745;
wire n_475;
wire n_896;
wire n_409;
wire n_519;
wire n_902;
wire n_384;
wire n_468;
wire n_853;
wire n_526;
wire n_716;
wire n_742;
wire n_696;
wire n_674;
wire n_482;
wire n_316;
wire n_798;
wire n_769;
wire n_820;
wire n_577;
wire n_407;
wire n_774;
wire n_872;
wire n_254;
wire n_596;
wire n_476;
wire n_460;
wire n_219;
wire n_832;
wire n_535;
wire n_231;
wire n_366;
wire n_744;
wire n_762;
wire n_656;
wire n_555;
wire n_234;
wire n_492;
wire n_574;
wire n_848;
wire n_804;
wire n_280;
wire n_252;
wire n_215;
wire n_629;
wire n_664;
wire n_454;
wire n_298;
wire n_532;
wire n_415;
wire n_794;
wire n_763;
wire n_655;
wire n_544;
wire n_216;
wire n_540;
wire n_692;
wire n_599;
wire n_768;
wire n_514;
wire n_418;
wire n_537;
wire n_223;
wire n_403;
wire n_750;
wire n_834;
wire n_389;
wire n_800;
wire n_657;
wire n_513;
wire n_837;
wire n_288;
wire n_812;
wire n_395;
wire n_621;
wire n_606;
wire n_213;
wire n_862;
wire n_304;
wire n_895;
wire n_659;
wire n_509;
wire n_583;
wire n_724;
wire n_306;
wire n_666;
wire n_313;
wire n_430;
wire n_626;
wire n_493;
wire n_722;
wire n_203;
wire n_378;
wire n_436;
wire n_757;
wire n_375;
wire n_324;
wire n_585;
wire n_875;
wire n_669;
wire n_785;
wire n_827;
wire n_619;
wire n_337;
wire n_437;
wire n_274;
wire n_622;
wire n_697;
wire n_472;
wire n_296;
wire n_265;
wire n_746;
wire n_208;
wire n_456;
wire n_292;
wire n_880;
wire n_852;
wire n_793;
wire n_275;
wire n_704;
wire n_204;
wire n_751;
wire n_615;
wire n_521;
wire n_873;
wire n_496;
wire n_739;
wire n_342;
wire n_866;
wire n_246;
wire n_517;
wire n_530;
wire n_792;
wire n_824;
wire n_428;
wire n_358;
wire n_580;
wire n_892;
wire n_608;
wire n_494;
wire n_719;
wire n_263;
wire n_434;
wire n_360;
wire n_563;
wire n_229;
wire n_394;
wire n_250;
wire n_773;
wire n_882;
wire n_317;
wire n_867;
wire n_243;
wire n_803;
wire n_329;
wire n_718;
wire n_340;
wire n_749;
wire n_289;
wire n_548;
wire n_542;
wire n_815;
wire n_523;
wire n_268;
wire n_266;
wire n_470;
wire n_457;
wire n_632;
wire n_477;
wire n_364;
wire n_258;
wire n_650;
wire n_782;
wire n_856;
wire n_425;
wire n_431;
wire n_811;
wire n_508;
wire n_624;
wire n_791;
wire n_876;
wire n_618;
wire n_411;
wire n_484;
wire n_712;
wire n_849;
wire n_353;
wire n_736;
wire n_767;
wire n_241;
wire n_357;
wire n_412;
wire n_687;
wire n_447;
wire n_382;
wire n_797;
wire n_489;
wire n_480;
wire n_211;
wire n_642;
wire n_408;
wire n_828;
wire n_595;
wire n_322;
wire n_251;
wire n_506;
wire n_893;
wire n_602;
wire n_799;
wire n_558;
wire n_592;
wire n_397;
wire n_841;
wire n_854;
wire n_471;
wire n_351;
wire n_886;
wire n_393;
wire n_474;
wire n_653;
wire n_359;
wire n_573;
wire n_796;
wire n_805;
wire n_531;
wire n_783;
wire n_675;

CKINVDCx16_ASAP7_75t_R g200 ( 
.A(n_168),
.Y(n_200)
);

CKINVDCx5p33_ASAP7_75t_R g201 ( 
.A(n_33),
.Y(n_201)
);

CKINVDCx5p33_ASAP7_75t_R g202 ( 
.A(n_53),
.Y(n_202)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_60),
.Y(n_203)
);

BUFx2_ASAP7_75t_L g204 ( 
.A(n_157),
.Y(n_204)
);

INVx2_ASAP7_75t_SL g205 ( 
.A(n_181),
.Y(n_205)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_67),
.Y(n_206)
);

INVx1_ASAP7_75t_SL g207 ( 
.A(n_47),
.Y(n_207)
);

CKINVDCx5p33_ASAP7_75t_R g208 ( 
.A(n_193),
.Y(n_208)
);

CKINVDCx5p33_ASAP7_75t_R g209 ( 
.A(n_127),
.Y(n_209)
);

CKINVDCx20_ASAP7_75t_R g210 ( 
.A(n_174),
.Y(n_210)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_191),
.Y(n_211)
);

CKINVDCx5p33_ASAP7_75t_R g212 ( 
.A(n_173),
.Y(n_212)
);

CKINVDCx5p33_ASAP7_75t_R g213 ( 
.A(n_123),
.Y(n_213)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_21),
.Y(n_214)
);

CKINVDCx5p33_ASAP7_75t_R g215 ( 
.A(n_198),
.Y(n_215)
);

INVx2_ASAP7_75t_L g216 ( 
.A(n_29),
.Y(n_216)
);

CKINVDCx5p33_ASAP7_75t_R g217 ( 
.A(n_12),
.Y(n_217)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_86),
.Y(n_218)
);

CKINVDCx5p33_ASAP7_75t_R g219 ( 
.A(n_72),
.Y(n_219)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_84),
.Y(n_220)
);

CKINVDCx5p33_ASAP7_75t_R g221 ( 
.A(n_175),
.Y(n_221)
);

CKINVDCx5p33_ASAP7_75t_R g222 ( 
.A(n_137),
.Y(n_222)
);

CKINVDCx5p33_ASAP7_75t_R g223 ( 
.A(n_59),
.Y(n_223)
);

CKINVDCx5p33_ASAP7_75t_R g224 ( 
.A(n_143),
.Y(n_224)
);

BUFx6f_ASAP7_75t_L g225 ( 
.A(n_41),
.Y(n_225)
);

INVx2_ASAP7_75t_SL g226 ( 
.A(n_139),
.Y(n_226)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_113),
.Y(n_227)
);

INVx2_ASAP7_75t_SL g228 ( 
.A(n_76),
.Y(n_228)
);

CKINVDCx5p33_ASAP7_75t_R g229 ( 
.A(n_153),
.Y(n_229)
);

CKINVDCx5p33_ASAP7_75t_R g230 ( 
.A(n_5),
.Y(n_230)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_36),
.Y(n_231)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_70),
.Y(n_232)
);

CKINVDCx5p33_ASAP7_75t_R g233 ( 
.A(n_54),
.Y(n_233)
);

CKINVDCx5p33_ASAP7_75t_R g234 ( 
.A(n_21),
.Y(n_234)
);

CKINVDCx5p33_ASAP7_75t_R g235 ( 
.A(n_99),
.Y(n_235)
);

CKINVDCx5p33_ASAP7_75t_R g236 ( 
.A(n_11),
.Y(n_236)
);

CKINVDCx5p33_ASAP7_75t_R g237 ( 
.A(n_188),
.Y(n_237)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_23),
.Y(n_238)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_38),
.Y(n_239)
);

INVx2_ASAP7_75t_SL g240 ( 
.A(n_195),
.Y(n_240)
);

CKINVDCx5p33_ASAP7_75t_R g241 ( 
.A(n_176),
.Y(n_241)
);

CKINVDCx5p33_ASAP7_75t_R g242 ( 
.A(n_151),
.Y(n_242)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_75),
.Y(n_243)
);

CKINVDCx5p33_ASAP7_75t_R g244 ( 
.A(n_116),
.Y(n_244)
);

CKINVDCx5p33_ASAP7_75t_R g245 ( 
.A(n_39),
.Y(n_245)
);

BUFx3_ASAP7_75t_L g246 ( 
.A(n_18),
.Y(n_246)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_125),
.Y(n_247)
);

CKINVDCx5p33_ASAP7_75t_R g248 ( 
.A(n_122),
.Y(n_248)
);

CKINVDCx5p33_ASAP7_75t_R g249 ( 
.A(n_140),
.Y(n_249)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_138),
.Y(n_250)
);

CKINVDCx5p33_ASAP7_75t_R g251 ( 
.A(n_179),
.Y(n_251)
);

CKINVDCx5p33_ASAP7_75t_R g252 ( 
.A(n_57),
.Y(n_252)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_82),
.Y(n_253)
);

BUFx3_ASAP7_75t_L g254 ( 
.A(n_199),
.Y(n_254)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_196),
.Y(n_255)
);

CKINVDCx5p33_ASAP7_75t_R g256 ( 
.A(n_78),
.Y(n_256)
);

CKINVDCx5p33_ASAP7_75t_R g257 ( 
.A(n_144),
.Y(n_257)
);

CKINVDCx5p33_ASAP7_75t_R g258 ( 
.A(n_32),
.Y(n_258)
);

CKINVDCx20_ASAP7_75t_R g259 ( 
.A(n_128),
.Y(n_259)
);

CKINVDCx5p33_ASAP7_75t_R g260 ( 
.A(n_7),
.Y(n_260)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_158),
.Y(n_261)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_40),
.Y(n_262)
);

CKINVDCx5p33_ASAP7_75t_R g263 ( 
.A(n_190),
.Y(n_263)
);

INVx2_ASAP7_75t_SL g264 ( 
.A(n_50),
.Y(n_264)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_149),
.Y(n_265)
);

CKINVDCx5p33_ASAP7_75t_R g266 ( 
.A(n_109),
.Y(n_266)
);

CKINVDCx5p33_ASAP7_75t_R g267 ( 
.A(n_43),
.Y(n_267)
);

CKINVDCx5p33_ASAP7_75t_R g268 ( 
.A(n_169),
.Y(n_268)
);

CKINVDCx5p33_ASAP7_75t_R g269 ( 
.A(n_197),
.Y(n_269)
);

CKINVDCx5p33_ASAP7_75t_R g270 ( 
.A(n_189),
.Y(n_270)
);

CKINVDCx5p33_ASAP7_75t_R g271 ( 
.A(n_73),
.Y(n_271)
);

CKINVDCx5p33_ASAP7_75t_R g272 ( 
.A(n_10),
.Y(n_272)
);

CKINVDCx5p33_ASAP7_75t_R g273 ( 
.A(n_96),
.Y(n_273)
);

CKINVDCx5p33_ASAP7_75t_R g274 ( 
.A(n_0),
.Y(n_274)
);

INVx3_ASAP7_75t_L g275 ( 
.A(n_92),
.Y(n_275)
);

CKINVDCx20_ASAP7_75t_R g276 ( 
.A(n_63),
.Y(n_276)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_65),
.Y(n_277)
);

CKINVDCx14_ASAP7_75t_R g278 ( 
.A(n_26),
.Y(n_278)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_42),
.Y(n_279)
);

INVx2_ASAP7_75t_L g280 ( 
.A(n_27),
.Y(n_280)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_246),
.Y(n_281)
);

NAND2xp5_ASAP7_75t_L g282 ( 
.A(n_204),
.B(n_0),
.Y(n_282)
);

INVxp67_ASAP7_75t_L g283 ( 
.A(n_214),
.Y(n_283)
);

INVx2_ASAP7_75t_L g284 ( 
.A(n_254),
.Y(n_284)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_246),
.Y(n_285)
);

INVx3_ASAP7_75t_L g286 ( 
.A(n_238),
.Y(n_286)
);

INVx5_ASAP7_75t_L g287 ( 
.A(n_225),
.Y(n_287)
);

HB1xp67_ASAP7_75t_L g288 ( 
.A(n_274),
.Y(n_288)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_203),
.Y(n_289)
);

INVx5_ASAP7_75t_L g290 ( 
.A(n_225),
.Y(n_290)
);

CKINVDCx5p33_ASAP7_75t_R g291 ( 
.A(n_200),
.Y(n_291)
);

BUFx6f_ASAP7_75t_L g292 ( 
.A(n_225),
.Y(n_292)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_206),
.Y(n_293)
);

NAND2xp5_ASAP7_75t_SL g294 ( 
.A(n_216),
.B(n_1),
.Y(n_294)
);

BUFx3_ASAP7_75t_L g295 ( 
.A(n_254),
.Y(n_295)
);

INVx3_ASAP7_75t_L g296 ( 
.A(n_280),
.Y(n_296)
);

BUFx6f_ASAP7_75t_L g297 ( 
.A(n_225),
.Y(n_297)
);

AND2x2_ASAP7_75t_L g298 ( 
.A(n_278),
.B(n_1),
.Y(n_298)
);

INVx5_ASAP7_75t_L g299 ( 
.A(n_275),
.Y(n_299)
);

BUFx2_ASAP7_75t_L g300 ( 
.A(n_274),
.Y(n_300)
);

INVx5_ASAP7_75t_L g301 ( 
.A(n_275),
.Y(n_301)
);

INVx3_ASAP7_75t_L g302 ( 
.A(n_280),
.Y(n_302)
);

NAND2xp5_ASAP7_75t_L g303 ( 
.A(n_211),
.B(n_2),
.Y(n_303)
);

INVx2_ASAP7_75t_L g304 ( 
.A(n_218),
.Y(n_304)
);

BUFx3_ASAP7_75t_L g305 ( 
.A(n_220),
.Y(n_305)
);

BUFx6f_ASAP7_75t_L g306 ( 
.A(n_275),
.Y(n_306)
);

NOR2xp33_ASAP7_75t_L g307 ( 
.A(n_227),
.B(n_2),
.Y(n_307)
);

AND2x4_ASAP7_75t_L g308 ( 
.A(n_216),
.B(n_3),
.Y(n_308)
);

BUFx6f_ASAP7_75t_L g309 ( 
.A(n_231),
.Y(n_309)
);

XNOR2x2_ASAP7_75t_L g310 ( 
.A(n_207),
.B(n_3),
.Y(n_310)
);

BUFx6f_ASAP7_75t_L g311 ( 
.A(n_232),
.Y(n_311)
);

NOR2xp33_ASAP7_75t_L g312 ( 
.A(n_239),
.B(n_4),
.Y(n_312)
);

BUFx2_ASAP7_75t_L g313 ( 
.A(n_217),
.Y(n_313)
);

AND2x2_ASAP7_75t_L g314 ( 
.A(n_278),
.B(n_4),
.Y(n_314)
);

BUFx6f_ASAP7_75t_L g315 ( 
.A(n_243),
.Y(n_315)
);

NAND2xp5_ASAP7_75t_L g316 ( 
.A(n_247),
.B(n_5),
.Y(n_316)
);

INVx2_ASAP7_75t_L g317 ( 
.A(n_250),
.Y(n_317)
);

AND2x2_ASAP7_75t_L g318 ( 
.A(n_230),
.B(n_6),
.Y(n_318)
);

BUFx6f_ASAP7_75t_L g319 ( 
.A(n_253),
.Y(n_319)
);

NAND2xp5_ASAP7_75t_L g320 ( 
.A(n_255),
.B(n_6),
.Y(n_320)
);

INVx5_ASAP7_75t_L g321 ( 
.A(n_205),
.Y(n_321)
);

NOR2xp33_ASAP7_75t_L g322 ( 
.A(n_261),
.B(n_7),
.Y(n_322)
);

HB1xp67_ASAP7_75t_L g323 ( 
.A(n_234),
.Y(n_323)
);

INVx5_ASAP7_75t_L g324 ( 
.A(n_226),
.Y(n_324)
);

BUFx2_ASAP7_75t_L g325 ( 
.A(n_236),
.Y(n_325)
);

AND2x2_ASAP7_75t_L g326 ( 
.A(n_260),
.B(n_8),
.Y(n_326)
);

NAND2xp5_ASAP7_75t_L g327 ( 
.A(n_262),
.B(n_8),
.Y(n_327)
);

BUFx12f_ASAP7_75t_L g328 ( 
.A(n_228),
.Y(n_328)
);

AND2x2_ASAP7_75t_L g329 ( 
.A(n_272),
.B(n_9),
.Y(n_329)
);

INVx2_ASAP7_75t_L g330 ( 
.A(n_265),
.Y(n_330)
);

AND2x4_ASAP7_75t_L g331 ( 
.A(n_240),
.B(n_9),
.Y(n_331)
);

AND2x4_ASAP7_75t_L g332 ( 
.A(n_264),
.B(n_10),
.Y(n_332)
);

BUFx6f_ASAP7_75t_L g333 ( 
.A(n_277),
.Y(n_333)
);

BUFx6f_ASAP7_75t_L g334 ( 
.A(n_279),
.Y(n_334)
);

BUFx2_ASAP7_75t_L g335 ( 
.A(n_210),
.Y(n_335)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_201),
.Y(n_336)
);

AND2x4_ASAP7_75t_L g337 ( 
.A(n_210),
.B(n_11),
.Y(n_337)
);

AND2x2_ASAP7_75t_L g338 ( 
.A(n_313),
.B(n_259),
.Y(n_338)
);

OAI22xp33_ASAP7_75t_L g339 ( 
.A1(n_337),
.A2(n_276),
.B1(n_259),
.B2(n_271),
.Y(n_339)
);

NAND3x1_ASAP7_75t_L g340 ( 
.A(n_310),
.B(n_276),
.C(n_12),
.Y(n_340)
);

OAI22xp33_ASAP7_75t_SL g341 ( 
.A1(n_337),
.A2(n_273),
.B1(n_270),
.B2(n_269),
.Y(n_341)
);

AND2x2_ASAP7_75t_L g342 ( 
.A(n_325),
.B(n_202),
.Y(n_342)
);

AND2x2_ASAP7_75t_L g343 ( 
.A(n_300),
.B(n_208),
.Y(n_343)
);

OAI22xp5_ASAP7_75t_L g344 ( 
.A1(n_291),
.A2(n_268),
.B1(n_267),
.B2(n_266),
.Y(n_344)
);

AND2x4_ASAP7_75t_L g345 ( 
.A(n_295),
.B(n_209),
.Y(n_345)
);

OAI22xp33_ASAP7_75t_SL g346 ( 
.A1(n_337),
.A2(n_263),
.B1(n_258),
.B2(n_257),
.Y(n_346)
);

AND2x2_ASAP7_75t_L g347 ( 
.A(n_323),
.B(n_212),
.Y(n_347)
);

INVx2_ASAP7_75t_L g348 ( 
.A(n_292),
.Y(n_348)
);

INVx1_ASAP7_75t_L g349 ( 
.A(n_309),
.Y(n_349)
);

AO22x2_ASAP7_75t_L g350 ( 
.A1(n_298),
.A2(n_13),
.B1(n_14),
.B2(n_15),
.Y(n_350)
);

AO22x2_ASAP7_75t_L g351 ( 
.A1(n_314),
.A2(n_13),
.B1(n_14),
.B2(n_15),
.Y(n_351)
);

INVx2_ASAP7_75t_L g352 ( 
.A(n_292),
.Y(n_352)
);

INVx2_ASAP7_75t_L g353 ( 
.A(n_292),
.Y(n_353)
);

AOI22xp5_ASAP7_75t_L g354 ( 
.A1(n_291),
.A2(n_256),
.B1(n_252),
.B2(n_251),
.Y(n_354)
);

OAI22xp33_ASAP7_75t_L g355 ( 
.A1(n_282),
.A2(n_249),
.B1(n_248),
.B2(n_245),
.Y(n_355)
);

BUFx2_ASAP7_75t_L g356 ( 
.A(n_323),
.Y(n_356)
);

INVx1_ASAP7_75t_SL g357 ( 
.A(n_335),
.Y(n_357)
);

OAI22xp33_ASAP7_75t_L g358 ( 
.A1(n_288),
.A2(n_244),
.B1(n_242),
.B2(n_241),
.Y(n_358)
);

INVx1_ASAP7_75t_L g359 ( 
.A(n_306),
.Y(n_359)
);

CKINVDCx5p33_ASAP7_75t_R g360 ( 
.A(n_328),
.Y(n_360)
);

OAI22xp5_ASAP7_75t_SL g361 ( 
.A1(n_310),
.A2(n_237),
.B1(n_235),
.B2(n_233),
.Y(n_361)
);

INVx1_ASAP7_75t_L g362 ( 
.A(n_309),
.Y(n_362)
);

NAND2xp5_ASAP7_75t_L g363 ( 
.A(n_336),
.B(n_213),
.Y(n_363)
);

NAND2xp5_ASAP7_75t_L g364 ( 
.A(n_295),
.B(n_284),
.Y(n_364)
);

AOI22xp5_ASAP7_75t_L g365 ( 
.A1(n_288),
.A2(n_229),
.B1(n_224),
.B2(n_223),
.Y(n_365)
);

BUFx10_ASAP7_75t_L g366 ( 
.A(n_331),
.Y(n_366)
);

OR2x6_ASAP7_75t_L g367 ( 
.A(n_328),
.B(n_16),
.Y(n_367)
);

INVx1_ASAP7_75t_SL g368 ( 
.A(n_318),
.Y(n_368)
);

OAI22xp33_ASAP7_75t_SL g369 ( 
.A1(n_294),
.A2(n_222),
.B1(n_221),
.B2(n_219),
.Y(n_369)
);

AND2x2_ASAP7_75t_L g370 ( 
.A(n_281),
.B(n_215),
.Y(n_370)
);

OAI22xp33_ASAP7_75t_L g371 ( 
.A1(n_283),
.A2(n_16),
.B1(n_17),
.B2(n_18),
.Y(n_371)
);

OAI22xp33_ASAP7_75t_L g372 ( 
.A1(n_294),
.A2(n_17),
.B1(n_19),
.B2(n_20),
.Y(n_372)
);

INVx1_ASAP7_75t_L g373 ( 
.A(n_309),
.Y(n_373)
);

INVx1_ASAP7_75t_L g374 ( 
.A(n_306),
.Y(n_374)
);

INVx2_ASAP7_75t_L g375 ( 
.A(n_292),
.Y(n_375)
);

AND3x1_ASAP7_75t_L g376 ( 
.A(n_307),
.B(n_19),
.C(n_20),
.Y(n_376)
);

AND2x2_ASAP7_75t_L g377 ( 
.A(n_285),
.B(n_22),
.Y(n_377)
);

OR2x6_ASAP7_75t_L g378 ( 
.A(n_304),
.B(n_317),
.Y(n_378)
);

OAI22xp33_ASAP7_75t_SL g379 ( 
.A1(n_303),
.A2(n_22),
.B1(n_23),
.B2(n_24),
.Y(n_379)
);

AOI22xp5_ASAP7_75t_L g380 ( 
.A1(n_331),
.A2(n_24),
.B1(n_25),
.B2(n_28),
.Y(n_380)
);

AOI22xp5_ASAP7_75t_L g381 ( 
.A1(n_331),
.A2(n_30),
.B1(n_31),
.B2(n_34),
.Y(n_381)
);

AO22x2_ASAP7_75t_L g382 ( 
.A1(n_308),
.A2(n_35),
.B1(n_37),
.B2(n_44),
.Y(n_382)
);

INVx1_ASAP7_75t_L g383 ( 
.A(n_309),
.Y(n_383)
);

AOI22xp5_ASAP7_75t_L g384 ( 
.A1(n_332),
.A2(n_45),
.B1(n_46),
.B2(n_48),
.Y(n_384)
);

INVx2_ASAP7_75t_L g385 ( 
.A(n_297),
.Y(n_385)
);

OAI22xp33_ASAP7_75t_L g386 ( 
.A1(n_316),
.A2(n_49),
.B1(n_51),
.B2(n_52),
.Y(n_386)
);

AOI22xp5_ASAP7_75t_L g387 ( 
.A1(n_332),
.A2(n_55),
.B1(n_56),
.B2(n_58),
.Y(n_387)
);

AOI22xp5_ASAP7_75t_L g388 ( 
.A1(n_332),
.A2(n_61),
.B1(n_62),
.B2(n_64),
.Y(n_388)
);

INVx2_ASAP7_75t_L g389 ( 
.A(n_297),
.Y(n_389)
);

NOR2xp33_ASAP7_75t_L g390 ( 
.A(n_321),
.B(n_66),
.Y(n_390)
);

AOI22xp5_ASAP7_75t_L g391 ( 
.A1(n_326),
.A2(n_68),
.B1(n_69),
.B2(n_71),
.Y(n_391)
);

INVx8_ASAP7_75t_L g392 ( 
.A(n_321),
.Y(n_392)
);

INVx1_ASAP7_75t_L g393 ( 
.A(n_359),
.Y(n_393)
);

AND2x4_ASAP7_75t_L g394 ( 
.A(n_345),
.B(n_305),
.Y(n_394)
);

INVx2_ASAP7_75t_L g395 ( 
.A(n_359),
.Y(n_395)
);

NAND2x1p5_ASAP7_75t_L g396 ( 
.A(n_380),
.B(n_308),
.Y(n_396)
);

INVx3_ASAP7_75t_L g397 ( 
.A(n_378),
.Y(n_397)
);

CKINVDCx20_ASAP7_75t_R g398 ( 
.A(n_357),
.Y(n_398)
);

BUFx3_ASAP7_75t_L g399 ( 
.A(n_364),
.Y(n_399)
);

INVx2_ASAP7_75t_L g400 ( 
.A(n_374),
.Y(n_400)
);

OAI21xp5_ASAP7_75t_L g401 ( 
.A1(n_363),
.A2(n_320),
.B(n_327),
.Y(n_401)
);

INVx1_ASAP7_75t_L g402 ( 
.A(n_374),
.Y(n_402)
);

HB1xp67_ASAP7_75t_L g403 ( 
.A(n_356),
.Y(n_403)
);

OR2x2_ASAP7_75t_L g404 ( 
.A(n_338),
.B(n_305),
.Y(n_404)
);

NOR2xp33_ASAP7_75t_L g405 ( 
.A(n_366),
.B(n_321),
.Y(n_405)
);

OAI21xp5_ASAP7_75t_L g406 ( 
.A1(n_370),
.A2(n_308),
.B(n_289),
.Y(n_406)
);

INVx1_ASAP7_75t_L g407 ( 
.A(n_349),
.Y(n_407)
);

AND2x2_ASAP7_75t_L g408 ( 
.A(n_368),
.B(n_293),
.Y(n_408)
);

INVx1_ASAP7_75t_L g409 ( 
.A(n_362),
.Y(n_409)
);

BUFx3_ASAP7_75t_L g410 ( 
.A(n_378),
.Y(n_410)
);

INVxp33_ASAP7_75t_L g411 ( 
.A(n_347),
.Y(n_411)
);

OAI21xp5_ASAP7_75t_L g412 ( 
.A1(n_345),
.A2(n_307),
.B(n_312),
.Y(n_412)
);

CKINVDCx5p33_ASAP7_75t_R g413 ( 
.A(n_360),
.Y(n_413)
);

INVx1_ASAP7_75t_L g414 ( 
.A(n_373),
.Y(n_414)
);

INVx1_ASAP7_75t_L g415 ( 
.A(n_383),
.Y(n_415)
);

INVx1_ASAP7_75t_L g416 ( 
.A(n_377),
.Y(n_416)
);

CKINVDCx16_ASAP7_75t_R g417 ( 
.A(n_354),
.Y(n_417)
);

AND2x2_ASAP7_75t_L g418 ( 
.A(n_343),
.B(n_284),
.Y(n_418)
);

CKINVDCx20_ASAP7_75t_R g419 ( 
.A(n_361),
.Y(n_419)
);

OR2x2_ASAP7_75t_L g420 ( 
.A(n_339),
.B(n_304),
.Y(n_420)
);

XOR2xp5_ASAP7_75t_L g421 ( 
.A(n_382),
.B(n_329),
.Y(n_421)
);

INVx2_ASAP7_75t_SL g422 ( 
.A(n_342),
.Y(n_422)
);

AND2x2_ASAP7_75t_L g423 ( 
.A(n_366),
.B(n_286),
.Y(n_423)
);

INVx1_ASAP7_75t_L g424 ( 
.A(n_348),
.Y(n_424)
);

INVx1_ASAP7_75t_L g425 ( 
.A(n_352),
.Y(n_425)
);

XOR2xp5_ASAP7_75t_L g426 ( 
.A(n_382),
.B(n_311),
.Y(n_426)
);

INVx1_ASAP7_75t_L g427 ( 
.A(n_353),
.Y(n_427)
);

INVx1_ASAP7_75t_L g428 ( 
.A(n_375),
.Y(n_428)
);

CKINVDCx20_ASAP7_75t_R g429 ( 
.A(n_367),
.Y(n_429)
);

INVx1_ASAP7_75t_L g430 ( 
.A(n_385),
.Y(n_430)
);

INVx1_ASAP7_75t_L g431 ( 
.A(n_389),
.Y(n_431)
);

OAI21xp5_ASAP7_75t_L g432 ( 
.A1(n_381),
.A2(n_312),
.B(n_322),
.Y(n_432)
);

INVx1_ASAP7_75t_L g433 ( 
.A(n_384),
.Y(n_433)
);

INVx1_ASAP7_75t_L g434 ( 
.A(n_387),
.Y(n_434)
);

INVx1_ASAP7_75t_L g435 ( 
.A(n_388),
.Y(n_435)
);

XOR2xp5_ASAP7_75t_L g436 ( 
.A(n_344),
.B(n_311),
.Y(n_436)
);

CKINVDCx16_ASAP7_75t_R g437 ( 
.A(n_367),
.Y(n_437)
);

INVx1_ASAP7_75t_L g438 ( 
.A(n_372),
.Y(n_438)
);

INVx1_ASAP7_75t_L g439 ( 
.A(n_392),
.Y(n_439)
);

INVx1_ASAP7_75t_L g440 ( 
.A(n_392),
.Y(n_440)
);

XNOR2xp5_ASAP7_75t_L g441 ( 
.A(n_340),
.B(n_317),
.Y(n_441)
);

INVx1_ASAP7_75t_L g442 ( 
.A(n_365),
.Y(n_442)
);

NOR2xp33_ASAP7_75t_L g443 ( 
.A(n_358),
.B(n_355),
.Y(n_443)
);

INVx2_ASAP7_75t_L g444 ( 
.A(n_391),
.Y(n_444)
);

INVx2_ASAP7_75t_SL g445 ( 
.A(n_350),
.Y(n_445)
);

INVx1_ASAP7_75t_L g446 ( 
.A(n_379),
.Y(n_446)
);

INVx1_ASAP7_75t_L g447 ( 
.A(n_350),
.Y(n_447)
);

NOR2xp33_ASAP7_75t_L g448 ( 
.A(n_369),
.B(n_321),
.Y(n_448)
);

CKINVDCx5p33_ASAP7_75t_R g449 ( 
.A(n_341),
.Y(n_449)
);

INVx2_ASAP7_75t_L g450 ( 
.A(n_390),
.Y(n_450)
);

AND2x2_ASAP7_75t_L g451 ( 
.A(n_351),
.B(n_286),
.Y(n_451)
);

NOR2xp33_ASAP7_75t_L g452 ( 
.A(n_346),
.B(n_324),
.Y(n_452)
);

NOR2xp33_ASAP7_75t_L g453 ( 
.A(n_371),
.B(n_324),
.Y(n_453)
);

AND2x2_ASAP7_75t_L g454 ( 
.A(n_351),
.B(n_286),
.Y(n_454)
);

INVx4_ASAP7_75t_SL g455 ( 
.A(n_386),
.Y(n_455)
);

AND2x2_ASAP7_75t_L g456 ( 
.A(n_376),
.B(n_330),
.Y(n_456)
);

INVx1_ASAP7_75t_L g457 ( 
.A(n_359),
.Y(n_457)
);

INVx1_ASAP7_75t_L g458 ( 
.A(n_359),
.Y(n_458)
);

BUFx3_ASAP7_75t_L g459 ( 
.A(n_364),
.Y(n_459)
);

NAND2xp5_ASAP7_75t_SL g460 ( 
.A(n_369),
.B(n_306),
.Y(n_460)
);

INVxp33_ASAP7_75t_L g461 ( 
.A(n_338),
.Y(n_461)
);

CKINVDCx20_ASAP7_75t_R g462 ( 
.A(n_357),
.Y(n_462)
);

XNOR2x2_ASAP7_75t_L g463 ( 
.A(n_350),
.B(n_322),
.Y(n_463)
);

BUFx6f_ASAP7_75t_L g464 ( 
.A(n_349),
.Y(n_464)
);

INVx1_ASAP7_75t_L g465 ( 
.A(n_393),
.Y(n_465)
);

BUFx3_ASAP7_75t_L g466 ( 
.A(n_410),
.Y(n_466)
);

AND2x2_ASAP7_75t_L g467 ( 
.A(n_408),
.B(n_456),
.Y(n_467)
);

INVx1_ASAP7_75t_L g468 ( 
.A(n_402),
.Y(n_468)
);

AND2x2_ASAP7_75t_L g469 ( 
.A(n_406),
.B(n_330),
.Y(n_469)
);

AND2x2_ASAP7_75t_L g470 ( 
.A(n_418),
.B(n_296),
.Y(n_470)
);

AND2x2_ASAP7_75t_L g471 ( 
.A(n_394),
.B(n_296),
.Y(n_471)
);

INVx2_ASAP7_75t_L g472 ( 
.A(n_395),
.Y(n_472)
);

NAND2xp5_ASAP7_75t_L g473 ( 
.A(n_423),
.B(n_296),
.Y(n_473)
);

BUFx6f_ASAP7_75t_L g474 ( 
.A(n_464),
.Y(n_474)
);

INVx2_ASAP7_75t_L g475 ( 
.A(n_400),
.Y(n_475)
);

AND2x2_ASAP7_75t_L g476 ( 
.A(n_394),
.B(n_302),
.Y(n_476)
);

BUFx6f_ASAP7_75t_L g477 ( 
.A(n_464),
.Y(n_477)
);

INVx3_ASAP7_75t_L g478 ( 
.A(n_464),
.Y(n_478)
);

HB1xp67_ASAP7_75t_L g479 ( 
.A(n_403),
.Y(n_479)
);

NAND2xp5_ASAP7_75t_L g480 ( 
.A(n_399),
.B(n_302),
.Y(n_480)
);

AND2x2_ASAP7_75t_L g481 ( 
.A(n_451),
.B(n_302),
.Y(n_481)
);

BUFx6f_ASAP7_75t_L g482 ( 
.A(n_464),
.Y(n_482)
);

OAI21xp5_ASAP7_75t_L g483 ( 
.A1(n_401),
.A2(n_299),
.B(n_301),
.Y(n_483)
);

NAND2xp5_ASAP7_75t_SL g484 ( 
.A(n_422),
.B(n_324),
.Y(n_484)
);

BUFx6f_ASAP7_75t_L g485 ( 
.A(n_399),
.Y(n_485)
);

AND2x6_ASAP7_75t_L g486 ( 
.A(n_454),
.B(n_306),
.Y(n_486)
);

AND2x2_ASAP7_75t_L g487 ( 
.A(n_420),
.B(n_412),
.Y(n_487)
);

AND2x2_ASAP7_75t_L g488 ( 
.A(n_411),
.B(n_311),
.Y(n_488)
);

INVx1_ASAP7_75t_L g489 ( 
.A(n_457),
.Y(n_489)
);

BUFx6f_ASAP7_75t_L g490 ( 
.A(n_459),
.Y(n_490)
);

INVx3_ASAP7_75t_L g491 ( 
.A(n_459),
.Y(n_491)
);

INVxp33_ASAP7_75t_L g492 ( 
.A(n_403),
.Y(n_492)
);

INVxp67_ASAP7_75t_L g493 ( 
.A(n_404),
.Y(n_493)
);

INVx2_ASAP7_75t_L g494 ( 
.A(n_458),
.Y(n_494)
);

NAND2xp5_ASAP7_75t_L g495 ( 
.A(n_433),
.B(n_311),
.Y(n_495)
);

INVx3_ASAP7_75t_L g496 ( 
.A(n_407),
.Y(n_496)
);

INVx2_ASAP7_75t_L g497 ( 
.A(n_409),
.Y(n_497)
);

NAND2xp5_ASAP7_75t_L g498 ( 
.A(n_434),
.B(n_315),
.Y(n_498)
);

INVx1_ASAP7_75t_L g499 ( 
.A(n_414),
.Y(n_499)
);

AND2x2_ASAP7_75t_L g500 ( 
.A(n_411),
.B(n_315),
.Y(n_500)
);

AND2x4_ASAP7_75t_L g501 ( 
.A(n_445),
.B(n_315),
.Y(n_501)
);

NAND2xp5_ASAP7_75t_L g502 ( 
.A(n_435),
.B(n_315),
.Y(n_502)
);

OAI21xp5_ASAP7_75t_L g503 ( 
.A1(n_432),
.A2(n_301),
.B(n_299),
.Y(n_503)
);

AND2x2_ASAP7_75t_L g504 ( 
.A(n_397),
.B(n_319),
.Y(n_504)
);

INVx1_ASAP7_75t_L g505 ( 
.A(n_415),
.Y(n_505)
);

AND2x2_ASAP7_75t_L g506 ( 
.A(n_397),
.B(n_319),
.Y(n_506)
);

NAND2xp5_ASAP7_75t_L g507 ( 
.A(n_443),
.B(n_319),
.Y(n_507)
);

AND2x2_ASAP7_75t_L g508 ( 
.A(n_438),
.B(n_319),
.Y(n_508)
);

AND2x2_ASAP7_75t_L g509 ( 
.A(n_416),
.B(n_333),
.Y(n_509)
);

AND2x2_ASAP7_75t_L g510 ( 
.A(n_446),
.B(n_333),
.Y(n_510)
);

NAND2xp5_ASAP7_75t_L g511 ( 
.A(n_443),
.B(n_333),
.Y(n_511)
);

INVx1_ASAP7_75t_L g512 ( 
.A(n_424),
.Y(n_512)
);

NAND2xp5_ASAP7_75t_L g513 ( 
.A(n_444),
.B(n_333),
.Y(n_513)
);

NAND2xp5_ASAP7_75t_L g514 ( 
.A(n_442),
.B(n_334),
.Y(n_514)
);

INVx2_ASAP7_75t_L g515 ( 
.A(n_425),
.Y(n_515)
);

NAND2xp5_ASAP7_75t_L g516 ( 
.A(n_405),
.B(n_334),
.Y(n_516)
);

INVxp67_ASAP7_75t_L g517 ( 
.A(n_436),
.Y(n_517)
);

INVx2_ASAP7_75t_L g518 ( 
.A(n_427),
.Y(n_518)
);

NAND2xp5_ASAP7_75t_L g519 ( 
.A(n_405),
.B(n_334),
.Y(n_519)
);

AND2x6_ASAP7_75t_L g520 ( 
.A(n_447),
.B(n_334),
.Y(n_520)
);

INVx2_ASAP7_75t_L g521 ( 
.A(n_428),
.Y(n_521)
);

BUFx6f_ASAP7_75t_L g522 ( 
.A(n_430),
.Y(n_522)
);

INVx2_ASAP7_75t_L g523 ( 
.A(n_431),
.Y(n_523)
);

INVx2_ASAP7_75t_L g524 ( 
.A(n_450),
.Y(n_524)
);

HB1xp67_ASAP7_75t_L g525 ( 
.A(n_398),
.Y(n_525)
);

NAND2xp5_ASAP7_75t_L g526 ( 
.A(n_396),
.B(n_324),
.Y(n_526)
);

NOR2xp33_ASAP7_75t_R g527 ( 
.A(n_413),
.B(n_299),
.Y(n_527)
);

INVx2_ASAP7_75t_L g528 ( 
.A(n_460),
.Y(n_528)
);

BUFx3_ASAP7_75t_L g529 ( 
.A(n_398),
.Y(n_529)
);

AND2x2_ASAP7_75t_SL g530 ( 
.A(n_463),
.B(n_297),
.Y(n_530)
);

AND2x2_ASAP7_75t_L g531 ( 
.A(n_461),
.B(n_453),
.Y(n_531)
);

AND2x2_ASAP7_75t_L g532 ( 
.A(n_461),
.B(n_299),
.Y(n_532)
);

INVx4_ASAP7_75t_L g533 ( 
.A(n_455),
.Y(n_533)
);

INVx2_ASAP7_75t_L g534 ( 
.A(n_460),
.Y(n_534)
);

INVx1_ASAP7_75t_L g535 ( 
.A(n_396),
.Y(n_535)
);

INVx1_ASAP7_75t_L g536 ( 
.A(n_455),
.Y(n_536)
);

NAND2xp5_ASAP7_75t_L g537 ( 
.A(n_448),
.B(n_301),
.Y(n_537)
);

NAND2xp5_ASAP7_75t_L g538 ( 
.A(n_448),
.B(n_301),
.Y(n_538)
);

OR2x2_ASAP7_75t_L g539 ( 
.A(n_525),
.B(n_417),
.Y(n_539)
);

INVx2_ASAP7_75t_L g540 ( 
.A(n_494),
.Y(n_540)
);

NAND2xp5_ASAP7_75t_L g541 ( 
.A(n_487),
.B(n_453),
.Y(n_541)
);

BUFx12f_ASAP7_75t_L g542 ( 
.A(n_529),
.Y(n_542)
);

INVx1_ASAP7_75t_L g543 ( 
.A(n_465),
.Y(n_543)
);

INVx2_ASAP7_75t_SL g544 ( 
.A(n_529),
.Y(n_544)
);

NAND2xp5_ASAP7_75t_L g545 ( 
.A(n_487),
.B(n_426),
.Y(n_545)
);

NOR2xp33_ASAP7_75t_L g546 ( 
.A(n_492),
.B(n_421),
.Y(n_546)
);

INVx1_ASAP7_75t_L g547 ( 
.A(n_465),
.Y(n_547)
);

AND2x2_ASAP7_75t_L g548 ( 
.A(n_467),
.B(n_531),
.Y(n_548)
);

HB1xp67_ASAP7_75t_L g549 ( 
.A(n_479),
.Y(n_549)
);

OR2x6_ASAP7_75t_L g550 ( 
.A(n_533),
.B(n_462),
.Y(n_550)
);

BUFx2_ASAP7_75t_L g551 ( 
.A(n_466),
.Y(n_551)
);

AND2x4_ASAP7_75t_L g552 ( 
.A(n_533),
.B(n_439),
.Y(n_552)
);

INVx1_ASAP7_75t_L g553 ( 
.A(n_468),
.Y(n_553)
);

AND2x2_ASAP7_75t_SL g554 ( 
.A(n_530),
.B(n_437),
.Y(n_554)
);

OR2x2_ASAP7_75t_L g555 ( 
.A(n_493),
.B(n_441),
.Y(n_555)
);

OR2x6_ASAP7_75t_L g556 ( 
.A(n_533),
.B(n_466),
.Y(n_556)
);

AND2x2_ASAP7_75t_L g557 ( 
.A(n_467),
.B(n_462),
.Y(n_557)
);

NAND2xp5_ASAP7_75t_SL g558 ( 
.A(n_527),
.B(n_485),
.Y(n_558)
);

BUFx4f_ASAP7_75t_L g559 ( 
.A(n_536),
.Y(n_559)
);

INVx5_ASAP7_75t_L g560 ( 
.A(n_520),
.Y(n_560)
);

NAND2xp5_ASAP7_75t_L g561 ( 
.A(n_469),
.B(n_455),
.Y(n_561)
);

INVx4_ASAP7_75t_L g562 ( 
.A(n_485),
.Y(n_562)
);

INVx2_ASAP7_75t_L g563 ( 
.A(n_494),
.Y(n_563)
);

NAND2x1p5_ASAP7_75t_L g564 ( 
.A(n_535),
.B(n_440),
.Y(n_564)
);

BUFx6f_ASAP7_75t_L g565 ( 
.A(n_474),
.Y(n_565)
);

NAND2xp5_ASAP7_75t_L g566 ( 
.A(n_469),
.B(n_507),
.Y(n_566)
);

AND2x4_ASAP7_75t_L g567 ( 
.A(n_535),
.B(n_449),
.Y(n_567)
);

INVx4_ASAP7_75t_L g568 ( 
.A(n_485),
.Y(n_568)
);

NAND2x1p5_ASAP7_75t_L g569 ( 
.A(n_536),
.B(n_452),
.Y(n_569)
);

NOR2xp33_ASAP7_75t_L g570 ( 
.A(n_531),
.B(n_419),
.Y(n_570)
);

AND2x6_ASAP7_75t_L g571 ( 
.A(n_501),
.B(n_452),
.Y(n_571)
);

NAND2xp5_ASAP7_75t_L g572 ( 
.A(n_511),
.B(n_419),
.Y(n_572)
);

NAND2xp5_ASAP7_75t_L g573 ( 
.A(n_481),
.B(n_524),
.Y(n_573)
);

NAND2xp5_ASAP7_75t_L g574 ( 
.A(n_481),
.B(n_429),
.Y(n_574)
);

AND2x4_ASAP7_75t_L g575 ( 
.A(n_471),
.B(n_429),
.Y(n_575)
);

NAND2xp5_ASAP7_75t_L g576 ( 
.A(n_524),
.B(n_297),
.Y(n_576)
);

OR2x6_ASAP7_75t_L g577 ( 
.A(n_517),
.B(n_74),
.Y(n_577)
);

INVx5_ASAP7_75t_L g578 ( 
.A(n_520),
.Y(n_578)
);

INVx1_ASAP7_75t_L g579 ( 
.A(n_468),
.Y(n_579)
);

BUFx3_ASAP7_75t_L g580 ( 
.A(n_471),
.Y(n_580)
);

INVxp67_ASAP7_75t_SL g581 ( 
.A(n_474),
.Y(n_581)
);

INVx1_ASAP7_75t_SL g582 ( 
.A(n_476),
.Y(n_582)
);

NAND2x1p5_ASAP7_75t_L g583 ( 
.A(n_476),
.B(n_287),
.Y(n_583)
);

BUFx4f_ASAP7_75t_L g584 ( 
.A(n_520),
.Y(n_584)
);

OR2x6_ASAP7_75t_L g585 ( 
.A(n_501),
.B(n_77),
.Y(n_585)
);

NAND2x1p5_ASAP7_75t_L g586 ( 
.A(n_485),
.B(n_287),
.Y(n_586)
);

NAND2xp5_ASAP7_75t_L g587 ( 
.A(n_528),
.B(n_287),
.Y(n_587)
);

INVx2_ASAP7_75t_L g588 ( 
.A(n_472),
.Y(n_588)
);

INVx2_ASAP7_75t_L g589 ( 
.A(n_472),
.Y(n_589)
);

AND2x2_ASAP7_75t_L g590 ( 
.A(n_470),
.B(n_287),
.Y(n_590)
);

AND2x4_ASAP7_75t_L g591 ( 
.A(n_470),
.B(n_79),
.Y(n_591)
);

BUFx3_ASAP7_75t_L g592 ( 
.A(n_488),
.Y(n_592)
);

BUFx2_ASAP7_75t_L g593 ( 
.A(n_486),
.Y(n_593)
);

NAND2xp5_ASAP7_75t_L g594 ( 
.A(n_508),
.B(n_290),
.Y(n_594)
);

INVx1_ASAP7_75t_L g595 ( 
.A(n_489),
.Y(n_595)
);

INVx2_ASAP7_75t_L g596 ( 
.A(n_475),
.Y(n_596)
);

BUFx3_ASAP7_75t_L g597 ( 
.A(n_488),
.Y(n_597)
);

BUFx8_ASAP7_75t_SL g598 ( 
.A(n_485),
.Y(n_598)
);

OR2x2_ASAP7_75t_L g599 ( 
.A(n_500),
.B(n_80),
.Y(n_599)
);

BUFx2_ASAP7_75t_L g600 ( 
.A(n_549),
.Y(n_600)
);

AND2x2_ASAP7_75t_L g601 ( 
.A(n_541),
.B(n_530),
.Y(n_601)
);

BUFx12f_ASAP7_75t_L g602 ( 
.A(n_542),
.Y(n_602)
);

BUFx2_ASAP7_75t_L g603 ( 
.A(n_580),
.Y(n_603)
);

AND2x2_ASAP7_75t_L g604 ( 
.A(n_548),
.B(n_530),
.Y(n_604)
);

INVx6_ASAP7_75t_SL g605 ( 
.A(n_550),
.Y(n_605)
);

INVx3_ASAP7_75t_L g606 ( 
.A(n_565),
.Y(n_606)
);

BUFx3_ASAP7_75t_L g607 ( 
.A(n_598),
.Y(n_607)
);

BUFx4_ASAP7_75t_SL g608 ( 
.A(n_550),
.Y(n_608)
);

INVx1_ASAP7_75t_L g609 ( 
.A(n_543),
.Y(n_609)
);

BUFx2_ASAP7_75t_L g610 ( 
.A(n_557),
.Y(n_610)
);

INVx3_ASAP7_75t_L g611 ( 
.A(n_565),
.Y(n_611)
);

BUFx12f_ASAP7_75t_L g612 ( 
.A(n_551),
.Y(n_612)
);

BUFx2_ASAP7_75t_L g613 ( 
.A(n_592),
.Y(n_613)
);

BUFx2_ASAP7_75t_SL g614 ( 
.A(n_560),
.Y(n_614)
);

INVx2_ASAP7_75t_L g615 ( 
.A(n_588),
.Y(n_615)
);

BUFx3_ASAP7_75t_L g616 ( 
.A(n_556),
.Y(n_616)
);

OR2x6_ASAP7_75t_L g617 ( 
.A(n_585),
.B(n_490),
.Y(n_617)
);

BUFx2_ASAP7_75t_L g618 ( 
.A(n_597),
.Y(n_618)
);

BUFx2_ASAP7_75t_SL g619 ( 
.A(n_560),
.Y(n_619)
);

INVx1_ASAP7_75t_L g620 ( 
.A(n_543),
.Y(n_620)
);

BUFx12f_ASAP7_75t_L g621 ( 
.A(n_544),
.Y(n_621)
);

INVx1_ASAP7_75t_L g622 ( 
.A(n_547),
.Y(n_622)
);

OR2x2_ASAP7_75t_L g623 ( 
.A(n_545),
.B(n_473),
.Y(n_623)
);

INVx3_ASAP7_75t_L g624 ( 
.A(n_565),
.Y(n_624)
);

BUFx6f_ASAP7_75t_L g625 ( 
.A(n_584),
.Y(n_625)
);

INVx4_ASAP7_75t_L g626 ( 
.A(n_584),
.Y(n_626)
);

BUFx4f_ASAP7_75t_SL g627 ( 
.A(n_575),
.Y(n_627)
);

INVx8_ASAP7_75t_L g628 ( 
.A(n_585),
.Y(n_628)
);

INVx6_ASAP7_75t_L g629 ( 
.A(n_556),
.Y(n_629)
);

INVx2_ASAP7_75t_L g630 ( 
.A(n_589),
.Y(n_630)
);

BUFx3_ASAP7_75t_L g631 ( 
.A(n_552),
.Y(n_631)
);

INVx5_ASAP7_75t_L g632 ( 
.A(n_560),
.Y(n_632)
);

BUFx2_ASAP7_75t_SL g633 ( 
.A(n_578),
.Y(n_633)
);

BUFx2_ASAP7_75t_L g634 ( 
.A(n_575),
.Y(n_634)
);

INVx3_ASAP7_75t_L g635 ( 
.A(n_578),
.Y(n_635)
);

BUFx3_ASAP7_75t_L g636 ( 
.A(n_552),
.Y(n_636)
);

INVx1_ASAP7_75t_SL g637 ( 
.A(n_539),
.Y(n_637)
);

AOI22xp33_ASAP7_75t_L g638 ( 
.A1(n_570),
.A2(n_528),
.B1(n_534),
.B2(n_532),
.Y(n_638)
);

BUFx12f_ASAP7_75t_L g639 ( 
.A(n_577),
.Y(n_639)
);

BUFx3_ASAP7_75t_L g640 ( 
.A(n_559),
.Y(n_640)
);

INVx4_ASAP7_75t_L g641 ( 
.A(n_578),
.Y(n_641)
);

INVx5_ASAP7_75t_SL g642 ( 
.A(n_577),
.Y(n_642)
);

INVx1_ASAP7_75t_L g643 ( 
.A(n_547),
.Y(n_643)
);

BUFx12f_ASAP7_75t_L g644 ( 
.A(n_567),
.Y(n_644)
);

NAND2x1p5_ASAP7_75t_L g645 ( 
.A(n_559),
.B(n_474),
.Y(n_645)
);

BUFx3_ASAP7_75t_L g646 ( 
.A(n_571),
.Y(n_646)
);

INVx6_ASAP7_75t_L g647 ( 
.A(n_612),
.Y(n_647)
);

AOI22xp33_ASAP7_75t_L g648 ( 
.A1(n_601),
.A2(n_572),
.B1(n_554),
.B2(n_546),
.Y(n_648)
);

AOI22xp5_ASAP7_75t_L g649 ( 
.A1(n_604),
.A2(n_582),
.B1(n_571),
.B2(n_561),
.Y(n_649)
);

OAI22xp5_ASAP7_75t_SL g650 ( 
.A1(n_639),
.A2(n_555),
.B1(n_574),
.B2(n_582),
.Y(n_650)
);

INVx1_ASAP7_75t_L g651 ( 
.A(n_609),
.Y(n_651)
);

HB1xp67_ASAP7_75t_SL g652 ( 
.A(n_607),
.Y(n_652)
);

NAND2xp5_ASAP7_75t_L g653 ( 
.A(n_600),
.B(n_553),
.Y(n_653)
);

NAND2xp5_ASAP7_75t_L g654 ( 
.A(n_600),
.B(n_553),
.Y(n_654)
);

CKINVDCx5p33_ASAP7_75t_R g655 ( 
.A(n_602),
.Y(n_655)
);

BUFx2_ASAP7_75t_R g656 ( 
.A(n_607),
.Y(n_656)
);

INVx3_ASAP7_75t_L g657 ( 
.A(n_625),
.Y(n_657)
);

INVx1_ASAP7_75t_L g658 ( 
.A(n_622),
.Y(n_658)
);

INVx2_ASAP7_75t_SL g659 ( 
.A(n_612),
.Y(n_659)
);

OR2x2_ASAP7_75t_L g660 ( 
.A(n_610),
.B(n_567),
.Y(n_660)
);

OAI22xp5_ASAP7_75t_L g661 ( 
.A1(n_620),
.A2(n_595),
.B1(n_579),
.B2(n_643),
.Y(n_661)
);

INVx1_ASAP7_75t_L g662 ( 
.A(n_620),
.Y(n_662)
);

INVx1_ASAP7_75t_L g663 ( 
.A(n_615),
.Y(n_663)
);

BUFx6f_ASAP7_75t_SL g664 ( 
.A(n_616),
.Y(n_664)
);

BUFx12f_ASAP7_75t_L g665 ( 
.A(n_602),
.Y(n_665)
);

BUFx3_ASAP7_75t_L g666 ( 
.A(n_621),
.Y(n_666)
);

AOI22xp33_ASAP7_75t_L g667 ( 
.A1(n_601),
.A2(n_571),
.B1(n_540),
.B2(n_563),
.Y(n_667)
);

OAI22xp33_ASAP7_75t_L g668 ( 
.A1(n_610),
.A2(n_595),
.B1(n_579),
.B2(n_491),
.Y(n_668)
);

BUFx2_ASAP7_75t_L g669 ( 
.A(n_605),
.Y(n_669)
);

CKINVDCx5p33_ASAP7_75t_R g670 ( 
.A(n_608),
.Y(n_670)
);

CKINVDCx20_ASAP7_75t_R g671 ( 
.A(n_627),
.Y(n_671)
);

INVx6_ASAP7_75t_L g672 ( 
.A(n_621),
.Y(n_672)
);

AOI22xp33_ASAP7_75t_L g673 ( 
.A1(n_623),
.A2(n_571),
.B1(n_534),
.B2(n_532),
.Y(n_673)
);

BUFx3_ASAP7_75t_L g674 ( 
.A(n_644),
.Y(n_674)
);

CKINVDCx6p67_ASAP7_75t_R g675 ( 
.A(n_639),
.Y(n_675)
);

INVx6_ASAP7_75t_L g676 ( 
.A(n_644),
.Y(n_676)
);

OAI22xp33_ASAP7_75t_L g677 ( 
.A1(n_628),
.A2(n_491),
.B1(n_573),
.B2(n_599),
.Y(n_677)
);

INVx1_ASAP7_75t_L g678 ( 
.A(n_615),
.Y(n_678)
);

CKINVDCx20_ASAP7_75t_R g679 ( 
.A(n_642),
.Y(n_679)
);

BUFx12f_ASAP7_75t_L g680 ( 
.A(n_634),
.Y(n_680)
);

CKINVDCx11_ASAP7_75t_R g681 ( 
.A(n_637),
.Y(n_681)
);

INVx1_ASAP7_75t_L g682 ( 
.A(n_630),
.Y(n_682)
);

BUFx6f_ASAP7_75t_L g683 ( 
.A(n_631),
.Y(n_683)
);

BUFx8_ASAP7_75t_L g684 ( 
.A(n_634),
.Y(n_684)
);

INVxp67_ASAP7_75t_SL g685 ( 
.A(n_631),
.Y(n_685)
);

BUFx2_ASAP7_75t_SL g686 ( 
.A(n_640),
.Y(n_686)
);

INVx2_ASAP7_75t_L g687 ( 
.A(n_630),
.Y(n_687)
);

AOI22xp33_ASAP7_75t_L g688 ( 
.A1(n_623),
.A2(n_500),
.B1(n_566),
.B2(n_596),
.Y(n_688)
);

AND2x2_ASAP7_75t_L g689 ( 
.A(n_660),
.B(n_604),
.Y(n_689)
);

OR2x2_ASAP7_75t_L g690 ( 
.A(n_653),
.B(n_642),
.Y(n_690)
);

INVx2_ASAP7_75t_SL g691 ( 
.A(n_676),
.Y(n_691)
);

OAI22xp5_ASAP7_75t_L g692 ( 
.A1(n_668),
.A2(n_617),
.B1(n_642),
.B2(n_638),
.Y(n_692)
);

AOI22xp33_ASAP7_75t_SL g693 ( 
.A1(n_650),
.A2(n_628),
.B1(n_642),
.B2(n_617),
.Y(n_693)
);

NOR2x1_ASAP7_75t_L g694 ( 
.A(n_666),
.B(n_613),
.Y(n_694)
);

AOI22xp33_ASAP7_75t_L g695 ( 
.A1(n_648),
.A2(n_628),
.B1(n_605),
.B2(n_508),
.Y(n_695)
);

NOR2xp33_ASAP7_75t_L g696 ( 
.A(n_681),
.B(n_603),
.Y(n_696)
);

INVx2_ASAP7_75t_L g697 ( 
.A(n_687),
.Y(n_697)
);

INVx1_ASAP7_75t_L g698 ( 
.A(n_651),
.Y(n_698)
);

INVx1_ASAP7_75t_L g699 ( 
.A(n_658),
.Y(n_699)
);

OAI22xp5_ASAP7_75t_L g700 ( 
.A1(n_654),
.A2(n_617),
.B1(n_628),
.B2(n_591),
.Y(n_700)
);

AOI22xp33_ASAP7_75t_L g701 ( 
.A1(n_650),
.A2(n_605),
.B1(n_617),
.B2(n_497),
.Y(n_701)
);

AOI22xp33_ASAP7_75t_L g702 ( 
.A1(n_688),
.A2(n_673),
.B1(n_649),
.B2(n_497),
.Y(n_702)
);

INVx5_ASAP7_75t_SL g703 ( 
.A(n_675),
.Y(n_703)
);

BUFx6f_ASAP7_75t_L g704 ( 
.A(n_683),
.Y(n_704)
);

CKINVDCx5p33_ASAP7_75t_R g705 ( 
.A(n_670),
.Y(n_705)
);

BUFx2_ASAP7_75t_L g706 ( 
.A(n_684),
.Y(n_706)
);

CKINVDCx5p33_ASAP7_75t_R g707 ( 
.A(n_665),
.Y(n_707)
);

BUFx2_ASAP7_75t_L g708 ( 
.A(n_684),
.Y(n_708)
);

BUFx2_ASAP7_75t_L g709 ( 
.A(n_680),
.Y(n_709)
);

OAI21xp5_ASAP7_75t_SL g710 ( 
.A1(n_677),
.A2(n_503),
.B(n_591),
.Y(n_710)
);

CKINVDCx20_ASAP7_75t_R g711 ( 
.A(n_671),
.Y(n_711)
);

INVx2_ASAP7_75t_L g712 ( 
.A(n_663),
.Y(n_712)
);

OAI22xp5_ASAP7_75t_L g713 ( 
.A1(n_661),
.A2(n_636),
.B1(n_603),
.B2(n_618),
.Y(n_713)
);

INVx1_ASAP7_75t_L g714 ( 
.A(n_662),
.Y(n_714)
);

OAI22xp5_ASAP7_75t_L g715 ( 
.A1(n_661),
.A2(n_636),
.B1(n_618),
.B2(n_613),
.Y(n_715)
);

OAI21xp5_ASAP7_75t_SL g716 ( 
.A1(n_669),
.A2(n_483),
.B(n_509),
.Y(n_716)
);

AND2x4_ASAP7_75t_L g717 ( 
.A(n_683),
.B(n_646),
.Y(n_717)
);

AOI22xp33_ASAP7_75t_L g718 ( 
.A1(n_649),
.A2(n_646),
.B1(n_515),
.B2(n_523),
.Y(n_718)
);

INVx1_ASAP7_75t_L g719 ( 
.A(n_678),
.Y(n_719)
);

NOR2xp33_ASAP7_75t_L g720 ( 
.A(n_652),
.B(n_640),
.Y(n_720)
);

HB1xp67_ASAP7_75t_L g721 ( 
.A(n_682),
.Y(n_721)
);

CKINVDCx5p33_ASAP7_75t_R g722 ( 
.A(n_655),
.Y(n_722)
);

AOI22xp33_ASAP7_75t_SL g723 ( 
.A1(n_679),
.A2(n_629),
.B1(n_616),
.B2(n_520),
.Y(n_723)
);

OAI21xp5_ASAP7_75t_SL g724 ( 
.A1(n_659),
.A2(n_509),
.B(n_558),
.Y(n_724)
);

AOI22xp33_ASAP7_75t_L g725 ( 
.A1(n_667),
.A2(n_521),
.B1(n_515),
.B2(n_518),
.Y(n_725)
);

CKINVDCx5p33_ASAP7_75t_R g726 ( 
.A(n_656),
.Y(n_726)
);

OAI21xp5_ASAP7_75t_SL g727 ( 
.A1(n_657),
.A2(n_645),
.B(n_564),
.Y(n_727)
);

INVx2_ASAP7_75t_L g728 ( 
.A(n_683),
.Y(n_728)
);

AND2x2_ASAP7_75t_L g729 ( 
.A(n_674),
.B(n_504),
.Y(n_729)
);

NAND2xp5_ASAP7_75t_L g730 ( 
.A(n_685),
.B(n_510),
.Y(n_730)
);

INVx1_ASAP7_75t_L g731 ( 
.A(n_664),
.Y(n_731)
);

NAND2xp5_ASAP7_75t_L g732 ( 
.A(n_686),
.B(n_510),
.Y(n_732)
);

OAI222xp33_ASAP7_75t_L g733 ( 
.A1(n_657),
.A2(n_569),
.B1(n_502),
.B2(n_495),
.C1(n_498),
.C2(n_514),
.Y(n_733)
);

INVx2_ASAP7_75t_L g734 ( 
.A(n_664),
.Y(n_734)
);

OAI22xp5_ASAP7_75t_L g735 ( 
.A1(n_676),
.A2(n_489),
.B1(n_499),
.B2(n_505),
.Y(n_735)
);

INVx1_ASAP7_75t_L g736 ( 
.A(n_647),
.Y(n_736)
);

AOI22xp33_ASAP7_75t_L g737 ( 
.A1(n_647),
.A2(n_523),
.B1(n_518),
.B2(n_521),
.Y(n_737)
);

AOI22xp33_ASAP7_75t_L g738 ( 
.A1(n_695),
.A2(n_490),
.B1(n_475),
.B2(n_537),
.Y(n_738)
);

AOI22xp33_ASAP7_75t_L g739 ( 
.A1(n_695),
.A2(n_702),
.B1(n_701),
.B2(n_693),
.Y(n_739)
);

OAI21xp5_ASAP7_75t_L g740 ( 
.A1(n_710),
.A2(n_519),
.B(n_516),
.Y(n_740)
);

AOI22xp33_ASAP7_75t_L g741 ( 
.A1(n_702),
.A2(n_490),
.B1(n_538),
.B2(n_512),
.Y(n_741)
);

AOI22xp33_ASAP7_75t_SL g742 ( 
.A1(n_692),
.A2(n_629),
.B1(n_672),
.B2(n_520),
.Y(n_742)
);

HB1xp67_ASAP7_75t_L g743 ( 
.A(n_721),
.Y(n_743)
);

OAI22xp5_ASAP7_75t_L g744 ( 
.A1(n_735),
.A2(n_672),
.B1(n_629),
.B2(n_505),
.Y(n_744)
);

NAND3xp33_ASAP7_75t_L g745 ( 
.A(n_716),
.B(n_506),
.C(n_504),
.Y(n_745)
);

NAND2xp5_ASAP7_75t_L g746 ( 
.A(n_689),
.B(n_606),
.Y(n_746)
);

NAND2xp5_ASAP7_75t_L g747 ( 
.A(n_698),
.B(n_606),
.Y(n_747)
);

AOI22xp33_ASAP7_75t_L g748 ( 
.A1(n_701),
.A2(n_490),
.B1(n_512),
.B2(n_499),
.Y(n_748)
);

AOI22xp33_ASAP7_75t_L g749 ( 
.A1(n_718),
.A2(n_490),
.B1(n_522),
.B2(n_513),
.Y(n_749)
);

OAI22xp5_ASAP7_75t_L g750 ( 
.A1(n_713),
.A2(n_629),
.B1(n_496),
.B2(n_645),
.Y(n_750)
);

AOI22xp5_ASAP7_75t_L g751 ( 
.A1(n_700),
.A2(n_520),
.B1(n_486),
.B2(n_593),
.Y(n_751)
);

AOI22xp33_ASAP7_75t_L g752 ( 
.A1(n_693),
.A2(n_522),
.B1(n_491),
.B2(n_526),
.Y(n_752)
);

AOI22xp33_ASAP7_75t_SL g753 ( 
.A1(n_715),
.A2(n_520),
.B1(n_614),
.B2(n_619),
.Y(n_753)
);

AOI22xp33_ASAP7_75t_L g754 ( 
.A1(n_725),
.A2(n_522),
.B1(n_496),
.B2(n_506),
.Y(n_754)
);

OAI22xp5_ASAP7_75t_L g755 ( 
.A1(n_690),
.A2(n_496),
.B1(n_645),
.B2(n_606),
.Y(n_755)
);

AOI22xp33_ASAP7_75t_SL g756 ( 
.A1(n_732),
.A2(n_614),
.B1(n_633),
.B2(n_619),
.Y(n_756)
);

AND2x2_ASAP7_75t_L g757 ( 
.A(n_699),
.B(n_611),
.Y(n_757)
);

AOI22xp5_ASAP7_75t_L g758 ( 
.A1(n_724),
.A2(n_486),
.B1(n_501),
.B2(n_626),
.Y(n_758)
);

OAI22xp5_ASAP7_75t_L g759 ( 
.A1(n_696),
.A2(n_624),
.B1(n_611),
.B2(n_626),
.Y(n_759)
);

NOR3xp33_ASAP7_75t_L g760 ( 
.A(n_694),
.B(n_484),
.C(n_611),
.Y(n_760)
);

NAND2xp5_ASAP7_75t_L g761 ( 
.A(n_714),
.B(n_624),
.Y(n_761)
);

AOI22xp33_ASAP7_75t_L g762 ( 
.A1(n_712),
.A2(n_522),
.B1(n_590),
.B2(n_480),
.Y(n_762)
);

NAND2xp5_ASAP7_75t_L g763 ( 
.A(n_721),
.B(n_624),
.Y(n_763)
);

AOI22xp33_ASAP7_75t_L g764 ( 
.A1(n_730),
.A2(n_522),
.B1(n_594),
.B2(n_478),
.Y(n_764)
);

AOI221xp5_ASAP7_75t_L g765 ( 
.A1(n_729),
.A2(n_733),
.B1(n_736),
.B2(n_731),
.C(n_737),
.Y(n_765)
);

AOI22xp33_ASAP7_75t_L g766 ( 
.A1(n_723),
.A2(n_478),
.B1(n_562),
.B2(n_568),
.Y(n_766)
);

AOI22xp5_ASAP7_75t_L g767 ( 
.A1(n_723),
.A2(n_486),
.B1(n_626),
.B2(n_625),
.Y(n_767)
);

AOI22xp33_ASAP7_75t_L g768 ( 
.A1(n_697),
.A2(n_478),
.B1(n_562),
.B2(n_568),
.Y(n_768)
);

NAND2xp5_ASAP7_75t_L g769 ( 
.A(n_728),
.B(n_581),
.Y(n_769)
);

AND2x2_ASAP7_75t_L g770 ( 
.A(n_704),
.B(n_583),
.Y(n_770)
);

AOI22xp33_ASAP7_75t_SL g771 ( 
.A1(n_734),
.A2(n_633),
.B1(n_632),
.B2(n_625),
.Y(n_771)
);

OAI221xp5_ASAP7_75t_SL g772 ( 
.A1(n_727),
.A2(n_576),
.B1(n_635),
.B2(n_587),
.C(n_486),
.Y(n_772)
);

AOI22xp33_ASAP7_75t_SL g773 ( 
.A1(n_717),
.A2(n_632),
.B1(n_625),
.B2(n_641),
.Y(n_773)
);

AOI22xp33_ASAP7_75t_L g774 ( 
.A1(n_726),
.A2(n_706),
.B1(n_708),
.B2(n_719),
.Y(n_774)
);

AOI221xp5_ASAP7_75t_L g775 ( 
.A1(n_733),
.A2(n_587),
.B1(n_474),
.B2(n_477),
.C(n_482),
.Y(n_775)
);

AOI22xp33_ASAP7_75t_SL g776 ( 
.A1(n_717),
.A2(n_632),
.B1(n_625),
.B2(n_641),
.Y(n_776)
);

NAND2xp5_ASAP7_75t_L g777 ( 
.A(n_704),
.B(n_486),
.Y(n_777)
);

NAND2xp5_ASAP7_75t_L g778 ( 
.A(n_743),
.B(n_704),
.Y(n_778)
);

AOI211xp5_ASAP7_75t_L g779 ( 
.A1(n_745),
.A2(n_720),
.B(n_691),
.C(n_709),
.Y(n_779)
);

NAND2xp5_ASAP7_75t_L g780 ( 
.A(n_743),
.B(n_703),
.Y(n_780)
);

NAND3xp33_ASAP7_75t_L g781 ( 
.A(n_765),
.B(n_722),
.C(n_707),
.Y(n_781)
);

NAND2xp5_ASAP7_75t_L g782 ( 
.A(n_757),
.B(n_703),
.Y(n_782)
);

OAI21xp5_ASAP7_75t_SL g783 ( 
.A1(n_739),
.A2(n_703),
.B(n_635),
.Y(n_783)
);

OA21x2_ASAP7_75t_L g784 ( 
.A1(n_775),
.A2(n_705),
.B(n_586),
.Y(n_784)
);

NOR2xp33_ASAP7_75t_L g785 ( 
.A(n_759),
.B(n_711),
.Y(n_785)
);

NAND2xp5_ASAP7_75t_SL g786 ( 
.A(n_756),
.B(n_632),
.Y(n_786)
);

AND2x2_ASAP7_75t_SL g787 ( 
.A(n_739),
.B(n_763),
.Y(n_787)
);

INVx2_ASAP7_75t_L g788 ( 
.A(n_747),
.Y(n_788)
);

INVx1_ASAP7_75t_L g789 ( 
.A(n_761),
.Y(n_789)
);

NAND3xp33_ASAP7_75t_L g790 ( 
.A(n_760),
.B(n_482),
.C(n_477),
.Y(n_790)
);

NAND2xp5_ASAP7_75t_L g791 ( 
.A(n_746),
.B(n_635),
.Y(n_791)
);

NAND2xp5_ASAP7_75t_L g792 ( 
.A(n_774),
.B(n_474),
.Y(n_792)
);

OAI22xp5_ASAP7_75t_L g793 ( 
.A1(n_758),
.A2(n_632),
.B1(n_641),
.B2(n_482),
.Y(n_793)
);

NAND2xp5_ASAP7_75t_SL g794 ( 
.A(n_753),
.B(n_477),
.Y(n_794)
);

AND2x2_ASAP7_75t_L g795 ( 
.A(n_774),
.B(n_477),
.Y(n_795)
);

AND2x2_ASAP7_75t_SL g796 ( 
.A(n_767),
.B(n_477),
.Y(n_796)
);

AND2x2_ASAP7_75t_L g797 ( 
.A(n_770),
.B(n_482),
.Y(n_797)
);

OAI21xp5_ASAP7_75t_SL g798 ( 
.A1(n_744),
.A2(n_482),
.B(n_83),
.Y(n_798)
);

OAI21xp5_ASAP7_75t_SL g799 ( 
.A1(n_742),
.A2(n_81),
.B(n_85),
.Y(n_799)
);

NAND3xp33_ASAP7_75t_L g800 ( 
.A(n_764),
.B(n_290),
.C(n_88),
.Y(n_800)
);

NAND2xp5_ASAP7_75t_L g801 ( 
.A(n_750),
.B(n_87),
.Y(n_801)
);

NAND2xp5_ASAP7_75t_L g802 ( 
.A(n_755),
.B(n_89),
.Y(n_802)
);

NAND2xp5_ASAP7_75t_L g803 ( 
.A(n_769),
.B(n_90),
.Y(n_803)
);

AND2x2_ASAP7_75t_L g804 ( 
.A(n_777),
.B(n_91),
.Y(n_804)
);

NAND3xp33_ASAP7_75t_L g805 ( 
.A(n_740),
.B(n_290),
.C(n_94),
.Y(n_805)
);

OAI221xp5_ASAP7_75t_L g806 ( 
.A1(n_748),
.A2(n_290),
.B1(n_95),
.B2(n_97),
.C(n_98),
.Y(n_806)
);

AND2x2_ASAP7_75t_L g807 ( 
.A(n_780),
.B(n_752),
.Y(n_807)
);

HB1xp67_ASAP7_75t_L g808 ( 
.A(n_789),
.Y(n_808)
);

AND2x2_ASAP7_75t_L g809 ( 
.A(n_778),
.B(n_773),
.Y(n_809)
);

AOI22xp33_ASAP7_75t_L g810 ( 
.A1(n_787),
.A2(n_741),
.B1(n_738),
.B2(n_762),
.Y(n_810)
);

NAND3xp33_ASAP7_75t_L g811 ( 
.A(n_779),
.B(n_772),
.C(n_768),
.Y(n_811)
);

NAND3xp33_ASAP7_75t_L g812 ( 
.A(n_805),
.B(n_771),
.C(n_749),
.Y(n_812)
);

OR2x2_ASAP7_75t_L g813 ( 
.A(n_788),
.B(n_766),
.Y(n_813)
);

AND2x2_ASAP7_75t_L g814 ( 
.A(n_782),
.B(n_776),
.Y(n_814)
);

NAND3xp33_ASAP7_75t_L g815 ( 
.A(n_781),
.B(n_751),
.C(n_754),
.Y(n_815)
);

OR2x2_ASAP7_75t_L g816 ( 
.A(n_791),
.B(n_93),
.Y(n_816)
);

INVx2_ASAP7_75t_L g817 ( 
.A(n_787),
.Y(n_817)
);

NAND3xp33_ASAP7_75t_L g818 ( 
.A(n_783),
.B(n_798),
.C(n_784),
.Y(n_818)
);

NAND3xp33_ASAP7_75t_L g819 ( 
.A(n_784),
.B(n_100),
.C(n_101),
.Y(n_819)
);

AND2x2_ASAP7_75t_L g820 ( 
.A(n_785),
.B(n_102),
.Y(n_820)
);

INVx2_ASAP7_75t_L g821 ( 
.A(n_797),
.Y(n_821)
);

HB1xp67_ASAP7_75t_L g822 ( 
.A(n_792),
.Y(n_822)
);

NAND2xp5_ASAP7_75t_SL g823 ( 
.A(n_796),
.B(n_103),
.Y(n_823)
);

INVx1_ASAP7_75t_L g824 ( 
.A(n_795),
.Y(n_824)
);

NAND4xp25_ASAP7_75t_L g825 ( 
.A(n_785),
.B(n_104),
.C(n_105),
.D(n_106),
.Y(n_825)
);

XNOR2x2_ASAP7_75t_L g826 ( 
.A(n_794),
.B(n_107),
.Y(n_826)
);

INVx1_ASAP7_75t_L g827 ( 
.A(n_808),
.Y(n_827)
);

AND2x2_ASAP7_75t_L g828 ( 
.A(n_822),
.B(n_796),
.Y(n_828)
);

NOR2xp33_ASAP7_75t_SL g829 ( 
.A(n_825),
.B(n_799),
.Y(n_829)
);

INVx1_ASAP7_75t_L g830 ( 
.A(n_808),
.Y(n_830)
);

INVx2_ASAP7_75t_SL g831 ( 
.A(n_822),
.Y(n_831)
);

INVx1_ASAP7_75t_L g832 ( 
.A(n_824),
.Y(n_832)
);

OR2x2_ASAP7_75t_L g833 ( 
.A(n_821),
.B(n_786),
.Y(n_833)
);

XNOR2xp5_ASAP7_75t_L g834 ( 
.A(n_820),
.B(n_814),
.Y(n_834)
);

AND2x2_ASAP7_75t_L g835 ( 
.A(n_807),
.B(n_786),
.Y(n_835)
);

INVx3_ASAP7_75t_L g836 ( 
.A(n_809),
.Y(n_836)
);

NOR4xp25_ASAP7_75t_L g837 ( 
.A(n_818),
.B(n_806),
.C(n_794),
.D(n_801),
.Y(n_837)
);

INVx2_ASAP7_75t_L g838 ( 
.A(n_817),
.Y(n_838)
);

INVx2_ASAP7_75t_L g839 ( 
.A(n_838),
.Y(n_839)
);

XNOR2x1_ASAP7_75t_L g840 ( 
.A(n_834),
.B(n_826),
.Y(n_840)
);

INVx3_ASAP7_75t_L g841 ( 
.A(n_831),
.Y(n_841)
);

XOR2x2_ASAP7_75t_L g842 ( 
.A(n_834),
.B(n_815),
.Y(n_842)
);

INVx1_ASAP7_75t_L g843 ( 
.A(n_827),
.Y(n_843)
);

XOR2x2_ASAP7_75t_L g844 ( 
.A(n_835),
.B(n_811),
.Y(n_844)
);

AOI22xp33_ASAP7_75t_L g845 ( 
.A1(n_840),
.A2(n_842),
.B1(n_844),
.B2(n_829),
.Y(n_845)
);

XOR2x2_ASAP7_75t_L g846 ( 
.A(n_840),
.B(n_835),
.Y(n_846)
);

INVx1_ASAP7_75t_L g847 ( 
.A(n_843),
.Y(n_847)
);

HB1xp67_ASAP7_75t_L g848 ( 
.A(n_841),
.Y(n_848)
);

OA22x2_ASAP7_75t_L g849 ( 
.A1(n_842),
.A2(n_836),
.B1(n_828),
.B2(n_831),
.Y(n_849)
);

INVx1_ASAP7_75t_L g850 ( 
.A(n_847),
.Y(n_850)
);

OAI322xp33_ASAP7_75t_L g851 ( 
.A1(n_849),
.A2(n_836),
.A3(n_830),
.B1(n_832),
.B2(n_841),
.C1(n_828),
.C2(n_833),
.Y(n_851)
);

OAI322xp33_ASAP7_75t_L g852 ( 
.A1(n_849),
.A2(n_836),
.A3(n_833),
.B1(n_823),
.B2(n_839),
.C1(n_838),
.C2(n_837),
.Y(n_852)
);

INVx1_ASAP7_75t_L g853 ( 
.A(n_848),
.Y(n_853)
);

AOI22x1_ASAP7_75t_L g854 ( 
.A1(n_853),
.A2(n_845),
.B1(n_846),
.B2(n_816),
.Y(n_854)
);

INVx1_ASAP7_75t_L g855 ( 
.A(n_850),
.Y(n_855)
);

BUFx4_ASAP7_75t_R g856 ( 
.A(n_851),
.Y(n_856)
);

INVx2_ASAP7_75t_L g857 ( 
.A(n_855),
.Y(n_857)
);

OAI211xp5_ASAP7_75t_SL g858 ( 
.A1(n_856),
.A2(n_852),
.B(n_823),
.C(n_810),
.Y(n_858)
);

OAI22xp33_ASAP7_75t_L g859 ( 
.A1(n_854),
.A2(n_819),
.B1(n_812),
.B2(n_839),
.Y(n_859)
);

INVx1_ASAP7_75t_L g860 ( 
.A(n_855),
.Y(n_860)
);

NOR2x1_ASAP7_75t_L g861 ( 
.A(n_858),
.B(n_800),
.Y(n_861)
);

OA22x2_ASAP7_75t_L g862 ( 
.A1(n_857),
.A2(n_802),
.B1(n_793),
.B2(n_803),
.Y(n_862)
);

NAND2xp5_ASAP7_75t_L g863 ( 
.A(n_860),
.B(n_810),
.Y(n_863)
);

OAI22xp5_ASAP7_75t_SL g864 ( 
.A1(n_859),
.A2(n_790),
.B1(n_813),
.B2(n_804),
.Y(n_864)
);

OR2x6_ASAP7_75t_L g865 ( 
.A(n_857),
.B(n_108),
.Y(n_865)
);

NOR3xp33_ASAP7_75t_L g866 ( 
.A(n_858),
.B(n_110),
.C(n_111),
.Y(n_866)
);

NOR4xp25_ASAP7_75t_L g867 ( 
.A(n_858),
.B(n_112),
.C(n_114),
.D(n_115),
.Y(n_867)
);

NOR2xp33_ASAP7_75t_L g868 ( 
.A(n_863),
.B(n_117),
.Y(n_868)
);

NOR2x1_ASAP7_75t_L g869 ( 
.A(n_861),
.B(n_118),
.Y(n_869)
);

INVx1_ASAP7_75t_L g870 ( 
.A(n_862),
.Y(n_870)
);

INVx1_ASAP7_75t_L g871 ( 
.A(n_865),
.Y(n_871)
);

NAND2xp5_ASAP7_75t_L g872 ( 
.A(n_867),
.B(n_866),
.Y(n_872)
);

NOR2x1_ASAP7_75t_L g873 ( 
.A(n_864),
.B(n_119),
.Y(n_873)
);

AOI22xp5_ASAP7_75t_L g874 ( 
.A1(n_861),
.A2(n_120),
.B1(n_121),
.B2(n_124),
.Y(n_874)
);

NAND4xp25_ASAP7_75t_L g875 ( 
.A(n_870),
.B(n_126),
.C(n_129),
.D(n_130),
.Y(n_875)
);

NAND4xp25_ASAP7_75t_L g876 ( 
.A(n_872),
.B(n_131),
.C(n_132),
.D(n_133),
.Y(n_876)
);

AO22x2_ASAP7_75t_L g877 ( 
.A1(n_871),
.A2(n_134),
.B1(n_135),
.B2(n_136),
.Y(n_877)
);

OR3x2_ASAP7_75t_L g878 ( 
.A(n_869),
.B(n_873),
.C(n_874),
.Y(n_878)
);

INVxp67_ASAP7_75t_SL g879 ( 
.A(n_868),
.Y(n_879)
);

OAI22xp5_ASAP7_75t_L g880 ( 
.A1(n_872),
.A2(n_141),
.B1(n_142),
.B2(n_145),
.Y(n_880)
);

NAND4xp25_ASAP7_75t_L g881 ( 
.A(n_870),
.B(n_146),
.C(n_147),
.D(n_148),
.Y(n_881)
);

INVx1_ASAP7_75t_L g882 ( 
.A(n_879),
.Y(n_882)
);

INVx1_ASAP7_75t_L g883 ( 
.A(n_878),
.Y(n_883)
);

INVxp67_ASAP7_75t_L g884 ( 
.A(n_876),
.Y(n_884)
);

INVx1_ASAP7_75t_L g885 ( 
.A(n_875),
.Y(n_885)
);

INVx2_ASAP7_75t_L g886 ( 
.A(n_877),
.Y(n_886)
);

OAI22xp5_ASAP7_75t_L g887 ( 
.A1(n_880),
.A2(n_150),
.B1(n_152),
.B2(n_154),
.Y(n_887)
);

AND3x1_ASAP7_75t_L g888 ( 
.A(n_881),
.B(n_877),
.C(n_156),
.Y(n_888)
);

INVx1_ASAP7_75t_L g889 ( 
.A(n_879),
.Y(n_889)
);

OAI22xp5_ASAP7_75t_L g890 ( 
.A1(n_882),
.A2(n_155),
.B1(n_159),
.B2(n_160),
.Y(n_890)
);

INVx1_ASAP7_75t_L g891 ( 
.A(n_889),
.Y(n_891)
);

INVx1_ASAP7_75t_L g892 ( 
.A(n_883),
.Y(n_892)
);

AO22x1_ASAP7_75t_L g893 ( 
.A1(n_885),
.A2(n_161),
.B1(n_162),
.B2(n_163),
.Y(n_893)
);

INVx1_ASAP7_75t_SL g894 ( 
.A(n_888),
.Y(n_894)
);

AO22x2_ASAP7_75t_L g895 ( 
.A1(n_886),
.A2(n_164),
.B1(n_165),
.B2(n_166),
.Y(n_895)
);

AOI22xp5_ASAP7_75t_L g896 ( 
.A1(n_884),
.A2(n_167),
.B1(n_170),
.B2(n_171),
.Y(n_896)
);

INVx1_ASAP7_75t_L g897 ( 
.A(n_891),
.Y(n_897)
);

INVx4_ASAP7_75t_L g898 ( 
.A(n_892),
.Y(n_898)
);

HB1xp67_ASAP7_75t_L g899 ( 
.A(n_894),
.Y(n_899)
);

INVx1_ASAP7_75t_L g900 ( 
.A(n_895),
.Y(n_900)
);

AOI22xp5_ASAP7_75t_L g901 ( 
.A1(n_899),
.A2(n_896),
.B1(n_887),
.B2(n_893),
.Y(n_901)
);

OAI22xp33_ASAP7_75t_L g902 ( 
.A1(n_898),
.A2(n_890),
.B1(n_177),
.B2(n_178),
.Y(n_902)
);

OAI221xp5_ASAP7_75t_L g903 ( 
.A1(n_897),
.A2(n_172),
.B1(n_180),
.B2(n_182),
.C(n_183),
.Y(n_903)
);

INVx1_ASAP7_75t_L g904 ( 
.A(n_901),
.Y(n_904)
);

AO22x2_ASAP7_75t_L g905 ( 
.A1(n_904),
.A2(n_898),
.B1(n_900),
.B2(n_902),
.Y(n_905)
);

INVx1_ASAP7_75t_L g906 ( 
.A(n_905),
.Y(n_906)
);

AOI221xp5_ASAP7_75t_L g907 ( 
.A1(n_906),
.A2(n_903),
.B1(n_185),
.B2(n_186),
.C(n_187),
.Y(n_907)
);

AOI211xp5_ASAP7_75t_L g908 ( 
.A1(n_907),
.A2(n_184),
.B(n_192),
.C(n_194),
.Y(n_908)
);


endmodule