module fake_ariane_450_n_2858 (n_295, n_356, n_556, n_170, n_190, n_160, n_64, n_180, n_119, n_124, n_386, n_307, n_516, n_332, n_581, n_294, n_197, n_463, n_176, n_34, n_404, n_172, n_347, n_423, n_183, n_469, n_479, n_373, n_299, n_541, n_499, n_12, n_564, n_133, n_66, n_205, n_341, n_71, n_109, n_245, n_421, n_96, n_549, n_522, n_319, n_49, n_20, n_416, n_283, n_50, n_187, n_525, n_367, n_345, n_374, n_318, n_103, n_244, n_226, n_220, n_261, n_36, n_370, n_189, n_72, n_286, n_443, n_57, n_424, n_528, n_387, n_406, n_117, n_139, n_524, n_85, n_130, n_349, n_391, n_466, n_346, n_214, n_348, n_552, n_2, n_462, n_32, n_410, n_379, n_445, n_515, n_138, n_162, n_264, n_137, n_122, n_198, n_232, n_52, n_441, n_568, n_385, n_73, n_327, n_77, n_372, n_377, n_15, n_396, n_23, n_399, n_554, n_520, n_87, n_279, n_207, n_363, n_354, n_41, n_140, n_419, n_151, n_28, n_146, n_230, n_270, n_194, n_154, n_338, n_142, n_285, n_473, n_186, n_202, n_145, n_193, n_500, n_59, n_336, n_315, n_311, n_239, n_402, n_35, n_272, n_54, n_8, n_339, n_487, n_167, n_90, n_38, n_422, n_47, n_153, n_18, n_269, n_75, n_158, n_69, n_259, n_95, n_446, n_553, n_143, n_566, n_578, n_152, n_405, n_557, n_120, n_169, n_106, n_173, n_242, n_309, n_320, n_115, n_331, n_559, n_401, n_485, n_267, n_495, n_504, n_483, n_335, n_435, n_350, n_291, n_344, n_381, n_426, n_433, n_481, n_398, n_62, n_210, n_200, n_529, n_502, n_166, n_253, n_561, n_218, n_79, n_3, n_271, n_465, n_486, n_507, n_247, n_569, n_567, n_91, n_240, n_369, n_128, n_224, n_44, n_82, n_31, n_547, n_420, n_562, n_518, n_439, n_222, n_478, n_510, n_256, n_326, n_227, n_48, n_188, n_323, n_550, n_330, n_400, n_11, n_129, n_126, n_282, n_328, n_368, n_277, n_248, n_301, n_467, n_432, n_545, n_536, n_293, n_228, n_325, n_276, n_93, n_427, n_108, n_497, n_303, n_442, n_168, n_81, n_1, n_206, n_352, n_538, n_576, n_511, n_238, n_365, n_429, n_455, n_136, n_334, n_192, n_488, n_300, n_533, n_505, n_14, n_163, n_88, n_141, n_390, n_498, n_104, n_501, n_438, n_314, n_16, n_440, n_273, n_305, n_539, n_312, n_233, n_56, n_60, n_388, n_333, n_449, n_413, n_392, n_376, n_512, n_579, n_459, n_221, n_321, n_86, n_361, n_458, n_89, n_149, n_383, n_237, n_175, n_453, n_74, n_491, n_19, n_40, n_181, n_570, n_53, n_260, n_362, n_543, n_310, n_236, n_565, n_281, n_24, n_7, n_461, n_209, n_262, n_490, n_17, n_225, n_235, n_464, n_575, n_546, n_297, n_503, n_290, n_527, n_46, n_84, n_371, n_199, n_107, n_217, n_452, n_178, n_42, n_551, n_308, n_417, n_201, n_70, n_572, n_343, n_10, n_414, n_571, n_287, n_302, n_380, n_6, n_582, n_94, n_284, n_4, n_448, n_249, n_534, n_37, n_58, n_65, n_123, n_212, n_355, n_444, n_278, n_255, n_560, n_450, n_257, n_148, n_451, n_475, n_135, n_409, n_171, n_519, n_384, n_468, n_61, n_526, n_102, n_182, n_482, n_316, n_196, n_125, n_43, n_577, n_407, n_13, n_27, n_254, n_476, n_460, n_219, n_55, n_535, n_231, n_366, n_555, n_234, n_492, n_574, n_280, n_215, n_252, n_161, n_454, n_298, n_532, n_68, n_415, n_78, n_63, n_99, n_540, n_216, n_544, n_5, n_514, n_418, n_537, n_223, n_403, n_25, n_83, n_389, n_513, n_288, n_179, n_395, n_195, n_213, n_110, n_304, n_67, n_509, n_306, n_313, n_92, n_430, n_493, n_203, n_378, n_436, n_150, n_98, n_375, n_113, n_114, n_33, n_324, n_337, n_437, n_111, n_21, n_274, n_472, n_296, n_265, n_208, n_456, n_156, n_292, n_174, n_275, n_100, n_132, n_147, n_204, n_521, n_51, n_496, n_76, n_342, n_26, n_246, n_517, n_530, n_0, n_428, n_159, n_358, n_105, n_580, n_30, n_494, n_131, n_263, n_434, n_360, n_563, n_229, n_394, n_250, n_165, n_144, n_317, n_101, n_243, n_134, n_329, n_185, n_340, n_289, n_9, n_112, n_45, n_542, n_548, n_523, n_268, n_266, n_470, n_457, n_164, n_157, n_184, n_177, n_477, n_364, n_258, n_425, n_431, n_508, n_118, n_121, n_411, n_484, n_353, n_22, n_241, n_29, n_357, n_412, n_447, n_191, n_382, n_489, n_80, n_480, n_211, n_97, n_408, n_322, n_251, n_506, n_558, n_116, n_397, n_471, n_351, n_39, n_393, n_474, n_359, n_155, n_573, n_127, n_531, n_2858);

input n_295;
input n_356;
input n_556;
input n_170;
input n_190;
input n_160;
input n_64;
input n_180;
input n_119;
input n_124;
input n_386;
input n_307;
input n_516;
input n_332;
input n_581;
input n_294;
input n_197;
input n_463;
input n_176;
input n_34;
input n_404;
input n_172;
input n_347;
input n_423;
input n_183;
input n_469;
input n_479;
input n_373;
input n_299;
input n_541;
input n_499;
input n_12;
input n_564;
input n_133;
input n_66;
input n_205;
input n_341;
input n_71;
input n_109;
input n_245;
input n_421;
input n_96;
input n_549;
input n_522;
input n_319;
input n_49;
input n_20;
input n_416;
input n_283;
input n_50;
input n_187;
input n_525;
input n_367;
input n_345;
input n_374;
input n_318;
input n_103;
input n_244;
input n_226;
input n_220;
input n_261;
input n_36;
input n_370;
input n_189;
input n_72;
input n_286;
input n_443;
input n_57;
input n_424;
input n_528;
input n_387;
input n_406;
input n_117;
input n_139;
input n_524;
input n_85;
input n_130;
input n_349;
input n_391;
input n_466;
input n_346;
input n_214;
input n_348;
input n_552;
input n_2;
input n_462;
input n_32;
input n_410;
input n_379;
input n_445;
input n_515;
input n_138;
input n_162;
input n_264;
input n_137;
input n_122;
input n_198;
input n_232;
input n_52;
input n_441;
input n_568;
input n_385;
input n_73;
input n_327;
input n_77;
input n_372;
input n_377;
input n_15;
input n_396;
input n_23;
input n_399;
input n_554;
input n_520;
input n_87;
input n_279;
input n_207;
input n_363;
input n_354;
input n_41;
input n_140;
input n_419;
input n_151;
input n_28;
input n_146;
input n_230;
input n_270;
input n_194;
input n_154;
input n_338;
input n_142;
input n_285;
input n_473;
input n_186;
input n_202;
input n_145;
input n_193;
input n_500;
input n_59;
input n_336;
input n_315;
input n_311;
input n_239;
input n_402;
input n_35;
input n_272;
input n_54;
input n_8;
input n_339;
input n_487;
input n_167;
input n_90;
input n_38;
input n_422;
input n_47;
input n_153;
input n_18;
input n_269;
input n_75;
input n_158;
input n_69;
input n_259;
input n_95;
input n_446;
input n_553;
input n_143;
input n_566;
input n_578;
input n_152;
input n_405;
input n_557;
input n_120;
input n_169;
input n_106;
input n_173;
input n_242;
input n_309;
input n_320;
input n_115;
input n_331;
input n_559;
input n_401;
input n_485;
input n_267;
input n_495;
input n_504;
input n_483;
input n_335;
input n_435;
input n_350;
input n_291;
input n_344;
input n_381;
input n_426;
input n_433;
input n_481;
input n_398;
input n_62;
input n_210;
input n_200;
input n_529;
input n_502;
input n_166;
input n_253;
input n_561;
input n_218;
input n_79;
input n_3;
input n_271;
input n_465;
input n_486;
input n_507;
input n_247;
input n_569;
input n_567;
input n_91;
input n_240;
input n_369;
input n_128;
input n_224;
input n_44;
input n_82;
input n_31;
input n_547;
input n_420;
input n_562;
input n_518;
input n_439;
input n_222;
input n_478;
input n_510;
input n_256;
input n_326;
input n_227;
input n_48;
input n_188;
input n_323;
input n_550;
input n_330;
input n_400;
input n_11;
input n_129;
input n_126;
input n_282;
input n_328;
input n_368;
input n_277;
input n_248;
input n_301;
input n_467;
input n_432;
input n_545;
input n_536;
input n_293;
input n_228;
input n_325;
input n_276;
input n_93;
input n_427;
input n_108;
input n_497;
input n_303;
input n_442;
input n_168;
input n_81;
input n_1;
input n_206;
input n_352;
input n_538;
input n_576;
input n_511;
input n_238;
input n_365;
input n_429;
input n_455;
input n_136;
input n_334;
input n_192;
input n_488;
input n_300;
input n_533;
input n_505;
input n_14;
input n_163;
input n_88;
input n_141;
input n_390;
input n_498;
input n_104;
input n_501;
input n_438;
input n_314;
input n_16;
input n_440;
input n_273;
input n_305;
input n_539;
input n_312;
input n_233;
input n_56;
input n_60;
input n_388;
input n_333;
input n_449;
input n_413;
input n_392;
input n_376;
input n_512;
input n_579;
input n_459;
input n_221;
input n_321;
input n_86;
input n_361;
input n_458;
input n_89;
input n_149;
input n_383;
input n_237;
input n_175;
input n_453;
input n_74;
input n_491;
input n_19;
input n_40;
input n_181;
input n_570;
input n_53;
input n_260;
input n_362;
input n_543;
input n_310;
input n_236;
input n_565;
input n_281;
input n_24;
input n_7;
input n_461;
input n_209;
input n_262;
input n_490;
input n_17;
input n_225;
input n_235;
input n_464;
input n_575;
input n_546;
input n_297;
input n_503;
input n_290;
input n_527;
input n_46;
input n_84;
input n_371;
input n_199;
input n_107;
input n_217;
input n_452;
input n_178;
input n_42;
input n_551;
input n_308;
input n_417;
input n_201;
input n_70;
input n_572;
input n_343;
input n_10;
input n_414;
input n_571;
input n_287;
input n_302;
input n_380;
input n_6;
input n_582;
input n_94;
input n_284;
input n_4;
input n_448;
input n_249;
input n_534;
input n_37;
input n_58;
input n_65;
input n_123;
input n_212;
input n_355;
input n_444;
input n_278;
input n_255;
input n_560;
input n_450;
input n_257;
input n_148;
input n_451;
input n_475;
input n_135;
input n_409;
input n_171;
input n_519;
input n_384;
input n_468;
input n_61;
input n_526;
input n_102;
input n_182;
input n_482;
input n_316;
input n_196;
input n_125;
input n_43;
input n_577;
input n_407;
input n_13;
input n_27;
input n_254;
input n_476;
input n_460;
input n_219;
input n_55;
input n_535;
input n_231;
input n_366;
input n_555;
input n_234;
input n_492;
input n_574;
input n_280;
input n_215;
input n_252;
input n_161;
input n_454;
input n_298;
input n_532;
input n_68;
input n_415;
input n_78;
input n_63;
input n_99;
input n_540;
input n_216;
input n_544;
input n_5;
input n_514;
input n_418;
input n_537;
input n_223;
input n_403;
input n_25;
input n_83;
input n_389;
input n_513;
input n_288;
input n_179;
input n_395;
input n_195;
input n_213;
input n_110;
input n_304;
input n_67;
input n_509;
input n_306;
input n_313;
input n_92;
input n_430;
input n_493;
input n_203;
input n_378;
input n_436;
input n_150;
input n_98;
input n_375;
input n_113;
input n_114;
input n_33;
input n_324;
input n_337;
input n_437;
input n_111;
input n_21;
input n_274;
input n_472;
input n_296;
input n_265;
input n_208;
input n_456;
input n_156;
input n_292;
input n_174;
input n_275;
input n_100;
input n_132;
input n_147;
input n_204;
input n_521;
input n_51;
input n_496;
input n_76;
input n_342;
input n_26;
input n_246;
input n_517;
input n_530;
input n_0;
input n_428;
input n_159;
input n_358;
input n_105;
input n_580;
input n_30;
input n_494;
input n_131;
input n_263;
input n_434;
input n_360;
input n_563;
input n_229;
input n_394;
input n_250;
input n_165;
input n_144;
input n_317;
input n_101;
input n_243;
input n_134;
input n_329;
input n_185;
input n_340;
input n_289;
input n_9;
input n_112;
input n_45;
input n_542;
input n_548;
input n_523;
input n_268;
input n_266;
input n_470;
input n_457;
input n_164;
input n_157;
input n_184;
input n_177;
input n_477;
input n_364;
input n_258;
input n_425;
input n_431;
input n_508;
input n_118;
input n_121;
input n_411;
input n_484;
input n_353;
input n_22;
input n_241;
input n_29;
input n_357;
input n_412;
input n_447;
input n_191;
input n_382;
input n_489;
input n_80;
input n_480;
input n_211;
input n_97;
input n_408;
input n_322;
input n_251;
input n_506;
input n_558;
input n_116;
input n_397;
input n_471;
input n_351;
input n_39;
input n_393;
input n_474;
input n_359;
input n_155;
input n_573;
input n_127;
input n_531;

output n_2858;

wire n_2752;
wire n_913;
wire n_1681;
wire n_2163;
wire n_1486;
wire n_1507;
wire n_1938;
wire n_589;
wire n_2484;
wire n_1174;
wire n_2346;
wire n_1469;
wire n_691;
wire n_1353;
wire n_2679;
wire n_1355;
wire n_2131;
wire n_2559;
wire n_2500;
wire n_2509;
wire n_1383;
wire n_2182;
wire n_603;
wire n_2135;
wire n_2334;
wire n_2680;
wire n_1250;
wire n_2030;
wire n_1169;
wire n_789;
wire n_850;
wire n_1916;
wire n_610;
wire n_1713;
wire n_1436;
wire n_2407;
wire n_690;
wire n_2818;
wire n_1109;
wire n_1430;
wire n_2537;
wire n_2002;
wire n_1463;
wire n_2243;
wire n_1238;
wire n_2694;
wire n_2011;
wire n_2729;
wire n_1515;
wire n_817;
wire n_1837;
wire n_924;
wire n_781;
wire n_2013;
wire n_2786;
wire n_1566;
wire n_2837;
wire n_717;
wire n_2006;
wire n_952;
wire n_864;
wire n_2446;
wire n_1096;
wire n_1379;
wire n_2436;
wire n_2376;
wire n_2367;
wire n_2671;
wire n_2790;
wire n_1706;
wire n_2207;
wire n_2461;
wire n_2702;
wire n_2731;
wire n_634;
wire n_1214;
wire n_1839;
wire n_1246;
wire n_1138;
wire n_2042;
wire n_2123;
wire n_1853;
wire n_764;
wire n_1503;
wire n_2238;
wire n_2529;
wire n_2374;
wire n_1196;
wire n_1181;
wire n_1999;
wire n_2380;
wire n_1187;
wire n_1131;
wire n_1225;
wire n_2646;
wire n_737;
wire n_1298;
wire n_2653;
wire n_1745;
wire n_1366;
wire n_2084;
wire n_2278;
wire n_1088;
wire n_1424;
wire n_766;
wire n_1835;
wire n_1457;
wire n_2482;
wire n_1682;
wire n_2750;
wire n_1836;
wire n_870;
wire n_2547;
wire n_1453;
wire n_945;
wire n_958;
wire n_2554;
wire n_2248;
wire n_813;
wire n_1985;
wire n_2288;
wire n_2621;
wire n_995;
wire n_2579;
wire n_1909;
wire n_2156;
wire n_1184;
wire n_1961;
wire n_1535;
wire n_754;
wire n_665;
wire n_903;
wire n_871;
wire n_2323;
wire n_1073;
wire n_2844;
wire n_1979;
wire n_1277;
wire n_2107;
wire n_1746;
wire n_829;
wire n_1761;
wire n_1062;
wire n_738;
wire n_1690;
wire n_2221;
wire n_2807;
wire n_672;
wire n_740;
wire n_1283;
wire n_2317;
wire n_2838;
wire n_1974;
wire n_1736;
wire n_1018;
wire n_2342;
wire n_2200;
wire n_2781;
wire n_2442;
wire n_2735;
wire n_953;
wire n_1364;
wire n_2390;
wire n_1888;
wire n_1224;
wire n_2109;
wire n_1425;
wire n_2634;
wire n_2709;
wire n_625;
wire n_2322;
wire n_2746;
wire n_1107;
wire n_2832;
wire n_1688;
wire n_989;
wire n_645;
wire n_1944;
wire n_2370;
wire n_2233;
wire n_2663;
wire n_1988;
wire n_795;
wire n_721;
wire n_1084;
wire n_1718;
wire n_1276;
wire n_1936;
wire n_2149;
wire n_2277;
wire n_1428;
wire n_1284;
wire n_1241;
wire n_821;
wire n_770;
wire n_1514;
wire n_2539;
wire n_1528;
wire n_901;
wire n_2782;
wire n_2078;
wire n_1145;
wire n_971;
wire n_2359;
wire n_2201;
wire n_787;
wire n_1650;
wire n_1519;
wire n_1195;
wire n_2049;
wire n_1522;
wire n_1207;
wire n_786;
wire n_1404;
wire n_868;
wire n_2232;
wire n_1847;
wire n_2458;
wire n_2779;
wire n_1542;
wire n_1314;
wire n_1512;
wire n_2227;
wire n_2301;
wire n_1539;
wire n_2847;
wire n_884;
wire n_1851;
wire n_2162;
wire n_1415;
wire n_1034;
wire n_1652;
wire n_2192;
wire n_1676;
wire n_1085;
wire n_1636;
wire n_823;
wire n_1900;
wire n_620;
wire n_1074;
wire n_859;
wire n_1765;
wire n_1889;
wire n_587;
wire n_1977;
wire n_693;
wire n_863;
wire n_2650;
wire n_1254;
wire n_929;
wire n_2433;
wire n_1703;
wire n_899;
wire n_2332;
wire n_2391;
wire n_611;
wire n_1295;
wire n_2060;
wire n_1850;
wire n_2004;
wire n_1013;
wire n_1495;
wire n_1637;
wire n_2571;
wire n_2427;
wire n_661;
wire n_2098;
wire n_2616;
wire n_1751;
wire n_1917;
wire n_2456;
wire n_2769;
wire n_1924;
wire n_1560;
wire n_1654;
wire n_2341;
wire n_1548;
wire n_1811;
wire n_2045;
wire n_2575;
wire n_2722;
wire n_1396;
wire n_1230;
wire n_612;
wire n_1840;
wire n_2739;
wire n_1597;
wire n_1771;
wire n_1544;
wire n_844;
wire n_1012;
wire n_1267;
wire n_2061;
wire n_2685;
wire n_2094;
wire n_2512;
wire n_1354;
wire n_1790;
wire n_1213;
wire n_2382;
wire n_2043;
wire n_780;
wire n_2349;
wire n_1918;
wire n_2788;
wire n_1021;
wire n_1443;
wire n_2595;
wire n_1465;
wire n_2686;
wire n_1949;
wire n_1595;
wire n_1142;
wire n_1140;
wire n_705;
wire n_2727;
wire n_942;
wire n_1437;
wire n_2077;
wire n_1378;
wire n_1121;
wire n_1416;
wire n_1461;
wire n_2717;
wire n_1391;
wire n_1947;
wire n_1599;
wire n_1876;
wire n_1006;
wire n_1830;
wire n_2527;
wire n_1112;
wire n_700;
wire n_1159;
wire n_772;
wire n_1216;
wire n_2759;
wire n_1245;
wire n_2743;
wire n_1669;
wire n_1675;
wire n_2466;
wire n_676;
wire n_2038;
wire n_2263;
wire n_2800;
wire n_2568;
wire n_2116;
wire n_2271;
wire n_2145;
wire n_2326;
wire n_1838;
wire n_1594;
wire n_680;
wire n_1935;
wire n_2806;
wire n_1716;
wire n_1872;
wire n_1585;
wire n_2281;
wire n_1432;
wire n_2245;
wire n_1108;
wire n_851;
wire n_1590;
wire n_1351;
wire n_2216;
wire n_1274;
wire n_2426;
wire n_652;
wire n_1819;
wire n_947;
wire n_2134;
wire n_930;
wire n_1260;
wire n_1179;
wire n_2703;
wire n_696;
wire n_1442;
wire n_2620;
wire n_798;
wire n_1833;
wire n_1691;
wire n_916;
wire n_1386;
wire n_2810;
wire n_912;
wire n_1884;
wire n_1555;
wire n_1842;
wire n_2499;
wire n_2549;
wire n_762;
wire n_1253;
wire n_1468;
wire n_1661;
wire n_2791;
wire n_2683;
wire n_804;
wire n_1656;
wire n_1382;
wire n_992;
wire n_966;
wire n_955;
wire n_1182;
wire n_794;
wire n_2855;
wire n_2166;
wire n_2848;
wire n_1692;
wire n_2611;
wire n_1562;
wire n_2748;
wire n_2185;
wire n_2398;
wire n_1376;
wire n_1292;
wire n_1178;
wire n_1972;
wire n_2015;
wire n_1435;
wire n_1750;
wire n_1026;
wire n_1506;
wire n_1610;
wire n_2202;
wire n_2072;
wire n_2415;
wire n_2693;
wire n_2745;
wire n_2087;
wire n_931;
wire n_669;
wire n_1491;
wire n_2628;
wire n_619;
wire n_967;
wire n_1083;
wire n_2161;
wire n_1418;
wire n_746;
wire n_1357;
wire n_1079;
wire n_1787;
wire n_2462;
wire n_1389;
wire n_2155;
wire n_2659;
wire n_615;
wire n_1139;
wire n_2836;
wire n_2439;
wire n_1312;
wire n_1717;
wire n_1812;
wire n_824;
wire n_2172;
wire n_2601;
wire n_892;
wire n_1880;
wire n_959;
wire n_2365;
wire n_2257;
wire n_1399;
wire n_1101;
wire n_1567;
wire n_1343;
wire n_2219;
wire n_1855;
wire n_2100;
wire n_2333;
wire n_990;
wire n_1623;
wire n_1903;
wire n_867;
wire n_2147;
wire n_2435;
wire n_1226;
wire n_2224;
wire n_944;
wire n_749;
wire n_1932;
wire n_1780;
wire n_2825;
wire n_1970;
wire n_1920;
wire n_2083;
wire n_815;
wire n_2167;
wire n_2293;
wire n_2753;
wire n_1340;
wire n_2668;
wire n_1240;
wire n_1087;
wire n_2701;
wire n_2400;
wire n_632;
wire n_650;
wire n_2388;
wire n_2273;
wire n_2712;
wire n_1433;
wire n_1911;
wire n_2567;
wire n_2557;
wire n_2695;
wire n_1825;
wire n_1908;
wire n_1155;
wire n_2598;
wire n_1071;
wire n_2755;
wire n_712;
wire n_976;
wire n_909;
wire n_1392;
wire n_767;
wire n_1832;
wire n_2795;
wire n_2682;
wire n_1841;
wire n_1680;
wire n_2066;
wire n_2302;
wire n_2762;
wire n_964;
wire n_1627;
wire n_2220;
wire n_2294;
wire n_2274;
wire n_974;
wire n_1731;
wire n_799;
wire n_1147;
wire n_2829;
wire n_2378;
wire n_2467;
wire n_2768;
wire n_965;
wire n_1914;
wire n_2253;
wire n_934;
wire n_2213;
wire n_1447;
wire n_2363;
wire n_1220;
wire n_2019;
wire n_698;
wire n_2728;
wire n_2130;
wire n_1674;
wire n_2021;
wire n_2025;
wire n_2160;
wire n_1992;
wire n_1209;
wire n_1020;
wire n_1563;
wire n_646;
wire n_2507;
wire n_2142;
wire n_1633;
wire n_2625;
wire n_1913;
wire n_2069;
wire n_2495;
wire n_1058;
wire n_2328;
wire n_2434;
wire n_1042;
wire n_1234;
wire n_2311;
wire n_1578;
wire n_2261;
wire n_1455;
wire n_2287;
wire n_836;
wire n_2223;
wire n_1279;
wire n_2473;
wire n_2144;
wire n_2511;
wire n_1029;
wire n_2649;
wire n_1247;
wire n_760;
wire n_2438;
wire n_1568;
wire n_1483;
wire n_1363;
wire n_2681;
wire n_1111;
wire n_970;
wire n_1689;
wire n_2535;
wire n_713;
wire n_1255;
wire n_2632;
wire n_1646;
wire n_598;
wire n_2262;
wire n_2565;
wire n_1237;
wire n_927;
wire n_1095;
wire n_1728;
wire n_2335;
wire n_706;
wire n_2120;
wire n_2631;
wire n_1401;
wire n_1419;
wire n_1531;
wire n_776;
wire n_2041;
wire n_2113;
wire n_1933;
wire n_1651;
wire n_2697;
wire n_1387;
wire n_1263;
wire n_1817;
wire n_2404;
wire n_2168;
wire n_2757;
wire n_2312;
wire n_670;
wire n_2677;
wire n_1826;
wire n_2834;
wire n_2483;
wire n_1951;
wire n_2490;
wire n_1032;
wire n_1217;
wire n_2558;
wire n_1496;
wire n_637;
wire n_1592;
wire n_2812;
wire n_2662;
wire n_1259;
wire n_2801;
wire n_1177;
wire n_2655;
wire n_1231;
wire n_2132;
wire n_980;
wire n_1618;
wire n_1869;
wire n_1743;
wire n_905;
wire n_2718;
wire n_720;
wire n_926;
wire n_1943;
wire n_2687;
wire n_2296;
wire n_1802;
wire n_2178;
wire n_2112;
wire n_2765;
wire n_1163;
wire n_2640;
wire n_2811;
wire n_1795;
wire n_1384;
wire n_2237;
wire n_2146;
wire n_1868;
wire n_1501;
wire n_2241;
wire n_2373;
wire n_1173;
wire n_2350;
wire n_1068;
wire n_1198;
wire n_2531;
wire n_1570;
wire n_2099;
wire n_1518;
wire n_1456;
wire n_1879;
wire n_1886;
wire n_1648;
wire n_2187;
wire n_1413;
wire n_2617;
wire n_2481;
wire n_2129;
wire n_855;
wire n_2327;
wire n_808;
wire n_1365;
wire n_2476;
wire n_2814;
wire n_2059;
wire n_2437;
wire n_2636;
wire n_1439;
wire n_814;
wire n_2074;
wire n_1665;
wire n_1287;
wire n_2841;
wire n_1611;
wire n_2122;
wire n_2399;
wire n_1414;
wire n_1134;
wire n_2067;
wire n_1484;
wire n_1901;
wire n_647;
wire n_2055;
wire n_2027;
wire n_1423;
wire n_2117;
wire n_600;
wire n_1053;
wire n_1609;
wire n_2822;
wire n_1939;
wire n_2308;
wire n_2242;
wire n_1906;
wire n_1899;
wire n_2195;
wire n_2194;
wire n_1467;
wire n_1828;
wire n_2159;
wire n_1798;
wire n_1304;
wire n_1608;
wire n_1744;
wire n_2267;
wire n_1105;
wire n_677;
wire n_604;
wire n_703;
wire n_1349;
wire n_1709;
wire n_1061;
wire n_2102;
wire n_681;
wire n_874;
wire n_2286;
wire n_2023;
wire n_1278;
wire n_707;
wire n_983;
wire n_2783;
wire n_2599;
wire n_699;
wire n_590;
wire n_727;
wire n_2075;
wire n_1726;
wire n_2523;
wire n_1945;
wire n_1015;
wire n_2418;
wire n_1377;
wire n_1162;
wire n_1614;
wire n_2031;
wire n_2496;
wire n_2118;
wire n_1740;
wire n_1602;
wire n_688;
wire n_636;
wire n_2853;
wire n_1098;
wire n_1490;
wire n_2338;
wire n_777;
wire n_1553;
wire n_1080;
wire n_920;
wire n_1760;
wire n_1086;
wire n_1092;
wire n_2225;
wire n_986;
wire n_1104;
wire n_1963;
wire n_2802;
wire n_729;
wire n_887;
wire n_2057;
wire n_2218;
wire n_1122;
wire n_1205;
wire n_1408;
wire n_2593;
wire n_1693;
wire n_2125;
wire n_2716;
wire n_1132;
wire n_1156;
wire n_2741;
wire n_2184;
wire n_2714;
wire n_1823;
wire n_2780;
wire n_1120;
wire n_1202;
wire n_627;
wire n_2254;
wire n_1188;
wire n_1498;
wire n_1371;
wire n_2033;
wire n_2618;
wire n_957;
wire n_1402;
wire n_1242;
wire n_2754;
wire n_2707;
wire n_2774;
wire n_2849;
wire n_1607;
wire n_1489;
wire n_2799;
wire n_1218;
wire n_2756;
wire n_2217;
wire n_2226;
wire n_1586;
wire n_861;
wire n_1543;
wire n_1431;
wire n_877;
wire n_1119;
wire n_1863;
wire n_1763;
wire n_1666;
wire n_1500;
wire n_616;
wire n_2214;
wire n_1055;
wire n_1395;
wire n_1346;
wire n_2763;
wire n_2256;
wire n_1189;
wire n_1089;
wire n_1859;
wire n_2660;
wire n_1502;
wire n_1523;
wire n_2190;
wire n_1478;
wire n_2732;
wire n_1883;
wire n_2516;
wire n_2776;
wire n_2555;
wire n_1969;
wire n_2708;
wire n_735;
wire n_1005;
wire n_2379;
wire n_1294;
wire n_2661;
wire n_1667;
wire n_845;
wire n_888;
wire n_2300;
wire n_1649;
wire n_2452;
wire n_1677;
wire n_2470;
wire n_1927;
wire n_1297;
wire n_2827;
wire n_1708;
wire n_1222;
wire n_2284;
wire n_1844;
wire n_2283;
wire n_2526;
wire n_1957;
wire n_1953;
wire n_2643;
wire n_755;
wire n_1097;
wire n_1219;
wire n_1711;
wire n_710;
wire n_1919;
wire n_1791;
wire n_2508;
wire n_2124;
wire n_1894;
wire n_1460;
wire n_1239;
wire n_2594;
wire n_2266;
wire n_2449;
wire n_890;
wire n_842;
wire n_1898;
wire n_1741;
wire n_745;
wire n_1572;
wire n_1907;
wire n_1793;
wire n_742;
wire n_1373;
wire n_1081;
wire n_1975;
wire n_1388;
wire n_1266;
wire n_1540;
wire n_1719;
wire n_2119;
wire n_2742;
wire n_769;
wire n_1797;
wire n_2366;
wire n_2493;
wire n_1753;
wire n_1990;
wire n_1372;
wire n_832;
wire n_744;
wire n_1895;
wire n_2821;
wire n_2690;
wire n_2474;
wire n_2623;
wire n_982;
wire n_1800;
wire n_915;
wire n_1075;
wire n_2008;
wire n_1331;
wire n_1890;
wire n_1529;
wire n_1227;
wire n_2127;
wire n_655;
wire n_1860;
wire n_1734;
wire n_2785;
wire n_2460;
wire n_2840;
wire n_1007;
wire n_1580;
wire n_1319;
wire n_657;
wire n_837;
wire n_812;
wire n_2448;
wire n_2211;
wire n_2292;
wire n_2480;
wire n_606;
wire n_951;
wire n_2772;
wire n_862;
wire n_1700;
wire n_2637;
wire n_659;
wire n_1332;
wire n_2306;
wire n_1854;
wire n_666;
wire n_1747;
wire n_2071;
wire n_2424;
wire n_1206;
wire n_1729;
wire n_722;
wire n_1508;
wire n_2414;
wire n_2082;
wire n_1532;
wire n_1171;
wire n_1030;
wire n_785;
wire n_2389;
wire n_1309;
wire n_999;
wire n_2280;
wire n_1766;
wire n_1338;
wire n_1342;
wire n_2737;
wire n_1867;
wire n_852;
wire n_1394;
wire n_2576;
wire n_704;
wire n_1060;
wire n_1044;
wire n_1714;
wire n_2696;
wire n_2140;
wire n_873;
wire n_1301;
wire n_1748;
wire n_2157;
wire n_1966;
wire n_1243;
wire n_2171;
wire n_2468;
wire n_1400;
wire n_2035;
wire n_2614;
wire n_1466;
wire n_1527;
wire n_1513;
wire n_2581;
wire n_1783;
wire n_608;
wire n_2494;
wire n_1538;
wire n_2831;
wire n_2457;
wire n_2128;
wire n_1037;
wire n_1329;
wire n_1993;
wire n_1545;
wire n_2629;
wire n_1257;
wire n_1480;
wire n_1954;
wire n_1668;
wire n_1878;
wire n_2540;
wire n_1605;
wire n_1078;
wire n_2486;
wire n_1897;
wire n_2520;
wire n_2137;
wire n_1161;
wire n_2489;
wire n_811;
wire n_624;
wire n_876;
wire n_791;
wire n_1191;
wire n_618;
wire n_2492;
wire n_736;
wire n_1025;
wire n_1215;
wire n_1449;
wire n_2337;
wire n_2265;
wire n_687;
wire n_797;
wire n_2026;
wire n_1786;
wire n_2627;
wire n_1327;
wire n_1475;
wire n_642;
wire n_1804;
wire n_2106;
wire n_1406;
wire n_595;
wire n_1405;
wire n_2684;
wire n_2726;
wire n_602;
wire n_2622;
wire n_2272;
wire n_1757;
wire n_592;
wire n_1499;
wire n_854;
wire n_1318;
wire n_2091;
wire n_1632;
wire n_1769;
wire n_1929;
wire n_1950;
wire n_2264;
wire n_2691;
wire n_805;
wire n_2032;
wire n_2090;
wire n_1658;
wire n_2249;
wire n_1072;
wire n_695;
wire n_1526;
wire n_1305;
wire n_730;
wire n_1596;
wire n_2348;
wire n_2656;
wire n_1281;
wire n_2574;
wire n_2364;
wire n_1997;
wire n_1137;
wire n_1873;
wire n_1258;
wire n_640;
wire n_1733;
wire n_1476;
wire n_1524;
wire n_1856;
wire n_2016;
wire n_2667;
wire n_2723;
wire n_2725;
wire n_943;
wire n_1118;
wire n_678;
wire n_651;
wire n_2850;
wire n_1874;
wire n_1293;
wire n_961;
wire n_1046;
wire n_1807;
wire n_1123;
wire n_726;
wire n_1657;
wire n_878;
wire n_2857;
wire n_1784;
wire n_771;
wire n_1321;
wire n_752;
wire n_2307;
wire n_1488;
wire n_985;
wire n_1330;
wire n_906;
wire n_1180;
wire n_1697;
wire n_2295;
wire n_2730;
wire n_806;
wire n_1984;
wire n_1350;
wire n_1556;
wire n_649;
wire n_1561;
wire n_2412;
wire n_2720;
wire n_1352;
wire n_2405;
wire n_2815;
wire n_1824;
wire n_643;
wire n_2606;
wire n_2700;
wire n_1492;
wire n_2383;
wire n_2764;
wire n_1441;
wire n_1822;
wire n_682;
wire n_1616;
wire n_2633;
wire n_2416;
wire n_819;
wire n_2386;
wire n_1971;
wire n_586;
wire n_1324;
wire n_1429;
wire n_2064;
wire n_2353;
wire n_2528;
wire n_1778;
wire n_1776;
wire n_686;
wire n_605;
wire n_1154;
wire n_584;
wire n_1557;
wire n_1759;
wire n_1829;
wire n_2325;
wire n_1130;
wire n_1450;
wire n_756;
wire n_2022;
wire n_1016;
wire n_2298;
wire n_1149;
wire n_1505;
wire n_2408;
wire n_2698;
wire n_2320;
wire n_979;
wire n_2329;
wire n_2570;
wire n_1642;
wire n_2417;
wire n_2789;
wire n_2525;
wire n_1815;
wire n_2813;
wire n_897;
wire n_2546;
wire n_949;
wire n_2454;
wire n_1493;
wire n_807;
wire n_891;
wire n_885;
wire n_1659;
wire n_2354;
wire n_1864;
wire n_2760;
wire n_1887;
wire n_1208;
wire n_1987;
wire n_2368;
wire n_802;
wire n_1151;
wire n_960;
wire n_2352;
wire n_2502;
wire n_1256;
wire n_714;
wire n_2170;
wire n_790;
wire n_2244;
wire n_2143;
wire n_2393;
wire n_725;
wire n_2377;
wire n_1577;
wire n_1448;
wire n_2198;
wire n_1009;
wire n_2652;
wire n_1133;
wire n_883;
wire n_1852;
wire n_801;
wire n_1286;
wire n_2612;
wire n_818;
wire n_1685;
wire n_779;
wire n_2410;
wire n_2314;
wire n_2477;
wire n_2279;
wire n_594;
wire n_2222;
wire n_1995;
wire n_1877;
wire n_1397;
wire n_1052;
wire n_1333;
wire n_1306;
wire n_1849;
wire n_2076;
wire n_2133;
wire n_2203;
wire n_833;
wire n_1426;
wire n_2250;
wire n_2497;
wire n_2247;
wire n_2230;
wire n_879;
wire n_1117;
wire n_1269;
wire n_1303;
wire n_1547;
wire n_1438;
wire n_1541;
wire n_597;
wire n_2001;
wire n_1047;
wire n_2506;
wire n_1472;
wire n_2413;
wire n_1593;
wire n_2610;
wire n_1050;
wire n_2626;
wire n_2158;
wire n_2578;
wire n_2607;
wire n_2285;
wire n_1201;
wire n_1288;
wire n_2605;
wire n_858;
wire n_2796;
wire n_1185;
wire n_2475;
wire n_2804;
wire n_2173;
wire n_2715;
wire n_1035;
wire n_1143;
wire n_2665;
wire n_2070;
wire n_2136;
wire n_2771;
wire n_1090;
wire n_2403;
wire n_1367;
wire n_2044;
wire n_928;
wire n_1153;
wire n_1103;
wire n_825;
wire n_732;
wire n_2619;
wire n_1565;
wire n_1192;
wire n_894;
wire n_1380;
wire n_1624;
wire n_1801;
wire n_2854;
wire n_1291;
wire n_2020;
wire n_748;
wire n_2310;
wire n_1045;
wire n_1160;
wire n_1882;
wire n_1976;
wire n_1023;
wire n_2711;
wire n_1881;
wire n_2635;
wire n_988;
wire n_914;
wire n_689;
wire n_1116;
wire n_1958;
wire n_2747;
wire n_1511;
wire n_2177;
wire n_2713;
wire n_1422;
wire n_2766;
wire n_1965;
wire n_644;
wire n_1197;
wire n_2820;
wire n_2613;
wire n_1165;
wire n_1641;
wire n_2845;
wire n_1517;
wire n_2036;
wire n_843;
wire n_2647;
wire n_588;
wire n_638;
wire n_2003;
wire n_2533;
wire n_2210;
wire n_1307;
wire n_1128;
wire n_2053;
wire n_1671;
wire n_1417;
wire n_1048;
wire n_2343;
wire n_775;
wire n_667;
wire n_2419;
wire n_1049;
wire n_2330;
wire n_2826;
wire n_869;
wire n_846;
wire n_1398;
wire n_1921;
wire n_2777;
wire n_2450;
wire n_2411;
wire n_1356;
wire n_1341;
wire n_2234;
wire n_2309;
wire n_1504;
wire n_1955;
wire n_2110;
wire n_2431;
wire n_1773;
wire n_1440;
wire n_2666;
wire n_1370;
wire n_1603;
wire n_728;
wire n_2401;
wire n_715;
wire n_889;
wire n_1066;
wire n_1549;
wire n_2588;
wire n_2331;
wire n_935;
wire n_2478;
wire n_685;
wire n_911;
wire n_2658;
wire n_623;
wire n_2608;
wire n_1712;
wire n_1403;
wire n_1065;
wire n_1534;
wire n_1948;
wire n_2767;
wire n_810;
wire n_1290;
wire n_1959;
wire n_617;
wire n_2396;
wire n_1362;
wire n_1559;
wire n_2121;
wire n_2692;
wire n_601;
wire n_683;
wire n_628;
wire n_1300;
wire n_1960;
wire n_2068;
wire n_743;
wire n_1194;
wire n_1647;
wire n_1546;
wire n_1420;
wire n_2553;
wire n_2645;
wire n_907;
wire n_2749;
wire n_1454;
wire n_2592;
wire n_660;
wire n_2459;
wire n_962;
wire n_941;
wire n_1210;
wire n_847;
wire n_747;
wire n_1622;
wire n_1135;
wire n_2566;
wire n_2751;
wire n_918;
wire n_1968;
wire n_1885;
wire n_639;
wire n_673;
wire n_2842;
wire n_2833;
wire n_2196;
wire n_1038;
wire n_2371;
wire n_1978;
wire n_1521;
wire n_1694;
wire n_1940;
wire n_593;
wire n_1695;
wire n_2560;
wire n_1164;
wire n_2313;
wire n_609;
wire n_1193;
wire n_1345;
wire n_613;
wire n_1022;
wire n_1336;
wire n_1033;
wire n_1774;
wire n_2609;
wire n_2561;
wire n_1166;
wire n_1056;
wire n_2007;
wire n_1994;
wire n_1767;
wire n_1040;
wire n_674;
wire n_1158;
wire n_1973;
wire n_1444;
wire n_1803;
wire n_820;
wire n_1749;
wire n_872;
wire n_1653;
wire n_2303;
wire n_2669;
wire n_1157;
wire n_1584;
wire n_848;
wire n_1664;
wire n_629;
wire n_1739;
wire n_2642;
wire n_1814;
wire n_2154;
wire n_2441;
wire n_2236;
wire n_1789;
wire n_763;
wire n_1986;
wire n_2174;
wire n_2688;
wire n_692;
wire n_2624;
wire n_2054;
wire n_1857;
wire n_2315;
wire n_984;
wire n_1687;
wire n_2073;
wire n_2150;
wire n_1552;
wire n_750;
wire n_834;
wire n_1612;
wire n_2498;
wire n_800;
wire n_2638;
wire n_2046;
wire n_1816;
wire n_1910;
wire n_2803;
wire n_1756;
wire n_1606;
wire n_2189;
wire n_621;
wire n_2648;
wire n_1587;
wire n_2093;
wire n_2340;
wire n_2018;
wire n_2672;
wire n_1772;
wire n_2444;
wire n_2602;
wire n_1014;
wire n_724;
wire n_2204;
wire n_1427;
wire n_1481;
wire n_2040;
wire n_1311;
wire n_2199;
wire n_1956;
wire n_1589;
wire n_2151;
wire n_1100;
wire n_585;
wire n_875;
wire n_1617;
wire n_2455;
wire n_827;
wire n_2600;
wire n_2231;
wire n_697;
wire n_2828;
wire n_622;
wire n_1626;
wire n_1962;
wire n_1335;
wire n_1715;
wire n_2305;
wire n_880;
wire n_793;
wire n_2114;
wire n_1175;
wire n_2289;
wire n_2530;
wire n_2299;
wire n_751;
wire n_1027;
wire n_1070;
wire n_2406;
wire n_1621;
wire n_739;
wire n_1485;
wire n_1028;
wire n_1221;
wire n_1785;
wire n_1262;
wire n_792;
wire n_1942;
wire n_2180;
wire n_1579;
wire n_2809;
wire n_2181;
wire n_2014;
wire n_975;
wire n_1645;
wire n_923;
wire n_1124;
wire n_1381;
wire n_1494;
wire n_932;
wire n_1893;
wire n_1183;
wire n_1326;
wire n_2276;
wire n_1805;
wire n_2282;
wire n_981;
wire n_2141;
wire n_1110;
wire n_1758;
wire n_2503;
wire n_2270;
wire n_2443;
wire n_1407;
wire n_2465;
wire n_1204;
wire n_1554;
wire n_994;
wire n_2428;
wire n_2586;
wire n_1360;
wire n_973;
wire n_972;
wire n_2251;
wire n_2843;
wire n_856;
wire n_2572;
wire n_1248;
wire n_1176;
wire n_1564;
wire n_2010;
wire n_1054;
wire n_1679;
wire n_2126;
wire n_1952;
wire n_2425;
wire n_2394;
wire n_1858;
wire n_1678;
wire n_2589;
wire n_1482;
wire n_1361;
wire n_2356;
wire n_1601;
wire n_1057;
wire n_2487;
wire n_1834;
wire n_978;
wire n_1011;
wire n_1520;
wire n_2534;
wire n_2488;
wire n_1509;
wire n_828;
wire n_1411;
wire n_1359;
wire n_1721;
wire n_2564;
wire n_2591;
wire n_653;
wire n_1445;
wire n_1317;
wire n_2050;
wire n_2197;
wire n_783;
wire n_2550;
wire n_1127;
wire n_1536;
wire n_1471;
wire n_2385;
wire n_2387;
wire n_1008;
wire n_1024;
wire n_830;
wire n_2291;
wire n_2816;
wire n_1980;
wire n_2518;
wire n_987;
wire n_936;
wire n_2510;
wire n_1620;
wire n_2501;
wire n_2542;
wire n_1385;
wire n_1525;
wire n_2793;
wire n_1998;
wire n_2165;
wire n_2675;
wire n_2604;
wire n_1775;
wire n_788;
wire n_908;
wire n_2639;
wire n_1036;
wire n_2169;
wire n_2603;
wire n_1270;
wire n_1167;
wire n_1272;
wire n_2630;
wire n_591;
wire n_2794;
wire n_969;
wire n_2028;
wire n_919;
wire n_1663;
wire n_2092;
wire n_2175;
wire n_1625;
wire n_2086;
wire n_2773;
wire n_2817;
wire n_1926;
wire n_2402;
wire n_1458;
wire n_679;
wire n_1630;
wire n_663;
wire n_1720;
wire n_2409;
wire n_2176;
wire n_1412;
wire n_1738;
wire n_1550;
wire n_1358;
wire n_1200;
wire n_826;
wire n_2808;
wire n_2453;
wire n_2344;
wire n_1922;
wire n_1735;
wire n_1788;
wire n_940;
wire n_2392;
wire n_1537;
wire n_2138;
wire n_2065;
wire n_2543;
wire n_2321;
wire n_1077;
wire n_2597;
wire n_607;
wire n_956;
wire n_1930;
wire n_765;
wire n_1809;
wire n_2787;
wire n_1843;
wire n_1904;
wire n_2000;
wire n_2805;
wire n_1268;
wire n_2676;
wire n_2758;
wire n_2395;
wire n_917;
wire n_1271;
wire n_2096;
wire n_2440;
wire n_2556;
wire n_2186;
wire n_1530;
wire n_2215;
wire n_2770;
wire n_631;
wire n_1170;
wire n_2724;
wire n_2258;
wire n_1261;
wire n_2471;
wire n_702;
wire n_857;
wire n_898;
wire n_968;
wire n_1067;
wire n_1235;
wire n_1323;
wire n_2584;
wire n_2375;
wire n_1462;
wire n_1937;
wire n_2012;
wire n_1064;
wire n_633;
wire n_900;
wire n_1446;
wire n_1282;
wire n_1701;
wire n_1093;
wire n_1551;
wire n_2039;
wire n_1755;
wire n_1285;
wire n_733;
wire n_761;
wire n_2212;
wire n_731;
wire n_1813;
wire n_2268;
wire n_1452;
wire n_2835;
wire n_1573;
wire n_2734;
wire n_668;
wire n_2569;
wire n_758;
wire n_2252;
wire n_2111;
wire n_2420;
wire n_1996;
wire n_1106;
wire n_2009;
wire n_648;
wire n_784;
wire n_816;
wire n_1322;
wire n_2583;
wire n_1473;
wire n_835;
wire n_1076;
wire n_2024;
wire n_1348;
wire n_2651;
wire n_753;
wire n_2445;
wire n_2733;
wire n_1770;
wire n_1003;
wire n_701;
wire n_2469;
wire n_1125;
wire n_2103;
wire n_2358;
wire n_1710;
wire n_1865;
wire n_2522;
wire n_2641;
wire n_2463;
wire n_1344;
wire n_2355;
wire n_1390;
wire n_2580;
wire n_2699;
wire n_1792;
wire n_2062;
wire n_1141;
wire n_1629;
wire n_1640;
wire n_822;
wire n_1094;
wire n_840;
wire n_1459;
wire n_2153;
wire n_2324;
wire n_1510;
wire n_2710;
wire n_2505;
wire n_2139;
wire n_1099;
wire n_839;
wire n_1754;
wire n_759;
wire n_2397;
wire n_2521;
wire n_1727;
wire n_2740;
wire n_2235;
wire n_1991;
wire n_1575;
wire n_2721;
wire n_1848;
wire n_1892;
wire n_1172;
wire n_2615;
wire n_614;
wire n_2775;
wire n_1212;
wire n_831;
wire n_778;
wire n_1619;
wire n_2351;
wire n_2260;
wire n_1315;
wire n_1660;
wire n_1902;
wire n_997;
wire n_635;
wire n_2206;
wire n_2784;
wire n_2541;
wire n_694;
wire n_1643;
wire n_1320;
wire n_1113;
wire n_2347;
wire n_1152;
wire n_2657;
wire n_2447;
wire n_2034;
wire n_1845;
wire n_2538;
wire n_1934;
wire n_2101;
wire n_2577;
wire n_921;
wire n_2362;
wire n_1615;
wire n_1236;
wire n_2104;
wire n_1265;
wire n_1576;
wire n_2105;
wire n_1470;
wire n_671;
wire n_1533;
wire n_1806;
wire n_2372;
wire n_2552;
wire n_1409;
wire n_1148;
wire n_1588;
wire n_1684;
wire n_1673;
wire n_2422;
wire n_2704;
wire n_1334;
wire n_654;
wire n_2290;
wire n_2856;
wire n_2088;
wire n_1275;
wire n_904;
wire n_2005;
wire n_2048;
wire n_1696;
wire n_1875;
wire n_1059;
wire n_684;
wire n_2429;
wire n_2108;
wire n_2736;
wire n_1039;
wire n_2246;
wire n_1150;
wire n_977;
wire n_2339;
wire n_1628;
wire n_1289;
wire n_1831;
wire n_2532;
wire n_2191;
wire n_1497;
wire n_1866;
wire n_2472;
wire n_2664;
wire n_2705;
wire n_2056;
wire n_2852;
wire n_1136;
wire n_2515;
wire n_1782;
wire n_1190;
wire n_1600;
wire n_1144;
wire n_838;
wire n_1558;
wire n_1941;
wire n_1316;
wire n_2519;
wire n_950;
wire n_1017;
wire n_711;
wire n_734;
wire n_1915;
wire n_2360;
wire n_723;
wire n_1393;
wire n_2240;
wire n_658;
wire n_630;
wire n_1369;
wire n_2846;
wire n_1781;
wire n_709;
wire n_2544;
wire n_809;
wire n_2085;
wire n_2432;
wire n_1686;
wire n_1964;
wire n_881;
wire n_1019;
wire n_1477;
wire n_1777;
wire n_2188;
wire n_1982;
wire n_2097;
wire n_662;
wire n_641;
wire n_2430;
wire n_2504;
wire n_910;
wire n_741;
wire n_939;
wire n_1410;
wire n_2297;
wire n_1114;
wire n_1325;
wire n_1742;
wire n_708;
wire n_1223;
wire n_2545;
wire n_1768;
wire n_2513;
wire n_2193;
wire n_2369;
wire n_1199;
wire n_865;
wire n_1273;
wire n_1983;
wire n_1041;
wire n_2451;
wire n_2115;
wire n_993;
wire n_1862;
wire n_948;
wire n_2017;
wire n_922;
wire n_1004;
wire n_1810;
wire n_2587;
wire n_1347;
wire n_2839;
wire n_860;
wire n_1043;
wire n_1923;
wire n_2670;
wire n_1764;
wire n_2674;
wire n_896;
wire n_1737;
wire n_1479;
wire n_1613;
wire n_2644;
wire n_902;
wire n_1031;
wire n_1723;
wire n_1638;
wire n_853;
wire n_716;
wire n_1571;
wire n_1698;
wire n_1337;
wire n_774;
wire n_1946;
wire n_2148;
wire n_933;
wire n_1779;
wire n_2562;
wire n_954;
wire n_596;
wire n_2051;
wire n_1168;
wire n_1821;
wire n_1310;
wire n_656;
wire n_2673;
wire n_664;
wire n_1591;
wire n_2585;
wire n_1229;
wire n_1683;
wire n_2582;
wire n_2548;
wire n_1896;
wire n_2164;
wire n_1732;
wire n_2381;
wire n_2744;
wire n_1967;
wire n_2384;
wire n_2678;
wire n_2179;
wire n_1280;
wire n_1516;
wire n_1186;
wire n_1705;
wire n_599;
wire n_768;
wire n_1091;
wire n_2052;
wire n_2485;
wire n_1063;
wire n_991;
wire n_2183;
wire n_2205;
wire n_2275;
wire n_2563;
wire n_1724;
wire n_1670;
wire n_1799;
wire n_1707;
wire n_2080;
wire n_2058;
wire n_1126;
wire n_2761;
wire n_2357;
wire n_2029;
wire n_1846;
wire n_1912;
wire n_938;
wire n_1891;
wire n_1328;
wire n_895;
wire n_1639;
wire n_583;
wire n_2209;
wire n_2421;
wire n_1302;
wire n_1000;
wire n_626;
wire n_1581;
wire n_1928;
wire n_946;
wire n_757;
wire n_2047;
wire n_1655;
wire n_1818;
wire n_1146;
wire n_2792;
wire n_1634;
wire n_2596;
wire n_1203;
wire n_998;
wire n_1699;
wire n_1598;
wire n_2269;
wire n_2081;
wire n_937;
wire n_1474;
wire n_2536;
wire n_2524;
wire n_1583;
wire n_1604;
wire n_1631;
wire n_1702;
wire n_1794;
wire n_1375;
wire n_1232;
wire n_996;
wire n_1211;
wire n_1368;
wire n_963;
wire n_1264;
wire n_1082;
wire n_1725;
wire n_2318;
wire n_1827;
wire n_866;
wire n_925;
wire n_1752;
wire n_1313;
wire n_1001;
wire n_1722;
wire n_2361;
wire n_1115;
wire n_2229;
wire n_2819;
wire n_1339;
wire n_1002;
wire n_1644;
wire n_1051;
wire n_2551;
wire n_719;
wire n_1102;
wire n_2255;
wire n_1129;
wire n_1252;
wire n_2239;
wire n_1464;
wire n_1296;
wire n_773;
wire n_2798;
wire n_2316;
wire n_2464;
wire n_1010;
wire n_2830;
wire n_882;
wire n_2706;
wire n_2304;
wire n_1249;
wire n_803;
wire n_1871;
wire n_2514;
wire n_718;
wire n_1434;
wire n_1905;
wire n_1569;
wire n_2573;
wire n_2336;
wire n_1662;
wire n_1299;
wire n_1870;
wire n_2063;
wire n_1925;
wire n_782;
wire n_2654;
wire n_2491;
wire n_1861;
wire n_2079;
wire n_1228;
wire n_2319;
wire n_2152;
wire n_2517;
wire n_1931;
wire n_1244;
wire n_1796;
wire n_2259;
wire n_849;
wire n_2095;
wire n_2719;
wire n_2738;
wire n_1820;
wire n_2590;
wire n_2797;
wire n_1251;
wire n_1989;
wire n_1421;
wire n_2208;
wire n_2423;
wire n_2689;
wire n_2778;
wire n_1762;
wire n_1233;
wire n_1808;
wire n_1574;
wire n_1672;
wire n_2228;
wire n_1635;
wire n_1704;
wire n_893;
wire n_1582;
wire n_841;
wire n_2479;
wire n_886;
wire n_1069;
wire n_1981;
wire n_2824;
wire n_2037;
wire n_1308;
wire n_796;
wire n_2851;
wire n_2823;
wire n_2345;
wire n_1730;
wire n_1374;
wire n_1451;
wire n_2089;
wire n_1487;
wire n_675;

INVx2_ASAP7_75t_L g583 ( 
.A(n_271),
.Y(n_583)
);

CKINVDCx5p33_ASAP7_75t_R g584 ( 
.A(n_412),
.Y(n_584)
);

CKINVDCx5p33_ASAP7_75t_R g585 ( 
.A(n_158),
.Y(n_585)
);

CKINVDCx5p33_ASAP7_75t_R g586 ( 
.A(n_534),
.Y(n_586)
);

CKINVDCx16_ASAP7_75t_R g587 ( 
.A(n_535),
.Y(n_587)
);

CKINVDCx20_ASAP7_75t_R g588 ( 
.A(n_497),
.Y(n_588)
);

CKINVDCx5p33_ASAP7_75t_R g589 ( 
.A(n_562),
.Y(n_589)
);

CKINVDCx5p33_ASAP7_75t_R g590 ( 
.A(n_442),
.Y(n_590)
);

CKINVDCx5p33_ASAP7_75t_R g591 ( 
.A(n_256),
.Y(n_591)
);

INVx1_ASAP7_75t_L g592 ( 
.A(n_134),
.Y(n_592)
);

INVx1_ASAP7_75t_L g593 ( 
.A(n_568),
.Y(n_593)
);

INVx1_ASAP7_75t_L g594 ( 
.A(n_476),
.Y(n_594)
);

CKINVDCx5p33_ASAP7_75t_R g595 ( 
.A(n_11),
.Y(n_595)
);

CKINVDCx5p33_ASAP7_75t_R g596 ( 
.A(n_529),
.Y(n_596)
);

CKINVDCx5p33_ASAP7_75t_R g597 ( 
.A(n_544),
.Y(n_597)
);

INVx1_ASAP7_75t_L g598 ( 
.A(n_309),
.Y(n_598)
);

CKINVDCx5p33_ASAP7_75t_R g599 ( 
.A(n_471),
.Y(n_599)
);

CKINVDCx5p33_ASAP7_75t_R g600 ( 
.A(n_550),
.Y(n_600)
);

CKINVDCx5p33_ASAP7_75t_R g601 ( 
.A(n_18),
.Y(n_601)
);

INVx1_ASAP7_75t_L g602 ( 
.A(n_37),
.Y(n_602)
);

CKINVDCx5p33_ASAP7_75t_R g603 ( 
.A(n_427),
.Y(n_603)
);

INVx1_ASAP7_75t_SL g604 ( 
.A(n_16),
.Y(n_604)
);

BUFx10_ASAP7_75t_L g605 ( 
.A(n_38),
.Y(n_605)
);

CKINVDCx5p33_ASAP7_75t_R g606 ( 
.A(n_563),
.Y(n_606)
);

CKINVDCx20_ASAP7_75t_R g607 ( 
.A(n_551),
.Y(n_607)
);

INVx1_ASAP7_75t_L g608 ( 
.A(n_468),
.Y(n_608)
);

CKINVDCx16_ASAP7_75t_R g609 ( 
.A(n_230),
.Y(n_609)
);

CKINVDCx16_ASAP7_75t_R g610 ( 
.A(n_407),
.Y(n_610)
);

INVx1_ASAP7_75t_L g611 ( 
.A(n_580),
.Y(n_611)
);

BUFx3_ASAP7_75t_L g612 ( 
.A(n_536),
.Y(n_612)
);

CKINVDCx5p33_ASAP7_75t_R g613 ( 
.A(n_564),
.Y(n_613)
);

CKINVDCx5p33_ASAP7_75t_R g614 ( 
.A(n_64),
.Y(n_614)
);

CKINVDCx5p33_ASAP7_75t_R g615 ( 
.A(n_549),
.Y(n_615)
);

CKINVDCx5p33_ASAP7_75t_R g616 ( 
.A(n_421),
.Y(n_616)
);

INVx1_ASAP7_75t_L g617 ( 
.A(n_181),
.Y(n_617)
);

CKINVDCx5p33_ASAP7_75t_R g618 ( 
.A(n_411),
.Y(n_618)
);

CKINVDCx5p33_ASAP7_75t_R g619 ( 
.A(n_391),
.Y(n_619)
);

CKINVDCx5p33_ASAP7_75t_R g620 ( 
.A(n_156),
.Y(n_620)
);

CKINVDCx5p33_ASAP7_75t_R g621 ( 
.A(n_322),
.Y(n_621)
);

INVx1_ASAP7_75t_L g622 ( 
.A(n_203),
.Y(n_622)
);

CKINVDCx5p33_ASAP7_75t_R g623 ( 
.A(n_64),
.Y(n_623)
);

BUFx3_ASAP7_75t_L g624 ( 
.A(n_287),
.Y(n_624)
);

CKINVDCx5p33_ASAP7_75t_R g625 ( 
.A(n_226),
.Y(n_625)
);

CKINVDCx5p33_ASAP7_75t_R g626 ( 
.A(n_298),
.Y(n_626)
);

INVx1_ASAP7_75t_L g627 ( 
.A(n_225),
.Y(n_627)
);

CKINVDCx5p33_ASAP7_75t_R g628 ( 
.A(n_413),
.Y(n_628)
);

CKINVDCx5p33_ASAP7_75t_R g629 ( 
.A(n_388),
.Y(n_629)
);

INVx1_ASAP7_75t_L g630 ( 
.A(n_51),
.Y(n_630)
);

INVx2_ASAP7_75t_L g631 ( 
.A(n_515),
.Y(n_631)
);

CKINVDCx5p33_ASAP7_75t_R g632 ( 
.A(n_34),
.Y(n_632)
);

INVx2_ASAP7_75t_L g633 ( 
.A(n_279),
.Y(n_633)
);

CKINVDCx20_ASAP7_75t_R g634 ( 
.A(n_218),
.Y(n_634)
);

CKINVDCx20_ASAP7_75t_R g635 ( 
.A(n_293),
.Y(n_635)
);

CKINVDCx16_ASAP7_75t_R g636 ( 
.A(n_540),
.Y(n_636)
);

INVx1_ASAP7_75t_L g637 ( 
.A(n_292),
.Y(n_637)
);

INVx1_ASAP7_75t_L g638 ( 
.A(n_334),
.Y(n_638)
);

CKINVDCx5p33_ASAP7_75t_R g639 ( 
.A(n_344),
.Y(n_639)
);

INVx1_ASAP7_75t_L g640 ( 
.A(n_173),
.Y(n_640)
);

INVxp33_ASAP7_75t_R g641 ( 
.A(n_554),
.Y(n_641)
);

CKINVDCx5p33_ASAP7_75t_R g642 ( 
.A(n_578),
.Y(n_642)
);

BUFx10_ASAP7_75t_L g643 ( 
.A(n_325),
.Y(n_643)
);

CKINVDCx5p33_ASAP7_75t_R g644 ( 
.A(n_268),
.Y(n_644)
);

INVx2_ASAP7_75t_L g645 ( 
.A(n_572),
.Y(n_645)
);

CKINVDCx5p33_ASAP7_75t_R g646 ( 
.A(n_265),
.Y(n_646)
);

INVx2_ASAP7_75t_L g647 ( 
.A(n_161),
.Y(n_647)
);

BUFx3_ASAP7_75t_L g648 ( 
.A(n_106),
.Y(n_648)
);

CKINVDCx5p33_ASAP7_75t_R g649 ( 
.A(n_324),
.Y(n_649)
);

BUFx3_ASAP7_75t_L g650 ( 
.A(n_530),
.Y(n_650)
);

CKINVDCx5p33_ASAP7_75t_R g651 ( 
.A(n_288),
.Y(n_651)
);

INVx1_ASAP7_75t_L g652 ( 
.A(n_299),
.Y(n_652)
);

CKINVDCx5p33_ASAP7_75t_R g653 ( 
.A(n_581),
.Y(n_653)
);

HB1xp67_ASAP7_75t_L g654 ( 
.A(n_566),
.Y(n_654)
);

INVx2_ASAP7_75t_L g655 ( 
.A(n_398),
.Y(n_655)
);

INVx1_ASAP7_75t_L g656 ( 
.A(n_503),
.Y(n_656)
);

CKINVDCx5p33_ASAP7_75t_R g657 ( 
.A(n_42),
.Y(n_657)
);

CKINVDCx5p33_ASAP7_75t_R g658 ( 
.A(n_571),
.Y(n_658)
);

CKINVDCx5p33_ASAP7_75t_R g659 ( 
.A(n_515),
.Y(n_659)
);

CKINVDCx5p33_ASAP7_75t_R g660 ( 
.A(n_380),
.Y(n_660)
);

BUFx3_ASAP7_75t_L g661 ( 
.A(n_575),
.Y(n_661)
);

CKINVDCx5p33_ASAP7_75t_R g662 ( 
.A(n_116),
.Y(n_662)
);

INVx1_ASAP7_75t_L g663 ( 
.A(n_310),
.Y(n_663)
);

BUFx3_ASAP7_75t_L g664 ( 
.A(n_79),
.Y(n_664)
);

CKINVDCx5p33_ASAP7_75t_R g665 ( 
.A(n_242),
.Y(n_665)
);

CKINVDCx5p33_ASAP7_75t_R g666 ( 
.A(n_204),
.Y(n_666)
);

INVx1_ASAP7_75t_L g667 ( 
.A(n_445),
.Y(n_667)
);

INVx1_ASAP7_75t_L g668 ( 
.A(n_156),
.Y(n_668)
);

CKINVDCx5p33_ASAP7_75t_R g669 ( 
.A(n_399),
.Y(n_669)
);

INVx1_ASAP7_75t_L g670 ( 
.A(n_175),
.Y(n_670)
);

CKINVDCx20_ASAP7_75t_R g671 ( 
.A(n_152),
.Y(n_671)
);

INVx2_ASAP7_75t_SL g672 ( 
.A(n_270),
.Y(n_672)
);

INVx1_ASAP7_75t_L g673 ( 
.A(n_561),
.Y(n_673)
);

CKINVDCx5p33_ASAP7_75t_R g674 ( 
.A(n_325),
.Y(n_674)
);

CKINVDCx5p33_ASAP7_75t_R g675 ( 
.A(n_526),
.Y(n_675)
);

INVx1_ASAP7_75t_L g676 ( 
.A(n_303),
.Y(n_676)
);

INVx1_ASAP7_75t_L g677 ( 
.A(n_400),
.Y(n_677)
);

INVx1_ASAP7_75t_L g678 ( 
.A(n_546),
.Y(n_678)
);

CKINVDCx5p33_ASAP7_75t_R g679 ( 
.A(n_314),
.Y(n_679)
);

INVx2_ASAP7_75t_SL g680 ( 
.A(n_212),
.Y(n_680)
);

CKINVDCx5p33_ASAP7_75t_R g681 ( 
.A(n_481),
.Y(n_681)
);

CKINVDCx5p33_ASAP7_75t_R g682 ( 
.A(n_112),
.Y(n_682)
);

CKINVDCx5p33_ASAP7_75t_R g683 ( 
.A(n_75),
.Y(n_683)
);

CKINVDCx5p33_ASAP7_75t_R g684 ( 
.A(n_29),
.Y(n_684)
);

CKINVDCx5p33_ASAP7_75t_R g685 ( 
.A(n_302),
.Y(n_685)
);

CKINVDCx5p33_ASAP7_75t_R g686 ( 
.A(n_247),
.Y(n_686)
);

CKINVDCx20_ASAP7_75t_R g687 ( 
.A(n_214),
.Y(n_687)
);

CKINVDCx5p33_ASAP7_75t_R g688 ( 
.A(n_71),
.Y(n_688)
);

CKINVDCx5p33_ASAP7_75t_R g689 ( 
.A(n_88),
.Y(n_689)
);

CKINVDCx5p33_ASAP7_75t_R g690 ( 
.A(n_279),
.Y(n_690)
);

CKINVDCx5p33_ASAP7_75t_R g691 ( 
.A(n_96),
.Y(n_691)
);

BUFx2_ASAP7_75t_L g692 ( 
.A(n_234),
.Y(n_692)
);

CKINVDCx20_ASAP7_75t_R g693 ( 
.A(n_361),
.Y(n_693)
);

CKINVDCx5p33_ASAP7_75t_R g694 ( 
.A(n_455),
.Y(n_694)
);

INVx1_ASAP7_75t_L g695 ( 
.A(n_108),
.Y(n_695)
);

INVx2_ASAP7_75t_L g696 ( 
.A(n_406),
.Y(n_696)
);

CKINVDCx5p33_ASAP7_75t_R g697 ( 
.A(n_201),
.Y(n_697)
);

CKINVDCx5p33_ASAP7_75t_R g698 ( 
.A(n_136),
.Y(n_698)
);

BUFx10_ASAP7_75t_L g699 ( 
.A(n_179),
.Y(n_699)
);

INVx1_ASAP7_75t_SL g700 ( 
.A(n_552),
.Y(n_700)
);

CKINVDCx5p33_ASAP7_75t_R g701 ( 
.A(n_383),
.Y(n_701)
);

BUFx10_ASAP7_75t_L g702 ( 
.A(n_505),
.Y(n_702)
);

INVx2_ASAP7_75t_L g703 ( 
.A(n_470),
.Y(n_703)
);

CKINVDCx5p33_ASAP7_75t_R g704 ( 
.A(n_570),
.Y(n_704)
);

BUFx10_ASAP7_75t_L g705 ( 
.A(n_246),
.Y(n_705)
);

HB1xp67_ASAP7_75t_L g706 ( 
.A(n_187),
.Y(n_706)
);

BUFx6f_ASAP7_75t_L g707 ( 
.A(n_49),
.Y(n_707)
);

CKINVDCx16_ASAP7_75t_R g708 ( 
.A(n_192),
.Y(n_708)
);

CKINVDCx5p33_ASAP7_75t_R g709 ( 
.A(n_560),
.Y(n_709)
);

CKINVDCx5p33_ASAP7_75t_R g710 ( 
.A(n_423),
.Y(n_710)
);

INVx1_ASAP7_75t_L g711 ( 
.A(n_507),
.Y(n_711)
);

INVx1_ASAP7_75t_L g712 ( 
.A(n_35),
.Y(n_712)
);

INVx1_ASAP7_75t_L g713 ( 
.A(n_406),
.Y(n_713)
);

CKINVDCx5p33_ASAP7_75t_R g714 ( 
.A(n_574),
.Y(n_714)
);

BUFx6f_ASAP7_75t_L g715 ( 
.A(n_461),
.Y(n_715)
);

CKINVDCx5p33_ASAP7_75t_R g716 ( 
.A(n_375),
.Y(n_716)
);

BUFx10_ASAP7_75t_L g717 ( 
.A(n_71),
.Y(n_717)
);

CKINVDCx16_ASAP7_75t_R g718 ( 
.A(n_558),
.Y(n_718)
);

BUFx6f_ASAP7_75t_L g719 ( 
.A(n_433),
.Y(n_719)
);

CKINVDCx5p33_ASAP7_75t_R g720 ( 
.A(n_316),
.Y(n_720)
);

INVx1_ASAP7_75t_L g721 ( 
.A(n_196),
.Y(n_721)
);

CKINVDCx5p33_ASAP7_75t_R g722 ( 
.A(n_430),
.Y(n_722)
);

INVx2_ASAP7_75t_L g723 ( 
.A(n_337),
.Y(n_723)
);

INVx1_ASAP7_75t_L g724 ( 
.A(n_576),
.Y(n_724)
);

INVx1_ASAP7_75t_L g725 ( 
.A(n_345),
.Y(n_725)
);

CKINVDCx5p33_ASAP7_75t_R g726 ( 
.A(n_278),
.Y(n_726)
);

CKINVDCx5p33_ASAP7_75t_R g727 ( 
.A(n_418),
.Y(n_727)
);

CKINVDCx5p33_ASAP7_75t_R g728 ( 
.A(n_255),
.Y(n_728)
);

CKINVDCx20_ASAP7_75t_R g729 ( 
.A(n_271),
.Y(n_729)
);

CKINVDCx5p33_ASAP7_75t_R g730 ( 
.A(n_467),
.Y(n_730)
);

CKINVDCx5p33_ASAP7_75t_R g731 ( 
.A(n_385),
.Y(n_731)
);

HB1xp67_ASAP7_75t_L g732 ( 
.A(n_278),
.Y(n_732)
);

INVx1_ASAP7_75t_L g733 ( 
.A(n_153),
.Y(n_733)
);

BUFx10_ASAP7_75t_L g734 ( 
.A(n_169),
.Y(n_734)
);

INVx1_ASAP7_75t_L g735 ( 
.A(n_14),
.Y(n_735)
);

INVx1_ASAP7_75t_L g736 ( 
.A(n_84),
.Y(n_736)
);

INVx1_ASAP7_75t_L g737 ( 
.A(n_465),
.Y(n_737)
);

CKINVDCx5p33_ASAP7_75t_R g738 ( 
.A(n_555),
.Y(n_738)
);

INVx1_ASAP7_75t_L g739 ( 
.A(n_527),
.Y(n_739)
);

CKINVDCx16_ASAP7_75t_R g740 ( 
.A(n_470),
.Y(n_740)
);

CKINVDCx5p33_ASAP7_75t_R g741 ( 
.A(n_52),
.Y(n_741)
);

INVx1_ASAP7_75t_L g742 ( 
.A(n_158),
.Y(n_742)
);

CKINVDCx5p33_ASAP7_75t_R g743 ( 
.A(n_567),
.Y(n_743)
);

CKINVDCx5p33_ASAP7_75t_R g744 ( 
.A(n_547),
.Y(n_744)
);

CKINVDCx5p33_ASAP7_75t_R g745 ( 
.A(n_525),
.Y(n_745)
);

CKINVDCx5p33_ASAP7_75t_R g746 ( 
.A(n_302),
.Y(n_746)
);

CKINVDCx5p33_ASAP7_75t_R g747 ( 
.A(n_582),
.Y(n_747)
);

CKINVDCx5p33_ASAP7_75t_R g748 ( 
.A(n_215),
.Y(n_748)
);

CKINVDCx5p33_ASAP7_75t_R g749 ( 
.A(n_378),
.Y(n_749)
);

BUFx6f_ASAP7_75t_L g750 ( 
.A(n_553),
.Y(n_750)
);

INVx2_ASAP7_75t_SL g751 ( 
.A(n_84),
.Y(n_751)
);

CKINVDCx5p33_ASAP7_75t_R g752 ( 
.A(n_579),
.Y(n_752)
);

CKINVDCx5p33_ASAP7_75t_R g753 ( 
.A(n_20),
.Y(n_753)
);

INVx2_ASAP7_75t_L g754 ( 
.A(n_94),
.Y(n_754)
);

BUFx6f_ASAP7_75t_L g755 ( 
.A(n_426),
.Y(n_755)
);

BUFx2_ASAP7_75t_L g756 ( 
.A(n_288),
.Y(n_756)
);

INVx1_ASAP7_75t_L g757 ( 
.A(n_4),
.Y(n_757)
);

INVx1_ASAP7_75t_L g758 ( 
.A(n_429),
.Y(n_758)
);

CKINVDCx5p33_ASAP7_75t_R g759 ( 
.A(n_403),
.Y(n_759)
);

CKINVDCx16_ASAP7_75t_R g760 ( 
.A(n_373),
.Y(n_760)
);

CKINVDCx5p33_ASAP7_75t_R g761 ( 
.A(n_382),
.Y(n_761)
);

INVx1_ASAP7_75t_L g762 ( 
.A(n_498),
.Y(n_762)
);

INVx1_ASAP7_75t_L g763 ( 
.A(n_15),
.Y(n_763)
);

CKINVDCx5p33_ASAP7_75t_R g764 ( 
.A(n_484),
.Y(n_764)
);

CKINVDCx5p33_ASAP7_75t_R g765 ( 
.A(n_205),
.Y(n_765)
);

CKINVDCx5p33_ASAP7_75t_R g766 ( 
.A(n_569),
.Y(n_766)
);

CKINVDCx5p33_ASAP7_75t_R g767 ( 
.A(n_161),
.Y(n_767)
);

CKINVDCx5p33_ASAP7_75t_R g768 ( 
.A(n_514),
.Y(n_768)
);

INVx1_ASAP7_75t_SL g769 ( 
.A(n_565),
.Y(n_769)
);

CKINVDCx5p33_ASAP7_75t_R g770 ( 
.A(n_77),
.Y(n_770)
);

CKINVDCx5p33_ASAP7_75t_R g771 ( 
.A(n_12),
.Y(n_771)
);

CKINVDCx5p33_ASAP7_75t_R g772 ( 
.A(n_371),
.Y(n_772)
);

INVx1_ASAP7_75t_L g773 ( 
.A(n_277),
.Y(n_773)
);

INVx1_ASAP7_75t_SL g774 ( 
.A(n_137),
.Y(n_774)
);

INVx2_ASAP7_75t_L g775 ( 
.A(n_227),
.Y(n_775)
);

INVx1_ASAP7_75t_L g776 ( 
.A(n_107),
.Y(n_776)
);

CKINVDCx5p33_ASAP7_75t_R g777 ( 
.A(n_214),
.Y(n_777)
);

CKINVDCx5p33_ASAP7_75t_R g778 ( 
.A(n_413),
.Y(n_778)
);

CKINVDCx5p33_ASAP7_75t_R g779 ( 
.A(n_291),
.Y(n_779)
);

INVx2_ASAP7_75t_L g780 ( 
.A(n_127),
.Y(n_780)
);

CKINVDCx5p33_ASAP7_75t_R g781 ( 
.A(n_459),
.Y(n_781)
);

CKINVDCx5p33_ASAP7_75t_R g782 ( 
.A(n_354),
.Y(n_782)
);

BUFx8_ASAP7_75t_SL g783 ( 
.A(n_258),
.Y(n_783)
);

CKINVDCx5p33_ASAP7_75t_R g784 ( 
.A(n_245),
.Y(n_784)
);

INVx2_ASAP7_75t_L g785 ( 
.A(n_421),
.Y(n_785)
);

CKINVDCx5p33_ASAP7_75t_R g786 ( 
.A(n_134),
.Y(n_786)
);

CKINVDCx20_ASAP7_75t_R g787 ( 
.A(n_236),
.Y(n_787)
);

INVx1_ASAP7_75t_L g788 ( 
.A(n_25),
.Y(n_788)
);

CKINVDCx5p33_ASAP7_75t_R g789 ( 
.A(n_317),
.Y(n_789)
);

INVx1_ASAP7_75t_L g790 ( 
.A(n_433),
.Y(n_790)
);

CKINVDCx5p33_ASAP7_75t_R g791 ( 
.A(n_273),
.Y(n_791)
);

CKINVDCx5p33_ASAP7_75t_R g792 ( 
.A(n_14),
.Y(n_792)
);

BUFx10_ASAP7_75t_L g793 ( 
.A(n_285),
.Y(n_793)
);

CKINVDCx5p33_ASAP7_75t_R g794 ( 
.A(n_556),
.Y(n_794)
);

INVx1_ASAP7_75t_SL g795 ( 
.A(n_318),
.Y(n_795)
);

CKINVDCx5p33_ASAP7_75t_R g796 ( 
.A(n_420),
.Y(n_796)
);

INVx1_ASAP7_75t_SL g797 ( 
.A(n_62),
.Y(n_797)
);

INVx2_ASAP7_75t_SL g798 ( 
.A(n_273),
.Y(n_798)
);

INVxp67_ASAP7_75t_L g799 ( 
.A(n_457),
.Y(n_799)
);

CKINVDCx5p33_ASAP7_75t_R g800 ( 
.A(n_573),
.Y(n_800)
);

INVx1_ASAP7_75t_L g801 ( 
.A(n_290),
.Y(n_801)
);

INVx1_ASAP7_75t_L g802 ( 
.A(n_100),
.Y(n_802)
);

INVx1_ASAP7_75t_L g803 ( 
.A(n_454),
.Y(n_803)
);

CKINVDCx5p33_ASAP7_75t_R g804 ( 
.A(n_497),
.Y(n_804)
);

CKINVDCx5p33_ASAP7_75t_R g805 ( 
.A(n_289),
.Y(n_805)
);

CKINVDCx20_ASAP7_75t_R g806 ( 
.A(n_85),
.Y(n_806)
);

INVx1_ASAP7_75t_L g807 ( 
.A(n_414),
.Y(n_807)
);

INVx2_ASAP7_75t_SL g808 ( 
.A(n_383),
.Y(n_808)
);

CKINVDCx5p33_ASAP7_75t_R g809 ( 
.A(n_88),
.Y(n_809)
);

CKINVDCx5p33_ASAP7_75t_R g810 ( 
.A(n_364),
.Y(n_810)
);

CKINVDCx5p33_ASAP7_75t_R g811 ( 
.A(n_559),
.Y(n_811)
);

INVx2_ASAP7_75t_L g812 ( 
.A(n_136),
.Y(n_812)
);

INVxp67_ASAP7_75t_L g813 ( 
.A(n_262),
.Y(n_813)
);

INVx1_ASAP7_75t_L g814 ( 
.A(n_541),
.Y(n_814)
);

INVx1_ASAP7_75t_L g815 ( 
.A(n_40),
.Y(n_815)
);

BUFx6f_ASAP7_75t_L g816 ( 
.A(n_368),
.Y(n_816)
);

INVx1_ASAP7_75t_L g817 ( 
.A(n_237),
.Y(n_817)
);

BUFx10_ASAP7_75t_L g818 ( 
.A(n_54),
.Y(n_818)
);

BUFx6f_ASAP7_75t_L g819 ( 
.A(n_520),
.Y(n_819)
);

CKINVDCx5p33_ASAP7_75t_R g820 ( 
.A(n_557),
.Y(n_820)
);

CKINVDCx5p33_ASAP7_75t_R g821 ( 
.A(n_67),
.Y(n_821)
);

CKINVDCx14_ASAP7_75t_R g822 ( 
.A(n_450),
.Y(n_822)
);

INVx1_ASAP7_75t_L g823 ( 
.A(n_60),
.Y(n_823)
);

CKINVDCx5p33_ASAP7_75t_R g824 ( 
.A(n_449),
.Y(n_824)
);

CKINVDCx5p33_ASAP7_75t_R g825 ( 
.A(n_217),
.Y(n_825)
);

INVx1_ASAP7_75t_L g826 ( 
.A(n_548),
.Y(n_826)
);

CKINVDCx5p33_ASAP7_75t_R g827 ( 
.A(n_86),
.Y(n_827)
);

CKINVDCx5p33_ASAP7_75t_R g828 ( 
.A(n_255),
.Y(n_828)
);

INVx1_ASAP7_75t_SL g829 ( 
.A(n_512),
.Y(n_829)
);

CKINVDCx20_ASAP7_75t_R g830 ( 
.A(n_297),
.Y(n_830)
);

CKINVDCx5p33_ASAP7_75t_R g831 ( 
.A(n_114),
.Y(n_831)
);

CKINVDCx5p33_ASAP7_75t_R g832 ( 
.A(n_283),
.Y(n_832)
);

CKINVDCx5p33_ASAP7_75t_R g833 ( 
.A(n_524),
.Y(n_833)
);

INVx1_ASAP7_75t_L g834 ( 
.A(n_624),
.Y(n_834)
);

INVx2_ASAP7_75t_L g835 ( 
.A(n_707),
.Y(n_835)
);

INVxp33_ASAP7_75t_SL g836 ( 
.A(n_706),
.Y(n_836)
);

INVx1_ASAP7_75t_SL g837 ( 
.A(n_783),
.Y(n_837)
);

CKINVDCx5p33_ASAP7_75t_R g838 ( 
.A(n_822),
.Y(n_838)
);

INVx1_ASAP7_75t_L g839 ( 
.A(n_624),
.Y(n_839)
);

INVx1_ASAP7_75t_L g840 ( 
.A(n_648),
.Y(n_840)
);

INVxp67_ASAP7_75t_L g841 ( 
.A(n_692),
.Y(n_841)
);

INVx1_ASAP7_75t_L g842 ( 
.A(n_648),
.Y(n_842)
);

BUFx6f_ASAP7_75t_L g843 ( 
.A(n_750),
.Y(n_843)
);

BUFx3_ASAP7_75t_L g844 ( 
.A(n_612),
.Y(n_844)
);

INVx1_ASAP7_75t_L g845 ( 
.A(n_664),
.Y(n_845)
);

INVxp33_ASAP7_75t_SL g846 ( 
.A(n_732),
.Y(n_846)
);

CKINVDCx16_ASAP7_75t_R g847 ( 
.A(n_609),
.Y(n_847)
);

INVx1_ASAP7_75t_L g848 ( 
.A(n_664),
.Y(n_848)
);

INVxp67_ASAP7_75t_SL g849 ( 
.A(n_707),
.Y(n_849)
);

CKINVDCx20_ASAP7_75t_R g850 ( 
.A(n_588),
.Y(n_850)
);

INVxp33_ASAP7_75t_L g851 ( 
.A(n_783),
.Y(n_851)
);

INVx1_ASAP7_75t_L g852 ( 
.A(n_592),
.Y(n_852)
);

INVx1_ASAP7_75t_L g853 ( 
.A(n_594),
.Y(n_853)
);

INVx1_ASAP7_75t_L g854 ( 
.A(n_598),
.Y(n_854)
);

INVx1_ASAP7_75t_L g855 ( 
.A(n_602),
.Y(n_855)
);

CKINVDCx5p33_ASAP7_75t_R g856 ( 
.A(n_587),
.Y(n_856)
);

CKINVDCx5p33_ASAP7_75t_R g857 ( 
.A(n_636),
.Y(n_857)
);

CKINVDCx5p33_ASAP7_75t_R g858 ( 
.A(n_610),
.Y(n_858)
);

INVx1_ASAP7_75t_L g859 ( 
.A(n_608),
.Y(n_859)
);

INVxp67_ASAP7_75t_SL g860 ( 
.A(n_707),
.Y(n_860)
);

INVx1_ASAP7_75t_L g861 ( 
.A(n_617),
.Y(n_861)
);

CKINVDCx5p33_ASAP7_75t_R g862 ( 
.A(n_718),
.Y(n_862)
);

INVx1_ASAP7_75t_L g863 ( 
.A(n_622),
.Y(n_863)
);

INVx1_ASAP7_75t_L g864 ( 
.A(n_627),
.Y(n_864)
);

INVx1_ASAP7_75t_L g865 ( 
.A(n_630),
.Y(n_865)
);

INVx1_ASAP7_75t_L g866 ( 
.A(n_637),
.Y(n_866)
);

INVx1_ASAP7_75t_L g867 ( 
.A(n_638),
.Y(n_867)
);

CKINVDCx16_ASAP7_75t_R g868 ( 
.A(n_708),
.Y(n_868)
);

INVx1_ASAP7_75t_L g869 ( 
.A(n_640),
.Y(n_869)
);

INVxp33_ASAP7_75t_SL g870 ( 
.A(n_654),
.Y(n_870)
);

INVx1_ASAP7_75t_L g871 ( 
.A(n_652),
.Y(n_871)
);

INVx1_ASAP7_75t_L g872 ( 
.A(n_656),
.Y(n_872)
);

INVx1_ASAP7_75t_L g873 ( 
.A(n_663),
.Y(n_873)
);

INVx2_ASAP7_75t_L g874 ( 
.A(n_707),
.Y(n_874)
);

INVx1_ASAP7_75t_L g875 ( 
.A(n_667),
.Y(n_875)
);

INVx1_ASAP7_75t_L g876 ( 
.A(n_668),
.Y(n_876)
);

INVx1_ASAP7_75t_L g877 ( 
.A(n_670),
.Y(n_877)
);

INVx1_ASAP7_75t_SL g878 ( 
.A(n_588),
.Y(n_878)
);

BUFx3_ASAP7_75t_L g879 ( 
.A(n_612),
.Y(n_879)
);

CKINVDCx20_ASAP7_75t_R g880 ( 
.A(n_634),
.Y(n_880)
);

INVx1_ASAP7_75t_L g881 ( 
.A(n_676),
.Y(n_881)
);

CKINVDCx16_ASAP7_75t_R g882 ( 
.A(n_740),
.Y(n_882)
);

CKINVDCx20_ASAP7_75t_R g883 ( 
.A(n_634),
.Y(n_883)
);

CKINVDCx5p33_ASAP7_75t_R g884 ( 
.A(n_607),
.Y(n_884)
);

INVx1_ASAP7_75t_L g885 ( 
.A(n_677),
.Y(n_885)
);

INVx1_ASAP7_75t_L g886 ( 
.A(n_695),
.Y(n_886)
);

BUFx6f_ASAP7_75t_L g887 ( 
.A(n_750),
.Y(n_887)
);

INVx1_ASAP7_75t_L g888 ( 
.A(n_711),
.Y(n_888)
);

INVx1_ASAP7_75t_L g889 ( 
.A(n_712),
.Y(n_889)
);

INVxp33_ASAP7_75t_SL g890 ( 
.A(n_599),
.Y(n_890)
);

CKINVDCx5p33_ASAP7_75t_R g891 ( 
.A(n_607),
.Y(n_891)
);

INVx2_ASAP7_75t_SL g892 ( 
.A(n_605),
.Y(n_892)
);

INVx1_ASAP7_75t_L g893 ( 
.A(n_713),
.Y(n_893)
);

INVx1_ASAP7_75t_L g894 ( 
.A(n_721),
.Y(n_894)
);

INVx1_ASAP7_75t_L g895 ( 
.A(n_725),
.Y(n_895)
);

INVxp33_ASAP7_75t_SL g896 ( 
.A(n_599),
.Y(n_896)
);

INVx1_ASAP7_75t_L g897 ( 
.A(n_733),
.Y(n_897)
);

INVx1_ASAP7_75t_L g898 ( 
.A(n_735),
.Y(n_898)
);

INVxp33_ASAP7_75t_L g899 ( 
.A(n_756),
.Y(n_899)
);

INVx1_ASAP7_75t_L g900 ( 
.A(n_736),
.Y(n_900)
);

CKINVDCx5p33_ASAP7_75t_R g901 ( 
.A(n_600),
.Y(n_901)
);

INVx1_ASAP7_75t_L g902 ( 
.A(n_737),
.Y(n_902)
);

INVx1_ASAP7_75t_L g903 ( 
.A(n_739),
.Y(n_903)
);

BUFx6f_ASAP7_75t_L g904 ( 
.A(n_750),
.Y(n_904)
);

INVx1_ASAP7_75t_L g905 ( 
.A(n_742),
.Y(n_905)
);

INVx1_ASAP7_75t_L g906 ( 
.A(n_757),
.Y(n_906)
);

INVx1_ASAP7_75t_L g907 ( 
.A(n_758),
.Y(n_907)
);

INVx1_ASAP7_75t_L g908 ( 
.A(n_762),
.Y(n_908)
);

INVxp67_ASAP7_75t_SL g909 ( 
.A(n_715),
.Y(n_909)
);

CKINVDCx5p33_ASAP7_75t_R g910 ( 
.A(n_600),
.Y(n_910)
);

INVx1_ASAP7_75t_L g911 ( 
.A(n_763),
.Y(n_911)
);

INVx4_ASAP7_75t_R g912 ( 
.A(n_641),
.Y(n_912)
);

CKINVDCx5p33_ASAP7_75t_R g913 ( 
.A(n_606),
.Y(n_913)
);

CKINVDCx16_ASAP7_75t_R g914 ( 
.A(n_760),
.Y(n_914)
);

HB1xp67_ASAP7_75t_L g915 ( 
.A(n_601),
.Y(n_915)
);

INVx1_ASAP7_75t_L g916 ( 
.A(n_773),
.Y(n_916)
);

CKINVDCx16_ASAP7_75t_R g917 ( 
.A(n_605),
.Y(n_917)
);

CKINVDCx5p33_ASAP7_75t_R g918 ( 
.A(n_606),
.Y(n_918)
);

HB1xp67_ASAP7_75t_L g919 ( 
.A(n_601),
.Y(n_919)
);

INVx1_ASAP7_75t_L g920 ( 
.A(n_776),
.Y(n_920)
);

INVx1_ASAP7_75t_L g921 ( 
.A(n_788),
.Y(n_921)
);

INVx1_ASAP7_75t_L g922 ( 
.A(n_790),
.Y(n_922)
);

INVx1_ASAP7_75t_L g923 ( 
.A(n_801),
.Y(n_923)
);

INVx1_ASAP7_75t_L g924 ( 
.A(n_802),
.Y(n_924)
);

INVx1_ASAP7_75t_L g925 ( 
.A(n_803),
.Y(n_925)
);

CKINVDCx5p33_ASAP7_75t_R g926 ( 
.A(n_584),
.Y(n_926)
);

INVx1_ASAP7_75t_L g927 ( 
.A(n_807),
.Y(n_927)
);

INVx1_ASAP7_75t_L g928 ( 
.A(n_815),
.Y(n_928)
);

BUFx2_ASAP7_75t_L g929 ( 
.A(n_833),
.Y(n_929)
);

NAND2xp5_ASAP7_75t_L g930 ( 
.A(n_593),
.B(n_0),
.Y(n_930)
);

INVx1_ASAP7_75t_L g931 ( 
.A(n_817),
.Y(n_931)
);

INVx1_ASAP7_75t_L g932 ( 
.A(n_823),
.Y(n_932)
);

CKINVDCx5p33_ASAP7_75t_R g933 ( 
.A(n_585),
.Y(n_933)
);

INVx1_ASAP7_75t_L g934 ( 
.A(n_583),
.Y(n_934)
);

CKINVDCx14_ASAP7_75t_R g935 ( 
.A(n_586),
.Y(n_935)
);

INVx1_ASAP7_75t_L g936 ( 
.A(n_583),
.Y(n_936)
);

INVxp67_ASAP7_75t_L g937 ( 
.A(n_672),
.Y(n_937)
);

BUFx12f_ASAP7_75t_L g938 ( 
.A(n_838),
.Y(n_938)
);

INVx2_ASAP7_75t_L g939 ( 
.A(n_843),
.Y(n_939)
);

INVx1_ASAP7_75t_L g940 ( 
.A(n_835),
.Y(n_940)
);

INVx4_ASAP7_75t_L g941 ( 
.A(n_843),
.Y(n_941)
);

OAI22x1_ASAP7_75t_SL g942 ( 
.A1(n_850),
.A2(n_729),
.B1(n_635),
.B2(n_687),
.Y(n_942)
);

BUFx12f_ASAP7_75t_L g943 ( 
.A(n_838),
.Y(n_943)
);

NOR2xp33_ASAP7_75t_SL g944 ( 
.A(n_856),
.B(n_729),
.Y(n_944)
);

CKINVDCx6p67_ASAP7_75t_R g945 ( 
.A(n_847),
.Y(n_945)
);

NAND2xp5_ASAP7_75t_L g946 ( 
.A(n_935),
.B(n_611),
.Y(n_946)
);

INVx2_ASAP7_75t_L g947 ( 
.A(n_843),
.Y(n_947)
);

BUFx8_ASAP7_75t_SL g948 ( 
.A(n_850),
.Y(n_948)
);

INVx1_ASAP7_75t_L g949 ( 
.A(n_835),
.Y(n_949)
);

INVxp33_ASAP7_75t_SL g950 ( 
.A(n_856),
.Y(n_950)
);

BUFx6f_ASAP7_75t_L g951 ( 
.A(n_843),
.Y(n_951)
);

BUFx6f_ASAP7_75t_L g952 ( 
.A(n_887),
.Y(n_952)
);

INVx1_ASAP7_75t_L g953 ( 
.A(n_874),
.Y(n_953)
);

INVx2_ASAP7_75t_L g954 ( 
.A(n_887),
.Y(n_954)
);

INVx1_ASAP7_75t_L g955 ( 
.A(n_874),
.Y(n_955)
);

AND2x4_ASAP7_75t_L g956 ( 
.A(n_844),
.B(n_672),
.Y(n_956)
);

INVx1_ASAP7_75t_L g957 ( 
.A(n_849),
.Y(n_957)
);

BUFx6f_ASAP7_75t_L g958 ( 
.A(n_887),
.Y(n_958)
);

BUFx6f_ASAP7_75t_L g959 ( 
.A(n_887),
.Y(n_959)
);

BUFx6f_ASAP7_75t_L g960 ( 
.A(n_904),
.Y(n_960)
);

CKINVDCx5p33_ASAP7_75t_R g961 ( 
.A(n_884),
.Y(n_961)
);

BUFx6f_ASAP7_75t_L g962 ( 
.A(n_904),
.Y(n_962)
);

NAND2xp5_ASAP7_75t_L g963 ( 
.A(n_935),
.B(n_673),
.Y(n_963)
);

BUFx8_ASAP7_75t_SL g964 ( 
.A(n_880),
.Y(n_964)
);

OAI22xp5_ASAP7_75t_L g965 ( 
.A1(n_870),
.A2(n_671),
.B1(n_687),
.B2(n_635),
.Y(n_965)
);

BUFx6f_ASAP7_75t_L g966 ( 
.A(n_904),
.Y(n_966)
);

INVx1_ASAP7_75t_L g967 ( 
.A(n_860),
.Y(n_967)
);

AND2x4_ASAP7_75t_L g968 ( 
.A(n_844),
.B(n_680),
.Y(n_968)
);

BUFx6f_ASAP7_75t_L g969 ( 
.A(n_904),
.Y(n_969)
);

INVx1_ASAP7_75t_L g970 ( 
.A(n_909),
.Y(n_970)
);

NAND2xp5_ASAP7_75t_L g971 ( 
.A(n_879),
.B(n_678),
.Y(n_971)
);

INVx5_ASAP7_75t_L g972 ( 
.A(n_879),
.Y(n_972)
);

BUFx12f_ASAP7_75t_L g973 ( 
.A(n_857),
.Y(n_973)
);

INVx1_ASAP7_75t_L g974 ( 
.A(n_934),
.Y(n_974)
);

BUFx3_ASAP7_75t_L g975 ( 
.A(n_834),
.Y(n_975)
);

BUFx6f_ASAP7_75t_L g976 ( 
.A(n_930),
.Y(n_976)
);

HB1xp67_ASAP7_75t_L g977 ( 
.A(n_858),
.Y(n_977)
);

NOR2x1_ASAP7_75t_L g978 ( 
.A(n_839),
.B(n_650),
.Y(n_978)
);

BUFx3_ASAP7_75t_L g979 ( 
.A(n_840),
.Y(n_979)
);

BUFx8_ASAP7_75t_SL g980 ( 
.A(n_880),
.Y(n_980)
);

OA21x2_ASAP7_75t_L g981 ( 
.A1(n_936),
.A2(n_814),
.B(n_724),
.Y(n_981)
);

OAI21x1_ASAP7_75t_L g982 ( 
.A1(n_842),
.A2(n_826),
.B(n_645),
.Y(n_982)
);

CKINVDCx20_ASAP7_75t_R g983 ( 
.A(n_883),
.Y(n_983)
);

BUFx6f_ASAP7_75t_L g984 ( 
.A(n_852),
.Y(n_984)
);

OAI22xp5_ASAP7_75t_SL g985 ( 
.A1(n_883),
.A2(n_671),
.B1(n_787),
.B2(n_693),
.Y(n_985)
);

BUFx6f_ASAP7_75t_L g986 ( 
.A(n_853),
.Y(n_986)
);

INVx1_ASAP7_75t_L g987 ( 
.A(n_854),
.Y(n_987)
);

INVx3_ASAP7_75t_L g988 ( 
.A(n_855),
.Y(n_988)
);

BUFx12f_ASAP7_75t_L g989 ( 
.A(n_857),
.Y(n_989)
);

BUFx12f_ASAP7_75t_L g990 ( 
.A(n_862),
.Y(n_990)
);

BUFx3_ASAP7_75t_L g991 ( 
.A(n_845),
.Y(n_991)
);

INVx2_ASAP7_75t_L g992 ( 
.A(n_859),
.Y(n_992)
);

INVx1_ASAP7_75t_L g993 ( 
.A(n_861),
.Y(n_993)
);

INVx4_ASAP7_75t_L g994 ( 
.A(n_901),
.Y(n_994)
);

INVx1_ASAP7_75t_SL g995 ( 
.A(n_878),
.Y(n_995)
);

INVx1_ASAP7_75t_L g996 ( 
.A(n_863),
.Y(n_996)
);

INVx2_ASAP7_75t_L g997 ( 
.A(n_864),
.Y(n_997)
);

BUFx8_ASAP7_75t_SL g998 ( 
.A(n_884),
.Y(n_998)
);

OAI21x1_ASAP7_75t_L g999 ( 
.A1(n_848),
.A2(n_645),
.B(n_633),
.Y(n_999)
);

INVx1_ASAP7_75t_L g1000 ( 
.A(n_865),
.Y(n_1000)
);

BUFx6f_ASAP7_75t_L g1001 ( 
.A(n_866),
.Y(n_1001)
);

NAND2xp5_ASAP7_75t_L g1002 ( 
.A(n_901),
.B(n_650),
.Y(n_1002)
);

INVx2_ASAP7_75t_L g1003 ( 
.A(n_867),
.Y(n_1003)
);

BUFx2_ASAP7_75t_L g1004 ( 
.A(n_929),
.Y(n_1004)
);

BUFx6f_ASAP7_75t_L g1005 ( 
.A(n_984),
.Y(n_1005)
);

INVx1_ASAP7_75t_L g1006 ( 
.A(n_999),
.Y(n_1006)
);

INVx2_ASAP7_75t_L g1007 ( 
.A(n_940),
.Y(n_1007)
);

BUFx3_ASAP7_75t_L g1008 ( 
.A(n_957),
.Y(n_1008)
);

INVx2_ASAP7_75t_L g1009 ( 
.A(n_940),
.Y(n_1009)
);

AND2x4_ASAP7_75t_L g1010 ( 
.A(n_956),
.B(n_892),
.Y(n_1010)
);

HB1xp67_ASAP7_75t_L g1011 ( 
.A(n_995),
.Y(n_1011)
);

AND2x4_ASAP7_75t_L g1012 ( 
.A(n_956),
.B(n_892),
.Y(n_1012)
);

AND2x2_ASAP7_75t_L g1013 ( 
.A(n_988),
.B(n_899),
.Y(n_1013)
);

INVx1_ASAP7_75t_L g1014 ( 
.A(n_999),
.Y(n_1014)
);

BUFx6f_ASAP7_75t_L g1015 ( 
.A(n_984),
.Y(n_1015)
);

INVx2_ASAP7_75t_L g1016 ( 
.A(n_949),
.Y(n_1016)
);

INVx1_ASAP7_75t_L g1017 ( 
.A(n_992),
.Y(n_1017)
);

OR2x2_ASAP7_75t_L g1018 ( 
.A(n_1004),
.B(n_868),
.Y(n_1018)
);

AND2x2_ASAP7_75t_L g1019 ( 
.A(n_988),
.B(n_899),
.Y(n_1019)
);

INVx1_ASAP7_75t_L g1020 ( 
.A(n_982),
.Y(n_1020)
);

NAND2xp5_ASAP7_75t_L g1021 ( 
.A(n_976),
.B(n_957),
.Y(n_1021)
);

BUFx8_ASAP7_75t_L g1022 ( 
.A(n_938),
.Y(n_1022)
);

NAND2xp5_ASAP7_75t_SL g1023 ( 
.A(n_994),
.B(n_910),
.Y(n_1023)
);

INVx3_ASAP7_75t_L g1024 ( 
.A(n_941),
.Y(n_1024)
);

INVx2_ASAP7_75t_L g1025 ( 
.A(n_949),
.Y(n_1025)
);

INVx1_ASAP7_75t_L g1026 ( 
.A(n_982),
.Y(n_1026)
);

INVx2_ASAP7_75t_L g1027 ( 
.A(n_953),
.Y(n_1027)
);

NOR2xp33_ASAP7_75t_L g1028 ( 
.A(n_1002),
.B(n_862),
.Y(n_1028)
);

NAND2xp5_ASAP7_75t_L g1029 ( 
.A(n_976),
.B(n_910),
.Y(n_1029)
);

NAND2xp5_ASAP7_75t_L g1030 ( 
.A(n_976),
.B(n_913),
.Y(n_1030)
);

NAND2xp5_ASAP7_75t_L g1031 ( 
.A(n_976),
.B(n_913),
.Y(n_1031)
);

INVx4_ASAP7_75t_L g1032 ( 
.A(n_972),
.Y(n_1032)
);

HB1xp67_ASAP7_75t_L g1033 ( 
.A(n_1004),
.Y(n_1033)
);

BUFx6f_ASAP7_75t_L g1034 ( 
.A(n_984),
.Y(n_1034)
);

OAI21x1_ASAP7_75t_L g1035 ( 
.A1(n_981),
.A2(n_871),
.B(n_869),
.Y(n_1035)
);

INVx2_ASAP7_75t_L g1036 ( 
.A(n_953),
.Y(n_1036)
);

NAND2xp5_ASAP7_75t_L g1037 ( 
.A(n_976),
.B(n_918),
.Y(n_1037)
);

CKINVDCx8_ASAP7_75t_R g1038 ( 
.A(n_961),
.Y(n_1038)
);

INVx1_ASAP7_75t_L g1039 ( 
.A(n_955),
.Y(n_1039)
);

INVx2_ASAP7_75t_L g1040 ( 
.A(n_955),
.Y(n_1040)
);

AND2x4_ASAP7_75t_L g1041 ( 
.A(n_956),
.B(n_872),
.Y(n_1041)
);

AND2x2_ASAP7_75t_L g1042 ( 
.A(n_988),
.B(n_917),
.Y(n_1042)
);

INVx2_ASAP7_75t_L g1043 ( 
.A(n_939),
.Y(n_1043)
);

INVx1_ASAP7_75t_L g1044 ( 
.A(n_981),
.Y(n_1044)
);

INVx1_ASAP7_75t_L g1045 ( 
.A(n_992),
.Y(n_1045)
);

NAND2xp5_ASAP7_75t_L g1046 ( 
.A(n_967),
.B(n_918),
.Y(n_1046)
);

NOR2xp33_ASAP7_75t_L g1047 ( 
.A(n_946),
.B(n_870),
.Y(n_1047)
);

INVx2_ASAP7_75t_L g1048 ( 
.A(n_939),
.Y(n_1048)
);

OAI22xp5_ASAP7_75t_SL g1049 ( 
.A1(n_985),
.A2(n_693),
.B1(n_806),
.B2(n_787),
.Y(n_1049)
);

AND2x2_ASAP7_75t_L g1050 ( 
.A(n_997),
.B(n_937),
.Y(n_1050)
);

INVx1_ASAP7_75t_L g1051 ( 
.A(n_997),
.Y(n_1051)
);

AND2x4_ASAP7_75t_L g1052 ( 
.A(n_956),
.B(n_873),
.Y(n_1052)
);

INVx3_ASAP7_75t_L g1053 ( 
.A(n_941),
.Y(n_1053)
);

OA21x2_ASAP7_75t_L g1054 ( 
.A1(n_947),
.A2(n_876),
.B(n_875),
.Y(n_1054)
);

INVx1_ASAP7_75t_L g1055 ( 
.A(n_981),
.Y(n_1055)
);

INVx1_ASAP7_75t_L g1056 ( 
.A(n_981),
.Y(n_1056)
);

INVx1_ASAP7_75t_L g1057 ( 
.A(n_984),
.Y(n_1057)
);

BUFx6f_ASAP7_75t_L g1058 ( 
.A(n_984),
.Y(n_1058)
);

NAND2xp5_ASAP7_75t_SL g1059 ( 
.A(n_994),
.B(n_926),
.Y(n_1059)
);

INVx1_ASAP7_75t_L g1060 ( 
.A(n_986),
.Y(n_1060)
);

INVx1_ASAP7_75t_L g1061 ( 
.A(n_986),
.Y(n_1061)
);

AND2x4_ASAP7_75t_L g1062 ( 
.A(n_968),
.B(n_877),
.Y(n_1062)
);

OAI21x1_ASAP7_75t_L g1063 ( 
.A1(n_963),
.A2(n_978),
.B(n_971),
.Y(n_1063)
);

AND2x2_ASAP7_75t_SL g1064 ( 
.A(n_994),
.B(n_631),
.Y(n_1064)
);

CKINVDCx5p33_ASAP7_75t_R g1065 ( 
.A(n_998),
.Y(n_1065)
);

INVx2_ASAP7_75t_L g1066 ( 
.A(n_947),
.Y(n_1066)
);

INVx1_ASAP7_75t_L g1067 ( 
.A(n_986),
.Y(n_1067)
);

AND3x1_ASAP7_75t_L g1068 ( 
.A(n_944),
.B(n_919),
.C(n_915),
.Y(n_1068)
);

BUFx6f_ASAP7_75t_L g1069 ( 
.A(n_986),
.Y(n_1069)
);

INVx2_ASAP7_75t_L g1070 ( 
.A(n_954),
.Y(n_1070)
);

AND2x4_ASAP7_75t_L g1071 ( 
.A(n_968),
.B(n_881),
.Y(n_1071)
);

AND2x4_ASAP7_75t_L g1072 ( 
.A(n_968),
.B(n_885),
.Y(n_1072)
);

INVx2_ASAP7_75t_L g1073 ( 
.A(n_954),
.Y(n_1073)
);

AND2x2_ASAP7_75t_L g1074 ( 
.A(n_1003),
.B(n_886),
.Y(n_1074)
);

NAND2xp5_ASAP7_75t_L g1075 ( 
.A(n_967),
.B(n_970),
.Y(n_1075)
);

INVx1_ASAP7_75t_L g1076 ( 
.A(n_986),
.Y(n_1076)
);

HB1xp67_ASAP7_75t_L g1077 ( 
.A(n_961),
.Y(n_1077)
);

BUFx6f_ASAP7_75t_L g1078 ( 
.A(n_1001),
.Y(n_1078)
);

NAND2xp5_ASAP7_75t_L g1079 ( 
.A(n_970),
.B(n_1001),
.Y(n_1079)
);

BUFx6f_ASAP7_75t_L g1080 ( 
.A(n_1001),
.Y(n_1080)
);

INVxp67_ASAP7_75t_L g1081 ( 
.A(n_977),
.Y(n_1081)
);

INVx3_ASAP7_75t_L g1082 ( 
.A(n_941),
.Y(n_1082)
);

HB1xp67_ASAP7_75t_L g1083 ( 
.A(n_965),
.Y(n_1083)
);

NAND2xp5_ASAP7_75t_L g1084 ( 
.A(n_1001),
.B(n_926),
.Y(n_1084)
);

INVx1_ASAP7_75t_L g1085 ( 
.A(n_1001),
.Y(n_1085)
);

INVx1_ASAP7_75t_L g1086 ( 
.A(n_974),
.Y(n_1086)
);

INVx1_ASAP7_75t_L g1087 ( 
.A(n_974),
.Y(n_1087)
);

AND2x2_ASAP7_75t_L g1088 ( 
.A(n_1003),
.B(n_888),
.Y(n_1088)
);

NAND2xp33_ASAP7_75t_L g1089 ( 
.A(n_987),
.B(n_715),
.Y(n_1089)
);

AND2x4_ASAP7_75t_L g1090 ( 
.A(n_975),
.B(n_889),
.Y(n_1090)
);

INVx3_ASAP7_75t_L g1091 ( 
.A(n_951),
.Y(n_1091)
);

INVx1_ASAP7_75t_L g1092 ( 
.A(n_1000),
.Y(n_1092)
);

BUFx2_ASAP7_75t_L g1093 ( 
.A(n_973),
.Y(n_1093)
);

BUFx6f_ASAP7_75t_L g1094 ( 
.A(n_1005),
.Y(n_1094)
);

INVx1_ASAP7_75t_L g1095 ( 
.A(n_1039),
.Y(n_1095)
);

INVx4_ASAP7_75t_L g1096 ( 
.A(n_1005),
.Y(n_1096)
);

NOR3xp33_ASAP7_75t_L g1097 ( 
.A(n_1047),
.B(n_1042),
.C(n_1030),
.Y(n_1097)
);

INVx1_ASAP7_75t_L g1098 ( 
.A(n_1039),
.Y(n_1098)
);

NAND2xp5_ASAP7_75t_SL g1099 ( 
.A(n_1064),
.B(n_950),
.Y(n_1099)
);

BUFx6f_ASAP7_75t_L g1100 ( 
.A(n_1005),
.Y(n_1100)
);

NAND2xp5_ASAP7_75t_L g1101 ( 
.A(n_1064),
.B(n_1008),
.Y(n_1101)
);

INVx3_ASAP7_75t_L g1102 ( 
.A(n_1024),
.Y(n_1102)
);

INVx1_ASAP7_75t_L g1103 ( 
.A(n_1092),
.Y(n_1103)
);

AOI22xp5_ASAP7_75t_L g1104 ( 
.A1(n_1042),
.A2(n_950),
.B1(n_896),
.B2(n_890),
.Y(n_1104)
);

NOR2xp33_ASAP7_75t_L g1105 ( 
.A(n_1029),
.B(n_890),
.Y(n_1105)
);

AOI22xp5_ASAP7_75t_L g1106 ( 
.A1(n_1031),
.A2(n_896),
.B1(n_846),
.B2(n_836),
.Y(n_1106)
);

OR2x6_ASAP7_75t_L g1107 ( 
.A(n_1093),
.B(n_973),
.Y(n_1107)
);

CKINVDCx5p33_ASAP7_75t_R g1108 ( 
.A(n_1065),
.Y(n_1108)
);

INVx2_ASAP7_75t_L g1109 ( 
.A(n_1007),
.Y(n_1109)
);

NAND2xp5_ASAP7_75t_L g1110 ( 
.A(n_1008),
.B(n_991),
.Y(n_1110)
);

NAND2xp5_ASAP7_75t_SL g1111 ( 
.A(n_1037),
.B(n_972),
.Y(n_1111)
);

INVx2_ASAP7_75t_L g1112 ( 
.A(n_1007),
.Y(n_1112)
);

INVx2_ASAP7_75t_L g1113 ( 
.A(n_1009),
.Y(n_1113)
);

INVx2_ASAP7_75t_L g1114 ( 
.A(n_1009),
.Y(n_1114)
);

INVx1_ASAP7_75t_L g1115 ( 
.A(n_1092),
.Y(n_1115)
);

INVx1_ASAP7_75t_L g1116 ( 
.A(n_1079),
.Y(n_1116)
);

AND2x2_ASAP7_75t_L g1117 ( 
.A(n_1011),
.B(n_882),
.Y(n_1117)
);

INVx8_ASAP7_75t_L g1118 ( 
.A(n_1010),
.Y(n_1118)
);

BUFx6f_ASAP7_75t_L g1119 ( 
.A(n_1005),
.Y(n_1119)
);

INVxp33_ASAP7_75t_L g1120 ( 
.A(n_1033),
.Y(n_1120)
);

OR2x6_ASAP7_75t_L g1121 ( 
.A(n_1093),
.B(n_989),
.Y(n_1121)
);

NOR2xp33_ASAP7_75t_R g1122 ( 
.A(n_1038),
.B(n_945),
.Y(n_1122)
);

INVx1_ASAP7_75t_L g1123 ( 
.A(n_1086),
.Y(n_1123)
);

OAI22xp33_ASAP7_75t_L g1124 ( 
.A1(n_1083),
.A2(n_830),
.B1(n_806),
.B2(n_751),
.Y(n_1124)
);

INVx1_ASAP7_75t_L g1125 ( 
.A(n_1086),
.Y(n_1125)
);

BUFx2_ASAP7_75t_L g1126 ( 
.A(n_1018),
.Y(n_1126)
);

INVx2_ASAP7_75t_L g1127 ( 
.A(n_1016),
.Y(n_1127)
);

INVx3_ASAP7_75t_L g1128 ( 
.A(n_1024),
.Y(n_1128)
);

INVx2_ASAP7_75t_SL g1129 ( 
.A(n_1018),
.Y(n_1129)
);

INVx3_ASAP7_75t_L g1130 ( 
.A(n_1024),
.Y(n_1130)
);

INVx1_ASAP7_75t_L g1131 ( 
.A(n_1087),
.Y(n_1131)
);

INVx2_ASAP7_75t_L g1132 ( 
.A(n_1016),
.Y(n_1132)
);

AND2x2_ASAP7_75t_L g1133 ( 
.A(n_1013),
.B(n_914),
.Y(n_1133)
);

INVx1_ASAP7_75t_L g1134 ( 
.A(n_1087),
.Y(n_1134)
);

INVx1_ASAP7_75t_L g1135 ( 
.A(n_1074),
.Y(n_1135)
);

NOR2xp33_ASAP7_75t_L g1136 ( 
.A(n_1046),
.B(n_975),
.Y(n_1136)
);

OAI22xp5_ASAP7_75t_L g1137 ( 
.A1(n_1028),
.A2(n_1084),
.B1(n_1023),
.B2(n_1059),
.Y(n_1137)
);

INVx1_ASAP7_75t_SL g1138 ( 
.A(n_1013),
.Y(n_1138)
);

INVx1_ASAP7_75t_L g1139 ( 
.A(n_1074),
.Y(n_1139)
);

NOR3xp33_ASAP7_75t_L g1140 ( 
.A(n_1019),
.B(n_813),
.C(n_799),
.Y(n_1140)
);

NOR2xp33_ASAP7_75t_L g1141 ( 
.A(n_1021),
.B(n_979),
.Y(n_1141)
);

INVx1_ASAP7_75t_L g1142 ( 
.A(n_1088),
.Y(n_1142)
);

BUFx10_ASAP7_75t_L g1143 ( 
.A(n_1065),
.Y(n_1143)
);

INVx2_ASAP7_75t_L g1144 ( 
.A(n_1025),
.Y(n_1144)
);

BUFx6f_ASAP7_75t_L g1145 ( 
.A(n_1005),
.Y(n_1145)
);

INVx5_ASAP7_75t_L g1146 ( 
.A(n_1015),
.Y(n_1146)
);

AND3x1_ASAP7_75t_L g1147 ( 
.A(n_1077),
.B(n_751),
.C(n_680),
.Y(n_1147)
);

INVx2_ASAP7_75t_L g1148 ( 
.A(n_1025),
.Y(n_1148)
);

INVx1_ASAP7_75t_L g1149 ( 
.A(n_1088),
.Y(n_1149)
);

INVx1_ASAP7_75t_L g1150 ( 
.A(n_1017),
.Y(n_1150)
);

INVx1_ASAP7_75t_L g1151 ( 
.A(n_1045),
.Y(n_1151)
);

AOI22xp33_ASAP7_75t_L g1152 ( 
.A1(n_1044),
.A2(n_836),
.B1(n_846),
.B2(n_830),
.Y(n_1152)
);

INVx2_ASAP7_75t_L g1153 ( 
.A(n_1027),
.Y(n_1153)
);

INVx2_ASAP7_75t_L g1154 ( 
.A(n_1027),
.Y(n_1154)
);

OR2x6_ASAP7_75t_L g1155 ( 
.A(n_1049),
.B(n_989),
.Y(n_1155)
);

AOI21x1_ASAP7_75t_L g1156 ( 
.A1(n_1020),
.A2(n_978),
.B(n_987),
.Y(n_1156)
);

INVx1_ASAP7_75t_L g1157 ( 
.A(n_1051),
.Y(n_1157)
);

INVx4_ASAP7_75t_L g1158 ( 
.A(n_1015),
.Y(n_1158)
);

INVx2_ASAP7_75t_L g1159 ( 
.A(n_1036),
.Y(n_1159)
);

NAND2xp5_ASAP7_75t_L g1160 ( 
.A(n_1019),
.B(n_1075),
.Y(n_1160)
);

INVx3_ASAP7_75t_L g1161 ( 
.A(n_1053),
.Y(n_1161)
);

INVx2_ASAP7_75t_SL g1162 ( 
.A(n_1010),
.Y(n_1162)
);

INVx2_ASAP7_75t_L g1163 ( 
.A(n_1036),
.Y(n_1163)
);

INVx1_ASAP7_75t_L g1164 ( 
.A(n_1040),
.Y(n_1164)
);

AOI22xp33_ASAP7_75t_L g1165 ( 
.A1(n_1044),
.A2(n_996),
.B1(n_1000),
.B2(n_993),
.Y(n_1165)
);

BUFx8_ASAP7_75t_SL g1166 ( 
.A(n_1022),
.Y(n_1166)
);

NAND2xp5_ASAP7_75t_L g1167 ( 
.A(n_1010),
.B(n_991),
.Y(n_1167)
);

NAND2xp5_ASAP7_75t_SL g1168 ( 
.A(n_1015),
.B(n_972),
.Y(n_1168)
);

INVx1_ASAP7_75t_L g1169 ( 
.A(n_1040),
.Y(n_1169)
);

INVx2_ASAP7_75t_L g1170 ( 
.A(n_1054),
.Y(n_1170)
);

AOI22xp33_ASAP7_75t_L g1171 ( 
.A1(n_1055),
.A2(n_996),
.B1(n_993),
.B2(n_808),
.Y(n_1171)
);

INVx2_ASAP7_75t_L g1172 ( 
.A(n_1054),
.Y(n_1172)
);

NAND2xp5_ASAP7_75t_SL g1173 ( 
.A(n_1015),
.B(n_972),
.Y(n_1173)
);

NAND2xp5_ASAP7_75t_L g1174 ( 
.A(n_1012),
.B(n_979),
.Y(n_1174)
);

NAND2xp5_ASAP7_75t_SL g1175 ( 
.A(n_1015),
.B(n_972),
.Y(n_1175)
);

INVx2_ASAP7_75t_L g1176 ( 
.A(n_1054),
.Y(n_1176)
);

INVx1_ASAP7_75t_L g1177 ( 
.A(n_1054),
.Y(n_1177)
);

NAND2xp5_ASAP7_75t_SL g1178 ( 
.A(n_1034),
.B(n_972),
.Y(n_1178)
);

AO21x2_ASAP7_75t_L g1179 ( 
.A1(n_1055),
.A2(n_1056),
.B(n_1063),
.Y(n_1179)
);

NOR2xp33_ASAP7_75t_L g1180 ( 
.A(n_1012),
.B(n_933),
.Y(n_1180)
);

NAND2xp5_ASAP7_75t_SL g1181 ( 
.A(n_1034),
.B(n_990),
.Y(n_1181)
);

BUFx6f_ASAP7_75t_L g1182 ( 
.A(n_1034),
.Y(n_1182)
);

OR2x2_ASAP7_75t_L g1183 ( 
.A(n_1081),
.B(n_891),
.Y(n_1183)
);

INVx2_ASAP7_75t_L g1184 ( 
.A(n_1043),
.Y(n_1184)
);

INVx2_ASAP7_75t_L g1185 ( 
.A(n_1043),
.Y(n_1185)
);

INVx1_ASAP7_75t_SL g1186 ( 
.A(n_1050),
.Y(n_1186)
);

BUFx6f_ASAP7_75t_SL g1187 ( 
.A(n_1012),
.Y(n_1187)
);

INVx1_ASAP7_75t_L g1188 ( 
.A(n_1090),
.Y(n_1188)
);

AO21x2_ASAP7_75t_L g1189 ( 
.A1(n_1056),
.A2(n_894),
.B(n_893),
.Y(n_1189)
);

AND2x2_ASAP7_75t_L g1190 ( 
.A(n_1050),
.B(n_945),
.Y(n_1190)
);

INVx2_ASAP7_75t_L g1191 ( 
.A(n_1048),
.Y(n_1191)
);

AOI22xp33_ASAP7_75t_L g1192 ( 
.A1(n_1041),
.A2(n_808),
.B1(n_798),
.B2(n_841),
.Y(n_1192)
);

INVx2_ASAP7_75t_L g1193 ( 
.A(n_1048),
.Y(n_1193)
);

INVx4_ASAP7_75t_L g1194 ( 
.A(n_1034),
.Y(n_1194)
);

INVx2_ASAP7_75t_L g1195 ( 
.A(n_1066),
.Y(n_1195)
);

INVx1_ASAP7_75t_L g1196 ( 
.A(n_1090),
.Y(n_1196)
);

INVx1_ASAP7_75t_L g1197 ( 
.A(n_1090),
.Y(n_1197)
);

INVx1_ASAP7_75t_L g1198 ( 
.A(n_1035),
.Y(n_1198)
);

OAI22xp5_ASAP7_75t_L g1199 ( 
.A1(n_1053),
.A2(n_779),
.B1(n_781),
.B2(n_603),
.Y(n_1199)
);

AND2x6_ASAP7_75t_L g1200 ( 
.A(n_1020),
.B(n_661),
.Y(n_1200)
);

INVx1_ASAP7_75t_L g1201 ( 
.A(n_1035),
.Y(n_1201)
);

INVx1_ASAP7_75t_L g1202 ( 
.A(n_1041),
.Y(n_1202)
);

NAND2xp5_ASAP7_75t_SL g1203 ( 
.A(n_1034),
.B(n_990),
.Y(n_1203)
);

NOR2x1p5_ASAP7_75t_L g1204 ( 
.A(n_1022),
.B(n_938),
.Y(n_1204)
);

INVx2_ASAP7_75t_L g1205 ( 
.A(n_1066),
.Y(n_1205)
);

INVx1_ASAP7_75t_L g1206 ( 
.A(n_1041),
.Y(n_1206)
);

INVx2_ASAP7_75t_L g1207 ( 
.A(n_1070),
.Y(n_1207)
);

INVx3_ASAP7_75t_L g1208 ( 
.A(n_1053),
.Y(n_1208)
);

INVx3_ASAP7_75t_L g1209 ( 
.A(n_1082),
.Y(n_1209)
);

INVx1_ASAP7_75t_L g1210 ( 
.A(n_1052),
.Y(n_1210)
);

INVx2_ASAP7_75t_L g1211 ( 
.A(n_1070),
.Y(n_1211)
);

NAND2xp5_ASAP7_75t_L g1212 ( 
.A(n_1052),
.B(n_933),
.Y(n_1212)
);

AOI22xp33_ASAP7_75t_L g1213 ( 
.A1(n_1052),
.A2(n_798),
.B1(n_633),
.B2(n_647),
.Y(n_1213)
);

INVx1_ASAP7_75t_L g1214 ( 
.A(n_1057),
.Y(n_1214)
);

INVx2_ASAP7_75t_L g1215 ( 
.A(n_1073),
.Y(n_1215)
);

INVx1_ASAP7_75t_L g1216 ( 
.A(n_1057),
.Y(n_1216)
);

CKINVDCx5p33_ASAP7_75t_R g1217 ( 
.A(n_1022),
.Y(n_1217)
);

INVx2_ASAP7_75t_SL g1218 ( 
.A(n_1062),
.Y(n_1218)
);

OR2x2_ASAP7_75t_L g1219 ( 
.A(n_1062),
.B(n_891),
.Y(n_1219)
);

OR2x2_ASAP7_75t_L g1220 ( 
.A(n_1062),
.B(n_837),
.Y(n_1220)
);

INVx1_ASAP7_75t_L g1221 ( 
.A(n_1060),
.Y(n_1221)
);

NAND2xp5_ASAP7_75t_L g1222 ( 
.A(n_1071),
.B(n_700),
.Y(n_1222)
);

AND2x2_ASAP7_75t_L g1223 ( 
.A(n_1071),
.B(n_851),
.Y(n_1223)
);

BUFx3_ASAP7_75t_L g1224 ( 
.A(n_1058),
.Y(n_1224)
);

AND3x1_ASAP7_75t_L g1225 ( 
.A(n_1038),
.B(n_647),
.C(n_631),
.Y(n_1225)
);

INVx1_ASAP7_75t_L g1226 ( 
.A(n_1060),
.Y(n_1226)
);

NAND2xp5_ASAP7_75t_L g1227 ( 
.A(n_1071),
.B(n_1072),
.Y(n_1227)
);

NAND2xp5_ASAP7_75t_L g1228 ( 
.A(n_1072),
.B(n_1082),
.Y(n_1228)
);

BUFx3_ASAP7_75t_L g1229 ( 
.A(n_1058),
.Y(n_1229)
);

NAND2xp5_ASAP7_75t_L g1230 ( 
.A(n_1072),
.B(n_769),
.Y(n_1230)
);

AOI22xp33_ASAP7_75t_SL g1231 ( 
.A1(n_1068),
.A2(n_643),
.B1(n_699),
.B2(n_605),
.Y(n_1231)
);

HB1xp67_ASAP7_75t_L g1232 ( 
.A(n_1126),
.Y(n_1232)
);

INVx2_ASAP7_75t_L g1233 ( 
.A(n_1184),
.Y(n_1233)
);

NAND2xp5_ASAP7_75t_SL g1234 ( 
.A(n_1097),
.B(n_1218),
.Y(n_1234)
);

NAND2xp5_ASAP7_75t_L g1235 ( 
.A(n_1116),
.B(n_1063),
.Y(n_1235)
);

INVx2_ASAP7_75t_L g1236 ( 
.A(n_1184),
.Y(n_1236)
);

AND2x2_ASAP7_75t_L g1237 ( 
.A(n_1186),
.B(n_851),
.Y(n_1237)
);

INVx1_ASAP7_75t_L g1238 ( 
.A(n_1103),
.Y(n_1238)
);

AND2x4_ASAP7_75t_L g1239 ( 
.A(n_1227),
.B(n_1082),
.Y(n_1239)
);

HB1xp67_ASAP7_75t_L g1240 ( 
.A(n_1129),
.Y(n_1240)
);

INVx1_ASAP7_75t_L g1241 ( 
.A(n_1115),
.Y(n_1241)
);

INVx1_ASAP7_75t_L g1242 ( 
.A(n_1123),
.Y(n_1242)
);

INVx2_ASAP7_75t_SL g1243 ( 
.A(n_1190),
.Y(n_1243)
);

NOR2xp33_ASAP7_75t_L g1244 ( 
.A(n_1105),
.B(n_983),
.Y(n_1244)
);

INVx1_ASAP7_75t_L g1245 ( 
.A(n_1125),
.Y(n_1245)
);

INVx2_ASAP7_75t_L g1246 ( 
.A(n_1185),
.Y(n_1246)
);

INVx2_ASAP7_75t_L g1247 ( 
.A(n_1185),
.Y(n_1247)
);

NOR2xp33_ASAP7_75t_L g1248 ( 
.A(n_1105),
.B(n_943),
.Y(n_1248)
);

BUFx4f_ASAP7_75t_L g1249 ( 
.A(n_1107),
.Y(n_1249)
);

NAND2x1p5_ASAP7_75t_L g1250 ( 
.A(n_1204),
.B(n_1061),
.Y(n_1250)
);

INVx2_ASAP7_75t_L g1251 ( 
.A(n_1191),
.Y(n_1251)
);

INVx2_ASAP7_75t_L g1252 ( 
.A(n_1191),
.Y(n_1252)
);

INVx1_ASAP7_75t_L g1253 ( 
.A(n_1131),
.Y(n_1253)
);

INVx3_ASAP7_75t_L g1254 ( 
.A(n_1096),
.Y(n_1254)
);

NAND2xp5_ASAP7_75t_L g1255 ( 
.A(n_1160),
.B(n_1061),
.Y(n_1255)
);

NAND2xp5_ASAP7_75t_L g1256 ( 
.A(n_1097),
.B(n_1067),
.Y(n_1256)
);

INVxp67_ASAP7_75t_L g1257 ( 
.A(n_1117),
.Y(n_1257)
);

NAND2xp5_ASAP7_75t_SL g1258 ( 
.A(n_1162),
.B(n_1058),
.Y(n_1258)
);

BUFx3_ASAP7_75t_L g1259 ( 
.A(n_1166),
.Y(n_1259)
);

OAI21xp33_ASAP7_75t_L g1260 ( 
.A1(n_1180),
.A2(n_696),
.B(n_655),
.Y(n_1260)
);

BUFx3_ASAP7_75t_L g1261 ( 
.A(n_1166),
.Y(n_1261)
);

INVx8_ASAP7_75t_L g1262 ( 
.A(n_1118),
.Y(n_1262)
);

INVx1_ASAP7_75t_L g1263 ( 
.A(n_1134),
.Y(n_1263)
);

INVx4_ASAP7_75t_L g1264 ( 
.A(n_1118),
.Y(n_1264)
);

NOR2xp33_ASAP7_75t_L g1265 ( 
.A(n_1099),
.B(n_943),
.Y(n_1265)
);

NOR2xp33_ASAP7_75t_L g1266 ( 
.A(n_1099),
.B(n_948),
.Y(n_1266)
);

BUFx8_ASAP7_75t_SL g1267 ( 
.A(n_1108),
.Y(n_1267)
);

INVx1_ASAP7_75t_L g1268 ( 
.A(n_1095),
.Y(n_1268)
);

BUFx10_ASAP7_75t_L g1269 ( 
.A(n_1180),
.Y(n_1269)
);

INVx1_ASAP7_75t_L g1270 ( 
.A(n_1098),
.Y(n_1270)
);

INVx5_ASAP7_75t_L g1271 ( 
.A(n_1118),
.Y(n_1271)
);

AND2x2_ASAP7_75t_SL g1272 ( 
.A(n_1152),
.B(n_942),
.Y(n_1272)
);

INVx2_ASAP7_75t_L g1273 ( 
.A(n_1211),
.Y(n_1273)
);

AND2x6_ASAP7_75t_L g1274 ( 
.A(n_1202),
.B(n_1026),
.Y(n_1274)
);

INVx1_ASAP7_75t_L g1275 ( 
.A(n_1164),
.Y(n_1275)
);

NAND2x1p5_ASAP7_75t_L g1276 ( 
.A(n_1146),
.B(n_1058),
.Y(n_1276)
);

INVx2_ASAP7_75t_L g1277 ( 
.A(n_1211),
.Y(n_1277)
);

INVx1_ASAP7_75t_L g1278 ( 
.A(n_1169),
.Y(n_1278)
);

INVx1_ASAP7_75t_L g1279 ( 
.A(n_1150),
.Y(n_1279)
);

INVx1_ASAP7_75t_SL g1280 ( 
.A(n_1133),
.Y(n_1280)
);

INVx1_ASAP7_75t_L g1281 ( 
.A(n_1151),
.Y(n_1281)
);

NAND2x1p5_ASAP7_75t_L g1282 ( 
.A(n_1146),
.B(n_1058),
.Y(n_1282)
);

AND2x2_ASAP7_75t_L g1283 ( 
.A(n_1138),
.B(n_895),
.Y(n_1283)
);

INVx2_ASAP7_75t_L g1284 ( 
.A(n_1215),
.Y(n_1284)
);

INVx1_ASAP7_75t_L g1285 ( 
.A(n_1157),
.Y(n_1285)
);

AND2x2_ASAP7_75t_L g1286 ( 
.A(n_1223),
.B(n_897),
.Y(n_1286)
);

AND2x6_ASAP7_75t_L g1287 ( 
.A(n_1206),
.B(n_1026),
.Y(n_1287)
);

AND2x6_ASAP7_75t_L g1288 ( 
.A(n_1210),
.B(n_1006),
.Y(n_1288)
);

OR2x2_ASAP7_75t_L g1289 ( 
.A(n_1183),
.B(n_964),
.Y(n_1289)
);

AND2x4_ASAP7_75t_L g1290 ( 
.A(n_1188),
.B(n_1067),
.Y(n_1290)
);

BUFx6f_ASAP7_75t_L g1291 ( 
.A(n_1094),
.Y(n_1291)
);

INVx2_ASAP7_75t_L g1292 ( 
.A(n_1215),
.Y(n_1292)
);

INVx4_ASAP7_75t_L g1293 ( 
.A(n_1107),
.Y(n_1293)
);

AND2x6_ASAP7_75t_L g1294 ( 
.A(n_1177),
.B(n_1006),
.Y(n_1294)
);

INVx1_ASAP7_75t_L g1295 ( 
.A(n_1135),
.Y(n_1295)
);

BUFx3_ASAP7_75t_L g1296 ( 
.A(n_1143),
.Y(n_1296)
);

BUFx6f_ASAP7_75t_L g1297 ( 
.A(n_1094),
.Y(n_1297)
);

HB1xp67_ASAP7_75t_L g1298 ( 
.A(n_1187),
.Y(n_1298)
);

INVx4_ASAP7_75t_L g1299 ( 
.A(n_1107),
.Y(n_1299)
);

BUFx6f_ASAP7_75t_L g1300 ( 
.A(n_1094),
.Y(n_1300)
);

NAND2xp5_ASAP7_75t_L g1301 ( 
.A(n_1136),
.B(n_1076),
.Y(n_1301)
);

AND2x6_ASAP7_75t_L g1302 ( 
.A(n_1170),
.B(n_1014),
.Y(n_1302)
);

INVx1_ASAP7_75t_L g1303 ( 
.A(n_1139),
.Y(n_1303)
);

INVx3_ASAP7_75t_L g1304 ( 
.A(n_1096),
.Y(n_1304)
);

NAND2xp5_ASAP7_75t_L g1305 ( 
.A(n_1136),
.B(n_1076),
.Y(n_1305)
);

AND2x4_ASAP7_75t_L g1306 ( 
.A(n_1196),
.B(n_1085),
.Y(n_1306)
);

BUFx6f_ASAP7_75t_L g1307 ( 
.A(n_1094),
.Y(n_1307)
);

INVx1_ASAP7_75t_L g1308 ( 
.A(n_1142),
.Y(n_1308)
);

AND2x6_ASAP7_75t_L g1309 ( 
.A(n_1170),
.B(n_1014),
.Y(n_1309)
);

AND2x4_ASAP7_75t_L g1310 ( 
.A(n_1197),
.B(n_1085),
.Y(n_1310)
);

BUFx3_ASAP7_75t_L g1311 ( 
.A(n_1143),
.Y(n_1311)
);

NAND2xp5_ASAP7_75t_SL g1312 ( 
.A(n_1101),
.B(n_1069),
.Y(n_1312)
);

BUFx3_ASAP7_75t_L g1313 ( 
.A(n_1217),
.Y(n_1313)
);

BUFx2_ASAP7_75t_L g1314 ( 
.A(n_1122),
.Y(n_1314)
);

NOR2xp33_ASAP7_75t_L g1315 ( 
.A(n_1120),
.B(n_980),
.Y(n_1315)
);

NOR2xp33_ASAP7_75t_L g1316 ( 
.A(n_1120),
.B(n_942),
.Y(n_1316)
);

INVx3_ASAP7_75t_L g1317 ( 
.A(n_1158),
.Y(n_1317)
);

AND2x4_ASAP7_75t_L g1318 ( 
.A(n_1121),
.B(n_898),
.Y(n_1318)
);

BUFx6f_ASAP7_75t_L g1319 ( 
.A(n_1100),
.Y(n_1319)
);

NAND2xp5_ASAP7_75t_L g1320 ( 
.A(n_1141),
.B(n_1069),
.Y(n_1320)
);

INVx1_ASAP7_75t_L g1321 ( 
.A(n_1149),
.Y(n_1321)
);

AND2x4_ASAP7_75t_L g1322 ( 
.A(n_1121),
.B(n_900),
.Y(n_1322)
);

INVx3_ASAP7_75t_L g1323 ( 
.A(n_1158),
.Y(n_1323)
);

INVx1_ASAP7_75t_L g1324 ( 
.A(n_1109),
.Y(n_1324)
);

AND2x2_ASAP7_75t_L g1325 ( 
.A(n_1152),
.B(n_902),
.Y(n_1325)
);

INVx3_ASAP7_75t_L g1326 ( 
.A(n_1194),
.Y(n_1326)
);

AOI22xp5_ASAP7_75t_L g1327 ( 
.A1(n_1140),
.A2(n_1089),
.B1(n_1078),
.B2(n_1080),
.Y(n_1327)
);

NAND2xp5_ASAP7_75t_SL g1328 ( 
.A(n_1137),
.B(n_1069),
.Y(n_1328)
);

BUFx3_ASAP7_75t_L g1329 ( 
.A(n_1121),
.Y(n_1329)
);

INVx1_ASAP7_75t_L g1330 ( 
.A(n_1109),
.Y(n_1330)
);

INVx1_ASAP7_75t_L g1331 ( 
.A(n_1112),
.Y(n_1331)
);

INVx2_ASAP7_75t_L g1332 ( 
.A(n_1112),
.Y(n_1332)
);

INVx3_ASAP7_75t_L g1333 ( 
.A(n_1194),
.Y(n_1333)
);

AND2x2_ASAP7_75t_L g1334 ( 
.A(n_1104),
.B(n_903),
.Y(n_1334)
);

BUFx6f_ASAP7_75t_L g1335 ( 
.A(n_1100),
.Y(n_1335)
);

AND2x4_ASAP7_75t_L g1336 ( 
.A(n_1181),
.B(n_905),
.Y(n_1336)
);

AOI22xp5_ASAP7_75t_L g1337 ( 
.A1(n_1140),
.A2(n_1089),
.B1(n_1078),
.B2(n_1080),
.Y(n_1337)
);

INVx1_ASAP7_75t_L g1338 ( 
.A(n_1113),
.Y(n_1338)
);

BUFx6f_ASAP7_75t_L g1339 ( 
.A(n_1100),
.Y(n_1339)
);

BUFx6f_ASAP7_75t_L g1340 ( 
.A(n_1100),
.Y(n_1340)
);

INVx2_ASAP7_75t_L g1341 ( 
.A(n_1113),
.Y(n_1341)
);

BUFx2_ASAP7_75t_L g1342 ( 
.A(n_1122),
.Y(n_1342)
);

NOR2xp33_ASAP7_75t_L g1343 ( 
.A(n_1220),
.B(n_1069),
.Y(n_1343)
);

INVx1_ASAP7_75t_L g1344 ( 
.A(n_1127),
.Y(n_1344)
);

INVx1_ASAP7_75t_L g1345 ( 
.A(n_1127),
.Y(n_1345)
);

BUFx3_ASAP7_75t_L g1346 ( 
.A(n_1155),
.Y(n_1346)
);

NAND2xp33_ASAP7_75t_L g1347 ( 
.A(n_1228),
.B(n_1069),
.Y(n_1347)
);

NAND2xp5_ASAP7_75t_L g1348 ( 
.A(n_1141),
.B(n_1165),
.Y(n_1348)
);

AND2x2_ASAP7_75t_L g1349 ( 
.A(n_1106),
.B(n_906),
.Y(n_1349)
);

AND2x4_ASAP7_75t_L g1350 ( 
.A(n_1181),
.B(n_907),
.Y(n_1350)
);

INVx1_ASAP7_75t_L g1351 ( 
.A(n_1132),
.Y(n_1351)
);

INVx2_ASAP7_75t_L g1352 ( 
.A(n_1132),
.Y(n_1352)
);

INVx1_ASAP7_75t_L g1353 ( 
.A(n_1148),
.Y(n_1353)
);

NOR2xp33_ASAP7_75t_SL g1354 ( 
.A(n_1187),
.B(n_793),
.Y(n_1354)
);

INVx1_ASAP7_75t_L g1355 ( 
.A(n_1148),
.Y(n_1355)
);

NOR2xp33_ASAP7_75t_L g1356 ( 
.A(n_1219),
.B(n_1078),
.Y(n_1356)
);

INVx3_ASAP7_75t_L g1357 ( 
.A(n_1224),
.Y(n_1357)
);

AND2x2_ASAP7_75t_L g1358 ( 
.A(n_1212),
.B(n_908),
.Y(n_1358)
);

BUFx3_ASAP7_75t_L g1359 ( 
.A(n_1155),
.Y(n_1359)
);

INVx2_ASAP7_75t_L g1360 ( 
.A(n_1153),
.Y(n_1360)
);

OR2x6_ASAP7_75t_L g1361 ( 
.A(n_1155),
.B(n_1078),
.Y(n_1361)
);

NAND2xp5_ASAP7_75t_L g1362 ( 
.A(n_1165),
.B(n_1078),
.Y(n_1362)
);

BUFx3_ASAP7_75t_L g1363 ( 
.A(n_1224),
.Y(n_1363)
);

INVx4_ASAP7_75t_L g1364 ( 
.A(n_1146),
.Y(n_1364)
);

NAND2xp5_ASAP7_75t_L g1365 ( 
.A(n_1153),
.B(n_1080),
.Y(n_1365)
);

AOI22xp5_ASAP7_75t_L g1366 ( 
.A1(n_1171),
.A2(n_1080),
.B1(n_774),
.B2(n_795),
.Y(n_1366)
);

BUFx3_ASAP7_75t_L g1367 ( 
.A(n_1229),
.Y(n_1367)
);

NAND2xp5_ASAP7_75t_L g1368 ( 
.A(n_1154),
.B(n_1080),
.Y(n_1368)
);

INVx4_ASAP7_75t_L g1369 ( 
.A(n_1146),
.Y(n_1369)
);

NAND2xp5_ASAP7_75t_L g1370 ( 
.A(n_1159),
.B(n_1073),
.Y(n_1370)
);

NOR2xp33_ASAP7_75t_L g1371 ( 
.A(n_1124),
.B(n_1091),
.Y(n_1371)
);

INVx1_ASAP7_75t_L g1372 ( 
.A(n_1159),
.Y(n_1372)
);

AND2x2_ASAP7_75t_L g1373 ( 
.A(n_1192),
.B(n_911),
.Y(n_1373)
);

AND2x4_ASAP7_75t_L g1374 ( 
.A(n_1203),
.B(n_916),
.Y(n_1374)
);

OAI221xp5_ASAP7_75t_L g1375 ( 
.A1(n_1213),
.A2(n_655),
.B1(n_723),
.B2(n_703),
.C(n_696),
.Y(n_1375)
);

NOR2xp33_ASAP7_75t_L g1376 ( 
.A(n_1124),
.B(n_1091),
.Y(n_1376)
);

NAND3xp33_ASAP7_75t_L g1377 ( 
.A(n_1171),
.B(n_816),
.C(n_719),
.Y(n_1377)
);

INVx1_ASAP7_75t_L g1378 ( 
.A(n_1163),
.Y(n_1378)
);

AOI22xp5_ASAP7_75t_L g1379 ( 
.A1(n_1225),
.A2(n_797),
.B1(n_829),
.B2(n_604),
.Y(n_1379)
);

INVx3_ASAP7_75t_L g1380 ( 
.A(n_1229),
.Y(n_1380)
);

INVx4_ASAP7_75t_L g1381 ( 
.A(n_1119),
.Y(n_1381)
);

INVx2_ASAP7_75t_L g1382 ( 
.A(n_1163),
.Y(n_1382)
);

BUFx6f_ASAP7_75t_L g1383 ( 
.A(n_1119),
.Y(n_1383)
);

NAND2xp5_ASAP7_75t_SL g1384 ( 
.A(n_1167),
.B(n_1091),
.Y(n_1384)
);

BUFx3_ASAP7_75t_L g1385 ( 
.A(n_1214),
.Y(n_1385)
);

CKINVDCx5p33_ASAP7_75t_R g1386 ( 
.A(n_1203),
.Y(n_1386)
);

INVx2_ASAP7_75t_L g1387 ( 
.A(n_1193),
.Y(n_1387)
);

AND2x4_ASAP7_75t_L g1388 ( 
.A(n_1174),
.B(n_920),
.Y(n_1388)
);

NAND2xp5_ASAP7_75t_L g1389 ( 
.A(n_1114),
.B(n_1032),
.Y(n_1389)
);

INVx1_ASAP7_75t_L g1390 ( 
.A(n_1144),
.Y(n_1390)
);

AND2x2_ASAP7_75t_L g1391 ( 
.A(n_1192),
.B(n_921),
.Y(n_1391)
);

INVx2_ASAP7_75t_SL g1392 ( 
.A(n_1222),
.Y(n_1392)
);

NAND2xp5_ASAP7_75t_L g1393 ( 
.A(n_1189),
.B(n_1032),
.Y(n_1393)
);

HB1xp67_ASAP7_75t_L g1394 ( 
.A(n_1230),
.Y(n_1394)
);

AND2x2_ASAP7_75t_L g1395 ( 
.A(n_1213),
.B(n_922),
.Y(n_1395)
);

AND2x4_ASAP7_75t_L g1396 ( 
.A(n_1110),
.B(n_923),
.Y(n_1396)
);

INVx1_ASAP7_75t_L g1397 ( 
.A(n_1216),
.Y(n_1397)
);

INVx3_ASAP7_75t_L g1398 ( 
.A(n_1119),
.Y(n_1398)
);

INVx1_ASAP7_75t_L g1399 ( 
.A(n_1221),
.Y(n_1399)
);

INVx1_ASAP7_75t_L g1400 ( 
.A(n_1226),
.Y(n_1400)
);

INVx1_ASAP7_75t_L g1401 ( 
.A(n_1195),
.Y(n_1401)
);

AND2x2_ASAP7_75t_L g1402 ( 
.A(n_1231),
.B(n_924),
.Y(n_1402)
);

INVx3_ASAP7_75t_L g1403 ( 
.A(n_1119),
.Y(n_1403)
);

NAND3xp33_ASAP7_75t_L g1404 ( 
.A(n_1147),
.B(n_819),
.C(n_719),
.Y(n_1404)
);

INVx1_ASAP7_75t_L g1405 ( 
.A(n_1205),
.Y(n_1405)
);

AOI22xp33_ASAP7_75t_L g1406 ( 
.A1(n_1231),
.A2(n_1207),
.B1(n_1189),
.B2(n_1176),
.Y(n_1406)
);

INVx1_ASAP7_75t_SL g1407 ( 
.A(n_1145),
.Y(n_1407)
);

INVx8_ASAP7_75t_L g1408 ( 
.A(n_1200),
.Y(n_1408)
);

INVxp67_ASAP7_75t_SL g1409 ( 
.A(n_1145),
.Y(n_1409)
);

INVx2_ASAP7_75t_L g1410 ( 
.A(n_1172),
.Y(n_1410)
);

NAND2xp33_ASAP7_75t_L g1411 ( 
.A(n_1102),
.B(n_603),
.Y(n_1411)
);

NAND2xp5_ASAP7_75t_L g1412 ( 
.A(n_1209),
.B(n_1032),
.Y(n_1412)
);

CKINVDCx20_ASAP7_75t_R g1413 ( 
.A(n_1199),
.Y(n_1413)
);

INVx1_ASAP7_75t_L g1414 ( 
.A(n_1156),
.Y(n_1414)
);

INVxp67_ASAP7_75t_L g1415 ( 
.A(n_1179),
.Y(n_1415)
);

INVx2_ASAP7_75t_L g1416 ( 
.A(n_1172),
.Y(n_1416)
);

AND2x2_ASAP7_75t_L g1417 ( 
.A(n_1176),
.B(n_925),
.Y(n_1417)
);

NAND2xp5_ASAP7_75t_L g1418 ( 
.A(n_1209),
.B(n_703),
.Y(n_1418)
);

OR2x2_ASAP7_75t_SL g1419 ( 
.A(n_1145),
.B(n_912),
.Y(n_1419)
);

AND3x4_ASAP7_75t_L g1420 ( 
.A(n_1102),
.B(n_754),
.C(n_723),
.Y(n_1420)
);

INVx1_ASAP7_75t_L g1421 ( 
.A(n_1208),
.Y(n_1421)
);

OAI22xp5_ASAP7_75t_L g1422 ( 
.A1(n_1128),
.A2(n_1161),
.B1(n_1130),
.B2(n_1208),
.Y(n_1422)
);

INVx1_ASAP7_75t_SL g1423 ( 
.A(n_1145),
.Y(n_1423)
);

INVx1_ASAP7_75t_L g1424 ( 
.A(n_1128),
.Y(n_1424)
);

BUFx6f_ASAP7_75t_L g1425 ( 
.A(n_1182),
.Y(n_1425)
);

NOR2xp33_ASAP7_75t_L g1426 ( 
.A(n_1130),
.B(n_779),
.Y(n_1426)
);

AOI22xp33_ASAP7_75t_L g1427 ( 
.A1(n_1200),
.A2(n_699),
.B1(n_702),
.B2(n_643),
.Y(n_1427)
);

INVx1_ASAP7_75t_L g1428 ( 
.A(n_1161),
.Y(n_1428)
);

NAND2xp5_ASAP7_75t_L g1429 ( 
.A(n_1179),
.B(n_754),
.Y(n_1429)
);

BUFx2_ASAP7_75t_L g1430 ( 
.A(n_1200),
.Y(n_1430)
);

INVx5_ASAP7_75t_L g1431 ( 
.A(n_1182),
.Y(n_1431)
);

BUFx3_ASAP7_75t_L g1432 ( 
.A(n_1182),
.Y(n_1432)
);

NOR2xp33_ASAP7_75t_L g1433 ( 
.A(n_1248),
.B(n_1111),
.Y(n_1433)
);

INVx8_ASAP7_75t_L g1434 ( 
.A(n_1262),
.Y(n_1434)
);

NOR2xp33_ASAP7_75t_L g1435 ( 
.A(n_1244),
.B(n_1111),
.Y(n_1435)
);

NAND2xp5_ASAP7_75t_SL g1436 ( 
.A(n_1271),
.B(n_831),
.Y(n_1436)
);

NOR2xp33_ASAP7_75t_L g1437 ( 
.A(n_1280),
.B(n_831),
.Y(n_1437)
);

INVx4_ASAP7_75t_L g1438 ( 
.A(n_1262),
.Y(n_1438)
);

NOR3xp33_ASAP7_75t_L g1439 ( 
.A(n_1315),
.B(n_833),
.C(n_780),
.Y(n_1439)
);

AOI22xp33_ASAP7_75t_L g1440 ( 
.A1(n_1272),
.A2(n_1200),
.B1(n_699),
.B2(n_702),
.Y(n_1440)
);

BUFx3_ASAP7_75t_L g1441 ( 
.A(n_1267),
.Y(n_1441)
);

NAND2xp5_ASAP7_75t_L g1442 ( 
.A(n_1348),
.B(n_1200),
.Y(n_1442)
);

AOI22xp33_ASAP7_75t_L g1443 ( 
.A1(n_1413),
.A2(n_702),
.B1(n_705),
.B2(n_643),
.Y(n_1443)
);

AND2x2_ASAP7_75t_L g1444 ( 
.A(n_1280),
.B(n_1286),
.Y(n_1444)
);

OAI22xp5_ASAP7_75t_L g1445 ( 
.A1(n_1348),
.A2(n_1201),
.B1(n_1198),
.B2(n_780),
.Y(n_1445)
);

AND2x6_ASAP7_75t_SL g1446 ( 
.A(n_1266),
.B(n_927),
.Y(n_1446)
);

INVx2_ASAP7_75t_L g1447 ( 
.A(n_1332),
.Y(n_1447)
);

NAND2xp5_ASAP7_75t_SL g1448 ( 
.A(n_1271),
.B(n_590),
.Y(n_1448)
);

OAI22xp33_ASAP7_75t_L g1449 ( 
.A1(n_1379),
.A2(n_591),
.B1(n_614),
.B2(n_595),
.Y(n_1449)
);

AOI22xp5_ASAP7_75t_L g1450 ( 
.A1(n_1420),
.A2(n_618),
.B1(n_619),
.B2(n_616),
.Y(n_1450)
);

NOR2xp33_ASAP7_75t_L g1451 ( 
.A(n_1232),
.B(n_620),
.Y(n_1451)
);

INVx2_ASAP7_75t_L g1452 ( 
.A(n_1341),
.Y(n_1452)
);

NAND2xp5_ASAP7_75t_L g1453 ( 
.A(n_1358),
.B(n_928),
.Y(n_1453)
);

INVx1_ASAP7_75t_L g1454 ( 
.A(n_1238),
.Y(n_1454)
);

NAND2xp5_ASAP7_75t_L g1455 ( 
.A(n_1283),
.B(n_931),
.Y(n_1455)
);

AND2x4_ASAP7_75t_L g1456 ( 
.A(n_1264),
.B(n_1168),
.Y(n_1456)
);

NOR2xp33_ASAP7_75t_L g1457 ( 
.A(n_1243),
.B(n_621),
.Y(n_1457)
);

NAND2xp5_ASAP7_75t_L g1458 ( 
.A(n_1395),
.B(n_932),
.Y(n_1458)
);

INVx2_ASAP7_75t_SL g1459 ( 
.A(n_1249),
.Y(n_1459)
);

BUFx3_ASAP7_75t_L g1460 ( 
.A(n_1259),
.Y(n_1460)
);

NAND2xp5_ASAP7_75t_SL g1461 ( 
.A(n_1269),
.B(n_1318),
.Y(n_1461)
);

NAND2xp5_ASAP7_75t_L g1462 ( 
.A(n_1373),
.B(n_623),
.Y(n_1462)
);

INVx1_ASAP7_75t_L g1463 ( 
.A(n_1241),
.Y(n_1463)
);

AND2x2_ASAP7_75t_L g1464 ( 
.A(n_1349),
.B(n_705),
.Y(n_1464)
);

NAND2xp5_ASAP7_75t_L g1465 ( 
.A(n_1391),
.B(n_625),
.Y(n_1465)
);

NAND2xp5_ASAP7_75t_L g1466 ( 
.A(n_1394),
.B(n_626),
.Y(n_1466)
);

AND2x6_ASAP7_75t_SL g1467 ( 
.A(n_1316),
.B(n_705),
.Y(n_1467)
);

AND2x6_ASAP7_75t_L g1468 ( 
.A(n_1254),
.B(n_661),
.Y(n_1468)
);

A2O1A1Ixp33_ASAP7_75t_L g1469 ( 
.A1(n_1260),
.A2(n_1371),
.B(n_1376),
.C(n_1256),
.Y(n_1469)
);

NAND2xp5_ASAP7_75t_SL g1470 ( 
.A(n_1269),
.B(n_628),
.Y(n_1470)
);

INVx1_ASAP7_75t_L g1471 ( 
.A(n_1242),
.Y(n_1471)
);

OR2x6_ASAP7_75t_L g1472 ( 
.A(n_1262),
.B(n_1168),
.Y(n_1472)
);

NOR2xp33_ASAP7_75t_L g1473 ( 
.A(n_1257),
.B(n_629),
.Y(n_1473)
);

AO21x1_ASAP7_75t_L g1474 ( 
.A1(n_1256),
.A2(n_1178),
.B(n_1175),
.Y(n_1474)
);

NOR2xp33_ASAP7_75t_L g1475 ( 
.A(n_1265),
.B(n_632),
.Y(n_1475)
);

AND2x4_ASAP7_75t_L g1476 ( 
.A(n_1264),
.B(n_1173),
.Y(n_1476)
);

NAND2xp5_ASAP7_75t_L g1477 ( 
.A(n_1255),
.B(n_1173),
.Y(n_1477)
);

AND2x6_ASAP7_75t_SL g1478 ( 
.A(n_1361),
.B(n_1318),
.Y(n_1478)
);

NAND2xp5_ASAP7_75t_L g1479 ( 
.A(n_1392),
.B(n_824),
.Y(n_1479)
);

NAND2xp5_ASAP7_75t_L g1480 ( 
.A(n_1325),
.B(n_825),
.Y(n_1480)
);

INVx1_ASAP7_75t_L g1481 ( 
.A(n_1245),
.Y(n_1481)
);

NAND3xp33_ASAP7_75t_SL g1482 ( 
.A(n_1289),
.B(n_646),
.C(n_644),
.Y(n_1482)
);

AOI21xp5_ASAP7_75t_L g1483 ( 
.A1(n_1301),
.A2(n_1178),
.B(n_1175),
.Y(n_1483)
);

INVx2_ASAP7_75t_L g1484 ( 
.A(n_1352),
.Y(n_1484)
);

INVx2_ASAP7_75t_L g1485 ( 
.A(n_1360),
.Y(n_1485)
);

OR2x6_ASAP7_75t_L g1486 ( 
.A(n_1408),
.B(n_775),
.Y(n_1486)
);

NOR2xp33_ASAP7_75t_L g1487 ( 
.A(n_1240),
.B(n_639),
.Y(n_1487)
);

NAND2xp5_ASAP7_75t_L g1488 ( 
.A(n_1334),
.B(n_649),
.Y(n_1488)
);

BUFx6f_ASAP7_75t_L g1489 ( 
.A(n_1431),
.Y(n_1489)
);

NAND2xp5_ASAP7_75t_SL g1490 ( 
.A(n_1322),
.B(n_1354),
.Y(n_1490)
);

NOR2xp33_ASAP7_75t_L g1491 ( 
.A(n_1386),
.B(n_651),
.Y(n_1491)
);

NAND3xp33_ASAP7_75t_L g1492 ( 
.A(n_1234),
.B(n_719),
.C(n_715),
.Y(n_1492)
);

NOR2x1p5_ASAP7_75t_L g1493 ( 
.A(n_1261),
.B(n_657),
.Y(n_1493)
);

NAND2xp5_ASAP7_75t_SL g1494 ( 
.A(n_1322),
.B(n_659),
.Y(n_1494)
);

INVx1_ASAP7_75t_L g1495 ( 
.A(n_1253),
.Y(n_1495)
);

INVx1_ASAP7_75t_L g1496 ( 
.A(n_1263),
.Y(n_1496)
);

INVx1_ASAP7_75t_L g1497 ( 
.A(n_1268),
.Y(n_1497)
);

AOI22xp33_ASAP7_75t_L g1498 ( 
.A1(n_1402),
.A2(n_734),
.B1(n_793),
.B2(n_717),
.Y(n_1498)
);

INVx2_ASAP7_75t_SL g1499 ( 
.A(n_1249),
.Y(n_1499)
);

NAND2xp5_ASAP7_75t_L g1500 ( 
.A(n_1388),
.B(n_660),
.Y(n_1500)
);

NAND2xp5_ASAP7_75t_L g1501 ( 
.A(n_1388),
.B(n_662),
.Y(n_1501)
);

OAI21xp5_ASAP7_75t_L g1502 ( 
.A1(n_1235),
.A2(n_785),
.B(n_775),
.Y(n_1502)
);

INVx1_ASAP7_75t_L g1503 ( 
.A(n_1270),
.Y(n_1503)
);

NAND2xp5_ASAP7_75t_SL g1504 ( 
.A(n_1354),
.B(n_1314),
.Y(n_1504)
);

INVx2_ASAP7_75t_L g1505 ( 
.A(n_1382),
.Y(n_1505)
);

NAND2xp5_ASAP7_75t_L g1506 ( 
.A(n_1343),
.B(n_665),
.Y(n_1506)
);

AND2x4_ASAP7_75t_L g1507 ( 
.A(n_1293),
.B(n_785),
.Y(n_1507)
);

INVx1_ASAP7_75t_L g1508 ( 
.A(n_1279),
.Y(n_1508)
);

NOR3xp33_ASAP7_75t_L g1509 ( 
.A(n_1404),
.B(n_812),
.C(n_669),
.Y(n_1509)
);

NAND2xp5_ASAP7_75t_L g1510 ( 
.A(n_1396),
.B(n_821),
.Y(n_1510)
);

INVx2_ASAP7_75t_L g1511 ( 
.A(n_1233),
.Y(n_1511)
);

NAND2xp5_ASAP7_75t_L g1512 ( 
.A(n_1255),
.B(n_1417),
.Y(n_1512)
);

OAI21xp5_ASAP7_75t_L g1513 ( 
.A1(n_1235),
.A2(n_812),
.B(n_674),
.Y(n_1513)
);

NAND2xp5_ASAP7_75t_L g1514 ( 
.A(n_1239),
.B(n_666),
.Y(n_1514)
);

NAND2xp5_ASAP7_75t_L g1515 ( 
.A(n_1239),
.B(n_675),
.Y(n_1515)
);

NAND2xp5_ASAP7_75t_L g1516 ( 
.A(n_1410),
.B(n_679),
.Y(n_1516)
);

BUFx6f_ASAP7_75t_L g1517 ( 
.A(n_1431),
.Y(n_1517)
);

INVx2_ASAP7_75t_L g1518 ( 
.A(n_1236),
.Y(n_1518)
);

NAND2xp5_ASAP7_75t_L g1519 ( 
.A(n_1396),
.B(n_681),
.Y(n_1519)
);

AOI22xp33_ASAP7_75t_L g1520 ( 
.A1(n_1379),
.A2(n_734),
.B1(n_793),
.B2(n_717),
.Y(n_1520)
);

BUFx3_ASAP7_75t_L g1521 ( 
.A(n_1296),
.Y(n_1521)
);

NAND2xp5_ASAP7_75t_SL g1522 ( 
.A(n_1342),
.B(n_682),
.Y(n_1522)
);

OAI221xp5_ASAP7_75t_L g1523 ( 
.A1(n_1404),
.A2(n_685),
.B1(n_686),
.B2(n_684),
.C(n_683),
.Y(n_1523)
);

NAND2xp5_ASAP7_75t_L g1524 ( 
.A(n_1416),
.B(n_688),
.Y(n_1524)
);

INVx1_ASAP7_75t_L g1525 ( 
.A(n_1281),
.Y(n_1525)
);

NAND2xp5_ASAP7_75t_SL g1526 ( 
.A(n_1431),
.B(n_689),
.Y(n_1526)
);

INVx2_ASAP7_75t_L g1527 ( 
.A(n_1246),
.Y(n_1527)
);

NAND2xp5_ASAP7_75t_L g1528 ( 
.A(n_1356),
.B(n_827),
.Y(n_1528)
);

NAND2xp5_ASAP7_75t_L g1529 ( 
.A(n_1275),
.B(n_690),
.Y(n_1529)
);

NAND2xp5_ASAP7_75t_SL g1530 ( 
.A(n_1366),
.B(n_691),
.Y(n_1530)
);

NAND2xp5_ASAP7_75t_SL g1531 ( 
.A(n_1366),
.B(n_694),
.Y(n_1531)
);

INVx2_ASAP7_75t_L g1532 ( 
.A(n_1247),
.Y(n_1532)
);

INVx2_ASAP7_75t_L g1533 ( 
.A(n_1251),
.Y(n_1533)
);

OR2x6_ASAP7_75t_SL g1534 ( 
.A(n_1295),
.B(n_697),
.Y(n_1534)
);

OAI22xp5_ASAP7_75t_SL g1535 ( 
.A1(n_1361),
.A2(n_698),
.B1(n_710),
.B2(n_701),
.Y(n_1535)
);

NAND2xp5_ASAP7_75t_SL g1536 ( 
.A(n_1363),
.B(n_716),
.Y(n_1536)
);

OAI21xp5_ASAP7_75t_L g1537 ( 
.A1(n_1415),
.A2(n_1305),
.B(n_1301),
.Y(n_1537)
);

NAND2xp5_ASAP7_75t_L g1538 ( 
.A(n_1303),
.B(n_720),
.Y(n_1538)
);

INVx2_ASAP7_75t_L g1539 ( 
.A(n_1252),
.Y(n_1539)
);

AND2x2_ASAP7_75t_L g1540 ( 
.A(n_1237),
.B(n_717),
.Y(n_1540)
);

NAND2xp5_ASAP7_75t_L g1541 ( 
.A(n_1308),
.B(n_722),
.Y(n_1541)
);

AOI22xp5_ASAP7_75t_L g1542 ( 
.A1(n_1411),
.A2(n_727),
.B1(n_728),
.B2(n_726),
.Y(n_1542)
);

AND2x4_ASAP7_75t_L g1543 ( 
.A(n_1293),
.B(n_715),
.Y(n_1543)
);

NAND2xp5_ASAP7_75t_L g1544 ( 
.A(n_1321),
.B(n_828),
.Y(n_1544)
);

NAND2xp5_ASAP7_75t_L g1545 ( 
.A(n_1278),
.B(n_730),
.Y(n_1545)
);

INVx1_ASAP7_75t_L g1546 ( 
.A(n_1285),
.Y(n_1546)
);

INVx1_ASAP7_75t_L g1547 ( 
.A(n_1397),
.Y(n_1547)
);

AOI22xp33_ASAP7_75t_L g1548 ( 
.A1(n_1336),
.A2(n_818),
.B1(n_734),
.B2(n_741),
.Y(n_1548)
);

NOR2xp33_ASAP7_75t_L g1549 ( 
.A(n_1385),
.B(n_731),
.Y(n_1549)
);

INVx3_ASAP7_75t_L g1550 ( 
.A(n_1364),
.Y(n_1550)
);

NAND2xp5_ASAP7_75t_SL g1551 ( 
.A(n_1367),
.B(n_745),
.Y(n_1551)
);

INVx2_ASAP7_75t_L g1552 ( 
.A(n_1273),
.Y(n_1552)
);

BUFx8_ASAP7_75t_L g1553 ( 
.A(n_1313),
.Y(n_1553)
);

NAND2xp5_ASAP7_75t_SL g1554 ( 
.A(n_1311),
.B(n_746),
.Y(n_1554)
);

AOI22xp5_ASAP7_75t_L g1555 ( 
.A1(n_1336),
.A2(n_749),
.B1(n_753),
.B2(n_748),
.Y(n_1555)
);

NAND2xp5_ASAP7_75t_L g1556 ( 
.A(n_1305),
.B(n_759),
.Y(n_1556)
);

AOI21xp5_ASAP7_75t_L g1557 ( 
.A1(n_1320),
.A2(n_596),
.B(n_589),
.Y(n_1557)
);

AOI22xp33_ASAP7_75t_L g1558 ( 
.A1(n_1350),
.A2(n_818),
.B1(n_764),
.B2(n_765),
.Y(n_1558)
);

AND2x2_ASAP7_75t_L g1559 ( 
.A(n_1346),
.B(n_818),
.Y(n_1559)
);

INVx4_ASAP7_75t_L g1560 ( 
.A(n_1299),
.Y(n_1560)
);

INVx2_ASAP7_75t_L g1561 ( 
.A(n_1277),
.Y(n_1561)
);

NAND2xp5_ASAP7_75t_SL g1562 ( 
.A(n_1350),
.B(n_761),
.Y(n_1562)
);

NAND2xp5_ASAP7_75t_L g1563 ( 
.A(n_1374),
.B(n_810),
.Y(n_1563)
);

NAND2xp5_ASAP7_75t_L g1564 ( 
.A(n_1374),
.B(n_832),
.Y(n_1564)
);

NAND3xp33_ASAP7_75t_L g1565 ( 
.A(n_1426),
.B(n_755),
.C(n_719),
.Y(n_1565)
);

NAND2xp5_ASAP7_75t_SL g1566 ( 
.A(n_1299),
.B(n_767),
.Y(n_1566)
);

NAND2xp5_ASAP7_75t_L g1567 ( 
.A(n_1399),
.B(n_1400),
.Y(n_1567)
);

NAND2xp5_ASAP7_75t_L g1568 ( 
.A(n_1260),
.B(n_768),
.Y(n_1568)
);

AND2x4_ASAP7_75t_L g1569 ( 
.A(n_1329),
.B(n_755),
.Y(n_1569)
);

NOR2xp33_ASAP7_75t_L g1570 ( 
.A(n_1361),
.B(n_770),
.Y(n_1570)
);

NAND2xp33_ASAP7_75t_L g1571 ( 
.A(n_1274),
.B(n_771),
.Y(n_1571)
);

NAND2xp5_ASAP7_75t_L g1572 ( 
.A(n_1290),
.B(n_772),
.Y(n_1572)
);

NOR2xp33_ASAP7_75t_L g1573 ( 
.A(n_1298),
.B(n_777),
.Y(n_1573)
);

INVx2_ASAP7_75t_L g1574 ( 
.A(n_1284),
.Y(n_1574)
);

NAND2xp5_ASAP7_75t_L g1575 ( 
.A(n_1290),
.B(n_778),
.Y(n_1575)
);

NAND2xp5_ASAP7_75t_SL g1576 ( 
.A(n_1357),
.B(n_782),
.Y(n_1576)
);

INVx3_ASAP7_75t_L g1577 ( 
.A(n_1364),
.Y(n_1577)
);

INVx1_ASAP7_75t_L g1578 ( 
.A(n_1390),
.Y(n_1578)
);

AOI21xp5_ASAP7_75t_L g1579 ( 
.A1(n_1320),
.A2(n_613),
.B(n_597),
.Y(n_1579)
);

NAND2xp5_ASAP7_75t_L g1580 ( 
.A(n_1306),
.B(n_1310),
.Y(n_1580)
);

NAND2xp5_ASAP7_75t_L g1581 ( 
.A(n_1306),
.B(n_784),
.Y(n_1581)
);

NAND2xp5_ASAP7_75t_L g1582 ( 
.A(n_1310),
.B(n_786),
.Y(n_1582)
);

INVx1_ASAP7_75t_L g1583 ( 
.A(n_1401),
.Y(n_1583)
);

AND2x2_ASAP7_75t_L g1584 ( 
.A(n_1359),
.B(n_1250),
.Y(n_1584)
);

NAND2xp5_ASAP7_75t_L g1585 ( 
.A(n_1418),
.B(n_804),
.Y(n_1585)
);

INVx2_ASAP7_75t_L g1586 ( 
.A(n_1292),
.Y(n_1586)
);

NAND2xp5_ASAP7_75t_SL g1587 ( 
.A(n_1357),
.B(n_789),
.Y(n_1587)
);

AND2x6_ASAP7_75t_SL g1588 ( 
.A(n_1418),
.B(n_791),
.Y(n_1588)
);

NAND2xp5_ASAP7_75t_SL g1589 ( 
.A(n_1380),
.B(n_792),
.Y(n_1589)
);

AOI22xp33_ASAP7_75t_L g1590 ( 
.A1(n_1375),
.A2(n_805),
.B1(n_809),
.B2(n_796),
.Y(n_1590)
);

AOI22xp5_ASAP7_75t_L g1591 ( 
.A1(n_1427),
.A2(n_1337),
.B1(n_1327),
.B2(n_1287),
.Y(n_1591)
);

INVx1_ASAP7_75t_L g1592 ( 
.A(n_1405),
.Y(n_1592)
);

NOR2xp33_ASAP7_75t_L g1593 ( 
.A(n_1421),
.B(n_615),
.Y(n_1593)
);

NAND2xp5_ASAP7_75t_L g1594 ( 
.A(n_1324),
.B(n_755),
.Y(n_1594)
);

AOI22xp5_ASAP7_75t_L g1595 ( 
.A1(n_1327),
.A2(n_653),
.B1(n_658),
.B2(n_642),
.Y(n_1595)
);

NOR2x2_ASAP7_75t_L g1596 ( 
.A(n_1419),
.B(n_0),
.Y(n_1596)
);

INVx2_ASAP7_75t_L g1597 ( 
.A(n_1330),
.Y(n_1597)
);

AOI22xp5_ASAP7_75t_L g1598 ( 
.A1(n_1337),
.A2(n_709),
.B1(n_714),
.B2(n_704),
.Y(n_1598)
);

NOR2xp33_ASAP7_75t_L g1599 ( 
.A(n_1424),
.B(n_738),
.Y(n_1599)
);

AND2x6_ASAP7_75t_L g1600 ( 
.A(n_1254),
.B(n_750),
.Y(n_1600)
);

NAND2xp5_ASAP7_75t_L g1601 ( 
.A(n_1331),
.B(n_755),
.Y(n_1601)
);

INVx2_ASAP7_75t_L g1602 ( 
.A(n_1338),
.Y(n_1602)
);

NAND2xp5_ASAP7_75t_SL g1603 ( 
.A(n_1380),
.B(n_800),
.Y(n_1603)
);

INVx2_ASAP7_75t_L g1604 ( 
.A(n_1344),
.Y(n_1604)
);

NAND2xp5_ASAP7_75t_L g1605 ( 
.A(n_1345),
.B(n_816),
.Y(n_1605)
);

AOI22xp5_ASAP7_75t_L g1606 ( 
.A1(n_1274),
.A2(n_744),
.B1(n_747),
.B2(n_743),
.Y(n_1606)
);

INVx2_ASAP7_75t_L g1607 ( 
.A(n_1351),
.Y(n_1607)
);

AOI22xp5_ASAP7_75t_L g1608 ( 
.A1(n_1274),
.A2(n_766),
.B1(n_794),
.B2(n_752),
.Y(n_1608)
);

AND2x6_ASAP7_75t_SL g1609 ( 
.A(n_1429),
.B(n_1),
.Y(n_1609)
);

NOR2xp33_ASAP7_75t_L g1610 ( 
.A(n_1428),
.B(n_811),
.Y(n_1610)
);

AND2x6_ASAP7_75t_SL g1611 ( 
.A(n_1429),
.B(n_1),
.Y(n_1611)
);

BUFx6f_ASAP7_75t_L g1612 ( 
.A(n_1291),
.Y(n_1612)
);

NAND2xp5_ASAP7_75t_L g1613 ( 
.A(n_1353),
.B(n_816),
.Y(n_1613)
);

INVx2_ASAP7_75t_L g1614 ( 
.A(n_1355),
.Y(n_1614)
);

NAND2xp5_ASAP7_75t_L g1615 ( 
.A(n_1372),
.B(n_1378),
.Y(n_1615)
);

NAND2xp5_ASAP7_75t_SL g1616 ( 
.A(n_1291),
.B(n_820),
.Y(n_1616)
);

BUFx8_ASAP7_75t_L g1617 ( 
.A(n_1291),
.Y(n_1617)
);

INVx1_ASAP7_75t_L g1618 ( 
.A(n_1387),
.Y(n_1618)
);

INVx2_ASAP7_75t_L g1619 ( 
.A(n_1370),
.Y(n_1619)
);

NAND2xp5_ASAP7_75t_SL g1620 ( 
.A(n_1297),
.B(n_816),
.Y(n_1620)
);

INVx1_ASAP7_75t_L g1621 ( 
.A(n_1370),
.Y(n_1621)
);

NOR2xp33_ASAP7_75t_L g1622 ( 
.A(n_1384),
.B(n_2),
.Y(n_1622)
);

NAND2xp5_ASAP7_75t_L g1623 ( 
.A(n_1362),
.B(n_1422),
.Y(n_1623)
);

NAND2xp5_ASAP7_75t_L g1624 ( 
.A(n_1362),
.B(n_819),
.Y(n_1624)
);

AOI22xp33_ASAP7_75t_L g1625 ( 
.A1(n_1375),
.A2(n_819),
.B1(n_952),
.B2(n_951),
.Y(n_1625)
);

O2A1O1Ixp5_ASAP7_75t_L g1626 ( 
.A1(n_1328),
.A2(n_819),
.B(n_4),
.C(n_2),
.Y(n_1626)
);

AND2x2_ASAP7_75t_L g1627 ( 
.A(n_1406),
.B(n_3),
.Y(n_1627)
);

BUFx3_ASAP7_75t_L g1628 ( 
.A(n_1432),
.Y(n_1628)
);

NAND2xp5_ASAP7_75t_L g1629 ( 
.A(n_1422),
.B(n_3),
.Y(n_1629)
);

AOI22xp33_ASAP7_75t_L g1630 ( 
.A1(n_1377),
.A2(n_952),
.B1(n_958),
.B2(n_951),
.Y(n_1630)
);

AND2x2_ASAP7_75t_L g1631 ( 
.A(n_1407),
.B(n_5),
.Y(n_1631)
);

INVx5_ASAP7_75t_L g1632 ( 
.A(n_1274),
.Y(n_1632)
);

BUFx3_ASAP7_75t_L g1633 ( 
.A(n_1297),
.Y(n_1633)
);

O2A1O1Ixp5_ASAP7_75t_L g1634 ( 
.A1(n_1258),
.A2(n_7),
.B(n_5),
.C(n_6),
.Y(n_1634)
);

NAND2xp5_ASAP7_75t_L g1635 ( 
.A(n_1407),
.B(n_1423),
.Y(n_1635)
);

INVx2_ASAP7_75t_L g1636 ( 
.A(n_1365),
.Y(n_1636)
);

INVx2_ASAP7_75t_SL g1637 ( 
.A(n_1297),
.Y(n_1637)
);

INVx2_ASAP7_75t_SL g1638 ( 
.A(n_1300),
.Y(n_1638)
);

AND2x2_ASAP7_75t_SL g1639 ( 
.A(n_1430),
.B(n_7),
.Y(n_1639)
);

OR2x6_ASAP7_75t_L g1640 ( 
.A(n_1486),
.B(n_1408),
.Y(n_1640)
);

NOR2xp33_ASAP7_75t_L g1641 ( 
.A(n_1475),
.B(n_1398),
.Y(n_1641)
);

NAND2xp5_ASAP7_75t_L g1642 ( 
.A(n_1444),
.B(n_1398),
.Y(n_1642)
);

NAND2xp5_ASAP7_75t_L g1643 ( 
.A(n_1464),
.B(n_1403),
.Y(n_1643)
);

NAND2xp5_ASAP7_75t_SL g1644 ( 
.A(n_1433),
.B(n_1300),
.Y(n_1644)
);

INVx1_ASAP7_75t_L g1645 ( 
.A(n_1508),
.Y(n_1645)
);

INVx2_ASAP7_75t_L g1646 ( 
.A(n_1597),
.Y(n_1646)
);

NAND2xp5_ASAP7_75t_L g1647 ( 
.A(n_1512),
.B(n_1403),
.Y(n_1647)
);

INVx2_ASAP7_75t_L g1648 ( 
.A(n_1602),
.Y(n_1648)
);

INVx2_ASAP7_75t_L g1649 ( 
.A(n_1604),
.Y(n_1649)
);

INVx1_ASAP7_75t_L g1650 ( 
.A(n_1525),
.Y(n_1650)
);

AND2x4_ASAP7_75t_L g1651 ( 
.A(n_1459),
.B(n_1381),
.Y(n_1651)
);

INVx1_ASAP7_75t_L g1652 ( 
.A(n_1546),
.Y(n_1652)
);

INVx5_ASAP7_75t_L g1653 ( 
.A(n_1434),
.Y(n_1653)
);

INVx3_ASAP7_75t_L g1654 ( 
.A(n_1434),
.Y(n_1654)
);

OR2x6_ASAP7_75t_L g1655 ( 
.A(n_1486),
.B(n_1408),
.Y(n_1655)
);

BUFx6f_ASAP7_75t_L g1656 ( 
.A(n_1434),
.Y(n_1656)
);

NAND2xp5_ASAP7_75t_L g1657 ( 
.A(n_1512),
.B(n_1319),
.Y(n_1657)
);

INVx1_ASAP7_75t_L g1658 ( 
.A(n_1454),
.Y(n_1658)
);

INVx1_ASAP7_75t_L g1659 ( 
.A(n_1463),
.Y(n_1659)
);

INVx1_ASAP7_75t_L g1660 ( 
.A(n_1471),
.Y(n_1660)
);

INVx2_ASAP7_75t_L g1661 ( 
.A(n_1607),
.Y(n_1661)
);

AND2x2_ASAP7_75t_L g1662 ( 
.A(n_1540),
.B(n_6),
.Y(n_1662)
);

INVx1_ASAP7_75t_L g1663 ( 
.A(n_1481),
.Y(n_1663)
);

BUFx3_ASAP7_75t_L g1664 ( 
.A(n_1521),
.Y(n_1664)
);

NAND2xp5_ASAP7_75t_L g1665 ( 
.A(n_1455),
.B(n_1300),
.Y(n_1665)
);

INVx2_ASAP7_75t_L g1666 ( 
.A(n_1614),
.Y(n_1666)
);

INVx2_ASAP7_75t_L g1667 ( 
.A(n_1447),
.Y(n_1667)
);

NAND2xp5_ASAP7_75t_SL g1668 ( 
.A(n_1435),
.B(n_1307),
.Y(n_1668)
);

INVx1_ASAP7_75t_L g1669 ( 
.A(n_1495),
.Y(n_1669)
);

NAND2xp5_ASAP7_75t_SL g1670 ( 
.A(n_1639),
.B(n_1307),
.Y(n_1670)
);

NOR2x1p5_ASAP7_75t_L g1671 ( 
.A(n_1441),
.B(n_1304),
.Y(n_1671)
);

NAND2xp5_ASAP7_75t_SL g1672 ( 
.A(n_1489),
.B(n_1307),
.Y(n_1672)
);

INVx1_ASAP7_75t_L g1673 ( 
.A(n_1496),
.Y(n_1673)
);

AND2x4_ASAP7_75t_SL g1674 ( 
.A(n_1438),
.B(n_1319),
.Y(n_1674)
);

NAND2xp5_ASAP7_75t_L g1675 ( 
.A(n_1453),
.B(n_1319),
.Y(n_1675)
);

NAND2xp5_ASAP7_75t_SL g1676 ( 
.A(n_1489),
.B(n_1335),
.Y(n_1676)
);

NOR2xp33_ASAP7_75t_L g1677 ( 
.A(n_1491),
.B(n_1335),
.Y(n_1677)
);

AND2x6_ASAP7_75t_SL g1678 ( 
.A(n_1437),
.B(n_1365),
.Y(n_1678)
);

BUFx3_ASAP7_75t_L g1679 ( 
.A(n_1460),
.Y(n_1679)
);

NAND2xp5_ASAP7_75t_SL g1680 ( 
.A(n_1489),
.B(n_1335),
.Y(n_1680)
);

BUFx6f_ASAP7_75t_L g1681 ( 
.A(n_1517),
.Y(n_1681)
);

INVx2_ASAP7_75t_L g1682 ( 
.A(n_1452),
.Y(n_1682)
);

NAND2xp5_ASAP7_75t_L g1683 ( 
.A(n_1488),
.B(n_1339),
.Y(n_1683)
);

AND2x4_ASAP7_75t_L g1684 ( 
.A(n_1499),
.B(n_1381),
.Y(n_1684)
);

BUFx6f_ASAP7_75t_L g1685 ( 
.A(n_1517),
.Y(n_1685)
);

BUFx6f_ASAP7_75t_L g1686 ( 
.A(n_1517),
.Y(n_1686)
);

INVx1_ASAP7_75t_L g1687 ( 
.A(n_1497),
.Y(n_1687)
);

NOR2xp67_ASAP7_75t_L g1688 ( 
.A(n_1632),
.B(n_1369),
.Y(n_1688)
);

OAI21xp5_ASAP7_75t_L g1689 ( 
.A1(n_1469),
.A2(n_1414),
.B(n_1377),
.Y(n_1689)
);

OR2x6_ASAP7_75t_L g1690 ( 
.A(n_1486),
.B(n_1369),
.Y(n_1690)
);

INVx4_ASAP7_75t_L g1691 ( 
.A(n_1438),
.Y(n_1691)
);

AOI22xp5_ASAP7_75t_L g1692 ( 
.A1(n_1449),
.A2(n_1287),
.B1(n_1288),
.B2(n_1294),
.Y(n_1692)
);

INVx2_ASAP7_75t_L g1693 ( 
.A(n_1484),
.Y(n_1693)
);

NOR2xp33_ASAP7_75t_L g1694 ( 
.A(n_1446),
.B(n_1339),
.Y(n_1694)
);

INVx1_ASAP7_75t_L g1695 ( 
.A(n_1503),
.Y(n_1695)
);

NAND2xp5_ASAP7_75t_L g1696 ( 
.A(n_1458),
.B(n_1339),
.Y(n_1696)
);

INVx2_ASAP7_75t_L g1697 ( 
.A(n_1485),
.Y(n_1697)
);

AOI22xp33_ASAP7_75t_L g1698 ( 
.A1(n_1627),
.A2(n_1312),
.B1(n_1294),
.B2(n_1287),
.Y(n_1698)
);

INVx1_ASAP7_75t_L g1699 ( 
.A(n_1547),
.Y(n_1699)
);

NAND2xp5_ASAP7_75t_L g1700 ( 
.A(n_1480),
.B(n_1567),
.Y(n_1700)
);

BUFx2_ASAP7_75t_L g1701 ( 
.A(n_1617),
.Y(n_1701)
);

AOI22xp33_ASAP7_75t_L g1702 ( 
.A1(n_1530),
.A2(n_1294),
.B1(n_1287),
.B2(n_1288),
.Y(n_1702)
);

CKINVDCx11_ASAP7_75t_R g1703 ( 
.A(n_1534),
.Y(n_1703)
);

AND2x6_ASAP7_75t_SL g1704 ( 
.A(n_1573),
.B(n_1368),
.Y(n_1704)
);

INVx2_ASAP7_75t_L g1705 ( 
.A(n_1505),
.Y(n_1705)
);

AOI22xp33_ASAP7_75t_L g1706 ( 
.A1(n_1531),
.A2(n_1294),
.B1(n_1288),
.B2(n_1393),
.Y(n_1706)
);

INVx1_ASAP7_75t_L g1707 ( 
.A(n_1578),
.Y(n_1707)
);

INVx1_ASAP7_75t_L g1708 ( 
.A(n_1583),
.Y(n_1708)
);

AOI22xp33_ASAP7_75t_L g1709 ( 
.A1(n_1520),
.A2(n_1288),
.B1(n_1393),
.B2(n_1309),
.Y(n_1709)
);

INVx1_ASAP7_75t_L g1710 ( 
.A(n_1592),
.Y(n_1710)
);

CKINVDCx5p33_ASAP7_75t_R g1711 ( 
.A(n_1553),
.Y(n_1711)
);

NAND2xp5_ASAP7_75t_SL g1712 ( 
.A(n_1632),
.B(n_1340),
.Y(n_1712)
);

INVx2_ASAP7_75t_SL g1713 ( 
.A(n_1553),
.Y(n_1713)
);

INVx1_ASAP7_75t_L g1714 ( 
.A(n_1618),
.Y(n_1714)
);

NAND2xp5_ASAP7_75t_SL g1715 ( 
.A(n_1632),
.B(n_1340),
.Y(n_1715)
);

BUFx2_ASAP7_75t_L g1716 ( 
.A(n_1617),
.Y(n_1716)
);

AND2x4_ASAP7_75t_L g1717 ( 
.A(n_1580),
.B(n_1340),
.Y(n_1717)
);

INVx1_ASAP7_75t_L g1718 ( 
.A(n_1511),
.Y(n_1718)
);

NAND2xp5_ASAP7_75t_L g1719 ( 
.A(n_1556),
.B(n_1462),
.Y(n_1719)
);

INVx1_ASAP7_75t_L g1720 ( 
.A(n_1518),
.Y(n_1720)
);

INVx2_ASAP7_75t_L g1721 ( 
.A(n_1527),
.Y(n_1721)
);

HB1xp67_ASAP7_75t_L g1722 ( 
.A(n_1631),
.Y(n_1722)
);

BUFx6f_ASAP7_75t_L g1723 ( 
.A(n_1612),
.Y(n_1723)
);

BUFx2_ASAP7_75t_L g1724 ( 
.A(n_1628),
.Y(n_1724)
);

HB1xp67_ASAP7_75t_L g1725 ( 
.A(n_1461),
.Y(n_1725)
);

INVx2_ASAP7_75t_L g1726 ( 
.A(n_1532),
.Y(n_1726)
);

INVx3_ASAP7_75t_L g1727 ( 
.A(n_1612),
.Y(n_1727)
);

INVx3_ASAP7_75t_L g1728 ( 
.A(n_1612),
.Y(n_1728)
);

INVx1_ASAP7_75t_L g1729 ( 
.A(n_1533),
.Y(n_1729)
);

INVx1_ASAP7_75t_L g1730 ( 
.A(n_1539),
.Y(n_1730)
);

NOR2xp33_ASAP7_75t_L g1731 ( 
.A(n_1490),
.B(n_1383),
.Y(n_1731)
);

INVx1_ASAP7_75t_L g1732 ( 
.A(n_1552),
.Y(n_1732)
);

INVx2_ASAP7_75t_L g1733 ( 
.A(n_1561),
.Y(n_1733)
);

INVx1_ASAP7_75t_L g1734 ( 
.A(n_1574),
.Y(n_1734)
);

BUFx2_ASAP7_75t_L g1735 ( 
.A(n_1584),
.Y(n_1735)
);

BUFx4f_ASAP7_75t_L g1736 ( 
.A(n_1472),
.Y(n_1736)
);

NOR2xp67_ASAP7_75t_L g1737 ( 
.A(n_1550),
.B(n_1304),
.Y(n_1737)
);

INVx2_ASAP7_75t_L g1738 ( 
.A(n_1586),
.Y(n_1738)
);

INVx2_ASAP7_75t_L g1739 ( 
.A(n_1636),
.Y(n_1739)
);

INVx1_ASAP7_75t_L g1740 ( 
.A(n_1615),
.Y(n_1740)
);

HB1xp67_ASAP7_75t_L g1741 ( 
.A(n_1633),
.Y(n_1741)
);

AND2x2_ASAP7_75t_L g1742 ( 
.A(n_1451),
.B(n_8),
.Y(n_1742)
);

NAND2xp5_ASAP7_75t_SL g1743 ( 
.A(n_1535),
.B(n_1383),
.Y(n_1743)
);

NAND2xp5_ASAP7_75t_L g1744 ( 
.A(n_1556),
.B(n_1383),
.Y(n_1744)
);

INVx2_ASAP7_75t_L g1745 ( 
.A(n_1619),
.Y(n_1745)
);

AND2x4_ASAP7_75t_L g1746 ( 
.A(n_1560),
.B(n_1425),
.Y(n_1746)
);

NAND2xp5_ASAP7_75t_L g1747 ( 
.A(n_1621),
.B(n_1537),
.Y(n_1747)
);

INVx2_ASAP7_75t_SL g1748 ( 
.A(n_1493),
.Y(n_1748)
);

OAI22xp5_ASAP7_75t_SL g1749 ( 
.A1(n_1440),
.A2(n_1323),
.B1(n_1326),
.B2(n_1317),
.Y(n_1749)
);

INVx1_ASAP7_75t_L g1750 ( 
.A(n_1594),
.Y(n_1750)
);

NOR2xp33_ASAP7_75t_L g1751 ( 
.A(n_1549),
.B(n_1504),
.Y(n_1751)
);

NAND2xp5_ASAP7_75t_SL g1752 ( 
.A(n_1591),
.B(n_1456),
.Y(n_1752)
);

INVx2_ASAP7_75t_L g1753 ( 
.A(n_1635),
.Y(n_1753)
);

NOR2xp33_ASAP7_75t_L g1754 ( 
.A(n_1562),
.B(n_1425),
.Y(n_1754)
);

NOR2xp67_ASAP7_75t_L g1755 ( 
.A(n_1550),
.B(n_1317),
.Y(n_1755)
);

OR2x2_ASAP7_75t_L g1756 ( 
.A(n_1465),
.B(n_1368),
.Y(n_1756)
);

INVx2_ASAP7_75t_L g1757 ( 
.A(n_1624),
.Y(n_1757)
);

BUFx2_ASAP7_75t_L g1758 ( 
.A(n_1560),
.Y(n_1758)
);

BUFx4f_ASAP7_75t_L g1759 ( 
.A(n_1472),
.Y(n_1759)
);

BUFx6f_ASAP7_75t_L g1760 ( 
.A(n_1472),
.Y(n_1760)
);

INVx2_ASAP7_75t_L g1761 ( 
.A(n_1624),
.Y(n_1761)
);

AND2x6_ASAP7_75t_L g1762 ( 
.A(n_1456),
.B(n_1323),
.Y(n_1762)
);

INVx1_ASAP7_75t_L g1763 ( 
.A(n_1629),
.Y(n_1763)
);

INVx2_ASAP7_75t_L g1764 ( 
.A(n_1601),
.Y(n_1764)
);

INVx1_ASAP7_75t_L g1765 ( 
.A(n_1629),
.Y(n_1765)
);

NAND2xp5_ASAP7_75t_L g1766 ( 
.A(n_1487),
.B(n_1425),
.Y(n_1766)
);

INVx1_ASAP7_75t_L g1767 ( 
.A(n_1516),
.Y(n_1767)
);

INVx2_ASAP7_75t_L g1768 ( 
.A(n_1605),
.Y(n_1768)
);

INVx1_ASAP7_75t_L g1769 ( 
.A(n_1516),
.Y(n_1769)
);

INVx2_ASAP7_75t_L g1770 ( 
.A(n_1613),
.Y(n_1770)
);

BUFx2_ASAP7_75t_L g1771 ( 
.A(n_1637),
.Y(n_1771)
);

OR2x6_ASAP7_75t_L g1772 ( 
.A(n_1476),
.B(n_1276),
.Y(n_1772)
);

NAND2xp5_ASAP7_75t_L g1773 ( 
.A(n_1473),
.B(n_1326),
.Y(n_1773)
);

INVx3_ASAP7_75t_L g1774 ( 
.A(n_1577),
.Y(n_1774)
);

AOI22xp33_ASAP7_75t_L g1775 ( 
.A1(n_1498),
.A2(n_1309),
.B1(n_1302),
.B2(n_1389),
.Y(n_1775)
);

BUFx4f_ASAP7_75t_L g1776 ( 
.A(n_1468),
.Y(n_1776)
);

NAND2xp5_ASAP7_75t_L g1777 ( 
.A(n_1457),
.B(n_1333),
.Y(n_1777)
);

INVx3_ASAP7_75t_L g1778 ( 
.A(n_1577),
.Y(n_1778)
);

NAND2xp5_ASAP7_75t_L g1779 ( 
.A(n_1559),
.B(n_1333),
.Y(n_1779)
);

NAND2xp5_ASAP7_75t_L g1780 ( 
.A(n_1537),
.B(n_1302),
.Y(n_1780)
);

BUFx6f_ASAP7_75t_L g1781 ( 
.A(n_1478),
.Y(n_1781)
);

INVx1_ASAP7_75t_L g1782 ( 
.A(n_1524),
.Y(n_1782)
);

INVx2_ASAP7_75t_L g1783 ( 
.A(n_1524),
.Y(n_1783)
);

INVx1_ASAP7_75t_L g1784 ( 
.A(n_1529),
.Y(n_1784)
);

NAND2xp5_ASAP7_75t_SL g1785 ( 
.A(n_1476),
.B(n_1409),
.Y(n_1785)
);

AND2x4_ASAP7_75t_L g1786 ( 
.A(n_1543),
.B(n_1302),
.Y(n_1786)
);

NAND2xp5_ASAP7_75t_SL g1787 ( 
.A(n_1570),
.B(n_1276),
.Y(n_1787)
);

AO22x1_ASAP7_75t_L g1788 ( 
.A1(n_1439),
.A2(n_1309),
.B1(n_1302),
.B2(n_1412),
.Y(n_1788)
);

OAI22xp33_ASAP7_75t_L g1789 ( 
.A1(n_1555),
.A2(n_1389),
.B1(n_1412),
.B2(n_1282),
.Y(n_1789)
);

INVx1_ASAP7_75t_L g1790 ( 
.A(n_1529),
.Y(n_1790)
);

AOI22xp5_ASAP7_75t_L g1791 ( 
.A1(n_1509),
.A2(n_1309),
.B1(n_1347),
.B2(n_1282),
.Y(n_1791)
);

INVx1_ASAP7_75t_L g1792 ( 
.A(n_1545),
.Y(n_1792)
);

INVx1_ASAP7_75t_L g1793 ( 
.A(n_1545),
.Y(n_1793)
);

AOI22xp5_ASAP7_75t_L g1794 ( 
.A1(n_1590),
.A2(n_952),
.B1(n_958),
.B2(n_951),
.Y(n_1794)
);

OA22x2_ASAP7_75t_L g1795 ( 
.A1(n_1494),
.A2(n_10),
.B1(n_8),
.B2(n_9),
.Y(n_1795)
);

AOI22xp33_ASAP7_75t_L g1796 ( 
.A1(n_1548),
.A2(n_952),
.B1(n_958),
.B2(n_951),
.Y(n_1796)
);

NOR2xp33_ASAP7_75t_L g1797 ( 
.A(n_1482),
.B(n_9),
.Y(n_1797)
);

INVx1_ASAP7_75t_L g1798 ( 
.A(n_1622),
.Y(n_1798)
);

INVx1_ASAP7_75t_L g1799 ( 
.A(n_1514),
.Y(n_1799)
);

INVxp33_ASAP7_75t_L g1800 ( 
.A(n_1569),
.Y(n_1800)
);

INVx2_ASAP7_75t_L g1801 ( 
.A(n_1477),
.Y(n_1801)
);

INVx1_ASAP7_75t_L g1802 ( 
.A(n_1514),
.Y(n_1802)
);

INVx1_ASAP7_75t_L g1803 ( 
.A(n_1515),
.Y(n_1803)
);

INVx1_ASAP7_75t_L g1804 ( 
.A(n_1515),
.Y(n_1804)
);

BUFx6f_ASAP7_75t_L g1805 ( 
.A(n_1638),
.Y(n_1805)
);

INVxp67_ASAP7_75t_SL g1806 ( 
.A(n_1623),
.Y(n_1806)
);

NAND2xp5_ASAP7_75t_L g1807 ( 
.A(n_1563),
.B(n_10),
.Y(n_1807)
);

AND2x4_ASAP7_75t_L g1808 ( 
.A(n_1543),
.B(n_528),
.Y(n_1808)
);

AND2x2_ASAP7_75t_L g1809 ( 
.A(n_1450),
.B(n_11),
.Y(n_1809)
);

INVx4_ASAP7_75t_L g1810 ( 
.A(n_1507),
.Y(n_1810)
);

NAND2xp5_ASAP7_75t_SL g1811 ( 
.A(n_1595),
.B(n_960),
.Y(n_1811)
);

INVx1_ASAP7_75t_L g1812 ( 
.A(n_1477),
.Y(n_1812)
);

BUFx6f_ASAP7_75t_L g1813 ( 
.A(n_1507),
.Y(n_1813)
);

NAND2xp5_ASAP7_75t_L g1814 ( 
.A(n_1564),
.B(n_12),
.Y(n_1814)
);

INVx5_ASAP7_75t_L g1815 ( 
.A(n_1600),
.Y(n_1815)
);

BUFx6f_ASAP7_75t_L g1816 ( 
.A(n_1569),
.Y(n_1816)
);

INVx4_ASAP7_75t_L g1817 ( 
.A(n_1588),
.Y(n_1817)
);

BUFx2_ASAP7_75t_L g1818 ( 
.A(n_1596),
.Y(n_1818)
);

BUFx12f_ASAP7_75t_L g1819 ( 
.A(n_1609),
.Y(n_1819)
);

BUFx6f_ASAP7_75t_L g1820 ( 
.A(n_1600),
.Y(n_1820)
);

INVx4_ASAP7_75t_L g1821 ( 
.A(n_1611),
.Y(n_1821)
);

BUFx6f_ASAP7_75t_L g1822 ( 
.A(n_1600),
.Y(n_1822)
);

OAI22xp33_ASAP7_75t_L g1823 ( 
.A1(n_1542),
.A2(n_22),
.B1(n_30),
.B2(n_13),
.Y(n_1823)
);

NOR2x1_ASAP7_75t_L g1824 ( 
.A(n_1571),
.B(n_958),
.Y(n_1824)
);

AOI22xp33_ASAP7_75t_L g1825 ( 
.A1(n_1558),
.A2(n_1519),
.B1(n_1510),
.B2(n_1501),
.Y(n_1825)
);

INVx2_ASAP7_75t_L g1826 ( 
.A(n_1626),
.Y(n_1826)
);

CKINVDCx5p33_ASAP7_75t_R g1827 ( 
.A(n_1467),
.Y(n_1827)
);

INVx1_ASAP7_75t_L g1828 ( 
.A(n_1538),
.Y(n_1828)
);

INVx2_ASAP7_75t_L g1829 ( 
.A(n_1634),
.Y(n_1829)
);

INVx1_ASAP7_75t_L g1830 ( 
.A(n_1541),
.Y(n_1830)
);

INVx1_ASAP7_75t_L g1831 ( 
.A(n_1544),
.Y(n_1831)
);

BUFx2_ASAP7_75t_L g1832 ( 
.A(n_1468),
.Y(n_1832)
);

NAND2x1p5_ASAP7_75t_L g1833 ( 
.A(n_1448),
.B(n_958),
.Y(n_1833)
);

OAI22xp5_ASAP7_75t_L g1834 ( 
.A1(n_1623),
.A2(n_16),
.B1(n_13),
.B2(n_15),
.Y(n_1834)
);

NAND2xp5_ASAP7_75t_L g1835 ( 
.A(n_1700),
.B(n_1719),
.Y(n_1835)
);

NOR3xp33_ASAP7_75t_SL g1836 ( 
.A(n_1711),
.B(n_1470),
.C(n_1554),
.Y(n_1836)
);

NAND2xp5_ASAP7_75t_L g1837 ( 
.A(n_1784),
.B(n_1513),
.Y(n_1837)
);

INVx3_ASAP7_75t_L g1838 ( 
.A(n_1723),
.Y(n_1838)
);

AOI21xp5_ASAP7_75t_L g1839 ( 
.A1(n_1806),
.A2(n_1445),
.B(n_1483),
.Y(n_1839)
);

OAI22xp5_ASAP7_75t_L g1840 ( 
.A1(n_1798),
.A2(n_1598),
.B1(n_1528),
.B2(n_1513),
.Y(n_1840)
);

AOI22xp5_ASAP7_75t_L g1841 ( 
.A1(n_1809),
.A2(n_1500),
.B1(n_1523),
.B2(n_1442),
.Y(n_1841)
);

INVx1_ASAP7_75t_L g1842 ( 
.A(n_1645),
.Y(n_1842)
);

AOI21xp5_ASAP7_75t_L g1843 ( 
.A1(n_1747),
.A2(n_1789),
.B(n_1765),
.Y(n_1843)
);

OAI22xp5_ASAP7_75t_L g1844 ( 
.A1(n_1692),
.A2(n_1608),
.B1(n_1606),
.B2(n_1593),
.Y(n_1844)
);

AOI21xp5_ASAP7_75t_L g1845 ( 
.A1(n_1747),
.A2(n_1502),
.B(n_1474),
.Y(n_1845)
);

INVx2_ASAP7_75t_SL g1846 ( 
.A(n_1664),
.Y(n_1846)
);

INVx2_ASAP7_75t_L g1847 ( 
.A(n_1646),
.Y(n_1847)
);

NOR2xp33_ASAP7_75t_L g1848 ( 
.A(n_1821),
.B(n_1677),
.Y(n_1848)
);

NAND2xp5_ASAP7_75t_L g1849 ( 
.A(n_1790),
.B(n_1506),
.Y(n_1849)
);

NAND2xp5_ASAP7_75t_L g1850 ( 
.A(n_1792),
.B(n_1585),
.Y(n_1850)
);

INVx1_ASAP7_75t_L g1851 ( 
.A(n_1650),
.Y(n_1851)
);

A2O1A1Ixp33_ASAP7_75t_L g1852 ( 
.A1(n_1751),
.A2(n_1797),
.B(n_1641),
.C(n_1807),
.Y(n_1852)
);

INVx2_ASAP7_75t_L g1853 ( 
.A(n_1648),
.Y(n_1853)
);

OR2x6_ASAP7_75t_L g1854 ( 
.A(n_1640),
.B(n_1502),
.Y(n_1854)
);

NOR2xp33_ASAP7_75t_SL g1855 ( 
.A(n_1776),
.B(n_1468),
.Y(n_1855)
);

INVx1_ASAP7_75t_L g1856 ( 
.A(n_1652),
.Y(n_1856)
);

NAND2xp5_ASAP7_75t_L g1857 ( 
.A(n_1793),
.B(n_1763),
.Y(n_1857)
);

INVx5_ASAP7_75t_L g1858 ( 
.A(n_1820),
.Y(n_1858)
);

INVx3_ASAP7_75t_L g1859 ( 
.A(n_1723),
.Y(n_1859)
);

OAI22xp5_ASAP7_75t_L g1860 ( 
.A1(n_1692),
.A2(n_1610),
.B1(n_1599),
.B2(n_1443),
.Y(n_1860)
);

AO22x1_ASAP7_75t_L g1861 ( 
.A1(n_1694),
.A2(n_1468),
.B1(n_1600),
.B2(n_1568),
.Y(n_1861)
);

INVx1_ASAP7_75t_L g1862 ( 
.A(n_1658),
.Y(n_1862)
);

OAI22x1_ASAP7_75t_L g1863 ( 
.A1(n_1821),
.A2(n_1566),
.B1(n_1522),
.B2(n_1436),
.Y(n_1863)
);

AOI21xp5_ASAP7_75t_L g1864 ( 
.A1(n_1780),
.A2(n_1565),
.B(n_1492),
.Y(n_1864)
);

NOR2xp33_ASAP7_75t_R g1865 ( 
.A(n_1701),
.B(n_1572),
.Y(n_1865)
);

INVx2_ASAP7_75t_L g1866 ( 
.A(n_1649),
.Y(n_1866)
);

NOR3xp33_ASAP7_75t_SL g1867 ( 
.A(n_1834),
.B(n_1587),
.C(n_1576),
.Y(n_1867)
);

NAND2xp5_ASAP7_75t_L g1868 ( 
.A(n_1740),
.B(n_1575),
.Y(n_1868)
);

INVx1_ASAP7_75t_L g1869 ( 
.A(n_1659),
.Y(n_1869)
);

NOR2xp33_ASAP7_75t_L g1870 ( 
.A(n_1818),
.B(n_1536),
.Y(n_1870)
);

NOR3xp33_ASAP7_75t_L g1871 ( 
.A(n_1823),
.B(n_1526),
.C(n_1551),
.Y(n_1871)
);

AOI21xp5_ASAP7_75t_L g1872 ( 
.A1(n_1780),
.A2(n_1565),
.B(n_1492),
.Y(n_1872)
);

NAND2xp5_ASAP7_75t_SL g1873 ( 
.A(n_1820),
.B(n_1822),
.Y(n_1873)
);

INVx1_ASAP7_75t_L g1874 ( 
.A(n_1660),
.Y(n_1874)
);

OAI21x1_ASAP7_75t_L g1875 ( 
.A1(n_1750),
.A2(n_1620),
.B(n_1579),
.Y(n_1875)
);

BUFx6f_ASAP7_75t_L g1876 ( 
.A(n_1656),
.Y(n_1876)
);

HB1xp67_ASAP7_75t_L g1877 ( 
.A(n_1722),
.Y(n_1877)
);

A2O1A1Ixp33_ASAP7_75t_L g1878 ( 
.A1(n_1814),
.A2(n_1557),
.B(n_1589),
.C(n_1625),
.Y(n_1878)
);

OAI21xp5_ASAP7_75t_L g1879 ( 
.A1(n_1834),
.A2(n_1582),
.B(n_1581),
.Y(n_1879)
);

AOI21xp5_ASAP7_75t_L g1880 ( 
.A1(n_1644),
.A2(n_1668),
.B(n_1815),
.Y(n_1880)
);

CKINVDCx6p67_ASAP7_75t_R g1881 ( 
.A(n_1679),
.Y(n_1881)
);

NAND3xp33_ASAP7_75t_L g1882 ( 
.A(n_1742),
.B(n_1616),
.C(n_1479),
.Y(n_1882)
);

A2O1A1Ixp33_ASAP7_75t_L g1883 ( 
.A1(n_1828),
.A2(n_1603),
.B(n_1466),
.C(n_1630),
.Y(n_1883)
);

NAND2xp5_ASAP7_75t_L g1884 ( 
.A(n_1830),
.B(n_17),
.Y(n_1884)
);

NAND3xp33_ASAP7_75t_L g1885 ( 
.A(n_1825),
.B(n_960),
.C(n_959),
.Y(n_1885)
);

NOR2xp33_ASAP7_75t_SL g1886 ( 
.A(n_1776),
.B(n_1817),
.Y(n_1886)
);

AOI21xp5_ASAP7_75t_L g1887 ( 
.A1(n_1815),
.A2(n_960),
.B(n_959),
.Y(n_1887)
);

NAND2xp5_ASAP7_75t_SL g1888 ( 
.A(n_1820),
.B(n_959),
.Y(n_1888)
);

INVxp67_ASAP7_75t_SL g1889 ( 
.A(n_1657),
.Y(n_1889)
);

AOI21xp5_ASAP7_75t_L g1890 ( 
.A1(n_1815),
.A2(n_960),
.B(n_959),
.Y(n_1890)
);

NAND2xp5_ASAP7_75t_SL g1891 ( 
.A(n_1822),
.B(n_959),
.Y(n_1891)
);

INVx2_ASAP7_75t_L g1892 ( 
.A(n_1661),
.Y(n_1892)
);

O2A1O1Ixp33_ASAP7_75t_L g1893 ( 
.A1(n_1831),
.A2(n_19),
.B(n_17),
.C(n_18),
.Y(n_1893)
);

NOR2xp33_ASAP7_75t_L g1894 ( 
.A(n_1703),
.B(n_19),
.Y(n_1894)
);

NAND2xp5_ASAP7_75t_SL g1895 ( 
.A(n_1822),
.B(n_960),
.Y(n_1895)
);

O2A1O1Ixp33_ASAP7_75t_L g1896 ( 
.A1(n_1777),
.A2(n_22),
.B(n_20),
.C(n_21),
.Y(n_1896)
);

O2A1O1Ixp33_ASAP7_75t_L g1897 ( 
.A1(n_1773),
.A2(n_24),
.B(n_21),
.C(n_23),
.Y(n_1897)
);

INVx1_ASAP7_75t_L g1898 ( 
.A(n_1663),
.Y(n_1898)
);

AOI21xp5_ASAP7_75t_L g1899 ( 
.A1(n_1811),
.A2(n_966),
.B(n_962),
.Y(n_1899)
);

AND2x2_ASAP7_75t_L g1900 ( 
.A(n_1662),
.B(n_23),
.Y(n_1900)
);

NOR2xp33_ASAP7_75t_L g1901 ( 
.A(n_1704),
.B(n_24),
.Y(n_1901)
);

O2A1O1Ixp33_ASAP7_75t_L g1902 ( 
.A1(n_1766),
.A2(n_27),
.B(n_25),
.C(n_26),
.Y(n_1902)
);

INVx2_ASAP7_75t_L g1903 ( 
.A(n_1666),
.Y(n_1903)
);

BUFx6f_ASAP7_75t_L g1904 ( 
.A(n_1656),
.Y(n_1904)
);

CKINVDCx20_ASAP7_75t_R g1905 ( 
.A(n_1716),
.Y(n_1905)
);

INVx2_ASAP7_75t_L g1906 ( 
.A(n_1667),
.Y(n_1906)
);

INVx4_ASAP7_75t_L g1907 ( 
.A(n_1653),
.Y(n_1907)
);

BUFx6f_ASAP7_75t_SL g1908 ( 
.A(n_1713),
.Y(n_1908)
);

BUFx2_ASAP7_75t_L g1909 ( 
.A(n_1724),
.Y(n_1909)
);

NAND2xp5_ASAP7_75t_L g1910 ( 
.A(n_1753),
.B(n_26),
.Y(n_1910)
);

NAND2xp5_ASAP7_75t_L g1911 ( 
.A(n_1799),
.B(n_27),
.Y(n_1911)
);

NAND2xp5_ASAP7_75t_SL g1912 ( 
.A(n_1756),
.B(n_962),
.Y(n_1912)
);

A2O1A1Ixp33_ASAP7_75t_L g1913 ( 
.A1(n_1767),
.A2(n_30),
.B(n_28),
.C(n_29),
.Y(n_1913)
);

BUFx2_ASAP7_75t_L g1914 ( 
.A(n_1741),
.Y(n_1914)
);

INVx3_ASAP7_75t_L g1915 ( 
.A(n_1723),
.Y(n_1915)
);

AND2x2_ASAP7_75t_L g1916 ( 
.A(n_1735),
.B(n_28),
.Y(n_1916)
);

NAND2xp5_ASAP7_75t_SL g1917 ( 
.A(n_1736),
.B(n_962),
.Y(n_1917)
);

INVx1_ASAP7_75t_L g1918 ( 
.A(n_1669),
.Y(n_1918)
);

NAND2xp5_ASAP7_75t_L g1919 ( 
.A(n_1802),
.B(n_1803),
.Y(n_1919)
);

INVx2_ASAP7_75t_L g1920 ( 
.A(n_1682),
.Y(n_1920)
);

OAI22xp5_ASAP7_75t_L g1921 ( 
.A1(n_1709),
.A2(n_1744),
.B1(n_1643),
.B2(n_1702),
.Y(n_1921)
);

INVx2_ASAP7_75t_L g1922 ( 
.A(n_1693),
.Y(n_1922)
);

OR2x6_ASAP7_75t_L g1923 ( 
.A(n_1640),
.B(n_962),
.Y(n_1923)
);

NAND2xp5_ASAP7_75t_L g1924 ( 
.A(n_1804),
.B(n_31),
.Y(n_1924)
);

NOR2x1_ASAP7_75t_L g1925 ( 
.A(n_1671),
.B(n_962),
.Y(n_1925)
);

BUFx6f_ASAP7_75t_L g1926 ( 
.A(n_1656),
.Y(n_1926)
);

OAI21x1_ASAP7_75t_L g1927 ( 
.A1(n_1689),
.A2(n_532),
.B(n_531),
.Y(n_1927)
);

AOI21xp5_ASAP7_75t_L g1928 ( 
.A1(n_1689),
.A2(n_969),
.B(n_966),
.Y(n_1928)
);

NAND2xp5_ASAP7_75t_SL g1929 ( 
.A(n_1736),
.B(n_966),
.Y(n_1929)
);

AOI21xp5_ASAP7_75t_L g1930 ( 
.A1(n_1788),
.A2(n_969),
.B(n_966),
.Y(n_1930)
);

BUFx6f_ASAP7_75t_L g1931 ( 
.A(n_1653),
.Y(n_1931)
);

A2O1A1Ixp33_ASAP7_75t_L g1932 ( 
.A1(n_1769),
.A2(n_33),
.B(n_31),
.C(n_32),
.Y(n_1932)
);

AOI33xp33_ASAP7_75t_L g1933 ( 
.A1(n_1782),
.A2(n_34),
.A3(n_36),
.B1(n_37),
.B2(n_33),
.B3(n_35),
.Y(n_1933)
);

BUFx3_ASAP7_75t_L g1934 ( 
.A(n_1748),
.Y(n_1934)
);

NOR2xp33_ASAP7_75t_L g1935 ( 
.A(n_1704),
.B(n_32),
.Y(n_1935)
);

OAI21xp5_ASAP7_75t_L g1936 ( 
.A1(n_1794),
.A2(n_36),
.B(n_38),
.Y(n_1936)
);

NOR2xp33_ASAP7_75t_L g1937 ( 
.A(n_1819),
.B(n_39),
.Y(n_1937)
);

INVx2_ASAP7_75t_L g1938 ( 
.A(n_1697),
.Y(n_1938)
);

NOR2xp33_ASAP7_75t_L g1939 ( 
.A(n_1817),
.B(n_39),
.Y(n_1939)
);

INVx3_ASAP7_75t_L g1940 ( 
.A(n_1762),
.Y(n_1940)
);

NAND2xp5_ASAP7_75t_SL g1941 ( 
.A(n_1759),
.B(n_966),
.Y(n_1941)
);

INVxp67_ASAP7_75t_L g1942 ( 
.A(n_1771),
.Y(n_1942)
);

OAI22xp5_ASAP7_75t_L g1943 ( 
.A1(n_1775),
.A2(n_42),
.B1(n_40),
.B2(n_41),
.Y(n_1943)
);

INVx1_ASAP7_75t_L g1944 ( 
.A(n_1673),
.Y(n_1944)
);

BUFx3_ASAP7_75t_L g1945 ( 
.A(n_1805),
.Y(n_1945)
);

BUFx2_ASAP7_75t_L g1946 ( 
.A(n_1810),
.Y(n_1946)
);

NAND2xp5_ASAP7_75t_L g1947 ( 
.A(n_1783),
.B(n_41),
.Y(n_1947)
);

CKINVDCx16_ASAP7_75t_R g1948 ( 
.A(n_1810),
.Y(n_1948)
);

OAI21xp5_ASAP7_75t_L g1949 ( 
.A1(n_1794),
.A2(n_43),
.B(n_44),
.Y(n_1949)
);

NAND2xp33_ASAP7_75t_R g1950 ( 
.A(n_1827),
.B(n_577),
.Y(n_1950)
);

CKINVDCx5p33_ASAP7_75t_R g1951 ( 
.A(n_1678),
.Y(n_1951)
);

AOI21xp5_ASAP7_75t_L g1952 ( 
.A1(n_1812),
.A2(n_969),
.B(n_43),
.Y(n_1952)
);

OAI21xp5_ASAP7_75t_L g1953 ( 
.A1(n_1829),
.A2(n_44),
.B(n_45),
.Y(n_1953)
);

AOI22x1_ASAP7_75t_L g1954 ( 
.A1(n_1691),
.A2(n_969),
.B1(n_47),
.B2(n_45),
.Y(n_1954)
);

NAND2xp5_ASAP7_75t_L g1955 ( 
.A(n_1642),
.B(n_46),
.Y(n_1955)
);

NAND2x1p5_ASAP7_75t_L g1956 ( 
.A(n_1681),
.B(n_533),
.Y(n_1956)
);

AOI22xp5_ASAP7_75t_L g1957 ( 
.A1(n_1752),
.A2(n_48),
.B1(n_46),
.B2(n_47),
.Y(n_1957)
);

NAND2xp5_ASAP7_75t_L g1958 ( 
.A(n_1801),
.B(n_48),
.Y(n_1958)
);

O2A1O1Ixp33_ASAP7_75t_L g1959 ( 
.A1(n_1779),
.A2(n_51),
.B(n_49),
.C(n_50),
.Y(n_1959)
);

NOR2xp33_ASAP7_75t_L g1960 ( 
.A(n_1743),
.B(n_1725),
.Y(n_1960)
);

NAND2xp5_ASAP7_75t_L g1961 ( 
.A(n_1687),
.B(n_50),
.Y(n_1961)
);

NOR2xp33_ASAP7_75t_L g1962 ( 
.A(n_1678),
.B(n_52),
.Y(n_1962)
);

NOR2xp33_ASAP7_75t_L g1963 ( 
.A(n_1670),
.B(n_53),
.Y(n_1963)
);

HB1xp67_ASAP7_75t_L g1964 ( 
.A(n_1657),
.Y(n_1964)
);

OAI22xp5_ASAP7_75t_SL g1965 ( 
.A1(n_1749),
.A2(n_1698),
.B1(n_1781),
.B2(n_1795),
.Y(n_1965)
);

NOR2xp33_ASAP7_75t_L g1966 ( 
.A(n_1754),
.B(n_53),
.Y(n_1966)
);

INVx3_ASAP7_75t_L g1967 ( 
.A(n_1762),
.Y(n_1967)
);

OAI22xp5_ASAP7_75t_L g1968 ( 
.A1(n_1706),
.A2(n_56),
.B1(n_54),
.B2(n_55),
.Y(n_1968)
);

INVx1_ASAP7_75t_L g1969 ( 
.A(n_1695),
.Y(n_1969)
);

AOI21xp5_ASAP7_75t_L g1970 ( 
.A1(n_1647),
.A2(n_55),
.B(n_56),
.Y(n_1970)
);

NAND3xp33_ASAP7_75t_SL g1971 ( 
.A(n_1683),
.B(n_57),
.C(n_58),
.Y(n_1971)
);

INVx1_ASAP7_75t_L g1972 ( 
.A(n_1699),
.Y(n_1972)
);

INVx2_ASAP7_75t_L g1973 ( 
.A(n_1705),
.Y(n_1973)
);

NAND2xp5_ASAP7_75t_SL g1974 ( 
.A(n_1759),
.B(n_57),
.Y(n_1974)
);

INVx2_ASAP7_75t_L g1975 ( 
.A(n_1721),
.Y(n_1975)
);

O2A1O1Ixp33_ASAP7_75t_L g1976 ( 
.A1(n_1787),
.A2(n_60),
.B(n_58),
.C(n_59),
.Y(n_1976)
);

OAI22xp5_ASAP7_75t_L g1977 ( 
.A1(n_1675),
.A2(n_62),
.B1(n_59),
.B2(n_61),
.Y(n_1977)
);

BUFx12f_ASAP7_75t_L g1978 ( 
.A(n_1781),
.Y(n_1978)
);

NOR2xp33_ASAP7_75t_L g1979 ( 
.A(n_1805),
.B(n_61),
.Y(n_1979)
);

BUFx4f_ASAP7_75t_L g1980 ( 
.A(n_1762),
.Y(n_1980)
);

AOI21xp5_ASAP7_75t_L g1981 ( 
.A1(n_1647),
.A2(n_63),
.B(n_65),
.Y(n_1981)
);

BUFx2_ASAP7_75t_L g1982 ( 
.A(n_1681),
.Y(n_1982)
);

NAND2xp5_ASAP7_75t_L g1983 ( 
.A(n_1707),
.B(n_63),
.Y(n_1983)
);

NAND2xp5_ASAP7_75t_L g1984 ( 
.A(n_1708),
.B(n_65),
.Y(n_1984)
);

INVx1_ASAP7_75t_L g1985 ( 
.A(n_1710),
.Y(n_1985)
);

NAND2xp5_ASAP7_75t_L g1986 ( 
.A(n_1745),
.B(n_66),
.Y(n_1986)
);

AOI22xp33_ASAP7_75t_L g1987 ( 
.A1(n_1781),
.A2(n_1739),
.B1(n_1733),
.B2(n_1738),
.Y(n_1987)
);

OAI22xp5_ASAP7_75t_L g1988 ( 
.A1(n_1691),
.A2(n_1749),
.B1(n_1655),
.B2(n_1640),
.Y(n_1988)
);

NAND2xp5_ASAP7_75t_SL g1989 ( 
.A(n_1813),
.B(n_66),
.Y(n_1989)
);

AOI22xp33_ASAP7_75t_L g1990 ( 
.A1(n_1726),
.A2(n_69),
.B1(n_67),
.B2(n_68),
.Y(n_1990)
);

OAI21xp33_ASAP7_75t_SL g1991 ( 
.A1(n_1791),
.A2(n_70),
.B(n_69),
.Y(n_1991)
);

INVx1_ASAP7_75t_L g1992 ( 
.A(n_1714),
.Y(n_1992)
);

INVx3_ASAP7_75t_L g1993 ( 
.A(n_1762),
.Y(n_1993)
);

NAND2xp5_ASAP7_75t_L g1994 ( 
.A(n_1816),
.B(n_68),
.Y(n_1994)
);

OR2x2_ASAP7_75t_SL g1995 ( 
.A(n_1813),
.B(n_70),
.Y(n_1995)
);

AOI21xp5_ASAP7_75t_L g1996 ( 
.A1(n_1824),
.A2(n_72),
.B(n_73),
.Y(n_1996)
);

INVx2_ASAP7_75t_L g1997 ( 
.A(n_1718),
.Y(n_1997)
);

INVx1_ASAP7_75t_L g1998 ( 
.A(n_1720),
.Y(n_1998)
);

O2A1O1Ixp5_ASAP7_75t_L g1999 ( 
.A1(n_1826),
.A2(n_74),
.B(n_72),
.C(n_73),
.Y(n_1999)
);

AOI21xp5_ASAP7_75t_L g2000 ( 
.A1(n_1824),
.A2(n_74),
.B(n_75),
.Y(n_2000)
);

NAND2xp5_ASAP7_75t_SL g2001 ( 
.A(n_1813),
.B(n_76),
.Y(n_2001)
);

INVx1_ASAP7_75t_SL g2002 ( 
.A(n_1816),
.Y(n_2002)
);

AOI21xp5_ASAP7_75t_L g2003 ( 
.A1(n_1737),
.A2(n_76),
.B(n_77),
.Y(n_2003)
);

AOI22xp33_ASAP7_75t_L g2004 ( 
.A1(n_1729),
.A2(n_80),
.B1(n_78),
.B2(n_79),
.Y(n_2004)
);

INVx1_ASAP7_75t_L g2005 ( 
.A(n_1730),
.Y(n_2005)
);

NAND2xp5_ASAP7_75t_L g2006 ( 
.A(n_1816),
.B(n_78),
.Y(n_2006)
);

NAND2xp5_ASAP7_75t_L g2007 ( 
.A(n_1717),
.B(n_80),
.Y(n_2007)
);

BUFx6f_ASAP7_75t_L g2008 ( 
.A(n_1931),
.Y(n_2008)
);

NAND2xp5_ASAP7_75t_L g2009 ( 
.A(n_1835),
.B(n_1717),
.Y(n_2009)
);

AOI21xp5_ASAP7_75t_L g2010 ( 
.A1(n_1839),
.A2(n_1715),
.B(n_1712),
.Y(n_2010)
);

INVx1_ASAP7_75t_L g2011 ( 
.A(n_1842),
.Y(n_2011)
);

NOR2xp33_ASAP7_75t_R g2012 ( 
.A(n_1905),
.B(n_1948),
.Y(n_2012)
);

AND2x2_ASAP7_75t_L g2013 ( 
.A(n_1914),
.B(n_1786),
.Y(n_2013)
);

OR2x6_ASAP7_75t_L g2014 ( 
.A(n_1854),
.B(n_1655),
.Y(n_2014)
);

NAND2xp5_ASAP7_75t_L g2015 ( 
.A(n_1889),
.B(n_1757),
.Y(n_2015)
);

INVx2_ASAP7_75t_SL g2016 ( 
.A(n_1846),
.Y(n_2016)
);

NAND3xp33_ASAP7_75t_L g2017 ( 
.A(n_1962),
.B(n_1731),
.C(n_1665),
.Y(n_2017)
);

INVx2_ASAP7_75t_L g2018 ( 
.A(n_1997),
.Y(n_2018)
);

INVx2_ASAP7_75t_L g2019 ( 
.A(n_1847),
.Y(n_2019)
);

INVx1_ASAP7_75t_L g2020 ( 
.A(n_1851),
.Y(n_2020)
);

BUFx2_ASAP7_75t_L g2021 ( 
.A(n_1909),
.Y(n_2021)
);

INVx8_ASAP7_75t_L g2022 ( 
.A(n_1908),
.Y(n_2022)
);

NAND2xp5_ASAP7_75t_L g2023 ( 
.A(n_1964),
.B(n_1761),
.Y(n_2023)
);

INVx2_ASAP7_75t_L g2024 ( 
.A(n_1853),
.Y(n_2024)
);

BUFx8_ASAP7_75t_SL g2025 ( 
.A(n_1908),
.Y(n_2025)
);

INVx1_ASAP7_75t_L g2026 ( 
.A(n_1856),
.Y(n_2026)
);

INVx5_ASAP7_75t_L g2027 ( 
.A(n_1923),
.Y(n_2027)
);

BUFx6f_ASAP7_75t_L g2028 ( 
.A(n_1931),
.Y(n_2028)
);

AOI22xp5_ASAP7_75t_L g2029 ( 
.A1(n_1860),
.A2(n_1808),
.B1(n_1786),
.B2(n_1696),
.Y(n_2029)
);

HB1xp67_ASAP7_75t_L g2030 ( 
.A(n_1877),
.Y(n_2030)
);

BUFx3_ASAP7_75t_L g2031 ( 
.A(n_1881),
.Y(n_2031)
);

NAND2xp5_ASAP7_75t_L g2032 ( 
.A(n_1857),
.B(n_1805),
.Y(n_2032)
);

INVx2_ASAP7_75t_L g2033 ( 
.A(n_1866),
.Y(n_2033)
);

NAND2xp5_ASAP7_75t_L g2034 ( 
.A(n_1919),
.B(n_1681),
.Y(n_2034)
);

CKINVDCx11_ASAP7_75t_R g2035 ( 
.A(n_1978),
.Y(n_2035)
);

INVx2_ASAP7_75t_L g2036 ( 
.A(n_1892),
.Y(n_2036)
);

NOR2xp33_ASAP7_75t_L g2037 ( 
.A(n_1848),
.B(n_1758),
.Y(n_2037)
);

CKINVDCx5p33_ASAP7_75t_R g2038 ( 
.A(n_1865),
.Y(n_2038)
);

INVx2_ASAP7_75t_L g2039 ( 
.A(n_1903),
.Y(n_2039)
);

HB1xp67_ASAP7_75t_L g2040 ( 
.A(n_1862),
.Y(n_2040)
);

AOI222xp33_ASAP7_75t_L g2041 ( 
.A1(n_1965),
.A2(n_1808),
.B1(n_1796),
.B2(n_1800),
.C1(n_1760),
.C2(n_1832),
.Y(n_2041)
);

OAI22x1_ASAP7_75t_L g2042 ( 
.A1(n_1951),
.A2(n_1791),
.B1(n_1785),
.B2(n_1768),
.Y(n_2042)
);

AOI21xp5_ASAP7_75t_L g2043 ( 
.A1(n_1936),
.A2(n_1655),
.B(n_1737),
.Y(n_2043)
);

HB1xp67_ASAP7_75t_L g2044 ( 
.A(n_1869),
.Y(n_2044)
);

INVx2_ASAP7_75t_L g2045 ( 
.A(n_1906),
.Y(n_2045)
);

AOI22xp33_ASAP7_75t_L g2046 ( 
.A1(n_1965),
.A2(n_1732),
.B1(n_1734),
.B2(n_1764),
.Y(n_2046)
);

INVx2_ASAP7_75t_L g2047 ( 
.A(n_1920),
.Y(n_2047)
);

INVx1_ASAP7_75t_L g2048 ( 
.A(n_1874),
.Y(n_2048)
);

NAND2xp5_ASAP7_75t_L g2049 ( 
.A(n_1849),
.B(n_1685),
.Y(n_2049)
);

INVx1_ASAP7_75t_L g2050 ( 
.A(n_1898),
.Y(n_2050)
);

NAND2xp5_ASAP7_75t_L g2051 ( 
.A(n_1868),
.B(n_1685),
.Y(n_2051)
);

CKINVDCx16_ASAP7_75t_R g2052 ( 
.A(n_1886),
.Y(n_2052)
);

INVx3_ASAP7_75t_L g2053 ( 
.A(n_1931),
.Y(n_2053)
);

AOI22xp5_ASAP7_75t_L g2054 ( 
.A1(n_1901),
.A2(n_1690),
.B1(n_1760),
.B2(n_1772),
.Y(n_2054)
);

INVx1_ASAP7_75t_L g2055 ( 
.A(n_1918),
.Y(n_2055)
);

NAND2xp5_ASAP7_75t_SL g2056 ( 
.A(n_1980),
.B(n_1760),
.Y(n_2056)
);

AOI21xp33_ASAP7_75t_L g2057 ( 
.A1(n_1949),
.A2(n_1770),
.B(n_1772),
.Y(n_2057)
);

AOI22xp33_ASAP7_75t_L g2058 ( 
.A1(n_1935),
.A2(n_1772),
.B1(n_1690),
.B2(n_1684),
.Y(n_2058)
);

OAI22xp5_ASAP7_75t_L g2059 ( 
.A1(n_1957),
.A2(n_1690),
.B1(n_1778),
.B2(n_1774),
.Y(n_2059)
);

BUFx3_ASAP7_75t_L g2060 ( 
.A(n_1934),
.Y(n_2060)
);

AND2x2_ASAP7_75t_L g2061 ( 
.A(n_1916),
.B(n_1727),
.Y(n_2061)
);

AOI21xp5_ASAP7_75t_L g2062 ( 
.A1(n_1843),
.A2(n_1755),
.B(n_1688),
.Y(n_2062)
);

AOI22xp33_ASAP7_75t_L g2063 ( 
.A1(n_1844),
.A2(n_1684),
.B1(n_1651),
.B2(n_1833),
.Y(n_2063)
);

AOI21xp5_ASAP7_75t_L g2064 ( 
.A1(n_1980),
.A2(n_1755),
.B(n_1688),
.Y(n_2064)
);

INVx1_ASAP7_75t_L g2065 ( 
.A(n_1944),
.Y(n_2065)
);

INVx3_ASAP7_75t_L g2066 ( 
.A(n_1907),
.Y(n_2066)
);

INVx2_ASAP7_75t_SL g2067 ( 
.A(n_1945),
.Y(n_2067)
);

INVx5_ASAP7_75t_SL g2068 ( 
.A(n_1876),
.Y(n_2068)
);

CKINVDCx5p33_ASAP7_75t_R g2069 ( 
.A(n_1836),
.Y(n_2069)
);

NAND2xp5_ASAP7_75t_L g2070 ( 
.A(n_1850),
.B(n_1685),
.Y(n_2070)
);

INVx2_ASAP7_75t_L g2071 ( 
.A(n_1922),
.Y(n_2071)
);

NAND2xp5_ASAP7_75t_L g2072 ( 
.A(n_1837),
.B(n_1969),
.Y(n_2072)
);

BUFx6f_ASAP7_75t_L g2073 ( 
.A(n_1876),
.Y(n_2073)
);

BUFx3_ASAP7_75t_L g2074 ( 
.A(n_1876),
.Y(n_2074)
);

INVx1_ASAP7_75t_L g2075 ( 
.A(n_1972),
.Y(n_2075)
);

NAND2xp5_ASAP7_75t_L g2076 ( 
.A(n_1985),
.B(n_1992),
.Y(n_2076)
);

INVx2_ASAP7_75t_SL g2077 ( 
.A(n_1904),
.Y(n_2077)
);

AND2x2_ASAP7_75t_L g2078 ( 
.A(n_1900),
.B(n_1727),
.Y(n_2078)
);

BUFx4f_ASAP7_75t_L g2079 ( 
.A(n_1904),
.Y(n_2079)
);

OAI22xp5_ASAP7_75t_SL g2080 ( 
.A1(n_1995),
.A2(n_1778),
.B1(n_1774),
.B2(n_1654),
.Y(n_2080)
);

INVx2_ASAP7_75t_SL g2081 ( 
.A(n_1904),
.Y(n_2081)
);

NAND2xp5_ASAP7_75t_L g2082 ( 
.A(n_1852),
.B(n_1686),
.Y(n_2082)
);

NAND2xp5_ASAP7_75t_L g2083 ( 
.A(n_1845),
.B(n_1998),
.Y(n_2083)
);

INVx1_ASAP7_75t_L g2084 ( 
.A(n_2005),
.Y(n_2084)
);

INVx2_ASAP7_75t_L g2085 ( 
.A(n_1938),
.Y(n_2085)
);

INVx4_ASAP7_75t_L g2086 ( 
.A(n_1926),
.Y(n_2086)
);

BUFx2_ASAP7_75t_L g2087 ( 
.A(n_1982),
.Y(n_2087)
);

BUFx6f_ASAP7_75t_L g2088 ( 
.A(n_1926),
.Y(n_2088)
);

BUFx3_ASAP7_75t_L g2089 ( 
.A(n_1926),
.Y(n_2089)
);

AOI22xp5_ASAP7_75t_L g2090 ( 
.A1(n_1957),
.A2(n_1651),
.B1(n_1746),
.B2(n_1676),
.Y(n_2090)
);

HB1xp67_ASAP7_75t_L g2091 ( 
.A(n_1942),
.Y(n_2091)
);

AND2x2_ASAP7_75t_L g2092 ( 
.A(n_1966),
.B(n_1728),
.Y(n_2092)
);

INVx5_ASAP7_75t_L g2093 ( 
.A(n_1923),
.Y(n_2093)
);

CKINVDCx20_ASAP7_75t_R g2094 ( 
.A(n_1870),
.Y(n_2094)
);

INVx1_ASAP7_75t_L g2095 ( 
.A(n_1973),
.Y(n_2095)
);

HB1xp67_ASAP7_75t_L g2096 ( 
.A(n_1921),
.Y(n_2096)
);

INVx5_ASAP7_75t_L g2097 ( 
.A(n_1923),
.Y(n_2097)
);

NAND2xp5_ASAP7_75t_L g2098 ( 
.A(n_1960),
.B(n_1686),
.Y(n_2098)
);

NAND2xp5_ASAP7_75t_L g2099 ( 
.A(n_1879),
.B(n_1686),
.Y(n_2099)
);

INVx2_ASAP7_75t_L g2100 ( 
.A(n_1975),
.Y(n_2100)
);

INVx1_ASAP7_75t_L g2101 ( 
.A(n_1961),
.Y(n_2101)
);

AND2x2_ASAP7_75t_L g2102 ( 
.A(n_1979),
.B(n_1728),
.Y(n_2102)
);

INVx2_ASAP7_75t_L g2103 ( 
.A(n_1986),
.Y(n_2103)
);

BUFx6f_ASAP7_75t_L g2104 ( 
.A(n_1858),
.Y(n_2104)
);

INVx2_ASAP7_75t_L g2105 ( 
.A(n_1958),
.Y(n_2105)
);

OAI22xp5_ASAP7_75t_L g2106 ( 
.A1(n_1840),
.A2(n_1841),
.B1(n_1953),
.B2(n_1932),
.Y(n_2106)
);

INVx3_ASAP7_75t_L g2107 ( 
.A(n_1907),
.Y(n_2107)
);

BUFx2_ASAP7_75t_L g2108 ( 
.A(n_1946),
.Y(n_2108)
);

AOI22xp33_ASAP7_75t_L g2109 ( 
.A1(n_1882),
.A2(n_1746),
.B1(n_1672),
.B2(n_1680),
.Y(n_2109)
);

NAND2xp5_ASAP7_75t_L g2110 ( 
.A(n_1955),
.B(n_1654),
.Y(n_2110)
);

INVx4_ASAP7_75t_L g2111 ( 
.A(n_1838),
.Y(n_2111)
);

OR2x2_ASAP7_75t_L g2112 ( 
.A(n_1983),
.B(n_81),
.Y(n_2112)
);

AOI221xp5_ASAP7_75t_L g2113 ( 
.A1(n_1893),
.A2(n_1674),
.B1(n_83),
.B2(n_81),
.C(n_82),
.Y(n_2113)
);

BUFx6f_ASAP7_75t_L g2114 ( 
.A(n_1858),
.Y(n_2114)
);

INVx3_ASAP7_75t_L g2115 ( 
.A(n_1940),
.Y(n_2115)
);

NAND2xp5_ASAP7_75t_L g2116 ( 
.A(n_1911),
.B(n_82),
.Y(n_2116)
);

BUFx2_ASAP7_75t_L g2117 ( 
.A(n_1838),
.Y(n_2117)
);

INVx4_ASAP7_75t_L g2118 ( 
.A(n_1859),
.Y(n_2118)
);

INVx2_ASAP7_75t_SL g2119 ( 
.A(n_1859),
.Y(n_2119)
);

AND2x4_ASAP7_75t_L g2120 ( 
.A(n_1940),
.B(n_1967),
.Y(n_2120)
);

NOR2xp33_ASAP7_75t_L g2121 ( 
.A(n_1894),
.B(n_83),
.Y(n_2121)
);

OAI22xp5_ASAP7_75t_L g2122 ( 
.A1(n_1841),
.A2(n_94),
.B1(n_102),
.B2(n_85),
.Y(n_2122)
);

INVx2_ASAP7_75t_L g2123 ( 
.A(n_1910),
.Y(n_2123)
);

INVxp67_ASAP7_75t_L g2124 ( 
.A(n_1884),
.Y(n_2124)
);

INVx1_ASAP7_75t_L g2125 ( 
.A(n_1984),
.Y(n_2125)
);

AOI22xp33_ASAP7_75t_SL g2126 ( 
.A1(n_1991),
.A2(n_96),
.B1(n_104),
.B2(n_86),
.Y(n_2126)
);

NAND2xp5_ASAP7_75t_L g2127 ( 
.A(n_1924),
.B(n_87),
.Y(n_2127)
);

INVx1_ASAP7_75t_L g2128 ( 
.A(n_1947),
.Y(n_2128)
);

AND2x4_ASAP7_75t_L g2129 ( 
.A(n_1967),
.B(n_537),
.Y(n_2129)
);

NOR2xp33_ASAP7_75t_SL g2130 ( 
.A(n_2038),
.B(n_1855),
.Y(n_2130)
);

AO32x2_ASAP7_75t_L g2131 ( 
.A1(n_2106),
.A2(n_1988),
.A3(n_1977),
.B1(n_1943),
.B2(n_1968),
.Y(n_2131)
);

AO31x2_ASAP7_75t_L g2132 ( 
.A1(n_2106),
.A2(n_2042),
.A3(n_2083),
.B(n_2015),
.Y(n_2132)
);

NAND2xp5_ASAP7_75t_L g2133 ( 
.A(n_2030),
.B(n_1933),
.Y(n_2133)
);

INVx2_ASAP7_75t_L g2134 ( 
.A(n_2018),
.Y(n_2134)
);

INVx1_ASAP7_75t_L g2135 ( 
.A(n_2040),
.Y(n_2135)
);

A2O1A1Ixp33_ASAP7_75t_L g2136 ( 
.A1(n_2096),
.A2(n_1867),
.B(n_1897),
.C(n_1896),
.Y(n_2136)
);

A2O1A1Ixp33_ASAP7_75t_L g2137 ( 
.A1(n_2122),
.A2(n_1991),
.B(n_1902),
.C(n_1959),
.Y(n_2137)
);

A2O1A1Ixp33_ASAP7_75t_L g2138 ( 
.A1(n_2122),
.A2(n_1882),
.B(n_2113),
.C(n_1939),
.Y(n_2138)
);

A2O1A1Ixp33_ASAP7_75t_L g2139 ( 
.A1(n_2029),
.A2(n_1963),
.B(n_1871),
.C(n_1883),
.Y(n_2139)
);

A2O1A1Ixp33_ASAP7_75t_L g2140 ( 
.A1(n_2029),
.A2(n_1913),
.B(n_1976),
.C(n_1937),
.Y(n_2140)
);

AOI21xp5_ASAP7_75t_L g2141 ( 
.A1(n_2062),
.A2(n_2010),
.B(n_2043),
.Y(n_2141)
);

INVx1_ASAP7_75t_L g2142 ( 
.A(n_2044),
.Y(n_2142)
);

AO31x2_ASAP7_75t_L g2143 ( 
.A1(n_2083),
.A2(n_2015),
.A3(n_2059),
.B(n_1864),
.Y(n_2143)
);

A2O1A1Ixp33_ASAP7_75t_L g2144 ( 
.A1(n_2046),
.A2(n_1981),
.B(n_1970),
.C(n_2003),
.Y(n_2144)
);

A2O1A1Ixp33_ASAP7_75t_L g2145 ( 
.A1(n_2121),
.A2(n_1999),
.B(n_1974),
.C(n_1996),
.Y(n_2145)
);

AOI21xp5_ASAP7_75t_L g2146 ( 
.A1(n_2059),
.A2(n_1928),
.B(n_1885),
.Y(n_2146)
);

BUFx12f_ASAP7_75t_L g2147 ( 
.A(n_2035),
.Y(n_2147)
);

AOI22xp33_ASAP7_75t_L g2148 ( 
.A1(n_2041),
.A2(n_1987),
.B1(n_1854),
.B2(n_1971),
.Y(n_2148)
);

OAI22xp33_ASAP7_75t_L g2149 ( 
.A1(n_2052),
.A2(n_1854),
.B1(n_1950),
.B2(n_1993),
.Y(n_2149)
);

NOR2xp33_ASAP7_75t_L g2150 ( 
.A(n_2069),
.B(n_1915),
.Y(n_2150)
);

AND2x2_ASAP7_75t_L g2151 ( 
.A(n_2013),
.B(n_1915),
.Y(n_2151)
);

A2O1A1Ixp33_ASAP7_75t_L g2152 ( 
.A1(n_2124),
.A2(n_2000),
.B(n_1878),
.C(n_1952),
.Y(n_2152)
);

CKINVDCx5p33_ASAP7_75t_R g2153 ( 
.A(n_2025),
.Y(n_2153)
);

AOI21xp5_ASAP7_75t_L g2154 ( 
.A1(n_2064),
.A2(n_1885),
.B(n_1872),
.Y(n_2154)
);

INVx2_ASAP7_75t_SL g2155 ( 
.A(n_2022),
.Y(n_2155)
);

NAND2xp5_ASAP7_75t_L g2156 ( 
.A(n_2072),
.B(n_1912),
.Y(n_2156)
);

NOR2xp33_ASAP7_75t_L g2157 ( 
.A(n_2037),
.B(n_1994),
.Y(n_2157)
);

NAND2xp5_ASAP7_75t_L g2158 ( 
.A(n_2091),
.B(n_2007),
.Y(n_2158)
);

HB1xp67_ASAP7_75t_L g2159 ( 
.A(n_2021),
.Y(n_2159)
);

A2O1A1Ixp33_ASAP7_75t_L g2160 ( 
.A1(n_2126),
.A2(n_2004),
.B(n_1990),
.C(n_1993),
.Y(n_2160)
);

NOR2xp67_ASAP7_75t_SL g2161 ( 
.A(n_2104),
.B(n_1858),
.Y(n_2161)
);

INVx2_ASAP7_75t_L g2162 ( 
.A(n_2084),
.Y(n_2162)
);

AOI221x1_ASAP7_75t_L g2163 ( 
.A1(n_2017),
.A2(n_2082),
.B1(n_2125),
.B2(n_2101),
.C(n_1863),
.Y(n_2163)
);

HB1xp67_ASAP7_75t_L g2164 ( 
.A(n_2087),
.Y(n_2164)
);

OAI22xp33_ASAP7_75t_L g2165 ( 
.A1(n_2090),
.A2(n_1954),
.B1(n_2006),
.B2(n_2001),
.Y(n_2165)
);

CKINVDCx11_ASAP7_75t_R g2166 ( 
.A(n_2094),
.Y(n_2166)
);

OAI22xp5_ASAP7_75t_L g2167 ( 
.A1(n_2080),
.A2(n_1989),
.B1(n_1925),
.B2(n_1956),
.Y(n_2167)
);

AOI21xp5_ASAP7_75t_L g2168 ( 
.A1(n_2099),
.A2(n_2080),
.B(n_1930),
.Y(n_2168)
);

OAI22xp5_ASAP7_75t_L g2169 ( 
.A1(n_2112),
.A2(n_1880),
.B1(n_1929),
.B2(n_1917),
.Y(n_2169)
);

INVx2_ASAP7_75t_SL g2170 ( 
.A(n_2022),
.Y(n_2170)
);

AOI221x1_ASAP7_75t_L g2171 ( 
.A1(n_2017),
.A2(n_1899),
.B1(n_1887),
.B2(n_1890),
.C(n_1861),
.Y(n_2171)
);

AOI21xp5_ASAP7_75t_L g2172 ( 
.A1(n_2099),
.A2(n_1927),
.B(n_1941),
.Y(n_2172)
);

AOI22xp33_ASAP7_75t_L g2173 ( 
.A1(n_2041),
.A2(n_1873),
.B1(n_2002),
.B2(n_1875),
.Y(n_2173)
);

INVx4_ASAP7_75t_L g2174 ( 
.A(n_2073),
.Y(n_2174)
);

INVx1_ASAP7_75t_L g2175 ( 
.A(n_2076),
.Y(n_2175)
);

O2A1O1Ixp33_ASAP7_75t_SL g2176 ( 
.A1(n_2116),
.A2(n_90),
.B(n_87),
.C(n_89),
.Y(n_2176)
);

OAI21x1_ASAP7_75t_L g2177 ( 
.A1(n_2066),
.A2(n_1891),
.B(n_1888),
.Y(n_2177)
);

A2O1A1Ixp33_ASAP7_75t_L g2178 ( 
.A1(n_2127),
.A2(n_1895),
.B(n_91),
.C(n_89),
.Y(n_2178)
);

BUFx12f_ASAP7_75t_L g2179 ( 
.A(n_2031),
.Y(n_2179)
);

A2O1A1Ixp33_ASAP7_75t_L g2180 ( 
.A1(n_2054),
.A2(n_92),
.B(n_90),
.C(n_91),
.Y(n_2180)
);

OAI22xp5_ASAP7_75t_L g2181 ( 
.A1(n_2063),
.A2(n_95),
.B1(n_92),
.B2(n_93),
.Y(n_2181)
);

O2A1O1Ixp33_ASAP7_75t_SL g2182 ( 
.A1(n_2110),
.A2(n_97),
.B(n_93),
.C(n_95),
.Y(n_2182)
);

A2O1A1Ixp33_ASAP7_75t_L g2183 ( 
.A1(n_2054),
.A2(n_99),
.B(n_97),
.C(n_98),
.Y(n_2183)
);

AOI22xp33_ASAP7_75t_L g2184 ( 
.A1(n_2123),
.A2(n_100),
.B1(n_98),
.B2(n_99),
.Y(n_2184)
);

AOI21xp5_ASAP7_75t_SL g2185 ( 
.A1(n_2129),
.A2(n_2014),
.B(n_2056),
.Y(n_2185)
);

NAND3xp33_ASAP7_75t_SL g2186 ( 
.A(n_2012),
.B(n_101),
.C(n_102),
.Y(n_2186)
);

OAI21x1_ASAP7_75t_L g2187 ( 
.A1(n_2066),
.A2(n_2107),
.B(n_2053),
.Y(n_2187)
);

OAI21x1_ASAP7_75t_L g2188 ( 
.A1(n_2107),
.A2(n_539),
.B(n_538),
.Y(n_2188)
);

OR2x6_ASAP7_75t_L g2189 ( 
.A(n_2022),
.B(n_542),
.Y(n_2189)
);

INVx1_ASAP7_75t_L g2190 ( 
.A(n_2076),
.Y(n_2190)
);

NAND2xp5_ASAP7_75t_L g2191 ( 
.A(n_2032),
.B(n_101),
.Y(n_2191)
);

OAI22xp5_ASAP7_75t_L g2192 ( 
.A1(n_2090),
.A2(n_2109),
.B1(n_2058),
.B2(n_2060),
.Y(n_2192)
);

INVx1_ASAP7_75t_L g2193 ( 
.A(n_2011),
.Y(n_2193)
);

NAND2xp5_ASAP7_75t_L g2194 ( 
.A(n_2108),
.B(n_103),
.Y(n_2194)
);

O2A1O1Ixp33_ASAP7_75t_SL g2195 ( 
.A1(n_2016),
.A2(n_105),
.B(n_103),
.C(n_104),
.Y(n_2195)
);

OAI21x1_ASAP7_75t_L g2196 ( 
.A1(n_2053),
.A2(n_545),
.B(n_543),
.Y(n_2196)
);

INVx1_ASAP7_75t_L g2197 ( 
.A(n_2020),
.Y(n_2197)
);

INVx2_ASAP7_75t_L g2198 ( 
.A(n_2019),
.Y(n_2198)
);

AOI21xp5_ASAP7_75t_L g2199 ( 
.A1(n_2027),
.A2(n_105),
.B(n_106),
.Y(n_2199)
);

AO32x2_ASAP7_75t_L g2200 ( 
.A1(n_2067),
.A2(n_109),
.A3(n_107),
.B1(n_108),
.B2(n_110),
.Y(n_2200)
);

A2O1A1Ixp33_ASAP7_75t_L g2201 ( 
.A1(n_2057),
.A2(n_111),
.B(n_109),
.C(n_110),
.Y(n_2201)
);

BUFx2_ASAP7_75t_L g2202 ( 
.A(n_2117),
.Y(n_2202)
);

OAI22xp5_ASAP7_75t_L g2203 ( 
.A1(n_2138),
.A2(n_2014),
.B1(n_2079),
.B2(n_2092),
.Y(n_2203)
);

HB1xp67_ASAP7_75t_L g2204 ( 
.A(n_2135),
.Y(n_2204)
);

CKINVDCx5p33_ASAP7_75t_R g2205 ( 
.A(n_2166),
.Y(n_2205)
);

CKINVDCx5p33_ASAP7_75t_R g2206 ( 
.A(n_2147),
.Y(n_2206)
);

AOI22xp33_ASAP7_75t_L g2207 ( 
.A1(n_2148),
.A2(n_2105),
.B1(n_2103),
.B2(n_2057),
.Y(n_2207)
);

O2A1O1Ixp5_ASAP7_75t_L g2208 ( 
.A1(n_2139),
.A2(n_2128),
.B(n_2034),
.C(n_2098),
.Y(n_2208)
);

INVx1_ASAP7_75t_L g2209 ( 
.A(n_2142),
.Y(n_2209)
);

AOI22xp33_ASAP7_75t_SL g2210 ( 
.A1(n_2192),
.A2(n_2061),
.B1(n_2078),
.B2(n_2009),
.Y(n_2210)
);

OAI221xp5_ASAP7_75t_L g2211 ( 
.A1(n_2136),
.A2(n_2049),
.B1(n_2051),
.B2(n_2070),
.C(n_2050),
.Y(n_2211)
);

INVx1_ASAP7_75t_L g2212 ( 
.A(n_2193),
.Y(n_2212)
);

AOI21xp33_ASAP7_75t_L g2213 ( 
.A1(n_2165),
.A2(n_2023),
.B(n_2026),
.Y(n_2213)
);

A2O1A1Ixp33_ASAP7_75t_L g2214 ( 
.A1(n_2140),
.A2(n_2129),
.B(n_2102),
.C(n_2055),
.Y(n_2214)
);

INVxp67_ASAP7_75t_L g2215 ( 
.A(n_2202),
.Y(n_2215)
);

AOI22xp33_ASAP7_75t_L g2216 ( 
.A1(n_2186),
.A2(n_2014),
.B1(n_2095),
.B2(n_2033),
.Y(n_2216)
);

OAI22xp33_ASAP7_75t_L g2217 ( 
.A1(n_2133),
.A2(n_2093),
.B1(n_2097),
.B2(n_2027),
.Y(n_2217)
);

OR2x2_ASAP7_75t_L g2218 ( 
.A(n_2159),
.B(n_2048),
.Y(n_2218)
);

INVx2_ASAP7_75t_L g2219 ( 
.A(n_2162),
.Y(n_2219)
);

OAI221xp5_ASAP7_75t_L g2220 ( 
.A1(n_2137),
.A2(n_2075),
.B1(n_2065),
.B2(n_2023),
.C(n_2119),
.Y(n_2220)
);

INVx1_ASAP7_75t_L g2221 ( 
.A(n_2197),
.Y(n_2221)
);

AOI22xp33_ASAP7_75t_L g2222 ( 
.A1(n_2181),
.A2(n_2120),
.B1(n_2024),
.B2(n_2039),
.Y(n_2222)
);

OAI22xp33_ASAP7_75t_L g2223 ( 
.A1(n_2163),
.A2(n_2146),
.B1(n_2154),
.B2(n_2189),
.Y(n_2223)
);

NAND2xp5_ASAP7_75t_L g2224 ( 
.A(n_2175),
.B(n_2115),
.Y(n_2224)
);

CKINVDCx6p67_ASAP7_75t_R g2225 ( 
.A(n_2179),
.Y(n_2225)
);

OAI22xp33_ASAP7_75t_L g2226 ( 
.A1(n_2189),
.A2(n_2027),
.B1(n_2097),
.B2(n_2093),
.Y(n_2226)
);

INVx2_ASAP7_75t_L g2227 ( 
.A(n_2134),
.Y(n_2227)
);

INVx2_ASAP7_75t_L g2228 ( 
.A(n_2198),
.Y(n_2228)
);

INVx2_ASAP7_75t_L g2229 ( 
.A(n_2190),
.Y(n_2229)
);

INVx1_ASAP7_75t_L g2230 ( 
.A(n_2164),
.Y(n_2230)
);

OAI22xp5_ASAP7_75t_L g2231 ( 
.A1(n_2145),
.A2(n_2079),
.B1(n_2115),
.B2(n_2068),
.Y(n_2231)
);

OAI22xp5_ASAP7_75t_L g2232 ( 
.A1(n_2180),
.A2(n_2068),
.B1(n_2097),
.B2(n_2093),
.Y(n_2232)
);

AO31x2_ASAP7_75t_L g2233 ( 
.A1(n_2141),
.A2(n_2045),
.A3(n_2047),
.B(n_2036),
.Y(n_2233)
);

AND2x2_ASAP7_75t_L g2234 ( 
.A(n_2151),
.B(n_2158),
.Y(n_2234)
);

OAI22xp5_ASAP7_75t_L g2235 ( 
.A1(n_2183),
.A2(n_2118),
.B1(n_2111),
.B2(n_2120),
.Y(n_2235)
);

AND2x4_ASAP7_75t_L g2236 ( 
.A(n_2143),
.B(n_2074),
.Y(n_2236)
);

AOI22xp33_ASAP7_75t_L g2237 ( 
.A1(n_2149),
.A2(n_2173),
.B1(n_2199),
.B2(n_2085),
.Y(n_2237)
);

INVx2_ASAP7_75t_L g2238 ( 
.A(n_2132),
.Y(n_2238)
);

AOI22xp33_ASAP7_75t_L g2239 ( 
.A1(n_2157),
.A2(n_2100),
.B1(n_2071),
.B2(n_2169),
.Y(n_2239)
);

OAI22xp5_ASAP7_75t_L g2240 ( 
.A1(n_2144),
.A2(n_2111),
.B1(n_2118),
.B2(n_2089),
.Y(n_2240)
);

OAI21xp33_ASAP7_75t_L g2241 ( 
.A1(n_2152),
.A2(n_2081),
.B(n_2077),
.Y(n_2241)
);

NAND2xp5_ASAP7_75t_L g2242 ( 
.A(n_2156),
.B(n_2073),
.Y(n_2242)
);

NAND2xp5_ASAP7_75t_L g2243 ( 
.A(n_2143),
.B(n_2073),
.Y(n_2243)
);

INVx1_ASAP7_75t_L g2244 ( 
.A(n_2132),
.Y(n_2244)
);

INVx2_ASAP7_75t_L g2245 ( 
.A(n_2132),
.Y(n_2245)
);

OAI22xp5_ASAP7_75t_L g2246 ( 
.A1(n_2201),
.A2(n_2160),
.B1(n_2184),
.B2(n_2178),
.Y(n_2246)
);

INVx1_ASAP7_75t_L g2247 ( 
.A(n_2143),
.Y(n_2247)
);

INVx2_ASAP7_75t_SL g2248 ( 
.A(n_2155),
.Y(n_2248)
);

AOI22xp5_ASAP7_75t_L g2249 ( 
.A1(n_2130),
.A2(n_2114),
.B1(n_2104),
.B2(n_2028),
.Y(n_2249)
);

OAI22xp5_ASAP7_75t_L g2250 ( 
.A1(n_2194),
.A2(n_2167),
.B1(n_2191),
.B2(n_2168),
.Y(n_2250)
);

AO31x2_ASAP7_75t_L g2251 ( 
.A1(n_2238),
.A2(n_2171),
.A3(n_2172),
.B(n_2174),
.Y(n_2251)
);

NOR2xp33_ASAP7_75t_L g2252 ( 
.A(n_2205),
.B(n_2153),
.Y(n_2252)
);

OAI22xp33_ASAP7_75t_L g2253 ( 
.A1(n_2220),
.A2(n_2200),
.B1(n_2131),
.B2(n_2114),
.Y(n_2253)
);

INVx2_ASAP7_75t_L g2254 ( 
.A(n_2233),
.Y(n_2254)
);

OAI21xp5_ASAP7_75t_L g2255 ( 
.A1(n_2223),
.A2(n_2182),
.B(n_2176),
.Y(n_2255)
);

INVx1_ASAP7_75t_L g2256 ( 
.A(n_2204),
.Y(n_2256)
);

NAND2xp5_ASAP7_75t_L g2257 ( 
.A(n_2204),
.B(n_2229),
.Y(n_2257)
);

OAI21xp5_ASAP7_75t_L g2258 ( 
.A1(n_2223),
.A2(n_2208),
.B(n_2246),
.Y(n_2258)
);

INVx3_ASAP7_75t_L g2259 ( 
.A(n_2236),
.Y(n_2259)
);

INVx2_ASAP7_75t_L g2260 ( 
.A(n_2233),
.Y(n_2260)
);

HB1xp67_ASAP7_75t_L g2261 ( 
.A(n_2247),
.Y(n_2261)
);

BUFx3_ASAP7_75t_L g2262 ( 
.A(n_2206),
.Y(n_2262)
);

INVx2_ASAP7_75t_L g2263 ( 
.A(n_2233),
.Y(n_2263)
);

AOI21x1_ASAP7_75t_L g2264 ( 
.A1(n_2244),
.A2(n_2187),
.B(n_2161),
.Y(n_2264)
);

BUFx4f_ASAP7_75t_SL g2265 ( 
.A(n_2225),
.Y(n_2265)
);

AND2x2_ASAP7_75t_L g2266 ( 
.A(n_2234),
.B(n_2174),
.Y(n_2266)
);

INVx11_ASAP7_75t_L g2267 ( 
.A(n_2248),
.Y(n_2267)
);

INVx1_ASAP7_75t_L g2268 ( 
.A(n_2212),
.Y(n_2268)
);

AOI22xp33_ASAP7_75t_L g2269 ( 
.A1(n_2207),
.A2(n_2150),
.B1(n_2131),
.B2(n_2170),
.Y(n_2269)
);

INVx1_ASAP7_75t_L g2270 ( 
.A(n_2221),
.Y(n_2270)
);

INVx2_ASAP7_75t_L g2271 ( 
.A(n_2233),
.Y(n_2271)
);

AOI22xp5_ASAP7_75t_L g2272 ( 
.A1(n_2250),
.A2(n_2195),
.B1(n_2131),
.B2(n_2200),
.Y(n_2272)
);

INVx1_ASAP7_75t_L g2273 ( 
.A(n_2209),
.Y(n_2273)
);

AOI22xp33_ASAP7_75t_L g2274 ( 
.A1(n_2237),
.A2(n_2216),
.B1(n_2210),
.B2(n_2211),
.Y(n_2274)
);

INVx1_ASAP7_75t_L g2275 ( 
.A(n_2219),
.Y(n_2275)
);

BUFx2_ASAP7_75t_L g2276 ( 
.A(n_2236),
.Y(n_2276)
);

AND2x2_ASAP7_75t_L g2277 ( 
.A(n_2215),
.B(n_2200),
.Y(n_2277)
);

INVx4_ASAP7_75t_L g2278 ( 
.A(n_2218),
.Y(n_2278)
);

OAI221xp5_ASAP7_75t_L g2279 ( 
.A1(n_2258),
.A2(n_2208),
.B1(n_2210),
.B2(n_2214),
.C(n_2239),
.Y(n_2279)
);

OAI22xp5_ASAP7_75t_L g2280 ( 
.A1(n_2269),
.A2(n_2272),
.B1(n_2258),
.B2(n_2253),
.Y(n_2280)
);

OAI22xp5_ASAP7_75t_L g2281 ( 
.A1(n_2272),
.A2(n_2203),
.B1(n_2215),
.B2(n_2231),
.Y(n_2281)
);

AOI22xp33_ASAP7_75t_SL g2282 ( 
.A1(n_2255),
.A2(n_2232),
.B1(n_2245),
.B2(n_2243),
.Y(n_2282)
);

OAI22xp5_ASAP7_75t_L g2283 ( 
.A1(n_2253),
.A2(n_2240),
.B1(n_2235),
.B2(n_2230),
.Y(n_2283)
);

INVxp67_ASAP7_75t_L g2284 ( 
.A(n_2277),
.Y(n_2284)
);

AND2x4_ASAP7_75t_L g2285 ( 
.A(n_2278),
.B(n_2224),
.Y(n_2285)
);

OAI211xp5_ASAP7_75t_L g2286 ( 
.A1(n_2255),
.A2(n_2213),
.B(n_2241),
.C(n_2222),
.Y(n_2286)
);

AOI22x1_ASAP7_75t_L g2287 ( 
.A1(n_2278),
.A2(n_2086),
.B1(n_2088),
.B2(n_2028),
.Y(n_2287)
);

BUFx3_ASAP7_75t_L g2288 ( 
.A(n_2262),
.Y(n_2288)
);

OR2x2_ASAP7_75t_L g2289 ( 
.A(n_2257),
.B(n_2242),
.Y(n_2289)
);

OAI22xp5_ASAP7_75t_L g2290 ( 
.A1(n_2274),
.A2(n_2222),
.B1(n_2249),
.B2(n_2185),
.Y(n_2290)
);

NOR3xp33_ASAP7_75t_L g2291 ( 
.A(n_2280),
.B(n_2277),
.C(n_2278),
.Y(n_2291)
);

INVx2_ASAP7_75t_L g2292 ( 
.A(n_2289),
.Y(n_2292)
);

INVx2_ASAP7_75t_L g2293 ( 
.A(n_2285),
.Y(n_2293)
);

INVx1_ASAP7_75t_L g2294 ( 
.A(n_2284),
.Y(n_2294)
);

OR2x2_ASAP7_75t_L g2295 ( 
.A(n_2283),
.B(n_2257),
.Y(n_2295)
);

HB1xp67_ASAP7_75t_L g2296 ( 
.A(n_2281),
.Y(n_2296)
);

INVx2_ASAP7_75t_SL g2297 ( 
.A(n_2288),
.Y(n_2297)
);

OR2x2_ASAP7_75t_L g2298 ( 
.A(n_2285),
.B(n_2256),
.Y(n_2298)
);

NAND4xp25_ASAP7_75t_L g2299 ( 
.A(n_2291),
.B(n_2286),
.C(n_2279),
.D(n_2282),
.Y(n_2299)
);

NAND3xp33_ASAP7_75t_L g2300 ( 
.A(n_2296),
.B(n_2261),
.C(n_2290),
.Y(n_2300)
);

AND2x2_ASAP7_75t_L g2301 ( 
.A(n_2297),
.B(n_2278),
.Y(n_2301)
);

AOI221xp5_ASAP7_75t_L g2302 ( 
.A1(n_2291),
.A2(n_2261),
.B1(n_2276),
.B2(n_2273),
.C(n_2270),
.Y(n_2302)
);

INVx2_ASAP7_75t_L g2303 ( 
.A(n_2298),
.Y(n_2303)
);

AOI211xp5_ASAP7_75t_L g2304 ( 
.A1(n_2296),
.A2(n_2295),
.B(n_2294),
.C(n_2293),
.Y(n_2304)
);

AND2x4_ASAP7_75t_L g2305 ( 
.A(n_2292),
.B(n_2262),
.Y(n_2305)
);

INVx1_ASAP7_75t_L g2306 ( 
.A(n_2294),
.Y(n_2306)
);

AND2x2_ASAP7_75t_L g2307 ( 
.A(n_2297),
.B(n_2266),
.Y(n_2307)
);

INVx1_ASAP7_75t_L g2308 ( 
.A(n_2294),
.Y(n_2308)
);

NAND2xp5_ASAP7_75t_L g2309 ( 
.A(n_2304),
.B(n_2256),
.Y(n_2309)
);

NAND2xp5_ASAP7_75t_L g2310 ( 
.A(n_2304),
.B(n_2268),
.Y(n_2310)
);

AND2x2_ASAP7_75t_L g2311 ( 
.A(n_2307),
.B(n_2262),
.Y(n_2311)
);

NAND2x1p5_ASAP7_75t_L g2312 ( 
.A(n_2305),
.B(n_2287),
.Y(n_2312)
);

NAND2xp5_ASAP7_75t_L g2313 ( 
.A(n_2306),
.B(n_2273),
.Y(n_2313)
);

OR2x2_ASAP7_75t_SL g2314 ( 
.A(n_2300),
.B(n_2265),
.Y(n_2314)
);

INVx3_ASAP7_75t_L g2315 ( 
.A(n_2305),
.Y(n_2315)
);

AND2x2_ASAP7_75t_L g2316 ( 
.A(n_2301),
.B(n_2252),
.Y(n_2316)
);

INVx2_ASAP7_75t_L g2317 ( 
.A(n_2303),
.Y(n_2317)
);

INVx1_ASAP7_75t_L g2318 ( 
.A(n_2308),
.Y(n_2318)
);

INVx1_ASAP7_75t_L g2319 ( 
.A(n_2299),
.Y(n_2319)
);

NAND2xp5_ASAP7_75t_L g2320 ( 
.A(n_2302),
.B(n_2268),
.Y(n_2320)
);

AND2x2_ASAP7_75t_L g2321 ( 
.A(n_2315),
.B(n_2266),
.Y(n_2321)
);

HB1xp67_ASAP7_75t_L g2322 ( 
.A(n_2315),
.Y(n_2322)
);

INVx1_ASAP7_75t_L g2323 ( 
.A(n_2313),
.Y(n_2323)
);

AND2x2_ASAP7_75t_L g2324 ( 
.A(n_2311),
.B(n_2276),
.Y(n_2324)
);

AOI21xp33_ASAP7_75t_L g2325 ( 
.A1(n_2310),
.A2(n_2260),
.B(n_2254),
.Y(n_2325)
);

INVx1_ASAP7_75t_L g2326 ( 
.A(n_2318),
.Y(n_2326)
);

INVx3_ASAP7_75t_L g2327 ( 
.A(n_2312),
.Y(n_2327)
);

AND2x2_ASAP7_75t_L g2328 ( 
.A(n_2316),
.B(n_2259),
.Y(n_2328)
);

OR2x2_ASAP7_75t_L g2329 ( 
.A(n_2309),
.B(n_2270),
.Y(n_2329)
);

NAND2xp5_ASAP7_75t_L g2330 ( 
.A(n_2322),
.B(n_2319),
.Y(n_2330)
);

OR2x2_ASAP7_75t_L g2331 ( 
.A(n_2323),
.B(n_2310),
.Y(n_2331)
);

AND2x2_ASAP7_75t_L g2332 ( 
.A(n_2321),
.B(n_2312),
.Y(n_2332)
);

INVx1_ASAP7_75t_L g2333 ( 
.A(n_2326),
.Y(n_2333)
);

INVx1_ASAP7_75t_L g2334 ( 
.A(n_2330),
.Y(n_2334)
);

CKINVDCx5p33_ASAP7_75t_R g2335 ( 
.A(n_2330),
.Y(n_2335)
);

OR2x2_ASAP7_75t_L g2336 ( 
.A(n_2331),
.B(n_2309),
.Y(n_2336)
);

INVx1_ASAP7_75t_L g2337 ( 
.A(n_2333),
.Y(n_2337)
);

AND2x2_ASAP7_75t_L g2338 ( 
.A(n_2335),
.B(n_2332),
.Y(n_2338)
);

OAI22xp33_ASAP7_75t_L g2339 ( 
.A1(n_2335),
.A2(n_2327),
.B1(n_2320),
.B2(n_2317),
.Y(n_2339)
);

AOI22xp5_ASAP7_75t_L g2340 ( 
.A1(n_2334),
.A2(n_2327),
.B1(n_2324),
.B2(n_2321),
.Y(n_2340)
);

NAND2xp5_ASAP7_75t_L g2341 ( 
.A(n_2337),
.B(n_2327),
.Y(n_2341)
);

OR2x2_ASAP7_75t_L g2342 ( 
.A(n_2336),
.B(n_2329),
.Y(n_2342)
);

AOI211x1_ASAP7_75t_L g2343 ( 
.A1(n_2334),
.A2(n_2324),
.B(n_2328),
.C(n_2325),
.Y(n_2343)
);

INVx1_ASAP7_75t_SL g2344 ( 
.A(n_2338),
.Y(n_2344)
);

NOR2xp33_ASAP7_75t_SL g2345 ( 
.A(n_2342),
.B(n_2265),
.Y(n_2345)
);

NAND2xp5_ASAP7_75t_L g2346 ( 
.A(n_2340),
.B(n_2328),
.Y(n_2346)
);

INVx1_ASAP7_75t_L g2347 ( 
.A(n_2341),
.Y(n_2347)
);

OR2x2_ASAP7_75t_L g2348 ( 
.A(n_2339),
.B(n_2314),
.Y(n_2348)
);

OR2x2_ASAP7_75t_L g2349 ( 
.A(n_2343),
.B(n_2259),
.Y(n_2349)
);

AND2x4_ASAP7_75t_SL g2350 ( 
.A(n_2338),
.B(n_2267),
.Y(n_2350)
);

INVx1_ASAP7_75t_L g2351 ( 
.A(n_2342),
.Y(n_2351)
);

BUFx2_ASAP7_75t_L g2352 ( 
.A(n_2338),
.Y(n_2352)
);

NOR2xp33_ASAP7_75t_L g2353 ( 
.A(n_2338),
.B(n_2267),
.Y(n_2353)
);

AOI322xp5_ASAP7_75t_L g2354 ( 
.A1(n_2351),
.A2(n_2217),
.A3(n_2271),
.B1(n_2260),
.B2(n_2263),
.C1(n_2254),
.C2(n_2226),
.Y(n_2354)
);

AND2x2_ASAP7_75t_L g2355 ( 
.A(n_2352),
.B(n_2259),
.Y(n_2355)
);

NAND2xp5_ASAP7_75t_L g2356 ( 
.A(n_2344),
.B(n_2259),
.Y(n_2356)
);

NAND2xp5_ASAP7_75t_L g2357 ( 
.A(n_2347),
.B(n_2251),
.Y(n_2357)
);

INVx2_ASAP7_75t_SL g2358 ( 
.A(n_2350),
.Y(n_2358)
);

O2A1O1Ixp33_ASAP7_75t_L g2359 ( 
.A1(n_2346),
.A2(n_2217),
.B(n_2226),
.C(n_113),
.Y(n_2359)
);

INVx2_ASAP7_75t_L g2360 ( 
.A(n_2348),
.Y(n_2360)
);

NAND4xp25_ASAP7_75t_L g2361 ( 
.A(n_2345),
.B(n_2086),
.C(n_113),
.D(n_111),
.Y(n_2361)
);

INVx1_ASAP7_75t_L g2362 ( 
.A(n_2349),
.Y(n_2362)
);

NOR2xp33_ASAP7_75t_L g2363 ( 
.A(n_2353),
.B(n_2264),
.Y(n_2363)
);

A2O1A1Ixp33_ASAP7_75t_L g2364 ( 
.A1(n_2351),
.A2(n_2254),
.B(n_2263),
.C(n_2260),
.Y(n_2364)
);

INVx1_ASAP7_75t_L g2365 ( 
.A(n_2352),
.Y(n_2365)
);

NAND2x1p5_ASAP7_75t_SL g2366 ( 
.A(n_2352),
.B(n_112),
.Y(n_2366)
);

OR2x2_ASAP7_75t_L g2367 ( 
.A(n_2365),
.B(n_114),
.Y(n_2367)
);

XNOR2x1_ASAP7_75t_L g2368 ( 
.A(n_2360),
.B(n_115),
.Y(n_2368)
);

NAND3x1_ASAP7_75t_L g2369 ( 
.A(n_2362),
.B(n_2264),
.C(n_115),
.Y(n_2369)
);

INVx1_ASAP7_75t_L g2370 ( 
.A(n_2366),
.Y(n_2370)
);

INVxp67_ASAP7_75t_L g2371 ( 
.A(n_2358),
.Y(n_2371)
);

NAND2x1p5_ASAP7_75t_L g2372 ( 
.A(n_2355),
.B(n_2356),
.Y(n_2372)
);

NAND2xp5_ASAP7_75t_L g2373 ( 
.A(n_2361),
.B(n_2251),
.Y(n_2373)
);

INVx1_ASAP7_75t_L g2374 ( 
.A(n_2357),
.Y(n_2374)
);

INVx1_ASAP7_75t_L g2375 ( 
.A(n_2359),
.Y(n_2375)
);

NAND2xp5_ASAP7_75t_L g2376 ( 
.A(n_2363),
.B(n_2251),
.Y(n_2376)
);

NOR2xp33_ASAP7_75t_SL g2377 ( 
.A(n_2364),
.B(n_2088),
.Y(n_2377)
);

NAND2xp5_ASAP7_75t_L g2378 ( 
.A(n_2354),
.B(n_2251),
.Y(n_2378)
);

NAND2xp5_ASAP7_75t_L g2379 ( 
.A(n_2365),
.B(n_2251),
.Y(n_2379)
);

INVxp67_ASAP7_75t_SL g2380 ( 
.A(n_2365),
.Y(n_2380)
);

INVx2_ASAP7_75t_SL g2381 ( 
.A(n_2355),
.Y(n_2381)
);

INVx1_ASAP7_75t_L g2382 ( 
.A(n_2380),
.Y(n_2382)
);

NAND2xp5_ASAP7_75t_L g2383 ( 
.A(n_2370),
.B(n_2368),
.Y(n_2383)
);

AND2x2_ASAP7_75t_L g2384 ( 
.A(n_2371),
.B(n_2251),
.Y(n_2384)
);

INVxp33_ASAP7_75t_L g2385 ( 
.A(n_2372),
.Y(n_2385)
);

NAND2x1p5_ASAP7_75t_L g2386 ( 
.A(n_2381),
.B(n_2188),
.Y(n_2386)
);

INVx1_ASAP7_75t_SL g2387 ( 
.A(n_2367),
.Y(n_2387)
);

NOR2xp33_ASAP7_75t_L g2388 ( 
.A(n_2375),
.B(n_116),
.Y(n_2388)
);

NAND2xp5_ASAP7_75t_L g2389 ( 
.A(n_2369),
.B(n_117),
.Y(n_2389)
);

INVx1_ASAP7_75t_L g2390 ( 
.A(n_2379),
.Y(n_2390)
);

AND2x2_ASAP7_75t_SL g2391 ( 
.A(n_2374),
.B(n_2088),
.Y(n_2391)
);

AOI22xp5_ASAP7_75t_L g2392 ( 
.A1(n_2373),
.A2(n_2271),
.B1(n_2263),
.B2(n_2275),
.Y(n_2392)
);

AOI22xp5_ASAP7_75t_L g2393 ( 
.A1(n_2376),
.A2(n_2271),
.B1(n_2275),
.B2(n_2028),
.Y(n_2393)
);

NAND2xp5_ASAP7_75t_L g2394 ( 
.A(n_2378),
.B(n_2377),
.Y(n_2394)
);

OAI21xp5_ASAP7_75t_L g2395 ( 
.A1(n_2380),
.A2(n_2196),
.B(n_2177),
.Y(n_2395)
);

INVx2_ASAP7_75t_L g2396 ( 
.A(n_2386),
.Y(n_2396)
);

NAND2xp5_ASAP7_75t_SL g2397 ( 
.A(n_2385),
.B(n_2008),
.Y(n_2397)
);

INVx1_ASAP7_75t_SL g2398 ( 
.A(n_2382),
.Y(n_2398)
);

AOI221x1_ASAP7_75t_SL g2399 ( 
.A1(n_2383),
.A2(n_119),
.B1(n_117),
.B2(n_118),
.C(n_120),
.Y(n_2399)
);

XNOR2x1_ASAP7_75t_L g2400 ( 
.A(n_2387),
.B(n_118),
.Y(n_2400)
);

AOI22xp33_ASAP7_75t_L g2401 ( 
.A1(n_2390),
.A2(n_2008),
.B1(n_2228),
.B2(n_2227),
.Y(n_2401)
);

NOR3x1_ASAP7_75t_L g2402 ( 
.A(n_2389),
.B(n_119),
.C(n_120),
.Y(n_2402)
);

NOR2xp33_ASAP7_75t_L g2403 ( 
.A(n_2388),
.B(n_121),
.Y(n_2403)
);

INVx1_ASAP7_75t_L g2404 ( 
.A(n_2391),
.Y(n_2404)
);

AND2x2_ASAP7_75t_L g2405 ( 
.A(n_2384),
.B(n_121),
.Y(n_2405)
);

AOI21xp5_ASAP7_75t_SL g2406 ( 
.A1(n_2394),
.A2(n_122),
.B(n_123),
.Y(n_2406)
);

INVx1_ASAP7_75t_L g2407 ( 
.A(n_2392),
.Y(n_2407)
);

AND2x4_ASAP7_75t_L g2408 ( 
.A(n_2395),
.B(n_122),
.Y(n_2408)
);

INVx2_ASAP7_75t_L g2409 ( 
.A(n_2393),
.Y(n_2409)
);

INVx1_ASAP7_75t_L g2410 ( 
.A(n_2389),
.Y(n_2410)
);

INVx1_ASAP7_75t_L g2411 ( 
.A(n_2389),
.Y(n_2411)
);

A2O1A1Ixp33_ASAP7_75t_L g2412 ( 
.A1(n_2382),
.A2(n_125),
.B(n_123),
.C(n_124),
.Y(n_2412)
);

NAND2xp5_ASAP7_75t_SL g2413 ( 
.A(n_2385),
.B(n_2008),
.Y(n_2413)
);

XOR2x2_ASAP7_75t_L g2414 ( 
.A(n_2383),
.B(n_124),
.Y(n_2414)
);

INVx1_ASAP7_75t_L g2415 ( 
.A(n_2389),
.Y(n_2415)
);

INVx2_ASAP7_75t_L g2416 ( 
.A(n_2386),
.Y(n_2416)
);

OR2x2_ASAP7_75t_L g2417 ( 
.A(n_2382),
.B(n_125),
.Y(n_2417)
);

NAND3xp33_ASAP7_75t_L g2418 ( 
.A(n_2400),
.B(n_126),
.C(n_127),
.Y(n_2418)
);

XNOR2xp5_ASAP7_75t_L g2419 ( 
.A(n_2414),
.B(n_126),
.Y(n_2419)
);

XNOR2xp5_ASAP7_75t_L g2420 ( 
.A(n_2399),
.B(n_2398),
.Y(n_2420)
);

OR2x2_ASAP7_75t_L g2421 ( 
.A(n_2417),
.B(n_128),
.Y(n_2421)
);

NAND2xp5_ASAP7_75t_SL g2422 ( 
.A(n_2412),
.B(n_2396),
.Y(n_2422)
);

AOI22x1_ASAP7_75t_SL g2423 ( 
.A1(n_2410),
.A2(n_130),
.B1(n_128),
.B2(n_129),
.Y(n_2423)
);

OAI21xp33_ASAP7_75t_SL g2424 ( 
.A1(n_2397),
.A2(n_129),
.B(n_130),
.Y(n_2424)
);

AND2x2_ASAP7_75t_L g2425 ( 
.A(n_2411),
.B(n_131),
.Y(n_2425)
);

NOR2x1_ASAP7_75t_L g2426 ( 
.A(n_2406),
.B(n_131),
.Y(n_2426)
);

AO22x2_ASAP7_75t_L g2427 ( 
.A1(n_2415),
.A2(n_135),
.B1(n_132),
.B2(n_133),
.Y(n_2427)
);

NOR5xp2_ASAP7_75t_L g2428 ( 
.A(n_2404),
.B(n_135),
.C(n_132),
.D(n_133),
.E(n_137),
.Y(n_2428)
);

NAND2xp5_ASAP7_75t_L g2429 ( 
.A(n_2402),
.B(n_138),
.Y(n_2429)
);

AO22x1_ASAP7_75t_L g2430 ( 
.A1(n_2416),
.A2(n_140),
.B1(n_138),
.B2(n_139),
.Y(n_2430)
);

A2O1A1Ixp33_ASAP7_75t_L g2431 ( 
.A1(n_2408),
.A2(n_141),
.B(n_139),
.C(n_140),
.Y(n_2431)
);

NOR2x1_ASAP7_75t_L g2432 ( 
.A(n_2403),
.B(n_141),
.Y(n_2432)
);

NAND2xp5_ASAP7_75t_L g2433 ( 
.A(n_2405),
.B(n_142),
.Y(n_2433)
);

OR2x2_ASAP7_75t_L g2434 ( 
.A(n_2413),
.B(n_142),
.Y(n_2434)
);

NAND5xp2_ASAP7_75t_L g2435 ( 
.A(n_2407),
.B(n_145),
.C(n_143),
.D(n_144),
.E(n_146),
.Y(n_2435)
);

OAI22xp5_ASAP7_75t_L g2436 ( 
.A1(n_2408),
.A2(n_2114),
.B1(n_2104),
.B2(n_145),
.Y(n_2436)
);

AND4x1_ASAP7_75t_L g2437 ( 
.A(n_2407),
.B(n_146),
.C(n_143),
.D(n_144),
.Y(n_2437)
);

AOI21xp5_ASAP7_75t_L g2438 ( 
.A1(n_2409),
.A2(n_147),
.B(n_148),
.Y(n_2438)
);

NOR2xp33_ASAP7_75t_L g2439 ( 
.A(n_2401),
.B(n_147),
.Y(n_2439)
);

NOR3xp33_ASAP7_75t_L g2440 ( 
.A(n_2398),
.B(n_148),
.C(n_149),
.Y(n_2440)
);

NAND4xp25_ASAP7_75t_L g2441 ( 
.A(n_2402),
.B(n_151),
.C(n_149),
.D(n_150),
.Y(n_2441)
);

NOR2x1_ASAP7_75t_L g2442 ( 
.A(n_2417),
.B(n_150),
.Y(n_2442)
);

AND2x2_ASAP7_75t_L g2443 ( 
.A(n_2398),
.B(n_151),
.Y(n_2443)
);

NOR3xp33_ASAP7_75t_SL g2444 ( 
.A(n_2410),
.B(n_152),
.C(n_153),
.Y(n_2444)
);

AND2x2_ASAP7_75t_L g2445 ( 
.A(n_2398),
.B(n_154),
.Y(n_2445)
);

NAND2xp5_ASAP7_75t_L g2446 ( 
.A(n_2399),
.B(n_154),
.Y(n_2446)
);

NOR2xp33_ASAP7_75t_SL g2447 ( 
.A(n_2398),
.B(n_155),
.Y(n_2447)
);

NOR2xp33_ASAP7_75t_L g2448 ( 
.A(n_2398),
.B(n_155),
.Y(n_2448)
);

NAND2xp5_ASAP7_75t_L g2449 ( 
.A(n_2399),
.B(n_157),
.Y(n_2449)
);

NAND2x1_ASAP7_75t_SL g2450 ( 
.A(n_2396),
.B(n_157),
.Y(n_2450)
);

NOR3xp33_ASAP7_75t_L g2451 ( 
.A(n_2398),
.B(n_159),
.C(n_160),
.Y(n_2451)
);

NAND4xp25_ASAP7_75t_SL g2452 ( 
.A(n_2398),
.B(n_162),
.C(n_159),
.D(n_160),
.Y(n_2452)
);

NOR4xp75_ASAP7_75t_L g2453 ( 
.A(n_2397),
.B(n_164),
.C(n_162),
.D(n_163),
.Y(n_2453)
);

AOI211x1_ASAP7_75t_SL g2454 ( 
.A1(n_2396),
.A2(n_165),
.B(n_163),
.C(n_164),
.Y(n_2454)
);

OAI31xp33_ASAP7_75t_L g2455 ( 
.A1(n_2420),
.A2(n_167),
.A3(n_165),
.B(n_166),
.Y(n_2455)
);

NOR2xp33_ASAP7_75t_SL g2456 ( 
.A(n_2443),
.B(n_166),
.Y(n_2456)
);

OAI21xp5_ASAP7_75t_L g2457 ( 
.A1(n_2424),
.A2(n_2449),
.B(n_2446),
.Y(n_2457)
);

AOI21xp33_ASAP7_75t_L g2458 ( 
.A1(n_2419),
.A2(n_167),
.B(n_168),
.Y(n_2458)
);

OR2x2_ASAP7_75t_L g2459 ( 
.A(n_2441),
.B(n_168),
.Y(n_2459)
);

XNOR2x1_ASAP7_75t_L g2460 ( 
.A(n_2426),
.B(n_169),
.Y(n_2460)
);

OAI21xp5_ASAP7_75t_L g2461 ( 
.A1(n_2418),
.A2(n_170),
.B(n_171),
.Y(n_2461)
);

OAI22xp5_ASAP7_75t_L g2462 ( 
.A1(n_2448),
.A2(n_172),
.B1(n_170),
.B2(n_171),
.Y(n_2462)
);

CKINVDCx5p33_ASAP7_75t_R g2463 ( 
.A(n_2444),
.Y(n_2463)
);

NAND3xp33_ASAP7_75t_SL g2464 ( 
.A(n_2454),
.B(n_172),
.C(n_173),
.Y(n_2464)
);

OR2x2_ASAP7_75t_L g2465 ( 
.A(n_2435),
.B(n_174),
.Y(n_2465)
);

AND2x2_ASAP7_75t_L g2466 ( 
.A(n_2445),
.B(n_174),
.Y(n_2466)
);

AOI21xp5_ASAP7_75t_L g2467 ( 
.A1(n_2422),
.A2(n_175),
.B(n_176),
.Y(n_2467)
);

OAI21xp5_ASAP7_75t_L g2468 ( 
.A1(n_2429),
.A2(n_176),
.B(n_177),
.Y(n_2468)
);

OAI21xp33_ASAP7_75t_SL g2469 ( 
.A1(n_2450),
.A2(n_177),
.B(n_178),
.Y(n_2469)
);

INVx1_ASAP7_75t_L g2470 ( 
.A(n_2427),
.Y(n_2470)
);

AOI221xp5_ASAP7_75t_L g2471 ( 
.A1(n_2436),
.A2(n_180),
.B1(n_178),
.B2(n_179),
.C(n_181),
.Y(n_2471)
);

OAI21xp5_ASAP7_75t_L g2472 ( 
.A1(n_2438),
.A2(n_180),
.B(n_182),
.Y(n_2472)
);

INVx1_ASAP7_75t_L g2473 ( 
.A(n_2427),
.Y(n_2473)
);

OAI221xp5_ASAP7_75t_L g2474 ( 
.A1(n_2447),
.A2(n_184),
.B1(n_182),
.B2(n_183),
.C(n_185),
.Y(n_2474)
);

INVx1_ASAP7_75t_L g2475 ( 
.A(n_2423),
.Y(n_2475)
);

AND2x4_ASAP7_75t_L g2476 ( 
.A(n_2425),
.B(n_2453),
.Y(n_2476)
);

INVx1_ASAP7_75t_L g2477 ( 
.A(n_2442),
.Y(n_2477)
);

INVx1_ASAP7_75t_L g2478 ( 
.A(n_2437),
.Y(n_2478)
);

INVxp67_ASAP7_75t_SL g2479 ( 
.A(n_2428),
.Y(n_2479)
);

INVx1_ASAP7_75t_L g2480 ( 
.A(n_2432),
.Y(n_2480)
);

NOR2xp67_ASAP7_75t_L g2481 ( 
.A(n_2452),
.B(n_183),
.Y(n_2481)
);

XNOR2xp5_ASAP7_75t_L g2482 ( 
.A(n_2433),
.B(n_184),
.Y(n_2482)
);

INVx1_ASAP7_75t_SL g2483 ( 
.A(n_2421),
.Y(n_2483)
);

XOR2xp5_ASAP7_75t_L g2484 ( 
.A(n_2434),
.B(n_185),
.Y(n_2484)
);

NOR2x1_ASAP7_75t_SL g2485 ( 
.A(n_2430),
.B(n_186),
.Y(n_2485)
);

INVxp67_ASAP7_75t_L g2486 ( 
.A(n_2439),
.Y(n_2486)
);

AOI221x1_ASAP7_75t_L g2487 ( 
.A1(n_2451),
.A2(n_188),
.B1(n_186),
.B2(n_187),
.C(n_189),
.Y(n_2487)
);

AOI22xp33_ASAP7_75t_L g2488 ( 
.A1(n_2440),
.A2(n_190),
.B1(n_188),
.B2(n_189),
.Y(n_2488)
);

NOR3xp33_ASAP7_75t_SL g2489 ( 
.A(n_2431),
.B(n_190),
.C(n_191),
.Y(n_2489)
);

OAI211xp5_ASAP7_75t_L g2490 ( 
.A1(n_2448),
.A2(n_193),
.B(n_191),
.C(n_192),
.Y(n_2490)
);

INVx2_ASAP7_75t_L g2491 ( 
.A(n_2427),
.Y(n_2491)
);

XNOR2xp5_ASAP7_75t_L g2492 ( 
.A(n_2419),
.B(n_193),
.Y(n_2492)
);

NOR2xp33_ASAP7_75t_L g2493 ( 
.A(n_2469),
.B(n_194),
.Y(n_2493)
);

NOR3x1_ASAP7_75t_L g2494 ( 
.A(n_2479),
.B(n_2474),
.C(n_2490),
.Y(n_2494)
);

NAND3xp33_ASAP7_75t_SL g2495 ( 
.A(n_2483),
.B(n_2463),
.C(n_2475),
.Y(n_2495)
);

AOI211x1_ASAP7_75t_L g2496 ( 
.A1(n_2457),
.A2(n_196),
.B(n_194),
.C(n_195),
.Y(n_2496)
);

NOR3xp33_ASAP7_75t_L g2497 ( 
.A(n_2477),
.B(n_195),
.C(n_197),
.Y(n_2497)
);

NAND4xp25_ASAP7_75t_L g2498 ( 
.A(n_2481),
.B(n_2487),
.C(n_2455),
.D(n_2464),
.Y(n_2498)
);

NAND2xp5_ASAP7_75t_L g2499 ( 
.A(n_2476),
.B(n_197),
.Y(n_2499)
);

AND2x2_ASAP7_75t_L g2500 ( 
.A(n_2466),
.B(n_198),
.Y(n_2500)
);

NOR3x1_ASAP7_75t_L g2501 ( 
.A(n_2468),
.B(n_198),
.C(n_199),
.Y(n_2501)
);

AND2x2_ASAP7_75t_L g2502 ( 
.A(n_2476),
.B(n_199),
.Y(n_2502)
);

INVx1_ASAP7_75t_L g2503 ( 
.A(n_2465),
.Y(n_2503)
);

NOR2xp67_ASAP7_75t_L g2504 ( 
.A(n_2467),
.B(n_200),
.Y(n_2504)
);

NAND2xp5_ASAP7_75t_L g2505 ( 
.A(n_2485),
.B(n_200),
.Y(n_2505)
);

NAND2xp5_ASAP7_75t_SL g2506 ( 
.A(n_2471),
.B(n_201),
.Y(n_2506)
);

AND2x2_ASAP7_75t_L g2507 ( 
.A(n_2478),
.B(n_202),
.Y(n_2507)
);

AOI21xp5_ASAP7_75t_L g2508 ( 
.A1(n_2492),
.A2(n_202),
.B(n_203),
.Y(n_2508)
);

NOR3xp33_ASAP7_75t_L g2509 ( 
.A(n_2480),
.B(n_204),
.C(n_205),
.Y(n_2509)
);

NAND4xp75_ASAP7_75t_L g2510 ( 
.A(n_2470),
.B(n_208),
.C(n_206),
.D(n_207),
.Y(n_2510)
);

NOR4xp25_ASAP7_75t_L g2511 ( 
.A(n_2473),
.B(n_2491),
.C(n_2486),
.D(n_2458),
.Y(n_2511)
);

NAND3xp33_ASAP7_75t_SL g2512 ( 
.A(n_2456),
.B(n_2459),
.C(n_2461),
.Y(n_2512)
);

NAND4xp75_ASAP7_75t_L g2513 ( 
.A(n_2472),
.B(n_2489),
.C(n_2460),
.D(n_2484),
.Y(n_2513)
);

NOR2x1_ASAP7_75t_L g2514 ( 
.A(n_2462),
.B(n_206),
.Y(n_2514)
);

NAND2xp5_ASAP7_75t_SL g2515 ( 
.A(n_2488),
.B(n_207),
.Y(n_2515)
);

INVx2_ASAP7_75t_SL g2516 ( 
.A(n_2482),
.Y(n_2516)
);

NAND3xp33_ASAP7_75t_L g2517 ( 
.A(n_2477),
.B(n_208),
.C(n_209),
.Y(n_2517)
);

NOR2x1_ASAP7_75t_L g2518 ( 
.A(n_2475),
.B(n_209),
.Y(n_2518)
);

NOR2x1_ASAP7_75t_L g2519 ( 
.A(n_2475),
.B(n_210),
.Y(n_2519)
);

NOR3xp33_ASAP7_75t_L g2520 ( 
.A(n_2483),
.B(n_210),
.C(n_211),
.Y(n_2520)
);

NAND2xp5_ASAP7_75t_L g2521 ( 
.A(n_2476),
.B(n_211),
.Y(n_2521)
);

NAND4xp75_ASAP7_75t_L g2522 ( 
.A(n_2469),
.B(n_215),
.C(n_212),
.D(n_213),
.Y(n_2522)
);

INVx1_ASAP7_75t_L g2523 ( 
.A(n_2465),
.Y(n_2523)
);

NAND2xp5_ASAP7_75t_L g2524 ( 
.A(n_2476),
.B(n_213),
.Y(n_2524)
);

NAND2xp5_ASAP7_75t_SL g2525 ( 
.A(n_2481),
.B(n_216),
.Y(n_2525)
);

NOR2x1_ASAP7_75t_L g2526 ( 
.A(n_2475),
.B(n_216),
.Y(n_2526)
);

INVx1_ASAP7_75t_L g2527 ( 
.A(n_2465),
.Y(n_2527)
);

NAND2xp5_ASAP7_75t_L g2528 ( 
.A(n_2476),
.B(n_217),
.Y(n_2528)
);

INVx1_ASAP7_75t_L g2529 ( 
.A(n_2465),
.Y(n_2529)
);

INVx1_ASAP7_75t_L g2530 ( 
.A(n_2465),
.Y(n_2530)
);

NAND4xp25_ASAP7_75t_L g2531 ( 
.A(n_2475),
.B(n_220),
.C(n_218),
.D(n_219),
.Y(n_2531)
);

NAND4xp75_ASAP7_75t_L g2532 ( 
.A(n_2469),
.B(n_221),
.C(n_219),
.D(n_220),
.Y(n_2532)
);

NAND4xp75_ASAP7_75t_L g2533 ( 
.A(n_2469),
.B(n_223),
.C(n_221),
.D(n_222),
.Y(n_2533)
);

AOI31xp33_ASAP7_75t_L g2534 ( 
.A1(n_2479),
.A2(n_224),
.A3(n_222),
.B(n_223),
.Y(n_2534)
);

AND5x1_ASAP7_75t_L g2535 ( 
.A(n_2456),
.B(n_226),
.C(n_224),
.D(n_225),
.E(n_227),
.Y(n_2535)
);

NAND3xp33_ASAP7_75t_L g2536 ( 
.A(n_2477),
.B(n_228),
.C(n_229),
.Y(n_2536)
);

NOR3xp33_ASAP7_75t_SL g2537 ( 
.A(n_2463),
.B(n_228),
.C(n_229),
.Y(n_2537)
);

NOR2xp33_ASAP7_75t_L g2538 ( 
.A(n_2469),
.B(n_230),
.Y(n_2538)
);

AOI211xp5_ASAP7_75t_L g2539 ( 
.A1(n_2457),
.A2(n_233),
.B(n_231),
.C(n_232),
.Y(n_2539)
);

NAND2xp5_ASAP7_75t_SL g2540 ( 
.A(n_2481),
.B(n_231),
.Y(n_2540)
);

NAND4xp75_ASAP7_75t_L g2541 ( 
.A(n_2469),
.B(n_234),
.C(n_232),
.D(n_233),
.Y(n_2541)
);

NOR3xp33_ASAP7_75t_L g2542 ( 
.A(n_2483),
.B(n_235),
.C(n_236),
.Y(n_2542)
);

NOR3xp33_ASAP7_75t_L g2543 ( 
.A(n_2483),
.B(n_235),
.C(n_237),
.Y(n_2543)
);

NAND2xp5_ASAP7_75t_L g2544 ( 
.A(n_2476),
.B(n_238),
.Y(n_2544)
);

INVx2_ASAP7_75t_L g2545 ( 
.A(n_2485),
.Y(n_2545)
);

NAND3x1_ASAP7_75t_L g2546 ( 
.A(n_2457),
.B(n_238),
.C(n_239),
.Y(n_2546)
);

OAI21xp5_ASAP7_75t_L g2547 ( 
.A1(n_2469),
.A2(n_239),
.B(n_240),
.Y(n_2547)
);

NOR3xp33_ASAP7_75t_L g2548 ( 
.A(n_2483),
.B(n_240),
.C(n_241),
.Y(n_2548)
);

INVx1_ASAP7_75t_L g2549 ( 
.A(n_2465),
.Y(n_2549)
);

NOR2x1p5_ASAP7_75t_L g2550 ( 
.A(n_2479),
.B(n_241),
.Y(n_2550)
);

NOR2x1_ASAP7_75t_L g2551 ( 
.A(n_2475),
.B(n_242),
.Y(n_2551)
);

NOR2x1_ASAP7_75t_L g2552 ( 
.A(n_2475),
.B(n_243),
.Y(n_2552)
);

O2A1O1Ixp33_ASAP7_75t_L g2553 ( 
.A1(n_2475),
.A2(n_245),
.B(n_243),
.C(n_244),
.Y(n_2553)
);

NAND4xp75_ASAP7_75t_L g2554 ( 
.A(n_2469),
.B(n_247),
.C(n_244),
.D(n_246),
.Y(n_2554)
);

NOR3xp33_ASAP7_75t_L g2555 ( 
.A(n_2495),
.B(n_248),
.C(n_249),
.Y(n_2555)
);

INVx1_ASAP7_75t_L g2556 ( 
.A(n_2518),
.Y(n_2556)
);

O2A1O1Ixp33_ASAP7_75t_SL g2557 ( 
.A1(n_2499),
.A2(n_250),
.B(n_248),
.C(n_249),
.Y(n_2557)
);

OAI21xp5_ASAP7_75t_L g2558 ( 
.A1(n_2493),
.A2(n_2538),
.B(n_2505),
.Y(n_2558)
);

NAND2xp33_ASAP7_75t_SL g2559 ( 
.A(n_2537),
.B(n_250),
.Y(n_2559)
);

CKINVDCx16_ASAP7_75t_R g2560 ( 
.A(n_2502),
.Y(n_2560)
);

AOI221xp5_ASAP7_75t_L g2561 ( 
.A1(n_2511),
.A2(n_253),
.B1(n_251),
.B2(n_252),
.C(n_254),
.Y(n_2561)
);

AND2x4_ASAP7_75t_L g2562 ( 
.A(n_2545),
.B(n_251),
.Y(n_2562)
);

XNOR2x1_ASAP7_75t_L g2563 ( 
.A(n_2513),
.B(n_252),
.Y(n_2563)
);

AOI21xp33_ASAP7_75t_SL g2564 ( 
.A1(n_2534),
.A2(n_253),
.B(n_254),
.Y(n_2564)
);

INVx1_ASAP7_75t_L g2565 ( 
.A(n_2519),
.Y(n_2565)
);

AND2x4_ASAP7_75t_L g2566 ( 
.A(n_2550),
.B(n_256),
.Y(n_2566)
);

NOR3xp33_ASAP7_75t_L g2567 ( 
.A(n_2503),
.B(n_257),
.C(n_258),
.Y(n_2567)
);

INVx1_ASAP7_75t_SL g2568 ( 
.A(n_2500),
.Y(n_2568)
);

OAI211xp5_ASAP7_75t_SL g2569 ( 
.A1(n_2523),
.A2(n_260),
.B(n_257),
.C(n_259),
.Y(n_2569)
);

NAND3xp33_ASAP7_75t_SL g2570 ( 
.A(n_2521),
.B(n_259),
.C(n_260),
.Y(n_2570)
);

AO22x2_ASAP7_75t_L g2571 ( 
.A1(n_2522),
.A2(n_263),
.B1(n_261),
.B2(n_262),
.Y(n_2571)
);

OAI221xp5_ASAP7_75t_L g2572 ( 
.A1(n_2527),
.A2(n_264),
.B1(n_261),
.B2(n_263),
.C(n_265),
.Y(n_2572)
);

NOR3x1_ASAP7_75t_L g2573 ( 
.A(n_2532),
.B(n_264),
.C(n_266),
.Y(n_2573)
);

AOI211xp5_ASAP7_75t_L g2574 ( 
.A1(n_2529),
.A2(n_2549),
.B(n_2530),
.C(n_2524),
.Y(n_2574)
);

AOI221xp5_ASAP7_75t_L g2575 ( 
.A1(n_2496),
.A2(n_268),
.B1(n_266),
.B2(n_267),
.C(n_269),
.Y(n_2575)
);

AOI21xp5_ASAP7_75t_L g2576 ( 
.A1(n_2528),
.A2(n_2544),
.B(n_2553),
.Y(n_2576)
);

OAI21xp33_ASAP7_75t_L g2577 ( 
.A1(n_2498),
.A2(n_267),
.B(n_269),
.Y(n_2577)
);

OAI22xp5_ASAP7_75t_SL g2578 ( 
.A1(n_2547),
.A2(n_274),
.B1(n_270),
.B2(n_272),
.Y(n_2578)
);

AND2x2_ASAP7_75t_L g2579 ( 
.A(n_2526),
.B(n_272),
.Y(n_2579)
);

OAI22xp33_ASAP7_75t_L g2580 ( 
.A1(n_2516),
.A2(n_276),
.B1(n_274),
.B2(n_275),
.Y(n_2580)
);

INVxp33_ASAP7_75t_SL g2581 ( 
.A(n_2494),
.Y(n_2581)
);

OAI22xp33_ASAP7_75t_L g2582 ( 
.A1(n_2517),
.A2(n_277),
.B1(n_275),
.B2(n_276),
.Y(n_2582)
);

AOI221xp5_ASAP7_75t_L g2583 ( 
.A1(n_2512),
.A2(n_282),
.B1(n_280),
.B2(n_281),
.C(n_283),
.Y(n_2583)
);

NAND4xp25_ASAP7_75t_L g2584 ( 
.A(n_2501),
.B(n_282),
.C(n_280),
.D(n_281),
.Y(n_2584)
);

INVx1_ASAP7_75t_L g2585 ( 
.A(n_2551),
.Y(n_2585)
);

AOI322xp5_ASAP7_75t_L g2586 ( 
.A1(n_2552),
.A2(n_284),
.A3(n_285),
.B1(n_286),
.B2(n_287),
.C1(n_289),
.C2(n_290),
.Y(n_2586)
);

INVx1_ASAP7_75t_L g2587 ( 
.A(n_2533),
.Y(n_2587)
);

OAI221xp5_ASAP7_75t_L g2588 ( 
.A1(n_2520),
.A2(n_291),
.B1(n_284),
.B2(n_286),
.C(n_292),
.Y(n_2588)
);

AOI211xp5_ASAP7_75t_L g2589 ( 
.A1(n_2542),
.A2(n_295),
.B(n_293),
.C(n_294),
.Y(n_2589)
);

AOI322xp5_ASAP7_75t_L g2590 ( 
.A1(n_2525),
.A2(n_294),
.A3(n_295),
.B1(n_296),
.B2(n_297),
.C1(n_298),
.C2(n_299),
.Y(n_2590)
);

OAI21xp33_ASAP7_75t_L g2591 ( 
.A1(n_2531),
.A2(n_296),
.B(n_300),
.Y(n_2591)
);

AND4x1_ASAP7_75t_L g2592 ( 
.A(n_2539),
.B(n_303),
.C(n_300),
.D(n_301),
.Y(n_2592)
);

NAND3xp33_ASAP7_75t_SL g2593 ( 
.A(n_2540),
.B(n_301),
.C(n_304),
.Y(n_2593)
);

NOR2x1_ASAP7_75t_L g2594 ( 
.A(n_2536),
.B(n_304),
.Y(n_2594)
);

INVx1_ASAP7_75t_L g2595 ( 
.A(n_2541),
.Y(n_2595)
);

AOI21xp5_ASAP7_75t_L g2596 ( 
.A1(n_2508),
.A2(n_305),
.B(n_306),
.Y(n_2596)
);

AOI22xp5_ASAP7_75t_L g2597 ( 
.A1(n_2504),
.A2(n_307),
.B1(n_305),
.B2(n_306),
.Y(n_2597)
);

XNOR2xp5_ASAP7_75t_L g2598 ( 
.A(n_2546),
.B(n_2554),
.Y(n_2598)
);

AND2x4_ASAP7_75t_L g2599 ( 
.A(n_2535),
.B(n_307),
.Y(n_2599)
);

INVx1_ASAP7_75t_L g2600 ( 
.A(n_2507),
.Y(n_2600)
);

NAND5xp2_ASAP7_75t_L g2601 ( 
.A(n_2543),
.B(n_310),
.C(n_308),
.D(n_309),
.E(n_311),
.Y(n_2601)
);

AOI21xp5_ASAP7_75t_L g2602 ( 
.A1(n_2506),
.A2(n_308),
.B(n_311),
.Y(n_2602)
);

AOI211x1_ASAP7_75t_L g2603 ( 
.A1(n_2515),
.A2(n_314),
.B(n_312),
.C(n_313),
.Y(n_2603)
);

AOI221xp5_ASAP7_75t_L g2604 ( 
.A1(n_2548),
.A2(n_315),
.B1(n_312),
.B2(n_313),
.C(n_316),
.Y(n_2604)
);

OAI311xp33_ASAP7_75t_L g2605 ( 
.A1(n_2514),
.A2(n_318),
.A3(n_315),
.B1(n_317),
.C1(n_319),
.Y(n_2605)
);

OAI21xp5_ASAP7_75t_L g2606 ( 
.A1(n_2510),
.A2(n_319),
.B(n_320),
.Y(n_2606)
);

NAND3xp33_ASAP7_75t_SL g2607 ( 
.A(n_2497),
.B(n_320),
.C(n_321),
.Y(n_2607)
);

NAND4xp25_ASAP7_75t_L g2608 ( 
.A(n_2539),
.B(n_323),
.C(n_321),
.D(n_322),
.Y(n_2608)
);

OAI22xp5_ASAP7_75t_L g2609 ( 
.A1(n_2509),
.A2(n_326),
.B1(n_323),
.B2(n_324),
.Y(n_2609)
);

NOR2x1_ASAP7_75t_L g2610 ( 
.A(n_2495),
.B(n_326),
.Y(n_2610)
);

AOI211xp5_ASAP7_75t_L g2611 ( 
.A1(n_2495),
.A2(n_329),
.B(n_327),
.C(n_328),
.Y(n_2611)
);

XNOR2xp5_ASAP7_75t_L g2612 ( 
.A(n_2513),
.B(n_327),
.Y(n_2612)
);

OR2x2_ASAP7_75t_L g2613 ( 
.A(n_2545),
.B(n_328),
.Y(n_2613)
);

AOI211xp5_ASAP7_75t_L g2614 ( 
.A1(n_2495),
.A2(n_331),
.B(n_329),
.C(n_330),
.Y(n_2614)
);

NAND2xp5_ASAP7_75t_L g2615 ( 
.A(n_2545),
.B(n_330),
.Y(n_2615)
);

AOI22xp5_ASAP7_75t_L g2616 ( 
.A1(n_2503),
.A2(n_333),
.B1(n_331),
.B2(n_332),
.Y(n_2616)
);

INVx2_ASAP7_75t_SL g2617 ( 
.A(n_2502),
.Y(n_2617)
);

AOI211xp5_ASAP7_75t_L g2618 ( 
.A1(n_2495),
.A2(n_334),
.B(n_332),
.C(n_333),
.Y(n_2618)
);

AOI311xp33_ASAP7_75t_L g2619 ( 
.A1(n_2503),
.A2(n_337),
.A3(n_335),
.B(n_336),
.C(n_338),
.Y(n_2619)
);

OAI22xp5_ASAP7_75t_L g2620 ( 
.A1(n_2499),
.A2(n_338),
.B1(n_335),
.B2(n_336),
.Y(n_2620)
);

OAI22xp5_ASAP7_75t_L g2621 ( 
.A1(n_2499),
.A2(n_341),
.B1(n_339),
.B2(n_340),
.Y(n_2621)
);

INVx2_ASAP7_75t_SL g2622 ( 
.A(n_2579),
.Y(n_2622)
);

INVx1_ASAP7_75t_L g2623 ( 
.A(n_2599),
.Y(n_2623)
);

INVx1_ASAP7_75t_L g2624 ( 
.A(n_2599),
.Y(n_2624)
);

INVx1_ASAP7_75t_L g2625 ( 
.A(n_2610),
.Y(n_2625)
);

NAND4xp75_ASAP7_75t_L g2626 ( 
.A(n_2556),
.B(n_341),
.C(n_339),
.D(n_340),
.Y(n_2626)
);

AOI22xp5_ASAP7_75t_L g2627 ( 
.A1(n_2581),
.A2(n_344),
.B1(n_342),
.B2(n_343),
.Y(n_2627)
);

NAND2xp5_ASAP7_75t_L g2628 ( 
.A(n_2560),
.B(n_342),
.Y(n_2628)
);

OR2x2_ASAP7_75t_L g2629 ( 
.A(n_2568),
.B(n_2565),
.Y(n_2629)
);

OAI22xp5_ASAP7_75t_L g2630 ( 
.A1(n_2611),
.A2(n_346),
.B1(n_343),
.B2(n_345),
.Y(n_2630)
);

OAI21x1_ASAP7_75t_SL g2631 ( 
.A1(n_2606),
.A2(n_346),
.B(n_347),
.Y(n_2631)
);

OA22x2_ASAP7_75t_L g2632 ( 
.A1(n_2597),
.A2(n_349),
.B1(n_347),
.B2(n_348),
.Y(n_2632)
);

NAND2xp5_ASAP7_75t_L g2633 ( 
.A(n_2585),
.B(n_348),
.Y(n_2633)
);

NAND4xp75_ASAP7_75t_L g2634 ( 
.A(n_2573),
.B(n_351),
.C(n_349),
.D(n_350),
.Y(n_2634)
);

NOR2xp33_ASAP7_75t_L g2635 ( 
.A(n_2566),
.B(n_350),
.Y(n_2635)
);

NAND2xp5_ASAP7_75t_SL g2636 ( 
.A(n_2566),
.B(n_351),
.Y(n_2636)
);

HB1xp67_ASAP7_75t_L g2637 ( 
.A(n_2562),
.Y(n_2637)
);

OAI31xp33_ASAP7_75t_L g2638 ( 
.A1(n_2605),
.A2(n_354),
.A3(n_352),
.B(n_353),
.Y(n_2638)
);

AOI211x1_ASAP7_75t_SL g2639 ( 
.A1(n_2558),
.A2(n_355),
.B(n_352),
.C(n_353),
.Y(n_2639)
);

OR2x2_ASAP7_75t_L g2640 ( 
.A(n_2584),
.B(n_355),
.Y(n_2640)
);

XNOR2xp5_ASAP7_75t_L g2641 ( 
.A(n_2563),
.B(n_356),
.Y(n_2641)
);

NAND4xp75_ASAP7_75t_L g2642 ( 
.A(n_2617),
.B(n_358),
.C(n_356),
.D(n_357),
.Y(n_2642)
);

A2O1A1Ixp33_ASAP7_75t_L g2643 ( 
.A1(n_2577),
.A2(n_359),
.B(n_357),
.C(n_358),
.Y(n_2643)
);

AND2x2_ASAP7_75t_L g2644 ( 
.A(n_2619),
.B(n_359),
.Y(n_2644)
);

AOI211x1_ASAP7_75t_L g2645 ( 
.A1(n_2591),
.A2(n_362),
.B(n_360),
.C(n_361),
.Y(n_2645)
);

O2A1O1Ixp33_ASAP7_75t_L g2646 ( 
.A1(n_2574),
.A2(n_363),
.B(n_360),
.C(n_362),
.Y(n_2646)
);

OR2x2_ASAP7_75t_L g2647 ( 
.A(n_2601),
.B(n_2613),
.Y(n_2647)
);

NAND4xp25_ASAP7_75t_L g2648 ( 
.A(n_2614),
.B(n_365),
.C(n_363),
.D(n_364),
.Y(n_2648)
);

OAI211xp5_ASAP7_75t_SL g2649 ( 
.A1(n_2561),
.A2(n_367),
.B(n_365),
.C(n_366),
.Y(n_2649)
);

OAI221xp5_ASAP7_75t_L g2650 ( 
.A1(n_2618),
.A2(n_366),
.B1(n_367),
.B2(n_368),
.C(n_369),
.Y(n_2650)
);

INVx1_ASAP7_75t_L g2651 ( 
.A(n_2571),
.Y(n_2651)
);

NAND2xp5_ASAP7_75t_L g2652 ( 
.A(n_2562),
.B(n_369),
.Y(n_2652)
);

NAND4xp25_ASAP7_75t_L g2653 ( 
.A(n_2559),
.B(n_372),
.C(n_370),
.D(n_371),
.Y(n_2653)
);

AND2x4_ASAP7_75t_L g2654 ( 
.A(n_2594),
.B(n_370),
.Y(n_2654)
);

INVx1_ASAP7_75t_L g2655 ( 
.A(n_2571),
.Y(n_2655)
);

AND3x4_ASAP7_75t_L g2656 ( 
.A(n_2592),
.B(n_372),
.C(n_373),
.Y(n_2656)
);

AOI221xp5_ASAP7_75t_SL g2657 ( 
.A1(n_2564),
.A2(n_374),
.B1(n_375),
.B2(n_376),
.C(n_377),
.Y(n_2657)
);

NOR2xp67_ASAP7_75t_L g2658 ( 
.A(n_2608),
.B(n_374),
.Y(n_2658)
);

NAND2xp5_ASAP7_75t_L g2659 ( 
.A(n_2600),
.B(n_376),
.Y(n_2659)
);

CKINVDCx5p33_ASAP7_75t_R g2660 ( 
.A(n_2612),
.Y(n_2660)
);

NAND4xp75_ASAP7_75t_L g2661 ( 
.A(n_2603),
.B(n_379),
.C(n_377),
.D(n_378),
.Y(n_2661)
);

NAND2xp5_ASAP7_75t_L g2662 ( 
.A(n_2598),
.B(n_379),
.Y(n_2662)
);

CKINVDCx16_ASAP7_75t_R g2663 ( 
.A(n_2587),
.Y(n_2663)
);

NAND2xp5_ASAP7_75t_SL g2664 ( 
.A(n_2575),
.B(n_380),
.Y(n_2664)
);

NAND3xp33_ASAP7_75t_SL g2665 ( 
.A(n_2555),
.B(n_381),
.C(n_382),
.Y(n_2665)
);

AND2x4_ASAP7_75t_L g2666 ( 
.A(n_2595),
.B(n_381),
.Y(n_2666)
);

NOR3xp33_ASAP7_75t_L g2667 ( 
.A(n_2570),
.B(n_384),
.C(n_385),
.Y(n_2667)
);

NOR3xp33_ASAP7_75t_L g2668 ( 
.A(n_2576),
.B(n_2593),
.C(n_2615),
.Y(n_2668)
);

NOR3xp33_ASAP7_75t_SL g2669 ( 
.A(n_2607),
.B(n_384),
.C(n_386),
.Y(n_2669)
);

INVx1_ASAP7_75t_L g2670 ( 
.A(n_2557),
.Y(n_2670)
);

CKINVDCx5p33_ASAP7_75t_R g2671 ( 
.A(n_2578),
.Y(n_2671)
);

INVx2_ASAP7_75t_SL g2672 ( 
.A(n_2620),
.Y(n_2672)
);

OAI22xp5_ASAP7_75t_L g2673 ( 
.A1(n_2588),
.A2(n_388),
.B1(n_386),
.B2(n_387),
.Y(n_2673)
);

AND3x1_ASAP7_75t_L g2674 ( 
.A(n_2567),
.B(n_387),
.C(n_389),
.Y(n_2674)
);

AOI221x1_ASAP7_75t_L g2675 ( 
.A1(n_2602),
.A2(n_389),
.B1(n_390),
.B2(n_391),
.C(n_392),
.Y(n_2675)
);

BUFx3_ASAP7_75t_L g2676 ( 
.A(n_2616),
.Y(n_2676)
);

INVx1_ASAP7_75t_L g2677 ( 
.A(n_2569),
.Y(n_2677)
);

NAND4xp75_ASAP7_75t_L g2678 ( 
.A(n_2596),
.B(n_393),
.C(n_390),
.D(n_392),
.Y(n_2678)
);

NOR2xp33_ASAP7_75t_L g2679 ( 
.A(n_2621),
.B(n_393),
.Y(n_2679)
);

CKINVDCx5p33_ASAP7_75t_R g2680 ( 
.A(n_2609),
.Y(n_2680)
);

INVx1_ASAP7_75t_L g2681 ( 
.A(n_2589),
.Y(n_2681)
);

NOR2x1_ASAP7_75t_L g2682 ( 
.A(n_2580),
.B(n_394),
.Y(n_2682)
);

INVx1_ASAP7_75t_SL g2683 ( 
.A(n_2586),
.Y(n_2683)
);

AND2x4_ASAP7_75t_SL g2684 ( 
.A(n_2590),
.B(n_394),
.Y(n_2684)
);

INVx1_ASAP7_75t_L g2685 ( 
.A(n_2582),
.Y(n_2685)
);

NAND4xp25_ASAP7_75t_L g2686 ( 
.A(n_2604),
.B(n_397),
.C(n_395),
.D(n_396),
.Y(n_2686)
);

OAI211xp5_ASAP7_75t_L g2687 ( 
.A1(n_2629),
.A2(n_2583),
.B(n_2572),
.C(n_397),
.Y(n_2687)
);

INVx1_ASAP7_75t_L g2688 ( 
.A(n_2637),
.Y(n_2688)
);

AOI22xp5_ASAP7_75t_L g2689 ( 
.A1(n_2663),
.A2(n_398),
.B1(n_395),
.B2(n_396),
.Y(n_2689)
);

OAI311xp33_ASAP7_75t_L g2690 ( 
.A1(n_2623),
.A2(n_399),
.A3(n_400),
.B1(n_401),
.C1(n_402),
.Y(n_2690)
);

NAND5xp2_ASAP7_75t_L g2691 ( 
.A(n_2624),
.B(n_401),
.C(n_402),
.D(n_403),
.E(n_404),
.Y(n_2691)
);

NAND4xp25_ASAP7_75t_L g2692 ( 
.A(n_2639),
.B(n_407),
.C(n_404),
.D(n_405),
.Y(n_2692)
);

NAND5xp2_ASAP7_75t_L g2693 ( 
.A(n_2638),
.B(n_405),
.C(n_408),
.D(n_409),
.E(n_410),
.Y(n_2693)
);

AOI311xp33_ASAP7_75t_L g2694 ( 
.A1(n_2651),
.A2(n_408),
.A3(n_409),
.B(n_410),
.C(n_411),
.Y(n_2694)
);

OAI22xp5_ASAP7_75t_L g2695 ( 
.A1(n_2627),
.A2(n_415),
.B1(n_412),
.B2(n_414),
.Y(n_2695)
);

OAI22xp5_ASAP7_75t_L g2696 ( 
.A1(n_2662),
.A2(n_417),
.B1(n_415),
.B2(n_416),
.Y(n_2696)
);

AND2x2_ASAP7_75t_L g2697 ( 
.A(n_2644),
.B(n_2625),
.Y(n_2697)
);

NAND5xp2_ASAP7_75t_L g2698 ( 
.A(n_2668),
.B(n_416),
.C(n_417),
.D(n_418),
.E(n_419),
.Y(n_2698)
);

XNOR2xp5_ASAP7_75t_L g2699 ( 
.A(n_2641),
.B(n_419),
.Y(n_2699)
);

A2O1A1Ixp33_ASAP7_75t_L g2700 ( 
.A1(n_2646),
.A2(n_423),
.B(n_420),
.C(n_422),
.Y(n_2700)
);

INVx1_ASAP7_75t_L g2701 ( 
.A(n_2656),
.Y(n_2701)
);

INVx1_ASAP7_75t_L g2702 ( 
.A(n_2647),
.Y(n_2702)
);

INVx1_ASAP7_75t_L g2703 ( 
.A(n_2652),
.Y(n_2703)
);

AOI22xp5_ASAP7_75t_L g2704 ( 
.A1(n_2660),
.A2(n_2683),
.B1(n_2622),
.B2(n_2628),
.Y(n_2704)
);

INVx2_ASAP7_75t_SL g2705 ( 
.A(n_2654),
.Y(n_2705)
);

AND3x1_ASAP7_75t_L g2706 ( 
.A(n_2635),
.B(n_422),
.C(n_424),
.Y(n_2706)
);

NOR3xp33_ASAP7_75t_L g2707 ( 
.A(n_2655),
.B(n_424),
.C(n_425),
.Y(n_2707)
);

NOR3xp33_ASAP7_75t_SL g2708 ( 
.A(n_2671),
.B(n_425),
.C(n_426),
.Y(n_2708)
);

AND4x1_ASAP7_75t_L g2709 ( 
.A(n_2669),
.B(n_427),
.C(n_428),
.D(n_429),
.Y(n_2709)
);

HB1xp67_ASAP7_75t_L g2710 ( 
.A(n_2654),
.Y(n_2710)
);

OAI21xp5_ASAP7_75t_L g2711 ( 
.A1(n_2658),
.A2(n_428),
.B(n_430),
.Y(n_2711)
);

AOI22xp33_ASAP7_75t_SL g2712 ( 
.A1(n_2670),
.A2(n_431),
.B1(n_432),
.B2(n_434),
.Y(n_2712)
);

XOR2xp5_ASAP7_75t_L g2713 ( 
.A(n_2634),
.B(n_431),
.Y(n_2713)
);

AOI22xp5_ASAP7_75t_L g2714 ( 
.A1(n_2665),
.A2(n_432),
.B1(n_434),
.B2(n_435),
.Y(n_2714)
);

OR2x2_ASAP7_75t_L g2715 ( 
.A(n_2653),
.B(n_435),
.Y(n_2715)
);

INVx1_ASAP7_75t_L g2716 ( 
.A(n_2666),
.Y(n_2716)
);

NAND3xp33_ASAP7_75t_L g2717 ( 
.A(n_2636),
.B(n_2680),
.C(n_2659),
.Y(n_2717)
);

INVx1_ASAP7_75t_L g2718 ( 
.A(n_2666),
.Y(n_2718)
);

NOR2xp33_ASAP7_75t_L g2719 ( 
.A(n_2677),
.B(n_436),
.Y(n_2719)
);

NAND5xp2_ASAP7_75t_L g2720 ( 
.A(n_2657),
.B(n_436),
.C(n_437),
.D(n_438),
.E(n_439),
.Y(n_2720)
);

NOR3xp33_ASAP7_75t_L g2721 ( 
.A(n_2672),
.B(n_437),
.C(n_438),
.Y(n_2721)
);

AOI22xp5_ASAP7_75t_L g2722 ( 
.A1(n_2630),
.A2(n_439),
.B1(n_440),
.B2(n_441),
.Y(n_2722)
);

AOI22xp33_ASAP7_75t_L g2723 ( 
.A1(n_2667),
.A2(n_2632),
.B1(n_2676),
.B2(n_2682),
.Y(n_2723)
);

AOI211xp5_ASAP7_75t_L g2724 ( 
.A1(n_2640),
.A2(n_440),
.B(n_441),
.C(n_442),
.Y(n_2724)
);

NOR4xp25_ASAP7_75t_L g2725 ( 
.A(n_2685),
.B(n_443),
.C(n_444),
.D(n_445),
.Y(n_2725)
);

NAND3xp33_ASAP7_75t_L g2726 ( 
.A(n_2681),
.B(n_443),
.C(n_444),
.Y(n_2726)
);

HB1xp67_ASAP7_75t_L g2727 ( 
.A(n_2674),
.Y(n_2727)
);

AOI211x1_ASAP7_75t_L g2728 ( 
.A1(n_2664),
.A2(n_2650),
.B(n_2648),
.C(n_2686),
.Y(n_2728)
);

OAI221xp5_ASAP7_75t_L g2729 ( 
.A1(n_2643),
.A2(n_446),
.B1(n_447),
.B2(n_448),
.C(n_449),
.Y(n_2729)
);

INVx2_ASAP7_75t_L g2730 ( 
.A(n_2661),
.Y(n_2730)
);

INVx1_ASAP7_75t_L g2731 ( 
.A(n_2633),
.Y(n_2731)
);

BUFx2_ASAP7_75t_L g2732 ( 
.A(n_2710),
.Y(n_2732)
);

XNOR2x1_ASAP7_75t_L g2733 ( 
.A(n_2688),
.B(n_2678),
.Y(n_2733)
);

NOR4xp25_ASAP7_75t_L g2734 ( 
.A(n_2705),
.B(n_2649),
.C(n_2679),
.D(n_2673),
.Y(n_2734)
);

INVx2_ASAP7_75t_L g2735 ( 
.A(n_2697),
.Y(n_2735)
);

AOI222xp33_ASAP7_75t_L g2736 ( 
.A1(n_2702),
.A2(n_2684),
.B1(n_2631),
.B2(n_2645),
.C1(n_2675),
.C2(n_2642),
.Y(n_2736)
);

INVxp33_ASAP7_75t_L g2737 ( 
.A(n_2699),
.Y(n_2737)
);

AND2x4_ASAP7_75t_L g2738 ( 
.A(n_2716),
.B(n_2626),
.Y(n_2738)
);

NOR2xp33_ASAP7_75t_L g2739 ( 
.A(n_2718),
.B(n_446),
.Y(n_2739)
);

NAND4xp75_ASAP7_75t_L g2740 ( 
.A(n_2704),
.B(n_447),
.C(n_448),
.D(n_450),
.Y(n_2740)
);

INVx1_ASAP7_75t_L g2741 ( 
.A(n_2727),
.Y(n_2741)
);

AOI21xp5_ASAP7_75t_L g2742 ( 
.A1(n_2701),
.A2(n_451),
.B(n_452),
.Y(n_2742)
);

INVx1_ASAP7_75t_L g2743 ( 
.A(n_2706),
.Y(n_2743)
);

HB1xp67_ASAP7_75t_L g2744 ( 
.A(n_2709),
.Y(n_2744)
);

XNOR2xp5_ASAP7_75t_L g2745 ( 
.A(n_2717),
.B(n_2713),
.Y(n_2745)
);

AOI21xp5_ASAP7_75t_L g2746 ( 
.A1(n_2711),
.A2(n_451),
.B(n_452),
.Y(n_2746)
);

INVx2_ASAP7_75t_L g2747 ( 
.A(n_2715),
.Y(n_2747)
);

NOR4xp25_ASAP7_75t_L g2748 ( 
.A(n_2703),
.B(n_453),
.C(n_454),
.D(n_455),
.Y(n_2748)
);

NAND2xp5_ASAP7_75t_L g2749 ( 
.A(n_2731),
.B(n_453),
.Y(n_2749)
);

AOI22xp5_ASAP7_75t_L g2750 ( 
.A1(n_2721),
.A2(n_2707),
.B1(n_2730),
.B2(n_2696),
.Y(n_2750)
);

NAND4xp75_ASAP7_75t_L g2751 ( 
.A(n_2708),
.B(n_456),
.C(n_457),
.D(n_458),
.Y(n_2751)
);

AOI22xp5_ASAP7_75t_L g2752 ( 
.A1(n_2695),
.A2(n_456),
.B1(n_458),
.B2(n_459),
.Y(n_2752)
);

OAI211xp5_ASAP7_75t_SL g2753 ( 
.A1(n_2723),
.A2(n_460),
.B(n_461),
.C(n_462),
.Y(n_2753)
);

HB1xp67_ASAP7_75t_L g2754 ( 
.A(n_2719),
.Y(n_2754)
);

NOR2xp33_ASAP7_75t_L g2755 ( 
.A(n_2691),
.B(n_2698),
.Y(n_2755)
);

INVx1_ASAP7_75t_L g2756 ( 
.A(n_2720),
.Y(n_2756)
);

NAND2xp5_ASAP7_75t_L g2757 ( 
.A(n_2728),
.B(n_460),
.Y(n_2757)
);

INVx1_ASAP7_75t_L g2758 ( 
.A(n_2693),
.Y(n_2758)
);

AOI22xp5_ASAP7_75t_L g2759 ( 
.A1(n_2687),
.A2(n_462),
.B1(n_463),
.B2(n_464),
.Y(n_2759)
);

INVxp67_ASAP7_75t_L g2760 ( 
.A(n_2726),
.Y(n_2760)
);

AO22x1_ASAP7_75t_L g2761 ( 
.A1(n_2694),
.A2(n_463),
.B1(n_464),
.B2(n_465),
.Y(n_2761)
);

NAND4xp25_ASAP7_75t_L g2762 ( 
.A(n_2692),
.B(n_2724),
.C(n_2714),
.D(n_2722),
.Y(n_2762)
);

INVx1_ASAP7_75t_SL g2763 ( 
.A(n_2712),
.Y(n_2763)
);

INVx2_ASAP7_75t_L g2764 ( 
.A(n_2689),
.Y(n_2764)
);

INVx1_ASAP7_75t_SL g2765 ( 
.A(n_2725),
.Y(n_2765)
);

INVx2_ASAP7_75t_L g2766 ( 
.A(n_2729),
.Y(n_2766)
);

OAI211xp5_ASAP7_75t_L g2767 ( 
.A1(n_2724),
.A2(n_466),
.B(n_467),
.C(n_468),
.Y(n_2767)
);

NAND2xp5_ASAP7_75t_L g2768 ( 
.A(n_2732),
.B(n_2700),
.Y(n_2768)
);

NOR2x1p5_ASAP7_75t_L g2769 ( 
.A(n_2751),
.B(n_2690),
.Y(n_2769)
);

NAND2xp5_ASAP7_75t_L g2770 ( 
.A(n_2735),
.B(n_466),
.Y(n_2770)
);

AOI221xp5_ASAP7_75t_SL g2771 ( 
.A1(n_2741),
.A2(n_469),
.B1(n_471),
.B2(n_472),
.C(n_473),
.Y(n_2771)
);

A2O1A1Ixp33_ASAP7_75t_SL g2772 ( 
.A1(n_2747),
.A2(n_469),
.B(n_472),
.C(n_473),
.Y(n_2772)
);

OR4x2_ASAP7_75t_L g2773 ( 
.A(n_2736),
.B(n_474),
.C(n_475),
.D(n_476),
.Y(n_2773)
);

AOI21xp5_ASAP7_75t_L g2774 ( 
.A1(n_2757),
.A2(n_474),
.B(n_475),
.Y(n_2774)
);

OR2x2_ASAP7_75t_L g2775 ( 
.A(n_2758),
.B(n_477),
.Y(n_2775)
);

AND2x2_ASAP7_75t_L g2776 ( 
.A(n_2756),
.B(n_477),
.Y(n_2776)
);

AO22x2_ASAP7_75t_L g2777 ( 
.A1(n_2733),
.A2(n_478),
.B1(n_479),
.B2(n_480),
.Y(n_2777)
);

OAI22x1_ASAP7_75t_L g2778 ( 
.A1(n_2759),
.A2(n_2765),
.B1(n_2743),
.B2(n_2744),
.Y(n_2778)
);

HB1xp67_ASAP7_75t_L g2779 ( 
.A(n_2755),
.Y(n_2779)
);

INVx1_ASAP7_75t_L g2780 ( 
.A(n_2754),
.Y(n_2780)
);

INVx1_ASAP7_75t_L g2781 ( 
.A(n_2745),
.Y(n_2781)
);

NAND2xp5_ASAP7_75t_L g2782 ( 
.A(n_2737),
.B(n_478),
.Y(n_2782)
);

INVx2_ASAP7_75t_L g2783 ( 
.A(n_2740),
.Y(n_2783)
);

OAI22x1_ASAP7_75t_L g2784 ( 
.A1(n_2750),
.A2(n_479),
.B1(n_480),
.B2(n_481),
.Y(n_2784)
);

NOR3xp33_ASAP7_75t_L g2785 ( 
.A(n_2738),
.B(n_482),
.C(n_483),
.Y(n_2785)
);

NOR3xp33_ASAP7_75t_L g2786 ( 
.A(n_2738),
.B(n_482),
.C(n_483),
.Y(n_2786)
);

XNOR2xp5_ASAP7_75t_L g2787 ( 
.A(n_2734),
.B(n_484),
.Y(n_2787)
);

AOI21xp5_ASAP7_75t_L g2788 ( 
.A1(n_2763),
.A2(n_485),
.B(n_486),
.Y(n_2788)
);

OAI22xp5_ASAP7_75t_L g2789 ( 
.A1(n_2752),
.A2(n_485),
.B1(n_486),
.B2(n_487),
.Y(n_2789)
);

INVx1_ASAP7_75t_L g2790 ( 
.A(n_2749),
.Y(n_2790)
);

INVx4_ASAP7_75t_L g2791 ( 
.A(n_2764),
.Y(n_2791)
);

INVx1_ASAP7_75t_L g2792 ( 
.A(n_2739),
.Y(n_2792)
);

NOR2x2_ASAP7_75t_L g2793 ( 
.A(n_2766),
.B(n_487),
.Y(n_2793)
);

AND2x2_ASAP7_75t_L g2794 ( 
.A(n_2748),
.B(n_488),
.Y(n_2794)
);

INVx3_ASAP7_75t_L g2795 ( 
.A(n_2791),
.Y(n_2795)
);

AOI22xp5_ASAP7_75t_L g2796 ( 
.A1(n_2780),
.A2(n_2753),
.B1(n_2760),
.B2(n_2762),
.Y(n_2796)
);

XNOR2xp5_ASAP7_75t_L g2797 ( 
.A(n_2779),
.B(n_2761),
.Y(n_2797)
);

INVx2_ASAP7_75t_L g2798 ( 
.A(n_2793),
.Y(n_2798)
);

AO22x2_ASAP7_75t_L g2799 ( 
.A1(n_2775),
.A2(n_2767),
.B1(n_2746),
.B2(n_2742),
.Y(n_2799)
);

NOR3xp33_ASAP7_75t_L g2800 ( 
.A(n_2781),
.B(n_2790),
.C(n_2768),
.Y(n_2800)
);

INVx1_ASAP7_75t_L g2801 ( 
.A(n_2787),
.Y(n_2801)
);

AOI22xp5_ASAP7_75t_L g2802 ( 
.A1(n_2769),
.A2(n_488),
.B1(n_489),
.B2(n_490),
.Y(n_2802)
);

AND2x4_ASAP7_75t_L g2803 ( 
.A(n_2792),
.B(n_489),
.Y(n_2803)
);

OAI22xp33_ASAP7_75t_SL g2804 ( 
.A1(n_2770),
.A2(n_490),
.B1(n_491),
.B2(n_492),
.Y(n_2804)
);

NAND2xp5_ASAP7_75t_SL g2805 ( 
.A(n_2776),
.B(n_491),
.Y(n_2805)
);

INVx1_ASAP7_75t_L g2806 ( 
.A(n_2773),
.Y(n_2806)
);

XOR2x1_ASAP7_75t_L g2807 ( 
.A(n_2794),
.B(n_492),
.Y(n_2807)
);

OAI22xp5_ASAP7_75t_SL g2808 ( 
.A1(n_2783),
.A2(n_493),
.B1(n_494),
.B2(n_495),
.Y(n_2808)
);

INVx2_ASAP7_75t_L g2809 ( 
.A(n_2777),
.Y(n_2809)
);

INVx3_ASAP7_75t_L g2810 ( 
.A(n_2777),
.Y(n_2810)
);

INVx1_ASAP7_75t_L g2811 ( 
.A(n_2782),
.Y(n_2811)
);

AOI22xp5_ASAP7_75t_L g2812 ( 
.A1(n_2778),
.A2(n_493),
.B1(n_494),
.B2(n_495),
.Y(n_2812)
);

INVx4_ASAP7_75t_L g2813 ( 
.A(n_2774),
.Y(n_2813)
);

INVx2_ASAP7_75t_SL g2814 ( 
.A(n_2784),
.Y(n_2814)
);

INVx1_ASAP7_75t_L g2815 ( 
.A(n_2795),
.Y(n_2815)
);

INVx1_ASAP7_75t_L g2816 ( 
.A(n_2798),
.Y(n_2816)
);

INVx2_ASAP7_75t_L g2817 ( 
.A(n_2806),
.Y(n_2817)
);

AOI22xp33_ASAP7_75t_SL g2818 ( 
.A1(n_2810),
.A2(n_2789),
.B1(n_2788),
.B2(n_2772),
.Y(n_2818)
);

AND3x4_ASAP7_75t_L g2819 ( 
.A(n_2800),
.B(n_2786),
.C(n_2785),
.Y(n_2819)
);

NOR3xp33_ASAP7_75t_L g2820 ( 
.A(n_2801),
.B(n_2811),
.C(n_2813),
.Y(n_2820)
);

NAND4xp25_ASAP7_75t_L g2821 ( 
.A(n_2796),
.B(n_2771),
.C(n_498),
.D(n_499),
.Y(n_2821)
);

INVx1_ASAP7_75t_L g2822 ( 
.A(n_2797),
.Y(n_2822)
);

AOI221xp5_ASAP7_75t_SL g2823 ( 
.A1(n_2809),
.A2(n_496),
.B1(n_499),
.B2(n_500),
.C(n_501),
.Y(n_2823)
);

OAI321xp33_ASAP7_75t_L g2824 ( 
.A1(n_2814),
.A2(n_496),
.A3(n_500),
.B1(n_501),
.B2(n_502),
.C(n_503),
.Y(n_2824)
);

INVx1_ASAP7_75t_L g2825 ( 
.A(n_2807),
.Y(n_2825)
);

NOR3xp33_ASAP7_75t_SL g2826 ( 
.A(n_2805),
.B(n_502),
.C(n_504),
.Y(n_2826)
);

OAI221xp5_ASAP7_75t_L g2827 ( 
.A1(n_2812),
.A2(n_504),
.B1(n_505),
.B2(n_506),
.C(n_507),
.Y(n_2827)
);

AOI22xp5_ASAP7_75t_L g2828 ( 
.A1(n_2817),
.A2(n_2799),
.B1(n_2804),
.B2(n_2802),
.Y(n_2828)
);

INVx1_ASAP7_75t_L g2829 ( 
.A(n_2816),
.Y(n_2829)
);

NAND2xp5_ASAP7_75t_L g2830 ( 
.A(n_2825),
.B(n_2803),
.Y(n_2830)
);

HB1xp67_ASAP7_75t_L g2831 ( 
.A(n_2815),
.Y(n_2831)
);

INVx1_ASAP7_75t_L g2832 ( 
.A(n_2822),
.Y(n_2832)
);

INVx1_ASAP7_75t_L g2833 ( 
.A(n_2820),
.Y(n_2833)
);

XOR2xp5_ASAP7_75t_L g2834 ( 
.A(n_2818),
.B(n_2808),
.Y(n_2834)
);

OAI22xp5_ASAP7_75t_L g2835 ( 
.A1(n_2819),
.A2(n_506),
.B1(n_508),
.B2(n_509),
.Y(n_2835)
);

HB1xp67_ASAP7_75t_L g2836 ( 
.A(n_2821),
.Y(n_2836)
);

HB1xp67_ASAP7_75t_L g2837 ( 
.A(n_2831),
.Y(n_2837)
);

INVx1_ASAP7_75t_L g2838 ( 
.A(n_2832),
.Y(n_2838)
);

OAI22x1_ASAP7_75t_L g2839 ( 
.A1(n_2829),
.A2(n_2826),
.B1(n_2823),
.B2(n_2824),
.Y(n_2839)
);

HB1xp67_ASAP7_75t_L g2840 ( 
.A(n_2833),
.Y(n_2840)
);

NOR2x1_ASAP7_75t_L g2841 ( 
.A(n_2830),
.B(n_2827),
.Y(n_2841)
);

INVx1_ASAP7_75t_L g2842 ( 
.A(n_2834),
.Y(n_2842)
);

AOI222xp33_ASAP7_75t_SL g2843 ( 
.A1(n_2837),
.A2(n_2838),
.B1(n_2840),
.B2(n_2842),
.C1(n_2836),
.C2(n_2828),
.Y(n_2843)
);

AOI221xp5_ASAP7_75t_L g2844 ( 
.A1(n_2839),
.A2(n_2835),
.B1(n_509),
.B2(n_510),
.C(n_511),
.Y(n_2844)
);

NAND2xp5_ASAP7_75t_L g2845 ( 
.A(n_2841),
.B(n_508),
.Y(n_2845)
);

XNOR2xp5_ASAP7_75t_L g2846 ( 
.A(n_2837),
.B(n_510),
.Y(n_2846)
);

BUFx2_ASAP7_75t_L g2847 ( 
.A(n_2845),
.Y(n_2847)
);

AOI222xp33_ASAP7_75t_L g2848 ( 
.A1(n_2844),
.A2(n_511),
.B1(n_512),
.B2(n_513),
.C1(n_514),
.C2(n_516),
.Y(n_2848)
);

AND2x2_ASAP7_75t_SL g2849 ( 
.A(n_2843),
.B(n_513),
.Y(n_2849)
);

OR2x2_ASAP7_75t_L g2850 ( 
.A(n_2847),
.B(n_2846),
.Y(n_2850)
);

AO21x2_ASAP7_75t_L g2851 ( 
.A1(n_2849),
.A2(n_516),
.B(n_517),
.Y(n_2851)
);

AOI22xp33_ASAP7_75t_L g2852 ( 
.A1(n_2848),
.A2(n_517),
.B1(n_518),
.B2(n_519),
.Y(n_2852)
);

AOI22xp5_ASAP7_75t_L g2853 ( 
.A1(n_2849),
.A2(n_518),
.B1(n_519),
.B2(n_520),
.Y(n_2853)
);

BUFx2_ASAP7_75t_L g2854 ( 
.A(n_2850),
.Y(n_2854)
);

INVx1_ASAP7_75t_L g2855 ( 
.A(n_2851),
.Y(n_2855)
);

OR2x6_ASAP7_75t_L g2856 ( 
.A(n_2854),
.B(n_2853),
.Y(n_2856)
);

AOI221xp5_ASAP7_75t_L g2857 ( 
.A1(n_2856),
.A2(n_2855),
.B1(n_2852),
.B2(n_523),
.C(n_524),
.Y(n_2857)
);

AOI211xp5_ASAP7_75t_L g2858 ( 
.A1(n_2857),
.A2(n_521),
.B(n_522),
.C(n_523),
.Y(n_2858)
);


endmodule