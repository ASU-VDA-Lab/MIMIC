module fake_jpeg_19826_n_228 (n_3, n_2, n_1, n_0, n_10, n_4, n_8, n_9, n_6, n_5, n_7, n_228);

input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_228;

wire n_159;
wire n_117;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_14;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_13;
wire n_175;
wire n_187;
wire n_57;
wire n_21;
wire n_223;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_24;
wire n_44;
wire n_143;
wire n_202;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_121;
wire n_130;
wire n_99;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_11;
wire n_131;
wire n_56;
wire n_212;
wire n_211;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_12;
wire n_132;
wire n_133;
wire n_67;
wire n_216;
wire n_217;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

BUFx6f_ASAP7_75t_L g11 ( 
.A(n_4),
.Y(n_11)
);

CKINVDCx20_ASAP7_75t_R g12 ( 
.A(n_2),
.Y(n_12)
);

BUFx4f_ASAP7_75t_SL g13 ( 
.A(n_10),
.Y(n_13)
);

BUFx6f_ASAP7_75t_L g14 ( 
.A(n_4),
.Y(n_14)
);

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_1),
.Y(n_15)
);

BUFx12f_ASAP7_75t_L g16 ( 
.A(n_10),
.Y(n_16)
);

INVx1_ASAP7_75t_SL g17 ( 
.A(n_10),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_0),
.Y(n_18)
);

INVx2_ASAP7_75t_L g19 ( 
.A(n_4),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_8),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_0),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_4),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_6),
.Y(n_23)
);

INVx8_ASAP7_75t_L g24 ( 
.A(n_16),
.Y(n_24)
);

INVx5_ASAP7_75t_L g35 ( 
.A(n_24),
.Y(n_35)
);

AOI21xp33_ASAP7_75t_L g25 ( 
.A1(n_12),
.A2(n_0),
.B(n_1),
.Y(n_25)
);

NOR2xp33_ASAP7_75t_L g37 ( 
.A(n_25),
.B(n_27),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_11),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_26),
.Y(n_36)
);

NAND2xp5_ASAP7_75t_SL g27 ( 
.A(n_16),
.B(n_9),
.Y(n_27)
);

INVx5_ASAP7_75t_L g28 ( 
.A(n_16),
.Y(n_28)
);

INVx4_ASAP7_75t_L g40 ( 
.A(n_28),
.Y(n_40)
);

BUFx5_ASAP7_75t_L g29 ( 
.A(n_11),
.Y(n_29)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_29),
.Y(n_39)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_13),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_30),
.Y(n_41)
);

INVx3_ASAP7_75t_L g31 ( 
.A(n_16),
.Y(n_31)
);

OA22x2_ASAP7_75t_L g38 ( 
.A1(n_31),
.A2(n_32),
.B1(n_17),
.B2(n_19),
.Y(n_38)
);

INVx4_ASAP7_75t_L g32 ( 
.A(n_16),
.Y(n_32)
);

AOI22xp33_ASAP7_75t_L g33 ( 
.A1(n_27),
.A2(n_19),
.B1(n_17),
.B2(n_22),
.Y(n_33)
);

AOI22xp5_ASAP7_75t_L g42 ( 
.A1(n_33),
.A2(n_27),
.B1(n_30),
.B2(n_32),
.Y(n_42)
);

AND2x2_ASAP7_75t_SL g34 ( 
.A(n_32),
.B(n_17),
.Y(n_34)
);

NAND2xp5_ASAP7_75t_SL g51 ( 
.A(n_34),
.B(n_30),
.Y(n_51)
);

AND2x2_ASAP7_75t_L g52 ( 
.A(n_38),
.B(n_32),
.Y(n_52)
);

OAI22xp5_ASAP7_75t_SL g64 ( 
.A1(n_42),
.A2(n_24),
.B1(n_28),
.B2(n_31),
.Y(n_64)
);

INVx6_ASAP7_75t_L g43 ( 
.A(n_35),
.Y(n_43)
);

AOI22xp33_ASAP7_75t_SL g71 ( 
.A1(n_43),
.A2(n_53),
.B1(n_54),
.B2(n_55),
.Y(n_71)
);

INVx3_ASAP7_75t_L g44 ( 
.A(n_40),
.Y(n_44)
);

INVx2_ASAP7_75t_L g78 ( 
.A(n_44),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_L g45 ( 
.A(n_37),
.B(n_26),
.Y(n_45)
);

NAND2xp5_ASAP7_75t_L g68 ( 
.A(n_45),
.B(n_51),
.Y(n_68)
);

OAI22xp5_ASAP7_75t_L g46 ( 
.A1(n_37),
.A2(n_19),
.B1(n_32),
.B2(n_30),
.Y(n_46)
);

AOI22xp5_ASAP7_75t_L g70 ( 
.A1(n_46),
.A2(n_59),
.B1(n_34),
.B2(n_39),
.Y(n_70)
);

INVx2_ASAP7_75t_L g47 ( 
.A(n_36),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_47),
.B(n_48),
.Y(n_72)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_39),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_36),
.Y(n_49)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_49),
.Y(n_65)
);

XOR2xp5_ASAP7_75t_SL g50 ( 
.A(n_34),
.B(n_33),
.Y(n_50)
);

A2O1A1Ixp33_ASAP7_75t_L g60 ( 
.A1(n_50),
.A2(n_45),
.B(n_34),
.C(n_51),
.Y(n_60)
);

AOI22xp5_ASAP7_75t_L g74 ( 
.A1(n_52),
.A2(n_34),
.B1(n_24),
.B2(n_31),
.Y(n_74)
);

INVx8_ASAP7_75t_L g53 ( 
.A(n_36),
.Y(n_53)
);

INVx5_ASAP7_75t_L g54 ( 
.A(n_36),
.Y(n_54)
);

AOI22xp33_ASAP7_75t_SL g55 ( 
.A1(n_41),
.A2(n_28),
.B1(n_24),
.B2(n_31),
.Y(n_55)
);

INVx3_ASAP7_75t_L g56 ( 
.A(n_40),
.Y(n_56)
);

CKINVDCx16_ASAP7_75t_R g61 ( 
.A(n_56),
.Y(n_61)
);

CKINVDCx20_ASAP7_75t_R g57 ( 
.A(n_39),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_SL g62 ( 
.A(n_57),
.B(n_41),
.Y(n_62)
);

HB1xp67_ASAP7_75t_L g58 ( 
.A(n_40),
.Y(n_58)
);

CKINVDCx20_ASAP7_75t_R g69 ( 
.A(n_58),
.Y(n_69)
);

OAI22xp5_ASAP7_75t_SL g59 ( 
.A1(n_41),
.A2(n_31),
.B1(n_28),
.B2(n_24),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_L g83 ( 
.A(n_60),
.B(n_76),
.Y(n_83)
);

CKINVDCx14_ASAP7_75t_R g96 ( 
.A(n_62),
.Y(n_96)
);

INVxp67_ASAP7_75t_L g63 ( 
.A(n_46),
.Y(n_63)
);

INVxp67_ASAP7_75t_SL g90 ( 
.A(n_63),
.Y(n_90)
);

AOI22xp5_ASAP7_75t_L g94 ( 
.A1(n_64),
.A2(n_75),
.B1(n_35),
.B2(n_26),
.Y(n_94)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_59),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_SL g84 ( 
.A(n_66),
.B(n_73),
.Y(n_84)
);

OAI21xp5_ASAP7_75t_L g67 ( 
.A1(n_50),
.A2(n_34),
.B(n_38),
.Y(n_67)
);

OAI21xp5_ASAP7_75t_SL g95 ( 
.A1(n_67),
.A2(n_74),
.B(n_29),
.Y(n_95)
);

OAI22xp5_ASAP7_75t_SL g80 ( 
.A1(n_70),
.A2(n_24),
.B1(n_28),
.B2(n_38),
.Y(n_80)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_49),
.Y(n_73)
);

AOI22xp33_ASAP7_75t_L g75 ( 
.A1(n_52),
.A2(n_42),
.B1(n_57),
.B2(n_48),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_SL g76 ( 
.A(n_52),
.B(n_38),
.Y(n_76)
);

CKINVDCx16_ASAP7_75t_R g77 ( 
.A(n_43),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_77),
.B(n_35),
.Y(n_92)
);

CKINVDCx20_ASAP7_75t_R g79 ( 
.A(n_72),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_79),
.B(n_89),
.Y(n_98)
);

AOI22xp5_ASAP7_75t_L g106 ( 
.A1(n_80),
.A2(n_81),
.B1(n_88),
.B2(n_91),
.Y(n_106)
);

OAI22xp5_ASAP7_75t_L g81 ( 
.A1(n_70),
.A2(n_66),
.B1(n_76),
.B2(n_67),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_SL g82 ( 
.A(n_62),
.B(n_23),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_SL g108 ( 
.A(n_82),
.B(n_87),
.Y(n_108)
);

AOI22xp5_ASAP7_75t_SL g85 ( 
.A1(n_67),
.A2(n_43),
.B1(n_38),
.B2(n_20),
.Y(n_85)
);

INVxp67_ASAP7_75t_L g97 ( 
.A(n_85),
.Y(n_97)
);

AOI22xp5_ASAP7_75t_SL g86 ( 
.A1(n_75),
.A2(n_38),
.B1(n_22),
.B2(n_20),
.Y(n_86)
);

INVx1_ASAP7_75t_SL g115 ( 
.A(n_86),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_SL g87 ( 
.A(n_68),
.B(n_38),
.Y(n_87)
);

OAI22xp5_ASAP7_75t_SL g88 ( 
.A1(n_74),
.A2(n_47),
.B1(n_53),
.B2(n_54),
.Y(n_88)
);

INVx5_ASAP7_75t_L g89 ( 
.A(n_77),
.Y(n_89)
);

OAI22xp5_ASAP7_75t_SL g91 ( 
.A1(n_74),
.A2(n_53),
.B1(n_40),
.B2(n_26),
.Y(n_91)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_92),
.Y(n_99)
);

AOI22xp33_ASAP7_75t_SL g93 ( 
.A1(n_71),
.A2(n_35),
.B1(n_56),
.B2(n_44),
.Y(n_93)
);

INVx13_ASAP7_75t_L g111 ( 
.A(n_93),
.Y(n_111)
);

OAI22xp5_ASAP7_75t_L g109 ( 
.A1(n_94),
.A2(n_73),
.B1(n_65),
.B2(n_72),
.Y(n_109)
);

HB1xp67_ASAP7_75t_L g107 ( 
.A(n_95),
.Y(n_107)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_84),
.Y(n_100)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_100),
.Y(n_123)
);

AOI22x1_ASAP7_75t_SL g101 ( 
.A1(n_90),
.A2(n_60),
.B1(n_71),
.B2(n_68),
.Y(n_101)
);

MAJIxp5_ASAP7_75t_SL g120 ( 
.A(n_101),
.B(n_104),
.C(n_114),
.Y(n_120)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_84),
.Y(n_102)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_102),
.Y(n_141)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_92),
.Y(n_103)
);

INVx1_ASAP7_75t_SL g144 ( 
.A(n_103),
.Y(n_144)
);

CKINVDCx20_ASAP7_75t_R g104 ( 
.A(n_82),
.Y(n_104)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_88),
.Y(n_105)
);

CKINVDCx20_ASAP7_75t_R g126 ( 
.A(n_105),
.Y(n_126)
);

AOI22xp5_ASAP7_75t_L g130 ( 
.A1(n_109),
.A2(n_60),
.B1(n_65),
.B2(n_61),
.Y(n_130)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_91),
.Y(n_110)
);

CKINVDCx20_ASAP7_75t_R g136 ( 
.A(n_110),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_L g112 ( 
.A(n_79),
.B(n_69),
.Y(n_112)
);

CKINVDCx14_ASAP7_75t_R g134 ( 
.A(n_112),
.Y(n_134)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_81),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_L g125 ( 
.A(n_113),
.B(n_116),
.Y(n_125)
);

CKINVDCx20_ASAP7_75t_R g114 ( 
.A(n_90),
.Y(n_114)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_94),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_89),
.B(n_69),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_L g140 ( 
.A(n_117),
.B(n_118),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_L g118 ( 
.A(n_89),
.B(n_61),
.Y(n_118)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_80),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_119),
.B(n_110),
.Y(n_127)
);

XOR2xp5_ASAP7_75t_L g121 ( 
.A(n_107),
.B(n_83),
.Y(n_121)
);

XOR2xp5_ASAP7_75t_L g148 ( 
.A(n_121),
.B(n_103),
.Y(n_148)
);

OAI21xp5_ASAP7_75t_L g122 ( 
.A1(n_97),
.A2(n_83),
.B(n_96),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_L g145 ( 
.A(n_122),
.B(n_128),
.Y(n_145)
);

OAI21xp5_ASAP7_75t_SL g124 ( 
.A1(n_97),
.A2(n_95),
.B(n_96),
.Y(n_124)
);

OAI21xp5_ASAP7_75t_SL g163 ( 
.A1(n_124),
.A2(n_138),
.B(n_2),
.Y(n_163)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_127),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_L g128 ( 
.A(n_100),
.B(n_87),
.Y(n_128)
);

OAI22xp5_ASAP7_75t_L g129 ( 
.A1(n_119),
.A2(n_85),
.B1(n_86),
.B2(n_64),
.Y(n_129)
);

AOI22xp5_ASAP7_75t_L g161 ( 
.A1(n_129),
.A2(n_133),
.B1(n_139),
.B2(n_1),
.Y(n_161)
);

NOR2xp33_ASAP7_75t_L g147 ( 
.A(n_130),
.B(n_142),
.Y(n_147)
);

MAJIxp5_ASAP7_75t_L g131 ( 
.A(n_113),
.B(n_26),
.C(n_78),
.Y(n_131)
);

MAJIxp5_ASAP7_75t_L g146 ( 
.A(n_131),
.B(n_137),
.C(n_98),
.Y(n_146)
);

AOI22xp5_ASAP7_75t_L g132 ( 
.A1(n_105),
.A2(n_116),
.B1(n_115),
.B2(n_109),
.Y(n_132)
);

AOI22xp33_ASAP7_75t_L g160 ( 
.A1(n_132),
.A2(n_143),
.B1(n_18),
.B2(n_15),
.Y(n_160)
);

OAI22xp5_ASAP7_75t_SL g133 ( 
.A1(n_106),
.A2(n_78),
.B1(n_49),
.B2(n_22),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_L g135 ( 
.A(n_102),
.B(n_108),
.Y(n_135)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_135),
.Y(n_162)
);

MAJIxp5_ASAP7_75t_L g137 ( 
.A(n_101),
.B(n_26),
.C(n_16),
.Y(n_137)
);

AOI21xp5_ASAP7_75t_L g138 ( 
.A1(n_115),
.A2(n_0),
.B(n_1),
.Y(n_138)
);

OAI22xp5_ASAP7_75t_L g139 ( 
.A1(n_106),
.A2(n_20),
.B1(n_23),
.B2(n_12),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_L g142 ( 
.A(n_108),
.B(n_13),
.Y(n_142)
);

AOI22xp5_ASAP7_75t_L g143 ( 
.A1(n_99),
.A2(n_29),
.B1(n_18),
.B2(n_15),
.Y(n_143)
);

XOR2xp5_ASAP7_75t_L g171 ( 
.A(n_146),
.B(n_152),
.Y(n_171)
);

XNOR2xp5_ASAP7_75t_SL g172 ( 
.A(n_148),
.B(n_154),
.Y(n_172)
);

MAJIxp5_ASAP7_75t_L g149 ( 
.A(n_134),
.B(n_121),
.C(n_140),
.Y(n_149)
);

NOR2xp33_ASAP7_75t_L g170 ( 
.A(n_149),
.B(n_150),
.Y(n_170)
);

MAJIxp5_ASAP7_75t_L g150 ( 
.A(n_130),
.B(n_137),
.C(n_122),
.Y(n_150)
);

XNOR2xp5_ASAP7_75t_SL g152 ( 
.A(n_120),
.B(n_99),
.Y(n_152)
);

AOI22xp33_ASAP7_75t_SL g153 ( 
.A1(n_136),
.A2(n_111),
.B1(n_114),
.B2(n_104),
.Y(n_153)
);

OAI22xp5_ASAP7_75t_L g175 ( 
.A1(n_153),
.A2(n_161),
.B1(n_138),
.B2(n_144),
.Y(n_175)
);

XNOR2xp5_ASAP7_75t_SL g154 ( 
.A(n_120),
.B(n_135),
.Y(n_154)
);

XNOR2xp5_ASAP7_75t_L g155 ( 
.A(n_124),
.B(n_111),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_L g173 ( 
.A(n_155),
.B(n_156),
.Y(n_173)
);

XNOR2xp5_ASAP7_75t_L g156 ( 
.A(n_123),
.B(n_111),
.Y(n_156)
);

XNOR2xp5_ASAP7_75t_L g157 ( 
.A(n_123),
.B(n_13),
.Y(n_157)
);

CKINVDCx16_ASAP7_75t_R g168 ( 
.A(n_157),
.Y(n_168)
);

XNOR2xp5_ASAP7_75t_L g158 ( 
.A(n_141),
.B(n_13),
.Y(n_158)
);

NOR2xp33_ASAP7_75t_SL g174 ( 
.A(n_158),
.B(n_144),
.Y(n_174)
);

XOR2xp5_ASAP7_75t_L g159 ( 
.A(n_128),
.B(n_13),
.Y(n_159)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_159),
.Y(n_164)
);

OR2x2_ASAP7_75t_L g167 ( 
.A(n_160),
.B(n_143),
.Y(n_167)
);

OAI21xp5_ASAP7_75t_SL g176 ( 
.A1(n_163),
.A2(n_141),
.B(n_125),
.Y(n_176)
);

AOI22xp5_ASAP7_75t_L g165 ( 
.A1(n_151),
.A2(n_129),
.B1(n_136),
.B2(n_126),
.Y(n_165)
);

OAI22xp5_ASAP7_75t_SL g183 ( 
.A1(n_165),
.A2(n_166),
.B1(n_167),
.B2(n_146),
.Y(n_183)
);

AOI22xp5_ASAP7_75t_L g166 ( 
.A1(n_152),
.A2(n_126),
.B1(n_125),
.B2(n_127),
.Y(n_166)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_162),
.Y(n_169)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_169),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_L g185 ( 
.A(n_174),
.B(n_176),
.Y(n_185)
);

AOI22xp5_ASAP7_75t_L g180 ( 
.A1(n_175),
.A2(n_133),
.B1(n_147),
.B2(n_153),
.Y(n_180)
);

AOI21xp5_ASAP7_75t_L g177 ( 
.A1(n_145),
.A2(n_132),
.B(n_139),
.Y(n_177)
);

OAI21xp5_ASAP7_75t_SL g187 ( 
.A1(n_177),
.A2(n_29),
.B(n_3),
.Y(n_187)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_154),
.Y(n_178)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_178),
.Y(n_188)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_180),
.Y(n_192)
);

XOR2x2_ASAP7_75t_L g181 ( 
.A(n_178),
.B(n_150),
.Y(n_181)
);

INVxp67_ASAP7_75t_L g197 ( 
.A(n_181),
.Y(n_197)
);

NOR3xp33_ASAP7_75t_SL g182 ( 
.A(n_170),
.B(n_160),
.C(n_148),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_L g193 ( 
.A(n_182),
.B(n_186),
.Y(n_193)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_183),
.Y(n_196)
);

MAJIxp5_ASAP7_75t_L g184 ( 
.A(n_171),
.B(n_159),
.C(n_131),
.Y(n_184)
);

MAJIxp5_ASAP7_75t_L g198 ( 
.A(n_184),
.B(n_166),
.C(n_176),
.Y(n_198)
);

XNOR2xp5_ASAP7_75t_L g186 ( 
.A(n_171),
.B(n_29),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_L g200 ( 
.A(n_187),
.B(n_190),
.Y(n_200)
);

XOR2x2_ASAP7_75t_SL g189 ( 
.A(n_177),
.B(n_21),
.Y(n_189)
);

NOR2xp33_ASAP7_75t_L g191 ( 
.A(n_189),
.B(n_167),
.Y(n_191)
);

AOI22xp5_ASAP7_75t_SL g190 ( 
.A1(n_168),
.A2(n_164),
.B1(n_169),
.B2(n_172),
.Y(n_190)
);

INVxp67_ASAP7_75t_L g207 ( 
.A(n_191),
.Y(n_207)
);

NOR2xp33_ASAP7_75t_L g194 ( 
.A(n_185),
.B(n_165),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_L g202 ( 
.A(n_194),
.B(n_199),
.Y(n_202)
);

AOI22xp5_ASAP7_75t_L g195 ( 
.A1(n_181),
.A2(n_164),
.B1(n_173),
.B2(n_172),
.Y(n_195)
);

OAI22xp5_ASAP7_75t_SL g206 ( 
.A1(n_195),
.A2(n_2),
.B1(n_3),
.B2(n_5),
.Y(n_206)
);

XOR2xp5_ASAP7_75t_L g208 ( 
.A(n_198),
.B(n_21),
.Y(n_208)
);

NOR2xp33_ASAP7_75t_L g199 ( 
.A(n_188),
.B(n_174),
.Y(n_199)
);

AOI21xp5_ASAP7_75t_L g201 ( 
.A1(n_197),
.A2(n_179),
.B(n_186),
.Y(n_201)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_201),
.Y(n_214)
);

OAI21xp5_ASAP7_75t_L g203 ( 
.A1(n_197),
.A2(n_190),
.B(n_184),
.Y(n_203)
);

OAI21xp5_ASAP7_75t_L g215 ( 
.A1(n_203),
.A2(n_204),
.B(n_3),
.Y(n_215)
);

OAI21xp5_ASAP7_75t_L g204 ( 
.A1(n_193),
.A2(n_182),
.B(n_189),
.Y(n_204)
);

NOR2xp33_ASAP7_75t_L g205 ( 
.A(n_196),
.B(n_21),
.Y(n_205)
);

NOR2xp33_ASAP7_75t_L g210 ( 
.A(n_205),
.B(n_14),
.Y(n_210)
);

NOR2xp33_ASAP7_75t_L g213 ( 
.A(n_206),
.B(n_208),
.Y(n_213)
);

AOI322xp5_ASAP7_75t_L g209 ( 
.A1(n_207),
.A2(n_192),
.A3(n_198),
.B1(n_200),
.B2(n_195),
.C1(n_11),
.C2(n_21),
.Y(n_209)
);

AOI21xp5_ASAP7_75t_L g219 ( 
.A1(n_209),
.A2(n_211),
.B(n_215),
.Y(n_219)
);

XOR2xp5_ASAP7_75t_L g217 ( 
.A(n_210),
.B(n_14),
.Y(n_217)
);

NAND5xp2_ASAP7_75t_L g211 ( 
.A(n_202),
.B(n_14),
.C(n_11),
.D(n_5),
.E(n_6),
.Y(n_211)
);

NOR2xp33_ASAP7_75t_SL g212 ( 
.A(n_205),
.B(n_2),
.Y(n_212)
);

NOR2xp33_ASAP7_75t_SL g216 ( 
.A(n_212),
.B(n_3),
.Y(n_216)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_216),
.Y(n_222)
);

MAJIxp5_ASAP7_75t_L g221 ( 
.A(n_217),
.B(n_220),
.C(n_210),
.Y(n_221)
);

NAND3xp33_ASAP7_75t_L g218 ( 
.A(n_214),
.B(n_5),
.C(n_6),
.Y(n_218)
);

AOI21xp33_ASAP7_75t_L g223 ( 
.A1(n_218),
.A2(n_5),
.B(n_7),
.Y(n_223)
);

OAI21xp5_ASAP7_75t_SL g220 ( 
.A1(n_213),
.A2(n_14),
.B(n_6),
.Y(n_220)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_221),
.Y(n_224)
);

OAI21xp5_ASAP7_75t_L g225 ( 
.A1(n_223),
.A2(n_219),
.B(n_8),
.Y(n_225)
);

AOI322xp5_ASAP7_75t_L g226 ( 
.A1(n_225),
.A2(n_7),
.A3(n_8),
.B1(n_9),
.B2(n_222),
.C1(n_224),
.C2(n_216),
.Y(n_226)
);

AOI22x1_ASAP7_75t_SL g227 ( 
.A1(n_226),
.A2(n_7),
.B1(n_8),
.B2(n_9),
.Y(n_227)
);

NAND2xp5_ASAP7_75t_L g228 ( 
.A(n_227),
.B(n_7),
.Y(n_228)
);


endmodule