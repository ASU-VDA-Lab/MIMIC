module fake_jpeg_14089_n_632 (n_13, n_1, n_10, n_6, n_14, n_18, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_632);

input n_13;
input n_1;
input n_10;
input n_6;
input n_14;
input n_18;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_632;

wire n_529;
wire n_595;
wire n_390;
wire n_552;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_525;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_586;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_620;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_611;
wire n_44;
wire n_355;
wire n_519;
wire n_276;
wire n_143;
wire n_431;
wire n_102;
wire n_549;
wire n_196;
wire n_66;
wire n_374;
wire n_566;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_597;
wire n_172;
wire n_547;
wire n_345;
wire n_591;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_513;
wire n_283;
wire n_107;
wire n_490;
wire n_517;
wire n_629;
wire n_415;
wire n_479;
wire n_543;
wire n_357;
wire n_89;
wire n_131;
wire n_607;
wire n_294;
wire n_230;
wire n_170;
wire n_602;
wire n_313;
wire n_542;
wire n_574;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_559;
wire n_48;
wire n_465;
wire n_200;
wire n_582;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_623;
wire n_579;
wire n_416;
wire n_221;
wire n_256;
wire n_454;
wire n_540;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_571;
wire n_82;
wire n_155;
wire n_508;
wire n_309;
wire n_624;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_606;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_569;
wire n_596;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_544;
wire n_31;
wire n_277;
wire n_255;
wire n_605;
wire n_601;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_349;
wire n_21;
wire n_393;
wire n_288;
wire n_234;
wire n_530;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_557;
wire n_408;
wire n_80;
wire n_562;
wire n_204;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_298;
wire n_106;
wire n_545;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_584;
wire n_254;
wire n_608;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_622;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_474;
wire n_539;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_626;
wire n_300;
wire n_442;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_575;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_511;
wire n_305;
wire n_161;
wire n_441;
wire n_555;
wire n_342;
wire n_101;
wire n_226;
wire n_509;
wire n_149;
wire n_87;
wire n_46;
wire n_578;
wire n_589;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_614;
wire n_97;
wire n_573;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_610;
wire n_174;
wire n_198;
wire n_422;
wire n_560;
wire n_190;
wire n_510;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_536;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_537;
wire n_110;
wire n_594;
wire n_590;
wire n_531;
wire n_76;
wire n_278;
wire n_343;
wire n_577;
wire n_26;
wire n_88;
wire n_397;
wire n_592;
wire n_363;
wire n_570;
wire n_238;
wire n_598;
wire n_615;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_554;
wire n_301;
wire n_609;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_523;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_533;
wire n_612;
wire n_296;
wire n_384;
wire n_588;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_585;
wire n_491;
wire n_24;
wire n_526;
wire n_467;
wire n_269;
wire n_572;
wire n_546;
wire n_287;
wire n_219;
wire n_452;
wire n_631;
wire n_433;
wire n_77;
wire n_473;
wire n_45;
wire n_520;
wire n_476;
wire n_337;
wire n_317;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_599;
wire n_239;
wire n_243;
wire n_481;
wire n_628;
wire n_619;
wire n_348;
wire n_587;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_583;
wire n_522;
wire n_333;
wire n_518;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_565;
wire n_302;
wire n_216;
wire n_528;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_199;
wire n_260;
wire n_550;
wire n_413;
wire n_275;
wire n_494;
wire n_604;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_551;
wire n_36;
wire n_62;
wire n_600;
wire n_492;
wire n_603;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_567;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_515;
wire n_347;
wire n_521;
wire n_424;
wire n_55;
wire n_358;
wire n_312;
wire n_47;
wire n_538;
wire n_625;
wire n_147;
wire n_449;
wire n_627;
wire n_98;
wire n_251;
wire n_534;
wire n_472;
wire n_279;
wire n_593;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_618;
wire n_356;
wire n_119;
wire n_484;
wire n_568;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_576;
wire n_469;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_553;
wire n_257;
wire n_61;
wire n_173;
wire n_561;
wire n_244;
wire n_232;
wire n_527;
wire n_482;
wire n_58;
wire n_41;
wire n_613;
wire n_630;
wire n_266;
wire n_548;
wire n_72;
wire n_512;
wire n_445;
wire n_443;
wire n_617;
wire n_215;
wire n_212;
wire n_516;
wire n_183;
wire n_409;
wire n_532;
wire n_249;
wire n_412;
wire n_581;
wire n_217;
wire n_471;
wire n_580;
wire n_541;
wire n_53;
wire n_372;
wire n_558;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_535;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_556;
wire n_524;
wire n_402;
wire n_563;
wire n_504;
wire n_438;
wire n_475;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_616;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_514;
wire n_564;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_621;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

INVx8_ASAP7_75t_L g19 ( 
.A(n_1),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_8),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_4),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_16),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_4),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_13),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_13),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_14),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_9),
.Y(n_27)
);

INVx4_ASAP7_75t_L g28 ( 
.A(n_11),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_3),
.Y(n_29)
);

BUFx12f_ASAP7_75t_L g30 ( 
.A(n_4),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_3),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_9),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_18),
.Y(n_33)
);

BUFx5_ASAP7_75t_L g34 ( 
.A(n_10),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_2),
.Y(n_35)
);

CKINVDCx16_ASAP7_75t_R g36 ( 
.A(n_7),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_9),
.Y(n_37)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_11),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_14),
.Y(n_39)
);

INVx8_ASAP7_75t_L g40 ( 
.A(n_12),
.Y(n_40)
);

INVx6_ASAP7_75t_SL g41 ( 
.A(n_4),
.Y(n_41)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_16),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_7),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_10),
.Y(n_44)
);

BUFx3_ASAP7_75t_L g45 ( 
.A(n_18),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_16),
.Y(n_46)
);

BUFx12f_ASAP7_75t_L g47 ( 
.A(n_2),
.Y(n_47)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_3),
.Y(n_48)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_7),
.Y(n_49)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_8),
.Y(n_50)
);

INVx2_ASAP7_75t_L g51 ( 
.A(n_8),
.Y(n_51)
);

INVx13_ASAP7_75t_L g52 ( 
.A(n_1),
.Y(n_52)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_3),
.Y(n_53)
);

INVx3_ASAP7_75t_L g54 ( 
.A(n_8),
.Y(n_54)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_13),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_6),
.Y(n_56)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_6),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_0),
.Y(n_58)
);

BUFx10_ASAP7_75t_L g59 ( 
.A(n_18),
.Y(n_59)
);

BUFx5_ASAP7_75t_L g60 ( 
.A(n_15),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_10),
.Y(n_61)
);

INVx6_ASAP7_75t_L g62 ( 
.A(n_61),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g159 ( 
.A(n_62),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_SL g63 ( 
.A(n_22),
.B(n_17),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_L g158 ( 
.A(n_63),
.B(n_80),
.Y(n_158)
);

INVx2_ASAP7_75t_L g64 ( 
.A(n_51),
.Y(n_64)
);

INVx2_ASAP7_75t_L g131 ( 
.A(n_64),
.Y(n_131)
);

INVx8_ASAP7_75t_L g65 ( 
.A(n_41),
.Y(n_65)
);

INVx5_ASAP7_75t_L g185 ( 
.A(n_65),
.Y(n_185)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_20),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g164 ( 
.A(n_66),
.Y(n_164)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_33),
.Y(n_67)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_67),
.Y(n_132)
);

BUFx3_ASAP7_75t_L g68 ( 
.A(n_34),
.Y(n_68)
);

BUFx12f_ASAP7_75t_L g135 ( 
.A(n_68),
.Y(n_135)
);

INVx8_ASAP7_75t_L g69 ( 
.A(n_41),
.Y(n_69)
);

INVx5_ASAP7_75t_L g196 ( 
.A(n_69),
.Y(n_196)
);

CKINVDCx20_ASAP7_75t_R g70 ( 
.A(n_59),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g136 ( 
.A(n_70),
.B(n_83),
.Y(n_136)
);

BUFx6f_ASAP7_75t_L g71 ( 
.A(n_20),
.Y(n_71)
);

BUFx6f_ASAP7_75t_L g167 ( 
.A(n_71),
.Y(n_167)
);

BUFx6f_ASAP7_75t_L g72 ( 
.A(n_20),
.Y(n_72)
);

BUFx6f_ASAP7_75t_L g179 ( 
.A(n_72),
.Y(n_179)
);

BUFx6f_ASAP7_75t_L g73 ( 
.A(n_23),
.Y(n_73)
);

BUFx6f_ASAP7_75t_L g188 ( 
.A(n_73),
.Y(n_188)
);

BUFx12f_ASAP7_75t_L g74 ( 
.A(n_34),
.Y(n_74)
);

BUFx3_ASAP7_75t_L g130 ( 
.A(n_74),
.Y(n_130)
);

BUFx3_ASAP7_75t_L g75 ( 
.A(n_34),
.Y(n_75)
);

BUFx12f_ASAP7_75t_L g141 ( 
.A(n_75),
.Y(n_141)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_33),
.Y(n_76)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_76),
.Y(n_140)
);

BUFx12f_ASAP7_75t_L g77 ( 
.A(n_60),
.Y(n_77)
);

BUFx3_ASAP7_75t_L g137 ( 
.A(n_77),
.Y(n_137)
);

INVx11_ASAP7_75t_L g78 ( 
.A(n_52),
.Y(n_78)
);

BUFx10_ASAP7_75t_L g149 ( 
.A(n_78),
.Y(n_149)
);

INVx4_ASAP7_75t_L g79 ( 
.A(n_28),
.Y(n_79)
);

INVx3_ASAP7_75t_L g146 ( 
.A(n_79),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_L g80 ( 
.A(n_22),
.B(n_17),
.Y(n_80)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_42),
.Y(n_81)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_81),
.Y(n_142)
);

BUFx3_ASAP7_75t_L g82 ( 
.A(n_30),
.Y(n_82)
);

BUFx12f_ASAP7_75t_L g172 ( 
.A(n_82),
.Y(n_172)
);

CKINVDCx20_ASAP7_75t_R g83 ( 
.A(n_59),
.Y(n_83)
);

INVx4_ASAP7_75t_L g84 ( 
.A(n_28),
.Y(n_84)
);

INVx3_ASAP7_75t_L g150 ( 
.A(n_84),
.Y(n_150)
);

INVx4_ASAP7_75t_L g85 ( 
.A(n_28),
.Y(n_85)
);

INVx3_ASAP7_75t_L g189 ( 
.A(n_85),
.Y(n_189)
);

BUFx6f_ASAP7_75t_L g86 ( 
.A(n_23),
.Y(n_86)
);

INVx6_ASAP7_75t_L g154 ( 
.A(n_86),
.Y(n_154)
);

BUFx6f_ASAP7_75t_L g87 ( 
.A(n_23),
.Y(n_87)
);

INVx6_ASAP7_75t_L g165 ( 
.A(n_87),
.Y(n_165)
);

INVx2_ASAP7_75t_L g88 ( 
.A(n_51),
.Y(n_88)
);

INVx2_ASAP7_75t_L g133 ( 
.A(n_88),
.Y(n_133)
);

BUFx5_ASAP7_75t_L g89 ( 
.A(n_60),
.Y(n_89)
);

BUFx12f_ASAP7_75t_L g177 ( 
.A(n_89),
.Y(n_177)
);

INVx3_ASAP7_75t_L g90 ( 
.A(n_60),
.Y(n_90)
);

INVx3_ASAP7_75t_L g191 ( 
.A(n_90),
.Y(n_191)
);

INVx11_ASAP7_75t_SL g91 ( 
.A(n_52),
.Y(n_91)
);

BUFx24_ASAP7_75t_L g201 ( 
.A(n_91),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_L g92 ( 
.A(n_21),
.B(n_17),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_L g173 ( 
.A(n_92),
.B(n_120),
.Y(n_173)
);

BUFx6f_ASAP7_75t_L g93 ( 
.A(n_25),
.Y(n_93)
);

INVx6_ASAP7_75t_L g166 ( 
.A(n_93),
.Y(n_166)
);

INVx3_ASAP7_75t_L g94 ( 
.A(n_45),
.Y(n_94)
);

INVx3_ASAP7_75t_L g200 ( 
.A(n_94),
.Y(n_200)
);

BUFx16f_ASAP7_75t_L g95 ( 
.A(n_30),
.Y(n_95)
);

INVx6_ASAP7_75t_SL g195 ( 
.A(n_95),
.Y(n_195)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_42),
.B(n_15),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_SL g148 ( 
.A(n_96),
.B(n_99),
.Y(n_148)
);

CKINVDCx20_ASAP7_75t_R g97 ( 
.A(n_59),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g151 ( 
.A(n_97),
.B(n_112),
.Y(n_151)
);

BUFx3_ASAP7_75t_L g98 ( 
.A(n_30),
.Y(n_98)
);

BUFx12f_ASAP7_75t_L g180 ( 
.A(n_98),
.Y(n_180)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_45),
.B(n_15),
.Y(n_99)
);

INVx5_ASAP7_75t_L g100 ( 
.A(n_19),
.Y(n_100)
);

INVx2_ASAP7_75t_SL g181 ( 
.A(n_100),
.Y(n_181)
);

BUFx6f_ASAP7_75t_L g101 ( 
.A(n_25),
.Y(n_101)
);

INVx6_ASAP7_75t_L g175 ( 
.A(n_101),
.Y(n_175)
);

BUFx3_ASAP7_75t_L g102 ( 
.A(n_30),
.Y(n_102)
);

BUFx12f_ASAP7_75t_L g197 ( 
.A(n_102),
.Y(n_197)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_31),
.Y(n_103)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_103),
.Y(n_143)
);

BUFx6f_ASAP7_75t_L g104 ( 
.A(n_25),
.Y(n_104)
);

INVx6_ASAP7_75t_L g184 ( 
.A(n_104),
.Y(n_184)
);

BUFx6f_ASAP7_75t_L g105 ( 
.A(n_37),
.Y(n_105)
);

INVx8_ASAP7_75t_L g182 ( 
.A(n_105),
.Y(n_182)
);

INVx2_ASAP7_75t_L g106 ( 
.A(n_54),
.Y(n_106)
);

INVx2_ASAP7_75t_L g145 ( 
.A(n_106),
.Y(n_145)
);

INVx8_ASAP7_75t_L g107 ( 
.A(n_37),
.Y(n_107)
);

INVx2_ASAP7_75t_L g169 ( 
.A(n_107),
.Y(n_169)
);

INVx6_ASAP7_75t_L g108 ( 
.A(n_37),
.Y(n_108)
);

BUFx3_ASAP7_75t_L g205 ( 
.A(n_108),
.Y(n_205)
);

INVx2_ASAP7_75t_L g109 ( 
.A(n_54),
.Y(n_109)
);

INVx2_ASAP7_75t_L g186 ( 
.A(n_109),
.Y(n_186)
);

BUFx6f_ASAP7_75t_L g110 ( 
.A(n_39),
.Y(n_110)
);

BUFx12f_ASAP7_75t_L g207 ( 
.A(n_110),
.Y(n_207)
);

BUFx6f_ASAP7_75t_L g111 ( 
.A(n_39),
.Y(n_111)
);

INVx2_ASAP7_75t_L g190 ( 
.A(n_111),
.Y(n_190)
);

INVx2_ASAP7_75t_R g112 ( 
.A(n_59),
.Y(n_112)
);

BUFx6f_ASAP7_75t_L g113 ( 
.A(n_39),
.Y(n_113)
);

INVx2_ASAP7_75t_L g193 ( 
.A(n_113),
.Y(n_193)
);

INVx4_ASAP7_75t_L g114 ( 
.A(n_30),
.Y(n_114)
);

HB1xp67_ASAP7_75t_L g139 ( 
.A(n_114),
.Y(n_139)
);

BUFx5_ASAP7_75t_L g115 ( 
.A(n_59),
.Y(n_115)
);

BUFx10_ASAP7_75t_L g203 ( 
.A(n_115),
.Y(n_203)
);

CKINVDCx20_ASAP7_75t_R g116 ( 
.A(n_45),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_L g155 ( 
.A(n_116),
.B(n_122),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_21),
.B(n_0),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_SL g156 ( 
.A(n_117),
.B(n_36),
.Y(n_156)
);

INVx2_ASAP7_75t_L g118 ( 
.A(n_54),
.Y(n_118)
);

INVx2_ASAP7_75t_L g199 ( 
.A(n_118),
.Y(n_199)
);

BUFx2_ASAP7_75t_L g119 ( 
.A(n_19),
.Y(n_119)
);

INVx2_ASAP7_75t_L g209 ( 
.A(n_119),
.Y(n_209)
);

NAND2xp5_ASAP7_75t_SL g120 ( 
.A(n_24),
.B(n_0),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_SL g121 ( 
.A(n_24),
.B(n_0),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_L g174 ( 
.A(n_121),
.B(n_1),
.Y(n_174)
);

CKINVDCx20_ASAP7_75t_R g122 ( 
.A(n_52),
.Y(n_122)
);

INVx3_ASAP7_75t_L g123 ( 
.A(n_47),
.Y(n_123)
);

INVx2_ASAP7_75t_L g210 ( 
.A(n_123),
.Y(n_210)
);

BUFx6f_ASAP7_75t_L g124 ( 
.A(n_43),
.Y(n_124)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_124),
.Y(n_152)
);

CKINVDCx20_ASAP7_75t_R g125 ( 
.A(n_31),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_L g161 ( 
.A(n_125),
.B(n_128),
.Y(n_161)
);

INVx11_ASAP7_75t_L g126 ( 
.A(n_36),
.Y(n_126)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_126),
.Y(n_176)
);

INVx3_ASAP7_75t_L g127 ( 
.A(n_47),
.Y(n_127)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_127),
.Y(n_178)
);

INVxp67_ASAP7_75t_L g128 ( 
.A(n_32),
.Y(n_128)
);

AOI22xp33_ASAP7_75t_L g129 ( 
.A1(n_62),
.A2(n_61),
.B1(n_58),
.B2(n_43),
.Y(n_129)
);

OAI22xp5_ASAP7_75t_SL g241 ( 
.A1(n_129),
.A2(n_162),
.B1(n_192),
.B2(n_44),
.Y(n_241)
);

CKINVDCx20_ASAP7_75t_R g134 ( 
.A(n_78),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_SL g227 ( 
.A(n_134),
.B(n_138),
.Y(n_227)
);

CKINVDCx20_ASAP7_75t_R g138 ( 
.A(n_126),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_SL g144 ( 
.A(n_112),
.B(n_35),
.Y(n_144)
);

NOR2xp33_ASAP7_75t_SL g258 ( 
.A(n_144),
.B(n_156),
.Y(n_258)
);

AND2x2_ASAP7_75t_SL g147 ( 
.A(n_79),
.B(n_84),
.Y(n_147)
);

MAJIxp5_ASAP7_75t_L g240 ( 
.A(n_147),
.B(n_194),
.C(n_32),
.Y(n_240)
);

AOI22xp5_ASAP7_75t_SL g153 ( 
.A1(n_68),
.A2(n_46),
.B1(n_58),
.B2(n_56),
.Y(n_153)
);

AOI21xp5_ASAP7_75t_L g274 ( 
.A1(n_153),
.A2(n_38),
.B(n_40),
.Y(n_274)
);

NOR2xp33_ASAP7_75t_SL g157 ( 
.A(n_128),
.B(n_35),
.Y(n_157)
);

NOR2xp33_ASAP7_75t_SL g268 ( 
.A(n_157),
.B(n_168),
.Y(n_268)
);

NAND2xp5_ASAP7_75t_SL g160 ( 
.A(n_65),
.B(n_29),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_L g217 ( 
.A(n_160),
.B(n_174),
.Y(n_217)
);

AOI22xp33_ASAP7_75t_L g162 ( 
.A1(n_108),
.A2(n_61),
.B1(n_58),
.B2(n_56),
.Y(n_162)
);

BUFx12_ASAP7_75t_L g163 ( 
.A(n_91),
.Y(n_163)
);

CKINVDCx6p67_ASAP7_75t_R g228 ( 
.A(n_163),
.Y(n_228)
);

CKINVDCx20_ASAP7_75t_R g168 ( 
.A(n_95),
.Y(n_168)
);

NOR2xp33_ASAP7_75t_L g170 ( 
.A(n_69),
.B(n_29),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_SL g230 ( 
.A(n_170),
.B(n_171),
.Y(n_230)
);

NOR2xp33_ASAP7_75t_L g171 ( 
.A(n_77),
.B(n_53),
.Y(n_171)
);

NOR2xp33_ASAP7_75t_SL g183 ( 
.A(n_77),
.B(n_53),
.Y(n_183)
);

NOR2xp33_ASAP7_75t_L g214 ( 
.A(n_183),
.B(n_202),
.Y(n_214)
);

OAI22xp5_ASAP7_75t_L g187 ( 
.A1(n_66),
.A2(n_46),
.B1(n_124),
.B2(n_86),
.Y(n_187)
);

AOI22xp5_ASAP7_75t_L g278 ( 
.A1(n_187),
.A2(n_208),
.B1(n_104),
.B2(n_101),
.Y(n_278)
);

AOI22xp33_ASAP7_75t_L g192 ( 
.A1(n_71),
.A2(n_44),
.B1(n_56),
.B2(n_43),
.Y(n_192)
);

MAJIxp5_ASAP7_75t_L g194 ( 
.A(n_127),
.B(n_57),
.C(n_55),
.Y(n_194)
);

NOR2xp33_ASAP7_75t_L g198 ( 
.A(n_82),
.B(n_26),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_L g245 ( 
.A(n_198),
.B(n_204),
.Y(n_245)
);

OR2x2_ASAP7_75t_L g202 ( 
.A(n_85),
.B(n_57),
.Y(n_202)
);

NOR2xp33_ASAP7_75t_L g204 ( 
.A(n_98),
.B(n_26),
.Y(n_204)
);

NOR2xp33_ASAP7_75t_L g206 ( 
.A(n_102),
.B(n_27),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_L g247 ( 
.A(n_206),
.B(n_74),
.Y(n_247)
);

OAI22xp5_ASAP7_75t_L g208 ( 
.A1(n_72),
.A2(n_46),
.B1(n_44),
.B2(n_48),
.Y(n_208)
);

AOI21xp33_ASAP7_75t_L g211 ( 
.A1(n_74),
.A2(n_49),
.B(n_48),
.Y(n_211)
);

NOR2xp33_ASAP7_75t_L g221 ( 
.A(n_211),
.B(n_47),
.Y(n_221)
);

BUFx6f_ASAP7_75t_L g212 ( 
.A(n_164),
.Y(n_212)
);

INVx5_ASAP7_75t_L g317 ( 
.A(n_212),
.Y(n_317)
);

CKINVDCx12_ASAP7_75t_R g213 ( 
.A(n_201),
.Y(n_213)
);

INVx4_ASAP7_75t_SL g300 ( 
.A(n_213),
.Y(n_300)
);

INVx2_ASAP7_75t_L g215 ( 
.A(n_143),
.Y(n_215)
);

INVx2_ASAP7_75t_L g286 ( 
.A(n_215),
.Y(n_286)
);

CKINVDCx20_ASAP7_75t_R g216 ( 
.A(n_136),
.Y(n_216)
);

NOR2xp33_ASAP7_75t_L g297 ( 
.A(n_216),
.B(n_236),
.Y(n_297)
);

INVx4_ASAP7_75t_L g218 ( 
.A(n_207),
.Y(n_218)
);

INVx3_ASAP7_75t_L g324 ( 
.A(n_218),
.Y(n_324)
);

AND2x2_ASAP7_75t_SL g219 ( 
.A(n_131),
.B(n_114),
.Y(n_219)
);

AND2x2_ASAP7_75t_L g289 ( 
.A(n_219),
.B(n_221),
.Y(n_289)
);

OAI22xp33_ASAP7_75t_SL g220 ( 
.A1(n_202),
.A2(n_87),
.B1(n_113),
.B2(n_111),
.Y(n_220)
);

AOI22xp5_ASAP7_75t_L g326 ( 
.A1(n_220),
.A2(n_241),
.B1(n_243),
.B2(n_205),
.Y(n_326)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_132),
.Y(n_222)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_222),
.Y(n_293)
);

INVx3_ASAP7_75t_L g223 ( 
.A(n_209),
.Y(n_223)
);

INVx3_ASAP7_75t_L g341 ( 
.A(n_223),
.Y(n_341)
);

INVx4_ASAP7_75t_L g224 ( 
.A(n_207),
.Y(n_224)
);

INVx2_ASAP7_75t_L g288 ( 
.A(n_224),
.Y(n_288)
);

INVx2_ASAP7_75t_L g225 ( 
.A(n_140),
.Y(n_225)
);

INVx2_ASAP7_75t_L g299 ( 
.A(n_225),
.Y(n_299)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_142),
.Y(n_226)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_226),
.Y(n_294)
);

AOI22xp33_ASAP7_75t_SL g229 ( 
.A1(n_177),
.A2(n_119),
.B1(n_19),
.B2(n_40),
.Y(n_229)
);

AOI22xp33_ASAP7_75t_SL g308 ( 
.A1(n_229),
.A2(n_257),
.B1(n_265),
.B2(n_266),
.Y(n_308)
);

INVx6_ASAP7_75t_L g231 ( 
.A(n_164),
.Y(n_231)
);

INVx2_ASAP7_75t_L g322 ( 
.A(n_231),
.Y(n_322)
);

NOR2xp33_ASAP7_75t_L g232 ( 
.A(n_161),
.B(n_50),
.Y(n_232)
);

INVxp67_ASAP7_75t_L g302 ( 
.A(n_232),
.Y(n_302)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_155),
.Y(n_233)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_233),
.Y(n_316)
);

INVx2_ASAP7_75t_L g234 ( 
.A(n_145),
.Y(n_234)
);

INVx2_ASAP7_75t_L g344 ( 
.A(n_234),
.Y(n_344)
);

INVx2_ASAP7_75t_L g235 ( 
.A(n_186),
.Y(n_235)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_235),
.Y(n_319)
);

CKINVDCx20_ASAP7_75t_R g236 ( 
.A(n_201),
.Y(n_236)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_178),
.Y(n_237)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_237),
.Y(n_334)
);

INVx2_ASAP7_75t_L g238 ( 
.A(n_199),
.Y(n_238)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_238),
.Y(n_337)
);

INVx4_ASAP7_75t_L g239 ( 
.A(n_207),
.Y(n_239)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_239),
.Y(n_292)
);

AND2x2_ASAP7_75t_L g290 ( 
.A(n_240),
.B(n_261),
.Y(n_290)
);

INVx6_ASAP7_75t_SL g242 ( 
.A(n_201),
.Y(n_242)
);

CKINVDCx16_ASAP7_75t_R g303 ( 
.A(n_242),
.Y(n_303)
);

OAI22xp33_ASAP7_75t_L g243 ( 
.A1(n_192),
.A2(n_110),
.B1(n_73),
.B2(n_105),
.Y(n_243)
);

BUFx6f_ASAP7_75t_L g244 ( 
.A(n_167),
.Y(n_244)
);

BUFx3_ASAP7_75t_L g330 ( 
.A(n_244),
.Y(n_330)
);

OAI21xp33_ASAP7_75t_SL g246 ( 
.A1(n_129),
.A2(n_100),
.B(n_49),
.Y(n_246)
);

AOI21xp5_ASAP7_75t_SL g307 ( 
.A1(n_246),
.A2(n_203),
.B(n_182),
.Y(n_307)
);

NOR2xp33_ASAP7_75t_L g298 ( 
.A(n_247),
.B(n_249),
.Y(n_298)
);

NOR2xp33_ASAP7_75t_L g248 ( 
.A(n_148),
.B(n_55),
.Y(n_248)
);

INVxp67_ASAP7_75t_L g312 ( 
.A(n_248),
.Y(n_312)
);

CKINVDCx12_ASAP7_75t_R g249 ( 
.A(n_195),
.Y(n_249)
);

INVx6_ASAP7_75t_L g250 ( 
.A(n_167),
.Y(n_250)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_250),
.Y(n_325)
);

BUFx3_ASAP7_75t_L g251 ( 
.A(n_172),
.Y(n_251)
);

INVx2_ASAP7_75t_SL g331 ( 
.A(n_251),
.Y(n_331)
);

INVx5_ASAP7_75t_L g252 ( 
.A(n_135),
.Y(n_252)
);

INVx11_ASAP7_75t_L g340 ( 
.A(n_252),
.Y(n_340)
);

INVx2_ASAP7_75t_L g253 ( 
.A(n_190),
.Y(n_253)
);

NOR2xp33_ASAP7_75t_L g309 ( 
.A(n_253),
.B(n_254),
.Y(n_309)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_139),
.Y(n_254)
);

BUFx3_ASAP7_75t_L g255 ( 
.A(n_172),
.Y(n_255)
);

NOR2xp33_ASAP7_75t_L g314 ( 
.A(n_255),
.B(n_256),
.Y(n_314)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_139),
.Y(n_256)
);

AOI22xp33_ASAP7_75t_SL g257 ( 
.A1(n_177),
.A2(n_40),
.B1(n_75),
.B2(n_107),
.Y(n_257)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_152),
.Y(n_259)
);

NOR2xp33_ASAP7_75t_L g320 ( 
.A(n_259),
.B(n_260),
.Y(n_320)
);

INVx2_ASAP7_75t_L g260 ( 
.A(n_193),
.Y(n_260)
);

NOR2xp33_ASAP7_75t_L g261 ( 
.A(n_151),
.B(n_50),
.Y(n_261)
);

NAND2xp5_ASAP7_75t_L g262 ( 
.A(n_158),
.B(n_27),
.Y(n_262)
);

NAND2xp5_ASAP7_75t_L g304 ( 
.A(n_262),
.B(n_271),
.Y(n_304)
);

INVx3_ASAP7_75t_L g263 ( 
.A(n_169),
.Y(n_263)
);

AND2x2_ASAP7_75t_L g339 ( 
.A(n_263),
.B(n_264),
.Y(n_339)
);

CKINVDCx20_ASAP7_75t_R g264 ( 
.A(n_163),
.Y(n_264)
);

INVx6_ASAP7_75t_L g265 ( 
.A(n_179),
.Y(n_265)
);

BUFx3_ASAP7_75t_L g266 ( 
.A(n_172),
.Y(n_266)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_200),
.Y(n_267)
);

AOI22xp33_ASAP7_75t_SL g335 ( 
.A1(n_267),
.A2(n_269),
.B1(n_270),
.B2(n_272),
.Y(n_335)
);

BUFx6f_ASAP7_75t_L g269 ( 
.A(n_179),
.Y(n_269)
);

BUFx6f_ASAP7_75t_L g270 ( 
.A(n_188),
.Y(n_270)
);

NAND2xp5_ASAP7_75t_L g271 ( 
.A(n_173),
.B(n_133),
.Y(n_271)
);

INVx2_ASAP7_75t_L g272 ( 
.A(n_210),
.Y(n_272)
);

INVx13_ASAP7_75t_L g273 ( 
.A(n_163),
.Y(n_273)
);

AOI22xp33_ASAP7_75t_SL g338 ( 
.A1(n_273),
.A2(n_276),
.B1(n_277),
.B2(n_279),
.Y(n_338)
);

OAI22xp5_ASAP7_75t_L g291 ( 
.A1(n_274),
.A2(n_278),
.B1(n_162),
.B2(n_181),
.Y(n_291)
);

NOR2xp33_ASAP7_75t_L g275 ( 
.A(n_196),
.B(n_38),
.Y(n_275)
);

NAND2xp5_ASAP7_75t_L g327 ( 
.A(n_275),
.B(n_280),
.Y(n_327)
);

INVx3_ASAP7_75t_L g276 ( 
.A(n_185),
.Y(n_276)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_146),
.Y(n_277)
);

AOI22xp33_ASAP7_75t_SL g279 ( 
.A1(n_177),
.A2(n_47),
.B1(n_93),
.B2(n_5),
.Y(n_279)
);

CKINVDCx20_ASAP7_75t_R g280 ( 
.A(n_149),
.Y(n_280)
);

NAND2xp5_ASAP7_75t_L g281 ( 
.A(n_147),
.B(n_176),
.Y(n_281)
);

NAND2xp5_ASAP7_75t_L g333 ( 
.A(n_281),
.B(n_282),
.Y(n_333)
);

NOR2xp33_ASAP7_75t_L g282 ( 
.A(n_185),
.B(n_47),
.Y(n_282)
);

INVx2_ASAP7_75t_L g283 ( 
.A(n_150),
.Y(n_283)
);

AOI22xp33_ASAP7_75t_SL g342 ( 
.A1(n_283),
.A2(n_284),
.B1(n_285),
.B2(n_2),
.Y(n_342)
);

INVx4_ASAP7_75t_L g284 ( 
.A(n_180),
.Y(n_284)
);

INVx3_ASAP7_75t_L g285 ( 
.A(n_149),
.Y(n_285)
);

AOI22xp5_ASAP7_75t_SL g287 ( 
.A1(n_220),
.A2(n_130),
.B1(n_181),
.B2(n_135),
.Y(n_287)
);

INVxp67_ASAP7_75t_L g357 ( 
.A(n_287),
.Y(n_357)
);

AOI22xp5_ASAP7_75t_L g347 ( 
.A1(n_291),
.A2(n_295),
.B1(n_296),
.B2(n_301),
.Y(n_347)
);

OAI22xp5_ASAP7_75t_SL g295 ( 
.A1(n_278),
.A2(n_159),
.B1(n_175),
.B2(n_166),
.Y(n_295)
);

OAI22xp5_ASAP7_75t_L g296 ( 
.A1(n_274),
.A2(n_175),
.B1(n_154),
.B2(n_184),
.Y(n_296)
);

OAI22xp5_ASAP7_75t_L g301 ( 
.A1(n_214),
.A2(n_166),
.B1(n_154),
.B2(n_165),
.Y(n_301)
);

OAI22xp5_ASAP7_75t_L g305 ( 
.A1(n_240),
.A2(n_184),
.B1(n_165),
.B2(n_188),
.Y(n_305)
);

AOI22xp5_ASAP7_75t_L g349 ( 
.A1(n_305),
.A2(n_318),
.B1(n_295),
.B2(n_321),
.Y(n_349)
);

A2O1A1Ixp33_ASAP7_75t_L g306 ( 
.A1(n_217),
.A2(n_149),
.B(n_203),
.C(n_189),
.Y(n_306)
);

NAND2xp5_ASAP7_75t_L g346 ( 
.A(n_306),
.B(n_336),
.Y(n_346)
);

AND2x2_ASAP7_75t_L g362 ( 
.A(n_307),
.B(n_310),
.Y(n_362)
);

AND2x2_ASAP7_75t_SL g310 ( 
.A(n_245),
.B(n_130),
.Y(n_310)
);

OA22x2_ASAP7_75t_L g311 ( 
.A1(n_246),
.A2(n_241),
.B1(n_243),
.B2(n_219),
.Y(n_311)
);

A2O1A1Ixp33_ASAP7_75t_SL g376 ( 
.A1(n_311),
.A2(n_315),
.B(n_321),
.C(n_328),
.Y(n_376)
);

FAx1_ASAP7_75t_SL g313 ( 
.A(n_227),
.B(n_258),
.CI(n_230),
.CON(n_313),
.SN(n_313)
);

NOR2xp33_ASAP7_75t_L g345 ( 
.A(n_313),
.B(n_332),
.Y(n_345)
);

AOI21xp5_ASAP7_75t_L g315 ( 
.A1(n_257),
.A2(n_203),
.B(n_191),
.Y(n_315)
);

OAI22xp5_ASAP7_75t_SL g318 ( 
.A1(n_229),
.A2(n_159),
.B1(n_205),
.B2(n_182),
.Y(n_318)
);

O2A1O1Ixp33_ASAP7_75t_L g321 ( 
.A1(n_219),
.A2(n_141),
.B(n_135),
.C(n_137),
.Y(n_321)
);

MAJx2_ASAP7_75t_L g323 ( 
.A(n_268),
.B(n_137),
.C(n_141),
.Y(n_323)
);

XOR2xp5_ASAP7_75t_L g359 ( 
.A(n_323),
.B(n_343),
.Y(n_359)
);

OAI22xp5_ASAP7_75t_L g372 ( 
.A1(n_326),
.A2(n_329),
.B1(n_270),
.B2(n_239),
.Y(n_372)
);

AOI22xp5_ASAP7_75t_SL g328 ( 
.A1(n_276),
.A2(n_141),
.B1(n_197),
.B2(n_180),
.Y(n_328)
);

AOI22xp5_ASAP7_75t_L g329 ( 
.A1(n_263),
.A2(n_197),
.B1(n_180),
.B2(n_5),
.Y(n_329)
);

FAx1_ASAP7_75t_SL g332 ( 
.A(n_242),
.B(n_197),
.CI(n_2),
.CON(n_332),
.SN(n_332)
);

NAND2xp5_ASAP7_75t_L g336 ( 
.A(n_223),
.B(n_1),
.Y(n_336)
);

HB1xp67_ASAP7_75t_L g377 ( 
.A(n_342),
.Y(n_377)
);

XNOR2xp5_ASAP7_75t_L g343 ( 
.A(n_279),
.B(n_5),
.Y(n_343)
);

INVx1_ASAP7_75t_SL g348 ( 
.A(n_339),
.Y(n_348)
);

AND2x2_ASAP7_75t_L g427 ( 
.A(n_348),
.B(n_360),
.Y(n_427)
);

OAI22xp5_ASAP7_75t_L g393 ( 
.A1(n_349),
.A2(n_373),
.B1(n_287),
.B2(n_308),
.Y(n_393)
);

INVx2_ASAP7_75t_L g350 ( 
.A(n_325),
.Y(n_350)
);

INVx1_ASAP7_75t_L g392 ( 
.A(n_350),
.Y(n_392)
);

INVx1_ASAP7_75t_L g351 ( 
.A(n_309),
.Y(n_351)
);

INVx1_ASAP7_75t_L g397 ( 
.A(n_351),
.Y(n_397)
);

INVx1_ASAP7_75t_L g352 ( 
.A(n_319),
.Y(n_352)
);

INVx1_ASAP7_75t_L g405 ( 
.A(n_352),
.Y(n_405)
);

NAND2xp5_ASAP7_75t_L g353 ( 
.A(n_304),
.B(n_231),
.Y(n_353)
);

NAND2xp5_ASAP7_75t_L g400 ( 
.A(n_353),
.B(n_363),
.Y(n_400)
);

INVx13_ASAP7_75t_L g354 ( 
.A(n_300),
.Y(n_354)
);

CKINVDCx14_ASAP7_75t_R g428 ( 
.A(n_354),
.Y(n_428)
);

CKINVDCx14_ASAP7_75t_R g355 ( 
.A(n_300),
.Y(n_355)
);

NOR2xp33_ASAP7_75t_L g396 ( 
.A(n_355),
.B(n_361),
.Y(n_396)
);

NOR2xp33_ASAP7_75t_L g356 ( 
.A(n_297),
.B(n_228),
.Y(n_356)
);

NAND2xp5_ASAP7_75t_SL g401 ( 
.A(n_356),
.B(n_364),
.Y(n_401)
);

OAI21xp33_ASAP7_75t_SL g358 ( 
.A1(n_327),
.A2(n_252),
.B(n_228),
.Y(n_358)
);

OAI21xp5_ASAP7_75t_SL g403 ( 
.A1(n_358),
.A2(n_382),
.B(n_385),
.Y(n_403)
);

INVx1_ASAP7_75t_SL g360 ( 
.A(n_339),
.Y(n_360)
);

AND2x6_ASAP7_75t_L g361 ( 
.A(n_313),
.B(n_228),
.Y(n_361)
);

NAND2xp5_ASAP7_75t_L g363 ( 
.A(n_304),
.B(n_265),
.Y(n_363)
);

NAND2xp5_ASAP7_75t_SL g364 ( 
.A(n_312),
.B(n_250),
.Y(n_364)
);

BUFx6f_ASAP7_75t_L g365 ( 
.A(n_330),
.Y(n_365)
);

BUFx2_ASAP7_75t_L g429 ( 
.A(n_365),
.Y(n_429)
);

AOI22xp33_ASAP7_75t_SL g366 ( 
.A1(n_318),
.A2(n_285),
.B1(n_284),
.B2(n_266),
.Y(n_366)
);

INVxp67_ASAP7_75t_L g414 ( 
.A(n_366),
.Y(n_414)
);

INVx11_ASAP7_75t_L g367 ( 
.A(n_340),
.Y(n_367)
);

INVxp67_ASAP7_75t_L g415 ( 
.A(n_367),
.Y(n_415)
);

BUFx12_ASAP7_75t_L g368 ( 
.A(n_340),
.Y(n_368)
);

CKINVDCx20_ASAP7_75t_R g391 ( 
.A(n_368),
.Y(n_391)
);

INVx3_ASAP7_75t_L g369 ( 
.A(n_330),
.Y(n_369)
);

INVx4_ASAP7_75t_L g426 ( 
.A(n_369),
.Y(n_426)
);

NAND3xp33_ASAP7_75t_L g370 ( 
.A(n_298),
.B(n_273),
.C(n_6),
.Y(n_370)
);

NAND2xp5_ASAP7_75t_SL g417 ( 
.A(n_370),
.B(n_374),
.Y(n_417)
);

OAI22xp5_ASAP7_75t_SL g371 ( 
.A1(n_326),
.A2(n_212),
.B1(n_269),
.B2(n_244),
.Y(n_371)
);

AOI22xp33_ASAP7_75t_SL g416 ( 
.A1(n_371),
.A2(n_384),
.B1(n_317),
.B2(n_325),
.Y(n_416)
);

INVx1_ASAP7_75t_L g409 ( 
.A(n_372),
.Y(n_409)
);

AOI22xp5_ASAP7_75t_L g373 ( 
.A1(n_289),
.A2(n_311),
.B1(n_333),
.B2(n_307),
.Y(n_373)
);

NOR2xp33_ASAP7_75t_L g374 ( 
.A(n_316),
.B(n_255),
.Y(n_374)
);

NOR2xp33_ASAP7_75t_L g375 ( 
.A(n_313),
.B(n_251),
.Y(n_375)
);

NAND2xp5_ASAP7_75t_SL g421 ( 
.A(n_375),
.B(n_379),
.Y(n_421)
);

INVx8_ASAP7_75t_L g378 ( 
.A(n_303),
.Y(n_378)
);

INVx1_ASAP7_75t_L g410 ( 
.A(n_378),
.Y(n_410)
);

NOR2xp33_ASAP7_75t_L g379 ( 
.A(n_327),
.B(n_218),
.Y(n_379)
);

NOR2xp33_ASAP7_75t_L g380 ( 
.A(n_293),
.B(n_224),
.Y(n_380)
);

NAND2xp5_ASAP7_75t_SL g423 ( 
.A(n_380),
.B(n_381),
.Y(n_423)
);

CKINVDCx20_ASAP7_75t_R g381 ( 
.A(n_320),
.Y(n_381)
);

OR2x2_ASAP7_75t_L g382 ( 
.A(n_332),
.B(n_5),
.Y(n_382)
);

INVx1_ASAP7_75t_L g383 ( 
.A(n_337),
.Y(n_383)
);

INVx1_ASAP7_75t_L g412 ( 
.A(n_383),
.Y(n_412)
);

OAI22xp5_ASAP7_75t_SL g384 ( 
.A1(n_311),
.A2(n_6),
.B1(n_7),
.B2(n_9),
.Y(n_384)
);

AND2x2_ASAP7_75t_L g385 ( 
.A(n_289),
.B(n_10),
.Y(n_385)
);

NAND2xp5_ASAP7_75t_L g386 ( 
.A(n_336),
.B(n_11),
.Y(n_386)
);

XNOR2xp5_ASAP7_75t_L g395 ( 
.A(n_386),
.B(n_387),
.Y(n_395)
);

NAND2xp5_ASAP7_75t_L g387 ( 
.A(n_289),
.B(n_11),
.Y(n_387)
);

CKINVDCx5p33_ASAP7_75t_R g388 ( 
.A(n_332),
.Y(n_388)
);

OAI21xp5_ASAP7_75t_L g399 ( 
.A1(n_388),
.A2(n_389),
.B(n_390),
.Y(n_399)
);

AOI22xp5_ASAP7_75t_SL g389 ( 
.A1(n_310),
.A2(n_12),
.B1(n_13),
.B2(n_14),
.Y(n_389)
);

OR2x2_ASAP7_75t_L g390 ( 
.A(n_333),
.B(n_306),
.Y(n_390)
);

AOI22xp5_ASAP7_75t_L g431 ( 
.A1(n_393),
.A2(n_394),
.B1(n_398),
.B2(n_422),
.Y(n_431)
);

OAI22xp5_ASAP7_75t_SL g394 ( 
.A1(n_373),
.A2(n_311),
.B1(n_315),
.B2(n_338),
.Y(n_394)
);

OAI22xp5_ASAP7_75t_SL g398 ( 
.A1(n_349),
.A2(n_302),
.B1(n_312),
.B2(n_343),
.Y(n_398)
);

OAI21xp5_ASAP7_75t_L g402 ( 
.A1(n_362),
.A2(n_390),
.B(n_346),
.Y(n_402)
);

AOI21xp5_ASAP7_75t_L g433 ( 
.A1(n_402),
.A2(n_419),
.B(n_388),
.Y(n_433)
);

CKINVDCx20_ASAP7_75t_R g404 ( 
.A(n_354),
.Y(n_404)
);

INVx13_ASAP7_75t_L g435 ( 
.A(n_404),
.Y(n_435)
);

XOR2xp5_ASAP7_75t_L g406 ( 
.A(n_359),
.B(n_290),
.Y(n_406)
);

XNOR2xp5_ASAP7_75t_SL g441 ( 
.A(n_406),
.B(n_411),
.Y(n_441)
);

CKINVDCx20_ASAP7_75t_R g407 ( 
.A(n_368),
.Y(n_407)
);

NOR2xp33_ASAP7_75t_L g439 ( 
.A(n_407),
.B(n_378),
.Y(n_439)
);

MAJx2_ASAP7_75t_L g408 ( 
.A(n_359),
.B(n_290),
.C(n_310),
.Y(n_408)
);

XNOR2xp5_ASAP7_75t_L g465 ( 
.A(n_408),
.B(n_413),
.Y(n_465)
);

XOR2xp5_ASAP7_75t_L g411 ( 
.A(n_387),
.B(n_290),
.Y(n_411)
);

MAJIxp5_ASAP7_75t_L g413 ( 
.A(n_362),
.B(n_323),
.C(n_339),
.Y(n_413)
);

OAI22xp33_ASAP7_75t_SL g451 ( 
.A1(n_416),
.A2(n_377),
.B1(n_357),
.B2(n_347),
.Y(n_451)
);

INVx1_ASAP7_75t_L g418 ( 
.A(n_350),
.Y(n_418)
);

INVx1_ASAP7_75t_L g437 ( 
.A(n_418),
.Y(n_437)
);

AOI21xp5_ASAP7_75t_L g419 ( 
.A1(n_362),
.A2(n_328),
.B(n_314),
.Y(n_419)
);

XOR2xp5_ASAP7_75t_L g420 ( 
.A(n_385),
.B(n_302),
.Y(n_420)
);

AND2x2_ASAP7_75t_L g436 ( 
.A(n_420),
.B(n_425),
.Y(n_436)
);

OAI22xp5_ASAP7_75t_L g422 ( 
.A1(n_347),
.A2(n_335),
.B1(n_329),
.B2(n_294),
.Y(n_422)
);

INVx1_ASAP7_75t_L g424 ( 
.A(n_352),
.Y(n_424)
);

INVx1_ASAP7_75t_L g446 ( 
.A(n_424),
.Y(n_446)
);

XOR2xp5_ASAP7_75t_L g425 ( 
.A(n_385),
.B(n_334),
.Y(n_425)
);

INVx3_ASAP7_75t_L g430 ( 
.A(n_426),
.Y(n_430)
);

INVx1_ASAP7_75t_L g476 ( 
.A(n_430),
.Y(n_476)
);

BUFx3_ASAP7_75t_L g432 ( 
.A(n_429),
.Y(n_432)
);

NOR2xp33_ASAP7_75t_L g482 ( 
.A(n_432),
.B(n_464),
.Y(n_482)
);

OAI21xp5_ASAP7_75t_L g474 ( 
.A1(n_433),
.A2(n_449),
.B(n_403),
.Y(n_474)
);

OAI21xp5_ASAP7_75t_SL g434 ( 
.A1(n_419),
.A2(n_346),
.B(n_345),
.Y(n_434)
);

OR2x2_ASAP7_75t_L g495 ( 
.A(n_434),
.B(n_459),
.Y(n_495)
);

NAND2xp5_ASAP7_75t_L g438 ( 
.A(n_400),
.B(n_353),
.Y(n_438)
);

INVx1_ASAP7_75t_L g485 ( 
.A(n_438),
.Y(n_485)
);

NAND2xp5_ASAP7_75t_L g468 ( 
.A(n_439),
.B(n_440),
.Y(n_468)
);

CKINVDCx20_ASAP7_75t_R g440 ( 
.A(n_423),
.Y(n_440)
);

CKINVDCx16_ASAP7_75t_R g442 ( 
.A(n_427),
.Y(n_442)
);

NAND2xp5_ASAP7_75t_SL g487 ( 
.A(n_442),
.B(n_444),
.Y(n_487)
);

NAND2xp5_ASAP7_75t_L g443 ( 
.A(n_400),
.B(n_363),
.Y(n_443)
);

INVx1_ASAP7_75t_L g489 ( 
.A(n_443),
.Y(n_489)
);

CKINVDCx16_ASAP7_75t_R g444 ( 
.A(n_427),
.Y(n_444)
);

CKINVDCx20_ASAP7_75t_R g445 ( 
.A(n_404),
.Y(n_445)
);

NAND2xp5_ASAP7_75t_L g469 ( 
.A(n_445),
.B(n_453),
.Y(n_469)
);

INVx1_ASAP7_75t_L g447 ( 
.A(n_405),
.Y(n_447)
);

INVx1_ASAP7_75t_L g490 ( 
.A(n_447),
.Y(n_490)
);

INVx1_ASAP7_75t_L g448 ( 
.A(n_405),
.Y(n_448)
);

INVx1_ASAP7_75t_L g491 ( 
.A(n_448),
.Y(n_491)
);

AOI21xp5_ASAP7_75t_L g449 ( 
.A1(n_402),
.A2(n_414),
.B(n_396),
.Y(n_449)
);

NAND2xp5_ASAP7_75t_L g450 ( 
.A(n_397),
.B(n_386),
.Y(n_450)
);

INVx1_ASAP7_75t_L g497 ( 
.A(n_450),
.Y(n_497)
);

AOI22xp5_ASAP7_75t_L g478 ( 
.A1(n_451),
.A2(n_452),
.B1(n_414),
.B2(n_376),
.Y(n_478)
);

OAI22xp5_ASAP7_75t_L g452 ( 
.A1(n_409),
.A2(n_357),
.B1(n_384),
.B2(n_348),
.Y(n_452)
);

INVx1_ASAP7_75t_L g453 ( 
.A(n_412),
.Y(n_453)
);

NAND2xp5_ASAP7_75t_SL g454 ( 
.A(n_397),
.B(n_381),
.Y(n_454)
);

NAND2xp5_ASAP7_75t_SL g493 ( 
.A(n_454),
.B(n_460),
.Y(n_493)
);

INVx1_ASAP7_75t_L g455 ( 
.A(n_412),
.Y(n_455)
);

NAND2xp5_ASAP7_75t_L g475 ( 
.A(n_455),
.B(n_456),
.Y(n_475)
);

CKINVDCx20_ASAP7_75t_R g456 ( 
.A(n_428),
.Y(n_456)
);

CKINVDCx20_ASAP7_75t_R g457 ( 
.A(n_401),
.Y(n_457)
);

NAND2xp5_ASAP7_75t_L g477 ( 
.A(n_457),
.B(n_458),
.Y(n_477)
);

INVx1_ASAP7_75t_L g458 ( 
.A(n_424),
.Y(n_458)
);

NOR2xp33_ASAP7_75t_SL g459 ( 
.A(n_421),
.B(n_351),
.Y(n_459)
);

NAND2xp5_ASAP7_75t_SL g460 ( 
.A(n_398),
.B(n_383),
.Y(n_460)
);

INVx2_ASAP7_75t_L g461 ( 
.A(n_392),
.Y(n_461)
);

NAND2xp5_ASAP7_75t_L g480 ( 
.A(n_461),
.B(n_462),
.Y(n_480)
);

NAND2xp5_ASAP7_75t_L g462 ( 
.A(n_392),
.B(n_360),
.Y(n_462)
);

CKINVDCx10_ASAP7_75t_R g463 ( 
.A(n_415),
.Y(n_463)
);

CKINVDCx20_ASAP7_75t_R g498 ( 
.A(n_463),
.Y(n_498)
);

NOR2x1_ASAP7_75t_L g464 ( 
.A(n_413),
.B(n_361),
.Y(n_464)
);

BUFx24_ASAP7_75t_SL g466 ( 
.A(n_459),
.Y(n_466)
);

NOR2xp33_ASAP7_75t_L g506 ( 
.A(n_466),
.B(n_395),
.Y(n_506)
);

NOR2xp33_ASAP7_75t_SL g467 ( 
.A(n_440),
.B(n_399),
.Y(n_467)
);

NAND3xp33_ASAP7_75t_L g521 ( 
.A(n_467),
.B(n_479),
.C(n_486),
.Y(n_521)
);

OA21x2_ASAP7_75t_L g470 ( 
.A1(n_431),
.A2(n_394),
.B(n_409),
.Y(n_470)
);

AOI22xp5_ASAP7_75t_L g508 ( 
.A1(n_470),
.A2(n_372),
.B1(n_371),
.B2(n_376),
.Y(n_508)
);

XOR2xp5_ASAP7_75t_L g471 ( 
.A(n_441),
.B(n_406),
.Y(n_471)
);

XOR2xp5_ASAP7_75t_L g516 ( 
.A(n_471),
.B(n_472),
.Y(n_516)
);

XNOR2xp5_ASAP7_75t_L g472 ( 
.A(n_441),
.B(n_408),
.Y(n_472)
);

AO21x1_ASAP7_75t_L g473 ( 
.A1(n_464),
.A2(n_399),
.B(n_427),
.Y(n_473)
);

AOI21xp5_ASAP7_75t_L g520 ( 
.A1(n_473),
.A2(n_474),
.B(n_487),
.Y(n_520)
);

OAI22xp5_ASAP7_75t_L g523 ( 
.A1(n_478),
.A2(n_376),
.B1(n_430),
.B2(n_426),
.Y(n_523)
);

NOR2xp33_ASAP7_75t_SL g479 ( 
.A(n_457),
.B(n_417),
.Y(n_479)
);

MAJIxp5_ASAP7_75t_L g481 ( 
.A(n_465),
.B(n_411),
.C(n_420),
.Y(n_481)
);

MAJIxp5_ASAP7_75t_L g511 ( 
.A(n_481),
.B(n_448),
.C(n_458),
.Y(n_511)
);

XNOR2xp5_ASAP7_75t_SL g483 ( 
.A(n_465),
.B(n_425),
.Y(n_483)
);

XNOR2xp5_ASAP7_75t_SL g526 ( 
.A(n_483),
.B(n_435),
.Y(n_526)
);

OAI22xp5_ASAP7_75t_L g484 ( 
.A1(n_431),
.A2(n_382),
.B1(n_389),
.B2(n_410),
.Y(n_484)
);

INVx1_ASAP7_75t_L g503 ( 
.A(n_484),
.Y(n_503)
);

NOR2xp33_ASAP7_75t_L g486 ( 
.A(n_456),
.B(n_410),
.Y(n_486)
);

OAI22xp5_ASAP7_75t_L g488 ( 
.A1(n_449),
.A2(n_418),
.B1(n_376),
.B2(n_415),
.Y(n_488)
);

INVx1_ASAP7_75t_L g504 ( 
.A(n_488),
.Y(n_504)
);

XNOR2xp5_ASAP7_75t_L g492 ( 
.A(n_436),
.B(n_395),
.Y(n_492)
);

XOR2xp5_ASAP7_75t_L g527 ( 
.A(n_492),
.B(n_292),
.Y(n_527)
);

NOR2xp33_ASAP7_75t_L g494 ( 
.A(n_450),
.B(n_407),
.Y(n_494)
);

INVx1_ASAP7_75t_L g509 ( 
.A(n_494),
.Y(n_509)
);

NAND2xp5_ASAP7_75t_L g496 ( 
.A(n_438),
.B(n_391),
.Y(n_496)
);

INVx1_ASAP7_75t_L g515 ( 
.A(n_496),
.Y(n_515)
);

OAI22xp5_ASAP7_75t_SL g499 ( 
.A1(n_478),
.A2(n_433),
.B1(n_443),
.B2(n_442),
.Y(n_499)
);

AOI22xp5_ASAP7_75t_L g552 ( 
.A1(n_499),
.A2(n_523),
.B1(n_367),
.B2(n_365),
.Y(n_552)
);

INVx3_ASAP7_75t_L g500 ( 
.A(n_476),
.Y(n_500)
);

INVx1_ASAP7_75t_L g530 ( 
.A(n_500),
.Y(n_530)
);

AOI22xp5_ASAP7_75t_SL g501 ( 
.A1(n_467),
.A2(n_444),
.B1(n_436),
.B2(n_452),
.Y(n_501)
);

OAI22xp5_ASAP7_75t_SL g531 ( 
.A1(n_501),
.A2(n_514),
.B1(n_525),
.B2(n_475),
.Y(n_531)
);

OAI21xp5_ASAP7_75t_SL g502 ( 
.A1(n_482),
.A2(n_445),
.B(n_462),
.Y(n_502)
);

INVx1_ASAP7_75t_L g547 ( 
.A(n_502),
.Y(n_547)
);

OAI21xp5_ASAP7_75t_SL g505 ( 
.A1(n_495),
.A2(n_463),
.B(n_434),
.Y(n_505)
);

NOR2xp33_ASAP7_75t_L g536 ( 
.A(n_505),
.B(n_506),
.Y(n_536)
);

XNOR2xp5_ASAP7_75t_L g507 ( 
.A(n_492),
.B(n_436),
.Y(n_507)
);

XOR2xp5_ASAP7_75t_L g529 ( 
.A(n_507),
.B(n_511),
.Y(n_529)
);

OAI22xp5_ASAP7_75t_L g543 ( 
.A1(n_508),
.A2(n_498),
.B1(n_491),
.B2(n_490),
.Y(n_543)
);

FAx1_ASAP7_75t_SL g510 ( 
.A(n_495),
.B(n_403),
.CI(n_376),
.CON(n_510),
.SN(n_510)
);

NOR2xp33_ASAP7_75t_L g551 ( 
.A(n_510),
.B(n_518),
.Y(n_551)
);

MAJIxp5_ASAP7_75t_L g512 ( 
.A(n_481),
.B(n_391),
.C(n_437),
.Y(n_512)
);

MAJIxp5_ASAP7_75t_L g532 ( 
.A(n_512),
.B(n_513),
.C(n_517),
.Y(n_532)
);

MAJIxp5_ASAP7_75t_L g513 ( 
.A(n_471),
.B(n_483),
.C(n_472),
.Y(n_513)
);

AOI22xp5_ASAP7_75t_L g514 ( 
.A1(n_470),
.A2(n_447),
.B1(n_455),
.B2(n_446),
.Y(n_514)
);

MAJIxp5_ASAP7_75t_L g517 ( 
.A(n_473),
.B(n_437),
.C(n_461),
.Y(n_517)
);

OAI22xp5_ASAP7_75t_SL g518 ( 
.A1(n_493),
.A2(n_497),
.B1(n_479),
.B2(n_477),
.Y(n_518)
);

CKINVDCx20_ASAP7_75t_R g519 ( 
.A(n_469),
.Y(n_519)
);

CKINVDCx20_ASAP7_75t_R g541 ( 
.A(n_519),
.Y(n_541)
);

OAI21xp5_ASAP7_75t_SL g540 ( 
.A1(n_520),
.A2(n_468),
.B(n_477),
.Y(n_540)
);

MAJIxp5_ASAP7_75t_L g522 ( 
.A(n_473),
.B(n_453),
.C(n_446),
.Y(n_522)
);

MAJIxp5_ASAP7_75t_L g535 ( 
.A(n_522),
.B(n_527),
.C(n_475),
.Y(n_535)
);

XNOR2xp5_ASAP7_75t_L g524 ( 
.A(n_474),
.B(n_292),
.Y(n_524)
);

XOR2xp5_ASAP7_75t_L g534 ( 
.A(n_524),
.B(n_526),
.Y(n_534)
);

AOI22xp5_ASAP7_75t_L g525 ( 
.A1(n_470),
.A2(n_429),
.B1(n_432),
.B2(n_435),
.Y(n_525)
);

INVx1_ASAP7_75t_L g528 ( 
.A(n_469),
.Y(n_528)
);

INVx1_ASAP7_75t_L g544 ( 
.A(n_528),
.Y(n_544)
);

AOI22xp33_ASAP7_75t_SL g566 ( 
.A1(n_531),
.A2(n_514),
.B1(n_510),
.B2(n_521),
.Y(n_566)
);

OAI22xp5_ASAP7_75t_SL g533 ( 
.A1(n_504),
.A2(n_497),
.B1(n_489),
.B2(n_485),
.Y(n_533)
);

AOI22xp5_ASAP7_75t_L g569 ( 
.A1(n_533),
.A2(n_537),
.B1(n_543),
.B2(n_545),
.Y(n_569)
);

MAJx2_ASAP7_75t_L g568 ( 
.A(n_535),
.B(n_553),
.C(n_331),
.Y(n_568)
);

OAI22xp5_ASAP7_75t_SL g537 ( 
.A1(n_503),
.A2(n_489),
.B1(n_485),
.B2(n_496),
.Y(n_537)
);

MAJIxp5_ASAP7_75t_L g538 ( 
.A(n_512),
.B(n_468),
.C(n_480),
.Y(n_538)
);

NAND2xp5_ASAP7_75t_L g558 ( 
.A(n_538),
.B(n_539),
.Y(n_558)
);

CKINVDCx16_ASAP7_75t_R g539 ( 
.A(n_522),
.Y(n_539)
);

AOI21xp5_ASAP7_75t_L g557 ( 
.A1(n_540),
.A2(n_517),
.B(n_524),
.Y(n_557)
);

MAJIxp5_ASAP7_75t_L g542 ( 
.A(n_511),
.B(n_480),
.C(n_498),
.Y(n_542)
);

MAJIxp5_ASAP7_75t_L g573 ( 
.A(n_542),
.B(n_546),
.C(n_548),
.Y(n_573)
);

OAI22xp5_ASAP7_75t_SL g545 ( 
.A1(n_501),
.A2(n_491),
.B1(n_490),
.B2(n_476),
.Y(n_545)
);

MAJIxp5_ASAP7_75t_L g546 ( 
.A(n_516),
.B(n_527),
.C(n_507),
.Y(n_546)
);

MAJIxp5_ASAP7_75t_L g548 ( 
.A(n_516),
.B(n_369),
.C(n_288),
.Y(n_548)
);

INVx1_ASAP7_75t_L g549 ( 
.A(n_515),
.Y(n_549)
);

INVx1_ASAP7_75t_L g556 ( 
.A(n_549),
.Y(n_556)
);

MAJIxp5_ASAP7_75t_L g550 ( 
.A(n_513),
.B(n_288),
.C(n_331),
.Y(n_550)
);

NOR2xp33_ASAP7_75t_L g565 ( 
.A(n_550),
.B(n_500),
.Y(n_565)
);

OAI22xp5_ASAP7_75t_SL g555 ( 
.A1(n_552),
.A2(n_508),
.B1(n_525),
.B2(n_509),
.Y(n_555)
);

XOR2xp5_ASAP7_75t_SL g553 ( 
.A(n_499),
.B(n_368),
.Y(n_553)
);

CKINVDCx16_ASAP7_75t_R g554 ( 
.A(n_542),
.Y(n_554)
);

NAND2xp5_ASAP7_75t_SL g589 ( 
.A(n_554),
.B(n_563),
.Y(n_589)
);

INVx1_ASAP7_75t_L g574 ( 
.A(n_555),
.Y(n_574)
);

AOI21xp5_ASAP7_75t_L g584 ( 
.A1(n_557),
.A2(n_534),
.B(n_529),
.Y(n_584)
);

INVx1_ASAP7_75t_L g559 ( 
.A(n_537),
.Y(n_559)
);

INVx1_ASAP7_75t_L g575 ( 
.A(n_559),
.Y(n_575)
);

INVxp67_ASAP7_75t_SL g560 ( 
.A(n_547),
.Y(n_560)
);

INVx1_ASAP7_75t_L g579 ( 
.A(n_560),
.Y(n_579)
);

INVx1_ASAP7_75t_L g561 ( 
.A(n_530),
.Y(n_561)
);

INVx1_ASAP7_75t_L g580 ( 
.A(n_561),
.Y(n_580)
);

XNOR2xp5_ASAP7_75t_L g562 ( 
.A(n_532),
.B(n_526),
.Y(n_562)
);

XNOR2xp5_ASAP7_75t_L g582 ( 
.A(n_562),
.B(n_565),
.Y(n_582)
);

BUFx24_ASAP7_75t_SL g563 ( 
.A(n_536),
.Y(n_563)
);

INVxp67_ASAP7_75t_L g564 ( 
.A(n_540),
.Y(n_564)
);

INVx1_ASAP7_75t_L g583 ( 
.A(n_564),
.Y(n_583)
);

HB1xp67_ASAP7_75t_L g578 ( 
.A(n_566),
.Y(n_578)
);

FAx1_ASAP7_75t_SL g567 ( 
.A(n_538),
.B(n_510),
.CI(n_368),
.CON(n_567),
.SN(n_567)
);

MAJx2_ASAP7_75t_L g581 ( 
.A(n_567),
.B(n_568),
.C(n_550),
.Y(n_581)
);

XOR2xp5_ASAP7_75t_L g570 ( 
.A(n_546),
.B(n_331),
.Y(n_570)
);

XNOR2xp5_ASAP7_75t_L g590 ( 
.A(n_570),
.B(n_572),
.Y(n_590)
);

BUFx24_ASAP7_75t_SL g571 ( 
.A(n_541),
.Y(n_571)
);

INVx1_ASAP7_75t_L g587 ( 
.A(n_571),
.Y(n_587)
);

XOR2xp5_ASAP7_75t_L g572 ( 
.A(n_532),
.B(n_324),
.Y(n_572)
);

AOI21x1_ASAP7_75t_L g576 ( 
.A1(n_564),
.A2(n_551),
.B(n_535),
.Y(n_576)
);

OAI21xp5_ASAP7_75t_L g600 ( 
.A1(n_576),
.A2(n_567),
.B(n_544),
.Y(n_600)
);

MAJIxp5_ASAP7_75t_L g577 ( 
.A(n_573),
.B(n_529),
.C(n_548),
.Y(n_577)
);

NAND2xp5_ASAP7_75t_L g595 ( 
.A(n_577),
.B(n_562),
.Y(n_595)
);

XNOR2xp5_ASAP7_75t_L g597 ( 
.A(n_581),
.B(n_568),
.Y(n_597)
);

AOI21xp5_ASAP7_75t_L g604 ( 
.A1(n_584),
.A2(n_585),
.B(n_530),
.Y(n_604)
);

OAI21xp5_ASAP7_75t_SL g585 ( 
.A1(n_558),
.A2(n_544),
.B(n_549),
.Y(n_585)
);

AOI22xp5_ASAP7_75t_SL g586 ( 
.A1(n_567),
.A2(n_531),
.B1(n_545),
.B2(n_533),
.Y(n_586)
);

XNOR2xp5_ASAP7_75t_L g598 ( 
.A(n_586),
.B(n_553),
.Y(n_598)
);

INVx1_ASAP7_75t_L g588 ( 
.A(n_556),
.Y(n_588)
);

INVx1_ASAP7_75t_L g591 ( 
.A(n_588),
.Y(n_591)
);

NAND2xp5_ASAP7_75t_SL g592 ( 
.A(n_589),
.B(n_573),
.Y(n_592)
);

NAND2xp5_ASAP7_75t_L g606 ( 
.A(n_592),
.B(n_593),
.Y(n_606)
);

MAJIxp5_ASAP7_75t_L g593 ( 
.A(n_577),
.B(n_572),
.C(n_570),
.Y(n_593)
);

NOR2xp33_ASAP7_75t_L g594 ( 
.A(n_582),
.B(n_569),
.Y(n_594)
);

NAND2xp5_ASAP7_75t_L g610 ( 
.A(n_594),
.B(n_595),
.Y(n_610)
);

NAND2xp5_ASAP7_75t_L g596 ( 
.A(n_580),
.B(n_583),
.Y(n_596)
);

NAND2xp5_ASAP7_75t_SL g614 ( 
.A(n_596),
.B(n_599),
.Y(n_614)
);

AOI21xp5_ASAP7_75t_L g607 ( 
.A1(n_597),
.A2(n_600),
.B(n_601),
.Y(n_607)
);

XNOR2xp5_ASAP7_75t_L g612 ( 
.A(n_598),
.B(n_322),
.Y(n_612)
);

XNOR2xp5_ASAP7_75t_L g599 ( 
.A(n_582),
.B(n_534),
.Y(n_599)
);

MAJIxp5_ASAP7_75t_L g601 ( 
.A(n_574),
.B(n_590),
.C(n_584),
.Y(n_601)
);

AND2x2_ASAP7_75t_L g602 ( 
.A(n_578),
.B(n_552),
.Y(n_602)
);

AOI22xp5_ASAP7_75t_L g608 ( 
.A1(n_602),
.A2(n_586),
.B1(n_581),
.B2(n_590),
.Y(n_608)
);

NOR2xp33_ASAP7_75t_L g603 ( 
.A(n_579),
.B(n_575),
.Y(n_603)
);

NOR2xp33_ASAP7_75t_SL g609 ( 
.A(n_603),
.B(n_604),
.Y(n_609)
);

HB1xp67_ASAP7_75t_L g605 ( 
.A(n_601),
.Y(n_605)
);

CKINVDCx20_ASAP7_75t_R g619 ( 
.A(n_605),
.Y(n_619)
);

NAND2xp33_ASAP7_75t_SL g616 ( 
.A(n_608),
.B(n_611),
.Y(n_616)
);

OA21x2_ASAP7_75t_SL g611 ( 
.A1(n_591),
.A2(n_587),
.B(n_324),
.Y(n_611)
);

INVxp67_ASAP7_75t_L g617 ( 
.A(n_612),
.Y(n_617)
);

MAJIxp5_ASAP7_75t_L g613 ( 
.A(n_593),
.B(n_322),
.C(n_341),
.Y(n_613)
);

NOR2xp33_ASAP7_75t_L g618 ( 
.A(n_613),
.B(n_341),
.Y(n_618)
);

AOI22xp5_ASAP7_75t_SL g615 ( 
.A1(n_605),
.A2(n_602),
.B1(n_598),
.B2(n_317),
.Y(n_615)
);

AOI21xp5_ASAP7_75t_L g624 ( 
.A1(n_615),
.A2(n_616),
.B(n_613),
.Y(n_624)
);

NAND2xp5_ASAP7_75t_SL g622 ( 
.A(n_618),
.B(n_621),
.Y(n_622)
);

O2A1O1Ixp33_ASAP7_75t_L g620 ( 
.A1(n_607),
.A2(n_344),
.B(n_14),
.C(n_12),
.Y(n_620)
);

OR2x2_ASAP7_75t_L g623 ( 
.A(n_620),
.B(n_609),
.Y(n_623)
);

NOR2xp33_ASAP7_75t_L g621 ( 
.A(n_614),
.B(n_344),
.Y(n_621)
);

INVx1_ASAP7_75t_L g627 ( 
.A(n_623),
.Y(n_627)
);

AOI322xp5_ASAP7_75t_L g626 ( 
.A1(n_624),
.A2(n_625),
.A3(n_622),
.B1(n_617),
.B2(n_620),
.C1(n_286),
.C2(n_299),
.Y(n_626)
);

MAJIxp5_ASAP7_75t_L g625 ( 
.A(n_619),
.B(n_606),
.C(n_610),
.Y(n_625)
);

BUFx24_ASAP7_75t_SL g628 ( 
.A(n_626),
.Y(n_628)
);

MAJIxp5_ASAP7_75t_L g629 ( 
.A(n_628),
.B(n_627),
.C(n_286),
.Y(n_629)
);

INVx1_ASAP7_75t_L g630 ( 
.A(n_629),
.Y(n_630)
);

MAJx2_ASAP7_75t_L g631 ( 
.A(n_630),
.B(n_299),
.C(n_12),
.Y(n_631)
);

CKINVDCx20_ASAP7_75t_R g632 ( 
.A(n_631),
.Y(n_632)
);


endmodule