module fake_jpeg_7191_n_297 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_297);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_297;

wire n_159;
wire n_117;
wire n_253;
wire n_286;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_251;
wire n_252;
wire n_273;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_279;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_278;
wire n_205;
wire n_295;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_293;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_281;
wire n_31;
wire n_155;
wire n_207;
wire n_277;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_291;
wire n_236;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_223;
wire n_21;
wire n_57;
wire n_187;
wire n_234;
wire n_284;
wire n_272;
wire n_288;
wire n_280;
wire n_171;
wire n_263;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_289;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_267;
wire n_248;
wire n_30;
wire n_296;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_274;
wire n_186;
wire n_24;
wire n_44;
wire n_276;
wire n_143;
wire n_202;
wire n_25;
wire n_17;
wire n_269;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_287;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_266;
wire n_34;
wire n_283;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_285;
wire n_215;
wire n_262;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_294;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_271;
wire n_217;
wire n_216;
wire n_264;
wire n_184;
wire n_53;
wire n_268;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_265;
wire n_176;
wire n_199;
wire n_112;
wire n_260;
wire n_270;
wire n_222;
wire n_95;
wire n_275;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_290;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_292;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_118;
wire n_100;
wire n_82;
wire n_128;
wire n_140;
wire n_258;
wire n_282;
wire n_96;

BUFx6f_ASAP7_75t_L g17 ( 
.A(n_11),
.Y(n_17)
);

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_0),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_16),
.Y(n_19)
);

INVx3_ASAP7_75t_L g20 ( 
.A(n_2),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_12),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_12),
.Y(n_22)
);

BUFx24_ASAP7_75t_L g23 ( 
.A(n_8),
.Y(n_23)
);

BUFx12f_ASAP7_75t_L g24 ( 
.A(n_6),
.Y(n_24)
);

BUFx10_ASAP7_75t_L g25 ( 
.A(n_7),
.Y(n_25)
);

BUFx3_ASAP7_75t_L g26 ( 
.A(n_16),
.Y(n_26)
);

INVx2_ASAP7_75t_L g27 ( 
.A(n_9),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_13),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_14),
.Y(n_29)
);

BUFx12_ASAP7_75t_L g30 ( 
.A(n_14),
.Y(n_30)
);

BUFx3_ASAP7_75t_L g31 ( 
.A(n_14),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_7),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_3),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_10),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_L g35 ( 
.A(n_19),
.B(n_15),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_SL g54 ( 
.A(n_35),
.B(n_21),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_24),
.Y(n_36)
);

INVx3_ASAP7_75t_L g65 ( 
.A(n_36),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_SL g37 ( 
.A(n_27),
.B(n_0),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g46 ( 
.A(n_37),
.B(n_39),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_L g38 ( 
.A(n_27),
.B(n_0),
.Y(n_38)
);

NAND2xp5_ASAP7_75t_L g58 ( 
.A(n_38),
.B(n_33),
.Y(n_58)
);

INVx2_ASAP7_75t_L g39 ( 
.A(n_25),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_24),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_40),
.Y(n_62)
);

INVx8_ASAP7_75t_L g41 ( 
.A(n_23),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g47 ( 
.A(n_41),
.B(n_44),
.Y(n_47)
);

INVx6_ASAP7_75t_SL g42 ( 
.A(n_26),
.Y(n_42)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_42),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_24),
.Y(n_43)
);

INVx5_ASAP7_75t_L g53 ( 
.A(n_43),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_SL g44 ( 
.A(n_23),
.B(n_1),
.Y(n_44)
);

INVx2_ASAP7_75t_L g45 ( 
.A(n_42),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_45),
.B(n_48),
.Y(n_82)
);

INVx2_ASAP7_75t_L g48 ( 
.A(n_42),
.Y(n_48)
);

INVx2_ASAP7_75t_L g49 ( 
.A(n_39),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_49),
.B(n_54),
.Y(n_74)
);

AOI22xp33_ASAP7_75t_SL g50 ( 
.A1(n_41),
.A2(n_20),
.B1(n_28),
.B2(n_21),
.Y(n_50)
);

INVxp67_ASAP7_75t_L g87 ( 
.A(n_50),
.Y(n_87)
);

OAI22xp5_ASAP7_75t_SL g51 ( 
.A1(n_38),
.A2(n_37),
.B1(n_20),
.B2(n_44),
.Y(n_51)
);

AOI22xp5_ASAP7_75t_L g88 ( 
.A1(n_51),
.A2(n_18),
.B1(n_17),
.B2(n_25),
.Y(n_88)
);

INVx4_ASAP7_75t_L g52 ( 
.A(n_39),
.Y(n_52)
);

INVx4_ASAP7_75t_L g76 ( 
.A(n_52),
.Y(n_76)
);

AOI22xp33_ASAP7_75t_SL g55 ( 
.A1(n_41),
.A2(n_28),
.B1(n_32),
.B2(n_34),
.Y(n_55)
);

OAI22xp5_ASAP7_75t_SL g78 ( 
.A1(n_55),
.A2(n_64),
.B1(n_68),
.B2(n_69),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_38),
.B(n_19),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_SL g75 ( 
.A(n_56),
.B(n_57),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g57 ( 
.A(n_37),
.B(n_34),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_L g73 ( 
.A(n_58),
.B(n_67),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_35),
.B(n_44),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_60),
.B(n_61),
.Y(n_86)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_36),
.Y(n_61)
);

AOI22xp33_ASAP7_75t_SL g63 ( 
.A1(n_41),
.A2(n_22),
.B1(n_32),
.B2(n_26),
.Y(n_63)
);

INVxp67_ASAP7_75t_L g91 ( 
.A(n_63),
.Y(n_91)
);

OAI22xp5_ASAP7_75t_L g64 ( 
.A1(n_36),
.A2(n_22),
.B1(n_17),
.B2(n_29),
.Y(n_64)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_36),
.Y(n_66)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_66),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g67 ( 
.A(n_43),
.B(n_24),
.Y(n_67)
);

AOI22xp33_ASAP7_75t_SL g68 ( 
.A1(n_36),
.A2(n_26),
.B1(n_31),
.B2(n_29),
.Y(n_68)
);

AOI22xp33_ASAP7_75t_SL g69 ( 
.A1(n_40),
.A2(n_31),
.B1(n_33),
.B2(n_29),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_SL g70 ( 
.A(n_40),
.B(n_30),
.Y(n_70)
);

CKINVDCx20_ASAP7_75t_R g94 ( 
.A(n_70),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_L g71 ( 
.A(n_40),
.B(n_33),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_71),
.B(n_18),
.Y(n_89)
);

AND2x2_ASAP7_75t_SL g72 ( 
.A(n_58),
.B(n_43),
.Y(n_72)
);

MAJIxp5_ASAP7_75t_L g112 ( 
.A(n_72),
.B(n_90),
.C(n_70),
.Y(n_112)
);

BUFx2_ASAP7_75t_L g77 ( 
.A(n_62),
.Y(n_77)
);

CKINVDCx20_ASAP7_75t_R g97 ( 
.A(n_77),
.Y(n_97)
);

INVx5_ASAP7_75t_L g79 ( 
.A(n_53),
.Y(n_79)
);

INVx2_ASAP7_75t_L g106 ( 
.A(n_79),
.Y(n_106)
);

INVx2_ASAP7_75t_L g80 ( 
.A(n_53),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_80),
.B(n_81),
.Y(n_105)
);

INVx5_ASAP7_75t_SL g81 ( 
.A(n_53),
.Y(n_81)
);

INVx2_ASAP7_75t_L g83 ( 
.A(n_64),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g116 ( 
.A(n_83),
.B(n_93),
.Y(n_116)
);

BUFx3_ASAP7_75t_L g85 ( 
.A(n_61),
.Y(n_85)
);

INVx8_ASAP7_75t_L g111 ( 
.A(n_85),
.Y(n_111)
);

XNOR2xp5_ASAP7_75t_L g120 ( 
.A(n_88),
.B(n_18),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_L g103 ( 
.A(n_89),
.B(n_56),
.Y(n_103)
);

MAJIxp5_ASAP7_75t_L g90 ( 
.A(n_51),
.B(n_43),
.C(n_40),
.Y(n_90)
);

BUFx6f_ASAP7_75t_L g92 ( 
.A(n_62),
.Y(n_92)
);

INVx2_ASAP7_75t_L g114 ( 
.A(n_92),
.Y(n_114)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_71),
.Y(n_93)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_86),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g143 ( 
.A(n_95),
.B(n_96),
.Y(n_143)
);

CKINVDCx11_ASAP7_75t_R g96 ( 
.A(n_81),
.Y(n_96)
);

CKINVDCx20_ASAP7_75t_R g98 ( 
.A(n_77),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g121 ( 
.A(n_98),
.B(n_107),
.Y(n_121)
);

OAI22xp5_ASAP7_75t_SL g99 ( 
.A1(n_90),
.A2(n_69),
.B1(n_46),
.B2(n_55),
.Y(n_99)
);

OAI22xp5_ASAP7_75t_SL g123 ( 
.A1(n_99),
.A2(n_109),
.B1(n_118),
.B2(n_87),
.Y(n_123)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_86),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_SL g132 ( 
.A(n_100),
.B(n_103),
.Y(n_132)
);

OAI21xp5_ASAP7_75t_L g101 ( 
.A1(n_91),
.A2(n_47),
.B(n_46),
.Y(n_101)
);

OAI21xp5_ASAP7_75t_SL g136 ( 
.A1(n_101),
.A2(n_102),
.B(n_75),
.Y(n_136)
);

AND2x2_ASAP7_75t_L g102 ( 
.A(n_93),
.B(n_47),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_L g104 ( 
.A(n_73),
.B(n_72),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_SL g138 ( 
.A(n_104),
.B(n_108),
.Y(n_138)
);

CKINVDCx20_ASAP7_75t_R g107 ( 
.A(n_77),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_L g108 ( 
.A(n_73),
.B(n_60),
.Y(n_108)
);

OAI22xp5_ASAP7_75t_SL g109 ( 
.A1(n_88),
.A2(n_67),
.B1(n_52),
.B2(n_59),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_L g110 ( 
.A(n_72),
.B(n_57),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_SL g139 ( 
.A(n_110),
.B(n_113),
.Y(n_139)
);

MAJIxp5_ASAP7_75t_L g141 ( 
.A(n_112),
.B(n_84),
.C(n_76),
.Y(n_141)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_74),
.Y(n_113)
);

OA22x2_ASAP7_75t_L g115 ( 
.A1(n_78),
.A2(n_65),
.B1(n_43),
.B2(n_66),
.Y(n_115)
);

A2O1A1Ixp33_ASAP7_75t_SL g147 ( 
.A1(n_115),
.A2(n_117),
.B(n_84),
.C(n_79),
.Y(n_147)
);

OAI22xp5_ASAP7_75t_L g117 ( 
.A1(n_83),
.A2(n_49),
.B1(n_59),
.B2(n_48),
.Y(n_117)
);

AOI22xp33_ASAP7_75t_L g118 ( 
.A1(n_78),
.A2(n_52),
.B1(n_65),
.B2(n_45),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_L g119 ( 
.A(n_72),
.B(n_54),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_SL g144 ( 
.A(n_119),
.B(n_120),
.Y(n_144)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_105),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_SL g155 ( 
.A(n_122),
.B(n_126),
.Y(n_155)
);

AOI22xp5_ASAP7_75t_L g151 ( 
.A1(n_123),
.A2(n_125),
.B1(n_147),
.B2(n_113),
.Y(n_151)
);

OAI21xp5_ASAP7_75t_L g124 ( 
.A1(n_101),
.A2(n_94),
.B(n_74),
.Y(n_124)
);

OAI21xp5_ASAP7_75t_SL g159 ( 
.A1(n_124),
.A2(n_134),
.B(n_25),
.Y(n_159)
);

OAI22xp5_ASAP7_75t_SL g125 ( 
.A1(n_112),
.A2(n_89),
.B1(n_94),
.B2(n_81),
.Y(n_125)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_116),
.Y(n_126)
);

CKINVDCx16_ASAP7_75t_R g127 ( 
.A(n_96),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_L g161 ( 
.A(n_127),
.B(n_135),
.Y(n_161)
);

INVxp67_ASAP7_75t_L g128 ( 
.A(n_99),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_SL g165 ( 
.A(n_128),
.B(n_129),
.Y(n_165)
);

INVxp67_ASAP7_75t_L g129 ( 
.A(n_109),
.Y(n_129)
);

BUFx2_ASAP7_75t_L g130 ( 
.A(n_106),
.Y(n_130)
);

CKINVDCx20_ASAP7_75t_R g148 ( 
.A(n_130),
.Y(n_148)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_115),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_SL g170 ( 
.A(n_131),
.B(n_133),
.Y(n_170)
);

INVxp67_ASAP7_75t_L g133 ( 
.A(n_106),
.Y(n_133)
);

HAxp5_ASAP7_75t_SL g134 ( 
.A(n_119),
.B(n_75),
.CON(n_134),
.SN(n_134)
);

CKINVDCx20_ASAP7_75t_R g135 ( 
.A(n_102),
.Y(n_135)
);

AOI21xp5_ASAP7_75t_L g149 ( 
.A1(n_136),
.A2(n_95),
.B(n_100),
.Y(n_149)
);

XOR2xp5_ASAP7_75t_L g137 ( 
.A(n_104),
.B(n_82),
.Y(n_137)
);

XOR2xp5_ASAP7_75t_L g153 ( 
.A(n_137),
.B(n_141),
.Y(n_153)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_115),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_SL g171 ( 
.A(n_140),
.B(n_142),
.Y(n_171)
);

INVxp67_ASAP7_75t_L g142 ( 
.A(n_111),
.Y(n_142)
);

CKINVDCx20_ASAP7_75t_R g145 ( 
.A(n_102),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_L g168 ( 
.A(n_145),
.B(n_146),
.Y(n_168)
);

CKINVDCx20_ASAP7_75t_R g146 ( 
.A(n_108),
.Y(n_146)
);

OAI21xp5_ASAP7_75t_SL g184 ( 
.A1(n_149),
.A2(n_151),
.B(n_145),
.Y(n_184)
);

CKINVDCx20_ASAP7_75t_R g150 ( 
.A(n_121),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_SL g182 ( 
.A(n_150),
.B(n_162),
.Y(n_182)
);

NOR2xp33_ASAP7_75t_SL g152 ( 
.A(n_146),
.B(n_103),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_SL g192 ( 
.A(n_152),
.B(n_159),
.Y(n_192)
);

AOI22xp5_ASAP7_75t_L g154 ( 
.A1(n_123),
.A2(n_115),
.B1(n_120),
.B2(n_110),
.Y(n_154)
);

AOI22xp5_ASAP7_75t_L g188 ( 
.A1(n_154),
.A2(n_166),
.B1(n_175),
.B2(n_125),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_L g156 ( 
.A(n_138),
.B(n_107),
.Y(n_156)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_156),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_L g157 ( 
.A(n_138),
.B(n_98),
.Y(n_157)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_157),
.Y(n_194)
);

BUFx5_ASAP7_75t_L g158 ( 
.A(n_130),
.Y(n_158)
);

INVx2_ASAP7_75t_L g189 ( 
.A(n_158),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_L g160 ( 
.A(n_132),
.B(n_97),
.Y(n_160)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_160),
.Y(n_199)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_143),
.Y(n_162)
);

INVx2_ASAP7_75t_SL g163 ( 
.A(n_130),
.Y(n_163)
);

NOR2xp33_ASAP7_75t_L g197 ( 
.A(n_163),
.B(n_172),
.Y(n_197)
);

CKINVDCx20_ASAP7_75t_R g164 ( 
.A(n_143),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_SL g200 ( 
.A(n_164),
.B(n_169),
.Y(n_200)
);

AOI22xp5_ASAP7_75t_L g166 ( 
.A1(n_131),
.A2(n_80),
.B1(n_76),
.B2(n_65),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_L g167 ( 
.A(n_132),
.B(n_97),
.Y(n_167)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_167),
.Y(n_201)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_139),
.Y(n_169)
);

CKINVDCx20_ASAP7_75t_R g172 ( 
.A(n_139),
.Y(n_172)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_127),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_L g178 ( 
.A(n_173),
.B(n_122),
.Y(n_178)
);

INVxp67_ASAP7_75t_L g174 ( 
.A(n_141),
.Y(n_174)
);

INVx1_ASAP7_75t_SL g177 ( 
.A(n_174),
.Y(n_177)
);

AOI22xp5_ASAP7_75t_L g175 ( 
.A1(n_140),
.A2(n_111),
.B1(n_114),
.B2(n_85),
.Y(n_175)
);

NOR2xp33_ASAP7_75t_L g176 ( 
.A(n_126),
.B(n_114),
.Y(n_176)
);

CKINVDCx20_ASAP7_75t_R g187 ( 
.A(n_176),
.Y(n_187)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_178),
.Y(n_203)
);

XOR2xp5_ASAP7_75t_L g179 ( 
.A(n_153),
.B(n_137),
.Y(n_179)
);

MAJIxp5_ASAP7_75t_L g202 ( 
.A(n_179),
.B(n_193),
.C(n_198),
.Y(n_202)
);

NAND2xp5_ASAP7_75t_L g180 ( 
.A(n_152),
.B(n_144),
.Y(n_180)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_180),
.Y(n_205)
);

NAND2xp5_ASAP7_75t_L g183 ( 
.A(n_156),
.B(n_144),
.Y(n_183)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_183),
.Y(n_216)
);

CKINVDCx14_ASAP7_75t_R g209 ( 
.A(n_184),
.Y(n_209)
);

OR2x2_ASAP7_75t_L g185 ( 
.A(n_164),
.B(n_135),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_L g206 ( 
.A(n_185),
.B(n_170),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_L g186 ( 
.A(n_157),
.B(n_124),
.Y(n_186)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_186),
.Y(n_219)
);

OAI22xp5_ASAP7_75t_SL g211 ( 
.A1(n_188),
.A2(n_191),
.B1(n_175),
.B2(n_154),
.Y(n_211)
);

NAND2xp5_ASAP7_75t_L g190 ( 
.A(n_172),
.B(n_136),
.Y(n_190)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_190),
.Y(n_221)
);

AOI22xp5_ASAP7_75t_L g191 ( 
.A1(n_165),
.A2(n_147),
.B1(n_62),
.B2(n_92),
.Y(n_191)
);

MAJIxp5_ASAP7_75t_L g193 ( 
.A(n_153),
.B(n_147),
.C(n_92),
.Y(n_193)
);

CKINVDCx20_ASAP7_75t_R g195 ( 
.A(n_155),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_L g204 ( 
.A(n_195),
.B(n_167),
.Y(n_204)
);

AOI21xp5_ASAP7_75t_L g196 ( 
.A1(n_171),
.A2(n_147),
.B(n_23),
.Y(n_196)
);

NOR2xp33_ASAP7_75t_L g213 ( 
.A(n_196),
.B(n_166),
.Y(n_213)
);

MAJIxp5_ASAP7_75t_L g198 ( 
.A(n_151),
.B(n_147),
.C(n_25),
.Y(n_198)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_204),
.Y(n_231)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_206),
.Y(n_237)
);

NAND2xp5_ASAP7_75t_SL g207 ( 
.A(n_178),
.B(n_150),
.Y(n_207)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_207),
.Y(n_239)
);

AOI22xp5_ASAP7_75t_L g208 ( 
.A1(n_199),
.A2(n_165),
.B1(n_171),
.B2(n_170),
.Y(n_208)
);

OAI22xp5_ASAP7_75t_SL g226 ( 
.A1(n_208),
.A2(n_212),
.B1(n_213),
.B2(n_195),
.Y(n_226)
);

MAJIxp5_ASAP7_75t_L g210 ( 
.A(n_179),
.B(n_177),
.C(n_193),
.Y(n_210)
);

MAJIxp5_ASAP7_75t_L g227 ( 
.A(n_210),
.B(n_214),
.C(n_215),
.Y(n_227)
);

AOI22xp5_ASAP7_75t_L g229 ( 
.A1(n_211),
.A2(n_217),
.B1(n_222),
.B2(n_219),
.Y(n_229)
);

AOI22xp5_ASAP7_75t_L g212 ( 
.A1(n_199),
.A2(n_168),
.B1(n_169),
.B2(n_162),
.Y(n_212)
);

MAJIxp5_ASAP7_75t_L g214 ( 
.A(n_177),
.B(n_149),
.C(n_159),
.Y(n_214)
);

XNOR2xp5_ASAP7_75t_L g215 ( 
.A(n_184),
.B(n_160),
.Y(n_215)
);

OAI22xp5_ASAP7_75t_SL g217 ( 
.A1(n_188),
.A2(n_161),
.B1(n_155),
.B2(n_173),
.Y(n_217)
);

NAND2xp5_ASAP7_75t_L g218 ( 
.A(n_182),
.B(n_148),
.Y(n_218)
);

NAND2xp5_ASAP7_75t_SL g241 ( 
.A(n_218),
.B(n_223),
.Y(n_241)
);

XNOR2xp5_ASAP7_75t_L g220 ( 
.A(n_192),
.B(n_158),
.Y(n_220)
);

MAJIxp5_ASAP7_75t_L g235 ( 
.A(n_220),
.B(n_198),
.C(n_190),
.Y(n_235)
);

OAI22xp5_ASAP7_75t_SL g222 ( 
.A1(n_191),
.A2(n_148),
.B1(n_163),
.B2(n_17),
.Y(n_222)
);

NAND2xp5_ASAP7_75t_L g223 ( 
.A(n_181),
.B(n_163),
.Y(n_223)
);

CKINVDCx20_ASAP7_75t_R g224 ( 
.A(n_197),
.Y(n_224)
);

INVxp67_ASAP7_75t_L g225 ( 
.A(n_224),
.Y(n_225)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_226),
.Y(n_256)
);

XNOR2xp5_ASAP7_75t_L g228 ( 
.A(n_202),
.B(n_210),
.Y(n_228)
);

MAJIxp5_ASAP7_75t_L g246 ( 
.A(n_228),
.B(n_235),
.C(n_236),
.Y(n_246)
);

NAND2xp5_ASAP7_75t_SL g244 ( 
.A(n_229),
.B(n_230),
.Y(n_244)
);

AOI22xp5_ASAP7_75t_L g230 ( 
.A1(n_211),
.A2(n_192),
.B1(n_201),
.B2(n_194),
.Y(n_230)
);

XOR2xp5_ASAP7_75t_L g232 ( 
.A(n_202),
.B(n_186),
.Y(n_232)
);

XOR2xp5_ASAP7_75t_L g249 ( 
.A(n_232),
.B(n_233),
.Y(n_249)
);

XOR2xp5_ASAP7_75t_L g233 ( 
.A(n_215),
.B(n_183),
.Y(n_233)
);

AOI22xp5_ASAP7_75t_L g234 ( 
.A1(n_217),
.A2(n_201),
.B1(n_194),
.B2(n_181),
.Y(n_234)
);

NAND2xp5_ASAP7_75t_L g253 ( 
.A(n_234),
.B(n_242),
.Y(n_253)
);

XNOR2xp5_ASAP7_75t_L g236 ( 
.A(n_214),
.B(n_200),
.Y(n_236)
);

XOR2xp5_ASAP7_75t_L g238 ( 
.A(n_220),
.B(n_180),
.Y(n_238)
);

XOR2xp5_ASAP7_75t_L g255 ( 
.A(n_238),
.B(n_30),
.Y(n_255)
);

OAI321xp33_ASAP7_75t_L g240 ( 
.A1(n_212),
.A2(n_196),
.A3(n_206),
.B1(n_205),
.B2(n_185),
.C(n_208),
.Y(n_240)
);

AOI21xp5_ASAP7_75t_L g250 ( 
.A1(n_240),
.A2(n_237),
.B(n_231),
.Y(n_250)
);

OAI22xp5_ASAP7_75t_SL g242 ( 
.A1(n_209),
.A2(n_221),
.B1(n_203),
.B2(n_223),
.Y(n_242)
);

BUFx2_ASAP7_75t_L g243 ( 
.A(n_222),
.Y(n_243)
);

INVxp33_ASAP7_75t_L g245 ( 
.A(n_243),
.Y(n_245)
);

XNOR2xp5_ASAP7_75t_L g247 ( 
.A(n_228),
.B(n_187),
.Y(n_247)
);

XNOR2xp5_ASAP7_75t_L g268 ( 
.A(n_247),
.B(n_254),
.Y(n_268)
);

MAJIxp5_ASAP7_75t_L g248 ( 
.A(n_232),
.B(n_216),
.C(n_187),
.Y(n_248)
);

MAJIxp5_ASAP7_75t_L g258 ( 
.A(n_248),
.B(n_251),
.C(n_252),
.Y(n_258)
);

OAI321xp33_ASAP7_75t_L g261 ( 
.A1(n_250),
.A2(n_245),
.A3(n_239),
.B1(n_243),
.B2(n_241),
.C(n_225),
.Y(n_261)
);

MAJIxp5_ASAP7_75t_L g251 ( 
.A(n_227),
.B(n_185),
.C(n_189),
.Y(n_251)
);

MAJIxp5_ASAP7_75t_L g252 ( 
.A(n_227),
.B(n_189),
.C(n_25),
.Y(n_252)
);

XNOR2xp5_ASAP7_75t_L g254 ( 
.A(n_235),
.B(n_238),
.Y(n_254)
);

XOR2xp5_ASAP7_75t_L g267 ( 
.A(n_255),
.B(n_257),
.Y(n_267)
);

XOR2xp5_ASAP7_75t_L g257 ( 
.A(n_233),
.B(n_30),
.Y(n_257)
);

XNOR2xp5_ASAP7_75t_L g259 ( 
.A(n_251),
.B(n_248),
.Y(n_259)
);

MAJIxp5_ASAP7_75t_L g277 ( 
.A(n_259),
.B(n_265),
.C(n_4),
.Y(n_277)
);

NAND2xp5_ASAP7_75t_L g260 ( 
.A(n_253),
.B(n_225),
.Y(n_260)
);

NAND2xp5_ASAP7_75t_SL g271 ( 
.A(n_260),
.B(n_261),
.Y(n_271)
);

NAND2xp5_ASAP7_75t_SL g262 ( 
.A(n_244),
.B(n_1),
.Y(n_262)
);

NAND2xp5_ASAP7_75t_L g274 ( 
.A(n_262),
.B(n_263),
.Y(n_274)
);

NOR2xp33_ASAP7_75t_SL g263 ( 
.A(n_246),
.B(n_1),
.Y(n_263)
);

NAND2xp5_ASAP7_75t_L g264 ( 
.A(n_256),
.B(n_2),
.Y(n_264)
);

CKINVDCx16_ASAP7_75t_R g275 ( 
.A(n_264),
.Y(n_275)
);

AOI22xp5_ASAP7_75t_L g265 ( 
.A1(n_245),
.A2(n_2),
.B1(n_3),
.B2(n_4),
.Y(n_265)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_255),
.Y(n_266)
);

NOR2xp33_ASAP7_75t_L g270 ( 
.A(n_266),
.B(n_269),
.Y(n_270)
);

NOR2xp33_ASAP7_75t_SL g269 ( 
.A(n_257),
.B(n_3),
.Y(n_269)
);

NOR2xp33_ASAP7_75t_SL g272 ( 
.A(n_259),
.B(n_268),
.Y(n_272)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_272),
.Y(n_280)
);

OAI21xp5_ASAP7_75t_L g273 ( 
.A1(n_258),
.A2(n_249),
.B(n_5),
.Y(n_273)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_273),
.Y(n_283)
);

OAI21xp5_ASAP7_75t_SL g276 ( 
.A1(n_258),
.A2(n_249),
.B(n_5),
.Y(n_276)
);

NAND2xp5_ASAP7_75t_SL g284 ( 
.A(n_276),
.B(n_277),
.Y(n_284)
);

NOR2xp33_ASAP7_75t_SL g278 ( 
.A(n_267),
.B(n_4),
.Y(n_278)
);

NOR2xp33_ASAP7_75t_L g285 ( 
.A(n_278),
.B(n_6),
.Y(n_285)
);

NOR2xp33_ASAP7_75t_SL g279 ( 
.A(n_275),
.B(n_267),
.Y(n_279)
);

NOR2xp33_ASAP7_75t_L g289 ( 
.A(n_279),
.B(n_281),
.Y(n_289)
);

NAND2xp5_ASAP7_75t_L g281 ( 
.A(n_271),
.B(n_5),
.Y(n_281)
);

AOI31xp67_ASAP7_75t_L g282 ( 
.A1(n_271),
.A2(n_6),
.A3(n_7),
.B(n_8),
.Y(n_282)
);

OAI22xp5_ASAP7_75t_L g290 ( 
.A1(n_282),
.A2(n_285),
.B1(n_283),
.B2(n_13),
.Y(n_290)
);

AOI322xp5_ASAP7_75t_L g288 ( 
.A1(n_285),
.A2(n_9),
.A3(n_10),
.B1(n_11),
.B2(n_12),
.C1(n_13),
.C2(n_15),
.Y(n_288)
);

OAI21xp5_ASAP7_75t_L g286 ( 
.A1(n_280),
.A2(n_270),
.B(n_274),
.Y(n_286)
);

CKINVDCx20_ASAP7_75t_R g291 ( 
.A(n_286),
.Y(n_291)
);

OAI21xp5_ASAP7_75t_SL g287 ( 
.A1(n_284),
.A2(n_8),
.B(n_9),
.Y(n_287)
);

NAND2xp5_ASAP7_75t_SL g293 ( 
.A(n_287),
.B(n_290),
.Y(n_293)
);

AO221x1_ASAP7_75t_L g292 ( 
.A1(n_288),
.A2(n_289),
.B1(n_11),
.B2(n_15),
.C(n_10),
.Y(n_292)
);

BUFx24_ASAP7_75t_SL g294 ( 
.A(n_292),
.Y(n_294)
);

MAJIxp5_ASAP7_75t_L g295 ( 
.A(n_291),
.B(n_30),
.C(n_23),
.Y(n_295)
);

NAND2xp5_ASAP7_75t_SL g296 ( 
.A(n_295),
.B(n_293),
.Y(n_296)
);

XNOR2xp5_ASAP7_75t_L g297 ( 
.A(n_296),
.B(n_294),
.Y(n_297)
);


endmodule