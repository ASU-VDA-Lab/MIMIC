module fake_jpeg_15373_n_142 (n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_142);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_142;

wire n_117;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_29;
wire n_103;
wire n_50;
wire n_15;
wire n_124;
wire n_141;
wire n_13;
wire n_57;
wire n_21;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_30;
wire n_106;
wire n_111;
wire n_44;
wire n_24;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_121;
wire n_99;
wire n_102;
wire n_130;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_78;
wire n_18;
wire n_20;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_97;
wire n_135;
wire n_36;
wire n_62;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

BUFx16f_ASAP7_75t_L g13 ( 
.A(n_12),
.Y(n_13)
);

INVx1_ASAP7_75t_L g14 ( 
.A(n_4),
.Y(n_14)
);

CKINVDCx16_ASAP7_75t_R g15 ( 
.A(n_8),
.Y(n_15)
);

BUFx6f_ASAP7_75t_L g16 ( 
.A(n_2),
.Y(n_16)
);

BUFx16f_ASAP7_75t_L g17 ( 
.A(n_12),
.Y(n_17)
);

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_5),
.Y(n_18)
);

HB1xp67_ASAP7_75t_L g19 ( 
.A(n_7),
.Y(n_19)
);

INVx8_ASAP7_75t_SL g20 ( 
.A(n_1),
.Y(n_20)
);

BUFx12_ASAP7_75t_L g21 ( 
.A(n_5),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_9),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_8),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_5),
.Y(n_24)
);

INVx6_ASAP7_75t_L g25 ( 
.A(n_4),
.Y(n_25)
);

INVx6_ASAP7_75t_L g26 ( 
.A(n_1),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_7),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_4),
.Y(n_28)
);

INVx6_ASAP7_75t_SL g29 ( 
.A(n_13),
.Y(n_29)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_29),
.B(n_30),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g30 ( 
.A(n_22),
.B(n_0),
.Y(n_30)
);

BUFx4f_ASAP7_75t_SL g31 ( 
.A(n_13),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_31),
.Y(n_46)
);

INVx6_ASAP7_75t_L g32 ( 
.A(n_13),
.Y(n_32)
);

INVx2_ASAP7_75t_L g45 ( 
.A(n_32),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g33 ( 
.A(n_22),
.B(n_0),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_33),
.B(n_34),
.Y(n_60)
);

BUFx12_ASAP7_75t_L g34 ( 
.A(n_13),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_L g35 ( 
.A(n_27),
.B(n_0),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_35),
.B(n_40),
.Y(n_64)
);

INVx3_ASAP7_75t_L g36 ( 
.A(n_16),
.Y(n_36)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_36),
.Y(n_54)
);

BUFx24_ASAP7_75t_L g37 ( 
.A(n_17),
.Y(n_37)
);

INVxp67_ASAP7_75t_L g59 ( 
.A(n_37),
.Y(n_59)
);

INVx2_ASAP7_75t_L g38 ( 
.A(n_16),
.Y(n_38)
);

INVx2_ASAP7_75t_L g50 ( 
.A(n_38),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_16),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_39),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g40 ( 
.A(n_27),
.B(n_1),
.Y(n_40)
);

INVx8_ASAP7_75t_L g41 ( 
.A(n_25),
.Y(n_41)
);

INVx4_ASAP7_75t_L g55 ( 
.A(n_41),
.Y(n_55)
);

BUFx3_ASAP7_75t_L g42 ( 
.A(n_16),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_42),
.B(n_19),
.Y(n_65)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_18),
.Y(n_43)
);

INVx3_ASAP7_75t_L g47 ( 
.A(n_43),
.Y(n_47)
);

BUFx12f_ASAP7_75t_L g44 ( 
.A(n_18),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g63 ( 
.A(n_44),
.Y(n_63)
);

INVx3_ASAP7_75t_L g48 ( 
.A(n_36),
.Y(n_48)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_48),
.Y(n_81)
);

OAI22xp5_ASAP7_75t_SL g49 ( 
.A1(n_41),
.A2(n_26),
.B1(n_25),
.B2(n_17),
.Y(n_49)
);

OAI22xp5_ASAP7_75t_L g80 ( 
.A1(n_49),
.A2(n_53),
.B1(n_57),
.B2(n_62),
.Y(n_80)
);

AOI21xp5_ASAP7_75t_L g52 ( 
.A1(n_37),
.A2(n_17),
.B(n_3),
.Y(n_52)
);

A2O1A1Ixp33_ASAP7_75t_L g82 ( 
.A1(n_52),
.A2(n_14),
.B(n_28),
.C(n_15),
.Y(n_82)
);

OAI22xp5_ASAP7_75t_SL g53 ( 
.A1(n_38),
.A2(n_26),
.B1(n_25),
.B2(n_17),
.Y(n_53)
);

OAI22xp5_ASAP7_75t_L g57 ( 
.A1(n_32),
.A2(n_26),
.B1(n_28),
.B2(n_24),
.Y(n_57)
);

INVx3_ASAP7_75t_L g58 ( 
.A(n_39),
.Y(n_58)
);

INVx8_ASAP7_75t_L g70 ( 
.A(n_58),
.Y(n_70)
);

CKINVDCx12_ASAP7_75t_R g61 ( 
.A(n_31),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_61),
.B(n_66),
.Y(n_68)
);

OAI22xp33_ASAP7_75t_SL g62 ( 
.A1(n_43),
.A2(n_18),
.B1(n_19),
.B2(n_20),
.Y(n_62)
);

CKINVDCx16_ASAP7_75t_R g77 ( 
.A(n_65),
.Y(n_77)
);

INVx3_ASAP7_75t_L g66 ( 
.A(n_42),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_L g67 ( 
.A(n_52),
.B(n_31),
.Y(n_67)
);

MAJIxp5_ASAP7_75t_L g87 ( 
.A(n_67),
.B(n_73),
.C(n_74),
.Y(n_87)
);

OR2x4_ASAP7_75t_L g69 ( 
.A(n_53),
.B(n_20),
.Y(n_69)
);

AOI21xp5_ASAP7_75t_L g94 ( 
.A1(n_69),
.A2(n_71),
.B(n_82),
.Y(n_94)
);

AOI21xp33_ASAP7_75t_L g71 ( 
.A1(n_64),
.A2(n_23),
.B(n_24),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_SL g72 ( 
.A(n_56),
.B(n_23),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_72),
.B(n_75),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g73 ( 
.A(n_46),
.B(n_54),
.Y(n_73)
);

MAJIxp5_ASAP7_75t_L g74 ( 
.A(n_63),
.B(n_37),
.C(n_44),
.Y(n_74)
);

INVx1_ASAP7_75t_SL g75 ( 
.A(n_51),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_L g76 ( 
.A(n_54),
.B(n_44),
.Y(n_76)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_76),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_60),
.B(n_21),
.Y(n_78)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_78),
.Y(n_95)
);

AOI32xp33_ASAP7_75t_L g79 ( 
.A1(n_59),
.A2(n_49),
.A3(n_55),
.B1(n_29),
.B2(n_34),
.Y(n_79)
);

AOI22xp5_ASAP7_75t_L g86 ( 
.A1(n_79),
.A2(n_59),
.B1(n_55),
.B2(n_58),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_L g83 ( 
.A(n_50),
.B(n_44),
.Y(n_83)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_83),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_SL g84 ( 
.A(n_45),
.B(n_14),
.Y(n_84)
);

OAI22xp5_ASAP7_75t_L g89 ( 
.A1(n_84),
.A2(n_85),
.B1(n_81),
.B2(n_15),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_45),
.B(n_21),
.Y(n_85)
);

XNOR2xp5_ASAP7_75t_SL g104 ( 
.A(n_86),
.B(n_79),
.Y(n_104)
);

OAI22xp5_ASAP7_75t_SL g88 ( 
.A1(n_67),
.A2(n_50),
.B1(n_48),
.B2(n_47),
.Y(n_88)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_88),
.Y(n_102)
);

CKINVDCx16_ASAP7_75t_R g109 ( 
.A(n_89),
.Y(n_109)
);

INVx3_ASAP7_75t_L g91 ( 
.A(n_70),
.Y(n_91)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_91),
.Y(n_112)
);

OAI22xp5_ASAP7_75t_SL g92 ( 
.A1(n_69),
.A2(n_47),
.B1(n_66),
.B2(n_51),
.Y(n_92)
);

INVxp67_ASAP7_75t_L g105 ( 
.A(n_92),
.Y(n_105)
);

OAI22xp5_ASAP7_75t_SL g93 ( 
.A1(n_80),
.A2(n_18),
.B1(n_21),
.B2(n_34),
.Y(n_93)
);

XOR2xp5_ASAP7_75t_L g107 ( 
.A(n_93),
.B(n_74),
.Y(n_107)
);

OAI22xp5_ASAP7_75t_L g96 ( 
.A1(n_77),
.A2(n_21),
.B1(n_3),
.B2(n_6),
.Y(n_96)
);

CKINVDCx20_ASAP7_75t_R g111 ( 
.A(n_96),
.Y(n_111)
);

INVx1_ASAP7_75t_SL g98 ( 
.A(n_75),
.Y(n_98)
);

AO221x1_ASAP7_75t_L g110 ( 
.A1(n_98),
.A2(n_70),
.B1(n_81),
.B2(n_21),
.C(n_82),
.Y(n_110)
);

INVx13_ASAP7_75t_L g100 ( 
.A(n_68),
.Y(n_100)
);

INVx13_ASAP7_75t_L g103 ( 
.A(n_100),
.Y(n_103)
);

OAI21xp5_ASAP7_75t_L g101 ( 
.A1(n_94),
.A2(n_73),
.B(n_84),
.Y(n_101)
);

AO21x1_ASAP7_75t_L g118 ( 
.A1(n_101),
.A2(n_95),
.B(n_99),
.Y(n_118)
);

XNOR2xp5_ASAP7_75t_SL g119 ( 
.A(n_104),
.B(n_92),
.Y(n_119)
);

BUFx12f_ASAP7_75t_SL g106 ( 
.A(n_94),
.Y(n_106)
);

NAND2xp33_ASAP7_75t_SL g114 ( 
.A(n_106),
.B(n_86),
.Y(n_114)
);

AOI22xp5_ASAP7_75t_L g116 ( 
.A1(n_107),
.A2(n_87),
.B1(n_97),
.B2(n_90),
.Y(n_116)
);

MAJIxp5_ASAP7_75t_L g108 ( 
.A(n_87),
.B(n_83),
.C(n_76),
.Y(n_108)
);

MAJIxp5_ASAP7_75t_L g120 ( 
.A(n_108),
.B(n_88),
.C(n_95),
.Y(n_120)
);

AO221x1_ASAP7_75t_L g121 ( 
.A1(n_110),
.A2(n_98),
.B1(n_91),
.B2(n_93),
.C(n_100),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_L g113 ( 
.A(n_108),
.B(n_90),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_L g126 ( 
.A(n_113),
.B(n_115),
.Y(n_126)
);

OAI21xp5_ASAP7_75t_L g122 ( 
.A1(n_114),
.A2(n_117),
.B(n_118),
.Y(n_122)
);

CKINVDCx20_ASAP7_75t_R g115 ( 
.A(n_112),
.Y(n_115)
);

MAJIxp5_ASAP7_75t_L g124 ( 
.A(n_116),
.B(n_119),
.C(n_120),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_L g117 ( 
.A(n_101),
.B(n_97),
.Y(n_117)
);

OAI21xp5_ASAP7_75t_L g123 ( 
.A1(n_121),
.A2(n_110),
.B(n_105),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_SL g133 ( 
.A(n_123),
.B(n_112),
.Y(n_133)
);

AND2x2_ASAP7_75t_L g125 ( 
.A(n_120),
.B(n_106),
.Y(n_125)
);

OAI21xp5_ASAP7_75t_SL g132 ( 
.A1(n_125),
.A2(n_127),
.B(n_128),
.Y(n_132)
);

A2O1A1O1Ixp25_ASAP7_75t_L g127 ( 
.A1(n_119),
.A2(n_104),
.B(n_107),
.C(n_109),
.D(n_105),
.Y(n_127)
);

AOI21xp5_ASAP7_75t_L g128 ( 
.A1(n_117),
.A2(n_102),
.B(n_109),
.Y(n_128)
);

INVxp67_ASAP7_75t_L g129 ( 
.A(n_126),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_L g135 ( 
.A(n_129),
.B(n_130),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_L g130 ( 
.A(n_122),
.B(n_118),
.Y(n_130)
);

OAI21xp33_ASAP7_75t_L g131 ( 
.A1(n_124),
.A2(n_113),
.B(n_102),
.Y(n_131)
);

OAI211xp5_ASAP7_75t_L g136 ( 
.A1(n_131),
.A2(n_133),
.B(n_111),
.C(n_103),
.Y(n_136)
);

MAJIxp5_ASAP7_75t_L g134 ( 
.A(n_132),
.B(n_116),
.C(n_111),
.Y(n_134)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_134),
.Y(n_138)
);

NOR2x1_ASAP7_75t_L g137 ( 
.A(n_136),
.B(n_103),
.Y(n_137)
);

A2O1A1Ixp33_ASAP7_75t_L g139 ( 
.A1(n_137),
.A2(n_135),
.B(n_3),
.C(n_6),
.Y(n_139)
);

MAJIxp5_ASAP7_75t_L g141 ( 
.A(n_139),
.B(n_140),
.C(n_138),
.Y(n_141)
);

MAJx2_ASAP7_75t_L g140 ( 
.A(n_137),
.B(n_9),
.C(n_10),
.Y(n_140)
);

AOI322xp5_ASAP7_75t_L g142 ( 
.A1(n_141),
.A2(n_2),
.A3(n_6),
.B1(n_10),
.B2(n_11),
.C1(n_103),
.C2(n_137),
.Y(n_142)
);


endmodule