module real_jpeg_4896_n_15 (n_108, n_8, n_0, n_2, n_10, n_9, n_12, n_107, n_6, n_104, n_100, n_106, n_11, n_14, n_7, n_3, n_99, n_5, n_4, n_102, n_105, n_101, n_1, n_13, n_103, n_15);

input n_108;
input n_8;
input n_0;
input n_2;
input n_10;
input n_9;
input n_12;
input n_107;
input n_6;
input n_104;
input n_100;
input n_106;
input n_11;
input n_14;
input n_7;
input n_3;
input n_99;
input n_5;
input n_4;
input n_102;
input n_105;
input n_101;
input n_1;
input n_13;
input n_103;

output n_15;

wire n_54;
wire n_37;
wire n_73;
wire n_35;
wire n_38;
wire n_29;
wire n_91;
wire n_49;
wire n_68;
wire n_83;
wire n_78;
wire n_64;
wire n_47;
wire n_22;
wire n_87;
wire n_40;
wire n_27;
wire n_56;
wire n_48;
wire n_93;
wire n_95;
wire n_65;
wire n_33;
wire n_76;
wire n_67;
wire n_79;
wire n_66;
wire n_28;
wire n_44;
wire n_62;
wire n_45;
wire n_42;
wire n_18;
wire n_77;
wire n_39;
wire n_94;
wire n_26;
wire n_19;
wire n_17;
wire n_21;
wire n_50;
wire n_69;
wire n_31;
wire n_72;
wire n_23;
wire n_51;
wire n_71;
wire n_90;
wire n_61;
wire n_86;
wire n_70;
wire n_41;
wire n_74;
wire n_80;
wire n_32;
wire n_20;
wire n_30;
wire n_43;
wire n_57;
wire n_84;
wire n_82;
wire n_55;
wire n_58;
wire n_52;
wire n_63;
wire n_24;
wire n_92;
wire n_75;
wire n_97;
wire n_34;
wire n_60;
wire n_46;
wire n_88;
wire n_59;
wire n_25;
wire n_53;
wire n_36;
wire n_81;
wire n_85;
wire n_96;
wire n_89;
wire n_16;

INVx5_ASAP7_75t_L g24 ( 
.A(n_0),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_0),
.Y(n_40)
);

BUFx5_ASAP7_75t_L g58 ( 
.A(n_0),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_SL g71 ( 
.A(n_0),
.B(n_72),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g35 ( 
.A(n_1),
.B(n_36),
.Y(n_35)
);

NAND2xp5_ASAP7_75t_L g94 ( 
.A(n_1),
.B(n_36),
.Y(n_94)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_2),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_3),
.B(n_71),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_L g73 ( 
.A(n_3),
.B(n_71),
.Y(n_73)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_4),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_5),
.Y(n_30)
);

NOR2xp33_ASAP7_75t_L g18 ( 
.A(n_6),
.B(n_19),
.Y(n_18)
);

AND2x2_ASAP7_75t_L g26 ( 
.A(n_6),
.B(n_19),
.Y(n_26)
);

NOR2xp33_ASAP7_75t_SL g28 ( 
.A(n_7),
.B(n_29),
.Y(n_28)
);

AND2x2_ASAP7_75t_L g97 ( 
.A(n_7),
.B(n_29),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_SL g46 ( 
.A(n_8),
.B(n_47),
.Y(n_46)
);

AND2x2_ASAP7_75t_L g76 ( 
.A(n_8),
.B(n_47),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_SL g51 ( 
.A(n_9),
.B(n_52),
.Y(n_51)
);

AND2x2_ASAP7_75t_L g77 ( 
.A(n_9),
.B(n_52),
.Y(n_77)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_10),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_11),
.B(n_84),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g88 ( 
.A(n_11),
.B(n_84),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_SL g90 ( 
.A(n_12),
.B(n_91),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_L g95 ( 
.A(n_12),
.B(n_91),
.Y(n_95)
);

AND2x2_ASAP7_75t_L g62 ( 
.A(n_13),
.B(n_63),
.Y(n_62)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_14),
.Y(n_68)
);

XOR2xp5_ASAP7_75t_L g15 ( 
.A(n_16),
.B(n_27),
.Y(n_15)
);

NAND2xp5_ASAP7_75t_SL g16 ( 
.A(n_17),
.B(n_25),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_18),
.Y(n_17)
);

NOR2xp33_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_21),
.Y(n_19)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_21),
.B(n_92),
.Y(n_91)
);

INVx8_ASAP7_75t_L g21 ( 
.A(n_22),
.Y(n_21)
);

INVx6_ASAP7_75t_L g22 ( 
.A(n_23),
.Y(n_22)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_23),
.B(n_64),
.Y(n_63)
);

INVx4_ASAP7_75t_L g23 ( 
.A(n_24),
.Y(n_23)
);

BUFx3_ASAP7_75t_L g32 ( 
.A(n_24),
.Y(n_32)
);

INVx5_ASAP7_75t_L g50 ( 
.A(n_24),
.Y(n_50)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_26),
.Y(n_25)
);

OAI21xp5_ASAP7_75t_L g27 ( 
.A1(n_28),
.A2(n_33),
.B(n_96),
.Y(n_27)
);

NOR2xp33_ASAP7_75t_L g29 ( 
.A(n_30),
.B(n_31),
.Y(n_29)
);

INVx3_ASAP7_75t_L g31 ( 
.A(n_32),
.Y(n_31)
);

AOI21xp5_ASAP7_75t_L g33 ( 
.A1(n_34),
.A2(n_89),
.B(n_93),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_L g34 ( 
.A(n_35),
.B(n_41),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_L g36 ( 
.A(n_37),
.B(n_38),
.Y(n_36)
);

BUFx8_ASAP7_75t_L g38 ( 
.A(n_39),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_39),
.B(n_53),
.Y(n_52)
);

BUFx12f_ASAP7_75t_L g39 ( 
.A(n_40),
.Y(n_39)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_42),
.Y(n_41)
);

OAI21x1_ASAP7_75t_L g42 ( 
.A1(n_43),
.A2(n_83),
.B(n_88),
.Y(n_42)
);

AOI21xp5_ASAP7_75t_L g43 ( 
.A1(n_44),
.A2(n_78),
.B(n_82),
.Y(n_43)
);

AO221x1_ASAP7_75t_L g44 ( 
.A1(n_45),
.A2(n_54),
.B1(n_75),
.B2(n_76),
.C(n_77),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g45 ( 
.A(n_46),
.B(n_51),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g47 ( 
.A(n_48),
.B(n_49),
.Y(n_47)
);

OR2x2_ASAP7_75t_L g79 ( 
.A(n_49),
.B(n_80),
.Y(n_79)
);

BUFx12_ASAP7_75t_L g49 ( 
.A(n_50),
.Y(n_49)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_51),
.Y(n_75)
);

AO21x1_ASAP7_75t_L g54 ( 
.A1(n_55),
.A2(n_60),
.B(n_74),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_SL g55 ( 
.A(n_56),
.B(n_59),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_56),
.B(n_59),
.Y(n_74)
);

OR2x2_ASAP7_75t_L g56 ( 
.A(n_57),
.B(n_58),
.Y(n_56)
);

OR2x2_ASAP7_75t_L g66 ( 
.A(n_58),
.B(n_67),
.Y(n_66)
);

INVx2_ASAP7_75t_L g87 ( 
.A(n_58),
.Y(n_87)
);

OAI21xp5_ASAP7_75t_L g60 ( 
.A1(n_61),
.A2(n_70),
.B(n_73),
.Y(n_60)
);

AOI21xp5_ASAP7_75t_L g61 ( 
.A1(n_62),
.A2(n_65),
.B(n_69),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_SL g65 ( 
.A(n_66),
.B(n_68),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_66),
.B(n_68),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_SL g78 ( 
.A(n_79),
.B(n_81),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_79),
.B(n_81),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_85),
.B(n_86),
.Y(n_84)
);

INVx4_ASAP7_75t_L g86 ( 
.A(n_87),
.Y(n_86)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_90),
.Y(n_89)
);

OAI21xp5_ASAP7_75t_L g93 ( 
.A1(n_90),
.A2(n_94),
.B(n_95),
.Y(n_93)
);

CKINVDCx20_ASAP7_75t_R g96 ( 
.A(n_97),
.Y(n_96)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_99),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_100),
.Y(n_48)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_101),
.Y(n_53)
);

CKINVDCx20_ASAP7_75t_R g57 ( 
.A(n_102),
.Y(n_57)
);

CKINVDCx20_ASAP7_75t_R g64 ( 
.A(n_103),
.Y(n_64)
);

CKINVDCx20_ASAP7_75t_R g67 ( 
.A(n_104),
.Y(n_67)
);

CKINVDCx20_ASAP7_75t_R g72 ( 
.A(n_105),
.Y(n_72)
);

CKINVDCx20_ASAP7_75t_R g80 ( 
.A(n_106),
.Y(n_80)
);

CKINVDCx20_ASAP7_75t_R g85 ( 
.A(n_107),
.Y(n_85)
);

CKINVDCx20_ASAP7_75t_R g92 ( 
.A(n_108),
.Y(n_92)
);


endmodule