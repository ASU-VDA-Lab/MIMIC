module fake_jpeg_20726_n_151 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_151);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_151;

wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_147;
wire n_73;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_15;
wire n_124;
wire n_141;
wire n_21;
wire n_57;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_106;
wire n_111;
wire n_24;
wire n_44;
wire n_143;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_78;
wire n_18;
wire n_20;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_33;
wire n_91;
wire n_93;
wire n_54;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_149;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_97;
wire n_135;
wire n_36;
wire n_62;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

INVx4_ASAP7_75t_L g15 ( 
.A(n_9),
.Y(n_15)
);

NOR2xp33_ASAP7_75t_L g16 ( 
.A(n_8),
.B(n_0),
.Y(n_16)
);

BUFx6f_ASAP7_75t_L g17 ( 
.A(n_14),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_0),
.Y(n_18)
);

BUFx3_ASAP7_75t_L g19 ( 
.A(n_6),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_11),
.Y(n_20)
);

INVx2_ASAP7_75t_L g21 ( 
.A(n_13),
.Y(n_21)
);

INVx11_ASAP7_75t_SL g22 ( 
.A(n_13),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_12),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_12),
.Y(n_24)
);

CKINVDCx16_ASAP7_75t_R g25 ( 
.A(n_4),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_1),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_7),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_1),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_10),
.Y(n_29)
);

NOR2xp33_ASAP7_75t_L g30 ( 
.A(n_9),
.B(n_6),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_2),
.Y(n_31)
);

AOI21xp33_ASAP7_75t_L g32 ( 
.A1(n_16),
.A2(n_0),
.B(n_1),
.Y(n_32)
);

NOR2xp33_ASAP7_75t_L g51 ( 
.A(n_32),
.B(n_34),
.Y(n_51)
);

INVx4_ASAP7_75t_L g33 ( 
.A(n_19),
.Y(n_33)
);

INVx3_ASAP7_75t_L g52 ( 
.A(n_33),
.Y(n_52)
);

INVx5_ASAP7_75t_L g34 ( 
.A(n_31),
.Y(n_34)
);

BUFx12f_ASAP7_75t_L g35 ( 
.A(n_31),
.Y(n_35)
);

INVx11_ASAP7_75t_L g54 ( 
.A(n_35),
.Y(n_54)
);

BUFx5_ASAP7_75t_L g36 ( 
.A(n_31),
.Y(n_36)
);

INVx13_ASAP7_75t_L g47 ( 
.A(n_36),
.Y(n_47)
);

INVx11_ASAP7_75t_L g37 ( 
.A(n_22),
.Y(n_37)
);

AO22x1_ASAP7_75t_L g46 ( 
.A1(n_37),
.A2(n_38),
.B1(n_25),
.B2(n_19),
.Y(n_46)
);

INVx2_ASAP7_75t_SL g38 ( 
.A(n_17),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_L g39 ( 
.A(n_16),
.B(n_2),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_39),
.B(n_41),
.Y(n_60)
);

INVx8_ASAP7_75t_L g40 ( 
.A(n_17),
.Y(n_40)
);

INVx3_ASAP7_75t_L g59 ( 
.A(n_40),
.Y(n_59)
);

BUFx12f_ASAP7_75t_L g41 ( 
.A(n_17),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g42 ( 
.A(n_30),
.B(n_2),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_42),
.B(n_43),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g43 ( 
.A(n_30),
.B(n_3),
.Y(n_43)
);

NAND3xp33_ASAP7_75t_SL g44 ( 
.A(n_39),
.B(n_29),
.C(n_24),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_44),
.B(n_55),
.Y(n_69)
);

AOI22xp33_ASAP7_75t_L g45 ( 
.A1(n_38),
.A2(n_40),
.B1(n_21),
.B2(n_34),
.Y(n_45)
);

AOI22xp33_ASAP7_75t_L g68 ( 
.A1(n_45),
.A2(n_53),
.B1(n_59),
.B2(n_48),
.Y(n_68)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_46),
.Y(n_71)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_33),
.Y(n_48)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_48),
.Y(n_77)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_33),
.Y(n_49)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_49),
.Y(n_80)
);

AOI21xp33_ASAP7_75t_L g50 ( 
.A1(n_42),
.A2(n_27),
.B(n_26),
.Y(n_50)
);

AOI21xp5_ASAP7_75t_L g79 ( 
.A1(n_50),
.A2(n_56),
.B(n_23),
.Y(n_79)
);

OAI22xp5_ASAP7_75t_SL g53 ( 
.A1(n_40),
.A2(n_21),
.B1(n_15),
.B2(n_18),
.Y(n_53)
);

OAI22xp5_ASAP7_75t_SL g83 ( 
.A1(n_53),
.A2(n_57),
.B1(n_58),
.B2(n_37),
.Y(n_83)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_36),
.Y(n_55)
);

O2A1O1Ixp33_ASAP7_75t_SL g56 ( 
.A1(n_38),
.A2(n_25),
.B(n_28),
.C(n_18),
.Y(n_56)
);

OAI22xp33_ASAP7_75t_SL g57 ( 
.A1(n_38),
.A2(n_34),
.B1(n_15),
.B2(n_28),
.Y(n_57)
);

OAI22xp5_ASAP7_75t_SL g58 ( 
.A1(n_43),
.A2(n_27),
.B1(n_26),
.B2(n_29),
.Y(n_58)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_35),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_61),
.B(n_47),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_L g63 ( 
.A(n_35),
.B(n_3),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_L g65 ( 
.A(n_63),
.B(n_35),
.Y(n_65)
);

AOI21xp5_ASAP7_75t_L g64 ( 
.A1(n_41),
.A2(n_3),
.B(n_4),
.Y(n_64)
);

OAI21xp5_ASAP7_75t_L g74 ( 
.A1(n_64),
.A2(n_23),
.B(n_20),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_SL g89 ( 
.A(n_65),
.B(n_67),
.Y(n_89)
);

AOI22xp33_ASAP7_75t_SL g66 ( 
.A1(n_52),
.A2(n_37),
.B1(n_20),
.B2(n_24),
.Y(n_66)
);

AOI22xp5_ASAP7_75t_SL g95 ( 
.A1(n_66),
.A2(n_68),
.B1(n_74),
.B2(n_83),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g67 ( 
.A(n_63),
.B(n_35),
.Y(n_67)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_52),
.Y(n_70)
);

BUFx6f_ASAP7_75t_L g98 ( 
.A(n_70),
.Y(n_98)
);

AND2x2_ASAP7_75t_L g97 ( 
.A(n_72),
.B(n_84),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g73 ( 
.A(n_58),
.B(n_41),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_SL g93 ( 
.A(n_73),
.B(n_75),
.Y(n_93)
);

CKINVDCx16_ASAP7_75t_R g75 ( 
.A(n_49),
.Y(n_75)
);

INVxp67_ASAP7_75t_L g76 ( 
.A(n_60),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_SL g103 ( 
.A(n_76),
.B(n_78),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_L g78 ( 
.A(n_64),
.B(n_41),
.Y(n_78)
);

OAI22xp5_ASAP7_75t_SL g100 ( 
.A1(n_79),
.A2(n_87),
.B1(n_56),
.B2(n_61),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_L g81 ( 
.A(n_60),
.B(n_41),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_81),
.B(n_82),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_62),
.B(n_4),
.Y(n_82)
);

AND2x2_ASAP7_75t_L g84 ( 
.A(n_51),
.B(n_5),
.Y(n_84)
);

NAND3xp33_ASAP7_75t_SL g85 ( 
.A(n_51),
.B(n_8),
.C(n_10),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_85),
.B(n_86),
.Y(n_94)
);

AND2x2_ASAP7_75t_L g86 ( 
.A(n_62),
.B(n_5),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_L g87 ( 
.A(n_50),
.B(n_5),
.Y(n_87)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_77),
.Y(n_88)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_88),
.Y(n_106)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_77),
.Y(n_91)
);

CKINVDCx16_ASAP7_75t_R g109 ( 
.A(n_91),
.Y(n_109)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_80),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_L g104 ( 
.A(n_92),
.B(n_96),
.Y(n_104)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_72),
.Y(n_96)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_71),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g113 ( 
.A(n_99),
.B(n_100),
.Y(n_113)
);

OAI22xp5_ASAP7_75t_SL g101 ( 
.A1(n_79),
.A2(n_56),
.B1(n_59),
.B2(n_55),
.Y(n_101)
);

OAI22xp5_ASAP7_75t_SL g115 ( 
.A1(n_101),
.A2(n_84),
.B1(n_82),
.B2(n_70),
.Y(n_115)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_71),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_L g116 ( 
.A(n_102),
.B(n_46),
.Y(n_116)
);

INVxp67_ASAP7_75t_L g105 ( 
.A(n_103),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_L g128 ( 
.A(n_105),
.B(n_116),
.Y(n_128)
);

MAJIxp5_ASAP7_75t_L g107 ( 
.A(n_89),
.B(n_78),
.C(n_87),
.Y(n_107)
);

MAJIxp5_ASAP7_75t_L g121 ( 
.A(n_107),
.B(n_110),
.C(n_111),
.Y(n_121)
);

AOI21xp5_ASAP7_75t_L g108 ( 
.A1(n_101),
.A2(n_74),
.B(n_73),
.Y(n_108)
);

INVxp67_ASAP7_75t_L g129 ( 
.A(n_108),
.Y(n_129)
);

XOR2xp5_ASAP7_75t_L g110 ( 
.A(n_100),
.B(n_67),
.Y(n_110)
);

MAJIxp5_ASAP7_75t_L g111 ( 
.A(n_96),
.B(n_65),
.C(n_81),
.Y(n_111)
);

OAI22xp5_ASAP7_75t_L g112 ( 
.A1(n_99),
.A2(n_83),
.B1(n_69),
.B2(n_75),
.Y(n_112)
);

AOI22xp5_ASAP7_75t_L g119 ( 
.A1(n_112),
.A2(n_95),
.B1(n_97),
.B2(n_88),
.Y(n_119)
);

BUFx12f_ASAP7_75t_L g114 ( 
.A(n_98),
.Y(n_114)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_114),
.Y(n_122)
);

AOI22xp5_ASAP7_75t_L g120 ( 
.A1(n_115),
.A2(n_97),
.B1(n_90),
.B2(n_95),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_L g117 ( 
.A(n_93),
.B(n_84),
.Y(n_117)
);

OAI211xp5_ASAP7_75t_SL g127 ( 
.A1(n_117),
.A2(n_105),
.B(n_108),
.C(n_118),
.Y(n_127)
);

AOI21xp5_ASAP7_75t_L g118 ( 
.A1(n_102),
.A2(n_86),
.B(n_47),
.Y(n_118)
);

AOI21xp5_ASAP7_75t_L g125 ( 
.A1(n_118),
.A2(n_46),
.B(n_47),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_L g133 ( 
.A(n_119),
.B(n_120),
.Y(n_133)
);

MAJIxp5_ASAP7_75t_L g123 ( 
.A(n_110),
.B(n_97),
.C(n_92),
.Y(n_123)
);

XNOR2xp5_ASAP7_75t_L g132 ( 
.A(n_123),
.B(n_125),
.Y(n_132)
);

AOI22xp5_ASAP7_75t_L g124 ( 
.A1(n_112),
.A2(n_91),
.B1(n_86),
.B2(n_94),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_L g137 ( 
.A(n_124),
.B(n_117),
.Y(n_137)
);

MAJIxp5_ASAP7_75t_L g126 ( 
.A(n_111),
.B(n_98),
.C(n_54),
.Y(n_126)
);

XNOR2xp5_ASAP7_75t_L g136 ( 
.A(n_126),
.B(n_119),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_L g134 ( 
.A(n_127),
.B(n_113),
.Y(n_134)
);

AO221x1_ASAP7_75t_L g130 ( 
.A1(n_122),
.A2(n_114),
.B1(n_109),
.B2(n_104),
.C(n_106),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_SL g139 ( 
.A(n_130),
.B(n_131),
.Y(n_139)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_128),
.Y(n_131)
);

OAI22xp5_ASAP7_75t_L g142 ( 
.A1(n_134),
.A2(n_135),
.B1(n_137),
.B2(n_123),
.Y(n_142)
);

AOI22xp5_ASAP7_75t_L g135 ( 
.A1(n_129),
.A2(n_113),
.B1(n_115),
.B2(n_116),
.Y(n_135)
);

XOR2xp5_ASAP7_75t_L g141 ( 
.A(n_136),
.B(n_121),
.Y(n_141)
);

BUFx3_ASAP7_75t_L g138 ( 
.A(n_135),
.Y(n_138)
);

AND2x2_ASAP7_75t_L g140 ( 
.A(n_132),
.B(n_136),
.Y(n_140)
);

MAJIxp5_ASAP7_75t_L g144 ( 
.A(n_141),
.B(n_132),
.C(n_126),
.Y(n_144)
);

AOI211xp5_ASAP7_75t_L g145 ( 
.A1(n_142),
.A2(n_133),
.B(n_129),
.C(n_106),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_SL g143 ( 
.A(n_139),
.B(n_104),
.Y(n_143)
);

NOR2xp33_ASAP7_75t_L g147 ( 
.A(n_143),
.B(n_138),
.Y(n_147)
);

MAJIxp5_ASAP7_75t_L g146 ( 
.A(n_144),
.B(n_145),
.C(n_141),
.Y(n_146)
);

OAI21xp5_ASAP7_75t_L g149 ( 
.A1(n_146),
.A2(n_147),
.B(n_148),
.Y(n_149)
);

XNOR2xp5_ASAP7_75t_L g148 ( 
.A(n_144),
.B(n_140),
.Y(n_148)
);

BUFx24_ASAP7_75t_SL g150 ( 
.A(n_149),
.Y(n_150)
);

XOR2xp5_ASAP7_75t_L g151 ( 
.A(n_150),
.B(n_7),
.Y(n_151)
);


endmodule