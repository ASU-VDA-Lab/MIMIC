module fake_jpeg_21508_n_61 (n_3, n_2, n_1, n_0, n_4, n_6, n_5, n_61);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_6;
input n_5;

output n_61;

wire n_13;
wire n_21;
wire n_57;
wire n_53;
wire n_33;
wire n_54;
wire n_45;
wire n_10;
wire n_23;
wire n_27;
wire n_55;
wire n_22;
wire n_47;
wire n_51;
wire n_14;
wire n_40;
wire n_19;
wire n_18;
wire n_20;
wire n_59;
wire n_35;
wire n_48;
wire n_52;
wire n_46;
wire n_58;
wire n_41;
wire n_60;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_16;
wire n_49;
wire n_24;
wire n_28;
wire n_38;
wire n_26;
wire n_44;
wire n_9;
wire n_36;
wire n_11;
wire n_17;
wire n_25;
wire n_31;
wire n_56;
wire n_29;
wire n_43;
wire n_37;
wire n_50;
wire n_12;
wire n_32;
wire n_8;
wire n_15;
wire n_7;

CKINVDCx20_ASAP7_75t_R g7 ( 
.A(n_2),
.Y(n_7)
);

BUFx5_ASAP7_75t_L g8 ( 
.A(n_2),
.Y(n_8)
);

BUFx3_ASAP7_75t_L g9 ( 
.A(n_0),
.Y(n_9)
);

BUFx6f_ASAP7_75t_L g10 ( 
.A(n_6),
.Y(n_10)
);

INVx1_ASAP7_75t_L g11 ( 
.A(n_3),
.Y(n_11)
);

BUFx6f_ASAP7_75t_L g12 ( 
.A(n_2),
.Y(n_12)
);

BUFx6f_ASAP7_75t_L g13 ( 
.A(n_6),
.Y(n_13)
);

NOR2xp33_ASAP7_75t_L g14 ( 
.A(n_5),
.B(n_1),
.Y(n_14)
);

INVx1_ASAP7_75t_L g15 ( 
.A(n_11),
.Y(n_15)
);

INVx5_ASAP7_75t_SL g21 ( 
.A(n_15),
.Y(n_21)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_10),
.Y(n_16)
);

NAND2xp5_ASAP7_75t_L g20 ( 
.A(n_16),
.B(n_18),
.Y(n_20)
);

INVx5_ASAP7_75t_L g17 ( 
.A(n_12),
.Y(n_17)
);

INVx6_ASAP7_75t_L g22 ( 
.A(n_17),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_12),
.Y(n_18)
);

INVx2_ASAP7_75t_L g19 ( 
.A(n_9),
.Y(n_19)
);

AOI22xp33_ASAP7_75t_L g24 ( 
.A1(n_19),
.A2(n_8),
.B1(n_9),
.B2(n_10),
.Y(n_24)
);

OAI22xp5_ASAP7_75t_L g23 ( 
.A1(n_17),
.A2(n_7),
.B1(n_14),
.B2(n_13),
.Y(n_23)
);

OAI22xp5_ASAP7_75t_SL g27 ( 
.A1(n_23),
.A2(n_19),
.B1(n_13),
.B2(n_18),
.Y(n_27)
);

CKINVDCx16_ASAP7_75t_R g28 ( 
.A(n_24),
.Y(n_28)
);

INVx3_ASAP7_75t_L g25 ( 
.A(n_22),
.Y(n_25)
);

NOR2xp33_ASAP7_75t_L g34 ( 
.A(n_25),
.B(n_22),
.Y(n_34)
);

INVx13_ASAP7_75t_L g26 ( 
.A(n_20),
.Y(n_26)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_26),
.Y(n_30)
);

NAND2xp5_ASAP7_75t_L g31 ( 
.A(n_27),
.B(n_29),
.Y(n_31)
);

NAND2xp5_ASAP7_75t_SL g29 ( 
.A(n_20),
.B(n_0),
.Y(n_29)
);

NAND2xp5_ASAP7_75t_SL g32 ( 
.A(n_29),
.B(n_23),
.Y(n_32)
);

NOR2xp33_ASAP7_75t_L g40 ( 
.A(n_32),
.B(n_28),
.Y(n_40)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_26),
.Y(n_33)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_33),
.Y(n_37)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_34),
.Y(n_39)
);

MAJIxp5_ASAP7_75t_SL g35 ( 
.A(n_27),
.B(n_24),
.C(n_21),
.Y(n_35)
);

XNOR2xp5_ASAP7_75t_SL g38 ( 
.A(n_35),
.B(n_20),
.Y(n_38)
);

OAI22xp5_ASAP7_75t_SL g36 ( 
.A1(n_31),
.A2(n_28),
.B1(n_27),
.B2(n_26),
.Y(n_36)
);

INVxp67_ASAP7_75t_L g44 ( 
.A(n_36),
.Y(n_44)
);

A2O1A1O1Ixp25_ASAP7_75t_L g42 ( 
.A1(n_38),
.A2(n_26),
.B(n_35),
.C(n_21),
.D(n_8),
.Y(n_42)
);

NAND2xp5_ASAP7_75t_SL g45 ( 
.A(n_40),
.B(n_41),
.Y(n_45)
);

BUFx5_ASAP7_75t_L g41 ( 
.A(n_30),
.Y(n_41)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_42),
.Y(n_47)
);

AOI21xp5_ASAP7_75t_L g43 ( 
.A1(n_39),
.A2(n_21),
.B(n_0),
.Y(n_43)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_43),
.Y(n_48)
);

AOI21xp5_ASAP7_75t_L g46 ( 
.A1(n_37),
.A2(n_21),
.B(n_1),
.Y(n_46)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_46),
.Y(n_50)
);

INVx2_ASAP7_75t_L g49 ( 
.A(n_45),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_49),
.B(n_25),
.Y(n_52)
);

XOR2xp5_ASAP7_75t_L g51 ( 
.A(n_47),
.B(n_38),
.Y(n_51)
);

XNOR2xp5_ASAP7_75t_L g54 ( 
.A(n_51),
.B(n_50),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_SL g55 ( 
.A(n_52),
.B(n_53),
.Y(n_55)
);

AOI321xp33_ASAP7_75t_L g53 ( 
.A1(n_48),
.A2(n_44),
.A3(n_36),
.B1(n_41),
.B2(n_5),
.C(n_4),
.Y(n_53)
);

XNOR2xp5_ASAP7_75t_L g56 ( 
.A(n_54),
.B(n_25),
.Y(n_56)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_56),
.Y(n_58)
);

OAI21xp5_ASAP7_75t_L g57 ( 
.A1(n_55),
.A2(n_3),
.B(n_4),
.Y(n_57)
);

AOI21xp5_ASAP7_75t_SL g59 ( 
.A1(n_58),
.A2(n_57),
.B(n_1),
.Y(n_59)
);

NAND2xp33_ASAP7_75t_SL g60 ( 
.A(n_59),
.B(n_22),
.Y(n_60)
);

XOR2xp5_ASAP7_75t_L g61 ( 
.A(n_60),
.B(n_22),
.Y(n_61)
);


endmodule