module fake_netlist_5_709_n_2173 (n_137, n_294, n_431, n_318, n_380, n_419, n_444, n_469, n_82, n_194, n_316, n_389, n_418, n_248, n_124, n_86, n_136, n_146, n_315, n_268, n_451, n_408, n_61, n_376, n_503, n_127, n_75, n_235, n_226, n_74, n_57, n_353, n_351, n_367, n_452, n_397, n_493, n_111, n_483, n_155, n_43, n_116, n_22, n_467, n_423, n_284, n_46, n_245, n_21, n_501, n_139, n_38, n_105, n_280, n_4, n_378, n_17, n_382, n_254, n_33, n_23, n_302, n_265, n_293, n_372, n_443, n_244, n_47, n_173, n_198, n_447, n_247, n_314, n_368, n_433, n_8, n_321, n_292, n_100, n_455, n_417, n_212, n_385, n_498, n_507, n_119, n_497, n_275, n_252, n_26, n_295, n_133, n_330, n_508, n_506, n_2, n_6, n_509, n_39, n_147, n_373, n_67, n_307, n_439, n_87, n_150, n_106, n_209, n_259, n_448, n_375, n_301, n_68, n_93, n_186, n_134, n_191, n_51, n_63, n_492, n_171, n_153, n_399, n_341, n_204, n_394, n_250, n_260, n_298, n_320, n_505, n_286, n_122, n_282, n_331, n_10, n_24, n_406, n_470, n_325, n_449, n_132, n_90, n_101, n_281, n_240, n_381, n_189, n_220, n_291, n_231, n_257, n_390, n_31, n_456, n_13, n_371, n_481, n_152, n_317, n_9, n_323, n_195, n_42, n_356, n_227, n_45, n_271, n_94, n_335, n_123, n_370, n_167, n_234, n_343, n_308, n_379, n_428, n_267, n_514, n_457, n_297, n_156, n_5, n_225, n_377, n_484, n_219, n_442, n_157, n_131, n_192, n_223, n_392, n_158, n_138, n_264, n_109, n_472, n_454, n_387, n_374, n_163, n_276, n_339, n_95, n_183, n_185, n_243, n_398, n_396, n_347, n_169, n_59, n_255, n_215, n_350, n_196, n_459, n_211, n_218, n_400, n_181, n_436, n_3, n_290, n_221, n_178, n_386, n_287, n_344, n_473, n_422, n_475, n_72, n_104, n_41, n_415, n_56, n_141, n_485, n_496, n_355, n_486, n_15, n_336, n_145, n_48, n_50, n_337, n_430, n_313, n_88, n_479, n_510, n_216, n_168, n_395, n_164, n_432, n_311, n_208, n_142, n_214, n_328, n_140, n_299, n_303, n_369, n_296, n_241, n_357, n_184, n_446, n_445, n_65, n_78, n_144, n_114, n_96, n_165, n_468, n_499, n_213, n_129, n_342, n_482, n_98, n_361, n_464, n_363, n_402, n_413, n_197, n_107, n_69, n_236, n_388, n_1, n_249, n_304, n_329, n_203, n_274, n_384, n_460, n_80, n_35, n_73, n_277, n_92, n_19, n_338, n_149, n_477, n_461, n_333, n_309, n_30, n_512, n_14, n_84, n_462, n_130, n_322, n_258, n_29, n_79, n_151, n_25, n_306, n_458, n_288, n_188, n_190, n_201, n_263, n_471, n_44, n_224, n_40, n_34, n_228, n_283, n_383, n_474, n_112, n_85, n_463, n_488, n_502, n_239, n_466, n_420, n_489, n_55, n_49, n_310, n_54, n_504, n_511, n_12, n_465, n_76, n_358, n_362, n_170, n_332, n_27, n_77, n_102, n_161, n_273, n_349, n_270, n_230, n_81, n_118, n_279, n_70, n_253, n_261, n_174, n_289, n_172, n_206, n_217, n_440, n_478, n_441, n_450, n_312, n_476, n_429, n_345, n_210, n_494, n_365, n_91, n_176, n_182, n_143, n_83, n_354, n_480, n_237, n_425, n_513, n_407, n_180, n_340, n_207, n_37, n_346, n_393, n_229, n_108, n_487, n_495, n_437, n_66, n_177, n_60, n_403, n_453, n_421, n_16, n_0, n_58, n_405, n_18, n_359, n_490, n_117, n_326, n_233, n_404, n_205, n_366, n_113, n_246, n_179, n_125, n_410, n_269, n_128, n_285, n_412, n_120, n_232, n_327, n_135, n_126, n_202, n_266, n_272, n_491, n_427, n_193, n_251, n_352, n_53, n_160, n_426, n_409, n_500, n_154, n_62, n_148, n_71, n_300, n_435, n_159, n_334, n_391, n_434, n_175, n_262, n_238, n_99, n_411, n_414, n_319, n_364, n_20, n_121, n_242, n_360, n_36, n_200, n_162, n_64, n_222, n_28, n_89, n_438, n_115, n_324, n_416, n_199, n_187, n_32, n_401, n_103, n_348, n_97, n_166, n_11, n_424, n_7, n_256, n_305, n_52, n_278, n_110, n_2173);

input n_137;
input n_294;
input n_431;
input n_318;
input n_380;
input n_419;
input n_444;
input n_469;
input n_82;
input n_194;
input n_316;
input n_389;
input n_418;
input n_248;
input n_124;
input n_86;
input n_136;
input n_146;
input n_315;
input n_268;
input n_451;
input n_408;
input n_61;
input n_376;
input n_503;
input n_127;
input n_75;
input n_235;
input n_226;
input n_74;
input n_57;
input n_353;
input n_351;
input n_367;
input n_452;
input n_397;
input n_493;
input n_111;
input n_483;
input n_155;
input n_43;
input n_116;
input n_22;
input n_467;
input n_423;
input n_284;
input n_46;
input n_245;
input n_21;
input n_501;
input n_139;
input n_38;
input n_105;
input n_280;
input n_4;
input n_378;
input n_17;
input n_382;
input n_254;
input n_33;
input n_23;
input n_302;
input n_265;
input n_293;
input n_372;
input n_443;
input n_244;
input n_47;
input n_173;
input n_198;
input n_447;
input n_247;
input n_314;
input n_368;
input n_433;
input n_8;
input n_321;
input n_292;
input n_100;
input n_455;
input n_417;
input n_212;
input n_385;
input n_498;
input n_507;
input n_119;
input n_497;
input n_275;
input n_252;
input n_26;
input n_295;
input n_133;
input n_330;
input n_508;
input n_506;
input n_2;
input n_6;
input n_509;
input n_39;
input n_147;
input n_373;
input n_67;
input n_307;
input n_439;
input n_87;
input n_150;
input n_106;
input n_209;
input n_259;
input n_448;
input n_375;
input n_301;
input n_68;
input n_93;
input n_186;
input n_134;
input n_191;
input n_51;
input n_63;
input n_492;
input n_171;
input n_153;
input n_399;
input n_341;
input n_204;
input n_394;
input n_250;
input n_260;
input n_298;
input n_320;
input n_505;
input n_286;
input n_122;
input n_282;
input n_331;
input n_10;
input n_24;
input n_406;
input n_470;
input n_325;
input n_449;
input n_132;
input n_90;
input n_101;
input n_281;
input n_240;
input n_381;
input n_189;
input n_220;
input n_291;
input n_231;
input n_257;
input n_390;
input n_31;
input n_456;
input n_13;
input n_371;
input n_481;
input n_152;
input n_317;
input n_9;
input n_323;
input n_195;
input n_42;
input n_356;
input n_227;
input n_45;
input n_271;
input n_94;
input n_335;
input n_123;
input n_370;
input n_167;
input n_234;
input n_343;
input n_308;
input n_379;
input n_428;
input n_267;
input n_514;
input n_457;
input n_297;
input n_156;
input n_5;
input n_225;
input n_377;
input n_484;
input n_219;
input n_442;
input n_157;
input n_131;
input n_192;
input n_223;
input n_392;
input n_158;
input n_138;
input n_264;
input n_109;
input n_472;
input n_454;
input n_387;
input n_374;
input n_163;
input n_276;
input n_339;
input n_95;
input n_183;
input n_185;
input n_243;
input n_398;
input n_396;
input n_347;
input n_169;
input n_59;
input n_255;
input n_215;
input n_350;
input n_196;
input n_459;
input n_211;
input n_218;
input n_400;
input n_181;
input n_436;
input n_3;
input n_290;
input n_221;
input n_178;
input n_386;
input n_287;
input n_344;
input n_473;
input n_422;
input n_475;
input n_72;
input n_104;
input n_41;
input n_415;
input n_56;
input n_141;
input n_485;
input n_496;
input n_355;
input n_486;
input n_15;
input n_336;
input n_145;
input n_48;
input n_50;
input n_337;
input n_430;
input n_313;
input n_88;
input n_479;
input n_510;
input n_216;
input n_168;
input n_395;
input n_164;
input n_432;
input n_311;
input n_208;
input n_142;
input n_214;
input n_328;
input n_140;
input n_299;
input n_303;
input n_369;
input n_296;
input n_241;
input n_357;
input n_184;
input n_446;
input n_445;
input n_65;
input n_78;
input n_144;
input n_114;
input n_96;
input n_165;
input n_468;
input n_499;
input n_213;
input n_129;
input n_342;
input n_482;
input n_98;
input n_361;
input n_464;
input n_363;
input n_402;
input n_413;
input n_197;
input n_107;
input n_69;
input n_236;
input n_388;
input n_1;
input n_249;
input n_304;
input n_329;
input n_203;
input n_274;
input n_384;
input n_460;
input n_80;
input n_35;
input n_73;
input n_277;
input n_92;
input n_19;
input n_338;
input n_149;
input n_477;
input n_461;
input n_333;
input n_309;
input n_30;
input n_512;
input n_14;
input n_84;
input n_462;
input n_130;
input n_322;
input n_258;
input n_29;
input n_79;
input n_151;
input n_25;
input n_306;
input n_458;
input n_288;
input n_188;
input n_190;
input n_201;
input n_263;
input n_471;
input n_44;
input n_224;
input n_40;
input n_34;
input n_228;
input n_283;
input n_383;
input n_474;
input n_112;
input n_85;
input n_463;
input n_488;
input n_502;
input n_239;
input n_466;
input n_420;
input n_489;
input n_55;
input n_49;
input n_310;
input n_54;
input n_504;
input n_511;
input n_12;
input n_465;
input n_76;
input n_358;
input n_362;
input n_170;
input n_332;
input n_27;
input n_77;
input n_102;
input n_161;
input n_273;
input n_349;
input n_270;
input n_230;
input n_81;
input n_118;
input n_279;
input n_70;
input n_253;
input n_261;
input n_174;
input n_289;
input n_172;
input n_206;
input n_217;
input n_440;
input n_478;
input n_441;
input n_450;
input n_312;
input n_476;
input n_429;
input n_345;
input n_210;
input n_494;
input n_365;
input n_91;
input n_176;
input n_182;
input n_143;
input n_83;
input n_354;
input n_480;
input n_237;
input n_425;
input n_513;
input n_407;
input n_180;
input n_340;
input n_207;
input n_37;
input n_346;
input n_393;
input n_229;
input n_108;
input n_487;
input n_495;
input n_437;
input n_66;
input n_177;
input n_60;
input n_403;
input n_453;
input n_421;
input n_16;
input n_0;
input n_58;
input n_405;
input n_18;
input n_359;
input n_490;
input n_117;
input n_326;
input n_233;
input n_404;
input n_205;
input n_366;
input n_113;
input n_246;
input n_179;
input n_125;
input n_410;
input n_269;
input n_128;
input n_285;
input n_412;
input n_120;
input n_232;
input n_327;
input n_135;
input n_126;
input n_202;
input n_266;
input n_272;
input n_491;
input n_427;
input n_193;
input n_251;
input n_352;
input n_53;
input n_160;
input n_426;
input n_409;
input n_500;
input n_154;
input n_62;
input n_148;
input n_71;
input n_300;
input n_435;
input n_159;
input n_334;
input n_391;
input n_434;
input n_175;
input n_262;
input n_238;
input n_99;
input n_411;
input n_414;
input n_319;
input n_364;
input n_20;
input n_121;
input n_242;
input n_360;
input n_36;
input n_200;
input n_162;
input n_64;
input n_222;
input n_28;
input n_89;
input n_438;
input n_115;
input n_324;
input n_416;
input n_199;
input n_187;
input n_32;
input n_401;
input n_103;
input n_348;
input n_97;
input n_166;
input n_11;
input n_424;
input n_7;
input n_256;
input n_305;
input n_52;
input n_278;
input n_110;

output n_2173;

wire n_924;
wire n_1263;
wire n_977;
wire n_1378;
wire n_611;
wire n_1126;
wire n_1423;
wire n_1729;
wire n_1166;
wire n_1751;
wire n_1508;
wire n_785;
wire n_549;
wire n_532;
wire n_1161;
wire n_1859;
wire n_1677;
wire n_1150;
wire n_1780;
wire n_1488;
wire n_667;
wire n_790;
wire n_1055;
wire n_1501;
wire n_880;
wire n_544;
wire n_1007;
wire n_552;
wire n_1528;
wire n_1370;
wire n_1292;
wire n_1198;
wire n_1360;
wire n_1099;
wire n_956;
wire n_564;
wire n_1738;
wire n_2021;
wire n_2134;
wire n_1021;
wire n_1960;
wire n_551;
wire n_2143;
wire n_2059;
wire n_1323;
wire n_1466;
wire n_688;
wire n_1695;
wire n_1353;
wire n_800;
wire n_1347;
wire n_1535;
wire n_1789;
wire n_1666;
wire n_671;
wire n_819;
wire n_1451;
wire n_1022;
wire n_915;
wire n_1545;
wire n_864;
wire n_859;
wire n_951;
wire n_1947;
wire n_1264;
wire n_2114;
wire n_2001;
wire n_1494;
wire n_625;
wire n_854;
wire n_1462;
wire n_1799;
wire n_2069;
wire n_1580;
wire n_674;
wire n_1939;
wire n_1806;
wire n_516;
wire n_933;
wire n_1152;
wire n_1869;
wire n_1607;
wire n_1563;
wire n_606;
wire n_2011;
wire n_2096;
wire n_877;
wire n_2105;
wire n_2024;
wire n_1696;
wire n_755;
wire n_1118;
wire n_1686;
wire n_947;
wire n_1285;
wire n_1860;
wire n_1359;
wire n_530;
wire n_1107;
wire n_1728;
wire n_556;
wire n_2031;
wire n_2076;
wire n_1230;
wire n_668;
wire n_1896;
wire n_2165;
wire n_2147;
wire n_929;
wire n_1124;
wire n_1818;
wire n_2127;
wire n_902;
wire n_1576;
wire n_1104;
wire n_1294;
wire n_659;
wire n_1705;
wire n_1257;
wire n_1182;
wire n_579;
wire n_1698;
wire n_1261;
wire n_938;
wire n_1098;
wire n_2142;
wire n_1154;
wire n_1242;
wire n_1135;
wire n_519;
wire n_1016;
wire n_1243;
wire n_546;
wire n_2047;
wire n_1280;
wire n_1845;
wire n_2052;
wire n_2058;
wire n_731;
wire n_1483;
wire n_1314;
wire n_1512;
wire n_709;
wire n_1490;
wire n_1236;
wire n_1633;
wire n_569;
wire n_2144;
wire n_1778;
wire n_920;
wire n_1289;
wire n_1517;
wire n_2091;
wire n_2085;
wire n_1669;
wire n_976;
wire n_1949;
wire n_1449;
wire n_1946;
wire n_1566;
wire n_2032;
wire n_2149;
wire n_1078;
wire n_1670;
wire n_775;
wire n_600;
wire n_1484;
wire n_2071;
wire n_1374;
wire n_1328;
wire n_2141;
wire n_1948;
wire n_1984;
wire n_2099;
wire n_1877;
wire n_1831;
wire n_1598;
wire n_1723;
wire n_955;
wire n_1850;
wire n_1146;
wire n_882;
wire n_1036;
wire n_1097;
wire n_1749;
wire n_550;
wire n_696;
wire n_897;
wire n_798;
wire n_646;
wire n_1428;
wire n_1394;
wire n_1414;
wire n_1216;
wire n_580;
wire n_1040;
wire n_1872;
wire n_1852;
wire n_2159;
wire n_578;
wire n_926;
wire n_1218;
wire n_1931;
wire n_1547;
wire n_1070;
wire n_777;
wire n_2089;
wire n_1030;
wire n_1755;
wire n_1561;
wire n_1071;
wire n_1165;
wire n_1267;
wire n_1801;
wire n_1391;
wire n_958;
wire n_1034;
wire n_670;
wire n_1513;
wire n_1600;
wire n_521;
wire n_663;
wire n_845;
wire n_1862;
wire n_673;
wire n_837;
wire n_1239;
wire n_528;
wire n_1796;
wire n_680;
wire n_1473;
wire n_1587;
wire n_553;
wire n_901;
wire n_813;
wire n_1521;
wire n_1284;
wire n_1590;
wire n_1748;
wire n_1672;
wire n_675;
wire n_888;
wire n_1880;
wire n_1167;
wire n_1626;
wire n_637;
wire n_1384;
wire n_1556;
wire n_1863;
wire n_1064;
wire n_858;
wire n_2079;
wire n_923;
wire n_2118;
wire n_691;
wire n_1151;
wire n_881;
wire n_1405;
wire n_1706;
wire n_1582;
wire n_1069;
wire n_1784;
wire n_1075;
wire n_1836;
wire n_1450;
wire n_1322;
wire n_2101;
wire n_1471;
wire n_1986;
wire n_2072;
wire n_1750;
wire n_1459;
wire n_889;
wire n_973;
wire n_1700;
wire n_571;
wire n_1585;
wire n_1971;
wire n_1599;
wire n_1211;
wire n_1197;
wire n_1523;
wire n_1950;
wire n_907;
wire n_1447;
wire n_1377;
wire n_989;
wire n_1039;
wire n_2055;
wire n_1403;
wire n_736;
wire n_892;
wire n_1000;
wire n_1202;
wire n_1278;
wire n_2062;
wire n_1002;
wire n_1463;
wire n_1581;
wire n_2100;
wire n_593;
wire n_748;
wire n_586;
wire n_1058;
wire n_1667;
wire n_838;
wire n_1053;
wire n_1224;
wire n_1926;
wire n_1248;
wire n_1331;
wire n_953;
wire n_1014;
wire n_1241;
wire n_2150;
wire n_2152;
wire n_963;
wire n_1052;
wire n_954;
wire n_627;
wire n_1385;
wire n_793;
wire n_2140;
wire n_1819;
wire n_2139;
wire n_1527;
wire n_2042;
wire n_534;
wire n_1882;
wire n_884;
wire n_944;
wire n_1754;
wire n_1623;
wire n_1854;
wire n_1565;
wire n_1809;
wire n_1856;
wire n_647;
wire n_1072;
wire n_857;
wire n_832;
wire n_1319;
wire n_561;
wire n_2154;
wire n_1825;
wire n_1951;
wire n_1883;
wire n_1906;
wire n_1712;
wire n_1387;
wire n_1532;
wire n_1027;
wire n_971;
wire n_1156;
wire n_794;
wire n_686;
wire n_847;
wire n_1393;
wire n_596;
wire n_1775;
wire n_2028;
wire n_1368;
wire n_558;
wire n_702;
wire n_1276;
wire n_822;
wire n_1412;
wire n_1709;
wire n_2108;
wire n_728;
wire n_1162;
wire n_1538;
wire n_1838;
wire n_1199;
wire n_1847;
wire n_1779;
wire n_1884;
wire n_1038;
wire n_520;
wire n_1369;
wire n_1841;
wire n_1660;
wire n_887;
wire n_1905;
wire n_809;
wire n_870;
wire n_931;
wire n_599;
wire n_1711;
wire n_1662;
wire n_1891;
wire n_1481;
wire n_1942;
wire n_1978;
wire n_1544;
wire n_868;
wire n_639;
wire n_914;
wire n_2120;
wire n_1629;
wire n_1293;
wire n_965;
wire n_1876;
wire n_1743;
wire n_935;
wire n_817;
wire n_1175;
wire n_1479;
wire n_1810;
wire n_1888;
wire n_2009;
wire n_759;
wire n_1892;
wire n_806;
wire n_1997;
wire n_1766;
wire n_1477;
wire n_1635;
wire n_1963;
wire n_1571;
wire n_1189;
wire n_1259;
wire n_1690;
wire n_706;
wire n_746;
wire n_1649;
wire n_747;
wire n_2064;
wire n_784;
wire n_1733;
wire n_1244;
wire n_1194;
wire n_1925;
wire n_1815;
wire n_851;
wire n_615;
wire n_1759;
wire n_843;
wire n_1788;
wire n_523;
wire n_913;
wire n_1537;
wire n_705;
wire n_865;
wire n_678;
wire n_697;
wire n_1222;
wire n_1679;
wire n_776;
wire n_2022;
wire n_1798;
wire n_1790;
wire n_1415;
wire n_525;
wire n_1260;
wire n_1746;
wire n_1647;
wire n_1829;
wire n_1464;
wire n_649;
wire n_547;
wire n_1444;
wire n_1191;
wire n_1674;
wire n_1833;
wire n_1830;
wire n_2073;
wire n_1710;
wire n_1128;
wire n_1734;
wire n_744;
wire n_590;
wire n_629;
wire n_1308;
wire n_1767;
wire n_1680;
wire n_1233;
wire n_1615;
wire n_1529;
wire n_2005;
wire n_526;
wire n_1916;
wire n_677;
wire n_1333;
wire n_1121;
wire n_604;
wire n_2007;
wire n_949;
wire n_1443;
wire n_1008;
wire n_946;
wire n_1539;
wire n_1001;
wire n_1503;
wire n_2054;
wire n_1468;
wire n_1559;
wire n_1765;
wire n_1866;
wire n_689;
wire n_738;
wire n_1624;
wire n_640;
wire n_1510;
wire n_624;
wire n_1380;
wire n_1744;
wire n_1617;
wire n_1010;
wire n_1994;
wire n_1231;
wire n_739;
wire n_1279;
wire n_1406;
wire n_1195;
wire n_1837;
wire n_1839;
wire n_610;
wire n_1760;
wire n_936;
wire n_568;
wire n_1500;
wire n_1090;
wire n_757;
wire n_633;
wire n_1832;
wire n_1851;
wire n_758;
wire n_999;
wire n_2046;
wire n_1933;
wire n_1656;
wire n_1158;
wire n_2045;
wire n_1509;
wire n_1874;
wire n_2040;
wire n_563;
wire n_2060;
wire n_1987;
wire n_1145;
wire n_878;
wire n_524;
wire n_1678;
wire n_1049;
wire n_1153;
wire n_2145;
wire n_741;
wire n_1639;
wire n_1306;
wire n_1068;
wire n_1871;
wire n_1964;
wire n_1163;
wire n_906;
wire n_2039;
wire n_1207;
wire n_919;
wire n_908;
wire n_724;
wire n_1781;
wire n_2084;
wire n_2035;
wire n_658;
wire n_2061;
wire n_1740;
wire n_1362;
wire n_1586;
wire n_959;
wire n_535;
wire n_940;
wire n_1445;
wire n_1492;
wire n_2155;
wire n_1923;
wire n_1773;
wire n_592;
wire n_1169;
wire n_1692;
wire n_1596;
wire n_1017;
wire n_2171;
wire n_978;
wire n_2116;
wire n_1434;
wire n_1054;
wire n_1474;
wire n_1665;
wire n_1269;
wire n_1095;
wire n_1828;
wire n_1614;
wire n_1079;
wire n_2093;
wire n_1045;
wire n_1208;
wire n_2038;
wire n_2137;
wire n_603;
wire n_1431;
wire n_1593;
wire n_1033;
wire n_636;
wire n_660;
wire n_2087;
wire n_1640;
wire n_2162;
wire n_1732;
wire n_1009;
wire n_1148;
wire n_2051;
wire n_742;
wire n_750;
wire n_2029;
wire n_995;
wire n_2168;
wire n_1609;
wire n_1989;
wire n_1887;
wire n_1383;
wire n_1073;
wire n_662;
wire n_962;
wire n_1215;
wire n_1171;
wire n_1578;
wire n_723;
wire n_1920;
wire n_1065;
wire n_1592;
wire n_1336;
wire n_1721;
wire n_1959;
wire n_1758;
wire n_1574;
wire n_2048;
wire n_2133;
wire n_1921;
wire n_1309;
wire n_1878;
wire n_1426;
wire n_1043;
wire n_1800;
wire n_1548;
wire n_614;
wire n_1421;
wire n_1286;
wire n_1177;
wire n_1355;
wire n_974;
wire n_727;
wire n_1159;
wire n_957;
wire n_773;
wire n_2124;
wire n_743;
wire n_2081;
wire n_613;
wire n_1119;
wire n_2156;
wire n_1240;
wire n_1820;
wire n_829;
wire n_1612;
wire n_1416;
wire n_2077;
wire n_1724;
wire n_2111;
wire n_700;
wire n_1237;
wire n_573;
wire n_1420;
wire n_1132;
wire n_1366;
wire n_1300;
wire n_1127;
wire n_761;
wire n_1785;
wire n_1568;
wire n_1006;
wire n_2110;
wire n_1270;
wire n_1664;
wire n_1486;
wire n_582;
wire n_1332;
wire n_1390;
wire n_2017;
wire n_2090;
wire n_1870;
wire n_1591;
wire n_2033;
wire n_1682;
wire n_1980;
wire n_1249;
wire n_652;
wire n_1111;
wire n_1365;
wire n_1927;
wire n_2132;
wire n_1349;
wire n_1093;
wire n_1031;
wire n_609;
wire n_1041;
wire n_1265;
wire n_1909;
wire n_1562;
wire n_834;
wire n_765;
wire n_893;
wire n_1015;
wire n_1140;
wire n_891;
wire n_1651;
wire n_1965;
wire n_630;
wire n_1902;
wire n_2151;
wire n_1941;
wire n_2106;
wire n_1913;
wire n_1823;
wire n_874;
wire n_1101;
wire n_1106;
wire n_1456;
wire n_2015;
wire n_1982;
wire n_1875;
wire n_1304;
wire n_1324;
wire n_987;
wire n_1846;
wire n_2066;
wire n_1885;
wire n_1455;
wire n_767;
wire n_993;
wire n_1903;
wire n_1407;
wire n_1551;
wire n_545;
wire n_860;
wire n_1805;
wire n_1816;
wire n_948;
wire n_1217;
wire n_628;
wire n_1849;
wire n_729;
wire n_1131;
wire n_1084;
wire n_1961;
wire n_970;
wire n_1935;
wire n_911;
wire n_1430;
wire n_1094;
wire n_1354;
wire n_560;
wire n_1534;
wire n_1351;
wire n_1044;
wire n_1205;
wire n_1209;
wire n_1552;
wire n_602;
wire n_574;
wire n_1435;
wire n_879;
wire n_623;
wire n_2088;
wire n_824;
wire n_1645;
wire n_1327;
wire n_996;
wire n_921;
wire n_1684;
wire n_1717;
wire n_572;
wire n_815;
wire n_1795;
wire n_2128;
wire n_1821;
wire n_1381;
wire n_1611;
wire n_1037;
wire n_1080;
wire n_1274;
wire n_1316;
wire n_1708;
wire n_1438;
wire n_1082;
wire n_1840;
wire n_589;
wire n_716;
wire n_1630;
wire n_2122;
wire n_562;
wire n_1436;
wire n_1691;
wire n_952;
wire n_2092;
wire n_1229;
wire n_701;
wire n_1437;
wire n_1023;
wire n_2075;
wire n_645;
wire n_539;
wire n_803;
wire n_1092;
wire n_1776;
wire n_2131;
wire n_531;
wire n_1757;
wire n_890;
wire n_1897;
wire n_764;
wire n_1919;
wire n_1056;
wire n_1424;
wire n_960;
wire n_1893;
wire n_1290;
wire n_1123;
wire n_1467;
wire n_1047;
wire n_2053;
wire n_2163;
wire n_634;
wire n_1958;
wire n_1252;
wire n_1382;
wire n_1029;
wire n_925;
wire n_1206;
wire n_1311;
wire n_1519;
wire n_950;
wire n_1553;
wire n_1811;
wire n_1346;
wire n_1299;
wire n_2158;
wire n_1808;
wire n_1060;
wire n_1141;
wire n_912;
wire n_968;
wire n_619;
wire n_1386;
wire n_1699;
wire n_967;
wire n_1442;
wire n_1139;
wire n_515;
wire n_885;
wire n_1432;
wire n_1357;
wire n_2125;
wire n_683;
wire n_1632;
wire n_1057;
wire n_1051;
wire n_1085;
wire n_1066;
wire n_721;
wire n_1157;
wire n_1050;
wire n_841;
wire n_802;
wire n_1954;
wire n_1608;
wire n_983;
wire n_1844;
wire n_1305;
wire n_873;
wire n_1826;
wire n_1112;
wire n_762;
wire n_1283;
wire n_1644;
wire n_690;
wire n_1974;
wire n_583;
wire n_2086;
wire n_1343;
wire n_1203;
wire n_1631;
wire n_821;
wire n_1763;
wire n_1966;
wire n_1768;
wire n_1179;
wire n_621;
wire n_753;
wire n_1048;
wire n_1719;
wire n_1288;
wire n_1560;
wire n_1605;
wire n_1228;
wire n_2123;
wire n_972;
wire n_692;
wire n_2037;
wire n_1953;
wire n_1938;
wire n_820;
wire n_1200;
wire n_1911;
wire n_1363;
wire n_1301;
wire n_1668;
wire n_1185;
wire n_991;
wire n_828;
wire n_1967;
wire n_779;
wire n_576;
wire n_1143;
wire n_1579;
wire n_1329;
wire n_1312;
wire n_1439;
wire n_804;
wire n_537;
wire n_1688;
wire n_945;
wire n_1504;
wire n_943;
wire n_992;
wire n_1932;
wire n_543;
wire n_842;
wire n_650;
wire n_984;
wire n_694;
wire n_2082;
wire n_1992;
wire n_1643;
wire n_883;
wire n_1983;
wire n_1594;
wire n_1214;
wire n_1342;
wire n_1400;
wire n_900;
wire n_856;
wire n_1793;
wire n_1976;
wire n_918;
wire n_942;
wire n_2169;
wire n_1804;
wire n_1147;
wire n_1557;
wire n_1977;
wire n_2153;
wire n_1610;
wire n_1077;
wire n_1422;
wire n_540;
wire n_618;
wire n_896;
wire n_894;
wire n_1636;
wire n_2056;
wire n_1730;
wire n_831;
wire n_964;
wire n_1373;
wire n_1350;
wire n_1511;
wire n_1865;
wire n_1470;
wire n_1096;
wire n_2094;
wire n_1735;
wire n_1697;
wire n_1575;
wire n_833;
wire n_2020;
wire n_1646;
wire n_1307;
wire n_1881;
wire n_988;
wire n_2043;
wire n_1940;
wire n_814;
wire n_1549;
wire n_1934;
wire n_1201;
wire n_1114;
wire n_655;
wire n_2025;
wire n_1616;
wire n_1446;
wire n_669;
wire n_1458;
wire n_1176;
wire n_1472;
wire n_1807;
wire n_1149;
wire n_1671;
wire n_635;
wire n_763;
wire n_1020;
wire n_1062;
wire n_1824;
wire n_1917;
wire n_1219;
wire n_1204;
wire n_1814;
wire n_1035;
wire n_783;
wire n_555;
wire n_1928;
wire n_1848;
wire n_2126;
wire n_1188;
wire n_1722;
wire n_661;
wire n_1802;
wire n_849;
wire n_584;
wire n_681;
wire n_1638;
wire n_1786;
wire n_2002;
wire n_830;
wire n_2098;
wire n_1296;
wire n_1413;
wire n_801;
wire n_2080;
wire n_2068;
wire n_875;
wire n_1110;
wire n_1655;
wire n_749;
wire n_1895;
wire n_1134;
wire n_1358;
wire n_717;
wire n_939;
wire n_1088;
wire n_588;
wire n_1173;
wire n_789;
wire n_1232;
wire n_1603;
wire n_734;
wire n_638;
wire n_866;
wire n_969;
wire n_1401;
wire n_1019;
wire n_1105;
wire n_1998;
wire n_1338;
wire n_577;
wire n_2016;
wire n_1522;
wire n_1687;
wire n_1637;
wire n_2034;
wire n_1419;
wire n_1653;
wire n_693;
wire n_1506;
wire n_836;
wire n_990;
wire n_1886;
wire n_1389;
wire n_1894;
wire n_975;
wire n_1908;
wire n_1256;
wire n_1702;
wire n_567;
wire n_1465;
wire n_778;
wire n_1122;
wire n_770;
wire n_1375;
wire n_1102;
wire n_1843;
wire n_711;
wire n_1499;
wire n_1187;
wire n_1441;
wire n_1392;
wire n_1597;
wire n_1929;
wire n_1164;
wire n_1659;
wire n_1834;
wire n_2097;
wire n_1174;
wire n_1371;
wire n_617;
wire n_1303;
wire n_2063;
wire n_1572;
wire n_1968;
wire n_876;
wire n_1516;
wire n_1190;
wire n_1736;
wire n_1685;
wire n_917;
wire n_601;
wire n_1714;
wire n_966;
wire n_1116;
wire n_2000;
wire n_1661;
wire n_1212;
wire n_2074;
wire n_1541;
wire n_726;
wire n_982;
wire n_1573;
wire n_1453;
wire n_1731;
wire n_818;
wire n_1970;
wire n_861;
wire n_1713;
wire n_1183;
wire n_1658;
wire n_899;
wire n_1253;
wire n_1737;
wire n_2117;
wire n_1904;
wire n_1993;
wire n_774;
wire n_1628;
wire n_1335;
wire n_1514;
wire n_1777;
wire n_1957;
wire n_1059;
wire n_1345;
wire n_1133;
wire n_1912;
wire n_1771;
wire n_1899;
wire n_557;
wire n_1410;
wire n_1005;
wire n_607;
wire n_1003;
wire n_679;
wire n_710;
wire n_2067;
wire n_527;
wire n_707;
wire n_1168;
wire n_2148;
wire n_937;
wire n_1427;
wire n_1584;
wire n_665;
wire n_1726;
wire n_1835;
wire n_1440;
wire n_2164;
wire n_1988;
wire n_2115;
wire n_1853;
wire n_1356;
wire n_1787;
wire n_910;
wire n_1657;
wire n_768;
wire n_1475;
wire n_1302;
wire n_1774;
wire n_1725;
wire n_1313;
wire n_1136;
wire n_1491;
wire n_754;
wire n_1496;
wire n_1125;
wire n_708;
wire n_529;
wire n_1812;
wire n_735;
wire n_1915;
wire n_1109;
wire n_895;
wire n_1310;
wire n_2121;
wire n_1803;
wire n_1399;
wire n_1543;
wire n_1991;
wire n_1979;
wire n_791;
wire n_732;
wire n_1533;
wire n_808;
wire n_797;
wire n_1025;
wire n_1930;
wire n_1955;
wire n_1067;
wire n_1720;
wire n_2003;
wire n_766;
wire n_1457;
wire n_541;
wire n_538;
wire n_2008;
wire n_1117;
wire n_799;
wire n_687;
wire n_715;
wire n_1742;
wire n_1480;
wire n_1482;
wire n_1213;
wire n_1266;
wire n_536;
wire n_872;
wire n_2012;
wire n_594;
wire n_1291;
wire n_1297;
wire n_1753;
wire n_1782;
wire n_1155;
wire n_1418;
wire n_1972;
wire n_1524;
wire n_1689;
wire n_1485;
wire n_1011;
wire n_1184;
wire n_985;
wire n_1855;
wire n_869;
wire n_810;
wire n_827;
wire n_1703;
wire n_1352;
wire n_626;
wire n_1650;
wire n_1144;
wire n_1137;
wire n_1570;
wire n_1170;
wire n_2023;
wire n_2095;
wire n_676;
wire n_2103;
wire n_653;
wire n_2160;
wire n_642;
wire n_1602;
wire n_855;
wire n_1178;
wire n_1461;
wire n_850;
wire n_684;
wire n_664;
wire n_1999;
wire n_2065;
wire n_2136;
wire n_1372;
wire n_605;
wire n_1273;
wire n_1822;
wire n_620;
wire n_643;
wire n_916;
wire n_1081;
wire n_1235;
wire n_980;
wire n_698;
wire n_703;
wire n_1115;
wire n_1282;
wire n_1318;
wire n_1783;
wire n_780;
wire n_998;
wire n_1454;
wire n_1227;
wire n_1531;
wire n_840;
wire n_1334;
wire n_1907;
wire n_823;
wire n_725;
wire n_1388;
wire n_1417;
wire n_1295;
wire n_672;
wire n_1985;
wire n_1898;
wire n_2107;
wire n_581;
wire n_554;
wire n_1625;
wire n_2130;
wire n_898;
wire n_1762;
wire n_1013;
wire n_1452;
wire n_718;
wire n_1120;
wire n_719;
wire n_1791;
wire n_1890;
wire n_1747;
wire n_714;
wire n_1683;
wire n_1944;
wire n_909;
wire n_1817;
wire n_1530;
wire n_1497;
wire n_997;
wire n_932;
wire n_612;
wire n_2078;
wire n_1409;
wire n_788;
wire n_1326;
wire n_1268;
wire n_559;
wire n_825;
wire n_1981;
wire n_1320;
wire n_1663;
wire n_737;
wire n_1718;
wire n_986;
wire n_1317;
wire n_1518;
wire n_1715;
wire n_2102;
wire n_1281;
wire n_1952;
wire n_1192;
wire n_1024;
wire n_1063;
wire n_1889;
wire n_1792;
wire n_1564;
wire n_1868;
wire n_1613;
wire n_733;
wire n_1489;
wire n_1922;
wire n_1376;
wire n_941;
wire n_981;
wire n_1569;
wire n_867;
wire n_587;
wire n_792;
wire n_756;
wire n_1429;
wire n_1238;
wire n_548;
wire n_812;
wire n_2104;
wire n_518;
wire n_2057;
wire n_1772;
wire n_752;
wire n_905;
wire n_1476;
wire n_1108;
wire n_782;
wire n_1100;
wire n_1861;
wire n_2129;
wire n_1395;
wire n_862;
wire n_1425;
wire n_760;
wire n_1901;
wire n_1900;
wire n_1620;
wire n_1330;
wire n_1867;
wire n_1945;
wire n_1675;
wire n_1924;
wire n_1727;
wire n_1554;
wire n_1745;
wire n_769;
wire n_2006;
wire n_1995;
wire n_2138;
wire n_1046;
wire n_934;
wire n_1618;
wire n_826;
wire n_1813;
wire n_886;
wire n_2014;
wire n_1221;
wire n_654;
wire n_1172;
wire n_1341;
wire n_570;
wire n_1641;
wire n_1361;
wire n_1707;
wire n_853;
wire n_751;
wire n_2172;
wire n_1973;
wire n_786;
wire n_1083;
wire n_1142;
wire n_1129;
wire n_704;
wire n_787;
wire n_1770;
wire n_961;
wire n_1756;
wire n_771;
wire n_1716;
wire n_1225;
wire n_1520;
wire n_522;
wire n_1287;
wire n_1262;
wire n_930;
wire n_1873;
wire n_1411;
wire n_622;
wire n_1962;
wire n_1577;
wire n_1087;
wire n_994;
wire n_1701;
wire n_848;
wire n_1550;
wire n_1498;
wire n_2167;
wire n_1223;
wire n_1272;
wire n_682;
wire n_1567;
wire n_1247;
wire n_922;
wire n_816;
wire n_1648;
wire n_591;
wire n_1536;
wire n_1857;
wire n_1344;
wire n_2041;
wire n_631;
wire n_1246;
wire n_1339;
wire n_1478;
wire n_1797;
wire n_1769;
wire n_839;
wire n_1210;
wire n_1364;
wire n_1250;
wire n_1842;
wire n_871;
wire n_685;
wire n_598;
wire n_608;
wire n_928;
wire n_1367;
wire n_1943;
wire n_1460;
wire n_772;
wire n_2018;
wire n_1555;
wire n_1589;
wire n_517;
wire n_1086;
wire n_796;
wire n_1858;
wire n_1619;
wire n_2119;
wire n_1502;
wire n_2157;
wire n_1469;
wire n_1012;
wire n_1396;
wire n_1348;
wire n_2030;
wire n_903;
wire n_1525;
wire n_1752;
wire n_740;
wire n_1404;
wire n_1794;
wire n_1315;
wire n_1061;
wire n_1910;
wire n_1298;
wire n_1652;
wire n_2050;
wire n_1193;
wire n_1676;
wire n_1255;
wire n_1113;
wire n_1226;
wire n_722;
wire n_1277;
wire n_2146;
wire n_844;
wire n_852;
wire n_1487;
wire n_1864;
wire n_1028;
wire n_1601;
wire n_781;
wire n_542;
wire n_1546;
wire n_595;
wire n_1337;
wire n_1495;
wire n_632;
wire n_699;
wire n_979;
wire n_1515;
wire n_1627;
wire n_1245;
wire n_846;
wire n_1673;
wire n_1321;
wire n_1975;
wire n_2070;
wire n_1937;
wire n_585;
wire n_2112;
wire n_1739;
wire n_616;
wire n_1914;
wire n_2135;
wire n_745;
wire n_1654;
wire n_1103;
wire n_648;
wire n_1379;
wire n_2170;
wire n_1076;
wire n_1091;
wire n_1408;
wire n_1761;
wire n_641;
wire n_730;
wire n_2036;
wire n_1325;
wire n_1595;
wire n_2161;
wire n_575;
wire n_795;
wire n_2083;
wire n_695;
wire n_656;
wire n_1606;
wire n_1220;
wire n_1694;
wire n_1540;
wire n_1936;
wire n_1956;
wire n_1642;
wire n_2027;
wire n_1130;
wire n_720;
wire n_1918;
wire n_1526;
wire n_863;
wire n_805;
wire n_1604;
wire n_1275;
wire n_1764;
wire n_712;
wire n_1583;
wire n_1042;
wire n_1402;
wire n_2049;
wire n_1493;
wire n_657;
wire n_644;
wire n_1741;
wire n_1160;
wire n_1397;
wire n_1258;
wire n_1074;
wire n_2004;
wire n_1621;
wire n_2113;
wire n_566;
wire n_565;
wire n_1448;
wire n_1507;
wire n_1398;
wire n_1879;
wire n_597;
wire n_1996;
wire n_1181;
wire n_1505;
wire n_1634;
wire n_1196;
wire n_2019;
wire n_651;
wire n_1340;
wire n_811;
wire n_1558;
wire n_807;
wire n_2166;
wire n_835;
wire n_666;
wire n_1433;
wire n_1704;
wire n_1254;
wire n_1026;
wire n_2026;
wire n_1969;
wire n_1234;
wire n_2109;
wire n_1138;
wire n_927;
wire n_1089;
wire n_2013;
wire n_1990;
wire n_2044;
wire n_1004;
wire n_1186;
wire n_1032;
wire n_1681;
wire n_2010;
wire n_1018;
wire n_1693;
wire n_713;
wire n_904;
wire n_1588;
wire n_1622;
wire n_1180;
wire n_1827;
wire n_1271;
wire n_533;
wire n_1542;
wire n_1251;

INVx2_ASAP7_75t_L g515 ( 
.A(n_157),
.Y(n_515)
);

INVx1_ASAP7_75t_L g516 ( 
.A(n_391),
.Y(n_516)
);

CKINVDCx5p33_ASAP7_75t_R g517 ( 
.A(n_298),
.Y(n_517)
);

INVx1_ASAP7_75t_L g518 ( 
.A(n_450),
.Y(n_518)
);

CKINVDCx20_ASAP7_75t_R g519 ( 
.A(n_281),
.Y(n_519)
);

CKINVDCx5p33_ASAP7_75t_R g520 ( 
.A(n_47),
.Y(n_520)
);

INVx1_ASAP7_75t_L g521 ( 
.A(n_494),
.Y(n_521)
);

INVx1_ASAP7_75t_L g522 ( 
.A(n_51),
.Y(n_522)
);

INVx1_ASAP7_75t_L g523 ( 
.A(n_230),
.Y(n_523)
);

INVx1_ASAP7_75t_L g524 ( 
.A(n_301),
.Y(n_524)
);

INVx1_ASAP7_75t_L g525 ( 
.A(n_231),
.Y(n_525)
);

CKINVDCx5p33_ASAP7_75t_R g526 ( 
.A(n_454),
.Y(n_526)
);

CKINVDCx5p33_ASAP7_75t_R g527 ( 
.A(n_36),
.Y(n_527)
);

INVx1_ASAP7_75t_L g528 ( 
.A(n_146),
.Y(n_528)
);

CKINVDCx5p33_ASAP7_75t_R g529 ( 
.A(n_164),
.Y(n_529)
);

CKINVDCx20_ASAP7_75t_R g530 ( 
.A(n_315),
.Y(n_530)
);

CKINVDCx5p33_ASAP7_75t_R g531 ( 
.A(n_380),
.Y(n_531)
);

CKINVDCx20_ASAP7_75t_R g532 ( 
.A(n_362),
.Y(n_532)
);

CKINVDCx16_ASAP7_75t_R g533 ( 
.A(n_152),
.Y(n_533)
);

INVx1_ASAP7_75t_L g534 ( 
.A(n_411),
.Y(n_534)
);

CKINVDCx5p33_ASAP7_75t_R g535 ( 
.A(n_273),
.Y(n_535)
);

INVx1_ASAP7_75t_L g536 ( 
.A(n_79),
.Y(n_536)
);

CKINVDCx5p33_ASAP7_75t_R g537 ( 
.A(n_348),
.Y(n_537)
);

CKINVDCx5p33_ASAP7_75t_R g538 ( 
.A(n_198),
.Y(n_538)
);

INVx2_ASAP7_75t_SL g539 ( 
.A(n_505),
.Y(n_539)
);

CKINVDCx16_ASAP7_75t_R g540 ( 
.A(n_473),
.Y(n_540)
);

CKINVDCx5p33_ASAP7_75t_R g541 ( 
.A(n_58),
.Y(n_541)
);

CKINVDCx5p33_ASAP7_75t_R g542 ( 
.A(n_408),
.Y(n_542)
);

CKINVDCx5p33_ASAP7_75t_R g543 ( 
.A(n_268),
.Y(n_543)
);

CKINVDCx20_ASAP7_75t_R g544 ( 
.A(n_350),
.Y(n_544)
);

CKINVDCx5p33_ASAP7_75t_R g545 ( 
.A(n_44),
.Y(n_545)
);

CKINVDCx5p33_ASAP7_75t_R g546 ( 
.A(n_352),
.Y(n_546)
);

CKINVDCx5p33_ASAP7_75t_R g547 ( 
.A(n_172),
.Y(n_547)
);

BUFx6f_ASAP7_75t_L g548 ( 
.A(n_510),
.Y(n_548)
);

CKINVDCx20_ASAP7_75t_R g549 ( 
.A(n_198),
.Y(n_549)
);

CKINVDCx5p33_ASAP7_75t_R g550 ( 
.A(n_125),
.Y(n_550)
);

BUFx10_ASAP7_75t_L g551 ( 
.A(n_493),
.Y(n_551)
);

INVx1_ASAP7_75t_L g552 ( 
.A(n_99),
.Y(n_552)
);

INVx1_ASAP7_75t_L g553 ( 
.A(n_307),
.Y(n_553)
);

CKINVDCx5p33_ASAP7_75t_R g554 ( 
.A(n_73),
.Y(n_554)
);

CKINVDCx5p33_ASAP7_75t_R g555 ( 
.A(n_328),
.Y(n_555)
);

CKINVDCx5p33_ASAP7_75t_R g556 ( 
.A(n_138),
.Y(n_556)
);

CKINVDCx20_ASAP7_75t_R g557 ( 
.A(n_444),
.Y(n_557)
);

INVx1_ASAP7_75t_L g558 ( 
.A(n_335),
.Y(n_558)
);

BUFx3_ASAP7_75t_L g559 ( 
.A(n_455),
.Y(n_559)
);

CKINVDCx5p33_ASAP7_75t_R g560 ( 
.A(n_316),
.Y(n_560)
);

CKINVDCx5p33_ASAP7_75t_R g561 ( 
.A(n_253),
.Y(n_561)
);

BUFx10_ASAP7_75t_L g562 ( 
.A(n_126),
.Y(n_562)
);

CKINVDCx5p33_ASAP7_75t_R g563 ( 
.A(n_324),
.Y(n_563)
);

INVx1_ASAP7_75t_L g564 ( 
.A(n_246),
.Y(n_564)
);

CKINVDCx5p33_ASAP7_75t_R g565 ( 
.A(n_141),
.Y(n_565)
);

INVx1_ASAP7_75t_L g566 ( 
.A(n_395),
.Y(n_566)
);

CKINVDCx5p33_ASAP7_75t_R g567 ( 
.A(n_490),
.Y(n_567)
);

INVx1_ASAP7_75t_L g568 ( 
.A(n_92),
.Y(n_568)
);

BUFx6f_ASAP7_75t_L g569 ( 
.A(n_318),
.Y(n_569)
);

INVx1_ASAP7_75t_L g570 ( 
.A(n_68),
.Y(n_570)
);

CKINVDCx5p33_ASAP7_75t_R g571 ( 
.A(n_159),
.Y(n_571)
);

INVx1_ASAP7_75t_L g572 ( 
.A(n_500),
.Y(n_572)
);

INVx1_ASAP7_75t_L g573 ( 
.A(n_32),
.Y(n_573)
);

CKINVDCx5p33_ASAP7_75t_R g574 ( 
.A(n_135),
.Y(n_574)
);

CKINVDCx20_ASAP7_75t_R g575 ( 
.A(n_385),
.Y(n_575)
);

BUFx3_ASAP7_75t_L g576 ( 
.A(n_400),
.Y(n_576)
);

BUFx6f_ASAP7_75t_L g577 ( 
.A(n_122),
.Y(n_577)
);

INVx1_ASAP7_75t_L g578 ( 
.A(n_249),
.Y(n_578)
);

CKINVDCx5p33_ASAP7_75t_R g579 ( 
.A(n_487),
.Y(n_579)
);

INVx1_ASAP7_75t_L g580 ( 
.A(n_241),
.Y(n_580)
);

INVx2_ASAP7_75t_L g581 ( 
.A(n_274),
.Y(n_581)
);

CKINVDCx5p33_ASAP7_75t_R g582 ( 
.A(n_44),
.Y(n_582)
);

CKINVDCx5p33_ASAP7_75t_R g583 ( 
.A(n_488),
.Y(n_583)
);

INVx1_ASAP7_75t_L g584 ( 
.A(n_492),
.Y(n_584)
);

INVx1_ASAP7_75t_L g585 ( 
.A(n_491),
.Y(n_585)
);

INVx1_ASAP7_75t_L g586 ( 
.A(n_203),
.Y(n_586)
);

CKINVDCx5p33_ASAP7_75t_R g587 ( 
.A(n_50),
.Y(n_587)
);

CKINVDCx5p33_ASAP7_75t_R g588 ( 
.A(n_451),
.Y(n_588)
);

CKINVDCx5p33_ASAP7_75t_R g589 ( 
.A(n_293),
.Y(n_589)
);

INVx1_ASAP7_75t_L g590 ( 
.A(n_367),
.Y(n_590)
);

CKINVDCx5p33_ASAP7_75t_R g591 ( 
.A(n_167),
.Y(n_591)
);

CKINVDCx20_ASAP7_75t_R g592 ( 
.A(n_428),
.Y(n_592)
);

CKINVDCx5p33_ASAP7_75t_R g593 ( 
.A(n_122),
.Y(n_593)
);

INVx2_ASAP7_75t_L g594 ( 
.A(n_419),
.Y(n_594)
);

INVx1_ASAP7_75t_L g595 ( 
.A(n_381),
.Y(n_595)
);

INVx1_ASAP7_75t_L g596 ( 
.A(n_10),
.Y(n_596)
);

INVx2_ASAP7_75t_L g597 ( 
.A(n_113),
.Y(n_597)
);

CKINVDCx5p33_ASAP7_75t_R g598 ( 
.A(n_453),
.Y(n_598)
);

CKINVDCx20_ASAP7_75t_R g599 ( 
.A(n_175),
.Y(n_599)
);

CKINVDCx5p33_ASAP7_75t_R g600 ( 
.A(n_247),
.Y(n_600)
);

CKINVDCx5p33_ASAP7_75t_R g601 ( 
.A(n_6),
.Y(n_601)
);

INVx1_ASAP7_75t_L g602 ( 
.A(n_250),
.Y(n_602)
);

INVx1_ASAP7_75t_L g603 ( 
.A(n_503),
.Y(n_603)
);

INVx1_ASAP7_75t_L g604 ( 
.A(n_407),
.Y(n_604)
);

INVx1_ASAP7_75t_L g605 ( 
.A(n_248),
.Y(n_605)
);

INVx1_ASAP7_75t_L g606 ( 
.A(n_277),
.Y(n_606)
);

INVx1_ASAP7_75t_L g607 ( 
.A(n_48),
.Y(n_607)
);

INVx2_ASAP7_75t_SL g608 ( 
.A(n_512),
.Y(n_608)
);

CKINVDCx5p33_ASAP7_75t_R g609 ( 
.A(n_364),
.Y(n_609)
);

CKINVDCx5p33_ASAP7_75t_R g610 ( 
.A(n_351),
.Y(n_610)
);

INVx1_ASAP7_75t_L g611 ( 
.A(n_93),
.Y(n_611)
);

BUFx3_ASAP7_75t_L g612 ( 
.A(n_311),
.Y(n_612)
);

CKINVDCx5p33_ASAP7_75t_R g613 ( 
.A(n_43),
.Y(n_613)
);

INVx1_ASAP7_75t_L g614 ( 
.A(n_346),
.Y(n_614)
);

CKINVDCx5p33_ASAP7_75t_R g615 ( 
.A(n_495),
.Y(n_615)
);

INVx1_ASAP7_75t_L g616 ( 
.A(n_464),
.Y(n_616)
);

BUFx10_ASAP7_75t_L g617 ( 
.A(n_412),
.Y(n_617)
);

CKINVDCx5p33_ASAP7_75t_R g618 ( 
.A(n_235),
.Y(n_618)
);

CKINVDCx20_ASAP7_75t_R g619 ( 
.A(n_341),
.Y(n_619)
);

INVx1_ASAP7_75t_L g620 ( 
.A(n_4),
.Y(n_620)
);

BUFx10_ASAP7_75t_L g621 ( 
.A(n_363),
.Y(n_621)
);

INVx3_ASAP7_75t_L g622 ( 
.A(n_449),
.Y(n_622)
);

CKINVDCx16_ASAP7_75t_R g623 ( 
.A(n_479),
.Y(n_623)
);

CKINVDCx5p33_ASAP7_75t_R g624 ( 
.A(n_80),
.Y(n_624)
);

CKINVDCx5p33_ASAP7_75t_R g625 ( 
.A(n_257),
.Y(n_625)
);

INVx1_ASAP7_75t_SL g626 ( 
.A(n_285),
.Y(n_626)
);

CKINVDCx5p33_ASAP7_75t_R g627 ( 
.A(n_71),
.Y(n_627)
);

CKINVDCx5p33_ASAP7_75t_R g628 ( 
.A(n_152),
.Y(n_628)
);

CKINVDCx5p33_ASAP7_75t_R g629 ( 
.A(n_471),
.Y(n_629)
);

CKINVDCx5p33_ASAP7_75t_R g630 ( 
.A(n_137),
.Y(n_630)
);

INVx1_ASAP7_75t_L g631 ( 
.A(n_459),
.Y(n_631)
);

INVx1_ASAP7_75t_L g632 ( 
.A(n_489),
.Y(n_632)
);

INVx1_ASAP7_75t_L g633 ( 
.A(n_448),
.Y(n_633)
);

CKINVDCx5p33_ASAP7_75t_R g634 ( 
.A(n_470),
.Y(n_634)
);

CKINVDCx5p33_ASAP7_75t_R g635 ( 
.A(n_251),
.Y(n_635)
);

CKINVDCx20_ASAP7_75t_R g636 ( 
.A(n_24),
.Y(n_636)
);

INVx2_ASAP7_75t_L g637 ( 
.A(n_374),
.Y(n_637)
);

CKINVDCx5p33_ASAP7_75t_R g638 ( 
.A(n_14),
.Y(n_638)
);

CKINVDCx5p33_ASAP7_75t_R g639 ( 
.A(n_420),
.Y(n_639)
);

INVx1_ASAP7_75t_SL g640 ( 
.A(n_460),
.Y(n_640)
);

INVx1_ASAP7_75t_L g641 ( 
.A(n_462),
.Y(n_641)
);

INVx1_ASAP7_75t_L g642 ( 
.A(n_33),
.Y(n_642)
);

INVx2_ASAP7_75t_L g643 ( 
.A(n_394),
.Y(n_643)
);

CKINVDCx5p33_ASAP7_75t_R g644 ( 
.A(n_163),
.Y(n_644)
);

CKINVDCx5p33_ASAP7_75t_R g645 ( 
.A(n_514),
.Y(n_645)
);

INVx1_ASAP7_75t_L g646 ( 
.A(n_238),
.Y(n_646)
);

INVx1_ASAP7_75t_SL g647 ( 
.A(n_182),
.Y(n_647)
);

CKINVDCx5p33_ASAP7_75t_R g648 ( 
.A(n_47),
.Y(n_648)
);

INVx1_ASAP7_75t_L g649 ( 
.A(n_17),
.Y(n_649)
);

BUFx3_ASAP7_75t_L g650 ( 
.A(n_112),
.Y(n_650)
);

INVx1_ASAP7_75t_L g651 ( 
.A(n_21),
.Y(n_651)
);

INVx1_ASAP7_75t_L g652 ( 
.A(n_313),
.Y(n_652)
);

CKINVDCx20_ASAP7_75t_R g653 ( 
.A(n_5),
.Y(n_653)
);

CKINVDCx5p33_ASAP7_75t_R g654 ( 
.A(n_210),
.Y(n_654)
);

INVx2_ASAP7_75t_L g655 ( 
.A(n_279),
.Y(n_655)
);

INVx1_ASAP7_75t_L g656 ( 
.A(n_17),
.Y(n_656)
);

CKINVDCx5p33_ASAP7_75t_R g657 ( 
.A(n_427),
.Y(n_657)
);

INVx2_ASAP7_75t_L g658 ( 
.A(n_347),
.Y(n_658)
);

INVx1_ASAP7_75t_L g659 ( 
.A(n_349),
.Y(n_659)
);

BUFx10_ASAP7_75t_L g660 ( 
.A(n_233),
.Y(n_660)
);

CKINVDCx5p33_ASAP7_75t_R g661 ( 
.A(n_266),
.Y(n_661)
);

INVx1_ASAP7_75t_SL g662 ( 
.A(n_323),
.Y(n_662)
);

INVx1_ASAP7_75t_L g663 ( 
.A(n_147),
.Y(n_663)
);

INVx1_ASAP7_75t_L g664 ( 
.A(n_144),
.Y(n_664)
);

INVx1_ASAP7_75t_L g665 ( 
.A(n_320),
.Y(n_665)
);

CKINVDCx5p33_ASAP7_75t_R g666 ( 
.A(n_357),
.Y(n_666)
);

INVx1_ASAP7_75t_L g667 ( 
.A(n_111),
.Y(n_667)
);

INVx1_ASAP7_75t_L g668 ( 
.A(n_439),
.Y(n_668)
);

CKINVDCx5p33_ASAP7_75t_R g669 ( 
.A(n_221),
.Y(n_669)
);

CKINVDCx5p33_ASAP7_75t_R g670 ( 
.A(n_234),
.Y(n_670)
);

BUFx2_ASAP7_75t_L g671 ( 
.A(n_339),
.Y(n_671)
);

CKINVDCx5p33_ASAP7_75t_R g672 ( 
.A(n_498),
.Y(n_672)
);

CKINVDCx20_ASAP7_75t_R g673 ( 
.A(n_458),
.Y(n_673)
);

CKINVDCx5p33_ASAP7_75t_R g674 ( 
.A(n_221),
.Y(n_674)
);

CKINVDCx5p33_ASAP7_75t_R g675 ( 
.A(n_138),
.Y(n_675)
);

INVx1_ASAP7_75t_L g676 ( 
.A(n_329),
.Y(n_676)
);

CKINVDCx14_ASAP7_75t_R g677 ( 
.A(n_343),
.Y(n_677)
);

CKINVDCx5p33_ASAP7_75t_R g678 ( 
.A(n_366),
.Y(n_678)
);

CKINVDCx5p33_ASAP7_75t_R g679 ( 
.A(n_446),
.Y(n_679)
);

CKINVDCx5p33_ASAP7_75t_R g680 ( 
.A(n_452),
.Y(n_680)
);

BUFx2_ASAP7_75t_L g681 ( 
.A(n_226),
.Y(n_681)
);

CKINVDCx5p33_ASAP7_75t_R g682 ( 
.A(n_0),
.Y(n_682)
);

CKINVDCx20_ASAP7_75t_R g683 ( 
.A(n_398),
.Y(n_683)
);

BUFx8_ASAP7_75t_SL g684 ( 
.A(n_319),
.Y(n_684)
);

INVx1_ASAP7_75t_L g685 ( 
.A(n_466),
.Y(n_685)
);

CKINVDCx5p33_ASAP7_75t_R g686 ( 
.A(n_206),
.Y(n_686)
);

INVx1_ASAP7_75t_L g687 ( 
.A(n_305),
.Y(n_687)
);

INVx1_ASAP7_75t_L g688 ( 
.A(n_93),
.Y(n_688)
);

BUFx3_ASAP7_75t_L g689 ( 
.A(n_124),
.Y(n_689)
);

INVx2_ASAP7_75t_L g690 ( 
.A(n_299),
.Y(n_690)
);

INVx1_ASAP7_75t_L g691 ( 
.A(n_239),
.Y(n_691)
);

BUFx10_ASAP7_75t_L g692 ( 
.A(n_159),
.Y(n_692)
);

HB1xp67_ASAP7_75t_L g693 ( 
.A(n_128),
.Y(n_693)
);

CKINVDCx20_ASAP7_75t_R g694 ( 
.A(n_45),
.Y(n_694)
);

INVx1_ASAP7_75t_L g695 ( 
.A(n_61),
.Y(n_695)
);

CKINVDCx5p33_ASAP7_75t_R g696 ( 
.A(n_110),
.Y(n_696)
);

INVx1_ASAP7_75t_L g697 ( 
.A(n_10),
.Y(n_697)
);

CKINVDCx5p33_ASAP7_75t_R g698 ( 
.A(n_402),
.Y(n_698)
);

INVx1_ASAP7_75t_L g699 ( 
.A(n_496),
.Y(n_699)
);

CKINVDCx14_ASAP7_75t_R g700 ( 
.A(n_265),
.Y(n_700)
);

INVx2_ASAP7_75t_L g701 ( 
.A(n_497),
.Y(n_701)
);

INVx1_ASAP7_75t_SL g702 ( 
.A(n_282),
.Y(n_702)
);

CKINVDCx5p33_ASAP7_75t_R g703 ( 
.A(n_263),
.Y(n_703)
);

INVx1_ASAP7_75t_L g704 ( 
.A(n_354),
.Y(n_704)
);

CKINVDCx5p33_ASAP7_75t_R g705 ( 
.A(n_147),
.Y(n_705)
);

INVx1_ASAP7_75t_L g706 ( 
.A(n_372),
.Y(n_706)
);

CKINVDCx5p33_ASAP7_75t_R g707 ( 
.A(n_486),
.Y(n_707)
);

INVx1_ASAP7_75t_L g708 ( 
.A(n_172),
.Y(n_708)
);

CKINVDCx5p33_ASAP7_75t_R g709 ( 
.A(n_43),
.Y(n_709)
);

CKINVDCx5p33_ASAP7_75t_R g710 ( 
.A(n_340),
.Y(n_710)
);

CKINVDCx5p33_ASAP7_75t_R g711 ( 
.A(n_361),
.Y(n_711)
);

INVx1_ASAP7_75t_L g712 ( 
.A(n_396),
.Y(n_712)
);

BUFx2_ASAP7_75t_SL g713 ( 
.A(n_264),
.Y(n_713)
);

INVx1_ASAP7_75t_L g714 ( 
.A(n_297),
.Y(n_714)
);

BUFx2_ASAP7_75t_L g715 ( 
.A(n_204),
.Y(n_715)
);

CKINVDCx16_ASAP7_75t_R g716 ( 
.A(n_94),
.Y(n_716)
);

CKINVDCx5p33_ASAP7_75t_R g717 ( 
.A(n_392),
.Y(n_717)
);

CKINVDCx5p33_ASAP7_75t_R g718 ( 
.A(n_227),
.Y(n_718)
);

INVx2_ASAP7_75t_SL g719 ( 
.A(n_166),
.Y(n_719)
);

INVx1_ASAP7_75t_L g720 ( 
.A(n_24),
.Y(n_720)
);

INVx1_ASAP7_75t_L g721 ( 
.A(n_650),
.Y(n_721)
);

BUFx6f_ASAP7_75t_L g722 ( 
.A(n_548),
.Y(n_722)
);

INVx1_ASAP7_75t_L g723 ( 
.A(n_650),
.Y(n_723)
);

INVx1_ASAP7_75t_L g724 ( 
.A(n_689),
.Y(n_724)
);

INVx1_ASAP7_75t_L g725 ( 
.A(n_689),
.Y(n_725)
);

INVx1_ASAP7_75t_SL g726 ( 
.A(n_715),
.Y(n_726)
);

INVx1_ASAP7_75t_L g727 ( 
.A(n_577),
.Y(n_727)
);

BUFx2_ASAP7_75t_SL g728 ( 
.A(n_619),
.Y(n_728)
);

INVx1_ASAP7_75t_L g729 ( 
.A(n_577),
.Y(n_729)
);

INVxp33_ASAP7_75t_SL g730 ( 
.A(n_693),
.Y(n_730)
);

INVx1_ASAP7_75t_L g731 ( 
.A(n_577),
.Y(n_731)
);

CKINVDCx16_ASAP7_75t_R g732 ( 
.A(n_533),
.Y(n_732)
);

INVx1_ASAP7_75t_L g733 ( 
.A(n_522),
.Y(n_733)
);

INVx1_ASAP7_75t_L g734 ( 
.A(n_528),
.Y(n_734)
);

INVx1_ASAP7_75t_L g735 ( 
.A(n_536),
.Y(n_735)
);

INVxp67_ASAP7_75t_SL g736 ( 
.A(n_671),
.Y(n_736)
);

INVxp67_ASAP7_75t_SL g737 ( 
.A(n_681),
.Y(n_737)
);

INVx1_ASAP7_75t_L g738 ( 
.A(n_552),
.Y(n_738)
);

INVxp67_ASAP7_75t_SL g739 ( 
.A(n_559),
.Y(n_739)
);

CKINVDCx20_ASAP7_75t_R g740 ( 
.A(n_599),
.Y(n_740)
);

CKINVDCx16_ASAP7_75t_R g741 ( 
.A(n_716),
.Y(n_741)
);

INVx1_ASAP7_75t_L g742 ( 
.A(n_568),
.Y(n_742)
);

INVx1_ASAP7_75t_L g743 ( 
.A(n_570),
.Y(n_743)
);

INVx1_ASAP7_75t_L g744 ( 
.A(n_573),
.Y(n_744)
);

INVx1_ASAP7_75t_L g745 ( 
.A(n_586),
.Y(n_745)
);

INVx1_ASAP7_75t_L g746 ( 
.A(n_596),
.Y(n_746)
);

INVx1_ASAP7_75t_L g747 ( 
.A(n_607),
.Y(n_747)
);

INVx1_ASAP7_75t_L g748 ( 
.A(n_611),
.Y(n_748)
);

CKINVDCx20_ASAP7_75t_R g749 ( 
.A(n_599),
.Y(n_749)
);

INVx1_ASAP7_75t_L g750 ( 
.A(n_620),
.Y(n_750)
);

INVxp33_ASAP7_75t_SL g751 ( 
.A(n_520),
.Y(n_751)
);

INVx2_ASAP7_75t_L g752 ( 
.A(n_515),
.Y(n_752)
);

INVx1_ASAP7_75t_L g753 ( 
.A(n_642),
.Y(n_753)
);

HB1xp67_ASAP7_75t_L g754 ( 
.A(n_527),
.Y(n_754)
);

CKINVDCx5p33_ASAP7_75t_R g755 ( 
.A(n_517),
.Y(n_755)
);

INVxp67_ASAP7_75t_L g756 ( 
.A(n_562),
.Y(n_756)
);

INVxp33_ASAP7_75t_SL g757 ( 
.A(n_529),
.Y(n_757)
);

INVxp33_ASAP7_75t_SL g758 ( 
.A(n_538),
.Y(n_758)
);

INVx1_ASAP7_75t_L g759 ( 
.A(n_649),
.Y(n_759)
);

INVxp67_ASAP7_75t_SL g760 ( 
.A(n_559),
.Y(n_760)
);

INVxp33_ASAP7_75t_L g761 ( 
.A(n_515),
.Y(n_761)
);

INVx1_ASAP7_75t_L g762 ( 
.A(n_651),
.Y(n_762)
);

INVx1_ASAP7_75t_L g763 ( 
.A(n_656),
.Y(n_763)
);

BUFx6f_ASAP7_75t_L g764 ( 
.A(n_548),
.Y(n_764)
);

INVxp67_ASAP7_75t_SL g765 ( 
.A(n_576),
.Y(n_765)
);

INVx1_ASAP7_75t_L g766 ( 
.A(n_663),
.Y(n_766)
);

INVx1_ASAP7_75t_L g767 ( 
.A(n_664),
.Y(n_767)
);

INVxp33_ASAP7_75t_SL g768 ( 
.A(n_541),
.Y(n_768)
);

INVx1_ASAP7_75t_L g769 ( 
.A(n_667),
.Y(n_769)
);

CKINVDCx5p33_ASAP7_75t_R g770 ( 
.A(n_526),
.Y(n_770)
);

INVx1_ASAP7_75t_SL g771 ( 
.A(n_549),
.Y(n_771)
);

INVxp67_ASAP7_75t_L g772 ( 
.A(n_562),
.Y(n_772)
);

CKINVDCx20_ASAP7_75t_R g773 ( 
.A(n_636),
.Y(n_773)
);

INVxp33_ASAP7_75t_L g774 ( 
.A(n_597),
.Y(n_774)
);

INVx2_ASAP7_75t_L g775 ( 
.A(n_597),
.Y(n_775)
);

INVx1_ASAP7_75t_L g776 ( 
.A(n_688),
.Y(n_776)
);

INVx1_ASAP7_75t_L g777 ( 
.A(n_695),
.Y(n_777)
);

INVx1_ASAP7_75t_L g778 ( 
.A(n_697),
.Y(n_778)
);

INVx1_ASAP7_75t_L g779 ( 
.A(n_708),
.Y(n_779)
);

INVxp33_ASAP7_75t_L g780 ( 
.A(n_720),
.Y(n_780)
);

INVxp67_ASAP7_75t_SL g781 ( 
.A(n_576),
.Y(n_781)
);

BUFx3_ASAP7_75t_L g782 ( 
.A(n_612),
.Y(n_782)
);

INVxp33_ASAP7_75t_L g783 ( 
.A(n_684),
.Y(n_783)
);

CKINVDCx16_ASAP7_75t_R g784 ( 
.A(n_540),
.Y(n_784)
);

INVxp67_ASAP7_75t_SL g785 ( 
.A(n_612),
.Y(n_785)
);

INVx1_ASAP7_75t_L g786 ( 
.A(n_516),
.Y(n_786)
);

INVx1_ASAP7_75t_L g787 ( 
.A(n_518),
.Y(n_787)
);

INVxp67_ASAP7_75t_SL g788 ( 
.A(n_622),
.Y(n_788)
);

INVx1_ASAP7_75t_L g789 ( 
.A(n_521),
.Y(n_789)
);

INVxp67_ASAP7_75t_SL g790 ( 
.A(n_622),
.Y(n_790)
);

INVx1_ASAP7_75t_L g791 ( 
.A(n_523),
.Y(n_791)
);

CKINVDCx20_ASAP7_75t_R g792 ( 
.A(n_636),
.Y(n_792)
);

INVxp67_ASAP7_75t_SL g793 ( 
.A(n_524),
.Y(n_793)
);

CKINVDCx5p33_ASAP7_75t_R g794 ( 
.A(n_531),
.Y(n_794)
);

HB1xp67_ASAP7_75t_L g795 ( 
.A(n_545),
.Y(n_795)
);

CKINVDCx20_ASAP7_75t_R g796 ( 
.A(n_653),
.Y(n_796)
);

INVx1_ASAP7_75t_L g797 ( 
.A(n_525),
.Y(n_797)
);

INVx1_ASAP7_75t_L g798 ( 
.A(n_534),
.Y(n_798)
);

INVx1_ASAP7_75t_L g799 ( 
.A(n_553),
.Y(n_799)
);

CKINVDCx5p33_ASAP7_75t_R g800 ( 
.A(n_535),
.Y(n_800)
);

INVxp33_ASAP7_75t_SL g801 ( 
.A(n_547),
.Y(n_801)
);

INVx1_ASAP7_75t_L g802 ( 
.A(n_558),
.Y(n_802)
);

CKINVDCx20_ASAP7_75t_R g803 ( 
.A(n_694),
.Y(n_803)
);

INVx1_ASAP7_75t_L g804 ( 
.A(n_564),
.Y(n_804)
);

CKINVDCx5p33_ASAP7_75t_R g805 ( 
.A(n_537),
.Y(n_805)
);

INVx1_ASAP7_75t_L g806 ( 
.A(n_566),
.Y(n_806)
);

INVx1_ASAP7_75t_L g807 ( 
.A(n_572),
.Y(n_807)
);

CKINVDCx20_ASAP7_75t_R g808 ( 
.A(n_619),
.Y(n_808)
);

INVx1_ASAP7_75t_L g809 ( 
.A(n_578),
.Y(n_809)
);

INVx1_ASAP7_75t_L g810 ( 
.A(n_580),
.Y(n_810)
);

INVx1_ASAP7_75t_L g811 ( 
.A(n_584),
.Y(n_811)
);

INVxp33_ASAP7_75t_L g812 ( 
.A(n_684),
.Y(n_812)
);

INVx1_ASAP7_75t_L g813 ( 
.A(n_585),
.Y(n_813)
);

HB1xp67_ASAP7_75t_L g814 ( 
.A(n_550),
.Y(n_814)
);

INVx1_ASAP7_75t_L g815 ( 
.A(n_590),
.Y(n_815)
);

INVx1_ASAP7_75t_L g816 ( 
.A(n_595),
.Y(n_816)
);

BUFx8_ASAP7_75t_L g817 ( 
.A(n_782),
.Y(n_817)
);

INVx2_ASAP7_75t_L g818 ( 
.A(n_722),
.Y(n_818)
);

INVx1_ASAP7_75t_L g819 ( 
.A(n_727),
.Y(n_819)
);

OAI22xp5_ASAP7_75t_SL g820 ( 
.A1(n_740),
.A2(n_673),
.B1(n_647),
.B2(n_556),
.Y(n_820)
);

BUFx2_ASAP7_75t_L g821 ( 
.A(n_756),
.Y(n_821)
);

BUFx2_ASAP7_75t_L g822 ( 
.A(n_772),
.Y(n_822)
);

NAND2xp5_ASAP7_75t_L g823 ( 
.A(n_755),
.B(n_539),
.Y(n_823)
);

AND2x4_ASAP7_75t_L g824 ( 
.A(n_788),
.B(n_608),
.Y(n_824)
);

BUFx6f_ASAP7_75t_L g825 ( 
.A(n_722),
.Y(n_825)
);

BUFx3_ASAP7_75t_L g826 ( 
.A(n_782),
.Y(n_826)
);

INVx2_ASAP7_75t_L g827 ( 
.A(n_722),
.Y(n_827)
);

AOI22xp5_ASAP7_75t_L g828 ( 
.A1(n_730),
.A2(n_677),
.B1(n_700),
.B2(n_623),
.Y(n_828)
);

BUFx12f_ASAP7_75t_L g829 ( 
.A(n_770),
.Y(n_829)
);

INVx1_ASAP7_75t_L g830 ( 
.A(n_729),
.Y(n_830)
);

OAI22x1_ASAP7_75t_L g831 ( 
.A1(n_726),
.A2(n_719),
.B1(n_565),
.B2(n_571),
.Y(n_831)
);

INVx2_ASAP7_75t_L g832 ( 
.A(n_722),
.Y(n_832)
);

INVx2_ASAP7_75t_L g833 ( 
.A(n_764),
.Y(n_833)
);

INVx1_ASAP7_75t_L g834 ( 
.A(n_731),
.Y(n_834)
);

BUFx3_ASAP7_75t_L g835 ( 
.A(n_721),
.Y(n_835)
);

INVx3_ASAP7_75t_L g836 ( 
.A(n_764),
.Y(n_836)
);

INVx2_ASAP7_75t_SL g837 ( 
.A(n_754),
.Y(n_837)
);

BUFx6f_ASAP7_75t_L g838 ( 
.A(n_764),
.Y(n_838)
);

CKINVDCx20_ASAP7_75t_R g839 ( 
.A(n_808),
.Y(n_839)
);

AND2x2_ASAP7_75t_SL g840 ( 
.A(n_784),
.B(n_581),
.Y(n_840)
);

BUFx6f_ASAP7_75t_L g841 ( 
.A(n_764),
.Y(n_841)
);

INVx2_ASAP7_75t_L g842 ( 
.A(n_752),
.Y(n_842)
);

AND2x2_ASAP7_75t_L g843 ( 
.A(n_739),
.B(n_700),
.Y(n_843)
);

NAND2xp5_ASAP7_75t_L g844 ( 
.A(n_794),
.B(n_581),
.Y(n_844)
);

BUFx6f_ASAP7_75t_L g845 ( 
.A(n_752),
.Y(n_845)
);

NOR2xp33_ASAP7_75t_L g846 ( 
.A(n_757),
.B(n_626),
.Y(n_846)
);

BUFx6f_ASAP7_75t_L g847 ( 
.A(n_775),
.Y(n_847)
);

AND2x4_ASAP7_75t_L g848 ( 
.A(n_790),
.B(n_594),
.Y(n_848)
);

BUFx6f_ASAP7_75t_L g849 ( 
.A(n_775),
.Y(n_849)
);

INVx2_ASAP7_75t_L g850 ( 
.A(n_786),
.Y(n_850)
);

INVx1_ASAP7_75t_L g851 ( 
.A(n_787),
.Y(n_851)
);

INVx1_ASAP7_75t_L g852 ( 
.A(n_789),
.Y(n_852)
);

NAND2xp5_ASAP7_75t_L g853 ( 
.A(n_800),
.B(n_594),
.Y(n_853)
);

HB1xp67_ASAP7_75t_L g854 ( 
.A(n_732),
.Y(n_854)
);

NOR2x1_ASAP7_75t_L g855 ( 
.A(n_791),
.B(n_713),
.Y(n_855)
);

AOI22xp5_ASAP7_75t_L g856 ( 
.A1(n_741),
.A2(n_673),
.B1(n_530),
.B2(n_532),
.Y(n_856)
);

BUFx3_ASAP7_75t_L g857 ( 
.A(n_723),
.Y(n_857)
);

OA21x2_ASAP7_75t_L g858 ( 
.A1(n_797),
.A2(n_643),
.B(n_637),
.Y(n_858)
);

INVx2_ASAP7_75t_L g859 ( 
.A(n_798),
.Y(n_859)
);

BUFx6f_ASAP7_75t_L g860 ( 
.A(n_799),
.Y(n_860)
);

CKINVDCx5p33_ASAP7_75t_R g861 ( 
.A(n_728),
.Y(n_861)
);

AND2x2_ASAP7_75t_L g862 ( 
.A(n_760),
.B(n_551),
.Y(n_862)
);

INVx2_ASAP7_75t_L g863 ( 
.A(n_802),
.Y(n_863)
);

OAI21x1_ASAP7_75t_L g864 ( 
.A1(n_804),
.A2(n_643),
.B(n_637),
.Y(n_864)
);

OA21x2_ASAP7_75t_L g865 ( 
.A1(n_806),
.A2(n_658),
.B(n_655),
.Y(n_865)
);

OAI22x1_ASAP7_75t_R g866 ( 
.A1(n_740),
.A2(n_773),
.B1(n_792),
.B2(n_749),
.Y(n_866)
);

AND2x4_ASAP7_75t_L g867 ( 
.A(n_793),
.B(n_655),
.Y(n_867)
);

CKINVDCx5p33_ASAP7_75t_R g868 ( 
.A(n_805),
.Y(n_868)
);

AND2x4_ASAP7_75t_L g869 ( 
.A(n_765),
.B(n_658),
.Y(n_869)
);

AND2x2_ASAP7_75t_L g870 ( 
.A(n_781),
.B(n_551),
.Y(n_870)
);

INVx2_ASAP7_75t_L g871 ( 
.A(n_807),
.Y(n_871)
);

BUFx6f_ASAP7_75t_L g872 ( 
.A(n_809),
.Y(n_872)
);

INVx2_ASAP7_75t_L g873 ( 
.A(n_810),
.Y(n_873)
);

INVx2_ASAP7_75t_L g874 ( 
.A(n_811),
.Y(n_874)
);

INVx1_ASAP7_75t_L g875 ( 
.A(n_813),
.Y(n_875)
);

INVx1_ASAP7_75t_L g876 ( 
.A(n_815),
.Y(n_876)
);

OAI21x1_ASAP7_75t_L g877 ( 
.A1(n_816),
.A2(n_701),
.B(n_690),
.Y(n_877)
);

INVx3_ASAP7_75t_L g878 ( 
.A(n_733),
.Y(n_878)
);

INVx1_ASAP7_75t_L g879 ( 
.A(n_851),
.Y(n_879)
);

INVx2_ASAP7_75t_L g880 ( 
.A(n_845),
.Y(n_880)
);

INVx2_ASAP7_75t_L g881 ( 
.A(n_845),
.Y(n_881)
);

INVx1_ASAP7_75t_L g882 ( 
.A(n_852),
.Y(n_882)
);

BUFx8_ASAP7_75t_L g883 ( 
.A(n_829),
.Y(n_883)
);

INVx2_ASAP7_75t_L g884 ( 
.A(n_845),
.Y(n_884)
);

INVx1_ASAP7_75t_SL g885 ( 
.A(n_821),
.Y(n_885)
);

BUFx6f_ASAP7_75t_L g886 ( 
.A(n_825),
.Y(n_886)
);

INVx2_ASAP7_75t_L g887 ( 
.A(n_845),
.Y(n_887)
);

OAI22xp5_ASAP7_75t_L g888 ( 
.A1(n_828),
.A2(n_737),
.B1(n_736),
.B2(n_761),
.Y(n_888)
);

BUFx6f_ASAP7_75t_L g889 ( 
.A(n_825),
.Y(n_889)
);

BUFx6f_ASAP7_75t_L g890 ( 
.A(n_825),
.Y(n_890)
);

INVx1_ASAP7_75t_L g891 ( 
.A(n_875),
.Y(n_891)
);

NAND2xp5_ASAP7_75t_L g892 ( 
.A(n_858),
.B(n_785),
.Y(n_892)
);

AND2x4_ASAP7_75t_L g893 ( 
.A(n_826),
.B(n_724),
.Y(n_893)
);

BUFx2_ASAP7_75t_L g894 ( 
.A(n_854),
.Y(n_894)
);

NAND2xp5_ASAP7_75t_L g895 ( 
.A(n_858),
.B(n_690),
.Y(n_895)
);

INVx1_ASAP7_75t_L g896 ( 
.A(n_876),
.Y(n_896)
);

INVx2_ASAP7_75t_L g897 ( 
.A(n_845),
.Y(n_897)
);

INVx2_ASAP7_75t_L g898 ( 
.A(n_847),
.Y(n_898)
);

INVx3_ASAP7_75t_L g899 ( 
.A(n_825),
.Y(n_899)
);

CKINVDCx16_ASAP7_75t_R g900 ( 
.A(n_866),
.Y(n_900)
);

INVx2_ASAP7_75t_L g901 ( 
.A(n_847),
.Y(n_901)
);

INVx1_ASAP7_75t_L g902 ( 
.A(n_835),
.Y(n_902)
);

BUFx6f_ASAP7_75t_L g903 ( 
.A(n_825),
.Y(n_903)
);

INVx1_ASAP7_75t_L g904 ( 
.A(n_857),
.Y(n_904)
);

NAND2x1p5_ASAP7_75t_L g905 ( 
.A(n_869),
.B(n_640),
.Y(n_905)
);

OAI22xp5_ASAP7_75t_L g906 ( 
.A1(n_846),
.A2(n_774),
.B1(n_761),
.B2(n_780),
.Y(n_906)
);

INVx1_ASAP7_75t_L g907 ( 
.A(n_857),
.Y(n_907)
);

INVx2_ASAP7_75t_L g908 ( 
.A(n_847),
.Y(n_908)
);

INVx1_ASAP7_75t_L g909 ( 
.A(n_860),
.Y(n_909)
);

INVxp67_ASAP7_75t_L g910 ( 
.A(n_821),
.Y(n_910)
);

NAND2xp33_ASAP7_75t_SL g911 ( 
.A(n_831),
.B(n_519),
.Y(n_911)
);

INVx2_ASAP7_75t_L g912 ( 
.A(n_847),
.Y(n_912)
);

INVxp67_ASAP7_75t_L g913 ( 
.A(n_822),
.Y(n_913)
);

NAND2xp5_ASAP7_75t_L g914 ( 
.A(n_858),
.B(n_701),
.Y(n_914)
);

NAND2xp5_ASAP7_75t_L g915 ( 
.A(n_865),
.B(n_725),
.Y(n_915)
);

INVx1_ASAP7_75t_SL g916 ( 
.A(n_822),
.Y(n_916)
);

INVx1_ASAP7_75t_L g917 ( 
.A(n_860),
.Y(n_917)
);

AND2x2_ASAP7_75t_L g918 ( 
.A(n_843),
.B(n_795),
.Y(n_918)
);

INVx2_ASAP7_75t_L g919 ( 
.A(n_849),
.Y(n_919)
);

CKINVDCx20_ASAP7_75t_R g920 ( 
.A(n_839),
.Y(n_920)
);

INVx1_ASAP7_75t_L g921 ( 
.A(n_860),
.Y(n_921)
);

INVx1_ASAP7_75t_L g922 ( 
.A(n_872),
.Y(n_922)
);

OA21x2_ASAP7_75t_L g923 ( 
.A1(n_864),
.A2(n_603),
.B(n_602),
.Y(n_923)
);

INVx2_ASAP7_75t_L g924 ( 
.A(n_849),
.Y(n_924)
);

INVx1_ASAP7_75t_L g925 ( 
.A(n_872),
.Y(n_925)
);

OA21x2_ASAP7_75t_L g926 ( 
.A1(n_864),
.A2(n_605),
.B(n_604),
.Y(n_926)
);

AND2x4_ASAP7_75t_L g927 ( 
.A(n_826),
.B(n_734),
.Y(n_927)
);

AOI22xp5_ASAP7_75t_L g928 ( 
.A1(n_840),
.A2(n_758),
.B1(n_768),
.B2(n_751),
.Y(n_928)
);

INVx2_ASAP7_75t_L g929 ( 
.A(n_849),
.Y(n_929)
);

OAI22xp5_ASAP7_75t_SL g930 ( 
.A1(n_820),
.A2(n_808),
.B1(n_773),
.B2(n_792),
.Y(n_930)
);

INVx2_ASAP7_75t_L g931 ( 
.A(n_849),
.Y(n_931)
);

NAND2xp5_ASAP7_75t_L g932 ( 
.A(n_865),
.B(n_606),
.Y(n_932)
);

NAND2xp5_ASAP7_75t_SL g933 ( 
.A(n_840),
.B(n_869),
.Y(n_933)
);

INVx2_ASAP7_75t_L g934 ( 
.A(n_836),
.Y(n_934)
);

INVx2_ASAP7_75t_L g935 ( 
.A(n_836),
.Y(n_935)
);

AND2x4_ASAP7_75t_L g936 ( 
.A(n_848),
.B(n_735),
.Y(n_936)
);

INVx2_ASAP7_75t_L g937 ( 
.A(n_818),
.Y(n_937)
);

INVx1_ASAP7_75t_L g938 ( 
.A(n_872),
.Y(n_938)
);

INVxp67_ASAP7_75t_L g939 ( 
.A(n_843),
.Y(n_939)
);

INVx1_ASAP7_75t_L g940 ( 
.A(n_850),
.Y(n_940)
);

BUFx6f_ASAP7_75t_L g941 ( 
.A(n_838),
.Y(n_941)
);

INVxp67_ASAP7_75t_L g942 ( 
.A(n_862),
.Y(n_942)
);

AND2x2_ASAP7_75t_L g943 ( 
.A(n_837),
.B(n_814),
.Y(n_943)
);

AND2x2_ASAP7_75t_L g944 ( 
.A(n_837),
.B(n_774),
.Y(n_944)
);

AND2x6_ASAP7_75t_L g945 ( 
.A(n_848),
.B(n_548),
.Y(n_945)
);

OAI22xp5_ASAP7_75t_L g946 ( 
.A1(n_856),
.A2(n_780),
.B1(n_554),
.B2(n_582),
.Y(n_946)
);

NAND2xp5_ASAP7_75t_L g947 ( 
.A(n_865),
.B(n_614),
.Y(n_947)
);

NOR2xp33_ASAP7_75t_SL g948 ( 
.A(n_868),
.B(n_544),
.Y(n_948)
);

NAND2xp5_ASAP7_75t_SL g949 ( 
.A(n_869),
.B(n_548),
.Y(n_949)
);

BUFx6f_ASAP7_75t_L g950 ( 
.A(n_838),
.Y(n_950)
);

CKINVDCx20_ASAP7_75t_R g951 ( 
.A(n_839),
.Y(n_951)
);

CKINVDCx16_ASAP7_75t_R g952 ( 
.A(n_829),
.Y(n_952)
);

NAND2xp5_ASAP7_75t_L g953 ( 
.A(n_848),
.B(n_616),
.Y(n_953)
);

NAND2xp5_ASAP7_75t_L g954 ( 
.A(n_867),
.B(n_631),
.Y(n_954)
);

AND2x6_ASAP7_75t_L g955 ( 
.A(n_867),
.B(n_862),
.Y(n_955)
);

INVx1_ASAP7_75t_L g956 ( 
.A(n_850),
.Y(n_956)
);

INVx2_ASAP7_75t_L g957 ( 
.A(n_940),
.Y(n_957)
);

INVx4_ASAP7_75t_L g958 ( 
.A(n_893),
.Y(n_958)
);

INVx1_ASAP7_75t_L g959 ( 
.A(n_879),
.Y(n_959)
);

NOR2xp33_ASAP7_75t_L g960 ( 
.A(n_942),
.B(n_868),
.Y(n_960)
);

INVx1_ASAP7_75t_L g961 ( 
.A(n_882),
.Y(n_961)
);

NOR2xp33_ASAP7_75t_L g962 ( 
.A(n_942),
.B(n_801),
.Y(n_962)
);

NOR2xp33_ASAP7_75t_L g963 ( 
.A(n_939),
.B(n_751),
.Y(n_963)
);

INVx2_ASAP7_75t_SL g964 ( 
.A(n_944),
.Y(n_964)
);

INVx1_ASAP7_75t_L g965 ( 
.A(n_891),
.Y(n_965)
);

BUFx10_ASAP7_75t_L g966 ( 
.A(n_893),
.Y(n_966)
);

AND2x6_ASAP7_75t_L g967 ( 
.A(n_915),
.B(n_870),
.Y(n_967)
);

OR2x2_ASAP7_75t_L g968 ( 
.A(n_885),
.B(n_771),
.Y(n_968)
);

INVx1_ASAP7_75t_L g969 ( 
.A(n_896),
.Y(n_969)
);

NAND2xp5_ASAP7_75t_L g970 ( 
.A(n_955),
.B(n_824),
.Y(n_970)
);

INVx4_ASAP7_75t_SL g971 ( 
.A(n_945),
.Y(n_971)
);

INVx1_ASAP7_75t_L g972 ( 
.A(n_956),
.Y(n_972)
);

AOI22xp5_ASAP7_75t_L g973 ( 
.A1(n_955),
.A2(n_824),
.B1(n_853),
.B2(n_844),
.Y(n_973)
);

NAND2xp5_ASAP7_75t_L g974 ( 
.A(n_955),
.B(n_824),
.Y(n_974)
);

INVx5_ASAP7_75t_L g975 ( 
.A(n_945),
.Y(n_975)
);

NAND2xp5_ASAP7_75t_SL g976 ( 
.A(n_906),
.B(n_861),
.Y(n_976)
);

CKINVDCx5p33_ASAP7_75t_R g977 ( 
.A(n_952),
.Y(n_977)
);

CKINVDCx5p33_ASAP7_75t_R g978 ( 
.A(n_920),
.Y(n_978)
);

INVxp33_ASAP7_75t_L g979 ( 
.A(n_943),
.Y(n_979)
);

AND2x2_ASAP7_75t_L g980 ( 
.A(n_885),
.B(n_870),
.Y(n_980)
);

BUFx4f_ASAP7_75t_L g981 ( 
.A(n_894),
.Y(n_981)
);

OAI22xp33_ASAP7_75t_L g982 ( 
.A1(n_933),
.A2(n_823),
.B1(n_861),
.B2(n_812),
.Y(n_982)
);

NAND2xp5_ASAP7_75t_L g983 ( 
.A(n_955),
.B(n_867),
.Y(n_983)
);

INVx2_ASAP7_75t_L g984 ( 
.A(n_937),
.Y(n_984)
);

INVx1_ASAP7_75t_L g985 ( 
.A(n_927),
.Y(n_985)
);

AND2x2_ASAP7_75t_L g986 ( 
.A(n_916),
.B(n_918),
.Y(n_986)
);

NAND2xp5_ASAP7_75t_SL g987 ( 
.A(n_905),
.B(n_768),
.Y(n_987)
);

AO22x2_ASAP7_75t_L g988 ( 
.A1(n_888),
.A2(n_831),
.B1(n_702),
.B2(n_662),
.Y(n_988)
);

NOR2xp33_ASAP7_75t_SL g989 ( 
.A(n_916),
.B(n_557),
.Y(n_989)
);

OR2x6_ASAP7_75t_L g990 ( 
.A(n_930),
.B(n_738),
.Y(n_990)
);

INVx2_ASAP7_75t_L g991 ( 
.A(n_934),
.Y(n_991)
);

INVx2_ASAP7_75t_L g992 ( 
.A(n_935),
.Y(n_992)
);

INVx1_ASAP7_75t_L g993 ( 
.A(n_927),
.Y(n_993)
);

AOI22xp33_ASAP7_75t_L g994 ( 
.A1(n_892),
.A2(n_633),
.B1(n_641),
.B2(n_632),
.Y(n_994)
);

INVx1_ASAP7_75t_L g995 ( 
.A(n_902),
.Y(n_995)
);

INVx1_ASAP7_75t_L g996 ( 
.A(n_904),
.Y(n_996)
);

INVx1_ASAP7_75t_L g997 ( 
.A(n_907),
.Y(n_997)
);

INVx2_ASAP7_75t_L g998 ( 
.A(n_899),
.Y(n_998)
);

INVx2_ASAP7_75t_L g999 ( 
.A(n_886),
.Y(n_999)
);

OR2x2_ASAP7_75t_L g1000 ( 
.A(n_910),
.B(n_783),
.Y(n_1000)
);

INVx2_ASAP7_75t_SL g1001 ( 
.A(n_936),
.Y(n_1001)
);

NOR2xp33_ASAP7_75t_L g1002 ( 
.A(n_910),
.B(n_783),
.Y(n_1002)
);

BUFx6f_ASAP7_75t_L g1003 ( 
.A(n_886),
.Y(n_1003)
);

NAND2xp5_ASAP7_75t_L g1004 ( 
.A(n_892),
.B(n_855),
.Y(n_1004)
);

INVx2_ASAP7_75t_L g1005 ( 
.A(n_889),
.Y(n_1005)
);

INVx6_ASAP7_75t_L g1006 ( 
.A(n_883),
.Y(n_1006)
);

INVx2_ASAP7_75t_L g1007 ( 
.A(n_889),
.Y(n_1007)
);

BUFx6f_ASAP7_75t_SL g1008 ( 
.A(n_883),
.Y(n_1008)
);

INVxp67_ASAP7_75t_L g1009 ( 
.A(n_948),
.Y(n_1009)
);

INVx1_ASAP7_75t_L g1010 ( 
.A(n_915),
.Y(n_1010)
);

INVx2_ASAP7_75t_SL g1011 ( 
.A(n_905),
.Y(n_1011)
);

AND2x4_ASAP7_75t_L g1012 ( 
.A(n_953),
.B(n_859),
.Y(n_1012)
);

INVx2_ASAP7_75t_SL g1013 ( 
.A(n_954),
.Y(n_1013)
);

INVx1_ASAP7_75t_L g1014 ( 
.A(n_953),
.Y(n_1014)
);

INVx5_ASAP7_75t_L g1015 ( 
.A(n_945),
.Y(n_1015)
);

INVx2_ASAP7_75t_L g1016 ( 
.A(n_889),
.Y(n_1016)
);

NAND2xp5_ASAP7_75t_SL g1017 ( 
.A(n_928),
.B(n_817),
.Y(n_1017)
);

INVx1_ASAP7_75t_L g1018 ( 
.A(n_954),
.Y(n_1018)
);

INVx4_ASAP7_75t_L g1019 ( 
.A(n_890),
.Y(n_1019)
);

BUFx3_ASAP7_75t_L g1020 ( 
.A(n_920),
.Y(n_1020)
);

NAND2xp5_ASAP7_75t_L g1021 ( 
.A(n_895),
.B(n_878),
.Y(n_1021)
);

NOR2xp33_ASAP7_75t_L g1022 ( 
.A(n_913),
.B(n_796),
.Y(n_1022)
);

NAND2xp33_ASAP7_75t_L g1023 ( 
.A(n_945),
.B(n_542),
.Y(n_1023)
);

AND2x6_ASAP7_75t_L g1024 ( 
.A(n_895),
.B(n_569),
.Y(n_1024)
);

BUFx2_ASAP7_75t_L g1025 ( 
.A(n_951),
.Y(n_1025)
);

AND2x6_ASAP7_75t_L g1026 ( 
.A(n_914),
.B(n_569),
.Y(n_1026)
);

INVx1_ASAP7_75t_L g1027 ( 
.A(n_949),
.Y(n_1027)
);

BUFx3_ASAP7_75t_L g1028 ( 
.A(n_951),
.Y(n_1028)
);

INVx4_ASAP7_75t_L g1029 ( 
.A(n_890),
.Y(n_1029)
);

INVx5_ASAP7_75t_L g1030 ( 
.A(n_945),
.Y(n_1030)
);

INVx3_ASAP7_75t_L g1031 ( 
.A(n_903),
.Y(n_1031)
);

INVx6_ASAP7_75t_L g1032 ( 
.A(n_900),
.Y(n_1032)
);

NOR2xp33_ASAP7_75t_L g1033 ( 
.A(n_888),
.B(n_796),
.Y(n_1033)
);

INVx4_ASAP7_75t_L g1034 ( 
.A(n_903),
.Y(n_1034)
);

NOR2xp33_ASAP7_75t_L g1035 ( 
.A(n_948),
.B(n_803),
.Y(n_1035)
);

INVx1_ASAP7_75t_L g1036 ( 
.A(n_949),
.Y(n_1036)
);

NAND2xp5_ASAP7_75t_SL g1037 ( 
.A(n_946),
.B(n_817),
.Y(n_1037)
);

NAND2xp5_ASAP7_75t_SL g1038 ( 
.A(n_946),
.B(n_817),
.Y(n_1038)
);

INVx4_ASAP7_75t_L g1039 ( 
.A(n_903),
.Y(n_1039)
);

AOI22xp33_ASAP7_75t_L g1040 ( 
.A1(n_932),
.A2(n_652),
.B1(n_659),
.B2(n_646),
.Y(n_1040)
);

AOI22xp33_ASAP7_75t_L g1041 ( 
.A1(n_932),
.A2(n_668),
.B1(n_676),
.B2(n_665),
.Y(n_1041)
);

BUFx4f_ASAP7_75t_L g1042 ( 
.A(n_923),
.Y(n_1042)
);

INVx2_ASAP7_75t_L g1043 ( 
.A(n_941),
.Y(n_1043)
);

CKINVDCx20_ASAP7_75t_R g1044 ( 
.A(n_911),
.Y(n_1044)
);

INVx1_ASAP7_75t_L g1045 ( 
.A(n_947),
.Y(n_1045)
);

NAND2xp5_ASAP7_75t_L g1046 ( 
.A(n_947),
.B(n_827),
.Y(n_1046)
);

NOR2x1p5_ASAP7_75t_L g1047 ( 
.A(n_909),
.B(n_574),
.Y(n_1047)
);

AOI22xp33_ASAP7_75t_L g1048 ( 
.A1(n_917),
.A2(n_687),
.B1(n_691),
.B2(n_685),
.Y(n_1048)
);

AND3x2_ASAP7_75t_L g1049 ( 
.A(n_921),
.B(n_704),
.C(n_699),
.Y(n_1049)
);

INVxp67_ASAP7_75t_L g1050 ( 
.A(n_926),
.Y(n_1050)
);

NAND2xp5_ASAP7_75t_L g1051 ( 
.A(n_922),
.B(n_827),
.Y(n_1051)
);

NOR2xp33_ASAP7_75t_L g1052 ( 
.A(n_925),
.B(n_575),
.Y(n_1052)
);

OR2x6_ASAP7_75t_L g1053 ( 
.A(n_880),
.B(n_742),
.Y(n_1053)
);

AND2x2_ASAP7_75t_L g1054 ( 
.A(n_938),
.B(n_863),
.Y(n_1054)
);

INVx1_ASAP7_75t_L g1055 ( 
.A(n_881),
.Y(n_1055)
);

INVx5_ASAP7_75t_L g1056 ( 
.A(n_941),
.Y(n_1056)
);

INVx3_ASAP7_75t_L g1057 ( 
.A(n_941),
.Y(n_1057)
);

INVx2_ASAP7_75t_L g1058 ( 
.A(n_950),
.Y(n_1058)
);

INVxp67_ASAP7_75t_SL g1059 ( 
.A(n_950),
.Y(n_1059)
);

NOR2xp33_ASAP7_75t_L g1060 ( 
.A(n_884),
.B(n_592),
.Y(n_1060)
);

AND2x6_ASAP7_75t_L g1061 ( 
.A(n_887),
.B(n_569),
.Y(n_1061)
);

INVx1_ASAP7_75t_L g1062 ( 
.A(n_897),
.Y(n_1062)
);

AND2x4_ASAP7_75t_L g1063 ( 
.A(n_898),
.B(n_863),
.Y(n_1063)
);

BUFx10_ASAP7_75t_L g1064 ( 
.A(n_901),
.Y(n_1064)
);

INVx1_ASAP7_75t_L g1065 ( 
.A(n_908),
.Y(n_1065)
);

INVx2_ASAP7_75t_L g1066 ( 
.A(n_912),
.Y(n_1066)
);

AND2x6_ASAP7_75t_L g1067 ( 
.A(n_919),
.B(n_569),
.Y(n_1067)
);

INVx1_ASAP7_75t_L g1068 ( 
.A(n_924),
.Y(n_1068)
);

NAND2xp5_ASAP7_75t_L g1069 ( 
.A(n_929),
.B(n_832),
.Y(n_1069)
);

NOR2xp33_ASAP7_75t_L g1070 ( 
.A(n_979),
.B(n_683),
.Y(n_1070)
);

INVx2_ASAP7_75t_L g1071 ( 
.A(n_1063),
.Y(n_1071)
);

INVxp67_ASAP7_75t_L g1072 ( 
.A(n_968),
.Y(n_1072)
);

NAND2xp5_ASAP7_75t_L g1073 ( 
.A(n_1014),
.B(n_931),
.Y(n_1073)
);

NAND2xp5_ASAP7_75t_L g1074 ( 
.A(n_1018),
.B(n_706),
.Y(n_1074)
);

NOR2xp33_ASAP7_75t_L g1075 ( 
.A(n_960),
.B(n_587),
.Y(n_1075)
);

NAND2xp5_ASAP7_75t_L g1076 ( 
.A(n_1045),
.B(n_1013),
.Y(n_1076)
);

INVx1_ASAP7_75t_L g1077 ( 
.A(n_1054),
.Y(n_1077)
);

NAND2xp5_ASAP7_75t_L g1078 ( 
.A(n_1010),
.B(n_712),
.Y(n_1078)
);

NAND2xp5_ASAP7_75t_L g1079 ( 
.A(n_1012),
.B(n_714),
.Y(n_1079)
);

NAND2xp5_ASAP7_75t_L g1080 ( 
.A(n_1012),
.B(n_871),
.Y(n_1080)
);

INVx1_ASAP7_75t_L g1081 ( 
.A(n_959),
.Y(n_1081)
);

INVx1_ASAP7_75t_L g1082 ( 
.A(n_961),
.Y(n_1082)
);

NAND2xp5_ASAP7_75t_L g1083 ( 
.A(n_1004),
.B(n_871),
.Y(n_1083)
);

AOI22x1_ASAP7_75t_SL g1084 ( 
.A1(n_978),
.A2(n_593),
.B1(n_601),
.B2(n_591),
.Y(n_1084)
);

BUFx10_ASAP7_75t_L g1085 ( 
.A(n_1022),
.Y(n_1085)
);

NAND2xp33_ASAP7_75t_L g1086 ( 
.A(n_967),
.B(n_543),
.Y(n_1086)
);

INVx2_ASAP7_75t_L g1087 ( 
.A(n_1063),
.Y(n_1087)
);

NAND2xp5_ASAP7_75t_L g1088 ( 
.A(n_967),
.B(n_873),
.Y(n_1088)
);

NOR2xp33_ASAP7_75t_L g1089 ( 
.A(n_963),
.B(n_613),
.Y(n_1089)
);

NAND2xp5_ASAP7_75t_L g1090 ( 
.A(n_967),
.B(n_873),
.Y(n_1090)
);

NAND2xp5_ASAP7_75t_L g1091 ( 
.A(n_967),
.B(n_874),
.Y(n_1091)
);

INVx1_ASAP7_75t_L g1092 ( 
.A(n_965),
.Y(n_1092)
);

INVx2_ASAP7_75t_L g1093 ( 
.A(n_957),
.Y(n_1093)
);

INVx3_ASAP7_75t_L g1094 ( 
.A(n_1064),
.Y(n_1094)
);

INVx1_ASAP7_75t_L g1095 ( 
.A(n_969),
.Y(n_1095)
);

OR2x2_ASAP7_75t_L g1096 ( 
.A(n_986),
.B(n_874),
.Y(n_1096)
);

NAND2xp5_ASAP7_75t_SL g1097 ( 
.A(n_980),
.B(n_546),
.Y(n_1097)
);

HB1xp67_ASAP7_75t_L g1098 ( 
.A(n_964),
.Y(n_1098)
);

BUFx4_ASAP7_75t_L g1099 ( 
.A(n_1008),
.Y(n_1099)
);

BUFx6f_ASAP7_75t_L g1100 ( 
.A(n_1003),
.Y(n_1100)
);

INVx1_ASAP7_75t_L g1101 ( 
.A(n_972),
.Y(n_1101)
);

NAND2xp5_ASAP7_75t_L g1102 ( 
.A(n_1027),
.B(n_842),
.Y(n_1102)
);

NAND2xp5_ASAP7_75t_L g1103 ( 
.A(n_1036),
.B(n_842),
.Y(n_1103)
);

INVx2_ASAP7_75t_L g1104 ( 
.A(n_984),
.Y(n_1104)
);

INVx1_ASAP7_75t_L g1105 ( 
.A(n_995),
.Y(n_1105)
);

INVx1_ASAP7_75t_L g1106 ( 
.A(n_996),
.Y(n_1106)
);

NAND2xp5_ASAP7_75t_SL g1107 ( 
.A(n_962),
.B(n_555),
.Y(n_1107)
);

INVxp67_ASAP7_75t_L g1108 ( 
.A(n_989),
.Y(n_1108)
);

AND2x4_ASAP7_75t_SL g1109 ( 
.A(n_966),
.B(n_551),
.Y(n_1109)
);

NAND2xp5_ASAP7_75t_SL g1110 ( 
.A(n_1009),
.B(n_560),
.Y(n_1110)
);

NAND2xp5_ASAP7_75t_L g1111 ( 
.A(n_994),
.B(n_819),
.Y(n_1111)
);

NAND2xp5_ASAP7_75t_SL g1112 ( 
.A(n_1011),
.B(n_982),
.Y(n_1112)
);

NAND2xp5_ASAP7_75t_SL g1113 ( 
.A(n_973),
.B(n_1001),
.Y(n_1113)
);

NOR2xp33_ASAP7_75t_L g1114 ( 
.A(n_976),
.B(n_624),
.Y(n_1114)
);

INVx2_ASAP7_75t_SL g1115 ( 
.A(n_981),
.Y(n_1115)
);

NAND2xp5_ASAP7_75t_L g1116 ( 
.A(n_1052),
.B(n_830),
.Y(n_1116)
);

NAND2xp5_ASAP7_75t_L g1117 ( 
.A(n_1040),
.B(n_834),
.Y(n_1117)
);

NOR2xp33_ASAP7_75t_L g1118 ( 
.A(n_1002),
.B(n_627),
.Y(n_1118)
);

INVxp67_ASAP7_75t_L g1119 ( 
.A(n_1000),
.Y(n_1119)
);

BUFx6f_ASAP7_75t_SL g1120 ( 
.A(n_1020),
.Y(n_1120)
);

NAND2xp5_ASAP7_75t_L g1121 ( 
.A(n_1041),
.B(n_832),
.Y(n_1121)
);

AOI22xp5_ASAP7_75t_L g1122 ( 
.A1(n_1033),
.A2(n_970),
.B1(n_974),
.B2(n_983),
.Y(n_1122)
);

CKINVDCx5p33_ASAP7_75t_R g1123 ( 
.A(n_977),
.Y(n_1123)
);

INVx4_ASAP7_75t_L g1124 ( 
.A(n_1003),
.Y(n_1124)
);

NAND2xp5_ASAP7_75t_SL g1125 ( 
.A(n_975),
.B(n_1015),
.Y(n_1125)
);

OAI22xp5_ASAP7_75t_L g1126 ( 
.A1(n_1021),
.A2(n_563),
.B1(n_567),
.B2(n_561),
.Y(n_1126)
);

NAND3x1_ASAP7_75t_L g1127 ( 
.A(n_1035),
.B(n_744),
.C(n_743),
.Y(n_1127)
);

NOR2xp33_ASAP7_75t_L g1128 ( 
.A(n_987),
.B(n_628),
.Y(n_1128)
);

INVx2_ASAP7_75t_L g1129 ( 
.A(n_997),
.Y(n_1129)
);

NAND2xp5_ASAP7_75t_L g1130 ( 
.A(n_1060),
.B(n_833),
.Y(n_1130)
);

AND2x2_ASAP7_75t_L g1131 ( 
.A(n_966),
.B(n_562),
.Y(n_1131)
);

BUFx6f_ASAP7_75t_L g1132 ( 
.A(n_1064),
.Y(n_1132)
);

NAND2xp5_ASAP7_75t_SL g1133 ( 
.A(n_975),
.B(n_579),
.Y(n_1133)
);

NOR2xp33_ASAP7_75t_SL g1134 ( 
.A(n_1008),
.B(n_617),
.Y(n_1134)
);

AO22x1_ASAP7_75t_L g1135 ( 
.A1(n_985),
.A2(n_638),
.B1(n_644),
.B2(n_630),
.Y(n_1135)
);

NAND2xp5_ASAP7_75t_L g1136 ( 
.A(n_1046),
.B(n_583),
.Y(n_1136)
);

NAND3xp33_ASAP7_75t_L g1137 ( 
.A(n_993),
.B(n_654),
.C(n_648),
.Y(n_1137)
);

OAI221xp5_ASAP7_75t_L g1138 ( 
.A1(n_1037),
.A2(n_1038),
.B1(n_1048),
.B2(n_990),
.C(n_1017),
.Y(n_1138)
);

NAND2xp5_ASAP7_75t_L g1139 ( 
.A(n_1024),
.B(n_588),
.Y(n_1139)
);

NAND2xp5_ASAP7_75t_L g1140 ( 
.A(n_1024),
.B(n_589),
.Y(n_1140)
);

NAND2xp5_ASAP7_75t_SL g1141 ( 
.A(n_975),
.B(n_1015),
.Y(n_1141)
);

NAND2xp5_ASAP7_75t_L g1142 ( 
.A(n_1024),
.B(n_598),
.Y(n_1142)
);

O2A1O1Ixp33_ASAP7_75t_L g1143 ( 
.A1(n_1050),
.A2(n_746),
.B(n_747),
.C(n_745),
.Y(n_1143)
);

BUFx3_ASAP7_75t_L g1144 ( 
.A(n_1028),
.Y(n_1144)
);

OAI21xp5_ASAP7_75t_L g1145 ( 
.A1(n_1042),
.A2(n_877),
.B(n_609),
.Y(n_1145)
);

INVx1_ASAP7_75t_L g1146 ( 
.A(n_991),
.Y(n_1146)
);

NAND2xp5_ASAP7_75t_L g1147 ( 
.A(n_1024),
.B(n_600),
.Y(n_1147)
);

INVx1_ASAP7_75t_L g1148 ( 
.A(n_992),
.Y(n_1148)
);

AND2x4_ASAP7_75t_SL g1149 ( 
.A(n_958),
.B(n_617),
.Y(n_1149)
);

NAND2xp33_ASAP7_75t_L g1150 ( 
.A(n_1015),
.B(n_610),
.Y(n_1150)
);

INVxp67_ASAP7_75t_L g1151 ( 
.A(n_1025),
.Y(n_1151)
);

NAND2xp5_ASAP7_75t_L g1152 ( 
.A(n_1026),
.B(n_615),
.Y(n_1152)
);

NOR2xp33_ASAP7_75t_L g1153 ( 
.A(n_1044),
.B(n_669),
.Y(n_1153)
);

NAND2xp5_ASAP7_75t_L g1154 ( 
.A(n_1026),
.B(n_618),
.Y(n_1154)
);

NOR2x1p5_ASAP7_75t_L g1155 ( 
.A(n_958),
.B(n_674),
.Y(n_1155)
);

NOR2xp33_ASAP7_75t_L g1156 ( 
.A(n_990),
.B(n_675),
.Y(n_1156)
);

BUFx6f_ASAP7_75t_L g1157 ( 
.A(n_1053),
.Y(n_1157)
);

NOR2xp33_ASAP7_75t_L g1158 ( 
.A(n_1053),
.B(n_682),
.Y(n_1158)
);

BUFx6f_ASAP7_75t_L g1159 ( 
.A(n_999),
.Y(n_1159)
);

NAND2xp5_ASAP7_75t_SL g1160 ( 
.A(n_1030),
.B(n_625),
.Y(n_1160)
);

NAND2xp5_ASAP7_75t_L g1161 ( 
.A(n_1026),
.B(n_1059),
.Y(n_1161)
);

NOR2xp33_ASAP7_75t_SL g1162 ( 
.A(n_1032),
.B(n_617),
.Y(n_1162)
);

AOI22xp33_ASAP7_75t_L g1163 ( 
.A1(n_988),
.A2(n_660),
.B1(n_621),
.B2(n_877),
.Y(n_1163)
);

INVxp67_ASAP7_75t_SL g1164 ( 
.A(n_1031),
.Y(n_1164)
);

NAND2xp5_ASAP7_75t_L g1165 ( 
.A(n_1055),
.B(n_1062),
.Y(n_1165)
);

NOR2xp33_ASAP7_75t_L g1166 ( 
.A(n_1032),
.B(n_686),
.Y(n_1166)
);

NAND2xp5_ASAP7_75t_L g1167 ( 
.A(n_1065),
.B(n_629),
.Y(n_1167)
);

INVxp67_ASAP7_75t_L g1168 ( 
.A(n_1047),
.Y(n_1168)
);

NAND2xp5_ASAP7_75t_L g1169 ( 
.A(n_1068),
.B(n_634),
.Y(n_1169)
);

NAND2xp5_ASAP7_75t_L g1170 ( 
.A(n_1066),
.B(n_635),
.Y(n_1170)
);

NAND2xp5_ASAP7_75t_L g1171 ( 
.A(n_998),
.B(n_639),
.Y(n_1171)
);

NAND2xp33_ASAP7_75t_L g1172 ( 
.A(n_1030),
.B(n_645),
.Y(n_1172)
);

NAND2xp5_ASAP7_75t_SL g1173 ( 
.A(n_1056),
.B(n_657),
.Y(n_1173)
);

INVx2_ASAP7_75t_L g1174 ( 
.A(n_1005),
.Y(n_1174)
);

NAND2xp5_ASAP7_75t_L g1175 ( 
.A(n_1007),
.B(n_1016),
.Y(n_1175)
);

NAND2xp5_ASAP7_75t_L g1176 ( 
.A(n_1043),
.B(n_661),
.Y(n_1176)
);

AOI21xp5_ASAP7_75t_L g1177 ( 
.A1(n_1056),
.A2(n_841),
.B(n_838),
.Y(n_1177)
);

AOI22xp33_ASAP7_75t_L g1178 ( 
.A1(n_1051),
.A2(n_660),
.B1(n_621),
.B2(n_666),
.Y(n_1178)
);

OR2x6_ASAP7_75t_L g1179 ( 
.A(n_1006),
.B(n_748),
.Y(n_1179)
);

NAND2xp5_ASAP7_75t_L g1180 ( 
.A(n_1058),
.B(n_670),
.Y(n_1180)
);

INVx1_ASAP7_75t_L g1181 ( 
.A(n_1069),
.Y(n_1181)
);

NAND2xp5_ASAP7_75t_SL g1182 ( 
.A(n_1056),
.B(n_672),
.Y(n_1182)
);

OAI22xp5_ASAP7_75t_L g1183 ( 
.A1(n_1057),
.A2(n_679),
.B1(n_680),
.B2(n_678),
.Y(n_1183)
);

BUFx6f_ASAP7_75t_L g1184 ( 
.A(n_1019),
.Y(n_1184)
);

AND2x2_ASAP7_75t_L g1185 ( 
.A(n_1006),
.B(n_692),
.Y(n_1185)
);

AOI22xp33_ASAP7_75t_L g1186 ( 
.A1(n_1023),
.A2(n_660),
.B1(n_621),
.B2(n_698),
.Y(n_1186)
);

O2A1O1Ixp33_ASAP7_75t_L g1187 ( 
.A1(n_1049),
.A2(n_753),
.B(n_759),
.C(n_750),
.Y(n_1187)
);

INVx2_ASAP7_75t_L g1188 ( 
.A(n_1029),
.Y(n_1188)
);

NAND2xp33_ASAP7_75t_L g1189 ( 
.A(n_1061),
.B(n_703),
.Y(n_1189)
);

INVx1_ASAP7_75t_L g1190 ( 
.A(n_1029),
.Y(n_1190)
);

BUFx6f_ASAP7_75t_L g1191 ( 
.A(n_1034),
.Y(n_1191)
);

HB1xp67_ASAP7_75t_L g1192 ( 
.A(n_971),
.Y(n_1192)
);

NAND2xp5_ASAP7_75t_SL g1193 ( 
.A(n_1034),
.B(n_707),
.Y(n_1193)
);

INVxp67_ASAP7_75t_L g1194 ( 
.A(n_1061),
.Y(n_1194)
);

NAND2xp5_ASAP7_75t_L g1195 ( 
.A(n_1039),
.B(n_710),
.Y(n_1195)
);

NAND2xp5_ASAP7_75t_L g1196 ( 
.A(n_1039),
.B(n_971),
.Y(n_1196)
);

INVx1_ASAP7_75t_L g1197 ( 
.A(n_1061),
.Y(n_1197)
);

OAI22xp5_ASAP7_75t_L g1198 ( 
.A1(n_1061),
.A2(n_717),
.B1(n_718),
.B2(n_711),
.Y(n_1198)
);

INVx1_ASAP7_75t_L g1199 ( 
.A(n_1067),
.Y(n_1199)
);

NOR2xp33_ASAP7_75t_L g1200 ( 
.A(n_1067),
.B(n_696),
.Y(n_1200)
);

AOI21xp5_ASAP7_75t_L g1201 ( 
.A1(n_1067),
.A2(n_841),
.B(n_838),
.Y(n_1201)
);

AOI22xp5_ASAP7_75t_L g1202 ( 
.A1(n_1014),
.A2(n_763),
.B1(n_766),
.B2(n_762),
.Y(n_1202)
);

NAND2xp5_ASAP7_75t_SL g1203 ( 
.A(n_980),
.B(n_838),
.Y(n_1203)
);

AOI22xp33_ASAP7_75t_SL g1204 ( 
.A1(n_989),
.A2(n_692),
.B1(n_709),
.B2(n_705),
.Y(n_1204)
);

NAND2xp5_ASAP7_75t_L g1205 ( 
.A(n_1014),
.B(n_841),
.Y(n_1205)
);

AOI22xp33_ASAP7_75t_L g1206 ( 
.A1(n_967),
.A2(n_767),
.B1(n_776),
.B2(n_769),
.Y(n_1206)
);

NOR2xp33_ASAP7_75t_L g1207 ( 
.A(n_979),
.B(n_692),
.Y(n_1207)
);

NAND2xp5_ASAP7_75t_L g1208 ( 
.A(n_1014),
.B(n_841),
.Y(n_1208)
);

NOR2xp33_ASAP7_75t_L g1209 ( 
.A(n_979),
.B(n_777),
.Y(n_1209)
);

HB1xp67_ASAP7_75t_L g1210 ( 
.A(n_986),
.Y(n_1210)
);

INVx1_ASAP7_75t_L g1211 ( 
.A(n_1054),
.Y(n_1211)
);

INVx3_ASAP7_75t_L g1212 ( 
.A(n_1064),
.Y(n_1212)
);

AND2x2_ASAP7_75t_L g1213 ( 
.A(n_980),
.B(n_778),
.Y(n_1213)
);

INVx1_ASAP7_75t_L g1214 ( 
.A(n_1054),
.Y(n_1214)
);

NAND2xp5_ASAP7_75t_L g1215 ( 
.A(n_1014),
.B(n_779),
.Y(n_1215)
);

NAND2xp5_ASAP7_75t_L g1216 ( 
.A(n_1014),
.B(n_0),
.Y(n_1216)
);

INVx1_ASAP7_75t_L g1217 ( 
.A(n_1054),
.Y(n_1217)
);

NOR2xp67_ASAP7_75t_SL g1218 ( 
.A(n_975),
.B(n_1),
.Y(n_1218)
);

AOI22xp5_ASAP7_75t_L g1219 ( 
.A1(n_1045),
.A2(n_229),
.B1(n_232),
.B2(n_228),
.Y(n_1219)
);

NAND2xp5_ASAP7_75t_L g1220 ( 
.A(n_1014),
.B(n_2),
.Y(n_1220)
);

INVx2_ASAP7_75t_L g1221 ( 
.A(n_1063),
.Y(n_1221)
);

INVx3_ASAP7_75t_L g1222 ( 
.A(n_1064),
.Y(n_1222)
);

AOI21xp5_ASAP7_75t_L g1223 ( 
.A1(n_983),
.A2(n_237),
.B(n_236),
.Y(n_1223)
);

NAND2xp5_ASAP7_75t_L g1224 ( 
.A(n_1014),
.B(n_2),
.Y(n_1224)
);

NAND2xp5_ASAP7_75t_L g1225 ( 
.A(n_1014),
.B(n_3),
.Y(n_1225)
);

BUFx6f_ASAP7_75t_L g1226 ( 
.A(n_1003),
.Y(n_1226)
);

INVx1_ASAP7_75t_L g1227 ( 
.A(n_1054),
.Y(n_1227)
);

INVx1_ASAP7_75t_L g1228 ( 
.A(n_1054),
.Y(n_1228)
);

OR2x2_ASAP7_75t_L g1229 ( 
.A(n_968),
.B(n_6),
.Y(n_1229)
);

NAND2xp5_ASAP7_75t_L g1230 ( 
.A(n_1014),
.B(n_7),
.Y(n_1230)
);

OR2x2_ASAP7_75t_L g1231 ( 
.A(n_968),
.B(n_7),
.Y(n_1231)
);

NAND2xp5_ASAP7_75t_L g1232 ( 
.A(n_1076),
.B(n_8),
.Y(n_1232)
);

BUFx12f_ASAP7_75t_SL g1233 ( 
.A(n_1179),
.Y(n_1233)
);

AND2x6_ASAP7_75t_L g1234 ( 
.A(n_1122),
.B(n_240),
.Y(n_1234)
);

INVx1_ASAP7_75t_L g1235 ( 
.A(n_1081),
.Y(n_1235)
);

INVx2_ASAP7_75t_SL g1236 ( 
.A(n_1098),
.Y(n_1236)
);

INVx1_ASAP7_75t_L g1237 ( 
.A(n_1082),
.Y(n_1237)
);

AND2x6_ASAP7_75t_L g1238 ( 
.A(n_1122),
.B(n_242),
.Y(n_1238)
);

NOR3xp33_ASAP7_75t_SL g1239 ( 
.A(n_1138),
.B(n_9),
.C(n_11),
.Y(n_1239)
);

AOI22xp5_ASAP7_75t_L g1240 ( 
.A1(n_1075),
.A2(n_244),
.B1(n_245),
.B2(n_243),
.Y(n_1240)
);

BUFx3_ASAP7_75t_L g1241 ( 
.A(n_1144),
.Y(n_1241)
);

NAND2xp5_ASAP7_75t_L g1242 ( 
.A(n_1089),
.B(n_9),
.Y(n_1242)
);

AND2x2_ASAP7_75t_L g1243 ( 
.A(n_1210),
.B(n_11),
.Y(n_1243)
);

INVx2_ASAP7_75t_L g1244 ( 
.A(n_1071),
.Y(n_1244)
);

INVx2_ASAP7_75t_L g1245 ( 
.A(n_1087),
.Y(n_1245)
);

BUFx3_ASAP7_75t_L g1246 ( 
.A(n_1132),
.Y(n_1246)
);

INVx2_ASAP7_75t_L g1247 ( 
.A(n_1221),
.Y(n_1247)
);

CKINVDCx8_ASAP7_75t_R g1248 ( 
.A(n_1123),
.Y(n_1248)
);

INVx2_ASAP7_75t_SL g1249 ( 
.A(n_1157),
.Y(n_1249)
);

AND2x6_ASAP7_75t_L g1250 ( 
.A(n_1219),
.B(n_252),
.Y(n_1250)
);

NAND2x1p5_ASAP7_75t_L g1251 ( 
.A(n_1094),
.B(n_254),
.Y(n_1251)
);

AND2x2_ASAP7_75t_L g1252 ( 
.A(n_1213),
.B(n_12),
.Y(n_1252)
);

NAND2xp5_ASAP7_75t_L g1253 ( 
.A(n_1077),
.B(n_13),
.Y(n_1253)
);

AND2x4_ASAP7_75t_L g1254 ( 
.A(n_1168),
.B(n_1129),
.Y(n_1254)
);

NOR2x1p5_ASAP7_75t_L g1255 ( 
.A(n_1094),
.B(n_255),
.Y(n_1255)
);

BUFx6f_ASAP7_75t_L g1256 ( 
.A(n_1100),
.Y(n_1256)
);

INVx1_ASAP7_75t_L g1257 ( 
.A(n_1092),
.Y(n_1257)
);

AND2x6_ASAP7_75t_SL g1258 ( 
.A(n_1153),
.B(n_13),
.Y(n_1258)
);

AND2x6_ASAP7_75t_SL g1259 ( 
.A(n_1179),
.B(n_14),
.Y(n_1259)
);

OR2x4_ASAP7_75t_L g1260 ( 
.A(n_1156),
.B(n_15),
.Y(n_1260)
);

INVx2_ASAP7_75t_L g1261 ( 
.A(n_1104),
.Y(n_1261)
);

AOI21x1_ASAP7_75t_L g1262 ( 
.A1(n_1088),
.A2(n_258),
.B(n_256),
.Y(n_1262)
);

INVx2_ASAP7_75t_SL g1263 ( 
.A(n_1157),
.Y(n_1263)
);

NAND2xp5_ASAP7_75t_L g1264 ( 
.A(n_1211),
.B(n_15),
.Y(n_1264)
);

BUFx3_ASAP7_75t_L g1265 ( 
.A(n_1115),
.Y(n_1265)
);

AND2x2_ASAP7_75t_L g1266 ( 
.A(n_1072),
.B(n_16),
.Y(n_1266)
);

AND2x6_ASAP7_75t_L g1267 ( 
.A(n_1219),
.B(n_259),
.Y(n_1267)
);

NAND2xp5_ASAP7_75t_L g1268 ( 
.A(n_1214),
.B(n_18),
.Y(n_1268)
);

AND2x2_ASAP7_75t_L g1269 ( 
.A(n_1118),
.B(n_18),
.Y(n_1269)
);

AOI22xp5_ASAP7_75t_L g1270 ( 
.A1(n_1114),
.A2(n_261),
.B1(n_262),
.B2(n_260),
.Y(n_1270)
);

HB1xp67_ASAP7_75t_L g1271 ( 
.A(n_1119),
.Y(n_1271)
);

INVx2_ASAP7_75t_SL g1272 ( 
.A(n_1157),
.Y(n_1272)
);

AND2x2_ASAP7_75t_L g1273 ( 
.A(n_1209),
.B(n_19),
.Y(n_1273)
);

NAND3xp33_ASAP7_75t_SL g1274 ( 
.A(n_1204),
.B(n_19),
.C(n_20),
.Y(n_1274)
);

AND2x4_ASAP7_75t_L g1275 ( 
.A(n_1212),
.B(n_267),
.Y(n_1275)
);

INVx2_ASAP7_75t_L g1276 ( 
.A(n_1101),
.Y(n_1276)
);

NAND2xp5_ASAP7_75t_L g1277 ( 
.A(n_1217),
.B(n_1227),
.Y(n_1277)
);

AOI21xp5_ASAP7_75t_L g1278 ( 
.A1(n_1113),
.A2(n_1145),
.B(n_1161),
.Y(n_1278)
);

INVxp67_ASAP7_75t_SL g1279 ( 
.A(n_1184),
.Y(n_1279)
);

AND2x4_ASAP7_75t_L g1280 ( 
.A(n_1212),
.B(n_269),
.Y(n_1280)
);

NAND2xp5_ASAP7_75t_L g1281 ( 
.A(n_1228),
.B(n_21),
.Y(n_1281)
);

NAND2xp5_ASAP7_75t_L g1282 ( 
.A(n_1083),
.B(n_22),
.Y(n_1282)
);

NAND2xp5_ASAP7_75t_SL g1283 ( 
.A(n_1222),
.B(n_270),
.Y(n_1283)
);

NAND2xp5_ASAP7_75t_SL g1284 ( 
.A(n_1222),
.B(n_271),
.Y(n_1284)
);

AOI22xp33_ASAP7_75t_L g1285 ( 
.A1(n_1112),
.A2(n_25),
.B1(n_22),
.B2(n_23),
.Y(n_1285)
);

INVx1_ASAP7_75t_L g1286 ( 
.A(n_1095),
.Y(n_1286)
);

INVx3_ASAP7_75t_L g1287 ( 
.A(n_1100),
.Y(n_1287)
);

INVx2_ASAP7_75t_L g1288 ( 
.A(n_1093),
.Y(n_1288)
);

NAND2xp5_ASAP7_75t_SL g1289 ( 
.A(n_1184),
.B(n_272),
.Y(n_1289)
);

NAND2xp5_ASAP7_75t_L g1290 ( 
.A(n_1215),
.B(n_1116),
.Y(n_1290)
);

INVx1_ASAP7_75t_L g1291 ( 
.A(n_1105),
.Y(n_1291)
);

NAND2xp5_ASAP7_75t_L g1292 ( 
.A(n_1080),
.B(n_23),
.Y(n_1292)
);

INVx1_ASAP7_75t_L g1293 ( 
.A(n_1106),
.Y(n_1293)
);

INVx5_ASAP7_75t_L g1294 ( 
.A(n_1184),
.Y(n_1294)
);

NAND2xp5_ASAP7_75t_L g1295 ( 
.A(n_1216),
.B(n_25),
.Y(n_1295)
);

NAND2xp5_ASAP7_75t_SL g1296 ( 
.A(n_1191),
.B(n_275),
.Y(n_1296)
);

INVx1_ASAP7_75t_L g1297 ( 
.A(n_1102),
.Y(n_1297)
);

BUFx6f_ASAP7_75t_L g1298 ( 
.A(n_1100),
.Y(n_1298)
);

NAND2xp5_ASAP7_75t_L g1299 ( 
.A(n_1220),
.B(n_26),
.Y(n_1299)
);

NAND2xp5_ASAP7_75t_L g1300 ( 
.A(n_1224),
.B(n_26),
.Y(n_1300)
);

INVx1_ASAP7_75t_L g1301 ( 
.A(n_1103),
.Y(n_1301)
);

INVxp67_ASAP7_75t_SL g1302 ( 
.A(n_1191),
.Y(n_1302)
);

BUFx6f_ASAP7_75t_L g1303 ( 
.A(n_1226),
.Y(n_1303)
);

INVx2_ASAP7_75t_SL g1304 ( 
.A(n_1096),
.Y(n_1304)
);

AOI22xp5_ASAP7_75t_L g1305 ( 
.A1(n_1070),
.A2(n_278),
.B1(n_280),
.B2(n_276),
.Y(n_1305)
);

INVx2_ASAP7_75t_L g1306 ( 
.A(n_1146),
.Y(n_1306)
);

INVx2_ASAP7_75t_L g1307 ( 
.A(n_1148),
.Y(n_1307)
);

INVx1_ASAP7_75t_L g1308 ( 
.A(n_1165),
.Y(n_1308)
);

BUFx2_ASAP7_75t_L g1309 ( 
.A(n_1151),
.Y(n_1309)
);

BUFx2_ASAP7_75t_L g1310 ( 
.A(n_1179),
.Y(n_1310)
);

INVx2_ASAP7_75t_SL g1311 ( 
.A(n_1229),
.Y(n_1311)
);

NAND2xp5_ASAP7_75t_L g1312 ( 
.A(n_1225),
.B(n_27),
.Y(n_1312)
);

NAND2xp5_ASAP7_75t_L g1313 ( 
.A(n_1230),
.B(n_28),
.Y(n_1313)
);

NOR2xp33_ASAP7_75t_L g1314 ( 
.A(n_1108),
.B(n_28),
.Y(n_1314)
);

BUFx3_ASAP7_75t_L g1315 ( 
.A(n_1185),
.Y(n_1315)
);

AOI22xp33_ASAP7_75t_L g1316 ( 
.A1(n_1206),
.A2(n_31),
.B1(n_29),
.B2(n_30),
.Y(n_1316)
);

INVx1_ASAP7_75t_L g1317 ( 
.A(n_1073),
.Y(n_1317)
);

AOI22xp5_ASAP7_75t_L g1318 ( 
.A1(n_1107),
.A2(n_284),
.B1(n_286),
.B2(n_283),
.Y(n_1318)
);

AND2x6_ASAP7_75t_L g1319 ( 
.A(n_1196),
.B(n_287),
.Y(n_1319)
);

INVx1_ASAP7_75t_L g1320 ( 
.A(n_1175),
.Y(n_1320)
);

NAND2xp5_ASAP7_75t_SL g1321 ( 
.A(n_1191),
.B(n_288),
.Y(n_1321)
);

NAND2xp5_ASAP7_75t_L g1322 ( 
.A(n_1074),
.B(n_29),
.Y(n_1322)
);

NAND2xp5_ASAP7_75t_SL g1323 ( 
.A(n_1085),
.B(n_289),
.Y(n_1323)
);

INVx1_ASAP7_75t_L g1324 ( 
.A(n_1174),
.Y(n_1324)
);

AND2x2_ASAP7_75t_L g1325 ( 
.A(n_1207),
.B(n_30),
.Y(n_1325)
);

INVx5_ASAP7_75t_L g1326 ( 
.A(n_1226),
.Y(n_1326)
);

BUFx2_ASAP7_75t_L g1327 ( 
.A(n_1131),
.Y(n_1327)
);

INVxp67_ASAP7_75t_L g1328 ( 
.A(n_1231),
.Y(n_1328)
);

NAND2xp5_ASAP7_75t_L g1329 ( 
.A(n_1181),
.B(n_31),
.Y(n_1329)
);

BUFx2_ASAP7_75t_L g1330 ( 
.A(n_1127),
.Y(n_1330)
);

INVx1_ASAP7_75t_L g1331 ( 
.A(n_1205),
.Y(n_1331)
);

INVx1_ASAP7_75t_L g1332 ( 
.A(n_1208),
.Y(n_1332)
);

AND2x2_ASAP7_75t_L g1333 ( 
.A(n_1085),
.B(n_1128),
.Y(n_1333)
);

NAND2xp5_ASAP7_75t_L g1334 ( 
.A(n_1136),
.B(n_32),
.Y(n_1334)
);

AND2x4_ASAP7_75t_L g1335 ( 
.A(n_1155),
.B(n_290),
.Y(n_1335)
);

AND2x4_ASAP7_75t_L g1336 ( 
.A(n_1192),
.B(n_291),
.Y(n_1336)
);

BUFx2_ASAP7_75t_L g1337 ( 
.A(n_1226),
.Y(n_1337)
);

AND2x4_ASAP7_75t_L g1338 ( 
.A(n_1137),
.B(n_292),
.Y(n_1338)
);

AND2x2_ASAP7_75t_L g1339 ( 
.A(n_1158),
.B(n_33),
.Y(n_1339)
);

AOI21x1_ASAP7_75t_L g1340 ( 
.A1(n_1090),
.A2(n_295),
.B(n_294),
.Y(n_1340)
);

AND2x4_ASAP7_75t_L g1341 ( 
.A(n_1188),
.B(n_296),
.Y(n_1341)
);

INVx2_ASAP7_75t_L g1342 ( 
.A(n_1159),
.Y(n_1342)
);

BUFx6f_ASAP7_75t_L g1343 ( 
.A(n_1124),
.Y(n_1343)
);

BUFx3_ASAP7_75t_L g1344 ( 
.A(n_1166),
.Y(n_1344)
);

INVx6_ASAP7_75t_L g1345 ( 
.A(n_1159),
.Y(n_1345)
);

NOR2xp33_ASAP7_75t_L g1346 ( 
.A(n_1097),
.B(n_34),
.Y(n_1346)
);

AOI22xp5_ASAP7_75t_L g1347 ( 
.A1(n_1110),
.A2(n_302),
.B1(n_303),
.B2(n_300),
.Y(n_1347)
);

BUFx2_ASAP7_75t_L g1348 ( 
.A(n_1159),
.Y(n_1348)
);

NAND2xp5_ASAP7_75t_L g1349 ( 
.A(n_1079),
.B(n_34),
.Y(n_1349)
);

INVx2_ASAP7_75t_L g1350 ( 
.A(n_1190),
.Y(n_1350)
);

HB1xp67_ASAP7_75t_L g1351 ( 
.A(n_1203),
.Y(n_1351)
);

AND2x2_ASAP7_75t_L g1352 ( 
.A(n_1109),
.B(n_35),
.Y(n_1352)
);

AND2x6_ASAP7_75t_L g1353 ( 
.A(n_1091),
.B(n_304),
.Y(n_1353)
);

NAND2x1p5_ASAP7_75t_L g1354 ( 
.A(n_1125),
.B(n_306),
.Y(n_1354)
);

INVx1_ASAP7_75t_L g1355 ( 
.A(n_1143),
.Y(n_1355)
);

INVx2_ASAP7_75t_L g1356 ( 
.A(n_1121),
.Y(n_1356)
);

INVx1_ASAP7_75t_L g1357 ( 
.A(n_1164),
.Y(n_1357)
);

NAND2xp5_ASAP7_75t_L g1358 ( 
.A(n_1078),
.B(n_35),
.Y(n_1358)
);

CKINVDCx6p67_ASAP7_75t_R g1359 ( 
.A(n_1120),
.Y(n_1359)
);

CKINVDCx14_ASAP7_75t_R g1360 ( 
.A(n_1099),
.Y(n_1360)
);

CKINVDCx20_ASAP7_75t_R g1361 ( 
.A(n_1084),
.Y(n_1361)
);

INVx1_ASAP7_75t_L g1362 ( 
.A(n_1202),
.Y(n_1362)
);

INVx1_ASAP7_75t_L g1363 ( 
.A(n_1111),
.Y(n_1363)
);

NAND2x1p5_ASAP7_75t_L g1364 ( 
.A(n_1141),
.B(n_308),
.Y(n_1364)
);

INVx2_ASAP7_75t_L g1365 ( 
.A(n_1130),
.Y(n_1365)
);

AOI22xp33_ASAP7_75t_L g1366 ( 
.A1(n_1186),
.A2(n_39),
.B1(n_37),
.B2(n_38),
.Y(n_1366)
);

OR2x2_ASAP7_75t_L g1367 ( 
.A(n_1135),
.B(n_1176),
.Y(n_1367)
);

INVx2_ASAP7_75t_L g1368 ( 
.A(n_1117),
.Y(n_1368)
);

INVx2_ASAP7_75t_SL g1369 ( 
.A(n_1149),
.Y(n_1369)
);

BUFx6f_ASAP7_75t_L g1370 ( 
.A(n_1133),
.Y(n_1370)
);

NAND2xp5_ASAP7_75t_L g1371 ( 
.A(n_1195),
.B(n_40),
.Y(n_1371)
);

INVx1_ASAP7_75t_L g1372 ( 
.A(n_1180),
.Y(n_1372)
);

AND2x4_ASAP7_75t_L g1373 ( 
.A(n_1173),
.B(n_309),
.Y(n_1373)
);

INVx5_ASAP7_75t_L g1374 ( 
.A(n_1218),
.Y(n_1374)
);

AND2x2_ASAP7_75t_L g1375 ( 
.A(n_1162),
.B(n_41),
.Y(n_1375)
);

NAND2xp5_ASAP7_75t_L g1376 ( 
.A(n_1126),
.B(n_41),
.Y(n_1376)
);

NAND2xp5_ASAP7_75t_L g1377 ( 
.A(n_1163),
.B(n_42),
.Y(n_1377)
);

AND2x4_ASAP7_75t_L g1378 ( 
.A(n_1182),
.B(n_310),
.Y(n_1378)
);

NAND2xp5_ASAP7_75t_L g1379 ( 
.A(n_1167),
.B(n_42),
.Y(n_1379)
);

HB1xp67_ASAP7_75t_L g1380 ( 
.A(n_1169),
.Y(n_1380)
);

NOR2xp33_ASAP7_75t_R g1381 ( 
.A(n_1086),
.B(n_1150),
.Y(n_1381)
);

INVx1_ASAP7_75t_L g1382 ( 
.A(n_1170),
.Y(n_1382)
);

OR2x6_ASAP7_75t_L g1383 ( 
.A(n_1223),
.B(n_45),
.Y(n_1383)
);

INVx1_ASAP7_75t_L g1384 ( 
.A(n_1171),
.Y(n_1384)
);

HB1xp67_ASAP7_75t_L g1385 ( 
.A(n_1193),
.Y(n_1385)
);

BUFx6f_ASAP7_75t_L g1386 ( 
.A(n_1160),
.Y(n_1386)
);

BUFx6f_ASAP7_75t_L g1387 ( 
.A(n_1197),
.Y(n_1387)
);

INVx1_ASAP7_75t_L g1388 ( 
.A(n_1199),
.Y(n_1388)
);

INVx1_ASAP7_75t_L g1389 ( 
.A(n_1187),
.Y(n_1389)
);

INVx1_ASAP7_75t_L g1390 ( 
.A(n_1194),
.Y(n_1390)
);

CKINVDCx5p33_ASAP7_75t_R g1391 ( 
.A(n_1183),
.Y(n_1391)
);

NAND2xp5_ASAP7_75t_SL g1392 ( 
.A(n_1178),
.B(n_1139),
.Y(n_1392)
);

INVx1_ASAP7_75t_L g1393 ( 
.A(n_1140),
.Y(n_1393)
);

NOR2xp33_ASAP7_75t_L g1394 ( 
.A(n_1134),
.B(n_46),
.Y(n_1394)
);

NAND2xp5_ASAP7_75t_L g1395 ( 
.A(n_1200),
.B(n_46),
.Y(n_1395)
);

BUFx6f_ASAP7_75t_L g1396 ( 
.A(n_1142),
.Y(n_1396)
);

NOR3xp33_ASAP7_75t_SL g1397 ( 
.A(n_1198),
.B(n_48),
.C(n_49),
.Y(n_1397)
);

INVx2_ASAP7_75t_SL g1398 ( 
.A(n_1147),
.Y(n_1398)
);

AND2x2_ASAP7_75t_L g1399 ( 
.A(n_1152),
.B(n_49),
.Y(n_1399)
);

INVx1_ASAP7_75t_L g1400 ( 
.A(n_1154),
.Y(n_1400)
);

BUFx6f_ASAP7_75t_L g1401 ( 
.A(n_1256),
.Y(n_1401)
);

NAND2xp5_ASAP7_75t_L g1402 ( 
.A(n_1290),
.B(n_1172),
.Y(n_1402)
);

INVx1_ASAP7_75t_L g1403 ( 
.A(n_1235),
.Y(n_1403)
);

INVx3_ASAP7_75t_L g1404 ( 
.A(n_1294),
.Y(n_1404)
);

BUFx8_ASAP7_75t_L g1405 ( 
.A(n_1310),
.Y(n_1405)
);

AND2x6_ASAP7_75t_L g1406 ( 
.A(n_1341),
.B(n_312),
.Y(n_1406)
);

NOR2xp33_ASAP7_75t_L g1407 ( 
.A(n_1344),
.B(n_1189),
.Y(n_1407)
);

HB1xp67_ASAP7_75t_L g1408 ( 
.A(n_1271),
.Y(n_1408)
);

NAND2xp5_ASAP7_75t_L g1409 ( 
.A(n_1308),
.B(n_1177),
.Y(n_1409)
);

INVx3_ASAP7_75t_L g1410 ( 
.A(n_1294),
.Y(n_1410)
);

INVx1_ASAP7_75t_L g1411 ( 
.A(n_1237),
.Y(n_1411)
);

NAND2xp5_ASAP7_75t_L g1412 ( 
.A(n_1365),
.B(n_50),
.Y(n_1412)
);

BUFx6f_ASAP7_75t_L g1413 ( 
.A(n_1256),
.Y(n_1413)
);

NAND2xp5_ASAP7_75t_L g1414 ( 
.A(n_1317),
.B(n_52),
.Y(n_1414)
);

AOI22xp33_ASAP7_75t_L g1415 ( 
.A1(n_1269),
.A2(n_1201),
.B1(n_54),
.B2(n_52),
.Y(n_1415)
);

AOI22xp33_ASAP7_75t_L g1416 ( 
.A1(n_1250),
.A2(n_55),
.B1(n_53),
.B2(n_54),
.Y(n_1416)
);

INVx2_ASAP7_75t_SL g1417 ( 
.A(n_1246),
.Y(n_1417)
);

CKINVDCx5p33_ASAP7_75t_R g1418 ( 
.A(n_1248),
.Y(n_1418)
);

O2A1O1Ixp33_ASAP7_75t_L g1419 ( 
.A1(n_1242),
.A2(n_56),
.B(n_53),
.C(n_55),
.Y(n_1419)
);

NAND2xp5_ASAP7_75t_L g1420 ( 
.A(n_1363),
.B(n_56),
.Y(n_1420)
);

NAND2xp5_ASAP7_75t_L g1421 ( 
.A(n_1297),
.B(n_57),
.Y(n_1421)
);

NAND2xp5_ASAP7_75t_SL g1422 ( 
.A(n_1304),
.B(n_57),
.Y(n_1422)
);

INVx1_ASAP7_75t_SL g1423 ( 
.A(n_1309),
.Y(n_1423)
);

BUFx6f_ASAP7_75t_L g1424 ( 
.A(n_1256),
.Y(n_1424)
);

AND3x1_ASAP7_75t_SL g1425 ( 
.A(n_1258),
.B(n_58),
.C(n_59),
.Y(n_1425)
);

NAND2xp5_ASAP7_75t_L g1426 ( 
.A(n_1301),
.B(n_59),
.Y(n_1426)
);

AND2x4_ASAP7_75t_L g1427 ( 
.A(n_1254),
.B(n_513),
.Y(n_1427)
);

BUFx2_ASAP7_75t_L g1428 ( 
.A(n_1233),
.Y(n_1428)
);

AND2x4_ASAP7_75t_L g1429 ( 
.A(n_1254),
.B(n_314),
.Y(n_1429)
);

INVx6_ASAP7_75t_L g1430 ( 
.A(n_1241),
.Y(n_1430)
);

INVx1_ASAP7_75t_L g1431 ( 
.A(n_1257),
.Y(n_1431)
);

AND2x2_ASAP7_75t_L g1432 ( 
.A(n_1273),
.B(n_60),
.Y(n_1432)
);

NAND2xp5_ASAP7_75t_L g1433 ( 
.A(n_1382),
.B(n_60),
.Y(n_1433)
);

INVx2_ASAP7_75t_L g1434 ( 
.A(n_1276),
.Y(n_1434)
);

CKINVDCx20_ASAP7_75t_R g1435 ( 
.A(n_1360),
.Y(n_1435)
);

INVx1_ASAP7_75t_L g1436 ( 
.A(n_1286),
.Y(n_1436)
);

BUFx3_ASAP7_75t_L g1437 ( 
.A(n_1265),
.Y(n_1437)
);

AND2x4_ASAP7_75t_L g1438 ( 
.A(n_1336),
.B(n_511),
.Y(n_1438)
);

NAND2xp5_ASAP7_75t_L g1439 ( 
.A(n_1368),
.B(n_61),
.Y(n_1439)
);

BUFx6f_ASAP7_75t_L g1440 ( 
.A(n_1298),
.Y(n_1440)
);

NOR2xp33_ASAP7_75t_L g1441 ( 
.A(n_1380),
.B(n_62),
.Y(n_1441)
);

BUFx6f_ASAP7_75t_L g1442 ( 
.A(n_1298),
.Y(n_1442)
);

INVx2_ASAP7_75t_L g1443 ( 
.A(n_1291),
.Y(n_1443)
);

AOI211xp5_ASAP7_75t_L g1444 ( 
.A1(n_1339),
.A2(n_64),
.B(n_62),
.C(n_63),
.Y(n_1444)
);

INVx2_ASAP7_75t_SL g1445 ( 
.A(n_1315),
.Y(n_1445)
);

INVx1_ASAP7_75t_L g1446 ( 
.A(n_1293),
.Y(n_1446)
);

OR2x6_ASAP7_75t_L g1447 ( 
.A(n_1369),
.B(n_317),
.Y(n_1447)
);

NAND2xp5_ASAP7_75t_L g1448 ( 
.A(n_1372),
.B(n_63),
.Y(n_1448)
);

INVx1_ASAP7_75t_L g1449 ( 
.A(n_1277),
.Y(n_1449)
);

NOR2xp33_ASAP7_75t_L g1450 ( 
.A(n_1333),
.B(n_65),
.Y(n_1450)
);

BUFx4f_ASAP7_75t_SL g1451 ( 
.A(n_1359),
.Y(n_1451)
);

INVx2_ASAP7_75t_L g1452 ( 
.A(n_1306),
.Y(n_1452)
);

BUFx3_ASAP7_75t_L g1453 ( 
.A(n_1249),
.Y(n_1453)
);

INVxp67_ASAP7_75t_SL g1454 ( 
.A(n_1236),
.Y(n_1454)
);

CKINVDCx5p33_ASAP7_75t_R g1455 ( 
.A(n_1327),
.Y(n_1455)
);

NAND2xp5_ASAP7_75t_L g1456 ( 
.A(n_1384),
.B(n_66),
.Y(n_1456)
);

AND2x4_ASAP7_75t_L g1457 ( 
.A(n_1336),
.B(n_509),
.Y(n_1457)
);

NOR2xp33_ASAP7_75t_L g1458 ( 
.A(n_1391),
.B(n_67),
.Y(n_1458)
);

BUFx3_ASAP7_75t_L g1459 ( 
.A(n_1263),
.Y(n_1459)
);

NAND2xp5_ASAP7_75t_L g1460 ( 
.A(n_1362),
.B(n_69),
.Y(n_1460)
);

INVx2_ASAP7_75t_L g1461 ( 
.A(n_1307),
.Y(n_1461)
);

AOI21xp5_ASAP7_75t_L g1462 ( 
.A1(n_1278),
.A2(n_322),
.B(n_321),
.Y(n_1462)
);

BUFx2_ASAP7_75t_L g1463 ( 
.A(n_1337),
.Y(n_1463)
);

NAND2xp5_ASAP7_75t_L g1464 ( 
.A(n_1320),
.B(n_69),
.Y(n_1464)
);

AOI22xp5_ASAP7_75t_L g1465 ( 
.A1(n_1250),
.A2(n_72),
.B1(n_70),
.B2(n_71),
.Y(n_1465)
);

INVx2_ASAP7_75t_L g1466 ( 
.A(n_1288),
.Y(n_1466)
);

NOR2xp67_ASAP7_75t_L g1467 ( 
.A(n_1294),
.B(n_508),
.Y(n_1467)
);

NAND2xp5_ASAP7_75t_L g1468 ( 
.A(n_1252),
.B(n_74),
.Y(n_1468)
);

INVx4_ASAP7_75t_L g1469 ( 
.A(n_1326),
.Y(n_1469)
);

NOR2xp33_ASAP7_75t_L g1470 ( 
.A(n_1330),
.B(n_75),
.Y(n_1470)
);

AND3x1_ASAP7_75t_SL g1471 ( 
.A(n_1255),
.B(n_75),
.C(n_76),
.Y(n_1471)
);

BUFx2_ASAP7_75t_L g1472 ( 
.A(n_1348),
.Y(n_1472)
);

INVx2_ASAP7_75t_L g1473 ( 
.A(n_1261),
.Y(n_1473)
);

BUFx4f_ASAP7_75t_L g1474 ( 
.A(n_1343),
.Y(n_1474)
);

HB1xp67_ASAP7_75t_L g1475 ( 
.A(n_1311),
.Y(n_1475)
);

AND3x2_ASAP7_75t_SL g1476 ( 
.A(n_1342),
.B(n_76),
.C(n_77),
.Y(n_1476)
);

BUFx6f_ASAP7_75t_L g1477 ( 
.A(n_1298),
.Y(n_1477)
);

NAND2xp5_ASAP7_75t_L g1478 ( 
.A(n_1232),
.B(n_77),
.Y(n_1478)
);

CKINVDCx5p33_ASAP7_75t_R g1479 ( 
.A(n_1259),
.Y(n_1479)
);

INVx1_ASAP7_75t_L g1480 ( 
.A(n_1356),
.Y(n_1480)
);

BUFx5_ASAP7_75t_L g1481 ( 
.A(n_1353),
.Y(n_1481)
);

AND2x6_ASAP7_75t_SL g1482 ( 
.A(n_1314),
.B(n_78),
.Y(n_1482)
);

NAND2xp5_ASAP7_75t_L g1483 ( 
.A(n_1325),
.B(n_78),
.Y(n_1483)
);

INVx2_ASAP7_75t_SL g1484 ( 
.A(n_1272),
.Y(n_1484)
);

INVx2_ASAP7_75t_L g1485 ( 
.A(n_1244),
.Y(n_1485)
);

INVx2_ASAP7_75t_SL g1486 ( 
.A(n_1345),
.Y(n_1486)
);

INVx2_ASAP7_75t_L g1487 ( 
.A(n_1245),
.Y(n_1487)
);

NAND2xp5_ASAP7_75t_L g1488 ( 
.A(n_1329),
.B(n_79),
.Y(n_1488)
);

BUFx3_ASAP7_75t_L g1489 ( 
.A(n_1345),
.Y(n_1489)
);

HB1xp67_ASAP7_75t_L g1490 ( 
.A(n_1326),
.Y(n_1490)
);

INVx1_ASAP7_75t_L g1491 ( 
.A(n_1388),
.Y(n_1491)
);

INVx2_ASAP7_75t_L g1492 ( 
.A(n_1247),
.Y(n_1492)
);

NAND2xp5_ASAP7_75t_L g1493 ( 
.A(n_1331),
.B(n_80),
.Y(n_1493)
);

AND2x2_ASAP7_75t_L g1494 ( 
.A(n_1243),
.B(n_81),
.Y(n_1494)
);

AND2x2_ASAP7_75t_L g1495 ( 
.A(n_1328),
.B(n_81),
.Y(n_1495)
);

INVx3_ASAP7_75t_L g1496 ( 
.A(n_1343),
.Y(n_1496)
);

NAND2xp5_ASAP7_75t_SL g1497 ( 
.A(n_1275),
.B(n_82),
.Y(n_1497)
);

INVx1_ASAP7_75t_L g1498 ( 
.A(n_1332),
.Y(n_1498)
);

NAND2xp5_ASAP7_75t_SL g1499 ( 
.A(n_1275),
.B(n_82),
.Y(n_1499)
);

OR2x2_ASAP7_75t_L g1500 ( 
.A(n_1292),
.B(n_83),
.Y(n_1500)
);

NAND2xp5_ASAP7_75t_SL g1501 ( 
.A(n_1280),
.B(n_83),
.Y(n_1501)
);

NAND2xp5_ASAP7_75t_L g1502 ( 
.A(n_1346),
.B(n_84),
.Y(n_1502)
);

AND2x4_ASAP7_75t_L g1503 ( 
.A(n_1390),
.B(n_325),
.Y(n_1503)
);

INVx1_ASAP7_75t_L g1504 ( 
.A(n_1324),
.Y(n_1504)
);

NAND2xp5_ASAP7_75t_SL g1505 ( 
.A(n_1280),
.B(n_84),
.Y(n_1505)
);

BUFx2_ASAP7_75t_L g1506 ( 
.A(n_1303),
.Y(n_1506)
);

INVxp67_ASAP7_75t_SL g1507 ( 
.A(n_1279),
.Y(n_1507)
);

NOR2xp33_ASAP7_75t_L g1508 ( 
.A(n_1385),
.B(n_85),
.Y(n_1508)
);

NAND2xp5_ASAP7_75t_L g1509 ( 
.A(n_1282),
.B(n_85),
.Y(n_1509)
);

BUFx12f_ASAP7_75t_L g1510 ( 
.A(n_1370),
.Y(n_1510)
);

NOR2xp33_ASAP7_75t_L g1511 ( 
.A(n_1393),
.B(n_86),
.Y(n_1511)
);

CKINVDCx16_ASAP7_75t_R g1512 ( 
.A(n_1361),
.Y(n_1512)
);

INVx2_ASAP7_75t_L g1513 ( 
.A(n_1350),
.Y(n_1513)
);

BUFx2_ASAP7_75t_L g1514 ( 
.A(n_1303),
.Y(n_1514)
);

INVx5_ASAP7_75t_L g1515 ( 
.A(n_1343),
.Y(n_1515)
);

AND2x2_ASAP7_75t_L g1516 ( 
.A(n_1266),
.B(n_86),
.Y(n_1516)
);

CKINVDCx6p67_ASAP7_75t_R g1517 ( 
.A(n_1326),
.Y(n_1517)
);

BUFx2_ASAP7_75t_L g1518 ( 
.A(n_1287),
.Y(n_1518)
);

BUFx3_ASAP7_75t_L g1519 ( 
.A(n_1370),
.Y(n_1519)
);

INVx1_ASAP7_75t_L g1520 ( 
.A(n_1351),
.Y(n_1520)
);

INVx2_ASAP7_75t_L g1521 ( 
.A(n_1357),
.Y(n_1521)
);

INVx2_ASAP7_75t_L g1522 ( 
.A(n_1387),
.Y(n_1522)
);

AND3x1_ASAP7_75t_SL g1523 ( 
.A(n_1260),
.B(n_1389),
.C(n_1400),
.Y(n_1523)
);

NOR2xp33_ASAP7_75t_SL g1524 ( 
.A(n_1394),
.B(n_326),
.Y(n_1524)
);

BUFx2_ASAP7_75t_L g1525 ( 
.A(n_1370),
.Y(n_1525)
);

A2O1A1Ixp33_ASAP7_75t_L g1526 ( 
.A1(n_1334),
.A2(n_89),
.B(n_87),
.C(n_88),
.Y(n_1526)
);

INVx2_ASAP7_75t_L g1527 ( 
.A(n_1387),
.Y(n_1527)
);

NAND2xp5_ASAP7_75t_L g1528 ( 
.A(n_1355),
.B(n_88),
.Y(n_1528)
);

AOI22xp33_ASAP7_75t_L g1529 ( 
.A1(n_1250),
.A2(n_91),
.B1(n_89),
.B2(n_90),
.Y(n_1529)
);

INVx1_ASAP7_75t_L g1530 ( 
.A(n_1253),
.Y(n_1530)
);

NAND2xp5_ASAP7_75t_L g1531 ( 
.A(n_1349),
.B(n_90),
.Y(n_1531)
);

NAND2xp33_ASAP7_75t_SL g1532 ( 
.A(n_1239),
.B(n_91),
.Y(n_1532)
);

AND2x4_ASAP7_75t_L g1533 ( 
.A(n_1386),
.B(n_327),
.Y(n_1533)
);

INVx2_ASAP7_75t_SL g1534 ( 
.A(n_1386),
.Y(n_1534)
);

AND2x2_ASAP7_75t_L g1535 ( 
.A(n_1375),
.B(n_92),
.Y(n_1535)
);

NAND2xp5_ASAP7_75t_L g1536 ( 
.A(n_1295),
.B(n_94),
.Y(n_1536)
);

AND2x4_ASAP7_75t_L g1537 ( 
.A(n_1386),
.B(n_507),
.Y(n_1537)
);

BUFx3_ASAP7_75t_L g1538 ( 
.A(n_1335),
.Y(n_1538)
);

INVx1_ASAP7_75t_L g1539 ( 
.A(n_1264),
.Y(n_1539)
);

BUFx6f_ASAP7_75t_L g1540 ( 
.A(n_1396),
.Y(n_1540)
);

AND2x4_ASAP7_75t_L g1541 ( 
.A(n_1302),
.B(n_330),
.Y(n_1541)
);

AOI221xp5_ASAP7_75t_L g1542 ( 
.A1(n_1274),
.A2(n_97),
.B1(n_95),
.B2(n_96),
.C(n_98),
.Y(n_1542)
);

CKINVDCx5p33_ASAP7_75t_R g1543 ( 
.A(n_1396),
.Y(n_1543)
);

INVx2_ASAP7_75t_L g1544 ( 
.A(n_1341),
.Y(n_1544)
);

NAND2xp5_ASAP7_75t_L g1545 ( 
.A(n_1299),
.B(n_95),
.Y(n_1545)
);

BUFx3_ASAP7_75t_L g1546 ( 
.A(n_1335),
.Y(n_1546)
);

BUFx3_ASAP7_75t_L g1547 ( 
.A(n_1352),
.Y(n_1547)
);

BUFx6f_ASAP7_75t_L g1548 ( 
.A(n_1373),
.Y(n_1548)
);

HB1xp67_ASAP7_75t_L g1549 ( 
.A(n_1399),
.Y(n_1549)
);

INVx4_ASAP7_75t_L g1550 ( 
.A(n_1374),
.Y(n_1550)
);

NAND2xp5_ASAP7_75t_SL g1551 ( 
.A(n_1367),
.B(n_96),
.Y(n_1551)
);

OR2x2_ASAP7_75t_L g1552 ( 
.A(n_1300),
.B(n_1312),
.Y(n_1552)
);

INVx3_ASAP7_75t_L g1553 ( 
.A(n_1354),
.Y(n_1553)
);

NAND2xp5_ASAP7_75t_L g1554 ( 
.A(n_1313),
.B(n_97),
.Y(n_1554)
);

BUFx4f_ASAP7_75t_L g1555 ( 
.A(n_1234),
.Y(n_1555)
);

NAND2xp5_ASAP7_75t_SL g1556 ( 
.A(n_1373),
.B(n_98),
.Y(n_1556)
);

INVx1_ASAP7_75t_SL g1557 ( 
.A(n_1268),
.Y(n_1557)
);

NAND2xp5_ASAP7_75t_L g1558 ( 
.A(n_1322),
.B(n_99),
.Y(n_1558)
);

INVx3_ASAP7_75t_L g1559 ( 
.A(n_1364),
.Y(n_1559)
);

BUFx6f_ASAP7_75t_L g1560 ( 
.A(n_1378),
.Y(n_1560)
);

AND2x4_ASAP7_75t_L g1561 ( 
.A(n_1398),
.B(n_331),
.Y(n_1561)
);

NAND2xp5_ASAP7_75t_SL g1562 ( 
.A(n_1378),
.B(n_100),
.Y(n_1562)
);

OR2x2_ASAP7_75t_L g1563 ( 
.A(n_1281),
.B(n_100),
.Y(n_1563)
);

NAND2xp5_ASAP7_75t_L g1564 ( 
.A(n_1449),
.B(n_1358),
.Y(n_1564)
);

INVxp67_ASAP7_75t_SL g1565 ( 
.A(n_1408),
.Y(n_1565)
);

AOI21x1_ASAP7_75t_L g1566 ( 
.A1(n_1402),
.A2(n_1392),
.B(n_1371),
.Y(n_1566)
);

INVx1_ASAP7_75t_L g1567 ( 
.A(n_1498),
.Y(n_1567)
);

BUFx6f_ASAP7_75t_L g1568 ( 
.A(n_1474),
.Y(n_1568)
);

OAI22x1_ASAP7_75t_L g1569 ( 
.A1(n_1465),
.A2(n_1551),
.B1(n_1502),
.B2(n_1458),
.Y(n_1569)
);

NOR2xp33_ASAP7_75t_L g1570 ( 
.A(n_1423),
.B(n_1338),
.Y(n_1570)
);

NAND3xp33_ASAP7_75t_L g1571 ( 
.A(n_1444),
.B(n_1397),
.C(n_1366),
.Y(n_1571)
);

BUFx2_ASAP7_75t_L g1572 ( 
.A(n_1455),
.Y(n_1572)
);

OAI21x1_ASAP7_75t_L g1573 ( 
.A1(n_1462),
.A2(n_1340),
.B(n_1262),
.Y(n_1573)
);

INVx2_ASAP7_75t_SL g1574 ( 
.A(n_1430),
.Y(n_1574)
);

AOI21x1_ASAP7_75t_L g1575 ( 
.A1(n_1509),
.A2(n_1340),
.B(n_1395),
.Y(n_1575)
);

NAND2xp5_ASAP7_75t_L g1576 ( 
.A(n_1530),
.B(n_1377),
.Y(n_1576)
);

INVx2_ASAP7_75t_L g1577 ( 
.A(n_1443),
.Y(n_1577)
);

OAI21x1_ASAP7_75t_SL g1578 ( 
.A1(n_1528),
.A2(n_1379),
.B(n_1376),
.Y(n_1578)
);

AOI21xp5_ASAP7_75t_L g1579 ( 
.A1(n_1555),
.A2(n_1383),
.B(n_1284),
.Y(n_1579)
);

NOR2xp67_ASAP7_75t_SL g1580 ( 
.A(n_1550),
.B(n_1374),
.Y(n_1580)
);

OAI22xp5_ASAP7_75t_L g1581 ( 
.A1(n_1557),
.A2(n_1285),
.B1(n_1316),
.B2(n_1374),
.Y(n_1581)
);

AND2x2_ASAP7_75t_L g1582 ( 
.A(n_1549),
.B(n_1494),
.Y(n_1582)
);

INVx1_ASAP7_75t_L g1583 ( 
.A(n_1491),
.Y(n_1583)
);

AOI21xp5_ASAP7_75t_L g1584 ( 
.A1(n_1409),
.A2(n_1383),
.B(n_1283),
.Y(n_1584)
);

BUFx2_ASAP7_75t_L g1585 ( 
.A(n_1463),
.Y(n_1585)
);

OAI21x1_ASAP7_75t_L g1586 ( 
.A1(n_1491),
.A2(n_1296),
.B(n_1289),
.Y(n_1586)
);

AOI22xp33_ASAP7_75t_L g1587 ( 
.A1(n_1532),
.A2(n_1267),
.B1(n_1238),
.B2(n_1234),
.Y(n_1587)
);

NOR2x1_ASAP7_75t_L g1588 ( 
.A(n_1550),
.B(n_1323),
.Y(n_1588)
);

NOR2xp33_ASAP7_75t_L g1589 ( 
.A(n_1552),
.B(n_1338),
.Y(n_1589)
);

INVx3_ASAP7_75t_L g1590 ( 
.A(n_1474),
.Y(n_1590)
);

OAI21x1_ASAP7_75t_L g1591 ( 
.A1(n_1480),
.A2(n_1321),
.B(n_1251),
.Y(n_1591)
);

OAI22xp5_ASAP7_75t_L g1592 ( 
.A1(n_1539),
.A2(n_1240),
.B1(n_1305),
.B2(n_1270),
.Y(n_1592)
);

O2A1O1Ixp33_ASAP7_75t_L g1593 ( 
.A1(n_1556),
.A2(n_1267),
.B(n_1238),
.C(n_1234),
.Y(n_1593)
);

OAI21xp33_ASAP7_75t_L g1594 ( 
.A1(n_1511),
.A2(n_1318),
.B(n_1347),
.Y(n_1594)
);

OAI22xp33_ASAP7_75t_L g1595 ( 
.A1(n_1524),
.A2(n_1267),
.B1(n_1238),
.B2(n_1234),
.Y(n_1595)
);

INVx5_ASAP7_75t_L g1596 ( 
.A(n_1469),
.Y(n_1596)
);

OAI22xp5_ASAP7_75t_L g1597 ( 
.A1(n_1548),
.A2(n_1238),
.B1(n_1381),
.B2(n_1319),
.Y(n_1597)
);

INVx3_ASAP7_75t_L g1598 ( 
.A(n_1515),
.Y(n_1598)
);

INVx1_ASAP7_75t_L g1599 ( 
.A(n_1403),
.Y(n_1599)
);

AOI211x1_ASAP7_75t_L g1600 ( 
.A1(n_1562),
.A2(n_103),
.B(n_101),
.C(n_102),
.Y(n_1600)
);

AOI21x1_ASAP7_75t_SL g1601 ( 
.A1(n_1488),
.A2(n_1353),
.B(n_1319),
.Y(n_1601)
);

CKINVDCx5p33_ASAP7_75t_R g1602 ( 
.A(n_1418),
.Y(n_1602)
);

BUFx2_ASAP7_75t_L g1603 ( 
.A(n_1472),
.Y(n_1603)
);

INVx1_ASAP7_75t_L g1604 ( 
.A(n_1446),
.Y(n_1604)
);

AOI21x1_ASAP7_75t_L g1605 ( 
.A1(n_1478),
.A2(n_1319),
.B(n_333),
.Y(n_1605)
);

BUFx6f_ASAP7_75t_L g1606 ( 
.A(n_1515),
.Y(n_1606)
);

OAI21x1_ASAP7_75t_L g1607 ( 
.A1(n_1553),
.A2(n_334),
.B(n_332),
.Y(n_1607)
);

AO31x2_ASAP7_75t_L g1608 ( 
.A1(n_1526),
.A2(n_1558),
.A3(n_1531),
.B(n_1446),
.Y(n_1608)
);

AND2x2_ASAP7_75t_L g1609 ( 
.A(n_1535),
.B(n_102),
.Y(n_1609)
);

AND2x2_ASAP7_75t_L g1610 ( 
.A(n_1516),
.B(n_103),
.Y(n_1610)
);

AND2x2_ASAP7_75t_L g1611 ( 
.A(n_1432),
.B(n_104),
.Y(n_1611)
);

OAI21xp5_ASAP7_75t_L g1612 ( 
.A1(n_1536),
.A2(n_104),
.B(n_105),
.Y(n_1612)
);

NAND2xp5_ASAP7_75t_L g1613 ( 
.A(n_1460),
.B(n_105),
.Y(n_1613)
);

AOI21xp5_ASAP7_75t_L g1614 ( 
.A1(n_1544),
.A2(n_337),
.B(n_336),
.Y(n_1614)
);

BUFx3_ASAP7_75t_L g1615 ( 
.A(n_1430),
.Y(n_1615)
);

NAND3xp33_ASAP7_75t_L g1616 ( 
.A(n_1542),
.B(n_106),
.C(n_107),
.Y(n_1616)
);

INVx4_ASAP7_75t_L g1617 ( 
.A(n_1515),
.Y(n_1617)
);

OAI21x1_ASAP7_75t_L g1618 ( 
.A1(n_1559),
.A2(n_342),
.B(n_338),
.Y(n_1618)
);

BUFx2_ASAP7_75t_L g1619 ( 
.A(n_1543),
.Y(n_1619)
);

OAI21x1_ASAP7_75t_L g1620 ( 
.A1(n_1559),
.A2(n_345),
.B(n_344),
.Y(n_1620)
);

AO31x2_ASAP7_75t_L g1621 ( 
.A1(n_1545),
.A2(n_108),
.A3(n_106),
.B(n_107),
.Y(n_1621)
);

NAND2xp5_ASAP7_75t_SL g1622 ( 
.A(n_1548),
.B(n_108),
.Y(n_1622)
);

OAI21x1_ASAP7_75t_SL g1623 ( 
.A1(n_1439),
.A2(n_109),
.B(n_110),
.Y(n_1623)
);

AO21x2_ASAP7_75t_L g1624 ( 
.A1(n_1554),
.A2(n_355),
.B(n_353),
.Y(n_1624)
);

INVxp67_ASAP7_75t_L g1625 ( 
.A(n_1475),
.Y(n_1625)
);

OAI21x1_ASAP7_75t_L g1626 ( 
.A1(n_1504),
.A2(n_358),
.B(n_356),
.Y(n_1626)
);

OAI21xp5_ASAP7_75t_L g1627 ( 
.A1(n_1419),
.A2(n_109),
.B(n_111),
.Y(n_1627)
);

AND2x2_ASAP7_75t_L g1628 ( 
.A(n_1495),
.B(n_113),
.Y(n_1628)
);

AOI21xp5_ASAP7_75t_L g1629 ( 
.A1(n_1507),
.A2(n_360),
.B(n_359),
.Y(n_1629)
);

INVx3_ASAP7_75t_L g1630 ( 
.A(n_1496),
.Y(n_1630)
);

AO31x2_ASAP7_75t_L g1631 ( 
.A1(n_1420),
.A2(n_116),
.A3(n_114),
.B(n_115),
.Y(n_1631)
);

NAND2xp5_ASAP7_75t_L g1632 ( 
.A(n_1548),
.B(n_1560),
.Y(n_1632)
);

BUFx3_ASAP7_75t_L g1633 ( 
.A(n_1437),
.Y(n_1633)
);

OAI21xp5_ASAP7_75t_L g1634 ( 
.A1(n_1433),
.A2(n_115),
.B(n_116),
.Y(n_1634)
);

OAI21xp5_ASAP7_75t_L g1635 ( 
.A1(n_1448),
.A2(n_117),
.B(n_118),
.Y(n_1635)
);

AOI21xp5_ASAP7_75t_L g1636 ( 
.A1(n_1521),
.A2(n_506),
.B(n_368),
.Y(n_1636)
);

OAI21x1_ASAP7_75t_L g1637 ( 
.A1(n_1411),
.A2(n_369),
.B(n_365),
.Y(n_1637)
);

NAND2xp5_ASAP7_75t_L g1638 ( 
.A(n_1560),
.B(n_117),
.Y(n_1638)
);

OAI22xp5_ASAP7_75t_L g1639 ( 
.A1(n_1560),
.A2(n_120),
.B1(n_118),
.B2(n_119),
.Y(n_1639)
);

OAI21x1_ASAP7_75t_L g1640 ( 
.A1(n_1431),
.A2(n_371),
.B(n_370),
.Y(n_1640)
);

OAI22xp5_ASAP7_75t_L g1641 ( 
.A1(n_1416),
.A2(n_121),
.B1(n_119),
.B2(n_120),
.Y(n_1641)
);

OAI21x1_ASAP7_75t_L g1642 ( 
.A1(n_1436),
.A2(n_375),
.B(n_373),
.Y(n_1642)
);

NAND2xp5_ASAP7_75t_L g1643 ( 
.A(n_1456),
.B(n_121),
.Y(n_1643)
);

AOI221xp5_ASAP7_75t_SL g1644 ( 
.A1(n_1529),
.A2(n_1450),
.B1(n_1483),
.B2(n_1415),
.C(n_1422),
.Y(n_1644)
);

AOI21x1_ASAP7_75t_L g1645 ( 
.A1(n_1493),
.A2(n_377),
.B(n_376),
.Y(n_1645)
);

AOI21xp5_ASAP7_75t_SL g1646 ( 
.A1(n_1438),
.A2(n_379),
.B(n_378),
.Y(n_1646)
);

NAND2xp5_ASAP7_75t_L g1647 ( 
.A(n_1414),
.B(n_123),
.Y(n_1647)
);

OAI21x1_ASAP7_75t_L g1648 ( 
.A1(n_1522),
.A2(n_383),
.B(n_382),
.Y(n_1648)
);

AOI21xp5_ASAP7_75t_L g1649 ( 
.A1(n_1438),
.A2(n_386),
.B(n_384),
.Y(n_1649)
);

AND2x2_ASAP7_75t_L g1650 ( 
.A(n_1457),
.B(n_123),
.Y(n_1650)
);

OAI21x1_ASAP7_75t_SL g1651 ( 
.A1(n_1421),
.A2(n_124),
.B(n_125),
.Y(n_1651)
);

NAND2x1p5_ASAP7_75t_L g1652 ( 
.A(n_1469),
.B(n_387),
.Y(n_1652)
);

HB1xp67_ASAP7_75t_L g1653 ( 
.A(n_1454),
.Y(n_1653)
);

NAND2xp5_ASAP7_75t_SL g1654 ( 
.A(n_1561),
.B(n_126),
.Y(n_1654)
);

OAI22xp5_ASAP7_75t_L g1655 ( 
.A1(n_1407),
.A2(n_127),
.B1(n_128),
.B2(n_129),
.Y(n_1655)
);

AND2x2_ASAP7_75t_L g1656 ( 
.A(n_1457),
.B(n_127),
.Y(n_1656)
);

AOI21xp5_ASAP7_75t_L g1657 ( 
.A1(n_1541),
.A2(n_504),
.B(n_389),
.Y(n_1657)
);

INVx1_ASAP7_75t_SL g1658 ( 
.A(n_1525),
.Y(n_1658)
);

AOI21xp5_ASAP7_75t_L g1659 ( 
.A1(n_1541),
.A2(n_502),
.B(n_390),
.Y(n_1659)
);

AND2x2_ASAP7_75t_L g1660 ( 
.A(n_1427),
.B(n_129),
.Y(n_1660)
);

OR2x2_ASAP7_75t_L g1661 ( 
.A(n_1500),
.B(n_130),
.Y(n_1661)
);

OAI21xp5_ASAP7_75t_L g1662 ( 
.A1(n_1412),
.A2(n_130),
.B(n_131),
.Y(n_1662)
);

OAI21x1_ASAP7_75t_L g1663 ( 
.A1(n_1527),
.A2(n_393),
.B(n_388),
.Y(n_1663)
);

NAND2x1p5_ASAP7_75t_L g1664 ( 
.A(n_1404),
.B(n_397),
.Y(n_1664)
);

CKINVDCx5p33_ASAP7_75t_R g1665 ( 
.A(n_1435),
.Y(n_1665)
);

NAND2xp5_ASAP7_75t_L g1666 ( 
.A(n_1464),
.B(n_1426),
.Y(n_1666)
);

NAND2xp5_ASAP7_75t_L g1667 ( 
.A(n_1434),
.B(n_131),
.Y(n_1667)
);

AOI22xp5_ASAP7_75t_L g1668 ( 
.A1(n_1523),
.A2(n_1499),
.B1(n_1501),
.B2(n_1497),
.Y(n_1668)
);

OAI21x1_ASAP7_75t_L g1669 ( 
.A1(n_1452),
.A2(n_401),
.B(n_399),
.Y(n_1669)
);

INVx1_ASAP7_75t_L g1670 ( 
.A(n_1461),
.Y(n_1670)
);

AO21x1_ASAP7_75t_L g1671 ( 
.A1(n_1468),
.A2(n_132),
.B(n_133),
.Y(n_1671)
);

NAND2xp5_ASAP7_75t_L g1672 ( 
.A(n_1520),
.B(n_132),
.Y(n_1672)
);

NAND2xp5_ASAP7_75t_L g1673 ( 
.A(n_1505),
.B(n_133),
.Y(n_1673)
);

CKINVDCx8_ASAP7_75t_R g1674 ( 
.A(n_1428),
.Y(n_1674)
);

NAND2xp5_ASAP7_75t_L g1675 ( 
.A(n_1563),
.B(n_134),
.Y(n_1675)
);

INVx3_ASAP7_75t_L g1676 ( 
.A(n_1496),
.Y(n_1676)
);

NAND2xp5_ASAP7_75t_L g1677 ( 
.A(n_1427),
.B(n_1429),
.Y(n_1677)
);

A2O1A1Ixp33_ASAP7_75t_L g1678 ( 
.A1(n_1508),
.A2(n_1441),
.B(n_1503),
.C(n_1561),
.Y(n_1678)
);

AOI22xp5_ASAP7_75t_L g1679 ( 
.A1(n_1429),
.A2(n_134),
.B1(n_135),
.B2(n_136),
.Y(n_1679)
);

INVx4_ASAP7_75t_L g1680 ( 
.A(n_1517),
.Y(n_1680)
);

NAND2xp5_ASAP7_75t_L g1681 ( 
.A(n_1466),
.B(n_136),
.Y(n_1681)
);

OAI22xp5_ASAP7_75t_L g1682 ( 
.A1(n_1538),
.A2(n_137),
.B1(n_139),
.B2(n_140),
.Y(n_1682)
);

NAND2xp5_ASAP7_75t_L g1683 ( 
.A(n_1473),
.B(n_139),
.Y(n_1683)
);

INVx1_ASAP7_75t_L g1684 ( 
.A(n_1513),
.Y(n_1684)
);

OAI21x1_ASAP7_75t_L g1685 ( 
.A1(n_1485),
.A2(n_404),
.B(n_403),
.Y(n_1685)
);

NAND2xp5_ASAP7_75t_L g1686 ( 
.A(n_1547),
.B(n_140),
.Y(n_1686)
);

AND2x2_ASAP7_75t_L g1687 ( 
.A(n_1503),
.B(n_141),
.Y(n_1687)
);

OAI21x1_ASAP7_75t_SL g1688 ( 
.A1(n_1487),
.A2(n_142),
.B(n_143),
.Y(n_1688)
);

HB1xp67_ASAP7_75t_L g1689 ( 
.A(n_1445),
.Y(n_1689)
);

INVx1_ASAP7_75t_L g1690 ( 
.A(n_1481),
.Y(n_1690)
);

OAI21x1_ASAP7_75t_L g1691 ( 
.A1(n_1492),
.A2(n_406),
.B(n_405),
.Y(n_1691)
);

INVx2_ASAP7_75t_L g1692 ( 
.A(n_1540),
.Y(n_1692)
);

AO21x2_ASAP7_75t_L g1693 ( 
.A1(n_1467),
.A2(n_410),
.B(n_409),
.Y(n_1693)
);

NAND2xp5_ASAP7_75t_L g1694 ( 
.A(n_1546),
.B(n_142),
.Y(n_1694)
);

AOI21xp5_ASAP7_75t_L g1695 ( 
.A1(n_1533),
.A2(n_501),
.B(n_414),
.Y(n_1695)
);

AOI21xp5_ASAP7_75t_L g1696 ( 
.A1(n_1533),
.A2(n_499),
.B(n_415),
.Y(n_1696)
);

CKINVDCx5p33_ASAP7_75t_R g1697 ( 
.A(n_1451),
.Y(n_1697)
);

CKINVDCx6p67_ASAP7_75t_R g1698 ( 
.A(n_1489),
.Y(n_1698)
);

INVx1_ASAP7_75t_L g1699 ( 
.A(n_1481),
.Y(n_1699)
);

NAND2xp5_ASAP7_75t_SL g1700 ( 
.A(n_1540),
.B(n_143),
.Y(n_1700)
);

INVx1_ASAP7_75t_L g1701 ( 
.A(n_1583),
.Y(n_1701)
);

OAI21xp5_ASAP7_75t_L g1702 ( 
.A1(n_1594),
.A2(n_1406),
.B(n_1470),
.Y(n_1702)
);

NAND2xp5_ASAP7_75t_L g1703 ( 
.A(n_1589),
.B(n_1540),
.Y(n_1703)
);

OAI21x1_ASAP7_75t_SL g1704 ( 
.A1(n_1578),
.A2(n_1534),
.B(n_1471),
.Y(n_1704)
);

BUFx6f_ASAP7_75t_L g1705 ( 
.A(n_1568),
.Y(n_1705)
);

HB1xp67_ASAP7_75t_L g1706 ( 
.A(n_1653),
.Y(n_1706)
);

AOI21xp5_ASAP7_75t_L g1707 ( 
.A1(n_1595),
.A2(n_1593),
.B(n_1584),
.Y(n_1707)
);

OAI21xp33_ASAP7_75t_L g1708 ( 
.A1(n_1627),
.A2(n_1537),
.B(n_1447),
.Y(n_1708)
);

AOI21xp5_ASAP7_75t_L g1709 ( 
.A1(n_1592),
.A2(n_1410),
.B(n_1404),
.Y(n_1709)
);

INVx5_ASAP7_75t_L g1710 ( 
.A(n_1606),
.Y(n_1710)
);

AOI21xp5_ASAP7_75t_L g1711 ( 
.A1(n_1597),
.A2(n_1481),
.B(n_1447),
.Y(n_1711)
);

INVx2_ASAP7_75t_L g1712 ( 
.A(n_1577),
.Y(n_1712)
);

OR2x2_ASAP7_75t_L g1713 ( 
.A(n_1565),
.B(n_1519),
.Y(n_1713)
);

AND2x4_ASAP7_75t_L g1714 ( 
.A(n_1692),
.B(n_1506),
.Y(n_1714)
);

NAND2xp5_ASAP7_75t_L g1715 ( 
.A(n_1666),
.B(n_1406),
.Y(n_1715)
);

CKINVDCx5p33_ASAP7_75t_R g1716 ( 
.A(n_1602),
.Y(n_1716)
);

A2O1A1Ixp33_ASAP7_75t_L g1717 ( 
.A1(n_1678),
.A2(n_1571),
.B(n_1587),
.C(n_1616),
.Y(n_1717)
);

INVx1_ASAP7_75t_SL g1718 ( 
.A(n_1572),
.Y(n_1718)
);

NOR2xp67_ASAP7_75t_L g1719 ( 
.A(n_1574),
.B(n_1510),
.Y(n_1719)
);

AND2x4_ASAP7_75t_L g1720 ( 
.A(n_1632),
.B(n_1514),
.Y(n_1720)
);

CKINVDCx5p33_ASAP7_75t_R g1721 ( 
.A(n_1665),
.Y(n_1721)
);

AOI22xp33_ASAP7_75t_L g1722 ( 
.A1(n_1569),
.A2(n_1406),
.B1(n_1405),
.B2(n_1481),
.Y(n_1722)
);

BUFx3_ASAP7_75t_L g1723 ( 
.A(n_1615),
.Y(n_1723)
);

AND2x2_ASAP7_75t_L g1724 ( 
.A(n_1582),
.B(n_1518),
.Y(n_1724)
);

NAND2xp5_ASAP7_75t_L g1725 ( 
.A(n_1564),
.B(n_1406),
.Y(n_1725)
);

O2A1O1Ixp33_ASAP7_75t_SL g1726 ( 
.A1(n_1612),
.A2(n_1476),
.B(n_1490),
.C(n_1484),
.Y(n_1726)
);

BUFx12f_ASAP7_75t_L g1727 ( 
.A(n_1697),
.Y(n_1727)
);

BUFx6f_ASAP7_75t_L g1728 ( 
.A(n_1568),
.Y(n_1728)
);

OAI22xp5_ASAP7_75t_L g1729 ( 
.A1(n_1668),
.A2(n_1479),
.B1(n_1453),
.B2(n_1459),
.Y(n_1729)
);

BUFx2_ASAP7_75t_L g1730 ( 
.A(n_1585),
.Y(n_1730)
);

BUFx12f_ASAP7_75t_L g1731 ( 
.A(n_1568),
.Y(n_1731)
);

OAI22xp5_ASAP7_75t_L g1732 ( 
.A1(n_1570),
.A2(n_1417),
.B1(n_1486),
.B2(n_1512),
.Y(n_1732)
);

INVx1_ASAP7_75t_L g1733 ( 
.A(n_1583),
.Y(n_1733)
);

AOI21xp5_ASAP7_75t_L g1734 ( 
.A1(n_1579),
.A2(n_1413),
.B(n_1401),
.Y(n_1734)
);

INVx1_ASAP7_75t_SL g1735 ( 
.A(n_1603),
.Y(n_1735)
);

AND2x2_ASAP7_75t_L g1736 ( 
.A(n_1609),
.B(n_1401),
.Y(n_1736)
);

O2A1O1Ixp33_ASAP7_75t_L g1737 ( 
.A1(n_1634),
.A2(n_1482),
.B(n_1425),
.C(n_1405),
.Y(n_1737)
);

INVx1_ASAP7_75t_L g1738 ( 
.A(n_1567),
.Y(n_1738)
);

AND2x2_ASAP7_75t_L g1739 ( 
.A(n_1610),
.B(n_1413),
.Y(n_1739)
);

AOI22xp33_ASAP7_75t_L g1740 ( 
.A1(n_1635),
.A2(n_1477),
.B1(n_1442),
.B2(n_1440),
.Y(n_1740)
);

INVx3_ASAP7_75t_SL g1741 ( 
.A(n_1698),
.Y(n_1741)
);

INVx2_ASAP7_75t_SL g1742 ( 
.A(n_1633),
.Y(n_1742)
);

NOR2xp33_ASAP7_75t_L g1743 ( 
.A(n_1677),
.B(n_1413),
.Y(n_1743)
);

NOR2xp33_ASAP7_75t_L g1744 ( 
.A(n_1576),
.B(n_1619),
.Y(n_1744)
);

BUFx3_ASAP7_75t_L g1745 ( 
.A(n_1674),
.Y(n_1745)
);

HB1xp67_ASAP7_75t_L g1746 ( 
.A(n_1567),
.Y(n_1746)
);

NOR2xp33_ASAP7_75t_R g1747 ( 
.A(n_1590),
.B(n_1424),
.Y(n_1747)
);

NAND2xp5_ASAP7_75t_SL g1748 ( 
.A(n_1644),
.B(n_1424),
.Y(n_1748)
);

CKINVDCx8_ASAP7_75t_R g1749 ( 
.A(n_1606),
.Y(n_1749)
);

AOI22xp33_ASAP7_75t_L g1750 ( 
.A1(n_1662),
.A2(n_1477),
.B1(n_1442),
.B2(n_1440),
.Y(n_1750)
);

BUFx6f_ASAP7_75t_L g1751 ( 
.A(n_1606),
.Y(n_1751)
);

NOR2xp33_ASAP7_75t_L g1752 ( 
.A(n_1625),
.B(n_1442),
.Y(n_1752)
);

BUFx3_ASAP7_75t_L g1753 ( 
.A(n_1689),
.Y(n_1753)
);

INVx2_ASAP7_75t_L g1754 ( 
.A(n_1670),
.Y(n_1754)
);

OAI21xp5_ASAP7_75t_L g1755 ( 
.A1(n_1566),
.A2(n_1477),
.B(n_144),
.Y(n_1755)
);

NOR2x1_ASAP7_75t_SL g1756 ( 
.A(n_1690),
.B(n_413),
.Y(n_1756)
);

AOI22xp5_ASAP7_75t_L g1757 ( 
.A1(n_1654),
.A2(n_145),
.B1(n_146),
.B2(n_148),
.Y(n_1757)
);

AND2x4_ASAP7_75t_L g1758 ( 
.A(n_1590),
.B(n_416),
.Y(n_1758)
);

CKINVDCx20_ASAP7_75t_R g1759 ( 
.A(n_1658),
.Y(n_1759)
);

AOI21xp5_ASAP7_75t_L g1760 ( 
.A1(n_1573),
.A2(n_418),
.B(n_417),
.Y(n_1760)
);

AND2x2_ASAP7_75t_L g1761 ( 
.A(n_1660),
.B(n_421),
.Y(n_1761)
);

NAND2xp5_ASAP7_75t_L g1762 ( 
.A(n_1684),
.B(n_145),
.Y(n_1762)
);

AOI21xp5_ASAP7_75t_L g1763 ( 
.A1(n_1629),
.A2(n_423),
.B(n_422),
.Y(n_1763)
);

NAND2xp5_ASAP7_75t_L g1764 ( 
.A(n_1684),
.B(n_148),
.Y(n_1764)
);

BUFx8_ASAP7_75t_SL g1765 ( 
.A(n_1598),
.Y(n_1765)
);

OAI22xp5_ASAP7_75t_L g1766 ( 
.A1(n_1679),
.A2(n_149),
.B1(n_150),
.B2(n_151),
.Y(n_1766)
);

OR2x6_ASAP7_75t_L g1767 ( 
.A(n_1646),
.B(n_424),
.Y(n_1767)
);

INVx2_ASAP7_75t_SL g1768 ( 
.A(n_1680),
.Y(n_1768)
);

INVx4_ASAP7_75t_L g1769 ( 
.A(n_1617),
.Y(n_1769)
);

BUFx6f_ASAP7_75t_L g1770 ( 
.A(n_1598),
.Y(n_1770)
);

BUFx3_ASAP7_75t_L g1771 ( 
.A(n_1680),
.Y(n_1771)
);

NAND2xp5_ASAP7_75t_L g1772 ( 
.A(n_1613),
.B(n_149),
.Y(n_1772)
);

OAI22xp5_ASAP7_75t_L g1773 ( 
.A1(n_1581),
.A2(n_151),
.B1(n_153),
.B2(n_154),
.Y(n_1773)
);

AND2x2_ASAP7_75t_L g1774 ( 
.A(n_1611),
.B(n_425),
.Y(n_1774)
);

AND2x4_ASAP7_75t_L g1775 ( 
.A(n_1630),
.B(n_426),
.Y(n_1775)
);

NAND2x1p5_ASAP7_75t_L g1776 ( 
.A(n_1596),
.B(n_429),
.Y(n_1776)
);

NAND2xp5_ASAP7_75t_L g1777 ( 
.A(n_1608),
.B(n_153),
.Y(n_1777)
);

BUFx5_ASAP7_75t_L g1778 ( 
.A(n_1690),
.Y(n_1778)
);

BUFx3_ASAP7_75t_L g1779 ( 
.A(n_1630),
.Y(n_1779)
);

AND2x2_ASAP7_75t_L g1780 ( 
.A(n_1628),
.B(n_430),
.Y(n_1780)
);

AND2x2_ASAP7_75t_L g1781 ( 
.A(n_1650),
.B(n_431),
.Y(n_1781)
);

INVx4_ASAP7_75t_L g1782 ( 
.A(n_1617),
.Y(n_1782)
);

NAND2xp5_ASAP7_75t_L g1783 ( 
.A(n_1608),
.B(n_1643),
.Y(n_1783)
);

CKINVDCx16_ASAP7_75t_R g1784 ( 
.A(n_1656),
.Y(n_1784)
);

NAND2xp5_ASAP7_75t_L g1785 ( 
.A(n_1608),
.B(n_154),
.Y(n_1785)
);

OAI22xp5_ASAP7_75t_L g1786 ( 
.A1(n_1647),
.A2(n_155),
.B1(n_156),
.B2(n_157),
.Y(n_1786)
);

INVx3_ASAP7_75t_L g1787 ( 
.A(n_1676),
.Y(n_1787)
);

NAND2xp5_ASAP7_75t_SL g1788 ( 
.A(n_1588),
.B(n_432),
.Y(n_1788)
);

AOI21xp33_ASAP7_75t_SL g1789 ( 
.A1(n_1661),
.A2(n_156),
.B(n_158),
.Y(n_1789)
);

NAND2x1p5_ASAP7_75t_L g1790 ( 
.A(n_1596),
.B(n_433),
.Y(n_1790)
);

NAND3xp33_ASAP7_75t_L g1791 ( 
.A(n_1655),
.B(n_158),
.C(n_160),
.Y(n_1791)
);

BUFx12f_ASAP7_75t_L g1792 ( 
.A(n_1687),
.Y(n_1792)
);

BUFx3_ASAP7_75t_L g1793 ( 
.A(n_1765),
.Y(n_1793)
);

OR2x2_ASAP7_75t_L g1794 ( 
.A(n_1706),
.B(n_1675),
.Y(n_1794)
);

AOI21xp5_ASAP7_75t_SL g1795 ( 
.A1(n_1767),
.A2(n_1652),
.B(n_1657),
.Y(n_1795)
);

NAND2xp5_ASAP7_75t_L g1796 ( 
.A(n_1744),
.B(n_1599),
.Y(n_1796)
);

A2O1A1Ixp33_ASAP7_75t_L g1797 ( 
.A1(n_1708),
.A2(n_1659),
.B(n_1641),
.C(n_1696),
.Y(n_1797)
);

A2O1A1Ixp33_ASAP7_75t_SL g1798 ( 
.A1(n_1755),
.A2(n_1580),
.B(n_1649),
.C(n_1695),
.Y(n_1798)
);

NOR2xp33_ASAP7_75t_SL g1799 ( 
.A(n_1716),
.B(n_1596),
.Y(n_1799)
);

HB1xp67_ASAP7_75t_L g1800 ( 
.A(n_1746),
.Y(n_1800)
);

AND2x2_ASAP7_75t_L g1801 ( 
.A(n_1736),
.B(n_1604),
.Y(n_1801)
);

AND2x2_ASAP7_75t_L g1802 ( 
.A(n_1739),
.B(n_1621),
.Y(n_1802)
);

A2O1A1Ixp33_ASAP7_75t_L g1803 ( 
.A1(n_1702),
.A2(n_1673),
.B(n_1639),
.C(n_1636),
.Y(n_1803)
);

INVx2_ASAP7_75t_L g1804 ( 
.A(n_1738),
.Y(n_1804)
);

INVx1_ASAP7_75t_L g1805 ( 
.A(n_1701),
.Y(n_1805)
);

A2O1A1Ixp33_ASAP7_75t_SL g1806 ( 
.A1(n_1763),
.A2(n_1614),
.B(n_1699),
.C(n_1682),
.Y(n_1806)
);

AND2x2_ASAP7_75t_L g1807 ( 
.A(n_1724),
.B(n_1621),
.Y(n_1807)
);

OR2x2_ASAP7_75t_L g1808 ( 
.A(n_1783),
.B(n_1733),
.Y(n_1808)
);

A2O1A1Ixp33_ASAP7_75t_L g1809 ( 
.A1(n_1707),
.A2(n_1622),
.B(n_1700),
.C(n_1640),
.Y(n_1809)
);

NAND2xp5_ASAP7_75t_L g1810 ( 
.A(n_1754),
.B(n_1621),
.Y(n_1810)
);

AND2x2_ASAP7_75t_L g1811 ( 
.A(n_1730),
.B(n_1631),
.Y(n_1811)
);

CKINVDCx5p33_ASAP7_75t_R g1812 ( 
.A(n_1721),
.Y(n_1812)
);

A2O1A1Ixp33_ASAP7_75t_L g1813 ( 
.A1(n_1717),
.A2(n_1642),
.B(n_1637),
.C(n_1626),
.Y(n_1813)
);

AND2x4_ASAP7_75t_L g1814 ( 
.A(n_1753),
.B(n_1631),
.Y(n_1814)
);

BUFx2_ASAP7_75t_L g1815 ( 
.A(n_1747),
.Y(n_1815)
);

NAND2xp5_ASAP7_75t_L g1816 ( 
.A(n_1735),
.B(n_1671),
.Y(n_1816)
);

AND2x2_ASAP7_75t_L g1817 ( 
.A(n_1720),
.B(n_1686),
.Y(n_1817)
);

INVxp67_ASAP7_75t_SL g1818 ( 
.A(n_1777),
.Y(n_1818)
);

OA21x2_ASAP7_75t_L g1819 ( 
.A1(n_1785),
.A2(n_1575),
.B(n_1586),
.Y(n_1819)
);

NAND2xp5_ASAP7_75t_SL g1820 ( 
.A(n_1725),
.B(n_1605),
.Y(n_1820)
);

NAND2xp5_ASAP7_75t_L g1821 ( 
.A(n_1712),
.B(n_1600),
.Y(n_1821)
);

O2A1O1Ixp33_ASAP7_75t_L g1822 ( 
.A1(n_1726),
.A2(n_1651),
.B(n_1623),
.C(n_1638),
.Y(n_1822)
);

BUFx3_ASAP7_75t_L g1823 ( 
.A(n_1751),
.Y(n_1823)
);

NAND2xp5_ASAP7_75t_L g1824 ( 
.A(n_1715),
.B(n_1703),
.Y(n_1824)
);

OR2x2_ASAP7_75t_L g1825 ( 
.A(n_1713),
.B(n_1672),
.Y(n_1825)
);

O2A1O1Ixp33_ASAP7_75t_L g1826 ( 
.A1(n_1737),
.A2(n_1694),
.B(n_1688),
.C(n_1667),
.Y(n_1826)
);

AND2x4_ASAP7_75t_L g1827 ( 
.A(n_1710),
.B(n_1591),
.Y(n_1827)
);

NOR2xp33_ASAP7_75t_L g1828 ( 
.A(n_1748),
.B(n_1624),
.Y(n_1828)
);

INVx1_ASAP7_75t_L g1829 ( 
.A(n_1778),
.Y(n_1829)
);

BUFx2_ASAP7_75t_L g1830 ( 
.A(n_1731),
.Y(n_1830)
);

HB1xp67_ASAP7_75t_L g1831 ( 
.A(n_1778),
.Y(n_1831)
);

AND2x2_ASAP7_75t_L g1832 ( 
.A(n_1743),
.B(n_1681),
.Y(n_1832)
);

NAND2xp5_ASAP7_75t_L g1833 ( 
.A(n_1718),
.B(n_1683),
.Y(n_1833)
);

HB1xp67_ASAP7_75t_L g1834 ( 
.A(n_1778),
.Y(n_1834)
);

OR2x2_ASAP7_75t_L g1835 ( 
.A(n_1732),
.B(n_1762),
.Y(n_1835)
);

AND2x2_ASAP7_75t_L g1836 ( 
.A(n_1784),
.B(n_1645),
.Y(n_1836)
);

INVx2_ASAP7_75t_L g1837 ( 
.A(n_1804),
.Y(n_1837)
);

INVx1_ASAP7_75t_L g1838 ( 
.A(n_1804),
.Y(n_1838)
);

AND2x2_ASAP7_75t_L g1839 ( 
.A(n_1802),
.B(n_1778),
.Y(n_1839)
);

INVx5_ASAP7_75t_L g1840 ( 
.A(n_1827),
.Y(n_1840)
);

AND2x4_ASAP7_75t_L g1841 ( 
.A(n_1829),
.B(n_1711),
.Y(n_1841)
);

INVx1_ASAP7_75t_L g1842 ( 
.A(n_1805),
.Y(n_1842)
);

AND2x2_ASAP7_75t_L g1843 ( 
.A(n_1807),
.B(n_1722),
.Y(n_1843)
);

INVx1_ASAP7_75t_SL g1844 ( 
.A(n_1794),
.Y(n_1844)
);

INVx2_ASAP7_75t_SL g1845 ( 
.A(n_1831),
.Y(n_1845)
);

INVx3_ASAP7_75t_L g1846 ( 
.A(n_1827),
.Y(n_1846)
);

HB1xp67_ASAP7_75t_L g1847 ( 
.A(n_1800),
.Y(n_1847)
);

INVx1_ASAP7_75t_L g1848 ( 
.A(n_1800),
.Y(n_1848)
);

NAND2xp5_ASAP7_75t_L g1849 ( 
.A(n_1818),
.B(n_1709),
.Y(n_1849)
);

OAI21x1_ASAP7_75t_L g1850 ( 
.A1(n_1820),
.A2(n_1760),
.B(n_1601),
.Y(n_1850)
);

HB1xp67_ASAP7_75t_L g1851 ( 
.A(n_1814),
.Y(n_1851)
);

AND2x2_ASAP7_75t_L g1852 ( 
.A(n_1811),
.B(n_1787),
.Y(n_1852)
);

INVx1_ASAP7_75t_L g1853 ( 
.A(n_1810),
.Y(n_1853)
);

HB1xp67_ASAP7_75t_L g1854 ( 
.A(n_1818),
.Y(n_1854)
);

INVx2_ASAP7_75t_SL g1855 ( 
.A(n_1831),
.Y(n_1855)
);

INVx1_ASAP7_75t_L g1856 ( 
.A(n_1808),
.Y(n_1856)
);

INVx2_ASAP7_75t_L g1857 ( 
.A(n_1819),
.Y(n_1857)
);

BUFx3_ASAP7_75t_L g1858 ( 
.A(n_1815),
.Y(n_1858)
);

NOR2xp33_ASAP7_75t_L g1859 ( 
.A(n_1824),
.B(n_1759),
.Y(n_1859)
);

NAND2xp33_ASAP7_75t_SL g1860 ( 
.A(n_1796),
.B(n_1741),
.Y(n_1860)
);

INVx1_ASAP7_75t_L g1861 ( 
.A(n_1837),
.Y(n_1861)
);

AOI22xp33_ASAP7_75t_L g1862 ( 
.A1(n_1860),
.A2(n_1836),
.B1(n_1791),
.B2(n_1766),
.Y(n_1862)
);

BUFx3_ASAP7_75t_L g1863 ( 
.A(n_1858),
.Y(n_1863)
);

INVx2_ASAP7_75t_L g1864 ( 
.A(n_1837),
.Y(n_1864)
);

INVx1_ASAP7_75t_L g1865 ( 
.A(n_1838),
.Y(n_1865)
);

HB1xp67_ASAP7_75t_L g1866 ( 
.A(n_1854),
.Y(n_1866)
);

BUFx2_ASAP7_75t_L g1867 ( 
.A(n_1846),
.Y(n_1867)
);

AND2x2_ASAP7_75t_L g1868 ( 
.A(n_1851),
.B(n_1834),
.Y(n_1868)
);

AND2x2_ASAP7_75t_L g1869 ( 
.A(n_1839),
.B(n_1834),
.Y(n_1869)
);

INVx1_ASAP7_75t_L g1870 ( 
.A(n_1838),
.Y(n_1870)
);

AND2x2_ASAP7_75t_L g1871 ( 
.A(n_1839),
.B(n_1846),
.Y(n_1871)
);

BUFx2_ASAP7_75t_L g1872 ( 
.A(n_1846),
.Y(n_1872)
);

NAND2xp5_ASAP7_75t_L g1873 ( 
.A(n_1844),
.B(n_1814),
.Y(n_1873)
);

INVx1_ASAP7_75t_L g1874 ( 
.A(n_1854),
.Y(n_1874)
);

AND2x2_ASAP7_75t_L g1875 ( 
.A(n_1846),
.B(n_1852),
.Y(n_1875)
);

INVx2_ASAP7_75t_L g1876 ( 
.A(n_1857),
.Y(n_1876)
);

AND2x2_ASAP7_75t_L g1877 ( 
.A(n_1844),
.B(n_1801),
.Y(n_1877)
);

INVx3_ASAP7_75t_L g1878 ( 
.A(n_1840),
.Y(n_1878)
);

OAI22xp5_ASAP7_75t_L g1879 ( 
.A1(n_1858),
.A2(n_1797),
.B1(n_1803),
.B2(n_1835),
.Y(n_1879)
);

OR2x2_ASAP7_75t_L g1880 ( 
.A(n_1847),
.B(n_1825),
.Y(n_1880)
);

INVx2_ASAP7_75t_L g1881 ( 
.A(n_1857),
.Y(n_1881)
);

INVx1_ASAP7_75t_L g1882 ( 
.A(n_1865),
.Y(n_1882)
);

NAND2xp5_ASAP7_75t_L g1883 ( 
.A(n_1880),
.B(n_1856),
.Y(n_1883)
);

INVx1_ASAP7_75t_L g1884 ( 
.A(n_1865),
.Y(n_1884)
);

BUFx3_ASAP7_75t_L g1885 ( 
.A(n_1863),
.Y(n_1885)
);

INVx1_ASAP7_75t_L g1886 ( 
.A(n_1870),
.Y(n_1886)
);

HB1xp67_ASAP7_75t_L g1887 ( 
.A(n_1866),
.Y(n_1887)
);

HB1xp67_ASAP7_75t_L g1888 ( 
.A(n_1874),
.Y(n_1888)
);

INVx1_ASAP7_75t_L g1889 ( 
.A(n_1870),
.Y(n_1889)
);

AND2x2_ASAP7_75t_L g1890 ( 
.A(n_1871),
.B(n_1840),
.Y(n_1890)
);

AND2x2_ASAP7_75t_L g1891 ( 
.A(n_1871),
.B(n_1840),
.Y(n_1891)
);

BUFx3_ASAP7_75t_L g1892 ( 
.A(n_1863),
.Y(n_1892)
);

INVx1_ASAP7_75t_L g1893 ( 
.A(n_1874),
.Y(n_1893)
);

INVx2_ASAP7_75t_L g1894 ( 
.A(n_1885),
.Y(n_1894)
);

INVx1_ASAP7_75t_SL g1895 ( 
.A(n_1885),
.Y(n_1895)
);

INVx1_ASAP7_75t_L g1896 ( 
.A(n_1884),
.Y(n_1896)
);

OR2x2_ASAP7_75t_L g1897 ( 
.A(n_1883),
.B(n_1880),
.Y(n_1897)
);

AND2x4_ASAP7_75t_L g1898 ( 
.A(n_1892),
.B(n_1863),
.Y(n_1898)
);

OAI22xp5_ASAP7_75t_L g1899 ( 
.A1(n_1892),
.A2(n_1862),
.B1(n_1879),
.B2(n_1858),
.Y(n_1899)
);

INVx1_ASAP7_75t_SL g1900 ( 
.A(n_1895),
.Y(n_1900)
);

OR2x2_ASAP7_75t_L g1901 ( 
.A(n_1897),
.B(n_1887),
.Y(n_1901)
);

AND2x2_ASAP7_75t_L g1902 ( 
.A(n_1898),
.B(n_1890),
.Y(n_1902)
);

AND2x2_ASAP7_75t_L g1903 ( 
.A(n_1894),
.B(n_1890),
.Y(n_1903)
);

INVx1_ASAP7_75t_L g1904 ( 
.A(n_1896),
.Y(n_1904)
);

INVx2_ASAP7_75t_L g1905 ( 
.A(n_1898),
.Y(n_1905)
);

INVx1_ASAP7_75t_L g1906 ( 
.A(n_1899),
.Y(n_1906)
);

AOI22xp33_ASAP7_75t_L g1907 ( 
.A1(n_1899),
.A2(n_1786),
.B1(n_1773),
.B2(n_1828),
.Y(n_1907)
);

INVx1_ASAP7_75t_L g1908 ( 
.A(n_1896),
.Y(n_1908)
);

NAND3xp33_ASAP7_75t_SL g1909 ( 
.A(n_1899),
.B(n_1799),
.C(n_1849),
.Y(n_1909)
);

AND2x4_ASAP7_75t_L g1910 ( 
.A(n_1905),
.B(n_1793),
.Y(n_1910)
);

OR2x2_ASAP7_75t_L g1911 ( 
.A(n_1900),
.B(n_1873),
.Y(n_1911)
);

AND2x2_ASAP7_75t_L g1912 ( 
.A(n_1902),
.B(n_1891),
.Y(n_1912)
);

AND2x2_ASAP7_75t_L g1913 ( 
.A(n_1902),
.B(n_1891),
.Y(n_1913)
);

INVx1_ASAP7_75t_L g1914 ( 
.A(n_1904),
.Y(n_1914)
);

INVx2_ASAP7_75t_L g1915 ( 
.A(n_1905),
.Y(n_1915)
);

INVx1_ASAP7_75t_L g1916 ( 
.A(n_1908),
.Y(n_1916)
);

INVx2_ASAP7_75t_L g1917 ( 
.A(n_1903),
.Y(n_1917)
);

NAND2xp5_ASAP7_75t_L g1918 ( 
.A(n_1906),
.B(n_1888),
.Y(n_1918)
);

INVx1_ASAP7_75t_L g1919 ( 
.A(n_1901),
.Y(n_1919)
);

INVx1_ASAP7_75t_L g1920 ( 
.A(n_1909),
.Y(n_1920)
);

OAI21xp33_ASAP7_75t_L g1921 ( 
.A1(n_1920),
.A2(n_1907),
.B(n_1849),
.Y(n_1921)
);

AND2x2_ASAP7_75t_L g1922 ( 
.A(n_1910),
.B(n_1793),
.Y(n_1922)
);

INVx1_ASAP7_75t_L g1923 ( 
.A(n_1915),
.Y(n_1923)
);

INVx1_ASAP7_75t_L g1924 ( 
.A(n_1915),
.Y(n_1924)
);

INVx1_ASAP7_75t_L g1925 ( 
.A(n_1919),
.Y(n_1925)
);

INVx1_ASAP7_75t_L g1926 ( 
.A(n_1914),
.Y(n_1926)
);

NAND2xp5_ASAP7_75t_L g1927 ( 
.A(n_1917),
.B(n_1907),
.Y(n_1927)
);

NAND2xp5_ASAP7_75t_L g1928 ( 
.A(n_1918),
.B(n_1893),
.Y(n_1928)
);

INVx1_ASAP7_75t_L g1929 ( 
.A(n_1923),
.Y(n_1929)
);

NOR3xp33_ASAP7_75t_L g1930 ( 
.A(n_1927),
.B(n_1918),
.C(n_1916),
.Y(n_1930)
);

AND2x2_ASAP7_75t_L g1931 ( 
.A(n_1922),
.B(n_1910),
.Y(n_1931)
);

NAND2xp5_ASAP7_75t_L g1932 ( 
.A(n_1925),
.B(n_1917),
.Y(n_1932)
);

OAI22xp5_ASAP7_75t_L g1933 ( 
.A1(n_1930),
.A2(n_1911),
.B1(n_1921),
.B2(n_1928),
.Y(n_1933)
);

INVx1_ASAP7_75t_L g1934 ( 
.A(n_1932),
.Y(n_1934)
);

AND2x2_ASAP7_75t_L g1935 ( 
.A(n_1931),
.B(n_1912),
.Y(n_1935)
);

INVx1_ASAP7_75t_L g1936 ( 
.A(n_1929),
.Y(n_1936)
);

INVx1_ASAP7_75t_L g1937 ( 
.A(n_1934),
.Y(n_1937)
);

AOI32xp33_ASAP7_75t_L g1938 ( 
.A1(n_1933),
.A2(n_1935),
.A3(n_1926),
.B1(n_1924),
.B2(n_1936),
.Y(n_1938)
);

AND2x2_ASAP7_75t_L g1939 ( 
.A(n_1935),
.B(n_1913),
.Y(n_1939)
);

NOR2x1_ASAP7_75t_L g1940 ( 
.A(n_1934),
.B(n_1928),
.Y(n_1940)
);

INVx2_ASAP7_75t_L g1941 ( 
.A(n_1935),
.Y(n_1941)
);

AND2x2_ASAP7_75t_L g1942 ( 
.A(n_1939),
.B(n_1812),
.Y(n_1942)
);

NAND2xp5_ASAP7_75t_L g1943 ( 
.A(n_1941),
.B(n_1859),
.Y(n_1943)
);

INVx1_ASAP7_75t_L g1944 ( 
.A(n_1940),
.Y(n_1944)
);

INVx2_ASAP7_75t_L g1945 ( 
.A(n_1937),
.Y(n_1945)
);

INVx1_ASAP7_75t_L g1946 ( 
.A(n_1938),
.Y(n_1946)
);

INVx2_ASAP7_75t_L g1947 ( 
.A(n_1939),
.Y(n_1947)
);

NAND2xp5_ASAP7_75t_L g1948 ( 
.A(n_1939),
.B(n_1882),
.Y(n_1948)
);

NAND2xp5_ASAP7_75t_L g1949 ( 
.A(n_1939),
.B(n_1884),
.Y(n_1949)
);

INVx1_ASAP7_75t_L g1950 ( 
.A(n_1941),
.Y(n_1950)
);

NAND2xp5_ASAP7_75t_L g1951 ( 
.A(n_1941),
.B(n_1886),
.Y(n_1951)
);

INVxp67_ASAP7_75t_SL g1952 ( 
.A(n_1944),
.Y(n_1952)
);

HB1xp67_ASAP7_75t_L g1953 ( 
.A(n_1947),
.Y(n_1953)
);

AND3x1_ASAP7_75t_L g1954 ( 
.A(n_1946),
.B(n_1772),
.C(n_1768),
.Y(n_1954)
);

OR2x2_ASAP7_75t_L g1955 ( 
.A(n_1950),
.B(n_1943),
.Y(n_1955)
);

INVx1_ASAP7_75t_L g1956 ( 
.A(n_1951),
.Y(n_1956)
);

INVx1_ASAP7_75t_SL g1957 ( 
.A(n_1942),
.Y(n_1957)
);

NAND2xp5_ASAP7_75t_L g1958 ( 
.A(n_1945),
.B(n_1889),
.Y(n_1958)
);

INVx2_ASAP7_75t_L g1959 ( 
.A(n_1949),
.Y(n_1959)
);

INVxp67_ASAP7_75t_SL g1960 ( 
.A(n_1951),
.Y(n_1960)
);

INVx3_ASAP7_75t_L g1961 ( 
.A(n_1948),
.Y(n_1961)
);

AND2x2_ASAP7_75t_L g1962 ( 
.A(n_1942),
.B(n_1727),
.Y(n_1962)
);

INVx1_ASAP7_75t_L g1963 ( 
.A(n_1944),
.Y(n_1963)
);

AND2x2_ASAP7_75t_L g1964 ( 
.A(n_1942),
.B(n_1723),
.Y(n_1964)
);

BUFx2_ASAP7_75t_L g1965 ( 
.A(n_1953),
.Y(n_1965)
);

NAND2xp5_ASAP7_75t_L g1966 ( 
.A(n_1957),
.B(n_1886),
.Y(n_1966)
);

NOR3xp33_ASAP7_75t_L g1967 ( 
.A(n_1957),
.B(n_1789),
.C(n_1745),
.Y(n_1967)
);

AOI211xp5_ASAP7_75t_L g1968 ( 
.A1(n_1963),
.A2(n_1719),
.B(n_1771),
.C(n_1729),
.Y(n_1968)
);

NAND2xp5_ASAP7_75t_L g1969 ( 
.A(n_1952),
.B(n_1889),
.Y(n_1969)
);

NOR2xp33_ASAP7_75t_SL g1970 ( 
.A(n_1955),
.B(n_1749),
.Y(n_1970)
);

INVx1_ASAP7_75t_L g1971 ( 
.A(n_1954),
.Y(n_1971)
);

NAND3xp33_ASAP7_75t_L g1972 ( 
.A(n_1959),
.B(n_1757),
.C(n_1764),
.Y(n_1972)
);

O2A1O1Ixp33_ASAP7_75t_SL g1973 ( 
.A1(n_1958),
.A2(n_1742),
.B(n_1833),
.C(n_1816),
.Y(n_1973)
);

NAND4xp25_ASAP7_75t_L g1974 ( 
.A(n_1962),
.B(n_1830),
.C(n_1826),
.D(n_1822),
.Y(n_1974)
);

INVx1_ASAP7_75t_L g1975 ( 
.A(n_1960),
.Y(n_1975)
);

NAND2xp5_ASAP7_75t_L g1976 ( 
.A(n_1961),
.B(n_1867),
.Y(n_1976)
);

INVx1_ASAP7_75t_L g1977 ( 
.A(n_1958),
.Y(n_1977)
);

NAND3xp33_ASAP7_75t_SL g1978 ( 
.A(n_1965),
.B(n_1956),
.C(n_1964),
.Y(n_1978)
);

NOR2x1_ASAP7_75t_L g1979 ( 
.A(n_1975),
.B(n_1961),
.Y(n_1979)
);

OR3x1_ASAP7_75t_L g1980 ( 
.A(n_1971),
.B(n_1752),
.C(n_1828),
.Y(n_1980)
);

NOR2xp67_ASAP7_75t_L g1981 ( 
.A(n_1976),
.B(n_160),
.Y(n_1981)
);

NOR3xp33_ASAP7_75t_L g1982 ( 
.A(n_1977),
.B(n_1774),
.C(n_1780),
.Y(n_1982)
);

OAI221xp5_ASAP7_75t_L g1983 ( 
.A1(n_1970),
.A2(n_1790),
.B1(n_1776),
.B2(n_1767),
.C(n_1878),
.Y(n_1983)
);

NOR3x1_ASAP7_75t_L g1984 ( 
.A(n_1969),
.B(n_1872),
.C(n_1867),
.Y(n_1984)
);

HB1xp67_ASAP7_75t_L g1985 ( 
.A(n_1966),
.Y(n_1985)
);

AOI221xp5_ASAP7_75t_L g1986 ( 
.A1(n_1967),
.A2(n_1878),
.B1(n_1781),
.B2(n_1761),
.C(n_1788),
.Y(n_1986)
);

AND2x2_ASAP7_75t_SL g1987 ( 
.A(n_1968),
.B(n_1758),
.Y(n_1987)
);

NAND3xp33_ASAP7_75t_L g1988 ( 
.A(n_1972),
.B(n_1973),
.C(n_1974),
.Y(n_1988)
);

NAND4xp25_ASAP7_75t_L g1989 ( 
.A(n_1970),
.B(n_1758),
.C(n_1795),
.D(n_1832),
.Y(n_1989)
);

NAND2xp5_ASAP7_75t_L g1990 ( 
.A(n_1981),
.B(n_1792),
.Y(n_1990)
);

AND2x4_ASAP7_75t_L g1991 ( 
.A(n_1979),
.B(n_1878),
.Y(n_1991)
);

INVx1_ASAP7_75t_L g1992 ( 
.A(n_1985),
.Y(n_1992)
);

NOR3xp33_ASAP7_75t_L g1993 ( 
.A(n_1978),
.B(n_1988),
.C(n_1989),
.Y(n_1993)
);

AOI211xp5_ASAP7_75t_L g1994 ( 
.A1(n_1986),
.A2(n_1728),
.B(n_1705),
.C(n_163),
.Y(n_1994)
);

INVx1_ASAP7_75t_L g1995 ( 
.A(n_1980),
.Y(n_1995)
);

O2A1O1Ixp33_ASAP7_75t_L g1996 ( 
.A1(n_1982),
.A2(n_164),
.B(n_161),
.C(n_162),
.Y(n_1996)
);

NAND3xp33_ASAP7_75t_L g1997 ( 
.A(n_1987),
.B(n_1983),
.C(n_1984),
.Y(n_1997)
);

NAND2xp5_ASAP7_75t_SL g1998 ( 
.A(n_1981),
.B(n_1705),
.Y(n_1998)
);

INVx1_ASAP7_75t_L g1999 ( 
.A(n_1979),
.Y(n_1999)
);

INVx1_ASAP7_75t_L g2000 ( 
.A(n_1979),
.Y(n_2000)
);

NAND3xp33_ASAP7_75t_L g2001 ( 
.A(n_1979),
.B(n_1728),
.C(n_1705),
.Y(n_2001)
);

INVx2_ASAP7_75t_SL g2002 ( 
.A(n_1979),
.Y(n_2002)
);

NAND2xp5_ASAP7_75t_SL g2003 ( 
.A(n_1981),
.B(n_1728),
.Y(n_2003)
);

AOI22xp5_ASAP7_75t_L g2004 ( 
.A1(n_1978),
.A2(n_1878),
.B1(n_1872),
.B2(n_1868),
.Y(n_2004)
);

INVx1_ASAP7_75t_SL g2005 ( 
.A(n_1979),
.Y(n_2005)
);

OR2x2_ASAP7_75t_L g2006 ( 
.A(n_2002),
.B(n_161),
.Y(n_2006)
);

INVx1_ASAP7_75t_L g2007 ( 
.A(n_1999),
.Y(n_2007)
);

AOI21xp33_ASAP7_75t_SL g2008 ( 
.A1(n_2000),
.A2(n_162),
.B(n_165),
.Y(n_2008)
);

NOR2x1_ASAP7_75t_L g2009 ( 
.A(n_2005),
.B(n_165),
.Y(n_2009)
);

NOR2x1_ASAP7_75t_L g2010 ( 
.A(n_1992),
.B(n_2001),
.Y(n_2010)
);

NOR2x1_ASAP7_75t_L g2011 ( 
.A(n_1998),
.B(n_166),
.Y(n_2011)
);

NOR2xp33_ASAP7_75t_L g2012 ( 
.A(n_2003),
.B(n_1990),
.Y(n_2012)
);

INVx2_ASAP7_75t_L g2013 ( 
.A(n_1991),
.Y(n_2013)
);

NOR3x2_ASAP7_75t_L g2014 ( 
.A(n_1993),
.B(n_167),
.C(n_168),
.Y(n_2014)
);

AND2x2_ASAP7_75t_SL g2015 ( 
.A(n_1995),
.B(n_1775),
.Y(n_2015)
);

NOR3xp33_ASAP7_75t_L g2016 ( 
.A(n_1997),
.B(n_1782),
.C(n_1769),
.Y(n_2016)
);

AND2x2_ASAP7_75t_L g2017 ( 
.A(n_2004),
.B(n_1877),
.Y(n_2017)
);

INVx1_ASAP7_75t_L g2018 ( 
.A(n_1996),
.Y(n_2018)
);

NOR2x1_ASAP7_75t_L g2019 ( 
.A(n_1994),
.B(n_168),
.Y(n_2019)
);

NOR2xp33_ASAP7_75t_L g2020 ( 
.A(n_2005),
.B(n_169),
.Y(n_2020)
);

NAND3xp33_ASAP7_75t_L g2021 ( 
.A(n_1993),
.B(n_1710),
.C(n_169),
.Y(n_2021)
);

AND2x4_ASAP7_75t_L g2022 ( 
.A(n_2002),
.B(n_1710),
.Y(n_2022)
);

NOR3xp33_ASAP7_75t_L g2023 ( 
.A(n_1993),
.B(n_1782),
.C(n_1769),
.Y(n_2023)
);

NAND4xp75_ASAP7_75t_L g2024 ( 
.A(n_2002),
.B(n_170),
.C(n_171),
.D(n_173),
.Y(n_2024)
);

OR2x2_ASAP7_75t_L g2025 ( 
.A(n_2002),
.B(n_170),
.Y(n_2025)
);

NAND2xp5_ASAP7_75t_L g2026 ( 
.A(n_1991),
.B(n_171),
.Y(n_2026)
);

INVx1_ASAP7_75t_L g2027 ( 
.A(n_2002),
.Y(n_2027)
);

NOR3xp33_ASAP7_75t_SL g2028 ( 
.A(n_1999),
.B(n_173),
.C(n_174),
.Y(n_2028)
);

NOR2xp33_ASAP7_75t_L g2029 ( 
.A(n_2005),
.B(n_174),
.Y(n_2029)
);

NAND2xp5_ASAP7_75t_SL g2030 ( 
.A(n_2002),
.B(n_1751),
.Y(n_2030)
);

OAI21xp5_ASAP7_75t_SL g2031 ( 
.A1(n_2004),
.A2(n_1664),
.B(n_1775),
.Y(n_2031)
);

INVx1_ASAP7_75t_L g2032 ( 
.A(n_2002),
.Y(n_2032)
);

NAND2xp5_ASAP7_75t_L g2033 ( 
.A(n_2022),
.B(n_175),
.Y(n_2033)
);

AOI21xp5_ASAP7_75t_L g2034 ( 
.A1(n_2027),
.A2(n_1803),
.B(n_1693),
.Y(n_2034)
);

INVx1_ASAP7_75t_L g2035 ( 
.A(n_2009),
.Y(n_2035)
);

NOR3x2_ASAP7_75t_L g2036 ( 
.A(n_2024),
.B(n_176),
.C(n_177),
.Y(n_2036)
);

OAI21xp5_ASAP7_75t_L g2037 ( 
.A1(n_2021),
.A2(n_1618),
.B(n_1607),
.Y(n_2037)
);

NAND2x1p5_ASAP7_75t_L g2038 ( 
.A(n_2011),
.B(n_1751),
.Y(n_2038)
);

INVx2_ASAP7_75t_L g2039 ( 
.A(n_2006),
.Y(n_2039)
);

NOR2x1_ASAP7_75t_L g2040 ( 
.A(n_2025),
.B(n_176),
.Y(n_2040)
);

BUFx6f_ASAP7_75t_L g2041 ( 
.A(n_2032),
.Y(n_2041)
);

NAND5xp2_ASAP7_75t_L g2042 ( 
.A(n_2023),
.B(n_1740),
.C(n_1750),
.D(n_179),
.E(n_180),
.Y(n_2042)
);

AND3x4_ASAP7_75t_L g2043 ( 
.A(n_2016),
.B(n_1823),
.C(n_1779),
.Y(n_2043)
);

NAND2xp5_ASAP7_75t_L g2044 ( 
.A(n_2022),
.B(n_177),
.Y(n_2044)
);

AO22x2_ASAP7_75t_L g2045 ( 
.A1(n_2013),
.A2(n_1881),
.B1(n_1876),
.B2(n_1704),
.Y(n_2045)
);

NAND3xp33_ASAP7_75t_L g2046 ( 
.A(n_2028),
.B(n_178),
.C(n_179),
.Y(n_2046)
);

OAI221xp5_ASAP7_75t_L g2047 ( 
.A1(n_2007),
.A2(n_1798),
.B1(n_1809),
.B2(n_1797),
.C(n_1734),
.Y(n_2047)
);

NOR2x1_ASAP7_75t_L g2048 ( 
.A(n_2010),
.B(n_178),
.Y(n_2048)
);

OAI211xp5_ASAP7_75t_SL g2049 ( 
.A1(n_2018),
.A2(n_180),
.B(n_181),
.C(n_182),
.Y(n_2049)
);

INVx2_ASAP7_75t_L g2050 ( 
.A(n_2014),
.Y(n_2050)
);

NAND2x1p5_ASAP7_75t_L g2051 ( 
.A(n_2030),
.B(n_1770),
.Y(n_2051)
);

OAI311xp33_ASAP7_75t_L g2052 ( 
.A1(n_2026),
.A2(n_181),
.A3(n_183),
.B1(n_184),
.C1(n_185),
.Y(n_2052)
);

NAND2x1p5_ASAP7_75t_L g2053 ( 
.A(n_2019),
.B(n_1770),
.Y(n_2053)
);

NAND2xp5_ASAP7_75t_L g2054 ( 
.A(n_2008),
.B(n_183),
.Y(n_2054)
);

INVx1_ASAP7_75t_L g2055 ( 
.A(n_2048),
.Y(n_2055)
);

NAND2xp5_ASAP7_75t_L g2056 ( 
.A(n_2035),
.B(n_2020),
.Y(n_2056)
);

INVx1_ASAP7_75t_L g2057 ( 
.A(n_2040),
.Y(n_2057)
);

OR2x6_ASAP7_75t_L g2058 ( 
.A(n_2050),
.B(n_2029),
.Y(n_2058)
);

INVx2_ASAP7_75t_L g2059 ( 
.A(n_2041),
.Y(n_2059)
);

INVx1_ASAP7_75t_L g2060 ( 
.A(n_2033),
.Y(n_2060)
);

NAND2xp5_ASAP7_75t_L g2061 ( 
.A(n_2041),
.B(n_2015),
.Y(n_2061)
);

INVx1_ASAP7_75t_L g2062 ( 
.A(n_2044),
.Y(n_2062)
);

INVxp67_ASAP7_75t_L g2063 ( 
.A(n_2054),
.Y(n_2063)
);

INVx2_ASAP7_75t_L g2064 ( 
.A(n_2036),
.Y(n_2064)
);

AOI22xp5_ASAP7_75t_L g2065 ( 
.A1(n_2043),
.A2(n_2012),
.B1(n_2017),
.B2(n_2031),
.Y(n_2065)
);

AOI22xp5_ASAP7_75t_L g2066 ( 
.A1(n_2046),
.A2(n_1868),
.B1(n_1877),
.B2(n_1875),
.Y(n_2066)
);

HB1xp67_ASAP7_75t_L g2067 ( 
.A(n_2038),
.Y(n_2067)
);

INVx2_ASAP7_75t_L g2068 ( 
.A(n_2053),
.Y(n_2068)
);

NOR2xp33_ASAP7_75t_L g2069 ( 
.A(n_2049),
.B(n_184),
.Y(n_2069)
);

NAND2xp5_ASAP7_75t_L g2070 ( 
.A(n_2039),
.B(n_2051),
.Y(n_2070)
);

INVx2_ASAP7_75t_L g2071 ( 
.A(n_2045),
.Y(n_2071)
);

NAND2xp5_ASAP7_75t_L g2072 ( 
.A(n_2034),
.B(n_186),
.Y(n_2072)
);

NOR2xp67_ASAP7_75t_L g2073 ( 
.A(n_2042),
.B(n_186),
.Y(n_2073)
);

INVx2_ASAP7_75t_L g2074 ( 
.A(n_2037),
.Y(n_2074)
);

AND2x2_ASAP7_75t_L g2075 ( 
.A(n_2052),
.B(n_1875),
.Y(n_2075)
);

INVx3_ASAP7_75t_L g2076 ( 
.A(n_2047),
.Y(n_2076)
);

INVx1_ASAP7_75t_L g2077 ( 
.A(n_2048),
.Y(n_2077)
);

INVx1_ASAP7_75t_L g2078 ( 
.A(n_2048),
.Y(n_2078)
);

OR2x2_ASAP7_75t_L g2079 ( 
.A(n_2057),
.B(n_2055),
.Y(n_2079)
);

AND4x1_ASAP7_75t_L g2080 ( 
.A(n_2061),
.B(n_187),
.C(n_188),
.D(n_189),
.Y(n_2080)
);

AO22x2_ASAP7_75t_L g2081 ( 
.A1(n_2077),
.A2(n_2078),
.B1(n_2059),
.B2(n_2064),
.Y(n_2081)
);

INVx1_ASAP7_75t_L g2082 ( 
.A(n_2075),
.Y(n_2082)
);

OAI221xp5_ASAP7_75t_L g2083 ( 
.A1(n_2065),
.A2(n_187),
.B1(n_188),
.B2(n_189),
.C(n_190),
.Y(n_2083)
);

OAI21x1_ASAP7_75t_L g2084 ( 
.A1(n_2056),
.A2(n_1620),
.B(n_1648),
.Y(n_2084)
);

AND2x4_ASAP7_75t_L g2085 ( 
.A(n_2058),
.B(n_1823),
.Y(n_2085)
);

AOI21xp5_ASAP7_75t_L g2086 ( 
.A1(n_2070),
.A2(n_191),
.B(n_192),
.Y(n_2086)
);

XNOR2x1_ASAP7_75t_L g2087 ( 
.A(n_2073),
.B(n_191),
.Y(n_2087)
);

NAND2xp5_ASAP7_75t_L g2088 ( 
.A(n_2069),
.B(n_192),
.Y(n_2088)
);

XNOR2x1_ASAP7_75t_L g2089 ( 
.A(n_2058),
.B(n_193),
.Y(n_2089)
);

AOI22xp33_ASAP7_75t_SL g2090 ( 
.A1(n_2067),
.A2(n_1756),
.B1(n_1770),
.B2(n_1693),
.Y(n_2090)
);

AOI22xp5_ASAP7_75t_L g2091 ( 
.A1(n_2060),
.A2(n_1817),
.B1(n_1869),
.B2(n_1848),
.Y(n_2091)
);

OA22x2_ASAP7_75t_L g2092 ( 
.A1(n_2068),
.A2(n_1881),
.B1(n_1876),
.B2(n_1855),
.Y(n_2092)
);

OAI22xp5_ASAP7_75t_L g2093 ( 
.A1(n_2063),
.A2(n_2066),
.B1(n_2062),
.B2(n_2071),
.Y(n_2093)
);

INVx2_ASAP7_75t_L g2094 ( 
.A(n_2072),
.Y(n_2094)
);

BUFx6f_ASAP7_75t_L g2095 ( 
.A(n_2076),
.Y(n_2095)
);

AOI22xp5_ASAP7_75t_L g2096 ( 
.A1(n_2074),
.A2(n_1869),
.B1(n_1848),
.B2(n_1845),
.Y(n_2096)
);

INVx3_ASAP7_75t_L g2097 ( 
.A(n_2055),
.Y(n_2097)
);

BUFx2_ASAP7_75t_L g2098 ( 
.A(n_2055),
.Y(n_2098)
);

OAI22xp5_ASAP7_75t_L g2099 ( 
.A1(n_2082),
.A2(n_1881),
.B1(n_1876),
.B2(n_1847),
.Y(n_2099)
);

OR2x2_ASAP7_75t_L g2100 ( 
.A(n_2089),
.B(n_193),
.Y(n_2100)
);

AOI221xp5_ASAP7_75t_L g2101 ( 
.A1(n_2093),
.A2(n_2081),
.B1(n_2098),
.B2(n_2097),
.C(n_2085),
.Y(n_2101)
);

OAI21xp5_ASAP7_75t_L g2102 ( 
.A1(n_2087),
.A2(n_1663),
.B(n_1850),
.Y(n_2102)
);

NOR2xp33_ASAP7_75t_L g2103 ( 
.A(n_2080),
.B(n_194),
.Y(n_2103)
);

NAND4xp75_ASAP7_75t_L g2104 ( 
.A(n_2088),
.B(n_194),
.C(n_195),
.D(n_196),
.Y(n_2104)
);

INVx1_ASAP7_75t_L g2105 ( 
.A(n_2079),
.Y(n_2105)
);

NOR2xp33_ASAP7_75t_L g2106 ( 
.A(n_2083),
.B(n_195),
.Y(n_2106)
);

INVx1_ASAP7_75t_L g2107 ( 
.A(n_2086),
.Y(n_2107)
);

NAND2xp5_ASAP7_75t_L g2108 ( 
.A(n_2094),
.B(n_196),
.Y(n_2108)
);

INVx1_ASAP7_75t_L g2109 ( 
.A(n_2095),
.Y(n_2109)
);

AOI21xp33_ASAP7_75t_SL g2110 ( 
.A1(n_2092),
.A2(n_197),
.B(n_199),
.Y(n_2110)
);

NAND4xp75_ASAP7_75t_L g2111 ( 
.A(n_2095),
.B(n_197),
.C(n_199),
.D(n_200),
.Y(n_2111)
);

AND2x4_ASAP7_75t_L g2112 ( 
.A(n_2091),
.B(n_200),
.Y(n_2112)
);

OAI22xp5_ASAP7_75t_L g2113 ( 
.A1(n_2096),
.A2(n_1855),
.B1(n_1845),
.B2(n_1840),
.Y(n_2113)
);

OAI221xp5_ASAP7_75t_L g2114 ( 
.A1(n_2090),
.A2(n_201),
.B1(n_202),
.B2(n_203),
.C(n_204),
.Y(n_2114)
);

OAI31xp33_ASAP7_75t_SL g2115 ( 
.A1(n_2084),
.A2(n_201),
.A3(n_202),
.B(n_205),
.Y(n_2115)
);

NAND3xp33_ASAP7_75t_SL g2116 ( 
.A(n_2098),
.B(n_205),
.C(n_206),
.Y(n_2116)
);

NAND2x1p5_ASAP7_75t_SL g2117 ( 
.A(n_2094),
.B(n_207),
.Y(n_2117)
);

O2A1O1Ixp33_ASAP7_75t_L g2118 ( 
.A1(n_2082),
.A2(n_207),
.B(n_208),
.C(n_209),
.Y(n_2118)
);

NOR3xp33_ASAP7_75t_L g2119 ( 
.A(n_2101),
.B(n_208),
.C(n_209),
.Y(n_2119)
);

OAI221xp5_ASAP7_75t_L g2120 ( 
.A1(n_2115),
.A2(n_210),
.B1(n_211),
.B2(n_212),
.C(n_213),
.Y(n_2120)
);

NAND2xp5_ASAP7_75t_L g2121 ( 
.A(n_2103),
.B(n_211),
.Y(n_2121)
);

NOR4xp75_ASAP7_75t_L g2122 ( 
.A(n_2116),
.B(n_212),
.C(n_213),
.D(n_214),
.Y(n_2122)
);

NOR2x2_ASAP7_75t_L g2123 ( 
.A(n_2104),
.B(n_214),
.Y(n_2123)
);

NAND3xp33_ASAP7_75t_L g2124 ( 
.A(n_2105),
.B(n_215),
.C(n_216),
.Y(n_2124)
);

AOI222xp33_ASAP7_75t_L g2125 ( 
.A1(n_2109),
.A2(n_215),
.B1(n_216),
.B2(n_217),
.C1(n_218),
.C2(n_219),
.Y(n_2125)
);

AOI221xp5_ASAP7_75t_L g2126 ( 
.A1(n_2110),
.A2(n_217),
.B1(n_218),
.B2(n_219),
.C(n_220),
.Y(n_2126)
);

AOI31xp33_ASAP7_75t_L g2127 ( 
.A1(n_2100),
.A2(n_220),
.A3(n_222),
.B(n_223),
.Y(n_2127)
);

OAI222xp33_ASAP7_75t_L g2128 ( 
.A1(n_2114),
.A2(n_222),
.B1(n_223),
.B2(n_224),
.C1(n_225),
.C2(n_1845),
.Y(n_2128)
);

AOI221xp5_ASAP7_75t_L g2129 ( 
.A1(n_2117),
.A2(n_224),
.B1(n_225),
.B2(n_1855),
.C(n_1861),
.Y(n_2129)
);

NAND5xp2_ASAP7_75t_L g2130 ( 
.A(n_2106),
.B(n_1809),
.C(n_1843),
.D(n_436),
.E(n_437),
.Y(n_2130)
);

NOR3xp33_ASAP7_75t_L g2131 ( 
.A(n_2107),
.B(n_434),
.C(n_435),
.Y(n_2131)
);

AOI22xp5_ASAP7_75t_L g2132 ( 
.A1(n_2112),
.A2(n_1841),
.B1(n_1843),
.B2(n_1856),
.Y(n_2132)
);

NOR3xp33_ASAP7_75t_L g2133 ( 
.A(n_2118),
.B(n_438),
.C(n_440),
.Y(n_2133)
);

BUFx2_ASAP7_75t_SL g2134 ( 
.A(n_2123),
.Y(n_2134)
);

NAND2xp5_ASAP7_75t_L g2135 ( 
.A(n_2127),
.B(n_2112),
.Y(n_2135)
);

NAND2x1p5_ASAP7_75t_L g2136 ( 
.A(n_2121),
.B(n_2108),
.Y(n_2136)
);

INVx1_ASAP7_75t_L g2137 ( 
.A(n_2122),
.Y(n_2137)
);

OAI22x1_ASAP7_75t_L g2138 ( 
.A1(n_2124),
.A2(n_2111),
.B1(n_2113),
.B2(n_2102),
.Y(n_2138)
);

INVx1_ASAP7_75t_L g2139 ( 
.A(n_2120),
.Y(n_2139)
);

AO22x2_ASAP7_75t_L g2140 ( 
.A1(n_2119),
.A2(n_2099),
.B1(n_1861),
.B2(n_1864),
.Y(n_2140)
);

INVx1_ASAP7_75t_L g2141 ( 
.A(n_2126),
.Y(n_2141)
);

INVx1_ASAP7_75t_L g2142 ( 
.A(n_2133),
.Y(n_2142)
);

OA22x2_ASAP7_75t_L g2143 ( 
.A1(n_2132),
.A2(n_2128),
.B1(n_2129),
.B2(n_2130),
.Y(n_2143)
);

AO21x2_ASAP7_75t_L g2144 ( 
.A1(n_2131),
.A2(n_1756),
.B(n_442),
.Y(n_2144)
);

OR4x2_ASAP7_75t_L g2145 ( 
.A(n_2143),
.B(n_2125),
.C(n_1813),
.D(n_445),
.Y(n_2145)
);

XNOR2xp5_ASAP7_75t_L g2146 ( 
.A(n_2137),
.B(n_441),
.Y(n_2146)
);

OR5x1_ASAP7_75t_L g2147 ( 
.A(n_2134),
.B(n_2138),
.C(n_2135),
.D(n_2136),
.E(n_2139),
.Y(n_2147)
);

NOR3xp33_ASAP7_75t_L g2148 ( 
.A(n_2141),
.B(n_443),
.C(n_447),
.Y(n_2148)
);

OAI221xp5_ASAP7_75t_L g2149 ( 
.A1(n_2142),
.A2(n_1798),
.B1(n_1806),
.B2(n_1813),
.C(n_463),
.Y(n_2149)
);

AOI21xp33_ASAP7_75t_L g2150 ( 
.A1(n_2140),
.A2(n_456),
.B(n_457),
.Y(n_2150)
);

INVx2_ASAP7_75t_L g2151 ( 
.A(n_2144),
.Y(n_2151)
);

INVx2_ASAP7_75t_L g2152 ( 
.A(n_2136),
.Y(n_2152)
);

INVx2_ASAP7_75t_L g2153 ( 
.A(n_2136),
.Y(n_2153)
);

INVx1_ASAP7_75t_L g2154 ( 
.A(n_2135),
.Y(n_2154)
);

AOI222xp33_ASAP7_75t_L g2155 ( 
.A1(n_2154),
.A2(n_1841),
.B1(n_1714),
.B2(n_1853),
.C1(n_1842),
.C2(n_1806),
.Y(n_2155)
);

OR3x2_ASAP7_75t_L g2156 ( 
.A(n_2147),
.B(n_461),
.C(n_465),
.Y(n_2156)
);

AOI222xp33_ASAP7_75t_SL g2157 ( 
.A1(n_2152),
.A2(n_467),
.B1(n_468),
.B2(n_469),
.C1(n_472),
.C2(n_474),
.Y(n_2157)
);

INVx1_ASAP7_75t_L g2158 ( 
.A(n_2146),
.Y(n_2158)
);

OAI22xp5_ASAP7_75t_L g2159 ( 
.A1(n_2153),
.A2(n_1840),
.B1(n_1821),
.B2(n_1853),
.Y(n_2159)
);

AND3x4_ASAP7_75t_L g2160 ( 
.A(n_2151),
.B(n_1714),
.C(n_476),
.Y(n_2160)
);

NOR4xp25_ASAP7_75t_L g2161 ( 
.A(n_2150),
.B(n_475),
.C(n_477),
.D(n_478),
.Y(n_2161)
);

INVxp67_ASAP7_75t_SL g2162 ( 
.A(n_2148),
.Y(n_2162)
);

AOI21xp5_ASAP7_75t_L g2163 ( 
.A1(n_2162),
.A2(n_2158),
.B(n_2161),
.Y(n_2163)
);

OAI21xp5_ASAP7_75t_L g2164 ( 
.A1(n_2156),
.A2(n_2145),
.B(n_2149),
.Y(n_2164)
);

OAI21xp5_ASAP7_75t_L g2165 ( 
.A1(n_2160),
.A2(n_1669),
.B(n_1685),
.Y(n_2165)
);

OAI22xp5_ASAP7_75t_L g2166 ( 
.A1(n_2159),
.A2(n_1840),
.B1(n_1841),
.B2(n_1864),
.Y(n_2166)
);

NAND2xp5_ASAP7_75t_L g2167 ( 
.A(n_2157),
.B(n_480),
.Y(n_2167)
);

OAI21xp5_ASAP7_75t_L g2168 ( 
.A1(n_2163),
.A2(n_2155),
.B(n_1691),
.Y(n_2168)
);

NAND2xp5_ASAP7_75t_L g2169 ( 
.A(n_2167),
.B(n_481),
.Y(n_2169)
);

INVx1_ASAP7_75t_L g2170 ( 
.A(n_2169),
.Y(n_2170)
);

OR2x6_ASAP7_75t_L g2171 ( 
.A(n_2170),
.B(n_2164),
.Y(n_2171)
);

AOI221xp5_ASAP7_75t_L g2172 ( 
.A1(n_2171),
.A2(n_2168),
.B1(n_2166),
.B2(n_2165),
.C(n_485),
.Y(n_2172)
);

AOI211xp5_ASAP7_75t_L g2173 ( 
.A1(n_2172),
.A2(n_482),
.B(n_483),
.C(n_484),
.Y(n_2173)
);


endmodule