module fake_jpeg_5361_n_126 (n_11, n_3, n_2, n_1, n_0, n_10, n_4, n_8, n_9, n_6, n_5, n_7, n_126);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_126;

wire n_117;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_114;
wire n_74;
wire n_31;
wire n_29;
wire n_103;
wire n_50;
wire n_15;
wire n_124;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_109;
wire n_113;
wire n_30;
wire n_106;
wire n_111;
wire n_24;
wire n_44;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_20;
wire n_18;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_56;
wire n_79;
wire n_12;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_22;
wire n_101;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_97;
wire n_36;
wire n_62;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_96;

CKINVDCx20_ASAP7_75t_R g12 ( 
.A(n_9),
.Y(n_12)
);

BUFx16f_ASAP7_75t_L g13 ( 
.A(n_2),
.Y(n_13)
);

BUFx3_ASAP7_75t_L g14 ( 
.A(n_7),
.Y(n_14)
);

BUFx6f_ASAP7_75t_L g15 ( 
.A(n_5),
.Y(n_15)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_7),
.Y(n_16)
);

BUFx6f_ASAP7_75t_L g17 ( 
.A(n_5),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_4),
.Y(n_18)
);

INVx3_ASAP7_75t_L g19 ( 
.A(n_0),
.Y(n_19)
);

INVx11_ASAP7_75t_SL g20 ( 
.A(n_6),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_6),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_2),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_0),
.Y(n_23)
);

BUFx12_ASAP7_75t_L g24 ( 
.A(n_8),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_1),
.Y(n_25)
);

BUFx10_ASAP7_75t_L g26 ( 
.A(n_3),
.Y(n_26)
);

AND2x2_ASAP7_75t_L g27 ( 
.A(n_13),
.B(n_0),
.Y(n_27)
);

NOR2xp33_ASAP7_75t_SL g42 ( 
.A(n_27),
.B(n_31),
.Y(n_42)
);

BUFx12f_ASAP7_75t_L g28 ( 
.A(n_13),
.Y(n_28)
);

INVx6_ASAP7_75t_L g43 ( 
.A(n_28),
.Y(n_43)
);

INVx6_ASAP7_75t_L g29 ( 
.A(n_13),
.Y(n_29)
);

INVx8_ASAP7_75t_L g49 ( 
.A(n_29),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_20),
.Y(n_30)
);

NOR2xp33_ASAP7_75t_L g51 ( 
.A(n_30),
.B(n_34),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g31 ( 
.A(n_12),
.B(n_1),
.Y(n_31)
);

INVx6_ASAP7_75t_SL g32 ( 
.A(n_24),
.Y(n_32)
);

INVx1_ASAP7_75t_SL g52 ( 
.A(n_32),
.Y(n_52)
);

INVx8_ASAP7_75t_L g33 ( 
.A(n_14),
.Y(n_33)
);

AOI22xp33_ASAP7_75t_SL g57 ( 
.A1(n_33),
.A2(n_19),
.B1(n_25),
.B2(n_23),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_17),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_L g35 ( 
.A(n_12),
.B(n_1),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_SL g48 ( 
.A(n_35),
.B(n_18),
.Y(n_48)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_26),
.Y(n_36)
);

NAND2xp5_ASAP7_75t_L g44 ( 
.A(n_36),
.B(n_39),
.Y(n_44)
);

INVx5_ASAP7_75t_L g37 ( 
.A(n_26),
.Y(n_37)
);

INVx3_ASAP7_75t_L g55 ( 
.A(n_37),
.Y(n_55)
);

INVx2_ASAP7_75t_L g38 ( 
.A(n_14),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_38),
.B(n_17),
.Y(n_53)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_26),
.Y(n_39)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_32),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_40),
.B(n_45),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_SL g41 ( 
.A(n_27),
.B(n_18),
.Y(n_41)
);

NAND2xp5_ASAP7_75t_L g68 ( 
.A(n_41),
.B(n_60),
.Y(n_68)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_37),
.Y(n_45)
);

INVx2_ASAP7_75t_SL g46 ( 
.A(n_38),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_46),
.B(n_47),
.Y(n_70)
);

INVx2_ASAP7_75t_L g47 ( 
.A(n_30),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_48),
.B(n_56),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_L g50 ( 
.A(n_27),
.B(n_25),
.Y(n_50)
);

AND2x2_ASAP7_75t_L g71 ( 
.A(n_50),
.B(n_24),
.Y(n_71)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_53),
.Y(n_72)
);

OAI22xp5_ASAP7_75t_L g54 ( 
.A1(n_33),
.A2(n_19),
.B1(n_21),
.B2(n_23),
.Y(n_54)
);

AOI22xp5_ASAP7_75t_L g76 ( 
.A1(n_54),
.A2(n_15),
.B1(n_22),
.B2(n_24),
.Y(n_76)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_34),
.Y(n_56)
);

INVxp67_ASAP7_75t_L g63 ( 
.A(n_57),
.Y(n_63)
);

INVx3_ASAP7_75t_L g58 ( 
.A(n_36),
.Y(n_58)
);

INVx1_ASAP7_75t_SL g73 ( 
.A(n_58),
.Y(n_73)
);

INVx2_ASAP7_75t_L g59 ( 
.A(n_39),
.Y(n_59)
);

INVx3_ASAP7_75t_L g78 ( 
.A(n_59),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_SL g60 ( 
.A(n_29),
.B(n_16),
.Y(n_60)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_47),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_61),
.B(n_66),
.Y(n_83)
);

OAI22xp33_ASAP7_75t_SL g62 ( 
.A1(n_50),
.A2(n_21),
.B1(n_16),
.B2(n_17),
.Y(n_62)
);

AOI22xp5_ASAP7_75t_SL g90 ( 
.A1(n_62),
.A2(n_43),
.B1(n_15),
.B2(n_22),
.Y(n_90)
);

XOR2xp5_ASAP7_75t_L g64 ( 
.A(n_44),
.B(n_28),
.Y(n_64)
);

XNOR2xp5_ASAP7_75t_L g87 ( 
.A(n_64),
.B(n_67),
.Y(n_87)
);

BUFx5_ASAP7_75t_L g66 ( 
.A(n_43),
.Y(n_66)
);

MAJIxp5_ASAP7_75t_L g67 ( 
.A(n_44),
.B(n_28),
.C(n_26),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_L g69 ( 
.A(n_42),
.B(n_2),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_69),
.B(n_75),
.Y(n_89)
);

XNOR2xp5_ASAP7_75t_SL g91 ( 
.A(n_71),
.B(n_24),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_L g75 ( 
.A(n_59),
.B(n_3),
.Y(n_75)
);

OAI22xp5_ASAP7_75t_SL g82 ( 
.A1(n_76),
.A2(n_55),
.B1(n_49),
.B2(n_56),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_L g77 ( 
.A(n_46),
.B(n_4),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_L g92 ( 
.A(n_77),
.B(n_8),
.Y(n_92)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_70),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_79),
.B(n_80),
.Y(n_98)
);

INVx2_ASAP7_75t_L g80 ( 
.A(n_66),
.Y(n_80)
);

CKINVDCx20_ASAP7_75t_R g81 ( 
.A(n_65),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_81),
.B(n_88),
.Y(n_102)
);

AOI22xp5_ASAP7_75t_L g100 ( 
.A1(n_82),
.A2(n_90),
.B1(n_63),
.B2(n_73),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_SL g84 ( 
.A(n_74),
.B(n_58),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_SL g93 ( 
.A(n_84),
.B(n_72),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_SL g85 ( 
.A(n_68),
.B(n_51),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_L g95 ( 
.A(n_85),
.B(n_92),
.Y(n_95)
);

OA22x2_ASAP7_75t_SL g86 ( 
.A1(n_64),
.A2(n_46),
.B1(n_55),
.B2(n_49),
.Y(n_86)
);

AO21x1_ASAP7_75t_L g96 ( 
.A1(n_86),
.A2(n_91),
.B(n_71),
.Y(n_96)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_73),
.Y(n_88)
);

MAJIxp5_ASAP7_75t_L g97 ( 
.A(n_91),
.B(n_67),
.C(n_71),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g105 ( 
.A(n_93),
.B(n_99),
.Y(n_105)
);

BUFx12_ASAP7_75t_L g94 ( 
.A(n_86),
.Y(n_94)
);

CKINVDCx20_ASAP7_75t_R g104 ( 
.A(n_94),
.Y(n_104)
);

A2O1A1O1Ixp25_ASAP7_75t_L g106 ( 
.A1(n_96),
.A2(n_94),
.B(n_101),
.C(n_97),
.D(n_90),
.Y(n_106)
);

MAJIxp5_ASAP7_75t_L g107 ( 
.A(n_97),
.B(n_101),
.C(n_82),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_SL g99 ( 
.A(n_89),
.B(n_63),
.Y(n_99)
);

XNOR2xp5_ASAP7_75t_L g109 ( 
.A(n_100),
.B(n_52),
.Y(n_109)
);

XOR2xp5_ASAP7_75t_L g101 ( 
.A(n_87),
.B(n_76),
.Y(n_101)
);

MAJx2_ASAP7_75t_L g103 ( 
.A(n_96),
.B(n_87),
.C(n_86),
.Y(n_103)
);

MAJIxp5_ASAP7_75t_L g112 ( 
.A(n_103),
.B(n_107),
.C(n_108),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_SL g110 ( 
.A(n_106),
.B(n_94),
.Y(n_110)
);

MAJIxp5_ASAP7_75t_L g108 ( 
.A(n_95),
.B(n_83),
.C(n_52),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_L g113 ( 
.A(n_109),
.B(n_98),
.Y(n_113)
);

AND2x2_ASAP7_75t_L g117 ( 
.A(n_110),
.B(n_113),
.Y(n_117)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_105),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_L g118 ( 
.A(n_111),
.B(n_114),
.Y(n_118)
);

AOI21xp5_ASAP7_75t_L g114 ( 
.A1(n_104),
.A2(n_103),
.B(n_106),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_SL g115 ( 
.A(n_112),
.B(n_102),
.Y(n_115)
);

CKINVDCx16_ASAP7_75t_R g121 ( 
.A(n_115),
.Y(n_121)
);

CKINVDCx20_ASAP7_75t_R g116 ( 
.A(n_112),
.Y(n_116)
);

NOR2xp67_ASAP7_75t_SL g119 ( 
.A(n_116),
.B(n_80),
.Y(n_119)
);

HB1xp67_ASAP7_75t_L g122 ( 
.A(n_119),
.Y(n_122)
);

AOI322xp5_ASAP7_75t_L g120 ( 
.A1(n_117),
.A2(n_9),
.A3(n_10),
.B1(n_11),
.B2(n_78),
.C1(n_115),
.C2(n_118),
.Y(n_120)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_120),
.Y(n_123)
);

AOI21xp5_ASAP7_75t_L g124 ( 
.A1(n_122),
.A2(n_121),
.B(n_11),
.Y(n_124)
);

MAJIxp5_ASAP7_75t_L g125 ( 
.A(n_124),
.B(n_123),
.C(n_10),
.Y(n_125)
);

XOR2xp5_ASAP7_75t_L g126 ( 
.A(n_125),
.B(n_78),
.Y(n_126)
);


endmodule