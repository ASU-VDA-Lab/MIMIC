module fake_netlist_6_136_n_1980 (n_52, n_16, n_1, n_91, n_119, n_46, n_146, n_163, n_18, n_21, n_193, n_147, n_154, n_191, n_88, n_3, n_209, n_98, n_113, n_39, n_63, n_73, n_4, n_148, n_199, n_138, n_22, n_161, n_208, n_68, n_166, n_28, n_184, n_50, n_158, n_49, n_7, n_83, n_206, n_5, n_101, n_167, n_144, n_174, n_127, n_125, n_153, n_168, n_178, n_77, n_156, n_149, n_152, n_106, n_92, n_145, n_42, n_133, n_96, n_8, n_90, n_160, n_24, n_105, n_131, n_54, n_132, n_188, n_102, n_186, n_204, n_0, n_87, n_195, n_189, n_32, n_66, n_85, n_99, n_78, n_84, n_130, n_164, n_100, n_129, n_13, n_121, n_197, n_11, n_137, n_17, n_23, n_203, n_142, n_20, n_143, n_207, n_2, n_180, n_19, n_47, n_62, n_29, n_155, n_75, n_109, n_150, n_122, n_45, n_205, n_34, n_140, n_70, n_120, n_37, n_15, n_67, n_33, n_82, n_27, n_38, n_110, n_151, n_61, n_112, n_172, n_81, n_59, n_181, n_76, n_36, n_182, n_26, n_124, n_55, n_126, n_202, n_94, n_97, n_108, n_58, n_116, n_64, n_117, n_118, n_175, n_48, n_65, n_25, n_40, n_93, n_80, n_141, n_135, n_196, n_200, n_165, n_139, n_41, n_134, n_177, n_176, n_114, n_86, n_198, n_104, n_95, n_179, n_9, n_107, n_10, n_71, n_74, n_6, n_190, n_14, n_123, n_136, n_72, n_187, n_89, n_173, n_201, n_103, n_111, n_60, n_159, n_157, n_162, n_170, n_185, n_35, n_183, n_115, n_12, n_69, n_128, n_30, n_79, n_43, n_194, n_171, n_31, n_192, n_57, n_169, n_53, n_51, n_44, n_56, n_1980);

input n_52;
input n_16;
input n_1;
input n_91;
input n_119;
input n_46;
input n_146;
input n_163;
input n_18;
input n_21;
input n_193;
input n_147;
input n_154;
input n_191;
input n_88;
input n_3;
input n_209;
input n_98;
input n_113;
input n_39;
input n_63;
input n_73;
input n_4;
input n_148;
input n_199;
input n_138;
input n_22;
input n_161;
input n_208;
input n_68;
input n_166;
input n_28;
input n_184;
input n_50;
input n_158;
input n_49;
input n_7;
input n_83;
input n_206;
input n_5;
input n_101;
input n_167;
input n_144;
input n_174;
input n_127;
input n_125;
input n_153;
input n_168;
input n_178;
input n_77;
input n_156;
input n_149;
input n_152;
input n_106;
input n_92;
input n_145;
input n_42;
input n_133;
input n_96;
input n_8;
input n_90;
input n_160;
input n_24;
input n_105;
input n_131;
input n_54;
input n_132;
input n_188;
input n_102;
input n_186;
input n_204;
input n_0;
input n_87;
input n_195;
input n_189;
input n_32;
input n_66;
input n_85;
input n_99;
input n_78;
input n_84;
input n_130;
input n_164;
input n_100;
input n_129;
input n_13;
input n_121;
input n_197;
input n_11;
input n_137;
input n_17;
input n_23;
input n_203;
input n_142;
input n_20;
input n_143;
input n_207;
input n_2;
input n_180;
input n_19;
input n_47;
input n_62;
input n_29;
input n_155;
input n_75;
input n_109;
input n_150;
input n_122;
input n_45;
input n_205;
input n_34;
input n_140;
input n_70;
input n_120;
input n_37;
input n_15;
input n_67;
input n_33;
input n_82;
input n_27;
input n_38;
input n_110;
input n_151;
input n_61;
input n_112;
input n_172;
input n_81;
input n_59;
input n_181;
input n_76;
input n_36;
input n_182;
input n_26;
input n_124;
input n_55;
input n_126;
input n_202;
input n_94;
input n_97;
input n_108;
input n_58;
input n_116;
input n_64;
input n_117;
input n_118;
input n_175;
input n_48;
input n_65;
input n_25;
input n_40;
input n_93;
input n_80;
input n_141;
input n_135;
input n_196;
input n_200;
input n_165;
input n_139;
input n_41;
input n_134;
input n_177;
input n_176;
input n_114;
input n_86;
input n_198;
input n_104;
input n_95;
input n_179;
input n_9;
input n_107;
input n_10;
input n_71;
input n_74;
input n_6;
input n_190;
input n_14;
input n_123;
input n_136;
input n_72;
input n_187;
input n_89;
input n_173;
input n_201;
input n_103;
input n_111;
input n_60;
input n_159;
input n_157;
input n_162;
input n_170;
input n_185;
input n_35;
input n_183;
input n_115;
input n_12;
input n_69;
input n_128;
input n_30;
input n_79;
input n_43;
input n_194;
input n_171;
input n_31;
input n_192;
input n_57;
input n_169;
input n_53;
input n_51;
input n_44;
input n_56;

output n_1980;

wire n_992;
wire n_1671;
wire n_801;
wire n_1613;
wire n_1234;
wire n_1458;
wire n_1199;
wire n_1674;
wire n_741;
wire n_1027;
wire n_1351;
wire n_625;
wire n_1189;
wire n_223;
wire n_1212;
wire n_226;
wire n_726;
wire n_212;
wire n_700;
wire n_1307;
wire n_1038;
wire n_578;
wire n_1581;
wire n_1003;
wire n_365;
wire n_1237;
wire n_1061;
wire n_1357;
wire n_1853;
wire n_783;
wire n_1738;
wire n_798;
wire n_1575;
wire n_1854;
wire n_1923;
wire n_509;
wire n_1342;
wire n_245;
wire n_1209;
wire n_1348;
wire n_1387;
wire n_677;
wire n_1708;
wire n_805;
wire n_1151;
wire n_396;
wire n_1739;
wire n_350;
wire n_1380;
wire n_442;
wire n_480;
wire n_1402;
wire n_1688;
wire n_1691;
wire n_1975;
wire n_1009;
wire n_1743;
wire n_1930;
wire n_1160;
wire n_883;
wire n_1238;
wire n_1724;
wire n_1032;
wire n_1247;
wire n_1547;
wire n_1553;
wire n_893;
wire n_1099;
wire n_1264;
wire n_1192;
wire n_471;
wire n_1844;
wire n_424;
wire n_1700;
wire n_1555;
wire n_1415;
wire n_1370;
wire n_1786;
wire n_369;
wire n_287;
wire n_415;
wire n_830;
wire n_230;
wire n_461;
wire n_873;
wire n_383;
wire n_1285;
wire n_1371;
wire n_447;
wire n_1803;
wire n_1172;
wire n_852;
wire n_229;
wire n_1590;
wire n_1532;
wire n_1393;
wire n_1517;
wire n_1867;
wire n_1704;
wire n_1078;
wire n_250;
wire n_544;
wire n_1711;
wire n_1140;
wire n_1444;
wire n_1670;
wire n_1603;
wire n_1579;
wire n_1263;
wire n_836;
wire n_375;
wire n_522;
wire n_1261;
wire n_945;
wire n_1649;
wire n_1903;
wire n_1511;
wire n_1143;
wire n_1422;
wire n_1232;
wire n_1772;
wire n_1572;
wire n_616;
wire n_658;
wire n_1874;
wire n_1119;
wire n_428;
wire n_1433;
wire n_1902;
wire n_1842;
wire n_1620;
wire n_1954;
wire n_1735;
wire n_1541;
wire n_1300;
wire n_641;
wire n_822;
wire n_693;
wire n_1313;
wire n_1056;
wire n_758;
wire n_516;
wire n_1455;
wire n_1163;
wire n_1180;
wire n_943;
wire n_1798;
wire n_1550;
wire n_491;
wire n_1591;
wire n_772;
wire n_1344;
wire n_666;
wire n_371;
wire n_940;
wire n_770;
wire n_567;
wire n_1781;
wire n_1971;
wire n_405;
wire n_213;
wire n_538;
wire n_1106;
wire n_886;
wire n_1471;
wire n_343;
wire n_1094;
wire n_953;
wire n_1345;
wire n_1820;
wire n_494;
wire n_539;
wire n_493;
wire n_454;
wire n_1421;
wire n_1936;
wire n_638;
wire n_1404;
wire n_1211;
wire n_381;
wire n_887;
wire n_1660;
wire n_1961;
wire n_1280;
wire n_713;
wire n_1400;
wire n_1467;
wire n_976;
wire n_224;
wire n_1445;
wire n_1526;
wire n_1560;
wire n_734;
wire n_1088;
wire n_1894;
wire n_1231;
wire n_1978;
wire n_917;
wire n_574;
wire n_907;
wire n_1446;
wire n_659;
wire n_1815;
wire n_407;
wire n_913;
wire n_1658;
wire n_808;
wire n_867;
wire n_1230;
wire n_473;
wire n_1193;
wire n_1967;
wire n_1054;
wire n_559;
wire n_1333;
wire n_1648;
wire n_1911;
wire n_1956;
wire n_1644;
wire n_1558;
wire n_1732;
wire n_281;
wire n_551;
wire n_699;
wire n_564;
wire n_451;
wire n_824;
wire n_279;
wire n_686;
wire n_757;
wire n_594;
wire n_1641;
wire n_1918;
wire n_577;
wire n_1843;
wire n_619;
wire n_1367;
wire n_1336;
wire n_521;
wire n_572;
wire n_395;
wire n_813;
wire n_1909;
wire n_1481;
wire n_323;
wire n_606;
wire n_1441;
wire n_818;
wire n_1123;
wire n_1309;
wire n_513;
wire n_645;
wire n_1381;
wire n_331;
wire n_1699;
wire n_916;
wire n_483;
wire n_1970;
wire n_608;
wire n_261;
wire n_630;
wire n_541;
wire n_512;
wire n_433;
wire n_792;
wire n_476;
wire n_1328;
wire n_1957;
wire n_219;
wire n_1907;
wire n_264;
wire n_263;
wire n_1162;
wire n_860;
wire n_1530;
wire n_788;
wire n_939;
wire n_1543;
wire n_821;
wire n_938;
wire n_1302;
wire n_1068;
wire n_1599;
wire n_329;
wire n_982;
wire n_549;
wire n_1762;
wire n_1910;
wire n_1075;
wire n_408;
wire n_932;
wire n_237;
wire n_1876;
wire n_1895;
wire n_1697;
wire n_243;
wire n_979;
wire n_1873;
wire n_905;
wire n_1866;
wire n_1680;
wire n_322;
wire n_993;
wire n_689;
wire n_354;
wire n_1413;
wire n_1330;
wire n_1605;
wire n_1278;
wire n_547;
wire n_558;
wire n_1064;
wire n_1396;
wire n_634;
wire n_966;
wire n_764;
wire n_1663;
wire n_692;
wire n_733;
wire n_1793;
wire n_1233;
wire n_1289;
wire n_487;
wire n_241;
wire n_1107;
wire n_1014;
wire n_1290;
wire n_1703;
wire n_882;
wire n_1354;
wire n_586;
wire n_423;
wire n_1865;
wire n_1875;
wire n_1701;
wire n_318;
wire n_1111;
wire n_1713;
wire n_715;
wire n_1251;
wire n_1265;
wire n_1726;
wire n_1950;
wire n_530;
wire n_1563;
wire n_1912;
wire n_277;
wire n_618;
wire n_1297;
wire n_1662;
wire n_1312;
wire n_1167;
wire n_1359;
wire n_674;
wire n_871;
wire n_922;
wire n_268;
wire n_1335;
wire n_1760;
wire n_1927;
wire n_210;
wire n_1069;
wire n_1722;
wire n_1664;
wire n_612;
wire n_247;
wire n_1165;
wire n_355;
wire n_702;
wire n_347;
wire n_1926;
wire n_1175;
wire n_328;
wire n_1386;
wire n_1896;
wire n_429;
wire n_1747;
wire n_1012;
wire n_780;
wire n_675;
wire n_903;
wire n_1540;
wire n_1977;
wire n_1802;
wire n_1504;
wire n_286;
wire n_254;
wire n_1655;
wire n_242;
wire n_835;
wire n_1214;
wire n_928;
wire n_690;
wire n_850;
wire n_1886;
wire n_1801;
wire n_1654;
wire n_816;
wire n_1157;
wire n_1750;
wire n_1462;
wire n_1188;
wire n_1752;
wire n_877;
wire n_1813;
wire n_604;
wire n_825;
wire n_728;
wire n_1063;
wire n_1588;
wire n_267;
wire n_1124;
wire n_1624;
wire n_515;
wire n_1965;
wire n_598;
wire n_696;
wire n_1515;
wire n_961;
wire n_437;
wire n_1082;
wire n_1317;
wire n_593;
wire n_514;
wire n_687;
wire n_697;
wire n_890;
wire n_637;
wire n_295;
wire n_701;
wire n_950;
wire n_388;
wire n_484;
wire n_1709;
wire n_1825;
wire n_1757;
wire n_1796;
wire n_1792;
wire n_891;
wire n_1412;
wire n_949;
wire n_1630;
wire n_678;
wire n_283;
wire n_507;
wire n_968;
wire n_909;
wire n_1369;
wire n_881;
wire n_1008;
wire n_760;
wire n_1546;
wire n_590;
wire n_362;
wire n_462;
wire n_1052;
wire n_1033;
wire n_1296;
wire n_304;
wire n_694;
wire n_1294;
wire n_1420;
wire n_1634;
wire n_595;
wire n_627;
wire n_297;
wire n_1767;
wire n_1779;
wire n_524;
wire n_1465;
wire n_342;
wire n_1858;
wire n_1044;
wire n_1712;
wire n_1391;
wire n_449;
wire n_1523;
wire n_1208;
wire n_1164;
wire n_1295;
wire n_1627;
wire n_1072;
wire n_1527;
wire n_1495;
wire n_1438;
wire n_495;
wire n_815;
wire n_1100;
wire n_585;
wire n_1487;
wire n_840;
wire n_874;
wire n_1756;
wire n_1128;
wire n_382;
wire n_673;
wire n_1969;
wire n_1071;
wire n_1067;
wire n_1565;
wire n_1493;
wire n_1968;
wire n_898;
wire n_255;
wire n_284;
wire n_1952;
wire n_865;
wire n_925;
wire n_1932;
wire n_1101;
wire n_1026;
wire n_1880;
wire n_289;
wire n_1364;
wire n_615;
wire n_1249;
wire n_1293;
wire n_1127;
wire n_1512;
wire n_1451;
wire n_320;
wire n_639;
wire n_963;
wire n_794;
wire n_727;
wire n_894;
wire n_1839;
wire n_685;
wire n_1765;
wire n_353;
wire n_605;
wire n_1514;
wire n_1863;
wire n_826;
wire n_1646;
wire n_872;
wire n_1139;
wire n_1714;
wire n_718;
wire n_1018;
wire n_1521;
wire n_1366;
wire n_542;
wire n_847;
wire n_644;
wire n_682;
wire n_851;
wire n_305;
wire n_996;
wire n_532;
wire n_1308;
wire n_1376;
wire n_1513;
wire n_413;
wire n_791;
wire n_1913;
wire n_510;
wire n_837;
wire n_1488;
wire n_1808;
wire n_948;
wire n_704;
wire n_977;
wire n_1005;
wire n_1947;
wire n_536;
wire n_1788;
wire n_622;
wire n_1469;
wire n_1838;
wire n_1835;
wire n_1776;
wire n_1766;
wire n_1959;
wire n_581;
wire n_765;
wire n_432;
wire n_987;
wire n_1492;
wire n_1340;
wire n_1771;
wire n_631;
wire n_720;
wire n_842;
wire n_1707;
wire n_1432;
wire n_843;
wire n_656;
wire n_989;
wire n_1277;
wire n_797;
wire n_1473;
wire n_1723;
wire n_1246;
wire n_1878;
wire n_899;
wire n_738;
wire n_1304;
wire n_1035;
wire n_294;
wire n_499;
wire n_1426;
wire n_705;
wire n_1004;
wire n_1176;
wire n_1529;
wire n_1022;
wire n_614;
wire n_529;
wire n_425;
wire n_684;
wire n_1431;
wire n_1615;
wire n_1474;
wire n_1571;
wire n_1809;
wire n_1577;
wire n_1181;
wire n_1822;
wire n_486;
wire n_947;
wire n_1117;
wire n_1087;
wire n_1448;
wire n_648;
wire n_657;
wire n_1049;
wire n_1666;
wire n_1505;
wire n_803;
wire n_290;
wire n_1717;
wire n_926;
wire n_1817;
wire n_927;
wire n_1849;
wire n_919;
wire n_1698;
wire n_478;
wire n_929;
wire n_1228;
wire n_417;
wire n_446;
wire n_1568;
wire n_1490;
wire n_777;
wire n_1299;
wire n_272;
wire n_526;
wire n_1183;
wire n_1436;
wire n_1384;
wire n_293;
wire n_458;
wire n_1070;
wire n_998;
wire n_717;
wire n_1665;
wire n_1383;
wire n_1178;
wire n_1424;
wire n_1073;
wire n_1000;
wire n_796;
wire n_252;
wire n_1195;
wire n_1626;
wire n_1507;
wire n_552;
wire n_1358;
wire n_1811;
wire n_1388;
wire n_216;
wire n_912;
wire n_1857;
wire n_1519;
wire n_745;
wire n_1284;
wire n_1604;
wire n_1142;
wire n_716;
wire n_1475;
wire n_623;
wire n_1048;
wire n_1201;
wire n_1398;
wire n_884;
wire n_1774;
wire n_1395;
wire n_731;
wire n_1502;
wire n_1659;
wire n_1955;
wire n_755;
wire n_1021;
wire n_931;
wire n_527;
wire n_474;
wire n_683;
wire n_811;
wire n_1207;
wire n_312;
wire n_1791;
wire n_1368;
wire n_1418;
wire n_958;
wire n_292;
wire n_1250;
wire n_1137;
wire n_1897;
wire n_880;
wire n_889;
wire n_1478;
wire n_589;
wire n_1310;
wire n_819;
wire n_1363;
wire n_1334;
wire n_1942;
wire n_1966;
wire n_767;
wire n_1314;
wire n_600;
wire n_964;
wire n_831;
wire n_1837;
wire n_477;
wire n_954;
wire n_864;
wire n_1110;
wire n_1410;
wire n_399;
wire n_1440;
wire n_1382;
wire n_1534;
wire n_1564;
wire n_1736;
wire n_211;
wire n_1483;
wire n_1834;
wire n_1372;
wire n_231;
wire n_1457;
wire n_505;
wire n_1719;
wire n_319;
wire n_1339;
wire n_1787;
wire n_537;
wire n_1427;
wire n_311;
wire n_1466;
wire n_403;
wire n_1919;
wire n_1080;
wire n_723;
wire n_1877;
wire n_596;
wire n_546;
wire n_562;
wire n_1141;
wire n_1268;
wire n_386;
wire n_1939;
wire n_1769;
wire n_1220;
wire n_1893;
wire n_556;
wire n_1755;
wire n_1602;
wire n_1136;
wire n_1125;
wire n_970;
wire n_642;
wire n_1159;
wire n_276;
wire n_995;
wire n_1092;
wire n_441;
wire n_221;
wire n_1060;
wire n_1951;
wire n_444;
wire n_1252;
wire n_1784;
wire n_1223;
wire n_303;
wire n_511;
wire n_1286;
wire n_1775;
wire n_1773;
wire n_1053;
wire n_416;
wire n_1681;
wire n_520;
wire n_418;
wire n_1093;
wire n_1783;
wire n_1533;
wire n_1597;
wire n_266;
wire n_296;
wire n_775;
wire n_651;
wire n_1153;
wire n_439;
wire n_1618;
wire n_217;
wire n_518;
wire n_1531;
wire n_1185;
wire n_453;
wire n_215;
wire n_1745;
wire n_914;
wire n_759;
wire n_1831;
wire n_426;
wire n_317;
wire n_1653;
wire n_1679;
wire n_1625;
wire n_1453;
wire n_488;
wire n_497;
wire n_773;
wire n_1901;
wire n_920;
wire n_1374;
wire n_1315;
wire n_1647;
wire n_1224;
wire n_1614;
wire n_1459;
wire n_1892;
wire n_1933;
wire n_1135;
wire n_1179;
wire n_1169;
wire n_401;
wire n_324;
wire n_1617;
wire n_335;
wire n_1470;
wire n_463;
wire n_1243;
wire n_848;
wire n_301;
wire n_274;
wire n_1096;
wire n_1091;
wire n_1917;
wire n_1580;
wire n_1425;
wire n_1881;
wire n_1267;
wire n_1281;
wire n_1806;
wire n_983;
wire n_427;
wire n_1520;
wire n_496;
wire n_906;
wire n_1390;
wire n_688;
wire n_1077;
wire n_1733;
wire n_1419;
wire n_351;
wire n_259;
wire n_1731;
wire n_1855;
wire n_1636;
wire n_1437;
wire n_1645;
wire n_1832;
wire n_385;
wire n_1687;
wire n_1439;
wire n_1323;
wire n_858;
wire n_1331;
wire n_613;
wire n_736;
wire n_501;
wire n_956;
wire n_960;
wire n_663;
wire n_856;
wire n_379;
wire n_778;
wire n_1668;
wire n_1134;
wire n_410;
wire n_1129;
wire n_554;
wire n_602;
wire n_1696;
wire n_1594;
wire n_664;
wire n_1869;
wire n_1764;
wire n_1429;
wire n_1610;
wire n_1889;
wire n_435;
wire n_1905;
wire n_793;
wire n_326;
wire n_587;
wire n_1593;
wire n_580;
wire n_762;
wire n_1030;
wire n_1202;
wire n_1937;
wire n_465;
wire n_1790;
wire n_1778;
wire n_1635;
wire n_1079;
wire n_341;
wire n_1744;
wire n_828;
wire n_607;
wire n_316;
wire n_419;
wire n_1551;
wire n_1103;
wire n_1203;
wire n_820;
wire n_951;
wire n_725;
wire n_952;
wire n_999;
wire n_358;
wire n_1254;
wire n_575;
wire n_368;
wire n_994;
wire n_1508;
wire n_732;
wire n_974;
wire n_392;
wire n_724;
wire n_1934;
wire n_1020;
wire n_1042;
wire n_628;
wire n_1273;
wire n_1434;
wire n_1573;
wire n_1728;
wire n_557;
wire n_1871;
wire n_349;
wire n_617;
wire n_845;
wire n_807;
wire n_1036;
wire n_1138;
wire n_1661;
wire n_1275;
wire n_485;
wire n_1549;
wire n_443;
wire n_1510;
wire n_892;
wire n_768;
wire n_421;
wire n_1468;
wire n_1859;
wire n_238;
wire n_1095;
wire n_1595;
wire n_1718;
wire n_1749;
wire n_1683;
wire n_1916;
wire n_597;
wire n_280;
wire n_1270;
wire n_1187;
wire n_610;
wire n_1403;
wire n_1669;
wire n_1852;
wire n_1024;
wire n_1768;
wire n_1847;
wire n_248;
wire n_517;
wire n_1667;
wire n_667;
wire n_1206;
wire n_621;
wire n_1037;
wire n_1397;
wire n_1279;
wire n_1115;
wire n_750;
wire n_901;
wire n_1499;
wire n_468;
wire n_923;
wire n_504;
wire n_1409;
wire n_1841;
wire n_1639;
wire n_1623;
wire n_1015;
wire n_1503;
wire n_466;
wire n_1057;
wire n_603;
wire n_991;
wire n_1657;
wire n_235;
wire n_1126;
wire n_340;
wire n_710;
wire n_1108;
wire n_1818;
wire n_1182;
wire n_1298;
wire n_1611;
wire n_785;
wire n_746;
wire n_609;
wire n_1601;
wire n_1960;
wire n_1686;
wire n_1356;
wire n_1589;
wire n_1740;
wire n_1497;
wire n_1168;
wire n_1216;
wire n_1943;
wire n_1320;
wire n_1430;
wire n_1316;
wire n_1287;
wire n_1452;
wire n_1622;
wire n_1586;
wire n_302;
wire n_1694;
wire n_380;
wire n_1535;
wire n_1596;
wire n_1190;
wire n_1734;
wire n_397;
wire n_1938;
wire n_1262;
wire n_218;
wire n_1891;
wire n_1213;
wire n_1350;
wire n_1673;
wire n_1715;
wire n_1443;
wire n_1272;
wire n_239;
wire n_782;
wire n_1539;
wire n_490;
wire n_220;
wire n_809;
wire n_1043;
wire n_1797;
wire n_1608;
wire n_986;
wire n_1472;
wire n_1081;
wire n_402;
wire n_1870;
wire n_352;
wire n_1692;
wire n_800;
wire n_1084;
wire n_1171;
wire n_460;
wire n_1827;
wire n_1361;
wire n_1864;
wire n_1491;
wire n_662;
wire n_374;
wire n_1152;
wire n_1840;
wire n_1705;
wire n_450;
wire n_1684;
wire n_921;
wire n_1346;
wire n_711;
wire n_1642;
wire n_579;
wire n_1352;
wire n_937;
wire n_1682;
wire n_370;
wire n_1695;
wire n_1828;
wire n_650;
wire n_1046;
wire n_1940;
wire n_1979;
wire n_1145;
wire n_330;
wire n_1121;
wire n_1102;
wire n_1963;
wire n_972;
wire n_1405;
wire n_258;
wire n_1406;
wire n_456;
wire n_1332;
wire n_260;
wire n_313;
wire n_624;
wire n_962;
wire n_1041;
wire n_565;
wire n_356;
wire n_1569;
wire n_936;
wire n_1883;
wire n_1288;
wire n_1186;
wire n_1062;
wire n_885;
wire n_896;
wire n_654;
wire n_411;
wire n_1222;
wire n_599;
wire n_776;
wire n_321;
wire n_1823;
wire n_227;
wire n_1974;
wire n_1720;
wire n_482;
wire n_934;
wire n_1637;
wire n_1407;
wire n_1795;
wire n_420;
wire n_1341;
wire n_394;
wire n_1456;
wire n_1845;
wire n_1489;
wire n_942;
wire n_1524;
wire n_543;
wire n_1964;
wire n_1920;
wire n_1496;
wire n_1271;
wire n_1545;
wire n_1946;
wire n_1355;
wire n_1225;
wire n_1544;
wire n_1485;
wire n_325;
wire n_1640;
wire n_804;
wire n_464;
wire n_1846;
wire n_533;
wire n_806;
wire n_879;
wire n_959;
wire n_584;
wire n_244;
wire n_1343;
wire n_1522;
wire n_548;
wire n_1782;
wire n_282;
wire n_1676;
wire n_833;
wire n_1830;
wire n_1567;
wire n_523;
wire n_1319;
wire n_707;
wire n_345;
wire n_1900;
wire n_799;
wire n_1548;
wire n_1155;
wire n_273;
wire n_1633;
wire n_787;
wire n_1416;
wire n_1528;
wire n_1146;
wire n_1086;
wire n_1066;
wire n_1948;
wire n_1282;
wire n_550;
wire n_275;
wire n_652;
wire n_560;
wire n_1906;
wire n_1484;
wire n_1241;
wire n_1321;
wire n_1672;
wire n_569;
wire n_1758;
wire n_1925;
wire n_737;
wire n_1318;
wire n_1914;
wire n_1235;
wire n_1229;
wire n_306;
wire n_1292;
wire n_1373;
wire n_346;
wire n_1029;
wire n_1447;
wire n_790;
wire n_1706;
wire n_1498;
wire n_1210;
wire n_299;
wire n_1248;
wire n_1556;
wire n_902;
wire n_333;
wire n_1047;
wire n_1385;
wire n_431;
wire n_459;
wire n_1269;
wire n_1931;
wire n_502;
wire n_672;
wire n_1257;
wire n_1751;
wire n_285;
wire n_1375;
wire n_1941;
wire n_655;
wire n_706;
wire n_1045;
wire n_1650;
wire n_786;
wire n_1794;
wire n_1236;
wire n_1962;
wire n_1559;
wire n_1725;
wire n_1928;
wire n_1872;
wire n_834;
wire n_743;
wire n_766;
wire n_430;
wire n_1746;
wire n_1325;
wire n_1002;
wire n_1741;
wire n_1949;
wire n_545;
wire n_489;
wire n_1804;
wire n_1727;
wire n_251;
wire n_1019;
wire n_636;
wire n_729;
wire n_876;
wire n_774;
wire n_1337;
wire n_660;
wire n_438;
wire n_1477;
wire n_1360;
wire n_1860;
wire n_1904;
wire n_1200;
wire n_479;
wire n_1607;
wire n_1353;
wire n_1777;
wire n_1908;
wire n_1454;
wire n_869;
wire n_1154;
wire n_1113;
wire n_1600;
wire n_646;
wire n_528;
wire n_391;
wire n_1098;
wire n_1329;
wire n_817;
wire n_262;
wire n_897;
wire n_846;
wire n_841;
wire n_1476;
wire n_1001;
wire n_508;
wire n_1800;
wire n_1050;
wire n_1411;
wire n_1463;
wire n_1177;
wire n_332;
wire n_1150;
wire n_1742;
wire n_1562;
wire n_1690;
wire n_398;
wire n_1191;
wire n_1826;
wire n_566;
wire n_1023;
wire n_1882;
wire n_1076;
wire n_1118;
wire n_1007;
wire n_1929;
wire n_1807;
wire n_1378;
wire n_855;
wire n_1592;
wire n_1759;
wire n_1814;
wire n_1631;
wire n_591;
wire n_1377;
wire n_1879;
wire n_256;
wire n_853;
wire n_440;
wire n_695;
wire n_1542;
wire n_875;
wire n_367;
wire n_680;
wire n_1678;
wire n_661;
wire n_1716;
wire n_278;
wire n_1256;
wire n_671;
wire n_1953;
wire n_933;
wire n_740;
wire n_703;
wire n_978;
wire n_384;
wire n_1976;
wire n_1291;
wire n_1217;
wire n_751;
wire n_749;
wire n_1824;
wire n_310;
wire n_1628;
wire n_1324;
wire n_1399;
wire n_1435;
wire n_969;
wire n_988;
wire n_1065;
wire n_1401;
wire n_1255;
wire n_568;
wire n_1516;
wire n_1536;
wire n_1204;
wire n_823;
wire n_1132;
wire n_643;
wire n_233;
wire n_698;
wire n_1074;
wire n_1394;
wire n_1327;
wire n_1326;
wire n_739;
wire n_400;
wire n_955;
wire n_337;
wire n_1379;
wire n_214;
wire n_246;
wire n_1338;
wire n_1097;
wire n_935;
wire n_781;
wire n_789;
wire n_1554;
wire n_1130;
wire n_1810;
wire n_573;
wire n_769;
wire n_676;
wire n_327;
wire n_1120;
wire n_832;
wire n_1583;
wire n_1730;
wire n_555;
wire n_389;
wire n_814;
wire n_1643;
wire n_1729;
wire n_669;
wire n_300;
wire n_222;
wire n_747;
wire n_1389;
wire n_1105;
wire n_721;
wire n_1461;
wire n_742;
wire n_535;
wire n_691;
wire n_372;
wire n_314;
wire n_1408;
wire n_378;
wire n_1196;
wire n_377;
wire n_1598;
wire n_863;
wire n_601;
wire n_338;
wire n_1283;
wire n_918;
wire n_748;
wire n_506;
wire n_1114;
wire n_1785;
wire n_763;
wire n_1147;
wire n_1848;
wire n_360;
wire n_1754;
wire n_1506;
wire n_1652;
wire n_1812;
wire n_957;
wire n_895;
wire n_866;
wire n_1227;
wire n_387;
wire n_452;
wire n_744;
wire n_971;
wire n_946;
wire n_344;
wire n_761;
wire n_1303;
wire n_1205;
wire n_1258;
wire n_1392;
wire n_1173;
wire n_1924;
wire n_525;
wire n_1677;
wire n_1116;
wire n_611;
wire n_1570;
wire n_1702;
wire n_1219;
wire n_1780;
wire n_1689;
wire n_1174;
wire n_1944;
wire n_1016;
wire n_1347;
wire n_795;
wire n_1501;
wire n_1221;
wire n_1245;
wire n_838;
wire n_647;
wire n_844;
wire n_448;
wire n_1017;
wire n_1083;
wire n_445;
wire n_1561;
wire n_930;
wire n_888;
wire n_1112;
wire n_234;
wire n_1945;
wire n_910;
wire n_1656;
wire n_1721;
wire n_1460;
wire n_911;
wire n_1464;
wire n_236;
wire n_653;
wire n_1737;
wire n_1414;
wire n_752;
wire n_908;
wire n_944;
wire n_576;
wire n_1028;
wire n_472;
wire n_270;
wire n_414;
wire n_1922;
wire n_563;
wire n_1011;
wire n_1566;
wire n_1215;
wire n_839;
wire n_708;
wire n_1973;
wire n_668;
wire n_626;
wire n_990;
wire n_1500;
wire n_779;
wire n_1537;
wire n_1821;
wire n_1104;
wire n_854;
wire n_1058;
wire n_498;
wire n_1122;
wire n_870;
wire n_904;
wire n_1253;
wire n_709;
wire n_1266;
wire n_366;
wire n_1509;
wire n_1693;
wire n_1109;
wire n_712;
wire n_348;
wire n_1276;
wire n_376;
wire n_390;
wire n_1148;
wire n_334;
wire n_1161;
wire n_1085;
wire n_232;
wire n_1239;
wire n_771;
wire n_1584;
wire n_470;
wire n_475;
wire n_924;
wire n_298;
wire n_1582;
wire n_492;
wire n_1149;
wire n_265;
wire n_1184;
wire n_228;
wire n_719;
wire n_1972;
wire n_1525;
wire n_455;
wire n_1585;
wire n_1851;
wire n_363;
wire n_1799;
wire n_1090;
wire n_592;
wire n_1816;
wire n_1518;
wire n_829;
wire n_1156;
wire n_1362;
wire n_393;
wire n_984;
wire n_1829;
wire n_503;
wire n_1450;
wire n_1638;
wire n_868;
wire n_570;
wire n_859;
wire n_406;
wire n_735;
wire n_1789;
wire n_1770;
wire n_878;
wire n_620;
wire n_519;
wire n_307;
wire n_469;
wire n_1218;
wire n_500;
wire n_1482;
wire n_981;
wire n_714;
wire n_1349;
wire n_291;
wire n_1144;
wire n_357;
wire n_985;
wire n_481;
wire n_997;
wire n_1710;
wire n_1301;
wire n_802;
wire n_561;
wire n_980;
wire n_1306;
wire n_1651;
wire n_1198;
wire n_1609;
wire n_436;
wire n_409;
wire n_1244;
wire n_1685;
wire n_1763;
wire n_1574;
wire n_240;
wire n_756;
wire n_1619;
wire n_1606;
wire n_810;
wire n_1133;
wire n_635;
wire n_1194;
wire n_1051;
wire n_253;
wire n_1552;
wire n_583;
wire n_249;
wire n_1039;
wire n_1442;
wire n_1034;
wire n_1480;
wire n_1158;
wire n_754;
wire n_941;
wire n_975;
wire n_1031;
wire n_1305;
wire n_553;
wire n_849;
wire n_753;
wire n_1753;
wire n_467;
wire n_269;
wire n_359;
wire n_973;
wire n_1921;
wire n_1479;
wire n_1055;
wire n_1675;
wire n_582;
wire n_861;
wire n_857;
wire n_967;
wire n_571;
wire n_404;
wire n_271;
wire n_1884;
wire n_679;
wire n_633;
wire n_1170;
wire n_665;
wire n_1629;
wire n_588;
wire n_225;
wire n_1260;
wire n_308;
wire n_309;
wire n_1819;
wire n_1010;
wire n_1040;
wire n_915;
wire n_632;
wire n_1166;
wire n_812;
wire n_1131;
wire n_1761;
wire n_534;
wire n_1578;
wire n_1006;
wire n_1861;
wire n_373;
wire n_1632;
wire n_1890;
wire n_1805;
wire n_257;
wire n_1557;
wire n_1888;
wire n_1833;
wire n_730;
wire n_1311;
wire n_1494;
wire n_670;
wire n_1850;
wire n_1898;
wire n_1868;
wire n_1089;
wire n_1887;
wire n_1587;
wire n_1365;
wire n_1417;
wire n_1242;
wire n_1836;
wire n_681;
wire n_1226;
wire n_1274;
wire n_1486;
wire n_412;
wire n_640;
wire n_1322;
wire n_965;
wire n_1899;
wire n_1428;
wire n_1616;
wire n_1576;
wire n_1862;
wire n_1856;
wire n_1958;
wire n_339;
wire n_784;
wire n_434;
wire n_315;
wire n_288;
wire n_1059;
wire n_1197;
wire n_422;
wire n_722;
wire n_862;
wire n_540;
wire n_1423;
wire n_1935;
wire n_457;
wire n_364;
wire n_1915;
wire n_629;
wire n_1621;
wire n_1748;
wire n_900;
wire n_1449;
wire n_531;
wire n_827;
wire n_361;
wire n_1025;
wire n_336;
wire n_1885;
wire n_1013;
wire n_1259;
wire n_1538;
wire n_649;
wire n_1612;
wire n_1240;

CKINVDCx5p33_ASAP7_75t_R g210 ( 
.A(n_100),
.Y(n_210)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_182),
.Y(n_211)
);

CKINVDCx5p33_ASAP7_75t_R g212 ( 
.A(n_71),
.Y(n_212)
);

CKINVDCx5p33_ASAP7_75t_R g213 ( 
.A(n_0),
.Y(n_213)
);

CKINVDCx20_ASAP7_75t_R g214 ( 
.A(n_16),
.Y(n_214)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_87),
.Y(n_215)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_52),
.Y(n_216)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_90),
.Y(n_217)
);

CKINVDCx5p33_ASAP7_75t_R g218 ( 
.A(n_207),
.Y(n_218)
);

INVx2_ASAP7_75t_L g219 ( 
.A(n_54),
.Y(n_219)
);

CKINVDCx5p33_ASAP7_75t_R g220 ( 
.A(n_53),
.Y(n_220)
);

BUFx6f_ASAP7_75t_L g221 ( 
.A(n_57),
.Y(n_221)
);

INVx2_ASAP7_75t_L g222 ( 
.A(n_74),
.Y(n_222)
);

CKINVDCx5p33_ASAP7_75t_R g223 ( 
.A(n_181),
.Y(n_223)
);

CKINVDCx5p33_ASAP7_75t_R g224 ( 
.A(n_111),
.Y(n_224)
);

CKINVDCx5p33_ASAP7_75t_R g225 ( 
.A(n_195),
.Y(n_225)
);

CKINVDCx5p33_ASAP7_75t_R g226 ( 
.A(n_67),
.Y(n_226)
);

CKINVDCx5p33_ASAP7_75t_R g227 ( 
.A(n_80),
.Y(n_227)
);

CKINVDCx5p33_ASAP7_75t_R g228 ( 
.A(n_143),
.Y(n_228)
);

CKINVDCx5p33_ASAP7_75t_R g229 ( 
.A(n_179),
.Y(n_229)
);

CKINVDCx5p33_ASAP7_75t_R g230 ( 
.A(n_96),
.Y(n_230)
);

INVx2_ASAP7_75t_L g231 ( 
.A(n_89),
.Y(n_231)
);

CKINVDCx5p33_ASAP7_75t_R g232 ( 
.A(n_165),
.Y(n_232)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_159),
.Y(n_233)
);

CKINVDCx5p33_ASAP7_75t_R g234 ( 
.A(n_156),
.Y(n_234)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_92),
.Y(n_235)
);

INVx1_ASAP7_75t_SL g236 ( 
.A(n_180),
.Y(n_236)
);

CKINVDCx5p33_ASAP7_75t_R g237 ( 
.A(n_185),
.Y(n_237)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_99),
.Y(n_238)
);

CKINVDCx5p33_ASAP7_75t_R g239 ( 
.A(n_164),
.Y(n_239)
);

INVx2_ASAP7_75t_L g240 ( 
.A(n_57),
.Y(n_240)
);

CKINVDCx5p33_ASAP7_75t_R g241 ( 
.A(n_79),
.Y(n_241)
);

CKINVDCx5p33_ASAP7_75t_R g242 ( 
.A(n_128),
.Y(n_242)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_101),
.Y(n_243)
);

CKINVDCx5p33_ASAP7_75t_R g244 ( 
.A(n_161),
.Y(n_244)
);

INVx2_ASAP7_75t_L g245 ( 
.A(n_201),
.Y(n_245)
);

CKINVDCx5p33_ASAP7_75t_R g246 ( 
.A(n_98),
.Y(n_246)
);

INVx1_ASAP7_75t_SL g247 ( 
.A(n_162),
.Y(n_247)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_64),
.Y(n_248)
);

CKINVDCx5p33_ASAP7_75t_R g249 ( 
.A(n_6),
.Y(n_249)
);

CKINVDCx5p33_ASAP7_75t_R g250 ( 
.A(n_86),
.Y(n_250)
);

HB1xp67_ASAP7_75t_L g251 ( 
.A(n_37),
.Y(n_251)
);

CKINVDCx5p33_ASAP7_75t_R g252 ( 
.A(n_91),
.Y(n_252)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_103),
.Y(n_253)
);

CKINVDCx5p33_ASAP7_75t_R g254 ( 
.A(n_83),
.Y(n_254)
);

INVx2_ASAP7_75t_L g255 ( 
.A(n_157),
.Y(n_255)
);

BUFx3_ASAP7_75t_L g256 ( 
.A(n_85),
.Y(n_256)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_48),
.Y(n_257)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_15),
.Y(n_258)
);

BUFx10_ASAP7_75t_L g259 ( 
.A(n_30),
.Y(n_259)
);

CKINVDCx5p33_ASAP7_75t_R g260 ( 
.A(n_123),
.Y(n_260)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_39),
.Y(n_261)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_134),
.Y(n_262)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_29),
.Y(n_263)
);

CKINVDCx5p33_ASAP7_75t_R g264 ( 
.A(n_55),
.Y(n_264)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_137),
.Y(n_265)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_112),
.Y(n_266)
);

CKINVDCx5p33_ASAP7_75t_R g267 ( 
.A(n_142),
.Y(n_267)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_78),
.Y(n_268)
);

BUFx6f_ASAP7_75t_L g269 ( 
.A(n_19),
.Y(n_269)
);

CKINVDCx20_ASAP7_75t_R g270 ( 
.A(n_202),
.Y(n_270)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_7),
.Y(n_271)
);

INVx2_ASAP7_75t_SL g272 ( 
.A(n_65),
.Y(n_272)
);

CKINVDCx5p33_ASAP7_75t_R g273 ( 
.A(n_38),
.Y(n_273)
);

CKINVDCx5p33_ASAP7_75t_R g274 ( 
.A(n_43),
.Y(n_274)
);

INVx2_ASAP7_75t_L g275 ( 
.A(n_146),
.Y(n_275)
);

CKINVDCx5p33_ASAP7_75t_R g276 ( 
.A(n_94),
.Y(n_276)
);

CKINVDCx5p33_ASAP7_75t_R g277 ( 
.A(n_3),
.Y(n_277)
);

CKINVDCx5p33_ASAP7_75t_R g278 ( 
.A(n_51),
.Y(n_278)
);

CKINVDCx20_ASAP7_75t_R g279 ( 
.A(n_204),
.Y(n_279)
);

CKINVDCx5p33_ASAP7_75t_R g280 ( 
.A(n_132),
.Y(n_280)
);

CKINVDCx5p33_ASAP7_75t_R g281 ( 
.A(n_42),
.Y(n_281)
);

CKINVDCx5p33_ASAP7_75t_R g282 ( 
.A(n_194),
.Y(n_282)
);

BUFx10_ASAP7_75t_L g283 ( 
.A(n_23),
.Y(n_283)
);

CKINVDCx5p33_ASAP7_75t_R g284 ( 
.A(n_63),
.Y(n_284)
);

BUFx10_ASAP7_75t_L g285 ( 
.A(n_135),
.Y(n_285)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_205),
.Y(n_286)
);

CKINVDCx5p33_ASAP7_75t_R g287 ( 
.A(n_84),
.Y(n_287)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_44),
.Y(n_288)
);

CKINVDCx5p33_ASAP7_75t_R g289 ( 
.A(n_51),
.Y(n_289)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_7),
.Y(n_290)
);

CKINVDCx20_ASAP7_75t_R g291 ( 
.A(n_47),
.Y(n_291)
);

CKINVDCx5p33_ASAP7_75t_R g292 ( 
.A(n_77),
.Y(n_292)
);

HB1xp67_ASAP7_75t_L g293 ( 
.A(n_196),
.Y(n_293)
);

BUFx8_ASAP7_75t_SL g294 ( 
.A(n_174),
.Y(n_294)
);

INVx1_ASAP7_75t_SL g295 ( 
.A(n_109),
.Y(n_295)
);

INVx2_ASAP7_75t_SL g296 ( 
.A(n_38),
.Y(n_296)
);

CKINVDCx5p33_ASAP7_75t_R g297 ( 
.A(n_170),
.Y(n_297)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_141),
.Y(n_298)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_151),
.Y(n_299)
);

INVx1_ASAP7_75t_SL g300 ( 
.A(n_187),
.Y(n_300)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_198),
.Y(n_301)
);

CKINVDCx5p33_ASAP7_75t_R g302 ( 
.A(n_155),
.Y(n_302)
);

CKINVDCx5p33_ASAP7_75t_R g303 ( 
.A(n_62),
.Y(n_303)
);

CKINVDCx5p33_ASAP7_75t_R g304 ( 
.A(n_48),
.Y(n_304)
);

CKINVDCx5p33_ASAP7_75t_R g305 ( 
.A(n_102),
.Y(n_305)
);

INVx2_ASAP7_75t_L g306 ( 
.A(n_24),
.Y(n_306)
);

CKINVDCx5p33_ASAP7_75t_R g307 ( 
.A(n_36),
.Y(n_307)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_54),
.Y(n_308)
);

INVx2_ASAP7_75t_SL g309 ( 
.A(n_150),
.Y(n_309)
);

HB1xp67_ASAP7_75t_L g310 ( 
.A(n_158),
.Y(n_310)
);

CKINVDCx5p33_ASAP7_75t_R g311 ( 
.A(n_183),
.Y(n_311)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_148),
.Y(n_312)
);

BUFx6f_ASAP7_75t_L g313 ( 
.A(n_175),
.Y(n_313)
);

CKINVDCx5p33_ASAP7_75t_R g314 ( 
.A(n_61),
.Y(n_314)
);

CKINVDCx5p33_ASAP7_75t_R g315 ( 
.A(n_163),
.Y(n_315)
);

CKINVDCx5p33_ASAP7_75t_R g316 ( 
.A(n_208),
.Y(n_316)
);

CKINVDCx5p33_ASAP7_75t_R g317 ( 
.A(n_177),
.Y(n_317)
);

CKINVDCx5p33_ASAP7_75t_R g318 ( 
.A(n_76),
.Y(n_318)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_172),
.Y(n_319)
);

CKINVDCx5p33_ASAP7_75t_R g320 ( 
.A(n_115),
.Y(n_320)
);

CKINVDCx5p33_ASAP7_75t_R g321 ( 
.A(n_88),
.Y(n_321)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_118),
.Y(n_322)
);

INVx1_ASAP7_75t_SL g323 ( 
.A(n_152),
.Y(n_323)
);

BUFx6f_ASAP7_75t_L g324 ( 
.A(n_160),
.Y(n_324)
);

CKINVDCx5p33_ASAP7_75t_R g325 ( 
.A(n_34),
.Y(n_325)
);

BUFx6f_ASAP7_75t_L g326 ( 
.A(n_27),
.Y(n_326)
);

INVx1_ASAP7_75t_SL g327 ( 
.A(n_28),
.Y(n_327)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_22),
.Y(n_328)
);

CKINVDCx20_ASAP7_75t_R g329 ( 
.A(n_144),
.Y(n_329)
);

CKINVDCx5p33_ASAP7_75t_R g330 ( 
.A(n_178),
.Y(n_330)
);

INVx1_ASAP7_75t_SL g331 ( 
.A(n_121),
.Y(n_331)
);

CKINVDCx5p33_ASAP7_75t_R g332 ( 
.A(n_139),
.Y(n_332)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_81),
.Y(n_333)
);

CKINVDCx16_ASAP7_75t_R g334 ( 
.A(n_116),
.Y(n_334)
);

CKINVDCx5p33_ASAP7_75t_R g335 ( 
.A(n_43),
.Y(n_335)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_131),
.Y(n_336)
);

CKINVDCx5p33_ASAP7_75t_R g337 ( 
.A(n_136),
.Y(n_337)
);

INVx1_ASAP7_75t_L g338 ( 
.A(n_0),
.Y(n_338)
);

CKINVDCx5p33_ASAP7_75t_R g339 ( 
.A(n_107),
.Y(n_339)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_29),
.Y(n_340)
);

CKINVDCx5p33_ASAP7_75t_R g341 ( 
.A(n_140),
.Y(n_341)
);

CKINVDCx5p33_ASAP7_75t_R g342 ( 
.A(n_10),
.Y(n_342)
);

CKINVDCx5p33_ASAP7_75t_R g343 ( 
.A(n_120),
.Y(n_343)
);

INVx1_ASAP7_75t_L g344 ( 
.A(n_93),
.Y(n_344)
);

HB1xp67_ASAP7_75t_L g345 ( 
.A(n_40),
.Y(n_345)
);

CKINVDCx5p33_ASAP7_75t_R g346 ( 
.A(n_56),
.Y(n_346)
);

CKINVDCx5p33_ASAP7_75t_R g347 ( 
.A(n_44),
.Y(n_347)
);

INVx1_ASAP7_75t_L g348 ( 
.A(n_2),
.Y(n_348)
);

CKINVDCx5p33_ASAP7_75t_R g349 ( 
.A(n_73),
.Y(n_349)
);

CKINVDCx5p33_ASAP7_75t_R g350 ( 
.A(n_129),
.Y(n_350)
);

CKINVDCx5p33_ASAP7_75t_R g351 ( 
.A(n_3),
.Y(n_351)
);

CKINVDCx5p33_ASAP7_75t_R g352 ( 
.A(n_19),
.Y(n_352)
);

CKINVDCx5p33_ASAP7_75t_R g353 ( 
.A(n_133),
.Y(n_353)
);

INVx1_ASAP7_75t_L g354 ( 
.A(n_11),
.Y(n_354)
);

INVx1_ASAP7_75t_L g355 ( 
.A(n_70),
.Y(n_355)
);

INVx2_ASAP7_75t_L g356 ( 
.A(n_190),
.Y(n_356)
);

HB1xp67_ASAP7_75t_L g357 ( 
.A(n_82),
.Y(n_357)
);

CKINVDCx5p33_ASAP7_75t_R g358 ( 
.A(n_16),
.Y(n_358)
);

CKINVDCx5p33_ASAP7_75t_R g359 ( 
.A(n_49),
.Y(n_359)
);

BUFx5_ASAP7_75t_L g360 ( 
.A(n_125),
.Y(n_360)
);

INVx1_ASAP7_75t_L g361 ( 
.A(n_153),
.Y(n_361)
);

CKINVDCx5p33_ASAP7_75t_R g362 ( 
.A(n_122),
.Y(n_362)
);

INVx1_ASAP7_75t_L g363 ( 
.A(n_33),
.Y(n_363)
);

INVx1_ASAP7_75t_L g364 ( 
.A(n_199),
.Y(n_364)
);

CKINVDCx5p33_ASAP7_75t_R g365 ( 
.A(n_31),
.Y(n_365)
);

INVx1_ASAP7_75t_L g366 ( 
.A(n_104),
.Y(n_366)
);

INVx1_ASAP7_75t_L g367 ( 
.A(n_23),
.Y(n_367)
);

CKINVDCx5p33_ASAP7_75t_R g368 ( 
.A(n_18),
.Y(n_368)
);

CKINVDCx5p33_ASAP7_75t_R g369 ( 
.A(n_188),
.Y(n_369)
);

CKINVDCx5p33_ASAP7_75t_R g370 ( 
.A(n_30),
.Y(n_370)
);

CKINVDCx5p33_ASAP7_75t_R g371 ( 
.A(n_56),
.Y(n_371)
);

INVx1_ASAP7_75t_L g372 ( 
.A(n_72),
.Y(n_372)
);

BUFx2_ASAP7_75t_L g373 ( 
.A(n_49),
.Y(n_373)
);

CKINVDCx5p33_ASAP7_75t_R g374 ( 
.A(n_110),
.Y(n_374)
);

CKINVDCx5p33_ASAP7_75t_R g375 ( 
.A(n_192),
.Y(n_375)
);

CKINVDCx5p33_ASAP7_75t_R g376 ( 
.A(n_14),
.Y(n_376)
);

INVx1_ASAP7_75t_SL g377 ( 
.A(n_127),
.Y(n_377)
);

BUFx3_ASAP7_75t_L g378 ( 
.A(n_28),
.Y(n_378)
);

CKINVDCx5p33_ASAP7_75t_R g379 ( 
.A(n_11),
.Y(n_379)
);

INVx1_ASAP7_75t_L g380 ( 
.A(n_75),
.Y(n_380)
);

CKINVDCx5p33_ASAP7_75t_R g381 ( 
.A(n_169),
.Y(n_381)
);

CKINVDCx20_ASAP7_75t_R g382 ( 
.A(n_95),
.Y(n_382)
);

INVx1_ASAP7_75t_L g383 ( 
.A(n_18),
.Y(n_383)
);

CKINVDCx5p33_ASAP7_75t_R g384 ( 
.A(n_138),
.Y(n_384)
);

INVx1_ASAP7_75t_L g385 ( 
.A(n_47),
.Y(n_385)
);

CKINVDCx5p33_ASAP7_75t_R g386 ( 
.A(n_147),
.Y(n_386)
);

INVx1_ASAP7_75t_L g387 ( 
.A(n_45),
.Y(n_387)
);

CKINVDCx20_ASAP7_75t_R g388 ( 
.A(n_68),
.Y(n_388)
);

INVx1_ASAP7_75t_L g389 ( 
.A(n_32),
.Y(n_389)
);

CKINVDCx20_ASAP7_75t_R g390 ( 
.A(n_130),
.Y(n_390)
);

INVx1_ASAP7_75t_L g391 ( 
.A(n_113),
.Y(n_391)
);

INVx1_ASAP7_75t_L g392 ( 
.A(n_191),
.Y(n_392)
);

CKINVDCx20_ASAP7_75t_R g393 ( 
.A(n_119),
.Y(n_393)
);

BUFx2_ASAP7_75t_L g394 ( 
.A(n_189),
.Y(n_394)
);

BUFx10_ASAP7_75t_L g395 ( 
.A(n_45),
.Y(n_395)
);

INVx1_ASAP7_75t_L g396 ( 
.A(n_53),
.Y(n_396)
);

INVx1_ASAP7_75t_L g397 ( 
.A(n_106),
.Y(n_397)
);

CKINVDCx5p33_ASAP7_75t_R g398 ( 
.A(n_1),
.Y(n_398)
);

CKINVDCx5p33_ASAP7_75t_R g399 ( 
.A(n_117),
.Y(n_399)
);

CKINVDCx5p33_ASAP7_75t_R g400 ( 
.A(n_114),
.Y(n_400)
);

CKINVDCx5p33_ASAP7_75t_R g401 ( 
.A(n_176),
.Y(n_401)
);

CKINVDCx5p33_ASAP7_75t_R g402 ( 
.A(n_26),
.Y(n_402)
);

CKINVDCx20_ASAP7_75t_R g403 ( 
.A(n_203),
.Y(n_403)
);

CKINVDCx20_ASAP7_75t_R g404 ( 
.A(n_173),
.Y(n_404)
);

INVx1_ASAP7_75t_L g405 ( 
.A(n_66),
.Y(n_405)
);

INVx1_ASAP7_75t_L g406 ( 
.A(n_27),
.Y(n_406)
);

INVx1_ASAP7_75t_L g407 ( 
.A(n_168),
.Y(n_407)
);

CKINVDCx20_ASAP7_75t_R g408 ( 
.A(n_22),
.Y(n_408)
);

CKINVDCx20_ASAP7_75t_R g409 ( 
.A(n_50),
.Y(n_409)
);

CKINVDCx5p33_ASAP7_75t_R g410 ( 
.A(n_25),
.Y(n_410)
);

CKINVDCx5p33_ASAP7_75t_R g411 ( 
.A(n_55),
.Y(n_411)
);

CKINVDCx5p33_ASAP7_75t_R g412 ( 
.A(n_145),
.Y(n_412)
);

CKINVDCx5p33_ASAP7_75t_R g413 ( 
.A(n_200),
.Y(n_413)
);

INVx1_ASAP7_75t_L g414 ( 
.A(n_12),
.Y(n_414)
);

INVx2_ASAP7_75t_L g415 ( 
.A(n_8),
.Y(n_415)
);

INVx1_ASAP7_75t_L g416 ( 
.A(n_124),
.Y(n_416)
);

INVx1_ASAP7_75t_L g417 ( 
.A(n_154),
.Y(n_417)
);

INVx1_ASAP7_75t_L g418 ( 
.A(n_221),
.Y(n_418)
);

HB1xp67_ASAP7_75t_L g419 ( 
.A(n_251),
.Y(n_419)
);

HB1xp67_ASAP7_75t_L g420 ( 
.A(n_345),
.Y(n_420)
);

CKINVDCx20_ASAP7_75t_R g421 ( 
.A(n_270),
.Y(n_421)
);

INVx1_ASAP7_75t_L g422 ( 
.A(n_221),
.Y(n_422)
);

INVx1_ASAP7_75t_L g423 ( 
.A(n_378),
.Y(n_423)
);

INVxp67_ASAP7_75t_SL g424 ( 
.A(n_293),
.Y(n_424)
);

CKINVDCx5p33_ASAP7_75t_R g425 ( 
.A(n_249),
.Y(n_425)
);

CKINVDCx20_ASAP7_75t_R g426 ( 
.A(n_279),
.Y(n_426)
);

INVx1_ASAP7_75t_L g427 ( 
.A(n_378),
.Y(n_427)
);

CKINVDCx20_ASAP7_75t_R g428 ( 
.A(n_329),
.Y(n_428)
);

CKINVDCx16_ASAP7_75t_R g429 ( 
.A(n_334),
.Y(n_429)
);

CKINVDCx16_ASAP7_75t_R g430 ( 
.A(n_259),
.Y(n_430)
);

CKINVDCx20_ASAP7_75t_R g431 ( 
.A(n_382),
.Y(n_431)
);

CKINVDCx20_ASAP7_75t_R g432 ( 
.A(n_388),
.Y(n_432)
);

INVx1_ASAP7_75t_L g433 ( 
.A(n_221),
.Y(n_433)
);

CKINVDCx5p33_ASAP7_75t_R g434 ( 
.A(n_264),
.Y(n_434)
);

CKINVDCx16_ASAP7_75t_R g435 ( 
.A(n_259),
.Y(n_435)
);

INVx1_ASAP7_75t_L g436 ( 
.A(n_221),
.Y(n_436)
);

CKINVDCx20_ASAP7_75t_R g437 ( 
.A(n_390),
.Y(n_437)
);

CKINVDCx5p33_ASAP7_75t_R g438 ( 
.A(n_273),
.Y(n_438)
);

INVx1_ASAP7_75t_L g439 ( 
.A(n_221),
.Y(n_439)
);

CKINVDCx20_ASAP7_75t_R g440 ( 
.A(n_393),
.Y(n_440)
);

CKINVDCx20_ASAP7_75t_R g441 ( 
.A(n_403),
.Y(n_441)
);

CKINVDCx20_ASAP7_75t_R g442 ( 
.A(n_404),
.Y(n_442)
);

CKINVDCx20_ASAP7_75t_R g443 ( 
.A(n_294),
.Y(n_443)
);

INVx1_ASAP7_75t_L g444 ( 
.A(n_269),
.Y(n_444)
);

INVx1_ASAP7_75t_L g445 ( 
.A(n_269),
.Y(n_445)
);

INVxp33_ASAP7_75t_SL g446 ( 
.A(n_213),
.Y(n_446)
);

CKINVDCx20_ASAP7_75t_R g447 ( 
.A(n_210),
.Y(n_447)
);

INVx1_ASAP7_75t_L g448 ( 
.A(n_269),
.Y(n_448)
);

HB1xp67_ASAP7_75t_L g449 ( 
.A(n_373),
.Y(n_449)
);

INVx1_ASAP7_75t_L g450 ( 
.A(n_269),
.Y(n_450)
);

INVx1_ASAP7_75t_L g451 ( 
.A(n_269),
.Y(n_451)
);

INVx1_ASAP7_75t_L g452 ( 
.A(n_326),
.Y(n_452)
);

CKINVDCx5p33_ASAP7_75t_R g453 ( 
.A(n_274),
.Y(n_453)
);

CKINVDCx5p33_ASAP7_75t_R g454 ( 
.A(n_277),
.Y(n_454)
);

INVx2_ASAP7_75t_L g455 ( 
.A(n_326),
.Y(n_455)
);

BUFx3_ASAP7_75t_L g456 ( 
.A(n_256),
.Y(n_456)
);

INVxp67_ASAP7_75t_L g457 ( 
.A(n_259),
.Y(n_457)
);

CKINVDCx5p33_ASAP7_75t_R g458 ( 
.A(n_278),
.Y(n_458)
);

INVx1_ASAP7_75t_L g459 ( 
.A(n_326),
.Y(n_459)
);

INVx1_ASAP7_75t_L g460 ( 
.A(n_326),
.Y(n_460)
);

INVx1_ASAP7_75t_L g461 ( 
.A(n_326),
.Y(n_461)
);

CKINVDCx14_ASAP7_75t_R g462 ( 
.A(n_394),
.Y(n_462)
);

INVx1_ASAP7_75t_L g463 ( 
.A(n_216),
.Y(n_463)
);

CKINVDCx20_ASAP7_75t_R g464 ( 
.A(n_246),
.Y(n_464)
);

CKINVDCx5p33_ASAP7_75t_R g465 ( 
.A(n_281),
.Y(n_465)
);

INVxp33_ASAP7_75t_L g466 ( 
.A(n_257),
.Y(n_466)
);

CKINVDCx5p33_ASAP7_75t_R g467 ( 
.A(n_289),
.Y(n_467)
);

INVx1_ASAP7_75t_L g468 ( 
.A(n_258),
.Y(n_468)
);

INVx1_ASAP7_75t_L g469 ( 
.A(n_261),
.Y(n_469)
);

INVx1_ASAP7_75t_L g470 ( 
.A(n_263),
.Y(n_470)
);

INVx1_ASAP7_75t_L g471 ( 
.A(n_219),
.Y(n_471)
);

INVxp67_ASAP7_75t_SL g472 ( 
.A(n_310),
.Y(n_472)
);

INVx1_ASAP7_75t_L g473 ( 
.A(n_271),
.Y(n_473)
);

INVx1_ASAP7_75t_L g474 ( 
.A(n_288),
.Y(n_474)
);

HB1xp67_ASAP7_75t_L g475 ( 
.A(n_213),
.Y(n_475)
);

CKINVDCx5p33_ASAP7_75t_R g476 ( 
.A(n_304),
.Y(n_476)
);

CKINVDCx5p33_ASAP7_75t_R g477 ( 
.A(n_307),
.Y(n_477)
);

INVx1_ASAP7_75t_L g478 ( 
.A(n_290),
.Y(n_478)
);

INVxp67_ASAP7_75t_SL g479 ( 
.A(n_357),
.Y(n_479)
);

INVx1_ASAP7_75t_L g480 ( 
.A(n_308),
.Y(n_480)
);

INVxp67_ASAP7_75t_SL g481 ( 
.A(n_256),
.Y(n_481)
);

INVxp67_ASAP7_75t_SL g482 ( 
.A(n_211),
.Y(n_482)
);

BUFx2_ASAP7_75t_L g483 ( 
.A(n_220),
.Y(n_483)
);

INVx1_ASAP7_75t_L g484 ( 
.A(n_328),
.Y(n_484)
);

INVx1_ASAP7_75t_L g485 ( 
.A(n_338),
.Y(n_485)
);

CKINVDCx20_ASAP7_75t_R g486 ( 
.A(n_250),
.Y(n_486)
);

INVxp67_ASAP7_75t_L g487 ( 
.A(n_283),
.Y(n_487)
);

CKINVDCx20_ASAP7_75t_R g488 ( 
.A(n_252),
.Y(n_488)
);

INVx1_ASAP7_75t_L g489 ( 
.A(n_340),
.Y(n_489)
);

INVx1_ASAP7_75t_L g490 ( 
.A(n_348),
.Y(n_490)
);

INVx1_ASAP7_75t_L g491 ( 
.A(n_354),
.Y(n_491)
);

CKINVDCx16_ASAP7_75t_R g492 ( 
.A(n_283),
.Y(n_492)
);

CKINVDCx20_ASAP7_75t_R g493 ( 
.A(n_254),
.Y(n_493)
);

HB1xp67_ASAP7_75t_L g494 ( 
.A(n_220),
.Y(n_494)
);

CKINVDCx16_ASAP7_75t_R g495 ( 
.A(n_283),
.Y(n_495)
);

INVxp67_ASAP7_75t_SL g496 ( 
.A(n_215),
.Y(n_496)
);

CKINVDCx5p33_ASAP7_75t_R g497 ( 
.A(n_325),
.Y(n_497)
);

INVx1_ASAP7_75t_L g498 ( 
.A(n_363),
.Y(n_498)
);

INVx1_ASAP7_75t_L g499 ( 
.A(n_219),
.Y(n_499)
);

INVx1_ASAP7_75t_L g500 ( 
.A(n_240),
.Y(n_500)
);

INVxp33_ASAP7_75t_SL g501 ( 
.A(n_376),
.Y(n_501)
);

INVx1_ASAP7_75t_SL g502 ( 
.A(n_214),
.Y(n_502)
);

INVxp67_ASAP7_75t_SL g503 ( 
.A(n_217),
.Y(n_503)
);

CKINVDCx5p33_ASAP7_75t_R g504 ( 
.A(n_335),
.Y(n_504)
);

CKINVDCx5p33_ASAP7_75t_R g505 ( 
.A(n_342),
.Y(n_505)
);

INVx1_ASAP7_75t_L g506 ( 
.A(n_240),
.Y(n_506)
);

INVx1_ASAP7_75t_L g507 ( 
.A(n_306),
.Y(n_507)
);

INVx1_ASAP7_75t_L g508 ( 
.A(n_306),
.Y(n_508)
);

INVx1_ASAP7_75t_L g509 ( 
.A(n_415),
.Y(n_509)
);

INVx1_ASAP7_75t_L g510 ( 
.A(n_415),
.Y(n_510)
);

CKINVDCx5p33_ASAP7_75t_R g511 ( 
.A(n_346),
.Y(n_511)
);

INVx1_ASAP7_75t_L g512 ( 
.A(n_367),
.Y(n_512)
);

INVx2_ASAP7_75t_L g513 ( 
.A(n_360),
.Y(n_513)
);

CKINVDCx20_ASAP7_75t_R g514 ( 
.A(n_260),
.Y(n_514)
);

CKINVDCx5p33_ASAP7_75t_R g515 ( 
.A(n_347),
.Y(n_515)
);

CKINVDCx16_ASAP7_75t_R g516 ( 
.A(n_395),
.Y(n_516)
);

HB1xp67_ASAP7_75t_L g517 ( 
.A(n_376),
.Y(n_517)
);

INVx2_ASAP7_75t_L g518 ( 
.A(n_360),
.Y(n_518)
);

CKINVDCx20_ASAP7_75t_R g519 ( 
.A(n_267),
.Y(n_519)
);

INVx1_ASAP7_75t_L g520 ( 
.A(n_383),
.Y(n_520)
);

INVxp67_ASAP7_75t_SL g521 ( 
.A(n_233),
.Y(n_521)
);

HB1xp67_ASAP7_75t_L g522 ( 
.A(n_379),
.Y(n_522)
);

CKINVDCx5p33_ASAP7_75t_R g523 ( 
.A(n_351),
.Y(n_523)
);

INVxp67_ASAP7_75t_SL g524 ( 
.A(n_235),
.Y(n_524)
);

INVx1_ASAP7_75t_L g525 ( 
.A(n_418),
.Y(n_525)
);

NAND2xp5_ASAP7_75t_L g526 ( 
.A(n_481),
.B(n_272),
.Y(n_526)
);

BUFx3_ASAP7_75t_L g527 ( 
.A(n_456),
.Y(n_527)
);

INVx2_ASAP7_75t_L g528 ( 
.A(n_455),
.Y(n_528)
);

INVx1_ASAP7_75t_L g529 ( 
.A(n_418),
.Y(n_529)
);

INVx1_ASAP7_75t_L g530 ( 
.A(n_422),
.Y(n_530)
);

CKINVDCx5p33_ASAP7_75t_R g531 ( 
.A(n_443),
.Y(n_531)
);

NAND2xp5_ASAP7_75t_L g532 ( 
.A(n_482),
.B(n_272),
.Y(n_532)
);

INVx1_ASAP7_75t_L g533 ( 
.A(n_422),
.Y(n_533)
);

INVx1_ASAP7_75t_L g534 ( 
.A(n_433),
.Y(n_534)
);

INVx2_ASAP7_75t_L g535 ( 
.A(n_455),
.Y(n_535)
);

INVxp67_ASAP7_75t_L g536 ( 
.A(n_475),
.Y(n_536)
);

INVx1_ASAP7_75t_L g537 ( 
.A(n_433),
.Y(n_537)
);

NAND2xp5_ASAP7_75t_SL g538 ( 
.A(n_429),
.B(n_285),
.Y(n_538)
);

HB1xp67_ASAP7_75t_L g539 ( 
.A(n_425),
.Y(n_539)
);

BUFx6f_ASAP7_75t_L g540 ( 
.A(n_436),
.Y(n_540)
);

BUFx8_ASAP7_75t_L g541 ( 
.A(n_483),
.Y(n_541)
);

BUFx6f_ASAP7_75t_L g542 ( 
.A(n_436),
.Y(n_542)
);

NAND2xp5_ASAP7_75t_L g543 ( 
.A(n_496),
.B(n_309),
.Y(n_543)
);

INVx1_ASAP7_75t_L g544 ( 
.A(n_439),
.Y(n_544)
);

AND2x2_ASAP7_75t_L g545 ( 
.A(n_456),
.B(n_296),
.Y(n_545)
);

AND2x2_ASAP7_75t_L g546 ( 
.A(n_423),
.B(n_427),
.Y(n_546)
);

AND2x2_ASAP7_75t_L g547 ( 
.A(n_503),
.B(n_296),
.Y(n_547)
);

INVx1_ASAP7_75t_L g548 ( 
.A(n_439),
.Y(n_548)
);

NAND2xp5_ASAP7_75t_L g549 ( 
.A(n_521),
.B(n_309),
.Y(n_549)
);

BUFx6f_ASAP7_75t_L g550 ( 
.A(n_444),
.Y(n_550)
);

NAND2xp5_ASAP7_75t_L g551 ( 
.A(n_524),
.B(n_222),
.Y(n_551)
);

AND2x6_ASAP7_75t_L g552 ( 
.A(n_513),
.B(n_313),
.Y(n_552)
);

AND2x2_ASAP7_75t_L g553 ( 
.A(n_424),
.B(n_285),
.Y(n_553)
);

INVx1_ASAP7_75t_L g554 ( 
.A(n_444),
.Y(n_554)
);

AND2x4_ASAP7_75t_L g555 ( 
.A(n_445),
.B(n_222),
.Y(n_555)
);

BUFx8_ASAP7_75t_L g556 ( 
.A(n_483),
.Y(n_556)
);

INVx1_ASAP7_75t_L g557 ( 
.A(n_445),
.Y(n_557)
);

AND2x2_ASAP7_75t_L g558 ( 
.A(n_472),
.B(n_285),
.Y(n_558)
);

INVx1_ASAP7_75t_L g559 ( 
.A(n_448),
.Y(n_559)
);

NAND2xp5_ASAP7_75t_L g560 ( 
.A(n_479),
.B(n_231),
.Y(n_560)
);

INVx2_ASAP7_75t_L g561 ( 
.A(n_448),
.Y(n_561)
);

INVx4_ASAP7_75t_L g562 ( 
.A(n_513),
.Y(n_562)
);

NAND2xp5_ASAP7_75t_L g563 ( 
.A(n_462),
.B(n_231),
.Y(n_563)
);

AND2x2_ASAP7_75t_L g564 ( 
.A(n_463),
.B(n_385),
.Y(n_564)
);

INVx6_ASAP7_75t_L g565 ( 
.A(n_459),
.Y(n_565)
);

AND2x6_ASAP7_75t_L g566 ( 
.A(n_518),
.B(n_313),
.Y(n_566)
);

AND2x4_ASAP7_75t_L g567 ( 
.A(n_450),
.B(n_245),
.Y(n_567)
);

INVx1_ASAP7_75t_L g568 ( 
.A(n_450),
.Y(n_568)
);

NOR2xp33_ASAP7_75t_R g569 ( 
.A(n_447),
.B(n_276),
.Y(n_569)
);

INVx3_ASAP7_75t_L g570 ( 
.A(n_518),
.Y(n_570)
);

HB1xp67_ASAP7_75t_L g571 ( 
.A(n_425),
.Y(n_571)
);

XOR2x2_ASAP7_75t_L g572 ( 
.A(n_502),
.B(n_327),
.Y(n_572)
);

HB1xp67_ASAP7_75t_L g573 ( 
.A(n_434),
.Y(n_573)
);

INVx3_ASAP7_75t_L g574 ( 
.A(n_451),
.Y(n_574)
);

BUFx2_ASAP7_75t_L g575 ( 
.A(n_434),
.Y(n_575)
);

CKINVDCx8_ASAP7_75t_R g576 ( 
.A(n_430),
.Y(n_576)
);

INVx1_ASAP7_75t_L g577 ( 
.A(n_451),
.Y(n_577)
);

CKINVDCx20_ASAP7_75t_R g578 ( 
.A(n_421),
.Y(n_578)
);

NAND2xp5_ASAP7_75t_L g579 ( 
.A(n_460),
.B(n_461),
.Y(n_579)
);

INVx3_ASAP7_75t_L g580 ( 
.A(n_452),
.Y(n_580)
);

BUFx6f_ASAP7_75t_L g581 ( 
.A(n_452),
.Y(n_581)
);

INVx2_ASAP7_75t_L g582 ( 
.A(n_471),
.Y(n_582)
);

INVx1_ASAP7_75t_L g583 ( 
.A(n_512),
.Y(n_583)
);

AND2x2_ASAP7_75t_L g584 ( 
.A(n_468),
.B(n_387),
.Y(n_584)
);

INVx1_ASAP7_75t_L g585 ( 
.A(n_512),
.Y(n_585)
);

CKINVDCx5p33_ASAP7_75t_R g586 ( 
.A(n_464),
.Y(n_586)
);

INVx1_ASAP7_75t_L g587 ( 
.A(n_520),
.Y(n_587)
);

INVx2_ASAP7_75t_L g588 ( 
.A(n_471),
.Y(n_588)
);

AND2x2_ASAP7_75t_L g589 ( 
.A(n_469),
.B(n_389),
.Y(n_589)
);

CKINVDCx16_ASAP7_75t_R g590 ( 
.A(n_435),
.Y(n_590)
);

CKINVDCx16_ASAP7_75t_R g591 ( 
.A(n_492),
.Y(n_591)
);

INVx2_ASAP7_75t_L g592 ( 
.A(n_499),
.Y(n_592)
);

BUFx6f_ASAP7_75t_L g593 ( 
.A(n_499),
.Y(n_593)
);

INVx1_ASAP7_75t_L g594 ( 
.A(n_520),
.Y(n_594)
);

CKINVDCx20_ASAP7_75t_R g595 ( 
.A(n_426),
.Y(n_595)
);

CKINVDCx5p33_ASAP7_75t_R g596 ( 
.A(n_486),
.Y(n_596)
);

AND2x2_ASAP7_75t_L g597 ( 
.A(n_470),
.B(n_396),
.Y(n_597)
);

BUFx3_ASAP7_75t_L g598 ( 
.A(n_473),
.Y(n_598)
);

NOR2xp33_ASAP7_75t_L g599 ( 
.A(n_446),
.B(n_236),
.Y(n_599)
);

OAI22xp5_ASAP7_75t_SL g600 ( 
.A1(n_495),
.A2(n_408),
.B1(n_291),
.B2(n_409),
.Y(n_600)
);

NAND2xp5_ASAP7_75t_L g601 ( 
.A(n_523),
.B(n_438),
.Y(n_601)
);

INVx2_ASAP7_75t_L g602 ( 
.A(n_500),
.Y(n_602)
);

INVx3_ASAP7_75t_L g603 ( 
.A(n_500),
.Y(n_603)
);

INVx1_ASAP7_75t_L g604 ( 
.A(n_506),
.Y(n_604)
);

INVx3_ASAP7_75t_L g605 ( 
.A(n_506),
.Y(n_605)
);

INVx1_ASAP7_75t_L g606 ( 
.A(n_507),
.Y(n_606)
);

INVx1_ASAP7_75t_L g607 ( 
.A(n_507),
.Y(n_607)
);

INVx2_ASAP7_75t_L g608 ( 
.A(n_508),
.Y(n_608)
);

INVx1_ASAP7_75t_L g609 ( 
.A(n_508),
.Y(n_609)
);

INVx3_ASAP7_75t_L g610 ( 
.A(n_562),
.Y(n_610)
);

AND2x2_ASAP7_75t_L g611 ( 
.A(n_547),
.B(n_509),
.Y(n_611)
);

NOR2xp33_ASAP7_75t_L g612 ( 
.A(n_599),
.B(n_501),
.Y(n_612)
);

AND2x4_ASAP7_75t_L g613 ( 
.A(n_527),
.B(n_474),
.Y(n_613)
);

INVx3_ASAP7_75t_L g614 ( 
.A(n_562),
.Y(n_614)
);

INVx2_ASAP7_75t_L g615 ( 
.A(n_528),
.Y(n_615)
);

BUFx6f_ASAP7_75t_L g616 ( 
.A(n_540),
.Y(n_616)
);

INVx3_ASAP7_75t_L g617 ( 
.A(n_562),
.Y(n_617)
);

INVx2_ASAP7_75t_L g618 ( 
.A(n_528),
.Y(n_618)
);

INVx1_ASAP7_75t_L g619 ( 
.A(n_562),
.Y(n_619)
);

INVx2_ASAP7_75t_SL g620 ( 
.A(n_527),
.Y(n_620)
);

NOR2xp33_ASAP7_75t_L g621 ( 
.A(n_601),
.B(n_488),
.Y(n_621)
);

OR2x6_ASAP7_75t_L g622 ( 
.A(n_527),
.B(n_406),
.Y(n_622)
);

INVx2_ASAP7_75t_L g623 ( 
.A(n_528),
.Y(n_623)
);

INVx2_ASAP7_75t_SL g624 ( 
.A(n_545),
.Y(n_624)
);

NAND2xp5_ASAP7_75t_SL g625 ( 
.A(n_553),
.B(n_516),
.Y(n_625)
);

INVx5_ASAP7_75t_L g626 ( 
.A(n_552),
.Y(n_626)
);

INVx3_ASAP7_75t_L g627 ( 
.A(n_570),
.Y(n_627)
);

INVx1_ASAP7_75t_L g628 ( 
.A(n_579),
.Y(n_628)
);

NAND2xp33_ASAP7_75t_R g629 ( 
.A(n_575),
.B(n_438),
.Y(n_629)
);

BUFx6f_ASAP7_75t_L g630 ( 
.A(n_540),
.Y(n_630)
);

NOR2xp33_ASAP7_75t_L g631 ( 
.A(n_563),
.B(n_493),
.Y(n_631)
);

NAND2xp5_ASAP7_75t_L g632 ( 
.A(n_547),
.B(n_453),
.Y(n_632)
);

INVx1_ASAP7_75t_L g633 ( 
.A(n_525),
.Y(n_633)
);

AOI21x1_ASAP7_75t_L g634 ( 
.A1(n_525),
.A2(n_255),
.B(n_245),
.Y(n_634)
);

INVx2_ASAP7_75t_L g635 ( 
.A(n_535),
.Y(n_635)
);

INVx2_ASAP7_75t_L g636 ( 
.A(n_535),
.Y(n_636)
);

INVx2_ASAP7_75t_L g637 ( 
.A(n_535),
.Y(n_637)
);

INVx2_ASAP7_75t_SL g638 ( 
.A(n_545),
.Y(n_638)
);

INVx2_ASAP7_75t_L g639 ( 
.A(n_561),
.Y(n_639)
);

AOI22xp33_ASAP7_75t_L g640 ( 
.A1(n_551),
.A2(n_449),
.B1(n_419),
.B2(n_420),
.Y(n_640)
);

NAND3xp33_ASAP7_75t_L g641 ( 
.A(n_560),
.B(n_454),
.C(n_453),
.Y(n_641)
);

INVx2_ASAP7_75t_L g642 ( 
.A(n_561),
.Y(n_642)
);

INVx2_ASAP7_75t_L g643 ( 
.A(n_561),
.Y(n_643)
);

INVx2_ASAP7_75t_SL g644 ( 
.A(n_553),
.Y(n_644)
);

NOR2xp33_ASAP7_75t_L g645 ( 
.A(n_536),
.B(n_514),
.Y(n_645)
);

BUFx3_ASAP7_75t_L g646 ( 
.A(n_546),
.Y(n_646)
);

INVx2_ASAP7_75t_L g647 ( 
.A(n_593),
.Y(n_647)
);

INVx1_ASAP7_75t_L g648 ( 
.A(n_529),
.Y(n_648)
);

AND3x2_ASAP7_75t_L g649 ( 
.A(n_575),
.B(n_275),
.C(n_255),
.Y(n_649)
);

INVx2_ASAP7_75t_L g650 ( 
.A(n_593),
.Y(n_650)
);

AND2x4_ASAP7_75t_L g651 ( 
.A(n_564),
.B(n_478),
.Y(n_651)
);

NOR2xp33_ASAP7_75t_L g652 ( 
.A(n_526),
.B(n_519),
.Y(n_652)
);

NAND2xp5_ASAP7_75t_SL g653 ( 
.A(n_558),
.B(n_454),
.Y(n_653)
);

INVx2_ASAP7_75t_L g654 ( 
.A(n_593),
.Y(n_654)
);

INVx5_ASAP7_75t_L g655 ( 
.A(n_552),
.Y(n_655)
);

INVx5_ASAP7_75t_L g656 ( 
.A(n_552),
.Y(n_656)
);

INVx1_ASAP7_75t_L g657 ( 
.A(n_598),
.Y(n_657)
);

NOR2x1p5_ASAP7_75t_L g658 ( 
.A(n_586),
.B(n_458),
.Y(n_658)
);

INVx4_ASAP7_75t_L g659 ( 
.A(n_552),
.Y(n_659)
);

INVx1_ASAP7_75t_L g660 ( 
.A(n_529),
.Y(n_660)
);

OR2x6_ASAP7_75t_L g661 ( 
.A(n_538),
.B(n_414),
.Y(n_661)
);

INVx2_ASAP7_75t_L g662 ( 
.A(n_593),
.Y(n_662)
);

INVx1_ASAP7_75t_L g663 ( 
.A(n_598),
.Y(n_663)
);

BUFx6f_ASAP7_75t_L g664 ( 
.A(n_540),
.Y(n_664)
);

BUFx3_ASAP7_75t_L g665 ( 
.A(n_546),
.Y(n_665)
);

INVx1_ASAP7_75t_L g666 ( 
.A(n_598),
.Y(n_666)
);

INVx1_ASAP7_75t_L g667 ( 
.A(n_583),
.Y(n_667)
);

INVx2_ASAP7_75t_L g668 ( 
.A(n_593),
.Y(n_668)
);

INVx2_ASAP7_75t_L g669 ( 
.A(n_593),
.Y(n_669)
);

INVx1_ASAP7_75t_L g670 ( 
.A(n_530),
.Y(n_670)
);

INVx4_ASAP7_75t_L g671 ( 
.A(n_552),
.Y(n_671)
);

INVx2_ASAP7_75t_L g672 ( 
.A(n_530),
.Y(n_672)
);

NAND2xp5_ASAP7_75t_SL g673 ( 
.A(n_558),
.B(n_458),
.Y(n_673)
);

NAND3xp33_ASAP7_75t_L g674 ( 
.A(n_532),
.B(n_467),
.C(n_465),
.Y(n_674)
);

INVx1_ASAP7_75t_L g675 ( 
.A(n_533),
.Y(n_675)
);

INVx1_ASAP7_75t_L g676 ( 
.A(n_533),
.Y(n_676)
);

NAND2xp5_ASAP7_75t_SL g677 ( 
.A(n_569),
.B(n_465),
.Y(n_677)
);

INVx2_ASAP7_75t_L g678 ( 
.A(n_534),
.Y(n_678)
);

BUFx6f_ASAP7_75t_L g679 ( 
.A(n_540),
.Y(n_679)
);

OAI22xp33_ASAP7_75t_L g680 ( 
.A1(n_543),
.A2(n_358),
.B1(n_359),
.B2(n_352),
.Y(n_680)
);

INVx2_ASAP7_75t_SL g681 ( 
.A(n_549),
.Y(n_681)
);

INVxp67_ASAP7_75t_SL g682 ( 
.A(n_570),
.Y(n_682)
);

INVx2_ASAP7_75t_L g683 ( 
.A(n_534),
.Y(n_683)
);

NAND2xp5_ASAP7_75t_SL g684 ( 
.A(n_590),
.B(n_467),
.Y(n_684)
);

INVx2_ASAP7_75t_L g685 ( 
.A(n_537),
.Y(n_685)
);

INVx2_ASAP7_75t_L g686 ( 
.A(n_537),
.Y(n_686)
);

INVx3_ASAP7_75t_L g687 ( 
.A(n_570),
.Y(n_687)
);

AND3x2_ASAP7_75t_L g688 ( 
.A(n_539),
.B(n_356),
.C(n_275),
.Y(n_688)
);

CKINVDCx5p33_ASAP7_75t_R g689 ( 
.A(n_596),
.Y(n_689)
);

INVx1_ASAP7_75t_L g690 ( 
.A(n_544),
.Y(n_690)
);

OR2x6_ASAP7_75t_L g691 ( 
.A(n_571),
.B(n_573),
.Y(n_691)
);

INVx1_ASAP7_75t_SL g692 ( 
.A(n_572),
.Y(n_692)
);

BUFx3_ASAP7_75t_L g693 ( 
.A(n_555),
.Y(n_693)
);

OAI22xp33_ASAP7_75t_L g694 ( 
.A1(n_576),
.A2(n_370),
.B1(n_365),
.B2(n_368),
.Y(n_694)
);

BUFx6f_ASAP7_75t_L g695 ( 
.A(n_540),
.Y(n_695)
);

INVx2_ASAP7_75t_L g696 ( 
.A(n_544),
.Y(n_696)
);

NAND2xp33_ASAP7_75t_L g697 ( 
.A(n_552),
.B(n_313),
.Y(n_697)
);

INVx1_ASAP7_75t_L g698 ( 
.A(n_548),
.Y(n_698)
);

INVx1_ASAP7_75t_L g699 ( 
.A(n_548),
.Y(n_699)
);

INVx1_ASAP7_75t_L g700 ( 
.A(n_554),
.Y(n_700)
);

OAI22xp5_ASAP7_75t_L g701 ( 
.A1(n_583),
.A2(n_476),
.B1(n_497),
.B2(n_477),
.Y(n_701)
);

INVx2_ASAP7_75t_L g702 ( 
.A(n_554),
.Y(n_702)
);

INVx3_ASAP7_75t_L g703 ( 
.A(n_570),
.Y(n_703)
);

INVx2_ASAP7_75t_L g704 ( 
.A(n_557),
.Y(n_704)
);

INVx5_ASAP7_75t_L g705 ( 
.A(n_552),
.Y(n_705)
);

INVx2_ASAP7_75t_L g706 ( 
.A(n_557),
.Y(n_706)
);

INVxp33_ASAP7_75t_L g707 ( 
.A(n_572),
.Y(n_707)
);

AOI22xp5_ASAP7_75t_L g708 ( 
.A1(n_564),
.A2(n_523),
.B1(n_476),
.B2(n_477),
.Y(n_708)
);

NOR3xp33_ASAP7_75t_L g709 ( 
.A(n_600),
.B(n_487),
.C(n_457),
.Y(n_709)
);

INVx1_ASAP7_75t_L g710 ( 
.A(n_585),
.Y(n_710)
);

INVx2_ASAP7_75t_L g711 ( 
.A(n_559),
.Y(n_711)
);

INVxp33_ASAP7_75t_L g712 ( 
.A(n_584),
.Y(n_712)
);

AND2x2_ASAP7_75t_SL g713 ( 
.A(n_555),
.B(n_356),
.Y(n_713)
);

NOR3xp33_ASAP7_75t_L g714 ( 
.A(n_590),
.B(n_517),
.C(n_494),
.Y(n_714)
);

INVx2_ASAP7_75t_L g715 ( 
.A(n_559),
.Y(n_715)
);

BUFx2_ASAP7_75t_L g716 ( 
.A(n_541),
.Y(n_716)
);

INVx1_ASAP7_75t_L g717 ( 
.A(n_568),
.Y(n_717)
);

INVx1_ASAP7_75t_L g718 ( 
.A(n_568),
.Y(n_718)
);

INVx1_ASAP7_75t_L g719 ( 
.A(n_577),
.Y(n_719)
);

INVx5_ASAP7_75t_L g720 ( 
.A(n_552),
.Y(n_720)
);

NOR2xp33_ASAP7_75t_L g721 ( 
.A(n_585),
.B(n_497),
.Y(n_721)
);

BUFx3_ASAP7_75t_L g722 ( 
.A(n_555),
.Y(n_722)
);

BUFx6f_ASAP7_75t_SL g723 ( 
.A(n_555),
.Y(n_723)
);

AND2x2_ASAP7_75t_L g724 ( 
.A(n_584),
.B(n_509),
.Y(n_724)
);

NAND2xp5_ASAP7_75t_SL g725 ( 
.A(n_591),
.B(n_504),
.Y(n_725)
);

CKINVDCx20_ASAP7_75t_R g726 ( 
.A(n_578),
.Y(n_726)
);

INVx1_ASAP7_75t_L g727 ( 
.A(n_577),
.Y(n_727)
);

NAND2xp5_ASAP7_75t_L g728 ( 
.A(n_574),
.B(n_580),
.Y(n_728)
);

NOR2xp33_ASAP7_75t_L g729 ( 
.A(n_587),
.B(n_504),
.Y(n_729)
);

INVx1_ASAP7_75t_L g730 ( 
.A(n_567),
.Y(n_730)
);

AOI22xp33_ASAP7_75t_SL g731 ( 
.A1(n_541),
.A2(n_432),
.B1(n_437),
.B2(n_428),
.Y(n_731)
);

NOR2xp33_ASAP7_75t_L g732 ( 
.A(n_587),
.B(n_505),
.Y(n_732)
);

OAI22xp33_ASAP7_75t_L g733 ( 
.A1(n_576),
.A2(n_371),
.B1(n_466),
.B2(n_379),
.Y(n_733)
);

INVx2_ASAP7_75t_L g734 ( 
.A(n_574),
.Y(n_734)
);

INVx1_ASAP7_75t_L g735 ( 
.A(n_567),
.Y(n_735)
);

AND2x2_ASAP7_75t_L g736 ( 
.A(n_589),
.B(n_510),
.Y(n_736)
);

BUFx3_ASAP7_75t_L g737 ( 
.A(n_567),
.Y(n_737)
);

NAND2xp5_ASAP7_75t_SL g738 ( 
.A(n_591),
.B(n_505),
.Y(n_738)
);

NOR2xp33_ASAP7_75t_L g739 ( 
.A(n_594),
.B(n_511),
.Y(n_739)
);

INVx1_ASAP7_75t_L g740 ( 
.A(n_567),
.Y(n_740)
);

INVx2_ASAP7_75t_L g741 ( 
.A(n_574),
.Y(n_741)
);

INVx2_ASAP7_75t_L g742 ( 
.A(n_574),
.Y(n_742)
);

CKINVDCx6p67_ASAP7_75t_R g743 ( 
.A(n_595),
.Y(n_743)
);

INVxp67_ASAP7_75t_SL g744 ( 
.A(n_540),
.Y(n_744)
);

INVx2_ASAP7_75t_L g745 ( 
.A(n_580),
.Y(n_745)
);

INVx2_ASAP7_75t_SL g746 ( 
.A(n_589),
.Y(n_746)
);

INVx2_ASAP7_75t_L g747 ( 
.A(n_580),
.Y(n_747)
);

NAND2xp5_ASAP7_75t_SL g748 ( 
.A(n_541),
.B(n_511),
.Y(n_748)
);

INVx2_ASAP7_75t_L g749 ( 
.A(n_580),
.Y(n_749)
);

NAND2xp5_ASAP7_75t_L g750 ( 
.A(n_542),
.B(n_515),
.Y(n_750)
);

NOR2xp33_ASAP7_75t_L g751 ( 
.A(n_594),
.B(n_515),
.Y(n_751)
);

INVx2_ASAP7_75t_L g752 ( 
.A(n_542),
.Y(n_752)
);

INVx1_ASAP7_75t_L g753 ( 
.A(n_604),
.Y(n_753)
);

INVx2_ASAP7_75t_SL g754 ( 
.A(n_597),
.Y(n_754)
);

AND2x2_ASAP7_75t_L g755 ( 
.A(n_597),
.B(n_604),
.Y(n_755)
);

NAND2xp5_ASAP7_75t_SL g756 ( 
.A(n_541),
.B(n_212),
.Y(n_756)
);

CKINVDCx20_ASAP7_75t_R g757 ( 
.A(n_556),
.Y(n_757)
);

INVx2_ASAP7_75t_L g758 ( 
.A(n_542),
.Y(n_758)
);

INVx3_ASAP7_75t_L g759 ( 
.A(n_542),
.Y(n_759)
);

NAND2xp5_ASAP7_75t_SL g760 ( 
.A(n_556),
.B(n_212),
.Y(n_760)
);

INVx3_ASAP7_75t_L g761 ( 
.A(n_542),
.Y(n_761)
);

AOI22xp5_ASAP7_75t_L g762 ( 
.A1(n_556),
.A2(n_522),
.B1(n_442),
.B2(n_441),
.Y(n_762)
);

OAI22xp33_ASAP7_75t_L g763 ( 
.A1(n_644),
.A2(n_398),
.B1(n_411),
.B2(n_410),
.Y(n_763)
);

AND2x2_ASAP7_75t_L g764 ( 
.A(n_624),
.B(n_431),
.Y(n_764)
);

INVxp67_ASAP7_75t_L g765 ( 
.A(n_632),
.Y(n_765)
);

BUFx3_ASAP7_75t_L g766 ( 
.A(n_726),
.Y(n_766)
);

NAND2xp5_ASAP7_75t_SL g767 ( 
.A(n_644),
.B(n_556),
.Y(n_767)
);

INVx1_ASAP7_75t_L g768 ( 
.A(n_693),
.Y(n_768)
);

INVx1_ASAP7_75t_L g769 ( 
.A(n_693),
.Y(n_769)
);

INVx2_ASAP7_75t_L g770 ( 
.A(n_627),
.Y(n_770)
);

INVx2_ASAP7_75t_L g771 ( 
.A(n_627),
.Y(n_771)
);

NAND2xp5_ASAP7_75t_L g772 ( 
.A(n_681),
.B(n_603),
.Y(n_772)
);

NOR2xp33_ASAP7_75t_L g773 ( 
.A(n_681),
.B(n_247),
.Y(n_773)
);

NAND2xp5_ASAP7_75t_L g774 ( 
.A(n_610),
.B(n_603),
.Y(n_774)
);

INVx2_ASAP7_75t_L g775 ( 
.A(n_627),
.Y(n_775)
);

NAND2xp5_ASAP7_75t_L g776 ( 
.A(n_610),
.B(n_614),
.Y(n_776)
);

INVx1_ASAP7_75t_L g777 ( 
.A(n_722),
.Y(n_777)
);

NAND3xp33_ASAP7_75t_L g778 ( 
.A(n_612),
.B(n_223),
.C(n_218),
.Y(n_778)
);

INVx2_ASAP7_75t_L g779 ( 
.A(n_687),
.Y(n_779)
);

OAI22xp5_ASAP7_75t_L g780 ( 
.A1(n_713),
.A2(n_624),
.B1(n_638),
.B2(n_746),
.Y(n_780)
);

NOR2xp33_ASAP7_75t_L g781 ( 
.A(n_712),
.B(n_721),
.Y(n_781)
);

BUFx2_ASAP7_75t_L g782 ( 
.A(n_726),
.Y(n_782)
);

NAND2xp5_ASAP7_75t_SL g783 ( 
.A(n_638),
.B(n_218),
.Y(n_783)
);

OR2x6_ASAP7_75t_L g784 ( 
.A(n_716),
.B(n_480),
.Y(n_784)
);

NOR2xp33_ASAP7_75t_L g785 ( 
.A(n_729),
.B(n_295),
.Y(n_785)
);

AOI22xp5_ASAP7_75t_L g786 ( 
.A1(n_652),
.A2(n_440),
.B1(n_323),
.B2(n_331),
.Y(n_786)
);

NAND2xp5_ASAP7_75t_L g787 ( 
.A(n_610),
.B(n_603),
.Y(n_787)
);

AOI22xp5_ASAP7_75t_L g788 ( 
.A1(n_713),
.A2(n_377),
.B1(n_300),
.B2(n_302),
.Y(n_788)
);

NAND2xp5_ASAP7_75t_L g789 ( 
.A(n_614),
.B(n_617),
.Y(n_789)
);

NAND2xp5_ASAP7_75t_L g790 ( 
.A(n_614),
.B(n_603),
.Y(n_790)
);

INVx2_ASAP7_75t_L g791 ( 
.A(n_687),
.Y(n_791)
);

AOI22xp33_ASAP7_75t_L g792 ( 
.A1(n_611),
.A2(n_313),
.B1(n_324),
.B2(n_360),
.Y(n_792)
);

BUFx3_ASAP7_75t_L g793 ( 
.A(n_613),
.Y(n_793)
);

NAND2xp5_ASAP7_75t_L g794 ( 
.A(n_617),
.B(n_605),
.Y(n_794)
);

NOR2xp33_ASAP7_75t_R g795 ( 
.A(n_689),
.B(n_531),
.Y(n_795)
);

AOI22xp5_ASAP7_75t_L g796 ( 
.A1(n_746),
.A2(n_320),
.B1(n_305),
.B2(n_297),
.Y(n_796)
);

NAND2xp5_ASAP7_75t_SL g797 ( 
.A(n_754),
.B(n_223),
.Y(n_797)
);

CKINVDCx20_ASAP7_75t_R g798 ( 
.A(n_743),
.Y(n_798)
);

NOR2xp67_ASAP7_75t_SL g799 ( 
.A(n_626),
.B(n_313),
.Y(n_799)
);

BUFx6f_ASAP7_75t_L g800 ( 
.A(n_722),
.Y(n_800)
);

INVx1_ASAP7_75t_L g801 ( 
.A(n_737),
.Y(n_801)
);

NAND2xp5_ASAP7_75t_L g802 ( 
.A(n_617),
.B(n_605),
.Y(n_802)
);

NAND2xp5_ASAP7_75t_L g803 ( 
.A(n_628),
.B(n_605),
.Y(n_803)
);

OR2x2_ASAP7_75t_L g804 ( 
.A(n_692),
.B(n_484),
.Y(n_804)
);

INVx2_ASAP7_75t_L g805 ( 
.A(n_687),
.Y(n_805)
);

NAND2xp5_ASAP7_75t_L g806 ( 
.A(n_628),
.B(n_619),
.Y(n_806)
);

INVx1_ASAP7_75t_L g807 ( 
.A(n_737),
.Y(n_807)
);

INVxp67_ASAP7_75t_L g808 ( 
.A(n_732),
.Y(n_808)
);

NAND2xp5_ASAP7_75t_L g809 ( 
.A(n_619),
.B(n_605),
.Y(n_809)
);

INVx2_ASAP7_75t_L g810 ( 
.A(n_703),
.Y(n_810)
);

NOR3xp33_ASAP7_75t_L g811 ( 
.A(n_653),
.B(n_243),
.C(n_238),
.Y(n_811)
);

NAND2xp5_ASAP7_75t_SL g812 ( 
.A(n_754),
.B(n_739),
.Y(n_812)
);

AOI22xp33_ASAP7_75t_L g813 ( 
.A1(n_611),
.A2(n_324),
.B1(n_360),
.B2(n_366),
.Y(n_813)
);

INVx2_ASAP7_75t_L g814 ( 
.A(n_703),
.Y(n_814)
);

AO221x1_ASAP7_75t_L g815 ( 
.A1(n_680),
.A2(n_324),
.B1(n_248),
.B2(n_380),
.C(n_253),
.Y(n_815)
);

NAND2xp5_ASAP7_75t_L g816 ( 
.A(n_682),
.B(n_542),
.Y(n_816)
);

NAND2xp5_ASAP7_75t_L g817 ( 
.A(n_667),
.B(n_550),
.Y(n_817)
);

NAND2xp5_ASAP7_75t_L g818 ( 
.A(n_710),
.B(n_550),
.Y(n_818)
);

NAND2xp5_ASAP7_75t_L g819 ( 
.A(n_755),
.B(n_550),
.Y(n_819)
);

INVx1_ASAP7_75t_SL g820 ( 
.A(n_689),
.Y(n_820)
);

NAND2xp5_ASAP7_75t_SL g821 ( 
.A(n_751),
.B(n_224),
.Y(n_821)
);

NAND2xp33_ASAP7_75t_L g822 ( 
.A(n_750),
.B(n_360),
.Y(n_822)
);

NAND2xp33_ASAP7_75t_L g823 ( 
.A(n_620),
.B(n_657),
.Y(n_823)
);

NAND2xp5_ASAP7_75t_L g824 ( 
.A(n_755),
.B(n_730),
.Y(n_824)
);

NAND2xp5_ASAP7_75t_L g825 ( 
.A(n_735),
.B(n_550),
.Y(n_825)
);

NAND2xp5_ASAP7_75t_SL g826 ( 
.A(n_708),
.B(n_224),
.Y(n_826)
);

NAND2xp5_ASAP7_75t_L g827 ( 
.A(n_735),
.B(n_740),
.Y(n_827)
);

NAND2xp5_ASAP7_75t_SL g828 ( 
.A(n_641),
.B(n_225),
.Y(n_828)
);

NAND2xp5_ASAP7_75t_SL g829 ( 
.A(n_674),
.B(n_225),
.Y(n_829)
);

NAND2xp5_ASAP7_75t_SL g830 ( 
.A(n_631),
.B(n_646),
.Y(n_830)
);

NOR2xp33_ASAP7_75t_L g831 ( 
.A(n_621),
.B(n_226),
.Y(n_831)
);

NAND2xp5_ASAP7_75t_L g832 ( 
.A(n_753),
.B(n_550),
.Y(n_832)
);

NAND2xp5_ASAP7_75t_L g833 ( 
.A(n_753),
.B(n_550),
.Y(n_833)
);

NAND2xp5_ASAP7_75t_L g834 ( 
.A(n_663),
.B(n_581),
.Y(n_834)
);

OAI22xp33_ASAP7_75t_L g835 ( 
.A1(n_661),
.A2(n_398),
.B1(n_402),
.B2(n_410),
.Y(n_835)
);

INVx8_ASAP7_75t_L g836 ( 
.A(n_691),
.Y(n_836)
);

NOR2xp33_ASAP7_75t_L g837 ( 
.A(n_673),
.B(n_226),
.Y(n_837)
);

NOR2xp33_ASAP7_75t_L g838 ( 
.A(n_701),
.B(n_625),
.Y(n_838)
);

OR2x6_ASAP7_75t_L g839 ( 
.A(n_716),
.B(n_485),
.Y(n_839)
);

INVx1_ASAP7_75t_L g840 ( 
.A(n_666),
.Y(n_840)
);

OAI22xp33_ASAP7_75t_L g841 ( 
.A1(n_661),
.A2(n_402),
.B1(n_411),
.B2(n_265),
.Y(n_841)
);

NAND2xp5_ASAP7_75t_L g842 ( 
.A(n_620),
.B(n_581),
.Y(n_842)
);

A2O1A1Ixp33_ASAP7_75t_L g843 ( 
.A1(n_633),
.A2(n_660),
.B(n_670),
.C(n_648),
.Y(n_843)
);

AND2x6_ASAP7_75t_L g844 ( 
.A(n_734),
.B(n_324),
.Y(n_844)
);

O2A1O1Ixp5_ASAP7_75t_L g845 ( 
.A1(n_633),
.A2(n_372),
.B(n_364),
.C(n_262),
.Y(n_845)
);

INVx8_ASAP7_75t_L g846 ( 
.A(n_691),
.Y(n_846)
);

INVx2_ASAP7_75t_L g847 ( 
.A(n_703),
.Y(n_847)
);

INVx2_ASAP7_75t_L g848 ( 
.A(n_615),
.Y(n_848)
);

NAND2xp5_ASAP7_75t_L g849 ( 
.A(n_648),
.B(n_581),
.Y(n_849)
);

INVx2_ASAP7_75t_SL g850 ( 
.A(n_613),
.Y(n_850)
);

NAND2xp5_ASAP7_75t_L g851 ( 
.A(n_660),
.B(n_581),
.Y(n_851)
);

INVx2_ASAP7_75t_L g852 ( 
.A(n_615),
.Y(n_852)
);

AOI22xp5_ASAP7_75t_L g853 ( 
.A1(n_723),
.A2(n_287),
.B1(n_284),
.B2(n_282),
.Y(n_853)
);

NAND2xp5_ASAP7_75t_SL g854 ( 
.A(n_646),
.B(n_227),
.Y(n_854)
);

INVx2_ASAP7_75t_L g855 ( 
.A(n_618),
.Y(n_855)
);

NAND2xp5_ASAP7_75t_L g856 ( 
.A(n_670),
.B(n_581),
.Y(n_856)
);

BUFx6f_ASAP7_75t_L g857 ( 
.A(n_665),
.Y(n_857)
);

INVx2_ASAP7_75t_L g858 ( 
.A(n_618),
.Y(n_858)
);

AOI22xp5_ASAP7_75t_L g859 ( 
.A1(n_723),
.A2(n_292),
.B1(n_303),
.B2(n_311),
.Y(n_859)
);

NAND2xp5_ASAP7_75t_L g860 ( 
.A(n_675),
.B(n_676),
.Y(n_860)
);

NAND2xp5_ASAP7_75t_L g861 ( 
.A(n_675),
.B(n_581),
.Y(n_861)
);

NOR2xp33_ASAP7_75t_L g862 ( 
.A(n_665),
.B(n_227),
.Y(n_862)
);

INVx2_ASAP7_75t_L g863 ( 
.A(n_623),
.Y(n_863)
);

INVx2_ASAP7_75t_L g864 ( 
.A(n_623),
.Y(n_864)
);

INVx1_ASAP7_75t_L g865 ( 
.A(n_724),
.Y(n_865)
);

NAND2xp5_ASAP7_75t_L g866 ( 
.A(n_676),
.B(n_266),
.Y(n_866)
);

INVx2_ASAP7_75t_L g867 ( 
.A(n_635),
.Y(n_867)
);

NAND2xp5_ASAP7_75t_L g868 ( 
.A(n_690),
.B(n_698),
.Y(n_868)
);

NAND2xp5_ASAP7_75t_SL g869 ( 
.A(n_651),
.B(n_228),
.Y(n_869)
);

NAND2xp5_ASAP7_75t_SL g870 ( 
.A(n_651),
.B(n_228),
.Y(n_870)
);

AOI221xp5_ASAP7_75t_L g871 ( 
.A1(n_733),
.A2(n_489),
.B1(n_498),
.B2(n_491),
.C(n_490),
.Y(n_871)
);

NOR2xp33_ASAP7_75t_L g872 ( 
.A(n_661),
.B(n_229),
.Y(n_872)
);

NAND2xp5_ASAP7_75t_SL g873 ( 
.A(n_651),
.B(n_229),
.Y(n_873)
);

NAND2xp5_ASAP7_75t_SL g874 ( 
.A(n_613),
.B(n_230),
.Y(n_874)
);

INVx1_ASAP7_75t_L g875 ( 
.A(n_736),
.Y(n_875)
);

NAND2xp5_ASAP7_75t_SL g876 ( 
.A(n_677),
.B(n_230),
.Y(n_876)
);

INVx2_ASAP7_75t_L g877 ( 
.A(n_635),
.Y(n_877)
);

AOI22xp33_ASAP7_75t_L g878 ( 
.A1(n_690),
.A2(n_324),
.B1(n_360),
.B2(n_417),
.Y(n_878)
);

NAND2xp5_ASAP7_75t_SL g879 ( 
.A(n_694),
.B(n_232),
.Y(n_879)
);

AOI22xp5_ASAP7_75t_L g880 ( 
.A1(n_723),
.A2(n_661),
.B1(n_629),
.B2(n_622),
.Y(n_880)
);

NOR2xp33_ASAP7_75t_R g881 ( 
.A(n_757),
.B(n_280),
.Y(n_881)
);

NAND2xp5_ASAP7_75t_SL g882 ( 
.A(n_645),
.B(n_232),
.Y(n_882)
);

INVx3_ASAP7_75t_L g883 ( 
.A(n_734),
.Y(n_883)
);

INVx2_ASAP7_75t_L g884 ( 
.A(n_636),
.Y(n_884)
);

NAND2xp5_ASAP7_75t_L g885 ( 
.A(n_699),
.B(n_268),
.Y(n_885)
);

INVxp67_ASAP7_75t_L g886 ( 
.A(n_699),
.Y(n_886)
);

NAND2xp5_ASAP7_75t_SL g887 ( 
.A(n_700),
.B(n_234),
.Y(n_887)
);

NAND2xp5_ASAP7_75t_L g888 ( 
.A(n_700),
.B(n_286),
.Y(n_888)
);

INVx2_ASAP7_75t_L g889 ( 
.A(n_636),
.Y(n_889)
);

NAND2xp5_ASAP7_75t_SL g890 ( 
.A(n_717),
.B(n_234),
.Y(n_890)
);

INVx4_ASAP7_75t_L g891 ( 
.A(n_616),
.Y(n_891)
);

INVxp67_ASAP7_75t_L g892 ( 
.A(n_717),
.Y(n_892)
);

NAND2x1p5_ASAP7_75t_L g893 ( 
.A(n_659),
.B(n_298),
.Y(n_893)
);

HB1xp67_ASAP7_75t_L g894 ( 
.A(n_622),
.Y(n_894)
);

OAI22xp5_ASAP7_75t_L g895 ( 
.A1(n_718),
.A2(n_299),
.B1(n_301),
.B2(n_416),
.Y(n_895)
);

INVx1_ASAP7_75t_L g896 ( 
.A(n_718),
.Y(n_896)
);

BUFx5_ASAP7_75t_L g897 ( 
.A(n_719),
.Y(n_897)
);

OR2x2_ASAP7_75t_L g898 ( 
.A(n_707),
.B(n_609),
.Y(n_898)
);

INVx2_ASAP7_75t_L g899 ( 
.A(n_637),
.Y(n_899)
);

NOR2xp33_ASAP7_75t_L g900 ( 
.A(n_684),
.B(n_237),
.Y(n_900)
);

CKINVDCx5p33_ASAP7_75t_R g901 ( 
.A(n_743),
.Y(n_901)
);

NAND2xp5_ASAP7_75t_L g902 ( 
.A(n_719),
.B(n_312),
.Y(n_902)
);

AOI22xp33_ASAP7_75t_L g903 ( 
.A1(n_727),
.A2(n_360),
.B1(n_319),
.B2(n_392),
.Y(n_903)
);

NOR2xp33_ASAP7_75t_L g904 ( 
.A(n_725),
.B(n_237),
.Y(n_904)
);

INVx1_ASAP7_75t_L g905 ( 
.A(n_727),
.Y(n_905)
);

NAND2xp5_ASAP7_75t_L g906 ( 
.A(n_672),
.B(n_322),
.Y(n_906)
);

INVx1_ASAP7_75t_L g907 ( 
.A(n_672),
.Y(n_907)
);

NAND2xp5_ASAP7_75t_L g908 ( 
.A(n_678),
.B(n_333),
.Y(n_908)
);

INVx2_ASAP7_75t_L g909 ( 
.A(n_637),
.Y(n_909)
);

BUFx6f_ASAP7_75t_L g910 ( 
.A(n_616),
.Y(n_910)
);

NAND2x1p5_ASAP7_75t_L g911 ( 
.A(n_659),
.B(n_671),
.Y(n_911)
);

NAND2xp5_ASAP7_75t_SL g912 ( 
.A(n_640),
.B(n_659),
.Y(n_912)
);

NAND2xp5_ASAP7_75t_L g913 ( 
.A(n_678),
.B(n_336),
.Y(n_913)
);

NAND2xp5_ASAP7_75t_L g914 ( 
.A(n_683),
.B(n_344),
.Y(n_914)
);

NAND2xp5_ASAP7_75t_SL g915 ( 
.A(n_671),
.B(n_239),
.Y(n_915)
);

AND2x2_ASAP7_75t_SL g916 ( 
.A(n_697),
.B(n_355),
.Y(n_916)
);

NAND2xp5_ASAP7_75t_L g917 ( 
.A(n_683),
.B(n_361),
.Y(n_917)
);

NAND2xp5_ASAP7_75t_L g918 ( 
.A(n_685),
.B(n_391),
.Y(n_918)
);

AND2x4_ASAP7_75t_L g919 ( 
.A(n_622),
.B(n_606),
.Y(n_919)
);

NOR2xp33_ASAP7_75t_L g920 ( 
.A(n_738),
.B(n_756),
.Y(n_920)
);

NAND2xp5_ASAP7_75t_SL g921 ( 
.A(n_671),
.B(n_239),
.Y(n_921)
);

NAND2xp5_ASAP7_75t_L g922 ( 
.A(n_685),
.B(n_397),
.Y(n_922)
);

NAND2xp5_ASAP7_75t_L g923 ( 
.A(n_686),
.B(n_405),
.Y(n_923)
);

NAND2xp5_ASAP7_75t_L g924 ( 
.A(n_686),
.B(n_696),
.Y(n_924)
);

NAND2xp5_ASAP7_75t_L g925 ( 
.A(n_696),
.B(n_407),
.Y(n_925)
);

NOR2xp33_ASAP7_75t_L g926 ( 
.A(n_760),
.B(n_241),
.Y(n_926)
);

NOR2xp33_ASAP7_75t_L g927 ( 
.A(n_622),
.B(n_241),
.Y(n_927)
);

NAND2xp5_ASAP7_75t_SL g928 ( 
.A(n_709),
.B(n_242),
.Y(n_928)
);

NAND2xp5_ASAP7_75t_L g929 ( 
.A(n_785),
.B(n_702),
.Y(n_929)
);

INVx5_ASAP7_75t_L g930 ( 
.A(n_910),
.Y(n_930)
);

INVx3_ASAP7_75t_L g931 ( 
.A(n_800),
.Y(n_931)
);

INVx3_ASAP7_75t_L g932 ( 
.A(n_800),
.Y(n_932)
);

NAND2xp5_ASAP7_75t_SL g933 ( 
.A(n_897),
.B(n_626),
.Y(n_933)
);

NAND2xp33_ASAP7_75t_SL g934 ( 
.A(n_795),
.B(n_748),
.Y(n_934)
);

NAND2xp5_ASAP7_75t_L g935 ( 
.A(n_785),
.B(n_702),
.Y(n_935)
);

AND2x2_ASAP7_75t_L g936 ( 
.A(n_781),
.B(n_691),
.Y(n_936)
);

NOR2xp33_ASAP7_75t_L g937 ( 
.A(n_808),
.B(n_691),
.Y(n_937)
);

OAI21xp5_ASAP7_75t_L g938 ( 
.A1(n_776),
.A2(n_728),
.B(n_744),
.Y(n_938)
);

AND2x6_ASAP7_75t_SL g939 ( 
.A(n_900),
.B(n_510),
.Y(n_939)
);

AOI22xp33_ASAP7_75t_L g940 ( 
.A1(n_792),
.A2(n_704),
.B1(n_706),
.B2(n_711),
.Y(n_940)
);

BUFx2_ASAP7_75t_L g941 ( 
.A(n_764),
.Y(n_941)
);

AOI21xp5_ASAP7_75t_L g942 ( 
.A1(n_789),
.A2(n_655),
.B(n_626),
.Y(n_942)
);

NAND2xp5_ASAP7_75t_SL g943 ( 
.A(n_897),
.B(n_626),
.Y(n_943)
);

HB1xp67_ASAP7_75t_L g944 ( 
.A(n_898),
.Y(n_944)
);

CKINVDCx6p67_ASAP7_75t_R g945 ( 
.A(n_766),
.Y(n_945)
);

NAND2xp5_ASAP7_75t_L g946 ( 
.A(n_773),
.B(n_704),
.Y(n_946)
);

NAND2xp5_ASAP7_75t_L g947 ( 
.A(n_773),
.B(n_706),
.Y(n_947)
);

INVx2_ASAP7_75t_L g948 ( 
.A(n_883),
.Y(n_948)
);

INVx2_ASAP7_75t_L g949 ( 
.A(n_883),
.Y(n_949)
);

INVx4_ASAP7_75t_L g950 ( 
.A(n_857),
.Y(n_950)
);

INVx5_ASAP7_75t_L g951 ( 
.A(n_910),
.Y(n_951)
);

INVx2_ASAP7_75t_L g952 ( 
.A(n_907),
.Y(n_952)
);

NAND2xp5_ASAP7_75t_SL g953 ( 
.A(n_897),
.B(n_626),
.Y(n_953)
);

NAND2xp5_ASAP7_75t_L g954 ( 
.A(n_886),
.B(n_711),
.Y(n_954)
);

INVx2_ASAP7_75t_SL g955 ( 
.A(n_804),
.Y(n_955)
);

NOR3xp33_ASAP7_75t_SL g956 ( 
.A(n_835),
.B(n_244),
.C(n_242),
.Y(n_956)
);

INVx1_ASAP7_75t_L g957 ( 
.A(n_896),
.Y(n_957)
);

INVx5_ASAP7_75t_L g958 ( 
.A(n_910),
.Y(n_958)
);

AND2x6_ASAP7_75t_SL g959 ( 
.A(n_904),
.B(n_658),
.Y(n_959)
);

INVx1_ASAP7_75t_L g960 ( 
.A(n_905),
.Y(n_960)
);

OR2x2_ASAP7_75t_L g961 ( 
.A(n_765),
.B(n_762),
.Y(n_961)
);

NAND2xp5_ASAP7_75t_SL g962 ( 
.A(n_897),
.B(n_655),
.Y(n_962)
);

INVx1_ASAP7_75t_L g963 ( 
.A(n_924),
.Y(n_963)
);

NAND2xp5_ASAP7_75t_L g964 ( 
.A(n_886),
.B(n_715),
.Y(n_964)
);

HB1xp67_ASAP7_75t_L g965 ( 
.A(n_857),
.Y(n_965)
);

INVx1_ASAP7_75t_L g966 ( 
.A(n_827),
.Y(n_966)
);

INVx2_ASAP7_75t_L g967 ( 
.A(n_848),
.Y(n_967)
);

NAND3xp33_ASAP7_75t_SL g968 ( 
.A(n_786),
.B(n_714),
.C(n_731),
.Y(n_968)
);

NAND2xp5_ASAP7_75t_SL g969 ( 
.A(n_897),
.B(n_655),
.Y(n_969)
);

NAND2xp5_ASAP7_75t_L g970 ( 
.A(n_892),
.B(n_715),
.Y(n_970)
);

INVxp67_ASAP7_75t_L g971 ( 
.A(n_781),
.Y(n_971)
);

BUFx3_ASAP7_75t_L g972 ( 
.A(n_857),
.Y(n_972)
);

NOR2xp33_ASAP7_75t_R g973 ( 
.A(n_901),
.B(n_757),
.Y(n_973)
);

NAND2xp5_ASAP7_75t_L g974 ( 
.A(n_892),
.B(n_741),
.Y(n_974)
);

NAND2xp5_ASAP7_75t_L g975 ( 
.A(n_806),
.B(n_741),
.Y(n_975)
);

NAND2xp5_ASAP7_75t_L g976 ( 
.A(n_808),
.B(n_765),
.Y(n_976)
);

NOR2xp33_ASAP7_75t_L g977 ( 
.A(n_831),
.B(n_649),
.Y(n_977)
);

A2O1A1Ixp33_ASAP7_75t_L g978 ( 
.A1(n_838),
.A2(n_749),
.B(n_747),
.C(n_745),
.Y(n_978)
);

INVx1_ASAP7_75t_L g979 ( 
.A(n_819),
.Y(n_979)
);

NAND2xp5_ASAP7_75t_L g980 ( 
.A(n_824),
.B(n_742),
.Y(n_980)
);

NAND2xp5_ASAP7_75t_L g981 ( 
.A(n_772),
.B(n_742),
.Y(n_981)
);

NAND2xp5_ASAP7_75t_L g982 ( 
.A(n_803),
.B(n_745),
.Y(n_982)
);

HB1xp67_ASAP7_75t_L g983 ( 
.A(n_857),
.Y(n_983)
);

INVx2_ASAP7_75t_L g984 ( 
.A(n_852),
.Y(n_984)
);

INVx2_ASAP7_75t_SL g985 ( 
.A(n_782),
.Y(n_985)
);

NAND2xp5_ASAP7_75t_SL g986 ( 
.A(n_897),
.B(n_655),
.Y(n_986)
);

NAND2xp5_ASAP7_75t_SL g987 ( 
.A(n_800),
.B(n_655),
.Y(n_987)
);

AND2x4_ASAP7_75t_L g988 ( 
.A(n_793),
.B(n_688),
.Y(n_988)
);

NAND2xp5_ASAP7_75t_SL g989 ( 
.A(n_800),
.B(n_656),
.Y(n_989)
);

INVx2_ASAP7_75t_L g990 ( 
.A(n_855),
.Y(n_990)
);

BUFx3_ASAP7_75t_L g991 ( 
.A(n_836),
.Y(n_991)
);

INVxp67_ASAP7_75t_L g992 ( 
.A(n_862),
.Y(n_992)
);

AND2x4_ASAP7_75t_L g993 ( 
.A(n_850),
.B(n_606),
.Y(n_993)
);

AOI22xp5_ASAP7_75t_L g994 ( 
.A1(n_780),
.A2(n_669),
.B1(n_650),
.B2(n_654),
.Y(n_994)
);

INVx2_ASAP7_75t_L g995 ( 
.A(n_858),
.Y(n_995)
);

INVx2_ASAP7_75t_L g996 ( 
.A(n_863),
.Y(n_996)
);

NOR2x2_ASAP7_75t_L g997 ( 
.A(n_784),
.B(n_395),
.Y(n_997)
);

OAI22xp33_ASAP7_75t_L g998 ( 
.A1(n_865),
.A2(n_401),
.B1(n_314),
.B2(n_381),
.Y(n_998)
);

INVx1_ASAP7_75t_L g999 ( 
.A(n_768),
.Y(n_999)
);

INVx2_ASAP7_75t_L g1000 ( 
.A(n_864),
.Y(n_1000)
);

NAND2xp5_ASAP7_75t_SL g1001 ( 
.A(n_911),
.B(n_656),
.Y(n_1001)
);

CKINVDCx5p33_ASAP7_75t_R g1002 ( 
.A(n_881),
.Y(n_1002)
);

INVx4_ASAP7_75t_L g1003 ( 
.A(n_910),
.Y(n_1003)
);

BUFx4f_ASAP7_75t_L g1004 ( 
.A(n_836),
.Y(n_1004)
);

INVx1_ASAP7_75t_L g1005 ( 
.A(n_769),
.Y(n_1005)
);

CKINVDCx5p33_ASAP7_75t_R g1006 ( 
.A(n_820),
.Y(n_1006)
);

BUFx4f_ASAP7_75t_L g1007 ( 
.A(n_836),
.Y(n_1007)
);

AOI21xp5_ASAP7_75t_L g1008 ( 
.A1(n_911),
.A2(n_656),
.B(n_705),
.Y(n_1008)
);

NAND2xp5_ASAP7_75t_SL g1009 ( 
.A(n_838),
.B(n_656),
.Y(n_1009)
);

NOR2xp33_ASAP7_75t_L g1010 ( 
.A(n_830),
.B(n_747),
.Y(n_1010)
);

INVx1_ASAP7_75t_L g1011 ( 
.A(n_777),
.Y(n_1011)
);

INVx4_ASAP7_75t_L g1012 ( 
.A(n_846),
.Y(n_1012)
);

CKINVDCx12_ASAP7_75t_R g1013 ( 
.A(n_784),
.Y(n_1013)
);

INVx1_ASAP7_75t_L g1014 ( 
.A(n_801),
.Y(n_1014)
);

INVx2_ASAP7_75t_L g1015 ( 
.A(n_867),
.Y(n_1015)
);

INVx2_ASAP7_75t_L g1016 ( 
.A(n_877),
.Y(n_1016)
);

AND2x4_ASAP7_75t_L g1017 ( 
.A(n_919),
.B(n_607),
.Y(n_1017)
);

AOI22xp5_ASAP7_75t_L g1018 ( 
.A1(n_912),
.A2(n_669),
.B1(n_650),
.B2(n_654),
.Y(n_1018)
);

INVx1_ASAP7_75t_L g1019 ( 
.A(n_807),
.Y(n_1019)
);

OAI21xp5_ASAP7_75t_L g1020 ( 
.A1(n_843),
.A2(n_749),
.B(n_662),
.Y(n_1020)
);

INVx1_ASAP7_75t_L g1021 ( 
.A(n_840),
.Y(n_1021)
);

OR2x2_ASAP7_75t_L g1022 ( 
.A(n_875),
.B(n_607),
.Y(n_1022)
);

NOR2xp33_ASAP7_75t_R g1023 ( 
.A(n_798),
.B(n_244),
.Y(n_1023)
);

NAND2xp5_ASAP7_75t_L g1024 ( 
.A(n_860),
.B(n_759),
.Y(n_1024)
);

AOI22xp33_ASAP7_75t_L g1025 ( 
.A1(n_792),
.A2(n_360),
.B1(n_395),
.B2(n_642),
.Y(n_1025)
);

INVx1_ASAP7_75t_L g1026 ( 
.A(n_868),
.Y(n_1026)
);

NAND2xp5_ASAP7_75t_L g1027 ( 
.A(n_862),
.B(n_759),
.Y(n_1027)
);

AND2x4_ASAP7_75t_L g1028 ( 
.A(n_919),
.B(n_609),
.Y(n_1028)
);

NAND2xp5_ASAP7_75t_L g1029 ( 
.A(n_812),
.B(n_759),
.Y(n_1029)
);

BUFx3_ASAP7_75t_L g1030 ( 
.A(n_846),
.Y(n_1030)
);

INVx1_ASAP7_75t_L g1031 ( 
.A(n_770),
.Y(n_1031)
);

NAND2xp5_ASAP7_75t_L g1032 ( 
.A(n_866),
.B(n_761),
.Y(n_1032)
);

INVx1_ASAP7_75t_L g1033 ( 
.A(n_771),
.Y(n_1033)
);

AOI22xp33_ASAP7_75t_L g1034 ( 
.A1(n_813),
.A2(n_643),
.B1(n_642),
.B2(n_639),
.Y(n_1034)
);

INVx2_ASAP7_75t_SL g1035 ( 
.A(n_846),
.Y(n_1035)
);

AOI22xp5_ASAP7_75t_L g1036 ( 
.A1(n_920),
.A2(n_647),
.B1(n_668),
.B2(n_662),
.Y(n_1036)
);

INVx2_ASAP7_75t_L g1037 ( 
.A(n_884),
.Y(n_1037)
);

AOI21xp5_ASAP7_75t_L g1038 ( 
.A1(n_774),
.A2(n_656),
.B(n_705),
.Y(n_1038)
);

BUFx6f_ASAP7_75t_L g1039 ( 
.A(n_891),
.Y(n_1039)
);

INVx1_ASAP7_75t_L g1040 ( 
.A(n_775),
.Y(n_1040)
);

NAND2xp5_ASAP7_75t_L g1041 ( 
.A(n_885),
.B(n_888),
.Y(n_1041)
);

INVx1_ASAP7_75t_SL g1042 ( 
.A(n_783),
.Y(n_1042)
);

INVx1_ASAP7_75t_L g1043 ( 
.A(n_779),
.Y(n_1043)
);

NAND2xp5_ASAP7_75t_L g1044 ( 
.A(n_902),
.B(n_788),
.Y(n_1044)
);

NAND2xp5_ASAP7_75t_L g1045 ( 
.A(n_837),
.B(n_761),
.Y(n_1045)
);

CKINVDCx5p33_ASAP7_75t_R g1046 ( 
.A(n_784),
.Y(n_1046)
);

INVx2_ASAP7_75t_L g1047 ( 
.A(n_889),
.Y(n_1047)
);

AOI21xp5_ASAP7_75t_L g1048 ( 
.A1(n_787),
.A2(n_705),
.B(n_720),
.Y(n_1048)
);

AOI22xp5_ASAP7_75t_L g1049 ( 
.A1(n_837),
.A2(n_647),
.B1(n_668),
.B2(n_761),
.Y(n_1049)
);

INVx3_ASAP7_75t_L g1050 ( 
.A(n_791),
.Y(n_1050)
);

OR2x2_ASAP7_75t_L g1051 ( 
.A(n_797),
.B(n_314),
.Y(n_1051)
);

NAND2xp5_ASAP7_75t_SL g1052 ( 
.A(n_880),
.B(n_705),
.Y(n_1052)
);

HB1xp67_ASAP7_75t_L g1053 ( 
.A(n_894),
.Y(n_1053)
);

CKINVDCx5p33_ASAP7_75t_R g1054 ( 
.A(n_839),
.Y(n_1054)
);

NAND2xp5_ASAP7_75t_L g1055 ( 
.A(n_809),
.B(n_752),
.Y(n_1055)
);

AND2x2_ASAP7_75t_L g1056 ( 
.A(n_872),
.B(n_582),
.Y(n_1056)
);

AOI22xp33_ASAP7_75t_L g1057 ( 
.A1(n_813),
.A2(n_815),
.B1(n_878),
.B2(n_841),
.Y(n_1057)
);

AND3x1_ASAP7_75t_SL g1058 ( 
.A(n_871),
.B(n_1),
.C(n_2),
.Y(n_1058)
);

AND2x2_ASAP7_75t_L g1059 ( 
.A(n_872),
.B(n_582),
.Y(n_1059)
);

NOR2xp67_ASAP7_75t_L g1060 ( 
.A(n_778),
.B(n_752),
.Y(n_1060)
);

INVx2_ASAP7_75t_L g1061 ( 
.A(n_899),
.Y(n_1061)
);

INVx1_ASAP7_75t_L g1062 ( 
.A(n_805),
.Y(n_1062)
);

NAND2xp5_ASAP7_75t_L g1063 ( 
.A(n_821),
.B(n_758),
.Y(n_1063)
);

NAND2xp5_ASAP7_75t_L g1064 ( 
.A(n_810),
.B(n_758),
.Y(n_1064)
);

INVx2_ASAP7_75t_L g1065 ( 
.A(n_909),
.Y(n_1065)
);

NAND2xp5_ASAP7_75t_L g1066 ( 
.A(n_814),
.B(n_847),
.Y(n_1066)
);

INVx2_ASAP7_75t_L g1067 ( 
.A(n_825),
.Y(n_1067)
);

INVx2_ASAP7_75t_L g1068 ( 
.A(n_832),
.Y(n_1068)
);

INVx2_ASAP7_75t_L g1069 ( 
.A(n_833),
.Y(n_1069)
);

NAND2xp5_ASAP7_75t_SL g1070 ( 
.A(n_790),
.B(n_705),
.Y(n_1070)
);

AND2x2_ASAP7_75t_L g1071 ( 
.A(n_882),
.B(n_582),
.Y(n_1071)
);

AOI22xp5_ASAP7_75t_L g1072 ( 
.A1(n_926),
.A2(n_315),
.B1(n_375),
.B2(n_316),
.Y(n_1072)
);

INVx3_ASAP7_75t_L g1073 ( 
.A(n_891),
.Y(n_1073)
);

INVx1_ASAP7_75t_L g1074 ( 
.A(n_849),
.Y(n_1074)
);

NAND2xp5_ASAP7_75t_L g1075 ( 
.A(n_794),
.B(n_643),
.Y(n_1075)
);

INVx3_ASAP7_75t_L g1076 ( 
.A(n_842),
.Y(n_1076)
);

INVx1_ASAP7_75t_L g1077 ( 
.A(n_851),
.Y(n_1077)
);

INVxp67_ASAP7_75t_SL g1078 ( 
.A(n_802),
.Y(n_1078)
);

INVx1_ASAP7_75t_L g1079 ( 
.A(n_856),
.Y(n_1079)
);

NOR3xp33_ASAP7_75t_SL g1080 ( 
.A(n_835),
.B(n_413),
.C(n_412),
.Y(n_1080)
);

NAND2xp5_ASAP7_75t_L g1081 ( 
.A(n_861),
.B(n_816),
.Y(n_1081)
);

NOR2xp33_ASAP7_75t_L g1082 ( 
.A(n_879),
.B(n_381),
.Y(n_1082)
);

INVx1_ASAP7_75t_L g1083 ( 
.A(n_817),
.Y(n_1083)
);

INVx1_ASAP7_75t_SL g1084 ( 
.A(n_854),
.Y(n_1084)
);

OAI21xp5_ASAP7_75t_L g1085 ( 
.A1(n_893),
.A2(n_634),
.B(n_697),
.Y(n_1085)
);

INVx1_ASAP7_75t_L g1086 ( 
.A(n_818),
.Y(n_1086)
);

NAND2xp5_ASAP7_75t_L g1087 ( 
.A(n_811),
.B(n_616),
.Y(n_1087)
);

INVx2_ASAP7_75t_L g1088 ( 
.A(n_834),
.Y(n_1088)
);

INVx1_ASAP7_75t_L g1089 ( 
.A(n_906),
.Y(n_1089)
);

INVx2_ASAP7_75t_L g1090 ( 
.A(n_908),
.Y(n_1090)
);

NOR2xp33_ASAP7_75t_L g1091 ( 
.A(n_841),
.B(n_384),
.Y(n_1091)
);

NAND2xp5_ASAP7_75t_SL g1092 ( 
.A(n_893),
.B(n_720),
.Y(n_1092)
);

BUFx6f_ASAP7_75t_L g1093 ( 
.A(n_916),
.Y(n_1093)
);

NOR3xp33_ASAP7_75t_SL g1094 ( 
.A(n_763),
.B(n_413),
.C(n_412),
.Y(n_1094)
);

INVx2_ASAP7_75t_L g1095 ( 
.A(n_913),
.Y(n_1095)
);

NAND2xp5_ASAP7_75t_L g1096 ( 
.A(n_811),
.B(n_616),
.Y(n_1096)
);

NAND2xp5_ASAP7_75t_SL g1097 ( 
.A(n_796),
.B(n_720),
.Y(n_1097)
);

INVx2_ASAP7_75t_L g1098 ( 
.A(n_914),
.Y(n_1098)
);

AOI22xp33_ASAP7_75t_L g1099 ( 
.A1(n_878),
.A2(n_566),
.B1(n_592),
.B2(n_588),
.Y(n_1099)
);

INVx1_ASAP7_75t_L g1100 ( 
.A(n_917),
.Y(n_1100)
);

INVx5_ASAP7_75t_L g1101 ( 
.A(n_844),
.Y(n_1101)
);

BUFx3_ASAP7_75t_L g1102 ( 
.A(n_839),
.Y(n_1102)
);

INVx2_ASAP7_75t_L g1103 ( 
.A(n_918),
.Y(n_1103)
);

INVx2_ASAP7_75t_L g1104 ( 
.A(n_922),
.Y(n_1104)
);

INVx2_ASAP7_75t_L g1105 ( 
.A(n_923),
.Y(n_1105)
);

AND2x2_ASAP7_75t_L g1106 ( 
.A(n_927),
.B(n_839),
.Y(n_1106)
);

INVx1_ASAP7_75t_L g1107 ( 
.A(n_925),
.Y(n_1107)
);

NAND2xp5_ASAP7_75t_SL g1108 ( 
.A(n_916),
.B(n_720),
.Y(n_1108)
);

BUFx2_ASAP7_75t_L g1109 ( 
.A(n_927),
.Y(n_1109)
);

INVx1_ASAP7_75t_L g1110 ( 
.A(n_823),
.Y(n_1110)
);

INVx1_ASAP7_75t_SL g1111 ( 
.A(n_869),
.Y(n_1111)
);

INVx1_ASAP7_75t_L g1112 ( 
.A(n_887),
.Y(n_1112)
);

AOI22xp33_ASAP7_75t_L g1113 ( 
.A1(n_903),
.A2(n_566),
.B1(n_592),
.B2(n_588),
.Y(n_1113)
);

AND2x2_ASAP7_75t_L g1114 ( 
.A(n_870),
.B(n_592),
.Y(n_1114)
);

INVx1_ASAP7_75t_L g1115 ( 
.A(n_890),
.Y(n_1115)
);

NAND2xp5_ASAP7_75t_L g1116 ( 
.A(n_1026),
.B(n_966),
.Y(n_1116)
);

OAI22xp5_ASAP7_75t_L g1117 ( 
.A1(n_1057),
.A2(n_903),
.B1(n_763),
.B2(n_826),
.Y(n_1117)
);

AOI21xp5_ASAP7_75t_L g1118 ( 
.A1(n_1081),
.A2(n_921),
.B(n_915),
.Y(n_1118)
);

OAI22xp5_ASAP7_75t_L g1119 ( 
.A1(n_1057),
.A2(n_767),
.B1(n_828),
.B2(n_829),
.Y(n_1119)
);

AND2x2_ASAP7_75t_L g1120 ( 
.A(n_971),
.B(n_873),
.Y(n_1120)
);

NOR2xp33_ASAP7_75t_L g1121 ( 
.A(n_992),
.B(n_976),
.Y(n_1121)
);

HB1xp67_ASAP7_75t_L g1122 ( 
.A(n_1053),
.Y(n_1122)
);

O2A1O1Ixp5_ASAP7_75t_L g1123 ( 
.A1(n_929),
.A2(n_876),
.B(n_845),
.C(n_928),
.Y(n_1123)
);

A2O1A1Ixp33_ASAP7_75t_L g1124 ( 
.A1(n_1082),
.A2(n_874),
.B(n_859),
.C(n_853),
.Y(n_1124)
);

NOR3xp33_ASAP7_75t_SL g1125 ( 
.A(n_968),
.B(n_384),
.C(n_386),
.Y(n_1125)
);

CKINVDCx10_ASAP7_75t_R g1126 ( 
.A(n_973),
.Y(n_1126)
);

NAND2x1_ASAP7_75t_L g1127 ( 
.A(n_1039),
.B(n_616),
.Y(n_1127)
);

BUFx2_ASAP7_75t_L g1128 ( 
.A(n_1006),
.Y(n_1128)
);

O2A1O1Ixp33_ASAP7_75t_SL g1129 ( 
.A1(n_1009),
.A2(n_895),
.B(n_822),
.C(n_845),
.Y(n_1129)
);

AOI21xp5_ASAP7_75t_L g1130 ( 
.A1(n_930),
.A2(n_720),
.B(n_630),
.Y(n_1130)
);

BUFx12f_ASAP7_75t_L g1131 ( 
.A(n_1046),
.Y(n_1131)
);

OAI21xp33_ASAP7_75t_L g1132 ( 
.A1(n_1091),
.A2(n_401),
.B(n_400),
.Y(n_1132)
);

BUFx2_ASAP7_75t_L g1133 ( 
.A(n_985),
.Y(n_1133)
);

AOI21xp5_ASAP7_75t_L g1134 ( 
.A1(n_930),
.A2(n_630),
.B(n_695),
.Y(n_1134)
);

INVx1_ASAP7_75t_L g1135 ( 
.A(n_957),
.Y(n_1135)
);

OAI22xp5_ASAP7_75t_L g1136 ( 
.A1(n_1093),
.A2(n_400),
.B1(n_399),
.B2(n_386),
.Y(n_1136)
);

OAI22xp5_ASAP7_75t_L g1137 ( 
.A1(n_1093),
.A2(n_399),
.B1(n_634),
.B2(n_602),
.Y(n_1137)
);

HB1xp67_ASAP7_75t_L g1138 ( 
.A(n_1053),
.Y(n_1138)
);

INVx2_ASAP7_75t_L g1139 ( 
.A(n_967),
.Y(n_1139)
);

NAND2xp5_ASAP7_75t_SL g1140 ( 
.A(n_936),
.B(n_317),
.Y(n_1140)
);

NAND2xp5_ASAP7_75t_L g1141 ( 
.A(n_935),
.B(n_602),
.Y(n_1141)
);

INVx1_ASAP7_75t_L g1142 ( 
.A(n_960),
.Y(n_1142)
);

O2A1O1Ixp33_ASAP7_75t_L g1143 ( 
.A1(n_1091),
.A2(n_602),
.B(n_608),
.C(n_6),
.Y(n_1143)
);

OAI22x1_ASAP7_75t_L g1144 ( 
.A1(n_1109),
.A2(n_937),
.B1(n_1111),
.B2(n_1054),
.Y(n_1144)
);

NOR3xp33_ASAP7_75t_SL g1145 ( 
.A(n_937),
.B(n_318),
.C(n_321),
.Y(n_1145)
);

INVx1_ASAP7_75t_L g1146 ( 
.A(n_952),
.Y(n_1146)
);

NAND2xp5_ASAP7_75t_SL g1147 ( 
.A(n_1084),
.B(n_330),
.Y(n_1147)
);

OAI21xp33_ASAP7_75t_L g1148 ( 
.A1(n_955),
.A2(n_1082),
.B(n_944),
.Y(n_1148)
);

OAI22xp5_ASAP7_75t_L g1149 ( 
.A1(n_1093),
.A2(n_1025),
.B1(n_940),
.B2(n_1099),
.Y(n_1149)
);

INVx1_ASAP7_75t_SL g1150 ( 
.A(n_944),
.Y(n_1150)
);

AOI22xp5_ASAP7_75t_L g1151 ( 
.A1(n_977),
.A2(n_369),
.B1(n_337),
.B2(n_339),
.Y(n_1151)
);

CKINVDCx5p33_ASAP7_75t_R g1152 ( 
.A(n_1002),
.Y(n_1152)
);

INVx2_ASAP7_75t_L g1153 ( 
.A(n_996),
.Y(n_1153)
);

AOI21x1_ASAP7_75t_L g1154 ( 
.A1(n_1009),
.A2(n_799),
.B(n_608),
.Y(n_1154)
);

INVx1_ASAP7_75t_L g1155 ( 
.A(n_952),
.Y(n_1155)
);

NAND2xp5_ASAP7_75t_L g1156 ( 
.A(n_979),
.B(n_608),
.Y(n_1156)
);

AOI22xp5_ASAP7_75t_L g1157 ( 
.A1(n_977),
.A2(n_374),
.B1(n_341),
.B2(n_343),
.Y(n_1157)
);

NAND3xp33_ASAP7_75t_SL g1158 ( 
.A(n_1023),
.B(n_362),
.C(n_353),
.Y(n_1158)
);

INVx4_ASAP7_75t_L g1159 ( 
.A(n_1039),
.Y(n_1159)
);

OAI22xp5_ASAP7_75t_L g1160 ( 
.A1(n_1093),
.A2(n_332),
.B1(n_349),
.B2(n_350),
.Y(n_1160)
);

NAND2xp5_ASAP7_75t_L g1161 ( 
.A(n_963),
.B(n_695),
.Y(n_1161)
);

INVx4_ASAP7_75t_L g1162 ( 
.A(n_1039),
.Y(n_1162)
);

INVx2_ASAP7_75t_L g1163 ( 
.A(n_996),
.Y(n_1163)
);

OAI22xp5_ASAP7_75t_L g1164 ( 
.A1(n_1025),
.A2(n_695),
.B1(n_679),
.B2(n_664),
.Y(n_1164)
);

OR2x2_ASAP7_75t_L g1165 ( 
.A(n_961),
.B(n_941),
.Y(n_1165)
);

NAND2xp5_ASAP7_75t_L g1166 ( 
.A(n_946),
.B(n_679),
.Y(n_1166)
);

OAI22xp5_ASAP7_75t_SL g1167 ( 
.A1(n_1013),
.A2(n_4),
.B1(n_5),
.B2(n_8),
.Y(n_1167)
);

INVxp67_ASAP7_75t_L g1168 ( 
.A(n_1112),
.Y(n_1168)
);

NOR2xp33_ASAP7_75t_L g1169 ( 
.A(n_1042),
.B(n_679),
.Y(n_1169)
);

NAND2xp5_ASAP7_75t_L g1170 ( 
.A(n_947),
.B(n_679),
.Y(n_1170)
);

O2A1O1Ixp33_ASAP7_75t_L g1171 ( 
.A1(n_1044),
.A2(n_4),
.B(n_5),
.C(n_9),
.Y(n_1171)
);

NAND2xp5_ASAP7_75t_L g1172 ( 
.A(n_1056),
.B(n_679),
.Y(n_1172)
);

A2O1A1Ixp33_ASAP7_75t_L g1173 ( 
.A1(n_1115),
.A2(n_664),
.B(n_630),
.C(n_844),
.Y(n_1173)
);

OAI21xp5_ASAP7_75t_L g1174 ( 
.A1(n_978),
.A2(n_844),
.B(n_566),
.Y(n_1174)
);

NAND2xp5_ASAP7_75t_L g1175 ( 
.A(n_1059),
.B(n_664),
.Y(n_1175)
);

AND2x4_ASAP7_75t_L g1176 ( 
.A(n_1012),
.B(n_664),
.Y(n_1176)
);

OAI21xp5_ASAP7_75t_L g1177 ( 
.A1(n_978),
.A2(n_844),
.B(n_566),
.Y(n_1177)
);

NAND2xp5_ASAP7_75t_L g1178 ( 
.A(n_954),
.B(n_664),
.Y(n_1178)
);

CKINVDCx14_ASAP7_75t_R g1179 ( 
.A(n_973),
.Y(n_1179)
);

AOI21xp5_ASAP7_75t_L g1180 ( 
.A1(n_951),
.A2(n_566),
.B(n_844),
.Y(n_1180)
);

NOR2xp33_ASAP7_75t_L g1181 ( 
.A(n_1051),
.B(n_9),
.Y(n_1181)
);

AOI21xp5_ASAP7_75t_L g1182 ( 
.A1(n_951),
.A2(n_566),
.B(n_167),
.Y(n_1182)
);

OAI22xp5_ASAP7_75t_SL g1183 ( 
.A1(n_1102),
.A2(n_10),
.B1(n_12),
.B2(n_13),
.Y(n_1183)
);

BUFx6f_ASAP7_75t_SL g1184 ( 
.A(n_1102),
.Y(n_1184)
);

BUFx8_ASAP7_75t_SL g1185 ( 
.A(n_1004),
.Y(n_1185)
);

OAI21x1_ASAP7_75t_L g1186 ( 
.A1(n_1020),
.A2(n_171),
.B(n_69),
.Y(n_1186)
);

INVx3_ASAP7_75t_L g1187 ( 
.A(n_1039),
.Y(n_1187)
);

NAND2xp5_ASAP7_75t_L g1188 ( 
.A(n_1067),
.B(n_1089),
.Y(n_1188)
);

AOI21xp33_ASAP7_75t_L g1189 ( 
.A1(n_1041),
.A2(n_13),
.B(n_14),
.Y(n_1189)
);

NAND2xp5_ASAP7_75t_SL g1190 ( 
.A(n_1017),
.B(n_209),
.Y(n_1190)
);

INVx3_ASAP7_75t_SL g1191 ( 
.A(n_945),
.Y(n_1191)
);

OAI22x1_ASAP7_75t_L g1192 ( 
.A1(n_1106),
.A2(n_15),
.B1(n_17),
.B2(n_20),
.Y(n_1192)
);

NAND2x1p5_ASAP7_75t_L g1193 ( 
.A(n_950),
.B(n_166),
.Y(n_1193)
);

A2O1A1Ixp33_ASAP7_75t_L g1194 ( 
.A1(n_1100),
.A2(n_17),
.B(n_20),
.C(n_21),
.Y(n_1194)
);

NAND2xp5_ASAP7_75t_L g1195 ( 
.A(n_964),
.B(n_566),
.Y(n_1195)
);

BUFx3_ASAP7_75t_L g1196 ( 
.A(n_991),
.Y(n_1196)
);

BUFx6f_ASAP7_75t_L g1197 ( 
.A(n_972),
.Y(n_1197)
);

NAND2xp5_ASAP7_75t_SL g1198 ( 
.A(n_1017),
.B(n_1028),
.Y(n_1198)
);

INVx1_ASAP7_75t_L g1199 ( 
.A(n_1021),
.Y(n_1199)
);

OAI21xp5_ASAP7_75t_L g1200 ( 
.A1(n_1075),
.A2(n_566),
.B(n_565),
.Y(n_1200)
);

CKINVDCx5p33_ASAP7_75t_R g1201 ( 
.A(n_959),
.Y(n_1201)
);

CKINVDCx20_ASAP7_75t_R g1202 ( 
.A(n_1023),
.Y(n_1202)
);

AOI21xp5_ASAP7_75t_L g1203 ( 
.A1(n_951),
.A2(n_149),
.B(n_206),
.Y(n_1203)
);

INVx1_ASAP7_75t_L g1204 ( 
.A(n_1000),
.Y(n_1204)
);

NAND2xp5_ASAP7_75t_L g1205 ( 
.A(n_970),
.B(n_565),
.Y(n_1205)
);

INVx1_ASAP7_75t_L g1206 ( 
.A(n_1000),
.Y(n_1206)
);

AOI21xp5_ASAP7_75t_L g1207 ( 
.A1(n_951),
.A2(n_126),
.B(n_197),
.Y(n_1207)
);

NAND2xp33_ASAP7_75t_R g1208 ( 
.A(n_956),
.B(n_1080),
.Y(n_1208)
);

NAND2xp5_ASAP7_75t_L g1209 ( 
.A(n_1067),
.B(n_565),
.Y(n_1209)
);

BUFx6f_ASAP7_75t_L g1210 ( 
.A(n_972),
.Y(n_1210)
);

AND2x2_ASAP7_75t_L g1211 ( 
.A(n_1028),
.B(n_21),
.Y(n_1211)
);

OAI22xp5_ASAP7_75t_SL g1212 ( 
.A1(n_988),
.A2(n_24),
.B1(n_25),
.B2(n_26),
.Y(n_1212)
);

A2O1A1Ixp33_ASAP7_75t_L g1213 ( 
.A1(n_1107),
.A2(n_31),
.B(n_32),
.C(n_33),
.Y(n_1213)
);

NAND2xp5_ASAP7_75t_L g1214 ( 
.A(n_1068),
.B(n_565),
.Y(n_1214)
);

NAND3xp33_ASAP7_75t_L g1215 ( 
.A(n_1094),
.B(n_34),
.C(n_35),
.Y(n_1215)
);

INVx6_ASAP7_75t_L g1216 ( 
.A(n_1012),
.Y(n_1216)
);

AOI21xp5_ASAP7_75t_L g1217 ( 
.A1(n_958),
.A2(n_108),
.B(n_193),
.Y(n_1217)
);

AOI21xp5_ASAP7_75t_L g1218 ( 
.A1(n_958),
.A2(n_1001),
.B(n_1078),
.Y(n_1218)
);

INVx3_ASAP7_75t_L g1219 ( 
.A(n_1073),
.Y(n_1219)
);

NAND2xp5_ASAP7_75t_SL g1220 ( 
.A(n_958),
.B(n_950),
.Y(n_1220)
);

AND2x4_ASAP7_75t_L g1221 ( 
.A(n_991),
.B(n_186),
.Y(n_1221)
);

INVx1_ASAP7_75t_L g1222 ( 
.A(n_1015),
.Y(n_1222)
);

NAND2xp5_ASAP7_75t_SL g1223 ( 
.A(n_958),
.B(n_184),
.Y(n_1223)
);

OAI22xp5_ASAP7_75t_L g1224 ( 
.A1(n_940),
.A2(n_1099),
.B1(n_1034),
.B2(n_1113),
.Y(n_1224)
);

NAND2xp33_ASAP7_75t_R g1225 ( 
.A(n_988),
.B(n_105),
.Y(n_1225)
);

NAND2x1p5_ASAP7_75t_L g1226 ( 
.A(n_1073),
.B(n_97),
.Y(n_1226)
);

A2O1A1Ixp33_ASAP7_75t_L g1227 ( 
.A1(n_1010),
.A2(n_35),
.B(n_36),
.C(n_37),
.Y(n_1227)
);

INVx1_ASAP7_75t_L g1228 ( 
.A(n_1015),
.Y(n_1228)
);

NAND3xp33_ASAP7_75t_SL g1229 ( 
.A(n_1072),
.B(n_39),
.C(n_40),
.Y(n_1229)
);

INVx2_ASAP7_75t_L g1230 ( 
.A(n_1016),
.Y(n_1230)
);

INVx2_ASAP7_75t_L g1231 ( 
.A(n_1016),
.Y(n_1231)
);

INVx3_ASAP7_75t_L g1232 ( 
.A(n_1003),
.Y(n_1232)
);

OAI22x1_ASAP7_75t_L g1233 ( 
.A1(n_1035),
.A2(n_41),
.B1(n_42),
.B2(n_46),
.Y(n_1233)
);

OAI21xp33_ASAP7_75t_L g1234 ( 
.A1(n_1022),
.A2(n_41),
.B(n_46),
.Y(n_1234)
);

O2A1O1Ixp5_ASAP7_75t_L g1235 ( 
.A1(n_1108),
.A2(n_565),
.B(n_52),
.C(n_58),
.Y(n_1235)
);

NAND2xp5_ASAP7_75t_L g1236 ( 
.A(n_1068),
.B(n_1069),
.Y(n_1236)
);

AOI21xp5_ASAP7_75t_L g1237 ( 
.A1(n_1001),
.A2(n_50),
.B(n_58),
.Y(n_1237)
);

AOI21xp5_ASAP7_75t_L g1238 ( 
.A1(n_938),
.A2(n_59),
.B(n_60),
.Y(n_1238)
);

O2A1O1Ixp33_ASAP7_75t_L g1239 ( 
.A1(n_998),
.A2(n_59),
.B(n_60),
.C(n_999),
.Y(n_1239)
);

AND2x2_ASAP7_75t_L g1240 ( 
.A(n_993),
.B(n_1114),
.Y(n_1240)
);

INVx1_ASAP7_75t_L g1241 ( 
.A(n_1065),
.Y(n_1241)
);

AOI21xp5_ASAP7_75t_L g1242 ( 
.A1(n_975),
.A2(n_1092),
.B(n_1027),
.Y(n_1242)
);

BUFx6f_ASAP7_75t_L g1243 ( 
.A(n_1030),
.Y(n_1243)
);

NAND2xp5_ASAP7_75t_L g1244 ( 
.A(n_1069),
.B(n_1074),
.Y(n_1244)
);

AOI21xp5_ASAP7_75t_L g1245 ( 
.A1(n_1092),
.A2(n_986),
.B(n_969),
.Y(n_1245)
);

AND2x2_ASAP7_75t_L g1246 ( 
.A(n_1071),
.B(n_1090),
.Y(n_1246)
);

AND2x2_ASAP7_75t_L g1247 ( 
.A(n_1090),
.B(n_1095),
.Y(n_1247)
);

NAND2xp33_ASAP7_75t_SL g1248 ( 
.A(n_965),
.B(n_983),
.Y(n_1248)
);

AOI21xp5_ASAP7_75t_L g1249 ( 
.A1(n_933),
.A2(n_969),
.B(n_986),
.Y(n_1249)
);

NOR2xp33_ASAP7_75t_L g1250 ( 
.A(n_939),
.B(n_998),
.Y(n_1250)
);

HB1xp67_ASAP7_75t_L g1251 ( 
.A(n_983),
.Y(n_1251)
);

NAND2xp5_ASAP7_75t_SL g1252 ( 
.A(n_934),
.B(n_1095),
.Y(n_1252)
);

INVx1_ASAP7_75t_L g1253 ( 
.A(n_1065),
.Y(n_1253)
);

INVx2_ASAP7_75t_L g1254 ( 
.A(n_948),
.Y(n_1254)
);

CKINVDCx5p33_ASAP7_75t_R g1255 ( 
.A(n_1030),
.Y(n_1255)
);

AOI21xp5_ASAP7_75t_L g1256 ( 
.A1(n_933),
.A2(n_943),
.B(n_962),
.Y(n_1256)
);

OAI22xp5_ASAP7_75t_L g1257 ( 
.A1(n_1034),
.A2(n_1113),
.B1(n_1098),
.B2(n_1105),
.Y(n_1257)
);

OAI22xp5_ASAP7_75t_L g1258 ( 
.A1(n_1098),
.A2(n_1105),
.B1(n_1104),
.B2(n_1103),
.Y(n_1258)
);

NOR3xp33_ASAP7_75t_SL g1259 ( 
.A(n_1005),
.B(n_1019),
.C(n_1011),
.Y(n_1259)
);

O2A1O1Ixp5_ASAP7_75t_L g1260 ( 
.A1(n_1108),
.A2(n_1085),
.B(n_1045),
.C(n_1097),
.Y(n_1260)
);

NOR2xp33_ASAP7_75t_SL g1261 ( 
.A(n_1004),
.B(n_1007),
.Y(n_1261)
);

BUFx12f_ASAP7_75t_L g1262 ( 
.A(n_1003),
.Y(n_1262)
);

AND2x2_ASAP7_75t_L g1263 ( 
.A(n_1103),
.B(n_1104),
.Y(n_1263)
);

BUFx3_ASAP7_75t_L g1264 ( 
.A(n_1007),
.Y(n_1264)
);

INVx5_ASAP7_75t_L g1265 ( 
.A(n_931),
.Y(n_1265)
);

AND2x2_ASAP7_75t_L g1266 ( 
.A(n_1014),
.B(n_1086),
.Y(n_1266)
);

INVx3_ASAP7_75t_L g1267 ( 
.A(n_931),
.Y(n_1267)
);

NAND2xp5_ASAP7_75t_L g1268 ( 
.A(n_1077),
.B(n_1079),
.Y(n_1268)
);

A2O1A1Ixp33_ASAP7_75t_L g1269 ( 
.A1(n_1010),
.A2(n_1110),
.B(n_1083),
.C(n_1063),
.Y(n_1269)
);

OAI21x1_ASAP7_75t_L g1270 ( 
.A1(n_1245),
.A2(n_1076),
.B(n_1055),
.Y(n_1270)
);

NOR2xp33_ASAP7_75t_L g1271 ( 
.A(n_1121),
.B(n_1029),
.Y(n_1271)
);

A2O1A1Ixp33_ASAP7_75t_L g1272 ( 
.A1(n_1124),
.A2(n_1060),
.B(n_1096),
.C(n_1087),
.Y(n_1272)
);

NAND2xp5_ASAP7_75t_L g1273 ( 
.A(n_1116),
.B(n_1088),
.Y(n_1273)
);

AOI21xp5_ASAP7_75t_L g1274 ( 
.A1(n_1118),
.A2(n_1032),
.B(n_1024),
.Y(n_1274)
);

OAI21xp5_ASAP7_75t_L g1275 ( 
.A1(n_1260),
.A2(n_1242),
.B(n_1238),
.Y(n_1275)
);

O2A1O1Ixp5_ASAP7_75t_L g1276 ( 
.A1(n_1252),
.A2(n_1052),
.B(n_1097),
.C(n_1070),
.Y(n_1276)
);

O2A1O1Ixp33_ASAP7_75t_SL g1277 ( 
.A1(n_1117),
.A2(n_1052),
.B(n_1070),
.C(n_974),
.Y(n_1277)
);

INVx1_ASAP7_75t_L g1278 ( 
.A(n_1199),
.Y(n_1278)
);

NAND2xp5_ASAP7_75t_L g1279 ( 
.A(n_1247),
.B(n_1088),
.Y(n_1279)
);

INVx4_ASAP7_75t_L g1280 ( 
.A(n_1216),
.Y(n_1280)
);

AND2x2_ASAP7_75t_L g1281 ( 
.A(n_1240),
.B(n_1037),
.Y(n_1281)
);

AOI21xp5_ASAP7_75t_L g1282 ( 
.A1(n_1224),
.A2(n_982),
.B(n_980),
.Y(n_1282)
);

NAND2xp5_ASAP7_75t_L g1283 ( 
.A(n_1263),
.B(n_1116),
.Y(n_1283)
);

OAI21x1_ASAP7_75t_L g1284 ( 
.A1(n_1249),
.A2(n_1076),
.B(n_1018),
.Y(n_1284)
);

INVx3_ASAP7_75t_SL g1285 ( 
.A(n_1191),
.Y(n_1285)
);

OAI21x1_ASAP7_75t_L g1286 ( 
.A1(n_1256),
.A2(n_1064),
.B(n_994),
.Y(n_1286)
);

BUFx6f_ASAP7_75t_L g1287 ( 
.A(n_1243),
.Y(n_1287)
);

AOI21xp5_ASAP7_75t_L g1288 ( 
.A1(n_1224),
.A2(n_953),
.B(n_943),
.Y(n_1288)
);

NAND2xp5_ASAP7_75t_L g1289 ( 
.A(n_1246),
.B(n_932),
.Y(n_1289)
);

INVx3_ASAP7_75t_L g1290 ( 
.A(n_1159),
.Y(n_1290)
);

NAND2x1p5_ASAP7_75t_L g1291 ( 
.A(n_1159),
.B(n_932),
.Y(n_1291)
);

OAI21x1_ASAP7_75t_L g1292 ( 
.A1(n_1154),
.A2(n_981),
.B(n_1066),
.Y(n_1292)
);

INVx6_ASAP7_75t_SL g1293 ( 
.A(n_1221),
.Y(n_1293)
);

BUFx3_ASAP7_75t_L g1294 ( 
.A(n_1133),
.Y(n_1294)
);

NOR2x1_ASAP7_75t_R g1295 ( 
.A(n_1152),
.B(n_997),
.Y(n_1295)
);

AOI21xp5_ASAP7_75t_L g1296 ( 
.A1(n_1149),
.A2(n_953),
.B(n_962),
.Y(n_1296)
);

NAND2x1_ASAP7_75t_L g1297 ( 
.A(n_1162),
.B(n_1050),
.Y(n_1297)
);

NAND2xp5_ASAP7_75t_L g1298 ( 
.A(n_1188),
.B(n_1268),
.Y(n_1298)
);

AO31x2_ASAP7_75t_L g1299 ( 
.A1(n_1137),
.A2(n_949),
.A3(n_948),
.B(n_1031),
.Y(n_1299)
);

NAND2xp5_ASAP7_75t_L g1300 ( 
.A(n_1188),
.B(n_1266),
.Y(n_1300)
);

NAND2xp5_ASAP7_75t_L g1301 ( 
.A(n_1258),
.B(n_995),
.Y(n_1301)
);

NAND2xp5_ASAP7_75t_L g1302 ( 
.A(n_1258),
.B(n_1047),
.Y(n_1302)
);

NAND2xp5_ASAP7_75t_L g1303 ( 
.A(n_1244),
.B(n_990),
.Y(n_1303)
);

NOR2xp67_ASAP7_75t_L g1304 ( 
.A(n_1162),
.B(n_1050),
.Y(n_1304)
);

INVx1_ASAP7_75t_L g1305 ( 
.A(n_1135),
.Y(n_1305)
);

OAI21x1_ASAP7_75t_L g1306 ( 
.A1(n_1218),
.A2(n_1036),
.B(n_1049),
.Y(n_1306)
);

AOI21xp5_ASAP7_75t_L g1307 ( 
.A1(n_1149),
.A2(n_1008),
.B(n_989),
.Y(n_1307)
);

NAND2xp5_ASAP7_75t_L g1308 ( 
.A(n_1120),
.B(n_1061),
.Y(n_1308)
);

OAI21x1_ASAP7_75t_L g1309 ( 
.A1(n_1186),
.A2(n_942),
.B(n_1038),
.Y(n_1309)
);

INVx1_ASAP7_75t_L g1310 ( 
.A(n_1142),
.Y(n_1310)
);

OAI21xp5_ASAP7_75t_L g1311 ( 
.A1(n_1123),
.A2(n_1040),
.B(n_1062),
.Y(n_1311)
);

INVx1_ASAP7_75t_L g1312 ( 
.A(n_1146),
.Y(n_1312)
);

OAI21x1_ASAP7_75t_L g1313 ( 
.A1(n_1174),
.A2(n_1048),
.B(n_949),
.Y(n_1313)
);

OAI21x1_ASAP7_75t_L g1314 ( 
.A1(n_1174),
.A2(n_1033),
.B(n_1043),
.Y(n_1314)
);

NAND2xp5_ASAP7_75t_L g1315 ( 
.A(n_1236),
.B(n_984),
.Y(n_1315)
);

O2A1O1Ixp5_ASAP7_75t_SL g1316 ( 
.A1(n_1189),
.A2(n_1119),
.B(n_1137),
.C(n_1117),
.Y(n_1316)
);

NAND2xp5_ASAP7_75t_L g1317 ( 
.A(n_1168),
.B(n_987),
.Y(n_1317)
);

CKINVDCx5p33_ASAP7_75t_R g1318 ( 
.A(n_1126),
.Y(n_1318)
);

CKINVDCx20_ASAP7_75t_R g1319 ( 
.A(n_1179),
.Y(n_1319)
);

NAND2xp5_ASAP7_75t_L g1320 ( 
.A(n_1181),
.B(n_987),
.Y(n_1320)
);

INVx2_ASAP7_75t_SL g1321 ( 
.A(n_1196),
.Y(n_1321)
);

AOI21xp5_ASAP7_75t_L g1322 ( 
.A1(n_1257),
.A2(n_989),
.B(n_1101),
.Y(n_1322)
);

OAI21x1_ASAP7_75t_L g1323 ( 
.A1(n_1177),
.A2(n_1101),
.B(n_1058),
.Y(n_1323)
);

A2O1A1Ixp33_ASAP7_75t_L g1324 ( 
.A1(n_1119),
.A2(n_1058),
.B(n_1101),
.C(n_1250),
.Y(n_1324)
);

INVx3_ASAP7_75t_L g1325 ( 
.A(n_1187),
.Y(n_1325)
);

AND2x2_ASAP7_75t_L g1326 ( 
.A(n_1165),
.B(n_1101),
.Y(n_1326)
);

OAI21x1_ASAP7_75t_SL g1327 ( 
.A1(n_1237),
.A2(n_1239),
.B(n_1143),
.Y(n_1327)
);

NOR2x1_ASAP7_75t_SL g1328 ( 
.A(n_1257),
.B(n_1265),
.Y(n_1328)
);

AOI21xp5_ASAP7_75t_SL g1329 ( 
.A1(n_1164),
.A2(n_1269),
.B(n_1172),
.Y(n_1329)
);

INVx2_ASAP7_75t_SL g1330 ( 
.A(n_1255),
.Y(n_1330)
);

AOI21xp5_ASAP7_75t_L g1331 ( 
.A1(n_1175),
.A2(n_1141),
.B(n_1170),
.Y(n_1331)
);

AO21x1_ASAP7_75t_L g1332 ( 
.A1(n_1171),
.A2(n_1248),
.B(n_1189),
.Y(n_1332)
);

NAND2xp5_ASAP7_75t_L g1333 ( 
.A(n_1155),
.B(n_1204),
.Y(n_1333)
);

A2O1A1Ixp33_ASAP7_75t_L g1334 ( 
.A1(n_1125),
.A2(n_1148),
.B(n_1132),
.C(n_1259),
.Y(n_1334)
);

AOI221xp5_ASAP7_75t_L g1335 ( 
.A1(n_1229),
.A2(n_1234),
.B1(n_1192),
.B2(n_1144),
.C(n_1215),
.Y(n_1335)
);

NAND2xp5_ASAP7_75t_L g1336 ( 
.A(n_1150),
.B(n_1251),
.Y(n_1336)
);

CKINVDCx5p33_ASAP7_75t_R g1337 ( 
.A(n_1128),
.Y(n_1337)
);

OAI21x1_ASAP7_75t_L g1338 ( 
.A1(n_1134),
.A2(n_1164),
.B(n_1209),
.Y(n_1338)
);

INVxp67_ASAP7_75t_SL g1339 ( 
.A(n_1122),
.Y(n_1339)
);

NAND2xp5_ASAP7_75t_L g1340 ( 
.A(n_1150),
.B(n_1169),
.Y(n_1340)
);

AO21x2_ASAP7_75t_L g1341 ( 
.A1(n_1173),
.A2(n_1166),
.B(n_1129),
.Y(n_1341)
);

OAI21x1_ASAP7_75t_L g1342 ( 
.A1(n_1214),
.A2(n_1178),
.B(n_1200),
.Y(n_1342)
);

NAND2xp5_ASAP7_75t_L g1343 ( 
.A(n_1206),
.B(n_1222),
.Y(n_1343)
);

NAND2xp5_ASAP7_75t_L g1344 ( 
.A(n_1198),
.B(n_1156),
.Y(n_1344)
);

NAND2xp5_ASAP7_75t_L g1345 ( 
.A(n_1140),
.B(n_1230),
.Y(n_1345)
);

AO31x2_ASAP7_75t_L g1346 ( 
.A1(n_1227),
.A2(n_1213),
.A3(n_1194),
.B(n_1205),
.Y(n_1346)
);

NOR2xp33_ASAP7_75t_L g1347 ( 
.A(n_1138),
.B(n_1147),
.Y(n_1347)
);

OR2x6_ASAP7_75t_L g1348 ( 
.A(n_1216),
.B(n_1264),
.Y(n_1348)
);

NAND2x1p5_ASAP7_75t_L g1349 ( 
.A(n_1197),
.B(n_1210),
.Y(n_1349)
);

OAI21x1_ASAP7_75t_L g1350 ( 
.A1(n_1200),
.A2(n_1161),
.B(n_1127),
.Y(n_1350)
);

NAND2xp5_ASAP7_75t_L g1351 ( 
.A(n_1139),
.B(n_1153),
.Y(n_1351)
);

NAND2xp5_ASAP7_75t_L g1352 ( 
.A(n_1163),
.B(n_1231),
.Y(n_1352)
);

A2O1A1Ixp33_ASAP7_75t_L g1353 ( 
.A1(n_1145),
.A2(n_1235),
.B(n_1157),
.C(n_1151),
.Y(n_1353)
);

OAI21x1_ASAP7_75t_L g1354 ( 
.A1(n_1130),
.A2(n_1254),
.B(n_1241),
.Y(n_1354)
);

A2O1A1Ixp33_ASAP7_75t_L g1355 ( 
.A1(n_1190),
.A2(n_1228),
.B(n_1253),
.C(n_1261),
.Y(n_1355)
);

AOI21xp5_ASAP7_75t_L g1356 ( 
.A1(n_1195),
.A2(n_1219),
.B(n_1220),
.Y(n_1356)
);

NOR2xp33_ASAP7_75t_L g1357 ( 
.A(n_1136),
.B(n_1158),
.Y(n_1357)
);

O2A1O1Ixp5_ASAP7_75t_L g1358 ( 
.A1(n_1223),
.A2(n_1160),
.B(n_1136),
.C(n_1207),
.Y(n_1358)
);

NAND2xp5_ASAP7_75t_L g1359 ( 
.A(n_1221),
.B(n_1211),
.Y(n_1359)
);

OAI21xp5_ASAP7_75t_L g1360 ( 
.A1(n_1203),
.A2(n_1217),
.B(n_1182),
.Y(n_1360)
);

OAI22x1_ASAP7_75t_L g1361 ( 
.A1(n_1201),
.A2(n_1226),
.B1(n_1183),
.B2(n_1167),
.Y(n_1361)
);

O2A1O1Ixp5_ASAP7_75t_SL g1362 ( 
.A1(n_1160),
.A2(n_1267),
.B(n_1219),
.C(n_1187),
.Y(n_1362)
);

INVx3_ASAP7_75t_L g1363 ( 
.A(n_1176),
.Y(n_1363)
);

OAI21x1_ASAP7_75t_L g1364 ( 
.A1(n_1180),
.A2(n_1226),
.B(n_1267),
.Y(n_1364)
);

CKINVDCx5p33_ASAP7_75t_R g1365 ( 
.A(n_1185),
.Y(n_1365)
);

NAND2xp5_ASAP7_75t_L g1366 ( 
.A(n_1197),
.B(n_1210),
.Y(n_1366)
);

OA21x2_ASAP7_75t_L g1367 ( 
.A1(n_1176),
.A2(n_1193),
.B(n_1265),
.Y(n_1367)
);

BUFx6f_ASAP7_75t_L g1368 ( 
.A(n_1262),
.Y(n_1368)
);

INVx3_ASAP7_75t_L g1369 ( 
.A(n_1232),
.Y(n_1369)
);

AOI21xp5_ASAP7_75t_L g1370 ( 
.A1(n_1232),
.A2(n_1265),
.B(n_1261),
.Y(n_1370)
);

NOR2xp33_ASAP7_75t_L g1371 ( 
.A(n_1202),
.B(n_1184),
.Y(n_1371)
);

AOI21xp5_ASAP7_75t_L g1372 ( 
.A1(n_1265),
.A2(n_1193),
.B(n_1233),
.Y(n_1372)
);

AOI22xp5_ASAP7_75t_L g1373 ( 
.A1(n_1208),
.A2(n_1225),
.B1(n_1212),
.B2(n_1184),
.Y(n_1373)
);

NAND2xp5_ASAP7_75t_L g1374 ( 
.A(n_1131),
.B(n_971),
.Y(n_1374)
);

AND2x2_ASAP7_75t_L g1375 ( 
.A(n_1240),
.B(n_781),
.Y(n_1375)
);

OR2x2_ASAP7_75t_L g1376 ( 
.A(n_1165),
.B(n_944),
.Y(n_1376)
);

BUFx12f_ASAP7_75t_L g1377 ( 
.A(n_1128),
.Y(n_1377)
);

OAI21x1_ASAP7_75t_L g1378 ( 
.A1(n_1245),
.A2(n_1256),
.B(n_1249),
.Y(n_1378)
);

AOI21xp5_ASAP7_75t_L g1379 ( 
.A1(n_1118),
.A2(n_911),
.B(n_789),
.Y(n_1379)
);

AO31x2_ASAP7_75t_L g1380 ( 
.A1(n_1238),
.A2(n_978),
.A3(n_1137),
.B(n_1119),
.Y(n_1380)
);

NAND2xp5_ASAP7_75t_L g1381 ( 
.A(n_1116),
.B(n_971),
.Y(n_1381)
);

OAI21x1_ASAP7_75t_L g1382 ( 
.A1(n_1245),
.A2(n_1256),
.B(n_1249),
.Y(n_1382)
);

NOR2xp67_ASAP7_75t_L g1383 ( 
.A(n_1159),
.B(n_1162),
.Y(n_1383)
);

NAND2xp5_ASAP7_75t_L g1384 ( 
.A(n_1116),
.B(n_971),
.Y(n_1384)
);

NAND2xp5_ASAP7_75t_L g1385 ( 
.A(n_1116),
.B(n_971),
.Y(n_1385)
);

NAND2xp5_ASAP7_75t_L g1386 ( 
.A(n_1116),
.B(n_971),
.Y(n_1386)
);

NAND2xp5_ASAP7_75t_L g1387 ( 
.A(n_1116),
.B(n_971),
.Y(n_1387)
);

AOI21xp33_ASAP7_75t_L g1388 ( 
.A1(n_1119),
.A2(n_785),
.B(n_831),
.Y(n_1388)
);

NAND2xp5_ASAP7_75t_L g1389 ( 
.A(n_1116),
.B(n_971),
.Y(n_1389)
);

NOR2xp33_ASAP7_75t_L g1390 ( 
.A(n_1121),
.B(n_971),
.Y(n_1390)
);

AND2x4_ASAP7_75t_L g1391 ( 
.A(n_1264),
.B(n_1012),
.Y(n_1391)
);

INVx1_ASAP7_75t_L g1392 ( 
.A(n_1199),
.Y(n_1392)
);

NAND2xp5_ASAP7_75t_L g1393 ( 
.A(n_1116),
.B(n_971),
.Y(n_1393)
);

O2A1O1Ixp5_ASAP7_75t_L g1394 ( 
.A1(n_1238),
.A2(n_831),
.B(n_785),
.C(n_1252),
.Y(n_1394)
);

INVx1_ASAP7_75t_L g1395 ( 
.A(n_1199),
.Y(n_1395)
);

INVxp67_ASAP7_75t_SL g1396 ( 
.A(n_1122),
.Y(n_1396)
);

INVxp67_ASAP7_75t_L g1397 ( 
.A(n_1128),
.Y(n_1397)
);

AOI221xp5_ASAP7_75t_L g1398 ( 
.A1(n_1250),
.A2(n_968),
.B1(n_785),
.B2(n_612),
.C(n_838),
.Y(n_1398)
);

A2O1A1Ixp33_ASAP7_75t_L g1399 ( 
.A1(n_1124),
.A2(n_785),
.B(n_831),
.C(n_838),
.Y(n_1399)
);

BUFx6f_ASAP7_75t_L g1400 ( 
.A(n_1243),
.Y(n_1400)
);

AND3x4_ASAP7_75t_L g1401 ( 
.A(n_1264),
.B(n_766),
.C(n_714),
.Y(n_1401)
);

OAI21x1_ASAP7_75t_SL g1402 ( 
.A1(n_1238),
.A2(n_1237),
.B(n_1239),
.Y(n_1402)
);

AOI21xp5_ASAP7_75t_L g1403 ( 
.A1(n_1118),
.A2(n_911),
.B(n_789),
.Y(n_1403)
);

CKINVDCx11_ASAP7_75t_R g1404 ( 
.A(n_1191),
.Y(n_1404)
);

BUFx6f_ASAP7_75t_L g1405 ( 
.A(n_1243),
.Y(n_1405)
);

NAND2xp5_ASAP7_75t_L g1406 ( 
.A(n_1116),
.B(n_971),
.Y(n_1406)
);

AO32x2_ASAP7_75t_L g1407 ( 
.A1(n_1117),
.A2(n_1119),
.A3(n_1137),
.B1(n_1258),
.B2(n_1257),
.Y(n_1407)
);

NAND2xp5_ASAP7_75t_L g1408 ( 
.A(n_1116),
.B(n_971),
.Y(n_1408)
);

NOR2xp33_ASAP7_75t_R g1409 ( 
.A(n_1179),
.B(n_726),
.Y(n_1409)
);

INVx1_ASAP7_75t_L g1410 ( 
.A(n_1199),
.Y(n_1410)
);

NAND2xp5_ASAP7_75t_L g1411 ( 
.A(n_1116),
.B(n_971),
.Y(n_1411)
);

NAND2xp5_ASAP7_75t_L g1412 ( 
.A(n_1247),
.B(n_1263),
.Y(n_1412)
);

INVx1_ASAP7_75t_SL g1413 ( 
.A(n_1150),
.Y(n_1413)
);

OA21x2_ASAP7_75t_L g1414 ( 
.A1(n_1260),
.A2(n_1242),
.B(n_978),
.Y(n_1414)
);

INVx1_ASAP7_75t_L g1415 ( 
.A(n_1199),
.Y(n_1415)
);

NAND2xp5_ASAP7_75t_L g1416 ( 
.A(n_1116),
.B(n_971),
.Y(n_1416)
);

NAND2xp5_ASAP7_75t_L g1417 ( 
.A(n_1116),
.B(n_971),
.Y(n_1417)
);

CKINVDCx5p33_ASAP7_75t_R g1418 ( 
.A(n_1152),
.Y(n_1418)
);

O2A1O1Ixp33_ASAP7_75t_L g1419 ( 
.A1(n_1181),
.A2(n_785),
.B(n_612),
.C(n_808),
.Y(n_1419)
);

OA21x2_ASAP7_75t_L g1420 ( 
.A1(n_1260),
.A2(n_1242),
.B(n_978),
.Y(n_1420)
);

NAND2x1p5_ASAP7_75t_L g1421 ( 
.A(n_1367),
.B(n_1413),
.Y(n_1421)
);

OAI21xp5_ASAP7_75t_L g1422 ( 
.A1(n_1399),
.A2(n_1388),
.B(n_1316),
.Y(n_1422)
);

OR2x6_ASAP7_75t_L g1423 ( 
.A(n_1372),
.B(n_1370),
.Y(n_1423)
);

AND2x2_ASAP7_75t_L g1424 ( 
.A(n_1375),
.B(n_1281),
.Y(n_1424)
);

OAI21x1_ASAP7_75t_L g1425 ( 
.A1(n_1270),
.A2(n_1313),
.B(n_1338),
.Y(n_1425)
);

OA21x2_ASAP7_75t_L g1426 ( 
.A1(n_1275),
.A2(n_1306),
.B(n_1342),
.Y(n_1426)
);

NAND2xp5_ASAP7_75t_L g1427 ( 
.A(n_1298),
.B(n_1283),
.Y(n_1427)
);

OR2x6_ASAP7_75t_L g1428 ( 
.A(n_1327),
.B(n_1329),
.Y(n_1428)
);

CKINVDCx8_ASAP7_75t_R g1429 ( 
.A(n_1418),
.Y(n_1429)
);

CKINVDCx6p67_ASAP7_75t_R g1430 ( 
.A(n_1285),
.Y(n_1430)
);

AND2x2_ASAP7_75t_L g1431 ( 
.A(n_1390),
.B(n_1271),
.Y(n_1431)
);

BUFx6f_ASAP7_75t_L g1432 ( 
.A(n_1348),
.Y(n_1432)
);

OAI21x1_ASAP7_75t_L g1433 ( 
.A1(n_1284),
.A2(n_1286),
.B(n_1292),
.Y(n_1433)
);

NAND2xp5_ASAP7_75t_L g1434 ( 
.A(n_1283),
.B(n_1273),
.Y(n_1434)
);

NAND2x1p5_ASAP7_75t_L g1435 ( 
.A(n_1367),
.B(n_1413),
.Y(n_1435)
);

O2A1O1Ixp33_ASAP7_75t_SL g1436 ( 
.A1(n_1388),
.A2(n_1324),
.B(n_1353),
.C(n_1398),
.Y(n_1436)
);

OAI21x1_ASAP7_75t_SL g1437 ( 
.A1(n_1402),
.A2(n_1332),
.B(n_1328),
.Y(n_1437)
);

NAND2x1p5_ASAP7_75t_L g1438 ( 
.A(n_1280),
.B(n_1290),
.Y(n_1438)
);

CKINVDCx5p33_ASAP7_75t_R g1439 ( 
.A(n_1404),
.Y(n_1439)
);

OA21x2_ASAP7_75t_L g1440 ( 
.A1(n_1275),
.A2(n_1274),
.B(n_1311),
.Y(n_1440)
);

NAND2xp5_ASAP7_75t_L g1441 ( 
.A(n_1300),
.B(n_1279),
.Y(n_1441)
);

NAND2xp5_ASAP7_75t_L g1442 ( 
.A(n_1279),
.B(n_1412),
.Y(n_1442)
);

OA21x2_ASAP7_75t_L g1443 ( 
.A1(n_1311),
.A2(n_1331),
.B(n_1394),
.Y(n_1443)
);

OAI21x1_ASAP7_75t_L g1444 ( 
.A1(n_1307),
.A2(n_1364),
.B(n_1350),
.Y(n_1444)
);

AO21x2_ASAP7_75t_L g1445 ( 
.A1(n_1360),
.A2(n_1272),
.B(n_1341),
.Y(n_1445)
);

INVx4_ASAP7_75t_L g1446 ( 
.A(n_1280),
.Y(n_1446)
);

OAI21x1_ASAP7_75t_L g1447 ( 
.A1(n_1360),
.A2(n_1314),
.B(n_1354),
.Y(n_1447)
);

OR2x6_ASAP7_75t_L g1448 ( 
.A(n_1301),
.B(n_1302),
.Y(n_1448)
);

OAI21x1_ASAP7_75t_L g1449 ( 
.A1(n_1296),
.A2(n_1356),
.B(n_1282),
.Y(n_1449)
);

AOI221xp5_ASAP7_75t_L g1450 ( 
.A1(n_1419),
.A2(n_1335),
.B1(n_1357),
.B2(n_1361),
.C(n_1384),
.Y(n_1450)
);

INVx1_ASAP7_75t_L g1451 ( 
.A(n_1305),
.Y(n_1451)
);

OAI21x1_ASAP7_75t_L g1452 ( 
.A1(n_1288),
.A2(n_1276),
.B(n_1322),
.Y(n_1452)
);

INVx1_ASAP7_75t_L g1453 ( 
.A(n_1310),
.Y(n_1453)
);

CKINVDCx11_ASAP7_75t_R g1454 ( 
.A(n_1319),
.Y(n_1454)
);

AND2x2_ASAP7_75t_L g1455 ( 
.A(n_1359),
.B(n_1326),
.Y(n_1455)
);

HB1xp67_ASAP7_75t_L g1456 ( 
.A(n_1299),
.Y(n_1456)
);

OAI21x1_ASAP7_75t_L g1457 ( 
.A1(n_1362),
.A2(n_1358),
.B(n_1323),
.Y(n_1457)
);

O2A1O1Ixp33_ASAP7_75t_SL g1458 ( 
.A1(n_1334),
.A2(n_1355),
.B(n_1320),
.C(n_1344),
.Y(n_1458)
);

OAI21x1_ASAP7_75t_L g1459 ( 
.A1(n_1414),
.A2(n_1420),
.B(n_1343),
.Y(n_1459)
);

O2A1O1Ixp33_ASAP7_75t_SL g1460 ( 
.A1(n_1345),
.A2(n_1317),
.B(n_1373),
.C(n_1333),
.Y(n_1460)
);

BUFx6f_ASAP7_75t_L g1461 ( 
.A(n_1287),
.Y(n_1461)
);

AOI22xp5_ASAP7_75t_L g1462 ( 
.A1(n_1401),
.A2(n_1373),
.B1(n_1347),
.B2(n_1397),
.Y(n_1462)
);

NAND2xp5_ASAP7_75t_L g1463 ( 
.A(n_1412),
.B(n_1381),
.Y(n_1463)
);

OA21x2_ASAP7_75t_L g1464 ( 
.A1(n_1333),
.A2(n_1312),
.B(n_1315),
.Y(n_1464)
);

OAI21x1_ASAP7_75t_L g1465 ( 
.A1(n_1351),
.A2(n_1352),
.B(n_1297),
.Y(n_1465)
);

OAI21x1_ASAP7_75t_L g1466 ( 
.A1(n_1289),
.A2(n_1303),
.B(n_1369),
.Y(n_1466)
);

BUFx2_ASAP7_75t_L g1467 ( 
.A(n_1294),
.Y(n_1467)
);

INVx1_ASAP7_75t_L g1468 ( 
.A(n_1392),
.Y(n_1468)
);

OA21x2_ASAP7_75t_L g1469 ( 
.A1(n_1395),
.A2(n_1415),
.B(n_1410),
.Y(n_1469)
);

NAND2xp5_ASAP7_75t_L g1470 ( 
.A(n_1385),
.B(n_1406),
.Y(n_1470)
);

AOI22xp5_ASAP7_75t_L g1471 ( 
.A1(n_1374),
.A2(n_1337),
.B1(n_1371),
.B2(n_1377),
.Y(n_1471)
);

INVx1_ASAP7_75t_L g1472 ( 
.A(n_1308),
.Y(n_1472)
);

AOI22xp5_ASAP7_75t_L g1473 ( 
.A1(n_1330),
.A2(n_1387),
.B1(n_1417),
.B2(n_1416),
.Y(n_1473)
);

CKINVDCx5p33_ASAP7_75t_R g1474 ( 
.A(n_1318),
.Y(n_1474)
);

NAND2xp5_ASAP7_75t_SL g1475 ( 
.A(n_1386),
.B(n_1408),
.Y(n_1475)
);

O2A1O1Ixp33_ASAP7_75t_SL g1476 ( 
.A1(n_1389),
.A2(n_1393),
.B(n_1411),
.C(n_1340),
.Y(n_1476)
);

NAND2xp5_ASAP7_75t_L g1477 ( 
.A(n_1277),
.B(n_1380),
.Y(n_1477)
);

OAI21x1_ASAP7_75t_L g1478 ( 
.A1(n_1325),
.A2(n_1291),
.B(n_1363),
.Y(n_1478)
);

AOI22xp33_ASAP7_75t_L g1479 ( 
.A1(n_1339),
.A2(n_1396),
.B1(n_1293),
.B2(n_1409),
.Y(n_1479)
);

NOR2xp67_ASAP7_75t_L g1480 ( 
.A(n_1321),
.B(n_1366),
.Y(n_1480)
);

NAND2xp5_ASAP7_75t_L g1481 ( 
.A(n_1380),
.B(n_1346),
.Y(n_1481)
);

OAI21x1_ASAP7_75t_L g1482 ( 
.A1(n_1325),
.A2(n_1290),
.B(n_1304),
.Y(n_1482)
);

OAI21x1_ASAP7_75t_L g1483 ( 
.A1(n_1304),
.A2(n_1349),
.B(n_1383),
.Y(n_1483)
);

NOR2xp67_ASAP7_75t_SL g1484 ( 
.A(n_1368),
.B(n_1365),
.Y(n_1484)
);

INVx2_ASAP7_75t_L g1485 ( 
.A(n_1299),
.Y(n_1485)
);

OAI21x1_ASAP7_75t_L g1486 ( 
.A1(n_1383),
.A2(n_1407),
.B(n_1293),
.Y(n_1486)
);

O2A1O1Ixp33_ASAP7_75t_SL g1487 ( 
.A1(n_1407),
.A2(n_1295),
.B(n_1400),
.C(n_1405),
.Y(n_1487)
);

AO31x2_ASAP7_75t_L g1488 ( 
.A1(n_1368),
.A2(n_1399),
.A3(n_1328),
.B(n_1332),
.Y(n_1488)
);

NAND2xp5_ASAP7_75t_L g1489 ( 
.A(n_1298),
.B(n_1283),
.Y(n_1489)
);

O2A1O1Ixp33_ASAP7_75t_L g1490 ( 
.A1(n_1399),
.A2(n_1419),
.B(n_1388),
.C(n_1398),
.Y(n_1490)
);

INVx1_ASAP7_75t_L g1491 ( 
.A(n_1278),
.Y(n_1491)
);

NOR2xp33_ASAP7_75t_L g1492 ( 
.A(n_1419),
.B(n_1398),
.Y(n_1492)
);

O2A1O1Ixp33_ASAP7_75t_SL g1493 ( 
.A1(n_1399),
.A2(n_1388),
.B(n_1324),
.C(n_1124),
.Y(n_1493)
);

INVx1_ASAP7_75t_SL g1494 ( 
.A(n_1413),
.Y(n_1494)
);

AOI21x1_ASAP7_75t_L g1495 ( 
.A1(n_1307),
.A2(n_1282),
.B(n_1379),
.Y(n_1495)
);

OAI21xp5_ASAP7_75t_L g1496 ( 
.A1(n_1399),
.A2(n_1388),
.B(n_1316),
.Y(n_1496)
);

AO21x2_ASAP7_75t_L g1497 ( 
.A1(n_1388),
.A2(n_1275),
.B(n_1399),
.Y(n_1497)
);

BUFx12f_ASAP7_75t_L g1498 ( 
.A(n_1404),
.Y(n_1498)
);

OR2x2_ASAP7_75t_L g1499 ( 
.A(n_1376),
.B(n_1336),
.Y(n_1499)
);

NAND2xp5_ASAP7_75t_L g1500 ( 
.A(n_1298),
.B(n_1283),
.Y(n_1500)
);

NAND2xp5_ASAP7_75t_L g1501 ( 
.A(n_1298),
.B(n_1283),
.Y(n_1501)
);

BUFx6f_ASAP7_75t_L g1502 ( 
.A(n_1348),
.Y(n_1502)
);

AO21x2_ASAP7_75t_L g1503 ( 
.A1(n_1388),
.A2(n_1275),
.B(n_1399),
.Y(n_1503)
);

AOI21xp5_ASAP7_75t_L g1504 ( 
.A1(n_1399),
.A2(n_1403),
.B(n_1379),
.Y(n_1504)
);

OR2x2_ASAP7_75t_L g1505 ( 
.A(n_1376),
.B(n_1336),
.Y(n_1505)
);

OAI21x1_ASAP7_75t_L g1506 ( 
.A1(n_1309),
.A2(n_1382),
.B(n_1378),
.Y(n_1506)
);

INVx1_ASAP7_75t_L g1507 ( 
.A(n_1278),
.Y(n_1507)
);

BUFx10_ASAP7_75t_L g1508 ( 
.A(n_1418),
.Y(n_1508)
);

INVx1_ASAP7_75t_L g1509 ( 
.A(n_1278),
.Y(n_1509)
);

OAI21xp5_ASAP7_75t_L g1510 ( 
.A1(n_1399),
.A2(n_1388),
.B(n_1316),
.Y(n_1510)
);

AO21x2_ASAP7_75t_L g1511 ( 
.A1(n_1388),
.A2(n_1275),
.B(n_1399),
.Y(n_1511)
);

BUFx3_ASAP7_75t_L g1512 ( 
.A(n_1377),
.Y(n_1512)
);

AOI22xp5_ASAP7_75t_L g1513 ( 
.A1(n_1398),
.A2(n_785),
.B1(n_612),
.B2(n_426),
.Y(n_1513)
);

AOI22xp33_ASAP7_75t_L g1514 ( 
.A1(n_1398),
.A2(n_1388),
.B1(n_1229),
.B2(n_785),
.Y(n_1514)
);

INVx1_ASAP7_75t_L g1515 ( 
.A(n_1278),
.Y(n_1515)
);

AOI222xp33_ASAP7_75t_SL g1516 ( 
.A1(n_1398),
.A2(n_692),
.B1(n_1167),
.B2(n_1183),
.C1(n_1212),
.C2(n_707),
.Y(n_1516)
);

AND2x2_ASAP7_75t_L g1517 ( 
.A(n_1375),
.B(n_1281),
.Y(n_1517)
);

NAND2xp5_ASAP7_75t_L g1518 ( 
.A(n_1298),
.B(n_1283),
.Y(n_1518)
);

NAND2xp5_ASAP7_75t_SL g1519 ( 
.A(n_1398),
.B(n_1399),
.Y(n_1519)
);

INVx1_ASAP7_75t_L g1520 ( 
.A(n_1278),
.Y(n_1520)
);

CKINVDCx8_ASAP7_75t_R g1521 ( 
.A(n_1418),
.Y(n_1521)
);

AOI21x1_ASAP7_75t_L g1522 ( 
.A1(n_1307),
.A2(n_1282),
.B(n_1379),
.Y(n_1522)
);

AND2x4_ASAP7_75t_L g1523 ( 
.A(n_1391),
.B(n_1348),
.Y(n_1523)
);

NAND2xp5_ASAP7_75t_L g1524 ( 
.A(n_1298),
.B(n_1283),
.Y(n_1524)
);

AOI21xp5_ASAP7_75t_L g1525 ( 
.A1(n_1399),
.A2(n_1403),
.B(n_1379),
.Y(n_1525)
);

AOI22xp5_ASAP7_75t_L g1526 ( 
.A1(n_1398),
.A2(n_785),
.B1(n_612),
.B2(n_426),
.Y(n_1526)
);

AO31x2_ASAP7_75t_L g1527 ( 
.A1(n_1399),
.A2(n_1328),
.A3(n_1332),
.B(n_1272),
.Y(n_1527)
);

OAI21x1_ASAP7_75t_SL g1528 ( 
.A1(n_1372),
.A2(n_1327),
.B(n_1402),
.Y(n_1528)
);

AOI222xp33_ASAP7_75t_L g1529 ( 
.A1(n_1398),
.A2(n_1212),
.B1(n_1167),
.B2(n_1183),
.C1(n_1250),
.C2(n_1091),
.Y(n_1529)
);

OR2x2_ASAP7_75t_L g1530 ( 
.A(n_1376),
.B(n_1336),
.Y(n_1530)
);

AOI22xp33_ASAP7_75t_L g1531 ( 
.A1(n_1398),
.A2(n_1388),
.B1(n_1229),
.B2(n_785),
.Y(n_1531)
);

OAI22xp5_ASAP7_75t_L g1532 ( 
.A1(n_1398),
.A2(n_1399),
.B1(n_1224),
.B2(n_785),
.Y(n_1532)
);

NAND3xp33_ASAP7_75t_SL g1533 ( 
.A(n_1398),
.B(n_1419),
.C(n_1399),
.Y(n_1533)
);

AOI22xp33_ASAP7_75t_SL g1534 ( 
.A1(n_1357),
.A2(n_1183),
.B1(n_1212),
.B2(n_1250),
.Y(n_1534)
);

AO21x2_ASAP7_75t_L g1535 ( 
.A1(n_1388),
.A2(n_1275),
.B(n_1399),
.Y(n_1535)
);

AO21x2_ASAP7_75t_L g1536 ( 
.A1(n_1388),
.A2(n_1275),
.B(n_1399),
.Y(n_1536)
);

AOI22xp33_ASAP7_75t_SL g1537 ( 
.A1(n_1357),
.A2(n_1183),
.B1(n_1212),
.B2(n_1250),
.Y(n_1537)
);

OA21x2_ASAP7_75t_L g1538 ( 
.A1(n_1275),
.A2(n_1306),
.B(n_1378),
.Y(n_1538)
);

AOI322xp5_ASAP7_75t_L g1539 ( 
.A1(n_1398),
.A2(n_1250),
.A3(n_692),
.B1(n_835),
.B2(n_1091),
.C1(n_841),
.C2(n_763),
.Y(n_1539)
);

CKINVDCx5p33_ASAP7_75t_R g1540 ( 
.A(n_1418),
.Y(n_1540)
);

AO21x2_ASAP7_75t_L g1541 ( 
.A1(n_1388),
.A2(n_1275),
.B(n_1399),
.Y(n_1541)
);

INVx1_ASAP7_75t_L g1542 ( 
.A(n_1278),
.Y(n_1542)
);

INVx1_ASAP7_75t_L g1543 ( 
.A(n_1278),
.Y(n_1543)
);

NAND2xp5_ASAP7_75t_L g1544 ( 
.A(n_1298),
.B(n_1283),
.Y(n_1544)
);

AND2x2_ASAP7_75t_L g1545 ( 
.A(n_1455),
.B(n_1424),
.Y(n_1545)
);

O2A1O1Ixp33_ASAP7_75t_L g1546 ( 
.A1(n_1492),
.A2(n_1519),
.B(n_1533),
.C(n_1532),
.Y(n_1546)
);

NOR2xp33_ASAP7_75t_L g1547 ( 
.A(n_1431),
.B(n_1517),
.Y(n_1547)
);

BUFx3_ASAP7_75t_L g1548 ( 
.A(n_1467),
.Y(n_1548)
);

AND2x2_ASAP7_75t_L g1549 ( 
.A(n_1470),
.B(n_1450),
.Y(n_1549)
);

BUFx8_ASAP7_75t_SL g1550 ( 
.A(n_1498),
.Y(n_1550)
);

OA21x2_ASAP7_75t_L g1551 ( 
.A1(n_1457),
.A2(n_1452),
.B(n_1422),
.Y(n_1551)
);

HB1xp67_ASAP7_75t_L g1552 ( 
.A(n_1456),
.Y(n_1552)
);

AND2x2_ASAP7_75t_L g1553 ( 
.A(n_1450),
.B(n_1472),
.Y(n_1553)
);

O2A1O1Ixp5_ASAP7_75t_L g1554 ( 
.A1(n_1519),
.A2(n_1496),
.B(n_1510),
.C(n_1492),
.Y(n_1554)
);

CKINVDCx5p33_ASAP7_75t_R g1555 ( 
.A(n_1540),
.Y(n_1555)
);

AOI21xp5_ASAP7_75t_L g1556 ( 
.A1(n_1504),
.A2(n_1525),
.B(n_1493),
.Y(n_1556)
);

AND2x2_ASAP7_75t_L g1557 ( 
.A(n_1463),
.B(n_1462),
.Y(n_1557)
);

OAI22xp5_ASAP7_75t_L g1558 ( 
.A1(n_1534),
.A2(n_1537),
.B1(n_1513),
.B2(n_1526),
.Y(n_1558)
);

OAI22xp5_ASAP7_75t_L g1559 ( 
.A1(n_1534),
.A2(n_1537),
.B1(n_1531),
.B2(n_1514),
.Y(n_1559)
);

OR2x2_ASAP7_75t_L g1560 ( 
.A(n_1499),
.B(n_1505),
.Y(n_1560)
);

OA21x2_ASAP7_75t_L g1561 ( 
.A1(n_1504),
.A2(n_1525),
.B(n_1447),
.Y(n_1561)
);

AOI21xp5_ASAP7_75t_SL g1562 ( 
.A1(n_1532),
.A2(n_1490),
.B(n_1533),
.Y(n_1562)
);

OA21x2_ASAP7_75t_L g1563 ( 
.A1(n_1449),
.A2(n_1433),
.B(n_1425),
.Y(n_1563)
);

NAND2xp5_ASAP7_75t_L g1564 ( 
.A(n_1475),
.B(n_1427),
.Y(n_1564)
);

AND2x2_ASAP7_75t_L g1565 ( 
.A(n_1530),
.B(n_1475),
.Y(n_1565)
);

O2A1O1Ixp33_ASAP7_75t_L g1566 ( 
.A1(n_1490),
.A2(n_1436),
.B(n_1493),
.C(n_1531),
.Y(n_1566)
);

O2A1O1Ixp33_ASAP7_75t_L g1567 ( 
.A1(n_1436),
.A2(n_1514),
.B(n_1529),
.C(n_1476),
.Y(n_1567)
);

AOI21xp5_ASAP7_75t_SL g1568 ( 
.A1(n_1427),
.A2(n_1544),
.B(n_1518),
.Y(n_1568)
);

HB1xp67_ASAP7_75t_L g1569 ( 
.A(n_1456),
.Y(n_1569)
);

OAI22xp5_ASAP7_75t_L g1570 ( 
.A1(n_1479),
.A2(n_1544),
.B1(n_1489),
.B2(n_1500),
.Y(n_1570)
);

O2A1O1Ixp33_ASAP7_75t_L g1571 ( 
.A1(n_1529),
.A2(n_1476),
.B(n_1460),
.C(n_1458),
.Y(n_1571)
);

NAND2xp5_ASAP7_75t_L g1572 ( 
.A(n_1489),
.B(n_1500),
.Y(n_1572)
);

OAI211xp5_ASAP7_75t_L g1573 ( 
.A1(n_1539),
.A2(n_1460),
.B(n_1458),
.C(n_1516),
.Y(n_1573)
);

OAI22xp5_ASAP7_75t_L g1574 ( 
.A1(n_1479),
.A2(n_1524),
.B1(n_1501),
.B2(n_1428),
.Y(n_1574)
);

O2A1O1Ixp33_ASAP7_75t_L g1575 ( 
.A1(n_1501),
.A2(n_1524),
.B(n_1528),
.C(n_1487),
.Y(n_1575)
);

AOI21xp5_ASAP7_75t_SL g1576 ( 
.A1(n_1434),
.A2(n_1428),
.B(n_1523),
.Y(n_1576)
);

AOI21xp5_ASAP7_75t_L g1577 ( 
.A1(n_1440),
.A2(n_1445),
.B(n_1443),
.Y(n_1577)
);

NAND2xp5_ASAP7_75t_L g1578 ( 
.A(n_1441),
.B(n_1434),
.Y(n_1578)
);

NOR2xp33_ASAP7_75t_R g1579 ( 
.A(n_1429),
.B(n_1521),
.Y(n_1579)
);

AOI22xp5_ASAP7_75t_L g1580 ( 
.A1(n_1516),
.A2(n_1471),
.B1(n_1523),
.B2(n_1484),
.Y(n_1580)
);

AOI22xp5_ASAP7_75t_L g1581 ( 
.A1(n_1480),
.A2(n_1430),
.B1(n_1502),
.B2(n_1432),
.Y(n_1581)
);

CKINVDCx5p33_ASAP7_75t_R g1582 ( 
.A(n_1474),
.Y(n_1582)
);

CKINVDCx20_ASAP7_75t_R g1583 ( 
.A(n_1454),
.Y(n_1583)
);

OR2x2_ASAP7_75t_L g1584 ( 
.A(n_1442),
.B(n_1451),
.Y(n_1584)
);

INVx1_ASAP7_75t_L g1585 ( 
.A(n_1453),
.Y(n_1585)
);

O2A1O1Ixp33_ASAP7_75t_L g1586 ( 
.A1(n_1487),
.A2(n_1437),
.B(n_1448),
.C(n_1542),
.Y(n_1586)
);

INVxp33_ASAP7_75t_SL g1587 ( 
.A(n_1454),
.Y(n_1587)
);

OAI22xp5_ASAP7_75t_L g1588 ( 
.A1(n_1446),
.A2(n_1543),
.B1(n_1491),
.B2(n_1520),
.Y(n_1588)
);

OAI22xp5_ASAP7_75t_L g1589 ( 
.A1(n_1468),
.A2(n_1507),
.B1(n_1509),
.B2(n_1515),
.Y(n_1589)
);

NAND2xp5_ASAP7_75t_L g1590 ( 
.A(n_1448),
.B(n_1464),
.Y(n_1590)
);

OAI22xp5_ASAP7_75t_L g1591 ( 
.A1(n_1423),
.A2(n_1438),
.B1(n_1435),
.B2(n_1421),
.Y(n_1591)
);

O2A1O1Ixp5_ASAP7_75t_L g1592 ( 
.A1(n_1495),
.A2(n_1522),
.B(n_1485),
.C(n_1535),
.Y(n_1592)
);

BUFx3_ASAP7_75t_L g1593 ( 
.A(n_1512),
.Y(n_1593)
);

OAI22xp5_ASAP7_75t_L g1594 ( 
.A1(n_1423),
.A2(n_1438),
.B1(n_1435),
.B2(n_1421),
.Y(n_1594)
);

O2A1O1Ixp33_ASAP7_75t_L g1595 ( 
.A1(n_1448),
.A2(n_1541),
.B(n_1503),
.C(n_1511),
.Y(n_1595)
);

AOI21xp5_ASAP7_75t_L g1596 ( 
.A1(n_1440),
.A2(n_1445),
.B(n_1443),
.Y(n_1596)
);

OR2x2_ASAP7_75t_L g1597 ( 
.A(n_1497),
.B(n_1541),
.Y(n_1597)
);

INVx1_ASAP7_75t_L g1598 ( 
.A(n_1464),
.Y(n_1598)
);

O2A1O1Ixp33_ASAP7_75t_L g1599 ( 
.A1(n_1536),
.A2(n_1426),
.B(n_1538),
.C(n_1488),
.Y(n_1599)
);

NOR2xp67_ASAP7_75t_L g1600 ( 
.A(n_1439),
.B(n_1461),
.Y(n_1600)
);

AND2x4_ASAP7_75t_L g1601 ( 
.A(n_1478),
.B(n_1486),
.Y(n_1601)
);

AND2x2_ASAP7_75t_L g1602 ( 
.A(n_1488),
.B(n_1466),
.Y(n_1602)
);

BUFx3_ASAP7_75t_L g1603 ( 
.A(n_1508),
.Y(n_1603)
);

AND2x4_ASAP7_75t_L g1604 ( 
.A(n_1482),
.B(n_1483),
.Y(n_1604)
);

AOI21x1_ASAP7_75t_SL g1605 ( 
.A1(n_1527),
.A2(n_1444),
.B(n_1459),
.Y(n_1605)
);

INVx4_ASAP7_75t_L g1606 ( 
.A(n_1508),
.Y(n_1606)
);

NAND2xp5_ASAP7_75t_L g1607 ( 
.A(n_1527),
.B(n_1465),
.Y(n_1607)
);

INVx1_ASAP7_75t_L g1608 ( 
.A(n_1506),
.Y(n_1608)
);

O2A1O1Ixp33_ASAP7_75t_L g1609 ( 
.A1(n_1492),
.A2(n_1419),
.B(n_1399),
.C(n_1388),
.Y(n_1609)
);

OAI22xp5_ASAP7_75t_L g1610 ( 
.A1(n_1534),
.A2(n_1537),
.B1(n_1513),
.B2(n_1526),
.Y(n_1610)
);

NAND2xp5_ASAP7_75t_L g1611 ( 
.A(n_1470),
.B(n_1463),
.Y(n_1611)
);

NOR2xp67_ASAP7_75t_L g1612 ( 
.A(n_1473),
.B(n_1330),
.Y(n_1612)
);

NAND2xp5_ASAP7_75t_L g1613 ( 
.A(n_1470),
.B(n_1463),
.Y(n_1613)
);

O2A1O1Ixp33_ASAP7_75t_L g1614 ( 
.A1(n_1492),
.A2(n_1419),
.B(n_1399),
.C(n_1388),
.Y(n_1614)
);

O2A1O1Ixp5_ASAP7_75t_L g1615 ( 
.A1(n_1519),
.A2(n_1388),
.B(n_1399),
.C(n_1422),
.Y(n_1615)
);

NAND2xp5_ASAP7_75t_L g1616 ( 
.A(n_1470),
.B(n_1463),
.Y(n_1616)
);

CKINVDCx20_ASAP7_75t_R g1617 ( 
.A(n_1454),
.Y(n_1617)
);

O2A1O1Ixp5_ASAP7_75t_L g1618 ( 
.A1(n_1519),
.A2(n_1388),
.B(n_1399),
.C(n_1422),
.Y(n_1618)
);

HB1xp67_ASAP7_75t_L g1619 ( 
.A(n_1494),
.Y(n_1619)
);

OR2x2_ASAP7_75t_L g1620 ( 
.A(n_1499),
.B(n_1505),
.Y(n_1620)
);

AND2x2_ASAP7_75t_L g1621 ( 
.A(n_1455),
.B(n_1424),
.Y(n_1621)
);

AND2x2_ASAP7_75t_L g1622 ( 
.A(n_1455),
.B(n_1424),
.Y(n_1622)
);

CKINVDCx16_ASAP7_75t_R g1623 ( 
.A(n_1498),
.Y(n_1623)
);

INVx1_ASAP7_75t_L g1624 ( 
.A(n_1469),
.Y(n_1624)
);

AOI21xp5_ASAP7_75t_SL g1625 ( 
.A1(n_1532),
.A2(n_1399),
.B(n_1149),
.Y(n_1625)
);

NAND2xp5_ASAP7_75t_L g1626 ( 
.A(n_1470),
.B(n_1463),
.Y(n_1626)
);

BUFx6f_ASAP7_75t_L g1627 ( 
.A(n_1432),
.Y(n_1627)
);

OAI22xp5_ASAP7_75t_L g1628 ( 
.A1(n_1534),
.A2(n_1537),
.B1(n_1513),
.B2(n_1526),
.Y(n_1628)
);

NOR2xp33_ASAP7_75t_L g1629 ( 
.A(n_1431),
.B(n_421),
.Y(n_1629)
);

OAI22xp5_ASAP7_75t_L g1630 ( 
.A1(n_1534),
.A2(n_1537),
.B1(n_1513),
.B2(n_1526),
.Y(n_1630)
);

AND2x6_ASAP7_75t_L g1631 ( 
.A(n_1477),
.B(n_1481),
.Y(n_1631)
);

NAND2xp5_ASAP7_75t_L g1632 ( 
.A(n_1470),
.B(n_1463),
.Y(n_1632)
);

O2A1O1Ixp5_ASAP7_75t_L g1633 ( 
.A1(n_1519),
.A2(n_1388),
.B(n_1399),
.C(n_1422),
.Y(n_1633)
);

AOI21xp5_ASAP7_75t_L g1634 ( 
.A1(n_1504),
.A2(n_1399),
.B(n_1525),
.Y(n_1634)
);

NAND2xp5_ASAP7_75t_L g1635 ( 
.A(n_1470),
.B(n_1463),
.Y(n_1635)
);

AND2x2_ASAP7_75t_L g1636 ( 
.A(n_1455),
.B(n_1424),
.Y(n_1636)
);

AND2x2_ASAP7_75t_L g1637 ( 
.A(n_1455),
.B(n_1424),
.Y(n_1637)
);

OA21x2_ASAP7_75t_L g1638 ( 
.A1(n_1457),
.A2(n_1452),
.B(n_1422),
.Y(n_1638)
);

INVx1_ASAP7_75t_L g1639 ( 
.A(n_1469),
.Y(n_1639)
);

AOI21xp5_ASAP7_75t_L g1640 ( 
.A1(n_1504),
.A2(n_1399),
.B(n_1525),
.Y(n_1640)
);

O2A1O1Ixp33_ASAP7_75t_L g1641 ( 
.A1(n_1492),
.A2(n_1419),
.B(n_1399),
.C(n_1388),
.Y(n_1641)
);

OR2x2_ASAP7_75t_L g1642 ( 
.A(n_1499),
.B(n_1505),
.Y(n_1642)
);

INVxp67_ASAP7_75t_SL g1643 ( 
.A(n_1590),
.Y(n_1643)
);

HB1xp67_ASAP7_75t_L g1644 ( 
.A(n_1565),
.Y(n_1644)
);

OR2x6_ASAP7_75t_L g1645 ( 
.A(n_1634),
.B(n_1640),
.Y(n_1645)
);

OAI21x1_ASAP7_75t_L g1646 ( 
.A1(n_1605),
.A2(n_1592),
.B(n_1577),
.Y(n_1646)
);

INVx2_ASAP7_75t_L g1647 ( 
.A(n_1624),
.Y(n_1647)
);

INVx3_ASAP7_75t_L g1648 ( 
.A(n_1604),
.Y(n_1648)
);

AOI21xp33_ASAP7_75t_L g1649 ( 
.A1(n_1609),
.A2(n_1641),
.B(n_1614),
.Y(n_1649)
);

INVx2_ASAP7_75t_L g1650 ( 
.A(n_1639),
.Y(n_1650)
);

OR2x2_ASAP7_75t_L g1651 ( 
.A(n_1597),
.B(n_1598),
.Y(n_1651)
);

NAND2xp5_ASAP7_75t_L g1652 ( 
.A(n_1611),
.B(n_1613),
.Y(n_1652)
);

OR2x2_ASAP7_75t_L g1653 ( 
.A(n_1552),
.B(n_1569),
.Y(n_1653)
);

AO21x2_ASAP7_75t_L g1654 ( 
.A1(n_1596),
.A2(n_1640),
.B(n_1556),
.Y(n_1654)
);

INVx3_ASAP7_75t_L g1655 ( 
.A(n_1604),
.Y(n_1655)
);

INVxp67_ASAP7_75t_L g1656 ( 
.A(n_1547),
.Y(n_1656)
);

INVx2_ASAP7_75t_L g1657 ( 
.A(n_1608),
.Y(n_1657)
);

INVx2_ASAP7_75t_L g1658 ( 
.A(n_1551),
.Y(n_1658)
);

NAND2xp5_ASAP7_75t_L g1659 ( 
.A(n_1616),
.B(n_1626),
.Y(n_1659)
);

HB1xp67_ASAP7_75t_L g1660 ( 
.A(n_1619),
.Y(n_1660)
);

HB1xp67_ASAP7_75t_L g1661 ( 
.A(n_1588),
.Y(n_1661)
);

OR2x2_ASAP7_75t_L g1662 ( 
.A(n_1552),
.B(n_1569),
.Y(n_1662)
);

OA21x2_ASAP7_75t_L g1663 ( 
.A1(n_1592),
.A2(n_1556),
.B(n_1554),
.Y(n_1663)
);

INVxp67_ASAP7_75t_SL g1664 ( 
.A(n_1575),
.Y(n_1664)
);

NAND2xp5_ASAP7_75t_L g1665 ( 
.A(n_1632),
.B(n_1635),
.Y(n_1665)
);

AND2x2_ASAP7_75t_L g1666 ( 
.A(n_1602),
.B(n_1585),
.Y(n_1666)
);

HB1xp67_ASAP7_75t_L g1667 ( 
.A(n_1584),
.Y(n_1667)
);

INVx3_ASAP7_75t_L g1668 ( 
.A(n_1601),
.Y(n_1668)
);

AOI21xp5_ASAP7_75t_SL g1669 ( 
.A1(n_1571),
.A2(n_1567),
.B(n_1566),
.Y(n_1669)
);

INVx1_ASAP7_75t_L g1670 ( 
.A(n_1631),
.Y(n_1670)
);

AOI22xp5_ASAP7_75t_L g1671 ( 
.A1(n_1558),
.A2(n_1610),
.B1(n_1628),
.B2(n_1630),
.Y(n_1671)
);

HB1xp67_ASAP7_75t_L g1672 ( 
.A(n_1560),
.Y(n_1672)
);

OR2x6_ASAP7_75t_L g1673 ( 
.A(n_1576),
.B(n_1625),
.Y(n_1673)
);

AOI22xp33_ASAP7_75t_L g1674 ( 
.A1(n_1559),
.A2(n_1549),
.B1(n_1553),
.B2(n_1557),
.Y(n_1674)
);

AND2x2_ASAP7_75t_L g1675 ( 
.A(n_1638),
.B(n_1545),
.Y(n_1675)
);

AND2x2_ASAP7_75t_L g1676 ( 
.A(n_1638),
.B(n_1621),
.Y(n_1676)
);

INVx2_ASAP7_75t_L g1677 ( 
.A(n_1563),
.Y(n_1677)
);

NOR2x1_ASAP7_75t_R g1678 ( 
.A(n_1555),
.B(n_1582),
.Y(n_1678)
);

INVx3_ASAP7_75t_L g1679 ( 
.A(n_1601),
.Y(n_1679)
);

INVx1_ASAP7_75t_L g1680 ( 
.A(n_1589),
.Y(n_1680)
);

INVx3_ASAP7_75t_L g1681 ( 
.A(n_1563),
.Y(n_1681)
);

INVx3_ASAP7_75t_L g1682 ( 
.A(n_1561),
.Y(n_1682)
);

INVx1_ASAP7_75t_L g1683 ( 
.A(n_1607),
.Y(n_1683)
);

INVx1_ASAP7_75t_L g1684 ( 
.A(n_1554),
.Y(n_1684)
);

OA21x2_ASAP7_75t_L g1685 ( 
.A1(n_1615),
.A2(n_1618),
.B(n_1633),
.Y(n_1685)
);

AO21x2_ASAP7_75t_L g1686 ( 
.A1(n_1599),
.A2(n_1595),
.B(n_1562),
.Y(n_1686)
);

NAND2xp5_ASAP7_75t_L g1687 ( 
.A(n_1578),
.B(n_1572),
.Y(n_1687)
);

INVx1_ASAP7_75t_L g1688 ( 
.A(n_1564),
.Y(n_1688)
);

INVx1_ASAP7_75t_L g1689 ( 
.A(n_1591),
.Y(n_1689)
);

OR2x2_ASAP7_75t_L g1690 ( 
.A(n_1620),
.B(n_1642),
.Y(n_1690)
);

INVx1_ASAP7_75t_L g1691 ( 
.A(n_1594),
.Y(n_1691)
);

AO21x2_ASAP7_75t_L g1692 ( 
.A1(n_1595),
.A2(n_1641),
.B(n_1614),
.Y(n_1692)
);

INVx1_ASAP7_75t_L g1693 ( 
.A(n_1586),
.Y(n_1693)
);

INVx2_ASAP7_75t_L g1694 ( 
.A(n_1615),
.Y(n_1694)
);

INVx1_ASAP7_75t_L g1695 ( 
.A(n_1586),
.Y(n_1695)
);

OAI21xp5_ASAP7_75t_L g1696 ( 
.A1(n_1609),
.A2(n_1546),
.B(n_1633),
.Y(n_1696)
);

NAND2xp5_ASAP7_75t_L g1697 ( 
.A(n_1643),
.B(n_1546),
.Y(n_1697)
);

INVx1_ASAP7_75t_L g1698 ( 
.A(n_1647),
.Y(n_1698)
);

INVx2_ASAP7_75t_L g1699 ( 
.A(n_1657),
.Y(n_1699)
);

INVx1_ASAP7_75t_L g1700 ( 
.A(n_1647),
.Y(n_1700)
);

AOI22xp33_ASAP7_75t_L g1701 ( 
.A1(n_1671),
.A2(n_1574),
.B1(n_1570),
.B2(n_1612),
.Y(n_1701)
);

HB1xp67_ASAP7_75t_L g1702 ( 
.A(n_1651),
.Y(n_1702)
);

INVx1_ASAP7_75t_L g1703 ( 
.A(n_1650),
.Y(n_1703)
);

NAND2xp5_ASAP7_75t_L g1704 ( 
.A(n_1684),
.B(n_1688),
.Y(n_1704)
);

AND2x2_ASAP7_75t_L g1705 ( 
.A(n_1675),
.B(n_1618),
.Y(n_1705)
);

AND2x2_ASAP7_75t_L g1706 ( 
.A(n_1675),
.B(n_1637),
.Y(n_1706)
);

INVx3_ASAP7_75t_L g1707 ( 
.A(n_1648),
.Y(n_1707)
);

AND2x4_ASAP7_75t_L g1708 ( 
.A(n_1668),
.B(n_1679),
.Y(n_1708)
);

NAND2xp5_ASAP7_75t_L g1709 ( 
.A(n_1684),
.B(n_1568),
.Y(n_1709)
);

BUFx6f_ASAP7_75t_L g1710 ( 
.A(n_1645),
.Y(n_1710)
);

BUFx2_ASAP7_75t_L g1711 ( 
.A(n_1670),
.Y(n_1711)
);

AND2x2_ASAP7_75t_L g1712 ( 
.A(n_1676),
.B(n_1622),
.Y(n_1712)
);

AND2x2_ASAP7_75t_L g1713 ( 
.A(n_1676),
.B(n_1636),
.Y(n_1713)
);

BUFx3_ASAP7_75t_L g1714 ( 
.A(n_1668),
.Y(n_1714)
);

INVx4_ASAP7_75t_R g1715 ( 
.A(n_1670),
.Y(n_1715)
);

INVx4_ASAP7_75t_L g1716 ( 
.A(n_1673),
.Y(n_1716)
);

OA21x2_ASAP7_75t_L g1717 ( 
.A1(n_1646),
.A2(n_1573),
.B(n_1605),
.Y(n_1717)
);

NAND2xp5_ASAP7_75t_L g1718 ( 
.A(n_1688),
.B(n_1575),
.Y(n_1718)
);

OR2x2_ASAP7_75t_L g1719 ( 
.A(n_1653),
.B(n_1548),
.Y(n_1719)
);

HB1xp67_ASAP7_75t_L g1720 ( 
.A(n_1662),
.Y(n_1720)
);

AND2x2_ASAP7_75t_L g1721 ( 
.A(n_1666),
.B(n_1566),
.Y(n_1721)
);

OAI22xp5_ASAP7_75t_SL g1722 ( 
.A1(n_1671),
.A2(n_1580),
.B1(n_1583),
.B2(n_1617),
.Y(n_1722)
);

INVx2_ASAP7_75t_L g1723 ( 
.A(n_1677),
.Y(n_1723)
);

AOI22xp5_ASAP7_75t_L g1724 ( 
.A1(n_1674),
.A2(n_1573),
.B1(n_1629),
.B2(n_1581),
.Y(n_1724)
);

AND2x2_ASAP7_75t_L g1725 ( 
.A(n_1648),
.B(n_1655),
.Y(n_1725)
);

INVx1_ASAP7_75t_L g1726 ( 
.A(n_1698),
.Y(n_1726)
);

INVx1_ASAP7_75t_L g1727 ( 
.A(n_1698),
.Y(n_1727)
);

INVx2_ASAP7_75t_SL g1728 ( 
.A(n_1714),
.Y(n_1728)
);

AND2x2_ASAP7_75t_L g1729 ( 
.A(n_1706),
.B(n_1644),
.Y(n_1729)
);

OAI31xp33_ASAP7_75t_L g1730 ( 
.A1(n_1722),
.A2(n_1649),
.A3(n_1567),
.B(n_1664),
.Y(n_1730)
);

AOI22xp33_ASAP7_75t_L g1731 ( 
.A1(n_1722),
.A2(n_1696),
.B1(n_1673),
.B2(n_1645),
.Y(n_1731)
);

OAI22xp33_ASAP7_75t_L g1732 ( 
.A1(n_1724),
.A2(n_1673),
.B1(n_1645),
.B2(n_1685),
.Y(n_1732)
);

AOI22xp33_ASAP7_75t_L g1733 ( 
.A1(n_1701),
.A2(n_1673),
.B1(n_1645),
.B2(n_1692),
.Y(n_1733)
);

AND2x2_ASAP7_75t_L g1734 ( 
.A(n_1706),
.B(n_1672),
.Y(n_1734)
);

INVx1_ASAP7_75t_L g1735 ( 
.A(n_1698),
.Y(n_1735)
);

AOI22xp33_ASAP7_75t_L g1736 ( 
.A1(n_1701),
.A2(n_1673),
.B1(n_1645),
.B2(n_1692),
.Y(n_1736)
);

INVx1_ASAP7_75t_L g1737 ( 
.A(n_1700),
.Y(n_1737)
);

AOI22xp33_ASAP7_75t_L g1738 ( 
.A1(n_1697),
.A2(n_1692),
.B1(n_1685),
.B2(n_1689),
.Y(n_1738)
);

INVx1_ASAP7_75t_L g1739 ( 
.A(n_1700),
.Y(n_1739)
);

NOR4xp25_ASAP7_75t_SL g1740 ( 
.A(n_1711),
.B(n_1695),
.C(n_1693),
.D(n_1689),
.Y(n_1740)
);

AND2x4_ASAP7_75t_L g1741 ( 
.A(n_1708),
.B(n_1714),
.Y(n_1741)
);

BUFx2_ASAP7_75t_L g1742 ( 
.A(n_1714),
.Y(n_1742)
);

OAI221xp5_ASAP7_75t_L g1743 ( 
.A1(n_1724),
.A2(n_1669),
.B1(n_1685),
.B2(n_1694),
.C(n_1661),
.Y(n_1743)
);

HB1xp67_ASAP7_75t_L g1744 ( 
.A(n_1720),
.Y(n_1744)
);

NOR2xp33_ASAP7_75t_R g1745 ( 
.A(n_1697),
.B(n_1623),
.Y(n_1745)
);

CKINVDCx5p33_ASAP7_75t_R g1746 ( 
.A(n_1719),
.Y(n_1746)
);

NAND2xp5_ASAP7_75t_L g1747 ( 
.A(n_1704),
.B(n_1694),
.Y(n_1747)
);

OAI211xp5_ASAP7_75t_L g1748 ( 
.A1(n_1709),
.A2(n_1669),
.B(n_1685),
.C(n_1718),
.Y(n_1748)
);

AOI221xp5_ASAP7_75t_L g1749 ( 
.A1(n_1709),
.A2(n_1656),
.B1(n_1694),
.B2(n_1695),
.C(n_1693),
.Y(n_1749)
);

BUFx2_ASAP7_75t_L g1750 ( 
.A(n_1714),
.Y(n_1750)
);

OA21x2_ASAP7_75t_L g1751 ( 
.A1(n_1723),
.A2(n_1646),
.B(n_1658),
.Y(n_1751)
);

OAI21xp5_ASAP7_75t_L g1752 ( 
.A1(n_1718),
.A2(n_1691),
.B(n_1680),
.Y(n_1752)
);

NOR2x1_ASAP7_75t_L g1753 ( 
.A(n_1704),
.B(n_1716),
.Y(n_1753)
);

AND2x2_ASAP7_75t_L g1754 ( 
.A(n_1712),
.B(n_1713),
.Y(n_1754)
);

AND2x2_ASAP7_75t_L g1755 ( 
.A(n_1712),
.B(n_1655),
.Y(n_1755)
);

AOI222xp33_ASAP7_75t_L g1756 ( 
.A1(n_1721),
.A2(n_1587),
.B1(n_1652),
.B2(n_1665),
.C1(n_1659),
.C2(n_1687),
.Y(n_1756)
);

NAND2xp5_ASAP7_75t_L g1757 ( 
.A(n_1705),
.B(n_1667),
.Y(n_1757)
);

AOI22xp33_ASAP7_75t_L g1758 ( 
.A1(n_1710),
.A2(n_1691),
.B1(n_1686),
.B2(n_1690),
.Y(n_1758)
);

AND2x2_ASAP7_75t_L g1759 ( 
.A(n_1713),
.B(n_1655),
.Y(n_1759)
);

OAI21x1_ASAP7_75t_L g1760 ( 
.A1(n_1707),
.A2(n_1682),
.B(n_1681),
.Y(n_1760)
);

NAND3xp33_ASAP7_75t_L g1761 ( 
.A(n_1717),
.B(n_1660),
.C(n_1663),
.Y(n_1761)
);

INVx2_ASAP7_75t_L g1762 ( 
.A(n_1699),
.Y(n_1762)
);

NAND2xp5_ASAP7_75t_L g1763 ( 
.A(n_1705),
.B(n_1683),
.Y(n_1763)
);

INVx1_ASAP7_75t_L g1764 ( 
.A(n_1726),
.Y(n_1764)
);

AND2x2_ASAP7_75t_L g1765 ( 
.A(n_1754),
.B(n_1713),
.Y(n_1765)
);

AND2x2_ASAP7_75t_L g1766 ( 
.A(n_1754),
.B(n_1725),
.Y(n_1766)
);

INVx2_ASAP7_75t_L g1767 ( 
.A(n_1751),
.Y(n_1767)
);

OA21x2_ASAP7_75t_L g1768 ( 
.A1(n_1760),
.A2(n_1761),
.B(n_1738),
.Y(n_1768)
);

NOR2xp33_ASAP7_75t_L g1769 ( 
.A(n_1746),
.B(n_1606),
.Y(n_1769)
);

AOI21xp5_ASAP7_75t_L g1770 ( 
.A1(n_1732),
.A2(n_1686),
.B(n_1654),
.Y(n_1770)
);

AOI21x1_ASAP7_75t_L g1771 ( 
.A1(n_1742),
.A2(n_1711),
.B(n_1703),
.Y(n_1771)
);

INVx1_ASAP7_75t_L g1772 ( 
.A(n_1726),
.Y(n_1772)
);

INVx1_ASAP7_75t_L g1773 ( 
.A(n_1727),
.Y(n_1773)
);

INVx4_ASAP7_75t_L g1774 ( 
.A(n_1742),
.Y(n_1774)
);

BUFx3_ASAP7_75t_L g1775 ( 
.A(n_1750),
.Y(n_1775)
);

BUFx2_ASAP7_75t_L g1776 ( 
.A(n_1753),
.Y(n_1776)
);

INVx2_ASAP7_75t_L g1777 ( 
.A(n_1751),
.Y(n_1777)
);

OAI21xp5_ASAP7_75t_L g1778 ( 
.A1(n_1730),
.A2(n_1721),
.B(n_1717),
.Y(n_1778)
);

OR2x2_ASAP7_75t_L g1779 ( 
.A(n_1763),
.B(n_1702),
.Y(n_1779)
);

INVx1_ASAP7_75t_L g1780 ( 
.A(n_1727),
.Y(n_1780)
);

INVx1_ASAP7_75t_L g1781 ( 
.A(n_1735),
.Y(n_1781)
);

INVx2_ASAP7_75t_L g1782 ( 
.A(n_1751),
.Y(n_1782)
);

INVx1_ASAP7_75t_L g1783 ( 
.A(n_1735),
.Y(n_1783)
);

INVx1_ASAP7_75t_L g1784 ( 
.A(n_1737),
.Y(n_1784)
);

INVx2_ASAP7_75t_L g1785 ( 
.A(n_1751),
.Y(n_1785)
);

NOR2x1p5_ASAP7_75t_L g1786 ( 
.A(n_1757),
.B(n_1716),
.Y(n_1786)
);

INVx4_ASAP7_75t_SL g1787 ( 
.A(n_1750),
.Y(n_1787)
);

INVx4_ASAP7_75t_SL g1788 ( 
.A(n_1728),
.Y(n_1788)
);

INVx4_ASAP7_75t_SL g1789 ( 
.A(n_1741),
.Y(n_1789)
);

INVxp67_ASAP7_75t_SL g1790 ( 
.A(n_1747),
.Y(n_1790)
);

NAND2x1_ASAP7_75t_L g1791 ( 
.A(n_1739),
.B(n_1715),
.Y(n_1791)
);

HB1xp67_ASAP7_75t_L g1792 ( 
.A(n_1764),
.Y(n_1792)
);

NAND2xp5_ASAP7_75t_L g1793 ( 
.A(n_1790),
.B(n_1763),
.Y(n_1793)
);

INVx2_ASAP7_75t_L g1794 ( 
.A(n_1767),
.Y(n_1794)
);

INVx2_ASAP7_75t_SL g1795 ( 
.A(n_1791),
.Y(n_1795)
);

INVx1_ASAP7_75t_L g1796 ( 
.A(n_1764),
.Y(n_1796)
);

BUFx3_ASAP7_75t_L g1797 ( 
.A(n_1775),
.Y(n_1797)
);

INVx3_ASAP7_75t_SL g1798 ( 
.A(n_1787),
.Y(n_1798)
);

NAND2xp5_ASAP7_75t_L g1799 ( 
.A(n_1790),
.B(n_1757),
.Y(n_1799)
);

AND2x2_ASAP7_75t_L g1800 ( 
.A(n_1787),
.B(n_1755),
.Y(n_1800)
);

AND2x2_ASAP7_75t_L g1801 ( 
.A(n_1787),
.B(n_1759),
.Y(n_1801)
);

INVx2_ASAP7_75t_SL g1802 ( 
.A(n_1791),
.Y(n_1802)
);

AND2x2_ASAP7_75t_L g1803 ( 
.A(n_1787),
.B(n_1759),
.Y(n_1803)
);

INVx2_ASAP7_75t_L g1804 ( 
.A(n_1767),
.Y(n_1804)
);

INVx2_ASAP7_75t_L g1805 ( 
.A(n_1767),
.Y(n_1805)
);

INVx2_ASAP7_75t_L g1806 ( 
.A(n_1777),
.Y(n_1806)
);

AND2x2_ASAP7_75t_L g1807 ( 
.A(n_1787),
.B(n_1762),
.Y(n_1807)
);

NAND2xp5_ASAP7_75t_L g1808 ( 
.A(n_1765),
.B(n_1779),
.Y(n_1808)
);

INVx3_ASAP7_75t_L g1809 ( 
.A(n_1771),
.Y(n_1809)
);

INVx1_ASAP7_75t_L g1810 ( 
.A(n_1772),
.Y(n_1810)
);

INVx2_ASAP7_75t_L g1811 ( 
.A(n_1777),
.Y(n_1811)
);

INVx2_ASAP7_75t_L g1812 ( 
.A(n_1777),
.Y(n_1812)
);

AND2x2_ASAP7_75t_L g1813 ( 
.A(n_1788),
.B(n_1744),
.Y(n_1813)
);

NAND2xp5_ASAP7_75t_L g1814 ( 
.A(n_1765),
.B(n_1752),
.Y(n_1814)
);

OAI22xp5_ASAP7_75t_L g1815 ( 
.A1(n_1778),
.A2(n_1743),
.B1(n_1736),
.B2(n_1733),
.Y(n_1815)
);

NAND4xp25_ASAP7_75t_L g1816 ( 
.A(n_1778),
.B(n_1730),
.C(n_1756),
.D(n_1743),
.Y(n_1816)
);

INVx2_ASAP7_75t_L g1817 ( 
.A(n_1782),
.Y(n_1817)
);

AND2x2_ASAP7_75t_L g1818 ( 
.A(n_1788),
.B(n_1729),
.Y(n_1818)
);

NAND2xp5_ASAP7_75t_L g1819 ( 
.A(n_1779),
.B(n_1752),
.Y(n_1819)
);

NAND2xp5_ASAP7_75t_L g1820 ( 
.A(n_1779),
.B(n_1756),
.Y(n_1820)
);

AND2x2_ASAP7_75t_L g1821 ( 
.A(n_1788),
.B(n_1729),
.Y(n_1821)
);

INVx2_ASAP7_75t_L g1822 ( 
.A(n_1782),
.Y(n_1822)
);

HB1xp67_ASAP7_75t_L g1823 ( 
.A(n_1772),
.Y(n_1823)
);

INVx2_ASAP7_75t_L g1824 ( 
.A(n_1785),
.Y(n_1824)
);

INVx1_ASAP7_75t_L g1825 ( 
.A(n_1773),
.Y(n_1825)
);

NAND2xp5_ASAP7_75t_L g1826 ( 
.A(n_1780),
.B(n_1734),
.Y(n_1826)
);

INVx2_ASAP7_75t_L g1827 ( 
.A(n_1785),
.Y(n_1827)
);

OAI22xp5_ASAP7_75t_L g1828 ( 
.A1(n_1770),
.A2(n_1731),
.B1(n_1748),
.B2(n_1740),
.Y(n_1828)
);

AND2x2_ASAP7_75t_L g1829 ( 
.A(n_1798),
.B(n_1789),
.Y(n_1829)
);

NAND2xp5_ASAP7_75t_L g1830 ( 
.A(n_1820),
.B(n_1749),
.Y(n_1830)
);

AND2x2_ASAP7_75t_L g1831 ( 
.A(n_1798),
.B(n_1818),
.Y(n_1831)
);

OR2x2_ASAP7_75t_L g1832 ( 
.A(n_1814),
.B(n_1781),
.Y(n_1832)
);

NAND2x1p5_ASAP7_75t_L g1833 ( 
.A(n_1797),
.B(n_1776),
.Y(n_1833)
);

INVx1_ASAP7_75t_L g1834 ( 
.A(n_1792),
.Y(n_1834)
);

NAND2xp5_ASAP7_75t_L g1835 ( 
.A(n_1820),
.B(n_1766),
.Y(n_1835)
);

OR2x2_ASAP7_75t_L g1836 ( 
.A(n_1814),
.B(n_1781),
.Y(n_1836)
);

AND2x2_ASAP7_75t_L g1837 ( 
.A(n_1798),
.B(n_1789),
.Y(n_1837)
);

INVxp33_ASAP7_75t_L g1838 ( 
.A(n_1816),
.Y(n_1838)
);

INVx2_ASAP7_75t_L g1839 ( 
.A(n_1797),
.Y(n_1839)
);

INVx1_ASAP7_75t_L g1840 ( 
.A(n_1792),
.Y(n_1840)
);

INVx1_ASAP7_75t_L g1841 ( 
.A(n_1823),
.Y(n_1841)
);

HB1xp67_ASAP7_75t_L g1842 ( 
.A(n_1797),
.Y(n_1842)
);

OR2x2_ASAP7_75t_L g1843 ( 
.A(n_1819),
.B(n_1783),
.Y(n_1843)
);

INVx1_ASAP7_75t_L g1844 ( 
.A(n_1823),
.Y(n_1844)
);

OR2x2_ASAP7_75t_L g1845 ( 
.A(n_1819),
.B(n_1783),
.Y(n_1845)
);

AND2x2_ASAP7_75t_L g1846 ( 
.A(n_1798),
.B(n_1789),
.Y(n_1846)
);

AND2x4_ASAP7_75t_SL g1847 ( 
.A(n_1800),
.B(n_1774),
.Y(n_1847)
);

INVx2_ASAP7_75t_L g1848 ( 
.A(n_1797),
.Y(n_1848)
);

OR2x2_ASAP7_75t_L g1849 ( 
.A(n_1808),
.B(n_1784),
.Y(n_1849)
);

NAND2xp5_ASAP7_75t_L g1850 ( 
.A(n_1816),
.B(n_1766),
.Y(n_1850)
);

INVx1_ASAP7_75t_L g1851 ( 
.A(n_1796),
.Y(n_1851)
);

AND2x2_ASAP7_75t_L g1852 ( 
.A(n_1818),
.B(n_1789),
.Y(n_1852)
);

AND2x2_ASAP7_75t_L g1853 ( 
.A(n_1818),
.B(n_1821),
.Y(n_1853)
);

NAND2x1p5_ASAP7_75t_L g1854 ( 
.A(n_1795),
.B(n_1776),
.Y(n_1854)
);

INVx1_ASAP7_75t_L g1855 ( 
.A(n_1796),
.Y(n_1855)
);

OR2x2_ASAP7_75t_L g1856 ( 
.A(n_1808),
.B(n_1784),
.Y(n_1856)
);

INVx1_ASAP7_75t_L g1857 ( 
.A(n_1796),
.Y(n_1857)
);

HB1xp67_ASAP7_75t_L g1858 ( 
.A(n_1810),
.Y(n_1858)
);

INVx2_ASAP7_75t_L g1859 ( 
.A(n_1794),
.Y(n_1859)
);

AND2x2_ASAP7_75t_L g1860 ( 
.A(n_1821),
.B(n_1789),
.Y(n_1860)
);

AOI31xp33_ASAP7_75t_L g1861 ( 
.A1(n_1828),
.A2(n_1678),
.A3(n_1769),
.B(n_1758),
.Y(n_1861)
);

INVx1_ASAP7_75t_SL g1862 ( 
.A(n_1800),
.Y(n_1862)
);

INVx1_ASAP7_75t_L g1863 ( 
.A(n_1810),
.Y(n_1863)
);

NOR2xp33_ASAP7_75t_L g1864 ( 
.A(n_1815),
.B(n_1550),
.Y(n_1864)
);

OAI22xp33_ASAP7_75t_SL g1865 ( 
.A1(n_1815),
.A2(n_1776),
.B1(n_1774),
.B2(n_1775),
.Y(n_1865)
);

INVxp67_ASAP7_75t_L g1866 ( 
.A(n_1842),
.Y(n_1866)
);

INVx1_ASAP7_75t_SL g1867 ( 
.A(n_1847),
.Y(n_1867)
);

INVx1_ASAP7_75t_L g1868 ( 
.A(n_1858),
.Y(n_1868)
);

INVx3_ASAP7_75t_L g1869 ( 
.A(n_1854),
.Y(n_1869)
);

INVx1_ASAP7_75t_L g1870 ( 
.A(n_1855),
.Y(n_1870)
);

NAND2xp5_ASAP7_75t_L g1871 ( 
.A(n_1830),
.B(n_1826),
.Y(n_1871)
);

CKINVDCx16_ASAP7_75t_R g1872 ( 
.A(n_1864),
.Y(n_1872)
);

AND2x2_ASAP7_75t_L g1873 ( 
.A(n_1853),
.B(n_1795),
.Y(n_1873)
);

AOI22xp33_ASAP7_75t_SL g1874 ( 
.A1(n_1865),
.A2(n_1828),
.B1(n_1745),
.B2(n_1770),
.Y(n_1874)
);

AND2x2_ASAP7_75t_L g1875 ( 
.A(n_1853),
.B(n_1795),
.Y(n_1875)
);

NOR2x1p5_ASAP7_75t_L g1876 ( 
.A(n_1850),
.B(n_1835),
.Y(n_1876)
);

INVx2_ASAP7_75t_SL g1877 ( 
.A(n_1847),
.Y(n_1877)
);

AND2x2_ASAP7_75t_L g1878 ( 
.A(n_1852),
.B(n_1795),
.Y(n_1878)
);

NAND2xp5_ASAP7_75t_L g1879 ( 
.A(n_1838),
.B(n_1826),
.Y(n_1879)
);

INVx1_ASAP7_75t_L g1880 ( 
.A(n_1855),
.Y(n_1880)
);

CKINVDCx16_ASAP7_75t_R g1881 ( 
.A(n_1831),
.Y(n_1881)
);

INVx1_ASAP7_75t_L g1882 ( 
.A(n_1851),
.Y(n_1882)
);

NAND2x1_ASAP7_75t_SL g1883 ( 
.A(n_1829),
.B(n_1809),
.Y(n_1883)
);

INVx1_ASAP7_75t_L g1884 ( 
.A(n_1841),
.Y(n_1884)
);

INVx1_ASAP7_75t_SL g1885 ( 
.A(n_1831),
.Y(n_1885)
);

INVx1_ASAP7_75t_SL g1886 ( 
.A(n_1829),
.Y(n_1886)
);

INVx1_ASAP7_75t_L g1887 ( 
.A(n_1841),
.Y(n_1887)
);

INVx1_ASAP7_75t_L g1888 ( 
.A(n_1857),
.Y(n_1888)
);

HB1xp67_ASAP7_75t_L g1889 ( 
.A(n_1833),
.Y(n_1889)
);

AND2x2_ASAP7_75t_L g1890 ( 
.A(n_1852),
.B(n_1802),
.Y(n_1890)
);

INVxp67_ASAP7_75t_SL g1891 ( 
.A(n_1833),
.Y(n_1891)
);

OAI22xp5_ASAP7_75t_L g1892 ( 
.A1(n_1861),
.A2(n_1802),
.B1(n_1786),
.B2(n_1740),
.Y(n_1892)
);

INVx1_ASAP7_75t_L g1893 ( 
.A(n_1844),
.Y(n_1893)
);

NOR2xp33_ASAP7_75t_L g1894 ( 
.A(n_1872),
.B(n_1678),
.Y(n_1894)
);

AOI22xp33_ASAP7_75t_L g1895 ( 
.A1(n_1874),
.A2(n_1862),
.B1(n_1860),
.B2(n_1837),
.Y(n_1895)
);

AOI22xp5_ASAP7_75t_L g1896 ( 
.A1(n_1881),
.A2(n_1860),
.B1(n_1837),
.B2(n_1846),
.Y(n_1896)
);

INVx1_ASAP7_75t_L g1897 ( 
.A(n_1870),
.Y(n_1897)
);

NOR4xp25_ASAP7_75t_L g1898 ( 
.A(n_1866),
.B(n_1839),
.C(n_1848),
.D(n_1840),
.Y(n_1898)
);

INVx1_ASAP7_75t_L g1899 ( 
.A(n_1870),
.Y(n_1899)
);

INVx1_ASAP7_75t_L g1900 ( 
.A(n_1868),
.Y(n_1900)
);

AOI322xp5_ASAP7_75t_L g1901 ( 
.A1(n_1879),
.A2(n_1834),
.A3(n_1844),
.B1(n_1809),
.B2(n_1799),
.C1(n_1793),
.C2(n_1848),
.Y(n_1901)
);

OR2x2_ASAP7_75t_L g1902 ( 
.A(n_1885),
.B(n_1839),
.Y(n_1902)
);

AOI22xp5_ASAP7_75t_L g1903 ( 
.A1(n_1867),
.A2(n_1846),
.B1(n_1802),
.B2(n_1800),
.Y(n_1903)
);

AOI321xp33_ASAP7_75t_SL g1904 ( 
.A1(n_1886),
.A2(n_1769),
.A3(n_1833),
.B1(n_1854),
.B2(n_1856),
.C(n_1849),
.Y(n_1904)
);

NAND2xp5_ASAP7_75t_L g1905 ( 
.A(n_1868),
.B(n_1876),
.Y(n_1905)
);

INVx1_ASAP7_75t_L g1906 ( 
.A(n_1880),
.Y(n_1906)
);

AOI21xp5_ASAP7_75t_L g1907 ( 
.A1(n_1871),
.A2(n_1854),
.B(n_1802),
.Y(n_1907)
);

INVx1_ASAP7_75t_L g1908 ( 
.A(n_1884),
.Y(n_1908)
);

OAI22xp5_ASAP7_75t_L g1909 ( 
.A1(n_1891),
.A2(n_1809),
.B1(n_1768),
.B2(n_1774),
.Y(n_1909)
);

O2A1O1Ixp5_ASAP7_75t_SL g1910 ( 
.A1(n_1884),
.A2(n_1863),
.B(n_1809),
.C(n_1825),
.Y(n_1910)
);

INVx1_ASAP7_75t_L g1911 ( 
.A(n_1887),
.Y(n_1911)
);

NOR2xp33_ASAP7_75t_L g1912 ( 
.A(n_1877),
.B(n_1606),
.Y(n_1912)
);

AOI32xp33_ASAP7_75t_L g1913 ( 
.A1(n_1892),
.A2(n_1809),
.A3(n_1801),
.B1(n_1803),
.B2(n_1813),
.Y(n_1913)
);

INVx1_ASAP7_75t_L g1914 ( 
.A(n_1887),
.Y(n_1914)
);

INVx2_ASAP7_75t_L g1915 ( 
.A(n_1869),
.Y(n_1915)
);

NOR2xp33_ASAP7_75t_L g1916 ( 
.A(n_1894),
.B(n_1877),
.Y(n_1916)
);

NAND2xp5_ASAP7_75t_L g1917 ( 
.A(n_1898),
.B(n_1878),
.Y(n_1917)
);

AND2x4_ASAP7_75t_L g1918 ( 
.A(n_1896),
.B(n_1878),
.Y(n_1918)
);

INVx1_ASAP7_75t_L g1919 ( 
.A(n_1897),
.Y(n_1919)
);

INVx2_ASAP7_75t_L g1920 ( 
.A(n_1915),
.Y(n_1920)
);

OR2x2_ASAP7_75t_L g1921 ( 
.A(n_1902),
.B(n_1893),
.Y(n_1921)
);

INVx1_ASAP7_75t_L g1922 ( 
.A(n_1899),
.Y(n_1922)
);

OR2x2_ASAP7_75t_L g1923 ( 
.A(n_1905),
.B(n_1893),
.Y(n_1923)
);

INVx1_ASAP7_75t_L g1924 ( 
.A(n_1908),
.Y(n_1924)
);

NOR2x1_ASAP7_75t_L g1925 ( 
.A(n_1911),
.B(n_1869),
.Y(n_1925)
);

NAND2xp5_ASAP7_75t_L g1926 ( 
.A(n_1905),
.B(n_1890),
.Y(n_1926)
);

AND2x2_ASAP7_75t_L g1927 ( 
.A(n_1903),
.B(n_1890),
.Y(n_1927)
);

NAND2xp5_ASAP7_75t_L g1928 ( 
.A(n_1895),
.B(n_1873),
.Y(n_1928)
);

NOR2xp33_ASAP7_75t_L g1929 ( 
.A(n_1912),
.B(n_1889),
.Y(n_1929)
);

AOI211xp5_ASAP7_75t_L g1930 ( 
.A1(n_1917),
.A2(n_1907),
.B(n_1904),
.C(n_1909),
.Y(n_1930)
);

AOI22xp5_ASAP7_75t_L g1931 ( 
.A1(n_1918),
.A2(n_1873),
.B1(n_1875),
.B2(n_1900),
.Y(n_1931)
);

AOI221x1_ASAP7_75t_SL g1932 ( 
.A1(n_1926),
.A2(n_1914),
.B1(n_1906),
.B2(n_1909),
.C(n_1882),
.Y(n_1932)
);

AOI221xp5_ASAP7_75t_L g1933 ( 
.A1(n_1928),
.A2(n_1913),
.B1(n_1888),
.B2(n_1869),
.C(n_1875),
.Y(n_1933)
);

NOR4xp25_ASAP7_75t_L g1934 ( 
.A(n_1923),
.B(n_1910),
.C(n_1901),
.D(n_1809),
.Y(n_1934)
);

AOI21xp5_ASAP7_75t_L g1935 ( 
.A1(n_1925),
.A2(n_1799),
.B(n_1843),
.Y(n_1935)
);

OAI22xp33_ASAP7_75t_L g1936 ( 
.A1(n_1925),
.A2(n_1768),
.B1(n_1774),
.B2(n_1775),
.Y(n_1936)
);

A2O1A1Ixp33_ASAP7_75t_L g1937 ( 
.A1(n_1916),
.A2(n_1883),
.B(n_1918),
.C(n_1927),
.Y(n_1937)
);

NAND4xp25_ASAP7_75t_L g1938 ( 
.A(n_1929),
.B(n_1600),
.C(n_1603),
.D(n_1843),
.Y(n_1938)
);

OAI221xp5_ASAP7_75t_L g1939 ( 
.A1(n_1921),
.A2(n_1920),
.B1(n_1883),
.B2(n_1924),
.C(n_1919),
.Y(n_1939)
);

NAND4xp25_ASAP7_75t_L g1940 ( 
.A(n_1922),
.B(n_1845),
.C(n_1593),
.D(n_1832),
.Y(n_1940)
);

INVxp67_ASAP7_75t_L g1941 ( 
.A(n_1916),
.Y(n_1941)
);

OAI21xp5_ASAP7_75t_L g1942 ( 
.A1(n_1917),
.A2(n_1845),
.B(n_1768),
.Y(n_1942)
);

OR2x2_ASAP7_75t_L g1943 ( 
.A(n_1931),
.B(n_1849),
.Y(n_1943)
);

INVxp67_ASAP7_75t_L g1944 ( 
.A(n_1939),
.Y(n_1944)
);

INVx1_ASAP7_75t_SL g1945 ( 
.A(n_1935),
.Y(n_1945)
);

INVx1_ASAP7_75t_L g1946 ( 
.A(n_1941),
.Y(n_1946)
);

AOI22xp5_ASAP7_75t_L g1947 ( 
.A1(n_1930),
.A2(n_1803),
.B1(n_1801),
.B2(n_1768),
.Y(n_1947)
);

INVx1_ASAP7_75t_L g1948 ( 
.A(n_1940),
.Y(n_1948)
);

OAI22xp33_ASAP7_75t_L g1949 ( 
.A1(n_1942),
.A2(n_1774),
.B1(n_1768),
.B2(n_1856),
.Y(n_1949)
);

INVxp67_ASAP7_75t_L g1950 ( 
.A(n_1943),
.Y(n_1950)
);

AND2x2_ASAP7_75t_L g1951 ( 
.A(n_1946),
.B(n_1937),
.Y(n_1951)
);

INVx2_ASAP7_75t_SL g1952 ( 
.A(n_1948),
.Y(n_1952)
);

INVx1_ASAP7_75t_L g1953 ( 
.A(n_1945),
.Y(n_1953)
);

INVx2_ASAP7_75t_L g1954 ( 
.A(n_1944),
.Y(n_1954)
);

INVxp67_ASAP7_75t_L g1955 ( 
.A(n_1947),
.Y(n_1955)
);

NAND2xp5_ASAP7_75t_L g1956 ( 
.A(n_1949),
.B(n_1932),
.Y(n_1956)
);

NAND2xp5_ASAP7_75t_L g1957 ( 
.A(n_1945),
.B(n_1934),
.Y(n_1957)
);

NAND2xp5_ASAP7_75t_L g1958 ( 
.A(n_1950),
.B(n_1933),
.Y(n_1958)
);

NOR2x1_ASAP7_75t_L g1959 ( 
.A(n_1957),
.B(n_1938),
.Y(n_1959)
);

AOI322xp5_ASAP7_75t_L g1960 ( 
.A1(n_1957),
.A2(n_1936),
.A3(n_1859),
.B1(n_1794),
.B2(n_1804),
.C1(n_1805),
.C2(n_1812),
.Y(n_1960)
);

NAND3xp33_ASAP7_75t_SL g1961 ( 
.A(n_1956),
.B(n_1579),
.C(n_1832),
.Y(n_1961)
);

O2A1O1Ixp33_ASAP7_75t_L g1962 ( 
.A1(n_1955),
.A2(n_1953),
.B(n_1954),
.C(n_1951),
.Y(n_1962)
);

NAND2xp5_ASAP7_75t_L g1963 ( 
.A(n_1952),
.B(n_1836),
.Y(n_1963)
);

INVx4_ASAP7_75t_L g1964 ( 
.A(n_1962),
.Y(n_1964)
);

INVx3_ASAP7_75t_L g1965 ( 
.A(n_1963),
.Y(n_1965)
);

AND2x4_ASAP7_75t_L g1966 ( 
.A(n_1959),
.B(n_1859),
.Y(n_1966)
);

OAI22xp33_ASAP7_75t_L g1967 ( 
.A1(n_1964),
.A2(n_1958),
.B1(n_1961),
.B2(n_1836),
.Y(n_1967)
);

OAI211xp5_ASAP7_75t_L g1968 ( 
.A1(n_1967),
.A2(n_1964),
.B(n_1965),
.C(n_1960),
.Y(n_1968)
);

OAI31xp33_ASAP7_75t_L g1969 ( 
.A1(n_1968),
.A2(n_1966),
.A3(n_1965),
.B(n_1807),
.Y(n_1969)
);

CKINVDCx12_ASAP7_75t_R g1970 ( 
.A(n_1968),
.Y(n_1970)
);

XOR2x2_ASAP7_75t_L g1971 ( 
.A(n_1970),
.B(n_1966),
.Y(n_1971)
);

XNOR2xp5_ASAP7_75t_L g1972 ( 
.A(n_1969),
.B(n_1786),
.Y(n_1972)
);

OAI22xp5_ASAP7_75t_L g1973 ( 
.A1(n_1972),
.A2(n_1827),
.B1(n_1805),
.B2(n_1804),
.Y(n_1973)
);

OAI22xp5_ASAP7_75t_SL g1974 ( 
.A1(n_1971),
.A2(n_1793),
.B1(n_1812),
.B2(n_1827),
.Y(n_1974)
);

XOR2xp5_ASAP7_75t_L g1975 ( 
.A(n_1974),
.B(n_1627),
.Y(n_1975)
);

AOI22xp33_ASAP7_75t_SL g1976 ( 
.A1(n_1975),
.A2(n_1973),
.B1(n_1827),
.B2(n_1811),
.Y(n_1976)
);

AOI22xp5_ASAP7_75t_L g1977 ( 
.A1(n_1976),
.A2(n_1827),
.B1(n_1794),
.B2(n_1804),
.Y(n_1977)
);

AOI322xp5_ASAP7_75t_L g1978 ( 
.A1(n_1977),
.A2(n_1811),
.A3(n_1806),
.B1(n_1805),
.B2(n_1812),
.C1(n_1804),
.C2(n_1824),
.Y(n_1978)
);

OAI22xp5_ASAP7_75t_L g1979 ( 
.A1(n_1978),
.A2(n_1794),
.B1(n_1822),
.B2(n_1812),
.Y(n_1979)
);

AOI211xp5_ASAP7_75t_L g1980 ( 
.A1(n_1979),
.A2(n_1811),
.B(n_1817),
.C(n_1822),
.Y(n_1980)
);


endmodule