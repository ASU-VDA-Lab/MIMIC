module fake_netlist_1_464_n_29 (n_11, n_1, n_2, n_12, n_6, n_4, n_3, n_9, n_5, n_7, n_10, n_8, n_0, n_29);
input n_11;
input n_1;
input n_2;
input n_12;
input n_6;
input n_4;
input n_3;
input n_9;
input n_5;
input n_7;
input n_10;
input n_8;
input n_0;
output n_29;
wire n_20;
wire n_23;
wire n_28;
wire n_22;
wire n_25;
wire n_16;
wire n_26;
wire n_13;
wire n_18;
wire n_17;
wire n_14;
wire n_15;
wire n_24;
wire n_19;
wire n_21;
wire n_27;
INVx2_ASAP7_75t_SL g13 ( .A(n_1), .Y(n_13) );
INVx2_ASAP7_75t_L g14 ( .A(n_3), .Y(n_14) );
INVx1_ASAP7_75t_L g15 ( .A(n_4), .Y(n_15) );
AND2x4_ASAP7_75t_L g16 ( .A(n_6), .B(n_8), .Y(n_16) );
NOR2xp67_ASAP7_75t_L g17 ( .A(n_10), .B(n_12), .Y(n_17) );
HB1xp67_ASAP7_75t_L g18 ( .A(n_11), .Y(n_18) );
INVx2_ASAP7_75t_L g19 ( .A(n_13), .Y(n_19) );
OAI22xp5_ASAP7_75t_L g20 ( .A1(n_14), .A2(n_0), .B1(n_1), .B2(n_2), .Y(n_20) );
INVx2_ASAP7_75t_L g21 ( .A(n_19), .Y(n_21) );
INVx2_ASAP7_75t_L g22 ( .A(n_21), .Y(n_22) );
AOI21xp33_ASAP7_75t_L g23 ( .A1(n_22), .A2(n_20), .B(n_18), .Y(n_23) );
INVxp33_ASAP7_75t_L g24 ( .A(n_23), .Y(n_24) );
INVx1_ASAP7_75t_L g25 ( .A(n_24), .Y(n_25) );
CKINVDCx5p33_ASAP7_75t_R g26 ( .A(n_25), .Y(n_26) );
OAI22xp5_ASAP7_75t_L g27 ( .A1(n_26), .A2(n_18), .B1(n_14), .B2(n_16), .Y(n_27) );
AOI22xp5_ASAP7_75t_L g28 ( .A1(n_27), .A2(n_16), .B1(n_17), .B2(n_15), .Y(n_28) );
AOI322xp5_ASAP7_75t_L g29 ( .A1(n_28), .A2(n_0), .A3(n_2), .B1(n_3), .B2(n_5), .C1(n_7), .C2(n_9), .Y(n_29) );
endmodule