module fake_jpeg_24069_n_333 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_333);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_333;

wire n_253;
wire n_330;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

BUFx3_ASAP7_75t_L g17 ( 
.A(n_3),
.Y(n_17)
);

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_6),
.Y(n_18)
);

NOR2xp33_ASAP7_75t_L g19 ( 
.A(n_15),
.B(n_5),
.Y(n_19)
);

BUFx12f_ASAP7_75t_L g20 ( 
.A(n_6),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_1),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_11),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_10),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_15),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_12),
.Y(n_25)
);

INVx6_ASAP7_75t_L g26 ( 
.A(n_4),
.Y(n_26)
);

BUFx5_ASAP7_75t_L g27 ( 
.A(n_12),
.Y(n_27)
);

BUFx3_ASAP7_75t_L g28 ( 
.A(n_9),
.Y(n_28)
);

INVx4_ASAP7_75t_L g29 ( 
.A(n_14),
.Y(n_29)
);

INVx8_ASAP7_75t_L g30 ( 
.A(n_2),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_0),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_0),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_1),
.Y(n_33)
);

INVx6_ASAP7_75t_L g34 ( 
.A(n_5),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_7),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_3),
.Y(n_36)
);

INVx11_ASAP7_75t_L g37 ( 
.A(n_2),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_8),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_20),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_39),
.Y(n_56)
);

BUFx5_ASAP7_75t_L g40 ( 
.A(n_20),
.Y(n_40)
);

INVx3_ASAP7_75t_SL g59 ( 
.A(n_40),
.Y(n_59)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_21),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_41),
.B(n_43),
.Y(n_54)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_21),
.Y(n_42)
);

NAND2xp5_ASAP7_75t_L g62 ( 
.A(n_42),
.B(n_35),
.Y(n_62)
);

INVx2_ASAP7_75t_L g43 ( 
.A(n_30),
.Y(n_43)
);

BUFx5_ASAP7_75t_L g44 ( 
.A(n_20),
.Y(n_44)
);

INVx1_ASAP7_75t_SL g68 ( 
.A(n_44),
.Y(n_68)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_20),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g80 ( 
.A(n_45),
.Y(n_80)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_20),
.Y(n_46)
);

INVx3_ASAP7_75t_L g58 ( 
.A(n_46),
.Y(n_58)
);

INVx3_ASAP7_75t_L g47 ( 
.A(n_37),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_47),
.B(n_48),
.Y(n_60)
);

INVx2_ASAP7_75t_L g48 ( 
.A(n_30),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_SL g49 ( 
.A(n_19),
.B(n_8),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_49),
.B(n_50),
.Y(n_83)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_32),
.Y(n_50)
);

BUFx12_ASAP7_75t_L g51 ( 
.A(n_20),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_51),
.B(n_17),
.Y(n_85)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_40),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_52),
.B(n_63),
.Y(n_92)
);

INVx2_ASAP7_75t_L g53 ( 
.A(n_51),
.Y(n_53)
);

INVx6_ASAP7_75t_L g109 ( 
.A(n_53),
.Y(n_109)
);

OAI22xp5_ASAP7_75t_L g55 ( 
.A1(n_41),
.A2(n_26),
.B1(n_34),
.B2(n_29),
.Y(n_55)
);

AOI22xp5_ASAP7_75t_L g99 ( 
.A1(n_55),
.A2(n_25),
.B1(n_31),
.B2(n_36),
.Y(n_99)
);

OAI22xp33_ASAP7_75t_L g57 ( 
.A1(n_40),
.A2(n_30),
.B1(n_29),
.B2(n_37),
.Y(n_57)
);

OAI22xp5_ASAP7_75t_SL g98 ( 
.A1(n_57),
.A2(n_67),
.B1(n_31),
.B2(n_23),
.Y(n_98)
);

BUFx3_ASAP7_75t_L g61 ( 
.A(n_44),
.Y(n_61)
);

INVx5_ASAP7_75t_L g108 ( 
.A(n_61),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_L g91 ( 
.A(n_62),
.B(n_74),
.Y(n_91)
);

INVx3_ASAP7_75t_L g63 ( 
.A(n_44),
.Y(n_63)
);

AOI22xp33_ASAP7_75t_SL g64 ( 
.A1(n_47),
.A2(n_26),
.B1(n_34),
.B2(n_29),
.Y(n_64)
);

AOI22xp33_ASAP7_75t_SL g105 ( 
.A1(n_64),
.A2(n_78),
.B1(n_79),
.B2(n_25),
.Y(n_105)
);

INVx2_ASAP7_75t_L g65 ( 
.A(n_51),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g114 ( 
.A(n_65),
.B(n_69),
.Y(n_114)
);

AOI22xp5_ASAP7_75t_SL g66 ( 
.A1(n_42),
.A2(n_26),
.B1(n_34),
.B2(n_30),
.Y(n_66)
);

A2O1A1Ixp33_ASAP7_75t_L g95 ( 
.A1(n_66),
.A2(n_82),
.B(n_18),
.C(n_38),
.Y(n_95)
);

AOI22xp5_ASAP7_75t_L g67 ( 
.A1(n_47),
.A2(n_26),
.B1(n_37),
.B2(n_28),
.Y(n_67)
);

INVx2_ASAP7_75t_L g69 ( 
.A(n_51),
.Y(n_69)
);

AND2x2_ASAP7_75t_SL g70 ( 
.A(n_51),
.B(n_27),
.Y(n_70)
);

AND2x2_ASAP7_75t_L g103 ( 
.A(n_70),
.B(n_14),
.Y(n_103)
);

INVx2_ASAP7_75t_L g71 ( 
.A(n_43),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g121 ( 
.A(n_71),
.B(n_72),
.Y(n_121)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_50),
.Y(n_72)
);

INVx2_ASAP7_75t_L g73 ( 
.A(n_43),
.Y(n_73)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_73),
.Y(n_89)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_39),
.Y(n_74)
);

INVx3_ASAP7_75t_L g75 ( 
.A(n_48),
.Y(n_75)
);

INVx4_ASAP7_75t_SL g117 ( 
.A(n_75),
.Y(n_117)
);

BUFx12f_ASAP7_75t_L g76 ( 
.A(n_39),
.Y(n_76)
);

INVx1_ASAP7_75t_SL g88 ( 
.A(n_76),
.Y(n_88)
);

INVx3_ASAP7_75t_L g77 ( 
.A(n_48),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_L g97 ( 
.A(n_77),
.B(n_81),
.Y(n_97)
);

AOI22xp33_ASAP7_75t_SL g78 ( 
.A1(n_42),
.A2(n_27),
.B1(n_23),
.B2(n_35),
.Y(n_78)
);

AOI22xp33_ASAP7_75t_SL g79 ( 
.A1(n_49),
.A2(n_27),
.B1(n_23),
.B2(n_35),
.Y(n_79)
);

INVx3_ASAP7_75t_L g81 ( 
.A(n_39),
.Y(n_81)
);

OAI21xp33_ASAP7_75t_L g82 ( 
.A1(n_45),
.A2(n_17),
.B(n_28),
.Y(n_82)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_45),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g116 ( 
.A(n_84),
.B(n_38),
.Y(n_116)
);

CKINVDCx16_ASAP7_75t_R g96 ( 
.A(n_85),
.Y(n_96)
);

INVx3_ASAP7_75t_L g86 ( 
.A(n_76),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g136 ( 
.A(n_86),
.B(n_94),
.Y(n_136)
);

BUFx12f_ASAP7_75t_L g87 ( 
.A(n_61),
.Y(n_87)
);

BUFx3_ASAP7_75t_L g132 ( 
.A(n_87),
.Y(n_132)
);

INVx2_ASAP7_75t_L g90 ( 
.A(n_76),
.Y(n_90)
);

INVx6_ASAP7_75t_L g128 ( 
.A(n_90),
.Y(n_128)
);

AOI22xp5_ASAP7_75t_SL g93 ( 
.A1(n_66),
.A2(n_28),
.B1(n_17),
.B2(n_19),
.Y(n_93)
);

INVxp67_ASAP7_75t_L g123 ( 
.A(n_93),
.Y(n_123)
);

INVx3_ASAP7_75t_L g94 ( 
.A(n_75),
.Y(n_94)
);

OAI22xp5_ASAP7_75t_L g133 ( 
.A1(n_95),
.A2(n_99),
.B1(n_105),
.B2(n_32),
.Y(n_133)
);

AOI22xp5_ASAP7_75t_L g148 ( 
.A1(n_98),
.A2(n_104),
.B1(n_113),
.B2(n_18),
.Y(n_148)
);

INVx2_ASAP7_75t_L g100 ( 
.A(n_77),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g149 ( 
.A(n_100),
.B(n_110),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_L g101 ( 
.A(n_62),
.B(n_46),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_L g140 ( 
.A(n_101),
.B(n_102),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_L g102 ( 
.A(n_54),
.B(n_46),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_L g141 ( 
.A(n_103),
.B(n_120),
.Y(n_141)
);

OAI22xp5_ASAP7_75t_SL g104 ( 
.A1(n_67),
.A2(n_31),
.B1(n_25),
.B2(n_33),
.Y(n_104)
);

A2O1A1Ixp33_ASAP7_75t_L g106 ( 
.A1(n_83),
.A2(n_22),
.B(n_36),
.C(n_24),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_SL g125 ( 
.A(n_106),
.B(n_107),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_SL g107 ( 
.A(n_63),
.B(n_22),
.Y(n_107)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_60),
.Y(n_110)
);

AND2x4_ASAP7_75t_SL g111 ( 
.A(n_70),
.B(n_46),
.Y(n_111)
);

AOI21xp33_ASAP7_75t_L g135 ( 
.A1(n_111),
.A2(n_0),
.B(n_1),
.Y(n_135)
);

BUFx3_ASAP7_75t_L g112 ( 
.A(n_68),
.Y(n_112)
);

BUFx3_ASAP7_75t_L g145 ( 
.A(n_112),
.Y(n_145)
);

O2A1O1Ixp33_ASAP7_75t_SL g113 ( 
.A1(n_70),
.A2(n_38),
.B(n_18),
.C(n_45),
.Y(n_113)
);

INVx4_ASAP7_75t_L g115 ( 
.A(n_68),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_L g153 ( 
.A(n_115),
.B(n_118),
.Y(n_153)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_116),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_SL g118 ( 
.A(n_58),
.B(n_24),
.Y(n_118)
);

BUFx6f_ASAP7_75t_L g119 ( 
.A(n_56),
.Y(n_119)
);

CKINVDCx16_ASAP7_75t_R g134 ( 
.A(n_119),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_L g120 ( 
.A(n_58),
.B(n_38),
.Y(n_120)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_71),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_L g156 ( 
.A(n_122),
.B(n_8),
.Y(n_156)
);

CKINVDCx14_ASAP7_75t_R g126 ( 
.A(n_114),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_L g164 ( 
.A(n_126),
.B(n_130),
.Y(n_164)
);

CKINVDCx5p33_ASAP7_75t_R g127 ( 
.A(n_112),
.Y(n_127)
);

CKINVDCx16_ASAP7_75t_R g187 ( 
.A(n_127),
.Y(n_187)
);

MAJIxp5_ASAP7_75t_L g129 ( 
.A(n_111),
.B(n_101),
.C(n_102),
.Y(n_129)
);

MAJIxp5_ASAP7_75t_L g177 ( 
.A(n_129),
.B(n_147),
.C(n_154),
.Y(n_177)
);

INVx3_ASAP7_75t_SL g130 ( 
.A(n_87),
.Y(n_130)
);

OAI22xp5_ASAP7_75t_SL g131 ( 
.A1(n_95),
.A2(n_93),
.B1(n_111),
.B2(n_99),
.Y(n_131)
);

AOI22xp5_ASAP7_75t_L g169 ( 
.A1(n_131),
.A2(n_133),
.B1(n_137),
.B2(n_143),
.Y(n_169)
);

OAI21xp5_ASAP7_75t_SL g178 ( 
.A1(n_135),
.A2(n_10),
.B(n_3),
.Y(n_178)
);

OAI22xp5_ASAP7_75t_SL g137 ( 
.A1(n_98),
.A2(n_73),
.B1(n_57),
.B2(n_81),
.Y(n_137)
);

INVxp67_ASAP7_75t_L g138 ( 
.A(n_92),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_L g171 ( 
.A(n_138),
.B(n_142),
.Y(n_171)
);

AOI32xp33_ASAP7_75t_L g139 ( 
.A1(n_113),
.A2(n_82),
.A3(n_59),
.B1(n_69),
.B2(n_65),
.Y(n_139)
);

MAJIxp5_ASAP7_75t_SL g170 ( 
.A(n_139),
.B(n_108),
.C(n_88),
.Y(n_170)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_97),
.Y(n_142)
);

OAI22xp5_ASAP7_75t_SL g143 ( 
.A1(n_120),
.A2(n_53),
.B1(n_33),
.B2(n_18),
.Y(n_143)
);

HB1xp67_ASAP7_75t_L g144 ( 
.A(n_87),
.Y(n_144)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_144),
.Y(n_174)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_121),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_L g172 ( 
.A(n_146),
.B(n_152),
.Y(n_172)
);

XOR2xp5_ASAP7_75t_L g147 ( 
.A(n_91),
.B(n_59),
.Y(n_147)
);

OAI22xp33_ASAP7_75t_SL g159 ( 
.A1(n_148),
.A2(n_117),
.B1(n_100),
.B2(n_109),
.Y(n_159)
);

OAI22xp5_ASAP7_75t_L g150 ( 
.A1(n_106),
.A2(n_9),
.B1(n_16),
.B2(n_15),
.Y(n_150)
);

AOI22xp5_ASAP7_75t_L g179 ( 
.A1(n_150),
.A2(n_11),
.B1(n_4),
.B2(n_5),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_L g151 ( 
.A(n_103),
.B(n_80),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_L g168 ( 
.A(n_151),
.B(n_155),
.Y(n_168)
);

INVx2_ASAP7_75t_L g152 ( 
.A(n_94),
.Y(n_152)
);

MAJIxp5_ASAP7_75t_L g154 ( 
.A(n_96),
.B(n_80),
.C(n_56),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_L g155 ( 
.A(n_103),
.B(n_0),
.Y(n_155)
);

CKINVDCx16_ASAP7_75t_R g188 ( 
.A(n_156),
.Y(n_188)
);

CKINVDCx20_ASAP7_75t_R g157 ( 
.A(n_104),
.Y(n_157)
);

NOR2xp33_ASAP7_75t_L g186 ( 
.A(n_157),
.B(n_158),
.Y(n_186)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_115),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_SL g203 ( 
.A(n_159),
.B(n_162),
.Y(n_203)
);

NOR2xp33_ASAP7_75t_SL g160 ( 
.A(n_125),
.B(n_13),
.Y(n_160)
);

NOR2xp33_ASAP7_75t_SL g208 ( 
.A(n_160),
.B(n_166),
.Y(n_208)
);

AOI32xp33_ASAP7_75t_L g161 ( 
.A1(n_123),
.A2(n_86),
.A3(n_109),
.B1(n_108),
.B2(n_117),
.Y(n_161)
);

XOR2xp5_ASAP7_75t_L g204 ( 
.A(n_161),
.B(n_127),
.Y(n_204)
);

INVxp67_ASAP7_75t_L g162 ( 
.A(n_136),
.Y(n_162)
);

CKINVDCx20_ASAP7_75t_R g163 ( 
.A(n_149),
.Y(n_163)
);

CKINVDCx20_ASAP7_75t_R g211 ( 
.A(n_163),
.Y(n_211)
);

AND2x2_ASAP7_75t_L g165 ( 
.A(n_151),
.B(n_1),
.Y(n_165)
);

OAI21xp5_ASAP7_75t_SL g201 ( 
.A1(n_165),
.A2(n_167),
.B(n_170),
.Y(n_201)
);

NOR2xp33_ASAP7_75t_SL g166 ( 
.A(n_125),
.B(n_12),
.Y(n_166)
);

OAI21xp5_ASAP7_75t_L g167 ( 
.A1(n_141),
.A2(n_89),
.B(n_88),
.Y(n_167)
);

NOR2xp33_ASAP7_75t_SL g173 ( 
.A(n_141),
.B(n_10),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_SL g206 ( 
.A(n_173),
.B(n_179),
.Y(n_206)
);

INVx2_ASAP7_75t_L g175 ( 
.A(n_145),
.Y(n_175)
);

NOR2xp33_ASAP7_75t_L g210 ( 
.A(n_175),
.B(n_176),
.Y(n_210)
);

INVx3_ASAP7_75t_L g176 ( 
.A(n_145),
.Y(n_176)
);

OAI21xp5_ASAP7_75t_SL g212 ( 
.A1(n_178),
.A2(n_190),
.B(n_191),
.Y(n_212)
);

OAI22xp33_ASAP7_75t_SL g180 ( 
.A1(n_157),
.A2(n_137),
.B1(n_139),
.B2(n_148),
.Y(n_180)
);

INVxp67_ASAP7_75t_L g198 ( 
.A(n_180),
.Y(n_198)
);

OAI22xp5_ASAP7_75t_SL g181 ( 
.A1(n_123),
.A2(n_90),
.B1(n_119),
.B2(n_2),
.Y(n_181)
);

OAI22xp5_ASAP7_75t_SL g209 ( 
.A1(n_181),
.A2(n_182),
.B1(n_134),
.B2(n_128),
.Y(n_209)
);

AOI22xp5_ASAP7_75t_L g182 ( 
.A1(n_131),
.A2(n_2),
.B1(n_4),
.B2(n_6),
.Y(n_182)
);

MAJIxp5_ASAP7_75t_L g183 ( 
.A(n_129),
.B(n_7),
.C(n_9),
.Y(n_183)
);

MAJIxp5_ASAP7_75t_L g193 ( 
.A(n_183),
.B(n_184),
.C(n_185),
.Y(n_193)
);

XOR2xp5_ASAP7_75t_L g184 ( 
.A(n_147),
.B(n_16),
.Y(n_184)
);

MAJIxp5_ASAP7_75t_L g185 ( 
.A(n_140),
.B(n_7),
.C(n_11),
.Y(n_185)
);

MAJIxp5_ASAP7_75t_L g189 ( 
.A(n_140),
.B(n_13),
.C(n_14),
.Y(n_189)
);

MAJIxp5_ASAP7_75t_L g195 ( 
.A(n_189),
.B(n_124),
.C(n_143),
.Y(n_195)
);

OAI21xp5_ASAP7_75t_L g190 ( 
.A1(n_155),
.A2(n_13),
.B(n_16),
.Y(n_190)
);

AOI21xp5_ASAP7_75t_L g191 ( 
.A1(n_142),
.A2(n_124),
.B(n_154),
.Y(n_191)
);

INVxp67_ASAP7_75t_L g192 ( 
.A(n_132),
.Y(n_192)
);

INVxp67_ASAP7_75t_L g217 ( 
.A(n_192),
.Y(n_217)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_172),
.Y(n_194)
);

NOR2xp33_ASAP7_75t_L g248 ( 
.A(n_194),
.B(n_202),
.Y(n_248)
);

MAJIxp5_ASAP7_75t_L g229 ( 
.A(n_195),
.B(n_199),
.C(n_188),
.Y(n_229)
);

NAND2xp5_ASAP7_75t_L g196 ( 
.A(n_168),
.B(n_153),
.Y(n_196)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_196),
.Y(n_230)
);

AND2x2_ASAP7_75t_L g197 ( 
.A(n_170),
.B(n_132),
.Y(n_197)
);

OAI21xp5_ASAP7_75t_SL g238 ( 
.A1(n_197),
.A2(n_200),
.B(n_218),
.Y(n_238)
);

MAJIxp5_ASAP7_75t_L g199 ( 
.A(n_177),
.B(n_146),
.C(n_158),
.Y(n_199)
);

AOI21xp5_ASAP7_75t_L g200 ( 
.A1(n_186),
.A2(n_152),
.B(n_138),
.Y(n_200)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_171),
.Y(n_202)
);

XOR2xp5_ASAP7_75t_L g240 ( 
.A(n_204),
.B(n_215),
.Y(n_240)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_164),
.Y(n_205)
);

AOI22xp33_ASAP7_75t_L g226 ( 
.A1(n_205),
.A2(n_209),
.B1(n_216),
.B2(n_197),
.Y(n_226)
);

INVx3_ASAP7_75t_L g207 ( 
.A(n_176),
.Y(n_207)
);

INVx3_ASAP7_75t_L g228 ( 
.A(n_207),
.Y(n_228)
);

OAI32xp33_ASAP7_75t_L g213 ( 
.A1(n_169),
.A2(n_128),
.A3(n_130),
.B1(n_168),
.B2(n_182),
.Y(n_213)
);

NAND2xp5_ASAP7_75t_L g224 ( 
.A(n_213),
.B(n_216),
.Y(n_224)
);

NAND2xp5_ASAP7_75t_L g214 ( 
.A(n_184),
.B(n_130),
.Y(n_214)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_214),
.Y(n_231)
);

XNOR2xp5_ASAP7_75t_L g215 ( 
.A(n_177),
.B(n_167),
.Y(n_215)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_181),
.Y(n_216)
);

AOI21xp5_ASAP7_75t_L g218 ( 
.A1(n_161),
.A2(n_178),
.B(n_191),
.Y(n_218)
);

OAI22xp5_ASAP7_75t_SL g219 ( 
.A1(n_169),
.A2(n_179),
.B1(n_165),
.B2(n_183),
.Y(n_219)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_219),
.Y(n_233)
);

OAI22xp5_ASAP7_75t_SL g220 ( 
.A1(n_165),
.A2(n_162),
.B1(n_163),
.B2(n_187),
.Y(n_220)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_220),
.Y(n_235)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_173),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_L g227 ( 
.A(n_221),
.B(n_160),
.Y(n_227)
);

AOI21xp5_ASAP7_75t_L g222 ( 
.A1(n_187),
.A2(n_174),
.B(n_190),
.Y(n_222)
);

AOI21xp5_ASAP7_75t_L g241 ( 
.A1(n_222),
.A2(n_201),
.B(n_212),
.Y(n_241)
);

NAND2xp5_ASAP7_75t_L g223 ( 
.A(n_185),
.B(n_189),
.Y(n_223)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_223),
.Y(n_239)
);

AOI22xp5_ASAP7_75t_SL g225 ( 
.A1(n_198),
.A2(n_188),
.B1(n_174),
.B2(n_192),
.Y(n_225)
);

OAI22xp5_ASAP7_75t_SL g264 ( 
.A1(n_225),
.A2(n_208),
.B1(n_217),
.B2(n_224),
.Y(n_264)
);

INVxp67_ASAP7_75t_L g252 ( 
.A(n_226),
.Y(n_252)
);

NAND2xp5_ASAP7_75t_L g251 ( 
.A(n_227),
.B(n_246),
.Y(n_251)
);

MAJIxp5_ASAP7_75t_L g260 ( 
.A(n_229),
.B(n_237),
.C(n_223),
.Y(n_260)
);

NAND2xp5_ASAP7_75t_L g232 ( 
.A(n_196),
.B(n_166),
.Y(n_232)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_232),
.Y(n_249)
);

NAND2xp5_ASAP7_75t_L g234 ( 
.A(n_214),
.B(n_213),
.Y(n_234)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_234),
.Y(n_263)
);

OAI21xp5_ASAP7_75t_L g236 ( 
.A1(n_218),
.A2(n_175),
.B(n_222),
.Y(n_236)
);

AOI21xp5_ASAP7_75t_L g258 ( 
.A1(n_236),
.A2(n_241),
.B(n_244),
.Y(n_258)
);

MAJIxp5_ASAP7_75t_L g237 ( 
.A(n_199),
.B(n_215),
.C(n_201),
.Y(n_237)
);

XOR2xp5_ASAP7_75t_L g242 ( 
.A(n_204),
.B(n_193),
.Y(n_242)
);

XOR2xp5_ASAP7_75t_L g257 ( 
.A(n_242),
.B(n_247),
.Y(n_257)
);

NAND2xp5_ASAP7_75t_L g243 ( 
.A(n_220),
.B(n_219),
.Y(n_243)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_243),
.Y(n_266)
);

OAI21xp5_ASAP7_75t_L g244 ( 
.A1(n_198),
.A2(n_197),
.B(n_203),
.Y(n_244)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_210),
.Y(n_245)
);

NOR2xp33_ASAP7_75t_L g262 ( 
.A(n_245),
.B(n_200),
.Y(n_262)
);

NAND2xp5_ASAP7_75t_L g246 ( 
.A(n_212),
.B(n_221),
.Y(n_246)
);

XOR2xp5_ASAP7_75t_L g247 ( 
.A(n_193),
.B(n_195),
.Y(n_247)
);

INVx3_ASAP7_75t_SL g250 ( 
.A(n_228),
.Y(n_250)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_250),
.Y(n_284)
);

OAI22xp5_ASAP7_75t_L g253 ( 
.A1(n_224),
.A2(n_235),
.B1(n_234),
.B2(n_233),
.Y(n_253)
);

AOI22xp5_ASAP7_75t_L g272 ( 
.A1(n_253),
.A2(n_264),
.B1(n_244),
.B2(n_238),
.Y(n_272)
);

CKINVDCx20_ASAP7_75t_R g254 ( 
.A(n_248),
.Y(n_254)
);

CKINVDCx20_ASAP7_75t_R g283 ( 
.A(n_254),
.Y(n_283)
);

NAND2xp5_ASAP7_75t_L g255 ( 
.A(n_230),
.B(n_206),
.Y(n_255)
);

NAND2xp5_ASAP7_75t_L g281 ( 
.A(n_255),
.B(n_256),
.Y(n_281)
);

NAND2xp5_ASAP7_75t_L g256 ( 
.A(n_230),
.B(n_194),
.Y(n_256)
);

AOI22xp5_ASAP7_75t_L g259 ( 
.A1(n_233),
.A2(n_209),
.B1(n_207),
.B2(n_217),
.Y(n_259)
);

OAI22xp5_ASAP7_75t_SL g277 ( 
.A1(n_259),
.A2(n_248),
.B1(n_240),
.B2(n_242),
.Y(n_277)
);

MAJIxp5_ASAP7_75t_L g275 ( 
.A(n_260),
.B(n_257),
.C(n_237),
.Y(n_275)
);

NAND2xp5_ASAP7_75t_L g261 ( 
.A(n_232),
.B(n_211),
.Y(n_261)
);

NOR2xp33_ASAP7_75t_L g274 ( 
.A(n_261),
.B(n_265),
.Y(n_274)
);

NAND2xp5_ASAP7_75t_SL g273 ( 
.A(n_262),
.B(n_267),
.Y(n_273)
);

NAND2xp5_ASAP7_75t_L g265 ( 
.A(n_239),
.B(n_231),
.Y(n_265)
);

NAND2xp5_ASAP7_75t_L g267 ( 
.A(n_239),
.B(n_231),
.Y(n_267)
);

NAND2xp5_ASAP7_75t_L g268 ( 
.A(n_246),
.B(n_227),
.Y(n_268)
);

NAND2xp5_ASAP7_75t_SL g279 ( 
.A(n_268),
.B(n_249),
.Y(n_279)
);

OAI22xp5_ASAP7_75t_L g269 ( 
.A1(n_259),
.A2(n_225),
.B1(n_235),
.B2(n_243),
.Y(n_269)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_269),
.Y(n_287)
);

AND2x2_ASAP7_75t_L g270 ( 
.A(n_251),
.B(n_240),
.Y(n_270)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_270),
.Y(n_288)
);

OAI22xp5_ASAP7_75t_L g271 ( 
.A1(n_259),
.A2(n_238),
.B1(n_241),
.B2(n_236),
.Y(n_271)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_271),
.Y(n_297)
);

NAND2xp5_ASAP7_75t_L g300 ( 
.A(n_272),
.B(n_285),
.Y(n_300)
);

MAJIxp5_ASAP7_75t_L g290 ( 
.A(n_275),
.B(n_282),
.C(n_260),
.Y(n_290)
);

AOI22xp5_ASAP7_75t_L g276 ( 
.A1(n_266),
.A2(n_245),
.B1(n_229),
.B2(n_228),
.Y(n_276)
);

AOI22xp5_ASAP7_75t_L g291 ( 
.A1(n_276),
.A2(n_277),
.B1(n_278),
.B2(n_286),
.Y(n_291)
);

OAI22xp5_ASAP7_75t_L g278 ( 
.A1(n_252),
.A2(n_247),
.B1(n_266),
.B2(n_263),
.Y(n_278)
);

NAND2xp5_ASAP7_75t_L g293 ( 
.A(n_279),
.B(n_255),
.Y(n_293)
);

NOR2xp33_ASAP7_75t_SL g280 ( 
.A(n_254),
.B(n_261),
.Y(n_280)
);

NAND2xp5_ASAP7_75t_SL g292 ( 
.A(n_280),
.B(n_249),
.Y(n_292)
);

MAJIxp5_ASAP7_75t_L g282 ( 
.A(n_257),
.B(n_260),
.C(n_267),
.Y(n_282)
);

AOI22xp5_ASAP7_75t_SL g285 ( 
.A1(n_251),
.A2(n_268),
.B1(n_262),
.B2(n_263),
.Y(n_285)
);

XOR2xp5_ASAP7_75t_L g294 ( 
.A(n_285),
.B(n_264),
.Y(n_294)
);

AOI21xp5_ASAP7_75t_L g286 ( 
.A1(n_258),
.A2(n_265),
.B(n_256),
.Y(n_286)
);

MAJx2_ASAP7_75t_L g289 ( 
.A(n_270),
.B(n_257),
.C(n_258),
.Y(n_289)
);

XOR2xp5_ASAP7_75t_L g302 ( 
.A(n_289),
.B(n_294),
.Y(n_302)
);

MAJIxp5_ASAP7_75t_L g306 ( 
.A(n_290),
.B(n_298),
.C(n_299),
.Y(n_306)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_292),
.Y(n_303)
);

NOR2xp33_ASAP7_75t_L g304 ( 
.A(n_293),
.B(n_295),
.Y(n_304)
);

NAND2xp5_ASAP7_75t_SL g295 ( 
.A(n_274),
.B(n_283),
.Y(n_295)
);

AO21x1_ASAP7_75t_L g296 ( 
.A1(n_283),
.A2(n_253),
.B(n_250),
.Y(n_296)
);

OAI22xp5_ASAP7_75t_SL g301 ( 
.A1(n_296),
.A2(n_300),
.B1(n_286),
.B2(n_272),
.Y(n_301)
);

MAJIxp5_ASAP7_75t_L g298 ( 
.A(n_282),
.B(n_250),
.C(n_275),
.Y(n_298)
);

MAJIxp5_ASAP7_75t_L g299 ( 
.A(n_276),
.B(n_250),
.C(n_277),
.Y(n_299)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_301),
.Y(n_312)
);

XNOR2xp5_ASAP7_75t_L g305 ( 
.A(n_299),
.B(n_273),
.Y(n_305)
);

XOR2xp5_ASAP7_75t_L g315 ( 
.A(n_305),
.B(n_298),
.Y(n_315)
);

AOI22xp5_ASAP7_75t_L g307 ( 
.A1(n_297),
.A2(n_284),
.B1(n_281),
.B2(n_270),
.Y(n_307)
);

NAND2xp5_ASAP7_75t_L g311 ( 
.A(n_307),
.B(n_308),
.Y(n_311)
);

NOR2xp33_ASAP7_75t_L g308 ( 
.A(n_293),
.B(n_284),
.Y(n_308)
);

INVx11_ASAP7_75t_L g309 ( 
.A(n_296),
.Y(n_309)
);

NAND2xp5_ASAP7_75t_L g316 ( 
.A(n_309),
.B(n_310),
.Y(n_316)
);

BUFx24_ASAP7_75t_SL g310 ( 
.A(n_294),
.Y(n_310)
);

NOR2xp67_ASAP7_75t_L g313 ( 
.A(n_302),
.B(n_288),
.Y(n_313)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_313),
.Y(n_319)
);

INVx6_ASAP7_75t_L g314 ( 
.A(n_306),
.Y(n_314)
);

NOR2xp33_ASAP7_75t_L g322 ( 
.A(n_314),
.B(n_309),
.Y(n_322)
);

MAJIxp5_ASAP7_75t_L g323 ( 
.A(n_315),
.B(n_317),
.C(n_302),
.Y(n_323)
);

MAJIxp5_ASAP7_75t_L g317 ( 
.A(n_306),
.B(n_290),
.C(n_291),
.Y(n_317)
);

XNOR2xp5_ASAP7_75t_L g318 ( 
.A(n_305),
.B(n_291),
.Y(n_318)
);

XNOR2xp5_ASAP7_75t_L g320 ( 
.A(n_318),
.B(n_304),
.Y(n_320)
);

NAND2xp5_ASAP7_75t_SL g325 ( 
.A(n_320),
.B(n_321),
.Y(n_325)
);

NAND2xp5_ASAP7_75t_L g321 ( 
.A(n_311),
.B(n_303),
.Y(n_321)
);

AOI21xp5_ASAP7_75t_SL g324 ( 
.A1(n_322),
.A2(n_312),
.B(n_281),
.Y(n_324)
);

NOR2xp33_ASAP7_75t_L g326 ( 
.A(n_323),
.B(n_315),
.Y(n_326)
);

NOR2xp33_ASAP7_75t_L g327 ( 
.A(n_324),
.B(n_326),
.Y(n_327)
);

AOI21x1_ASAP7_75t_L g328 ( 
.A1(n_325),
.A2(n_322),
.B(n_318),
.Y(n_328)
);

INVxp67_ASAP7_75t_L g329 ( 
.A(n_328),
.Y(n_329)
);

OAI22xp5_ASAP7_75t_SL g330 ( 
.A1(n_329),
.A2(n_327),
.B1(n_319),
.B2(n_314),
.Y(n_330)
);

AOI22xp5_ASAP7_75t_L g331 ( 
.A1(n_330),
.A2(n_317),
.B1(n_287),
.B2(n_316),
.Y(n_331)
);

INVxp67_ASAP7_75t_L g332 ( 
.A(n_331),
.Y(n_332)
);

XNOR2xp5_ASAP7_75t_L g333 ( 
.A(n_332),
.B(n_289),
.Y(n_333)
);


endmodule