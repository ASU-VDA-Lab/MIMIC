module fake_jpeg_28909_n_435 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_435);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_435;

wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_385;
wire n_228;
wire n_134;
wire n_428;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_377;
wire n_291;
wire n_236;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_17;
wire n_431;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_415;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_429;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_305;
wire n_161;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_382;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_389;
wire n_339;
wire n_109;
wire n_267;
wire n_384;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_433;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_413;
wire n_275;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_379;
wire n_114;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_202;
wire n_430;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_409;
wire n_249;
wire n_412;
wire n_217;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_391;
wire n_209;
wire n_22;
wire n_138;
wire n_402;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVx8_ASAP7_75t_L g16 ( 
.A(n_15),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_2),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_0),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_9),
.Y(n_19)
);

BUFx4f_ASAP7_75t_SL g20 ( 
.A(n_2),
.Y(n_20)
);

BUFx4f_ASAP7_75t_SL g21 ( 
.A(n_12),
.Y(n_21)
);

INVxp67_ASAP7_75t_L g22 ( 
.A(n_14),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_8),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_6),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_4),
.Y(n_25)
);

BUFx12f_ASAP7_75t_L g26 ( 
.A(n_11),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_10),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_1),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_12),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_13),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_6),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_14),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_3),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_14),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_12),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_12),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_1),
.Y(n_37)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_4),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_5),
.Y(n_39)
);

BUFx3_ASAP7_75t_L g40 ( 
.A(n_14),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_15),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_15),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_3),
.Y(n_43)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_0),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_1),
.Y(n_45)
);

INVx2_ASAP7_75t_L g46 ( 
.A(n_27),
.Y(n_46)
);

INVx2_ASAP7_75t_L g92 ( 
.A(n_46),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g47 ( 
.A(n_22),
.B(n_7),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g123 ( 
.A(n_47),
.B(n_53),
.Y(n_123)
);

BUFx5_ASAP7_75t_L g48 ( 
.A(n_26),
.Y(n_48)
);

INVx3_ASAP7_75t_SL g126 ( 
.A(n_48),
.Y(n_126)
);

BUFx3_ASAP7_75t_L g49 ( 
.A(n_40),
.Y(n_49)
);

INVx4_ASAP7_75t_L g96 ( 
.A(n_49),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_SL g50 ( 
.A(n_17),
.B(n_7),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_SL g104 ( 
.A(n_50),
.B(n_91),
.Y(n_104)
);

INVx2_ASAP7_75t_L g51 ( 
.A(n_27),
.Y(n_51)
);

INVx2_ASAP7_75t_L g94 ( 
.A(n_51),
.Y(n_94)
);

HAxp5_ASAP7_75t_SL g52 ( 
.A(n_18),
.B(n_7),
.CON(n_52),
.SN(n_52)
);

A2O1A1Ixp33_ASAP7_75t_L g119 ( 
.A1(n_52),
.A2(n_38),
.B(n_34),
.C(n_32),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_17),
.B(n_7),
.Y(n_53)
);

INVx13_ASAP7_75t_L g54 ( 
.A(n_16),
.Y(n_54)
);

BUFx12f_ASAP7_75t_L g111 ( 
.A(n_54),
.Y(n_111)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_27),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g101 ( 
.A(n_55),
.Y(n_101)
);

INVx3_ASAP7_75t_L g56 ( 
.A(n_40),
.Y(n_56)
);

INVx3_ASAP7_75t_L g127 ( 
.A(n_56),
.Y(n_127)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_27),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g112 ( 
.A(n_57),
.Y(n_112)
);

BUFx12f_ASAP7_75t_L g58 ( 
.A(n_31),
.Y(n_58)
);

INVx3_ASAP7_75t_L g128 ( 
.A(n_58),
.Y(n_128)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_31),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g124 ( 
.A(n_59),
.Y(n_124)
);

BUFx5_ASAP7_75t_L g60 ( 
.A(n_26),
.Y(n_60)
);

INVx5_ASAP7_75t_L g93 ( 
.A(n_60),
.Y(n_93)
);

AND2x2_ASAP7_75t_L g61 ( 
.A(n_19),
.B(n_6),
.Y(n_61)
);

MAJIxp5_ASAP7_75t_L g134 ( 
.A(n_61),
.B(n_44),
.C(n_18),
.Y(n_134)
);

BUFx5_ASAP7_75t_L g62 ( 
.A(n_26),
.Y(n_62)
);

INVx5_ASAP7_75t_L g135 ( 
.A(n_62),
.Y(n_135)
);

INVx6_ASAP7_75t_L g63 ( 
.A(n_31),
.Y(n_63)
);

INVx6_ASAP7_75t_L g100 ( 
.A(n_63),
.Y(n_100)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_31),
.Y(n_64)
);

INVx6_ASAP7_75t_L g120 ( 
.A(n_64),
.Y(n_120)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_19),
.Y(n_65)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_65),
.Y(n_99)
);

BUFx3_ASAP7_75t_L g66 ( 
.A(n_40),
.Y(n_66)
);

INVx4_ASAP7_75t_L g117 ( 
.A(n_66),
.Y(n_117)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_33),
.Y(n_67)
);

INVx8_ASAP7_75t_L g143 ( 
.A(n_67),
.Y(n_143)
);

INVx3_ASAP7_75t_L g68 ( 
.A(n_26),
.Y(n_68)
);

INVx3_ASAP7_75t_L g133 ( 
.A(n_68),
.Y(n_133)
);

INVx2_ASAP7_75t_L g69 ( 
.A(n_33),
.Y(n_69)
);

INVx2_ASAP7_75t_L g95 ( 
.A(n_69),
.Y(n_95)
);

BUFx6f_ASAP7_75t_L g70 ( 
.A(n_33),
.Y(n_70)
);

BUFx2_ASAP7_75t_L g114 ( 
.A(n_70),
.Y(n_114)
);

INVx6_ASAP7_75t_L g71 ( 
.A(n_33),
.Y(n_71)
);

BUFx2_ASAP7_75t_L g115 ( 
.A(n_71),
.Y(n_115)
);

INVx6_ASAP7_75t_L g72 ( 
.A(n_45),
.Y(n_72)
);

BUFx2_ASAP7_75t_L g122 ( 
.A(n_72),
.Y(n_122)
);

INVx3_ASAP7_75t_SL g73 ( 
.A(n_45),
.Y(n_73)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_73),
.Y(n_102)
);

INVx8_ASAP7_75t_L g74 ( 
.A(n_16),
.Y(n_74)
);

INVx3_ASAP7_75t_L g141 ( 
.A(n_74),
.Y(n_141)
);

BUFx6f_ASAP7_75t_L g75 ( 
.A(n_45),
.Y(n_75)
);

INVx4_ASAP7_75t_L g106 ( 
.A(n_75),
.Y(n_106)
);

BUFx6f_ASAP7_75t_L g76 ( 
.A(n_45),
.Y(n_76)
);

INVx4_ASAP7_75t_L g144 ( 
.A(n_76),
.Y(n_144)
);

BUFx6f_ASAP7_75t_L g77 ( 
.A(n_16),
.Y(n_77)
);

BUFx3_ASAP7_75t_L g98 ( 
.A(n_77),
.Y(n_98)
);

INVx2_ASAP7_75t_L g78 ( 
.A(n_29),
.Y(n_78)
);

INVx2_ASAP7_75t_L g116 ( 
.A(n_78),
.Y(n_116)
);

BUFx6f_ASAP7_75t_L g79 ( 
.A(n_20),
.Y(n_79)
);

BUFx3_ASAP7_75t_L g107 ( 
.A(n_79),
.Y(n_107)
);

INVx2_ASAP7_75t_L g80 ( 
.A(n_29),
.Y(n_80)
);

INVx2_ASAP7_75t_L g131 ( 
.A(n_80),
.Y(n_131)
);

INVx4_ASAP7_75t_L g81 ( 
.A(n_20),
.Y(n_81)
);

HB1xp67_ASAP7_75t_L g132 ( 
.A(n_81),
.Y(n_132)
);

INVx8_ASAP7_75t_L g82 ( 
.A(n_20),
.Y(n_82)
);

BUFx3_ASAP7_75t_L g129 ( 
.A(n_82),
.Y(n_129)
);

BUFx6f_ASAP7_75t_L g83 ( 
.A(n_20),
.Y(n_83)
);

BUFx3_ASAP7_75t_L g140 ( 
.A(n_83),
.Y(n_140)
);

INVx2_ASAP7_75t_L g84 ( 
.A(n_30),
.Y(n_84)
);

INVx2_ASAP7_75t_L g139 ( 
.A(n_84),
.Y(n_139)
);

INVx2_ASAP7_75t_L g85 ( 
.A(n_30),
.Y(n_85)
);

HB1xp67_ASAP7_75t_L g137 ( 
.A(n_85),
.Y(n_137)
);

INVx4_ASAP7_75t_L g86 ( 
.A(n_20),
.Y(n_86)
);

HB1xp67_ASAP7_75t_L g138 ( 
.A(n_86),
.Y(n_138)
);

INVx5_ASAP7_75t_L g87 ( 
.A(n_21),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g130 ( 
.A(n_87),
.B(n_89),
.Y(n_130)
);

BUFx6f_ASAP7_75t_L g88 ( 
.A(n_21),
.Y(n_88)
);

INVx6_ASAP7_75t_SL g121 ( 
.A(n_88),
.Y(n_121)
);

INVx5_ASAP7_75t_L g89 ( 
.A(n_21),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_23),
.B(n_6),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_SL g110 ( 
.A(n_90),
.B(n_39),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_SL g91 ( 
.A(n_23),
.B(n_8),
.Y(n_91)
);

O2A1O1Ixp33_ASAP7_75t_L g97 ( 
.A1(n_52),
.A2(n_24),
.B(n_43),
.C(n_42),
.Y(n_97)
);

O2A1O1Ixp33_ASAP7_75t_L g161 ( 
.A1(n_97),
.A2(n_21),
.B(n_88),
.C(n_79),
.Y(n_161)
);

CKINVDCx20_ASAP7_75t_R g103 ( 
.A(n_61),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g183 ( 
.A(n_103),
.B(n_108),
.Y(n_183)
);

OAI22xp5_ASAP7_75t_SL g105 ( 
.A1(n_55),
.A2(n_24),
.B1(n_43),
.B2(n_42),
.Y(n_105)
);

AOI22xp5_ASAP7_75t_L g163 ( 
.A1(n_105),
.A2(n_75),
.B1(n_70),
.B2(n_67),
.Y(n_163)
);

CKINVDCx20_ASAP7_75t_R g108 ( 
.A(n_49),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_SL g109 ( 
.A(n_86),
.B(n_39),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_L g156 ( 
.A(n_109),
.B(n_110),
.Y(n_156)
);

AOI22xp33_ASAP7_75t_SL g113 ( 
.A1(n_73),
.A2(n_66),
.B1(n_26),
.B2(n_74),
.Y(n_113)
);

AOI22xp33_ASAP7_75t_SL g168 ( 
.A1(n_113),
.A2(n_118),
.B1(n_0),
.B2(n_1),
.Y(n_168)
);

AOI22xp33_ASAP7_75t_SL g118 ( 
.A1(n_77),
.A2(n_25),
.B1(n_38),
.B2(n_32),
.Y(n_118)
);

A2O1A1Ixp33_ASAP7_75t_L g153 ( 
.A1(n_119),
.A2(n_125),
.B(n_35),
.C(n_41),
.Y(n_153)
);

A2O1A1Ixp33_ASAP7_75t_L g125 ( 
.A1(n_54),
.A2(n_36),
.B(n_38),
.C(n_25),
.Y(n_125)
);

AND2x2_ASAP7_75t_L g149 ( 
.A(n_134),
.B(n_36),
.Y(n_149)
);

CKINVDCx12_ASAP7_75t_R g136 ( 
.A(n_82),
.Y(n_136)
);

INVx4_ASAP7_75t_SL g160 ( 
.A(n_136),
.Y(n_160)
);

AOI22xp33_ASAP7_75t_L g142 ( 
.A1(n_63),
.A2(n_34),
.B1(n_25),
.B2(n_32),
.Y(n_142)
);

OAI22xp5_ASAP7_75t_SL g176 ( 
.A1(n_142),
.A2(n_0),
.B1(n_3),
.B2(n_4),
.Y(n_176)
);

CKINVDCx20_ASAP7_75t_R g145 ( 
.A(n_97),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_L g195 ( 
.A(n_145),
.B(n_165),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_L g146 ( 
.A(n_99),
.B(n_44),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_L g196 ( 
.A(n_146),
.B(n_148),
.Y(n_196)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_137),
.Y(n_147)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_147),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_L g148 ( 
.A(n_104),
.B(n_34),
.Y(n_148)
);

AND2x2_ASAP7_75t_L g222 ( 
.A(n_149),
.B(n_151),
.Y(n_222)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_137),
.Y(n_150)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_150),
.Y(n_201)
);

OA22x2_ASAP7_75t_L g151 ( 
.A1(n_118),
.A2(n_71),
.B1(n_72),
.B2(n_58),
.Y(n_151)
);

INVx5_ASAP7_75t_SL g152 ( 
.A(n_96),
.Y(n_152)
);

INVx3_ASAP7_75t_L g236 ( 
.A(n_152),
.Y(n_236)
);

OR2x2_ASAP7_75t_L g218 ( 
.A(n_153),
.B(n_154),
.Y(n_218)
);

AOI22xp5_ASAP7_75t_SL g154 ( 
.A1(n_116),
.A2(n_35),
.B1(n_41),
.B2(n_37),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_L g155 ( 
.A(n_131),
.B(n_28),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_L g215 ( 
.A(n_155),
.B(n_191),
.Y(n_215)
);

AOI22xp5_ASAP7_75t_SL g157 ( 
.A1(n_139),
.A2(n_28),
.B1(n_37),
.B2(n_21),
.Y(n_157)
);

INVxp67_ASAP7_75t_L g211 ( 
.A(n_157),
.Y(n_211)
);

AOI22xp5_ASAP7_75t_SL g158 ( 
.A1(n_141),
.A2(n_127),
.B1(n_113),
.B2(n_117),
.Y(n_158)
);

AND2x4_ASAP7_75t_L g228 ( 
.A(n_158),
.B(n_162),
.Y(n_228)
);

BUFx3_ASAP7_75t_L g159 ( 
.A(n_93),
.Y(n_159)
);

INVx4_ASAP7_75t_L g216 ( 
.A(n_159),
.Y(n_216)
);

CKINVDCx16_ASAP7_75t_R g205 ( 
.A(n_161),
.Y(n_205)
);

OAI21xp33_ASAP7_75t_SL g162 ( 
.A1(n_123),
.A2(n_58),
.B(n_76),
.Y(n_162)
);

OAI22xp5_ASAP7_75t_SL g200 ( 
.A1(n_163),
.A2(n_124),
.B1(n_101),
.B2(n_112),
.Y(n_200)
);

AOI22xp5_ASAP7_75t_L g164 ( 
.A1(n_100),
.A2(n_64),
.B1(n_59),
.B2(n_57),
.Y(n_164)
);

OAI22xp5_ASAP7_75t_L g234 ( 
.A1(n_164),
.A2(n_168),
.B1(n_184),
.B2(n_157),
.Y(n_234)
);

CKINVDCx20_ASAP7_75t_R g165 ( 
.A(n_129),
.Y(n_165)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_102),
.Y(n_166)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_166),
.Y(n_213)
);

NOR2xp33_ASAP7_75t_L g167 ( 
.A(n_130),
.B(n_83),
.Y(n_167)
);

NOR2xp33_ASAP7_75t_L g212 ( 
.A(n_167),
.B(n_170),
.Y(n_212)
);

INVx2_ASAP7_75t_L g169 ( 
.A(n_92),
.Y(n_169)
);

INVx2_ASAP7_75t_L g223 ( 
.A(n_169),
.Y(n_223)
);

INVxp67_ASAP7_75t_L g170 ( 
.A(n_138),
.Y(n_170)
);

MAJIxp5_ASAP7_75t_L g171 ( 
.A(n_94),
.B(n_95),
.C(n_133),
.Y(n_171)
);

NOR2xp33_ASAP7_75t_L g204 ( 
.A(n_171),
.B(n_175),
.Y(n_204)
);

FAx1_ASAP7_75t_SL g172 ( 
.A(n_142),
.B(n_8),
.CI(n_2),
.CON(n_172),
.SN(n_172)
);

MAJIxp5_ASAP7_75t_SL g203 ( 
.A(n_172),
.B(n_177),
.C(n_11),
.Y(n_203)
);

AOI22xp33_ASAP7_75t_SL g173 ( 
.A1(n_114),
.A2(n_8),
.B1(n_2),
.B2(n_3),
.Y(n_173)
);

AOI22xp33_ASAP7_75t_SL g198 ( 
.A1(n_173),
.A2(n_111),
.B1(n_143),
.B2(n_144),
.Y(n_198)
);

INVxp67_ASAP7_75t_L g174 ( 
.A(n_138),
.Y(n_174)
);

CKINVDCx14_ASAP7_75t_R g217 ( 
.A(n_174),
.Y(n_217)
);

CKINVDCx20_ASAP7_75t_R g175 ( 
.A(n_129),
.Y(n_175)
);

AOI22xp5_ASAP7_75t_L g197 ( 
.A1(n_176),
.A2(n_179),
.B1(n_193),
.B2(n_10),
.Y(n_197)
);

A2O1A1Ixp33_ASAP7_75t_L g177 ( 
.A1(n_111),
.A2(n_132),
.B(n_126),
.C(n_121),
.Y(n_177)
);

AND2x2_ASAP7_75t_L g178 ( 
.A(n_126),
.B(n_0),
.Y(n_178)
);

AND2x2_ASAP7_75t_SL g210 ( 
.A(n_178),
.B(n_180),
.Y(n_210)
);

OAI22xp5_ASAP7_75t_L g179 ( 
.A1(n_120),
.A2(n_4),
.B1(n_5),
.B2(n_9),
.Y(n_179)
);

AND2x2_ASAP7_75t_L g180 ( 
.A(n_132),
.B(n_5),
.Y(n_180)
);

INVx2_ASAP7_75t_L g181 ( 
.A(n_106),
.Y(n_181)
);

INVx2_ASAP7_75t_L g226 ( 
.A(n_181),
.Y(n_226)
);

INVx2_ASAP7_75t_L g182 ( 
.A(n_106),
.Y(n_182)
);

INVx2_ASAP7_75t_L g233 ( 
.A(n_182),
.Y(n_233)
);

AOI22xp5_ASAP7_75t_L g184 ( 
.A1(n_100),
.A2(n_5),
.B1(n_9),
.B2(n_10),
.Y(n_184)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_115),
.Y(n_185)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_185),
.Y(n_214)
);

CKINVDCx16_ASAP7_75t_R g186 ( 
.A(n_111),
.Y(n_186)
);

NOR2xp33_ASAP7_75t_L g207 ( 
.A(n_186),
.B(n_188),
.Y(n_207)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_115),
.Y(n_187)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_187),
.Y(n_227)
);

INVxp67_ASAP7_75t_L g188 ( 
.A(n_128),
.Y(n_188)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_122),
.Y(n_189)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_189),
.Y(n_229)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_122),
.Y(n_190)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_190),
.Y(n_235)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_114),
.Y(n_191)
);

INVx1_ASAP7_75t_SL g192 ( 
.A(n_135),
.Y(n_192)
);

NAND2xp33_ASAP7_75t_SL g232 ( 
.A(n_192),
.B(n_160),
.Y(n_232)
);

OAI22xp5_ASAP7_75t_SL g193 ( 
.A1(n_120),
.A2(n_9),
.B1(n_10),
.B2(n_11),
.Y(n_193)
);

BUFx3_ASAP7_75t_L g194 ( 
.A(n_107),
.Y(n_194)
);

INVx4_ASAP7_75t_L g231 ( 
.A(n_194),
.Y(n_231)
);

OAI22xp5_ASAP7_75t_L g248 ( 
.A1(n_197),
.A2(n_184),
.B1(n_166),
.B2(n_150),
.Y(n_248)
);

INVxp67_ASAP7_75t_L g260 ( 
.A(n_198),
.Y(n_260)
);

AOI22xp5_ASAP7_75t_L g251 ( 
.A1(n_200),
.A2(n_208),
.B1(n_219),
.B2(n_234),
.Y(n_251)
);

AOI22xp5_ASAP7_75t_L g202 ( 
.A1(n_145),
.A2(n_144),
.B1(n_124),
.B2(n_101),
.Y(n_202)
);

OAI22xp5_ASAP7_75t_SL g243 ( 
.A1(n_202),
.A2(n_206),
.B1(n_209),
.B2(n_220),
.Y(n_243)
);

AO21x1_ASAP7_75t_L g261 ( 
.A1(n_203),
.A2(n_232),
.B(n_186),
.Y(n_261)
);

AOI22xp5_ASAP7_75t_L g206 ( 
.A1(n_176),
.A2(n_112),
.B1(n_143),
.B2(n_98),
.Y(n_206)
);

OAI22xp5_ASAP7_75t_SL g208 ( 
.A1(n_163),
.A2(n_98),
.B1(n_107),
.B2(n_140),
.Y(n_208)
);

AOI22xp5_ASAP7_75t_L g209 ( 
.A1(n_179),
.A2(n_140),
.B1(n_13),
.B2(n_15),
.Y(n_209)
);

OAI22xp5_ASAP7_75t_SL g219 ( 
.A1(n_158),
.A2(n_11),
.B1(n_13),
.B2(n_164),
.Y(n_219)
);

AOI22xp5_ASAP7_75t_L g220 ( 
.A1(n_151),
.A2(n_13),
.B1(n_172),
.B2(n_153),
.Y(n_220)
);

NOR2xp33_ASAP7_75t_L g221 ( 
.A(n_156),
.B(n_183),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_SL g272 ( 
.A(n_221),
.B(n_224),
.Y(n_272)
);

NOR2xp33_ASAP7_75t_L g224 ( 
.A(n_183),
.B(n_146),
.Y(n_224)
);

AOI22xp5_ASAP7_75t_L g225 ( 
.A1(n_151),
.A2(n_172),
.B1(n_193),
.B2(n_161),
.Y(n_225)
);

OAI22xp5_ASAP7_75t_SL g255 ( 
.A1(n_225),
.A2(n_177),
.B1(n_152),
.B2(n_192),
.Y(n_255)
);

NOR2xp33_ASAP7_75t_L g230 ( 
.A(n_149),
.B(n_148),
.Y(n_230)
);

NOR2xp33_ASAP7_75t_L g241 ( 
.A(n_230),
.B(n_218),
.Y(n_241)
);

OAI21xp5_ASAP7_75t_L g237 ( 
.A1(n_218),
.A2(n_154),
.B(n_155),
.Y(n_237)
);

INVxp67_ASAP7_75t_L g303 ( 
.A(n_237),
.Y(n_303)
);

NAND2xp5_ASAP7_75t_SL g238 ( 
.A(n_196),
.B(n_171),
.Y(n_238)
);

NAND2xp5_ASAP7_75t_L g275 ( 
.A(n_238),
.B(n_240),
.Y(n_275)
);

AO22x1_ASAP7_75t_L g239 ( 
.A1(n_203),
.A2(n_205),
.B1(n_225),
.B2(n_228),
.Y(n_239)
);

OR2x2_ASAP7_75t_L g287 ( 
.A(n_239),
.B(n_261),
.Y(n_287)
);

NAND2xp5_ASAP7_75t_L g240 ( 
.A(n_196),
.B(n_180),
.Y(n_240)
);

NOR2xp33_ASAP7_75t_L g280 ( 
.A(n_241),
.B(n_244),
.Y(n_280)
);

NAND2xp5_ASAP7_75t_L g242 ( 
.A(n_215),
.B(n_180),
.Y(n_242)
);

NAND2xp5_ASAP7_75t_L g279 ( 
.A(n_242),
.B(n_245),
.Y(n_279)
);

BUFx12_ASAP7_75t_L g244 ( 
.A(n_231),
.Y(n_244)
);

NAND2xp5_ASAP7_75t_L g245 ( 
.A(n_215),
.B(n_178),
.Y(n_245)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_199),
.Y(n_246)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_246),
.Y(n_281)
);

INVx2_ASAP7_75t_L g247 ( 
.A(n_223),
.Y(n_247)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_247),
.Y(n_290)
);

AOI22xp5_ASAP7_75t_L g274 ( 
.A1(n_248),
.A2(n_255),
.B1(n_270),
.B2(n_273),
.Y(n_274)
);

NOR2xp33_ASAP7_75t_SL g249 ( 
.A(n_195),
.B(n_149),
.Y(n_249)
);

NOR2xp33_ASAP7_75t_SL g298 ( 
.A(n_249),
.B(n_232),
.Y(n_298)
);

CKINVDCx20_ASAP7_75t_R g250 ( 
.A(n_195),
.Y(n_250)
);

CKINVDCx5p33_ASAP7_75t_R g297 ( 
.A(n_250),
.Y(n_297)
);

AOI22xp5_ASAP7_75t_L g252 ( 
.A1(n_234),
.A2(n_151),
.B1(n_178),
.B2(n_147),
.Y(n_252)
);

OAI22xp5_ASAP7_75t_L g276 ( 
.A1(n_252),
.A2(n_258),
.B1(n_263),
.B2(n_268),
.Y(n_276)
);

NOR2xp33_ASAP7_75t_L g253 ( 
.A(n_212),
.B(n_160),
.Y(n_253)
);

NAND2xp5_ASAP7_75t_SL g278 ( 
.A(n_253),
.B(n_259),
.Y(n_278)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_199),
.Y(n_254)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_254),
.Y(n_292)
);

BUFx2_ASAP7_75t_L g256 ( 
.A(n_236),
.Y(n_256)
);

CKINVDCx20_ASAP7_75t_R g277 ( 
.A(n_256),
.Y(n_277)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_201),
.Y(n_257)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_257),
.Y(n_293)
);

A2O1A1Ixp33_ASAP7_75t_SL g258 ( 
.A1(n_228),
.A2(n_222),
.B(n_205),
.C(n_220),
.Y(n_258)
);

NOR2xp33_ASAP7_75t_L g259 ( 
.A(n_212),
.B(n_160),
.Y(n_259)
);

NAND2xp5_ASAP7_75t_SL g262 ( 
.A(n_218),
.B(n_169),
.Y(n_262)
);

NAND2xp5_ASAP7_75t_L g286 ( 
.A(n_262),
.B(n_269),
.Y(n_286)
);

AOI22xp5_ASAP7_75t_L g263 ( 
.A1(n_222),
.A2(n_190),
.B1(n_189),
.B2(n_187),
.Y(n_263)
);

INVx2_ASAP7_75t_L g264 ( 
.A(n_223),
.Y(n_264)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_264),
.Y(n_296)
);

MAJIxp5_ASAP7_75t_L g265 ( 
.A(n_204),
.B(n_175),
.C(n_165),
.Y(n_265)
);

MAJIxp5_ASAP7_75t_L g283 ( 
.A(n_265),
.B(n_210),
.C(n_201),
.Y(n_283)
);

BUFx5_ASAP7_75t_L g266 ( 
.A(n_226),
.Y(n_266)
);

NOR2xp33_ASAP7_75t_L g282 ( 
.A(n_266),
.B(n_236),
.Y(n_282)
);

NOR2xp33_ASAP7_75t_L g267 ( 
.A(n_207),
.B(n_170),
.Y(n_267)
);

NAND2xp5_ASAP7_75t_SL g305 ( 
.A(n_267),
.B(n_271),
.Y(n_305)
);

AOI22xp5_ASAP7_75t_L g268 ( 
.A1(n_222),
.A2(n_185),
.B1(n_191),
.B2(n_152),
.Y(n_268)
);

NAND2xp5_ASAP7_75t_SL g269 ( 
.A(n_210),
.B(n_213),
.Y(n_269)
);

OAI22xp33_ASAP7_75t_SL g270 ( 
.A1(n_211),
.A2(n_181),
.B1(n_182),
.B2(n_159),
.Y(n_270)
);

NOR2xp33_ASAP7_75t_L g271 ( 
.A(n_217),
.B(n_174),
.Y(n_271)
);

OAI22xp5_ASAP7_75t_SL g273 ( 
.A1(n_197),
.A2(n_188),
.B1(n_194),
.B2(n_211),
.Y(n_273)
);

CKINVDCx16_ASAP7_75t_R g308 ( 
.A(n_282),
.Y(n_308)
);

MAJIxp5_ASAP7_75t_L g310 ( 
.A(n_283),
.B(n_284),
.C(n_285),
.Y(n_310)
);

MAJIxp5_ASAP7_75t_L g284 ( 
.A(n_265),
.B(n_210),
.C(n_213),
.Y(n_284)
);

MAJIxp5_ASAP7_75t_L g285 ( 
.A(n_238),
.B(n_210),
.C(n_214),
.Y(n_285)
);

XNOR2xp5_ASAP7_75t_L g288 ( 
.A(n_240),
.B(n_228),
.Y(n_288)
);

XNOR2xp5_ASAP7_75t_SL g317 ( 
.A(n_288),
.B(n_304),
.Y(n_317)
);

AND2x6_ASAP7_75t_L g289 ( 
.A(n_239),
.B(n_228),
.Y(n_289)
);

NOR3xp33_ASAP7_75t_L g324 ( 
.A(n_289),
.B(n_242),
.C(n_266),
.Y(n_324)
);

NOR2xp33_ASAP7_75t_L g291 ( 
.A(n_249),
.B(n_216),
.Y(n_291)
);

NOR2xp33_ASAP7_75t_L g312 ( 
.A(n_291),
.B(n_295),
.Y(n_312)
);

AOI22xp5_ASAP7_75t_L g294 ( 
.A1(n_243),
.A2(n_219),
.B1(n_228),
.B2(n_200),
.Y(n_294)
);

OAI22xp5_ASAP7_75t_SL g321 ( 
.A1(n_294),
.A2(n_268),
.B1(n_263),
.B2(n_258),
.Y(n_321)
);

NOR2xp33_ASAP7_75t_L g295 ( 
.A(n_272),
.B(n_216),
.Y(n_295)
);

NAND2xp5_ASAP7_75t_SL g332 ( 
.A(n_298),
.B(n_233),
.Y(n_332)
);

OAI32xp33_ASAP7_75t_L g299 ( 
.A1(n_239),
.A2(n_202),
.A3(n_206),
.B1(n_208),
.B2(n_209),
.Y(n_299)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_299),
.Y(n_309)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_246),
.Y(n_300)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_300),
.Y(n_330)
);

NAND2xp5_ASAP7_75t_L g301 ( 
.A(n_250),
.B(n_214),
.Y(n_301)
);

NAND2xp5_ASAP7_75t_L g315 ( 
.A(n_301),
.B(n_237),
.Y(n_315)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_254),
.Y(n_302)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_302),
.Y(n_333)
);

XOR2x2_ASAP7_75t_L g304 ( 
.A(n_258),
.B(n_227),
.Y(n_304)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_257),
.Y(n_306)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_306),
.Y(n_334)
);

AOI22xp5_ASAP7_75t_L g307 ( 
.A1(n_276),
.A2(n_243),
.B1(n_248),
.B2(n_255),
.Y(n_307)
);

OAI22xp5_ASAP7_75t_SL g335 ( 
.A1(n_307),
.A2(n_314),
.B1(n_319),
.B2(n_326),
.Y(n_335)
);

NOR2xp33_ASAP7_75t_SL g311 ( 
.A(n_278),
.B(n_262),
.Y(n_311)
);

CKINVDCx14_ASAP7_75t_R g352 ( 
.A(n_311),
.Y(n_352)
);

NOR2xp33_ASAP7_75t_L g313 ( 
.A(n_297),
.B(n_256),
.Y(n_313)
);

NAND2xp5_ASAP7_75t_L g346 ( 
.A(n_313),
.B(n_315),
.Y(n_346)
);

AOI22xp5_ASAP7_75t_L g314 ( 
.A1(n_276),
.A2(n_273),
.B1(n_251),
.B2(n_260),
.Y(n_314)
);

NOR2xp33_ASAP7_75t_L g316 ( 
.A(n_297),
.B(n_256),
.Y(n_316)
);

NAND2xp5_ASAP7_75t_L g351 ( 
.A(n_316),
.B(n_324),
.Y(n_351)
);

OAI21xp33_ASAP7_75t_SL g318 ( 
.A1(n_301),
.A2(n_261),
.B(n_258),
.Y(n_318)
);

AOI22xp5_ASAP7_75t_L g341 ( 
.A1(n_318),
.A2(n_321),
.B1(n_287),
.B2(n_306),
.Y(n_341)
);

AOI22xp5_ASAP7_75t_L g319 ( 
.A1(n_299),
.A2(n_251),
.B1(n_260),
.B2(n_252),
.Y(n_319)
);

OAI21xp5_ASAP7_75t_SL g320 ( 
.A1(n_303),
.A2(n_258),
.B(n_261),
.Y(n_320)
);

AOI21xp5_ASAP7_75t_L g358 ( 
.A1(n_320),
.A2(n_322),
.B(n_332),
.Y(n_358)
);

OAI21xp5_ASAP7_75t_SL g322 ( 
.A1(n_303),
.A2(n_287),
.B(n_298),
.Y(n_322)
);

MAJIxp5_ASAP7_75t_L g323 ( 
.A(n_285),
.B(n_269),
.C(n_245),
.Y(n_323)
);

MAJIxp5_ASAP7_75t_L g336 ( 
.A(n_323),
.B(n_327),
.C(n_284),
.Y(n_336)
);

CKINVDCx20_ASAP7_75t_R g325 ( 
.A(n_305),
.Y(n_325)
);

NOR2xp33_ASAP7_75t_L g350 ( 
.A(n_325),
.B(n_292),
.Y(n_350)
);

AOI22xp5_ASAP7_75t_L g326 ( 
.A1(n_294),
.A2(n_227),
.B1(n_229),
.B2(n_235),
.Y(n_326)
);

MAJIxp5_ASAP7_75t_L g327 ( 
.A(n_283),
.B(n_235),
.C(n_229),
.Y(n_327)
);

AOI22xp5_ASAP7_75t_L g328 ( 
.A1(n_274),
.A2(n_231),
.B1(n_247),
.B2(n_264),
.Y(n_328)
);

OAI22xp5_ASAP7_75t_SL g337 ( 
.A1(n_328),
.A2(n_329),
.B1(n_331),
.B2(n_286),
.Y(n_337)
);

AOI22xp5_ASAP7_75t_L g329 ( 
.A1(n_274),
.A2(n_288),
.B1(n_280),
.B2(n_304),
.Y(n_329)
);

AOI22xp5_ASAP7_75t_L g331 ( 
.A1(n_289),
.A2(n_226),
.B1(n_233),
.B2(n_244),
.Y(n_331)
);

NAND2xp5_ASAP7_75t_L g355 ( 
.A(n_332),
.B(n_281),
.Y(n_355)
);

MAJIxp5_ASAP7_75t_L g360 ( 
.A(n_336),
.B(n_347),
.C(n_317),
.Y(n_360)
);

AOI22xp5_ASAP7_75t_L g377 ( 
.A1(n_337),
.A2(n_314),
.B1(n_326),
.B2(n_328),
.Y(n_377)
);

OAI22xp5_ASAP7_75t_L g338 ( 
.A1(n_309),
.A2(n_287),
.B1(n_286),
.B2(n_275),
.Y(n_338)
);

CKINVDCx14_ASAP7_75t_R g371 ( 
.A(n_338),
.Y(n_371)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_313),
.Y(n_339)
);

INVx1_ASAP7_75t_L g359 ( 
.A(n_339),
.Y(n_359)
);

INVx6_ASAP7_75t_L g340 ( 
.A(n_308),
.Y(n_340)
);

INVx1_ASAP7_75t_L g361 ( 
.A(n_340),
.Y(n_361)
);

OAI22xp5_ASAP7_75t_SL g369 ( 
.A1(n_341),
.A2(n_319),
.B1(n_307),
.B2(n_309),
.Y(n_369)
);

INVx1_ASAP7_75t_L g342 ( 
.A(n_316),
.Y(n_342)
);

INVx1_ASAP7_75t_L g363 ( 
.A(n_342),
.Y(n_363)
);

XOR2xp5_ASAP7_75t_L g343 ( 
.A(n_310),
.B(n_275),
.Y(n_343)
);

XOR2xp5_ASAP7_75t_L g375 ( 
.A(n_343),
.B(n_345),
.Y(n_375)
);

INVx1_ASAP7_75t_SL g344 ( 
.A(n_330),
.Y(n_344)
);

NAND2xp5_ASAP7_75t_L g364 ( 
.A(n_344),
.B(n_349),
.Y(n_364)
);

XOR2xp5_ASAP7_75t_L g345 ( 
.A(n_310),
.B(n_279),
.Y(n_345)
);

MAJIxp5_ASAP7_75t_L g347 ( 
.A(n_327),
.B(n_279),
.C(n_302),
.Y(n_347)
);

INVx1_ASAP7_75t_L g348 ( 
.A(n_330),
.Y(n_348)
);

INVx1_ASAP7_75t_L g365 ( 
.A(n_348),
.Y(n_365)
);

INVx1_ASAP7_75t_L g349 ( 
.A(n_333),
.Y(n_349)
);

NOR2xp33_ASAP7_75t_SL g362 ( 
.A(n_350),
.B(n_311),
.Y(n_362)
);

NAND2xp5_ASAP7_75t_SL g353 ( 
.A(n_325),
.B(n_292),
.Y(n_353)
);

NOR2xp33_ASAP7_75t_L g366 ( 
.A(n_353),
.B(n_354),
.Y(n_366)
);

BUFx6f_ASAP7_75t_L g354 ( 
.A(n_308),
.Y(n_354)
);

NOR2xp33_ASAP7_75t_L g370 ( 
.A(n_355),
.B(n_356),
.Y(n_370)
);

NAND2xp5_ASAP7_75t_L g356 ( 
.A(n_312),
.B(n_281),
.Y(n_356)
);

AND2x2_ASAP7_75t_L g357 ( 
.A(n_312),
.B(n_293),
.Y(n_357)
);

OAI21xp5_ASAP7_75t_SL g368 ( 
.A1(n_357),
.A2(n_358),
.B(n_315),
.Y(n_368)
);

MAJIxp5_ASAP7_75t_L g390 ( 
.A(n_360),
.B(n_367),
.C(n_373),
.Y(n_390)
);

NAND2xp5_ASAP7_75t_L g382 ( 
.A(n_362),
.B(n_369),
.Y(n_382)
);

MAJIxp5_ASAP7_75t_L g367 ( 
.A(n_336),
.B(n_323),
.C(n_329),
.Y(n_367)
);

CKINVDCx20_ASAP7_75t_R g380 ( 
.A(n_368),
.Y(n_380)
);

XOR2x2_ASAP7_75t_L g372 ( 
.A(n_345),
.B(n_317),
.Y(n_372)
);

AOI21xp5_ASAP7_75t_L g381 ( 
.A1(n_372),
.A2(n_378),
.B(n_346),
.Y(n_381)
);

MAJIxp5_ASAP7_75t_L g373 ( 
.A(n_343),
.B(n_322),
.C(n_331),
.Y(n_373)
);

MAJIxp5_ASAP7_75t_L g374 ( 
.A(n_347),
.B(n_320),
.C(n_321),
.Y(n_374)
);

NAND2xp5_ASAP7_75t_SL g394 ( 
.A(n_374),
.B(n_344),
.Y(n_394)
);

XNOR2xp5_ASAP7_75t_L g376 ( 
.A(n_346),
.B(n_337),
.Y(n_376)
);

XOR2xp5_ASAP7_75t_L g379 ( 
.A(n_376),
.B(n_341),
.Y(n_379)
);

OAI22xp5_ASAP7_75t_SL g383 ( 
.A1(n_377),
.A2(n_342),
.B1(n_339),
.B2(n_355),
.Y(n_383)
);

OAI21xp33_ASAP7_75t_L g378 ( 
.A1(n_352),
.A2(n_334),
.B(n_333),
.Y(n_378)
);

NOR2xp33_ASAP7_75t_L g395 ( 
.A(n_379),
.B(n_381),
.Y(n_395)
);

NAND2xp5_ASAP7_75t_L g403 ( 
.A(n_383),
.B(n_385),
.Y(n_403)
);

XOR2xp5_ASAP7_75t_L g384 ( 
.A(n_375),
.B(n_351),
.Y(n_384)
);

NOR2xp33_ASAP7_75t_L g399 ( 
.A(n_384),
.B(n_388),
.Y(n_399)
);

AND2x2_ASAP7_75t_L g385 ( 
.A(n_366),
.B(n_351),
.Y(n_385)
);

A2O1A1Ixp33_ASAP7_75t_L g386 ( 
.A1(n_368),
.A2(n_358),
.B(n_356),
.C(n_357),
.Y(n_386)
);

OAI21xp5_ASAP7_75t_SL g406 ( 
.A1(n_386),
.A2(n_382),
.B(n_387),
.Y(n_406)
);

NOR3xp33_ASAP7_75t_SL g387 ( 
.A(n_370),
.B(n_357),
.C(n_340),
.Y(n_387)
);

NOR3xp33_ASAP7_75t_L g398 ( 
.A(n_387),
.B(n_365),
.C(n_364),
.Y(n_398)
);

XOR2xp5_ASAP7_75t_L g388 ( 
.A(n_375),
.B(n_335),
.Y(n_388)
);

XOR2xp5_ASAP7_75t_L g389 ( 
.A(n_373),
.B(n_335),
.Y(n_389)
);

NAND2xp5_ASAP7_75t_SL g397 ( 
.A(n_389),
.B(n_394),
.Y(n_397)
);

AND2x2_ASAP7_75t_L g391 ( 
.A(n_359),
.B(n_354),
.Y(n_391)
);

NAND2xp5_ASAP7_75t_L g405 ( 
.A(n_391),
.B(n_393),
.Y(n_405)
);

NAND2xp5_ASAP7_75t_L g392 ( 
.A(n_359),
.B(n_354),
.Y(n_392)
);

INVx1_ASAP7_75t_L g400 ( 
.A(n_392),
.Y(n_400)
);

NOR2xp33_ASAP7_75t_SL g393 ( 
.A(n_363),
.B(n_349),
.Y(n_393)
);

OAI21xp33_ASAP7_75t_L g396 ( 
.A1(n_380),
.A2(n_363),
.B(n_371),
.Y(n_396)
);

CKINVDCx16_ASAP7_75t_R g414 ( 
.A(n_396),
.Y(n_414)
);

NAND2xp5_ASAP7_75t_L g408 ( 
.A(n_398),
.B(n_401),
.Y(n_408)
);

OAI21xp5_ASAP7_75t_L g401 ( 
.A1(n_385),
.A2(n_374),
.B(n_377),
.Y(n_401)
);

INVx1_ASAP7_75t_L g402 ( 
.A(n_391),
.Y(n_402)
);

NAND2xp5_ASAP7_75t_L g409 ( 
.A(n_402),
.B(n_404),
.Y(n_409)
);

AOI21xp5_ASAP7_75t_L g404 ( 
.A1(n_383),
.A2(n_369),
.B(n_376),
.Y(n_404)
);

NOR2xp33_ASAP7_75t_L g407 ( 
.A(n_406),
.B(n_384),
.Y(n_407)
);

AOI21x1_ASAP7_75t_L g418 ( 
.A1(n_407),
.A2(n_401),
.B(n_403),
.Y(n_418)
);

MAJIxp5_ASAP7_75t_L g410 ( 
.A(n_397),
.B(n_390),
.C(n_389),
.Y(n_410)
);

NAND2xp5_ASAP7_75t_L g421 ( 
.A(n_410),
.B(n_411),
.Y(n_421)
);

NOR2xp33_ASAP7_75t_L g411 ( 
.A(n_405),
.B(n_361),
.Y(n_411)
);

HB1xp67_ASAP7_75t_L g412 ( 
.A(n_406),
.Y(n_412)
);

NAND2xp5_ASAP7_75t_L g422 ( 
.A(n_412),
.B(n_413),
.Y(n_422)
);

NAND2xp5_ASAP7_75t_L g413 ( 
.A(n_400),
.B(n_361),
.Y(n_413)
);

NOR2xp33_ASAP7_75t_SL g415 ( 
.A(n_395),
.B(n_390),
.Y(n_415)
);

NOR2xp33_ASAP7_75t_L g417 ( 
.A(n_415),
.B(n_388),
.Y(n_417)
);

XNOR2xp5_ASAP7_75t_L g416 ( 
.A(n_399),
.B(n_367),
.Y(n_416)
);

NOR2xp33_ASAP7_75t_SL g420 ( 
.A(n_416),
.B(n_360),
.Y(n_420)
);

NAND2xp5_ASAP7_75t_L g427 ( 
.A(n_417),
.B(n_418),
.Y(n_427)
);

OAI22xp5_ASAP7_75t_L g419 ( 
.A1(n_412),
.A2(n_404),
.B1(n_396),
.B2(n_364),
.Y(n_419)
);

INVxp67_ASAP7_75t_L g424 ( 
.A(n_419),
.Y(n_424)
);

OAI22xp5_ASAP7_75t_L g425 ( 
.A1(n_420),
.A2(n_421),
.B1(n_410),
.B2(n_417),
.Y(n_425)
);

AOI321xp33_ASAP7_75t_L g423 ( 
.A1(n_408),
.A2(n_386),
.A3(n_372),
.B1(n_365),
.B2(n_348),
.C(n_379),
.Y(n_423)
);

FAx1_ASAP7_75t_SL g426 ( 
.A(n_423),
.B(n_409),
.CI(n_414),
.CON(n_426),
.SN(n_426)
);

NAND2xp5_ASAP7_75t_L g429 ( 
.A(n_425),
.B(n_426),
.Y(n_429)
);

NOR2xp33_ASAP7_75t_SL g428 ( 
.A(n_427),
.B(n_422),
.Y(n_428)
);

AOI321xp33_ASAP7_75t_L g431 ( 
.A1(n_428),
.A2(n_426),
.A3(n_300),
.B1(n_277),
.B2(n_296),
.C(n_290),
.Y(n_431)
);

MAJIxp5_ASAP7_75t_L g430 ( 
.A(n_424),
.B(n_334),
.C(n_293),
.Y(n_430)
);

XOR2xp5_ASAP7_75t_L g432 ( 
.A(n_430),
.B(n_290),
.Y(n_432)
);

OAI22xp5_ASAP7_75t_L g433 ( 
.A1(n_431),
.A2(n_432),
.B1(n_429),
.B2(n_277),
.Y(n_433)
);

OAI21xp5_ASAP7_75t_L g434 ( 
.A1(n_433),
.A2(n_296),
.B(n_244),
.Y(n_434)
);

XOR2xp5_ASAP7_75t_L g435 ( 
.A(n_434),
.B(n_244),
.Y(n_435)
);


endmodule