module fake_jpeg_3274_n_75 (n_3, n_2, n_1, n_0, n_4, n_8, n_6, n_5, n_7, n_75);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_8;
input n_6;
input n_5;
input n_7;

output n_75;

wire n_13;
wire n_21;
wire n_57;
wire n_53;
wire n_33;
wire n_54;
wire n_61;
wire n_45;
wire n_23;
wire n_10;
wire n_69;
wire n_27;
wire n_55;
wire n_64;
wire n_22;
wire n_47;
wire n_51;
wire n_14;
wire n_40;
wire n_73;
wire n_19;
wire n_20;
wire n_18;
wire n_59;
wire n_35;
wire n_48;
wire n_68;
wire n_52;
wire n_71;
wire n_46;
wire n_58;
wire n_41;
wire n_60;
wire n_65;
wire n_63;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_16;
wire n_49;
wire n_72;
wire n_24;
wire n_28;
wire n_44;
wire n_26;
wire n_38;
wire n_9;
wire n_36;
wire n_74;
wire n_11;
wire n_62;
wire n_17;
wire n_25;
wire n_31;
wire n_56;
wire n_67;
wire n_29;
wire n_43;
wire n_50;
wire n_37;
wire n_12;
wire n_32;
wire n_70;
wire n_15;
wire n_66;

INVx4_ASAP7_75t_L g9 ( 
.A(n_3),
.Y(n_9)
);

NAND2xp5_ASAP7_75t_L g10 ( 
.A(n_1),
.B(n_3),
.Y(n_10)
);

INVx1_ASAP7_75t_L g11 ( 
.A(n_0),
.Y(n_11)
);

INVx4_ASAP7_75t_L g12 ( 
.A(n_5),
.Y(n_12)
);

CKINVDCx20_ASAP7_75t_R g13 ( 
.A(n_1),
.Y(n_13)
);

NAND2xp5_ASAP7_75t_L g14 ( 
.A(n_6),
.B(n_4),
.Y(n_14)
);

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_8),
.Y(n_15)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_2),
.Y(n_16)
);

BUFx3_ASAP7_75t_L g17 ( 
.A(n_2),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_7),
.Y(n_18)
);

OR2x2_ASAP7_75t_L g19 ( 
.A(n_0),
.B(n_4),
.Y(n_19)
);

INVx2_ASAP7_75t_L g20 ( 
.A(n_9),
.Y(n_20)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_20),
.Y(n_40)
);

INVx5_ASAP7_75t_L g21 ( 
.A(n_9),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_21),
.Y(n_31)
);

NOR2xp33_ASAP7_75t_L g22 ( 
.A(n_14),
.B(n_18),
.Y(n_22)
);

NOR2xp33_ASAP7_75t_L g33 ( 
.A(n_22),
.B(n_23),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_10),
.Y(n_23)
);

INVx6_ASAP7_75t_L g24 ( 
.A(n_17),
.Y(n_24)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_24),
.Y(n_32)
);

INVx4_ASAP7_75t_L g25 ( 
.A(n_9),
.Y(n_25)
);

AND2x2_ASAP7_75t_L g36 ( 
.A(n_25),
.B(n_27),
.Y(n_36)
);

INVx2_ASAP7_75t_L g26 ( 
.A(n_12),
.Y(n_26)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_26),
.Y(n_38)
);

INVx2_ASAP7_75t_L g27 ( 
.A(n_12),
.Y(n_27)
);

NAND2xp5_ASAP7_75t_L g28 ( 
.A(n_10),
.B(n_14),
.Y(n_28)
);

NAND2xp5_ASAP7_75t_L g30 ( 
.A(n_28),
.B(n_14),
.Y(n_30)
);

INVx4_ASAP7_75t_L g29 ( 
.A(n_17),
.Y(n_29)
);

CKINVDCx16_ASAP7_75t_R g37 ( 
.A(n_29),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_SL g46 ( 
.A(n_30),
.B(n_39),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_L g34 ( 
.A(n_28),
.B(n_19),
.Y(n_34)
);

OAI21xp5_ASAP7_75t_SL g47 ( 
.A1(n_34),
.A2(n_20),
.B(n_21),
.Y(n_47)
);

MAJIxp5_ASAP7_75t_L g35 ( 
.A(n_23),
.B(n_19),
.C(n_17),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_35),
.B(n_29),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g39 ( 
.A(n_26),
.B(n_18),
.Y(n_39)
);

AOI22xp5_ASAP7_75t_L g41 ( 
.A1(n_30),
.A2(n_35),
.B1(n_34),
.B2(n_36),
.Y(n_41)
);

NAND2xp5_ASAP7_75t_L g51 ( 
.A(n_41),
.B(n_50),
.Y(n_51)
);

OAI22xp5_ASAP7_75t_L g42 ( 
.A1(n_33),
.A2(n_19),
.B1(n_12),
.B2(n_27),
.Y(n_42)
);

AOI22xp33_ASAP7_75t_L g57 ( 
.A1(n_42),
.A2(n_13),
.B1(n_25),
.B2(n_16),
.Y(n_57)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_36),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_SL g55 ( 
.A(n_43),
.B(n_47),
.Y(n_55)
);

A2O1A1Ixp33_ASAP7_75t_SL g44 ( 
.A1(n_36),
.A2(n_19),
.B(n_24),
.C(n_16),
.Y(n_44)
);

OAI21xp5_ASAP7_75t_L g54 ( 
.A1(n_44),
.A2(n_37),
.B(n_13),
.Y(n_54)
);

BUFx3_ASAP7_75t_L g45 ( 
.A(n_31),
.Y(n_45)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_45),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_SL g48 ( 
.A(n_38),
.B(n_15),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_L g56 ( 
.A(n_48),
.B(n_49),
.Y(n_56)
);

INVx2_ASAP7_75t_L g49 ( 
.A(n_32),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_L g52 ( 
.A(n_41),
.B(n_40),
.Y(n_52)
);

MAJIxp5_ASAP7_75t_L g59 ( 
.A(n_52),
.B(n_49),
.C(n_44),
.Y(n_59)
);

AOI22xp5_ASAP7_75t_L g60 ( 
.A1(n_54),
.A2(n_57),
.B1(n_11),
.B2(n_15),
.Y(n_60)
);

AND2x6_ASAP7_75t_L g58 ( 
.A(n_51),
.B(n_46),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_58),
.B(n_59),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_L g63 ( 
.A(n_60),
.B(n_61),
.Y(n_63)
);

AOI22xp5_ASAP7_75t_L g61 ( 
.A1(n_52),
.A2(n_44),
.B1(n_11),
.B2(n_45),
.Y(n_61)
);

AOI21xp5_ASAP7_75t_SL g62 ( 
.A1(n_58),
.A2(n_55),
.B(n_51),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_L g67 ( 
.A(n_62),
.B(n_64),
.Y(n_67)
);

CKINVDCx20_ASAP7_75t_R g64 ( 
.A(n_61),
.Y(n_64)
);

MAJIxp5_ASAP7_75t_L g66 ( 
.A(n_65),
.B(n_56),
.C(n_54),
.Y(n_66)
);

MAJIxp5_ASAP7_75t_L g69 ( 
.A(n_66),
.B(n_53),
.C(n_44),
.Y(n_69)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_63),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_SL g70 ( 
.A(n_68),
.B(n_31),
.Y(n_70)
);

OAI21xp5_ASAP7_75t_L g71 ( 
.A1(n_69),
.A2(n_67),
.B(n_1),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_L g72 ( 
.A(n_70),
.B(n_0),
.Y(n_72)
);

XNOR2xp5_ASAP7_75t_L g73 ( 
.A(n_71),
.B(n_72),
.Y(n_73)
);

XNOR2xp5_ASAP7_75t_L g74 ( 
.A(n_73),
.B(n_5),
.Y(n_74)
);

OAI221xp5_ASAP7_75t_SL g75 ( 
.A1(n_74),
.A2(n_6),
.B1(n_7),
.B2(n_8),
.C(n_3),
.Y(n_75)
);


endmodule