module fake_jpeg_6348_n_341 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_341);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_341;

wire n_253;
wire n_330;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_340;
wire n_291;
wire n_236;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_260;
wire n_199;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

BUFx6f_ASAP7_75t_L g17 ( 
.A(n_1),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_7),
.Y(n_18)
);

BUFx12f_ASAP7_75t_L g19 ( 
.A(n_15),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_7),
.Y(n_20)
);

BUFx12f_ASAP7_75t_L g21 ( 
.A(n_11),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_12),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_16),
.Y(n_23)
);

BUFx8_ASAP7_75t_L g24 ( 
.A(n_0),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_16),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_12),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_1),
.Y(n_27)
);

CKINVDCx16_ASAP7_75t_R g28 ( 
.A(n_1),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_6),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_8),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_9),
.Y(n_31)
);

INVx4_ASAP7_75t_L g32 ( 
.A(n_11),
.Y(n_32)
);

BUFx2_ASAP7_75t_L g33 ( 
.A(n_4),
.Y(n_33)
);

BUFx3_ASAP7_75t_L g34 ( 
.A(n_11),
.Y(n_34)
);

BUFx3_ASAP7_75t_L g35 ( 
.A(n_1),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_10),
.Y(n_36)
);

BUFx12_ASAP7_75t_L g37 ( 
.A(n_24),
.Y(n_37)
);

INVx3_ASAP7_75t_L g52 ( 
.A(n_37),
.Y(n_52)
);

BUFx3_ASAP7_75t_L g38 ( 
.A(n_19),
.Y(n_38)
);

INVx4_ASAP7_75t_L g58 ( 
.A(n_38),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g39 ( 
.A(n_33),
.B(n_32),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g51 ( 
.A(n_39),
.B(n_40),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g40 ( 
.A(n_33),
.B(n_8),
.Y(n_40)
);

INVx2_ASAP7_75t_L g41 ( 
.A(n_33),
.Y(n_41)
);

INVx6_ASAP7_75t_L g63 ( 
.A(n_41),
.Y(n_63)
);

INVx11_ASAP7_75t_L g42 ( 
.A(n_17),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_42),
.B(n_43),
.Y(n_62)
);

INVx6_ASAP7_75t_SL g43 ( 
.A(n_19),
.Y(n_43)
);

NAND2xp5_ASAP7_75t_L g44 ( 
.A(n_24),
.B(n_0),
.Y(n_44)
);

NAND2xp5_ASAP7_75t_SL g59 ( 
.A(n_44),
.B(n_45),
.Y(n_59)
);

AND2x2_ASAP7_75t_L g45 ( 
.A(n_24),
.B(n_0),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_33),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_46),
.Y(n_55)
);

INVx11_ASAP7_75t_L g47 ( 
.A(n_17),
.Y(n_47)
);

AOI22xp33_ASAP7_75t_SL g50 ( 
.A1(n_47),
.A2(n_32),
.B1(n_28),
.B2(n_18),
.Y(n_50)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_34),
.Y(n_48)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_48),
.Y(n_54)
);

HB1xp67_ASAP7_75t_L g49 ( 
.A(n_43),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_49),
.B(n_53),
.Y(n_90)
);

INVxp67_ASAP7_75t_L g93 ( 
.A(n_50),
.Y(n_93)
);

INVx2_ASAP7_75t_L g53 ( 
.A(n_38),
.Y(n_53)
);

INVx2_ASAP7_75t_SL g56 ( 
.A(n_43),
.Y(n_56)
);

INVx11_ASAP7_75t_L g84 ( 
.A(n_56),
.Y(n_84)
);

INVx6_ASAP7_75t_SL g57 ( 
.A(n_43),
.Y(n_57)
);

BUFx2_ASAP7_75t_SL g97 ( 
.A(n_57),
.Y(n_97)
);

INVx3_ASAP7_75t_L g60 ( 
.A(n_37),
.Y(n_60)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_60),
.Y(n_68)
);

AOI22xp33_ASAP7_75t_SL g61 ( 
.A1(n_42),
.A2(n_32),
.B1(n_28),
.B2(n_27),
.Y(n_61)
);

AOI21xp5_ASAP7_75t_L g87 ( 
.A1(n_61),
.A2(n_34),
.B(n_35),
.Y(n_87)
);

AOI22xp33_ASAP7_75t_L g64 ( 
.A1(n_42),
.A2(n_36),
.B1(n_31),
.B2(n_30),
.Y(n_64)
);

OAI22xp5_ASAP7_75t_L g101 ( 
.A1(n_64),
.A2(n_66),
.B1(n_67),
.B2(n_23),
.Y(n_101)
);

BUFx12f_ASAP7_75t_L g65 ( 
.A(n_37),
.Y(n_65)
);

BUFx3_ASAP7_75t_L g80 ( 
.A(n_65),
.Y(n_80)
);

OAI22xp5_ASAP7_75t_L g66 ( 
.A1(n_42),
.A2(n_27),
.B1(n_31),
.B2(n_30),
.Y(n_66)
);

AOI22xp5_ASAP7_75t_L g67 ( 
.A1(n_47),
.A2(n_36),
.B1(n_23),
.B2(n_25),
.Y(n_67)
);

XNOR2xp5_ASAP7_75t_L g69 ( 
.A(n_59),
.B(n_44),
.Y(n_69)
);

XNOR2xp5_ASAP7_75t_SL g109 ( 
.A(n_69),
.B(n_45),
.Y(n_109)
);

INVx3_ASAP7_75t_L g70 ( 
.A(n_57),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g106 ( 
.A(n_70),
.B(n_73),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_SL g71 ( 
.A(n_51),
.B(n_40),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_SL g105 ( 
.A(n_71),
.B(n_89),
.Y(n_105)
);

AOI22xp33_ASAP7_75t_L g72 ( 
.A1(n_63),
.A2(n_47),
.B1(n_41),
.B2(n_48),
.Y(n_72)
);

AOI22xp33_ASAP7_75t_SL g102 ( 
.A1(n_72),
.A2(n_76),
.B1(n_83),
.B2(n_87),
.Y(n_102)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_66),
.Y(n_73)
);

INVx4_ASAP7_75t_L g74 ( 
.A(n_63),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g115 ( 
.A(n_74),
.B(n_75),
.Y(n_115)
);

INVx3_ASAP7_75t_L g75 ( 
.A(n_55),
.Y(n_75)
);

AOI22xp33_ASAP7_75t_SL g76 ( 
.A1(n_56),
.A2(n_47),
.B1(n_41),
.B2(n_25),
.Y(n_76)
);

INVx2_ASAP7_75t_L g77 ( 
.A(n_63),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g121 ( 
.A(n_77),
.B(n_78),
.Y(n_121)
);

INVx2_ASAP7_75t_L g78 ( 
.A(n_55),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_L g79 ( 
.A(n_59),
.B(n_44),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_SL g107 ( 
.A(n_79),
.B(n_81),
.Y(n_107)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_67),
.Y(n_81)
);

OA22x2_ASAP7_75t_L g82 ( 
.A1(n_49),
.A2(n_45),
.B1(n_41),
.B2(n_46),
.Y(n_82)
);

AOI22xp5_ASAP7_75t_SL g125 ( 
.A1(n_82),
.A2(n_60),
.B1(n_52),
.B2(n_46),
.Y(n_125)
);

AOI22xp33_ASAP7_75t_L g83 ( 
.A1(n_54),
.A2(n_48),
.B1(n_39),
.B2(n_45),
.Y(n_83)
);

OAI21xp5_ASAP7_75t_SL g85 ( 
.A1(n_51),
.A2(n_39),
.B(n_40),
.Y(n_85)
);

INVxp67_ASAP7_75t_L g103 ( 
.A(n_85),
.Y(n_103)
);

INVx3_ASAP7_75t_L g86 ( 
.A(n_53),
.Y(n_86)
);

BUFx6f_ASAP7_75t_L g104 ( 
.A(n_86),
.Y(n_104)
);

INVx2_ASAP7_75t_L g88 ( 
.A(n_55),
.Y(n_88)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_88),
.Y(n_123)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_62),
.Y(n_89)
);

BUFx12_ASAP7_75t_L g91 ( 
.A(n_65),
.Y(n_91)
);

INVx3_ASAP7_75t_L g114 ( 
.A(n_91),
.Y(n_114)
);

INVx2_ASAP7_75t_L g92 ( 
.A(n_54),
.Y(n_92)
);

CKINVDCx20_ASAP7_75t_R g111 ( 
.A(n_92),
.Y(n_111)
);

INVx2_ASAP7_75t_L g94 ( 
.A(n_58),
.Y(n_94)
);

INVx3_ASAP7_75t_L g120 ( 
.A(n_94),
.Y(n_120)
);

INVxp67_ASAP7_75t_L g95 ( 
.A(n_62),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_SL g119 ( 
.A(n_95),
.B(n_99),
.Y(n_119)
);

INVx3_ASAP7_75t_L g96 ( 
.A(n_58),
.Y(n_96)
);

INVx5_ASAP7_75t_L g110 ( 
.A(n_96),
.Y(n_110)
);

INVx6_ASAP7_75t_L g98 ( 
.A(n_65),
.Y(n_98)
);

BUFx6f_ASAP7_75t_L g113 ( 
.A(n_98),
.Y(n_113)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_58),
.Y(n_99)
);

INVx6_ASAP7_75t_L g100 ( 
.A(n_65),
.Y(n_100)
);

INVx5_ASAP7_75t_L g130 ( 
.A(n_100),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_SL g122 ( 
.A(n_101),
.B(n_26),
.Y(n_122)
);

AND2x2_ASAP7_75t_L g108 ( 
.A(n_82),
.B(n_45),
.Y(n_108)
);

OAI21xp5_ASAP7_75t_SL g160 ( 
.A1(n_108),
.A2(n_126),
.B(n_127),
.Y(n_160)
);

XNOR2xp5_ASAP7_75t_SL g137 ( 
.A(n_109),
.B(n_37),
.Y(n_137)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_90),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_L g139 ( 
.A(n_112),
.B(n_117),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_L g116 ( 
.A(n_95),
.B(n_45),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_L g148 ( 
.A(n_116),
.B(n_118),
.Y(n_148)
);

INVxp67_ASAP7_75t_L g117 ( 
.A(n_72),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_L g118 ( 
.A(n_82),
.B(n_56),
.Y(n_118)
);

AOI22xp5_ASAP7_75t_L g154 ( 
.A1(n_122),
.A2(n_22),
.B1(n_20),
.B2(n_17),
.Y(n_154)
);

INVxp67_ASAP7_75t_L g124 ( 
.A(n_97),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_L g152 ( 
.A(n_124),
.B(n_128),
.Y(n_152)
);

OAI22xp5_ASAP7_75t_SL g134 ( 
.A1(n_125),
.A2(n_74),
.B1(n_86),
.B2(n_52),
.Y(n_134)
);

AND2x2_ASAP7_75t_L g126 ( 
.A(n_83),
.B(n_24),
.Y(n_126)
);

AND2x2_ASAP7_75t_L g127 ( 
.A(n_93),
.B(n_24),
.Y(n_127)
);

INVxp67_ASAP7_75t_L g128 ( 
.A(n_76),
.Y(n_128)
);

INVx2_ASAP7_75t_L g129 ( 
.A(n_80),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_L g161 ( 
.A(n_129),
.B(n_104),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_SL g131 ( 
.A(n_68),
.B(n_26),
.Y(n_131)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_131),
.Y(n_138)
);

INVx4_ASAP7_75t_L g132 ( 
.A(n_130),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_L g170 ( 
.A(n_132),
.B(n_135),
.Y(n_170)
);

MAJIxp5_ASAP7_75t_L g133 ( 
.A(n_109),
.B(n_93),
.C(n_38),
.Y(n_133)
);

MAJIxp5_ASAP7_75t_L g174 ( 
.A(n_133),
.B(n_142),
.C(n_145),
.Y(n_174)
);

AOI22xp5_ASAP7_75t_L g183 ( 
.A1(n_134),
.A2(n_140),
.B1(n_144),
.B2(n_149),
.Y(n_183)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_121),
.Y(n_135)
);

AOI22xp33_ASAP7_75t_L g136 ( 
.A1(n_102),
.A2(n_128),
.B1(n_125),
.B2(n_127),
.Y(n_136)
);

CKINVDCx16_ASAP7_75t_R g162 ( 
.A(n_136),
.Y(n_162)
);

XNOR2xp5_ASAP7_75t_L g163 ( 
.A(n_137),
.B(n_153),
.Y(n_163)
);

OAI22xp5_ASAP7_75t_SL g140 ( 
.A1(n_118),
.A2(n_84),
.B1(n_46),
.B2(n_18),
.Y(n_140)
);

INVxp67_ASAP7_75t_L g141 ( 
.A(n_130),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_SL g173 ( 
.A(n_141),
.B(n_146),
.Y(n_173)
);

XOR2xp5_ASAP7_75t_L g142 ( 
.A(n_116),
.B(n_108),
.Y(n_142)
);

BUFx2_ASAP7_75t_L g143 ( 
.A(n_110),
.Y(n_143)
);

INVx3_ASAP7_75t_L g167 ( 
.A(n_143),
.Y(n_167)
);

OAI22xp5_ASAP7_75t_SL g144 ( 
.A1(n_117),
.A2(n_84),
.B1(n_46),
.B2(n_29),
.Y(n_144)
);

MAJIxp5_ASAP7_75t_L g145 ( 
.A(n_107),
.B(n_38),
.C(n_65),
.Y(n_145)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_115),
.Y(n_146)
);

INVxp67_ASAP7_75t_L g147 ( 
.A(n_110),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_SL g181 ( 
.A(n_147),
.B(n_154),
.Y(n_181)
);

OAI22xp5_ASAP7_75t_SL g149 ( 
.A1(n_103),
.A2(n_29),
.B1(n_98),
.B2(n_100),
.Y(n_149)
);

AOI22xp5_ASAP7_75t_SL g150 ( 
.A1(n_103),
.A2(n_20),
.B1(n_22),
.B2(n_21),
.Y(n_150)
);

OAI21xp5_ASAP7_75t_L g165 ( 
.A1(n_150),
.A2(n_155),
.B(n_160),
.Y(n_165)
);

OAI21xp5_ASAP7_75t_L g151 ( 
.A1(n_105),
.A2(n_37),
.B(n_19),
.Y(n_151)
);

OAI21xp5_ASAP7_75t_SL g169 ( 
.A1(n_151),
.A2(n_158),
.B(n_111),
.Y(n_169)
);

MAJIxp5_ASAP7_75t_L g153 ( 
.A(n_108),
.B(n_91),
.C(n_37),
.Y(n_153)
);

AOI22xp5_ASAP7_75t_L g155 ( 
.A1(n_126),
.A2(n_22),
.B1(n_20),
.B2(n_37),
.Y(n_155)
);

OAI22xp5_ASAP7_75t_SL g164 ( 
.A1(n_155),
.A2(n_124),
.B1(n_120),
.B2(n_112),
.Y(n_164)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_106),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_SL g191 ( 
.A(n_156),
.B(n_113),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_L g157 ( 
.A(n_119),
.B(n_21),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_L g168 ( 
.A(n_157),
.B(n_148),
.Y(n_168)
);

OAI21xp5_ASAP7_75t_L g158 ( 
.A1(n_126),
.A2(n_21),
.B(n_19),
.Y(n_158)
);

INVx2_ASAP7_75t_L g159 ( 
.A(n_104),
.Y(n_159)
);

CKINVDCx20_ASAP7_75t_R g185 ( 
.A(n_159),
.Y(n_185)
);

CKINVDCx20_ASAP7_75t_R g192 ( 
.A(n_161),
.Y(n_192)
);

AOI22xp5_ASAP7_75t_L g208 ( 
.A1(n_164),
.A2(n_2),
.B1(n_3),
.B2(n_4),
.Y(n_208)
);

NOR2xp33_ASAP7_75t_L g226 ( 
.A(n_165),
.B(n_175),
.Y(n_226)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_139),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_SL g200 ( 
.A(n_166),
.B(n_171),
.Y(n_200)
);

NAND2xp5_ASAP7_75t_L g196 ( 
.A(n_168),
.B(n_179),
.Y(n_196)
);

OAI21xp5_ASAP7_75t_L g215 ( 
.A1(n_169),
.A2(n_177),
.B(n_178),
.Y(n_215)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_157),
.Y(n_171)
);

XNOR2xp5_ASAP7_75t_L g172 ( 
.A(n_137),
.B(n_127),
.Y(n_172)
);

XNOR2xp5_ASAP7_75t_L g212 ( 
.A(n_172),
.B(n_182),
.Y(n_212)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_149),
.Y(n_175)
);

INVx2_ASAP7_75t_L g176 ( 
.A(n_143),
.Y(n_176)
);

CKINVDCx20_ASAP7_75t_R g199 ( 
.A(n_176),
.Y(n_199)
);

AND2x2_ASAP7_75t_SL g177 ( 
.A(n_160),
.B(n_19),
.Y(n_177)
);

OAI21xp5_ASAP7_75t_SL g178 ( 
.A1(n_148),
.A2(n_129),
.B(n_123),
.Y(n_178)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_144),
.Y(n_179)
);

CKINVDCx16_ASAP7_75t_R g180 ( 
.A(n_154),
.Y(n_180)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_180),
.Y(n_197)
);

OAI21xp5_ASAP7_75t_SL g182 ( 
.A1(n_153),
.A2(n_21),
.B(n_35),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_L g184 ( 
.A(n_142),
.B(n_21),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_L g204 ( 
.A(n_184),
.B(n_189),
.Y(n_204)
);

AOI322xp5_ASAP7_75t_L g186 ( 
.A1(n_158),
.A2(n_34),
.A3(n_35),
.B1(n_91),
.B2(n_113),
.C1(n_120),
.C2(n_114),
.Y(n_186)
);

MAJIxp5_ASAP7_75t_L g224 ( 
.A(n_186),
.B(n_187),
.C(n_190),
.Y(n_224)
);

XNOR2xp5_ASAP7_75t_SL g187 ( 
.A(n_140),
.B(n_10),
.Y(n_187)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_150),
.Y(n_188)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_188),
.Y(n_202)
);

NAND2xp5_ASAP7_75t_L g189 ( 
.A(n_145),
.B(n_0),
.Y(n_189)
);

XNOR2xp5_ASAP7_75t_L g190 ( 
.A(n_133),
.B(n_80),
.Y(n_190)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_191),
.Y(n_217)
);

CKINVDCx20_ASAP7_75t_R g193 ( 
.A(n_159),
.Y(n_193)
);

CKINVDCx20_ASAP7_75t_R g216 ( 
.A(n_193),
.Y(n_216)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_134),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_L g207 ( 
.A(n_194),
.B(n_195),
.Y(n_207)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_152),
.Y(n_195)
);

OAI22xp5_ASAP7_75t_SL g198 ( 
.A1(n_194),
.A2(n_146),
.B1(n_135),
.B2(n_151),
.Y(n_198)
);

AOI22xp5_ASAP7_75t_L g239 ( 
.A1(n_198),
.A2(n_203),
.B1(n_222),
.B2(n_167),
.Y(n_239)
);

AND2x2_ASAP7_75t_L g201 ( 
.A(n_177),
.B(n_141),
.Y(n_201)
);

OAI21xp5_ASAP7_75t_SL g230 ( 
.A1(n_201),
.A2(n_169),
.B(n_182),
.Y(n_230)
);

OAI22xp5_ASAP7_75t_L g203 ( 
.A1(n_183),
.A2(n_138),
.B1(n_147),
.B2(n_114),
.Y(n_203)
);

INVxp67_ASAP7_75t_L g205 ( 
.A(n_170),
.Y(n_205)
);

NAND2xp5_ASAP7_75t_SL g236 ( 
.A(n_205),
.B(n_220),
.Y(n_236)
);

AOI22xp5_ASAP7_75t_SL g206 ( 
.A1(n_177),
.A2(n_132),
.B1(n_3),
.B2(n_4),
.Y(n_206)
);

OAI22xp5_ASAP7_75t_SL g231 ( 
.A1(n_206),
.A2(n_213),
.B1(n_223),
.B2(n_187),
.Y(n_231)
);

CKINVDCx14_ASAP7_75t_R g237 ( 
.A(n_208),
.Y(n_237)
);

NAND2xp5_ASAP7_75t_L g209 ( 
.A(n_168),
.B(n_2),
.Y(n_209)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_209),
.Y(n_227)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_173),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_L g233 ( 
.A(n_210),
.B(n_214),
.Y(n_233)
);

NAND2xp5_ASAP7_75t_L g211 ( 
.A(n_178),
.B(n_2),
.Y(n_211)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_211),
.Y(n_228)
);

AOI22xp5_ASAP7_75t_L g213 ( 
.A1(n_162),
.A2(n_3),
.B1(n_5),
.B2(n_6),
.Y(n_213)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_164),
.Y(n_214)
);

CKINVDCx20_ASAP7_75t_R g218 ( 
.A(n_185),
.Y(n_218)
);

NOR2xp33_ASAP7_75t_SL g247 ( 
.A(n_218),
.B(n_221),
.Y(n_247)
);

BUFx3_ASAP7_75t_L g219 ( 
.A(n_176),
.Y(n_219)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_219),
.Y(n_229)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_183),
.Y(n_220)
);

CKINVDCx16_ASAP7_75t_R g221 ( 
.A(n_181),
.Y(n_221)
);

OAI22xp5_ASAP7_75t_SL g222 ( 
.A1(n_179),
.A2(n_5),
.B1(n_6),
.B2(n_7),
.Y(n_222)
);

AOI22xp5_ASAP7_75t_L g223 ( 
.A1(n_165),
.A2(n_174),
.B1(n_195),
.B2(n_189),
.Y(n_223)
);

MAJIxp5_ASAP7_75t_L g225 ( 
.A(n_174),
.B(n_16),
.C(n_8),
.Y(n_225)
);

MAJIxp5_ASAP7_75t_L g234 ( 
.A(n_225),
.B(n_184),
.C(n_192),
.Y(n_234)
);

MAJIxp5_ASAP7_75t_L g257 ( 
.A(n_230),
.B(n_241),
.C(n_243),
.Y(n_257)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_231),
.Y(n_254)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_200),
.Y(n_232)
);

NAND2xp5_ASAP7_75t_L g268 ( 
.A(n_232),
.B(n_250),
.Y(n_268)
);

NOR2xp33_ASAP7_75t_SL g271 ( 
.A(n_234),
.B(n_201),
.Y(n_271)
);

XNOR2xp5_ASAP7_75t_L g235 ( 
.A(n_212),
.B(n_163),
.Y(n_235)
);

XOR2xp5_ASAP7_75t_L g258 ( 
.A(n_235),
.B(n_238),
.Y(n_258)
);

XOR2xp5_ASAP7_75t_L g238 ( 
.A(n_212),
.B(n_163),
.Y(n_238)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_239),
.Y(n_255)
);

AOI22xp5_ASAP7_75t_L g240 ( 
.A1(n_214),
.A2(n_172),
.B1(n_190),
.B2(n_167),
.Y(n_240)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_240),
.Y(n_256)
);

MAJIxp5_ASAP7_75t_L g241 ( 
.A(n_223),
.B(n_15),
.C(n_9),
.Y(n_241)
);

AOI21xp5_ASAP7_75t_L g242 ( 
.A1(n_215),
.A2(n_5),
.B(n_9),
.Y(n_242)
);

XNOR2xp5_ASAP7_75t_L g253 ( 
.A(n_242),
.B(n_211),
.Y(n_253)
);

XOR2xp5_ASAP7_75t_L g243 ( 
.A(n_215),
.B(n_15),
.Y(n_243)
);

XOR2xp5_ASAP7_75t_L g244 ( 
.A(n_204),
.B(n_10),
.Y(n_244)
);

MAJIxp5_ASAP7_75t_L g260 ( 
.A(n_244),
.B(n_245),
.C(n_246),
.Y(n_260)
);

MAJIxp5_ASAP7_75t_L g245 ( 
.A(n_204),
.B(n_12),
.C(n_13),
.Y(n_245)
);

MAJIxp5_ASAP7_75t_L g246 ( 
.A(n_224),
.B(n_13),
.C(n_14),
.Y(n_246)
);

NOR2xp33_ASAP7_75t_SL g248 ( 
.A(n_210),
.B(n_13),
.Y(n_248)
);

NAND2xp5_ASAP7_75t_SL g266 ( 
.A(n_248),
.B(n_222),
.Y(n_266)
);

XNOR2xp5_ASAP7_75t_SL g249 ( 
.A(n_196),
.B(n_14),
.Y(n_249)
);

XNOR2xp5_ASAP7_75t_SL g270 ( 
.A(n_249),
.B(n_209),
.Y(n_270)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_219),
.Y(n_250)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_207),
.Y(n_251)
);

NAND2xp5_ASAP7_75t_L g269 ( 
.A(n_251),
.B(n_207),
.Y(n_269)
);

CKINVDCx20_ASAP7_75t_R g252 ( 
.A(n_247),
.Y(n_252)
);

OAI21xp5_ASAP7_75t_SL g283 ( 
.A1(n_252),
.A2(n_227),
.B(n_245),
.Y(n_283)
);

XNOR2xp5_ASAP7_75t_L g274 ( 
.A(n_253),
.B(n_263),
.Y(n_274)
);

XNOR2xp5_ASAP7_75t_L g259 ( 
.A(n_235),
.B(n_224),
.Y(n_259)
);

XOR2xp5_ASAP7_75t_L g275 ( 
.A(n_259),
.B(n_234),
.Y(n_275)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_233),
.Y(n_261)
);

NAND2xp5_ASAP7_75t_L g284 ( 
.A(n_261),
.B(n_262),
.Y(n_284)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_249),
.Y(n_262)
);

MAJIxp5_ASAP7_75t_L g263 ( 
.A(n_238),
.B(n_225),
.C(n_196),
.Y(n_263)
);

AOI21x1_ASAP7_75t_L g264 ( 
.A1(n_230),
.A2(n_201),
.B(n_243),
.Y(n_264)
);

XNOR2x1_ASAP7_75t_L g273 ( 
.A(n_264),
.B(n_240),
.Y(n_273)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_239),
.Y(n_265)
);

NAND2xp5_ASAP7_75t_L g287 ( 
.A(n_265),
.B(n_266),
.Y(n_287)
);

INVxp33_ASAP7_75t_SL g267 ( 
.A(n_236),
.Y(n_267)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_267),
.Y(n_278)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_269),
.Y(n_286)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_270),
.Y(n_290)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_271),
.Y(n_288)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_244),
.Y(n_272)
);

NAND2xp5_ASAP7_75t_L g289 ( 
.A(n_272),
.B(n_226),
.Y(n_289)
);

XOR2xp5_ASAP7_75t_L g301 ( 
.A(n_273),
.B(n_275),
.Y(n_301)
);

NOR2xp33_ASAP7_75t_SL g276 ( 
.A(n_268),
.B(n_228),
.Y(n_276)
);

NAND2xp5_ASAP7_75t_SL g292 ( 
.A(n_276),
.B(n_205),
.Y(n_292)
);

HB1xp67_ASAP7_75t_L g277 ( 
.A(n_267),
.Y(n_277)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_277),
.Y(n_297)
);

XOR2xp5_ASAP7_75t_L g279 ( 
.A(n_258),
.B(n_231),
.Y(n_279)
);

XOR2xp5_ASAP7_75t_L g305 ( 
.A(n_279),
.B(n_280),
.Y(n_305)
);

XOR2xp5_ASAP7_75t_L g280 ( 
.A(n_258),
.B(n_241),
.Y(n_280)
);

XOR2xp5_ASAP7_75t_L g281 ( 
.A(n_259),
.B(n_242),
.Y(n_281)
);

MAJIxp5_ASAP7_75t_L g303 ( 
.A(n_281),
.B(n_282),
.C(n_260),
.Y(n_303)
);

XOR2xp5_ASAP7_75t_L g282 ( 
.A(n_263),
.B(n_246),
.Y(n_282)
);

OAI21xp5_ASAP7_75t_SL g304 ( 
.A1(n_283),
.A2(n_289),
.B(n_217),
.Y(n_304)
);

AND2x2_ASAP7_75t_SL g285 ( 
.A(n_264),
.B(n_254),
.Y(n_285)
);

AOI21xp5_ASAP7_75t_L g291 ( 
.A1(n_285),
.A2(n_256),
.B(n_255),
.Y(n_291)
);

AOI21xp5_ASAP7_75t_L g308 ( 
.A1(n_291),
.A2(n_295),
.B(n_298),
.Y(n_308)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_292),
.Y(n_309)
);

XNOR2xp5_ASAP7_75t_L g293 ( 
.A(n_279),
.B(n_270),
.Y(n_293)
);

XOR2xp5_ASAP7_75t_L g315 ( 
.A(n_293),
.B(n_303),
.Y(n_315)
);

BUFx24_ASAP7_75t_SL g294 ( 
.A(n_288),
.Y(n_294)
);

NOR2xp33_ASAP7_75t_L g310 ( 
.A(n_294),
.B(n_296),
.Y(n_310)
);

CKINVDCx20_ASAP7_75t_R g295 ( 
.A(n_287),
.Y(n_295)
);

INVx11_ASAP7_75t_L g296 ( 
.A(n_278),
.Y(n_296)
);

AOI21xp5_ASAP7_75t_L g298 ( 
.A1(n_285),
.A2(n_197),
.B(n_257),
.Y(n_298)
);

NAND2xp5_ASAP7_75t_L g299 ( 
.A(n_286),
.B(n_216),
.Y(n_299)
);

AOI21xp5_ASAP7_75t_L g311 ( 
.A1(n_299),
.A2(n_300),
.B(n_302),
.Y(n_311)
);

AOI21xp5_ASAP7_75t_L g300 ( 
.A1(n_285),
.A2(n_257),
.B(n_199),
.Y(n_300)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_284),
.Y(n_302)
);

NAND2xp5_ASAP7_75t_L g307 ( 
.A(n_304),
.B(n_253),
.Y(n_307)
);

NAND2xp5_ASAP7_75t_SL g306 ( 
.A(n_297),
.B(n_229),
.Y(n_306)
);

OAI21xp5_ASAP7_75t_SL g322 ( 
.A1(n_306),
.A2(n_307),
.B(n_298),
.Y(n_322)
);

AND2x2_ASAP7_75t_L g312 ( 
.A(n_301),
.B(n_273),
.Y(n_312)
);

NAND2xp5_ASAP7_75t_L g326 ( 
.A(n_312),
.B(n_316),
.Y(n_326)
);

XNOR2xp5_ASAP7_75t_L g313 ( 
.A(n_303),
.B(n_274),
.Y(n_313)
);

XOR2xp5_ASAP7_75t_L g321 ( 
.A(n_313),
.B(n_305),
.Y(n_321)
);

OAI22xp5_ASAP7_75t_SL g314 ( 
.A1(n_296),
.A2(n_290),
.B1(n_237),
.B2(n_202),
.Y(n_314)
);

INVxp67_ASAP7_75t_L g325 ( 
.A(n_314),
.Y(n_325)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_300),
.Y(n_316)
);

HB1xp67_ASAP7_75t_L g317 ( 
.A(n_291),
.Y(n_317)
);

NOR2xp33_ASAP7_75t_L g324 ( 
.A(n_317),
.B(n_198),
.Y(n_324)
);

NOR2xp33_ASAP7_75t_SL g318 ( 
.A(n_310),
.B(n_311),
.Y(n_318)
);

AOI21xp5_ASAP7_75t_L g328 ( 
.A1(n_318),
.A2(n_319),
.B(n_322),
.Y(n_328)
);

NOR2xp67_ASAP7_75t_SL g319 ( 
.A(n_312),
.B(n_301),
.Y(n_319)
);

MAJIxp5_ASAP7_75t_L g320 ( 
.A(n_315),
.B(n_305),
.C(n_275),
.Y(n_320)
);

MAJIxp5_ASAP7_75t_L g329 ( 
.A(n_320),
.B(n_321),
.C(n_315),
.Y(n_329)
);

NOR2xp33_ASAP7_75t_L g323 ( 
.A(n_317),
.B(n_208),
.Y(n_323)
);

NAND2xp5_ASAP7_75t_SL g331 ( 
.A(n_323),
.B(n_324),
.Y(n_331)
);

NAND2xp5_ASAP7_75t_L g327 ( 
.A(n_325),
.B(n_309),
.Y(n_327)
);

AOI21xp5_ASAP7_75t_L g334 ( 
.A1(n_327),
.A2(n_330),
.B(n_260),
.Y(n_334)
);

MAJIxp5_ASAP7_75t_L g333 ( 
.A(n_329),
.B(n_332),
.C(n_280),
.Y(n_333)
);

NAND2xp5_ASAP7_75t_L g330 ( 
.A(n_324),
.B(n_308),
.Y(n_330)
);

XOR2xp5_ASAP7_75t_L g332 ( 
.A(n_326),
.B(n_293),
.Y(n_332)
);

INVxp67_ASAP7_75t_L g336 ( 
.A(n_333),
.Y(n_336)
);

NAND2xp5_ASAP7_75t_SL g335 ( 
.A(n_328),
.B(n_282),
.Y(n_335)
);

NOR3xp33_ASAP7_75t_L g337 ( 
.A(n_336),
.B(n_334),
.C(n_335),
.Y(n_337)
);

MAJIxp5_ASAP7_75t_L g338 ( 
.A(n_337),
.B(n_331),
.C(n_281),
.Y(n_338)
);

MAJIxp5_ASAP7_75t_L g339 ( 
.A(n_338),
.B(n_331),
.C(n_206),
.Y(n_339)
);

XNOR2xp5_ASAP7_75t_L g340 ( 
.A(n_339),
.B(n_213),
.Y(n_340)
);

NOR2xp33_ASAP7_75t_L g341 ( 
.A(n_340),
.B(n_14),
.Y(n_341)
);


endmodule