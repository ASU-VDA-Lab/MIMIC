module fake_jpeg_17568_n_161 (n_13, n_21, n_33, n_1, n_45, n_10, n_23, n_27, n_6, n_22, n_14, n_40, n_19, n_18, n_20, n_35, n_46, n_41, n_4, n_34, n_30, n_39, n_42, n_16, n_3, n_0, n_24, n_28, n_38, n_26, n_44, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_43, n_12, n_32, n_8, n_15, n_7, n_161);

input n_13;
input n_21;
input n_33;
input n_1;
input n_45;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_46;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_42;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_44;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_43;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_161;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_84;
wire n_59;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_155;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_57;
wire n_119;
wire n_69;
wire n_83;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_106;
wire n_111;
wire n_143;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_77;
wire n_136;
wire n_61;
wire n_139;
wire n_78;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_91;
wire n_54;
wire n_93;
wire n_138;
wire n_101;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_153;
wire n_135;
wire n_62;
wire n_120;
wire n_118;
wire n_100;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_8),
.Y(n_47)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_11),
.Y(n_48)
);

BUFx4f_ASAP7_75t_L g49 ( 
.A(n_2),
.Y(n_49)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_32),
.Y(n_50)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_20),
.Y(n_51)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_12),
.Y(n_52)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_38),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_11),
.Y(n_54)
);

INVx11_ASAP7_75t_L g55 ( 
.A(n_10),
.Y(n_55)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_9),
.Y(n_56)
);

CKINVDCx20_ASAP7_75t_R g57 ( 
.A(n_44),
.Y(n_57)
);

INVx8_ASAP7_75t_L g58 ( 
.A(n_10),
.Y(n_58)
);

INVx8_ASAP7_75t_L g59 ( 
.A(n_3),
.Y(n_59)
);

CKINVDCx20_ASAP7_75t_R g60 ( 
.A(n_24),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_15),
.Y(n_61)
);

CKINVDCx20_ASAP7_75t_R g62 ( 
.A(n_13),
.Y(n_62)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_45),
.Y(n_63)
);

INVx3_ASAP7_75t_L g64 ( 
.A(n_28),
.Y(n_64)
);

CKINVDCx16_ASAP7_75t_R g65 ( 
.A(n_14),
.Y(n_65)
);

INVx11_ASAP7_75t_L g66 ( 
.A(n_49),
.Y(n_66)
);

HB1xp67_ASAP7_75t_L g76 ( 
.A(n_66),
.Y(n_76)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_52),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_67),
.B(n_56),
.Y(n_83)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_61),
.Y(n_68)
);

BUFx6f_ASAP7_75t_L g75 ( 
.A(n_68),
.Y(n_75)
);

INVx3_ASAP7_75t_L g69 ( 
.A(n_49),
.Y(n_69)
);

INVx3_ASAP7_75t_L g81 ( 
.A(n_69),
.Y(n_81)
);

BUFx6f_ASAP7_75t_L g70 ( 
.A(n_61),
.Y(n_70)
);

BUFx6f_ASAP7_75t_L g82 ( 
.A(n_70),
.Y(n_82)
);

BUFx6f_ASAP7_75t_L g71 ( 
.A(n_49),
.Y(n_71)
);

BUFx6f_ASAP7_75t_L g90 ( 
.A(n_71),
.Y(n_90)
);

INVx6_ASAP7_75t_L g72 ( 
.A(n_54),
.Y(n_72)
);

INVx2_ASAP7_75t_L g77 ( 
.A(n_72),
.Y(n_77)
);

BUFx3_ASAP7_75t_L g73 ( 
.A(n_54),
.Y(n_73)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_73),
.Y(n_80)
);

INVx6_ASAP7_75t_L g74 ( 
.A(n_68),
.Y(n_74)
);

INVx2_ASAP7_75t_L g94 ( 
.A(n_74),
.Y(n_94)
);

INVx2_ASAP7_75t_L g78 ( 
.A(n_70),
.Y(n_78)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_78),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g79 ( 
.A(n_67),
.B(n_52),
.Y(n_79)
);

AND2x2_ASAP7_75t_L g100 ( 
.A(n_79),
.B(n_85),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_L g92 ( 
.A(n_83),
.B(n_87),
.Y(n_92)
);

INVx3_ASAP7_75t_L g84 ( 
.A(n_69),
.Y(n_84)
);

INVx3_ASAP7_75t_L g95 ( 
.A(n_84),
.Y(n_95)
);

AND2x2_ASAP7_75t_L g85 ( 
.A(n_66),
.B(n_47),
.Y(n_85)
);

INVx3_ASAP7_75t_L g86 ( 
.A(n_71),
.Y(n_86)
);

INVx3_ASAP7_75t_L g108 ( 
.A(n_86),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_73),
.B(n_56),
.Y(n_87)
);

INVx3_ASAP7_75t_L g88 ( 
.A(n_72),
.Y(n_88)
);

INVx3_ASAP7_75t_L g109 ( 
.A(n_88),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_67),
.B(n_48),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_SL g106 ( 
.A(n_89),
.B(n_91),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_67),
.B(n_50),
.Y(n_91)
);

AOI21xp5_ASAP7_75t_L g93 ( 
.A1(n_87),
.A2(n_64),
.B(n_50),
.Y(n_93)
);

OAI22xp5_ASAP7_75t_SL g121 ( 
.A1(n_93),
.A2(n_103),
.B1(n_104),
.B2(n_107),
.Y(n_121)
);

INVx5_ASAP7_75t_SL g97 ( 
.A(n_76),
.Y(n_97)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_97),
.Y(n_115)
);

CKINVDCx20_ASAP7_75t_R g98 ( 
.A(n_91),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g123 ( 
.A(n_98),
.B(n_99),
.Y(n_123)
);

CKINVDCx20_ASAP7_75t_R g99 ( 
.A(n_83),
.Y(n_99)
);

BUFx2_ASAP7_75t_L g101 ( 
.A(n_76),
.Y(n_101)
);

INVx3_ASAP7_75t_L g113 ( 
.A(n_101),
.Y(n_113)
);

HB1xp67_ASAP7_75t_L g102 ( 
.A(n_80),
.Y(n_102)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_102),
.Y(n_116)
);

AOI22xp33_ASAP7_75t_SL g103 ( 
.A1(n_77),
.A2(n_64),
.B1(n_55),
.B2(n_59),
.Y(n_103)
);

OA22x2_ASAP7_75t_L g104 ( 
.A1(n_90),
.A2(n_55),
.B1(n_58),
.B2(n_59),
.Y(n_104)
);

INVx2_ASAP7_75t_L g105 ( 
.A(n_75),
.Y(n_105)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_105),
.Y(n_119)
);

AOI22xp33_ASAP7_75t_SL g107 ( 
.A1(n_81),
.A2(n_58),
.B1(n_65),
.B2(n_62),
.Y(n_107)
);

INVx4_ASAP7_75t_L g110 ( 
.A(n_82),
.Y(n_110)
);

INVx2_ASAP7_75t_L g114 ( 
.A(n_110),
.Y(n_114)
);

AOI22xp33_ASAP7_75t_SL g111 ( 
.A1(n_74),
.A2(n_60),
.B1(n_57),
.B2(n_53),
.Y(n_111)
);

AOI22xp5_ASAP7_75t_L g122 ( 
.A1(n_111),
.A2(n_112),
.B1(n_0),
.B2(n_1),
.Y(n_122)
);

OA22x2_ASAP7_75t_SL g112 ( 
.A1(n_77),
.A2(n_51),
.B1(n_25),
.B2(n_46),
.Y(n_112)
);

INVx2_ASAP7_75t_L g117 ( 
.A(n_96),
.Y(n_117)
);

INVx2_ASAP7_75t_L g130 ( 
.A(n_117),
.Y(n_130)
);

AO22x2_ASAP7_75t_L g118 ( 
.A1(n_104),
.A2(n_22),
.B1(n_43),
.B2(n_42),
.Y(n_118)
);

AOI22xp5_ASAP7_75t_L g128 ( 
.A1(n_118),
.A2(n_120),
.B1(n_100),
.B2(n_3),
.Y(n_128)
);

AOI22xp33_ASAP7_75t_L g120 ( 
.A1(n_94),
.A2(n_63),
.B1(n_1),
.B2(n_2),
.Y(n_120)
);

OAI22xp5_ASAP7_75t_L g126 ( 
.A1(n_122),
.A2(n_92),
.B1(n_106),
.B2(n_103),
.Y(n_126)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_95),
.Y(n_124)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_124),
.Y(n_129)
);

INVx3_ASAP7_75t_L g125 ( 
.A(n_108),
.Y(n_125)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_125),
.Y(n_131)
);

AOI22xp33_ASAP7_75t_L g135 ( 
.A1(n_126),
.A2(n_118),
.B1(n_121),
.B2(n_109),
.Y(n_135)
);

AND2x2_ASAP7_75t_L g127 ( 
.A(n_123),
.B(n_112),
.Y(n_127)
);

XNOR2xp5_ASAP7_75t_L g134 ( 
.A(n_127),
.B(n_132),
.Y(n_134)
);

OAI22xp5_ASAP7_75t_SL g133 ( 
.A1(n_128),
.A2(n_120),
.B1(n_118),
.B2(n_100),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_L g132 ( 
.A(n_115),
.B(n_106),
.Y(n_132)
);

OAI22xp5_ASAP7_75t_L g141 ( 
.A1(n_133),
.A2(n_135),
.B1(n_136),
.B2(n_114),
.Y(n_141)
);

OA21x2_ASAP7_75t_L g136 ( 
.A1(n_128),
.A2(n_113),
.B(n_116),
.Y(n_136)
);

MAJIxp5_ASAP7_75t_L g137 ( 
.A(n_129),
.B(n_119),
.C(n_26),
.Y(n_137)
);

MAJIxp5_ASAP7_75t_L g142 ( 
.A(n_137),
.B(n_23),
.C(n_41),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_L g138 ( 
.A(n_136),
.B(n_131),
.Y(n_138)
);

CKINVDCx20_ASAP7_75t_R g146 ( 
.A(n_138),
.Y(n_146)
);

AOI21xp5_ASAP7_75t_L g139 ( 
.A1(n_134),
.A2(n_127),
.B(n_27),
.Y(n_139)
);

OAI22xp5_ASAP7_75t_SL g144 ( 
.A1(n_139),
.A2(n_140),
.B1(n_141),
.B2(n_130),
.Y(n_144)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_135),
.Y(n_140)
);

MAJIxp5_ASAP7_75t_L g147 ( 
.A(n_142),
.B(n_143),
.C(n_17),
.Y(n_147)
);

MAJx2_ASAP7_75t_L g143 ( 
.A(n_134),
.B(n_21),
.C(n_30),
.Y(n_143)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_144),
.Y(n_148)
);

AOI22xp5_ASAP7_75t_L g145 ( 
.A1(n_138),
.A2(n_130),
.B1(n_19),
.B2(n_29),
.Y(n_145)
);

MAJIxp5_ASAP7_75t_L g149 ( 
.A(n_145),
.B(n_147),
.C(n_18),
.Y(n_149)
);

XOR2xp5_ASAP7_75t_L g150 ( 
.A(n_149),
.B(n_147),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_L g151 ( 
.A(n_150),
.B(n_148),
.Y(n_151)
);

OAI22xp33_ASAP7_75t_SL g152 ( 
.A1(n_151),
.A2(n_146),
.B1(n_145),
.B2(n_31),
.Y(n_152)
);

AO21x1_ASAP7_75t_L g153 ( 
.A1(n_152),
.A2(n_16),
.B(n_40),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_L g154 ( 
.A(n_153),
.B(n_39),
.Y(n_154)
);

OAI21xp5_ASAP7_75t_SL g155 ( 
.A1(n_154),
.A2(n_37),
.B(n_36),
.Y(n_155)
);

OAI21xp5_ASAP7_75t_SL g156 ( 
.A1(n_155),
.A2(n_35),
.B(n_34),
.Y(n_156)
);

NOR2xp33_ASAP7_75t_L g157 ( 
.A(n_156),
.B(n_33),
.Y(n_157)
);

MAJIxp5_ASAP7_75t_L g158 ( 
.A(n_157),
.B(n_0),
.C(n_4),
.Y(n_158)
);

OAI321xp33_ASAP7_75t_L g159 ( 
.A1(n_158),
.A2(n_4),
.A3(n_5),
.B1(n_6),
.B2(n_7),
.C(n_8),
.Y(n_159)
);

OAI22xp5_ASAP7_75t_L g160 ( 
.A1(n_159),
.A2(n_5),
.B1(n_6),
.B2(n_7),
.Y(n_160)
);

BUFx24_ASAP7_75t_SL g161 ( 
.A(n_160),
.Y(n_161)
);


endmodule