module fake_jpeg_25278_n_250 (n_11, n_3, n_2, n_1, n_0, n_10, n_4, n_8, n_9, n_6, n_5, n_7, n_250);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_250;

wire n_159;
wire n_117;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_14;
wire n_152;
wire n_19;
wire n_182;
wire n_84;
wire n_59;
wire n_98;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_16;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_13;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_223;
wire n_234;
wire n_171;
wire n_119;
wire n_23;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_44;
wire n_24;
wire n_143;
wire n_202;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_102;
wire n_121;
wire n_99;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_170;
wire n_162;
wire n_12;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_216;
wire n_217;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_48;
wire n_35;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

CKINVDCx20_ASAP7_75t_R g12 ( 
.A(n_5),
.Y(n_12)
);

INVx1_ASAP7_75t_L g13 ( 
.A(n_11),
.Y(n_13)
);

INVx1_ASAP7_75t_L g14 ( 
.A(n_1),
.Y(n_14)
);

BUFx6f_ASAP7_75t_L g15 ( 
.A(n_2),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_9),
.Y(n_16)
);

INVx8_ASAP7_75t_L g17 ( 
.A(n_8),
.Y(n_17)
);

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_10),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_0),
.Y(n_19)
);

INVx2_ASAP7_75t_L g20 ( 
.A(n_4),
.Y(n_20)
);

INVx8_ASAP7_75t_L g21 ( 
.A(n_6),
.Y(n_21)
);

INVx3_ASAP7_75t_L g22 ( 
.A(n_8),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_3),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_4),
.Y(n_24)
);

NAND2xp5_ASAP7_75t_SL g25 ( 
.A(n_20),
.B(n_0),
.Y(n_25)
);

NOR2xp33_ASAP7_75t_L g34 ( 
.A(n_25),
.B(n_28),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_20),
.Y(n_26)
);

INVx2_ASAP7_75t_L g35 ( 
.A(n_26),
.Y(n_35)
);

BUFx4f_ASAP7_75t_L g27 ( 
.A(n_15),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_27),
.Y(n_39)
);

BUFx5_ASAP7_75t_L g28 ( 
.A(n_15),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_20),
.Y(n_29)
);

INVx2_ASAP7_75t_L g38 ( 
.A(n_29),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_L g30 ( 
.A(n_12),
.B(n_6),
.Y(n_30)
);

NOR2xp33_ASAP7_75t_L g42 ( 
.A(n_30),
.B(n_32),
.Y(n_42)
);

INVx11_ASAP7_75t_L g31 ( 
.A(n_15),
.Y(n_31)
);

INVx8_ASAP7_75t_L g37 ( 
.A(n_31),
.Y(n_37)
);

INVx3_ASAP7_75t_L g32 ( 
.A(n_18),
.Y(n_32)
);

INVx2_ASAP7_75t_SL g33 ( 
.A(n_15),
.Y(n_33)
);

INVx4_ASAP7_75t_SL g36 ( 
.A(n_33),
.Y(n_36)
);

CKINVDCx16_ASAP7_75t_R g40 ( 
.A(n_25),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_40),
.B(n_43),
.Y(n_56)
);

AOI22xp5_ASAP7_75t_L g41 ( 
.A1(n_32),
.A2(n_22),
.B1(n_17),
.B2(n_21),
.Y(n_41)
);

OAI22xp5_ASAP7_75t_L g55 ( 
.A1(n_41),
.A2(n_32),
.B1(n_33),
.B2(n_31),
.Y(n_55)
);

INVx3_ASAP7_75t_L g43 ( 
.A(n_29),
.Y(n_43)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_30),
.Y(n_44)
);

NAND2xp5_ASAP7_75t_L g49 ( 
.A(n_44),
.B(n_30),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_L g45 ( 
.A(n_34),
.B(n_25),
.Y(n_45)
);

NAND2xp5_ASAP7_75t_L g63 ( 
.A(n_45),
.B(n_52),
.Y(n_63)
);

INVx2_ASAP7_75t_L g46 ( 
.A(n_38),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_46),
.Y(n_64)
);

INVx4_ASAP7_75t_L g47 ( 
.A(n_39),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_47),
.B(n_51),
.Y(n_62)
);

INVx3_ASAP7_75t_L g48 ( 
.A(n_37),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_48),
.B(n_57),
.Y(n_78)
);

AND2x2_ASAP7_75t_L g72 ( 
.A(n_49),
.B(n_55),
.Y(n_72)
);

AOI22xp33_ASAP7_75t_SL g50 ( 
.A1(n_44),
.A2(n_17),
.B1(n_21),
.B2(n_22),
.Y(n_50)
);

AOI22xp33_ASAP7_75t_SL g65 ( 
.A1(n_50),
.A2(n_33),
.B1(n_36),
.B2(n_22),
.Y(n_65)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_42),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_L g52 ( 
.A(n_40),
.B(n_26),
.Y(n_52)
);

OR2x2_ASAP7_75t_L g53 ( 
.A(n_34),
.B(n_29),
.Y(n_53)
);

OR2x2_ASAP7_75t_L g75 ( 
.A(n_53),
.B(n_39),
.Y(n_75)
);

OAI22xp33_ASAP7_75t_SL g54 ( 
.A1(n_35),
.A2(n_32),
.B1(n_33),
.B2(n_31),
.Y(n_54)
);

OA22x2_ASAP7_75t_L g67 ( 
.A1(n_54),
.A2(n_36),
.B1(n_33),
.B2(n_43),
.Y(n_67)
);

INVx4_ASAP7_75t_L g57 ( 
.A(n_39),
.Y(n_57)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_38),
.Y(n_58)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_58),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_L g59 ( 
.A(n_42),
.B(n_26),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_L g71 ( 
.A(n_59),
.B(n_29),
.Y(n_71)
);

INVx2_ASAP7_75t_SL g60 ( 
.A(n_39),
.Y(n_60)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_60),
.Y(n_66)
);

AOI22xp33_ASAP7_75t_L g84 ( 
.A1(n_65),
.A2(n_69),
.B1(n_36),
.B2(n_60),
.Y(n_84)
);

AND2x2_ASAP7_75t_L g85 ( 
.A(n_67),
.B(n_27),
.Y(n_85)
);

AOI22xp33_ASAP7_75t_SL g68 ( 
.A1(n_51),
.A2(n_12),
.B1(n_16),
.B2(n_21),
.Y(n_68)
);

INVxp67_ASAP7_75t_L g80 ( 
.A(n_68),
.Y(n_80)
);

AOI22xp33_ASAP7_75t_SL g69 ( 
.A1(n_48),
.A2(n_12),
.B1(n_16),
.B2(n_17),
.Y(n_69)
);

CKINVDCx20_ASAP7_75t_R g70 ( 
.A(n_59),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_70),
.B(n_73),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_L g87 ( 
.A(n_71),
.B(n_76),
.Y(n_87)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_56),
.Y(n_73)
);

FAx1_ASAP7_75t_SL g74 ( 
.A(n_45),
.B(n_52),
.CI(n_56),
.CON(n_74),
.SN(n_74)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_74),
.B(n_77),
.Y(n_90)
);

OR2x2_ASAP7_75t_L g82 ( 
.A(n_75),
.B(n_28),
.Y(n_82)
);

OAI21xp5_ASAP7_75t_SL g76 ( 
.A1(n_53),
.A2(n_41),
.B(n_14),
.Y(n_76)
);

INVxp67_ASAP7_75t_L g77 ( 
.A(n_50),
.Y(n_77)
);

OAI22xp5_ASAP7_75t_SL g79 ( 
.A1(n_75),
.A2(n_53),
.B1(n_41),
.B2(n_55),
.Y(n_79)
);

OAI22xp5_ASAP7_75t_SL g99 ( 
.A1(n_79),
.A2(n_81),
.B1(n_83),
.B2(n_88),
.Y(n_99)
);

AOI22xp5_ASAP7_75t_L g81 ( 
.A1(n_72),
.A2(n_53),
.B1(n_54),
.B2(n_45),
.Y(n_81)
);

OAI21xp5_ASAP7_75t_L g110 ( 
.A1(n_82),
.A2(n_85),
.B(n_76),
.Y(n_110)
);

OAI22xp5_ASAP7_75t_SL g83 ( 
.A1(n_75),
.A2(n_49),
.B1(n_35),
.B2(n_33),
.Y(n_83)
);

INVxp67_ASAP7_75t_L g109 ( 
.A(n_84),
.Y(n_109)
);

OAI22xp5_ASAP7_75t_SL g88 ( 
.A1(n_70),
.A2(n_35),
.B1(n_43),
.B2(n_31),
.Y(n_88)
);

OAI22xp5_ASAP7_75t_SL g89 ( 
.A1(n_63),
.A2(n_31),
.B1(n_58),
.B2(n_46),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g103 ( 
.A(n_89),
.B(n_67),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_SL g91 ( 
.A(n_63),
.B(n_16),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_SL g106 ( 
.A(n_91),
.B(n_92),
.Y(n_106)
);

AND2x6_ASAP7_75t_L g92 ( 
.A(n_74),
.B(n_11),
.Y(n_92)
);

INVx13_ASAP7_75t_L g93 ( 
.A(n_64),
.Y(n_93)
);

INVx4_ASAP7_75t_L g113 ( 
.A(n_93),
.Y(n_113)
);

INVx11_ASAP7_75t_SL g94 ( 
.A(n_78),
.Y(n_94)
);

INVx2_ASAP7_75t_L g108 ( 
.A(n_94),
.Y(n_108)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_78),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_SL g111 ( 
.A(n_95),
.B(n_62),
.Y(n_111)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_88),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_SL g116 ( 
.A(n_96),
.B(n_111),
.Y(n_116)
);

CKINVDCx20_ASAP7_75t_R g97 ( 
.A(n_86),
.Y(n_97)
);

CKINVDCx20_ASAP7_75t_R g115 ( 
.A(n_97),
.Y(n_115)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_89),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_SL g130 ( 
.A(n_98),
.B(n_107),
.Y(n_130)
);

XNOR2xp5_ASAP7_75t_L g100 ( 
.A(n_90),
.B(n_74),
.Y(n_100)
);

MAJIxp5_ASAP7_75t_L g114 ( 
.A(n_100),
.B(n_112),
.C(n_87),
.Y(n_114)
);

AND2x2_ASAP7_75t_L g101 ( 
.A(n_90),
.B(n_83),
.Y(n_101)
);

OAI21xp5_ASAP7_75t_SL g129 ( 
.A1(n_101),
.A2(n_104),
.B(n_105),
.Y(n_129)
);

CKINVDCx20_ASAP7_75t_R g102 ( 
.A(n_86),
.Y(n_102)
);

CKINVDCx20_ASAP7_75t_R g120 ( 
.A(n_102),
.Y(n_120)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_103),
.Y(n_125)
);

AOI22xp33_ASAP7_75t_SL g104 ( 
.A1(n_95),
.A2(n_73),
.B1(n_48),
.B2(n_57),
.Y(n_104)
);

AOI22xp33_ASAP7_75t_SL g105 ( 
.A1(n_80),
.A2(n_93),
.B1(n_47),
.B2(n_57),
.Y(n_105)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_85),
.Y(n_107)
);

AOI21xp5_ASAP7_75t_SL g123 ( 
.A1(n_110),
.A2(n_82),
.B(n_72),
.Y(n_123)
);

XNOR2xp5_ASAP7_75t_L g112 ( 
.A(n_87),
.B(n_74),
.Y(n_112)
);

XNOR2xp5_ASAP7_75t_L g136 ( 
.A(n_114),
.B(n_110),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_108),
.B(n_62),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_SL g148 ( 
.A(n_117),
.B(n_119),
.Y(n_148)
);

OAI22xp5_ASAP7_75t_SL g118 ( 
.A1(n_98),
.A2(n_81),
.B1(n_92),
.B2(n_79),
.Y(n_118)
);

AOI22xp5_ASAP7_75t_L g154 ( 
.A1(n_118),
.A2(n_121),
.B1(n_122),
.B2(n_125),
.Y(n_154)
);

NOR2xp33_ASAP7_75t_L g119 ( 
.A(n_108),
.B(n_91),
.Y(n_119)
);

OAI22xp5_ASAP7_75t_L g121 ( 
.A1(n_103),
.A2(n_92),
.B1(n_85),
.B2(n_71),
.Y(n_121)
);

OAI22xp5_ASAP7_75t_SL g122 ( 
.A1(n_109),
.A2(n_85),
.B1(n_82),
.B2(n_72),
.Y(n_122)
);

OAI21xp5_ASAP7_75t_SL g138 ( 
.A1(n_123),
.A2(n_101),
.B(n_67),
.Y(n_138)
);

AND2x6_ASAP7_75t_L g124 ( 
.A(n_106),
.B(n_67),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_L g142 ( 
.A(n_124),
.B(n_133),
.Y(n_142)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_99),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_L g135 ( 
.A(n_126),
.B(n_107),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_112),
.B(n_61),
.Y(n_127)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_127),
.Y(n_156)
);

MAJIxp5_ASAP7_75t_L g128 ( 
.A(n_100),
.B(n_61),
.C(n_64),
.Y(n_128)
);

MAJIxp5_ASAP7_75t_L g137 ( 
.A(n_128),
.B(n_122),
.C(n_115),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_L g131 ( 
.A(n_99),
.B(n_64),
.Y(n_131)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_131),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_L g132 ( 
.A(n_113),
.B(n_93),
.Y(n_132)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_132),
.Y(n_144)
);

INVx13_ASAP7_75t_L g133 ( 
.A(n_113),
.Y(n_133)
);

INVx3_ASAP7_75t_L g134 ( 
.A(n_109),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_L g155 ( 
.A(n_134),
.B(n_47),
.Y(n_155)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_135),
.Y(n_171)
);

XNOR2xp5_ASAP7_75t_L g163 ( 
.A(n_136),
.B(n_140),
.Y(n_163)
);

MAJIxp5_ASAP7_75t_L g159 ( 
.A(n_137),
.B(n_128),
.C(n_121),
.Y(n_159)
);

AO21x1_ASAP7_75t_L g161 ( 
.A1(n_138),
.A2(n_66),
.B(n_28),
.Y(n_161)
);

INVx2_ASAP7_75t_L g139 ( 
.A(n_133),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_L g162 ( 
.A(n_139),
.B(n_145),
.Y(n_162)
);

XOR2xp5_ASAP7_75t_L g140 ( 
.A(n_114),
.B(n_101),
.Y(n_140)
);

A2O1A1Ixp33_ASAP7_75t_L g143 ( 
.A1(n_126),
.A2(n_13),
.B(n_24),
.C(n_23),
.Y(n_143)
);

OAI21xp5_ASAP7_75t_L g158 ( 
.A1(n_143),
.A2(n_153),
.B(n_123),
.Y(n_158)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_130),
.Y(n_145)
);

CKINVDCx20_ASAP7_75t_R g146 ( 
.A(n_115),
.Y(n_146)
);

CKINVDCx20_ASAP7_75t_R g165 ( 
.A(n_146),
.Y(n_165)
);

NOR4xp25_ASAP7_75t_L g147 ( 
.A(n_120),
.B(n_17),
.C(n_21),
.D(n_23),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_L g166 ( 
.A(n_147),
.B(n_149),
.Y(n_166)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_130),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_L g150 ( 
.A(n_120),
.B(n_58),
.Y(n_150)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_150),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_L g151 ( 
.A(n_116),
.B(n_46),
.Y(n_151)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_151),
.Y(n_175)
);

NOR2xp33_ASAP7_75t_L g152 ( 
.A(n_118),
.B(n_18),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_L g168 ( 
.A(n_152),
.B(n_155),
.Y(n_168)
);

AND2x2_ASAP7_75t_L g153 ( 
.A(n_129),
.B(n_67),
.Y(n_153)
);

OAI22xp5_ASAP7_75t_SL g169 ( 
.A1(n_154),
.A2(n_60),
.B1(n_36),
.B2(n_37),
.Y(n_169)
);

AOI22xp5_ASAP7_75t_SL g157 ( 
.A1(n_153),
.A2(n_134),
.B1(n_129),
.B2(n_125),
.Y(n_157)
);

OAI22xp5_ASAP7_75t_SL g187 ( 
.A1(n_157),
.A2(n_167),
.B1(n_24),
.B2(n_19),
.Y(n_187)
);

AO21x1_ASAP7_75t_L g177 ( 
.A1(n_158),
.A2(n_148),
.B(n_151),
.Y(n_177)
);

XOR2xp5_ASAP7_75t_L g185 ( 
.A(n_159),
.B(n_28),
.Y(n_185)
);

OAI22xp5_ASAP7_75t_L g160 ( 
.A1(n_142),
.A2(n_124),
.B1(n_127),
.B2(n_66),
.Y(n_160)
);

AOI22xp5_ASAP7_75t_L g181 ( 
.A1(n_160),
.A2(n_164),
.B1(n_169),
.B2(n_60),
.Y(n_181)
);

AOI21xp5_ASAP7_75t_L g176 ( 
.A1(n_161),
.A2(n_150),
.B(n_143),
.Y(n_176)
);

OAI22xp5_ASAP7_75t_SL g164 ( 
.A1(n_154),
.A2(n_135),
.B1(n_137),
.B2(n_141),
.Y(n_164)
);

AOI22xp5_ASAP7_75t_L g167 ( 
.A1(n_153),
.A2(n_156),
.B1(n_138),
.B2(n_144),
.Y(n_167)
);

XNOR2xp5_ASAP7_75t_L g170 ( 
.A(n_136),
.B(n_13),
.Y(n_170)
);

XNOR2xp5_ASAP7_75t_L g182 ( 
.A(n_170),
.B(n_14),
.Y(n_182)
);

MAJIxp5_ASAP7_75t_L g172 ( 
.A(n_140),
.B(n_29),
.C(n_26),
.Y(n_172)
);

MAJIxp5_ASAP7_75t_L g180 ( 
.A(n_172),
.B(n_174),
.C(n_37),
.Y(n_180)
);

MAJIxp5_ASAP7_75t_L g174 ( 
.A(n_156),
.B(n_29),
.C(n_26),
.Y(n_174)
);

HAxp5_ASAP7_75t_SL g199 ( 
.A(n_176),
.B(n_161),
.CON(n_199),
.SN(n_199)
);

AOI21xp5_ASAP7_75t_L g195 ( 
.A1(n_177),
.A2(n_178),
.B(n_183),
.Y(n_195)
);

OAI21xp5_ASAP7_75t_L g178 ( 
.A1(n_166),
.A2(n_139),
.B(n_13),
.Y(n_178)
);

INVx2_ASAP7_75t_SL g179 ( 
.A(n_165),
.Y(n_179)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_179),
.Y(n_196)
);

MAJIxp5_ASAP7_75t_L g198 ( 
.A(n_180),
.B(n_190),
.C(n_172),
.Y(n_198)
);

XOR2xp5_ASAP7_75t_L g201 ( 
.A(n_181),
.B(n_185),
.Y(n_201)
);

XNOR2xp5_ASAP7_75t_SL g202 ( 
.A(n_182),
.B(n_187),
.Y(n_202)
);

XNOR2xp5_ASAP7_75t_L g183 ( 
.A(n_159),
.B(n_14),
.Y(n_183)
);

AOI22xp5_ASAP7_75t_L g184 ( 
.A1(n_164),
.A2(n_24),
.B1(n_23),
.B2(n_18),
.Y(n_184)
);

BUFx2_ASAP7_75t_L g200 ( 
.A(n_184),
.Y(n_200)
);

HB1xp67_ASAP7_75t_L g186 ( 
.A(n_162),
.Y(n_186)
);

CKINVDCx20_ASAP7_75t_R g193 ( 
.A(n_186),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_L g188 ( 
.A(n_171),
.B(n_7),
.Y(n_188)
);

CKINVDCx20_ASAP7_75t_R g194 ( 
.A(n_188),
.Y(n_194)
);

OAI22xp5_ASAP7_75t_SL g189 ( 
.A1(n_167),
.A2(n_18),
.B1(n_27),
.B2(n_7),
.Y(n_189)
);

INVx13_ASAP7_75t_L g197 ( 
.A(n_189),
.Y(n_197)
);

XNOR2xp5_ASAP7_75t_L g190 ( 
.A(n_163),
.B(n_7),
.Y(n_190)
);

OAI22xp5_ASAP7_75t_L g191 ( 
.A1(n_168),
.A2(n_6),
.B1(n_11),
.B2(n_10),
.Y(n_191)
);

CKINVDCx20_ASAP7_75t_R g204 ( 
.A(n_191),
.Y(n_204)
);

XNOR2x1_ASAP7_75t_L g192 ( 
.A(n_163),
.B(n_157),
.Y(n_192)
);

XNOR2xp5_ASAP7_75t_SL g205 ( 
.A(n_192),
.B(n_158),
.Y(n_205)
);

NOR2xp33_ASAP7_75t_L g209 ( 
.A(n_198),
.B(n_180),
.Y(n_209)
);

A2O1A1Ixp33_ASAP7_75t_L g211 ( 
.A1(n_199),
.A2(n_190),
.B(n_8),
.C(n_9),
.Y(n_211)
);

MAJIxp5_ASAP7_75t_L g203 ( 
.A(n_185),
.B(n_173),
.C(n_174),
.Y(n_203)
);

MAJIxp5_ASAP7_75t_L g208 ( 
.A(n_203),
.B(n_198),
.C(n_196),
.Y(n_208)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_205),
.Y(n_207)
);

AO21x1_ASAP7_75t_L g206 ( 
.A1(n_177),
.A2(n_175),
.B(n_170),
.Y(n_206)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_206),
.Y(n_214)
);

MAJIxp5_ASAP7_75t_L g226 ( 
.A(n_208),
.B(n_215),
.C(n_216),
.Y(n_226)
);

NAND2xp5_ASAP7_75t_L g224 ( 
.A(n_209),
.B(n_210),
.Y(n_224)
);

OAI22xp5_ASAP7_75t_SL g210 ( 
.A1(n_197),
.A2(n_192),
.B1(n_179),
.B2(n_186),
.Y(n_210)
);

OAI21xp5_ASAP7_75t_L g220 ( 
.A1(n_211),
.A2(n_213),
.B(n_194),
.Y(n_220)
);

NAND2xp5_ASAP7_75t_L g212 ( 
.A(n_193),
.B(n_5),
.Y(n_212)
);

NOR2xp33_ASAP7_75t_L g219 ( 
.A(n_212),
.B(n_217),
.Y(n_219)
);

OAI21xp5_ASAP7_75t_SL g213 ( 
.A1(n_195),
.A2(n_5),
.B(n_10),
.Y(n_213)
);

MAJIxp5_ASAP7_75t_L g215 ( 
.A(n_203),
.B(n_19),
.C(n_27),
.Y(n_215)
);

MAJIxp5_ASAP7_75t_L g216 ( 
.A(n_201),
.B(n_19),
.C(n_27),
.Y(n_216)
);

CKINVDCx16_ASAP7_75t_R g217 ( 
.A(n_200),
.Y(n_217)
);

INVxp67_ASAP7_75t_L g218 ( 
.A(n_208),
.Y(n_218)
);

NAND2xp5_ASAP7_75t_L g235 ( 
.A(n_218),
.B(n_227),
.Y(n_235)
);

NAND2xp5_ASAP7_75t_SL g229 ( 
.A(n_220),
.B(n_221),
.Y(n_229)
);

XNOR2xp5_ASAP7_75t_L g221 ( 
.A(n_215),
.B(n_201),
.Y(n_221)
);

OAI22xp5_ASAP7_75t_SL g222 ( 
.A1(n_214),
.A2(n_197),
.B1(n_204),
.B2(n_206),
.Y(n_222)
);

NOR2xp33_ASAP7_75t_L g228 ( 
.A(n_222),
.B(n_223),
.Y(n_228)
);

XOR2xp5_ASAP7_75t_L g223 ( 
.A(n_216),
.B(n_205),
.Y(n_223)
);

XNOR2xp5_ASAP7_75t_L g225 ( 
.A(n_207),
.B(n_202),
.Y(n_225)
);

AND2x2_ASAP7_75t_SL g234 ( 
.A(n_225),
.B(n_0),
.Y(n_234)
);

XOR2xp5_ASAP7_75t_L g227 ( 
.A(n_211),
.B(n_202),
.Y(n_227)
);

NOR2x1_ASAP7_75t_L g230 ( 
.A(n_218),
.B(n_199),
.Y(n_230)
);

HB1xp67_ASAP7_75t_L g239 ( 
.A(n_230),
.Y(n_239)
);

INVx11_ASAP7_75t_L g231 ( 
.A(n_219),
.Y(n_231)
);

XOR2xp5_ASAP7_75t_L g237 ( 
.A(n_231),
.B(n_0),
.Y(n_237)
);

NOR2xp67_ASAP7_75t_L g232 ( 
.A(n_227),
.B(n_200),
.Y(n_232)
);

OAI21xp5_ASAP7_75t_L g236 ( 
.A1(n_232),
.A2(n_226),
.B(n_223),
.Y(n_236)
);

OAI22xp5_ASAP7_75t_L g233 ( 
.A1(n_224),
.A2(n_27),
.B1(n_19),
.B2(n_9),
.Y(n_233)
);

MAJIxp5_ASAP7_75t_L g240 ( 
.A(n_233),
.B(n_234),
.C(n_1),
.Y(n_240)
);

AOI21xp5_ASAP7_75t_L g243 ( 
.A1(n_236),
.A2(n_229),
.B(n_2),
.Y(n_243)
);

MAJIxp5_ASAP7_75t_L g242 ( 
.A(n_237),
.B(n_238),
.C(n_235),
.Y(n_242)
);

XOR2xp5_ASAP7_75t_L g238 ( 
.A(n_235),
.B(n_27),
.Y(n_238)
);

OR2x2_ASAP7_75t_L g241 ( 
.A(n_240),
.B(n_228),
.Y(n_241)
);

NAND2xp5_ASAP7_75t_L g245 ( 
.A(n_241),
.B(n_242),
.Y(n_245)
);

AOI31xp67_ASAP7_75t_SL g244 ( 
.A1(n_243),
.A2(n_239),
.A3(n_2),
.B(n_3),
.Y(n_244)
);

MAJx2_ASAP7_75t_L g246 ( 
.A(n_244),
.B(n_1),
.C(n_2),
.Y(n_246)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_246),
.Y(n_247)
);

AOI31xp33_ASAP7_75t_L g248 ( 
.A1(n_247),
.A2(n_245),
.A3(n_3),
.B(n_4),
.Y(n_248)
);

XNOR2xp5_ASAP7_75t_L g249 ( 
.A(n_248),
.B(n_1),
.Y(n_249)
);

AOI21xp5_ASAP7_75t_L g250 ( 
.A1(n_249),
.A2(n_3),
.B(n_4),
.Y(n_250)
);


endmodule