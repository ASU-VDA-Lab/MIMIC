module fake_jpeg_22402_n_187 (n_13, n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_187);

input n_13;
input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_187;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_14;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_175;
wire n_21;
wire n_57;
wire n_171;
wire n_119;
wire n_23;
wire n_69;
wire n_27;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_186;
wire n_24;
wire n_44;
wire n_143;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_177;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_128;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_161;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_176;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_36;
wire n_62;
wire n_167;
wire n_174;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_140;
wire n_96;

INVx1_ASAP7_75t_L g14 ( 
.A(n_13),
.Y(n_14)
);

BUFx6f_ASAP7_75t_L g15 ( 
.A(n_2),
.Y(n_15)
);

BUFx12f_ASAP7_75t_L g16 ( 
.A(n_11),
.Y(n_16)
);

BUFx6f_ASAP7_75t_L g17 ( 
.A(n_0),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_6),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_13),
.Y(n_19)
);

INVx11_ASAP7_75t_L g20 ( 
.A(n_4),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_2),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_11),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_1),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_6),
.Y(n_24)
);

INVx3_ASAP7_75t_L g25 ( 
.A(n_12),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_1),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_11),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_16),
.Y(n_28)
);

INVx6_ASAP7_75t_L g51 ( 
.A(n_28),
.Y(n_51)
);

BUFx3_ASAP7_75t_L g29 ( 
.A(n_16),
.Y(n_29)
);

BUFx2_ASAP7_75t_L g45 ( 
.A(n_29),
.Y(n_45)
);

INVx8_ASAP7_75t_L g30 ( 
.A(n_15),
.Y(n_30)
);

AOI22xp33_ASAP7_75t_SL g54 ( 
.A1(n_30),
.A2(n_35),
.B1(n_20),
.B2(n_25),
.Y(n_54)
);

BUFx3_ASAP7_75t_L g31 ( 
.A(n_16),
.Y(n_31)
);

INVx4_ASAP7_75t_L g44 ( 
.A(n_31),
.Y(n_44)
);

NAND2xp5_ASAP7_75t_L g32 ( 
.A(n_21),
.B(n_0),
.Y(n_32)
);

NOR2xp33_ASAP7_75t_L g41 ( 
.A(n_32),
.B(n_36),
.Y(n_41)
);

NAND2xp5_ASAP7_75t_SL g33 ( 
.A(n_21),
.B(n_0),
.Y(n_33)
);

NAND2xp33_ASAP7_75t_SL g42 ( 
.A(n_33),
.B(n_20),
.Y(n_42)
);

INVx6_ASAP7_75t_L g34 ( 
.A(n_15),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_34),
.Y(n_53)
);

INVx6_ASAP7_75t_L g35 ( 
.A(n_15),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_16),
.Y(n_36)
);

INVx5_ASAP7_75t_L g37 ( 
.A(n_16),
.Y(n_37)
);

INVx4_ASAP7_75t_L g52 ( 
.A(n_37),
.Y(n_52)
);

OA22x2_ASAP7_75t_SL g38 ( 
.A1(n_29),
.A2(n_16),
.B1(n_27),
.B2(n_15),
.Y(n_38)
);

OA22x2_ASAP7_75t_L g62 ( 
.A1(n_38),
.A2(n_37),
.B1(n_28),
.B2(n_27),
.Y(n_62)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_32),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_39),
.B(n_40),
.Y(n_58)
);

INVx3_ASAP7_75t_L g40 ( 
.A(n_29),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_SL g65 ( 
.A(n_42),
.B(n_43),
.Y(n_65)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_33),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g46 ( 
.A(n_36),
.B(n_19),
.Y(n_46)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_46),
.Y(n_61)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_31),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_SL g70 ( 
.A(n_47),
.B(n_49),
.Y(n_70)
);

OAI22xp5_ASAP7_75t_L g48 ( 
.A1(n_34),
.A2(n_25),
.B1(n_20),
.B2(n_21),
.Y(n_48)
);

AOI22xp5_ASAP7_75t_L g60 ( 
.A1(n_48),
.A2(n_35),
.B1(n_30),
.B2(n_14),
.Y(n_60)
);

OR2x2_ASAP7_75t_L g49 ( 
.A(n_31),
.B(n_24),
.Y(n_49)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_34),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_50),
.B(n_14),
.Y(n_67)
);

CKINVDCx16_ASAP7_75t_R g66 ( 
.A(n_54),
.Y(n_66)
);

INVx3_ASAP7_75t_L g55 ( 
.A(n_48),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_55),
.B(n_68),
.Y(n_83)
);

BUFx2_ASAP7_75t_L g56 ( 
.A(n_53),
.Y(n_56)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_56),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_L g57 ( 
.A(n_39),
.B(n_28),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_57),
.B(n_69),
.Y(n_89)
);

OAI22xp5_ASAP7_75t_L g59 ( 
.A1(n_38),
.A2(n_35),
.B1(n_30),
.B2(n_25),
.Y(n_59)
);

OAI22xp5_ASAP7_75t_SL g72 ( 
.A1(n_59),
.A2(n_60),
.B1(n_64),
.B2(n_50),
.Y(n_72)
);

NAND2xp33_ASAP7_75t_SL g74 ( 
.A(n_62),
.B(n_53),
.Y(n_74)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_41),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_SL g82 ( 
.A(n_63),
.B(n_71),
.Y(n_82)
);

OAI22xp33_ASAP7_75t_SL g64 ( 
.A1(n_38),
.A2(n_37),
.B1(n_14),
.B2(n_19),
.Y(n_64)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_67),
.Y(n_77)
);

INVx2_ASAP7_75t_L g68 ( 
.A(n_38),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_L g69 ( 
.A(n_43),
.B(n_27),
.Y(n_69)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_45),
.Y(n_71)
);

AOI22xp5_ASAP7_75t_L g106 ( 
.A1(n_72),
.A2(n_73),
.B1(n_62),
.B2(n_40),
.Y(n_106)
);

OAI22xp5_ASAP7_75t_SL g73 ( 
.A1(n_55),
.A2(n_52),
.B1(n_42),
.B2(n_51),
.Y(n_73)
);

AOI22xp33_ASAP7_75t_L g104 ( 
.A1(n_74),
.A2(n_81),
.B1(n_88),
.B2(n_51),
.Y(n_104)
);

INVxp67_ASAP7_75t_L g76 ( 
.A(n_67),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_76),
.B(n_78),
.Y(n_96)
);

INVx4_ASAP7_75t_L g78 ( 
.A(n_71),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_SL g79 ( 
.A(n_65),
.B(n_49),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_SL g91 ( 
.A(n_79),
.B(n_84),
.Y(n_91)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_58),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_80),
.B(n_90),
.Y(n_98)
);

AND2x2_ASAP7_75t_L g81 ( 
.A(n_57),
.B(n_47),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_SL g84 ( 
.A(n_58),
.B(n_24),
.Y(n_84)
);

CKINVDCx14_ASAP7_75t_R g85 ( 
.A(n_70),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_85),
.B(n_86),
.Y(n_101)
);

INVx3_ASAP7_75t_L g86 ( 
.A(n_56),
.Y(n_86)
);

CKINVDCx20_ASAP7_75t_R g87 ( 
.A(n_69),
.Y(n_87)
);

CKINVDCx20_ASAP7_75t_R g93 ( 
.A(n_87),
.Y(n_93)
);

AND2x2_ASAP7_75t_L g88 ( 
.A(n_65),
.B(n_49),
.Y(n_88)
);

INVx2_ASAP7_75t_L g90 ( 
.A(n_56),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_L g92 ( 
.A(n_89),
.B(n_70),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_L g115 ( 
.A(n_92),
.B(n_102),
.Y(n_115)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_78),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_SL g117 ( 
.A(n_94),
.B(n_95),
.Y(n_117)
);

INVxp67_ASAP7_75t_L g95 ( 
.A(n_82),
.Y(n_95)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_89),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_SL g119 ( 
.A(n_97),
.B(n_77),
.Y(n_119)
);

CKINVDCx20_ASAP7_75t_R g99 ( 
.A(n_81),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g112 ( 
.A(n_99),
.B(n_76),
.Y(n_112)
);

O2A1O1Ixp33_ASAP7_75t_L g100 ( 
.A1(n_73),
.A2(n_59),
.B(n_62),
.C(n_68),
.Y(n_100)
);

AOI22xp5_ASAP7_75t_L g110 ( 
.A1(n_100),
.A2(n_106),
.B1(n_107),
.B2(n_86),
.Y(n_110)
);

OAI32xp33_ASAP7_75t_L g102 ( 
.A1(n_83),
.A2(n_62),
.A3(n_63),
.B1(n_60),
.B2(n_66),
.Y(n_102)
);

AOI22xp33_ASAP7_75t_SL g103 ( 
.A1(n_80),
.A2(n_66),
.B1(n_52),
.B2(n_51),
.Y(n_103)
);

AO21x1_ASAP7_75t_L g120 ( 
.A1(n_103),
.A2(n_104),
.B(n_99),
.Y(n_120)
);

XNOR2xp5_ASAP7_75t_L g105 ( 
.A(n_88),
.B(n_62),
.Y(n_105)
);

MAJIxp5_ASAP7_75t_L g116 ( 
.A(n_105),
.B(n_81),
.C(n_88),
.Y(n_116)
);

AOI22xp5_ASAP7_75t_L g107 ( 
.A1(n_72),
.A2(n_44),
.B1(n_53),
.B2(n_18),
.Y(n_107)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_98),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_L g135 ( 
.A(n_108),
.B(n_109),
.Y(n_135)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_98),
.Y(n_109)
);

OAI22xp5_ASAP7_75t_L g138 ( 
.A1(n_110),
.A2(n_111),
.B1(n_124),
.B2(n_121),
.Y(n_138)
);

AOI22xp5_ASAP7_75t_L g111 ( 
.A1(n_100),
.A2(n_74),
.B1(n_87),
.B2(n_79),
.Y(n_111)
);

AOI21xp5_ASAP7_75t_L g126 ( 
.A1(n_112),
.A2(n_120),
.B(n_123),
.Y(n_126)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_96),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_SL g132 ( 
.A(n_113),
.B(n_114),
.Y(n_132)
);

CKINVDCx16_ASAP7_75t_R g114 ( 
.A(n_101),
.Y(n_114)
);

XNOR2xp5_ASAP7_75t_L g125 ( 
.A(n_116),
.B(n_105),
.Y(n_125)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_92),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_118),
.B(n_121),
.Y(n_128)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_119),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g121 ( 
.A(n_97),
.B(n_77),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_L g122 ( 
.A(n_93),
.B(n_75),
.Y(n_122)
);

CKINVDCx16_ASAP7_75t_R g137 ( 
.A(n_122),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_L g123 ( 
.A(n_95),
.B(n_61),
.Y(n_123)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_107),
.Y(n_124)
);

XOR2xp5_ASAP7_75t_L g143 ( 
.A(n_125),
.B(n_127),
.Y(n_143)
);

XNOR2xp5_ASAP7_75t_L g127 ( 
.A(n_116),
.B(n_106),
.Y(n_127)
);

XOR2xp5_ASAP7_75t_L g129 ( 
.A(n_115),
.B(n_102),
.Y(n_129)
);

MAJIxp5_ASAP7_75t_L g139 ( 
.A(n_129),
.B(n_136),
.C(n_122),
.Y(n_139)
);

OAI22xp5_ASAP7_75t_SL g130 ( 
.A1(n_115),
.A2(n_93),
.B1(n_91),
.B2(n_75),
.Y(n_130)
);

OAI22xp5_ASAP7_75t_SL g149 ( 
.A1(n_130),
.A2(n_134),
.B1(n_26),
.B2(n_23),
.Y(n_149)
);

AOI21xp5_ASAP7_75t_SL g133 ( 
.A1(n_118),
.A2(n_91),
.B(n_94),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_SL g147 ( 
.A(n_133),
.B(n_124),
.Y(n_147)
);

OAI22xp5_ASAP7_75t_SL g134 ( 
.A1(n_110),
.A2(n_90),
.B1(n_44),
.B2(n_61),
.Y(n_134)
);

XOR2xp5_ASAP7_75t_L g136 ( 
.A(n_111),
.B(n_45),
.Y(n_136)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_138),
.Y(n_144)
);

MAJIxp5_ASAP7_75t_L g154 ( 
.A(n_139),
.B(n_142),
.C(n_145),
.Y(n_154)
);

XOR2x2_ASAP7_75t_L g140 ( 
.A(n_136),
.B(n_120),
.Y(n_140)
);

OAI21xp5_ASAP7_75t_SL g151 ( 
.A1(n_140),
.A2(n_146),
.B(n_45),
.Y(n_151)
);

INVxp33_ASAP7_75t_SL g141 ( 
.A(n_132),
.Y(n_141)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_141),
.Y(n_158)
);

OAI322xp33_ASAP7_75t_L g142 ( 
.A1(n_133),
.A2(n_120),
.A3(n_117),
.B1(n_114),
.B2(n_113),
.C1(n_109),
.C2(n_108),
.Y(n_142)
);

OAI322xp33_ASAP7_75t_L g145 ( 
.A1(n_125),
.A2(n_137),
.A3(n_128),
.B1(n_135),
.B2(n_130),
.C1(n_127),
.C2(n_126),
.Y(n_145)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_134),
.Y(n_146)
);

AOI22xp5_ASAP7_75t_L g152 ( 
.A1(n_147),
.A2(n_149),
.B1(n_26),
.B2(n_23),
.Y(n_152)
);

CKINVDCx5p33_ASAP7_75t_R g148 ( 
.A(n_131),
.Y(n_148)
);

NOR2xp33_ASAP7_75t_L g156 ( 
.A(n_148),
.B(n_1),
.Y(n_156)
);

HB1xp67_ASAP7_75t_L g150 ( 
.A(n_129),
.Y(n_150)
);

HB1xp67_ASAP7_75t_L g153 ( 
.A(n_150),
.Y(n_153)
);

XOR2xp5_ASAP7_75t_L g161 ( 
.A(n_151),
.B(n_149),
.Y(n_161)
);

NOR2xp33_ASAP7_75t_L g164 ( 
.A(n_152),
.B(n_3),
.Y(n_164)
);

MAJIxp5_ASAP7_75t_L g155 ( 
.A(n_143),
.B(n_139),
.C(n_148),
.Y(n_155)
);

MAJIxp5_ASAP7_75t_L g168 ( 
.A(n_155),
.B(n_159),
.C(n_160),
.Y(n_168)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_156),
.Y(n_167)
);

AOI22xp5_ASAP7_75t_L g157 ( 
.A1(n_144),
.A2(n_22),
.B1(n_18),
.B2(n_27),
.Y(n_157)
);

INVxp67_ASAP7_75t_L g165 ( 
.A(n_157),
.Y(n_165)
);

MAJIxp5_ASAP7_75t_L g159 ( 
.A(n_143),
.B(n_22),
.C(n_17),
.Y(n_159)
);

MAJIxp5_ASAP7_75t_L g160 ( 
.A(n_140),
.B(n_17),
.C(n_3),
.Y(n_160)
);

AND2x2_ASAP7_75t_L g171 ( 
.A(n_161),
.B(n_4),
.Y(n_171)
);

AOI22xp5_ASAP7_75t_L g162 ( 
.A1(n_158),
.A2(n_146),
.B1(n_153),
.B2(n_154),
.Y(n_162)
);

AOI22xp5_ASAP7_75t_L g170 ( 
.A1(n_162),
.A2(n_4),
.B1(n_5),
.B2(n_7),
.Y(n_170)
);

OAI21xp5_ASAP7_75t_L g163 ( 
.A1(n_153),
.A2(n_2),
.B(n_3),
.Y(n_163)
);

MAJIxp5_ASAP7_75t_L g174 ( 
.A(n_163),
.B(n_166),
.C(n_12),
.Y(n_174)
);

NOR2xp33_ASAP7_75t_L g172 ( 
.A(n_164),
.B(n_5),
.Y(n_172)
);

XNOR2xp5_ASAP7_75t_L g166 ( 
.A(n_156),
.B(n_17),
.Y(n_166)
);

AOI22xp5_ASAP7_75t_SL g169 ( 
.A1(n_165),
.A2(n_17),
.B1(n_5),
.B2(n_6),
.Y(n_169)
);

OAI22xp5_ASAP7_75t_SL g179 ( 
.A1(n_169),
.A2(n_172),
.B1(n_7),
.B2(n_8),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_L g176 ( 
.A(n_170),
.B(n_171),
.Y(n_176)
);

AOI31xp33_ASAP7_75t_L g173 ( 
.A1(n_161),
.A2(n_7),
.A3(n_8),
.B(n_9),
.Y(n_173)
);

OAI21xp5_ASAP7_75t_L g175 ( 
.A1(n_173),
.A2(n_167),
.B(n_165),
.Y(n_175)
);

MAJIxp5_ASAP7_75t_L g178 ( 
.A(n_174),
.B(n_168),
.C(n_8),
.Y(n_178)
);

NOR2xp33_ASAP7_75t_L g180 ( 
.A(n_175),
.B(n_177),
.Y(n_180)
);

MAJIxp5_ASAP7_75t_L g177 ( 
.A(n_171),
.B(n_168),
.C(n_172),
.Y(n_177)
);

MAJIxp5_ASAP7_75t_L g182 ( 
.A(n_177),
.B(n_9),
.C(n_10),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_L g181 ( 
.A(n_178),
.B(n_179),
.Y(n_181)
);

OR2x2_ASAP7_75t_L g183 ( 
.A(n_180),
.B(n_182),
.Y(n_183)
);

AOI22xp5_ASAP7_75t_SL g184 ( 
.A1(n_181),
.A2(n_176),
.B1(n_10),
.B2(n_12),
.Y(n_184)
);

INVxp67_ASAP7_75t_L g185 ( 
.A(n_184),
.Y(n_185)
);

OAI21xp5_ASAP7_75t_SL g186 ( 
.A1(n_185),
.A2(n_183),
.B(n_9),
.Y(n_186)
);

XNOR2xp5_ASAP7_75t_L g187 ( 
.A(n_186),
.B(n_10),
.Y(n_187)
);


endmodule