module fake_aes_12576_n_515 (n_44, n_69, n_22, n_57, n_52, n_26, n_50, n_33, n_73, n_49, n_60, n_41, n_35, n_65, n_9, n_10, n_19, n_74, n_7, n_29, n_45, n_62, n_36, n_47, n_37, n_34, n_5, n_23, n_8, n_16, n_13, n_70, n_17, n_63, n_14, n_71, n_56, n_42, n_24, n_6, n_4, n_40, n_38, n_64, n_46, n_31, n_58, n_32, n_0, n_55, n_12, n_75, n_72, n_43, n_76, n_68, n_27, n_53, n_67, n_20, n_2, n_54, n_28, n_48, n_11, n_25, n_30, n_59, n_3, n_18, n_66, n_1, n_15, n_61, n_21, n_51, n_39, n_515);
input n_44;
input n_69;
input n_22;
input n_57;
input n_52;
input n_26;
input n_50;
input n_33;
input n_73;
input n_49;
input n_60;
input n_41;
input n_35;
input n_65;
input n_9;
input n_10;
input n_19;
input n_74;
input n_7;
input n_29;
input n_45;
input n_62;
input n_36;
input n_47;
input n_37;
input n_34;
input n_5;
input n_23;
input n_8;
input n_16;
input n_13;
input n_70;
input n_17;
input n_63;
input n_14;
input n_71;
input n_56;
input n_42;
input n_24;
input n_6;
input n_4;
input n_40;
input n_38;
input n_64;
input n_46;
input n_31;
input n_58;
input n_32;
input n_0;
input n_55;
input n_12;
input n_75;
input n_72;
input n_43;
input n_76;
input n_68;
input n_27;
input n_53;
input n_67;
input n_20;
input n_2;
input n_54;
input n_28;
input n_48;
input n_11;
input n_25;
input n_30;
input n_59;
input n_3;
input n_18;
input n_66;
input n_1;
input n_15;
input n_61;
input n_21;
input n_51;
input n_39;
output n_515;
wire n_117;
wire n_361;
wire n_513;
wire n_185;
wire n_407;
wire n_284;
wire n_278;
wire n_500;
wire n_114;
wire n_94;
wire n_125;
wire n_431;
wire n_484;
wire n_161;
wire n_496;
wire n_177;
wire n_130;
wire n_189;
wire n_311;
wire n_292;
wire n_309;
wire n_160;
wire n_154;
wire n_328;
wire n_468;
wire n_229;
wire n_336;
wire n_464;
wire n_448;
wire n_348;
wire n_252;
wire n_152;
wire n_113;
wire n_353;
wire n_206;
wire n_288;
wire n_383;
wire n_400;
wire n_296;
wire n_157;
wire n_79;
wire n_202;
wire n_386;
wire n_432;
wire n_142;
wire n_232;
wire n_462;
wire n_316;
wire n_211;
wire n_334;
wire n_389;
wire n_436;
wire n_275;
wire n_463;
wire n_131;
wire n_112;
wire n_205;
wire n_330;
wire n_162;
wire n_387;
wire n_163;
wire n_434;
wire n_105;
wire n_227;
wire n_384;
wire n_476;
wire n_231;
wire n_452;
wire n_298;
wire n_411;
wire n_144;
wire n_183;
wire n_489;
wire n_199;
wire n_351;
wire n_83;
wire n_401;
wire n_100;
wire n_305;
wire n_461;
wire n_228;
wire n_345;
wire n_360;
wire n_236;
wire n_340;
wire n_481;
wire n_443;
wire n_150;
wire n_373;
wire n_301;
wire n_222;
wire n_234;
wire n_465;
wire n_366;
wire n_286;
wire n_190;
wire n_246;
wire n_321;
wire n_324;
wire n_392;
wire n_279;
wire n_303;
wire n_437;
wire n_512;
wire n_326;
wire n_289;
wire n_333;
wire n_249;
wire n_244;
wire n_119;
wire n_141;
wire n_479;
wire n_97;
wire n_167;
wire n_447;
wire n_171;
wire n_196;
wire n_192;
wire n_502;
wire n_312;
wire n_455;
wire n_137;
wire n_511;
wire n_277;
wire n_467;
wire n_367;
wire n_250;
wire n_85;
wire n_314;
wire n_237;
wire n_181;
wire n_101;
wire n_255;
wire n_426;
wire n_91;
wire n_108;
wire n_116;
wire n_230;
wire n_209;
wire n_274;
wire n_282;
wire n_319;
wire n_499;
wire n_417;
wire n_241;
wire n_95;
wire n_238;
wire n_318;
wire n_471;
wire n_293;
wire n_506;
wire n_135;
wire n_393;
wire n_247;
wire n_490;
wire n_381;
wire n_304;
wire n_399;
wire n_294;
wire n_459;
wire n_313;
wire n_210;
wire n_184;
wire n_322;
wire n_310;
wire n_191;
wire n_307;
wire n_474;
wire n_354;
wire n_402;
wire n_413;
wire n_391;
wire n_427;
wire n_460;
wire n_478;
wire n_243;
wire n_235;
wire n_415;
wire n_394;
wire n_482;
wire n_442;
wire n_331;
wire n_485;
wire n_352;
wire n_268;
wire n_174;
wire n_501;
wire n_248;
wire n_299;
wire n_89;
wire n_338;
wire n_256;
wire n_77;
wire n_404;
wire n_369;
wire n_509;
wire n_172;
wire n_329;
wire n_251;
wire n_218;
wire n_507;
wire n_271;
wire n_302;
wire n_466;
wire n_270;
wire n_362;
wire n_153;
wire n_259;
wire n_308;
wire n_93;
wire n_412;
wire n_140;
wire n_207;
wire n_224;
wire n_96;
wire n_219;
wire n_475;
wire n_133;
wire n_149;
wire n_81;
wire n_214;
wire n_204;
wire n_430;
wire n_88;
wire n_450;
wire n_107;
wire n_403;
wire n_254;
wire n_262;
wire n_239;
wire n_439;
wire n_87;
wire n_379;
wire n_98;
wire n_276;
wire n_320;
wire n_285;
wire n_195;
wire n_165;
wire n_420;
wire n_423;
wire n_342;
wire n_446;
wire n_370;
wire n_217;
wire n_139;
wire n_388;
wire n_454;
wire n_193;
wire n_273;
wire n_505;
wire n_390;
wire n_120;
wire n_514;
wire n_486;
wire n_245;
wire n_357;
wire n_90;
wire n_260;
wire n_78;
wire n_197;
wire n_201;
wire n_317;
wire n_416;
wire n_374;
wire n_111;
wire n_265;
wire n_264;
wire n_200;
wire n_208;
wire n_126;
wire n_178;
wire n_118;
wire n_365;
wire n_179;
wire n_315;
wire n_363;
wire n_409;
wire n_86;
wire n_143;
wire n_295;
wire n_263;
wire n_166;
wire n_495;
wire n_186;
wire n_364;
wire n_428;
wire n_376;
wire n_344;
wire n_136;
wire n_503;
wire n_283;
wire n_435;
wire n_216;
wire n_147;
wire n_148;
wire n_212;
wire n_472;
wire n_92;
wire n_419;
wire n_396;
wire n_168;
wire n_477;
wire n_508;
wire n_398;
wire n_445;
wire n_438;
wire n_134;
wire n_429;
wire n_488;
wire n_233;
wire n_82;
wire n_106;
wire n_440;
wire n_173;
wire n_422;
wire n_327;
wire n_325;
wire n_349;
wire n_498;
wire n_225;
wire n_220;
wire n_358;
wire n_267;
wire n_221;
wire n_456;
wire n_203;
wire n_102;
wire n_449;
wire n_115;
wire n_80;
wire n_300;
wire n_158;
wire n_121;
wire n_497;
wire n_339;
wire n_240;
wire n_378;
wire n_359;
wire n_346;
wire n_103;
wire n_180;
wire n_441;
wire n_104;
wire n_335;
wire n_272;
wire n_146;
wire n_397;
wire n_306;
wire n_215;
wire n_242;
wire n_155;
wire n_198;
wire n_169;
wire n_424;
wire n_156;
wire n_124;
wire n_297;
wire n_128;
wire n_129;
wire n_410;
wire n_188;
wire n_377;
wire n_510;
wire n_343;
wire n_127;
wire n_291;
wire n_170;
wire n_504;
wire n_458;
wire n_418;
wire n_493;
wire n_380;
wire n_356;
wire n_281;
wire n_341;
wire n_470;
wire n_122;
wire n_187;
wire n_375;
wire n_138;
wire n_451;
wire n_487;
wire n_371;
wire n_323;
wire n_473;
wire n_347;
wire n_258;
wire n_253;
wire n_84;
wire n_266;
wire n_213;
wire n_182;
wire n_492;
wire n_368;
wire n_355;
wire n_226;
wire n_382;
wire n_159;
wire n_337;
wire n_444;
wire n_176;
wire n_469;
wire n_123;
wire n_457;
wire n_223;
wire n_494;
wire n_480;
wire n_372;
wire n_453;
wire n_194;
wire n_287;
wire n_110;
wire n_261;
wire n_425;
wire n_332;
wire n_414;
wire n_350;
wire n_433;
wire n_164;
wire n_421;
wire n_175;
wire n_145;
wire n_483;
wire n_408;
wire n_290;
wire n_405;
wire n_280;
wire n_132;
wire n_99;
wire n_109;
wire n_406;
wire n_395;
wire n_491;
wire n_151;
wire n_385;
wire n_257;
wire n_269;
CKINVDCx20_ASAP7_75t_R g77 ( .A(n_33), .Y(n_77) );
INVx1_ASAP7_75t_L g78 ( .A(n_52), .Y(n_78) );
INVxp67_ASAP7_75t_SL g79 ( .A(n_16), .Y(n_79) );
INVx1_ASAP7_75t_L g80 ( .A(n_43), .Y(n_80) );
INVx1_ASAP7_75t_L g81 ( .A(n_5), .Y(n_81) );
INVx1_ASAP7_75t_L g82 ( .A(n_40), .Y(n_82) );
INVx1_ASAP7_75t_L g83 ( .A(n_13), .Y(n_83) );
INVxp33_ASAP7_75t_L g84 ( .A(n_49), .Y(n_84) );
INVx1_ASAP7_75t_L g85 ( .A(n_50), .Y(n_85) );
BUFx3_ASAP7_75t_L g86 ( .A(n_42), .Y(n_86) );
INVx1_ASAP7_75t_L g87 ( .A(n_35), .Y(n_87) );
INVx1_ASAP7_75t_L g88 ( .A(n_71), .Y(n_88) );
INVxp67_ASAP7_75t_L g89 ( .A(n_57), .Y(n_89) );
CKINVDCx5p33_ASAP7_75t_R g90 ( .A(n_4), .Y(n_90) );
INVx1_ASAP7_75t_L g91 ( .A(n_39), .Y(n_91) );
INVxp67_ASAP7_75t_L g92 ( .A(n_63), .Y(n_92) );
CKINVDCx5p33_ASAP7_75t_R g93 ( .A(n_68), .Y(n_93) );
BUFx3_ASAP7_75t_L g94 ( .A(n_60), .Y(n_94) );
INVx1_ASAP7_75t_L g95 ( .A(n_31), .Y(n_95) );
INVx1_ASAP7_75t_L g96 ( .A(n_53), .Y(n_96) );
INVx1_ASAP7_75t_L g97 ( .A(n_8), .Y(n_97) );
INVx2_ASAP7_75t_L g98 ( .A(n_73), .Y(n_98) );
INVx1_ASAP7_75t_L g99 ( .A(n_28), .Y(n_99) );
INVxp67_ASAP7_75t_L g100 ( .A(n_37), .Y(n_100) );
INVx1_ASAP7_75t_SL g101 ( .A(n_4), .Y(n_101) );
INVx1_ASAP7_75t_L g102 ( .A(n_69), .Y(n_102) );
INVx1_ASAP7_75t_L g103 ( .A(n_19), .Y(n_103) );
BUFx3_ASAP7_75t_L g104 ( .A(n_19), .Y(n_104) );
INVx2_ASAP7_75t_L g105 ( .A(n_58), .Y(n_105) );
INVx1_ASAP7_75t_L g106 ( .A(n_27), .Y(n_106) );
INVx1_ASAP7_75t_L g107 ( .A(n_10), .Y(n_107) );
INVx1_ASAP7_75t_L g108 ( .A(n_20), .Y(n_108) );
INVx1_ASAP7_75t_L g109 ( .A(n_18), .Y(n_109) );
INVx1_ASAP7_75t_L g110 ( .A(n_65), .Y(n_110) );
CKINVDCx16_ASAP7_75t_R g111 ( .A(n_66), .Y(n_111) );
CKINVDCx5p33_ASAP7_75t_R g112 ( .A(n_17), .Y(n_112) );
CKINVDCx16_ASAP7_75t_R g113 ( .A(n_64), .Y(n_113) );
INVx1_ASAP7_75t_L g114 ( .A(n_9), .Y(n_114) );
AND2x2_ASAP7_75t_L g115 ( .A(n_84), .B(n_0), .Y(n_115) );
INVx1_ASAP7_75t_L g116 ( .A(n_78), .Y(n_116) );
INVx3_ASAP7_75t_L g117 ( .A(n_104), .Y(n_117) );
BUFx6f_ASAP7_75t_L g118 ( .A(n_86), .Y(n_118) );
AND2x4_ASAP7_75t_L g119 ( .A(n_104), .B(n_0), .Y(n_119) );
BUFx6f_ASAP7_75t_L g120 ( .A(n_86), .Y(n_120) );
INVx2_ASAP7_75t_L g121 ( .A(n_98), .Y(n_121) );
BUFx6f_ASAP7_75t_L g122 ( .A(n_94), .Y(n_122) );
INVx1_ASAP7_75t_L g123 ( .A(n_78), .Y(n_123) );
INVx1_ASAP7_75t_L g124 ( .A(n_80), .Y(n_124) );
NAND2xp5_ASAP7_75t_L g125 ( .A(n_81), .B(n_1), .Y(n_125) );
AND2x4_ASAP7_75t_L g126 ( .A(n_81), .B(n_1), .Y(n_126) );
AND2x2_ASAP7_75t_L g127 ( .A(n_111), .B(n_2), .Y(n_127) );
NAND2xp5_ASAP7_75t_L g128 ( .A(n_83), .B(n_2), .Y(n_128) );
INVxp67_ASAP7_75t_L g129 ( .A(n_83), .Y(n_129) );
AND2x4_ASAP7_75t_L g130 ( .A(n_97), .B(n_3), .Y(n_130) );
INVx2_ASAP7_75t_L g131 ( .A(n_98), .Y(n_131) );
AND2x2_ASAP7_75t_L g132 ( .A(n_113), .B(n_3), .Y(n_132) );
BUFx6f_ASAP7_75t_L g133 ( .A(n_94), .Y(n_133) );
NAND2xp5_ASAP7_75t_L g134 ( .A(n_97), .B(n_5), .Y(n_134) );
INVx2_ASAP7_75t_L g135 ( .A(n_105), .Y(n_135) );
INVx1_ASAP7_75t_L g136 ( .A(n_80), .Y(n_136) );
NOR2xp33_ASAP7_75t_L g137 ( .A(n_129), .B(n_89), .Y(n_137) );
AND2x4_ASAP7_75t_L g138 ( .A(n_119), .B(n_103), .Y(n_138) );
INVx3_ASAP7_75t_L g139 ( .A(n_126), .Y(n_139) );
NOR2xp33_ASAP7_75t_L g140 ( .A(n_129), .B(n_92), .Y(n_140) );
AND2x4_ASAP7_75t_L g141 ( .A(n_119), .B(n_103), .Y(n_141) );
AOI22xp5_ASAP7_75t_L g142 ( .A1(n_126), .A2(n_77), .B1(n_112), .B2(n_90), .Y(n_142) );
NAND2xp5_ASAP7_75t_L g143 ( .A(n_115), .B(n_93), .Y(n_143) );
NAND2x1p5_ASAP7_75t_L g144 ( .A(n_126), .B(n_82), .Y(n_144) );
INVx2_ASAP7_75t_SL g145 ( .A(n_115), .Y(n_145) );
BUFx2_ASAP7_75t_L g146 ( .A(n_127), .Y(n_146) );
CKINVDCx5p33_ASAP7_75t_R g147 ( .A(n_127), .Y(n_147) );
INVx1_ASAP7_75t_L g148 ( .A(n_121), .Y(n_148) );
INVx1_ASAP7_75t_SL g149 ( .A(n_127), .Y(n_149) );
INVx1_ASAP7_75t_L g150 ( .A(n_121), .Y(n_150) );
INVx1_ASAP7_75t_L g151 ( .A(n_121), .Y(n_151) );
AO22x2_ASAP7_75t_L g152 ( .A1(n_119), .A2(n_102), .B1(n_110), .B2(n_91), .Y(n_152) );
INVx4_ASAP7_75t_L g153 ( .A(n_119), .Y(n_153) );
AND2x4_ASAP7_75t_L g154 ( .A(n_126), .B(n_107), .Y(n_154) );
NAND2x1p5_ASAP7_75t_L g155 ( .A(n_130), .B(n_82), .Y(n_155) );
NAND2xp5_ASAP7_75t_L g156 ( .A(n_115), .B(n_100), .Y(n_156) );
NAND2xp5_ASAP7_75t_SL g157 ( .A(n_116), .B(n_102), .Y(n_157) );
INVx2_ASAP7_75t_L g158 ( .A(n_118), .Y(n_158) );
INVx1_ASAP7_75t_L g159 ( .A(n_131), .Y(n_159) );
BUFx3_ASAP7_75t_L g160 ( .A(n_117), .Y(n_160) );
AND2x4_ASAP7_75t_L g161 ( .A(n_130), .B(n_114), .Y(n_161) );
BUFx6f_ASAP7_75t_L g162 ( .A(n_160), .Y(n_162) );
INVx3_ASAP7_75t_L g163 ( .A(n_153), .Y(n_163) );
BUFx6f_ASAP7_75t_L g164 ( .A(n_160), .Y(n_164) );
AOI21xp5_ASAP7_75t_L g165 ( .A1(n_139), .A2(n_136), .B(n_124), .Y(n_165) );
NAND2xp33_ASAP7_75t_L g166 ( .A(n_144), .B(n_132), .Y(n_166) );
AOI22xp33_ASAP7_75t_L g167 ( .A1(n_152), .A2(n_130), .B1(n_132), .B2(n_123), .Y(n_167) );
INVx2_ASAP7_75t_L g168 ( .A(n_158), .Y(n_168) );
NOR2xp33_ASAP7_75t_L g169 ( .A(n_156), .B(n_116), .Y(n_169) );
INVx1_ASAP7_75t_L g170 ( .A(n_139), .Y(n_170) );
BUFx4f_ASAP7_75t_L g171 ( .A(n_144), .Y(n_171) );
AND2x4_ASAP7_75t_L g172 ( .A(n_145), .B(n_132), .Y(n_172) );
BUFx12f_ASAP7_75t_L g173 ( .A(n_146), .Y(n_173) );
CKINVDCx8_ASAP7_75t_R g174 ( .A(n_146), .Y(n_174) );
NAND2xp5_ASAP7_75t_SL g175 ( .A(n_145), .B(n_130), .Y(n_175) );
INVx5_ASAP7_75t_L g176 ( .A(n_153), .Y(n_176) );
INVx2_ASAP7_75t_SL g177 ( .A(n_144), .Y(n_177) );
OR2x2_ASAP7_75t_L g178 ( .A(n_149), .B(n_125), .Y(n_178) );
NAND2xp5_ASAP7_75t_L g179 ( .A(n_137), .B(n_123), .Y(n_179) );
BUFx3_ASAP7_75t_L g180 ( .A(n_155), .Y(n_180) );
INVx1_ASAP7_75t_L g181 ( .A(n_139), .Y(n_181) );
INVx1_ASAP7_75t_L g182 ( .A(n_139), .Y(n_182) );
INVx5_ASAP7_75t_L g183 ( .A(n_153), .Y(n_183) );
NAND2xp5_ASAP7_75t_L g184 ( .A(n_140), .B(n_124), .Y(n_184) );
INVx4_ASAP7_75t_L g185 ( .A(n_153), .Y(n_185) );
NAND2x1p5_ASAP7_75t_L g186 ( .A(n_138), .B(n_136), .Y(n_186) );
NAND2x1p5_ASAP7_75t_L g187 ( .A(n_138), .B(n_85), .Y(n_187) );
INVx2_ASAP7_75t_SL g188 ( .A(n_155), .Y(n_188) );
INVx1_ASAP7_75t_L g189 ( .A(n_148), .Y(n_189) );
INVx2_ASAP7_75t_L g190 ( .A(n_158), .Y(n_190) );
INVx1_ASAP7_75t_L g191 ( .A(n_148), .Y(n_191) );
BUFx6f_ASAP7_75t_L g192 ( .A(n_155), .Y(n_192) );
INVx2_ASAP7_75t_L g193 ( .A(n_150), .Y(n_193) );
INVx3_ASAP7_75t_L g194 ( .A(n_192), .Y(n_194) );
CKINVDCx16_ASAP7_75t_R g195 ( .A(n_173), .Y(n_195) );
INVx4_ASAP7_75t_L g196 ( .A(n_171), .Y(n_196) );
AND2x2_ASAP7_75t_L g197 ( .A(n_178), .B(n_147), .Y(n_197) );
HB1xp67_ASAP7_75t_L g198 ( .A(n_174), .Y(n_198) );
NAND2xp5_ASAP7_75t_L g199 ( .A(n_169), .B(n_152), .Y(n_199) );
AOI22xp5_ASAP7_75t_L g200 ( .A1(n_166), .A2(n_152), .B1(n_141), .B2(n_138), .Y(n_200) );
AOI22xp33_ASAP7_75t_L g201 ( .A1(n_167), .A2(n_152), .B1(n_138), .B2(n_141), .Y(n_201) );
BUFx2_ASAP7_75t_L g202 ( .A(n_180), .Y(n_202) );
INVx1_ASAP7_75t_L g203 ( .A(n_193), .Y(n_203) );
NAND2xp5_ASAP7_75t_L g204 ( .A(n_178), .B(n_154), .Y(n_204) );
INVx2_ASAP7_75t_L g205 ( .A(n_193), .Y(n_205) );
INVx1_ASAP7_75t_SL g206 ( .A(n_192), .Y(n_206) );
BUFx3_ASAP7_75t_L g207 ( .A(n_180), .Y(n_207) );
OAI22xp5_ASAP7_75t_SL g208 ( .A1(n_174), .A2(n_142), .B1(n_79), .B2(n_101), .Y(n_208) );
BUFx8_ASAP7_75t_SL g209 ( .A(n_173), .Y(n_209) );
NAND2xp5_ASAP7_75t_L g210 ( .A(n_186), .B(n_154), .Y(n_210) );
O2A1O1Ixp33_ASAP7_75t_L g211 ( .A1(n_179), .A2(n_157), .B(n_128), .C(n_134), .Y(n_211) );
AOI21xp5_ASAP7_75t_L g212 ( .A1(n_175), .A2(n_161), .B(n_154), .Y(n_212) );
INVx1_ASAP7_75t_L g213 ( .A(n_193), .Y(n_213) );
OR2x2_ASAP7_75t_L g214 ( .A(n_172), .B(n_142), .Y(n_214) );
INVx2_ASAP7_75t_SL g215 ( .A(n_171), .Y(n_215) );
INVx2_ASAP7_75t_L g216 ( .A(n_189), .Y(n_216) );
BUFx6f_ASAP7_75t_L g217 ( .A(n_192), .Y(n_217) );
BUFx12f_ASAP7_75t_L g218 ( .A(n_192), .Y(n_218) );
INVx2_ASAP7_75t_SL g219 ( .A(n_171), .Y(n_219) );
INVx1_ASAP7_75t_L g220 ( .A(n_189), .Y(n_220) );
INVx1_ASAP7_75t_L g221 ( .A(n_191), .Y(n_221) );
A2O1A1Ixp33_ASAP7_75t_L g222 ( .A1(n_165), .A2(n_141), .B(n_161), .C(n_154), .Y(n_222) );
INVx2_ASAP7_75t_L g223 ( .A(n_191), .Y(n_223) );
BUFx8_ASAP7_75t_L g224 ( .A(n_180), .Y(n_224) );
INVx1_ASAP7_75t_L g225 ( .A(n_170), .Y(n_225) );
AND2x2_ASAP7_75t_L g226 ( .A(n_197), .B(n_172), .Y(n_226) );
AOI221x1_ASAP7_75t_L g227 ( .A1(n_199), .A2(n_118), .B1(n_120), .B2(n_122), .C(n_133), .Y(n_227) );
BUFx6f_ASAP7_75t_L g228 ( .A(n_218), .Y(n_228) );
OAI21xp5_ASAP7_75t_L g229 ( .A1(n_222), .A2(n_182), .B(n_170), .Y(n_229) );
CKINVDCx5p33_ASAP7_75t_R g230 ( .A(n_209), .Y(n_230) );
INVx1_ASAP7_75t_L g231 ( .A(n_203), .Y(n_231) );
AOI22xp5_ASAP7_75t_L g232 ( .A1(n_200), .A2(n_171), .B1(n_172), .B2(n_188), .Y(n_232) );
INVx1_ASAP7_75t_L g233 ( .A(n_203), .Y(n_233) );
OAI22xp5_ASAP7_75t_L g234 ( .A1(n_200), .A2(n_187), .B1(n_188), .B2(n_177), .Y(n_234) );
INVx3_ASAP7_75t_L g235 ( .A(n_218), .Y(n_235) );
AOI22xp33_ASAP7_75t_L g236 ( .A1(n_208), .A2(n_172), .B1(n_177), .B2(n_187), .Y(n_236) );
BUFx6f_ASAP7_75t_L g237 ( .A(n_218), .Y(n_237) );
AOI22xp33_ASAP7_75t_SL g238 ( .A1(n_208), .A2(n_192), .B1(n_187), .B2(n_186), .Y(n_238) );
OAI22xp33_ASAP7_75t_SL g239 ( .A1(n_214), .A2(n_186), .B1(n_134), .B2(n_128), .Y(n_239) );
AOI22xp33_ASAP7_75t_L g240 ( .A1(n_197), .A2(n_192), .B1(n_185), .B2(n_141), .Y(n_240) );
INVx2_ASAP7_75t_L g241 ( .A(n_205), .Y(n_241) );
OAI22xp33_ASAP7_75t_L g242 ( .A1(n_195), .A2(n_143), .B1(n_184), .B2(n_185), .Y(n_242) );
BUFx12f_ASAP7_75t_L g243 ( .A(n_224), .Y(n_243) );
OAI22xp5_ASAP7_75t_L g244 ( .A1(n_201), .A2(n_161), .B1(n_185), .B2(n_182), .Y(n_244) );
CKINVDCx5p33_ASAP7_75t_R g245 ( .A(n_195), .Y(n_245) );
INVx2_ASAP7_75t_L g246 ( .A(n_205), .Y(n_246) );
CKINVDCx20_ASAP7_75t_R g247 ( .A(n_224), .Y(n_247) );
OAI22xp33_ASAP7_75t_L g248 ( .A1(n_214), .A2(n_185), .B1(n_183), .B2(n_176), .Y(n_248) );
AOI22xp33_ASAP7_75t_L g249 ( .A1(n_199), .A2(n_163), .B1(n_161), .B2(n_181), .Y(n_249) );
INVx1_ASAP7_75t_L g250 ( .A(n_213), .Y(n_250) );
OAI22xp5_ASAP7_75t_L g251 ( .A1(n_204), .A2(n_181), .B1(n_183), .B2(n_176), .Y(n_251) );
AOI22xp33_ASAP7_75t_SL g252 ( .A1(n_224), .A2(n_125), .B1(n_163), .B2(n_176), .Y(n_252) );
AOI22xp33_ASAP7_75t_L g253 ( .A1(n_238), .A2(n_198), .B1(n_224), .B2(n_204), .Y(n_253) );
AND2x4_ASAP7_75t_L g254 ( .A(n_228), .B(n_196), .Y(n_254) );
AND2x2_ASAP7_75t_L g255 ( .A(n_231), .B(n_213), .Y(n_255) );
OAI31xp33_ASAP7_75t_L g256 ( .A1(n_242), .A2(n_210), .A3(n_108), .B(n_109), .Y(n_256) );
AOI22xp33_ASAP7_75t_L g257 ( .A1(n_236), .A2(n_196), .B1(n_221), .B2(n_220), .Y(n_257) );
OAI21xp33_ASAP7_75t_L g258 ( .A1(n_239), .A2(n_205), .B(n_223), .Y(n_258) );
INVx2_ASAP7_75t_L g259 ( .A(n_241), .Y(n_259) );
BUFx2_ASAP7_75t_L g260 ( .A(n_228), .Y(n_260) );
NAND2xp5_ASAP7_75t_L g261 ( .A(n_231), .B(n_233), .Y(n_261) );
AOI22xp33_ASAP7_75t_L g262 ( .A1(n_226), .A2(n_196), .B1(n_221), .B2(n_220), .Y(n_262) );
AO21x2_ASAP7_75t_L g263 ( .A1(n_229), .A2(n_223), .B(n_216), .Y(n_263) );
AOI22xp33_ASAP7_75t_L g264 ( .A1(n_226), .A2(n_196), .B1(n_202), .B2(n_223), .Y(n_264) );
NAND2xp5_ASAP7_75t_L g265 ( .A(n_233), .B(n_216), .Y(n_265) );
AOI221xp5_ASAP7_75t_L g266 ( .A1(n_240), .A2(n_211), .B1(n_212), .B2(n_216), .C(n_108), .Y(n_266) );
NAND3xp33_ASAP7_75t_L g267 ( .A(n_227), .B(n_217), .C(n_118), .Y(n_267) );
AOI221xp5_ASAP7_75t_L g268 ( .A1(n_248), .A2(n_107), .B1(n_109), .B2(n_114), .C(n_135), .Y(n_268) );
AOI22xp33_ASAP7_75t_L g269 ( .A1(n_243), .A2(n_202), .B1(n_207), .B2(n_210), .Y(n_269) );
INVx2_ASAP7_75t_L g270 ( .A(n_241), .Y(n_270) );
OAI22xp5_ASAP7_75t_L g271 ( .A1(n_232), .A2(n_207), .B1(n_206), .B2(n_217), .Y(n_271) );
OAI211xp5_ASAP7_75t_L g272 ( .A1(n_232), .A2(n_135), .B(n_131), .C(n_117), .Y(n_272) );
INVx2_ASAP7_75t_L g273 ( .A(n_246), .Y(n_273) );
AOI22xp33_ASAP7_75t_L g274 ( .A1(n_243), .A2(n_207), .B1(n_225), .B2(n_215), .Y(n_274) );
OAI221xp5_ASAP7_75t_L g275 ( .A1(n_256), .A2(n_252), .B1(n_249), .B2(n_234), .C(n_244), .Y(n_275) );
OA21x2_ASAP7_75t_L g276 ( .A1(n_267), .A2(n_227), .B(n_250), .Y(n_276) );
AOI221xp5_ASAP7_75t_L g277 ( .A1(n_256), .A2(n_250), .B1(n_247), .B2(n_245), .C(n_117), .Y(n_277) );
AND2x2_ASAP7_75t_SL g278 ( .A(n_253), .B(n_228), .Y(n_278) );
AND2x2_ASAP7_75t_L g279 ( .A(n_255), .B(n_246), .Y(n_279) );
OAI221xp5_ASAP7_75t_L g280 ( .A1(n_268), .A2(n_235), .B1(n_251), .B2(n_237), .C(n_228), .Y(n_280) );
OAI221xp5_ASAP7_75t_SL g281 ( .A1(n_268), .A2(n_235), .B1(n_87), .B2(n_85), .C(n_88), .Y(n_281) );
BUFx2_ASAP7_75t_L g282 ( .A(n_260), .Y(n_282) );
INVx1_ASAP7_75t_L g283 ( .A(n_261), .Y(n_283) );
AOI221xp5_ASAP7_75t_L g284 ( .A1(n_266), .A2(n_245), .B1(n_131), .B2(n_135), .C(n_117), .Y(n_284) );
AOI22xp33_ASAP7_75t_L g285 ( .A1(n_257), .A2(n_237), .B1(n_228), .B2(n_235), .Y(n_285) );
INVx2_ASAP7_75t_L g286 ( .A(n_259), .Y(n_286) );
OAI211xp5_ASAP7_75t_L g287 ( .A1(n_269), .A2(n_230), .B(n_87), .C(n_88), .Y(n_287) );
NOR2x1_ASAP7_75t_R g288 ( .A(n_260), .B(n_230), .Y(n_288) );
OAI21xp33_ASAP7_75t_L g289 ( .A1(n_258), .A2(n_237), .B(n_91), .Y(n_289) );
AOI211xp5_ASAP7_75t_SL g290 ( .A1(n_271), .A2(n_194), .B(n_96), .C(n_99), .Y(n_290) );
INVx2_ASAP7_75t_L g291 ( .A(n_259), .Y(n_291) );
AND2x2_ASAP7_75t_L g292 ( .A(n_255), .B(n_237), .Y(n_292) );
NOR2xp33_ASAP7_75t_R g293 ( .A(n_254), .B(n_237), .Y(n_293) );
AOI221xp5_ASAP7_75t_L g294 ( .A1(n_258), .A2(n_159), .B1(n_150), .B2(n_151), .C(n_225), .Y(n_294) );
INVx2_ASAP7_75t_L g295 ( .A(n_259), .Y(n_295) );
NOR2xp33_ASAP7_75t_L g296 ( .A(n_254), .B(n_215), .Y(n_296) );
AND2x2_ASAP7_75t_L g297 ( .A(n_279), .B(n_270), .Y(n_297) );
OAI31xp33_ASAP7_75t_SL g298 ( .A1(n_277), .A2(n_271), .A3(n_267), .B(n_254), .Y(n_298) );
INVx2_ASAP7_75t_L g299 ( .A(n_286), .Y(n_299) );
NAND4xp25_ASAP7_75t_L g300 ( .A(n_277), .B(n_262), .C(n_96), .D(n_99), .Y(n_300) );
BUFx2_ASAP7_75t_L g301 ( .A(n_282), .Y(n_301) );
NAND3xp33_ASAP7_75t_L g302 ( .A(n_290), .B(n_272), .C(n_95), .Y(n_302) );
INVx4_ASAP7_75t_L g303 ( .A(n_278), .Y(n_303) );
OAI31xp33_ASAP7_75t_L g304 ( .A1(n_281), .A2(n_261), .A3(n_254), .B(n_264), .Y(n_304) );
AND2x2_ASAP7_75t_L g305 ( .A(n_279), .B(n_270), .Y(n_305) );
AO22x1_ASAP7_75t_L g306 ( .A1(n_282), .A2(n_265), .B1(n_273), .B2(n_270), .Y(n_306) );
INVx2_ASAP7_75t_L g307 ( .A(n_286), .Y(n_307) );
HB1xp67_ASAP7_75t_L g308 ( .A(n_286), .Y(n_308) );
OR2x2_ASAP7_75t_L g309 ( .A(n_283), .B(n_265), .Y(n_309) );
INVx2_ASAP7_75t_SL g310 ( .A(n_291), .Y(n_310) );
INVx2_ASAP7_75t_L g311 ( .A(n_291), .Y(n_311) );
INVx1_ASAP7_75t_L g312 ( .A(n_291), .Y(n_312) );
AND2x4_ASAP7_75t_L g313 ( .A(n_295), .B(n_263), .Y(n_313) );
AND2x2_ASAP7_75t_L g314 ( .A(n_292), .B(n_273), .Y(n_314) );
AND2x2_ASAP7_75t_L g315 ( .A(n_292), .B(n_273), .Y(n_315) );
OAI31xp33_ASAP7_75t_L g316 ( .A1(n_280), .A2(n_219), .A3(n_274), .B(n_95), .Y(n_316) );
AND2x2_ASAP7_75t_L g317 ( .A(n_295), .B(n_263), .Y(n_317) );
INVx2_ASAP7_75t_L g318 ( .A(n_295), .Y(n_318) );
INVx2_ASAP7_75t_SL g319 ( .A(n_293), .Y(n_319) );
OAI221xp5_ASAP7_75t_L g320 ( .A1(n_280), .A2(n_110), .B1(n_106), .B2(n_219), .C(n_105), .Y(n_320) );
HB1xp67_ASAP7_75t_L g321 ( .A(n_283), .Y(n_321) );
OAI221xp5_ASAP7_75t_L g322 ( .A1(n_275), .A2(n_106), .B1(n_206), .B2(n_159), .C(n_151), .Y(n_322) );
OAI31xp33_ASAP7_75t_L g323 ( .A1(n_275), .A2(n_194), .A3(n_163), .B(n_8), .Y(n_323) );
INVx1_ASAP7_75t_L g324 ( .A(n_276), .Y(n_324) );
OAI221xp5_ASAP7_75t_L g325 ( .A1(n_290), .A2(n_194), .B1(n_217), .B2(n_118), .C(n_120), .Y(n_325) );
AND2x4_ASAP7_75t_SL g326 ( .A(n_303), .B(n_319), .Y(n_326) );
NAND2xp5_ASAP7_75t_SL g327 ( .A(n_319), .B(n_278), .Y(n_327) );
AND2x2_ASAP7_75t_L g328 ( .A(n_310), .B(n_276), .Y(n_328) );
INVx1_ASAP7_75t_L g329 ( .A(n_312), .Y(n_329) );
INVx2_ASAP7_75t_L g330 ( .A(n_299), .Y(n_330) );
INVx1_ASAP7_75t_L g331 ( .A(n_321), .Y(n_331) );
NAND2xp5_ASAP7_75t_L g332 ( .A(n_297), .B(n_288), .Y(n_332) );
NAND2xp5_ASAP7_75t_L g333 ( .A(n_297), .B(n_288), .Y(n_333) );
INVx2_ASAP7_75t_L g334 ( .A(n_299), .Y(n_334) );
INVx2_ASAP7_75t_L g335 ( .A(n_299), .Y(n_335) );
OR2x2_ASAP7_75t_L g336 ( .A(n_301), .B(n_263), .Y(n_336) );
INVx1_ASAP7_75t_L g337 ( .A(n_321), .Y(n_337) );
AND2x2_ASAP7_75t_L g338 ( .A(n_310), .B(n_276), .Y(n_338) );
INVx1_ASAP7_75t_L g339 ( .A(n_308), .Y(n_339) );
AND2x2_ASAP7_75t_L g340 ( .A(n_310), .B(n_276), .Y(n_340) );
NAND4xp25_ASAP7_75t_L g341 ( .A(n_323), .B(n_287), .C(n_284), .D(n_289), .Y(n_341) );
HB1xp67_ASAP7_75t_L g342 ( .A(n_308), .Y(n_342) );
INVx2_ASAP7_75t_L g343 ( .A(n_307), .Y(n_343) );
AOI21xp5_ASAP7_75t_L g344 ( .A1(n_306), .A2(n_289), .B(n_263), .Y(n_344) );
INVx1_ASAP7_75t_L g345 ( .A(n_307), .Y(n_345) );
OR2x6_ASAP7_75t_L g346 ( .A(n_306), .B(n_296), .Y(n_346) );
NAND2xp5_ASAP7_75t_L g347 ( .A(n_305), .B(n_285), .Y(n_347) );
INVxp67_ASAP7_75t_L g348 ( .A(n_314), .Y(n_348) );
INVx1_ASAP7_75t_L g349 ( .A(n_307), .Y(n_349) );
AND2x2_ASAP7_75t_L g350 ( .A(n_314), .B(n_133), .Y(n_350) );
AND2x2_ASAP7_75t_L g351 ( .A(n_315), .B(n_133), .Y(n_351) );
AND2x2_ASAP7_75t_L g352 ( .A(n_315), .B(n_133), .Y(n_352) );
AND2x2_ASAP7_75t_L g353 ( .A(n_317), .B(n_133), .Y(n_353) );
AND2x2_ASAP7_75t_L g354 ( .A(n_317), .B(n_133), .Y(n_354) );
INVx1_ASAP7_75t_L g355 ( .A(n_311), .Y(n_355) );
AND2x2_ASAP7_75t_L g356 ( .A(n_305), .B(n_133), .Y(n_356) );
INVx1_ASAP7_75t_L g357 ( .A(n_311), .Y(n_357) );
AND2x2_ASAP7_75t_L g358 ( .A(n_311), .B(n_318), .Y(n_358) );
NOR3xp33_ASAP7_75t_L g359 ( .A(n_322), .B(n_294), .C(n_194), .Y(n_359) );
AND2x2_ASAP7_75t_L g360 ( .A(n_318), .B(n_118), .Y(n_360) );
AND2x2_ASAP7_75t_L g361 ( .A(n_318), .B(n_118), .Y(n_361) );
INVx1_ASAP7_75t_L g362 ( .A(n_313), .Y(n_362) );
INVx1_ASAP7_75t_SL g363 ( .A(n_309), .Y(n_363) );
INVx1_ASAP7_75t_L g364 ( .A(n_313), .Y(n_364) );
OAI22xp5_ASAP7_75t_L g365 ( .A1(n_322), .A2(n_217), .B1(n_183), .B2(n_176), .Y(n_365) );
INVxp67_ASAP7_75t_L g366 ( .A(n_309), .Y(n_366) );
OR2x2_ASAP7_75t_L g367 ( .A(n_363), .B(n_348), .Y(n_367) );
NOR2x1_ASAP7_75t_L g368 ( .A(n_346), .B(n_325), .Y(n_368) );
OR2x2_ASAP7_75t_L g369 ( .A(n_363), .B(n_303), .Y(n_369) );
NAND2xp5_ASAP7_75t_L g370 ( .A(n_366), .B(n_324), .Y(n_370) );
NAND2xp5_ASAP7_75t_L g371 ( .A(n_331), .B(n_324), .Y(n_371) );
NAND2xp5_ASAP7_75t_L g372 ( .A(n_331), .B(n_313), .Y(n_372) );
OR2x2_ASAP7_75t_L g373 ( .A(n_342), .B(n_303), .Y(n_373) );
AO211x2_ASAP7_75t_L g374 ( .A1(n_341), .A2(n_333), .B(n_332), .C(n_302), .Y(n_374) );
AND2x2_ASAP7_75t_L g375 ( .A(n_353), .B(n_313), .Y(n_375) );
INVx2_ASAP7_75t_L g376 ( .A(n_358), .Y(n_376) );
OR2x2_ASAP7_75t_L g377 ( .A(n_337), .B(n_320), .Y(n_377) );
AND5x1_ASAP7_75t_L g378 ( .A(n_344), .B(n_298), .C(n_323), .D(n_304), .E(n_316), .Y(n_378) );
OR2x2_ASAP7_75t_L g379 ( .A(n_337), .B(n_320), .Y(n_379) );
NAND2xp5_ASAP7_75t_SL g380 ( .A(n_326), .B(n_298), .Y(n_380) );
INVxp67_ASAP7_75t_L g381 ( .A(n_353), .Y(n_381) );
INVx11_ASAP7_75t_L g382 ( .A(n_326), .Y(n_382) );
OAI322xp33_ASAP7_75t_L g383 ( .A1(n_336), .A2(n_325), .A3(n_302), .B1(n_122), .B2(n_120), .C1(n_118), .C2(n_304), .Y(n_383) );
AND2x2_ASAP7_75t_L g384 ( .A(n_354), .B(n_316), .Y(n_384) );
AOI22xp33_ASAP7_75t_L g385 ( .A1(n_341), .A2(n_300), .B1(n_359), .B2(n_327), .Y(n_385) );
AND2x2_ASAP7_75t_L g386 ( .A(n_354), .B(n_6), .Y(n_386) );
NAND2xp5_ASAP7_75t_L g387 ( .A(n_329), .B(n_300), .Y(n_387) );
AND2x2_ASAP7_75t_L g388 ( .A(n_350), .B(n_6), .Y(n_388) );
NAND2xp5_ASAP7_75t_L g389 ( .A(n_339), .B(n_345), .Y(n_389) );
INVx2_ASAP7_75t_L g390 ( .A(n_330), .Y(n_390) );
INVx1_ASAP7_75t_L g391 ( .A(n_339), .Y(n_391) );
A2O1A1Ixp33_ASAP7_75t_L g392 ( .A1(n_326), .A2(n_122), .B(n_120), .C(n_217), .Y(n_392) );
OAI22xp5_ASAP7_75t_SL g393 ( .A1(n_346), .A2(n_7), .B1(n_9), .B2(n_10), .Y(n_393) );
AND2x2_ASAP7_75t_L g394 ( .A(n_351), .B(n_7), .Y(n_394) );
OAI32xp33_ASAP7_75t_L g395 ( .A1(n_365), .A2(n_11), .A3(n_12), .B1(n_13), .B2(n_14), .Y(n_395) );
HB1xp67_ASAP7_75t_L g396 ( .A(n_330), .Y(n_396) );
AND2x2_ASAP7_75t_L g397 ( .A(n_351), .B(n_11), .Y(n_397) );
INVx1_ASAP7_75t_L g398 ( .A(n_352), .Y(n_398) );
AOI32xp33_ASAP7_75t_L g399 ( .A1(n_356), .A2(n_12), .A3(n_14), .B1(n_15), .B2(n_16), .Y(n_399) );
NOR2x1p5_ASAP7_75t_L g400 ( .A(n_347), .B(n_122), .Y(n_400) );
NAND4xp25_ASAP7_75t_L g401 ( .A(n_362), .B(n_15), .C(n_17), .D(n_18), .Y(n_401) );
NAND2xp5_ASAP7_75t_L g402 ( .A(n_345), .B(n_122), .Y(n_402) );
NOR2xp33_ASAP7_75t_R g403 ( .A(n_356), .B(n_20), .Y(n_403) );
INVx1_ASAP7_75t_L g404 ( .A(n_352), .Y(n_404) );
OR2x2_ASAP7_75t_L g405 ( .A(n_362), .B(n_120), .Y(n_405) );
INVx1_ASAP7_75t_SL g406 ( .A(n_346), .Y(n_406) );
NAND2xp5_ASAP7_75t_L g407 ( .A(n_349), .B(n_21), .Y(n_407) );
AND2x4_ASAP7_75t_L g408 ( .A(n_346), .B(n_22), .Y(n_408) );
BUFx2_ASAP7_75t_L g409 ( .A(n_346), .Y(n_409) );
NAND2x1p5_ASAP7_75t_L g410 ( .A(n_360), .B(n_183), .Y(n_410) );
NAND2xp5_ASAP7_75t_L g411 ( .A(n_370), .B(n_364), .Y(n_411) );
OAI21xp5_ASAP7_75t_L g412 ( .A1(n_401), .A2(n_361), .B(n_360), .Y(n_412) );
INVx1_ASAP7_75t_L g413 ( .A(n_391), .Y(n_413) );
NAND2xp5_ASAP7_75t_L g414 ( .A(n_370), .B(n_364), .Y(n_414) );
NAND2xp5_ASAP7_75t_L g415 ( .A(n_398), .B(n_340), .Y(n_415) );
INVx1_ASAP7_75t_L g416 ( .A(n_389), .Y(n_416) );
AOI31xp33_ASAP7_75t_L g417 ( .A1(n_380), .A2(n_336), .A3(n_328), .B(n_338), .Y(n_417) );
INVx2_ASAP7_75t_SL g418 ( .A(n_382), .Y(n_418) );
INVx1_ASAP7_75t_L g419 ( .A(n_389), .Y(n_419) );
AOI21xp5_ASAP7_75t_L g420 ( .A1(n_380), .A2(n_349), .B(n_357), .Y(n_420) );
A2O1A1Ixp33_ASAP7_75t_L g421 ( .A1(n_385), .A2(n_338), .B(n_328), .C(n_340), .Y(n_421) );
OR2x2_ASAP7_75t_L g422 ( .A(n_367), .B(n_357), .Y(n_422) );
NAND2xp5_ASAP7_75t_L g423 ( .A(n_404), .B(n_372), .Y(n_423) );
AND2x2_ASAP7_75t_L g424 ( .A(n_381), .B(n_355), .Y(n_424) );
INVxp67_ASAP7_75t_L g425 ( .A(n_371), .Y(n_425) );
NAND3xp33_ASAP7_75t_L g426 ( .A(n_385), .B(n_361), .C(n_343), .Y(n_426) );
OAI21xp33_ASAP7_75t_L g427 ( .A1(n_368), .A2(n_343), .B(n_335), .Y(n_427) );
NAND4xp25_ASAP7_75t_L g428 ( .A(n_399), .B(n_343), .C(n_335), .D(n_334), .Y(n_428) );
AND2x2_ASAP7_75t_L g429 ( .A(n_381), .B(n_335), .Y(n_429) );
XOR2x2_ASAP7_75t_L g430 ( .A(n_393), .B(n_23), .Y(n_430) );
OR2x2_ASAP7_75t_L g431 ( .A(n_376), .B(n_24), .Y(n_431) );
NOR2xp33_ASAP7_75t_SL g432 ( .A(n_408), .B(n_183), .Y(n_432) );
HB1xp67_ASAP7_75t_L g433 ( .A(n_396), .Y(n_433) );
INVxp67_ASAP7_75t_L g434 ( .A(n_371), .Y(n_434) );
NOR2xp33_ASAP7_75t_L g435 ( .A(n_387), .B(n_25), .Y(n_435) );
NOR2xp33_ASAP7_75t_L g436 ( .A(n_387), .B(n_26), .Y(n_436) );
INVx1_ASAP7_75t_SL g437 ( .A(n_403), .Y(n_437) );
NAND2xp5_ASAP7_75t_L g438 ( .A(n_377), .B(n_29), .Y(n_438) );
AND2x2_ASAP7_75t_L g439 ( .A(n_409), .B(n_30), .Y(n_439) );
OR2x2_ASAP7_75t_L g440 ( .A(n_369), .B(n_373), .Y(n_440) );
AOI21xp5_ASAP7_75t_L g441 ( .A1(n_383), .A2(n_164), .B(n_162), .Y(n_441) );
XNOR2x1_ASAP7_75t_L g442 ( .A(n_374), .B(n_32), .Y(n_442) );
NAND2xp5_ASAP7_75t_L g443 ( .A(n_379), .B(n_34), .Y(n_443) );
AND2x2_ASAP7_75t_L g444 ( .A(n_406), .B(n_36), .Y(n_444) );
XNOR2xp5_ASAP7_75t_L g445 ( .A(n_386), .B(n_38), .Y(n_445) );
NAND2xp5_ASAP7_75t_L g446 ( .A(n_390), .B(n_41), .Y(n_446) );
NAND2xp5_ASAP7_75t_L g447 ( .A(n_384), .B(n_44), .Y(n_447) );
NAND2xp5_ASAP7_75t_L g448 ( .A(n_405), .B(n_45), .Y(n_448) );
AOI21xp33_ASAP7_75t_SL g449 ( .A1(n_408), .A2(n_46), .B(n_47), .Y(n_449) );
NAND2xp5_ASAP7_75t_L g450 ( .A(n_388), .B(n_48), .Y(n_450) );
HB1xp67_ASAP7_75t_L g451 ( .A(n_402), .Y(n_451) );
AOI211xp5_ASAP7_75t_L g452 ( .A1(n_403), .A2(n_164), .B(n_162), .C(n_55), .Y(n_452) );
OAI211xp5_ASAP7_75t_L g453 ( .A1(n_395), .A2(n_183), .B(n_176), .C(n_163), .Y(n_453) );
INVx1_ASAP7_75t_L g454 ( .A(n_402), .Y(n_454) );
NAND4xp75_ASAP7_75t_L g455 ( .A(n_394), .B(n_51), .C(n_54), .D(n_56), .Y(n_455) );
OAI21xp33_ASAP7_75t_L g456 ( .A1(n_397), .A2(n_190), .B(n_168), .Y(n_456) );
A2O1A1Ixp33_ASAP7_75t_L g457 ( .A1(n_400), .A2(n_59), .B(n_61), .C(n_62), .Y(n_457) );
INVx3_ASAP7_75t_L g458 ( .A(n_410), .Y(n_458) );
XNOR2x1_ASAP7_75t_L g459 ( .A(n_410), .B(n_67), .Y(n_459) );
INVx1_ASAP7_75t_L g460 ( .A(n_407), .Y(n_460) );
INVx2_ASAP7_75t_SL g461 ( .A(n_407), .Y(n_461) );
XNOR2x1_ASAP7_75t_L g462 ( .A(n_378), .B(n_70), .Y(n_462) );
NAND2xp5_ASAP7_75t_SL g463 ( .A(n_392), .B(n_162), .Y(n_463) );
O2A1O1Ixp5_ASAP7_75t_SL g464 ( .A1(n_380), .A2(n_72), .B(n_74), .C(n_75), .Y(n_464) );
INVx2_ASAP7_75t_L g465 ( .A(n_396), .Y(n_465) );
INVx1_ASAP7_75t_L g466 ( .A(n_391), .Y(n_466) );
AND2x2_ASAP7_75t_L g467 ( .A(n_375), .B(n_76), .Y(n_467) );
NAND2x1p5_ASAP7_75t_L g468 ( .A(n_408), .B(n_162), .Y(n_468) );
A2O1A1Ixp33_ASAP7_75t_L g469 ( .A1(n_380), .A2(n_162), .B(n_164), .C(n_168), .Y(n_469) );
XNOR2x1_ASAP7_75t_L g470 ( .A(n_374), .B(n_162), .Y(n_470) );
INVx1_ASAP7_75t_L g471 ( .A(n_391), .Y(n_471) );
AOI22xp33_ASAP7_75t_SL g472 ( .A1(n_403), .A2(n_164), .B1(n_190), .B2(n_409), .Y(n_472) );
OAI22xp33_ASAP7_75t_L g473 ( .A1(n_380), .A2(n_164), .B1(n_401), .B2(n_346), .Y(n_473) );
INVx1_ASAP7_75t_L g474 ( .A(n_416), .Y(n_474) );
NOR2x1_ASAP7_75t_SL g475 ( .A(n_418), .B(n_426), .Y(n_475) );
OAI211xp5_ASAP7_75t_L g476 ( .A1(n_437), .A2(n_472), .B(n_421), .C(n_427), .Y(n_476) );
INVx1_ASAP7_75t_L g477 ( .A(n_419), .Y(n_477) );
NAND2xp5_ASAP7_75t_L g478 ( .A(n_425), .B(n_434), .Y(n_478) );
NAND2xp5_ASAP7_75t_L g479 ( .A(n_425), .B(n_434), .Y(n_479) );
AOI211xp5_ASAP7_75t_SL g480 ( .A1(n_473), .A2(n_417), .B(n_432), .C(n_452), .Y(n_480) );
AOI22xp5_ASAP7_75t_L g481 ( .A1(n_473), .A2(n_421), .B1(n_428), .B2(n_423), .Y(n_481) );
INVxp67_ASAP7_75t_L g482 ( .A(n_433), .Y(n_482) );
NOR2x1_ASAP7_75t_L g483 ( .A(n_459), .B(n_469), .Y(n_483) );
INVx2_ASAP7_75t_SL g484 ( .A(n_440), .Y(n_484) );
AOI21xp5_ASAP7_75t_L g485 ( .A1(n_420), .A2(n_469), .B(n_463), .Y(n_485) );
INVx1_ASAP7_75t_L g486 ( .A(n_424), .Y(n_486) );
AOI22xp33_ASAP7_75t_L g487 ( .A1(n_430), .A2(n_436), .B1(n_435), .B2(n_451), .Y(n_487) );
OAI221xp5_ASAP7_75t_L g488 ( .A1(n_472), .A2(n_442), .B1(n_462), .B2(n_470), .C(n_430), .Y(n_488) );
NAND2xp5_ASAP7_75t_L g489 ( .A(n_451), .B(n_460), .Y(n_489) );
AOI22xp33_ASAP7_75t_L g490 ( .A1(n_442), .A2(n_458), .B1(n_461), .B2(n_454), .Y(n_490) );
AOI22xp5_ASAP7_75t_L g491 ( .A1(n_435), .A2(n_436), .B1(n_415), .B2(n_414), .Y(n_491) );
OAI211xp5_ASAP7_75t_L g492 ( .A1(n_490), .A2(n_449), .B(n_456), .C(n_447), .Y(n_492) );
INVx2_ASAP7_75t_L g493 ( .A(n_484), .Y(n_493) );
NAND4xp25_ASAP7_75t_L g494 ( .A(n_480), .B(n_488), .C(n_487), .D(n_483), .Y(n_494) );
OAI221xp5_ASAP7_75t_SL g495 ( .A1(n_487), .A2(n_445), .B1(n_443), .B2(n_438), .C(n_450), .Y(n_495) );
NAND4xp25_ASAP7_75t_L g496 ( .A(n_481), .B(n_439), .C(n_412), .D(n_457), .Y(n_496) );
NOR3xp33_ASAP7_75t_SL g497 ( .A(n_476), .B(n_453), .C(n_455), .Y(n_497) );
OAI211xp5_ASAP7_75t_SL g498 ( .A1(n_485), .A2(n_457), .B(n_453), .C(n_463), .Y(n_498) );
NAND3xp33_ASAP7_75t_L g499 ( .A(n_482), .B(n_464), .C(n_433), .Y(n_499) );
INVx1_ASAP7_75t_L g500 ( .A(n_489), .Y(n_500) );
OAI21xp5_ASAP7_75t_L g501 ( .A1(n_482), .A2(n_468), .B(n_458), .Y(n_501) );
INVx1_ASAP7_75t_SL g502 ( .A(n_493), .Y(n_502) );
OAI22xp5_ASAP7_75t_SL g503 ( .A1(n_494), .A2(n_475), .B1(n_468), .B2(n_491), .Y(n_503) );
NOR3xp33_ASAP7_75t_L g504 ( .A(n_499), .B(n_448), .C(n_479), .Y(n_504) );
AOI22xp5_ASAP7_75t_L g505 ( .A1(n_496), .A2(n_478), .B1(n_486), .B2(n_477), .Y(n_505) );
AOI211xp5_ASAP7_75t_SL g506 ( .A1(n_492), .A2(n_444), .B(n_467), .C(n_431), .Y(n_506) );
OR3x1_ASAP7_75t_L g507 ( .A(n_503), .B(n_498), .C(n_500), .Y(n_507) );
OR4x2_ASAP7_75t_L g508 ( .A(n_506), .B(n_495), .C(n_497), .D(n_501), .Y(n_508) );
NAND4xp25_ASAP7_75t_L g509 ( .A(n_504), .B(n_441), .C(n_446), .D(n_474), .Y(n_509) );
NOR3xp33_ASAP7_75t_L g510 ( .A(n_509), .B(n_502), .C(n_505), .Y(n_510) );
INVxp67_ASAP7_75t_SL g511 ( .A(n_507), .Y(n_511) );
OR3x2_ASAP7_75t_L g512 ( .A(n_511), .B(n_508), .C(n_422), .Y(n_512) );
NOR2xp67_ASAP7_75t_L g513 ( .A(n_512), .B(n_510), .Y(n_513) );
O2A1O1Ixp33_ASAP7_75t_L g514 ( .A1(n_513), .A2(n_471), .B(n_466), .C(n_413), .Y(n_514) );
AOI22xp33_ASAP7_75t_L g515 ( .A1(n_514), .A2(n_429), .B1(n_411), .B2(n_465), .Y(n_515) );
endmodule