module real_aes_2539_n_77 (n_17, n_28, n_76, n_56, n_34, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_43, n_54, n_35, n_42, n_15, n_9, n_23, n_72, n_44, n_7, n_4, n_6, n_12, n_68, n_69, n_46, n_59, n_25, n_73, n_48, n_37, n_70, n_50, n_26, n_13, n_24, n_2, n_55, n_62, n_67, n_33, n_14, n_11, n_16, n_39, n_5, n_45, n_60, n_38, n_0, n_63, n_1, n_53, n_36, n_77);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_43;
input n_54;
input n_35;
input n_42;
input n_15;
input n_9;
input n_23;
input n_72;
input n_44;
input n_7;
input n_4;
input n_6;
input n_12;
input n_68;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_48;
input n_37;
input n_70;
input n_50;
input n_26;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_67;
input n_33;
input n_14;
input n_11;
input n_16;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_0;
input n_63;
input n_1;
input n_53;
input n_36;
output n_77;
wire n_480;
wire n_113;
wire n_476;
wire n_187;
wire n_436;
wire n_90;
wire n_257;
wire n_390;
wire n_185;
wire n_285;
wire n_522;
wire n_485;
wire n_222;
wire n_287;
wire n_357;
wire n_503;
wire n_386;
wire n_518;
wire n_254;
wire n_207;
wire n_469;
wire n_83;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_445;
wire n_540;
wire n_299;
wire n_322;
wire n_328;
wire n_318;
wire n_355;
wire n_239;
wire n_100;
wire n_423;
wire n_458;
wire n_444;
wire n_112;
wire n_319;
wire n_421;
wire n_364;
wire n_329;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_169;
wire n_242;
wire n_376;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_448;
wire n_545;
wire n_341;
wire n_232;
wire n_460;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_537;
wire n_320;
wire n_260;
wire n_97;
wire n_186;
wire n_138;
wire n_379;
wire n_374;
wire n_453;
wire n_235;
wire n_399;
wire n_378;
wire n_245;
wire n_161;
wire n_189;
wire n_271;
wire n_489;
wire n_427;
wire n_145;
wire n_415;
wire n_227;
wire n_92;
wire n_519;
wire n_510;
wire n_330;
wire n_388;
wire n_512;
wire n_395;
wire n_332;
wire n_292;
wire n_539;
wire n_400;
wire n_116;
wire n_94;
wire n_289;
wire n_462;
wire n_280;
wire n_333;
wire n_213;
wire n_478;
wire n_356;
wire n_408;
wire n_184;
wire n_372;
wire n_528;
wire n_202;
wire n_495;
wire n_370;
wire n_98;
wire n_384;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_82;
wire n_467;
wire n_327;
wire n_106;
wire n_466;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_517;
wire n_174;
wire n_530;
wire n_104;
wire n_535;
wire n_211;
wire n_281;
wire n_496;
wire n_173;
wire n_468;
wire n_234;
wire n_284;
wire n_153;
wire n_316;
wire n_532;
wire n_178;
wire n_409;
wire n_298;
wire n_523;
wire n_439;
wire n_506;
wire n_513;
wire n_297;
wire n_383;
wire n_529;
wire n_119;
wire n_310;
wire n_455;
wire n_504;
wire n_164;
wire n_231;
wire n_102;
wire n_454;
wire n_122;
wire n_443;
wire n_534;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_80;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_367;
wire n_267;
wire n_218;
wire n_204;
wire n_339;
wire n_398;
wire n_89;
wire n_277;
wire n_425;
wire n_331;
wire n_93;
wire n_182;
wire n_363;
wire n_417;
wire n_449;
wire n_323;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_142;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_368;
wire n_527;
wire n_434;
wire n_502;
wire n_505;
wire n_250;
wire n_85;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_402;
wire n_171;
wire n_87;
wire n_78;
wire n_531;
wire n_451;
wire n_146;
wire n_432;
wire n_226;
wire n_255;
wire n_286;
wire n_416;
wire n_410;
wire n_120;
wire n_490;
wire n_261;
wire n_238;
wire n_391;
wire n_360;
wire n_165;
wire n_361;
wire n_246;
wire n_176;
wire n_412;
wire n_163;
wire n_542;
wire n_488;
wire n_501;
wire n_251;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_115;
wire n_96;
wire n_110;
wire n_392;
wire n_150;
wire n_147;
wire n_288;
wire n_404;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_95;
wire n_188;
wire n_269;
wire n_430;
wire n_201;
wire n_413;
wire n_471;
wire n_306;
wire n_158;
wire n_533;
wire n_366;
wire n_346;
wire n_193;
wire n_397;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_109;
wire n_536;
wire n_203;
wire n_470;
wire n_81;
wire n_133;
wire n_494;
wire n_377;
wire n_273;
wire n_114;
wire n_276;
wire n_295;
wire n_382;
wire n_265;
wire n_354;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_486;
wire n_411;
wire n_291;
wire n_148;
wire n_481;
wire n_498;
wire n_88;
wire n_159;
wire n_108;
wire n_373;
wire n_233;
wire n_487;
wire n_290;
wire n_365;
wire n_526;
wire n_155;
wire n_243;
wire n_544;
wire n_268;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_101;
wire n_309;
wire n_344;
wire n_229;
wire n_107;
wire n_482;
wire n_520;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_262;
wire n_134;
wire n_349;
wire n_420;
wire n_336;
wire n_195;
wire n_438;
wire n_300;
wire n_252;
wire n_283;
wire n_314;
wire n_249;
wire n_446;
wire n_221;
wire n_156;
wire n_359;
wire n_456;
wire n_312;
wire n_183;
wire n_266;
wire n_205;
wire n_433;
wire n_335;
wire n_177;
wire n_516;
wire n_313;
wire n_140;
wire n_418;
wire n_521;
wire n_422;
wire n_219;
wire n_524;
wire n_180;
wire n_212;
wire n_210;
wire n_325;
wire n_338;
wire n_479;
wire n_442;
wire n_371;
wire n_103;
wire n_166;
wire n_541;
wire n_224;
wire n_151;
wire n_130;
wire n_253;
wire n_459;
wire n_99;
wire n_440;
wire n_525;
wire n_152;
wire n_198;
wire n_228;
wire n_272;
wire n_196;
wire n_347;
wire n_315;
wire n_414;
wire n_123;
wire n_279;
wire n_79;
wire n_543;
wire n_497;
wire n_514;
wire n_270;
wire n_507;
wire n_305;
wire n_450;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_465;
wire n_473;
wire n_474;
wire n_170;
wire n_86;
wire n_375;
wire n_340;
wire n_483;
wire n_380;
wire n_394;
wire n_168;
wire n_175;
wire n_241;
wire n_105;
wire n_84;
wire n_294;
wire n_393;
wire n_258;
wire n_206;
wire n_307;
wire n_500;
wire n_463;
wire n_396;
wire n_447;
wire n_342;
wire n_348;
wire n_403;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_143;
wire n_192;
wire n_475;
wire n_264;
wire n_237;
wire n_91;
AOI22xp33_ASAP7_75t_L g120 ( .A1(n_0), .A2(n_57), .B1(n_121), .B2(n_124), .Y(n_120) );
AOI22xp5_ASAP7_75t_L g149 ( .A1(n_1), .A2(n_150), .B1(n_151), .B2(n_152), .Y(n_149) );
INVx1_ASAP7_75t_L g150 ( .A(n_1), .Y(n_150) );
AO22x2_ASAP7_75t_L g102 ( .A1(n_2), .A2(n_52), .B1(n_92), .B2(n_103), .Y(n_102) );
INVx1_ASAP7_75t_L g168 ( .A(n_3), .Y(n_168) );
NAND2xp5_ASAP7_75t_SL g296 ( .A(n_4), .B(n_213), .Y(n_296) );
INVx1_ASAP7_75t_L g276 ( .A(n_5), .Y(n_276) );
AO22x2_ASAP7_75t_L g99 ( .A1(n_6), .A2(n_18), .B1(n_92), .B2(n_100), .Y(n_99) );
CKINVDCx5p33_ASAP7_75t_R g241 ( .A(n_7), .Y(n_241) );
AOI22xp5_ASAP7_75t_L g132 ( .A1(n_8), .A2(n_22), .B1(n_133), .B2(n_137), .Y(n_132) );
INVx2_ASAP7_75t_L g186 ( .A(n_9), .Y(n_186) );
AOI22xp5_ASAP7_75t_L g79 ( .A1(n_10), .A2(n_80), .B1(n_81), .B2(n_147), .Y(n_79) );
INVx1_ASAP7_75t_L g147 ( .A(n_10), .Y(n_147) );
INVx1_ASAP7_75t_L g305 ( .A(n_11), .Y(n_305) );
INVx1_ASAP7_75t_L g302 ( .A(n_12), .Y(n_302) );
INVx1_ASAP7_75t_SL g223 ( .A(n_13), .Y(n_223) );
NAND2xp5_ASAP7_75t_SL g292 ( .A(n_14), .B(n_201), .Y(n_292) );
AOI22xp5_ASAP7_75t_L g536 ( .A1(n_15), .A2(n_80), .B1(n_81), .B2(n_537), .Y(n_536) );
CKINVDCx20_ASAP7_75t_R g537 ( .A(n_15), .Y(n_537) );
AOI33xp33_ASAP7_75t_L g262 ( .A1(n_16), .A2(n_38), .A3(n_191), .B1(n_199), .B2(n_263), .B3(n_264), .Y(n_262) );
OAI22xp5_ASAP7_75t_SL g152 ( .A1(n_17), .A2(n_75), .B1(n_153), .B2(n_154), .Y(n_152) );
INVx1_ASAP7_75t_L g154 ( .A(n_17), .Y(n_154) );
OAI221xp5_ASAP7_75t_L g160 ( .A1(n_18), .A2(n_52), .B1(n_55), .B2(n_161), .C(n_163), .Y(n_160) );
OA21x2_ASAP7_75t_L g185 ( .A1(n_19), .A2(n_68), .B(n_186), .Y(n_185) );
OR2x2_ASAP7_75t_L g214 ( .A(n_19), .B(n_68), .Y(n_214) );
NAND2xp5_ASAP7_75t_L g220 ( .A(n_20), .B(n_209), .Y(n_220) );
INVx3_ASAP7_75t_L g92 ( .A(n_21), .Y(n_92) );
INVx1_ASAP7_75t_SL g93 ( .A(n_23), .Y(n_93) );
INVx1_ASAP7_75t_L g170 ( .A(n_24), .Y(n_170) );
AND2x2_ASAP7_75t_L g207 ( .A(n_24), .B(n_168), .Y(n_207) );
AND2x2_ASAP7_75t_L g212 ( .A(n_24), .B(n_193), .Y(n_212) );
CKINVDCx20_ASAP7_75t_R g236 ( .A(n_25), .Y(n_236) );
NAND2xp5_ASAP7_75t_L g248 ( .A(n_26), .B(n_209), .Y(n_248) );
INVx1_ASAP7_75t_L g545 ( .A(n_26), .Y(n_545) );
AOI22xp33_ASAP7_75t_L g104 ( .A1(n_27), .A2(n_37), .B1(n_105), .B2(n_109), .Y(n_104) );
AOI22xp33_ASAP7_75t_L g139 ( .A1(n_28), .A2(n_41), .B1(n_140), .B2(n_141), .Y(n_139) );
AOI22xp5_ASAP7_75t_L g285 ( .A1(n_29), .A2(n_184), .B1(n_213), .B2(n_286), .Y(n_285) );
NAND2xp5_ASAP7_75t_L g293 ( .A(n_30), .B(n_294), .Y(n_293) );
NAND2xp5_ASAP7_75t_L g224 ( .A(n_31), .B(n_201), .Y(n_224) );
NAND2xp5_ASAP7_75t_SL g278 ( .A(n_32), .B(n_257), .Y(n_278) );
NAND2xp5_ASAP7_75t_L g277 ( .A(n_33), .B(n_201), .Y(n_277) );
AOI22xp33_ASAP7_75t_SL g128 ( .A1(n_34), .A2(n_49), .B1(n_129), .B2(n_130), .Y(n_128) );
AO22x2_ASAP7_75t_L g95 ( .A1(n_35), .A2(n_55), .B1(n_92), .B2(n_96), .Y(n_95) );
CKINVDCx5p33_ASAP7_75t_R g289 ( .A(n_36), .Y(n_289) );
NAND2xp5_ASAP7_75t_L g252 ( .A(n_39), .B(n_201), .Y(n_252) );
AOI22xp5_ASAP7_75t_L g528 ( .A1(n_39), .A2(n_80), .B1(n_81), .B2(n_529), .Y(n_528) );
INVx1_ASAP7_75t_L g529 ( .A(n_39), .Y(n_529) );
INVx1_ASAP7_75t_L g195 ( .A(n_40), .Y(n_195) );
INVx1_ASAP7_75t_L g203 ( .A(n_40), .Y(n_203) );
AND2x2_ASAP7_75t_L g253 ( .A(n_42), .B(n_217), .Y(n_253) );
AOI221xp5_ASAP7_75t_L g274 ( .A1(n_43), .A2(n_59), .B1(n_189), .B2(n_209), .C(n_275), .Y(n_274) );
NAND2xp5_ASAP7_75t_L g208 ( .A(n_44), .B(n_209), .Y(n_208) );
INVx1_ASAP7_75t_L g94 ( .A(n_45), .Y(n_94) );
NAND2xp5_ASAP7_75t_L g243 ( .A(n_46), .B(n_184), .Y(n_243) );
AOI21xp5_ASAP7_75t_SL g188 ( .A1(n_47), .A2(n_189), .B(n_196), .Y(n_188) );
INVx1_ASAP7_75t_L g299 ( .A(n_48), .Y(n_299) );
INVx1_ASAP7_75t_L g251 ( .A(n_50), .Y(n_251) );
AOI21xp5_ASAP7_75t_L g249 ( .A1(n_51), .A2(n_189), .B(n_250), .Y(n_249) );
INVxp33_ASAP7_75t_L g165 ( .A(n_52), .Y(n_165) );
INVx1_ASAP7_75t_L g193 ( .A(n_53), .Y(n_193) );
INVx1_ASAP7_75t_L g205 ( .A(n_53), .Y(n_205) );
AOI22xp33_ASAP7_75t_SL g113 ( .A1(n_54), .A2(n_58), .B1(n_114), .B2(n_117), .Y(n_113) );
INVxp67_ASAP7_75t_L g164 ( .A(n_55), .Y(n_164) );
NAND2xp5_ASAP7_75t_L g265 ( .A(n_56), .B(n_209), .Y(n_265) );
AND2x2_ASAP7_75t_L g225 ( .A(n_60), .B(n_183), .Y(n_225) );
INVx1_ASAP7_75t_L g300 ( .A(n_61), .Y(n_300) );
AOI21xp5_ASAP7_75t_L g221 ( .A1(n_62), .A2(n_189), .B(n_222), .Y(n_221) );
A2O1A1Ixp33_ASAP7_75t_L g290 ( .A1(n_63), .A2(n_189), .B(n_256), .C(n_291), .Y(n_290) );
AND2x2_ASAP7_75t_SL g182 ( .A(n_64), .B(n_183), .Y(n_182) );
AOI22xp5_ASAP7_75t_L g259 ( .A1(n_65), .A2(n_189), .B1(n_260), .B2(n_261), .Y(n_259) );
AOI22xp5_ASAP7_75t_L g148 ( .A1(n_66), .A2(n_149), .B1(n_155), .B2(n_156), .Y(n_148) );
INVx1_ASAP7_75t_L g155 ( .A(n_66), .Y(n_155) );
AOI22xp33_ASAP7_75t_L g142 ( .A1(n_67), .A2(n_73), .B1(n_143), .B2(n_144), .Y(n_142) );
INVx1_ASAP7_75t_L g197 ( .A(n_69), .Y(n_197) );
AND2x2_ASAP7_75t_L g266 ( .A(n_70), .B(n_183), .Y(n_266) );
A2O1A1Ixp33_ASAP7_75t_L g231 ( .A1(n_71), .A2(n_232), .B(n_233), .C(n_235), .Y(n_231) );
NAND2xp5_ASAP7_75t_SL g85 ( .A(n_72), .B(n_86), .Y(n_85) );
BUFx2_ASAP7_75t_SL g162 ( .A(n_74), .Y(n_162) );
INVx1_ASAP7_75t_L g153 ( .A(n_75), .Y(n_153) );
NAND2xp5_ASAP7_75t_L g200 ( .A(n_76), .B(n_201), .Y(n_200) );
AOI221xp5_ASAP7_75t_L g77 ( .A1(n_78), .A2(n_157), .B1(n_171), .B2(n_525), .C(n_527), .Y(n_77) );
XOR2xp5_ASAP7_75t_L g78 ( .A(n_79), .B(n_148), .Y(n_78) );
CKINVDCx20_ASAP7_75t_R g80 ( .A(n_81), .Y(n_80) );
HB1xp67_ASAP7_75t_L g81 ( .A(n_82), .Y(n_81) );
NAND2x1_ASAP7_75t_L g82 ( .A(n_83), .B(n_126), .Y(n_82) );
NOR2x1_ASAP7_75t_L g83 ( .A(n_84), .B(n_112), .Y(n_83) );
NAND2xp5_ASAP7_75t_L g84 ( .A(n_85), .B(n_104), .Y(n_84) );
INVx4_ASAP7_75t_SL g86 ( .A(n_87), .Y(n_86) );
INVx6_ASAP7_75t_L g87 ( .A(n_88), .Y(n_87) );
AND2x2_ASAP7_75t_L g88 ( .A(n_89), .B(n_97), .Y(n_88) );
AND2x2_ASAP7_75t_L g117 ( .A(n_89), .B(n_118), .Y(n_117) );
AND2x2_ASAP7_75t_L g124 ( .A(n_89), .B(n_125), .Y(n_124) );
AND2x2_ASAP7_75t_L g89 ( .A(n_90), .B(n_95), .Y(n_89) );
AND2x2_ASAP7_75t_L g107 ( .A(n_90), .B(n_108), .Y(n_107) );
HB1xp67_ASAP7_75t_L g110 ( .A(n_90), .Y(n_110) );
INVx2_ASAP7_75t_L g123 ( .A(n_90), .Y(n_123) );
OAI22x1_ASAP7_75t_L g90 ( .A1(n_91), .A2(n_92), .B1(n_93), .B2(n_94), .Y(n_90) );
INVx1_ASAP7_75t_L g91 ( .A(n_92), .Y(n_91) );
INVx1_ASAP7_75t_L g96 ( .A(n_92), .Y(n_96) );
INVx2_ASAP7_75t_L g100 ( .A(n_92), .Y(n_100) );
INVx1_ASAP7_75t_L g103 ( .A(n_92), .Y(n_103) );
INVx2_ASAP7_75t_L g108 ( .A(n_95), .Y(n_108) );
AND2x2_ASAP7_75t_L g122 ( .A(n_95), .B(n_123), .Y(n_122) );
BUFx2_ASAP7_75t_L g131 ( .A(n_95), .Y(n_131) );
AND2x4_ASAP7_75t_L g135 ( .A(n_97), .B(n_136), .Y(n_135) );
AND2x2_ASAP7_75t_L g140 ( .A(n_97), .B(n_107), .Y(n_140) );
AND2x6_ASAP7_75t_L g143 ( .A(n_97), .B(n_122), .Y(n_143) );
AND2x4_ASAP7_75t_L g97 ( .A(n_98), .B(n_101), .Y(n_97) );
INVx1_ASAP7_75t_L g98 ( .A(n_99), .Y(n_98) );
AND2x4_ASAP7_75t_L g106 ( .A(n_99), .B(n_101), .Y(n_106) );
AND2x2_ASAP7_75t_L g111 ( .A(n_99), .B(n_102), .Y(n_111) );
INVx1_ASAP7_75t_L g116 ( .A(n_99), .Y(n_116) );
INVxp67_ASAP7_75t_L g125 ( .A(n_101), .Y(n_125) );
INVx2_ASAP7_75t_L g101 ( .A(n_102), .Y(n_101) );
AND2x2_ASAP7_75t_L g115 ( .A(n_102), .B(n_116), .Y(n_115) );
AND2x4_ASAP7_75t_L g105 ( .A(n_106), .B(n_107), .Y(n_105) );
AND2x2_ASAP7_75t_L g121 ( .A(n_106), .B(n_122), .Y(n_121) );
AND2x4_ASAP7_75t_L g146 ( .A(n_106), .B(n_136), .Y(n_146) );
AND2x4_ASAP7_75t_L g114 ( .A(n_107), .B(n_115), .Y(n_114) );
AND2x4_ASAP7_75t_L g136 ( .A(n_108), .B(n_123), .Y(n_136) );
AND2x2_ASAP7_75t_SL g109 ( .A(n_110), .B(n_111), .Y(n_109) );
AND2x4_ASAP7_75t_L g130 ( .A(n_111), .B(n_131), .Y(n_130) );
AND2x4_ASAP7_75t_L g141 ( .A(n_111), .B(n_136), .Y(n_141) );
NAND2xp5_ASAP7_75t_L g112 ( .A(n_113), .B(n_120), .Y(n_112) );
AND2x2_ASAP7_75t_SL g129 ( .A(n_115), .B(n_122), .Y(n_129) );
AND2x6_ASAP7_75t_L g137 ( .A(n_115), .B(n_136), .Y(n_137) );
HB1xp67_ASAP7_75t_L g119 ( .A(n_116), .Y(n_119) );
INVx1_ASAP7_75t_L g118 ( .A(n_119), .Y(n_118) );
NOR2x1_ASAP7_75t_L g126 ( .A(n_127), .B(n_138), .Y(n_126) );
NAND2xp5_ASAP7_75t_L g127 ( .A(n_128), .B(n_132), .Y(n_127) );
INVx3_ASAP7_75t_L g133 ( .A(n_134), .Y(n_133) );
INVx8_ASAP7_75t_L g134 ( .A(n_135), .Y(n_134) );
NAND2xp5_ASAP7_75t_L g138 ( .A(n_139), .B(n_142), .Y(n_138) );
INVx1_ASAP7_75t_L g144 ( .A(n_145), .Y(n_144) );
INVx2_ASAP7_75t_L g145 ( .A(n_146), .Y(n_145) );
CKINVDCx20_ASAP7_75t_R g156 ( .A(n_149), .Y(n_156) );
CKINVDCx20_ASAP7_75t_R g151 ( .A(n_152), .Y(n_151) );
NOR2xp33_ASAP7_75t_L g233 ( .A(n_154), .B(n_234), .Y(n_233) );
INVx1_ASAP7_75t_SL g157 ( .A(n_158), .Y(n_157) );
CKINVDCx20_ASAP7_75t_R g158 ( .A(n_159), .Y(n_158) );
AND3x1_ASAP7_75t_SL g159 ( .A(n_160), .B(n_166), .C(n_169), .Y(n_159) );
INVxp67_ASAP7_75t_L g535 ( .A(n_160), .Y(n_535) );
CKINVDCx8_ASAP7_75t_R g161 ( .A(n_162), .Y(n_161) );
NOR2xp33_ASAP7_75t_L g163 ( .A(n_164), .B(n_165), .Y(n_163) );
CKINVDCx16_ASAP7_75t_R g533 ( .A(n_166), .Y(n_533) );
AOI21xp33_ASAP7_75t_L g542 ( .A1(n_166), .A2(n_543), .B(n_544), .Y(n_542) );
INVx1_ASAP7_75t_L g166 ( .A(n_167), .Y(n_166) );
AND2x2_ASAP7_75t_L g210 ( .A(n_167), .B(n_199), .Y(n_210) );
OR2x2_ASAP7_75t_SL g540 ( .A(n_167), .B(n_169), .Y(n_540) );
HB1xp67_ASAP7_75t_L g167 ( .A(n_168), .Y(n_167) );
AND2x2_ASAP7_75t_L g194 ( .A(n_168), .B(n_195), .Y(n_194) );
NAND2xp5_ASAP7_75t_L g534 ( .A(n_169), .B(n_535), .Y(n_534) );
INVx1_ASAP7_75t_L g169 ( .A(n_170), .Y(n_169) );
NOR2x1p5_ASAP7_75t_L g190 ( .A(n_170), .B(n_191), .Y(n_190) );
HB1xp67_ASAP7_75t_L g171 ( .A(n_172), .Y(n_171) );
INVx1_ASAP7_75t_SL g172 ( .A(n_173), .Y(n_172) );
AND3x2_ASAP7_75t_L g173 ( .A(n_174), .B(n_415), .C(n_478), .Y(n_173) );
INVx1_ASAP7_75t_L g174 ( .A(n_175), .Y(n_174) );
NAND2xp5_ASAP7_75t_L g175 ( .A(n_176), .B(n_379), .Y(n_175) );
NOR3xp33_ASAP7_75t_L g176 ( .A(n_177), .B(n_320), .C(n_349), .Y(n_176) );
NAND2xp5_ASAP7_75t_SL g177 ( .A(n_178), .B(n_309), .Y(n_177) );
AOI22xp5_ASAP7_75t_L g178 ( .A1(n_179), .A2(n_226), .B1(n_267), .B2(n_279), .Y(n_178) );
NAND2x1_ASAP7_75t_L g464 ( .A(n_179), .B(n_310), .Y(n_464) );
INVx2_ASAP7_75t_SL g179 ( .A(n_180), .Y(n_179) );
OR2x2_ASAP7_75t_L g180 ( .A(n_181), .B(n_215), .Y(n_180) );
INVx2_ASAP7_75t_L g281 ( .A(n_181), .Y(n_281) );
INVx4_ASAP7_75t_L g325 ( .A(n_181), .Y(n_325) );
BUFx6f_ASAP7_75t_L g345 ( .A(n_181), .Y(n_345) );
AND2x4_ASAP7_75t_L g356 ( .A(n_181), .B(n_324), .Y(n_356) );
AND2x2_ASAP7_75t_L g362 ( .A(n_181), .B(n_284), .Y(n_362) );
NOR2x1_ASAP7_75t_SL g492 ( .A(n_181), .B(n_295), .Y(n_492) );
OR2x6_ASAP7_75t_L g181 ( .A(n_182), .B(n_187), .Y(n_181) );
OAI22xp5_ASAP7_75t_L g230 ( .A1(n_183), .A2(n_231), .B1(n_236), .B2(n_237), .Y(n_230) );
INVx3_ASAP7_75t_L g237 ( .A(n_183), .Y(n_237) );
INVx4_ASAP7_75t_L g183 ( .A(n_184), .Y(n_183) );
NAND2xp5_ASAP7_75t_L g239 ( .A(n_184), .B(n_240), .Y(n_239) );
INVx3_ASAP7_75t_L g184 ( .A(n_185), .Y(n_184) );
BUFx4f_ASAP7_75t_L g257 ( .A(n_185), .Y(n_257) );
AND2x4_ASAP7_75t_L g213 ( .A(n_186), .B(n_214), .Y(n_213) );
AND2x2_ASAP7_75t_SL g218 ( .A(n_186), .B(n_214), .Y(n_218) );
AOI21xp5_ASAP7_75t_L g187 ( .A1(n_188), .A2(n_208), .B(n_213), .Y(n_187) );
INVxp67_ASAP7_75t_L g242 ( .A(n_189), .Y(n_242) );
AND2x4_ASAP7_75t_L g189 ( .A(n_190), .B(n_194), .Y(n_189) );
INVx1_ASAP7_75t_L g264 ( .A(n_191), .Y(n_264) );
INVx3_ASAP7_75t_L g191 ( .A(n_192), .Y(n_191) );
OR2x6_ASAP7_75t_L g198 ( .A(n_192), .B(n_199), .Y(n_198) );
INVx2_ASAP7_75t_L g192 ( .A(n_193), .Y(n_192) );
AND2x6_ASAP7_75t_L g304 ( .A(n_193), .B(n_202), .Y(n_304) );
INVx2_ASAP7_75t_L g199 ( .A(n_195), .Y(n_199) );
AND2x4_ASAP7_75t_L g307 ( .A(n_195), .B(n_204), .Y(n_307) );
O2A1O1Ixp33_ASAP7_75t_L g196 ( .A1(n_197), .A2(n_198), .B(n_200), .C(n_206), .Y(n_196) );
O2A1O1Ixp33_ASAP7_75t_SL g222 ( .A1(n_198), .A2(n_206), .B(n_223), .C(n_224), .Y(n_222) );
INVxp67_ASAP7_75t_L g232 ( .A(n_198), .Y(n_232) );
O2A1O1Ixp33_ASAP7_75t_L g250 ( .A1(n_198), .A2(n_206), .B(n_251), .C(n_252), .Y(n_250) );
O2A1O1Ixp33_ASAP7_75t_SL g275 ( .A1(n_198), .A2(n_206), .B(n_276), .C(n_277), .Y(n_275) );
INVx2_ASAP7_75t_L g294 ( .A(n_198), .Y(n_294) );
OAI22xp5_ASAP7_75t_L g298 ( .A1(n_198), .A2(n_234), .B1(n_299), .B2(n_300), .Y(n_298) );
INVxp33_ASAP7_75t_L g263 ( .A(n_199), .Y(n_263) );
HB1xp67_ASAP7_75t_L g543 ( .A(n_199), .Y(n_543) );
INVx1_ASAP7_75t_L g234 ( .A(n_201), .Y(n_234) );
AND2x4_ASAP7_75t_L g201 ( .A(n_202), .B(n_204), .Y(n_201) );
INVx2_ASAP7_75t_L g202 ( .A(n_203), .Y(n_202) );
INVx2_ASAP7_75t_L g204 ( .A(n_205), .Y(n_204) );
INVx1_ASAP7_75t_L g260 ( .A(n_206), .Y(n_260) );
AOI21xp5_ASAP7_75t_L g291 ( .A1(n_206), .A2(n_292), .B(n_293), .Y(n_291) );
NOR2xp33_ASAP7_75t_L g308 ( .A(n_206), .B(n_213), .Y(n_308) );
INVx5_ASAP7_75t_L g206 ( .A(n_207), .Y(n_206) );
HB1xp67_ASAP7_75t_L g235 ( .A(n_207), .Y(n_235) );
INVx1_ASAP7_75t_L g244 ( .A(n_209), .Y(n_244) );
AND2x4_ASAP7_75t_L g209 ( .A(n_210), .B(n_211), .Y(n_209) );
INVx1_ASAP7_75t_L g287 ( .A(n_210), .Y(n_287) );
INVx1_ASAP7_75t_L g288 ( .A(n_211), .Y(n_288) );
BUFx3_ASAP7_75t_L g211 ( .A(n_212), .Y(n_211) );
INVx2_ASAP7_75t_L g328 ( .A(n_215), .Y(n_328) );
HB1xp67_ASAP7_75t_L g342 ( .A(n_215), .Y(n_342) );
INVx1_ASAP7_75t_L g353 ( .A(n_215), .Y(n_353) );
HB1xp67_ASAP7_75t_L g365 ( .A(n_215), .Y(n_365) );
AND2x2_ASAP7_75t_L g397 ( .A(n_215), .B(n_295), .Y(n_397) );
AND2x2_ASAP7_75t_L g429 ( .A(n_215), .B(n_313), .Y(n_429) );
INVx1_ASAP7_75t_L g436 ( .A(n_215), .Y(n_436) );
AO21x2_ASAP7_75t_L g215 ( .A1(n_216), .A2(n_219), .B(n_225), .Y(n_215) );
CKINVDCx5p33_ASAP7_75t_R g216 ( .A(n_217), .Y(n_216) );
BUFx6f_ASAP7_75t_L g217 ( .A(n_218), .Y(n_217) );
NAND2xp5_ASAP7_75t_L g219 ( .A(n_220), .B(n_221), .Y(n_219) );
AND2x2_ASAP7_75t_L g226 ( .A(n_227), .B(n_245), .Y(n_226) );
INVx1_ASAP7_75t_L g227 ( .A(n_228), .Y(n_227) );
AND2x2_ASAP7_75t_L g378 ( .A(n_228), .B(n_317), .Y(n_378) );
INVx2_ASAP7_75t_L g452 ( .A(n_228), .Y(n_452) );
AND2x2_ASAP7_75t_L g475 ( .A(n_228), .B(n_245), .Y(n_475) );
INVx1_ASAP7_75t_L g228 ( .A(n_229), .Y(n_228) );
NAND2xp5_ASAP7_75t_L g316 ( .A(n_229), .B(n_270), .Y(n_316) );
INVx2_ASAP7_75t_L g337 ( .A(n_229), .Y(n_337) );
AND2x4_ASAP7_75t_L g359 ( .A(n_229), .B(n_360), .Y(n_359) );
INVx1_ASAP7_75t_L g394 ( .A(n_229), .Y(n_394) );
AND2x2_ASAP7_75t_L g471 ( .A(n_229), .B(n_273), .Y(n_471) );
OR2x2_ASAP7_75t_L g229 ( .A(n_230), .B(n_238), .Y(n_229) );
AO21x2_ASAP7_75t_L g246 ( .A1(n_237), .A2(n_247), .B(n_253), .Y(n_246) );
AO21x2_ASAP7_75t_L g270 ( .A1(n_237), .A2(n_247), .B(n_253), .Y(n_270) );
OAI22xp5_ASAP7_75t_L g238 ( .A1(n_239), .A2(n_242), .B1(n_243), .B2(n_244), .Y(n_238) );
INVx1_ASAP7_75t_L g240 ( .A(n_241), .Y(n_240) );
HB1xp67_ASAP7_75t_L g526 ( .A(n_244), .Y(n_526) );
INVx1_ASAP7_75t_L g442 ( .A(n_245), .Y(n_442) );
AND2x2_ASAP7_75t_L g245 ( .A(n_246), .B(n_254), .Y(n_245) );
NOR2xp67_ASAP7_75t_L g367 ( .A(n_246), .B(n_337), .Y(n_367) );
AND2x2_ASAP7_75t_L g372 ( .A(n_246), .B(n_337), .Y(n_372) );
INVx2_ASAP7_75t_L g385 ( .A(n_246), .Y(n_385) );
NOR2x1_ASAP7_75t_L g433 ( .A(n_246), .B(n_434), .Y(n_433) );
NAND2xp5_ASAP7_75t_L g247 ( .A(n_248), .B(n_249), .Y(n_247) );
AND2x4_ASAP7_75t_L g358 ( .A(n_254), .B(n_269), .Y(n_358) );
AND2x2_ASAP7_75t_L g373 ( .A(n_254), .B(n_374), .Y(n_373) );
INVx1_ASAP7_75t_L g426 ( .A(n_254), .Y(n_426) );
INVx2_ASAP7_75t_L g254 ( .A(n_255), .Y(n_254) );
NAND2xp5_ASAP7_75t_L g348 ( .A(n_255), .B(n_273), .Y(n_348) );
NAND2xp5_ASAP7_75t_L g430 ( .A(n_255), .B(n_270), .Y(n_430) );
AO21x2_ASAP7_75t_L g255 ( .A1(n_256), .A2(n_258), .B(n_266), .Y(n_255) );
AO21x2_ASAP7_75t_L g319 ( .A1(n_256), .A2(n_258), .B(n_266), .Y(n_319) );
INVx2_ASAP7_75t_SL g256 ( .A(n_257), .Y(n_256) );
OA21x2_ASAP7_75t_L g273 ( .A1(n_257), .A2(n_274), .B(n_278), .Y(n_273) );
NAND2xp5_ASAP7_75t_SL g258 ( .A(n_259), .B(n_265), .Y(n_258) );
INVx1_ASAP7_75t_L g261 ( .A(n_262), .Y(n_261) );
INVxp33_ASAP7_75t_L g267 ( .A(n_268), .Y(n_267) );
NAND2x1p5_ASAP7_75t_L g268 ( .A(n_269), .B(n_271), .Y(n_268) );
INVx3_ASAP7_75t_L g334 ( .A(n_269), .Y(n_334) );
INVx3_ASAP7_75t_L g269 ( .A(n_270), .Y(n_269) );
HB1xp67_ASAP7_75t_L g332 ( .A(n_270), .Y(n_332) );
AND2x2_ASAP7_75t_L g501 ( .A(n_270), .B(n_502), .Y(n_501) );
INVx3_ASAP7_75t_L g389 ( .A(n_271), .Y(n_389) );
NAND2xp5_ASAP7_75t_L g521 ( .A(n_271), .B(n_426), .Y(n_521) );
BUFx3_ASAP7_75t_L g271 ( .A(n_272), .Y(n_271) );
AND2x2_ASAP7_75t_L g336 ( .A(n_272), .B(n_337), .Y(n_336) );
INVx1_ASAP7_75t_L g272 ( .A(n_273), .Y(n_272) );
AND2x4_ASAP7_75t_L g317 ( .A(n_273), .B(n_318), .Y(n_317) );
INVx2_ASAP7_75t_L g360 ( .A(n_273), .Y(n_360) );
INVxp67_ASAP7_75t_L g374 ( .A(n_273), .Y(n_374) );
INVx1_ASAP7_75t_L g434 ( .A(n_273), .Y(n_434) );
HB1xp67_ASAP7_75t_L g502 ( .A(n_273), .Y(n_502) );
INVx1_ASAP7_75t_L g486 ( .A(n_279), .Y(n_486) );
NOR2x1_ASAP7_75t_L g279 ( .A(n_280), .B(n_282), .Y(n_279) );
NOR2x1_ASAP7_75t_L g406 ( .A(n_280), .B(n_407), .Y(n_406) );
INVx1_ASAP7_75t_L g280 ( .A(n_281), .Y(n_280) );
AND2x2_ASAP7_75t_L g440 ( .A(n_281), .B(n_312), .Y(n_440) );
OR2x2_ASAP7_75t_L g476 ( .A(n_282), .B(n_477), .Y(n_476) );
INVx2_ASAP7_75t_L g282 ( .A(n_283), .Y(n_282) );
AND2x2_ASAP7_75t_L g458 ( .A(n_283), .B(n_436), .Y(n_458) );
AND2x2_ASAP7_75t_L g510 ( .A(n_283), .B(n_345), .Y(n_510) );
AND2x2_ASAP7_75t_L g283 ( .A(n_284), .B(n_295), .Y(n_283) );
AND2x4_ASAP7_75t_L g312 ( .A(n_284), .B(n_313), .Y(n_312) );
INVx1_ASAP7_75t_L g324 ( .A(n_284), .Y(n_324) );
INVx2_ASAP7_75t_L g341 ( .A(n_284), .Y(n_341) );
HB1xp67_ASAP7_75t_L g519 ( .A(n_284), .Y(n_519) );
AND2x2_ASAP7_75t_L g284 ( .A(n_285), .B(n_290), .Y(n_284) );
NOR3xp33_ASAP7_75t_L g286 ( .A(n_287), .B(n_288), .C(n_289), .Y(n_286) );
INVxp67_ASAP7_75t_L g544 ( .A(n_288), .Y(n_544) );
INVx3_ASAP7_75t_L g313 ( .A(n_295), .Y(n_313) );
INVx2_ASAP7_75t_L g407 ( .A(n_295), .Y(n_407) );
AND2x4_ASAP7_75t_L g295 ( .A(n_296), .B(n_297), .Y(n_295) );
OAI21xp5_ASAP7_75t_L g297 ( .A1(n_298), .A2(n_301), .B(n_308), .Y(n_297) );
OAI22xp5_ASAP7_75t_L g301 ( .A1(n_302), .A2(n_303), .B1(n_305), .B2(n_306), .Y(n_301) );
INVxp67_ASAP7_75t_L g303 ( .A(n_304), .Y(n_303) );
INVxp67_ASAP7_75t_L g306 ( .A(n_307), .Y(n_306) );
NAND2xp5_ASAP7_75t_L g309 ( .A(n_310), .B(n_314), .Y(n_309) );
INVx2_ASAP7_75t_L g310 ( .A(n_311), .Y(n_310) );
NOR2xp33_ASAP7_75t_L g404 ( .A(n_311), .B(n_387), .Y(n_404) );
NOR2x1_ASAP7_75t_L g446 ( .A(n_311), .B(n_325), .Y(n_446) );
INVx4_ASAP7_75t_L g311 ( .A(n_312), .Y(n_311) );
NAND2xp5_ASAP7_75t_L g524 ( .A(n_312), .B(n_387), .Y(n_524) );
AND2x2_ASAP7_75t_L g340 ( .A(n_313), .B(n_341), .Y(n_340) );
INVx1_ASAP7_75t_L g354 ( .A(n_313), .Y(n_354) );
AOI22xp5_ASAP7_75t_SL g402 ( .A1(n_314), .A2(n_403), .B1(n_404), .B2(n_405), .Y(n_402) );
AND2x2_ASAP7_75t_L g314 ( .A(n_315), .B(n_317), .Y(n_314) );
NAND2x1p5_ASAP7_75t_L g399 ( .A(n_315), .B(n_373), .Y(n_399) );
INVx2_ASAP7_75t_SL g315 ( .A(n_316), .Y(n_315) );
OR2x2_ASAP7_75t_L g460 ( .A(n_316), .B(n_348), .Y(n_460) );
AND2x2_ASAP7_75t_L g330 ( .A(n_317), .B(n_331), .Y(n_330) );
AND2x4_ASAP7_75t_L g366 ( .A(n_317), .B(n_367), .Y(n_366) );
AND2x2_ASAP7_75t_L g462 ( .A(n_317), .B(n_452), .Y(n_462) );
INVx2_ASAP7_75t_L g318 ( .A(n_319), .Y(n_318) );
AND2x4_ASAP7_75t_L g384 ( .A(n_319), .B(n_385), .Y(n_384) );
INVx1_ASAP7_75t_L g410 ( .A(n_319), .Y(n_410) );
AND2x2_ASAP7_75t_L g500 ( .A(n_319), .B(n_337), .Y(n_500) );
OAI221xp5_ASAP7_75t_L g320 ( .A1(n_321), .A2(n_329), .B1(n_333), .B2(n_338), .C(n_343), .Y(n_320) );
INVx1_ASAP7_75t_L g321 ( .A(n_322), .Y(n_321) );
AND2x2_ASAP7_75t_L g322 ( .A(n_323), .B(n_326), .Y(n_322) );
INVx1_ASAP7_75t_L g401 ( .A(n_323), .Y(n_401) );
NAND2xp5_ASAP7_75t_L g428 ( .A(n_323), .B(n_429), .Y(n_428) );
NAND2xp5_ASAP7_75t_L g516 ( .A(n_323), .B(n_397), .Y(n_516) );
AND2x4_ASAP7_75t_L g323 ( .A(n_324), .B(n_325), .Y(n_323) );
NOR2xp67_ASAP7_75t_SL g369 ( .A(n_325), .B(n_370), .Y(n_369) );
HB1xp67_ASAP7_75t_L g382 ( .A(n_325), .Y(n_382) );
OR2x2_ASAP7_75t_L g466 ( .A(n_325), .B(n_467), .Y(n_466) );
AND2x4_ASAP7_75t_SL g518 ( .A(n_325), .B(n_519), .Y(n_518) );
HB1xp67_ASAP7_75t_L g326 ( .A(n_327), .Y(n_326) );
INVx3_ASAP7_75t_L g387 ( .A(n_327), .Y(n_387) );
INVx2_ASAP7_75t_L g327 ( .A(n_328), .Y(n_327) );
HB1xp67_ASAP7_75t_L g477 ( .A(n_328), .Y(n_477) );
INVx1_ASAP7_75t_L g329 ( .A(n_330), .Y(n_329) );
AOI221x1_ASAP7_75t_L g417 ( .A1(n_330), .A2(n_418), .B1(n_420), .B2(n_423), .C(n_427), .Y(n_417) );
AND2x2_ASAP7_75t_L g403 ( .A(n_331), .B(n_359), .Y(n_403) );
INVx1_ASAP7_75t_L g331 ( .A(n_332), .Y(n_331) );
OR2x2_ASAP7_75t_L g333 ( .A(n_334), .B(n_335), .Y(n_333) );
AND2x2_ASAP7_75t_L g346 ( .A(n_334), .B(n_347), .Y(n_346) );
NAND2xp5_ASAP7_75t_L g473 ( .A(n_334), .B(n_336), .Y(n_473) );
INVx2_ASAP7_75t_L g335 ( .A(n_336), .Y(n_335) );
INVx2_ASAP7_75t_L g338 ( .A(n_339), .Y(n_338) );
AND2x2_ASAP7_75t_L g339 ( .A(n_340), .B(n_342), .Y(n_339) );
AND2x2_ASAP7_75t_SL g344 ( .A(n_340), .B(n_345), .Y(n_344) );
NAND2xp5_ASAP7_75t_L g370 ( .A(n_340), .B(n_353), .Y(n_370) );
INVx2_ASAP7_75t_L g377 ( .A(n_340), .Y(n_377) );
INVx1_ASAP7_75t_L g422 ( .A(n_341), .Y(n_422) );
BUFx2_ASAP7_75t_L g511 ( .A(n_342), .Y(n_511) );
NAND2xp33_ASAP7_75t_SL g343 ( .A(n_344), .B(n_346), .Y(n_343) );
OR2x6_ASAP7_75t_L g376 ( .A(n_345), .B(n_377), .Y(n_376) );
AND2x2_ASAP7_75t_L g457 ( .A(n_345), .B(n_397), .Y(n_457) );
INVx2_ASAP7_75t_L g347 ( .A(n_348), .Y(n_347) );
NAND2xp5_ASAP7_75t_L g349 ( .A(n_350), .B(n_368), .Y(n_349) );
AOI22xp5_ASAP7_75t_L g350 ( .A1(n_351), .A2(n_357), .B1(n_361), .B2(n_366), .Y(n_350) );
NOR2xp33_ASAP7_75t_L g351 ( .A(n_352), .B(n_355), .Y(n_351) );
AND2x2_ASAP7_75t_SL g414 ( .A(n_352), .B(n_356), .Y(n_414) );
AND2x4_ASAP7_75t_L g420 ( .A(n_352), .B(n_421), .Y(n_420) );
AND2x4_ASAP7_75t_SL g352 ( .A(n_353), .B(n_354), .Y(n_352) );
HB1xp67_ASAP7_75t_L g445 ( .A(n_353), .Y(n_445) );
INVx2_ASAP7_75t_L g355 ( .A(n_356), .Y(n_355) );
NOR2xp33_ASAP7_75t_L g395 ( .A(n_356), .B(n_396), .Y(n_395) );
NAND2xp5_ASAP7_75t_L g419 ( .A(n_356), .B(n_387), .Y(n_419) );
HB1xp67_ASAP7_75t_L g503 ( .A(n_356), .Y(n_503) );
AND2x2_ASAP7_75t_L g357 ( .A(n_358), .B(n_359), .Y(n_357) );
AND2x2_ASAP7_75t_L g450 ( .A(n_358), .B(n_451), .Y(n_450) );
INVx3_ASAP7_75t_L g411 ( .A(n_359), .Y(n_411) );
NAND2x1_ASAP7_75t_SL g455 ( .A(n_359), .B(n_410), .Y(n_455) );
AND2x2_ASAP7_75t_L g489 ( .A(n_359), .B(n_384), .Y(n_489) );
AND2x2_ASAP7_75t_L g361 ( .A(n_362), .B(n_363), .Y(n_361) );
INVx1_ASAP7_75t_L g363 ( .A(n_364), .Y(n_363) );
INVx1_ASAP7_75t_L g364 ( .A(n_365), .Y(n_364) );
AOI22xp5_ASAP7_75t_L g368 ( .A1(n_369), .A2(n_371), .B1(n_375), .B2(n_378), .Y(n_368) );
BUFx2_ASAP7_75t_L g484 ( .A(n_370), .Y(n_484) );
AOI22xp33_ASAP7_75t_L g522 ( .A1(n_371), .A2(n_440), .B1(n_514), .B2(n_523), .Y(n_522) );
AND2x2_ASAP7_75t_L g371 ( .A(n_372), .B(n_373), .Y(n_371) );
NAND2x1p5_ASAP7_75t_L g425 ( .A(n_372), .B(n_426), .Y(n_425) );
AND2x2_ASAP7_75t_L g392 ( .A(n_373), .B(n_393), .Y(n_392) );
INVx2_ASAP7_75t_L g375 ( .A(n_376), .Y(n_375) );
NAND3xp33_ASAP7_75t_L g508 ( .A(n_377), .B(n_509), .C(n_511), .Y(n_508) );
INVx1_ASAP7_75t_L g412 ( .A(n_378), .Y(n_412) );
AOI211x1_ASAP7_75t_L g379 ( .A1(n_380), .A2(n_388), .B(n_390), .C(n_408), .Y(n_379) );
INVx1_ASAP7_75t_L g380 ( .A(n_381), .Y(n_380) );
NAND2xp5_ASAP7_75t_L g381 ( .A(n_382), .B(n_383), .Y(n_381) );
NAND2xp5_ASAP7_75t_SL g439 ( .A(n_383), .B(n_440), .Y(n_439) );
AND2x2_ASAP7_75t_L g383 ( .A(n_384), .B(n_386), .Y(n_383) );
AND2x2_ASAP7_75t_L g470 ( .A(n_384), .B(n_471), .Y(n_470) );
NAND2xp5_ASAP7_75t_L g482 ( .A(n_384), .B(n_451), .Y(n_482) );
AND2x2_ASAP7_75t_L g514 ( .A(n_384), .B(n_452), .Y(n_514) );
INVx1_ASAP7_75t_L g386 ( .A(n_387), .Y(n_386) );
INVx1_ASAP7_75t_L g495 ( .A(n_387), .Y(n_495) );
INVx1_ASAP7_75t_L g388 ( .A(n_389), .Y(n_388) );
OR2x2_ASAP7_75t_L g424 ( .A(n_389), .B(n_425), .Y(n_424) );
NAND2xp5_ASAP7_75t_L g390 ( .A(n_391), .B(n_402), .Y(n_390) );
AOI22xp5_ASAP7_75t_SL g391 ( .A1(n_392), .A2(n_395), .B1(n_398), .B2(n_400), .Y(n_391) );
BUFx2_ASAP7_75t_L g393 ( .A(n_394), .Y(n_393) );
AND2x2_ASAP7_75t_L g432 ( .A(n_394), .B(n_433), .Y(n_432) );
INVx1_ASAP7_75t_SL g447 ( .A(n_394), .Y(n_447) );
INVx1_ASAP7_75t_L g396 ( .A(n_397), .Y(n_396) );
AND2x2_ASAP7_75t_SL g517 ( .A(n_397), .B(n_518), .Y(n_517) );
INVx3_ASAP7_75t_L g398 ( .A(n_399), .Y(n_398) );
INVxp67_ASAP7_75t_L g400 ( .A(n_401), .Y(n_400) );
HB1xp67_ASAP7_75t_L g405 ( .A(n_406), .Y(n_405) );
AND2x2_ASAP7_75t_L g453 ( .A(n_406), .B(n_436), .Y(n_453) );
AOI21xp5_ASAP7_75t_L g408 ( .A1(n_409), .A2(n_412), .B(n_413), .Y(n_408) );
OR2x2_ASAP7_75t_L g409 ( .A(n_410), .B(n_411), .Y(n_409) );
NAND2xp5_ASAP7_75t_L g507 ( .A(n_410), .B(n_432), .Y(n_507) );
OR2x2_ASAP7_75t_L g485 ( .A(n_411), .B(n_430), .Y(n_485) );
INVx1_ASAP7_75t_SL g413 ( .A(n_414), .Y(n_413) );
INVx1_ASAP7_75t_L g415 ( .A(n_416), .Y(n_415) );
NAND3x1_ASAP7_75t_L g416 ( .A(n_417), .B(n_437), .C(n_461), .Y(n_416) );
INVx1_ASAP7_75t_L g418 ( .A(n_419), .Y(n_418) );
AOI22xp5_ASAP7_75t_L g449 ( .A1(n_420), .A2(n_450), .B1(n_453), .B2(n_454), .Y(n_449) );
NAND2xp5_ASAP7_75t_SL g435 ( .A(n_421), .B(n_436), .Y(n_435) );
INVx2_ASAP7_75t_SL g494 ( .A(n_421), .Y(n_494) );
NAND2xp5_ASAP7_75t_L g498 ( .A(n_421), .B(n_495), .Y(n_498) );
INVx2_ASAP7_75t_L g421 ( .A(n_422), .Y(n_421) );
INVx1_ASAP7_75t_L g423 ( .A(n_424), .Y(n_423) );
OAI222xp33_ASAP7_75t_L g481 ( .A1(n_425), .A2(n_482), .B1(n_483), .B2(n_484), .C1(n_485), .C2(n_486), .Y(n_481) );
OAI22xp5_ASAP7_75t_L g427 ( .A1(n_428), .A2(n_430), .B1(n_431), .B2(n_435), .Y(n_427) );
INVx1_ASAP7_75t_SL g467 ( .A(n_429), .Y(n_467) );
INVx1_ASAP7_75t_L g431 ( .A(n_432), .Y(n_431) );
AND2x2_ASAP7_75t_L g504 ( .A(n_433), .B(n_500), .Y(n_504) );
NOR2x1_ASAP7_75t_L g437 ( .A(n_438), .B(n_448), .Y(n_437) );
AOI21xp5_ASAP7_75t_SL g438 ( .A1(n_439), .A2(n_441), .B(n_447), .Y(n_438) );
NAND2xp5_ASAP7_75t_L g441 ( .A(n_442), .B(n_443), .Y(n_441) );
INVx1_ASAP7_75t_L g443 ( .A(n_444), .Y(n_443) );
NAND2xp5_ASAP7_75t_L g444 ( .A(n_445), .B(n_446), .Y(n_444) );
NAND2xp5_ASAP7_75t_L g448 ( .A(n_449), .B(n_456), .Y(n_448) );
INVx1_ASAP7_75t_L g451 ( .A(n_452), .Y(n_451) );
INVx2_ASAP7_75t_SL g454 ( .A(n_455), .Y(n_454) );
NAND2xp5_ASAP7_75t_L g468 ( .A(n_455), .B(n_469), .Y(n_468) );
OAI21xp5_ASAP7_75t_SL g456 ( .A1(n_457), .A2(n_458), .B(n_459), .Y(n_456) );
INVx1_ASAP7_75t_L g483 ( .A(n_458), .Y(n_483) );
INVx1_ASAP7_75t_SL g459 ( .A(n_460), .Y(n_459) );
AOI221xp5_ASAP7_75t_L g461 ( .A1(n_462), .A2(n_463), .B1(n_465), .B2(n_468), .C(n_472), .Y(n_461) );
INVx1_ASAP7_75t_L g463 ( .A(n_464), .Y(n_463) );
INVxp67_ASAP7_75t_L g465 ( .A(n_466), .Y(n_465) );
INVx2_ASAP7_75t_L g469 ( .A(n_470), .Y(n_469) );
AOI21xp5_ASAP7_75t_L g472 ( .A1(n_473), .A2(n_474), .B(n_476), .Y(n_472) );
INVx1_ASAP7_75t_L g474 ( .A(n_475), .Y(n_474) );
INVxp67_ASAP7_75t_SL g478 ( .A(n_479), .Y(n_478) );
NAND3x1_ASAP7_75t_L g479 ( .A(n_480), .B(n_505), .C(n_512), .Y(n_479) );
NOR2x1_ASAP7_75t_L g480 ( .A(n_481), .B(n_487), .Y(n_480) );
NAND2xp5_ASAP7_75t_L g487 ( .A(n_488), .B(n_496), .Y(n_487) );
NAND2xp5_ASAP7_75t_SL g488 ( .A(n_489), .B(n_490), .Y(n_488) );
NAND2xp5_ASAP7_75t_L g490 ( .A(n_491), .B(n_493), .Y(n_490) );
NAND2xp5_ASAP7_75t_L g497 ( .A(n_491), .B(n_498), .Y(n_497) );
INVx1_ASAP7_75t_L g491 ( .A(n_492), .Y(n_491) );
NAND2xp5_ASAP7_75t_L g493 ( .A(n_494), .B(n_495), .Y(n_493) );
AOI22xp5_ASAP7_75t_L g496 ( .A1(n_497), .A2(n_499), .B1(n_503), .B2(n_504), .Y(n_496) );
AND2x4_ASAP7_75t_L g499 ( .A(n_500), .B(n_501), .Y(n_499) );
NAND2xp5_ASAP7_75t_SL g505 ( .A(n_506), .B(n_508), .Y(n_505) );
INVx1_ASAP7_75t_L g506 ( .A(n_507), .Y(n_506) );
INVx1_ASAP7_75t_L g509 ( .A(n_510), .Y(n_509) );
AND2x2_ASAP7_75t_L g512 ( .A(n_513), .B(n_522), .Y(n_512) );
AOI22xp5_ASAP7_75t_SL g513 ( .A1(n_514), .A2(n_515), .B1(n_517), .B2(n_520), .Y(n_513) );
INVx1_ASAP7_75t_L g515 ( .A(n_516), .Y(n_515) );
INVxp67_ASAP7_75t_L g520 ( .A(n_521), .Y(n_520) );
INVx1_ASAP7_75t_L g523 ( .A(n_524), .Y(n_523) );
CKINVDCx20_ASAP7_75t_R g525 ( .A(n_526), .Y(n_525) );
OAI222xp33_ASAP7_75t_L g527 ( .A1(n_528), .A2(n_530), .B1(n_536), .B2(n_538), .C1(n_541), .C2(n_545), .Y(n_527) );
CKINVDCx20_ASAP7_75t_R g530 ( .A(n_531), .Y(n_530) );
CKINVDCx20_ASAP7_75t_R g531 ( .A(n_532), .Y(n_531) );
OR2x2_ASAP7_75t_L g532 ( .A(n_533), .B(n_534), .Y(n_532) );
CKINVDCx20_ASAP7_75t_R g538 ( .A(n_539), .Y(n_538) );
INVx2_ASAP7_75t_L g539 ( .A(n_540), .Y(n_539) );
CKINVDCx20_ASAP7_75t_R g541 ( .A(n_542), .Y(n_541) );
endmodule