module fake_ibex_98_n_2003 (n_151, n_85, n_395, n_84, n_64, n_171, n_103, n_389, n_204, n_274, n_387, n_130, n_177, n_76, n_273, n_309, n_330, n_9, n_328, n_293, n_341, n_372, n_124, n_37, n_256, n_418, n_193, n_446, n_108, n_350, n_165, n_86, n_70, n_255, n_175, n_398, n_59, n_28, n_125, n_304, n_191, n_5, n_62, n_71, n_153, n_194, n_249, n_334, n_312, n_239, n_94, n_134, n_432, n_371, n_403, n_423, n_357, n_88, n_412, n_142, n_226, n_336, n_258, n_40, n_90, n_17, n_74, n_176, n_58, n_43, n_216, n_33, n_421, n_166, n_163, n_114, n_236, n_34, n_376, n_377, n_15, n_24, n_189, n_280, n_317, n_340, n_375, n_105, n_187, n_1, n_154, n_182, n_196, n_326, n_327, n_89, n_50, n_144, n_170, n_270, n_346, n_383, n_113, n_117, n_417, n_265, n_158, n_259, n_276, n_339, n_210, n_348, n_220, n_91, n_287, n_54, n_243, n_19, n_228, n_147, n_251, n_384, n_373, n_244, n_73, n_343, n_310, n_426, n_323, n_143, n_106, n_386, n_8, n_224, n_183, n_67, n_333, n_110, n_306, n_400, n_47, n_169, n_10, n_21, n_242, n_278, n_316, n_16, n_404, n_60, n_7, n_109, n_127, n_121, n_48, n_325, n_57, n_301, n_434, n_296, n_120, n_168, n_155, n_315, n_441, n_13, n_122, n_116, n_370, n_431, n_0, n_289, n_12, n_150, n_286, n_321, n_133, n_51, n_215, n_279, n_49, n_374, n_235, n_22, n_136, n_261, n_30, n_367, n_221, n_437, n_355, n_407, n_102, n_52, n_448, n_99, n_269, n_156, n_126, n_356, n_25, n_104, n_45, n_420, n_141, n_222, n_186, n_349, n_295, n_331, n_230, n_96, n_185, n_388, n_352, n_290, n_174, n_427, n_157, n_219, n_246, n_31, n_442, n_146, n_207, n_438, n_167, n_128, n_253, n_208, n_234, n_3, n_152, n_300, n_145, n_65, n_358, n_205, n_139, n_429, n_275, n_98, n_129, n_267, n_245, n_229, n_209, n_347, n_445, n_335, n_413, n_82, n_263, n_27, n_353, n_359, n_299, n_87, n_262, n_433, n_75, n_439, n_137, n_338, n_173, n_363, n_402, n_180, n_369, n_201, n_14, n_351, n_368, n_257, n_77, n_44, n_401, n_66, n_305, n_307, n_192, n_140, n_416, n_365, n_4, n_6, n_100, n_179, n_354, n_206, n_392, n_329, n_447, n_26, n_188, n_200, n_444, n_199, n_410, n_308, n_411, n_135, n_283, n_366, n_397, n_111, n_36, n_18, n_322, n_53, n_227, n_115, n_11, n_248, n_92, n_101, n_190, n_138, n_409, n_214, n_238, n_332, n_211, n_218, n_314, n_132, n_277, n_337, n_225, n_360, n_272, n_23, n_223, n_381, n_382, n_95, n_405, n_415, n_285, n_288, n_247, n_320, n_379, n_55, n_291, n_318, n_63, n_161, n_237, n_29, n_203, n_268, n_440, n_148, n_2, n_342, n_233, n_385, n_414, n_430, n_118, n_378, n_422, n_164, n_38, n_198, n_264, n_217, n_324, n_391, n_78, n_20, n_69, n_390, n_39, n_178, n_303, n_362, n_93, n_162, n_240, n_282, n_61, n_266, n_42, n_294, n_112, n_46, n_284, n_80, n_172, n_250, n_313, n_345, n_408, n_119, n_361, n_419, n_72, n_319, n_195, n_212, n_311, n_406, n_97, n_197, n_181, n_131, n_123, n_260, n_302, n_443, n_344, n_393, n_436, n_428, n_297, n_435, n_41, n_252, n_396, n_83, n_32, n_107, n_149, n_399, n_254, n_213, n_424, n_271, n_241, n_68, n_292, n_394, n_79, n_81, n_35, n_364, n_159, n_202, n_231, n_298, n_160, n_184, n_56, n_232, n_380, n_281, n_425, n_2003);

input n_151;
input n_85;
input n_395;
input n_84;
input n_64;
input n_171;
input n_103;
input n_389;
input n_204;
input n_274;
input n_387;
input n_130;
input n_177;
input n_76;
input n_273;
input n_309;
input n_330;
input n_9;
input n_328;
input n_293;
input n_341;
input n_372;
input n_124;
input n_37;
input n_256;
input n_418;
input n_193;
input n_446;
input n_108;
input n_350;
input n_165;
input n_86;
input n_70;
input n_255;
input n_175;
input n_398;
input n_59;
input n_28;
input n_125;
input n_304;
input n_191;
input n_5;
input n_62;
input n_71;
input n_153;
input n_194;
input n_249;
input n_334;
input n_312;
input n_239;
input n_94;
input n_134;
input n_432;
input n_371;
input n_403;
input n_423;
input n_357;
input n_88;
input n_412;
input n_142;
input n_226;
input n_336;
input n_258;
input n_40;
input n_90;
input n_17;
input n_74;
input n_176;
input n_58;
input n_43;
input n_216;
input n_33;
input n_421;
input n_166;
input n_163;
input n_114;
input n_236;
input n_34;
input n_376;
input n_377;
input n_15;
input n_24;
input n_189;
input n_280;
input n_317;
input n_340;
input n_375;
input n_105;
input n_187;
input n_1;
input n_154;
input n_182;
input n_196;
input n_326;
input n_327;
input n_89;
input n_50;
input n_144;
input n_170;
input n_270;
input n_346;
input n_383;
input n_113;
input n_117;
input n_417;
input n_265;
input n_158;
input n_259;
input n_276;
input n_339;
input n_210;
input n_348;
input n_220;
input n_91;
input n_287;
input n_54;
input n_243;
input n_19;
input n_228;
input n_147;
input n_251;
input n_384;
input n_373;
input n_244;
input n_73;
input n_343;
input n_310;
input n_426;
input n_323;
input n_143;
input n_106;
input n_386;
input n_8;
input n_224;
input n_183;
input n_67;
input n_333;
input n_110;
input n_306;
input n_400;
input n_47;
input n_169;
input n_10;
input n_21;
input n_242;
input n_278;
input n_316;
input n_16;
input n_404;
input n_60;
input n_7;
input n_109;
input n_127;
input n_121;
input n_48;
input n_325;
input n_57;
input n_301;
input n_434;
input n_296;
input n_120;
input n_168;
input n_155;
input n_315;
input n_441;
input n_13;
input n_122;
input n_116;
input n_370;
input n_431;
input n_0;
input n_289;
input n_12;
input n_150;
input n_286;
input n_321;
input n_133;
input n_51;
input n_215;
input n_279;
input n_49;
input n_374;
input n_235;
input n_22;
input n_136;
input n_261;
input n_30;
input n_367;
input n_221;
input n_437;
input n_355;
input n_407;
input n_102;
input n_52;
input n_448;
input n_99;
input n_269;
input n_156;
input n_126;
input n_356;
input n_25;
input n_104;
input n_45;
input n_420;
input n_141;
input n_222;
input n_186;
input n_349;
input n_295;
input n_331;
input n_230;
input n_96;
input n_185;
input n_388;
input n_352;
input n_290;
input n_174;
input n_427;
input n_157;
input n_219;
input n_246;
input n_31;
input n_442;
input n_146;
input n_207;
input n_438;
input n_167;
input n_128;
input n_253;
input n_208;
input n_234;
input n_3;
input n_152;
input n_300;
input n_145;
input n_65;
input n_358;
input n_205;
input n_139;
input n_429;
input n_275;
input n_98;
input n_129;
input n_267;
input n_245;
input n_229;
input n_209;
input n_347;
input n_445;
input n_335;
input n_413;
input n_82;
input n_263;
input n_27;
input n_353;
input n_359;
input n_299;
input n_87;
input n_262;
input n_433;
input n_75;
input n_439;
input n_137;
input n_338;
input n_173;
input n_363;
input n_402;
input n_180;
input n_369;
input n_201;
input n_14;
input n_351;
input n_368;
input n_257;
input n_77;
input n_44;
input n_401;
input n_66;
input n_305;
input n_307;
input n_192;
input n_140;
input n_416;
input n_365;
input n_4;
input n_6;
input n_100;
input n_179;
input n_354;
input n_206;
input n_392;
input n_329;
input n_447;
input n_26;
input n_188;
input n_200;
input n_444;
input n_199;
input n_410;
input n_308;
input n_411;
input n_135;
input n_283;
input n_366;
input n_397;
input n_111;
input n_36;
input n_18;
input n_322;
input n_53;
input n_227;
input n_115;
input n_11;
input n_248;
input n_92;
input n_101;
input n_190;
input n_138;
input n_409;
input n_214;
input n_238;
input n_332;
input n_211;
input n_218;
input n_314;
input n_132;
input n_277;
input n_337;
input n_225;
input n_360;
input n_272;
input n_23;
input n_223;
input n_381;
input n_382;
input n_95;
input n_405;
input n_415;
input n_285;
input n_288;
input n_247;
input n_320;
input n_379;
input n_55;
input n_291;
input n_318;
input n_63;
input n_161;
input n_237;
input n_29;
input n_203;
input n_268;
input n_440;
input n_148;
input n_2;
input n_342;
input n_233;
input n_385;
input n_414;
input n_430;
input n_118;
input n_378;
input n_422;
input n_164;
input n_38;
input n_198;
input n_264;
input n_217;
input n_324;
input n_391;
input n_78;
input n_20;
input n_69;
input n_390;
input n_39;
input n_178;
input n_303;
input n_362;
input n_93;
input n_162;
input n_240;
input n_282;
input n_61;
input n_266;
input n_42;
input n_294;
input n_112;
input n_46;
input n_284;
input n_80;
input n_172;
input n_250;
input n_313;
input n_345;
input n_408;
input n_119;
input n_361;
input n_419;
input n_72;
input n_319;
input n_195;
input n_212;
input n_311;
input n_406;
input n_97;
input n_197;
input n_181;
input n_131;
input n_123;
input n_260;
input n_302;
input n_443;
input n_344;
input n_393;
input n_436;
input n_428;
input n_297;
input n_435;
input n_41;
input n_252;
input n_396;
input n_83;
input n_32;
input n_107;
input n_149;
input n_399;
input n_254;
input n_213;
input n_424;
input n_271;
input n_241;
input n_68;
input n_292;
input n_394;
input n_79;
input n_81;
input n_35;
input n_364;
input n_159;
input n_202;
input n_231;
input n_298;
input n_160;
input n_184;
input n_56;
input n_232;
input n_380;
input n_281;
input n_425;

output n_2003;

wire n_1084;
wire n_1474;
wire n_1295;
wire n_507;
wire n_1983;
wire n_992;
wire n_1582;
wire n_766;
wire n_1110;
wire n_1382;
wire n_1998;
wire n_1596;
wire n_926;
wire n_1079;
wire n_1100;
wire n_845;
wire n_1930;
wire n_452;
wire n_1234;
wire n_1594;
wire n_1944;
wire n_1802;
wire n_773;
wire n_1469;
wire n_821;
wire n_873;
wire n_1227;
wire n_962;
wire n_1080;
wire n_862;
wire n_909;
wire n_957;
wire n_1652;
wire n_969;
wire n_678;
wire n_1859;
wire n_1954;
wire n_1883;
wire n_1125;
wire n_733;
wire n_622;
wire n_1226;
wire n_1034;
wire n_1765;
wire n_872;
wire n_1873;
wire n_1619;
wire n_457;
wire n_1666;
wire n_494;
wire n_930;
wire n_1044;
wire n_1492;
wire n_1134;
wire n_1478;
wire n_1684;
wire n_1796;
wire n_1614;
wire n_1722;
wire n_911;
wire n_652;
wire n_781;
wire n_475;
wire n_802;
wire n_1233;
wire n_1045;
wire n_1856;
wire n_500;
wire n_963;
wire n_1782;
wire n_531;
wire n_1308;
wire n_556;
wire n_1138;
wire n_498;
wire n_708;
wire n_1096;
wire n_1391;
wire n_667;
wire n_884;
wire n_850;
wire n_1971;
wire n_879;
wire n_1957;
wire n_723;
wire n_1144;
wire n_1392;
wire n_1268;
wire n_739;
wire n_853;
wire n_948;
wire n_504;
wire n_1752;
wire n_1829;
wire n_1338;
wire n_1730;
wire n_875;
wire n_1307;
wire n_1327;
wire n_481;
wire n_876;
wire n_497;
wire n_711;
wire n_1840;
wire n_671;
wire n_989;
wire n_1908;
wire n_1668;
wire n_1641;
wire n_829;
wire n_825;
wire n_1480;
wire n_1463;
wire n_1823;
wire n_1681;
wire n_939;
wire n_1636;
wire n_1687;
wire n_655;
wire n_1766;
wire n_550;
wire n_1922;
wire n_557;
wire n_641;
wire n_1937;
wire n_893;
wire n_527;
wire n_1654;
wire n_496;
wire n_1258;
wire n_1344;
wire n_1929;
wire n_1749;
wire n_1680;
wire n_835;
wire n_1981;
wire n_1195;
wire n_824;
wire n_1945;
wire n_694;
wire n_523;
wire n_787;
wire n_614;
wire n_1130;
wire n_1228;
wire n_1081;
wire n_538;
wire n_1155;
wire n_1292;
wire n_459;
wire n_1576;
wire n_1664;
wire n_518;
wire n_852;
wire n_1427;
wire n_1133;
wire n_1926;
wire n_904;
wire n_1970;
wire n_1778;
wire n_646;
wire n_466;
wire n_1030;
wire n_1698;
wire n_1094;
wire n_1496;
wire n_1910;
wire n_715;
wire n_530;
wire n_1663;
wire n_1214;
wire n_1274;
wire n_1606;
wire n_769;
wire n_1595;
wire n_1509;
wire n_1618;
wire n_1648;
wire n_1886;
wire n_857;
wire n_765;
wire n_1070;
wire n_1841;
wire n_777;
wire n_1955;
wire n_917;
wire n_968;
wire n_1253;
wire n_1306;
wire n_1484;
wire n_1493;
wire n_1313;
wire n_558;
wire n_666;
wire n_1638;
wire n_1071;
wire n_1449;
wire n_1723;
wire n_1960;
wire n_793;
wire n_937;
wire n_1645;
wire n_973;
wire n_1038;
wire n_618;
wire n_1943;
wire n_1863;
wire n_1269;
wire n_662;
wire n_979;
wire n_1309;
wire n_1999;
wire n_1316;
wire n_1562;
wire n_1215;
wire n_629;
wire n_1445;
wire n_573;
wire n_1716;
wire n_1466;
wire n_1412;
wire n_1672;
wire n_1007;
wire n_643;
wire n_1276;
wire n_1637;
wire n_841;
wire n_772;
wire n_810;
wire n_1401;
wire n_1817;
wire n_1588;
wire n_1301;
wire n_869;
wire n_1620;
wire n_1561;
wire n_718;
wire n_554;
wire n_553;
wire n_1078;
wire n_1219;
wire n_713;
wire n_1865;
wire n_1252;
wire n_1170;
wire n_1927;
wire n_605;
wire n_539;
wire n_630;
wire n_1869;
wire n_567;
wire n_1853;
wire n_745;
wire n_1753;
wire n_562;
wire n_564;
wire n_1322;
wire n_1305;
wire n_795;
wire n_592;
wire n_1248;
wire n_762;
wire n_1388;
wire n_800;
wire n_706;
wire n_784;
wire n_684;
wire n_1653;
wire n_1375;
wire n_1356;
wire n_894;
wire n_1118;
wire n_692;
wire n_1881;
wire n_1969;
wire n_709;
wire n_1296;
wire n_499;
wire n_971;
wire n_702;
wire n_1326;
wire n_451;
wire n_1350;
wire n_906;
wire n_1093;
wire n_1764;
wire n_978;
wire n_579;
wire n_899;
wire n_1799;
wire n_1019;
wire n_902;
wire n_1689;
wire n_1250;
wire n_1190;
wire n_1304;
wire n_744;
wire n_563;
wire n_1506;
wire n_881;
wire n_1702;
wire n_734;
wire n_1558;
wire n_1650;
wire n_1520;
wire n_1073;
wire n_1453;
wire n_1108;
wire n_1794;
wire n_1423;
wire n_1239;
wire n_1370;
wire n_1209;
wire n_1708;
wire n_551;
wire n_1616;
wire n_729;
wire n_1569;
wire n_1434;
wire n_603;
wire n_1649;
wire n_1936;
wire n_1717;
wire n_1609;
wire n_1613;
wire n_820;
wire n_805;
wire n_1988;
wire n_670;
wire n_1132;
wire n_892;
wire n_1467;
wire n_1803;
wire n_544;
wire n_1787;
wire n_1281;
wire n_1447;
wire n_695;
wire n_1549;
wire n_639;
wire n_1867;
wire n_1531;
wire n_1332;
wire n_482;
wire n_1424;
wire n_1742;
wire n_1818;
wire n_870;
wire n_1709;
wire n_1610;
wire n_1298;
wire n_1844;
wire n_1387;
wire n_609;
wire n_1040;
wire n_476;
wire n_1159;
wire n_1368;
wire n_1154;
wire n_455;
wire n_1701;
wire n_1243;
wire n_1121;
wire n_693;
wire n_606;
wire n_737;
wire n_1571;
wire n_1980;
wire n_462;
wire n_1407;
wire n_1235;
wire n_1821;
wire n_1003;
wire n_889;
wire n_816;
wire n_1058;
wire n_1835;
wire n_1862;
wire n_1543;
wire n_823;
wire n_1504;
wire n_1519;
wire n_1425;
wire n_1781;
wire n_1441;
wire n_1924;
wire n_1921;
wire n_657;
wire n_1156;
wire n_1293;
wire n_1360;
wire n_749;
wire n_1555;
wire n_1394;
wire n_1347;
wire n_819;
wire n_822;
wire n_1042;
wire n_1888;
wire n_743;
wire n_754;
wire n_1786;
wire n_1319;
wire n_1553;
wire n_1041;
wire n_1964;
wire n_1090;
wire n_1196;
wire n_1182;
wire n_1271;
wire n_1731;
wire n_1905;
wire n_1031;
wire n_981;
wire n_1591;
wire n_583;
wire n_1671;
wire n_1795;
wire n_1409;
wire n_1015;
wire n_663;
wire n_1377;
wire n_1583;
wire n_1521;
wire n_1152;
wire n_974;
wire n_1036;
wire n_1831;
wire n_864;
wire n_608;
wire n_1987;
wire n_959;
wire n_1106;
wire n_1312;
wire n_1129;
wire n_1244;
wire n_449;
wire n_1733;
wire n_1634;
wire n_1932;
wire n_1452;
wire n_1552;
wire n_1318;
wire n_1508;
wire n_738;
wire n_1217;
wire n_1715;
wire n_1189;
wire n_761;
wire n_748;
wire n_1713;
wire n_901;
wire n_1577;
wire n_1255;
wire n_1700;
wire n_1218;
wire n_1181;
wire n_1140;
wire n_1985;
wire n_1772;
wire n_1056;
wire n_1283;
wire n_1446;
wire n_1487;
wire n_840;
wire n_1203;
wire n_1421;
wire n_561;
wire n_471;
wire n_846;
wire n_1793;
wire n_1237;
wire n_859;
wire n_965;
wire n_1109;
wire n_1633;
wire n_1711;
wire n_1051;
wire n_1008;
wire n_458;
wire n_1498;
wire n_1053;
wire n_1656;
wire n_1207;
wire n_1735;
wire n_1076;
wire n_1032;
wire n_936;
wire n_469;
wire n_1884;
wire n_1825;
wire n_1589;
wire n_1210;
wire n_591;
wire n_1933;
wire n_1996;
wire n_1510;
wire n_1201;
wire n_1842;
wire n_1246;
wire n_1677;
wire n_732;
wire n_1236;
wire n_832;
wire n_1792;
wire n_1712;
wire n_1984;
wire n_590;
wire n_1568;
wire n_1877;
wire n_1184;
wire n_1477;
wire n_1724;
wire n_1364;
wire n_1540;
wire n_1676;
wire n_1013;
wire n_929;
wire n_637;
wire n_1136;
wire n_1890;
wire n_1075;
wire n_1249;
wire n_1918;
wire n_574;
wire n_515;
wire n_1229;
wire n_1440;
wire n_1490;
wire n_907;
wire n_1179;
wire n_1990;
wire n_1153;
wire n_1751;
wire n_669;
wire n_1737;
wire n_521;
wire n_1117;
wire n_1273;
wire n_1748;
wire n_1083;
wire n_1014;
wire n_724;
wire n_938;
wire n_1178;
wire n_474;
wire n_878;
wire n_594;
wire n_1464;
wire n_1566;
wire n_944;
wire n_1848;
wire n_623;
wire n_585;
wire n_1982;
wire n_1334;
wire n_1963;
wire n_483;
wire n_1695;
wire n_1418;
wire n_1137;
wire n_660;
wire n_524;
wire n_1977;
wire n_1200;
wire n_1120;
wire n_576;
wire n_1602;
wire n_1776;
wire n_1852;
wire n_1522;
wire n_1279;
wire n_931;
wire n_607;
wire n_827;
wire n_1064;
wire n_1408;
wire n_1028;
wire n_1264;
wire n_1935;
wire n_1146;
wire n_488;
wire n_705;
wire n_1548;
wire n_1682;
wire n_1608;
wire n_1009;
wire n_1260;
wire n_589;
wire n_1896;
wire n_472;
wire n_1704;
wire n_847;
wire n_1436;
wire n_1069;
wire n_1485;
wire n_1465;
wire n_1352;
wire n_1171;
wire n_1126;
wire n_1232;
wire n_1979;
wire n_679;
wire n_1345;
wire n_696;
wire n_837;
wire n_1590;
wire n_640;
wire n_954;
wire n_1628;
wire n_725;
wire n_1773;
wire n_596;
wire n_1545;
wire n_456;
wire n_1471;
wire n_1738;
wire n_998;
wire n_1115;
wire n_1395;
wire n_1729;
wire n_801;
wire n_1479;
wire n_1046;
wire n_882;
wire n_942;
wire n_1627;
wire n_1431;
wire n_651;
wire n_721;
wire n_814;
wire n_1864;
wire n_943;
wire n_1086;
wire n_1523;
wire n_1756;
wire n_1470;
wire n_1761;
wire n_1836;
wire n_1593;
wire n_986;
wire n_495;
wire n_1420;
wire n_1750;
wire n_1775;
wire n_1699;
wire n_927;
wire n_1563;
wire n_615;
wire n_803;
wire n_1875;
wire n_1615;
wire n_1087;
wire n_757;
wire n_1400;
wire n_712;
wire n_1599;
wire n_1806;
wire n_1539;
wire n_650;
wire n_1575;
wire n_1448;
wire n_517;
wire n_817;
wire n_555;
wire n_951;
wire n_468;
wire n_1580;
wire n_1574;
wire n_780;
wire n_502;
wire n_1705;
wire n_633;
wire n_1746;
wire n_532;
wire n_726;
wire n_1439;
wire n_863;
wire n_597;
wire n_1832;
wire n_1128;
wire n_1266;
wire n_1300;
wire n_807;
wire n_741;
wire n_1785;
wire n_486;
wire n_1870;
wire n_1405;
wire n_997;
wire n_1428;
wire n_891;
wire n_1528;
wire n_1495;
wire n_717;
wire n_1357;
wire n_1512;
wire n_668;
wire n_871;
wire n_1339;
wire n_1544;
wire n_1426;
wire n_485;
wire n_1315;
wire n_1413;
wire n_811;
wire n_808;
wire n_945;
wire n_460;
wire n_1706;
wire n_1560;
wire n_1592;
wire n_1461;
wire n_461;
wire n_903;
wire n_1967;
wire n_1095;
wire n_1328;
wire n_1265;
wire n_1378;
wire n_1048;
wire n_774;
wire n_1925;
wire n_588;
wire n_1430;
wire n_1251;
wire n_1247;
wire n_528;
wire n_836;
wire n_1475;
wire n_1263;
wire n_1185;
wire n_1683;
wire n_1122;
wire n_890;
wire n_628;
wire n_874;
wire n_1505;
wire n_1163;
wire n_677;
wire n_1514;
wire n_964;
wire n_916;
wire n_503;
wire n_895;
wire n_687;
wire n_1035;
wire n_1535;
wire n_751;
wire n_1127;
wire n_932;
wire n_1972;
wire n_947;
wire n_1004;
wire n_831;
wire n_778;
wire n_1898;
wire n_1254;
wire n_1148;
wire n_540;
wire n_1667;
wire n_1104;
wire n_1845;
wire n_1011;
wire n_1437;
wire n_529;
wire n_626;
wire n_1707;
wire n_1941;
wire n_1679;
wire n_1497;
wire n_2002;
wire n_1578;
wire n_1143;
wire n_1783;
wire n_510;
wire n_972;
wire n_1815;
wire n_601;
wire n_610;
wire n_1917;
wire n_1444;
wire n_920;
wire n_664;
wire n_1067;
wire n_994;
wire n_2000;
wire n_1857;
wire n_1920;
wire n_545;
wire n_887;
wire n_1162;
wire n_1997;
wire n_1894;
wire n_961;
wire n_991;
wire n_634;
wire n_1223;
wire n_1349;
wire n_1331;
wire n_1323;
wire n_578;
wire n_1739;
wire n_1777;
wire n_1353;
wire n_1429;
wire n_1546;
wire n_1432;
wire n_1950;
wire n_1320;
wire n_996;
wire n_915;
wire n_1174;
wire n_1874;
wire n_1834;
wire n_1727;
wire n_1286;
wire n_1657;
wire n_1741;
wire n_542;
wire n_1294;
wire n_1601;
wire n_900;
wire n_1351;
wire n_647;
wire n_1380;
wire n_1367;
wire n_1291;
wire n_1914;
wire n_1458;
wire n_1694;
wire n_1460;
wire n_1830;
wire n_1629;
wire n_1826;
wire n_1855;
wire n_1662;
wire n_1340;
wire n_1626;
wire n_674;
wire n_1660;
wire n_1850;
wire n_1643;
wire n_1670;
wire n_1789;
wire n_552;
wire n_1112;
wire n_1267;
wire n_1384;
wire n_1376;
wire n_1537;
wire n_1858;
wire n_1816;
wire n_1612;
wire n_703;
wire n_1172;
wire n_1099;
wire n_598;
wire n_1422;
wire n_508;
wire n_453;
wire n_1527;
wire n_1055;
wire n_1524;
wire n_673;
wire n_798;
wire n_1754;
wire n_1177;
wire n_1025;
wire n_1991;
wire n_1517;
wire n_690;
wire n_1225;
wire n_1962;
wire n_982;
wire n_1624;
wire n_785;
wire n_1952;
wire n_604;
wire n_1598;
wire n_977;
wire n_1895;
wire n_719;
wire n_1491;
wire n_1860;
wire n_716;
wire n_1810;
wire n_1763;
wire n_923;
wire n_642;
wire n_1607;
wire n_1625;
wire n_933;
wire n_1774;
wire n_1797;
wire n_1037;
wire n_1899;
wire n_464;
wire n_1289;
wire n_838;
wire n_1348;
wire n_1021;
wire n_746;
wire n_1557;
wire n_1188;
wire n_1567;
wire n_742;
wire n_1191;
wire n_1503;
wire n_1052;
wire n_789;
wire n_1942;
wire n_656;
wire n_602;
wire n_842;
wire n_767;
wire n_1617;
wire n_1839;
wire n_1587;
wire n_636;
wire n_1259;
wire n_490;
wire n_595;
wire n_1001;
wire n_570;
wire n_1396;
wire n_1224;
wire n_1923;
wire n_1538;
wire n_487;
wire n_454;
wire n_1017;
wire n_730;
wire n_1456;
wire n_1889;
wire n_625;
wire n_619;
wire n_1124;
wire n_611;
wire n_1690;
wire n_1673;
wire n_922;
wire n_1790;
wire n_851;
wire n_993;
wire n_1725;
wire n_1135;
wire n_2001;
wire n_1820;
wire n_1800;
wire n_541;
wire n_613;
wire n_659;
wire n_1494;
wire n_1550;
wire n_1066;
wire n_648;
wire n_571;
wire n_1169;
wire n_1726;
wire n_1946;
wire n_1938;
wire n_830;
wire n_473;
wire n_1241;
wire n_1072;
wire n_1231;
wire n_1173;
wire n_1208;
wire n_1639;
wire n_1604;
wire n_826;
wire n_1976;
wire n_1337;
wire n_1906;
wire n_1647;
wire n_1901;
wire n_768;
wire n_839;
wire n_1278;
wire n_796;
wire n_797;
wire n_1006;
wire n_1238;
wire n_1415;
wire n_976;
wire n_1710;
wire n_1063;
wire n_1270;
wire n_834;
wire n_1476;
wire n_935;
wire n_1603;
wire n_925;
wire n_1054;
wire n_722;
wire n_1644;
wire n_1406;
wire n_1489;
wire n_1880;
wire n_1993;
wire n_804;
wire n_484;
wire n_1455;
wire n_1642;
wire n_1871;
wire n_480;
wire n_1057;
wire n_1473;
wire n_516;
wire n_1403;
wire n_1149;
wire n_1176;
wire n_1502;
wire n_1605;
wire n_506;
wire n_868;
wire n_1202;
wire n_1065;
wire n_1897;
wire n_1457;
wire n_905;
wire n_975;
wire n_675;
wire n_463;
wire n_624;
wire n_520;
wire n_934;
wire n_775;
wire n_512;
wire n_950;
wire n_685;
wire n_1222;
wire n_1630;
wire n_1879;
wire n_1959;
wire n_1198;
wire n_1311;
wire n_1261;
wire n_776;
wire n_1114;
wire n_818;
wire n_1167;
wire n_1282;
wire n_1321;
wire n_700;
wire n_1779;
wire n_1770;
wire n_1107;
wire n_1846;
wire n_1573;
wire n_525;
wire n_815;
wire n_919;
wire n_535;
wire n_1956;
wire n_681;
wire n_1718;
wire n_1411;
wire n_1139;
wire n_1018;
wire n_858;
wire n_1324;
wire n_1669;
wire n_1501;
wire n_782;
wire n_616;
wire n_1885;
wire n_1740;
wire n_1989;
wire n_1838;
wire n_833;
wire n_1343;
wire n_1801;
wire n_1371;
wire n_1513;
wire n_728;
wire n_1788;
wire n_786;
wire n_505;
wire n_1621;
wire n_1919;
wire n_1342;
wire n_501;
wire n_752;
wire n_958;
wire n_1175;
wire n_1416;
wire n_1659;
wire n_1221;
wire n_1047;
wire n_1878;
wire n_1515;
wire n_1374;
wire n_1435;
wire n_1688;
wire n_792;
wire n_1433;
wire n_1314;
wire n_575;
wire n_1242;
wire n_1119;
wire n_1085;
wire n_1907;
wire n_885;
wire n_1530;
wire n_513;
wire n_877;
wire n_1088;
wire n_896;
wire n_1813;
wire n_1451;
wire n_1005;
wire n_1102;
wire n_631;
wire n_794;
wire n_1288;
wire n_1275;
wire n_985;
wire n_1165;
wire n_897;
wire n_1622;
wire n_697;
wire n_1105;
wire n_1459;
wire n_912;
wire n_1893;
wire n_1570;
wire n_701;
wire n_995;
wire n_1000;
wire n_1931;
wire n_1256;
wire n_587;
wire n_1303;
wire n_1994;
wire n_1771;
wire n_1526;
wire n_764;
wire n_1507;
wire n_1206;
wire n_1809;
wire n_855;
wire n_812;
wire n_1961;
wire n_1050;
wire n_599;
wire n_1769;
wire n_1060;
wire n_1372;
wire n_1847;
wire n_756;
wire n_1565;
wire n_1257;
wire n_1632;
wire n_688;
wire n_1547;
wire n_946;
wire n_1542;
wire n_707;
wire n_1362;
wire n_1586;
wire n_1097;
wire n_1909;
wire n_621;
wire n_956;
wire n_790;
wire n_1541;
wire n_1812;
wire n_1951;
wire n_586;
wire n_1330;
wire n_638;
wire n_1697;
wire n_1872;
wire n_1940;
wire n_593;
wire n_1747;
wire n_1212;
wire n_1887;
wire n_1199;
wire n_1978;
wire n_1767;
wire n_1939;
wire n_1768;
wire n_1443;
wire n_478;
wire n_1585;
wire n_1861;
wire n_1564;
wire n_1995;
wire n_1631;
wire n_1623;
wire n_861;
wire n_1828;
wire n_1389;
wire n_1131;
wire n_547;
wire n_1798;
wire n_727;
wire n_1077;
wire n_1554;
wire n_1584;
wire n_1481;
wire n_1928;
wire n_828;
wire n_1438;
wire n_1973;
wire n_753;
wire n_747;
wire n_645;
wire n_1147;
wire n_1363;
wire n_1691;
wire n_1098;
wire n_584;
wire n_1366;
wire n_1518;
wire n_1187;
wire n_1361;
wire n_1693;
wire n_698;
wire n_1892;
wire n_1061;
wire n_682;
wire n_1373;
wire n_1686;
wire n_1302;
wire n_886;
wire n_1010;
wire n_883;
wire n_755;
wire n_1029;
wire n_470;
wire n_770;
wire n_1572;
wire n_1635;
wire n_941;
wire n_1245;
wire n_1317;
wire n_632;
wire n_1329;
wire n_854;
wire n_1369;
wire n_714;
wire n_1297;
wire n_1912;
wire n_1734;
wire n_1876;
wire n_740;
wire n_549;
wire n_533;
wire n_1811;
wire n_928;
wire n_898;
wire n_1285;
wire n_967;
wire n_736;
wire n_1529;
wire n_1381;
wire n_1824;
wire n_1597;
wire n_1103;
wire n_1161;
wire n_465;
wire n_1486;
wire n_1068;
wire n_617;
wire n_1833;
wire n_914;
wire n_1986;
wire n_526;
wire n_1024;
wire n_1141;
wire n_1949;
wire n_1197;
wire n_1168;
wire n_865;
wire n_569;
wire n_600;
wire n_1556;
wire n_1192;
wire n_1646;
wire n_1290;
wire n_1759;
wire n_987;
wire n_750;
wire n_1299;
wire n_665;
wire n_1101;
wire n_1720;
wire n_880;
wire n_654;
wire n_1911;
wire n_731;
wire n_1336;
wire n_1166;
wire n_758;
wire n_720;
wire n_710;
wire n_1390;
wire n_1023;
wire n_568;
wire n_1358;
wire n_813;
wire n_1211;
wire n_1397;
wire n_1284;
wire n_1359;
wire n_1116;
wire n_1758;
wire n_791;
wire n_1532;
wire n_1419;
wire n_543;
wire n_580;
wire n_1784;
wire n_1685;
wire n_1992;
wire n_1082;
wire n_1213;
wire n_980;
wire n_1193;
wire n_849;
wire n_1488;
wire n_1074;
wire n_759;
wire n_1379;
wire n_1721;
wire n_1827;
wire n_953;
wire n_1180;
wire n_1462;
wire n_536;
wire n_1866;
wire n_1220;
wire n_467;
wire n_1398;
wire n_1262;
wire n_1904;
wire n_1692;
wire n_1012;
wire n_1805;
wire n_689;
wire n_960;
wire n_1022;
wire n_1760;
wire n_676;
wire n_1240;
wire n_1183;
wire n_1204;
wire n_1151;
wire n_1814;
wire n_771;
wire n_999;
wire n_514;
wire n_1092;
wire n_1808;
wire n_560;
wire n_1658;
wire n_1386;
wire n_910;
wire n_635;
wire n_844;
wire n_1728;
wire n_1020;
wire n_783;
wire n_1142;
wire n_1385;
wire n_1062;
wire n_1230;
wire n_1027;
wire n_1516;
wire n_1499;
wire n_1500;
wire n_1868;
wire n_966;
wire n_949;
wire n_704;
wire n_924;
wire n_1600;
wire n_477;
wire n_1661;
wire n_1965;
wire n_1757;
wire n_699;
wire n_918;
wire n_1913;
wire n_672;
wire n_1039;
wire n_1043;
wire n_1402;
wire n_735;
wire n_1450;
wire n_566;
wire n_581;
wire n_1365;
wire n_1472;
wire n_1089;
wire n_1536;
wire n_1049;
wire n_1719;
wire n_1974;
wire n_548;
wire n_1158;
wire n_763;
wire n_1882;
wire n_1915;
wire n_940;
wire n_1762;
wire n_1404;
wire n_546;
wire n_788;
wire n_1736;
wire n_1160;
wire n_1442;
wire n_658;
wire n_1948;
wire n_1216;
wire n_1891;
wire n_1026;
wire n_1454;
wire n_1033;
wire n_627;
wire n_990;
wire n_1383;
wire n_1968;
wire n_888;
wire n_1325;
wire n_582;
wire n_1483;
wire n_1703;
wire n_653;
wire n_1205;
wire n_1822;
wire n_843;
wire n_1953;
wire n_1059;
wire n_799;
wire n_691;
wire n_1804;
wire n_1581;
wire n_522;
wire n_479;
wire n_534;
wire n_1837;
wire n_511;
wire n_1744;
wire n_1975;
wire n_1414;
wire n_1002;
wire n_1851;
wire n_1755;
wire n_1111;
wire n_1819;
wire n_1341;
wire n_1807;
wire n_1310;
wire n_1745;
wire n_1714;
wire n_612;
wire n_1958;
wire n_1611;
wire n_955;
wire n_1333;
wire n_1916;
wire n_952;
wire n_1675;
wire n_1947;
wire n_1640;
wire n_1551;
wire n_1145;
wire n_1533;
wire n_1511;
wire n_1791;
wire n_537;
wire n_1113;
wire n_1651;
wire n_1966;
wire n_1468;
wire n_913;
wire n_509;
wire n_1164;
wire n_1732;
wire n_1354;
wire n_1277;
wire n_1696;
wire n_1016;
wire n_680;
wire n_1355;
wire n_809;
wire n_856;
wire n_779;
wire n_1559;
wire n_1579;
wire n_1280;
wire n_493;
wire n_1335;
wire n_1934;
wire n_1900;
wire n_519;
wire n_1843;
wire n_1665;
wire n_1091;
wire n_1678;
wire n_1780;
wire n_1287;
wire n_1482;
wire n_860;
wire n_1525;
wire n_661;
wire n_848;
wire n_1902;
wire n_683;
wire n_1150;
wire n_1194;
wire n_620;
wire n_1399;
wire n_450;
wire n_1903;
wire n_1674;
wire n_1849;
wire n_686;
wire n_572;
wire n_867;
wire n_983;
wire n_1417;
wire n_644;
wire n_577;
wire n_970;
wire n_491;
wire n_921;
wire n_489;
wire n_1534;
wire n_908;
wire n_1346;
wire n_565;
wire n_1123;
wire n_1272;
wire n_1393;
wire n_984;
wire n_1655;
wire n_1410;
wire n_988;
wire n_760;
wire n_1157;
wire n_806;
wire n_1186;
wire n_1743;
wire n_492;
wire n_649;
wire n_1854;
wire n_866;
wire n_559;

BUFx3_ASAP7_75t_L g449 ( 
.A(n_345),
.Y(n_449)
);

BUFx10_ASAP7_75t_L g450 ( 
.A(n_434),
.Y(n_450)
);

CKINVDCx5p33_ASAP7_75t_R g451 ( 
.A(n_217),
.Y(n_451)
);

INVx1_ASAP7_75t_L g452 ( 
.A(n_31),
.Y(n_452)
);

INVx1_ASAP7_75t_L g453 ( 
.A(n_124),
.Y(n_453)
);

CKINVDCx5p33_ASAP7_75t_R g454 ( 
.A(n_12),
.Y(n_454)
);

INVx2_ASAP7_75t_L g455 ( 
.A(n_388),
.Y(n_455)
);

CKINVDCx5p33_ASAP7_75t_R g456 ( 
.A(n_275),
.Y(n_456)
);

CKINVDCx5p33_ASAP7_75t_R g457 ( 
.A(n_398),
.Y(n_457)
);

INVx1_ASAP7_75t_L g458 ( 
.A(n_359),
.Y(n_458)
);

CKINVDCx5p33_ASAP7_75t_R g459 ( 
.A(n_346),
.Y(n_459)
);

INVx2_ASAP7_75t_L g460 ( 
.A(n_328),
.Y(n_460)
);

BUFx6f_ASAP7_75t_L g461 ( 
.A(n_370),
.Y(n_461)
);

CKINVDCx5p33_ASAP7_75t_R g462 ( 
.A(n_277),
.Y(n_462)
);

CKINVDCx20_ASAP7_75t_R g463 ( 
.A(n_421),
.Y(n_463)
);

CKINVDCx5p33_ASAP7_75t_R g464 ( 
.A(n_439),
.Y(n_464)
);

CKINVDCx5p33_ASAP7_75t_R g465 ( 
.A(n_1),
.Y(n_465)
);

CKINVDCx5p33_ASAP7_75t_R g466 ( 
.A(n_406),
.Y(n_466)
);

CKINVDCx5p33_ASAP7_75t_R g467 ( 
.A(n_435),
.Y(n_467)
);

CKINVDCx5p33_ASAP7_75t_R g468 ( 
.A(n_376),
.Y(n_468)
);

CKINVDCx5p33_ASAP7_75t_R g469 ( 
.A(n_48),
.Y(n_469)
);

CKINVDCx5p33_ASAP7_75t_R g470 ( 
.A(n_223),
.Y(n_470)
);

CKINVDCx5p33_ASAP7_75t_R g471 ( 
.A(n_109),
.Y(n_471)
);

CKINVDCx5p33_ASAP7_75t_R g472 ( 
.A(n_318),
.Y(n_472)
);

BUFx2_ASAP7_75t_SL g473 ( 
.A(n_412),
.Y(n_473)
);

INVx1_ASAP7_75t_L g474 ( 
.A(n_441),
.Y(n_474)
);

CKINVDCx5p33_ASAP7_75t_R g475 ( 
.A(n_19),
.Y(n_475)
);

CKINVDCx5p33_ASAP7_75t_R g476 ( 
.A(n_331),
.Y(n_476)
);

CKINVDCx5p33_ASAP7_75t_R g477 ( 
.A(n_126),
.Y(n_477)
);

INVx1_ASAP7_75t_L g478 ( 
.A(n_14),
.Y(n_478)
);

CKINVDCx5p33_ASAP7_75t_R g479 ( 
.A(n_12),
.Y(n_479)
);

CKINVDCx5p33_ASAP7_75t_R g480 ( 
.A(n_105),
.Y(n_480)
);

INVx1_ASAP7_75t_L g481 ( 
.A(n_299),
.Y(n_481)
);

CKINVDCx5p33_ASAP7_75t_R g482 ( 
.A(n_79),
.Y(n_482)
);

CKINVDCx5p33_ASAP7_75t_R g483 ( 
.A(n_240),
.Y(n_483)
);

INVx1_ASAP7_75t_L g484 ( 
.A(n_140),
.Y(n_484)
);

CKINVDCx20_ASAP7_75t_R g485 ( 
.A(n_43),
.Y(n_485)
);

CKINVDCx5p33_ASAP7_75t_R g486 ( 
.A(n_177),
.Y(n_486)
);

CKINVDCx5p33_ASAP7_75t_R g487 ( 
.A(n_55),
.Y(n_487)
);

INVx3_ASAP7_75t_L g488 ( 
.A(n_46),
.Y(n_488)
);

INVx1_ASAP7_75t_L g489 ( 
.A(n_160),
.Y(n_489)
);

INVx2_ASAP7_75t_SL g490 ( 
.A(n_62),
.Y(n_490)
);

INVx1_ASAP7_75t_SL g491 ( 
.A(n_99),
.Y(n_491)
);

CKINVDCx5p33_ASAP7_75t_R g492 ( 
.A(n_40),
.Y(n_492)
);

INVx2_ASAP7_75t_L g493 ( 
.A(n_237),
.Y(n_493)
);

CKINVDCx5p33_ASAP7_75t_R g494 ( 
.A(n_407),
.Y(n_494)
);

CKINVDCx5p33_ASAP7_75t_R g495 ( 
.A(n_404),
.Y(n_495)
);

INVx2_ASAP7_75t_L g496 ( 
.A(n_372),
.Y(n_496)
);

CKINVDCx5p33_ASAP7_75t_R g497 ( 
.A(n_416),
.Y(n_497)
);

CKINVDCx5p33_ASAP7_75t_R g498 ( 
.A(n_70),
.Y(n_498)
);

INVx2_ASAP7_75t_L g499 ( 
.A(n_105),
.Y(n_499)
);

INVx1_ASAP7_75t_L g500 ( 
.A(n_429),
.Y(n_500)
);

INVx1_ASAP7_75t_L g501 ( 
.A(n_227),
.Y(n_501)
);

CKINVDCx5p33_ASAP7_75t_R g502 ( 
.A(n_231),
.Y(n_502)
);

CKINVDCx5p33_ASAP7_75t_R g503 ( 
.A(n_24),
.Y(n_503)
);

CKINVDCx5p33_ASAP7_75t_R g504 ( 
.A(n_375),
.Y(n_504)
);

CKINVDCx5p33_ASAP7_75t_R g505 ( 
.A(n_149),
.Y(n_505)
);

INVx2_ASAP7_75t_SL g506 ( 
.A(n_443),
.Y(n_506)
);

CKINVDCx5p33_ASAP7_75t_R g507 ( 
.A(n_432),
.Y(n_507)
);

CKINVDCx5p33_ASAP7_75t_R g508 ( 
.A(n_168),
.Y(n_508)
);

INVx2_ASAP7_75t_SL g509 ( 
.A(n_233),
.Y(n_509)
);

CKINVDCx5p33_ASAP7_75t_R g510 ( 
.A(n_293),
.Y(n_510)
);

CKINVDCx5p33_ASAP7_75t_R g511 ( 
.A(n_107),
.Y(n_511)
);

INVx1_ASAP7_75t_L g512 ( 
.A(n_273),
.Y(n_512)
);

CKINVDCx5p33_ASAP7_75t_R g513 ( 
.A(n_280),
.Y(n_513)
);

BUFx10_ASAP7_75t_L g514 ( 
.A(n_396),
.Y(n_514)
);

BUFx6f_ASAP7_75t_L g515 ( 
.A(n_52),
.Y(n_515)
);

INVx1_ASAP7_75t_SL g516 ( 
.A(n_63),
.Y(n_516)
);

CKINVDCx5p33_ASAP7_75t_R g517 ( 
.A(n_73),
.Y(n_517)
);

INVx1_ASAP7_75t_L g518 ( 
.A(n_199),
.Y(n_518)
);

BUFx10_ASAP7_75t_L g519 ( 
.A(n_313),
.Y(n_519)
);

BUFx3_ASAP7_75t_L g520 ( 
.A(n_236),
.Y(n_520)
);

CKINVDCx5p33_ASAP7_75t_R g521 ( 
.A(n_377),
.Y(n_521)
);

CKINVDCx5p33_ASAP7_75t_R g522 ( 
.A(n_369),
.Y(n_522)
);

BUFx2_ASAP7_75t_L g523 ( 
.A(n_334),
.Y(n_523)
);

CKINVDCx20_ASAP7_75t_R g524 ( 
.A(n_191),
.Y(n_524)
);

CKINVDCx5p33_ASAP7_75t_R g525 ( 
.A(n_213),
.Y(n_525)
);

BUFx3_ASAP7_75t_L g526 ( 
.A(n_363),
.Y(n_526)
);

BUFx6f_ASAP7_75t_L g527 ( 
.A(n_145),
.Y(n_527)
);

CKINVDCx5p33_ASAP7_75t_R g528 ( 
.A(n_425),
.Y(n_528)
);

INVx1_ASAP7_75t_L g529 ( 
.A(n_408),
.Y(n_529)
);

INVx1_ASAP7_75t_L g530 ( 
.A(n_129),
.Y(n_530)
);

CKINVDCx5p33_ASAP7_75t_R g531 ( 
.A(n_29),
.Y(n_531)
);

CKINVDCx5p33_ASAP7_75t_R g532 ( 
.A(n_117),
.Y(n_532)
);

INVx1_ASAP7_75t_L g533 ( 
.A(n_218),
.Y(n_533)
);

INVx2_ASAP7_75t_L g534 ( 
.A(n_226),
.Y(n_534)
);

HB1xp67_ASAP7_75t_L g535 ( 
.A(n_186),
.Y(n_535)
);

BUFx3_ASAP7_75t_L g536 ( 
.A(n_57),
.Y(n_536)
);

INVx1_ASAP7_75t_L g537 ( 
.A(n_103),
.Y(n_537)
);

CKINVDCx20_ASAP7_75t_R g538 ( 
.A(n_360),
.Y(n_538)
);

CKINVDCx20_ASAP7_75t_R g539 ( 
.A(n_63),
.Y(n_539)
);

CKINVDCx5p33_ASAP7_75t_R g540 ( 
.A(n_9),
.Y(n_540)
);

CKINVDCx5p33_ASAP7_75t_R g541 ( 
.A(n_23),
.Y(n_541)
);

INVx1_ASAP7_75t_L g542 ( 
.A(n_302),
.Y(n_542)
);

INVx1_ASAP7_75t_L g543 ( 
.A(n_176),
.Y(n_543)
);

INVx2_ASAP7_75t_SL g544 ( 
.A(n_437),
.Y(n_544)
);

CKINVDCx5p33_ASAP7_75t_R g545 ( 
.A(n_120),
.Y(n_545)
);

CKINVDCx5p33_ASAP7_75t_R g546 ( 
.A(n_224),
.Y(n_546)
);

INVx2_ASAP7_75t_SL g547 ( 
.A(n_389),
.Y(n_547)
);

CKINVDCx5p33_ASAP7_75t_R g548 ( 
.A(n_113),
.Y(n_548)
);

CKINVDCx5p33_ASAP7_75t_R g549 ( 
.A(n_1),
.Y(n_549)
);

CKINVDCx5p33_ASAP7_75t_R g550 ( 
.A(n_246),
.Y(n_550)
);

CKINVDCx5p33_ASAP7_75t_R g551 ( 
.A(n_14),
.Y(n_551)
);

CKINVDCx16_ASAP7_75t_R g552 ( 
.A(n_316),
.Y(n_552)
);

INVx1_ASAP7_75t_L g553 ( 
.A(n_303),
.Y(n_553)
);

CKINVDCx5p33_ASAP7_75t_R g554 ( 
.A(n_68),
.Y(n_554)
);

INVxp67_ASAP7_75t_L g555 ( 
.A(n_138),
.Y(n_555)
);

BUFx3_ASAP7_75t_L g556 ( 
.A(n_326),
.Y(n_556)
);

INVx1_ASAP7_75t_L g557 ( 
.A(n_400),
.Y(n_557)
);

CKINVDCx5p33_ASAP7_75t_R g558 ( 
.A(n_243),
.Y(n_558)
);

INVx2_ASAP7_75t_SL g559 ( 
.A(n_265),
.Y(n_559)
);

INVx1_ASAP7_75t_L g560 ( 
.A(n_201),
.Y(n_560)
);

INVx2_ASAP7_75t_SL g561 ( 
.A(n_353),
.Y(n_561)
);

CKINVDCx5p33_ASAP7_75t_R g562 ( 
.A(n_16),
.Y(n_562)
);

CKINVDCx14_ASAP7_75t_R g563 ( 
.A(n_254),
.Y(n_563)
);

INVx1_ASAP7_75t_L g564 ( 
.A(n_419),
.Y(n_564)
);

BUFx10_ASAP7_75t_L g565 ( 
.A(n_357),
.Y(n_565)
);

CKINVDCx5p33_ASAP7_75t_R g566 ( 
.A(n_445),
.Y(n_566)
);

CKINVDCx5p33_ASAP7_75t_R g567 ( 
.A(n_430),
.Y(n_567)
);

CKINVDCx5p33_ASAP7_75t_R g568 ( 
.A(n_127),
.Y(n_568)
);

CKINVDCx5p33_ASAP7_75t_R g569 ( 
.A(n_269),
.Y(n_569)
);

INVx1_ASAP7_75t_L g570 ( 
.A(n_200),
.Y(n_570)
);

INVx1_ASAP7_75t_L g571 ( 
.A(n_208),
.Y(n_571)
);

CKINVDCx5p33_ASAP7_75t_R g572 ( 
.A(n_319),
.Y(n_572)
);

CKINVDCx5p33_ASAP7_75t_R g573 ( 
.A(n_151),
.Y(n_573)
);

CKINVDCx5p33_ASAP7_75t_R g574 ( 
.A(n_381),
.Y(n_574)
);

INVx2_ASAP7_75t_L g575 ( 
.A(n_431),
.Y(n_575)
);

INVx2_ASAP7_75t_L g576 ( 
.A(n_390),
.Y(n_576)
);

INVx2_ASAP7_75t_SL g577 ( 
.A(n_433),
.Y(n_577)
);

CKINVDCx5p33_ASAP7_75t_R g578 ( 
.A(n_436),
.Y(n_578)
);

INVx1_ASAP7_75t_L g579 ( 
.A(n_317),
.Y(n_579)
);

CKINVDCx5p33_ASAP7_75t_R g580 ( 
.A(n_26),
.Y(n_580)
);

INVx1_ASAP7_75t_L g581 ( 
.A(n_397),
.Y(n_581)
);

BUFx6f_ASAP7_75t_L g582 ( 
.A(n_194),
.Y(n_582)
);

INVx1_ASAP7_75t_SL g583 ( 
.A(n_148),
.Y(n_583)
);

CKINVDCx20_ASAP7_75t_R g584 ( 
.A(n_8),
.Y(n_584)
);

CKINVDCx5p33_ASAP7_75t_R g585 ( 
.A(n_215),
.Y(n_585)
);

BUFx6f_ASAP7_75t_L g586 ( 
.A(n_73),
.Y(n_586)
);

BUFx6f_ASAP7_75t_L g587 ( 
.A(n_378),
.Y(n_587)
);

CKINVDCx5p33_ASAP7_75t_R g588 ( 
.A(n_150),
.Y(n_588)
);

INVx1_ASAP7_75t_L g589 ( 
.A(n_36),
.Y(n_589)
);

INVx1_ASAP7_75t_L g590 ( 
.A(n_66),
.Y(n_590)
);

CKINVDCx5p33_ASAP7_75t_R g591 ( 
.A(n_25),
.Y(n_591)
);

INVx1_ASAP7_75t_L g592 ( 
.A(n_411),
.Y(n_592)
);

CKINVDCx5p33_ASAP7_75t_R g593 ( 
.A(n_181),
.Y(n_593)
);

CKINVDCx5p33_ASAP7_75t_R g594 ( 
.A(n_415),
.Y(n_594)
);

CKINVDCx5p33_ASAP7_75t_R g595 ( 
.A(n_391),
.Y(n_595)
);

INVx1_ASAP7_75t_L g596 ( 
.A(n_402),
.Y(n_596)
);

CKINVDCx5p33_ASAP7_75t_R g597 ( 
.A(n_179),
.Y(n_597)
);

CKINVDCx5p33_ASAP7_75t_R g598 ( 
.A(n_324),
.Y(n_598)
);

INVx1_ASAP7_75t_L g599 ( 
.A(n_395),
.Y(n_599)
);

CKINVDCx5p33_ASAP7_75t_R g600 ( 
.A(n_290),
.Y(n_600)
);

CKINVDCx5p33_ASAP7_75t_R g601 ( 
.A(n_85),
.Y(n_601)
);

CKINVDCx5p33_ASAP7_75t_R g602 ( 
.A(n_77),
.Y(n_602)
);

CKINVDCx20_ASAP7_75t_R g603 ( 
.A(n_348),
.Y(n_603)
);

CKINVDCx5p33_ASAP7_75t_R g604 ( 
.A(n_95),
.Y(n_604)
);

INVx1_ASAP7_75t_L g605 ( 
.A(n_337),
.Y(n_605)
);

CKINVDCx5p33_ASAP7_75t_R g606 ( 
.A(n_38),
.Y(n_606)
);

INVx1_ASAP7_75t_L g607 ( 
.A(n_7),
.Y(n_607)
);

INVx1_ASAP7_75t_L g608 ( 
.A(n_329),
.Y(n_608)
);

INVx1_ASAP7_75t_L g609 ( 
.A(n_4),
.Y(n_609)
);

BUFx6f_ASAP7_75t_L g610 ( 
.A(n_420),
.Y(n_610)
);

CKINVDCx5p33_ASAP7_75t_R g611 ( 
.A(n_250),
.Y(n_611)
);

INVx2_ASAP7_75t_L g612 ( 
.A(n_320),
.Y(n_612)
);

INVx1_ASAP7_75t_L g613 ( 
.A(n_392),
.Y(n_613)
);

BUFx6f_ASAP7_75t_L g614 ( 
.A(n_245),
.Y(n_614)
);

INVx1_ASAP7_75t_L g615 ( 
.A(n_394),
.Y(n_615)
);

BUFx3_ASAP7_75t_L g616 ( 
.A(n_136),
.Y(n_616)
);

CKINVDCx5p33_ASAP7_75t_R g617 ( 
.A(n_60),
.Y(n_617)
);

CKINVDCx5p33_ASAP7_75t_R g618 ( 
.A(n_285),
.Y(n_618)
);

CKINVDCx5p33_ASAP7_75t_R g619 ( 
.A(n_386),
.Y(n_619)
);

BUFx2_ASAP7_75t_L g620 ( 
.A(n_118),
.Y(n_620)
);

CKINVDCx5p33_ASAP7_75t_R g621 ( 
.A(n_110),
.Y(n_621)
);

CKINVDCx5p33_ASAP7_75t_R g622 ( 
.A(n_159),
.Y(n_622)
);

CKINVDCx5p33_ASAP7_75t_R g623 ( 
.A(n_242),
.Y(n_623)
);

CKINVDCx5p33_ASAP7_75t_R g624 ( 
.A(n_75),
.Y(n_624)
);

CKINVDCx5p33_ASAP7_75t_R g625 ( 
.A(n_384),
.Y(n_625)
);

BUFx6f_ASAP7_75t_L g626 ( 
.A(n_428),
.Y(n_626)
);

CKINVDCx5p33_ASAP7_75t_R g627 ( 
.A(n_383),
.Y(n_627)
);

CKINVDCx5p33_ASAP7_75t_R g628 ( 
.A(n_427),
.Y(n_628)
);

CKINVDCx5p33_ASAP7_75t_R g629 ( 
.A(n_64),
.Y(n_629)
);

CKINVDCx5p33_ASAP7_75t_R g630 ( 
.A(n_296),
.Y(n_630)
);

INVx1_ASAP7_75t_L g631 ( 
.A(n_409),
.Y(n_631)
);

INVx1_ASAP7_75t_L g632 ( 
.A(n_368),
.Y(n_632)
);

INVx1_ASAP7_75t_L g633 ( 
.A(n_382),
.Y(n_633)
);

CKINVDCx5p33_ASAP7_75t_R g634 ( 
.A(n_321),
.Y(n_634)
);

INVx1_ASAP7_75t_L g635 ( 
.A(n_60),
.Y(n_635)
);

CKINVDCx5p33_ASAP7_75t_R g636 ( 
.A(n_210),
.Y(n_636)
);

INVx1_ASAP7_75t_L g637 ( 
.A(n_56),
.Y(n_637)
);

BUFx10_ASAP7_75t_L g638 ( 
.A(n_162),
.Y(n_638)
);

CKINVDCx5p33_ASAP7_75t_R g639 ( 
.A(n_255),
.Y(n_639)
);

CKINVDCx5p33_ASAP7_75t_R g640 ( 
.A(n_291),
.Y(n_640)
);

CKINVDCx5p33_ASAP7_75t_R g641 ( 
.A(n_157),
.Y(n_641)
);

CKINVDCx5p33_ASAP7_75t_R g642 ( 
.A(n_414),
.Y(n_642)
);

CKINVDCx5p33_ASAP7_75t_R g643 ( 
.A(n_34),
.Y(n_643)
);

CKINVDCx5p33_ASAP7_75t_R g644 ( 
.A(n_222),
.Y(n_644)
);

CKINVDCx5p33_ASAP7_75t_R g645 ( 
.A(n_352),
.Y(n_645)
);

BUFx10_ASAP7_75t_L g646 ( 
.A(n_354),
.Y(n_646)
);

INVx2_ASAP7_75t_L g647 ( 
.A(n_410),
.Y(n_647)
);

INVx1_ASAP7_75t_L g648 ( 
.A(n_164),
.Y(n_648)
);

CKINVDCx5p33_ASAP7_75t_R g649 ( 
.A(n_211),
.Y(n_649)
);

CKINVDCx5p33_ASAP7_75t_R g650 ( 
.A(n_424),
.Y(n_650)
);

INVx2_ASAP7_75t_SL g651 ( 
.A(n_64),
.Y(n_651)
);

CKINVDCx5p33_ASAP7_75t_R g652 ( 
.A(n_0),
.Y(n_652)
);

CKINVDCx5p33_ASAP7_75t_R g653 ( 
.A(n_216),
.Y(n_653)
);

CKINVDCx5p33_ASAP7_75t_R g654 ( 
.A(n_289),
.Y(n_654)
);

CKINVDCx20_ASAP7_75t_R g655 ( 
.A(n_17),
.Y(n_655)
);

INVx1_ASAP7_75t_L g656 ( 
.A(n_342),
.Y(n_656)
);

INVx2_ASAP7_75t_L g657 ( 
.A(n_442),
.Y(n_657)
);

CKINVDCx5p33_ASAP7_75t_R g658 ( 
.A(n_86),
.Y(n_658)
);

INVx1_ASAP7_75t_SL g659 ( 
.A(n_309),
.Y(n_659)
);

CKINVDCx5p33_ASAP7_75t_R g660 ( 
.A(n_438),
.Y(n_660)
);

INVx1_ASAP7_75t_L g661 ( 
.A(n_80),
.Y(n_661)
);

CKINVDCx5p33_ASAP7_75t_R g662 ( 
.A(n_125),
.Y(n_662)
);

INVx1_ASAP7_75t_L g663 ( 
.A(n_221),
.Y(n_663)
);

INVx1_ASAP7_75t_L g664 ( 
.A(n_362),
.Y(n_664)
);

INVx1_ASAP7_75t_SL g665 ( 
.A(n_365),
.Y(n_665)
);

INVx1_ASAP7_75t_L g666 ( 
.A(n_88),
.Y(n_666)
);

CKINVDCx5p33_ASAP7_75t_R g667 ( 
.A(n_121),
.Y(n_667)
);

CKINVDCx5p33_ASAP7_75t_R g668 ( 
.A(n_335),
.Y(n_668)
);

INVx1_ASAP7_75t_L g669 ( 
.A(n_287),
.Y(n_669)
);

INVx1_ASAP7_75t_L g670 ( 
.A(n_2),
.Y(n_670)
);

CKINVDCx5p33_ASAP7_75t_R g671 ( 
.A(n_209),
.Y(n_671)
);

INVx1_ASAP7_75t_L g672 ( 
.A(n_40),
.Y(n_672)
);

CKINVDCx5p33_ASAP7_75t_R g673 ( 
.A(n_413),
.Y(n_673)
);

INVxp67_ASAP7_75t_L g674 ( 
.A(n_248),
.Y(n_674)
);

CKINVDCx5p33_ASAP7_75t_R g675 ( 
.A(n_417),
.Y(n_675)
);

CKINVDCx5p33_ASAP7_75t_R g676 ( 
.A(n_28),
.Y(n_676)
);

CKINVDCx5p33_ASAP7_75t_R g677 ( 
.A(n_238),
.Y(n_677)
);

CKINVDCx5p33_ASAP7_75t_R g678 ( 
.A(n_153),
.Y(n_678)
);

INVx1_ASAP7_75t_L g679 ( 
.A(n_288),
.Y(n_679)
);

CKINVDCx5p33_ASAP7_75t_R g680 ( 
.A(n_350),
.Y(n_680)
);

INVx1_ASAP7_75t_L g681 ( 
.A(n_77),
.Y(n_681)
);

INVx2_ASAP7_75t_SL g682 ( 
.A(n_48),
.Y(n_682)
);

CKINVDCx5p33_ASAP7_75t_R g683 ( 
.A(n_122),
.Y(n_683)
);

INVx2_ASAP7_75t_SL g684 ( 
.A(n_446),
.Y(n_684)
);

INVx1_ASAP7_75t_SL g685 ( 
.A(n_380),
.Y(n_685)
);

CKINVDCx20_ASAP7_75t_R g686 ( 
.A(n_399),
.Y(n_686)
);

INVx1_ASAP7_75t_L g687 ( 
.A(n_9),
.Y(n_687)
);

INVx1_ASAP7_75t_L g688 ( 
.A(n_158),
.Y(n_688)
);

CKINVDCx5p33_ASAP7_75t_R g689 ( 
.A(n_103),
.Y(n_689)
);

BUFx2_ASAP7_75t_SL g690 ( 
.A(n_423),
.Y(n_690)
);

CKINVDCx5p33_ASAP7_75t_R g691 ( 
.A(n_6),
.Y(n_691)
);

CKINVDCx20_ASAP7_75t_R g692 ( 
.A(n_146),
.Y(n_692)
);

CKINVDCx5p33_ASAP7_75t_R g693 ( 
.A(n_418),
.Y(n_693)
);

CKINVDCx5p33_ASAP7_75t_R g694 ( 
.A(n_235),
.Y(n_694)
);

CKINVDCx5p33_ASAP7_75t_R g695 ( 
.A(n_161),
.Y(n_695)
);

CKINVDCx20_ASAP7_75t_R g696 ( 
.A(n_100),
.Y(n_696)
);

CKINVDCx20_ASAP7_75t_R g697 ( 
.A(n_327),
.Y(n_697)
);

CKINVDCx5p33_ASAP7_75t_R g698 ( 
.A(n_403),
.Y(n_698)
);

INVx1_ASAP7_75t_L g699 ( 
.A(n_351),
.Y(n_699)
);

CKINVDCx20_ASAP7_75t_R g700 ( 
.A(n_272),
.Y(n_700)
);

INVx2_ASAP7_75t_L g701 ( 
.A(n_178),
.Y(n_701)
);

INVx1_ASAP7_75t_L g702 ( 
.A(n_204),
.Y(n_702)
);

INVxp67_ASAP7_75t_L g703 ( 
.A(n_447),
.Y(n_703)
);

INVx2_ASAP7_75t_L g704 ( 
.A(n_100),
.Y(n_704)
);

INVx2_ASAP7_75t_SL g705 ( 
.A(n_203),
.Y(n_705)
);

CKINVDCx5p33_ASAP7_75t_R g706 ( 
.A(n_27),
.Y(n_706)
);

INVx1_ASAP7_75t_L g707 ( 
.A(n_42),
.Y(n_707)
);

CKINVDCx5p33_ASAP7_75t_R g708 ( 
.A(n_379),
.Y(n_708)
);

CKINVDCx20_ASAP7_75t_R g709 ( 
.A(n_99),
.Y(n_709)
);

CKINVDCx5p33_ASAP7_75t_R g710 ( 
.A(n_11),
.Y(n_710)
);

INVx1_ASAP7_75t_L g711 ( 
.A(n_278),
.Y(n_711)
);

CKINVDCx16_ASAP7_75t_R g712 ( 
.A(n_267),
.Y(n_712)
);

INVx1_ASAP7_75t_L g713 ( 
.A(n_172),
.Y(n_713)
);

CKINVDCx5p33_ASAP7_75t_R g714 ( 
.A(n_440),
.Y(n_714)
);

CKINVDCx5p33_ASAP7_75t_R g715 ( 
.A(n_156),
.Y(n_715)
);

INVx1_ASAP7_75t_L g716 ( 
.A(n_271),
.Y(n_716)
);

BUFx6f_ASAP7_75t_L g717 ( 
.A(n_385),
.Y(n_717)
);

CKINVDCx5p33_ASAP7_75t_R g718 ( 
.A(n_230),
.Y(n_718)
);

CKINVDCx5p33_ASAP7_75t_R g719 ( 
.A(n_207),
.Y(n_719)
);

CKINVDCx16_ASAP7_75t_R g720 ( 
.A(n_27),
.Y(n_720)
);

BUFx5_ASAP7_75t_L g721 ( 
.A(n_393),
.Y(n_721)
);

INVx1_ASAP7_75t_L g722 ( 
.A(n_422),
.Y(n_722)
);

CKINVDCx5p33_ASAP7_75t_R g723 ( 
.A(n_256),
.Y(n_723)
);

BUFx2_ASAP7_75t_L g724 ( 
.A(n_307),
.Y(n_724)
);

INVx1_ASAP7_75t_L g725 ( 
.A(n_333),
.Y(n_725)
);

INVx1_ASAP7_75t_L g726 ( 
.A(n_387),
.Y(n_726)
);

BUFx10_ASAP7_75t_L g727 ( 
.A(n_88),
.Y(n_727)
);

INVx1_ASAP7_75t_L g728 ( 
.A(n_305),
.Y(n_728)
);

CKINVDCx5p33_ASAP7_75t_R g729 ( 
.A(n_102),
.Y(n_729)
);

CKINVDCx5p33_ASAP7_75t_R g730 ( 
.A(n_22),
.Y(n_730)
);

INVx1_ASAP7_75t_L g731 ( 
.A(n_42),
.Y(n_731)
);

INVx2_ASAP7_75t_L g732 ( 
.A(n_58),
.Y(n_732)
);

INVx1_ASAP7_75t_L g733 ( 
.A(n_84),
.Y(n_733)
);

CKINVDCx5p33_ASAP7_75t_R g734 ( 
.A(n_7),
.Y(n_734)
);

INVx1_ASAP7_75t_L g735 ( 
.A(n_109),
.Y(n_735)
);

INVx1_ASAP7_75t_L g736 ( 
.A(n_374),
.Y(n_736)
);

CKINVDCx5p33_ASAP7_75t_R g737 ( 
.A(n_121),
.Y(n_737)
);

INVx1_ASAP7_75t_L g738 ( 
.A(n_426),
.Y(n_738)
);

CKINVDCx5p33_ASAP7_75t_R g739 ( 
.A(n_405),
.Y(n_739)
);

INVx2_ASAP7_75t_L g740 ( 
.A(n_401),
.Y(n_740)
);

CKINVDCx5p33_ASAP7_75t_R g741 ( 
.A(n_71),
.Y(n_741)
);

CKINVDCx5p33_ASAP7_75t_R g742 ( 
.A(n_189),
.Y(n_742)
);

CKINVDCx5p33_ASAP7_75t_R g743 ( 
.A(n_463),
.Y(n_743)
);

INVx1_ASAP7_75t_L g744 ( 
.A(n_535),
.Y(n_744)
);

INVx2_ASAP7_75t_L g745 ( 
.A(n_721),
.Y(n_745)
);

INVx1_ASAP7_75t_L g746 ( 
.A(n_535),
.Y(n_746)
);

INVx1_ASAP7_75t_L g747 ( 
.A(n_488),
.Y(n_747)
);

INVxp67_ASAP7_75t_SL g748 ( 
.A(n_488),
.Y(n_748)
);

CKINVDCx16_ASAP7_75t_R g749 ( 
.A(n_720),
.Y(n_749)
);

HB1xp67_ASAP7_75t_L g750 ( 
.A(n_620),
.Y(n_750)
);

CKINVDCx20_ASAP7_75t_R g751 ( 
.A(n_485),
.Y(n_751)
);

BUFx3_ASAP7_75t_L g752 ( 
.A(n_449),
.Y(n_752)
);

CKINVDCx5p33_ASAP7_75t_R g753 ( 
.A(n_524),
.Y(n_753)
);

INVx2_ASAP7_75t_L g754 ( 
.A(n_721),
.Y(n_754)
);

INVx1_ASAP7_75t_L g755 ( 
.A(n_523),
.Y(n_755)
);

INVx1_ASAP7_75t_L g756 ( 
.A(n_724),
.Y(n_756)
);

HB1xp67_ASAP7_75t_L g757 ( 
.A(n_536),
.Y(n_757)
);

INVx1_ASAP7_75t_L g758 ( 
.A(n_536),
.Y(n_758)
);

CKINVDCx20_ASAP7_75t_R g759 ( 
.A(n_539),
.Y(n_759)
);

CKINVDCx5p33_ASAP7_75t_R g760 ( 
.A(n_538),
.Y(n_760)
);

INVxp67_ASAP7_75t_SL g761 ( 
.A(n_555),
.Y(n_761)
);

INVx1_ASAP7_75t_L g762 ( 
.A(n_499),
.Y(n_762)
);

INVx1_ASAP7_75t_L g763 ( 
.A(n_704),
.Y(n_763)
);

INVx2_ASAP7_75t_L g764 ( 
.A(n_721),
.Y(n_764)
);

INVx1_ASAP7_75t_L g765 ( 
.A(n_732),
.Y(n_765)
);

CKINVDCx5p33_ASAP7_75t_R g766 ( 
.A(n_603),
.Y(n_766)
);

INVx1_ASAP7_75t_L g767 ( 
.A(n_490),
.Y(n_767)
);

INVx1_ASAP7_75t_L g768 ( 
.A(n_651),
.Y(n_768)
);

INVx1_ASAP7_75t_L g769 ( 
.A(n_682),
.Y(n_769)
);

INVx1_ASAP7_75t_L g770 ( 
.A(n_452),
.Y(n_770)
);

INVx1_ASAP7_75t_L g771 ( 
.A(n_478),
.Y(n_771)
);

INVx1_ASAP7_75t_L g772 ( 
.A(n_537),
.Y(n_772)
);

CKINVDCx16_ASAP7_75t_R g773 ( 
.A(n_552),
.Y(n_773)
);

INVx1_ASAP7_75t_L g774 ( 
.A(n_589),
.Y(n_774)
);

HB1xp67_ASAP7_75t_L g775 ( 
.A(n_454),
.Y(n_775)
);

INVx1_ASAP7_75t_L g776 ( 
.A(n_590),
.Y(n_776)
);

INVx1_ASAP7_75t_L g777 ( 
.A(n_607),
.Y(n_777)
);

CKINVDCx20_ASAP7_75t_R g778 ( 
.A(n_584),
.Y(n_778)
);

CKINVDCx5p33_ASAP7_75t_R g779 ( 
.A(n_686),
.Y(n_779)
);

CKINVDCx20_ASAP7_75t_R g780 ( 
.A(n_655),
.Y(n_780)
);

CKINVDCx20_ASAP7_75t_R g781 ( 
.A(n_696),
.Y(n_781)
);

INVxp33_ASAP7_75t_L g782 ( 
.A(n_609),
.Y(n_782)
);

CKINVDCx5p33_ASAP7_75t_R g783 ( 
.A(n_692),
.Y(n_783)
);

INVx1_ASAP7_75t_L g784 ( 
.A(n_635),
.Y(n_784)
);

INVxp67_ASAP7_75t_SL g785 ( 
.A(n_555),
.Y(n_785)
);

INVx1_ASAP7_75t_L g786 ( 
.A(n_637),
.Y(n_786)
);

INVxp33_ASAP7_75t_SL g787 ( 
.A(n_465),
.Y(n_787)
);

INVx1_ASAP7_75t_L g788 ( 
.A(n_661),
.Y(n_788)
);

INVx1_ASAP7_75t_L g789 ( 
.A(n_666),
.Y(n_789)
);

CKINVDCx20_ASAP7_75t_R g790 ( 
.A(n_709),
.Y(n_790)
);

INVx1_ASAP7_75t_L g791 ( 
.A(n_670),
.Y(n_791)
);

CKINVDCx20_ASAP7_75t_R g792 ( 
.A(n_697),
.Y(n_792)
);

INVx1_ASAP7_75t_L g793 ( 
.A(n_672),
.Y(n_793)
);

INVx1_ASAP7_75t_L g794 ( 
.A(n_681),
.Y(n_794)
);

INVx1_ASAP7_75t_L g795 ( 
.A(n_687),
.Y(n_795)
);

INVx1_ASAP7_75t_L g796 ( 
.A(n_707),
.Y(n_796)
);

INVx1_ASAP7_75t_L g797 ( 
.A(n_731),
.Y(n_797)
);

INVx1_ASAP7_75t_L g798 ( 
.A(n_733),
.Y(n_798)
);

INVxp67_ASAP7_75t_SL g799 ( 
.A(n_674),
.Y(n_799)
);

INVxp67_ASAP7_75t_SL g800 ( 
.A(n_674),
.Y(n_800)
);

INVx1_ASAP7_75t_L g801 ( 
.A(n_735),
.Y(n_801)
);

INVx1_ASAP7_75t_L g802 ( 
.A(n_450),
.Y(n_802)
);

INVx2_ASAP7_75t_L g803 ( 
.A(n_721),
.Y(n_803)
);

CKINVDCx20_ASAP7_75t_R g804 ( 
.A(n_700),
.Y(n_804)
);

INVxp33_ASAP7_75t_L g805 ( 
.A(n_515),
.Y(n_805)
);

INVxp67_ASAP7_75t_L g806 ( 
.A(n_727),
.Y(n_806)
);

INVx1_ASAP7_75t_L g807 ( 
.A(n_450),
.Y(n_807)
);

INVx1_ASAP7_75t_L g808 ( 
.A(n_514),
.Y(n_808)
);

INVx1_ASAP7_75t_L g809 ( 
.A(n_514),
.Y(n_809)
);

INVx1_ASAP7_75t_L g810 ( 
.A(n_519),
.Y(n_810)
);

INVx1_ASAP7_75t_L g811 ( 
.A(n_519),
.Y(n_811)
);

INVx1_ASAP7_75t_L g812 ( 
.A(n_565),
.Y(n_812)
);

INVx1_ASAP7_75t_SL g813 ( 
.A(n_469),
.Y(n_813)
);

INVx1_ASAP7_75t_L g814 ( 
.A(n_565),
.Y(n_814)
);

CKINVDCx20_ASAP7_75t_R g815 ( 
.A(n_712),
.Y(n_815)
);

CKINVDCx5p33_ASAP7_75t_R g816 ( 
.A(n_563),
.Y(n_816)
);

INVx1_ASAP7_75t_L g817 ( 
.A(n_638),
.Y(n_817)
);

INVx1_ASAP7_75t_L g818 ( 
.A(n_638),
.Y(n_818)
);

INVx1_ASAP7_75t_L g819 ( 
.A(n_646),
.Y(n_819)
);

INVx1_ASAP7_75t_L g820 ( 
.A(n_646),
.Y(n_820)
);

BUFx3_ASAP7_75t_L g821 ( 
.A(n_449),
.Y(n_821)
);

CKINVDCx5p33_ASAP7_75t_R g822 ( 
.A(n_563),
.Y(n_822)
);

INVxp33_ASAP7_75t_L g823 ( 
.A(n_515),
.Y(n_823)
);

INVx1_ASAP7_75t_L g824 ( 
.A(n_453),
.Y(n_824)
);

INVx1_ASAP7_75t_L g825 ( 
.A(n_458),
.Y(n_825)
);

CKINVDCx5p33_ASAP7_75t_R g826 ( 
.A(n_471),
.Y(n_826)
);

INVx1_ASAP7_75t_L g827 ( 
.A(n_474),
.Y(n_827)
);

INVx1_ASAP7_75t_L g828 ( 
.A(n_481),
.Y(n_828)
);

INVx1_ASAP7_75t_L g829 ( 
.A(n_484),
.Y(n_829)
);

BUFx3_ASAP7_75t_L g830 ( 
.A(n_520),
.Y(n_830)
);

HB1xp67_ASAP7_75t_L g831 ( 
.A(n_475),
.Y(n_831)
);

INVxp67_ASAP7_75t_SL g832 ( 
.A(n_703),
.Y(n_832)
);

INVxp33_ASAP7_75t_SL g833 ( 
.A(n_479),
.Y(n_833)
);

BUFx3_ASAP7_75t_L g834 ( 
.A(n_520),
.Y(n_834)
);

CKINVDCx5p33_ASAP7_75t_R g835 ( 
.A(n_480),
.Y(n_835)
);

INVx1_ASAP7_75t_L g836 ( 
.A(n_489),
.Y(n_836)
);

CKINVDCx5p33_ASAP7_75t_R g837 ( 
.A(n_482),
.Y(n_837)
);

CKINVDCx5p33_ASAP7_75t_R g838 ( 
.A(n_487),
.Y(n_838)
);

INVx1_ASAP7_75t_L g839 ( 
.A(n_500),
.Y(n_839)
);

INVx1_ASAP7_75t_L g840 ( 
.A(n_501),
.Y(n_840)
);

CKINVDCx20_ASAP7_75t_R g841 ( 
.A(n_727),
.Y(n_841)
);

INVxp67_ASAP7_75t_L g842 ( 
.A(n_492),
.Y(n_842)
);

INVx1_ASAP7_75t_L g843 ( 
.A(n_512),
.Y(n_843)
);

INVx1_ASAP7_75t_L g844 ( 
.A(n_518),
.Y(n_844)
);

CKINVDCx20_ASAP7_75t_R g845 ( 
.A(n_751),
.Y(n_845)
);

OA21x2_ASAP7_75t_L g846 ( 
.A1(n_745),
.A2(n_701),
.B(n_460),
.Y(n_846)
);

HB1xp67_ASAP7_75t_L g847 ( 
.A(n_750),
.Y(n_847)
);

AND2x2_ASAP7_75t_L g848 ( 
.A(n_782),
.B(n_498),
.Y(n_848)
);

INVx2_ASAP7_75t_L g849 ( 
.A(n_752),
.Y(n_849)
);

INVx2_ASAP7_75t_L g850 ( 
.A(n_752),
.Y(n_850)
);

BUFx6f_ASAP7_75t_L g851 ( 
.A(n_821),
.Y(n_851)
);

AND2x4_ASAP7_75t_L g852 ( 
.A(n_744),
.B(n_515),
.Y(n_852)
);

NAND2xp5_ASAP7_75t_L g853 ( 
.A(n_761),
.B(n_506),
.Y(n_853)
);

NOR2xp33_ASAP7_75t_L g854 ( 
.A(n_755),
.B(n_509),
.Y(n_854)
);

INVx6_ASAP7_75t_L g855 ( 
.A(n_821),
.Y(n_855)
);

INVx1_ASAP7_75t_L g856 ( 
.A(n_767),
.Y(n_856)
);

BUFx3_ASAP7_75t_L g857 ( 
.A(n_830),
.Y(n_857)
);

AND2x4_ASAP7_75t_L g858 ( 
.A(n_746),
.B(n_515),
.Y(n_858)
);

INVx3_ASAP7_75t_L g859 ( 
.A(n_830),
.Y(n_859)
);

CKINVDCx20_ASAP7_75t_R g860 ( 
.A(n_751),
.Y(n_860)
);

AND2x2_ASAP7_75t_L g861 ( 
.A(n_782),
.B(n_503),
.Y(n_861)
);

INVx1_ASAP7_75t_L g862 ( 
.A(n_768),
.Y(n_862)
);

OAI22xp5_ASAP7_75t_SL g863 ( 
.A1(n_759),
.A2(n_511),
.B1(n_531),
.B2(n_517),
.Y(n_863)
);

BUFx6f_ASAP7_75t_L g864 ( 
.A(n_834),
.Y(n_864)
);

AND2x4_ASAP7_75t_L g865 ( 
.A(n_756),
.B(n_802),
.Y(n_865)
);

BUFx6f_ASAP7_75t_L g866 ( 
.A(n_834),
.Y(n_866)
);

OAI22xp5_ASAP7_75t_SL g867 ( 
.A1(n_759),
.A2(n_540),
.B1(n_541),
.B2(n_532),
.Y(n_867)
);

INVx1_ASAP7_75t_L g868 ( 
.A(n_769),
.Y(n_868)
);

INVx1_ASAP7_75t_L g869 ( 
.A(n_748),
.Y(n_869)
);

AND2x4_ASAP7_75t_L g870 ( 
.A(n_807),
.B(n_586),
.Y(n_870)
);

INVx1_ASAP7_75t_L g871 ( 
.A(n_747),
.Y(n_871)
);

INVx1_ASAP7_75t_L g872 ( 
.A(n_757),
.Y(n_872)
);

INVx3_ASAP7_75t_L g873 ( 
.A(n_745),
.Y(n_873)
);

AOI22xp5_ASAP7_75t_L g874 ( 
.A1(n_785),
.A2(n_548),
.B1(n_549),
.B2(n_545),
.Y(n_874)
);

INVx1_ASAP7_75t_L g875 ( 
.A(n_758),
.Y(n_875)
);

BUFx3_ASAP7_75t_L g876 ( 
.A(n_808),
.Y(n_876)
);

HB1xp67_ASAP7_75t_L g877 ( 
.A(n_775),
.Y(n_877)
);

AND2x2_ASAP7_75t_L g878 ( 
.A(n_773),
.B(n_551),
.Y(n_878)
);

BUFx2_ASAP7_75t_L g879 ( 
.A(n_826),
.Y(n_879)
);

BUFx3_ASAP7_75t_L g880 ( 
.A(n_809),
.Y(n_880)
);

BUFx6f_ASAP7_75t_L g881 ( 
.A(n_754),
.Y(n_881)
);

NAND2x1_ASAP7_75t_L g882 ( 
.A(n_810),
.B(n_544),
.Y(n_882)
);

BUFx6f_ASAP7_75t_L g883 ( 
.A(n_754),
.Y(n_883)
);

CKINVDCx5p33_ASAP7_75t_R g884 ( 
.A(n_743),
.Y(n_884)
);

INVx5_ASAP7_75t_L g885 ( 
.A(n_764),
.Y(n_885)
);

NAND2xp5_ASAP7_75t_L g886 ( 
.A(n_799),
.B(n_547),
.Y(n_886)
);

INVx2_ASAP7_75t_L g887 ( 
.A(n_764),
.Y(n_887)
);

NAND2xp5_ASAP7_75t_L g888 ( 
.A(n_800),
.B(n_559),
.Y(n_888)
);

BUFx6f_ASAP7_75t_L g889 ( 
.A(n_803),
.Y(n_889)
);

BUFx6f_ASAP7_75t_L g890 ( 
.A(n_803),
.Y(n_890)
);

BUFx2_ASAP7_75t_L g891 ( 
.A(n_835),
.Y(n_891)
);

INVx1_ASAP7_75t_L g892 ( 
.A(n_770),
.Y(n_892)
);

INVx2_ASAP7_75t_L g893 ( 
.A(n_762),
.Y(n_893)
);

INVx2_ASAP7_75t_L g894 ( 
.A(n_763),
.Y(n_894)
);

AND2x4_ASAP7_75t_L g895 ( 
.A(n_811),
.B(n_586),
.Y(n_895)
);

INVx1_ASAP7_75t_L g896 ( 
.A(n_771),
.Y(n_896)
);

OA21x2_ASAP7_75t_L g897 ( 
.A1(n_824),
.A2(n_701),
.B(n_460),
.Y(n_897)
);

INVx1_ASAP7_75t_L g898 ( 
.A(n_772),
.Y(n_898)
);

INVx2_ASAP7_75t_L g899 ( 
.A(n_765),
.Y(n_899)
);

INVx1_ASAP7_75t_L g900 ( 
.A(n_774),
.Y(n_900)
);

INVxp67_ASAP7_75t_L g901 ( 
.A(n_831),
.Y(n_901)
);

INVx1_ASAP7_75t_L g902 ( 
.A(n_776),
.Y(n_902)
);

AND2x2_ASAP7_75t_L g903 ( 
.A(n_749),
.B(n_554),
.Y(n_903)
);

INVx1_ASAP7_75t_L g904 ( 
.A(n_777),
.Y(n_904)
);

AOI22xp5_ASAP7_75t_L g905 ( 
.A1(n_832),
.A2(n_833),
.B1(n_787),
.B2(n_837),
.Y(n_905)
);

INVx2_ASAP7_75t_L g906 ( 
.A(n_784),
.Y(n_906)
);

NAND2xp5_ASAP7_75t_SL g907 ( 
.A(n_816),
.B(n_561),
.Y(n_907)
);

BUFx6f_ASAP7_75t_L g908 ( 
.A(n_786),
.Y(n_908)
);

NAND2xp5_ASAP7_75t_SL g909 ( 
.A(n_822),
.B(n_812),
.Y(n_909)
);

BUFx3_ASAP7_75t_L g910 ( 
.A(n_814),
.Y(n_910)
);

INVx2_ASAP7_75t_L g911 ( 
.A(n_788),
.Y(n_911)
);

AND2x2_ASAP7_75t_L g912 ( 
.A(n_813),
.B(n_562),
.Y(n_912)
);

AOI22xp5_ASAP7_75t_L g913 ( 
.A1(n_838),
.A2(n_591),
.B1(n_601),
.B2(n_580),
.Y(n_913)
);

INVx1_ASAP7_75t_L g914 ( 
.A(n_789),
.Y(n_914)
);

INVx2_ASAP7_75t_L g915 ( 
.A(n_791),
.Y(n_915)
);

INVx1_ASAP7_75t_L g916 ( 
.A(n_793),
.Y(n_916)
);

OA21x2_ASAP7_75t_L g917 ( 
.A1(n_825),
.A2(n_530),
.B(n_529),
.Y(n_917)
);

INVx1_ASAP7_75t_L g918 ( 
.A(n_794),
.Y(n_918)
);

INVx2_ASAP7_75t_L g919 ( 
.A(n_795),
.Y(n_919)
);

AND2x2_ASAP7_75t_L g920 ( 
.A(n_842),
.B(n_602),
.Y(n_920)
);

CKINVDCx5p33_ASAP7_75t_R g921 ( 
.A(n_753),
.Y(n_921)
);

INVx1_ASAP7_75t_L g922 ( 
.A(n_796),
.Y(n_922)
);

AND2x2_ASAP7_75t_L g923 ( 
.A(n_806),
.B(n_817),
.Y(n_923)
);

INVx1_ASAP7_75t_L g924 ( 
.A(n_797),
.Y(n_924)
);

INVx2_ASAP7_75t_L g925 ( 
.A(n_798),
.Y(n_925)
);

CKINVDCx20_ASAP7_75t_R g926 ( 
.A(n_778),
.Y(n_926)
);

INVx1_ASAP7_75t_L g927 ( 
.A(n_801),
.Y(n_927)
);

BUFx8_ASAP7_75t_L g928 ( 
.A(n_818),
.Y(n_928)
);

HB1xp67_ASAP7_75t_L g929 ( 
.A(n_827),
.Y(n_929)
);

INVx1_ASAP7_75t_L g930 ( 
.A(n_828),
.Y(n_930)
);

AND2x6_ASAP7_75t_L g931 ( 
.A(n_829),
.B(n_526),
.Y(n_931)
);

INVx1_ASAP7_75t_L g932 ( 
.A(n_836),
.Y(n_932)
);

CKINVDCx5p33_ASAP7_75t_R g933 ( 
.A(n_760),
.Y(n_933)
);

INVx1_ASAP7_75t_L g934 ( 
.A(n_839),
.Y(n_934)
);

INVx2_ASAP7_75t_L g935 ( 
.A(n_840),
.Y(n_935)
);

NAND2xp5_ASAP7_75t_L g936 ( 
.A(n_843),
.B(n_844),
.Y(n_936)
);

INVx2_ASAP7_75t_L g937 ( 
.A(n_819),
.Y(n_937)
);

NAND2xp5_ASAP7_75t_L g938 ( 
.A(n_820),
.B(n_577),
.Y(n_938)
);

OA21x2_ASAP7_75t_L g939 ( 
.A1(n_805),
.A2(n_542),
.B(n_533),
.Y(n_939)
);

INVx2_ASAP7_75t_L g940 ( 
.A(n_805),
.Y(n_940)
);

INVx1_ASAP7_75t_L g941 ( 
.A(n_823),
.Y(n_941)
);

BUFx6f_ASAP7_75t_L g942 ( 
.A(n_823),
.Y(n_942)
);

INVxp67_ASAP7_75t_L g943 ( 
.A(n_766),
.Y(n_943)
);

NOR2xp33_ASAP7_75t_L g944 ( 
.A(n_815),
.B(n_684),
.Y(n_944)
);

INVx2_ASAP7_75t_L g945 ( 
.A(n_841),
.Y(n_945)
);

INVx2_ASAP7_75t_L g946 ( 
.A(n_841),
.Y(n_946)
);

INVx2_ASAP7_75t_L g947 ( 
.A(n_815),
.Y(n_947)
);

NAND2xp5_ASAP7_75t_L g948 ( 
.A(n_779),
.B(n_705),
.Y(n_948)
);

OR2x2_ASAP7_75t_L g949 ( 
.A(n_783),
.B(n_491),
.Y(n_949)
);

INVx3_ASAP7_75t_L g950 ( 
.A(n_792),
.Y(n_950)
);

AND2x2_ASAP7_75t_L g951 ( 
.A(n_792),
.B(n_604),
.Y(n_951)
);

INVx2_ASAP7_75t_L g952 ( 
.A(n_804),
.Y(n_952)
);

INVx1_ASAP7_75t_L g953 ( 
.A(n_804),
.Y(n_953)
);

NAND2xp5_ASAP7_75t_L g954 ( 
.A(n_778),
.B(n_455),
.Y(n_954)
);

INVx3_ASAP7_75t_L g955 ( 
.A(n_780),
.Y(n_955)
);

INVx3_ASAP7_75t_L g956 ( 
.A(n_780),
.Y(n_956)
);

BUFx6f_ASAP7_75t_L g957 ( 
.A(n_781),
.Y(n_957)
);

INVx1_ASAP7_75t_L g958 ( 
.A(n_781),
.Y(n_958)
);

INVx1_ASAP7_75t_L g959 ( 
.A(n_790),
.Y(n_959)
);

INVx1_ASAP7_75t_L g960 ( 
.A(n_790),
.Y(n_960)
);

BUFx6f_ASAP7_75t_L g961 ( 
.A(n_752),
.Y(n_961)
);

OAI22xp5_ASAP7_75t_L g962 ( 
.A1(n_782),
.A2(n_617),
.B1(n_621),
.B2(n_606),
.Y(n_962)
);

AND2x2_ASAP7_75t_L g963 ( 
.A(n_750),
.B(n_624),
.Y(n_963)
);

INVx2_ASAP7_75t_L g964 ( 
.A(n_752),
.Y(n_964)
);

NAND2xp5_ASAP7_75t_SL g965 ( 
.A(n_816),
.B(n_703),
.Y(n_965)
);

INVxp67_ASAP7_75t_L g966 ( 
.A(n_750),
.Y(n_966)
);

OA21x2_ASAP7_75t_L g967 ( 
.A1(n_745),
.A2(n_553),
.B(n_543),
.Y(n_967)
);

INVx1_ASAP7_75t_L g968 ( 
.A(n_767),
.Y(n_968)
);

AND2x2_ASAP7_75t_L g969 ( 
.A(n_750),
.B(n_629),
.Y(n_969)
);

BUFx6f_ASAP7_75t_L g970 ( 
.A(n_752),
.Y(n_970)
);

INVx1_ASAP7_75t_L g971 ( 
.A(n_767),
.Y(n_971)
);

INVxp67_ASAP7_75t_L g972 ( 
.A(n_750),
.Y(n_972)
);

CKINVDCx5p33_ASAP7_75t_R g973 ( 
.A(n_743),
.Y(n_973)
);

BUFx8_ASAP7_75t_L g974 ( 
.A(n_744),
.Y(n_974)
);

AND2x2_ASAP7_75t_L g975 ( 
.A(n_750),
.B(n_643),
.Y(n_975)
);

INVx3_ASAP7_75t_L g976 ( 
.A(n_752),
.Y(n_976)
);

BUFx6f_ASAP7_75t_L g977 ( 
.A(n_752),
.Y(n_977)
);

INVx1_ASAP7_75t_L g978 ( 
.A(n_767),
.Y(n_978)
);

INVx2_ASAP7_75t_L g979 ( 
.A(n_752),
.Y(n_979)
);

INVx1_ASAP7_75t_L g980 ( 
.A(n_767),
.Y(n_980)
);

INVx2_ASAP7_75t_L g981 ( 
.A(n_752),
.Y(n_981)
);

INVx1_ASAP7_75t_L g982 ( 
.A(n_767),
.Y(n_982)
);

HB1xp67_ASAP7_75t_L g983 ( 
.A(n_750),
.Y(n_983)
);

CKINVDCx5p33_ASAP7_75t_R g984 ( 
.A(n_743),
.Y(n_984)
);

INVx2_ASAP7_75t_L g985 ( 
.A(n_752),
.Y(n_985)
);

OAI22xp5_ASAP7_75t_L g986 ( 
.A1(n_782),
.A2(n_658),
.B1(n_667),
.B2(n_652),
.Y(n_986)
);

INVx2_ASAP7_75t_L g987 ( 
.A(n_752),
.Y(n_987)
);

INVx1_ASAP7_75t_L g988 ( 
.A(n_767),
.Y(n_988)
);

INVx1_ASAP7_75t_L g989 ( 
.A(n_767),
.Y(n_989)
);

AND2x4_ASAP7_75t_L g990 ( 
.A(n_744),
.B(n_586),
.Y(n_990)
);

INVx2_ASAP7_75t_L g991 ( 
.A(n_752),
.Y(n_991)
);

INVx3_ASAP7_75t_L g992 ( 
.A(n_752),
.Y(n_992)
);

INVx2_ASAP7_75t_L g993 ( 
.A(n_752),
.Y(n_993)
);

CKINVDCx5p33_ASAP7_75t_R g994 ( 
.A(n_743),
.Y(n_994)
);

INVx2_ASAP7_75t_L g995 ( 
.A(n_752),
.Y(n_995)
);

INVx4_ASAP7_75t_L g996 ( 
.A(n_752),
.Y(n_996)
);

INVx1_ASAP7_75t_L g997 ( 
.A(n_767),
.Y(n_997)
);

INVx2_ASAP7_75t_L g998 ( 
.A(n_752),
.Y(n_998)
);

INVx1_ASAP7_75t_L g999 ( 
.A(n_767),
.Y(n_999)
);

HB1xp67_ASAP7_75t_L g1000 ( 
.A(n_750),
.Y(n_1000)
);

INVx2_ASAP7_75t_L g1001 ( 
.A(n_752),
.Y(n_1001)
);

HB1xp67_ASAP7_75t_L g1002 ( 
.A(n_813),
.Y(n_1002)
);

NAND2xp5_ASAP7_75t_L g1003 ( 
.A(n_761),
.B(n_493),
.Y(n_1003)
);

BUFx6f_ASAP7_75t_L g1004 ( 
.A(n_752),
.Y(n_1004)
);

INVx1_ASAP7_75t_L g1005 ( 
.A(n_767),
.Y(n_1005)
);

INVx1_ASAP7_75t_L g1006 ( 
.A(n_767),
.Y(n_1006)
);

NAND3xp33_ASAP7_75t_L g1007 ( 
.A(n_917),
.B(n_560),
.C(n_557),
.Y(n_1007)
);

INVx1_ASAP7_75t_L g1008 ( 
.A(n_940),
.Y(n_1008)
);

INVx2_ASAP7_75t_SL g1009 ( 
.A(n_1002),
.Y(n_1009)
);

INVx4_ASAP7_75t_L g1010 ( 
.A(n_942),
.Y(n_1010)
);

INVx2_ASAP7_75t_L g1011 ( 
.A(n_851),
.Y(n_1011)
);

INVx2_ASAP7_75t_L g1012 ( 
.A(n_851),
.Y(n_1012)
);

CKINVDCx5p33_ASAP7_75t_R g1013 ( 
.A(n_845),
.Y(n_1013)
);

BUFx3_ASAP7_75t_L g1014 ( 
.A(n_942),
.Y(n_1014)
);

NAND2xp33_ASAP7_75t_L g1015 ( 
.A(n_931),
.B(n_929),
.Y(n_1015)
);

AOI22xp5_ASAP7_75t_L g1016 ( 
.A1(n_929),
.A2(n_689),
.B1(n_691),
.B2(n_676),
.Y(n_1016)
);

INVx2_ASAP7_75t_L g1017 ( 
.A(n_851),
.Y(n_1017)
);

INVx2_ASAP7_75t_L g1018 ( 
.A(n_864),
.Y(n_1018)
);

INVx2_ASAP7_75t_L g1019 ( 
.A(n_864),
.Y(n_1019)
);

INVx5_ASAP7_75t_L g1020 ( 
.A(n_942),
.Y(n_1020)
);

INVx2_ASAP7_75t_L g1021 ( 
.A(n_864),
.Y(n_1021)
);

INVx2_ASAP7_75t_L g1022 ( 
.A(n_866),
.Y(n_1022)
);

INVx2_ASAP7_75t_L g1023 ( 
.A(n_866),
.Y(n_1023)
);

INVx3_ASAP7_75t_L g1024 ( 
.A(n_852),
.Y(n_1024)
);

INVx1_ASAP7_75t_L g1025 ( 
.A(n_941),
.Y(n_1025)
);

AND3x2_ASAP7_75t_L g1026 ( 
.A(n_943),
.B(n_570),
.C(n_564),
.Y(n_1026)
);

INVx1_ASAP7_75t_L g1027 ( 
.A(n_870),
.Y(n_1027)
);

NAND2xp33_ASAP7_75t_SL g1028 ( 
.A(n_879),
.B(n_706),
.Y(n_1028)
);

INVx1_ASAP7_75t_L g1029 ( 
.A(n_870),
.Y(n_1029)
);

INVx2_ASAP7_75t_L g1030 ( 
.A(n_866),
.Y(n_1030)
);

AND2x6_ASAP7_75t_L g1031 ( 
.A(n_869),
.B(n_526),
.Y(n_1031)
);

INVx1_ASAP7_75t_L g1032 ( 
.A(n_895),
.Y(n_1032)
);

INVx3_ASAP7_75t_L g1033 ( 
.A(n_852),
.Y(n_1033)
);

BUFx10_ASAP7_75t_L g1034 ( 
.A(n_944),
.Y(n_1034)
);

INVx2_ASAP7_75t_L g1035 ( 
.A(n_961),
.Y(n_1035)
);

NAND2xp5_ASAP7_75t_SL g1036 ( 
.A(n_848),
.B(n_861),
.Y(n_1036)
);

INVx1_ASAP7_75t_L g1037 ( 
.A(n_895),
.Y(n_1037)
);

INVx2_ASAP7_75t_L g1038 ( 
.A(n_961),
.Y(n_1038)
);

INVx2_ASAP7_75t_L g1039 ( 
.A(n_961),
.Y(n_1039)
);

BUFx16f_ASAP7_75t_R g1040 ( 
.A(n_974),
.Y(n_1040)
);

INVx2_ASAP7_75t_L g1041 ( 
.A(n_970),
.Y(n_1041)
);

INVx1_ASAP7_75t_L g1042 ( 
.A(n_858),
.Y(n_1042)
);

INVx1_ASAP7_75t_L g1043 ( 
.A(n_858),
.Y(n_1043)
);

BUFx6f_ASAP7_75t_L g1044 ( 
.A(n_970),
.Y(n_1044)
);

INVx2_ASAP7_75t_L g1045 ( 
.A(n_970),
.Y(n_1045)
);

INVx2_ASAP7_75t_L g1046 ( 
.A(n_977),
.Y(n_1046)
);

INVx1_ASAP7_75t_L g1047 ( 
.A(n_990),
.Y(n_1047)
);

INVx2_ASAP7_75t_L g1048 ( 
.A(n_977),
.Y(n_1048)
);

INVx2_ASAP7_75t_SL g1049 ( 
.A(n_847),
.Y(n_1049)
);

NAND2xp5_ASAP7_75t_L g1050 ( 
.A(n_930),
.B(n_571),
.Y(n_1050)
);

BUFx3_ASAP7_75t_L g1051 ( 
.A(n_891),
.Y(n_1051)
);

OAI22xp5_ASAP7_75t_L g1052 ( 
.A1(n_905),
.A2(n_729),
.B1(n_730),
.B2(n_710),
.Y(n_1052)
);

INVx1_ASAP7_75t_L g1053 ( 
.A(n_990),
.Y(n_1053)
);

INVx2_ASAP7_75t_L g1054 ( 
.A(n_977),
.Y(n_1054)
);

INVx4_ASAP7_75t_L g1055 ( 
.A(n_855),
.Y(n_1055)
);

CKINVDCx5p33_ASAP7_75t_R g1056 ( 
.A(n_860),
.Y(n_1056)
);

NOR2xp33_ASAP7_75t_L g1057 ( 
.A(n_965),
.B(n_583),
.Y(n_1057)
);

INVx1_ASAP7_75t_L g1058 ( 
.A(n_856),
.Y(n_1058)
);

INVx3_ASAP7_75t_L g1059 ( 
.A(n_859),
.Y(n_1059)
);

NOR2x1p5_ASAP7_75t_L g1060 ( 
.A(n_884),
.B(n_734),
.Y(n_1060)
);

INVx2_ASAP7_75t_L g1061 ( 
.A(n_1004),
.Y(n_1061)
);

INVx2_ASAP7_75t_L g1062 ( 
.A(n_1004),
.Y(n_1062)
);

INVx1_ASAP7_75t_L g1063 ( 
.A(n_862),
.Y(n_1063)
);

INVx2_ASAP7_75t_L g1064 ( 
.A(n_1004),
.Y(n_1064)
);

INVx1_ASAP7_75t_L g1065 ( 
.A(n_868),
.Y(n_1065)
);

NAND2xp5_ASAP7_75t_L g1066 ( 
.A(n_932),
.B(n_451),
.Y(n_1066)
);

HB1xp67_ASAP7_75t_L g1067 ( 
.A(n_847),
.Y(n_1067)
);

AND2x2_ASAP7_75t_L g1068 ( 
.A(n_966),
.B(n_737),
.Y(n_1068)
);

OR2x2_ASAP7_75t_L g1069 ( 
.A(n_983),
.B(n_516),
.Y(n_1069)
);

AND2x4_ASAP7_75t_L g1070 ( 
.A(n_876),
.B(n_741),
.Y(n_1070)
);

BUFx10_ASAP7_75t_L g1071 ( 
.A(n_983),
.Y(n_1071)
);

BUFx3_ASAP7_75t_L g1072 ( 
.A(n_855),
.Y(n_1072)
);

INVx2_ASAP7_75t_L g1073 ( 
.A(n_859),
.Y(n_1073)
);

INVx1_ASAP7_75t_L g1074 ( 
.A(n_1006),
.Y(n_1074)
);

INVx1_ASAP7_75t_L g1075 ( 
.A(n_968),
.Y(n_1075)
);

INVx2_ASAP7_75t_SL g1076 ( 
.A(n_1000),
.Y(n_1076)
);

AOI22xp33_ASAP7_75t_SL g1077 ( 
.A1(n_974),
.A2(n_690),
.B1(n_473),
.B2(n_586),
.Y(n_1077)
);

CKINVDCx5p33_ASAP7_75t_R g1078 ( 
.A(n_926),
.Y(n_1078)
);

INVx2_ASAP7_75t_SL g1079 ( 
.A(n_1000),
.Y(n_1079)
);

NOR2xp33_ASAP7_75t_L g1080 ( 
.A(n_907),
.B(n_659),
.Y(n_1080)
);

NOR2xp33_ASAP7_75t_L g1081 ( 
.A(n_909),
.B(n_665),
.Y(n_1081)
);

NAND3xp33_ASAP7_75t_L g1082 ( 
.A(n_917),
.B(n_581),
.C(n_579),
.Y(n_1082)
);

NAND2xp5_ASAP7_75t_L g1083 ( 
.A(n_934),
.B(n_456),
.Y(n_1083)
);

INVx2_ASAP7_75t_SL g1084 ( 
.A(n_877),
.Y(n_1084)
);

INVx2_ASAP7_75t_L g1085 ( 
.A(n_976),
.Y(n_1085)
);

INVx2_ASAP7_75t_L g1086 ( 
.A(n_976),
.Y(n_1086)
);

INVx1_ASAP7_75t_L g1087 ( 
.A(n_1005),
.Y(n_1087)
);

INVxp33_ASAP7_75t_L g1088 ( 
.A(n_877),
.Y(n_1088)
);

INVx2_ASAP7_75t_L g1089 ( 
.A(n_992),
.Y(n_1089)
);

INVx2_ASAP7_75t_L g1090 ( 
.A(n_992),
.Y(n_1090)
);

BUFx10_ASAP7_75t_L g1091 ( 
.A(n_865),
.Y(n_1091)
);

INVx1_ASAP7_75t_L g1092 ( 
.A(n_971),
.Y(n_1092)
);

AOI22xp33_ASAP7_75t_SL g1093 ( 
.A1(n_863),
.A2(n_616),
.B1(n_556),
.B2(n_459),
.Y(n_1093)
);

NOR2xp33_ASAP7_75t_L g1094 ( 
.A(n_923),
.B(n_685),
.Y(n_1094)
);

INVx1_ASAP7_75t_L g1095 ( 
.A(n_978),
.Y(n_1095)
);

INVx2_ASAP7_75t_L g1096 ( 
.A(n_849),
.Y(n_1096)
);

INVx2_ASAP7_75t_L g1097 ( 
.A(n_850),
.Y(n_1097)
);

INVx2_ASAP7_75t_L g1098 ( 
.A(n_964),
.Y(n_1098)
);

NAND2xp33_ASAP7_75t_R g1099 ( 
.A(n_921),
.B(n_457),
.Y(n_1099)
);

INVx1_ASAP7_75t_L g1100 ( 
.A(n_980),
.Y(n_1100)
);

INVx2_ASAP7_75t_L g1101 ( 
.A(n_979),
.Y(n_1101)
);

INVx2_ASAP7_75t_L g1102 ( 
.A(n_981),
.Y(n_1102)
);

INVx5_ASAP7_75t_L g1103 ( 
.A(n_931),
.Y(n_1103)
);

INVx1_ASAP7_75t_L g1104 ( 
.A(n_982),
.Y(n_1104)
);

INVx1_ASAP7_75t_L g1105 ( 
.A(n_988),
.Y(n_1105)
);

INVx1_ASAP7_75t_L g1106 ( 
.A(n_989),
.Y(n_1106)
);

AND3x2_ASAP7_75t_L g1107 ( 
.A(n_943),
.B(n_596),
.C(n_592),
.Y(n_1107)
);

INVx8_ASAP7_75t_L g1108 ( 
.A(n_931),
.Y(n_1108)
);

INVx1_ASAP7_75t_L g1109 ( 
.A(n_997),
.Y(n_1109)
);

CKINVDCx5p33_ASAP7_75t_R g1110 ( 
.A(n_933),
.Y(n_1110)
);

INVx1_ASAP7_75t_L g1111 ( 
.A(n_999),
.Y(n_1111)
);

AND2x2_ASAP7_75t_L g1112 ( 
.A(n_966),
.B(n_556),
.Y(n_1112)
);

INVx5_ASAP7_75t_L g1113 ( 
.A(n_931),
.Y(n_1113)
);

CKINVDCx5p33_ASAP7_75t_R g1114 ( 
.A(n_973),
.Y(n_1114)
);

OAI22xp33_ASAP7_75t_L g1115 ( 
.A1(n_905),
.A2(n_605),
.B1(n_608),
.B2(n_599),
.Y(n_1115)
);

INVx1_ASAP7_75t_L g1116 ( 
.A(n_908),
.Y(n_1116)
);

INVx1_ASAP7_75t_L g1117 ( 
.A(n_908),
.Y(n_1117)
);

INVx2_ASAP7_75t_SL g1118 ( 
.A(n_865),
.Y(n_1118)
);

INVx4_ASAP7_75t_L g1119 ( 
.A(n_996),
.Y(n_1119)
);

NOR2x1p5_ASAP7_75t_L g1120 ( 
.A(n_984),
.B(n_462),
.Y(n_1120)
);

INVx2_ASAP7_75t_L g1121 ( 
.A(n_985),
.Y(n_1121)
);

OAI22xp33_ASAP7_75t_L g1122 ( 
.A1(n_972),
.A2(n_615),
.B1(n_631),
.B2(n_613),
.Y(n_1122)
);

NAND2xp5_ASAP7_75t_SL g1123 ( 
.A(n_937),
.B(n_464),
.Y(n_1123)
);

NAND2xp33_ASAP7_75t_L g1124 ( 
.A(n_881),
.B(n_721),
.Y(n_1124)
);

INVx3_ASAP7_75t_L g1125 ( 
.A(n_908),
.Y(n_1125)
);

INVx1_ASAP7_75t_L g1126 ( 
.A(n_893),
.Y(n_1126)
);

NAND2xp5_ASAP7_75t_SL g1127 ( 
.A(n_920),
.B(n_466),
.Y(n_1127)
);

CKINVDCx5p33_ASAP7_75t_R g1128 ( 
.A(n_994),
.Y(n_1128)
);

CKINVDCx6p67_ASAP7_75t_R g1129 ( 
.A(n_957),
.Y(n_1129)
);

CKINVDCx5p33_ASAP7_75t_R g1130 ( 
.A(n_928),
.Y(n_1130)
);

NAND2xp5_ASAP7_75t_SL g1131 ( 
.A(n_901),
.B(n_467),
.Y(n_1131)
);

INVx1_ASAP7_75t_L g1132 ( 
.A(n_894),
.Y(n_1132)
);

NAND2xp5_ASAP7_75t_L g1133 ( 
.A(n_892),
.B(n_632),
.Y(n_1133)
);

INVx1_ASAP7_75t_L g1134 ( 
.A(n_899),
.Y(n_1134)
);

INVx1_ASAP7_75t_L g1135 ( 
.A(n_875),
.Y(n_1135)
);

CKINVDCx5p33_ASAP7_75t_R g1136 ( 
.A(n_928),
.Y(n_1136)
);

INVx2_ASAP7_75t_SL g1137 ( 
.A(n_963),
.Y(n_1137)
);

AND2x2_ASAP7_75t_L g1138 ( 
.A(n_972),
.B(n_616),
.Y(n_1138)
);

INVx1_ASAP7_75t_L g1139 ( 
.A(n_871),
.Y(n_1139)
);

NAND2xp5_ASAP7_75t_SL g1140 ( 
.A(n_901),
.B(n_468),
.Y(n_1140)
);

NAND2xp5_ASAP7_75t_L g1141 ( 
.A(n_896),
.B(n_633),
.Y(n_1141)
);

NAND2xp5_ASAP7_75t_SL g1142 ( 
.A(n_912),
.B(n_470),
.Y(n_1142)
);

OAI22xp5_ASAP7_75t_L g1143 ( 
.A1(n_936),
.A2(n_656),
.B1(n_663),
.B2(n_648),
.Y(n_1143)
);

INVx2_ASAP7_75t_L g1144 ( 
.A(n_987),
.Y(n_1144)
);

INVx1_ASAP7_75t_L g1145 ( 
.A(n_906),
.Y(n_1145)
);

NAND2xp5_ASAP7_75t_SL g1146 ( 
.A(n_857),
.B(n_472),
.Y(n_1146)
);

NAND2xp5_ASAP7_75t_L g1147 ( 
.A(n_898),
.B(n_664),
.Y(n_1147)
);

INVx1_ASAP7_75t_L g1148 ( 
.A(n_911),
.Y(n_1148)
);

NAND2xp5_ASAP7_75t_SL g1149 ( 
.A(n_880),
.B(n_476),
.Y(n_1149)
);

INVx2_ASAP7_75t_L g1150 ( 
.A(n_991),
.Y(n_1150)
);

AND2x6_ASAP7_75t_L g1151 ( 
.A(n_910),
.B(n_669),
.Y(n_1151)
);

INVx2_ASAP7_75t_L g1152 ( 
.A(n_993),
.Y(n_1152)
);

INVx1_ASAP7_75t_L g1153 ( 
.A(n_915),
.Y(n_1153)
);

INVx2_ASAP7_75t_L g1154 ( 
.A(n_995),
.Y(n_1154)
);

INVxp67_ASAP7_75t_SL g1155 ( 
.A(n_936),
.Y(n_1155)
);

NAND2xp5_ASAP7_75t_SL g1156 ( 
.A(n_948),
.B(n_477),
.Y(n_1156)
);

INVx1_ASAP7_75t_L g1157 ( 
.A(n_919),
.Y(n_1157)
);

INVx2_ASAP7_75t_L g1158 ( 
.A(n_998),
.Y(n_1158)
);

AOI22xp33_ASAP7_75t_L g1159 ( 
.A1(n_872),
.A2(n_688),
.B1(n_699),
.B2(n_679),
.Y(n_1159)
);

NAND2xp5_ASAP7_75t_L g1160 ( 
.A(n_900),
.B(n_702),
.Y(n_1160)
);

INVx2_ASAP7_75t_L g1161 ( 
.A(n_1001),
.Y(n_1161)
);

INVx3_ASAP7_75t_L g1162 ( 
.A(n_996),
.Y(n_1162)
);

INVx2_ASAP7_75t_L g1163 ( 
.A(n_881),
.Y(n_1163)
);

BUFx6f_ASAP7_75t_SL g1164 ( 
.A(n_957),
.Y(n_1164)
);

INVxp67_ASAP7_75t_SL g1165 ( 
.A(n_967),
.Y(n_1165)
);

INVx2_ASAP7_75t_L g1166 ( 
.A(n_881),
.Y(n_1166)
);

INVx5_ASAP7_75t_L g1167 ( 
.A(n_883),
.Y(n_1167)
);

NAND3xp33_ASAP7_75t_L g1168 ( 
.A(n_967),
.B(n_713),
.C(n_711),
.Y(n_1168)
);

OR2x6_ASAP7_75t_L g1169 ( 
.A(n_863),
.B(n_716),
.Y(n_1169)
);

INVx2_ASAP7_75t_L g1170 ( 
.A(n_883),
.Y(n_1170)
);

NOR2x1p5_ASAP7_75t_L g1171 ( 
.A(n_945),
.B(n_483),
.Y(n_1171)
);

BUFx6f_ASAP7_75t_L g1172 ( 
.A(n_883),
.Y(n_1172)
);

INVx2_ASAP7_75t_L g1173 ( 
.A(n_889),
.Y(n_1173)
);

INVx1_ASAP7_75t_L g1174 ( 
.A(n_925),
.Y(n_1174)
);

NAND2xp33_ASAP7_75t_SL g1175 ( 
.A(n_882),
.B(n_486),
.Y(n_1175)
);

INVx1_ASAP7_75t_L g1176 ( 
.A(n_935),
.Y(n_1176)
);

AOI21x1_ASAP7_75t_L g1177 ( 
.A1(n_939),
.A2(n_725),
.B(n_722),
.Y(n_1177)
);

NOR2xp33_ASAP7_75t_L g1178 ( 
.A(n_853),
.B(n_494),
.Y(n_1178)
);

BUFx3_ASAP7_75t_L g1179 ( 
.A(n_885),
.Y(n_1179)
);

BUFx6f_ASAP7_75t_L g1180 ( 
.A(n_889),
.Y(n_1180)
);

AOI22xp33_ASAP7_75t_L g1181 ( 
.A1(n_902),
.A2(n_728),
.B1(n_736),
.B2(n_726),
.Y(n_1181)
);

NAND2xp5_ASAP7_75t_L g1182 ( 
.A(n_904),
.B(n_495),
.Y(n_1182)
);

INVx2_ASAP7_75t_L g1183 ( 
.A(n_889),
.Y(n_1183)
);

AOI22xp5_ASAP7_75t_L g1184 ( 
.A1(n_914),
.A2(n_738),
.B1(n_502),
.B2(n_504),
.Y(n_1184)
);

OR2x6_ASAP7_75t_L g1185 ( 
.A(n_867),
.B(n_946),
.Y(n_1185)
);

NAND3xp33_ASAP7_75t_L g1186 ( 
.A(n_897),
.B(n_534),
.C(n_496),
.Y(n_1186)
);

INVx2_ASAP7_75t_SL g1187 ( 
.A(n_969),
.Y(n_1187)
);

AOI22xp33_ASAP7_75t_L g1188 ( 
.A1(n_916),
.A2(n_576),
.B1(n_612),
.B2(n_575),
.Y(n_1188)
);

INVx2_ASAP7_75t_L g1189 ( 
.A(n_890),
.Y(n_1189)
);

NAND2xp33_ASAP7_75t_L g1190 ( 
.A(n_890),
.B(n_721),
.Y(n_1190)
);

INVx1_ASAP7_75t_L g1191 ( 
.A(n_918),
.Y(n_1191)
);

NAND3xp33_ASAP7_75t_L g1192 ( 
.A(n_897),
.B(n_657),
.C(n_647),
.Y(n_1192)
);

NAND2xp5_ASAP7_75t_SL g1193 ( 
.A(n_948),
.B(n_497),
.Y(n_1193)
);

NOR2x1p5_ASAP7_75t_L g1194 ( 
.A(n_950),
.B(n_505),
.Y(n_1194)
);

INVx1_ASAP7_75t_L g1195 ( 
.A(n_922),
.Y(n_1195)
);

INVx1_ASAP7_75t_L g1196 ( 
.A(n_924),
.Y(n_1196)
);

NAND3xp33_ASAP7_75t_L g1197 ( 
.A(n_846),
.B(n_740),
.C(n_508),
.Y(n_1197)
);

CKINVDCx6p67_ASAP7_75t_R g1198 ( 
.A(n_957),
.Y(n_1198)
);

AND2x4_ASAP7_75t_L g1199 ( 
.A(n_938),
.B(n_507),
.Y(n_1199)
);

AOI22xp33_ASAP7_75t_L g1200 ( 
.A1(n_927),
.A2(n_510),
.B1(n_521),
.B2(n_513),
.Y(n_1200)
);

NOR2xp33_ASAP7_75t_L g1201 ( 
.A(n_853),
.B(n_522),
.Y(n_1201)
);

NAND2xp5_ASAP7_75t_SL g1202 ( 
.A(n_962),
.B(n_525),
.Y(n_1202)
);

INVx1_ASAP7_75t_L g1203 ( 
.A(n_938),
.Y(n_1203)
);

NAND2xp5_ASAP7_75t_SL g1204 ( 
.A(n_962),
.B(n_528),
.Y(n_1204)
);

CKINVDCx5p33_ASAP7_75t_R g1205 ( 
.A(n_986),
.Y(n_1205)
);

INVx2_ASAP7_75t_L g1206 ( 
.A(n_890),
.Y(n_1206)
);

BUFx3_ASAP7_75t_L g1207 ( 
.A(n_885),
.Y(n_1207)
);

INVx2_ASAP7_75t_L g1208 ( 
.A(n_873),
.Y(n_1208)
);

INVx1_ASAP7_75t_L g1209 ( 
.A(n_886),
.Y(n_1209)
);

AND2x2_ASAP7_75t_SL g1210 ( 
.A(n_951),
.B(n_461),
.Y(n_1210)
);

NAND2xp5_ASAP7_75t_SL g1211 ( 
.A(n_986),
.B(n_546),
.Y(n_1211)
);

INVx1_ASAP7_75t_L g1212 ( 
.A(n_886),
.Y(n_1212)
);

INVx4_ASAP7_75t_L g1213 ( 
.A(n_873),
.Y(n_1213)
);

INVx1_ASAP7_75t_L g1214 ( 
.A(n_888),
.Y(n_1214)
);

OAI21xp33_ASAP7_75t_SL g1215 ( 
.A1(n_1003),
.A2(n_0),
.B(n_2),
.Y(n_1215)
);

INVx3_ASAP7_75t_L g1216 ( 
.A(n_846),
.Y(n_1216)
);

NOR3xp33_ASAP7_75t_L g1217 ( 
.A(n_867),
.B(n_558),
.C(n_550),
.Y(n_1217)
);

INVx4_ASAP7_75t_L g1218 ( 
.A(n_885),
.Y(n_1218)
);

INVx1_ASAP7_75t_L g1219 ( 
.A(n_888),
.Y(n_1219)
);

INVx2_ASAP7_75t_L g1220 ( 
.A(n_887),
.Y(n_1220)
);

NAND2xp5_ASAP7_75t_SL g1221 ( 
.A(n_1003),
.B(n_566),
.Y(n_1221)
);

OAI22xp33_ASAP7_75t_R g1222 ( 
.A1(n_958),
.A2(n_5),
.B1(n_3),
.B2(n_4),
.Y(n_1222)
);

INVx2_ASAP7_75t_SL g1223 ( 
.A(n_975),
.Y(n_1223)
);

NOR2xp33_ASAP7_75t_L g1224 ( 
.A(n_854),
.B(n_567),
.Y(n_1224)
);

INVx2_ASAP7_75t_L g1225 ( 
.A(n_939),
.Y(n_1225)
);

OAI22xp33_ASAP7_75t_SL g1226 ( 
.A1(n_954),
.A2(n_569),
.B1(n_572),
.B2(n_568),
.Y(n_1226)
);

NOR2xp33_ASAP7_75t_L g1227 ( 
.A(n_878),
.B(n_573),
.Y(n_1227)
);

BUFx3_ASAP7_75t_L g1228 ( 
.A(n_903),
.Y(n_1228)
);

NAND2xp5_ASAP7_75t_L g1229 ( 
.A(n_874),
.B(n_574),
.Y(n_1229)
);

INVx1_ASAP7_75t_L g1230 ( 
.A(n_874),
.Y(n_1230)
);

CKINVDCx5p33_ASAP7_75t_R g1231 ( 
.A(n_955),
.Y(n_1231)
);

AND2x2_ASAP7_75t_L g1232 ( 
.A(n_913),
.B(n_742),
.Y(n_1232)
);

INVx1_ASAP7_75t_L g1233 ( 
.A(n_954),
.Y(n_1233)
);

AOI22xp33_ASAP7_75t_L g1234 ( 
.A1(n_913),
.A2(n_585),
.B1(n_588),
.B2(n_578),
.Y(n_1234)
);

INVx2_ASAP7_75t_L g1235 ( 
.A(n_949),
.Y(n_1235)
);

INVx2_ASAP7_75t_L g1236 ( 
.A(n_947),
.Y(n_1236)
);

NOR2xp33_ASAP7_75t_L g1237 ( 
.A(n_1088),
.B(n_952),
.Y(n_1237)
);

INVxp67_ASAP7_75t_L g1238 ( 
.A(n_1009),
.Y(n_1238)
);

INVx1_ASAP7_75t_L g1239 ( 
.A(n_1155),
.Y(n_1239)
);

HB1xp67_ASAP7_75t_L g1240 ( 
.A(n_1067),
.Y(n_1240)
);

INVx2_ASAP7_75t_L g1241 ( 
.A(n_1044),
.Y(n_1241)
);

NAND2xp5_ASAP7_75t_L g1242 ( 
.A(n_1209),
.B(n_593),
.Y(n_1242)
);

BUFx3_ASAP7_75t_L g1243 ( 
.A(n_1051),
.Y(n_1243)
);

AOI22xp5_ASAP7_75t_L g1244 ( 
.A1(n_1203),
.A2(n_953),
.B1(n_960),
.B2(n_959),
.Y(n_1244)
);

NOR2xp33_ASAP7_75t_L g1245 ( 
.A(n_1049),
.B(n_950),
.Y(n_1245)
);

NAND2xp5_ASAP7_75t_L g1246 ( 
.A(n_1212),
.B(n_594),
.Y(n_1246)
);

INVx1_ASAP7_75t_L g1247 ( 
.A(n_1191),
.Y(n_1247)
);

INVx1_ASAP7_75t_L g1248 ( 
.A(n_1195),
.Y(n_1248)
);

INVx2_ASAP7_75t_L g1249 ( 
.A(n_1044),
.Y(n_1249)
);

NAND2xp5_ASAP7_75t_L g1250 ( 
.A(n_1214),
.B(n_595),
.Y(n_1250)
);

NAND2xp5_ASAP7_75t_SL g1251 ( 
.A(n_1071),
.B(n_597),
.Y(n_1251)
);

INVx3_ASAP7_75t_L g1252 ( 
.A(n_1213),
.Y(n_1252)
);

INVx1_ASAP7_75t_L g1253 ( 
.A(n_1196),
.Y(n_1253)
);

AND2x2_ASAP7_75t_L g1254 ( 
.A(n_1071),
.B(n_955),
.Y(n_1254)
);

INVx4_ASAP7_75t_L g1255 ( 
.A(n_1091),
.Y(n_1255)
);

NAND2xp5_ASAP7_75t_SL g1256 ( 
.A(n_1076),
.B(n_598),
.Y(n_1256)
);

INVx1_ASAP7_75t_L g1257 ( 
.A(n_1058),
.Y(n_1257)
);

INVx1_ASAP7_75t_L g1258 ( 
.A(n_1063),
.Y(n_1258)
);

NAND2xp5_ASAP7_75t_L g1259 ( 
.A(n_1219),
.B(n_600),
.Y(n_1259)
);

AOI22xp5_ASAP7_75t_L g1260 ( 
.A1(n_1233),
.A2(n_618),
.B1(n_619),
.B2(n_611),
.Y(n_1260)
);

NAND2xp5_ASAP7_75t_L g1261 ( 
.A(n_1199),
.B(n_622),
.Y(n_1261)
);

NAND3xp33_ASAP7_75t_L g1262 ( 
.A(n_1186),
.B(n_527),
.C(n_461),
.Y(n_1262)
);

INVx1_ASAP7_75t_L g1263 ( 
.A(n_1065),
.Y(n_1263)
);

NAND2xp33_ASAP7_75t_L g1264 ( 
.A(n_1108),
.B(n_623),
.Y(n_1264)
);

NOR2xp33_ASAP7_75t_L g1265 ( 
.A(n_1079),
.B(n_956),
.Y(n_1265)
);

NAND3xp33_ASAP7_75t_L g1266 ( 
.A(n_1186),
.B(n_527),
.C(n_461),
.Y(n_1266)
);

NAND2xp5_ASAP7_75t_L g1267 ( 
.A(n_1199),
.B(n_625),
.Y(n_1267)
);

NAND2xp33_ASAP7_75t_L g1268 ( 
.A(n_1108),
.B(n_1151),
.Y(n_1268)
);

NAND2xp5_ASAP7_75t_L g1269 ( 
.A(n_1112),
.B(n_627),
.Y(n_1269)
);

BUFx6f_ASAP7_75t_L g1270 ( 
.A(n_1108),
.Y(n_1270)
);

HB1xp67_ASAP7_75t_L g1271 ( 
.A(n_1084),
.Y(n_1271)
);

NAND2xp5_ASAP7_75t_L g1272 ( 
.A(n_1139),
.B(n_628),
.Y(n_1272)
);

NAND2xp5_ASAP7_75t_L g1273 ( 
.A(n_1138),
.B(n_630),
.Y(n_1273)
);

OR2x2_ASAP7_75t_L g1274 ( 
.A(n_1069),
.B(n_956),
.Y(n_1274)
);

AND2x2_ASAP7_75t_L g1275 ( 
.A(n_1235),
.B(n_3),
.Y(n_1275)
);

INVx2_ASAP7_75t_L g1276 ( 
.A(n_1044),
.Y(n_1276)
);

BUFx3_ASAP7_75t_L g1277 ( 
.A(n_1129),
.Y(n_1277)
);

NOR2x1p5_ASAP7_75t_L g1278 ( 
.A(n_1130),
.B(n_634),
.Y(n_1278)
);

NAND2xp5_ASAP7_75t_SL g1279 ( 
.A(n_1091),
.B(n_636),
.Y(n_1279)
);

NAND2xp5_ASAP7_75t_L g1280 ( 
.A(n_1178),
.B(n_639),
.Y(n_1280)
);

NOR2xp33_ASAP7_75t_SL g1281 ( 
.A(n_1165),
.B(n_640),
.Y(n_1281)
);

NAND2xp5_ASAP7_75t_L g1282 ( 
.A(n_1201),
.B(n_641),
.Y(n_1282)
);

INVx2_ASAP7_75t_L g1283 ( 
.A(n_1096),
.Y(n_1283)
);

INVxp67_ASAP7_75t_SL g1284 ( 
.A(n_1118),
.Y(n_1284)
);

A2O1A1Ixp33_ASAP7_75t_L g1285 ( 
.A1(n_1074),
.A2(n_527),
.B(n_582),
.C(n_461),
.Y(n_1285)
);

INVx2_ASAP7_75t_L g1286 ( 
.A(n_1097),
.Y(n_1286)
);

NOR2xp33_ASAP7_75t_L g1287 ( 
.A(n_1137),
.B(n_642),
.Y(n_1287)
);

INVx1_ASAP7_75t_L g1288 ( 
.A(n_1075),
.Y(n_1288)
);

INVx2_ASAP7_75t_L g1289 ( 
.A(n_1098),
.Y(n_1289)
);

NAND2xp5_ASAP7_75t_SL g1290 ( 
.A(n_1103),
.B(n_644),
.Y(n_1290)
);

NAND2xp5_ASAP7_75t_SL g1291 ( 
.A(n_1103),
.B(n_739),
.Y(n_1291)
);

NOR2xp33_ASAP7_75t_SL g1292 ( 
.A(n_1103),
.B(n_645),
.Y(n_1292)
);

NAND2xp33_ASAP7_75t_L g1293 ( 
.A(n_1151),
.B(n_649),
.Y(n_1293)
);

INVx1_ASAP7_75t_L g1294 ( 
.A(n_1087),
.Y(n_1294)
);

NAND2xp5_ASAP7_75t_L g1295 ( 
.A(n_1092),
.B(n_650),
.Y(n_1295)
);

INVx2_ASAP7_75t_SL g1296 ( 
.A(n_1070),
.Y(n_1296)
);

NOR2xp33_ASAP7_75t_L g1297 ( 
.A(n_1187),
.B(n_653),
.Y(n_1297)
);

NOR3xp33_ASAP7_75t_SL g1298 ( 
.A(n_1136),
.B(n_660),
.C(n_654),
.Y(n_1298)
);

NOR2xp33_ASAP7_75t_SL g1299 ( 
.A(n_1113),
.B(n_662),
.Y(n_1299)
);

INVx1_ASAP7_75t_L g1300 ( 
.A(n_1095),
.Y(n_1300)
);

NOR3xp33_ASAP7_75t_L g1301 ( 
.A(n_1052),
.B(n_671),
.C(n_668),
.Y(n_1301)
);

BUFx6f_ASAP7_75t_L g1302 ( 
.A(n_1113),
.Y(n_1302)
);

INVx1_ASAP7_75t_L g1303 ( 
.A(n_1100),
.Y(n_1303)
);

OR2x2_ASAP7_75t_L g1304 ( 
.A(n_1052),
.B(n_5),
.Y(n_1304)
);

INVx2_ASAP7_75t_SL g1305 ( 
.A(n_1070),
.Y(n_1305)
);

INVx2_ASAP7_75t_L g1306 ( 
.A(n_1101),
.Y(n_1306)
);

NOR2xp67_ASAP7_75t_L g1307 ( 
.A(n_1110),
.B(n_6),
.Y(n_1307)
);

INVx2_ASAP7_75t_L g1308 ( 
.A(n_1102),
.Y(n_1308)
);

AOI22xp33_ASAP7_75t_L g1309 ( 
.A1(n_1230),
.A2(n_1205),
.B1(n_1036),
.B2(n_1210),
.Y(n_1309)
);

INVxp67_ASAP7_75t_L g1310 ( 
.A(n_1068),
.Y(n_1310)
);

INVx2_ASAP7_75t_L g1311 ( 
.A(n_1121),
.Y(n_1311)
);

INVx1_ASAP7_75t_L g1312 ( 
.A(n_1104),
.Y(n_1312)
);

INVx2_ASAP7_75t_L g1313 ( 
.A(n_1144),
.Y(n_1313)
);

INVx2_ASAP7_75t_L g1314 ( 
.A(n_1150),
.Y(n_1314)
);

NOR2xp33_ASAP7_75t_L g1315 ( 
.A(n_1223),
.B(n_673),
.Y(n_1315)
);

NAND2xp5_ASAP7_75t_L g1316 ( 
.A(n_1105),
.B(n_675),
.Y(n_1316)
);

CKINVDCx5p33_ASAP7_75t_R g1317 ( 
.A(n_1114),
.Y(n_1317)
);

NOR2xp33_ASAP7_75t_L g1318 ( 
.A(n_1232),
.B(n_677),
.Y(n_1318)
);

INVx2_ASAP7_75t_L g1319 ( 
.A(n_1152),
.Y(n_1319)
);

INVx2_ASAP7_75t_L g1320 ( 
.A(n_1154),
.Y(n_1320)
);

NOR2x1p5_ASAP7_75t_L g1321 ( 
.A(n_1040),
.B(n_678),
.Y(n_1321)
);

AO221x1_ASAP7_75t_L g1322 ( 
.A1(n_1040),
.A2(n_587),
.B1(n_610),
.B2(n_582),
.C(n_527),
.Y(n_1322)
);

NAND2xp5_ASAP7_75t_SL g1323 ( 
.A(n_1113),
.B(n_680),
.Y(n_1323)
);

OAI22xp33_ASAP7_75t_L g1324 ( 
.A1(n_1169),
.A2(n_1185),
.B1(n_1016),
.B2(n_1128),
.Y(n_1324)
);

NAND2xp5_ASAP7_75t_L g1325 ( 
.A(n_1106),
.B(n_683),
.Y(n_1325)
);

INVx1_ASAP7_75t_L g1326 ( 
.A(n_1109),
.Y(n_1326)
);

INVx2_ASAP7_75t_L g1327 ( 
.A(n_1158),
.Y(n_1327)
);

NOR2xp33_ASAP7_75t_L g1328 ( 
.A(n_1229),
.B(n_693),
.Y(n_1328)
);

AND2x2_ASAP7_75t_L g1329 ( 
.A(n_1016),
.B(n_8),
.Y(n_1329)
);

AND2x2_ASAP7_75t_L g1330 ( 
.A(n_1228),
.B(n_10),
.Y(n_1330)
);

NAND2xp5_ASAP7_75t_SL g1331 ( 
.A(n_1213),
.B(n_1226),
.Y(n_1331)
);

INVxp67_ASAP7_75t_L g1332 ( 
.A(n_1099),
.Y(n_1332)
);

INVx1_ASAP7_75t_L g1333 ( 
.A(n_1111),
.Y(n_1333)
);

NAND2xp5_ASAP7_75t_L g1334 ( 
.A(n_1025),
.B(n_1135),
.Y(n_1334)
);

NAND2xp5_ASAP7_75t_L g1335 ( 
.A(n_1145),
.B(n_694),
.Y(n_1335)
);

NAND2xp5_ASAP7_75t_L g1336 ( 
.A(n_1148),
.B(n_1153),
.Y(n_1336)
);

NAND2xp5_ASAP7_75t_SL g1337 ( 
.A(n_1226),
.B(n_723),
.Y(n_1337)
);

INVx1_ASAP7_75t_L g1338 ( 
.A(n_1024),
.Y(n_1338)
);

INVx1_ASAP7_75t_L g1339 ( 
.A(n_1024),
.Y(n_1339)
);

NAND2xp5_ASAP7_75t_L g1340 ( 
.A(n_1157),
.B(n_695),
.Y(n_1340)
);

INVx2_ASAP7_75t_L g1341 ( 
.A(n_1161),
.Y(n_1341)
);

NAND2xp5_ASAP7_75t_L g1342 ( 
.A(n_1174),
.B(n_698),
.Y(n_1342)
);

AOI22xp33_ASAP7_75t_L g1343 ( 
.A1(n_1202),
.A2(n_714),
.B1(n_715),
.B2(n_708),
.Y(n_1343)
);

BUFx6f_ASAP7_75t_L g1344 ( 
.A(n_1172),
.Y(n_1344)
);

AOI22xp5_ASAP7_75t_L g1345 ( 
.A1(n_1222),
.A2(n_719),
.B1(n_718),
.B2(n_587),
.Y(n_1345)
);

NAND2xp5_ASAP7_75t_L g1346 ( 
.A(n_1176),
.B(n_10),
.Y(n_1346)
);

AND2x2_ASAP7_75t_L g1347 ( 
.A(n_1034),
.B(n_11),
.Y(n_1347)
);

NAND2xp5_ASAP7_75t_SL g1348 ( 
.A(n_1028),
.B(n_582),
.Y(n_1348)
);

NAND2xp5_ASAP7_75t_L g1349 ( 
.A(n_1151),
.B(n_13),
.Y(n_1349)
);

INVx2_ASAP7_75t_L g1350 ( 
.A(n_1208),
.Y(n_1350)
);

INVx1_ASAP7_75t_L g1351 ( 
.A(n_1033),
.Y(n_1351)
);

INVx1_ASAP7_75t_L g1352 ( 
.A(n_1033),
.Y(n_1352)
);

AND2x2_ASAP7_75t_L g1353 ( 
.A(n_1034),
.B(n_13),
.Y(n_1353)
);

INVxp67_ASAP7_75t_SL g1354 ( 
.A(n_1015),
.Y(n_1354)
);

INVx1_ASAP7_75t_L g1355 ( 
.A(n_1027),
.Y(n_1355)
);

NAND2xp5_ASAP7_75t_SL g1356 ( 
.A(n_1020),
.B(n_582),
.Y(n_1356)
);

INVx2_ASAP7_75t_L g1357 ( 
.A(n_1073),
.Y(n_1357)
);

NOR2xp33_ASAP7_75t_L g1358 ( 
.A(n_1229),
.B(n_15),
.Y(n_1358)
);

OAI22xp5_ASAP7_75t_L g1359 ( 
.A1(n_1050),
.A2(n_717),
.B1(n_610),
.B2(n_614),
.Y(n_1359)
);

NAND2xp5_ASAP7_75t_SL g1360 ( 
.A(n_1020),
.B(n_587),
.Y(n_1360)
);

NAND2xp5_ASAP7_75t_L g1361 ( 
.A(n_1151),
.B(n_15),
.Y(n_1361)
);

BUFx6f_ASAP7_75t_L g1362 ( 
.A(n_1172),
.Y(n_1362)
);

AOI22xp33_ASAP7_75t_L g1363 ( 
.A1(n_1204),
.A2(n_610),
.B1(n_614),
.B2(n_587),
.Y(n_1363)
);

NAND2xp5_ASAP7_75t_L g1364 ( 
.A(n_1126),
.B(n_16),
.Y(n_1364)
);

INVx2_ASAP7_75t_L g1365 ( 
.A(n_1085),
.Y(n_1365)
);

NOR3xp33_ASAP7_75t_L g1366 ( 
.A(n_1115),
.B(n_17),
.C(n_18),
.Y(n_1366)
);

NOR2x1p5_ASAP7_75t_L g1367 ( 
.A(n_1013),
.B(n_610),
.Y(n_1367)
);

INVx1_ASAP7_75t_L g1368 ( 
.A(n_1029),
.Y(n_1368)
);

INVx1_ASAP7_75t_L g1369 ( 
.A(n_1032),
.Y(n_1369)
);

NAND3xp33_ASAP7_75t_L g1370 ( 
.A(n_1192),
.B(n_626),
.C(n_614),
.Y(n_1370)
);

INVx2_ASAP7_75t_L g1371 ( 
.A(n_1086),
.Y(n_1371)
);

NAND2xp5_ASAP7_75t_L g1372 ( 
.A(n_1132),
.B(n_18),
.Y(n_1372)
);

NAND2x1p5_ASAP7_75t_L g1373 ( 
.A(n_1020),
.B(n_614),
.Y(n_1373)
);

AND2x4_ASAP7_75t_L g1374 ( 
.A(n_1194),
.B(n_19),
.Y(n_1374)
);

BUFx3_ASAP7_75t_L g1375 ( 
.A(n_1198),
.Y(n_1375)
);

NAND2xp5_ASAP7_75t_L g1376 ( 
.A(n_1134),
.B(n_20),
.Y(n_1376)
);

NOR2x1_ASAP7_75t_L g1377 ( 
.A(n_1060),
.B(n_626),
.Y(n_1377)
);

INVx2_ASAP7_75t_L g1378 ( 
.A(n_1089),
.Y(n_1378)
);

OAI22xp5_ASAP7_75t_L g1379 ( 
.A1(n_1050),
.A2(n_717),
.B1(n_626),
.B2(n_22),
.Y(n_1379)
);

INVxp67_ASAP7_75t_L g1380 ( 
.A(n_1094),
.Y(n_1380)
);

NAND2xp5_ASAP7_75t_SL g1381 ( 
.A(n_1184),
.B(n_626),
.Y(n_1381)
);

CKINVDCx5p33_ASAP7_75t_R g1382 ( 
.A(n_1056),
.Y(n_1382)
);

INVx2_ASAP7_75t_L g1383 ( 
.A(n_1090),
.Y(n_1383)
);

INVx2_ASAP7_75t_L g1384 ( 
.A(n_1059),
.Y(n_1384)
);

NAND2xp5_ASAP7_75t_L g1385 ( 
.A(n_1184),
.B(n_20),
.Y(n_1385)
);

NAND2xp5_ASAP7_75t_L g1386 ( 
.A(n_1008),
.B(n_21),
.Y(n_1386)
);

OR2x2_ASAP7_75t_L g1387 ( 
.A(n_1078),
.B(n_21),
.Y(n_1387)
);

INVxp67_ASAP7_75t_L g1388 ( 
.A(n_1227),
.Y(n_1388)
);

NAND2xp5_ASAP7_75t_L g1389 ( 
.A(n_1143),
.B(n_23),
.Y(n_1389)
);

INVx3_ASAP7_75t_L g1390 ( 
.A(n_1119),
.Y(n_1390)
);

INVx2_ASAP7_75t_L g1391 ( 
.A(n_1059),
.Y(n_1391)
);

NAND2xp5_ASAP7_75t_SL g1392 ( 
.A(n_1119),
.B(n_717),
.Y(n_1392)
);

INVx2_ASAP7_75t_L g1393 ( 
.A(n_1216),
.Y(n_1393)
);

INVxp67_ASAP7_75t_L g1394 ( 
.A(n_1164),
.Y(n_1394)
);

NOR2xp33_ASAP7_75t_L g1395 ( 
.A(n_1142),
.B(n_24),
.Y(n_1395)
);

CKINVDCx5p33_ASAP7_75t_R g1396 ( 
.A(n_1164),
.Y(n_1396)
);

NOR2xp33_ASAP7_75t_L g1397 ( 
.A(n_1131),
.B(n_25),
.Y(n_1397)
);

NAND2xp5_ASAP7_75t_L g1398 ( 
.A(n_1143),
.B(n_26),
.Y(n_1398)
);

BUFx4f_ASAP7_75t_L g1399 ( 
.A(n_1169),
.Y(n_1399)
);

AOI22xp5_ASAP7_75t_L g1400 ( 
.A1(n_1215),
.A2(n_717),
.B1(n_30),
.B2(n_28),
.Y(n_1400)
);

AOI22xp5_ASAP7_75t_L g1401 ( 
.A1(n_1215),
.A2(n_31),
.B1(n_29),
.B2(n_30),
.Y(n_1401)
);

NAND2xp5_ASAP7_75t_SL g1402 ( 
.A(n_1218),
.B(n_32),
.Y(n_1402)
);

INVx1_ASAP7_75t_L g1403 ( 
.A(n_1037),
.Y(n_1403)
);

BUFx6f_ASAP7_75t_L g1404 ( 
.A(n_1172),
.Y(n_1404)
);

NAND2xp5_ASAP7_75t_SL g1405 ( 
.A(n_1218),
.B(n_32),
.Y(n_1405)
);

NAND2xp5_ASAP7_75t_L g1406 ( 
.A(n_1133),
.B(n_33),
.Y(n_1406)
);

NOR2xp67_ASAP7_75t_L g1407 ( 
.A(n_1231),
.B(n_33),
.Y(n_1407)
);

NOR2xp33_ASAP7_75t_L g1408 ( 
.A(n_1140),
.B(n_34),
.Y(n_1408)
);

OR2x2_ASAP7_75t_L g1409 ( 
.A(n_1185),
.B(n_35),
.Y(n_1409)
);

INVx2_ASAP7_75t_L g1410 ( 
.A(n_1216),
.Y(n_1410)
);

INVx1_ASAP7_75t_L g1411 ( 
.A(n_1042),
.Y(n_1411)
);

INVx1_ASAP7_75t_L g1412 ( 
.A(n_1043),
.Y(n_1412)
);

INVx2_ASAP7_75t_L g1413 ( 
.A(n_1162),
.Y(n_1413)
);

NOR3xp33_ASAP7_75t_L g1414 ( 
.A(n_1217),
.B(n_35),
.C(n_36),
.Y(n_1414)
);

NAND2xp5_ASAP7_75t_L g1415 ( 
.A(n_1133),
.B(n_37),
.Y(n_1415)
);

AND2x4_ASAP7_75t_L g1416 ( 
.A(n_1194),
.B(n_37),
.Y(n_1416)
);

INVx2_ASAP7_75t_L g1417 ( 
.A(n_1162),
.Y(n_1417)
);

AOI22xp33_ASAP7_75t_L g1418 ( 
.A1(n_1211),
.A2(n_41),
.B1(n_38),
.B2(n_39),
.Y(n_1418)
);

AOI22xp33_ASAP7_75t_L g1419 ( 
.A1(n_1169),
.A2(n_43),
.B1(n_39),
.B2(n_41),
.Y(n_1419)
);

NAND2xp5_ASAP7_75t_SL g1420 ( 
.A(n_1066),
.B(n_44),
.Y(n_1420)
);

NOR2xp33_ASAP7_75t_L g1421 ( 
.A(n_1127),
.B(n_44),
.Y(n_1421)
);

AOI22xp33_ASAP7_75t_L g1422 ( 
.A1(n_1236),
.A2(n_47),
.B1(n_45),
.B2(n_46),
.Y(n_1422)
);

NAND2xp5_ASAP7_75t_L g1423 ( 
.A(n_1141),
.B(n_45),
.Y(n_1423)
);

INVx2_ASAP7_75t_L g1424 ( 
.A(n_1220),
.Y(n_1424)
);

NOR2xp33_ASAP7_75t_L g1425 ( 
.A(n_1156),
.B(n_47),
.Y(n_1425)
);

INVx2_ASAP7_75t_L g1426 ( 
.A(n_1125),
.Y(n_1426)
);

NAND2xp5_ASAP7_75t_L g1427 ( 
.A(n_1141),
.B(n_1147),
.Y(n_1427)
);

INVx2_ASAP7_75t_L g1428 ( 
.A(n_1125),
.Y(n_1428)
);

NAND2xp5_ASAP7_75t_L g1429 ( 
.A(n_1147),
.B(n_49),
.Y(n_1429)
);

INVxp67_ASAP7_75t_L g1430 ( 
.A(n_1031),
.Y(n_1430)
);

AND2x2_ASAP7_75t_SL g1431 ( 
.A(n_1234),
.B(n_1055),
.Y(n_1431)
);

NAND2xp5_ASAP7_75t_L g1432 ( 
.A(n_1160),
.B(n_49),
.Y(n_1432)
);

INVx1_ASAP7_75t_L g1433 ( 
.A(n_1047),
.Y(n_1433)
);

AOI22xp5_ASAP7_75t_L g1434 ( 
.A1(n_1380),
.A2(n_1185),
.B1(n_1060),
.B2(n_1122),
.Y(n_1434)
);

INVx1_ASAP7_75t_L g1435 ( 
.A(n_1239),
.Y(n_1435)
);

INVx4_ASAP7_75t_L g1436 ( 
.A(n_1255),
.Y(n_1436)
);

INVx1_ASAP7_75t_SL g1437 ( 
.A(n_1243),
.Y(n_1437)
);

INVx1_ASAP7_75t_L g1438 ( 
.A(n_1247),
.Y(n_1438)
);

NAND2xp5_ASAP7_75t_L g1439 ( 
.A(n_1427),
.B(n_1159),
.Y(n_1439)
);

O2A1O1Ixp33_ASAP7_75t_L g1440 ( 
.A1(n_1389),
.A2(n_1160),
.B(n_1193),
.C(n_1221),
.Y(n_1440)
);

INVx5_ASAP7_75t_L g1441 ( 
.A(n_1255),
.Y(n_1441)
);

BUFx6f_ASAP7_75t_L g1442 ( 
.A(n_1344),
.Y(n_1442)
);

INVx2_ASAP7_75t_SL g1443 ( 
.A(n_1277),
.Y(n_1443)
);

OAI22xp5_ASAP7_75t_L g1444 ( 
.A1(n_1309),
.A2(n_1225),
.B1(n_1053),
.B2(n_1181),
.Y(n_1444)
);

HB1xp67_ASAP7_75t_L g1445 ( 
.A(n_1240),
.Y(n_1445)
);

INVx2_ASAP7_75t_L g1446 ( 
.A(n_1248),
.Y(n_1446)
);

BUFx2_ASAP7_75t_L g1447 ( 
.A(n_1271),
.Y(n_1447)
);

NAND2xp5_ASAP7_75t_L g1448 ( 
.A(n_1253),
.B(n_1057),
.Y(n_1448)
);

INVx2_ASAP7_75t_L g1449 ( 
.A(n_1257),
.Y(n_1449)
);

INVx2_ASAP7_75t_L g1450 ( 
.A(n_1258),
.Y(n_1450)
);

AOI22xp33_ASAP7_75t_L g1451 ( 
.A1(n_1399),
.A2(n_1093),
.B1(n_1171),
.B2(n_1031),
.Y(n_1451)
);

BUFx3_ASAP7_75t_L g1452 ( 
.A(n_1375),
.Y(n_1452)
);

NAND2xp5_ASAP7_75t_SL g1453 ( 
.A(n_1238),
.B(n_1077),
.Y(n_1453)
);

BUFx6f_ASAP7_75t_L g1454 ( 
.A(n_1344),
.Y(n_1454)
);

INVx2_ASAP7_75t_SL g1455 ( 
.A(n_1396),
.Y(n_1455)
);

NAND2xp5_ASAP7_75t_SL g1456 ( 
.A(n_1281),
.B(n_1200),
.Y(n_1456)
);

NAND2xp5_ASAP7_75t_L g1457 ( 
.A(n_1263),
.B(n_1081),
.Y(n_1457)
);

AOI21xp5_ASAP7_75t_L g1458 ( 
.A1(n_1334),
.A2(n_1192),
.B(n_1197),
.Y(n_1458)
);

INVx3_ASAP7_75t_L g1459 ( 
.A(n_1270),
.Y(n_1459)
);

INVx1_ASAP7_75t_L g1460 ( 
.A(n_1288),
.Y(n_1460)
);

INVx2_ASAP7_75t_L g1461 ( 
.A(n_1294),
.Y(n_1461)
);

INVx1_ASAP7_75t_L g1462 ( 
.A(n_1300),
.Y(n_1462)
);

AND3x2_ASAP7_75t_SL g1463 ( 
.A(n_1321),
.B(n_1120),
.C(n_1107),
.Y(n_1463)
);

AOI22xp33_ASAP7_75t_L g1464 ( 
.A1(n_1399),
.A2(n_1171),
.B1(n_1031),
.B2(n_1120),
.Y(n_1464)
);

OR2x2_ASAP7_75t_L g1465 ( 
.A(n_1274),
.B(n_1072),
.Y(n_1465)
);

AOI22xp33_ASAP7_75t_L g1466 ( 
.A1(n_1329),
.A2(n_1031),
.B1(n_1080),
.B2(n_1224),
.Y(n_1466)
);

INVx2_ASAP7_75t_L g1467 ( 
.A(n_1303),
.Y(n_1467)
);

OR2x6_ASAP7_75t_L g1468 ( 
.A(n_1409),
.B(n_1055),
.Y(n_1468)
);

INVx2_ASAP7_75t_L g1469 ( 
.A(n_1312),
.Y(n_1469)
);

AOI22xp5_ASAP7_75t_L g1470 ( 
.A1(n_1237),
.A2(n_1182),
.B1(n_1083),
.B2(n_1175),
.Y(n_1470)
);

INVx1_ASAP7_75t_L g1471 ( 
.A(n_1326),
.Y(n_1471)
);

NAND2xp5_ASAP7_75t_L g1472 ( 
.A(n_1333),
.B(n_1188),
.Y(n_1472)
);

AOI22xp33_ASAP7_75t_L g1473 ( 
.A1(n_1301),
.A2(n_1179),
.B1(n_1207),
.B2(n_1123),
.Y(n_1473)
);

NAND2xp5_ASAP7_75t_L g1474 ( 
.A(n_1310),
.B(n_1026),
.Y(n_1474)
);

NAND2xp5_ASAP7_75t_L g1475 ( 
.A(n_1275),
.B(n_1149),
.Y(n_1475)
);

INVx5_ASAP7_75t_L g1476 ( 
.A(n_1302),
.Y(n_1476)
);

NAND2xp5_ASAP7_75t_SL g1477 ( 
.A(n_1281),
.B(n_1010),
.Y(n_1477)
);

INVx3_ASAP7_75t_L g1478 ( 
.A(n_1270),
.Y(n_1478)
);

AOI21xp5_ASAP7_75t_L g1479 ( 
.A1(n_1393),
.A2(n_1197),
.B(n_1168),
.Y(n_1479)
);

NAND2xp5_ASAP7_75t_L g1480 ( 
.A(n_1388),
.B(n_1146),
.Y(n_1480)
);

AOI22xp33_ASAP7_75t_L g1481 ( 
.A1(n_1366),
.A2(n_1010),
.B1(n_1014),
.B2(n_1007),
.Y(n_1481)
);

NAND2x1p5_ASAP7_75t_L g1482 ( 
.A(n_1254),
.B(n_1167),
.Y(n_1482)
);

INVx3_ASAP7_75t_L g1483 ( 
.A(n_1270),
.Y(n_1483)
);

NAND2xp5_ASAP7_75t_SL g1484 ( 
.A(n_1324),
.B(n_1167),
.Y(n_1484)
);

BUFx3_ASAP7_75t_L g1485 ( 
.A(n_1317),
.Y(n_1485)
);

INVx2_ASAP7_75t_L g1486 ( 
.A(n_1424),
.Y(n_1486)
);

NAND2xp5_ASAP7_75t_L g1487 ( 
.A(n_1244),
.B(n_1168),
.Y(n_1487)
);

NOR2x1p5_ASAP7_75t_L g1488 ( 
.A(n_1304),
.B(n_1382),
.Y(n_1488)
);

AOI22xp33_ASAP7_75t_L g1489 ( 
.A1(n_1296),
.A2(n_1082),
.B1(n_1007),
.B2(n_1116),
.Y(n_1489)
);

INVx2_ASAP7_75t_SL g1490 ( 
.A(n_1278),
.Y(n_1490)
);

HB1xp67_ASAP7_75t_L g1491 ( 
.A(n_1305),
.Y(n_1491)
);

AND2x2_ASAP7_75t_SL g1492 ( 
.A(n_1268),
.B(n_1180),
.Y(n_1492)
);

NOR2x1_ASAP7_75t_R g1493 ( 
.A(n_1374),
.B(n_1167),
.Y(n_1493)
);

INVx2_ASAP7_75t_SL g1494 ( 
.A(n_1367),
.Y(n_1494)
);

AND2x2_ASAP7_75t_L g1495 ( 
.A(n_1345),
.B(n_1318),
.Y(n_1495)
);

AND2x2_ASAP7_75t_L g1496 ( 
.A(n_1345),
.B(n_1011),
.Y(n_1496)
);

NAND2xp5_ASAP7_75t_SL g1497 ( 
.A(n_1292),
.B(n_1180),
.Y(n_1497)
);

INVx1_ASAP7_75t_L g1498 ( 
.A(n_1336),
.Y(n_1498)
);

AND2x2_ASAP7_75t_L g1499 ( 
.A(n_1244),
.B(n_1012),
.Y(n_1499)
);

AOI22xp33_ASAP7_75t_L g1500 ( 
.A1(n_1358),
.A2(n_1082),
.B1(n_1117),
.B2(n_1018),
.Y(n_1500)
);

NOR2xp33_ASAP7_75t_L g1501 ( 
.A(n_1245),
.B(n_1017),
.Y(n_1501)
);

INVx2_ASAP7_75t_L g1502 ( 
.A(n_1355),
.Y(n_1502)
);

BUFx6f_ASAP7_75t_L g1503 ( 
.A(n_1344),
.Y(n_1503)
);

AND2x2_ASAP7_75t_L g1504 ( 
.A(n_1330),
.B(n_1347),
.Y(n_1504)
);

NAND2xp5_ASAP7_75t_L g1505 ( 
.A(n_1368),
.B(n_1019),
.Y(n_1505)
);

INVx1_ASAP7_75t_L g1506 ( 
.A(n_1369),
.Y(n_1506)
);

AOI22xp5_ASAP7_75t_L g1507 ( 
.A1(n_1265),
.A2(n_1022),
.B1(n_1023),
.B2(n_1021),
.Y(n_1507)
);

BUFx3_ASAP7_75t_L g1508 ( 
.A(n_1374),
.Y(n_1508)
);

AND2x4_ASAP7_75t_SL g1509 ( 
.A(n_1416),
.B(n_1030),
.Y(n_1509)
);

INVx2_ASAP7_75t_L g1510 ( 
.A(n_1403),
.Y(n_1510)
);

AND2x4_ASAP7_75t_L g1511 ( 
.A(n_1284),
.B(n_1377),
.Y(n_1511)
);

NAND2xp5_ASAP7_75t_SL g1512 ( 
.A(n_1292),
.B(n_1180),
.Y(n_1512)
);

AOI22xp5_ASAP7_75t_L g1513 ( 
.A1(n_1431),
.A2(n_1038),
.B1(n_1039),
.B2(n_1035),
.Y(n_1513)
);

INVx1_ASAP7_75t_L g1514 ( 
.A(n_1411),
.Y(n_1514)
);

AND2x4_ASAP7_75t_L g1515 ( 
.A(n_1353),
.B(n_1041),
.Y(n_1515)
);

INVx2_ASAP7_75t_SL g1516 ( 
.A(n_1416),
.Y(n_1516)
);

HB1xp67_ASAP7_75t_L g1517 ( 
.A(n_1394),
.Y(n_1517)
);

BUFx3_ASAP7_75t_L g1518 ( 
.A(n_1373),
.Y(n_1518)
);

NOR3xp33_ASAP7_75t_SL g1519 ( 
.A(n_1337),
.B(n_50),
.C(n_51),
.Y(n_1519)
);

BUFx6f_ASAP7_75t_L g1520 ( 
.A(n_1362),
.Y(n_1520)
);

NOR2x1p5_ASAP7_75t_L g1521 ( 
.A(n_1387),
.B(n_1177),
.Y(n_1521)
);

AOI22xp5_ASAP7_75t_L g1522 ( 
.A1(n_1260),
.A2(n_1046),
.B1(n_1048),
.B2(n_1045),
.Y(n_1522)
);

CKINVDCx5p33_ASAP7_75t_R g1523 ( 
.A(n_1298),
.Y(n_1523)
);

INVx1_ASAP7_75t_L g1524 ( 
.A(n_1412),
.Y(n_1524)
);

NOR2xp33_ASAP7_75t_SL g1525 ( 
.A(n_1332),
.B(n_1054),
.Y(n_1525)
);

BUFx2_ASAP7_75t_L g1526 ( 
.A(n_1390),
.Y(n_1526)
);

AND2x4_ASAP7_75t_L g1527 ( 
.A(n_1252),
.B(n_1061),
.Y(n_1527)
);

O2A1O1Ixp33_ASAP7_75t_L g1528 ( 
.A1(n_1398),
.A2(n_1379),
.B(n_1385),
.C(n_1415),
.Y(n_1528)
);

NAND2xp5_ASAP7_75t_L g1529 ( 
.A(n_1433),
.B(n_1062),
.Y(n_1529)
);

NAND2xp5_ASAP7_75t_L g1530 ( 
.A(n_1328),
.B(n_1064),
.Y(n_1530)
);

NOR2x1p5_ASAP7_75t_L g1531 ( 
.A(n_1261),
.B(n_50),
.Y(n_1531)
);

AND2x4_ASAP7_75t_L g1532 ( 
.A(n_1252),
.B(n_1206),
.Y(n_1532)
);

INVx2_ASAP7_75t_L g1533 ( 
.A(n_1283),
.Y(n_1533)
);

NAND2xp5_ASAP7_75t_SL g1534 ( 
.A(n_1299),
.B(n_1163),
.Y(n_1534)
);

NOR2xp33_ASAP7_75t_L g1535 ( 
.A(n_1267),
.B(n_1166),
.Y(n_1535)
);

AND2x2_ASAP7_75t_L g1536 ( 
.A(n_1260),
.B(n_51),
.Y(n_1536)
);

AOI22xp5_ASAP7_75t_L g1537 ( 
.A1(n_1421),
.A2(n_1190),
.B1(n_1124),
.B2(n_1173),
.Y(n_1537)
);

NAND2xp5_ASAP7_75t_SL g1538 ( 
.A(n_1299),
.B(n_1362),
.Y(n_1538)
);

BUFx6f_ASAP7_75t_L g1539 ( 
.A(n_1362),
.Y(n_1539)
);

NOR2xp33_ASAP7_75t_L g1540 ( 
.A(n_1251),
.B(n_1287),
.Y(n_1540)
);

INVx1_ASAP7_75t_L g1541 ( 
.A(n_1415),
.Y(n_1541)
);

INVx1_ASAP7_75t_L g1542 ( 
.A(n_1386),
.Y(n_1542)
);

BUFx3_ASAP7_75t_L g1543 ( 
.A(n_1373),
.Y(n_1543)
);

INVx2_ASAP7_75t_L g1544 ( 
.A(n_1286),
.Y(n_1544)
);

A2O1A1Ixp33_ASAP7_75t_L g1545 ( 
.A1(n_1406),
.A2(n_1183),
.B(n_1189),
.C(n_1170),
.Y(n_1545)
);

INVx1_ASAP7_75t_L g1546 ( 
.A(n_1289),
.Y(n_1546)
);

NAND2x1p5_ASAP7_75t_L g1547 ( 
.A(n_1390),
.B(n_52),
.Y(n_1547)
);

NAND2xp5_ASAP7_75t_SL g1548 ( 
.A(n_1404),
.B(n_53),
.Y(n_1548)
);

INVx1_ASAP7_75t_L g1549 ( 
.A(n_1423),
.Y(n_1549)
);

NAND2xp5_ASAP7_75t_SL g1550 ( 
.A(n_1404),
.B(n_1297),
.Y(n_1550)
);

CKINVDCx5p33_ASAP7_75t_R g1551 ( 
.A(n_1400),
.Y(n_1551)
);

BUFx2_ASAP7_75t_L g1552 ( 
.A(n_1349),
.Y(n_1552)
);

NAND2xp5_ASAP7_75t_SL g1553 ( 
.A(n_1404),
.B(n_53),
.Y(n_1553)
);

AOI22xp33_ASAP7_75t_L g1554 ( 
.A1(n_1414),
.A2(n_56),
.B1(n_54),
.B2(n_55),
.Y(n_1554)
);

INVx1_ASAP7_75t_L g1555 ( 
.A(n_1429),
.Y(n_1555)
);

AND2x2_ASAP7_75t_L g1556 ( 
.A(n_1315),
.B(n_54),
.Y(n_1556)
);

NOR2xp33_ASAP7_75t_L g1557 ( 
.A(n_1256),
.B(n_57),
.Y(n_1557)
);

NAND2xp5_ASAP7_75t_L g1558 ( 
.A(n_1272),
.B(n_58),
.Y(n_1558)
);

NAND2xp5_ASAP7_75t_SL g1559 ( 
.A(n_1407),
.B(n_1272),
.Y(n_1559)
);

INVx1_ASAP7_75t_L g1560 ( 
.A(n_1432),
.Y(n_1560)
);

NAND2xp5_ASAP7_75t_L g1561 ( 
.A(n_1242),
.B(n_59),
.Y(n_1561)
);

NAND2xp5_ASAP7_75t_L g1562 ( 
.A(n_1246),
.B(n_59),
.Y(n_1562)
);

INVx1_ASAP7_75t_L g1563 ( 
.A(n_1346),
.Y(n_1563)
);

AND2x4_ASAP7_75t_L g1564 ( 
.A(n_1331),
.B(n_61),
.Y(n_1564)
);

INVx2_ASAP7_75t_SL g1565 ( 
.A(n_1279),
.Y(n_1565)
);

NOR2xp33_ASAP7_75t_L g1566 ( 
.A(n_1250),
.B(n_61),
.Y(n_1566)
);

NAND2xp5_ASAP7_75t_SL g1567 ( 
.A(n_1259),
.B(n_62),
.Y(n_1567)
);

NAND3xp33_ASAP7_75t_SL g1568 ( 
.A(n_1401),
.B(n_65),
.C(n_66),
.Y(n_1568)
);

INVx1_ASAP7_75t_L g1569 ( 
.A(n_1364),
.Y(n_1569)
);

HB1xp67_ASAP7_75t_L g1570 ( 
.A(n_1379),
.Y(n_1570)
);

AOI22xp33_ASAP7_75t_L g1571 ( 
.A1(n_1381),
.A2(n_68),
.B1(n_65),
.B2(n_67),
.Y(n_1571)
);

NAND2xp5_ASAP7_75t_SL g1572 ( 
.A(n_1307),
.B(n_67),
.Y(n_1572)
);

HB1xp67_ASAP7_75t_L g1573 ( 
.A(n_1361),
.Y(n_1573)
);

NOR3xp33_ASAP7_75t_SL g1574 ( 
.A(n_1395),
.B(n_69),
.C(n_70),
.Y(n_1574)
);

NAND2xp5_ASAP7_75t_SL g1575 ( 
.A(n_1302),
.B(n_69),
.Y(n_1575)
);

BUFx2_ASAP7_75t_L g1576 ( 
.A(n_1430),
.Y(n_1576)
);

NAND3xp33_ASAP7_75t_SL g1577 ( 
.A(n_1401),
.B(n_71),
.C(n_72),
.Y(n_1577)
);

AND2x6_ASAP7_75t_L g1578 ( 
.A(n_1302),
.B(n_72),
.Y(n_1578)
);

AND2x4_ASAP7_75t_SL g1579 ( 
.A(n_1400),
.B(n_74),
.Y(n_1579)
);

NOR2xp67_ASAP7_75t_L g1580 ( 
.A(n_1397),
.B(n_74),
.Y(n_1580)
);

NAND2xp5_ASAP7_75t_SL g1581 ( 
.A(n_1269),
.B(n_75),
.Y(n_1581)
);

INVxp67_ASAP7_75t_L g1582 ( 
.A(n_1408),
.Y(n_1582)
);

BUFx4f_ASAP7_75t_SL g1583 ( 
.A(n_1402),
.Y(n_1583)
);

NAND2xp5_ASAP7_75t_L g1584 ( 
.A(n_1273),
.B(n_76),
.Y(n_1584)
);

AO21x1_ASAP7_75t_L g1585 ( 
.A1(n_1564),
.A2(n_1359),
.B(n_1405),
.Y(n_1585)
);

NAND2xp5_ASAP7_75t_L g1586 ( 
.A(n_1498),
.B(n_1425),
.Y(n_1586)
);

AOI21xp5_ASAP7_75t_L g1587 ( 
.A1(n_1458),
.A2(n_1354),
.B(n_1266),
.Y(n_1587)
);

OAI22xp5_ASAP7_75t_L g1588 ( 
.A1(n_1551),
.A2(n_1419),
.B1(n_1372),
.B2(n_1376),
.Y(n_1588)
);

INVx3_ASAP7_75t_SL g1589 ( 
.A(n_1437),
.Y(n_1589)
);

AOI21xp5_ASAP7_75t_L g1590 ( 
.A1(n_1479),
.A2(n_1266),
.B(n_1262),
.Y(n_1590)
);

OR2x2_ASAP7_75t_L g1591 ( 
.A(n_1445),
.B(n_1295),
.Y(n_1591)
);

AOI21xp5_ASAP7_75t_L g1592 ( 
.A1(n_1528),
.A2(n_1370),
.B(n_1262),
.Y(n_1592)
);

O2A1O1Ixp33_ASAP7_75t_L g1593 ( 
.A1(n_1582),
.A2(n_1420),
.B(n_1348),
.C(n_1325),
.Y(n_1593)
);

INVx2_ASAP7_75t_L g1594 ( 
.A(n_1435),
.Y(n_1594)
);

AOI21xp5_ASAP7_75t_L g1595 ( 
.A1(n_1541),
.A2(n_1370),
.B(n_1293),
.Y(n_1595)
);

INVx2_ASAP7_75t_L g1596 ( 
.A(n_1435),
.Y(n_1596)
);

AOI22x1_ASAP7_75t_L g1597 ( 
.A1(n_1521),
.A2(n_1410),
.B1(n_1417),
.B2(n_1413),
.Y(n_1597)
);

NOR2xp33_ASAP7_75t_L g1598 ( 
.A(n_1495),
.B(n_1316),
.Y(n_1598)
);

OAI21xp5_ASAP7_75t_L g1599 ( 
.A1(n_1487),
.A2(n_1340),
.B(n_1335),
.Y(n_1599)
);

AOI22x1_ASAP7_75t_L g1600 ( 
.A1(n_1570),
.A2(n_1249),
.B1(n_1276),
.B2(n_1241),
.Y(n_1600)
);

NAND3xp33_ASAP7_75t_L g1601 ( 
.A(n_1574),
.B(n_1418),
.C(n_1363),
.Y(n_1601)
);

NAND3xp33_ASAP7_75t_SL g1602 ( 
.A(n_1434),
.B(n_1422),
.C(n_1343),
.Y(n_1602)
);

CKINVDCx11_ASAP7_75t_R g1603 ( 
.A(n_1485),
.Y(n_1603)
);

AO32x2_ASAP7_75t_L g1604 ( 
.A1(n_1444),
.A2(n_1359),
.A3(n_1322),
.B1(n_1285),
.B2(n_1356),
.Y(n_1604)
);

AND2x2_ASAP7_75t_L g1605 ( 
.A(n_1488),
.B(n_1306),
.Y(n_1605)
);

NOR3xp33_ASAP7_75t_L g1606 ( 
.A(n_1568),
.B(n_1282),
.C(n_1280),
.Y(n_1606)
);

INVx4_ASAP7_75t_L g1607 ( 
.A(n_1441),
.Y(n_1607)
);

AOI22xp5_ASAP7_75t_L g1608 ( 
.A1(n_1579),
.A2(n_1264),
.B1(n_1342),
.B2(n_1339),
.Y(n_1608)
);

HB1xp67_ASAP7_75t_L g1609 ( 
.A(n_1447),
.Y(n_1609)
);

AOI21xp5_ASAP7_75t_L g1610 ( 
.A1(n_1559),
.A2(n_1440),
.B(n_1549),
.Y(n_1610)
);

OR2x2_ASAP7_75t_L g1611 ( 
.A(n_1465),
.B(n_1308),
.Y(n_1611)
);

HB1xp67_ASAP7_75t_L g1612 ( 
.A(n_1441),
.Y(n_1612)
);

INVx4_ASAP7_75t_L g1613 ( 
.A(n_1441),
.Y(n_1613)
);

INVx1_ASAP7_75t_L g1614 ( 
.A(n_1446),
.Y(n_1614)
);

AOI22x1_ASAP7_75t_L g1615 ( 
.A1(n_1531),
.A2(n_1391),
.B1(n_1384),
.B2(n_1365),
.Y(n_1615)
);

AOI21xp5_ASAP7_75t_L g1616 ( 
.A1(n_1555),
.A2(n_1392),
.B(n_1371),
.Y(n_1616)
);

BUFx6f_ASAP7_75t_L g1617 ( 
.A(n_1442),
.Y(n_1617)
);

NAND2xp5_ASAP7_75t_L g1618 ( 
.A(n_1439),
.B(n_1338),
.Y(n_1618)
);

AOI21x1_ASAP7_75t_L g1619 ( 
.A1(n_1538),
.A2(n_1360),
.B(n_1291),
.Y(n_1619)
);

AOI21xp5_ASAP7_75t_L g1620 ( 
.A1(n_1560),
.A2(n_1378),
.B(n_1357),
.Y(n_1620)
);

OAI22xp5_ASAP7_75t_L g1621 ( 
.A1(n_1508),
.A2(n_1311),
.B1(n_1314),
.B2(n_1313),
.Y(n_1621)
);

NAND2xp5_ASAP7_75t_SL g1622 ( 
.A(n_1476),
.B(n_1319),
.Y(n_1622)
);

AOI21xp5_ASAP7_75t_L g1623 ( 
.A1(n_1545),
.A2(n_1383),
.B(n_1327),
.Y(n_1623)
);

NOR2xp33_ASAP7_75t_L g1624 ( 
.A(n_1516),
.B(n_1351),
.Y(n_1624)
);

OAI22xp5_ASAP7_75t_L g1625 ( 
.A1(n_1466),
.A2(n_1468),
.B1(n_1451),
.B2(n_1547),
.Y(n_1625)
);

O2A1O1Ixp33_ASAP7_75t_L g1626 ( 
.A1(n_1453),
.A2(n_1352),
.B(n_1350),
.C(n_1323),
.Y(n_1626)
);

NAND2xp5_ASAP7_75t_SL g1627 ( 
.A(n_1476),
.B(n_1320),
.Y(n_1627)
);

BUFx8_ASAP7_75t_L g1628 ( 
.A(n_1455),
.Y(n_1628)
);

OAI22x1_ASAP7_75t_L g1629 ( 
.A1(n_1564),
.A2(n_79),
.B1(n_76),
.B2(n_78),
.Y(n_1629)
);

NAND2xp5_ASAP7_75t_SL g1630 ( 
.A(n_1476),
.B(n_1341),
.Y(n_1630)
);

AND2x4_ASAP7_75t_L g1631 ( 
.A(n_1436),
.B(n_1290),
.Y(n_1631)
);

NAND2xp5_ASAP7_75t_SL g1632 ( 
.A(n_1436),
.B(n_1426),
.Y(n_1632)
);

NOR2x1_ASAP7_75t_R g1633 ( 
.A(n_1452),
.B(n_1428),
.Y(n_1633)
);

OAI21xp5_ASAP7_75t_L g1634 ( 
.A1(n_1457),
.A2(n_78),
.B(n_80),
.Y(n_1634)
);

INVx3_ASAP7_75t_L g1635 ( 
.A(n_1482),
.Y(n_1635)
);

INVxp67_ASAP7_75t_L g1636 ( 
.A(n_1493),
.Y(n_1636)
);

INVx1_ASAP7_75t_L g1637 ( 
.A(n_1449),
.Y(n_1637)
);

HB1xp67_ASAP7_75t_L g1638 ( 
.A(n_1546),
.Y(n_1638)
);

INVx1_ASAP7_75t_L g1639 ( 
.A(n_1450),
.Y(n_1639)
);

NAND2xp5_ASAP7_75t_L g1640 ( 
.A(n_1438),
.B(n_81),
.Y(n_1640)
);

INVx5_ASAP7_75t_L g1641 ( 
.A(n_1578),
.Y(n_1641)
);

NOR2xp33_ASAP7_75t_L g1642 ( 
.A(n_1474),
.B(n_81),
.Y(n_1642)
);

NAND2x1p5_ASAP7_75t_L g1643 ( 
.A(n_1518),
.B(n_82),
.Y(n_1643)
);

OAI22xp5_ASAP7_75t_SL g1644 ( 
.A1(n_1464),
.A2(n_84),
.B1(n_82),
.B2(n_83),
.Y(n_1644)
);

HB1xp67_ASAP7_75t_L g1645 ( 
.A(n_1546),
.Y(n_1645)
);

NAND2xp5_ASAP7_75t_SL g1646 ( 
.A(n_1511),
.B(n_83),
.Y(n_1646)
);

BUFx3_ASAP7_75t_L g1647 ( 
.A(n_1443),
.Y(n_1647)
);

NAND2xp5_ASAP7_75t_L g1648 ( 
.A(n_1460),
.B(n_85),
.Y(n_1648)
);

AOI22xp5_ASAP7_75t_L g1649 ( 
.A1(n_1536),
.A2(n_89),
.B1(n_86),
.B2(n_87),
.Y(n_1649)
);

INVx3_ASAP7_75t_L g1650 ( 
.A(n_1543),
.Y(n_1650)
);

OAI22x1_ASAP7_75t_L g1651 ( 
.A1(n_1484),
.A2(n_90),
.B1(n_87),
.B2(n_89),
.Y(n_1651)
);

INVx2_ASAP7_75t_L g1652 ( 
.A(n_1461),
.Y(n_1652)
);

NAND2xp5_ASAP7_75t_SL g1653 ( 
.A(n_1511),
.B(n_90),
.Y(n_1653)
);

OR2x6_ASAP7_75t_L g1654 ( 
.A(n_1490),
.B(n_91),
.Y(n_1654)
);

INVx4_ASAP7_75t_L g1655 ( 
.A(n_1578),
.Y(n_1655)
);

NOR2xp33_ASAP7_75t_L g1656 ( 
.A(n_1468),
.B(n_91),
.Y(n_1656)
);

INVx1_ASAP7_75t_L g1657 ( 
.A(n_1467),
.Y(n_1657)
);

AND2x2_ASAP7_75t_L g1658 ( 
.A(n_1504),
.B(n_92),
.Y(n_1658)
);

NAND2xp5_ASAP7_75t_L g1659 ( 
.A(n_1462),
.B(n_92),
.Y(n_1659)
);

AOI22xp33_ASAP7_75t_L g1660 ( 
.A1(n_1577),
.A2(n_95),
.B1(n_93),
.B2(n_94),
.Y(n_1660)
);

NOR2xp33_ASAP7_75t_L g1661 ( 
.A(n_1540),
.B(n_93),
.Y(n_1661)
);

A2O1A1Ixp33_ASAP7_75t_L g1662 ( 
.A1(n_1566),
.A2(n_97),
.B(n_94),
.C(n_96),
.Y(n_1662)
);

OAI21xp33_ASAP7_75t_L g1663 ( 
.A1(n_1470),
.A2(n_96),
.B(n_97),
.Y(n_1663)
);

INVx2_ASAP7_75t_SL g1664 ( 
.A(n_1517),
.Y(n_1664)
);

INVx1_ASAP7_75t_L g1665 ( 
.A(n_1469),
.Y(n_1665)
);

AND2x2_ASAP7_75t_L g1666 ( 
.A(n_1471),
.B(n_98),
.Y(n_1666)
);

NAND2xp5_ASAP7_75t_L g1667 ( 
.A(n_1506),
.B(n_98),
.Y(n_1667)
);

NAND2xp5_ASAP7_75t_L g1668 ( 
.A(n_1514),
.B(n_101),
.Y(n_1668)
);

NAND2xp5_ASAP7_75t_L g1669 ( 
.A(n_1524),
.B(n_101),
.Y(n_1669)
);

NOR2xp33_ASAP7_75t_L g1670 ( 
.A(n_1480),
.B(n_102),
.Y(n_1670)
);

INVx3_ASAP7_75t_L g1671 ( 
.A(n_1583),
.Y(n_1671)
);

BUFx8_ASAP7_75t_L g1672 ( 
.A(n_1578),
.Y(n_1672)
);

AOI21xp5_ASAP7_75t_L g1673 ( 
.A1(n_1542),
.A2(n_128),
.B(n_123),
.Y(n_1673)
);

AND2x2_ASAP7_75t_L g1674 ( 
.A(n_1502),
.B(n_104),
.Y(n_1674)
);

A2O1A1Ixp33_ASAP7_75t_SL g1675 ( 
.A1(n_1557),
.A2(n_107),
.B(n_104),
.C(n_106),
.Y(n_1675)
);

NAND2xp5_ASAP7_75t_L g1676 ( 
.A(n_1448),
.B(n_106),
.Y(n_1676)
);

NAND2xp5_ASAP7_75t_L g1677 ( 
.A(n_1598),
.B(n_1510),
.Y(n_1677)
);

INVx1_ASAP7_75t_SL g1678 ( 
.A(n_1589),
.Y(n_1678)
);

AOI21xp5_ASAP7_75t_L g1679 ( 
.A1(n_1592),
.A2(n_1512),
.B(n_1497),
.Y(n_1679)
);

AOI21xp5_ASAP7_75t_L g1680 ( 
.A1(n_1587),
.A2(n_1534),
.B(n_1477),
.Y(n_1680)
);

BUFx2_ASAP7_75t_L g1681 ( 
.A(n_1613),
.Y(n_1681)
);

AOI221xp5_ASAP7_75t_SL g1682 ( 
.A1(n_1629),
.A2(n_1554),
.B1(n_1581),
.B2(n_1567),
.C(n_1558),
.Y(n_1682)
);

INVx2_ASAP7_75t_L g1683 ( 
.A(n_1652),
.Y(n_1683)
);

BUFx3_ASAP7_75t_L g1684 ( 
.A(n_1628),
.Y(n_1684)
);

NOR4xp25_ASAP7_75t_L g1685 ( 
.A(n_1634),
.B(n_1572),
.C(n_1496),
.D(n_1575),
.Y(n_1685)
);

OAI21x1_ASAP7_75t_L g1686 ( 
.A1(n_1600),
.A2(n_1597),
.B(n_1590),
.Y(n_1686)
);

AOI21xp5_ASAP7_75t_SL g1687 ( 
.A1(n_1655),
.A2(n_1578),
.B(n_1456),
.Y(n_1687)
);

HB1xp67_ASAP7_75t_L g1688 ( 
.A(n_1609),
.Y(n_1688)
);

AOI21xp5_ASAP7_75t_L g1689 ( 
.A1(n_1595),
.A2(n_1454),
.B(n_1442),
.Y(n_1689)
);

BUFx6f_ASAP7_75t_L g1690 ( 
.A(n_1617),
.Y(n_1690)
);

INVx1_ASAP7_75t_L g1691 ( 
.A(n_1614),
.Y(n_1691)
);

NAND2xp5_ASAP7_75t_L g1692 ( 
.A(n_1594),
.B(n_1596),
.Y(n_1692)
);

NAND2xp5_ASAP7_75t_L g1693 ( 
.A(n_1586),
.B(n_1499),
.Y(n_1693)
);

NOR2xp33_ASAP7_75t_SL g1694 ( 
.A(n_1672),
.B(n_1523),
.Y(n_1694)
);

NAND2x1p5_ASAP7_75t_L g1695 ( 
.A(n_1613),
.B(n_1459),
.Y(n_1695)
);

NAND3xp33_ASAP7_75t_L g1696 ( 
.A(n_1606),
.B(n_1519),
.C(n_1571),
.Y(n_1696)
);

INVx1_ASAP7_75t_L g1697 ( 
.A(n_1637),
.Y(n_1697)
);

NAND2xp5_ASAP7_75t_L g1698 ( 
.A(n_1639),
.B(n_1472),
.Y(n_1698)
);

NAND2xp5_ASAP7_75t_L g1699 ( 
.A(n_1657),
.B(n_1556),
.Y(n_1699)
);

NOR2xp33_ASAP7_75t_L g1700 ( 
.A(n_1605),
.B(n_1565),
.Y(n_1700)
);

NOR2xp67_ASAP7_75t_L g1701 ( 
.A(n_1655),
.B(n_1494),
.Y(n_1701)
);

NAND3x1_ASAP7_75t_L g1702 ( 
.A(n_1656),
.B(n_1463),
.C(n_1584),
.Y(n_1702)
);

AOI21xp5_ASAP7_75t_L g1703 ( 
.A1(n_1610),
.A2(n_1454),
.B(n_1442),
.Y(n_1703)
);

INVx1_ASAP7_75t_L g1704 ( 
.A(n_1665),
.Y(n_1704)
);

INVx1_ASAP7_75t_L g1705 ( 
.A(n_1638),
.Y(n_1705)
);

OAI21x1_ASAP7_75t_L g1706 ( 
.A1(n_1623),
.A2(n_1550),
.B(n_1548),
.Y(n_1706)
);

INVx1_ASAP7_75t_L g1707 ( 
.A(n_1645),
.Y(n_1707)
);

INVx1_ASAP7_75t_L g1708 ( 
.A(n_1611),
.Y(n_1708)
);

OAI21x1_ASAP7_75t_L g1709 ( 
.A1(n_1619),
.A2(n_1553),
.B(n_1513),
.Y(n_1709)
);

OA21x2_ASAP7_75t_L g1710 ( 
.A1(n_1585),
.A2(n_1500),
.B(n_1489),
.Y(n_1710)
);

AND2x2_ASAP7_75t_L g1711 ( 
.A(n_1658),
.B(n_1491),
.Y(n_1711)
);

BUFx12f_ASAP7_75t_L g1712 ( 
.A(n_1603),
.Y(n_1712)
);

AOI21x1_ASAP7_75t_L g1713 ( 
.A1(n_1625),
.A2(n_1580),
.B(n_1573),
.Y(n_1713)
);

INVx1_ASAP7_75t_L g1714 ( 
.A(n_1666),
.Y(n_1714)
);

AOI21xp5_ASAP7_75t_L g1715 ( 
.A1(n_1599),
.A2(n_1503),
.B(n_1454),
.Y(n_1715)
);

INVx1_ASAP7_75t_L g1716 ( 
.A(n_1674),
.Y(n_1716)
);

AO31x2_ASAP7_75t_L g1717 ( 
.A1(n_1651),
.A2(n_1569),
.A3(n_1563),
.B(n_1561),
.Y(n_1717)
);

OAI21x1_ASAP7_75t_L g1718 ( 
.A1(n_1616),
.A2(n_1620),
.B(n_1673),
.Y(n_1718)
);

INVx2_ASAP7_75t_SL g1719 ( 
.A(n_1628),
.Y(n_1719)
);

AOI21xp5_ASAP7_75t_L g1720 ( 
.A1(n_1588),
.A2(n_1520),
.B(n_1503),
.Y(n_1720)
);

AND2x4_ASAP7_75t_L g1721 ( 
.A(n_1641),
.B(n_1552),
.Y(n_1721)
);

BUFx12f_ASAP7_75t_L g1722 ( 
.A(n_1672),
.Y(n_1722)
);

NAND2xp5_ASAP7_75t_SL g1723 ( 
.A(n_1641),
.B(n_1492),
.Y(n_1723)
);

AOI22xp5_ASAP7_75t_L g1724 ( 
.A1(n_1602),
.A2(n_1562),
.B1(n_1475),
.B2(n_1535),
.Y(n_1724)
);

NAND2xp5_ASAP7_75t_L g1725 ( 
.A(n_1661),
.B(n_1486),
.Y(n_1725)
);

AOI21xp5_ASAP7_75t_L g1726 ( 
.A1(n_1618),
.A2(n_1520),
.B(n_1503),
.Y(n_1726)
);

OAI22xp5_ASAP7_75t_L g1727 ( 
.A1(n_1724),
.A2(n_1641),
.B1(n_1649),
.B2(n_1693),
.Y(n_1727)
);

OAI22xp33_ASAP7_75t_L g1728 ( 
.A1(n_1684),
.A2(n_1654),
.B1(n_1608),
.B2(n_1643),
.Y(n_1728)
);

INVx1_ASAP7_75t_L g1729 ( 
.A(n_1691),
.Y(n_1729)
);

OAI21x1_ASAP7_75t_L g1730 ( 
.A1(n_1686),
.A2(n_1615),
.B(n_1622),
.Y(n_1730)
);

INVx1_ASAP7_75t_L g1731 ( 
.A(n_1697),
.Y(n_1731)
);

INVxp67_ASAP7_75t_L g1732 ( 
.A(n_1681),
.Y(n_1732)
);

INVx3_ASAP7_75t_L g1733 ( 
.A(n_1721),
.Y(n_1733)
);

AO21x2_ASAP7_75t_L g1734 ( 
.A1(n_1679),
.A2(n_1663),
.B(n_1675),
.Y(n_1734)
);

INVx1_ASAP7_75t_L g1735 ( 
.A(n_1704),
.Y(n_1735)
);

OAI22xp33_ASAP7_75t_L g1736 ( 
.A1(n_1678),
.A2(n_1654),
.B1(n_1612),
.B2(n_1653),
.Y(n_1736)
);

AO31x2_ASAP7_75t_L g1737 ( 
.A1(n_1680),
.A2(n_1662),
.A3(n_1621),
.B(n_1670),
.Y(n_1737)
);

AOI22xp33_ASAP7_75t_L g1738 ( 
.A1(n_1696),
.A2(n_1644),
.B1(n_1642),
.B2(n_1601),
.Y(n_1738)
);

NAND2xp5_ASAP7_75t_L g1739 ( 
.A(n_1698),
.B(n_1640),
.Y(n_1739)
);

INVx1_ASAP7_75t_L g1740 ( 
.A(n_1705),
.Y(n_1740)
);

INVx1_ASAP7_75t_L g1741 ( 
.A(n_1707),
.Y(n_1741)
);

OAI21xp5_ASAP7_75t_L g1742 ( 
.A1(n_1724),
.A2(n_1696),
.B(n_1685),
.Y(n_1742)
);

OAI21x1_ASAP7_75t_L g1743 ( 
.A1(n_1689),
.A2(n_1630),
.B(n_1627),
.Y(n_1743)
);

NAND2xp5_ASAP7_75t_L g1744 ( 
.A(n_1692),
.B(n_1716),
.Y(n_1744)
);

OAI21x1_ASAP7_75t_L g1745 ( 
.A1(n_1703),
.A2(n_1626),
.B(n_1632),
.Y(n_1745)
);

NAND2x1p5_ASAP7_75t_L g1746 ( 
.A(n_1719),
.B(n_1607),
.Y(n_1746)
);

AND2x2_ASAP7_75t_L g1747 ( 
.A(n_1708),
.B(n_1664),
.Y(n_1747)
);

NAND2x1p5_ASAP7_75t_L g1748 ( 
.A(n_1721),
.B(n_1650),
.Y(n_1748)
);

AOI22xp33_ASAP7_75t_L g1749 ( 
.A1(n_1711),
.A2(n_1646),
.B1(n_1660),
.B2(n_1676),
.Y(n_1749)
);

AND2x2_ASAP7_75t_L g1750 ( 
.A(n_1677),
.B(n_1591),
.Y(n_1750)
);

INVx1_ASAP7_75t_L g1751 ( 
.A(n_1683),
.Y(n_1751)
);

NAND2xp5_ASAP7_75t_L g1752 ( 
.A(n_1714),
.B(n_1685),
.Y(n_1752)
);

AO21x2_ASAP7_75t_L g1753 ( 
.A1(n_1713),
.A2(n_1659),
.B(n_1648),
.Y(n_1753)
);

OR2x2_ASAP7_75t_L g1754 ( 
.A(n_1688),
.B(n_1647),
.Y(n_1754)
);

AO21x2_ASAP7_75t_L g1755 ( 
.A1(n_1720),
.A2(n_1668),
.B(n_1667),
.Y(n_1755)
);

OAI22xp5_ASAP7_75t_L g1756 ( 
.A1(n_1702),
.A2(n_1669),
.B1(n_1636),
.B2(n_1481),
.Y(n_1756)
);

A2O1A1Ixp33_ASAP7_75t_L g1757 ( 
.A1(n_1682),
.A2(n_1593),
.B(n_1635),
.C(n_1631),
.Y(n_1757)
);

BUFx2_ASAP7_75t_L g1758 ( 
.A(n_1695),
.Y(n_1758)
);

AOI22xp5_ASAP7_75t_L g1759 ( 
.A1(n_1725),
.A2(n_1624),
.B1(n_1501),
.B2(n_1671),
.Y(n_1759)
);

INVx1_ASAP7_75t_L g1760 ( 
.A(n_1699),
.Y(n_1760)
);

OA21x2_ASAP7_75t_L g1761 ( 
.A1(n_1709),
.A2(n_1530),
.B(n_1522),
.Y(n_1761)
);

AND2x4_ASAP7_75t_L g1762 ( 
.A(n_1733),
.B(n_1701),
.Y(n_1762)
);

OAI22xp5_ASAP7_75t_L g1763 ( 
.A1(n_1727),
.A2(n_1687),
.B1(n_1723),
.B2(n_1701),
.Y(n_1763)
);

AND2x2_ASAP7_75t_L g1764 ( 
.A(n_1750),
.B(n_1700),
.Y(n_1764)
);

O2A1O1Ixp33_ASAP7_75t_L g1765 ( 
.A1(n_1728),
.A2(n_1756),
.B(n_1736),
.C(n_1757),
.Y(n_1765)
);

INVxp67_ASAP7_75t_L g1766 ( 
.A(n_1754),
.Y(n_1766)
);

AOI21xp5_ASAP7_75t_L g1767 ( 
.A1(n_1742),
.A2(n_1715),
.B(n_1726),
.Y(n_1767)
);

AOI21xp5_ASAP7_75t_L g1768 ( 
.A1(n_1742),
.A2(n_1710),
.B(n_1718),
.Y(n_1768)
);

BUFx3_ASAP7_75t_L g1769 ( 
.A(n_1746),
.Y(n_1769)
);

O2A1O1Ixp5_ASAP7_75t_L g1770 ( 
.A1(n_1756),
.A2(n_1631),
.B(n_1515),
.C(n_1478),
.Y(n_1770)
);

INVxp67_ASAP7_75t_L g1771 ( 
.A(n_1732),
.Y(n_1771)
);

O2A1O1Ixp5_ASAP7_75t_L g1772 ( 
.A1(n_1752),
.A2(n_1515),
.B(n_1478),
.C(n_1483),
.Y(n_1772)
);

OA21x2_ASAP7_75t_L g1773 ( 
.A1(n_1730),
.A2(n_1706),
.B(n_1682),
.Y(n_1773)
);

O2A1O1Ixp5_ASAP7_75t_L g1774 ( 
.A1(n_1752),
.A2(n_1727),
.B(n_1733),
.C(n_1739),
.Y(n_1774)
);

AOI211xp5_ASAP7_75t_L g1775 ( 
.A1(n_1732),
.A2(n_1633),
.B(n_1694),
.C(n_1526),
.Y(n_1775)
);

AOI21xp5_ASAP7_75t_SL g1776 ( 
.A1(n_1748),
.A2(n_1710),
.B(n_1690),
.Y(n_1776)
);

OAI22xp5_ASAP7_75t_L g1777 ( 
.A1(n_1738),
.A2(n_1722),
.B1(n_1690),
.B2(n_1712),
.Y(n_1777)
);

AOI21x1_ASAP7_75t_SL g1778 ( 
.A1(n_1739),
.A2(n_1527),
.B(n_1532),
.Y(n_1778)
);

OR2x2_ASAP7_75t_L g1779 ( 
.A(n_1740),
.B(n_1717),
.Y(n_1779)
);

INVx2_ASAP7_75t_L g1780 ( 
.A(n_1751),
.Y(n_1780)
);

INVx1_ASAP7_75t_L g1781 ( 
.A(n_1729),
.Y(n_1781)
);

NAND2xp5_ASAP7_75t_L g1782 ( 
.A(n_1760),
.B(n_1717),
.Y(n_1782)
);

A2O1A1Ixp33_ASAP7_75t_L g1783 ( 
.A1(n_1758),
.A2(n_1759),
.B(n_1749),
.C(n_1741),
.Y(n_1783)
);

OR2x2_ASAP7_75t_L g1784 ( 
.A(n_1744),
.B(n_1717),
.Y(n_1784)
);

AND2x4_ASAP7_75t_L g1785 ( 
.A(n_1731),
.B(n_1690),
.Y(n_1785)
);

INVx1_ASAP7_75t_L g1786 ( 
.A(n_1735),
.Y(n_1786)
);

OAI22xp5_ASAP7_75t_L g1787 ( 
.A1(n_1744),
.A2(n_1544),
.B1(n_1533),
.B2(n_1617),
.Y(n_1787)
);

INVx3_ASAP7_75t_L g1788 ( 
.A(n_1748),
.Y(n_1788)
);

OAI22xp5_ASAP7_75t_L g1789 ( 
.A1(n_1746),
.A2(n_1473),
.B1(n_1509),
.B2(n_1617),
.Y(n_1789)
);

INVx2_ASAP7_75t_L g1790 ( 
.A(n_1747),
.Y(n_1790)
);

AND2x4_ASAP7_75t_L g1791 ( 
.A(n_1755),
.B(n_1459),
.Y(n_1791)
);

INVx2_ASAP7_75t_L g1792 ( 
.A(n_1780),
.Y(n_1792)
);

AOI22xp33_ASAP7_75t_L g1793 ( 
.A1(n_1777),
.A2(n_1755),
.B1(n_1753),
.B2(n_1734),
.Y(n_1793)
);

AND2x2_ASAP7_75t_L g1794 ( 
.A(n_1784),
.B(n_1761),
.Y(n_1794)
);

BUFx3_ASAP7_75t_L g1795 ( 
.A(n_1769),
.Y(n_1795)
);

OR2x2_ASAP7_75t_L g1796 ( 
.A(n_1782),
.B(n_1753),
.Y(n_1796)
);

OA21x2_ASAP7_75t_L g1797 ( 
.A1(n_1768),
.A2(n_1745),
.B(n_1743),
.Y(n_1797)
);

INVx2_ASAP7_75t_R g1798 ( 
.A(n_1778),
.Y(n_1798)
);

BUFx2_ASAP7_75t_L g1799 ( 
.A(n_1762),
.Y(n_1799)
);

INVx1_ASAP7_75t_L g1800 ( 
.A(n_1781),
.Y(n_1800)
);

NAND3xp33_ASAP7_75t_L g1801 ( 
.A(n_1775),
.B(n_1761),
.C(n_1525),
.Y(n_1801)
);

INVx3_ASAP7_75t_L g1802 ( 
.A(n_1791),
.Y(n_1802)
);

AND2x2_ASAP7_75t_L g1803 ( 
.A(n_1786),
.B(n_1737),
.Y(n_1803)
);

INVx1_ASAP7_75t_L g1804 ( 
.A(n_1779),
.Y(n_1804)
);

INVx1_ASAP7_75t_L g1805 ( 
.A(n_1791),
.Y(n_1805)
);

NAND2xp5_ASAP7_75t_L g1806 ( 
.A(n_1771),
.B(n_1737),
.Y(n_1806)
);

OAI21x1_ASAP7_75t_L g1807 ( 
.A1(n_1767),
.A2(n_1483),
.B(n_1505),
.Y(n_1807)
);

AND2x2_ASAP7_75t_L g1808 ( 
.A(n_1790),
.B(n_1737),
.Y(n_1808)
);

OR2x6_ASAP7_75t_L g1809 ( 
.A(n_1763),
.B(n_1776),
.Y(n_1809)
);

AO21x2_ASAP7_75t_L g1810 ( 
.A1(n_1787),
.A2(n_1734),
.B(n_1507),
.Y(n_1810)
);

OAI21xp5_ASAP7_75t_L g1811 ( 
.A1(n_1770),
.A2(n_1529),
.B(n_1576),
.Y(n_1811)
);

OR2x2_ASAP7_75t_L g1812 ( 
.A(n_1766),
.B(n_108),
.Y(n_1812)
);

INVx2_ASAP7_75t_L g1813 ( 
.A(n_1773),
.Y(n_1813)
);

AO21x2_ASAP7_75t_L g1814 ( 
.A1(n_1787),
.A2(n_1537),
.B(n_1604),
.Y(n_1814)
);

AND2x2_ASAP7_75t_L g1815 ( 
.A(n_1785),
.B(n_1604),
.Y(n_1815)
);

AND2x2_ASAP7_75t_L g1816 ( 
.A(n_1808),
.B(n_1794),
.Y(n_1816)
);

NAND2xp5_ASAP7_75t_L g1817 ( 
.A(n_1808),
.B(n_1783),
.Y(n_1817)
);

INVx2_ASAP7_75t_L g1818 ( 
.A(n_1792),
.Y(n_1818)
);

AND2x2_ASAP7_75t_L g1819 ( 
.A(n_1794),
.B(n_1773),
.Y(n_1819)
);

A2O1A1Ixp33_ASAP7_75t_L g1820 ( 
.A1(n_1795),
.A2(n_1775),
.B(n_1765),
.C(n_1777),
.Y(n_1820)
);

HB1xp67_ASAP7_75t_L g1821 ( 
.A(n_1792),
.Y(n_1821)
);

INVx3_ASAP7_75t_L g1822 ( 
.A(n_1802),
.Y(n_1822)
);

INVx1_ASAP7_75t_L g1823 ( 
.A(n_1792),
.Y(n_1823)
);

INVx1_ASAP7_75t_L g1824 ( 
.A(n_1804),
.Y(n_1824)
);

INVx2_ASAP7_75t_L g1825 ( 
.A(n_1800),
.Y(n_1825)
);

AND2x2_ASAP7_75t_L g1826 ( 
.A(n_1805),
.B(n_1785),
.Y(n_1826)
);

BUFx3_ASAP7_75t_L g1827 ( 
.A(n_1795),
.Y(n_1827)
);

AND2x2_ASAP7_75t_L g1828 ( 
.A(n_1805),
.B(n_1764),
.Y(n_1828)
);

INVx2_ASAP7_75t_L g1829 ( 
.A(n_1800),
.Y(n_1829)
);

INVx2_ASAP7_75t_SL g1830 ( 
.A(n_1795),
.Y(n_1830)
);

AND2x4_ASAP7_75t_L g1831 ( 
.A(n_1802),
.B(n_1762),
.Y(n_1831)
);

AND2x2_ASAP7_75t_L g1832 ( 
.A(n_1815),
.B(n_1774),
.Y(n_1832)
);

BUFx3_ASAP7_75t_L g1833 ( 
.A(n_1799),
.Y(n_1833)
);

AND2x2_ASAP7_75t_L g1834 ( 
.A(n_1815),
.B(n_1772),
.Y(n_1834)
);

INVx2_ASAP7_75t_L g1835 ( 
.A(n_1804),
.Y(n_1835)
);

BUFx24_ASAP7_75t_SL g1836 ( 
.A(n_1820),
.Y(n_1836)
);

NAND4xp75_ASAP7_75t_L g1837 ( 
.A(n_1830),
.B(n_1806),
.C(n_1811),
.D(n_1803),
.Y(n_1837)
);

AND2x4_ASAP7_75t_L g1838 ( 
.A(n_1827),
.B(n_1802),
.Y(n_1838)
);

AND2x2_ASAP7_75t_L g1839 ( 
.A(n_1816),
.B(n_1799),
.Y(n_1839)
);

OAI22xp5_ASAP7_75t_L g1840 ( 
.A1(n_1827),
.A2(n_1801),
.B1(n_1809),
.B2(n_1812),
.Y(n_1840)
);

AND2x2_ASAP7_75t_L g1841 ( 
.A(n_1816),
.B(n_1802),
.Y(n_1841)
);

BUFx3_ASAP7_75t_L g1842 ( 
.A(n_1827),
.Y(n_1842)
);

INVx1_ASAP7_75t_L g1843 ( 
.A(n_1824),
.Y(n_1843)
);

AND2x2_ASAP7_75t_L g1844 ( 
.A(n_1828),
.B(n_1803),
.Y(n_1844)
);

OAI22xp5_ASAP7_75t_L g1845 ( 
.A1(n_1830),
.A2(n_1801),
.B1(n_1809),
.B2(n_1812),
.Y(n_1845)
);

AOI22xp33_ASAP7_75t_L g1846 ( 
.A1(n_1832),
.A2(n_1809),
.B1(n_1798),
.B2(n_1806),
.Y(n_1846)
);

AOI221xp5_ASAP7_75t_L g1847 ( 
.A1(n_1832),
.A2(n_1793),
.B1(n_1763),
.B2(n_1796),
.C(n_1789),
.Y(n_1847)
);

OR2x2_ASAP7_75t_L g1848 ( 
.A(n_1835),
.B(n_1796),
.Y(n_1848)
);

AOI22xp33_ASAP7_75t_SL g1849 ( 
.A1(n_1833),
.A2(n_1809),
.B1(n_1788),
.B2(n_1810),
.Y(n_1849)
);

NOR2x2_ASAP7_75t_L g1850 ( 
.A(n_1835),
.B(n_1809),
.Y(n_1850)
);

AOI22xp33_ASAP7_75t_SL g1851 ( 
.A1(n_1833),
.A2(n_1788),
.B1(n_1810),
.B2(n_1811),
.Y(n_1851)
);

BUFx3_ASAP7_75t_L g1852 ( 
.A(n_1833),
.Y(n_1852)
);

NOR3xp33_ASAP7_75t_L g1853 ( 
.A(n_1817),
.B(n_1807),
.C(n_1813),
.Y(n_1853)
);

INVx4_ASAP7_75t_SL g1854 ( 
.A(n_1831),
.Y(n_1854)
);

OAI221xp5_ASAP7_75t_L g1855 ( 
.A1(n_1822),
.A2(n_1813),
.B1(n_1797),
.B2(n_1798),
.C(n_1810),
.Y(n_1855)
);

BUFx2_ASAP7_75t_L g1856 ( 
.A(n_1831),
.Y(n_1856)
);

INVx2_ASAP7_75t_L g1857 ( 
.A(n_1852),
.Y(n_1857)
);

AOI21x1_ASAP7_75t_L g1858 ( 
.A1(n_1845),
.A2(n_1831),
.B(n_1821),
.Y(n_1858)
);

INVx2_ASAP7_75t_L g1859 ( 
.A(n_1848),
.Y(n_1859)
);

INVx5_ASAP7_75t_L g1860 ( 
.A(n_1842),
.Y(n_1860)
);

NAND2xp5_ASAP7_75t_L g1861 ( 
.A(n_1847),
.B(n_1819),
.Y(n_1861)
);

INVx1_ASAP7_75t_L g1862 ( 
.A(n_1843),
.Y(n_1862)
);

NAND2xp5_ASAP7_75t_L g1863 ( 
.A(n_1844),
.B(n_1819),
.Y(n_1863)
);

INVx2_ASAP7_75t_L g1864 ( 
.A(n_1841),
.Y(n_1864)
);

INVx2_ASAP7_75t_L g1865 ( 
.A(n_1860),
.Y(n_1865)
);

NAND2xp5_ASAP7_75t_L g1866 ( 
.A(n_1861),
.B(n_1853),
.Y(n_1866)
);

AND2x4_ASAP7_75t_L g1867 ( 
.A(n_1860),
.B(n_1854),
.Y(n_1867)
);

INVx1_ASAP7_75t_L g1868 ( 
.A(n_1862),
.Y(n_1868)
);

AND2x2_ASAP7_75t_L g1869 ( 
.A(n_1865),
.B(n_1858),
.Y(n_1869)
);

INVx1_ASAP7_75t_L g1870 ( 
.A(n_1868),
.Y(n_1870)
);

INVx1_ASAP7_75t_SL g1871 ( 
.A(n_1870),
.Y(n_1871)
);

AOI222xp33_ASAP7_75t_L g1872 ( 
.A1(n_1869),
.A2(n_1866),
.B1(n_1867),
.B2(n_1840),
.C1(n_1845),
.C2(n_1836),
.Y(n_1872)
);

INVx1_ASAP7_75t_L g1873 ( 
.A(n_1869),
.Y(n_1873)
);

NAND3xp33_ASAP7_75t_L g1874 ( 
.A(n_1869),
.B(n_1851),
.C(n_1849),
.Y(n_1874)
);

OAI21xp33_ASAP7_75t_SL g1875 ( 
.A1(n_1873),
.A2(n_1863),
.B(n_1857),
.Y(n_1875)
);

OR2x2_ASAP7_75t_L g1876 ( 
.A(n_1871),
.B(n_1859),
.Y(n_1876)
);

AOI322xp5_ASAP7_75t_L g1877 ( 
.A1(n_1872),
.A2(n_1867),
.A3(n_1846),
.B1(n_1856),
.B2(n_1828),
.C1(n_1839),
.C2(n_1864),
.Y(n_1877)
);

OR2x2_ASAP7_75t_L g1878 ( 
.A(n_1874),
.B(n_1824),
.Y(n_1878)
);

NOR2xp33_ASAP7_75t_L g1879 ( 
.A(n_1873),
.B(n_1860),
.Y(n_1879)
);

AOI21xp5_ASAP7_75t_L g1880 ( 
.A1(n_1873),
.A2(n_1840),
.B(n_1855),
.Y(n_1880)
);

NAND2xp5_ASAP7_75t_L g1881 ( 
.A(n_1873),
.B(n_1834),
.Y(n_1881)
);

NAND2xp5_ASAP7_75t_L g1882 ( 
.A(n_1877),
.B(n_1834),
.Y(n_1882)
);

INVx1_ASAP7_75t_L g1883 ( 
.A(n_1876),
.Y(n_1883)
);

NOR2xp33_ASAP7_75t_L g1884 ( 
.A(n_1875),
.B(n_1837),
.Y(n_1884)
);

NAND2xp5_ASAP7_75t_L g1885 ( 
.A(n_1879),
.B(n_1826),
.Y(n_1885)
);

NOR2xp67_ASAP7_75t_L g1886 ( 
.A(n_1881),
.B(n_108),
.Y(n_1886)
);

INVx1_ASAP7_75t_L g1887 ( 
.A(n_1878),
.Y(n_1887)
);

INVx1_ASAP7_75t_L g1888 ( 
.A(n_1880),
.Y(n_1888)
);

INVx1_ASAP7_75t_L g1889 ( 
.A(n_1876),
.Y(n_1889)
);

INVx1_ASAP7_75t_L g1890 ( 
.A(n_1876),
.Y(n_1890)
);

CKINVDCx16_ASAP7_75t_R g1891 ( 
.A(n_1876),
.Y(n_1891)
);

NOR3xp33_ASAP7_75t_L g1892 ( 
.A(n_1891),
.B(n_1822),
.C(n_110),
.Y(n_1892)
);

AOI222xp33_ASAP7_75t_L g1893 ( 
.A1(n_1888),
.A2(n_1854),
.B1(n_1838),
.B2(n_1822),
.C1(n_1831),
.C2(n_1813),
.Y(n_1893)
);

NOR2xp33_ASAP7_75t_L g1894 ( 
.A(n_1883),
.B(n_1838),
.Y(n_1894)
);

AOI211xp5_ASAP7_75t_L g1895 ( 
.A1(n_1890),
.A2(n_1822),
.B(n_1850),
.C(n_1854),
.Y(n_1895)
);

AOI221xp5_ASAP7_75t_L g1896 ( 
.A1(n_1889),
.A2(n_1829),
.B1(n_1825),
.B2(n_1810),
.C(n_1823),
.Y(n_1896)
);

INVx1_ASAP7_75t_L g1897 ( 
.A(n_1887),
.Y(n_1897)
);

AOI21xp33_ASAP7_75t_SL g1898 ( 
.A1(n_1884),
.A2(n_111),
.B(n_112),
.Y(n_1898)
);

NAND2xp5_ASAP7_75t_L g1899 ( 
.A(n_1886),
.B(n_1825),
.Y(n_1899)
);

AOI221xp5_ASAP7_75t_L g1900 ( 
.A1(n_1882),
.A2(n_1829),
.B1(n_1823),
.B2(n_1826),
.C(n_1818),
.Y(n_1900)
);

INVx1_ASAP7_75t_L g1901 ( 
.A(n_1885),
.Y(n_1901)
);

AOI211xp5_ASAP7_75t_L g1902 ( 
.A1(n_1888),
.A2(n_1807),
.B(n_113),
.C(n_111),
.Y(n_1902)
);

NAND4xp25_ASAP7_75t_SL g1903 ( 
.A(n_1888),
.B(n_1798),
.C(n_1818),
.D(n_115),
.Y(n_1903)
);

AOI221xp5_ASAP7_75t_L g1904 ( 
.A1(n_1888),
.A2(n_1814),
.B1(n_1527),
.B2(n_115),
.C(n_116),
.Y(n_1904)
);

NOR2xp33_ASAP7_75t_L g1905 ( 
.A(n_1888),
.B(n_112),
.Y(n_1905)
);

AOI211xp5_ASAP7_75t_L g1906 ( 
.A1(n_1888),
.A2(n_117),
.B(n_114),
.C(n_116),
.Y(n_1906)
);

AOI221xp5_ASAP7_75t_L g1907 ( 
.A1(n_1888),
.A2(n_1814),
.B1(n_118),
.B2(n_119),
.C(n_120),
.Y(n_1907)
);

OAI311xp33_ASAP7_75t_L g1908 ( 
.A1(n_1888),
.A2(n_114),
.A3(n_119),
.B1(n_1814),
.C1(n_1604),
.Y(n_1908)
);

INVx3_ASAP7_75t_SL g1909 ( 
.A(n_1897),
.Y(n_1909)
);

AOI22xp5_ASAP7_75t_L g1910 ( 
.A1(n_1894),
.A2(n_1814),
.B1(n_1797),
.B2(n_1532),
.Y(n_1910)
);

O2A1O1Ixp33_ASAP7_75t_L g1911 ( 
.A1(n_1905),
.A2(n_1797),
.B(n_131),
.C(n_132),
.Y(n_1911)
);

INVx1_ASAP7_75t_L g1912 ( 
.A(n_1899),
.Y(n_1912)
);

INVx2_ASAP7_75t_L g1913 ( 
.A(n_1901),
.Y(n_1913)
);

AOI321xp33_ASAP7_75t_L g1914 ( 
.A1(n_1898),
.A2(n_1797),
.A3(n_133),
.B1(n_134),
.B2(n_135),
.C(n_137),
.Y(n_1914)
);

AOI21xp5_ASAP7_75t_L g1915 ( 
.A1(n_1906),
.A2(n_1539),
.B(n_1520),
.Y(n_1915)
);

AOI221xp5_ASAP7_75t_L g1916 ( 
.A1(n_1903),
.A2(n_1539),
.B1(n_139),
.B2(n_141),
.C(n_142),
.Y(n_1916)
);

BUFx6f_ASAP7_75t_L g1917 ( 
.A(n_1892),
.Y(n_1917)
);

A2O1A1Ixp33_ASAP7_75t_L g1918 ( 
.A1(n_1902),
.A2(n_1539),
.B(n_143),
.C(n_144),
.Y(n_1918)
);

AOI21xp33_ASAP7_75t_SL g1919 ( 
.A1(n_1893),
.A2(n_130),
.B(n_147),
.Y(n_1919)
);

INVx1_ASAP7_75t_L g1920 ( 
.A(n_1907),
.Y(n_1920)
);

INVx1_ASAP7_75t_L g1921 ( 
.A(n_1900),
.Y(n_1921)
);

INVx1_ASAP7_75t_L g1922 ( 
.A(n_1904),
.Y(n_1922)
);

NAND2xp33_ASAP7_75t_R g1923 ( 
.A(n_1908),
.B(n_1895),
.Y(n_1923)
);

AOI221xp5_ASAP7_75t_L g1924 ( 
.A1(n_1896),
.A2(n_152),
.B1(n_154),
.B2(n_155),
.C(n_163),
.Y(n_1924)
);

OAI222xp33_ASAP7_75t_L g1925 ( 
.A1(n_1897),
.A2(n_165),
.B1(n_166),
.B2(n_167),
.C1(n_169),
.C2(n_170),
.Y(n_1925)
);

INVx1_ASAP7_75t_L g1926 ( 
.A(n_1899),
.Y(n_1926)
);

INVxp67_ASAP7_75t_SL g1927 ( 
.A(n_1906),
.Y(n_1927)
);

NAND2xp5_ASAP7_75t_SL g1928 ( 
.A(n_1919),
.B(n_171),
.Y(n_1928)
);

NAND2xp5_ASAP7_75t_L g1929 ( 
.A(n_1916),
.B(n_173),
.Y(n_1929)
);

NAND2xp5_ASAP7_75t_L g1930 ( 
.A(n_1927),
.B(n_174),
.Y(n_1930)
);

NAND3xp33_ASAP7_75t_L g1931 ( 
.A(n_1913),
.B(n_1920),
.C(n_1917),
.Y(n_1931)
);

INVx1_ASAP7_75t_L g1932 ( 
.A(n_1917),
.Y(n_1932)
);

OR2x2_ASAP7_75t_L g1933 ( 
.A(n_1909),
.B(n_175),
.Y(n_1933)
);

NOR2x1_ASAP7_75t_L g1934 ( 
.A(n_1922),
.B(n_180),
.Y(n_1934)
);

AND2x2_ASAP7_75t_L g1935 ( 
.A(n_1921),
.B(n_182),
.Y(n_1935)
);

INVx1_ASAP7_75t_L g1936 ( 
.A(n_1912),
.Y(n_1936)
);

AND2x4_ASAP7_75t_L g1937 ( 
.A(n_1926),
.B(n_183),
.Y(n_1937)
);

NOR3xp33_ASAP7_75t_L g1938 ( 
.A(n_1925),
.B(n_184),
.C(n_185),
.Y(n_1938)
);

NAND2xp5_ASAP7_75t_L g1939 ( 
.A(n_1918),
.B(n_187),
.Y(n_1939)
);

NAND2xp5_ASAP7_75t_L g1940 ( 
.A(n_1924),
.B(n_188),
.Y(n_1940)
);

NOR3x1_ASAP7_75t_L g1941 ( 
.A(n_1923),
.B(n_190),
.C(n_192),
.Y(n_1941)
);

INVx1_ASAP7_75t_L g1942 ( 
.A(n_1914),
.Y(n_1942)
);

INVxp67_ASAP7_75t_L g1943 ( 
.A(n_1915),
.Y(n_1943)
);

INVx1_ASAP7_75t_SL g1944 ( 
.A(n_1910),
.Y(n_1944)
);

INVxp67_ASAP7_75t_L g1945 ( 
.A(n_1911),
.Y(n_1945)
);

AND2x2_ASAP7_75t_L g1946 ( 
.A(n_1927),
.B(n_193),
.Y(n_1946)
);

AOI221xp5_ASAP7_75t_L g1947 ( 
.A1(n_1942),
.A2(n_195),
.B1(n_196),
.B2(n_197),
.C(n_198),
.Y(n_1947)
);

INVx1_ASAP7_75t_L g1948 ( 
.A(n_1930),
.Y(n_1948)
);

NOR2xp33_ASAP7_75t_L g1949 ( 
.A(n_1945),
.B(n_202),
.Y(n_1949)
);

INVx1_ASAP7_75t_L g1950 ( 
.A(n_1936),
.Y(n_1950)
);

AND2x2_ASAP7_75t_SL g1951 ( 
.A(n_1941),
.B(n_1946),
.Y(n_1951)
);

O2A1O1Ixp33_ASAP7_75t_L g1952 ( 
.A1(n_1943),
.A2(n_205),
.B(n_206),
.C(n_212),
.Y(n_1952)
);

OR2x2_ASAP7_75t_L g1953 ( 
.A(n_1931),
.B(n_214),
.Y(n_1953)
);

XNOR2xp5_ASAP7_75t_L g1954 ( 
.A(n_1928),
.B(n_219),
.Y(n_1954)
);

AOI222xp33_ASAP7_75t_L g1955 ( 
.A1(n_1935),
.A2(n_220),
.B1(n_225),
.B2(n_228),
.C1(n_229),
.C2(n_232),
.Y(n_1955)
);

O2A1O1Ixp5_ASAP7_75t_L g1956 ( 
.A1(n_1932),
.A2(n_234),
.B(n_239),
.C(n_241),
.Y(n_1956)
);

INVx3_ASAP7_75t_L g1957 ( 
.A(n_1937),
.Y(n_1957)
);

INVx1_ASAP7_75t_SL g1958 ( 
.A(n_1937),
.Y(n_1958)
);

INVx2_ASAP7_75t_SL g1959 ( 
.A(n_1933),
.Y(n_1959)
);

AOI211xp5_ASAP7_75t_L g1960 ( 
.A1(n_1938),
.A2(n_244),
.B(n_247),
.C(n_249),
.Y(n_1960)
);

AOI22xp5_ASAP7_75t_L g1961 ( 
.A1(n_1951),
.A2(n_1944),
.B1(n_1934),
.B2(n_1929),
.Y(n_1961)
);

AND2x4_ASAP7_75t_L g1962 ( 
.A(n_1957),
.B(n_1939),
.Y(n_1962)
);

AOI21xp5_ASAP7_75t_L g1963 ( 
.A1(n_1958),
.A2(n_1940),
.B(n_251),
.Y(n_1963)
);

NAND2xp5_ASAP7_75t_L g1964 ( 
.A(n_1947),
.B(n_252),
.Y(n_1964)
);

NOR2xp67_ASAP7_75t_L g1965 ( 
.A(n_1953),
.B(n_1950),
.Y(n_1965)
);

NOR2xp33_ASAP7_75t_L g1966 ( 
.A(n_1949),
.B(n_253),
.Y(n_1966)
);

OAI221xp5_ASAP7_75t_L g1967 ( 
.A1(n_1960),
.A2(n_257),
.B1(n_258),
.B2(n_259),
.C(n_260),
.Y(n_1967)
);

NAND4xp75_ASAP7_75t_L g1968 ( 
.A(n_1956),
.B(n_448),
.C(n_262),
.D(n_263),
.Y(n_1968)
);

OAI21xp5_ASAP7_75t_L g1969 ( 
.A1(n_1959),
.A2(n_261),
.B(n_264),
.Y(n_1969)
);

NAND4xp75_ASAP7_75t_L g1970 ( 
.A(n_1948),
.B(n_266),
.C(n_268),
.D(n_270),
.Y(n_1970)
);

O2A1O1Ixp33_ASAP7_75t_L g1971 ( 
.A1(n_1952),
.A2(n_274),
.B(n_276),
.C(n_279),
.Y(n_1971)
);

INVx5_ASAP7_75t_L g1972 ( 
.A(n_1954),
.Y(n_1972)
);

NOR2x1p5_ASAP7_75t_L g1973 ( 
.A(n_1968),
.B(n_1955),
.Y(n_1973)
);

AND2x2_ASAP7_75t_L g1974 ( 
.A(n_1962),
.B(n_281),
.Y(n_1974)
);

AND4x2_ASAP7_75t_L g1975 ( 
.A(n_1963),
.B(n_282),
.C(n_283),
.D(n_284),
.Y(n_1975)
);

BUFx12f_ASAP7_75t_L g1976 ( 
.A(n_1972),
.Y(n_1976)
);

NAND4xp75_ASAP7_75t_L g1977 ( 
.A(n_1965),
.B(n_286),
.C(n_292),
.D(n_294),
.Y(n_1977)
);

NAND4xp75_ASAP7_75t_L g1978 ( 
.A(n_1969),
.B(n_295),
.C(n_297),
.D(n_298),
.Y(n_1978)
);

NOR2x1_ASAP7_75t_L g1979 ( 
.A(n_1964),
.B(n_1970),
.Y(n_1979)
);

AND2x2_ASAP7_75t_L g1980 ( 
.A(n_1972),
.B(n_300),
.Y(n_1980)
);

NOR3xp33_ASAP7_75t_L g1981 ( 
.A(n_1967),
.B(n_301),
.C(n_304),
.Y(n_1981)
);

INVx2_ASAP7_75t_L g1982 ( 
.A(n_1974),
.Y(n_1982)
);

AOI322xp5_ASAP7_75t_L g1983 ( 
.A1(n_1979),
.A2(n_1961),
.A3(n_1966),
.B1(n_1971),
.B2(n_311),
.C1(n_312),
.C2(n_314),
.Y(n_1983)
);

NOR3xp33_ASAP7_75t_L g1984 ( 
.A(n_1977),
.B(n_306),
.C(n_308),
.Y(n_1984)
);

AOI322xp5_ASAP7_75t_L g1985 ( 
.A1(n_1981),
.A2(n_310),
.A3(n_315),
.B1(n_322),
.B2(n_323),
.C1(n_325),
.C2(n_330),
.Y(n_1985)
);

INVx1_ASAP7_75t_L g1986 ( 
.A(n_1980),
.Y(n_1986)
);

NOR2xp33_ASAP7_75t_L g1987 ( 
.A(n_1976),
.B(n_332),
.Y(n_1987)
);

INVx1_ASAP7_75t_L g1988 ( 
.A(n_1987),
.Y(n_1988)
);

OR5x1_ASAP7_75t_L g1989 ( 
.A(n_1983),
.B(n_1973),
.C(n_1975),
.D(n_1978),
.E(n_340),
.Y(n_1989)
);

INVx1_ASAP7_75t_SL g1990 ( 
.A(n_1982),
.Y(n_1990)
);

AOI21xp5_ASAP7_75t_SL g1991 ( 
.A1(n_1988),
.A2(n_1986),
.B(n_1985),
.Y(n_1991)
);

INVx1_ASAP7_75t_L g1992 ( 
.A(n_1990),
.Y(n_1992)
);

INVx1_ASAP7_75t_L g1993 ( 
.A(n_1989),
.Y(n_1993)
);

INVx1_ASAP7_75t_L g1994 ( 
.A(n_1992),
.Y(n_1994)
);

AOI22x1_ASAP7_75t_L g1995 ( 
.A1(n_1993),
.A2(n_1984),
.B1(n_338),
.B2(n_339),
.Y(n_1995)
);

OAI22xp5_ASAP7_75t_L g1996 ( 
.A1(n_1991),
.A2(n_336),
.B1(n_341),
.B2(n_343),
.Y(n_1996)
);

HB1xp67_ASAP7_75t_L g1997 ( 
.A(n_1994),
.Y(n_1997)
);

INVx1_ASAP7_75t_L g1998 ( 
.A(n_1996),
.Y(n_1998)
);

OA21x2_ASAP7_75t_L g1999 ( 
.A1(n_1998),
.A2(n_1995),
.B(n_347),
.Y(n_1999)
);

AOI21xp5_ASAP7_75t_L g2000 ( 
.A1(n_1999),
.A2(n_1997),
.B(n_349),
.Y(n_2000)
);

AOI222xp33_ASAP7_75t_L g2001 ( 
.A1(n_2000),
.A2(n_344),
.B1(n_355),
.B2(n_356),
.C1(n_358),
.C2(n_361),
.Y(n_2001)
);

AOI22xp5_ASAP7_75t_L g2002 ( 
.A1(n_2001),
.A2(n_364),
.B1(n_366),
.B2(n_367),
.Y(n_2002)
);

AOI211xp5_ASAP7_75t_L g2003 ( 
.A1(n_2002),
.A2(n_444),
.B(n_371),
.C(n_373),
.Y(n_2003)
);


endmodule