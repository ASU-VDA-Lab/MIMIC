module fake_jpeg_3420_n_654 (n_13, n_1, n_10, n_6, n_14, n_18, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_654);

input n_13;
input n_1;
input n_10;
input n_6;
input n_14;
input n_18;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_654;

wire n_529;
wire n_595;
wire n_390;
wire n_552;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_525;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_586;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_620;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_611;
wire n_44;
wire n_355;
wire n_519;
wire n_276;
wire n_143;
wire n_431;
wire n_102;
wire n_549;
wire n_196;
wire n_66;
wire n_374;
wire n_566;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_597;
wire n_172;
wire n_547;
wire n_345;
wire n_591;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_513;
wire n_283;
wire n_107;
wire n_490;
wire n_635;
wire n_517;
wire n_629;
wire n_415;
wire n_479;
wire n_543;
wire n_357;
wire n_89;
wire n_131;
wire n_607;
wire n_294;
wire n_230;
wire n_643;
wire n_170;
wire n_602;
wire n_313;
wire n_542;
wire n_574;
wire n_264;
wire n_647;
wire n_437;
wire n_93;
wire n_227;
wire n_559;
wire n_641;
wire n_48;
wire n_465;
wire n_638;
wire n_200;
wire n_582;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_623;
wire n_579;
wire n_416;
wire n_256;
wire n_221;
wire n_454;
wire n_540;
wire n_292;
wire n_213;
wire n_135;
wire n_435;
wire n_189;
wire n_637;
wire n_370;
wire n_410;
wire n_571;
wire n_82;
wire n_155;
wire n_508;
wire n_309;
wire n_624;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_606;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_569;
wire n_596;
wire n_400;
wire n_646;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_544;
wire n_31;
wire n_277;
wire n_255;
wire n_605;
wire n_601;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_349;
wire n_21;
wire n_393;
wire n_288;
wire n_234;
wire n_530;
wire n_634;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_557;
wire n_408;
wire n_80;
wire n_562;
wire n_204;
wire n_639;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_645;
wire n_298;
wire n_106;
wire n_545;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_584;
wire n_254;
wire n_608;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_622;
wire n_463;
wire n_92;
wire n_332;
wire n_640;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_653;
wire n_474;
wire n_539;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_626;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_575;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_511;
wire n_305;
wire n_161;
wire n_441;
wire n_555;
wire n_342;
wire n_642;
wire n_101;
wire n_226;
wire n_509;
wire n_644;
wire n_149;
wire n_87;
wire n_46;
wire n_578;
wire n_589;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_614;
wire n_97;
wire n_649;
wire n_573;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_610;
wire n_174;
wire n_198;
wire n_422;
wire n_560;
wire n_190;
wire n_510;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_536;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_537;
wire n_110;
wire n_594;
wire n_590;
wire n_531;
wire n_76;
wire n_278;
wire n_343;
wire n_577;
wire n_26;
wire n_88;
wire n_397;
wire n_592;
wire n_363;
wire n_570;
wire n_238;
wire n_598;
wire n_615;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_554;
wire n_301;
wire n_609;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_648;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_523;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_533;
wire n_612;
wire n_384;
wire n_296;
wire n_588;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_585;
wire n_491;
wire n_24;
wire n_526;
wire n_467;
wire n_269;
wire n_572;
wire n_546;
wire n_287;
wire n_219;
wire n_452;
wire n_631;
wire n_433;
wire n_636;
wire n_77;
wire n_473;
wire n_45;
wire n_520;
wire n_476;
wire n_337;
wire n_317;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_650;
wire n_218;
wire n_63;
wire n_652;
wire n_599;
wire n_239;
wire n_243;
wire n_481;
wire n_628;
wire n_619;
wire n_348;
wire n_587;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_583;
wire n_522;
wire n_333;
wire n_518;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_565;
wire n_302;
wire n_216;
wire n_528;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_199;
wire n_260;
wire n_550;
wire n_413;
wire n_275;
wire n_494;
wire n_604;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_551;
wire n_36;
wire n_62;
wire n_600;
wire n_492;
wire n_603;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_567;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_515;
wire n_347;
wire n_521;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_538;
wire n_625;
wire n_147;
wire n_449;
wire n_627;
wire n_98;
wire n_251;
wire n_534;
wire n_472;
wire n_279;
wire n_593;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_618;
wire n_356;
wire n_119;
wire n_484;
wire n_568;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_576;
wire n_469;
wire n_111;
wire n_197;
wire n_396;
wire n_375;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_553;
wire n_257;
wire n_61;
wire n_173;
wire n_561;
wire n_244;
wire n_232;
wire n_527;
wire n_482;
wire n_58;
wire n_41;
wire n_613;
wire n_630;
wire n_266;
wire n_548;
wire n_72;
wire n_512;
wire n_445;
wire n_443;
wire n_617;
wire n_215;
wire n_212;
wire n_516;
wire n_183;
wire n_409;
wire n_532;
wire n_249;
wire n_412;
wire n_581;
wire n_217;
wire n_471;
wire n_580;
wire n_541;
wire n_53;
wire n_372;
wire n_558;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_535;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_556;
wire n_524;
wire n_402;
wire n_563;
wire n_504;
wire n_438;
wire n_475;
wire n_247;
wire n_157;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_633;
wire n_112;
wire n_632;
wire n_616;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_514;
wire n_651;
wire n_564;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_621;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

BUFx8_ASAP7_75t_L g19 ( 
.A(n_4),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_18),
.Y(n_20)
);

BUFx3_ASAP7_75t_L g21 ( 
.A(n_0),
.Y(n_21)
);

BUFx5_ASAP7_75t_L g22 ( 
.A(n_0),
.Y(n_22)
);

NOR2xp33_ASAP7_75t_L g23 ( 
.A(n_1),
.B(n_5),
.Y(n_23)
);

BUFx5_ASAP7_75t_L g24 ( 
.A(n_0),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_11),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_13),
.Y(n_26)
);

BUFx12_ASAP7_75t_L g27 ( 
.A(n_3),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_15),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_16),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_18),
.Y(n_30)
);

BUFx16f_ASAP7_75t_L g31 ( 
.A(n_18),
.Y(n_31)
);

INVx4_ASAP7_75t_L g32 ( 
.A(n_6),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_3),
.Y(n_33)
);

BUFx5_ASAP7_75t_L g34 ( 
.A(n_14),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_17),
.Y(n_35)
);

BUFx12f_ASAP7_75t_L g36 ( 
.A(n_1),
.Y(n_36)
);

BUFx12_ASAP7_75t_L g37 ( 
.A(n_16),
.Y(n_37)
);

INVx6_ASAP7_75t_L g38 ( 
.A(n_8),
.Y(n_38)
);

BUFx3_ASAP7_75t_L g39 ( 
.A(n_2),
.Y(n_39)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_9),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g41 ( 
.A(n_11),
.B(n_7),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_14),
.Y(n_42)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_8),
.Y(n_43)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_2),
.Y(n_44)
);

BUFx3_ASAP7_75t_L g45 ( 
.A(n_4),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_12),
.Y(n_46)
);

INVx6_ASAP7_75t_L g47 ( 
.A(n_2),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_17),
.Y(n_48)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_8),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_5),
.Y(n_50)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_16),
.Y(n_51)
);

BUFx4f_ASAP7_75t_SL g52 ( 
.A(n_2),
.Y(n_52)
);

BUFx24_ASAP7_75t_L g53 ( 
.A(n_13),
.Y(n_53)
);

INVx3_ASAP7_75t_L g54 ( 
.A(n_4),
.Y(n_54)
);

BUFx12f_ASAP7_75t_L g55 ( 
.A(n_13),
.Y(n_55)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_1),
.Y(n_56)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_8),
.Y(n_57)
);

BUFx3_ASAP7_75t_L g58 ( 
.A(n_18),
.Y(n_58)
);

BUFx24_ASAP7_75t_L g59 ( 
.A(n_16),
.Y(n_59)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_52),
.Y(n_60)
);

INVx2_ASAP7_75t_L g130 ( 
.A(n_60),
.Y(n_130)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_20),
.Y(n_61)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_61),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_SL g62 ( 
.A(n_41),
.B(n_9),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g145 ( 
.A(n_62),
.B(n_83),
.Y(n_145)
);

INVx5_ASAP7_75t_L g63 ( 
.A(n_21),
.Y(n_63)
);

BUFx3_ASAP7_75t_L g203 ( 
.A(n_63),
.Y(n_203)
);

INVx2_ASAP7_75t_L g64 ( 
.A(n_52),
.Y(n_64)
);

INVx2_ASAP7_75t_L g131 ( 
.A(n_64),
.Y(n_131)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_26),
.Y(n_65)
);

BUFx6f_ASAP7_75t_L g124 ( 
.A(n_65),
.Y(n_124)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_26),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g139 ( 
.A(n_66),
.Y(n_139)
);

BUFx3_ASAP7_75t_L g67 ( 
.A(n_45),
.Y(n_67)
);

BUFx2_ASAP7_75t_L g159 ( 
.A(n_67),
.Y(n_159)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_26),
.Y(n_68)
);

BUFx6f_ASAP7_75t_L g152 ( 
.A(n_68),
.Y(n_152)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_20),
.Y(n_69)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_69),
.Y(n_162)
);

BUFx6f_ASAP7_75t_L g70 ( 
.A(n_28),
.Y(n_70)
);

BUFx6f_ASAP7_75t_L g156 ( 
.A(n_70),
.Y(n_156)
);

INVx2_ASAP7_75t_L g71 ( 
.A(n_52),
.Y(n_71)
);

INVx2_ASAP7_75t_L g133 ( 
.A(n_71),
.Y(n_133)
);

INVx2_ASAP7_75t_L g72 ( 
.A(n_52),
.Y(n_72)
);

INVx2_ASAP7_75t_L g136 ( 
.A(n_72),
.Y(n_136)
);

BUFx6f_ASAP7_75t_L g73 ( 
.A(n_28),
.Y(n_73)
);

BUFx6f_ASAP7_75t_L g161 ( 
.A(n_73),
.Y(n_161)
);

BUFx6f_ASAP7_75t_L g74 ( 
.A(n_28),
.Y(n_74)
);

BUFx6f_ASAP7_75t_L g178 ( 
.A(n_74),
.Y(n_178)
);

INVx6_ASAP7_75t_L g75 ( 
.A(n_42),
.Y(n_75)
);

INVx3_ASAP7_75t_SL g144 ( 
.A(n_75),
.Y(n_144)
);

BUFx6f_ASAP7_75t_L g76 ( 
.A(n_42),
.Y(n_76)
);

INVx6_ASAP7_75t_L g128 ( 
.A(n_76),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_41),
.B(n_9),
.Y(n_77)
);

A2O1A1Ixp33_ASAP7_75t_L g153 ( 
.A1(n_77),
.A2(n_29),
.B(n_35),
.C(n_46),
.Y(n_153)
);

INVx2_ASAP7_75t_L g78 ( 
.A(n_32),
.Y(n_78)
);

INVx2_ASAP7_75t_L g143 ( 
.A(n_78),
.Y(n_143)
);

BUFx3_ASAP7_75t_L g79 ( 
.A(n_58),
.Y(n_79)
);

BUFx2_ASAP7_75t_L g170 ( 
.A(n_79),
.Y(n_170)
);

HB1xp67_ASAP7_75t_L g80 ( 
.A(n_36),
.Y(n_80)
);

INVx2_ASAP7_75t_L g151 ( 
.A(n_80),
.Y(n_151)
);

INVx2_ASAP7_75t_L g81 ( 
.A(n_32),
.Y(n_81)
);

INVx2_ASAP7_75t_L g163 ( 
.A(n_81),
.Y(n_163)
);

BUFx6f_ASAP7_75t_L g82 ( 
.A(n_42),
.Y(n_82)
);

INVx6_ASAP7_75t_L g183 ( 
.A(n_82),
.Y(n_183)
);

NOR2xp33_ASAP7_75t_SL g83 ( 
.A(n_23),
.B(n_9),
.Y(n_83)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_40),
.Y(n_84)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_84),
.Y(n_164)
);

BUFx6f_ASAP7_75t_L g85 ( 
.A(n_48),
.Y(n_85)
);

INVx8_ASAP7_75t_L g171 ( 
.A(n_85),
.Y(n_171)
);

INVx13_ASAP7_75t_L g86 ( 
.A(n_19),
.Y(n_86)
);

INVx2_ASAP7_75t_SL g146 ( 
.A(n_86),
.Y(n_146)
);

INVx4_ASAP7_75t_L g87 ( 
.A(n_22),
.Y(n_87)
);

INVx2_ASAP7_75t_SL g200 ( 
.A(n_87),
.Y(n_200)
);

BUFx6f_ASAP7_75t_L g88 ( 
.A(n_48),
.Y(n_88)
);

INVx8_ASAP7_75t_L g196 ( 
.A(n_88),
.Y(n_196)
);

INVx2_ASAP7_75t_L g89 ( 
.A(n_54),
.Y(n_89)
);

INVx2_ASAP7_75t_L g167 ( 
.A(n_89),
.Y(n_167)
);

INVx11_ASAP7_75t_L g90 ( 
.A(n_19),
.Y(n_90)
);

INVx4_ASAP7_75t_L g138 ( 
.A(n_90),
.Y(n_138)
);

INVx4_ASAP7_75t_L g91 ( 
.A(n_22),
.Y(n_91)
);

INVx3_ASAP7_75t_L g134 ( 
.A(n_91),
.Y(n_134)
);

INVx3_ASAP7_75t_L g92 ( 
.A(n_31),
.Y(n_92)
);

INVx3_ASAP7_75t_L g142 ( 
.A(n_92),
.Y(n_142)
);

INVx2_ASAP7_75t_L g93 ( 
.A(n_54),
.Y(n_93)
);

INVx2_ASAP7_75t_L g181 ( 
.A(n_93),
.Y(n_181)
);

BUFx12f_ASAP7_75t_L g94 ( 
.A(n_19),
.Y(n_94)
);

INVx5_ASAP7_75t_L g132 ( 
.A(n_94),
.Y(n_132)
);

BUFx6f_ASAP7_75t_L g95 ( 
.A(n_48),
.Y(n_95)
);

INVx5_ASAP7_75t_L g148 ( 
.A(n_95),
.Y(n_148)
);

BUFx3_ASAP7_75t_L g96 ( 
.A(n_58),
.Y(n_96)
);

INVx5_ASAP7_75t_L g149 ( 
.A(n_96),
.Y(n_149)
);

INVx2_ASAP7_75t_L g97 ( 
.A(n_47),
.Y(n_97)
);

INVx2_ASAP7_75t_L g185 ( 
.A(n_97),
.Y(n_185)
);

INVx3_ASAP7_75t_L g98 ( 
.A(n_31),
.Y(n_98)
);

INVx3_ASAP7_75t_L g154 ( 
.A(n_98),
.Y(n_154)
);

INVx3_ASAP7_75t_L g99 ( 
.A(n_31),
.Y(n_99)
);

INVx3_ASAP7_75t_L g160 ( 
.A(n_99),
.Y(n_160)
);

INVx6_ASAP7_75t_L g100 ( 
.A(n_33),
.Y(n_100)
);

INVx2_ASAP7_75t_L g187 ( 
.A(n_100),
.Y(n_187)
);

AND2x2_ASAP7_75t_L g101 ( 
.A(n_23),
.B(n_7),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_L g173 ( 
.A(n_101),
.B(n_29),
.Y(n_173)
);

INVx2_ASAP7_75t_L g102 ( 
.A(n_47),
.Y(n_102)
);

INVx2_ASAP7_75t_L g191 ( 
.A(n_102),
.Y(n_191)
);

INVx4_ASAP7_75t_L g103 ( 
.A(n_24),
.Y(n_103)
);

INVx3_ASAP7_75t_L g176 ( 
.A(n_103),
.Y(n_176)
);

INVx3_ASAP7_75t_L g104 ( 
.A(n_31),
.Y(n_104)
);

INVx3_ASAP7_75t_L g188 ( 
.A(n_104),
.Y(n_188)
);

INVx2_ASAP7_75t_L g105 ( 
.A(n_47),
.Y(n_105)
);

INVx2_ASAP7_75t_L g192 ( 
.A(n_105),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_L g106 ( 
.A(n_25),
.B(n_17),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_L g125 ( 
.A(n_106),
.B(n_121),
.Y(n_125)
);

INVx3_ASAP7_75t_L g107 ( 
.A(n_36),
.Y(n_107)
);

INVx3_ASAP7_75t_L g189 ( 
.A(n_107),
.Y(n_189)
);

BUFx6f_ASAP7_75t_L g108 ( 
.A(n_33),
.Y(n_108)
);

INVx5_ASAP7_75t_L g158 ( 
.A(n_108),
.Y(n_158)
);

INVx8_ASAP7_75t_L g109 ( 
.A(n_36),
.Y(n_109)
);

INVx5_ASAP7_75t_L g175 ( 
.A(n_109),
.Y(n_175)
);

INVx8_ASAP7_75t_L g110 ( 
.A(n_36),
.Y(n_110)
);

INVx3_ASAP7_75t_L g190 ( 
.A(n_110),
.Y(n_190)
);

BUFx5_ASAP7_75t_L g111 ( 
.A(n_19),
.Y(n_111)
);

INVx4_ASAP7_75t_L g140 ( 
.A(n_111),
.Y(n_140)
);

INVx4_ASAP7_75t_L g112 ( 
.A(n_24),
.Y(n_112)
);

INVx4_ASAP7_75t_L g141 ( 
.A(n_112),
.Y(n_141)
);

INVx8_ASAP7_75t_L g113 ( 
.A(n_55),
.Y(n_113)
);

INVx4_ASAP7_75t_L g147 ( 
.A(n_113),
.Y(n_147)
);

AOI22xp33_ASAP7_75t_SL g114 ( 
.A1(n_39),
.A2(n_7),
.B1(n_15),
.B2(n_14),
.Y(n_114)
);

AOI22xp33_ASAP7_75t_SL g127 ( 
.A1(n_114),
.A2(n_30),
.B1(n_50),
.B2(n_46),
.Y(n_127)
);

INVx3_ASAP7_75t_SL g115 ( 
.A(n_33),
.Y(n_115)
);

INVx2_ASAP7_75t_L g193 ( 
.A(n_115),
.Y(n_193)
);

BUFx6f_ASAP7_75t_L g116 ( 
.A(n_38),
.Y(n_116)
);

INVx2_ASAP7_75t_L g194 ( 
.A(n_116),
.Y(n_194)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_40),
.Y(n_117)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_117),
.Y(n_177)
);

BUFx6f_ASAP7_75t_L g118 ( 
.A(n_38),
.Y(n_118)
);

INVx2_ASAP7_75t_L g197 ( 
.A(n_118),
.Y(n_197)
);

INVx3_ASAP7_75t_L g119 ( 
.A(n_39),
.Y(n_119)
);

INVx4_ASAP7_75t_L g155 ( 
.A(n_119),
.Y(n_155)
);

INVx4_ASAP7_75t_L g120 ( 
.A(n_34),
.Y(n_120)
);

INVx4_ASAP7_75t_L g157 ( 
.A(n_120),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_L g121 ( 
.A(n_25),
.B(n_17),
.Y(n_121)
);

BUFx6f_ASAP7_75t_L g122 ( 
.A(n_38),
.Y(n_122)
);

INVx2_ASAP7_75t_L g198 ( 
.A(n_122),
.Y(n_198)
);

BUFx3_ASAP7_75t_L g123 ( 
.A(n_45),
.Y(n_123)
);

INVx4_ASAP7_75t_L g168 ( 
.A(n_123),
.Y(n_168)
);

AOI21xp5_ASAP7_75t_L g241 ( 
.A1(n_127),
.A2(n_114),
.B(n_59),
.Y(n_241)
);

CKINVDCx14_ASAP7_75t_SL g129 ( 
.A(n_86),
.Y(n_129)
);

BUFx10_ASAP7_75t_L g258 ( 
.A(n_129),
.Y(n_258)
);

NAND2xp5_ASAP7_75t_L g135 ( 
.A(n_77),
.B(n_51),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_L g239 ( 
.A(n_135),
.B(n_153),
.Y(n_239)
);

CKINVDCx20_ASAP7_75t_R g137 ( 
.A(n_80),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_L g211 ( 
.A(n_137),
.B(n_165),
.Y(n_211)
);

MAJIxp5_ASAP7_75t_L g150 ( 
.A(n_101),
.B(n_45),
.C(n_39),
.Y(n_150)
);

MAJIxp5_ASAP7_75t_L g269 ( 
.A(n_150),
.B(n_59),
.C(n_53),
.Y(n_269)
);

NOR2xp33_ASAP7_75t_SL g165 ( 
.A(n_67),
.B(n_35),
.Y(n_165)
);

AOI22xp33_ASAP7_75t_SL g166 ( 
.A1(n_94),
.A2(n_21),
.B1(n_55),
.B2(n_49),
.Y(n_166)
);

AOI22xp5_ASAP7_75t_SL g275 ( 
.A1(n_166),
.A2(n_53),
.B1(n_59),
.B2(n_34),
.Y(n_275)
);

NAND2xp5_ASAP7_75t_L g169 ( 
.A(n_115),
.B(n_43),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_L g225 ( 
.A(n_169),
.B(n_174),
.Y(n_225)
);

OAI22xp5_ASAP7_75t_L g172 ( 
.A1(n_75),
.A2(n_55),
.B1(n_30),
.B2(n_50),
.Y(n_172)
);

AOI22xp5_ASAP7_75t_L g233 ( 
.A1(n_172),
.A2(n_186),
.B1(n_70),
.B2(n_95),
.Y(n_233)
);

AND2x2_ASAP7_75t_L g210 ( 
.A(n_173),
.B(n_44),
.Y(n_210)
);

NOR2xp33_ASAP7_75t_L g174 ( 
.A(n_94),
.B(n_43),
.Y(n_174)
);

INVx4_ASAP7_75t_L g179 ( 
.A(n_109),
.Y(n_179)
);

INVx1_ASAP7_75t_SL g234 ( 
.A(n_179),
.Y(n_234)
);

INVx4_ASAP7_75t_L g180 ( 
.A(n_110),
.Y(n_180)
);

INVx4_ASAP7_75t_L g267 ( 
.A(n_180),
.Y(n_267)
);

INVx4_ASAP7_75t_L g182 ( 
.A(n_113),
.Y(n_182)
);

INVx3_ASAP7_75t_SL g219 ( 
.A(n_182),
.Y(n_219)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_100),
.Y(n_184)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_184),
.Y(n_206)
);

OAI22xp5_ASAP7_75t_L g186 ( 
.A1(n_65),
.A2(n_55),
.B1(n_57),
.B2(n_51),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_L g195 ( 
.A(n_108),
.B(n_57),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_L g235 ( 
.A(n_195),
.B(n_204),
.Y(n_235)
);

INVx2_ASAP7_75t_L g199 ( 
.A(n_116),
.Y(n_199)
);

INVx2_ASAP7_75t_L g207 ( 
.A(n_199),
.Y(n_207)
);

INVx2_ASAP7_75t_L g201 ( 
.A(n_118),
.Y(n_201)
);

INVx2_ASAP7_75t_L g213 ( 
.A(n_201),
.Y(n_213)
);

INVx4_ASAP7_75t_L g202 ( 
.A(n_123),
.Y(n_202)
);

BUFx2_ASAP7_75t_L g260 ( 
.A(n_202),
.Y(n_260)
);

NOR2xp33_ASAP7_75t_L g204 ( 
.A(n_122),
.B(n_49),
.Y(n_204)
);

INVx2_ASAP7_75t_L g205 ( 
.A(n_66),
.Y(n_205)
);

INVx2_ASAP7_75t_L g221 ( 
.A(n_205),
.Y(n_221)
);

INVx8_ASAP7_75t_L g208 ( 
.A(n_129),
.Y(n_208)
);

INVx3_ASAP7_75t_L g293 ( 
.A(n_208),
.Y(n_293)
);

CKINVDCx20_ASAP7_75t_R g209 ( 
.A(n_204),
.Y(n_209)
);

NOR2xp33_ASAP7_75t_SL g334 ( 
.A(n_209),
.B(n_210),
.Y(n_334)
);

NOR2xp33_ASAP7_75t_L g212 ( 
.A(n_126),
.B(n_56),
.Y(n_212)
);

NOR2xp33_ASAP7_75t_L g283 ( 
.A(n_212),
.B(n_217),
.Y(n_283)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_162),
.Y(n_214)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_214),
.Y(n_297)
);

INVx5_ASAP7_75t_L g215 ( 
.A(n_132),
.Y(n_215)
);

INVx4_ASAP7_75t_L g319 ( 
.A(n_215),
.Y(n_319)
);

BUFx6f_ASAP7_75t_L g216 ( 
.A(n_124),
.Y(n_216)
);

BUFx6f_ASAP7_75t_L g322 ( 
.A(n_216),
.Y(n_322)
);

CKINVDCx20_ASAP7_75t_R g217 ( 
.A(n_174),
.Y(n_217)
);

NOR2xp33_ASAP7_75t_L g218 ( 
.A(n_164),
.B(n_56),
.Y(n_218)
);

NOR2xp33_ASAP7_75t_L g284 ( 
.A(n_218),
.B(n_222),
.Y(n_284)
);

INVx8_ASAP7_75t_L g220 ( 
.A(n_124),
.Y(n_220)
);

INVx2_ASAP7_75t_L g285 ( 
.A(n_220),
.Y(n_285)
);

NOR2xp33_ASAP7_75t_L g222 ( 
.A(n_177),
.B(n_44),
.Y(n_222)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_146),
.Y(n_223)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_223),
.Y(n_323)
);

BUFx3_ASAP7_75t_L g224 ( 
.A(n_175),
.Y(n_224)
);

INVx2_ASAP7_75t_L g287 ( 
.A(n_224),
.Y(n_287)
);

BUFx6f_ASAP7_75t_L g226 ( 
.A(n_139),
.Y(n_226)
);

INVx2_ASAP7_75t_L g288 ( 
.A(n_226),
.Y(n_288)
);

NOR2xp33_ASAP7_75t_L g227 ( 
.A(n_145),
.B(n_74),
.Y(n_227)
);

NOR2xp33_ASAP7_75t_L g306 ( 
.A(n_227),
.B(n_230),
.Y(n_306)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_146),
.Y(n_228)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_228),
.Y(n_330)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_151),
.Y(n_229)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_229),
.Y(n_282)
);

NOR2xp33_ASAP7_75t_L g230 ( 
.A(n_145),
.B(n_73),
.Y(n_230)
);

INVx2_ASAP7_75t_L g231 ( 
.A(n_187),
.Y(n_231)
);

INVx2_ASAP7_75t_L g311 ( 
.A(n_231),
.Y(n_311)
);

INVx3_ASAP7_75t_L g232 ( 
.A(n_147),
.Y(n_232)
);

INVx4_ASAP7_75t_SL g337 ( 
.A(n_232),
.Y(n_337)
);

OA22x2_ASAP7_75t_L g286 ( 
.A1(n_233),
.A2(n_275),
.B1(n_166),
.B2(n_138),
.Y(n_286)
);

NAND2xp33_ASAP7_75t_SL g236 ( 
.A(n_170),
.B(n_0),
.Y(n_236)
);

OAI21xp5_ASAP7_75t_SL g292 ( 
.A1(n_236),
.A2(n_241),
.B(n_53),
.Y(n_292)
);

INVx8_ASAP7_75t_L g237 ( 
.A(n_139),
.Y(n_237)
);

INVx2_ASAP7_75t_L g321 ( 
.A(n_237),
.Y(n_321)
);

NOR2xp33_ASAP7_75t_L g238 ( 
.A(n_125),
.B(n_68),
.Y(n_238)
);

NOR2xp33_ASAP7_75t_L g314 ( 
.A(n_238),
.B(n_242),
.Y(n_314)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_130),
.Y(n_240)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_240),
.Y(n_289)
);

NOR2xp33_ASAP7_75t_L g242 ( 
.A(n_173),
.B(n_85),
.Y(n_242)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_131),
.Y(n_243)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_243),
.Y(n_290)
);

CKINVDCx20_ASAP7_75t_R g244 ( 
.A(n_159),
.Y(n_244)
);

NOR2xp33_ASAP7_75t_L g320 ( 
.A(n_244),
.B(n_247),
.Y(n_320)
);

INVx2_ASAP7_75t_L g245 ( 
.A(n_193),
.Y(n_245)
);

INVx2_ASAP7_75t_L g327 ( 
.A(n_245),
.Y(n_327)
);

AOI22xp33_ASAP7_75t_L g246 ( 
.A1(n_172),
.A2(n_186),
.B1(n_82),
.B2(n_76),
.Y(n_246)
);

OAI22xp33_ASAP7_75t_SL g329 ( 
.A1(n_246),
.A2(n_27),
.B1(n_37),
.B2(n_3),
.Y(n_329)
);

NOR2xp33_ASAP7_75t_L g247 ( 
.A(n_142),
.B(n_88),
.Y(n_247)
);

INVx2_ASAP7_75t_L g248 ( 
.A(n_185),
.Y(n_248)
);

INVx2_ASAP7_75t_L g328 ( 
.A(n_248),
.Y(n_328)
);

INVx2_ASAP7_75t_L g249 ( 
.A(n_191),
.Y(n_249)
);

INVx2_ASAP7_75t_L g332 ( 
.A(n_249),
.Y(n_332)
);

INVx2_ASAP7_75t_L g250 ( 
.A(n_192),
.Y(n_250)
);

INVx2_ASAP7_75t_L g339 ( 
.A(n_250),
.Y(n_339)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_133),
.Y(n_251)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_251),
.Y(n_294)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_136),
.Y(n_252)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_252),
.Y(n_304)
);

INVx6_ASAP7_75t_L g253 ( 
.A(n_152),
.Y(n_253)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_253),
.Y(n_305)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_143),
.Y(n_254)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_254),
.Y(n_316)
);

CKINVDCx20_ASAP7_75t_R g255 ( 
.A(n_159),
.Y(n_255)
);

NOR2xp33_ASAP7_75t_L g342 ( 
.A(n_255),
.B(n_264),
.Y(n_342)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_163),
.Y(n_256)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_256),
.Y(n_335)
);

INVx2_ASAP7_75t_L g257 ( 
.A(n_194),
.Y(n_257)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_257),
.Y(n_341)
);

INVx2_ASAP7_75t_L g259 ( 
.A(n_197),
.Y(n_259)
);

INVx1_ASAP7_75t_L g346 ( 
.A(n_259),
.Y(n_346)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_167),
.Y(n_261)
);

INVxp67_ASAP7_75t_L g296 ( 
.A(n_261),
.Y(n_296)
);

BUFx3_ASAP7_75t_L g262 ( 
.A(n_149),
.Y(n_262)
);

BUFx5_ASAP7_75t_L g310 ( 
.A(n_262),
.Y(n_310)
);

BUFx2_ASAP7_75t_L g263 ( 
.A(n_170),
.Y(n_263)
);

CKINVDCx16_ASAP7_75t_R g309 ( 
.A(n_263),
.Y(n_309)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_181),
.Y(n_264)
);

CKINVDCx20_ASAP7_75t_R g265 ( 
.A(n_148),
.Y(n_265)
);

CKINVDCx20_ASAP7_75t_R g295 ( 
.A(n_265),
.Y(n_295)
);

BUFx6f_ASAP7_75t_L g266 ( 
.A(n_152),
.Y(n_266)
);

CKINVDCx20_ASAP7_75t_R g307 ( 
.A(n_266),
.Y(n_307)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_154),
.Y(n_268)
);

AND2x2_ASAP7_75t_L g303 ( 
.A(n_268),
.B(n_272),
.Y(n_303)
);

XNOR2x1_ASAP7_75t_L g336 ( 
.A(n_269),
.B(n_37),
.Y(n_336)
);

BUFx6f_ASAP7_75t_L g270 ( 
.A(n_156),
.Y(n_270)
);

CKINVDCx20_ASAP7_75t_R g343 ( 
.A(n_270),
.Y(n_343)
);

BUFx8_ASAP7_75t_L g271 ( 
.A(n_140),
.Y(n_271)
);

BUFx5_ASAP7_75t_L g344 ( 
.A(n_271),
.Y(n_344)
);

INVx3_ASAP7_75t_L g272 ( 
.A(n_190),
.Y(n_272)
);

INVx2_ASAP7_75t_L g273 ( 
.A(n_198),
.Y(n_273)
);

CKINVDCx16_ASAP7_75t_R g318 ( 
.A(n_273),
.Y(n_318)
);

INVx5_ASAP7_75t_L g274 ( 
.A(n_196),
.Y(n_274)
);

AOI22xp33_ASAP7_75t_SL g302 ( 
.A1(n_274),
.A2(n_279),
.B1(n_281),
.B2(n_203),
.Y(n_302)
);

NOR2xp33_ASAP7_75t_L g276 ( 
.A(n_160),
.B(n_11),
.Y(n_276)
);

NAND2xp5_ASAP7_75t_L g291 ( 
.A(n_276),
.B(n_277),
.Y(n_291)
);

NAND2xp5_ASAP7_75t_L g277 ( 
.A(n_189),
.B(n_0),
.Y(n_277)
);

OAI22xp5_ASAP7_75t_SL g278 ( 
.A1(n_127),
.A2(n_59),
.B1(n_53),
.B2(n_27),
.Y(n_278)
);

AOI22xp5_ASAP7_75t_L g325 ( 
.A1(n_278),
.A2(n_171),
.B1(n_161),
.B2(n_27),
.Y(n_325)
);

BUFx2_ASAP7_75t_SL g279 ( 
.A(n_156),
.Y(n_279)
);

NAND2xp5_ASAP7_75t_L g280 ( 
.A(n_155),
.B(n_1),
.Y(n_280)
);

NAND2xp5_ASAP7_75t_L g298 ( 
.A(n_280),
.B(n_1),
.Y(n_298)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_188),
.Y(n_281)
);

OAI21xp33_ASAP7_75t_SL g377 ( 
.A1(n_286),
.A2(n_292),
.B(n_312),
.Y(n_377)
);

NAND2xp5_ASAP7_75t_SL g375 ( 
.A(n_298),
.B(n_249),
.Y(n_375)
);

AOI21xp5_ASAP7_75t_L g299 ( 
.A1(n_241),
.A2(n_200),
.B(n_176),
.Y(n_299)
);

AOI21xp5_ASAP7_75t_L g365 ( 
.A1(n_299),
.A2(n_267),
.B(n_260),
.Y(n_365)
);

OAI22xp5_ASAP7_75t_SL g300 ( 
.A1(n_233),
.A2(n_144),
.B1(n_128),
.B2(n_183),
.Y(n_300)
);

AOI22xp5_ASAP7_75t_L g361 ( 
.A1(n_300),
.A2(n_325),
.B1(n_333),
.B2(n_263),
.Y(n_361)
);

NAND2xp5_ASAP7_75t_L g301 ( 
.A(n_235),
.B(n_134),
.Y(n_301)
);

NAND2xp5_ASAP7_75t_L g372 ( 
.A(n_301),
.B(n_308),
.Y(n_372)
);

BUFx2_ASAP7_75t_L g387 ( 
.A(n_302),
.Y(n_387)
);

NAND2xp5_ASAP7_75t_L g308 ( 
.A(n_235),
.B(n_168),
.Y(n_308)
);

OA22x2_ASAP7_75t_L g312 ( 
.A1(n_275),
.A2(n_158),
.B1(n_200),
.B2(n_141),
.Y(n_312)
);

NAND2xp5_ASAP7_75t_L g313 ( 
.A(n_277),
.B(n_144),
.Y(n_313)
);

NAND2xp5_ASAP7_75t_L g391 ( 
.A(n_313),
.B(n_317),
.Y(n_391)
);

XOR2xp5_ASAP7_75t_L g315 ( 
.A(n_225),
.B(n_157),
.Y(n_315)
);

MAJIxp5_ASAP7_75t_L g347 ( 
.A(n_315),
.B(n_336),
.C(n_234),
.Y(n_347)
);

NAND2xp5_ASAP7_75t_L g317 ( 
.A(n_280),
.B(n_178),
.Y(n_317)
);

AOI22xp33_ASAP7_75t_SL g324 ( 
.A1(n_278),
.A2(n_171),
.B1(n_161),
.B2(n_178),
.Y(n_324)
);

AOI22xp33_ASAP7_75t_SL g358 ( 
.A1(n_324),
.A2(n_338),
.B1(n_208),
.B2(n_271),
.Y(n_358)
);

AOI22xp33_ASAP7_75t_L g326 ( 
.A1(n_225),
.A2(n_27),
.B1(n_37),
.B2(n_2),
.Y(n_326)
);

OAI22xp33_ASAP7_75t_SL g367 ( 
.A1(n_326),
.A2(n_270),
.B1(n_226),
.B2(n_216),
.Y(n_367)
);

AOI22xp33_ASAP7_75t_L g350 ( 
.A1(n_329),
.A2(n_274),
.B1(n_301),
.B2(n_266),
.Y(n_350)
);

AOI22xp5_ASAP7_75t_L g331 ( 
.A1(n_269),
.A2(n_37),
.B1(n_4),
.B2(n_5),
.Y(n_331)
);

OAI22xp5_ASAP7_75t_L g364 ( 
.A1(n_331),
.A2(n_234),
.B1(n_271),
.B2(n_215),
.Y(n_364)
);

OAI22xp5_ASAP7_75t_SL g333 ( 
.A1(n_239),
.A2(n_210),
.B1(n_211),
.B2(n_213),
.Y(n_333)
);

AOI22xp33_ASAP7_75t_SL g338 ( 
.A1(n_272),
.A2(n_11),
.B1(n_5),
.B2(n_6),
.Y(n_338)
);

NAND2xp5_ASAP7_75t_L g340 ( 
.A(n_210),
.B(n_3),
.Y(n_340)
);

NAND2xp5_ASAP7_75t_L g394 ( 
.A(n_340),
.B(n_345),
.Y(n_394)
);

NAND2xp5_ASAP7_75t_L g345 ( 
.A(n_236),
.B(n_3),
.Y(n_345)
);

XNOR2xp5_ASAP7_75t_L g440 ( 
.A(n_347),
.B(n_341),
.Y(n_440)
);

CKINVDCx16_ASAP7_75t_R g348 ( 
.A(n_303),
.Y(n_348)
);

INVx1_ASAP7_75t_L g401 ( 
.A(n_348),
.Y(n_401)
);

OAI22xp5_ASAP7_75t_SL g349 ( 
.A1(n_299),
.A2(n_253),
.B1(n_273),
.B2(n_259),
.Y(n_349)
);

AOI22xp5_ASAP7_75t_L g412 ( 
.A1(n_349),
.A2(n_361),
.B1(n_364),
.B2(n_367),
.Y(n_412)
);

AOI22xp33_ASAP7_75t_SL g422 ( 
.A1(n_350),
.A2(n_358),
.B1(n_374),
.B2(n_396),
.Y(n_422)
);

INVx3_ASAP7_75t_L g351 ( 
.A(n_285),
.Y(n_351)
);

INVx2_ASAP7_75t_L g435 ( 
.A(n_351),
.Y(n_435)
);

INVx1_ASAP7_75t_L g352 ( 
.A(n_289),
.Y(n_352)
);

INVx1_ASAP7_75t_L g403 ( 
.A(n_352),
.Y(n_403)
);

NOR2xp33_ASAP7_75t_SL g353 ( 
.A(n_283),
.B(n_206),
.Y(n_353)
);

NAND2xp5_ASAP7_75t_SL g409 ( 
.A(n_353),
.B(n_360),
.Y(n_409)
);

INVx2_ASAP7_75t_L g354 ( 
.A(n_305),
.Y(n_354)
);

INVx1_ASAP7_75t_L g410 ( 
.A(n_354),
.Y(n_410)
);

INVx1_ASAP7_75t_L g355 ( 
.A(n_289),
.Y(n_355)
);

INVx1_ASAP7_75t_L g413 ( 
.A(n_355),
.Y(n_413)
);

INVx1_ASAP7_75t_L g356 ( 
.A(n_290),
.Y(n_356)
);

INVx1_ASAP7_75t_L g423 ( 
.A(n_356),
.Y(n_423)
);

CKINVDCx14_ASAP7_75t_R g357 ( 
.A(n_345),
.Y(n_357)
);

INVx11_ASAP7_75t_L g425 ( 
.A(n_357),
.Y(n_425)
);

INVx1_ASAP7_75t_L g359 ( 
.A(n_290),
.Y(n_359)
);

INVx1_ASAP7_75t_L g424 ( 
.A(n_359),
.Y(n_424)
);

NOR2xp33_ASAP7_75t_SL g360 ( 
.A(n_334),
.B(n_232),
.Y(n_360)
);

INVx2_ASAP7_75t_L g362 ( 
.A(n_305),
.Y(n_362)
);

INVx1_ASAP7_75t_L g429 ( 
.A(n_362),
.Y(n_429)
);

CKINVDCx20_ASAP7_75t_R g363 ( 
.A(n_303),
.Y(n_363)
);

NOR2xp33_ASAP7_75t_L g421 ( 
.A(n_363),
.B(n_366),
.Y(n_421)
);

OAI21xp5_ASAP7_75t_SL g404 ( 
.A1(n_365),
.A2(n_369),
.B(n_370),
.Y(n_404)
);

INVxp67_ASAP7_75t_L g366 ( 
.A(n_342),
.Y(n_366)
);

OAI22xp33_ASAP7_75t_SL g368 ( 
.A1(n_306),
.A2(n_267),
.B1(n_224),
.B2(n_260),
.Y(n_368)
);

AOI22xp5_ASAP7_75t_L g430 ( 
.A1(n_368),
.A2(n_388),
.B1(n_392),
.B2(n_395),
.Y(n_430)
);

NAND2xp33_ASAP7_75t_SL g369 ( 
.A(n_292),
.B(n_262),
.Y(n_369)
);

AOI22xp5_ASAP7_75t_SL g370 ( 
.A1(n_308),
.A2(n_219),
.B1(n_231),
.B2(n_250),
.Y(n_370)
);

AOI22xp5_ASAP7_75t_L g371 ( 
.A1(n_300),
.A2(n_221),
.B1(n_257),
.B2(n_207),
.Y(n_371)
);

OAI22xp5_ASAP7_75t_SL g419 ( 
.A1(n_371),
.A2(n_379),
.B1(n_382),
.B2(n_346),
.Y(n_419)
);

INVx3_ASAP7_75t_L g373 ( 
.A(n_285),
.Y(n_373)
);

INVx1_ASAP7_75t_L g431 ( 
.A(n_373),
.Y(n_431)
);

AOI22xp33_ASAP7_75t_L g374 ( 
.A1(n_307),
.A2(n_343),
.B1(n_314),
.B2(n_320),
.Y(n_374)
);

NAND2xp5_ASAP7_75t_L g415 ( 
.A(n_375),
.B(n_383),
.Y(n_415)
);

MAJIxp5_ASAP7_75t_L g376 ( 
.A(n_315),
.B(n_248),
.C(n_245),
.Y(n_376)
);

MAJIxp5_ASAP7_75t_L g405 ( 
.A(n_376),
.B(n_282),
.C(n_335),
.Y(n_405)
);

CKINVDCx20_ASAP7_75t_R g378 ( 
.A(n_303),
.Y(n_378)
);

NOR2xp33_ASAP7_75t_L g427 ( 
.A(n_378),
.B(n_381),
.Y(n_427)
);

AOI22xp5_ASAP7_75t_L g379 ( 
.A1(n_313),
.A2(n_221),
.B1(n_207),
.B2(n_213),
.Y(n_379)
);

OAI21xp5_ASAP7_75t_L g380 ( 
.A1(n_291),
.A2(n_219),
.B(n_237),
.Y(n_380)
);

OAI21xp5_ASAP7_75t_SL g406 ( 
.A1(n_380),
.A2(n_384),
.B(n_389),
.Y(n_406)
);

CKINVDCx20_ASAP7_75t_R g381 ( 
.A(n_296),
.Y(n_381)
);

AOI22xp5_ASAP7_75t_L g382 ( 
.A1(n_317),
.A2(n_220),
.B1(n_258),
.B2(n_10),
.Y(n_382)
);

NOR2xp33_ASAP7_75t_L g383 ( 
.A(n_284),
.B(n_333),
.Y(n_383)
);

OAI21xp5_ASAP7_75t_L g384 ( 
.A1(n_291),
.A2(n_258),
.B(n_7),
.Y(n_384)
);

INVx3_ASAP7_75t_L g385 ( 
.A(n_321),
.Y(n_385)
);

INVx1_ASAP7_75t_L g433 ( 
.A(n_385),
.Y(n_433)
);

CKINVDCx20_ASAP7_75t_R g386 ( 
.A(n_296),
.Y(n_386)
);

NOR2xp33_ASAP7_75t_L g428 ( 
.A(n_386),
.B(n_337),
.Y(n_428)
);

OAI22xp5_ASAP7_75t_SL g388 ( 
.A1(n_325),
.A2(n_258),
.B1(n_10),
.B2(n_12),
.Y(n_388)
);

OAI21xp5_ASAP7_75t_L g389 ( 
.A1(n_331),
.A2(n_258),
.B(n_10),
.Y(n_389)
);

NOR2xp33_ASAP7_75t_L g390 ( 
.A(n_323),
.B(n_6),
.Y(n_390)
);

NAND2xp5_ASAP7_75t_L g434 ( 
.A(n_390),
.B(n_393),
.Y(n_434)
);

OAI22xp5_ASAP7_75t_L g392 ( 
.A1(n_298),
.A2(n_6),
.B1(n_10),
.B2(n_12),
.Y(n_392)
);

OAI32xp33_ASAP7_75t_L g393 ( 
.A1(n_340),
.A2(n_12),
.A3(n_13),
.B1(n_14),
.B2(n_15),
.Y(n_393)
);

OAI22xp5_ASAP7_75t_L g395 ( 
.A1(n_286),
.A2(n_15),
.B1(n_336),
.B2(n_312),
.Y(n_395)
);

AOI22xp33_ASAP7_75t_L g396 ( 
.A1(n_286),
.A2(n_295),
.B1(n_312),
.B2(n_337),
.Y(n_396)
);

AOI21xp33_ASAP7_75t_L g397 ( 
.A1(n_312),
.A2(n_286),
.B(n_282),
.Y(n_397)
);

MAJx2_ASAP7_75t_L g399 ( 
.A(n_397),
.B(n_395),
.C(n_377),
.Y(n_399)
);

INVx2_ASAP7_75t_SL g398 ( 
.A(n_321),
.Y(n_398)
);

INVx1_ASAP7_75t_L g443 ( 
.A(n_398),
.Y(n_443)
);

INVx1_ASAP7_75t_SL g469 ( 
.A(n_399),
.Y(n_469)
);

CKINVDCx20_ASAP7_75t_R g400 ( 
.A(n_353),
.Y(n_400)
);

NAND2xp5_ASAP7_75t_L g471 ( 
.A(n_400),
.B(n_411),
.Y(n_471)
);

AOI21xp5_ASAP7_75t_L g402 ( 
.A1(n_397),
.A2(n_287),
.B(n_319),
.Y(n_402)
);

OAI21xp5_ASAP7_75t_SL g470 ( 
.A1(n_402),
.A2(n_351),
.B(n_373),
.Y(n_470)
);

MAJIxp5_ASAP7_75t_L g444 ( 
.A(n_405),
.B(n_440),
.C(n_348),
.Y(n_444)
);

XNOR2xp5_ASAP7_75t_SL g407 ( 
.A(n_347),
.B(n_297),
.Y(n_407)
);

XOR2xp5_ASAP7_75t_L g467 ( 
.A(n_407),
.B(n_392),
.Y(n_467)
);

OAI21x1_ASAP7_75t_L g408 ( 
.A1(n_369),
.A2(n_330),
.B(n_294),
.Y(n_408)
);

OR2x2_ASAP7_75t_L g465 ( 
.A(n_408),
.B(n_432),
.Y(n_465)
);

CKINVDCx20_ASAP7_75t_R g411 ( 
.A(n_390),
.Y(n_411)
);

BUFx24_ASAP7_75t_SL g414 ( 
.A(n_383),
.Y(n_414)
);

NOR2xp33_ASAP7_75t_L g457 ( 
.A(n_414),
.B(n_416),
.Y(n_457)
);

AOI322xp5_ASAP7_75t_L g416 ( 
.A1(n_372),
.A2(n_322),
.A3(n_316),
.B1(n_294),
.B2(n_335),
.C1(n_304),
.C2(n_341),
.Y(n_416)
);

CKINVDCx20_ASAP7_75t_R g417 ( 
.A(n_360),
.Y(n_417)
);

NAND2xp5_ASAP7_75t_L g478 ( 
.A(n_417),
.B(n_420),
.Y(n_478)
);

CKINVDCx16_ASAP7_75t_R g418 ( 
.A(n_370),
.Y(n_418)
);

INVx1_ASAP7_75t_L g445 ( 
.A(n_418),
.Y(n_445)
);

INVx1_ASAP7_75t_L g451 ( 
.A(n_419),
.Y(n_451)
);

CKINVDCx20_ASAP7_75t_R g420 ( 
.A(n_380),
.Y(n_420)
);

CKINVDCx20_ASAP7_75t_R g426 ( 
.A(n_379),
.Y(n_426)
);

NAND2xp5_ASAP7_75t_L g479 ( 
.A(n_426),
.B(n_428),
.Y(n_479)
);

FAx1_ASAP7_75t_SL g432 ( 
.A(n_376),
.B(n_304),
.CI(n_316),
.CON(n_432),
.SN(n_432)
);

CKINVDCx20_ASAP7_75t_R g436 ( 
.A(n_381),
.Y(n_436)
);

NOR2xp33_ASAP7_75t_L g458 ( 
.A(n_436),
.B(n_327),
.Y(n_458)
);

NAND2xp5_ASAP7_75t_L g437 ( 
.A(n_391),
.B(n_346),
.Y(n_437)
);

INVx1_ASAP7_75t_L g461 ( 
.A(n_437),
.Y(n_461)
);

AOI22xp5_ASAP7_75t_L g438 ( 
.A1(n_377),
.A2(n_372),
.B1(n_361),
.B2(n_357),
.Y(n_438)
);

OAI22xp5_ASAP7_75t_L g454 ( 
.A1(n_438),
.A2(n_441),
.B1(n_386),
.B2(n_359),
.Y(n_454)
);

OAI211xp5_ASAP7_75t_SL g439 ( 
.A1(n_391),
.A2(n_287),
.B(n_327),
.C(n_339),
.Y(n_439)
);

INVx1_ASAP7_75t_L g464 ( 
.A(n_439),
.Y(n_464)
);

AOI22xp5_ASAP7_75t_L g441 ( 
.A1(n_349),
.A2(n_288),
.B1(n_322),
.B2(n_318),
.Y(n_441)
);

NAND2xp5_ASAP7_75t_SL g442 ( 
.A(n_394),
.B(n_339),
.Y(n_442)
);

NAND3xp33_ASAP7_75t_L g456 ( 
.A(n_442),
.B(n_393),
.C(n_355),
.Y(n_456)
);

MAJIxp5_ASAP7_75t_L g494 ( 
.A(n_444),
.B(n_446),
.C(n_463),
.Y(n_494)
);

MAJIxp5_ASAP7_75t_L g446 ( 
.A(n_407),
.B(n_363),
.C(n_378),
.Y(n_446)
);

CKINVDCx20_ASAP7_75t_R g447 ( 
.A(n_427),
.Y(n_447)
);

NOR2xp33_ASAP7_75t_SL g503 ( 
.A(n_447),
.B(n_400),
.Y(n_503)
);

CKINVDCx16_ASAP7_75t_R g448 ( 
.A(n_421),
.Y(n_448)
);

NOR2xp33_ASAP7_75t_L g487 ( 
.A(n_448),
.B(n_456),
.Y(n_487)
);

AOI22xp5_ASAP7_75t_L g449 ( 
.A1(n_438),
.A2(n_365),
.B1(n_364),
.B2(n_388),
.Y(n_449)
);

OAI22xp5_ASAP7_75t_SL g504 ( 
.A1(n_449),
.A2(n_483),
.B1(n_412),
.B2(n_441),
.Y(n_504)
);

OAI22xp5_ASAP7_75t_SL g450 ( 
.A1(n_420),
.A2(n_375),
.B1(n_394),
.B2(n_382),
.Y(n_450)
);

AOI22xp5_ASAP7_75t_L g518 ( 
.A1(n_450),
.A2(n_453),
.B1(n_454),
.B2(n_455),
.Y(n_518)
);

INVxp67_ASAP7_75t_L g452 ( 
.A(n_404),
.Y(n_452)
);

NAND2xp5_ASAP7_75t_L g492 ( 
.A(n_452),
.B(n_458),
.Y(n_492)
);

OAI22xp5_ASAP7_75t_SL g453 ( 
.A1(n_430),
.A2(n_389),
.B1(n_371),
.B2(n_384),
.Y(n_453)
);

OAI22xp5_ASAP7_75t_SL g455 ( 
.A1(n_430),
.A2(n_387),
.B1(n_352),
.B2(n_356),
.Y(n_455)
);

OAI21xp5_ASAP7_75t_L g459 ( 
.A1(n_402),
.A2(n_387),
.B(n_398),
.Y(n_459)
);

OAI21xp5_ASAP7_75t_SL g511 ( 
.A1(n_459),
.A2(n_470),
.B(n_477),
.Y(n_511)
);

CKINVDCx16_ASAP7_75t_R g460 ( 
.A(n_409),
.Y(n_460)
);

NOR2xp33_ASAP7_75t_L g493 ( 
.A(n_460),
.B(n_462),
.Y(n_493)
);

CKINVDCx20_ASAP7_75t_R g462 ( 
.A(n_409),
.Y(n_462)
);

MAJIxp5_ASAP7_75t_L g463 ( 
.A(n_440),
.B(n_354),
.C(n_362),
.Y(n_463)
);

XNOR2xp5_ASAP7_75t_L g466 ( 
.A(n_415),
.B(n_332),
.Y(n_466)
);

XOR2xp5_ASAP7_75t_L g506 ( 
.A(n_466),
.B(n_406),
.Y(n_506)
);

XOR2xp5_ASAP7_75t_L g490 ( 
.A(n_467),
.B(n_399),
.Y(n_490)
);

AOI22x1_ASAP7_75t_L g468 ( 
.A1(n_399),
.A2(n_387),
.B1(n_398),
.B2(n_385),
.Y(n_468)
);

NAND2xp5_ASAP7_75t_L g505 ( 
.A(n_468),
.B(n_482),
.Y(n_505)
);

AOI22xp33_ASAP7_75t_L g472 ( 
.A1(n_417),
.A2(n_288),
.B1(n_319),
.B2(n_293),
.Y(n_472)
);

INVxp67_ASAP7_75t_L g491 ( 
.A(n_472),
.Y(n_491)
);

INVx1_ASAP7_75t_L g473 ( 
.A(n_403),
.Y(n_473)
);

INVx1_ASAP7_75t_L g484 ( 
.A(n_473),
.Y(n_484)
);

OAI22xp5_ASAP7_75t_L g474 ( 
.A1(n_422),
.A2(n_293),
.B1(n_328),
.B2(n_332),
.Y(n_474)
);

INVx1_ASAP7_75t_L g495 ( 
.A(n_474),
.Y(n_495)
);

INVx1_ASAP7_75t_L g475 ( 
.A(n_403),
.Y(n_475)
);

INVx1_ASAP7_75t_L g501 ( 
.A(n_475),
.Y(n_501)
);

INVx6_ASAP7_75t_L g476 ( 
.A(n_439),
.Y(n_476)
);

CKINVDCx20_ASAP7_75t_R g488 ( 
.A(n_476),
.Y(n_488)
);

OAI21xp5_ASAP7_75t_L g477 ( 
.A1(n_404),
.A2(n_309),
.B(n_328),
.Y(n_477)
);

MAJIxp5_ASAP7_75t_L g480 ( 
.A(n_405),
.B(n_311),
.C(n_310),
.Y(n_480)
);

MAJIxp5_ASAP7_75t_L g498 ( 
.A(n_480),
.B(n_481),
.C(n_429),
.Y(n_498)
);

MAJIxp5_ASAP7_75t_L g481 ( 
.A(n_415),
.B(n_401),
.C(n_437),
.Y(n_481)
);

INVx1_ASAP7_75t_SL g482 ( 
.A(n_401),
.Y(n_482)
);

AOI22xp5_ASAP7_75t_L g483 ( 
.A1(n_434),
.A2(n_311),
.B1(n_310),
.B2(n_344),
.Y(n_483)
);

CKINVDCx16_ASAP7_75t_R g485 ( 
.A(n_478),
.Y(n_485)
);

INVx1_ASAP7_75t_L g520 ( 
.A(n_485),
.Y(n_520)
);

CKINVDCx16_ASAP7_75t_R g486 ( 
.A(n_478),
.Y(n_486)
);

INVx1_ASAP7_75t_L g532 ( 
.A(n_486),
.Y(n_532)
);

AOI22xp5_ASAP7_75t_L g489 ( 
.A1(n_451),
.A2(n_434),
.B1(n_436),
.B2(n_418),
.Y(n_489)
);

OAI22xp5_ASAP7_75t_L g519 ( 
.A1(n_489),
.A2(n_496),
.B1(n_449),
.B2(n_518),
.Y(n_519)
);

XOR2xp5_ASAP7_75t_L g526 ( 
.A(n_490),
.B(n_497),
.Y(n_526)
);

AOI22xp5_ASAP7_75t_L g496 ( 
.A1(n_451),
.A2(n_426),
.B1(n_412),
.B2(n_419),
.Y(n_496)
);

XOR2xp5_ASAP7_75t_L g497 ( 
.A(n_444),
.B(n_446),
.Y(n_497)
);

MAJIxp5_ASAP7_75t_L g522 ( 
.A(n_498),
.B(n_480),
.C(n_469),
.Y(n_522)
);

AOI21xp5_ASAP7_75t_L g499 ( 
.A1(n_452),
.A2(n_408),
.B(n_406),
.Y(n_499)
);

OAI21xp5_ASAP7_75t_L g530 ( 
.A1(n_499),
.A2(n_513),
.B(n_514),
.Y(n_530)
);

NAND2xp5_ASAP7_75t_SL g500 ( 
.A(n_462),
.B(n_442),
.Y(n_500)
);

OR2x2_ASAP7_75t_L g534 ( 
.A(n_500),
.B(n_503),
.Y(n_534)
);

INVx1_ASAP7_75t_L g502 ( 
.A(n_473),
.Y(n_502)
);

INVx1_ASAP7_75t_L g540 ( 
.A(n_502),
.Y(n_540)
);

AOI22xp5_ASAP7_75t_L g523 ( 
.A1(n_504),
.A2(n_453),
.B1(n_464),
.B2(n_455),
.Y(n_523)
);

HB1xp67_ASAP7_75t_L g521 ( 
.A(n_506),
.Y(n_521)
);

XOR2xp5_ASAP7_75t_L g507 ( 
.A(n_467),
.B(n_463),
.Y(n_507)
);

XOR2xp5_ASAP7_75t_L g542 ( 
.A(n_507),
.B(n_431),
.Y(n_542)
);

INVx1_ASAP7_75t_L g508 ( 
.A(n_475),
.Y(n_508)
);

INVx1_ASAP7_75t_L g543 ( 
.A(n_508),
.Y(n_543)
);

INVx1_ASAP7_75t_L g509 ( 
.A(n_479),
.Y(n_509)
);

INVx1_ASAP7_75t_L g547 ( 
.A(n_509),
.Y(n_547)
);

INVx1_ASAP7_75t_L g510 ( 
.A(n_479),
.Y(n_510)
);

INVx1_ASAP7_75t_L g549 ( 
.A(n_510),
.Y(n_549)
);

NAND2xp5_ASAP7_75t_L g512 ( 
.A(n_471),
.B(n_411),
.Y(n_512)
);

INVx1_ASAP7_75t_L g528 ( 
.A(n_512),
.Y(n_528)
);

OAI21xp5_ASAP7_75t_SL g513 ( 
.A1(n_465),
.A2(n_432),
.B(n_425),
.Y(n_513)
);

OAI21xp5_ASAP7_75t_SL g514 ( 
.A1(n_465),
.A2(n_432),
.B(n_425),
.Y(n_514)
);

CKINVDCx20_ASAP7_75t_R g515 ( 
.A(n_471),
.Y(n_515)
);

NAND2xp5_ASAP7_75t_L g525 ( 
.A(n_515),
.B(n_517),
.Y(n_525)
);

OAI21xp5_ASAP7_75t_L g516 ( 
.A1(n_469),
.A2(n_413),
.B(n_423),
.Y(n_516)
);

OAI21xp5_ASAP7_75t_L g546 ( 
.A1(n_516),
.A2(n_443),
.B(n_431),
.Y(n_546)
);

INVx1_ASAP7_75t_L g517 ( 
.A(n_461),
.Y(n_517)
);

AOI21xp5_ASAP7_75t_SL g565 ( 
.A1(n_519),
.A2(n_511),
.B(n_512),
.Y(n_565)
);

MAJIxp5_ASAP7_75t_L g550 ( 
.A(n_522),
.B(n_524),
.C(n_527),
.Y(n_550)
);

OAI22xp5_ASAP7_75t_L g569 ( 
.A1(n_523),
.A2(n_533),
.B1(n_495),
.B2(n_504),
.Y(n_569)
);

MAJIxp5_ASAP7_75t_L g524 ( 
.A(n_494),
.B(n_481),
.C(n_466),
.Y(n_524)
);

MAJIxp5_ASAP7_75t_L g527 ( 
.A(n_494),
.B(n_482),
.C(n_461),
.Y(n_527)
);

MAJIxp5_ASAP7_75t_L g529 ( 
.A(n_497),
.B(n_445),
.C(n_470),
.Y(n_529)
);

MAJIxp5_ASAP7_75t_L g557 ( 
.A(n_529),
.B(n_531),
.C(n_535),
.Y(n_557)
);

MAJIxp5_ASAP7_75t_L g531 ( 
.A(n_498),
.B(n_445),
.C(n_450),
.Y(n_531)
);

AOI22xp5_ASAP7_75t_L g533 ( 
.A1(n_518),
.A2(n_464),
.B1(n_459),
.B2(n_483),
.Y(n_533)
);

MAJIxp5_ASAP7_75t_L g535 ( 
.A(n_507),
.B(n_477),
.C(n_468),
.Y(n_535)
);

XNOR2xp5_ASAP7_75t_L g536 ( 
.A(n_490),
.B(n_468),
.Y(n_536)
);

XNOR2xp5_ASAP7_75t_L g553 ( 
.A(n_536),
.B(n_548),
.Y(n_553)
);

NOR2x1_ASAP7_75t_R g537 ( 
.A(n_509),
.B(n_476),
.Y(n_537)
);

INVxp67_ASAP7_75t_L g568 ( 
.A(n_537),
.Y(n_568)
);

OAI22xp5_ASAP7_75t_SL g538 ( 
.A1(n_485),
.A2(n_457),
.B1(n_424),
.B2(n_413),
.Y(n_538)
);

INVx1_ASAP7_75t_L g563 ( 
.A(n_538),
.Y(n_563)
);

MAJIxp5_ASAP7_75t_L g539 ( 
.A(n_506),
.B(n_429),
.C(n_410),
.Y(n_539)
);

MAJIxp5_ASAP7_75t_L g558 ( 
.A(n_539),
.B(n_499),
.C(n_506),
.Y(n_558)
);

OAI22xp5_ASAP7_75t_SL g541 ( 
.A1(n_486),
.A2(n_423),
.B1(n_424),
.B2(n_410),
.Y(n_541)
);

NAND2xp5_ASAP7_75t_L g551 ( 
.A(n_541),
.B(n_515),
.Y(n_551)
);

XNOR2xp5_ASAP7_75t_SL g573 ( 
.A(n_542),
.B(n_484),
.Y(n_573)
);

CKINVDCx20_ASAP7_75t_R g544 ( 
.A(n_503),
.Y(n_544)
);

OAI22xp33_ASAP7_75t_SL g555 ( 
.A1(n_544),
.A2(n_545),
.B1(n_493),
.B2(n_510),
.Y(n_555)
);

CKINVDCx20_ASAP7_75t_R g545 ( 
.A(n_493),
.Y(n_545)
);

OR2x2_ASAP7_75t_L g552 ( 
.A(n_546),
.B(n_516),
.Y(n_552)
);

XNOR2xp5_ASAP7_75t_L g548 ( 
.A(n_513),
.B(n_433),
.Y(n_548)
);

INVx1_ASAP7_75t_L g580 ( 
.A(n_551),
.Y(n_580)
);

INVx1_ASAP7_75t_L g582 ( 
.A(n_552),
.Y(n_582)
);

AOI21xp5_ASAP7_75t_L g554 ( 
.A1(n_530),
.A2(n_534),
.B(n_505),
.Y(n_554)
);

OAI21xp5_ASAP7_75t_SL g593 ( 
.A1(n_554),
.A2(n_565),
.B(n_567),
.Y(n_593)
);

INVx1_ASAP7_75t_L g590 ( 
.A(n_555),
.Y(n_590)
);

INVx1_ASAP7_75t_L g556 ( 
.A(n_534),
.Y(n_556)
);

INVx1_ASAP7_75t_L g576 ( 
.A(n_556),
.Y(n_576)
);

XNOR2xp5_ASAP7_75t_L g577 ( 
.A(n_558),
.B(n_570),
.Y(n_577)
);

INVx1_ASAP7_75t_SL g559 ( 
.A(n_546),
.Y(n_559)
);

INVx1_ASAP7_75t_L g597 ( 
.A(n_559),
.Y(n_597)
);

MAJIxp5_ASAP7_75t_L g560 ( 
.A(n_524),
.B(n_492),
.C(n_514),
.Y(n_560)
);

NAND2xp5_ASAP7_75t_SL g581 ( 
.A(n_560),
.B(n_561),
.Y(n_581)
);

MAJIxp5_ASAP7_75t_L g561 ( 
.A(n_542),
.B(n_492),
.C(n_517),
.Y(n_561)
);

MAJIxp5_ASAP7_75t_L g562 ( 
.A(n_527),
.B(n_511),
.C(n_489),
.Y(n_562)
);

NAND2xp5_ASAP7_75t_SL g592 ( 
.A(n_562),
.B(n_574),
.Y(n_592)
);

OAI22xp5_ASAP7_75t_SL g564 ( 
.A1(n_523),
.A2(n_488),
.B1(n_505),
.B2(n_496),
.Y(n_564)
);

AOI22xp33_ASAP7_75t_SL g578 ( 
.A1(n_564),
.A2(n_569),
.B1(n_571),
.B2(n_572),
.Y(n_578)
);

NAND2xp5_ASAP7_75t_L g566 ( 
.A(n_541),
.B(n_500),
.Y(n_566)
);

CKINVDCx20_ASAP7_75t_R g585 ( 
.A(n_566),
.Y(n_585)
);

OAI21xp5_ASAP7_75t_SL g567 ( 
.A1(n_530),
.A2(n_488),
.B(n_487),
.Y(n_567)
);

XNOR2xp5_ASAP7_75t_L g570 ( 
.A(n_522),
.B(n_487),
.Y(n_570)
);

OAI22xp5_ASAP7_75t_L g571 ( 
.A1(n_533),
.A2(n_495),
.B1(n_491),
.B2(n_508),
.Y(n_571)
);

INVx1_ASAP7_75t_L g572 ( 
.A(n_525),
.Y(n_572)
);

XNOR2xp5_ASAP7_75t_SL g586 ( 
.A(n_573),
.B(n_526),
.Y(n_586)
);

INVx1_ASAP7_75t_L g574 ( 
.A(n_525),
.Y(n_574)
);

OAI21xp5_ASAP7_75t_SL g575 ( 
.A1(n_528),
.A2(n_502),
.B(n_484),
.Y(n_575)
);

NAND2xp5_ASAP7_75t_SL g596 ( 
.A(n_575),
.B(n_501),
.Y(n_596)
);

OAI221xp5_ASAP7_75t_L g579 ( 
.A1(n_554),
.A2(n_549),
.B1(n_547),
.B2(n_528),
.C(n_532),
.Y(n_579)
);

INVx1_ASAP7_75t_L g607 ( 
.A(n_579),
.Y(n_607)
);

NOR2xp33_ASAP7_75t_SL g583 ( 
.A(n_570),
.B(n_538),
.Y(n_583)
);

NAND2xp5_ASAP7_75t_L g603 ( 
.A(n_583),
.B(n_588),
.Y(n_603)
);

NAND2xp5_ASAP7_75t_L g584 ( 
.A(n_566),
.B(n_520),
.Y(n_584)
);

INVx1_ASAP7_75t_L g612 ( 
.A(n_584),
.Y(n_612)
);

XNOR2xp5_ASAP7_75t_L g601 ( 
.A(n_586),
.B(n_587),
.Y(n_601)
);

XNOR2xp5_ASAP7_75t_L g587 ( 
.A(n_550),
.B(n_531),
.Y(n_587)
);

AND2x2_ASAP7_75t_L g588 ( 
.A(n_559),
.B(n_548),
.Y(n_588)
);

MAJIxp5_ASAP7_75t_L g589 ( 
.A(n_550),
.B(n_526),
.C(n_539),
.Y(n_589)
);

NAND2xp5_ASAP7_75t_L g605 ( 
.A(n_589),
.B(n_596),
.Y(n_605)
);

XNOR2xp5_ASAP7_75t_SL g591 ( 
.A(n_573),
.B(n_521),
.Y(n_591)
);

XNOR2xp5_ASAP7_75t_L g604 ( 
.A(n_591),
.B(n_594),
.Y(n_604)
);

XNOR2xp5_ASAP7_75t_L g594 ( 
.A(n_557),
.B(n_535),
.Y(n_594)
);

OAI22xp5_ASAP7_75t_SL g595 ( 
.A1(n_563),
.A2(n_537),
.B1(n_536),
.B2(n_543),
.Y(n_595)
);

AOI22xp5_ASAP7_75t_SL g602 ( 
.A1(n_595),
.A2(n_568),
.B1(n_563),
.B2(n_564),
.Y(n_602)
);

HB1xp67_ASAP7_75t_L g598 ( 
.A(n_593),
.Y(n_598)
);

NAND2xp5_ASAP7_75t_L g621 ( 
.A(n_598),
.B(n_600),
.Y(n_621)
);

XOR2xp5_ASAP7_75t_L g599 ( 
.A(n_594),
.B(n_558),
.Y(n_599)
);

XOR2xp5_ASAP7_75t_L g618 ( 
.A(n_599),
.B(n_614),
.Y(n_618)
);

NOR2xp33_ASAP7_75t_L g600 ( 
.A(n_587),
.B(n_567),
.Y(n_600)
);

OAI22xp5_ASAP7_75t_SL g623 ( 
.A1(n_602),
.A2(n_610),
.B1(n_588),
.B2(n_585),
.Y(n_623)
);

NAND2xp5_ASAP7_75t_L g606 ( 
.A(n_592),
.B(n_561),
.Y(n_606)
);

NAND2xp5_ASAP7_75t_L g625 ( 
.A(n_606),
.B(n_608),
.Y(n_625)
);

MAJIxp5_ASAP7_75t_L g608 ( 
.A(n_589),
.B(n_557),
.C(n_560),
.Y(n_608)
);

MAJIxp5_ASAP7_75t_L g609 ( 
.A(n_577),
.B(n_562),
.C(n_565),
.Y(n_609)
);

MAJIxp5_ASAP7_75t_L g620 ( 
.A(n_609),
.B(n_597),
.C(n_591),
.Y(n_620)
);

AOI22xp33_ASAP7_75t_SL g610 ( 
.A1(n_582),
.A2(n_568),
.B1(n_551),
.B2(n_552),
.Y(n_610)
);

NOR2xp33_ASAP7_75t_L g611 ( 
.A(n_590),
.B(n_575),
.Y(n_611)
);

NOR2xp33_ASAP7_75t_SL g616 ( 
.A(n_611),
.B(n_613),
.Y(n_616)
);

NOR2xp33_ASAP7_75t_L g613 ( 
.A(n_576),
.B(n_433),
.Y(n_613)
);

XNOR2xp5_ASAP7_75t_L g614 ( 
.A(n_577),
.B(n_553),
.Y(n_614)
);

XNOR2xp5_ASAP7_75t_L g615 ( 
.A(n_581),
.B(n_553),
.Y(n_615)
);

XOR2xp5_ASAP7_75t_L g619 ( 
.A(n_615),
.B(n_593),
.Y(n_619)
);

OAI22xp5_ASAP7_75t_L g617 ( 
.A1(n_607),
.A2(n_576),
.B1(n_578),
.B2(n_580),
.Y(n_617)
);

OR2x2_ASAP7_75t_L g638 ( 
.A(n_617),
.B(n_619),
.Y(n_638)
);

INVx1_ASAP7_75t_L g635 ( 
.A(n_620),
.Y(n_635)
);

MAJIxp5_ASAP7_75t_L g622 ( 
.A(n_599),
.B(n_597),
.C(n_588),
.Y(n_622)
);

NOR2xp67_ASAP7_75t_SL g637 ( 
.A(n_622),
.B(n_627),
.Y(n_637)
);

NAND2xp5_ASAP7_75t_SL g632 ( 
.A(n_623),
.B(n_624),
.Y(n_632)
);

OAI21xp5_ASAP7_75t_SL g624 ( 
.A1(n_610),
.A2(n_584),
.B(n_595),
.Y(n_624)
);

OAI22xp5_ASAP7_75t_SL g626 ( 
.A1(n_602),
.A2(n_540),
.B1(n_501),
.B2(n_586),
.Y(n_626)
);

NAND2xp5_ASAP7_75t_L g631 ( 
.A(n_626),
.B(n_628),
.Y(n_631)
);

MAJIxp5_ASAP7_75t_L g627 ( 
.A(n_608),
.B(n_529),
.C(n_443),
.Y(n_627)
);

MAJIxp5_ASAP7_75t_L g628 ( 
.A(n_609),
.B(n_435),
.C(n_344),
.Y(n_628)
);

NAND2x1_ASAP7_75t_L g629 ( 
.A(n_603),
.B(n_435),
.Y(n_629)
);

OAI21x1_ASAP7_75t_L g639 ( 
.A1(n_629),
.A2(n_601),
.B(n_619),
.Y(n_639)
);

NOR2xp33_ASAP7_75t_L g630 ( 
.A(n_616),
.B(n_605),
.Y(n_630)
);

NAND2xp5_ASAP7_75t_SL g640 ( 
.A(n_630),
.B(n_633),
.Y(n_640)
);

NAND2xp5_ASAP7_75t_L g633 ( 
.A(n_625),
.B(n_612),
.Y(n_633)
);

NOR2xp33_ASAP7_75t_L g634 ( 
.A(n_622),
.B(n_615),
.Y(n_634)
);

NAND2xp5_ASAP7_75t_SL g644 ( 
.A(n_634),
.B(n_636),
.Y(n_644)
);

NOR2xp33_ASAP7_75t_L g636 ( 
.A(n_621),
.B(n_604),
.Y(n_636)
);

AO21x1_ASAP7_75t_L g641 ( 
.A1(n_639),
.A2(n_624),
.B(n_629),
.Y(n_641)
);

INVx1_ASAP7_75t_L g648 ( 
.A(n_641),
.Y(n_648)
);

AND2x2_ASAP7_75t_L g642 ( 
.A(n_635),
.B(n_618),
.Y(n_642)
);

OAI21xp5_ASAP7_75t_L g646 ( 
.A1(n_642),
.A2(n_645),
.B(n_632),
.Y(n_646)
);

NOR2xp33_ASAP7_75t_L g643 ( 
.A(n_631),
.B(n_620),
.Y(n_643)
);

NAND2xp5_ASAP7_75t_L g647 ( 
.A(n_643),
.B(n_637),
.Y(n_647)
);

OAI21xp5_ASAP7_75t_SL g645 ( 
.A1(n_632),
.A2(n_618),
.B(n_623),
.Y(n_645)
);

AOI21xp5_ASAP7_75t_L g649 ( 
.A1(n_646),
.A2(n_647),
.B(n_644),
.Y(n_649)
);

CKINVDCx20_ASAP7_75t_R g651 ( 
.A(n_649),
.Y(n_651)
);

MAJIxp5_ASAP7_75t_L g650 ( 
.A(n_648),
.B(n_640),
.C(n_638),
.Y(n_650)
);

MAJIxp5_ASAP7_75t_L g652 ( 
.A(n_651),
.B(n_650),
.C(n_628),
.Y(n_652)
);

XOR2xp5_ASAP7_75t_L g653 ( 
.A(n_652),
.B(n_627),
.Y(n_653)
);

AOI21xp5_ASAP7_75t_L g654 ( 
.A1(n_653),
.A2(n_629),
.B(n_626),
.Y(n_654)
);


endmodule