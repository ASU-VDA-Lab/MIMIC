module fake_jpeg_16702_n_305 (n_11, n_3, n_2, n_1, n_0, n_10, n_4, n_8, n_9, n_6, n_5, n_7, n_305);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_305;

wire n_159;
wire n_117;
wire n_253;
wire n_286;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_14;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_252;
wire n_251;
wire n_273;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_279;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_278;
wire n_205;
wire n_295;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_293;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_281;
wire n_31;
wire n_155;
wire n_207;
wire n_277;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_291;
wire n_236;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_13;
wire n_175;
wire n_187;
wire n_57;
wire n_21;
wire n_223;
wire n_234;
wire n_284;
wire n_272;
wire n_288;
wire n_280;
wire n_171;
wire n_263;
wire n_23;
wire n_119;
wire n_301;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_289;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_267;
wire n_248;
wire n_30;
wire n_296;
wire n_168;
wire n_298;
wire n_106;
wire n_111;
wire n_197;
wire n_274;
wire n_186;
wire n_24;
wire n_44;
wire n_276;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_269;
wire n_122;
wire n_75;
wire n_246;
wire n_37;
wire n_233;
wire n_287;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_20;
wire n_145;
wire n_18;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_303;
wire n_90;
wire n_304;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_266;
wire n_34;
wire n_283;
wire n_107;
wire n_39;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_285;
wire n_215;
wire n_262;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_294;
wire n_299;
wire n_211;
wire n_300;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_12;
wire n_132;
wire n_133;
wire n_249;
wire n_302;
wire n_67;
wire n_271;
wire n_216;
wire n_217;
wire n_264;
wire n_184;
wire n_53;
wire n_268;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_297;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_265;
wire n_176;
wire n_199;
wire n_112;
wire n_260;
wire n_270;
wire n_222;
wire n_95;
wire n_275;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_290;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_292;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_140;
wire n_82;
wire n_128;
wire n_118;
wire n_258;
wire n_282;
wire n_96;

CKINVDCx20_ASAP7_75t_R g12 ( 
.A(n_4),
.Y(n_12)
);

BUFx12f_ASAP7_75t_L g13 ( 
.A(n_9),
.Y(n_13)
);

CKINVDCx20_ASAP7_75t_R g14 ( 
.A(n_11),
.Y(n_14)
);

BUFx12_ASAP7_75t_L g15 ( 
.A(n_9),
.Y(n_15)
);

NOR2xp33_ASAP7_75t_SL g16 ( 
.A(n_11),
.B(n_7),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_2),
.Y(n_17)
);

BUFx24_ASAP7_75t_L g18 ( 
.A(n_7),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_10),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_3),
.Y(n_20)
);

BUFx24_ASAP7_75t_L g21 ( 
.A(n_9),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_10),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_7),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_11),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_1),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_19),
.Y(n_26)
);

INVx3_ASAP7_75t_L g43 ( 
.A(n_26),
.Y(n_43)
);

INVx6_ASAP7_75t_SL g27 ( 
.A(n_13),
.Y(n_27)
);

INVx6_ASAP7_75t_SL g42 ( 
.A(n_27),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g28 ( 
.A(n_16),
.B(n_0),
.Y(n_28)
);

NOR2xp33_ASAP7_75t_SL g36 ( 
.A(n_28),
.B(n_16),
.Y(n_36)
);

BUFx12f_ASAP7_75t_L g29 ( 
.A(n_13),
.Y(n_29)
);

INVx6_ASAP7_75t_SL g44 ( 
.A(n_29),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_19),
.Y(n_30)
);

INVx3_ASAP7_75t_L g41 ( 
.A(n_30),
.Y(n_41)
);

INVx8_ASAP7_75t_L g31 ( 
.A(n_13),
.Y(n_31)
);

INVx11_ASAP7_75t_L g39 ( 
.A(n_31),
.Y(n_39)
);

INVx2_ASAP7_75t_L g32 ( 
.A(n_24),
.Y(n_32)
);

INVx3_ASAP7_75t_L g46 ( 
.A(n_32),
.Y(n_46)
);

INVx3_ASAP7_75t_L g33 ( 
.A(n_24),
.Y(n_33)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_33),
.Y(n_37)
);

BUFx3_ASAP7_75t_L g34 ( 
.A(n_13),
.Y(n_34)
);

INVx11_ASAP7_75t_L g40 ( 
.A(n_34),
.Y(n_40)
);

BUFx3_ASAP7_75t_L g35 ( 
.A(n_13),
.Y(n_35)
);

INVx8_ASAP7_75t_L g47 ( 
.A(n_35),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_SL g57 ( 
.A(n_36),
.B(n_38),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_SL g38 ( 
.A(n_28),
.B(n_17),
.Y(n_38)
);

NAND2xp5_ASAP7_75t_L g45 ( 
.A(n_26),
.B(n_13),
.Y(n_45)
);

AND2x2_ASAP7_75t_L g52 ( 
.A(n_45),
.B(n_17),
.Y(n_52)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_29),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_48),
.B(n_27),
.Y(n_58)
);

AOI22xp33_ASAP7_75t_SL g49 ( 
.A1(n_41),
.A2(n_33),
.B1(n_17),
.B2(n_32),
.Y(n_49)
);

AOI21xp5_ASAP7_75t_L g89 ( 
.A1(n_49),
.A2(n_51),
.B(n_59),
.Y(n_89)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_37),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_50),
.B(n_54),
.Y(n_78)
);

OAI21xp33_ASAP7_75t_L g51 ( 
.A1(n_45),
.A2(n_19),
.B(n_24),
.Y(n_51)
);

AND2x2_ASAP7_75t_L g82 ( 
.A(n_52),
.B(n_56),
.Y(n_82)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_46),
.Y(n_53)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_53),
.Y(n_70)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_37),
.Y(n_54)
);

AOI22xp33_ASAP7_75t_L g55 ( 
.A1(n_46),
.A2(n_33),
.B1(n_30),
.B2(n_26),
.Y(n_55)
);

AOI22xp33_ASAP7_75t_SL g75 ( 
.A1(n_55),
.A2(n_65),
.B1(n_66),
.B2(n_67),
.Y(n_75)
);

AOI22xp5_ASAP7_75t_SL g56 ( 
.A1(n_42),
.A2(n_27),
.B1(n_12),
.B2(n_31),
.Y(n_56)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_58),
.Y(n_71)
);

OAI22xp5_ASAP7_75t_L g59 ( 
.A1(n_45),
.A2(n_31),
.B1(n_30),
.B2(n_24),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_38),
.B(n_14),
.Y(n_60)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_60),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_38),
.B(n_14),
.Y(n_61)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_61),
.Y(n_79)
);

OA22x2_ASAP7_75t_SL g62 ( 
.A1(n_48),
.A2(n_29),
.B1(n_35),
.B2(n_34),
.Y(n_62)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_62),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g63 ( 
.A(n_45),
.B(n_29),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_L g73 ( 
.A(n_63),
.B(n_48),
.Y(n_73)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_46),
.Y(n_64)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_64),
.Y(n_83)
);

OAI22xp33_ASAP7_75t_L g65 ( 
.A1(n_46),
.A2(n_19),
.B1(n_12),
.B2(n_25),
.Y(n_65)
);

AOI22xp33_ASAP7_75t_L g66 ( 
.A1(n_41),
.A2(n_12),
.B1(n_25),
.B2(n_23),
.Y(n_66)
);

OAI22xp33_ASAP7_75t_L g67 ( 
.A1(n_41),
.A2(n_22),
.B1(n_20),
.B2(n_23),
.Y(n_67)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_37),
.Y(n_68)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_68),
.Y(n_87)
);

INVxp67_ASAP7_75t_L g69 ( 
.A(n_58),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_69),
.B(n_80),
.Y(n_95)
);

INVx2_ASAP7_75t_L g72 ( 
.A(n_53),
.Y(n_72)
);

INVx3_ASAP7_75t_L g90 ( 
.A(n_72),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_L g91 ( 
.A(n_73),
.B(n_74),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_SL g74 ( 
.A(n_52),
.B(n_57),
.Y(n_74)
);

INVx2_ASAP7_75t_L g77 ( 
.A(n_64),
.Y(n_77)
);

INVx3_ASAP7_75t_L g110 ( 
.A(n_77),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_60),
.B(n_61),
.Y(n_80)
);

CKINVDCx20_ASAP7_75t_R g84 ( 
.A(n_68),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_84),
.B(n_54),
.Y(n_99)
);

AND2x2_ASAP7_75t_L g85 ( 
.A(n_63),
.B(n_37),
.Y(n_85)
);

AOI22xp5_ASAP7_75t_SL g94 ( 
.A1(n_85),
.A2(n_52),
.B1(n_51),
.B2(n_50),
.Y(n_94)
);

MAJIxp5_ASAP7_75t_L g86 ( 
.A(n_63),
.B(n_48),
.C(n_29),
.Y(n_86)
);

XOR2xp5_ASAP7_75t_L g93 ( 
.A(n_86),
.B(n_52),
.Y(n_93)
);

OR2x2_ASAP7_75t_L g88 ( 
.A(n_56),
.B(n_42),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_L g97 ( 
.A(n_88),
.B(n_56),
.Y(n_97)
);

INVx8_ASAP7_75t_L g92 ( 
.A(n_72),
.Y(n_92)
);

INVx4_ASAP7_75t_L g118 ( 
.A(n_92),
.Y(n_118)
);

MAJIxp5_ASAP7_75t_L g111 ( 
.A(n_93),
.B(n_86),
.C(n_71),
.Y(n_111)
);

AND2x2_ASAP7_75t_L g134 ( 
.A(n_94),
.B(n_62),
.Y(n_134)
);

CKINVDCx20_ASAP7_75t_R g96 ( 
.A(n_78),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_SL g131 ( 
.A(n_96),
.B(n_105),
.Y(n_131)
);

OAI21xp5_ASAP7_75t_L g117 ( 
.A1(n_97),
.A2(n_102),
.B(n_82),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_L g98 ( 
.A(n_78),
.B(n_57),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g133 ( 
.A(n_98),
.B(n_101),
.Y(n_133)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_99),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_76),
.B(n_38),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_SL g115 ( 
.A(n_100),
.B(n_103),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_SL g101 ( 
.A(n_74),
.B(n_73),
.Y(n_101)
);

NAND3xp33_ASAP7_75t_L g102 ( 
.A(n_84),
.B(n_62),
.C(n_36),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_76),
.B(n_66),
.Y(n_103)
);

AOI22xp33_ASAP7_75t_SL g104 ( 
.A1(n_81),
.A2(n_44),
.B1(n_42),
.B2(n_47),
.Y(n_104)
);

AOI21xp5_ASAP7_75t_L g122 ( 
.A1(n_104),
.A2(n_43),
.B(n_41),
.Y(n_122)
);

CKINVDCx20_ASAP7_75t_R g105 ( 
.A(n_70),
.Y(n_105)
);

INVxp33_ASAP7_75t_L g106 ( 
.A(n_77),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g116 ( 
.A(n_106),
.B(n_108),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_79),
.B(n_36),
.Y(n_107)
);

INVxp33_ASAP7_75t_L g123 ( 
.A(n_107),
.Y(n_123)
);

CKINVDCx20_ASAP7_75t_R g108 ( 
.A(n_70),
.Y(n_108)
);

OA22x2_ASAP7_75t_L g109 ( 
.A1(n_89),
.A2(n_62),
.B1(n_59),
.B2(n_49),
.Y(n_109)
);

AOI22xp5_ASAP7_75t_L g125 ( 
.A1(n_109),
.A2(n_82),
.B1(n_81),
.B2(n_85),
.Y(n_125)
);

MAJIxp5_ASAP7_75t_L g137 ( 
.A(n_111),
.B(n_93),
.C(n_94),
.Y(n_137)
);

CKINVDCx20_ASAP7_75t_R g112 ( 
.A(n_99),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_L g136 ( 
.A(n_112),
.B(n_113),
.Y(n_136)
);

CKINVDCx20_ASAP7_75t_R g113 ( 
.A(n_95),
.Y(n_113)
);

CKINVDCx20_ASAP7_75t_R g114 ( 
.A(n_95),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g153 ( 
.A(n_114),
.B(n_121),
.Y(n_153)
);

OAI21xp5_ASAP7_75t_L g140 ( 
.A1(n_117),
.A2(n_122),
.B(n_124),
.Y(n_140)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_90),
.Y(n_120)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_120),
.Y(n_154)
);

CKINVDCx20_ASAP7_75t_R g121 ( 
.A(n_98),
.Y(n_121)
);

OAI21xp5_ASAP7_75t_L g124 ( 
.A1(n_97),
.A2(n_82),
.B(n_88),
.Y(n_124)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_125),
.Y(n_156)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_90),
.Y(n_126)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_126),
.Y(n_158)
);

AOI21xp5_ASAP7_75t_L g127 ( 
.A1(n_96),
.A2(n_85),
.B(n_88),
.Y(n_127)
);

OAI21xp5_ASAP7_75t_L g151 ( 
.A1(n_127),
.A2(n_134),
.B(n_87),
.Y(n_151)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_110),
.B(n_71),
.Y(n_128)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_128),
.Y(n_159)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_110),
.Y(n_129)
);

CKINVDCx16_ASAP7_75t_R g147 ( 
.A(n_129),
.Y(n_147)
);

INVx2_ASAP7_75t_SL g130 ( 
.A(n_92),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_L g149 ( 
.A(n_130),
.B(n_132),
.Y(n_149)
);

INVx6_ASAP7_75t_L g132 ( 
.A(n_92),
.Y(n_132)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_105),
.Y(n_135)
);

CKINVDCx20_ASAP7_75t_R g161 ( 
.A(n_135),
.Y(n_161)
);

NOR2xp33_ASAP7_75t_L g168 ( 
.A(n_137),
.B(n_139),
.Y(n_168)
);

XNOR2xp5_ASAP7_75t_L g138 ( 
.A(n_111),
.B(n_91),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_SL g185 ( 
.A(n_138),
.B(n_150),
.Y(n_185)
);

MAJIxp5_ASAP7_75t_L g139 ( 
.A(n_125),
.B(n_91),
.C(n_101),
.Y(n_139)
);

OR2x2_ASAP7_75t_L g141 ( 
.A(n_112),
.B(n_121),
.Y(n_141)
);

OAI21xp5_ASAP7_75t_L g172 ( 
.A1(n_141),
.A2(n_144),
.B(n_151),
.Y(n_172)
);

MAJIxp5_ASAP7_75t_L g142 ( 
.A(n_127),
.B(n_89),
.C(n_79),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_L g171 ( 
.A(n_142),
.B(n_145),
.Y(n_171)
);

NOR2xp33_ASAP7_75t_SL g143 ( 
.A(n_123),
.B(n_107),
.Y(n_143)
);

NOR2xp33_ASAP7_75t_SL g169 ( 
.A(n_143),
.B(n_103),
.Y(n_169)
);

OR2x6_ASAP7_75t_L g144 ( 
.A(n_117),
.B(n_102),
.Y(n_144)
);

MAJIxp5_ASAP7_75t_L g145 ( 
.A(n_124),
.B(n_87),
.C(n_83),
.Y(n_145)
);

HB1xp67_ASAP7_75t_L g146 ( 
.A(n_120),
.Y(n_146)
);

CKINVDCx20_ASAP7_75t_R g167 ( 
.A(n_146),
.Y(n_167)
);

HB1xp67_ASAP7_75t_L g148 ( 
.A(n_126),
.Y(n_148)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_148),
.Y(n_165)
);

INVx1_ASAP7_75t_SL g150 ( 
.A(n_134),
.Y(n_150)
);

HB1xp67_ASAP7_75t_L g152 ( 
.A(n_129),
.Y(n_152)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_152),
.Y(n_174)
);

NOR2xp33_ASAP7_75t_L g155 ( 
.A(n_113),
.B(n_108),
.Y(n_155)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_155),
.Y(n_164)
);

MAJIxp5_ASAP7_75t_L g157 ( 
.A(n_133),
.B(n_114),
.C(n_119),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_L g186 ( 
.A(n_157),
.B(n_162),
.Y(n_186)
);

XOR2xp5_ASAP7_75t_L g160 ( 
.A(n_133),
.B(n_100),
.Y(n_160)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_160),
.Y(n_175)
);

CKINVDCx5p33_ASAP7_75t_R g162 ( 
.A(n_119),
.Y(n_162)
);

INVx13_ASAP7_75t_L g163 ( 
.A(n_149),
.Y(n_163)
);

NOR2xp33_ASAP7_75t_L g192 ( 
.A(n_163),
.B(n_161),
.Y(n_192)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_136),
.Y(n_166)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_166),
.Y(n_189)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_169),
.Y(n_191)
);

NOR2xp33_ASAP7_75t_SL g170 ( 
.A(n_141),
.B(n_36),
.Y(n_170)
);

NOR2xp33_ASAP7_75t_SL g202 ( 
.A(n_170),
.B(n_182),
.Y(n_202)
);

AOI21xp5_ASAP7_75t_L g173 ( 
.A1(n_140),
.A2(n_134),
.B(n_131),
.Y(n_173)
);

OAI22xp5_ASAP7_75t_L g206 ( 
.A1(n_173),
.A2(n_44),
.B1(n_47),
.B2(n_40),
.Y(n_206)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_153),
.Y(n_176)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_176),
.Y(n_199)
);

A2O1A1O1Ixp25_ASAP7_75t_L g177 ( 
.A1(n_144),
.A2(n_115),
.B(n_109),
.C(n_135),
.D(n_122),
.Y(n_177)
);

XNOR2xp5_ASAP7_75t_SL g201 ( 
.A(n_177),
.B(n_188),
.Y(n_201)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_154),
.Y(n_178)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_178),
.Y(n_208)
);

OAI22xp5_ASAP7_75t_SL g179 ( 
.A1(n_156),
.A2(n_109),
.B1(n_116),
.B2(n_75),
.Y(n_179)
);

OAI22xp5_ASAP7_75t_SL g195 ( 
.A1(n_179),
.A2(n_181),
.B1(n_183),
.B2(n_187),
.Y(n_195)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_158),
.Y(n_180)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_180),
.Y(n_210)
);

AOI22xp5_ASAP7_75t_L g181 ( 
.A1(n_142),
.A2(n_109),
.B1(n_132),
.B2(n_118),
.Y(n_181)
);

NOR2xp33_ASAP7_75t_SL g182 ( 
.A(n_159),
.B(n_115),
.Y(n_182)
);

OAI22xp5_ASAP7_75t_SL g183 ( 
.A1(n_150),
.A2(n_109),
.B1(n_118),
.B2(n_130),
.Y(n_183)
);

INVx1_ASAP7_75t_SL g184 ( 
.A(n_162),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_L g203 ( 
.A(n_184),
.B(n_151),
.Y(n_203)
);

AOI22xp5_ASAP7_75t_L g187 ( 
.A1(n_144),
.A2(n_130),
.B1(n_83),
.B2(n_43),
.Y(n_187)
);

A2O1A1O1Ixp25_ASAP7_75t_L g188 ( 
.A1(n_144),
.A2(n_62),
.B(n_42),
.C(n_44),
.D(n_34),
.Y(n_188)
);

CKINVDCx16_ASAP7_75t_R g190 ( 
.A(n_164),
.Y(n_190)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_190),
.Y(n_220)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_192),
.Y(n_221)
);

MAJIxp5_ASAP7_75t_L g193 ( 
.A(n_168),
.B(n_138),
.C(n_137),
.Y(n_193)
);

MAJIxp5_ASAP7_75t_L g213 ( 
.A(n_193),
.B(n_205),
.C(n_207),
.Y(n_213)
);

XOR2xp5_ASAP7_75t_L g194 ( 
.A(n_185),
.B(n_140),
.Y(n_194)
);

XOR2xp5_ASAP7_75t_L g224 ( 
.A(n_194),
.B(n_204),
.Y(n_224)
);

NOR2xp33_ASAP7_75t_L g196 ( 
.A(n_167),
.B(n_160),
.Y(n_196)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_196),
.Y(n_228)
);

AOI22xp5_ASAP7_75t_L g197 ( 
.A1(n_186),
.A2(n_157),
.B1(n_144),
.B2(n_145),
.Y(n_197)
);

OAI22xp5_ASAP7_75t_L g219 ( 
.A1(n_197),
.A2(n_174),
.B1(n_165),
.B2(n_180),
.Y(n_219)
);

CKINVDCx20_ASAP7_75t_R g198 ( 
.A(n_176),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_L g218 ( 
.A(n_198),
.B(n_200),
.Y(n_218)
);

NOR2xp33_ASAP7_75t_L g200 ( 
.A(n_163),
.B(n_147),
.Y(n_200)
);

NAND2xp5_ASAP7_75t_L g222 ( 
.A(n_203),
.B(n_209),
.Y(n_222)
);

XNOR2xp5_ASAP7_75t_SL g204 ( 
.A(n_172),
.B(n_139),
.Y(n_204)
);

MAJIxp5_ASAP7_75t_L g205 ( 
.A(n_171),
.B(n_35),
.C(n_47),
.Y(n_205)
);

AOI21xp5_ASAP7_75t_L g225 ( 
.A1(n_206),
.A2(n_21),
.B(n_18),
.Y(n_225)
);

MAJIxp5_ASAP7_75t_L g207 ( 
.A(n_186),
.B(n_175),
.C(n_181),
.Y(n_207)
);

INVx1_ASAP7_75t_SL g209 ( 
.A(n_184),
.Y(n_209)
);

XNOR2x2_ASAP7_75t_SL g211 ( 
.A(n_173),
.B(n_44),
.Y(n_211)
);

OAI22xp5_ASAP7_75t_SL g215 ( 
.A1(n_211),
.A2(n_188),
.B1(n_187),
.B2(n_172),
.Y(n_215)
);

XNOR2xp5_ASAP7_75t_L g212 ( 
.A(n_204),
.B(n_183),
.Y(n_212)
);

MAJIxp5_ASAP7_75t_L g233 ( 
.A(n_212),
.B(n_223),
.C(n_226),
.Y(n_233)
);

BUFx3_ASAP7_75t_L g214 ( 
.A(n_209),
.Y(n_214)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_214),
.Y(n_237)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_215),
.Y(n_240)
);

OAI21xp5_ASAP7_75t_L g216 ( 
.A1(n_203),
.A2(n_177),
.B(n_179),
.Y(n_216)
);

AOI21xp5_ASAP7_75t_L g239 ( 
.A1(n_216),
.A2(n_230),
.B(n_218),
.Y(n_239)
);

AOI22xp5_ASAP7_75t_L g217 ( 
.A1(n_189),
.A2(n_175),
.B1(n_174),
.B2(n_165),
.Y(n_217)
);

NAND2xp5_ASAP7_75t_SL g235 ( 
.A(n_217),
.B(n_199),
.Y(n_235)
);

AOI22xp5_ASAP7_75t_L g243 ( 
.A1(n_219),
.A2(n_195),
.B1(n_201),
.B2(n_43),
.Y(n_243)
);

XNOR2xp5_ASAP7_75t_L g223 ( 
.A(n_197),
.B(n_178),
.Y(n_223)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_225),
.Y(n_248)
);

MAJIxp5_ASAP7_75t_L g226 ( 
.A(n_207),
.B(n_47),
.C(n_40),
.Y(n_226)
);

XNOR2xp5_ASAP7_75t_L g227 ( 
.A(n_193),
.B(n_47),
.Y(n_227)
);

MAJIxp5_ASAP7_75t_L g238 ( 
.A(n_227),
.B(n_231),
.C(n_208),
.Y(n_238)
);

NOR2xp33_ASAP7_75t_L g229 ( 
.A(n_202),
.B(n_15),
.Y(n_229)
);

NAND2xp5_ASAP7_75t_L g234 ( 
.A(n_229),
.B(n_221),
.Y(n_234)
);

OAI21xp5_ASAP7_75t_L g230 ( 
.A1(n_211),
.A2(n_22),
.B(n_20),
.Y(n_230)
);

MAJIxp5_ASAP7_75t_L g231 ( 
.A(n_199),
.B(n_40),
.C(n_39),
.Y(n_231)
);

NOR2xp33_ASAP7_75t_L g232 ( 
.A(n_214),
.B(n_191),
.Y(n_232)
);

NAND2xp5_ASAP7_75t_SL g254 ( 
.A(n_232),
.B(n_234),
.Y(n_254)
);

XNOR2xp5_ASAP7_75t_L g249 ( 
.A(n_235),
.B(n_236),
.Y(n_249)
);

NAND2xp5_ASAP7_75t_L g236 ( 
.A(n_222),
.B(n_210),
.Y(n_236)
);

MAJIxp5_ASAP7_75t_L g250 ( 
.A(n_238),
.B(n_242),
.C(n_244),
.Y(n_250)
);

OAI22xp5_ASAP7_75t_L g257 ( 
.A1(n_239),
.A2(n_243),
.B1(n_245),
.B2(n_39),
.Y(n_257)
);

NAND2xp5_ASAP7_75t_L g241 ( 
.A(n_220),
.B(n_205),
.Y(n_241)
);

XNOR2xp5_ASAP7_75t_L g251 ( 
.A(n_241),
.B(n_246),
.Y(n_251)
);

XNOR2xp5_ASAP7_75t_L g242 ( 
.A(n_212),
.B(n_194),
.Y(n_242)
);

MAJIxp5_ASAP7_75t_L g244 ( 
.A(n_213),
.B(n_195),
.C(n_201),
.Y(n_244)
);

NOR2xp33_ASAP7_75t_SL g245 ( 
.A(n_228),
.B(n_227),
.Y(n_245)
);

NAND2xp5_ASAP7_75t_SL g246 ( 
.A(n_223),
.B(n_40),
.Y(n_246)
);

NAND2xp5_ASAP7_75t_SL g247 ( 
.A(n_226),
.B(n_40),
.Y(n_247)
);

XNOR2xp5_ASAP7_75t_L g256 ( 
.A(n_247),
.B(n_236),
.Y(n_256)
);

MAJIxp5_ASAP7_75t_L g252 ( 
.A(n_233),
.B(n_213),
.C(n_224),
.Y(n_252)
);

MAJIxp5_ASAP7_75t_L g265 ( 
.A(n_252),
.B(n_261),
.C(n_21),
.Y(n_265)
);

AOI22xp5_ASAP7_75t_L g253 ( 
.A1(n_240),
.A2(n_231),
.B1(n_216),
.B2(n_224),
.Y(n_253)
);

OAI22xp5_ASAP7_75t_SL g272 ( 
.A1(n_253),
.A2(n_255),
.B1(n_260),
.B2(n_2),
.Y(n_272)
);

AOI22xp5_ASAP7_75t_SL g255 ( 
.A1(n_237),
.A2(n_230),
.B1(n_43),
.B2(n_55),
.Y(n_255)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_256),
.Y(n_267)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_257),
.Y(n_274)
);

XNOR2xp5_ASAP7_75t_L g258 ( 
.A(n_242),
.B(n_39),
.Y(n_258)
);

NAND2xp5_ASAP7_75t_SL g273 ( 
.A(n_258),
.B(n_259),
.Y(n_273)
);

OAI22xp5_ASAP7_75t_SL g259 ( 
.A1(n_239),
.A2(n_39),
.B1(n_43),
.B2(n_2),
.Y(n_259)
);

AOI22xp5_ASAP7_75t_L g260 ( 
.A1(n_244),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_260)
);

MAJIxp5_ASAP7_75t_L g261 ( 
.A(n_233),
.B(n_21),
.C(n_18),
.Y(n_261)
);

XNOR2xp5_ASAP7_75t_L g262 ( 
.A(n_238),
.B(n_39),
.Y(n_262)
);

NAND2xp5_ASAP7_75t_L g271 ( 
.A(n_262),
.B(n_0),
.Y(n_271)
);

XOR2xp5_ASAP7_75t_SL g263 ( 
.A(n_249),
.B(n_243),
.Y(n_263)
);

AOI21xp5_ASAP7_75t_L g278 ( 
.A1(n_263),
.A2(n_261),
.B(n_4),
.Y(n_278)
);

OAI21xp5_ASAP7_75t_L g264 ( 
.A1(n_250),
.A2(n_248),
.B(n_1),
.Y(n_264)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_264),
.Y(n_275)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_265),
.Y(n_280)
);

AOI21xp5_ASAP7_75t_L g266 ( 
.A1(n_251),
.A2(n_0),
.B(n_1),
.Y(n_266)
);

CKINVDCx20_ASAP7_75t_R g276 ( 
.A(n_266),
.Y(n_276)
);

NOR2xp33_ASAP7_75t_L g268 ( 
.A(n_254),
.B(n_15),
.Y(n_268)
);

NAND2xp5_ASAP7_75t_L g279 ( 
.A(n_268),
.B(n_3),
.Y(n_279)
);

MAJIxp5_ASAP7_75t_L g269 ( 
.A(n_250),
.B(n_21),
.C(n_18),
.Y(n_269)
);

MAJIxp5_ASAP7_75t_L g283 ( 
.A(n_269),
.B(n_270),
.C(n_18),
.Y(n_283)
);

MAJIxp5_ASAP7_75t_L g270 ( 
.A(n_252),
.B(n_21),
.C(n_18),
.Y(n_270)
);

NOR2xp33_ASAP7_75t_SL g277 ( 
.A(n_271),
.B(n_255),
.Y(n_277)
);

XOR2xp5_ASAP7_75t_L g282 ( 
.A(n_272),
.B(n_273),
.Y(n_282)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_277),
.Y(n_291)
);

XNOR2xp5_ASAP7_75t_L g289 ( 
.A(n_278),
.B(n_282),
.Y(n_289)
);

NOR2xp33_ASAP7_75t_L g288 ( 
.A(n_279),
.B(n_281),
.Y(n_288)
);

AOI22xp5_ASAP7_75t_L g281 ( 
.A1(n_274),
.A2(n_3),
.B1(n_4),
.B2(n_5),
.Y(n_281)
);

MAJIxp5_ASAP7_75t_L g285 ( 
.A(n_283),
.B(n_284),
.C(n_270),
.Y(n_285)
);

OAI22xp5_ASAP7_75t_L g284 ( 
.A1(n_267),
.A2(n_263),
.B1(n_269),
.B2(n_265),
.Y(n_284)
);

MAJIxp5_ASAP7_75t_L g294 ( 
.A(n_285),
.B(n_286),
.C(n_290),
.Y(n_294)
);

MAJIxp5_ASAP7_75t_L g286 ( 
.A(n_282),
.B(n_15),
.C(n_4),
.Y(n_286)
);

OAI21xp33_ASAP7_75t_L g287 ( 
.A1(n_275),
.A2(n_3),
.B(n_5),
.Y(n_287)
);

NAND2xp5_ASAP7_75t_L g293 ( 
.A(n_287),
.B(n_281),
.Y(n_293)
);

MAJIxp5_ASAP7_75t_L g290 ( 
.A(n_280),
.B(n_15),
.C(n_6),
.Y(n_290)
);

NOR2xp33_ASAP7_75t_L g292 ( 
.A(n_289),
.B(n_276),
.Y(n_292)
);

AOI322xp5_ASAP7_75t_L g296 ( 
.A1(n_292),
.A2(n_293),
.A3(n_295),
.B1(n_288),
.B2(n_283),
.C1(n_15),
.C2(n_8),
.Y(n_296)
);

NAND2xp5_ASAP7_75t_L g295 ( 
.A(n_288),
.B(n_291),
.Y(n_295)
);

MAJIxp5_ASAP7_75t_L g298 ( 
.A(n_296),
.B(n_297),
.C(n_5),
.Y(n_298)
);

INVx11_ASAP7_75t_L g297 ( 
.A(n_294),
.Y(n_297)
);

OAI21xp5_ASAP7_75t_SL g299 ( 
.A1(n_298),
.A2(n_5),
.B(n_6),
.Y(n_299)
);

OAI21xp5_ASAP7_75t_L g300 ( 
.A1(n_299),
.A2(n_6),
.B(n_7),
.Y(n_300)
);

MAJIxp5_ASAP7_75t_L g301 ( 
.A(n_300),
.B(n_6),
.C(n_8),
.Y(n_301)
);

MAJIxp5_ASAP7_75t_L g302 ( 
.A(n_301),
.B(n_8),
.C(n_9),
.Y(n_302)
);

CKINVDCx20_ASAP7_75t_R g303 ( 
.A(n_302),
.Y(n_303)
);

NAND2xp5_ASAP7_75t_L g304 ( 
.A(n_303),
.B(n_297),
.Y(n_304)
);

AOI22xp5_ASAP7_75t_L g305 ( 
.A1(n_304),
.A2(n_8),
.B1(n_10),
.B2(n_303),
.Y(n_305)
);


endmodule