module real_aes_6816_n_101 (n_17, n_28, n_76, n_56, n_34, n_98, n_90, n_82, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_83, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_91, n_100, n_43, n_96, n_54, n_35, n_42, n_99, n_15, n_9, n_23, n_72, n_95, n_44, n_7, n_4, n_80, n_6, n_12, n_68, n_79, n_69, n_46, n_59, n_25, n_73, n_77, n_81, n_48, n_37, n_97, n_70, n_50, n_89, n_26, n_86, n_93, n_13, n_24, n_2, n_55, n_62, n_84, n_67, n_92, n_33, n_88, n_14, n_11, n_85, n_16, n_94, n_39, n_5, n_45, n_60, n_38, n_87, n_0, n_78, n_63, n_1, n_53, n_36, n_101);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_98;
input n_90;
input n_82;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_83;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_91;
input n_100;
input n_43;
input n_96;
input n_54;
input n_35;
input n_42;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_95;
input n_44;
input n_7;
input n_4;
input n_80;
input n_6;
input n_12;
input n_68;
input n_79;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_81;
input n_48;
input n_37;
input n_97;
input n_70;
input n_50;
input n_89;
input n_26;
input n_86;
input n_93;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_84;
input n_67;
input n_92;
input n_33;
input n_88;
input n_14;
input n_11;
input n_85;
input n_16;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_87;
input n_0;
input n_78;
input n_63;
input n_1;
input n_53;
input n_36;
output n_101;
wire n_480;
wire n_113;
wire n_476;
wire n_599;
wire n_187;
wire n_436;
wire n_684;
wire n_257;
wire n_390;
wire n_185;
wire n_285;
wire n_624;
wire n_618;
wire n_522;
wire n_485;
wire n_222;
wire n_750;
wire n_631;
wire n_287;
wire n_357;
wire n_503;
wire n_635;
wire n_386;
wire n_673;
wire n_518;
wire n_254;
wire n_207;
wire n_665;
wire n_667;
wire n_577;
wire n_580;
wire n_469;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_718;
wire n_318;
wire n_355;
wire n_239;
wire n_669;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_742;
wire n_112;
wire n_319;
wire n_364;
wire n_421;
wire n_555;
wire n_329;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_169;
wire n_242;
wire n_376;
wire n_549;
wire n_571;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_752;
wire n_448;
wire n_545;
wire n_341;
wire n_556;
wire n_593;
wire n_232;
wire n_460;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_666;
wire n_320;
wire n_537;
wire n_551;
wire n_560;
wire n_260;
wire n_660;
wire n_594;
wire n_186;
wire n_138;
wire n_696;
wire n_704;
wire n_379;
wire n_374;
wire n_453;
wire n_647;
wire n_235;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_161;
wire n_189;
wire n_271;
wire n_489;
wire n_427;
wire n_548;
wire n_678;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_519;
wire n_564;
wire n_638;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_512;
wire n_395;
wire n_332;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_116;
wire n_625;
wire n_462;
wire n_289;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_716;
wire n_213;
wire n_356;
wire n_478;
wire n_584;
wire n_408;
wire n_553;
wire n_184;
wire n_372;
wire n_528;
wire n_578;
wire n_202;
wire n_495;
wire n_370;
wire n_744;
wire n_384;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_467;
wire n_327;
wire n_106;
wire n_466;
wire n_559;
wire n_636;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_726;
wire n_369;
wire n_343;
wire n_517;
wire n_683;
wire n_174;
wire n_570;
wire n_675;
wire n_530;
wire n_104;
wire n_535;
wire n_732;
wire n_211;
wire n_281;
wire n_496;
wire n_693;
wire n_173;
wire n_468;
wire n_234;
wire n_746;
wire n_284;
wire n_153;
wire n_316;
wire n_532;
wire n_656;
wire n_178;
wire n_409;
wire n_748;
wire n_523;
wire n_298;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_297;
wire n_383;
wire n_529;
wire n_119;
wire n_725;
wire n_310;
wire n_455;
wire n_504;
wire n_164;
wire n_671;
wire n_231;
wire n_102;
wire n_547;
wire n_659;
wire n_682;
wire n_634;
wire n_454;
wire n_122;
wire n_443;
wire n_565;
wire n_608;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_267;
wire n_218;
wire n_737;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_722;
wire n_745;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_331;
wire n_449;
wire n_182;
wire n_363;
wire n_417;
wire n_607;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_142;
wire n_561;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_655;
wire n_654;
wire n_527;
wire n_434;
wire n_502;
wire n_505;
wire n_600;
wire n_731;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_602;
wire n_402;
wire n_552;
wire n_617;
wire n_733;
wire n_171;
wire n_676;
wire n_658;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_146;
wire n_432;
wire n_226;
wire n_255;
wire n_286;
wire n_416;
wire n_410;
wire n_120;
wire n_751;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_695;
wire n_685;
wire n_165;
wire n_361;
wire n_632;
wire n_246;
wire n_176;
wire n_412;
wire n_163;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_501;
wire n_488;
wire n_251;
wire n_642;
wire n_613;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_702;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_734;
wire n_110;
wire n_392;
wire n_562;
wire n_150;
wire n_147;
wire n_288;
wire n_404;
wire n_598;
wire n_713;
wire n_728;
wire n_735;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_569;
wire n_563;
wire n_188;
wire n_269;
wire n_430;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_193;
wire n_397;
wire n_293;
wire n_749;
wire n_162;
wire n_385;
wire n_275;
wire n_214;
wire n_358;
wire n_649;
wire n_663;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_707;
wire n_622;
wire n_470;
wire n_133;
wire n_494;
wire n_711;
wire n_377;
wire n_273;
wire n_723;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_265;
wire n_354;
wire n_720;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_730;
wire n_643;
wire n_747;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_481;
wire n_148;
wire n_498;
wire n_691;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_233;
wire n_487;
wire n_290;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_155;
wire n_243;
wire n_692;
wire n_544;
wire n_268;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_738;
wire n_701;
wire n_309;
wire n_344;
wire n_107;
wire n_229;
wire n_482;
wire n_520;
wire n_633;
wire n_679;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_262;
wire n_630;
wire n_689;
wire n_715;
wire n_134;
wire n_349;
wire n_336;
wire n_420;
wire n_612;
wire n_195;
wire n_438;
wire n_300;
wire n_753;
wire n_252;
wire n_283;
wire n_314;
wire n_741;
wire n_249;
wire n_623;
wire n_446;
wire n_721;
wire n_221;
wire n_681;
wire n_156;
wire n_359;
wire n_717;
wire n_456;
wire n_312;
wire n_183;
wire n_266;
wire n_712;
wire n_205;
wire n_433;
wire n_516;
wire n_177;
wire n_335;
wire n_313;
wire n_627;
wire n_739;
wire n_140;
wire n_521;
wire n_418;
wire n_422;
wire n_524;
wire n_219;
wire n_705;
wire n_180;
wire n_212;
wire n_210;
wire n_575;
wire n_325;
wire n_338;
wire n_479;
wire n_442;
wire n_698;
wire n_371;
wire n_740;
wire n_103;
wire n_166;
wire n_541;
wire n_224;
wire n_151;
wire n_546;
wire n_587;
wire n_639;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_724;
wire n_440;
wire n_525;
wire n_674;
wire n_644;
wire n_152;
wire n_198;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_414;
wire n_123;
wire n_279;
wire n_686;
wire n_543;
wire n_497;
wire n_514;
wire n_507;
wire n_270;
wire n_614;
wire n_305;
wire n_586;
wire n_450;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_465;
wire n_473;
wire n_719;
wire n_566;
wire n_474;
wire n_170;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_168;
wire n_729;
wire n_241;
wire n_175;
wire n_687;
wire n_646;
wire n_650;
wire n_710;
wire n_743;
wire n_105;
wire n_294;
wire n_393;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_307;
wire n_500;
wire n_601;
wire n_661;
wire n_463;
wire n_396;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_143;
wire n_192;
wire n_475;
wire n_554;
wire n_264;
wire n_237;
wire n_668;
A2O1A1Ixp33_ASAP7_75t_SL g512 ( .A1(n_0), .A2(n_155), .B(n_513), .C(n_514), .Y(n_512) );
NAND2xp5_ASAP7_75t_L g516 ( .A(n_1), .B(n_174), .Y(n_516) );
INVx1_ASAP7_75t_L g110 ( .A(n_2), .Y(n_110) );
A2O1A1Ixp33_ASAP7_75t_L g183 ( .A1(n_3), .A2(n_141), .B(n_146), .C(n_184), .Y(n_183) );
AOI21xp5_ASAP7_75t_L g232 ( .A1(n_4), .A2(n_136), .B(n_233), .Y(n_232) );
NAND2xp5_ASAP7_75t_SL g503 ( .A(n_5), .B(n_211), .Y(n_503) );
AOI21xp5_ASAP7_75t_L g457 ( .A1(n_6), .A2(n_136), .B(n_458), .Y(n_457) );
NAND2xp5_ASAP7_75t_L g240 ( .A(n_7), .B(n_174), .Y(n_240) );
AO21x2_ASAP7_75t_L g466 ( .A1(n_8), .A2(n_159), .B(n_467), .Y(n_466) );
AND2x6_ASAP7_75t_L g141 ( .A(n_9), .B(n_142), .Y(n_141) );
A2O1A1Ixp33_ASAP7_75t_L g523 ( .A1(n_10), .A2(n_141), .B(n_146), .C(n_524), .Y(n_523) );
INVx1_ASAP7_75t_L g153 ( .A(n_11), .Y(n_153) );
NAND2xp5_ASAP7_75t_L g107 ( .A(n_12), .B(n_42), .Y(n_107) );
NOR2xp33_ASAP7_75t_L g123 ( .A(n_12), .B(n_42), .Y(n_123) );
NAND2xp5_ASAP7_75t_SL g188 ( .A(n_13), .B(n_151), .Y(n_188) );
INVx1_ASAP7_75t_L g134 ( .A(n_14), .Y(n_134) );
NAND2xp5_ASAP7_75t_SL g473 ( .A(n_15), .B(n_211), .Y(n_473) );
A2O1A1Ixp33_ASAP7_75t_L g167 ( .A1(n_16), .A2(n_154), .B(n_168), .C(n_172), .Y(n_167) );
NAND2xp5_ASAP7_75t_L g173 ( .A(n_17), .B(n_174), .Y(n_173) );
CKINVDCx20_ASAP7_75t_R g735 ( .A(n_18), .Y(n_735) );
NAND2xp5_ASAP7_75t_L g279 ( .A(n_19), .B(n_280), .Y(n_279) );
A2O1A1Ixp33_ASAP7_75t_L g197 ( .A1(n_20), .A2(n_198), .B(n_199), .C(n_201), .Y(n_197) );
A2O1A1Ixp33_ASAP7_75t_L g491 ( .A1(n_21), .A2(n_146), .B(n_215), .C(n_492), .Y(n_491) );
NAND2xp5_ASAP7_75t_SL g226 ( .A(n_22), .B(n_151), .Y(n_226) );
NAND2xp5_ASAP7_75t_SL g212 ( .A(n_23), .B(n_151), .Y(n_212) );
CKINVDCx16_ASAP7_75t_R g222 ( .A(n_24), .Y(n_222) );
INVx1_ASAP7_75t_L g210 ( .A(n_25), .Y(n_210) );
A2O1A1Ixp33_ASAP7_75t_L g469 ( .A1(n_26), .A2(n_146), .B(n_215), .C(n_470), .Y(n_469) );
BUFx6f_ASAP7_75t_L g140 ( .A(n_27), .Y(n_140) );
CKINVDCx20_ASAP7_75t_R g181 ( .A(n_28), .Y(n_181) );
AOI22xp33_ASAP7_75t_L g101 ( .A1(n_29), .A2(n_102), .B1(n_115), .B2(n_753), .Y(n_101) );
INVx1_ASAP7_75t_L g276 ( .A(n_30), .Y(n_276) );
AOI21xp5_ASAP7_75t_L g509 ( .A1(n_31), .A2(n_136), .B(n_510), .Y(n_509) );
INVx2_ASAP7_75t_L g139 ( .A(n_32), .Y(n_139) );
A2O1A1Ixp33_ASAP7_75t_L g481 ( .A1(n_33), .A2(n_227), .B(n_448), .C(n_482), .Y(n_481) );
CKINVDCx20_ASAP7_75t_R g191 ( .A(n_34), .Y(n_191) );
A2O1A1Ixp33_ASAP7_75t_L g235 ( .A1(n_35), .A2(n_198), .B(n_236), .C(n_238), .Y(n_235) );
INVxp67_ASAP7_75t_L g277 ( .A(n_36), .Y(n_277) );
NAND2xp5_ASAP7_75t_L g471 ( .A(n_37), .B(n_472), .Y(n_471) );
A2O1A1Ixp33_ASAP7_75t_L g208 ( .A1(n_38), .A2(n_146), .B(n_209), .C(n_215), .Y(n_208) );
CKINVDCx14_ASAP7_75t_R g234 ( .A(n_39), .Y(n_234) );
OAI22xp5_ASAP7_75t_SL g742 ( .A1(n_40), .A2(n_47), .B1(n_743), .B2(n_744), .Y(n_742) );
INVx1_ASAP7_75t_L g743 ( .A(n_40), .Y(n_743) );
OAI22xp5_ASAP7_75t_L g726 ( .A1(n_41), .A2(n_46), .B1(n_727), .B2(n_728), .Y(n_726) );
INVx1_ASAP7_75t_L g728 ( .A(n_41), .Y(n_728) );
A2O1A1Ixp33_ASAP7_75t_L g149 ( .A1(n_43), .A2(n_150), .B(n_152), .C(n_155), .Y(n_149) );
NAND2xp5_ASAP7_75t_L g490 ( .A(n_44), .B(n_271), .Y(n_490) );
CKINVDCx20_ASAP7_75t_R g528 ( .A(n_45), .Y(n_528) );
CKINVDCx20_ASAP7_75t_R g727 ( .A(n_46), .Y(n_727) );
INVx1_ASAP7_75t_L g744 ( .A(n_47), .Y(n_744) );
NAND2xp5_ASAP7_75t_L g451 ( .A(n_48), .B(n_211), .Y(n_451) );
CKINVDCx20_ASAP7_75t_R g750 ( .A(n_49), .Y(n_750) );
NAND2xp5_ASAP7_75t_L g468 ( .A(n_50), .B(n_136), .Y(n_468) );
CKINVDCx20_ASAP7_75t_R g217 ( .A(n_51), .Y(n_217) );
CKINVDCx20_ASAP7_75t_R g273 ( .A(n_52), .Y(n_273) );
A2O1A1Ixp33_ASAP7_75t_L g447 ( .A1(n_53), .A2(n_227), .B(n_448), .C(n_449), .Y(n_447) );
INVx1_ASAP7_75t_L g515 ( .A(n_54), .Y(n_515) );
INVx1_ASAP7_75t_L g450 ( .A(n_55), .Y(n_450) );
INVx1_ASAP7_75t_L g196 ( .A(n_56), .Y(n_196) );
NAND2xp5_ASAP7_75t_L g446 ( .A(n_57), .B(n_136), .Y(n_446) );
CKINVDCx20_ASAP7_75t_R g496 ( .A(n_58), .Y(n_496) );
CKINVDCx14_ASAP7_75t_R g144 ( .A(n_59), .Y(n_144) );
INVx1_ASAP7_75t_L g142 ( .A(n_60), .Y(n_142) );
NAND2xp5_ASAP7_75t_L g505 ( .A(n_61), .B(n_136), .Y(n_505) );
NAND2xp5_ASAP7_75t_L g464 ( .A(n_62), .B(n_174), .Y(n_464) );
A2O1A1Ixp33_ASAP7_75t_L g460 ( .A1(n_63), .A2(n_214), .B(n_461), .C(n_462), .Y(n_460) );
INVx1_ASAP7_75t_L g133 ( .A(n_64), .Y(n_133) );
INVx1_ASAP7_75t_SL g237 ( .A(n_65), .Y(n_237) );
CKINVDCx20_ASAP7_75t_R g738 ( .A(n_66), .Y(n_738) );
NAND2xp5_ASAP7_75t_SL g484 ( .A(n_67), .B(n_211), .Y(n_484) );
NAND2xp5_ASAP7_75t_L g203 ( .A(n_68), .B(n_174), .Y(n_203) );
NAND2xp5_ASAP7_75t_L g525 ( .A(n_69), .B(n_154), .Y(n_525) );
INVx1_ASAP7_75t_L g225 ( .A(n_70), .Y(n_225) );
CKINVDCx16_ASAP7_75t_R g511 ( .A(n_71), .Y(n_511) );
NAND2xp5_ASAP7_75t_L g493 ( .A(n_72), .B(n_187), .Y(n_493) );
A2O1A1Ixp33_ASAP7_75t_L g500 ( .A1(n_73), .A2(n_146), .B(n_227), .C(n_501), .Y(n_500) );
CKINVDCx16_ASAP7_75t_R g459 ( .A(n_74), .Y(n_459) );
INVx1_ASAP7_75t_L g114 ( .A(n_75), .Y(n_114) );
AOI21xp5_ASAP7_75t_L g135 ( .A1(n_76), .A2(n_136), .B(n_143), .Y(n_135) );
CKINVDCx20_ASAP7_75t_R g229 ( .A(n_77), .Y(n_229) );
AOI21xp5_ASAP7_75t_L g164 ( .A1(n_78), .A2(n_136), .B(n_165), .Y(n_164) );
AOI21xp5_ASAP7_75t_L g270 ( .A1(n_79), .A2(n_271), .B(n_272), .Y(n_270) );
INVx1_ASAP7_75t_L g166 ( .A(n_80), .Y(n_166) );
CKINVDCx16_ASAP7_75t_R g207 ( .A(n_81), .Y(n_207) );
NAND2xp5_ASAP7_75t_SL g494 ( .A(n_82), .B(n_186), .Y(n_494) );
CKINVDCx20_ASAP7_75t_R g486 ( .A(n_83), .Y(n_486) );
AOI21xp5_ASAP7_75t_L g194 ( .A1(n_84), .A2(n_136), .B(n_195), .Y(n_194) );
INVx1_ASAP7_75t_L g169 ( .A(n_85), .Y(n_169) );
INVx2_ASAP7_75t_L g131 ( .A(n_86), .Y(n_131) );
INVx1_ASAP7_75t_L g185 ( .A(n_87), .Y(n_185) );
CKINVDCx20_ASAP7_75t_R g507 ( .A(n_88), .Y(n_507) );
NAND2xp5_ASAP7_75t_SL g526 ( .A(n_89), .B(n_151), .Y(n_526) );
INVx2_ASAP7_75t_L g111 ( .A(n_90), .Y(n_111) );
OR2x2_ASAP7_75t_L g439 ( .A(n_90), .B(n_122), .Y(n_439) );
OR2x2_ASAP7_75t_L g746 ( .A(n_90), .B(n_734), .Y(n_746) );
A2O1A1Ixp33_ASAP7_75t_L g223 ( .A1(n_91), .A2(n_146), .B(n_224), .C(n_227), .Y(n_223) );
NAND2xp5_ASAP7_75t_L g480 ( .A(n_92), .B(n_136), .Y(n_480) );
INVx1_ASAP7_75t_L g483 ( .A(n_93), .Y(n_483) );
INVxp67_ASAP7_75t_L g463 ( .A(n_94), .Y(n_463) );
NAND2xp5_ASAP7_75t_L g158 ( .A(n_95), .B(n_159), .Y(n_158) );
NAND2xp5_ASAP7_75t_L g113 ( .A(n_96), .B(n_114), .Y(n_113) );
INVx2_ASAP7_75t_L g200 ( .A(n_97), .Y(n_200) );
INVx1_ASAP7_75t_L g502 ( .A(n_98), .Y(n_502) );
INVx1_ASAP7_75t_L g522 ( .A(n_99), .Y(n_522) );
AND2x2_ASAP7_75t_L g453 ( .A(n_100), .B(n_130), .Y(n_453) );
INVx1_ASAP7_75t_SL g102 ( .A(n_103), .Y(n_102) );
INVx1_ASAP7_75t_L g103 ( .A(n_104), .Y(n_103) );
INVx2_ASAP7_75t_L g753 ( .A(n_104), .Y(n_753) );
CKINVDCx9p33_ASAP7_75t_R g104 ( .A(n_105), .Y(n_104) );
NAND2xp5_ASAP7_75t_L g105 ( .A(n_106), .B(n_108), .Y(n_105) );
CKINVDCx20_ASAP7_75t_R g106 ( .A(n_107), .Y(n_106) );
CKINVDCx14_ASAP7_75t_R g108 ( .A(n_109), .Y(n_108) );
NAND3xp33_ASAP7_75t_SL g109 ( .A(n_110), .B(n_111), .C(n_112), .Y(n_109) );
AND2x2_ASAP7_75t_L g122 ( .A(n_110), .B(n_123), .Y(n_122) );
OR2x2_ASAP7_75t_L g121 ( .A(n_111), .B(n_122), .Y(n_121) );
NOR2x2_ASAP7_75t_L g733 ( .A(n_111), .B(n_734), .Y(n_733) );
INVx1_ASAP7_75t_SL g112 ( .A(n_113), .Y(n_112) );
AO221x1_ASAP7_75t_L g115 ( .A1(n_116), .A2(n_736), .B1(n_739), .B2(n_747), .C(n_749), .Y(n_115) );
OAI222xp33_ASAP7_75t_L g116 ( .A1(n_117), .A2(n_725), .B1(n_726), .B2(n_729), .C1(n_732), .C2(n_735), .Y(n_116) );
AOI22xp5_ASAP7_75t_L g117 ( .A1(n_118), .A2(n_124), .B1(n_436), .B2(n_440), .Y(n_117) );
AOI22x1_ASAP7_75t_SL g729 ( .A1(n_118), .A2(n_436), .B1(n_730), .B2(n_731), .Y(n_729) );
INVx1_ASAP7_75t_L g118 ( .A(n_119), .Y(n_118) );
INVx2_ASAP7_75t_L g119 ( .A(n_120), .Y(n_119) );
INVx1_ASAP7_75t_L g120 ( .A(n_121), .Y(n_120) );
INVx2_ASAP7_75t_L g734 ( .A(n_122), .Y(n_734) );
INVx2_ASAP7_75t_L g730 ( .A(n_124), .Y(n_730) );
OR2x2_ASAP7_75t_L g124 ( .A(n_125), .B(n_366), .Y(n_124) );
NAND5xp2_ASAP7_75t_L g125 ( .A(n_126), .B(n_281), .C(n_313), .D(n_330), .E(n_353), .Y(n_125) );
AOI221xp5_ASAP7_75t_L g126 ( .A1(n_127), .A2(n_204), .B1(n_241), .B2(n_245), .C(n_249), .Y(n_126) );
INVx1_ASAP7_75t_L g393 ( .A(n_127), .Y(n_393) );
AND2x2_ASAP7_75t_L g127 ( .A(n_128), .B(n_176), .Y(n_127) );
AND3x2_ASAP7_75t_L g368 ( .A(n_128), .B(n_178), .C(n_369), .Y(n_368) );
AND2x2_ASAP7_75t_L g128 ( .A(n_129), .B(n_161), .Y(n_128) );
NAND2xp5_ASAP7_75t_L g246 ( .A(n_129), .B(n_247), .Y(n_246) );
BUFx3_ASAP7_75t_L g256 ( .A(n_129), .Y(n_256) );
AND2x2_ASAP7_75t_L g260 ( .A(n_129), .B(n_192), .Y(n_260) );
INVx2_ASAP7_75t_L g290 ( .A(n_129), .Y(n_290) );
OR2x2_ASAP7_75t_L g301 ( .A(n_129), .B(n_193), .Y(n_301) );
NOR2xp33_ASAP7_75t_L g320 ( .A(n_129), .B(n_177), .Y(n_320) );
NAND2xp5_ASAP7_75t_L g338 ( .A(n_129), .B(n_339), .Y(n_338) );
AND2x2_ASAP7_75t_L g380 ( .A(n_129), .B(n_193), .Y(n_380) );
OA21x2_ASAP7_75t_L g129 ( .A1(n_130), .A2(n_135), .B(n_158), .Y(n_129) );
INVx1_ASAP7_75t_L g179 ( .A(n_130), .Y(n_179) );
O2A1O1Ixp33_ASAP7_75t_L g206 ( .A1(n_130), .A2(n_182), .B(n_207), .C(n_208), .Y(n_206) );
INVx2_ASAP7_75t_L g230 ( .A(n_130), .Y(n_230) );
AOI21xp5_ASAP7_75t_L g445 ( .A1(n_130), .A2(n_446), .B(n_447), .Y(n_445) );
AOI21xp5_ASAP7_75t_L g479 ( .A1(n_130), .A2(n_480), .B(n_481), .Y(n_479) );
AND2x2_ASAP7_75t_SL g130 ( .A(n_131), .B(n_132), .Y(n_130) );
AND2x2_ASAP7_75t_L g160 ( .A(n_131), .B(n_132), .Y(n_160) );
NAND2xp5_ASAP7_75t_L g132 ( .A(n_133), .B(n_134), .Y(n_132) );
BUFx2_ASAP7_75t_L g271 ( .A(n_136), .Y(n_271) );
AND2x4_ASAP7_75t_L g136 ( .A(n_137), .B(n_141), .Y(n_136) );
NAND2x1p5_ASAP7_75t_L g182 ( .A(n_137), .B(n_141), .Y(n_182) );
AND2x2_ASAP7_75t_L g137 ( .A(n_138), .B(n_140), .Y(n_137) );
INVx1_ASAP7_75t_L g214 ( .A(n_138), .Y(n_214) );
INVx1_ASAP7_75t_L g138 ( .A(n_139), .Y(n_138) );
INVx2_ASAP7_75t_L g147 ( .A(n_139), .Y(n_147) );
INVx1_ASAP7_75t_L g202 ( .A(n_139), .Y(n_202) );
INVx1_ASAP7_75t_L g148 ( .A(n_140), .Y(n_148) );
BUFx6f_ASAP7_75t_L g151 ( .A(n_140), .Y(n_151) );
INVx3_ASAP7_75t_L g154 ( .A(n_140), .Y(n_154) );
BUFx6f_ASAP7_75t_L g171 ( .A(n_140), .Y(n_171) );
INVx1_ASAP7_75t_L g472 ( .A(n_140), .Y(n_472) );
INVx4_ASAP7_75t_SL g157 ( .A(n_141), .Y(n_157) );
BUFx3_ASAP7_75t_L g215 ( .A(n_141), .Y(n_215) );
O2A1O1Ixp33_ASAP7_75t_SL g143 ( .A1(n_144), .A2(n_145), .B(n_149), .C(n_157), .Y(n_143) );
O2A1O1Ixp33_ASAP7_75t_SL g165 ( .A1(n_145), .A2(n_157), .B(n_166), .C(n_167), .Y(n_165) );
O2A1O1Ixp33_ASAP7_75t_SL g195 ( .A1(n_145), .A2(n_157), .B(n_196), .C(n_197), .Y(n_195) );
O2A1O1Ixp33_ASAP7_75t_L g233 ( .A1(n_145), .A2(n_157), .B(n_234), .C(n_235), .Y(n_233) );
O2A1O1Ixp33_ASAP7_75t_SL g272 ( .A1(n_145), .A2(n_157), .B(n_273), .C(n_274), .Y(n_272) );
INVx2_ASAP7_75t_L g448 ( .A(n_145), .Y(n_448) );
O2A1O1Ixp33_ASAP7_75t_L g458 ( .A1(n_145), .A2(n_157), .B(n_459), .C(n_460), .Y(n_458) );
O2A1O1Ixp33_ASAP7_75t_SL g510 ( .A1(n_145), .A2(n_157), .B(n_511), .C(n_512), .Y(n_510) );
INVx5_ASAP7_75t_L g145 ( .A(n_146), .Y(n_145) );
AND2x6_ASAP7_75t_L g146 ( .A(n_147), .B(n_148), .Y(n_146) );
BUFx3_ASAP7_75t_L g156 ( .A(n_147), .Y(n_156) );
BUFx6f_ASAP7_75t_L g239 ( .A(n_147), .Y(n_239) );
INVx2_ASAP7_75t_L g150 ( .A(n_151), .Y(n_150) );
INVx4_ASAP7_75t_L g198 ( .A(n_151), .Y(n_198) );
NOR2xp33_ASAP7_75t_L g152 ( .A(n_153), .B(n_154), .Y(n_152) );
INVx5_ASAP7_75t_L g211 ( .A(n_154), .Y(n_211) );
INVx2_ASAP7_75t_L g189 ( .A(n_155), .Y(n_189) );
INVx2_ASAP7_75t_L g155 ( .A(n_156), .Y(n_155) );
INVx1_ASAP7_75t_L g172 ( .A(n_156), .Y(n_172) );
HB1xp67_ASAP7_75t_L g452 ( .A(n_156), .Y(n_452) );
INVx1_ASAP7_75t_L g227 ( .A(n_157), .Y(n_227) );
HB1xp67_ASAP7_75t_L g163 ( .A(n_159), .Y(n_163) );
INVx4_ASAP7_75t_L g175 ( .A(n_159), .Y(n_175) );
AOI21xp5_ASAP7_75t_L g467 ( .A1(n_159), .A2(n_468), .B(n_469), .Y(n_467) );
BUFx6f_ASAP7_75t_L g159 ( .A(n_160), .Y(n_159) );
INVx1_ASAP7_75t_L g268 ( .A(n_160), .Y(n_268) );
HB1xp67_ASAP7_75t_L g259 ( .A(n_161), .Y(n_259) );
AND2x2_ASAP7_75t_L g321 ( .A(n_161), .B(n_322), .Y(n_321) );
NAND2xp5_ASAP7_75t_L g340 ( .A(n_161), .B(n_177), .Y(n_340) );
INVx1_ASAP7_75t_SL g161 ( .A(n_162), .Y(n_161) );
OR2x2_ASAP7_75t_L g248 ( .A(n_162), .B(n_177), .Y(n_248) );
HB1xp67_ASAP7_75t_L g255 ( .A(n_162), .Y(n_255) );
AND2x2_ASAP7_75t_L g307 ( .A(n_162), .B(n_193), .Y(n_307) );
NAND3xp33_ASAP7_75t_L g332 ( .A(n_162), .B(n_176), .C(n_290), .Y(n_332) );
AND2x2_ASAP7_75t_L g397 ( .A(n_162), .B(n_178), .Y(n_397) );
AND2x2_ASAP7_75t_L g431 ( .A(n_162), .B(n_177), .Y(n_431) );
OA21x2_ASAP7_75t_L g162 ( .A1(n_163), .A2(n_164), .B(n_173), .Y(n_162) );
OA21x2_ASAP7_75t_L g193 ( .A1(n_163), .A2(n_194), .B(n_203), .Y(n_193) );
OA21x2_ASAP7_75t_L g231 ( .A1(n_163), .A2(n_232), .B(n_240), .Y(n_231) );
OA21x2_ASAP7_75t_L g456 ( .A1(n_163), .A2(n_457), .B(n_464), .Y(n_456) );
NOR2xp33_ASAP7_75t_L g168 ( .A(n_169), .B(n_170), .Y(n_168) );
NOR2xp33_ASAP7_75t_L g199 ( .A(n_170), .B(n_200), .Y(n_199) );
OAI22xp33_ASAP7_75t_L g275 ( .A1(n_170), .A2(n_211), .B1(n_276), .B2(n_277), .Y(n_275) );
INVx1_ASAP7_75t_L g461 ( .A(n_170), .Y(n_461) );
INVx4_ASAP7_75t_L g170 ( .A(n_171), .Y(n_170) );
INVx2_ASAP7_75t_L g187 ( .A(n_171), .Y(n_187) );
OA21x2_ASAP7_75t_L g508 ( .A1(n_174), .A2(n_509), .B(n_516), .Y(n_508) );
INVx3_ASAP7_75t_L g174 ( .A(n_175), .Y(n_174) );
NOR2xp33_ASAP7_75t_L g190 ( .A(n_175), .B(n_191), .Y(n_190) );
NOR2xp33_ASAP7_75t_L g216 ( .A(n_175), .B(n_217), .Y(n_216) );
AO21x2_ASAP7_75t_L g220 ( .A1(n_175), .A2(n_221), .B(n_228), .Y(n_220) );
NOR2xp33_ASAP7_75t_L g485 ( .A(n_175), .B(n_486), .Y(n_485) );
AO21x2_ASAP7_75t_L g498 ( .A1(n_175), .A2(n_499), .B(n_506), .Y(n_498) );
NOR2xp33_ASAP7_75t_L g506 ( .A(n_175), .B(n_507), .Y(n_506) );
AO21x2_ASAP7_75t_L g520 ( .A1(n_175), .A2(n_521), .B(n_527), .Y(n_520) );
INVxp67_ASAP7_75t_L g257 ( .A(n_176), .Y(n_257) );
AND2x2_ASAP7_75t_L g176 ( .A(n_177), .B(n_192), .Y(n_176) );
NAND2xp5_ASAP7_75t_L g308 ( .A(n_177), .B(n_290), .Y(n_308) );
NAND2xp5_ASAP7_75t_L g329 ( .A(n_177), .B(n_321), .Y(n_329) );
AND2x2_ASAP7_75t_L g379 ( .A(n_177), .B(n_380), .Y(n_379) );
INVx1_ASAP7_75t_L g407 ( .A(n_177), .Y(n_407) );
INVx4_ASAP7_75t_L g177 ( .A(n_178), .Y(n_177) );
AND2x2_ASAP7_75t_L g314 ( .A(n_178), .B(n_307), .Y(n_314) );
BUFx3_ASAP7_75t_L g346 ( .A(n_178), .Y(n_346) );
AO21x2_ASAP7_75t_L g178 ( .A1(n_179), .A2(n_180), .B(n_190), .Y(n_178) );
NOR2xp33_ASAP7_75t_L g495 ( .A(n_179), .B(n_496), .Y(n_495) );
OAI21xp5_ASAP7_75t_L g180 ( .A1(n_181), .A2(n_182), .B(n_183), .Y(n_180) );
OAI21xp5_ASAP7_75t_L g221 ( .A1(n_182), .A2(n_222), .B(n_223), .Y(n_221) );
OAI21xp5_ASAP7_75t_L g521 ( .A1(n_182), .A2(n_522), .B(n_523), .Y(n_521) );
O2A1O1Ixp5_ASAP7_75t_L g184 ( .A1(n_185), .A2(n_186), .B(n_188), .C(n_189), .Y(n_184) );
O2A1O1Ixp33_ASAP7_75t_L g224 ( .A1(n_186), .A2(n_189), .B(n_225), .C(n_226), .Y(n_224) );
O2A1O1Ixp33_ASAP7_75t_L g449 ( .A1(n_186), .A2(n_450), .B(n_451), .C(n_452), .Y(n_449) );
O2A1O1Ixp33_ASAP7_75t_L g482 ( .A1(n_186), .A2(n_452), .B(n_483), .C(n_484), .Y(n_482) );
INVx2_ASAP7_75t_L g186 ( .A(n_187), .Y(n_186) );
INVx2_ASAP7_75t_L g322 ( .A(n_192), .Y(n_322) );
INVx2_ASAP7_75t_L g192 ( .A(n_193), .Y(n_192) );
HB1xp67_ASAP7_75t_L g291 ( .A(n_193), .Y(n_291) );
NOR2xp33_ASAP7_75t_L g236 ( .A(n_198), .B(n_237), .Y(n_236) );
NOR2xp33_ASAP7_75t_L g514 ( .A(n_198), .B(n_515), .Y(n_514) );
INVx2_ASAP7_75t_L g474 ( .A(n_201), .Y(n_474) );
INVx3_ASAP7_75t_L g201 ( .A(n_202), .Y(n_201) );
AOI22xp33_ASAP7_75t_L g381 ( .A1(n_204), .A2(n_382), .B1(n_384), .B2(n_385), .Y(n_381) );
AND2x2_ASAP7_75t_L g204 ( .A(n_205), .B(n_218), .Y(n_204) );
AND2x2_ASAP7_75t_L g241 ( .A(n_205), .B(n_242), .Y(n_241) );
INVx3_ASAP7_75t_SL g252 ( .A(n_205), .Y(n_252) );
NAND2xp5_ASAP7_75t_L g317 ( .A(n_205), .B(n_285), .Y(n_317) );
OR2x2_ASAP7_75t_L g336 ( .A(n_205), .B(n_219), .Y(n_336) );
AND2x2_ASAP7_75t_L g341 ( .A(n_205), .B(n_293), .Y(n_341) );
AND2x2_ASAP7_75t_L g344 ( .A(n_205), .B(n_286), .Y(n_344) );
AND2x2_ASAP7_75t_L g356 ( .A(n_205), .B(n_231), .Y(n_356) );
AND2x2_ASAP7_75t_L g372 ( .A(n_205), .B(n_220), .Y(n_372) );
AND2x4_ASAP7_75t_L g375 ( .A(n_205), .B(n_243), .Y(n_375) );
OR2x2_ASAP7_75t_L g392 ( .A(n_205), .B(n_328), .Y(n_392) );
OR2x2_ASAP7_75t_L g423 ( .A(n_205), .B(n_265), .Y(n_423) );
NAND2xp5_ASAP7_75t_SL g425 ( .A(n_205), .B(n_351), .Y(n_425) );
OR2x6_ASAP7_75t_L g205 ( .A(n_206), .B(n_216), .Y(n_205) );
O2A1O1Ixp33_ASAP7_75t_L g209 ( .A1(n_210), .A2(n_211), .B(n_212), .C(n_213), .Y(n_209) );
NOR2xp33_ASAP7_75t_L g462 ( .A(n_211), .B(n_463), .Y(n_462) );
INVx2_ASAP7_75t_L g513 ( .A(n_211), .Y(n_513) );
AOI21xp5_ASAP7_75t_L g492 ( .A1(n_213), .A2(n_493), .B(n_494), .Y(n_492) );
INVx2_ASAP7_75t_L g213 ( .A(n_214), .Y(n_213) );
NAND2xp5_ASAP7_75t_SL g274 ( .A(n_214), .B(n_275), .Y(n_274) );
AND2x2_ASAP7_75t_L g299 ( .A(n_218), .B(n_263), .Y(n_299) );
NAND2xp5_ASAP7_75t_L g418 ( .A(n_218), .B(n_286), .Y(n_418) );
AND2x2_ASAP7_75t_L g218 ( .A(n_219), .B(n_231), .Y(n_218) );
AND2x2_ASAP7_75t_L g251 ( .A(n_219), .B(n_252), .Y(n_251) );
AND2x2_ASAP7_75t_L g285 ( .A(n_219), .B(n_286), .Y(n_285) );
AND2x2_ASAP7_75t_L g293 ( .A(n_219), .B(n_265), .Y(n_293) );
AND2x2_ASAP7_75t_L g311 ( .A(n_219), .B(n_243), .Y(n_311) );
OR2x2_ASAP7_75t_L g328 ( .A(n_219), .B(n_286), .Y(n_328) );
INVx2_ASAP7_75t_SL g219 ( .A(n_220), .Y(n_219) );
BUFx2_ASAP7_75t_L g244 ( .A(n_220), .Y(n_244) );
AND2x2_ASAP7_75t_L g351 ( .A(n_220), .B(n_231), .Y(n_351) );
NOR2xp33_ASAP7_75t_L g228 ( .A(n_229), .B(n_230), .Y(n_228) );
INVx1_ASAP7_75t_L g280 ( .A(n_230), .Y(n_280) );
INVx2_ASAP7_75t_L g243 ( .A(n_231), .Y(n_243) );
INVx1_ASAP7_75t_L g363 ( .A(n_231), .Y(n_363) );
AND2x2_ASAP7_75t_L g413 ( .A(n_231), .B(n_252), .Y(n_413) );
INVx3_ASAP7_75t_L g238 ( .A(n_239), .Y(n_238) );
HB1xp67_ASAP7_75t_L g504 ( .A(n_239), .Y(n_504) );
AND2x2_ASAP7_75t_L g262 ( .A(n_242), .B(n_263), .Y(n_262) );
AND2x2_ASAP7_75t_L g297 ( .A(n_242), .B(n_252), .Y(n_297) );
NAND2xp5_ASAP7_75t_L g343 ( .A(n_242), .B(n_344), .Y(n_343) );
AND2x2_ASAP7_75t_L g242 ( .A(n_243), .B(n_244), .Y(n_242) );
AND2x2_ASAP7_75t_L g284 ( .A(n_243), .B(n_252), .Y(n_284) );
OR2x2_ASAP7_75t_L g400 ( .A(n_244), .B(n_374), .Y(n_400) );
INVx1_ASAP7_75t_L g245 ( .A(n_246), .Y(n_245) );
NAND2xp5_ASAP7_75t_L g386 ( .A(n_247), .B(n_380), .Y(n_386) );
INVx2_ASAP7_75t_SL g247 ( .A(n_248), .Y(n_247) );
OAI32xp33_ASAP7_75t_L g342 ( .A1(n_248), .A2(n_343), .A3(n_345), .B1(n_347), .B2(n_348), .Y(n_342) );
OR2x2_ASAP7_75t_L g359 ( .A(n_248), .B(n_301), .Y(n_359) );
OAI21xp33_ASAP7_75t_SL g384 ( .A1(n_248), .A2(n_258), .B(n_289), .Y(n_384) );
OAI22xp33_ASAP7_75t_L g249 ( .A1(n_250), .A2(n_253), .B1(n_258), .B2(n_261), .Y(n_249) );
INVxp33_ASAP7_75t_L g250 ( .A(n_251), .Y(n_250) );
NAND2xp5_ASAP7_75t_L g324 ( .A(n_251), .B(n_325), .Y(n_324) );
NAND2xp5_ASAP7_75t_L g292 ( .A(n_252), .B(n_293), .Y(n_292) );
AND2x2_ASAP7_75t_L g310 ( .A(n_252), .B(n_311), .Y(n_310) );
AND2x2_ASAP7_75t_L g410 ( .A(n_252), .B(n_351), .Y(n_410) );
OR2x2_ASAP7_75t_L g434 ( .A(n_252), .B(n_328), .Y(n_434) );
AOI21xp33_ASAP7_75t_L g417 ( .A1(n_253), .A2(n_316), .B(n_418), .Y(n_417) );
OR2x2_ASAP7_75t_L g253 ( .A(n_254), .B(n_257), .Y(n_253) );
NAND2xp5_ASAP7_75t_L g254 ( .A(n_255), .B(n_256), .Y(n_254) );
INVx1_ASAP7_75t_L g294 ( .A(n_255), .Y(n_294) );
NAND2xp5_ASAP7_75t_L g312 ( .A(n_255), .B(n_260), .Y(n_312) );
AND2x2_ASAP7_75t_L g334 ( .A(n_256), .B(n_307), .Y(n_334) );
INVx1_ASAP7_75t_L g347 ( .A(n_256), .Y(n_347) );
OR2x2_ASAP7_75t_L g352 ( .A(n_256), .B(n_286), .Y(n_352) );
NAND2xp5_ASAP7_75t_L g258 ( .A(n_259), .B(n_260), .Y(n_258) );
NOR2xp33_ASAP7_75t_L g300 ( .A(n_259), .B(n_301), .Y(n_300) );
OAI22xp33_ASAP7_75t_L g282 ( .A1(n_260), .A2(n_283), .B1(n_288), .B2(n_292), .Y(n_282) );
INVx1_ASAP7_75t_L g261 ( .A(n_262), .Y(n_261) );
OAI22xp5_ASAP7_75t_L g331 ( .A1(n_263), .A2(n_325), .B1(n_332), .B2(n_333), .Y(n_331) );
AND2x2_ASAP7_75t_L g409 ( .A(n_263), .B(n_410), .Y(n_409) );
INVx2_ASAP7_75t_L g263 ( .A(n_264), .Y(n_263) );
INVx1_ASAP7_75t_SL g264 ( .A(n_265), .Y(n_264) );
NAND2xp5_ASAP7_75t_L g362 ( .A(n_265), .B(n_363), .Y(n_362) );
AND2x2_ASAP7_75t_L g428 ( .A(n_265), .B(n_311), .Y(n_428) );
AO21x2_ASAP7_75t_L g265 ( .A1(n_266), .A2(n_269), .B(n_278), .Y(n_265) );
INVx1_ASAP7_75t_L g287 ( .A(n_266), .Y(n_287) );
INVx1_ASAP7_75t_L g266 ( .A(n_267), .Y(n_266) );
INVx2_ASAP7_75t_L g267 ( .A(n_268), .Y(n_267) );
NOR2xp33_ASAP7_75t_L g527 ( .A(n_268), .B(n_528), .Y(n_527) );
INVx1_ASAP7_75t_L g269 ( .A(n_270), .Y(n_269) );
OA21x2_ASAP7_75t_L g286 ( .A1(n_270), .A2(n_279), .B(n_287), .Y(n_286) );
INVx1_ASAP7_75t_L g278 ( .A(n_279), .Y(n_278) );
AOI21xp5_ASAP7_75t_SL g489 ( .A1(n_280), .A2(n_490), .B(n_491), .Y(n_489) );
AOI221xp5_ASAP7_75t_L g281 ( .A1(n_282), .A2(n_294), .B1(n_295), .B2(n_300), .C(n_302), .Y(n_281) );
NAND2xp5_ASAP7_75t_L g283 ( .A(n_284), .B(n_285), .Y(n_283) );
NAND2xp5_ASAP7_75t_L g316 ( .A(n_284), .B(n_286), .Y(n_316) );
NAND2xp5_ASAP7_75t_L g326 ( .A(n_284), .B(n_327), .Y(n_326) );
INVx1_ASAP7_75t_L g303 ( .A(n_285), .Y(n_303) );
O2A1O1Ixp33_ASAP7_75t_L g390 ( .A1(n_285), .A2(n_391), .B(n_392), .C(n_393), .Y(n_390) );
AND2x2_ASAP7_75t_L g395 ( .A(n_285), .B(n_375), .Y(n_395) );
O2A1O1Ixp33_ASAP7_75t_SL g433 ( .A1(n_285), .A2(n_374), .B(n_434), .C(n_435), .Y(n_433) );
BUFx3_ASAP7_75t_L g325 ( .A(n_286), .Y(n_325) );
INVx1_ASAP7_75t_L g288 ( .A(n_289), .Y(n_288) );
NAND2xp5_ASAP7_75t_L g389 ( .A(n_289), .B(n_346), .Y(n_389) );
AOI211xp5_ASAP7_75t_L g408 ( .A1(n_289), .A2(n_409), .B(n_411), .C(n_417), .Y(n_408) );
AND2x2_ASAP7_75t_L g289 ( .A(n_290), .B(n_291), .Y(n_289) );
INVxp67_ASAP7_75t_L g369 ( .A(n_291), .Y(n_369) );
NAND2xp5_ASAP7_75t_L g412 ( .A(n_293), .B(n_413), .Y(n_412) );
NAND2xp5_ASAP7_75t_SL g295 ( .A(n_296), .B(n_298), .Y(n_295) );
INVx1_ASAP7_75t_SL g296 ( .A(n_297), .Y(n_296) );
AOI211xp5_ASAP7_75t_L g313 ( .A1(n_297), .A2(n_314), .B(n_315), .C(n_323), .Y(n_313) );
INVx1_ASAP7_75t_L g298 ( .A(n_299), .Y(n_298) );
INVx1_ASAP7_75t_L g398 ( .A(n_301), .Y(n_398) );
OR2x2_ASAP7_75t_L g415 ( .A(n_301), .B(n_345), .Y(n_415) );
OAI22xp5_ASAP7_75t_L g302 ( .A1(n_303), .A2(n_304), .B1(n_309), .B2(n_312), .Y(n_302) );
OAI22xp33_ASAP7_75t_L g315 ( .A1(n_304), .A2(n_316), .B1(n_317), .B2(n_318), .Y(n_315) );
INVx1_ASAP7_75t_L g304 ( .A(n_305), .Y(n_304) );
NOR2xp33_ASAP7_75t_L g305 ( .A(n_306), .B(n_308), .Y(n_305) );
OR2x2_ASAP7_75t_L g402 ( .A(n_306), .B(n_346), .Y(n_402) );
INVx1_ASAP7_75t_SL g306 ( .A(n_307), .Y(n_306) );
AND2x2_ASAP7_75t_L g357 ( .A(n_307), .B(n_347), .Y(n_357) );
INVx1_ASAP7_75t_L g365 ( .A(n_308), .Y(n_365) );
INVx1_ASAP7_75t_L g309 ( .A(n_310), .Y(n_309) );
NAND2xp5_ASAP7_75t_L g373 ( .A(n_311), .B(n_325), .Y(n_373) );
INVx1_ASAP7_75t_L g318 ( .A(n_319), .Y(n_318) );
AND2x2_ASAP7_75t_L g319 ( .A(n_320), .B(n_321), .Y(n_319) );
NAND2xp5_ASAP7_75t_SL g364 ( .A(n_321), .B(n_365), .Y(n_364) );
INVx2_ASAP7_75t_L g430 ( .A(n_322), .Y(n_430) );
AOI21xp33_ASAP7_75t_L g323 ( .A1(n_324), .A2(n_326), .B(n_329), .Y(n_323) );
INVx1_ASAP7_75t_L g360 ( .A(n_324), .Y(n_360) );
NAND2xp5_ASAP7_75t_SL g335 ( .A(n_325), .B(n_336), .Y(n_335) );
NAND2xp5_ASAP7_75t_L g355 ( .A(n_325), .B(n_356), .Y(n_355) );
NAND2x1p5_ASAP7_75t_L g376 ( .A(n_325), .B(n_351), .Y(n_376) );
NAND2xp5_ASAP7_75t_SL g383 ( .A(n_325), .B(n_372), .Y(n_383) );
OAI211xp5_ASAP7_75t_L g387 ( .A1(n_325), .A2(n_335), .B(n_375), .C(n_388), .Y(n_387) );
INVx1_ASAP7_75t_SL g327 ( .A(n_328), .Y(n_327) );
AOI221xp5_ASAP7_75t_SL g330 ( .A1(n_331), .A2(n_335), .B1(n_337), .B2(n_341), .C(n_342), .Y(n_330) );
INVx1_ASAP7_75t_L g333 ( .A(n_334), .Y(n_333) );
INVxp67_ASAP7_75t_L g337 ( .A(n_338), .Y(n_337) );
NAND2xp5_ASAP7_75t_L g421 ( .A(n_339), .B(n_347), .Y(n_421) );
INVx1_ASAP7_75t_L g339 ( .A(n_340), .Y(n_339) );
O2A1O1Ixp33_ASAP7_75t_L g432 ( .A1(n_341), .A2(n_356), .B(n_358), .C(n_433), .Y(n_432) );
NAND2xp5_ASAP7_75t_L g416 ( .A(n_344), .B(n_351), .Y(n_416) );
NAND2xp5_ASAP7_75t_SL g435 ( .A(n_345), .B(n_398), .Y(n_435) );
CKINVDCx16_ASAP7_75t_R g345 ( .A(n_346), .Y(n_345) );
INVxp33_ASAP7_75t_L g348 ( .A(n_349), .Y(n_348) );
NOR2xp33_ASAP7_75t_L g349 ( .A(n_350), .B(n_352), .Y(n_349) );
AOI21xp33_ASAP7_75t_SL g361 ( .A1(n_350), .A2(n_362), .B(n_364), .Y(n_361) );
NOR2xp33_ASAP7_75t_L g422 ( .A(n_350), .B(n_423), .Y(n_422) );
INVx2_ASAP7_75t_SL g350 ( .A(n_351), .Y(n_350) );
NAND2xp5_ASAP7_75t_L g404 ( .A(n_351), .B(n_405), .Y(n_404) );
AOI221xp5_ASAP7_75t_L g353 ( .A1(n_354), .A2(n_357), .B1(n_358), .B2(n_360), .C(n_361), .Y(n_353) );
INVx1_ASAP7_75t_L g354 ( .A(n_355), .Y(n_354) );
NAND2xp5_ASAP7_75t_L g406 ( .A(n_357), .B(n_407), .Y(n_406) );
INVx1_ASAP7_75t_L g358 ( .A(n_359), .Y(n_358) );
INVx1_ASAP7_75t_L g391 ( .A(n_363), .Y(n_391) );
NAND5xp2_ASAP7_75t_L g366 ( .A(n_367), .B(n_394), .C(n_408), .D(n_419), .E(n_432), .Y(n_366) );
AOI211xp5_ASAP7_75t_L g367 ( .A1(n_368), .A2(n_370), .B(n_377), .C(n_390), .Y(n_367) );
INVx2_ASAP7_75t_SL g414 ( .A(n_368), .Y(n_414) );
NAND4xp25_ASAP7_75t_SL g370 ( .A(n_371), .B(n_373), .C(n_374), .D(n_376), .Y(n_370) );
INVx1_ASAP7_75t_L g371 ( .A(n_372), .Y(n_371) );
INVx3_ASAP7_75t_L g374 ( .A(n_375), .Y(n_374) );
OAI211xp5_ASAP7_75t_SL g377 ( .A1(n_376), .A2(n_378), .B(n_381), .C(n_387), .Y(n_377) );
CKINVDCx20_ASAP7_75t_R g378 ( .A(n_379), .Y(n_378) );
AOI221xp5_ASAP7_75t_L g419 ( .A1(n_379), .A2(n_420), .B1(n_422), .B2(n_424), .C(n_426), .Y(n_419) );
INVx1_ASAP7_75t_L g382 ( .A(n_383), .Y(n_382) );
INVx1_ASAP7_75t_L g385 ( .A(n_386), .Y(n_385) );
INVx1_ASAP7_75t_L g388 ( .A(n_389), .Y(n_388) );
AOI221xp5_ASAP7_75t_SL g394 ( .A1(n_395), .A2(n_396), .B1(n_399), .B2(n_401), .C(n_403), .Y(n_394) );
AND2x2_ASAP7_75t_L g396 ( .A(n_397), .B(n_398), .Y(n_396) );
INVx1_ASAP7_75t_L g399 ( .A(n_400), .Y(n_399) );
INVx1_ASAP7_75t_L g401 ( .A(n_402), .Y(n_401) );
OAI22xp5_ASAP7_75t_L g426 ( .A1(n_402), .A2(n_425), .B1(n_427), .B2(n_429), .Y(n_426) );
INVx1_ASAP7_75t_L g403 ( .A(n_404), .Y(n_403) );
INVx1_ASAP7_75t_SL g405 ( .A(n_406), .Y(n_405) );
OAI22xp5_ASAP7_75t_L g411 ( .A1(n_412), .A2(n_414), .B1(n_415), .B2(n_416), .Y(n_411) );
INVx1_ASAP7_75t_L g420 ( .A(n_421), .Y(n_420) );
INVx1_ASAP7_75t_L g424 ( .A(n_425), .Y(n_424) );
INVx1_ASAP7_75t_SL g427 ( .A(n_428), .Y(n_427) );
NAND2xp5_ASAP7_75t_L g429 ( .A(n_430), .B(n_431), .Y(n_429) );
INVx1_ASAP7_75t_SL g436 ( .A(n_437), .Y(n_436) );
INVx2_ASAP7_75t_L g437 ( .A(n_438), .Y(n_437) );
INVx1_ASAP7_75t_L g438 ( .A(n_439), .Y(n_438) );
INVx4_ASAP7_75t_L g731 ( .A(n_440), .Y(n_731) );
XOR2xp5_ASAP7_75t_L g741 ( .A(n_440), .B(n_742), .Y(n_741) );
BUFx6f_ASAP7_75t_L g440 ( .A(n_441), .Y(n_440) );
OR5x1_ASAP7_75t_L g441 ( .A(n_442), .B(n_598), .C(n_676), .D(n_700), .E(n_717), .Y(n_441) );
OAI211xp5_ASAP7_75t_SL g442 ( .A1(n_443), .A2(n_475), .B(n_517), .C(n_575), .Y(n_442) );
NAND2xp5_ASAP7_75t_L g443 ( .A(n_444), .B(n_454), .Y(n_443) );
AND2x2_ASAP7_75t_L g529 ( .A(n_444), .B(n_456), .Y(n_529) );
INVx5_ASAP7_75t_SL g557 ( .A(n_444), .Y(n_557) );
AND2x2_ASAP7_75t_L g593 ( .A(n_444), .B(n_578), .Y(n_593) );
OR2x2_ASAP7_75t_L g632 ( .A(n_444), .B(n_455), .Y(n_632) );
OR2x2_ASAP7_75t_L g663 ( .A(n_444), .B(n_554), .Y(n_663) );
NOR2xp33_ASAP7_75t_L g699 ( .A(n_444), .B(n_567), .Y(n_699) );
AND2x2_ASAP7_75t_L g711 ( .A(n_444), .B(n_554), .Y(n_711) );
OR2x6_ASAP7_75t_L g444 ( .A(n_445), .B(n_453), .Y(n_444) );
AND2x2_ASAP7_75t_L g710 ( .A(n_454), .B(n_711), .Y(n_710) );
INVx1_ASAP7_75t_SL g454 ( .A(n_455), .Y(n_454) );
OR2x2_ASAP7_75t_L g573 ( .A(n_455), .B(n_574), .Y(n_573) );
OR2x2_ASAP7_75t_L g455 ( .A(n_456), .B(n_465), .Y(n_455) );
NAND2xp5_ASAP7_75t_L g553 ( .A(n_456), .B(n_554), .Y(n_553) );
HB1xp67_ASAP7_75t_L g566 ( .A(n_456), .Y(n_566) );
INVx3_ASAP7_75t_L g581 ( .A(n_456), .Y(n_581) );
NAND2xp5_ASAP7_75t_L g605 ( .A(n_456), .B(n_465), .Y(n_605) );
OR2x2_ASAP7_75t_L g614 ( .A(n_456), .B(n_557), .Y(n_614) );
AND2x2_ASAP7_75t_L g618 ( .A(n_456), .B(n_578), .Y(n_618) );
AND2x2_ASAP7_75t_L g624 ( .A(n_456), .B(n_625), .Y(n_624) );
INVxp67_ASAP7_75t_L g661 ( .A(n_456), .Y(n_661) );
NAND2xp5_ASAP7_75t_L g675 ( .A(n_456), .B(n_520), .Y(n_675) );
O2A1O1Ixp33_ASAP7_75t_L g501 ( .A1(n_461), .A2(n_502), .B(n_503), .C(n_504), .Y(n_501) );
OR2x2_ASAP7_75t_L g567 ( .A(n_465), .B(n_520), .Y(n_567) );
AND2x2_ASAP7_75t_L g578 ( .A(n_465), .B(n_554), .Y(n_578) );
AND2x2_ASAP7_75t_L g590 ( .A(n_465), .B(n_581), .Y(n_590) );
NAND2xp5_ASAP7_75t_SL g613 ( .A(n_465), .B(n_520), .Y(n_613) );
INVx1_ASAP7_75t_SL g625 ( .A(n_465), .Y(n_625) );
INVx2_ASAP7_75t_L g465 ( .A(n_466), .Y(n_465) );
AND2x2_ASAP7_75t_L g519 ( .A(n_466), .B(n_520), .Y(n_519) );
NAND2xp5_ASAP7_75t_L g556 ( .A(n_466), .B(n_557), .Y(n_556) );
AOI21xp5_ASAP7_75t_L g470 ( .A1(n_471), .A2(n_473), .B(n_474), .Y(n_470) );
AOI21xp5_ASAP7_75t_L g524 ( .A1(n_474), .A2(n_525), .B(n_526), .Y(n_524) );
INVx1_ASAP7_75t_L g475 ( .A(n_476), .Y(n_475) );
AND2x2_ASAP7_75t_L g476 ( .A(n_477), .B(n_487), .Y(n_476) );
AND2x2_ASAP7_75t_L g538 ( .A(n_477), .B(n_539), .Y(n_538) );
NAND2xp5_ASAP7_75t_L g542 ( .A(n_477), .B(n_497), .Y(n_542) );
AND2x2_ASAP7_75t_L g545 ( .A(n_477), .B(n_546), .Y(n_545) );
NAND2xp5_ASAP7_75t_L g547 ( .A(n_477), .B(n_548), .Y(n_547) );
OR2x2_ASAP7_75t_L g570 ( .A(n_477), .B(n_561), .Y(n_570) );
HB1xp67_ASAP7_75t_L g589 ( .A(n_477), .Y(n_589) );
AND2x2_ASAP7_75t_L g610 ( .A(n_477), .B(n_611), .Y(n_610) );
OR2x2_ASAP7_75t_L g620 ( .A(n_477), .B(n_621), .Y(n_620) );
AND2x2_ASAP7_75t_L g666 ( .A(n_477), .B(n_549), .Y(n_666) );
NAND2xp5_ASAP7_75t_L g693 ( .A(n_477), .B(n_572), .Y(n_693) );
INVx5_ASAP7_75t_L g477 ( .A(n_478), .Y(n_477) );
BUFx2_ASAP7_75t_L g563 ( .A(n_478), .Y(n_563) );
AND2x2_ASAP7_75t_L g629 ( .A(n_478), .B(n_561), .Y(n_629) );
AND2x2_ASAP7_75t_L g713 ( .A(n_478), .B(n_581), .Y(n_713) );
OR2x6_ASAP7_75t_L g478 ( .A(n_479), .B(n_485), .Y(n_478) );
NAND2xp5_ASAP7_75t_L g698 ( .A(n_487), .B(n_699), .Y(n_698) );
INVx1_ASAP7_75t_L g702 ( .A(n_487), .Y(n_702) );
AND2x2_ASAP7_75t_L g487 ( .A(n_488), .B(n_497), .Y(n_487) );
AND2x2_ASAP7_75t_L g532 ( .A(n_488), .B(n_533), .Y(n_532) );
AND2x4_ASAP7_75t_L g541 ( .A(n_488), .B(n_539), .Y(n_541) );
INVx5_ASAP7_75t_L g549 ( .A(n_488), .Y(n_549) );
AND2x2_ASAP7_75t_L g572 ( .A(n_488), .B(n_508), .Y(n_572) );
HB1xp67_ASAP7_75t_L g609 ( .A(n_488), .Y(n_609) );
OR2x6_ASAP7_75t_L g488 ( .A(n_489), .B(n_495), .Y(n_488) );
INVx1_ASAP7_75t_L g650 ( .A(n_497), .Y(n_650) );
NAND2xp5_ASAP7_75t_L g665 ( .A(n_497), .B(n_666), .Y(n_665) );
AND2x2_ASAP7_75t_L g683 ( .A(n_497), .B(n_549), .Y(n_683) );
A2O1A1Ixp33_ASAP7_75t_L g712 ( .A1(n_497), .A2(n_606), .B(n_713), .C(n_714), .Y(n_712) );
AND2x2_ASAP7_75t_L g497 ( .A(n_498), .B(n_508), .Y(n_497) );
BUFx2_ASAP7_75t_L g533 ( .A(n_498), .Y(n_533) );
INVx2_ASAP7_75t_L g537 ( .A(n_498), .Y(n_537) );
NAND2xp5_ASAP7_75t_L g499 ( .A(n_500), .B(n_505), .Y(n_499) );
INVx2_ASAP7_75t_L g539 ( .A(n_508), .Y(n_539) );
AND2x2_ASAP7_75t_L g546 ( .A(n_508), .B(n_537), .Y(n_546) );
AND2x2_ASAP7_75t_L g637 ( .A(n_508), .B(n_549), .Y(n_637) );
AOI211x1_ASAP7_75t_SL g517 ( .A1(n_518), .A2(n_530), .B(n_543), .C(n_568), .Y(n_517) );
INVx1_ASAP7_75t_L g634 ( .A(n_518), .Y(n_634) );
AND2x2_ASAP7_75t_L g518 ( .A(n_519), .B(n_529), .Y(n_518) );
INVx5_ASAP7_75t_SL g554 ( .A(n_520), .Y(n_554) );
NAND2xp5_ASAP7_75t_L g623 ( .A(n_520), .B(n_624), .Y(n_623) );
AOI311xp33_ASAP7_75t_L g642 ( .A1(n_520), .A2(n_643), .A3(n_645), .B(n_646), .C(n_652), .Y(n_642) );
A2O1A1Ixp33_ASAP7_75t_L g677 ( .A1(n_520), .A2(n_590), .B(n_678), .C(n_681), .Y(n_677) );
INVxp67_ASAP7_75t_L g597 ( .A(n_529), .Y(n_597) );
NAND4xp25_ASAP7_75t_SL g530 ( .A(n_531), .B(n_534), .C(n_540), .D(n_542), .Y(n_530) );
NOR2xp33_ASAP7_75t_L g595 ( .A(n_531), .B(n_596), .Y(n_595) );
INVx2_ASAP7_75t_L g531 ( .A(n_532), .Y(n_531) );
AND2x2_ASAP7_75t_L g588 ( .A(n_532), .B(n_589), .Y(n_588) );
NAND2xp5_ASAP7_75t_L g534 ( .A(n_535), .B(n_538), .Y(n_534) );
NAND2xp5_ASAP7_75t_L g584 ( .A(n_535), .B(n_541), .Y(n_584) );
NAND2xp5_ASAP7_75t_L g668 ( .A(n_535), .B(n_548), .Y(n_668) );
BUFx2_ASAP7_75t_L g535 ( .A(n_536), .Y(n_535) );
NAND2xp5_ASAP7_75t_L g686 ( .A(n_536), .B(n_549), .Y(n_686) );
HB1xp67_ASAP7_75t_L g536 ( .A(n_537), .Y(n_536) );
INVx2_ASAP7_75t_L g561 ( .A(n_537), .Y(n_561) );
INVxp67_ASAP7_75t_L g596 ( .A(n_538), .Y(n_596) );
AND2x4_ASAP7_75t_L g548 ( .A(n_539), .B(n_549), .Y(n_548) );
AND2x2_ASAP7_75t_L g622 ( .A(n_539), .B(n_561), .Y(n_622) );
INVx1_ASAP7_75t_L g649 ( .A(n_539), .Y(n_649) );
NAND2xp5_ASAP7_75t_L g696 ( .A(n_539), .B(n_636), .Y(n_696) );
NOR2xp33_ASAP7_75t_L g630 ( .A(n_540), .B(n_610), .Y(n_630) );
INVx1_ASAP7_75t_SL g540 ( .A(n_541), .Y(n_540) );
NAND2xp5_ASAP7_75t_L g707 ( .A(n_541), .B(n_563), .Y(n_707) );
NAND2xp5_ASAP7_75t_L g709 ( .A(n_541), .B(n_610), .Y(n_709) );
INVx1_ASAP7_75t_L g720 ( .A(n_542), .Y(n_720) );
A2O1A1Ixp33_ASAP7_75t_L g543 ( .A1(n_544), .A2(n_547), .B(n_550), .C(n_558), .Y(n_543) );
INVx1_ASAP7_75t_SL g544 ( .A(n_545), .Y(n_544) );
AND2x2_ASAP7_75t_L g562 ( .A(n_546), .B(n_563), .Y(n_562) );
AND2x2_ASAP7_75t_L g600 ( .A(n_546), .B(n_601), .Y(n_600) );
INVx1_ASAP7_75t_L g582 ( .A(n_547), .Y(n_582) );
AND2x2_ASAP7_75t_L g559 ( .A(n_548), .B(n_560), .Y(n_559) );
NAND2xp5_ASAP7_75t_L g644 ( .A(n_548), .B(n_610), .Y(n_644) );
NAND2xp5_ASAP7_75t_L g653 ( .A(n_548), .B(n_629), .Y(n_653) );
OR2x2_ASAP7_75t_L g569 ( .A(n_549), .B(n_570), .Y(n_569) );
INVx2_ASAP7_75t_L g601 ( .A(n_549), .Y(n_601) );
NAND2xp5_ASAP7_75t_L g616 ( .A(n_549), .B(n_561), .Y(n_616) );
AND2x2_ASAP7_75t_L g673 ( .A(n_549), .B(n_629), .Y(n_673) );
HB1xp67_ASAP7_75t_L g680 ( .A(n_549), .Y(n_680) );
INVx1_ASAP7_75t_L g550 ( .A(n_551), .Y(n_550) );
AOI221xp5_ASAP7_75t_L g684 ( .A1(n_551), .A2(n_563), .B1(n_685), .B2(n_687), .C(n_690), .Y(n_684) );
AND2x2_ASAP7_75t_L g551 ( .A(n_552), .B(n_555), .Y(n_551) );
INVx1_ASAP7_75t_SL g552 ( .A(n_553), .Y(n_552) );
OR2x2_ASAP7_75t_L g574 ( .A(n_554), .B(n_557), .Y(n_574) );
NAND2xp5_ASAP7_75t_L g670 ( .A(n_554), .B(n_624), .Y(n_670) );
NAND2xp5_ASAP7_75t_L g689 ( .A(n_554), .B(n_581), .Y(n_689) );
INVx1_ASAP7_75t_SL g555 ( .A(n_556), .Y(n_555) );
OR2x2_ASAP7_75t_L g674 ( .A(n_556), .B(n_675), .Y(n_674) );
OR2x2_ASAP7_75t_L g688 ( .A(n_556), .B(n_689), .Y(n_688) );
NAND2xp5_ASAP7_75t_L g580 ( .A(n_557), .B(n_581), .Y(n_580) );
AND2x2_ASAP7_75t_L g585 ( .A(n_557), .B(n_578), .Y(n_585) );
AND2x2_ASAP7_75t_L g655 ( .A(n_557), .B(n_656), .Y(n_655) );
NAND2xp5_ASAP7_75t_L g701 ( .A(n_557), .B(n_604), .Y(n_701) );
NOR2xp33_ASAP7_75t_L g704 ( .A(n_557), .B(n_705), .Y(n_704) );
OAI21xp5_ASAP7_75t_SL g558 ( .A1(n_559), .A2(n_562), .B(n_564), .Y(n_558) );
INVx2_ASAP7_75t_L g591 ( .A(n_559), .Y(n_591) );
HB1xp67_ASAP7_75t_L g560 ( .A(n_561), .Y(n_560) );
INVx1_ASAP7_75t_L g611 ( .A(n_561), .Y(n_611) );
OR2x2_ASAP7_75t_L g615 ( .A(n_563), .B(n_616), .Y(n_615) );
OR2x2_ASAP7_75t_L g718 ( .A(n_563), .B(n_686), .Y(n_718) );
INVx1_ASAP7_75t_SL g564 ( .A(n_565), .Y(n_564) );
OR2x2_ASAP7_75t_L g565 ( .A(n_566), .B(n_567), .Y(n_565) );
AOI21xp33_ASAP7_75t_SL g568 ( .A1(n_569), .A2(n_571), .B(n_573), .Y(n_568) );
INVx1_ASAP7_75t_L g722 ( .A(n_569), .Y(n_722) );
INVx2_ASAP7_75t_SL g636 ( .A(n_570), .Y(n_636) );
INVx1_ASAP7_75t_L g571 ( .A(n_572), .Y(n_571) );
A2O1A1Ixp33_ASAP7_75t_L g717 ( .A1(n_573), .A2(n_654), .B(n_718), .C(n_719), .Y(n_717) );
OAI322xp33_ASAP7_75t_SL g586 ( .A1(n_574), .A2(n_587), .A3(n_590), .B1(n_591), .B2(n_592), .C1(n_594), .C2(n_597), .Y(n_586) );
INVx2_ASAP7_75t_L g606 ( .A(n_574), .Y(n_606) );
AOI221xp5_ASAP7_75t_L g575 ( .A1(n_576), .A2(n_582), .B1(n_583), .B2(n_585), .C(n_586), .Y(n_575) );
INVx1_ASAP7_75t_L g576 ( .A(n_577), .Y(n_576) );
OAI22xp33_ASAP7_75t_SL g652 ( .A1(n_577), .A2(n_653), .B1(n_654), .B2(n_657), .Y(n_652) );
NAND2xp5_ASAP7_75t_L g577 ( .A(n_578), .B(n_579), .Y(n_577) );
NAND2xp5_ASAP7_75t_L g692 ( .A(n_578), .B(n_581), .Y(n_692) );
NAND2xp5_ASAP7_75t_L g715 ( .A(n_578), .B(n_716), .Y(n_715) );
INVx2_ASAP7_75t_L g579 ( .A(n_580), .Y(n_579) );
OR2x2_ASAP7_75t_L g651 ( .A(n_580), .B(n_613), .Y(n_651) );
INVx1_ASAP7_75t_L g641 ( .A(n_581), .Y(n_641) );
INVx1_ASAP7_75t_L g583 ( .A(n_584), .Y(n_583) );
AOI21xp5_ASAP7_75t_L g694 ( .A1(n_585), .A2(n_695), .B(n_697), .Y(n_694) );
AOI21xp33_ASAP7_75t_L g619 ( .A1(n_587), .A2(n_620), .B(n_623), .Y(n_619) );
INVx1_ASAP7_75t_L g587 ( .A(n_588), .Y(n_587) );
NOR2xp67_ASAP7_75t_SL g648 ( .A(n_589), .B(n_649), .Y(n_648) );
NOR2xp33_ASAP7_75t_L g681 ( .A(n_589), .B(n_682), .Y(n_681) );
INVx1_ASAP7_75t_SL g705 ( .A(n_590), .Y(n_705) );
INVx1_ASAP7_75t_SL g592 ( .A(n_593), .Y(n_592) );
INVx1_ASAP7_75t_L g594 ( .A(n_595), .Y(n_594) );
NAND4xp25_ASAP7_75t_L g598 ( .A(n_599), .B(n_626), .C(n_642), .D(n_658), .Y(n_598) );
AOI211xp5_ASAP7_75t_L g599 ( .A1(n_600), .A2(n_602), .B(n_607), .C(n_619), .Y(n_599) );
INVx1_ASAP7_75t_L g691 ( .A(n_600), .Y(n_691) );
AND2x2_ASAP7_75t_L g639 ( .A(n_601), .B(n_622), .Y(n_639) );
INVx1_ASAP7_75t_L g602 ( .A(n_603), .Y(n_602) );
NAND2xp5_ASAP7_75t_L g603 ( .A(n_604), .B(n_606), .Y(n_603) );
INVx1_ASAP7_75t_SL g604 ( .A(n_605), .Y(n_604) );
NAND2xp5_ASAP7_75t_L g640 ( .A(n_606), .B(n_641), .Y(n_640) );
OAI22xp33_ASAP7_75t_L g607 ( .A1(n_608), .A2(n_612), .B1(n_615), .B2(n_617), .Y(n_607) );
NAND2xp5_ASAP7_75t_L g608 ( .A(n_609), .B(n_610), .Y(n_608) );
NAND2xp5_ASAP7_75t_L g628 ( .A(n_609), .B(n_629), .Y(n_628) );
INVx1_ASAP7_75t_L g657 ( .A(n_610), .Y(n_657) );
O2A1O1Ixp33_ASAP7_75t_L g671 ( .A1(n_610), .A2(n_649), .B(n_672), .C(n_674), .Y(n_671) );
OR2x2_ASAP7_75t_L g612 ( .A(n_613), .B(n_614), .Y(n_612) );
INVx1_ASAP7_75t_L g656 ( .A(n_613), .Y(n_656) );
INVx1_ASAP7_75t_L g716 ( .A(n_614), .Y(n_716) );
NAND2xp33_ASAP7_75t_SL g706 ( .A(n_615), .B(n_707), .Y(n_706) );
INVx1_ASAP7_75t_SL g617 ( .A(n_618), .Y(n_617) );
INVx1_ASAP7_75t_L g621 ( .A(n_622), .Y(n_621) );
INVx2_ASAP7_75t_L g645 ( .A(n_624), .Y(n_645) );
O2A1O1Ixp33_ASAP7_75t_L g626 ( .A1(n_627), .A2(n_630), .B(n_631), .C(n_633), .Y(n_626) );
INVx1_ASAP7_75t_L g627 ( .A(n_628), .Y(n_627) );
INVx1_ASAP7_75t_L g631 ( .A(n_632), .Y(n_631) );
OAI22xp5_ASAP7_75t_L g633 ( .A1(n_634), .A2(n_635), .B1(n_638), .B2(n_640), .Y(n_633) );
NAND2xp5_ASAP7_75t_L g635 ( .A(n_636), .B(n_637), .Y(n_635) );
NAND2xp5_ASAP7_75t_L g679 ( .A(n_636), .B(n_680), .Y(n_679) );
INVx1_ASAP7_75t_L g638 ( .A(n_639), .Y(n_638) );
NAND2xp5_ASAP7_75t_L g724 ( .A(n_641), .B(n_662), .Y(n_724) );
INVx1_ASAP7_75t_L g643 ( .A(n_644), .Y(n_643) );
AOI21xp33_ASAP7_75t_SL g646 ( .A1(n_647), .A2(n_650), .B(n_651), .Y(n_646) );
INVx1_ASAP7_75t_L g647 ( .A(n_648), .Y(n_647) );
INVx1_ASAP7_75t_SL g654 ( .A(n_655), .Y(n_654) );
AOI221xp5_ASAP7_75t_L g658 ( .A1(n_659), .A2(n_664), .B1(n_667), .B2(n_669), .C(n_671), .Y(n_658) );
INVx1_ASAP7_75t_L g659 ( .A(n_660), .Y(n_659) );
NAND2xp5_ASAP7_75t_L g660 ( .A(n_661), .B(n_662), .Y(n_660) );
INVx1_ASAP7_75t_SL g662 ( .A(n_663), .Y(n_662) );
INVx1_ASAP7_75t_L g664 ( .A(n_665), .Y(n_664) );
INVx1_ASAP7_75t_L g667 ( .A(n_668), .Y(n_667) );
INVxp67_ASAP7_75t_L g669 ( .A(n_670), .Y(n_669) );
INVx1_ASAP7_75t_L g672 ( .A(n_673), .Y(n_672) );
OAI22xp5_ASAP7_75t_L g690 ( .A1(n_674), .A2(n_691), .B1(n_692), .B2(n_693), .Y(n_690) );
NAND3xp33_ASAP7_75t_SL g676 ( .A(n_677), .B(n_684), .C(n_694), .Y(n_676) );
INVx1_ASAP7_75t_L g678 ( .A(n_679), .Y(n_678) );
INVx1_ASAP7_75t_SL g682 ( .A(n_683), .Y(n_682) );
INVx1_ASAP7_75t_L g685 ( .A(n_686), .Y(n_685) );
CKINVDCx16_ASAP7_75t_R g687 ( .A(n_688), .Y(n_687) );
INVx1_ASAP7_75t_L g695 ( .A(n_696), .Y(n_695) );
INVxp67_ASAP7_75t_L g697 ( .A(n_698), .Y(n_697) );
OAI211xp5_ASAP7_75t_L g700 ( .A1(n_701), .A2(n_702), .B(n_703), .C(n_712), .Y(n_700) );
INVx1_ASAP7_75t_L g721 ( .A(n_701), .Y(n_721) );
AOI22xp33_ASAP7_75t_L g703 ( .A1(n_704), .A2(n_706), .B1(n_708), .B2(n_710), .Y(n_703) );
INVx1_ASAP7_75t_L g708 ( .A(n_709), .Y(n_708) );
INVx1_ASAP7_75t_L g714 ( .A(n_715), .Y(n_714) );
AOI22xp5_ASAP7_75t_L g719 ( .A1(n_720), .A2(n_721), .B1(n_722), .B2(n_723), .Y(n_719) );
INVx1_ASAP7_75t_L g723 ( .A(n_724), .Y(n_723) );
CKINVDCx16_ASAP7_75t_R g725 ( .A(n_726), .Y(n_725) );
INVx2_ASAP7_75t_L g732 ( .A(n_733), .Y(n_732) );
BUFx2_ASAP7_75t_L g736 ( .A(n_737), .Y(n_736) );
INVx2_ASAP7_75t_L g737 ( .A(n_738), .Y(n_737) );
INVx1_ASAP7_75t_L g748 ( .A(n_738), .Y(n_748) );
INVxp67_ASAP7_75t_L g739 ( .A(n_740), .Y(n_739) );
NAND2xp5_ASAP7_75t_L g740 ( .A(n_741), .B(n_745), .Y(n_740) );
BUFx2_ASAP7_75t_L g745 ( .A(n_746), .Y(n_745) );
INVx2_ASAP7_75t_L g752 ( .A(n_746), .Y(n_752) );
INVx1_ASAP7_75t_L g747 ( .A(n_748), .Y(n_747) );
NOR2xp33_ASAP7_75t_L g749 ( .A(n_750), .B(n_751), .Y(n_749) );
INVx1_ASAP7_75t_L g751 ( .A(n_752), .Y(n_751) );
endmodule