module fake_netlist_5_1872_n_1243 (n_137, n_294, n_318, n_82, n_194, n_316, n_248, n_124, n_86, n_136, n_146, n_315, n_268, n_61, n_127, n_75, n_235, n_226, n_74, n_57, n_111, n_155, n_43, n_116, n_22, n_284, n_46, n_245, n_21, n_139, n_38, n_105, n_280, n_4, n_17, n_254, n_33, n_23, n_302, n_265, n_293, n_244, n_47, n_173, n_198, n_247, n_314, n_8, n_321, n_292, n_100, n_212, n_119, n_275, n_252, n_26, n_295, n_133, n_330, n_2, n_6, n_39, n_147, n_67, n_307, n_87, n_150, n_106, n_209, n_259, n_301, n_68, n_93, n_186, n_134, n_191, n_51, n_63, n_171, n_153, n_204, n_250, n_260, n_298, n_320, n_286, n_122, n_282, n_331, n_10, n_24, n_325, n_132, n_90, n_101, n_281, n_240, n_189, n_220, n_291, n_231, n_257, n_31, n_13, n_152, n_317, n_9, n_323, n_195, n_42, n_227, n_45, n_271, n_94, n_123, n_167, n_234, n_308, n_267, n_297, n_156, n_5, n_225, n_219, n_157, n_131, n_192, n_223, n_158, n_138, n_264, n_109, n_163, n_276, n_95, n_183, n_185, n_243, n_169, n_59, n_255, n_215, n_196, n_211, n_218, n_181, n_3, n_290, n_221, n_178, n_287, n_72, n_104, n_41, n_56, n_141, n_15, n_145, n_48, n_50, n_313, n_88, n_216, n_168, n_164, n_311, n_208, n_142, n_214, n_328, n_140, n_299, n_303, n_296, n_241, n_184, n_65, n_78, n_144, n_114, n_96, n_165, n_213, n_129, n_98, n_197, n_107, n_69, n_236, n_1, n_249, n_304, n_329, n_203, n_274, n_80, n_35, n_73, n_277, n_92, n_19, n_149, n_309, n_30, n_14, n_84, n_130, n_322, n_258, n_29, n_79, n_151, n_25, n_306, n_288, n_188, n_190, n_201, n_263, n_44, n_224, n_40, n_34, n_228, n_283, n_112, n_85, n_239, n_55, n_49, n_310, n_54, n_12, n_76, n_170, n_27, n_77, n_102, n_161, n_273, n_270, n_230, n_81, n_118, n_279, n_70, n_253, n_261, n_174, n_289, n_172, n_206, n_217, n_312, n_210, n_91, n_176, n_182, n_143, n_83, n_237, n_180, n_207, n_37, n_229, n_108, n_66, n_177, n_60, n_16, n_0, n_58, n_18, n_117, n_326, n_233, n_205, n_113, n_246, n_179, n_125, n_269, n_128, n_285, n_120, n_232, n_327, n_135, n_126, n_202, n_266, n_272, n_193, n_251, n_53, n_160, n_154, n_62, n_148, n_71, n_300, n_159, n_175, n_262, n_238, n_99, n_319, n_20, n_121, n_242, n_36, n_200, n_162, n_64, n_222, n_28, n_89, n_115, n_324, n_199, n_187, n_32, n_103, n_97, n_166, n_11, n_7, n_256, n_305, n_52, n_278, n_110, n_1243);

input n_137;
input n_294;
input n_318;
input n_82;
input n_194;
input n_316;
input n_248;
input n_124;
input n_86;
input n_136;
input n_146;
input n_315;
input n_268;
input n_61;
input n_127;
input n_75;
input n_235;
input n_226;
input n_74;
input n_57;
input n_111;
input n_155;
input n_43;
input n_116;
input n_22;
input n_284;
input n_46;
input n_245;
input n_21;
input n_139;
input n_38;
input n_105;
input n_280;
input n_4;
input n_17;
input n_254;
input n_33;
input n_23;
input n_302;
input n_265;
input n_293;
input n_244;
input n_47;
input n_173;
input n_198;
input n_247;
input n_314;
input n_8;
input n_321;
input n_292;
input n_100;
input n_212;
input n_119;
input n_275;
input n_252;
input n_26;
input n_295;
input n_133;
input n_330;
input n_2;
input n_6;
input n_39;
input n_147;
input n_67;
input n_307;
input n_87;
input n_150;
input n_106;
input n_209;
input n_259;
input n_301;
input n_68;
input n_93;
input n_186;
input n_134;
input n_191;
input n_51;
input n_63;
input n_171;
input n_153;
input n_204;
input n_250;
input n_260;
input n_298;
input n_320;
input n_286;
input n_122;
input n_282;
input n_331;
input n_10;
input n_24;
input n_325;
input n_132;
input n_90;
input n_101;
input n_281;
input n_240;
input n_189;
input n_220;
input n_291;
input n_231;
input n_257;
input n_31;
input n_13;
input n_152;
input n_317;
input n_9;
input n_323;
input n_195;
input n_42;
input n_227;
input n_45;
input n_271;
input n_94;
input n_123;
input n_167;
input n_234;
input n_308;
input n_267;
input n_297;
input n_156;
input n_5;
input n_225;
input n_219;
input n_157;
input n_131;
input n_192;
input n_223;
input n_158;
input n_138;
input n_264;
input n_109;
input n_163;
input n_276;
input n_95;
input n_183;
input n_185;
input n_243;
input n_169;
input n_59;
input n_255;
input n_215;
input n_196;
input n_211;
input n_218;
input n_181;
input n_3;
input n_290;
input n_221;
input n_178;
input n_287;
input n_72;
input n_104;
input n_41;
input n_56;
input n_141;
input n_15;
input n_145;
input n_48;
input n_50;
input n_313;
input n_88;
input n_216;
input n_168;
input n_164;
input n_311;
input n_208;
input n_142;
input n_214;
input n_328;
input n_140;
input n_299;
input n_303;
input n_296;
input n_241;
input n_184;
input n_65;
input n_78;
input n_144;
input n_114;
input n_96;
input n_165;
input n_213;
input n_129;
input n_98;
input n_197;
input n_107;
input n_69;
input n_236;
input n_1;
input n_249;
input n_304;
input n_329;
input n_203;
input n_274;
input n_80;
input n_35;
input n_73;
input n_277;
input n_92;
input n_19;
input n_149;
input n_309;
input n_30;
input n_14;
input n_84;
input n_130;
input n_322;
input n_258;
input n_29;
input n_79;
input n_151;
input n_25;
input n_306;
input n_288;
input n_188;
input n_190;
input n_201;
input n_263;
input n_44;
input n_224;
input n_40;
input n_34;
input n_228;
input n_283;
input n_112;
input n_85;
input n_239;
input n_55;
input n_49;
input n_310;
input n_54;
input n_12;
input n_76;
input n_170;
input n_27;
input n_77;
input n_102;
input n_161;
input n_273;
input n_270;
input n_230;
input n_81;
input n_118;
input n_279;
input n_70;
input n_253;
input n_261;
input n_174;
input n_289;
input n_172;
input n_206;
input n_217;
input n_312;
input n_210;
input n_91;
input n_176;
input n_182;
input n_143;
input n_83;
input n_237;
input n_180;
input n_207;
input n_37;
input n_229;
input n_108;
input n_66;
input n_177;
input n_60;
input n_16;
input n_0;
input n_58;
input n_18;
input n_117;
input n_326;
input n_233;
input n_205;
input n_113;
input n_246;
input n_179;
input n_125;
input n_269;
input n_128;
input n_285;
input n_120;
input n_232;
input n_327;
input n_135;
input n_126;
input n_202;
input n_266;
input n_272;
input n_193;
input n_251;
input n_53;
input n_160;
input n_154;
input n_62;
input n_148;
input n_71;
input n_300;
input n_159;
input n_175;
input n_262;
input n_238;
input n_99;
input n_319;
input n_20;
input n_121;
input n_242;
input n_36;
input n_200;
input n_162;
input n_64;
input n_222;
input n_28;
input n_89;
input n_115;
input n_324;
input n_199;
input n_187;
input n_32;
input n_103;
input n_97;
input n_166;
input n_11;
input n_7;
input n_256;
input n_305;
input n_52;
input n_278;
input n_110;

output n_1243;

wire n_924;
wire n_977;
wire n_611;
wire n_1126;
wire n_1166;
wire n_469;
wire n_785;
wire n_549;
wire n_532;
wire n_1161;
wire n_1150;
wire n_667;
wire n_790;
wire n_1055;
wire n_880;
wire n_544;
wire n_1007;
wire n_552;
wire n_1198;
wire n_1099;
wire n_956;
wire n_564;
wire n_423;
wire n_1021;
wire n_551;
wire n_688;
wire n_800;
wire n_671;
wire n_819;
wire n_1022;
wire n_915;
wire n_864;
wire n_859;
wire n_951;
wire n_447;
wire n_625;
wire n_854;
wire n_674;
wire n_417;
wire n_516;
wire n_933;
wire n_1152;
wire n_497;
wire n_606;
wire n_877;
wire n_755;
wire n_1118;
wire n_947;
wire n_373;
wire n_530;
wire n_1107;
wire n_556;
wire n_1230;
wire n_668;
wire n_375;
wire n_929;
wire n_1124;
wire n_902;
wire n_1104;
wire n_659;
wire n_1182;
wire n_579;
wire n_938;
wire n_1098;
wire n_1154;
wire n_1242;
wire n_1135;
wire n_406;
wire n_519;
wire n_1016;
wire n_546;
wire n_731;
wire n_371;
wire n_709;
wire n_1236;
wire n_569;
wire n_920;
wire n_335;
wire n_370;
wire n_976;
wire n_343;
wire n_1078;
wire n_775;
wire n_600;
wire n_955;
wire n_339;
wire n_1146;
wire n_882;
wire n_1036;
wire n_1097;
wire n_347;
wire n_550;
wire n_696;
wire n_897;
wire n_798;
wire n_350;
wire n_646;
wire n_436;
wire n_1216;
wire n_580;
wire n_1040;
wire n_578;
wire n_926;
wire n_344;
wire n_1218;
wire n_475;
wire n_422;
wire n_777;
wire n_1070;
wire n_1030;
wire n_415;
wire n_1071;
wire n_485;
wire n_1165;
wire n_496;
wire n_958;
wire n_1034;
wire n_670;
wire n_521;
wire n_663;
wire n_845;
wire n_673;
wire n_837;
wire n_1239;
wire n_528;
wire n_680;
wire n_395;
wire n_553;
wire n_901;
wire n_813;
wire n_675;
wire n_888;
wire n_1167;
wire n_637;
wire n_446;
wire n_1064;
wire n_858;
wire n_923;
wire n_691;
wire n_1151;
wire n_881;
wire n_468;
wire n_342;
wire n_464;
wire n_363;
wire n_1069;
wire n_1075;
wire n_460;
wire n_889;
wire n_973;
wire n_477;
wire n_571;
wire n_461;
wire n_1211;
wire n_1197;
wire n_907;
wire n_989;
wire n_1039;
wire n_488;
wire n_736;
wire n_892;
wire n_1000;
wire n_1202;
wire n_1002;
wire n_593;
wire n_748;
wire n_586;
wire n_1058;
wire n_838;
wire n_332;
wire n_1053;
wire n_1224;
wire n_349;
wire n_953;
wire n_1014;
wire n_1241;
wire n_963;
wire n_1052;
wire n_954;
wire n_627;
wire n_440;
wire n_793;
wire n_478;
wire n_476;
wire n_534;
wire n_884;
wire n_345;
wire n_944;
wire n_647;
wire n_407;
wire n_1072;
wire n_832;
wire n_857;
wire n_561;
wire n_1027;
wire n_971;
wire n_1156;
wire n_794;
wire n_404;
wire n_686;
wire n_847;
wire n_596;
wire n_558;
wire n_702;
wire n_822;
wire n_728;
wire n_1162;
wire n_1199;
wire n_352;
wire n_1038;
wire n_520;
wire n_409;
wire n_887;
wire n_809;
wire n_870;
wire n_931;
wire n_599;
wire n_434;
wire n_868;
wire n_639;
wire n_914;
wire n_411;
wire n_414;
wire n_965;
wire n_935;
wire n_1175;
wire n_817;
wire n_360;
wire n_759;
wire n_806;
wire n_1189;
wire n_706;
wire n_746;
wire n_747;
wire n_784;
wire n_431;
wire n_1194;
wire n_615;
wire n_851;
wire n_843;
wire n_523;
wire n_913;
wire n_705;
wire n_865;
wire n_678;
wire n_697;
wire n_1222;
wire n_776;
wire n_367;
wire n_452;
wire n_525;
wire n_649;
wire n_547;
wire n_1191;
wire n_1128;
wire n_744;
wire n_590;
wire n_629;
wire n_1233;
wire n_526;
wire n_372;
wire n_677;
wire n_1121;
wire n_368;
wire n_433;
wire n_604;
wire n_949;
wire n_1008;
wire n_946;
wire n_1001;
wire n_498;
wire n_689;
wire n_738;
wire n_640;
wire n_624;
wire n_1010;
wire n_1231;
wire n_739;
wire n_1195;
wire n_610;
wire n_936;
wire n_568;
wire n_1090;
wire n_757;
wire n_633;
wire n_439;
wire n_448;
wire n_758;
wire n_999;
wire n_1158;
wire n_563;
wire n_1145;
wire n_878;
wire n_524;
wire n_394;
wire n_1049;
wire n_1153;
wire n_741;
wire n_1068;
wire n_906;
wire n_1163;
wire n_1207;
wire n_919;
wire n_908;
wire n_724;
wire n_658;
wire n_456;
wire n_959;
wire n_535;
wire n_940;
wire n_592;
wire n_1169;
wire n_1017;
wire n_978;
wire n_1054;
wire n_1095;
wire n_514;
wire n_457;
wire n_1079;
wire n_1045;
wire n_1208;
wire n_603;
wire n_484;
wire n_1033;
wire n_442;
wire n_636;
wire n_660;
wire n_1009;
wire n_1148;
wire n_750;
wire n_742;
wire n_995;
wire n_454;
wire n_374;
wire n_396;
wire n_1073;
wire n_662;
wire n_459;
wire n_962;
wire n_1215;
wire n_1171;
wire n_723;
wire n_1065;
wire n_473;
wire n_1043;
wire n_355;
wire n_486;
wire n_614;
wire n_337;
wire n_1177;
wire n_974;
wire n_727;
wire n_1159;
wire n_957;
wire n_773;
wire n_743;
wire n_613;
wire n_1119;
wire n_1240;
wire n_829;
wire n_361;
wire n_1237;
wire n_700;
wire n_573;
wire n_1132;
wire n_388;
wire n_1127;
wire n_761;
wire n_1006;
wire n_582;
wire n_512;
wire n_652;
wire n_1111;
wire n_1093;
wire n_1031;
wire n_609;
wire n_1041;
wire n_383;
wire n_834;
wire n_765;
wire n_893;
wire n_1015;
wire n_1140;
wire n_891;
wire n_630;
wire n_504;
wire n_511;
wire n_874;
wire n_358;
wire n_1101;
wire n_1106;
wire n_987;
wire n_767;
wire n_993;
wire n_545;
wire n_441;
wire n_860;
wire n_450;
wire n_429;
wire n_948;
wire n_1217;
wire n_628;
wire n_365;
wire n_729;
wire n_1131;
wire n_1084;
wire n_970;
wire n_911;
wire n_513;
wire n_1094;
wire n_560;
wire n_340;
wire n_1044;
wire n_1205;
wire n_346;
wire n_1209;
wire n_495;
wire n_602;
wire n_574;
wire n_879;
wire n_623;
wire n_405;
wire n_824;
wire n_359;
wire n_490;
wire n_996;
wire n_921;
wire n_572;
wire n_366;
wire n_815;
wire n_1037;
wire n_1080;
wire n_426;
wire n_1082;
wire n_589;
wire n_716;
wire n_562;
wire n_952;
wire n_1229;
wire n_391;
wire n_701;
wire n_1023;
wire n_645;
wire n_539;
wire n_803;
wire n_1092;
wire n_531;
wire n_890;
wire n_764;
wire n_1056;
wire n_960;
wire n_1123;
wire n_1047;
wire n_634;
wire n_348;
wire n_1029;
wire n_925;
wire n_1206;
wire n_424;
wire n_950;
wire n_380;
wire n_419;
wire n_444;
wire n_1060;
wire n_1141;
wire n_389;
wire n_418;
wire n_912;
wire n_968;
wire n_451;
wire n_619;
wire n_408;
wire n_376;
wire n_967;
wire n_1139;
wire n_515;
wire n_351;
wire n_885;
wire n_397;
wire n_483;
wire n_683;
wire n_1057;
wire n_1051;
wire n_1085;
wire n_1066;
wire n_721;
wire n_1157;
wire n_841;
wire n_1050;
wire n_802;
wire n_983;
wire n_873;
wire n_378;
wire n_1112;
wire n_762;
wire n_690;
wire n_583;
wire n_1203;
wire n_821;
wire n_1179;
wire n_621;
wire n_753;
wire n_455;
wire n_1048;
wire n_385;
wire n_507;
wire n_1228;
wire n_972;
wire n_692;
wire n_820;
wire n_1200;
wire n_1185;
wire n_991;
wire n_828;
wire n_779;
wire n_576;
wire n_1143;
wire n_804;
wire n_537;
wire n_945;
wire n_492;
wire n_943;
wire n_341;
wire n_992;
wire n_543;
wire n_842;
wire n_650;
wire n_984;
wire n_694;
wire n_883;
wire n_470;
wire n_449;
wire n_1214;
wire n_900;
wire n_856;
wire n_918;
wire n_942;
wire n_1147;
wire n_1077;
wire n_540;
wire n_618;
wire n_896;
wire n_356;
wire n_894;
wire n_831;
wire n_964;
wire n_1096;
wire n_833;
wire n_988;
wire n_814;
wire n_1201;
wire n_1114;
wire n_655;
wire n_669;
wire n_472;
wire n_1176;
wire n_387;
wire n_1149;
wire n_398;
wire n_635;
wire n_763;
wire n_1020;
wire n_1062;
wire n_1219;
wire n_1204;
wire n_1035;
wire n_555;
wire n_783;
wire n_1188;
wire n_661;
wire n_849;
wire n_336;
wire n_584;
wire n_681;
wire n_430;
wire n_510;
wire n_830;
wire n_801;
wire n_875;
wire n_357;
wire n_1110;
wire n_445;
wire n_749;
wire n_1134;
wire n_717;
wire n_939;
wire n_482;
wire n_1088;
wire n_588;
wire n_1173;
wire n_789;
wire n_1232;
wire n_734;
wire n_638;
wire n_866;
wire n_969;
wire n_1019;
wire n_1105;
wire n_577;
wire n_338;
wire n_693;
wire n_836;
wire n_990;
wire n_975;
wire n_567;
wire n_778;
wire n_1122;
wire n_458;
wire n_770;
wire n_1102;
wire n_711;
wire n_1187;
wire n_1164;
wire n_489;
wire n_1174;
wire n_617;
wire n_876;
wire n_1190;
wire n_601;
wire n_917;
wire n_966;
wire n_1116;
wire n_1212;
wire n_726;
wire n_982;
wire n_818;
wire n_861;
wire n_1183;
wire n_899;
wire n_774;
wire n_1059;
wire n_1133;
wire n_557;
wire n_1005;
wire n_607;
wire n_1003;
wire n_679;
wire n_710;
wire n_527;
wire n_1168;
wire n_707;
wire n_937;
wire n_393;
wire n_487;
wire n_665;
wire n_421;
wire n_910;
wire n_768;
wire n_1136;
wire n_754;
wire n_1125;
wire n_410;
wire n_708;
wire n_529;
wire n_735;
wire n_1109;
wire n_895;
wire n_427;
wire n_791;
wire n_732;
wire n_808;
wire n_797;
wire n_1025;
wire n_500;
wire n_1067;
wire n_435;
wire n_766;
wire n_541;
wire n_538;
wire n_1117;
wire n_799;
wire n_687;
wire n_715;
wire n_1213;
wire n_536;
wire n_872;
wire n_594;
wire n_1155;
wire n_1011;
wire n_1184;
wire n_985;
wire n_869;
wire n_810;
wire n_416;
wire n_827;
wire n_401;
wire n_626;
wire n_1144;
wire n_1137;
wire n_1170;
wire n_676;
wire n_653;
wire n_642;
wire n_855;
wire n_1178;
wire n_850;
wire n_684;
wire n_664;
wire n_503;
wire n_605;
wire n_353;
wire n_620;
wire n_643;
wire n_916;
wire n_1081;
wire n_493;
wire n_1235;
wire n_703;
wire n_698;
wire n_980;
wire n_1115;
wire n_780;
wire n_998;
wire n_467;
wire n_1227;
wire n_840;
wire n_501;
wire n_823;
wire n_725;
wire n_672;
wire n_581;
wire n_382;
wire n_554;
wire n_898;
wire n_1013;
wire n_718;
wire n_1120;
wire n_719;
wire n_443;
wire n_714;
wire n_909;
wire n_997;
wire n_932;
wire n_612;
wire n_788;
wire n_559;
wire n_825;
wire n_508;
wire n_506;
wire n_737;
wire n_986;
wire n_509;
wire n_1192;
wire n_1024;
wire n_1063;
wire n_733;
wire n_941;
wire n_981;
wire n_867;
wire n_587;
wire n_792;
wire n_756;
wire n_399;
wire n_1238;
wire n_548;
wire n_812;
wire n_518;
wire n_505;
wire n_752;
wire n_905;
wire n_1108;
wire n_782;
wire n_1100;
wire n_862;
wire n_760;
wire n_381;
wire n_390;
wire n_481;
wire n_769;
wire n_1046;
wire n_934;
wire n_826;
wire n_886;
wire n_1221;
wire n_654;
wire n_1172;
wire n_379;
wire n_428;
wire n_570;
wire n_853;
wire n_377;
wire n_751;
wire n_786;
wire n_1083;
wire n_1142;
wire n_1129;
wire n_392;
wire n_704;
wire n_787;
wire n_961;
wire n_771;
wire n_1225;
wire n_522;
wire n_400;
wire n_930;
wire n_622;
wire n_1087;
wire n_386;
wire n_994;
wire n_848;
wire n_1223;
wire n_682;
wire n_922;
wire n_816;
wire n_591;
wire n_631;
wire n_479;
wire n_432;
wire n_839;
wire n_1210;
wire n_369;
wire n_871;
wire n_598;
wire n_685;
wire n_608;
wire n_928;
wire n_772;
wire n_499;
wire n_517;
wire n_413;
wire n_402;
wire n_1086;
wire n_796;
wire n_1012;
wire n_903;
wire n_740;
wire n_384;
wire n_1061;
wire n_333;
wire n_462;
wire n_1193;
wire n_1113;
wire n_1226;
wire n_722;
wire n_844;
wire n_471;
wire n_852;
wire n_1028;
wire n_781;
wire n_474;
wire n_542;
wire n_463;
wire n_595;
wire n_502;
wire n_466;
wire n_420;
wire n_632;
wire n_699;
wire n_979;
wire n_846;
wire n_465;
wire n_362;
wire n_585;
wire n_616;
wire n_745;
wire n_1103;
wire n_648;
wire n_1076;
wire n_1091;
wire n_494;
wire n_641;
wire n_730;
wire n_354;
wire n_575;
wire n_480;
wire n_425;
wire n_795;
wire n_695;
wire n_656;
wire n_1220;
wire n_437;
wire n_453;
wire n_403;
wire n_1130;
wire n_720;
wire n_863;
wire n_805;
wire n_712;
wire n_1042;
wire n_412;
wire n_657;
wire n_644;
wire n_1160;
wire n_491;
wire n_1074;
wire n_566;
wire n_565;
wire n_597;
wire n_1181;
wire n_1196;
wire n_651;
wire n_334;
wire n_811;
wire n_807;
wire n_835;
wire n_666;
wire n_1026;
wire n_1234;
wire n_364;
wire n_1138;
wire n_927;
wire n_1089;
wire n_1004;
wire n_1186;
wire n_1032;
wire n_1018;
wire n_438;
wire n_713;
wire n_904;
wire n_1180;
wire n_533;

CKINVDCx5p33_ASAP7_75t_R g332 ( 
.A(n_194),
.Y(n_332)
);

CKINVDCx5p33_ASAP7_75t_R g333 ( 
.A(n_128),
.Y(n_333)
);

BUFx3_ASAP7_75t_L g334 ( 
.A(n_72),
.Y(n_334)
);

CKINVDCx5p33_ASAP7_75t_R g335 ( 
.A(n_134),
.Y(n_335)
);

INVxp67_ASAP7_75t_L g336 ( 
.A(n_11),
.Y(n_336)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_144),
.Y(n_337)
);

CKINVDCx5p33_ASAP7_75t_R g338 ( 
.A(n_266),
.Y(n_338)
);

INVx1_ASAP7_75t_SL g339 ( 
.A(n_262),
.Y(n_339)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_301),
.Y(n_340)
);

CKINVDCx5p33_ASAP7_75t_R g341 ( 
.A(n_253),
.Y(n_341)
);

BUFx2_ASAP7_75t_SL g342 ( 
.A(n_209),
.Y(n_342)
);

CKINVDCx5p33_ASAP7_75t_R g343 ( 
.A(n_305),
.Y(n_343)
);

INVx2_ASAP7_75t_L g344 ( 
.A(n_38),
.Y(n_344)
);

CKINVDCx5p33_ASAP7_75t_R g345 ( 
.A(n_32),
.Y(n_345)
);

INVx1_ASAP7_75t_L g346 ( 
.A(n_6),
.Y(n_346)
);

CKINVDCx5p33_ASAP7_75t_R g347 ( 
.A(n_193),
.Y(n_347)
);

CKINVDCx5p33_ASAP7_75t_R g348 ( 
.A(n_274),
.Y(n_348)
);

CKINVDCx5p33_ASAP7_75t_R g349 ( 
.A(n_250),
.Y(n_349)
);

CKINVDCx5p33_ASAP7_75t_R g350 ( 
.A(n_170),
.Y(n_350)
);

INVx1_ASAP7_75t_L g351 ( 
.A(n_57),
.Y(n_351)
);

INVx1_ASAP7_75t_SL g352 ( 
.A(n_242),
.Y(n_352)
);

CKINVDCx5p33_ASAP7_75t_R g353 ( 
.A(n_317),
.Y(n_353)
);

CKINVDCx5p33_ASAP7_75t_R g354 ( 
.A(n_55),
.Y(n_354)
);

HB1xp67_ASAP7_75t_L g355 ( 
.A(n_183),
.Y(n_355)
);

INVx2_ASAP7_75t_L g356 ( 
.A(n_184),
.Y(n_356)
);

CKINVDCx5p33_ASAP7_75t_R g357 ( 
.A(n_230),
.Y(n_357)
);

CKINVDCx5p33_ASAP7_75t_R g358 ( 
.A(n_91),
.Y(n_358)
);

INVx1_ASAP7_75t_L g359 ( 
.A(n_320),
.Y(n_359)
);

CKINVDCx5p33_ASAP7_75t_R g360 ( 
.A(n_64),
.Y(n_360)
);

CKINVDCx5p33_ASAP7_75t_R g361 ( 
.A(n_119),
.Y(n_361)
);

INVx1_ASAP7_75t_L g362 ( 
.A(n_16),
.Y(n_362)
);

BUFx3_ASAP7_75t_L g363 ( 
.A(n_24),
.Y(n_363)
);

CKINVDCx5p33_ASAP7_75t_R g364 ( 
.A(n_201),
.Y(n_364)
);

INVx1_ASAP7_75t_L g365 ( 
.A(n_34),
.Y(n_365)
);

BUFx10_ASAP7_75t_L g366 ( 
.A(n_312),
.Y(n_366)
);

CKINVDCx5p33_ASAP7_75t_R g367 ( 
.A(n_319),
.Y(n_367)
);

CKINVDCx5p33_ASAP7_75t_R g368 ( 
.A(n_27),
.Y(n_368)
);

CKINVDCx16_ASAP7_75t_R g369 ( 
.A(n_240),
.Y(n_369)
);

CKINVDCx5p33_ASAP7_75t_R g370 ( 
.A(n_143),
.Y(n_370)
);

CKINVDCx5p33_ASAP7_75t_R g371 ( 
.A(n_30),
.Y(n_371)
);

INVx1_ASAP7_75t_L g372 ( 
.A(n_152),
.Y(n_372)
);

INVx2_ASAP7_75t_L g373 ( 
.A(n_314),
.Y(n_373)
);

INVxp33_ASAP7_75t_SL g374 ( 
.A(n_155),
.Y(n_374)
);

BUFx10_ASAP7_75t_L g375 ( 
.A(n_115),
.Y(n_375)
);

CKINVDCx5p33_ASAP7_75t_R g376 ( 
.A(n_110),
.Y(n_376)
);

CKINVDCx5p33_ASAP7_75t_R g377 ( 
.A(n_4),
.Y(n_377)
);

CKINVDCx5p33_ASAP7_75t_R g378 ( 
.A(n_310),
.Y(n_378)
);

INVx1_ASAP7_75t_L g379 ( 
.A(n_5),
.Y(n_379)
);

CKINVDCx20_ASAP7_75t_R g380 ( 
.A(n_239),
.Y(n_380)
);

CKINVDCx20_ASAP7_75t_R g381 ( 
.A(n_59),
.Y(n_381)
);

CKINVDCx5p33_ASAP7_75t_R g382 ( 
.A(n_286),
.Y(n_382)
);

INVx1_ASAP7_75t_SL g383 ( 
.A(n_73),
.Y(n_383)
);

INVx1_ASAP7_75t_L g384 ( 
.A(n_225),
.Y(n_384)
);

CKINVDCx5p33_ASAP7_75t_R g385 ( 
.A(n_197),
.Y(n_385)
);

INVx2_ASAP7_75t_L g386 ( 
.A(n_185),
.Y(n_386)
);

CKINVDCx5p33_ASAP7_75t_R g387 ( 
.A(n_123),
.Y(n_387)
);

CKINVDCx5p33_ASAP7_75t_R g388 ( 
.A(n_200),
.Y(n_388)
);

BUFx6f_ASAP7_75t_L g389 ( 
.A(n_298),
.Y(n_389)
);

CKINVDCx5p33_ASAP7_75t_R g390 ( 
.A(n_112),
.Y(n_390)
);

CKINVDCx5p33_ASAP7_75t_R g391 ( 
.A(n_151),
.Y(n_391)
);

CKINVDCx5p33_ASAP7_75t_R g392 ( 
.A(n_148),
.Y(n_392)
);

INVx1_ASAP7_75t_L g393 ( 
.A(n_179),
.Y(n_393)
);

INVx1_ASAP7_75t_L g394 ( 
.A(n_39),
.Y(n_394)
);

INVx1_ASAP7_75t_L g395 ( 
.A(n_324),
.Y(n_395)
);

CKINVDCx5p33_ASAP7_75t_R g396 ( 
.A(n_133),
.Y(n_396)
);

BUFx10_ASAP7_75t_L g397 ( 
.A(n_2),
.Y(n_397)
);

CKINVDCx5p33_ASAP7_75t_R g398 ( 
.A(n_157),
.Y(n_398)
);

CKINVDCx5p33_ASAP7_75t_R g399 ( 
.A(n_63),
.Y(n_399)
);

CKINVDCx5p33_ASAP7_75t_R g400 ( 
.A(n_265),
.Y(n_400)
);

CKINVDCx5p33_ASAP7_75t_R g401 ( 
.A(n_279),
.Y(n_401)
);

CKINVDCx5p33_ASAP7_75t_R g402 ( 
.A(n_90),
.Y(n_402)
);

CKINVDCx20_ASAP7_75t_R g403 ( 
.A(n_273),
.Y(n_403)
);

INVx1_ASAP7_75t_L g404 ( 
.A(n_145),
.Y(n_404)
);

INVx2_ASAP7_75t_L g405 ( 
.A(n_294),
.Y(n_405)
);

INVx1_ASAP7_75t_L g406 ( 
.A(n_101),
.Y(n_406)
);

CKINVDCx5p33_ASAP7_75t_R g407 ( 
.A(n_211),
.Y(n_407)
);

CKINVDCx5p33_ASAP7_75t_R g408 ( 
.A(n_249),
.Y(n_408)
);

INVx1_ASAP7_75t_SL g409 ( 
.A(n_237),
.Y(n_409)
);

INVx2_ASAP7_75t_L g410 ( 
.A(n_236),
.Y(n_410)
);

CKINVDCx5p33_ASAP7_75t_R g411 ( 
.A(n_223),
.Y(n_411)
);

CKINVDCx5p33_ASAP7_75t_R g412 ( 
.A(n_244),
.Y(n_412)
);

INVx2_ASAP7_75t_SL g413 ( 
.A(n_280),
.Y(n_413)
);

INVx1_ASAP7_75t_L g414 ( 
.A(n_173),
.Y(n_414)
);

CKINVDCx5p33_ASAP7_75t_R g415 ( 
.A(n_272),
.Y(n_415)
);

CKINVDCx20_ASAP7_75t_R g416 ( 
.A(n_166),
.Y(n_416)
);

CKINVDCx5p33_ASAP7_75t_R g417 ( 
.A(n_214),
.Y(n_417)
);

CKINVDCx5p33_ASAP7_75t_R g418 ( 
.A(n_109),
.Y(n_418)
);

CKINVDCx5p33_ASAP7_75t_R g419 ( 
.A(n_330),
.Y(n_419)
);

CKINVDCx5p33_ASAP7_75t_R g420 ( 
.A(n_276),
.Y(n_420)
);

INVx1_ASAP7_75t_L g421 ( 
.A(n_247),
.Y(n_421)
);

CKINVDCx5p33_ASAP7_75t_R g422 ( 
.A(n_315),
.Y(n_422)
);

CKINVDCx5p33_ASAP7_75t_R g423 ( 
.A(n_231),
.Y(n_423)
);

CKINVDCx5p33_ASAP7_75t_R g424 ( 
.A(n_313),
.Y(n_424)
);

INVx1_ASAP7_75t_L g425 ( 
.A(n_259),
.Y(n_425)
);

INVx1_ASAP7_75t_L g426 ( 
.A(n_297),
.Y(n_426)
);

CKINVDCx5p33_ASAP7_75t_R g427 ( 
.A(n_178),
.Y(n_427)
);

CKINVDCx5p33_ASAP7_75t_R g428 ( 
.A(n_238),
.Y(n_428)
);

CKINVDCx5p33_ASAP7_75t_R g429 ( 
.A(n_227),
.Y(n_429)
);

CKINVDCx5p33_ASAP7_75t_R g430 ( 
.A(n_11),
.Y(n_430)
);

CKINVDCx5p33_ASAP7_75t_R g431 ( 
.A(n_160),
.Y(n_431)
);

CKINVDCx5p33_ASAP7_75t_R g432 ( 
.A(n_186),
.Y(n_432)
);

INVx1_ASAP7_75t_L g433 ( 
.A(n_191),
.Y(n_433)
);

CKINVDCx5p33_ASAP7_75t_R g434 ( 
.A(n_177),
.Y(n_434)
);

CKINVDCx5p33_ASAP7_75t_R g435 ( 
.A(n_52),
.Y(n_435)
);

INVx1_ASAP7_75t_L g436 ( 
.A(n_245),
.Y(n_436)
);

CKINVDCx20_ASAP7_75t_R g437 ( 
.A(n_210),
.Y(n_437)
);

CKINVDCx5p33_ASAP7_75t_R g438 ( 
.A(n_86),
.Y(n_438)
);

INVx2_ASAP7_75t_L g439 ( 
.A(n_203),
.Y(n_439)
);

CKINVDCx5p33_ASAP7_75t_R g440 ( 
.A(n_141),
.Y(n_440)
);

INVx1_ASAP7_75t_SL g441 ( 
.A(n_229),
.Y(n_441)
);

CKINVDCx5p33_ASAP7_75t_R g442 ( 
.A(n_41),
.Y(n_442)
);

CKINVDCx14_ASAP7_75t_R g443 ( 
.A(n_175),
.Y(n_443)
);

INVx1_ASAP7_75t_L g444 ( 
.A(n_278),
.Y(n_444)
);

INVx1_ASAP7_75t_L g445 ( 
.A(n_129),
.Y(n_445)
);

CKINVDCx20_ASAP7_75t_R g446 ( 
.A(n_327),
.Y(n_446)
);

CKINVDCx16_ASAP7_75t_R g447 ( 
.A(n_5),
.Y(n_447)
);

CKINVDCx5p33_ASAP7_75t_R g448 ( 
.A(n_31),
.Y(n_448)
);

CKINVDCx5p33_ASAP7_75t_R g449 ( 
.A(n_251),
.Y(n_449)
);

CKINVDCx5p33_ASAP7_75t_R g450 ( 
.A(n_147),
.Y(n_450)
);

CKINVDCx5p33_ASAP7_75t_R g451 ( 
.A(n_199),
.Y(n_451)
);

CKINVDCx5p33_ASAP7_75t_R g452 ( 
.A(n_292),
.Y(n_452)
);

CKINVDCx20_ASAP7_75t_R g453 ( 
.A(n_76),
.Y(n_453)
);

BUFx2_ASAP7_75t_L g454 ( 
.A(n_99),
.Y(n_454)
);

CKINVDCx5p33_ASAP7_75t_R g455 ( 
.A(n_84),
.Y(n_455)
);

INVx1_ASAP7_75t_L g456 ( 
.A(n_26),
.Y(n_456)
);

INVx1_ASAP7_75t_L g457 ( 
.A(n_118),
.Y(n_457)
);

CKINVDCx20_ASAP7_75t_R g458 ( 
.A(n_132),
.Y(n_458)
);

CKINVDCx20_ASAP7_75t_R g459 ( 
.A(n_2),
.Y(n_459)
);

CKINVDCx5p33_ASAP7_75t_R g460 ( 
.A(n_206),
.Y(n_460)
);

CKINVDCx5p33_ASAP7_75t_R g461 ( 
.A(n_15),
.Y(n_461)
);

CKINVDCx5p33_ASAP7_75t_R g462 ( 
.A(n_171),
.Y(n_462)
);

CKINVDCx5p33_ASAP7_75t_R g463 ( 
.A(n_331),
.Y(n_463)
);

INVx1_ASAP7_75t_SL g464 ( 
.A(n_78),
.Y(n_464)
);

INVx2_ASAP7_75t_L g465 ( 
.A(n_138),
.Y(n_465)
);

CKINVDCx20_ASAP7_75t_R g466 ( 
.A(n_208),
.Y(n_466)
);

CKINVDCx5p33_ASAP7_75t_R g467 ( 
.A(n_159),
.Y(n_467)
);

BUFx3_ASAP7_75t_L g468 ( 
.A(n_243),
.Y(n_468)
);

CKINVDCx20_ASAP7_75t_R g469 ( 
.A(n_174),
.Y(n_469)
);

CKINVDCx5p33_ASAP7_75t_R g470 ( 
.A(n_267),
.Y(n_470)
);

CKINVDCx20_ASAP7_75t_R g471 ( 
.A(n_6),
.Y(n_471)
);

CKINVDCx14_ASAP7_75t_R g472 ( 
.A(n_270),
.Y(n_472)
);

CKINVDCx20_ASAP7_75t_R g473 ( 
.A(n_1),
.Y(n_473)
);

CKINVDCx5p33_ASAP7_75t_R g474 ( 
.A(n_300),
.Y(n_474)
);

INVx1_ASAP7_75t_L g475 ( 
.A(n_311),
.Y(n_475)
);

CKINVDCx5p33_ASAP7_75t_R g476 ( 
.A(n_220),
.Y(n_476)
);

CKINVDCx5p33_ASAP7_75t_R g477 ( 
.A(n_43),
.Y(n_477)
);

BUFx6f_ASAP7_75t_L g478 ( 
.A(n_7),
.Y(n_478)
);

INVxp67_ASAP7_75t_SL g479 ( 
.A(n_303),
.Y(n_479)
);

INVx1_ASAP7_75t_L g480 ( 
.A(n_283),
.Y(n_480)
);

CKINVDCx5p33_ASAP7_75t_R g481 ( 
.A(n_309),
.Y(n_481)
);

CKINVDCx5p33_ASAP7_75t_R g482 ( 
.A(n_328),
.Y(n_482)
);

CKINVDCx20_ASAP7_75t_R g483 ( 
.A(n_82),
.Y(n_483)
);

CKINVDCx5p33_ASAP7_75t_R g484 ( 
.A(n_28),
.Y(n_484)
);

CKINVDCx5p33_ASAP7_75t_R g485 ( 
.A(n_61),
.Y(n_485)
);

CKINVDCx5p33_ASAP7_75t_R g486 ( 
.A(n_103),
.Y(n_486)
);

INVx1_ASAP7_75t_SL g487 ( 
.A(n_102),
.Y(n_487)
);

INVx1_ASAP7_75t_L g488 ( 
.A(n_45),
.Y(n_488)
);

CKINVDCx5p33_ASAP7_75t_R g489 ( 
.A(n_168),
.Y(n_489)
);

CKINVDCx5p33_ASAP7_75t_R g490 ( 
.A(n_135),
.Y(n_490)
);

CKINVDCx5p33_ASAP7_75t_R g491 ( 
.A(n_105),
.Y(n_491)
);

CKINVDCx5p33_ASAP7_75t_R g492 ( 
.A(n_321),
.Y(n_492)
);

INVx1_ASAP7_75t_SL g493 ( 
.A(n_121),
.Y(n_493)
);

CKINVDCx5p33_ASAP7_75t_R g494 ( 
.A(n_25),
.Y(n_494)
);

CKINVDCx5p33_ASAP7_75t_R g495 ( 
.A(n_88),
.Y(n_495)
);

INVx1_ASAP7_75t_L g496 ( 
.A(n_322),
.Y(n_496)
);

INVxp67_ASAP7_75t_L g497 ( 
.A(n_232),
.Y(n_497)
);

CKINVDCx5p33_ASAP7_75t_R g498 ( 
.A(n_19),
.Y(n_498)
);

CKINVDCx16_ASAP7_75t_R g499 ( 
.A(n_156),
.Y(n_499)
);

CKINVDCx5p33_ASAP7_75t_R g500 ( 
.A(n_154),
.Y(n_500)
);

INVx1_ASAP7_75t_L g501 ( 
.A(n_306),
.Y(n_501)
);

CKINVDCx5p33_ASAP7_75t_R g502 ( 
.A(n_18),
.Y(n_502)
);

INVx1_ASAP7_75t_L g503 ( 
.A(n_4),
.Y(n_503)
);

CKINVDCx5p33_ASAP7_75t_R g504 ( 
.A(n_95),
.Y(n_504)
);

CKINVDCx5p33_ASAP7_75t_R g505 ( 
.A(n_252),
.Y(n_505)
);

CKINVDCx5p33_ASAP7_75t_R g506 ( 
.A(n_285),
.Y(n_506)
);

CKINVDCx5p33_ASAP7_75t_R g507 ( 
.A(n_68),
.Y(n_507)
);

CKINVDCx20_ASAP7_75t_R g508 ( 
.A(n_167),
.Y(n_508)
);

CKINVDCx5p33_ASAP7_75t_R g509 ( 
.A(n_212),
.Y(n_509)
);

CKINVDCx5p33_ASAP7_75t_R g510 ( 
.A(n_16),
.Y(n_510)
);

CKINVDCx20_ASAP7_75t_R g511 ( 
.A(n_241),
.Y(n_511)
);

CKINVDCx5p33_ASAP7_75t_R g512 ( 
.A(n_326),
.Y(n_512)
);

INVx1_ASAP7_75t_SL g513 ( 
.A(n_113),
.Y(n_513)
);

CKINVDCx5p33_ASAP7_75t_R g514 ( 
.A(n_85),
.Y(n_514)
);

CKINVDCx5p33_ASAP7_75t_R g515 ( 
.A(n_165),
.Y(n_515)
);

CKINVDCx5p33_ASAP7_75t_R g516 ( 
.A(n_325),
.Y(n_516)
);

CKINVDCx5p33_ASAP7_75t_R g517 ( 
.A(n_120),
.Y(n_517)
);

CKINVDCx5p33_ASAP7_75t_R g518 ( 
.A(n_71),
.Y(n_518)
);

INVx2_ASAP7_75t_L g519 ( 
.A(n_221),
.Y(n_519)
);

CKINVDCx5p33_ASAP7_75t_R g520 ( 
.A(n_87),
.Y(n_520)
);

CKINVDCx5p33_ASAP7_75t_R g521 ( 
.A(n_146),
.Y(n_521)
);

CKINVDCx5p33_ASAP7_75t_R g522 ( 
.A(n_104),
.Y(n_522)
);

CKINVDCx14_ASAP7_75t_R g523 ( 
.A(n_295),
.Y(n_523)
);

CKINVDCx5p33_ASAP7_75t_R g524 ( 
.A(n_122),
.Y(n_524)
);

INVx1_ASAP7_75t_L g525 ( 
.A(n_281),
.Y(n_525)
);

BUFx3_ASAP7_75t_L g526 ( 
.A(n_188),
.Y(n_526)
);

BUFx3_ASAP7_75t_L g527 ( 
.A(n_58),
.Y(n_527)
);

CKINVDCx5p33_ASAP7_75t_R g528 ( 
.A(n_222),
.Y(n_528)
);

CKINVDCx5p33_ASAP7_75t_R g529 ( 
.A(n_49),
.Y(n_529)
);

INVx1_ASAP7_75t_L g530 ( 
.A(n_307),
.Y(n_530)
);

CKINVDCx5p33_ASAP7_75t_R g531 ( 
.A(n_195),
.Y(n_531)
);

CKINVDCx5p33_ASAP7_75t_R g532 ( 
.A(n_51),
.Y(n_532)
);

CKINVDCx5p33_ASAP7_75t_R g533 ( 
.A(n_304),
.Y(n_533)
);

INVx2_ASAP7_75t_L g534 ( 
.A(n_308),
.Y(n_534)
);

INVx1_ASAP7_75t_L g535 ( 
.A(n_40),
.Y(n_535)
);

CKINVDCx20_ASAP7_75t_R g536 ( 
.A(n_111),
.Y(n_536)
);

CKINVDCx5p33_ASAP7_75t_R g537 ( 
.A(n_1),
.Y(n_537)
);

INVx4_ASAP7_75t_R g538 ( 
.A(n_67),
.Y(n_538)
);

BUFx3_ASAP7_75t_L g539 ( 
.A(n_44),
.Y(n_539)
);

INVx1_ASAP7_75t_L g540 ( 
.A(n_106),
.Y(n_540)
);

CKINVDCx5p33_ASAP7_75t_R g541 ( 
.A(n_282),
.Y(n_541)
);

INVx2_ASAP7_75t_L g542 ( 
.A(n_10),
.Y(n_542)
);

INVx1_ASAP7_75t_SL g543 ( 
.A(n_3),
.Y(n_543)
);

CKINVDCx20_ASAP7_75t_R g544 ( 
.A(n_22),
.Y(n_544)
);

INVx1_ASAP7_75t_L g545 ( 
.A(n_478),
.Y(n_545)
);

CKINVDCx5p33_ASAP7_75t_R g546 ( 
.A(n_332),
.Y(n_546)
);

CKINVDCx20_ASAP7_75t_R g547 ( 
.A(n_380),
.Y(n_547)
);

INVxp67_ASAP7_75t_SL g548 ( 
.A(n_355),
.Y(n_548)
);

CKINVDCx5p33_ASAP7_75t_R g549 ( 
.A(n_333),
.Y(n_549)
);

INVx1_ASAP7_75t_L g550 ( 
.A(n_478),
.Y(n_550)
);

INVxp67_ASAP7_75t_L g551 ( 
.A(n_397),
.Y(n_551)
);

INVx1_ASAP7_75t_L g552 ( 
.A(n_478),
.Y(n_552)
);

CKINVDCx20_ASAP7_75t_R g553 ( 
.A(n_381),
.Y(n_553)
);

CKINVDCx5p33_ASAP7_75t_R g554 ( 
.A(n_335),
.Y(n_554)
);

CKINVDCx20_ASAP7_75t_R g555 ( 
.A(n_403),
.Y(n_555)
);

CKINVDCx5p33_ASAP7_75t_R g556 ( 
.A(n_338),
.Y(n_556)
);

INVx1_ASAP7_75t_L g557 ( 
.A(n_478),
.Y(n_557)
);

CKINVDCx5p33_ASAP7_75t_R g558 ( 
.A(n_341),
.Y(n_558)
);

INVx1_ASAP7_75t_L g559 ( 
.A(n_346),
.Y(n_559)
);

NOR2xp33_ASAP7_75t_L g560 ( 
.A(n_454),
.B(n_0),
.Y(n_560)
);

INVx1_ASAP7_75t_L g561 ( 
.A(n_362),
.Y(n_561)
);

INVx1_ASAP7_75t_L g562 ( 
.A(n_379),
.Y(n_562)
);

INVx1_ASAP7_75t_L g563 ( 
.A(n_503),
.Y(n_563)
);

CKINVDCx20_ASAP7_75t_R g564 ( 
.A(n_416),
.Y(n_564)
);

INVxp67_ASAP7_75t_L g565 ( 
.A(n_397),
.Y(n_565)
);

INVx1_ASAP7_75t_L g566 ( 
.A(n_334),
.Y(n_566)
);

CKINVDCx5p33_ASAP7_75t_R g567 ( 
.A(n_343),
.Y(n_567)
);

CKINVDCx5p33_ASAP7_75t_R g568 ( 
.A(n_345),
.Y(n_568)
);

CKINVDCx20_ASAP7_75t_R g569 ( 
.A(n_437),
.Y(n_569)
);

INVxp67_ASAP7_75t_SL g570 ( 
.A(n_334),
.Y(n_570)
);

CKINVDCx5p33_ASAP7_75t_R g571 ( 
.A(n_347),
.Y(n_571)
);

CKINVDCx5p33_ASAP7_75t_R g572 ( 
.A(n_348),
.Y(n_572)
);

INVx1_ASAP7_75t_L g573 ( 
.A(n_363),
.Y(n_573)
);

INVx1_ASAP7_75t_L g574 ( 
.A(n_363),
.Y(n_574)
);

NOR2xp33_ASAP7_75t_L g575 ( 
.A(n_497),
.B(n_339),
.Y(n_575)
);

CKINVDCx5p33_ASAP7_75t_R g576 ( 
.A(n_349),
.Y(n_576)
);

CKINVDCx5p33_ASAP7_75t_R g577 ( 
.A(n_350),
.Y(n_577)
);

INVx1_ASAP7_75t_L g578 ( 
.A(n_468),
.Y(n_578)
);

INVx1_ASAP7_75t_L g579 ( 
.A(n_468),
.Y(n_579)
);

INVx1_ASAP7_75t_L g580 ( 
.A(n_526),
.Y(n_580)
);

INVx1_ASAP7_75t_L g581 ( 
.A(n_526),
.Y(n_581)
);

INVxp67_ASAP7_75t_SL g582 ( 
.A(n_527),
.Y(n_582)
);

INVx2_ASAP7_75t_L g583 ( 
.A(n_542),
.Y(n_583)
);

INVxp67_ASAP7_75t_SL g584 ( 
.A(n_527),
.Y(n_584)
);

INVx2_ASAP7_75t_L g585 ( 
.A(n_389),
.Y(n_585)
);

CKINVDCx5p33_ASAP7_75t_R g586 ( 
.A(n_353),
.Y(n_586)
);

INVx2_ASAP7_75t_L g587 ( 
.A(n_389),
.Y(n_587)
);

CKINVDCx20_ASAP7_75t_R g588 ( 
.A(n_446),
.Y(n_588)
);

CKINVDCx5p33_ASAP7_75t_R g589 ( 
.A(n_354),
.Y(n_589)
);

INVx1_ASAP7_75t_L g590 ( 
.A(n_539),
.Y(n_590)
);

CKINVDCx5p33_ASAP7_75t_R g591 ( 
.A(n_357),
.Y(n_591)
);

CKINVDCx20_ASAP7_75t_R g592 ( 
.A(n_453),
.Y(n_592)
);

CKINVDCx5p33_ASAP7_75t_R g593 ( 
.A(n_358),
.Y(n_593)
);

CKINVDCx20_ASAP7_75t_R g594 ( 
.A(n_458),
.Y(n_594)
);

INVx1_ASAP7_75t_L g595 ( 
.A(n_539),
.Y(n_595)
);

INVx1_ASAP7_75t_L g596 ( 
.A(n_337),
.Y(n_596)
);

CKINVDCx16_ASAP7_75t_R g597 ( 
.A(n_447),
.Y(n_597)
);

HB1xp67_ASAP7_75t_L g598 ( 
.A(n_377),
.Y(n_598)
);

CKINVDCx20_ASAP7_75t_R g599 ( 
.A(n_466),
.Y(n_599)
);

INVx1_ASAP7_75t_L g600 ( 
.A(n_340),
.Y(n_600)
);

CKINVDCx5p33_ASAP7_75t_R g601 ( 
.A(n_360),
.Y(n_601)
);

INVx1_ASAP7_75t_L g602 ( 
.A(n_351),
.Y(n_602)
);

CKINVDCx20_ASAP7_75t_R g603 ( 
.A(n_469),
.Y(n_603)
);

INVx1_ASAP7_75t_L g604 ( 
.A(n_359),
.Y(n_604)
);

CKINVDCx20_ASAP7_75t_R g605 ( 
.A(n_483),
.Y(n_605)
);

HB1xp67_ASAP7_75t_L g606 ( 
.A(n_430),
.Y(n_606)
);

CKINVDCx16_ASAP7_75t_R g607 ( 
.A(n_369),
.Y(n_607)
);

INVx1_ASAP7_75t_L g608 ( 
.A(n_365),
.Y(n_608)
);

INVx1_ASAP7_75t_L g609 ( 
.A(n_372),
.Y(n_609)
);

CKINVDCx5p33_ASAP7_75t_R g610 ( 
.A(n_361),
.Y(n_610)
);

INVx1_ASAP7_75t_L g611 ( 
.A(n_384),
.Y(n_611)
);

CKINVDCx5p33_ASAP7_75t_R g612 ( 
.A(n_364),
.Y(n_612)
);

OR2x2_ASAP7_75t_L g613 ( 
.A(n_543),
.B(n_0),
.Y(n_613)
);

INVx1_ASAP7_75t_L g614 ( 
.A(n_393),
.Y(n_614)
);

INVx1_ASAP7_75t_L g615 ( 
.A(n_394),
.Y(n_615)
);

INVxp67_ASAP7_75t_L g616 ( 
.A(n_461),
.Y(n_616)
);

CKINVDCx20_ASAP7_75t_R g617 ( 
.A(n_508),
.Y(n_617)
);

INVx1_ASAP7_75t_L g618 ( 
.A(n_395),
.Y(n_618)
);

CKINVDCx20_ASAP7_75t_R g619 ( 
.A(n_511),
.Y(n_619)
);

CKINVDCx20_ASAP7_75t_R g620 ( 
.A(n_536),
.Y(n_620)
);

INVx1_ASAP7_75t_L g621 ( 
.A(n_404),
.Y(n_621)
);

CKINVDCx5p33_ASAP7_75t_R g622 ( 
.A(n_367),
.Y(n_622)
);

NOR2xp33_ASAP7_75t_L g623 ( 
.A(n_352),
.B(n_3),
.Y(n_623)
);

INVx1_ASAP7_75t_L g624 ( 
.A(n_406),
.Y(n_624)
);

NOR2xp33_ASAP7_75t_L g625 ( 
.A(n_383),
.B(n_409),
.Y(n_625)
);

INVxp67_ASAP7_75t_SL g626 ( 
.A(n_414),
.Y(n_626)
);

CKINVDCx16_ASAP7_75t_R g627 ( 
.A(n_499),
.Y(n_627)
);

CKINVDCx5p33_ASAP7_75t_R g628 ( 
.A(n_368),
.Y(n_628)
);

NOR2xp33_ASAP7_75t_R g629 ( 
.A(n_443),
.B(n_7),
.Y(n_629)
);

INVx1_ASAP7_75t_L g630 ( 
.A(n_421),
.Y(n_630)
);

INVx1_ASAP7_75t_L g631 ( 
.A(n_425),
.Y(n_631)
);

INVx1_ASAP7_75t_L g632 ( 
.A(n_426),
.Y(n_632)
);

CKINVDCx20_ASAP7_75t_R g633 ( 
.A(n_472),
.Y(n_633)
);

HB1xp67_ASAP7_75t_L g634 ( 
.A(n_498),
.Y(n_634)
);

INVx1_ASAP7_75t_L g635 ( 
.A(n_433),
.Y(n_635)
);

CKINVDCx20_ASAP7_75t_R g636 ( 
.A(n_523),
.Y(n_636)
);

HB1xp67_ASAP7_75t_L g637 ( 
.A(n_502),
.Y(n_637)
);

CKINVDCx16_ASAP7_75t_R g638 ( 
.A(n_366),
.Y(n_638)
);

INVxp67_ASAP7_75t_SL g639 ( 
.A(n_436),
.Y(n_639)
);

CKINVDCx5p33_ASAP7_75t_R g640 ( 
.A(n_370),
.Y(n_640)
);

INVx1_ASAP7_75t_SL g641 ( 
.A(n_459),
.Y(n_641)
);

INVxp67_ASAP7_75t_L g642 ( 
.A(n_510),
.Y(n_642)
);

INVx1_ASAP7_75t_L g643 ( 
.A(n_444),
.Y(n_643)
);

INVx1_ASAP7_75t_L g644 ( 
.A(n_445),
.Y(n_644)
);

INVx1_ASAP7_75t_L g645 ( 
.A(n_456),
.Y(n_645)
);

CKINVDCx20_ASAP7_75t_R g646 ( 
.A(n_371),
.Y(n_646)
);

CKINVDCx5p33_ASAP7_75t_R g647 ( 
.A(n_376),
.Y(n_647)
);

NAND2xp5_ASAP7_75t_L g648 ( 
.A(n_413),
.B(n_8),
.Y(n_648)
);

INVx1_ASAP7_75t_L g649 ( 
.A(n_457),
.Y(n_649)
);

CKINVDCx20_ASAP7_75t_R g650 ( 
.A(n_378),
.Y(n_650)
);

CKINVDCx5p33_ASAP7_75t_R g651 ( 
.A(n_382),
.Y(n_651)
);

INVxp67_ASAP7_75t_SL g652 ( 
.A(n_475),
.Y(n_652)
);

INVxp67_ASAP7_75t_L g653 ( 
.A(n_537),
.Y(n_653)
);

CKINVDCx5p33_ASAP7_75t_R g654 ( 
.A(n_385),
.Y(n_654)
);

CKINVDCx20_ASAP7_75t_R g655 ( 
.A(n_387),
.Y(n_655)
);

INVx1_ASAP7_75t_L g656 ( 
.A(n_480),
.Y(n_656)
);

INVxp33_ASAP7_75t_SL g657 ( 
.A(n_388),
.Y(n_657)
);

CKINVDCx5p33_ASAP7_75t_R g658 ( 
.A(n_390),
.Y(n_658)
);

INVxp33_ASAP7_75t_L g659 ( 
.A(n_488),
.Y(n_659)
);

INVx1_ASAP7_75t_L g660 ( 
.A(n_496),
.Y(n_660)
);

CKINVDCx20_ASAP7_75t_R g661 ( 
.A(n_391),
.Y(n_661)
);

INVx1_ASAP7_75t_L g662 ( 
.A(n_501),
.Y(n_662)
);

AND2x6_ASAP7_75t_L g663 ( 
.A(n_585),
.B(n_389),
.Y(n_663)
);

INVx1_ASAP7_75t_L g664 ( 
.A(n_545),
.Y(n_664)
);

NAND2xp5_ASAP7_75t_L g665 ( 
.A(n_625),
.B(n_534),
.Y(n_665)
);

INVx1_ASAP7_75t_L g666 ( 
.A(n_550),
.Y(n_666)
);

CKINVDCx5p33_ASAP7_75t_R g667 ( 
.A(n_546),
.Y(n_667)
);

CKINVDCx5p33_ASAP7_75t_R g668 ( 
.A(n_549),
.Y(n_668)
);

CKINVDCx5p33_ASAP7_75t_R g669 ( 
.A(n_554),
.Y(n_669)
);

CKINVDCx5p33_ASAP7_75t_R g670 ( 
.A(n_556),
.Y(n_670)
);

INVx1_ASAP7_75t_L g671 ( 
.A(n_552),
.Y(n_671)
);

NOR2xp33_ASAP7_75t_L g672 ( 
.A(n_625),
.B(n_374),
.Y(n_672)
);

INVx3_ASAP7_75t_L g673 ( 
.A(n_583),
.Y(n_673)
);

INVx2_ASAP7_75t_L g674 ( 
.A(n_557),
.Y(n_674)
);

CKINVDCx5p33_ASAP7_75t_R g675 ( 
.A(n_558),
.Y(n_675)
);

INVx2_ASAP7_75t_L g676 ( 
.A(n_585),
.Y(n_676)
);

CKINVDCx5p33_ASAP7_75t_R g677 ( 
.A(n_567),
.Y(n_677)
);

CKINVDCx5p33_ASAP7_75t_R g678 ( 
.A(n_568),
.Y(n_678)
);

INVx1_ASAP7_75t_L g679 ( 
.A(n_596),
.Y(n_679)
);

INVx1_ASAP7_75t_SL g680 ( 
.A(n_641),
.Y(n_680)
);

AND2x6_ASAP7_75t_L g681 ( 
.A(n_587),
.B(n_389),
.Y(n_681)
);

AND2x2_ASAP7_75t_L g682 ( 
.A(n_616),
.B(n_366),
.Y(n_682)
);

CKINVDCx20_ASAP7_75t_R g683 ( 
.A(n_547),
.Y(n_683)
);

INVx1_ASAP7_75t_L g684 ( 
.A(n_600),
.Y(n_684)
);

INVx2_ASAP7_75t_L g685 ( 
.A(n_587),
.Y(n_685)
);

INVx1_ASAP7_75t_L g686 ( 
.A(n_602),
.Y(n_686)
);

NOR2xp33_ASAP7_75t_L g687 ( 
.A(n_575),
.B(n_441),
.Y(n_687)
);

INVx1_ASAP7_75t_L g688 ( 
.A(n_604),
.Y(n_688)
);

INVx1_ASAP7_75t_L g689 ( 
.A(n_608),
.Y(n_689)
);

INVx2_ASAP7_75t_L g690 ( 
.A(n_559),
.Y(n_690)
);

INVx2_ASAP7_75t_L g691 ( 
.A(n_561),
.Y(n_691)
);

AND2x2_ASAP7_75t_L g692 ( 
.A(n_642),
.B(n_375),
.Y(n_692)
);

BUFx3_ASAP7_75t_L g693 ( 
.A(n_646),
.Y(n_693)
);

BUFx6f_ASAP7_75t_L g694 ( 
.A(n_562),
.Y(n_694)
);

INVx3_ASAP7_75t_L g695 ( 
.A(n_563),
.Y(n_695)
);

CKINVDCx5p33_ASAP7_75t_R g696 ( 
.A(n_571),
.Y(n_696)
);

CKINVDCx20_ASAP7_75t_R g697 ( 
.A(n_553),
.Y(n_697)
);

CKINVDCx5p33_ASAP7_75t_R g698 ( 
.A(n_572),
.Y(n_698)
);

INVx1_ASAP7_75t_L g699 ( 
.A(n_609),
.Y(n_699)
);

CKINVDCx5p33_ASAP7_75t_R g700 ( 
.A(n_576),
.Y(n_700)
);

AND2x4_ASAP7_75t_L g701 ( 
.A(n_570),
.B(n_479),
.Y(n_701)
);

NAND2xp5_ASAP7_75t_L g702 ( 
.A(n_577),
.B(n_534),
.Y(n_702)
);

INVx2_ASAP7_75t_L g703 ( 
.A(n_611),
.Y(n_703)
);

INVx1_ASAP7_75t_L g704 ( 
.A(n_614),
.Y(n_704)
);

INVx2_ASAP7_75t_L g705 ( 
.A(n_615),
.Y(n_705)
);

INVx3_ASAP7_75t_L g706 ( 
.A(n_618),
.Y(n_706)
);

CKINVDCx5p33_ASAP7_75t_R g707 ( 
.A(n_586),
.Y(n_707)
);

INVx1_ASAP7_75t_L g708 ( 
.A(n_621),
.Y(n_708)
);

INVx1_ASAP7_75t_L g709 ( 
.A(n_624),
.Y(n_709)
);

AND2x4_ASAP7_75t_L g710 ( 
.A(n_582),
.B(n_344),
.Y(n_710)
);

AND2x2_ASAP7_75t_L g711 ( 
.A(n_653),
.B(n_375),
.Y(n_711)
);

INVxp67_ASAP7_75t_L g712 ( 
.A(n_598),
.Y(n_712)
);

INVx1_ASAP7_75t_L g713 ( 
.A(n_630),
.Y(n_713)
);

NOR2xp33_ASAP7_75t_R g714 ( 
.A(n_633),
.B(n_392),
.Y(n_714)
);

INVx1_ASAP7_75t_L g715 ( 
.A(n_631),
.Y(n_715)
);

INVx1_ASAP7_75t_L g716 ( 
.A(n_632),
.Y(n_716)
);

INVx2_ASAP7_75t_L g717 ( 
.A(n_635),
.Y(n_717)
);

INVx2_ASAP7_75t_L g718 ( 
.A(n_662),
.Y(n_718)
);

CKINVDCx20_ASAP7_75t_R g719 ( 
.A(n_555),
.Y(n_719)
);

CKINVDCx5p33_ASAP7_75t_R g720 ( 
.A(n_589),
.Y(n_720)
);

HB1xp67_ASAP7_75t_L g721 ( 
.A(n_597),
.Y(n_721)
);

INVx3_ASAP7_75t_L g722 ( 
.A(n_566),
.Y(n_722)
);

INVx1_ASAP7_75t_L g723 ( 
.A(n_643),
.Y(n_723)
);

NAND2xp5_ASAP7_75t_SL g724 ( 
.A(n_638),
.B(n_464),
.Y(n_724)
);

CKINVDCx5p33_ASAP7_75t_R g725 ( 
.A(n_591),
.Y(n_725)
);

INVx1_ASAP7_75t_L g726 ( 
.A(n_644),
.Y(n_726)
);

NAND2xp5_ASAP7_75t_L g727 ( 
.A(n_593),
.B(n_356),
.Y(n_727)
);

INVx2_ASAP7_75t_L g728 ( 
.A(n_645),
.Y(n_728)
);

INVx1_ASAP7_75t_L g729 ( 
.A(n_649),
.Y(n_729)
);

INVx1_ASAP7_75t_L g730 ( 
.A(n_656),
.Y(n_730)
);

INVx4_ASAP7_75t_L g731 ( 
.A(n_601),
.Y(n_731)
);

OR2x2_ASAP7_75t_L g732 ( 
.A(n_613),
.B(n_336),
.Y(n_732)
);

CKINVDCx20_ASAP7_75t_R g733 ( 
.A(n_564),
.Y(n_733)
);

BUFx6f_ASAP7_75t_L g734 ( 
.A(n_660),
.Y(n_734)
);

NAND2xp5_ASAP7_75t_L g735 ( 
.A(n_610),
.B(n_373),
.Y(n_735)
);

NOR2xp33_ASAP7_75t_R g736 ( 
.A(n_636),
.B(n_396),
.Y(n_736)
);

CKINVDCx20_ASAP7_75t_R g737 ( 
.A(n_569),
.Y(n_737)
);

INVx2_ASAP7_75t_L g738 ( 
.A(n_573),
.Y(n_738)
);

CKINVDCx5p33_ASAP7_75t_R g739 ( 
.A(n_612),
.Y(n_739)
);

INVx1_ASAP7_75t_SL g740 ( 
.A(n_588),
.Y(n_740)
);

AND2x6_ASAP7_75t_L g741 ( 
.A(n_560),
.B(n_386),
.Y(n_741)
);

CKINVDCx5p33_ASAP7_75t_R g742 ( 
.A(n_622),
.Y(n_742)
);

INVx1_ASAP7_75t_L g743 ( 
.A(n_574),
.Y(n_743)
);

INVx2_ASAP7_75t_L g744 ( 
.A(n_578),
.Y(n_744)
);

INVx2_ASAP7_75t_L g745 ( 
.A(n_579),
.Y(n_745)
);

AND2x2_ASAP7_75t_L g746 ( 
.A(n_606),
.B(n_487),
.Y(n_746)
);

CKINVDCx5p33_ASAP7_75t_R g747 ( 
.A(n_628),
.Y(n_747)
);

INVx3_ASAP7_75t_L g748 ( 
.A(n_580),
.Y(n_748)
);

AND2x2_ASAP7_75t_L g749 ( 
.A(n_634),
.B(n_493),
.Y(n_749)
);

INVx1_ASAP7_75t_L g750 ( 
.A(n_581),
.Y(n_750)
);

INVx1_ASAP7_75t_L g751 ( 
.A(n_590),
.Y(n_751)
);

INVx1_ASAP7_75t_L g752 ( 
.A(n_595),
.Y(n_752)
);

NAND2xp5_ASAP7_75t_L g753 ( 
.A(n_672),
.B(n_640),
.Y(n_753)
);

INVx2_ASAP7_75t_L g754 ( 
.A(n_676),
.Y(n_754)
);

INVx1_ASAP7_75t_L g755 ( 
.A(n_679),
.Y(n_755)
);

AND2x2_ASAP7_75t_L g756 ( 
.A(n_687),
.B(n_637),
.Y(n_756)
);

AND2x6_ASAP7_75t_L g757 ( 
.A(n_743),
.B(n_560),
.Y(n_757)
);

BUFx2_ASAP7_75t_L g758 ( 
.A(n_680),
.Y(n_758)
);

INVx1_ASAP7_75t_SL g759 ( 
.A(n_740),
.Y(n_759)
);

HB1xp67_ASAP7_75t_L g760 ( 
.A(n_721),
.Y(n_760)
);

BUFx2_ASAP7_75t_L g761 ( 
.A(n_746),
.Y(n_761)
);

BUFx6f_ASAP7_75t_L g762 ( 
.A(n_734),
.Y(n_762)
);

NAND2xp5_ASAP7_75t_L g763 ( 
.A(n_701),
.B(n_647),
.Y(n_763)
);

AND2x2_ASAP7_75t_L g764 ( 
.A(n_749),
.B(n_607),
.Y(n_764)
);

BUFx2_ASAP7_75t_L g765 ( 
.A(n_712),
.Y(n_765)
);

INVx1_ASAP7_75t_SL g766 ( 
.A(n_683),
.Y(n_766)
);

INVx2_ASAP7_75t_L g767 ( 
.A(n_685),
.Y(n_767)
);

INVx2_ASAP7_75t_L g768 ( 
.A(n_674),
.Y(n_768)
);

INVx1_ASAP7_75t_SL g769 ( 
.A(n_697),
.Y(n_769)
);

NAND2xp5_ASAP7_75t_L g770 ( 
.A(n_701),
.B(n_651),
.Y(n_770)
);

INVx2_ASAP7_75t_L g771 ( 
.A(n_664),
.Y(n_771)
);

INVx2_ASAP7_75t_L g772 ( 
.A(n_666),
.Y(n_772)
);

NOR2xp33_ASAP7_75t_L g773 ( 
.A(n_727),
.B(n_657),
.Y(n_773)
);

INVx1_ASAP7_75t_L g774 ( 
.A(n_684),
.Y(n_774)
);

NAND2xp5_ASAP7_75t_L g775 ( 
.A(n_702),
.B(n_654),
.Y(n_775)
);

INVx1_ASAP7_75t_L g776 ( 
.A(n_671),
.Y(n_776)
);

INVx3_ASAP7_75t_L g777 ( 
.A(n_734),
.Y(n_777)
);

AND2x4_ASAP7_75t_L g778 ( 
.A(n_750),
.B(n_584),
.Y(n_778)
);

AND2x6_ASAP7_75t_L g779 ( 
.A(n_751),
.B(n_525),
.Y(n_779)
);

INVx2_ASAP7_75t_SL g780 ( 
.A(n_682),
.Y(n_780)
);

INVx5_ASAP7_75t_L g781 ( 
.A(n_663),
.Y(n_781)
);

NAND2xp5_ASAP7_75t_L g782 ( 
.A(n_741),
.B(n_658),
.Y(n_782)
);

BUFx6f_ASAP7_75t_L g783 ( 
.A(n_734),
.Y(n_783)
);

INVx2_ASAP7_75t_L g784 ( 
.A(n_703),
.Y(n_784)
);

NAND2xp5_ASAP7_75t_SL g785 ( 
.A(n_692),
.B(n_627),
.Y(n_785)
);

INVx4_ASAP7_75t_L g786 ( 
.A(n_748),
.Y(n_786)
);

INVx2_ASAP7_75t_L g787 ( 
.A(n_705),
.Y(n_787)
);

BUFx2_ASAP7_75t_L g788 ( 
.A(n_714),
.Y(n_788)
);

INVx4_ASAP7_75t_L g789 ( 
.A(n_748),
.Y(n_789)
);

INVx1_ASAP7_75t_L g790 ( 
.A(n_686),
.Y(n_790)
);

INVx4_ASAP7_75t_SL g791 ( 
.A(n_663),
.Y(n_791)
);

AND2x2_ASAP7_75t_L g792 ( 
.A(n_711),
.B(n_575),
.Y(n_792)
);

INVx2_ASAP7_75t_L g793 ( 
.A(n_717),
.Y(n_793)
);

INVx2_ASAP7_75t_L g794 ( 
.A(n_718),
.Y(n_794)
);

NAND2xp5_ASAP7_75t_SL g795 ( 
.A(n_667),
.B(n_629),
.Y(n_795)
);

NAND2xp5_ASAP7_75t_L g796 ( 
.A(n_741),
.B(n_626),
.Y(n_796)
);

INVx4_ASAP7_75t_L g797 ( 
.A(n_722),
.Y(n_797)
);

INVx4_ASAP7_75t_L g798 ( 
.A(n_694),
.Y(n_798)
);

INVx3_ASAP7_75t_L g799 ( 
.A(n_694),
.Y(n_799)
);

NAND2xp5_ASAP7_75t_L g800 ( 
.A(n_741),
.B(n_735),
.Y(n_800)
);

INVx2_ASAP7_75t_L g801 ( 
.A(n_728),
.Y(n_801)
);

BUFx6f_ASAP7_75t_L g802 ( 
.A(n_694),
.Y(n_802)
);

BUFx3_ASAP7_75t_L g803 ( 
.A(n_752),
.Y(n_803)
);

AND2x2_ASAP7_75t_L g804 ( 
.A(n_710),
.B(n_548),
.Y(n_804)
);

INVx2_ASAP7_75t_L g805 ( 
.A(n_690),
.Y(n_805)
);

BUFx10_ASAP7_75t_L g806 ( 
.A(n_668),
.Y(n_806)
);

AND2x2_ASAP7_75t_L g807 ( 
.A(n_710),
.B(n_665),
.Y(n_807)
);

NAND3x1_ASAP7_75t_L g808 ( 
.A(n_695),
.B(n_623),
.C(n_648),
.Y(n_808)
);

INVx3_ASAP7_75t_L g809 ( 
.A(n_673),
.Y(n_809)
);

AND3x4_ASAP7_75t_L g810 ( 
.A(n_693),
.B(n_594),
.C(n_592),
.Y(n_810)
);

INVx1_ASAP7_75t_L g811 ( 
.A(n_688),
.Y(n_811)
);

AND2x2_ASAP7_75t_L g812 ( 
.A(n_732),
.B(n_659),
.Y(n_812)
);

BUFx6f_ASAP7_75t_L g813 ( 
.A(n_738),
.Y(n_813)
);

INVx2_ASAP7_75t_L g814 ( 
.A(n_691),
.Y(n_814)
);

INVx3_ASAP7_75t_L g815 ( 
.A(n_744),
.Y(n_815)
);

AOI22xp33_ASAP7_75t_L g816 ( 
.A1(n_741),
.A2(n_639),
.B1(n_652),
.B2(n_629),
.Y(n_816)
);

AND2x6_ASAP7_75t_L g817 ( 
.A(n_745),
.B(n_530),
.Y(n_817)
);

INVx1_ASAP7_75t_L g818 ( 
.A(n_689),
.Y(n_818)
);

INVx4_ASAP7_75t_L g819 ( 
.A(n_706),
.Y(n_819)
);

OR2x2_ASAP7_75t_SL g820 ( 
.A(n_724),
.B(n_405),
.Y(n_820)
);

INVx1_ASAP7_75t_L g821 ( 
.A(n_699),
.Y(n_821)
);

AND2x2_ASAP7_75t_SL g822 ( 
.A(n_731),
.B(n_623),
.Y(n_822)
);

INVx1_ASAP7_75t_L g823 ( 
.A(n_704),
.Y(n_823)
);

AND2x2_ASAP7_75t_SL g824 ( 
.A(n_731),
.B(n_410),
.Y(n_824)
);

AOI22xp5_ASAP7_75t_L g825 ( 
.A1(n_669),
.A2(n_655),
.B1(n_661),
.B2(n_650),
.Y(n_825)
);

NAND2xp5_ASAP7_75t_L g826 ( 
.A(n_708),
.B(n_513),
.Y(n_826)
);

INVx4_ASAP7_75t_L g827 ( 
.A(n_706),
.Y(n_827)
);

NOR2xp33_ASAP7_75t_L g828 ( 
.A(n_670),
.B(n_551),
.Y(n_828)
);

INVx2_ASAP7_75t_L g829 ( 
.A(n_709),
.Y(n_829)
);

NAND2xp5_ASAP7_75t_SL g830 ( 
.A(n_675),
.B(n_565),
.Y(n_830)
);

INVx2_ASAP7_75t_L g831 ( 
.A(n_713),
.Y(n_831)
);

INVx1_ASAP7_75t_L g832 ( 
.A(n_715),
.Y(n_832)
);

NOR2xp33_ASAP7_75t_L g833 ( 
.A(n_677),
.B(n_599),
.Y(n_833)
);

NAND2xp5_ASAP7_75t_L g834 ( 
.A(n_716),
.B(n_398),
.Y(n_834)
);

OR2x2_ASAP7_75t_L g835 ( 
.A(n_723),
.B(n_535),
.Y(n_835)
);

INVx2_ASAP7_75t_L g836 ( 
.A(n_726),
.Y(n_836)
);

NAND2xp5_ASAP7_75t_L g837 ( 
.A(n_807),
.B(n_678),
.Y(n_837)
);

INVx1_ASAP7_75t_L g838 ( 
.A(n_776),
.Y(n_838)
);

BUFx6f_ASAP7_75t_L g839 ( 
.A(n_762),
.Y(n_839)
);

AOI22xp5_ASAP7_75t_L g840 ( 
.A1(n_824),
.A2(n_698),
.B1(n_700),
.B2(n_696),
.Y(n_840)
);

NOR2xp33_ASAP7_75t_L g841 ( 
.A(n_753),
.B(n_707),
.Y(n_841)
);

CKINVDCx5p33_ASAP7_75t_R g842 ( 
.A(n_788),
.Y(n_842)
);

NAND2xp33_ASAP7_75t_L g843 ( 
.A(n_800),
.B(n_782),
.Y(n_843)
);

INVx2_ASAP7_75t_L g844 ( 
.A(n_754),
.Y(n_844)
);

AOI22xp33_ASAP7_75t_L g845 ( 
.A1(n_756),
.A2(n_439),
.B1(n_519),
.B2(n_465),
.Y(n_845)
);

NAND2xp5_ASAP7_75t_SL g846 ( 
.A(n_792),
.B(n_720),
.Y(n_846)
);

AND2x2_ASAP7_75t_L g847 ( 
.A(n_761),
.B(n_725),
.Y(n_847)
);

CKINVDCx11_ASAP7_75t_R g848 ( 
.A(n_806),
.Y(n_848)
);

NAND2xp5_ASAP7_75t_L g849 ( 
.A(n_819),
.B(n_739),
.Y(n_849)
);

NAND2xp5_ASAP7_75t_L g850 ( 
.A(n_819),
.B(n_827),
.Y(n_850)
);

INVx2_ASAP7_75t_L g851 ( 
.A(n_767),
.Y(n_851)
);

INVx3_ASAP7_75t_L g852 ( 
.A(n_827),
.Y(n_852)
);

INVx1_ASAP7_75t_L g853 ( 
.A(n_776),
.Y(n_853)
);

INVx1_ASAP7_75t_L g854 ( 
.A(n_755),
.Y(n_854)
);

NAND2x1p5_ASAP7_75t_L g855 ( 
.A(n_761),
.B(n_695),
.Y(n_855)
);

INVx1_ASAP7_75t_L g856 ( 
.A(n_774),
.Y(n_856)
);

BUFx3_ASAP7_75t_L g857 ( 
.A(n_758),
.Y(n_857)
);

INVx1_ASAP7_75t_L g858 ( 
.A(n_790),
.Y(n_858)
);

INVx1_ASAP7_75t_L g859 ( 
.A(n_811),
.Y(n_859)
);

NAND2xp5_ASAP7_75t_SL g860 ( 
.A(n_780),
.B(n_742),
.Y(n_860)
);

NAND2xp5_ASAP7_75t_L g861 ( 
.A(n_773),
.B(n_747),
.Y(n_861)
);

NAND2xp5_ASAP7_75t_L g862 ( 
.A(n_786),
.B(n_729),
.Y(n_862)
);

NAND2xp5_ASAP7_75t_L g863 ( 
.A(n_786),
.B(n_730),
.Y(n_863)
);

AOI22xp5_ASAP7_75t_L g864 ( 
.A1(n_808),
.A2(n_605),
.B1(n_617),
.B2(n_603),
.Y(n_864)
);

NAND2xp5_ASAP7_75t_L g865 ( 
.A(n_789),
.B(n_775),
.Y(n_865)
);

NAND2xp5_ASAP7_75t_L g866 ( 
.A(n_789),
.B(n_540),
.Y(n_866)
);

AND2x6_ASAP7_75t_SL g867 ( 
.A(n_828),
.B(n_471),
.Y(n_867)
);

INVx1_ASAP7_75t_L g868 ( 
.A(n_818),
.Y(n_868)
);

NAND2xp5_ASAP7_75t_SL g869 ( 
.A(n_822),
.B(n_736),
.Y(n_869)
);

NAND2xp5_ASAP7_75t_L g870 ( 
.A(n_796),
.B(n_399),
.Y(n_870)
);

O2A1O1Ixp5_ASAP7_75t_L g871 ( 
.A1(n_821),
.A2(n_823),
.B(n_832),
.C(n_778),
.Y(n_871)
);

AOI22xp33_ASAP7_75t_L g872 ( 
.A1(n_757),
.A2(n_342),
.B1(n_681),
.B2(n_663),
.Y(n_872)
);

INVx2_ASAP7_75t_SL g873 ( 
.A(n_758),
.Y(n_873)
);

NOR2xp33_ASAP7_75t_L g874 ( 
.A(n_763),
.B(n_619),
.Y(n_874)
);

NAND2xp5_ASAP7_75t_L g875 ( 
.A(n_797),
.B(n_400),
.Y(n_875)
);

NOR2x1p5_ASAP7_75t_L g876 ( 
.A(n_764),
.B(n_401),
.Y(n_876)
);

AOI22xp5_ASAP7_75t_L g877 ( 
.A1(n_757),
.A2(n_544),
.B1(n_473),
.B2(n_620),
.Y(n_877)
);

NOR2xp33_ASAP7_75t_L g878 ( 
.A(n_770),
.B(n_719),
.Y(n_878)
);

NAND2xp5_ASAP7_75t_L g879 ( 
.A(n_797),
.B(n_402),
.Y(n_879)
);

NAND2xp5_ASAP7_75t_L g880 ( 
.A(n_804),
.B(n_407),
.Y(n_880)
);

NAND3xp33_ASAP7_75t_SL g881 ( 
.A(n_825),
.B(n_737),
.C(n_733),
.Y(n_881)
);

NAND2xp5_ASAP7_75t_L g882 ( 
.A(n_778),
.B(n_408),
.Y(n_882)
);

NOR2xp33_ASAP7_75t_L g883 ( 
.A(n_765),
.B(n_411),
.Y(n_883)
);

BUFx3_ASAP7_75t_L g884 ( 
.A(n_803),
.Y(n_884)
);

O2A1O1Ixp5_ASAP7_75t_L g885 ( 
.A1(n_834),
.A2(n_538),
.B(n_663),
.C(n_681),
.Y(n_885)
);

NAND2xp5_ASAP7_75t_L g886 ( 
.A(n_812),
.B(n_412),
.Y(n_886)
);

INVx3_ASAP7_75t_L g887 ( 
.A(n_784),
.Y(n_887)
);

NAND2xp5_ASAP7_75t_L g888 ( 
.A(n_829),
.B(n_415),
.Y(n_888)
);

AOI22xp33_ASAP7_75t_L g889 ( 
.A1(n_757),
.A2(n_681),
.B1(n_418),
.B2(n_419),
.Y(n_889)
);

INVx2_ASAP7_75t_L g890 ( 
.A(n_787),
.Y(n_890)
);

NAND2xp5_ASAP7_75t_L g891 ( 
.A(n_831),
.B(n_417),
.Y(n_891)
);

AOI22xp5_ASAP7_75t_L g892 ( 
.A1(n_816),
.A2(n_422),
.B1(n_423),
.B2(n_420),
.Y(n_892)
);

AND2x4_ASAP7_75t_L g893 ( 
.A(n_836),
.B(n_424),
.Y(n_893)
);

INVx3_ASAP7_75t_L g894 ( 
.A(n_793),
.Y(n_894)
);

NAND2xp5_ASAP7_75t_SL g895 ( 
.A(n_762),
.B(n_427),
.Y(n_895)
);

NAND2xp5_ASAP7_75t_L g896 ( 
.A(n_798),
.B(n_428),
.Y(n_896)
);

INVx1_ASAP7_75t_L g897 ( 
.A(n_794),
.Y(n_897)
);

NAND2xp5_ASAP7_75t_L g898 ( 
.A(n_798),
.B(n_801),
.Y(n_898)
);

OR2x6_ASAP7_75t_L g899 ( 
.A(n_788),
.B(n_8),
.Y(n_899)
);

AOI22xp33_ASAP7_75t_L g900 ( 
.A1(n_779),
.A2(n_681),
.B1(n_541),
.B2(n_533),
.Y(n_900)
);

NAND2xp5_ASAP7_75t_L g901 ( 
.A(n_805),
.B(n_814),
.Y(n_901)
);

AND2x6_ASAP7_75t_SL g902 ( 
.A(n_833),
.B(n_9),
.Y(n_902)
);

NAND2xp5_ASAP7_75t_L g903 ( 
.A(n_771),
.B(n_772),
.Y(n_903)
);

INVx1_ASAP7_75t_L g904 ( 
.A(n_809),
.Y(n_904)
);

XNOR2xp5_ASAP7_75t_L g905 ( 
.A(n_810),
.B(n_429),
.Y(n_905)
);

INVx1_ASAP7_75t_L g906 ( 
.A(n_768),
.Y(n_906)
);

AND2x2_ASAP7_75t_L g907 ( 
.A(n_765),
.B(n_431),
.Y(n_907)
);

INVx2_ASAP7_75t_L g908 ( 
.A(n_815),
.Y(n_908)
);

INVx1_ASAP7_75t_L g909 ( 
.A(n_835),
.Y(n_909)
);

O2A1O1Ixp33_ASAP7_75t_L g910 ( 
.A1(n_826),
.A2(n_532),
.B(n_531),
.C(n_529),
.Y(n_910)
);

NAND2xp5_ASAP7_75t_L g911 ( 
.A(n_762),
.B(n_432),
.Y(n_911)
);

INVx2_ASAP7_75t_L g912 ( 
.A(n_813),
.Y(n_912)
);

NAND2xp5_ASAP7_75t_SL g913 ( 
.A(n_783),
.B(n_434),
.Y(n_913)
);

NAND2xp33_ASAP7_75t_L g914 ( 
.A(n_779),
.B(n_528),
.Y(n_914)
);

NOR2xp33_ASAP7_75t_L g915 ( 
.A(n_830),
.B(n_435),
.Y(n_915)
);

NAND2xp5_ASAP7_75t_L g916 ( 
.A(n_783),
.B(n_438),
.Y(n_916)
);

INVx1_ASAP7_75t_L g917 ( 
.A(n_813),
.Y(n_917)
);

INVx2_ASAP7_75t_SL g918 ( 
.A(n_760),
.Y(n_918)
);

INVx4_ASAP7_75t_L g919 ( 
.A(n_839),
.Y(n_919)
);

AND2x2_ASAP7_75t_L g920 ( 
.A(n_873),
.B(n_759),
.Y(n_920)
);

NAND2xp5_ASAP7_75t_L g921 ( 
.A(n_841),
.B(n_783),
.Y(n_921)
);

HB1xp67_ASAP7_75t_L g922 ( 
.A(n_857),
.Y(n_922)
);

INVx3_ASAP7_75t_L g923 ( 
.A(n_839),
.Y(n_923)
);

AOI22xp33_ASAP7_75t_SL g924 ( 
.A1(n_861),
.A2(n_806),
.B1(n_769),
.B2(n_766),
.Y(n_924)
);

BUFx8_ASAP7_75t_L g925 ( 
.A(n_847),
.Y(n_925)
);

NAND2xp5_ASAP7_75t_SL g926 ( 
.A(n_837),
.B(n_802),
.Y(n_926)
);

NOR2xp33_ASAP7_75t_R g927 ( 
.A(n_842),
.B(n_777),
.Y(n_927)
);

BUFx3_ASAP7_75t_L g928 ( 
.A(n_884),
.Y(n_928)
);

INVx1_ASAP7_75t_L g929 ( 
.A(n_838),
.Y(n_929)
);

INVx1_ASAP7_75t_L g930 ( 
.A(n_853),
.Y(n_930)
);

BUFx6f_ASAP7_75t_L g931 ( 
.A(n_839),
.Y(n_931)
);

NAND3xp33_ASAP7_75t_SL g932 ( 
.A(n_877),
.B(n_795),
.C(n_785),
.Y(n_932)
);

INVx2_ASAP7_75t_L g933 ( 
.A(n_844),
.Y(n_933)
);

BUFx6f_ASAP7_75t_L g934 ( 
.A(n_855),
.Y(n_934)
);

BUFx2_ASAP7_75t_L g935 ( 
.A(n_918),
.Y(n_935)
);

NOR2xp33_ASAP7_75t_L g936 ( 
.A(n_846),
.B(n_820),
.Y(n_936)
);

INVx1_ASAP7_75t_L g937 ( 
.A(n_854),
.Y(n_937)
);

CKINVDCx5p33_ASAP7_75t_R g938 ( 
.A(n_848),
.Y(n_938)
);

BUFx3_ASAP7_75t_L g939 ( 
.A(n_904),
.Y(n_939)
);

INVx2_ASAP7_75t_L g940 ( 
.A(n_851),
.Y(n_940)
);

BUFx6f_ASAP7_75t_L g941 ( 
.A(n_912),
.Y(n_941)
);

BUFx6f_ASAP7_75t_L g942 ( 
.A(n_898),
.Y(n_942)
);

CKINVDCx5p33_ASAP7_75t_R g943 ( 
.A(n_840),
.Y(n_943)
);

INVx1_ASAP7_75t_SL g944 ( 
.A(n_907),
.Y(n_944)
);

NAND2xp5_ASAP7_75t_SL g945 ( 
.A(n_849),
.B(n_852),
.Y(n_945)
);

INVx2_ASAP7_75t_L g946 ( 
.A(n_890),
.Y(n_946)
);

INVx1_ASAP7_75t_L g947 ( 
.A(n_856),
.Y(n_947)
);

NAND2xp5_ASAP7_75t_SL g948 ( 
.A(n_852),
.B(n_802),
.Y(n_948)
);

INVx2_ASAP7_75t_L g949 ( 
.A(n_858),
.Y(n_949)
);

INVx3_ASAP7_75t_L g950 ( 
.A(n_887),
.Y(n_950)
);

NAND2xp5_ASAP7_75t_L g951 ( 
.A(n_865),
.B(n_802),
.Y(n_951)
);

INVx3_ASAP7_75t_L g952 ( 
.A(n_887),
.Y(n_952)
);

INVx2_ASAP7_75t_L g953 ( 
.A(n_859),
.Y(n_953)
);

NAND2xp5_ASAP7_75t_L g954 ( 
.A(n_862),
.B(n_779),
.Y(n_954)
);

NOR2x1p5_ASAP7_75t_L g955 ( 
.A(n_881),
.B(n_799),
.Y(n_955)
);

INVx1_ASAP7_75t_L g956 ( 
.A(n_868),
.Y(n_956)
);

INVx3_ASAP7_75t_L g957 ( 
.A(n_894),
.Y(n_957)
);

NAND3xp33_ASAP7_75t_SL g958 ( 
.A(n_877),
.B(n_442),
.C(n_440),
.Y(n_958)
);

INVx1_ASAP7_75t_L g959 ( 
.A(n_901),
.Y(n_959)
);

INVx1_ASAP7_75t_L g960 ( 
.A(n_897),
.Y(n_960)
);

BUFx6f_ASAP7_75t_L g961 ( 
.A(n_893),
.Y(n_961)
);

INVx6_ASAP7_75t_L g962 ( 
.A(n_899),
.Y(n_962)
);

NAND2xp5_ASAP7_75t_L g963 ( 
.A(n_863),
.B(n_813),
.Y(n_963)
);

CKINVDCx5p33_ASAP7_75t_R g964 ( 
.A(n_878),
.Y(n_964)
);

NOR3xp33_ASAP7_75t_SL g965 ( 
.A(n_869),
.B(n_449),
.C(n_448),
.Y(n_965)
);

HB1xp67_ASAP7_75t_L g966 ( 
.A(n_909),
.Y(n_966)
);

INVx2_ASAP7_75t_L g967 ( 
.A(n_894),
.Y(n_967)
);

INVx1_ASAP7_75t_L g968 ( 
.A(n_906),
.Y(n_968)
);

NOR3xp33_ASAP7_75t_SL g969 ( 
.A(n_874),
.B(n_451),
.C(n_450),
.Y(n_969)
);

INVx1_ASAP7_75t_L g970 ( 
.A(n_903),
.Y(n_970)
);

NAND2xp5_ASAP7_75t_L g971 ( 
.A(n_880),
.B(n_817),
.Y(n_971)
);

BUFx6f_ASAP7_75t_L g972 ( 
.A(n_893),
.Y(n_972)
);

INVx2_ASAP7_75t_L g973 ( 
.A(n_908),
.Y(n_973)
);

INVx1_ASAP7_75t_L g974 ( 
.A(n_917),
.Y(n_974)
);

INVx5_ASAP7_75t_L g975 ( 
.A(n_899),
.Y(n_975)
);

INVx3_ASAP7_75t_L g976 ( 
.A(n_850),
.Y(n_976)
);

INVx1_ASAP7_75t_L g977 ( 
.A(n_871),
.Y(n_977)
);

INVx2_ASAP7_75t_L g978 ( 
.A(n_866),
.Y(n_978)
);

OAI21xp5_ASAP7_75t_L g979 ( 
.A1(n_977),
.A2(n_843),
.B(n_870),
.Y(n_979)
);

BUFx4f_ASAP7_75t_L g980 ( 
.A(n_961),
.Y(n_980)
);

OAI21xp5_ASAP7_75t_L g981 ( 
.A1(n_970),
.A2(n_885),
.B(n_886),
.Y(n_981)
);

OAI21x1_ASAP7_75t_L g982 ( 
.A1(n_976),
.A2(n_916),
.B(n_911),
.Y(n_982)
);

AND2x4_ASAP7_75t_L g983 ( 
.A(n_934),
.B(n_876),
.Y(n_983)
);

OAI21xp5_ASAP7_75t_L g984 ( 
.A1(n_959),
.A2(n_889),
.B(n_892),
.Y(n_984)
);

NOR2xp33_ASAP7_75t_L g985 ( 
.A(n_964),
.B(n_883),
.Y(n_985)
);

NAND2xp5_ASAP7_75t_L g986 ( 
.A(n_978),
.B(n_915),
.Y(n_986)
);

INVx1_ASAP7_75t_L g987 ( 
.A(n_929),
.Y(n_987)
);

AO31x2_ASAP7_75t_L g988 ( 
.A1(n_951),
.A2(n_891),
.A3(n_888),
.B(n_875),
.Y(n_988)
);

INVx2_ASAP7_75t_L g989 ( 
.A(n_949),
.Y(n_989)
);

AOI21x1_ASAP7_75t_L g990 ( 
.A1(n_945),
.A2(n_896),
.B(n_879),
.Y(n_990)
);

AOI21x1_ASAP7_75t_L g991 ( 
.A1(n_971),
.A2(n_913),
.B(n_895),
.Y(n_991)
);

AOI21x1_ASAP7_75t_L g992 ( 
.A1(n_954),
.A2(n_882),
.B(n_860),
.Y(n_992)
);

AND2x4_ASAP7_75t_L g993 ( 
.A(n_934),
.B(n_961),
.Y(n_993)
);

OAI21x1_ASAP7_75t_L g994 ( 
.A1(n_976),
.A2(n_910),
.B(n_872),
.Y(n_994)
);

NAND2xp5_ASAP7_75t_L g995 ( 
.A(n_930),
.B(n_845),
.Y(n_995)
);

AO31x2_ASAP7_75t_L g996 ( 
.A1(n_963),
.A2(n_914),
.A3(n_900),
.B(n_817),
.Y(n_996)
);

AO31x2_ASAP7_75t_L g997 ( 
.A1(n_921),
.A2(n_817),
.A3(n_791),
.B(n_12),
.Y(n_997)
);

AND2x2_ASAP7_75t_L g998 ( 
.A(n_920),
.B(n_864),
.Y(n_998)
);

NAND2xp5_ASAP7_75t_L g999 ( 
.A(n_937),
.B(n_905),
.Y(n_999)
);

OAI21xp5_ASAP7_75t_L g1000 ( 
.A1(n_947),
.A2(n_781),
.B(n_455),
.Y(n_1000)
);

AOI31xp67_ASAP7_75t_L g1001 ( 
.A1(n_926),
.A2(n_791),
.A3(n_494),
.B(n_512),
.Y(n_1001)
);

OAI21x1_ASAP7_75t_L g1002 ( 
.A1(n_948),
.A2(n_29),
.B(n_23),
.Y(n_1002)
);

AOI21x1_ASAP7_75t_L g1003 ( 
.A1(n_974),
.A2(n_781),
.B(n_460),
.Y(n_1003)
);

NAND2xp5_ASAP7_75t_L g1004 ( 
.A(n_956),
.B(n_452),
.Y(n_1004)
);

AOI21xp5_ASAP7_75t_L g1005 ( 
.A1(n_942),
.A2(n_781),
.B(n_463),
.Y(n_1005)
);

OAI21x1_ASAP7_75t_L g1006 ( 
.A1(n_950),
.A2(n_35),
.B(n_33),
.Y(n_1006)
);

CKINVDCx5p33_ASAP7_75t_R g1007 ( 
.A(n_938),
.Y(n_1007)
);

AOI21xp33_ASAP7_75t_L g1008 ( 
.A1(n_944),
.A2(n_467),
.B(n_462),
.Y(n_1008)
);

OAI22xp5_ASAP7_75t_L g1009 ( 
.A1(n_943),
.A2(n_504),
.B1(n_474),
.B2(n_524),
.Y(n_1009)
);

BUFx2_ASAP7_75t_L g1010 ( 
.A(n_922),
.Y(n_1010)
);

BUFx2_ASAP7_75t_L g1011 ( 
.A(n_935),
.Y(n_1011)
);

OAI21x1_ASAP7_75t_L g1012 ( 
.A1(n_950),
.A2(n_37),
.B(n_36),
.Y(n_1012)
);

NAND2xp33_ASAP7_75t_L g1013 ( 
.A(n_934),
.B(n_470),
.Y(n_1013)
);

OAI21xp5_ASAP7_75t_L g1014 ( 
.A1(n_953),
.A2(n_477),
.B(n_476),
.Y(n_1014)
);

CKINVDCx5p33_ASAP7_75t_R g1015 ( 
.A(n_925),
.Y(n_1015)
);

INVx3_ASAP7_75t_L g1016 ( 
.A(n_928),
.Y(n_1016)
);

OAI21x1_ASAP7_75t_L g1017 ( 
.A1(n_952),
.A2(n_46),
.B(n_42),
.Y(n_1017)
);

OAI21x1_ASAP7_75t_L g1018 ( 
.A1(n_952),
.A2(n_48),
.B(n_47),
.Y(n_1018)
);

OAI21x1_ASAP7_75t_L g1019 ( 
.A1(n_957),
.A2(n_53),
.B(n_50),
.Y(n_1019)
);

NOR2xp33_ASAP7_75t_L g1020 ( 
.A(n_932),
.B(n_936),
.Y(n_1020)
);

INVx1_ASAP7_75t_L g1021 ( 
.A(n_960),
.Y(n_1021)
);

NAND3xp33_ASAP7_75t_L g1022 ( 
.A(n_924),
.B(n_482),
.C(n_481),
.Y(n_1022)
);

NAND2xp5_ASAP7_75t_L g1023 ( 
.A(n_942),
.B(n_957),
.Y(n_1023)
);

NAND2xp5_ASAP7_75t_L g1024 ( 
.A(n_942),
.B(n_484),
.Y(n_1024)
);

INVxp67_ASAP7_75t_L g1025 ( 
.A(n_1011),
.Y(n_1025)
);

BUFx4f_ASAP7_75t_L g1026 ( 
.A(n_983),
.Y(n_1026)
);

INVx1_ASAP7_75t_SL g1027 ( 
.A(n_1010),
.Y(n_1027)
);

INVx1_ASAP7_75t_SL g1028 ( 
.A(n_1016),
.Y(n_1028)
);

OAI21x1_ASAP7_75t_L g1029 ( 
.A1(n_982),
.A2(n_968),
.B(n_923),
.Y(n_1029)
);

INVx2_ASAP7_75t_L g1030 ( 
.A(n_987),
.Y(n_1030)
);

OAI21x1_ASAP7_75t_L g1031 ( 
.A1(n_990),
.A2(n_979),
.B(n_981),
.Y(n_1031)
);

OAI21x1_ASAP7_75t_SL g1032 ( 
.A1(n_992),
.A2(n_919),
.B(n_967),
.Y(n_1032)
);

NAND4xp25_ASAP7_75t_L g1033 ( 
.A(n_999),
.B(n_985),
.C(n_1020),
.D(n_998),
.Y(n_1033)
);

AO31x2_ASAP7_75t_L g1034 ( 
.A1(n_986),
.A2(n_946),
.A3(n_933),
.B(n_940),
.Y(n_1034)
);

INVx2_ASAP7_75t_L g1035 ( 
.A(n_1021),
.Y(n_1035)
);

AND2x2_ASAP7_75t_L g1036 ( 
.A(n_989),
.B(n_966),
.Y(n_1036)
);

INVx2_ASAP7_75t_L g1037 ( 
.A(n_1023),
.Y(n_1037)
);

NOR2xp33_ASAP7_75t_SL g1038 ( 
.A(n_1007),
.B(n_925),
.Y(n_1038)
);

OAI21xp5_ASAP7_75t_L g1039 ( 
.A1(n_984),
.A2(n_958),
.B(n_965),
.Y(n_1039)
);

OAI21x1_ASAP7_75t_L g1040 ( 
.A1(n_1002),
.A2(n_923),
.B(n_973),
.Y(n_1040)
);

CKINVDCx11_ASAP7_75t_R g1041 ( 
.A(n_983),
.Y(n_1041)
);

HB1xp67_ASAP7_75t_L g1042 ( 
.A(n_980),
.Y(n_1042)
);

BUFx4f_ASAP7_75t_SL g1043 ( 
.A(n_993),
.Y(n_1043)
);

AO31x2_ASAP7_75t_L g1044 ( 
.A1(n_995),
.A2(n_919),
.A3(n_969),
.B(n_955),
.Y(n_1044)
);

OAI21xp5_ASAP7_75t_L g1045 ( 
.A1(n_1000),
.A2(n_939),
.B(n_486),
.Y(n_1045)
);

OAI21x1_ASAP7_75t_L g1046 ( 
.A1(n_1006),
.A2(n_941),
.B(n_931),
.Y(n_1046)
);

BUFx3_ASAP7_75t_L g1047 ( 
.A(n_993),
.Y(n_1047)
);

OAI21x1_ASAP7_75t_L g1048 ( 
.A1(n_1012),
.A2(n_941),
.B(n_931),
.Y(n_1048)
);

INVx2_ASAP7_75t_L g1049 ( 
.A(n_997),
.Y(n_1049)
);

O2A1O1Ixp33_ASAP7_75t_SL g1050 ( 
.A1(n_1024),
.A2(n_867),
.B(n_972),
.C(n_961),
.Y(n_1050)
);

OA21x2_ASAP7_75t_L g1051 ( 
.A1(n_994),
.A2(n_489),
.B(n_485),
.Y(n_1051)
);

INVx1_ASAP7_75t_L g1052 ( 
.A(n_1017),
.Y(n_1052)
);

NAND2xp5_ASAP7_75t_L g1053 ( 
.A(n_1004),
.B(n_972),
.Y(n_1053)
);

INVx1_ASAP7_75t_L g1054 ( 
.A(n_1018),
.Y(n_1054)
);

INVx4_ASAP7_75t_SL g1055 ( 
.A(n_997),
.Y(n_1055)
);

OAI22xp33_ASAP7_75t_L g1056 ( 
.A1(n_1022),
.A2(n_975),
.B1(n_972),
.B2(n_962),
.Y(n_1056)
);

OA21x2_ASAP7_75t_L g1057 ( 
.A1(n_1019),
.A2(n_491),
.B(n_490),
.Y(n_1057)
);

AND2x4_ASAP7_75t_L g1058 ( 
.A(n_991),
.B(n_975),
.Y(n_1058)
);

AND2x4_ASAP7_75t_L g1059 ( 
.A(n_1005),
.B(n_975),
.Y(n_1059)
);

OA21x2_ASAP7_75t_L g1060 ( 
.A1(n_1003),
.A2(n_495),
.B(n_492),
.Y(n_1060)
);

OAI21x1_ASAP7_75t_L g1061 ( 
.A1(n_1014),
.A2(n_941),
.B(n_931),
.Y(n_1061)
);

INVx1_ASAP7_75t_L g1062 ( 
.A(n_997),
.Y(n_1062)
);

INVx2_ASAP7_75t_L g1063 ( 
.A(n_988),
.Y(n_1063)
);

NOR2x1_ASAP7_75t_R g1064 ( 
.A(n_1015),
.B(n_962),
.Y(n_1064)
);

AO32x2_ASAP7_75t_L g1065 ( 
.A1(n_1055),
.A2(n_1009),
.A3(n_1001),
.B1(n_988),
.B2(n_996),
.Y(n_1065)
);

AOI22xp33_ASAP7_75t_L g1066 ( 
.A1(n_1033),
.A2(n_1008),
.B1(n_1013),
.B2(n_927),
.Y(n_1066)
);

AND2x4_ASAP7_75t_L g1067 ( 
.A(n_1047),
.B(n_996),
.Y(n_1067)
);

AND2x6_ASAP7_75t_L g1068 ( 
.A(n_1059),
.B(n_996),
.Y(n_1068)
);

AND2x2_ASAP7_75t_L g1069 ( 
.A(n_1036),
.B(n_500),
.Y(n_1069)
);

BUFx2_ASAP7_75t_L g1070 ( 
.A(n_1034),
.Y(n_1070)
);

BUFx2_ASAP7_75t_L g1071 ( 
.A(n_1034),
.Y(n_1071)
);

INVx1_ASAP7_75t_SL g1072 ( 
.A(n_1027),
.Y(n_1072)
);

CKINVDCx6p67_ASAP7_75t_R g1073 ( 
.A(n_1041),
.Y(n_1073)
);

A2O1A1Ixp33_ASAP7_75t_L g1074 ( 
.A1(n_1039),
.A2(n_516),
.B(n_506),
.C(n_522),
.Y(n_1074)
);

OR2x6_ASAP7_75t_L g1075 ( 
.A(n_1042),
.B(n_902),
.Y(n_1075)
);

INVxp67_ASAP7_75t_L g1076 ( 
.A(n_1028),
.Y(n_1076)
);

OAI22xp33_ASAP7_75t_L g1077 ( 
.A1(n_1033),
.A2(n_515),
.B1(n_521),
.B2(n_520),
.Y(n_1077)
);

INVx1_ASAP7_75t_SL g1078 ( 
.A(n_1043),
.Y(n_1078)
);

NAND2xp33_ASAP7_75t_SL g1079 ( 
.A(n_1053),
.B(n_505),
.Y(n_1079)
);

AOI22xp33_ASAP7_75t_L g1080 ( 
.A1(n_1045),
.A2(n_518),
.B1(n_517),
.B2(n_514),
.Y(n_1080)
);

INVx1_ASAP7_75t_L g1081 ( 
.A(n_1030),
.Y(n_1081)
);

INVx2_ASAP7_75t_L g1082 ( 
.A(n_1035),
.Y(n_1082)
);

AOI22xp33_ASAP7_75t_L g1083 ( 
.A1(n_1058),
.A2(n_509),
.B1(n_507),
.B2(n_988),
.Y(n_1083)
);

INVx1_ASAP7_75t_L g1084 ( 
.A(n_1037),
.Y(n_1084)
);

INVx1_ASAP7_75t_L g1085 ( 
.A(n_1034),
.Y(n_1085)
);

AO21x2_ASAP7_75t_L g1086 ( 
.A1(n_1052),
.A2(n_176),
.B(n_323),
.Y(n_1086)
);

INVx1_ASAP7_75t_L g1087 ( 
.A(n_1062),
.Y(n_1087)
);

INVx1_ASAP7_75t_L g1088 ( 
.A(n_1062),
.Y(n_1088)
);

BUFx8_ASAP7_75t_L g1089 ( 
.A(n_1059),
.Y(n_1089)
);

BUFx3_ASAP7_75t_L g1090 ( 
.A(n_1026),
.Y(n_1090)
);

A2O1A1Ixp33_ASAP7_75t_L g1091 ( 
.A1(n_1058),
.A2(n_9),
.B(n_10),
.C(n_12),
.Y(n_1091)
);

OAI21x1_ASAP7_75t_L g1092 ( 
.A1(n_1046),
.A2(n_181),
.B(n_318),
.Y(n_1092)
);

NAND2xp33_ASAP7_75t_L g1093 ( 
.A(n_1052),
.B(n_13),
.Y(n_1093)
);

AND2x2_ASAP7_75t_SL g1094 ( 
.A(n_1038),
.B(n_13),
.Y(n_1094)
);

INVx2_ASAP7_75t_L g1095 ( 
.A(n_1029),
.Y(n_1095)
);

INVx3_ASAP7_75t_L g1096 ( 
.A(n_1026),
.Y(n_1096)
);

OR2x2_ASAP7_75t_L g1097 ( 
.A(n_1025),
.B(n_14),
.Y(n_1097)
);

NAND2xp5_ASAP7_75t_L g1098 ( 
.A(n_1056),
.B(n_14),
.Y(n_1098)
);

AND2x4_ASAP7_75t_L g1099 ( 
.A(n_1044),
.B(n_54),
.Y(n_1099)
);

INVx1_ASAP7_75t_L g1100 ( 
.A(n_1032),
.Y(n_1100)
);

AND2x4_ASAP7_75t_L g1101 ( 
.A(n_1044),
.B(n_56),
.Y(n_1101)
);

OAI22xp5_ASAP7_75t_L g1102 ( 
.A1(n_1063),
.A2(n_1054),
.B1(n_1049),
.B2(n_1051),
.Y(n_1102)
);

AND2x4_ASAP7_75t_L g1103 ( 
.A(n_1044),
.B(n_60),
.Y(n_1103)
);

OAI211xp5_ASAP7_75t_L g1104 ( 
.A1(n_1091),
.A2(n_1050),
.B(n_1060),
.C(n_1051),
.Y(n_1104)
);

OA21x2_ASAP7_75t_L g1105 ( 
.A1(n_1085),
.A2(n_1031),
.B(n_1054),
.Y(n_1105)
);

OAI211xp5_ASAP7_75t_SL g1106 ( 
.A1(n_1066),
.A2(n_1064),
.B(n_1055),
.C(n_1060),
.Y(n_1106)
);

INVx5_ASAP7_75t_L g1107 ( 
.A(n_1103),
.Y(n_1107)
);

AOI22xp33_ASAP7_75t_L g1108 ( 
.A1(n_1093),
.A2(n_1061),
.B1(n_1057),
.B2(n_1040),
.Y(n_1108)
);

OAI22xp5_ASAP7_75t_L g1109 ( 
.A1(n_1098),
.A2(n_1057),
.B1(n_1064),
.B2(n_1048),
.Y(n_1109)
);

AOI22xp33_ASAP7_75t_L g1110 ( 
.A1(n_1094),
.A2(n_15),
.B1(n_17),
.B2(n_18),
.Y(n_1110)
);

AOI221xp5_ASAP7_75t_L g1111 ( 
.A1(n_1077),
.A2(n_1080),
.B1(n_1074),
.B2(n_1083),
.C(n_1069),
.Y(n_1111)
);

AOI221xp5_ASAP7_75t_L g1112 ( 
.A1(n_1076),
.A2(n_17),
.B1(n_19),
.B2(n_20),
.C(n_21),
.Y(n_1112)
);

AND2x2_ASAP7_75t_L g1113 ( 
.A(n_1084),
.B(n_62),
.Y(n_1113)
);

OAI22xp33_ASAP7_75t_L g1114 ( 
.A1(n_1075),
.A2(n_20),
.B1(n_21),
.B2(n_22),
.Y(n_1114)
);

AOI22xp33_ASAP7_75t_L g1115 ( 
.A1(n_1103),
.A2(n_65),
.B1(n_66),
.B2(n_69),
.Y(n_1115)
);

AOI221xp5_ASAP7_75t_L g1116 ( 
.A1(n_1072),
.A2(n_70),
.B1(n_74),
.B2(n_75),
.C(n_77),
.Y(n_1116)
);

AOI211xp5_ASAP7_75t_L g1117 ( 
.A1(n_1079),
.A2(n_79),
.B(n_80),
.C(n_81),
.Y(n_1117)
);

OAI221xp5_ASAP7_75t_L g1118 ( 
.A1(n_1075),
.A2(n_83),
.B1(n_89),
.B2(n_92),
.C(n_93),
.Y(n_1118)
);

OR2x2_ASAP7_75t_L g1119 ( 
.A(n_1081),
.B(n_94),
.Y(n_1119)
);

AOI22xp33_ASAP7_75t_L g1120 ( 
.A1(n_1099),
.A2(n_96),
.B1(n_97),
.B2(n_98),
.Y(n_1120)
);

OAI22xp33_ASAP7_75t_L g1121 ( 
.A1(n_1073),
.A2(n_100),
.B1(n_107),
.B2(n_108),
.Y(n_1121)
);

OAI21xp5_ASAP7_75t_SL g1122 ( 
.A1(n_1101),
.A2(n_114),
.B(n_116),
.Y(n_1122)
);

OAI21x1_ASAP7_75t_L g1123 ( 
.A1(n_1092),
.A2(n_117),
.B(n_124),
.Y(n_1123)
);

OAI22xp5_ASAP7_75t_L g1124 ( 
.A1(n_1090),
.A2(n_125),
.B1(n_126),
.B2(n_127),
.Y(n_1124)
);

INVx1_ASAP7_75t_L g1125 ( 
.A(n_1087),
.Y(n_1125)
);

OA21x2_ASAP7_75t_L g1126 ( 
.A1(n_1070),
.A2(n_130),
.B(n_131),
.Y(n_1126)
);

OAI22xp5_ASAP7_75t_L g1127 ( 
.A1(n_1096),
.A2(n_136),
.B1(n_137),
.B2(n_139),
.Y(n_1127)
);

AOI22xp33_ASAP7_75t_L g1128 ( 
.A1(n_1067),
.A2(n_140),
.B1(n_142),
.B2(n_149),
.Y(n_1128)
);

INVx2_ASAP7_75t_L g1129 ( 
.A(n_1082),
.Y(n_1129)
);

AOI22xp33_ASAP7_75t_L g1130 ( 
.A1(n_1067),
.A2(n_150),
.B1(n_153),
.B2(n_158),
.Y(n_1130)
);

INVx5_ASAP7_75t_L g1131 ( 
.A(n_1068),
.Y(n_1131)
);

BUFx3_ASAP7_75t_L g1132 ( 
.A(n_1089),
.Y(n_1132)
);

AOI221xp5_ASAP7_75t_L g1133 ( 
.A1(n_1097),
.A2(n_161),
.B1(n_162),
.B2(n_163),
.C(n_164),
.Y(n_1133)
);

AOI22xp33_ASAP7_75t_L g1134 ( 
.A1(n_1068),
.A2(n_169),
.B1(n_172),
.B2(n_180),
.Y(n_1134)
);

BUFx4f_ASAP7_75t_SL g1135 ( 
.A(n_1078),
.Y(n_1135)
);

INVx2_ASAP7_75t_L g1136 ( 
.A(n_1088),
.Y(n_1136)
);

OAI22xp5_ASAP7_75t_L g1137 ( 
.A1(n_1100),
.A2(n_1071),
.B1(n_1070),
.B2(n_1102),
.Y(n_1137)
);

AO21x2_ASAP7_75t_L g1138 ( 
.A1(n_1095),
.A2(n_182),
.B(n_187),
.Y(n_1138)
);

OAI21xp33_ASAP7_75t_L g1139 ( 
.A1(n_1065),
.A2(n_329),
.B(n_190),
.Y(n_1139)
);

INVx3_ASAP7_75t_L g1140 ( 
.A(n_1129),
.Y(n_1140)
);

CKINVDCx20_ASAP7_75t_R g1141 ( 
.A(n_1135),
.Y(n_1141)
);

OR2x2_ASAP7_75t_L g1142 ( 
.A(n_1136),
.B(n_1071),
.Y(n_1142)
);

INVx2_ASAP7_75t_L g1143 ( 
.A(n_1125),
.Y(n_1143)
);

INVx3_ASAP7_75t_L g1144 ( 
.A(n_1107),
.Y(n_1144)
);

AND2x4_ASAP7_75t_L g1145 ( 
.A(n_1131),
.B(n_1068),
.Y(n_1145)
);

INVx2_ASAP7_75t_L g1146 ( 
.A(n_1105),
.Y(n_1146)
);

NOR2x1_ASAP7_75t_SL g1147 ( 
.A(n_1131),
.B(n_1086),
.Y(n_1147)
);

INVx2_ASAP7_75t_L g1148 ( 
.A(n_1105),
.Y(n_1148)
);

INVx1_ASAP7_75t_L g1149 ( 
.A(n_1137),
.Y(n_1149)
);

INVx1_ASAP7_75t_L g1150 ( 
.A(n_1126),
.Y(n_1150)
);

NOR2xp33_ASAP7_75t_L g1151 ( 
.A(n_1106),
.B(n_189),
.Y(n_1151)
);

INVx1_ASAP7_75t_L g1152 ( 
.A(n_1126),
.Y(n_1152)
);

INVx2_ASAP7_75t_L g1153 ( 
.A(n_1119),
.Y(n_1153)
);

INVx2_ASAP7_75t_L g1154 ( 
.A(n_1113),
.Y(n_1154)
);

HB1xp67_ASAP7_75t_L g1155 ( 
.A(n_1131),
.Y(n_1155)
);

AND2x2_ASAP7_75t_L g1156 ( 
.A(n_1107),
.B(n_1065),
.Y(n_1156)
);

OR2x2_ASAP7_75t_L g1157 ( 
.A(n_1109),
.B(n_192),
.Y(n_1157)
);

NAND2xp5_ASAP7_75t_L g1158 ( 
.A(n_1107),
.B(n_196),
.Y(n_1158)
);

AND2x2_ASAP7_75t_L g1159 ( 
.A(n_1108),
.B(n_198),
.Y(n_1159)
);

AND2x4_ASAP7_75t_SL g1160 ( 
.A(n_1115),
.B(n_202),
.Y(n_1160)
);

INVx2_ASAP7_75t_L g1161 ( 
.A(n_1138),
.Y(n_1161)
);

OR2x6_ASAP7_75t_L g1162 ( 
.A(n_1139),
.B(n_204),
.Y(n_1162)
);

AND2x4_ASAP7_75t_L g1163 ( 
.A(n_1132),
.B(n_316),
.Y(n_1163)
);

INVx1_ASAP7_75t_L g1164 ( 
.A(n_1123),
.Y(n_1164)
);

HB1xp67_ASAP7_75t_L g1165 ( 
.A(n_1142),
.Y(n_1165)
);

HB1xp67_ASAP7_75t_L g1166 ( 
.A(n_1150),
.Y(n_1166)
);

NAND2xp5_ASAP7_75t_L g1167 ( 
.A(n_1143),
.B(n_1112),
.Y(n_1167)
);

AND2x2_ASAP7_75t_L g1168 ( 
.A(n_1153),
.B(n_1134),
.Y(n_1168)
);

AND2x2_ASAP7_75t_L g1169 ( 
.A(n_1140),
.B(n_1130),
.Y(n_1169)
);

AO21x2_ASAP7_75t_L g1170 ( 
.A1(n_1152),
.A2(n_1104),
.B(n_1114),
.Y(n_1170)
);

AOI221xp5_ASAP7_75t_L g1171 ( 
.A1(n_1151),
.A2(n_1110),
.B1(n_1118),
.B2(n_1111),
.C(n_1121),
.Y(n_1171)
);

NOR3xp33_ASAP7_75t_L g1172 ( 
.A(n_1151),
.B(n_1122),
.C(n_1117),
.Y(n_1172)
);

AOI31xp33_ASAP7_75t_L g1173 ( 
.A1(n_1157),
.A2(n_1116),
.A3(n_1133),
.B(n_1120),
.Y(n_1173)
);

INVx2_ASAP7_75t_L g1174 ( 
.A(n_1140),
.Y(n_1174)
);

BUFx2_ASAP7_75t_L g1175 ( 
.A(n_1144),
.Y(n_1175)
);

BUFx3_ASAP7_75t_L g1176 ( 
.A(n_1141),
.Y(n_1176)
);

HB1xp67_ASAP7_75t_L g1177 ( 
.A(n_1166),
.Y(n_1177)
);

INVx1_ASAP7_75t_L g1178 ( 
.A(n_1165),
.Y(n_1178)
);

INVx3_ASAP7_75t_L g1179 ( 
.A(n_1175),
.Y(n_1179)
);

INVx2_ASAP7_75t_L g1180 ( 
.A(n_1174),
.Y(n_1180)
);

AND2x2_ASAP7_75t_L g1181 ( 
.A(n_1176),
.B(n_1156),
.Y(n_1181)
);

OR2x2_ASAP7_75t_L g1182 ( 
.A(n_1170),
.B(n_1149),
.Y(n_1182)
);

INVxp67_ASAP7_75t_SL g1183 ( 
.A(n_1168),
.Y(n_1183)
);

NAND2xp5_ASAP7_75t_L g1184 ( 
.A(n_1170),
.B(n_1146),
.Y(n_1184)
);

INVx1_ASAP7_75t_L g1185 ( 
.A(n_1167),
.Y(n_1185)
);

INVxp67_ASAP7_75t_L g1186 ( 
.A(n_1169),
.Y(n_1186)
);

NAND2xp5_ASAP7_75t_L g1187 ( 
.A(n_1186),
.B(n_1155),
.Y(n_1187)
);

NAND2x1_ASAP7_75t_SL g1188 ( 
.A(n_1177),
.B(n_1155),
.Y(n_1188)
);

INVx2_ASAP7_75t_SL g1189 ( 
.A(n_1179),
.Y(n_1189)
);

AOI22xp5_ASAP7_75t_L g1190 ( 
.A1(n_1186),
.A2(n_1172),
.B1(n_1171),
.B2(n_1162),
.Y(n_1190)
);

NAND2xp5_ASAP7_75t_L g1191 ( 
.A(n_1183),
.B(n_1164),
.Y(n_1191)
);

HB1xp67_ASAP7_75t_L g1192 ( 
.A(n_1182),
.Y(n_1192)
);

NOR2x1_ASAP7_75t_L g1193 ( 
.A(n_1185),
.B(n_1141),
.Y(n_1193)
);

CKINVDCx5p33_ASAP7_75t_R g1194 ( 
.A(n_1190),
.Y(n_1194)
);

INVx1_ASAP7_75t_L g1195 ( 
.A(n_1187),
.Y(n_1195)
);

AND2x2_ASAP7_75t_L g1196 ( 
.A(n_1193),
.B(n_1181),
.Y(n_1196)
);

OR2x2_ASAP7_75t_L g1197 ( 
.A(n_1191),
.B(n_1178),
.Y(n_1197)
);

OAI22xp5_ASAP7_75t_L g1198 ( 
.A1(n_1189),
.A2(n_1162),
.B1(n_1173),
.B2(n_1184),
.Y(n_1198)
);

NOR3xp33_ASAP7_75t_L g1199 ( 
.A(n_1192),
.B(n_1173),
.C(n_1184),
.Y(n_1199)
);

NAND2xp33_ASAP7_75t_SL g1200 ( 
.A(n_1188),
.B(n_1179),
.Y(n_1200)
);

AOI22xp33_ASAP7_75t_L g1201 ( 
.A1(n_1190),
.A2(n_1162),
.B1(n_1160),
.B2(n_1159),
.Y(n_1201)
);

INVx1_ASAP7_75t_L g1202 ( 
.A(n_1187),
.Y(n_1202)
);

INVx1_ASAP7_75t_SL g1203 ( 
.A(n_1193),
.Y(n_1203)
);

INVx1_ASAP7_75t_L g1204 ( 
.A(n_1197),
.Y(n_1204)
);

NAND2x1p5_ASAP7_75t_L g1205 ( 
.A(n_1203),
.B(n_1144),
.Y(n_1205)
);

AOI22xp5_ASAP7_75t_L g1206 ( 
.A1(n_1199),
.A2(n_1145),
.B1(n_1160),
.B2(n_1163),
.Y(n_1206)
);

INVxp67_ASAP7_75t_SL g1207 ( 
.A(n_1196),
.Y(n_1207)
);

AND2x2_ASAP7_75t_L g1208 ( 
.A(n_1195),
.B(n_1180),
.Y(n_1208)
);

OAI32xp33_ASAP7_75t_L g1209 ( 
.A1(n_1199),
.A2(n_1158),
.A3(n_1154),
.B1(n_1161),
.B2(n_1148),
.Y(n_1209)
);

NOR2xp33_ASAP7_75t_L g1210 ( 
.A(n_1207),
.B(n_1194),
.Y(n_1210)
);

NAND2xp5_ASAP7_75t_L g1211 ( 
.A(n_1204),
.B(n_1202),
.Y(n_1211)
);

AND2x4_ASAP7_75t_L g1212 ( 
.A(n_1206),
.B(n_1163),
.Y(n_1212)
);

NOR3xp33_ASAP7_75t_L g1213 ( 
.A(n_1209),
.B(n_1198),
.C(n_1200),
.Y(n_1213)
);

NAND3xp33_ASAP7_75t_L g1214 ( 
.A(n_1208),
.B(n_1201),
.C(n_1158),
.Y(n_1214)
);

OAI21xp5_ASAP7_75t_L g1215 ( 
.A1(n_1205),
.A2(n_1124),
.B(n_1127),
.Y(n_1215)
);

AND2x2_ASAP7_75t_L g1216 ( 
.A(n_1212),
.B(n_1145),
.Y(n_1216)
);

NAND2xp5_ASAP7_75t_L g1217 ( 
.A(n_1210),
.B(n_1161),
.Y(n_1217)
);

NOR2xp33_ASAP7_75t_L g1218 ( 
.A(n_1211),
.B(n_1147),
.Y(n_1218)
);

INVx1_ASAP7_75t_L g1219 ( 
.A(n_1214),
.Y(n_1219)
);

OAI32xp33_ASAP7_75t_L g1220 ( 
.A1(n_1219),
.A2(n_1213),
.A3(n_1215),
.B1(n_1128),
.B2(n_215),
.Y(n_1220)
);

INVx1_ASAP7_75t_L g1221 ( 
.A(n_1217),
.Y(n_1221)
);

INVx2_ASAP7_75t_L g1222 ( 
.A(n_1216),
.Y(n_1222)
);

AOI22xp5_ASAP7_75t_L g1223 ( 
.A1(n_1222),
.A2(n_1218),
.B1(n_207),
.B2(n_213),
.Y(n_1223)
);

AOI221xp5_ASAP7_75t_L g1224 ( 
.A1(n_1220),
.A2(n_205),
.B1(n_216),
.B2(n_217),
.C(n_218),
.Y(n_1224)
);

NAND4xp25_ASAP7_75t_L g1225 ( 
.A(n_1221),
.B(n_219),
.C(n_224),
.D(n_226),
.Y(n_1225)
);

INVx1_ASAP7_75t_L g1226 ( 
.A(n_1225),
.Y(n_1226)
);

AOI322xp5_ASAP7_75t_L g1227 ( 
.A1(n_1224),
.A2(n_228),
.A3(n_233),
.B1(n_234),
.B2(n_235),
.C1(n_246),
.C2(n_248),
.Y(n_1227)
);

INVx1_ASAP7_75t_L g1228 ( 
.A(n_1226),
.Y(n_1228)
);

AOI211xp5_ASAP7_75t_L g1229 ( 
.A1(n_1228),
.A2(n_1223),
.B(n_1227),
.C(n_256),
.Y(n_1229)
);

NOR4xp25_ASAP7_75t_L g1230 ( 
.A(n_1228),
.B(n_254),
.C(n_255),
.D(n_257),
.Y(n_1230)
);

HB1xp67_ASAP7_75t_L g1231 ( 
.A(n_1230),
.Y(n_1231)
);

XOR2xp5_ASAP7_75t_L g1232 ( 
.A(n_1229),
.B(n_258),
.Y(n_1232)
);

INVx2_ASAP7_75t_L g1233 ( 
.A(n_1232),
.Y(n_1233)
);

INVx1_ASAP7_75t_L g1234 ( 
.A(n_1231),
.Y(n_1234)
);

INVx2_ASAP7_75t_L g1235 ( 
.A(n_1232),
.Y(n_1235)
);

AOI21xp5_ASAP7_75t_L g1236 ( 
.A1(n_1234),
.A2(n_260),
.B(n_261),
.Y(n_1236)
);

XNOR2xp5_ASAP7_75t_L g1237 ( 
.A(n_1236),
.B(n_1235),
.Y(n_1237)
);

OAI22xp5_ASAP7_75t_L g1238 ( 
.A1(n_1237),
.A2(n_1233),
.B1(n_264),
.B2(n_268),
.Y(n_1238)
);

OAI22xp5_ASAP7_75t_SL g1239 ( 
.A1(n_1238),
.A2(n_263),
.B1(n_269),
.B2(n_271),
.Y(n_1239)
);

AOI22xp33_ASAP7_75t_SL g1240 ( 
.A1(n_1238),
.A2(n_275),
.B1(n_277),
.B2(n_284),
.Y(n_1240)
);

AOI22xp33_ASAP7_75t_L g1241 ( 
.A1(n_1239),
.A2(n_287),
.B1(n_288),
.B2(n_289),
.Y(n_1241)
);

OAI221xp5_ASAP7_75t_R g1242 ( 
.A1(n_1241),
.A2(n_1240),
.B1(n_291),
.B2(n_293),
.C(n_296),
.Y(n_1242)
);

AOI211xp5_ASAP7_75t_L g1243 ( 
.A1(n_1242),
.A2(n_290),
.B(n_299),
.C(n_302),
.Y(n_1243)
);


endmodule