module fake_jpeg_28739_n_122 (n_13, n_21, n_33, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_19, n_18, n_20, n_35, n_4, n_34, n_30, n_16, n_3, n_0, n_24, n_28, n_26, n_9, n_5, n_11, n_17, n_25, n_31, n_2, n_29, n_12, n_32, n_8, n_15, n_7, n_122);

input n_13;
input n_21;
input n_33;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_35;
input n_4;
input n_34;
input n_30;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_26;
input n_9;
input n_5;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_122;

wire n_117;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_73;
wire n_84;
wire n_59;
wire n_98;
wire n_65;
wire n_110;
wire n_42;
wire n_49;
wire n_76;
wire n_38;
wire n_88;
wire n_116;
wire n_114;
wire n_74;
wire n_103;
wire n_50;
wire n_57;
wire n_119;
wire n_69;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_109;
wire n_113;
wire n_106;
wire n_111;
wire n_44;
wire n_75;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_56;
wire n_79;
wire n_67;
wire n_53;
wire n_54;
wire n_93;
wire n_91;
wire n_101;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_112;
wire n_95;
wire n_97;
wire n_36;
wire n_62;
wire n_120;
wire n_43;
wire n_100;
wire n_118;
wire n_82;
wire n_96;

INVx1_ASAP7_75t_L g36 ( 
.A(n_34),
.Y(n_36)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_25),
.Y(n_37)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_1),
.Y(n_38)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_31),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_1),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_33),
.Y(n_41)
);

BUFx3_ASAP7_75t_L g42 ( 
.A(n_7),
.Y(n_42)
);

BUFx12f_ASAP7_75t_L g43 ( 
.A(n_7),
.Y(n_43)
);

BUFx5_ASAP7_75t_L g44 ( 
.A(n_2),
.Y(n_44)
);

INVx6_ASAP7_75t_SL g45 ( 
.A(n_21),
.Y(n_45)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_35),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_20),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_29),
.Y(n_48)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_9),
.Y(n_49)
);

BUFx6f_ASAP7_75t_SL g50 ( 
.A(n_32),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g51 ( 
.A(n_43),
.B(n_0),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_L g63 ( 
.A(n_51),
.B(n_49),
.Y(n_63)
);

INVx13_ASAP7_75t_L g52 ( 
.A(n_50),
.Y(n_52)
);

INVx3_ASAP7_75t_L g64 ( 
.A(n_52),
.Y(n_64)
);

INVx2_ASAP7_75t_L g53 ( 
.A(n_42),
.Y(n_53)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_53),
.Y(n_70)
);

INVx11_ASAP7_75t_L g54 ( 
.A(n_50),
.Y(n_54)
);

INVx2_ASAP7_75t_L g67 ( 
.A(n_54),
.Y(n_67)
);

CKINVDCx20_ASAP7_75t_R g55 ( 
.A(n_42),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_55),
.B(n_56),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_40),
.B(n_0),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_47),
.Y(n_57)
);

INVx2_ASAP7_75t_L g69 ( 
.A(n_57),
.Y(n_69)
);

INVx8_ASAP7_75t_L g58 ( 
.A(n_44),
.Y(n_58)
);

CKINVDCx16_ASAP7_75t_R g59 ( 
.A(n_58),
.Y(n_59)
);

CKINVDCx16_ASAP7_75t_R g60 ( 
.A(n_51),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_60),
.B(n_41),
.Y(n_71)
);

OAI22xp33_ASAP7_75t_SL g61 ( 
.A1(n_57),
.A2(n_48),
.B1(n_47),
.B2(n_45),
.Y(n_61)
);

AOI22xp5_ASAP7_75t_L g76 ( 
.A1(n_61),
.A2(n_62),
.B1(n_65),
.B2(n_66),
.Y(n_76)
);

OAI22xp5_ASAP7_75t_SL g62 ( 
.A1(n_57),
.A2(n_48),
.B1(n_43),
.B2(n_46),
.Y(n_62)
);

AND2x2_ASAP7_75t_L g81 ( 
.A(n_63),
.B(n_4),
.Y(n_81)
);

AOI22xp33_ASAP7_75t_L g65 ( 
.A1(n_53),
.A2(n_43),
.B1(n_44),
.B2(n_38),
.Y(n_65)
);

AOI22xp5_ASAP7_75t_L g66 ( 
.A1(n_55),
.A2(n_46),
.B1(n_36),
.B2(n_39),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_71),
.B(n_73),
.Y(n_90)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_66),
.Y(n_72)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_72),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_68),
.B(n_36),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_L g74 ( 
.A(n_70),
.B(n_37),
.Y(n_74)
);

OAI22xp5_ASAP7_75t_L g89 ( 
.A1(n_74),
.A2(n_77),
.B1(n_79),
.B2(n_82),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_SL g75 ( 
.A(n_61),
.B(n_2),
.Y(n_75)
);

OAI21xp5_ASAP7_75t_SL g93 ( 
.A1(n_75),
.A2(n_81),
.B(n_85),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_L g77 ( 
.A(n_62),
.B(n_3),
.Y(n_77)
);

BUFx3_ASAP7_75t_L g78 ( 
.A(n_64),
.Y(n_78)
);

INVx2_ASAP7_75t_SL g91 ( 
.A(n_78),
.Y(n_91)
);

AOI22xp33_ASAP7_75t_SL g79 ( 
.A1(n_69),
.A2(n_58),
.B1(n_45),
.B2(n_52),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_SL g80 ( 
.A(n_59),
.B(n_3),
.Y(n_80)
);

CKINVDCx20_ASAP7_75t_R g94 ( 
.A(n_80),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_L g82 ( 
.A(n_64),
.B(n_4),
.Y(n_82)
);

OAI21xp5_ASAP7_75t_L g83 ( 
.A1(n_67),
.A2(n_54),
.B(n_6),
.Y(n_83)
);

XNOR2xp5_ASAP7_75t_L g96 ( 
.A(n_83),
.B(n_10),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_63),
.B(n_5),
.Y(n_84)
);

CKINVDCx16_ASAP7_75t_R g97 ( 
.A(n_84),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_SL g85 ( 
.A(n_60),
.B(n_5),
.Y(n_85)
);

AOI22xp5_ASAP7_75t_L g86 ( 
.A1(n_76),
.A2(n_83),
.B1(n_81),
.B2(n_79),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_L g103 ( 
.A(n_86),
.B(n_92),
.Y(n_103)
);

CKINVDCx10_ASAP7_75t_R g87 ( 
.A(n_78),
.Y(n_87)
);

CKINVDCx20_ASAP7_75t_R g104 ( 
.A(n_87),
.Y(n_104)
);

OAI22xp5_ASAP7_75t_SL g92 ( 
.A1(n_76),
.A2(n_6),
.B1(n_8),
.B2(n_9),
.Y(n_92)
);

OAI22xp5_ASAP7_75t_L g95 ( 
.A1(n_72),
.A2(n_8),
.B1(n_10),
.B2(n_11),
.Y(n_95)
);

OAI21xp5_ASAP7_75t_SL g107 ( 
.A1(n_95),
.A2(n_101),
.B(n_15),
.Y(n_107)
);

XOR2xp5_ASAP7_75t_L g110 ( 
.A(n_96),
.B(n_18),
.Y(n_110)
);

INVxp67_ASAP7_75t_L g98 ( 
.A(n_83),
.Y(n_98)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_98),
.Y(n_105)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_74),
.Y(n_99)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_99),
.Y(n_106)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_74),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_SL g102 ( 
.A(n_100),
.B(n_14),
.Y(n_102)
);

OAI22xp5_ASAP7_75t_L g101 ( 
.A1(n_72),
.A2(n_11),
.B1(n_12),
.B2(n_13),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_SL g114 ( 
.A(n_102),
.B(n_107),
.Y(n_114)
);

OAI21xp5_ASAP7_75t_SL g108 ( 
.A1(n_98),
.A2(n_16),
.B(n_17),
.Y(n_108)
);

MAJIxp5_ASAP7_75t_L g113 ( 
.A(n_108),
.B(n_110),
.C(n_97),
.Y(n_113)
);

OAI21xp5_ASAP7_75t_L g109 ( 
.A1(n_88),
.A2(n_96),
.B(n_89),
.Y(n_109)
);

A2O1A1O1Ixp25_ASAP7_75t_L g111 ( 
.A1(n_109),
.A2(n_105),
.B(n_103),
.C(n_106),
.D(n_110),
.Y(n_111)
);

OAI22xp5_ASAP7_75t_SL g115 ( 
.A1(n_111),
.A2(n_112),
.B1(n_113),
.B2(n_109),
.Y(n_115)
);

CKINVDCx20_ASAP7_75t_R g112 ( 
.A(n_104),
.Y(n_112)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_115),
.Y(n_117)
);

OAI321xp33_ASAP7_75t_L g116 ( 
.A1(n_111),
.A2(n_93),
.A3(n_94),
.B1(n_90),
.B2(n_87),
.C(n_26),
.Y(n_116)
);

AOI221xp5_ASAP7_75t_L g118 ( 
.A1(n_117),
.A2(n_116),
.B1(n_114),
.B2(n_91),
.C(n_24),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_L g119 ( 
.A(n_118),
.B(n_19),
.Y(n_119)
);

CKINVDCx20_ASAP7_75t_R g120 ( 
.A(n_119),
.Y(n_120)
);

OAI321xp33_ASAP7_75t_L g121 ( 
.A1(n_120),
.A2(n_91),
.A3(n_23),
.B1(n_27),
.B2(n_28),
.C(n_30),
.Y(n_121)
);

XNOR2xp5_ASAP7_75t_L g122 ( 
.A(n_121),
.B(n_22),
.Y(n_122)
);


endmodule