module fake_jpeg_15839_n_109 (n_11, n_3, n_2, n_1, n_0, n_10, n_4, n_8, n_9, n_6, n_5, n_7, n_109);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_109;

wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_74;
wire n_31;
wire n_29;
wire n_103;
wire n_50;
wire n_15;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_30;
wire n_106;
wire n_24;
wire n_44;
wire n_25;
wire n_17;
wire n_75;
wire n_37;
wire n_102;
wire n_99;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_18;
wire n_20;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_56;
wire n_79;
wire n_12;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_22;
wire n_101;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_95;
wire n_97;
wire n_36;
wire n_62;
wire n_43;
wire n_32;
wire n_100;
wire n_82;
wire n_96;

INVx1_ASAP7_75t_SL g12 ( 
.A(n_7),
.Y(n_12)
);

INVx5_ASAP7_75t_L g13 ( 
.A(n_0),
.Y(n_13)
);

INVx1_ASAP7_75t_L g14 ( 
.A(n_11),
.Y(n_14)
);

INVx1_ASAP7_75t_L g15 ( 
.A(n_2),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_0),
.Y(n_16)
);

BUFx3_ASAP7_75t_L g17 ( 
.A(n_9),
.Y(n_17)
);

INVx2_ASAP7_75t_L g18 ( 
.A(n_10),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_3),
.Y(n_19)
);

BUFx3_ASAP7_75t_L g20 ( 
.A(n_2),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_11),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_9),
.Y(n_22)
);

INVx13_ASAP7_75t_L g23 ( 
.A(n_8),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_8),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_5),
.Y(n_25)
);

AOI22xp33_ASAP7_75t_SL g26 ( 
.A1(n_12),
.A2(n_6),
.B1(n_10),
.B2(n_2),
.Y(n_26)
);

AOI22xp33_ASAP7_75t_SL g47 ( 
.A1(n_26),
.A2(n_22),
.B1(n_13),
.B2(n_15),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g27 ( 
.A(n_12),
.B(n_11),
.Y(n_27)
);

NOR2xp33_ASAP7_75t_SL g38 ( 
.A(n_27),
.B(n_24),
.Y(n_38)
);

AOI22xp5_ASAP7_75t_L g28 ( 
.A1(n_18),
.A2(n_0),
.B1(n_1),
.B2(n_3),
.Y(n_28)
);

MAJIxp5_ASAP7_75t_L g41 ( 
.A(n_28),
.B(n_30),
.C(n_31),
.Y(n_41)
);

INVx2_ASAP7_75t_L g29 ( 
.A(n_18),
.Y(n_29)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_29),
.Y(n_39)
);

OAI22xp5_ASAP7_75t_SL g30 ( 
.A1(n_18),
.A2(n_0),
.B1(n_1),
.B2(n_3),
.Y(n_30)
);

OAI22xp5_ASAP7_75t_L g31 ( 
.A1(n_13),
.A2(n_1),
.B1(n_4),
.B2(n_5),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_14),
.Y(n_32)
);

NOR2xp33_ASAP7_75t_L g43 ( 
.A(n_32),
.B(n_33),
.Y(n_43)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_14),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_21),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_34),
.B(n_35),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_21),
.Y(n_35)
);

NAND2xp5_ASAP7_75t_L g36 ( 
.A(n_29),
.B(n_24),
.Y(n_36)
);

NAND2xp5_ASAP7_75t_L g62 ( 
.A(n_36),
.B(n_45),
.Y(n_62)
);

NOR2x1_ASAP7_75t_L g37 ( 
.A(n_32),
.B(n_12),
.Y(n_37)
);

NAND2xp5_ASAP7_75t_SL g60 ( 
.A(n_37),
.B(n_42),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g51 ( 
.A(n_38),
.B(n_50),
.Y(n_51)
);

INVx5_ASAP7_75t_L g40 ( 
.A(n_34),
.Y(n_40)
);

INVx5_ASAP7_75t_L g64 ( 
.A(n_40),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_SL g42 ( 
.A(n_33),
.B(n_15),
.Y(n_42)
);

OA22x2_ASAP7_75t_L g44 ( 
.A1(n_28),
.A2(n_13),
.B1(n_23),
.B2(n_16),
.Y(n_44)
);

AOI22xp5_ASAP7_75t_L g53 ( 
.A1(n_44),
.A2(n_46),
.B1(n_31),
.B2(n_23),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_L g45 ( 
.A(n_28),
.B(n_24),
.Y(n_45)
);

AOI21xp33_ASAP7_75t_L g46 ( 
.A1(n_27),
.A2(n_22),
.B(n_16),
.Y(n_46)
);

AOI22xp33_ASAP7_75t_SL g63 ( 
.A1(n_47),
.A2(n_19),
.B1(n_23),
.B2(n_5),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_L g49 ( 
.A(n_30),
.B(n_22),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_SL g66 ( 
.A(n_49),
.B(n_1),
.Y(n_66)
);

INVx5_ASAP7_75t_L g50 ( 
.A(n_34),
.Y(n_50)
);

CKINVDCx16_ASAP7_75t_R g52 ( 
.A(n_36),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_52),
.B(n_57),
.Y(n_71)
);

XNOR2xp5_ASAP7_75t_SL g74 ( 
.A(n_53),
.B(n_65),
.Y(n_74)
);

OAI22xp5_ASAP7_75t_L g54 ( 
.A1(n_41),
.A2(n_26),
.B1(n_34),
.B2(n_35),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_L g78 ( 
.A(n_54),
.B(n_55),
.Y(n_78)
);

CKINVDCx20_ASAP7_75t_R g55 ( 
.A(n_43),
.Y(n_55)
);

OAI22xp5_ASAP7_75t_SL g56 ( 
.A1(n_41),
.A2(n_23),
.B1(n_35),
.B2(n_25),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_56),
.B(n_59),
.Y(n_77)
);

OAI22xp5_ASAP7_75t_L g57 ( 
.A1(n_41),
.A2(n_35),
.B1(n_21),
.B2(n_25),
.Y(n_57)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_48),
.Y(n_58)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_58),
.Y(n_76)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_48),
.Y(n_59)
);

OAI22xp5_ASAP7_75t_L g61 ( 
.A1(n_45),
.A2(n_21),
.B1(n_19),
.B2(n_20),
.Y(n_61)
);

O2A1O1Ixp33_ASAP7_75t_L g75 ( 
.A1(n_61),
.A2(n_63),
.B(n_47),
.C(n_44),
.Y(n_75)
);

AOI22xp5_ASAP7_75t_L g65 ( 
.A1(n_49),
.A2(n_8),
.B1(n_4),
.B2(n_6),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_L g73 ( 
.A(n_66),
.B(n_44),
.Y(n_73)
);

MAJIxp5_ASAP7_75t_L g67 ( 
.A(n_62),
.B(n_39),
.C(n_37),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_L g79 ( 
.A(n_67),
.B(n_70),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_SL g68 ( 
.A(n_55),
.B(n_43),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_68),
.B(n_69),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_SL g69 ( 
.A(n_60),
.B(n_42),
.Y(n_69)
);

MAJIxp5_ASAP7_75t_L g70 ( 
.A(n_62),
.B(n_39),
.C(n_37),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_SL g72 ( 
.A(n_60),
.B(n_38),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_72),
.B(n_73),
.Y(n_87)
);

AOI22xp5_ASAP7_75t_SL g83 ( 
.A1(n_75),
.A2(n_44),
.B1(n_59),
.B2(n_64),
.Y(n_83)
);

OAI22xp5_ASAP7_75t_L g80 ( 
.A1(n_78),
.A2(n_53),
.B1(n_52),
.B2(n_54),
.Y(n_80)
);

OAI22xp5_ASAP7_75t_L g90 ( 
.A1(n_80),
.A2(n_81),
.B1(n_82),
.B2(n_83),
.Y(n_90)
);

OAI22xp5_ASAP7_75t_L g81 ( 
.A1(n_77),
.A2(n_56),
.B1(n_57),
.B2(n_50),
.Y(n_81)
);

AOI22xp5_ASAP7_75t_L g82 ( 
.A1(n_71),
.A2(n_61),
.B1(n_66),
.B2(n_58),
.Y(n_82)
);

HB1xp67_ASAP7_75t_L g84 ( 
.A(n_76),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_84),
.B(n_64),
.Y(n_93)
);

OAI22xp5_ASAP7_75t_L g85 ( 
.A1(n_75),
.A2(n_40),
.B1(n_50),
.B2(n_44),
.Y(n_85)
);

OAI22xp5_ASAP7_75t_L g94 ( 
.A1(n_85),
.A2(n_88),
.B1(n_51),
.B2(n_20),
.Y(n_94)
);

OAI22xp5_ASAP7_75t_SL g88 ( 
.A1(n_73),
.A2(n_44),
.B1(n_40),
.B2(n_65),
.Y(n_88)
);

MAJIxp5_ASAP7_75t_L g89 ( 
.A(n_79),
.B(n_80),
.C(n_74),
.Y(n_89)
);

XNOR2xp5_ASAP7_75t_L g98 ( 
.A(n_89),
.B(n_91),
.Y(n_98)
);

MAJIxp5_ASAP7_75t_L g91 ( 
.A(n_79),
.B(n_74),
.C(n_70),
.Y(n_91)
);

MAJx2_ASAP7_75t_L g92 ( 
.A(n_87),
.B(n_67),
.C(n_46),
.Y(n_92)
);

AND2x2_ASAP7_75t_L g96 ( 
.A(n_92),
.B(n_82),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g100 ( 
.A(n_93),
.B(n_95),
.Y(n_100)
);

AOI22xp5_ASAP7_75t_L g97 ( 
.A1(n_94),
.A2(n_85),
.B1(n_90),
.B2(n_81),
.Y(n_97)
);

CKINVDCx20_ASAP7_75t_R g95 ( 
.A(n_86),
.Y(n_95)
);

OAI321xp33_ASAP7_75t_L g103 ( 
.A1(n_97),
.A2(n_96),
.A3(n_100),
.B1(n_98),
.B2(n_17),
.C(n_4),
.Y(n_103)
);

AOI21xp5_ASAP7_75t_L g99 ( 
.A1(n_92),
.A2(n_83),
.B(n_86),
.Y(n_99)
);

MAJIxp5_ASAP7_75t_L g101 ( 
.A(n_99),
.B(n_89),
.C(n_91),
.Y(n_101)
);

MAJIxp5_ASAP7_75t_L g105 ( 
.A(n_101),
.B(n_102),
.C(n_6),
.Y(n_105)
);

MAJIxp5_ASAP7_75t_L g102 ( 
.A(n_98),
.B(n_88),
.C(n_20),
.Y(n_102)
);

OAI22xp5_ASAP7_75t_SL g104 ( 
.A1(n_103),
.A2(n_97),
.B1(n_17),
.B2(n_9),
.Y(n_104)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_104),
.Y(n_107)
);

OAI21x1_ASAP7_75t_L g106 ( 
.A1(n_103),
.A2(n_7),
.B(n_10),
.Y(n_106)
);

OAI21xp5_ASAP7_75t_L g108 ( 
.A1(n_107),
.A2(n_105),
.B(n_106),
.Y(n_108)
);

BUFx24_ASAP7_75t_SL g109 ( 
.A(n_108),
.Y(n_109)
);


endmodule