module fake_jpeg_1429_n_43 (n_11, n_3, n_2, n_1, n_0, n_10, n_4, n_8, n_9, n_6, n_5, n_7, n_43);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_43;

wire n_13;
wire n_21;
wire n_33;
wire n_23;
wire n_27;
wire n_22;
wire n_14;
wire n_40;
wire n_19;
wire n_18;
wire n_20;
wire n_35;
wire n_41;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_16;
wire n_24;
wire n_28;
wire n_38;
wire n_26;
wire n_36;
wire n_17;
wire n_25;
wire n_31;
wire n_29;
wire n_37;
wire n_12;
wire n_32;
wire n_15;

BUFx6f_ASAP7_75t_L g12 ( 
.A(n_3),
.Y(n_12)
);

INVx5_ASAP7_75t_L g13 ( 
.A(n_11),
.Y(n_13)
);

CKINVDCx20_ASAP7_75t_R g14 ( 
.A(n_6),
.Y(n_14)
);

INVx8_ASAP7_75t_L g15 ( 
.A(n_0),
.Y(n_15)
);

BUFx6f_ASAP7_75t_L g16 ( 
.A(n_4),
.Y(n_16)
);

AOI22xp5_ASAP7_75t_L g17 ( 
.A1(n_12),
.A2(n_10),
.B1(n_9),
.B2(n_2),
.Y(n_17)
);

AOI22xp5_ASAP7_75t_L g20 ( 
.A1(n_17),
.A2(n_14),
.B1(n_16),
.B2(n_12),
.Y(n_20)
);

INVx2_ASAP7_75t_SL g18 ( 
.A(n_13),
.Y(n_18)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_18),
.Y(n_23)
);

NAND2xp5_ASAP7_75t_L g19 ( 
.A(n_16),
.B(n_0),
.Y(n_19)
);

CKINVDCx14_ASAP7_75t_R g21 ( 
.A(n_19),
.Y(n_21)
);

OA21x2_ASAP7_75t_L g27 ( 
.A1(n_20),
.A2(n_22),
.B(n_17),
.Y(n_27)
);

AOI22xp5_ASAP7_75t_L g22 ( 
.A1(n_19),
.A2(n_16),
.B1(n_12),
.B2(n_15),
.Y(n_22)
);

AND2x6_ASAP7_75t_L g24 ( 
.A(n_21),
.B(n_1),
.Y(n_24)
);

MAJIxp5_ASAP7_75t_L g30 ( 
.A(n_24),
.B(n_1),
.C(n_2),
.Y(n_30)
);

NOR2xp33_ASAP7_75t_SL g25 ( 
.A(n_23),
.B(n_14),
.Y(n_25)
);

NAND2xp5_ASAP7_75t_L g31 ( 
.A(n_25),
.B(n_26),
.Y(n_31)
);

NAND2xp5_ASAP7_75t_SL g26 ( 
.A(n_22),
.B(n_18),
.Y(n_26)
);

AOI22xp5_ASAP7_75t_SL g29 ( 
.A1(n_27),
.A2(n_13),
.B1(n_15),
.B2(n_3),
.Y(n_29)
);

AOI21xp5_ASAP7_75t_L g28 ( 
.A1(n_25),
.A2(n_20),
.B(n_18),
.Y(n_28)
);

INVxp67_ASAP7_75t_L g33 ( 
.A(n_28),
.Y(n_33)
);

NAND2xp5_ASAP7_75t_SL g35 ( 
.A(n_29),
.B(n_30),
.Y(n_35)
);

XNOR2xp5_ASAP7_75t_SL g32 ( 
.A(n_31),
.B(n_4),
.Y(n_32)
);

MAJIxp5_ASAP7_75t_L g36 ( 
.A(n_32),
.B(n_34),
.C(n_5),
.Y(n_36)
);

XOR2xp5_ASAP7_75t_L g34 ( 
.A(n_31),
.B(n_5),
.Y(n_34)
);

NAND2xp5_ASAP7_75t_L g40 ( 
.A(n_36),
.B(n_37),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g37 ( 
.A(n_35),
.B(n_33),
.Y(n_37)
);

AND2x2_ASAP7_75t_L g38 ( 
.A(n_33),
.B(n_6),
.Y(n_38)
);

NAND2xp5_ASAP7_75t_SL g39 ( 
.A(n_38),
.B(n_7),
.Y(n_39)
);

NOR2x1_ASAP7_75t_L g41 ( 
.A(n_39),
.B(n_7),
.Y(n_41)
);

MAJIxp5_ASAP7_75t_L g42 ( 
.A(n_41),
.B(n_40),
.C(n_8),
.Y(n_42)
);

MAJIxp5_ASAP7_75t_L g43 ( 
.A(n_42),
.B(n_41),
.C(n_8),
.Y(n_43)
);


endmodule