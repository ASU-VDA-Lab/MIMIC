module fake_jpeg_29526_n_507 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_507);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_507;

wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_17;
wire n_431;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_490;
wire n_415;
wire n_479;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_48;
wire n_465;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_221;
wire n_256;
wire n_454;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_474;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_305;
wire n_161;
wire n_441;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_352;
wire n_350;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_296;
wire n_384;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_491;
wire n_24;
wire n_467;
wire n_269;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_473;
wire n_45;
wire n_476;
wire n_337;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_481;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_199;
wire n_260;
wire n_413;
wire n_275;
wire n_494;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_492;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_472;
wire n_279;
wire n_154;
wire n_495;
wire n_205;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_484;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_469;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_482;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_183;
wire n_409;
wire n_249;
wire n_412;
wire n_217;
wire n_471;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_402;
wire n_504;
wire n_438;
wire n_475;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

BUFx10_ASAP7_75t_L g17 ( 
.A(n_6),
.Y(n_17)
);

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_14),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_16),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_10),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_4),
.Y(n_21)
);

BUFx4f_ASAP7_75t_L g22 ( 
.A(n_5),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_15),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_10),
.Y(n_24)
);

BUFx4f_ASAP7_75t_SL g25 ( 
.A(n_14),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_0),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_0),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_9),
.Y(n_28)
);

BUFx3_ASAP7_75t_L g29 ( 
.A(n_9),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_16),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_8),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_8),
.Y(n_32)
);

BUFx12f_ASAP7_75t_L g33 ( 
.A(n_14),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_16),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_7),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_12),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_12),
.Y(n_37)
);

INVx2_ASAP7_75t_L g38 ( 
.A(n_6),
.Y(n_38)
);

BUFx12f_ASAP7_75t_L g39 ( 
.A(n_7),
.Y(n_39)
);

BUFx3_ASAP7_75t_L g40 ( 
.A(n_2),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_6),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_3),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_10),
.Y(n_43)
);

BUFx4f_ASAP7_75t_L g44 ( 
.A(n_0),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_15),
.Y(n_45)
);

BUFx10_ASAP7_75t_L g46 ( 
.A(n_16),
.Y(n_46)
);

HB1xp67_ASAP7_75t_L g47 ( 
.A(n_4),
.Y(n_47)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_3),
.Y(n_48)
);

CKINVDCx14_ASAP7_75t_R g49 ( 
.A(n_12),
.Y(n_49)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_11),
.Y(n_50)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_14),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_L g52 ( 
.A(n_24),
.B(n_7),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_L g149 ( 
.A(n_52),
.B(n_66),
.Y(n_149)
);

INVx4_ASAP7_75t_L g53 ( 
.A(n_29),
.Y(n_53)
);

INVx3_ASAP7_75t_SL g136 ( 
.A(n_53),
.Y(n_136)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_20),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g105 ( 
.A(n_54),
.Y(n_105)
);

INVx6_ASAP7_75t_SL g55 ( 
.A(n_22),
.Y(n_55)
);

CKINVDCx14_ASAP7_75t_R g109 ( 
.A(n_55),
.Y(n_109)
);

INVx5_ASAP7_75t_L g56 ( 
.A(n_29),
.Y(n_56)
);

INVx5_ASAP7_75t_L g104 ( 
.A(n_56),
.Y(n_104)
);

INVx4_ASAP7_75t_SL g57 ( 
.A(n_38),
.Y(n_57)
);

INVx2_ASAP7_75t_SL g145 ( 
.A(n_57),
.Y(n_145)
);

HAxp5_ASAP7_75t_SL g58 ( 
.A(n_44),
.B(n_15),
.CON(n_58),
.SN(n_58)
);

AND2x2_ASAP7_75t_L g123 ( 
.A(n_58),
.B(n_61),
.Y(n_123)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_38),
.Y(n_59)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_59),
.Y(n_110)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_47),
.Y(n_60)
);

INVx2_ASAP7_75t_L g114 ( 
.A(n_60),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_24),
.B(n_51),
.Y(n_61)
);

BUFx3_ASAP7_75t_L g62 ( 
.A(n_29),
.Y(n_62)
);

INVx5_ASAP7_75t_L g129 ( 
.A(n_62),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_SL g63 ( 
.A(n_28),
.B(n_7),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g122 ( 
.A(n_63),
.B(n_64),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_28),
.B(n_8),
.Y(n_64)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_47),
.Y(n_65)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_65),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_L g66 ( 
.A(n_32),
.B(n_8),
.Y(n_66)
);

BUFx24_ASAP7_75t_L g67 ( 
.A(n_22),
.Y(n_67)
);

BUFx2_ASAP7_75t_L g107 ( 
.A(n_67),
.Y(n_107)
);

BUFx5_ASAP7_75t_L g68 ( 
.A(n_33),
.Y(n_68)
);

INVx5_ASAP7_75t_L g140 ( 
.A(n_68),
.Y(n_140)
);

INVx2_ASAP7_75t_L g69 ( 
.A(n_40),
.Y(n_69)
);

INVx2_ASAP7_75t_L g124 ( 
.A(n_69),
.Y(n_124)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_40),
.Y(n_70)
);

INVx2_ASAP7_75t_L g130 ( 
.A(n_70),
.Y(n_130)
);

BUFx6f_ASAP7_75t_L g71 ( 
.A(n_20),
.Y(n_71)
);

BUFx6f_ASAP7_75t_L g111 ( 
.A(n_71),
.Y(n_111)
);

CKINVDCx20_ASAP7_75t_R g72 ( 
.A(n_17),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g126 ( 
.A(n_72),
.B(n_76),
.Y(n_126)
);

INVx2_ASAP7_75t_L g73 ( 
.A(n_40),
.Y(n_73)
);

INVx2_ASAP7_75t_L g131 ( 
.A(n_73),
.Y(n_131)
);

INVx6_ASAP7_75t_L g74 ( 
.A(n_20),
.Y(n_74)
);

BUFx6f_ASAP7_75t_L g138 ( 
.A(n_74),
.Y(n_138)
);

INVx2_ASAP7_75t_L g75 ( 
.A(n_20),
.Y(n_75)
);

INVx2_ASAP7_75t_L g146 ( 
.A(n_75),
.Y(n_146)
);

CKINVDCx20_ASAP7_75t_R g76 ( 
.A(n_17),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_L g77 ( 
.A(n_32),
.B(n_6),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_SL g102 ( 
.A(n_77),
.B(n_51),
.Y(n_102)
);

BUFx3_ASAP7_75t_L g78 ( 
.A(n_31),
.Y(n_78)
);

INVx5_ASAP7_75t_L g152 ( 
.A(n_78),
.Y(n_152)
);

BUFx6f_ASAP7_75t_L g79 ( 
.A(n_31),
.Y(n_79)
);

BUFx6f_ASAP7_75t_L g151 ( 
.A(n_79),
.Y(n_151)
);

INVx2_ASAP7_75t_L g80 ( 
.A(n_31),
.Y(n_80)
);

INVx2_ASAP7_75t_L g103 ( 
.A(n_80),
.Y(n_103)
);

BUFx6f_ASAP7_75t_L g81 ( 
.A(n_31),
.Y(n_81)
);

INVx6_ASAP7_75t_L g120 ( 
.A(n_81),
.Y(n_120)
);

BUFx6f_ASAP7_75t_L g82 ( 
.A(n_18),
.Y(n_82)
);

INVx6_ASAP7_75t_L g148 ( 
.A(n_82),
.Y(n_148)
);

INVx2_ASAP7_75t_L g83 ( 
.A(n_44),
.Y(n_83)
);

INVx2_ASAP7_75t_L g112 ( 
.A(n_83),
.Y(n_112)
);

BUFx16f_ASAP7_75t_L g84 ( 
.A(n_22),
.Y(n_84)
);

CKINVDCx16_ASAP7_75t_R g116 ( 
.A(n_84),
.Y(n_116)
);

INVx2_ASAP7_75t_L g85 ( 
.A(n_44),
.Y(n_85)
);

INVx2_ASAP7_75t_L g119 ( 
.A(n_85),
.Y(n_119)
);

INVx4_ASAP7_75t_L g86 ( 
.A(n_22),
.Y(n_86)
);

INVx4_ASAP7_75t_L g134 ( 
.A(n_86),
.Y(n_134)
);

CKINVDCx20_ASAP7_75t_R g87 ( 
.A(n_17),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g133 ( 
.A(n_87),
.B(n_89),
.Y(n_133)
);

INVx3_ASAP7_75t_L g88 ( 
.A(n_33),
.Y(n_88)
);

INVx3_ASAP7_75t_L g108 ( 
.A(n_88),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_37),
.B(n_9),
.Y(n_89)
);

BUFx6f_ASAP7_75t_L g90 ( 
.A(n_18),
.Y(n_90)
);

INVx4_ASAP7_75t_L g156 ( 
.A(n_90),
.Y(n_156)
);

BUFx6f_ASAP7_75t_L g91 ( 
.A(n_18),
.Y(n_91)
);

INVx3_ASAP7_75t_L g132 ( 
.A(n_91),
.Y(n_132)
);

INVx6_ASAP7_75t_L g92 ( 
.A(n_30),
.Y(n_92)
);

INVx3_ASAP7_75t_L g135 ( 
.A(n_92),
.Y(n_135)
);

BUFx6f_ASAP7_75t_L g93 ( 
.A(n_30),
.Y(n_93)
);

HB1xp67_ASAP7_75t_L g139 ( 
.A(n_93),
.Y(n_139)
);

CKINVDCx20_ASAP7_75t_R g94 ( 
.A(n_17),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g141 ( 
.A(n_94),
.B(n_95),
.Y(n_141)
);

BUFx3_ASAP7_75t_L g95 ( 
.A(n_30),
.Y(n_95)
);

CKINVDCx20_ASAP7_75t_R g96 ( 
.A(n_17),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g154 ( 
.A(n_96),
.B(n_97),
.Y(n_154)
);

CKINVDCx20_ASAP7_75t_R g97 ( 
.A(n_46),
.Y(n_97)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_19),
.Y(n_98)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_98),
.Y(n_125)
);

BUFx5_ASAP7_75t_L g99 ( 
.A(n_33),
.Y(n_99)
);

OR2x2_ASAP7_75t_L g106 ( 
.A(n_99),
.B(n_33),
.Y(n_106)
);

INVx4_ASAP7_75t_L g100 ( 
.A(n_41),
.Y(n_100)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_100),
.Y(n_127)
);

OAI21xp33_ASAP7_75t_L g101 ( 
.A1(n_58),
.A2(n_49),
.B(n_50),
.Y(n_101)
);

O2A1O1Ixp33_ASAP7_75t_L g183 ( 
.A1(n_101),
.A2(n_25),
.B(n_46),
.C(n_68),
.Y(n_183)
);

NOR2xp33_ASAP7_75t_L g170 ( 
.A(n_102),
.B(n_128),
.Y(n_170)
);

CKINVDCx16_ASAP7_75t_R g161 ( 
.A(n_106),
.Y(n_161)
);

OAI22xp5_ASAP7_75t_L g113 ( 
.A1(n_82),
.A2(n_41),
.B1(n_37),
.B2(n_45),
.Y(n_113)
);

AOI22xp5_ASAP7_75t_L g187 ( 
.A1(n_113),
.A2(n_115),
.B1(n_117),
.B2(n_121),
.Y(n_187)
);

OAI22xp5_ASAP7_75t_L g115 ( 
.A1(n_90),
.A2(n_41),
.B1(n_45),
.B2(n_43),
.Y(n_115)
);

OAI22xp33_ASAP7_75t_SL g117 ( 
.A1(n_92),
.A2(n_27),
.B1(n_44),
.B2(n_35),
.Y(n_117)
);

OAI22xp5_ASAP7_75t_L g121 ( 
.A1(n_91),
.A2(n_43),
.B1(n_42),
.B2(n_27),
.Y(n_121)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_60),
.Y(n_128)
);

OAI22xp5_ASAP7_75t_L g137 ( 
.A1(n_93),
.A2(n_42),
.B1(n_27),
.B2(n_49),
.Y(n_137)
);

AOI22xp33_ASAP7_75t_L g158 ( 
.A1(n_137),
.A2(n_21),
.B1(n_35),
.B2(n_36),
.Y(n_158)
);

AOI22xp33_ASAP7_75t_SL g142 ( 
.A1(n_55),
.A2(n_39),
.B1(n_33),
.B2(n_50),
.Y(n_142)
);

AOI22xp33_ASAP7_75t_SL g184 ( 
.A1(n_142),
.A2(n_155),
.B1(n_145),
.B2(n_109),
.Y(n_184)
);

AOI22xp33_ASAP7_75t_L g143 ( 
.A1(n_74),
.A2(n_39),
.B1(n_26),
.B2(n_48),
.Y(n_143)
);

OAI22xp5_ASAP7_75t_SL g169 ( 
.A1(n_143),
.A2(n_26),
.B1(n_23),
.B2(n_36),
.Y(n_169)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_57),
.Y(n_144)
);

NOR2xp33_ASAP7_75t_L g194 ( 
.A(n_144),
.B(n_150),
.Y(n_194)
);

A2O1A1Ixp33_ASAP7_75t_L g147 ( 
.A1(n_84),
.A2(n_48),
.B(n_34),
.C(n_19),
.Y(n_147)
);

OAI21xp5_ASAP7_75t_SL g207 ( 
.A1(n_147),
.A2(n_11),
.B(n_13),
.Y(n_207)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_75),
.Y(n_150)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_80),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_L g196 ( 
.A(n_153),
.B(n_157),
.Y(n_196)
);

AOI22xp33_ASAP7_75t_SL g155 ( 
.A1(n_95),
.A2(n_100),
.B1(n_78),
.B2(n_62),
.Y(n_155)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_69),
.Y(n_157)
);

OAI22xp5_ASAP7_75t_SL g224 ( 
.A1(n_158),
.A2(n_178),
.B1(n_206),
.B2(n_156),
.Y(n_224)
);

CKINVDCx20_ASAP7_75t_R g159 ( 
.A(n_126),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_SL g212 ( 
.A(n_159),
.B(n_163),
.Y(n_212)
);

AOI32xp33_ASAP7_75t_L g160 ( 
.A1(n_123),
.A2(n_53),
.A3(n_84),
.B1(n_86),
.B2(n_88),
.Y(n_160)
);

AOI32xp33_ASAP7_75t_L g250 ( 
.A1(n_160),
.A2(n_138),
.A3(n_111),
.B1(n_151),
.B2(n_1),
.Y(n_250)
);

OAI22xp5_ASAP7_75t_L g162 ( 
.A1(n_149),
.A2(n_54),
.B1(n_71),
.B2(n_79),
.Y(n_162)
);

AOI22xp5_ASAP7_75t_L g210 ( 
.A1(n_162),
.A2(n_164),
.B1(n_169),
.B2(n_180),
.Y(n_210)
);

CKINVDCx20_ASAP7_75t_R g163 ( 
.A(n_154),
.Y(n_163)
);

OAI22xp5_ASAP7_75t_L g164 ( 
.A1(n_123),
.A2(n_81),
.B1(n_70),
.B2(n_73),
.Y(n_164)
);

INVx2_ASAP7_75t_L g165 ( 
.A(n_112),
.Y(n_165)
);

INVx2_ASAP7_75t_L g213 ( 
.A(n_165),
.Y(n_213)
);

CKINVDCx20_ASAP7_75t_R g166 ( 
.A(n_141),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_SL g235 ( 
.A(n_166),
.B(n_179),
.Y(n_235)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_110),
.Y(n_167)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_167),
.Y(n_211)
);

NAND2xp5_ASAP7_75t_SL g168 ( 
.A(n_147),
.B(n_85),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_L g233 ( 
.A(n_168),
.B(n_175),
.Y(n_233)
);

BUFx6f_ASAP7_75t_L g171 ( 
.A(n_105),
.Y(n_171)
);

INVx5_ASAP7_75t_L g214 ( 
.A(n_171),
.Y(n_214)
);

INVx1_ASAP7_75t_SL g172 ( 
.A(n_106),
.Y(n_172)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_172),
.Y(n_216)
);

A2O1A1Ixp33_ASAP7_75t_L g173 ( 
.A1(n_101),
.A2(n_21),
.B(n_23),
.C(n_34),
.Y(n_173)
);

O2A1O1Ixp33_ASAP7_75t_SL g244 ( 
.A1(n_173),
.A2(n_176),
.B(n_199),
.C(n_1),
.Y(n_244)
);

INVx8_ASAP7_75t_L g174 ( 
.A(n_105),
.Y(n_174)
);

INVx3_ASAP7_75t_L g220 ( 
.A(n_174),
.Y(n_220)
);

NAND2xp5_ASAP7_75t_SL g175 ( 
.A(n_125),
.B(n_83),
.Y(n_175)
);

A2O1A1Ixp33_ASAP7_75t_L g176 ( 
.A1(n_133),
.A2(n_67),
.B(n_25),
.C(n_46),
.Y(n_176)
);

OAI21xp33_ASAP7_75t_L g177 ( 
.A1(n_122),
.A2(n_39),
.B(n_25),
.Y(n_177)
);

CKINVDCx16_ASAP7_75t_R g230 ( 
.A(n_177),
.Y(n_230)
);

AOI22xp33_ASAP7_75t_L g178 ( 
.A1(n_148),
.A2(n_56),
.B1(n_39),
.B2(n_99),
.Y(n_178)
);

CKINVDCx20_ASAP7_75t_R g179 ( 
.A(n_107),
.Y(n_179)
);

OAI22xp5_ASAP7_75t_SL g180 ( 
.A1(n_143),
.A2(n_39),
.B1(n_67),
.B2(n_46),
.Y(n_180)
);

CKINVDCx20_ASAP7_75t_R g181 ( 
.A(n_107),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_SL g238 ( 
.A(n_181),
.B(n_201),
.Y(n_238)
);

CKINVDCx16_ASAP7_75t_R g182 ( 
.A(n_142),
.Y(n_182)
);

NOR2xp33_ASAP7_75t_L g227 ( 
.A(n_182),
.B(n_202),
.Y(n_227)
);

INVxp67_ASAP7_75t_L g231 ( 
.A(n_183),
.Y(n_231)
);

AOI22xp5_ASAP7_75t_SL g246 ( 
.A1(n_184),
.A2(n_134),
.B1(n_104),
.B2(n_152),
.Y(n_246)
);

HB1xp67_ASAP7_75t_L g185 ( 
.A(n_108),
.Y(n_185)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_185),
.Y(n_229)
);

AND2x2_ASAP7_75t_L g186 ( 
.A(n_114),
.B(n_25),
.Y(n_186)
);

FAx1_ASAP7_75t_SL g215 ( 
.A(n_186),
.B(n_195),
.CI(n_136),
.CON(n_215),
.SN(n_215)
);

INVx3_ASAP7_75t_L g188 ( 
.A(n_108),
.Y(n_188)
);

INVx3_ASAP7_75t_L g226 ( 
.A(n_188),
.Y(n_226)
);

BUFx2_ASAP7_75t_SL g189 ( 
.A(n_140),
.Y(n_189)
);

INVx2_ASAP7_75t_SL g236 ( 
.A(n_189),
.Y(n_236)
);

BUFx6f_ASAP7_75t_L g190 ( 
.A(n_111),
.Y(n_190)
);

INVx2_ASAP7_75t_L g221 ( 
.A(n_190),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_L g191 ( 
.A(n_118),
.B(n_46),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_L g245 ( 
.A(n_191),
.B(n_193),
.Y(n_245)
);

AOI22xp5_ASAP7_75t_SL g192 ( 
.A1(n_117),
.A2(n_25),
.B1(n_9),
.B2(n_10),
.Y(n_192)
);

XNOR2xp5_ASAP7_75t_L g248 ( 
.A(n_192),
.B(n_207),
.Y(n_248)
);

NAND2xp5_ASAP7_75t_L g193 ( 
.A(n_103),
.B(n_5),
.Y(n_193)
);

AND2x2_ASAP7_75t_L g195 ( 
.A(n_103),
.B(n_0),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_L g197 ( 
.A(n_124),
.B(n_5),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_L g252 ( 
.A(n_197),
.B(n_203),
.Y(n_252)
);

INVx11_ASAP7_75t_L g198 ( 
.A(n_140),
.Y(n_198)
);

INVx2_ASAP7_75t_L g223 ( 
.A(n_198),
.Y(n_223)
);

A2O1A1Ixp33_ASAP7_75t_L g199 ( 
.A1(n_116),
.A2(n_5),
.B(n_13),
.C(n_12),
.Y(n_199)
);

INVx11_ASAP7_75t_L g200 ( 
.A(n_152),
.Y(n_200)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_200),
.Y(n_237)
);

CKINVDCx14_ASAP7_75t_R g201 ( 
.A(n_145),
.Y(n_201)
);

CKINVDCx16_ASAP7_75t_R g202 ( 
.A(n_127),
.Y(n_202)
);

NAND2xp5_ASAP7_75t_SL g203 ( 
.A(n_130),
.B(n_4),
.Y(n_203)
);

OAI22xp5_ASAP7_75t_L g204 ( 
.A1(n_155),
.A2(n_4),
.B1(n_13),
.B2(n_11),
.Y(n_204)
);

AOI22xp5_ASAP7_75t_L g222 ( 
.A1(n_204),
.A2(n_208),
.B1(n_0),
.B2(n_1),
.Y(n_222)
);

NOR2xp33_ASAP7_75t_L g205 ( 
.A(n_136),
.B(n_3),
.Y(n_205)
);

NOR2xp33_ASAP7_75t_L g241 ( 
.A(n_205),
.B(n_1),
.Y(n_241)
);

AOI22xp33_ASAP7_75t_L g206 ( 
.A1(n_148),
.A2(n_3),
.B1(n_11),
.B2(n_13),
.Y(n_206)
);

OAI22xp5_ASAP7_75t_L g208 ( 
.A1(n_139),
.A2(n_15),
.B1(n_1),
.B2(n_2),
.Y(n_208)
);

INVx1_ASAP7_75t_SL g209 ( 
.A(n_129),
.Y(n_209)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_209),
.Y(n_249)
);

AND2x2_ASAP7_75t_L g265 ( 
.A(n_215),
.B(n_224),
.Y(n_265)
);

MAJIxp5_ASAP7_75t_L g217 ( 
.A(n_161),
.B(n_131),
.C(n_119),
.Y(n_217)
);

MAJIxp5_ASAP7_75t_L g255 ( 
.A(n_217),
.B(n_232),
.C(n_234),
.Y(n_255)
);

AOI22xp33_ASAP7_75t_L g218 ( 
.A1(n_168),
.A2(n_182),
.B1(n_161),
.B2(n_172),
.Y(n_218)
);

OAI22xp5_ASAP7_75t_SL g274 ( 
.A1(n_218),
.A2(n_175),
.B1(n_192),
.B2(n_191),
.Y(n_274)
);

OAI22xp5_ASAP7_75t_L g219 ( 
.A1(n_187),
.A2(n_120),
.B1(n_138),
.B2(n_132),
.Y(n_219)
);

AOI22xp5_ASAP7_75t_L g263 ( 
.A1(n_219),
.A2(n_239),
.B1(n_162),
.B2(n_164),
.Y(n_263)
);

OAI22xp5_ASAP7_75t_L g291 ( 
.A1(n_222),
.A2(n_246),
.B1(n_205),
.B2(n_209),
.Y(n_291)
);

CKINVDCx20_ASAP7_75t_R g225 ( 
.A(n_196),
.Y(n_225)
);

NOR2xp33_ASAP7_75t_L g257 ( 
.A(n_225),
.B(n_228),
.Y(n_257)
);

CKINVDCx20_ASAP7_75t_R g228 ( 
.A(n_196),
.Y(n_228)
);

MAJIxp5_ASAP7_75t_L g232 ( 
.A(n_176),
.B(n_112),
.C(n_119),
.Y(n_232)
);

XOR2xp5_ASAP7_75t_L g234 ( 
.A(n_160),
.B(n_146),
.Y(n_234)
);

OAI22xp5_ASAP7_75t_L g239 ( 
.A1(n_187),
.A2(n_120),
.B1(n_132),
.B2(n_151),
.Y(n_239)
);

MAJIxp5_ASAP7_75t_L g240 ( 
.A(n_176),
.B(n_134),
.C(n_135),
.Y(n_240)
);

MAJIxp5_ASAP7_75t_L g285 ( 
.A(n_240),
.B(n_186),
.C(n_195),
.Y(n_285)
);

NOR2xp33_ASAP7_75t_L g262 ( 
.A(n_241),
.B(n_243),
.Y(n_262)
);

AOI22xp33_ASAP7_75t_SL g242 ( 
.A1(n_172),
.A2(n_156),
.B1(n_135),
.B2(n_129),
.Y(n_242)
);

INVxp67_ASAP7_75t_L g276 ( 
.A(n_242),
.Y(n_276)
);

CKINVDCx20_ASAP7_75t_R g243 ( 
.A(n_194),
.Y(n_243)
);

OAI21xp5_ASAP7_75t_SL g288 ( 
.A1(n_244),
.A2(n_250),
.B(n_199),
.Y(n_288)
);

NOR2xp33_ASAP7_75t_L g247 ( 
.A(n_159),
.B(n_104),
.Y(n_247)
);

NOR2xp33_ASAP7_75t_L g269 ( 
.A(n_247),
.B(n_201),
.Y(n_269)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_165),
.Y(n_251)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_251),
.Y(n_256)
);

INVx2_ASAP7_75t_SL g253 ( 
.A(n_220),
.Y(n_253)
);

INVx2_ASAP7_75t_SL g314 ( 
.A(n_253),
.Y(n_314)
);

AOI22xp5_ASAP7_75t_SL g254 ( 
.A1(n_230),
.A2(n_231),
.B1(n_219),
.B2(n_216),
.Y(n_254)
);

INVxp67_ASAP7_75t_L g302 ( 
.A(n_254),
.Y(n_302)
);

AOI22xp33_ASAP7_75t_L g258 ( 
.A1(n_227),
.A2(n_216),
.B1(n_224),
.B2(n_210),
.Y(n_258)
);

AOI22xp33_ASAP7_75t_L g307 ( 
.A1(n_258),
.A2(n_208),
.B1(n_249),
.B2(n_202),
.Y(n_307)
);

INVx3_ASAP7_75t_L g259 ( 
.A(n_226),
.Y(n_259)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_259),
.Y(n_292)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_211),
.Y(n_260)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_260),
.Y(n_293)
);

NAND2xp5_ASAP7_75t_L g261 ( 
.A(n_252),
.B(n_203),
.Y(n_261)
);

NAND2xp5_ASAP7_75t_L g312 ( 
.A(n_261),
.B(n_264),
.Y(n_312)
);

OAI22xp5_ASAP7_75t_L g297 ( 
.A1(n_263),
.A2(n_266),
.B1(n_287),
.B2(n_246),
.Y(n_297)
);

NAND2xp5_ASAP7_75t_L g264 ( 
.A(n_252),
.B(n_193),
.Y(n_264)
);

AOI22xp5_ASAP7_75t_L g266 ( 
.A1(n_234),
.A2(n_204),
.B1(n_180),
.B2(n_169),
.Y(n_266)
);

BUFx6f_ASAP7_75t_L g267 ( 
.A(n_221),
.Y(n_267)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_267),
.Y(n_296)
);

OAI21xp5_ASAP7_75t_L g268 ( 
.A1(n_233),
.A2(n_183),
.B(n_207),
.Y(n_268)
);

OAI21xp5_ASAP7_75t_L g327 ( 
.A1(n_268),
.A2(n_185),
.B(n_213),
.Y(n_327)
);

NOR2xp33_ASAP7_75t_L g313 ( 
.A(n_269),
.B(n_270),
.Y(n_313)
);

CKINVDCx16_ASAP7_75t_R g270 ( 
.A(n_238),
.Y(n_270)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_211),
.Y(n_271)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_271),
.Y(n_299)
);

XNOR2xp5_ASAP7_75t_SL g272 ( 
.A(n_245),
.B(n_170),
.Y(n_272)
);

XOR2xp5_ASAP7_75t_L g301 ( 
.A(n_272),
.B(n_285),
.Y(n_301)
);

INVx2_ASAP7_75t_L g273 ( 
.A(n_213),
.Y(n_273)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_273),
.Y(n_300)
);

AOI22xp5_ASAP7_75t_L g294 ( 
.A1(n_274),
.A2(n_286),
.B1(n_291),
.B2(n_265),
.Y(n_294)
);

INVx3_ASAP7_75t_L g275 ( 
.A(n_226),
.Y(n_275)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_275),
.Y(n_306)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_251),
.Y(n_277)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_277),
.Y(n_319)
);

NAND2xp5_ASAP7_75t_L g278 ( 
.A(n_245),
.B(n_197),
.Y(n_278)
);

NAND2xp5_ASAP7_75t_L g326 ( 
.A(n_278),
.B(n_279),
.Y(n_326)
);

INVx2_ASAP7_75t_SL g279 ( 
.A(n_220),
.Y(n_279)
);

NOR2xp33_ASAP7_75t_SL g280 ( 
.A(n_225),
.B(n_170),
.Y(n_280)
);

NAND2xp5_ASAP7_75t_SL g315 ( 
.A(n_280),
.B(n_282),
.Y(n_315)
);

NOR2xp33_ASAP7_75t_L g281 ( 
.A(n_243),
.B(n_163),
.Y(n_281)
);

NOR2xp33_ASAP7_75t_L g295 ( 
.A(n_281),
.B(n_283),
.Y(n_295)
);

NOR2xp33_ASAP7_75t_SL g282 ( 
.A(n_228),
.B(n_166),
.Y(n_282)
);

NAND2xp5_ASAP7_75t_SL g283 ( 
.A(n_233),
.B(n_173),
.Y(n_283)
);

XNOR2xp5_ASAP7_75t_L g284 ( 
.A(n_232),
.B(n_173),
.Y(n_284)
);

MAJIxp5_ASAP7_75t_L g303 ( 
.A(n_284),
.B(n_217),
.C(n_215),
.Y(n_303)
);

OAI22xp5_ASAP7_75t_SL g286 ( 
.A1(n_210),
.A2(n_183),
.B1(n_167),
.B2(n_195),
.Y(n_286)
);

AOI22xp5_ASAP7_75t_L g287 ( 
.A1(n_231),
.A2(n_248),
.B1(n_244),
.B2(n_250),
.Y(n_287)
);

AOI21xp5_ASAP7_75t_L g316 ( 
.A1(n_288),
.A2(n_199),
.B(n_236),
.Y(n_316)
);

NOR2xp33_ASAP7_75t_L g289 ( 
.A(n_212),
.B(n_235),
.Y(n_289)
);

CKINVDCx20_ASAP7_75t_R g310 ( 
.A(n_289),
.Y(n_310)
);

XNOR2xp5_ASAP7_75t_SL g290 ( 
.A(n_248),
.B(n_195),
.Y(n_290)
);

XOR2xp5_ASAP7_75t_L g305 ( 
.A(n_290),
.B(n_186),
.Y(n_305)
);

OAI22xp5_ASAP7_75t_SL g352 ( 
.A1(n_294),
.A2(n_307),
.B1(n_263),
.B2(n_253),
.Y(n_352)
);

NAND2xp5_ASAP7_75t_L g342 ( 
.A(n_297),
.B(n_323),
.Y(n_342)
);

OAI32xp33_ASAP7_75t_L g298 ( 
.A1(n_283),
.A2(n_244),
.A3(n_240),
.B1(n_194),
.B2(n_215),
.Y(n_298)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_298),
.Y(n_332)
);

MAJIxp5_ASAP7_75t_L g330 ( 
.A(n_303),
.B(n_304),
.C(n_255),
.Y(n_330)
);

MAJIxp5_ASAP7_75t_L g304 ( 
.A(n_255),
.B(n_290),
.C(n_272),
.Y(n_304)
);

XNOR2xp5_ASAP7_75t_L g333 ( 
.A(n_305),
.B(n_285),
.Y(n_333)
);

OA21x2_ASAP7_75t_L g308 ( 
.A1(n_288),
.A2(n_249),
.B(n_222),
.Y(n_308)
);

CKINVDCx20_ASAP7_75t_R g331 ( 
.A(n_308),
.Y(n_331)
);

BUFx24_ASAP7_75t_SL g309 ( 
.A(n_282),
.Y(n_309)
);

NOR2xp33_ASAP7_75t_L g338 ( 
.A(n_309),
.B(n_320),
.Y(n_338)
);

AOI22xp33_ASAP7_75t_SL g311 ( 
.A1(n_276),
.A2(n_236),
.B1(n_223),
.B2(n_229),
.Y(n_311)
);

INVxp67_ASAP7_75t_L g329 ( 
.A(n_311),
.Y(n_329)
);

OAI21xp5_ASAP7_75t_SL g350 ( 
.A1(n_316),
.A2(n_321),
.B(n_279),
.Y(n_350)
);

CKINVDCx20_ASAP7_75t_R g317 ( 
.A(n_257),
.Y(n_317)
);

NOR2xp33_ASAP7_75t_L g356 ( 
.A(n_317),
.B(n_322),
.Y(n_356)
);

NOR2xp67_ASAP7_75t_SL g318 ( 
.A(n_268),
.B(n_284),
.Y(n_318)
);

OAI21xp5_ASAP7_75t_L g354 ( 
.A1(n_318),
.A2(n_327),
.B(n_256),
.Y(n_354)
);

BUFx24_ASAP7_75t_SL g320 ( 
.A(n_280),
.Y(n_320)
);

AOI21xp5_ASAP7_75t_L g321 ( 
.A1(n_276),
.A2(n_236),
.B(n_237),
.Y(n_321)
);

CKINVDCx20_ASAP7_75t_R g322 ( 
.A(n_262),
.Y(n_322)
);

O2A1O1Ixp33_ASAP7_75t_L g323 ( 
.A1(n_287),
.A2(n_181),
.B(n_179),
.C(n_237),
.Y(n_323)
);

OAI21xp5_ASAP7_75t_SL g324 ( 
.A1(n_265),
.A2(n_229),
.B(n_209),
.Y(n_324)
);

AOI21xp5_ASAP7_75t_L g349 ( 
.A1(n_324),
.A2(n_274),
.B(n_253),
.Y(n_349)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_260),
.Y(n_325)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_325),
.Y(n_334)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_271),
.Y(n_328)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_328),
.Y(n_336)
);

MAJIxp5_ASAP7_75t_L g368 ( 
.A(n_330),
.B(n_346),
.C(n_355),
.Y(n_368)
);

XNOR2xp5_ASAP7_75t_SL g383 ( 
.A(n_333),
.B(n_308),
.Y(n_383)
);

HB1xp67_ASAP7_75t_L g335 ( 
.A(n_292),
.Y(n_335)
);

INVx1_ASAP7_75t_L g371 ( 
.A(n_335),
.Y(n_371)
);

CKINVDCx16_ASAP7_75t_R g337 ( 
.A(n_313),
.Y(n_337)
);

NAND2xp5_ASAP7_75t_SL g370 ( 
.A(n_337),
.B(n_348),
.Y(n_370)
);

NOR2xp33_ASAP7_75t_L g339 ( 
.A(n_310),
.B(n_270),
.Y(n_339)
);

CKINVDCx14_ASAP7_75t_R g385 ( 
.A(n_339),
.Y(n_385)
);

CKINVDCx20_ASAP7_75t_R g340 ( 
.A(n_315),
.Y(n_340)
);

CKINVDCx20_ASAP7_75t_R g363 ( 
.A(n_340),
.Y(n_363)
);

OAI22xp33_ASAP7_75t_SL g341 ( 
.A1(n_302),
.A2(n_291),
.B1(n_266),
.B2(n_254),
.Y(n_341)
);

AOI22xp5_ASAP7_75t_L g367 ( 
.A1(n_341),
.A2(n_352),
.B1(n_297),
.B2(n_321),
.Y(n_367)
);

NAND2xp5_ASAP7_75t_L g343 ( 
.A(n_315),
.B(n_278),
.Y(n_343)
);

INVx1_ASAP7_75t_L g365 ( 
.A(n_343),
.Y(n_365)
);

XNOR2xp5_ASAP7_75t_L g344 ( 
.A(n_301),
.B(n_264),
.Y(n_344)
);

XNOR2xp5_ASAP7_75t_L g369 ( 
.A(n_344),
.B(n_345),
.Y(n_369)
);

XNOR2xp5_ASAP7_75t_L g345 ( 
.A(n_301),
.B(n_261),
.Y(n_345)
);

XOR2xp5_ASAP7_75t_L g346 ( 
.A(n_304),
.B(n_286),
.Y(n_346)
);

NAND2xp5_ASAP7_75t_L g347 ( 
.A(n_326),
.B(n_265),
.Y(n_347)
);

INVx1_ASAP7_75t_L g377 ( 
.A(n_347),
.Y(n_377)
);

NOR2xp33_ASAP7_75t_L g348 ( 
.A(n_310),
.B(n_317),
.Y(n_348)
);

OAI21xp5_ASAP7_75t_SL g381 ( 
.A1(n_349),
.A2(n_323),
.B(n_324),
.Y(n_381)
);

AOI21xp5_ASAP7_75t_L g364 ( 
.A1(n_350),
.A2(n_354),
.B(n_327),
.Y(n_364)
);

NOR2xp33_ASAP7_75t_L g351 ( 
.A(n_295),
.B(n_275),
.Y(n_351)
);

NAND2xp5_ASAP7_75t_SL g389 ( 
.A(n_351),
.B(n_306),
.Y(n_389)
);

NAND2xp5_ASAP7_75t_L g353 ( 
.A(n_326),
.B(n_277),
.Y(n_353)
);

INVx1_ASAP7_75t_L g390 ( 
.A(n_353),
.Y(n_390)
);

MAJIxp5_ASAP7_75t_L g355 ( 
.A(n_303),
.B(n_256),
.C(n_259),
.Y(n_355)
);

NAND2xp5_ASAP7_75t_L g357 ( 
.A(n_312),
.B(n_279),
.Y(n_357)
);

NAND2xp5_ASAP7_75t_L g373 ( 
.A(n_357),
.B(n_358),
.Y(n_373)
);

NAND2xp5_ASAP7_75t_L g358 ( 
.A(n_312),
.B(n_273),
.Y(n_358)
);

INVx1_ASAP7_75t_L g359 ( 
.A(n_293),
.Y(n_359)
);

CKINVDCx16_ASAP7_75t_R g362 ( 
.A(n_359),
.Y(n_362)
);

XNOR2xp5_ASAP7_75t_L g360 ( 
.A(n_305),
.B(n_189),
.Y(n_360)
);

XNOR2xp5_ASAP7_75t_L g372 ( 
.A(n_360),
.B(n_298),
.Y(n_372)
);

INVx2_ASAP7_75t_L g361 ( 
.A(n_296),
.Y(n_361)
);

NAND2xp5_ASAP7_75t_L g380 ( 
.A(n_361),
.B(n_296),
.Y(n_380)
);

CKINVDCx14_ASAP7_75t_R g417 ( 
.A(n_364),
.Y(n_417)
);

XOR2xp5_ASAP7_75t_L g366 ( 
.A(n_346),
.B(n_318),
.Y(n_366)
);

XOR2xp5_ASAP7_75t_L g392 ( 
.A(n_366),
.B(n_372),
.Y(n_392)
);

OAI22xp5_ASAP7_75t_L g393 ( 
.A1(n_367),
.A2(n_375),
.B1(n_387),
.B2(n_342),
.Y(n_393)
);

XNOR2xp5_ASAP7_75t_L g374 ( 
.A(n_344),
.B(n_294),
.Y(n_374)
);

XNOR2xp5_ASAP7_75t_L g399 ( 
.A(n_374),
.B(n_379),
.Y(n_399)
);

OAI22xp5_ASAP7_75t_L g375 ( 
.A1(n_340),
.A2(n_322),
.B1(n_313),
.B2(n_316),
.Y(n_375)
);

NOR2xp33_ASAP7_75t_SL g376 ( 
.A(n_356),
.B(n_293),
.Y(n_376)
);

NAND2xp5_ASAP7_75t_SL g397 ( 
.A(n_376),
.B(n_378),
.Y(n_397)
);

NOR2xp33_ASAP7_75t_SL g378 ( 
.A(n_356),
.B(n_338),
.Y(n_378)
);

XNOR2xp5_ASAP7_75t_L g379 ( 
.A(n_330),
.B(n_308),
.Y(n_379)
);

NAND2xp5_ASAP7_75t_L g402 ( 
.A(n_380),
.B(n_388),
.Y(n_402)
);

INVx1_ASAP7_75t_L g395 ( 
.A(n_381),
.Y(n_395)
);

AOI22xp5_ASAP7_75t_L g382 ( 
.A1(n_352),
.A2(n_308),
.B1(n_323),
.B2(n_325),
.Y(n_382)
);

OAI22xp5_ASAP7_75t_SL g396 ( 
.A1(n_382),
.A2(n_386),
.B1(n_391),
.B2(n_354),
.Y(n_396)
);

XOR2xp5_ASAP7_75t_L g398 ( 
.A(n_383),
.B(n_384),
.Y(n_398)
);

XOR2xp5_ASAP7_75t_L g384 ( 
.A(n_333),
.B(n_328),
.Y(n_384)
);

AOI22xp5_ASAP7_75t_L g386 ( 
.A1(n_331),
.A2(n_299),
.B1(n_319),
.B2(n_314),
.Y(n_386)
);

OAI22xp5_ASAP7_75t_L g387 ( 
.A1(n_337),
.A2(n_299),
.B1(n_319),
.B2(n_314),
.Y(n_387)
);

OA21x2_ASAP7_75t_L g388 ( 
.A1(n_342),
.A2(n_306),
.B(n_292),
.Y(n_388)
);

NAND2xp5_ASAP7_75t_SL g404 ( 
.A(n_389),
.B(n_385),
.Y(n_404)
);

AOI22xp5_ASAP7_75t_L g391 ( 
.A1(n_331),
.A2(n_332),
.B1(n_349),
.B2(n_329),
.Y(n_391)
);

AOI22xp5_ASAP7_75t_SL g432 ( 
.A1(n_393),
.A2(n_396),
.B1(n_221),
.B2(n_174),
.Y(n_432)
);

FAx1_ASAP7_75t_SL g394 ( 
.A(n_383),
.B(n_347),
.CI(n_343),
.CON(n_394),
.SN(n_394)
);

NAND2xp5_ASAP7_75t_L g429 ( 
.A(n_394),
.B(n_405),
.Y(n_429)
);

XOR2xp5_ASAP7_75t_L g400 ( 
.A(n_366),
.B(n_369),
.Y(n_400)
);

XOR2xp5_ASAP7_75t_L g421 ( 
.A(n_400),
.B(n_410),
.Y(n_421)
);

INVx1_ASAP7_75t_L g401 ( 
.A(n_373),
.Y(n_401)
);

INVx1_ASAP7_75t_L g422 ( 
.A(n_401),
.Y(n_422)
);

NAND2xp5_ASAP7_75t_L g403 ( 
.A(n_363),
.B(n_353),
.Y(n_403)
);

INVx1_ASAP7_75t_L g436 ( 
.A(n_403),
.Y(n_436)
);

CKINVDCx14_ASAP7_75t_R g428 ( 
.A(n_404),
.Y(n_428)
);

INVx1_ASAP7_75t_L g405 ( 
.A(n_373),
.Y(n_405)
);

MAJIxp5_ASAP7_75t_L g406 ( 
.A(n_368),
.B(n_355),
.C(n_345),
.Y(n_406)
);

MAJIxp5_ASAP7_75t_L g423 ( 
.A(n_406),
.B(n_407),
.C(n_369),
.Y(n_423)
);

MAJIxp5_ASAP7_75t_L g407 ( 
.A(n_368),
.B(n_332),
.C(n_360),
.Y(n_407)
);

NAND2xp5_ASAP7_75t_L g408 ( 
.A(n_370),
.B(n_357),
.Y(n_408)
);

INVx2_ASAP7_75t_L g433 ( 
.A(n_408),
.Y(n_433)
);

OAI21xp33_ASAP7_75t_L g409 ( 
.A1(n_377),
.A2(n_358),
.B(n_350),
.Y(n_409)
);

AOI321xp33_ASAP7_75t_L g425 ( 
.A1(n_409),
.A2(n_381),
.A3(n_388),
.B1(n_362),
.B2(n_380),
.C(n_371),
.Y(n_425)
);

NAND2xp5_ASAP7_75t_L g410 ( 
.A(n_365),
.B(n_359),
.Y(n_410)
);

NOR2xp33_ASAP7_75t_SL g411 ( 
.A(n_365),
.B(n_336),
.Y(n_411)
);

OR2x2_ASAP7_75t_L g435 ( 
.A(n_411),
.B(n_412),
.Y(n_435)
);

INVx1_ASAP7_75t_L g412 ( 
.A(n_390),
.Y(n_412)
);

INVx1_ASAP7_75t_L g413 ( 
.A(n_390),
.Y(n_413)
);

AOI22xp33_ASAP7_75t_SL g419 ( 
.A1(n_413),
.A2(n_414),
.B1(n_361),
.B2(n_334),
.Y(n_419)
);

INVx1_ASAP7_75t_L g414 ( 
.A(n_377),
.Y(n_414)
);

NAND2xp5_ASAP7_75t_SL g415 ( 
.A(n_379),
.B(n_336),
.Y(n_415)
);

OAI22xp5_ASAP7_75t_L g424 ( 
.A1(n_415),
.A2(n_374),
.B1(n_386),
.B2(n_384),
.Y(n_424)
);

MAJx2_ASAP7_75t_L g416 ( 
.A(n_372),
.B(n_334),
.C(n_329),
.Y(n_416)
);

XOR2xp5_ASAP7_75t_L g427 ( 
.A(n_416),
.B(n_392),
.Y(n_427)
);

NOR2xp67_ASAP7_75t_SL g418 ( 
.A(n_417),
.B(n_364),
.Y(n_418)
);

OAI21xp5_ASAP7_75t_L g445 ( 
.A1(n_418),
.A2(n_426),
.B(n_431),
.Y(n_445)
);

INVx1_ASAP7_75t_L g439 ( 
.A(n_419),
.Y(n_439)
);

OAI22xp5_ASAP7_75t_SL g420 ( 
.A1(n_402),
.A2(n_367),
.B1(n_382),
.B2(n_391),
.Y(n_420)
);

AOI22xp5_ASAP7_75t_L g441 ( 
.A1(n_420),
.A2(n_438),
.B1(n_413),
.B2(n_405),
.Y(n_441)
);

XNOR2xp5_ASAP7_75t_L g442 ( 
.A(n_423),
.B(n_424),
.Y(n_442)
);

AOI21x1_ASAP7_75t_SL g443 ( 
.A1(n_425),
.A2(n_416),
.B(n_394),
.Y(n_443)
);

AOI21xp5_ASAP7_75t_L g426 ( 
.A1(n_395),
.A2(n_396),
.B(n_402),
.Y(n_426)
);

NOR2xp33_ASAP7_75t_L g448 ( 
.A(n_427),
.B(n_399),
.Y(n_448)
);

A2O1A1Ixp33_ASAP7_75t_L g430 ( 
.A1(n_395),
.A2(n_388),
.B(n_300),
.C(n_314),
.Y(n_430)
);

INVx1_ASAP7_75t_L g446 ( 
.A(n_430),
.Y(n_446)
);

AOI21xp5_ASAP7_75t_L g431 ( 
.A1(n_403),
.A2(n_300),
.B(n_223),
.Y(n_431)
);

OAI22xp5_ASAP7_75t_SL g444 ( 
.A1(n_432),
.A2(n_401),
.B1(n_414),
.B2(n_408),
.Y(n_444)
);

MAJIxp5_ASAP7_75t_L g434 ( 
.A(n_406),
.B(n_267),
.C(n_188),
.Y(n_434)
);

MAJIxp5_ASAP7_75t_L g449 ( 
.A(n_434),
.B(n_421),
.C(n_423),
.Y(n_449)
);

OAI22xp5_ASAP7_75t_L g437 ( 
.A1(n_397),
.A2(n_267),
.B1(n_214),
.B2(n_190),
.Y(n_437)
);

INVx1_ASAP7_75t_L g447 ( 
.A(n_437),
.Y(n_447)
);

OAI22xp5_ASAP7_75t_L g438 ( 
.A1(n_412),
.A2(n_214),
.B1(n_171),
.B2(n_190),
.Y(n_438)
);

NAND2xp5_ASAP7_75t_L g440 ( 
.A(n_435),
.B(n_411),
.Y(n_440)
);

INVx1_ASAP7_75t_L g456 ( 
.A(n_440),
.Y(n_456)
);

OAI22xp5_ASAP7_75t_L g461 ( 
.A1(n_441),
.A2(n_429),
.B1(n_433),
.B2(n_430),
.Y(n_461)
);

INVx1_ASAP7_75t_L g457 ( 
.A(n_443),
.Y(n_457)
);

AOI22xp5_ASAP7_75t_L g458 ( 
.A1(n_444),
.A2(n_420),
.B1(n_436),
.B2(n_431),
.Y(n_458)
);

XOR2xp5_ASAP7_75t_L g465 ( 
.A(n_448),
.B(n_398),
.Y(n_465)
);

MAJIxp5_ASAP7_75t_L g466 ( 
.A(n_449),
.B(n_451),
.C(n_398),
.Y(n_466)
);

NAND2xp5_ASAP7_75t_SL g450 ( 
.A(n_428),
.B(n_407),
.Y(n_450)
);

NAND2xp5_ASAP7_75t_SL g467 ( 
.A(n_450),
.B(n_452),
.Y(n_467)
);

MAJIxp5_ASAP7_75t_L g451 ( 
.A(n_434),
.B(n_399),
.C(n_400),
.Y(n_451)
);

NOR2xp33_ASAP7_75t_L g452 ( 
.A(n_435),
.B(n_394),
.Y(n_452)
);

NOR2xp33_ASAP7_75t_L g453 ( 
.A(n_426),
.B(n_410),
.Y(n_453)
);

CKINVDCx16_ASAP7_75t_R g463 ( 
.A(n_453),
.Y(n_463)
);

INVxp67_ASAP7_75t_L g454 ( 
.A(n_418),
.Y(n_454)
);

NOR2xp33_ASAP7_75t_L g462 ( 
.A(n_454),
.B(n_429),
.Y(n_462)
);

NAND2xp5_ASAP7_75t_L g455 ( 
.A(n_436),
.B(n_392),
.Y(n_455)
);

INVx1_ASAP7_75t_L g469 ( 
.A(n_455),
.Y(n_469)
);

NAND2xp5_ASAP7_75t_L g476 ( 
.A(n_458),
.B(n_461),
.Y(n_476)
);

AOI21xp5_ASAP7_75t_L g459 ( 
.A1(n_454),
.A2(n_422),
.B(n_425),
.Y(n_459)
);

AOI21xp5_ASAP7_75t_L g482 ( 
.A1(n_459),
.A2(n_468),
.B(n_470),
.Y(n_482)
);

AOI22xp5_ASAP7_75t_L g460 ( 
.A1(n_447),
.A2(n_422),
.B1(n_433),
.B2(n_432),
.Y(n_460)
);

INVx1_ASAP7_75t_L g474 ( 
.A(n_460),
.Y(n_474)
);

OR2x2_ASAP7_75t_L g481 ( 
.A(n_462),
.B(n_445),
.Y(n_481)
);

OAI22xp5_ASAP7_75t_L g464 ( 
.A1(n_446),
.A2(n_438),
.B1(n_421),
.B2(n_427),
.Y(n_464)
);

NAND2xp5_ASAP7_75t_L g477 ( 
.A(n_464),
.B(n_465),
.Y(n_477)
);

NAND2xp5_ASAP7_75t_L g479 ( 
.A(n_466),
.B(n_451),
.Y(n_479)
);

OAI21xp5_ASAP7_75t_SL g468 ( 
.A1(n_440),
.A2(n_198),
.B(n_174),
.Y(n_468)
);

OAI21xp5_ASAP7_75t_SL g470 ( 
.A1(n_439),
.A2(n_198),
.B(n_171),
.Y(n_470)
);

INVxp33_ASAP7_75t_L g471 ( 
.A(n_467),
.Y(n_471)
);

INVx1_ASAP7_75t_L g484 ( 
.A(n_471),
.Y(n_484)
);

NAND2xp5_ASAP7_75t_L g472 ( 
.A(n_456),
.B(n_444),
.Y(n_472)
);

NAND2xp5_ASAP7_75t_L g487 ( 
.A(n_472),
.B(n_473),
.Y(n_487)
);

NOR2xp33_ASAP7_75t_SL g473 ( 
.A(n_457),
.B(n_442),
.Y(n_473)
);

OAI21xp5_ASAP7_75t_SL g475 ( 
.A1(n_459),
.A2(n_443),
.B(n_445),
.Y(n_475)
);

AOI21xp5_ASAP7_75t_L g492 ( 
.A1(n_475),
.A2(n_458),
.B(n_469),
.Y(n_492)
);

CKINVDCx16_ASAP7_75t_R g478 ( 
.A(n_456),
.Y(n_478)
);

BUFx2_ASAP7_75t_L g485 ( 
.A(n_478),
.Y(n_485)
);

XNOR2xp5_ASAP7_75t_L g491 ( 
.A(n_479),
.B(n_480),
.Y(n_491)
);

NAND2xp5_ASAP7_75t_L g480 ( 
.A(n_463),
.B(n_441),
.Y(n_480)
);

INVxp67_ASAP7_75t_L g489 ( 
.A(n_481),
.Y(n_489)
);

MAJIxp5_ASAP7_75t_L g483 ( 
.A(n_466),
.B(n_449),
.C(n_442),
.Y(n_483)
);

XNOR2xp5_ASAP7_75t_L g493 ( 
.A(n_483),
.B(n_465),
.Y(n_493)
);

OAI21xp5_ASAP7_75t_SL g486 ( 
.A1(n_483),
.A2(n_457),
.B(n_481),
.Y(n_486)
);

AO21x1_ASAP7_75t_L g496 ( 
.A1(n_486),
.A2(n_490),
.B(n_468),
.Y(n_496)
);

A2O1A1Ixp33_ASAP7_75t_L g488 ( 
.A1(n_475),
.A2(n_472),
.B(n_476),
.C(n_471),
.Y(n_488)
);

INVx1_ASAP7_75t_L g497 ( 
.A(n_488),
.Y(n_497)
);

AND2x2_ASAP7_75t_L g490 ( 
.A(n_477),
.B(n_469),
.Y(n_490)
);

OA21x2_ASAP7_75t_L g495 ( 
.A1(n_492),
.A2(n_482),
.B(n_474),
.Y(n_495)
);

NAND2xp5_ASAP7_75t_L g498 ( 
.A(n_493),
.B(n_455),
.Y(n_498)
);

AOI21xp5_ASAP7_75t_L g494 ( 
.A1(n_489),
.A2(n_484),
.B(n_491),
.Y(n_494)
);

OAI21xp5_ASAP7_75t_L g500 ( 
.A1(n_494),
.A2(n_495),
.B(n_489),
.Y(n_500)
);

AOI21xp5_ASAP7_75t_L g501 ( 
.A1(n_496),
.A2(n_490),
.B(n_487),
.Y(n_501)
);

NAND2xp5_ASAP7_75t_SL g502 ( 
.A(n_498),
.B(n_499),
.Y(n_502)
);

NOR2xp33_ASAP7_75t_L g499 ( 
.A(n_485),
.B(n_460),
.Y(n_499)
);

AO21x1_ASAP7_75t_L g504 ( 
.A1(n_500),
.A2(n_501),
.B(n_470),
.Y(n_504)
);

NOR3xp33_ASAP7_75t_L g503 ( 
.A(n_502),
.B(n_497),
.C(n_485),
.Y(n_503)
);

AOI22xp5_ASAP7_75t_SL g505 ( 
.A1(n_503),
.A2(n_504),
.B1(n_482),
.B2(n_200),
.Y(n_505)
);

OAI21xp5_ASAP7_75t_L g506 ( 
.A1(n_505),
.A2(n_200),
.B(n_2),
.Y(n_506)
);

MAJIxp5_ASAP7_75t_L g507 ( 
.A(n_506),
.B(n_2),
.C(n_489),
.Y(n_507)
);


endmodule