module fake_jpeg_18642_n_71 (n_3, n_2, n_1, n_0, n_4, n_8, n_9, n_6, n_5, n_7, n_71);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_71;

wire n_13;
wire n_21;
wire n_57;
wire n_53;
wire n_33;
wire n_54;
wire n_61;
wire n_45;
wire n_23;
wire n_10;
wire n_69;
wire n_27;
wire n_55;
wire n_64;
wire n_22;
wire n_47;
wire n_51;
wire n_14;
wire n_40;
wire n_19;
wire n_20;
wire n_18;
wire n_59;
wire n_35;
wire n_48;
wire n_68;
wire n_52;
wire n_46;
wire n_58;
wire n_41;
wire n_60;
wire n_63;
wire n_65;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_16;
wire n_49;
wire n_24;
wire n_28;
wire n_38;
wire n_26;
wire n_44;
wire n_36;
wire n_11;
wire n_62;
wire n_25;
wire n_17;
wire n_31;
wire n_56;
wire n_67;
wire n_29;
wire n_37;
wire n_43;
wire n_50;
wire n_12;
wire n_32;
wire n_70;
wire n_15;
wire n_66;

INVx6_ASAP7_75t_L g10 ( 
.A(n_0),
.Y(n_10)
);

AOI21xp5_ASAP7_75t_L g11 ( 
.A1(n_0),
.A2(n_3),
.B(n_5),
.Y(n_11)
);

INVx4_ASAP7_75t_L g12 ( 
.A(n_3),
.Y(n_12)
);

BUFx4f_ASAP7_75t_L g13 ( 
.A(n_6),
.Y(n_13)
);

INVx6_ASAP7_75t_L g14 ( 
.A(n_6),
.Y(n_14)
);

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_7),
.Y(n_15)
);

INVx6_ASAP7_75t_L g16 ( 
.A(n_4),
.Y(n_16)
);

INVx5_ASAP7_75t_L g17 ( 
.A(n_0),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_5),
.Y(n_18)
);

BUFx5_ASAP7_75t_L g19 ( 
.A(n_9),
.Y(n_19)
);

INVx2_ASAP7_75t_L g20 ( 
.A(n_1),
.Y(n_20)
);

NAND2xp5_ASAP7_75t_L g21 ( 
.A(n_20),
.B(n_1),
.Y(n_21)
);

NAND2xp5_ASAP7_75t_L g33 ( 
.A(n_21),
.B(n_28),
.Y(n_33)
);

INVx6_ASAP7_75t_L g22 ( 
.A(n_20),
.Y(n_22)
);

INVx11_ASAP7_75t_L g32 ( 
.A(n_22),
.Y(n_32)
);

OAI22xp5_ASAP7_75t_L g23 ( 
.A1(n_11),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_23)
);

AOI22xp5_ASAP7_75t_L g37 ( 
.A1(n_23),
.A2(n_26),
.B1(n_27),
.B2(n_7),
.Y(n_37)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_18),
.Y(n_24)
);

INVx1_ASAP7_75t_SL g31 ( 
.A(n_24),
.Y(n_31)
);

INVxp33_ASAP7_75t_L g25 ( 
.A(n_19),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_25),
.Y(n_35)
);

OAI22xp33_ASAP7_75t_L g26 ( 
.A1(n_14),
.A2(n_2),
.B1(n_4),
.B2(n_5),
.Y(n_26)
);

OA22x2_ASAP7_75t_SL g27 ( 
.A1(n_11),
.A2(n_2),
.B1(n_4),
.B2(n_6),
.Y(n_27)
);

NOR2xp33_ASAP7_75t_L g28 ( 
.A(n_15),
.B(n_7),
.Y(n_28)
);

OAI22xp5_ASAP7_75t_SL g29 ( 
.A1(n_22),
.A2(n_14),
.B1(n_16),
.B2(n_10),
.Y(n_29)
);

AOI22xp5_ASAP7_75t_L g44 ( 
.A1(n_29),
.A2(n_36),
.B1(n_34),
.B2(n_35),
.Y(n_44)
);

AOI22xp33_ASAP7_75t_SL g30 ( 
.A1(n_22),
.A2(n_14),
.B1(n_10),
.B2(n_16),
.Y(n_30)
);

OAI22xp5_ASAP7_75t_SL g46 ( 
.A1(n_30),
.A2(n_37),
.B1(n_18),
.B2(n_28),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_L g34 ( 
.A(n_21),
.B(n_27),
.Y(n_34)
);

NAND2xp5_ASAP7_75t_L g43 ( 
.A(n_34),
.B(n_13),
.Y(n_43)
);

OAI22xp5_ASAP7_75t_SL g36 ( 
.A1(n_27),
.A2(n_12),
.B1(n_17),
.B2(n_15),
.Y(n_36)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_29),
.Y(n_38)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_38),
.Y(n_53)
);

AOI22xp5_ASAP7_75t_SL g39 ( 
.A1(n_36),
.A2(n_27),
.B1(n_17),
.B2(n_12),
.Y(n_39)
);

XNOR2xp5_ASAP7_75t_L g52 ( 
.A(n_39),
.B(n_40),
.Y(n_52)
);

XNOR2xp5_ASAP7_75t_L g40 ( 
.A(n_33),
.B(n_23),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_31),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g49 ( 
.A(n_41),
.B(n_44),
.Y(n_49)
);

INVxp67_ASAP7_75t_L g42 ( 
.A(n_30),
.Y(n_42)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_42),
.Y(n_48)
);

XNOR2xp5_ASAP7_75t_L g54 ( 
.A(n_43),
.B(n_45),
.Y(n_54)
);

XNOR2xp5_ASAP7_75t_L g45 ( 
.A(n_33),
.B(n_24),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g51 ( 
.A(n_46),
.B(n_47),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g47 ( 
.A(n_35),
.B(n_8),
.Y(n_47)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_44),
.Y(n_50)
);

OAI22xp5_ASAP7_75t_L g59 ( 
.A1(n_50),
.A2(n_31),
.B1(n_32),
.B2(n_13),
.Y(n_59)
);

MAJIxp5_ASAP7_75t_L g55 ( 
.A(n_52),
.B(n_45),
.C(n_40),
.Y(n_55)
);

XOR2xp5_ASAP7_75t_L g61 ( 
.A(n_55),
.B(n_54),
.Y(n_61)
);

OAI21xp33_ASAP7_75t_SL g56 ( 
.A1(n_48),
.A2(n_37),
.B(n_42),
.Y(n_56)
);

XOR2xp5_ASAP7_75t_L g63 ( 
.A(n_56),
.B(n_52),
.Y(n_63)
);

OAI22xp5_ASAP7_75t_L g57 ( 
.A1(n_50),
.A2(n_46),
.B1(n_37),
.B2(n_39),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_L g64 ( 
.A(n_57),
.B(n_58),
.Y(n_64)
);

OAI22xp5_ASAP7_75t_SL g58 ( 
.A1(n_49),
.A2(n_31),
.B1(n_29),
.B2(n_32),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_59),
.B(n_60),
.Y(n_62)
);

OAI22xp5_ASAP7_75t_SL g60 ( 
.A1(n_51),
.A2(n_32),
.B1(n_13),
.B2(n_19),
.Y(n_60)
);

XOR2xp5_ASAP7_75t_L g66 ( 
.A(n_61),
.B(n_63),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_L g65 ( 
.A(n_61),
.B(n_53),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_SL g69 ( 
.A(n_65),
.B(n_67),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_L g67 ( 
.A(n_64),
.B(n_54),
.Y(n_67)
);

AOI322xp5_ASAP7_75t_L g68 ( 
.A1(n_66),
.A2(n_57),
.A3(n_62),
.B1(n_55),
.B2(n_48),
.C1(n_60),
.C2(n_58),
.Y(n_68)
);

OAI21xp5_ASAP7_75t_L g70 ( 
.A1(n_68),
.A2(n_66),
.B(n_13),
.Y(n_70)
);

OAI31xp33_ASAP7_75t_SL g71 ( 
.A1(n_70),
.A2(n_69),
.A3(n_8),
.B(n_9),
.Y(n_71)
);


endmodule