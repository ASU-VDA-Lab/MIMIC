module real_jpeg_26439_n_12 (n_5, n_4, n_8, n_0, n_1, n_11, n_2, n_6, n_7, n_3, n_10, n_9, n_12);

input n_5;
input n_4;
input n_8;
input n_0;
input n_1;
input n_11;
input n_2;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_12;

wire n_37;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_300;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_13;
wire n_199;
wire n_95;
wire n_238;
wire n_67;
wire n_235;
wire n_107;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_123;
wire n_50;
wire n_186;
wire n_137;
wire n_72;
wire n_171;
wire n_151;
wire n_272;
wire n_203;
wire n_198;
wire n_23;
wire n_71;
wire n_61;
wire n_99;
wire n_80;
wire n_30;
wire n_149;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_230;
wire n_128;
wire n_202;
wire n_216;
wire n_127;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_252;
wire n_310;
wire n_78;
wire n_83;
wire n_288;
wire n_221;
wire n_104;
wire n_153;
wire n_131;
wire n_87;
wire n_40;
wire n_98;
wire n_200;
wire n_214;
wire n_113;
wire n_251;
wire n_139;
wire n_33;
wire n_175;
wire n_156;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_77;
wire n_219;
wire n_122;
wire n_19;
wire n_262;
wire n_17;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_20;
wire n_314;
wire n_278;
wire n_103;
wire n_232;
wire n_212;
wire n_284;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_213;
wire n_25;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_49;
wire n_68;
wire n_146;
wire n_286;
wire n_166;
wire n_176;
wire n_215;
wire n_312;
wire n_307;
wire n_316;
wire n_161;
wire n_207;
wire n_237;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_140;
wire n_126;
wire n_120;
wire n_155;
wire n_319;
wire n_93;
wire n_242;
wire n_142;
wire n_76;
wire n_79;
wire n_282;
wire n_147;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_18;
wire n_145;
wire n_266;
wire n_109;
wire n_148;
wire n_196;
wire n_298;
wire n_152;
wire n_270;
wire n_159;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_258;
wire n_150;
wire n_41;
wire n_74;
wire n_158;
wire n_204;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_75;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_119;
wire n_283;
wire n_181;
wire n_256;
wire n_253;
wire n_273;
wire n_16;
wire n_54;
wire n_168;
wire n_38;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_292;
wire n_64;
wire n_291;
wire n_236;
wire n_276;
wire n_287;
wire n_174;
wire n_255;
wire n_243;
wire n_299;
wire n_56;
wire n_293;
wire n_275;
wire n_227;
wire n_229;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_45;
wire n_268;
wire n_42;
wire n_313;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_143;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_303;
wire n_100;
wire n_51;
wire n_14;
wire n_205;
wire n_261;
wire n_86;
wire n_70;
wire n_32;
wire n_228;
wire n_15;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_133;
wire n_257;
wire n_210;
wire n_206;
wire n_85;
wire n_96;
wire n_308;

INVx3_ASAP7_75t_L g109 ( 
.A(n_0),
.Y(n_109)
);

INVx2_ASAP7_75t_L g110 ( 
.A(n_0),
.Y(n_110)
);

INVx6_ASAP7_75t_L g131 ( 
.A(n_0),
.Y(n_131)
);

INVx6_ASAP7_75t_L g262 ( 
.A(n_0),
.Y(n_262)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_1),
.Y(n_44)
);

AOI22xp33_ASAP7_75t_L g49 ( 
.A1(n_2),
.A2(n_43),
.B1(n_45),
.B2(n_50),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_2),
.Y(n_50)
);

OAI22xp5_ASAP7_75t_SL g67 ( 
.A1(n_2),
.A2(n_50),
.B1(n_68),
.B2(n_69),
.Y(n_67)
);

OAI22xp5_ASAP7_75t_L g94 ( 
.A1(n_2),
.A2(n_22),
.B1(n_27),
.B2(n_50),
.Y(n_94)
);

AOI22xp5_ASAP7_75t_L g134 ( 
.A1(n_2),
.A2(n_29),
.B1(n_31),
.B2(n_50),
.Y(n_134)
);

BUFx12f_ASAP7_75t_L g26 ( 
.A(n_3),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_4),
.Y(n_30)
);

BUFx10_ASAP7_75t_L g60 ( 
.A(n_5),
.Y(n_60)
);

OAI22xp33_ASAP7_75t_SL g142 ( 
.A1(n_6),
.A2(n_9),
.B1(n_54),
.B2(n_143),
.Y(n_142)
);

CKINVDCx20_ASAP7_75t_R g143 ( 
.A(n_6),
.Y(n_143)
);

OAI22xp33_ASAP7_75t_SL g190 ( 
.A1(n_6),
.A2(n_43),
.B1(n_45),
.B2(n_143),
.Y(n_190)
);

OAI22xp5_ASAP7_75t_L g230 ( 
.A1(n_6),
.A2(n_22),
.B1(n_27),
.B2(n_143),
.Y(n_230)
);

OAI22xp5_ASAP7_75t_SL g255 ( 
.A1(n_6),
.A2(n_29),
.B1(n_31),
.B2(n_143),
.Y(n_255)
);

OAI22xp5_ASAP7_75t_SL g52 ( 
.A1(n_7),
.A2(n_53),
.B1(n_55),
.B2(n_56),
.Y(n_52)
);

CKINVDCx20_ASAP7_75t_R g55 ( 
.A(n_7),
.Y(n_55)
);

OAI22xp5_ASAP7_75t_SL g88 ( 
.A1(n_7),
.A2(n_43),
.B1(n_45),
.B2(n_55),
.Y(n_88)
);

AOI22xp5_ASAP7_75t_SL g114 ( 
.A1(n_7),
.A2(n_22),
.B1(n_27),
.B2(n_55),
.Y(n_114)
);

AOI22xp5_ASAP7_75t_SL g167 ( 
.A1(n_7),
.A2(n_29),
.B1(n_31),
.B2(n_55),
.Y(n_167)
);

BUFx5_ASAP7_75t_L g39 ( 
.A(n_8),
.Y(n_39)
);

INVx13_ASAP7_75t_L g54 ( 
.A(n_9),
.Y(n_54)
);

BUFx12f_ASAP7_75t_L g23 ( 
.A(n_10),
.Y(n_23)
);

OAI22xp5_ASAP7_75t_SL g34 ( 
.A1(n_11),
.A2(n_22),
.B1(n_27),
.B2(n_35),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_11),
.Y(n_35)
);

OAI22xp5_ASAP7_75t_L g42 ( 
.A1(n_11),
.A2(n_35),
.B1(n_43),
.B2(n_45),
.Y(n_42)
);

OAI22xp5_ASAP7_75t_SL g79 ( 
.A1(n_11),
.A2(n_35),
.B1(n_54),
.B2(n_65),
.Y(n_79)
);

AOI22xp5_ASAP7_75t_L g111 ( 
.A1(n_11),
.A2(n_29),
.B1(n_31),
.B2(n_35),
.Y(n_111)
);

O2A1O1Ixp33_ASAP7_75t_L g202 ( 
.A1(n_11),
.A2(n_60),
.B(n_69),
.C(n_203),
.Y(n_202)
);

NAND2xp5_ASAP7_75t_L g215 ( 
.A(n_11),
.B(n_58),
.Y(n_215)
);

O2A1O1Ixp33_ASAP7_75t_L g225 ( 
.A1(n_11),
.A2(n_39),
.B(n_45),
.C(n_226),
.Y(n_225)
);

MAJIxp5_ASAP7_75t_L g243 ( 
.A(n_11),
.B(n_25),
.C(n_29),
.Y(n_243)
);

NAND2xp5_ASAP7_75t_SL g247 ( 
.A(n_11),
.B(n_89),
.Y(n_247)
);

NAND2xp5_ASAP7_75t_L g268 ( 
.A(n_11),
.B(n_269),
.Y(n_268)
);

NAND2xp5_ASAP7_75t_SL g273 ( 
.A(n_11),
.B(n_28),
.Y(n_273)
);

XNOR2xp5_ASAP7_75t_L g12 ( 
.A(n_13),
.B(n_82),
.Y(n_12)
);

NAND2xp5_ASAP7_75t_L g13 ( 
.A(n_14),
.B(n_80),
.Y(n_13)
);

NAND2xp5_ASAP7_75t_SL g14 ( 
.A(n_15),
.B(n_76),
.Y(n_14)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_15),
.B(n_76),
.Y(n_81)
);

MAJIxp5_ASAP7_75t_L g15 ( 
.A(n_16),
.B(n_70),
.C(n_71),
.Y(n_15)
);

AOI22xp33_ASAP7_75t_SL g316 ( 
.A1(n_16),
.A2(n_17),
.B1(n_317),
.B2(n_318),
.Y(n_316)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_17),
.Y(n_16)
);

MAJIxp5_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_36),
.C(n_51),
.Y(n_17)
);

OAI22xp5_ASAP7_75t_L g98 ( 
.A1(n_18),
.A2(n_99),
.B1(n_100),
.B2(n_103),
.Y(n_98)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_18),
.Y(n_103)
);

OAI22xp5_ASAP7_75t_SL g149 ( 
.A1(n_18),
.A2(n_36),
.B1(n_103),
.B2(n_150),
.Y(n_149)
);

OAI22xp5_ASAP7_75t_SL g211 ( 
.A1(n_18),
.A2(n_103),
.B1(n_187),
.B2(n_212),
.Y(n_211)
);

AOI21xp5_ASAP7_75t_SL g18 ( 
.A1(n_19),
.A2(n_32),
.B(n_33),
.Y(n_18)
);

OAI21xp5_ASAP7_75t_SL g113 ( 
.A1(n_19),
.A2(n_114),
.B(n_115),
.Y(n_113)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_20),
.Y(n_19)
);

NAND2xp5_ASAP7_75t_SL g93 ( 
.A(n_20),
.B(n_94),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_SL g171 ( 
.A(n_20),
.B(n_34),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_L g229 ( 
.A(n_20),
.B(n_230),
.Y(n_229)
);

NOR2xp33_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_28),
.Y(n_20)
);

AOI22xp33_ASAP7_75t_L g21 ( 
.A1(n_22),
.A2(n_24),
.B1(n_25),
.B2(n_27),
.Y(n_21)
);

INVx4_ASAP7_75t_L g27 ( 
.A(n_22),
.Y(n_27)
);

AOI22xp5_ASAP7_75t_L g38 ( 
.A1(n_22),
.A2(n_27),
.B1(n_39),
.B2(n_40),
.Y(n_38)
);

NAND2xp5_ASAP7_75t_L g242 ( 
.A(n_22),
.B(n_243),
.Y(n_242)
);

BUFx12f_ASAP7_75t_L g22 ( 
.A(n_23),
.Y(n_22)
);

OAI22xp5_ASAP7_75t_SL g28 ( 
.A1(n_24),
.A2(n_25),
.B1(n_29),
.B2(n_31),
.Y(n_28)
);

INVx13_ASAP7_75t_L g24 ( 
.A(n_25),
.Y(n_24)
);

BUFx24_ASAP7_75t_L g25 ( 
.A(n_26),
.Y(n_25)
);

OAI21xp33_ASAP7_75t_L g226 ( 
.A1(n_27),
.A2(n_35),
.B(n_40),
.Y(n_226)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_28),
.Y(n_32)
);

NAND2xp5_ASAP7_75t_L g115 ( 
.A(n_28),
.B(n_94),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_SL g240 ( 
.A(n_28),
.B(n_230),
.Y(n_240)
);

INVx6_ASAP7_75t_SL g31 ( 
.A(n_29),
.Y(n_31)
);

NAND2xp5_ASAP7_75t_L g108 ( 
.A(n_29),
.B(n_109),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_SL g267 ( 
.A(n_29),
.B(n_268),
.Y(n_267)
);

BUFx12f_ASAP7_75t_L g29 ( 
.A(n_30),
.Y(n_29)
);

NOR2xp33_ASAP7_75t_SL g91 ( 
.A(n_32),
.B(n_33),
.Y(n_91)
);

OAI21xp5_ASAP7_75t_L g135 ( 
.A1(n_32),
.A2(n_93),
.B(n_114),
.Y(n_135)
);

CKINVDCx16_ASAP7_75t_R g33 ( 
.A(n_34),
.Y(n_33)
);

OAI21xp33_ASAP7_75t_L g203 ( 
.A1(n_35),
.A2(n_45),
.B(n_59),
.Y(n_203)
);

CKINVDCx20_ASAP7_75t_R g150 ( 
.A(n_36),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_L g36 ( 
.A(n_37),
.B(n_46),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_SL g195 ( 
.A(n_37),
.B(n_196),
.Y(n_195)
);

NOR2xp33_ASAP7_75t_L g37 ( 
.A(n_38),
.B(n_41),
.Y(n_37)
);

NAND2xp5_ASAP7_75t_L g47 ( 
.A(n_38),
.B(n_48),
.Y(n_47)
);

AOI21xp5_ASAP7_75t_L g70 ( 
.A1(n_38),
.A2(n_41),
.B(n_47),
.Y(n_70)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_38),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_SL g102 ( 
.A(n_38),
.B(n_49),
.Y(n_102)
);

INVx2_ASAP7_75t_L g40 ( 
.A(n_39),
.Y(n_40)
);

OAI22xp5_ASAP7_75t_L g48 ( 
.A1(n_39),
.A2(n_40),
.B1(n_43),
.B2(n_45),
.Y(n_48)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_42),
.Y(n_41)
);

NAND2xp5_ASAP7_75t_SL g138 ( 
.A(n_42),
.B(n_101),
.Y(n_138)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_43),
.Y(n_45)
);

OAI22xp5_ASAP7_75t_L g58 ( 
.A1(n_43),
.A2(n_45),
.B1(n_59),
.B2(n_60),
.Y(n_58)
);

BUFx12f_ASAP7_75t_L g43 ( 
.A(n_44),
.Y(n_43)
);

AOI21xp5_ASAP7_75t_L g87 ( 
.A1(n_46),
.A2(n_88),
.B(n_89),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_SL g187 ( 
.A(n_46),
.B(n_188),
.Y(n_187)
);

NOR2xp33_ASAP7_75t_SL g46 ( 
.A(n_47),
.B(n_49),
.Y(n_46)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_47),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_SL g196 ( 
.A(n_47),
.B(n_197),
.Y(n_196)
);

XNOR2xp5_ASAP7_75t_L g148 ( 
.A(n_51),
.B(n_149),
.Y(n_148)
);

AOI21xp5_ASAP7_75t_L g51 ( 
.A1(n_52),
.A2(n_58),
.B(n_61),
.Y(n_51)
);

CKINVDCx20_ASAP7_75t_R g74 ( 
.A(n_52),
.Y(n_74)
);

INVx8_ASAP7_75t_L g66 ( 
.A(n_53),
.Y(n_66)
);

INVx11_ASAP7_75t_L g53 ( 
.A(n_54),
.Y(n_53)
);

INVx8_ASAP7_75t_L g57 ( 
.A(n_54),
.Y(n_57)
);

INVx8_ASAP7_75t_L g65 ( 
.A(n_54),
.Y(n_65)
);

INVx6_ASAP7_75t_L g68 ( 
.A(n_54),
.Y(n_68)
);

INVx11_ASAP7_75t_L g56 ( 
.A(n_57),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_58),
.B(n_64),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_L g75 ( 
.A(n_58),
.B(n_67),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_SL g78 ( 
.A(n_58),
.B(n_79),
.Y(n_78)
);

INVxp67_ASAP7_75t_L g118 ( 
.A(n_58),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_L g173 ( 
.A(n_58),
.B(n_142),
.Y(n_173)
);

AOI22xp33_ASAP7_75t_L g64 ( 
.A1(n_59),
.A2(n_60),
.B1(n_65),
.B2(n_66),
.Y(n_64)
);

INVx4_ASAP7_75t_L g59 ( 
.A(n_60),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_SL g76 ( 
.A(n_61),
.B(n_77),
.Y(n_76)
);

CKINVDCx14_ASAP7_75t_R g61 ( 
.A(n_62),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_L g172 ( 
.A(n_62),
.B(n_173),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_SL g62 ( 
.A(n_63),
.B(n_67),
.Y(n_62)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_63),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_L g97 ( 
.A(n_63),
.B(n_79),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g141 ( 
.A(n_63),
.B(n_142),
.Y(n_141)
);

INVx4_ASAP7_75t_L g69 ( 
.A(n_65),
.Y(n_69)
);

MAJIxp5_ASAP7_75t_L g163 ( 
.A(n_70),
.B(n_164),
.C(n_172),
.Y(n_163)
);

OAI22xp5_ASAP7_75t_SL g301 ( 
.A1(n_70),
.A2(n_172),
.B1(n_302),
.B2(n_303),
.Y(n_301)
);

CKINVDCx14_ASAP7_75t_R g302 ( 
.A(n_70),
.Y(n_302)
);

OAI22xp5_ASAP7_75t_L g317 ( 
.A1(n_70),
.A2(n_71),
.B1(n_72),
.B2(n_302),
.Y(n_317)
);

CKINVDCx20_ASAP7_75t_R g71 ( 
.A(n_72),
.Y(n_71)
);

OAI21xp5_ASAP7_75t_SL g72 ( 
.A1(n_73),
.A2(n_74),
.B(n_75),
.Y(n_72)
);

AOI21xp5_ASAP7_75t_SL g117 ( 
.A1(n_73),
.A2(n_118),
.B(n_119),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_SL g96 ( 
.A(n_75),
.B(n_97),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g198 ( 
.A(n_75),
.B(n_141),
.Y(n_198)
);

INVxp33_ASAP7_75t_L g77 ( 
.A(n_78),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_L g140 ( 
.A(n_78),
.B(n_141),
.Y(n_140)
);

INVxp67_ASAP7_75t_L g119 ( 
.A(n_79),
.Y(n_119)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_81),
.Y(n_80)
);

AOI21xp5_ASAP7_75t_L g82 ( 
.A1(n_83),
.A2(n_315),
.B(n_320),
.Y(n_82)
);

OAI211xp5_ASAP7_75t_L g83 ( 
.A1(n_84),
.A2(n_144),
.B(n_153),
.C(n_314),
.Y(n_83)
);

OR2x2_ASAP7_75t_L g84 ( 
.A(n_85),
.B(n_120),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g145 ( 
.A(n_85),
.B(n_146),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_L g154 ( 
.A(n_85),
.B(n_120),
.Y(n_154)
);

OR2x2_ASAP7_75t_L g314 ( 
.A(n_85),
.B(n_146),
.Y(n_314)
);

FAx1_ASAP7_75t_L g85 ( 
.A(n_86),
.B(n_95),
.CI(n_106),
.CON(n_85),
.SN(n_85)
);

OAI21xp5_ASAP7_75t_SL g125 ( 
.A1(n_86),
.A2(n_87),
.B(n_90),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_L g86 ( 
.A(n_87),
.B(n_90),
.Y(n_86)
);

AOI21xp5_ASAP7_75t_L g100 ( 
.A1(n_88),
.A2(n_101),
.B(n_102),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_L g189 ( 
.A(n_89),
.B(n_190),
.Y(n_189)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_91),
.B(n_92),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g227 ( 
.A(n_91),
.B(n_228),
.Y(n_227)
);

INVxp33_ASAP7_75t_L g92 ( 
.A(n_93),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_L g283 ( 
.A(n_93),
.B(n_240),
.Y(n_283)
);

OAI22xp5_ASAP7_75t_L g95 ( 
.A1(n_96),
.A2(n_98),
.B1(n_104),
.B2(n_105),
.Y(n_95)
);

CKINVDCx20_ASAP7_75t_R g104 ( 
.A(n_96),
.Y(n_104)
);

OAI22xp5_ASAP7_75t_L g147 ( 
.A1(n_96),
.A2(n_104),
.B1(n_148),
.B2(n_151),
.Y(n_147)
);

MAJIxp5_ASAP7_75t_L g152 ( 
.A(n_96),
.B(n_100),
.C(n_103),
.Y(n_152)
);

MAJIxp5_ASAP7_75t_L g319 ( 
.A(n_96),
.B(n_148),
.C(n_152),
.Y(n_319)
);

NAND2xp5_ASAP7_75t_L g186 ( 
.A(n_97),
.B(n_173),
.Y(n_186)
);

CKINVDCx16_ASAP7_75t_R g105 ( 
.A(n_98),
.Y(n_105)
);

CKINVDCx16_ASAP7_75t_R g99 ( 
.A(n_100),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g136 ( 
.A(n_102),
.B(n_137),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_L g218 ( 
.A(n_102),
.B(n_196),
.Y(n_218)
);

MAJIxp5_ASAP7_75t_L g184 ( 
.A(n_103),
.B(n_185),
.C(n_187),
.Y(n_184)
);

AOI21xp33_ASAP7_75t_L g106 ( 
.A1(n_107),
.A2(n_112),
.B(n_116),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_L g112 ( 
.A(n_107),
.B(n_113),
.Y(n_112)
);

OAI22xp5_ASAP7_75t_L g123 ( 
.A1(n_107),
.A2(n_116),
.B1(n_117),
.B2(n_124),
.Y(n_123)
);

CKINVDCx16_ASAP7_75t_R g124 ( 
.A(n_107),
.Y(n_124)
);

AOI22xp5_ASAP7_75t_L g161 ( 
.A1(n_107),
.A2(n_113),
.B1(n_124),
.B2(n_162),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_L g224 ( 
.A(n_107),
.B(n_225),
.Y(n_224)
);

OAI22xp5_ASAP7_75t_L g284 ( 
.A1(n_107),
.A2(n_124),
.B1(n_225),
.B2(n_285),
.Y(n_284)
);

AOI21xp5_ASAP7_75t_L g107 ( 
.A1(n_108),
.A2(n_110),
.B(n_111),
.Y(n_107)
);

OR2x2_ASAP7_75t_L g133 ( 
.A(n_108),
.B(n_134),
.Y(n_133)
);

OAI21xp5_ASAP7_75t_SL g166 ( 
.A1(n_108),
.A2(n_167),
.B(n_168),
.Y(n_166)
);

NOR2xp33_ASAP7_75t_SL g217 ( 
.A(n_108),
.B(n_111),
.Y(n_217)
);

NOR2xp33_ASAP7_75t_SL g253 ( 
.A(n_108),
.B(n_254),
.Y(n_253)
);

NOR2xp33_ASAP7_75t_L g169 ( 
.A(n_110),
.B(n_134),
.Y(n_169)
);

BUFx2_ASAP7_75t_L g205 ( 
.A(n_110),
.Y(n_205)
);

INVxp67_ASAP7_75t_L g132 ( 
.A(n_111),
.Y(n_132)
);

XOR2xp5_ASAP7_75t_L g122 ( 
.A(n_112),
.B(n_123),
.Y(n_122)
);

CKINVDCx20_ASAP7_75t_R g162 ( 
.A(n_113),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_SL g170 ( 
.A(n_115),
.B(n_171),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_SL g248 ( 
.A(n_115),
.B(n_229),
.Y(n_248)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_117),
.Y(n_116)
);

MAJIxp5_ASAP7_75t_L g120 ( 
.A(n_121),
.B(n_125),
.C(n_126),
.Y(n_120)
);

OAI22xp5_ASAP7_75t_SL g175 ( 
.A1(n_121),
.A2(n_122),
.B1(n_125),
.B2(n_176),
.Y(n_175)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_122),
.Y(n_121)
);

CKINVDCx20_ASAP7_75t_R g176 ( 
.A(n_125),
.Y(n_176)
);

XOR2xp5_ASAP7_75t_L g174 ( 
.A(n_126),
.B(n_175),
.Y(n_174)
);

MAJIxp5_ASAP7_75t_L g126 ( 
.A(n_127),
.B(n_136),
.C(n_139),
.Y(n_126)
);

XOR2xp5_ASAP7_75t_L g158 ( 
.A(n_127),
.B(n_159),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_128),
.B(n_135),
.Y(n_127)
);

XOR2xp5_ASAP7_75t_L g305 ( 
.A(n_128),
.B(n_135),
.Y(n_305)
);

NAND2xp5_ASAP7_75t_L g128 ( 
.A(n_129),
.B(n_133),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_L g251 ( 
.A(n_129),
.B(n_252),
.Y(n_251)
);

NAND2xp5_ASAP7_75t_L g129 ( 
.A(n_130),
.B(n_132),
.Y(n_129)
);

INVx2_ASAP7_75t_L g130 ( 
.A(n_131),
.Y(n_130)
);

OAI21xp5_ASAP7_75t_L g204 ( 
.A1(n_133),
.A2(n_167),
.B(n_205),
.Y(n_204)
);

NAND2xp5_ASAP7_75t_L g259 ( 
.A(n_133),
.B(n_260),
.Y(n_259)
);

OAI22xp5_ASAP7_75t_SL g159 ( 
.A1(n_136),
.A2(n_139),
.B1(n_140),
.B2(n_160),
.Y(n_159)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_136),
.Y(n_160)
);

CKINVDCx14_ASAP7_75t_R g137 ( 
.A(n_138),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_L g282 ( 
.A(n_138),
.B(n_189),
.Y(n_282)
);

CKINVDCx20_ASAP7_75t_R g139 ( 
.A(n_140),
.Y(n_139)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_145),
.Y(n_144)
);

NAND3xp33_ASAP7_75t_SL g153 ( 
.A(n_145),
.B(n_154),
.C(n_155),
.Y(n_153)
);

XNOR2xp5_ASAP7_75t_L g146 ( 
.A(n_147),
.B(n_152),
.Y(n_146)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_148),
.Y(n_151)
);

OAI21xp5_ASAP7_75t_L g155 ( 
.A1(n_156),
.A2(n_177),
.B(n_313),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_L g156 ( 
.A(n_157),
.B(n_174),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_SL g313 ( 
.A(n_157),
.B(n_174),
.Y(n_313)
);

MAJIxp5_ASAP7_75t_L g157 ( 
.A(n_158),
.B(n_161),
.C(n_163),
.Y(n_157)
);

XOR2xp5_ASAP7_75t_L g311 ( 
.A(n_158),
.B(n_161),
.Y(n_311)
);

XOR2xp5_ASAP7_75t_L g310 ( 
.A(n_163),
.B(n_311),
.Y(n_310)
);

AOI22xp5_ASAP7_75t_L g299 ( 
.A1(n_164),
.A2(n_165),
.B1(n_300),
.B2(n_301),
.Y(n_299)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_165),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_L g165 ( 
.A(n_166),
.B(n_170),
.Y(n_165)
);

XNOR2xp5_ASAP7_75t_L g183 ( 
.A(n_166),
.B(n_170),
.Y(n_183)
);

INVxp67_ASAP7_75t_L g168 ( 
.A(n_169),
.Y(n_168)
);

NOR2xp33_ASAP7_75t_L g216 ( 
.A(n_169),
.B(n_217),
.Y(n_216)
);

NOR2xp33_ASAP7_75t_L g274 ( 
.A(n_169),
.B(n_253),
.Y(n_274)
);

NAND2xp5_ASAP7_75t_L g239 ( 
.A(n_171),
.B(n_240),
.Y(n_239)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_172),
.Y(n_303)
);

AOI21xp5_ASAP7_75t_L g177 ( 
.A1(n_178),
.A2(n_308),
.B(n_312),
.Y(n_177)
);

A2O1A1Ixp33_ASAP7_75t_SL g178 ( 
.A1(n_179),
.A2(n_219),
.B(n_294),
.C(n_307),
.Y(n_178)
);

OR2x2_ASAP7_75t_L g179 ( 
.A(n_180),
.B(n_207),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_L g293 ( 
.A(n_180),
.B(n_207),
.Y(n_293)
);

AOI22xp5_ASAP7_75t_SL g180 ( 
.A1(n_181),
.A2(n_182),
.B1(n_193),
.B2(n_206),
.Y(n_180)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_182),
.Y(n_181)
);

OAI22xp5_ASAP7_75t_L g182 ( 
.A1(n_183),
.A2(n_184),
.B1(n_191),
.B2(n_192),
.Y(n_182)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_183),
.Y(n_191)
);

MAJIxp5_ASAP7_75t_L g295 ( 
.A(n_183),
.B(n_192),
.C(n_206),
.Y(n_295)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_184),
.Y(n_192)
);

AOI22xp5_ASAP7_75t_L g209 ( 
.A1(n_185),
.A2(n_186),
.B1(n_210),
.B2(n_211),
.Y(n_209)
);

CKINVDCx20_ASAP7_75t_R g185 ( 
.A(n_186),
.Y(n_185)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_187),
.Y(n_212)
);

CKINVDCx16_ASAP7_75t_R g188 ( 
.A(n_189),
.Y(n_188)
);

INVxp67_ASAP7_75t_SL g197 ( 
.A(n_190),
.Y(n_197)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_193),
.Y(n_206)
);

XOR2xp5_ASAP7_75t_L g193 ( 
.A(n_194),
.B(n_201),
.Y(n_193)
);

AOI22xp5_ASAP7_75t_L g194 ( 
.A1(n_195),
.A2(n_198),
.B1(n_199),
.B2(n_200),
.Y(n_194)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_195),
.Y(n_199)
);

MAJIxp5_ASAP7_75t_L g306 ( 
.A(n_195),
.B(n_200),
.C(n_201),
.Y(n_306)
);

CKINVDCx20_ASAP7_75t_R g200 ( 
.A(n_198),
.Y(n_200)
);

NAND2xp5_ASAP7_75t_L g201 ( 
.A(n_202),
.B(n_204),
.Y(n_201)
);

XOR2xp5_ASAP7_75t_L g213 ( 
.A(n_202),
.B(n_204),
.Y(n_213)
);

MAJIxp5_ASAP7_75t_L g207 ( 
.A(n_208),
.B(n_213),
.C(n_214),
.Y(n_207)
);

OAI22xp5_ASAP7_75t_SL g231 ( 
.A1(n_208),
.A2(n_209),
.B1(n_232),
.B2(n_233),
.Y(n_231)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_209),
.Y(n_208)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_211),
.Y(n_210)
);

XOR2xp5_ASAP7_75t_L g233 ( 
.A(n_213),
.B(n_214),
.Y(n_233)
);

CKINVDCx5p33_ASAP7_75t_R g223 ( 
.A(n_214),
.Y(n_223)
);

FAx1_ASAP7_75t_L g214 ( 
.A(n_215),
.B(n_216),
.CI(n_218),
.CON(n_214),
.SN(n_214)
);

NOR2xp33_ASAP7_75t_L g270 ( 
.A(n_217),
.B(n_271),
.Y(n_270)
);

NAND2xp5_ASAP7_75t_SL g219 ( 
.A(n_220),
.B(n_293),
.Y(n_219)
);

OAI21xp5_ASAP7_75t_L g220 ( 
.A1(n_221),
.A2(n_234),
.B(n_292),
.Y(n_220)
);

NOR2xp33_ASAP7_75t_L g221 ( 
.A(n_222),
.B(n_231),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_SL g292 ( 
.A(n_222),
.B(n_231),
.Y(n_292)
);

MAJIxp5_ASAP7_75t_L g222 ( 
.A(n_223),
.B(n_224),
.C(n_227),
.Y(n_222)
);

XOR2xp5_ASAP7_75t_L g289 ( 
.A(n_223),
.B(n_290),
.Y(n_289)
);

XOR2xp5_ASAP7_75t_L g290 ( 
.A(n_224),
.B(n_227),
.Y(n_290)
);

CKINVDCx16_ASAP7_75t_R g285 ( 
.A(n_225),
.Y(n_285)
);

INVxp33_ASAP7_75t_L g228 ( 
.A(n_229),
.Y(n_228)
);

CKINVDCx14_ASAP7_75t_R g232 ( 
.A(n_233),
.Y(n_232)
);

AOI21xp5_ASAP7_75t_L g234 ( 
.A1(n_235),
.A2(n_287),
.B(n_291),
.Y(n_234)
);

OAI21xp5_ASAP7_75t_SL g235 ( 
.A1(n_236),
.A2(n_278),
.B(n_286),
.Y(n_235)
);

AOI21xp5_ASAP7_75t_L g236 ( 
.A1(n_237),
.A2(n_257),
.B(n_277),
.Y(n_236)
);

NAND2xp5_ASAP7_75t_L g237 ( 
.A(n_238),
.B(n_244),
.Y(n_237)
);

NOR2xp33_ASAP7_75t_SL g277 ( 
.A(n_238),
.B(n_244),
.Y(n_277)
);

NAND2xp5_ASAP7_75t_SL g238 ( 
.A(n_239),
.B(n_241),
.Y(n_238)
);

OAI22xp5_ASAP7_75t_SL g263 ( 
.A1(n_239),
.A2(n_241),
.B1(n_242),
.B2(n_264),
.Y(n_263)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_239),
.Y(n_264)
);

CKINVDCx20_ASAP7_75t_R g241 ( 
.A(n_242),
.Y(n_241)
);

AOI22xp5_ASAP7_75t_SL g244 ( 
.A1(n_245),
.A2(n_246),
.B1(n_251),
.B2(n_256),
.Y(n_244)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_246),
.Y(n_245)
);

OAI22xp5_ASAP7_75t_L g246 ( 
.A1(n_247),
.A2(n_248),
.B1(n_249),
.B2(n_250),
.Y(n_246)
);

CKINVDCx14_ASAP7_75t_R g249 ( 
.A(n_247),
.Y(n_249)
);

MAJIxp5_ASAP7_75t_L g279 ( 
.A(n_247),
.B(n_250),
.C(n_256),
.Y(n_279)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_248),
.Y(n_250)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_251),
.Y(n_256)
);

INVxp67_ASAP7_75t_L g252 ( 
.A(n_253),
.Y(n_252)
);

CKINVDCx16_ASAP7_75t_R g254 ( 
.A(n_255),
.Y(n_254)
);

NAND2xp5_ASAP7_75t_SL g260 ( 
.A(n_255),
.B(n_261),
.Y(n_260)
);

OAI21xp5_ASAP7_75t_SL g257 ( 
.A1(n_258),
.A2(n_265),
.B(n_276),
.Y(n_257)
);

NOR2xp33_ASAP7_75t_L g258 ( 
.A(n_259),
.B(n_263),
.Y(n_258)
);

NAND2xp5_ASAP7_75t_SL g276 ( 
.A(n_259),
.B(n_263),
.Y(n_276)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_260),
.Y(n_271)
);

INVx3_ASAP7_75t_SL g261 ( 
.A(n_262),
.Y(n_261)
);

INVx8_ASAP7_75t_L g269 ( 
.A(n_262),
.Y(n_269)
);

AOI21xp5_ASAP7_75t_L g265 ( 
.A1(n_266),
.A2(n_272),
.B(n_275),
.Y(n_265)
);

NOR2xp33_ASAP7_75t_L g266 ( 
.A(n_267),
.B(n_270),
.Y(n_266)
);

NAND2xp5_ASAP7_75t_L g272 ( 
.A(n_273),
.B(n_274),
.Y(n_272)
);

NOR2xp33_ASAP7_75t_SL g275 ( 
.A(n_273),
.B(n_274),
.Y(n_275)
);

NOR2xp33_ASAP7_75t_L g278 ( 
.A(n_279),
.B(n_280),
.Y(n_278)
);

NAND2xp5_ASAP7_75t_SL g286 ( 
.A(n_279),
.B(n_280),
.Y(n_286)
);

XNOR2xp5_ASAP7_75t_L g280 ( 
.A(n_281),
.B(n_284),
.Y(n_280)
);

XNOR2xp5_ASAP7_75t_L g281 ( 
.A(n_282),
.B(n_283),
.Y(n_281)
);

MAJIxp5_ASAP7_75t_L g288 ( 
.A(n_282),
.B(n_283),
.C(n_284),
.Y(n_288)
);

NAND2xp5_ASAP7_75t_L g287 ( 
.A(n_288),
.B(n_289),
.Y(n_287)
);

NOR2xp33_ASAP7_75t_SL g291 ( 
.A(n_288),
.B(n_289),
.Y(n_291)
);

NOR2xp33_ASAP7_75t_L g294 ( 
.A(n_295),
.B(n_296),
.Y(n_294)
);

NAND2xp5_ASAP7_75t_SL g307 ( 
.A(n_295),
.B(n_296),
.Y(n_307)
);

XOR2xp5_ASAP7_75t_L g296 ( 
.A(n_297),
.B(n_306),
.Y(n_296)
);

OAI22xp5_ASAP7_75t_SL g297 ( 
.A1(n_298),
.A2(n_299),
.B1(n_304),
.B2(n_305),
.Y(n_297)
);

MAJIxp5_ASAP7_75t_L g309 ( 
.A(n_298),
.B(n_305),
.C(n_306),
.Y(n_309)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_299),
.Y(n_298)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_301),
.Y(n_300)
);

CKINVDCx16_ASAP7_75t_R g304 ( 
.A(n_305),
.Y(n_304)
);

NAND2xp5_ASAP7_75t_L g308 ( 
.A(n_309),
.B(n_310),
.Y(n_308)
);

NOR2xp33_ASAP7_75t_SL g312 ( 
.A(n_309),
.B(n_310),
.Y(n_312)
);

NAND2xp5_ASAP7_75t_L g315 ( 
.A(n_316),
.B(n_319),
.Y(n_315)
);

NOR2xp33_ASAP7_75t_SL g320 ( 
.A(n_316),
.B(n_319),
.Y(n_320)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_317),
.Y(n_318)
);


endmodule