module fake_netlist_5_1367_n_80 (n_16, n_0, n_12, n_9, n_18, n_1, n_8, n_10, n_4, n_11, n_17, n_19, n_7, n_15, n_5, n_14, n_2, n_13, n_3, n_6, n_80);

input n_16;
input n_0;
input n_12;
input n_9;
input n_18;
input n_1;
input n_8;
input n_10;
input n_4;
input n_11;
input n_17;
input n_19;
input n_7;
input n_15;
input n_5;
input n_14;
input n_2;
input n_13;
input n_3;
input n_6;

output n_80;

wire n_24;
wire n_61;
wire n_75;
wire n_65;
wire n_78;
wire n_74;
wire n_57;
wire n_37;
wire n_31;
wire n_66;
wire n_60;
wire n_43;
wire n_58;
wire n_69;
wire n_42;
wire n_22;
wire n_45;
wire n_46;
wire n_21;
wire n_38;
wire n_35;
wire n_73;
wire n_30;
wire n_33;
wire n_23;
wire n_29;
wire n_79;
wire n_47;
wire n_25;
wire n_53;
wire n_44;
wire n_40;
wire n_34;
wire n_62;
wire n_71;
wire n_59;
wire n_26;
wire n_55;
wire n_49;
wire n_20;
wire n_39;
wire n_54;
wire n_67;
wire n_36;
wire n_76;
wire n_27;
wire n_64;
wire n_77;
wire n_28;
wire n_70;
wire n_68;
wire n_72;
wire n_32;
wire n_41;
wire n_56;
wire n_51;
wire n_63;
wire n_48;
wire n_50;
wire n_52;

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_1),
.Y(n_20)
);

AOI22xp5_ASAP7_75t_SL g21 ( 
.A1(n_2),
.A2(n_15),
.B1(n_18),
.B2(n_14),
.Y(n_21)
);

HB1xp67_ASAP7_75t_L g22 ( 
.A(n_9),
.Y(n_22)
);

OAI21x1_ASAP7_75t_L g23 ( 
.A1(n_10),
.A2(n_13),
.B(n_3),
.Y(n_23)
);

INVx5_ASAP7_75t_L g24 ( 
.A(n_8),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_17),
.Y(n_25)
);

INVx2_ASAP7_75t_L g26 ( 
.A(n_19),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_2),
.Y(n_27)
);

BUFx3_ASAP7_75t_L g28 ( 
.A(n_3),
.Y(n_28)
);

INVx6_ASAP7_75t_L g29 ( 
.A(n_5),
.Y(n_29)
);

AOI22xp5_ASAP7_75t_L g30 ( 
.A1(n_7),
.A2(n_12),
.B1(n_6),
.B2(n_0),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_1),
.Y(n_31)
);

NOR2xp33_ASAP7_75t_L g32 ( 
.A(n_11),
.B(n_4),
.Y(n_32)
);

BUFx12f_ASAP7_75t_L g33 ( 
.A(n_0),
.Y(n_33)
);

NAND2xp5_ASAP7_75t_SL g34 ( 
.A(n_22),
.B(n_4),
.Y(n_34)
);

NAND2xp5_ASAP7_75t_SL g35 ( 
.A(n_20),
.B(n_27),
.Y(n_35)
);

NAND2xp5_ASAP7_75t_SL g36 ( 
.A(n_20),
.B(n_16),
.Y(n_36)
);

AOI22xp33_ASAP7_75t_L g37 ( 
.A1(n_28),
.A2(n_29),
.B1(n_33),
.B2(n_20),
.Y(n_37)
);

NAND2xp5_ASAP7_75t_SL g38 ( 
.A(n_20),
.B(n_27),
.Y(n_38)
);

INVxp67_ASAP7_75t_L g39 ( 
.A(n_31),
.Y(n_39)
);

NAND2xp5_ASAP7_75t_L g40 ( 
.A(n_26),
.B(n_27),
.Y(n_40)
);

OAI21xp5_ASAP7_75t_L g41 ( 
.A1(n_35),
.A2(n_23),
.B(n_30),
.Y(n_41)
);

AOI21xp5_ASAP7_75t_L g42 ( 
.A1(n_38),
.A2(n_32),
.B(n_24),
.Y(n_42)
);

O2A1O1Ixp5_ASAP7_75t_L g43 ( 
.A1(n_40),
.A2(n_32),
.B(n_21),
.C(n_29),
.Y(n_43)
);

AND2x2_ASAP7_75t_L g44 ( 
.A(n_39),
.B(n_28),
.Y(n_44)
);

BUFx2_ASAP7_75t_L g45 ( 
.A(n_37),
.Y(n_45)
);

NAND2xp5_ASAP7_75t_L g46 ( 
.A(n_36),
.B(n_24),
.Y(n_46)
);

INVx2_ASAP7_75t_L g47 ( 
.A(n_46),
.Y(n_47)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_44),
.Y(n_48)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_44),
.Y(n_49)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_42),
.Y(n_50)
);

INVx2_ASAP7_75t_SL g51 ( 
.A(n_45),
.Y(n_51)
);

AND2x4_ASAP7_75t_L g52 ( 
.A(n_41),
.B(n_34),
.Y(n_52)
);

AND2x2_ASAP7_75t_L g53 ( 
.A(n_45),
.B(n_29),
.Y(n_53)
);

INVx2_ASAP7_75t_L g54 ( 
.A(n_50),
.Y(n_54)
);

INVxp67_ASAP7_75t_L g55 ( 
.A(n_51),
.Y(n_55)
);

NAND2x1p5_ASAP7_75t_L g56 ( 
.A(n_52),
.B(n_24),
.Y(n_56)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_48),
.Y(n_57)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_49),
.Y(n_58)
);

INVxp67_ASAP7_75t_SL g59 ( 
.A(n_52),
.Y(n_59)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_54),
.Y(n_60)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_57),
.Y(n_61)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_58),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_SL g63 ( 
.A(n_55),
.B(n_51),
.Y(n_63)
);

AND2x2_ASAP7_75t_L g64 ( 
.A(n_59),
.B(n_52),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_L g65 ( 
.A(n_64),
.B(n_59),
.Y(n_65)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_60),
.Y(n_66)
);

INVxp67_ASAP7_75t_L g67 ( 
.A(n_63),
.Y(n_67)
);

AND2x2_ASAP7_75t_L g68 ( 
.A(n_64),
.B(n_55),
.Y(n_68)
);

AOI221xp5_ASAP7_75t_L g69 ( 
.A1(n_67),
.A2(n_43),
.B1(n_53),
.B2(n_62),
.C(n_61),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_68),
.B(n_56),
.Y(n_70)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_66),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_L g72 ( 
.A(n_65),
.B(n_56),
.Y(n_72)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_71),
.Y(n_73)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_69),
.Y(n_74)
);

BUFx12f_ASAP7_75t_L g75 ( 
.A(n_70),
.Y(n_75)
);

NOR2x1_ASAP7_75t_L g76 ( 
.A(n_74),
.B(n_72),
.Y(n_76)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_73),
.Y(n_77)
);

OAI22x1_ASAP7_75t_L g78 ( 
.A1(n_76),
.A2(n_75),
.B1(n_24),
.B2(n_47),
.Y(n_78)
);

OAI21xp33_ASAP7_75t_L g79 ( 
.A1(n_78),
.A2(n_77),
.B(n_25),
.Y(n_79)
);

OR2x6_ASAP7_75t_L g80 ( 
.A(n_79),
.B(n_25),
.Y(n_80)
);


endmodule