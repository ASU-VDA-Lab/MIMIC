module fake_netlist_6_3276_n_1376 (n_52, n_16, n_1, n_91, n_119, n_46, n_146, n_163, n_235, n_303, n_256, n_298, n_18, n_21, n_193, n_147, n_269, n_258, n_281, n_154, n_191, n_88, n_3, n_209, n_98, n_277, n_260, n_265, n_283, n_113, n_39, n_63, n_223, n_278, n_270, n_73, n_279, n_4, n_148, n_199, n_138, n_22, n_161, n_208, n_68, n_226, n_228, n_252, n_266, n_296, n_166, n_28, n_184, n_304, n_212, n_268, n_271, n_50, n_158, n_49, n_7, n_210, n_216, n_83, n_206, n_217, n_299, n_5, n_101, n_167, n_144, n_174, n_127, n_125, n_153, n_168, n_215, n_297, n_178, n_247, n_225, n_77, n_156, n_149, n_152, n_106, n_92, n_145, n_42, n_133, n_96, n_8, n_90, n_160, n_24, n_105, n_131, n_54, n_227, n_132, n_188, n_102, n_186, n_204, n_245, n_0, n_87, n_195, n_285, n_261, n_189, n_32, n_66, n_85, n_99, n_78, n_84, n_130, n_213, n_164, n_257, n_100, n_292, n_129, n_13, n_121, n_294, n_302, n_197, n_11, n_137, n_17, n_23, n_203, n_254, n_142, n_286, n_20, n_143, n_207, n_2, n_242, n_180, n_19, n_47, n_62, n_29, n_155, n_219, n_291, n_75, n_109, n_150, n_233, n_263, n_122, n_264, n_45, n_255, n_284, n_205, n_34, n_140, n_218, n_70, n_120, n_234, n_251, n_301, n_214, n_274, n_37, n_15, n_67, n_33, n_82, n_27, n_236, n_246, n_38, n_110, n_151, n_289, n_61, n_112, n_172, n_237, n_81, n_59, n_244, n_181, n_76, n_36, n_182, n_26, n_124, n_238, n_239, n_55, n_126, n_202, n_94, n_97, n_108, n_267, n_282, n_58, n_116, n_280, n_211, n_287, n_64, n_220, n_288, n_290, n_117, n_118, n_175, n_224, n_48, n_231, n_65, n_230, n_25, n_40, n_93, n_80, n_141, n_240, n_135, n_196, n_200, n_165, n_139, n_41, n_134, n_259, n_177, n_176, n_273, n_114, n_86, n_198, n_104, n_222, n_95, n_179, n_243, n_9, n_248, n_300, n_107, n_10, n_295, n_71, n_74, n_229, n_253, n_6, n_190, n_14, n_123, n_262, n_136, n_72, n_187, n_89, n_249, n_173, n_201, n_250, n_103, n_111, n_60, n_159, n_272, n_157, n_162, n_170, n_185, n_35, n_183, n_232, n_115, n_12, n_69, n_128, n_241, n_30, n_79, n_275, n_43, n_194, n_171, n_293, n_31, n_192, n_57, n_169, n_53, n_276, n_51, n_44, n_56, n_221, n_1376);

input n_52;
input n_16;
input n_1;
input n_91;
input n_119;
input n_46;
input n_146;
input n_163;
input n_235;
input n_303;
input n_256;
input n_298;
input n_18;
input n_21;
input n_193;
input n_147;
input n_269;
input n_258;
input n_281;
input n_154;
input n_191;
input n_88;
input n_3;
input n_209;
input n_98;
input n_277;
input n_260;
input n_265;
input n_283;
input n_113;
input n_39;
input n_63;
input n_223;
input n_278;
input n_270;
input n_73;
input n_279;
input n_4;
input n_148;
input n_199;
input n_138;
input n_22;
input n_161;
input n_208;
input n_68;
input n_226;
input n_228;
input n_252;
input n_266;
input n_296;
input n_166;
input n_28;
input n_184;
input n_304;
input n_212;
input n_268;
input n_271;
input n_50;
input n_158;
input n_49;
input n_7;
input n_210;
input n_216;
input n_83;
input n_206;
input n_217;
input n_299;
input n_5;
input n_101;
input n_167;
input n_144;
input n_174;
input n_127;
input n_125;
input n_153;
input n_168;
input n_215;
input n_297;
input n_178;
input n_247;
input n_225;
input n_77;
input n_156;
input n_149;
input n_152;
input n_106;
input n_92;
input n_145;
input n_42;
input n_133;
input n_96;
input n_8;
input n_90;
input n_160;
input n_24;
input n_105;
input n_131;
input n_54;
input n_227;
input n_132;
input n_188;
input n_102;
input n_186;
input n_204;
input n_245;
input n_0;
input n_87;
input n_195;
input n_285;
input n_261;
input n_189;
input n_32;
input n_66;
input n_85;
input n_99;
input n_78;
input n_84;
input n_130;
input n_213;
input n_164;
input n_257;
input n_100;
input n_292;
input n_129;
input n_13;
input n_121;
input n_294;
input n_302;
input n_197;
input n_11;
input n_137;
input n_17;
input n_23;
input n_203;
input n_254;
input n_142;
input n_286;
input n_20;
input n_143;
input n_207;
input n_2;
input n_242;
input n_180;
input n_19;
input n_47;
input n_62;
input n_29;
input n_155;
input n_219;
input n_291;
input n_75;
input n_109;
input n_150;
input n_233;
input n_263;
input n_122;
input n_264;
input n_45;
input n_255;
input n_284;
input n_205;
input n_34;
input n_140;
input n_218;
input n_70;
input n_120;
input n_234;
input n_251;
input n_301;
input n_214;
input n_274;
input n_37;
input n_15;
input n_67;
input n_33;
input n_82;
input n_27;
input n_236;
input n_246;
input n_38;
input n_110;
input n_151;
input n_289;
input n_61;
input n_112;
input n_172;
input n_237;
input n_81;
input n_59;
input n_244;
input n_181;
input n_76;
input n_36;
input n_182;
input n_26;
input n_124;
input n_238;
input n_239;
input n_55;
input n_126;
input n_202;
input n_94;
input n_97;
input n_108;
input n_267;
input n_282;
input n_58;
input n_116;
input n_280;
input n_211;
input n_287;
input n_64;
input n_220;
input n_288;
input n_290;
input n_117;
input n_118;
input n_175;
input n_224;
input n_48;
input n_231;
input n_65;
input n_230;
input n_25;
input n_40;
input n_93;
input n_80;
input n_141;
input n_240;
input n_135;
input n_196;
input n_200;
input n_165;
input n_139;
input n_41;
input n_134;
input n_259;
input n_177;
input n_176;
input n_273;
input n_114;
input n_86;
input n_198;
input n_104;
input n_222;
input n_95;
input n_179;
input n_243;
input n_9;
input n_248;
input n_300;
input n_107;
input n_10;
input n_295;
input n_71;
input n_74;
input n_229;
input n_253;
input n_6;
input n_190;
input n_14;
input n_123;
input n_262;
input n_136;
input n_72;
input n_187;
input n_89;
input n_249;
input n_173;
input n_201;
input n_250;
input n_103;
input n_111;
input n_60;
input n_159;
input n_272;
input n_157;
input n_162;
input n_170;
input n_185;
input n_35;
input n_183;
input n_232;
input n_115;
input n_12;
input n_69;
input n_128;
input n_241;
input n_30;
input n_79;
input n_275;
input n_43;
input n_194;
input n_171;
input n_293;
input n_31;
input n_192;
input n_57;
input n_169;
input n_53;
input n_276;
input n_51;
input n_44;
input n_56;
input n_221;

output n_1376;

wire n_992;
wire n_801;
wire n_1234;
wire n_1199;
wire n_741;
wire n_1027;
wire n_1351;
wire n_625;
wire n_1189;
wire n_1212;
wire n_726;
wire n_700;
wire n_1307;
wire n_1038;
wire n_578;
wire n_1003;
wire n_365;
wire n_1237;
wire n_1061;
wire n_1357;
wire n_783;
wire n_798;
wire n_509;
wire n_1342;
wire n_1209;
wire n_1348;
wire n_677;
wire n_805;
wire n_1151;
wire n_396;
wire n_350;
wire n_442;
wire n_480;
wire n_1009;
wire n_1160;
wire n_883;
wire n_1238;
wire n_1032;
wire n_1247;
wire n_893;
wire n_1099;
wire n_1264;
wire n_1192;
wire n_471;
wire n_424;
wire n_1370;
wire n_369;
wire n_415;
wire n_830;
wire n_461;
wire n_873;
wire n_383;
wire n_1285;
wire n_1371;
wire n_447;
wire n_1172;
wire n_852;
wire n_1078;
wire n_544;
wire n_1140;
wire n_1263;
wire n_836;
wire n_375;
wire n_522;
wire n_1261;
wire n_945;
wire n_1143;
wire n_1232;
wire n_658;
wire n_616;
wire n_1119;
wire n_428;
wire n_1300;
wire n_641;
wire n_822;
wire n_693;
wire n_1313;
wire n_1056;
wire n_758;
wire n_516;
wire n_1163;
wire n_1180;
wire n_943;
wire n_491;
wire n_772;
wire n_1344;
wire n_666;
wire n_371;
wire n_940;
wire n_770;
wire n_567;
wire n_405;
wire n_538;
wire n_1106;
wire n_886;
wire n_343;
wire n_953;
wire n_1094;
wire n_1345;
wire n_494;
wire n_539;
wire n_493;
wire n_454;
wire n_638;
wire n_1211;
wire n_381;
wire n_887;
wire n_1280;
wire n_713;
wire n_976;
wire n_734;
wire n_1088;
wire n_1231;
wire n_917;
wire n_574;
wire n_907;
wire n_659;
wire n_407;
wire n_913;
wire n_808;
wire n_867;
wire n_1230;
wire n_473;
wire n_1193;
wire n_1054;
wire n_559;
wire n_1333;
wire n_551;
wire n_699;
wire n_564;
wire n_451;
wire n_824;
wire n_686;
wire n_757;
wire n_594;
wire n_577;
wire n_619;
wire n_1367;
wire n_1336;
wire n_521;
wire n_572;
wire n_395;
wire n_813;
wire n_323;
wire n_606;
wire n_818;
wire n_1123;
wire n_1309;
wire n_513;
wire n_645;
wire n_331;
wire n_916;
wire n_483;
wire n_608;
wire n_630;
wire n_541;
wire n_512;
wire n_433;
wire n_792;
wire n_476;
wire n_1328;
wire n_1162;
wire n_860;
wire n_788;
wire n_939;
wire n_821;
wire n_938;
wire n_1302;
wire n_1068;
wire n_329;
wire n_982;
wire n_549;
wire n_1075;
wire n_408;
wire n_932;
wire n_979;
wire n_905;
wire n_322;
wire n_993;
wire n_689;
wire n_354;
wire n_1330;
wire n_1278;
wire n_547;
wire n_558;
wire n_1064;
wire n_634;
wire n_966;
wire n_764;
wire n_692;
wire n_733;
wire n_1233;
wire n_1289;
wire n_487;
wire n_1107;
wire n_1014;
wire n_1290;
wire n_882;
wire n_1354;
wire n_586;
wire n_423;
wire n_318;
wire n_1111;
wire n_715;
wire n_1251;
wire n_1265;
wire n_530;
wire n_618;
wire n_1297;
wire n_1312;
wire n_1167;
wire n_1359;
wire n_674;
wire n_871;
wire n_922;
wire n_1335;
wire n_1069;
wire n_612;
wire n_1165;
wire n_355;
wire n_702;
wire n_347;
wire n_1175;
wire n_328;
wire n_429;
wire n_1012;
wire n_780;
wire n_675;
wire n_903;
wire n_835;
wire n_928;
wire n_1214;
wire n_690;
wire n_850;
wire n_816;
wire n_1157;
wire n_1188;
wire n_877;
wire n_604;
wire n_825;
wire n_728;
wire n_1063;
wire n_1124;
wire n_515;
wire n_598;
wire n_696;
wire n_961;
wire n_437;
wire n_1082;
wire n_1317;
wire n_593;
wire n_514;
wire n_687;
wire n_697;
wire n_890;
wire n_637;
wire n_701;
wire n_950;
wire n_388;
wire n_484;
wire n_891;
wire n_949;
wire n_678;
wire n_507;
wire n_968;
wire n_909;
wire n_1369;
wire n_881;
wire n_1008;
wire n_760;
wire n_590;
wire n_362;
wire n_462;
wire n_1033;
wire n_1052;
wire n_1296;
wire n_694;
wire n_1294;
wire n_627;
wire n_595;
wire n_524;
wire n_342;
wire n_1044;
wire n_449;
wire n_1208;
wire n_1164;
wire n_1295;
wire n_1072;
wire n_495;
wire n_815;
wire n_1100;
wire n_585;
wire n_840;
wire n_874;
wire n_1128;
wire n_673;
wire n_382;
wire n_1071;
wire n_1067;
wire n_898;
wire n_865;
wire n_925;
wire n_1101;
wire n_1026;
wire n_1364;
wire n_615;
wire n_1249;
wire n_1293;
wire n_1127;
wire n_320;
wire n_639;
wire n_963;
wire n_794;
wire n_727;
wire n_894;
wire n_685;
wire n_353;
wire n_605;
wire n_826;
wire n_872;
wire n_1139;
wire n_718;
wire n_1018;
wire n_1366;
wire n_542;
wire n_847;
wire n_644;
wire n_682;
wire n_851;
wire n_305;
wire n_996;
wire n_532;
wire n_1308;
wire n_413;
wire n_791;
wire n_510;
wire n_837;
wire n_948;
wire n_704;
wire n_977;
wire n_1005;
wire n_536;
wire n_622;
wire n_581;
wire n_765;
wire n_432;
wire n_987;
wire n_1340;
wire n_631;
wire n_720;
wire n_842;
wire n_843;
wire n_656;
wire n_989;
wire n_1277;
wire n_797;
wire n_1246;
wire n_899;
wire n_738;
wire n_1304;
wire n_1035;
wire n_499;
wire n_705;
wire n_1004;
wire n_1176;
wire n_1022;
wire n_614;
wire n_529;
wire n_425;
wire n_684;
wire n_1181;
wire n_486;
wire n_947;
wire n_1117;
wire n_1087;
wire n_648;
wire n_657;
wire n_1049;
wire n_803;
wire n_926;
wire n_927;
wire n_919;
wire n_478;
wire n_929;
wire n_1228;
wire n_417;
wire n_446;
wire n_777;
wire n_1299;
wire n_526;
wire n_1183;
wire n_458;
wire n_1070;
wire n_998;
wire n_717;
wire n_1178;
wire n_1073;
wire n_1000;
wire n_796;
wire n_1195;
wire n_552;
wire n_1358;
wire n_912;
wire n_745;
wire n_1284;
wire n_1142;
wire n_716;
wire n_623;
wire n_1048;
wire n_1201;
wire n_884;
wire n_731;
wire n_755;
wire n_931;
wire n_1021;
wire n_527;
wire n_683;
wire n_811;
wire n_474;
wire n_1207;
wire n_312;
wire n_1368;
wire n_958;
wire n_1250;
wire n_1137;
wire n_880;
wire n_889;
wire n_589;
wire n_1310;
wire n_819;
wire n_1363;
wire n_1334;
wire n_767;
wire n_1314;
wire n_600;
wire n_964;
wire n_831;
wire n_477;
wire n_954;
wire n_864;
wire n_1110;
wire n_399;
wire n_1372;
wire n_505;
wire n_319;
wire n_1339;
wire n_537;
wire n_311;
wire n_403;
wire n_1080;
wire n_723;
wire n_596;
wire n_546;
wire n_562;
wire n_1141;
wire n_1268;
wire n_386;
wire n_1220;
wire n_556;
wire n_1136;
wire n_1125;
wire n_970;
wire n_642;
wire n_995;
wire n_1159;
wire n_1092;
wire n_441;
wire n_1060;
wire n_444;
wire n_1252;
wire n_1223;
wire n_511;
wire n_1286;
wire n_1053;
wire n_416;
wire n_520;
wire n_418;
wire n_1093;
wire n_775;
wire n_651;
wire n_1153;
wire n_439;
wire n_518;
wire n_1185;
wire n_453;
wire n_914;
wire n_759;
wire n_426;
wire n_317;
wire n_488;
wire n_497;
wire n_773;
wire n_920;
wire n_1374;
wire n_1315;
wire n_1224;
wire n_1135;
wire n_1179;
wire n_1169;
wire n_401;
wire n_324;
wire n_335;
wire n_463;
wire n_1243;
wire n_848;
wire n_1096;
wire n_1091;
wire n_1281;
wire n_1267;
wire n_983;
wire n_427;
wire n_496;
wire n_906;
wire n_688;
wire n_1077;
wire n_351;
wire n_385;
wire n_1323;
wire n_858;
wire n_1331;
wire n_613;
wire n_736;
wire n_501;
wire n_956;
wire n_960;
wire n_663;
wire n_856;
wire n_379;
wire n_778;
wire n_1134;
wire n_410;
wire n_1129;
wire n_554;
wire n_602;
wire n_664;
wire n_435;
wire n_793;
wire n_326;
wire n_587;
wire n_580;
wire n_762;
wire n_1030;
wire n_1202;
wire n_465;
wire n_1079;
wire n_341;
wire n_828;
wire n_607;
wire n_316;
wire n_419;
wire n_1103;
wire n_1203;
wire n_820;
wire n_951;
wire n_725;
wire n_952;
wire n_999;
wire n_358;
wire n_1254;
wire n_368;
wire n_575;
wire n_994;
wire n_732;
wire n_974;
wire n_392;
wire n_724;
wire n_1020;
wire n_1042;
wire n_628;
wire n_1273;
wire n_557;
wire n_349;
wire n_617;
wire n_845;
wire n_807;
wire n_1036;
wire n_1138;
wire n_1275;
wire n_485;
wire n_443;
wire n_892;
wire n_768;
wire n_421;
wire n_1095;
wire n_597;
wire n_1270;
wire n_1187;
wire n_610;
wire n_1024;
wire n_517;
wire n_667;
wire n_1206;
wire n_621;
wire n_1037;
wire n_1279;
wire n_1115;
wire n_750;
wire n_901;
wire n_468;
wire n_923;
wire n_504;
wire n_1015;
wire n_466;
wire n_1057;
wire n_603;
wire n_991;
wire n_1126;
wire n_340;
wire n_710;
wire n_1108;
wire n_1182;
wire n_1298;
wire n_785;
wire n_746;
wire n_609;
wire n_1356;
wire n_1168;
wire n_1216;
wire n_1320;
wire n_1316;
wire n_1287;
wire n_380;
wire n_1190;
wire n_397;
wire n_1262;
wire n_1213;
wire n_1350;
wire n_1272;
wire n_782;
wire n_490;
wire n_809;
wire n_1043;
wire n_986;
wire n_1081;
wire n_402;
wire n_352;
wire n_800;
wire n_1084;
wire n_1171;
wire n_460;
wire n_1361;
wire n_662;
wire n_374;
wire n_1152;
wire n_450;
wire n_921;
wire n_1346;
wire n_711;
wire n_579;
wire n_1352;
wire n_937;
wire n_370;
wire n_650;
wire n_1046;
wire n_1145;
wire n_330;
wire n_1121;
wire n_1102;
wire n_972;
wire n_456;
wire n_1332;
wire n_313;
wire n_624;
wire n_962;
wire n_1041;
wire n_565;
wire n_356;
wire n_936;
wire n_1288;
wire n_1186;
wire n_1062;
wire n_885;
wire n_896;
wire n_654;
wire n_411;
wire n_1222;
wire n_599;
wire n_776;
wire n_321;
wire n_482;
wire n_934;
wire n_420;
wire n_1341;
wire n_394;
wire n_942;
wire n_543;
wire n_1271;
wire n_1355;
wire n_1225;
wire n_325;
wire n_804;
wire n_464;
wire n_533;
wire n_806;
wire n_879;
wire n_959;
wire n_584;
wire n_1343;
wire n_548;
wire n_833;
wire n_523;
wire n_1319;
wire n_707;
wire n_345;
wire n_799;
wire n_1155;
wire n_787;
wire n_1146;
wire n_1086;
wire n_1066;
wire n_1282;
wire n_550;
wire n_652;
wire n_560;
wire n_1321;
wire n_1241;
wire n_569;
wire n_737;
wire n_1318;
wire n_1235;
wire n_1229;
wire n_306;
wire n_1292;
wire n_1373;
wire n_346;
wire n_1029;
wire n_790;
wire n_1210;
wire n_1248;
wire n_902;
wire n_333;
wire n_1047;
wire n_431;
wire n_459;
wire n_1269;
wire n_502;
wire n_672;
wire n_1257;
wire n_1375;
wire n_655;
wire n_706;
wire n_1045;
wire n_786;
wire n_1236;
wire n_834;
wire n_743;
wire n_766;
wire n_430;
wire n_1325;
wire n_1002;
wire n_545;
wire n_489;
wire n_1019;
wire n_636;
wire n_729;
wire n_876;
wire n_774;
wire n_1337;
wire n_660;
wire n_438;
wire n_1360;
wire n_1200;
wire n_479;
wire n_1353;
wire n_869;
wire n_1154;
wire n_1113;
wire n_646;
wire n_528;
wire n_391;
wire n_1098;
wire n_1329;
wire n_817;
wire n_897;
wire n_846;
wire n_841;
wire n_1001;
wire n_508;
wire n_1050;
wire n_1177;
wire n_332;
wire n_1150;
wire n_398;
wire n_1191;
wire n_566;
wire n_1023;
wire n_1076;
wire n_1118;
wire n_1007;
wire n_855;
wire n_591;
wire n_853;
wire n_440;
wire n_695;
wire n_875;
wire n_367;
wire n_680;
wire n_661;
wire n_1256;
wire n_671;
wire n_933;
wire n_740;
wire n_703;
wire n_978;
wire n_384;
wire n_1291;
wire n_1217;
wire n_751;
wire n_749;
wire n_310;
wire n_1324;
wire n_969;
wire n_988;
wire n_1065;
wire n_1255;
wire n_568;
wire n_1204;
wire n_823;
wire n_1132;
wire n_643;
wire n_1074;
wire n_698;
wire n_1327;
wire n_1326;
wire n_739;
wire n_400;
wire n_955;
wire n_337;
wire n_1338;
wire n_1097;
wire n_935;
wire n_781;
wire n_789;
wire n_1130;
wire n_573;
wire n_769;
wire n_676;
wire n_327;
wire n_1120;
wire n_832;
wire n_555;
wire n_814;
wire n_389;
wire n_669;
wire n_747;
wire n_1105;
wire n_721;
wire n_742;
wire n_535;
wire n_691;
wire n_372;
wire n_314;
wire n_378;
wire n_1196;
wire n_377;
wire n_863;
wire n_601;
wire n_338;
wire n_1283;
wire n_918;
wire n_748;
wire n_506;
wire n_1114;
wire n_763;
wire n_1147;
wire n_360;
wire n_957;
wire n_895;
wire n_866;
wire n_1227;
wire n_387;
wire n_452;
wire n_744;
wire n_971;
wire n_946;
wire n_344;
wire n_761;
wire n_1303;
wire n_1205;
wire n_1258;
wire n_1173;
wire n_525;
wire n_1116;
wire n_611;
wire n_1219;
wire n_1174;
wire n_1016;
wire n_1347;
wire n_795;
wire n_1221;
wire n_1245;
wire n_838;
wire n_647;
wire n_844;
wire n_448;
wire n_1017;
wire n_1083;
wire n_445;
wire n_930;
wire n_888;
wire n_1112;
wire n_910;
wire n_911;
wire n_653;
wire n_752;
wire n_908;
wire n_944;
wire n_576;
wire n_1028;
wire n_472;
wire n_414;
wire n_563;
wire n_1011;
wire n_1215;
wire n_839;
wire n_708;
wire n_668;
wire n_626;
wire n_990;
wire n_779;
wire n_1104;
wire n_854;
wire n_1058;
wire n_498;
wire n_1122;
wire n_870;
wire n_904;
wire n_1253;
wire n_709;
wire n_1266;
wire n_366;
wire n_1109;
wire n_712;
wire n_348;
wire n_1276;
wire n_376;
wire n_390;
wire n_1148;
wire n_334;
wire n_1161;
wire n_1085;
wire n_1239;
wire n_771;
wire n_470;
wire n_924;
wire n_475;
wire n_492;
wire n_1149;
wire n_1184;
wire n_719;
wire n_455;
wire n_363;
wire n_1090;
wire n_592;
wire n_829;
wire n_1156;
wire n_1362;
wire n_393;
wire n_984;
wire n_503;
wire n_868;
wire n_859;
wire n_570;
wire n_406;
wire n_735;
wire n_878;
wire n_620;
wire n_519;
wire n_307;
wire n_469;
wire n_1218;
wire n_500;
wire n_981;
wire n_714;
wire n_1349;
wire n_1144;
wire n_357;
wire n_985;
wire n_481;
wire n_997;
wire n_1301;
wire n_802;
wire n_561;
wire n_980;
wire n_1306;
wire n_1198;
wire n_436;
wire n_409;
wire n_1244;
wire n_756;
wire n_810;
wire n_1133;
wire n_635;
wire n_1194;
wire n_1051;
wire n_583;
wire n_1039;
wire n_1034;
wire n_1158;
wire n_754;
wire n_941;
wire n_975;
wire n_1031;
wire n_1305;
wire n_553;
wire n_849;
wire n_753;
wire n_467;
wire n_359;
wire n_973;
wire n_1055;
wire n_582;
wire n_861;
wire n_857;
wire n_967;
wire n_571;
wire n_404;
wire n_679;
wire n_633;
wire n_1170;
wire n_665;
wire n_588;
wire n_1260;
wire n_308;
wire n_309;
wire n_1010;
wire n_1040;
wire n_915;
wire n_632;
wire n_1166;
wire n_812;
wire n_1131;
wire n_534;
wire n_1006;
wire n_373;
wire n_730;
wire n_1311;
wire n_670;
wire n_1089;
wire n_1365;
wire n_1242;
wire n_681;
wire n_1226;
wire n_1274;
wire n_412;
wire n_640;
wire n_1322;
wire n_965;
wire n_339;
wire n_784;
wire n_315;
wire n_434;
wire n_1059;
wire n_1197;
wire n_422;
wire n_722;
wire n_862;
wire n_540;
wire n_457;
wire n_364;
wire n_629;
wire n_900;
wire n_531;
wire n_827;
wire n_361;
wire n_1025;
wire n_336;
wire n_1013;
wire n_1259;
wire n_649;
wire n_1240;

CKINVDCx5p33_ASAP7_75t_R g305 ( 
.A(n_42),
.Y(n_305)
);

INVx2_ASAP7_75t_L g306 ( 
.A(n_22),
.Y(n_306)
);

INVx2_ASAP7_75t_L g307 ( 
.A(n_253),
.Y(n_307)
);

CKINVDCx5p33_ASAP7_75t_R g308 ( 
.A(n_29),
.Y(n_308)
);

CKINVDCx5p33_ASAP7_75t_R g309 ( 
.A(n_153),
.Y(n_309)
);

HB1xp67_ASAP7_75t_L g310 ( 
.A(n_220),
.Y(n_310)
);

CKINVDCx5p33_ASAP7_75t_R g311 ( 
.A(n_122),
.Y(n_311)
);

INVx2_ASAP7_75t_L g312 ( 
.A(n_302),
.Y(n_312)
);

CKINVDCx5p33_ASAP7_75t_R g313 ( 
.A(n_151),
.Y(n_313)
);

CKINVDCx16_ASAP7_75t_R g314 ( 
.A(n_268),
.Y(n_314)
);

CKINVDCx5p33_ASAP7_75t_R g315 ( 
.A(n_58),
.Y(n_315)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_275),
.Y(n_316)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_189),
.Y(n_317)
);

CKINVDCx5p33_ASAP7_75t_R g318 ( 
.A(n_182),
.Y(n_318)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_101),
.Y(n_319)
);

CKINVDCx5p33_ASAP7_75t_R g320 ( 
.A(n_121),
.Y(n_320)
);

CKINVDCx5p33_ASAP7_75t_R g321 ( 
.A(n_156),
.Y(n_321)
);

BUFx2_ASAP7_75t_L g322 ( 
.A(n_34),
.Y(n_322)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_173),
.Y(n_323)
);

CKINVDCx5p33_ASAP7_75t_R g324 ( 
.A(n_254),
.Y(n_324)
);

BUFx3_ASAP7_75t_L g325 ( 
.A(n_186),
.Y(n_325)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_201),
.Y(n_326)
);

CKINVDCx5p33_ASAP7_75t_R g327 ( 
.A(n_12),
.Y(n_327)
);

CKINVDCx5p33_ASAP7_75t_R g328 ( 
.A(n_240),
.Y(n_328)
);

INVx2_ASAP7_75t_L g329 ( 
.A(n_300),
.Y(n_329)
);

INVx1_ASAP7_75t_SL g330 ( 
.A(n_276),
.Y(n_330)
);

CKINVDCx5p33_ASAP7_75t_R g331 ( 
.A(n_175),
.Y(n_331)
);

INVx2_ASAP7_75t_L g332 ( 
.A(n_13),
.Y(n_332)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_228),
.Y(n_333)
);

CKINVDCx5p33_ASAP7_75t_R g334 ( 
.A(n_161),
.Y(n_334)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_67),
.Y(n_335)
);

CKINVDCx5p33_ASAP7_75t_R g336 ( 
.A(n_249),
.Y(n_336)
);

CKINVDCx5p33_ASAP7_75t_R g337 ( 
.A(n_279),
.Y(n_337)
);

CKINVDCx20_ASAP7_75t_R g338 ( 
.A(n_54),
.Y(n_338)
);

INVx2_ASAP7_75t_L g339 ( 
.A(n_208),
.Y(n_339)
);

BUFx6f_ASAP7_75t_L g340 ( 
.A(n_77),
.Y(n_340)
);

INVx2_ASAP7_75t_L g341 ( 
.A(n_71),
.Y(n_341)
);

INVx1_ASAP7_75t_L g342 ( 
.A(n_17),
.Y(n_342)
);

CKINVDCx5p33_ASAP7_75t_R g343 ( 
.A(n_277),
.Y(n_343)
);

CKINVDCx20_ASAP7_75t_R g344 ( 
.A(n_30),
.Y(n_344)
);

CKINVDCx5p33_ASAP7_75t_R g345 ( 
.A(n_165),
.Y(n_345)
);

INVx1_ASAP7_75t_L g346 ( 
.A(n_293),
.Y(n_346)
);

CKINVDCx5p33_ASAP7_75t_R g347 ( 
.A(n_140),
.Y(n_347)
);

INVxp67_ASAP7_75t_L g348 ( 
.A(n_114),
.Y(n_348)
);

CKINVDCx5p33_ASAP7_75t_R g349 ( 
.A(n_123),
.Y(n_349)
);

CKINVDCx5p33_ASAP7_75t_R g350 ( 
.A(n_143),
.Y(n_350)
);

CKINVDCx5p33_ASAP7_75t_R g351 ( 
.A(n_0),
.Y(n_351)
);

CKINVDCx5p33_ASAP7_75t_R g352 ( 
.A(n_272),
.Y(n_352)
);

CKINVDCx20_ASAP7_75t_R g353 ( 
.A(n_296),
.Y(n_353)
);

INVx1_ASAP7_75t_L g354 ( 
.A(n_200),
.Y(n_354)
);

INVx1_ASAP7_75t_L g355 ( 
.A(n_50),
.Y(n_355)
);

CKINVDCx5p33_ASAP7_75t_R g356 ( 
.A(n_292),
.Y(n_356)
);

INVx2_ASAP7_75t_L g357 ( 
.A(n_205),
.Y(n_357)
);

INVxp33_ASAP7_75t_SL g358 ( 
.A(n_93),
.Y(n_358)
);

CKINVDCx5p33_ASAP7_75t_R g359 ( 
.A(n_280),
.Y(n_359)
);

CKINVDCx5p33_ASAP7_75t_R g360 ( 
.A(n_301),
.Y(n_360)
);

CKINVDCx5p33_ASAP7_75t_R g361 ( 
.A(n_187),
.Y(n_361)
);

INVx1_ASAP7_75t_L g362 ( 
.A(n_40),
.Y(n_362)
);

CKINVDCx20_ASAP7_75t_R g363 ( 
.A(n_96),
.Y(n_363)
);

BUFx10_ASAP7_75t_L g364 ( 
.A(n_60),
.Y(n_364)
);

CKINVDCx5p33_ASAP7_75t_R g365 ( 
.A(n_204),
.Y(n_365)
);

NOR2xp67_ASAP7_75t_L g366 ( 
.A(n_181),
.B(n_243),
.Y(n_366)
);

CKINVDCx5p33_ASAP7_75t_R g367 ( 
.A(n_290),
.Y(n_367)
);

CKINVDCx5p33_ASAP7_75t_R g368 ( 
.A(n_124),
.Y(n_368)
);

INVx2_ASAP7_75t_L g369 ( 
.A(n_111),
.Y(n_369)
);

INVx1_ASAP7_75t_SL g370 ( 
.A(n_66),
.Y(n_370)
);

INVx2_ASAP7_75t_L g371 ( 
.A(n_285),
.Y(n_371)
);

INVx1_ASAP7_75t_L g372 ( 
.A(n_0),
.Y(n_372)
);

CKINVDCx5p33_ASAP7_75t_R g373 ( 
.A(n_82),
.Y(n_373)
);

CKINVDCx16_ASAP7_75t_R g374 ( 
.A(n_85),
.Y(n_374)
);

CKINVDCx5p33_ASAP7_75t_R g375 ( 
.A(n_263),
.Y(n_375)
);

CKINVDCx5p33_ASAP7_75t_R g376 ( 
.A(n_163),
.Y(n_376)
);

CKINVDCx5p33_ASAP7_75t_R g377 ( 
.A(n_86),
.Y(n_377)
);

INVx1_ASAP7_75t_L g378 ( 
.A(n_196),
.Y(n_378)
);

INVx1_ASAP7_75t_L g379 ( 
.A(n_230),
.Y(n_379)
);

CKINVDCx5p33_ASAP7_75t_R g380 ( 
.A(n_133),
.Y(n_380)
);

INVx1_ASAP7_75t_L g381 ( 
.A(n_256),
.Y(n_381)
);

CKINVDCx5p33_ASAP7_75t_R g382 ( 
.A(n_248),
.Y(n_382)
);

CKINVDCx16_ASAP7_75t_R g383 ( 
.A(n_144),
.Y(n_383)
);

INVx1_ASAP7_75t_L g384 ( 
.A(n_148),
.Y(n_384)
);

CKINVDCx5p33_ASAP7_75t_R g385 ( 
.A(n_110),
.Y(n_385)
);

INVx1_ASAP7_75t_L g386 ( 
.A(n_102),
.Y(n_386)
);

NAND2xp5_ASAP7_75t_L g387 ( 
.A(n_74),
.B(n_231),
.Y(n_387)
);

CKINVDCx5p33_ASAP7_75t_R g388 ( 
.A(n_190),
.Y(n_388)
);

CKINVDCx5p33_ASAP7_75t_R g389 ( 
.A(n_297),
.Y(n_389)
);

CKINVDCx5p33_ASAP7_75t_R g390 ( 
.A(n_198),
.Y(n_390)
);

INVx3_ASAP7_75t_L g391 ( 
.A(n_89),
.Y(n_391)
);

INVx2_ASAP7_75t_L g392 ( 
.A(n_49),
.Y(n_392)
);

CKINVDCx5p33_ASAP7_75t_R g393 ( 
.A(n_218),
.Y(n_393)
);

CKINVDCx5p33_ASAP7_75t_R g394 ( 
.A(n_19),
.Y(n_394)
);

INVx1_ASAP7_75t_L g395 ( 
.A(n_299),
.Y(n_395)
);

CKINVDCx5p33_ASAP7_75t_R g396 ( 
.A(n_91),
.Y(n_396)
);

CKINVDCx5p33_ASAP7_75t_R g397 ( 
.A(n_46),
.Y(n_397)
);

CKINVDCx5p33_ASAP7_75t_R g398 ( 
.A(n_295),
.Y(n_398)
);

INVx1_ASAP7_75t_L g399 ( 
.A(n_8),
.Y(n_399)
);

BUFx3_ASAP7_75t_L g400 ( 
.A(n_252),
.Y(n_400)
);

INVx1_ASAP7_75t_L g401 ( 
.A(n_69),
.Y(n_401)
);

HB1xp67_ASAP7_75t_L g402 ( 
.A(n_139),
.Y(n_402)
);

BUFx5_ASAP7_75t_L g403 ( 
.A(n_131),
.Y(n_403)
);

CKINVDCx5p33_ASAP7_75t_R g404 ( 
.A(n_168),
.Y(n_404)
);

INVx2_ASAP7_75t_L g405 ( 
.A(n_206),
.Y(n_405)
);

BUFx2_ASAP7_75t_L g406 ( 
.A(n_63),
.Y(n_406)
);

INVx1_ASAP7_75t_L g407 ( 
.A(n_132),
.Y(n_407)
);

INVx1_ASAP7_75t_L g408 ( 
.A(n_13),
.Y(n_408)
);

INVx1_ASAP7_75t_L g409 ( 
.A(n_194),
.Y(n_409)
);

INVx1_ASAP7_75t_L g410 ( 
.A(n_241),
.Y(n_410)
);

INVx1_ASAP7_75t_L g411 ( 
.A(n_53),
.Y(n_411)
);

CKINVDCx5p33_ASAP7_75t_R g412 ( 
.A(n_209),
.Y(n_412)
);

HB1xp67_ASAP7_75t_L g413 ( 
.A(n_213),
.Y(n_413)
);

BUFx10_ASAP7_75t_L g414 ( 
.A(n_4),
.Y(n_414)
);

CKINVDCx5p33_ASAP7_75t_R g415 ( 
.A(n_291),
.Y(n_415)
);

BUFx10_ASAP7_75t_L g416 ( 
.A(n_180),
.Y(n_416)
);

CKINVDCx5p33_ASAP7_75t_R g417 ( 
.A(n_108),
.Y(n_417)
);

CKINVDCx5p33_ASAP7_75t_R g418 ( 
.A(n_282),
.Y(n_418)
);

INVx1_ASAP7_75t_SL g419 ( 
.A(n_47),
.Y(n_419)
);

CKINVDCx5p33_ASAP7_75t_R g420 ( 
.A(n_141),
.Y(n_420)
);

CKINVDCx20_ASAP7_75t_R g421 ( 
.A(n_48),
.Y(n_421)
);

INVx1_ASAP7_75t_L g422 ( 
.A(n_298),
.Y(n_422)
);

CKINVDCx5p33_ASAP7_75t_R g423 ( 
.A(n_117),
.Y(n_423)
);

INVx1_ASAP7_75t_SL g424 ( 
.A(n_6),
.Y(n_424)
);

INVx1_ASAP7_75t_L g425 ( 
.A(n_45),
.Y(n_425)
);

INVx1_ASAP7_75t_L g426 ( 
.A(n_229),
.Y(n_426)
);

CKINVDCx5p33_ASAP7_75t_R g427 ( 
.A(n_179),
.Y(n_427)
);

CKINVDCx5p33_ASAP7_75t_R g428 ( 
.A(n_250),
.Y(n_428)
);

CKINVDCx5p33_ASAP7_75t_R g429 ( 
.A(n_2),
.Y(n_429)
);

INVx1_ASAP7_75t_L g430 ( 
.A(n_245),
.Y(n_430)
);

CKINVDCx5p33_ASAP7_75t_R g431 ( 
.A(n_171),
.Y(n_431)
);

CKINVDCx20_ASAP7_75t_R g432 ( 
.A(n_211),
.Y(n_432)
);

INVx1_ASAP7_75t_SL g433 ( 
.A(n_21),
.Y(n_433)
);

INVx1_ASAP7_75t_L g434 ( 
.A(n_83),
.Y(n_434)
);

INVx1_ASAP7_75t_L g435 ( 
.A(n_119),
.Y(n_435)
);

INVxp67_ASAP7_75t_L g436 ( 
.A(n_159),
.Y(n_436)
);

CKINVDCx5p33_ASAP7_75t_R g437 ( 
.A(n_2),
.Y(n_437)
);

CKINVDCx5p33_ASAP7_75t_R g438 ( 
.A(n_216),
.Y(n_438)
);

INVx1_ASAP7_75t_L g439 ( 
.A(n_146),
.Y(n_439)
);

CKINVDCx5p33_ASAP7_75t_R g440 ( 
.A(n_103),
.Y(n_440)
);

BUFx3_ASAP7_75t_L g441 ( 
.A(n_149),
.Y(n_441)
);

INVx1_ASAP7_75t_L g442 ( 
.A(n_262),
.Y(n_442)
);

INVx2_ASAP7_75t_SL g443 ( 
.A(n_162),
.Y(n_443)
);

INVx1_ASAP7_75t_L g444 ( 
.A(n_126),
.Y(n_444)
);

BUFx10_ASAP7_75t_L g445 ( 
.A(n_185),
.Y(n_445)
);

INVx2_ASAP7_75t_L g446 ( 
.A(n_287),
.Y(n_446)
);

CKINVDCx5p33_ASAP7_75t_R g447 ( 
.A(n_5),
.Y(n_447)
);

CKINVDCx5p33_ASAP7_75t_R g448 ( 
.A(n_169),
.Y(n_448)
);

INVx1_ASAP7_75t_L g449 ( 
.A(n_43),
.Y(n_449)
);

CKINVDCx20_ASAP7_75t_R g450 ( 
.A(n_157),
.Y(n_450)
);

INVx1_ASAP7_75t_L g451 ( 
.A(n_202),
.Y(n_451)
);

CKINVDCx5p33_ASAP7_75t_R g452 ( 
.A(n_81),
.Y(n_452)
);

INVx1_ASAP7_75t_L g453 ( 
.A(n_283),
.Y(n_453)
);

INVx1_ASAP7_75t_L g454 ( 
.A(n_274),
.Y(n_454)
);

INVx2_ASAP7_75t_L g455 ( 
.A(n_155),
.Y(n_455)
);

CKINVDCx5p33_ASAP7_75t_R g456 ( 
.A(n_113),
.Y(n_456)
);

CKINVDCx5p33_ASAP7_75t_R g457 ( 
.A(n_197),
.Y(n_457)
);

INVx2_ASAP7_75t_L g458 ( 
.A(n_183),
.Y(n_458)
);

CKINVDCx5p33_ASAP7_75t_R g459 ( 
.A(n_260),
.Y(n_459)
);

INVx1_ASAP7_75t_L g460 ( 
.A(n_23),
.Y(n_460)
);

INVx2_ASAP7_75t_L g461 ( 
.A(n_176),
.Y(n_461)
);

INVx1_ASAP7_75t_L g462 ( 
.A(n_238),
.Y(n_462)
);

CKINVDCx5p33_ASAP7_75t_R g463 ( 
.A(n_184),
.Y(n_463)
);

CKINVDCx20_ASAP7_75t_R g464 ( 
.A(n_214),
.Y(n_464)
);

CKINVDCx5p33_ASAP7_75t_R g465 ( 
.A(n_304),
.Y(n_465)
);

HB1xp67_ASAP7_75t_L g466 ( 
.A(n_212),
.Y(n_466)
);

CKINVDCx5p33_ASAP7_75t_R g467 ( 
.A(n_160),
.Y(n_467)
);

INVx2_ASAP7_75t_SL g468 ( 
.A(n_278),
.Y(n_468)
);

CKINVDCx5p33_ASAP7_75t_R g469 ( 
.A(n_62),
.Y(n_469)
);

BUFx6f_ASAP7_75t_L g470 ( 
.A(n_104),
.Y(n_470)
);

CKINVDCx5p33_ASAP7_75t_R g471 ( 
.A(n_137),
.Y(n_471)
);

BUFx3_ASAP7_75t_L g472 ( 
.A(n_147),
.Y(n_472)
);

INVx1_ASAP7_75t_L g473 ( 
.A(n_100),
.Y(n_473)
);

CKINVDCx5p33_ASAP7_75t_R g474 ( 
.A(n_172),
.Y(n_474)
);

CKINVDCx5p33_ASAP7_75t_R g475 ( 
.A(n_264),
.Y(n_475)
);

BUFx8_ASAP7_75t_SL g476 ( 
.A(n_289),
.Y(n_476)
);

CKINVDCx5p33_ASAP7_75t_R g477 ( 
.A(n_135),
.Y(n_477)
);

BUFx6f_ASAP7_75t_L g478 ( 
.A(n_36),
.Y(n_478)
);

BUFx6f_ASAP7_75t_L g479 ( 
.A(n_281),
.Y(n_479)
);

BUFx6f_ASAP7_75t_L g480 ( 
.A(n_35),
.Y(n_480)
);

CKINVDCx5p33_ASAP7_75t_R g481 ( 
.A(n_115),
.Y(n_481)
);

CKINVDCx20_ASAP7_75t_R g482 ( 
.A(n_78),
.Y(n_482)
);

CKINVDCx5p33_ASAP7_75t_R g483 ( 
.A(n_193),
.Y(n_483)
);

CKINVDCx5p33_ASAP7_75t_R g484 ( 
.A(n_188),
.Y(n_484)
);

CKINVDCx5p33_ASAP7_75t_R g485 ( 
.A(n_270),
.Y(n_485)
);

CKINVDCx5p33_ASAP7_75t_R g486 ( 
.A(n_136),
.Y(n_486)
);

INVx2_ASAP7_75t_L g487 ( 
.A(n_284),
.Y(n_487)
);

INVx1_ASAP7_75t_L g488 ( 
.A(n_6),
.Y(n_488)
);

CKINVDCx5p33_ASAP7_75t_R g489 ( 
.A(n_203),
.Y(n_489)
);

CKINVDCx5p33_ASAP7_75t_R g490 ( 
.A(n_224),
.Y(n_490)
);

CKINVDCx5p33_ASAP7_75t_R g491 ( 
.A(n_80),
.Y(n_491)
);

BUFx10_ASAP7_75t_L g492 ( 
.A(n_177),
.Y(n_492)
);

INVx1_ASAP7_75t_L g493 ( 
.A(n_134),
.Y(n_493)
);

CKINVDCx5p33_ASAP7_75t_R g494 ( 
.A(n_226),
.Y(n_494)
);

CKINVDCx5p33_ASAP7_75t_R g495 ( 
.A(n_35),
.Y(n_495)
);

INVx1_ASAP7_75t_L g496 ( 
.A(n_273),
.Y(n_496)
);

BUFx6f_ASAP7_75t_L g497 ( 
.A(n_99),
.Y(n_497)
);

CKINVDCx5p33_ASAP7_75t_R g498 ( 
.A(n_120),
.Y(n_498)
);

INVx2_ASAP7_75t_L g499 ( 
.A(n_44),
.Y(n_499)
);

CKINVDCx5p33_ASAP7_75t_R g500 ( 
.A(n_90),
.Y(n_500)
);

NOR2xp67_ASAP7_75t_L g501 ( 
.A(n_269),
.B(n_178),
.Y(n_501)
);

CKINVDCx5p33_ASAP7_75t_R g502 ( 
.A(n_52),
.Y(n_502)
);

INVx2_ASAP7_75t_L g503 ( 
.A(n_225),
.Y(n_503)
);

INVx1_ASAP7_75t_L g504 ( 
.A(n_84),
.Y(n_504)
);

INVx1_ASAP7_75t_L g505 ( 
.A(n_70),
.Y(n_505)
);

BUFx6f_ASAP7_75t_L g506 ( 
.A(n_1),
.Y(n_506)
);

CKINVDCx5p33_ASAP7_75t_R g507 ( 
.A(n_267),
.Y(n_507)
);

INVx1_ASAP7_75t_L g508 ( 
.A(n_255),
.Y(n_508)
);

INVx1_ASAP7_75t_L g509 ( 
.A(n_28),
.Y(n_509)
);

CKINVDCx5p33_ASAP7_75t_R g510 ( 
.A(n_38),
.Y(n_510)
);

BUFx10_ASAP7_75t_L g511 ( 
.A(n_39),
.Y(n_511)
);

CKINVDCx20_ASAP7_75t_R g512 ( 
.A(n_167),
.Y(n_512)
);

INVx1_ASAP7_75t_L g513 ( 
.A(n_303),
.Y(n_513)
);

BUFx10_ASAP7_75t_L g514 ( 
.A(n_19),
.Y(n_514)
);

CKINVDCx5p33_ASAP7_75t_R g515 ( 
.A(n_286),
.Y(n_515)
);

CKINVDCx5p33_ASAP7_75t_R g516 ( 
.A(n_207),
.Y(n_516)
);

CKINVDCx5p33_ASAP7_75t_R g517 ( 
.A(n_166),
.Y(n_517)
);

INVx1_ASAP7_75t_L g518 ( 
.A(n_88),
.Y(n_518)
);

INVx1_ASAP7_75t_L g519 ( 
.A(n_174),
.Y(n_519)
);

CKINVDCx5p33_ASAP7_75t_R g520 ( 
.A(n_33),
.Y(n_520)
);

INVx2_ASAP7_75t_SL g521 ( 
.A(n_191),
.Y(n_521)
);

CKINVDCx5p33_ASAP7_75t_R g522 ( 
.A(n_154),
.Y(n_522)
);

INVx1_ASAP7_75t_L g523 ( 
.A(n_145),
.Y(n_523)
);

INVx1_ASAP7_75t_L g524 ( 
.A(n_79),
.Y(n_524)
);

INVx1_ASAP7_75t_SL g525 ( 
.A(n_44),
.Y(n_525)
);

OAI22x1_ASAP7_75t_R g526 ( 
.A1(n_344),
.A2(n_1),
.B1(n_3),
.B2(n_4),
.Y(n_526)
);

NOR2xp33_ASAP7_75t_L g527 ( 
.A(n_310),
.B(n_3),
.Y(n_527)
);

BUFx3_ASAP7_75t_L g528 ( 
.A(n_364),
.Y(n_528)
);

INVx1_ASAP7_75t_L g529 ( 
.A(n_478),
.Y(n_529)
);

BUFx6f_ASAP7_75t_L g530 ( 
.A(n_340),
.Y(n_530)
);

INVx3_ASAP7_75t_L g531 ( 
.A(n_478),
.Y(n_531)
);

INVx3_ASAP7_75t_L g532 ( 
.A(n_478),
.Y(n_532)
);

INVx4_ASAP7_75t_L g533 ( 
.A(n_340),
.Y(n_533)
);

BUFx6f_ASAP7_75t_L g534 ( 
.A(n_340),
.Y(n_534)
);

BUFx2_ASAP7_75t_L g535 ( 
.A(n_322),
.Y(n_535)
);

BUFx6f_ASAP7_75t_L g536 ( 
.A(n_340),
.Y(n_536)
);

BUFx6f_ASAP7_75t_L g537 ( 
.A(n_470),
.Y(n_537)
);

INVx2_ASAP7_75t_L g538 ( 
.A(n_478),
.Y(n_538)
);

AOI22x1_ASAP7_75t_SL g539 ( 
.A1(n_305),
.A2(n_5),
.B1(n_7),
.B2(n_8),
.Y(n_539)
);

AND2x2_ASAP7_75t_L g540 ( 
.A(n_406),
.B(n_7),
.Y(n_540)
);

BUFx2_ASAP7_75t_L g541 ( 
.A(n_308),
.Y(n_541)
);

INVx1_ASAP7_75t_L g542 ( 
.A(n_480),
.Y(n_542)
);

BUFx6f_ASAP7_75t_L g543 ( 
.A(n_470),
.Y(n_543)
);

INVx1_ASAP7_75t_L g544 ( 
.A(n_480),
.Y(n_544)
);

BUFx3_ASAP7_75t_L g545 ( 
.A(n_364),
.Y(n_545)
);

NOR2xp33_ASAP7_75t_SL g546 ( 
.A(n_314),
.B(n_9),
.Y(n_546)
);

INVx1_ASAP7_75t_L g547 ( 
.A(n_480),
.Y(n_547)
);

INVx5_ASAP7_75t_L g548 ( 
.A(n_470),
.Y(n_548)
);

INVx1_ASAP7_75t_SL g549 ( 
.A(n_414),
.Y(n_549)
);

BUFx2_ASAP7_75t_L g550 ( 
.A(n_327),
.Y(n_550)
);

BUFx6f_ASAP7_75t_L g551 ( 
.A(n_470),
.Y(n_551)
);

BUFx3_ASAP7_75t_L g552 ( 
.A(n_416),
.Y(n_552)
);

BUFx2_ASAP7_75t_L g553 ( 
.A(n_351),
.Y(n_553)
);

BUFx6f_ASAP7_75t_L g554 ( 
.A(n_479),
.Y(n_554)
);

OAI22x1_ASAP7_75t_SL g555 ( 
.A1(n_394),
.A2(n_9),
.B1(n_10),
.B2(n_11),
.Y(n_555)
);

INVx3_ASAP7_75t_L g556 ( 
.A(n_506),
.Y(n_556)
);

CKINVDCx5p33_ASAP7_75t_R g557 ( 
.A(n_476),
.Y(n_557)
);

INVx2_ASAP7_75t_L g558 ( 
.A(n_506),
.Y(n_558)
);

BUFx6f_ASAP7_75t_L g559 ( 
.A(n_479),
.Y(n_559)
);

BUFx6f_ASAP7_75t_L g560 ( 
.A(n_479),
.Y(n_560)
);

INVx1_ASAP7_75t_L g561 ( 
.A(n_506),
.Y(n_561)
);

INVx1_ASAP7_75t_L g562 ( 
.A(n_506),
.Y(n_562)
);

AND2x4_ASAP7_75t_L g563 ( 
.A(n_325),
.B(n_10),
.Y(n_563)
);

INVx5_ASAP7_75t_L g564 ( 
.A(n_479),
.Y(n_564)
);

AOI22x1_ASAP7_75t_SL g565 ( 
.A1(n_397),
.A2(n_12),
.B1(n_14),
.B2(n_15),
.Y(n_565)
);

HB1xp67_ASAP7_75t_L g566 ( 
.A(n_429),
.Y(n_566)
);

CKINVDCx5p33_ASAP7_75t_R g567 ( 
.A(n_309),
.Y(n_567)
);

OA21x2_ASAP7_75t_L g568 ( 
.A1(n_316),
.A2(n_14),
.B(n_15),
.Y(n_568)
);

CKINVDCx20_ASAP7_75t_R g569 ( 
.A(n_338),
.Y(n_569)
);

BUFx6f_ASAP7_75t_L g570 ( 
.A(n_497),
.Y(n_570)
);

INVx1_ASAP7_75t_L g571 ( 
.A(n_342),
.Y(n_571)
);

INVx1_ASAP7_75t_L g572 ( 
.A(n_362),
.Y(n_572)
);

INVx5_ASAP7_75t_L g573 ( 
.A(n_497),
.Y(n_573)
);

AND2x4_ASAP7_75t_L g574 ( 
.A(n_400),
.B(n_16),
.Y(n_574)
);

BUFx6f_ASAP7_75t_L g575 ( 
.A(n_497),
.Y(n_575)
);

OAI21x1_ASAP7_75t_L g576 ( 
.A1(n_391),
.A2(n_55),
.B(n_51),
.Y(n_576)
);

INVx5_ASAP7_75t_L g577 ( 
.A(n_497),
.Y(n_577)
);

INVx2_ASAP7_75t_L g578 ( 
.A(n_403),
.Y(n_578)
);

INVx2_ASAP7_75t_L g579 ( 
.A(n_403),
.Y(n_579)
);

INVx1_ASAP7_75t_L g580 ( 
.A(n_372),
.Y(n_580)
);

AND2x4_ASAP7_75t_L g581 ( 
.A(n_441),
.B(n_18),
.Y(n_581)
);

CKINVDCx11_ASAP7_75t_R g582 ( 
.A(n_511),
.Y(n_582)
);

HB1xp67_ASAP7_75t_L g583 ( 
.A(n_437),
.Y(n_583)
);

BUFx8_ASAP7_75t_L g584 ( 
.A(n_306),
.Y(n_584)
);

CKINVDCx16_ASAP7_75t_R g585 ( 
.A(n_374),
.Y(n_585)
);

HB1xp67_ASAP7_75t_L g586 ( 
.A(n_447),
.Y(n_586)
);

BUFx3_ASAP7_75t_L g587 ( 
.A(n_416),
.Y(n_587)
);

INVx2_ASAP7_75t_L g588 ( 
.A(n_403),
.Y(n_588)
);

AND2x6_ASAP7_75t_L g589 ( 
.A(n_391),
.B(n_56),
.Y(n_589)
);

BUFx6f_ASAP7_75t_L g590 ( 
.A(n_472),
.Y(n_590)
);

BUFx6f_ASAP7_75t_L g591 ( 
.A(n_307),
.Y(n_591)
);

INVx1_ASAP7_75t_L g592 ( 
.A(n_399),
.Y(n_592)
);

BUFx6f_ASAP7_75t_L g593 ( 
.A(n_312),
.Y(n_593)
);

INVx1_ASAP7_75t_L g594 ( 
.A(n_408),
.Y(n_594)
);

BUFx12f_ASAP7_75t_L g595 ( 
.A(n_514),
.Y(n_595)
);

BUFx12f_ASAP7_75t_L g596 ( 
.A(n_514),
.Y(n_596)
);

INVx1_ASAP7_75t_L g597 ( 
.A(n_425),
.Y(n_597)
);

BUFx8_ASAP7_75t_SL g598 ( 
.A(n_353),
.Y(n_598)
);

HB1xp67_ASAP7_75t_L g599 ( 
.A(n_495),
.Y(n_599)
);

INVx1_ASAP7_75t_L g600 ( 
.A(n_449),
.Y(n_600)
);

BUFx6f_ASAP7_75t_L g601 ( 
.A(n_329),
.Y(n_601)
);

INVx2_ASAP7_75t_L g602 ( 
.A(n_403),
.Y(n_602)
);

AND2x4_ASAP7_75t_L g603 ( 
.A(n_310),
.B(n_20),
.Y(n_603)
);

INVx2_ASAP7_75t_L g604 ( 
.A(n_403),
.Y(n_604)
);

BUFx6f_ASAP7_75t_L g605 ( 
.A(n_339),
.Y(n_605)
);

AND2x6_ASAP7_75t_L g606 ( 
.A(n_341),
.B(n_57),
.Y(n_606)
);

BUFx6f_ASAP7_75t_L g607 ( 
.A(n_357),
.Y(n_607)
);

BUFx3_ASAP7_75t_L g608 ( 
.A(n_445),
.Y(n_608)
);

INVx3_ASAP7_75t_L g609 ( 
.A(n_332),
.Y(n_609)
);

BUFx8_ASAP7_75t_SL g610 ( 
.A(n_363),
.Y(n_610)
);

INVx2_ASAP7_75t_L g611 ( 
.A(n_403),
.Y(n_611)
);

AND2x6_ASAP7_75t_L g612 ( 
.A(n_369),
.B(n_59),
.Y(n_612)
);

BUFx12f_ASAP7_75t_L g613 ( 
.A(n_492),
.Y(n_613)
);

INVx2_ASAP7_75t_L g614 ( 
.A(n_460),
.Y(n_614)
);

AOI22xp5_ASAP7_75t_L g615 ( 
.A1(n_383),
.A2(n_23),
.B1(n_24),
.B2(n_25),
.Y(n_615)
);

NAND2xp5_ASAP7_75t_L g616 ( 
.A(n_402),
.B(n_24),
.Y(n_616)
);

BUFx8_ASAP7_75t_L g617 ( 
.A(n_499),
.Y(n_617)
);

INVx6_ASAP7_75t_L g618 ( 
.A(n_492),
.Y(n_618)
);

CKINVDCx5p33_ASAP7_75t_R g619 ( 
.A(n_311),
.Y(n_619)
);

INVx1_ASAP7_75t_L g620 ( 
.A(n_488),
.Y(n_620)
);

BUFx6f_ASAP7_75t_L g621 ( 
.A(n_371),
.Y(n_621)
);

INVx2_ASAP7_75t_L g622 ( 
.A(n_509),
.Y(n_622)
);

INVx5_ASAP7_75t_L g623 ( 
.A(n_443),
.Y(n_623)
);

BUFx6f_ASAP7_75t_L g624 ( 
.A(n_392),
.Y(n_624)
);

AND2x2_ASAP7_75t_L g625 ( 
.A(n_402),
.B(n_25),
.Y(n_625)
);

BUFx3_ASAP7_75t_L g626 ( 
.A(n_313),
.Y(n_626)
);

INVx1_ASAP7_75t_L g627 ( 
.A(n_317),
.Y(n_627)
);

OAI21x1_ASAP7_75t_L g628 ( 
.A1(n_405),
.A2(n_64),
.B(n_61),
.Y(n_628)
);

INVx3_ASAP7_75t_L g629 ( 
.A(n_510),
.Y(n_629)
);

INVx1_ASAP7_75t_L g630 ( 
.A(n_319),
.Y(n_630)
);

BUFx8_ASAP7_75t_SL g631 ( 
.A(n_421),
.Y(n_631)
);

OAI21x1_ASAP7_75t_L g632 ( 
.A1(n_446),
.A2(n_68),
.B(n_65),
.Y(n_632)
);

INVx1_ASAP7_75t_L g633 ( 
.A(n_323),
.Y(n_633)
);

INVx5_ASAP7_75t_L g634 ( 
.A(n_468),
.Y(n_634)
);

BUFx6f_ASAP7_75t_L g635 ( 
.A(n_455),
.Y(n_635)
);

NAND2xp5_ASAP7_75t_L g636 ( 
.A(n_413),
.B(n_26),
.Y(n_636)
);

HB1xp67_ASAP7_75t_L g637 ( 
.A(n_520),
.Y(n_637)
);

AND2x4_ASAP7_75t_L g638 ( 
.A(n_466),
.B(n_27),
.Y(n_638)
);

BUFx12f_ASAP7_75t_L g639 ( 
.A(n_315),
.Y(n_639)
);

INVx1_ASAP7_75t_L g640 ( 
.A(n_326),
.Y(n_640)
);

BUFx6f_ASAP7_75t_L g641 ( 
.A(n_458),
.Y(n_641)
);

AND2x4_ASAP7_75t_L g642 ( 
.A(n_466),
.B(n_28),
.Y(n_642)
);

INVx5_ASAP7_75t_L g643 ( 
.A(n_521),
.Y(n_643)
);

INVx5_ASAP7_75t_L g644 ( 
.A(n_461),
.Y(n_644)
);

AOI22xp5_ASAP7_75t_L g645 ( 
.A1(n_358),
.A2(n_30),
.B1(n_31),
.B2(n_32),
.Y(n_645)
);

INVx2_ASAP7_75t_L g646 ( 
.A(n_333),
.Y(n_646)
);

INVxp67_ASAP7_75t_L g647 ( 
.A(n_419),
.Y(n_647)
);

INVx2_ASAP7_75t_L g648 ( 
.A(n_335),
.Y(n_648)
);

NAND2xp5_ASAP7_75t_L g649 ( 
.A(n_487),
.B(n_31),
.Y(n_649)
);

INVx1_ASAP7_75t_L g650 ( 
.A(n_346),
.Y(n_650)
);

INVx1_ASAP7_75t_L g651 ( 
.A(n_354),
.Y(n_651)
);

BUFx3_ASAP7_75t_L g652 ( 
.A(n_318),
.Y(n_652)
);

INVx2_ASAP7_75t_L g653 ( 
.A(n_355),
.Y(n_653)
);

INVx5_ASAP7_75t_L g654 ( 
.A(n_503),
.Y(n_654)
);

INVx2_ASAP7_75t_L g655 ( 
.A(n_378),
.Y(n_655)
);

INVx2_ASAP7_75t_L g656 ( 
.A(n_379),
.Y(n_656)
);

INVx1_ASAP7_75t_L g657 ( 
.A(n_381),
.Y(n_657)
);

BUFx3_ASAP7_75t_L g658 ( 
.A(n_320),
.Y(n_658)
);

OAI21x1_ASAP7_75t_L g659 ( 
.A1(n_387),
.A2(n_73),
.B(n_72),
.Y(n_659)
);

BUFx6f_ASAP7_75t_L g660 ( 
.A(n_384),
.Y(n_660)
);

INVx2_ASAP7_75t_L g661 ( 
.A(n_386),
.Y(n_661)
);

INVx1_ASAP7_75t_L g662 ( 
.A(n_395),
.Y(n_662)
);

OAI21x1_ASAP7_75t_L g663 ( 
.A1(n_401),
.A2(n_409),
.B(n_407),
.Y(n_663)
);

INVx1_ASAP7_75t_L g664 ( 
.A(n_410),
.Y(n_664)
);

BUFx6f_ASAP7_75t_L g665 ( 
.A(n_411),
.Y(n_665)
);

BUFx12f_ASAP7_75t_L g666 ( 
.A(n_321),
.Y(n_666)
);

INVx2_ASAP7_75t_L g667 ( 
.A(n_422),
.Y(n_667)
);

AOI22xp5_ASAP7_75t_L g668 ( 
.A1(n_424),
.A2(n_37),
.B1(n_38),
.B2(n_39),
.Y(n_668)
);

AND2x2_ASAP7_75t_L g669 ( 
.A(n_525),
.B(n_433),
.Y(n_669)
);

INVx2_ASAP7_75t_L g670 ( 
.A(n_426),
.Y(n_670)
);

INVx1_ASAP7_75t_L g671 ( 
.A(n_430),
.Y(n_671)
);

AND2x2_ASAP7_75t_L g672 ( 
.A(n_566),
.B(n_330),
.Y(n_672)
);

INVx3_ASAP7_75t_L g673 ( 
.A(n_531),
.Y(n_673)
);

CKINVDCx5p33_ASAP7_75t_R g674 ( 
.A(n_598),
.Y(n_674)
);

BUFx2_ASAP7_75t_L g675 ( 
.A(n_647),
.Y(n_675)
);

BUFx3_ASAP7_75t_L g676 ( 
.A(n_590),
.Y(n_676)
);

CKINVDCx5p33_ASAP7_75t_R g677 ( 
.A(n_610),
.Y(n_677)
);

INVx2_ASAP7_75t_L g678 ( 
.A(n_538),
.Y(n_678)
);

INVx4_ASAP7_75t_L g679 ( 
.A(n_567),
.Y(n_679)
);

CKINVDCx5p33_ASAP7_75t_R g680 ( 
.A(n_631),
.Y(n_680)
);

CKINVDCx20_ASAP7_75t_R g681 ( 
.A(n_569),
.Y(n_681)
);

CKINVDCx5p33_ASAP7_75t_R g682 ( 
.A(n_619),
.Y(n_682)
);

BUFx10_ASAP7_75t_L g683 ( 
.A(n_557),
.Y(n_683)
);

CKINVDCx20_ASAP7_75t_R g684 ( 
.A(n_585),
.Y(n_684)
);

INVx2_ASAP7_75t_L g685 ( 
.A(n_558),
.Y(n_685)
);

CKINVDCx20_ASAP7_75t_R g686 ( 
.A(n_626),
.Y(n_686)
);

INVx1_ASAP7_75t_L g687 ( 
.A(n_529),
.Y(n_687)
);

CKINVDCx5p33_ASAP7_75t_R g688 ( 
.A(n_639),
.Y(n_688)
);

INVxp67_ASAP7_75t_L g689 ( 
.A(n_669),
.Y(n_689)
);

INVxp67_ASAP7_75t_L g690 ( 
.A(n_583),
.Y(n_690)
);

INVx1_ASAP7_75t_L g691 ( 
.A(n_542),
.Y(n_691)
);

BUFx2_ASAP7_75t_L g692 ( 
.A(n_528),
.Y(n_692)
);

CKINVDCx5p33_ASAP7_75t_R g693 ( 
.A(n_666),
.Y(n_693)
);

CKINVDCx20_ASAP7_75t_R g694 ( 
.A(n_652),
.Y(n_694)
);

INVx2_ASAP7_75t_L g695 ( 
.A(n_544),
.Y(n_695)
);

INVx1_ASAP7_75t_L g696 ( 
.A(n_547),
.Y(n_696)
);

NAND2xp33_ASAP7_75t_R g697 ( 
.A(n_541),
.B(n_324),
.Y(n_697)
);

CKINVDCx20_ASAP7_75t_R g698 ( 
.A(n_658),
.Y(n_698)
);

INVx1_ASAP7_75t_L g699 ( 
.A(n_561),
.Y(n_699)
);

INVx1_ASAP7_75t_L g700 ( 
.A(n_562),
.Y(n_700)
);

CKINVDCx5p33_ASAP7_75t_R g701 ( 
.A(n_582),
.Y(n_701)
);

NOR2xp33_ASAP7_75t_R g702 ( 
.A(n_629),
.B(n_432),
.Y(n_702)
);

INVx2_ASAP7_75t_L g703 ( 
.A(n_532),
.Y(n_703)
);

BUFx6f_ASAP7_75t_L g704 ( 
.A(n_530),
.Y(n_704)
);

CKINVDCx5p33_ASAP7_75t_R g705 ( 
.A(n_613),
.Y(n_705)
);

INVx2_ASAP7_75t_L g706 ( 
.A(n_556),
.Y(n_706)
);

INVx2_ASAP7_75t_L g707 ( 
.A(n_530),
.Y(n_707)
);

NAND2xp5_ASAP7_75t_L g708 ( 
.A(n_627),
.B(n_328),
.Y(n_708)
);

BUFx3_ASAP7_75t_L g709 ( 
.A(n_590),
.Y(n_709)
);

CKINVDCx5p33_ASAP7_75t_R g710 ( 
.A(n_595),
.Y(n_710)
);

NAND2xp5_ASAP7_75t_L g711 ( 
.A(n_630),
.B(n_331),
.Y(n_711)
);

CKINVDCx5p33_ASAP7_75t_R g712 ( 
.A(n_596),
.Y(n_712)
);

AND2x2_ASAP7_75t_L g713 ( 
.A(n_586),
.B(n_370),
.Y(n_713)
);

CKINVDCx20_ASAP7_75t_R g714 ( 
.A(n_599),
.Y(n_714)
);

CKINVDCx20_ASAP7_75t_R g715 ( 
.A(n_637),
.Y(n_715)
);

CKINVDCx5p33_ASAP7_75t_R g716 ( 
.A(n_541),
.Y(n_716)
);

CKINVDCx5p33_ASAP7_75t_R g717 ( 
.A(n_550),
.Y(n_717)
);

CKINVDCx5p33_ASAP7_75t_R g718 ( 
.A(n_550),
.Y(n_718)
);

CKINVDCx5p33_ASAP7_75t_R g719 ( 
.A(n_553),
.Y(n_719)
);

INVx1_ASAP7_75t_L g720 ( 
.A(n_646),
.Y(n_720)
);

NOR2xp33_ASAP7_75t_R g721 ( 
.A(n_546),
.B(n_450),
.Y(n_721)
);

NOR2xp67_ASAP7_75t_L g722 ( 
.A(n_623),
.B(n_348),
.Y(n_722)
);

INVx1_ASAP7_75t_L g723 ( 
.A(n_648),
.Y(n_723)
);

CKINVDCx5p33_ASAP7_75t_R g724 ( 
.A(n_545),
.Y(n_724)
);

CKINVDCx5p33_ASAP7_75t_R g725 ( 
.A(n_552),
.Y(n_725)
);

CKINVDCx20_ASAP7_75t_R g726 ( 
.A(n_535),
.Y(n_726)
);

CKINVDCx5p33_ASAP7_75t_R g727 ( 
.A(n_587),
.Y(n_727)
);

CKINVDCx5p33_ASAP7_75t_R g728 ( 
.A(n_608),
.Y(n_728)
);

INVx1_ASAP7_75t_L g729 ( 
.A(n_653),
.Y(n_729)
);

NOR2xp33_ASAP7_75t_R g730 ( 
.A(n_589),
.B(n_464),
.Y(n_730)
);

NOR2xp33_ASAP7_75t_R g731 ( 
.A(n_589),
.B(n_482),
.Y(n_731)
);

CKINVDCx5p33_ASAP7_75t_R g732 ( 
.A(n_618),
.Y(n_732)
);

CKINVDCx5p33_ASAP7_75t_R g733 ( 
.A(n_549),
.Y(n_733)
);

CKINVDCx5p33_ASAP7_75t_R g734 ( 
.A(n_590),
.Y(n_734)
);

INVx1_ASAP7_75t_L g735 ( 
.A(n_655),
.Y(n_735)
);

NAND2xp33_ASAP7_75t_R g736 ( 
.A(n_535),
.B(n_334),
.Y(n_736)
);

BUFx6f_ASAP7_75t_L g737 ( 
.A(n_530),
.Y(n_737)
);

CKINVDCx8_ASAP7_75t_R g738 ( 
.A(n_603),
.Y(n_738)
);

NOR2xp33_ASAP7_75t_R g739 ( 
.A(n_589),
.B(n_512),
.Y(n_739)
);

CKINVDCx5p33_ASAP7_75t_R g740 ( 
.A(n_584),
.Y(n_740)
);

CKINVDCx5p33_ASAP7_75t_R g741 ( 
.A(n_584),
.Y(n_741)
);

INVx1_ASAP7_75t_L g742 ( 
.A(n_656),
.Y(n_742)
);

INVx2_ASAP7_75t_L g743 ( 
.A(n_534),
.Y(n_743)
);

CKINVDCx5p33_ASAP7_75t_R g744 ( 
.A(n_617),
.Y(n_744)
);

CKINVDCx20_ASAP7_75t_R g745 ( 
.A(n_617),
.Y(n_745)
);

BUFx6f_ASAP7_75t_L g746 ( 
.A(n_534),
.Y(n_746)
);

CKINVDCx20_ASAP7_75t_R g747 ( 
.A(n_540),
.Y(n_747)
);

NAND2xp33_ASAP7_75t_R g748 ( 
.A(n_603),
.B(n_638),
.Y(n_748)
);

CKINVDCx20_ASAP7_75t_R g749 ( 
.A(n_625),
.Y(n_749)
);

CKINVDCx5p33_ASAP7_75t_R g750 ( 
.A(n_623),
.Y(n_750)
);

INVx1_ASAP7_75t_L g751 ( 
.A(n_661),
.Y(n_751)
);

INVx2_ASAP7_75t_SL g752 ( 
.A(n_571),
.Y(n_752)
);

BUFx6f_ASAP7_75t_L g753 ( 
.A(n_534),
.Y(n_753)
);

CKINVDCx5p33_ASAP7_75t_R g754 ( 
.A(n_623),
.Y(n_754)
);

CKINVDCx5p33_ASAP7_75t_R g755 ( 
.A(n_634),
.Y(n_755)
);

INVx2_ASAP7_75t_L g756 ( 
.A(n_536),
.Y(n_756)
);

CKINVDCx20_ASAP7_75t_R g757 ( 
.A(n_616),
.Y(n_757)
);

BUFx6f_ASAP7_75t_L g758 ( 
.A(n_536),
.Y(n_758)
);

BUFx3_ASAP7_75t_L g759 ( 
.A(n_591),
.Y(n_759)
);

CKINVDCx5p33_ASAP7_75t_R g760 ( 
.A(n_634),
.Y(n_760)
);

CKINVDCx5p33_ASAP7_75t_R g761 ( 
.A(n_634),
.Y(n_761)
);

CKINVDCx5p33_ASAP7_75t_R g762 ( 
.A(n_643),
.Y(n_762)
);

NOR2xp33_ASAP7_75t_R g763 ( 
.A(n_643),
.B(n_336),
.Y(n_763)
);

CKINVDCx5p33_ASAP7_75t_R g764 ( 
.A(n_643),
.Y(n_764)
);

AOI21x1_ASAP7_75t_L g765 ( 
.A1(n_649),
.A2(n_671),
.B(n_579),
.Y(n_765)
);

CKINVDCx5p33_ASAP7_75t_R g766 ( 
.A(n_591),
.Y(n_766)
);

HB1xp67_ASAP7_75t_L g767 ( 
.A(n_572),
.Y(n_767)
);

NAND2xp5_ASAP7_75t_SL g768 ( 
.A(n_733),
.B(n_675),
.Y(n_768)
);

NAND2xp5_ASAP7_75t_L g769 ( 
.A(n_765),
.B(n_578),
.Y(n_769)
);

HB1xp67_ASAP7_75t_L g770 ( 
.A(n_722),
.Y(n_770)
);

AND2x2_ASAP7_75t_L g771 ( 
.A(n_689),
.B(n_667),
.Y(n_771)
);

HB1xp67_ASAP7_75t_L g772 ( 
.A(n_689),
.Y(n_772)
);

NOR2xp67_ASAP7_75t_L g773 ( 
.A(n_679),
.B(n_548),
.Y(n_773)
);

NOR2xp33_ASAP7_75t_L g774 ( 
.A(n_690),
.B(n_638),
.Y(n_774)
);

INVx8_ASAP7_75t_L g775 ( 
.A(n_684),
.Y(n_775)
);

NOR2xp33_ASAP7_75t_L g776 ( 
.A(n_738),
.B(n_642),
.Y(n_776)
);

AND2x2_ASAP7_75t_L g777 ( 
.A(n_672),
.B(n_670),
.Y(n_777)
);

NOR2xp33_ASAP7_75t_L g778 ( 
.A(n_679),
.B(n_642),
.Y(n_778)
);

INVxp67_ASAP7_75t_L g779 ( 
.A(n_736),
.Y(n_779)
);

INVx2_ASAP7_75t_L g780 ( 
.A(n_707),
.Y(n_780)
);

CKINVDCx5p33_ASAP7_75t_R g781 ( 
.A(n_682),
.Y(n_781)
);

INVx2_ASAP7_75t_L g782 ( 
.A(n_743),
.Y(n_782)
);

NOR3xp33_ASAP7_75t_L g783 ( 
.A(n_716),
.B(n_636),
.C(n_527),
.Y(n_783)
);

INVx2_ASAP7_75t_L g784 ( 
.A(n_756),
.Y(n_784)
);

INVx1_ASAP7_75t_L g785 ( 
.A(n_767),
.Y(n_785)
);

NAND2xp5_ASAP7_75t_L g786 ( 
.A(n_678),
.B(n_588),
.Y(n_786)
);

INVx2_ASAP7_75t_L g787 ( 
.A(n_704),
.Y(n_787)
);

NAND2xp5_ASAP7_75t_L g788 ( 
.A(n_685),
.B(n_602),
.Y(n_788)
);

INVx1_ASAP7_75t_L g789 ( 
.A(n_673),
.Y(n_789)
);

NAND2xp5_ASAP7_75t_L g790 ( 
.A(n_766),
.B(n_644),
.Y(n_790)
);

NAND2xp5_ASAP7_75t_L g791 ( 
.A(n_687),
.B(n_604),
.Y(n_791)
);

NAND2xp5_ASAP7_75t_L g792 ( 
.A(n_708),
.B(n_644),
.Y(n_792)
);

NOR2xp33_ASAP7_75t_L g793 ( 
.A(n_708),
.B(n_563),
.Y(n_793)
);

BUFx6f_ASAP7_75t_L g794 ( 
.A(n_704),
.Y(n_794)
);

NOR2xp33_ASAP7_75t_L g795 ( 
.A(n_711),
.B(n_563),
.Y(n_795)
);

INVx2_ASAP7_75t_L g796 ( 
.A(n_704),
.Y(n_796)
);

NAND2xp5_ASAP7_75t_L g797 ( 
.A(n_711),
.B(n_644),
.Y(n_797)
);

INVx2_ASAP7_75t_L g798 ( 
.A(n_737),
.Y(n_798)
);

NAND2xp5_ASAP7_75t_L g799 ( 
.A(n_691),
.B(n_611),
.Y(n_799)
);

AND2x2_ASAP7_75t_L g800 ( 
.A(n_713),
.B(n_609),
.Y(n_800)
);

NAND2xp5_ASAP7_75t_L g801 ( 
.A(n_696),
.B(n_663),
.Y(n_801)
);

BUFx5_ASAP7_75t_L g802 ( 
.A(n_699),
.Y(n_802)
);

INVxp67_ASAP7_75t_L g803 ( 
.A(n_697),
.Y(n_803)
);

OAI22xp33_ASAP7_75t_L g804 ( 
.A1(n_748),
.A2(n_615),
.B1(n_645),
.B2(n_668),
.Y(n_804)
);

NOR3xp33_ASAP7_75t_L g805 ( 
.A(n_717),
.B(n_719),
.C(n_718),
.Y(n_805)
);

BUFx6f_ASAP7_75t_L g806 ( 
.A(n_737),
.Y(n_806)
);

AND2x2_ASAP7_75t_L g807 ( 
.A(n_692),
.B(n_734),
.Y(n_807)
);

INVx3_ASAP7_75t_L g808 ( 
.A(n_737),
.Y(n_808)
);

INVx2_ASAP7_75t_L g809 ( 
.A(n_746),
.Y(n_809)
);

INVx2_ASAP7_75t_L g810 ( 
.A(n_746),
.Y(n_810)
);

NAND3xp33_ASAP7_75t_L g811 ( 
.A(n_700),
.B(n_640),
.C(n_633),
.Y(n_811)
);

INVx2_ASAP7_75t_L g812 ( 
.A(n_746),
.Y(n_812)
);

INVx2_ASAP7_75t_L g813 ( 
.A(n_753),
.Y(n_813)
);

INVx2_ASAP7_75t_L g814 ( 
.A(n_753),
.Y(n_814)
);

NAND2xp5_ASAP7_75t_SL g815 ( 
.A(n_702),
.B(n_574),
.Y(n_815)
);

INVx1_ASAP7_75t_L g816 ( 
.A(n_673),
.Y(n_816)
);

NAND2xp5_ASAP7_75t_L g817 ( 
.A(n_759),
.B(n_654),
.Y(n_817)
);

NOR3xp33_ASAP7_75t_L g818 ( 
.A(n_752),
.B(n_436),
.C(n_348),
.Y(n_818)
);

INVx2_ASAP7_75t_SL g819 ( 
.A(n_732),
.Y(n_819)
);

NAND2xp33_ASAP7_75t_L g820 ( 
.A(n_730),
.B(n_606),
.Y(n_820)
);

NOR3xp33_ASAP7_75t_L g821 ( 
.A(n_720),
.B(n_651),
.C(n_650),
.Y(n_821)
);

NAND2xp5_ASAP7_75t_L g822 ( 
.A(n_695),
.B(n_593),
.Y(n_822)
);

NOR2xp67_ASAP7_75t_L g823 ( 
.A(n_750),
.B(n_548),
.Y(n_823)
);

NOR2xp67_ASAP7_75t_L g824 ( 
.A(n_754),
.B(n_548),
.Y(n_824)
);

BUFx6f_ASAP7_75t_L g825 ( 
.A(n_753),
.Y(n_825)
);

INVx2_ASAP7_75t_L g826 ( 
.A(n_758),
.Y(n_826)
);

AND2x2_ASAP7_75t_L g827 ( 
.A(n_755),
.B(n_657),
.Y(n_827)
);

NAND2xp5_ASAP7_75t_L g828 ( 
.A(n_723),
.B(n_593),
.Y(n_828)
);

AND2x2_ASAP7_75t_L g829 ( 
.A(n_760),
.B(n_662),
.Y(n_829)
);

INVx1_ASAP7_75t_L g830 ( 
.A(n_703),
.Y(n_830)
);

INVx2_ASAP7_75t_L g831 ( 
.A(n_758),
.Y(n_831)
);

INVx2_ASAP7_75t_SL g832 ( 
.A(n_724),
.Y(n_832)
);

BUFx3_ASAP7_75t_L g833 ( 
.A(n_676),
.Y(n_833)
);

NOR2xp67_ASAP7_75t_L g834 ( 
.A(n_761),
.B(n_564),
.Y(n_834)
);

NAND2xp5_ASAP7_75t_L g835 ( 
.A(n_758),
.B(n_654),
.Y(n_835)
);

NAND2xp33_ASAP7_75t_L g836 ( 
.A(n_731),
.B(n_606),
.Y(n_836)
);

INVxp67_ASAP7_75t_SL g837 ( 
.A(n_709),
.Y(n_837)
);

AOI22xp5_ASAP7_75t_L g838 ( 
.A1(n_757),
.A2(n_749),
.B1(n_747),
.B2(n_686),
.Y(n_838)
);

AO221x1_ASAP7_75t_L g839 ( 
.A1(n_729),
.A2(n_435),
.B1(n_442),
.B2(n_439),
.C(n_434),
.Y(n_839)
);

NOR2xp33_ASAP7_75t_L g840 ( 
.A(n_725),
.B(n_727),
.Y(n_840)
);

NAND2xp5_ASAP7_75t_L g841 ( 
.A(n_735),
.B(n_654),
.Y(n_841)
);

NOR2xp33_ASAP7_75t_L g842 ( 
.A(n_728),
.B(n_581),
.Y(n_842)
);

AND2x2_ASAP7_75t_SL g843 ( 
.A(n_721),
.B(n_581),
.Y(n_843)
);

NAND2xp5_ASAP7_75t_L g844 ( 
.A(n_742),
.B(n_564),
.Y(n_844)
);

INVx1_ASAP7_75t_L g845 ( 
.A(n_706),
.Y(n_845)
);

NOR2xp67_ASAP7_75t_SL g846 ( 
.A(n_762),
.B(n_564),
.Y(n_846)
);

NAND3xp33_ASAP7_75t_L g847 ( 
.A(n_751),
.B(n_664),
.C(n_671),
.Y(n_847)
);

NAND2xp5_ASAP7_75t_L g848 ( 
.A(n_764),
.B(n_593),
.Y(n_848)
);

NAND2xp5_ASAP7_75t_L g849 ( 
.A(n_739),
.B(n_601),
.Y(n_849)
);

INVx3_ASAP7_75t_L g850 ( 
.A(n_683),
.Y(n_850)
);

AND2x2_ASAP7_75t_L g851 ( 
.A(n_763),
.B(n_614),
.Y(n_851)
);

INVx2_ASAP7_75t_L g852 ( 
.A(n_694),
.Y(n_852)
);

NOR2xp33_ASAP7_75t_L g853 ( 
.A(n_698),
.B(n_660),
.Y(n_853)
);

NAND2xp5_ASAP7_75t_SL g854 ( 
.A(n_740),
.B(n_337),
.Y(n_854)
);

AND2x2_ASAP7_75t_L g855 ( 
.A(n_688),
.B(n_622),
.Y(n_855)
);

AND2x2_ASAP7_75t_SL g856 ( 
.A(n_843),
.B(n_568),
.Y(n_856)
);

NOR2xp33_ASAP7_75t_R g857 ( 
.A(n_781),
.B(n_674),
.Y(n_857)
);

CKINVDCx5p33_ASAP7_75t_R g858 ( 
.A(n_840),
.Y(n_858)
);

NAND2xp5_ASAP7_75t_SL g859 ( 
.A(n_803),
.B(n_693),
.Y(n_859)
);

NAND2xp5_ASAP7_75t_L g860 ( 
.A(n_793),
.B(n_795),
.Y(n_860)
);

BUFx3_ASAP7_75t_L g861 ( 
.A(n_833),
.Y(n_861)
);

INVx1_ASAP7_75t_L g862 ( 
.A(n_822),
.Y(n_862)
);

OR2x6_ASAP7_75t_L g863 ( 
.A(n_775),
.B(n_580),
.Y(n_863)
);

OR2x6_ASAP7_75t_L g864 ( 
.A(n_775),
.B(n_592),
.Y(n_864)
);

INVx1_ASAP7_75t_L g865 ( 
.A(n_786),
.Y(n_865)
);

NOR2xp33_ASAP7_75t_L g866 ( 
.A(n_779),
.B(n_714),
.Y(n_866)
);

NAND2xp5_ASAP7_75t_L g867 ( 
.A(n_778),
.B(n_777),
.Y(n_867)
);

BUFx3_ASAP7_75t_L g868 ( 
.A(n_775),
.Y(n_868)
);

BUFx3_ASAP7_75t_L g869 ( 
.A(n_852),
.Y(n_869)
);

INVx2_ASAP7_75t_L g870 ( 
.A(n_780),
.Y(n_870)
);

INVx1_ASAP7_75t_L g871 ( 
.A(n_822),
.Y(n_871)
);

INVxp67_ASAP7_75t_L g872 ( 
.A(n_800),
.Y(n_872)
);

OR2x6_ASAP7_75t_L g873 ( 
.A(n_850),
.B(n_594),
.Y(n_873)
);

BUFx2_ASAP7_75t_L g874 ( 
.A(n_772),
.Y(n_874)
);

NAND2xp5_ASAP7_75t_SL g875 ( 
.A(n_776),
.B(n_683),
.Y(n_875)
);

AOI22x1_ASAP7_75t_L g876 ( 
.A1(n_771),
.A2(n_451),
.B1(n_453),
.B2(n_444),
.Y(n_876)
);

INVx1_ASAP7_75t_L g877 ( 
.A(n_828),
.Y(n_877)
);

INVx2_ASAP7_75t_SL g878 ( 
.A(n_827),
.Y(n_878)
);

NOR2x2_ASAP7_75t_L g879 ( 
.A(n_804),
.B(n_526),
.Y(n_879)
);

INVx1_ASAP7_75t_L g880 ( 
.A(n_828),
.Y(n_880)
);

INVx1_ASAP7_75t_L g881 ( 
.A(n_789),
.Y(n_881)
);

NOR3xp33_ASAP7_75t_L g882 ( 
.A(n_768),
.B(n_805),
.C(n_783),
.Y(n_882)
);

INVx1_ASAP7_75t_L g883 ( 
.A(n_786),
.Y(n_883)
);

AND2x2_ASAP7_75t_L g884 ( 
.A(n_853),
.B(n_807),
.Y(n_884)
);

CKINVDCx5p33_ASAP7_75t_R g885 ( 
.A(n_850),
.Y(n_885)
);

BUFx2_ASAP7_75t_L g886 ( 
.A(n_838),
.Y(n_886)
);

BUFx3_ASAP7_75t_L g887 ( 
.A(n_785),
.Y(n_887)
);

NAND3xp33_ASAP7_75t_SL g888 ( 
.A(n_818),
.B(n_726),
.C(n_715),
.Y(n_888)
);

INVx2_ASAP7_75t_SL g889 ( 
.A(n_829),
.Y(n_889)
);

AOI22xp5_ASAP7_75t_L g890 ( 
.A1(n_774),
.A2(n_345),
.B1(n_347),
.B2(n_343),
.Y(n_890)
);

BUFx4f_ASAP7_75t_L g891 ( 
.A(n_819),
.Y(n_891)
);

NAND2xp5_ASAP7_75t_L g892 ( 
.A(n_802),
.B(n_601),
.Y(n_892)
);

INVx1_ASAP7_75t_L g893 ( 
.A(n_816),
.Y(n_893)
);

CKINVDCx5p33_ASAP7_75t_R g894 ( 
.A(n_832),
.Y(n_894)
);

BUFx6f_ASAP7_75t_L g895 ( 
.A(n_794),
.Y(n_895)
);

INVx2_ASAP7_75t_SL g896 ( 
.A(n_855),
.Y(n_896)
);

INVx4_ASAP7_75t_L g897 ( 
.A(n_794),
.Y(n_897)
);

NAND2xp5_ASAP7_75t_L g898 ( 
.A(n_802),
.B(n_605),
.Y(n_898)
);

INVx2_ASAP7_75t_SL g899 ( 
.A(n_848),
.Y(n_899)
);

CKINVDCx6p67_ASAP7_75t_R g900 ( 
.A(n_854),
.Y(n_900)
);

NAND2xp5_ASAP7_75t_L g901 ( 
.A(n_802),
.B(n_605),
.Y(n_901)
);

INVx2_ASAP7_75t_L g902 ( 
.A(n_782),
.Y(n_902)
);

INVx2_ASAP7_75t_L g903 ( 
.A(n_784),
.Y(n_903)
);

NAND2xp5_ASAP7_75t_SL g904 ( 
.A(n_849),
.B(n_705),
.Y(n_904)
);

CKINVDCx20_ASAP7_75t_R g905 ( 
.A(n_849),
.Y(n_905)
);

AOI22xp5_ASAP7_75t_L g906 ( 
.A1(n_820),
.A2(n_350),
.B1(n_352),
.B2(n_349),
.Y(n_906)
);

INVx2_ASAP7_75t_SL g907 ( 
.A(n_848),
.Y(n_907)
);

NOR2xp33_ASAP7_75t_L g908 ( 
.A(n_815),
.B(n_741),
.Y(n_908)
);

A2O1A1Ixp33_ASAP7_75t_L g909 ( 
.A1(n_769),
.A2(n_576),
.B(n_632),
.C(n_628),
.Y(n_909)
);

NOR2x2_ASAP7_75t_L g910 ( 
.A(n_787),
.B(n_555),
.Y(n_910)
);

INVx2_ASAP7_75t_SL g911 ( 
.A(n_851),
.Y(n_911)
);

NAND2xp5_ASAP7_75t_SL g912 ( 
.A(n_842),
.B(n_356),
.Y(n_912)
);

AOI22xp5_ASAP7_75t_L g913 ( 
.A1(n_836),
.A2(n_360),
.B1(n_361),
.B2(n_359),
.Y(n_913)
);

NAND2xp5_ASAP7_75t_SL g914 ( 
.A(n_773),
.B(n_365),
.Y(n_914)
);

NAND2xp5_ASAP7_75t_L g915 ( 
.A(n_792),
.B(n_607),
.Y(n_915)
);

OR2x2_ASAP7_75t_L g916 ( 
.A(n_837),
.B(n_677),
.Y(n_916)
);

AND2x2_ASAP7_75t_L g917 ( 
.A(n_770),
.B(n_701),
.Y(n_917)
);

NAND2xp5_ASAP7_75t_L g918 ( 
.A(n_797),
.B(n_607),
.Y(n_918)
);

INVx2_ASAP7_75t_L g919 ( 
.A(n_830),
.Y(n_919)
);

BUFx2_ASAP7_75t_L g920 ( 
.A(n_796),
.Y(n_920)
);

AOI21xp5_ASAP7_75t_L g921 ( 
.A1(n_769),
.A2(n_577),
.B(n_573),
.Y(n_921)
);

BUFx2_ASAP7_75t_L g922 ( 
.A(n_798),
.Y(n_922)
);

INVxp67_ASAP7_75t_L g923 ( 
.A(n_845),
.Y(n_923)
);

NAND2xp5_ASAP7_75t_L g924 ( 
.A(n_801),
.B(n_621),
.Y(n_924)
);

BUFx12f_ASAP7_75t_L g925 ( 
.A(n_794),
.Y(n_925)
);

INVx5_ASAP7_75t_L g926 ( 
.A(n_806),
.Y(n_926)
);

NAND2xp5_ASAP7_75t_L g927 ( 
.A(n_801),
.B(n_621),
.Y(n_927)
);

BUFx2_ASAP7_75t_L g928 ( 
.A(n_809),
.Y(n_928)
);

INVx1_ASAP7_75t_L g929 ( 
.A(n_788),
.Y(n_929)
);

INVx1_ASAP7_75t_L g930 ( 
.A(n_788),
.Y(n_930)
);

AOI22xp5_ASAP7_75t_L g931 ( 
.A1(n_839),
.A2(n_367),
.B1(n_373),
.B2(n_368),
.Y(n_931)
);

INVx1_ASAP7_75t_L g932 ( 
.A(n_791),
.Y(n_932)
);

OAI21xp33_ASAP7_75t_L g933 ( 
.A1(n_821),
.A2(n_600),
.B(n_597),
.Y(n_933)
);

NOR2xp33_ASAP7_75t_R g934 ( 
.A(n_808),
.B(n_680),
.Y(n_934)
);

AOI22xp5_ASAP7_75t_SL g935 ( 
.A1(n_790),
.A2(n_681),
.B1(n_745),
.B2(n_565),
.Y(n_935)
);

BUFx4f_ASAP7_75t_L g936 ( 
.A(n_806),
.Y(n_936)
);

AND2x4_ASAP7_75t_L g937 ( 
.A(n_810),
.B(n_620),
.Y(n_937)
);

INVx2_ASAP7_75t_L g938 ( 
.A(n_808),
.Y(n_938)
);

NAND2xp5_ASAP7_75t_L g939 ( 
.A(n_799),
.B(n_624),
.Y(n_939)
);

INVx1_ASAP7_75t_L g940 ( 
.A(n_812),
.Y(n_940)
);

INVx3_ASAP7_75t_L g941 ( 
.A(n_813),
.Y(n_941)
);

NAND2xp5_ASAP7_75t_L g942 ( 
.A(n_814),
.B(n_624),
.Y(n_942)
);

INVx2_ASAP7_75t_L g943 ( 
.A(n_826),
.Y(n_943)
);

AND2x4_ASAP7_75t_L g944 ( 
.A(n_831),
.B(n_454),
.Y(n_944)
);

NAND2xp5_ASAP7_75t_L g945 ( 
.A(n_806),
.B(n_624),
.Y(n_945)
);

AOI21x1_ASAP7_75t_L g946 ( 
.A1(n_921),
.A2(n_844),
.B(n_835),
.Y(n_946)
);

NAND2xp5_ASAP7_75t_L g947 ( 
.A(n_860),
.B(n_825),
.Y(n_947)
);

NAND2xp5_ASAP7_75t_L g948 ( 
.A(n_932),
.B(n_825),
.Y(n_948)
);

NOR2xp33_ASAP7_75t_L g949 ( 
.A(n_858),
.B(n_744),
.Y(n_949)
);

AOI21xp5_ASAP7_75t_L g950 ( 
.A1(n_924),
.A2(n_817),
.B(n_841),
.Y(n_950)
);

BUFx6f_ASAP7_75t_L g951 ( 
.A(n_895),
.Y(n_951)
);

AOI21xp5_ASAP7_75t_L g952 ( 
.A1(n_927),
.A2(n_577),
.B(n_573),
.Y(n_952)
);

NAND2xp5_ASAP7_75t_L g953 ( 
.A(n_929),
.B(n_825),
.Y(n_953)
);

NAND2xp5_ASAP7_75t_SL g954 ( 
.A(n_867),
.B(n_823),
.Y(n_954)
);

AOI221xp5_ASAP7_75t_L g955 ( 
.A1(n_908),
.A2(n_811),
.B1(n_847),
.B2(n_462),
.C(n_473),
.Y(n_955)
);

INVx3_ASAP7_75t_L g956 ( 
.A(n_941),
.Y(n_956)
);

NAND3xp33_ASAP7_75t_L g957 ( 
.A(n_866),
.B(n_811),
.C(n_847),
.Y(n_957)
);

A2O1A1Ixp33_ASAP7_75t_L g958 ( 
.A1(n_930),
.A2(n_659),
.B(n_501),
.C(n_366),
.Y(n_958)
);

BUFx2_ASAP7_75t_L g959 ( 
.A(n_874),
.Y(n_959)
);

NAND2xp5_ASAP7_75t_L g960 ( 
.A(n_865),
.B(n_493),
.Y(n_960)
);

BUFx6f_ASAP7_75t_L g961 ( 
.A(n_895),
.Y(n_961)
);

NAND2xp5_ASAP7_75t_L g962 ( 
.A(n_883),
.B(n_496),
.Y(n_962)
);

AOI22xp33_ASAP7_75t_L g963 ( 
.A1(n_856),
.A2(n_612),
.B1(n_606),
.B2(n_505),
.Y(n_963)
);

AOI21xp5_ASAP7_75t_L g964 ( 
.A1(n_883),
.A2(n_537),
.B(n_536),
.Y(n_964)
);

BUFx12f_ASAP7_75t_L g965 ( 
.A(n_885),
.Y(n_965)
);

NAND2xp5_ASAP7_75t_L g966 ( 
.A(n_877),
.B(n_504),
.Y(n_966)
);

AND2x4_ASAP7_75t_L g967 ( 
.A(n_861),
.B(n_508),
.Y(n_967)
);

OAI22xp5_ASAP7_75t_L g968 ( 
.A1(n_872),
.A2(n_518),
.B1(n_519),
.B2(n_513),
.Y(n_968)
);

NOR2xp33_ASAP7_75t_L g969 ( 
.A(n_884),
.B(n_539),
.Y(n_969)
);

AOI22xp33_ASAP7_75t_L g970 ( 
.A1(n_862),
.A2(n_612),
.B1(n_524),
.B2(n_523),
.Y(n_970)
);

NAND2xp5_ASAP7_75t_L g971 ( 
.A(n_880),
.B(n_824),
.Y(n_971)
);

NAND2xp5_ASAP7_75t_L g972 ( 
.A(n_871),
.B(n_834),
.Y(n_972)
);

INVx2_ASAP7_75t_L g973 ( 
.A(n_937),
.Y(n_973)
);

AOI21xp5_ASAP7_75t_L g974 ( 
.A1(n_892),
.A2(n_543),
.B(n_537),
.Y(n_974)
);

NAND2xp5_ASAP7_75t_SL g975 ( 
.A(n_911),
.B(n_375),
.Y(n_975)
);

NOR2x1_ASAP7_75t_L g976 ( 
.A(n_875),
.B(n_533),
.Y(n_976)
);

AOI21xp5_ASAP7_75t_L g977 ( 
.A1(n_898),
.A2(n_543),
.B(n_537),
.Y(n_977)
);

NAND2xp5_ASAP7_75t_SL g978 ( 
.A(n_899),
.B(n_376),
.Y(n_978)
);

AOI21xp5_ASAP7_75t_L g979 ( 
.A1(n_901),
.A2(n_551),
.B(n_543),
.Y(n_979)
);

NOR2xp33_ASAP7_75t_L g980 ( 
.A(n_907),
.B(n_710),
.Y(n_980)
);

A2O1A1Ixp33_ASAP7_75t_L g981 ( 
.A1(n_882),
.A2(n_471),
.B(n_380),
.C(n_382),
.Y(n_981)
);

OAI21xp33_ASAP7_75t_L g982 ( 
.A1(n_896),
.A2(n_712),
.B(n_385),
.Y(n_982)
);

INVx2_ASAP7_75t_L g983 ( 
.A(n_870),
.Y(n_983)
);

INVx1_ASAP7_75t_SL g984 ( 
.A(n_905),
.Y(n_984)
);

INVx1_ASAP7_75t_L g985 ( 
.A(n_881),
.Y(n_985)
);

AOI21xp5_ASAP7_75t_L g986 ( 
.A1(n_936),
.A2(n_559),
.B(n_554),
.Y(n_986)
);

NOR3xp33_ASAP7_75t_SL g987 ( 
.A(n_888),
.B(n_388),
.C(n_377),
.Y(n_987)
);

INVx2_ASAP7_75t_L g988 ( 
.A(n_902),
.Y(n_988)
);

AND2x2_ASAP7_75t_L g989 ( 
.A(n_878),
.B(n_660),
.Y(n_989)
);

O2A1O1Ixp33_ASAP7_75t_L g990 ( 
.A1(n_939),
.A2(n_635),
.B(n_641),
.C(n_389),
.Y(n_990)
);

AO22x1_ASAP7_75t_L g991 ( 
.A1(n_886),
.A2(n_481),
.B1(n_393),
.B2(n_396),
.Y(n_991)
);

NAND2x1p5_ASAP7_75t_L g992 ( 
.A(n_891),
.B(n_846),
.Y(n_992)
);

AO32x1_ASAP7_75t_L g993 ( 
.A1(n_940),
.A2(n_533),
.A3(n_41),
.B1(n_42),
.B2(n_43),
.Y(n_993)
);

OAI22xp5_ASAP7_75t_L g994 ( 
.A1(n_889),
.A2(n_474),
.B1(n_398),
.B2(n_404),
.Y(n_994)
);

INVx3_ASAP7_75t_SL g995 ( 
.A(n_894),
.Y(n_995)
);

AOI21xp5_ASAP7_75t_L g996 ( 
.A1(n_936),
.A2(n_909),
.B(n_915),
.Y(n_996)
);

AOI21xp5_ASAP7_75t_L g997 ( 
.A1(n_918),
.A2(n_560),
.B(n_559),
.Y(n_997)
);

AOI21xp5_ASAP7_75t_L g998 ( 
.A1(n_926),
.A2(n_897),
.B(n_893),
.Y(n_998)
);

NAND2xp5_ASAP7_75t_L g999 ( 
.A(n_903),
.B(n_635),
.Y(n_999)
);

NAND2xp5_ASAP7_75t_L g1000 ( 
.A(n_919),
.B(n_635),
.Y(n_1000)
);

INVx5_ASAP7_75t_L g1001 ( 
.A(n_925),
.Y(n_1001)
);

INVx6_ASAP7_75t_L g1002 ( 
.A(n_868),
.Y(n_1002)
);

NAND2xp5_ASAP7_75t_SL g1003 ( 
.A(n_891),
.B(n_390),
.Y(n_1003)
);

INVx3_ASAP7_75t_L g1004 ( 
.A(n_941),
.Y(n_1004)
);

NAND2xp5_ASAP7_75t_L g1005 ( 
.A(n_923),
.B(n_641),
.Y(n_1005)
);

INVx5_ASAP7_75t_L g1006 ( 
.A(n_873),
.Y(n_1006)
);

HB1xp67_ASAP7_75t_L g1007 ( 
.A(n_887),
.Y(n_1007)
);

INVx1_ASAP7_75t_L g1008 ( 
.A(n_945),
.Y(n_1008)
);

NAND2xp5_ASAP7_75t_L g1009 ( 
.A(n_920),
.B(n_641),
.Y(n_1009)
);

NAND2xp5_ASAP7_75t_L g1010 ( 
.A(n_922),
.B(n_412),
.Y(n_1010)
);

A2O1A1Ixp33_ASAP7_75t_L g1011 ( 
.A1(n_906),
.A2(n_475),
.B(n_417),
.C(n_418),
.Y(n_1011)
);

INVx1_ASAP7_75t_L g1012 ( 
.A(n_928),
.Y(n_1012)
);

NAND2xp5_ASAP7_75t_L g1013 ( 
.A(n_890),
.B(n_415),
.Y(n_1013)
);

INVx3_ASAP7_75t_L g1014 ( 
.A(n_895),
.Y(n_1014)
);

NAND2xp5_ASAP7_75t_L g1015 ( 
.A(n_938),
.B(n_420),
.Y(n_1015)
);

INVx2_ASAP7_75t_L g1016 ( 
.A(n_943),
.Y(n_1016)
);

INVx2_ASAP7_75t_L g1017 ( 
.A(n_944),
.Y(n_1017)
);

OAI221xp5_ASAP7_75t_L g1018 ( 
.A1(n_933),
.A2(n_876),
.B1(n_931),
.B2(n_873),
.C(n_913),
.Y(n_1018)
);

INVxp67_ASAP7_75t_L g1019 ( 
.A(n_869),
.Y(n_1019)
);

OAI22xp5_ASAP7_75t_SL g1020 ( 
.A1(n_879),
.A2(n_477),
.B1(n_522),
.B2(n_517),
.Y(n_1020)
);

CKINVDCx16_ASAP7_75t_R g1021 ( 
.A(n_965),
.Y(n_1021)
);

NOR2xp33_ASAP7_75t_L g1022 ( 
.A(n_969),
.B(n_859),
.Y(n_1022)
);

AO21x1_ASAP7_75t_L g1023 ( 
.A1(n_996),
.A2(n_944),
.B(n_942),
.Y(n_1023)
);

BUFx3_ASAP7_75t_L g1024 ( 
.A(n_1002),
.Y(n_1024)
);

INVx1_ASAP7_75t_SL g1025 ( 
.A(n_959),
.Y(n_1025)
);

OAI21x1_ASAP7_75t_L g1026 ( 
.A1(n_946),
.A2(n_876),
.B(n_912),
.Y(n_1026)
);

BUFx4f_ASAP7_75t_SL g1027 ( 
.A(n_995),
.Y(n_1027)
);

INVx2_ASAP7_75t_L g1028 ( 
.A(n_956),
.Y(n_1028)
);

INVx2_ASAP7_75t_L g1029 ( 
.A(n_956),
.Y(n_1029)
);

OAI21xp5_ASAP7_75t_L g1030 ( 
.A1(n_947),
.A2(n_962),
.B(n_960),
.Y(n_1030)
);

BUFx3_ASAP7_75t_L g1031 ( 
.A(n_1002),
.Y(n_1031)
);

INVx1_ASAP7_75t_L g1032 ( 
.A(n_985),
.Y(n_1032)
);

BUFx6f_ASAP7_75t_L g1033 ( 
.A(n_951),
.Y(n_1033)
);

INVx4_ASAP7_75t_L g1034 ( 
.A(n_951),
.Y(n_1034)
);

NAND2x1p5_ASAP7_75t_L g1035 ( 
.A(n_951),
.B(n_897),
.Y(n_1035)
);

INVx2_ASAP7_75t_L g1036 ( 
.A(n_1004),
.Y(n_1036)
);

INVx1_ASAP7_75t_L g1037 ( 
.A(n_983),
.Y(n_1037)
);

OAI21x1_ASAP7_75t_L g1038 ( 
.A1(n_950),
.A2(n_914),
.B(n_904),
.Y(n_1038)
);

BUFx3_ASAP7_75t_L g1039 ( 
.A(n_1001),
.Y(n_1039)
);

AOI22x1_ASAP7_75t_L g1040 ( 
.A1(n_1008),
.A2(n_1016),
.B1(n_988),
.B2(n_998),
.Y(n_1040)
);

INVx3_ASAP7_75t_L g1041 ( 
.A(n_961),
.Y(n_1041)
);

INVx3_ASAP7_75t_L g1042 ( 
.A(n_961),
.Y(n_1042)
);

INVx1_ASAP7_75t_L g1043 ( 
.A(n_953),
.Y(n_1043)
);

INVx2_ASAP7_75t_SL g1044 ( 
.A(n_961),
.Y(n_1044)
);

INVx1_ASAP7_75t_L g1045 ( 
.A(n_948),
.Y(n_1045)
);

AND2x4_ASAP7_75t_L g1046 ( 
.A(n_1017),
.B(n_916),
.Y(n_1046)
);

INVx2_ASAP7_75t_L g1047 ( 
.A(n_1004),
.Y(n_1047)
);

OAI21x1_ASAP7_75t_L g1048 ( 
.A1(n_974),
.A2(n_917),
.B(n_926),
.Y(n_1048)
);

OAI21x1_ASAP7_75t_L g1049 ( 
.A1(n_977),
.A2(n_926),
.B(n_900),
.Y(n_1049)
);

AO21x2_ASAP7_75t_L g1050 ( 
.A1(n_958),
.A2(n_934),
.B(n_857),
.Y(n_1050)
);

INVx2_ASAP7_75t_L g1051 ( 
.A(n_999),
.Y(n_1051)
);

INVx2_ASAP7_75t_SL g1052 ( 
.A(n_1007),
.Y(n_1052)
);

AOI22x1_ASAP7_75t_L g1053 ( 
.A1(n_964),
.A2(n_935),
.B1(n_485),
.B2(n_484),
.Y(n_1053)
);

INVx3_ASAP7_75t_L g1054 ( 
.A(n_1014),
.Y(n_1054)
);

INVx2_ASAP7_75t_SL g1055 ( 
.A(n_1012),
.Y(n_1055)
);

INVx1_ASAP7_75t_L g1056 ( 
.A(n_973),
.Y(n_1056)
);

INVx2_ASAP7_75t_L g1057 ( 
.A(n_1000),
.Y(n_1057)
);

AND2x4_ASAP7_75t_L g1058 ( 
.A(n_1006),
.B(n_863),
.Y(n_1058)
);

OAI21x1_ASAP7_75t_L g1059 ( 
.A1(n_979),
.A2(n_76),
.B(n_75),
.Y(n_1059)
);

INVx1_ASAP7_75t_L g1060 ( 
.A(n_1009),
.Y(n_1060)
);

OAI21x1_ASAP7_75t_L g1061 ( 
.A1(n_990),
.A2(n_92),
.B(n_87),
.Y(n_1061)
);

INVx2_ASAP7_75t_L g1062 ( 
.A(n_966),
.Y(n_1062)
);

AOI22xp33_ASAP7_75t_L g1063 ( 
.A1(n_1018),
.A2(n_665),
.B1(n_864),
.B2(n_863),
.Y(n_1063)
);

NAND2x1p5_ASAP7_75t_L g1064 ( 
.A(n_1001),
.B(n_559),
.Y(n_1064)
);

AO21x2_ASAP7_75t_L g1065 ( 
.A1(n_981),
.A2(n_665),
.B(n_427),
.Y(n_1065)
);

AO21x2_ASAP7_75t_L g1066 ( 
.A1(n_954),
.A2(n_428),
.B(n_423),
.Y(n_1066)
);

CKINVDCx16_ASAP7_75t_R g1067 ( 
.A(n_984),
.Y(n_1067)
);

INVx2_ASAP7_75t_L g1068 ( 
.A(n_989),
.Y(n_1068)
);

INVx4_ASAP7_75t_L g1069 ( 
.A(n_1001),
.Y(n_1069)
);

BUFx4f_ASAP7_75t_L g1070 ( 
.A(n_992),
.Y(n_1070)
);

INVx1_ASAP7_75t_L g1071 ( 
.A(n_1005),
.Y(n_1071)
);

INVx1_ASAP7_75t_L g1072 ( 
.A(n_1015),
.Y(n_1072)
);

BUFx3_ASAP7_75t_L g1073 ( 
.A(n_1006),
.Y(n_1073)
);

INVx1_ASAP7_75t_L g1074 ( 
.A(n_1019),
.Y(n_1074)
);

AO21x2_ASAP7_75t_L g1075 ( 
.A1(n_1011),
.A2(n_438),
.B(n_431),
.Y(n_1075)
);

AND2x4_ASAP7_75t_L g1076 ( 
.A(n_1006),
.B(n_864),
.Y(n_1076)
);

OAI21x1_ASAP7_75t_L g1077 ( 
.A1(n_997),
.A2(n_95),
.B(n_94),
.Y(n_1077)
);

INVx4_ASAP7_75t_L g1078 ( 
.A(n_967),
.Y(n_1078)
);

AO21x2_ASAP7_75t_L g1079 ( 
.A1(n_957),
.A2(n_1013),
.B(n_972),
.Y(n_1079)
);

AO21x2_ASAP7_75t_L g1080 ( 
.A1(n_971),
.A2(n_448),
.B(n_440),
.Y(n_1080)
);

INVx1_ASAP7_75t_SL g1081 ( 
.A(n_967),
.Y(n_1081)
);

BUFx2_ASAP7_75t_SL g1082 ( 
.A(n_1003),
.Y(n_1082)
);

INVx1_ASAP7_75t_L g1083 ( 
.A(n_968),
.Y(n_1083)
);

INVx2_ASAP7_75t_L g1084 ( 
.A(n_993),
.Y(n_1084)
);

INVx2_ASAP7_75t_L g1085 ( 
.A(n_993),
.Y(n_1085)
);

INVx1_ASAP7_75t_L g1086 ( 
.A(n_1010),
.Y(n_1086)
);

INVx1_ASAP7_75t_L g1087 ( 
.A(n_1032),
.Y(n_1087)
);

OA21x2_ASAP7_75t_L g1088 ( 
.A1(n_1023),
.A2(n_1030),
.B(n_1026),
.Y(n_1088)
);

INVx2_ASAP7_75t_L g1089 ( 
.A(n_1037),
.Y(n_1089)
);

INVx3_ASAP7_75t_L g1090 ( 
.A(n_1034),
.Y(n_1090)
);

AND2x2_ASAP7_75t_L g1091 ( 
.A(n_1022),
.B(n_987),
.Y(n_1091)
);

OAI22xp5_ASAP7_75t_L g1092 ( 
.A1(n_1062),
.A2(n_963),
.B1(n_980),
.B2(n_978),
.Y(n_1092)
);

INVx1_ASAP7_75t_L g1093 ( 
.A(n_1056),
.Y(n_1093)
);

BUFx2_ASAP7_75t_SL g1094 ( 
.A(n_1024),
.Y(n_1094)
);

INVx2_ASAP7_75t_L g1095 ( 
.A(n_1028),
.Y(n_1095)
);

INVx2_ASAP7_75t_L g1096 ( 
.A(n_1028),
.Y(n_1096)
);

INVx1_ASAP7_75t_L g1097 ( 
.A(n_1068),
.Y(n_1097)
);

CKINVDCx6p67_ASAP7_75t_R g1098 ( 
.A(n_1024),
.Y(n_1098)
);

INVx1_ASAP7_75t_SL g1099 ( 
.A(n_1025),
.Y(n_1099)
);

NAND2xp5_ASAP7_75t_L g1100 ( 
.A(n_1086),
.B(n_991),
.Y(n_1100)
);

INVxp67_ASAP7_75t_L g1101 ( 
.A(n_1055),
.Y(n_1101)
);

AOI22xp33_ASAP7_75t_L g1102 ( 
.A1(n_1022),
.A2(n_955),
.B1(n_976),
.B2(n_975),
.Y(n_1102)
);

OAI22xp33_ASAP7_75t_L g1103 ( 
.A1(n_1062),
.A2(n_949),
.B1(n_994),
.B2(n_491),
.Y(n_1103)
);

INVx1_ASAP7_75t_L g1104 ( 
.A(n_1068),
.Y(n_1104)
);

INVx1_ASAP7_75t_L g1105 ( 
.A(n_1043),
.Y(n_1105)
);

BUFx3_ASAP7_75t_L g1106 ( 
.A(n_1031),
.Y(n_1106)
);

OAI22xp5_ASAP7_75t_L g1107 ( 
.A1(n_1045),
.A2(n_970),
.B1(n_982),
.B2(n_1020),
.Y(n_1107)
);

INVx2_ASAP7_75t_L g1108 ( 
.A(n_1029),
.Y(n_1108)
);

AOI22xp33_ASAP7_75t_L g1109 ( 
.A1(n_1083),
.A2(n_489),
.B1(n_456),
.B2(n_457),
.Y(n_1109)
);

AOI22xp33_ASAP7_75t_SL g1110 ( 
.A1(n_1082),
.A2(n_910),
.B1(n_452),
.B2(n_498),
.Y(n_1110)
);

NAND2xp5_ASAP7_75t_L g1111 ( 
.A(n_1060),
.B(n_952),
.Y(n_1111)
);

HB1xp67_ASAP7_75t_L g1112 ( 
.A(n_1055),
.Y(n_1112)
);

AND2x2_ASAP7_75t_L g1113 ( 
.A(n_1046),
.B(n_459),
.Y(n_1113)
);

INVx2_ASAP7_75t_L g1114 ( 
.A(n_1029),
.Y(n_1114)
);

INVx2_ASAP7_75t_L g1115 ( 
.A(n_1036),
.Y(n_1115)
);

BUFx2_ASAP7_75t_R g1116 ( 
.A(n_1039),
.Y(n_1116)
);

CKINVDCx5p33_ASAP7_75t_R g1117 ( 
.A(n_1027),
.Y(n_1117)
);

INVx2_ASAP7_75t_L g1118 ( 
.A(n_1036),
.Y(n_1118)
);

AOI22xp33_ASAP7_75t_L g1119 ( 
.A1(n_1063),
.A2(n_500),
.B1(n_465),
.B2(n_467),
.Y(n_1119)
);

AO21x1_ASAP7_75t_L g1120 ( 
.A1(n_1084),
.A2(n_986),
.B(n_41),
.Y(n_1120)
);

INVx1_ASAP7_75t_L g1121 ( 
.A(n_1047),
.Y(n_1121)
);

BUFx6f_ASAP7_75t_L g1122 ( 
.A(n_1033),
.Y(n_1122)
);

INVx2_ASAP7_75t_L g1123 ( 
.A(n_1047),
.Y(n_1123)
);

OAI22xp5_ASAP7_75t_L g1124 ( 
.A1(n_1072),
.A2(n_1071),
.B1(n_1063),
.B2(n_1046),
.Y(n_1124)
);

HB1xp67_ASAP7_75t_L g1125 ( 
.A(n_1052),
.Y(n_1125)
);

BUFx8_ASAP7_75t_L g1126 ( 
.A(n_1058),
.Y(n_1126)
);

BUFx2_ASAP7_75t_R g1127 ( 
.A(n_1073),
.Y(n_1127)
);

OAI22xp5_ASAP7_75t_L g1128 ( 
.A1(n_1046),
.A2(n_502),
.B1(n_469),
.B2(n_483),
.Y(n_1128)
);

INVx6_ASAP7_75t_L g1129 ( 
.A(n_1069),
.Y(n_1129)
);

INVx4_ASAP7_75t_L g1130 ( 
.A(n_1069),
.Y(n_1130)
);

HB1xp67_ASAP7_75t_L g1131 ( 
.A(n_1052),
.Y(n_1131)
);

CKINVDCx20_ASAP7_75t_R g1132 ( 
.A(n_1027),
.Y(n_1132)
);

NOR2xp33_ASAP7_75t_L g1133 ( 
.A(n_1067),
.B(n_463),
.Y(n_1133)
);

OA21x2_ASAP7_75t_L g1134 ( 
.A1(n_1023),
.A2(n_515),
.B(n_490),
.Y(n_1134)
);

INVx1_ASAP7_75t_L g1135 ( 
.A(n_1040),
.Y(n_1135)
);

INVx2_ASAP7_75t_L g1136 ( 
.A(n_1051),
.Y(n_1136)
);

INVx2_ASAP7_75t_L g1137 ( 
.A(n_1051),
.Y(n_1137)
);

INVx1_ASAP7_75t_L g1138 ( 
.A(n_1057),
.Y(n_1138)
);

AOI22xp33_ASAP7_75t_L g1139 ( 
.A1(n_1079),
.A2(n_516),
.B1(n_507),
.B2(n_494),
.Y(n_1139)
);

INVx2_ASAP7_75t_L g1140 ( 
.A(n_1054),
.Y(n_1140)
);

INVx1_ASAP7_75t_L g1141 ( 
.A(n_1057),
.Y(n_1141)
);

INVx1_ASAP7_75t_L g1142 ( 
.A(n_1054),
.Y(n_1142)
);

BUFx12f_ASAP7_75t_L g1143 ( 
.A(n_1069),
.Y(n_1143)
);

OAI22xp5_ASAP7_75t_L g1144 ( 
.A1(n_1070),
.A2(n_486),
.B1(n_570),
.B2(n_560),
.Y(n_1144)
);

INVx2_ASAP7_75t_L g1145 ( 
.A(n_1054),
.Y(n_1145)
);

INVx2_ASAP7_75t_L g1146 ( 
.A(n_1041),
.Y(n_1146)
);

AND2x4_ASAP7_75t_SL g1147 ( 
.A(n_1098),
.B(n_1058),
.Y(n_1147)
);

NOR2xp33_ASAP7_75t_L g1148 ( 
.A(n_1091),
.B(n_1099),
.Y(n_1148)
);

INVx2_ASAP7_75t_SL g1149 ( 
.A(n_1106),
.Y(n_1149)
);

NAND2xp5_ASAP7_75t_L g1150 ( 
.A(n_1105),
.B(n_1081),
.Y(n_1150)
);

OR2x6_ASAP7_75t_L g1151 ( 
.A(n_1094),
.B(n_1076),
.Y(n_1151)
);

CKINVDCx5p33_ASAP7_75t_R g1152 ( 
.A(n_1132),
.Y(n_1152)
);

INVx2_ASAP7_75t_L g1153 ( 
.A(n_1089),
.Y(n_1153)
);

NOR2xp33_ASAP7_75t_R g1154 ( 
.A(n_1132),
.B(n_1021),
.Y(n_1154)
);

NOR2x1_ASAP7_75t_SL g1155 ( 
.A(n_1124),
.B(n_1079),
.Y(n_1155)
);

NOR3xp33_ASAP7_75t_SL g1156 ( 
.A(n_1100),
.B(n_1074),
.C(n_1053),
.Y(n_1156)
);

OR2x2_ASAP7_75t_L g1157 ( 
.A(n_1097),
.B(n_1078),
.Y(n_1157)
);

NOR2xp33_ASAP7_75t_R g1158 ( 
.A(n_1117),
.B(n_1106),
.Y(n_1158)
);

BUFx4f_ASAP7_75t_SL g1159 ( 
.A(n_1143),
.Y(n_1159)
);

INVx2_ASAP7_75t_L g1160 ( 
.A(n_1136),
.Y(n_1160)
);

INVx1_ASAP7_75t_L g1161 ( 
.A(n_1087),
.Y(n_1161)
);

AO32x2_ASAP7_75t_L g1162 ( 
.A1(n_1092),
.A2(n_1078),
.A3(n_1084),
.B1(n_1085),
.B2(n_1044),
.Y(n_1162)
);

CKINVDCx16_ASAP7_75t_R g1163 ( 
.A(n_1133),
.Y(n_1163)
);

AND2x2_ASAP7_75t_L g1164 ( 
.A(n_1113),
.B(n_1070),
.Y(n_1164)
);

NAND2x1_ASAP7_75t_L g1165 ( 
.A(n_1090),
.B(n_1034),
.Y(n_1165)
);

OR2x2_ASAP7_75t_L g1166 ( 
.A(n_1104),
.B(n_1050),
.Y(n_1166)
);

AND2x2_ASAP7_75t_L g1167 ( 
.A(n_1112),
.B(n_1125),
.Y(n_1167)
);

NAND2xp5_ASAP7_75t_L g1168 ( 
.A(n_1102),
.B(n_1050),
.Y(n_1168)
);

AOI22xp33_ASAP7_75t_L g1169 ( 
.A1(n_1102),
.A2(n_1066),
.B1(n_1080),
.B2(n_1075),
.Y(n_1169)
);

NAND2xp33_ASAP7_75t_R g1170 ( 
.A(n_1134),
.B(n_1041),
.Y(n_1170)
);

O2A1O1Ixp33_ASAP7_75t_L g1171 ( 
.A1(n_1107),
.A2(n_1080),
.B(n_1066),
.C(n_1064),
.Y(n_1171)
);

NAND2xp5_ASAP7_75t_SL g1172 ( 
.A(n_1103),
.B(n_1033),
.Y(n_1172)
);

BUFx6f_ASAP7_75t_L g1173 ( 
.A(n_1122),
.Y(n_1173)
);

NOR2xp33_ASAP7_75t_L g1174 ( 
.A(n_1133),
.B(n_1042),
.Y(n_1174)
);

INVx2_ASAP7_75t_L g1175 ( 
.A(n_1136),
.Y(n_1175)
);

NAND2xp5_ASAP7_75t_SL g1176 ( 
.A(n_1110),
.B(n_1033),
.Y(n_1176)
);

INVx1_ASAP7_75t_L g1177 ( 
.A(n_1138),
.Y(n_1177)
);

INVx2_ASAP7_75t_L g1178 ( 
.A(n_1137),
.Y(n_1178)
);

INVx2_ASAP7_75t_L g1179 ( 
.A(n_1137),
.Y(n_1179)
);

NOR2xp33_ASAP7_75t_R g1180 ( 
.A(n_1126),
.B(n_1042),
.Y(n_1180)
);

INVx1_ASAP7_75t_L g1181 ( 
.A(n_1141),
.Y(n_1181)
);

NAND3xp33_ASAP7_75t_SL g1182 ( 
.A(n_1110),
.B(n_1035),
.C(n_1085),
.Y(n_1182)
);

CKINVDCx5p33_ASAP7_75t_R g1183 ( 
.A(n_1116),
.Y(n_1183)
);

NOR3xp33_ASAP7_75t_SL g1184 ( 
.A(n_1128),
.B(n_1144),
.C(n_1111),
.Y(n_1184)
);

INVx2_ASAP7_75t_L g1185 ( 
.A(n_1095),
.Y(n_1185)
);

INVx2_ASAP7_75t_SL g1186 ( 
.A(n_1126),
.Y(n_1186)
);

OR2x6_ASAP7_75t_L g1187 ( 
.A(n_1129),
.B(n_1035),
.Y(n_1187)
);

AO31x2_ASAP7_75t_L g1188 ( 
.A1(n_1135),
.A2(n_1065),
.A3(n_1061),
.B(n_1038),
.Y(n_1188)
);

AND2x4_ASAP7_75t_L g1189 ( 
.A(n_1131),
.B(n_1044),
.Y(n_1189)
);

AO31x2_ASAP7_75t_L g1190 ( 
.A1(n_1120),
.A2(n_1061),
.A3(n_1059),
.B(n_1077),
.Y(n_1190)
);

INVx2_ASAP7_75t_L g1191 ( 
.A(n_1096),
.Y(n_1191)
);

AND2x2_ASAP7_75t_L g1192 ( 
.A(n_1101),
.B(n_1048),
.Y(n_1192)
);

NAND2xp5_ASAP7_75t_L g1193 ( 
.A(n_1101),
.B(n_1048),
.Y(n_1193)
);

NAND2xp5_ASAP7_75t_L g1194 ( 
.A(n_1093),
.B(n_1049),
.Y(n_1194)
);

CKINVDCx16_ASAP7_75t_R g1195 ( 
.A(n_1130),
.Y(n_1195)
);

OR2x6_ASAP7_75t_L g1196 ( 
.A(n_1122),
.B(n_1049),
.Y(n_1196)
);

AND2x4_ASAP7_75t_SL g1197 ( 
.A(n_1090),
.B(n_570),
.Y(n_1197)
);

NAND2xp5_ASAP7_75t_L g1198 ( 
.A(n_1109),
.B(n_40),
.Y(n_1198)
);

INVx2_ASAP7_75t_SL g1199 ( 
.A(n_1146),
.Y(n_1199)
);

AND2x2_ASAP7_75t_L g1200 ( 
.A(n_1192),
.B(n_1134),
.Y(n_1200)
);

AND2x2_ASAP7_75t_L g1201 ( 
.A(n_1167),
.B(n_1134),
.Y(n_1201)
);

AND2x2_ASAP7_75t_L g1202 ( 
.A(n_1168),
.B(n_1088),
.Y(n_1202)
);

INVx2_ASAP7_75t_L g1203 ( 
.A(n_1160),
.Y(n_1203)
);

INVx2_ASAP7_75t_L g1204 ( 
.A(n_1175),
.Y(n_1204)
);

AND2x2_ASAP7_75t_L g1205 ( 
.A(n_1162),
.B(n_1088),
.Y(n_1205)
);

AND2x4_ASAP7_75t_L g1206 ( 
.A(n_1196),
.B(n_1145),
.Y(n_1206)
);

INVx2_ASAP7_75t_L g1207 ( 
.A(n_1178),
.Y(n_1207)
);

INVx1_ASAP7_75t_L g1208 ( 
.A(n_1161),
.Y(n_1208)
);

AND2x4_ASAP7_75t_L g1209 ( 
.A(n_1196),
.B(n_1145),
.Y(n_1209)
);

OR2x2_ASAP7_75t_L g1210 ( 
.A(n_1166),
.B(n_1088),
.Y(n_1210)
);

OR2x2_ASAP7_75t_L g1211 ( 
.A(n_1150),
.B(n_1121),
.Y(n_1211)
);

INVx2_ASAP7_75t_L g1212 ( 
.A(n_1179),
.Y(n_1212)
);

AND2x4_ASAP7_75t_L g1213 ( 
.A(n_1177),
.B(n_1142),
.Y(n_1213)
);

AND2x2_ASAP7_75t_L g1214 ( 
.A(n_1162),
.B(n_1096),
.Y(n_1214)
);

NAND2xp5_ASAP7_75t_L g1215 ( 
.A(n_1174),
.B(n_1123),
.Y(n_1215)
);

INVx2_ASAP7_75t_L g1216 ( 
.A(n_1185),
.Y(n_1216)
);

INVx2_ASAP7_75t_L g1217 ( 
.A(n_1191),
.Y(n_1217)
);

NAND2xp5_ASAP7_75t_L g1218 ( 
.A(n_1153),
.B(n_1108),
.Y(n_1218)
);

INVx2_ASAP7_75t_L g1219 ( 
.A(n_1181),
.Y(n_1219)
);

INVx1_ASAP7_75t_L g1220 ( 
.A(n_1194),
.Y(n_1220)
);

OR2x2_ASAP7_75t_L g1221 ( 
.A(n_1193),
.B(n_1114),
.Y(n_1221)
);

INVx2_ASAP7_75t_L g1222 ( 
.A(n_1188),
.Y(n_1222)
);

OR2x2_ASAP7_75t_L g1223 ( 
.A(n_1188),
.B(n_1115),
.Y(n_1223)
);

INVx2_ASAP7_75t_L g1224 ( 
.A(n_1188),
.Y(n_1224)
);

INVx5_ASAP7_75t_L g1225 ( 
.A(n_1187),
.Y(n_1225)
);

AOI22xp5_ASAP7_75t_L g1226 ( 
.A1(n_1163),
.A2(n_1139),
.B1(n_1119),
.B2(n_1109),
.Y(n_1226)
);

OR2x2_ASAP7_75t_L g1227 ( 
.A(n_1148),
.B(n_1157),
.Y(n_1227)
);

INVx2_ASAP7_75t_L g1228 ( 
.A(n_1190),
.Y(n_1228)
);

AND2x2_ASAP7_75t_L g1229 ( 
.A(n_1155),
.B(n_1118),
.Y(n_1229)
);

INVx1_ASAP7_75t_L g1230 ( 
.A(n_1199),
.Y(n_1230)
);

AND2x2_ASAP7_75t_L g1231 ( 
.A(n_1169),
.B(n_1189),
.Y(n_1231)
);

OR2x2_ASAP7_75t_L g1232 ( 
.A(n_1198),
.B(n_1140),
.Y(n_1232)
);

INVx1_ASAP7_75t_L g1233 ( 
.A(n_1190),
.Y(n_1233)
);

BUFx2_ASAP7_75t_L g1234 ( 
.A(n_1151),
.Y(n_1234)
);

INVx1_ASAP7_75t_L g1235 ( 
.A(n_1190),
.Y(n_1235)
);

NAND2xp5_ASAP7_75t_L g1236 ( 
.A(n_1176),
.B(n_1119),
.Y(n_1236)
);

INVx1_ASAP7_75t_L g1237 ( 
.A(n_1172),
.Y(n_1237)
);

INVx1_ASAP7_75t_L g1238 ( 
.A(n_1171),
.Y(n_1238)
);

NOR2xp33_ASAP7_75t_L g1239 ( 
.A(n_1164),
.B(n_1127),
.Y(n_1239)
);

INVx1_ASAP7_75t_L g1240 ( 
.A(n_1173),
.Y(n_1240)
);

INVx2_ASAP7_75t_L g1241 ( 
.A(n_1165),
.Y(n_1241)
);

INVx3_ASAP7_75t_L g1242 ( 
.A(n_1187),
.Y(n_1242)
);

OR2x2_ASAP7_75t_L g1243 ( 
.A(n_1182),
.B(n_1149),
.Y(n_1243)
);

AND2x2_ASAP7_75t_L g1244 ( 
.A(n_1184),
.B(n_45),
.Y(n_1244)
);

OR2x6_ASAP7_75t_L g1245 ( 
.A(n_1186),
.B(n_575),
.Y(n_1245)
);

INVx2_ASAP7_75t_L g1246 ( 
.A(n_1197),
.Y(n_1246)
);

AND2x2_ASAP7_75t_L g1247 ( 
.A(n_1156),
.B(n_47),
.Y(n_1247)
);

BUFx2_ASAP7_75t_SL g1248 ( 
.A(n_1158),
.Y(n_1248)
);

AND2x2_ASAP7_75t_L g1249 ( 
.A(n_1195),
.B(n_97),
.Y(n_1249)
);

INVx3_ASAP7_75t_L g1250 ( 
.A(n_1147),
.Y(n_1250)
);

INVx2_ASAP7_75t_L g1251 ( 
.A(n_1219),
.Y(n_1251)
);

AND2x2_ASAP7_75t_L g1252 ( 
.A(n_1231),
.B(n_1152),
.Y(n_1252)
);

BUFx3_ASAP7_75t_L g1253 ( 
.A(n_1250),
.Y(n_1253)
);

AOI221xp5_ASAP7_75t_SL g1254 ( 
.A1(n_1244),
.A2(n_1170),
.B1(n_1180),
.B2(n_1154),
.C(n_1159),
.Y(n_1254)
);

INVxp67_ASAP7_75t_L g1255 ( 
.A(n_1201),
.Y(n_1255)
);

INVx1_ASAP7_75t_L g1256 ( 
.A(n_1208),
.Y(n_1256)
);

INVx2_ASAP7_75t_L g1257 ( 
.A(n_1219),
.Y(n_1257)
);

NAND2xp5_ASAP7_75t_L g1258 ( 
.A(n_1215),
.B(n_1183),
.Y(n_1258)
);

INVx1_ASAP7_75t_L g1259 ( 
.A(n_1220),
.Y(n_1259)
);

OR2x2_ASAP7_75t_L g1260 ( 
.A(n_1227),
.B(n_98),
.Y(n_1260)
);

INVx2_ASAP7_75t_L g1261 ( 
.A(n_1223),
.Y(n_1261)
);

AND2x2_ASAP7_75t_L g1262 ( 
.A(n_1231),
.B(n_294),
.Y(n_1262)
);

INVx2_ASAP7_75t_L g1263 ( 
.A(n_1221),
.Y(n_1263)
);

NAND3xp33_ASAP7_75t_L g1264 ( 
.A(n_1226),
.B(n_105),
.C(n_106),
.Y(n_1264)
);

INVx2_ASAP7_75t_L g1265 ( 
.A(n_1221),
.Y(n_1265)
);

HB1xp67_ASAP7_75t_L g1266 ( 
.A(n_1233),
.Y(n_1266)
);

NAND2xp5_ASAP7_75t_L g1267 ( 
.A(n_1211),
.B(n_107),
.Y(n_1267)
);

INVx1_ASAP7_75t_L g1268 ( 
.A(n_1203),
.Y(n_1268)
);

INVx1_ASAP7_75t_L g1269 ( 
.A(n_1203),
.Y(n_1269)
);

OR2x2_ASAP7_75t_L g1270 ( 
.A(n_1210),
.B(n_109),
.Y(n_1270)
);

INVx1_ASAP7_75t_L g1271 ( 
.A(n_1204),
.Y(n_1271)
);

INVx1_ASAP7_75t_L g1272 ( 
.A(n_1204),
.Y(n_1272)
);

INVx1_ASAP7_75t_L g1273 ( 
.A(n_1207),
.Y(n_1273)
);

AND2x4_ASAP7_75t_L g1274 ( 
.A(n_1229),
.B(n_112),
.Y(n_1274)
);

AND2x2_ASAP7_75t_L g1275 ( 
.A(n_1237),
.B(n_1200),
.Y(n_1275)
);

NOR2xp33_ASAP7_75t_L g1276 ( 
.A(n_1244),
.B(n_116),
.Y(n_1276)
);

INVx2_ASAP7_75t_L g1277 ( 
.A(n_1222),
.Y(n_1277)
);

NAND2xp5_ASAP7_75t_L g1278 ( 
.A(n_1232),
.B(n_118),
.Y(n_1278)
);

INVxp67_ASAP7_75t_L g1279 ( 
.A(n_1238),
.Y(n_1279)
);

HB1xp67_ASAP7_75t_L g1280 ( 
.A(n_1235),
.Y(n_1280)
);

NAND3xp33_ASAP7_75t_L g1281 ( 
.A(n_1236),
.B(n_125),
.C(n_127),
.Y(n_1281)
);

OR2x2_ASAP7_75t_L g1282 ( 
.A(n_1210),
.B(n_128),
.Y(n_1282)
);

NAND3xp33_ASAP7_75t_L g1283 ( 
.A(n_1247),
.B(n_129),
.C(n_130),
.Y(n_1283)
);

INVx3_ASAP7_75t_L g1284 ( 
.A(n_1206),
.Y(n_1284)
);

INVx1_ASAP7_75t_L g1285 ( 
.A(n_1212),
.Y(n_1285)
);

INVx2_ASAP7_75t_L g1286 ( 
.A(n_1224),
.Y(n_1286)
);

INVx2_ASAP7_75t_L g1287 ( 
.A(n_1251),
.Y(n_1287)
);

NAND2xp5_ASAP7_75t_L g1288 ( 
.A(n_1263),
.B(n_1202),
.Y(n_1288)
);

AND2x2_ASAP7_75t_L g1289 ( 
.A(n_1255),
.B(n_1214),
.Y(n_1289)
);

AND2x2_ASAP7_75t_L g1290 ( 
.A(n_1275),
.B(n_1265),
.Y(n_1290)
);

AND2x2_ASAP7_75t_L g1291 ( 
.A(n_1261),
.B(n_1214),
.Y(n_1291)
);

INVx1_ASAP7_75t_L g1292 ( 
.A(n_1256),
.Y(n_1292)
);

HB1xp67_ASAP7_75t_L g1293 ( 
.A(n_1279),
.Y(n_1293)
);

NAND2xp5_ASAP7_75t_SL g1294 ( 
.A(n_1254),
.B(n_1225),
.Y(n_1294)
);

INVx1_ASAP7_75t_L g1295 ( 
.A(n_1257),
.Y(n_1295)
);

INVx3_ASAP7_75t_L g1296 ( 
.A(n_1284),
.Y(n_1296)
);

INVx2_ASAP7_75t_L g1297 ( 
.A(n_1277),
.Y(n_1297)
);

OR2x2_ASAP7_75t_L g1298 ( 
.A(n_1261),
.B(n_1228),
.Y(n_1298)
);

INVx3_ASAP7_75t_L g1299 ( 
.A(n_1284),
.Y(n_1299)
);

INVx2_ASAP7_75t_L g1300 ( 
.A(n_1277),
.Y(n_1300)
);

INVx1_ASAP7_75t_L g1301 ( 
.A(n_1266),
.Y(n_1301)
);

INVx1_ASAP7_75t_L g1302 ( 
.A(n_1259),
.Y(n_1302)
);

AND2x2_ASAP7_75t_L g1303 ( 
.A(n_1268),
.B(n_1205),
.Y(n_1303)
);

AND2x2_ASAP7_75t_L g1304 ( 
.A(n_1269),
.B(n_1205),
.Y(n_1304)
);

AND2x2_ASAP7_75t_L g1305 ( 
.A(n_1271),
.B(n_1272),
.Y(n_1305)
);

INVx2_ASAP7_75t_L g1306 ( 
.A(n_1286),
.Y(n_1306)
);

NOR2xp33_ASAP7_75t_L g1307 ( 
.A(n_1258),
.B(n_1239),
.Y(n_1307)
);

AND2x2_ASAP7_75t_L g1308 ( 
.A(n_1273),
.B(n_1228),
.Y(n_1308)
);

INVx4_ASAP7_75t_L g1309 ( 
.A(n_1274),
.Y(n_1309)
);

INVx2_ASAP7_75t_L g1310 ( 
.A(n_1287),
.Y(n_1310)
);

INVx1_ASAP7_75t_L g1311 ( 
.A(n_1292),
.Y(n_1311)
);

AND2x4_ASAP7_75t_L g1312 ( 
.A(n_1296),
.B(n_1299),
.Y(n_1312)
);

INVx1_ASAP7_75t_L g1313 ( 
.A(n_1293),
.Y(n_1313)
);

INVx2_ASAP7_75t_L g1314 ( 
.A(n_1287),
.Y(n_1314)
);

OR2x6_ASAP7_75t_L g1315 ( 
.A(n_1294),
.B(n_1248),
.Y(n_1315)
);

AOI22xp5_ASAP7_75t_L g1316 ( 
.A1(n_1309),
.A2(n_1264),
.B1(n_1276),
.B2(n_1283),
.Y(n_1316)
);

AOI22xp33_ASAP7_75t_L g1317 ( 
.A1(n_1307),
.A2(n_1276),
.B1(n_1281),
.B2(n_1262),
.Y(n_1317)
);

NAND2xp5_ASAP7_75t_L g1318 ( 
.A(n_1288),
.B(n_1285),
.Y(n_1318)
);

NAND2xp5_ASAP7_75t_L g1319 ( 
.A(n_1290),
.B(n_1252),
.Y(n_1319)
);

OAI322xp33_ASAP7_75t_L g1320 ( 
.A1(n_1302),
.A2(n_1247),
.A3(n_1260),
.B1(n_1282),
.B2(n_1270),
.C1(n_1243),
.C2(n_1230),
.Y(n_1320)
);

NOR2xp67_ASAP7_75t_L g1321 ( 
.A(n_1296),
.B(n_1280),
.Y(n_1321)
);

NAND2xp5_ASAP7_75t_L g1322 ( 
.A(n_1313),
.B(n_1305),
.Y(n_1322)
);

NAND3xp33_ASAP7_75t_L g1323 ( 
.A(n_1317),
.B(n_1301),
.C(n_1267),
.Y(n_1323)
);

AOI21xp33_ASAP7_75t_L g1324 ( 
.A1(n_1315),
.A2(n_1278),
.B(n_1301),
.Y(n_1324)
);

OAI21xp5_ASAP7_75t_SL g1325 ( 
.A1(n_1316),
.A2(n_1239),
.B(n_1249),
.Y(n_1325)
);

INVxp67_ASAP7_75t_SL g1326 ( 
.A(n_1321),
.Y(n_1326)
);

INVx2_ASAP7_75t_L g1327 ( 
.A(n_1310),
.Y(n_1327)
);

AO22x2_ASAP7_75t_L g1328 ( 
.A1(n_1311),
.A2(n_1299),
.B1(n_1296),
.B2(n_1295),
.Y(n_1328)
);

AOI22xp5_ASAP7_75t_L g1329 ( 
.A1(n_1319),
.A2(n_1242),
.B1(n_1234),
.B2(n_1253),
.Y(n_1329)
);

O2A1O1Ixp33_ASAP7_75t_L g1330 ( 
.A1(n_1325),
.A2(n_1320),
.B(n_1245),
.C(n_1318),
.Y(n_1330)
);

OAI22xp5_ASAP7_75t_L g1331 ( 
.A1(n_1323),
.A2(n_1225),
.B1(n_1312),
.B2(n_1289),
.Y(n_1331)
);

OAI22xp33_ASAP7_75t_SL g1332 ( 
.A1(n_1326),
.A2(n_1312),
.B1(n_1314),
.B2(n_1245),
.Y(n_1332)
);

INVx2_ASAP7_75t_L g1333 ( 
.A(n_1328),
.Y(n_1333)
);

INVx2_ASAP7_75t_L g1334 ( 
.A(n_1328),
.Y(n_1334)
);

OAI21xp5_ASAP7_75t_SL g1335 ( 
.A1(n_1329),
.A2(n_1250),
.B(n_1291),
.Y(n_1335)
);

INVx1_ASAP7_75t_L g1336 ( 
.A(n_1322),
.Y(n_1336)
);

AND2x2_ASAP7_75t_L g1337 ( 
.A(n_1327),
.B(n_1303),
.Y(n_1337)
);

OAI21xp33_ASAP7_75t_SL g1338 ( 
.A1(n_1324),
.A2(n_1304),
.B(n_1308),
.Y(n_1338)
);

OR2x2_ASAP7_75t_L g1339 ( 
.A(n_1336),
.B(n_1298),
.Y(n_1339)
);

NOR3xp33_ASAP7_75t_L g1340 ( 
.A(n_1330),
.B(n_1240),
.C(n_1246),
.Y(n_1340)
);

AOI221xp5_ASAP7_75t_L g1341 ( 
.A1(n_1331),
.A2(n_1308),
.B1(n_1213),
.B2(n_1306),
.C(n_1300),
.Y(n_1341)
);

HB1xp67_ASAP7_75t_L g1342 ( 
.A(n_1333),
.Y(n_1342)
);

AOI221xp5_ASAP7_75t_L g1343 ( 
.A1(n_1338),
.A2(n_1213),
.B1(n_1306),
.B2(n_1300),
.C(n_1297),
.Y(n_1343)
);

O2A1O1Ixp33_ASAP7_75t_L g1344 ( 
.A1(n_1332),
.A2(n_1246),
.B(n_1241),
.C(n_1218),
.Y(n_1344)
);

NOR3xp33_ASAP7_75t_L g1345 ( 
.A(n_1342),
.B(n_1334),
.C(n_1335),
.Y(n_1345)
);

AND2x2_ASAP7_75t_L g1346 ( 
.A(n_1340),
.B(n_1337),
.Y(n_1346)
);

INVx1_ASAP7_75t_L g1347 ( 
.A(n_1339),
.Y(n_1347)
);

NAND4xp25_ASAP7_75t_L g1348 ( 
.A(n_1345),
.B(n_1341),
.C(n_1344),
.D(n_1343),
.Y(n_1348)
);

INVx1_ASAP7_75t_L g1349 ( 
.A(n_1347),
.Y(n_1349)
);

NAND3xp33_ASAP7_75t_L g1350 ( 
.A(n_1346),
.B(n_1209),
.C(n_1217),
.Y(n_1350)
);

AOI22xp5_ASAP7_75t_L g1351 ( 
.A1(n_1348),
.A2(n_1280),
.B1(n_1216),
.B2(n_1286),
.Y(n_1351)
);

CKINVDCx16_ASAP7_75t_R g1352 ( 
.A(n_1350),
.Y(n_1352)
);

OR2x2_ASAP7_75t_L g1353 ( 
.A(n_1349),
.B(n_138),
.Y(n_1353)
);

AND2x2_ASAP7_75t_L g1354 ( 
.A(n_1352),
.B(n_142),
.Y(n_1354)
);

INVx2_ASAP7_75t_L g1355 ( 
.A(n_1353),
.Y(n_1355)
);

NAND2xp5_ASAP7_75t_L g1356 ( 
.A(n_1351),
.B(n_150),
.Y(n_1356)
);

BUFx6f_ASAP7_75t_L g1357 ( 
.A(n_1354),
.Y(n_1357)
);

INVx1_ASAP7_75t_SL g1358 ( 
.A(n_1355),
.Y(n_1358)
);

HB1xp67_ASAP7_75t_L g1359 ( 
.A(n_1356),
.Y(n_1359)
);

INVxp67_ASAP7_75t_SL g1360 ( 
.A(n_1357),
.Y(n_1360)
);

XOR2xp5_ASAP7_75t_L g1361 ( 
.A(n_1359),
.B(n_152),
.Y(n_1361)
);

INVx1_ASAP7_75t_L g1362 ( 
.A(n_1358),
.Y(n_1362)
);

OAI31xp33_ASAP7_75t_L g1363 ( 
.A1(n_1362),
.A2(n_158),
.A3(n_164),
.B(n_170),
.Y(n_1363)
);

BUFx2_ASAP7_75t_L g1364 ( 
.A(n_1360),
.Y(n_1364)
);

HB1xp67_ASAP7_75t_L g1365 ( 
.A(n_1361),
.Y(n_1365)
);

AOI22xp5_ASAP7_75t_L g1366 ( 
.A1(n_1365),
.A2(n_192),
.B1(n_195),
.B2(n_199),
.Y(n_1366)
);

OAI22xp5_ASAP7_75t_L g1367 ( 
.A1(n_1363),
.A2(n_210),
.B1(n_215),
.B2(n_217),
.Y(n_1367)
);

NAND3xp33_ASAP7_75t_L g1368 ( 
.A(n_1364),
.B(n_219),
.C(n_221),
.Y(n_1368)
);

AOI222xp33_ASAP7_75t_L g1369 ( 
.A1(n_1367),
.A2(n_288),
.B1(n_223),
.B2(n_227),
.C1(n_232),
.C2(n_233),
.Y(n_1369)
);

INVx1_ASAP7_75t_L g1370 ( 
.A(n_1368),
.Y(n_1370)
);

AOI21xp5_ASAP7_75t_L g1371 ( 
.A1(n_1370),
.A2(n_1366),
.B(n_234),
.Y(n_1371)
);

AO22x2_ASAP7_75t_L g1372 ( 
.A1(n_1369),
.A2(n_222),
.B1(n_235),
.B2(n_236),
.Y(n_1372)
);

AOI22xp33_ASAP7_75t_L g1373 ( 
.A1(n_1372),
.A2(n_237),
.B1(n_239),
.B2(n_242),
.Y(n_1373)
);

AOI222xp33_ASAP7_75t_L g1374 ( 
.A1(n_1371),
.A2(n_244),
.B1(n_246),
.B2(n_247),
.C1(n_251),
.C2(n_257),
.Y(n_1374)
);

AOI221x1_ASAP7_75t_L g1375 ( 
.A1(n_1374),
.A2(n_258),
.B1(n_259),
.B2(n_261),
.C(n_265),
.Y(n_1375)
);

AOI211xp5_ASAP7_75t_L g1376 ( 
.A1(n_1375),
.A2(n_1373),
.B(n_266),
.C(n_271),
.Y(n_1376)
);


endmodule