module fake_jpeg_25200_n_310 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_310);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_310;

wire n_253;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_18;
wire n_20;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_208;
wire n_308;
wire n_297;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVx6_ASAP7_75t_L g16 ( 
.A(n_9),
.Y(n_16)
);

BUFx12f_ASAP7_75t_L g17 ( 
.A(n_0),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_9),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_5),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_5),
.Y(n_20)
);

BUFx16f_ASAP7_75t_L g21 ( 
.A(n_13),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_7),
.Y(n_22)
);

BUFx3_ASAP7_75t_L g23 ( 
.A(n_10),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_5),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_14),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_0),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_8),
.Y(n_27)
);

INVx8_ASAP7_75t_L g28 ( 
.A(n_10),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_1),
.Y(n_29)
);

INVx5_ASAP7_75t_L g30 ( 
.A(n_0),
.Y(n_30)
);

CKINVDCx16_ASAP7_75t_R g31 ( 
.A(n_11),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_12),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_0),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_28),
.Y(n_34)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_34),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_17),
.Y(n_35)
);

INVx6_ASAP7_75t_L g45 ( 
.A(n_35),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_17),
.Y(n_36)
);

INVx6_ASAP7_75t_L g60 ( 
.A(n_36),
.Y(n_60)
);

CKINVDCx16_ASAP7_75t_R g37 ( 
.A(n_17),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_37),
.B(n_19),
.Y(n_55)
);

INVx2_ASAP7_75t_L g38 ( 
.A(n_17),
.Y(n_38)
);

INVx2_ASAP7_75t_L g46 ( 
.A(n_38),
.Y(n_46)
);

INVx2_ASAP7_75t_SL g39 ( 
.A(n_30),
.Y(n_39)
);

BUFx2_ASAP7_75t_L g43 ( 
.A(n_39),
.Y(n_43)
);

INVx3_ASAP7_75t_L g40 ( 
.A(n_17),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_40),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_17),
.Y(n_41)
);

INVx2_ASAP7_75t_L g49 ( 
.A(n_41),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_30),
.Y(n_42)
);

INVx2_ASAP7_75t_L g53 ( 
.A(n_42),
.Y(n_53)
);

INVx8_ASAP7_75t_L g44 ( 
.A(n_42),
.Y(n_44)
);

INVx8_ASAP7_75t_L g89 ( 
.A(n_44),
.Y(n_89)
);

BUFx2_ASAP7_75t_L g47 ( 
.A(n_39),
.Y(n_47)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_47),
.Y(n_65)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_38),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_51),
.B(n_54),
.Y(n_78)
);

INVx3_ASAP7_75t_L g52 ( 
.A(n_42),
.Y(n_52)
);

INVx1_ASAP7_75t_SL g86 ( 
.A(n_52),
.Y(n_86)
);

INVx6_ASAP7_75t_SL g54 ( 
.A(n_39),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_L g74 ( 
.A(n_55),
.B(n_62),
.Y(n_74)
);

AOI22xp33_ASAP7_75t_L g56 ( 
.A1(n_39),
.A2(n_16),
.B1(n_28),
.B2(n_30),
.Y(n_56)
);

OA22x2_ASAP7_75t_L g77 ( 
.A1(n_56),
.A2(n_16),
.B1(n_28),
.B2(n_40),
.Y(n_77)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_38),
.Y(n_57)
);

INVx2_ASAP7_75t_L g63 ( 
.A(n_57),
.Y(n_63)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_40),
.Y(n_58)
);

INVx4_ASAP7_75t_L g84 ( 
.A(n_58),
.Y(n_84)
);

INVx2_ASAP7_75t_L g59 ( 
.A(n_35),
.Y(n_59)
);

INVx2_ASAP7_75t_L g82 ( 
.A(n_59),
.Y(n_82)
);

AND2x2_ASAP7_75t_L g61 ( 
.A(n_42),
.B(n_24),
.Y(n_61)
);

A2O1A1Ixp33_ASAP7_75t_L g69 ( 
.A1(n_61),
.A2(n_37),
.B(n_34),
.C(n_39),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_L g62 ( 
.A(n_37),
.B(n_26),
.Y(n_62)
);

INVx2_ASAP7_75t_L g64 ( 
.A(n_46),
.Y(n_64)
);

INVx2_ASAP7_75t_L g102 ( 
.A(n_64),
.Y(n_102)
);

INVx3_ASAP7_75t_L g66 ( 
.A(n_50),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_66),
.B(n_67),
.Y(n_96)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_62),
.Y(n_67)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_43),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_68),
.B(n_72),
.Y(n_105)
);

OAI21xp5_ASAP7_75t_L g90 ( 
.A1(n_69),
.A2(n_61),
.B(n_53),
.Y(n_90)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_46),
.Y(n_70)
);

INVx2_ASAP7_75t_L g107 ( 
.A(n_70),
.Y(n_107)
);

XNOR2xp5_ASAP7_75t_L g71 ( 
.A(n_48),
.B(n_34),
.Y(n_71)
);

XNOR2xp5_ASAP7_75t_L g115 ( 
.A(n_71),
.B(n_29),
.Y(n_115)
);

INVx3_ASAP7_75t_L g72 ( 
.A(n_50),
.Y(n_72)
);

CKINVDCx20_ASAP7_75t_R g73 ( 
.A(n_58),
.Y(n_73)
);

CKINVDCx20_ASAP7_75t_R g101 ( 
.A(n_73),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_L g75 ( 
.A(n_48),
.B(n_18),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_SL g103 ( 
.A(n_75),
.B(n_80),
.Y(n_103)
);

INVx3_ASAP7_75t_L g76 ( 
.A(n_44),
.Y(n_76)
);

BUFx2_ASAP7_75t_L g92 ( 
.A(n_76),
.Y(n_92)
);

AND2x2_ASAP7_75t_L g95 ( 
.A(n_77),
.B(n_83),
.Y(n_95)
);

INVx5_ASAP7_75t_L g79 ( 
.A(n_54),
.Y(n_79)
);

INVx2_ASAP7_75t_SL g104 ( 
.A(n_79),
.Y(n_104)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_43),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_SL g81 ( 
.A(n_57),
.B(n_20),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_SL g109 ( 
.A(n_81),
.B(n_18),
.Y(n_109)
);

OA22x2_ASAP7_75t_L g83 ( 
.A1(n_52),
.A2(n_16),
.B1(n_28),
.B2(n_26),
.Y(n_83)
);

BUFx2_ASAP7_75t_L g85 ( 
.A(n_47),
.Y(n_85)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_85),
.Y(n_93)
);

HB1xp67_ASAP7_75t_L g87 ( 
.A(n_49),
.Y(n_87)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_87),
.Y(n_108)
);

OA22x2_ASAP7_75t_L g88 ( 
.A1(n_61),
.A2(n_16),
.B1(n_27),
.B2(n_26),
.Y(n_88)
);

AND2x2_ASAP7_75t_L g98 ( 
.A(n_88),
.B(n_25),
.Y(n_98)
);

XOR2xp5_ASAP7_75t_L g140 ( 
.A(n_90),
.B(n_115),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_L g91 ( 
.A(n_71),
.B(n_53),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_SL g143 ( 
.A(n_91),
.B(n_97),
.Y(n_143)
);

OAI22xp5_ASAP7_75t_L g94 ( 
.A1(n_74),
.A2(n_45),
.B1(n_60),
.B2(n_49),
.Y(n_94)
);

AOI22xp5_ASAP7_75t_L g118 ( 
.A1(n_94),
.A2(n_100),
.B1(n_110),
.B2(n_66),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_L g97 ( 
.A(n_88),
.B(n_59),
.Y(n_97)
);

AOI22xp5_ASAP7_75t_SL g123 ( 
.A1(n_98),
.A2(n_84),
.B1(n_86),
.B2(n_29),
.Y(n_123)
);

OAI21xp5_ASAP7_75t_L g99 ( 
.A1(n_69),
.A2(n_88),
.B(n_78),
.Y(n_99)
);

AOI21xp5_ASAP7_75t_L g124 ( 
.A1(n_99),
.A2(n_32),
.B(n_31),
.Y(n_124)
);

OAI22xp5_ASAP7_75t_L g100 ( 
.A1(n_77),
.A2(n_45),
.B1(n_60),
.B2(n_29),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_L g106 ( 
.A(n_64),
.B(n_41),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g137 ( 
.A(n_106),
.B(n_109),
.Y(n_137)
);

OAI22xp5_ASAP7_75t_SL g110 ( 
.A1(n_77),
.A2(n_70),
.B1(n_63),
.B2(n_83),
.Y(n_110)
);

AOI22xp33_ASAP7_75t_SL g111 ( 
.A1(n_79),
.A2(n_18),
.B1(n_32),
.B2(n_33),
.Y(n_111)
);

OAI22xp5_ASAP7_75t_L g134 ( 
.A1(n_111),
.A2(n_31),
.B1(n_27),
.B2(n_22),
.Y(n_134)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_85),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_L g145 ( 
.A(n_112),
.B(n_114),
.Y(n_145)
);

CKINVDCx14_ASAP7_75t_R g113 ( 
.A(n_83),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_L g142 ( 
.A(n_113),
.B(n_41),
.Y(n_142)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_89),
.Y(n_114)
);

INVx2_ASAP7_75t_L g116 ( 
.A(n_82),
.Y(n_116)
);

INVx2_ASAP7_75t_L g129 ( 
.A(n_116),
.Y(n_129)
);

OAI22xp5_ASAP7_75t_SL g117 ( 
.A1(n_113),
.A2(n_89),
.B1(n_76),
.B2(n_72),
.Y(n_117)
);

AOI22xp5_ASAP7_75t_L g151 ( 
.A1(n_117),
.A2(n_119),
.B1(n_133),
.B2(n_138),
.Y(n_151)
);

AOI22xp33_ASAP7_75t_L g147 ( 
.A1(n_118),
.A2(n_130),
.B1(n_131),
.B2(n_104),
.Y(n_147)
);

OAI22xp5_ASAP7_75t_L g119 ( 
.A1(n_97),
.A2(n_84),
.B1(n_86),
.B2(n_65),
.Y(n_119)
);

BUFx3_ASAP7_75t_L g120 ( 
.A(n_116),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_L g158 ( 
.A(n_120),
.B(n_121),
.Y(n_158)
);

INVx3_ASAP7_75t_L g121 ( 
.A(n_92),
.Y(n_121)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_106),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_SL g148 ( 
.A(n_122),
.B(n_125),
.Y(n_148)
);

OAI21xp5_ASAP7_75t_SL g163 ( 
.A1(n_123),
.A2(n_124),
.B(n_134),
.Y(n_163)
);

CKINVDCx14_ASAP7_75t_R g125 ( 
.A(n_105),
.Y(n_125)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_105),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_SL g156 ( 
.A(n_126),
.B(n_127),
.Y(n_156)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_92),
.Y(n_127)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_92),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_SL g174 ( 
.A(n_128),
.B(n_132),
.Y(n_174)
);

OAI22xp33_ASAP7_75t_SL g130 ( 
.A1(n_98),
.A2(n_20),
.B1(n_33),
.B2(n_22),
.Y(n_130)
);

AOI22xp33_ASAP7_75t_L g131 ( 
.A1(n_99),
.A2(n_25),
.B1(n_19),
.B2(n_24),
.Y(n_131)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_94),
.Y(n_132)
);

OAI22xp5_ASAP7_75t_L g133 ( 
.A1(n_90),
.A2(n_32),
.B1(n_22),
.B2(n_27),
.Y(n_133)
);

INVx2_ASAP7_75t_L g135 ( 
.A(n_102),
.Y(n_135)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_135),
.Y(n_149)
);

MAJIxp5_ASAP7_75t_L g136 ( 
.A(n_91),
.B(n_36),
.C(n_35),
.Y(n_136)
);

MAJIxp5_ASAP7_75t_L g146 ( 
.A(n_136),
.B(n_100),
.C(n_98),
.Y(n_146)
);

OAI22xp5_ASAP7_75t_L g138 ( 
.A1(n_110),
.A2(n_41),
.B1(n_36),
.B2(n_35),
.Y(n_138)
);

INVx2_ASAP7_75t_L g139 ( 
.A(n_102),
.Y(n_139)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_139),
.Y(n_159)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_96),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_L g150 ( 
.A(n_141),
.B(n_103),
.Y(n_150)
);

CKINVDCx14_ASAP7_75t_R g153 ( 
.A(n_142),
.Y(n_153)
);

BUFx2_ASAP7_75t_L g144 ( 
.A(n_107),
.Y(n_144)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_144),
.Y(n_162)
);

MAJIxp5_ASAP7_75t_L g193 ( 
.A(n_146),
.B(n_154),
.C(n_25),
.Y(n_193)
);

OAI22xp5_ASAP7_75t_L g178 ( 
.A1(n_147),
.A2(n_165),
.B1(n_123),
.B2(n_128),
.Y(n_178)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_150),
.Y(n_180)
);

CKINVDCx16_ASAP7_75t_R g152 ( 
.A(n_145),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_L g199 ( 
.A(n_152),
.B(n_164),
.Y(n_199)
);

MAJIxp5_ASAP7_75t_L g154 ( 
.A(n_140),
.B(n_115),
.C(n_96),
.Y(n_154)
);

AOI22xp5_ASAP7_75t_L g155 ( 
.A1(n_132),
.A2(n_95),
.B1(n_103),
.B2(n_114),
.Y(n_155)
);

OAI22xp5_ASAP7_75t_SL g192 ( 
.A1(n_155),
.A2(n_161),
.B1(n_176),
.B2(n_129),
.Y(n_192)
);

XOR2xp5_ASAP7_75t_L g157 ( 
.A(n_140),
.B(n_95),
.Y(n_157)
);

XOR2xp5_ASAP7_75t_L g185 ( 
.A(n_157),
.B(n_21),
.Y(n_185)
);

XNOR2xp5_ASAP7_75t_L g160 ( 
.A(n_136),
.B(n_109),
.Y(n_160)
);

XNOR2xp5_ASAP7_75t_L g182 ( 
.A(n_160),
.B(n_175),
.Y(n_182)
);

AOI22xp5_ASAP7_75t_L g161 ( 
.A1(n_138),
.A2(n_95),
.B1(n_101),
.B2(n_108),
.Y(n_161)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_144),
.Y(n_164)
);

AOI22xp33_ASAP7_75t_SL g165 ( 
.A1(n_121),
.A2(n_104),
.B1(n_101),
.B2(n_112),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_L g166 ( 
.A(n_143),
.B(n_107),
.Y(n_166)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_166),
.Y(n_181)
);

AOI21xp5_ASAP7_75t_L g167 ( 
.A1(n_117),
.A2(n_93),
.B(n_108),
.Y(n_167)
);

OAI21xp5_ASAP7_75t_SL g183 ( 
.A1(n_167),
.A2(n_133),
.B(n_127),
.Y(n_183)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_144),
.Y(n_168)
);

OAI21xp5_ASAP7_75t_SL g186 ( 
.A1(n_168),
.A2(n_170),
.B(n_172),
.Y(n_186)
);

CKINVDCx14_ASAP7_75t_R g169 ( 
.A(n_119),
.Y(n_169)
);

AOI22xp5_ASAP7_75t_SL g197 ( 
.A1(n_169),
.A2(n_21),
.B1(n_23),
.B2(n_24),
.Y(n_197)
);

AOI22xp5_ASAP7_75t_SL g170 ( 
.A1(n_141),
.A2(n_104),
.B1(n_93),
.B2(n_23),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_L g171 ( 
.A(n_143),
.B(n_122),
.Y(n_171)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_171),
.Y(n_184)
);

NAND3xp33_ASAP7_75t_L g172 ( 
.A(n_124),
.B(n_11),
.C(n_15),
.Y(n_172)
);

CKINVDCx20_ASAP7_75t_R g173 ( 
.A(n_135),
.Y(n_173)
);

CKINVDCx20_ASAP7_75t_R g187 ( 
.A(n_173),
.Y(n_187)
);

XNOR2xp5_ASAP7_75t_L g175 ( 
.A(n_137),
.B(n_21),
.Y(n_175)
);

AOI22xp5_ASAP7_75t_L g176 ( 
.A1(n_118),
.A2(n_36),
.B1(n_25),
.B2(n_24),
.Y(n_176)
);

NOR2xp33_ASAP7_75t_SL g177 ( 
.A(n_126),
.B(n_23),
.Y(n_177)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_177),
.Y(n_195)
);

AOI22xp5_ASAP7_75t_L g226 ( 
.A1(n_178),
.A2(n_192),
.B1(n_194),
.B2(n_198),
.Y(n_226)
);

INVx6_ASAP7_75t_L g179 ( 
.A(n_158),
.Y(n_179)
);

NOR2xp33_ASAP7_75t_L g213 ( 
.A(n_179),
.B(n_204),
.Y(n_213)
);

OAI21xp5_ASAP7_75t_L g211 ( 
.A1(n_183),
.A2(n_190),
.B(n_159),
.Y(n_211)
);

XNOR2xp5_ASAP7_75t_L g209 ( 
.A(n_185),
.B(n_203),
.Y(n_209)
);

INVxp67_ASAP7_75t_L g188 ( 
.A(n_174),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_L g206 ( 
.A(n_188),
.B(n_189),
.Y(n_206)
);

INVxp67_ASAP7_75t_L g189 ( 
.A(n_170),
.Y(n_189)
);

AOI22xp33_ASAP7_75t_SL g190 ( 
.A1(n_173),
.A2(n_168),
.B1(n_164),
.B2(n_162),
.Y(n_190)
);

XOR2xp5_ASAP7_75t_L g191 ( 
.A(n_157),
.B(n_21),
.Y(n_191)
);

MAJIxp5_ASAP7_75t_L g229 ( 
.A(n_191),
.B(n_193),
.C(n_196),
.Y(n_229)
);

OAI22xp5_ASAP7_75t_SL g194 ( 
.A1(n_161),
.A2(n_129),
.B1(n_139),
.B2(n_120),
.Y(n_194)
);

XOR2xp5_ASAP7_75t_L g196 ( 
.A(n_154),
.B(n_160),
.Y(n_196)
);

INVx1_ASAP7_75t_SL g218 ( 
.A(n_197),
.Y(n_218)
);

OAI22xp5_ASAP7_75t_SL g198 ( 
.A1(n_151),
.A2(n_19),
.B1(n_21),
.B2(n_3),
.Y(n_198)
);

OA22x2_ASAP7_75t_L g200 ( 
.A1(n_167),
.A2(n_19),
.B1(n_2),
.B2(n_3),
.Y(n_200)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_200),
.Y(n_208)
);

INVx4_ASAP7_75t_L g201 ( 
.A(n_162),
.Y(n_201)
);

INVx2_ASAP7_75t_L g217 ( 
.A(n_201),
.Y(n_217)
);

OAI21xp5_ASAP7_75t_SL g202 ( 
.A1(n_163),
.A2(n_155),
.B(n_153),
.Y(n_202)
);

AOI21xp5_ASAP7_75t_L g207 ( 
.A1(n_202),
.A2(n_163),
.B(n_151),
.Y(n_207)
);

XNOR2xp5_ASAP7_75t_L g203 ( 
.A(n_175),
.B(n_15),
.Y(n_203)
);

INVxp33_ASAP7_75t_L g204 ( 
.A(n_156),
.Y(n_204)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_148),
.Y(n_205)
);

NAND2xp5_ASAP7_75t_SL g222 ( 
.A(n_205),
.B(n_150),
.Y(n_222)
);

XNOR2xp5_ASAP7_75t_SL g247 ( 
.A(n_207),
.B(n_203),
.Y(n_247)
);

NAND2xp5_ASAP7_75t_L g210 ( 
.A(n_188),
.B(n_171),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_L g239 ( 
.A(n_210),
.B(n_212),
.Y(n_239)
);

CKINVDCx14_ASAP7_75t_R g230 ( 
.A(n_211),
.Y(n_230)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_199),
.Y(n_212)
);

NAND2xp5_ASAP7_75t_L g214 ( 
.A(n_184),
.B(n_166),
.Y(n_214)
);

CKINVDCx20_ASAP7_75t_R g237 ( 
.A(n_214),
.Y(n_237)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_194),
.Y(n_215)
);

NOR2xp33_ASAP7_75t_L g235 ( 
.A(n_215),
.B(n_221),
.Y(n_235)
);

NOR2xp33_ASAP7_75t_L g216 ( 
.A(n_204),
.B(n_179),
.Y(n_216)
);

CKINVDCx14_ASAP7_75t_R g242 ( 
.A(n_216),
.Y(n_242)
);

CKINVDCx16_ASAP7_75t_R g219 ( 
.A(n_183),
.Y(n_219)
);

NAND2xp5_ASAP7_75t_SL g236 ( 
.A(n_219),
.B(n_222),
.Y(n_236)
);

HB1xp67_ASAP7_75t_L g220 ( 
.A(n_202),
.Y(n_220)
);

CKINVDCx20_ASAP7_75t_R g244 ( 
.A(n_220),
.Y(n_244)
);

AOI21xp5_ASAP7_75t_L g221 ( 
.A1(n_189),
.A2(n_159),
.B(n_149),
.Y(n_221)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_187),
.Y(n_223)
);

NOR2xp33_ASAP7_75t_L g238 ( 
.A(n_223),
.B(n_225),
.Y(n_238)
);

OAI21xp5_ASAP7_75t_L g224 ( 
.A1(n_181),
.A2(n_146),
.B(n_149),
.Y(n_224)
);

XNOR2xp5_ASAP7_75t_L g234 ( 
.A(n_224),
.B(n_182),
.Y(n_234)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_200),
.Y(n_225)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_200),
.Y(n_227)
);

OAI22xp5_ASAP7_75t_L g241 ( 
.A1(n_227),
.A2(n_197),
.B1(n_176),
.B2(n_200),
.Y(n_241)
);

INVx2_ASAP7_75t_SL g228 ( 
.A(n_201),
.Y(n_228)
);

INVx2_ASAP7_75t_L g231 ( 
.A(n_228),
.Y(n_231)
);

MAJIxp5_ASAP7_75t_L g232 ( 
.A(n_229),
.B(n_193),
.C(n_196),
.Y(n_232)
);

MAJIxp5_ASAP7_75t_L g249 ( 
.A(n_232),
.B(n_233),
.C(n_240),
.Y(n_249)
);

MAJIxp5_ASAP7_75t_L g233 ( 
.A(n_229),
.B(n_224),
.C(n_182),
.Y(n_233)
);

XNOR2xp5_ASAP7_75t_L g259 ( 
.A(n_234),
.B(n_247),
.Y(n_259)
);

MAJIxp5_ASAP7_75t_L g240 ( 
.A(n_209),
.B(n_185),
.C(n_191),
.Y(n_240)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_241),
.Y(n_251)
);

MAJIxp5_ASAP7_75t_L g243 ( 
.A(n_209),
.B(n_211),
.C(n_207),
.Y(n_243)
);

NAND2xp5_ASAP7_75t_L g257 ( 
.A(n_243),
.B(n_245),
.Y(n_257)
);

MAJIxp5_ASAP7_75t_L g245 ( 
.A(n_210),
.B(n_180),
.C(n_192),
.Y(n_245)
);

AOI22xp5_ASAP7_75t_L g246 ( 
.A1(n_215),
.A2(n_198),
.B1(n_195),
.B2(n_186),
.Y(n_246)
);

OAI22xp5_ASAP7_75t_SL g263 ( 
.A1(n_246),
.A2(n_218),
.B1(n_217),
.B2(n_3),
.Y(n_263)
);

OAI221xp5_ASAP7_75t_SL g248 ( 
.A1(n_214),
.A2(n_15),
.B1(n_14),
.B2(n_13),
.C(n_12),
.Y(n_248)
);

OAI22xp5_ASAP7_75t_L g252 ( 
.A1(n_248),
.A2(n_208),
.B1(n_227),
.B2(n_225),
.Y(n_252)
);

HB1xp67_ASAP7_75t_L g250 ( 
.A(n_245),
.Y(n_250)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_250),
.Y(n_268)
);

NOR2xp33_ASAP7_75t_L g266 ( 
.A(n_252),
.B(n_253),
.Y(n_266)
);

NOR2xp33_ASAP7_75t_L g253 ( 
.A(n_244),
.B(n_213),
.Y(n_253)
);

AOI22xp5_ASAP7_75t_L g254 ( 
.A1(n_230),
.A2(n_208),
.B1(n_226),
.B2(n_228),
.Y(n_254)
);

OAI22xp5_ASAP7_75t_SL g276 ( 
.A1(n_254),
.A2(n_255),
.B1(n_1),
.B2(n_2),
.Y(n_276)
);

AOI22xp5_ASAP7_75t_L g255 ( 
.A1(n_235),
.A2(n_226),
.B1(n_228),
.B2(n_221),
.Y(n_255)
);

NOR2xp33_ASAP7_75t_SL g256 ( 
.A(n_236),
.B(n_212),
.Y(n_256)
);

XNOR2xp5_ASAP7_75t_L g269 ( 
.A(n_256),
.B(n_258),
.Y(n_269)
);

AOI21xp5_ASAP7_75t_L g258 ( 
.A1(n_238),
.A2(n_206),
.B(n_218),
.Y(n_258)
);

XNOR2xp5_ASAP7_75t_L g260 ( 
.A(n_234),
.B(n_206),
.Y(n_260)
);

MAJIxp5_ASAP7_75t_L g264 ( 
.A(n_260),
.B(n_233),
.C(n_232),
.Y(n_264)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_239),
.Y(n_261)
);

AOI22xp5_ASAP7_75t_SL g270 ( 
.A1(n_261),
.A2(n_237),
.B1(n_231),
.B2(n_247),
.Y(n_270)
);

NOR2xp33_ASAP7_75t_L g262 ( 
.A(n_242),
.B(n_217),
.Y(n_262)
);

AOI22xp5_ASAP7_75t_L g265 ( 
.A1(n_262),
.A2(n_263),
.B1(n_231),
.B2(n_237),
.Y(n_265)
);

XNOR2xp5_ASAP7_75t_L g279 ( 
.A(n_264),
.B(n_270),
.Y(n_279)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_265),
.Y(n_281)
);

OAI22xp5_ASAP7_75t_SL g267 ( 
.A1(n_251),
.A2(n_246),
.B1(n_243),
.B2(n_239),
.Y(n_267)
);

AOI22xp5_ASAP7_75t_L g284 ( 
.A1(n_267),
.A2(n_276),
.B1(n_260),
.B2(n_259),
.Y(n_284)
);

MAJIxp5_ASAP7_75t_L g271 ( 
.A(n_249),
.B(n_240),
.C(n_14),
.Y(n_271)
);

OR2x2_ASAP7_75t_L g277 ( 
.A(n_271),
.B(n_272),
.Y(n_277)
);

MAJIxp5_ASAP7_75t_L g272 ( 
.A(n_249),
.B(n_13),
.C(n_12),
.Y(n_272)
);

MAJIxp5_ASAP7_75t_L g273 ( 
.A(n_257),
.B(n_11),
.C(n_10),
.Y(n_273)
);

OR2x2_ASAP7_75t_L g285 ( 
.A(n_273),
.B(n_272),
.Y(n_285)
);

INVxp67_ASAP7_75t_SL g274 ( 
.A(n_258),
.Y(n_274)
);

NOR2xp33_ASAP7_75t_L g282 ( 
.A(n_274),
.B(n_254),
.Y(n_282)
);

HB1xp67_ASAP7_75t_L g275 ( 
.A(n_263),
.Y(n_275)
);

XNOR2xp5_ASAP7_75t_L g280 ( 
.A(n_275),
.B(n_255),
.Y(n_280)
);

AOI21xp5_ASAP7_75t_L g278 ( 
.A1(n_268),
.A2(n_269),
.B(n_266),
.Y(n_278)
);

NAND2xp5_ASAP7_75t_L g290 ( 
.A(n_278),
.B(n_282),
.Y(n_290)
);

NAND2xp5_ASAP7_75t_SL g291 ( 
.A(n_280),
.B(n_284),
.Y(n_291)
);

BUFx24_ASAP7_75t_SL g283 ( 
.A(n_274),
.Y(n_283)
);

NAND2xp5_ASAP7_75t_L g294 ( 
.A(n_283),
.B(n_285),
.Y(n_294)
);

HB1xp67_ASAP7_75t_L g286 ( 
.A(n_273),
.Y(n_286)
);

XNOR2xp5_ASAP7_75t_L g292 ( 
.A(n_286),
.B(n_1),
.Y(n_292)
);

OAI21xp5_ASAP7_75t_L g287 ( 
.A1(n_271),
.A2(n_259),
.B(n_9),
.Y(n_287)
);

MAJIxp5_ASAP7_75t_L g295 ( 
.A(n_287),
.B(n_2),
.C(n_3),
.Y(n_295)
);

NOR2xp33_ASAP7_75t_SL g288 ( 
.A(n_277),
.B(n_264),
.Y(n_288)
);

NAND2xp5_ASAP7_75t_SL g298 ( 
.A(n_288),
.B(n_292),
.Y(n_298)
);

NOR2xp33_ASAP7_75t_SL g289 ( 
.A(n_279),
.B(n_1),
.Y(n_289)
);

NAND2xp5_ASAP7_75t_L g301 ( 
.A(n_289),
.B(n_293),
.Y(n_301)
);

AND2x2_ASAP7_75t_L g293 ( 
.A(n_282),
.B(n_2),
.Y(n_293)
);

NOR2xp33_ASAP7_75t_L g296 ( 
.A(n_295),
.B(n_4),
.Y(n_296)
);

NAND2xp5_ASAP7_75t_L g303 ( 
.A(n_296),
.B(n_300),
.Y(n_303)
);

XOR2xp5_ASAP7_75t_L g297 ( 
.A(n_291),
.B(n_281),
.Y(n_297)
);

NOR2xp33_ASAP7_75t_L g302 ( 
.A(n_297),
.B(n_299),
.Y(n_302)
);

INVx6_ASAP7_75t_L g299 ( 
.A(n_288),
.Y(n_299)
);

NOR2xp33_ASAP7_75t_L g300 ( 
.A(n_290),
.B(n_4),
.Y(n_300)
);

AOI21xp5_ASAP7_75t_L g304 ( 
.A1(n_298),
.A2(n_294),
.B(n_5),
.Y(n_304)
);

OAI21xp5_ASAP7_75t_SL g305 ( 
.A1(n_304),
.A2(n_301),
.B(n_298),
.Y(n_305)
);

OAI21xp5_ASAP7_75t_SL g306 ( 
.A1(n_305),
.A2(n_302),
.B(n_303),
.Y(n_306)
);

OAI321xp33_ASAP7_75t_L g307 ( 
.A1(n_306),
.A2(n_4),
.A3(n_6),
.B1(n_7),
.B2(n_8),
.C(n_298),
.Y(n_307)
);

OAI21xp5_ASAP7_75t_L g308 ( 
.A1(n_307),
.A2(n_4),
.B(n_6),
.Y(n_308)
);

AOI22xp5_ASAP7_75t_L g309 ( 
.A1(n_308),
.A2(n_6),
.B1(n_7),
.B2(n_8),
.Y(n_309)
);

AOI21xp5_ASAP7_75t_L g310 ( 
.A1(n_309),
.A2(n_6),
.B(n_7),
.Y(n_310)
);


endmodule