module fake_jpeg_2155_n_303 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_303);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_303;

wire n_159;
wire n_117;
wire n_253;
wire n_286;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_84;
wire n_59;
wire n_98;
wire n_251;
wire n_252;
wire n_273;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_279;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_278;
wire n_205;
wire n_295;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_293;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_281;
wire n_31;
wire n_155;
wire n_207;
wire n_277;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_291;
wire n_236;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_223;
wire n_21;
wire n_57;
wire n_187;
wire n_234;
wire n_288;
wire n_272;
wire n_284;
wire n_280;
wire n_171;
wire n_263;
wire n_23;
wire n_119;
wire n_301;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_289;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_267;
wire n_248;
wire n_30;
wire n_296;
wire n_168;
wire n_298;
wire n_106;
wire n_111;
wire n_197;
wire n_274;
wire n_186;
wire n_44;
wire n_24;
wire n_276;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_269;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_287;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_266;
wire n_34;
wire n_283;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_285;
wire n_215;
wire n_262;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_294;
wire n_300;
wire n_211;
wire n_299;
wire n_230;
wire n_183;
wire n_79;
wire n_170;
wire n_162;
wire n_132;
wire n_133;
wire n_249;
wire n_302;
wire n_67;
wire n_271;
wire n_216;
wire n_217;
wire n_264;
wire n_184;
wire n_53;
wire n_268;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_297;
wire n_226;
wire n_210;
wire n_48;
wire n_35;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_270;
wire n_176;
wire n_199;
wire n_112;
wire n_260;
wire n_265;
wire n_222;
wire n_95;
wire n_275;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_290;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_292;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_258;
wire n_282;
wire n_96;

BUFx6f_ASAP7_75t_L g16 ( 
.A(n_4),
.Y(n_16)
);

BUFx6f_ASAP7_75t_L g17 ( 
.A(n_2),
.Y(n_17)
);

INVx4_ASAP7_75t_L g18 ( 
.A(n_1),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_12),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_11),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_7),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_15),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_1),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_12),
.Y(n_24)
);

INVx4_ASAP7_75t_L g25 ( 
.A(n_11),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_13),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_6),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_1),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_13),
.Y(n_29)
);

INVx11_ASAP7_75t_L g30 ( 
.A(n_3),
.Y(n_30)
);

BUFx3_ASAP7_75t_L g31 ( 
.A(n_3),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_9),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_15),
.Y(n_33)
);

BUFx5_ASAP7_75t_L g34 ( 
.A(n_13),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_4),
.Y(n_35)
);

BUFx16f_ASAP7_75t_L g36 ( 
.A(n_12),
.Y(n_36)
);

INVx1_ASAP7_75t_SL g37 ( 
.A(n_4),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_0),
.Y(n_38)
);

BUFx3_ASAP7_75t_L g39 ( 
.A(n_11),
.Y(n_39)
);

INVx3_ASAP7_75t_L g40 ( 
.A(n_8),
.Y(n_40)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_6),
.Y(n_41)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_7),
.Y(n_42)
);

INVx11_ASAP7_75t_L g43 ( 
.A(n_10),
.Y(n_43)
);

AND2x2_ASAP7_75t_L g44 ( 
.A(n_37),
.B(n_0),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_44),
.B(n_76),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g45 ( 
.A(n_37),
.B(n_14),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_SL g118 ( 
.A(n_45),
.B(n_48),
.Y(n_118)
);

BUFx12f_ASAP7_75t_L g46 ( 
.A(n_36),
.Y(n_46)
);

BUFx10_ASAP7_75t_L g114 ( 
.A(n_46),
.Y(n_114)
);

BUFx3_ASAP7_75t_L g47 ( 
.A(n_36),
.Y(n_47)
);

BUFx3_ASAP7_75t_L g104 ( 
.A(n_47),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_37),
.B(n_14),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_16),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g88 ( 
.A(n_49),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_L g50 ( 
.A(n_21),
.B(n_0),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_L g94 ( 
.A(n_50),
.B(n_68),
.Y(n_94)
);

AOI21xp33_ASAP7_75t_L g51 ( 
.A1(n_19),
.A2(n_2),
.B(n_3),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_SL g131 ( 
.A(n_51),
.B(n_59),
.Y(n_131)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_16),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g105 ( 
.A(n_52),
.Y(n_105)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_19),
.Y(n_53)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_53),
.Y(n_97)
);

BUFx12_ASAP7_75t_L g54 ( 
.A(n_36),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g112 ( 
.A(n_54),
.Y(n_112)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_16),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g113 ( 
.A(n_55),
.Y(n_113)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_18),
.Y(n_56)
);

INVx2_ASAP7_75t_L g101 ( 
.A(n_56),
.Y(n_101)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_20),
.Y(n_57)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_57),
.Y(n_115)
);

INVx3_ASAP7_75t_L g58 ( 
.A(n_18),
.Y(n_58)
);

INVx3_ASAP7_75t_L g107 ( 
.A(n_58),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_21),
.B(n_2),
.Y(n_59)
);

INVx3_ASAP7_75t_L g60 ( 
.A(n_18),
.Y(n_60)
);

BUFx2_ASAP7_75t_L g89 ( 
.A(n_60),
.Y(n_89)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_17),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g135 ( 
.A(n_61),
.Y(n_135)
);

BUFx12_ASAP7_75t_L g62 ( 
.A(n_36),
.Y(n_62)
);

INVx5_ASAP7_75t_L g91 ( 
.A(n_62),
.Y(n_91)
);

BUFx3_ASAP7_75t_L g63 ( 
.A(n_25),
.Y(n_63)
);

INVx5_ASAP7_75t_L g108 ( 
.A(n_63),
.Y(n_108)
);

INVx5_ASAP7_75t_L g64 ( 
.A(n_31),
.Y(n_64)
);

INVx4_ASAP7_75t_L g109 ( 
.A(n_64),
.Y(n_109)
);

INVx8_ASAP7_75t_L g65 ( 
.A(n_17),
.Y(n_65)
);

INVx6_ASAP7_75t_L g90 ( 
.A(n_65),
.Y(n_90)
);

INVx11_ASAP7_75t_L g66 ( 
.A(n_30),
.Y(n_66)
);

INVx2_ASAP7_75t_L g119 ( 
.A(n_66),
.Y(n_119)
);

INVx6_ASAP7_75t_L g67 ( 
.A(n_17),
.Y(n_67)
);

INVx2_ASAP7_75t_L g121 ( 
.A(n_67),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_L g68 ( 
.A(n_23),
.B(n_5),
.Y(n_68)
);

INVx4_ASAP7_75t_SL g69 ( 
.A(n_40),
.Y(n_69)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_69),
.Y(n_116)
);

NAND2xp33_ASAP7_75t_SL g70 ( 
.A(n_25),
.B(n_5),
.Y(n_70)
);

AND2x2_ASAP7_75t_L g132 ( 
.A(n_70),
.B(n_73),
.Y(n_132)
);

BUFx3_ASAP7_75t_L g71 ( 
.A(n_25),
.Y(n_71)
);

INVx2_ASAP7_75t_L g124 ( 
.A(n_71),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_23),
.B(n_5),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_L g103 ( 
.A(n_72),
.B(n_77),
.Y(n_103)
);

INVx8_ASAP7_75t_L g73 ( 
.A(n_35),
.Y(n_73)
);

BUFx6f_ASAP7_75t_L g74 ( 
.A(n_35),
.Y(n_74)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_74),
.Y(n_129)
);

BUFx6f_ASAP7_75t_L g75 ( 
.A(n_35),
.Y(n_75)
);

AND2x2_ASAP7_75t_L g93 ( 
.A(n_75),
.B(n_79),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_SL g76 ( 
.A(n_24),
.B(n_6),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_SL g77 ( 
.A(n_20),
.B(n_7),
.Y(n_77)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_27),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_78),
.B(n_81),
.Y(n_95)
);

BUFx12f_ASAP7_75t_L g79 ( 
.A(n_40),
.Y(n_79)
);

BUFx6f_ASAP7_75t_L g80 ( 
.A(n_22),
.Y(n_80)
);

CKINVDCx20_ASAP7_75t_R g92 ( 
.A(n_80),
.Y(n_92)
);

INVx8_ASAP7_75t_L g81 ( 
.A(n_22),
.Y(n_81)
);

CKINVDCx20_ASAP7_75t_R g82 ( 
.A(n_22),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_82),
.B(n_83),
.Y(n_98)
);

BUFx3_ASAP7_75t_L g83 ( 
.A(n_31),
.Y(n_83)
);

INVx8_ASAP7_75t_L g84 ( 
.A(n_33),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_84),
.B(n_39),
.Y(n_99)
);

BUFx6f_ASAP7_75t_L g85 ( 
.A(n_33),
.Y(n_85)
);

CKINVDCx20_ASAP7_75t_R g111 ( 
.A(n_85),
.Y(n_111)
);

BUFx6f_ASAP7_75t_L g86 ( 
.A(n_33),
.Y(n_86)
);

CKINVDCx20_ASAP7_75t_R g127 ( 
.A(n_86),
.Y(n_127)
);

AOI22xp33_ASAP7_75t_SL g96 ( 
.A1(n_69),
.A2(n_30),
.B1(n_43),
.B2(n_31),
.Y(n_96)
);

AOI22xp33_ASAP7_75t_SL g140 ( 
.A1(n_96),
.A2(n_102),
.B1(n_122),
.B2(n_125),
.Y(n_140)
);

INVxp67_ASAP7_75t_L g155 ( 
.A(n_99),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_59),
.B(n_28),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_L g151 ( 
.A(n_100),
.B(n_106),
.Y(n_151)
);

AOI22xp33_ASAP7_75t_SL g102 ( 
.A1(n_79),
.A2(n_30),
.B1(n_43),
.B2(n_39),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_L g106 ( 
.A(n_72),
.B(n_27),
.Y(n_106)
);

AND2x2_ASAP7_75t_SL g110 ( 
.A(n_44),
.B(n_39),
.Y(n_110)
);

CKINVDCx14_ASAP7_75t_R g167 ( 
.A(n_110),
.Y(n_167)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_45),
.B(n_29),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_L g161 ( 
.A(n_117),
.B(n_120),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_L g120 ( 
.A(n_48),
.B(n_41),
.Y(n_120)
);

AOI22xp33_ASAP7_75t_SL g122 ( 
.A1(n_46),
.A2(n_43),
.B1(n_29),
.B2(n_32),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_L g123 ( 
.A(n_81),
.B(n_28),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_L g169 ( 
.A(n_123),
.B(n_133),
.Y(n_169)
);

AOI22xp33_ASAP7_75t_SL g125 ( 
.A1(n_65),
.A2(n_32),
.B1(n_38),
.B2(n_26),
.Y(n_125)
);

AOI22xp33_ASAP7_75t_SL g126 ( 
.A1(n_73),
.A2(n_26),
.B1(n_38),
.B2(n_24),
.Y(n_126)
);

AOI22xp33_ASAP7_75t_SL g144 ( 
.A1(n_126),
.A2(n_34),
.B1(n_9),
.B2(n_10),
.Y(n_144)
);

AOI22xp5_ASAP7_75t_L g128 ( 
.A1(n_80),
.A2(n_86),
.B1(n_85),
.B2(n_49),
.Y(n_128)
);

OAI22xp5_ASAP7_75t_SL g139 ( 
.A1(n_128),
.A2(n_75),
.B1(n_74),
.B2(n_61),
.Y(n_139)
);

CKINVDCx20_ASAP7_75t_R g130 ( 
.A(n_52),
.Y(n_130)
);

CKINVDCx5p33_ASAP7_75t_R g154 ( 
.A(n_130),
.Y(n_154)
);

NOR2xp33_ASAP7_75t_L g133 ( 
.A(n_84),
.B(n_41),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_L g134 ( 
.A(n_55),
.B(n_42),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_L g141 ( 
.A(n_134),
.B(n_42),
.Y(n_141)
);

AOI22xp5_ASAP7_75t_L g136 ( 
.A1(n_132),
.A2(n_128),
.B1(n_131),
.B2(n_127),
.Y(n_136)
);

OAI22xp5_ASAP7_75t_SL g178 ( 
.A1(n_136),
.A2(n_149),
.B1(n_105),
.B2(n_113),
.Y(n_178)
);

INVx2_ASAP7_75t_L g137 ( 
.A(n_121),
.Y(n_137)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_137),
.Y(n_176)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_97),
.Y(n_138)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_138),
.Y(n_185)
);

AOI22xp5_ASAP7_75t_L g190 ( 
.A1(n_139),
.A2(n_163),
.B1(n_135),
.B2(n_105),
.Y(n_190)
);

OAI21xp33_ASAP7_75t_L g193 ( 
.A1(n_141),
.A2(n_156),
.B(n_174),
.Y(n_193)
);

AOI22xp5_ASAP7_75t_SL g142 ( 
.A1(n_132),
.A2(n_34),
.B1(n_54),
.B2(n_62),
.Y(n_142)
);

INVxp67_ASAP7_75t_L g179 ( 
.A(n_142),
.Y(n_179)
);

BUFx6f_ASAP7_75t_L g143 ( 
.A(n_88),
.Y(n_143)
);

INVx5_ASAP7_75t_L g202 ( 
.A(n_143),
.Y(n_202)
);

INVxp67_ASAP7_75t_L g181 ( 
.A(n_144),
.Y(n_181)
);

INVx2_ASAP7_75t_L g145 ( 
.A(n_121),
.Y(n_145)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_145),
.Y(n_186)
);

INVx2_ASAP7_75t_L g146 ( 
.A(n_129),
.Y(n_146)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_146),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_L g147 ( 
.A(n_110),
.B(n_8),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_L g194 ( 
.A(n_147),
.B(n_170),
.Y(n_194)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_115),
.Y(n_148)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_148),
.Y(n_192)
);

AOI22xp5_ASAP7_75t_L g149 ( 
.A1(n_92),
.A2(n_8),
.B1(n_9),
.B2(n_10),
.Y(n_149)
);

INVx2_ASAP7_75t_L g150 ( 
.A(n_124),
.Y(n_150)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_150),
.Y(n_198)
);

NOR2xp33_ASAP7_75t_L g152 ( 
.A(n_118),
.B(n_87),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_SL g177 ( 
.A(n_152),
.B(n_157),
.Y(n_177)
);

MAJIxp5_ASAP7_75t_L g153 ( 
.A(n_110),
.B(n_94),
.C(n_101),
.Y(n_153)
);

XNOR2xp5_ASAP7_75t_L g188 ( 
.A(n_153),
.B(n_119),
.Y(n_188)
);

AND2x2_ASAP7_75t_L g156 ( 
.A(n_107),
.B(n_101),
.Y(n_156)
);

NOR2xp33_ASAP7_75t_L g157 ( 
.A(n_103),
.B(n_95),
.Y(n_157)
);

INVx4_ASAP7_75t_SL g158 ( 
.A(n_112),
.Y(n_158)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_158),
.Y(n_201)
);

NOR2xp33_ASAP7_75t_L g159 ( 
.A(n_98),
.B(n_116),
.Y(n_159)
);

NOR2xp33_ASAP7_75t_SL g205 ( 
.A(n_159),
.B(n_160),
.Y(n_205)
);

NOR2xp33_ASAP7_75t_L g160 ( 
.A(n_91),
.B(n_107),
.Y(n_160)
);

INVx3_ASAP7_75t_L g162 ( 
.A(n_109),
.Y(n_162)
);

NOR2xp33_ASAP7_75t_L g187 ( 
.A(n_162),
.B(n_164),
.Y(n_187)
);

OAI22xp5_ASAP7_75t_SL g163 ( 
.A1(n_125),
.A2(n_126),
.B1(n_102),
.B2(n_96),
.Y(n_163)
);

NOR2xp33_ASAP7_75t_L g164 ( 
.A(n_91),
.B(n_89),
.Y(n_164)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_89),
.Y(n_165)
);

NOR2xp33_ASAP7_75t_L g189 ( 
.A(n_165),
.B(n_166),
.Y(n_189)
);

NOR2xp33_ASAP7_75t_L g166 ( 
.A(n_112),
.B(n_124),
.Y(n_166)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_109),
.Y(n_168)
);

NOR2xp33_ASAP7_75t_L g197 ( 
.A(n_168),
.B(n_171),
.Y(n_197)
);

OAI32xp33_ASAP7_75t_L g170 ( 
.A1(n_93),
.A2(n_119),
.A3(n_122),
.B1(n_111),
.B2(n_90),
.Y(n_170)
);

INVxp67_ASAP7_75t_L g171 ( 
.A(n_93),
.Y(n_171)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_90),
.Y(n_172)
);

NOR2xp33_ASAP7_75t_L g200 ( 
.A(n_172),
.B(n_173),
.Y(n_200)
);

INVx2_ASAP7_75t_L g173 ( 
.A(n_88),
.Y(n_173)
);

AND2x2_ASAP7_75t_L g174 ( 
.A(n_93),
.B(n_108),
.Y(n_174)
);

INVx3_ASAP7_75t_L g175 ( 
.A(n_108),
.Y(n_175)
);

NOR2xp33_ASAP7_75t_L g204 ( 
.A(n_175),
.B(n_114),
.Y(n_204)
);

AOI22xp5_ASAP7_75t_L g222 ( 
.A1(n_178),
.A2(n_182),
.B1(n_190),
.B2(n_156),
.Y(n_222)
);

CKINVDCx20_ASAP7_75t_R g180 ( 
.A(n_154),
.Y(n_180)
);

INVxp67_ASAP7_75t_SL g213 ( 
.A(n_180),
.Y(n_213)
);

OAI22xp5_ASAP7_75t_SL g182 ( 
.A1(n_136),
.A2(n_167),
.B1(n_140),
.B2(n_155),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_SL g183 ( 
.A(n_161),
.B(n_104),
.Y(n_183)
);

NOR2xp33_ASAP7_75t_SL g220 ( 
.A(n_183),
.B(n_156),
.Y(n_220)
);

CKINVDCx20_ASAP7_75t_R g184 ( 
.A(n_154),
.Y(n_184)
);

NOR2xp33_ASAP7_75t_L g218 ( 
.A(n_184),
.B(n_158),
.Y(n_218)
);

XNOR2xp5_ASAP7_75t_L g208 ( 
.A(n_188),
.B(n_174),
.Y(n_208)
);

NAND2xp5_ASAP7_75t_L g195 ( 
.A(n_153),
.B(n_113),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_L g207 ( 
.A(n_195),
.B(n_196),
.Y(n_207)
);

NAND2xp5_ASAP7_75t_L g196 ( 
.A(n_155),
.B(n_135),
.Y(n_196)
);

AOI21xp5_ASAP7_75t_L g199 ( 
.A1(n_163),
.A2(n_114),
.B(n_104),
.Y(n_199)
);

AOI21xp5_ASAP7_75t_L g225 ( 
.A1(n_199),
.A2(n_175),
.B(n_162),
.Y(n_225)
);

NAND2xp5_ASAP7_75t_L g203 ( 
.A(n_147),
.B(n_114),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_L g217 ( 
.A(n_203),
.B(n_206),
.Y(n_217)
);

INVxp67_ASAP7_75t_L g224 ( 
.A(n_204),
.Y(n_224)
);

NAND2xp5_ASAP7_75t_SL g206 ( 
.A(n_169),
.B(n_151),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_L g246 ( 
.A(n_208),
.B(n_219),
.Y(n_246)
);

AOI22xp33_ASAP7_75t_L g209 ( 
.A1(n_199),
.A2(n_194),
.B1(n_180),
.B2(n_184),
.Y(n_209)
);

INVxp67_ASAP7_75t_L g229 ( 
.A(n_209),
.Y(n_229)
);

OAI22xp5_ASAP7_75t_SL g210 ( 
.A1(n_194),
.A2(n_171),
.B1(n_139),
.B2(n_170),
.Y(n_210)
);

AOI22xp5_ASAP7_75t_L g236 ( 
.A1(n_210),
.A2(n_222),
.B1(n_223),
.B2(n_226),
.Y(n_236)
);

CKINVDCx20_ASAP7_75t_R g211 ( 
.A(n_189),
.Y(n_211)
);

NOR2xp33_ASAP7_75t_L g235 ( 
.A(n_211),
.B(n_220),
.Y(n_235)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_200),
.Y(n_212)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_212),
.Y(n_231)
);

INVx4_ASAP7_75t_L g214 ( 
.A(n_202),
.Y(n_214)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_214),
.Y(n_239)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_191),
.Y(n_215)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_215),
.Y(n_241)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_191),
.Y(n_216)
);

NOR2xp33_ASAP7_75t_L g232 ( 
.A(n_216),
.B(n_221),
.Y(n_232)
);

NOR2xp33_ASAP7_75t_SL g230 ( 
.A(n_218),
.B(n_201),
.Y(n_230)
);

NAND2xp5_ASAP7_75t_L g219 ( 
.A(n_195),
.B(n_174),
.Y(n_219)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_185),
.Y(n_221)
);

OAI22xp5_ASAP7_75t_SL g223 ( 
.A1(n_190),
.A2(n_149),
.B1(n_142),
.B2(n_173),
.Y(n_223)
);

OAI21xp5_ASAP7_75t_SL g245 ( 
.A1(n_225),
.A2(n_201),
.B(n_181),
.Y(n_245)
);

OAI22xp5_ASAP7_75t_SL g226 ( 
.A1(n_182),
.A2(n_137),
.B1(n_145),
.B2(n_143),
.Y(n_226)
);

NOR2xp33_ASAP7_75t_L g227 ( 
.A(n_205),
.B(n_177),
.Y(n_227)
);

INVxp67_ASAP7_75t_L g234 ( 
.A(n_227),
.Y(n_234)
);

INVx2_ASAP7_75t_L g228 ( 
.A(n_176),
.Y(n_228)
);

CKINVDCx20_ASAP7_75t_R g237 ( 
.A(n_228),
.Y(n_237)
);

NAND2xp5_ASAP7_75t_L g248 ( 
.A(n_230),
.B(n_240),
.Y(n_248)
);

AOI221xp5_ASAP7_75t_L g233 ( 
.A1(n_217),
.A2(n_193),
.B1(n_206),
.B2(n_179),
.C(n_203),
.Y(n_233)
);

INVxp67_ASAP7_75t_L g249 ( 
.A(n_233),
.Y(n_249)
);

AOI22xp5_ASAP7_75t_L g238 ( 
.A1(n_210),
.A2(n_222),
.B1(n_226),
.B2(n_223),
.Y(n_238)
);

OAI22xp5_ASAP7_75t_SL g250 ( 
.A1(n_238),
.A2(n_225),
.B1(n_224),
.B2(n_212),
.Y(n_250)
);

NOR2xp33_ASAP7_75t_SL g240 ( 
.A(n_217),
.B(n_177),
.Y(n_240)
);

OAI32xp33_ASAP7_75t_L g242 ( 
.A1(n_207),
.A2(n_179),
.A3(n_196),
.B1(n_187),
.B2(n_197),
.Y(n_242)
);

OAI21xp5_ASAP7_75t_L g252 ( 
.A1(n_242),
.A2(n_245),
.B(n_205),
.Y(n_252)
);

AOI21xp5_ASAP7_75t_SL g243 ( 
.A1(n_213),
.A2(n_181),
.B(n_188),
.Y(n_243)
);

OA21x2_ASAP7_75t_L g260 ( 
.A1(n_243),
.A2(n_186),
.B(n_150),
.Y(n_260)
);

NAND2xp33_ASAP7_75t_L g244 ( 
.A(n_207),
.B(n_178),
.Y(n_244)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_244),
.Y(n_253)
);

MAJIxp5_ASAP7_75t_L g247 ( 
.A(n_246),
.B(n_208),
.C(n_219),
.Y(n_247)
);

XNOR2xp5_ASAP7_75t_L g272 ( 
.A(n_247),
.B(n_254),
.Y(n_272)
);

AOI22xp5_ASAP7_75t_L g268 ( 
.A1(n_250),
.A2(n_236),
.B1(n_238),
.B2(n_230),
.Y(n_268)
);

XNOR2x1_ASAP7_75t_L g251 ( 
.A(n_246),
.B(n_224),
.Y(n_251)
);

XNOR2xp5_ASAP7_75t_SL g266 ( 
.A(n_251),
.B(n_255),
.Y(n_266)
);

AOI22xp33_ASAP7_75t_L g267 ( 
.A1(n_252),
.A2(n_231),
.B1(n_240),
.B2(n_244),
.Y(n_267)
);

MAJIxp5_ASAP7_75t_L g254 ( 
.A(n_243),
.B(n_185),
.C(n_192),
.Y(n_254)
);

XOR2xp5_ASAP7_75t_L g255 ( 
.A(n_242),
.B(n_192),
.Y(n_255)
);

BUFx6f_ASAP7_75t_L g256 ( 
.A(n_231),
.Y(n_256)
);

INVx11_ASAP7_75t_L g263 ( 
.A(n_256),
.Y(n_263)
);

MAJIxp5_ASAP7_75t_L g257 ( 
.A(n_243),
.B(n_216),
.C(n_215),
.Y(n_257)
);

NAND2xp5_ASAP7_75t_SL g265 ( 
.A(n_257),
.B(n_258),
.Y(n_265)
);

A2O1A1Ixp33_ASAP7_75t_L g258 ( 
.A1(n_229),
.A2(n_228),
.B(n_198),
.C(n_176),
.Y(n_258)
);

AOI22xp5_ASAP7_75t_SL g259 ( 
.A1(n_234),
.A2(n_214),
.B1(n_202),
.B2(n_198),
.Y(n_259)
);

NAND2xp5_ASAP7_75t_SL g269 ( 
.A(n_259),
.B(n_245),
.Y(n_269)
);

CKINVDCx16_ASAP7_75t_R g262 ( 
.A(n_260),
.Y(n_262)
);

XNOR2xp5_ASAP7_75t_SL g261 ( 
.A(n_235),
.B(n_186),
.Y(n_261)
);

XNOR2xp5_ASAP7_75t_SL g270 ( 
.A(n_261),
.B(n_232),
.Y(n_270)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_256),
.Y(n_264)
);

NOR2xp33_ASAP7_75t_L g274 ( 
.A(n_264),
.B(n_267),
.Y(n_274)
);

AOI22xp5_ASAP7_75t_L g276 ( 
.A1(n_268),
.A2(n_253),
.B1(n_260),
.B2(n_236),
.Y(n_276)
);

CKINVDCx16_ASAP7_75t_R g278 ( 
.A(n_269),
.Y(n_278)
);

XNOR2xp5_ASAP7_75t_SL g273 ( 
.A(n_270),
.B(n_261),
.Y(n_273)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_248),
.Y(n_271)
);

NOR2xp33_ASAP7_75t_L g275 ( 
.A(n_271),
.B(n_255),
.Y(n_275)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_273),
.Y(n_285)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_275),
.Y(n_286)
);

AOI22xp5_ASAP7_75t_L g282 ( 
.A1(n_276),
.A2(n_262),
.B1(n_268),
.B2(n_258),
.Y(n_282)
);

NOR2xp33_ASAP7_75t_L g277 ( 
.A(n_272),
.B(n_247),
.Y(n_277)
);

NOR2xp33_ASAP7_75t_SL g284 ( 
.A(n_277),
.B(n_279),
.Y(n_284)
);

XOR2xp5_ASAP7_75t_L g279 ( 
.A(n_272),
.B(n_251),
.Y(n_279)
);

OAI21xp5_ASAP7_75t_SL g280 ( 
.A1(n_265),
.A2(n_260),
.B(n_249),
.Y(n_280)
);

AOI21xp5_ASAP7_75t_L g288 ( 
.A1(n_280),
.A2(n_281),
.B(n_266),
.Y(n_288)
);

OAI322xp33_ASAP7_75t_L g281 ( 
.A1(n_270),
.A2(n_249),
.A3(n_232),
.B1(n_254),
.B2(n_257),
.C1(n_237),
.C2(n_241),
.Y(n_281)
);

XOR2xp5_ASAP7_75t_L g293 ( 
.A(n_282),
.B(n_239),
.Y(n_293)
);

A2O1A1O1Ixp25_ASAP7_75t_L g283 ( 
.A1(n_274),
.A2(n_266),
.B(n_237),
.C(n_241),
.D(n_264),
.Y(n_283)
);

NAND2xp5_ASAP7_75t_L g290 ( 
.A(n_283),
.B(n_287),
.Y(n_290)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_280),
.Y(n_287)
);

OAI221xp5_ASAP7_75t_L g289 ( 
.A1(n_288),
.A2(n_273),
.B1(n_279),
.B2(n_276),
.C(n_278),
.Y(n_289)
);

NAND2xp5_ASAP7_75t_SL g297 ( 
.A(n_289),
.B(n_293),
.Y(n_297)
);

NAND2xp5_ASAP7_75t_L g291 ( 
.A(n_286),
.B(n_278),
.Y(n_291)
);

NAND2xp5_ASAP7_75t_L g296 ( 
.A(n_291),
.B(n_292),
.Y(n_296)
);

NOR2xp33_ASAP7_75t_L g292 ( 
.A(n_284),
.B(n_239),
.Y(n_292)
);

MAJIxp5_ASAP7_75t_L g294 ( 
.A(n_290),
.B(n_285),
.C(n_282),
.Y(n_294)
);

NOR2xp33_ASAP7_75t_L g299 ( 
.A(n_294),
.B(n_295),
.Y(n_299)
);

OAI21xp5_ASAP7_75t_SL g295 ( 
.A1(n_293),
.A2(n_283),
.B(n_263),
.Y(n_295)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_296),
.Y(n_298)
);

NAND2xp5_ASAP7_75t_L g301 ( 
.A(n_298),
.B(n_300),
.Y(n_301)
);

AOI21x1_ASAP7_75t_L g300 ( 
.A1(n_297),
.A2(n_263),
.B(n_146),
.Y(n_300)
);

BUFx24_ASAP7_75t_SL g302 ( 
.A(n_299),
.Y(n_302)
);

XOR2xp5_ASAP7_75t_L g303 ( 
.A(n_302),
.B(n_301),
.Y(n_303)
);


endmodule