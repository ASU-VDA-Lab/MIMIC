module fake_jpeg_121_n_675 (n_13, n_1, n_10, n_6, n_14, n_19, n_18, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_675);

input n_13;
input n_1;
input n_10;
input n_6;
input n_14;
input n_19;
input n_18;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_675;

wire n_529;
wire n_595;
wire n_390;
wire n_552;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_252;
wire n_182;
wire n_525;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_586;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_657;
wire n_27;
wire n_664;
wire n_365;
wire n_179;
wire n_620;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_611;
wire n_44;
wire n_519;
wire n_355;
wire n_276;
wire n_143;
wire n_431;
wire n_102;
wire n_549;
wire n_196;
wire n_66;
wire n_374;
wire n_566;
wire n_142;
wire n_417;
wire n_362;
wire n_470;
wire n_597;
wire n_172;
wire n_547;
wire n_345;
wire n_591;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_513;
wire n_283;
wire n_107;
wire n_490;
wire n_635;
wire n_517;
wire n_629;
wire n_415;
wire n_479;
wire n_543;
wire n_357;
wire n_89;
wire n_131;
wire n_607;
wire n_294;
wire n_230;
wire n_643;
wire n_170;
wire n_602;
wire n_313;
wire n_542;
wire n_574;
wire n_264;
wire n_647;
wire n_437;
wire n_93;
wire n_227;
wire n_559;
wire n_641;
wire n_48;
wire n_465;
wire n_638;
wire n_200;
wire n_582;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_623;
wire n_579;
wire n_416;
wire n_221;
wire n_256;
wire n_454;
wire n_540;
wire n_292;
wire n_213;
wire n_135;
wire n_435;
wire n_189;
wire n_637;
wire n_370;
wire n_410;
wire n_571;
wire n_82;
wire n_155;
wire n_508;
wire n_672;
wire n_309;
wire n_624;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_606;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_569;
wire n_596;
wire n_400;
wire n_646;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_544;
wire n_31;
wire n_277;
wire n_663;
wire n_255;
wire n_605;
wire n_601;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_530;
wire n_634;
wire n_23;
wire n_69;
wire n_658;
wire n_195;
wire n_450;
wire n_557;
wire n_408;
wire n_80;
wire n_562;
wire n_204;
wire n_666;
wire n_639;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_645;
wire n_298;
wire n_106;
wire n_545;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_584;
wire n_254;
wire n_608;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_622;
wire n_463;
wire n_667;
wire n_92;
wire n_332;
wire n_640;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_653;
wire n_474;
wire n_539;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_626;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_668;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_575;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_511;
wire n_305;
wire n_161;
wire n_441;
wire n_555;
wire n_342;
wire n_642;
wire n_101;
wire n_226;
wire n_509;
wire n_644;
wire n_149;
wire n_87;
wire n_46;
wire n_578;
wire n_656;
wire n_589;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_614;
wire n_97;
wire n_649;
wire n_573;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_610;
wire n_174;
wire n_198;
wire n_422;
wire n_560;
wire n_190;
wire n_510;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_536;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_537;
wire n_110;
wire n_594;
wire n_590;
wire n_531;
wire n_76;
wire n_278;
wire n_343;
wire n_577;
wire n_26;
wire n_88;
wire n_397;
wire n_592;
wire n_363;
wire n_570;
wire n_238;
wire n_598;
wire n_615;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_488;
wire n_662;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_554;
wire n_301;
wire n_609;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_648;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_523;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_533;
wire n_612;
wire n_296;
wire n_384;
wire n_588;
wire n_168;
wire n_670;
wire n_459;
wire n_274;
wire n_485;
wire n_585;
wire n_491;
wire n_24;
wire n_526;
wire n_467;
wire n_269;
wire n_572;
wire n_546;
wire n_287;
wire n_219;
wire n_452;
wire n_631;
wire n_433;
wire n_636;
wire n_77;
wire n_473;
wire n_45;
wire n_520;
wire n_476;
wire n_337;
wire n_317;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_344;
wire n_328;
wire n_650;
wire n_218;
wire n_63;
wire n_652;
wire n_599;
wire n_239;
wire n_674;
wire n_243;
wire n_481;
wire n_628;
wire n_619;
wire n_348;
wire n_587;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_583;
wire n_522;
wire n_333;
wire n_518;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_565;
wire n_302;
wire n_216;
wire n_528;
wire n_184;
wire n_655;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_199;
wire n_260;
wire n_550;
wire n_413;
wire n_275;
wire n_494;
wire n_604;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_551;
wire n_36;
wire n_62;
wire n_600;
wire n_492;
wire n_603;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_567;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_515;
wire n_347;
wire n_521;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_538;
wire n_625;
wire n_147;
wire n_449;
wire n_627;
wire n_98;
wire n_251;
wire n_534;
wire n_472;
wire n_279;
wire n_593;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_618;
wire n_356;
wire n_119;
wire n_484;
wire n_568;
wire n_83;
wire n_395;
wire n_659;
wire n_125;
wire n_661;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_576;
wire n_469;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_553;
wire n_257;
wire n_61;
wire n_173;
wire n_561;
wire n_244;
wire n_232;
wire n_527;
wire n_482;
wire n_673;
wire n_58;
wire n_41;
wire n_613;
wire n_630;
wire n_266;
wire n_548;
wire n_665;
wire n_72;
wire n_512;
wire n_654;
wire n_445;
wire n_443;
wire n_617;
wire n_215;
wire n_212;
wire n_516;
wire n_183;
wire n_409;
wire n_532;
wire n_249;
wire n_412;
wire n_581;
wire n_217;
wire n_471;
wire n_580;
wire n_541;
wire n_53;
wire n_372;
wire n_558;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_535;
wire n_671;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_556;
wire n_669;
wire n_524;
wire n_402;
wire n_563;
wire n_504;
wire n_438;
wire n_475;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_660;
wire n_373;
wire n_633;
wire n_112;
wire n_632;
wire n_616;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_514;
wire n_651;
wire n_564;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_621;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_16),
.Y(n_20)
);

INVx4_ASAP7_75t_L g21 ( 
.A(n_19),
.Y(n_21)
);

INVx3_ASAP7_75t_L g22 ( 
.A(n_8),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_17),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_9),
.Y(n_24)
);

INVx11_ASAP7_75t_L g25 ( 
.A(n_9),
.Y(n_25)
);

INVx3_ASAP7_75t_L g26 ( 
.A(n_1),
.Y(n_26)
);

BUFx5_ASAP7_75t_L g27 ( 
.A(n_17),
.Y(n_27)
);

BUFx5_ASAP7_75t_L g28 ( 
.A(n_15),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_4),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_10),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_12),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_13),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_10),
.Y(n_33)
);

BUFx5_ASAP7_75t_L g34 ( 
.A(n_1),
.Y(n_34)
);

INVx2_ASAP7_75t_L g35 ( 
.A(n_15),
.Y(n_35)
);

BUFx24_ASAP7_75t_L g36 ( 
.A(n_19),
.Y(n_36)
);

INVx2_ASAP7_75t_L g37 ( 
.A(n_1),
.Y(n_37)
);

INVxp67_ASAP7_75t_L g38 ( 
.A(n_16),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_2),
.Y(n_39)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_6),
.Y(n_40)
);

INVx4_ASAP7_75t_L g41 ( 
.A(n_15),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_2),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_2),
.Y(n_43)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_12),
.Y(n_44)
);

INVx4_ASAP7_75t_L g45 ( 
.A(n_10),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_13),
.Y(n_46)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_12),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_11),
.Y(n_48)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_7),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_1),
.Y(n_50)
);

BUFx12f_ASAP7_75t_L g51 ( 
.A(n_3),
.Y(n_51)
);

INVx3_ASAP7_75t_L g52 ( 
.A(n_8),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_7),
.Y(n_53)
);

BUFx3_ASAP7_75t_L g54 ( 
.A(n_15),
.Y(n_54)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_17),
.Y(n_55)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_3),
.Y(n_56)
);

INVx1_ASAP7_75t_SL g57 ( 
.A(n_12),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_18),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_38),
.B(n_49),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_L g134 ( 
.A(n_59),
.B(n_75),
.Y(n_134)
);

CKINVDCx20_ASAP7_75t_R g60 ( 
.A(n_24),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g133 ( 
.A(n_60),
.B(n_66),
.Y(n_133)
);

BUFx4f_ASAP7_75t_SL g61 ( 
.A(n_51),
.Y(n_61)
);

BUFx8_ASAP7_75t_L g167 ( 
.A(n_61),
.Y(n_167)
);

BUFx3_ASAP7_75t_L g62 ( 
.A(n_54),
.Y(n_62)
);

BUFx3_ASAP7_75t_L g170 ( 
.A(n_62),
.Y(n_170)
);

INVx2_ASAP7_75t_L g63 ( 
.A(n_37),
.Y(n_63)
);

INVx2_ASAP7_75t_L g137 ( 
.A(n_63),
.Y(n_137)
);

INVx3_ASAP7_75t_L g64 ( 
.A(n_21),
.Y(n_64)
);

INVx2_ASAP7_75t_SL g188 ( 
.A(n_64),
.Y(n_188)
);

INVx6_ASAP7_75t_L g65 ( 
.A(n_24),
.Y(n_65)
);

BUFx6f_ASAP7_75t_L g136 ( 
.A(n_65),
.Y(n_136)
);

CKINVDCx20_ASAP7_75t_R g66 ( 
.A(n_24),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_24),
.Y(n_67)
);

BUFx6f_ASAP7_75t_L g154 ( 
.A(n_67),
.Y(n_154)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_30),
.Y(n_68)
);

BUFx6f_ASAP7_75t_L g189 ( 
.A(n_68),
.Y(n_189)
);

INVx4_ASAP7_75t_L g69 ( 
.A(n_34),
.Y(n_69)
);

INVx3_ASAP7_75t_L g153 ( 
.A(n_69),
.Y(n_153)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_31),
.Y(n_70)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_70),
.Y(n_141)
);

INVx13_ASAP7_75t_L g71 ( 
.A(n_36),
.Y(n_71)
);

INVx5_ASAP7_75t_SL g217 ( 
.A(n_71),
.Y(n_217)
);

INVx3_ASAP7_75t_L g72 ( 
.A(n_21),
.Y(n_72)
);

INVx3_ASAP7_75t_L g190 ( 
.A(n_72),
.Y(n_190)
);

AND2x2_ASAP7_75t_L g73 ( 
.A(n_37),
.B(n_26),
.Y(n_73)
);

AND2x2_ASAP7_75t_SL g160 ( 
.A(n_73),
.B(n_92),
.Y(n_160)
);

INVx3_ASAP7_75t_L g74 ( 
.A(n_21),
.Y(n_74)
);

INVx3_ASAP7_75t_L g195 ( 
.A(n_74),
.Y(n_195)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_31),
.B(n_9),
.Y(n_75)
);

BUFx6f_ASAP7_75t_L g76 ( 
.A(n_30),
.Y(n_76)
);

BUFx6f_ASAP7_75t_L g199 ( 
.A(n_76),
.Y(n_199)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_40),
.Y(n_77)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_77),
.Y(n_159)
);

BUFx6f_ASAP7_75t_L g78 ( 
.A(n_30),
.Y(n_78)
);

BUFx6f_ASAP7_75t_L g222 ( 
.A(n_78),
.Y(n_222)
);

INVx2_ASAP7_75t_R g79 ( 
.A(n_41),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_SL g177 ( 
.A(n_79),
.B(n_23),
.Y(n_177)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_40),
.B(n_9),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_L g147 ( 
.A(n_80),
.B(n_88),
.Y(n_147)
);

CKINVDCx20_ASAP7_75t_R g81 ( 
.A(n_58),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g142 ( 
.A(n_81),
.B(n_84),
.Y(n_142)
);

INVx2_ASAP7_75t_L g82 ( 
.A(n_35),
.Y(n_82)
);

INVx2_ASAP7_75t_L g152 ( 
.A(n_82),
.Y(n_152)
);

BUFx6f_ASAP7_75t_L g83 ( 
.A(n_30),
.Y(n_83)
);

INVx6_ASAP7_75t_L g135 ( 
.A(n_83),
.Y(n_135)
);

CKINVDCx20_ASAP7_75t_R g84 ( 
.A(n_58),
.Y(n_84)
);

CKINVDCx20_ASAP7_75t_R g85 ( 
.A(n_58),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g157 ( 
.A(n_85),
.B(n_86),
.Y(n_157)
);

CKINVDCx20_ASAP7_75t_R g86 ( 
.A(n_58),
.Y(n_86)
);

INVx2_ASAP7_75t_L g87 ( 
.A(n_35),
.Y(n_87)
);

INVx2_ASAP7_75t_L g156 ( 
.A(n_87),
.Y(n_156)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_44),
.B(n_8),
.Y(n_88)
);

BUFx6f_ASAP7_75t_L g89 ( 
.A(n_48),
.Y(n_89)
);

INVx6_ASAP7_75t_L g211 ( 
.A(n_89),
.Y(n_211)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_44),
.Y(n_90)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_90),
.Y(n_193)
);

INVx3_ASAP7_75t_L g91 ( 
.A(n_41),
.Y(n_91)
);

INVx3_ASAP7_75t_L g201 ( 
.A(n_91),
.Y(n_201)
);

AND2x2_ASAP7_75t_L g92 ( 
.A(n_26),
.B(n_0),
.Y(n_92)
);

BUFx8_ASAP7_75t_L g93 ( 
.A(n_36),
.Y(n_93)
);

BUFx12f_ASAP7_75t_L g176 ( 
.A(n_93),
.Y(n_176)
);

AND2x2_ASAP7_75t_L g94 ( 
.A(n_26),
.B(n_0),
.Y(n_94)
);

AND2x2_ASAP7_75t_SL g164 ( 
.A(n_94),
.B(n_25),
.Y(n_164)
);

INVx6_ASAP7_75t_L g95 ( 
.A(n_48),
.Y(n_95)
);

INVx3_ASAP7_75t_SL g215 ( 
.A(n_95),
.Y(n_215)
);

BUFx12_ASAP7_75t_L g96 ( 
.A(n_36),
.Y(n_96)
);

INVx5_ASAP7_75t_L g191 ( 
.A(n_96),
.Y(n_191)
);

BUFx6f_ASAP7_75t_L g97 ( 
.A(n_48),
.Y(n_97)
);

INVx8_ASAP7_75t_L g204 ( 
.A(n_97),
.Y(n_204)
);

BUFx5_ASAP7_75t_L g98 ( 
.A(n_36),
.Y(n_98)
);

INVx4_ASAP7_75t_L g144 ( 
.A(n_98),
.Y(n_144)
);

BUFx6f_ASAP7_75t_L g99 ( 
.A(n_53),
.Y(n_99)
);

INVx5_ASAP7_75t_L g198 ( 
.A(n_99),
.Y(n_198)
);

CKINVDCx20_ASAP7_75t_R g100 ( 
.A(n_53),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g161 ( 
.A(n_100),
.B(n_113),
.Y(n_161)
);

BUFx6f_ASAP7_75t_L g101 ( 
.A(n_53),
.Y(n_101)
);

INVx5_ASAP7_75t_L g208 ( 
.A(n_101),
.Y(n_208)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_47),
.Y(n_102)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_102),
.Y(n_202)
);

INVx3_ASAP7_75t_L g103 ( 
.A(n_41),
.Y(n_103)
);

INVx3_ASAP7_75t_L g213 ( 
.A(n_103),
.Y(n_213)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_47),
.Y(n_104)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_104),
.Y(n_214)
);

BUFx5_ASAP7_75t_L g105 ( 
.A(n_36),
.Y(n_105)
);

INVx4_ASAP7_75t_L g145 ( 
.A(n_105),
.Y(n_145)
);

BUFx3_ASAP7_75t_L g106 ( 
.A(n_54),
.Y(n_106)
);

INVx5_ASAP7_75t_L g224 ( 
.A(n_106),
.Y(n_224)
);

INVx2_ASAP7_75t_L g107 ( 
.A(n_51),
.Y(n_107)
);

INVx2_ASAP7_75t_L g158 ( 
.A(n_107),
.Y(n_158)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_49),
.Y(n_108)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_108),
.Y(n_220)
);

INVx1_ASAP7_75t_SL g109 ( 
.A(n_51),
.Y(n_109)
);

INVx3_ASAP7_75t_L g223 ( 
.A(n_109),
.Y(n_223)
);

INVx2_ASAP7_75t_L g110 ( 
.A(n_51),
.Y(n_110)
);

INVx2_ASAP7_75t_L g169 ( 
.A(n_110),
.Y(n_169)
);

INVx2_ASAP7_75t_L g111 ( 
.A(n_51),
.Y(n_111)
);

INVx2_ASAP7_75t_L g178 ( 
.A(n_111),
.Y(n_178)
);

INVx11_ASAP7_75t_L g112 ( 
.A(n_34),
.Y(n_112)
);

INVx4_ASAP7_75t_L g173 ( 
.A(n_112),
.Y(n_173)
);

CKINVDCx20_ASAP7_75t_R g113 ( 
.A(n_39),
.Y(n_113)
);

BUFx6f_ASAP7_75t_L g114 ( 
.A(n_39),
.Y(n_114)
);

INVx3_ASAP7_75t_L g228 ( 
.A(n_114),
.Y(n_228)
);

CKINVDCx20_ASAP7_75t_R g115 ( 
.A(n_39),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_L g162 ( 
.A(n_115),
.B(n_120),
.Y(n_162)
);

BUFx5_ASAP7_75t_L g116 ( 
.A(n_27),
.Y(n_116)
);

INVx4_ASAP7_75t_L g187 ( 
.A(n_116),
.Y(n_187)
);

INVx6_ASAP7_75t_L g117 ( 
.A(n_39),
.Y(n_117)
);

INVx2_ASAP7_75t_L g179 ( 
.A(n_117),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_L g118 ( 
.A(n_22),
.B(n_0),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_L g168 ( 
.A(n_118),
.B(n_122),
.Y(n_168)
);

BUFx3_ASAP7_75t_L g119 ( 
.A(n_54),
.Y(n_119)
);

INVx4_ASAP7_75t_L g194 ( 
.A(n_119),
.Y(n_194)
);

CKINVDCx20_ASAP7_75t_R g120 ( 
.A(n_42),
.Y(n_120)
);

INVx11_ASAP7_75t_L g121 ( 
.A(n_34),
.Y(n_121)
);

INVx4_ASAP7_75t_L g200 ( 
.A(n_121),
.Y(n_200)
);

NAND2xp5_ASAP7_75t_L g122 ( 
.A(n_22),
.B(n_0),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_L g123 ( 
.A(n_22),
.B(n_0),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_L g174 ( 
.A(n_123),
.B(n_125),
.Y(n_174)
);

INVx13_ASAP7_75t_L g124 ( 
.A(n_57),
.Y(n_124)
);

INVx3_ASAP7_75t_L g230 ( 
.A(n_124),
.Y(n_230)
);

NOR2xp33_ASAP7_75t_L g125 ( 
.A(n_55),
.B(n_10),
.Y(n_125)
);

BUFx12f_ASAP7_75t_L g126 ( 
.A(n_52),
.Y(n_126)
);

HB1xp67_ASAP7_75t_L g151 ( 
.A(n_126),
.Y(n_151)
);

BUFx6f_ASAP7_75t_L g127 ( 
.A(n_42),
.Y(n_127)
);

INVx2_ASAP7_75t_L g182 ( 
.A(n_127),
.Y(n_182)
);

INVx8_ASAP7_75t_L g128 ( 
.A(n_42),
.Y(n_128)
);

INVx2_ASAP7_75t_L g184 ( 
.A(n_128),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_L g129 ( 
.A(n_52),
.B(n_1),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_L g185 ( 
.A(n_129),
.B(n_2),
.Y(n_185)
);

INVx13_ASAP7_75t_L g130 ( 
.A(n_57),
.Y(n_130)
);

HB1xp67_ASAP7_75t_L g172 ( 
.A(n_130),
.Y(n_172)
);

BUFx12_ASAP7_75t_L g131 ( 
.A(n_27),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_L g163 ( 
.A(n_131),
.B(n_61),
.Y(n_163)
);

BUFx3_ASAP7_75t_L g132 ( 
.A(n_45),
.Y(n_132)
);

INVx2_ASAP7_75t_L g186 ( 
.A(n_132),
.Y(n_186)
);

AOI22xp33_ASAP7_75t_L g138 ( 
.A1(n_118),
.A2(n_122),
.B1(n_129),
.B2(n_123),
.Y(n_138)
);

OAI22xp5_ASAP7_75t_L g252 ( 
.A1(n_138),
.A2(n_140),
.B1(n_146),
.B2(n_148),
.Y(n_252)
);

OAI22xp33_ASAP7_75t_SL g139 ( 
.A1(n_127),
.A2(n_52),
.B1(n_45),
.B2(n_50),
.Y(n_139)
);

AOI22xp5_ASAP7_75t_L g268 ( 
.A1(n_139),
.A2(n_181),
.B1(n_231),
.B2(n_5),
.Y(n_268)
);

AOI22xp5_ASAP7_75t_L g140 ( 
.A1(n_73),
.A2(n_45),
.B1(n_55),
.B2(n_46),
.Y(n_140)
);

CKINVDCx20_ASAP7_75t_R g143 ( 
.A(n_73),
.Y(n_143)
);

NOR2xp33_ASAP7_75t_SL g267 ( 
.A(n_143),
.B(n_171),
.Y(n_267)
);

AOI22xp33_ASAP7_75t_L g146 ( 
.A1(n_89),
.A2(n_57),
.B1(n_50),
.B2(n_43),
.Y(n_146)
);

AOI22xp33_ASAP7_75t_L g148 ( 
.A1(n_97),
.A2(n_43),
.B1(n_29),
.B2(n_56),
.Y(n_148)
);

AOI22xp5_ASAP7_75t_L g149 ( 
.A1(n_92),
.A2(n_20),
.B1(n_46),
.B2(n_33),
.Y(n_149)
);

OAI22xp5_ASAP7_75t_L g261 ( 
.A1(n_149),
.A2(n_150),
.B1(n_155),
.B2(n_165),
.Y(n_261)
);

AOI22xp33_ASAP7_75t_SL g150 ( 
.A1(n_93),
.A2(n_109),
.B1(n_25),
.B2(n_121),
.Y(n_150)
);

AOI22xp33_ASAP7_75t_SL g155 ( 
.A1(n_93),
.A2(n_25),
.B1(n_29),
.B2(n_56),
.Y(n_155)
);

CKINVDCx16_ASAP7_75t_R g246 ( 
.A(n_163),
.Y(n_246)
);

AND2x2_ASAP7_75t_L g235 ( 
.A(n_164),
.B(n_119),
.Y(n_235)
);

AOI22xp33_ASAP7_75t_SL g165 ( 
.A1(n_112),
.A2(n_33),
.B1(n_32),
.B2(n_23),
.Y(n_165)
);

AOI22xp5_ASAP7_75t_SL g166 ( 
.A1(n_92),
.A2(n_94),
.B1(n_72),
.B2(n_74),
.Y(n_166)
);

OR2x2_ASAP7_75t_L g304 ( 
.A(n_166),
.B(n_177),
.Y(n_304)
);

NOR2xp33_ASAP7_75t_L g171 ( 
.A(n_70),
.B(n_32),
.Y(n_171)
);

NOR2xp33_ASAP7_75t_L g175 ( 
.A(n_77),
.B(n_20),
.Y(n_175)
);

NOR2xp33_ASAP7_75t_SL g277 ( 
.A(n_175),
.B(n_180),
.Y(n_277)
);

NOR2xp33_ASAP7_75t_L g180 ( 
.A(n_90),
.B(n_13),
.Y(n_180)
);

OAI22xp33_ASAP7_75t_SL g181 ( 
.A1(n_99),
.A2(n_28),
.B1(n_27),
.B2(n_4),
.Y(n_181)
);

CKINVDCx20_ASAP7_75t_R g183 ( 
.A(n_117),
.Y(n_183)
);

NOR2xp33_ASAP7_75t_L g255 ( 
.A(n_183),
.B(n_210),
.Y(n_255)
);

NAND2xp5_ASAP7_75t_SL g247 ( 
.A(n_185),
.B(n_196),
.Y(n_247)
);

AOI22xp33_ASAP7_75t_L g192 ( 
.A1(n_101),
.A2(n_2),
.B1(n_3),
.B2(n_4),
.Y(n_192)
);

OAI22xp5_ASAP7_75t_L g283 ( 
.A1(n_192),
.A2(n_205),
.B1(n_206),
.B2(n_219),
.Y(n_283)
);

NAND2xp5_ASAP7_75t_SL g196 ( 
.A(n_102),
.B(n_13),
.Y(n_196)
);

INVx2_ASAP7_75t_L g197 ( 
.A(n_63),
.Y(n_197)
);

INVx2_ASAP7_75t_L g233 ( 
.A(n_197),
.Y(n_233)
);

NAND2xp5_ASAP7_75t_L g203 ( 
.A(n_104),
.B(n_11),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_SL g260 ( 
.A(n_203),
.B(n_207),
.Y(n_260)
);

AOI22xp33_ASAP7_75t_L g205 ( 
.A1(n_114),
.A2(n_87),
.B1(n_82),
.B2(n_78),
.Y(n_205)
);

AOI22xp33_ASAP7_75t_L g206 ( 
.A1(n_67),
.A2(n_3),
.B1(n_4),
.B2(n_5),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_L g207 ( 
.A(n_108),
.B(n_11),
.Y(n_207)
);

INVx2_ASAP7_75t_L g209 ( 
.A(n_107),
.Y(n_209)
);

INVx2_ASAP7_75t_L g240 ( 
.A(n_209),
.Y(n_240)
);

NOR2xp33_ASAP7_75t_L g210 ( 
.A(n_61),
.B(n_126),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_L g212 ( 
.A(n_94),
.B(n_11),
.Y(n_212)
);

OR2x2_ASAP7_75t_L g312 ( 
.A(n_212),
.B(n_218),
.Y(n_312)
);

INVx2_ASAP7_75t_L g216 ( 
.A(n_110),
.Y(n_216)
);

INVx2_ASAP7_75t_L g243 ( 
.A(n_216),
.Y(n_243)
);

AOI22xp5_ASAP7_75t_SL g218 ( 
.A1(n_64),
.A2(n_28),
.B1(n_14),
.B2(n_16),
.Y(n_218)
);

OAI22xp5_ASAP7_75t_L g219 ( 
.A1(n_95),
.A2(n_65),
.B1(n_76),
.B2(n_68),
.Y(n_219)
);

AOI22xp33_ASAP7_75t_SL g221 ( 
.A1(n_69),
.A2(n_28),
.B1(n_14),
.B2(n_16),
.Y(n_221)
);

AOI22xp33_ASAP7_75t_SL g239 ( 
.A1(n_221),
.A2(n_105),
.B1(n_98),
.B2(n_106),
.Y(n_239)
);

NAND2xp5_ASAP7_75t_L g225 ( 
.A(n_111),
.B(n_8),
.Y(n_225)
);

NAND2xp5_ASAP7_75t_L g253 ( 
.A(n_225),
.B(n_4),
.Y(n_253)
);

INVx2_ASAP7_75t_L g226 ( 
.A(n_91),
.Y(n_226)
);

INVx2_ASAP7_75t_L g269 ( 
.A(n_226),
.Y(n_269)
);

NOR2xp33_ASAP7_75t_L g227 ( 
.A(n_126),
.B(n_19),
.Y(n_227)
);

NOR2xp33_ASAP7_75t_L g262 ( 
.A(n_227),
.B(n_6),
.Y(n_262)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_103),
.Y(n_229)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_229),
.Y(n_241)
);

OAI22xp5_ASAP7_75t_SL g231 ( 
.A1(n_83),
.A2(n_7),
.B1(n_18),
.B2(n_17),
.Y(n_231)
);

HB1xp67_ASAP7_75t_L g232 ( 
.A(n_188),
.Y(n_232)
);

BUFx2_ASAP7_75t_L g356 ( 
.A(n_232),
.Y(n_356)
);

OR2x4_ASAP7_75t_L g234 ( 
.A(n_160),
.B(n_79),
.Y(n_234)
);

OR2x2_ASAP7_75t_L g320 ( 
.A(n_234),
.B(n_282),
.Y(n_320)
);

AND2x2_ASAP7_75t_L g357 ( 
.A(n_235),
.B(n_280),
.Y(n_357)
);

A2O1A1Ixp33_ASAP7_75t_L g236 ( 
.A1(n_174),
.A2(n_124),
.B(n_130),
.C(n_71),
.Y(n_236)
);

AOI21xp33_ASAP7_75t_L g324 ( 
.A1(n_236),
.A2(n_307),
.B(n_208),
.Y(n_324)
);

INVx13_ASAP7_75t_L g237 ( 
.A(n_167),
.Y(n_237)
);

CKINVDCx16_ASAP7_75t_R g328 ( 
.A(n_237),
.Y(n_328)
);

AND2x2_ASAP7_75t_L g238 ( 
.A(n_160),
.B(n_132),
.Y(n_238)
);

NAND2xp33_ASAP7_75t_SL g370 ( 
.A(n_238),
.B(n_248),
.Y(n_370)
);

INVxp67_ASAP7_75t_L g332 ( 
.A(n_239),
.Y(n_332)
);

INVx5_ASAP7_75t_L g242 ( 
.A(n_167),
.Y(n_242)
);

INVx4_ASAP7_75t_L g336 ( 
.A(n_242),
.Y(n_336)
);

AOI22xp33_ASAP7_75t_SL g244 ( 
.A1(n_230),
.A2(n_62),
.B1(n_128),
.B2(n_96),
.Y(n_244)
);

INVxp67_ASAP7_75t_L g369 ( 
.A(n_244),
.Y(n_369)
);

BUFx12f_ASAP7_75t_L g245 ( 
.A(n_167),
.Y(n_245)
);

INVx8_ASAP7_75t_L g338 ( 
.A(n_245),
.Y(n_338)
);

AND2x2_ASAP7_75t_L g248 ( 
.A(n_160),
.B(n_3),
.Y(n_248)
);

BUFx6f_ASAP7_75t_L g249 ( 
.A(n_154),
.Y(n_249)
);

INVx6_ASAP7_75t_L g327 ( 
.A(n_249),
.Y(n_327)
);

CKINVDCx20_ASAP7_75t_R g250 ( 
.A(n_162),
.Y(n_250)
);

NAND2xp5_ASAP7_75t_SL g360 ( 
.A(n_250),
.B(n_253),
.Y(n_360)
);

AOI21xp5_ASAP7_75t_L g251 ( 
.A1(n_181),
.A2(n_96),
.B(n_116),
.Y(n_251)
);

AOI21xp5_ASAP7_75t_L g361 ( 
.A1(n_251),
.A2(n_281),
.B(n_236),
.Y(n_361)
);

MAJIxp5_ASAP7_75t_L g254 ( 
.A(n_168),
.B(n_131),
.C(n_6),
.Y(n_254)
);

MAJIxp5_ASAP7_75t_L g318 ( 
.A(n_254),
.B(n_310),
.C(n_313),
.Y(n_318)
);

HB1xp67_ASAP7_75t_L g256 ( 
.A(n_188),
.Y(n_256)
);

CKINVDCx16_ASAP7_75t_R g342 ( 
.A(n_256),
.Y(n_342)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_133),
.Y(n_257)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_257),
.Y(n_322)
);

AOI22xp5_ASAP7_75t_SL g258 ( 
.A1(n_147),
.A2(n_139),
.B1(n_134),
.B2(n_193),
.Y(n_258)
);

OAI21xp5_ASAP7_75t_SL g352 ( 
.A1(n_258),
.A2(n_272),
.B(n_278),
.Y(n_352)
);

AOI22xp33_ASAP7_75t_SL g259 ( 
.A1(n_230),
.A2(n_131),
.B1(n_6),
.B2(n_7),
.Y(n_259)
);

AOI22xp5_ASAP7_75t_SL g333 ( 
.A1(n_259),
.A2(n_285),
.B1(n_294),
.B2(n_301),
.Y(n_333)
);

NOR2xp33_ASAP7_75t_L g317 ( 
.A(n_262),
.B(n_298),
.Y(n_317)
);

CKINVDCx20_ASAP7_75t_R g263 ( 
.A(n_142),
.Y(n_263)
);

NAND2xp5_ASAP7_75t_SL g366 ( 
.A(n_263),
.B(n_276),
.Y(n_366)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_141),
.Y(n_264)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_264),
.Y(n_325)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_159),
.Y(n_265)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_265),
.Y(n_335)
);

BUFx12f_ASAP7_75t_L g266 ( 
.A(n_223),
.Y(n_266)
);

INVx5_ASAP7_75t_L g339 ( 
.A(n_266),
.Y(n_339)
);

AOI22xp5_ASAP7_75t_L g344 ( 
.A1(n_268),
.A2(n_222),
.B1(n_283),
.B2(n_252),
.Y(n_344)
);

AOI22xp33_ASAP7_75t_L g270 ( 
.A1(n_148),
.A2(n_14),
.B1(n_18),
.B2(n_19),
.Y(n_270)
);

OAI22xp5_ASAP7_75t_SL g330 ( 
.A1(n_270),
.A2(n_284),
.B1(n_211),
.B2(n_189),
.Y(n_330)
);

INVx3_ASAP7_75t_L g271 ( 
.A(n_224),
.Y(n_271)
);

INVx3_ASAP7_75t_L g321 ( 
.A(n_271),
.Y(n_321)
);

AOI22xp5_ASAP7_75t_SL g272 ( 
.A1(n_202),
.A2(n_220),
.B1(n_214),
.B2(n_184),
.Y(n_272)
);

INVx2_ASAP7_75t_L g273 ( 
.A(n_179),
.Y(n_273)
);

INVx2_ASAP7_75t_L g351 ( 
.A(n_273),
.Y(n_351)
);

INVx6_ASAP7_75t_L g274 ( 
.A(n_204),
.Y(n_274)
);

INVx3_ASAP7_75t_L g323 ( 
.A(n_274),
.Y(n_323)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_172),
.Y(n_275)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_275),
.Y(n_341)
);

CKINVDCx16_ASAP7_75t_R g276 ( 
.A(n_151),
.Y(n_276)
);

OAI21xp5_ASAP7_75t_L g278 ( 
.A1(n_138),
.A2(n_5),
.B(n_14),
.Y(n_278)
);

INVx3_ASAP7_75t_L g279 ( 
.A(n_224),
.Y(n_279)
);

INVx3_ASAP7_75t_L g362 ( 
.A(n_279),
.Y(n_362)
);

INVx1_ASAP7_75t_SL g280 ( 
.A(n_176),
.Y(n_280)
);

OAI21xp33_ASAP7_75t_L g281 ( 
.A1(n_164),
.A2(n_18),
.B(n_5),
.Y(n_281)
);

NAND2xp67_ASAP7_75t_L g282 ( 
.A(n_164),
.B(n_5),
.Y(n_282)
);

AOI22xp5_ASAP7_75t_L g284 ( 
.A1(n_182),
.A2(n_166),
.B1(n_228),
.B2(n_152),
.Y(n_284)
);

AOI22xp33_ASAP7_75t_SL g285 ( 
.A1(n_223),
.A2(n_187),
.B1(n_176),
.B2(n_153),
.Y(n_285)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_137),
.Y(n_286)
);

INVx1_ASAP7_75t_L g345 ( 
.A(n_286),
.Y(n_345)
);

INVx5_ASAP7_75t_L g287 ( 
.A(n_176),
.Y(n_287)
);

INVx3_ASAP7_75t_L g367 ( 
.A(n_287),
.Y(n_367)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_157),
.Y(n_288)
);

INVx1_ASAP7_75t_L g348 ( 
.A(n_288),
.Y(n_348)
);

NAND2xp5_ASAP7_75t_L g289 ( 
.A(n_156),
.B(n_161),
.Y(n_289)
);

NAND2xp5_ASAP7_75t_L g329 ( 
.A(n_289),
.B(n_303),
.Y(n_329)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_158),
.Y(n_290)
);

INVx1_ASAP7_75t_L g358 ( 
.A(n_290),
.Y(n_358)
);

INVx4_ASAP7_75t_L g291 ( 
.A(n_191),
.Y(n_291)
);

INVx2_ASAP7_75t_L g355 ( 
.A(n_291),
.Y(n_355)
);

BUFx4f_ASAP7_75t_SL g292 ( 
.A(n_217),
.Y(n_292)
);

CKINVDCx16_ASAP7_75t_R g353 ( 
.A(n_292),
.Y(n_353)
);

BUFx6f_ASAP7_75t_L g293 ( 
.A(n_154),
.Y(n_293)
);

INVx2_ASAP7_75t_L g365 ( 
.A(n_293),
.Y(n_365)
);

OAI22xp33_ASAP7_75t_SL g294 ( 
.A1(n_146),
.A2(n_205),
.B1(n_192),
.B2(n_165),
.Y(n_294)
);

AND2x2_ASAP7_75t_SL g295 ( 
.A(n_169),
.B(n_178),
.Y(n_295)
);

CKINVDCx16_ASAP7_75t_R g359 ( 
.A(n_295),
.Y(n_359)
);

INVx3_ASAP7_75t_L g296 ( 
.A(n_194),
.Y(n_296)
);

INVx2_ASAP7_75t_L g374 ( 
.A(n_296),
.Y(n_374)
);

INVx4_ASAP7_75t_L g297 ( 
.A(n_191),
.Y(n_297)
);

INVx1_ASAP7_75t_L g372 ( 
.A(n_297),
.Y(n_372)
);

INVx2_ASAP7_75t_L g298 ( 
.A(n_215),
.Y(n_298)
);

INVx4_ASAP7_75t_L g299 ( 
.A(n_194),
.Y(n_299)
);

NOR2xp33_ASAP7_75t_L g340 ( 
.A(n_299),
.B(n_300),
.Y(n_340)
);

INVx2_ASAP7_75t_L g300 ( 
.A(n_215),
.Y(n_300)
);

AOI22xp5_ASAP7_75t_SL g301 ( 
.A1(n_170),
.A2(n_187),
.B1(n_153),
.B2(n_186),
.Y(n_301)
);

HB1xp67_ASAP7_75t_L g302 ( 
.A(n_190),
.Y(n_302)
);

CKINVDCx20_ASAP7_75t_R g334 ( 
.A(n_302),
.Y(n_334)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_228),
.Y(n_303)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_190),
.Y(n_305)
);

NOR2xp33_ASAP7_75t_L g363 ( 
.A(n_305),
.B(n_315),
.Y(n_363)
);

NAND2xp5_ASAP7_75t_L g306 ( 
.A(n_206),
.B(n_136),
.Y(n_306)
);

NAND2xp5_ASAP7_75t_L g347 ( 
.A(n_306),
.B(n_308),
.Y(n_347)
);

AOI22xp33_ASAP7_75t_SL g307 ( 
.A1(n_195),
.A2(n_201),
.B1(n_213),
.B2(n_144),
.Y(n_307)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_195),
.Y(n_308)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_201),
.Y(n_309)
);

NAND2xp5_ASAP7_75t_L g354 ( 
.A(n_309),
.B(n_295),
.Y(n_354)
);

MAJIxp5_ASAP7_75t_L g310 ( 
.A(n_213),
.B(n_170),
.C(n_221),
.Y(n_310)
);

OAI22xp33_ASAP7_75t_SL g311 ( 
.A1(n_155),
.A2(n_150),
.B1(n_136),
.B2(n_199),
.Y(n_311)
);

AOI22x1_ASAP7_75t_L g349 ( 
.A1(n_311),
.A2(n_314),
.B1(n_261),
.B2(n_251),
.Y(n_349)
);

AND2x2_ASAP7_75t_L g313 ( 
.A(n_173),
.B(n_200),
.Y(n_313)
);

AOI22xp5_ASAP7_75t_SL g314 ( 
.A1(n_198),
.A2(n_208),
.B1(n_144),
.B2(n_145),
.Y(n_314)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_198),
.Y(n_315)
);

NOR2xp33_ASAP7_75t_L g316 ( 
.A(n_217),
.B(n_200),
.Y(n_316)
);

NOR2xp33_ASAP7_75t_SL g326 ( 
.A(n_316),
.B(n_189),
.Y(n_326)
);

MAJIxp5_ASAP7_75t_L g319 ( 
.A(n_238),
.B(n_145),
.C(n_173),
.Y(n_319)
);

MAJIxp5_ASAP7_75t_L g383 ( 
.A(n_319),
.B(n_376),
.C(n_295),
.Y(n_383)
);

AOI21xp5_ASAP7_75t_L g421 ( 
.A1(n_324),
.A2(n_280),
.B(n_313),
.Y(n_421)
);

NOR2xp33_ASAP7_75t_L g379 ( 
.A(n_326),
.B(n_350),
.Y(n_379)
);

AND2x2_ASAP7_75t_L g395 ( 
.A(n_330),
.B(n_293),
.Y(n_395)
);

OAI22xp5_ASAP7_75t_SL g331 ( 
.A1(n_268),
.A2(n_211),
.B1(n_135),
.B2(n_199),
.Y(n_331)
);

AOI22xp5_ASAP7_75t_L g391 ( 
.A1(n_331),
.A2(n_344),
.B1(n_346),
.B2(n_292),
.Y(n_391)
);

BUFx12_ASAP7_75t_L g337 ( 
.A(n_237),
.Y(n_337)
);

INVxp67_ASAP7_75t_L g394 ( 
.A(n_337),
.Y(n_394)
);

AOI21xp33_ASAP7_75t_L g343 ( 
.A1(n_234),
.A2(n_204),
.B(n_135),
.Y(n_343)
);

NOR2xp33_ASAP7_75t_SL g387 ( 
.A(n_343),
.B(n_364),
.Y(n_387)
);

OAI22xp5_ASAP7_75t_SL g346 ( 
.A1(n_306),
.A2(n_222),
.B1(n_312),
.B2(n_258),
.Y(n_346)
);

OAI22xp33_ASAP7_75t_L g419 ( 
.A1(n_349),
.A2(n_297),
.B1(n_291),
.B2(n_279),
.Y(n_419)
);

CKINVDCx20_ASAP7_75t_R g350 ( 
.A(n_255),
.Y(n_350)
);

INVx1_ASAP7_75t_L g392 ( 
.A(n_354),
.Y(n_392)
);

CKINVDCx16_ASAP7_75t_R g390 ( 
.A(n_361),
.Y(n_390)
);

NOR2xp33_ASAP7_75t_L g364 ( 
.A(n_267),
.B(n_288),
.Y(n_364)
);

NAND2xp5_ASAP7_75t_L g368 ( 
.A(n_253),
.B(n_281),
.Y(n_368)
);

NAND2xp5_ASAP7_75t_L g398 ( 
.A(n_368),
.B(n_371),
.Y(n_398)
);

NAND2xp5_ASAP7_75t_L g371 ( 
.A(n_248),
.B(n_282),
.Y(n_371)
);

NOR2xp33_ASAP7_75t_L g373 ( 
.A(n_277),
.B(n_289),
.Y(n_373)
);

NOR2xp33_ASAP7_75t_SL g424 ( 
.A(n_373),
.B(n_378),
.Y(n_424)
);

AOI22x1_ASAP7_75t_L g375 ( 
.A1(n_238),
.A2(n_235),
.B1(n_278),
.B2(n_248),
.Y(n_375)
);

OAI22xp5_ASAP7_75t_L g389 ( 
.A1(n_375),
.A2(n_300),
.B1(n_298),
.B2(n_292),
.Y(n_389)
);

MAJIxp5_ASAP7_75t_L g376 ( 
.A(n_235),
.B(n_254),
.C(n_304),
.Y(n_376)
);

NAND2xp5_ASAP7_75t_L g377 ( 
.A(n_260),
.B(n_247),
.Y(n_377)
);

NAND2xp5_ASAP7_75t_L g409 ( 
.A(n_377),
.B(n_240),
.Y(n_409)
);

NOR2xp33_ASAP7_75t_L g378 ( 
.A(n_246),
.B(n_265),
.Y(n_378)
);

OR2x2_ASAP7_75t_L g380 ( 
.A(n_361),
.B(n_272),
.Y(n_380)
);

OAI21xp5_ASAP7_75t_L g431 ( 
.A1(n_380),
.A2(n_320),
.B(n_352),
.Y(n_431)
);

XNOR2xp5_ASAP7_75t_L g381 ( 
.A(n_376),
.B(n_304),
.Y(n_381)
);

MAJIxp5_ASAP7_75t_L g429 ( 
.A(n_381),
.B(n_383),
.C(n_401),
.Y(n_429)
);

NOR2xp33_ASAP7_75t_L g382 ( 
.A(n_350),
.B(n_264),
.Y(n_382)
);

NOR2xp33_ASAP7_75t_SL g448 ( 
.A(n_382),
.B(n_388),
.Y(n_448)
);

OAI22xp5_ASAP7_75t_SL g384 ( 
.A1(n_344),
.A2(n_312),
.B1(n_284),
.B2(n_301),
.Y(n_384)
);

AOI22xp5_ASAP7_75t_L g449 ( 
.A1(n_384),
.A2(n_386),
.B1(n_391),
.B2(n_395),
.Y(n_449)
);

CKINVDCx20_ASAP7_75t_R g385 ( 
.A(n_363),
.Y(n_385)
);

NOR2xp33_ASAP7_75t_L g463 ( 
.A(n_385),
.B(n_396),
.Y(n_463)
);

OAI22xp5_ASAP7_75t_SL g386 ( 
.A1(n_347),
.A2(n_314),
.B1(n_310),
.B2(n_286),
.Y(n_386)
);

NAND2xp5_ASAP7_75t_SL g388 ( 
.A(n_329),
.B(n_308),
.Y(n_388)
);

AND2x2_ASAP7_75t_L g465 ( 
.A(n_389),
.B(n_416),
.Y(n_465)
);

NOR2xp33_ASAP7_75t_L g393 ( 
.A(n_348),
.B(n_309),
.Y(n_393)
);

NAND2xp5_ASAP7_75t_SL g433 ( 
.A(n_393),
.B(n_409),
.Y(n_433)
);

CKINVDCx20_ASAP7_75t_R g396 ( 
.A(n_356),
.Y(n_396)
);

CKINVDCx20_ASAP7_75t_R g397 ( 
.A(n_356),
.Y(n_397)
);

NOR2xp33_ASAP7_75t_L g466 ( 
.A(n_397),
.B(n_410),
.Y(n_466)
);

OAI21xp5_ASAP7_75t_SL g399 ( 
.A1(n_320),
.A2(n_275),
.B(n_241),
.Y(n_399)
);

OAI21xp5_ASAP7_75t_SL g437 ( 
.A1(n_399),
.A2(n_421),
.B(n_354),
.Y(n_437)
);

INVx4_ASAP7_75t_L g400 ( 
.A(n_323),
.Y(n_400)
);

INVx2_ASAP7_75t_L g468 ( 
.A(n_400),
.Y(n_468)
);

MAJIxp5_ASAP7_75t_L g401 ( 
.A(n_318),
.B(n_233),
.C(n_240),
.Y(n_401)
);

INVx1_ASAP7_75t_L g402 ( 
.A(n_325),
.Y(n_402)
);

INVx1_ASAP7_75t_L g432 ( 
.A(n_402),
.Y(n_432)
);

AOI22xp5_ASAP7_75t_L g403 ( 
.A1(n_346),
.A2(n_303),
.B1(n_273),
.B2(n_233),
.Y(n_403)
);

OAI22xp5_ASAP7_75t_L g428 ( 
.A1(n_403),
.A2(n_391),
.B1(n_406),
.B2(n_402),
.Y(n_428)
);

INVx1_ASAP7_75t_L g404 ( 
.A(n_325),
.Y(n_404)
);

INVx1_ASAP7_75t_L g436 ( 
.A(n_404),
.Y(n_436)
);

INVx1_ASAP7_75t_L g405 ( 
.A(n_335),
.Y(n_405)
);

INVx1_ASAP7_75t_L g438 ( 
.A(n_405),
.Y(n_438)
);

INVx1_ASAP7_75t_L g406 ( 
.A(n_335),
.Y(n_406)
);

INVx1_ASAP7_75t_L g445 ( 
.A(n_406),
.Y(n_445)
);

OAI22xp5_ASAP7_75t_L g407 ( 
.A1(n_349),
.A2(n_274),
.B1(n_249),
.B2(n_271),
.Y(n_407)
);

AOI22xp5_ASAP7_75t_L g452 ( 
.A1(n_407),
.A2(n_412),
.B1(n_419),
.B2(n_330),
.Y(n_452)
);

INVx2_ASAP7_75t_L g408 ( 
.A(n_323),
.Y(n_408)
);

INVx1_ASAP7_75t_L g459 ( 
.A(n_408),
.Y(n_459)
);

CKINVDCx20_ASAP7_75t_R g410 ( 
.A(n_366),
.Y(n_410)
);

INVx3_ASAP7_75t_L g411 ( 
.A(n_321),
.Y(n_411)
);

INVx4_ASAP7_75t_L g435 ( 
.A(n_411),
.Y(n_435)
);

OAI22xp5_ASAP7_75t_SL g412 ( 
.A1(n_347),
.A2(n_243),
.B1(n_269),
.B2(n_296),
.Y(n_412)
);

NOR2xp33_ASAP7_75t_L g413 ( 
.A(n_348),
.B(n_269),
.Y(n_413)
);

NAND2xp5_ASAP7_75t_SL g439 ( 
.A(n_413),
.B(n_417),
.Y(n_439)
);

INVx1_ASAP7_75t_L g414 ( 
.A(n_345),
.Y(n_414)
);

INVx1_ASAP7_75t_L g462 ( 
.A(n_414),
.Y(n_462)
);

INVx2_ASAP7_75t_L g415 ( 
.A(n_365),
.Y(n_415)
);

INVx1_ASAP7_75t_L g464 ( 
.A(n_415),
.Y(n_464)
);

INVx1_ASAP7_75t_L g416 ( 
.A(n_345),
.Y(n_416)
);

NAND2xp5_ASAP7_75t_SL g417 ( 
.A(n_329),
.B(n_243),
.Y(n_417)
);

INVx4_ASAP7_75t_L g418 ( 
.A(n_365),
.Y(n_418)
);

AOI22xp33_ASAP7_75t_SL g442 ( 
.A1(n_418),
.A2(n_426),
.B1(n_369),
.B2(n_332),
.Y(n_442)
);

CKINVDCx20_ASAP7_75t_R g420 ( 
.A(n_340),
.Y(n_420)
);

CKINVDCx20_ASAP7_75t_R g454 ( 
.A(n_420),
.Y(n_454)
);

NAND2xp5_ASAP7_75t_SL g422 ( 
.A(n_377),
.B(n_299),
.Y(n_422)
);

NAND2xp5_ASAP7_75t_SL g440 ( 
.A(n_422),
.B(n_359),
.Y(n_440)
);

CKINVDCx20_ASAP7_75t_R g423 ( 
.A(n_339),
.Y(n_423)
);

CKINVDCx20_ASAP7_75t_R g456 ( 
.A(n_423),
.Y(n_456)
);

HB1xp67_ASAP7_75t_L g425 ( 
.A(n_321),
.Y(n_425)
);

CKINVDCx20_ASAP7_75t_R g458 ( 
.A(n_425),
.Y(n_458)
);

AOI22xp33_ASAP7_75t_L g426 ( 
.A1(n_349),
.A2(n_242),
.B1(n_287),
.B2(n_313),
.Y(n_426)
);

CKINVDCx20_ASAP7_75t_R g427 ( 
.A(n_339),
.Y(n_427)
);

CKINVDCx16_ASAP7_75t_R g469 ( 
.A(n_427),
.Y(n_469)
);

AOI22xp5_ASAP7_75t_L g490 ( 
.A1(n_428),
.A2(n_441),
.B1(n_444),
.B2(n_447),
.Y(n_490)
);

XNOR2xp5_ASAP7_75t_L g430 ( 
.A(n_381),
.B(n_318),
.Y(n_430)
);

XNOR2xp5_ASAP7_75t_SL g475 ( 
.A(n_430),
.B(n_446),
.Y(n_475)
);

OAI21xp5_ASAP7_75t_L g488 ( 
.A1(n_431),
.A2(n_434),
.B(n_393),
.Y(n_488)
);

OAI21xp5_ASAP7_75t_L g434 ( 
.A1(n_390),
.A2(n_352),
.B(n_375),
.Y(n_434)
);

NAND2xp5_ASAP7_75t_SL g500 ( 
.A(n_437),
.B(n_322),
.Y(n_500)
);

NAND2xp5_ASAP7_75t_L g477 ( 
.A(n_440),
.B(n_457),
.Y(n_477)
);

OAI22xp5_ASAP7_75t_SL g441 ( 
.A1(n_390),
.A2(n_333),
.B1(n_332),
.B2(n_368),
.Y(n_441)
);

INVx1_ASAP7_75t_SL g493 ( 
.A(n_442),
.Y(n_493)
);

AOI22xp5_ASAP7_75t_SL g443 ( 
.A1(n_407),
.A2(n_386),
.B1(n_387),
.B2(n_389),
.Y(n_443)
);

OAI22x1_ASAP7_75t_L g492 ( 
.A1(n_443),
.A2(n_413),
.B1(n_416),
.B2(n_414),
.Y(n_492)
);

OAI22xp5_ASAP7_75t_SL g444 ( 
.A1(n_380),
.A2(n_333),
.B1(n_331),
.B2(n_375),
.Y(n_444)
);

XNOR2xp5_ASAP7_75t_L g446 ( 
.A(n_383),
.B(n_370),
.Y(n_446)
);

OAI22xp5_ASAP7_75t_SL g447 ( 
.A1(n_380),
.A2(n_371),
.B1(n_317),
.B2(n_369),
.Y(n_447)
);

XNOR2xp5_ASAP7_75t_L g450 ( 
.A(n_398),
.B(n_360),
.Y(n_450)
);

MAJIxp5_ASAP7_75t_L g472 ( 
.A(n_450),
.B(n_451),
.C(n_461),
.Y(n_472)
);

XNOR2xp5_ASAP7_75t_L g451 ( 
.A(n_398),
.B(n_319),
.Y(n_451)
);

INVx1_ASAP7_75t_L g470 ( 
.A(n_452),
.Y(n_470)
);

AOI22xp5_ASAP7_75t_L g453 ( 
.A1(n_384),
.A2(n_357),
.B1(n_334),
.B2(n_362),
.Y(n_453)
);

OAI22xp5_ASAP7_75t_SL g473 ( 
.A1(n_453),
.A2(n_467),
.B1(n_403),
.B2(n_395),
.Y(n_473)
);

AOI21xp5_ASAP7_75t_L g455 ( 
.A1(n_421),
.A2(n_357),
.B(n_353),
.Y(n_455)
);

AOI21xp5_ASAP7_75t_L g471 ( 
.A1(n_455),
.A2(n_399),
.B(n_387),
.Y(n_471)
);

OAI22xp5_ASAP7_75t_SL g457 ( 
.A1(n_392),
.A2(n_357),
.B1(n_334),
.B2(n_327),
.Y(n_457)
);

OAI22xp5_ASAP7_75t_SL g460 ( 
.A1(n_392),
.A2(n_327),
.B1(n_358),
.B2(n_362),
.Y(n_460)
);

NAND2xp5_ASAP7_75t_L g480 ( 
.A(n_460),
.B(n_404),
.Y(n_480)
);

XNOR2xp5_ASAP7_75t_L g461 ( 
.A(n_401),
.B(n_322),
.Y(n_461)
);

AOI22xp5_ASAP7_75t_L g467 ( 
.A1(n_395),
.A2(n_358),
.B1(n_372),
.B2(n_341),
.Y(n_467)
);

AO21x1_ASAP7_75t_L g536 ( 
.A1(n_471),
.A2(n_488),
.B(n_491),
.Y(n_536)
);

AND2x2_ASAP7_75t_L g522 ( 
.A(n_473),
.B(n_479),
.Y(n_522)
);

INVx1_ASAP7_75t_L g474 ( 
.A(n_432),
.Y(n_474)
);

INVx1_ASAP7_75t_L g513 ( 
.A(n_474),
.Y(n_513)
);

CKINVDCx20_ASAP7_75t_R g476 ( 
.A(n_466),
.Y(n_476)
);

NAND2xp5_ASAP7_75t_L g510 ( 
.A(n_476),
.B(n_487),
.Y(n_510)
);

AOI21xp5_ASAP7_75t_L g478 ( 
.A1(n_434),
.A2(n_427),
.B(n_423),
.Y(n_478)
);

AOI21xp5_ASAP7_75t_L g509 ( 
.A1(n_478),
.A2(n_488),
.B(n_502),
.Y(n_509)
);

OA21x2_ASAP7_75t_L g479 ( 
.A1(n_465),
.A2(n_395),
.B(n_379),
.Y(n_479)
);

INVx1_ASAP7_75t_L g512 ( 
.A(n_480),
.Y(n_512)
);

CKINVDCx16_ASAP7_75t_R g481 ( 
.A(n_463),
.Y(n_481)
);

INVx1_ASAP7_75t_L g516 ( 
.A(n_481),
.Y(n_516)
);

INVx1_ASAP7_75t_L g482 ( 
.A(n_432),
.Y(n_482)
);

INVx1_ASAP7_75t_L g534 ( 
.A(n_482),
.Y(n_534)
);

OAI32xp33_ASAP7_75t_L g483 ( 
.A1(n_465),
.A2(n_409),
.A3(n_379),
.B1(n_382),
.B2(n_424),
.Y(n_483)
);

INVxp67_ASAP7_75t_L g535 ( 
.A(n_483),
.Y(n_535)
);

NAND2xp5_ASAP7_75t_L g484 ( 
.A(n_454),
.B(n_433),
.Y(n_484)
);

INVx1_ASAP7_75t_L g540 ( 
.A(n_484),
.Y(n_540)
);

OAI22xp5_ASAP7_75t_L g485 ( 
.A1(n_449),
.A2(n_388),
.B1(n_417),
.B2(n_422),
.Y(n_485)
);

OAI22xp5_ASAP7_75t_L g543 ( 
.A1(n_485),
.A2(n_495),
.B1(n_497),
.B2(n_508),
.Y(n_543)
);

INVx1_ASAP7_75t_L g486 ( 
.A(n_436),
.Y(n_486)
);

INVx1_ASAP7_75t_L g541 ( 
.A(n_486),
.Y(n_541)
);

NAND2xp5_ASAP7_75t_L g487 ( 
.A(n_454),
.B(n_420),
.Y(n_487)
);

CKINVDCx20_ASAP7_75t_R g489 ( 
.A(n_460),
.Y(n_489)
);

NOR2xp33_ASAP7_75t_L g525 ( 
.A(n_489),
.B(n_494),
.Y(n_525)
);

NAND2xp5_ASAP7_75t_L g491 ( 
.A(n_439),
.B(n_405),
.Y(n_491)
);

AOI22xp5_ASAP7_75t_SL g518 ( 
.A1(n_492),
.A2(n_457),
.B1(n_469),
.B2(n_453),
.Y(n_518)
);

BUFx24_ASAP7_75t_SL g494 ( 
.A(n_450),
.Y(n_494)
);

INVx1_ASAP7_75t_L g495 ( 
.A(n_436),
.Y(n_495)
);

XOR2xp5_ASAP7_75t_L g496 ( 
.A(n_429),
.B(n_424),
.Y(n_496)
);

MAJIxp5_ASAP7_75t_L g517 ( 
.A(n_496),
.B(n_498),
.C(n_499),
.Y(n_517)
);

INVx1_ASAP7_75t_L g497 ( 
.A(n_438),
.Y(n_497)
);

XOR2xp5_ASAP7_75t_L g498 ( 
.A(n_429),
.B(n_412),
.Y(n_498)
);

MAJIxp5_ASAP7_75t_L g499 ( 
.A(n_430),
.B(n_410),
.C(n_385),
.Y(n_499)
);

AOI21xp33_ASAP7_75t_L g532 ( 
.A1(n_500),
.A2(n_394),
.B(n_464),
.Y(n_532)
);

XNOR2xp5_ASAP7_75t_L g501 ( 
.A(n_446),
.B(n_341),
.Y(n_501)
);

XOR2xp5_ASAP7_75t_L g514 ( 
.A(n_501),
.B(n_447),
.Y(n_514)
);

NAND2xp5_ASAP7_75t_L g502 ( 
.A(n_448),
.B(n_456),
.Y(n_502)
);

CKINVDCx20_ASAP7_75t_R g539 ( 
.A(n_502),
.Y(n_539)
);

MAJIxp5_ASAP7_75t_L g503 ( 
.A(n_461),
.B(n_451),
.C(n_431),
.Y(n_503)
);

MAJIxp5_ASAP7_75t_L g528 ( 
.A(n_503),
.B(n_504),
.C(n_458),
.Y(n_528)
);

MAJIxp5_ASAP7_75t_L g504 ( 
.A(n_440),
.B(n_437),
.C(n_455),
.Y(n_504)
);

NOR2xp33_ASAP7_75t_L g505 ( 
.A(n_448),
.B(n_342),
.Y(n_505)
);

CKINVDCx16_ASAP7_75t_R g531 ( 
.A(n_505),
.Y(n_531)
);

CKINVDCx20_ASAP7_75t_R g506 ( 
.A(n_456),
.Y(n_506)
);

CKINVDCx20_ASAP7_75t_R g542 ( 
.A(n_506),
.Y(n_542)
);

OAI22xp5_ASAP7_75t_SL g507 ( 
.A1(n_449),
.A2(n_396),
.B1(n_397),
.B2(n_408),
.Y(n_507)
);

AOI22xp5_ASAP7_75t_L g511 ( 
.A1(n_507),
.A2(n_473),
.B1(n_428),
.B2(n_489),
.Y(n_511)
);

INVx1_ASAP7_75t_L g508 ( 
.A(n_438),
.Y(n_508)
);

AOI21xp33_ASAP7_75t_L g570 ( 
.A1(n_509),
.A2(n_532),
.B(n_474),
.Y(n_570)
);

OAI22xp5_ASAP7_75t_SL g546 ( 
.A1(n_511),
.A2(n_515),
.B1(n_518),
.B2(n_521),
.Y(n_546)
);

XNOR2xp5_ASAP7_75t_L g559 ( 
.A(n_514),
.B(n_528),
.Y(n_559)
);

AOI22xp5_ASAP7_75t_L g515 ( 
.A1(n_470),
.A2(n_444),
.B1(n_465),
.B2(n_441),
.Y(n_515)
);

XNOR2xp5_ASAP7_75t_SL g519 ( 
.A(n_475),
.B(n_443),
.Y(n_519)
);

XNOR2xp5_ASAP7_75t_SL g549 ( 
.A(n_519),
.B(n_504),
.Y(n_549)
);

FAx1_ASAP7_75t_SL g520 ( 
.A(n_503),
.B(n_445),
.CI(n_462),
.CON(n_520),
.SN(n_520)
);

NAND2xp5_ASAP7_75t_L g553 ( 
.A(n_520),
.B(n_523),
.Y(n_553)
);

AOI22xp5_ASAP7_75t_L g521 ( 
.A1(n_470),
.A2(n_452),
.B1(n_469),
.B2(n_458),
.Y(n_521)
);

OAI21xp5_ASAP7_75t_L g523 ( 
.A1(n_478),
.A2(n_467),
.B(n_462),
.Y(n_523)
);

XNOR2xp5_ASAP7_75t_L g524 ( 
.A(n_496),
.B(n_445),
.Y(n_524)
);

XOR2xp5_ASAP7_75t_L g550 ( 
.A(n_524),
.B(n_526),
.Y(n_550)
);

XOR2xp5_ASAP7_75t_L g526 ( 
.A(n_475),
.B(n_425),
.Y(n_526)
);

XOR2x2_ASAP7_75t_L g527 ( 
.A(n_498),
.B(n_459),
.Y(n_527)
);

NOR2xp33_ASAP7_75t_L g567 ( 
.A(n_527),
.B(n_508),
.Y(n_567)
);

AOI22xp5_ASAP7_75t_L g529 ( 
.A1(n_490),
.A2(n_459),
.B1(n_464),
.B2(n_468),
.Y(n_529)
);

AOI22xp5_ASAP7_75t_L g565 ( 
.A1(n_529),
.A2(n_530),
.B1(n_533),
.B2(n_545),
.Y(n_565)
);

AOI22xp5_ASAP7_75t_L g530 ( 
.A1(n_490),
.A2(n_492),
.B1(n_479),
.B2(n_485),
.Y(n_530)
);

AOI22xp5_ASAP7_75t_L g533 ( 
.A1(n_479),
.A2(n_468),
.B1(n_435),
.B2(n_400),
.Y(n_533)
);

MAJIxp5_ASAP7_75t_L g537 ( 
.A(n_472),
.B(n_372),
.C(n_355),
.Y(n_537)
);

MAJIxp5_ASAP7_75t_L g547 ( 
.A(n_537),
.B(n_544),
.C(n_506),
.Y(n_547)
);

XOR2xp5_ASAP7_75t_L g538 ( 
.A(n_472),
.B(n_355),
.Y(n_538)
);

XOR2xp5_ASAP7_75t_L g568 ( 
.A(n_538),
.B(n_497),
.Y(n_568)
);

MAJIxp5_ASAP7_75t_L g544 ( 
.A(n_501),
.B(n_374),
.C(n_411),
.Y(n_544)
);

AOI22xp5_ASAP7_75t_L g545 ( 
.A1(n_507),
.A2(n_435),
.B1(n_400),
.B2(n_415),
.Y(n_545)
);

MAJIxp5_ASAP7_75t_L g590 ( 
.A(n_547),
.B(n_555),
.C(n_558),
.Y(n_590)
);

INVx1_ASAP7_75t_L g548 ( 
.A(n_510),
.Y(n_548)
);

INVx1_ASAP7_75t_L g579 ( 
.A(n_548),
.Y(n_579)
);

XOR2xp5_ASAP7_75t_L g584 ( 
.A(n_549),
.B(n_557),
.Y(n_584)
);

CKINVDCx14_ASAP7_75t_R g551 ( 
.A(n_510),
.Y(n_551)
);

NAND2xp5_ASAP7_75t_L g578 ( 
.A(n_551),
.B(n_552),
.Y(n_578)
);

CKINVDCx14_ASAP7_75t_R g552 ( 
.A(n_542),
.Y(n_552)
);

INVx1_ASAP7_75t_L g554 ( 
.A(n_540),
.Y(n_554)
);

INVx1_ASAP7_75t_L g587 ( 
.A(n_554),
.Y(n_587)
);

MAJIxp5_ASAP7_75t_L g555 ( 
.A(n_517),
.B(n_499),
.C(n_471),
.Y(n_555)
);

AOI22xp5_ASAP7_75t_L g556 ( 
.A1(n_535),
.A2(n_477),
.B1(n_493),
.B2(n_476),
.Y(n_556)
);

OAI22xp5_ASAP7_75t_SL g577 ( 
.A1(n_556),
.A2(n_560),
.B1(n_533),
.B2(n_518),
.Y(n_577)
);

XNOR2xp5_ASAP7_75t_SL g557 ( 
.A(n_526),
.B(n_483),
.Y(n_557)
);

MAJIxp5_ASAP7_75t_L g558 ( 
.A(n_517),
.B(n_487),
.C(n_491),
.Y(n_558)
);

AOI22xp5_ASAP7_75t_L g560 ( 
.A1(n_535),
.A2(n_477),
.B1(n_493),
.B2(n_484),
.Y(n_560)
);

INVx1_ASAP7_75t_L g561 ( 
.A(n_540),
.Y(n_561)
);

INVx2_ASAP7_75t_L g585 ( 
.A(n_561),
.Y(n_585)
);

XNOR2xp5_ASAP7_75t_SL g562 ( 
.A(n_514),
.B(n_481),
.Y(n_562)
);

XOR2xp5_ASAP7_75t_L g597 ( 
.A(n_562),
.B(n_567),
.Y(n_597)
);

XNOR2xp5_ASAP7_75t_L g563 ( 
.A(n_538),
.B(n_480),
.Y(n_563)
);

XNOR2xp5_ASAP7_75t_L g582 ( 
.A(n_563),
.B(n_572),
.Y(n_582)
);

INVx1_ASAP7_75t_L g564 ( 
.A(n_541),
.Y(n_564)
);

NAND2xp5_ASAP7_75t_L g594 ( 
.A(n_564),
.B(n_571),
.Y(n_594)
);

BUFx6f_ASAP7_75t_L g566 ( 
.A(n_516),
.Y(n_566)
);

CKINVDCx20_ASAP7_75t_R g580 ( 
.A(n_566),
.Y(n_580)
);

XOR2xp5_ASAP7_75t_L g601 ( 
.A(n_568),
.B(n_534),
.Y(n_601)
);

AOI22xp5_ASAP7_75t_L g569 ( 
.A1(n_539),
.A2(n_495),
.B1(n_486),
.B2(n_482),
.Y(n_569)
);

INVxp67_ASAP7_75t_L g600 ( 
.A(n_569),
.Y(n_600)
);

OAI21xp5_ASAP7_75t_L g591 ( 
.A1(n_570),
.A2(n_523),
.B(n_530),
.Y(n_591)
);

INVx2_ASAP7_75t_L g571 ( 
.A(n_513),
.Y(n_571)
);

XNOR2xp5_ASAP7_75t_L g572 ( 
.A(n_524),
.B(n_528),
.Y(n_572)
);

INVx1_ASAP7_75t_L g573 ( 
.A(n_541),
.Y(n_573)
);

NOR2xp33_ASAP7_75t_SL g581 ( 
.A(n_573),
.B(n_512),
.Y(n_581)
);

MAJIxp5_ASAP7_75t_L g574 ( 
.A(n_537),
.B(n_374),
.C(n_367),
.Y(n_574)
);

MAJIxp5_ASAP7_75t_L g596 ( 
.A(n_574),
.B(n_575),
.C(n_576),
.Y(n_596)
);

MAJIxp5_ASAP7_75t_L g575 ( 
.A(n_527),
.B(n_367),
.C(n_336),
.Y(n_575)
);

MAJIxp5_ASAP7_75t_L g576 ( 
.A(n_519),
.B(n_336),
.C(n_328),
.Y(n_576)
);

AOI22xp5_ASAP7_75t_L g605 ( 
.A1(n_577),
.A2(n_588),
.B1(n_591),
.B2(n_595),
.Y(n_605)
);

INVx1_ASAP7_75t_L g604 ( 
.A(n_581),
.Y(n_604)
);

NOR2xp33_ASAP7_75t_SL g583 ( 
.A(n_558),
.B(n_525),
.Y(n_583)
);

NAND2xp5_ASAP7_75t_SL g607 ( 
.A(n_583),
.B(n_562),
.Y(n_607)
);

AOI21xp5_ASAP7_75t_L g586 ( 
.A1(n_553),
.A2(n_509),
.B(n_536),
.Y(n_586)
);

NAND2xp5_ASAP7_75t_L g608 ( 
.A(n_586),
.B(n_598),
.Y(n_608)
);

AOI22xp5_ASAP7_75t_L g588 ( 
.A1(n_546),
.A2(n_522),
.B1(n_512),
.B2(n_511),
.Y(n_588)
);

XNOR2xp5_ASAP7_75t_L g589 ( 
.A(n_555),
.B(n_536),
.Y(n_589)
);

XNOR2xp5_ASAP7_75t_L g610 ( 
.A(n_589),
.B(n_599),
.Y(n_610)
);

AND2x2_ASAP7_75t_L g592 ( 
.A(n_565),
.B(n_529),
.Y(n_592)
);

INVx1_ASAP7_75t_L g611 ( 
.A(n_592),
.Y(n_611)
);

INVx13_ASAP7_75t_L g593 ( 
.A(n_566),
.Y(n_593)
);

INVxp67_ASAP7_75t_SL g602 ( 
.A(n_593),
.Y(n_602)
);

AOI22xp5_ASAP7_75t_L g595 ( 
.A1(n_560),
.A2(n_522),
.B1(n_543),
.B2(n_515),
.Y(n_595)
);

MAJIxp5_ASAP7_75t_L g598 ( 
.A(n_559),
.B(n_544),
.C(n_520),
.Y(n_598)
);

AOI22xp5_ASAP7_75t_L g599 ( 
.A1(n_556),
.A2(n_522),
.B1(n_521),
.B2(n_575),
.Y(n_599)
);

XNOR2xp5_ASAP7_75t_L g618 ( 
.A(n_601),
.B(n_351),
.Y(n_618)
);

NOR2xp33_ASAP7_75t_L g603 ( 
.A(n_580),
.B(n_531),
.Y(n_603)
);

NOR2xp33_ASAP7_75t_SL g626 ( 
.A(n_603),
.B(n_607),
.Y(n_626)
);

MAJIxp5_ASAP7_75t_L g606 ( 
.A(n_590),
.B(n_547),
.C(n_572),
.Y(n_606)
);

MAJIxp5_ASAP7_75t_L g630 ( 
.A(n_606),
.B(n_609),
.C(n_613),
.Y(n_630)
);

MAJIxp5_ASAP7_75t_L g609 ( 
.A(n_590),
.B(n_559),
.C(n_574),
.Y(n_609)
);

NAND2xp5_ASAP7_75t_SL g612 ( 
.A(n_589),
.B(n_563),
.Y(n_612)
);

NOR2xp33_ASAP7_75t_SL g631 ( 
.A(n_612),
.B(n_616),
.Y(n_631)
);

MAJIxp5_ASAP7_75t_L g613 ( 
.A(n_582),
.B(n_568),
.C(n_550),
.Y(n_613)
);

MAJIxp5_ASAP7_75t_L g614 ( 
.A(n_582),
.B(n_550),
.C(n_557),
.Y(n_614)
);

MAJIxp5_ASAP7_75t_L g636 ( 
.A(n_614),
.B(n_617),
.C(n_620),
.Y(n_636)
);

XOR2xp5_ASAP7_75t_L g615 ( 
.A(n_586),
.B(n_576),
.Y(n_615)
);

XOR2xp5_ASAP7_75t_L g623 ( 
.A(n_615),
.B(n_618),
.Y(n_623)
);

NOR2xp33_ASAP7_75t_SL g616 ( 
.A(n_578),
.B(n_520),
.Y(n_616)
);

MAJIxp5_ASAP7_75t_L g617 ( 
.A(n_596),
.B(n_549),
.C(n_545),
.Y(n_617)
);

XOR2xp5_ASAP7_75t_L g619 ( 
.A(n_598),
.B(n_338),
.Y(n_619)
);

XOR2xp5_ASAP7_75t_L g633 ( 
.A(n_619),
.B(n_588),
.Y(n_633)
);

MAJIxp5_ASAP7_75t_L g620 ( 
.A(n_596),
.B(n_418),
.C(n_351),
.Y(n_620)
);

MAJIxp5_ASAP7_75t_L g621 ( 
.A(n_601),
.B(n_418),
.C(n_338),
.Y(n_621)
);

MAJIxp5_ASAP7_75t_L g637 ( 
.A(n_621),
.B(n_597),
.C(n_577),
.Y(n_637)
);

XNOR2xp5_ASAP7_75t_L g622 ( 
.A(n_597),
.B(n_337),
.Y(n_622)
);

NOR2xp33_ASAP7_75t_L g632 ( 
.A(n_622),
.B(n_584),
.Y(n_632)
);

OAI22xp5_ASAP7_75t_L g624 ( 
.A1(n_604),
.A2(n_579),
.B1(n_600),
.B2(n_595),
.Y(n_624)
);

NAND2xp5_ASAP7_75t_L g641 ( 
.A(n_624),
.B(n_625),
.Y(n_641)
);

INVx1_ASAP7_75t_L g625 ( 
.A(n_602),
.Y(n_625)
);

INVx1_ASAP7_75t_L g627 ( 
.A(n_611),
.Y(n_627)
);

NAND2xp5_ASAP7_75t_L g647 ( 
.A(n_627),
.B(n_628),
.Y(n_647)
);

AND2x2_ASAP7_75t_L g628 ( 
.A(n_621),
.B(n_592),
.Y(n_628)
);

NAND2xp5_ASAP7_75t_L g629 ( 
.A(n_610),
.B(n_585),
.Y(n_629)
);

NAND2xp5_ASAP7_75t_L g650 ( 
.A(n_629),
.B(n_632),
.Y(n_650)
);

XNOR2xp5_ASAP7_75t_L g640 ( 
.A(n_633),
.B(n_637),
.Y(n_640)
);

INVx6_ASAP7_75t_L g634 ( 
.A(n_608),
.Y(n_634)
);

NOR2xp33_ASAP7_75t_L g645 ( 
.A(n_634),
.B(n_620),
.Y(n_645)
);

OAI22xp5_ASAP7_75t_L g635 ( 
.A1(n_605),
.A2(n_600),
.B1(n_599),
.B2(n_587),
.Y(n_635)
);

NAND2xp5_ASAP7_75t_SL g646 ( 
.A(n_635),
.B(n_638),
.Y(n_646)
);

NOR2xp33_ASAP7_75t_L g638 ( 
.A(n_606),
.B(n_591),
.Y(n_638)
);

OAI21xp5_ASAP7_75t_L g639 ( 
.A1(n_610),
.A2(n_592),
.B(n_584),
.Y(n_639)
);

AOI21xp5_ASAP7_75t_L g652 ( 
.A1(n_639),
.A2(n_266),
.B(n_633),
.Y(n_652)
);

MAJIxp5_ASAP7_75t_L g642 ( 
.A(n_630),
.B(n_609),
.C(n_619),
.Y(n_642)
);

NAND2xp5_ASAP7_75t_L g653 ( 
.A(n_642),
.B(n_644),
.Y(n_653)
);

OAI22xp5_ASAP7_75t_L g643 ( 
.A1(n_634),
.A2(n_585),
.B1(n_617),
.B2(n_615),
.Y(n_643)
);

INVx1_ASAP7_75t_L g657 ( 
.A(n_643),
.Y(n_657)
);

OAI22xp5_ASAP7_75t_SL g644 ( 
.A1(n_627),
.A2(n_594),
.B1(n_614),
.B2(n_613),
.Y(n_644)
);

NAND2xp5_ASAP7_75t_L g654 ( 
.A(n_645),
.B(n_648),
.Y(n_654)
);

MAJIxp5_ASAP7_75t_L g648 ( 
.A(n_630),
.B(n_594),
.C(n_593),
.Y(n_648)
);

MAJIxp5_ASAP7_75t_L g649 ( 
.A(n_636),
.B(n_337),
.C(n_245),
.Y(n_649)
);

NAND2xp5_ASAP7_75t_L g659 ( 
.A(n_649),
.B(n_651),
.Y(n_659)
);

MAJIxp5_ASAP7_75t_L g651 ( 
.A(n_636),
.B(n_245),
.C(n_266),
.Y(n_651)
);

XOR2xp5_ASAP7_75t_L g656 ( 
.A(n_652),
.B(n_625),
.Y(n_656)
);

NOR2xp33_ASAP7_75t_L g655 ( 
.A(n_648),
.B(n_631),
.Y(n_655)
);

CKINVDCx20_ASAP7_75t_R g666 ( 
.A(n_655),
.Y(n_666)
);

XOR2xp5_ASAP7_75t_L g664 ( 
.A(n_656),
.B(n_660),
.Y(n_664)
);

NAND2xp5_ASAP7_75t_SL g658 ( 
.A(n_646),
.B(n_626),
.Y(n_658)
);

AOI21xp5_ASAP7_75t_L g667 ( 
.A1(n_658),
.A2(n_661),
.B(n_651),
.Y(n_667)
);

MAJIxp5_ASAP7_75t_L g660 ( 
.A(n_642),
.B(n_629),
.C(n_637),
.Y(n_660)
);

MAJIxp5_ASAP7_75t_L g661 ( 
.A(n_640),
.B(n_628),
.C(n_623),
.Y(n_661)
);

MAJIxp5_ASAP7_75t_L g662 ( 
.A(n_660),
.B(n_640),
.C(n_644),
.Y(n_662)
);

INVxp33_ASAP7_75t_L g669 ( 
.A(n_662),
.Y(n_669)
);

MAJIxp5_ASAP7_75t_L g663 ( 
.A(n_653),
.B(n_650),
.C(n_641),
.Y(n_663)
);

A2O1A1O1Ixp25_ASAP7_75t_L g670 ( 
.A1(n_663),
.A2(n_665),
.B(n_661),
.C(n_659),
.D(n_649),
.Y(n_670)
);

OAI211xp5_ASAP7_75t_L g665 ( 
.A1(n_657),
.A2(n_647),
.B(n_639),
.C(n_626),
.Y(n_665)
);

AO21x1_ASAP7_75t_L g668 ( 
.A1(n_667),
.A2(n_654),
.B(n_666),
.Y(n_668)
);

OAI21xp5_ASAP7_75t_L g671 ( 
.A1(n_668),
.A2(n_670),
.B(n_665),
.Y(n_671)
);

XNOR2xp5_ASAP7_75t_L g673 ( 
.A(n_671),
.B(n_672),
.Y(n_673)
);

MAJIxp5_ASAP7_75t_L g672 ( 
.A(n_669),
.B(n_664),
.C(n_656),
.Y(n_672)
);

XOR2xp5_ASAP7_75t_L g674 ( 
.A(n_673),
.B(n_628),
.Y(n_674)
);

XNOR2xp5_ASAP7_75t_L g675 ( 
.A(n_674),
.B(n_623),
.Y(n_675)
);


endmodule