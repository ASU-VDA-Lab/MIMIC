module fake_aes_12375_n_727 (n_44, n_81, n_69, n_22, n_57, n_88, n_52, n_26, n_50, n_33, n_73, n_49, n_80, n_60, n_41, n_35, n_94, n_65, n_9, n_10, n_19, n_87, n_74, n_7, n_29, n_45, n_85, n_62, n_36, n_47, n_37, n_34, n_5, n_23, n_8, n_91, n_16, n_13, n_70, n_17, n_63, n_14, n_71, n_90, n_56, n_42, n_24, n_78, n_6, n_4, n_40, n_79, n_38, n_64, n_46, n_31, n_58, n_32, n_0, n_84, n_55, n_12, n_86, n_75, n_72, n_43, n_76, n_89, n_68, n_27, n_53, n_67, n_77, n_20, n_2, n_54, n_83, n_28, n_48, n_92, n_11, n_25, n_30, n_59, n_3, n_18, n_66, n_1, n_82, n_15, n_61, n_21, n_93, n_51, n_39, n_727);
input n_44;
input n_81;
input n_69;
input n_22;
input n_57;
input n_88;
input n_52;
input n_26;
input n_50;
input n_33;
input n_73;
input n_49;
input n_80;
input n_60;
input n_41;
input n_35;
input n_94;
input n_65;
input n_9;
input n_10;
input n_19;
input n_87;
input n_74;
input n_7;
input n_29;
input n_45;
input n_85;
input n_62;
input n_36;
input n_47;
input n_37;
input n_34;
input n_5;
input n_23;
input n_8;
input n_91;
input n_16;
input n_13;
input n_70;
input n_17;
input n_63;
input n_14;
input n_71;
input n_90;
input n_56;
input n_42;
input n_24;
input n_78;
input n_6;
input n_4;
input n_40;
input n_79;
input n_38;
input n_64;
input n_46;
input n_31;
input n_58;
input n_32;
input n_0;
input n_84;
input n_55;
input n_12;
input n_86;
input n_75;
input n_72;
input n_43;
input n_76;
input n_89;
input n_68;
input n_27;
input n_53;
input n_67;
input n_77;
input n_20;
input n_2;
input n_54;
input n_83;
input n_28;
input n_48;
input n_92;
input n_11;
input n_25;
input n_30;
input n_59;
input n_3;
input n_18;
input n_66;
input n_1;
input n_82;
input n_15;
input n_61;
input n_21;
input n_93;
input n_51;
input n_39;
output n_727;
wire n_117;
wire n_663;
wire n_707;
wire n_361;
wire n_513;
wire n_185;
wire n_705;
wire n_603;
wire n_604;
wire n_590;
wire n_407;
wire n_646;
wire n_284;
wire n_278;
wire n_500;
wire n_114;
wire n_607;
wire n_125;
wire n_431;
wire n_484;
wire n_161;
wire n_496;
wire n_667;
wire n_177;
wire n_130;
wire n_189;
wire n_311;
wire n_292;
wire n_309;
wire n_160;
wire n_701;
wire n_612;
wire n_154;
wire n_328;
wire n_655;
wire n_468;
wire n_523;
wire n_229;
wire n_336;
wire n_464;
wire n_448;
wire n_645;
wire n_348;
wire n_252;
wire n_152;
wire n_113;
wire n_637;
wire n_353;
wire n_564;
wire n_528;
wire n_206;
wire n_288;
wire n_383;
wire n_661;
wire n_672;
wire n_532;
wire n_627;
wire n_544;
wire n_400;
wire n_296;
wire n_157;
wire n_202;
wire n_386;
wire n_432;
wire n_142;
wire n_659;
wire n_232;
wire n_462;
wire n_316;
wire n_545;
wire n_211;
wire n_334;
wire n_389;
wire n_548;
wire n_436;
wire n_588;
wire n_275;
wire n_715;
wire n_463;
wire n_131;
wire n_112;
wire n_205;
wire n_330;
wire n_587;
wire n_662;
wire n_162;
wire n_678;
wire n_387;
wire n_163;
wire n_434;
wire n_105;
wire n_227;
wire n_384;
wire n_476;
wire n_617;
wire n_231;
wire n_452;
wire n_518;
wire n_547;
wire n_298;
wire n_628;
wire n_411;
wire n_598;
wire n_144;
wire n_183;
wire n_489;
wire n_199;
wire n_351;
wire n_401;
wire n_100;
wire n_461;
wire n_305;
wire n_599;
wire n_228;
wire n_724;
wire n_360;
wire n_345;
wire n_236;
wire n_340;
wire n_481;
wire n_443;
wire n_150;
wire n_373;
wire n_576;
wire n_694;
wire n_301;
wire n_222;
wire n_234;
wire n_465;
wire n_609;
wire n_636;
wire n_366;
wire n_596;
wire n_286;
wire n_190;
wire n_246;
wire n_321;
wire n_702;
wire n_572;
wire n_324;
wire n_392;
wire n_668;
wire n_652;
wire n_279;
wire n_303;
wire n_437;
wire n_512;
wire n_326;
wire n_289;
wire n_333;
wire n_249;
wire n_680;
wire n_642;
wire n_586;
wire n_671;
wire n_244;
wire n_540;
wire n_563;
wire n_638;
wire n_119;
wire n_141;
wire n_517;
wire n_560;
wire n_479;
wire n_97;
wire n_167;
wire n_623;
wire n_593;
wire n_697;
wire n_554;
wire n_726;
wire n_712;
wire n_447;
wire n_608;
wire n_171;
wire n_567;
wire n_196;
wire n_580;
wire n_192;
wire n_502;
wire n_543;
wire n_312;
wire n_455;
wire n_529;
wire n_630;
wire n_137;
wire n_511;
wire n_277;
wire n_467;
wire n_692;
wire n_647;
wire n_367;
wire n_644;
wire n_250;
wire n_314;
wire n_237;
wire n_181;
wire n_101;
wire n_255;
wire n_426;
wire n_624;
wire n_725;
wire n_108;
wire n_116;
wire n_230;
wire n_209;
wire n_274;
wire n_282;
wire n_319;
wire n_499;
wire n_417;
wire n_241;
wire n_575;
wire n_95;
wire n_238;
wire n_711;
wire n_318;
wire n_471;
wire n_632;
wire n_293;
wire n_506;
wire n_533;
wire n_135;
wire n_393;
wire n_490;
wire n_247;
wire n_613;
wire n_648;
wire n_381;
wire n_550;
wire n_304;
wire n_399;
wire n_665;
wire n_571;
wire n_294;
wire n_459;
wire n_313;
wire n_210;
wire n_184;
wire n_322;
wire n_310;
wire n_708;
wire n_191;
wire n_307;
wire n_634;
wire n_610;
wire n_696;
wire n_474;
wire n_354;
wire n_402;
wire n_413;
wire n_676;
wire n_391;
wire n_427;
wire n_460;
wire n_478;
wire n_235;
wire n_243;
wire n_415;
wire n_394;
wire n_482;
wire n_442;
wire n_331;
wire n_485;
wire n_703;
wire n_352;
wire n_619;
wire n_268;
wire n_174;
wire n_501;
wire n_248;
wire n_299;
wire n_338;
wire n_519;
wire n_699;
wire n_693;
wire n_256;
wire n_551;
wire n_404;
wire n_369;
wire n_509;
wire n_651;
wire n_674;
wire n_172;
wire n_329;
wire n_251;
wire n_635;
wire n_689;
wire n_525;
wire n_218;
wire n_507;
wire n_605;
wire n_719;
wire n_611;
wire n_704;
wire n_633;
wire n_271;
wire n_626;
wire n_302;
wire n_466;
wire n_710;
wire n_270;
wire n_685;
wire n_362;
wire n_153;
wire n_259;
wire n_308;
wire n_546;
wire n_412;
wire n_664;
wire n_140;
wire n_207;
wire n_565;
wire n_224;
wire n_96;
wire n_219;
wire n_475;
wire n_578;
wire n_133;
wire n_149;
wire n_542;
wire n_537;
wire n_214;
wire n_204;
wire n_660;
wire n_430;
wire n_450;
wire n_579;
wire n_107;
wire n_403;
wire n_557;
wire n_516;
wire n_254;
wire n_549;
wire n_622;
wire n_262;
wire n_556;
wire n_239;
wire n_439;
wire n_601;
wire n_379;
wire n_641;
wire n_614;
wire n_527;
wire n_98;
wire n_526;
wire n_276;
wire n_649;
wire n_320;
wire n_285;
wire n_195;
wire n_165;
wire n_420;
wire n_423;
wire n_342;
wire n_446;
wire n_621;
wire n_666;
wire n_370;
wire n_589;
wire n_643;
wire n_574;
wire n_217;
wire n_139;
wire n_388;
wire n_454;
wire n_687;
wire n_193;
wire n_273;
wire n_505;
wire n_706;
wire n_390;
wire n_682;
wire n_120;
wire n_514;
wire n_486;
wire n_720;
wire n_568;
wire n_245;
wire n_357;
wire n_653;
wire n_716;
wire n_260;
wire n_539;
wire n_197;
wire n_201;
wire n_591;
wire n_317;
wire n_416;
wire n_374;
wire n_718;
wire n_111;
wire n_536;
wire n_265;
wire n_264;
wire n_522;
wire n_208;
wire n_200;
wire n_573;
wire n_126;
wire n_673;
wire n_669;
wire n_178;
wire n_616;
wire n_118;
wire n_365;
wire n_717;
wire n_541;
wire n_179;
wire n_315;
wire n_363;
wire n_409;
wire n_143;
wire n_295;
wire n_654;
wire n_263;
wire n_166;
wire n_495;
wire n_186;
wire n_364;
wire n_428;
wire n_566;
wire n_376;
wire n_639;
wire n_552;
wire n_677;
wire n_344;
wire n_136;
wire n_503;
wire n_283;
wire n_520;
wire n_681;
wire n_435;
wire n_216;
wire n_577;
wire n_147;
wire n_148;
wire n_615;
wire n_212;
wire n_472;
wire n_419;
wire n_396;
wire n_168;
wire n_477;
wire n_508;
wire n_570;
wire n_398;
wire n_445;
wire n_656;
wire n_438;
wire n_134;
wire n_721;
wire n_640;
wire n_429;
wire n_488;
wire n_233;
wire n_686;
wire n_684;
wire n_440;
wire n_106;
wire n_553;
wire n_173;
wire n_422;
wire n_679;
wire n_327;
wire n_325;
wire n_349;
wire n_498;
wire n_597;
wire n_723;
wire n_225;
wire n_535;
wire n_530;
wire n_220;
wire n_358;
wire n_267;
wire n_221;
wire n_456;
wire n_203;
wire n_102;
wire n_449;
wire n_115;
wire n_300;
wire n_158;
wire n_524;
wire n_121;
wire n_584;
wire n_497;
wire n_339;
wire n_657;
wire n_583;
wire n_620;
wire n_240;
wire n_378;
wire n_582;
wire n_359;
wire n_346;
wire n_103;
wire n_180;
wire n_441;
wire n_104;
wire n_561;
wire n_335;
wire n_272;
wire n_700;
wire n_594;
wire n_534;
wire n_531;
wire n_146;
wire n_397;
wire n_306;
wire n_215;
wire n_242;
wire n_155;
wire n_602;
wire n_198;
wire n_169;
wire n_424;
wire n_714;
wire n_629;
wire n_156;
wire n_124;
wire n_569;
wire n_297;
wire n_128;
wire n_129;
wire n_410;
wire n_188;
wire n_377;
wire n_510;
wire n_343;
wire n_127;
wire n_675;
wire n_291;
wire n_170;
wire n_504;
wire n_458;
wire n_581;
wire n_418;
wire n_493;
wire n_555;
wire n_698;
wire n_380;
wire n_722;
wire n_618;
wire n_690;
wire n_356;
wire n_281;
wire n_341;
wire n_470;
wire n_600;
wire n_122;
wire n_187;
wire n_375;
wire n_138;
wire n_451;
wire n_487;
wire n_371;
wire n_688;
wire n_323;
wire n_473;
wire n_347;
wire n_558;
wire n_258;
wire n_253;
wire n_515;
wire n_670;
wire n_266;
wire n_683;
wire n_213;
wire n_538;
wire n_182;
wire n_492;
wire n_592;
wire n_368;
wire n_355;
wire n_226;
wire n_382;
wire n_159;
wire n_337;
wire n_658;
wire n_691;
wire n_444;
wire n_176;
wire n_521;
wire n_625;
wire n_650;
wire n_695;
wire n_469;
wire n_585;
wire n_713;
wire n_123;
wire n_457;
wire n_595;
wire n_223;
wire n_494;
wire n_559;
wire n_480;
wire n_372;
wire n_453;
wire n_631;
wire n_194;
wire n_287;
wire n_261;
wire n_110;
wire n_606;
wire n_425;
wire n_332;
wire n_414;
wire n_562;
wire n_350;
wire n_433;
wire n_164;
wire n_421;
wire n_175;
wire n_709;
wire n_145;
wire n_483;
wire n_408;
wire n_290;
wire n_405;
wire n_280;
wire n_99;
wire n_109;
wire n_132;
wire n_406;
wire n_395;
wire n_491;
wire n_151;
wire n_385;
wire n_257;
wire n_269;
INVx1_ASAP7_75t_L g95 ( .A(n_70), .Y(n_95) );
INVx1_ASAP7_75t_L g96 ( .A(n_78), .Y(n_96) );
CKINVDCx5p33_ASAP7_75t_R g97 ( .A(n_42), .Y(n_97) );
INVx1_ASAP7_75t_L g98 ( .A(n_59), .Y(n_98) );
BUFx3_ASAP7_75t_L g99 ( .A(n_51), .Y(n_99) );
CKINVDCx5p33_ASAP7_75t_R g100 ( .A(n_53), .Y(n_100) );
INVx1_ASAP7_75t_L g101 ( .A(n_61), .Y(n_101) );
INVx1_ASAP7_75t_L g102 ( .A(n_88), .Y(n_102) );
INVx1_ASAP7_75t_L g103 ( .A(n_76), .Y(n_103) );
INVx1_ASAP7_75t_L g104 ( .A(n_92), .Y(n_104) );
INVx1_ASAP7_75t_L g105 ( .A(n_94), .Y(n_105) );
INVx1_ASAP7_75t_L g106 ( .A(n_20), .Y(n_106) );
INVx2_ASAP7_75t_L g107 ( .A(n_71), .Y(n_107) );
CKINVDCx5p33_ASAP7_75t_R g108 ( .A(n_89), .Y(n_108) );
INVx2_ASAP7_75t_L g109 ( .A(n_55), .Y(n_109) );
INVx2_ASAP7_75t_L g110 ( .A(n_41), .Y(n_110) );
CKINVDCx5p33_ASAP7_75t_R g111 ( .A(n_85), .Y(n_111) );
INVx1_ASAP7_75t_L g112 ( .A(n_47), .Y(n_112) );
INVx1_ASAP7_75t_L g113 ( .A(n_31), .Y(n_113) );
CKINVDCx5p33_ASAP7_75t_R g114 ( .A(n_23), .Y(n_114) );
INVx1_ASAP7_75t_L g115 ( .A(n_49), .Y(n_115) );
CKINVDCx5p33_ASAP7_75t_R g116 ( .A(n_40), .Y(n_116) );
INVx1_ASAP7_75t_L g117 ( .A(n_33), .Y(n_117) );
INVx1_ASAP7_75t_L g118 ( .A(n_43), .Y(n_118) );
INVx1_ASAP7_75t_L g119 ( .A(n_24), .Y(n_119) );
INVx1_ASAP7_75t_L g120 ( .A(n_3), .Y(n_120) );
INVx1_ASAP7_75t_L g121 ( .A(n_4), .Y(n_121) );
INVx1_ASAP7_75t_L g122 ( .A(n_7), .Y(n_122) );
INVx1_ASAP7_75t_L g123 ( .A(n_37), .Y(n_123) );
INVx1_ASAP7_75t_L g124 ( .A(n_62), .Y(n_124) );
INVx1_ASAP7_75t_L g125 ( .A(n_90), .Y(n_125) );
BUFx2_ASAP7_75t_SL g126 ( .A(n_67), .Y(n_126) );
BUFx3_ASAP7_75t_L g127 ( .A(n_5), .Y(n_127) );
CKINVDCx14_ASAP7_75t_R g128 ( .A(n_0), .Y(n_128) );
CKINVDCx5p33_ASAP7_75t_R g129 ( .A(n_66), .Y(n_129) );
INVx1_ASAP7_75t_L g130 ( .A(n_5), .Y(n_130) );
OR2x2_ASAP7_75t_L g131 ( .A(n_64), .B(n_39), .Y(n_131) );
INVx1_ASAP7_75t_SL g132 ( .A(n_50), .Y(n_132) );
INVx1_ASAP7_75t_L g133 ( .A(n_32), .Y(n_133) );
HB1xp67_ASAP7_75t_L g134 ( .A(n_79), .Y(n_134) );
INVxp67_ASAP7_75t_L g135 ( .A(n_11), .Y(n_135) );
BUFx6f_ASAP7_75t_L g136 ( .A(n_99), .Y(n_136) );
INVxp67_ASAP7_75t_L g137 ( .A(n_134), .Y(n_137) );
OA21x2_ASAP7_75t_L g138 ( .A1(n_95), .A2(n_0), .B(n_1), .Y(n_138) );
INVx3_ASAP7_75t_L g139 ( .A(n_107), .Y(n_139) );
INVx1_ASAP7_75t_L g140 ( .A(n_95), .Y(n_140) );
AOI22xp5_ASAP7_75t_L g141 ( .A1(n_128), .A2(n_120), .B1(n_121), .B2(n_122), .Y(n_141) );
INVx3_ASAP7_75t_L g142 ( .A(n_96), .Y(n_142) );
INVx2_ASAP7_75t_L g143 ( .A(n_107), .Y(n_143) );
INVx3_ASAP7_75t_L g144 ( .A(n_96), .Y(n_144) );
OA21x2_ASAP7_75t_L g145 ( .A1(n_98), .A2(n_1), .B(n_2), .Y(n_145) );
AND2x2_ASAP7_75t_SL g146 ( .A(n_131), .B(n_21), .Y(n_146) );
OAI22xp5_ASAP7_75t_L g147 ( .A1(n_120), .A2(n_2), .B1(n_3), .B2(n_4), .Y(n_147) );
NOR2xp33_ASAP7_75t_L g148 ( .A(n_135), .B(n_6), .Y(n_148) );
NAND2xp5_ASAP7_75t_L g149 ( .A(n_121), .B(n_6), .Y(n_149) );
AND2x2_ASAP7_75t_L g150 ( .A(n_127), .B(n_7), .Y(n_150) );
INVx1_ASAP7_75t_L g151 ( .A(n_98), .Y(n_151) );
BUFx6f_ASAP7_75t_L g152 ( .A(n_99), .Y(n_152) );
BUFx3_ASAP7_75t_L g153 ( .A(n_109), .Y(n_153) );
INVx1_ASAP7_75t_L g154 ( .A(n_101), .Y(n_154) );
INVx1_ASAP7_75t_L g155 ( .A(n_101), .Y(n_155) );
INVx2_ASAP7_75t_L g156 ( .A(n_136), .Y(n_156) );
INVx2_ASAP7_75t_L g157 ( .A(n_136), .Y(n_157) );
BUFx2_ASAP7_75t_L g158 ( .A(n_137), .Y(n_158) );
INVx2_ASAP7_75t_L g159 ( .A(n_136), .Y(n_159) );
NOR2x1p5_ASAP7_75t_L g160 ( .A(n_149), .B(n_127), .Y(n_160) );
NOR2xp33_ASAP7_75t_L g161 ( .A(n_137), .B(n_115), .Y(n_161) );
BUFx3_ASAP7_75t_L g162 ( .A(n_136), .Y(n_162) );
NAND2xp5_ASAP7_75t_SL g163 ( .A(n_141), .B(n_97), .Y(n_163) );
BUFx6f_ASAP7_75t_L g164 ( .A(n_136), .Y(n_164) );
NOR2xp33_ASAP7_75t_L g165 ( .A(n_140), .B(n_117), .Y(n_165) );
INVx2_ASAP7_75t_SL g166 ( .A(n_142), .Y(n_166) );
INVx2_ASAP7_75t_L g167 ( .A(n_136), .Y(n_167) );
INVx1_ASAP7_75t_L g168 ( .A(n_143), .Y(n_168) );
NAND3xp33_ASAP7_75t_L g169 ( .A(n_140), .B(n_133), .C(n_102), .Y(n_169) );
NAND2xp5_ASAP7_75t_L g170 ( .A(n_140), .B(n_100), .Y(n_170) );
XNOR2xp5_ASAP7_75t_L g171 ( .A(n_141), .B(n_146), .Y(n_171) );
NAND2xp5_ASAP7_75t_SL g172 ( .A(n_151), .B(n_108), .Y(n_172) );
AND2x2_ASAP7_75t_L g173 ( .A(n_150), .B(n_122), .Y(n_173) );
INVx3_ASAP7_75t_L g174 ( .A(n_153), .Y(n_174) );
INVx4_ASAP7_75t_L g175 ( .A(n_146), .Y(n_175) );
INVx2_ASAP7_75t_L g176 ( .A(n_136), .Y(n_176) );
NAND2xp5_ASAP7_75t_L g177 ( .A(n_151), .B(n_111), .Y(n_177) );
INVx2_ASAP7_75t_L g178 ( .A(n_136), .Y(n_178) );
INVx2_ASAP7_75t_L g179 ( .A(n_152), .Y(n_179) );
NOR2xp33_ASAP7_75t_L g180 ( .A(n_151), .B(n_118), .Y(n_180) );
BUFx6f_ASAP7_75t_L g181 ( .A(n_152), .Y(n_181) );
INVx1_ASAP7_75t_L g182 ( .A(n_143), .Y(n_182) );
INVx1_ASAP7_75t_L g183 ( .A(n_143), .Y(n_183) );
INVx2_ASAP7_75t_L g184 ( .A(n_152), .Y(n_184) );
NAND2xp5_ASAP7_75t_L g185 ( .A(n_154), .B(n_114), .Y(n_185) );
OR2x2_ASAP7_75t_SL g186 ( .A(n_171), .B(n_138), .Y(n_186) );
INVx1_ASAP7_75t_L g187 ( .A(n_168), .Y(n_187) );
NAND2xp5_ASAP7_75t_SL g188 ( .A(n_158), .B(n_146), .Y(n_188) );
AND2x2_ASAP7_75t_L g189 ( .A(n_158), .B(n_146), .Y(n_189) );
NOR2xp33_ASAP7_75t_L g190 ( .A(n_173), .B(n_148), .Y(n_190) );
INVx2_ASAP7_75t_L g191 ( .A(n_162), .Y(n_191) );
AOI22xp33_ASAP7_75t_L g192 ( .A1(n_175), .A2(n_150), .B1(n_145), .B2(n_138), .Y(n_192) );
NOR2xp33_ASAP7_75t_R g193 ( .A(n_171), .B(n_150), .Y(n_193) );
INVx2_ASAP7_75t_L g194 ( .A(n_162), .Y(n_194) );
INVx1_ASAP7_75t_L g195 ( .A(n_168), .Y(n_195) );
NAND2x1_ASAP7_75t_L g196 ( .A(n_175), .B(n_142), .Y(n_196) );
NAND2xp5_ASAP7_75t_L g197 ( .A(n_173), .B(n_154), .Y(n_197) );
INVxp67_ASAP7_75t_L g198 ( .A(n_161), .Y(n_198) );
INVx1_ASAP7_75t_L g199 ( .A(n_182), .Y(n_199) );
NOR2xp33_ASAP7_75t_SL g200 ( .A(n_175), .B(n_147), .Y(n_200) );
INVx1_ASAP7_75t_L g201 ( .A(n_182), .Y(n_201) );
NAND2xp5_ASAP7_75t_L g202 ( .A(n_170), .B(n_154), .Y(n_202) );
INVx2_ASAP7_75t_L g203 ( .A(n_162), .Y(n_203) );
INVx2_ASAP7_75t_L g204 ( .A(n_166), .Y(n_204) );
AND2x6_ASAP7_75t_SL g205 ( .A(n_165), .B(n_148), .Y(n_205) );
A2O1A1Ixp33_ASAP7_75t_L g206 ( .A1(n_180), .A2(n_142), .B(n_144), .C(n_155), .Y(n_206) );
NAND2xp5_ASAP7_75t_L g207 ( .A(n_177), .B(n_155), .Y(n_207) );
INVx2_ASAP7_75t_SL g208 ( .A(n_160), .Y(n_208) );
OAI22xp5_ASAP7_75t_L g209 ( .A1(n_175), .A2(n_149), .B1(n_155), .B2(n_147), .Y(n_209) );
CKINVDCx5p33_ASAP7_75t_R g210 ( .A(n_163), .Y(n_210) );
NOR2xp33_ASAP7_75t_L g211 ( .A(n_172), .B(n_142), .Y(n_211) );
NAND2xp5_ASAP7_75t_SL g212 ( .A(n_185), .B(n_116), .Y(n_212) );
AOI22xp5_ASAP7_75t_L g213 ( .A1(n_160), .A2(n_169), .B1(n_174), .B2(n_144), .Y(n_213) );
INVx2_ASAP7_75t_L g214 ( .A(n_166), .Y(n_214) );
BUFx3_ASAP7_75t_L g215 ( .A(n_174), .Y(n_215) );
AND2x2_ASAP7_75t_L g216 ( .A(n_183), .B(n_142), .Y(n_216) );
INVx1_ASAP7_75t_L g217 ( .A(n_183), .Y(n_217) );
NAND2x1p5_ASAP7_75t_L g218 ( .A(n_174), .B(n_138), .Y(n_218) );
NAND2xp5_ASAP7_75t_L g219 ( .A(n_174), .B(n_144), .Y(n_219) );
CKINVDCx5p33_ASAP7_75t_R g220 ( .A(n_169), .Y(n_220) );
INVx2_ASAP7_75t_L g221 ( .A(n_157), .Y(n_221) );
NAND2xp5_ASAP7_75t_L g222 ( .A(n_156), .B(n_144), .Y(n_222) );
NOR2xp33_ASAP7_75t_L g223 ( .A(n_164), .B(n_144), .Y(n_223) );
NAND2xp5_ASAP7_75t_L g224 ( .A(n_156), .B(n_153), .Y(n_224) );
AOI22xp33_ASAP7_75t_L g225 ( .A1(n_159), .A2(n_138), .B1(n_145), .B2(n_153), .Y(n_225) );
NOR2xp33_ASAP7_75t_L g226 ( .A(n_198), .B(n_130), .Y(n_226) );
OR2x2_ASAP7_75t_L g227 ( .A(n_209), .B(n_189), .Y(n_227) );
INVx1_ASAP7_75t_L g228 ( .A(n_216), .Y(n_228) );
OAI22xp5_ASAP7_75t_L g229 ( .A1(n_188), .A2(n_153), .B1(n_138), .B2(n_145), .Y(n_229) );
NOR3xp33_ASAP7_75t_L g230 ( .A(n_189), .B(n_125), .C(n_103), .Y(n_230) );
O2A1O1Ixp33_ASAP7_75t_L g231 ( .A1(n_206), .A2(n_143), .B(n_139), .C(n_104), .Y(n_231) );
INVx1_ASAP7_75t_L g232 ( .A(n_216), .Y(n_232) );
OR2x2_ASAP7_75t_L g233 ( .A(n_197), .B(n_138), .Y(n_233) );
NAND2xp5_ASAP7_75t_L g234 ( .A(n_190), .B(n_145), .Y(n_234) );
OAI21xp5_ASAP7_75t_L g235 ( .A1(n_192), .A2(n_179), .B(n_178), .Y(n_235) );
INVx2_ASAP7_75t_L g236 ( .A(n_187), .Y(n_236) );
BUFx4f_ASAP7_75t_L g237 ( .A(n_208), .Y(n_237) );
NAND2xp5_ASAP7_75t_SL g238 ( .A(n_220), .B(n_129), .Y(n_238) );
OA22x2_ASAP7_75t_L g239 ( .A1(n_210), .A2(n_126), .B1(n_102), .B2(n_112), .Y(n_239) );
INVx1_ASAP7_75t_L g240 ( .A(n_187), .Y(n_240) );
AOI21xp5_ASAP7_75t_L g241 ( .A1(n_202), .A2(n_159), .B(n_176), .Y(n_241) );
INVx1_ASAP7_75t_L g242 ( .A(n_195), .Y(n_242) );
NOR2xp33_ASAP7_75t_L g243 ( .A(n_208), .B(n_132), .Y(n_243) );
INVx2_ASAP7_75t_L g244 ( .A(n_195), .Y(n_244) );
INVx3_ASAP7_75t_L g245 ( .A(n_215), .Y(n_245) );
NAND2xp5_ASAP7_75t_L g246 ( .A(n_207), .B(n_145), .Y(n_246) );
INVx3_ASAP7_75t_L g247 ( .A(n_215), .Y(n_247) );
INVx3_ASAP7_75t_L g248 ( .A(n_215), .Y(n_248) );
OAI21xp33_ASAP7_75t_L g249 ( .A1(n_200), .A2(n_139), .B(n_104), .Y(n_249) );
BUFx6f_ASAP7_75t_L g250 ( .A(n_196), .Y(n_250) );
O2A1O1Ixp33_ASAP7_75t_L g251 ( .A1(n_199), .A2(n_139), .B(n_105), .C(n_106), .Y(n_251) );
HB1xp67_ASAP7_75t_L g252 ( .A(n_199), .Y(n_252) );
OAI22xp5_ASAP7_75t_L g253 ( .A1(n_186), .A2(n_145), .B1(n_131), .B2(n_139), .Y(n_253) );
CKINVDCx6p67_ASAP7_75t_R g254 ( .A(n_212), .Y(n_254) );
OR2x6_ASAP7_75t_SL g255 ( .A(n_193), .B(n_103), .Y(n_255) );
AOI21xp5_ASAP7_75t_L g256 ( .A1(n_196), .A2(n_176), .B(n_178), .Y(n_256) );
NAND2xp5_ASAP7_75t_SL g257 ( .A(n_201), .B(n_152), .Y(n_257) );
NAND2xp5_ASAP7_75t_SL g258 ( .A(n_201), .B(n_152), .Y(n_258) );
NOR2xp33_ASAP7_75t_L g259 ( .A(n_205), .B(n_139), .Y(n_259) );
BUFx3_ASAP7_75t_L g260 ( .A(n_250), .Y(n_260) );
AOI21xp5_ASAP7_75t_L g261 ( .A1(n_234), .A2(n_219), .B(n_204), .Y(n_261) );
AOI21xp5_ASAP7_75t_L g262 ( .A1(n_246), .A2(n_204), .B(n_214), .Y(n_262) );
BUFx2_ASAP7_75t_L g263 ( .A(n_255), .Y(n_263) );
AOI22xp33_ASAP7_75t_L g264 ( .A1(n_230), .A2(n_211), .B1(n_217), .B2(n_213), .Y(n_264) );
AOI21xp5_ASAP7_75t_L g265 ( .A1(n_241), .A2(n_204), .B(n_214), .Y(n_265) );
AND2x4_ASAP7_75t_L g266 ( .A(n_228), .B(n_217), .Y(n_266) );
AOI21xp5_ASAP7_75t_L g267 ( .A1(n_235), .A2(n_214), .B(n_203), .Y(n_267) );
AO31x2_ASAP7_75t_L g268 ( .A1(n_253), .A2(n_223), .A3(n_157), .B(n_167), .Y(n_268) );
AOI221xp5_ASAP7_75t_L g269 ( .A1(n_226), .A2(n_213), .B1(n_225), .B2(n_139), .C(n_205), .Y(n_269) );
INVx1_ASAP7_75t_L g270 ( .A(n_240), .Y(n_270) );
AOI21xp5_ASAP7_75t_SL g271 ( .A1(n_252), .A2(n_218), .B(n_106), .Y(n_271) );
OAI21x1_ASAP7_75t_L g272 ( .A1(n_229), .A2(n_218), .B(n_167), .Y(n_272) );
OAI21x1_ASAP7_75t_L g273 ( .A1(n_257), .A2(n_218), .B(n_167), .Y(n_273) );
AND2x2_ASAP7_75t_L g274 ( .A(n_252), .B(n_191), .Y(n_274) );
AOI211x1_ASAP7_75t_L g275 ( .A1(n_232), .A2(n_224), .B(n_123), .C(n_119), .Y(n_275) );
BUFx2_ASAP7_75t_L g276 ( .A(n_236), .Y(n_276) );
AOI21xp5_ASAP7_75t_L g277 ( .A1(n_256), .A2(n_203), .B(n_194), .Y(n_277) );
INVx1_ASAP7_75t_L g278 ( .A(n_242), .Y(n_278) );
OAI21x1_ASAP7_75t_L g279 ( .A1(n_257), .A2(n_184), .B(n_157), .Y(n_279) );
INVx1_ASAP7_75t_L g280 ( .A(n_244), .Y(n_280) );
OAI21x1_ASAP7_75t_L g281 ( .A1(n_258), .A2(n_184), .B(n_221), .Y(n_281) );
AO31x2_ASAP7_75t_L g282 ( .A1(n_259), .A2(n_184), .A3(n_179), .B(n_119), .Y(n_282) );
OAI21x1_ASAP7_75t_L g283 ( .A1(n_258), .A2(n_221), .B(n_222), .Y(n_283) );
AND2x2_ASAP7_75t_L g284 ( .A(n_266), .B(n_227), .Y(n_284) );
INVx1_ASAP7_75t_L g285 ( .A(n_270), .Y(n_285) );
AO31x2_ASAP7_75t_L g286 ( .A1(n_267), .A2(n_259), .A3(n_226), .B(n_105), .Y(n_286) );
NAND2x1p5_ASAP7_75t_L g287 ( .A(n_260), .B(n_245), .Y(n_287) );
NOR2xp33_ASAP7_75t_L g288 ( .A(n_263), .B(n_254), .Y(n_288) );
INVx1_ASAP7_75t_L g289 ( .A(n_278), .Y(n_289) );
A2O1A1Ixp33_ASAP7_75t_L g290 ( .A1(n_269), .A2(n_231), .B(n_249), .C(n_251), .Y(n_290) );
NOR2xp33_ASAP7_75t_L g291 ( .A(n_266), .B(n_243), .Y(n_291) );
AND2x2_ASAP7_75t_L g292 ( .A(n_266), .B(n_230), .Y(n_292) );
CKINVDCx20_ASAP7_75t_R g293 ( .A(n_276), .Y(n_293) );
AOI22xp33_ASAP7_75t_L g294 ( .A1(n_276), .A2(n_239), .B1(n_243), .B2(n_238), .Y(n_294) );
HB1xp67_ASAP7_75t_L g295 ( .A(n_280), .Y(n_295) );
AND2x2_ASAP7_75t_L g296 ( .A(n_274), .B(n_233), .Y(n_296) );
NOR2xp33_ASAP7_75t_L g297 ( .A(n_260), .B(n_237), .Y(n_297) );
INVx1_ASAP7_75t_L g298 ( .A(n_274), .Y(n_298) );
AOI21xp5_ASAP7_75t_L g299 ( .A1(n_271), .A2(n_194), .B(n_203), .Y(n_299) );
INVx1_ASAP7_75t_L g300 ( .A(n_275), .Y(n_300) );
AOI21xp5_ASAP7_75t_L g301 ( .A1(n_271), .A2(n_194), .B(n_191), .Y(n_301) );
INVx1_ASAP7_75t_L g302 ( .A(n_282), .Y(n_302) );
INVx3_ASAP7_75t_L g303 ( .A(n_282), .Y(n_303) );
AO31x2_ASAP7_75t_L g304 ( .A1(n_261), .A2(n_133), .A3(n_124), .B(n_112), .Y(n_304) );
OA21x2_ASAP7_75t_L g305 ( .A1(n_272), .A2(n_281), .B(n_283), .Y(n_305) );
OR2x2_ASAP7_75t_L g306 ( .A(n_284), .B(n_268), .Y(n_306) );
INVx1_ASAP7_75t_L g307 ( .A(n_302), .Y(n_307) );
AND2x2_ASAP7_75t_L g308 ( .A(n_284), .B(n_282), .Y(n_308) );
AND2x2_ASAP7_75t_L g309 ( .A(n_296), .B(n_282), .Y(n_309) );
INVx1_ASAP7_75t_L g310 ( .A(n_302), .Y(n_310) );
AND2x2_ASAP7_75t_L g311 ( .A(n_296), .B(n_282), .Y(n_311) );
AND2x2_ASAP7_75t_L g312 ( .A(n_292), .B(n_268), .Y(n_312) );
BUFx3_ASAP7_75t_L g313 ( .A(n_293), .Y(n_313) );
OAI31xp33_ASAP7_75t_SL g314 ( .A1(n_292), .A2(n_272), .A3(n_113), .B(n_123), .Y(n_314) );
OR2x6_ASAP7_75t_L g315 ( .A(n_303), .B(n_273), .Y(n_315) );
INVx2_ASAP7_75t_L g316 ( .A(n_305), .Y(n_316) );
NAND2xp5_ASAP7_75t_L g317 ( .A(n_298), .B(n_268), .Y(n_317) );
AND2x4_ASAP7_75t_L g318 ( .A(n_298), .B(n_268), .Y(n_318) );
INVx1_ASAP7_75t_L g319 ( .A(n_285), .Y(n_319) );
INVx1_ASAP7_75t_L g320 ( .A(n_285), .Y(n_320) );
HB1xp67_ASAP7_75t_L g321 ( .A(n_303), .Y(n_321) );
HB1xp67_ASAP7_75t_L g322 ( .A(n_303), .Y(n_322) );
INVx1_ASAP7_75t_L g323 ( .A(n_289), .Y(n_323) );
AND2x2_ASAP7_75t_L g324 ( .A(n_300), .B(n_268), .Y(n_324) );
AND2x2_ASAP7_75t_L g325 ( .A(n_300), .B(n_264), .Y(n_325) );
INVx2_ASAP7_75t_L g326 ( .A(n_305), .Y(n_326) );
OR2x6_ASAP7_75t_L g327 ( .A(n_287), .B(n_273), .Y(n_327) );
AO21x2_ASAP7_75t_L g328 ( .A1(n_299), .A2(n_262), .B(n_265), .Y(n_328) );
AO21x2_ASAP7_75t_L g329 ( .A1(n_301), .A2(n_283), .B(n_281), .Y(n_329) );
AO21x2_ASAP7_75t_L g330 ( .A1(n_290), .A2(n_277), .B(n_279), .Y(n_330) );
INVx1_ASAP7_75t_L g331 ( .A(n_289), .Y(n_331) );
INVx1_ASAP7_75t_L g332 ( .A(n_304), .Y(n_332) );
INVx1_ASAP7_75t_L g333 ( .A(n_304), .Y(n_333) );
NOR2xp33_ASAP7_75t_L g334 ( .A(n_288), .B(n_237), .Y(n_334) );
HB1xp67_ASAP7_75t_L g335 ( .A(n_295), .Y(n_335) );
INVx1_ASAP7_75t_L g336 ( .A(n_304), .Y(n_336) );
AOI22xp33_ASAP7_75t_L g337 ( .A1(n_312), .A2(n_291), .B1(n_239), .B2(n_294), .Y(n_337) );
BUFx2_ASAP7_75t_L g338 ( .A(n_327), .Y(n_338) );
AND2x2_ASAP7_75t_L g339 ( .A(n_312), .B(n_286), .Y(n_339) );
INVx2_ASAP7_75t_L g340 ( .A(n_316), .Y(n_340) );
NOR2x1p5_ASAP7_75t_L g341 ( .A(n_332), .B(n_286), .Y(n_341) );
INVx1_ASAP7_75t_L g342 ( .A(n_307), .Y(n_342) );
AND2x2_ASAP7_75t_L g343 ( .A(n_318), .B(n_286), .Y(n_343) );
HB1xp67_ASAP7_75t_L g344 ( .A(n_321), .Y(n_344) );
INVx1_ASAP7_75t_L g345 ( .A(n_307), .Y(n_345) );
INVx1_ASAP7_75t_L g346 ( .A(n_310), .Y(n_346) );
BUFx3_ASAP7_75t_L g347 ( .A(n_327), .Y(n_347) );
AND2x2_ASAP7_75t_L g348 ( .A(n_318), .B(n_286), .Y(n_348) );
AND2x2_ASAP7_75t_L g349 ( .A(n_318), .B(n_286), .Y(n_349) );
INVx2_ASAP7_75t_L g350 ( .A(n_316), .Y(n_350) );
INVx2_ASAP7_75t_L g351 ( .A(n_316), .Y(n_351) );
HB1xp67_ASAP7_75t_L g352 ( .A(n_321), .Y(n_352) );
AND2x2_ASAP7_75t_SL g353 ( .A(n_314), .B(n_305), .Y(n_353) );
HB1xp67_ASAP7_75t_L g354 ( .A(n_322), .Y(n_354) );
INVxp67_ASAP7_75t_L g355 ( .A(n_335), .Y(n_355) );
NAND2xp5_ASAP7_75t_L g356 ( .A(n_319), .B(n_304), .Y(n_356) );
BUFx6f_ASAP7_75t_L g357 ( .A(n_327), .Y(n_357) );
AND2x2_ASAP7_75t_L g358 ( .A(n_318), .B(n_304), .Y(n_358) );
HB1xp67_ASAP7_75t_L g359 ( .A(n_322), .Y(n_359) );
OR2x2_ASAP7_75t_L g360 ( .A(n_306), .B(n_305), .Y(n_360) );
AND2x2_ASAP7_75t_L g361 ( .A(n_308), .B(n_113), .Y(n_361) );
HB1xp67_ASAP7_75t_L g362 ( .A(n_335), .Y(n_362) );
INVx3_ASAP7_75t_L g363 ( .A(n_327), .Y(n_363) );
INVx1_ASAP7_75t_L g364 ( .A(n_310), .Y(n_364) );
INVx2_ASAP7_75t_L g365 ( .A(n_326), .Y(n_365) );
INVx2_ASAP7_75t_L g366 ( .A(n_326), .Y(n_366) );
NAND2xp5_ASAP7_75t_L g367 ( .A(n_319), .B(n_287), .Y(n_367) );
OR2x2_ASAP7_75t_SL g368 ( .A(n_306), .B(n_124), .Y(n_368) );
AND2x2_ASAP7_75t_L g369 ( .A(n_308), .B(n_287), .Y(n_369) );
INVx2_ASAP7_75t_L g370 ( .A(n_326), .Y(n_370) );
BUFx2_ASAP7_75t_L g371 ( .A(n_327), .Y(n_371) );
INVxp67_ASAP7_75t_SL g372 ( .A(n_336), .Y(n_372) );
INVx2_ASAP7_75t_L g373 ( .A(n_315), .Y(n_373) );
AND2x4_ASAP7_75t_L g374 ( .A(n_315), .B(n_279), .Y(n_374) );
INVxp67_ASAP7_75t_SL g375 ( .A(n_336), .Y(n_375) );
AND2x2_ASAP7_75t_L g376 ( .A(n_309), .B(n_126), .Y(n_376) );
INVx2_ASAP7_75t_SL g377 ( .A(n_327), .Y(n_377) );
INVxp67_ASAP7_75t_SL g378 ( .A(n_332), .Y(n_378) );
AND2x6_ASAP7_75t_L g379 ( .A(n_309), .B(n_297), .Y(n_379) );
OAI33xp33_ASAP7_75t_L g380 ( .A1(n_320), .A2(n_109), .A3(n_110), .B1(n_10), .B2(n_11), .B3(n_12), .Y(n_380) );
BUFx2_ASAP7_75t_L g381 ( .A(n_315), .Y(n_381) );
INVx1_ASAP7_75t_L g382 ( .A(n_333), .Y(n_382) );
INVx2_ASAP7_75t_L g383 ( .A(n_315), .Y(n_383) );
INVx2_ASAP7_75t_L g384 ( .A(n_315), .Y(n_384) );
INVx1_ASAP7_75t_L g385 ( .A(n_333), .Y(n_385) );
AND2x2_ASAP7_75t_L g386 ( .A(n_311), .B(n_110), .Y(n_386) );
NAND2xp5_ASAP7_75t_L g387 ( .A(n_320), .B(n_250), .Y(n_387) );
BUFx6f_ASAP7_75t_L g388 ( .A(n_315), .Y(n_388) );
HB1xp67_ASAP7_75t_L g389 ( .A(n_317), .Y(n_389) );
INVx2_ASAP7_75t_L g390 ( .A(n_340), .Y(n_390) );
AND2x2_ASAP7_75t_L g391 ( .A(n_343), .B(n_324), .Y(n_391) );
AND2x2_ASAP7_75t_L g392 ( .A(n_343), .B(n_324), .Y(n_392) );
OR2x2_ASAP7_75t_L g393 ( .A(n_389), .B(n_317), .Y(n_393) );
OR2x2_ASAP7_75t_L g394 ( .A(n_389), .B(n_311), .Y(n_394) );
AND2x2_ASAP7_75t_L g395 ( .A(n_348), .B(n_323), .Y(n_395) );
AND2x4_ASAP7_75t_L g396 ( .A(n_377), .B(n_323), .Y(n_396) );
NAND2xp5_ASAP7_75t_L g397 ( .A(n_361), .B(n_331), .Y(n_397) );
AND2x2_ASAP7_75t_L g398 ( .A(n_348), .B(n_331), .Y(n_398) );
NAND2xp5_ASAP7_75t_L g399 ( .A(n_361), .B(n_325), .Y(n_399) );
INVx1_ASAP7_75t_L g400 ( .A(n_362), .Y(n_400) );
INVx1_ASAP7_75t_SL g401 ( .A(n_362), .Y(n_401) );
NOR2xp33_ASAP7_75t_L g402 ( .A(n_355), .B(n_313), .Y(n_402) );
AND2x2_ASAP7_75t_L g403 ( .A(n_349), .B(n_325), .Y(n_403) );
NAND2xp5_ASAP7_75t_L g404 ( .A(n_386), .B(n_314), .Y(n_404) );
INVx1_ASAP7_75t_L g405 ( .A(n_355), .Y(n_405) );
OR2x2_ASAP7_75t_L g406 ( .A(n_360), .B(n_313), .Y(n_406) );
INVx2_ASAP7_75t_L g407 ( .A(n_340), .Y(n_407) );
AND2x2_ASAP7_75t_L g408 ( .A(n_349), .B(n_329), .Y(n_408) );
INVx2_ASAP7_75t_L g409 ( .A(n_340), .Y(n_409) );
AND2x2_ASAP7_75t_L g410 ( .A(n_358), .B(n_329), .Y(n_410) );
INVx1_ASAP7_75t_L g411 ( .A(n_342), .Y(n_411) );
INVx1_ASAP7_75t_L g412 ( .A(n_345), .Y(n_412) );
INVx1_ASAP7_75t_L g413 ( .A(n_345), .Y(n_413) );
INVx1_ASAP7_75t_L g414 ( .A(n_346), .Y(n_414) );
BUFx2_ASAP7_75t_L g415 ( .A(n_344), .Y(n_415) );
AND2x2_ASAP7_75t_L g416 ( .A(n_358), .B(n_329), .Y(n_416) );
INVx1_ASAP7_75t_L g417 ( .A(n_346), .Y(n_417) );
AND2x2_ASAP7_75t_L g418 ( .A(n_339), .B(n_329), .Y(n_418) );
OR2x2_ASAP7_75t_L g419 ( .A(n_360), .B(n_313), .Y(n_419) );
INVx2_ASAP7_75t_L g420 ( .A(n_350), .Y(n_420) );
OR2x2_ASAP7_75t_L g421 ( .A(n_344), .B(n_330), .Y(n_421) );
NAND2xp5_ASAP7_75t_L g422 ( .A(n_386), .B(n_330), .Y(n_422) );
INVx1_ASAP7_75t_L g423 ( .A(n_364), .Y(n_423) );
BUFx2_ASAP7_75t_L g424 ( .A(n_352), .Y(n_424) );
NAND2xp5_ASAP7_75t_L g425 ( .A(n_376), .B(n_330), .Y(n_425) );
INVx1_ASAP7_75t_L g426 ( .A(n_364), .Y(n_426) );
NAND2xp5_ASAP7_75t_L g427 ( .A(n_376), .B(n_330), .Y(n_427) );
NAND2xp5_ASAP7_75t_L g428 ( .A(n_339), .B(n_334), .Y(n_428) );
INVx1_ASAP7_75t_L g429 ( .A(n_387), .Y(n_429) );
INVx2_ASAP7_75t_L g430 ( .A(n_350), .Y(n_430) );
INVx1_ASAP7_75t_L g431 ( .A(n_387), .Y(n_431) );
INVx1_ASAP7_75t_SL g432 ( .A(n_369), .Y(n_432) );
INVx1_ASAP7_75t_L g433 ( .A(n_382), .Y(n_433) );
AND2x2_ASAP7_75t_L g434 ( .A(n_341), .B(n_328), .Y(n_434) );
INVx1_ASAP7_75t_L g435 ( .A(n_382), .Y(n_435) );
HB1xp67_ASAP7_75t_L g436 ( .A(n_352), .Y(n_436) );
INVx2_ASAP7_75t_L g437 ( .A(n_350), .Y(n_437) );
AND2x4_ASAP7_75t_L g438 ( .A(n_377), .B(n_328), .Y(n_438) );
INVx1_ASAP7_75t_L g439 ( .A(n_385), .Y(n_439) );
INVx1_ASAP7_75t_L g440 ( .A(n_385), .Y(n_440) );
INVx2_ASAP7_75t_L g441 ( .A(n_351), .Y(n_441) );
NOR2xp67_ASAP7_75t_L g442 ( .A(n_363), .B(n_8), .Y(n_442) );
INVx4_ASAP7_75t_L g443 ( .A(n_379), .Y(n_443) );
INVx1_ASAP7_75t_L g444 ( .A(n_367), .Y(n_444) );
INVx1_ASAP7_75t_L g445 ( .A(n_367), .Y(n_445) );
INVx2_ASAP7_75t_L g446 ( .A(n_351), .Y(n_446) );
INVx1_ASAP7_75t_L g447 ( .A(n_372), .Y(n_447) );
INVx1_ASAP7_75t_L g448 ( .A(n_372), .Y(n_448) );
OAI322xp33_ASAP7_75t_L g449 ( .A1(n_356), .A2(n_152), .A3(n_9), .B1(n_10), .B2(n_12), .C1(n_13), .C2(n_14), .Y(n_449) );
AND2x4_ASAP7_75t_L g450 ( .A(n_377), .B(n_363), .Y(n_450) );
AND2x2_ASAP7_75t_L g451 ( .A(n_341), .B(n_328), .Y(n_451) );
INVx2_ASAP7_75t_L g452 ( .A(n_351), .Y(n_452) );
AND2x4_ASAP7_75t_L g453 ( .A(n_363), .B(n_328), .Y(n_453) );
AND2x4_ASAP7_75t_L g454 ( .A(n_363), .B(n_152), .Y(n_454) );
AND2x2_ASAP7_75t_L g455 ( .A(n_369), .B(n_152), .Y(n_455) );
AND2x2_ASAP7_75t_L g456 ( .A(n_365), .B(n_8), .Y(n_456) );
AND2x2_ASAP7_75t_L g457 ( .A(n_365), .B(n_9), .Y(n_457) );
NAND2xp5_ASAP7_75t_L g458 ( .A(n_337), .B(n_13), .Y(n_458) );
NAND2xp5_ASAP7_75t_L g459 ( .A(n_356), .B(n_14), .Y(n_459) );
AND2x2_ASAP7_75t_L g460 ( .A(n_365), .B(n_15), .Y(n_460) );
BUFx2_ASAP7_75t_L g461 ( .A(n_354), .Y(n_461) );
INVx2_ASAP7_75t_L g462 ( .A(n_366), .Y(n_462) );
OR2x2_ASAP7_75t_L g463 ( .A(n_354), .B(n_186), .Y(n_463) );
AND2x2_ASAP7_75t_L g464 ( .A(n_366), .B(n_15), .Y(n_464) );
AND2x4_ASAP7_75t_SL g465 ( .A(n_357), .B(n_250), .Y(n_465) );
HB1xp67_ASAP7_75t_L g466 ( .A(n_359), .Y(n_466) );
AND2x2_ASAP7_75t_L g467 ( .A(n_366), .B(n_370), .Y(n_467) );
OR2x2_ASAP7_75t_L g468 ( .A(n_394), .B(n_359), .Y(n_468) );
AND2x2_ASAP7_75t_L g469 ( .A(n_432), .B(n_381), .Y(n_469) );
INVx1_ASAP7_75t_L g470 ( .A(n_405), .Y(n_470) );
AND2x2_ASAP7_75t_L g471 ( .A(n_391), .B(n_381), .Y(n_471) );
OR2x2_ASAP7_75t_L g472 ( .A(n_394), .B(n_375), .Y(n_472) );
NAND2xp5_ASAP7_75t_L g473 ( .A(n_403), .B(n_375), .Y(n_473) );
INVx2_ASAP7_75t_L g474 ( .A(n_467), .Y(n_474) );
AND2x2_ASAP7_75t_L g475 ( .A(n_391), .B(n_338), .Y(n_475) );
OR2x2_ASAP7_75t_L g476 ( .A(n_406), .B(n_378), .Y(n_476) );
INVx1_ASAP7_75t_L g477 ( .A(n_413), .Y(n_477) );
AND2x4_ASAP7_75t_L g478 ( .A(n_443), .B(n_338), .Y(n_478) );
HB1xp67_ASAP7_75t_L g479 ( .A(n_401), .Y(n_479) );
INVx1_ASAP7_75t_L g480 ( .A(n_413), .Y(n_480) );
HB1xp67_ASAP7_75t_L g481 ( .A(n_415), .Y(n_481) );
OR2x2_ASAP7_75t_L g482 ( .A(n_406), .B(n_378), .Y(n_482) );
OR2x2_ASAP7_75t_L g483 ( .A(n_419), .B(n_370), .Y(n_483) );
INVx1_ASAP7_75t_L g484 ( .A(n_414), .Y(n_484) );
NAND2xp5_ASAP7_75t_L g485 ( .A(n_403), .B(n_379), .Y(n_485) );
NAND2xp5_ASAP7_75t_L g486 ( .A(n_395), .B(n_379), .Y(n_486) );
AND2x2_ASAP7_75t_L g487 ( .A(n_392), .B(n_371), .Y(n_487) );
NAND2xp5_ASAP7_75t_L g488 ( .A(n_418), .B(n_370), .Y(n_488) );
AND2x2_ASAP7_75t_L g489 ( .A(n_395), .B(n_373), .Y(n_489) );
NAND2xp5_ASAP7_75t_L g490 ( .A(n_418), .B(n_353), .Y(n_490) );
INVx1_ASAP7_75t_L g491 ( .A(n_414), .Y(n_491) );
OR2x2_ASAP7_75t_L g492 ( .A(n_419), .B(n_368), .Y(n_492) );
AND2x2_ASAP7_75t_L g493 ( .A(n_398), .B(n_373), .Y(n_493) );
INVx2_ASAP7_75t_L g494 ( .A(n_467), .Y(n_494) );
NAND2xp5_ASAP7_75t_L g495 ( .A(n_429), .B(n_353), .Y(n_495) );
INVx1_ASAP7_75t_L g496 ( .A(n_417), .Y(n_496) );
AND2x2_ASAP7_75t_L g497 ( .A(n_398), .B(n_373), .Y(n_497) );
INVx1_ASAP7_75t_SL g498 ( .A(n_415), .Y(n_498) );
INVx1_ASAP7_75t_L g499 ( .A(n_417), .Y(n_499) );
INVx4_ASAP7_75t_L g500 ( .A(n_443), .Y(n_500) );
NAND2xp5_ASAP7_75t_L g501 ( .A(n_431), .B(n_353), .Y(n_501) );
AND2x2_ASAP7_75t_L g502 ( .A(n_402), .B(n_383), .Y(n_502) );
OR2x6_ASAP7_75t_L g503 ( .A(n_443), .B(n_347), .Y(n_503) );
INVx1_ASAP7_75t_L g504 ( .A(n_400), .Y(n_504) );
INVx1_ASAP7_75t_L g505 ( .A(n_411), .Y(n_505) );
AND2x4_ASAP7_75t_L g506 ( .A(n_450), .B(n_347), .Y(n_506) );
NAND2xp5_ASAP7_75t_L g507 ( .A(n_393), .B(n_383), .Y(n_507) );
AND2x2_ASAP7_75t_L g508 ( .A(n_455), .B(n_383), .Y(n_508) );
NAND2xp5_ASAP7_75t_L g509 ( .A(n_444), .B(n_379), .Y(n_509) );
OR2x2_ASAP7_75t_L g510 ( .A(n_393), .B(n_368), .Y(n_510) );
NAND2xp5_ASAP7_75t_SL g511 ( .A(n_442), .B(n_357), .Y(n_511) );
OR2x2_ASAP7_75t_L g512 ( .A(n_436), .B(n_347), .Y(n_512) );
INVx2_ASAP7_75t_L g513 ( .A(n_424), .Y(n_513) );
INVx2_ASAP7_75t_SL g514 ( .A(n_455), .Y(n_514) );
NAND2xp5_ASAP7_75t_L g515 ( .A(n_445), .B(n_384), .Y(n_515) );
INVx2_ASAP7_75t_L g516 ( .A(n_424), .Y(n_516) );
INVx1_ASAP7_75t_L g517 ( .A(n_412), .Y(n_517) );
INVx3_ASAP7_75t_L g518 ( .A(n_396), .Y(n_518) );
INVx1_ASAP7_75t_SL g519 ( .A(n_461), .Y(n_519) );
INVx2_ASAP7_75t_L g520 ( .A(n_461), .Y(n_520) );
INVx1_ASAP7_75t_L g521 ( .A(n_423), .Y(n_521) );
INVx2_ASAP7_75t_L g522 ( .A(n_390), .Y(n_522) );
OAI31xp33_ASAP7_75t_L g523 ( .A1(n_404), .A2(n_374), .A3(n_384), .B(n_379), .Y(n_523) );
INVx1_ASAP7_75t_L g524 ( .A(n_426), .Y(n_524) );
AND2x2_ASAP7_75t_L g525 ( .A(n_408), .B(n_384), .Y(n_525) );
AND2x2_ASAP7_75t_L g526 ( .A(n_408), .B(n_379), .Y(n_526) );
OR2x6_ASAP7_75t_L g527 ( .A(n_396), .B(n_357), .Y(n_527) );
INVx1_ASAP7_75t_L g528 ( .A(n_433), .Y(n_528) );
AND2x2_ASAP7_75t_L g529 ( .A(n_428), .B(n_379), .Y(n_529) );
NAND2xp67_ASAP7_75t_L g530 ( .A(n_434), .B(n_379), .Y(n_530) );
AND2x2_ASAP7_75t_L g531 ( .A(n_410), .B(n_388), .Y(n_531) );
NAND2xp5_ASAP7_75t_L g532 ( .A(n_435), .B(n_388), .Y(n_532) );
OR2x2_ASAP7_75t_L g533 ( .A(n_466), .B(n_357), .Y(n_533) );
NAND2xp5_ASAP7_75t_L g534 ( .A(n_439), .B(n_388), .Y(n_534) );
NAND2xp5_ASAP7_75t_L g535 ( .A(n_397), .B(n_388), .Y(n_535) );
INVx1_ASAP7_75t_L g536 ( .A(n_440), .Y(n_536) );
INVx1_ASAP7_75t_L g537 ( .A(n_447), .Y(n_537) );
NAND2xp5_ASAP7_75t_L g538 ( .A(n_399), .B(n_388), .Y(n_538) );
INVx1_ASAP7_75t_L g539 ( .A(n_448), .Y(n_539) );
INVxp67_ASAP7_75t_L g540 ( .A(n_456), .Y(n_540) );
OR2x2_ASAP7_75t_L g541 ( .A(n_463), .B(n_357), .Y(n_541) );
INVx1_ASAP7_75t_SL g542 ( .A(n_465), .Y(n_542) );
INVx1_ASAP7_75t_L g543 ( .A(n_456), .Y(n_543) );
AND2x2_ASAP7_75t_L g544 ( .A(n_410), .B(n_388), .Y(n_544) );
INVx1_ASAP7_75t_L g545 ( .A(n_457), .Y(n_545) );
AND2x2_ASAP7_75t_L g546 ( .A(n_416), .B(n_357), .Y(n_546) );
AND2x4_ASAP7_75t_L g547 ( .A(n_450), .B(n_374), .Y(n_547) );
NOR2xp33_ASAP7_75t_L g548 ( .A(n_458), .B(n_16), .Y(n_548) );
INVx1_ASAP7_75t_L g549 ( .A(n_457), .Y(n_549) );
INVx1_ASAP7_75t_L g550 ( .A(n_460), .Y(n_550) );
NAND2xp5_ASAP7_75t_L g551 ( .A(n_416), .B(n_374), .Y(n_551) );
INVx1_ASAP7_75t_L g552 ( .A(n_460), .Y(n_552) );
INVx1_ASAP7_75t_SL g553 ( .A(n_465), .Y(n_553) );
INVxp67_ASAP7_75t_L g554 ( .A(n_464), .Y(n_554) );
INVx1_ASAP7_75t_L g555 ( .A(n_464), .Y(n_555) );
AND2x2_ASAP7_75t_L g556 ( .A(n_471), .B(n_450), .Y(n_556) );
NAND2xp5_ASAP7_75t_L g557 ( .A(n_537), .B(n_434), .Y(n_557) );
NOR2xp33_ASAP7_75t_L g558 ( .A(n_479), .B(n_459), .Y(n_558) );
INVx1_ASAP7_75t_L g559 ( .A(n_470), .Y(n_559) );
OR2x2_ASAP7_75t_L g560 ( .A(n_473), .B(n_422), .Y(n_560) );
INVx2_ASAP7_75t_L g561 ( .A(n_483), .Y(n_561) );
INVx1_ASAP7_75t_L g562 ( .A(n_539), .Y(n_562) );
INVx1_ASAP7_75t_L g563 ( .A(n_504), .Y(n_563) );
OR2x2_ASAP7_75t_L g564 ( .A(n_473), .B(n_421), .Y(n_564) );
NAND2xp5_ASAP7_75t_L g565 ( .A(n_488), .B(n_451), .Y(n_565) );
NAND2x1p5_ASAP7_75t_L g566 ( .A(n_500), .B(n_454), .Y(n_566) );
AND2x2_ASAP7_75t_L g567 ( .A(n_475), .B(n_451), .Y(n_567) );
INVx1_ASAP7_75t_L g568 ( .A(n_505), .Y(n_568) );
NAND2xp5_ASAP7_75t_L g569 ( .A(n_507), .B(n_425), .Y(n_569) );
NAND2xp5_ASAP7_75t_L g570 ( .A(n_488), .B(n_427), .Y(n_570) );
NAND2xp5_ASAP7_75t_L g571 ( .A(n_481), .B(n_421), .Y(n_571) );
OR2x2_ASAP7_75t_L g572 ( .A(n_468), .B(n_507), .Y(n_572) );
INVx1_ASAP7_75t_L g573 ( .A(n_517), .Y(n_573) );
NAND2xp5_ASAP7_75t_SL g574 ( .A(n_500), .B(n_438), .Y(n_574) );
AND2x2_ASAP7_75t_L g575 ( .A(n_487), .B(n_453), .Y(n_575) );
INVx2_ASAP7_75t_L g576 ( .A(n_498), .Y(n_576) );
INVx1_ASAP7_75t_L g577 ( .A(n_521), .Y(n_577) );
NAND2xp5_ASAP7_75t_L g578 ( .A(n_524), .B(n_390), .Y(n_578) );
NAND2xp5_ASAP7_75t_L g579 ( .A(n_528), .B(n_407), .Y(n_579) );
AND2x2_ASAP7_75t_L g580 ( .A(n_489), .B(n_453), .Y(n_580) );
NAND2xp5_ASAP7_75t_L g581 ( .A(n_536), .B(n_407), .Y(n_581) );
AND2x2_ASAP7_75t_L g582 ( .A(n_493), .B(n_497), .Y(n_582) );
INVx1_ASAP7_75t_L g583 ( .A(n_477), .Y(n_583) );
INVx2_ASAP7_75t_L g584 ( .A(n_498), .Y(n_584) );
AOI211xp5_ASAP7_75t_L g585 ( .A1(n_523), .A2(n_449), .B(n_463), .C(n_438), .Y(n_585) );
OR2x2_ASAP7_75t_L g586 ( .A(n_472), .B(n_462), .Y(n_586) );
NAND2xp5_ASAP7_75t_L g587 ( .A(n_480), .B(n_409), .Y(n_587) );
INVx2_ASAP7_75t_L g588 ( .A(n_519), .Y(n_588) );
INVx1_ASAP7_75t_L g589 ( .A(n_484), .Y(n_589) );
NAND2xp33_ASAP7_75t_L g590 ( .A(n_510), .B(n_409), .Y(n_590) );
INVx1_ASAP7_75t_SL g591 ( .A(n_519), .Y(n_591) );
INVxp67_ASAP7_75t_SL g592 ( .A(n_513), .Y(n_592) );
INVx1_ASAP7_75t_L g593 ( .A(n_491), .Y(n_593) );
NOR4xp25_ASAP7_75t_L g594 ( .A(n_548), .B(n_490), .C(n_492), .D(n_495), .Y(n_594) );
INVx1_ASAP7_75t_L g595 ( .A(n_496), .Y(n_595) );
NAND2xp5_ASAP7_75t_L g596 ( .A(n_499), .B(n_420), .Y(n_596) );
NAND2xp5_ASAP7_75t_L g597 ( .A(n_515), .B(n_420), .Y(n_597) );
INVx1_ASAP7_75t_L g598 ( .A(n_515), .Y(n_598) );
AND2x2_ASAP7_75t_L g599 ( .A(n_526), .B(n_438), .Y(n_599) );
AND2x2_ASAP7_75t_L g600 ( .A(n_531), .B(n_454), .Y(n_600) );
INVx1_ASAP7_75t_L g601 ( .A(n_474), .Y(n_601) );
NAND2xp5_ASAP7_75t_L g602 ( .A(n_516), .B(n_430), .Y(n_602) );
NAND2xp5_ASAP7_75t_L g603 ( .A(n_520), .B(n_430), .Y(n_603) );
INVx1_ASAP7_75t_L g604 ( .A(n_494), .Y(n_604) );
NAND2xp5_ASAP7_75t_L g605 ( .A(n_490), .B(n_437), .Y(n_605) );
NAND4xp25_ASAP7_75t_L g606 ( .A(n_523), .B(n_454), .C(n_462), .D(n_452), .Y(n_606) );
INVx2_ASAP7_75t_L g607 ( .A(n_476), .Y(n_607) );
INVx1_ASAP7_75t_L g608 ( .A(n_532), .Y(n_608) );
NAND3xp33_ASAP7_75t_L g609 ( .A(n_495), .B(n_452), .C(n_446), .Y(n_609) );
NAND4xp25_ASAP7_75t_SL g610 ( .A(n_485), .B(n_446), .C(n_441), .D(n_437), .Y(n_610) );
AND2x2_ASAP7_75t_L g611 ( .A(n_544), .B(n_441), .Y(n_611) );
INVx1_ASAP7_75t_L g612 ( .A(n_532), .Y(n_612) );
INVx1_ASAP7_75t_L g613 ( .A(n_534), .Y(n_613) );
INVx1_ASAP7_75t_L g614 ( .A(n_534), .Y(n_614) );
NAND2xp5_ASAP7_75t_L g615 ( .A(n_525), .B(n_16), .Y(n_615) );
AND2x4_ASAP7_75t_L g616 ( .A(n_503), .B(n_17), .Y(n_616) );
AND2x2_ASAP7_75t_L g617 ( .A(n_546), .B(n_17), .Y(n_617) );
INVx1_ASAP7_75t_L g618 ( .A(n_502), .Y(n_618) );
INVx1_ASAP7_75t_L g619 ( .A(n_535), .Y(n_619) );
INVx2_ASAP7_75t_L g620 ( .A(n_482), .Y(n_620) );
CKINVDCx16_ASAP7_75t_R g621 ( .A(n_503), .Y(n_621) );
INVx2_ASAP7_75t_L g622 ( .A(n_522), .Y(n_622) );
NAND2xp5_ASAP7_75t_L g623 ( .A(n_543), .B(n_18), .Y(n_623) );
INVx1_ASAP7_75t_L g624 ( .A(n_538), .Y(n_624) );
INVx1_ASAP7_75t_L g625 ( .A(n_545), .Y(n_625) );
INVx1_ASAP7_75t_L g626 ( .A(n_549), .Y(n_626) );
AOI22xp5_ASAP7_75t_L g627 ( .A1(n_529), .A2(n_380), .B1(n_250), .B2(n_181), .Y(n_627) );
HB1xp67_ASAP7_75t_L g628 ( .A(n_576), .Y(n_628) );
INVx1_ASAP7_75t_SL g629 ( .A(n_591), .Y(n_629) );
NOR2x1_ASAP7_75t_L g630 ( .A(n_616), .B(n_503), .Y(n_630) );
AND2x2_ASAP7_75t_L g631 ( .A(n_621), .B(n_547), .Y(n_631) );
OAI22xp5_ASAP7_75t_L g632 ( .A1(n_616), .A2(n_486), .B1(n_478), .B2(n_514), .Y(n_632) );
INVx1_ASAP7_75t_L g633 ( .A(n_598), .Y(n_633) );
OR2x2_ASAP7_75t_L g634 ( .A(n_564), .B(n_551), .Y(n_634) );
INVx1_ASAP7_75t_L g635 ( .A(n_572), .Y(n_635) );
AOI221xp5_ASAP7_75t_L g636 ( .A1(n_594), .A2(n_551), .B1(n_554), .B2(n_540), .C(n_501), .Y(n_636) );
OR2x2_ASAP7_75t_L g637 ( .A(n_565), .B(n_501), .Y(n_637) );
INVxp33_ASAP7_75t_L g638 ( .A(n_566), .Y(n_638) );
INVx2_ASAP7_75t_L g639 ( .A(n_584), .Y(n_639) );
AND2x2_ASAP7_75t_L g640 ( .A(n_580), .B(n_547), .Y(n_640) );
NOR2xp33_ASAP7_75t_L g641 ( .A(n_558), .B(n_512), .Y(n_641) );
AND2x2_ASAP7_75t_L g642 ( .A(n_582), .B(n_469), .Y(n_642) );
OAI32xp33_ASAP7_75t_L g643 ( .A1(n_606), .A2(n_518), .A3(n_509), .B1(n_553), .B2(n_542), .Y(n_643) );
AND2x2_ASAP7_75t_L g644 ( .A(n_567), .B(n_506), .Y(n_644) );
OAI211xp5_ASAP7_75t_SL g645 ( .A1(n_585), .A2(n_511), .B(n_518), .C(n_542), .Y(n_645) );
INVx1_ASAP7_75t_SL g646 ( .A(n_566), .Y(n_646) );
A2O1A1Ixp33_ASAP7_75t_L g647 ( .A1(n_590), .A2(n_478), .B(n_506), .C(n_553), .Y(n_647) );
AOI22xp5_ASAP7_75t_L g648 ( .A1(n_610), .A2(n_508), .B1(n_552), .B2(n_550), .Y(n_648) );
NAND2xp5_ASAP7_75t_L g649 ( .A(n_557), .B(n_555), .Y(n_649) );
INVx2_ASAP7_75t_L g650 ( .A(n_588), .Y(n_650) );
INVx1_ASAP7_75t_L g651 ( .A(n_568), .Y(n_651) );
NOR2xp33_ASAP7_75t_L g652 ( .A(n_559), .B(n_533), .Y(n_652) );
NAND2xp5_ASAP7_75t_L g653 ( .A(n_557), .B(n_541), .Y(n_653) );
NAND2xp5_ASAP7_75t_L g654 ( .A(n_565), .B(n_530), .Y(n_654) );
HB1xp67_ASAP7_75t_L g655 ( .A(n_571), .Y(n_655) );
AOI221xp5_ASAP7_75t_L g656 ( .A1(n_570), .A2(n_380), .B1(n_181), .B2(n_164), .C(n_19), .Y(n_656) );
INVx1_ASAP7_75t_L g657 ( .A(n_573), .Y(n_657) );
NOR3xp33_ASAP7_75t_SL g658 ( .A(n_615), .B(n_19), .C(n_527), .Y(n_658) );
NAND2x1_ASAP7_75t_L g659 ( .A(n_609), .B(n_527), .Y(n_659) );
NAND2xp5_ASAP7_75t_SL g660 ( .A(n_574), .B(n_527), .Y(n_660) );
NOR2xp33_ASAP7_75t_L g661 ( .A(n_563), .B(n_22), .Y(n_661) );
OAI21xp5_ASAP7_75t_SL g662 ( .A1(n_627), .A2(n_181), .B(n_164), .Y(n_662) );
OAI22xp33_ASAP7_75t_L g663 ( .A1(n_615), .A2(n_248), .B1(n_247), .B2(n_245), .Y(n_663) );
NAND2xp5_ASAP7_75t_L g664 ( .A(n_571), .B(n_181), .Y(n_664) );
INVx1_ASAP7_75t_L g665 ( .A(n_577), .Y(n_665) );
AOI33xp33_ASAP7_75t_L g666 ( .A1(n_617), .A2(n_221), .A3(n_191), .B1(n_27), .B2(n_28), .B3(n_29), .Y(n_666) );
INVx1_ASAP7_75t_L g667 ( .A(n_562), .Y(n_667) );
AOI22xp5_ASAP7_75t_L g668 ( .A1(n_569), .A2(n_164), .B1(n_26), .B2(n_30), .Y(n_668) );
INVx2_ASAP7_75t_L g669 ( .A(n_608), .Y(n_669) );
INVx1_ASAP7_75t_L g670 ( .A(n_583), .Y(n_670) );
NOR3xp33_ASAP7_75t_L g671 ( .A(n_645), .B(n_623), .C(n_625), .Y(n_671) );
AOI22xp33_ASAP7_75t_L g672 ( .A1(n_645), .A2(n_560), .B1(n_600), .B2(n_618), .Y(n_672) );
OAI221xp5_ASAP7_75t_L g673 ( .A1(n_636), .A2(n_626), .B1(n_605), .B2(n_623), .C(n_624), .Y(n_673) );
AOI21xp33_ASAP7_75t_L g674 ( .A1(n_643), .A2(n_614), .B(n_613), .Y(n_674) );
INVx2_ASAP7_75t_SL g675 ( .A(n_631), .Y(n_675) );
AOI221xp5_ASAP7_75t_L g676 ( .A1(n_655), .A2(n_619), .B1(n_592), .B2(n_601), .C(n_604), .Y(n_676) );
AO22x1_ASAP7_75t_L g677 ( .A1(n_630), .A2(n_620), .B1(n_607), .B2(n_561), .Y(n_677) );
AOI221xp5_ASAP7_75t_L g678 ( .A1(n_655), .A2(n_612), .B1(n_593), .B2(n_595), .C(n_589), .Y(n_678) );
AOI22xp5_ASAP7_75t_L g679 ( .A1(n_632), .A2(n_658), .B1(n_641), .B2(n_629), .Y(n_679) );
NAND2xp5_ASAP7_75t_L g680 ( .A(n_635), .B(n_605), .Y(n_680) );
AOI221xp5_ASAP7_75t_L g681 ( .A1(n_652), .A2(n_597), .B1(n_581), .B2(n_578), .C(n_579), .Y(n_681) );
OAI221xp5_ASAP7_75t_L g682 ( .A1(n_647), .A2(n_597), .B1(n_579), .B2(n_581), .C(n_578), .Y(n_682) );
OAI21xp33_ASAP7_75t_SL g683 ( .A1(n_660), .A2(n_556), .B(n_599), .Y(n_683) );
AOI222xp33_ASAP7_75t_L g684 ( .A1(n_656), .A2(n_603), .B1(n_602), .B2(n_611), .C1(n_596), .C2(n_587), .Y(n_684) );
AOI221xp5_ASAP7_75t_L g685 ( .A1(n_652), .A2(n_575), .B1(n_603), .B2(n_602), .C(n_596), .Y(n_685) );
AND2x2_ASAP7_75t_L g686 ( .A(n_644), .B(n_586), .Y(n_686) );
AOI22xp33_ASAP7_75t_L g687 ( .A1(n_654), .A2(n_622), .B1(n_587), .B2(n_164), .Y(n_687) );
OAI221xp5_ASAP7_75t_SL g688 ( .A1(n_662), .A2(n_25), .B1(n_34), .B2(n_35), .C(n_36), .Y(n_688) );
AOI322xp5_ASAP7_75t_L g689 ( .A1(n_658), .A2(n_164), .A3(n_44), .B1(n_45), .B2(n_46), .C1(n_48), .C2(n_52), .Y(n_689) );
AND2x2_ASAP7_75t_L g690 ( .A(n_640), .B(n_38), .Y(n_690) );
OAI221xp5_ASAP7_75t_SL g691 ( .A1(n_646), .A2(n_54), .B1(n_56), .B2(n_57), .C(n_58), .Y(n_691) );
INVx1_ASAP7_75t_L g692 ( .A(n_633), .Y(n_692) );
NOR3xp33_ASAP7_75t_L g693 ( .A(n_664), .B(n_60), .C(n_63), .Y(n_693) );
AOI221x1_ASAP7_75t_L g694 ( .A1(n_651), .A2(n_65), .B1(n_68), .B2(n_69), .C(n_72), .Y(n_694) );
NOR3xp33_ASAP7_75t_L g695 ( .A(n_659), .B(n_663), .C(n_666), .Y(n_695) );
AOI22xp5_ASAP7_75t_L g696 ( .A1(n_648), .A2(n_73), .B1(n_74), .B2(n_75), .Y(n_696) );
AOI322xp5_ASAP7_75t_L g697 ( .A1(n_642), .A2(n_77), .A3(n_80), .B1(n_81), .B2(n_82), .C1(n_83), .C2(n_84), .Y(n_697) );
INVx1_ASAP7_75t_L g698 ( .A(n_670), .Y(n_698) );
AOI221xp5_ASAP7_75t_L g699 ( .A1(n_657), .A2(n_86), .B1(n_87), .B2(n_91), .C(n_93), .Y(n_699) );
NOR2xp33_ASAP7_75t_SL g700 ( .A(n_638), .B(n_661), .Y(n_700) );
AOI211xp5_ASAP7_75t_L g701 ( .A1(n_663), .A2(n_661), .B(n_628), .C(n_637), .Y(n_701) );
NAND2xp5_ASAP7_75t_L g702 ( .A(n_669), .B(n_649), .Y(n_702) );
NOR3xp33_ASAP7_75t_SL g703 ( .A(n_653), .B(n_665), .C(n_667), .Y(n_703) );
AOI211xp5_ASAP7_75t_L g704 ( .A1(n_628), .A2(n_634), .B(n_639), .C(n_650), .Y(n_704) );
OAI211xp5_ASAP7_75t_SL g705 ( .A1(n_668), .A2(n_658), .B(n_636), .C(n_630), .Y(n_705) );
NAND4xp25_ASAP7_75t_SL g706 ( .A(n_683), .B(n_679), .C(n_672), .D(n_701), .Y(n_706) );
AOI221x1_ASAP7_75t_L g707 ( .A1(n_705), .A2(n_695), .B1(n_671), .B2(n_674), .C(n_693), .Y(n_707) );
AND4x1_ASAP7_75t_L g708 ( .A(n_700), .B(n_703), .C(n_684), .D(n_696), .Y(n_708) );
AOI22xp5_ASAP7_75t_L g709 ( .A1(n_673), .A2(n_682), .B1(n_675), .B2(n_677), .Y(n_709) );
NAND2xp5_ASAP7_75t_L g710 ( .A(n_678), .B(n_681), .Y(n_710) );
NAND2xp5_ASAP7_75t_L g711 ( .A(n_676), .B(n_685), .Y(n_711) );
NOR2x1_ASAP7_75t_L g712 ( .A(n_706), .B(n_690), .Y(n_712) );
NAND4xp25_ASAP7_75t_L g713 ( .A(n_707), .B(n_689), .C(n_697), .D(n_691), .Y(n_713) );
INVx1_ASAP7_75t_L g714 ( .A(n_711), .Y(n_714) );
NAND2xp5_ASAP7_75t_L g715 ( .A(n_710), .B(n_698), .Y(n_715) );
INVx1_ASAP7_75t_L g716 ( .A(n_715), .Y(n_716) );
OR2x2_ASAP7_75t_L g717 ( .A(n_714), .B(n_709), .Y(n_717) );
NAND3xp33_ASAP7_75t_L g718 ( .A(n_712), .B(n_708), .C(n_691), .Y(n_718) );
AOI22xp5_ASAP7_75t_L g719 ( .A1(n_718), .A2(n_713), .B1(n_704), .B2(n_687), .Y(n_719) );
XOR2x2_ASAP7_75t_L g720 ( .A(n_717), .B(n_688), .Y(n_720) );
CKINVDCx5p33_ASAP7_75t_R g721 ( .A(n_720), .Y(n_721) );
AOI22x1_ASAP7_75t_L g722 ( .A1(n_719), .A2(n_716), .B1(n_692), .B2(n_686), .Y(n_722) );
INVx1_ASAP7_75t_L g723 ( .A(n_722), .Y(n_723) );
OAI22xp5_ASAP7_75t_L g724 ( .A1(n_723), .A2(n_721), .B1(n_680), .B2(n_702), .Y(n_724) );
INVx1_ASAP7_75t_L g725 ( .A(n_724), .Y(n_725) );
XNOR2xp5_ASAP7_75t_L g726 ( .A(n_725), .B(n_699), .Y(n_726) );
AOI21xp5_ASAP7_75t_L g727 ( .A1(n_726), .A2(n_688), .B(n_694), .Y(n_727) );
endmodule