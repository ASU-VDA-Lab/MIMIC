module fake_jpeg_24649_n_325 (n_13, n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_325);

input n_13;
input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_325;

wire n_253;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_15;
wire n_141;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_14;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

CKINVDCx16_ASAP7_75t_R g14 ( 
.A(n_7),
.Y(n_14)
);

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_4),
.Y(n_15)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_5),
.Y(n_16)
);

INVx3_ASAP7_75t_L g17 ( 
.A(n_10),
.Y(n_17)
);

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_1),
.Y(n_18)
);

INVx2_ASAP7_75t_L g19 ( 
.A(n_7),
.Y(n_19)
);

BUFx4f_ASAP7_75t_SL g20 ( 
.A(n_11),
.Y(n_20)
);

BUFx12_ASAP7_75t_L g21 ( 
.A(n_7),
.Y(n_21)
);

BUFx12f_ASAP7_75t_L g22 ( 
.A(n_13),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_13),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_3),
.Y(n_24)
);

CKINVDCx16_ASAP7_75t_R g25 ( 
.A(n_12),
.Y(n_25)
);

INVx8_ASAP7_75t_L g26 ( 
.A(n_11),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_2),
.Y(n_27)
);

BUFx12_ASAP7_75t_L g28 ( 
.A(n_9),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_8),
.Y(n_29)
);

INVx2_ASAP7_75t_L g30 ( 
.A(n_26),
.Y(n_30)
);

INVx6_ASAP7_75t_L g49 ( 
.A(n_30),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_20),
.Y(n_31)
);

INVx8_ASAP7_75t_L g60 ( 
.A(n_31),
.Y(n_60)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_27),
.Y(n_32)
);

NOR2xp33_ASAP7_75t_L g43 ( 
.A(n_32),
.B(n_33),
.Y(n_43)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_27),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_15),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_34),
.B(n_37),
.Y(n_53)
);

INVx1_ASAP7_75t_SL g35 ( 
.A(n_20),
.Y(n_35)
);

INVx4_ASAP7_75t_L g55 ( 
.A(n_35),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_20),
.Y(n_36)
);

BUFx2_ASAP7_75t_L g45 ( 
.A(n_36),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_15),
.Y(n_37)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_22),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_L g41 ( 
.A(n_38),
.B(n_19),
.Y(n_41)
);

BUFx5_ASAP7_75t_L g39 ( 
.A(n_22),
.Y(n_39)
);

INVx3_ASAP7_75t_L g50 ( 
.A(n_39),
.Y(n_50)
);

INVx11_ASAP7_75t_L g40 ( 
.A(n_20),
.Y(n_40)
);

AOI22xp33_ASAP7_75t_SL g42 ( 
.A1(n_40),
.A2(n_26),
.B1(n_20),
.B2(n_22),
.Y(n_42)
);

CKINVDCx16_ASAP7_75t_R g81 ( 
.A(n_41),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_42),
.B(n_54),
.Y(n_61)
);

OR2x2_ASAP7_75t_L g44 ( 
.A(n_34),
.B(n_22),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_SL g80 ( 
.A(n_44),
.B(n_47),
.Y(n_80)
);

AOI22xp33_ASAP7_75t_SL g46 ( 
.A1(n_40),
.A2(n_26),
.B1(n_17),
.B2(n_19),
.Y(n_46)
);

OAI22xp5_ASAP7_75t_L g82 ( 
.A1(n_46),
.A2(n_51),
.B1(n_30),
.B2(n_35),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g47 ( 
.A(n_34),
.B(n_29),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_37),
.B(n_29),
.Y(n_48)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_48),
.Y(n_64)
);

OAI22xp5_ASAP7_75t_L g51 ( 
.A1(n_30),
.A2(n_19),
.B1(n_17),
.B2(n_26),
.Y(n_51)
);

OR2x2_ASAP7_75t_L g52 ( 
.A(n_37),
.B(n_22),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_L g62 ( 
.A(n_52),
.B(n_56),
.Y(n_62)
);

INVx2_ASAP7_75t_L g54 ( 
.A(n_39),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_L g56 ( 
.A(n_38),
.B(n_18),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g57 ( 
.A(n_32),
.B(n_29),
.Y(n_57)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_57),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_SL g58 ( 
.A(n_32),
.B(n_23),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_L g66 ( 
.A(n_58),
.B(n_59),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_33),
.B(n_23),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_54),
.B(n_40),
.Y(n_63)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_63),
.Y(n_94)
);

INVx2_ASAP7_75t_L g65 ( 
.A(n_60),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_65),
.B(n_75),
.Y(n_89)
);

BUFx12f_ASAP7_75t_L g67 ( 
.A(n_50),
.Y(n_67)
);

BUFx3_ASAP7_75t_L g103 ( 
.A(n_67),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_54),
.B(n_40),
.Y(n_68)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_68),
.Y(n_96)
);

MAJIxp5_ASAP7_75t_L g69 ( 
.A(n_56),
.B(n_35),
.C(n_38),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_L g90 ( 
.A(n_69),
.B(n_70),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_L g70 ( 
.A(n_44),
.B(n_38),
.Y(n_70)
);

BUFx6f_ASAP7_75t_L g71 ( 
.A(n_60),
.Y(n_71)
);

INVxp67_ASAP7_75t_L g85 ( 
.A(n_71),
.Y(n_85)
);

BUFx6f_ASAP7_75t_L g72 ( 
.A(n_60),
.Y(n_72)
);

INVx2_ASAP7_75t_L g86 ( 
.A(n_72),
.Y(n_86)
);

OAI22xp33_ASAP7_75t_SL g73 ( 
.A1(n_51),
.A2(n_30),
.B1(n_17),
.B2(n_40),
.Y(n_73)
);

AOI22xp5_ASAP7_75t_SL g98 ( 
.A1(n_73),
.A2(n_55),
.B1(n_41),
.B2(n_50),
.Y(n_98)
);

BUFx6f_ASAP7_75t_L g74 ( 
.A(n_60),
.Y(n_74)
);

INVx2_ASAP7_75t_L g99 ( 
.A(n_74),
.Y(n_99)
);

INVx2_ASAP7_75t_L g75 ( 
.A(n_51),
.Y(n_75)
);

BUFx2_ASAP7_75t_L g76 ( 
.A(n_45),
.Y(n_76)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_76),
.Y(n_101)
);

BUFx6f_ASAP7_75t_L g78 ( 
.A(n_45),
.Y(n_78)
);

INVx2_ASAP7_75t_L g100 ( 
.A(n_78),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_50),
.B(n_21),
.Y(n_79)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_79),
.Y(n_104)
);

AOI22xp5_ASAP7_75t_L g95 ( 
.A1(n_82),
.A2(n_49),
.B1(n_41),
.B2(n_55),
.Y(n_95)
);

O2A1O1Ixp33_ASAP7_75t_SL g83 ( 
.A1(n_56),
.A2(n_39),
.B(n_22),
.C(n_35),
.Y(n_83)
);

AOI22xp5_ASAP7_75t_SL g109 ( 
.A1(n_83),
.A2(n_42),
.B1(n_44),
.B2(n_52),
.Y(n_109)
);

INVx2_ASAP7_75t_L g84 ( 
.A(n_49),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_84),
.B(n_49),
.Y(n_91)
);

CKINVDCx20_ASAP7_75t_R g87 ( 
.A(n_67),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g120 ( 
.A(n_87),
.B(n_95),
.Y(n_120)
);

AOI22xp33_ASAP7_75t_SL g88 ( 
.A1(n_75),
.A2(n_55),
.B1(n_50),
.B2(n_49),
.Y(n_88)
);

AOI21xp5_ASAP7_75t_L g131 ( 
.A1(n_88),
.A2(n_92),
.B(n_109),
.Y(n_131)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_91),
.Y(n_112)
);

OAI21xp33_ASAP7_75t_L g92 ( 
.A1(n_70),
.A2(n_44),
.B(n_52),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_64),
.B(n_58),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_SL g116 ( 
.A(n_93),
.B(n_97),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_64),
.B(n_58),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g121 ( 
.A(n_98),
.B(n_61),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_77),
.B(n_59),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_SL g117 ( 
.A(n_102),
.B(n_108),
.Y(n_117)
);

INVx2_ASAP7_75t_L g105 ( 
.A(n_67),
.Y(n_105)
);

INVx6_ASAP7_75t_L g115 ( 
.A(n_105),
.Y(n_115)
);

AOI22xp5_ASAP7_75t_L g106 ( 
.A1(n_82),
.A2(n_55),
.B1(n_46),
.B2(n_39),
.Y(n_106)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_106),
.Y(n_113)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_80),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_L g114 ( 
.A(n_107),
.B(n_66),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_SL g108 ( 
.A(n_66),
.B(n_43),
.Y(n_108)
);

INVx2_ASAP7_75t_L g110 ( 
.A(n_103),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_L g137 ( 
.A(n_110),
.B(n_111),
.Y(n_137)
);

INVx4_ASAP7_75t_L g111 ( 
.A(n_103),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_SL g150 ( 
.A(n_114),
.B(n_118),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_SL g118 ( 
.A(n_108),
.B(n_80),
.Y(n_118)
);

INVx3_ASAP7_75t_L g119 ( 
.A(n_103),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_L g146 ( 
.A(n_119),
.B(n_122),
.Y(n_146)
);

AOI22xp5_ASAP7_75t_L g143 ( 
.A1(n_121),
.A2(n_129),
.B1(n_83),
.B2(n_97),
.Y(n_143)
);

INVx4_ASAP7_75t_L g122 ( 
.A(n_87),
.Y(n_122)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_89),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_SL g151 ( 
.A(n_123),
.B(n_125),
.Y(n_151)
);

INVx2_ASAP7_75t_L g124 ( 
.A(n_105),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_L g148 ( 
.A(n_124),
.B(n_126),
.Y(n_148)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_89),
.Y(n_125)
);

INVx4_ASAP7_75t_L g126 ( 
.A(n_85),
.Y(n_126)
);

INVx8_ASAP7_75t_L g127 ( 
.A(n_86),
.Y(n_127)
);

INVx2_ASAP7_75t_L g154 ( 
.A(n_127),
.Y(n_154)
);

INVx8_ASAP7_75t_L g128 ( 
.A(n_86),
.Y(n_128)
);

CKINVDCx14_ASAP7_75t_R g160 ( 
.A(n_128),
.Y(n_160)
);

O2A1O1Ixp33_ASAP7_75t_SL g129 ( 
.A1(n_109),
.A2(n_62),
.B(n_83),
.C(n_81),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_L g130 ( 
.A(n_94),
.B(n_77),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_SL g161 ( 
.A(n_130),
.B(n_134),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_L g132 ( 
.A(n_90),
.B(n_62),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_L g144 ( 
.A(n_132),
.B(n_135),
.Y(n_144)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_91),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_SL g155 ( 
.A(n_133),
.B(n_101),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_L g134 ( 
.A(n_94),
.B(n_67),
.Y(n_134)
);

OR2x2_ASAP7_75t_L g135 ( 
.A(n_93),
.B(n_53),
.Y(n_135)
);

XOR2xp5_ASAP7_75t_L g136 ( 
.A(n_132),
.B(n_90),
.Y(n_136)
);

MAJIxp5_ASAP7_75t_L g180 ( 
.A(n_136),
.B(n_142),
.C(n_23),
.Y(n_180)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_122),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_SL g166 ( 
.A(n_138),
.B(n_140),
.Y(n_166)
);

OAI22xp5_ASAP7_75t_SL g139 ( 
.A1(n_113),
.A2(n_109),
.B1(n_106),
.B2(n_95),
.Y(n_139)
);

OAI22xp5_ASAP7_75t_SL g169 ( 
.A1(n_139),
.A2(n_133),
.B1(n_112),
.B2(n_43),
.Y(n_169)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_126),
.Y(n_140)
);

AND2x2_ASAP7_75t_L g141 ( 
.A(n_129),
.B(n_69),
.Y(n_141)
);

OAI21xp5_ASAP7_75t_SL g177 ( 
.A1(n_141),
.A2(n_153),
.B(n_57),
.Y(n_177)
);

MAJIxp5_ASAP7_75t_L g142 ( 
.A(n_131),
.B(n_104),
.C(n_107),
.Y(n_142)
);

OAI21xp5_ASAP7_75t_L g173 ( 
.A1(n_143),
.A2(n_144),
.B(n_159),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_L g145 ( 
.A(n_118),
.B(n_102),
.Y(n_145)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_145),
.Y(n_167)
);

NOR2xp67_ASAP7_75t_L g147 ( 
.A(n_135),
.B(n_98),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_L g168 ( 
.A(n_147),
.B(n_116),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_L g149 ( 
.A(n_117),
.B(n_96),
.Y(n_149)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_149),
.Y(n_170)
);

AOI22xp5_ASAP7_75t_L g152 ( 
.A1(n_113),
.A2(n_88),
.B1(n_96),
.B2(n_104),
.Y(n_152)
);

OAI22xp5_ASAP7_75t_L g187 ( 
.A1(n_152),
.A2(n_156),
.B1(n_159),
.B2(n_115),
.Y(n_187)
);

AND2x2_ASAP7_75t_L g153 ( 
.A(n_129),
.B(n_52),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_SL g175 ( 
.A(n_155),
.B(n_47),
.Y(n_175)
);

AOI22xp5_ASAP7_75t_L g156 ( 
.A1(n_120),
.A2(n_65),
.B1(n_84),
.B2(n_99),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_L g157 ( 
.A(n_117),
.B(n_53),
.Y(n_157)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_157),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_L g158 ( 
.A(n_114),
.B(n_48),
.Y(n_158)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_158),
.Y(n_185)
);

AOI22xp5_ASAP7_75t_L g159 ( 
.A1(n_131),
.A2(n_99),
.B1(n_101),
.B2(n_100),
.Y(n_159)
);

AOI22xp5_ASAP7_75t_SL g162 ( 
.A1(n_145),
.A2(n_125),
.B1(n_123),
.B2(n_135),
.Y(n_162)
);

OAI21xp5_ASAP7_75t_SL g192 ( 
.A1(n_162),
.A2(n_172),
.B(n_177),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_L g163 ( 
.A(n_144),
.B(n_116),
.Y(n_163)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_163),
.Y(n_198)
);

CKINVDCx20_ASAP7_75t_R g164 ( 
.A(n_148),
.Y(n_164)
);

CKINVDCx20_ASAP7_75t_R g202 ( 
.A(n_164),
.Y(n_202)
);

INVx2_ASAP7_75t_L g165 ( 
.A(n_154),
.Y(n_165)
);

NOR2xp33_ASAP7_75t_L g197 ( 
.A(n_165),
.B(n_178),
.Y(n_197)
);

OAI21xp5_ASAP7_75t_L g190 ( 
.A1(n_168),
.A2(n_173),
.B(n_151),
.Y(n_190)
);

AOI22xp5_ASAP7_75t_L g209 ( 
.A1(n_169),
.A2(n_187),
.B1(n_167),
.B2(n_179),
.Y(n_209)
);

NOR2xp33_ASAP7_75t_L g171 ( 
.A(n_154),
.B(n_111),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_SL g195 ( 
.A(n_171),
.B(n_175),
.Y(n_195)
);

AOI22xp5_ASAP7_75t_SL g172 ( 
.A1(n_157),
.A2(n_112),
.B1(n_59),
.B2(n_127),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_L g174 ( 
.A(n_150),
.B(n_47),
.Y(n_174)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_174),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_L g176 ( 
.A(n_150),
.B(n_48),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_L g203 ( 
.A(n_176),
.B(n_181),
.Y(n_203)
);

INVx2_ASAP7_75t_L g178 ( 
.A(n_160),
.Y(n_178)
);

XNOR2xp5_ASAP7_75t_L g191 ( 
.A(n_180),
.B(n_186),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_L g181 ( 
.A(n_136),
.B(n_128),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_L g182 ( 
.A(n_149),
.B(n_115),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_L g205 ( 
.A(n_182),
.B(n_156),
.Y(n_205)
);

A2O1A1Ixp33_ASAP7_75t_L g183 ( 
.A1(n_143),
.A2(n_153),
.B(n_141),
.C(n_158),
.Y(n_183)
);

OAI21xp5_ASAP7_75t_SL g196 ( 
.A1(n_183),
.A2(n_184),
.B(n_169),
.Y(n_196)
);

OA22x2_ASAP7_75t_L g184 ( 
.A1(n_152),
.A2(n_71),
.B1(n_72),
.B2(n_74),
.Y(n_184)
);

XNOR2xp5_ASAP7_75t_L g186 ( 
.A(n_142),
.B(n_36),
.Y(n_186)
);

NOR2xp33_ASAP7_75t_L g188 ( 
.A(n_137),
.B(n_119),
.Y(n_188)
);

NOR2xp33_ASAP7_75t_L g211 ( 
.A(n_188),
.B(n_76),
.Y(n_211)
);

INVxp33_ASAP7_75t_L g189 ( 
.A(n_166),
.Y(n_189)
);

NOR2xp33_ASAP7_75t_L g218 ( 
.A(n_189),
.B(n_199),
.Y(n_218)
);

NOR2xp33_ASAP7_75t_SL g214 ( 
.A(n_190),
.B(n_172),
.Y(n_214)
);

AND2x2_ASAP7_75t_L g193 ( 
.A(n_182),
.B(n_139),
.Y(n_193)
);

AOI21xp5_ASAP7_75t_L g232 ( 
.A1(n_193),
.A2(n_194),
.B(n_196),
.Y(n_232)
);

AOI21xp5_ASAP7_75t_L g194 ( 
.A1(n_177),
.A2(n_138),
.B(n_146),
.Y(n_194)
);

OAI21xp5_ASAP7_75t_L g199 ( 
.A1(n_173),
.A2(n_153),
.B(n_141),
.Y(n_199)
);

OAI22xp5_ASAP7_75t_SL g200 ( 
.A1(n_183),
.A2(n_181),
.B1(n_162),
.B2(n_163),
.Y(n_200)
);

AOI22xp5_ASAP7_75t_L g222 ( 
.A1(n_200),
.A2(n_208),
.B1(n_185),
.B2(n_176),
.Y(n_222)
);

INVx3_ASAP7_75t_L g201 ( 
.A(n_165),
.Y(n_201)
);

NOR2xp33_ASAP7_75t_L g220 ( 
.A(n_201),
.B(n_76),
.Y(n_220)
);

CKINVDCx20_ASAP7_75t_R g204 ( 
.A(n_164),
.Y(n_204)
);

CKINVDCx20_ASAP7_75t_R g219 ( 
.A(n_204),
.Y(n_219)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_205),
.Y(n_221)
);

AOI22xp5_ASAP7_75t_SL g206 ( 
.A1(n_170),
.A2(n_140),
.B1(n_110),
.B2(n_161),
.Y(n_206)
);

OAI22xp5_ASAP7_75t_L g217 ( 
.A1(n_206),
.A2(n_207),
.B1(n_209),
.B2(n_213),
.Y(n_217)
);

OAI21xp5_ASAP7_75t_SL g207 ( 
.A1(n_170),
.A2(n_124),
.B(n_100),
.Y(n_207)
);

OAI22xp5_ASAP7_75t_SL g208 ( 
.A1(n_167),
.A2(n_16),
.B1(n_33),
.B2(n_24),
.Y(n_208)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_211),
.Y(n_229)
);

BUFx3_ASAP7_75t_L g212 ( 
.A(n_178),
.Y(n_212)
);

CKINVDCx20_ASAP7_75t_R g228 ( 
.A(n_212),
.Y(n_228)
);

AOI22xp5_ASAP7_75t_L g213 ( 
.A1(n_179),
.A2(n_16),
.B1(n_15),
.B2(n_24),
.Y(n_213)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_214),
.Y(n_237)
);

CKINVDCx16_ASAP7_75t_R g215 ( 
.A(n_197),
.Y(n_215)
);

NAND2xp5_ASAP7_75t_L g245 ( 
.A(n_215),
.B(n_216),
.Y(n_245)
);

INVxp67_ASAP7_75t_L g216 ( 
.A(n_212),
.Y(n_216)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_220),
.Y(n_244)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_222),
.Y(n_246)
);

AO22x1_ASAP7_75t_L g223 ( 
.A1(n_193),
.A2(n_196),
.B1(n_205),
.B2(n_199),
.Y(n_223)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_223),
.Y(n_248)
);

OAI22xp5_ASAP7_75t_L g224 ( 
.A1(n_209),
.A2(n_184),
.B1(n_185),
.B2(n_174),
.Y(n_224)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_224),
.Y(n_255)
);

NOR2xp33_ASAP7_75t_L g225 ( 
.A(n_201),
.B(n_184),
.Y(n_225)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_225),
.Y(n_254)
);

NOR2xp33_ASAP7_75t_L g226 ( 
.A(n_202),
.B(n_184),
.Y(n_226)
);

CKINVDCx20_ASAP7_75t_R g249 ( 
.A(n_226),
.Y(n_249)
);

INVx8_ASAP7_75t_L g227 ( 
.A(n_193),
.Y(n_227)
);

AOI22xp5_ASAP7_75t_SL g252 ( 
.A1(n_227),
.A2(n_234),
.B1(n_235),
.B2(n_229),
.Y(n_252)
);

AOI22xp5_ASAP7_75t_SL g230 ( 
.A1(n_198),
.A2(n_186),
.B1(n_180),
.B2(n_16),
.Y(n_230)
);

OAI22xp5_ASAP7_75t_L g250 ( 
.A1(n_230),
.A2(n_208),
.B1(n_14),
.B2(n_25),
.Y(n_250)
);

OAI221xp5_ASAP7_75t_L g231 ( 
.A1(n_198),
.A2(n_36),
.B1(n_31),
.B2(n_24),
.C(n_45),
.Y(n_231)
);

XNOR2xp5_ASAP7_75t_L g236 ( 
.A(n_231),
.B(n_213),
.Y(n_236)
);

CKINVDCx16_ASAP7_75t_R g233 ( 
.A(n_207),
.Y(n_233)
);

BUFx24_ASAP7_75t_SL g240 ( 
.A(n_233),
.Y(n_240)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_203),
.Y(n_234)
);

NAND2xp5_ASAP7_75t_L g235 ( 
.A(n_210),
.B(n_0),
.Y(n_235)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_236),
.Y(n_262)
);

XNOR2xp5_ASAP7_75t_SL g238 ( 
.A(n_223),
.B(n_200),
.Y(n_238)
);

XOR2xp5_ASAP7_75t_L g265 ( 
.A(n_238),
.B(n_231),
.Y(n_265)
);

FAx1_ASAP7_75t_SL g239 ( 
.A(n_223),
.B(n_203),
.CI(n_190),
.CON(n_239),
.SN(n_239)
);

NOR2xp33_ASAP7_75t_L g272 ( 
.A(n_239),
.B(n_28),
.Y(n_272)
);

MAJIxp5_ASAP7_75t_L g241 ( 
.A(n_218),
.B(n_234),
.C(n_221),
.Y(n_241)
);

MAJIxp5_ASAP7_75t_L g256 ( 
.A(n_241),
.B(n_243),
.C(n_247),
.Y(n_256)
);

AOI22xp5_ASAP7_75t_L g242 ( 
.A1(n_227),
.A2(n_210),
.B1(n_192),
.B2(n_206),
.Y(n_242)
);

OAI22xp5_ASAP7_75t_SL g259 ( 
.A1(n_242),
.A2(n_251),
.B1(n_252),
.B2(n_253),
.Y(n_259)
);

MAJIxp5_ASAP7_75t_L g243 ( 
.A(n_221),
.B(n_194),
.C(n_192),
.Y(n_243)
);

MAJIxp5_ASAP7_75t_L g247 ( 
.A(n_232),
.B(n_191),
.C(n_195),
.Y(n_247)
);

XNOR2xp5_ASAP7_75t_L g271 ( 
.A(n_250),
.B(n_31),
.Y(n_271)
);

OAI22xp5_ASAP7_75t_L g251 ( 
.A1(n_232),
.A2(n_191),
.B1(n_25),
.B2(n_14),
.Y(n_251)
);

OAI22xp5_ASAP7_75t_L g253 ( 
.A1(n_222),
.A2(n_18),
.B1(n_11),
.B2(n_13),
.Y(n_253)
);

OAI21xp5_ASAP7_75t_L g257 ( 
.A1(n_248),
.A2(n_219),
.B(n_216),
.Y(n_257)
);

NAND2xp5_ASAP7_75t_L g282 ( 
.A(n_257),
.B(n_258),
.Y(n_282)
);

OR2x2_ASAP7_75t_L g258 ( 
.A(n_249),
.B(n_219),
.Y(n_258)
);

NAND2xp5_ASAP7_75t_L g260 ( 
.A(n_244),
.B(n_229),
.Y(n_260)
);

NOR2xp33_ASAP7_75t_SL g284 ( 
.A(n_260),
.B(n_263),
.Y(n_284)
);

XNOR2xp5_ASAP7_75t_SL g261 ( 
.A(n_242),
.B(n_217),
.Y(n_261)
);

MAJIxp5_ASAP7_75t_L g273 ( 
.A(n_261),
.B(n_265),
.C(n_267),
.Y(n_273)
);

NAND2xp5_ASAP7_75t_L g263 ( 
.A(n_245),
.B(n_235),
.Y(n_263)
);

OAI22xp5_ASAP7_75t_L g264 ( 
.A1(n_255),
.A2(n_214),
.B1(n_230),
.B2(n_228),
.Y(n_264)
);

AOI22xp5_ASAP7_75t_L g275 ( 
.A1(n_264),
.A2(n_271),
.B1(n_259),
.B2(n_246),
.Y(n_275)
);

NAND2xp5_ASAP7_75t_L g266 ( 
.A(n_252),
.B(n_228),
.Y(n_266)
);

INVxp67_ASAP7_75t_L g286 ( 
.A(n_266),
.Y(n_286)
);

MAJIxp5_ASAP7_75t_L g267 ( 
.A(n_247),
.B(n_78),
.C(n_45),
.Y(n_267)
);

MAJIxp5_ASAP7_75t_L g268 ( 
.A(n_241),
.B(n_45),
.C(n_36),
.Y(n_268)
);

MAJIxp5_ASAP7_75t_L g276 ( 
.A(n_268),
.B(n_269),
.C(n_238),
.Y(n_276)
);

MAJIxp5_ASAP7_75t_L g269 ( 
.A(n_243),
.B(n_36),
.C(n_31),
.Y(n_269)
);

NAND2xp5_ASAP7_75t_L g270 ( 
.A(n_254),
.B(n_31),
.Y(n_270)
);

OAI21xp5_ASAP7_75t_SL g285 ( 
.A1(n_270),
.A2(n_18),
.B(n_28),
.Y(n_285)
);

OAI22xp5_ASAP7_75t_SL g274 ( 
.A1(n_272),
.A2(n_237),
.B1(n_262),
.B2(n_240),
.Y(n_274)
);

AOI22xp5_ASAP7_75t_L g298 ( 
.A1(n_274),
.A2(n_279),
.B1(n_4),
.B2(n_5),
.Y(n_298)
);

OAI22xp5_ASAP7_75t_L g291 ( 
.A1(n_275),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_291)
);

AOI21xp5_ASAP7_75t_L g289 ( 
.A1(n_276),
.A2(n_281),
.B(n_285),
.Y(n_289)
);

BUFx12_ASAP7_75t_L g277 ( 
.A(n_258),
.Y(n_277)
);

NAND2xp5_ASAP7_75t_L g295 ( 
.A(n_277),
.B(n_2),
.Y(n_295)
);

AOI321xp33_ASAP7_75t_L g278 ( 
.A1(n_256),
.A2(n_239),
.A3(n_236),
.B1(n_9),
.B2(n_10),
.C(n_12),
.Y(n_278)
);

XNOR2xp5_ASAP7_75t_L g288 ( 
.A(n_278),
.B(n_268),
.Y(n_288)
);

OAI22xp5_ASAP7_75t_SL g279 ( 
.A1(n_256),
.A2(n_239),
.B1(n_8),
.B2(n_9),
.Y(n_279)
);

NAND3xp33_ASAP7_75t_L g280 ( 
.A(n_265),
.B(n_12),
.C(n_10),
.Y(n_280)
);

AO21x1_ASAP7_75t_L g299 ( 
.A1(n_280),
.A2(n_277),
.B(n_6),
.Y(n_299)
);

OAI21xp5_ASAP7_75t_L g281 ( 
.A1(n_267),
.A2(n_18),
.B(n_8),
.Y(n_281)
);

HB1xp67_ASAP7_75t_L g283 ( 
.A(n_261),
.Y(n_283)
);

CKINVDCx16_ASAP7_75t_R g292 ( 
.A(n_283),
.Y(n_292)
);

OAI21xp5_ASAP7_75t_L g287 ( 
.A1(n_269),
.A2(n_0),
.B(n_1),
.Y(n_287)
);

AOI21xp5_ASAP7_75t_L g290 ( 
.A1(n_287),
.A2(n_0),
.B(n_1),
.Y(n_290)
);

NAND2xp5_ASAP7_75t_SL g301 ( 
.A(n_288),
.B(n_291),
.Y(n_301)
);

NOR2xp33_ASAP7_75t_SL g300 ( 
.A(n_290),
.B(n_299),
.Y(n_300)
);

NAND2xp5_ASAP7_75t_SL g293 ( 
.A(n_284),
.B(n_28),
.Y(n_293)
);

NAND2xp5_ASAP7_75t_L g303 ( 
.A(n_293),
.B(n_277),
.Y(n_303)
);

AOI21xp5_ASAP7_75t_L g294 ( 
.A1(n_282),
.A2(n_2),
.B(n_3),
.Y(n_294)
);

AOI21xp5_ASAP7_75t_L g307 ( 
.A1(n_294),
.A2(n_286),
.B(n_6),
.Y(n_307)
);

CKINVDCx16_ASAP7_75t_R g305 ( 
.A(n_295),
.Y(n_305)
);

MAJIxp5_ASAP7_75t_L g296 ( 
.A(n_276),
.B(n_3),
.C(n_4),
.Y(n_296)
);

MAJIxp5_ASAP7_75t_L g304 ( 
.A(n_296),
.B(n_297),
.C(n_273),
.Y(n_304)
);

MAJIxp5_ASAP7_75t_L g297 ( 
.A(n_273),
.B(n_3),
.C(n_4),
.Y(n_297)
);

XNOR2xp5_ASAP7_75t_SL g302 ( 
.A(n_298),
.B(n_280),
.Y(n_302)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_302),
.Y(n_311)
);

NOR2xp33_ASAP7_75t_L g314 ( 
.A(n_303),
.B(n_304),
.Y(n_314)
);

XOR2xp5_ASAP7_75t_L g306 ( 
.A(n_289),
.B(n_286),
.Y(n_306)
);

MAJIxp5_ASAP7_75t_L g309 ( 
.A(n_306),
.B(n_296),
.C(n_292),
.Y(n_309)
);

OAI21xp5_ASAP7_75t_SL g313 ( 
.A1(n_307),
.A2(n_308),
.B(n_5),
.Y(n_313)
);

AOI21xp5_ASAP7_75t_L g308 ( 
.A1(n_297),
.A2(n_5),
.B(n_6),
.Y(n_308)
);

NAND2xp5_ASAP7_75t_L g316 ( 
.A(n_309),
.B(n_313),
.Y(n_316)
);

NOR2xp67_ASAP7_75t_SL g310 ( 
.A(n_301),
.B(n_288),
.Y(n_310)
);

OAI21xp5_ASAP7_75t_SL g315 ( 
.A1(n_310),
.A2(n_305),
.B(n_6),
.Y(n_315)
);

OR2x2_ASAP7_75t_L g312 ( 
.A(n_300),
.B(n_299),
.Y(n_312)
);

NOR2xp33_ASAP7_75t_SL g317 ( 
.A(n_312),
.B(n_314),
.Y(n_317)
);

NAND2xp5_ASAP7_75t_L g318 ( 
.A(n_315),
.B(n_317),
.Y(n_318)
);

AO21x1_ASAP7_75t_L g319 ( 
.A1(n_318),
.A2(n_311),
.B(n_316),
.Y(n_319)
);

CKINVDCx20_ASAP7_75t_R g320 ( 
.A(n_319),
.Y(n_320)
);

INVxp67_ASAP7_75t_L g321 ( 
.A(n_320),
.Y(n_321)
);

MAJIxp5_ASAP7_75t_L g322 ( 
.A(n_321),
.B(n_305),
.C(n_21),
.Y(n_322)
);

OAI21xp5_ASAP7_75t_SL g323 ( 
.A1(n_322),
.A2(n_21),
.B(n_28),
.Y(n_323)
);

XNOR2xp5_ASAP7_75t_L g324 ( 
.A(n_323),
.B(n_21),
.Y(n_324)
);

AOI21xp5_ASAP7_75t_L g325 ( 
.A1(n_324),
.A2(n_21),
.B(n_28),
.Y(n_325)
);


endmodule