module real_jpeg_23657_n_16 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_3, n_10, n_9, n_16);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_16;

wire n_108;
wire n_54;
wire n_37;
wire n_168;
wire n_73;
wire n_35;
wire n_38;
wire n_29;
wire n_91;
wire n_49;
wire n_114;
wire n_201;
wire n_68;
wire n_146;
wire n_78;
wire n_83;
wire n_166;
wire n_176;
wire n_104;
wire n_153;
wire n_194;
wire n_161;
wire n_207;
wire n_64;
wire n_177;
wire n_47;
wire n_131;
wire n_163;
wire n_22;
wire n_174;
wire n_87;
wire n_197;
wire n_40;
wire n_105;
wire n_173;
wire n_115;
wire n_98;
wire n_27;
wire n_184;
wire n_56;
wire n_48;
wire n_164;
wire n_200;
wire n_140;
wire n_126;
wire n_214;
wire n_113;
wire n_120;
wire n_155;
wire n_199;
wire n_93;
wire n_95;
wire n_141;
wire n_65;
wire n_33;
wire n_139;
wire n_188;
wire n_142;
wire n_175;
wire n_76;
wire n_178;
wire n_67;
wire n_79;
wire n_107;
wire n_156;
wire n_147;
wire n_189;
wire n_170;
wire n_66;
wire n_136;
wire n_28;
wire n_44;
wire n_208;
wire n_62;
wire n_162;
wire n_121;
wire n_106;
wire n_172;
wire n_211;
wire n_160;
wire n_45;
wire n_112;
wire n_42;
wire n_18;
wire n_145;
wire n_77;
wire n_109;
wire n_39;
wire n_122;
wire n_94;
wire n_26;
wire n_19;
wire n_148;
wire n_118;
wire n_17;
wire n_123;
wire n_116;
wire n_21;
wire n_50;
wire n_143;
wire n_196;
wire n_69;
wire n_186;
wire n_31;
wire n_137;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_165;
wire n_134;
wire n_72;
wire n_159;
wire n_171;
wire n_151;
wire n_183;
wire n_203;
wire n_192;
wire n_100;
wire n_198;
wire n_23;
wire n_51;
wire n_71;
wire n_90;
wire n_61;
wire n_110;
wire n_195;
wire n_205;
wire n_117;
wire n_99;
wire n_193;
wire n_86;
wire n_70;
wire n_41;
wire n_74;
wire n_80;
wire n_32;
wire n_20;
wire n_150;
wire n_30;
wire n_158;
wire n_204;
wire n_149;
wire n_144;
wire n_130;
wire n_103;
wire n_43;
wire n_57;
wire n_157;
wire n_84;
wire n_212;
wire n_82;
wire n_111;
wire n_132;
wire n_125;
wire n_185;
wire n_55;
wire n_209;
wire n_180;
wire n_58;
wire n_52;
wire n_191;
wire n_63;
wire n_124;
wire n_24;
wire n_92;
wire n_97;
wire n_75;
wire n_187;
wire n_34;
wire n_190;
wire n_60;
wire n_46;
wire n_169;
wire n_88;
wire n_59;
wire n_128;
wire n_167;
wire n_202;
wire n_179;
wire n_213;
wire n_133;
wire n_138;
wire n_25;
wire n_53;
wire n_127;
wire n_210;
wire n_206;
wire n_119;
wire n_36;
wire n_81;
wire n_102;
wire n_181;
wire n_85;
wire n_101;
wire n_182;
wire n_96;
wire n_89;

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_0),
.Y(n_28)
);

OAI22xp33_ASAP7_75t_SL g60 ( 
.A1(n_1),
.A2(n_27),
.B1(n_35),
.B2(n_61),
.Y(n_60)
);

CKINVDCx20_ASAP7_75t_R g61 ( 
.A(n_1),
.Y(n_61)
);

AOI22xp33_ASAP7_75t_L g72 ( 
.A1(n_1),
.A2(n_31),
.B1(n_61),
.B2(n_73),
.Y(n_72)
);

OAI22xp5_ASAP7_75t_SL g103 ( 
.A1(n_1),
.A2(n_51),
.B1(n_52),
.B2(n_61),
.Y(n_103)
);

OAI22xp5_ASAP7_75t_L g152 ( 
.A1(n_1),
.A2(n_38),
.B1(n_39),
.B2(n_61),
.Y(n_152)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_2),
.Y(n_30)
);

NAND2xp5_ASAP7_75t_L g125 ( 
.A(n_2),
.B(n_69),
.Y(n_125)
);

O2A1O1Ixp33_ASAP7_75t_L g148 ( 
.A1(n_2),
.A2(n_35),
.B(n_53),
.C(n_149),
.Y(n_148)
);

AOI22xp33_ASAP7_75t_L g161 ( 
.A1(n_2),
.A2(n_27),
.B1(n_30),
.B2(n_35),
.Y(n_161)
);

MAJIxp5_ASAP7_75t_L g169 ( 
.A(n_2),
.B(n_39),
.C(n_94),
.Y(n_169)
);

AOI22xp33_ASAP7_75t_L g172 ( 
.A1(n_2),
.A2(n_30),
.B1(n_51),
.B2(n_52),
.Y(n_172)
);

OAI21xp5_ASAP7_75t_SL g183 ( 
.A1(n_2),
.A2(n_81),
.B(n_184),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_L g195 ( 
.A(n_2),
.B(n_62),
.Y(n_195)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_3),
.Y(n_40)
);

BUFx12f_ASAP7_75t_L g95 ( 
.A(n_4),
.Y(n_95)
);

INVx8_ASAP7_75t_SL g26 ( 
.A(n_5),
.Y(n_26)
);

AOI22xp33_ASAP7_75t_SL g89 ( 
.A1(n_6),
.A2(n_51),
.B1(n_52),
.B2(n_90),
.Y(n_89)
);

CKINVDCx20_ASAP7_75t_R g90 ( 
.A(n_6),
.Y(n_90)
);

AOI22xp33_ASAP7_75t_L g127 ( 
.A1(n_6),
.A2(n_38),
.B1(n_39),
.B2(n_90),
.Y(n_127)
);

OAI22xp5_ASAP7_75t_L g65 ( 
.A1(n_7),
.A2(n_32),
.B1(n_66),
.B2(n_67),
.Y(n_65)
);

CKINVDCx20_ASAP7_75t_R g66 ( 
.A(n_7),
.Y(n_66)
);

OAI22xp5_ASAP7_75t_L g105 ( 
.A1(n_7),
.A2(n_27),
.B1(n_35),
.B2(n_66),
.Y(n_105)
);

AOI22xp33_ASAP7_75t_L g158 ( 
.A1(n_7),
.A2(n_51),
.B1(n_52),
.B2(n_66),
.Y(n_158)
);

AOI22xp5_ASAP7_75t_L g175 ( 
.A1(n_7),
.A2(n_38),
.B1(n_39),
.B2(n_66),
.Y(n_175)
);

BUFx5_ASAP7_75t_L g53 ( 
.A(n_8),
.Y(n_53)
);

OAI22xp5_ASAP7_75t_L g57 ( 
.A1(n_9),
.A2(n_27),
.B1(n_35),
.B2(n_58),
.Y(n_57)
);

CKINVDCx16_ASAP7_75t_R g58 ( 
.A(n_9),
.Y(n_58)
);

OAI22xp5_ASAP7_75t_L g143 ( 
.A1(n_9),
.A2(n_51),
.B1(n_52),
.B2(n_58),
.Y(n_143)
);

AOI22xp33_ASAP7_75t_L g177 ( 
.A1(n_9),
.A2(n_38),
.B1(n_39),
.B2(n_58),
.Y(n_177)
);

INVx13_ASAP7_75t_L g32 ( 
.A(n_10),
.Y(n_32)
);

AOI22xp5_ASAP7_75t_L g44 ( 
.A1(n_11),
.A2(n_38),
.B1(n_39),
.B2(n_45),
.Y(n_44)
);

CKINVDCx14_ASAP7_75t_R g45 ( 
.A(n_11),
.Y(n_45)
);

AOI22xp33_ASAP7_75t_L g98 ( 
.A1(n_11),
.A2(n_45),
.B1(n_51),
.B2(n_52),
.Y(n_98)
);

AOI22xp33_ASAP7_75t_SL g86 ( 
.A1(n_12),
.A2(n_38),
.B1(n_39),
.B2(n_87),
.Y(n_86)
);

CKINVDCx20_ASAP7_75t_R g87 ( 
.A(n_12),
.Y(n_87)
);

OAI22xp5_ASAP7_75t_L g46 ( 
.A1(n_13),
.A2(n_38),
.B1(n_39),
.B2(n_47),
.Y(n_46)
);

CKINVDCx16_ASAP7_75t_R g47 ( 
.A(n_13),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_14),
.Y(n_52)
);

AOI22xp5_ASAP7_75t_L g36 ( 
.A1(n_15),
.A2(n_37),
.B1(n_43),
.B2(n_46),
.Y(n_36)
);

INVx6_ASAP7_75t_L g42 ( 
.A(n_15),
.Y(n_42)
);

INVx6_ASAP7_75t_L g85 ( 
.A(n_15),
.Y(n_85)
);

INVx2_ASAP7_75t_L g128 ( 
.A(n_15),
.Y(n_128)
);

AOI22xp5_ASAP7_75t_L g173 ( 
.A1(n_15),
.A2(n_37),
.B1(n_174),
.B2(n_176),
.Y(n_173)
);

INVx3_ASAP7_75t_L g182 ( 
.A(n_15),
.Y(n_182)
);

XNOR2xp5_ASAP7_75t_L g16 ( 
.A(n_17),
.B(n_131),
.Y(n_16)
);

NAND2xp5_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_129),
.Y(n_17)
);

INVxp67_ASAP7_75t_L g18 ( 
.A(n_19),
.Y(n_18)
);

NOR2xp33_ASAP7_75t_SL g19 ( 
.A(n_20),
.B(n_112),
.Y(n_19)
);

AND2x2_ASAP7_75t_L g130 ( 
.A(n_20),
.B(n_112),
.Y(n_130)
);

OAI22xp5_ASAP7_75t_L g20 ( 
.A1(n_21),
.A2(n_77),
.B1(n_78),
.B2(n_111),
.Y(n_20)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_21),
.Y(n_111)
);

BUFx24_ASAP7_75t_SL g216 ( 
.A(n_21),
.Y(n_216)
);

FAx1_ASAP7_75t_SL g21 ( 
.A(n_22),
.B(n_48),
.CI(n_63),
.CON(n_21),
.SN(n_21)
);

NOR2xp33_ASAP7_75t_L g22 ( 
.A(n_23),
.B(n_36),
.Y(n_22)
);

OAI22xp5_ASAP7_75t_L g118 ( 
.A1(n_23),
.A2(n_24),
.B1(n_36),
.B2(n_119),
.Y(n_118)
);

CKINVDCx14_ASAP7_75t_R g23 ( 
.A(n_24),
.Y(n_23)
);

A2O1A1Ixp33_ASAP7_75t_L g24 ( 
.A1(n_25),
.A2(n_27),
.B(n_29),
.C(n_33),
.Y(n_24)
);

OAI22xp5_ASAP7_75t_L g69 ( 
.A1(n_25),
.A2(n_26),
.B1(n_27),
.B2(n_35),
.Y(n_69)
);

OAI22xp33_ASAP7_75t_L g76 ( 
.A1(n_25),
.A2(n_26),
.B1(n_32),
.B2(n_74),
.Y(n_76)
);

INVx8_ASAP7_75t_L g25 ( 
.A(n_26),
.Y(n_25)
);

NAND3xp33_ASAP7_75t_SL g33 ( 
.A(n_26),
.B(n_34),
.C(n_35),
.Y(n_33)
);

INVx5_ASAP7_75t_SL g35 ( 
.A(n_27),
.Y(n_35)
);

OAI22xp5_ASAP7_75t_L g55 ( 
.A1(n_27),
.A2(n_35),
.B1(n_53),
.B2(n_54),
.Y(n_55)
);

BUFx12f_ASAP7_75t_L g27 ( 
.A(n_28),
.Y(n_27)
);

OAI21xp33_ASAP7_75t_L g108 ( 
.A1(n_29),
.A2(n_30),
.B(n_109),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_SL g29 ( 
.A(n_30),
.B(n_31),
.Y(n_29)
);

OAI21xp33_ASAP7_75t_L g149 ( 
.A1(n_30),
.A2(n_51),
.B(n_54),
.Y(n_149)
);

NOR2xp33_ASAP7_75t_SL g181 ( 
.A(n_30),
.B(n_182),
.Y(n_181)
);

NOR2xp33_ASAP7_75t_L g188 ( 
.A(n_30),
.B(n_97),
.Y(n_188)
);

INVx11_ASAP7_75t_L g31 ( 
.A(n_32),
.Y(n_31)
);

INVx8_ASAP7_75t_L g34 ( 
.A(n_32),
.Y(n_34)
);

INVx8_ASAP7_75t_L g67 ( 
.A(n_32),
.Y(n_67)
);

INVx6_ASAP7_75t_L g74 ( 
.A(n_32),
.Y(n_74)
);

CKINVDCx14_ASAP7_75t_R g119 ( 
.A(n_36),
.Y(n_119)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_37),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g151 ( 
.A(n_37),
.B(n_152),
.Y(n_151)
);

NOR2xp33_ASAP7_75t_L g37 ( 
.A(n_38),
.B(n_41),
.Y(n_37)
);

OA22x2_ASAP7_75t_L g97 ( 
.A1(n_38),
.A2(n_39),
.B1(n_94),
.B2(n_96),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g180 ( 
.A(n_38),
.B(n_181),
.Y(n_180)
);

INVx6_ASAP7_75t_SL g38 ( 
.A(n_39),
.Y(n_38)
);

BUFx12f_ASAP7_75t_L g39 ( 
.A(n_40),
.Y(n_39)
);

INVx8_ASAP7_75t_L g41 ( 
.A(n_42),
.Y(n_41)
);

INVxp67_ASAP7_75t_L g43 ( 
.A(n_44),
.Y(n_43)
);

OAI22xp5_ASAP7_75t_SL g126 ( 
.A1(n_44),
.A2(n_81),
.B1(n_127),
.B2(n_128),
.Y(n_126)
);

INVxp67_ASAP7_75t_L g82 ( 
.A(n_46),
.Y(n_82)
);

OAI21xp5_ASAP7_75t_SL g48 ( 
.A1(n_49),
.A2(n_56),
.B(n_59),
.Y(n_48)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_49),
.Y(n_106)
);

OAI21xp33_ASAP7_75t_L g160 ( 
.A1(n_49),
.A2(n_59),
.B(n_161),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_L g49 ( 
.A(n_50),
.B(n_55),
.Y(n_49)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_50),
.Y(n_62)
);

OAI21xp5_ASAP7_75t_SL g121 ( 
.A1(n_50),
.A2(n_122),
.B(n_123),
.Y(n_121)
);

AOI22xp5_ASAP7_75t_SL g50 ( 
.A1(n_51),
.A2(n_52),
.B1(n_53),
.B2(n_54),
.Y(n_50)
);

OAI22xp33_ASAP7_75t_L g93 ( 
.A1(n_51),
.A2(n_52),
.B1(n_94),
.B2(n_96),
.Y(n_93)
);

INVx1_ASAP7_75t_SL g51 ( 
.A(n_52),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_L g168 ( 
.A(n_52),
.B(n_169),
.Y(n_168)
);

INVx2_ASAP7_75t_L g54 ( 
.A(n_53),
.Y(n_54)
);

CKINVDCx14_ASAP7_75t_R g56 ( 
.A(n_57),
.Y(n_56)
);

AOI22xp5_ASAP7_75t_L g104 ( 
.A1(n_57),
.A2(n_62),
.B1(n_105),
.B2(n_106),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_SL g59 ( 
.A(n_60),
.B(n_62),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_L g123 ( 
.A(n_60),
.B(n_106),
.Y(n_123)
);

OAI21xp5_ASAP7_75t_L g63 ( 
.A1(n_64),
.A2(n_68),
.B(n_70),
.Y(n_63)
);

CKINVDCx20_ASAP7_75t_R g64 ( 
.A(n_65),
.Y(n_64)
);

AND2x2_ASAP7_75t_L g75 ( 
.A(n_68),
.B(n_76),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_68),
.B(n_72),
.Y(n_110)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_69),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_L g70 ( 
.A(n_71),
.B(n_75),
.Y(n_70)
);

CKINVDCx14_ASAP7_75t_R g71 ( 
.A(n_72),
.Y(n_71)
);

INVx8_ASAP7_75t_L g109 ( 
.A(n_73),
.Y(n_109)
);

INVx8_ASAP7_75t_L g73 ( 
.A(n_74),
.Y(n_73)
);

AOI21xp5_ASAP7_75t_L g107 ( 
.A1(n_75),
.A2(n_108),
.B(n_110),
.Y(n_107)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_78),
.Y(n_77)
);

XNOR2xp5_ASAP7_75t_SL g78 ( 
.A(n_79),
.B(n_99),
.Y(n_78)
);

XOR2xp5_ASAP7_75t_L g79 ( 
.A(n_80),
.B(n_88),
.Y(n_79)
);

OAI22xp5_ASAP7_75t_L g80 ( 
.A1(n_81),
.A2(n_82),
.B1(n_83),
.B2(n_86),
.Y(n_80)
);

OAI21xp5_ASAP7_75t_L g198 ( 
.A1(n_81),
.A2(n_177),
.B(n_184),
.Y(n_198)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_84),
.Y(n_83)
);

INVx2_ASAP7_75t_L g84 ( 
.A(n_85),
.Y(n_84)
);

OAI22xp5_ASAP7_75t_L g88 ( 
.A1(n_89),
.A2(n_91),
.B1(n_97),
.B2(n_98),
.Y(n_88)
);

OAI21xp5_ASAP7_75t_L g101 ( 
.A1(n_89),
.A2(n_97),
.B(n_102),
.Y(n_101)
);

OAI21xp5_ASAP7_75t_SL g141 ( 
.A1(n_91),
.A2(n_142),
.B(n_144),
.Y(n_141)
);

OAI21xp5_ASAP7_75t_SL g171 ( 
.A1(n_91),
.A2(n_144),
.B(n_172),
.Y(n_171)
);

CKINVDCx20_ASAP7_75t_R g91 ( 
.A(n_92),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_SL g102 ( 
.A(n_92),
.B(n_103),
.Y(n_102)
);

AOI22xp5_ASAP7_75t_L g156 ( 
.A1(n_92),
.A2(n_143),
.B1(n_145),
.B2(n_157),
.Y(n_156)
);

AND2x2_ASAP7_75t_L g92 ( 
.A(n_93),
.B(n_97),
.Y(n_92)
);

INVx13_ASAP7_75t_L g96 ( 
.A(n_94),
.Y(n_96)
);

BUFx24_ASAP7_75t_L g94 ( 
.A(n_95),
.Y(n_94)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_97),
.Y(n_145)
);

OAI21xp5_ASAP7_75t_L g197 ( 
.A1(n_97),
.A2(n_102),
.B(n_158),
.Y(n_197)
);

MAJIxp5_ASAP7_75t_L g99 ( 
.A(n_100),
.B(n_104),
.C(n_107),
.Y(n_99)
);

AOI22xp5_ASAP7_75t_L g115 ( 
.A1(n_100),
.A2(n_101),
.B1(n_104),
.B2(n_116),
.Y(n_115)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_101),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_SL g144 ( 
.A(n_103),
.B(n_145),
.Y(n_144)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_104),
.Y(n_116)
);

CKINVDCx16_ASAP7_75t_R g122 ( 
.A(n_105),
.Y(n_122)
);

XOR2xp5_ASAP7_75t_L g114 ( 
.A(n_107),
.B(n_115),
.Y(n_114)
);

MAJIxp5_ASAP7_75t_L g112 ( 
.A(n_113),
.B(n_117),
.C(n_120),
.Y(n_112)
);

AOI22xp5_ASAP7_75t_L g209 ( 
.A1(n_113),
.A2(n_114),
.B1(n_210),
.B2(n_211),
.Y(n_209)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_114),
.Y(n_113)
);

AOI22xp5_ASAP7_75t_L g211 ( 
.A1(n_117),
.A2(n_118),
.B1(n_120),
.B2(n_212),
.Y(n_211)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_118),
.Y(n_117)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_120),
.Y(n_212)
);

MAJIxp5_ASAP7_75t_L g120 ( 
.A(n_121),
.B(n_124),
.C(n_126),
.Y(n_120)
);

XOR2xp5_ASAP7_75t_L g136 ( 
.A(n_121),
.B(n_137),
.Y(n_136)
);

AOI22xp5_ASAP7_75t_L g137 ( 
.A1(n_124),
.A2(n_125),
.B1(n_126),
.B2(n_138),
.Y(n_137)
);

CKINVDCx20_ASAP7_75t_R g124 ( 
.A(n_125),
.Y(n_124)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_126),
.Y(n_138)
);

OAI21xp5_ASAP7_75t_L g150 ( 
.A1(n_127),
.A2(n_128),
.B(n_151),
.Y(n_150)
);

CKINVDCx20_ASAP7_75t_R g129 ( 
.A(n_130),
.Y(n_129)
);

AOI21xp5_ASAP7_75t_SL g131 ( 
.A1(n_132),
.A2(n_208),
.B(n_214),
.Y(n_131)
);

OAI21xp5_ASAP7_75t_L g132 ( 
.A1(n_133),
.A2(n_162),
.B(n_207),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_SL g133 ( 
.A(n_134),
.B(n_154),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_L g207 ( 
.A(n_134),
.B(n_154),
.Y(n_207)
);

OAI22xp5_ASAP7_75t_SL g134 ( 
.A1(n_135),
.A2(n_136),
.B1(n_139),
.B2(n_153),
.Y(n_134)
);

MAJIxp5_ASAP7_75t_L g213 ( 
.A(n_135),
.B(n_141),
.C(n_146),
.Y(n_213)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_136),
.Y(n_135)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_139),
.Y(n_153)
);

AOI22xp5_ASAP7_75t_L g139 ( 
.A1(n_140),
.A2(n_141),
.B1(n_146),
.B2(n_147),
.Y(n_139)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_141),
.Y(n_140)
);

CKINVDCx20_ASAP7_75t_R g142 ( 
.A(n_143),
.Y(n_142)
);

CKINVDCx16_ASAP7_75t_R g146 ( 
.A(n_147),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_L g147 ( 
.A(n_148),
.B(n_150),
.Y(n_147)
);

XNOR2xp5_ASAP7_75t_SL g155 ( 
.A(n_148),
.B(n_150),
.Y(n_155)
);

OAI21xp5_ASAP7_75t_L g187 ( 
.A1(n_151),
.A2(n_175),
.B(n_182),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_L g184 ( 
.A(n_152),
.B(n_185),
.Y(n_184)
);

MAJIxp5_ASAP7_75t_L g154 ( 
.A(n_155),
.B(n_156),
.C(n_159),
.Y(n_154)
);

XNOR2xp5_ASAP7_75t_L g202 ( 
.A(n_155),
.B(n_203),
.Y(n_202)
);

AOI22xp5_ASAP7_75t_L g203 ( 
.A1(n_156),
.A2(n_159),
.B1(n_160),
.B2(n_204),
.Y(n_203)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_156),
.Y(n_204)
);

INVxp67_ASAP7_75t_L g157 ( 
.A(n_158),
.Y(n_157)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_160),
.Y(n_159)
);

AOI21xp5_ASAP7_75t_L g162 ( 
.A1(n_163),
.A2(n_201),
.B(n_206),
.Y(n_162)
);

OAI21xp5_ASAP7_75t_L g163 ( 
.A1(n_164),
.A2(n_191),
.B(n_200),
.Y(n_163)
);

AOI21xp5_ASAP7_75t_L g164 ( 
.A1(n_165),
.A2(n_178),
.B(n_190),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_SL g165 ( 
.A(n_166),
.B(n_173),
.Y(n_165)
);

NOR2xp33_ASAP7_75t_L g190 ( 
.A(n_166),
.B(n_173),
.Y(n_190)
);

AOI22xp5_ASAP7_75t_L g166 ( 
.A1(n_167),
.A2(n_168),
.B1(n_170),
.B2(n_171),
.Y(n_166)
);

CKINVDCx20_ASAP7_75t_R g167 ( 
.A(n_168),
.Y(n_167)
);

NOR2xp33_ASAP7_75t_L g199 ( 
.A(n_168),
.B(n_170),
.Y(n_199)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_171),
.Y(n_170)
);

CKINVDCx16_ASAP7_75t_R g174 ( 
.A(n_175),
.Y(n_174)
);

INVxp67_ASAP7_75t_L g176 ( 
.A(n_177),
.Y(n_176)
);

OAI21xp5_ASAP7_75t_L g178 ( 
.A1(n_179),
.A2(n_186),
.B(n_189),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_L g179 ( 
.A(n_180),
.B(n_183),
.Y(n_179)
);

INVx3_ASAP7_75t_L g185 ( 
.A(n_182),
.Y(n_185)
);

NOR2xp33_ASAP7_75t_SL g186 ( 
.A(n_187),
.B(n_188),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_L g189 ( 
.A(n_187),
.B(n_188),
.Y(n_189)
);

NOR2xp33_ASAP7_75t_SL g191 ( 
.A(n_192),
.B(n_199),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_L g200 ( 
.A(n_192),
.B(n_199),
.Y(n_200)
);

XNOR2xp5_ASAP7_75t_L g192 ( 
.A(n_193),
.B(n_198),
.Y(n_192)
);

AOI22xp5_ASAP7_75t_L g193 ( 
.A1(n_194),
.A2(n_195),
.B1(n_196),
.B2(n_197),
.Y(n_193)
);

MAJIxp5_ASAP7_75t_L g205 ( 
.A(n_194),
.B(n_197),
.C(n_198),
.Y(n_205)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_195),
.Y(n_194)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_197),
.Y(n_196)
);

NAND2xp5_ASAP7_75t_SL g201 ( 
.A(n_202),
.B(n_205),
.Y(n_201)
);

NOR2xp33_ASAP7_75t_L g206 ( 
.A(n_202),
.B(n_205),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_SL g208 ( 
.A(n_209),
.B(n_213),
.Y(n_208)
);

NOR2xp33_ASAP7_75t_L g214 ( 
.A(n_209),
.B(n_213),
.Y(n_214)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_211),
.Y(n_210)
);


endmodule