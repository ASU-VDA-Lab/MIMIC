module fake_jpeg_22508_n_272 (n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_272);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_272;

wire n_159;
wire n_117;
wire n_253;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_14;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_251;
wire n_252;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_154;
wire n_127;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_13;
wire n_175;
wire n_187;
wire n_57;
wire n_21;
wire n_223;
wire n_234;
wire n_171;
wire n_263;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_267;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_24;
wire n_44;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_269;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_128;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_266;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_262;
wire n_212;
wire n_131;
wire n_56;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_271;
wire n_216;
wire n_217;
wire n_264;
wire n_184;
wire n_53;
wire n_268;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_265;
wire n_176;
wire n_199;
wire n_112;
wire n_260;
wire n_270;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_140;
wire n_258;
wire n_96;

CKINVDCx20_ASAP7_75t_R g13 ( 
.A(n_5),
.Y(n_13)
);

INVx6_ASAP7_75t_L g14 ( 
.A(n_3),
.Y(n_14)
);

BUFx5_ASAP7_75t_L g15 ( 
.A(n_3),
.Y(n_15)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_5),
.Y(n_16)
);

BUFx12f_ASAP7_75t_L g17 ( 
.A(n_4),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_9),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_12),
.Y(n_19)
);

BUFx5_ASAP7_75t_L g20 ( 
.A(n_4),
.Y(n_20)
);

BUFx10_ASAP7_75t_L g21 ( 
.A(n_6),
.Y(n_21)
);

INVx11_ASAP7_75t_L g22 ( 
.A(n_2),
.Y(n_22)
);

INVx13_ASAP7_75t_L g23 ( 
.A(n_10),
.Y(n_23)
);

NOR2xp33_ASAP7_75t_L g24 ( 
.A(n_5),
.B(n_7),
.Y(n_24)
);

BUFx12_ASAP7_75t_L g25 ( 
.A(n_9),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_12),
.Y(n_26)
);

INVx3_ASAP7_75t_L g27 ( 
.A(n_12),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_17),
.Y(n_28)
);

NOR2xp33_ASAP7_75t_L g41 ( 
.A(n_28),
.B(n_30),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g29 ( 
.A(n_24),
.B(n_6),
.Y(n_29)
);

NOR2xp33_ASAP7_75t_SL g48 ( 
.A(n_29),
.B(n_34),
.Y(n_48)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_17),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_13),
.Y(n_31)
);

NOR2xp33_ASAP7_75t_L g43 ( 
.A(n_31),
.B(n_36),
.Y(n_43)
);

INVx2_ASAP7_75t_L g32 ( 
.A(n_25),
.Y(n_32)
);

INVx6_ASAP7_75t_L g49 ( 
.A(n_32),
.Y(n_49)
);

INVx4_ASAP7_75t_L g33 ( 
.A(n_23),
.Y(n_33)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_33),
.Y(n_44)
);

AND2x2_ASAP7_75t_L g34 ( 
.A(n_23),
.B(n_17),
.Y(n_34)
);

BUFx12f_ASAP7_75t_L g35 ( 
.A(n_17),
.Y(n_35)
);

BUFx3_ASAP7_75t_L g50 ( 
.A(n_35),
.Y(n_50)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_17),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_13),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g51 ( 
.A(n_37),
.B(n_13),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_L g38 ( 
.A(n_34),
.B(n_14),
.Y(n_38)
);

NAND2xp5_ASAP7_75t_L g60 ( 
.A(n_38),
.B(n_55),
.Y(n_60)
);

INVx2_ASAP7_75t_L g39 ( 
.A(n_35),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_39),
.B(n_42),
.Y(n_56)
);

AOI22xp33_ASAP7_75t_L g40 ( 
.A1(n_34),
.A2(n_14),
.B1(n_23),
.B2(n_22),
.Y(n_40)
);

AOI22xp5_ASAP7_75t_SL g59 ( 
.A1(n_40),
.A2(n_27),
.B1(n_15),
.B2(n_20),
.Y(n_59)
);

INVxp67_ASAP7_75t_L g42 ( 
.A(n_35),
.Y(n_42)
);

INVx3_ASAP7_75t_L g45 ( 
.A(n_35),
.Y(n_45)
);

INVx3_ASAP7_75t_SL g71 ( 
.A(n_45),
.Y(n_71)
);

AOI22xp33_ASAP7_75t_SL g46 ( 
.A1(n_35),
.A2(n_14),
.B1(n_27),
.B2(n_22),
.Y(n_46)
);

AOI21xp5_ASAP7_75t_L g70 ( 
.A1(n_46),
.A2(n_47),
.B(n_17),
.Y(n_70)
);

AOI22xp33_ASAP7_75t_SL g47 ( 
.A1(n_28),
.A2(n_14),
.B1(n_27),
.B2(n_22),
.Y(n_47)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_51),
.Y(n_58)
);

INVx2_ASAP7_75t_L g52 ( 
.A(n_32),
.Y(n_52)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_52),
.Y(n_61)
);

INVx3_ASAP7_75t_L g53 ( 
.A(n_33),
.Y(n_53)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_53),
.Y(n_66)
);

CKINVDCx14_ASAP7_75t_SL g54 ( 
.A(n_33),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_54),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_L g55 ( 
.A(n_34),
.B(n_16),
.Y(n_55)
);

AOI22xp33_ASAP7_75t_SL g57 ( 
.A1(n_49),
.A2(n_27),
.B1(n_22),
.B2(n_23),
.Y(n_57)
);

INVxp67_ASAP7_75t_L g82 ( 
.A(n_57),
.Y(n_82)
);

OAI22xp5_ASAP7_75t_SL g91 ( 
.A1(n_59),
.A2(n_46),
.B1(n_70),
.B2(n_32),
.Y(n_91)
);

AOI22xp33_ASAP7_75t_SL g62 ( 
.A1(n_49),
.A2(n_23),
.B1(n_18),
.B2(n_26),
.Y(n_62)
);

AOI22xp33_ASAP7_75t_SL g90 ( 
.A1(n_62),
.A2(n_70),
.B1(n_17),
.B2(n_53),
.Y(n_90)
);

INVx2_ASAP7_75t_L g63 ( 
.A(n_54),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_63),
.B(n_64),
.Y(n_87)
);

INVx2_ASAP7_75t_L g64 ( 
.A(n_50),
.Y(n_64)
);

INVx2_ASAP7_75t_L g67 ( 
.A(n_50),
.Y(n_67)
);

INVx2_ASAP7_75t_L g80 ( 
.A(n_67),
.Y(n_80)
);

INVx2_ASAP7_75t_L g68 ( 
.A(n_50),
.Y(n_68)
);

INVx3_ASAP7_75t_L g85 ( 
.A(n_68),
.Y(n_85)
);

MAJIxp5_ASAP7_75t_L g69 ( 
.A(n_38),
.B(n_30),
.C(n_36),
.Y(n_69)
);

MAJIxp5_ASAP7_75t_L g88 ( 
.A(n_69),
.B(n_55),
.C(n_48),
.Y(n_88)
);

CKINVDCx20_ASAP7_75t_R g72 ( 
.A(n_43),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_SL g97 ( 
.A(n_72),
.B(n_73),
.Y(n_97)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_43),
.Y(n_73)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_51),
.Y(n_74)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_74),
.Y(n_78)
);

INVx2_ASAP7_75t_L g75 ( 
.A(n_52),
.Y(n_75)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_75),
.Y(n_79)
);

BUFx6f_ASAP7_75t_L g76 ( 
.A(n_53),
.Y(n_76)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_76),
.Y(n_83)
);

AND2x2_ASAP7_75t_L g77 ( 
.A(n_60),
.B(n_38),
.Y(n_77)
);

OAI21xp5_ASAP7_75t_SL g116 ( 
.A1(n_77),
.A2(n_84),
.B(n_88),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_L g81 ( 
.A(n_60),
.B(n_69),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_81),
.B(n_93),
.Y(n_99)
);

OA21x2_ASAP7_75t_L g84 ( 
.A1(n_59),
.A2(n_40),
.B(n_47),
.Y(n_84)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_56),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_86),
.B(n_71),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_SL g89 ( 
.A(n_74),
.B(n_48),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_SL g100 ( 
.A(n_89),
.B(n_37),
.Y(n_100)
);

INVxp67_ASAP7_75t_L g104 ( 
.A(n_90),
.Y(n_104)
);

AOI22xp5_ASAP7_75t_L g111 ( 
.A1(n_91),
.A2(n_94),
.B1(n_96),
.B2(n_71),
.Y(n_111)
);

AOI22xp5_ASAP7_75t_L g92 ( 
.A1(n_73),
.A2(n_49),
.B1(n_52),
.B2(n_41),
.Y(n_92)
);

OAI22xp5_ASAP7_75t_SL g110 ( 
.A1(n_92),
.A2(n_63),
.B1(n_26),
.B2(n_18),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_L g93 ( 
.A(n_58),
.B(n_41),
.Y(n_93)
);

OAI22xp5_ASAP7_75t_SL g94 ( 
.A1(n_61),
.A2(n_28),
.B1(n_36),
.B2(n_45),
.Y(n_94)
);

MAJIxp5_ASAP7_75t_L g95 ( 
.A(n_61),
.B(n_44),
.C(n_39),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g101 ( 
.A(n_95),
.B(n_66),
.Y(n_101)
);

OAI22xp5_ASAP7_75t_SL g96 ( 
.A1(n_75),
.A2(n_45),
.B1(n_39),
.B2(n_44),
.Y(n_96)
);

OAI22xp33_ASAP7_75t_SL g98 ( 
.A1(n_84),
.A2(n_91),
.B1(n_78),
.B2(n_82),
.Y(n_98)
);

AOI22xp5_ASAP7_75t_L g122 ( 
.A1(n_98),
.A2(n_110),
.B1(n_114),
.B2(n_78),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_SL g125 ( 
.A(n_100),
.B(n_107),
.Y(n_125)
);

OAI21xp5_ASAP7_75t_SL g129 ( 
.A1(n_101),
.A2(n_112),
.B(n_109),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_L g102 ( 
.A(n_77),
.B(n_66),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_L g121 ( 
.A(n_102),
.B(n_109),
.Y(n_121)
);

AOI22xp33_ASAP7_75t_L g103 ( 
.A1(n_84),
.A2(n_20),
.B1(n_15),
.B2(n_76),
.Y(n_103)
);

OAI22xp5_ASAP7_75t_SL g123 ( 
.A1(n_103),
.A2(n_111),
.B1(n_92),
.B2(n_83),
.Y(n_123)
);

BUFx3_ASAP7_75t_L g105 ( 
.A(n_85),
.Y(n_105)
);

CKINVDCx16_ASAP7_75t_R g136 ( 
.A(n_105),
.Y(n_136)
);

BUFx3_ASAP7_75t_L g106 ( 
.A(n_85),
.Y(n_106)
);

CKINVDCx20_ASAP7_75t_R g126 ( 
.A(n_106),
.Y(n_126)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_87),
.Y(n_107)
);

INVx5_ASAP7_75t_L g108 ( 
.A(n_80),
.Y(n_108)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_108),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_L g109 ( 
.A(n_77),
.B(n_21),
.Y(n_109)
);

XOR2x1_ASAP7_75t_L g112 ( 
.A(n_84),
.B(n_15),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_L g113 ( 
.A(n_81),
.B(n_21),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_L g130 ( 
.A(n_113),
.B(n_86),
.Y(n_130)
);

OAI22xp5_ASAP7_75t_SL g114 ( 
.A1(n_82),
.A2(n_15),
.B1(n_20),
.B2(n_16),
.Y(n_114)
);

INVx13_ASAP7_75t_L g115 ( 
.A(n_80),
.Y(n_115)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_115),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_SL g142 ( 
.A(n_117),
.B(n_118),
.Y(n_142)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_96),
.Y(n_118)
);

INVxp67_ASAP7_75t_L g119 ( 
.A(n_95),
.Y(n_119)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_119),
.Y(n_132)
);

OAI32xp33_ASAP7_75t_L g120 ( 
.A1(n_112),
.A2(n_88),
.A3(n_93),
.B1(n_94),
.B2(n_89),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_L g157 ( 
.A(n_120),
.B(n_130),
.Y(n_157)
);

OAI22xp5_ASAP7_75t_L g152 ( 
.A1(n_122),
.A2(n_131),
.B1(n_141),
.B2(n_111),
.Y(n_152)
);

AOI22xp5_ASAP7_75t_L g151 ( 
.A1(n_123),
.A2(n_140),
.B1(n_114),
.B2(n_110),
.Y(n_151)
);

XOR2xp5_ASAP7_75t_L g124 ( 
.A(n_116),
.B(n_97),
.Y(n_124)
);

MAJIxp5_ASAP7_75t_L g147 ( 
.A(n_124),
.B(n_137),
.C(n_99),
.Y(n_147)
);

XNOR2xp5_ASAP7_75t_L g144 ( 
.A(n_129),
.B(n_99),
.Y(n_144)
);

AOI22xp5_ASAP7_75t_SL g131 ( 
.A1(n_104),
.A2(n_20),
.B1(n_18),
.B2(n_26),
.Y(n_131)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_117),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_SL g146 ( 
.A(n_133),
.B(n_107),
.Y(n_146)
);

OAI21xp5_ASAP7_75t_SL g134 ( 
.A1(n_112),
.A2(n_79),
.B(n_83),
.Y(n_134)
);

XOR2xp5_ASAP7_75t_L g155 ( 
.A(n_134),
.B(n_138),
.Y(n_155)
);

AND2x2_ASAP7_75t_L g135 ( 
.A(n_102),
.B(n_101),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_L g163 ( 
.A(n_135),
.B(n_21),
.Y(n_163)
);

MAJIxp5_ASAP7_75t_L g137 ( 
.A(n_116),
.B(n_79),
.C(n_68),
.Y(n_137)
);

XNOR2xp5_ASAP7_75t_L g138 ( 
.A(n_113),
.B(n_29),
.Y(n_138)
);

CKINVDCx20_ASAP7_75t_R g139 ( 
.A(n_105),
.Y(n_139)
);

CKINVDCx20_ASAP7_75t_R g156 ( 
.A(n_139),
.Y(n_156)
);

OAI22xp5_ASAP7_75t_SL g140 ( 
.A1(n_103),
.A2(n_64),
.B1(n_67),
.B2(n_31),
.Y(n_140)
);

OAI21xp5_ASAP7_75t_SL g141 ( 
.A1(n_118),
.A2(n_16),
.B(n_21),
.Y(n_141)
);

INVx1_ASAP7_75t_SL g143 ( 
.A(n_142),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_SL g177 ( 
.A(n_143),
.B(n_150),
.Y(n_177)
);

XNOR2xp5_ASAP7_75t_SL g187 ( 
.A(n_144),
.B(n_145),
.Y(n_187)
);

XNOR2x2_ASAP7_75t_L g145 ( 
.A(n_129),
.B(n_98),
.Y(n_145)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_146),
.Y(n_178)
);

MAJIxp5_ASAP7_75t_L g172 ( 
.A(n_147),
.B(n_153),
.C(n_137),
.Y(n_172)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_130),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_L g168 ( 
.A(n_148),
.B(n_149),
.Y(n_168)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_121),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_SL g150 ( 
.A(n_125),
.B(n_100),
.Y(n_150)
);

CKINVDCx16_ASAP7_75t_R g167 ( 
.A(n_151),
.Y(n_167)
);

AOI22xp5_ASAP7_75t_L g175 ( 
.A1(n_152),
.A2(n_154),
.B1(n_123),
.B2(n_135),
.Y(n_175)
);

MAJIxp5_ASAP7_75t_L g153 ( 
.A(n_132),
.B(n_106),
.C(n_105),
.Y(n_153)
);

OAI22xp5_ASAP7_75t_SL g154 ( 
.A1(n_134),
.A2(n_121),
.B1(n_122),
.B2(n_132),
.Y(n_154)
);

CKINVDCx20_ASAP7_75t_R g158 ( 
.A(n_126),
.Y(n_158)
);

CKINVDCx20_ASAP7_75t_R g173 ( 
.A(n_158),
.Y(n_173)
);

CKINVDCx16_ASAP7_75t_R g159 ( 
.A(n_140),
.Y(n_159)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_159),
.Y(n_182)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_141),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_L g169 ( 
.A(n_160),
.B(n_162),
.Y(n_169)
);

NOR2xp33_ASAP7_75t_SL g161 ( 
.A(n_133),
.B(n_108),
.Y(n_161)
);

CKINVDCx20_ASAP7_75t_R g171 ( 
.A(n_161),
.Y(n_171)
);

AO32x1_ASAP7_75t_L g162 ( 
.A1(n_120),
.A2(n_106),
.A3(n_19),
.B1(n_108),
.B2(n_115),
.Y(n_162)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_163),
.Y(n_188)
);

INVx3_ASAP7_75t_L g164 ( 
.A(n_136),
.Y(n_164)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_164),
.Y(n_183)
);

CKINVDCx20_ASAP7_75t_R g165 ( 
.A(n_127),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_L g180 ( 
.A(n_165),
.B(n_166),
.Y(n_180)
);

CKINVDCx20_ASAP7_75t_R g166 ( 
.A(n_128),
.Y(n_166)
);

INVx2_ASAP7_75t_L g170 ( 
.A(n_164),
.Y(n_170)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_170),
.Y(n_192)
);

MAJIxp5_ASAP7_75t_L g195 ( 
.A(n_172),
.B(n_181),
.C(n_185),
.Y(n_195)
);

A2O1A1Ixp33_ASAP7_75t_L g174 ( 
.A1(n_157),
.A2(n_135),
.B(n_131),
.C(n_124),
.Y(n_174)
);

OAI21xp5_ASAP7_75t_SL g198 ( 
.A1(n_174),
.A2(n_179),
.B(n_162),
.Y(n_198)
);

NOR2xp33_ASAP7_75t_L g190 ( 
.A(n_175),
.B(n_154),
.Y(n_190)
);

HB1xp67_ASAP7_75t_L g176 ( 
.A(n_145),
.Y(n_176)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_176),
.Y(n_201)
);

AOI21xp5_ASAP7_75t_L g179 ( 
.A1(n_160),
.A2(n_128),
.B(n_115),
.Y(n_179)
);

MAJIxp5_ASAP7_75t_L g181 ( 
.A(n_147),
.B(n_138),
.C(n_24),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_L g184 ( 
.A(n_148),
.B(n_21),
.Y(n_184)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_184),
.Y(n_193)
);

MAJIxp5_ASAP7_75t_L g185 ( 
.A(n_155),
.B(n_24),
.C(n_21),
.Y(n_185)
);

OAI22xp5_ASAP7_75t_SL g186 ( 
.A1(n_157),
.A2(n_19),
.B1(n_21),
.B2(n_2),
.Y(n_186)
);

AOI22xp5_ASAP7_75t_L g194 ( 
.A1(n_186),
.A2(n_143),
.B1(n_163),
.B2(n_156),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_L g189 ( 
.A(n_171),
.B(n_149),
.Y(n_189)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_189),
.Y(n_207)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_190),
.Y(n_208)
);

CKINVDCx16_ASAP7_75t_R g191 ( 
.A(n_180),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_SL g221 ( 
.A(n_191),
.B(n_202),
.Y(n_221)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_194),
.Y(n_216)
);

MAJIxp5_ASAP7_75t_L g196 ( 
.A(n_172),
.B(n_155),
.C(n_153),
.Y(n_196)
);

MAJIxp5_ASAP7_75t_L g211 ( 
.A(n_196),
.B(n_203),
.C(n_188),
.Y(n_211)
);

XOR2xp5_ASAP7_75t_L g197 ( 
.A(n_187),
.B(n_144),
.Y(n_197)
);

XOR2xp5_ASAP7_75t_L g213 ( 
.A(n_197),
.B(n_200),
.Y(n_213)
);

AOI21xp5_ASAP7_75t_L g210 ( 
.A1(n_198),
.A2(n_204),
.B(n_179),
.Y(n_210)
);

CKINVDCx20_ASAP7_75t_R g199 ( 
.A(n_180),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_L g215 ( 
.A(n_199),
.B(n_205),
.Y(n_215)
);

XNOR2xp5_ASAP7_75t_L g200 ( 
.A(n_187),
.B(n_151),
.Y(n_200)
);

CKINVDCx16_ASAP7_75t_R g202 ( 
.A(n_168),
.Y(n_202)
);

XOR2xp5_ASAP7_75t_L g203 ( 
.A(n_175),
.B(n_21),
.Y(n_203)
);

OAI21xp5_ASAP7_75t_L g204 ( 
.A1(n_169),
.A2(n_19),
.B(n_7),
.Y(n_204)
);

NAND2xp5_ASAP7_75t_SL g205 ( 
.A(n_183),
.B(n_25),
.Y(n_205)
);

NAND2xp5_ASAP7_75t_L g206 ( 
.A(n_171),
.B(n_0),
.Y(n_206)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_206),
.Y(n_217)
);

XNOR2xp5_ASAP7_75t_L g209 ( 
.A(n_196),
.B(n_169),
.Y(n_209)
);

XOR2xp5_ASAP7_75t_L g235 ( 
.A(n_209),
.B(n_25),
.Y(n_235)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_210),
.Y(n_230)
);

MAJIxp5_ASAP7_75t_L g223 ( 
.A(n_211),
.B(n_212),
.C(n_214),
.Y(n_223)
);

MAJIxp5_ASAP7_75t_L g212 ( 
.A(n_195),
.B(n_188),
.C(n_168),
.Y(n_212)
);

MAJIxp5_ASAP7_75t_L g214 ( 
.A(n_195),
.B(n_181),
.C(n_185),
.Y(n_214)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_189),
.Y(n_218)
);

NAND2xp5_ASAP7_75t_L g232 ( 
.A(n_218),
.B(n_220),
.Y(n_232)
);

NOR2xp33_ASAP7_75t_L g219 ( 
.A(n_194),
.B(n_173),
.Y(n_219)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_219),
.Y(n_233)
);

MAJIxp5_ASAP7_75t_L g220 ( 
.A(n_193),
.B(n_182),
.C(n_167),
.Y(n_220)
);

NAND3xp33_ASAP7_75t_L g222 ( 
.A(n_206),
.B(n_178),
.C(n_201),
.Y(n_222)
);

NOR2xp33_ASAP7_75t_L g229 ( 
.A(n_222),
.B(n_204),
.Y(n_229)
);

NAND2xp5_ASAP7_75t_SL g224 ( 
.A(n_208),
.B(n_178),
.Y(n_224)
);

NAND2xp5_ASAP7_75t_L g240 ( 
.A(n_224),
.B(n_226),
.Y(n_240)
);

AOI21xp5_ASAP7_75t_L g225 ( 
.A1(n_207),
.A2(n_198),
.B(n_182),
.Y(n_225)
);

AOI21xp5_ASAP7_75t_L g237 ( 
.A1(n_225),
.A2(n_227),
.B(n_236),
.Y(n_237)
);

OAI22xp5_ASAP7_75t_SL g226 ( 
.A1(n_216),
.A2(n_174),
.B1(n_193),
.B2(n_200),
.Y(n_226)
);

AOI21xp5_ASAP7_75t_L g227 ( 
.A1(n_221),
.A2(n_192),
.B(n_183),
.Y(n_227)
);

AOI22xp5_ASAP7_75t_SL g228 ( 
.A1(n_215),
.A2(n_203),
.B1(n_184),
.B2(n_197),
.Y(n_228)
);

AOI22xp33_ASAP7_75t_L g242 ( 
.A1(n_228),
.A2(n_234),
.B1(n_217),
.B2(n_214),
.Y(n_242)
);

OR2x2_ASAP7_75t_L g238 ( 
.A(n_229),
.B(n_231),
.Y(n_238)
);

NOR2xp33_ASAP7_75t_L g231 ( 
.A(n_209),
.B(n_170),
.Y(n_231)
);

AOI22xp5_ASAP7_75t_SL g234 ( 
.A1(n_210),
.A2(n_186),
.B1(n_177),
.B2(n_8),
.Y(n_234)
);

MAJIxp5_ASAP7_75t_L g243 ( 
.A(n_235),
.B(n_213),
.C(n_1),
.Y(n_243)
);

OAI21xp5_ASAP7_75t_SL g236 ( 
.A1(n_212),
.A2(n_7),
.B(n_11),
.Y(n_236)
);

CKINVDCx20_ASAP7_75t_R g239 ( 
.A(n_232),
.Y(n_239)
);

NAND2xp5_ASAP7_75t_L g253 ( 
.A(n_239),
.B(n_247),
.Y(n_253)
);

AOI21xp5_ASAP7_75t_L g241 ( 
.A1(n_230),
.A2(n_211),
.B(n_220),
.Y(n_241)
);

OAI21xp5_ASAP7_75t_SL g255 ( 
.A1(n_241),
.A2(n_245),
.B(n_9),
.Y(n_255)
);

NOR2xp33_ASAP7_75t_L g250 ( 
.A(n_242),
.B(n_247),
.Y(n_250)
);

XOR2xp5_ASAP7_75t_L g249 ( 
.A(n_243),
.B(n_244),
.Y(n_249)
);

XNOR2xp5_ASAP7_75t_L g244 ( 
.A(n_223),
.B(n_213),
.Y(n_244)
);

AOI21xp5_ASAP7_75t_L g245 ( 
.A1(n_225),
.A2(n_6),
.B(n_11),
.Y(n_245)
);

XNOR2xp5_ASAP7_75t_SL g246 ( 
.A(n_226),
.B(n_8),
.Y(n_246)
);

XOR2xp5_ASAP7_75t_L g254 ( 
.A(n_246),
.B(n_10),
.Y(n_254)
);

NAND3xp33_ASAP7_75t_L g247 ( 
.A(n_233),
.B(n_8),
.C(n_11),
.Y(n_247)
);

NOR2xp33_ASAP7_75t_SL g248 ( 
.A(n_238),
.B(n_234),
.Y(n_248)
);

NAND2xp5_ASAP7_75t_SL g261 ( 
.A(n_248),
.B(n_253),
.Y(n_261)
);

OAI21xp5_ASAP7_75t_L g251 ( 
.A1(n_237),
.A2(n_223),
.B(n_235),
.Y(n_251)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_251),
.Y(n_262)
);

AOI21xp5_ASAP7_75t_SL g252 ( 
.A1(n_240),
.A2(n_228),
.B(n_10),
.Y(n_252)
);

OAI21xp5_ASAP7_75t_SL g260 ( 
.A1(n_252),
.A2(n_0),
.B(n_1),
.Y(n_260)
);

AOI21x1_ASAP7_75t_SL g259 ( 
.A1(n_254),
.A2(n_255),
.B(n_256),
.Y(n_259)
);

AOI22xp5_ASAP7_75t_L g256 ( 
.A1(n_240),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_256)
);

NOR2x1_ASAP7_75t_SL g257 ( 
.A(n_250),
.B(n_0),
.Y(n_257)
);

NAND2xp5_ASAP7_75t_SL g266 ( 
.A(n_257),
.B(n_258),
.Y(n_266)
);

INVx1_ASAP7_75t_SL g258 ( 
.A(n_252),
.Y(n_258)
);

MAJIxp5_ASAP7_75t_L g263 ( 
.A(n_260),
.B(n_250),
.C(n_261),
.Y(n_263)
);

MAJIxp5_ASAP7_75t_L g267 ( 
.A(n_263),
.B(n_264),
.C(n_265),
.Y(n_267)
);

MAJIxp5_ASAP7_75t_L g264 ( 
.A(n_262),
.B(n_249),
.C(n_2),
.Y(n_264)
);

OAI21xp5_ASAP7_75t_L g265 ( 
.A1(n_259),
.A2(n_1),
.B(n_3),
.Y(n_265)
);

MAJIxp5_ASAP7_75t_L g268 ( 
.A(n_266),
.B(n_3),
.C(n_4),
.Y(n_268)
);

OAI21xp5_ASAP7_75t_SL g269 ( 
.A1(n_268),
.A2(n_4),
.B(n_5),
.Y(n_269)
);

MAJx2_ASAP7_75t_L g270 ( 
.A(n_269),
.B(n_267),
.C(n_25),
.Y(n_270)
);

AOI211xp5_ASAP7_75t_L g271 ( 
.A1(n_270),
.A2(n_25),
.B(n_65),
.C(n_260),
.Y(n_271)
);

XNOR2xp5_ASAP7_75t_L g272 ( 
.A(n_271),
.B(n_65),
.Y(n_272)
);


endmodule