module real_aes_8759_n_104 (n_17, n_28, n_76, n_56, n_34, n_98, n_90, n_82, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_83, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_91, n_100, n_43, n_103, n_96, n_54, n_35, n_42, n_99, n_15, n_9, n_23, n_72, n_95, n_44, n_102, n_7, n_4, n_80, n_6, n_12, n_68, n_79, n_69, n_46, n_59, n_25, n_73, n_77, n_81, n_48, n_37, n_97, n_70, n_50, n_89, n_26, n_86, n_93, n_13, n_24, n_2, n_55, n_62, n_84, n_67, n_92, n_33, n_88, n_14, n_11, n_85, n_16, n_94, n_39, n_5, n_45, n_60, n_38, n_87, n_0, n_78, n_101, n_63, n_1, n_53, n_36, n_104);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_98;
input n_90;
input n_82;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_83;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_91;
input n_100;
input n_43;
input n_103;
input n_96;
input n_54;
input n_35;
input n_42;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_95;
input n_44;
input n_102;
input n_7;
input n_4;
input n_80;
input n_6;
input n_12;
input n_68;
input n_79;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_81;
input n_48;
input n_37;
input n_97;
input n_70;
input n_50;
input n_89;
input n_26;
input n_86;
input n_93;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_84;
input n_67;
input n_92;
input n_33;
input n_88;
input n_14;
input n_11;
input n_85;
input n_16;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_87;
input n_0;
input n_78;
input n_101;
input n_63;
input n_1;
input n_53;
input n_36;
output n_104;
wire n_480;
wire n_113;
wire n_476;
wire n_599;
wire n_187;
wire n_436;
wire n_684;
wire n_257;
wire n_390;
wire n_185;
wire n_285;
wire n_624;
wire n_618;
wire n_522;
wire n_485;
wire n_222;
wire n_750;
wire n_631;
wire n_287;
wire n_357;
wire n_503;
wire n_635;
wire n_386;
wire n_673;
wire n_518;
wire n_254;
wire n_207;
wire n_665;
wire n_667;
wire n_577;
wire n_580;
wire n_469;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_718;
wire n_318;
wire n_355;
wire n_239;
wire n_669;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_742;
wire n_112;
wire n_364;
wire n_421;
wire n_319;
wire n_555;
wire n_329;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_169;
wire n_242;
wire n_376;
wire n_549;
wire n_571;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_752;
wire n_448;
wire n_545;
wire n_341;
wire n_556;
wire n_593;
wire n_232;
wire n_460;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_537;
wire n_320;
wire n_551;
wire n_666;
wire n_560;
wire n_260;
wire n_660;
wire n_594;
wire n_186;
wire n_138;
wire n_696;
wire n_704;
wire n_379;
wire n_374;
wire n_453;
wire n_647;
wire n_235;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_161;
wire n_189;
wire n_271;
wire n_489;
wire n_427;
wire n_548;
wire n_678;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_519;
wire n_564;
wire n_638;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_512;
wire n_395;
wire n_332;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_116;
wire n_625;
wire n_462;
wire n_289;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_716;
wire n_213;
wire n_478;
wire n_356;
wire n_584;
wire n_408;
wire n_553;
wire n_184;
wire n_372;
wire n_528;
wire n_578;
wire n_202;
wire n_495;
wire n_370;
wire n_384;
wire n_744;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_467;
wire n_327;
wire n_106;
wire n_559;
wire n_466;
wire n_636;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_726;
wire n_517;
wire n_683;
wire n_174;
wire n_570;
wire n_675;
wire n_530;
wire n_535;
wire n_732;
wire n_211;
wire n_281;
wire n_496;
wire n_693;
wire n_173;
wire n_468;
wire n_234;
wire n_746;
wire n_284;
wire n_153;
wire n_532;
wire n_316;
wire n_656;
wire n_178;
wire n_409;
wire n_748;
wire n_298;
wire n_523;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_297;
wire n_383;
wire n_529;
wire n_119;
wire n_310;
wire n_455;
wire n_504;
wire n_725;
wire n_164;
wire n_671;
wire n_231;
wire n_547;
wire n_659;
wire n_634;
wire n_682;
wire n_454;
wire n_122;
wire n_565;
wire n_443;
wire n_608;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_267;
wire n_218;
wire n_737;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_722;
wire n_745;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_331;
wire n_449;
wire n_182;
wire n_363;
wire n_754;
wire n_417;
wire n_607;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_142;
wire n_561;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_655;
wire n_654;
wire n_527;
wire n_505;
wire n_434;
wire n_502;
wire n_600;
wire n_731;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_602;
wire n_402;
wire n_617;
wire n_552;
wire n_733;
wire n_171;
wire n_676;
wire n_658;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_146;
wire n_432;
wire n_226;
wire n_255;
wire n_286;
wire n_416;
wire n_410;
wire n_120;
wire n_751;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_695;
wire n_685;
wire n_165;
wire n_361;
wire n_632;
wire n_246;
wire n_176;
wire n_412;
wire n_163;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_501;
wire n_488;
wire n_251;
wire n_642;
wire n_613;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_702;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_734;
wire n_110;
wire n_392;
wire n_562;
wire n_150;
wire n_147;
wire n_288;
wire n_404;
wire n_713;
wire n_598;
wire n_728;
wire n_735;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_569;
wire n_563;
wire n_188;
wire n_269;
wire n_430;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_193;
wire n_397;
wire n_293;
wire n_162;
wire n_749;
wire n_385;
wire n_358;
wire n_214;
wire n_275;
wire n_649;
wire n_663;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_707;
wire n_622;
wire n_470;
wire n_133;
wire n_494;
wire n_711;
wire n_377;
wire n_273;
wire n_723;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_265;
wire n_354;
wire n_720;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_730;
wire n_643;
wire n_747;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_148;
wire n_498;
wire n_481;
wire n_691;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_233;
wire n_487;
wire n_290;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_155;
wire n_243;
wire n_692;
wire n_544;
wire n_268;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_738;
wire n_701;
wire n_309;
wire n_344;
wire n_107;
wire n_229;
wire n_482;
wire n_520;
wire n_633;
wire n_679;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_262;
wire n_630;
wire n_689;
wire n_715;
wire n_134;
wire n_420;
wire n_336;
wire n_349;
wire n_612;
wire n_195;
wire n_438;
wire n_300;
wire n_252;
wire n_283;
wire n_314;
wire n_741;
wire n_753;
wire n_249;
wire n_623;
wire n_446;
wire n_721;
wire n_221;
wire n_681;
wire n_456;
wire n_156;
wire n_359;
wire n_717;
wire n_312;
wire n_183;
wire n_266;
wire n_712;
wire n_205;
wire n_433;
wire n_516;
wire n_177;
wire n_335;
wire n_313;
wire n_627;
wire n_739;
wire n_140;
wire n_521;
wire n_418;
wire n_422;
wire n_219;
wire n_524;
wire n_705;
wire n_180;
wire n_212;
wire n_210;
wire n_575;
wire n_325;
wire n_479;
wire n_338;
wire n_442;
wire n_698;
wire n_371;
wire n_740;
wire n_166;
wire n_541;
wire n_224;
wire n_151;
wire n_546;
wire n_587;
wire n_639;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_724;
wire n_440;
wire n_525;
wire n_644;
wire n_674;
wire n_152;
wire n_198;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_414;
wire n_123;
wire n_279;
wire n_686;
wire n_543;
wire n_497;
wire n_514;
wire n_507;
wire n_270;
wire n_614;
wire n_305;
wire n_586;
wire n_450;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_465;
wire n_473;
wire n_719;
wire n_566;
wire n_474;
wire n_170;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_168;
wire n_175;
wire n_241;
wire n_687;
wire n_729;
wire n_646;
wire n_650;
wire n_710;
wire n_105;
wire n_743;
wire n_393;
wire n_294;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_500;
wire n_307;
wire n_601;
wire n_661;
wire n_463;
wire n_396;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_143;
wire n_192;
wire n_475;
wire n_554;
wire n_264;
wire n_237;
wire n_668;
NAND3xp33_ASAP7_75t_SL g112 ( .A(n_0), .B(n_113), .C(n_114), .Y(n_112) );
INVx1_ASAP7_75t_L g127 ( .A(n_0), .Y(n_127) );
AOI22xp5_ASAP7_75t_L g460 ( .A1(n_1), .A2(n_461), .B1(n_462), .B2(n_463), .Y(n_460) );
INVx1_ASAP7_75t_L g461 ( .A(n_1), .Y(n_461) );
A2O1A1Ixp33_ASAP7_75t_L g194 ( .A1(n_2), .A2(n_152), .B(n_157), .C(n_195), .Y(n_194) );
AOI21xp5_ASAP7_75t_L g243 ( .A1(n_3), .A2(n_147), .B(n_244), .Y(n_243) );
INVx1_ASAP7_75t_L g509 ( .A(n_4), .Y(n_509) );
NAND2xp5_ASAP7_75t_L g251 ( .A(n_5), .B(n_185), .Y(n_251) );
AOI21xp33_ASAP7_75t_L g516 ( .A1(n_6), .A2(n_147), .B(n_517), .Y(n_516) );
AND2x6_ASAP7_75t_L g152 ( .A(n_7), .B(n_153), .Y(n_152) );
AOI21xp5_ASAP7_75t_L g495 ( .A1(n_8), .A2(n_282), .B(n_496), .Y(n_495) );
INVx1_ASAP7_75t_L g164 ( .A(n_9), .Y(n_164) );
INVx1_ASAP7_75t_L g110 ( .A(n_10), .Y(n_110) );
NOR2xp33_ASAP7_75t_L g128 ( .A(n_10), .B(n_43), .Y(n_128) );
OAI22xp5_ASAP7_75t_L g463 ( .A1(n_11), .A2(n_33), .B1(n_464), .B2(n_465), .Y(n_463) );
CKINVDCx20_ASAP7_75t_R g465 ( .A(n_11), .Y(n_465) );
NAND2xp5_ASAP7_75t_SL g199 ( .A(n_12), .B(n_162), .Y(n_199) );
NAND2xp5_ASAP7_75t_L g488 ( .A(n_13), .B(n_209), .Y(n_488) );
INVx1_ASAP7_75t_L g521 ( .A(n_14), .Y(n_521) );
INVx1_ASAP7_75t_L g145 ( .A(n_15), .Y(n_145) );
INVx1_ASAP7_75t_L g500 ( .A(n_16), .Y(n_500) );
A2O1A1Ixp33_ASAP7_75t_L g178 ( .A1(n_17), .A2(n_165), .B(n_179), .C(n_183), .Y(n_178) );
NAND2xp5_ASAP7_75t_L g184 ( .A(n_18), .B(n_185), .Y(n_184) );
NAND2xp5_ASAP7_75t_L g564 ( .A(n_19), .B(n_479), .Y(n_564) );
NAND2xp5_ASAP7_75t_SL g474 ( .A(n_20), .B(n_147), .Y(n_474) );
NAND2xp5_ASAP7_75t_L g290 ( .A(n_21), .B(n_291), .Y(n_290) );
A2O1A1Ixp33_ASAP7_75t_L g208 ( .A1(n_22), .A2(n_209), .B(n_210), .C(n_212), .Y(n_208) );
NAND2xp5_ASAP7_75t_L g540 ( .A(n_23), .B(n_185), .Y(n_540) );
NAND2xp5_ASAP7_75t_SL g237 ( .A(n_24), .B(n_162), .Y(n_237) );
A2O1A1Ixp33_ASAP7_75t_L g498 ( .A1(n_25), .A2(n_181), .B(n_183), .C(n_499), .Y(n_498) );
NAND2xp5_ASAP7_75t_SL g223 ( .A(n_26), .B(n_162), .Y(n_223) );
CKINVDCx16_ASAP7_75t_R g233 ( .A(n_27), .Y(n_233) );
INVx1_ASAP7_75t_L g221 ( .A(n_28), .Y(n_221) );
BUFx6f_ASAP7_75t_L g151 ( .A(n_29), .Y(n_151) );
CKINVDCx20_ASAP7_75t_R g192 ( .A(n_30), .Y(n_192) );
NAND2xp5_ASAP7_75t_L g510 ( .A(n_31), .B(n_162), .Y(n_510) );
NAND2xp5_ASAP7_75t_L g451 ( .A(n_32), .B(n_452), .Y(n_451) );
INVx1_ASAP7_75t_L g464 ( .A(n_33), .Y(n_464) );
INVx1_ASAP7_75t_L g287 ( .A(n_34), .Y(n_287) );
INVx1_ASAP7_75t_L g529 ( .A(n_35), .Y(n_529) );
INVx2_ASAP7_75t_L g150 ( .A(n_36), .Y(n_150) );
CKINVDCx20_ASAP7_75t_R g202 ( .A(n_37), .Y(n_202) );
A2O1A1Ixp33_ASAP7_75t_L g246 ( .A1(n_38), .A2(n_209), .B(n_247), .C(n_249), .Y(n_246) );
INVxp67_ASAP7_75t_L g288 ( .A(n_39), .Y(n_288) );
A2O1A1Ixp33_ASAP7_75t_L g219 ( .A1(n_40), .A2(n_157), .B(n_220), .C(n_226), .Y(n_219) );
CKINVDCx14_ASAP7_75t_R g245 ( .A(n_41), .Y(n_245) );
A2O1A1Ixp33_ASAP7_75t_L g475 ( .A1(n_42), .A2(n_152), .B(n_157), .C(n_476), .Y(n_475) );
NAND2xp5_ASAP7_75t_L g109 ( .A(n_43), .B(n_110), .Y(n_109) );
INVx1_ASAP7_75t_L g528 ( .A(n_44), .Y(n_528) );
A2O1A1Ixp33_ASAP7_75t_L g160 ( .A1(n_45), .A2(n_161), .B(n_163), .C(n_166), .Y(n_160) );
NAND2xp5_ASAP7_75t_SL g563 ( .A(n_46), .B(n_162), .Y(n_563) );
CKINVDCx20_ASAP7_75t_R g228 ( .A(n_47), .Y(n_228) );
CKINVDCx20_ASAP7_75t_R g284 ( .A(n_48), .Y(n_284) );
INVx1_ASAP7_75t_L g207 ( .A(n_49), .Y(n_207) );
CKINVDCx16_ASAP7_75t_R g530 ( .A(n_50), .Y(n_530) );
NAND2xp5_ASAP7_75t_L g490 ( .A(n_51), .B(n_147), .Y(n_490) );
AOI22xp5_ASAP7_75t_L g526 ( .A1(n_52), .A2(n_157), .B1(n_212), .B2(n_527), .Y(n_526) );
AOI22xp33_ASAP7_75t_L g104 ( .A1(n_53), .A2(n_105), .B1(n_117), .B2(n_754), .Y(n_104) );
CKINVDCx20_ASAP7_75t_R g481 ( .A(n_54), .Y(n_481) );
CKINVDCx16_ASAP7_75t_R g506 ( .A(n_55), .Y(n_506) );
CKINVDCx14_ASAP7_75t_R g155 ( .A(n_56), .Y(n_155) );
A2O1A1Ixp33_ASAP7_75t_L g519 ( .A1(n_57), .A2(n_161), .B(n_249), .C(n_520), .Y(n_519) );
CKINVDCx20_ASAP7_75t_R g566 ( .A(n_58), .Y(n_566) );
INVx1_ASAP7_75t_L g518 ( .A(n_59), .Y(n_518) );
INVx1_ASAP7_75t_L g153 ( .A(n_60), .Y(n_153) );
INVx1_ASAP7_75t_L g144 ( .A(n_61), .Y(n_144) );
INVx1_ASAP7_75t_SL g248 ( .A(n_62), .Y(n_248) );
CKINVDCx20_ASAP7_75t_R g121 ( .A(n_63), .Y(n_121) );
NAND2xp5_ASAP7_75t_L g214 ( .A(n_64), .B(n_185), .Y(n_214) );
INVx1_ASAP7_75t_L g236 ( .A(n_65), .Y(n_236) );
A2O1A1Ixp33_ASAP7_75t_SL g537 ( .A1(n_66), .A2(n_249), .B(n_479), .C(n_538), .Y(n_537) );
INVxp67_ASAP7_75t_L g539 ( .A(n_67), .Y(n_539) );
INVx1_ASAP7_75t_L g116 ( .A(n_68), .Y(n_116) );
AOI21xp5_ASAP7_75t_L g146 ( .A1(n_69), .A2(n_147), .B(n_154), .Y(n_146) );
CKINVDCx20_ASAP7_75t_R g240 ( .A(n_70), .Y(n_240) );
AOI21xp5_ASAP7_75t_L g175 ( .A1(n_71), .A2(n_147), .B(n_176), .Y(n_175) );
CKINVDCx20_ASAP7_75t_R g532 ( .A(n_72), .Y(n_532) );
INVx1_ASAP7_75t_L g560 ( .A(n_73), .Y(n_560) );
AOI21xp5_ASAP7_75t_L g281 ( .A1(n_74), .A2(n_282), .B(n_283), .Y(n_281) );
INVx1_ASAP7_75t_L g177 ( .A(n_75), .Y(n_177) );
CKINVDCx16_ASAP7_75t_R g218 ( .A(n_76), .Y(n_218) );
OAI22xp5_ASAP7_75t_SL g447 ( .A1(n_77), .A2(n_78), .B1(n_448), .B2(n_449), .Y(n_447) );
CKINVDCx20_ASAP7_75t_R g449 ( .A(n_77), .Y(n_449) );
CKINVDCx20_ASAP7_75t_R g448 ( .A(n_78), .Y(n_448) );
A2O1A1Ixp33_ASAP7_75t_L g561 ( .A1(n_79), .A2(n_152), .B(n_157), .C(n_562), .Y(n_561) );
AOI22xp5_ASAP7_75t_SL g455 ( .A1(n_80), .A2(n_125), .B1(n_456), .B2(n_749), .Y(n_455) );
AOI21xp5_ASAP7_75t_L g205 ( .A1(n_81), .A2(n_147), .B(n_206), .Y(n_205) );
INVx1_ASAP7_75t_L g180 ( .A(n_82), .Y(n_180) );
NAND2xp5_ASAP7_75t_SL g477 ( .A(n_83), .B(n_222), .Y(n_477) );
INVx2_ASAP7_75t_L g142 ( .A(n_84), .Y(n_142) );
INVx1_ASAP7_75t_L g196 ( .A(n_85), .Y(n_196) );
NAND2xp5_ASAP7_75t_L g478 ( .A(n_86), .B(n_479), .Y(n_478) );
A2O1A1Ixp33_ASAP7_75t_L g507 ( .A1(n_87), .A2(n_152), .B(n_157), .C(n_508), .Y(n_507) );
INVx2_ASAP7_75t_L g113 ( .A(n_88), .Y(n_113) );
OR2x2_ASAP7_75t_L g124 ( .A(n_88), .B(n_125), .Y(n_124) );
A2O1A1Ixp33_ASAP7_75t_L g234 ( .A1(n_89), .A2(n_157), .B(n_235), .C(n_238), .Y(n_234) );
OAI22xp5_ASAP7_75t_SL g130 ( .A1(n_90), .A2(n_92), .B1(n_131), .B2(n_132), .Y(n_130) );
CKINVDCx20_ASAP7_75t_R g132 ( .A(n_90), .Y(n_132) );
NAND2xp5_ASAP7_75t_L g522 ( .A(n_91), .B(n_141), .Y(n_522) );
CKINVDCx20_ASAP7_75t_R g131 ( .A(n_92), .Y(n_131) );
A2O1A1Ixp33_ASAP7_75t_L g485 ( .A1(n_93), .A2(n_152), .B(n_157), .C(n_486), .Y(n_485) );
CKINVDCx20_ASAP7_75t_R g492 ( .A(n_94), .Y(n_492) );
INVx1_ASAP7_75t_L g536 ( .A(n_95), .Y(n_536) );
CKINVDCx16_ASAP7_75t_R g497 ( .A(n_96), .Y(n_497) );
NAND2xp5_ASAP7_75t_SL g487 ( .A(n_97), .B(n_222), .Y(n_487) );
NAND2xp5_ASAP7_75t_L g169 ( .A(n_98), .B(n_170), .Y(n_169) );
NAND2xp5_ASAP7_75t_L g501 ( .A(n_99), .B(n_170), .Y(n_501) );
NAND2xp5_ASAP7_75t_L g115 ( .A(n_100), .B(n_116), .Y(n_115) );
INVx2_ASAP7_75t_L g211 ( .A(n_101), .Y(n_211) );
OAI22xp5_ASAP7_75t_L g457 ( .A1(n_102), .A2(n_458), .B1(n_459), .B2(n_460), .Y(n_457) );
CKINVDCx20_ASAP7_75t_R g458 ( .A(n_102), .Y(n_458) );
AOI21xp5_ASAP7_75t_L g534 ( .A1(n_103), .A2(n_147), .B(n_535), .Y(n_534) );
INVx1_ASAP7_75t_L g105 ( .A(n_106), .Y(n_105) );
INVx2_ASAP7_75t_L g106 ( .A(n_107), .Y(n_106) );
INVx2_ASAP7_75t_L g754 ( .A(n_107), .Y(n_754) );
AND2x2_ASAP7_75t_L g107 ( .A(n_108), .B(n_111), .Y(n_107) );
INVx1_ASAP7_75t_L g108 ( .A(n_109), .Y(n_108) );
INVx1_ASAP7_75t_L g111 ( .A(n_112), .Y(n_111) );
INVx1_ASAP7_75t_L g747 ( .A(n_113), .Y(n_747) );
NOR2x2_ASAP7_75t_L g751 ( .A(n_113), .B(n_125), .Y(n_751) );
INVx1_ASAP7_75t_SL g114 ( .A(n_115), .Y(n_114) );
OA21x2_ASAP7_75t_L g117 ( .A1(n_118), .A2(n_122), .B(n_454), .Y(n_117) );
BUFx2_ASAP7_75t_L g118 ( .A(n_119), .Y(n_118) );
BUFx2_ASAP7_75t_L g119 ( .A(n_120), .Y(n_119) );
INVx1_ASAP7_75t_L g753 ( .A(n_120), .Y(n_753) );
INVx2_ASAP7_75t_L g120 ( .A(n_121), .Y(n_120) );
OAI21xp5_ASAP7_75t_L g122 ( .A1(n_123), .A2(n_129), .B(n_451), .Y(n_122) );
INVx1_ASAP7_75t_SL g123 ( .A(n_124), .Y(n_123) );
HB1xp67_ASAP7_75t_L g453 ( .A(n_124), .Y(n_453) );
INVx2_ASAP7_75t_L g125 ( .A(n_126), .Y(n_125) );
AND2x2_ASAP7_75t_L g126 ( .A(n_127), .B(n_128), .Y(n_126) );
AOI22xp33_ASAP7_75t_L g129 ( .A1(n_130), .A2(n_133), .B1(n_134), .B2(n_450), .Y(n_129) );
CKINVDCx20_ASAP7_75t_R g450 ( .A(n_130), .Y(n_450) );
NOR2xp33_ASAP7_75t_L g512 ( .A(n_131), .B(n_190), .Y(n_512) );
INVx1_ASAP7_75t_L g133 ( .A(n_134), .Y(n_133) );
XOR2xp5_ASAP7_75t_L g134 ( .A(n_135), .B(n_447), .Y(n_134) );
INVx2_ASAP7_75t_L g748 ( .A(n_135), .Y(n_748) );
OR2x2_ASAP7_75t_L g135 ( .A(n_136), .B(n_377), .Y(n_135) );
NAND5xp2_ASAP7_75t_L g136 ( .A(n_137), .B(n_292), .C(n_324), .D(n_341), .E(n_364), .Y(n_136) );
AOI221xp5_ASAP7_75t_L g137 ( .A1(n_138), .A2(n_215), .B1(n_252), .B2(n_256), .C(n_260), .Y(n_137) );
INVx1_ASAP7_75t_L g404 ( .A(n_138), .Y(n_404) );
AND2x2_ASAP7_75t_L g138 ( .A(n_139), .B(n_187), .Y(n_138) );
AND3x2_ASAP7_75t_L g379 ( .A(n_139), .B(n_189), .C(n_380), .Y(n_379) );
AND2x2_ASAP7_75t_L g139 ( .A(n_140), .B(n_172), .Y(n_139) );
NAND2xp5_ASAP7_75t_L g257 ( .A(n_140), .B(n_258), .Y(n_257) );
BUFx3_ASAP7_75t_L g267 ( .A(n_140), .Y(n_267) );
AND2x2_ASAP7_75t_L g271 ( .A(n_140), .B(n_203), .Y(n_271) );
INVx2_ASAP7_75t_L g301 ( .A(n_140), .Y(n_301) );
OR2x2_ASAP7_75t_L g312 ( .A(n_140), .B(n_204), .Y(n_312) );
NOR2xp33_ASAP7_75t_L g331 ( .A(n_140), .B(n_188), .Y(n_331) );
NAND2xp5_ASAP7_75t_L g349 ( .A(n_140), .B(n_350), .Y(n_349) );
AND2x2_ASAP7_75t_L g391 ( .A(n_140), .B(n_204), .Y(n_391) );
OA21x2_ASAP7_75t_L g140 ( .A1(n_141), .A2(n_146), .B(n_169), .Y(n_140) );
INVx1_ASAP7_75t_L g190 ( .A(n_141), .Y(n_190) );
O2A1O1Ixp33_ASAP7_75t_L g217 ( .A1(n_141), .A2(n_193), .B(n_218), .C(n_219), .Y(n_217) );
INVx2_ASAP7_75t_L g241 ( .A(n_141), .Y(n_241) );
OA21x2_ASAP7_75t_L g494 ( .A1(n_141), .A2(n_495), .B(n_501), .Y(n_494) );
AND2x2_ASAP7_75t_SL g141 ( .A(n_142), .B(n_143), .Y(n_141) );
AND2x2_ASAP7_75t_L g171 ( .A(n_142), .B(n_143), .Y(n_171) );
NAND2xp5_ASAP7_75t_L g143 ( .A(n_144), .B(n_145), .Y(n_143) );
BUFx2_ASAP7_75t_L g282 ( .A(n_147), .Y(n_282) );
AND2x4_ASAP7_75t_L g147 ( .A(n_148), .B(n_152), .Y(n_147) );
NAND2x1p5_ASAP7_75t_L g193 ( .A(n_148), .B(n_152), .Y(n_193) );
AND2x2_ASAP7_75t_L g148 ( .A(n_149), .B(n_151), .Y(n_148) );
INVx1_ASAP7_75t_L g225 ( .A(n_149), .Y(n_225) );
INVx1_ASAP7_75t_L g149 ( .A(n_150), .Y(n_149) );
INVx2_ASAP7_75t_L g158 ( .A(n_150), .Y(n_158) );
INVx1_ASAP7_75t_L g213 ( .A(n_150), .Y(n_213) );
INVx1_ASAP7_75t_L g159 ( .A(n_151), .Y(n_159) );
BUFx6f_ASAP7_75t_L g162 ( .A(n_151), .Y(n_162) );
INVx3_ASAP7_75t_L g165 ( .A(n_151), .Y(n_165) );
BUFx6f_ASAP7_75t_L g182 ( .A(n_151), .Y(n_182) );
INVx1_ASAP7_75t_L g479 ( .A(n_151), .Y(n_479) );
INVx4_ASAP7_75t_SL g168 ( .A(n_152), .Y(n_168) );
BUFx3_ASAP7_75t_L g226 ( .A(n_152), .Y(n_226) );
O2A1O1Ixp33_ASAP7_75t_SL g154 ( .A1(n_155), .A2(n_156), .B(n_160), .C(n_168), .Y(n_154) );
O2A1O1Ixp33_ASAP7_75t_SL g176 ( .A1(n_156), .A2(n_168), .B(n_177), .C(n_178), .Y(n_176) );
O2A1O1Ixp33_ASAP7_75t_SL g206 ( .A1(n_156), .A2(n_168), .B(n_207), .C(n_208), .Y(n_206) );
O2A1O1Ixp33_ASAP7_75t_L g244 ( .A1(n_156), .A2(n_168), .B(n_245), .C(n_246), .Y(n_244) );
O2A1O1Ixp33_ASAP7_75t_SL g283 ( .A1(n_156), .A2(n_168), .B(n_284), .C(n_285), .Y(n_283) );
O2A1O1Ixp33_ASAP7_75t_L g496 ( .A1(n_156), .A2(n_168), .B(n_497), .C(n_498), .Y(n_496) );
O2A1O1Ixp33_ASAP7_75t_L g517 ( .A1(n_156), .A2(n_168), .B(n_518), .C(n_519), .Y(n_517) );
O2A1O1Ixp33_ASAP7_75t_L g535 ( .A1(n_156), .A2(n_168), .B(n_536), .C(n_537), .Y(n_535) );
INVx5_ASAP7_75t_L g156 ( .A(n_157), .Y(n_156) );
AND2x6_ASAP7_75t_L g157 ( .A(n_158), .B(n_159), .Y(n_157) );
BUFx3_ASAP7_75t_L g167 ( .A(n_158), .Y(n_167) );
BUFx6f_ASAP7_75t_L g250 ( .A(n_158), .Y(n_250) );
INVx2_ASAP7_75t_L g161 ( .A(n_162), .Y(n_161) );
INVx4_ASAP7_75t_L g209 ( .A(n_162), .Y(n_209) );
NOR2xp33_ASAP7_75t_L g163 ( .A(n_164), .B(n_165), .Y(n_163) );
INVx5_ASAP7_75t_L g222 ( .A(n_165), .Y(n_222) );
NOR2xp33_ASAP7_75t_L g520 ( .A(n_165), .B(n_521), .Y(n_520) );
NOR2xp33_ASAP7_75t_L g538 ( .A(n_165), .B(n_539), .Y(n_538) );
INVx2_ASAP7_75t_L g200 ( .A(n_166), .Y(n_200) );
INVx2_ASAP7_75t_L g166 ( .A(n_167), .Y(n_166) );
INVx1_ASAP7_75t_L g183 ( .A(n_167), .Y(n_183) );
INVx1_ASAP7_75t_L g238 ( .A(n_168), .Y(n_238) );
OAI22xp33_ASAP7_75t_L g525 ( .A1(n_168), .A2(n_193), .B1(n_526), .B2(n_530), .Y(n_525) );
HB1xp67_ASAP7_75t_L g174 ( .A(n_170), .Y(n_174) );
INVx4_ASAP7_75t_L g186 ( .A(n_170), .Y(n_186) );
OA21x2_ASAP7_75t_L g533 ( .A1(n_170), .A2(n_534), .B(n_540), .Y(n_533) );
BUFx6f_ASAP7_75t_L g170 ( .A(n_171), .Y(n_170) );
INVx1_ASAP7_75t_L g279 ( .A(n_171), .Y(n_279) );
HB1xp67_ASAP7_75t_L g270 ( .A(n_172), .Y(n_270) );
AND2x2_ASAP7_75t_L g332 ( .A(n_172), .B(n_333), .Y(n_332) );
NAND2xp5_ASAP7_75t_L g351 ( .A(n_172), .B(n_188), .Y(n_351) );
INVx1_ASAP7_75t_SL g172 ( .A(n_173), .Y(n_172) );
OR2x2_ASAP7_75t_L g259 ( .A(n_173), .B(n_188), .Y(n_259) );
HB1xp67_ASAP7_75t_L g266 ( .A(n_173), .Y(n_266) );
AND2x2_ASAP7_75t_L g318 ( .A(n_173), .B(n_204), .Y(n_318) );
NAND3xp33_ASAP7_75t_L g343 ( .A(n_173), .B(n_187), .C(n_301), .Y(n_343) );
AND2x2_ASAP7_75t_L g408 ( .A(n_173), .B(n_189), .Y(n_408) );
AND2x2_ASAP7_75t_L g442 ( .A(n_173), .B(n_188), .Y(n_442) );
OA21x2_ASAP7_75t_L g173 ( .A1(n_174), .A2(n_175), .B(n_184), .Y(n_173) );
OA21x2_ASAP7_75t_L g204 ( .A1(n_174), .A2(n_205), .B(n_214), .Y(n_204) );
OA21x2_ASAP7_75t_L g242 ( .A1(n_174), .A2(n_243), .B(n_251), .Y(n_242) );
NOR2xp33_ASAP7_75t_L g179 ( .A(n_180), .B(n_181), .Y(n_179) );
NOR2xp33_ASAP7_75t_L g210 ( .A(n_181), .B(n_211), .Y(n_210) );
OAI22xp33_ASAP7_75t_L g286 ( .A1(n_181), .A2(n_222), .B1(n_287), .B2(n_288), .Y(n_286) );
NOR2xp33_ASAP7_75t_L g499 ( .A(n_181), .B(n_500), .Y(n_499) );
INVx4_ASAP7_75t_L g181 ( .A(n_182), .Y(n_181) );
INVx2_ASAP7_75t_L g198 ( .A(n_182), .Y(n_198) );
OAI22xp5_ASAP7_75t_SL g527 ( .A1(n_182), .A2(n_198), .B1(n_528), .B2(n_529), .Y(n_527) );
OA21x2_ASAP7_75t_L g515 ( .A1(n_185), .A2(n_516), .B(n_522), .Y(n_515) );
INVx3_ASAP7_75t_L g185 ( .A(n_186), .Y(n_185) );
NOR2xp33_ASAP7_75t_L g201 ( .A(n_186), .B(n_202), .Y(n_201) );
NOR2xp33_ASAP7_75t_L g227 ( .A(n_186), .B(n_228), .Y(n_227) );
AO21x2_ASAP7_75t_L g231 ( .A1(n_186), .A2(n_232), .B(n_239), .Y(n_231) );
NOR2xp33_ASAP7_75t_SL g480 ( .A(n_186), .B(n_481), .Y(n_480) );
INVxp67_ASAP7_75t_L g268 ( .A(n_187), .Y(n_268) );
AND2x2_ASAP7_75t_L g187 ( .A(n_188), .B(n_203), .Y(n_187) );
NAND2xp5_ASAP7_75t_L g319 ( .A(n_188), .B(n_301), .Y(n_319) );
NAND2xp5_ASAP7_75t_L g340 ( .A(n_188), .B(n_332), .Y(n_340) );
AND2x2_ASAP7_75t_L g390 ( .A(n_188), .B(n_391), .Y(n_390) );
INVx1_ASAP7_75t_L g418 ( .A(n_188), .Y(n_418) );
INVx4_ASAP7_75t_L g188 ( .A(n_189), .Y(n_188) );
AND2x2_ASAP7_75t_L g325 ( .A(n_189), .B(n_318), .Y(n_325) );
BUFx3_ASAP7_75t_L g357 ( .A(n_189), .Y(n_357) );
AO21x2_ASAP7_75t_L g189 ( .A1(n_190), .A2(n_191), .B(n_201), .Y(n_189) );
NOR2xp33_ASAP7_75t_L g491 ( .A(n_190), .B(n_492), .Y(n_491) );
NOR2xp33_ASAP7_75t_L g565 ( .A(n_190), .B(n_566), .Y(n_565) );
OAI21xp5_ASAP7_75t_L g191 ( .A1(n_192), .A2(n_193), .B(n_194), .Y(n_191) );
OAI21xp5_ASAP7_75t_L g232 ( .A1(n_193), .A2(n_233), .B(n_234), .Y(n_232) );
OAI21xp5_ASAP7_75t_L g505 ( .A1(n_193), .A2(n_506), .B(n_507), .Y(n_505) );
OAI21xp5_ASAP7_75t_L g559 ( .A1(n_193), .A2(n_560), .B(n_561), .Y(n_559) );
O2A1O1Ixp5_ASAP7_75t_L g195 ( .A1(n_196), .A2(n_197), .B(n_199), .C(n_200), .Y(n_195) );
O2A1O1Ixp33_ASAP7_75t_L g235 ( .A1(n_197), .A2(n_200), .B(n_236), .C(n_237), .Y(n_235) );
INVx2_ASAP7_75t_L g197 ( .A(n_198), .Y(n_197) );
AOI21xp5_ASAP7_75t_L g476 ( .A1(n_200), .A2(n_477), .B(n_478), .Y(n_476) );
AOI21xp5_ASAP7_75t_L g562 ( .A1(n_200), .A2(n_563), .B(n_564), .Y(n_562) );
INVx2_ASAP7_75t_L g333 ( .A(n_203), .Y(n_333) );
INVx2_ASAP7_75t_L g203 ( .A(n_204), .Y(n_203) );
HB1xp67_ASAP7_75t_L g302 ( .A(n_204), .Y(n_302) );
NOR2xp33_ASAP7_75t_L g247 ( .A(n_209), .B(n_248), .Y(n_247) );
INVx2_ASAP7_75t_L g511 ( .A(n_212), .Y(n_511) );
INVx3_ASAP7_75t_L g212 ( .A(n_213), .Y(n_212) );
AOI22xp33_ASAP7_75t_L g392 ( .A1(n_215), .A2(n_393), .B1(n_395), .B2(n_396), .Y(n_392) );
AND2x2_ASAP7_75t_L g215 ( .A(n_216), .B(n_229), .Y(n_215) );
AND2x2_ASAP7_75t_L g252 ( .A(n_216), .B(n_253), .Y(n_252) );
INVx3_ASAP7_75t_SL g263 ( .A(n_216), .Y(n_263) );
NAND2xp5_ASAP7_75t_L g328 ( .A(n_216), .B(n_296), .Y(n_328) );
OR2x2_ASAP7_75t_L g347 ( .A(n_216), .B(n_230), .Y(n_347) );
AND2x2_ASAP7_75t_L g352 ( .A(n_216), .B(n_304), .Y(n_352) );
AND2x2_ASAP7_75t_L g355 ( .A(n_216), .B(n_297), .Y(n_355) );
AND2x2_ASAP7_75t_L g367 ( .A(n_216), .B(n_242), .Y(n_367) );
AND2x2_ASAP7_75t_L g383 ( .A(n_216), .B(n_231), .Y(n_383) );
AND2x4_ASAP7_75t_L g386 ( .A(n_216), .B(n_254), .Y(n_386) );
OR2x2_ASAP7_75t_L g403 ( .A(n_216), .B(n_339), .Y(n_403) );
OR2x2_ASAP7_75t_L g434 ( .A(n_216), .B(n_276), .Y(n_434) );
NAND2xp5_ASAP7_75t_SL g436 ( .A(n_216), .B(n_362), .Y(n_436) );
OR2x6_ASAP7_75t_L g216 ( .A(n_217), .B(n_227), .Y(n_216) );
O2A1O1Ixp33_ASAP7_75t_L g220 ( .A1(n_221), .A2(n_222), .B(n_223), .C(n_224), .Y(n_220) );
O2A1O1Ixp33_ASAP7_75t_L g508 ( .A1(n_222), .A2(n_509), .B(n_510), .C(n_511), .Y(n_508) );
INVx2_ASAP7_75t_L g224 ( .A(n_225), .Y(n_224) );
NAND2xp5_ASAP7_75t_SL g285 ( .A(n_225), .B(n_286), .Y(n_285) );
AND2x2_ASAP7_75t_L g310 ( .A(n_229), .B(n_274), .Y(n_310) );
NAND2xp5_ASAP7_75t_L g429 ( .A(n_229), .B(n_297), .Y(n_429) );
AND2x2_ASAP7_75t_L g229 ( .A(n_230), .B(n_242), .Y(n_229) );
AND2x2_ASAP7_75t_L g262 ( .A(n_230), .B(n_263), .Y(n_262) );
AND2x2_ASAP7_75t_L g296 ( .A(n_230), .B(n_297), .Y(n_296) );
AND2x2_ASAP7_75t_L g304 ( .A(n_230), .B(n_276), .Y(n_304) );
AND2x2_ASAP7_75t_L g322 ( .A(n_230), .B(n_254), .Y(n_322) );
OR2x2_ASAP7_75t_L g339 ( .A(n_230), .B(n_297), .Y(n_339) );
INVx2_ASAP7_75t_SL g230 ( .A(n_231), .Y(n_230) );
BUFx2_ASAP7_75t_L g255 ( .A(n_231), .Y(n_255) );
AND2x2_ASAP7_75t_L g362 ( .A(n_231), .B(n_242), .Y(n_362) );
NOR2xp33_ASAP7_75t_L g239 ( .A(n_240), .B(n_241), .Y(n_239) );
INVx1_ASAP7_75t_L g291 ( .A(n_241), .Y(n_291) );
AO21x2_ASAP7_75t_L g483 ( .A1(n_241), .A2(n_484), .B(n_491), .Y(n_483) );
INVx2_ASAP7_75t_L g254 ( .A(n_242), .Y(n_254) );
INVx1_ASAP7_75t_L g374 ( .A(n_242), .Y(n_374) );
AND2x2_ASAP7_75t_L g424 ( .A(n_242), .B(n_263), .Y(n_424) );
INVx3_ASAP7_75t_L g249 ( .A(n_250), .Y(n_249) );
HB1xp67_ASAP7_75t_L g489 ( .A(n_250), .Y(n_489) );
AND2x2_ASAP7_75t_L g273 ( .A(n_253), .B(n_274), .Y(n_273) );
AND2x2_ASAP7_75t_L g308 ( .A(n_253), .B(n_263), .Y(n_308) );
NAND2xp5_ASAP7_75t_L g354 ( .A(n_253), .B(n_355), .Y(n_354) );
AND2x2_ASAP7_75t_L g253 ( .A(n_254), .B(n_255), .Y(n_253) );
AND2x2_ASAP7_75t_L g295 ( .A(n_254), .B(n_263), .Y(n_295) );
OR2x2_ASAP7_75t_L g411 ( .A(n_255), .B(n_385), .Y(n_411) );
INVx1_ASAP7_75t_L g256 ( .A(n_257), .Y(n_256) );
NAND2xp5_ASAP7_75t_L g397 ( .A(n_258), .B(n_391), .Y(n_397) );
INVx2_ASAP7_75t_SL g258 ( .A(n_259), .Y(n_258) );
OAI32xp33_ASAP7_75t_L g353 ( .A1(n_259), .A2(n_354), .A3(n_356), .B1(n_358), .B2(n_359), .Y(n_353) );
OR2x2_ASAP7_75t_L g370 ( .A(n_259), .B(n_312), .Y(n_370) );
OAI21xp33_ASAP7_75t_SL g395 ( .A1(n_259), .A2(n_269), .B(n_300), .Y(n_395) );
OAI22xp33_ASAP7_75t_L g260 ( .A1(n_261), .A2(n_264), .B1(n_269), .B2(n_272), .Y(n_260) );
INVxp33_ASAP7_75t_L g261 ( .A(n_262), .Y(n_261) );
NAND2xp5_ASAP7_75t_L g335 ( .A(n_262), .B(n_336), .Y(n_335) );
NAND2xp5_ASAP7_75t_L g303 ( .A(n_263), .B(n_304), .Y(n_303) );
AND2x2_ASAP7_75t_L g321 ( .A(n_263), .B(n_322), .Y(n_321) );
AND2x2_ASAP7_75t_L g421 ( .A(n_263), .B(n_362), .Y(n_421) );
OR2x2_ASAP7_75t_L g445 ( .A(n_263), .B(n_339), .Y(n_445) );
AOI21xp33_ASAP7_75t_L g428 ( .A1(n_264), .A2(n_327), .B(n_429), .Y(n_428) );
OR2x2_ASAP7_75t_L g264 ( .A(n_265), .B(n_268), .Y(n_264) );
NAND2xp5_ASAP7_75t_L g265 ( .A(n_266), .B(n_267), .Y(n_265) );
INVx1_ASAP7_75t_L g305 ( .A(n_266), .Y(n_305) );
NAND2xp5_ASAP7_75t_L g323 ( .A(n_266), .B(n_271), .Y(n_323) );
AND2x2_ASAP7_75t_L g345 ( .A(n_267), .B(n_318), .Y(n_345) );
INVx1_ASAP7_75t_L g358 ( .A(n_267), .Y(n_358) );
OR2x2_ASAP7_75t_L g363 ( .A(n_267), .B(n_297), .Y(n_363) );
NAND2xp5_ASAP7_75t_L g269 ( .A(n_270), .B(n_271), .Y(n_269) );
NOR2xp33_ASAP7_75t_L g311 ( .A(n_270), .B(n_312), .Y(n_311) );
OAI22xp33_ASAP7_75t_L g293 ( .A1(n_271), .A2(n_294), .B1(n_299), .B2(n_303), .Y(n_293) );
INVx1_ASAP7_75t_L g272 ( .A(n_273), .Y(n_272) );
OAI22xp5_ASAP7_75t_L g342 ( .A1(n_274), .A2(n_336), .B1(n_343), .B2(n_344), .Y(n_342) );
AND2x2_ASAP7_75t_L g420 ( .A(n_274), .B(n_421), .Y(n_420) );
INVx2_ASAP7_75t_L g274 ( .A(n_275), .Y(n_274) );
INVx1_ASAP7_75t_SL g275 ( .A(n_276), .Y(n_275) );
NAND2xp5_ASAP7_75t_L g373 ( .A(n_276), .B(n_374), .Y(n_373) );
AND2x2_ASAP7_75t_L g439 ( .A(n_276), .B(n_322), .Y(n_439) );
AO21x2_ASAP7_75t_L g276 ( .A1(n_277), .A2(n_280), .B(n_289), .Y(n_276) );
INVx1_ASAP7_75t_L g298 ( .A(n_277), .Y(n_298) );
AO21x2_ASAP7_75t_L g558 ( .A1(n_277), .A2(n_559), .B(n_565), .Y(n_558) );
INVx1_ASAP7_75t_L g277 ( .A(n_278), .Y(n_277) );
AOI21xp5_ASAP7_75t_SL g473 ( .A1(n_278), .A2(n_474), .B(n_475), .Y(n_473) );
INVx2_ASAP7_75t_L g278 ( .A(n_279), .Y(n_278) );
AO21x2_ASAP7_75t_L g504 ( .A1(n_279), .A2(n_505), .B(n_512), .Y(n_504) );
AO21x2_ASAP7_75t_L g524 ( .A1(n_279), .A2(n_525), .B(n_531), .Y(n_524) );
NOR2xp33_ASAP7_75t_L g531 ( .A(n_279), .B(n_532), .Y(n_531) );
INVx1_ASAP7_75t_L g280 ( .A(n_281), .Y(n_280) );
OA21x2_ASAP7_75t_L g297 ( .A1(n_281), .A2(n_290), .B(n_298), .Y(n_297) );
INVx1_ASAP7_75t_L g289 ( .A(n_290), .Y(n_289) );
AOI221xp5_ASAP7_75t_L g292 ( .A1(n_293), .A2(n_305), .B1(n_306), .B2(n_311), .C(n_313), .Y(n_292) );
NAND2xp5_ASAP7_75t_L g294 ( .A(n_295), .B(n_296), .Y(n_294) );
NAND2xp5_ASAP7_75t_L g327 ( .A(n_295), .B(n_297), .Y(n_327) );
NAND2xp5_ASAP7_75t_L g337 ( .A(n_295), .B(n_338), .Y(n_337) );
INVx1_ASAP7_75t_L g314 ( .A(n_296), .Y(n_314) );
O2A1O1Ixp33_ASAP7_75t_L g401 ( .A1(n_296), .A2(n_402), .B(n_403), .C(n_404), .Y(n_401) );
AND2x2_ASAP7_75t_L g406 ( .A(n_296), .B(n_386), .Y(n_406) );
O2A1O1Ixp33_ASAP7_75t_SL g444 ( .A1(n_296), .A2(n_385), .B(n_445), .C(n_446), .Y(n_444) );
BUFx3_ASAP7_75t_L g336 ( .A(n_297), .Y(n_336) );
INVx1_ASAP7_75t_L g299 ( .A(n_300), .Y(n_299) );
NAND2xp5_ASAP7_75t_L g400 ( .A(n_300), .B(n_357), .Y(n_400) );
AOI211xp5_ASAP7_75t_L g419 ( .A1(n_300), .A2(n_420), .B(n_422), .C(n_428), .Y(n_419) );
AND2x2_ASAP7_75t_L g300 ( .A(n_301), .B(n_302), .Y(n_300) );
INVxp67_ASAP7_75t_L g380 ( .A(n_302), .Y(n_380) );
NAND2xp5_ASAP7_75t_L g423 ( .A(n_304), .B(n_424), .Y(n_423) );
NAND2xp5_ASAP7_75t_SL g306 ( .A(n_307), .B(n_309), .Y(n_306) );
INVx1_ASAP7_75t_SL g307 ( .A(n_308), .Y(n_307) );
AOI211xp5_ASAP7_75t_L g324 ( .A1(n_308), .A2(n_325), .B(n_326), .C(n_334), .Y(n_324) );
INVx1_ASAP7_75t_L g309 ( .A(n_310), .Y(n_309) );
INVx1_ASAP7_75t_L g409 ( .A(n_312), .Y(n_409) );
OR2x2_ASAP7_75t_L g426 ( .A(n_312), .B(n_356), .Y(n_426) );
OAI22xp5_ASAP7_75t_L g313 ( .A1(n_314), .A2(n_315), .B1(n_320), .B2(n_323), .Y(n_313) );
OAI22xp33_ASAP7_75t_L g326 ( .A1(n_315), .A2(n_327), .B1(n_328), .B2(n_329), .Y(n_326) );
INVx1_ASAP7_75t_L g315 ( .A(n_316), .Y(n_315) );
NOR2xp33_ASAP7_75t_L g316 ( .A(n_317), .B(n_319), .Y(n_316) );
OR2x2_ASAP7_75t_L g413 ( .A(n_317), .B(n_357), .Y(n_413) );
INVx1_ASAP7_75t_SL g317 ( .A(n_318), .Y(n_317) );
AND2x2_ASAP7_75t_L g368 ( .A(n_318), .B(n_358), .Y(n_368) );
INVx1_ASAP7_75t_L g376 ( .A(n_319), .Y(n_376) );
INVx1_ASAP7_75t_L g320 ( .A(n_321), .Y(n_320) );
NAND2xp5_ASAP7_75t_L g384 ( .A(n_322), .B(n_336), .Y(n_384) );
INVx1_ASAP7_75t_L g329 ( .A(n_330), .Y(n_329) );
AND2x2_ASAP7_75t_L g330 ( .A(n_331), .B(n_332), .Y(n_330) );
NAND2xp5_ASAP7_75t_SL g375 ( .A(n_332), .B(n_376), .Y(n_375) );
INVx2_ASAP7_75t_L g441 ( .A(n_333), .Y(n_441) );
AOI21xp33_ASAP7_75t_L g334 ( .A1(n_335), .A2(n_337), .B(n_340), .Y(n_334) );
INVx1_ASAP7_75t_L g371 ( .A(n_335), .Y(n_371) );
NAND2xp5_ASAP7_75t_SL g346 ( .A(n_336), .B(n_347), .Y(n_346) );
NAND2xp5_ASAP7_75t_L g366 ( .A(n_336), .B(n_367), .Y(n_366) );
NAND2x1p5_ASAP7_75t_L g387 ( .A(n_336), .B(n_362), .Y(n_387) );
NAND2xp5_ASAP7_75t_SL g394 ( .A(n_336), .B(n_383), .Y(n_394) );
OAI211xp5_ASAP7_75t_L g398 ( .A1(n_336), .A2(n_346), .B(n_386), .C(n_399), .Y(n_398) );
INVx1_ASAP7_75t_SL g338 ( .A(n_339), .Y(n_338) );
AOI221xp5_ASAP7_75t_SL g341 ( .A1(n_342), .A2(n_346), .B1(n_348), .B2(n_352), .C(n_353), .Y(n_341) );
INVx1_ASAP7_75t_L g344 ( .A(n_345), .Y(n_344) );
INVxp67_ASAP7_75t_L g348 ( .A(n_349), .Y(n_348) );
NAND2xp5_ASAP7_75t_L g432 ( .A(n_350), .B(n_358), .Y(n_432) );
INVx1_ASAP7_75t_L g350 ( .A(n_351), .Y(n_350) );
O2A1O1Ixp33_ASAP7_75t_L g443 ( .A1(n_352), .A2(n_367), .B(n_369), .C(n_444), .Y(n_443) );
NAND2xp5_ASAP7_75t_L g427 ( .A(n_355), .B(n_362), .Y(n_427) );
NAND2xp5_ASAP7_75t_SL g446 ( .A(n_356), .B(n_409), .Y(n_446) );
CKINVDCx16_ASAP7_75t_R g356 ( .A(n_357), .Y(n_356) );
INVxp33_ASAP7_75t_L g359 ( .A(n_360), .Y(n_359) );
NOR2xp33_ASAP7_75t_L g360 ( .A(n_361), .B(n_363), .Y(n_360) );
AOI21xp33_ASAP7_75t_SL g372 ( .A1(n_361), .A2(n_373), .B(n_375), .Y(n_372) );
NOR2xp33_ASAP7_75t_L g433 ( .A(n_361), .B(n_434), .Y(n_433) );
INVx2_ASAP7_75t_SL g361 ( .A(n_362), .Y(n_361) );
NAND2xp5_ASAP7_75t_L g415 ( .A(n_362), .B(n_416), .Y(n_415) );
AOI221xp5_ASAP7_75t_L g364 ( .A1(n_365), .A2(n_368), .B1(n_369), .B2(n_371), .C(n_372), .Y(n_364) );
INVx1_ASAP7_75t_L g365 ( .A(n_366), .Y(n_365) );
NAND2xp5_ASAP7_75t_L g417 ( .A(n_368), .B(n_418), .Y(n_417) );
INVx1_ASAP7_75t_L g369 ( .A(n_370), .Y(n_369) );
INVx1_ASAP7_75t_L g402 ( .A(n_374), .Y(n_402) );
NAND5xp2_ASAP7_75t_L g377 ( .A(n_378), .B(n_405), .C(n_419), .D(n_430), .E(n_443), .Y(n_377) );
AOI211xp5_ASAP7_75t_L g378 ( .A1(n_379), .A2(n_381), .B(n_388), .C(n_401), .Y(n_378) );
INVx2_ASAP7_75t_SL g425 ( .A(n_379), .Y(n_425) );
NAND4xp25_ASAP7_75t_SL g381 ( .A(n_382), .B(n_384), .C(n_385), .D(n_387), .Y(n_381) );
INVx1_ASAP7_75t_L g382 ( .A(n_383), .Y(n_382) );
INVx3_ASAP7_75t_L g385 ( .A(n_386), .Y(n_385) );
OAI211xp5_ASAP7_75t_SL g388 ( .A1(n_387), .A2(n_389), .B(n_392), .C(n_398), .Y(n_388) );
CKINVDCx20_ASAP7_75t_R g389 ( .A(n_390), .Y(n_389) );
AOI221xp5_ASAP7_75t_L g430 ( .A1(n_390), .A2(n_431), .B1(n_433), .B2(n_435), .C(n_437), .Y(n_430) );
INVx1_ASAP7_75t_L g393 ( .A(n_394), .Y(n_393) );
INVx1_ASAP7_75t_L g396 ( .A(n_397), .Y(n_396) );
INVx1_ASAP7_75t_L g399 ( .A(n_400), .Y(n_399) );
AOI221xp5_ASAP7_75t_SL g405 ( .A1(n_406), .A2(n_407), .B1(n_410), .B2(n_412), .C(n_414), .Y(n_405) );
AND2x2_ASAP7_75t_L g407 ( .A(n_408), .B(n_409), .Y(n_407) );
INVx1_ASAP7_75t_L g410 ( .A(n_411), .Y(n_410) );
INVx1_ASAP7_75t_L g412 ( .A(n_413), .Y(n_412) );
OAI22xp5_ASAP7_75t_L g437 ( .A1(n_413), .A2(n_436), .B1(n_438), .B2(n_440), .Y(n_437) );
INVx1_ASAP7_75t_L g414 ( .A(n_415), .Y(n_414) );
INVx1_ASAP7_75t_SL g416 ( .A(n_417), .Y(n_416) );
OAI22xp5_ASAP7_75t_L g422 ( .A1(n_423), .A2(n_425), .B1(n_426), .B2(n_427), .Y(n_422) );
INVx1_ASAP7_75t_L g431 ( .A(n_432), .Y(n_431) );
INVx1_ASAP7_75t_L g435 ( .A(n_436), .Y(n_435) );
INVx1_ASAP7_75t_SL g438 ( .A(n_439), .Y(n_438) );
NAND2xp5_ASAP7_75t_L g440 ( .A(n_441), .B(n_442), .Y(n_440) );
NAND3xp33_ASAP7_75t_L g454 ( .A(n_451), .B(n_455), .C(n_752), .Y(n_454) );
INVx1_ASAP7_75t_SL g452 ( .A(n_453), .Y(n_452) );
XOR2xp5_ASAP7_75t_L g456 ( .A(n_457), .B(n_466), .Y(n_456) );
INVx1_ASAP7_75t_L g459 ( .A(n_460), .Y(n_459) );
INVx1_ASAP7_75t_L g462 ( .A(n_463), .Y(n_462) );
OAI22xp5_ASAP7_75t_SL g466 ( .A1(n_467), .A2(n_746), .B1(n_747), .B2(n_748), .Y(n_466) );
AND2x2_ASAP7_75t_SL g467 ( .A(n_468), .B(n_715), .Y(n_467) );
NOR3xp33_ASAP7_75t_L g468 ( .A(n_469), .B(n_608), .C(n_681), .Y(n_468) );
OAI211xp5_ASAP7_75t_SL g469 ( .A1(n_470), .A2(n_502), .B(n_541), .C(n_592), .Y(n_469) );
INVxp67_ASAP7_75t_L g470 ( .A(n_471), .Y(n_470) );
AND2x2_ASAP7_75t_L g471 ( .A(n_472), .B(n_482), .Y(n_471) );
AND2x2_ASAP7_75t_L g557 ( .A(n_472), .B(n_558), .Y(n_557) );
INVx3_ASAP7_75t_L g575 ( .A(n_472), .Y(n_575) );
INVx2_ASAP7_75t_L g590 ( .A(n_472), .Y(n_590) );
INVx1_ASAP7_75t_L g620 ( .A(n_472), .Y(n_620) );
AND2x2_ASAP7_75t_L g670 ( .A(n_472), .B(n_591), .Y(n_670) );
AOI32xp33_ASAP7_75t_L g697 ( .A1(n_472), .A2(n_625), .A3(n_698), .B1(n_700), .B2(n_701), .Y(n_697) );
NAND2xp5_ASAP7_75t_L g703 ( .A(n_472), .B(n_547), .Y(n_703) );
AND2x2_ASAP7_75t_L g730 ( .A(n_472), .B(n_573), .Y(n_730) );
NOR2xp33_ASAP7_75t_L g738 ( .A(n_472), .B(n_739), .Y(n_738) );
OR2x6_ASAP7_75t_L g472 ( .A(n_473), .B(n_480), .Y(n_472) );
AND2x2_ASAP7_75t_L g619 ( .A(n_482), .B(n_620), .Y(n_619) );
INVx1_ASAP7_75t_L g641 ( .A(n_482), .Y(n_641) );
AND2x2_ASAP7_75t_L g726 ( .A(n_482), .B(n_557), .Y(n_726) );
AND2x2_ASAP7_75t_L g729 ( .A(n_482), .B(n_730), .Y(n_729) );
AND2x2_ASAP7_75t_L g482 ( .A(n_483), .B(n_493), .Y(n_482) );
INVx2_ASAP7_75t_L g549 ( .A(n_483), .Y(n_549) );
NAND2xp5_ASAP7_75t_L g579 ( .A(n_483), .B(n_573), .Y(n_579) );
AND2x2_ASAP7_75t_L g589 ( .A(n_483), .B(n_590), .Y(n_589) );
INVx1_ASAP7_75t_L g625 ( .A(n_483), .Y(n_625) );
NAND2xp5_ASAP7_75t_L g484 ( .A(n_485), .B(n_490), .Y(n_484) );
AOI21xp5_ASAP7_75t_L g486 ( .A1(n_487), .A2(n_488), .B(n_489), .Y(n_486) );
AND2x2_ASAP7_75t_L g567 ( .A(n_493), .B(n_549), .Y(n_567) );
INVx1_ASAP7_75t_L g493 ( .A(n_494), .Y(n_493) );
INVx2_ASAP7_75t_L g550 ( .A(n_494), .Y(n_550) );
AND2x2_ASAP7_75t_L g591 ( .A(n_494), .B(n_573), .Y(n_591) );
AND2x2_ASAP7_75t_L g660 ( .A(n_494), .B(n_558), .Y(n_660) );
NAND2xp5_ASAP7_75t_L g502 ( .A(n_503), .B(n_513), .Y(n_502) );
OR2x2_ASAP7_75t_L g555 ( .A(n_503), .B(n_524), .Y(n_555) );
INVx1_ASAP7_75t_L g633 ( .A(n_503), .Y(n_633) );
AND2x2_ASAP7_75t_L g647 ( .A(n_503), .B(n_648), .Y(n_647) );
NAND2xp5_ASAP7_75t_L g679 ( .A(n_503), .B(n_523), .Y(n_679) );
NAND2xp5_ASAP7_75t_L g699 ( .A(n_503), .B(n_645), .Y(n_699) );
AND2x2_ASAP7_75t_L g707 ( .A(n_503), .B(n_708), .Y(n_707) );
INVx3_ASAP7_75t_L g503 ( .A(n_504), .Y(n_503) );
INVx3_ASAP7_75t_L g545 ( .A(n_504), .Y(n_545) );
AND2x2_ASAP7_75t_L g614 ( .A(n_504), .B(n_524), .Y(n_614) );
NAND2xp5_ASAP7_75t_L g737 ( .A(n_513), .B(n_738), .Y(n_737) );
INVx2_ASAP7_75t_L g741 ( .A(n_513), .Y(n_741) );
AND2x2_ASAP7_75t_L g513 ( .A(n_514), .B(n_523), .Y(n_513) );
NAND2xp5_ASAP7_75t_L g607 ( .A(n_514), .B(n_585), .Y(n_607) );
OR2x2_ASAP7_75t_L g636 ( .A(n_514), .B(n_637), .Y(n_636) );
AND2x2_ASAP7_75t_L g668 ( .A(n_514), .B(n_648), .Y(n_668) );
INVx1_ASAP7_75t_SL g688 ( .A(n_514), .Y(n_688) );
AND2x2_ASAP7_75t_L g692 ( .A(n_514), .B(n_554), .Y(n_692) );
INVx2_ASAP7_75t_L g514 ( .A(n_515), .Y(n_514) );
AND2x2_ASAP7_75t_SL g546 ( .A(n_515), .B(n_523), .Y(n_546) );
AND2x2_ASAP7_75t_L g553 ( .A(n_515), .B(n_533), .Y(n_553) );
NAND2xp5_ASAP7_75t_L g576 ( .A(n_515), .B(n_577), .Y(n_576) );
OR2x2_ASAP7_75t_L g595 ( .A(n_515), .B(n_577), .Y(n_595) );
INVx1_ASAP7_75t_SL g602 ( .A(n_515), .Y(n_602) );
BUFx2_ASAP7_75t_L g613 ( .A(n_515), .Y(n_613) );
AND2x2_ASAP7_75t_L g629 ( .A(n_515), .B(n_545), .Y(n_629) );
AND2x2_ASAP7_75t_L g644 ( .A(n_515), .B(n_645), .Y(n_644) );
AND2x2_ASAP7_75t_L g708 ( .A(n_515), .B(n_524), .Y(n_708) );
NAND2xp5_ASAP7_75t_L g628 ( .A(n_523), .B(n_629), .Y(n_628) );
AND2x2_ASAP7_75t_L g632 ( .A(n_523), .B(n_633), .Y(n_632) );
AOI221xp5_ASAP7_75t_L g649 ( .A1(n_523), .A2(n_650), .B1(n_653), .B2(n_656), .C(n_661), .Y(n_649) );
NAND2xp5_ASAP7_75t_L g723 ( .A(n_523), .B(n_724), .Y(n_723) );
AND2x2_ASAP7_75t_L g523 ( .A(n_524), .B(n_533), .Y(n_523) );
INVx3_ASAP7_75t_L g577 ( .A(n_524), .Y(n_577) );
BUFx2_ASAP7_75t_L g587 ( .A(n_533), .Y(n_587) );
AND2x2_ASAP7_75t_L g601 ( .A(n_533), .B(n_602), .Y(n_601) );
INVx1_ASAP7_75t_L g618 ( .A(n_533), .Y(n_618) );
OR2x2_ASAP7_75t_L g637 ( .A(n_533), .B(n_577), .Y(n_637) );
INVx3_ASAP7_75t_L g645 ( .A(n_533), .Y(n_645) );
AND2x2_ASAP7_75t_L g648 ( .A(n_533), .B(n_577), .Y(n_648) );
AOI221xp5_ASAP7_75t_L g541 ( .A1(n_542), .A2(n_547), .B1(n_551), .B2(n_556), .C(n_568), .Y(n_541) );
INVx1_ASAP7_75t_L g542 ( .A(n_543), .Y(n_542) );
NAND2xp5_ASAP7_75t_L g543 ( .A(n_544), .B(n_546), .Y(n_543) );
NAND2xp5_ASAP7_75t_L g742 ( .A(n_544), .B(n_617), .Y(n_742) );
OR2x2_ASAP7_75t_L g745 ( .A(n_544), .B(n_576), .Y(n_745) );
INVx1_ASAP7_75t_SL g544 ( .A(n_545), .Y(n_544) );
OAI221xp5_ASAP7_75t_SL g568 ( .A1(n_545), .A2(n_569), .B1(n_576), .B2(n_578), .C(n_581), .Y(n_568) );
AND2x2_ASAP7_75t_L g585 ( .A(n_545), .B(n_577), .Y(n_585) );
AND2x2_ASAP7_75t_L g593 ( .A(n_545), .B(n_594), .Y(n_593) );
NAND2xp5_ASAP7_75t_L g600 ( .A(n_545), .B(n_601), .Y(n_600) );
NAND2x1_ASAP7_75t_L g643 ( .A(n_545), .B(n_644), .Y(n_643) );
OR2x2_ASAP7_75t_L g695 ( .A(n_545), .B(n_637), .Y(n_695) );
AOI22xp5_ASAP7_75t_L g683 ( .A1(n_547), .A2(n_655), .B1(n_684), .B2(n_686), .Y(n_683) );
INVx2_ASAP7_75t_L g547 ( .A(n_548), .Y(n_547) );
AOI322xp5_ASAP7_75t_L g592 ( .A1(n_548), .A2(n_557), .A3(n_593), .B1(n_596), .B2(n_599), .C1(n_603), .C2(n_606), .Y(n_592) );
OR2x2_ASAP7_75t_L g604 ( .A(n_548), .B(n_605), .Y(n_604) );
OR2x2_ASAP7_75t_L g548 ( .A(n_549), .B(n_550), .Y(n_548) );
NAND2xp5_ASAP7_75t_L g572 ( .A(n_549), .B(n_573), .Y(n_572) );
AND2x2_ASAP7_75t_L g583 ( .A(n_549), .B(n_558), .Y(n_583) );
INVx1_ASAP7_75t_L g598 ( .A(n_549), .Y(n_598) );
AND2x2_ASAP7_75t_L g664 ( .A(n_549), .B(n_665), .Y(n_664) );
AND2x2_ASAP7_75t_L g574 ( .A(n_550), .B(n_575), .Y(n_574) );
INVx2_ASAP7_75t_L g665 ( .A(n_550), .Y(n_665) );
NAND2xp5_ASAP7_75t_L g739 ( .A(n_550), .B(n_573), .Y(n_739) );
INVx1_ASAP7_75t_L g551 ( .A(n_552), .Y(n_551) );
NAND2xp5_ASAP7_75t_L g552 ( .A(n_553), .B(n_554), .Y(n_552) );
NAND2xp5_ASAP7_75t_L g687 ( .A(n_554), .B(n_688), .Y(n_687) );
INVx3_ASAP7_75t_SL g554 ( .A(n_555), .Y(n_554) );
OR2x2_ASAP7_75t_L g639 ( .A(n_555), .B(n_586), .Y(n_639) );
OR2x2_ASAP7_75t_L g736 ( .A(n_555), .B(n_587), .Y(n_736) );
INVx1_ASAP7_75t_L g717 ( .A(n_556), .Y(n_717) );
AND2x2_ASAP7_75t_L g556 ( .A(n_557), .B(n_567), .Y(n_556) );
INVx4_ASAP7_75t_L g605 ( .A(n_557), .Y(n_605) );
NAND2xp5_ASAP7_75t_L g630 ( .A(n_557), .B(n_624), .Y(n_630) );
INVx2_ASAP7_75t_L g573 ( .A(n_558), .Y(n_573) );
INVx1_ASAP7_75t_L g655 ( .A(n_567), .Y(n_655) );
NAND2xp5_ASAP7_75t_L g696 ( .A(n_567), .B(n_627), .Y(n_696) );
AOI21xp33_ASAP7_75t_L g642 ( .A1(n_569), .A2(n_643), .B(n_646), .Y(n_642) );
INVx2_ASAP7_75t_L g569 ( .A(n_570), .Y(n_569) );
AND2x2_ASAP7_75t_L g570 ( .A(n_571), .B(n_574), .Y(n_570) );
INVx1_ASAP7_75t_L g571 ( .A(n_572), .Y(n_571) );
INVx2_ASAP7_75t_L g627 ( .A(n_573), .Y(n_627) );
INVx1_ASAP7_75t_L g654 ( .A(n_573), .Y(n_654) );
INVx1_ASAP7_75t_L g580 ( .A(n_574), .Y(n_580) );
AND2x2_ASAP7_75t_L g582 ( .A(n_574), .B(n_583), .Y(n_582) );
AND2x2_ASAP7_75t_L g678 ( .A(n_575), .B(n_664), .Y(n_678) );
AND2x2_ASAP7_75t_L g700 ( .A(n_575), .B(n_660), .Y(n_700) );
BUFx2_ASAP7_75t_L g652 ( .A(n_577), .Y(n_652) );
OR2x2_ASAP7_75t_L g578 ( .A(n_579), .B(n_580), .Y(n_578) );
AOI32xp33_ASAP7_75t_L g581 ( .A1(n_582), .A2(n_584), .A3(n_585), .B1(n_586), .B2(n_588), .Y(n_581) );
INVx1_ASAP7_75t_L g662 ( .A(n_582), .Y(n_662) );
AOI22xp33_ASAP7_75t_L g709 ( .A1(n_582), .A2(n_710), .B1(n_711), .B2(n_713), .Y(n_709) );
INVx1_ASAP7_75t_L g584 ( .A(n_585), .Y(n_584) );
NOR2xp33_ASAP7_75t_L g615 ( .A(n_585), .B(n_616), .Y(n_615) );
NAND2xp5_ASAP7_75t_L g685 ( .A(n_585), .B(n_644), .Y(n_685) );
AND2x2_ASAP7_75t_L g732 ( .A(n_585), .B(n_617), .Y(n_732) );
NAND2xp5_ASAP7_75t_L g680 ( .A(n_586), .B(n_633), .Y(n_680) );
INVx1_ASAP7_75t_L g586 ( .A(n_587), .Y(n_586) );
INVx1_ASAP7_75t_L g733 ( .A(n_588), .Y(n_733) );
AND2x2_ASAP7_75t_L g588 ( .A(n_589), .B(n_591), .Y(n_588) );
INVx1_ASAP7_75t_L g658 ( .A(n_589), .Y(n_658) );
NAND2xp5_ASAP7_75t_L g597 ( .A(n_591), .B(n_598), .Y(n_597) );
AND2x2_ASAP7_75t_L g705 ( .A(n_591), .B(n_625), .Y(n_705) );
NAND2xp5_ASAP7_75t_L g712 ( .A(n_591), .B(n_620), .Y(n_712) );
INVx1_ASAP7_75t_SL g694 ( .A(n_593), .Y(n_694) );
NAND2xp5_ASAP7_75t_L g672 ( .A(n_594), .B(n_645), .Y(n_672) );
NOR4xp25_ASAP7_75t_L g718 ( .A(n_594), .B(n_617), .C(n_719), .D(n_722), .Y(n_718) );
INVx1_ASAP7_75t_L g594 ( .A(n_595), .Y(n_594) );
NOR2xp33_ASAP7_75t_L g698 ( .A(n_595), .B(n_699), .Y(n_698) );
INVx1_ASAP7_75t_L g596 ( .A(n_597), .Y(n_596) );
INVxp67_ASAP7_75t_L g675 ( .A(n_598), .Y(n_675) );
INVx1_ASAP7_75t_L g599 ( .A(n_600), .Y(n_599) );
OAI21xp33_ASAP7_75t_L g725 ( .A1(n_601), .A2(n_692), .B(n_726), .Y(n_725) );
AND2x4_ASAP7_75t_L g617 ( .A(n_602), .B(n_618), .Y(n_617) );
INVx1_ASAP7_75t_L g603 ( .A(n_604), .Y(n_603) );
INVx1_ASAP7_75t_L g666 ( .A(n_605), .Y(n_666) );
INVx1_ASAP7_75t_L g606 ( .A(n_607), .Y(n_606) );
NAND4xp25_ASAP7_75t_SL g608 ( .A(n_609), .B(n_634), .C(n_649), .D(n_669), .Y(n_608) );
O2A1O1Ixp33_ASAP7_75t_L g609 ( .A1(n_610), .A2(n_615), .B(n_619), .C(n_621), .Y(n_609) );
INVx1_ASAP7_75t_SL g610 ( .A(n_611), .Y(n_610) );
NAND2xp5_ASAP7_75t_L g611 ( .A(n_612), .B(n_614), .Y(n_611) );
INVx1_ASAP7_75t_SL g612 ( .A(n_613), .Y(n_612) );
AND2x2_ASAP7_75t_L g701 ( .A(n_614), .B(n_644), .Y(n_701) );
AND2x2_ASAP7_75t_L g710 ( .A(n_614), .B(n_688), .Y(n_710) );
INVx3_ASAP7_75t_SL g616 ( .A(n_617), .Y(n_616) );
NAND2xp5_ASAP7_75t_L g714 ( .A(n_617), .B(n_652), .Y(n_714) );
AND2x2_ASAP7_75t_L g626 ( .A(n_620), .B(n_627), .Y(n_626) );
OAI22xp5_ASAP7_75t_L g621 ( .A1(n_622), .A2(n_628), .B1(n_630), .B2(n_631), .Y(n_621) );
INVx1_ASAP7_75t_L g622 ( .A(n_623), .Y(n_622) );
AND2x2_ASAP7_75t_L g623 ( .A(n_624), .B(n_626), .Y(n_623) );
AND2x2_ASAP7_75t_L g724 ( .A(n_624), .B(n_670), .Y(n_724) );
INVx1_ASAP7_75t_L g624 ( .A(n_625), .Y(n_624) );
NAND2xp5_ASAP7_75t_L g691 ( .A(n_626), .B(n_675), .Y(n_691) );
NOR2xp33_ASAP7_75t_L g640 ( .A(n_627), .B(n_641), .Y(n_640) );
INVx1_ASAP7_75t_L g631 ( .A(n_632), .Y(n_631) );
O2A1O1Ixp33_ASAP7_75t_L g634 ( .A1(n_635), .A2(n_638), .B(n_640), .C(n_642), .Y(n_634) );
AOI221xp5_ASAP7_75t_L g669 ( .A1(n_635), .A2(n_670), .B1(n_671), .B2(n_673), .C(n_676), .Y(n_669) );
INVx1_ASAP7_75t_SL g635 ( .A(n_636), .Y(n_635) );
INVx1_ASAP7_75t_L g638 ( .A(n_639), .Y(n_638) );
OAI221xp5_ASAP7_75t_L g727 ( .A1(n_643), .A2(n_728), .B1(n_731), .B2(n_733), .C(n_734), .Y(n_727) );
NAND2xp5_ASAP7_75t_L g651 ( .A(n_644), .B(n_652), .Y(n_651) );
INVx1_ASAP7_75t_SL g646 ( .A(n_647), .Y(n_646) );
INVx1_ASAP7_75t_L g650 ( .A(n_651), .Y(n_650) );
NAND2xp5_ASAP7_75t_L g720 ( .A(n_652), .B(n_721), .Y(n_720) );
NOR2xp33_ASAP7_75t_L g653 ( .A(n_654), .B(n_655), .Y(n_653) );
INVx1_ASAP7_75t_L g682 ( .A(n_654), .Y(n_682) );
INVx1_ASAP7_75t_SL g656 ( .A(n_657), .Y(n_656) );
OAI22xp5_ASAP7_75t_L g676 ( .A1(n_657), .A2(n_677), .B1(n_679), .B2(n_680), .Y(n_676) );
OR2x2_ASAP7_75t_L g657 ( .A(n_658), .B(n_659), .Y(n_657) );
INVx1_ASAP7_75t_L g659 ( .A(n_660), .Y(n_659) );
AOI21xp33_ASAP7_75t_L g661 ( .A1(n_662), .A2(n_663), .B(n_667), .Y(n_661) );
NAND2xp5_ASAP7_75t_L g663 ( .A(n_664), .B(n_666), .Y(n_663) );
NAND2xp5_ASAP7_75t_L g674 ( .A(n_666), .B(n_675), .Y(n_674) );
INVx1_ASAP7_75t_L g667 ( .A(n_668), .Y(n_667) );
INVx1_ASAP7_75t_L g671 ( .A(n_672), .Y(n_671) );
INVx1_ASAP7_75t_L g673 ( .A(n_674), .Y(n_673) );
OAI221xp5_ASAP7_75t_L g740 ( .A1(n_677), .A2(n_703), .B1(n_741), .B2(n_742), .C(n_743), .Y(n_740) );
INVx1_ASAP7_75t_L g677 ( .A(n_678), .Y(n_677) );
INVx1_ASAP7_75t_L g722 ( .A(n_679), .Y(n_722) );
OAI211xp5_ASAP7_75t_SL g681 ( .A1(n_682), .A2(n_683), .B(n_689), .C(n_709), .Y(n_681) );
INVx1_ASAP7_75t_L g684 ( .A(n_685), .Y(n_684) );
INVx1_ASAP7_75t_L g686 ( .A(n_687), .Y(n_686) );
AOI211xp5_ASAP7_75t_L g689 ( .A1(n_690), .A2(n_692), .B(n_693), .C(n_702), .Y(n_689) );
INVx1_ASAP7_75t_L g690 ( .A(n_691), .Y(n_690) );
A2O1A1Ixp33_ASAP7_75t_L g693 ( .A1(n_694), .A2(n_695), .B(n_696), .C(n_697), .Y(n_693) );
INVx1_ASAP7_75t_L g721 ( .A(n_699), .Y(n_721) );
OAI21xp5_ASAP7_75t_SL g743 ( .A1(n_700), .A2(n_726), .B(n_744), .Y(n_743) );
AOI21xp33_ASAP7_75t_L g702 ( .A1(n_703), .A2(n_704), .B(n_706), .Y(n_702) );
INVx1_ASAP7_75t_SL g704 ( .A(n_705), .Y(n_704) );
INVxp67_ASAP7_75t_L g706 ( .A(n_707), .Y(n_706) );
INVx1_ASAP7_75t_L g711 ( .A(n_712), .Y(n_711) );
OAI21xp5_ASAP7_75t_SL g735 ( .A1(n_712), .A2(n_736), .B(n_737), .Y(n_735) );
INVx1_ASAP7_75t_L g713 ( .A(n_714), .Y(n_713) );
NOR3xp33_ASAP7_75t_L g715 ( .A(n_716), .B(n_727), .C(n_740), .Y(n_715) );
OAI211xp5_ASAP7_75t_L g716 ( .A1(n_717), .A2(n_718), .B(n_723), .C(n_725), .Y(n_716) );
INVx1_ASAP7_75t_L g719 ( .A(n_720), .Y(n_719) );
CKINVDCx14_ASAP7_75t_R g728 ( .A(n_729), .Y(n_728) );
INVx2_ASAP7_75t_L g731 ( .A(n_732), .Y(n_731) );
INVx1_ASAP7_75t_L g734 ( .A(n_735), .Y(n_734) );
INVx1_ASAP7_75t_L g744 ( .A(n_745), .Y(n_744) );
INVx1_ASAP7_75t_L g746 ( .A(n_747), .Y(n_746) );
INVx1_ASAP7_75t_L g749 ( .A(n_750), .Y(n_749) );
INVx2_ASAP7_75t_L g750 ( .A(n_751), .Y(n_750) );
CKINVDCx20_ASAP7_75t_R g752 ( .A(n_753), .Y(n_752) );
endmodule