module fake_netlist_5_135_n_1281 (n_137, n_294, n_318, n_380, n_82, n_194, n_316, n_248, n_124, n_86, n_136, n_146, n_315, n_268, n_61, n_376, n_127, n_75, n_235, n_226, n_74, n_57, n_353, n_351, n_367, n_111, n_155, n_43, n_116, n_22, n_284, n_46, n_245, n_21, n_139, n_38, n_105, n_280, n_4, n_378, n_17, n_382, n_254, n_33, n_23, n_302, n_265, n_293, n_372, n_244, n_47, n_173, n_198, n_247, n_314, n_368, n_8, n_321, n_292, n_100, n_212, n_385, n_119, n_275, n_252, n_26, n_295, n_133, n_330, n_2, n_6, n_39, n_147, n_373, n_67, n_307, n_87, n_150, n_106, n_209, n_259, n_375, n_301, n_68, n_93, n_186, n_134, n_191, n_51, n_63, n_171, n_153, n_341, n_204, n_250, n_260, n_298, n_320, n_286, n_122, n_282, n_331, n_10, n_24, n_325, n_132, n_90, n_101, n_281, n_240, n_381, n_189, n_220, n_291, n_231, n_257, n_31, n_13, n_371, n_152, n_317, n_9, n_323, n_195, n_42, n_356, n_227, n_45, n_271, n_94, n_335, n_123, n_370, n_167, n_234, n_343, n_308, n_379, n_267, n_297, n_156, n_5, n_225, n_377, n_219, n_157, n_131, n_192, n_223, n_158, n_138, n_264, n_109, n_387, n_374, n_163, n_276, n_339, n_95, n_183, n_185, n_243, n_347, n_169, n_59, n_255, n_215, n_350, n_196, n_211, n_218, n_181, n_3, n_290, n_221, n_178, n_386, n_287, n_344, n_72, n_104, n_41, n_56, n_141, n_355, n_15, n_336, n_145, n_48, n_50, n_337, n_313, n_88, n_216, n_168, n_164, n_311, n_208, n_142, n_214, n_328, n_140, n_299, n_303, n_369, n_296, n_241, n_357, n_184, n_65, n_78, n_144, n_114, n_96, n_165, n_213, n_129, n_342, n_98, n_361, n_363, n_197, n_107, n_69, n_236, n_388, n_1, n_249, n_304, n_329, n_203, n_274, n_384, n_80, n_35, n_73, n_277, n_92, n_19, n_338, n_149, n_333, n_309, n_30, n_14, n_84, n_130, n_322, n_258, n_29, n_79, n_151, n_25, n_306, n_288, n_188, n_190, n_201, n_263, n_44, n_224, n_40, n_34, n_228, n_283, n_383, n_112, n_85, n_239, n_55, n_49, n_310, n_54, n_12, n_76, n_358, n_362, n_170, n_332, n_27, n_77, n_102, n_161, n_273, n_349, n_270, n_230, n_81, n_118, n_279, n_70, n_253, n_261, n_174, n_289, n_172, n_206, n_217, n_312, n_345, n_210, n_365, n_91, n_176, n_182, n_143, n_83, n_354, n_237, n_180, n_340, n_207, n_37, n_346, n_229, n_108, n_66, n_177, n_60, n_16, n_0, n_58, n_18, n_359, n_117, n_326, n_233, n_205, n_366, n_113, n_246, n_179, n_125, n_269, n_128, n_285, n_120, n_232, n_327, n_135, n_126, n_202, n_266, n_272, n_193, n_251, n_352, n_53, n_160, n_154, n_62, n_148, n_71, n_300, n_159, n_334, n_175, n_262, n_238, n_99, n_319, n_364, n_20, n_121, n_242, n_360, n_36, n_200, n_162, n_64, n_222, n_28, n_89, n_115, n_324, n_199, n_187, n_32, n_103, n_348, n_97, n_166, n_11, n_7, n_256, n_305, n_52, n_278, n_110, n_1281);

input n_137;
input n_294;
input n_318;
input n_380;
input n_82;
input n_194;
input n_316;
input n_248;
input n_124;
input n_86;
input n_136;
input n_146;
input n_315;
input n_268;
input n_61;
input n_376;
input n_127;
input n_75;
input n_235;
input n_226;
input n_74;
input n_57;
input n_353;
input n_351;
input n_367;
input n_111;
input n_155;
input n_43;
input n_116;
input n_22;
input n_284;
input n_46;
input n_245;
input n_21;
input n_139;
input n_38;
input n_105;
input n_280;
input n_4;
input n_378;
input n_17;
input n_382;
input n_254;
input n_33;
input n_23;
input n_302;
input n_265;
input n_293;
input n_372;
input n_244;
input n_47;
input n_173;
input n_198;
input n_247;
input n_314;
input n_368;
input n_8;
input n_321;
input n_292;
input n_100;
input n_212;
input n_385;
input n_119;
input n_275;
input n_252;
input n_26;
input n_295;
input n_133;
input n_330;
input n_2;
input n_6;
input n_39;
input n_147;
input n_373;
input n_67;
input n_307;
input n_87;
input n_150;
input n_106;
input n_209;
input n_259;
input n_375;
input n_301;
input n_68;
input n_93;
input n_186;
input n_134;
input n_191;
input n_51;
input n_63;
input n_171;
input n_153;
input n_341;
input n_204;
input n_250;
input n_260;
input n_298;
input n_320;
input n_286;
input n_122;
input n_282;
input n_331;
input n_10;
input n_24;
input n_325;
input n_132;
input n_90;
input n_101;
input n_281;
input n_240;
input n_381;
input n_189;
input n_220;
input n_291;
input n_231;
input n_257;
input n_31;
input n_13;
input n_371;
input n_152;
input n_317;
input n_9;
input n_323;
input n_195;
input n_42;
input n_356;
input n_227;
input n_45;
input n_271;
input n_94;
input n_335;
input n_123;
input n_370;
input n_167;
input n_234;
input n_343;
input n_308;
input n_379;
input n_267;
input n_297;
input n_156;
input n_5;
input n_225;
input n_377;
input n_219;
input n_157;
input n_131;
input n_192;
input n_223;
input n_158;
input n_138;
input n_264;
input n_109;
input n_387;
input n_374;
input n_163;
input n_276;
input n_339;
input n_95;
input n_183;
input n_185;
input n_243;
input n_347;
input n_169;
input n_59;
input n_255;
input n_215;
input n_350;
input n_196;
input n_211;
input n_218;
input n_181;
input n_3;
input n_290;
input n_221;
input n_178;
input n_386;
input n_287;
input n_344;
input n_72;
input n_104;
input n_41;
input n_56;
input n_141;
input n_355;
input n_15;
input n_336;
input n_145;
input n_48;
input n_50;
input n_337;
input n_313;
input n_88;
input n_216;
input n_168;
input n_164;
input n_311;
input n_208;
input n_142;
input n_214;
input n_328;
input n_140;
input n_299;
input n_303;
input n_369;
input n_296;
input n_241;
input n_357;
input n_184;
input n_65;
input n_78;
input n_144;
input n_114;
input n_96;
input n_165;
input n_213;
input n_129;
input n_342;
input n_98;
input n_361;
input n_363;
input n_197;
input n_107;
input n_69;
input n_236;
input n_388;
input n_1;
input n_249;
input n_304;
input n_329;
input n_203;
input n_274;
input n_384;
input n_80;
input n_35;
input n_73;
input n_277;
input n_92;
input n_19;
input n_338;
input n_149;
input n_333;
input n_309;
input n_30;
input n_14;
input n_84;
input n_130;
input n_322;
input n_258;
input n_29;
input n_79;
input n_151;
input n_25;
input n_306;
input n_288;
input n_188;
input n_190;
input n_201;
input n_263;
input n_44;
input n_224;
input n_40;
input n_34;
input n_228;
input n_283;
input n_383;
input n_112;
input n_85;
input n_239;
input n_55;
input n_49;
input n_310;
input n_54;
input n_12;
input n_76;
input n_358;
input n_362;
input n_170;
input n_332;
input n_27;
input n_77;
input n_102;
input n_161;
input n_273;
input n_349;
input n_270;
input n_230;
input n_81;
input n_118;
input n_279;
input n_70;
input n_253;
input n_261;
input n_174;
input n_289;
input n_172;
input n_206;
input n_217;
input n_312;
input n_345;
input n_210;
input n_365;
input n_91;
input n_176;
input n_182;
input n_143;
input n_83;
input n_354;
input n_237;
input n_180;
input n_340;
input n_207;
input n_37;
input n_346;
input n_229;
input n_108;
input n_66;
input n_177;
input n_60;
input n_16;
input n_0;
input n_58;
input n_18;
input n_359;
input n_117;
input n_326;
input n_233;
input n_205;
input n_366;
input n_113;
input n_246;
input n_179;
input n_125;
input n_269;
input n_128;
input n_285;
input n_120;
input n_232;
input n_327;
input n_135;
input n_126;
input n_202;
input n_266;
input n_272;
input n_193;
input n_251;
input n_352;
input n_53;
input n_160;
input n_154;
input n_62;
input n_148;
input n_71;
input n_300;
input n_159;
input n_334;
input n_175;
input n_262;
input n_238;
input n_99;
input n_319;
input n_364;
input n_20;
input n_121;
input n_242;
input n_360;
input n_36;
input n_200;
input n_162;
input n_64;
input n_222;
input n_28;
input n_89;
input n_115;
input n_324;
input n_199;
input n_187;
input n_32;
input n_103;
input n_348;
input n_97;
input n_166;
input n_11;
input n_7;
input n_256;
input n_305;
input n_52;
input n_278;
input n_110;

output n_1281;

wire n_924;
wire n_1263;
wire n_977;
wire n_611;
wire n_1126;
wire n_1166;
wire n_469;
wire n_785;
wire n_549;
wire n_532;
wire n_1161;
wire n_1150;
wire n_667;
wire n_790;
wire n_1055;
wire n_880;
wire n_544;
wire n_1007;
wire n_552;
wire n_1198;
wire n_1099;
wire n_956;
wire n_564;
wire n_423;
wire n_1021;
wire n_551;
wire n_688;
wire n_800;
wire n_671;
wire n_819;
wire n_1022;
wire n_915;
wire n_864;
wire n_859;
wire n_951;
wire n_1264;
wire n_447;
wire n_625;
wire n_854;
wire n_674;
wire n_417;
wire n_516;
wire n_933;
wire n_1152;
wire n_497;
wire n_606;
wire n_877;
wire n_755;
wire n_1118;
wire n_947;
wire n_530;
wire n_1107;
wire n_556;
wire n_1230;
wire n_668;
wire n_929;
wire n_1124;
wire n_902;
wire n_1104;
wire n_659;
wire n_1257;
wire n_1182;
wire n_579;
wire n_1261;
wire n_938;
wire n_1098;
wire n_1154;
wire n_1242;
wire n_1135;
wire n_519;
wire n_406;
wire n_1016;
wire n_1243;
wire n_546;
wire n_1280;
wire n_731;
wire n_709;
wire n_1236;
wire n_569;
wire n_920;
wire n_976;
wire n_1078;
wire n_775;
wire n_600;
wire n_955;
wire n_1146;
wire n_882;
wire n_1036;
wire n_1097;
wire n_550;
wire n_696;
wire n_897;
wire n_798;
wire n_646;
wire n_436;
wire n_1216;
wire n_580;
wire n_1040;
wire n_578;
wire n_926;
wire n_1218;
wire n_422;
wire n_475;
wire n_777;
wire n_1070;
wire n_1030;
wire n_415;
wire n_1071;
wire n_485;
wire n_1165;
wire n_1267;
wire n_496;
wire n_958;
wire n_1034;
wire n_670;
wire n_521;
wire n_663;
wire n_845;
wire n_673;
wire n_837;
wire n_1239;
wire n_528;
wire n_680;
wire n_395;
wire n_553;
wire n_901;
wire n_813;
wire n_675;
wire n_888;
wire n_1167;
wire n_637;
wire n_446;
wire n_1064;
wire n_858;
wire n_923;
wire n_691;
wire n_1151;
wire n_881;
wire n_468;
wire n_464;
wire n_1069;
wire n_1075;
wire n_460;
wire n_889;
wire n_973;
wire n_477;
wire n_571;
wire n_461;
wire n_1211;
wire n_1197;
wire n_907;
wire n_989;
wire n_1039;
wire n_488;
wire n_736;
wire n_892;
wire n_1000;
wire n_1202;
wire n_1278;
wire n_1002;
wire n_593;
wire n_748;
wire n_586;
wire n_1058;
wire n_838;
wire n_1053;
wire n_1224;
wire n_1248;
wire n_953;
wire n_1014;
wire n_1241;
wire n_963;
wire n_1052;
wire n_954;
wire n_627;
wire n_440;
wire n_793;
wire n_478;
wire n_476;
wire n_534;
wire n_884;
wire n_944;
wire n_647;
wire n_407;
wire n_1072;
wire n_832;
wire n_857;
wire n_561;
wire n_1027;
wire n_971;
wire n_1156;
wire n_794;
wire n_404;
wire n_686;
wire n_847;
wire n_596;
wire n_558;
wire n_702;
wire n_1276;
wire n_822;
wire n_728;
wire n_1162;
wire n_1199;
wire n_1038;
wire n_520;
wire n_409;
wire n_887;
wire n_809;
wire n_931;
wire n_870;
wire n_599;
wire n_434;
wire n_868;
wire n_639;
wire n_914;
wire n_411;
wire n_414;
wire n_965;
wire n_935;
wire n_817;
wire n_1175;
wire n_759;
wire n_806;
wire n_1189;
wire n_1259;
wire n_706;
wire n_746;
wire n_747;
wire n_784;
wire n_1244;
wire n_431;
wire n_1194;
wire n_615;
wire n_851;
wire n_843;
wire n_523;
wire n_913;
wire n_705;
wire n_865;
wire n_678;
wire n_697;
wire n_1222;
wire n_776;
wire n_452;
wire n_525;
wire n_1260;
wire n_649;
wire n_547;
wire n_1191;
wire n_1128;
wire n_744;
wire n_629;
wire n_590;
wire n_1233;
wire n_526;
wire n_677;
wire n_1121;
wire n_433;
wire n_604;
wire n_949;
wire n_1008;
wire n_946;
wire n_1001;
wire n_498;
wire n_689;
wire n_738;
wire n_640;
wire n_624;
wire n_1010;
wire n_1231;
wire n_739;
wire n_1279;
wire n_1195;
wire n_610;
wire n_936;
wire n_568;
wire n_1090;
wire n_757;
wire n_633;
wire n_439;
wire n_448;
wire n_758;
wire n_999;
wire n_1158;
wire n_563;
wire n_1145;
wire n_878;
wire n_524;
wire n_394;
wire n_1049;
wire n_1153;
wire n_741;
wire n_1068;
wire n_906;
wire n_1163;
wire n_1207;
wire n_919;
wire n_908;
wire n_724;
wire n_658;
wire n_456;
wire n_959;
wire n_535;
wire n_940;
wire n_592;
wire n_1169;
wire n_1017;
wire n_978;
wire n_1054;
wire n_1269;
wire n_1095;
wire n_514;
wire n_457;
wire n_1079;
wire n_1045;
wire n_1208;
wire n_603;
wire n_484;
wire n_1033;
wire n_442;
wire n_636;
wire n_660;
wire n_1009;
wire n_1148;
wire n_742;
wire n_750;
wire n_995;
wire n_454;
wire n_396;
wire n_1073;
wire n_662;
wire n_459;
wire n_962;
wire n_1215;
wire n_1171;
wire n_723;
wire n_1065;
wire n_473;
wire n_1043;
wire n_486;
wire n_614;
wire n_1177;
wire n_974;
wire n_727;
wire n_1159;
wire n_957;
wire n_773;
wire n_743;
wire n_613;
wire n_1119;
wire n_1240;
wire n_829;
wire n_1237;
wire n_700;
wire n_573;
wire n_1132;
wire n_1127;
wire n_761;
wire n_1006;
wire n_1270;
wire n_582;
wire n_512;
wire n_1249;
wire n_652;
wire n_1111;
wire n_1093;
wire n_1031;
wire n_609;
wire n_1041;
wire n_1265;
wire n_834;
wire n_765;
wire n_893;
wire n_1015;
wire n_1140;
wire n_891;
wire n_630;
wire n_504;
wire n_511;
wire n_874;
wire n_1101;
wire n_1106;
wire n_987;
wire n_767;
wire n_993;
wire n_545;
wire n_441;
wire n_860;
wire n_450;
wire n_429;
wire n_948;
wire n_1217;
wire n_628;
wire n_729;
wire n_1131;
wire n_1084;
wire n_970;
wire n_911;
wire n_513;
wire n_1094;
wire n_560;
wire n_1044;
wire n_1205;
wire n_1209;
wire n_495;
wire n_602;
wire n_574;
wire n_879;
wire n_623;
wire n_405;
wire n_824;
wire n_490;
wire n_996;
wire n_921;
wire n_572;
wire n_815;
wire n_1037;
wire n_1080;
wire n_1274;
wire n_426;
wire n_1082;
wire n_589;
wire n_716;
wire n_562;
wire n_952;
wire n_1229;
wire n_391;
wire n_701;
wire n_1023;
wire n_645;
wire n_539;
wire n_803;
wire n_1092;
wire n_531;
wire n_890;
wire n_764;
wire n_1056;
wire n_960;
wire n_1123;
wire n_1047;
wire n_634;
wire n_1252;
wire n_1029;
wire n_925;
wire n_1206;
wire n_424;
wire n_950;
wire n_419;
wire n_444;
wire n_1060;
wire n_1141;
wire n_389;
wire n_418;
wire n_968;
wire n_912;
wire n_451;
wire n_619;
wire n_408;
wire n_967;
wire n_1139;
wire n_515;
wire n_885;
wire n_397;
wire n_483;
wire n_683;
wire n_1057;
wire n_1051;
wire n_1085;
wire n_1066;
wire n_721;
wire n_1157;
wire n_841;
wire n_1050;
wire n_802;
wire n_983;
wire n_873;
wire n_1112;
wire n_762;
wire n_690;
wire n_583;
wire n_1203;
wire n_821;
wire n_1179;
wire n_621;
wire n_753;
wire n_455;
wire n_1048;
wire n_507;
wire n_1228;
wire n_972;
wire n_692;
wire n_820;
wire n_1200;
wire n_1185;
wire n_991;
wire n_828;
wire n_779;
wire n_576;
wire n_1143;
wire n_804;
wire n_537;
wire n_945;
wire n_492;
wire n_943;
wire n_992;
wire n_543;
wire n_842;
wire n_650;
wire n_984;
wire n_694;
wire n_883;
wire n_470;
wire n_449;
wire n_1214;
wire n_900;
wire n_856;
wire n_918;
wire n_942;
wire n_1147;
wire n_1077;
wire n_540;
wire n_618;
wire n_896;
wire n_894;
wire n_831;
wire n_964;
wire n_1096;
wire n_833;
wire n_988;
wire n_814;
wire n_1201;
wire n_1114;
wire n_655;
wire n_669;
wire n_472;
wire n_1176;
wire n_1149;
wire n_398;
wire n_635;
wire n_763;
wire n_1020;
wire n_1062;
wire n_1219;
wire n_1204;
wire n_1035;
wire n_555;
wire n_783;
wire n_1188;
wire n_661;
wire n_849;
wire n_584;
wire n_681;
wire n_430;
wire n_510;
wire n_830;
wire n_801;
wire n_875;
wire n_1110;
wire n_445;
wire n_749;
wire n_1134;
wire n_717;
wire n_939;
wire n_482;
wire n_1088;
wire n_588;
wire n_1173;
wire n_789;
wire n_1232;
wire n_734;
wire n_638;
wire n_866;
wire n_969;
wire n_1019;
wire n_1105;
wire n_577;
wire n_693;
wire n_836;
wire n_990;
wire n_975;
wire n_1256;
wire n_567;
wire n_778;
wire n_1122;
wire n_458;
wire n_770;
wire n_1102;
wire n_711;
wire n_1187;
wire n_1164;
wire n_489;
wire n_1174;
wire n_617;
wire n_876;
wire n_1190;
wire n_601;
wire n_917;
wire n_966;
wire n_1116;
wire n_1212;
wire n_726;
wire n_982;
wire n_818;
wire n_861;
wire n_1183;
wire n_899;
wire n_1253;
wire n_774;
wire n_1059;
wire n_1133;
wire n_557;
wire n_1005;
wire n_607;
wire n_1003;
wire n_679;
wire n_710;
wire n_527;
wire n_1168;
wire n_707;
wire n_937;
wire n_393;
wire n_487;
wire n_665;
wire n_421;
wire n_910;
wire n_768;
wire n_1136;
wire n_754;
wire n_1125;
wire n_410;
wire n_708;
wire n_529;
wire n_735;
wire n_1109;
wire n_895;
wire n_427;
wire n_791;
wire n_732;
wire n_808;
wire n_797;
wire n_1025;
wire n_500;
wire n_1067;
wire n_435;
wire n_766;
wire n_541;
wire n_538;
wire n_1117;
wire n_799;
wire n_687;
wire n_715;
wire n_1213;
wire n_1266;
wire n_536;
wire n_872;
wire n_594;
wire n_1155;
wire n_1011;
wire n_1184;
wire n_985;
wire n_869;
wire n_810;
wire n_416;
wire n_827;
wire n_401;
wire n_626;
wire n_1144;
wire n_1137;
wire n_1170;
wire n_676;
wire n_653;
wire n_642;
wire n_855;
wire n_1178;
wire n_850;
wire n_684;
wire n_664;
wire n_503;
wire n_605;
wire n_1273;
wire n_620;
wire n_643;
wire n_916;
wire n_1081;
wire n_493;
wire n_1235;
wire n_703;
wire n_698;
wire n_980;
wire n_1115;
wire n_780;
wire n_998;
wire n_467;
wire n_1227;
wire n_840;
wire n_501;
wire n_823;
wire n_725;
wire n_672;
wire n_581;
wire n_554;
wire n_898;
wire n_1013;
wire n_718;
wire n_1120;
wire n_719;
wire n_443;
wire n_714;
wire n_909;
wire n_997;
wire n_932;
wire n_612;
wire n_788;
wire n_1268;
wire n_559;
wire n_825;
wire n_508;
wire n_506;
wire n_737;
wire n_986;
wire n_509;
wire n_1192;
wire n_1024;
wire n_1063;
wire n_733;
wire n_941;
wire n_981;
wire n_867;
wire n_587;
wire n_792;
wire n_756;
wire n_399;
wire n_1238;
wire n_548;
wire n_812;
wire n_518;
wire n_505;
wire n_752;
wire n_905;
wire n_1108;
wire n_782;
wire n_1100;
wire n_862;
wire n_760;
wire n_390;
wire n_481;
wire n_769;
wire n_1046;
wire n_934;
wire n_826;
wire n_886;
wire n_1221;
wire n_654;
wire n_1172;
wire n_428;
wire n_570;
wire n_853;
wire n_751;
wire n_786;
wire n_1083;
wire n_1142;
wire n_1129;
wire n_392;
wire n_704;
wire n_787;
wire n_961;
wire n_771;
wire n_1225;
wire n_522;
wire n_1262;
wire n_400;
wire n_930;
wire n_622;
wire n_1087;
wire n_994;
wire n_848;
wire n_1223;
wire n_1272;
wire n_682;
wire n_1247;
wire n_922;
wire n_816;
wire n_591;
wire n_631;
wire n_479;
wire n_1246;
wire n_432;
wire n_839;
wire n_1210;
wire n_1250;
wire n_871;
wire n_685;
wire n_598;
wire n_608;
wire n_928;
wire n_772;
wire n_499;
wire n_517;
wire n_413;
wire n_402;
wire n_1086;
wire n_796;
wire n_1012;
wire n_903;
wire n_740;
wire n_1061;
wire n_462;
wire n_1193;
wire n_1255;
wire n_1113;
wire n_1226;
wire n_722;
wire n_1277;
wire n_844;
wire n_471;
wire n_852;
wire n_1028;
wire n_781;
wire n_474;
wire n_542;
wire n_463;
wire n_595;
wire n_502;
wire n_466;
wire n_420;
wire n_632;
wire n_699;
wire n_979;
wire n_1245;
wire n_846;
wire n_465;
wire n_585;
wire n_616;
wire n_745;
wire n_1103;
wire n_648;
wire n_1076;
wire n_1091;
wire n_494;
wire n_641;
wire n_730;
wire n_575;
wire n_480;
wire n_425;
wire n_795;
wire n_695;
wire n_656;
wire n_1220;
wire n_437;
wire n_403;
wire n_453;
wire n_1130;
wire n_720;
wire n_863;
wire n_805;
wire n_1275;
wire n_712;
wire n_1042;
wire n_412;
wire n_657;
wire n_644;
wire n_1160;
wire n_491;
wire n_1258;
wire n_1074;
wire n_566;
wire n_565;
wire n_597;
wire n_1181;
wire n_1196;
wire n_651;
wire n_811;
wire n_807;
wire n_835;
wire n_666;
wire n_1254;
wire n_1026;
wire n_1234;
wire n_1138;
wire n_927;
wire n_1089;
wire n_1004;
wire n_1186;
wire n_1032;
wire n_1018;
wire n_438;
wire n_713;
wire n_904;
wire n_1180;
wire n_1271;
wire n_533;
wire n_1251;

CKINVDCx5p33_ASAP7_75t_R g389 ( 
.A(n_316),
.Y(n_389)
);

INVx1_ASAP7_75t_SL g390 ( 
.A(n_130),
.Y(n_390)
);

INVx2_ASAP7_75t_L g391 ( 
.A(n_152),
.Y(n_391)
);

CKINVDCx5p33_ASAP7_75t_R g392 ( 
.A(n_226),
.Y(n_392)
);

HB1xp67_ASAP7_75t_L g393 ( 
.A(n_111),
.Y(n_393)
);

CKINVDCx5p33_ASAP7_75t_R g394 ( 
.A(n_329),
.Y(n_394)
);

CKINVDCx5p33_ASAP7_75t_R g395 ( 
.A(n_158),
.Y(n_395)
);

CKINVDCx5p33_ASAP7_75t_R g396 ( 
.A(n_301),
.Y(n_396)
);

NOR2xp67_ASAP7_75t_L g397 ( 
.A(n_193),
.B(n_213),
.Y(n_397)
);

INVx1_ASAP7_75t_L g398 ( 
.A(n_381),
.Y(n_398)
);

CKINVDCx20_ASAP7_75t_R g399 ( 
.A(n_123),
.Y(n_399)
);

INVx2_ASAP7_75t_L g400 ( 
.A(n_208),
.Y(n_400)
);

CKINVDCx5p33_ASAP7_75t_R g401 ( 
.A(n_339),
.Y(n_401)
);

CKINVDCx5p33_ASAP7_75t_R g402 ( 
.A(n_140),
.Y(n_402)
);

CKINVDCx20_ASAP7_75t_R g403 ( 
.A(n_181),
.Y(n_403)
);

INVx2_ASAP7_75t_L g404 ( 
.A(n_242),
.Y(n_404)
);

CKINVDCx5p33_ASAP7_75t_R g405 ( 
.A(n_361),
.Y(n_405)
);

INVx1_ASAP7_75t_SL g406 ( 
.A(n_383),
.Y(n_406)
);

CKINVDCx14_ASAP7_75t_R g407 ( 
.A(n_294),
.Y(n_407)
);

CKINVDCx20_ASAP7_75t_R g408 ( 
.A(n_91),
.Y(n_408)
);

CKINVDCx5p33_ASAP7_75t_R g409 ( 
.A(n_188),
.Y(n_409)
);

CKINVDCx5p33_ASAP7_75t_R g410 ( 
.A(n_380),
.Y(n_410)
);

INVx2_ASAP7_75t_L g411 ( 
.A(n_212),
.Y(n_411)
);

CKINVDCx20_ASAP7_75t_R g412 ( 
.A(n_323),
.Y(n_412)
);

OR2x2_ASAP7_75t_L g413 ( 
.A(n_107),
.B(n_264),
.Y(n_413)
);

INVx1_ASAP7_75t_L g414 ( 
.A(n_3),
.Y(n_414)
);

CKINVDCx5p33_ASAP7_75t_R g415 ( 
.A(n_266),
.Y(n_415)
);

CKINVDCx5p33_ASAP7_75t_R g416 ( 
.A(n_309),
.Y(n_416)
);

BUFx2_ASAP7_75t_L g417 ( 
.A(n_85),
.Y(n_417)
);

CKINVDCx5p33_ASAP7_75t_R g418 ( 
.A(n_133),
.Y(n_418)
);

CKINVDCx5p33_ASAP7_75t_R g419 ( 
.A(n_279),
.Y(n_419)
);

INVx2_ASAP7_75t_L g420 ( 
.A(n_9),
.Y(n_420)
);

INVx1_ASAP7_75t_L g421 ( 
.A(n_37),
.Y(n_421)
);

HB1xp67_ASAP7_75t_L g422 ( 
.A(n_233),
.Y(n_422)
);

NOR2xp33_ASAP7_75t_L g423 ( 
.A(n_54),
.B(n_271),
.Y(n_423)
);

CKINVDCx5p33_ASAP7_75t_R g424 ( 
.A(n_250),
.Y(n_424)
);

CKINVDCx20_ASAP7_75t_R g425 ( 
.A(n_81),
.Y(n_425)
);

CKINVDCx5p33_ASAP7_75t_R g426 ( 
.A(n_254),
.Y(n_426)
);

CKINVDCx5p33_ASAP7_75t_R g427 ( 
.A(n_204),
.Y(n_427)
);

CKINVDCx5p33_ASAP7_75t_R g428 ( 
.A(n_368),
.Y(n_428)
);

CKINVDCx5p33_ASAP7_75t_R g429 ( 
.A(n_9),
.Y(n_429)
);

BUFx6f_ASAP7_75t_L g430 ( 
.A(n_377),
.Y(n_430)
);

CKINVDCx14_ASAP7_75t_R g431 ( 
.A(n_251),
.Y(n_431)
);

CKINVDCx20_ASAP7_75t_R g432 ( 
.A(n_131),
.Y(n_432)
);

CKINVDCx5p33_ASAP7_75t_R g433 ( 
.A(n_14),
.Y(n_433)
);

CKINVDCx5p33_ASAP7_75t_R g434 ( 
.A(n_313),
.Y(n_434)
);

INVx1_ASAP7_75t_L g435 ( 
.A(n_312),
.Y(n_435)
);

CKINVDCx5p33_ASAP7_75t_R g436 ( 
.A(n_268),
.Y(n_436)
);

INVx2_ASAP7_75t_L g437 ( 
.A(n_218),
.Y(n_437)
);

CKINVDCx20_ASAP7_75t_R g438 ( 
.A(n_365),
.Y(n_438)
);

CKINVDCx16_ASAP7_75t_R g439 ( 
.A(n_80),
.Y(n_439)
);

INVx2_ASAP7_75t_L g440 ( 
.A(n_159),
.Y(n_440)
);

INVx2_ASAP7_75t_L g441 ( 
.A(n_26),
.Y(n_441)
);

INVx1_ASAP7_75t_L g442 ( 
.A(n_168),
.Y(n_442)
);

INVx1_ASAP7_75t_L g443 ( 
.A(n_111),
.Y(n_443)
);

INVx1_ASAP7_75t_L g444 ( 
.A(n_52),
.Y(n_444)
);

INVx1_ASAP7_75t_L g445 ( 
.A(n_196),
.Y(n_445)
);

INVx1_ASAP7_75t_L g446 ( 
.A(n_335),
.Y(n_446)
);

CKINVDCx16_ASAP7_75t_R g447 ( 
.A(n_151),
.Y(n_447)
);

INVx1_ASAP7_75t_L g448 ( 
.A(n_263),
.Y(n_448)
);

CKINVDCx20_ASAP7_75t_R g449 ( 
.A(n_355),
.Y(n_449)
);

CKINVDCx16_ASAP7_75t_R g450 ( 
.A(n_387),
.Y(n_450)
);

CKINVDCx5p33_ASAP7_75t_R g451 ( 
.A(n_258),
.Y(n_451)
);

CKINVDCx5p33_ASAP7_75t_R g452 ( 
.A(n_13),
.Y(n_452)
);

CKINVDCx20_ASAP7_75t_R g453 ( 
.A(n_241),
.Y(n_453)
);

CKINVDCx5p33_ASAP7_75t_R g454 ( 
.A(n_47),
.Y(n_454)
);

CKINVDCx5p33_ASAP7_75t_R g455 ( 
.A(n_5),
.Y(n_455)
);

BUFx6f_ASAP7_75t_L g456 ( 
.A(n_297),
.Y(n_456)
);

INVx1_ASAP7_75t_L g457 ( 
.A(n_224),
.Y(n_457)
);

CKINVDCx5p33_ASAP7_75t_R g458 ( 
.A(n_359),
.Y(n_458)
);

CKINVDCx20_ASAP7_75t_R g459 ( 
.A(n_177),
.Y(n_459)
);

CKINVDCx5p33_ASAP7_75t_R g460 ( 
.A(n_246),
.Y(n_460)
);

CKINVDCx16_ASAP7_75t_R g461 ( 
.A(n_60),
.Y(n_461)
);

INVx2_ASAP7_75t_L g462 ( 
.A(n_369),
.Y(n_462)
);

INVx1_ASAP7_75t_L g463 ( 
.A(n_108),
.Y(n_463)
);

CKINVDCx5p33_ASAP7_75t_R g464 ( 
.A(n_17),
.Y(n_464)
);

CKINVDCx14_ASAP7_75t_R g465 ( 
.A(n_311),
.Y(n_465)
);

HB1xp67_ASAP7_75t_L g466 ( 
.A(n_214),
.Y(n_466)
);

INVx1_ASAP7_75t_SL g467 ( 
.A(n_170),
.Y(n_467)
);

INVx1_ASAP7_75t_SL g468 ( 
.A(n_103),
.Y(n_468)
);

CKINVDCx5p33_ASAP7_75t_R g469 ( 
.A(n_38),
.Y(n_469)
);

CKINVDCx5p33_ASAP7_75t_R g470 ( 
.A(n_44),
.Y(n_470)
);

INVx1_ASAP7_75t_SL g471 ( 
.A(n_277),
.Y(n_471)
);

INVx1_ASAP7_75t_L g472 ( 
.A(n_15),
.Y(n_472)
);

AND2x2_ASAP7_75t_L g473 ( 
.A(n_216),
.B(n_78),
.Y(n_473)
);

INVx1_ASAP7_75t_SL g474 ( 
.A(n_281),
.Y(n_474)
);

INVx1_ASAP7_75t_L g475 ( 
.A(n_142),
.Y(n_475)
);

INVx1_ASAP7_75t_L g476 ( 
.A(n_371),
.Y(n_476)
);

INVx1_ASAP7_75t_L g477 ( 
.A(n_65),
.Y(n_477)
);

INVx1_ASAP7_75t_L g478 ( 
.A(n_267),
.Y(n_478)
);

CKINVDCx14_ASAP7_75t_R g479 ( 
.A(n_282),
.Y(n_479)
);

BUFx2_ASAP7_75t_L g480 ( 
.A(n_319),
.Y(n_480)
);

INVx2_ASAP7_75t_L g481 ( 
.A(n_30),
.Y(n_481)
);

BUFx10_ASAP7_75t_L g482 ( 
.A(n_3),
.Y(n_482)
);

INVx1_ASAP7_75t_L g483 ( 
.A(n_363),
.Y(n_483)
);

CKINVDCx20_ASAP7_75t_R g484 ( 
.A(n_67),
.Y(n_484)
);

INVx1_ASAP7_75t_L g485 ( 
.A(n_46),
.Y(n_485)
);

BUFx2_ASAP7_75t_L g486 ( 
.A(n_6),
.Y(n_486)
);

CKINVDCx5p33_ASAP7_75t_R g487 ( 
.A(n_114),
.Y(n_487)
);

CKINVDCx5p33_ASAP7_75t_R g488 ( 
.A(n_382),
.Y(n_488)
);

INVxp67_ASAP7_75t_L g489 ( 
.A(n_174),
.Y(n_489)
);

CKINVDCx20_ASAP7_75t_R g490 ( 
.A(n_59),
.Y(n_490)
);

INVx1_ASAP7_75t_L g491 ( 
.A(n_200),
.Y(n_491)
);

BUFx2_ASAP7_75t_SL g492 ( 
.A(n_56),
.Y(n_492)
);

INVx2_ASAP7_75t_L g493 ( 
.A(n_331),
.Y(n_493)
);

INVx1_ASAP7_75t_L g494 ( 
.A(n_12),
.Y(n_494)
);

CKINVDCx5p33_ASAP7_75t_R g495 ( 
.A(n_203),
.Y(n_495)
);

CKINVDCx5p33_ASAP7_75t_R g496 ( 
.A(n_385),
.Y(n_496)
);

CKINVDCx20_ASAP7_75t_R g497 ( 
.A(n_149),
.Y(n_497)
);

CKINVDCx20_ASAP7_75t_R g498 ( 
.A(n_249),
.Y(n_498)
);

CKINVDCx5p33_ASAP7_75t_R g499 ( 
.A(n_135),
.Y(n_499)
);

INVx1_ASAP7_75t_L g500 ( 
.A(n_217),
.Y(n_500)
);

CKINVDCx5p33_ASAP7_75t_R g501 ( 
.A(n_215),
.Y(n_501)
);

INVx2_ASAP7_75t_L g502 ( 
.A(n_283),
.Y(n_502)
);

BUFx2_ASAP7_75t_L g503 ( 
.A(n_122),
.Y(n_503)
);

BUFx6f_ASAP7_75t_L g504 ( 
.A(n_73),
.Y(n_504)
);

CKINVDCx5p33_ASAP7_75t_R g505 ( 
.A(n_53),
.Y(n_505)
);

INVx1_ASAP7_75t_L g506 ( 
.A(n_11),
.Y(n_506)
);

CKINVDCx5p33_ASAP7_75t_R g507 ( 
.A(n_97),
.Y(n_507)
);

CKINVDCx5p33_ASAP7_75t_R g508 ( 
.A(n_291),
.Y(n_508)
);

CKINVDCx20_ASAP7_75t_R g509 ( 
.A(n_364),
.Y(n_509)
);

CKINVDCx5p33_ASAP7_75t_R g510 ( 
.A(n_52),
.Y(n_510)
);

INVx2_ASAP7_75t_L g511 ( 
.A(n_302),
.Y(n_511)
);

CKINVDCx5p33_ASAP7_75t_R g512 ( 
.A(n_354),
.Y(n_512)
);

BUFx2_ASAP7_75t_L g513 ( 
.A(n_64),
.Y(n_513)
);

INVx1_ASAP7_75t_L g514 ( 
.A(n_296),
.Y(n_514)
);

INVx1_ASAP7_75t_L g515 ( 
.A(n_169),
.Y(n_515)
);

HB1xp67_ASAP7_75t_L g516 ( 
.A(n_37),
.Y(n_516)
);

CKINVDCx20_ASAP7_75t_R g517 ( 
.A(n_328),
.Y(n_517)
);

CKINVDCx5p33_ASAP7_75t_R g518 ( 
.A(n_223),
.Y(n_518)
);

INVx2_ASAP7_75t_L g519 ( 
.A(n_54),
.Y(n_519)
);

CKINVDCx20_ASAP7_75t_R g520 ( 
.A(n_17),
.Y(n_520)
);

CKINVDCx5p33_ASAP7_75t_R g521 ( 
.A(n_38),
.Y(n_521)
);

INVx2_ASAP7_75t_L g522 ( 
.A(n_240),
.Y(n_522)
);

CKINVDCx5p33_ASAP7_75t_R g523 ( 
.A(n_259),
.Y(n_523)
);

INVx1_ASAP7_75t_L g524 ( 
.A(n_98),
.Y(n_524)
);

INVx1_ASAP7_75t_L g525 ( 
.A(n_85),
.Y(n_525)
);

CKINVDCx5p33_ASAP7_75t_R g526 ( 
.A(n_278),
.Y(n_526)
);

BUFx3_ASAP7_75t_L g527 ( 
.A(n_205),
.Y(n_527)
);

CKINVDCx5p33_ASAP7_75t_R g528 ( 
.A(n_307),
.Y(n_528)
);

CKINVDCx5p33_ASAP7_75t_R g529 ( 
.A(n_71),
.Y(n_529)
);

INVx3_ASAP7_75t_L g530 ( 
.A(n_284),
.Y(n_530)
);

CKINVDCx5p33_ASAP7_75t_R g531 ( 
.A(n_25),
.Y(n_531)
);

INVx1_ASAP7_75t_L g532 ( 
.A(n_247),
.Y(n_532)
);

CKINVDCx5p33_ASAP7_75t_R g533 ( 
.A(n_156),
.Y(n_533)
);

CKINVDCx5p33_ASAP7_75t_R g534 ( 
.A(n_146),
.Y(n_534)
);

BUFx2_ASAP7_75t_L g535 ( 
.A(n_327),
.Y(n_535)
);

INVx1_ASAP7_75t_L g536 ( 
.A(n_63),
.Y(n_536)
);

INVx2_ASAP7_75t_L g537 ( 
.A(n_375),
.Y(n_537)
);

CKINVDCx5p33_ASAP7_75t_R g538 ( 
.A(n_56),
.Y(n_538)
);

CKINVDCx5p33_ASAP7_75t_R g539 ( 
.A(n_351),
.Y(n_539)
);

INVx1_ASAP7_75t_L g540 ( 
.A(n_219),
.Y(n_540)
);

BUFx6f_ASAP7_75t_L g541 ( 
.A(n_340),
.Y(n_541)
);

CKINVDCx5p33_ASAP7_75t_R g542 ( 
.A(n_164),
.Y(n_542)
);

INVx1_ASAP7_75t_L g543 ( 
.A(n_157),
.Y(n_543)
);

BUFx6f_ASAP7_75t_L g544 ( 
.A(n_207),
.Y(n_544)
);

CKINVDCx20_ASAP7_75t_R g545 ( 
.A(n_187),
.Y(n_545)
);

INVx1_ASAP7_75t_L g546 ( 
.A(n_298),
.Y(n_546)
);

CKINVDCx5p33_ASAP7_75t_R g547 ( 
.A(n_357),
.Y(n_547)
);

HB1xp67_ASAP7_75t_L g548 ( 
.A(n_202),
.Y(n_548)
);

INVx1_ASAP7_75t_L g549 ( 
.A(n_384),
.Y(n_549)
);

BUFx2_ASAP7_75t_L g550 ( 
.A(n_285),
.Y(n_550)
);

CKINVDCx20_ASAP7_75t_R g551 ( 
.A(n_57),
.Y(n_551)
);

INVx1_ASAP7_75t_L g552 ( 
.A(n_50),
.Y(n_552)
);

CKINVDCx5p33_ASAP7_75t_R g553 ( 
.A(n_325),
.Y(n_553)
);

CKINVDCx5p33_ASAP7_75t_R g554 ( 
.A(n_209),
.Y(n_554)
);

CKINVDCx5p33_ASAP7_75t_R g555 ( 
.A(n_45),
.Y(n_555)
);

CKINVDCx5p33_ASAP7_75t_R g556 ( 
.A(n_244),
.Y(n_556)
);

BUFx6f_ASAP7_75t_L g557 ( 
.A(n_239),
.Y(n_557)
);

CKINVDCx5p33_ASAP7_75t_R g558 ( 
.A(n_172),
.Y(n_558)
);

CKINVDCx5p33_ASAP7_75t_R g559 ( 
.A(n_34),
.Y(n_559)
);

INVx1_ASAP7_75t_L g560 ( 
.A(n_260),
.Y(n_560)
);

CKINVDCx16_ASAP7_75t_R g561 ( 
.A(n_178),
.Y(n_561)
);

CKINVDCx5p33_ASAP7_75t_R g562 ( 
.A(n_275),
.Y(n_562)
);

CKINVDCx5p33_ASAP7_75t_R g563 ( 
.A(n_356),
.Y(n_563)
);

CKINVDCx5p33_ASAP7_75t_R g564 ( 
.A(n_347),
.Y(n_564)
);

NOR2xp67_ASAP7_75t_L g565 ( 
.A(n_287),
.B(n_243),
.Y(n_565)
);

INVx1_ASAP7_75t_SL g566 ( 
.A(n_21),
.Y(n_566)
);

CKINVDCx5p33_ASAP7_75t_R g567 ( 
.A(n_74),
.Y(n_567)
);

INVx1_ASAP7_75t_L g568 ( 
.A(n_144),
.Y(n_568)
);

INVx1_ASAP7_75t_L g569 ( 
.A(n_206),
.Y(n_569)
);

CKINVDCx5p33_ASAP7_75t_R g570 ( 
.A(n_175),
.Y(n_570)
);

INVx1_ASAP7_75t_L g571 ( 
.A(n_306),
.Y(n_571)
);

CKINVDCx20_ASAP7_75t_R g572 ( 
.A(n_171),
.Y(n_572)
);

INVx1_ASAP7_75t_L g573 ( 
.A(n_0),
.Y(n_573)
);

CKINVDCx5p33_ASAP7_75t_R g574 ( 
.A(n_341),
.Y(n_574)
);

BUFx6f_ASAP7_75t_L g575 ( 
.A(n_138),
.Y(n_575)
);

CKINVDCx5p33_ASAP7_75t_R g576 ( 
.A(n_386),
.Y(n_576)
);

NAND2xp5_ASAP7_75t_L g577 ( 
.A(n_530),
.B(n_0),
.Y(n_577)
);

OAI22xp5_ASAP7_75t_L g578 ( 
.A1(n_393),
.A2(n_4),
.B1(n_1),
.B2(n_2),
.Y(n_578)
);

AOI22xp5_ASAP7_75t_SL g579 ( 
.A1(n_399),
.A2(n_4),
.B1(n_1),
.B2(n_2),
.Y(n_579)
);

INVx1_ASAP7_75t_L g580 ( 
.A(n_504),
.Y(n_580)
);

AND2x2_ASAP7_75t_L g581 ( 
.A(n_417),
.B(n_5),
.Y(n_581)
);

NAND2xp5_ASAP7_75t_L g582 ( 
.A(n_530),
.B(n_6),
.Y(n_582)
);

INVx2_ASAP7_75t_L g583 ( 
.A(n_504),
.Y(n_583)
);

INVx3_ASAP7_75t_L g584 ( 
.A(n_504),
.Y(n_584)
);

CKINVDCx8_ASAP7_75t_R g585 ( 
.A(n_439),
.Y(n_585)
);

INVx5_ASAP7_75t_L g586 ( 
.A(n_430),
.Y(n_586)
);

INVxp67_ASAP7_75t_L g587 ( 
.A(n_393),
.Y(n_587)
);

NOR2x1_ASAP7_75t_L g588 ( 
.A(n_527),
.B(n_127),
.Y(n_588)
);

BUFx2_ASAP7_75t_L g589 ( 
.A(n_516),
.Y(n_589)
);

AOI22xp5_ASAP7_75t_L g590 ( 
.A1(n_407),
.A2(n_10),
.B1(n_7),
.B2(n_8),
.Y(n_590)
);

AOI22xp5_ASAP7_75t_L g591 ( 
.A1(n_407),
.A2(n_10),
.B1(n_7),
.B2(n_8),
.Y(n_591)
);

INVx2_ASAP7_75t_L g592 ( 
.A(n_504),
.Y(n_592)
);

OAI21x1_ASAP7_75t_L g593 ( 
.A1(n_391),
.A2(n_462),
.B(n_411),
.Y(n_593)
);

INVx2_ASAP7_75t_L g594 ( 
.A(n_441),
.Y(n_594)
);

AND2x2_ASAP7_75t_L g595 ( 
.A(n_486),
.B(n_11),
.Y(n_595)
);

BUFx6f_ASAP7_75t_L g596 ( 
.A(n_430),
.Y(n_596)
);

BUFx6f_ASAP7_75t_L g597 ( 
.A(n_430),
.Y(n_597)
);

OA21x2_ASAP7_75t_L g598 ( 
.A1(n_441),
.A2(n_12),
.B(n_13),
.Y(n_598)
);

INVx1_ASAP7_75t_L g599 ( 
.A(n_414),
.Y(n_599)
);

INVx1_ASAP7_75t_L g600 ( 
.A(n_421),
.Y(n_600)
);

INVx1_ASAP7_75t_L g601 ( 
.A(n_443),
.Y(n_601)
);

HB1xp67_ASAP7_75t_L g602 ( 
.A(n_516),
.Y(n_602)
);

INVx1_ASAP7_75t_L g603 ( 
.A(n_444),
.Y(n_603)
);

INVx2_ASAP7_75t_L g604 ( 
.A(n_463),
.Y(n_604)
);

INVx2_ASAP7_75t_L g605 ( 
.A(n_481),
.Y(n_605)
);

INVx1_ASAP7_75t_L g606 ( 
.A(n_472),
.Y(n_606)
);

INVx5_ASAP7_75t_L g607 ( 
.A(n_456),
.Y(n_607)
);

XOR2xp5_ASAP7_75t_L g608 ( 
.A(n_461),
.B(n_14),
.Y(n_608)
);

INVx1_ASAP7_75t_L g609 ( 
.A(n_477),
.Y(n_609)
);

AND2x4_ASAP7_75t_L g610 ( 
.A(n_527),
.B(n_16),
.Y(n_610)
);

INVx1_ASAP7_75t_L g611 ( 
.A(n_485),
.Y(n_611)
);

AND2x4_ASAP7_75t_L g612 ( 
.A(n_473),
.B(n_422),
.Y(n_612)
);

BUFx6f_ASAP7_75t_L g613 ( 
.A(n_456),
.Y(n_613)
);

BUFx3_ASAP7_75t_L g614 ( 
.A(n_480),
.Y(n_614)
);

INVx3_ASAP7_75t_L g615 ( 
.A(n_420),
.Y(n_615)
);

INVx1_ASAP7_75t_L g616 ( 
.A(n_494),
.Y(n_616)
);

BUFx6f_ASAP7_75t_L g617 ( 
.A(n_456),
.Y(n_617)
);

INVx2_ASAP7_75t_L g618 ( 
.A(n_506),
.Y(n_618)
);

BUFx6f_ASAP7_75t_L g619 ( 
.A(n_456),
.Y(n_619)
);

BUFx6f_ASAP7_75t_L g620 ( 
.A(n_541),
.Y(n_620)
);

INVx2_ASAP7_75t_SL g621 ( 
.A(n_482),
.Y(n_621)
);

AND2x2_ASAP7_75t_SL g622 ( 
.A(n_447),
.B(n_16),
.Y(n_622)
);

BUFx6f_ASAP7_75t_L g623 ( 
.A(n_541),
.Y(n_623)
);

AND2x4_ASAP7_75t_L g624 ( 
.A(n_422),
.B(n_18),
.Y(n_624)
);

NAND2xp5_ASAP7_75t_L g625 ( 
.A(n_466),
.B(n_18),
.Y(n_625)
);

NAND2xp5_ASAP7_75t_L g626 ( 
.A(n_466),
.B(n_19),
.Y(n_626)
);

BUFx6f_ASAP7_75t_L g627 ( 
.A(n_541),
.Y(n_627)
);

BUFx6f_ASAP7_75t_L g628 ( 
.A(n_541),
.Y(n_628)
);

AND2x4_ASAP7_75t_L g629 ( 
.A(n_548),
.B(n_19),
.Y(n_629)
);

AND2x2_ASAP7_75t_L g630 ( 
.A(n_503),
.B(n_20),
.Y(n_630)
);

INVx2_ASAP7_75t_L g631 ( 
.A(n_524),
.Y(n_631)
);

NAND2xp5_ASAP7_75t_L g632 ( 
.A(n_548),
.B(n_400),
.Y(n_632)
);

INVx2_ASAP7_75t_L g633 ( 
.A(n_525),
.Y(n_633)
);

INVx6_ASAP7_75t_L g634 ( 
.A(n_482),
.Y(n_634)
);

HB1xp67_ASAP7_75t_L g635 ( 
.A(n_519),
.Y(n_635)
);

BUFx8_ASAP7_75t_SL g636 ( 
.A(n_513),
.Y(n_636)
);

AND2x2_ASAP7_75t_L g637 ( 
.A(n_431),
.B(n_20),
.Y(n_637)
);

AND2x2_ASAP7_75t_L g638 ( 
.A(n_431),
.B(n_21),
.Y(n_638)
);

BUFx6f_ASAP7_75t_L g639 ( 
.A(n_544),
.Y(n_639)
);

AND2x4_ASAP7_75t_L g640 ( 
.A(n_535),
.B(n_22),
.Y(n_640)
);

INVx2_ASAP7_75t_L g641 ( 
.A(n_536),
.Y(n_641)
);

BUFx8_ASAP7_75t_SL g642 ( 
.A(n_408),
.Y(n_642)
);

INVx2_ASAP7_75t_L g643 ( 
.A(n_552),
.Y(n_643)
);

OAI22x1_ASAP7_75t_R g644 ( 
.A1(n_425),
.A2(n_24),
.B1(n_22),
.B2(n_23),
.Y(n_644)
);

OAI21x1_ASAP7_75t_L g645 ( 
.A1(n_493),
.A2(n_129),
.B(n_128),
.Y(n_645)
);

NAND2xp5_ASAP7_75t_L g646 ( 
.A(n_400),
.B(n_23),
.Y(n_646)
);

NAND2xp5_ASAP7_75t_SL g647 ( 
.A(n_450),
.B(n_24),
.Y(n_647)
);

INVx1_ASAP7_75t_L g648 ( 
.A(n_573),
.Y(n_648)
);

AOI22xp5_ASAP7_75t_L g649 ( 
.A1(n_465),
.A2(n_479),
.B1(n_561),
.B2(n_433),
.Y(n_649)
);

INVx2_ASAP7_75t_L g650 ( 
.A(n_544),
.Y(n_650)
);

INVx6_ASAP7_75t_L g651 ( 
.A(n_544),
.Y(n_651)
);

INVx2_ASAP7_75t_L g652 ( 
.A(n_583),
.Y(n_652)
);

INVx1_ASAP7_75t_L g653 ( 
.A(n_592),
.Y(n_653)
);

NOR2xp33_ASAP7_75t_L g654 ( 
.A(n_632),
.B(n_550),
.Y(n_654)
);

INVx1_ASAP7_75t_L g655 ( 
.A(n_580),
.Y(n_655)
);

OR2x2_ASAP7_75t_L g656 ( 
.A(n_621),
.B(n_468),
.Y(n_656)
);

INVx1_ASAP7_75t_L g657 ( 
.A(n_583),
.Y(n_657)
);

INVx3_ASAP7_75t_L g658 ( 
.A(n_584),
.Y(n_658)
);

INVx3_ASAP7_75t_L g659 ( 
.A(n_584),
.Y(n_659)
);

INVx2_ASAP7_75t_L g660 ( 
.A(n_650),
.Y(n_660)
);

NAND2xp33_ASAP7_75t_SL g661 ( 
.A(n_625),
.B(n_626),
.Y(n_661)
);

NAND2xp33_ASAP7_75t_L g662 ( 
.A(n_637),
.B(n_413),
.Y(n_662)
);

AND2x2_ASAP7_75t_L g663 ( 
.A(n_614),
.B(n_479),
.Y(n_663)
);

AND3x2_ASAP7_75t_L g664 ( 
.A(n_638),
.B(n_423),
.C(n_404),
.Y(n_664)
);

NAND2xp5_ASAP7_75t_SL g665 ( 
.A(n_622),
.B(n_423),
.Y(n_665)
);

NAND2xp5_ASAP7_75t_SL g666 ( 
.A(n_622),
.B(n_429),
.Y(n_666)
);

INVx1_ASAP7_75t_L g667 ( 
.A(n_651),
.Y(n_667)
);

CKINVDCx5p33_ASAP7_75t_R g668 ( 
.A(n_642),
.Y(n_668)
);

INVx2_ASAP7_75t_L g669 ( 
.A(n_650),
.Y(n_669)
);

INVx4_ASAP7_75t_L g670 ( 
.A(n_586),
.Y(n_670)
);

AND3x2_ASAP7_75t_L g671 ( 
.A(n_581),
.B(n_437),
.C(n_404),
.Y(n_671)
);

NAND2xp5_ASAP7_75t_L g672 ( 
.A(n_612),
.B(n_632),
.Y(n_672)
);

NAND2xp5_ASAP7_75t_SL g673 ( 
.A(n_649),
.B(n_452),
.Y(n_673)
);

NAND2xp5_ASAP7_75t_SL g674 ( 
.A(n_647),
.B(n_454),
.Y(n_674)
);

OAI22xp5_ASAP7_75t_L g675 ( 
.A1(n_625),
.A2(n_464),
.B1(n_469),
.B2(n_455),
.Y(n_675)
);

INVx1_ASAP7_75t_L g676 ( 
.A(n_651),
.Y(n_676)
);

BUFx6f_ASAP7_75t_L g677 ( 
.A(n_596),
.Y(n_677)
);

INVx2_ASAP7_75t_L g678 ( 
.A(n_596),
.Y(n_678)
);

NAND2xp5_ASAP7_75t_SL g679 ( 
.A(n_647),
.B(n_470),
.Y(n_679)
);

AOI22xp5_ASAP7_75t_L g680 ( 
.A1(n_640),
.A2(n_630),
.B1(n_595),
.B2(n_629),
.Y(n_680)
);

NAND2xp5_ASAP7_75t_L g681 ( 
.A(n_586),
.B(n_437),
.Y(n_681)
);

INVx1_ASAP7_75t_L g682 ( 
.A(n_651),
.Y(n_682)
);

INVx3_ASAP7_75t_L g683 ( 
.A(n_596),
.Y(n_683)
);

INVx1_ASAP7_75t_L g684 ( 
.A(n_635),
.Y(n_684)
);

NAND2xp5_ASAP7_75t_SL g685 ( 
.A(n_640),
.B(n_487),
.Y(n_685)
);

INVx1_ASAP7_75t_L g686 ( 
.A(n_635),
.Y(n_686)
);

INVx1_ASAP7_75t_L g687 ( 
.A(n_599),
.Y(n_687)
);

NAND2xp5_ASAP7_75t_L g688 ( 
.A(n_607),
.B(n_440),
.Y(n_688)
);

INVx1_ASAP7_75t_L g689 ( 
.A(n_600),
.Y(n_689)
);

NAND2xp5_ASAP7_75t_SL g690 ( 
.A(n_624),
.B(n_505),
.Y(n_690)
);

NAND2xp5_ASAP7_75t_L g691 ( 
.A(n_607),
.B(n_440),
.Y(n_691)
);

INVx3_ASAP7_75t_L g692 ( 
.A(n_597),
.Y(n_692)
);

INVx2_ASAP7_75t_L g693 ( 
.A(n_597),
.Y(n_693)
);

NAND2xp5_ASAP7_75t_SL g694 ( 
.A(n_624),
.B(n_507),
.Y(n_694)
);

BUFx6f_ASAP7_75t_L g695 ( 
.A(n_597),
.Y(n_695)
);

BUFx6f_ASAP7_75t_L g696 ( 
.A(n_597),
.Y(n_696)
);

INVx8_ASAP7_75t_L g697 ( 
.A(n_607),
.Y(n_697)
);

INVx2_ASAP7_75t_L g698 ( 
.A(n_613),
.Y(n_698)
);

INVx2_ASAP7_75t_L g699 ( 
.A(n_613),
.Y(n_699)
);

NAND2xp5_ASAP7_75t_SL g700 ( 
.A(n_654),
.B(n_672),
.Y(n_700)
);

BUFx2_ASAP7_75t_L g701 ( 
.A(n_656),
.Y(n_701)
);

AOI22xp5_ASAP7_75t_L g702 ( 
.A1(n_665),
.A2(n_626),
.B1(n_590),
.B2(n_591),
.Y(n_702)
);

INVx1_ASAP7_75t_L g703 ( 
.A(n_687),
.Y(n_703)
);

NAND2xp5_ASAP7_75t_L g704 ( 
.A(n_663),
.B(n_610),
.Y(n_704)
);

INVx1_ASAP7_75t_L g705 ( 
.A(n_689),
.Y(n_705)
);

NAND2xp5_ASAP7_75t_L g706 ( 
.A(n_680),
.B(n_593),
.Y(n_706)
);

NAND2xp5_ASAP7_75t_SL g707 ( 
.A(n_661),
.B(n_585),
.Y(n_707)
);

NOR2xp33_ASAP7_75t_L g708 ( 
.A(n_673),
.B(n_674),
.Y(n_708)
);

INVx2_ASAP7_75t_L g709 ( 
.A(n_683),
.Y(n_709)
);

INVx2_ASAP7_75t_L g710 ( 
.A(n_692),
.Y(n_710)
);

NAND2xp33_ASAP7_75t_L g711 ( 
.A(n_661),
.B(n_577),
.Y(n_711)
);

NAND2xp5_ASAP7_75t_SL g712 ( 
.A(n_674),
.B(n_679),
.Y(n_712)
);

AOI22xp33_ASAP7_75t_L g713 ( 
.A1(n_662),
.A2(n_629),
.B1(n_577),
.B2(n_582),
.Y(n_713)
);

CKINVDCx20_ASAP7_75t_R g714 ( 
.A(n_668),
.Y(n_714)
);

NAND2xp5_ASAP7_75t_SL g715 ( 
.A(n_679),
.B(n_614),
.Y(n_715)
);

NOR2xp33_ASAP7_75t_L g716 ( 
.A(n_673),
.B(n_634),
.Y(n_716)
);

OR2x2_ASAP7_75t_L g717 ( 
.A(n_684),
.B(n_589),
.Y(n_717)
);

BUFx8_ASAP7_75t_L g718 ( 
.A(n_686),
.Y(n_718)
);

NAND2xp5_ASAP7_75t_SL g719 ( 
.A(n_675),
.B(n_582),
.Y(n_719)
);

AOI22xp5_ASAP7_75t_L g720 ( 
.A1(n_665),
.A2(n_578),
.B1(n_490),
.B2(n_520),
.Y(n_720)
);

NAND2xp5_ASAP7_75t_L g721 ( 
.A(n_678),
.B(n_617),
.Y(n_721)
);

NAND2xp5_ASAP7_75t_SL g722 ( 
.A(n_685),
.B(n_690),
.Y(n_722)
);

AOI22xp5_ASAP7_75t_L g723 ( 
.A1(n_662),
.A2(n_666),
.B1(n_685),
.B2(n_690),
.Y(n_723)
);

AOI22xp5_ASAP7_75t_L g724 ( 
.A1(n_666),
.A2(n_578),
.B1(n_551),
.B2(n_484),
.Y(n_724)
);

NAND3xp33_ASAP7_75t_L g725 ( 
.A(n_694),
.B(n_587),
.C(n_602),
.Y(n_725)
);

INVx1_ASAP7_75t_L g726 ( 
.A(n_658),
.Y(n_726)
);

INVx1_ASAP7_75t_L g727 ( 
.A(n_658),
.Y(n_727)
);

CKINVDCx5p33_ASAP7_75t_R g728 ( 
.A(n_694),
.Y(n_728)
);

INVxp67_ASAP7_75t_L g729 ( 
.A(n_659),
.Y(n_729)
);

INVx1_ASAP7_75t_L g730 ( 
.A(n_659),
.Y(n_730)
);

AND2x4_ASAP7_75t_L g731 ( 
.A(n_667),
.B(n_604),
.Y(n_731)
);

BUFx3_ASAP7_75t_L g732 ( 
.A(n_676),
.Y(n_732)
);

BUFx6f_ASAP7_75t_L g733 ( 
.A(n_677),
.Y(n_733)
);

BUFx6f_ASAP7_75t_L g734 ( 
.A(n_677),
.Y(n_734)
);

NAND2xp5_ASAP7_75t_SL g735 ( 
.A(n_682),
.B(n_587),
.Y(n_735)
);

AND2x4_ASAP7_75t_L g736 ( 
.A(n_671),
.B(n_618),
.Y(n_736)
);

INVxp33_ASAP7_75t_L g737 ( 
.A(n_655),
.Y(n_737)
);

INVx3_ASAP7_75t_L g738 ( 
.A(n_677),
.Y(n_738)
);

BUFx3_ASAP7_75t_L g739 ( 
.A(n_653),
.Y(n_739)
);

OAI22xp5_ASAP7_75t_SL g740 ( 
.A1(n_664),
.A2(n_608),
.B1(n_644),
.B2(n_566),
.Y(n_740)
);

AND2x4_ASAP7_75t_L g741 ( 
.A(n_657),
.B(n_631),
.Y(n_741)
);

NAND2xp5_ASAP7_75t_L g742 ( 
.A(n_693),
.B(n_698),
.Y(n_742)
);

AOI22xp33_ASAP7_75t_L g743 ( 
.A1(n_652),
.A2(n_598),
.B1(n_646),
.B2(n_602),
.Y(n_743)
);

AOI221xp5_ASAP7_75t_L g744 ( 
.A1(n_652),
.A2(n_646),
.B1(n_521),
.B2(n_531),
.C(n_529),
.Y(n_744)
);

NAND3xp33_ASAP7_75t_L g745 ( 
.A(n_681),
.B(n_648),
.C(n_603),
.Y(n_745)
);

BUFx5_ASAP7_75t_L g746 ( 
.A(n_697),
.Y(n_746)
);

BUFx4f_ASAP7_75t_L g747 ( 
.A(n_677),
.Y(n_747)
);

NOR2xp33_ASAP7_75t_L g748 ( 
.A(n_699),
.B(n_634),
.Y(n_748)
);

AND2x4_ASAP7_75t_SL g749 ( 
.A(n_660),
.B(n_403),
.Y(n_749)
);

NAND2xp33_ASAP7_75t_L g750 ( 
.A(n_688),
.B(n_544),
.Y(n_750)
);

HB1xp67_ASAP7_75t_L g751 ( 
.A(n_691),
.Y(n_751)
);

INVx1_ASAP7_75t_L g752 ( 
.A(n_669),
.Y(n_752)
);

INVx1_ASAP7_75t_L g753 ( 
.A(n_695),
.Y(n_753)
);

OR2x2_ASAP7_75t_L g754 ( 
.A(n_695),
.B(n_633),
.Y(n_754)
);

NAND2xp5_ASAP7_75t_L g755 ( 
.A(n_695),
.B(n_619),
.Y(n_755)
);

NAND2xp5_ASAP7_75t_L g756 ( 
.A(n_696),
.B(n_619),
.Y(n_756)
);

BUFx2_ASAP7_75t_L g757 ( 
.A(n_696),
.Y(n_757)
);

NOR2xp33_ASAP7_75t_L g758 ( 
.A(n_696),
.B(n_634),
.Y(n_758)
);

NAND2xp33_ASAP7_75t_L g759 ( 
.A(n_696),
.B(n_557),
.Y(n_759)
);

INVx2_ASAP7_75t_L g760 ( 
.A(n_754),
.Y(n_760)
);

OAI22xp5_ASAP7_75t_L g761 ( 
.A1(n_713),
.A2(n_432),
.B1(n_438),
.B2(n_412),
.Y(n_761)
);

OAI21xp5_ASAP7_75t_L g762 ( 
.A1(n_706),
.A2(n_645),
.B(n_588),
.Y(n_762)
);

INVx1_ASAP7_75t_L g763 ( 
.A(n_705),
.Y(n_763)
);

OAI321xp33_ASAP7_75t_L g764 ( 
.A1(n_702),
.A2(n_719),
.A3(n_708),
.B1(n_723),
.B2(n_700),
.C(n_725),
.Y(n_764)
);

INVx2_ASAP7_75t_L g765 ( 
.A(n_731),
.Y(n_765)
);

INVx2_ASAP7_75t_L g766 ( 
.A(n_731),
.Y(n_766)
);

AOI21x1_ASAP7_75t_L g767 ( 
.A1(n_742),
.A2(n_565),
.B(n_397),
.Y(n_767)
);

NAND2xp5_ASAP7_75t_L g768 ( 
.A(n_743),
.B(n_511),
.Y(n_768)
);

OAI21xp5_ASAP7_75t_L g769 ( 
.A1(n_712),
.A2(n_489),
.B(n_598),
.Y(n_769)
);

OAI321xp33_ASAP7_75t_L g770 ( 
.A1(n_702),
.A2(n_611),
.A3(n_606),
.B1(n_616),
.B2(n_609),
.C(n_601),
.Y(n_770)
);

OAI22xp5_ASAP7_75t_L g771 ( 
.A1(n_722),
.A2(n_453),
.B1(n_459),
.B2(n_449),
.Y(n_771)
);

NAND2xp5_ASAP7_75t_L g772 ( 
.A(n_751),
.B(n_729),
.Y(n_772)
);

INVx1_ASAP7_75t_L g773 ( 
.A(n_726),
.Y(n_773)
);

INVx2_ASAP7_75t_L g774 ( 
.A(n_752),
.Y(n_774)
);

BUFx6f_ASAP7_75t_L g775 ( 
.A(n_732),
.Y(n_775)
);

INVx1_ASAP7_75t_L g776 ( 
.A(n_727),
.Y(n_776)
);

INVx2_ASAP7_75t_L g777 ( 
.A(n_741),
.Y(n_777)
);

INVx2_ASAP7_75t_L g778 ( 
.A(n_741),
.Y(n_778)
);

CKINVDCx14_ASAP7_75t_R g779 ( 
.A(n_714),
.Y(n_779)
);

OAI21xp5_ASAP7_75t_L g780 ( 
.A1(n_716),
.A2(n_598),
.B(n_522),
.Y(n_780)
);

NAND2xp5_ASAP7_75t_L g781 ( 
.A(n_730),
.B(n_511),
.Y(n_781)
);

NAND2xp5_ASAP7_75t_L g782 ( 
.A(n_757),
.B(n_522),
.Y(n_782)
);

AND2x4_ASAP7_75t_L g783 ( 
.A(n_739),
.B(n_641),
.Y(n_783)
);

AOI21xp5_ASAP7_75t_L g784 ( 
.A1(n_747),
.A2(n_670),
.B(n_620),
.Y(n_784)
);

AND2x2_ASAP7_75t_L g785 ( 
.A(n_701),
.B(n_749),
.Y(n_785)
);

NAND2xp5_ASAP7_75t_L g786 ( 
.A(n_709),
.B(n_398),
.Y(n_786)
);

NOR2xp33_ASAP7_75t_L g787 ( 
.A(n_728),
.B(n_636),
.Y(n_787)
);

AOI21xp5_ASAP7_75t_L g788 ( 
.A1(n_747),
.A2(n_756),
.B(n_755),
.Y(n_788)
);

BUFx6f_ASAP7_75t_L g789 ( 
.A(n_733),
.Y(n_789)
);

OR2x2_ASAP7_75t_L g790 ( 
.A(n_717),
.B(n_492),
.Y(n_790)
);

NOR2xp67_ASAP7_75t_L g791 ( 
.A(n_745),
.B(n_132),
.Y(n_791)
);

INVx1_ASAP7_75t_SL g792 ( 
.A(n_735),
.Y(n_792)
);

AND2x2_ASAP7_75t_L g793 ( 
.A(n_737),
.B(n_643),
.Y(n_793)
);

NOR2xp33_ASAP7_75t_L g794 ( 
.A(n_707),
.B(n_636),
.Y(n_794)
);

NAND2xp5_ASAP7_75t_L g795 ( 
.A(n_753),
.B(n_435),
.Y(n_795)
);

INVx3_ASAP7_75t_L g796 ( 
.A(n_738),
.Y(n_796)
);

O2A1O1Ixp33_ASAP7_75t_L g797 ( 
.A1(n_715),
.A2(n_750),
.B(n_744),
.C(n_759),
.Y(n_797)
);

NOR2xp67_ASAP7_75t_L g798 ( 
.A(n_710),
.B(n_134),
.Y(n_798)
);

A2O1A1Ixp33_ASAP7_75t_L g799 ( 
.A1(n_720),
.A2(n_445),
.B(n_446),
.C(n_442),
.Y(n_799)
);

AOI21xp5_ASAP7_75t_L g800 ( 
.A1(n_721),
.A2(n_627),
.B(n_623),
.Y(n_800)
);

OAI22xp5_ASAP7_75t_L g801 ( 
.A1(n_720),
.A2(n_498),
.B1(n_509),
.B2(n_497),
.Y(n_801)
);

NAND2xp5_ASAP7_75t_L g802 ( 
.A(n_738),
.B(n_448),
.Y(n_802)
);

HB1xp67_ASAP7_75t_L g803 ( 
.A(n_736),
.Y(n_803)
);

NOR2xp33_ASAP7_75t_L g804 ( 
.A(n_724),
.B(n_517),
.Y(n_804)
);

A2O1A1Ixp33_ASAP7_75t_L g805 ( 
.A1(n_748),
.A2(n_475),
.B(n_476),
.C(n_457),
.Y(n_805)
);

NAND2xp5_ASAP7_75t_L g806 ( 
.A(n_734),
.B(n_478),
.Y(n_806)
);

INVx1_ASAP7_75t_L g807 ( 
.A(n_758),
.Y(n_807)
);

A2O1A1Ixp33_ASAP7_75t_L g808 ( 
.A1(n_734),
.A2(n_491),
.B(n_500),
.C(n_483),
.Y(n_808)
);

AND2x4_ASAP7_75t_L g809 ( 
.A(n_740),
.B(n_594),
.Y(n_809)
);

AOI21xp5_ASAP7_75t_L g810 ( 
.A1(n_746),
.A2(n_639),
.B(n_628),
.Y(n_810)
);

NAND2xp5_ASAP7_75t_L g811 ( 
.A(n_746),
.B(n_514),
.Y(n_811)
);

INVx2_ASAP7_75t_L g812 ( 
.A(n_718),
.Y(n_812)
);

AOI21xp5_ASAP7_75t_L g813 ( 
.A1(n_746),
.A2(n_639),
.B(n_537),
.Y(n_813)
);

AND2x2_ASAP7_75t_L g814 ( 
.A(n_718),
.B(n_615),
.Y(n_814)
);

BUFx12f_ASAP7_75t_L g815 ( 
.A(n_746),
.Y(n_815)
);

NAND2xp5_ASAP7_75t_L g816 ( 
.A(n_746),
.B(n_515),
.Y(n_816)
);

OAI22xp5_ASAP7_75t_L g817 ( 
.A1(n_713),
.A2(n_572),
.B1(n_545),
.B2(n_390),
.Y(n_817)
);

AOI21xp5_ASAP7_75t_L g818 ( 
.A1(n_704),
.A2(n_502),
.B(n_532),
.Y(n_818)
);

NOR2xp33_ASAP7_75t_L g819 ( 
.A(n_700),
.B(n_406),
.Y(n_819)
);

AOI21xp5_ASAP7_75t_L g820 ( 
.A1(n_704),
.A2(n_543),
.B(n_540),
.Y(n_820)
);

INVx3_ASAP7_75t_L g821 ( 
.A(n_731),
.Y(n_821)
);

BUFx12f_ASAP7_75t_L g822 ( 
.A(n_718),
.Y(n_822)
);

AOI21xp5_ASAP7_75t_L g823 ( 
.A1(n_704),
.A2(n_549),
.B(n_546),
.Y(n_823)
);

BUFx6f_ASAP7_75t_L g824 ( 
.A(n_732),
.Y(n_824)
);

AOI21xp5_ASAP7_75t_L g825 ( 
.A1(n_704),
.A2(n_568),
.B(n_560),
.Y(n_825)
);

AOI21xp5_ASAP7_75t_L g826 ( 
.A1(n_704),
.A2(n_571),
.B(n_569),
.Y(n_826)
);

NAND2xp5_ASAP7_75t_L g827 ( 
.A(n_713),
.B(n_467),
.Y(n_827)
);

AOI21xp5_ASAP7_75t_L g828 ( 
.A1(n_704),
.A2(n_474),
.B(n_471),
.Y(n_828)
);

INVx1_ASAP7_75t_L g829 ( 
.A(n_703),
.Y(n_829)
);

NAND3xp33_ASAP7_75t_SL g830 ( 
.A(n_723),
.B(n_538),
.C(n_510),
.Y(n_830)
);

AOI21xp5_ASAP7_75t_L g831 ( 
.A1(n_704),
.A2(n_575),
.B(n_557),
.Y(n_831)
);

NAND2xp5_ASAP7_75t_L g832 ( 
.A(n_713),
.B(n_389),
.Y(n_832)
);

INVx1_ASAP7_75t_L g833 ( 
.A(n_703),
.Y(n_833)
);

NAND3xp33_ASAP7_75t_L g834 ( 
.A(n_708),
.B(n_579),
.C(n_559),
.Y(n_834)
);

NAND2xp5_ASAP7_75t_L g835 ( 
.A(n_713),
.B(n_392),
.Y(n_835)
);

AOI21xp5_ASAP7_75t_L g836 ( 
.A1(n_704),
.A2(n_575),
.B(n_557),
.Y(n_836)
);

NAND2xp5_ASAP7_75t_L g837 ( 
.A(n_713),
.B(n_394),
.Y(n_837)
);

OR2x6_ASAP7_75t_L g838 ( 
.A(n_701),
.B(n_605),
.Y(n_838)
);

NAND2xp5_ASAP7_75t_L g839 ( 
.A(n_713),
.B(n_395),
.Y(n_839)
);

AOI21xp5_ASAP7_75t_L g840 ( 
.A1(n_704),
.A2(n_575),
.B(n_401),
.Y(n_840)
);

CKINVDCx10_ASAP7_75t_R g841 ( 
.A(n_714),
.Y(n_841)
);

AOI22xp5_ASAP7_75t_L g842 ( 
.A1(n_708),
.A2(n_402),
.B1(n_405),
.B2(n_396),
.Y(n_842)
);

NOR2xp67_ASAP7_75t_L g843 ( 
.A(n_723),
.B(n_409),
.Y(n_843)
);

NAND2xp5_ASAP7_75t_SL g844 ( 
.A(n_723),
.B(n_410),
.Y(n_844)
);

AOI22xp33_ASAP7_75t_L g845 ( 
.A1(n_711),
.A2(n_567),
.B1(n_555),
.B2(n_416),
.Y(n_845)
);

INVx1_ASAP7_75t_SL g846 ( 
.A(n_701),
.Y(n_846)
);

OAI21xp5_ASAP7_75t_L g847 ( 
.A1(n_706),
.A2(n_418),
.B(n_415),
.Y(n_847)
);

AOI21xp5_ASAP7_75t_L g848 ( 
.A1(n_704),
.A2(n_424),
.B(n_419),
.Y(n_848)
);

AOI21xp5_ASAP7_75t_L g849 ( 
.A1(n_704),
.A2(n_427),
.B(n_426),
.Y(n_849)
);

INVx1_ASAP7_75t_L g850 ( 
.A(n_703),
.Y(n_850)
);

OAI21xp5_ASAP7_75t_L g851 ( 
.A1(n_780),
.A2(n_434),
.B(n_428),
.Y(n_851)
);

NAND2xp5_ASAP7_75t_L g852 ( 
.A(n_819),
.B(n_436),
.Y(n_852)
);

NAND2xp5_ASAP7_75t_L g853 ( 
.A(n_817),
.B(n_451),
.Y(n_853)
);

OAI21xp5_ASAP7_75t_L g854 ( 
.A1(n_762),
.A2(n_769),
.B(n_768),
.Y(n_854)
);

AOI21xp5_ASAP7_75t_L g855 ( 
.A1(n_811),
.A2(n_460),
.B(n_458),
.Y(n_855)
);

AO31x2_ASAP7_75t_L g856 ( 
.A1(n_799),
.A2(n_27),
.A3(n_25),
.B(n_26),
.Y(n_856)
);

AO31x2_ASAP7_75t_L g857 ( 
.A1(n_827),
.A2(n_29),
.A3(n_27),
.B(n_28),
.Y(n_857)
);

NAND2xp5_ASAP7_75t_L g858 ( 
.A(n_807),
.B(n_488),
.Y(n_858)
);

OAI22xp5_ASAP7_75t_L g859 ( 
.A1(n_843),
.A2(n_496),
.B1(n_499),
.B2(n_495),
.Y(n_859)
);

OAI22xp5_ASAP7_75t_L g860 ( 
.A1(n_832),
.A2(n_508),
.B1(n_512),
.B2(n_501),
.Y(n_860)
);

OAI22x1_ASAP7_75t_L g861 ( 
.A1(n_804),
.A2(n_523),
.B1(n_526),
.B2(n_518),
.Y(n_861)
);

NAND2xp5_ASAP7_75t_SL g862 ( 
.A(n_764),
.B(n_528),
.Y(n_862)
);

A2O1A1Ixp33_ASAP7_75t_L g863 ( 
.A1(n_797),
.A2(n_534),
.B(n_539),
.C(n_533),
.Y(n_863)
);

OAI21xp5_ASAP7_75t_L g864 ( 
.A1(n_847),
.A2(n_547),
.B(n_542),
.Y(n_864)
);

AOI221x1_ASAP7_75t_L g865 ( 
.A1(n_830),
.A2(n_576),
.B1(n_556),
.B2(n_558),
.C(n_554),
.Y(n_865)
);

AOI21xp5_ASAP7_75t_L g866 ( 
.A1(n_816),
.A2(n_562),
.B(n_553),
.Y(n_866)
);

OAI22xp5_ASAP7_75t_L g867 ( 
.A1(n_835),
.A2(n_564),
.B1(n_570),
.B2(n_563),
.Y(n_867)
);

NAND2xp5_ASAP7_75t_SL g868 ( 
.A(n_761),
.B(n_574),
.Y(n_868)
);

NOR2xp67_ASAP7_75t_L g869 ( 
.A(n_842),
.B(n_136),
.Y(n_869)
);

AOI21xp5_ASAP7_75t_L g870 ( 
.A1(n_810),
.A2(n_139),
.B(n_137),
.Y(n_870)
);

OA21x2_ASAP7_75t_L g871 ( 
.A1(n_818),
.A2(n_143),
.B(n_141),
.Y(n_871)
);

OAI21x1_ASAP7_75t_L g872 ( 
.A1(n_796),
.A2(n_388),
.B(n_147),
.Y(n_872)
);

OAI21xp5_ASAP7_75t_L g873 ( 
.A1(n_837),
.A2(n_148),
.B(n_145),
.Y(n_873)
);

AOI21xp5_ASAP7_75t_L g874 ( 
.A1(n_844),
.A2(n_153),
.B(n_150),
.Y(n_874)
);

BUFx3_ASAP7_75t_L g875 ( 
.A(n_775),
.Y(n_875)
);

NAND2xp5_ASAP7_75t_L g876 ( 
.A(n_763),
.B(n_31),
.Y(n_876)
);

BUFx6f_ASAP7_75t_L g877 ( 
.A(n_789),
.Y(n_877)
);

OAI21xp5_ASAP7_75t_L g878 ( 
.A1(n_839),
.A2(n_155),
.B(n_154),
.Y(n_878)
);

AND2x2_ASAP7_75t_SL g879 ( 
.A(n_787),
.B(n_32),
.Y(n_879)
);

BUFx2_ASAP7_75t_L g880 ( 
.A(n_785),
.Y(n_880)
);

NOR2x1_ASAP7_75t_SL g881 ( 
.A(n_815),
.B(n_160),
.Y(n_881)
);

OAI22xp5_ASAP7_75t_L g882 ( 
.A1(n_771),
.A2(n_162),
.B1(n_163),
.B2(n_161),
.Y(n_882)
);

AOI22x1_ASAP7_75t_L g883 ( 
.A1(n_829),
.A2(n_35),
.B1(n_33),
.B2(n_34),
.Y(n_883)
);

NOR2xp33_ASAP7_75t_L g884 ( 
.A(n_801),
.B(n_772),
.Y(n_884)
);

INVx3_ASAP7_75t_SL g885 ( 
.A(n_809),
.Y(n_885)
);

OAI22xp5_ASAP7_75t_L g886 ( 
.A1(n_833),
.A2(n_166),
.B1(n_167),
.B2(n_165),
.Y(n_886)
);

AOI22xp5_ASAP7_75t_L g887 ( 
.A1(n_850),
.A2(n_176),
.B1(n_179),
.B2(n_173),
.Y(n_887)
);

OAI21xp33_ASAP7_75t_L g888 ( 
.A1(n_845),
.A2(n_36),
.B(n_39),
.Y(n_888)
);

AOI21xp33_ASAP7_75t_L g889 ( 
.A1(n_803),
.A2(n_36),
.B(n_39),
.Y(n_889)
);

A2O1A1Ixp33_ASAP7_75t_L g890 ( 
.A1(n_828),
.A2(n_42),
.B(n_40),
.C(n_41),
.Y(n_890)
);

CKINVDCx20_ASAP7_75t_R g891 ( 
.A(n_779),
.Y(n_891)
);

AOI221x1_ASAP7_75t_L g892 ( 
.A1(n_820),
.A2(n_183),
.B1(n_184),
.B2(n_182),
.C(n_180),
.Y(n_892)
);

BUFx2_ASAP7_75t_L g893 ( 
.A(n_838),
.Y(n_893)
);

NAND2xp5_ASAP7_75t_L g894 ( 
.A(n_774),
.B(n_782),
.Y(n_894)
);

AOI21xp5_ASAP7_75t_L g895 ( 
.A1(n_789),
.A2(n_186),
.B(n_185),
.Y(n_895)
);

BUFx2_ASAP7_75t_L g896 ( 
.A(n_809),
.Y(n_896)
);

BUFx2_ASAP7_75t_SL g897 ( 
.A(n_775),
.Y(n_897)
);

NAND2xp5_ASAP7_75t_L g898 ( 
.A(n_773),
.B(n_41),
.Y(n_898)
);

NAND2xp5_ASAP7_75t_L g899 ( 
.A(n_776),
.B(n_42),
.Y(n_899)
);

NAND2xp5_ASAP7_75t_L g900 ( 
.A(n_823),
.B(n_43),
.Y(n_900)
);

NAND2xp5_ASAP7_75t_L g901 ( 
.A(n_825),
.B(n_43),
.Y(n_901)
);

OAI21xp5_ASAP7_75t_L g902 ( 
.A1(n_826),
.A2(n_190),
.B(n_189),
.Y(n_902)
);

NAND2xp5_ASAP7_75t_L g903 ( 
.A(n_821),
.B(n_44),
.Y(n_903)
);

OAI21xp5_ASAP7_75t_L g904 ( 
.A1(n_840),
.A2(n_192),
.B(n_191),
.Y(n_904)
);

OAI21xp5_ASAP7_75t_L g905 ( 
.A1(n_848),
.A2(n_195),
.B(n_194),
.Y(n_905)
);

OAI21xp5_ASAP7_75t_L g906 ( 
.A1(n_849),
.A2(n_198),
.B(n_197),
.Y(n_906)
);

NAND2xp5_ASAP7_75t_L g907 ( 
.A(n_821),
.B(n_45),
.Y(n_907)
);

NAND2xp5_ASAP7_75t_L g908 ( 
.A(n_777),
.B(n_778),
.Y(n_908)
);

INVx2_ASAP7_75t_SL g909 ( 
.A(n_783),
.Y(n_909)
);

NAND2xp5_ASAP7_75t_L g910 ( 
.A(n_781),
.B(n_46),
.Y(n_910)
);

BUFx4f_ASAP7_75t_SL g911 ( 
.A(n_822),
.Y(n_911)
);

OAI21xp5_ASAP7_75t_L g912 ( 
.A1(n_802),
.A2(n_201),
.B(n_199),
.Y(n_912)
);

OR2x6_ASAP7_75t_L g913 ( 
.A(n_812),
.B(n_814),
.Y(n_913)
);

OAI21xp5_ASAP7_75t_L g914 ( 
.A1(n_795),
.A2(n_211),
.B(n_210),
.Y(n_914)
);

NOR4xp25_ASAP7_75t_L g915 ( 
.A(n_770),
.B(n_49),
.C(n_47),
.D(n_48),
.Y(n_915)
);

OAI22xp5_ASAP7_75t_L g916 ( 
.A1(n_792),
.A2(n_221),
.B1(n_222),
.B2(n_220),
.Y(n_916)
);

A2O1A1Ixp33_ASAP7_75t_L g917 ( 
.A1(n_790),
.A2(n_50),
.B(n_48),
.C(n_49),
.Y(n_917)
);

OAI22xp5_ASAP7_75t_L g918 ( 
.A1(n_765),
.A2(n_227),
.B1(n_228),
.B2(n_225),
.Y(n_918)
);

AND2x2_ASAP7_75t_L g919 ( 
.A(n_783),
.B(n_51),
.Y(n_919)
);

OAI21xp5_ASAP7_75t_L g920 ( 
.A1(n_831),
.A2(n_230),
.B(n_229),
.Y(n_920)
);

NOR2xp67_ASAP7_75t_L g921 ( 
.A(n_794),
.B(n_231),
.Y(n_921)
);

OAI21xp5_ASAP7_75t_L g922 ( 
.A1(n_836),
.A2(n_234),
.B(n_232),
.Y(n_922)
);

AOI21xp5_ASAP7_75t_L g923 ( 
.A1(n_813),
.A2(n_236),
.B(n_235),
.Y(n_923)
);

OAI21x1_ASAP7_75t_SL g924 ( 
.A1(n_767),
.A2(n_238),
.B(n_237),
.Y(n_924)
);

NAND2x1_ASAP7_75t_L g925 ( 
.A(n_824),
.B(n_766),
.Y(n_925)
);

AOI21xp5_ASAP7_75t_L g926 ( 
.A1(n_784),
.A2(n_248),
.B(n_245),
.Y(n_926)
);

AOI21xp5_ASAP7_75t_L g927 ( 
.A1(n_806),
.A2(n_253),
.B(n_252),
.Y(n_927)
);

OR2x6_ASAP7_75t_L g928 ( 
.A(n_824),
.B(n_51),
.Y(n_928)
);

AO31x2_ASAP7_75t_L g929 ( 
.A1(n_805),
.A2(n_57),
.A3(n_53),
.B(n_55),
.Y(n_929)
);

NAND2xp5_ASAP7_75t_L g930 ( 
.A(n_786),
.B(n_55),
.Y(n_930)
);

NAND2xp5_ASAP7_75t_L g931 ( 
.A(n_791),
.B(n_58),
.Y(n_931)
);

OAI21xp5_ASAP7_75t_L g932 ( 
.A1(n_791),
.A2(n_256),
.B(n_255),
.Y(n_932)
);

NAND2xp5_ASAP7_75t_L g933 ( 
.A(n_798),
.B(n_58),
.Y(n_933)
);

AND2x6_ASAP7_75t_L g934 ( 
.A(n_834),
.B(n_257),
.Y(n_934)
);

OAI21xp5_ASAP7_75t_L g935 ( 
.A1(n_800),
.A2(n_262),
.B(n_261),
.Y(n_935)
);

A2O1A1Ixp33_ASAP7_75t_L g936 ( 
.A1(n_808),
.A2(n_59),
.B(n_60),
.C(n_61),
.Y(n_936)
);

BUFx6f_ASAP7_75t_L g937 ( 
.A(n_841),
.Y(n_937)
);

NAND2x1p5_ASAP7_75t_L g938 ( 
.A(n_775),
.B(n_265),
.Y(n_938)
);

OAI22xp5_ASAP7_75t_L g939 ( 
.A1(n_827),
.A2(n_292),
.B1(n_379),
.B2(n_378),
.Y(n_939)
);

OAI21xp5_ASAP7_75t_L g940 ( 
.A1(n_780),
.A2(n_270),
.B(n_269),
.Y(n_940)
);

NAND2xp5_ASAP7_75t_L g941 ( 
.A(n_819),
.B(n_62),
.Y(n_941)
);

OAI22x1_ASAP7_75t_L g942 ( 
.A1(n_804),
.A2(n_64),
.B1(n_65),
.B2(n_66),
.Y(n_942)
);

NAND3xp33_ASAP7_75t_SL g943 ( 
.A(n_804),
.B(n_66),
.C(n_67),
.Y(n_943)
);

NAND2xp5_ASAP7_75t_L g944 ( 
.A(n_819),
.B(n_68),
.Y(n_944)
);

NAND2xp5_ASAP7_75t_L g945 ( 
.A(n_819),
.B(n_68),
.Y(n_945)
);

NAND2x1_ASAP7_75t_L g946 ( 
.A(n_789),
.B(n_272),
.Y(n_946)
);

OAI21x1_ASAP7_75t_L g947 ( 
.A1(n_788),
.A2(n_274),
.B(n_273),
.Y(n_947)
);

OAI21xp5_ASAP7_75t_L g948 ( 
.A1(n_780),
.A2(n_280),
.B(n_276),
.Y(n_948)
);

OAI22xp5_ASAP7_75t_L g949 ( 
.A1(n_827),
.A2(n_300),
.B1(n_376),
.B2(n_374),
.Y(n_949)
);

NOR2xp33_ASAP7_75t_L g950 ( 
.A(n_764),
.B(n_69),
.Y(n_950)
);

AO31x2_ASAP7_75t_L g951 ( 
.A1(n_768),
.A2(n_69),
.A3(n_70),
.B(n_71),
.Y(n_951)
);

NOR2xp33_ASAP7_75t_L g952 ( 
.A(n_764),
.B(n_70),
.Y(n_952)
);

NAND2xp5_ASAP7_75t_L g953 ( 
.A(n_819),
.B(n_72),
.Y(n_953)
);

OAI21xp5_ASAP7_75t_L g954 ( 
.A1(n_780),
.A2(n_288),
.B(n_286),
.Y(n_954)
);

NAND2xp5_ASAP7_75t_L g955 ( 
.A(n_819),
.B(n_72),
.Y(n_955)
);

NAND2xp5_ASAP7_75t_L g956 ( 
.A(n_819),
.B(n_73),
.Y(n_956)
);

OA21x2_ASAP7_75t_L g957 ( 
.A1(n_780),
.A2(n_290),
.B(n_289),
.Y(n_957)
);

NAND2xp5_ASAP7_75t_L g958 ( 
.A(n_819),
.B(n_74),
.Y(n_958)
);

AOI21xp5_ASAP7_75t_L g959 ( 
.A1(n_768),
.A2(n_295),
.B(n_293),
.Y(n_959)
);

INVx2_ASAP7_75t_L g960 ( 
.A(n_760),
.Y(n_960)
);

OAI21xp33_ASAP7_75t_L g961 ( 
.A1(n_804),
.A2(n_75),
.B(n_76),
.Y(n_961)
);

AO32x2_ASAP7_75t_L g962 ( 
.A1(n_817),
.A2(n_76),
.A3(n_77),
.B1(n_78),
.B2(n_79),
.Y(n_962)
);

OAI22xp5_ASAP7_75t_L g963 ( 
.A1(n_827),
.A2(n_308),
.B1(n_373),
.B2(n_372),
.Y(n_963)
);

AND2x2_ASAP7_75t_L g964 ( 
.A(n_793),
.B(n_77),
.Y(n_964)
);

NAND2xp5_ASAP7_75t_L g965 ( 
.A(n_819),
.B(n_80),
.Y(n_965)
);

INVx1_ASAP7_75t_L g966 ( 
.A(n_760),
.Y(n_966)
);

AOI21xp5_ASAP7_75t_L g967 ( 
.A1(n_768),
.A2(n_310),
.B(n_367),
.Y(n_967)
);

OAI21xp5_ASAP7_75t_L g968 ( 
.A1(n_780),
.A2(n_305),
.B(n_366),
.Y(n_968)
);

CKINVDCx6p67_ASAP7_75t_R g969 ( 
.A(n_841),
.Y(n_969)
);

O2A1O1Ixp5_ASAP7_75t_SL g970 ( 
.A1(n_844),
.A2(n_81),
.B(n_82),
.C(n_83),
.Y(n_970)
);

BUFx3_ASAP7_75t_L g971 ( 
.A(n_775),
.Y(n_971)
);

NAND2xp5_ASAP7_75t_L g972 ( 
.A(n_819),
.B(n_82),
.Y(n_972)
);

AO21x1_ASAP7_75t_L g973 ( 
.A1(n_780),
.A2(n_83),
.B(n_84),
.Y(n_973)
);

NAND2xp5_ASAP7_75t_L g974 ( 
.A(n_819),
.B(n_86),
.Y(n_974)
);

BUFx4f_ASAP7_75t_SL g975 ( 
.A(n_969),
.Y(n_975)
);

INVx1_ASAP7_75t_SL g976 ( 
.A(n_880),
.Y(n_976)
);

AOI22xp33_ASAP7_75t_L g977 ( 
.A1(n_950),
.A2(n_952),
.B1(n_884),
.B2(n_888),
.Y(n_977)
);

NAND2xp5_ASAP7_75t_L g978 ( 
.A(n_852),
.B(n_87),
.Y(n_978)
);

AOI221xp5_ASAP7_75t_L g979 ( 
.A1(n_915),
.A2(n_961),
.B1(n_943),
.B2(n_942),
.C(n_944),
.Y(n_979)
);

OR2x6_ASAP7_75t_L g980 ( 
.A(n_897),
.B(n_88),
.Y(n_980)
);

AND2x2_ASAP7_75t_L g981 ( 
.A(n_964),
.B(n_89),
.Y(n_981)
);

INVx2_ASAP7_75t_L g982 ( 
.A(n_960),
.Y(n_982)
);

HB1xp67_ASAP7_75t_L g983 ( 
.A(n_893),
.Y(n_983)
);

OAI21xp5_ASAP7_75t_L g984 ( 
.A1(n_854),
.A2(n_304),
.B(n_362),
.Y(n_984)
);

AOI22xp33_ASAP7_75t_L g985 ( 
.A1(n_941),
.A2(n_89),
.B1(n_90),
.B2(n_91),
.Y(n_985)
);

AOI22xp33_ASAP7_75t_SL g986 ( 
.A1(n_879),
.A2(n_90),
.B1(n_92),
.B2(n_93),
.Y(n_986)
);

AOI22xp33_ASAP7_75t_SL g987 ( 
.A1(n_945),
.A2(n_92),
.B1(n_93),
.B2(n_94),
.Y(n_987)
);

AOI22xp33_ASAP7_75t_L g988 ( 
.A1(n_953),
.A2(n_94),
.B1(n_95),
.B2(n_96),
.Y(n_988)
);

OR2x6_ASAP7_75t_L g989 ( 
.A(n_928),
.B(n_95),
.Y(n_989)
);

OA21x2_ASAP7_75t_L g990 ( 
.A1(n_940),
.A2(n_315),
.B(n_360),
.Y(n_990)
);

HB1xp67_ASAP7_75t_L g991 ( 
.A(n_896),
.Y(n_991)
);

INVx1_ASAP7_75t_L g992 ( 
.A(n_908),
.Y(n_992)
);

OAI21xp5_ASAP7_75t_L g993 ( 
.A1(n_863),
.A2(n_317),
.B(n_358),
.Y(n_993)
);

INVx1_ASAP7_75t_L g994 ( 
.A(n_894),
.Y(n_994)
);

CKINVDCx5p33_ASAP7_75t_R g995 ( 
.A(n_891),
.Y(n_995)
);

OAI22xp5_ASAP7_75t_L g996 ( 
.A1(n_853),
.A2(n_956),
.B1(n_958),
.B2(n_955),
.Y(n_996)
);

AOI22xp33_ASAP7_75t_L g997 ( 
.A1(n_965),
.A2(n_99),
.B1(n_100),
.B2(n_101),
.Y(n_997)
);

OAI21xp5_ASAP7_75t_L g998 ( 
.A1(n_948),
.A2(n_314),
.B(n_353),
.Y(n_998)
);

OAI21x1_ASAP7_75t_L g999 ( 
.A1(n_947),
.A2(n_303),
.B(n_352),
.Y(n_999)
);

NAND2xp5_ASAP7_75t_L g1000 ( 
.A(n_972),
.B(n_100),
.Y(n_1000)
);

AOI22xp33_ASAP7_75t_L g1001 ( 
.A1(n_974),
.A2(n_101),
.B1(n_102),
.B2(n_103),
.Y(n_1001)
);

AOI22xp33_ASAP7_75t_L g1002 ( 
.A1(n_862),
.A2(n_102),
.B1(n_104),
.B2(n_105),
.Y(n_1002)
);

NOR2xp33_ASAP7_75t_L g1003 ( 
.A(n_858),
.B(n_104),
.Y(n_1003)
);

AND2x6_ASAP7_75t_SL g1004 ( 
.A(n_913),
.B(n_105),
.Y(n_1004)
);

AOI21x1_ASAP7_75t_L g1005 ( 
.A1(n_954),
.A2(n_318),
.B(n_350),
.Y(n_1005)
);

OAI21xp5_ASAP7_75t_L g1006 ( 
.A1(n_968),
.A2(n_320),
.B(n_349),
.Y(n_1006)
);

A2O1A1Ixp33_ASAP7_75t_L g1007 ( 
.A1(n_873),
.A2(n_878),
.B(n_864),
.C(n_851),
.Y(n_1007)
);

AND2x2_ASAP7_75t_L g1008 ( 
.A(n_966),
.B(n_106),
.Y(n_1008)
);

NAND2x1_ASAP7_75t_L g1009 ( 
.A(n_877),
.B(n_299),
.Y(n_1009)
);

AOI21xp33_ASAP7_75t_L g1010 ( 
.A1(n_868),
.A2(n_106),
.B(n_107),
.Y(n_1010)
);

OAI21xp5_ASAP7_75t_L g1011 ( 
.A1(n_970),
.A2(n_321),
.B(n_348),
.Y(n_1011)
);

OAI22xp5_ASAP7_75t_L g1012 ( 
.A1(n_869),
.A2(n_370),
.B1(n_346),
.B2(n_345),
.Y(n_1012)
);

NAND2xp5_ASAP7_75t_SL g1013 ( 
.A(n_909),
.B(n_344),
.Y(n_1013)
);

AOI21xp5_ASAP7_75t_L g1014 ( 
.A1(n_905),
.A2(n_343),
.B(n_342),
.Y(n_1014)
);

OAI22xp5_ASAP7_75t_L g1015 ( 
.A1(n_903),
.A2(n_338),
.B1(n_337),
.B2(n_336),
.Y(n_1015)
);

AND2x4_ASAP7_75t_L g1016 ( 
.A(n_919),
.B(n_334),
.Y(n_1016)
);

OAI22xp5_ASAP7_75t_L g1017 ( 
.A1(n_907),
.A2(n_333),
.B1(n_332),
.B2(n_330),
.Y(n_1017)
);

INVx2_ASAP7_75t_L g1018 ( 
.A(n_925),
.Y(n_1018)
);

AOI21xp33_ASAP7_75t_L g1019 ( 
.A1(n_860),
.A2(n_109),
.B(n_110),
.Y(n_1019)
);

INVx1_ASAP7_75t_L g1020 ( 
.A(n_910),
.Y(n_1020)
);

INVx2_ASAP7_75t_L g1021 ( 
.A(n_876),
.Y(n_1021)
);

OA21x2_ASAP7_75t_L g1022 ( 
.A1(n_912),
.A2(n_326),
.B(n_324),
.Y(n_1022)
);

AND2x2_ASAP7_75t_L g1023 ( 
.A(n_885),
.B(n_112),
.Y(n_1023)
);

OAI22xp5_ASAP7_75t_L g1024 ( 
.A1(n_932),
.A2(n_931),
.B1(n_921),
.B2(n_933),
.Y(n_1024)
);

AOI22x1_ASAP7_75t_L g1025 ( 
.A1(n_861),
.A2(n_322),
.B1(n_114),
.B2(n_115),
.Y(n_1025)
);

NOR2xp33_ASAP7_75t_L g1026 ( 
.A(n_898),
.B(n_113),
.Y(n_1026)
);

CKINVDCx11_ASAP7_75t_R g1027 ( 
.A(n_937),
.Y(n_1027)
);

AOI21xp5_ASAP7_75t_L g1028 ( 
.A1(n_906),
.A2(n_126),
.B(n_115),
.Y(n_1028)
);

INVx1_ASAP7_75t_L g1029 ( 
.A(n_899),
.Y(n_1029)
);

AOI21xp5_ASAP7_75t_L g1030 ( 
.A1(n_904),
.A2(n_113),
.B(n_116),
.Y(n_1030)
);

CKINVDCx11_ASAP7_75t_R g1031 ( 
.A(n_937),
.Y(n_1031)
);

OAI21x1_ASAP7_75t_SL g1032 ( 
.A1(n_881),
.A2(n_116),
.B(n_117),
.Y(n_1032)
);

BUFx6f_ASAP7_75t_L g1033 ( 
.A(n_946),
.Y(n_1033)
);

CKINVDCx20_ASAP7_75t_R g1034 ( 
.A(n_911),
.Y(n_1034)
);

BUFx12f_ASAP7_75t_L g1035 ( 
.A(n_913),
.Y(n_1035)
);

AO31x2_ASAP7_75t_L g1036 ( 
.A1(n_892),
.A2(n_117),
.A3(n_118),
.B(n_119),
.Y(n_1036)
);

OAI21x1_ASAP7_75t_L g1037 ( 
.A1(n_872),
.A2(n_118),
.B(n_119),
.Y(n_1037)
);

HB1xp67_ASAP7_75t_L g1038 ( 
.A(n_928),
.Y(n_1038)
);

AO21x2_ASAP7_75t_L g1039 ( 
.A1(n_914),
.A2(n_126),
.B(n_120),
.Y(n_1039)
);

OAI22xp5_ASAP7_75t_L g1040 ( 
.A1(n_902),
.A2(n_121),
.B1(n_122),
.B2(n_123),
.Y(n_1040)
);

AOI21xp5_ASAP7_75t_L g1041 ( 
.A1(n_957),
.A2(n_124),
.B(n_125),
.Y(n_1041)
);

CKINVDCx16_ASAP7_75t_R g1042 ( 
.A(n_934),
.Y(n_1042)
);

AOI22xp5_ASAP7_75t_L g1043 ( 
.A1(n_867),
.A2(n_859),
.B1(n_934),
.B2(n_882),
.Y(n_1043)
);

INVx4_ASAP7_75t_L g1044 ( 
.A(n_938),
.Y(n_1044)
);

INVx1_ASAP7_75t_L g1045 ( 
.A(n_930),
.Y(n_1045)
);

INVx2_ASAP7_75t_SL g1046 ( 
.A(n_857),
.Y(n_1046)
);

INVx4_ASAP7_75t_L g1047 ( 
.A(n_934),
.Y(n_1047)
);

AOI22xp33_ASAP7_75t_L g1048 ( 
.A1(n_900),
.A2(n_901),
.B1(n_883),
.B2(n_889),
.Y(n_1048)
);

OAI22xp5_ASAP7_75t_L g1049 ( 
.A1(n_957),
.A2(n_887),
.B1(n_917),
.B2(n_890),
.Y(n_1049)
);

INVx1_ASAP7_75t_L g1050 ( 
.A(n_951),
.Y(n_1050)
);

AO21x2_ASAP7_75t_L g1051 ( 
.A1(n_924),
.A2(n_935),
.B(n_922),
.Y(n_1051)
);

AO31x2_ASAP7_75t_L g1052 ( 
.A1(n_865),
.A2(n_936),
.A3(n_939),
.B(n_963),
.Y(n_1052)
);

AND2x2_ASAP7_75t_L g1053 ( 
.A(n_962),
.B(n_881),
.Y(n_1053)
);

AND2x2_ASAP7_75t_L g1054 ( 
.A(n_962),
.B(n_857),
.Y(n_1054)
);

NAND2xp5_ASAP7_75t_L g1055 ( 
.A(n_855),
.B(n_866),
.Y(n_1055)
);

AO32x2_ASAP7_75t_L g1056 ( 
.A1(n_962),
.A2(n_949),
.A3(n_916),
.B1(n_886),
.B2(n_918),
.Y(n_1056)
);

OAI22xp5_ASAP7_75t_L g1057 ( 
.A1(n_920),
.A2(n_874),
.B1(n_967),
.B2(n_959),
.Y(n_1057)
);

NOR2xp67_ASAP7_75t_L g1058 ( 
.A(n_895),
.B(n_927),
.Y(n_1058)
);

HB1xp67_ASAP7_75t_L g1059 ( 
.A(n_856),
.Y(n_1059)
);

OAI22xp5_ASAP7_75t_L g1060 ( 
.A1(n_871),
.A2(n_926),
.B1(n_870),
.B2(n_923),
.Y(n_1060)
);

INVx2_ASAP7_75t_R g1061 ( 
.A(n_929),
.Y(n_1061)
);

INVxp67_ASAP7_75t_SL g1062 ( 
.A(n_929),
.Y(n_1062)
);

INVx1_ASAP7_75t_L g1063 ( 
.A(n_857),
.Y(n_1063)
);

BUFx2_ASAP7_75t_L g1064 ( 
.A(n_896),
.Y(n_1064)
);

AO31x2_ASAP7_75t_L g1065 ( 
.A1(n_973),
.A2(n_952),
.A3(n_950),
.B(n_863),
.Y(n_1065)
);

AO21x2_ASAP7_75t_L g1066 ( 
.A1(n_854),
.A2(n_948),
.B(n_940),
.Y(n_1066)
);

AOI22xp33_ASAP7_75t_L g1067 ( 
.A1(n_950),
.A2(n_952),
.B1(n_708),
.B2(n_884),
.Y(n_1067)
);

AND2x4_ASAP7_75t_L g1068 ( 
.A(n_875),
.B(n_971),
.Y(n_1068)
);

OR2x2_ASAP7_75t_L g1069 ( 
.A(n_884),
.B(n_846),
.Y(n_1069)
);

CKINVDCx16_ASAP7_75t_R g1070 ( 
.A(n_891),
.Y(n_1070)
);

AOI21xp5_ASAP7_75t_L g1071 ( 
.A1(n_854),
.A2(n_948),
.B(n_940),
.Y(n_1071)
);

AND2x2_ASAP7_75t_L g1072 ( 
.A(n_884),
.B(n_701),
.Y(n_1072)
);

NAND2xp5_ASAP7_75t_L g1073 ( 
.A(n_884),
.B(n_819),
.Y(n_1073)
);

CKINVDCx5p33_ASAP7_75t_R g1074 ( 
.A(n_969),
.Y(n_1074)
);

NOR2xp33_ASAP7_75t_SL g1075 ( 
.A(n_969),
.B(n_937),
.Y(n_1075)
);

AOI22x1_ASAP7_75t_L g1076 ( 
.A1(n_940),
.A2(n_948),
.B1(n_968),
.B2(n_954),
.Y(n_1076)
);

INVx4_ASAP7_75t_L g1077 ( 
.A(n_877),
.Y(n_1077)
);

INVx4_ASAP7_75t_L g1078 ( 
.A(n_877),
.Y(n_1078)
);

CKINVDCx20_ASAP7_75t_R g1079 ( 
.A(n_891),
.Y(n_1079)
);

OR2x2_ASAP7_75t_L g1080 ( 
.A(n_1069),
.B(n_1072),
.Y(n_1080)
);

CKINVDCx5p33_ASAP7_75t_R g1081 ( 
.A(n_1027),
.Y(n_1081)
);

NAND2xp5_ASAP7_75t_L g1082 ( 
.A(n_1073),
.B(n_994),
.Y(n_1082)
);

AOI221xp5_ASAP7_75t_L g1083 ( 
.A1(n_1067),
.A2(n_977),
.B1(n_1040),
.B2(n_979),
.C(n_1019),
.Y(n_1083)
);

BUFx3_ASAP7_75t_L g1084 ( 
.A(n_1068),
.Y(n_1084)
);

AND2x2_ASAP7_75t_L g1085 ( 
.A(n_1021),
.B(n_981),
.Y(n_1085)
);

NAND2xp5_ASAP7_75t_L g1086 ( 
.A(n_992),
.B(n_1020),
.Y(n_1086)
);

AO21x1_ASAP7_75t_SL g1087 ( 
.A1(n_998),
.A2(n_1006),
.B(n_984),
.Y(n_1087)
);

CKINVDCx11_ASAP7_75t_R g1088 ( 
.A(n_1031),
.Y(n_1088)
);

INVx2_ASAP7_75t_L g1089 ( 
.A(n_982),
.Y(n_1089)
);

NAND2xp5_ASAP7_75t_L g1090 ( 
.A(n_992),
.B(n_1020),
.Y(n_1090)
);

CKINVDCx5p33_ASAP7_75t_R g1091 ( 
.A(n_1074),
.Y(n_1091)
);

INVxp33_ASAP7_75t_L g1092 ( 
.A(n_991),
.Y(n_1092)
);

HB1xp67_ASAP7_75t_L g1093 ( 
.A(n_983),
.Y(n_1093)
);

AOI21x1_ASAP7_75t_L g1094 ( 
.A1(n_1024),
.A2(n_1060),
.B(n_1057),
.Y(n_1094)
);

BUFx2_ASAP7_75t_L g1095 ( 
.A(n_1064),
.Y(n_1095)
);

INVx3_ASAP7_75t_L g1096 ( 
.A(n_1033),
.Y(n_1096)
);

AOI22xp33_ASAP7_75t_L g1097 ( 
.A1(n_1076),
.A2(n_986),
.B1(n_985),
.B2(n_988),
.Y(n_1097)
);

INVxp67_ASAP7_75t_L g1098 ( 
.A(n_976),
.Y(n_1098)
);

NAND2xp5_ASAP7_75t_L g1099 ( 
.A(n_1045),
.B(n_1029),
.Y(n_1099)
);

AOI22xp33_ASAP7_75t_L g1100 ( 
.A1(n_997),
.A2(n_1001),
.B1(n_1025),
.B2(n_1003),
.Y(n_1100)
);

BUFx2_ASAP7_75t_L g1101 ( 
.A(n_1038),
.Y(n_1101)
);

AND2x2_ASAP7_75t_L g1102 ( 
.A(n_1008),
.B(n_1016),
.Y(n_1102)
);

INVx1_ASAP7_75t_L g1103 ( 
.A(n_1059),
.Y(n_1103)
);

AOI22x1_ASAP7_75t_L g1104 ( 
.A1(n_1071),
.A2(n_1028),
.B1(n_1030),
.B2(n_1014),
.Y(n_1104)
);

AOI22xp33_ASAP7_75t_L g1105 ( 
.A1(n_1026),
.A2(n_1002),
.B1(n_1010),
.B2(n_987),
.Y(n_1105)
);

BUFx2_ASAP7_75t_R g1106 ( 
.A(n_995),
.Y(n_1106)
);

NAND3x1_ASAP7_75t_L g1107 ( 
.A(n_1023),
.B(n_1000),
.C(n_978),
.Y(n_1107)
);

INVx2_ASAP7_75t_L g1108 ( 
.A(n_1046),
.Y(n_1108)
);

INVx2_ASAP7_75t_L g1109 ( 
.A(n_1018),
.Y(n_1109)
);

OAI22xp5_ASAP7_75t_SL g1110 ( 
.A1(n_989),
.A2(n_980),
.B1(n_1042),
.B2(n_1079),
.Y(n_1110)
);

INVx3_ASAP7_75t_L g1111 ( 
.A(n_1033),
.Y(n_1111)
);

AOI21xp33_ASAP7_75t_L g1112 ( 
.A1(n_996),
.A2(n_1007),
.B(n_1048),
.Y(n_1112)
);

INVx1_ASAP7_75t_L g1113 ( 
.A(n_1063),
.Y(n_1113)
);

INVx1_ASAP7_75t_L g1114 ( 
.A(n_1063),
.Y(n_1114)
);

INVx1_ASAP7_75t_L g1115 ( 
.A(n_1050),
.Y(n_1115)
);

NAND2xp5_ASAP7_75t_L g1116 ( 
.A(n_1066),
.B(n_1065),
.Y(n_1116)
);

BUFx2_ASAP7_75t_L g1117 ( 
.A(n_1035),
.Y(n_1117)
);

OR2x2_ASAP7_75t_L g1118 ( 
.A(n_1070),
.B(n_1044),
.Y(n_1118)
);

NAND2xp5_ASAP7_75t_L g1119 ( 
.A(n_1066),
.B(n_1065),
.Y(n_1119)
);

HB1xp67_ASAP7_75t_L g1120 ( 
.A(n_1077),
.Y(n_1120)
);

OR2x2_ASAP7_75t_L g1121 ( 
.A(n_1078),
.B(n_1047),
.Y(n_1121)
);

HB1xp67_ASAP7_75t_L g1122 ( 
.A(n_1062),
.Y(n_1122)
);

CKINVDCx5p33_ASAP7_75t_R g1123 ( 
.A(n_975),
.Y(n_1123)
);

CKINVDCx11_ASAP7_75t_R g1124 ( 
.A(n_1034),
.Y(n_1124)
);

OAI22xp5_ASAP7_75t_L g1125 ( 
.A1(n_1043),
.A2(n_1049),
.B1(n_1047),
.B2(n_1053),
.Y(n_1125)
);

CKINVDCx20_ASAP7_75t_R g1126 ( 
.A(n_1075),
.Y(n_1126)
);

INVx2_ASAP7_75t_SL g1127 ( 
.A(n_1009),
.Y(n_1127)
);

INVx1_ASAP7_75t_L g1128 ( 
.A(n_1013),
.Y(n_1128)
);

OR2x6_ASAP7_75t_L g1129 ( 
.A(n_1012),
.B(n_993),
.Y(n_1129)
);

BUFx3_ASAP7_75t_L g1130 ( 
.A(n_1032),
.Y(n_1130)
);

NAND2xp5_ASAP7_75t_L g1131 ( 
.A(n_1054),
.B(n_1039),
.Y(n_1131)
);

HB1xp67_ASAP7_75t_SL g1132 ( 
.A(n_1015),
.Y(n_1132)
);

NOR2xp33_ASAP7_75t_L g1133 ( 
.A(n_1005),
.B(n_1004),
.Y(n_1133)
);

AO21x2_ASAP7_75t_L g1134 ( 
.A1(n_1051),
.A2(n_1041),
.B(n_1058),
.Y(n_1134)
);

OR2x2_ASAP7_75t_L g1135 ( 
.A(n_1052),
.B(n_1061),
.Y(n_1135)
);

AND2x2_ASAP7_75t_L g1136 ( 
.A(n_1052),
.B(n_1011),
.Y(n_1136)
);

HB1xp67_ASAP7_75t_L g1137 ( 
.A(n_1052),
.Y(n_1137)
);

HB1xp67_ASAP7_75t_L g1138 ( 
.A(n_1036),
.Y(n_1138)
);

AOI22xp33_ASAP7_75t_L g1139 ( 
.A1(n_990),
.A2(n_1022),
.B1(n_1017),
.B2(n_1037),
.Y(n_1139)
);

AND2x2_ASAP7_75t_L g1140 ( 
.A(n_1056),
.B(n_1022),
.Y(n_1140)
);

NAND2xp5_ASAP7_75t_L g1141 ( 
.A(n_990),
.B(n_1055),
.Y(n_1141)
);

INVx2_ASAP7_75t_L g1142 ( 
.A(n_999),
.Y(n_1142)
);

AND2x2_ASAP7_75t_L g1143 ( 
.A(n_1085),
.B(n_1102),
.Y(n_1143)
);

HB1xp67_ASAP7_75t_L g1144 ( 
.A(n_1122),
.Y(n_1144)
);

OR2x2_ASAP7_75t_L g1145 ( 
.A(n_1080),
.B(n_1099),
.Y(n_1145)
);

INVx1_ASAP7_75t_SL g1146 ( 
.A(n_1095),
.Y(n_1146)
);

BUFx2_ASAP7_75t_L g1147 ( 
.A(n_1098),
.Y(n_1147)
);

BUFx2_ASAP7_75t_L g1148 ( 
.A(n_1098),
.Y(n_1148)
);

OR2x2_ASAP7_75t_L g1149 ( 
.A(n_1099),
.B(n_1082),
.Y(n_1149)
);

OR2x2_ASAP7_75t_L g1150 ( 
.A(n_1082),
.B(n_1093),
.Y(n_1150)
);

BUFx6f_ASAP7_75t_L g1151 ( 
.A(n_1084),
.Y(n_1151)
);

NAND2xp5_ASAP7_75t_L g1152 ( 
.A(n_1086),
.B(n_1090),
.Y(n_1152)
);

INVx2_ASAP7_75t_SL g1153 ( 
.A(n_1118),
.Y(n_1153)
);

BUFx3_ASAP7_75t_L g1154 ( 
.A(n_1101),
.Y(n_1154)
);

NOR2x1_ASAP7_75t_SL g1155 ( 
.A(n_1129),
.B(n_1087),
.Y(n_1155)
);

INVxp67_ASAP7_75t_L g1156 ( 
.A(n_1093),
.Y(n_1156)
);

BUFx3_ASAP7_75t_L g1157 ( 
.A(n_1117),
.Y(n_1157)
);

AND2x2_ASAP7_75t_L g1158 ( 
.A(n_1092),
.B(n_1133),
.Y(n_1158)
);

AND2x2_ASAP7_75t_L g1159 ( 
.A(n_1133),
.B(n_1089),
.Y(n_1159)
);

INVx3_ASAP7_75t_SL g1160 ( 
.A(n_1081),
.Y(n_1160)
);

INVx1_ASAP7_75t_L g1161 ( 
.A(n_1113),
.Y(n_1161)
);

HB1xp67_ASAP7_75t_L g1162 ( 
.A(n_1103),
.Y(n_1162)
);

INVx1_ASAP7_75t_L g1163 ( 
.A(n_1114),
.Y(n_1163)
);

AOI22xp33_ASAP7_75t_L g1164 ( 
.A1(n_1083),
.A2(n_1105),
.B1(n_1097),
.B2(n_1100),
.Y(n_1164)
);

INVx1_ASAP7_75t_L g1165 ( 
.A(n_1115),
.Y(n_1165)
);

AND2x2_ASAP7_75t_L g1166 ( 
.A(n_1086),
.B(n_1090),
.Y(n_1166)
);

BUFx6f_ASAP7_75t_L g1167 ( 
.A(n_1121),
.Y(n_1167)
);

OR2x2_ASAP7_75t_L g1168 ( 
.A(n_1110),
.B(n_1131),
.Y(n_1168)
);

NAND2xp5_ASAP7_75t_L g1169 ( 
.A(n_1083),
.B(n_1097),
.Y(n_1169)
);

AO22x1_ASAP7_75t_L g1170 ( 
.A1(n_1128),
.A2(n_1111),
.B1(n_1096),
.B2(n_1091),
.Y(n_1170)
);

NAND2xp5_ASAP7_75t_L g1171 ( 
.A(n_1112),
.B(n_1125),
.Y(n_1171)
);

AND2x2_ASAP7_75t_L g1172 ( 
.A(n_1106),
.B(n_1120),
.Y(n_1172)
);

NAND2xp5_ASAP7_75t_L g1173 ( 
.A(n_1112),
.B(n_1125),
.Y(n_1173)
);

OR2x2_ASAP7_75t_L g1174 ( 
.A(n_1109),
.B(n_1116),
.Y(n_1174)
);

AND2x2_ASAP7_75t_L g1175 ( 
.A(n_1106),
.B(n_1100),
.Y(n_1175)
);

NAND2xp5_ASAP7_75t_L g1176 ( 
.A(n_1129),
.B(n_1136),
.Y(n_1176)
);

INVxp67_ASAP7_75t_SL g1177 ( 
.A(n_1108),
.Y(n_1177)
);

OR2x2_ASAP7_75t_L g1178 ( 
.A(n_1116),
.B(n_1119),
.Y(n_1178)
);

BUFx2_ASAP7_75t_L g1179 ( 
.A(n_1126),
.Y(n_1179)
);

INVx3_ASAP7_75t_L g1180 ( 
.A(n_1130),
.Y(n_1180)
);

AOI22xp5_ASAP7_75t_L g1181 ( 
.A1(n_1107),
.A2(n_1132),
.B1(n_1126),
.B2(n_1127),
.Y(n_1181)
);

BUFx6f_ASAP7_75t_L g1182 ( 
.A(n_1130),
.Y(n_1182)
);

AND2x2_ASAP7_75t_L g1183 ( 
.A(n_1124),
.B(n_1123),
.Y(n_1183)
);

BUFx6f_ASAP7_75t_SL g1184 ( 
.A(n_1088),
.Y(n_1184)
);

HB1xp67_ASAP7_75t_L g1185 ( 
.A(n_1150),
.Y(n_1185)
);

NAND2xp5_ASAP7_75t_L g1186 ( 
.A(n_1149),
.B(n_1119),
.Y(n_1186)
);

INVxp33_ASAP7_75t_L g1187 ( 
.A(n_1143),
.Y(n_1187)
);

HB1xp67_ASAP7_75t_L g1188 ( 
.A(n_1156),
.Y(n_1188)
);

NAND2xp5_ASAP7_75t_L g1189 ( 
.A(n_1166),
.B(n_1137),
.Y(n_1189)
);

NAND2xp5_ASAP7_75t_L g1190 ( 
.A(n_1145),
.B(n_1140),
.Y(n_1190)
);

INVx1_ASAP7_75t_L g1191 ( 
.A(n_1162),
.Y(n_1191)
);

HB1xp67_ASAP7_75t_L g1192 ( 
.A(n_1156),
.Y(n_1192)
);

OAI22xp5_ASAP7_75t_L g1193 ( 
.A1(n_1164),
.A2(n_1132),
.B1(n_1104),
.B2(n_1139),
.Y(n_1193)
);

INVx2_ASAP7_75t_SL g1194 ( 
.A(n_1182),
.Y(n_1194)
);

INVxp67_ASAP7_75t_L g1195 ( 
.A(n_1147),
.Y(n_1195)
);

INVx1_ASAP7_75t_L g1196 ( 
.A(n_1161),
.Y(n_1196)
);

INVx1_ASAP7_75t_L g1197 ( 
.A(n_1163),
.Y(n_1197)
);

BUFx2_ASAP7_75t_SL g1198 ( 
.A(n_1184),
.Y(n_1198)
);

INVx1_ASAP7_75t_L g1199 ( 
.A(n_1165),
.Y(n_1199)
);

BUFx2_ASAP7_75t_L g1200 ( 
.A(n_1154),
.Y(n_1200)
);

NOR2x1_ASAP7_75t_L g1201 ( 
.A(n_1180),
.B(n_1141),
.Y(n_1201)
);

AND2x2_ASAP7_75t_L g1202 ( 
.A(n_1176),
.B(n_1138),
.Y(n_1202)
);

INVxp67_ASAP7_75t_SL g1203 ( 
.A(n_1177),
.Y(n_1203)
);

OR2x2_ASAP7_75t_L g1204 ( 
.A(n_1178),
.B(n_1135),
.Y(n_1204)
);

INVx1_ASAP7_75t_L g1205 ( 
.A(n_1144),
.Y(n_1205)
);

CKINVDCx20_ASAP7_75t_R g1206 ( 
.A(n_1160),
.Y(n_1206)
);

OR2x2_ASAP7_75t_L g1207 ( 
.A(n_1168),
.B(n_1158),
.Y(n_1207)
);

BUFx12f_ASAP7_75t_L g1208 ( 
.A(n_1179),
.Y(n_1208)
);

AND2x2_ASAP7_75t_L g1209 ( 
.A(n_1171),
.B(n_1094),
.Y(n_1209)
);

NAND2xp5_ASAP7_75t_L g1210 ( 
.A(n_1152),
.B(n_1124),
.Y(n_1210)
);

AND2x2_ASAP7_75t_L g1211 ( 
.A(n_1173),
.B(n_1134),
.Y(n_1211)
);

BUFx2_ASAP7_75t_SL g1212 ( 
.A(n_1184),
.Y(n_1212)
);

BUFx2_ASAP7_75t_L g1213 ( 
.A(n_1154),
.Y(n_1213)
);

INVx2_ASAP7_75t_SL g1214 ( 
.A(n_1182),
.Y(n_1214)
);

NAND2xp5_ASAP7_75t_L g1215 ( 
.A(n_1159),
.B(n_1142),
.Y(n_1215)
);

BUFx3_ASAP7_75t_L g1216 ( 
.A(n_1148),
.Y(n_1216)
);

NAND2xp5_ASAP7_75t_L g1217 ( 
.A(n_1185),
.B(n_1164),
.Y(n_1217)
);

NAND2xp5_ASAP7_75t_L g1218 ( 
.A(n_1188),
.B(n_1169),
.Y(n_1218)
);

INVxp67_ASAP7_75t_L g1219 ( 
.A(n_1216),
.Y(n_1219)
);

NAND2xp5_ASAP7_75t_L g1220 ( 
.A(n_1192),
.B(n_1169),
.Y(n_1220)
);

NAND2xp5_ASAP7_75t_L g1221 ( 
.A(n_1186),
.B(n_1203),
.Y(n_1221)
);

INVx1_ASAP7_75t_L g1222 ( 
.A(n_1196),
.Y(n_1222)
);

OR2x2_ASAP7_75t_L g1223 ( 
.A(n_1204),
.B(n_1174),
.Y(n_1223)
);

AND2x2_ASAP7_75t_L g1224 ( 
.A(n_1202),
.B(n_1155),
.Y(n_1224)
);

INVx1_ASAP7_75t_L g1225 ( 
.A(n_1197),
.Y(n_1225)
);

INVx1_ASAP7_75t_L g1226 ( 
.A(n_1199),
.Y(n_1226)
);

NAND2x1p5_ASAP7_75t_L g1227 ( 
.A(n_1201),
.B(n_1180),
.Y(n_1227)
);

NAND2xp5_ASAP7_75t_L g1228 ( 
.A(n_1190),
.B(n_1167),
.Y(n_1228)
);

NAND2xp5_ASAP7_75t_L g1229 ( 
.A(n_1189),
.B(n_1191),
.Y(n_1229)
);

NOR2xp67_ASAP7_75t_L g1230 ( 
.A(n_1195),
.B(n_1153),
.Y(n_1230)
);

HB1xp67_ASAP7_75t_L g1231 ( 
.A(n_1205),
.Y(n_1231)
);

NAND2xp5_ASAP7_75t_L g1232 ( 
.A(n_1221),
.B(n_1211),
.Y(n_1232)
);

NAND2xp5_ASAP7_75t_L g1233 ( 
.A(n_1228),
.B(n_1207),
.Y(n_1233)
);

INVx1_ASAP7_75t_L g1234 ( 
.A(n_1222),
.Y(n_1234)
);

NAND2xp5_ASAP7_75t_SL g1235 ( 
.A(n_1217),
.B(n_1193),
.Y(n_1235)
);

INVx1_ASAP7_75t_L g1236 ( 
.A(n_1225),
.Y(n_1236)
);

OAI21xp33_ASAP7_75t_L g1237 ( 
.A1(n_1218),
.A2(n_1181),
.B(n_1175),
.Y(n_1237)
);

INVx1_ASAP7_75t_L g1238 ( 
.A(n_1225),
.Y(n_1238)
);

NOR3xp33_ASAP7_75t_L g1239 ( 
.A(n_1220),
.B(n_1170),
.C(n_1210),
.Y(n_1239)
);

CKINVDCx14_ASAP7_75t_R g1240 ( 
.A(n_1224),
.Y(n_1240)
);

INVx1_ASAP7_75t_L g1241 ( 
.A(n_1226),
.Y(n_1241)
);

INVx1_ASAP7_75t_L g1242 ( 
.A(n_1226),
.Y(n_1242)
);

INVx1_ASAP7_75t_L g1243 ( 
.A(n_1231),
.Y(n_1243)
);

AOI21xp33_ASAP7_75t_L g1244 ( 
.A1(n_1235),
.A2(n_1187),
.B(n_1215),
.Y(n_1244)
);

AOI22xp5_ASAP7_75t_L g1245 ( 
.A1(n_1235),
.A2(n_1239),
.B1(n_1237),
.B2(n_1209),
.Y(n_1245)
);

OAI21xp5_ASAP7_75t_L g1246 ( 
.A1(n_1243),
.A2(n_1230),
.B(n_1227),
.Y(n_1246)
);

INVx1_ASAP7_75t_L g1247 ( 
.A(n_1234),
.Y(n_1247)
);

AOI21xp33_ASAP7_75t_L g1248 ( 
.A1(n_1232),
.A2(n_1187),
.B(n_1223),
.Y(n_1248)
);

INVx1_ASAP7_75t_L g1249 ( 
.A(n_1236),
.Y(n_1249)
);

INVx1_ASAP7_75t_L g1250 ( 
.A(n_1238),
.Y(n_1250)
);

INVx1_ASAP7_75t_L g1251 ( 
.A(n_1241),
.Y(n_1251)
);

INVxp67_ASAP7_75t_L g1252 ( 
.A(n_1233),
.Y(n_1252)
);

INVx1_ASAP7_75t_L g1253 ( 
.A(n_1242),
.Y(n_1253)
);

OAI21xp5_ASAP7_75t_SL g1254 ( 
.A1(n_1240),
.A2(n_1224),
.B(n_1172),
.Y(n_1254)
);

INVx1_ASAP7_75t_L g1255 ( 
.A(n_1247),
.Y(n_1255)
);

INVxp67_ASAP7_75t_L g1256 ( 
.A(n_1249),
.Y(n_1256)
);

AOI221xp5_ASAP7_75t_L g1257 ( 
.A1(n_1245),
.A2(n_1219),
.B1(n_1146),
.B2(n_1216),
.C(n_1213),
.Y(n_1257)
);

INVx1_ASAP7_75t_L g1258 ( 
.A(n_1250),
.Y(n_1258)
);

NAND3xp33_ASAP7_75t_SL g1259 ( 
.A(n_1246),
.B(n_1206),
.C(n_1200),
.Y(n_1259)
);

INVx1_ASAP7_75t_L g1260 ( 
.A(n_1251),
.Y(n_1260)
);

INVx1_ASAP7_75t_L g1261 ( 
.A(n_1253),
.Y(n_1261)
);

AOI22xp5_ASAP7_75t_L g1262 ( 
.A1(n_1259),
.A2(n_1254),
.B1(n_1252),
.B2(n_1246),
.Y(n_1262)
);

OAI21xp5_ASAP7_75t_SL g1263 ( 
.A1(n_1259),
.A2(n_1244),
.B(n_1248),
.Y(n_1263)
);

NAND2xp33_ASAP7_75t_SL g1264 ( 
.A(n_1257),
.B(n_1206),
.Y(n_1264)
);

AOI21xp5_ASAP7_75t_L g1265 ( 
.A1(n_1256),
.A2(n_1244),
.B(n_1229),
.Y(n_1265)
);

INVx1_ASAP7_75t_L g1266 ( 
.A(n_1265),
.Y(n_1266)
);

AND2x2_ASAP7_75t_L g1267 ( 
.A(n_1262),
.B(n_1240),
.Y(n_1267)
);

AND2x4_ASAP7_75t_L g1268 ( 
.A(n_1264),
.B(n_1255),
.Y(n_1268)
);

NOR4xp25_ASAP7_75t_L g1269 ( 
.A(n_1263),
.B(n_1261),
.C(n_1260),
.D(n_1258),
.Y(n_1269)
);

NOR3xp33_ASAP7_75t_L g1270 ( 
.A(n_1266),
.B(n_1088),
.C(n_1183),
.Y(n_1270)
);

NAND3xp33_ASAP7_75t_L g1271 ( 
.A(n_1269),
.B(n_1182),
.C(n_1167),
.Y(n_1271)
);

AND2x4_ASAP7_75t_L g1272 ( 
.A(n_1270),
.B(n_1267),
.Y(n_1272)
);

XOR2xp5_ASAP7_75t_L g1273 ( 
.A(n_1272),
.B(n_1198),
.Y(n_1273)
);

INVx2_ASAP7_75t_L g1274 ( 
.A(n_1273),
.Y(n_1274)
);

NAND3xp33_ASAP7_75t_L g1275 ( 
.A(n_1274),
.B(n_1271),
.C(n_1268),
.Y(n_1275)
);

AOI22xp5_ASAP7_75t_L g1276 ( 
.A1(n_1275),
.A2(n_1212),
.B1(n_1208),
.B2(n_1160),
.Y(n_1276)
);

INVx2_ASAP7_75t_L g1277 ( 
.A(n_1276),
.Y(n_1277)
);

OAI21x1_ASAP7_75t_SL g1278 ( 
.A1(n_1277),
.A2(n_1157),
.B(n_1194),
.Y(n_1278)
);

NAND2xp5_ASAP7_75t_SL g1279 ( 
.A(n_1278),
.B(n_1151),
.Y(n_1279)
);

INVx1_ASAP7_75t_L g1280 ( 
.A(n_1279),
.Y(n_1280)
);

AOI22xp33_ASAP7_75t_L g1281 ( 
.A1(n_1280),
.A2(n_1151),
.B1(n_1214),
.B2(n_1194),
.Y(n_1281)
);


endmodule