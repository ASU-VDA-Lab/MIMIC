module fake_ariane_2318_n_667 (n_83, n_8, n_56, n_60, n_64, n_119, n_124, n_90, n_38, n_47, n_110, n_18, n_86, n_75, n_89, n_67, n_34, n_69, n_95, n_92, n_143, n_98, n_74, n_113, n_114, n_33, n_19, n_40, n_120, n_106, n_12, n_53, n_111, n_21, n_115, n_133, n_66, n_71, n_24, n_7, n_109, n_96, n_49, n_20, n_100, n_17, n_50, n_132, n_62, n_51, n_76, n_103, n_79, n_26, n_3, n_46, n_0, n_84, n_36, n_91, n_107, n_72, n_105, n_128, n_44, n_30, n_82, n_31, n_42, n_57, n_131, n_70, n_10, n_117, n_139, n_85, n_130, n_144, n_6, n_48, n_94, n_101, n_4, n_134, n_2, n_32, n_37, n_58, n_65, n_123, n_9, n_138, n_112, n_45, n_11, n_129, n_126, n_137, n_122, n_52, n_135, n_73, n_77, n_15, n_118, n_93, n_121, n_23, n_61, n_108, n_102, n_125, n_22, n_43, n_1, n_81, n_87, n_13, n_27, n_29, n_41, n_140, n_55, n_136, n_28, n_80, n_97, n_142, n_14, n_88, n_141, n_68, n_116, n_104, n_78, n_39, n_59, n_63, n_99, n_16, n_5, n_127, n_35, n_54, n_25, n_667);

input n_83;
input n_8;
input n_56;
input n_60;
input n_64;
input n_119;
input n_124;
input n_90;
input n_38;
input n_47;
input n_110;
input n_18;
input n_86;
input n_75;
input n_89;
input n_67;
input n_34;
input n_69;
input n_95;
input n_92;
input n_143;
input n_98;
input n_74;
input n_113;
input n_114;
input n_33;
input n_19;
input n_40;
input n_120;
input n_106;
input n_12;
input n_53;
input n_111;
input n_21;
input n_115;
input n_133;
input n_66;
input n_71;
input n_24;
input n_7;
input n_109;
input n_96;
input n_49;
input n_20;
input n_100;
input n_17;
input n_50;
input n_132;
input n_62;
input n_51;
input n_76;
input n_103;
input n_79;
input n_26;
input n_3;
input n_46;
input n_0;
input n_84;
input n_36;
input n_91;
input n_107;
input n_72;
input n_105;
input n_128;
input n_44;
input n_30;
input n_82;
input n_31;
input n_42;
input n_57;
input n_131;
input n_70;
input n_10;
input n_117;
input n_139;
input n_85;
input n_130;
input n_144;
input n_6;
input n_48;
input n_94;
input n_101;
input n_4;
input n_134;
input n_2;
input n_32;
input n_37;
input n_58;
input n_65;
input n_123;
input n_9;
input n_138;
input n_112;
input n_45;
input n_11;
input n_129;
input n_126;
input n_137;
input n_122;
input n_52;
input n_135;
input n_73;
input n_77;
input n_15;
input n_118;
input n_93;
input n_121;
input n_23;
input n_61;
input n_108;
input n_102;
input n_125;
input n_22;
input n_43;
input n_1;
input n_81;
input n_87;
input n_13;
input n_27;
input n_29;
input n_41;
input n_140;
input n_55;
input n_136;
input n_28;
input n_80;
input n_97;
input n_142;
input n_14;
input n_88;
input n_141;
input n_68;
input n_116;
input n_104;
input n_78;
input n_39;
input n_59;
input n_63;
input n_99;
input n_16;
input n_5;
input n_127;
input n_35;
input n_54;
input n_25;

output n_667;

wire n_295;
wire n_356;
wire n_556;
wire n_170;
wire n_190;
wire n_160;
wire n_180;
wire n_386;
wire n_307;
wire n_516;
wire n_589;
wire n_332;
wire n_581;
wire n_294;
wire n_646;
wire n_197;
wire n_640;
wire n_463;
wire n_176;
wire n_404;
wire n_172;
wire n_651;
wire n_347;
wire n_423;
wire n_183;
wire n_469;
wire n_479;
wire n_603;
wire n_373;
wire n_299;
wire n_541;
wire n_499;
wire n_564;
wire n_610;
wire n_205;
wire n_341;
wire n_421;
wire n_245;
wire n_549;
wire n_522;
wire n_319;
wire n_591;
wire n_416;
wire n_283;
wire n_525;
wire n_187;
wire n_367;
wire n_649;
wire n_598;
wire n_345;
wire n_374;
wire n_318;
wire n_244;
wire n_643;
wire n_226;
wire n_220;
wire n_261;
wire n_663;
wire n_370;
wire n_189;
wire n_286;
wire n_443;
wire n_586;
wire n_605;
wire n_424;
wire n_528;
wire n_584;
wire n_387;
wire n_406;
wire n_524;
wire n_391;
wire n_349;
wire n_634;
wire n_466;
wire n_346;
wire n_214;
wire n_348;
wire n_552;
wire n_462;
wire n_607;
wire n_410;
wire n_379;
wire n_445;
wire n_515;
wire n_162;
wire n_264;
wire n_198;
wire n_232;
wire n_441;
wire n_568;
wire n_385;
wire n_637;
wire n_327;
wire n_372;
wire n_377;
wire n_396;
wire n_631;
wire n_399;
wire n_554;
wire n_520;
wire n_279;
wire n_207;
wire n_363;
wire n_354;
wire n_419;
wire n_151;
wire n_146;
wire n_230;
wire n_270;
wire n_194;
wire n_633;
wire n_154;
wire n_338;
wire n_285;
wire n_473;
wire n_186;
wire n_202;
wire n_145;
wire n_193;
wire n_500;
wire n_665;
wire n_336;
wire n_315;
wire n_594;
wire n_311;
wire n_239;
wire n_402;
wire n_272;
wire n_339;
wire n_487;
wire n_167;
wire n_422;
wire n_153;
wire n_648;
wire n_269;
wire n_597;
wire n_158;
wire n_259;
wire n_446;
wire n_553;
wire n_566;
wire n_578;
wire n_625;
wire n_152;
wire n_405;
wire n_557;
wire n_169;
wire n_173;
wire n_242;
wire n_645;
wire n_309;
wire n_320;
wire n_331;
wire n_559;
wire n_401;
wire n_485;
wire n_267;
wire n_495;
wire n_504;
wire n_647;
wire n_483;
wire n_335;
wire n_435;
wire n_350;
wire n_291;
wire n_381;
wire n_344;
wire n_426;
wire n_481;
wire n_433;
wire n_600;
wire n_398;
wire n_210;
wire n_200;
wire n_529;
wire n_502;
wire n_166;
wire n_253;
wire n_561;
wire n_218;
wire n_271;
wire n_465;
wire n_507;
wire n_486;
wire n_247;
wire n_569;
wire n_567;
wire n_369;
wire n_240;
wire n_224;
wire n_547;
wire n_420;
wire n_562;
wire n_518;
wire n_439;
wire n_604;
wire n_614;
wire n_222;
wire n_478;
wire n_510;
wire n_256;
wire n_326;
wire n_227;
wire n_188;
wire n_323;
wire n_550;
wire n_635;
wire n_330;
wire n_400;
wire n_282;
wire n_328;
wire n_368;
wire n_590;
wire n_277;
wire n_248;
wire n_301;
wire n_467;
wire n_432;
wire n_545;
wire n_536;
wire n_644;
wire n_293;
wire n_620;
wire n_228;
wire n_325;
wire n_276;
wire n_636;
wire n_427;
wire n_587;
wire n_497;
wire n_303;
wire n_442;
wire n_168;
wire n_206;
wire n_352;
wire n_538;
wire n_576;
wire n_511;
wire n_611;
wire n_238;
wire n_365;
wire n_429;
wire n_455;
wire n_654;
wire n_588;
wire n_638;
wire n_334;
wire n_192;
wire n_661;
wire n_488;
wire n_300;
wire n_533;
wire n_505;
wire n_163;
wire n_390;
wire n_498;
wire n_501;
wire n_438;
wire n_314;
wire n_440;
wire n_627;
wire n_273;
wire n_305;
wire n_539;
wire n_312;
wire n_233;
wire n_388;
wire n_333;
wire n_449;
wire n_612;
wire n_413;
wire n_392;
wire n_376;
wire n_512;
wire n_579;
wire n_459;
wire n_221;
wire n_321;
wire n_361;
wire n_458;
wire n_149;
wire n_383;
wire n_623;
wire n_237;
wire n_175;
wire n_453;
wire n_491;
wire n_181;
wire n_616;
wire n_617;
wire n_658;
wire n_630;
wire n_570;
wire n_260;
wire n_362;
wire n_543;
wire n_310;
wire n_236;
wire n_601;
wire n_565;
wire n_281;
wire n_628;
wire n_461;
wire n_209;
wire n_262;
wire n_490;
wire n_225;
wire n_235;
wire n_660;
wire n_464;
wire n_575;
wire n_546;
wire n_297;
wire n_662;
wire n_641;
wire n_503;
wire n_290;
wire n_527;
wire n_371;
wire n_199;
wire n_639;
wire n_217;
wire n_452;
wire n_178;
wire n_551;
wire n_308;
wire n_417;
wire n_201;
wire n_572;
wire n_343;
wire n_414;
wire n_571;
wire n_287;
wire n_302;
wire n_380;
wire n_582;
wire n_284;
wire n_448;
wire n_593;
wire n_249;
wire n_534;
wire n_212;
wire n_355;
wire n_444;
wire n_609;
wire n_278;
wire n_255;
wire n_560;
wire n_450;
wire n_257;
wire n_148;
wire n_652;
wire n_451;
wire n_613;
wire n_475;
wire n_409;
wire n_171;
wire n_519;
wire n_384;
wire n_468;
wire n_526;
wire n_182;
wire n_482;
wire n_316;
wire n_196;
wire n_577;
wire n_407;
wire n_254;
wire n_596;
wire n_476;
wire n_460;
wire n_219;
wire n_535;
wire n_231;
wire n_366;
wire n_656;
wire n_555;
wire n_234;
wire n_492;
wire n_574;
wire n_280;
wire n_215;
wire n_252;
wire n_629;
wire n_664;
wire n_161;
wire n_454;
wire n_298;
wire n_532;
wire n_415;
wire n_655;
wire n_544;
wire n_216;
wire n_540;
wire n_599;
wire n_514;
wire n_418;
wire n_537;
wire n_223;
wire n_403;
wire n_389;
wire n_657;
wire n_513;
wire n_288;
wire n_179;
wire n_395;
wire n_621;
wire n_195;
wire n_606;
wire n_213;
wire n_304;
wire n_659;
wire n_509;
wire n_583;
wire n_306;
wire n_666;
wire n_313;
wire n_430;
wire n_626;
wire n_493;
wire n_203;
wire n_378;
wire n_436;
wire n_150;
wire n_375;
wire n_324;
wire n_585;
wire n_619;
wire n_437;
wire n_337;
wire n_274;
wire n_622;
wire n_472;
wire n_296;
wire n_265;
wire n_208;
wire n_456;
wire n_156;
wire n_292;
wire n_174;
wire n_275;
wire n_147;
wire n_204;
wire n_615;
wire n_521;
wire n_496;
wire n_342;
wire n_246;
wire n_517;
wire n_530;
wire n_428;
wire n_159;
wire n_358;
wire n_580;
wire n_608;
wire n_494;
wire n_263;
wire n_434;
wire n_360;
wire n_563;
wire n_229;
wire n_394;
wire n_250;
wire n_165;
wire n_317;
wire n_243;
wire n_329;
wire n_185;
wire n_340;
wire n_289;
wire n_548;
wire n_542;
wire n_523;
wire n_268;
wire n_266;
wire n_470;
wire n_457;
wire n_164;
wire n_157;
wire n_632;
wire n_184;
wire n_177;
wire n_477;
wire n_364;
wire n_258;
wire n_650;
wire n_425;
wire n_431;
wire n_508;
wire n_624;
wire n_618;
wire n_411;
wire n_484;
wire n_353;
wire n_241;
wire n_357;
wire n_412;
wire n_447;
wire n_191;
wire n_382;
wire n_489;
wire n_480;
wire n_211;
wire n_642;
wire n_408;
wire n_595;
wire n_322;
wire n_251;
wire n_506;
wire n_602;
wire n_558;
wire n_592;
wire n_397;
wire n_471;
wire n_351;
wire n_393;
wire n_474;
wire n_653;
wire n_359;
wire n_155;
wire n_573;
wire n_531;

CKINVDCx5p33_ASAP7_75t_R g145 ( 
.A(n_89),
.Y(n_145)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_23),
.Y(n_146)
);

CKINVDCx5p33_ASAP7_75t_R g147 ( 
.A(n_135),
.Y(n_147)
);

CKINVDCx5p33_ASAP7_75t_R g148 ( 
.A(n_143),
.Y(n_148)
);

CKINVDCx5p33_ASAP7_75t_R g149 ( 
.A(n_118),
.Y(n_149)
);

CKINVDCx5p33_ASAP7_75t_R g150 ( 
.A(n_133),
.Y(n_150)
);

CKINVDCx5p33_ASAP7_75t_R g151 ( 
.A(n_125),
.Y(n_151)
);

CKINVDCx5p33_ASAP7_75t_R g152 ( 
.A(n_108),
.Y(n_152)
);

INVx2_ASAP7_75t_L g153 ( 
.A(n_124),
.Y(n_153)
);

CKINVDCx5p33_ASAP7_75t_R g154 ( 
.A(n_37),
.Y(n_154)
);

INVx2_ASAP7_75t_L g155 ( 
.A(n_111),
.Y(n_155)
);

CKINVDCx5p33_ASAP7_75t_R g156 ( 
.A(n_44),
.Y(n_156)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_7),
.Y(n_157)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_105),
.Y(n_158)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_47),
.Y(n_159)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_1),
.Y(n_160)
);

CKINVDCx5p33_ASAP7_75t_R g161 ( 
.A(n_96),
.Y(n_161)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_119),
.Y(n_162)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_103),
.Y(n_163)
);

CKINVDCx5p33_ASAP7_75t_R g164 ( 
.A(n_60),
.Y(n_164)
);

CKINVDCx5p33_ASAP7_75t_R g165 ( 
.A(n_142),
.Y(n_165)
);

BUFx10_ASAP7_75t_L g166 ( 
.A(n_10),
.Y(n_166)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_38),
.Y(n_167)
);

CKINVDCx5p33_ASAP7_75t_R g168 ( 
.A(n_97),
.Y(n_168)
);

INVx2_ASAP7_75t_L g169 ( 
.A(n_112),
.Y(n_169)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_64),
.Y(n_170)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_59),
.Y(n_171)
);

CKINVDCx14_ASAP7_75t_R g172 ( 
.A(n_12),
.Y(n_172)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_6),
.Y(n_173)
);

HB1xp67_ASAP7_75t_L g174 ( 
.A(n_98),
.Y(n_174)
);

CKINVDCx5p33_ASAP7_75t_R g175 ( 
.A(n_93),
.Y(n_175)
);

INVx3_ASAP7_75t_L g176 ( 
.A(n_80),
.Y(n_176)
);

BUFx3_ASAP7_75t_L g177 ( 
.A(n_123),
.Y(n_177)
);

CKINVDCx20_ASAP7_75t_R g178 ( 
.A(n_71),
.Y(n_178)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_65),
.Y(n_179)
);

CKINVDCx20_ASAP7_75t_R g180 ( 
.A(n_100),
.Y(n_180)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_33),
.Y(n_181)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_95),
.Y(n_182)
);

CKINVDCx5p33_ASAP7_75t_R g183 ( 
.A(n_68),
.Y(n_183)
);

CKINVDCx5p33_ASAP7_75t_R g184 ( 
.A(n_82),
.Y(n_184)
);

CKINVDCx20_ASAP7_75t_R g185 ( 
.A(n_45),
.Y(n_185)
);

CKINVDCx5p33_ASAP7_75t_R g186 ( 
.A(n_85),
.Y(n_186)
);

CKINVDCx5p33_ASAP7_75t_R g187 ( 
.A(n_12),
.Y(n_187)
);

INVx3_ASAP7_75t_L g188 ( 
.A(n_101),
.Y(n_188)
);

CKINVDCx5p33_ASAP7_75t_R g189 ( 
.A(n_73),
.Y(n_189)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_28),
.Y(n_190)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_16),
.Y(n_191)
);

CKINVDCx5p33_ASAP7_75t_R g192 ( 
.A(n_137),
.Y(n_192)
);

CKINVDCx5p33_ASAP7_75t_R g193 ( 
.A(n_131),
.Y(n_193)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_127),
.Y(n_194)
);

CKINVDCx5p33_ASAP7_75t_R g195 ( 
.A(n_78),
.Y(n_195)
);

CKINVDCx5p33_ASAP7_75t_R g196 ( 
.A(n_63),
.Y(n_196)
);

CKINVDCx20_ASAP7_75t_R g197 ( 
.A(n_121),
.Y(n_197)
);

CKINVDCx5p33_ASAP7_75t_R g198 ( 
.A(n_53),
.Y(n_198)
);

BUFx6f_ASAP7_75t_L g199 ( 
.A(n_41),
.Y(n_199)
);

INVx2_ASAP7_75t_SL g200 ( 
.A(n_34),
.Y(n_200)
);

CKINVDCx5p33_ASAP7_75t_R g201 ( 
.A(n_104),
.Y(n_201)
);

CKINVDCx5p33_ASAP7_75t_R g202 ( 
.A(n_0),
.Y(n_202)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_77),
.Y(n_203)
);

CKINVDCx5p33_ASAP7_75t_R g204 ( 
.A(n_66),
.Y(n_204)
);

CKINVDCx5p33_ASAP7_75t_R g205 ( 
.A(n_107),
.Y(n_205)
);

CKINVDCx5p33_ASAP7_75t_R g206 ( 
.A(n_52),
.Y(n_206)
);

CKINVDCx5p33_ASAP7_75t_R g207 ( 
.A(n_144),
.Y(n_207)
);

CKINVDCx5p33_ASAP7_75t_R g208 ( 
.A(n_14),
.Y(n_208)
);

CKINVDCx5p33_ASAP7_75t_R g209 ( 
.A(n_99),
.Y(n_209)
);

CKINVDCx5p33_ASAP7_75t_R g210 ( 
.A(n_102),
.Y(n_210)
);

CKINVDCx5p33_ASAP7_75t_R g211 ( 
.A(n_54),
.Y(n_211)
);

CKINVDCx5p33_ASAP7_75t_R g212 ( 
.A(n_56),
.Y(n_212)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_14),
.Y(n_213)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_157),
.Y(n_214)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_160),
.Y(n_215)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_173),
.Y(n_216)
);

XNOR2xp5_ASAP7_75t_L g217 ( 
.A(n_178),
.B(n_0),
.Y(n_217)
);

CKINVDCx5p33_ASAP7_75t_R g218 ( 
.A(n_180),
.Y(n_218)
);

HB1xp67_ASAP7_75t_L g219 ( 
.A(n_172),
.Y(n_219)
);

NOR2xp67_ASAP7_75t_L g220 ( 
.A(n_176),
.B(n_1),
.Y(n_220)
);

INVxp67_ASAP7_75t_SL g221 ( 
.A(n_191),
.Y(n_221)
);

CKINVDCx20_ASAP7_75t_R g222 ( 
.A(n_172),
.Y(n_222)
);

CKINVDCx5p33_ASAP7_75t_R g223 ( 
.A(n_185),
.Y(n_223)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_213),
.Y(n_224)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_174),
.Y(n_225)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_166),
.Y(n_226)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_166),
.Y(n_227)
);

INVxp67_ASAP7_75t_SL g228 ( 
.A(n_176),
.Y(n_228)
);

BUFx6f_ASAP7_75t_SL g229 ( 
.A(n_166),
.Y(n_229)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_146),
.Y(n_230)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_158),
.Y(n_231)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_159),
.Y(n_232)
);

CKINVDCx5p33_ASAP7_75t_R g233 ( 
.A(n_197),
.Y(n_233)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_162),
.Y(n_234)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_163),
.Y(n_235)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_167),
.Y(n_236)
);

CKINVDCx5p33_ASAP7_75t_R g237 ( 
.A(n_187),
.Y(n_237)
);

CKINVDCx5p33_ASAP7_75t_R g238 ( 
.A(n_202),
.Y(n_238)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_170),
.Y(n_239)
);

HB1xp67_ASAP7_75t_L g240 ( 
.A(n_208),
.Y(n_240)
);

CKINVDCx16_ASAP7_75t_R g241 ( 
.A(n_178),
.Y(n_241)
);

INVxp67_ASAP7_75t_SL g242 ( 
.A(n_176),
.Y(n_242)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_171),
.Y(n_243)
);

BUFx3_ASAP7_75t_L g244 ( 
.A(n_177),
.Y(n_244)
);

CKINVDCx20_ASAP7_75t_R g245 ( 
.A(n_177),
.Y(n_245)
);

CKINVDCx5p33_ASAP7_75t_R g246 ( 
.A(n_145),
.Y(n_246)
);

BUFx5_ASAP7_75t_L g247 ( 
.A(n_179),
.Y(n_247)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_181),
.Y(n_248)
);

CKINVDCx5p33_ASAP7_75t_R g249 ( 
.A(n_147),
.Y(n_249)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_182),
.Y(n_250)
);

CKINVDCx20_ASAP7_75t_R g251 ( 
.A(n_148),
.Y(n_251)
);

CKINVDCx5p33_ASAP7_75t_R g252 ( 
.A(n_149),
.Y(n_252)
);

CKINVDCx20_ASAP7_75t_R g253 ( 
.A(n_212),
.Y(n_253)
);

CKINVDCx16_ASAP7_75t_R g254 ( 
.A(n_199),
.Y(n_254)
);

CKINVDCx20_ASAP7_75t_R g255 ( 
.A(n_150),
.Y(n_255)
);

INVx1_ASAP7_75t_SL g256 ( 
.A(n_151),
.Y(n_256)
);

CKINVDCx20_ASAP7_75t_R g257 ( 
.A(n_152),
.Y(n_257)
);

CKINVDCx5p33_ASAP7_75t_R g258 ( 
.A(n_154),
.Y(n_258)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_190),
.Y(n_259)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_194),
.Y(n_260)
);

NOR2xp33_ASAP7_75t_R g261 ( 
.A(n_246),
.B(n_156),
.Y(n_261)
);

HB1xp67_ASAP7_75t_L g262 ( 
.A(n_219),
.Y(n_262)
);

AND2x6_ASAP7_75t_L g263 ( 
.A(n_244),
.B(n_188),
.Y(n_263)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_214),
.Y(n_264)
);

BUFx2_ASAP7_75t_L g265 ( 
.A(n_237),
.Y(n_265)
);

AND2x4_ASAP7_75t_L g266 ( 
.A(n_219),
.B(n_188),
.Y(n_266)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_215),
.Y(n_267)
);

INVx3_ASAP7_75t_L g268 ( 
.A(n_244),
.Y(n_268)
);

BUFx6f_ASAP7_75t_L g269 ( 
.A(n_230),
.Y(n_269)
);

INVx2_ASAP7_75t_L g270 ( 
.A(n_247),
.Y(n_270)
);

OAI22xp5_ASAP7_75t_SL g271 ( 
.A1(n_217),
.A2(n_153),
.B1(n_155),
.B2(n_169),
.Y(n_271)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_216),
.Y(n_272)
);

CKINVDCx5p33_ASAP7_75t_R g273 ( 
.A(n_218),
.Y(n_273)
);

HB1xp67_ASAP7_75t_L g274 ( 
.A(n_240),
.Y(n_274)
);

CKINVDCx16_ASAP7_75t_R g275 ( 
.A(n_241),
.Y(n_275)
);

BUFx6f_ASAP7_75t_L g276 ( 
.A(n_231),
.Y(n_276)
);

INVx2_ASAP7_75t_L g277 ( 
.A(n_247),
.Y(n_277)
);

AND2x4_ASAP7_75t_L g278 ( 
.A(n_226),
.B(n_188),
.Y(n_278)
);

CKINVDCx5p33_ASAP7_75t_R g279 ( 
.A(n_223),
.Y(n_279)
);

CKINVDCx20_ASAP7_75t_R g280 ( 
.A(n_233),
.Y(n_280)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_224),
.Y(n_281)
);

CKINVDCx20_ASAP7_75t_R g282 ( 
.A(n_222),
.Y(n_282)
);

BUFx6f_ASAP7_75t_L g283 ( 
.A(n_232),
.Y(n_283)
);

CKINVDCx20_ASAP7_75t_R g284 ( 
.A(n_251),
.Y(n_284)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_221),
.Y(n_285)
);

INVx6_ASAP7_75t_L g286 ( 
.A(n_254),
.Y(n_286)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_260),
.Y(n_287)
);

INVx2_ASAP7_75t_L g288 ( 
.A(n_247),
.Y(n_288)
);

INVx2_ASAP7_75t_L g289 ( 
.A(n_247),
.Y(n_289)
);

CKINVDCx5p33_ASAP7_75t_R g290 ( 
.A(n_249),
.Y(n_290)
);

INVx2_ASAP7_75t_L g291 ( 
.A(n_247),
.Y(n_291)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_259),
.Y(n_292)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_234),
.Y(n_293)
);

NOR2xp33_ASAP7_75t_R g294 ( 
.A(n_252),
.B(n_161),
.Y(n_294)
);

CKINVDCx20_ASAP7_75t_R g295 ( 
.A(n_245),
.Y(n_295)
);

CKINVDCx5p33_ASAP7_75t_R g296 ( 
.A(n_258),
.Y(n_296)
);

AND2x2_ASAP7_75t_L g297 ( 
.A(n_256),
.B(n_200),
.Y(n_297)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_235),
.Y(n_298)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_236),
.Y(n_299)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_239),
.Y(n_300)
);

OAI21x1_ASAP7_75t_L g301 ( 
.A1(n_243),
.A2(n_203),
.B(n_155),
.Y(n_301)
);

CKINVDCx20_ASAP7_75t_R g302 ( 
.A(n_251),
.Y(n_302)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_248),
.Y(n_303)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_250),
.Y(n_304)
);

CKINVDCx20_ASAP7_75t_R g305 ( 
.A(n_245),
.Y(n_305)
);

CKINVDCx5p33_ASAP7_75t_R g306 ( 
.A(n_253),
.Y(n_306)
);

CKINVDCx5p33_ASAP7_75t_R g307 ( 
.A(n_255),
.Y(n_307)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_228),
.Y(n_308)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_242),
.Y(n_309)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_247),
.Y(n_310)
);

NAND2xp5_ASAP7_75t_L g311 ( 
.A(n_225),
.B(n_153),
.Y(n_311)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_220),
.Y(n_312)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_227),
.Y(n_313)
);

AND2x6_ASAP7_75t_L g314 ( 
.A(n_266),
.B(n_169),
.Y(n_314)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_264),
.Y(n_315)
);

NOR2xp33_ASAP7_75t_L g316 ( 
.A(n_308),
.B(n_238),
.Y(n_316)
);

OR2x2_ASAP7_75t_L g317 ( 
.A(n_274),
.B(n_262),
.Y(n_317)
);

INVx1_ASAP7_75t_SL g318 ( 
.A(n_286),
.Y(n_318)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_267),
.Y(n_319)
);

NAND2xp5_ASAP7_75t_L g320 ( 
.A(n_297),
.B(n_240),
.Y(n_320)
);

INVx3_ASAP7_75t_L g321 ( 
.A(n_269),
.Y(n_321)
);

NAND2xp5_ASAP7_75t_L g322 ( 
.A(n_310),
.B(n_270),
.Y(n_322)
);

INVx3_ASAP7_75t_L g323 ( 
.A(n_269),
.Y(n_323)
);

BUFx6f_ASAP7_75t_L g324 ( 
.A(n_269),
.Y(n_324)
);

AND2x4_ASAP7_75t_L g325 ( 
.A(n_268),
.B(n_257),
.Y(n_325)
);

AND2x2_ASAP7_75t_L g326 ( 
.A(n_286),
.B(n_229),
.Y(n_326)
);

AND2x2_ASAP7_75t_L g327 ( 
.A(n_286),
.B(n_229),
.Y(n_327)
);

NAND2xp5_ASAP7_75t_L g328 ( 
.A(n_268),
.B(n_266),
.Y(n_328)
);

BUFx2_ASAP7_75t_L g329 ( 
.A(n_273),
.Y(n_329)
);

AOI22xp5_ASAP7_75t_L g330 ( 
.A1(n_271),
.A2(n_211),
.B1(n_210),
.B2(n_209),
.Y(n_330)
);

INVx2_ASAP7_75t_L g331 ( 
.A(n_269),
.Y(n_331)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_272),
.Y(n_332)
);

INVx1_ASAP7_75t_SL g333 ( 
.A(n_280),
.Y(n_333)
);

INVx2_ASAP7_75t_L g334 ( 
.A(n_276),
.Y(n_334)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_281),
.Y(n_335)
);

AND2x4_ASAP7_75t_L g336 ( 
.A(n_278),
.B(n_199),
.Y(n_336)
);

NAND2xp5_ASAP7_75t_SL g337 ( 
.A(n_261),
.B(n_164),
.Y(n_337)
);

OR2x2_ASAP7_75t_L g338 ( 
.A(n_274),
.B(n_2),
.Y(n_338)
);

AND2x4_ASAP7_75t_L g339 ( 
.A(n_278),
.B(n_199),
.Y(n_339)
);

NAND2xp5_ASAP7_75t_SL g340 ( 
.A(n_261),
.B(n_165),
.Y(n_340)
);

AND2x2_ASAP7_75t_L g341 ( 
.A(n_262),
.B(n_168),
.Y(n_341)
);

INVx1_ASAP7_75t_L g342 ( 
.A(n_276),
.Y(n_342)
);

NAND2xp5_ASAP7_75t_L g343 ( 
.A(n_309),
.B(n_312),
.Y(n_343)
);

INVx1_ASAP7_75t_L g344 ( 
.A(n_276),
.Y(n_344)
);

AO22x2_ASAP7_75t_L g345 ( 
.A1(n_285),
.A2(n_2),
.B1(n_3),
.B2(n_4),
.Y(n_345)
);

INVx4_ASAP7_75t_L g346 ( 
.A(n_276),
.Y(n_346)
);

AOI22xp5_ASAP7_75t_L g347 ( 
.A1(n_313),
.A2(n_207),
.B1(n_206),
.B2(n_205),
.Y(n_347)
);

NOR2xp33_ASAP7_75t_L g348 ( 
.A(n_290),
.B(n_296),
.Y(n_348)
);

BUFx2_ASAP7_75t_L g349 ( 
.A(n_279),
.Y(n_349)
);

BUFx4f_ASAP7_75t_L g350 ( 
.A(n_265),
.Y(n_350)
);

NOR2xp33_ASAP7_75t_L g351 ( 
.A(n_287),
.B(n_175),
.Y(n_351)
);

NAND2xp33_ASAP7_75t_L g352 ( 
.A(n_263),
.B(n_183),
.Y(n_352)
);

NAND2xp5_ASAP7_75t_L g353 ( 
.A(n_283),
.B(n_263),
.Y(n_353)
);

INVx1_ASAP7_75t_L g354 ( 
.A(n_283),
.Y(n_354)
);

INVx1_ASAP7_75t_L g355 ( 
.A(n_283),
.Y(n_355)
);

BUFx2_ASAP7_75t_L g356 ( 
.A(n_284),
.Y(n_356)
);

BUFx6f_ASAP7_75t_L g357 ( 
.A(n_283),
.Y(n_357)
);

INVx8_ASAP7_75t_L g358 ( 
.A(n_263),
.Y(n_358)
);

OAI22xp5_ASAP7_75t_L g359 ( 
.A1(n_292),
.A2(n_204),
.B1(n_201),
.B2(n_198),
.Y(n_359)
);

INVx2_ASAP7_75t_L g360 ( 
.A(n_277),
.Y(n_360)
);

INVxp67_ASAP7_75t_L g361 ( 
.A(n_306),
.Y(n_361)
);

INVx1_ASAP7_75t_L g362 ( 
.A(n_293),
.Y(n_362)
);

INVx1_ASAP7_75t_L g363 ( 
.A(n_298),
.Y(n_363)
);

NAND2xp5_ASAP7_75t_L g364 ( 
.A(n_263),
.B(n_184),
.Y(n_364)
);

INVx1_ASAP7_75t_SL g365 ( 
.A(n_307),
.Y(n_365)
);

INVx1_ASAP7_75t_L g366 ( 
.A(n_299),
.Y(n_366)
);

INVx2_ASAP7_75t_L g367 ( 
.A(n_288),
.Y(n_367)
);

NOR2xp33_ASAP7_75t_L g368 ( 
.A(n_300),
.B(n_186),
.Y(n_368)
);

INVx1_ASAP7_75t_L g369 ( 
.A(n_303),
.Y(n_369)
);

INVx1_ASAP7_75t_SL g370 ( 
.A(n_295),
.Y(n_370)
);

CKINVDCx5p33_ASAP7_75t_R g371 ( 
.A(n_294),
.Y(n_371)
);

BUFx6f_ASAP7_75t_L g372 ( 
.A(n_301),
.Y(n_372)
);

INVx1_ASAP7_75t_SL g373 ( 
.A(n_295),
.Y(n_373)
);

INVx2_ASAP7_75t_L g374 ( 
.A(n_289),
.Y(n_374)
);

INVx2_ASAP7_75t_L g375 ( 
.A(n_291),
.Y(n_375)
);

INVx2_ASAP7_75t_L g376 ( 
.A(n_304),
.Y(n_376)
);

NAND2x1p5_ASAP7_75t_L g377 ( 
.A(n_311),
.B(n_199),
.Y(n_377)
);

INVx1_ASAP7_75t_L g378 ( 
.A(n_263),
.Y(n_378)
);

HB1xp67_ASAP7_75t_L g379 ( 
.A(n_275),
.Y(n_379)
);

AND3x2_ASAP7_75t_L g380 ( 
.A(n_282),
.B(n_3),
.C(n_4),
.Y(n_380)
);

INVx1_ASAP7_75t_L g381 ( 
.A(n_294),
.Y(n_381)
);

INVx2_ASAP7_75t_L g382 ( 
.A(n_376),
.Y(n_382)
);

NAND2xp5_ASAP7_75t_SL g383 ( 
.A(n_371),
.B(n_302),
.Y(n_383)
);

AND2x4_ASAP7_75t_L g384 ( 
.A(n_318),
.B(n_305),
.Y(n_384)
);

AOI22xp33_ASAP7_75t_L g385 ( 
.A1(n_345),
.A2(n_282),
.B1(n_305),
.B2(n_196),
.Y(n_385)
);

NAND2xp5_ASAP7_75t_L g386 ( 
.A(n_316),
.B(n_189),
.Y(n_386)
);

OAI21xp5_ASAP7_75t_L g387 ( 
.A1(n_322),
.A2(n_195),
.B(n_193),
.Y(n_387)
);

NAND2xp5_ASAP7_75t_L g388 ( 
.A(n_314),
.B(n_192),
.Y(n_388)
);

INVx1_ASAP7_75t_L g389 ( 
.A(n_315),
.Y(n_389)
);

INVx4_ASAP7_75t_L g390 ( 
.A(n_358),
.Y(n_390)
);

AOI22xp33_ASAP7_75t_L g391 ( 
.A1(n_345),
.A2(n_5),
.B1(n_6),
.B2(n_7),
.Y(n_391)
);

A2O1A1Ixp33_ASAP7_75t_SL g392 ( 
.A1(n_351),
.A2(n_5),
.B(n_8),
.C(n_9),
.Y(n_392)
);

OR2x2_ASAP7_75t_L g393 ( 
.A(n_317),
.B(n_8),
.Y(n_393)
);

AND2x4_ASAP7_75t_SL g394 ( 
.A(n_326),
.B(n_9),
.Y(n_394)
);

NOR2xp33_ASAP7_75t_SL g395 ( 
.A(n_348),
.B(n_10),
.Y(n_395)
);

INVx2_ASAP7_75t_L g396 ( 
.A(n_324),
.Y(n_396)
);

NAND2xp5_ASAP7_75t_SL g397 ( 
.A(n_350),
.B(n_11),
.Y(n_397)
);

AND2x2_ASAP7_75t_SL g398 ( 
.A(n_350),
.B(n_11),
.Y(n_398)
);

AND2x6_ASAP7_75t_SL g399 ( 
.A(n_325),
.B(n_13),
.Y(n_399)
);

AND2x2_ASAP7_75t_L g400 ( 
.A(n_318),
.B(n_13),
.Y(n_400)
);

NAND2xp5_ASAP7_75t_SL g401 ( 
.A(n_381),
.B(n_15),
.Y(n_401)
);

INVx1_ASAP7_75t_L g402 ( 
.A(n_319),
.Y(n_402)
);

AND2x6_ASAP7_75t_L g403 ( 
.A(n_378),
.B(n_18),
.Y(n_403)
);

AOI22xp33_ASAP7_75t_L g404 ( 
.A1(n_314),
.A2(n_15),
.B1(n_16),
.B2(n_17),
.Y(n_404)
);

OAI22xp5_ASAP7_75t_L g405 ( 
.A1(n_328),
.A2(n_17),
.B1(n_19),
.B2(n_20),
.Y(n_405)
);

NAND2xp5_ASAP7_75t_L g406 ( 
.A(n_314),
.B(n_141),
.Y(n_406)
);

INVx1_ASAP7_75t_L g407 ( 
.A(n_332),
.Y(n_407)
);

NAND2xp5_ASAP7_75t_L g408 ( 
.A(n_314),
.B(n_21),
.Y(n_408)
);

NAND2xp5_ASAP7_75t_L g409 ( 
.A(n_336),
.B(n_140),
.Y(n_409)
);

INVx2_ASAP7_75t_L g410 ( 
.A(n_324),
.Y(n_410)
);

INVx1_ASAP7_75t_L g411 ( 
.A(n_335),
.Y(n_411)
);

INVx2_ASAP7_75t_L g412 ( 
.A(n_324),
.Y(n_412)
);

INVx2_ASAP7_75t_L g413 ( 
.A(n_357),
.Y(n_413)
);

AOI21xp5_ASAP7_75t_L g414 ( 
.A1(n_322),
.A2(n_22),
.B(n_24),
.Y(n_414)
);

NAND2xp5_ASAP7_75t_L g415 ( 
.A(n_336),
.B(n_25),
.Y(n_415)
);

INVx1_ASAP7_75t_L g416 ( 
.A(n_362),
.Y(n_416)
);

NAND2xp5_ASAP7_75t_SL g417 ( 
.A(n_372),
.B(n_26),
.Y(n_417)
);

AOI22xp5_ASAP7_75t_L g418 ( 
.A1(n_320),
.A2(n_27),
.B1(n_29),
.B2(n_30),
.Y(n_418)
);

INVx3_ASAP7_75t_L g419 ( 
.A(n_346),
.Y(n_419)
);

NAND2xp5_ASAP7_75t_L g420 ( 
.A(n_339),
.B(n_139),
.Y(n_420)
);

NAND2xp5_ASAP7_75t_L g421 ( 
.A(n_339),
.B(n_31),
.Y(n_421)
);

AND2x2_ASAP7_75t_L g422 ( 
.A(n_341),
.B(n_32),
.Y(n_422)
);

NOR2xp33_ASAP7_75t_L g423 ( 
.A(n_343),
.B(n_35),
.Y(n_423)
);

OR2x6_ASAP7_75t_L g424 ( 
.A(n_329),
.B(n_349),
.Y(n_424)
);

NAND2xp5_ASAP7_75t_L g425 ( 
.A(n_363),
.B(n_138),
.Y(n_425)
);

INVx1_ASAP7_75t_L g426 ( 
.A(n_366),
.Y(n_426)
);

CKINVDCx5p33_ASAP7_75t_R g427 ( 
.A(n_365),
.Y(n_427)
);

INVx2_ASAP7_75t_L g428 ( 
.A(n_357),
.Y(n_428)
);

INVx1_ASAP7_75t_L g429 ( 
.A(n_369),
.Y(n_429)
);

INVx2_ASAP7_75t_SL g430 ( 
.A(n_379),
.Y(n_430)
);

NAND2xp5_ASAP7_75t_L g431 ( 
.A(n_368),
.B(n_346),
.Y(n_431)
);

INVx2_ASAP7_75t_SL g432 ( 
.A(n_327),
.Y(n_432)
);

INVx2_ASAP7_75t_L g433 ( 
.A(n_357),
.Y(n_433)
);

NAND2xp5_ASAP7_75t_SL g434 ( 
.A(n_372),
.B(n_36),
.Y(n_434)
);

INVx2_ASAP7_75t_L g435 ( 
.A(n_321),
.Y(n_435)
);

INVx1_ASAP7_75t_L g436 ( 
.A(n_342),
.Y(n_436)
);

AOI22xp5_ASAP7_75t_L g437 ( 
.A1(n_330),
.A2(n_352),
.B1(n_323),
.B2(n_321),
.Y(n_437)
);

AND2x2_ASAP7_75t_SL g438 ( 
.A(n_330),
.B(n_136),
.Y(n_438)
);

INVx2_ASAP7_75t_SL g439 ( 
.A(n_325),
.Y(n_439)
);

AOI22xp33_ASAP7_75t_L g440 ( 
.A1(n_358),
.A2(n_39),
.B1(n_40),
.B2(n_42),
.Y(n_440)
);

INVxp67_ASAP7_75t_L g441 ( 
.A(n_356),
.Y(n_441)
);

INVx2_ASAP7_75t_SL g442 ( 
.A(n_333),
.Y(n_442)
);

INVx2_ASAP7_75t_L g443 ( 
.A(n_323),
.Y(n_443)
);

INVx1_ASAP7_75t_L g444 ( 
.A(n_344),
.Y(n_444)
);

AOI22xp33_ASAP7_75t_L g445 ( 
.A1(n_358),
.A2(n_43),
.B1(n_46),
.B2(n_48),
.Y(n_445)
);

INVx2_ASAP7_75t_SL g446 ( 
.A(n_333),
.Y(n_446)
);

INVx4_ASAP7_75t_L g447 ( 
.A(n_372),
.Y(n_447)
);

INVxp67_ASAP7_75t_L g448 ( 
.A(n_370),
.Y(n_448)
);

INVx3_ASAP7_75t_L g449 ( 
.A(n_447),
.Y(n_449)
);

NAND2xp5_ASAP7_75t_L g450 ( 
.A(n_386),
.B(n_347),
.Y(n_450)
);

NOR2xp33_ASAP7_75t_L g451 ( 
.A(n_427),
.B(n_365),
.Y(n_451)
);

INVx2_ASAP7_75t_L g452 ( 
.A(n_436),
.Y(n_452)
);

NOR2xp33_ASAP7_75t_L g453 ( 
.A(n_448),
.B(n_370),
.Y(n_453)
);

NAND2x1p5_ASAP7_75t_L g454 ( 
.A(n_390),
.B(n_355),
.Y(n_454)
);

NOR2xp67_ASAP7_75t_L g455 ( 
.A(n_442),
.B(n_361),
.Y(n_455)
);

NAND2xp5_ASAP7_75t_L g456 ( 
.A(n_389),
.B(n_347),
.Y(n_456)
);

INVx1_ASAP7_75t_L g457 ( 
.A(n_402),
.Y(n_457)
);

HB1xp67_ASAP7_75t_L g458 ( 
.A(n_446),
.Y(n_458)
);

NOR2xp33_ASAP7_75t_L g459 ( 
.A(n_448),
.B(n_373),
.Y(n_459)
);

INVx2_ASAP7_75t_L g460 ( 
.A(n_444),
.Y(n_460)
);

CKINVDCx20_ASAP7_75t_R g461 ( 
.A(n_424),
.Y(n_461)
);

AND2x4_ASAP7_75t_L g462 ( 
.A(n_390),
.B(n_373),
.Y(n_462)
);

INVx1_ASAP7_75t_L g463 ( 
.A(n_407),
.Y(n_463)
);

BUFx2_ASAP7_75t_L g464 ( 
.A(n_384),
.Y(n_464)
);

INVx1_ASAP7_75t_L g465 ( 
.A(n_411),
.Y(n_465)
);

NOR2xp33_ASAP7_75t_L g466 ( 
.A(n_441),
.B(n_338),
.Y(n_466)
);

INVx1_ASAP7_75t_L g467 ( 
.A(n_416),
.Y(n_467)
);

INVx3_ASAP7_75t_L g468 ( 
.A(n_447),
.Y(n_468)
);

INVx1_ASAP7_75t_L g469 ( 
.A(n_426),
.Y(n_469)
);

INVx2_ASAP7_75t_L g470 ( 
.A(n_382),
.Y(n_470)
);

CKINVDCx5p33_ASAP7_75t_R g471 ( 
.A(n_424),
.Y(n_471)
);

AND2x2_ASAP7_75t_L g472 ( 
.A(n_438),
.B(n_377),
.Y(n_472)
);

BUFx2_ASAP7_75t_L g473 ( 
.A(n_384),
.Y(n_473)
);

NAND2x1p5_ASAP7_75t_L g474 ( 
.A(n_419),
.B(n_354),
.Y(n_474)
);

BUFx3_ASAP7_75t_L g475 ( 
.A(n_424),
.Y(n_475)
);

INVx1_ASAP7_75t_L g476 ( 
.A(n_429),
.Y(n_476)
);

OR2x6_ASAP7_75t_SL g477 ( 
.A(n_438),
.B(n_359),
.Y(n_477)
);

NOR2xp67_ASAP7_75t_L g478 ( 
.A(n_430),
.B(n_359),
.Y(n_478)
);

INVx1_ASAP7_75t_L g479 ( 
.A(n_435),
.Y(n_479)
);

NAND2xp5_ASAP7_75t_SL g480 ( 
.A(n_423),
.B(n_360),
.Y(n_480)
);

INVx3_ASAP7_75t_L g481 ( 
.A(n_403),
.Y(n_481)
);

INVx2_ASAP7_75t_L g482 ( 
.A(n_443),
.Y(n_482)
);

INVx3_ASAP7_75t_L g483 ( 
.A(n_403),
.Y(n_483)
);

AND2x4_ASAP7_75t_L g484 ( 
.A(n_439),
.B(n_331),
.Y(n_484)
);

AO22x1_ASAP7_75t_L g485 ( 
.A1(n_441),
.A2(n_380),
.B1(n_353),
.B2(n_364),
.Y(n_485)
);

AND2x4_ASAP7_75t_L g486 ( 
.A(n_432),
.B(n_334),
.Y(n_486)
);

INVx1_ASAP7_75t_L g487 ( 
.A(n_396),
.Y(n_487)
);

INVxp67_ASAP7_75t_L g488 ( 
.A(n_395),
.Y(n_488)
);

HB1xp67_ASAP7_75t_L g489 ( 
.A(n_400),
.Y(n_489)
);

AND2x4_ASAP7_75t_L g490 ( 
.A(n_422),
.B(n_419),
.Y(n_490)
);

BUFx6f_ASAP7_75t_L g491 ( 
.A(n_403),
.Y(n_491)
);

INVx1_ASAP7_75t_L g492 ( 
.A(n_410),
.Y(n_492)
);

BUFx12f_ASAP7_75t_L g493 ( 
.A(n_471),
.Y(n_493)
);

AO31x2_ASAP7_75t_L g494 ( 
.A1(n_450),
.A2(n_423),
.A3(n_425),
.B(n_414),
.Y(n_494)
);

INVx1_ASAP7_75t_L g495 ( 
.A(n_457),
.Y(n_495)
);

OAI21x1_ASAP7_75t_L g496 ( 
.A1(n_481),
.A2(n_483),
.B(n_417),
.Y(n_496)
);

AOI21xp5_ASAP7_75t_L g497 ( 
.A1(n_480),
.A2(n_431),
.B(n_417),
.Y(n_497)
);

NAND2xp5_ASAP7_75t_L g498 ( 
.A(n_451),
.B(n_398),
.Y(n_498)
);

NAND2xp5_ASAP7_75t_SL g499 ( 
.A(n_455),
.B(n_398),
.Y(n_499)
);

OAI21x1_ASAP7_75t_L g500 ( 
.A1(n_481),
.A2(n_483),
.B(n_434),
.Y(n_500)
);

NAND3xp33_ASAP7_75t_SL g501 ( 
.A(n_488),
.B(n_391),
.C(n_404),
.Y(n_501)
);

NAND2x1p5_ASAP7_75t_L g502 ( 
.A(n_475),
.B(n_383),
.Y(n_502)
);

NAND2xp5_ASAP7_75t_L g503 ( 
.A(n_456),
.B(n_393),
.Y(n_503)
);

AOI22xp33_ASAP7_75t_L g504 ( 
.A1(n_464),
.A2(n_385),
.B1(n_473),
.B2(n_459),
.Y(n_504)
);

AOI21xp33_ASAP7_75t_L g505 ( 
.A1(n_453),
.A2(n_387),
.B(n_388),
.Y(n_505)
);

OAI21xp5_ASAP7_75t_L g506 ( 
.A1(n_480),
.A2(n_434),
.B(n_437),
.Y(n_506)
);

AOI21x1_ASAP7_75t_L g507 ( 
.A1(n_490),
.A2(n_409),
.B(n_415),
.Y(n_507)
);

NAND2xp5_ASAP7_75t_L g508 ( 
.A(n_477),
.B(n_397),
.Y(n_508)
);

AND2x4_ASAP7_75t_L g509 ( 
.A(n_475),
.B(n_394),
.Y(n_509)
);

NAND2xp5_ASAP7_75t_SL g510 ( 
.A(n_478),
.B(n_397),
.Y(n_510)
);

AOI21x1_ASAP7_75t_L g511 ( 
.A1(n_490),
.A2(n_420),
.B(n_421),
.Y(n_511)
);

NOR2x1_ASAP7_75t_SL g512 ( 
.A(n_491),
.B(n_406),
.Y(n_512)
);

AOI21xp5_ASAP7_75t_L g513 ( 
.A1(n_490),
.A2(n_414),
.B(n_375),
.Y(n_513)
);

OAI21xp5_ASAP7_75t_L g514 ( 
.A1(n_463),
.A2(n_401),
.B(n_367),
.Y(n_514)
);

AOI21xp33_ASAP7_75t_L g515 ( 
.A1(n_466),
.A2(n_385),
.B(n_401),
.Y(n_515)
);

AO31x2_ASAP7_75t_L g516 ( 
.A1(n_452),
.A2(n_460),
.A3(n_470),
.B(n_482),
.Y(n_516)
);

AO31x2_ASAP7_75t_L g517 ( 
.A1(n_452),
.A2(n_408),
.A3(n_374),
.B(n_405),
.Y(n_517)
);

OAI21x1_ASAP7_75t_L g518 ( 
.A1(n_481),
.A2(n_412),
.B(n_413),
.Y(n_518)
);

INVx6_ASAP7_75t_L g519 ( 
.A(n_462),
.Y(n_519)
);

OAI21xp5_ASAP7_75t_L g520 ( 
.A1(n_465),
.A2(n_404),
.B(n_418),
.Y(n_520)
);

OAI21xp33_ASAP7_75t_SL g521 ( 
.A1(n_477),
.A2(n_391),
.B(n_440),
.Y(n_521)
);

BUFx3_ASAP7_75t_L g522 ( 
.A(n_461),
.Y(n_522)
);

AND2x2_ASAP7_75t_L g523 ( 
.A(n_521),
.B(n_472),
.Y(n_523)
);

NOR2x1_ASAP7_75t_L g524 ( 
.A(n_510),
.B(n_449),
.Y(n_524)
);

NAND2xp5_ASAP7_75t_L g525 ( 
.A(n_503),
.B(n_458),
.Y(n_525)
);

OA21x2_ASAP7_75t_L g526 ( 
.A1(n_506),
.A2(n_445),
.B(n_440),
.Y(n_526)
);

INVx2_ASAP7_75t_L g527 ( 
.A(n_516),
.Y(n_527)
);

AOI21xp5_ASAP7_75t_L g528 ( 
.A1(n_497),
.A2(n_483),
.B(n_491),
.Y(n_528)
);

OAI21x1_ASAP7_75t_L g529 ( 
.A1(n_496),
.A2(n_449),
.B(n_468),
.Y(n_529)
);

INVx1_ASAP7_75t_L g530 ( 
.A(n_516),
.Y(n_530)
);

AND2x2_ASAP7_75t_L g531 ( 
.A(n_521),
.B(n_472),
.Y(n_531)
);

AOI21xp5_ASAP7_75t_L g532 ( 
.A1(n_506),
.A2(n_491),
.B(n_468),
.Y(n_532)
);

BUFx6f_ASAP7_75t_L g533 ( 
.A(n_519),
.Y(n_533)
);

INVx2_ASAP7_75t_L g534 ( 
.A(n_516),
.Y(n_534)
);

AOI22xp33_ASAP7_75t_L g535 ( 
.A1(n_501),
.A2(n_473),
.B1(n_464),
.B2(n_489),
.Y(n_535)
);

AO21x2_ASAP7_75t_L g536 ( 
.A1(n_513),
.A2(n_392),
.B(n_492),
.Y(n_536)
);

INVx3_ASAP7_75t_L g537 ( 
.A(n_500),
.Y(n_537)
);

NAND2xp5_ASAP7_75t_L g538 ( 
.A(n_498),
.B(n_462),
.Y(n_538)
);

OAI21x1_ASAP7_75t_L g539 ( 
.A1(n_507),
.A2(n_449),
.B(n_468),
.Y(n_539)
);

OAI21x1_ASAP7_75t_L g540 ( 
.A1(n_511),
.A2(n_474),
.B(n_454),
.Y(n_540)
);

HB1xp67_ASAP7_75t_L g541 ( 
.A(n_522),
.Y(n_541)
);

OAI21x1_ASAP7_75t_L g542 ( 
.A1(n_518),
.A2(n_474),
.B(n_454),
.Y(n_542)
);

OAI21x1_ASAP7_75t_L g543 ( 
.A1(n_514),
.A2(n_460),
.B(n_445),
.Y(n_543)
);

AOI21xp5_ASAP7_75t_L g544 ( 
.A1(n_520),
.A2(n_491),
.B(n_469),
.Y(n_544)
);

OAI22xp5_ASAP7_75t_SL g545 ( 
.A1(n_508),
.A2(n_461),
.B1(n_471),
.B2(n_399),
.Y(n_545)
);

O2A1O1Ixp33_ASAP7_75t_SL g546 ( 
.A1(n_505),
.A2(n_392),
.B(n_467),
.C(n_476),
.Y(n_546)
);

INVx2_ASAP7_75t_L g547 ( 
.A(n_517),
.Y(n_547)
);

OAI21x1_ASAP7_75t_L g548 ( 
.A1(n_514),
.A2(n_482),
.B(n_428),
.Y(n_548)
);

OAI21xp5_ASAP7_75t_L g549 ( 
.A1(n_520),
.A2(n_479),
.B(n_403),
.Y(n_549)
);

AND2x2_ASAP7_75t_L g550 ( 
.A(n_525),
.B(n_509),
.Y(n_550)
);

INVx2_ASAP7_75t_L g551 ( 
.A(n_530),
.Y(n_551)
);

BUFx6f_ASAP7_75t_L g552 ( 
.A(n_533),
.Y(n_552)
);

OR2x2_ASAP7_75t_L g553 ( 
.A(n_523),
.B(n_495),
.Y(n_553)
);

AOI22xp33_ASAP7_75t_L g554 ( 
.A1(n_526),
.A2(n_515),
.B1(n_504),
.B2(n_519),
.Y(n_554)
);

INVx1_ASAP7_75t_L g555 ( 
.A(n_530),
.Y(n_555)
);

OAI21x1_ASAP7_75t_L g556 ( 
.A1(n_539),
.A2(n_433),
.B(n_487),
.Y(n_556)
);

INVx1_ASAP7_75t_SL g557 ( 
.A(n_541),
.Y(n_557)
);

INVx1_ASAP7_75t_SL g558 ( 
.A(n_533),
.Y(n_558)
);

OAI221xp5_ASAP7_75t_L g559 ( 
.A1(n_545),
.A2(n_499),
.B1(n_535),
.B2(n_502),
.C(n_538),
.Y(n_559)
);

INVx1_ASAP7_75t_L g560 ( 
.A(n_527),
.Y(n_560)
);

INVx4_ASAP7_75t_SL g561 ( 
.A(n_533),
.Y(n_561)
);

OA21x2_ASAP7_75t_L g562 ( 
.A1(n_547),
.A2(n_470),
.B(n_494),
.Y(n_562)
);

CKINVDCx5p33_ASAP7_75t_R g563 ( 
.A(n_545),
.Y(n_563)
);

OAI221xp5_ASAP7_75t_L g564 ( 
.A1(n_549),
.A2(n_337),
.B1(n_340),
.B2(n_485),
.C(n_494),
.Y(n_564)
);

AND2x4_ASAP7_75t_L g565 ( 
.A(n_533),
.B(n_509),
.Y(n_565)
);

OR2x6_ASAP7_75t_SL g566 ( 
.A(n_523),
.B(n_493),
.Y(n_566)
);

NAND2xp5_ASAP7_75t_L g567 ( 
.A(n_533),
.B(n_462),
.Y(n_567)
);

BUFx4f_ASAP7_75t_L g568 ( 
.A(n_531),
.Y(n_568)
);

CKINVDCx5p33_ASAP7_75t_R g569 ( 
.A(n_544),
.Y(n_569)
);

OAI22xp33_ASAP7_75t_L g570 ( 
.A1(n_526),
.A2(n_484),
.B1(n_486),
.B2(n_494),
.Y(n_570)
);

BUFx12f_ASAP7_75t_L g571 ( 
.A(n_531),
.Y(n_571)
);

AOI22xp33_ASAP7_75t_SL g572 ( 
.A1(n_526),
.A2(n_549),
.B1(n_543),
.B2(n_512),
.Y(n_572)
);

AOI21xp5_ASAP7_75t_L g573 ( 
.A1(n_526),
.A2(n_517),
.B(n_486),
.Y(n_573)
);

NAND2xp33_ASAP7_75t_SL g574 ( 
.A(n_536),
.B(n_486),
.Y(n_574)
);

OAI22xp5_ASAP7_75t_L g575 ( 
.A1(n_524),
.A2(n_484),
.B1(n_517),
.B2(n_403),
.Y(n_575)
);

NAND2xp5_ASAP7_75t_L g576 ( 
.A(n_524),
.B(n_484),
.Y(n_576)
);

AOI22xp5_ASAP7_75t_L g577 ( 
.A1(n_532),
.A2(n_49),
.B1(n_50),
.B2(n_51),
.Y(n_577)
);

AOI21xp5_ASAP7_75t_L g578 ( 
.A1(n_528),
.A2(n_134),
.B(n_57),
.Y(n_578)
);

AOI221xp5_ASAP7_75t_L g579 ( 
.A1(n_546),
.A2(n_55),
.B1(n_58),
.B2(n_61),
.C(n_62),
.Y(n_579)
);

OR2x2_ASAP7_75t_L g580 ( 
.A(n_527),
.B(n_67),
.Y(n_580)
);

INVx1_ASAP7_75t_L g581 ( 
.A(n_527),
.Y(n_581)
);

AND2x2_ASAP7_75t_L g582 ( 
.A(n_568),
.B(n_534),
.Y(n_582)
);

OAI211xp5_ASAP7_75t_L g583 ( 
.A1(n_579),
.A2(n_537),
.B(n_547),
.C(n_543),
.Y(n_583)
);

AND2x4_ASAP7_75t_SL g584 ( 
.A(n_552),
.B(n_534),
.Y(n_584)
);

INVx1_ASAP7_75t_L g585 ( 
.A(n_553),
.Y(n_585)
);

AOI22xp33_ASAP7_75t_L g586 ( 
.A1(n_554),
.A2(n_534),
.B1(n_547),
.B2(n_536),
.Y(n_586)
);

AOI221xp5_ASAP7_75t_L g587 ( 
.A1(n_563),
.A2(n_564),
.B1(n_559),
.B2(n_570),
.C(n_557),
.Y(n_587)
);

AND2x2_ASAP7_75t_L g588 ( 
.A(n_568),
.B(n_537),
.Y(n_588)
);

BUFx2_ASAP7_75t_L g589 ( 
.A(n_571),
.Y(n_589)
);

NAND2xp33_ASAP7_75t_L g590 ( 
.A(n_569),
.B(n_537),
.Y(n_590)
);

OAI22xp33_ASAP7_75t_SL g591 ( 
.A1(n_566),
.A2(n_537),
.B1(n_536),
.B2(n_548),
.Y(n_591)
);

AOI21xp5_ASAP7_75t_L g592 ( 
.A1(n_574),
.A2(n_540),
.B(n_539),
.Y(n_592)
);

BUFx2_ASAP7_75t_L g593 ( 
.A(n_562),
.Y(n_593)
);

AOI22xp33_ASAP7_75t_L g594 ( 
.A1(n_550),
.A2(n_548),
.B1(n_540),
.B2(n_542),
.Y(n_594)
);

AND2x2_ASAP7_75t_L g595 ( 
.A(n_555),
.B(n_529),
.Y(n_595)
);

AOI21xp5_ASAP7_75t_L g596 ( 
.A1(n_575),
.A2(n_529),
.B(n_542),
.Y(n_596)
);

NAND2xp5_ASAP7_75t_L g597 ( 
.A(n_558),
.B(n_69),
.Y(n_597)
);

OAI211xp5_ASAP7_75t_L g598 ( 
.A1(n_577),
.A2(n_70),
.B(n_72),
.C(n_74),
.Y(n_598)
);

OAI22xp5_ASAP7_75t_L g599 ( 
.A1(n_567),
.A2(n_75),
.B1(n_76),
.B2(n_79),
.Y(n_599)
);

OAI21xp5_ASAP7_75t_SL g600 ( 
.A1(n_572),
.A2(n_578),
.B(n_565),
.Y(n_600)
);

INVx4_ASAP7_75t_L g601 ( 
.A(n_552),
.Y(n_601)
);

NAND2xp5_ASAP7_75t_L g602 ( 
.A(n_552),
.B(n_81),
.Y(n_602)
);

CKINVDCx5p33_ASAP7_75t_R g603 ( 
.A(n_565),
.Y(n_603)
);

AOI22xp33_ASAP7_75t_L g604 ( 
.A1(n_576),
.A2(n_83),
.B1(n_84),
.B2(n_86),
.Y(n_604)
);

HB1xp67_ASAP7_75t_L g605 ( 
.A(n_595),
.Y(n_605)
);

NAND2xp5_ASAP7_75t_L g606 ( 
.A(n_585),
.B(n_573),
.Y(n_606)
);

HB1xp67_ASAP7_75t_L g607 ( 
.A(n_595),
.Y(n_607)
);

INVx1_ASAP7_75t_L g608 ( 
.A(n_582),
.Y(n_608)
);

INVx2_ASAP7_75t_L g609 ( 
.A(n_593),
.Y(n_609)
);

AND2x2_ASAP7_75t_L g610 ( 
.A(n_589),
.B(n_561),
.Y(n_610)
);

AND2x2_ASAP7_75t_L g611 ( 
.A(n_588),
.B(n_561),
.Y(n_611)
);

BUFx2_ASAP7_75t_L g612 ( 
.A(n_588),
.Y(n_612)
);

NAND2xp5_ASAP7_75t_L g613 ( 
.A(n_590),
.B(n_562),
.Y(n_613)
);

AOI22xp33_ASAP7_75t_L g614 ( 
.A1(n_587),
.A2(n_580),
.B1(n_551),
.B2(n_581),
.Y(n_614)
);

AO31x2_ASAP7_75t_L g615 ( 
.A1(n_593),
.A2(n_581),
.A3(n_560),
.B(n_556),
.Y(n_615)
);

NAND2xp5_ASAP7_75t_L g616 ( 
.A(n_590),
.B(n_87),
.Y(n_616)
);

INVx2_ASAP7_75t_L g617 ( 
.A(n_582),
.Y(n_617)
);

OR2x2_ASAP7_75t_L g618 ( 
.A(n_586),
.B(n_88),
.Y(n_618)
);

INVx1_ASAP7_75t_L g619 ( 
.A(n_584),
.Y(n_619)
);

AOI221xp5_ASAP7_75t_L g620 ( 
.A1(n_606),
.A2(n_583),
.B1(n_591),
.B2(n_600),
.C(n_599),
.Y(n_620)
);

OAI22xp5_ASAP7_75t_L g621 ( 
.A1(n_616),
.A2(n_598),
.B1(n_604),
.B2(n_601),
.Y(n_621)
);

INVx2_ASAP7_75t_L g622 ( 
.A(n_609),
.Y(n_622)
);

INVx2_ASAP7_75t_L g623 ( 
.A(n_617),
.Y(n_623)
);

AND2x2_ASAP7_75t_L g624 ( 
.A(n_612),
.B(n_601),
.Y(n_624)
);

NAND3xp33_ASAP7_75t_L g625 ( 
.A(n_614),
.B(n_596),
.C(n_601),
.Y(n_625)
);

INVx2_ASAP7_75t_L g626 ( 
.A(n_608),
.Y(n_626)
);

AND2x2_ASAP7_75t_L g627 ( 
.A(n_605),
.B(n_603),
.Y(n_627)
);

NAND2xp5_ASAP7_75t_L g628 ( 
.A(n_626),
.B(n_605),
.Y(n_628)
);

INVx1_ASAP7_75t_L g629 ( 
.A(n_622),
.Y(n_629)
);

NOR2xp33_ASAP7_75t_L g630 ( 
.A(n_627),
.B(n_610),
.Y(n_630)
);

INVxp67_ASAP7_75t_L g631 ( 
.A(n_624),
.Y(n_631)
);

NAND2x1p5_ASAP7_75t_L g632 ( 
.A(n_623),
.B(n_616),
.Y(n_632)
);

INVx1_ASAP7_75t_L g633 ( 
.A(n_625),
.Y(n_633)
);

AND2x2_ASAP7_75t_L g634 ( 
.A(n_625),
.B(n_607),
.Y(n_634)
);

NAND2xp5_ASAP7_75t_L g635 ( 
.A(n_633),
.B(n_620),
.Y(n_635)
);

AND2x2_ASAP7_75t_L g636 ( 
.A(n_634),
.B(n_611),
.Y(n_636)
);

INVx2_ASAP7_75t_L g637 ( 
.A(n_632),
.Y(n_637)
);

INVx1_ASAP7_75t_L g638 ( 
.A(n_628),
.Y(n_638)
);

NAND2xp5_ASAP7_75t_L g639 ( 
.A(n_632),
.B(n_606),
.Y(n_639)
);

OAI21xp33_ASAP7_75t_L g640 ( 
.A1(n_635),
.A2(n_631),
.B(n_630),
.Y(n_640)
);

NOR2x1p5_ASAP7_75t_L g641 ( 
.A(n_635),
.B(n_613),
.Y(n_641)
);

INVx2_ASAP7_75t_L g642 ( 
.A(n_637),
.Y(n_642)
);

OR2x2_ASAP7_75t_L g643 ( 
.A(n_638),
.B(n_629),
.Y(n_643)
);

OR2x2_ASAP7_75t_L g644 ( 
.A(n_639),
.B(n_619),
.Y(n_644)
);

OAI21xp5_ASAP7_75t_SL g645 ( 
.A1(n_640),
.A2(n_621),
.B(n_636),
.Y(n_645)
);

HB1xp67_ASAP7_75t_L g646 ( 
.A(n_644),
.Y(n_646)
);

INVx1_ASAP7_75t_L g647 ( 
.A(n_643),
.Y(n_647)
);

INVx1_ASAP7_75t_L g648 ( 
.A(n_647),
.Y(n_648)
);

INVxp67_ASAP7_75t_L g649 ( 
.A(n_646),
.Y(n_649)
);

INVx1_ASAP7_75t_L g650 ( 
.A(n_648),
.Y(n_650)
);

NOR2xp33_ASAP7_75t_L g651 ( 
.A(n_650),
.B(n_649),
.Y(n_651)
);

OAI211xp5_ASAP7_75t_L g652 ( 
.A1(n_651),
.A2(n_645),
.B(n_642),
.C(n_618),
.Y(n_652)
);

AOI211xp5_ASAP7_75t_L g653 ( 
.A1(n_652),
.A2(n_641),
.B(n_613),
.C(n_602),
.Y(n_653)
);

NAND2xp5_ASAP7_75t_SL g654 ( 
.A(n_653),
.B(n_597),
.Y(n_654)
);

XNOR2xp5_ASAP7_75t_L g655 ( 
.A(n_654),
.B(n_603),
.Y(n_655)
);

CKINVDCx5p33_ASAP7_75t_R g656 ( 
.A(n_655),
.Y(n_656)
);

INVxp67_ASAP7_75t_L g657 ( 
.A(n_656),
.Y(n_657)
);

OAI211xp5_ASAP7_75t_L g658 ( 
.A1(n_657),
.A2(n_592),
.B(n_91),
.C(n_92),
.Y(n_658)
);

NOR2xp33_ASAP7_75t_SL g659 ( 
.A(n_658),
.B(n_90),
.Y(n_659)
);

INVx1_ASAP7_75t_L g660 ( 
.A(n_659),
.Y(n_660)
);

NOR3xp33_ASAP7_75t_SL g661 ( 
.A(n_659),
.B(n_94),
.C(n_106),
.Y(n_661)
);

AOI22xp33_ASAP7_75t_L g662 ( 
.A1(n_660),
.A2(n_594),
.B1(n_584),
.B2(n_615),
.Y(n_662)
);

AOI22xp33_ASAP7_75t_R g663 ( 
.A1(n_661),
.A2(n_109),
.B1(n_110),
.B2(n_113),
.Y(n_663)
);

AOI22xp5_ASAP7_75t_L g664 ( 
.A1(n_662),
.A2(n_114),
.B1(n_115),
.B2(n_116),
.Y(n_664)
);

AOI22xp33_ASAP7_75t_L g665 ( 
.A1(n_663),
.A2(n_117),
.B1(n_120),
.B2(n_122),
.Y(n_665)
);

OAI221xp5_ASAP7_75t_L g666 ( 
.A1(n_665),
.A2(n_126),
.B1(n_128),
.B2(n_129),
.C(n_130),
.Y(n_666)
);

AOI211xp5_ASAP7_75t_L g667 ( 
.A1(n_666),
.A2(n_664),
.B(n_132),
.C(n_615),
.Y(n_667)
);


endmodule