module real_aes_2200_n_101 (n_17, n_28, n_76, n_56, n_34, n_98, n_90, n_82, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_784, n_10, n_83, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_91, n_100, n_43, n_96, n_54, n_35, n_42, n_99, n_15, n_9, n_23, n_72, n_95, n_44, n_7, n_4, n_80, n_6, n_12, n_68, n_79, n_69, n_46, n_59, n_25, n_73, n_77, n_81, n_48, n_37, n_97, n_70, n_50, n_89, n_26, n_86, n_93, n_13, n_24, n_2, n_55, n_62, n_84, n_67, n_92, n_33, n_88, n_14, n_11, n_85, n_16, n_94, n_39, n_5, n_45, n_60, n_38, n_87, n_0, n_78, n_63, n_1, n_53, n_36, n_101);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_98;
input n_90;
input n_82;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_784;
input n_10;
input n_83;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_91;
input n_100;
input n_43;
input n_96;
input n_54;
input n_35;
input n_42;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_95;
input n_44;
input n_7;
input n_4;
input n_80;
input n_6;
input n_12;
input n_68;
input n_79;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_81;
input n_48;
input n_37;
input n_97;
input n_70;
input n_50;
input n_89;
input n_26;
input n_86;
input n_93;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_84;
input n_67;
input n_92;
input n_33;
input n_88;
input n_14;
input n_11;
input n_85;
input n_16;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_87;
input n_0;
input n_78;
input n_63;
input n_1;
input n_53;
input n_36;
output n_101;
wire n_480;
wire n_113;
wire n_476;
wire n_758;
wire n_599;
wire n_187;
wire n_436;
wire n_684;
wire n_257;
wire n_390;
wire n_185;
wire n_285;
wire n_624;
wire n_618;
wire n_778;
wire n_522;
wire n_485;
wire n_222;
wire n_750;
wire n_631;
wire n_503;
wire n_287;
wire n_357;
wire n_635;
wire n_386;
wire n_673;
wire n_518;
wire n_254;
wire n_207;
wire n_665;
wire n_667;
wire n_577;
wire n_580;
wire n_469;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_759;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_718;
wire n_318;
wire n_355;
wire n_239;
wire n_669;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_761;
wire n_742;
wire n_112;
wire n_319;
wire n_421;
wire n_364;
wire n_555;
wire n_329;
wire n_766;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_242;
wire n_169;
wire n_376;
wire n_571;
wire n_549;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_752;
wire n_448;
wire n_556;
wire n_341;
wire n_545;
wire n_593;
wire n_232;
wire n_460;
wire n_773;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_537;
wire n_320;
wire n_551;
wire n_666;
wire n_560;
wire n_260;
wire n_660;
wire n_594;
wire n_186;
wire n_767;
wire n_138;
wire n_696;
wire n_704;
wire n_379;
wire n_374;
wire n_453;
wire n_647;
wire n_235;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_775;
wire n_161;
wire n_763;
wire n_189;
wire n_271;
wire n_489;
wire n_427;
wire n_548;
wire n_678;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_564;
wire n_519;
wire n_638;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_512;
wire n_395;
wire n_332;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_116;
wire n_625;
wire n_289;
wire n_462;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_716;
wire n_213;
wire n_478;
wire n_356;
wire n_584;
wire n_408;
wire n_553;
wire n_184;
wire n_372;
wire n_528;
wire n_578;
wire n_202;
wire n_495;
wire n_370;
wire n_384;
wire n_744;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_467;
wire n_327;
wire n_774;
wire n_106;
wire n_466;
wire n_559;
wire n_636;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_726;
wire n_517;
wire n_683;
wire n_780;
wire n_174;
wire n_570;
wire n_675;
wire n_530;
wire n_104;
wire n_535;
wire n_732;
wire n_211;
wire n_281;
wire n_496;
wire n_693;
wire n_173;
wire n_468;
wire n_234;
wire n_746;
wire n_284;
wire n_153;
wire n_316;
wire n_532;
wire n_656;
wire n_755;
wire n_178;
wire n_409;
wire n_748;
wire n_781;
wire n_523;
wire n_298;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_297;
wire n_383;
wire n_529;
wire n_119;
wire n_504;
wire n_310;
wire n_455;
wire n_725;
wire n_164;
wire n_671;
wire n_231;
wire n_102;
wire n_547;
wire n_659;
wire n_682;
wire n_634;
wire n_454;
wire n_122;
wire n_782;
wire n_443;
wire n_565;
wire n_760;
wire n_608;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_267;
wire n_218;
wire n_737;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_770;
wire n_745;
wire n_722;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_331;
wire n_449;
wire n_182;
wire n_363;
wire n_417;
wire n_607;
wire n_754;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_142;
wire n_561;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_655;
wire n_654;
wire n_502;
wire n_505;
wire n_769;
wire n_434;
wire n_527;
wire n_600;
wire n_731;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_602;
wire n_402;
wire n_552;
wire n_617;
wire n_733;
wire n_171;
wire n_658;
wire n_676;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_146;
wire n_432;
wire n_226;
wire n_255;
wire n_286;
wire n_416;
wire n_410;
wire n_120;
wire n_751;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_695;
wire n_685;
wire n_165;
wire n_361;
wire n_632;
wire n_246;
wire n_176;
wire n_768;
wire n_412;
wire n_163;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_777;
wire n_488;
wire n_501;
wire n_251;
wire n_642;
wire n_613;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_702;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_734;
wire n_110;
wire n_392;
wire n_562;
wire n_150;
wire n_147;
wire n_288;
wire n_404;
wire n_598;
wire n_713;
wire n_735;
wire n_728;
wire n_756;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_569;
wire n_563;
wire n_188;
wire n_269;
wire n_430;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_193;
wire n_397;
wire n_293;
wire n_162;
wire n_749;
wire n_385;
wire n_275;
wire n_214;
wire n_358;
wire n_649;
wire n_663;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_707;
wire n_622;
wire n_470;
wire n_133;
wire n_494;
wire n_711;
wire n_377;
wire n_273;
wire n_723;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_265;
wire n_354;
wire n_720;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_730;
wire n_643;
wire n_747;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_779;
wire n_148;
wire n_481;
wire n_498;
wire n_765;
wire n_691;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_233;
wire n_487;
wire n_290;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_155;
wire n_243;
wire n_692;
wire n_544;
wire n_268;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_738;
wire n_701;
wire n_309;
wire n_344;
wire n_229;
wire n_107;
wire n_482;
wire n_520;
wire n_633;
wire n_679;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_262;
wire n_630;
wire n_689;
wire n_715;
wire n_134;
wire n_349;
wire n_336;
wire n_420;
wire n_612;
wire n_195;
wire n_438;
wire n_764;
wire n_300;
wire n_252;
wire n_283;
wire n_314;
wire n_741;
wire n_753;
wire n_249;
wire n_623;
wire n_446;
wire n_721;
wire n_221;
wire n_681;
wire n_156;
wire n_359;
wire n_456;
wire n_717;
wire n_312;
wire n_183;
wire n_266;
wire n_712;
wire n_205;
wire n_433;
wire n_516;
wire n_177;
wire n_335;
wire n_313;
wire n_627;
wire n_739;
wire n_521;
wire n_140;
wire n_418;
wire n_422;
wire n_771;
wire n_219;
wire n_524;
wire n_705;
wire n_180;
wire n_212;
wire n_210;
wire n_575;
wire n_325;
wire n_762;
wire n_479;
wire n_338;
wire n_442;
wire n_698;
wire n_371;
wire n_740;
wire n_166;
wire n_103;
wire n_541;
wire n_224;
wire n_151;
wire n_546;
wire n_587;
wire n_639;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_724;
wire n_440;
wire n_525;
wire n_644;
wire n_674;
wire n_152;
wire n_198;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_414;
wire n_757;
wire n_123;
wire n_279;
wire n_686;
wire n_776;
wire n_543;
wire n_497;
wire n_514;
wire n_507;
wire n_270;
wire n_614;
wire n_305;
wire n_586;
wire n_772;
wire n_450;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_465;
wire n_473;
wire n_719;
wire n_566;
wire n_474;
wire n_170;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_168;
wire n_175;
wire n_241;
wire n_687;
wire n_729;
wire n_646;
wire n_650;
wire n_710;
wire n_105;
wire n_743;
wire n_294;
wire n_393;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_307;
wire n_500;
wire n_601;
wire n_661;
wire n_463;
wire n_396;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_143;
wire n_192;
wire n_475;
wire n_554;
wire n_264;
wire n_237;
wire n_668;
NAND2xp5_ASAP7_75t_L g229 ( .A(n_0), .B(n_166), .Y(n_229) );
NAND2xp5_ASAP7_75t_L g109 ( .A(n_1), .B(n_110), .Y(n_109) );
NAND2xp5_ASAP7_75t_L g536 ( .A(n_2), .B(n_142), .Y(n_536) );
NAND2xp5_ASAP7_75t_L g479 ( .A(n_3), .B(n_164), .Y(n_479) );
INVx1_ASAP7_75t_L g138 ( .A(n_4), .Y(n_138) );
NAND2xp5_ASAP7_75t_L g187 ( .A(n_5), .B(n_142), .Y(n_187) );
NAND2xp33_ASAP7_75t_SL g249 ( .A(n_6), .B(n_148), .Y(n_249) );
INVx1_ASAP7_75t_L g241 ( .A(n_7), .Y(n_241) );
AOI22xp5_ASAP7_75t_L g776 ( .A1(n_8), .A2(n_57), .B1(n_777), .B2(n_778), .Y(n_776) );
CKINVDCx20_ASAP7_75t_R g777 ( .A(n_8), .Y(n_777) );
CKINVDCx16_ASAP7_75t_R g110 ( .A(n_9), .Y(n_110) );
AND2x2_ASAP7_75t_L g185 ( .A(n_10), .B(n_171), .Y(n_185) );
AND2x2_ASAP7_75t_L g472 ( .A(n_11), .B(n_247), .Y(n_472) );
AND2x2_ASAP7_75t_L g481 ( .A(n_12), .B(n_128), .Y(n_481) );
INVx2_ASAP7_75t_L g130 ( .A(n_13), .Y(n_130) );
NAND2xp5_ASAP7_75t_L g506 ( .A(n_14), .B(n_164), .Y(n_506) );
CKINVDCx16_ASAP7_75t_R g111 ( .A(n_15), .Y(n_111) );
AOI221x1_ASAP7_75t_L g244 ( .A1(n_16), .A2(n_150), .B1(n_245), .B2(n_247), .C(n_248), .Y(n_244) );
NAND2xp5_ASAP7_75t_SL g209 ( .A(n_17), .B(n_142), .Y(n_209) );
OAI22xp5_ASAP7_75t_SL g746 ( .A1(n_18), .A2(n_69), .B1(n_747), .B2(n_748), .Y(n_746) );
CKINVDCx20_ASAP7_75t_R g748 ( .A(n_18), .Y(n_748) );
NAND2xp5_ASAP7_75t_SL g521 ( .A(n_19), .B(n_142), .Y(n_521) );
INVx1_ASAP7_75t_L g107 ( .A(n_20), .Y(n_107) );
AOI22xp33_ASAP7_75t_L g460 ( .A1(n_21), .A2(n_90), .B1(n_133), .B2(n_142), .Y(n_460) );
AOI21xp5_ASAP7_75t_L g188 ( .A1(n_22), .A2(n_150), .B(n_189), .Y(n_188) );
AOI221xp5_ASAP7_75t_SL g218 ( .A1(n_23), .A2(n_38), .B1(n_142), .B2(n_150), .C(n_219), .Y(n_218) );
NAND2xp5_ASAP7_75t_L g190 ( .A(n_24), .B(n_166), .Y(n_190) );
OA21x2_ASAP7_75t_L g129 ( .A1(n_25), .A2(n_89), .B(n_130), .Y(n_129) );
OR2x2_ASAP7_75t_L g172 ( .A(n_25), .B(n_89), .Y(n_172) );
NAND2xp5_ASAP7_75t_L g213 ( .A(n_26), .B(n_164), .Y(n_213) );
INVxp67_ASAP7_75t_L g243 ( .A(n_27), .Y(n_243) );
AND2x2_ASAP7_75t_L g182 ( .A(n_28), .B(n_170), .Y(n_182) );
CKINVDCx20_ASAP7_75t_R g780 ( .A(n_29), .Y(n_780) );
AOI21xp5_ASAP7_75t_L g227 ( .A1(n_30), .A2(n_150), .B(n_228), .Y(n_227) );
AO21x2_ASAP7_75t_L g501 ( .A1(n_31), .A2(n_247), .B(n_502), .Y(n_501) );
NAND2xp5_ASAP7_75t_L g220 ( .A(n_32), .B(n_164), .Y(n_220) );
AOI21xp5_ASAP7_75t_L g476 ( .A1(n_33), .A2(n_150), .B(n_477), .Y(n_476) );
CKINVDCx20_ASAP7_75t_R g759 ( .A(n_34), .Y(n_759) );
NAND2xp5_ASAP7_75t_L g535 ( .A(n_35), .B(n_164), .Y(n_535) );
AND2x2_ASAP7_75t_L g140 ( .A(n_36), .B(n_141), .Y(n_140) );
AND2x2_ASAP7_75t_L g148 ( .A(n_36), .B(n_138), .Y(n_148) );
INVx1_ASAP7_75t_L g154 ( .A(n_36), .Y(n_154) );
NOR3xp33_ASAP7_75t_L g108 ( .A(n_37), .B(n_109), .C(n_111), .Y(n_108) );
OR2x6_ASAP7_75t_L g118 ( .A(n_37), .B(n_119), .Y(n_118) );
NAND2xp5_ASAP7_75t_L g480 ( .A(n_39), .B(n_142), .Y(n_480) );
AOI22xp5_ASAP7_75t_L g149 ( .A1(n_40), .A2(n_82), .B1(n_150), .B2(n_152), .Y(n_149) );
NAND2xp5_ASAP7_75t_L g516 ( .A(n_41), .B(n_164), .Y(n_516) );
NAND2xp5_ASAP7_75t_L g488 ( .A(n_42), .B(n_142), .Y(n_488) );
NAND2xp5_ASAP7_75t_L g180 ( .A(n_43), .B(n_166), .Y(n_180) );
AOI21xp5_ASAP7_75t_L g467 ( .A1(n_44), .A2(n_150), .B(n_468), .Y(n_467) );
AND2x2_ASAP7_75t_L g232 ( .A(n_45), .B(n_170), .Y(n_232) );
NAND2xp5_ASAP7_75t_L g492 ( .A(n_46), .B(n_166), .Y(n_492) );
NAND2xp5_ASAP7_75t_L g222 ( .A(n_47), .B(n_170), .Y(n_222) );
NAND2xp5_ASAP7_75t_SL g503 ( .A(n_48), .B(n_142), .Y(n_503) );
INVx1_ASAP7_75t_L g136 ( .A(n_49), .Y(n_136) );
INVx1_ASAP7_75t_L g145 ( .A(n_49), .Y(n_145) );
NAND2xp5_ASAP7_75t_L g470 ( .A(n_50), .B(n_164), .Y(n_470) );
AND2x2_ASAP7_75t_L g511 ( .A(n_51), .B(n_170), .Y(n_511) );
NAND2xp5_ASAP7_75t_SL g181 ( .A(n_52), .B(n_142), .Y(n_181) );
NAND2xp5_ASAP7_75t_L g469 ( .A(n_53), .B(n_166), .Y(n_469) );
NAND2xp5_ASAP7_75t_L g534 ( .A(n_54), .B(n_166), .Y(n_534) );
AND2x2_ASAP7_75t_L g173 ( .A(n_55), .B(n_170), .Y(n_173) );
NAND2xp5_ASAP7_75t_SL g471 ( .A(n_56), .B(n_142), .Y(n_471) );
CKINVDCx20_ASAP7_75t_R g778 ( .A(n_57), .Y(n_778) );
NAND2xp5_ASAP7_75t_L g230 ( .A(n_58), .B(n_164), .Y(n_230) );
NAND2xp5_ASAP7_75t_SL g513 ( .A(n_59), .B(n_142), .Y(n_513) );
AOI21xp5_ASAP7_75t_L g532 ( .A1(n_60), .A2(n_150), .B(n_533), .Y(n_532) );
NAND2xp5_ASAP7_75t_L g165 ( .A(n_61), .B(n_166), .Y(n_165) );
AND2x2_ASAP7_75t_SL g214 ( .A(n_62), .B(n_171), .Y(n_214) );
AND2x2_ASAP7_75t_L g527 ( .A(n_63), .B(n_171), .Y(n_527) );
AOI21xp5_ASAP7_75t_L g177 ( .A1(n_64), .A2(n_150), .B(n_178), .Y(n_177) );
NAND2xp5_ASAP7_75t_L g191 ( .A(n_65), .B(n_164), .Y(n_191) );
AND2x2_ASAP7_75t_SL g157 ( .A(n_66), .B(n_128), .Y(n_157) );
NAND2xp5_ASAP7_75t_L g517 ( .A(n_67), .B(n_166), .Y(n_517) );
NAND2xp5_ASAP7_75t_L g507 ( .A(n_68), .B(n_166), .Y(n_507) );
CKINVDCx20_ASAP7_75t_R g747 ( .A(n_69), .Y(n_747) );
CKINVDCx20_ASAP7_75t_R g753 ( .A(n_70), .Y(n_753) );
AOI22xp5_ASAP7_75t_L g461 ( .A1(n_71), .A2(n_92), .B1(n_150), .B2(n_152), .Y(n_461) );
NAND2xp5_ASAP7_75t_L g524 ( .A(n_72), .B(n_164), .Y(n_524) );
INVx1_ASAP7_75t_L g141 ( .A(n_73), .Y(n_141) );
INVx1_ASAP7_75t_L g147 ( .A(n_73), .Y(n_147) );
NAND2xp5_ASAP7_75t_L g478 ( .A(n_74), .B(n_166), .Y(n_478) );
AOI21xp5_ASAP7_75t_L g514 ( .A1(n_75), .A2(n_150), .B(n_515), .Y(n_514) );
AOI21xp5_ASAP7_75t_L g489 ( .A1(n_76), .A2(n_150), .B(n_490), .Y(n_489) );
AOI21xp5_ASAP7_75t_L g504 ( .A1(n_77), .A2(n_150), .B(n_505), .Y(n_504) );
AND2x2_ASAP7_75t_L g537 ( .A(n_78), .B(n_171), .Y(n_537) );
NAND2xp5_ASAP7_75t_SL g458 ( .A(n_79), .B(n_170), .Y(n_458) );
AOI22xp5_ASAP7_75t_L g132 ( .A1(n_80), .A2(n_84), .B1(n_133), .B2(n_142), .Y(n_132) );
NAND2xp5_ASAP7_75t_SL g168 ( .A(n_81), .B(n_142), .Y(n_168) );
INVx1_ASAP7_75t_L g106 ( .A(n_83), .Y(n_106) );
NAND2xp5_ASAP7_75t_L g212 ( .A(n_85), .B(n_166), .Y(n_212) );
NAND2xp5_ASAP7_75t_L g221 ( .A(n_86), .B(n_166), .Y(n_221) );
AND2x2_ASAP7_75t_L g493 ( .A(n_87), .B(n_128), .Y(n_493) );
AOI21xp5_ASAP7_75t_L g161 ( .A1(n_88), .A2(n_150), .B(n_162), .Y(n_161) );
NAND2xp5_ASAP7_75t_L g163 ( .A(n_91), .B(n_164), .Y(n_163) );
AOI21xp5_ASAP7_75t_L g522 ( .A1(n_93), .A2(n_150), .B(n_523), .Y(n_522) );
NAND2xp5_ASAP7_75t_L g491 ( .A(n_94), .B(n_164), .Y(n_491) );
NAND2xp5_ASAP7_75t_L g231 ( .A(n_95), .B(n_142), .Y(n_231) );
INVxp67_ASAP7_75t_L g246 ( .A(n_96), .Y(n_246) );
NAND2xp5_ASAP7_75t_L g179 ( .A(n_97), .B(n_164), .Y(n_179) );
AOI21xp5_ASAP7_75t_L g210 ( .A1(n_98), .A2(n_150), .B(n_211), .Y(n_210) );
BUFx2_ASAP7_75t_L g526 ( .A(n_99), .Y(n_526) );
BUFx2_ASAP7_75t_L g768 ( .A(n_100), .Y(n_768) );
INVx1_ASAP7_75t_SL g771 ( .A(n_100), .Y(n_771) );
AOI21xp5_ASAP7_75t_L g101 ( .A1(n_102), .A2(n_112), .B(n_779), .Y(n_101) );
INVx2_ASAP7_75t_R g102 ( .A(n_103), .Y(n_102) );
CKINVDCx5p33_ASAP7_75t_R g782 ( .A(n_103), .Y(n_782) );
INVx3_ASAP7_75t_SL g103 ( .A(n_104), .Y(n_103) );
AND2x2_ASAP7_75t_SL g104 ( .A(n_105), .B(n_108), .Y(n_104) );
NOR2xp33_ASAP7_75t_L g105 ( .A(n_106), .B(n_107), .Y(n_105) );
NAND2xp5_ASAP7_75t_L g119 ( .A(n_106), .B(n_107), .Y(n_119) );
AND2x6_ASAP7_75t_SL g117 ( .A(n_111), .B(n_118), .Y(n_117) );
OR2x6_ASAP7_75t_SL g744 ( .A(n_111), .B(n_745), .Y(n_744) );
OR2x2_ASAP7_75t_L g756 ( .A(n_111), .B(n_118), .Y(n_756) );
NAND2xp5_ASAP7_75t_L g764 ( .A(n_111), .B(n_745), .Y(n_764) );
OR2x2_ASAP7_75t_L g112 ( .A(n_113), .B(n_769), .Y(n_112) );
AOI21xp5_ASAP7_75t_L g113 ( .A1(n_114), .A2(n_757), .B(n_765), .Y(n_113) );
AOI221xp5_ASAP7_75t_L g114 ( .A1(n_115), .A2(n_746), .B1(n_749), .B2(n_750), .C(n_752), .Y(n_114) );
OAI22xp5_ASAP7_75t_L g115 ( .A1(n_116), .A2(n_120), .B1(n_449), .B2(n_742), .Y(n_115) );
INVx3_ASAP7_75t_SL g751 ( .A(n_116), .Y(n_751) );
CKINVDCx5p33_ASAP7_75t_R g116 ( .A(n_117), .Y(n_116) );
CKINVDCx5p33_ASAP7_75t_R g745 ( .A(n_118), .Y(n_745) );
AO22x1_ASAP7_75t_L g750 ( .A1(n_120), .A2(n_449), .B1(n_743), .B2(n_751), .Y(n_750) );
XNOR2x1_ASAP7_75t_L g775 ( .A(n_120), .B(n_776), .Y(n_775) );
AND3x4_ASAP7_75t_L g120 ( .A(n_121), .B(n_320), .C(n_394), .Y(n_120) );
NOR3xp33_ASAP7_75t_L g121 ( .A(n_122), .B(n_262), .C(n_293), .Y(n_121) );
A2O1A1Ixp33_ASAP7_75t_L g122 ( .A1(n_123), .A2(n_195), .B(n_204), .C(n_233), .Y(n_122) );
AOI21x1_ASAP7_75t_SL g123 ( .A1(n_124), .A2(n_174), .B(n_193), .Y(n_123) );
AOI22xp33_ASAP7_75t_L g295 ( .A1(n_124), .A2(n_296), .B1(n_302), .B2(n_305), .Y(n_295) );
AND2x2_ASAP7_75t_L g429 ( .A(n_124), .B(n_197), .Y(n_429) );
AND2x2_ASAP7_75t_L g124 ( .A(n_125), .B(n_158), .Y(n_124) );
BUFx2_ASAP7_75t_L g200 ( .A(n_125), .Y(n_200) );
AND2x2_ASAP7_75t_L g288 ( .A(n_125), .B(n_159), .Y(n_288) );
AND2x2_ASAP7_75t_L g359 ( .A(n_125), .B(n_203), .Y(n_359) );
INVx2_ASAP7_75t_L g125 ( .A(n_126), .Y(n_125) );
BUFx6f_ASAP7_75t_L g253 ( .A(n_126), .Y(n_253) );
AOI21x1_ASAP7_75t_L g126 ( .A1(n_127), .A2(n_131), .B(n_157), .Y(n_126) );
INVx2_ASAP7_75t_SL g127 ( .A(n_128), .Y(n_127) );
AOI21xp5_ASAP7_75t_L g208 ( .A1(n_128), .A2(n_209), .B(n_210), .Y(n_208) );
AOI21xp5_ASAP7_75t_L g520 ( .A1(n_128), .A2(n_521), .B(n_522), .Y(n_520) );
BUFx4f_ASAP7_75t_L g128 ( .A(n_129), .Y(n_128) );
INVx3_ASAP7_75t_L g225 ( .A(n_129), .Y(n_225) );
AND2x2_ASAP7_75t_SL g171 ( .A(n_130), .B(n_172), .Y(n_171) );
AND2x4_ASAP7_75t_L g192 ( .A(n_130), .B(n_172), .Y(n_192) );
NAND2xp5_ASAP7_75t_L g131 ( .A(n_132), .B(n_149), .Y(n_131) );
AOI22xp5_ASAP7_75t_L g239 ( .A1(n_133), .A2(n_152), .B1(n_240), .B2(n_242), .Y(n_239) );
AND2x4_ASAP7_75t_L g133 ( .A(n_134), .B(n_139), .Y(n_133) );
AND2x2_ASAP7_75t_L g134 ( .A(n_135), .B(n_137), .Y(n_134) );
INVx2_ASAP7_75t_L g135 ( .A(n_136), .Y(n_135) );
AND2x2_ASAP7_75t_L g151 ( .A(n_136), .B(n_138), .Y(n_151) );
AND2x4_ASAP7_75t_L g164 ( .A(n_136), .B(n_146), .Y(n_164) );
HB1xp67_ASAP7_75t_L g137 ( .A(n_138), .Y(n_137) );
BUFx3_ASAP7_75t_L g139 ( .A(n_140), .Y(n_139) );
AND2x6_ASAP7_75t_L g150 ( .A(n_140), .B(n_151), .Y(n_150) );
INVx2_ASAP7_75t_L g156 ( .A(n_141), .Y(n_156) );
AND2x6_ASAP7_75t_L g166 ( .A(n_141), .B(n_144), .Y(n_166) );
AND2x4_ASAP7_75t_L g142 ( .A(n_143), .B(n_148), .Y(n_142) );
INVx1_ASAP7_75t_L g250 ( .A(n_143), .Y(n_250) );
AND2x4_ASAP7_75t_L g143 ( .A(n_144), .B(n_146), .Y(n_143) );
INVx2_ASAP7_75t_L g144 ( .A(n_145), .Y(n_144) );
INVx2_ASAP7_75t_L g146 ( .A(n_147), .Y(n_146) );
INVx5_ASAP7_75t_L g167 ( .A(n_148), .Y(n_167) );
AND2x4_ASAP7_75t_L g152 ( .A(n_151), .B(n_153), .Y(n_152) );
NOR2x1p5_ASAP7_75t_L g153 ( .A(n_154), .B(n_155), .Y(n_153) );
INVx3_ASAP7_75t_L g155 ( .A(n_156), .Y(n_155) );
AND2x4_ASAP7_75t_L g252 ( .A(n_158), .B(n_253), .Y(n_252) );
INVx2_ASAP7_75t_L g158 ( .A(n_159), .Y(n_158) );
AND2x2_ASAP7_75t_L g194 ( .A(n_159), .B(n_184), .Y(n_194) );
OR2x2_ASAP7_75t_L g202 ( .A(n_159), .B(n_203), .Y(n_202) );
AND2x4_ASAP7_75t_L g257 ( .A(n_159), .B(n_258), .Y(n_257) );
INVx1_ASAP7_75t_L g304 ( .A(n_159), .Y(n_304) );
NAND2xp5_ASAP7_75t_L g312 ( .A(n_159), .B(n_203), .Y(n_312) );
AND2x2_ASAP7_75t_L g349 ( .A(n_159), .B(n_253), .Y(n_349) );
HB1xp67_ASAP7_75t_L g358 ( .A(n_159), .Y(n_358) );
NAND2xp5_ASAP7_75t_L g390 ( .A(n_159), .B(n_183), .Y(n_390) );
AO21x2_ASAP7_75t_L g159 ( .A1(n_160), .A2(n_169), .B(n_173), .Y(n_159) );
NAND2xp5_ASAP7_75t_L g160 ( .A(n_161), .B(n_168), .Y(n_160) );
AOI21xp5_ASAP7_75t_L g162 ( .A1(n_163), .A2(n_165), .B(n_167), .Y(n_162) );
NAND2xp5_ASAP7_75t_L g525 ( .A(n_166), .B(n_526), .Y(n_525) );
AOI21xp5_ASAP7_75t_L g178 ( .A1(n_167), .A2(n_179), .B(n_180), .Y(n_178) );
AOI21xp5_ASAP7_75t_L g189 ( .A1(n_167), .A2(n_190), .B(n_191), .Y(n_189) );
AOI21xp5_ASAP7_75t_L g211 ( .A1(n_167), .A2(n_212), .B(n_213), .Y(n_211) );
AOI21xp5_ASAP7_75t_L g219 ( .A1(n_167), .A2(n_220), .B(n_221), .Y(n_219) );
AOI21xp5_ASAP7_75t_L g228 ( .A1(n_167), .A2(n_229), .B(n_230), .Y(n_228) );
AOI21xp5_ASAP7_75t_L g468 ( .A1(n_167), .A2(n_469), .B(n_470), .Y(n_468) );
AOI21xp5_ASAP7_75t_L g477 ( .A1(n_167), .A2(n_478), .B(n_479), .Y(n_477) );
AOI21xp5_ASAP7_75t_L g490 ( .A1(n_167), .A2(n_491), .B(n_492), .Y(n_490) );
AOI21xp5_ASAP7_75t_L g505 ( .A1(n_167), .A2(n_506), .B(n_507), .Y(n_505) );
AOI21xp5_ASAP7_75t_L g515 ( .A1(n_167), .A2(n_516), .B(n_517), .Y(n_515) );
AOI21xp5_ASAP7_75t_L g523 ( .A1(n_167), .A2(n_524), .B(n_525), .Y(n_523) );
AOI21xp5_ASAP7_75t_L g533 ( .A1(n_167), .A2(n_534), .B(n_535), .Y(n_533) );
AO21x2_ASAP7_75t_L g175 ( .A1(n_169), .A2(n_176), .B(n_182), .Y(n_175) );
AO21x2_ASAP7_75t_L g203 ( .A1(n_169), .A2(n_176), .B(n_182), .Y(n_203) );
AOI21x1_ASAP7_75t_L g474 ( .A1(n_169), .A2(n_475), .B(n_481), .Y(n_474) );
CKINVDCx5p33_ASAP7_75t_R g169 ( .A(n_170), .Y(n_169) );
OA21x2_ASAP7_75t_L g217 ( .A1(n_170), .A2(n_218), .B(n_222), .Y(n_217) );
AO21x2_ASAP7_75t_L g459 ( .A1(n_170), .A2(n_460), .B(n_461), .Y(n_459) );
AOI21xp5_ASAP7_75t_L g487 ( .A1(n_170), .A2(n_488), .B(n_489), .Y(n_487) );
BUFx6f_ASAP7_75t_L g170 ( .A(n_171), .Y(n_170) );
INVx2_ASAP7_75t_L g291 ( .A(n_174), .Y(n_291) );
NAND2xp5_ASAP7_75t_L g347 ( .A(n_174), .B(n_252), .Y(n_347) );
HB1xp67_ASAP7_75t_L g448 ( .A(n_174), .Y(n_448) );
AND2x4_ASAP7_75t_L g174 ( .A(n_175), .B(n_183), .Y(n_174) );
AND2x2_ASAP7_75t_L g193 ( .A(n_175), .B(n_194), .Y(n_193) );
OR2x2_ASAP7_75t_L g273 ( .A(n_175), .B(n_184), .Y(n_273) );
NAND2xp5_ASAP7_75t_L g387 ( .A(n_175), .B(n_304), .Y(n_387) );
NAND2xp5_ASAP7_75t_L g176 ( .A(n_177), .B(n_181), .Y(n_176) );
AND2x2_ASAP7_75t_L g340 ( .A(n_183), .B(n_257), .Y(n_340) );
NAND2xp5_ASAP7_75t_L g396 ( .A(n_183), .B(n_252), .Y(n_396) );
INVx5_ASAP7_75t_L g183 ( .A(n_184), .Y(n_183) );
INVx2_ASAP7_75t_L g198 ( .A(n_184), .Y(n_198) );
AND2x2_ASAP7_75t_L g267 ( .A(n_184), .B(n_258), .Y(n_267) );
HB1xp67_ASAP7_75t_L g287 ( .A(n_184), .Y(n_287) );
AND2x4_ASAP7_75t_L g294 ( .A(n_184), .B(n_203), .Y(n_294) );
AND2x2_ASAP7_75t_SL g441 ( .A(n_184), .B(n_253), .Y(n_441) );
OR2x6_ASAP7_75t_L g184 ( .A(n_185), .B(n_186), .Y(n_184) );
AOI21xp5_ASAP7_75t_L g186 ( .A1(n_187), .A2(n_188), .B(n_192), .Y(n_186) );
NOR2xp33_ASAP7_75t_L g240 ( .A(n_192), .B(n_241), .Y(n_240) );
NOR2xp33_ASAP7_75t_L g242 ( .A(n_192), .B(n_243), .Y(n_242) );
NOR2xp33_ASAP7_75t_L g245 ( .A(n_192), .B(n_246), .Y(n_245) );
NOR3xp33_ASAP7_75t_L g248 ( .A(n_192), .B(n_249), .C(n_250), .Y(n_248) );
AOI21xp5_ASAP7_75t_L g502 ( .A1(n_192), .A2(n_503), .B(n_504), .Y(n_502) );
AOI21xp5_ASAP7_75t_L g512 ( .A1(n_192), .A2(n_513), .B(n_514), .Y(n_512) );
INVx1_ASAP7_75t_L g420 ( .A(n_193), .Y(n_420) );
INVx1_ASAP7_75t_L g362 ( .A(n_194), .Y(n_362) );
INVx1_ASAP7_75t_L g195 ( .A(n_196), .Y(n_195) );
AND2x2_ASAP7_75t_L g196 ( .A(n_197), .B(n_199), .Y(n_196) );
INVx2_ASAP7_75t_L g197 ( .A(n_198), .Y(n_197) );
OR2x2_ASAP7_75t_L g284 ( .A(n_198), .B(n_202), .Y(n_284) );
NOR2xp33_ASAP7_75t_L g377 ( .A(n_198), .B(n_253), .Y(n_377) );
AND2x2_ASAP7_75t_L g379 ( .A(n_198), .B(n_201), .Y(n_379) );
AOI32xp33_ASAP7_75t_L g445 ( .A1(n_198), .A2(n_261), .A3(n_416), .B1(n_446), .B2(n_448), .Y(n_445) );
AND2x2_ASAP7_75t_L g199 ( .A(n_200), .B(n_201), .Y(n_199) );
AND2x2_ASAP7_75t_L g271 ( .A(n_200), .B(n_272), .Y(n_271) );
OR2x2_ASAP7_75t_L g389 ( .A(n_200), .B(n_390), .Y(n_389) );
OR2x2_ASAP7_75t_L g412 ( .A(n_200), .B(n_273), .Y(n_412) );
AND2x2_ASAP7_75t_L g439 ( .A(n_200), .B(n_340), .Y(n_439) );
AND2x2_ASAP7_75t_L g365 ( .A(n_201), .B(n_253), .Y(n_365) );
AND2x2_ASAP7_75t_L g440 ( .A(n_201), .B(n_441), .Y(n_440) );
INVx2_ASAP7_75t_L g201 ( .A(n_202), .Y(n_201) );
INVx2_ASAP7_75t_L g258 ( .A(n_203), .Y(n_258) );
INVx1_ASAP7_75t_L g204 ( .A(n_205), .Y(n_204) );
AND2x2_ASAP7_75t_L g205 ( .A(n_206), .B(n_215), .Y(n_205) );
NOR2x1p5_ASAP7_75t_L g298 ( .A(n_206), .B(n_299), .Y(n_298) );
INVx1_ASAP7_75t_L g316 ( .A(n_206), .Y(n_316) );
OR2x2_ASAP7_75t_L g344 ( .A(n_206), .B(n_345), .Y(n_344) );
INVx2_ASAP7_75t_L g206 ( .A(n_207), .Y(n_206) );
AND2x4_ASAP7_75t_SL g261 ( .A(n_207), .B(n_238), .Y(n_261) );
AND2x4_ASAP7_75t_L g277 ( .A(n_207), .B(n_278), .Y(n_277) );
OR2x2_ASAP7_75t_L g280 ( .A(n_207), .B(n_281), .Y(n_280) );
OR2x2_ASAP7_75t_L g308 ( .A(n_207), .B(n_217), .Y(n_308) );
OR2x2_ASAP7_75t_L g333 ( .A(n_207), .B(n_282), .Y(n_333) );
NAND2xp5_ASAP7_75t_L g337 ( .A(n_207), .B(n_338), .Y(n_337) );
NAND2xp5_ASAP7_75t_L g368 ( .A(n_207), .B(n_217), .Y(n_368) );
INVx2_ASAP7_75t_L g384 ( .A(n_207), .Y(n_384) );
AND2x2_ASAP7_75t_L g399 ( .A(n_207), .B(n_237), .Y(n_399) );
HB1xp67_ASAP7_75t_L g423 ( .A(n_207), .Y(n_423) );
INVx1_ASAP7_75t_L g428 ( .A(n_207), .Y(n_428) );
OR2x6_ASAP7_75t_L g207 ( .A(n_208), .B(n_214), .Y(n_207) );
AND2x2_ASAP7_75t_L g292 ( .A(n_215), .B(n_277), .Y(n_292) );
AND2x2_ASAP7_75t_L g313 ( .A(n_215), .B(n_261), .Y(n_313) );
INVx1_ASAP7_75t_L g345 ( .A(n_215), .Y(n_345) );
AND2x2_ASAP7_75t_L g215 ( .A(n_216), .B(n_223), .Y(n_215) );
INVx2_ASAP7_75t_L g216 ( .A(n_217), .Y(n_216) );
INVx1_ASAP7_75t_L g236 ( .A(n_217), .Y(n_236) );
INVx2_ASAP7_75t_L g282 ( .A(n_217), .Y(n_282) );
BUFx3_ASAP7_75t_L g299 ( .A(n_217), .Y(n_299) );
AND2x2_ASAP7_75t_L g338 ( .A(n_217), .B(n_223), .Y(n_338) );
HB1xp67_ASAP7_75t_L g436 ( .A(n_217), .Y(n_436) );
INVx2_ASAP7_75t_L g251 ( .A(n_223), .Y(n_251) );
HB1xp67_ASAP7_75t_L g260 ( .A(n_223), .Y(n_260) );
INVx1_ASAP7_75t_L g276 ( .A(n_223), .Y(n_276) );
OR2x2_ASAP7_75t_L g281 ( .A(n_223), .B(n_282), .Y(n_281) );
INVx1_ASAP7_75t_L g301 ( .A(n_223), .Y(n_301) );
NAND2xp5_ASAP7_75t_L g369 ( .A(n_223), .B(n_278), .Y(n_369) );
NAND2xp5_ASAP7_75t_L g383 ( .A(n_223), .B(n_384), .Y(n_383) );
INVx3_ASAP7_75t_L g223 ( .A(n_224), .Y(n_223) );
AOI21x1_ASAP7_75t_L g224 ( .A1(n_225), .A2(n_226), .B(n_232), .Y(n_224) );
INVx4_ASAP7_75t_L g247 ( .A(n_225), .Y(n_247) );
AO21x2_ASAP7_75t_L g465 ( .A1(n_225), .A2(n_466), .B(n_472), .Y(n_465) );
NAND2xp5_ASAP7_75t_L g226 ( .A(n_227), .B(n_231), .Y(n_226) );
AOI21xp5_ASAP7_75t_L g233 ( .A1(n_234), .A2(n_252), .B(n_254), .Y(n_233) );
AND2x2_ASAP7_75t_SL g234 ( .A(n_235), .B(n_237), .Y(n_234) );
HB1xp67_ASAP7_75t_L g444 ( .A(n_235), .Y(n_444) );
INVx1_ASAP7_75t_L g235 ( .A(n_236), .Y(n_235) );
INVxp67_ASAP7_75t_SL g270 ( .A(n_236), .Y(n_270) );
NAND2xp5_ASAP7_75t_L g318 ( .A(n_236), .B(n_276), .Y(n_318) );
HB1xp67_ASAP7_75t_L g433 ( .A(n_236), .Y(n_433) );
NAND2xp5_ASAP7_75t_L g306 ( .A(n_237), .B(n_307), .Y(n_306) );
AND2x2_ASAP7_75t_L g323 ( .A(n_237), .B(n_324), .Y(n_323) );
INVx1_ASAP7_75t_L g374 ( .A(n_237), .Y(n_374) );
AOI221xp5_ASAP7_75t_L g378 ( .A1(n_237), .A2(n_379), .B1(n_380), .B2(n_385), .C(n_388), .Y(n_378) );
NAND2xp5_ASAP7_75t_L g427 ( .A(n_237), .B(n_428), .Y(n_427) );
AND2x4_ASAP7_75t_L g237 ( .A(n_238), .B(n_251), .Y(n_237) );
INVx3_ASAP7_75t_L g278 ( .A(n_238), .Y(n_278) );
NAND2xp5_ASAP7_75t_L g382 ( .A(n_238), .B(n_282), .Y(n_382) );
AND2x2_ASAP7_75t_L g411 ( .A(n_238), .B(n_384), .Y(n_411) );
NOR2xp33_ASAP7_75t_L g442 ( .A(n_238), .B(n_443), .Y(n_442) );
AND2x4_ASAP7_75t_L g238 ( .A(n_239), .B(n_244), .Y(n_238) );
INVx3_ASAP7_75t_L g530 ( .A(n_247), .Y(n_530) );
AND2x2_ASAP7_75t_L g319 ( .A(n_252), .B(n_294), .Y(n_319) );
AOI21xp5_ASAP7_75t_L g355 ( .A1(n_252), .A2(n_272), .B(n_356), .Y(n_355) );
AND2x2_ASAP7_75t_L g256 ( .A(n_253), .B(n_257), .Y(n_256) );
INVx2_ASAP7_75t_L g265 ( .A(n_253), .Y(n_265) );
OR2x2_ASAP7_75t_L g311 ( .A(n_253), .B(n_312), .Y(n_311) );
NAND2xp5_ASAP7_75t_SL g403 ( .A(n_253), .B(n_294), .Y(n_403) );
OR2x2_ASAP7_75t_L g435 ( .A(n_253), .B(n_436), .Y(n_435) );
OR2x2_ASAP7_75t_L g447 ( .A(n_253), .B(n_353), .Y(n_447) );
INVxp67_ASAP7_75t_L g254 ( .A(n_255), .Y(n_254) );
NAND2xp5_ASAP7_75t_L g255 ( .A(n_256), .B(n_259), .Y(n_255) );
INVx2_ASAP7_75t_L g325 ( .A(n_256), .Y(n_325) );
INVx3_ASAP7_75t_SL g391 ( .A(n_257), .Y(n_391) );
INVxp67_ASAP7_75t_L g341 ( .A(n_259), .Y(n_341) );
AND2x2_ASAP7_75t_L g259 ( .A(n_260), .B(n_261), .Y(n_259) );
AOI322xp5_ASAP7_75t_L g263 ( .A1(n_261), .A2(n_264), .A3(n_268), .B1(n_271), .B2(n_274), .C1(n_279), .C2(n_283), .Y(n_263) );
INVx1_ASAP7_75t_SL g352 ( .A(n_261), .Y(n_352) );
AND2x4_ASAP7_75t_L g437 ( .A(n_261), .B(n_324), .Y(n_437) );
NAND2xp5_ASAP7_75t_L g262 ( .A(n_263), .B(n_285), .Y(n_262) );
NOR2x1_ASAP7_75t_L g264 ( .A(n_265), .B(n_266), .Y(n_264) );
OR2x2_ASAP7_75t_L g290 ( .A(n_265), .B(n_291), .Y(n_290) );
OR2x2_ASAP7_75t_L g386 ( .A(n_265), .B(n_387), .Y(n_386) );
AND2x2_ASAP7_75t_L g414 ( .A(n_265), .B(n_267), .Y(n_414) );
AOI32xp33_ASAP7_75t_L g415 ( .A1(n_265), .A2(n_266), .A3(n_416), .B1(n_418), .B2(n_421), .Y(n_415) );
OR2x2_ASAP7_75t_L g419 ( .A(n_265), .B(n_312), .Y(n_419) );
NAND3xp33_ASAP7_75t_L g375 ( .A(n_266), .B(n_291), .C(n_376), .Y(n_375) );
OAI22xp33_ASAP7_75t_SL g395 ( .A1(n_266), .A2(n_332), .B1(n_396), .B2(n_397), .Y(n_395) );
INVx2_ASAP7_75t_L g266 ( .A(n_267), .Y(n_266) );
INVxp67_ASAP7_75t_L g268 ( .A(n_269), .Y(n_268) );
AND2x2_ASAP7_75t_L g398 ( .A(n_269), .B(n_399), .Y(n_398) );
INVx1_ASAP7_75t_L g269 ( .A(n_270), .Y(n_269) );
INVx1_ASAP7_75t_SL g272 ( .A(n_273), .Y(n_272) );
NOR2xp33_ASAP7_75t_L g434 ( .A(n_273), .B(n_435), .Y(n_434) );
INVx1_ASAP7_75t_L g274 ( .A(n_275), .Y(n_274) );
NAND2xp5_ASAP7_75t_L g275 ( .A(n_276), .B(n_277), .Y(n_275) );
OAI322xp33_ASAP7_75t_L g321 ( .A1(n_277), .A2(n_281), .A3(n_290), .B1(n_322), .B2(n_325), .C1(n_326), .C2(n_327), .Y(n_321) );
NAND2xp5_ASAP7_75t_L g329 ( .A(n_277), .B(n_330), .Y(n_329) );
NAND2xp5_ASAP7_75t_L g392 ( .A(n_277), .B(n_393), .Y(n_392) );
AND2x2_ASAP7_75t_L g300 ( .A(n_278), .B(n_301), .Y(n_300) );
OR2x2_ASAP7_75t_L g332 ( .A(n_278), .B(n_333), .Y(n_332) );
NAND2xp5_ASAP7_75t_L g432 ( .A(n_278), .B(n_433), .Y(n_432) );
INVx1_ASAP7_75t_L g279 ( .A(n_280), .Y(n_279) );
INVx1_ASAP7_75t_L g393 ( .A(n_281), .Y(n_393) );
HB1xp67_ASAP7_75t_L g324 ( .A(n_282), .Y(n_324) );
INVx1_ASAP7_75t_L g283 ( .A(n_284), .Y(n_283) );
OAI21xp5_ASAP7_75t_L g285 ( .A1(n_286), .A2(n_289), .B(n_292), .Y(n_285) );
AND2x2_ASAP7_75t_L g286 ( .A(n_287), .B(n_288), .Y(n_286) );
NAND2xp5_ASAP7_75t_L g335 ( .A(n_288), .B(n_336), .Y(n_335) );
AOI322xp5_ASAP7_75t_SL g430 ( .A1(n_288), .A2(n_294), .A3(n_411), .B1(n_429), .B2(n_431), .C1(n_434), .C2(n_437), .Y(n_430) );
INVx1_ASAP7_75t_L g289 ( .A(n_290), .Y(n_289) );
OAI21xp33_ASAP7_75t_L g293 ( .A1(n_294), .A2(n_295), .B(n_309), .Y(n_293) );
NAND2xp5_ASAP7_75t_L g326 ( .A(n_294), .B(n_304), .Y(n_326) );
INVx2_ASAP7_75t_SL g336 ( .A(n_294), .Y(n_336) );
INVx1_ASAP7_75t_L g296 ( .A(n_297), .Y(n_296) );
NAND2xp5_ASAP7_75t_L g297 ( .A(n_298), .B(n_300), .Y(n_297) );
INVx1_ASAP7_75t_SL g361 ( .A(n_300), .Y(n_361) );
HB1xp67_ASAP7_75t_L g331 ( .A(n_301), .Y(n_331) );
INVx1_ASAP7_75t_L g302 ( .A(n_303), .Y(n_302) );
HB1xp67_ASAP7_75t_L g303 ( .A(n_304), .Y(n_303) );
INVx1_ASAP7_75t_L g305 ( .A(n_306), .Y(n_305) );
AND2x2_ASAP7_75t_L g406 ( .A(n_307), .B(n_407), .Y(n_406) );
INVx1_ASAP7_75t_SL g307 ( .A(n_308), .Y(n_307) );
OR2x2_ASAP7_75t_L g360 ( .A(n_308), .B(n_361), .Y(n_360) );
AOI22xp33_ASAP7_75t_L g309 ( .A1(n_310), .A2(n_313), .B1(n_314), .B2(n_319), .Y(n_309) );
INVx1_ASAP7_75t_SL g310 ( .A(n_311), .Y(n_310) );
INVx1_ASAP7_75t_L g314 ( .A(n_315), .Y(n_314) );
NAND2xp5_ASAP7_75t_L g315 ( .A(n_316), .B(n_317), .Y(n_315) );
INVx1_ASAP7_75t_L g317 ( .A(n_318), .Y(n_317) );
NOR4xp75_ASAP7_75t_L g320 ( .A(n_321), .B(n_334), .C(n_354), .D(n_370), .Y(n_320) );
INVx1_ASAP7_75t_SL g322 ( .A(n_323), .Y(n_322) );
INVxp67_ASAP7_75t_L g327 ( .A(n_328), .Y(n_327) );
NAND2xp5_ASAP7_75t_SL g328 ( .A(n_329), .B(n_332), .Y(n_328) );
INVxp67_ASAP7_75t_L g330 ( .A(n_331), .Y(n_330) );
OAI22xp5_ASAP7_75t_L g408 ( .A1(n_332), .A2(n_409), .B1(n_412), .B2(n_413), .Y(n_408) );
OR2x2_ASAP7_75t_L g373 ( .A(n_333), .B(n_374), .Y(n_373) );
INVx2_ASAP7_75t_L g417 ( .A(n_333), .Y(n_417) );
OAI221xp5_ASAP7_75t_L g334 ( .A1(n_335), .A2(n_337), .B1(n_339), .B2(n_341), .C(n_342), .Y(n_334) );
INVx2_ASAP7_75t_L g353 ( .A(n_338), .Y(n_353) );
AND2x2_ASAP7_75t_L g410 ( .A(n_338), .B(n_411), .Y(n_410) );
INVx2_ASAP7_75t_L g339 ( .A(n_340), .Y(n_339) );
AOI22xp5_ASAP7_75t_L g342 ( .A1(n_343), .A2(n_346), .B1(n_348), .B2(n_350), .Y(n_342) );
INVx1_ASAP7_75t_SL g343 ( .A(n_344), .Y(n_343) );
INVx1_ASAP7_75t_L g346 ( .A(n_347), .Y(n_346) );
BUFx2_ASAP7_75t_L g348 ( .A(n_349), .Y(n_348) );
INVx1_ASAP7_75t_L g405 ( .A(n_349), .Y(n_405) );
AOI22xp5_ASAP7_75t_L g371 ( .A1(n_350), .A2(n_356), .B1(n_372), .B2(n_375), .Y(n_371) );
INVx1_ASAP7_75t_SL g350 ( .A(n_351), .Y(n_350) );
OR2x2_ASAP7_75t_L g351 ( .A(n_352), .B(n_353), .Y(n_351) );
OAI221xp5_ASAP7_75t_L g354 ( .A1(n_355), .A2(n_360), .B1(n_362), .B2(n_363), .C(n_784), .Y(n_354) );
AND2x2_ASAP7_75t_SL g356 ( .A(n_357), .B(n_359), .Y(n_356) );
INVx1_ASAP7_75t_L g357 ( .A(n_358), .Y(n_357) );
OR2x2_ASAP7_75t_L g422 ( .A(n_361), .B(n_423), .Y(n_422) );
INVxp67_ASAP7_75t_L g363 ( .A(n_364), .Y(n_363) );
AND2x2_ASAP7_75t_L g364 ( .A(n_365), .B(n_366), .Y(n_364) );
INVx2_ASAP7_75t_L g366 ( .A(n_367), .Y(n_366) );
OR2x2_ASAP7_75t_L g367 ( .A(n_368), .B(n_369), .Y(n_367) );
INVx1_ASAP7_75t_L g407 ( .A(n_369), .Y(n_407) );
NAND2xp5_ASAP7_75t_L g370 ( .A(n_371), .B(n_378), .Y(n_370) );
INVx1_ASAP7_75t_L g372 ( .A(n_373), .Y(n_372) );
INVx1_ASAP7_75t_L g376 ( .A(n_377), .Y(n_376) );
INVx2_ASAP7_75t_SL g380 ( .A(n_381), .Y(n_380) );
OR2x2_ASAP7_75t_L g381 ( .A(n_382), .B(n_383), .Y(n_381) );
INVx1_ASAP7_75t_SL g385 ( .A(n_386), .Y(n_385) );
AOI21xp33_ASAP7_75t_L g388 ( .A1(n_389), .A2(n_391), .B(n_392), .Y(n_388) );
NOR3xp33_ASAP7_75t_SL g394 ( .A(n_395), .B(n_400), .C(n_424), .Y(n_394) );
INVx1_ASAP7_75t_L g397 ( .A(n_398), .Y(n_397) );
NAND2xp5_ASAP7_75t_L g400 ( .A(n_401), .B(n_415), .Y(n_400) );
O2A1O1Ixp33_ASAP7_75t_L g401 ( .A1(n_402), .A2(n_404), .B(n_406), .C(n_408), .Y(n_401) );
INVx1_ASAP7_75t_L g402 ( .A(n_403), .Y(n_402) );
INVx1_ASAP7_75t_L g404 ( .A(n_405), .Y(n_404) );
AND2x4_ASAP7_75t_L g416 ( .A(n_407), .B(n_417), .Y(n_416) );
INVx1_ASAP7_75t_SL g409 ( .A(n_410), .Y(n_409) );
INVx1_ASAP7_75t_SL g413 ( .A(n_414), .Y(n_413) );
NAND2xp5_ASAP7_75t_SL g418 ( .A(n_419), .B(n_420), .Y(n_418) );
INVx1_ASAP7_75t_SL g421 ( .A(n_422), .Y(n_421) );
NAND4xp25_ASAP7_75t_SL g424 ( .A(n_425), .B(n_430), .C(n_438), .D(n_445), .Y(n_424) );
NAND2xp5_ASAP7_75t_L g425 ( .A(n_426), .B(n_429), .Y(n_425) );
INVx1_ASAP7_75t_SL g426 ( .A(n_427), .Y(n_426) );
INVxp67_ASAP7_75t_SL g431 ( .A(n_432), .Y(n_431) );
OAI21xp5_ASAP7_75t_SL g438 ( .A1(n_439), .A2(n_440), .B(n_442), .Y(n_438) );
INVx1_ASAP7_75t_L g443 ( .A(n_444), .Y(n_443) );
INVx3_ASAP7_75t_L g446 ( .A(n_447), .Y(n_446) );
AND2x4_ASAP7_75t_L g449 ( .A(n_450), .B(n_667), .Y(n_449) );
NOR3xp33_ASAP7_75t_L g450 ( .A(n_451), .B(n_603), .C(n_650), .Y(n_450) );
NAND4xp25_ASAP7_75t_SL g451 ( .A(n_452), .B(n_538), .C(n_556), .D(n_582), .Y(n_451) );
OAI21xp33_ASAP7_75t_SL g452 ( .A1(n_453), .A2(n_497), .B(n_498), .Y(n_452) );
NAND2xp5_ASAP7_75t_SL g453 ( .A(n_454), .B(n_482), .Y(n_453) );
INVx1_ASAP7_75t_L g718 ( .A(n_454), .Y(n_718) );
OR2x2_ASAP7_75t_L g454 ( .A(n_455), .B(n_462), .Y(n_454) );
INVx2_ASAP7_75t_L g542 ( .A(n_455), .Y(n_542) );
AND2x2_ASAP7_75t_L g562 ( .A(n_455), .B(n_563), .Y(n_562) );
OR2x2_ASAP7_75t_L g664 ( .A(n_455), .B(n_484), .Y(n_664) );
AND2x2_ASAP7_75t_L g724 ( .A(n_455), .B(n_543), .Y(n_724) );
INVx2_ASAP7_75t_L g455 ( .A(n_456), .Y(n_455) );
NAND2xp5_ASAP7_75t_L g576 ( .A(n_456), .B(n_577), .Y(n_576) );
INVx2_ASAP7_75t_L g456 ( .A(n_457), .Y(n_456) );
OR2x2_ASAP7_75t_L g608 ( .A(n_457), .B(n_465), .Y(n_608) );
BUFx3_ASAP7_75t_L g618 ( .A(n_457), .Y(n_618) );
AND2x2_ASAP7_75t_L g681 ( .A(n_457), .B(n_682), .Y(n_681) );
AND2x4_ASAP7_75t_L g457 ( .A(n_458), .B(n_459), .Y(n_457) );
AND2x4_ASAP7_75t_L g496 ( .A(n_458), .B(n_459), .Y(n_496) );
INVx1_ASAP7_75t_SL g462 ( .A(n_463), .Y(n_462) );
INVx1_ASAP7_75t_L g727 ( .A(n_463), .Y(n_727) );
AND2x2_ASAP7_75t_L g463 ( .A(n_464), .B(n_473), .Y(n_463) );
AND2x2_ASAP7_75t_L g495 ( .A(n_464), .B(n_496), .Y(n_495) );
INVx1_ASAP7_75t_L g682 ( .A(n_464), .Y(n_682) );
INVx2_ASAP7_75t_L g464 ( .A(n_465), .Y(n_464) );
AND2x2_ASAP7_75t_L g497 ( .A(n_465), .B(n_486), .Y(n_497) );
AND2x2_ASAP7_75t_L g559 ( .A(n_465), .B(n_473), .Y(n_559) );
INVx2_ASAP7_75t_L g564 ( .A(n_465), .Y(n_564) );
AND2x2_ASAP7_75t_L g566 ( .A(n_465), .B(n_474), .Y(n_566) );
NAND2xp5_ASAP7_75t_L g466 ( .A(n_467), .B(n_471), .Y(n_466) );
INVx1_ASAP7_75t_L g544 ( .A(n_473), .Y(n_544) );
INVx2_ASAP7_75t_L g548 ( .A(n_473), .Y(n_548) );
AND2x4_ASAP7_75t_SL g579 ( .A(n_473), .B(n_486), .Y(n_579) );
HB1xp67_ASAP7_75t_L g611 ( .A(n_473), .Y(n_611) );
INVx3_ASAP7_75t_L g473 ( .A(n_474), .Y(n_473) );
HB1xp67_ASAP7_75t_L g494 ( .A(n_474), .Y(n_494) );
NAND2xp5_ASAP7_75t_L g475 ( .A(n_476), .B(n_480), .Y(n_475) );
NAND2xp5_ASAP7_75t_L g482 ( .A(n_483), .B(n_495), .Y(n_482) );
AND2x2_ASAP7_75t_L g645 ( .A(n_483), .B(n_590), .Y(n_645) );
INVx2_ASAP7_75t_SL g733 ( .A(n_483), .Y(n_733) );
INVx1_ASAP7_75t_L g483 ( .A(n_484), .Y(n_483) );
NAND2xp5_ASAP7_75t_L g484 ( .A(n_485), .B(n_494), .Y(n_484) );
NAND2x1p5_ASAP7_75t_L g546 ( .A(n_485), .B(n_547), .Y(n_546) );
AND2x2_ASAP7_75t_L g653 ( .A(n_485), .B(n_566), .Y(n_653) );
INVx4_ASAP7_75t_L g485 ( .A(n_486), .Y(n_485) );
BUFx2_ASAP7_75t_L g541 ( .A(n_486), .Y(n_541) );
AND2x4_ASAP7_75t_L g543 ( .A(n_486), .B(n_544), .Y(n_543) );
NOR2x1_ASAP7_75t_L g563 ( .A(n_486), .B(n_564), .Y(n_563) );
INVx1_ASAP7_75t_L g636 ( .A(n_486), .Y(n_636) );
AND2x2_ASAP7_75t_L g655 ( .A(n_486), .B(n_594), .Y(n_655) );
AND2x2_ASAP7_75t_L g686 ( .A(n_486), .B(n_595), .Y(n_686) );
OR2x6_ASAP7_75t_L g486 ( .A(n_487), .B(n_493), .Y(n_486) );
AND2x2_ASAP7_75t_L g625 ( .A(n_495), .B(n_579), .Y(n_625) );
NAND2xp5_ASAP7_75t_SL g661 ( .A(n_495), .B(n_636), .Y(n_661) );
AOI22xp5_ASAP7_75t_L g735 ( .A1(n_495), .A2(n_736), .B1(n_738), .B2(n_739), .Y(n_735) );
AND2x2_ASAP7_75t_L g738 ( .A(n_495), .B(n_545), .Y(n_738) );
INVx3_ASAP7_75t_L g591 ( .A(n_496), .Y(n_591) );
AND2x2_ASAP7_75t_L g594 ( .A(n_496), .B(n_595), .Y(n_594) );
AND2x2_ASAP7_75t_L g610 ( .A(n_497), .B(n_611), .Y(n_610) );
INVx1_ASAP7_75t_L g619 ( .A(n_497), .Y(n_619) );
AND2x4_ASAP7_75t_SL g498 ( .A(n_499), .B(n_508), .Y(n_498) );
NAND2xp5_ASAP7_75t_L g630 ( .A(n_499), .B(n_631), .Y(n_630) );
AND2x2_ASAP7_75t_L g670 ( .A(n_499), .B(n_671), .Y(n_670) );
NOR3xp33_ASAP7_75t_L g722 ( .A(n_499), .B(n_632), .C(n_723), .Y(n_722) );
OR2x2_ASAP7_75t_L g740 ( .A(n_499), .B(n_634), .Y(n_740) );
INVx3_ASAP7_75t_L g499 ( .A(n_500), .Y(n_499) );
INVx1_ASAP7_75t_L g500 ( .A(n_501), .Y(n_500) );
OR2x2_ASAP7_75t_L g555 ( .A(n_501), .B(n_519), .Y(n_555) );
INVx1_ASAP7_75t_L g572 ( .A(n_501), .Y(n_572) );
INVx2_ASAP7_75t_L g585 ( .A(n_501), .Y(n_585) );
HB1xp67_ASAP7_75t_L g600 ( .A(n_501), .Y(n_600) );
AND2x2_ASAP7_75t_L g614 ( .A(n_501), .B(n_587), .Y(n_614) );
AND2x2_ASAP7_75t_L g693 ( .A(n_501), .B(n_510), .Y(n_693) );
AOI221xp5_ASAP7_75t_L g556 ( .A1(n_508), .A2(n_557), .B1(n_560), .B2(n_567), .C(n_573), .Y(n_556) );
AOI221xp5_ASAP7_75t_L g685 ( .A1(n_508), .A2(n_686), .B1(n_687), .B2(n_688), .C(n_689), .Y(n_685) );
AND2x2_ASAP7_75t_L g508 ( .A(n_509), .B(n_518), .Y(n_508) );
INVx2_ASAP7_75t_L g627 ( .A(n_509), .Y(n_627) );
AND2x2_ASAP7_75t_L g687 ( .A(n_509), .B(n_571), .Y(n_687) );
AND2x2_ASAP7_75t_L g697 ( .A(n_509), .B(n_583), .Y(n_697) );
OR2x2_ASAP7_75t_L g737 ( .A(n_509), .B(n_621), .Y(n_737) );
INVx2_ASAP7_75t_L g509 ( .A(n_510), .Y(n_509) );
OR2x2_ASAP7_75t_SL g554 ( .A(n_510), .B(n_555), .Y(n_554) );
NAND2x1_ASAP7_75t_L g570 ( .A(n_510), .B(n_519), .Y(n_570) );
INVx4_ASAP7_75t_L g599 ( .A(n_510), .Y(n_599) );
OR2x2_ASAP7_75t_L g641 ( .A(n_510), .B(n_528), .Y(n_641) );
OR2x6_ASAP7_75t_L g510 ( .A(n_511), .B(n_512), .Y(n_510) );
AND2x2_ASAP7_75t_L g692 ( .A(n_518), .B(n_693), .Y(n_692) );
AND2x2_ASAP7_75t_L g518 ( .A(n_519), .B(n_528), .Y(n_518) );
INVx2_ASAP7_75t_SL g580 ( .A(n_519), .Y(n_580) );
NOR2x1_ASAP7_75t_SL g586 ( .A(n_519), .B(n_587), .Y(n_586) );
AND2x2_ASAP7_75t_L g601 ( .A(n_519), .B(n_602), .Y(n_601) );
OR2x2_ASAP7_75t_L g632 ( .A(n_519), .B(n_599), .Y(n_632) );
AND2x2_ASAP7_75t_L g639 ( .A(n_519), .B(n_585), .Y(n_639) );
BUFx2_ASAP7_75t_L g673 ( .A(n_519), .Y(n_673) );
AND2x2_ASAP7_75t_L g684 ( .A(n_519), .B(n_599), .Y(n_684) );
OR2x6_ASAP7_75t_L g519 ( .A(n_520), .B(n_527), .Y(n_519) );
HB1xp67_ASAP7_75t_L g552 ( .A(n_528), .Y(n_552) );
AND2x2_ASAP7_75t_L g571 ( .A(n_528), .B(n_572), .Y(n_571) );
INVx2_ASAP7_75t_L g602 ( .A(n_528), .Y(n_602) );
AND2x2_ASAP7_75t_L g628 ( .A(n_528), .B(n_584), .Y(n_628) );
INVx3_ASAP7_75t_L g528 ( .A(n_529), .Y(n_528) );
AO21x2_ASAP7_75t_L g529 ( .A1(n_530), .A2(n_531), .B(n_537), .Y(n_529) );
AO21x1_ASAP7_75t_SL g587 ( .A1(n_530), .A2(n_531), .B(n_537), .Y(n_587) );
NAND2xp5_ASAP7_75t_L g531 ( .A(n_532), .B(n_536), .Y(n_531) );
OAI31xp33_ASAP7_75t_L g538 ( .A1(n_539), .A2(n_543), .A3(n_545), .B(n_549), .Y(n_538) );
INVx1_ASAP7_75t_L g539 ( .A(n_540), .Y(n_539) );
NAND2xp5_ASAP7_75t_L g540 ( .A(n_541), .B(n_542), .Y(n_540) );
INVx2_ASAP7_75t_L g647 ( .A(n_541), .Y(n_647) );
NOR2xp67_ASAP7_75t_L g557 ( .A(n_542), .B(n_558), .Y(n_557) );
AOI322xp5_ASAP7_75t_L g637 ( .A1(n_542), .A2(n_631), .A3(n_638), .B1(n_642), .B2(n_643), .C1(n_645), .C2(n_646), .Y(n_637) );
AND2x2_ASAP7_75t_L g709 ( .A(n_542), .B(n_686), .Y(n_709) );
AOI221xp5_ASAP7_75t_SL g622 ( .A1(n_543), .A2(n_623), .B1(n_625), .B2(n_626), .C(n_629), .Y(n_622) );
INVx2_ASAP7_75t_L g642 ( .A(n_543), .Y(n_642) );
NAND2xp5_ASAP7_75t_L g606 ( .A(n_545), .B(n_607), .Y(n_606) );
NAND2xp5_ASAP7_75t_L g741 ( .A(n_545), .B(n_638), .Y(n_741) );
INVx1_ASAP7_75t_L g545 ( .A(n_546), .Y(n_545) );
OR2x2_ASAP7_75t_L g616 ( .A(n_546), .B(n_591), .Y(n_616) );
INVx1_ASAP7_75t_SL g547 ( .A(n_548), .Y(n_547) );
AND2x2_ASAP7_75t_L g595 ( .A(n_548), .B(n_564), .Y(n_595) );
AND2x4_ASAP7_75t_L g549 ( .A(n_550), .B(n_553), .Y(n_549) );
INVx1_ASAP7_75t_L g550 ( .A(n_551), .Y(n_550) );
INVx1_ASAP7_75t_L g551 ( .A(n_552), .Y(n_551) );
INVx1_ASAP7_75t_L g666 ( .A(n_552), .Y(n_666) );
O2A1O1Ixp5_ASAP7_75t_L g657 ( .A1(n_553), .A2(n_658), .B(n_660), .C(n_662), .Y(n_657) );
INVx2_ASAP7_75t_L g553 ( .A(n_554), .Y(n_553) );
OAI22xp5_ASAP7_75t_L g689 ( .A1(n_554), .A2(n_690), .B1(n_691), .B2(n_694), .Y(n_689) );
OR2x2_ASAP7_75t_L g644 ( .A(n_555), .B(n_641), .Y(n_644) );
INVx1_ASAP7_75t_L g558 ( .A(n_559), .Y(n_558) );
NAND2xp5_ASAP7_75t_SL g560 ( .A(n_561), .B(n_565), .Y(n_560) );
INVx1_ASAP7_75t_L g561 ( .A(n_562), .Y(n_561) );
INVx1_ASAP7_75t_L g577 ( .A(n_564), .Y(n_577) );
INVx1_ASAP7_75t_L g565 ( .A(n_566), .Y(n_565) );
NAND2xp5_ASAP7_75t_L g589 ( .A(n_566), .B(n_590), .Y(n_589) );
INVx1_ASAP7_75t_L g567 ( .A(n_568), .Y(n_567) );
NAND2xp5_ASAP7_75t_L g568 ( .A(n_569), .B(n_571), .Y(n_568) );
INVx3_ASAP7_75t_L g569 ( .A(n_570), .Y(n_569) );
OR2x2_ASAP7_75t_L g620 ( .A(n_570), .B(n_621), .Y(n_620) );
NAND2xp5_ASAP7_75t_L g663 ( .A(n_570), .B(n_571), .Y(n_663) );
OR2x2_ASAP7_75t_L g665 ( .A(n_570), .B(n_666), .Y(n_665) );
NOR2xp33_ASAP7_75t_L g713 ( .A(n_570), .B(n_714), .Y(n_713) );
BUFx2_ASAP7_75t_L g581 ( .A(n_572), .Y(n_581) );
NOR4xp25_ASAP7_75t_L g573 ( .A(n_574), .B(n_578), .C(n_580), .D(n_581), .Y(n_573) );
INVx1_ASAP7_75t_L g574 ( .A(n_575), .Y(n_574) );
AND2x2_ASAP7_75t_L g701 ( .A(n_575), .B(n_702), .Y(n_701) );
AND2x2_ASAP7_75t_L g729 ( .A(n_575), .B(n_578), .Y(n_729) );
INVx2_ASAP7_75t_L g575 ( .A(n_576), .Y(n_575) );
INVx1_ASAP7_75t_L g659 ( .A(n_577), .Y(n_659) );
NAND2xp5_ASAP7_75t_L g694 ( .A(n_578), .B(n_607), .Y(n_694) );
AOI321xp33_ASAP7_75t_L g696 ( .A1(n_578), .A2(n_697), .A3(n_698), .B1(n_699), .B2(n_701), .C(n_704), .Y(n_696) );
INVx2_ASAP7_75t_SL g578 ( .A(n_579), .Y(n_578) );
AND2x2_ASAP7_75t_SL g658 ( .A(n_579), .B(n_659), .Y(n_658) );
NAND2xp5_ASAP7_75t_L g680 ( .A(n_579), .B(n_618), .Y(n_680) );
NAND2xp5_ASAP7_75t_L g707 ( .A(n_580), .B(n_602), .Y(n_707) );
OR2x2_ASAP7_75t_L g734 ( .A(n_581), .B(n_618), .Y(n_734) );
AOI21xp5_ASAP7_75t_L g582 ( .A1(n_583), .A2(n_588), .B(n_592), .Y(n_582) );
AND2x2_ASAP7_75t_L g623 ( .A(n_583), .B(n_624), .Y(n_623) );
AND2x2_ASAP7_75t_L g583 ( .A(n_584), .B(n_586), .Y(n_583) );
INVx1_ASAP7_75t_L g584 ( .A(n_585), .Y(n_584) );
AND2x2_ASAP7_75t_L g649 ( .A(n_585), .B(n_587), .Y(n_649) );
INVx2_ASAP7_75t_L g634 ( .A(n_586), .Y(n_634) );
INVx1_ASAP7_75t_SL g588 ( .A(n_589), .Y(n_588) );
NOR2xp33_ASAP7_75t_L g704 ( .A(n_589), .B(n_705), .Y(n_704) );
OR2x2_ASAP7_75t_L g690 ( .A(n_590), .B(n_642), .Y(n_690) );
INVx2_ASAP7_75t_L g590 ( .A(n_591), .Y(n_590) );
AND2x2_ASAP7_75t_L g648 ( .A(n_591), .B(n_649), .Y(n_648) );
NOR2x1_ASAP7_75t_L g726 ( .A(n_591), .B(n_727), .Y(n_726) );
NOR2xp67_ASAP7_75t_L g592 ( .A(n_593), .B(n_596), .Y(n_592) );
INVx2_ASAP7_75t_L g593 ( .A(n_594), .Y(n_593) );
INVx1_ASAP7_75t_L g677 ( .A(n_595), .Y(n_677) );
INVx2_ASAP7_75t_L g596 ( .A(n_597), .Y(n_596) );
AND2x2_ASAP7_75t_L g597 ( .A(n_598), .B(n_601), .Y(n_597) );
NOR2xp67_ASAP7_75t_L g598 ( .A(n_599), .B(n_600), .Y(n_598) );
NAND2xp5_ASAP7_75t_L g613 ( .A(n_599), .B(n_614), .Y(n_613) );
INVx1_ASAP7_75t_L g624 ( .A(n_599), .Y(n_624) );
BUFx2_ASAP7_75t_L g706 ( .A(n_599), .Y(n_706) );
INVxp67_ASAP7_75t_L g714 ( .A(n_602), .Y(n_714) );
NAND3xp33_ASAP7_75t_L g603 ( .A(n_604), .B(n_622), .C(n_637), .Y(n_603) );
AOI21xp5_ASAP7_75t_L g604 ( .A1(n_605), .A2(n_612), .B(n_615), .Y(n_604) );
NAND2xp5_ASAP7_75t_L g605 ( .A(n_606), .B(n_609), .Y(n_605) );
INVx2_ASAP7_75t_SL g607 ( .A(n_608), .Y(n_607) );
OR2x2_ASAP7_75t_L g635 ( .A(n_608), .B(n_636), .Y(n_635) );
INVx2_ASAP7_75t_L g688 ( .A(n_609), .Y(n_688) );
INVx1_ASAP7_75t_L g609 ( .A(n_610), .Y(n_609) );
INVx2_ASAP7_75t_L g703 ( .A(n_611), .Y(n_703) );
AOI21xp5_ASAP7_75t_L g708 ( .A1(n_612), .A2(n_709), .B(n_710), .Y(n_708) );
INVx1_ASAP7_75t_SL g612 ( .A(n_613), .Y(n_612) );
INVx2_ASAP7_75t_SL g621 ( .A(n_614), .Y(n_621) );
AND2x2_ASAP7_75t_L g683 ( .A(n_614), .B(n_684), .Y(n_683) );
AOI21xp33_ASAP7_75t_L g615 ( .A1(n_616), .A2(n_617), .B(n_620), .Y(n_615) );
OAI22xp5_ASAP7_75t_L g662 ( .A1(n_616), .A2(n_663), .B1(n_664), .B2(n_665), .Y(n_662) );
OR2x2_ASAP7_75t_L g617 ( .A(n_618), .B(n_619), .Y(n_617) );
INVx1_ASAP7_75t_L g652 ( .A(n_618), .Y(n_652) );
OR2x2_ASAP7_75t_L g700 ( .A(n_621), .B(n_632), .Y(n_700) );
NOR4xp25_ASAP7_75t_L g732 ( .A(n_624), .B(n_673), .C(n_733), .D(n_734), .Y(n_732) );
AND2x2_ASAP7_75t_L g626 ( .A(n_627), .B(n_628), .Y(n_626) );
OR2x2_ASAP7_75t_L g633 ( .A(n_627), .B(n_634), .Y(n_633) );
NAND2xp5_ASAP7_75t_L g731 ( .A(n_627), .B(n_649), .Y(n_731) );
AOI21xp33_ASAP7_75t_SL g629 ( .A1(n_630), .A2(n_633), .B(n_635), .Y(n_629) );
INVx2_ASAP7_75t_SL g631 ( .A(n_632), .Y(n_631) );
OR2x2_ASAP7_75t_L g720 ( .A(n_632), .B(n_721), .Y(n_720) );
INVx1_ASAP7_75t_L g728 ( .A(n_634), .Y(n_728) );
AND2x4_ASAP7_75t_L g638 ( .A(n_639), .B(n_640), .Y(n_638) );
INVxp67_ASAP7_75t_L g656 ( .A(n_639), .Y(n_656) );
INVx1_ASAP7_75t_L g640 ( .A(n_641), .Y(n_640) );
OR2x2_ASAP7_75t_L g672 ( .A(n_641), .B(n_673), .Y(n_672) );
INVx1_ASAP7_75t_L g643 ( .A(n_644), .Y(n_643) );
AND2x2_ASAP7_75t_L g646 ( .A(n_647), .B(n_648), .Y(n_646) );
AND2x2_ASAP7_75t_L g675 ( .A(n_647), .B(n_676), .Y(n_675) );
INVx1_ASAP7_75t_L g721 ( .A(n_649), .Y(n_721) );
A2O1A1Ixp33_ASAP7_75t_L g650 ( .A1(n_651), .A2(n_654), .B(n_656), .C(n_657), .Y(n_650) );
NAND2xp5_ASAP7_75t_L g651 ( .A(n_652), .B(n_653), .Y(n_651) );
INVx1_ASAP7_75t_L g711 ( .A(n_653), .Y(n_711) );
INVx1_ASAP7_75t_L g654 ( .A(n_655), .Y(n_654) );
INVxp67_ASAP7_75t_L g715 ( .A(n_658), .Y(n_715) );
INVx1_ASAP7_75t_L g660 ( .A(n_661), .Y(n_660) );
NOR3xp33_ASAP7_75t_L g667 ( .A(n_668), .B(n_695), .C(n_716), .Y(n_667) );
OAI211xp5_ASAP7_75t_SL g668 ( .A1(n_669), .A2(n_674), .B(n_678), .C(n_685), .Y(n_668) );
INVx1_ASAP7_75t_L g669 ( .A(n_670), .Y(n_669) );
INVx1_ASAP7_75t_SL g671 ( .A(n_672), .Y(n_671) );
INVxp67_ASAP7_75t_L g674 ( .A(n_675), .Y(n_674) );
INVx2_ASAP7_75t_L g676 ( .A(n_677), .Y(n_676) );
OAI21xp5_ASAP7_75t_SL g678 ( .A1(n_679), .A2(n_681), .B(n_683), .Y(n_678) );
INVx1_ASAP7_75t_L g679 ( .A(n_680), .Y(n_679) );
O2A1O1Ixp33_ASAP7_75t_L g717 ( .A1(n_681), .A2(n_718), .B(n_719), .C(n_722), .Y(n_717) );
BUFx2_ASAP7_75t_L g698 ( .A(n_682), .Y(n_698) );
INVx2_ASAP7_75t_L g691 ( .A(n_692), .Y(n_691) );
NAND2xp5_ASAP7_75t_L g695 ( .A(n_696), .B(n_708), .Y(n_695) );
INVx2_ASAP7_75t_L g699 ( .A(n_700), .Y(n_699) );
INVx2_ASAP7_75t_L g702 ( .A(n_703), .Y(n_702) );
OAI22xp5_ASAP7_75t_L g710 ( .A1(n_705), .A2(n_711), .B1(n_712), .B2(n_715), .Y(n_710) );
OR2x2_ASAP7_75t_L g705 ( .A(n_706), .B(n_707), .Y(n_705) );
INVx1_ASAP7_75t_L g712 ( .A(n_713), .Y(n_712) );
NAND4xp25_ASAP7_75t_L g716 ( .A(n_717), .B(n_725), .C(n_735), .D(n_741), .Y(n_716) );
INVx2_ASAP7_75t_L g719 ( .A(n_720), .Y(n_719) );
INVx1_ASAP7_75t_L g723 ( .A(n_724), .Y(n_723) );
AOI221xp5_ASAP7_75t_L g725 ( .A1(n_726), .A2(n_728), .B1(n_729), .B2(n_730), .C(n_732), .Y(n_725) );
INVx1_ASAP7_75t_L g730 ( .A(n_731), .Y(n_730) );
INVx1_ASAP7_75t_L g736 ( .A(n_737), .Y(n_736) );
INVx1_ASAP7_75t_L g739 ( .A(n_740), .Y(n_739) );
INVx1_ASAP7_75t_SL g742 ( .A(n_743), .Y(n_742) );
CKINVDCx11_ASAP7_75t_R g743 ( .A(n_744), .Y(n_743) );
INVx1_ASAP7_75t_L g749 ( .A(n_746), .Y(n_749) );
NOR2xp33_ASAP7_75t_L g752 ( .A(n_753), .B(n_754), .Y(n_752) );
INVx1_ASAP7_75t_L g754 ( .A(n_755), .Y(n_754) );
INVx3_ASAP7_75t_L g755 ( .A(n_756), .Y(n_755) );
INVxp33_ASAP7_75t_L g757 ( .A(n_758), .Y(n_757) );
AOI21xp5_ASAP7_75t_L g772 ( .A1(n_758), .A2(n_773), .B(n_774), .Y(n_772) );
NOR2xp33_ASAP7_75t_L g758 ( .A(n_759), .B(n_760), .Y(n_758) );
INVx1_ASAP7_75t_SL g760 ( .A(n_761), .Y(n_760) );
BUFx2_ASAP7_75t_L g761 ( .A(n_762), .Y(n_761) );
CKINVDCx20_ASAP7_75t_R g762 ( .A(n_763), .Y(n_762) );
BUFx3_ASAP7_75t_L g763 ( .A(n_764), .Y(n_763) );
BUFx2_ASAP7_75t_R g773 ( .A(n_764), .Y(n_773) );
BUFx3_ASAP7_75t_L g765 ( .A(n_766), .Y(n_765) );
CKINVDCx20_ASAP7_75t_R g766 ( .A(n_767), .Y(n_766) );
HB1xp67_ASAP7_75t_L g767 ( .A(n_768), .Y(n_767) );
NOR2xp67_ASAP7_75t_L g769 ( .A(n_770), .B(n_772), .Y(n_769) );
INVx2_ASAP7_75t_SL g770 ( .A(n_771), .Y(n_770) );
INVx2_ASAP7_75t_L g774 ( .A(n_775), .Y(n_774) );
NOR2xp33_ASAP7_75t_L g779 ( .A(n_780), .B(n_781), .Y(n_779) );
HB1xp67_ASAP7_75t_L g781 ( .A(n_782), .Y(n_781) );
endmodule