module fake_jpeg_26797_n_226 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_226);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_226;

wire n_159;
wire n_117;
wire n_144;
wire n_225;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_84;
wire n_59;
wire n_98;
wire n_178;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_57;
wire n_21;
wire n_223;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_44;
wire n_24;
wire n_143;
wire n_202;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_37;
wire n_121;
wire n_99;
wire n_102;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_212;
wire n_131;
wire n_56;
wire n_211;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_216;
wire n_217;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_118;
wire n_100;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

NOR2xp33_ASAP7_75t_L g16 ( 
.A(n_6),
.B(n_2),
.Y(n_16)
);

BUFx24_ASAP7_75t_L g17 ( 
.A(n_6),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_0),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_6),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_9),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_10),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_14),
.Y(n_22)
);

BUFx5_ASAP7_75t_L g23 ( 
.A(n_12),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_14),
.Y(n_24)
);

INVx11_ASAP7_75t_L g25 ( 
.A(n_0),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_0),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_12),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_9),
.Y(n_28)
);

INVx3_ASAP7_75t_L g29 ( 
.A(n_9),
.Y(n_29)
);

BUFx3_ASAP7_75t_L g30 ( 
.A(n_10),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_8),
.Y(n_31)
);

BUFx5_ASAP7_75t_L g32 ( 
.A(n_15),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_1),
.Y(n_33)
);

INVx2_ASAP7_75t_L g34 ( 
.A(n_25),
.Y(n_34)
);

INVx2_ASAP7_75t_L g55 ( 
.A(n_34),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_17),
.Y(n_35)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_35),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_17),
.Y(n_36)
);

INVx4_ASAP7_75t_L g51 ( 
.A(n_36),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_17),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_37),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_SL g38 ( 
.A(n_16),
.B(n_1),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_SL g52 ( 
.A(n_38),
.B(n_40),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_17),
.Y(n_39)
);

BUFx12f_ASAP7_75t_L g48 ( 
.A(n_39),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g40 ( 
.A(n_16),
.B(n_1),
.Y(n_40)
);

BUFx5_ASAP7_75t_L g41 ( 
.A(n_17),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_41),
.B(n_44),
.Y(n_53)
);

INVx2_ASAP7_75t_L g42 ( 
.A(n_25),
.Y(n_42)
);

AND2x2_ASAP7_75t_L g62 ( 
.A(n_42),
.B(n_26),
.Y(n_62)
);

INVx8_ASAP7_75t_L g43 ( 
.A(n_25),
.Y(n_43)
);

INVx5_ASAP7_75t_L g65 ( 
.A(n_43),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g44 ( 
.A(n_22),
.B(n_15),
.Y(n_44)
);

INVx6_ASAP7_75t_L g45 ( 
.A(n_20),
.Y(n_45)
);

OAI21xp33_ASAP7_75t_L g47 ( 
.A1(n_45),
.A2(n_29),
.B(n_32),
.Y(n_47)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_43),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_46),
.B(n_49),
.Y(n_70)
);

OA22x2_ASAP7_75t_L g79 ( 
.A1(n_47),
.A2(n_39),
.B1(n_37),
.B2(n_36),
.Y(n_79)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_43),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_35),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_50),
.B(n_57),
.Y(n_77)
);

OAI22xp5_ASAP7_75t_SL g54 ( 
.A1(n_45),
.A2(n_29),
.B1(n_33),
.B2(n_18),
.Y(n_54)
);

AOI22xp5_ASAP7_75t_L g74 ( 
.A1(n_54),
.A2(n_60),
.B1(n_66),
.B2(n_62),
.Y(n_74)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_34),
.Y(n_57)
);

AOI22xp33_ASAP7_75t_L g59 ( 
.A1(n_45),
.A2(n_29),
.B1(n_19),
.B2(n_33),
.Y(n_59)
);

OAI22xp5_ASAP7_75t_L g71 ( 
.A1(n_59),
.A2(n_31),
.B1(n_26),
.B2(n_20),
.Y(n_71)
);

OAI22xp5_ASAP7_75t_L g60 ( 
.A1(n_38),
.A2(n_19),
.B1(n_18),
.B2(n_21),
.Y(n_60)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_42),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_SL g88 ( 
.A(n_61),
.B(n_39),
.Y(n_88)
);

CKINVDCx16_ASAP7_75t_R g76 ( 
.A(n_62),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_40),
.B(n_27),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_63),
.B(n_23),
.Y(n_69)
);

AOI21xp33_ASAP7_75t_L g64 ( 
.A1(n_41),
.A2(n_27),
.B(n_24),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_R g78 ( 
.A(n_64),
.B(n_30),
.Y(n_78)
);

OAI22xp33_ASAP7_75t_SL g66 ( 
.A1(n_35),
.A2(n_24),
.B1(n_22),
.B2(n_26),
.Y(n_66)
);

AOI22xp33_ASAP7_75t_SL g67 ( 
.A1(n_65),
.A2(n_21),
.B1(n_28),
.B2(n_32),
.Y(n_67)
);

CKINVDCx16_ASAP7_75t_R g104 ( 
.A(n_67),
.Y(n_104)
);

A2O1A1Ixp33_ASAP7_75t_L g68 ( 
.A1(n_52),
.A2(n_28),
.B(n_32),
.C(n_23),
.Y(n_68)
);

OAI21xp5_ASAP7_75t_L g93 ( 
.A1(n_68),
.A2(n_53),
.B(n_57),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_69),
.B(n_72),
.Y(n_90)
);

AOI22xp5_ASAP7_75t_L g91 ( 
.A1(n_71),
.A2(n_73),
.B1(n_58),
.B2(n_61),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_52),
.B(n_30),
.Y(n_72)
);

OAI22xp33_ASAP7_75t_SL g73 ( 
.A1(n_54),
.A2(n_31),
.B1(n_20),
.B2(n_30),
.Y(n_73)
);

OR2x2_ASAP7_75t_L g106 ( 
.A(n_74),
.B(n_78),
.Y(n_106)
);

BUFx2_ASAP7_75t_SL g75 ( 
.A(n_48),
.Y(n_75)
);

CKINVDCx16_ASAP7_75t_R g108 ( 
.A(n_75),
.Y(n_108)
);

OR2x2_ASAP7_75t_L g112 ( 
.A(n_79),
.B(n_48),
.Y(n_112)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_62),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_SL g92 ( 
.A(n_80),
.B(n_84),
.Y(n_92)
);

BUFx2_ASAP7_75t_L g81 ( 
.A(n_56),
.Y(n_81)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_81),
.Y(n_95)
);

INVx2_ASAP7_75t_L g82 ( 
.A(n_55),
.Y(n_82)
);

BUFx6f_ASAP7_75t_L g102 ( 
.A(n_82),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_L g83 ( 
.A(n_60),
.B(n_31),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g97 ( 
.A(n_83),
.B(n_37),
.Y(n_97)
);

CKINVDCx20_ASAP7_75t_R g84 ( 
.A(n_50),
.Y(n_84)
);

CKINVDCx20_ASAP7_75t_R g85 ( 
.A(n_56),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_SL g96 ( 
.A(n_85),
.B(n_49),
.Y(n_96)
);

INVx2_ASAP7_75t_L g86 ( 
.A(n_55),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_86),
.B(n_87),
.Y(n_94)
);

INVx6_ASAP7_75t_L g87 ( 
.A(n_56),
.Y(n_87)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_88),
.Y(n_99)
);

INVx2_ASAP7_75t_L g89 ( 
.A(n_58),
.Y(n_89)
);

CKINVDCx20_ASAP7_75t_R g100 ( 
.A(n_89),
.Y(n_100)
);

OAI22xp5_ASAP7_75t_L g118 ( 
.A1(n_91),
.A2(n_93),
.B1(n_97),
.B2(n_88),
.Y(n_118)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_96),
.Y(n_114)
);

INVx5_ASAP7_75t_L g98 ( 
.A(n_81),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g123 ( 
.A(n_98),
.B(n_89),
.Y(n_123)
);

OA22x2_ASAP7_75t_L g101 ( 
.A1(n_79),
.A2(n_51),
.B1(n_65),
.B2(n_36),
.Y(n_101)
);

OAI21xp5_ASAP7_75t_SL g127 ( 
.A1(n_101),
.A2(n_112),
.B(n_71),
.Y(n_127)
);

CKINVDCx20_ASAP7_75t_R g103 ( 
.A(n_84),
.Y(n_103)
);

CKINVDCx20_ASAP7_75t_R g126 ( 
.A(n_103),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_L g105 ( 
.A(n_76),
.B(n_46),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_L g115 ( 
.A(n_105),
.B(n_113),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_SL g107 ( 
.A(n_80),
.B(n_83),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_SL g133 ( 
.A(n_107),
.B(n_79),
.Y(n_133)
);

OAI22xp5_ASAP7_75t_SL g109 ( 
.A1(n_74),
.A2(n_51),
.B1(n_48),
.B2(n_4),
.Y(n_109)
);

AOI22xp5_ASAP7_75t_SL g120 ( 
.A1(n_109),
.A2(n_111),
.B1(n_87),
.B2(n_85),
.Y(n_120)
);

XNOR2xp5_ASAP7_75t_L g110 ( 
.A(n_78),
.B(n_2),
.Y(n_110)
);

XOR2xp5_ASAP7_75t_L g117 ( 
.A(n_110),
.B(n_68),
.Y(n_117)
);

OAI22xp5_ASAP7_75t_SL g111 ( 
.A1(n_76),
.A2(n_48),
.B1(n_3),
.B2(n_4),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_L g113 ( 
.A(n_77),
.B(n_2),
.Y(n_113)
);

INVxp67_ASAP7_75t_L g116 ( 
.A(n_94),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_SL g151 ( 
.A(n_116),
.B(n_119),
.Y(n_151)
);

XNOR2xp5_ASAP7_75t_L g150 ( 
.A(n_117),
.B(n_104),
.Y(n_150)
);

AOI22xp5_ASAP7_75t_L g140 ( 
.A1(n_118),
.A2(n_99),
.B1(n_104),
.B2(n_97),
.Y(n_140)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_103),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_L g137 ( 
.A(n_120),
.B(n_122),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_L g121 ( 
.A(n_106),
.B(n_77),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_L g139 ( 
.A(n_121),
.B(n_128),
.Y(n_139)
);

BUFx24_ASAP7_75t_L g122 ( 
.A(n_102),
.Y(n_122)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_123),
.Y(n_141)
);

NOR2x1_ASAP7_75t_L g124 ( 
.A(n_93),
.B(n_79),
.Y(n_124)
);

OR2x2_ASAP7_75t_L g155 ( 
.A(n_124),
.B(n_133),
.Y(n_155)
);

INVx2_ASAP7_75t_L g125 ( 
.A(n_102),
.Y(n_125)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_125),
.Y(n_143)
);

AOI21xp5_ASAP7_75t_L g152 ( 
.A1(n_127),
.A2(n_101),
.B(n_108),
.Y(n_152)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_109),
.Y(n_128)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_100),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_L g142 ( 
.A(n_129),
.B(n_130),
.Y(n_142)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_100),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_L g131 ( 
.A(n_90),
.B(n_70),
.Y(n_131)
);

CKINVDCx20_ASAP7_75t_R g138 ( 
.A(n_131),
.Y(n_138)
);

MAJIxp5_ASAP7_75t_L g132 ( 
.A(n_106),
.B(n_70),
.C(n_82),
.Y(n_132)
);

MAJIxp5_ASAP7_75t_L g154 ( 
.A(n_132),
.B(n_102),
.C(n_95),
.Y(n_154)
);

INVxp67_ASAP7_75t_L g134 ( 
.A(n_92),
.Y(n_134)
);

INVx2_ASAP7_75t_SL g153 ( 
.A(n_134),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_L g135 ( 
.A(n_107),
.B(n_86),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_L g144 ( 
.A(n_135),
.B(n_112),
.Y(n_144)
);

AOI322xp5_ASAP7_75t_SL g136 ( 
.A1(n_117),
.A2(n_110),
.A3(n_111),
.B1(n_113),
.B2(n_13),
.C1(n_105),
.C2(n_99),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_L g162 ( 
.A(n_136),
.B(n_147),
.Y(n_162)
);

OAI22xp5_ASAP7_75t_L g158 ( 
.A1(n_140),
.A2(n_128),
.B1(n_120),
.B2(n_115),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_L g170 ( 
.A(n_144),
.B(n_146),
.Y(n_170)
);

XNOR2x1_ASAP7_75t_SL g145 ( 
.A(n_121),
.B(n_101),
.Y(n_145)
);

OAI21xp5_ASAP7_75t_SL g166 ( 
.A1(n_145),
.A2(n_152),
.B(n_146),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_L g146 ( 
.A(n_126),
.B(n_101),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_L g147 ( 
.A(n_126),
.B(n_135),
.Y(n_147)
);

XOR2xp5_ASAP7_75t_L g148 ( 
.A(n_132),
.B(n_91),
.Y(n_148)
);

XOR2xp5_ASAP7_75t_L g169 ( 
.A(n_148),
.B(n_81),
.Y(n_169)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_129),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_L g168 ( 
.A(n_149),
.B(n_125),
.Y(n_168)
);

XNOR2xp5_ASAP7_75t_L g163 ( 
.A(n_150),
.B(n_127),
.Y(n_163)
);

MAJIxp5_ASAP7_75t_L g159 ( 
.A(n_154),
.B(n_156),
.C(n_119),
.Y(n_159)
);

MAJIxp5_ASAP7_75t_L g156 ( 
.A(n_115),
.B(n_95),
.C(n_98),
.Y(n_156)
);

HB1xp67_ASAP7_75t_L g157 ( 
.A(n_156),
.Y(n_157)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_157),
.Y(n_180)
);

AOI22xp5_ASAP7_75t_L g187 ( 
.A1(n_158),
.A2(n_152),
.B1(n_153),
.B2(n_141),
.Y(n_187)
);

XNOR2xp5_ASAP7_75t_L g176 ( 
.A(n_159),
.B(n_160),
.Y(n_176)
);

MAJIxp5_ASAP7_75t_L g160 ( 
.A(n_148),
.B(n_130),
.C(n_124),
.Y(n_160)
);

NOR2xp33_ASAP7_75t_SL g161 ( 
.A(n_138),
.B(n_114),
.Y(n_161)
);

NOR2xp33_ASAP7_75t_SL g174 ( 
.A(n_161),
.B(n_173),
.Y(n_174)
);

XOR2xp5_ASAP7_75t_L g182 ( 
.A(n_163),
.B(n_166),
.Y(n_182)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_142),
.Y(n_164)
);

NOR2xp33_ASAP7_75t_L g177 ( 
.A(n_164),
.B(n_165),
.Y(n_177)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_142),
.Y(n_165)
);

AOI22xp5_ASAP7_75t_L g167 ( 
.A1(n_145),
.A2(n_116),
.B1(n_134),
.B2(n_114),
.Y(n_167)
);

OAI22xp5_ASAP7_75t_SL g184 ( 
.A1(n_167),
.A2(n_172),
.B1(n_140),
.B2(n_139),
.Y(n_184)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_168),
.Y(n_181)
);

AND2x2_ASAP7_75t_L g179 ( 
.A(n_169),
.B(n_154),
.Y(n_179)
);

INVx1_ASAP7_75t_SL g171 ( 
.A(n_147),
.Y(n_171)
);

NOR2xp33_ASAP7_75t_L g185 ( 
.A(n_171),
.B(n_153),
.Y(n_185)
);

AOI22xp5_ASAP7_75t_L g172 ( 
.A1(n_137),
.A2(n_122),
.B1(n_13),
.B2(n_5),
.Y(n_172)
);

NOR2xp33_ASAP7_75t_L g173 ( 
.A(n_153),
.B(n_141),
.Y(n_173)
);

HB1xp67_ASAP7_75t_L g175 ( 
.A(n_159),
.Y(n_175)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_175),
.Y(n_191)
);

NAND3xp33_ASAP7_75t_L g178 ( 
.A(n_162),
.B(n_139),
.C(n_144),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_SL g190 ( 
.A(n_178),
.B(n_179),
.Y(n_190)
);

INVx1_ASAP7_75t_SL g183 ( 
.A(n_170),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_L g189 ( 
.A(n_183),
.B(n_186),
.Y(n_189)
);

AOI22xp5_ASAP7_75t_L g194 ( 
.A1(n_184),
.A2(n_151),
.B1(n_172),
.B2(n_155),
.Y(n_194)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_185),
.Y(n_196)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_170),
.Y(n_186)
);

OAI22xp5_ASAP7_75t_SL g188 ( 
.A1(n_187),
.A2(n_167),
.B1(n_171),
.B2(n_160),
.Y(n_188)
);

AOI22xp5_ASAP7_75t_L g201 ( 
.A1(n_188),
.A2(n_195),
.B1(n_196),
.B2(n_181),
.Y(n_201)
);

XOR2xp5_ASAP7_75t_L g192 ( 
.A(n_182),
.B(n_169),
.Y(n_192)
);

XNOR2xp5_ASAP7_75t_L g202 ( 
.A(n_192),
.B(n_197),
.Y(n_202)
);

AOI321xp33_ASAP7_75t_L g193 ( 
.A1(n_178),
.A2(n_166),
.A3(n_163),
.B1(n_155),
.B2(n_150),
.C(n_149),
.Y(n_193)
);

OAI21xp5_ASAP7_75t_SL g204 ( 
.A1(n_193),
.A2(n_198),
.B(n_183),
.Y(n_204)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_194),
.Y(n_206)
);

OAI22xp5_ASAP7_75t_SL g195 ( 
.A1(n_187),
.A2(n_143),
.B1(n_122),
.B2(n_5),
.Y(n_195)
);

XNOR2xp5_ASAP7_75t_L g197 ( 
.A(n_176),
.B(n_182),
.Y(n_197)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_174),
.Y(n_198)
);

AOI21xp5_ASAP7_75t_L g199 ( 
.A1(n_191),
.A2(n_180),
.B(n_179),
.Y(n_199)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_199),
.Y(n_212)
);

AND2x2_ASAP7_75t_L g200 ( 
.A(n_190),
.B(n_177),
.Y(n_200)
);

NAND2xp5_ASAP7_75t_L g207 ( 
.A(n_200),
.B(n_201),
.Y(n_207)
);

HB1xp67_ASAP7_75t_L g203 ( 
.A(n_189),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_L g209 ( 
.A(n_203),
.B(n_205),
.Y(n_209)
);

AOI31xp67_ASAP7_75t_SL g208 ( 
.A1(n_204),
.A2(n_193),
.A3(n_176),
.B(n_192),
.Y(n_208)
);

CKINVDCx20_ASAP7_75t_R g205 ( 
.A(n_194),
.Y(n_205)
);

OR2x2_ASAP7_75t_L g214 ( 
.A(n_208),
.B(n_211),
.Y(n_214)
);

OA22x2_ASAP7_75t_L g210 ( 
.A1(n_206),
.A2(n_197),
.B1(n_122),
.B2(n_143),
.Y(n_210)
);

NOR2xp33_ASAP7_75t_L g215 ( 
.A(n_210),
.B(n_213),
.Y(n_215)
);

AOI22xp5_ASAP7_75t_L g211 ( 
.A1(n_200),
.A2(n_3),
.B1(n_4),
.B2(n_5),
.Y(n_211)
);

AOI22xp5_ASAP7_75t_L g213 ( 
.A1(n_203),
.A2(n_3),
.B1(n_7),
.B2(n_8),
.Y(n_213)
);

AOI21xp5_ASAP7_75t_L g216 ( 
.A1(n_212),
.A2(n_207),
.B(n_209),
.Y(n_216)
);

NAND2xp5_ASAP7_75t_L g220 ( 
.A(n_216),
.B(n_217),
.Y(n_220)
);

AOI21xp5_ASAP7_75t_L g217 ( 
.A1(n_210),
.A2(n_202),
.B(n_8),
.Y(n_217)
);

XNOR2xp5_ASAP7_75t_L g218 ( 
.A(n_213),
.B(n_7),
.Y(n_218)
);

NOR2xp33_ASAP7_75t_L g219 ( 
.A(n_218),
.B(n_214),
.Y(n_219)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_219),
.Y(n_223)
);

MAJIxp5_ASAP7_75t_L g221 ( 
.A(n_215),
.B(n_210),
.C(n_10),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_L g222 ( 
.A(n_221),
.B(n_7),
.Y(n_222)
);

OA21x2_ASAP7_75t_L g224 ( 
.A1(n_222),
.A2(n_220),
.B(n_11),
.Y(n_224)
);

AOI21x1_ASAP7_75t_L g225 ( 
.A1(n_224),
.A2(n_11),
.B(n_223),
.Y(n_225)
);

XNOR2xp5_ASAP7_75t_L g226 ( 
.A(n_225),
.B(n_11),
.Y(n_226)
);


endmodule