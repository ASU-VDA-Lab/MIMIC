module fake_netlist_6_3279_n_2299 (n_52, n_16, n_1, n_91, n_119, n_46, n_146, n_163, n_18, n_21, n_193, n_147, n_154, n_191, n_88, n_3, n_209, n_98, n_113, n_39, n_63, n_223, n_73, n_4, n_148, n_199, n_138, n_22, n_161, n_208, n_68, n_226, n_228, n_166, n_28, n_184, n_212, n_50, n_158, n_49, n_7, n_210, n_216, n_83, n_206, n_217, n_5, n_101, n_167, n_144, n_174, n_127, n_125, n_153, n_168, n_215, n_178, n_225, n_77, n_156, n_149, n_152, n_106, n_92, n_145, n_42, n_133, n_96, n_8, n_90, n_160, n_24, n_105, n_131, n_54, n_227, n_132, n_188, n_102, n_186, n_204, n_0, n_87, n_195, n_189, n_32, n_66, n_85, n_99, n_78, n_84, n_130, n_213, n_164, n_100, n_129, n_13, n_121, n_197, n_11, n_137, n_17, n_23, n_203, n_142, n_20, n_143, n_207, n_2, n_180, n_19, n_47, n_62, n_29, n_155, n_219, n_75, n_109, n_150, n_122, n_45, n_205, n_34, n_140, n_218, n_70, n_120, n_214, n_37, n_15, n_67, n_33, n_82, n_27, n_38, n_110, n_151, n_61, n_112, n_172, n_81, n_59, n_181, n_76, n_36, n_182, n_26, n_124, n_55, n_126, n_202, n_94, n_97, n_108, n_58, n_116, n_211, n_64, n_220, n_117, n_118, n_175, n_224, n_48, n_65, n_25, n_40, n_93, n_80, n_141, n_135, n_196, n_200, n_165, n_139, n_41, n_134, n_177, n_176, n_114, n_86, n_198, n_104, n_222, n_95, n_179, n_9, n_107, n_10, n_71, n_74, n_229, n_6, n_190, n_14, n_123, n_136, n_72, n_187, n_89, n_173, n_201, n_103, n_111, n_60, n_159, n_157, n_162, n_170, n_185, n_35, n_183, n_115, n_12, n_69, n_128, n_30, n_79, n_43, n_194, n_171, n_31, n_192, n_57, n_169, n_53, n_51, n_44, n_56, n_221, n_2299);

input n_52;
input n_16;
input n_1;
input n_91;
input n_119;
input n_46;
input n_146;
input n_163;
input n_18;
input n_21;
input n_193;
input n_147;
input n_154;
input n_191;
input n_88;
input n_3;
input n_209;
input n_98;
input n_113;
input n_39;
input n_63;
input n_223;
input n_73;
input n_4;
input n_148;
input n_199;
input n_138;
input n_22;
input n_161;
input n_208;
input n_68;
input n_226;
input n_228;
input n_166;
input n_28;
input n_184;
input n_212;
input n_50;
input n_158;
input n_49;
input n_7;
input n_210;
input n_216;
input n_83;
input n_206;
input n_217;
input n_5;
input n_101;
input n_167;
input n_144;
input n_174;
input n_127;
input n_125;
input n_153;
input n_168;
input n_215;
input n_178;
input n_225;
input n_77;
input n_156;
input n_149;
input n_152;
input n_106;
input n_92;
input n_145;
input n_42;
input n_133;
input n_96;
input n_8;
input n_90;
input n_160;
input n_24;
input n_105;
input n_131;
input n_54;
input n_227;
input n_132;
input n_188;
input n_102;
input n_186;
input n_204;
input n_0;
input n_87;
input n_195;
input n_189;
input n_32;
input n_66;
input n_85;
input n_99;
input n_78;
input n_84;
input n_130;
input n_213;
input n_164;
input n_100;
input n_129;
input n_13;
input n_121;
input n_197;
input n_11;
input n_137;
input n_17;
input n_23;
input n_203;
input n_142;
input n_20;
input n_143;
input n_207;
input n_2;
input n_180;
input n_19;
input n_47;
input n_62;
input n_29;
input n_155;
input n_219;
input n_75;
input n_109;
input n_150;
input n_122;
input n_45;
input n_205;
input n_34;
input n_140;
input n_218;
input n_70;
input n_120;
input n_214;
input n_37;
input n_15;
input n_67;
input n_33;
input n_82;
input n_27;
input n_38;
input n_110;
input n_151;
input n_61;
input n_112;
input n_172;
input n_81;
input n_59;
input n_181;
input n_76;
input n_36;
input n_182;
input n_26;
input n_124;
input n_55;
input n_126;
input n_202;
input n_94;
input n_97;
input n_108;
input n_58;
input n_116;
input n_211;
input n_64;
input n_220;
input n_117;
input n_118;
input n_175;
input n_224;
input n_48;
input n_65;
input n_25;
input n_40;
input n_93;
input n_80;
input n_141;
input n_135;
input n_196;
input n_200;
input n_165;
input n_139;
input n_41;
input n_134;
input n_177;
input n_176;
input n_114;
input n_86;
input n_198;
input n_104;
input n_222;
input n_95;
input n_179;
input n_9;
input n_107;
input n_10;
input n_71;
input n_74;
input n_229;
input n_6;
input n_190;
input n_14;
input n_123;
input n_136;
input n_72;
input n_187;
input n_89;
input n_173;
input n_201;
input n_103;
input n_111;
input n_60;
input n_159;
input n_157;
input n_162;
input n_170;
input n_185;
input n_35;
input n_183;
input n_115;
input n_12;
input n_69;
input n_128;
input n_30;
input n_79;
input n_43;
input n_194;
input n_171;
input n_31;
input n_192;
input n_57;
input n_169;
input n_53;
input n_51;
input n_44;
input n_56;
input n_221;

output n_2299;

wire n_992;
wire n_1671;
wire n_801;
wire n_1613;
wire n_1234;
wire n_1458;
wire n_1199;
wire n_1674;
wire n_741;
wire n_1027;
wire n_1351;
wire n_625;
wire n_1189;
wire n_1212;
wire n_726;
wire n_2157;
wire n_700;
wire n_1307;
wire n_2003;
wire n_1038;
wire n_578;
wire n_1581;
wire n_1003;
wire n_365;
wire n_1237;
wire n_1061;
wire n_1357;
wire n_1853;
wire n_783;
wire n_1738;
wire n_2243;
wire n_798;
wire n_1575;
wire n_1854;
wire n_1923;
wire n_509;
wire n_1342;
wire n_245;
wire n_1209;
wire n_1348;
wire n_1387;
wire n_2260;
wire n_677;
wire n_1708;
wire n_805;
wire n_1151;
wire n_396;
wire n_1739;
wire n_350;
wire n_2051;
wire n_1380;
wire n_442;
wire n_480;
wire n_1402;
wire n_1688;
wire n_1691;
wire n_1975;
wire n_1009;
wire n_1743;
wire n_1930;
wire n_1160;
wire n_883;
wire n_1238;
wire n_1991;
wire n_2179;
wire n_1724;
wire n_1032;
wire n_1247;
wire n_1547;
wire n_1553;
wire n_893;
wire n_1099;
wire n_1264;
wire n_1192;
wire n_471;
wire n_1844;
wire n_424;
wire n_1700;
wire n_1555;
wire n_1415;
wire n_2211;
wire n_1370;
wire n_1786;
wire n_369;
wire n_287;
wire n_2291;
wire n_415;
wire n_830;
wire n_230;
wire n_461;
wire n_873;
wire n_383;
wire n_1285;
wire n_1371;
wire n_1985;
wire n_447;
wire n_2184;
wire n_1803;
wire n_1172;
wire n_852;
wire n_1590;
wire n_1532;
wire n_1393;
wire n_1517;
wire n_1867;
wire n_1704;
wire n_1078;
wire n_250;
wire n_544;
wire n_1711;
wire n_2247;
wire n_1140;
wire n_1444;
wire n_1670;
wire n_1603;
wire n_1579;
wire n_1263;
wire n_2019;
wire n_836;
wire n_375;
wire n_2074;
wire n_522;
wire n_2129;
wire n_1261;
wire n_945;
wire n_2286;
wire n_1649;
wire n_2018;
wire n_2094;
wire n_1903;
wire n_1511;
wire n_1143;
wire n_1422;
wire n_1232;
wire n_1772;
wire n_1572;
wire n_616;
wire n_658;
wire n_1874;
wire n_1119;
wire n_2013;
wire n_428;
wire n_1433;
wire n_1902;
wire n_1842;
wire n_1620;
wire n_2044;
wire n_1954;
wire n_1735;
wire n_1541;
wire n_1300;
wire n_641;
wire n_822;
wire n_693;
wire n_1313;
wire n_1056;
wire n_2212;
wire n_758;
wire n_516;
wire n_1455;
wire n_1163;
wire n_1180;
wire n_2256;
wire n_943;
wire n_1798;
wire n_1550;
wire n_491;
wire n_1591;
wire n_772;
wire n_1344;
wire n_666;
wire n_371;
wire n_940;
wire n_770;
wire n_567;
wire n_1781;
wire n_1971;
wire n_2058;
wire n_2090;
wire n_405;
wire n_538;
wire n_2173;
wire n_2004;
wire n_1106;
wire n_886;
wire n_1471;
wire n_953;
wire n_343;
wire n_1094;
wire n_1345;
wire n_1820;
wire n_494;
wire n_539;
wire n_493;
wire n_2108;
wire n_454;
wire n_1421;
wire n_1936;
wire n_638;
wire n_1404;
wire n_1211;
wire n_2124;
wire n_381;
wire n_887;
wire n_1660;
wire n_1961;
wire n_1280;
wire n_713;
wire n_1400;
wire n_1467;
wire n_976;
wire n_2155;
wire n_1445;
wire n_1526;
wire n_1560;
wire n_734;
wire n_1088;
wire n_1894;
wire n_1231;
wire n_1978;
wire n_2085;
wire n_917;
wire n_574;
wire n_907;
wire n_1446;
wire n_659;
wire n_1815;
wire n_2214;
wire n_913;
wire n_407;
wire n_1658;
wire n_808;
wire n_867;
wire n_1230;
wire n_473;
wire n_1193;
wire n_1967;
wire n_1054;
wire n_559;
wire n_1333;
wire n_1648;
wire n_1911;
wire n_1956;
wire n_1644;
wire n_2011;
wire n_2277;
wire n_1558;
wire n_1732;
wire n_281;
wire n_551;
wire n_699;
wire n_1986;
wire n_564;
wire n_451;
wire n_824;
wire n_279;
wire n_686;
wire n_757;
wire n_594;
wire n_1641;
wire n_2113;
wire n_1918;
wire n_2190;
wire n_577;
wire n_1843;
wire n_619;
wire n_2268;
wire n_1367;
wire n_1336;
wire n_521;
wire n_572;
wire n_813;
wire n_395;
wire n_1909;
wire n_2080;
wire n_1481;
wire n_323;
wire n_606;
wire n_1441;
wire n_818;
wire n_1123;
wire n_1309;
wire n_2104;
wire n_513;
wire n_645;
wire n_1381;
wire n_331;
wire n_1699;
wire n_916;
wire n_2093;
wire n_483;
wire n_2207;
wire n_1970;
wire n_608;
wire n_261;
wire n_2101;
wire n_630;
wire n_2059;
wire n_2198;
wire n_541;
wire n_512;
wire n_2073;
wire n_2273;
wire n_433;
wire n_792;
wire n_476;
wire n_1328;
wire n_1957;
wire n_1907;
wire n_264;
wire n_263;
wire n_1162;
wire n_860;
wire n_1530;
wire n_788;
wire n_939;
wire n_1543;
wire n_821;
wire n_938;
wire n_1302;
wire n_1068;
wire n_1599;
wire n_329;
wire n_982;
wire n_549;
wire n_1762;
wire n_1910;
wire n_1075;
wire n_408;
wire n_932;
wire n_237;
wire n_1876;
wire n_1895;
wire n_2123;
wire n_1697;
wire n_2143;
wire n_243;
wire n_979;
wire n_1873;
wire n_905;
wire n_1866;
wire n_1680;
wire n_322;
wire n_993;
wire n_689;
wire n_2031;
wire n_354;
wire n_2130;
wire n_1330;
wire n_1413;
wire n_1605;
wire n_2228;
wire n_1988;
wire n_1278;
wire n_547;
wire n_558;
wire n_1064;
wire n_1396;
wire n_634;
wire n_966;
wire n_764;
wire n_1663;
wire n_2009;
wire n_692;
wire n_733;
wire n_1793;
wire n_1233;
wire n_1289;
wire n_2245;
wire n_487;
wire n_241;
wire n_2068;
wire n_1107;
wire n_1014;
wire n_1290;
wire n_1703;
wire n_882;
wire n_2176;
wire n_2072;
wire n_1354;
wire n_586;
wire n_423;
wire n_1865;
wire n_1875;
wire n_1701;
wire n_318;
wire n_1111;
wire n_1713;
wire n_715;
wire n_1251;
wire n_1265;
wire n_1726;
wire n_1950;
wire n_530;
wire n_1563;
wire n_1912;
wire n_277;
wire n_1982;
wire n_618;
wire n_1297;
wire n_1662;
wire n_1312;
wire n_1167;
wire n_1359;
wire n_674;
wire n_871;
wire n_922;
wire n_268;
wire n_1335;
wire n_1760;
wire n_1927;
wire n_2028;
wire n_1069;
wire n_1664;
wire n_1722;
wire n_612;
wire n_247;
wire n_1165;
wire n_355;
wire n_702;
wire n_347;
wire n_2008;
wire n_2192;
wire n_2254;
wire n_1926;
wire n_1175;
wire n_328;
wire n_1386;
wire n_1896;
wire n_429;
wire n_1747;
wire n_1012;
wire n_780;
wire n_675;
wire n_903;
wire n_1540;
wire n_1977;
wire n_1802;
wire n_1504;
wire n_286;
wire n_254;
wire n_2193;
wire n_1655;
wire n_242;
wire n_835;
wire n_928;
wire n_1214;
wire n_690;
wire n_850;
wire n_1801;
wire n_1886;
wire n_2092;
wire n_1654;
wire n_816;
wire n_1157;
wire n_1750;
wire n_1462;
wire n_1188;
wire n_1752;
wire n_877;
wire n_1813;
wire n_2206;
wire n_604;
wire n_825;
wire n_728;
wire n_1063;
wire n_1588;
wire n_267;
wire n_1124;
wire n_1624;
wire n_515;
wire n_2096;
wire n_1965;
wire n_598;
wire n_696;
wire n_1515;
wire n_961;
wire n_437;
wire n_1082;
wire n_1317;
wire n_593;
wire n_514;
wire n_687;
wire n_697;
wire n_890;
wire n_637;
wire n_295;
wire n_701;
wire n_2178;
wire n_950;
wire n_388;
wire n_484;
wire n_2036;
wire n_2152;
wire n_1709;
wire n_1825;
wire n_1757;
wire n_1796;
wire n_1792;
wire n_891;
wire n_2067;
wire n_2136;
wire n_2082;
wire n_2252;
wire n_1412;
wire n_949;
wire n_1630;
wire n_678;
wire n_283;
wire n_2075;
wire n_2194;
wire n_1987;
wire n_507;
wire n_968;
wire n_909;
wire n_1369;
wire n_881;
wire n_2271;
wire n_1008;
wire n_760;
wire n_1546;
wire n_590;
wire n_362;
wire n_2279;
wire n_462;
wire n_1033;
wire n_1052;
wire n_1296;
wire n_1990;
wire n_304;
wire n_694;
wire n_2150;
wire n_1294;
wire n_1420;
wire n_1634;
wire n_2078;
wire n_297;
wire n_627;
wire n_595;
wire n_1767;
wire n_1779;
wire n_524;
wire n_1465;
wire n_342;
wire n_1858;
wire n_1044;
wire n_2165;
wire n_2133;
wire n_1712;
wire n_1391;
wire n_449;
wire n_1523;
wire n_1208;
wire n_1164;
wire n_1295;
wire n_1627;
wire n_1072;
wire n_1527;
wire n_1495;
wire n_1438;
wire n_495;
wire n_815;
wire n_1100;
wire n_585;
wire n_1487;
wire n_840;
wire n_874;
wire n_1756;
wire n_1128;
wire n_673;
wire n_382;
wire n_2230;
wire n_1969;
wire n_1071;
wire n_1067;
wire n_1565;
wire n_1493;
wire n_2145;
wire n_1968;
wire n_898;
wire n_255;
wire n_284;
wire n_1952;
wire n_865;
wire n_925;
wire n_1932;
wire n_1101;
wire n_1026;
wire n_1880;
wire n_289;
wire n_1364;
wire n_615;
wire n_1249;
wire n_1293;
wire n_1127;
wire n_1512;
wire n_2151;
wire n_1451;
wire n_320;
wire n_639;
wire n_963;
wire n_794;
wire n_727;
wire n_894;
wire n_1839;
wire n_685;
wire n_1765;
wire n_353;
wire n_605;
wire n_1514;
wire n_1863;
wire n_826;
wire n_1646;
wire n_872;
wire n_1139;
wire n_1714;
wire n_718;
wire n_1018;
wire n_1521;
wire n_1366;
wire n_542;
wire n_847;
wire n_851;
wire n_682;
wire n_644;
wire n_305;
wire n_996;
wire n_532;
wire n_1308;
wire n_2089;
wire n_1376;
wire n_1513;
wire n_413;
wire n_791;
wire n_1913;
wire n_510;
wire n_837;
wire n_2097;
wire n_2170;
wire n_1488;
wire n_1808;
wire n_948;
wire n_704;
wire n_2148;
wire n_977;
wire n_1005;
wire n_1947;
wire n_536;
wire n_1788;
wire n_1999;
wire n_622;
wire n_1469;
wire n_2060;
wire n_1838;
wire n_1835;
wire n_1766;
wire n_1776;
wire n_1959;
wire n_2002;
wire n_581;
wire n_2138;
wire n_765;
wire n_432;
wire n_987;
wire n_1492;
wire n_1340;
wire n_1771;
wire n_631;
wire n_720;
wire n_842;
wire n_2262;
wire n_1707;
wire n_2239;
wire n_1432;
wire n_2208;
wire n_843;
wire n_656;
wire n_989;
wire n_1277;
wire n_797;
wire n_1473;
wire n_2191;
wire n_1723;
wire n_1246;
wire n_1878;
wire n_899;
wire n_738;
wire n_2012;
wire n_1304;
wire n_1035;
wire n_294;
wire n_499;
wire n_1426;
wire n_705;
wire n_1004;
wire n_1176;
wire n_2134;
wire n_1529;
wire n_1022;
wire n_614;
wire n_529;
wire n_2069;
wire n_425;
wire n_684;
wire n_1431;
wire n_1615;
wire n_1474;
wire n_1571;
wire n_1809;
wire n_1577;
wire n_2297;
wire n_1181;
wire n_2119;
wire n_1822;
wire n_486;
wire n_947;
wire n_1117;
wire n_1087;
wire n_1448;
wire n_1992;
wire n_648;
wire n_657;
wire n_1049;
wire n_2057;
wire n_2103;
wire n_1666;
wire n_1505;
wire n_803;
wire n_290;
wire n_1717;
wire n_926;
wire n_1817;
wire n_927;
wire n_1849;
wire n_919;
wire n_1698;
wire n_478;
wire n_2231;
wire n_929;
wire n_1228;
wire n_417;
wire n_446;
wire n_1568;
wire n_1490;
wire n_777;
wire n_1299;
wire n_272;
wire n_526;
wire n_1183;
wire n_1436;
wire n_2251;
wire n_1384;
wire n_2238;
wire n_293;
wire n_458;
wire n_1070;
wire n_998;
wire n_717;
wire n_1665;
wire n_1383;
wire n_1178;
wire n_2127;
wire n_1424;
wire n_1073;
wire n_1000;
wire n_796;
wire n_252;
wire n_1195;
wire n_2137;
wire n_1626;
wire n_1507;
wire n_552;
wire n_1358;
wire n_1811;
wire n_1388;
wire n_912;
wire n_1857;
wire n_1519;
wire n_2144;
wire n_745;
wire n_1284;
wire n_1604;
wire n_2296;
wire n_1142;
wire n_716;
wire n_1475;
wire n_623;
wire n_1048;
wire n_1201;
wire n_1398;
wire n_884;
wire n_1774;
wire n_1395;
wire n_2110;
wire n_2199;
wire n_731;
wire n_1502;
wire n_1659;
wire n_1955;
wire n_755;
wire n_931;
wire n_1021;
wire n_527;
wire n_474;
wire n_683;
wire n_811;
wire n_1207;
wire n_312;
wire n_1791;
wire n_1368;
wire n_1418;
wire n_958;
wire n_292;
wire n_1250;
wire n_1137;
wire n_1897;
wire n_2064;
wire n_880;
wire n_2053;
wire n_2259;
wire n_2121;
wire n_889;
wire n_1478;
wire n_589;
wire n_1310;
wire n_819;
wire n_2294;
wire n_1363;
wire n_1334;
wire n_1966;
wire n_1942;
wire n_767;
wire n_1314;
wire n_600;
wire n_964;
wire n_831;
wire n_1837;
wire n_2218;
wire n_477;
wire n_954;
wire n_864;
wire n_1110;
wire n_2213;
wire n_1410;
wire n_399;
wire n_1440;
wire n_2132;
wire n_2063;
wire n_1382;
wire n_1534;
wire n_1564;
wire n_1736;
wire n_1483;
wire n_1834;
wire n_1372;
wire n_231;
wire n_2292;
wire n_1457;
wire n_505;
wire n_1719;
wire n_319;
wire n_1339;
wire n_1787;
wire n_537;
wire n_1993;
wire n_2281;
wire n_1427;
wire n_311;
wire n_1466;
wire n_403;
wire n_1919;
wire n_1080;
wire n_723;
wire n_1877;
wire n_596;
wire n_546;
wire n_562;
wire n_1141;
wire n_1268;
wire n_386;
wire n_1939;
wire n_2030;
wire n_1769;
wire n_1220;
wire n_1893;
wire n_556;
wire n_2209;
wire n_1755;
wire n_1602;
wire n_1136;
wire n_2025;
wire n_1125;
wire n_970;
wire n_2224;
wire n_1980;
wire n_642;
wire n_995;
wire n_276;
wire n_1159;
wire n_1092;
wire n_2237;
wire n_441;
wire n_1060;
wire n_1951;
wire n_2250;
wire n_444;
wire n_1252;
wire n_1784;
wire n_1223;
wire n_303;
wire n_511;
wire n_1286;
wire n_1773;
wire n_1775;
wire n_2115;
wire n_1053;
wire n_416;
wire n_1681;
wire n_520;
wire n_418;
wire n_1093;
wire n_1783;
wire n_1533;
wire n_1597;
wire n_266;
wire n_296;
wire n_2274;
wire n_775;
wire n_651;
wire n_1153;
wire n_439;
wire n_1618;
wire n_518;
wire n_1531;
wire n_1185;
wire n_453;
wire n_1745;
wire n_914;
wire n_759;
wire n_1831;
wire n_426;
wire n_317;
wire n_1653;
wire n_1679;
wire n_1625;
wire n_2160;
wire n_1453;
wire n_2146;
wire n_2226;
wire n_2131;
wire n_488;
wire n_497;
wire n_773;
wire n_1901;
wire n_920;
wire n_1374;
wire n_1315;
wire n_1647;
wire n_1224;
wire n_1614;
wire n_1459;
wire n_1892;
wire n_1933;
wire n_1135;
wire n_1169;
wire n_1179;
wire n_401;
wire n_324;
wire n_1617;
wire n_335;
wire n_1470;
wire n_463;
wire n_1243;
wire n_848;
wire n_301;
wire n_274;
wire n_1096;
wire n_2249;
wire n_1091;
wire n_1917;
wire n_2000;
wire n_1580;
wire n_2227;
wire n_2270;
wire n_1425;
wire n_1881;
wire n_1281;
wire n_1267;
wire n_1806;
wire n_983;
wire n_2023;
wire n_427;
wire n_2204;
wire n_1520;
wire n_496;
wire n_2159;
wire n_906;
wire n_1390;
wire n_688;
wire n_2289;
wire n_1077;
wire n_1733;
wire n_1419;
wire n_351;
wire n_259;
wire n_1731;
wire n_2158;
wire n_2087;
wire n_1855;
wire n_1636;
wire n_1437;
wire n_2135;
wire n_1645;
wire n_1832;
wire n_385;
wire n_1687;
wire n_1439;
wire n_1323;
wire n_2202;
wire n_858;
wire n_2049;
wire n_1331;
wire n_736;
wire n_613;
wire n_501;
wire n_956;
wire n_960;
wire n_2276;
wire n_663;
wire n_856;
wire n_2100;
wire n_379;
wire n_778;
wire n_1668;
wire n_1134;
wire n_410;
wire n_1129;
wire n_554;
wire n_602;
wire n_1696;
wire n_1995;
wire n_1594;
wire n_2181;
wire n_664;
wire n_1869;
wire n_1764;
wire n_1429;
wire n_1610;
wire n_1889;
wire n_435;
wire n_1905;
wire n_2016;
wire n_793;
wire n_326;
wire n_587;
wire n_1593;
wire n_580;
wire n_762;
wire n_1030;
wire n_1202;
wire n_1937;
wire n_465;
wire n_1790;
wire n_1778;
wire n_1635;
wire n_1079;
wire n_341;
wire n_1744;
wire n_828;
wire n_2139;
wire n_2142;
wire n_607;
wire n_316;
wire n_419;
wire n_1551;
wire n_1103;
wire n_2219;
wire n_1203;
wire n_820;
wire n_951;
wire n_2201;
wire n_725;
wire n_952;
wire n_999;
wire n_358;
wire n_1254;
wire n_368;
wire n_575;
wire n_994;
wire n_2263;
wire n_1508;
wire n_732;
wire n_974;
wire n_2240;
wire n_392;
wire n_2278;
wire n_724;
wire n_1934;
wire n_1020;
wire n_1042;
wire n_628;
wire n_1273;
wire n_1434;
wire n_1573;
wire n_1728;
wire n_557;
wire n_1871;
wire n_349;
wire n_617;
wire n_845;
wire n_807;
wire n_1036;
wire n_1138;
wire n_1661;
wire n_1275;
wire n_485;
wire n_1549;
wire n_443;
wire n_1510;
wire n_892;
wire n_768;
wire n_421;
wire n_1468;
wire n_1859;
wire n_2102;
wire n_238;
wire n_1095;
wire n_2024;
wire n_1595;
wire n_2156;
wire n_1718;
wire n_1749;
wire n_1683;
wire n_1916;
wire n_597;
wire n_280;
wire n_1270;
wire n_1187;
wire n_610;
wire n_1403;
wire n_1669;
wire n_1852;
wire n_1024;
wire n_1768;
wire n_2153;
wire n_2052;
wire n_1847;
wire n_248;
wire n_517;
wire n_1667;
wire n_667;
wire n_1206;
wire n_621;
wire n_1037;
wire n_1397;
wire n_1279;
wire n_1115;
wire n_750;
wire n_901;
wire n_1499;
wire n_468;
wire n_923;
wire n_504;
wire n_1409;
wire n_1841;
wire n_1639;
wire n_1623;
wire n_1015;
wire n_1503;
wire n_466;
wire n_1057;
wire n_603;
wire n_991;
wire n_1657;
wire n_235;
wire n_1126;
wire n_1997;
wire n_340;
wire n_710;
wire n_1108;
wire n_1818;
wire n_1182;
wire n_1298;
wire n_2177;
wire n_2088;
wire n_1611;
wire n_785;
wire n_746;
wire n_609;
wire n_1601;
wire n_1960;
wire n_2061;
wire n_1686;
wire n_1356;
wire n_1589;
wire n_1740;
wire n_1497;
wire n_1168;
wire n_1216;
wire n_1943;
wire n_1320;
wire n_1430;
wire n_1316;
wire n_1287;
wire n_1452;
wire n_1622;
wire n_1586;
wire n_2264;
wire n_302;
wire n_1694;
wire n_380;
wire n_1535;
wire n_1596;
wire n_1190;
wire n_1734;
wire n_397;
wire n_1983;
wire n_1938;
wire n_2220;
wire n_1262;
wire n_1891;
wire n_2171;
wire n_1213;
wire n_2235;
wire n_1350;
wire n_1673;
wire n_2232;
wire n_1715;
wire n_1443;
wire n_1272;
wire n_239;
wire n_2037;
wire n_2298;
wire n_782;
wire n_1539;
wire n_490;
wire n_809;
wire n_1043;
wire n_1797;
wire n_1608;
wire n_986;
wire n_2120;
wire n_1472;
wire n_2050;
wire n_2164;
wire n_2225;
wire n_1081;
wire n_402;
wire n_1870;
wire n_352;
wire n_1692;
wire n_800;
wire n_1084;
wire n_1171;
wire n_460;
wire n_2169;
wire n_1827;
wire n_1361;
wire n_1864;
wire n_2006;
wire n_1491;
wire n_2187;
wire n_662;
wire n_374;
wire n_1152;
wire n_1840;
wire n_1705;
wire n_450;
wire n_2244;
wire n_1684;
wire n_921;
wire n_1346;
wire n_711;
wire n_1642;
wire n_579;
wire n_1352;
wire n_937;
wire n_2257;
wire n_1682;
wire n_2017;
wire n_370;
wire n_1695;
wire n_1828;
wire n_2046;
wire n_2272;
wire n_2200;
wire n_650;
wire n_1046;
wire n_1940;
wire n_1979;
wire n_1145;
wire n_330;
wire n_1121;
wire n_1102;
wire n_1963;
wire n_972;
wire n_1405;
wire n_258;
wire n_1406;
wire n_456;
wire n_1332;
wire n_260;
wire n_313;
wire n_624;
wire n_962;
wire n_1041;
wire n_565;
wire n_356;
wire n_1569;
wire n_936;
wire n_1883;
wire n_1288;
wire n_1186;
wire n_1062;
wire n_885;
wire n_896;
wire n_2167;
wire n_2084;
wire n_654;
wire n_411;
wire n_1222;
wire n_599;
wire n_776;
wire n_321;
wire n_1823;
wire n_1974;
wire n_1720;
wire n_482;
wire n_934;
wire n_1637;
wire n_1407;
wire n_1795;
wire n_420;
wire n_1341;
wire n_394;
wire n_1456;
wire n_1845;
wire n_1489;
wire n_942;
wire n_1524;
wire n_543;
wire n_2229;
wire n_1964;
wire n_2288;
wire n_1920;
wire n_2099;
wire n_1496;
wire n_1271;
wire n_1545;
wire n_2007;
wire n_2039;
wire n_1946;
wire n_1355;
wire n_1225;
wire n_1544;
wire n_1485;
wire n_2258;
wire n_325;
wire n_1640;
wire n_804;
wire n_464;
wire n_1846;
wire n_533;
wire n_806;
wire n_959;
wire n_879;
wire n_584;
wire n_2141;
wire n_244;
wire n_1343;
wire n_1522;
wire n_548;
wire n_1782;
wire n_282;
wire n_1676;
wire n_833;
wire n_1830;
wire n_1567;
wire n_523;
wire n_1319;
wire n_707;
wire n_345;
wire n_1900;
wire n_799;
wire n_1548;
wire n_1155;
wire n_2196;
wire n_273;
wire n_1633;
wire n_2195;
wire n_787;
wire n_2172;
wire n_1416;
wire n_1528;
wire n_2293;
wire n_1146;
wire n_2021;
wire n_2114;
wire n_1086;
wire n_1066;
wire n_1948;
wire n_2125;
wire n_2026;
wire n_1282;
wire n_550;
wire n_275;
wire n_652;
wire n_2154;
wire n_560;
wire n_1906;
wire n_1484;
wire n_1321;
wire n_1241;
wire n_1672;
wire n_569;
wire n_1758;
wire n_2283;
wire n_1925;
wire n_737;
wire n_1318;
wire n_1914;
wire n_1235;
wire n_1229;
wire n_306;
wire n_1292;
wire n_1373;
wire n_2266;
wire n_346;
wire n_1029;
wire n_1447;
wire n_2056;
wire n_790;
wire n_1706;
wire n_1498;
wire n_1210;
wire n_299;
wire n_1248;
wire n_1556;
wire n_902;
wire n_333;
wire n_2189;
wire n_2246;
wire n_1047;
wire n_1984;
wire n_2236;
wire n_1385;
wire n_431;
wire n_459;
wire n_1269;
wire n_1931;
wire n_2083;
wire n_502;
wire n_672;
wire n_1257;
wire n_1751;
wire n_285;
wire n_1375;
wire n_1941;
wire n_2128;
wire n_655;
wire n_706;
wire n_1045;
wire n_1650;
wire n_786;
wire n_1794;
wire n_1236;
wire n_1962;
wire n_1559;
wire n_1725;
wire n_1928;
wire n_1872;
wire n_834;
wire n_743;
wire n_766;
wire n_430;
wire n_1741;
wire n_1325;
wire n_1002;
wire n_1746;
wire n_1949;
wire n_545;
wire n_489;
wire n_1804;
wire n_1727;
wire n_251;
wire n_1019;
wire n_636;
wire n_2054;
wire n_729;
wire n_876;
wire n_774;
wire n_1337;
wire n_660;
wire n_2062;
wire n_2041;
wire n_438;
wire n_1477;
wire n_1360;
wire n_1860;
wire n_1904;
wire n_1200;
wire n_2070;
wire n_479;
wire n_1607;
wire n_1353;
wire n_1777;
wire n_1908;
wire n_1454;
wire n_2126;
wire n_869;
wire n_1154;
wire n_1113;
wire n_1600;
wire n_2253;
wire n_646;
wire n_528;
wire n_391;
wire n_1098;
wire n_1329;
wire n_2045;
wire n_817;
wire n_2261;
wire n_2216;
wire n_2210;
wire n_262;
wire n_897;
wire n_846;
wire n_2066;
wire n_841;
wire n_1476;
wire n_1001;
wire n_508;
wire n_1800;
wire n_2241;
wire n_1050;
wire n_1411;
wire n_1463;
wire n_1177;
wire n_332;
wire n_1150;
wire n_1742;
wire n_1562;
wire n_1690;
wire n_398;
wire n_1191;
wire n_1826;
wire n_566;
wire n_1023;
wire n_1882;
wire n_1118;
wire n_1076;
wire n_1007;
wire n_1807;
wire n_1929;
wire n_1378;
wire n_855;
wire n_1592;
wire n_1759;
wire n_1814;
wire n_1631;
wire n_591;
wire n_1377;
wire n_1879;
wire n_256;
wire n_853;
wire n_440;
wire n_695;
wire n_1542;
wire n_875;
wire n_367;
wire n_680;
wire n_1678;
wire n_661;
wire n_1716;
wire n_278;
wire n_1256;
wire n_671;
wire n_1953;
wire n_933;
wire n_740;
wire n_703;
wire n_978;
wire n_384;
wire n_1976;
wire n_1291;
wire n_1217;
wire n_751;
wire n_749;
wire n_1824;
wire n_310;
wire n_1628;
wire n_1324;
wire n_1399;
wire n_2122;
wire n_2109;
wire n_1435;
wire n_969;
wire n_988;
wire n_2140;
wire n_1065;
wire n_1401;
wire n_1255;
wire n_568;
wire n_1516;
wire n_1536;
wire n_2186;
wire n_2163;
wire n_2029;
wire n_1204;
wire n_823;
wire n_1132;
wire n_643;
wire n_233;
wire n_698;
wire n_1074;
wire n_1394;
wire n_1327;
wire n_1326;
wire n_739;
wire n_400;
wire n_955;
wire n_337;
wire n_1379;
wire n_246;
wire n_1338;
wire n_1097;
wire n_935;
wire n_781;
wire n_789;
wire n_1554;
wire n_1130;
wire n_1810;
wire n_573;
wire n_769;
wire n_676;
wire n_327;
wire n_1120;
wire n_832;
wire n_1583;
wire n_1730;
wire n_2295;
wire n_555;
wire n_389;
wire n_814;
wire n_1643;
wire n_2020;
wire n_2269;
wire n_1729;
wire n_669;
wire n_2290;
wire n_2048;
wire n_300;
wire n_2005;
wire n_747;
wire n_1389;
wire n_1105;
wire n_721;
wire n_1461;
wire n_742;
wire n_535;
wire n_691;
wire n_372;
wire n_2076;
wire n_314;
wire n_1408;
wire n_378;
wire n_1196;
wire n_377;
wire n_1598;
wire n_863;
wire n_2175;
wire n_601;
wire n_2182;
wire n_338;
wire n_1283;
wire n_918;
wire n_748;
wire n_506;
wire n_1114;
wire n_1785;
wire n_763;
wire n_1147;
wire n_1848;
wire n_360;
wire n_1754;
wire n_2149;
wire n_1506;
wire n_1652;
wire n_1812;
wire n_957;
wire n_1994;
wire n_895;
wire n_866;
wire n_1227;
wire n_2284;
wire n_387;
wire n_2287;
wire n_452;
wire n_744;
wire n_971;
wire n_946;
wire n_344;
wire n_761;
wire n_1303;
wire n_1205;
wire n_1258;
wire n_1392;
wire n_1173;
wire n_1924;
wire n_525;
wire n_1677;
wire n_1116;
wire n_611;
wire n_1570;
wire n_1702;
wire n_1219;
wire n_1780;
wire n_1689;
wire n_2180;
wire n_1174;
wire n_1944;
wire n_1016;
wire n_1347;
wire n_795;
wire n_1501;
wire n_1221;
wire n_1245;
wire n_838;
wire n_647;
wire n_844;
wire n_448;
wire n_1017;
wire n_2117;
wire n_2234;
wire n_1083;
wire n_445;
wire n_1561;
wire n_930;
wire n_888;
wire n_2275;
wire n_1112;
wire n_2081;
wire n_2168;
wire n_234;
wire n_2022;
wire n_1945;
wire n_2203;
wire n_910;
wire n_1656;
wire n_1721;
wire n_1460;
wire n_911;
wire n_2112;
wire n_2255;
wire n_1464;
wire n_236;
wire n_653;
wire n_1737;
wire n_1414;
wire n_752;
wire n_908;
wire n_944;
wire n_2034;
wire n_576;
wire n_1028;
wire n_2106;
wire n_472;
wire n_270;
wire n_2265;
wire n_414;
wire n_1922;
wire n_563;
wire n_2032;
wire n_1011;
wire n_1566;
wire n_1215;
wire n_839;
wire n_708;
wire n_1973;
wire n_2267;
wire n_668;
wire n_626;
wire n_990;
wire n_1500;
wire n_779;
wire n_1537;
wire n_1821;
wire n_2205;
wire n_1104;
wire n_854;
wire n_1058;
wire n_498;
wire n_1122;
wire n_870;
wire n_904;
wire n_1253;
wire n_709;
wire n_1266;
wire n_366;
wire n_2242;
wire n_1509;
wire n_1693;
wire n_1109;
wire n_2222;
wire n_712;
wire n_348;
wire n_1276;
wire n_376;
wire n_2015;
wire n_2118;
wire n_2111;
wire n_390;
wire n_1148;
wire n_2188;
wire n_334;
wire n_1989;
wire n_1161;
wire n_1085;
wire n_232;
wire n_2014;
wire n_2042;
wire n_1239;
wire n_771;
wire n_1584;
wire n_470;
wire n_475;
wire n_924;
wire n_298;
wire n_1582;
wire n_492;
wire n_1149;
wire n_265;
wire n_1184;
wire n_719;
wire n_1972;
wire n_1525;
wire n_455;
wire n_1585;
wire n_1851;
wire n_363;
wire n_1799;
wire n_1090;
wire n_2147;
wire n_592;
wire n_1816;
wire n_1518;
wire n_829;
wire n_1156;
wire n_1362;
wire n_393;
wire n_984;
wire n_1829;
wire n_503;
wire n_2035;
wire n_1450;
wire n_1638;
wire n_868;
wire n_570;
wire n_859;
wire n_2033;
wire n_406;
wire n_735;
wire n_1789;
wire n_1770;
wire n_878;
wire n_620;
wire n_519;
wire n_307;
wire n_469;
wire n_1218;
wire n_500;
wire n_1482;
wire n_981;
wire n_714;
wire n_1349;
wire n_291;
wire n_1144;
wire n_2071;
wire n_357;
wire n_985;
wire n_2233;
wire n_481;
wire n_997;
wire n_1710;
wire n_2161;
wire n_1301;
wire n_802;
wire n_561;
wire n_980;
wire n_1306;
wire n_2010;
wire n_2282;
wire n_1651;
wire n_1198;
wire n_2047;
wire n_2095;
wire n_1609;
wire n_2174;
wire n_436;
wire n_409;
wire n_1244;
wire n_1685;
wire n_1763;
wire n_1998;
wire n_1574;
wire n_240;
wire n_756;
wire n_1619;
wire n_1981;
wire n_2285;
wire n_1606;
wire n_810;
wire n_1133;
wire n_635;
wire n_1194;
wire n_1051;
wire n_253;
wire n_1552;
wire n_583;
wire n_1996;
wire n_249;
wire n_1039;
wire n_1442;
wire n_1034;
wire n_2043;
wire n_1480;
wire n_1158;
wire n_2248;
wire n_754;
wire n_941;
wire n_975;
wire n_1031;
wire n_1305;
wire n_553;
wire n_849;
wire n_753;
wire n_1753;
wire n_467;
wire n_269;
wire n_359;
wire n_973;
wire n_1921;
wire n_1479;
wire n_1055;
wire n_1675;
wire n_2197;
wire n_2217;
wire n_582;
wire n_2065;
wire n_861;
wire n_857;
wire n_967;
wire n_571;
wire n_2215;
wire n_271;
wire n_404;
wire n_2001;
wire n_2107;
wire n_1884;
wire n_2040;
wire n_679;
wire n_633;
wire n_1170;
wire n_665;
wire n_1629;
wire n_2221;
wire n_588;
wire n_1260;
wire n_308;
wire n_309;
wire n_2055;
wire n_1819;
wire n_1010;
wire n_1040;
wire n_915;
wire n_632;
wire n_1166;
wire n_2038;
wire n_812;
wire n_1131;
wire n_1761;
wire n_534;
wire n_1578;
wire n_1006;
wire n_1861;
wire n_373;
wire n_1632;
wire n_1890;
wire n_1805;
wire n_257;
wire n_1557;
wire n_1888;
wire n_2280;
wire n_1833;
wire n_730;
wire n_1311;
wire n_1494;
wire n_670;
wire n_1850;
wire n_1898;
wire n_2162;
wire n_1868;
wire n_2079;
wire n_1089;
wire n_1887;
wire n_1587;
wire n_1365;
wire n_1417;
wire n_1242;
wire n_2086;
wire n_2185;
wire n_1836;
wire n_681;
wire n_1226;
wire n_1274;
wire n_1486;
wire n_2166;
wire n_412;
wire n_640;
wire n_1322;
wire n_965;
wire n_1899;
wire n_1428;
wire n_1616;
wire n_1576;
wire n_1856;
wire n_1862;
wire n_1958;
wire n_2077;
wire n_339;
wire n_784;
wire n_434;
wire n_315;
wire n_288;
wire n_1059;
wire n_1197;
wire n_422;
wire n_722;
wire n_862;
wire n_2105;
wire n_2098;
wire n_540;
wire n_1423;
wire n_1935;
wire n_2027;
wire n_457;
wire n_2223;
wire n_2091;
wire n_364;
wire n_1915;
wire n_629;
wire n_1621;
wire n_1748;
wire n_900;
wire n_1449;
wire n_531;
wire n_827;
wire n_361;
wire n_1025;
wire n_2116;
wire n_336;
wire n_1885;
wire n_1013;
wire n_1259;
wire n_2183;
wire n_1538;
wire n_649;
wire n_1612;
wire n_1240;

INVx1_ASAP7_75t_L g230 ( 
.A(n_138),
.Y(n_230)
);

CKINVDCx5p33_ASAP7_75t_R g231 ( 
.A(n_52),
.Y(n_231)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_126),
.Y(n_232)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_228),
.Y(n_233)
);

CKINVDCx5p33_ASAP7_75t_R g234 ( 
.A(n_30),
.Y(n_234)
);

CKINVDCx20_ASAP7_75t_R g235 ( 
.A(n_185),
.Y(n_235)
);

CKINVDCx5p33_ASAP7_75t_R g236 ( 
.A(n_107),
.Y(n_236)
);

CKINVDCx5p33_ASAP7_75t_R g237 ( 
.A(n_58),
.Y(n_237)
);

CKINVDCx5p33_ASAP7_75t_R g238 ( 
.A(n_85),
.Y(n_238)
);

CKINVDCx5p33_ASAP7_75t_R g239 ( 
.A(n_10),
.Y(n_239)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_207),
.Y(n_240)
);

CKINVDCx5p33_ASAP7_75t_R g241 ( 
.A(n_120),
.Y(n_241)
);

CKINVDCx5p33_ASAP7_75t_R g242 ( 
.A(n_95),
.Y(n_242)
);

CKINVDCx5p33_ASAP7_75t_R g243 ( 
.A(n_89),
.Y(n_243)
);

CKINVDCx5p33_ASAP7_75t_R g244 ( 
.A(n_49),
.Y(n_244)
);

INVx2_ASAP7_75t_L g245 ( 
.A(n_187),
.Y(n_245)
);

INVx2_ASAP7_75t_L g246 ( 
.A(n_83),
.Y(n_246)
);

INVx2_ASAP7_75t_L g247 ( 
.A(n_63),
.Y(n_247)
);

CKINVDCx20_ASAP7_75t_R g248 ( 
.A(n_48),
.Y(n_248)
);

CKINVDCx5p33_ASAP7_75t_R g249 ( 
.A(n_21),
.Y(n_249)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_28),
.Y(n_250)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_93),
.Y(n_251)
);

BUFx6f_ASAP7_75t_L g252 ( 
.A(n_151),
.Y(n_252)
);

CKINVDCx5p33_ASAP7_75t_R g253 ( 
.A(n_62),
.Y(n_253)
);

BUFx5_ASAP7_75t_L g254 ( 
.A(n_173),
.Y(n_254)
);

CKINVDCx5p33_ASAP7_75t_R g255 ( 
.A(n_216),
.Y(n_255)
);

CKINVDCx5p33_ASAP7_75t_R g256 ( 
.A(n_20),
.Y(n_256)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_145),
.Y(n_257)
);

CKINVDCx5p33_ASAP7_75t_R g258 ( 
.A(n_7),
.Y(n_258)
);

INVx1_ASAP7_75t_SL g259 ( 
.A(n_122),
.Y(n_259)
);

CKINVDCx5p33_ASAP7_75t_R g260 ( 
.A(n_104),
.Y(n_260)
);

CKINVDCx5p33_ASAP7_75t_R g261 ( 
.A(n_215),
.Y(n_261)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_188),
.Y(n_262)
);

CKINVDCx5p33_ASAP7_75t_R g263 ( 
.A(n_91),
.Y(n_263)
);

CKINVDCx20_ASAP7_75t_R g264 ( 
.A(n_5),
.Y(n_264)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_108),
.Y(n_265)
);

CKINVDCx16_ASAP7_75t_R g266 ( 
.A(n_190),
.Y(n_266)
);

CKINVDCx5p33_ASAP7_75t_R g267 ( 
.A(n_112),
.Y(n_267)
);

CKINVDCx5p33_ASAP7_75t_R g268 ( 
.A(n_118),
.Y(n_268)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_97),
.Y(n_269)
);

CKINVDCx5p33_ASAP7_75t_R g270 ( 
.A(n_103),
.Y(n_270)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_148),
.Y(n_271)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_87),
.Y(n_272)
);

CKINVDCx5p33_ASAP7_75t_R g273 ( 
.A(n_177),
.Y(n_273)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_149),
.Y(n_274)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_175),
.Y(n_275)
);

CKINVDCx5p33_ASAP7_75t_R g276 ( 
.A(n_17),
.Y(n_276)
);

CKINVDCx5p33_ASAP7_75t_R g277 ( 
.A(n_24),
.Y(n_277)
);

CKINVDCx20_ASAP7_75t_R g278 ( 
.A(n_152),
.Y(n_278)
);

CKINVDCx5p33_ASAP7_75t_R g279 ( 
.A(n_11),
.Y(n_279)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_181),
.Y(n_280)
);

INVx2_ASAP7_75t_L g281 ( 
.A(n_217),
.Y(n_281)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_159),
.Y(n_282)
);

CKINVDCx5p33_ASAP7_75t_R g283 ( 
.A(n_3),
.Y(n_283)
);

CKINVDCx5p33_ASAP7_75t_R g284 ( 
.A(n_130),
.Y(n_284)
);

BUFx6f_ASAP7_75t_L g285 ( 
.A(n_63),
.Y(n_285)
);

BUFx6f_ASAP7_75t_L g286 ( 
.A(n_227),
.Y(n_286)
);

CKINVDCx5p33_ASAP7_75t_R g287 ( 
.A(n_147),
.Y(n_287)
);

CKINVDCx5p33_ASAP7_75t_R g288 ( 
.A(n_72),
.Y(n_288)
);

CKINVDCx20_ASAP7_75t_R g289 ( 
.A(n_60),
.Y(n_289)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_74),
.Y(n_290)
);

CKINVDCx20_ASAP7_75t_R g291 ( 
.A(n_172),
.Y(n_291)
);

CKINVDCx5p33_ASAP7_75t_R g292 ( 
.A(n_77),
.Y(n_292)
);

CKINVDCx5p33_ASAP7_75t_R g293 ( 
.A(n_210),
.Y(n_293)
);

CKINVDCx5p33_ASAP7_75t_R g294 ( 
.A(n_22),
.Y(n_294)
);

HB1xp67_ASAP7_75t_L g295 ( 
.A(n_202),
.Y(n_295)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_110),
.Y(n_296)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_170),
.Y(n_297)
);

BUFx6f_ASAP7_75t_L g298 ( 
.A(n_85),
.Y(n_298)
);

CKINVDCx5p33_ASAP7_75t_R g299 ( 
.A(n_62),
.Y(n_299)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_33),
.Y(n_300)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_28),
.Y(n_301)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_10),
.Y(n_302)
);

CKINVDCx20_ASAP7_75t_R g303 ( 
.A(n_19),
.Y(n_303)
);

CKINVDCx5p33_ASAP7_75t_R g304 ( 
.A(n_15),
.Y(n_304)
);

CKINVDCx16_ASAP7_75t_R g305 ( 
.A(n_129),
.Y(n_305)
);

CKINVDCx5p33_ASAP7_75t_R g306 ( 
.A(n_2),
.Y(n_306)
);

CKINVDCx5p33_ASAP7_75t_R g307 ( 
.A(n_68),
.Y(n_307)
);

BUFx3_ASAP7_75t_L g308 ( 
.A(n_54),
.Y(n_308)
);

BUFx3_ASAP7_75t_L g309 ( 
.A(n_75),
.Y(n_309)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_213),
.Y(n_310)
);

CKINVDCx20_ASAP7_75t_R g311 ( 
.A(n_226),
.Y(n_311)
);

CKINVDCx5p33_ASAP7_75t_R g312 ( 
.A(n_34),
.Y(n_312)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_30),
.Y(n_313)
);

CKINVDCx5p33_ASAP7_75t_R g314 ( 
.A(n_34),
.Y(n_314)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_195),
.Y(n_315)
);

CKINVDCx20_ASAP7_75t_R g316 ( 
.A(n_182),
.Y(n_316)
);

CKINVDCx5p33_ASAP7_75t_R g317 ( 
.A(n_154),
.Y(n_317)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_171),
.Y(n_318)
);

BUFx3_ASAP7_75t_L g319 ( 
.A(n_163),
.Y(n_319)
);

CKINVDCx5p33_ASAP7_75t_R g320 ( 
.A(n_65),
.Y(n_320)
);

CKINVDCx5p33_ASAP7_75t_R g321 ( 
.A(n_121),
.Y(n_321)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_123),
.Y(n_322)
);

CKINVDCx5p33_ASAP7_75t_R g323 ( 
.A(n_67),
.Y(n_323)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_39),
.Y(n_324)
);

INVx2_ASAP7_75t_SL g325 ( 
.A(n_11),
.Y(n_325)
);

CKINVDCx5p33_ASAP7_75t_R g326 ( 
.A(n_41),
.Y(n_326)
);

BUFx2_ASAP7_75t_L g327 ( 
.A(n_105),
.Y(n_327)
);

BUFx2_ASAP7_75t_L g328 ( 
.A(n_132),
.Y(n_328)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_183),
.Y(n_329)
);

CKINVDCx5p33_ASAP7_75t_R g330 ( 
.A(n_55),
.Y(n_330)
);

CKINVDCx5p33_ASAP7_75t_R g331 ( 
.A(n_113),
.Y(n_331)
);

CKINVDCx5p33_ASAP7_75t_R g332 ( 
.A(n_40),
.Y(n_332)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_75),
.Y(n_333)
);

INVx1_ASAP7_75t_SL g334 ( 
.A(n_117),
.Y(n_334)
);

CKINVDCx5p33_ASAP7_75t_R g335 ( 
.A(n_83),
.Y(n_335)
);

CKINVDCx5p33_ASAP7_75t_R g336 ( 
.A(n_86),
.Y(n_336)
);

CKINVDCx5p33_ASAP7_75t_R g337 ( 
.A(n_124),
.Y(n_337)
);

CKINVDCx5p33_ASAP7_75t_R g338 ( 
.A(n_78),
.Y(n_338)
);

BUFx5_ASAP7_75t_L g339 ( 
.A(n_37),
.Y(n_339)
);

CKINVDCx5p33_ASAP7_75t_R g340 ( 
.A(n_0),
.Y(n_340)
);

CKINVDCx5p33_ASAP7_75t_R g341 ( 
.A(n_204),
.Y(n_341)
);

CKINVDCx5p33_ASAP7_75t_R g342 ( 
.A(n_26),
.Y(n_342)
);

CKINVDCx5p33_ASAP7_75t_R g343 ( 
.A(n_38),
.Y(n_343)
);

CKINVDCx20_ASAP7_75t_R g344 ( 
.A(n_193),
.Y(n_344)
);

CKINVDCx20_ASAP7_75t_R g345 ( 
.A(n_92),
.Y(n_345)
);

CKINVDCx5p33_ASAP7_75t_R g346 ( 
.A(n_101),
.Y(n_346)
);

BUFx8_ASAP7_75t_SL g347 ( 
.A(n_100),
.Y(n_347)
);

INVx2_ASAP7_75t_L g348 ( 
.A(n_48),
.Y(n_348)
);

CKINVDCx5p33_ASAP7_75t_R g349 ( 
.A(n_20),
.Y(n_349)
);

CKINVDCx5p33_ASAP7_75t_R g350 ( 
.A(n_66),
.Y(n_350)
);

CKINVDCx5p33_ASAP7_75t_R g351 ( 
.A(n_19),
.Y(n_351)
);

INVx1_ASAP7_75t_L g352 ( 
.A(n_214),
.Y(n_352)
);

CKINVDCx20_ASAP7_75t_R g353 ( 
.A(n_12),
.Y(n_353)
);

CKINVDCx5p33_ASAP7_75t_R g354 ( 
.A(n_102),
.Y(n_354)
);

BUFx6f_ASAP7_75t_L g355 ( 
.A(n_144),
.Y(n_355)
);

CKINVDCx5p33_ASAP7_75t_R g356 ( 
.A(n_109),
.Y(n_356)
);

CKINVDCx5p33_ASAP7_75t_R g357 ( 
.A(n_79),
.Y(n_357)
);

CKINVDCx5p33_ASAP7_75t_R g358 ( 
.A(n_160),
.Y(n_358)
);

INVx1_ASAP7_75t_L g359 ( 
.A(n_225),
.Y(n_359)
);

CKINVDCx20_ASAP7_75t_R g360 ( 
.A(n_197),
.Y(n_360)
);

CKINVDCx20_ASAP7_75t_R g361 ( 
.A(n_31),
.Y(n_361)
);

INVx1_ASAP7_75t_L g362 ( 
.A(n_198),
.Y(n_362)
);

CKINVDCx5p33_ASAP7_75t_R g363 ( 
.A(n_51),
.Y(n_363)
);

CKINVDCx5p33_ASAP7_75t_R g364 ( 
.A(n_69),
.Y(n_364)
);

CKINVDCx5p33_ASAP7_75t_R g365 ( 
.A(n_40),
.Y(n_365)
);

BUFx10_ASAP7_75t_L g366 ( 
.A(n_199),
.Y(n_366)
);

CKINVDCx5p33_ASAP7_75t_R g367 ( 
.A(n_150),
.Y(n_367)
);

CKINVDCx20_ASAP7_75t_R g368 ( 
.A(n_99),
.Y(n_368)
);

CKINVDCx5p33_ASAP7_75t_R g369 ( 
.A(n_70),
.Y(n_369)
);

INVx1_ASAP7_75t_L g370 ( 
.A(n_51),
.Y(n_370)
);

INVx1_ASAP7_75t_L g371 ( 
.A(n_42),
.Y(n_371)
);

CKINVDCx5p33_ASAP7_75t_R g372 ( 
.A(n_3),
.Y(n_372)
);

CKINVDCx5p33_ASAP7_75t_R g373 ( 
.A(n_80),
.Y(n_373)
);

CKINVDCx5p33_ASAP7_75t_R g374 ( 
.A(n_142),
.Y(n_374)
);

INVx1_ASAP7_75t_L g375 ( 
.A(n_26),
.Y(n_375)
);

CKINVDCx20_ASAP7_75t_R g376 ( 
.A(n_164),
.Y(n_376)
);

CKINVDCx20_ASAP7_75t_R g377 ( 
.A(n_82),
.Y(n_377)
);

INVx1_ASAP7_75t_L g378 ( 
.A(n_12),
.Y(n_378)
);

INVx2_ASAP7_75t_SL g379 ( 
.A(n_128),
.Y(n_379)
);

CKINVDCx20_ASAP7_75t_R g380 ( 
.A(n_9),
.Y(n_380)
);

INVx1_ASAP7_75t_L g381 ( 
.A(n_201),
.Y(n_381)
);

CKINVDCx5p33_ASAP7_75t_R g382 ( 
.A(n_55),
.Y(n_382)
);

CKINVDCx5p33_ASAP7_75t_R g383 ( 
.A(n_169),
.Y(n_383)
);

CKINVDCx20_ASAP7_75t_R g384 ( 
.A(n_88),
.Y(n_384)
);

CKINVDCx5p33_ASAP7_75t_R g385 ( 
.A(n_24),
.Y(n_385)
);

INVx1_ASAP7_75t_L g386 ( 
.A(n_156),
.Y(n_386)
);

INVx1_ASAP7_75t_L g387 ( 
.A(n_29),
.Y(n_387)
);

CKINVDCx5p33_ASAP7_75t_R g388 ( 
.A(n_178),
.Y(n_388)
);

INVx2_ASAP7_75t_L g389 ( 
.A(n_168),
.Y(n_389)
);

INVx1_ASAP7_75t_L g390 ( 
.A(n_71),
.Y(n_390)
);

INVx1_ASAP7_75t_L g391 ( 
.A(n_52),
.Y(n_391)
);

CKINVDCx5p33_ASAP7_75t_R g392 ( 
.A(n_179),
.Y(n_392)
);

INVx1_ASAP7_75t_L g393 ( 
.A(n_131),
.Y(n_393)
);

CKINVDCx5p33_ASAP7_75t_R g394 ( 
.A(n_73),
.Y(n_394)
);

CKINVDCx5p33_ASAP7_75t_R g395 ( 
.A(n_15),
.Y(n_395)
);

CKINVDCx5p33_ASAP7_75t_R g396 ( 
.A(n_23),
.Y(n_396)
);

CKINVDCx5p33_ASAP7_75t_R g397 ( 
.A(n_134),
.Y(n_397)
);

INVx1_ASAP7_75t_L g398 ( 
.A(n_66),
.Y(n_398)
);

BUFx3_ASAP7_75t_L g399 ( 
.A(n_65),
.Y(n_399)
);

BUFx2_ASAP7_75t_L g400 ( 
.A(n_115),
.Y(n_400)
);

CKINVDCx5p33_ASAP7_75t_R g401 ( 
.A(n_61),
.Y(n_401)
);

CKINVDCx5p33_ASAP7_75t_R g402 ( 
.A(n_16),
.Y(n_402)
);

CKINVDCx5p33_ASAP7_75t_R g403 ( 
.A(n_81),
.Y(n_403)
);

CKINVDCx5p33_ASAP7_75t_R g404 ( 
.A(n_54),
.Y(n_404)
);

CKINVDCx5p33_ASAP7_75t_R g405 ( 
.A(n_29),
.Y(n_405)
);

CKINVDCx5p33_ASAP7_75t_R g406 ( 
.A(n_5),
.Y(n_406)
);

CKINVDCx5p33_ASAP7_75t_R g407 ( 
.A(n_21),
.Y(n_407)
);

INVx1_ASAP7_75t_L g408 ( 
.A(n_139),
.Y(n_408)
);

CKINVDCx20_ASAP7_75t_R g409 ( 
.A(n_13),
.Y(n_409)
);

CKINVDCx20_ASAP7_75t_R g410 ( 
.A(n_44),
.Y(n_410)
);

BUFx6f_ASAP7_75t_L g411 ( 
.A(n_196),
.Y(n_411)
);

INVx3_ASAP7_75t_L g412 ( 
.A(n_98),
.Y(n_412)
);

BUFx6f_ASAP7_75t_L g413 ( 
.A(n_49),
.Y(n_413)
);

CKINVDCx5p33_ASAP7_75t_R g414 ( 
.A(n_96),
.Y(n_414)
);

INVx1_ASAP7_75t_L g415 ( 
.A(n_59),
.Y(n_415)
);

INVx1_ASAP7_75t_L g416 ( 
.A(n_184),
.Y(n_416)
);

CKINVDCx5p33_ASAP7_75t_R g417 ( 
.A(n_209),
.Y(n_417)
);

CKINVDCx12_ASAP7_75t_R g418 ( 
.A(n_167),
.Y(n_418)
);

INVx1_ASAP7_75t_L g419 ( 
.A(n_94),
.Y(n_419)
);

CKINVDCx5p33_ASAP7_75t_R g420 ( 
.A(n_17),
.Y(n_420)
);

CKINVDCx5p33_ASAP7_75t_R g421 ( 
.A(n_194),
.Y(n_421)
);

BUFx6f_ASAP7_75t_L g422 ( 
.A(n_44),
.Y(n_422)
);

CKINVDCx5p33_ASAP7_75t_R g423 ( 
.A(n_223),
.Y(n_423)
);

INVx1_ASAP7_75t_L g424 ( 
.A(n_219),
.Y(n_424)
);

CKINVDCx5p33_ASAP7_75t_R g425 ( 
.A(n_174),
.Y(n_425)
);

CKINVDCx20_ASAP7_75t_R g426 ( 
.A(n_191),
.Y(n_426)
);

BUFx6f_ASAP7_75t_L g427 ( 
.A(n_6),
.Y(n_427)
);

INVx2_ASAP7_75t_SL g428 ( 
.A(n_135),
.Y(n_428)
);

INVx1_ASAP7_75t_SL g429 ( 
.A(n_36),
.Y(n_429)
);

CKINVDCx5p33_ASAP7_75t_R g430 ( 
.A(n_8),
.Y(n_430)
);

CKINVDCx20_ASAP7_75t_R g431 ( 
.A(n_161),
.Y(n_431)
);

BUFx10_ASAP7_75t_L g432 ( 
.A(n_57),
.Y(n_432)
);

INVx1_ASAP7_75t_L g433 ( 
.A(n_56),
.Y(n_433)
);

CKINVDCx5p33_ASAP7_75t_R g434 ( 
.A(n_76),
.Y(n_434)
);

CKINVDCx5p33_ASAP7_75t_R g435 ( 
.A(n_218),
.Y(n_435)
);

INVx1_ASAP7_75t_L g436 ( 
.A(n_16),
.Y(n_436)
);

CKINVDCx5p33_ASAP7_75t_R g437 ( 
.A(n_111),
.Y(n_437)
);

CKINVDCx5p33_ASAP7_75t_R g438 ( 
.A(n_205),
.Y(n_438)
);

CKINVDCx5p33_ASAP7_75t_R g439 ( 
.A(n_176),
.Y(n_439)
);

CKINVDCx5p33_ASAP7_75t_R g440 ( 
.A(n_64),
.Y(n_440)
);

INVx1_ASAP7_75t_L g441 ( 
.A(n_90),
.Y(n_441)
);

INVx1_ASAP7_75t_SL g442 ( 
.A(n_206),
.Y(n_442)
);

CKINVDCx5p33_ASAP7_75t_R g443 ( 
.A(n_84),
.Y(n_443)
);

CKINVDCx20_ASAP7_75t_R g444 ( 
.A(n_36),
.Y(n_444)
);

CKINVDCx20_ASAP7_75t_R g445 ( 
.A(n_37),
.Y(n_445)
);

CKINVDCx5p33_ASAP7_75t_R g446 ( 
.A(n_189),
.Y(n_446)
);

INVx1_ASAP7_75t_L g447 ( 
.A(n_41),
.Y(n_447)
);

INVx1_ASAP7_75t_L g448 ( 
.A(n_106),
.Y(n_448)
);

INVx1_ASAP7_75t_L g449 ( 
.A(n_77),
.Y(n_449)
);

CKINVDCx5p33_ASAP7_75t_R g450 ( 
.A(n_155),
.Y(n_450)
);

HB1xp67_ASAP7_75t_L g451 ( 
.A(n_74),
.Y(n_451)
);

INVx1_ASAP7_75t_L g452 ( 
.A(n_339),
.Y(n_452)
);

INVx1_ASAP7_75t_L g453 ( 
.A(n_339),
.Y(n_453)
);

CKINVDCx20_ASAP7_75t_R g454 ( 
.A(n_235),
.Y(n_454)
);

INVx2_ASAP7_75t_L g455 ( 
.A(n_339),
.Y(n_455)
);

INVx1_ASAP7_75t_L g456 ( 
.A(n_339),
.Y(n_456)
);

INVxp67_ASAP7_75t_SL g457 ( 
.A(n_295),
.Y(n_457)
);

INVx1_ASAP7_75t_L g458 ( 
.A(n_339),
.Y(n_458)
);

INVxp67_ASAP7_75t_SL g459 ( 
.A(n_327),
.Y(n_459)
);

CKINVDCx5p33_ASAP7_75t_R g460 ( 
.A(n_347),
.Y(n_460)
);

NOR2xp67_ASAP7_75t_L g461 ( 
.A(n_412),
.B(n_0),
.Y(n_461)
);

CKINVDCx5p33_ASAP7_75t_R g462 ( 
.A(n_270),
.Y(n_462)
);

INVx1_ASAP7_75t_L g463 ( 
.A(n_339),
.Y(n_463)
);

CKINVDCx5p33_ASAP7_75t_R g464 ( 
.A(n_273),
.Y(n_464)
);

INVx1_ASAP7_75t_L g465 ( 
.A(n_339),
.Y(n_465)
);

CKINVDCx5p33_ASAP7_75t_R g466 ( 
.A(n_284),
.Y(n_466)
);

CKINVDCx20_ASAP7_75t_R g467 ( 
.A(n_278),
.Y(n_467)
);

CKINVDCx5p33_ASAP7_75t_R g468 ( 
.A(n_287),
.Y(n_468)
);

BUFx2_ASAP7_75t_L g469 ( 
.A(n_308),
.Y(n_469)
);

INVx1_ASAP7_75t_L g470 ( 
.A(n_339),
.Y(n_470)
);

CKINVDCx20_ASAP7_75t_R g471 ( 
.A(n_291),
.Y(n_471)
);

CKINVDCx20_ASAP7_75t_R g472 ( 
.A(n_311),
.Y(n_472)
);

CKINVDCx5p33_ASAP7_75t_R g473 ( 
.A(n_293),
.Y(n_473)
);

CKINVDCx5p33_ASAP7_75t_R g474 ( 
.A(n_317),
.Y(n_474)
);

NOR2xp33_ASAP7_75t_L g475 ( 
.A(n_328),
.B(n_1),
.Y(n_475)
);

CKINVDCx5p33_ASAP7_75t_R g476 ( 
.A(n_321),
.Y(n_476)
);

CKINVDCx5p33_ASAP7_75t_R g477 ( 
.A(n_331),
.Y(n_477)
);

INVx2_ASAP7_75t_L g478 ( 
.A(n_285),
.Y(n_478)
);

INVx1_ASAP7_75t_L g479 ( 
.A(n_285),
.Y(n_479)
);

INVx1_ASAP7_75t_L g480 ( 
.A(n_285),
.Y(n_480)
);

INVx1_ASAP7_75t_L g481 ( 
.A(n_285),
.Y(n_481)
);

CKINVDCx20_ASAP7_75t_R g482 ( 
.A(n_316),
.Y(n_482)
);

NOR2xp67_ASAP7_75t_L g483 ( 
.A(n_412),
.B(n_1),
.Y(n_483)
);

INVxp33_ASAP7_75t_SL g484 ( 
.A(n_451),
.Y(n_484)
);

INVx1_ASAP7_75t_L g485 ( 
.A(n_285),
.Y(n_485)
);

CKINVDCx5p33_ASAP7_75t_R g486 ( 
.A(n_336),
.Y(n_486)
);

INVx1_ASAP7_75t_L g487 ( 
.A(n_298),
.Y(n_487)
);

INVx1_ASAP7_75t_L g488 ( 
.A(n_298),
.Y(n_488)
);

INVx1_ASAP7_75t_L g489 ( 
.A(n_298),
.Y(n_489)
);

CKINVDCx5p33_ASAP7_75t_R g490 ( 
.A(n_337),
.Y(n_490)
);

CKINVDCx5p33_ASAP7_75t_R g491 ( 
.A(n_346),
.Y(n_491)
);

INVx1_ASAP7_75t_L g492 ( 
.A(n_308),
.Y(n_492)
);

INVx1_ASAP7_75t_L g493 ( 
.A(n_309),
.Y(n_493)
);

CKINVDCx5p33_ASAP7_75t_R g494 ( 
.A(n_354),
.Y(n_494)
);

NOR2xp33_ASAP7_75t_L g495 ( 
.A(n_400),
.B(n_2),
.Y(n_495)
);

CKINVDCx20_ASAP7_75t_R g496 ( 
.A(n_344),
.Y(n_496)
);

CKINVDCx20_ASAP7_75t_R g497 ( 
.A(n_345),
.Y(n_497)
);

INVx1_ASAP7_75t_L g498 ( 
.A(n_298),
.Y(n_498)
);

BUFx2_ASAP7_75t_SL g499 ( 
.A(n_379),
.Y(n_499)
);

BUFx3_ASAP7_75t_L g500 ( 
.A(n_319),
.Y(n_500)
);

INVx1_ASAP7_75t_L g501 ( 
.A(n_298),
.Y(n_501)
);

CKINVDCx20_ASAP7_75t_R g502 ( 
.A(n_360),
.Y(n_502)
);

NOR2xp33_ASAP7_75t_L g503 ( 
.A(n_379),
.B(n_4),
.Y(n_503)
);

HB1xp67_ASAP7_75t_L g504 ( 
.A(n_231),
.Y(n_504)
);

INVx1_ASAP7_75t_L g505 ( 
.A(n_413),
.Y(n_505)
);

INVx1_ASAP7_75t_L g506 ( 
.A(n_413),
.Y(n_506)
);

NOR2xp33_ASAP7_75t_R g507 ( 
.A(n_368),
.B(n_114),
.Y(n_507)
);

INVx1_ASAP7_75t_L g508 ( 
.A(n_413),
.Y(n_508)
);

HB1xp67_ASAP7_75t_L g509 ( 
.A(n_231),
.Y(n_509)
);

INVx1_ASAP7_75t_L g510 ( 
.A(n_413),
.Y(n_510)
);

INVx1_ASAP7_75t_L g511 ( 
.A(n_413),
.Y(n_511)
);

NOR2xp33_ASAP7_75t_L g512 ( 
.A(n_428),
.B(n_4),
.Y(n_512)
);

CKINVDCx20_ASAP7_75t_R g513 ( 
.A(n_376),
.Y(n_513)
);

INVx2_ASAP7_75t_L g514 ( 
.A(n_422),
.Y(n_514)
);

INVx1_ASAP7_75t_L g515 ( 
.A(n_422),
.Y(n_515)
);

BUFx2_ASAP7_75t_SL g516 ( 
.A(n_428),
.Y(n_516)
);

INVxp67_ASAP7_75t_L g517 ( 
.A(n_432),
.Y(n_517)
);

INVx1_ASAP7_75t_L g518 ( 
.A(n_422),
.Y(n_518)
);

CKINVDCx20_ASAP7_75t_R g519 ( 
.A(n_384),
.Y(n_519)
);

CKINVDCx20_ASAP7_75t_R g520 ( 
.A(n_426),
.Y(n_520)
);

INVx1_ASAP7_75t_L g521 ( 
.A(n_422),
.Y(n_521)
);

CKINVDCx20_ASAP7_75t_R g522 ( 
.A(n_431),
.Y(n_522)
);

INVx1_ASAP7_75t_L g523 ( 
.A(n_422),
.Y(n_523)
);

INVx1_ASAP7_75t_L g524 ( 
.A(n_427),
.Y(n_524)
);

BUFx6f_ASAP7_75t_L g525 ( 
.A(n_252),
.Y(n_525)
);

INVx1_ASAP7_75t_L g526 ( 
.A(n_427),
.Y(n_526)
);

NOR2xp33_ASAP7_75t_L g527 ( 
.A(n_412),
.B(n_6),
.Y(n_527)
);

CKINVDCx20_ASAP7_75t_R g528 ( 
.A(n_266),
.Y(n_528)
);

CKINVDCx5p33_ASAP7_75t_R g529 ( 
.A(n_356),
.Y(n_529)
);

CKINVDCx20_ASAP7_75t_R g530 ( 
.A(n_305),
.Y(n_530)
);

INVxp67_ASAP7_75t_L g531 ( 
.A(n_432),
.Y(n_531)
);

INVx1_ASAP7_75t_L g532 ( 
.A(n_427),
.Y(n_532)
);

NAND2xp5_ASAP7_75t_L g533 ( 
.A(n_245),
.B(n_7),
.Y(n_533)
);

CKINVDCx20_ASAP7_75t_R g534 ( 
.A(n_358),
.Y(n_534)
);

CKINVDCx5p33_ASAP7_75t_R g535 ( 
.A(n_367),
.Y(n_535)
);

INVx1_ASAP7_75t_L g536 ( 
.A(n_427),
.Y(n_536)
);

CKINVDCx16_ASAP7_75t_R g537 ( 
.A(n_432),
.Y(n_537)
);

INVx1_ASAP7_75t_L g538 ( 
.A(n_427),
.Y(n_538)
);

INVxp67_ASAP7_75t_L g539 ( 
.A(n_250),
.Y(n_539)
);

NAND2xp5_ASAP7_75t_L g540 ( 
.A(n_245),
.B(n_8),
.Y(n_540)
);

CKINVDCx5p33_ASAP7_75t_R g541 ( 
.A(n_374),
.Y(n_541)
);

CKINVDCx5p33_ASAP7_75t_R g542 ( 
.A(n_383),
.Y(n_542)
);

NAND2xp5_ASAP7_75t_L g543 ( 
.A(n_281),
.B(n_9),
.Y(n_543)
);

CKINVDCx5p33_ASAP7_75t_R g544 ( 
.A(n_388),
.Y(n_544)
);

CKINVDCx16_ASAP7_75t_R g545 ( 
.A(n_366),
.Y(n_545)
);

CKINVDCx5p33_ASAP7_75t_R g546 ( 
.A(n_392),
.Y(n_546)
);

CKINVDCx5p33_ASAP7_75t_R g547 ( 
.A(n_397),
.Y(n_547)
);

CKINVDCx5p33_ASAP7_75t_R g548 ( 
.A(n_276),
.Y(n_548)
);

CKINVDCx5p33_ASAP7_75t_R g549 ( 
.A(n_277),
.Y(n_549)
);

CKINVDCx20_ASAP7_75t_R g550 ( 
.A(n_418),
.Y(n_550)
);

INVx1_ASAP7_75t_L g551 ( 
.A(n_246),
.Y(n_551)
);

CKINVDCx5p33_ASAP7_75t_R g552 ( 
.A(n_279),
.Y(n_552)
);

NOR2xp33_ASAP7_75t_L g553 ( 
.A(n_281),
.B(n_13),
.Y(n_553)
);

CKINVDCx5p33_ASAP7_75t_R g554 ( 
.A(n_283),
.Y(n_554)
);

INVx1_ASAP7_75t_L g555 ( 
.A(n_246),
.Y(n_555)
);

CKINVDCx5p33_ASAP7_75t_R g556 ( 
.A(n_288),
.Y(n_556)
);

CKINVDCx5p33_ASAP7_75t_R g557 ( 
.A(n_292),
.Y(n_557)
);

BUFx3_ASAP7_75t_L g558 ( 
.A(n_319),
.Y(n_558)
);

INVx1_ASAP7_75t_L g559 ( 
.A(n_247),
.Y(n_559)
);

CKINVDCx20_ASAP7_75t_R g560 ( 
.A(n_236),
.Y(n_560)
);

INVx2_ASAP7_75t_L g561 ( 
.A(n_254),
.Y(n_561)
);

NOR2xp33_ASAP7_75t_L g562 ( 
.A(n_389),
.B(n_14),
.Y(n_562)
);

INVxp33_ASAP7_75t_SL g563 ( 
.A(n_234),
.Y(n_563)
);

CKINVDCx20_ASAP7_75t_R g564 ( 
.A(n_236),
.Y(n_564)
);

CKINVDCx20_ASAP7_75t_R g565 ( 
.A(n_241),
.Y(n_565)
);

INVx1_ASAP7_75t_L g566 ( 
.A(n_247),
.Y(n_566)
);

CKINVDCx20_ASAP7_75t_R g567 ( 
.A(n_241),
.Y(n_567)
);

INVx1_ASAP7_75t_L g568 ( 
.A(n_348),
.Y(n_568)
);

HB1xp67_ASAP7_75t_L g569 ( 
.A(n_234),
.Y(n_569)
);

INVxp67_ASAP7_75t_SL g570 ( 
.A(n_309),
.Y(n_570)
);

CKINVDCx5p33_ASAP7_75t_R g571 ( 
.A(n_294),
.Y(n_571)
);

INVx1_ASAP7_75t_L g572 ( 
.A(n_348),
.Y(n_572)
);

CKINVDCx5p33_ASAP7_75t_R g573 ( 
.A(n_299),
.Y(n_573)
);

BUFx2_ASAP7_75t_L g574 ( 
.A(n_548),
.Y(n_574)
);

INVx2_ASAP7_75t_L g575 ( 
.A(n_455),
.Y(n_575)
);

AND2x2_ASAP7_75t_L g576 ( 
.A(n_570),
.B(n_399),
.Y(n_576)
);

INVx3_ASAP7_75t_L g577 ( 
.A(n_525),
.Y(n_577)
);

INVx2_ASAP7_75t_L g578 ( 
.A(n_455),
.Y(n_578)
);

INVx1_ASAP7_75t_L g579 ( 
.A(n_479),
.Y(n_579)
);

INVx1_ASAP7_75t_L g580 ( 
.A(n_479),
.Y(n_580)
);

INVx1_ASAP7_75t_L g581 ( 
.A(n_480),
.Y(n_581)
);

INVx5_ASAP7_75t_L g582 ( 
.A(n_525),
.Y(n_582)
);

AND2x6_ASAP7_75t_L g583 ( 
.A(n_527),
.B(n_389),
.Y(n_583)
);

INVx3_ASAP7_75t_L g584 ( 
.A(n_525),
.Y(n_584)
);

INVx1_ASAP7_75t_L g585 ( 
.A(n_480),
.Y(n_585)
);

INVx1_ASAP7_75t_L g586 ( 
.A(n_481),
.Y(n_586)
);

INVx1_ASAP7_75t_L g587 ( 
.A(n_481),
.Y(n_587)
);

INVx1_ASAP7_75t_L g588 ( 
.A(n_485),
.Y(n_588)
);

INVx1_ASAP7_75t_L g589 ( 
.A(n_485),
.Y(n_589)
);

INVx2_ASAP7_75t_L g590 ( 
.A(n_452),
.Y(n_590)
);

NAND2xp5_ASAP7_75t_L g591 ( 
.A(n_503),
.B(n_242),
.Y(n_591)
);

INVx2_ASAP7_75t_L g592 ( 
.A(n_452),
.Y(n_592)
);

NAND2xp5_ASAP7_75t_L g593 ( 
.A(n_512),
.B(n_242),
.Y(n_593)
);

AND2x4_ASAP7_75t_L g594 ( 
.A(n_461),
.B(n_252),
.Y(n_594)
);

INVx1_ASAP7_75t_L g595 ( 
.A(n_487),
.Y(n_595)
);

NAND2xp5_ASAP7_75t_SL g596 ( 
.A(n_483),
.B(n_366),
.Y(n_596)
);

BUFx6f_ASAP7_75t_L g597 ( 
.A(n_525),
.Y(n_597)
);

INVx1_ASAP7_75t_L g598 ( 
.A(n_487),
.Y(n_598)
);

INVx2_ASAP7_75t_L g599 ( 
.A(n_453),
.Y(n_599)
);

INVx3_ASAP7_75t_L g600 ( 
.A(n_525),
.Y(n_600)
);

INVx1_ASAP7_75t_L g601 ( 
.A(n_488),
.Y(n_601)
);

BUFx6f_ASAP7_75t_L g602 ( 
.A(n_561),
.Y(n_602)
);

AND2x4_ASAP7_75t_L g603 ( 
.A(n_478),
.B(n_252),
.Y(n_603)
);

AND2x4_ASAP7_75t_L g604 ( 
.A(n_478),
.B(n_252),
.Y(n_604)
);

INVx1_ASAP7_75t_L g605 ( 
.A(n_488),
.Y(n_605)
);

INVx2_ASAP7_75t_L g606 ( 
.A(n_453),
.Y(n_606)
);

BUFx6f_ASAP7_75t_L g607 ( 
.A(n_561),
.Y(n_607)
);

INVx3_ASAP7_75t_L g608 ( 
.A(n_514),
.Y(n_608)
);

NOR2xp33_ASAP7_75t_L g609 ( 
.A(n_499),
.B(n_259),
.Y(n_609)
);

INVx3_ASAP7_75t_L g610 ( 
.A(n_514),
.Y(n_610)
);

INVx1_ASAP7_75t_L g611 ( 
.A(n_489),
.Y(n_611)
);

AND2x2_ASAP7_75t_L g612 ( 
.A(n_500),
.B(n_399),
.Y(n_612)
);

INVx1_ASAP7_75t_L g613 ( 
.A(n_489),
.Y(n_613)
);

HB1xp67_ASAP7_75t_L g614 ( 
.A(n_504),
.Y(n_614)
);

NAND2xp5_ASAP7_75t_L g615 ( 
.A(n_498),
.B(n_501),
.Y(n_615)
);

CKINVDCx20_ASAP7_75t_R g616 ( 
.A(n_454),
.Y(n_616)
);

INVx2_ASAP7_75t_L g617 ( 
.A(n_456),
.Y(n_617)
);

INVx1_ASAP7_75t_L g618 ( 
.A(n_498),
.Y(n_618)
);

NAND2xp5_ASAP7_75t_SL g619 ( 
.A(n_475),
.B(n_366),
.Y(n_619)
);

BUFx2_ASAP7_75t_L g620 ( 
.A(n_549),
.Y(n_620)
);

INVx1_ASAP7_75t_L g621 ( 
.A(n_501),
.Y(n_621)
);

INVx1_ASAP7_75t_L g622 ( 
.A(n_505),
.Y(n_622)
);

BUFx6f_ASAP7_75t_L g623 ( 
.A(n_456),
.Y(n_623)
);

BUFx6f_ASAP7_75t_L g624 ( 
.A(n_458),
.Y(n_624)
);

INVx2_ASAP7_75t_L g625 ( 
.A(n_458),
.Y(n_625)
);

NOR2xp33_ASAP7_75t_L g626 ( 
.A(n_499),
.B(n_334),
.Y(n_626)
);

INVx2_ASAP7_75t_L g627 ( 
.A(n_463),
.Y(n_627)
);

INVx1_ASAP7_75t_L g628 ( 
.A(n_505),
.Y(n_628)
);

AND2x4_ASAP7_75t_L g629 ( 
.A(n_506),
.B(n_252),
.Y(n_629)
);

INVx1_ASAP7_75t_L g630 ( 
.A(n_506),
.Y(n_630)
);

INVx1_ASAP7_75t_L g631 ( 
.A(n_508),
.Y(n_631)
);

BUFx3_ASAP7_75t_L g632 ( 
.A(n_508),
.Y(n_632)
);

INVx1_ASAP7_75t_SL g633 ( 
.A(n_560),
.Y(n_633)
);

INVx2_ASAP7_75t_L g634 ( 
.A(n_463),
.Y(n_634)
);

INVx1_ASAP7_75t_L g635 ( 
.A(n_510),
.Y(n_635)
);

AND2x4_ASAP7_75t_L g636 ( 
.A(n_510),
.B(n_286),
.Y(n_636)
);

INVx2_ASAP7_75t_L g637 ( 
.A(n_465),
.Y(n_637)
);

INVx1_ASAP7_75t_L g638 ( 
.A(n_511),
.Y(n_638)
);

OA21x2_ASAP7_75t_L g639 ( 
.A1(n_465),
.A2(n_300),
.B(n_290),
.Y(n_639)
);

AND2x2_ASAP7_75t_L g640 ( 
.A(n_500),
.B(n_325),
.Y(n_640)
);

NAND2xp5_ASAP7_75t_L g641 ( 
.A(n_511),
.B(n_243),
.Y(n_641)
);

INVx1_ASAP7_75t_L g642 ( 
.A(n_515),
.Y(n_642)
);

INVx1_ASAP7_75t_L g643 ( 
.A(n_515),
.Y(n_643)
);

INVx1_ASAP7_75t_L g644 ( 
.A(n_518),
.Y(n_644)
);

INVx1_ASAP7_75t_L g645 ( 
.A(n_518),
.Y(n_645)
);

BUFx3_ASAP7_75t_L g646 ( 
.A(n_521),
.Y(n_646)
);

INVx2_ASAP7_75t_L g647 ( 
.A(n_470),
.Y(n_647)
);

INVx1_ASAP7_75t_L g648 ( 
.A(n_521),
.Y(n_648)
);

INVx3_ASAP7_75t_L g649 ( 
.A(n_470),
.Y(n_649)
);

OAI21x1_ASAP7_75t_L g650 ( 
.A1(n_533),
.A2(n_232),
.B(n_230),
.Y(n_650)
);

INVx2_ASAP7_75t_L g651 ( 
.A(n_523),
.Y(n_651)
);

NAND2xp5_ASAP7_75t_L g652 ( 
.A(n_523),
.B(n_243),
.Y(n_652)
);

INVx3_ASAP7_75t_L g653 ( 
.A(n_524),
.Y(n_653)
);

INVx2_ASAP7_75t_L g654 ( 
.A(n_524),
.Y(n_654)
);

INVx3_ASAP7_75t_L g655 ( 
.A(n_526),
.Y(n_655)
);

INVx3_ASAP7_75t_L g656 ( 
.A(n_526),
.Y(n_656)
);

INVx1_ASAP7_75t_L g657 ( 
.A(n_532),
.Y(n_657)
);

INVx1_ASAP7_75t_L g658 ( 
.A(n_532),
.Y(n_658)
);

INVx1_ASAP7_75t_L g659 ( 
.A(n_536),
.Y(n_659)
);

OR2x6_ASAP7_75t_L g660 ( 
.A(n_540),
.B(n_325),
.Y(n_660)
);

INVx2_ASAP7_75t_L g661 ( 
.A(n_536),
.Y(n_661)
);

INVx1_ASAP7_75t_L g662 ( 
.A(n_538),
.Y(n_662)
);

INVx1_ASAP7_75t_L g663 ( 
.A(n_538),
.Y(n_663)
);

INVx1_ASAP7_75t_L g664 ( 
.A(n_551),
.Y(n_664)
);

INVx1_ASAP7_75t_L g665 ( 
.A(n_551),
.Y(n_665)
);

AND2x2_ASAP7_75t_L g666 ( 
.A(n_558),
.B(n_233),
.Y(n_666)
);

INVx1_ASAP7_75t_L g667 ( 
.A(n_555),
.Y(n_667)
);

BUFx6f_ASAP7_75t_L g668 ( 
.A(n_555),
.Y(n_668)
);

INVx2_ASAP7_75t_L g669 ( 
.A(n_575),
.Y(n_669)
);

INVx1_ASAP7_75t_L g670 ( 
.A(n_632),
.Y(n_670)
);

NAND2xp5_ASAP7_75t_L g671 ( 
.A(n_609),
.B(n_462),
.Y(n_671)
);

INVxp33_ASAP7_75t_L g672 ( 
.A(n_612),
.Y(n_672)
);

BUFx2_ASAP7_75t_L g673 ( 
.A(n_574),
.Y(n_673)
);

NOR2xp33_ASAP7_75t_L g674 ( 
.A(n_619),
.B(n_464),
.Y(n_674)
);

INVx2_ASAP7_75t_L g675 ( 
.A(n_575),
.Y(n_675)
);

INVx1_ASAP7_75t_L g676 ( 
.A(n_632),
.Y(n_676)
);

INVx1_ASAP7_75t_L g677 ( 
.A(n_632),
.Y(n_677)
);

NAND2xp5_ASAP7_75t_L g678 ( 
.A(n_609),
.B(n_466),
.Y(n_678)
);

INVx2_ASAP7_75t_L g679 ( 
.A(n_575),
.Y(n_679)
);

NOR2xp33_ASAP7_75t_L g680 ( 
.A(n_619),
.B(n_468),
.Y(n_680)
);

NOR2xp33_ASAP7_75t_L g681 ( 
.A(n_591),
.B(n_473),
.Y(n_681)
);

INVx1_ASAP7_75t_L g682 ( 
.A(n_632),
.Y(n_682)
);

CKINVDCx8_ASAP7_75t_R g683 ( 
.A(n_574),
.Y(n_683)
);

AND2x2_ASAP7_75t_L g684 ( 
.A(n_666),
.B(n_558),
.Y(n_684)
);

INVx1_ASAP7_75t_L g685 ( 
.A(n_646),
.Y(n_685)
);

INVx2_ASAP7_75t_SL g686 ( 
.A(n_612),
.Y(n_686)
);

CKINVDCx5p33_ASAP7_75t_R g687 ( 
.A(n_616),
.Y(n_687)
);

BUFx2_ASAP7_75t_L g688 ( 
.A(n_574),
.Y(n_688)
);

INVx1_ASAP7_75t_L g689 ( 
.A(n_646),
.Y(n_689)
);

NAND2xp5_ASAP7_75t_L g690 ( 
.A(n_626),
.B(n_474),
.Y(n_690)
);

INVx1_ASAP7_75t_L g691 ( 
.A(n_646),
.Y(n_691)
);

INVx1_ASAP7_75t_L g692 ( 
.A(n_646),
.Y(n_692)
);

NAND2xp33_ASAP7_75t_R g693 ( 
.A(n_620),
.B(n_552),
.Y(n_693)
);

INVxp67_ASAP7_75t_SL g694 ( 
.A(n_602),
.Y(n_694)
);

INVx3_ASAP7_75t_L g695 ( 
.A(n_597),
.Y(n_695)
);

OR2x2_ASAP7_75t_L g696 ( 
.A(n_614),
.B(n_509),
.Y(n_696)
);

INVx4_ASAP7_75t_L g697 ( 
.A(n_623),
.Y(n_697)
);

OR2x6_ASAP7_75t_L g698 ( 
.A(n_660),
.B(n_539),
.Y(n_698)
);

AOI22xp5_ASAP7_75t_L g699 ( 
.A1(n_626),
.A2(n_459),
.B1(n_534),
.B2(n_457),
.Y(n_699)
);

INVx1_ASAP7_75t_SL g700 ( 
.A(n_633),
.Y(n_700)
);

NOR2xp33_ASAP7_75t_L g701 ( 
.A(n_591),
.B(n_476),
.Y(n_701)
);

INVx2_ASAP7_75t_L g702 ( 
.A(n_575),
.Y(n_702)
);

BUFx6f_ASAP7_75t_L g703 ( 
.A(n_597),
.Y(n_703)
);

AOI22xp5_ASAP7_75t_L g704 ( 
.A1(n_576),
.A2(n_565),
.B1(n_567),
.B2(n_564),
.Y(n_704)
);

INVx1_ASAP7_75t_L g705 ( 
.A(n_649),
.Y(n_705)
);

AND2x6_ASAP7_75t_L g706 ( 
.A(n_594),
.B(n_286),
.Y(n_706)
);

AND2x6_ASAP7_75t_L g707 ( 
.A(n_594),
.B(n_286),
.Y(n_707)
);

NOR2xp33_ASAP7_75t_L g708 ( 
.A(n_593),
.B(n_477),
.Y(n_708)
);

INVx2_ASAP7_75t_L g709 ( 
.A(n_578),
.Y(n_709)
);

AOI22xp5_ASAP7_75t_L g710 ( 
.A1(n_576),
.A2(n_554),
.B1(n_557),
.B2(n_556),
.Y(n_710)
);

INVx3_ASAP7_75t_L g711 ( 
.A(n_597),
.Y(n_711)
);

INVx2_ASAP7_75t_L g712 ( 
.A(n_578),
.Y(n_712)
);

INVx1_ASAP7_75t_L g713 ( 
.A(n_649),
.Y(n_713)
);

NAND2xp5_ASAP7_75t_L g714 ( 
.A(n_593),
.B(n_486),
.Y(n_714)
);

INVx2_ASAP7_75t_L g715 ( 
.A(n_578),
.Y(n_715)
);

INVx1_ASAP7_75t_L g716 ( 
.A(n_649),
.Y(n_716)
);

INVx2_ASAP7_75t_L g717 ( 
.A(n_578),
.Y(n_717)
);

CKINVDCx5p33_ASAP7_75t_R g718 ( 
.A(n_616),
.Y(n_718)
);

INVx1_ASAP7_75t_L g719 ( 
.A(n_649),
.Y(n_719)
);

INVx2_ASAP7_75t_L g720 ( 
.A(n_651),
.Y(n_720)
);

INVx1_ASAP7_75t_L g721 ( 
.A(n_649),
.Y(n_721)
);

NAND2xp5_ASAP7_75t_SL g722 ( 
.A(n_594),
.B(n_571),
.Y(n_722)
);

INVx2_ASAP7_75t_L g723 ( 
.A(n_651),
.Y(n_723)
);

NOR2x1p5_ASAP7_75t_L g724 ( 
.A(n_640),
.B(n_460),
.Y(n_724)
);

INVxp33_ASAP7_75t_L g725 ( 
.A(n_612),
.Y(n_725)
);

INVx1_ASAP7_75t_L g726 ( 
.A(n_639),
.Y(n_726)
);

INVx2_ASAP7_75t_L g727 ( 
.A(n_651),
.Y(n_727)
);

AND2x4_ASAP7_75t_L g728 ( 
.A(n_666),
.B(n_492),
.Y(n_728)
);

INVx3_ASAP7_75t_L g729 ( 
.A(n_597),
.Y(n_729)
);

INVx4_ASAP7_75t_L g730 ( 
.A(n_623),
.Y(n_730)
);

INVx1_ASAP7_75t_L g731 ( 
.A(n_639),
.Y(n_731)
);

INVx2_ASAP7_75t_SL g732 ( 
.A(n_576),
.Y(n_732)
);

INVx1_ASAP7_75t_L g733 ( 
.A(n_639),
.Y(n_733)
);

NOR2xp33_ASAP7_75t_L g734 ( 
.A(n_596),
.B(n_490),
.Y(n_734)
);

INVx6_ASAP7_75t_L g735 ( 
.A(n_594),
.Y(n_735)
);

INVx2_ASAP7_75t_L g736 ( 
.A(n_651),
.Y(n_736)
);

NAND2xp5_ASAP7_75t_L g737 ( 
.A(n_583),
.B(n_491),
.Y(n_737)
);

INVx2_ASAP7_75t_L g738 ( 
.A(n_654),
.Y(n_738)
);

INVx3_ASAP7_75t_L g739 ( 
.A(n_597),
.Y(n_739)
);

AOI22xp33_ASAP7_75t_L g740 ( 
.A1(n_583),
.A2(n_553),
.B1(n_562),
.B2(n_484),
.Y(n_740)
);

INVx2_ASAP7_75t_L g741 ( 
.A(n_654),
.Y(n_741)
);

NAND2xp33_ASAP7_75t_L g742 ( 
.A(n_583),
.B(n_286),
.Y(n_742)
);

INVx2_ASAP7_75t_L g743 ( 
.A(n_654),
.Y(n_743)
);

NAND2xp5_ASAP7_75t_L g744 ( 
.A(n_583),
.B(n_494),
.Y(n_744)
);

INVx2_ASAP7_75t_L g745 ( 
.A(n_654),
.Y(n_745)
);

INVx1_ASAP7_75t_L g746 ( 
.A(n_639),
.Y(n_746)
);

NOR2xp33_ASAP7_75t_L g747 ( 
.A(n_596),
.B(n_529),
.Y(n_747)
);

INVx2_ASAP7_75t_L g748 ( 
.A(n_661),
.Y(n_748)
);

BUFx2_ASAP7_75t_L g749 ( 
.A(n_620),
.Y(n_749)
);

CKINVDCx5p33_ASAP7_75t_R g750 ( 
.A(n_633),
.Y(n_750)
);

NAND2xp5_ASAP7_75t_SL g751 ( 
.A(n_594),
.B(n_573),
.Y(n_751)
);

NOR2xp33_ASAP7_75t_L g752 ( 
.A(n_641),
.B(n_535),
.Y(n_752)
);

NAND3xp33_ASAP7_75t_L g753 ( 
.A(n_641),
.B(n_495),
.C(n_541),
.Y(n_753)
);

NOR2xp33_ASAP7_75t_L g754 ( 
.A(n_652),
.B(n_542),
.Y(n_754)
);

INVx1_ASAP7_75t_L g755 ( 
.A(n_639),
.Y(n_755)
);

INVx3_ASAP7_75t_L g756 ( 
.A(n_597),
.Y(n_756)
);

AND3x2_ASAP7_75t_L g757 ( 
.A(n_620),
.B(n_531),
.C(n_517),
.Y(n_757)
);

INVx3_ASAP7_75t_L g758 ( 
.A(n_597),
.Y(n_758)
);

NAND3xp33_ASAP7_75t_L g759 ( 
.A(n_652),
.B(n_546),
.C(n_544),
.Y(n_759)
);

INVxp67_ASAP7_75t_SL g760 ( 
.A(n_602),
.Y(n_760)
);

BUFx6f_ASAP7_75t_L g761 ( 
.A(n_597),
.Y(n_761)
);

AND2x2_ASAP7_75t_L g762 ( 
.A(n_666),
.B(n_516),
.Y(n_762)
);

NAND2xp5_ASAP7_75t_SL g763 ( 
.A(n_594),
.B(n_286),
.Y(n_763)
);

NAND2xp5_ASAP7_75t_SL g764 ( 
.A(n_629),
.B(n_355),
.Y(n_764)
);

OR2x2_ASAP7_75t_L g765 ( 
.A(n_614),
.B(n_569),
.Y(n_765)
);

INVxp67_ASAP7_75t_SL g766 ( 
.A(n_602),
.Y(n_766)
);

INVx1_ASAP7_75t_L g767 ( 
.A(n_639),
.Y(n_767)
);

NAND2xp5_ASAP7_75t_SL g768 ( 
.A(n_629),
.B(n_355),
.Y(n_768)
);

INVx5_ASAP7_75t_L g769 ( 
.A(n_583),
.Y(n_769)
);

INVx2_ASAP7_75t_L g770 ( 
.A(n_661),
.Y(n_770)
);

NAND2xp5_ASAP7_75t_SL g771 ( 
.A(n_629),
.B(n_355),
.Y(n_771)
);

INVx1_ASAP7_75t_L g772 ( 
.A(n_629),
.Y(n_772)
);

INVx2_ASAP7_75t_L g773 ( 
.A(n_661),
.Y(n_773)
);

INVx1_ASAP7_75t_L g774 ( 
.A(n_629),
.Y(n_774)
);

NOR2xp33_ASAP7_75t_L g775 ( 
.A(n_640),
.B(n_547),
.Y(n_775)
);

NAND2xp5_ASAP7_75t_SL g776 ( 
.A(n_636),
.B(n_355),
.Y(n_776)
);

INVx2_ASAP7_75t_L g777 ( 
.A(n_661),
.Y(n_777)
);

INVx1_ASAP7_75t_L g778 ( 
.A(n_636),
.Y(n_778)
);

INVx1_ASAP7_75t_L g779 ( 
.A(n_636),
.Y(n_779)
);

INVx2_ASAP7_75t_SL g780 ( 
.A(n_640),
.Y(n_780)
);

INVx5_ASAP7_75t_L g781 ( 
.A(n_583),
.Y(n_781)
);

NAND2xp33_ASAP7_75t_L g782 ( 
.A(n_583),
.B(n_355),
.Y(n_782)
);

AND2x2_ASAP7_75t_SL g783 ( 
.A(n_603),
.B(n_543),
.Y(n_783)
);

AND2x6_ASAP7_75t_L g784 ( 
.A(n_590),
.B(n_411),
.Y(n_784)
);

OR2x6_ASAP7_75t_L g785 ( 
.A(n_660),
.B(n_516),
.Y(n_785)
);

INVx4_ASAP7_75t_L g786 ( 
.A(n_623),
.Y(n_786)
);

AND2x2_ASAP7_75t_L g787 ( 
.A(n_664),
.B(n_493),
.Y(n_787)
);

INVx4_ASAP7_75t_SL g788 ( 
.A(n_583),
.Y(n_788)
);

INVx2_ASAP7_75t_SL g789 ( 
.A(n_660),
.Y(n_789)
);

INVx1_ASAP7_75t_L g790 ( 
.A(n_636),
.Y(n_790)
);

INVxp33_ASAP7_75t_L g791 ( 
.A(n_664),
.Y(n_791)
);

NOR2xp33_ASAP7_75t_L g792 ( 
.A(n_660),
.B(n_563),
.Y(n_792)
);

NAND2xp5_ASAP7_75t_SL g793 ( 
.A(n_636),
.B(n_411),
.Y(n_793)
);

INVx1_ASAP7_75t_L g794 ( 
.A(n_636),
.Y(n_794)
);

NOR2xp33_ASAP7_75t_L g795 ( 
.A(n_660),
.B(n_545),
.Y(n_795)
);

INVx1_ASAP7_75t_L g796 ( 
.A(n_603),
.Y(n_796)
);

INVx1_ASAP7_75t_L g797 ( 
.A(n_603),
.Y(n_797)
);

NAND3xp33_ASAP7_75t_L g798 ( 
.A(n_660),
.B(n_469),
.C(n_306),
.Y(n_798)
);

NAND3xp33_ASAP7_75t_L g799 ( 
.A(n_660),
.B(n_469),
.C(n_307),
.Y(n_799)
);

INVx2_ASAP7_75t_L g800 ( 
.A(n_590),
.Y(n_800)
);

INVx1_ASAP7_75t_L g801 ( 
.A(n_603),
.Y(n_801)
);

AND2x6_ASAP7_75t_L g802 ( 
.A(n_590),
.B(n_411),
.Y(n_802)
);

INVx4_ASAP7_75t_L g803 ( 
.A(n_623),
.Y(n_803)
);

OR2x6_ASAP7_75t_L g804 ( 
.A(n_650),
.B(n_301),
.Y(n_804)
);

INVx1_ASAP7_75t_L g805 ( 
.A(n_603),
.Y(n_805)
);

INVx2_ASAP7_75t_SL g806 ( 
.A(n_583),
.Y(n_806)
);

INVx2_ASAP7_75t_L g807 ( 
.A(n_590),
.Y(n_807)
);

NAND2xp5_ASAP7_75t_SL g808 ( 
.A(n_650),
.B(n_411),
.Y(n_808)
);

INVx2_ASAP7_75t_L g809 ( 
.A(n_592),
.Y(n_809)
);

INVx2_ASAP7_75t_L g810 ( 
.A(n_592),
.Y(n_810)
);

NAND2xp5_ASAP7_75t_L g811 ( 
.A(n_583),
.B(n_442),
.Y(n_811)
);

AND2x2_ASAP7_75t_L g812 ( 
.A(n_664),
.B(n_572),
.Y(n_812)
);

INVx1_ASAP7_75t_SL g813 ( 
.A(n_665),
.Y(n_813)
);

INVx6_ASAP7_75t_L g814 ( 
.A(n_603),
.Y(n_814)
);

HB1xp67_ASAP7_75t_L g815 ( 
.A(n_665),
.Y(n_815)
);

AOI22xp5_ASAP7_75t_L g816 ( 
.A1(n_583),
.A2(n_550),
.B1(n_530),
.B2(n_528),
.Y(n_816)
);

BUFx3_ASAP7_75t_L g817 ( 
.A(n_604),
.Y(n_817)
);

INVx2_ASAP7_75t_L g818 ( 
.A(n_592),
.Y(n_818)
);

NAND2xp5_ASAP7_75t_L g819 ( 
.A(n_592),
.B(n_240),
.Y(n_819)
);

AND2x2_ASAP7_75t_L g820 ( 
.A(n_665),
.B(n_572),
.Y(n_820)
);

NOR2xp33_ASAP7_75t_L g821 ( 
.A(n_667),
.B(n_537),
.Y(n_821)
);

INVx3_ASAP7_75t_L g822 ( 
.A(n_602),
.Y(n_822)
);

INVx2_ASAP7_75t_L g823 ( 
.A(n_599),
.Y(n_823)
);

NAND2xp5_ASAP7_75t_SL g824 ( 
.A(n_650),
.B(n_411),
.Y(n_824)
);

OR2x6_ASAP7_75t_L g825 ( 
.A(n_667),
.B(n_302),
.Y(n_825)
);

AOI22xp33_ASAP7_75t_L g826 ( 
.A1(n_599),
.A2(n_324),
.B1(n_333),
.B2(n_313),
.Y(n_826)
);

INVx2_ASAP7_75t_L g827 ( 
.A(n_726),
.Y(n_827)
);

AND2x4_ASAP7_75t_SL g828 ( 
.A(n_785),
.B(n_467),
.Y(n_828)
);

NAND2xp5_ASAP7_75t_SL g829 ( 
.A(n_732),
.B(n_507),
.Y(n_829)
);

BUFx6f_ASAP7_75t_SL g830 ( 
.A(n_698),
.Y(n_830)
);

BUFx3_ASAP7_75t_L g831 ( 
.A(n_817),
.Y(n_831)
);

AOI22xp33_ASAP7_75t_L g832 ( 
.A1(n_731),
.A2(n_371),
.B1(n_375),
.B2(n_370),
.Y(n_832)
);

INVx2_ASAP7_75t_L g833 ( 
.A(n_733),
.Y(n_833)
);

AOI22xp33_ASAP7_75t_L g834 ( 
.A1(n_746),
.A2(n_387),
.B1(n_390),
.B2(n_378),
.Y(n_834)
);

BUFx8_ASAP7_75t_L g835 ( 
.A(n_673),
.Y(n_835)
);

INVx1_ASAP7_75t_L g836 ( 
.A(n_815),
.Y(n_836)
);

HB1xp67_ASAP7_75t_L g837 ( 
.A(n_700),
.Y(n_837)
);

NAND2xp5_ASAP7_75t_SL g838 ( 
.A(n_732),
.B(n_623),
.Y(n_838)
);

INVx1_ASAP7_75t_L g839 ( 
.A(n_817),
.Y(n_839)
);

INVx1_ASAP7_75t_L g840 ( 
.A(n_796),
.Y(n_840)
);

INVx2_ASAP7_75t_L g841 ( 
.A(n_755),
.Y(n_841)
);

NAND2xp5_ASAP7_75t_L g842 ( 
.A(n_681),
.B(n_623),
.Y(n_842)
);

INVx2_ASAP7_75t_L g843 ( 
.A(n_767),
.Y(n_843)
);

NOR2xp67_ASAP7_75t_L g844 ( 
.A(n_674),
.B(n_667),
.Y(n_844)
);

OAI22xp5_ASAP7_75t_L g845 ( 
.A1(n_740),
.A2(n_472),
.B1(n_482),
.B2(n_471),
.Y(n_845)
);

NAND2xp5_ASAP7_75t_L g846 ( 
.A(n_701),
.B(n_623),
.Y(n_846)
);

NAND2xp5_ASAP7_75t_SL g847 ( 
.A(n_769),
.B(n_623),
.Y(n_847)
);

OR2x6_ASAP7_75t_L g848 ( 
.A(n_688),
.B(n_391),
.Y(n_848)
);

INVx2_ASAP7_75t_L g849 ( 
.A(n_669),
.Y(n_849)
);

AOI221xp5_ASAP7_75t_L g850 ( 
.A1(n_680),
.A2(n_429),
.B1(n_239),
.B2(n_244),
.C(n_238),
.Y(n_850)
);

NOR2xp33_ASAP7_75t_SL g851 ( 
.A(n_683),
.B(n_496),
.Y(n_851)
);

NAND2xp5_ASAP7_75t_SL g852 ( 
.A(n_769),
.B(n_624),
.Y(n_852)
);

AOI221xp5_ASAP7_75t_L g853 ( 
.A1(n_708),
.A2(n_258),
.B1(n_420),
.B2(n_434),
.C(n_335),
.Y(n_853)
);

INVx2_ASAP7_75t_SL g854 ( 
.A(n_684),
.Y(n_854)
);

NAND2xp5_ASAP7_75t_SL g855 ( 
.A(n_769),
.B(n_624),
.Y(n_855)
);

NAND2xp5_ASAP7_75t_SL g856 ( 
.A(n_769),
.B(n_624),
.Y(n_856)
);

NOR2x1p5_ASAP7_75t_L g857 ( 
.A(n_696),
.B(n_237),
.Y(n_857)
);

NAND2xp5_ASAP7_75t_L g858 ( 
.A(n_752),
.B(n_624),
.Y(n_858)
);

INVx1_ASAP7_75t_L g859 ( 
.A(n_797),
.Y(n_859)
);

OR2x2_ASAP7_75t_L g860 ( 
.A(n_696),
.B(n_237),
.Y(n_860)
);

NOR2xp33_ASAP7_75t_L g861 ( 
.A(n_672),
.B(n_725),
.Y(n_861)
);

NAND2xp5_ASAP7_75t_SL g862 ( 
.A(n_769),
.B(n_624),
.Y(n_862)
);

NAND2xp5_ASAP7_75t_L g863 ( 
.A(n_754),
.B(n_624),
.Y(n_863)
);

NAND2xp5_ASAP7_75t_L g864 ( 
.A(n_780),
.B(n_624),
.Y(n_864)
);

OAI22xp33_ASAP7_75t_L g865 ( 
.A1(n_780),
.A2(n_502),
.B1(n_513),
.B2(n_497),
.Y(n_865)
);

INVx2_ASAP7_75t_SL g866 ( 
.A(n_684),
.Y(n_866)
);

NAND2xp5_ASAP7_75t_L g867 ( 
.A(n_762),
.B(n_624),
.Y(n_867)
);

AOI22xp5_ASAP7_75t_L g868 ( 
.A1(n_789),
.A2(n_520),
.B1(n_522),
.B2(n_519),
.Y(n_868)
);

NAND2xp5_ASAP7_75t_L g869 ( 
.A(n_762),
.B(n_599),
.Y(n_869)
);

NAND2xp5_ASAP7_75t_SL g870 ( 
.A(n_781),
.B(n_599),
.Y(n_870)
);

INVx2_ASAP7_75t_L g871 ( 
.A(n_669),
.Y(n_871)
);

INVxp67_ASAP7_75t_L g872 ( 
.A(n_821),
.Y(n_872)
);

NAND2xp5_ASAP7_75t_L g873 ( 
.A(n_714),
.B(n_606),
.Y(n_873)
);

INVx3_ASAP7_75t_L g874 ( 
.A(n_814),
.Y(n_874)
);

NAND2xp5_ASAP7_75t_L g875 ( 
.A(n_813),
.B(n_606),
.Y(n_875)
);

INVx2_ASAP7_75t_L g876 ( 
.A(n_675),
.Y(n_876)
);

INVx4_ASAP7_75t_L g877 ( 
.A(n_735),
.Y(n_877)
);

NOR2xp33_ASAP7_75t_L g878 ( 
.A(n_672),
.B(n_255),
.Y(n_878)
);

NAND2xp5_ASAP7_75t_L g879 ( 
.A(n_686),
.B(n_606),
.Y(n_879)
);

NOR2xp67_ASAP7_75t_SL g880 ( 
.A(n_781),
.B(n_735),
.Y(n_880)
);

OAI221xp5_ASAP7_75t_L g881 ( 
.A1(n_826),
.A2(n_449),
.B1(n_398),
.B2(n_447),
.C(n_436),
.Y(n_881)
);

INVx3_ASAP7_75t_L g882 ( 
.A(n_814),
.Y(n_882)
);

NAND2xp5_ASAP7_75t_L g883 ( 
.A(n_686),
.B(n_606),
.Y(n_883)
);

OR2x2_ASAP7_75t_L g884 ( 
.A(n_765),
.B(n_238),
.Y(n_884)
);

NAND2xp5_ASAP7_75t_L g885 ( 
.A(n_775),
.B(n_617),
.Y(n_885)
);

INVx1_ASAP7_75t_L g886 ( 
.A(n_801),
.Y(n_886)
);

NAND2xp5_ASAP7_75t_SL g887 ( 
.A(n_781),
.B(n_617),
.Y(n_887)
);

INVx2_ASAP7_75t_L g888 ( 
.A(n_675),
.Y(n_888)
);

NOR2xp33_ASAP7_75t_L g889 ( 
.A(n_725),
.B(n_255),
.Y(n_889)
);

NAND2xp5_ASAP7_75t_L g890 ( 
.A(n_791),
.B(n_617),
.Y(n_890)
);

AOI21xp5_ASAP7_75t_L g891 ( 
.A1(n_694),
.A2(n_615),
.B(n_617),
.Y(n_891)
);

AOI22xp33_ASAP7_75t_L g892 ( 
.A1(n_804),
.A2(n_433),
.B1(n_415),
.B2(n_264),
.Y(n_892)
);

INVx1_ASAP7_75t_L g893 ( 
.A(n_805),
.Y(n_893)
);

BUFx6f_ASAP7_75t_SL g894 ( 
.A(n_698),
.Y(n_894)
);

NOR2xp67_ASAP7_75t_L g895 ( 
.A(n_759),
.B(n_710),
.Y(n_895)
);

NAND2xp5_ASAP7_75t_SL g896 ( 
.A(n_781),
.B(n_625),
.Y(n_896)
);

NAND2xp5_ASAP7_75t_SL g897 ( 
.A(n_781),
.B(n_625),
.Y(n_897)
);

NOR3xp33_ASAP7_75t_L g898 ( 
.A(n_792),
.B(n_312),
.C(n_304),
.Y(n_898)
);

NAND2xp5_ASAP7_75t_L g899 ( 
.A(n_791),
.B(n_625),
.Y(n_899)
);

NAND2xp5_ASAP7_75t_L g900 ( 
.A(n_671),
.B(n_625),
.Y(n_900)
);

NAND2xp5_ASAP7_75t_L g901 ( 
.A(n_678),
.B(n_627),
.Y(n_901)
);

INVx3_ASAP7_75t_L g902 ( 
.A(n_814),
.Y(n_902)
);

NAND2xp5_ASAP7_75t_L g903 ( 
.A(n_690),
.B(n_627),
.Y(n_903)
);

NOR2xp33_ASAP7_75t_L g904 ( 
.A(n_734),
.B(n_747),
.Y(n_904)
);

BUFx6f_ASAP7_75t_L g905 ( 
.A(n_735),
.Y(n_905)
);

AOI22xp5_ASAP7_75t_L g906 ( 
.A1(n_789),
.A2(n_261),
.B1(n_263),
.B2(n_260),
.Y(n_906)
);

INVx1_ASAP7_75t_L g907 ( 
.A(n_772),
.Y(n_907)
);

INVx2_ASAP7_75t_L g908 ( 
.A(n_679),
.Y(n_908)
);

NAND2xp5_ASAP7_75t_L g909 ( 
.A(n_774),
.B(n_627),
.Y(n_909)
);

NAND2xp5_ASAP7_75t_SL g910 ( 
.A(n_783),
.B(n_627),
.Y(n_910)
);

O2A1O1Ixp33_ASAP7_75t_L g911 ( 
.A1(n_811),
.A2(n_634),
.B(n_647),
.C(n_637),
.Y(n_911)
);

INVx2_ASAP7_75t_L g912 ( 
.A(n_679),
.Y(n_912)
);

AOI22xp5_ASAP7_75t_L g913 ( 
.A1(n_783),
.A2(n_261),
.B1(n_263),
.B2(n_260),
.Y(n_913)
);

AOI22xp5_ASAP7_75t_L g914 ( 
.A1(n_722),
.A2(n_268),
.B1(n_341),
.B2(n_267),
.Y(n_914)
);

INVxp67_ASAP7_75t_L g915 ( 
.A(n_765),
.Y(n_915)
);

HB1xp67_ASAP7_75t_L g916 ( 
.A(n_750),
.Y(n_916)
);

INVx2_ASAP7_75t_L g917 ( 
.A(n_702),
.Y(n_917)
);

NAND2xp5_ASAP7_75t_L g918 ( 
.A(n_778),
.B(n_634),
.Y(n_918)
);

INVx1_ASAP7_75t_L g919 ( 
.A(n_779),
.Y(n_919)
);

INVx2_ASAP7_75t_L g920 ( 
.A(n_702),
.Y(n_920)
);

NAND2xp5_ASAP7_75t_L g921 ( 
.A(n_790),
.B(n_634),
.Y(n_921)
);

NAND2xp5_ASAP7_75t_L g922 ( 
.A(n_794),
.B(n_634),
.Y(n_922)
);

INVx2_ASAP7_75t_SL g923 ( 
.A(n_728),
.Y(n_923)
);

NAND2xp5_ASAP7_75t_L g924 ( 
.A(n_670),
.B(n_637),
.Y(n_924)
);

O2A1O1Ixp5_ASAP7_75t_L g925 ( 
.A1(n_808),
.A2(n_604),
.B(n_647),
.C(n_637),
.Y(n_925)
);

AOI22xp33_ASAP7_75t_L g926 ( 
.A1(n_804),
.A2(n_289),
.B1(n_303),
.B2(n_248),
.Y(n_926)
);

INVxp33_ASAP7_75t_L g927 ( 
.A(n_704),
.Y(n_927)
);

INVx2_ASAP7_75t_L g928 ( 
.A(n_709),
.Y(n_928)
);

NAND2xp5_ASAP7_75t_SL g929 ( 
.A(n_806),
.B(n_637),
.Y(n_929)
);

NOR2xp33_ASAP7_75t_L g930 ( 
.A(n_753),
.B(n_267),
.Y(n_930)
);

NAND2xp5_ASAP7_75t_L g931 ( 
.A(n_676),
.B(n_647),
.Y(n_931)
);

NAND2x1_ASAP7_75t_L g932 ( 
.A(n_695),
.B(n_604),
.Y(n_932)
);

NAND2xp5_ASAP7_75t_L g933 ( 
.A(n_677),
.B(n_647),
.Y(n_933)
);

NAND2xp5_ASAP7_75t_SL g934 ( 
.A(n_806),
.B(n_602),
.Y(n_934)
);

NAND2xp5_ASAP7_75t_L g935 ( 
.A(n_682),
.B(n_602),
.Y(n_935)
);

NAND2xp33_ASAP7_75t_L g936 ( 
.A(n_737),
.B(n_254),
.Y(n_936)
);

NAND2xp5_ASAP7_75t_L g937 ( 
.A(n_685),
.B(n_689),
.Y(n_937)
);

NAND2xp33_ASAP7_75t_L g938 ( 
.A(n_744),
.B(n_254),
.Y(n_938)
);

NAND2xp5_ASAP7_75t_L g939 ( 
.A(n_691),
.B(n_602),
.Y(n_939)
);

OAI22xp33_ASAP7_75t_L g940 ( 
.A1(n_785),
.A2(n_257),
.B1(n_262),
.B2(n_251),
.Y(n_940)
);

INVx1_ASAP7_75t_L g941 ( 
.A(n_787),
.Y(n_941)
);

INVx1_ASAP7_75t_L g942 ( 
.A(n_787),
.Y(n_942)
);

INVx2_ASAP7_75t_SL g943 ( 
.A(n_728),
.Y(n_943)
);

NAND2xp5_ASAP7_75t_L g944 ( 
.A(n_692),
.B(n_602),
.Y(n_944)
);

INVx2_ASAP7_75t_L g945 ( 
.A(n_709),
.Y(n_945)
);

AND2x2_ASAP7_75t_L g946 ( 
.A(n_749),
.B(n_559),
.Y(n_946)
);

INVx2_ASAP7_75t_L g947 ( 
.A(n_712),
.Y(n_947)
);

AND2x2_ASAP7_75t_L g948 ( 
.A(n_699),
.B(n_559),
.Y(n_948)
);

INVx2_ASAP7_75t_SL g949 ( 
.A(n_728),
.Y(n_949)
);

OR2x2_ASAP7_75t_SL g950 ( 
.A(n_798),
.B(n_353),
.Y(n_950)
);

NAND2xp5_ASAP7_75t_L g951 ( 
.A(n_705),
.B(n_607),
.Y(n_951)
);

NAND2xp5_ASAP7_75t_SL g952 ( 
.A(n_788),
.B(n_607),
.Y(n_952)
);

INVxp33_ASAP7_75t_L g953 ( 
.A(n_795),
.Y(n_953)
);

NAND2xp5_ASAP7_75t_L g954 ( 
.A(n_713),
.B(n_607),
.Y(n_954)
);

NOR3xp33_ASAP7_75t_L g955 ( 
.A(n_799),
.B(n_320),
.C(n_314),
.Y(n_955)
);

AO22x2_ASAP7_75t_L g956 ( 
.A1(n_808),
.A2(n_824),
.B1(n_788),
.B2(n_751),
.Y(n_956)
);

BUFx6f_ASAP7_75t_L g957 ( 
.A(n_703),
.Y(n_957)
);

INVx2_ASAP7_75t_SL g958 ( 
.A(n_724),
.Y(n_958)
);

AND2x2_ASAP7_75t_L g959 ( 
.A(n_683),
.B(n_566),
.Y(n_959)
);

AOI22xp5_ASAP7_75t_L g960 ( 
.A1(n_722),
.A2(n_341),
.B1(n_414),
.B2(n_268),
.Y(n_960)
);

NAND3xp33_ASAP7_75t_L g961 ( 
.A(n_751),
.B(n_326),
.C(n_323),
.Y(n_961)
);

NAND2xp5_ASAP7_75t_L g962 ( 
.A(n_716),
.B(n_607),
.Y(n_962)
);

INVx1_ASAP7_75t_L g963 ( 
.A(n_812),
.Y(n_963)
);

AOI22xp33_ASAP7_75t_L g964 ( 
.A1(n_804),
.A2(n_361),
.B1(n_380),
.B2(n_377),
.Y(n_964)
);

INVx2_ASAP7_75t_SL g965 ( 
.A(n_750),
.Y(n_965)
);

NOR2xp33_ASAP7_75t_L g966 ( 
.A(n_698),
.B(n_414),
.Y(n_966)
);

AOI22xp5_ASAP7_75t_L g967 ( 
.A1(n_785),
.A2(n_421),
.B1(n_423),
.B2(n_417),
.Y(n_967)
);

INVx1_ASAP7_75t_L g968 ( 
.A(n_812),
.Y(n_968)
);

INVx2_ASAP7_75t_L g969 ( 
.A(n_712),
.Y(n_969)
);

INVx1_ASAP7_75t_L g970 ( 
.A(n_820),
.Y(n_970)
);

INVx1_ASAP7_75t_L g971 ( 
.A(n_820),
.Y(n_971)
);

INVx2_ASAP7_75t_L g972 ( 
.A(n_715),
.Y(n_972)
);

NAND2xp5_ASAP7_75t_L g973 ( 
.A(n_719),
.B(n_607),
.Y(n_973)
);

NOR2xp33_ASAP7_75t_L g974 ( 
.A(n_698),
.B(n_417),
.Y(n_974)
);

NOR3xp33_ASAP7_75t_L g975 ( 
.A(n_816),
.B(n_332),
.C(n_330),
.Y(n_975)
);

NAND2xp5_ASAP7_75t_SL g976 ( 
.A(n_788),
.B(n_607),
.Y(n_976)
);

NAND2xp5_ASAP7_75t_L g977 ( 
.A(n_721),
.B(n_760),
.Y(n_977)
);

INVx1_ASAP7_75t_L g978 ( 
.A(n_825),
.Y(n_978)
);

INVx1_ASAP7_75t_L g979 ( 
.A(n_825),
.Y(n_979)
);

NAND2xp5_ASAP7_75t_L g980 ( 
.A(n_766),
.B(n_607),
.Y(n_980)
);

INVx1_ASAP7_75t_L g981 ( 
.A(n_825),
.Y(n_981)
);

NAND2xp5_ASAP7_75t_L g982 ( 
.A(n_822),
.B(n_607),
.Y(n_982)
);

BUFx6f_ASAP7_75t_L g983 ( 
.A(n_703),
.Y(n_983)
);

O2A1O1Ixp33_ASAP7_75t_L g984 ( 
.A1(n_742),
.A2(n_615),
.B(n_580),
.C(n_581),
.Y(n_984)
);

BUFx6f_ASAP7_75t_L g985 ( 
.A(n_703),
.Y(n_985)
);

CKINVDCx5p33_ASAP7_75t_R g986 ( 
.A(n_693),
.Y(n_986)
);

NOR2xp33_ASAP7_75t_L g987 ( 
.A(n_785),
.B(n_421),
.Y(n_987)
);

BUFx5_ASAP7_75t_L g988 ( 
.A(n_706),
.Y(n_988)
);

INVx1_ASAP7_75t_L g989 ( 
.A(n_825),
.Y(n_989)
);

NAND2xp5_ASAP7_75t_SL g990 ( 
.A(n_788),
.B(n_254),
.Y(n_990)
);

BUFx3_ASAP7_75t_L g991 ( 
.A(n_804),
.Y(n_991)
);

INVx1_ASAP7_75t_L g992 ( 
.A(n_764),
.Y(n_992)
);

NAND2xp5_ASAP7_75t_SL g993 ( 
.A(n_822),
.B(n_800),
.Y(n_993)
);

INVx2_ASAP7_75t_L g994 ( 
.A(n_715),
.Y(n_994)
);

NAND2xp5_ASAP7_75t_L g995 ( 
.A(n_822),
.B(n_579),
.Y(n_995)
);

NAND2xp5_ASAP7_75t_L g996 ( 
.A(n_695),
.B(n_579),
.Y(n_996)
);

OA21x2_ASAP7_75t_L g997 ( 
.A1(n_819),
.A2(n_611),
.B(n_605),
.Y(n_997)
);

INVx3_ASAP7_75t_L g998 ( 
.A(n_905),
.Y(n_998)
);

INVx3_ASAP7_75t_L g999 ( 
.A(n_905),
.Y(n_999)
);

NAND2xp5_ASAP7_75t_L g1000 ( 
.A(n_904),
.B(n_800),
.Y(n_1000)
);

OAI22xp5_ASAP7_75t_L g1001 ( 
.A1(n_904),
.A2(n_763),
.B1(n_768),
.B2(n_764),
.Y(n_1001)
);

AOI21xp5_ASAP7_75t_L g1002 ( 
.A1(n_869),
.A2(n_867),
.B(n_873),
.Y(n_1002)
);

NOR2x1_ASAP7_75t_R g1003 ( 
.A(n_986),
.B(n_687),
.Y(n_1003)
);

INVx1_ASAP7_75t_L g1004 ( 
.A(n_840),
.Y(n_1004)
);

NAND2xp5_ASAP7_75t_L g1005 ( 
.A(n_844),
.B(n_807),
.Y(n_1005)
);

NAND2xp5_ASAP7_75t_L g1006 ( 
.A(n_885),
.B(n_807),
.Y(n_1006)
);

INVx2_ASAP7_75t_SL g1007 ( 
.A(n_837),
.Y(n_1007)
);

AOI21xp5_ASAP7_75t_L g1008 ( 
.A1(n_910),
.A2(n_782),
.B(n_742),
.Y(n_1008)
);

AND2x2_ASAP7_75t_L g1009 ( 
.A(n_959),
.B(n_687),
.Y(n_1009)
);

OAI21xp5_ASAP7_75t_L g1010 ( 
.A1(n_910),
.A2(n_782),
.B(n_809),
.Y(n_1010)
);

NAND2xp5_ASAP7_75t_L g1011 ( 
.A(n_861),
.B(n_809),
.Y(n_1011)
);

NAND2xp5_ASAP7_75t_L g1012 ( 
.A(n_861),
.B(n_810),
.Y(n_1012)
);

AOI22xp5_ASAP7_75t_L g1013 ( 
.A1(n_895),
.A2(n_763),
.B1(n_706),
.B2(n_707),
.Y(n_1013)
);

INVx3_ASAP7_75t_L g1014 ( 
.A(n_905),
.Y(n_1014)
);

HB1xp67_ASAP7_75t_L g1015 ( 
.A(n_916),
.Y(n_1015)
);

NAND2xp5_ASAP7_75t_L g1016 ( 
.A(n_875),
.B(n_810),
.Y(n_1016)
);

NAND2xp5_ASAP7_75t_SL g1017 ( 
.A(n_892),
.B(n_718),
.Y(n_1017)
);

NAND2xp5_ASAP7_75t_L g1018 ( 
.A(n_900),
.B(n_818),
.Y(n_1018)
);

AOI22xp33_ASAP7_75t_L g1019 ( 
.A1(n_892),
.A2(n_771),
.B1(n_776),
.B2(n_768),
.Y(n_1019)
);

A2O1A1Ixp33_ASAP7_75t_L g1020 ( 
.A1(n_930),
.A2(n_269),
.B(n_271),
.C(n_265),
.Y(n_1020)
);

NAND2xp5_ASAP7_75t_L g1021 ( 
.A(n_901),
.B(n_818),
.Y(n_1021)
);

A2O1A1Ixp33_ASAP7_75t_L g1022 ( 
.A1(n_930),
.A2(n_274),
.B(n_275),
.C(n_272),
.Y(n_1022)
);

NAND2xp5_ASAP7_75t_L g1023 ( 
.A(n_903),
.B(n_823),
.Y(n_1023)
);

AOI21xp5_ASAP7_75t_L g1024 ( 
.A1(n_858),
.A2(n_776),
.B(n_771),
.Y(n_1024)
);

CKINVDCx20_ASAP7_75t_R g1025 ( 
.A(n_868),
.Y(n_1025)
);

AOI21xp5_ASAP7_75t_L g1026 ( 
.A1(n_863),
.A2(n_793),
.B(n_730),
.Y(n_1026)
);

AOI21xp5_ASAP7_75t_L g1027 ( 
.A1(n_842),
.A2(n_793),
.B(n_730),
.Y(n_1027)
);

INVx1_ASAP7_75t_L g1028 ( 
.A(n_859),
.Y(n_1028)
);

NAND2xp5_ASAP7_75t_L g1029 ( 
.A(n_890),
.B(n_823),
.Y(n_1029)
);

INVx3_ASAP7_75t_L g1030 ( 
.A(n_905),
.Y(n_1030)
);

INVx1_ASAP7_75t_L g1031 ( 
.A(n_886),
.Y(n_1031)
);

AOI21xp5_ASAP7_75t_L g1032 ( 
.A1(n_846),
.A2(n_730),
.B(n_697),
.Y(n_1032)
);

OAI21xp5_ASAP7_75t_L g1033 ( 
.A1(n_925),
.A2(n_929),
.B(n_911),
.Y(n_1033)
);

INVx2_ASAP7_75t_L g1034 ( 
.A(n_849),
.Y(n_1034)
);

NAND2xp5_ASAP7_75t_L g1035 ( 
.A(n_899),
.B(n_695),
.Y(n_1035)
);

NAND2xp5_ASAP7_75t_L g1036 ( 
.A(n_963),
.B(n_711),
.Y(n_1036)
);

AOI21xp5_ASAP7_75t_L g1037 ( 
.A1(n_980),
.A2(n_786),
.B(n_697),
.Y(n_1037)
);

AOI21xp5_ASAP7_75t_L g1038 ( 
.A1(n_864),
.A2(n_786),
.B(n_697),
.Y(n_1038)
);

OAI21xp5_ASAP7_75t_L g1039 ( 
.A1(n_929),
.A2(n_717),
.B(n_786),
.Y(n_1039)
);

AND2x2_ASAP7_75t_L g1040 ( 
.A(n_946),
.B(n_718),
.Y(n_1040)
);

AOI22xp5_ASAP7_75t_L g1041 ( 
.A1(n_975),
.A2(n_707),
.B1(n_706),
.B2(n_803),
.Y(n_1041)
);

AO21x1_ASAP7_75t_L g1042 ( 
.A1(n_936),
.A2(n_282),
.B(n_280),
.Y(n_1042)
);

AND2x2_ASAP7_75t_L g1043 ( 
.A(n_872),
.B(n_757),
.Y(n_1043)
);

NAND2xp5_ASAP7_75t_L g1044 ( 
.A(n_968),
.B(n_970),
.Y(n_1044)
);

INVx1_ASAP7_75t_L g1045 ( 
.A(n_893),
.Y(n_1045)
);

O2A1O1Ixp33_ASAP7_75t_L g1046 ( 
.A1(n_971),
.A2(n_581),
.B(n_585),
.C(n_580),
.Y(n_1046)
);

AOI21xp5_ASAP7_75t_L g1047 ( 
.A1(n_838),
.A2(n_803),
.B(n_717),
.Y(n_1047)
);

INVx4_ASAP7_75t_L g1048 ( 
.A(n_831),
.Y(n_1048)
);

AOI21xp5_ASAP7_75t_L g1049 ( 
.A1(n_838),
.A2(n_803),
.B(n_729),
.Y(n_1049)
);

INVx2_ASAP7_75t_L g1050 ( 
.A(n_871),
.Y(n_1050)
);

NAND2xp5_ASAP7_75t_L g1051 ( 
.A(n_878),
.B(n_711),
.Y(n_1051)
);

AOI21xp5_ASAP7_75t_L g1052 ( 
.A1(n_934),
.A2(n_729),
.B(n_711),
.Y(n_1052)
);

AOI21xp5_ASAP7_75t_L g1053 ( 
.A1(n_934),
.A2(n_739),
.B(n_729),
.Y(n_1053)
);

HB1xp67_ASAP7_75t_L g1054 ( 
.A(n_965),
.Y(n_1054)
);

AOI21xp5_ASAP7_75t_L g1055 ( 
.A1(n_938),
.A2(n_756),
.B(n_739),
.Y(n_1055)
);

BUFx6f_ASAP7_75t_L g1056 ( 
.A(n_831),
.Y(n_1056)
);

INVx3_ASAP7_75t_L g1057 ( 
.A(n_874),
.Y(n_1057)
);

AOI22xp5_ASAP7_75t_L g1058 ( 
.A1(n_898),
.A2(n_707),
.B1(n_706),
.B2(n_296),
.Y(n_1058)
);

INVx2_ASAP7_75t_SL g1059 ( 
.A(n_857),
.Y(n_1059)
);

INVx1_ASAP7_75t_L g1060 ( 
.A(n_907),
.Y(n_1060)
);

NAND2xp5_ASAP7_75t_L g1061 ( 
.A(n_878),
.B(n_739),
.Y(n_1061)
);

NAND2xp5_ASAP7_75t_L g1062 ( 
.A(n_889),
.B(n_756),
.Y(n_1062)
);

INVx4_ASAP7_75t_L g1063 ( 
.A(n_874),
.Y(n_1063)
);

OR2x6_ASAP7_75t_L g1064 ( 
.A(n_958),
.B(n_848),
.Y(n_1064)
);

OAI21xp33_ASAP7_75t_L g1065 ( 
.A1(n_853),
.A2(n_850),
.B(n_926),
.Y(n_1065)
);

OAI21xp5_ASAP7_75t_L g1066 ( 
.A1(n_827),
.A2(n_758),
.B(n_756),
.Y(n_1066)
);

NAND2xp5_ASAP7_75t_L g1067 ( 
.A(n_889),
.B(n_758),
.Y(n_1067)
);

OR2x6_ASAP7_75t_L g1068 ( 
.A(n_848),
.B(n_297),
.Y(n_1068)
);

NOR2xp33_ASAP7_75t_L g1069 ( 
.A(n_953),
.B(n_409),
.Y(n_1069)
);

AOI21xp5_ASAP7_75t_L g1070 ( 
.A1(n_879),
.A2(n_758),
.B(n_723),
.Y(n_1070)
);

NAND2xp5_ASAP7_75t_L g1071 ( 
.A(n_941),
.B(n_703),
.Y(n_1071)
);

NAND2xp5_ASAP7_75t_L g1072 ( 
.A(n_942),
.B(n_761),
.Y(n_1072)
);

BUFx6f_ASAP7_75t_L g1073 ( 
.A(n_991),
.Y(n_1073)
);

NAND2xp5_ASAP7_75t_SL g1074 ( 
.A(n_854),
.B(n_423),
.Y(n_1074)
);

BUFx6f_ASAP7_75t_L g1075 ( 
.A(n_991),
.Y(n_1075)
);

NAND2xp5_ASAP7_75t_SL g1076 ( 
.A(n_866),
.B(n_425),
.Y(n_1076)
);

NAND2xp5_ASAP7_75t_L g1077 ( 
.A(n_827),
.B(n_761),
.Y(n_1077)
);

NAND2xp5_ASAP7_75t_L g1078 ( 
.A(n_833),
.B(n_761),
.Y(n_1078)
);

NAND2xp5_ASAP7_75t_L g1079 ( 
.A(n_833),
.B(n_761),
.Y(n_1079)
);

NAND2xp5_ASAP7_75t_L g1080 ( 
.A(n_841),
.B(n_720),
.Y(n_1080)
);

INVx2_ASAP7_75t_L g1081 ( 
.A(n_888),
.Y(n_1081)
);

NOR2xp33_ASAP7_75t_L g1082 ( 
.A(n_927),
.B(n_410),
.Y(n_1082)
);

NAND2xp5_ASAP7_75t_L g1083 ( 
.A(n_841),
.B(n_727),
.Y(n_1083)
);

AOI21xp5_ASAP7_75t_L g1084 ( 
.A1(n_883),
.A2(n_736),
.B(n_727),
.Y(n_1084)
);

OAI21xp5_ASAP7_75t_L g1085 ( 
.A1(n_843),
.A2(n_738),
.B(n_736),
.Y(n_1085)
);

NOR2xp33_ASAP7_75t_L g1086 ( 
.A(n_915),
.B(n_444),
.Y(n_1086)
);

NAND2xp5_ASAP7_75t_L g1087 ( 
.A(n_843),
.B(n_738),
.Y(n_1087)
);

NAND2xp5_ASAP7_75t_L g1088 ( 
.A(n_919),
.B(n_741),
.Y(n_1088)
);

AOI21xp5_ASAP7_75t_L g1089 ( 
.A1(n_977),
.A2(n_743),
.B(n_741),
.Y(n_1089)
);

INVx2_ASAP7_75t_L g1090 ( 
.A(n_888),
.Y(n_1090)
);

BUFx6f_ASAP7_75t_L g1091 ( 
.A(n_957),
.Y(n_1091)
);

NOR2xp33_ASAP7_75t_L g1092 ( 
.A(n_829),
.B(n_865),
.Y(n_1092)
);

NAND2xp5_ASAP7_75t_L g1093 ( 
.A(n_832),
.B(n_743),
.Y(n_1093)
);

INVx2_ASAP7_75t_SL g1094 ( 
.A(n_848),
.Y(n_1094)
);

INVx1_ASAP7_75t_L g1095 ( 
.A(n_839),
.Y(n_1095)
);

AND2x2_ASAP7_75t_L g1096 ( 
.A(n_948),
.B(n_566),
.Y(n_1096)
);

NAND2xp5_ASAP7_75t_L g1097 ( 
.A(n_832),
.B(n_834),
.Y(n_1097)
);

HB1xp67_ASAP7_75t_L g1098 ( 
.A(n_836),
.Y(n_1098)
);

NAND2xp5_ASAP7_75t_L g1099 ( 
.A(n_834),
.B(n_745),
.Y(n_1099)
);

INVx1_ASAP7_75t_L g1100 ( 
.A(n_937),
.Y(n_1100)
);

AND2x2_ASAP7_75t_L g1101 ( 
.A(n_860),
.B(n_568),
.Y(n_1101)
);

A2O1A1Ixp33_ASAP7_75t_L g1102 ( 
.A1(n_987),
.A2(n_424),
.B(n_329),
.C(n_322),
.Y(n_1102)
);

AND2x4_ASAP7_75t_L g1103 ( 
.A(n_923),
.B(n_568),
.Y(n_1103)
);

AOI21xp5_ASAP7_75t_L g1104 ( 
.A1(n_909),
.A2(n_921),
.B(n_918),
.Y(n_1104)
);

INVxp67_ASAP7_75t_L g1105 ( 
.A(n_829),
.Y(n_1105)
);

AOI22xp5_ASAP7_75t_L g1106 ( 
.A1(n_943),
.A2(n_949),
.B1(n_961),
.B2(n_978),
.Y(n_1106)
);

OAI21xp5_ASAP7_75t_L g1107 ( 
.A1(n_891),
.A2(n_770),
.B(n_748),
.Y(n_1107)
);

NAND2xp5_ASAP7_75t_L g1108 ( 
.A(n_992),
.B(n_770),
.Y(n_1108)
);

INVx3_ASAP7_75t_L g1109 ( 
.A(n_882),
.Y(n_1109)
);

INVx5_ASAP7_75t_L g1110 ( 
.A(n_957),
.Y(n_1110)
);

AND2x2_ASAP7_75t_L g1111 ( 
.A(n_884),
.B(n_239),
.Y(n_1111)
);

AND2x4_ASAP7_75t_L g1112 ( 
.A(n_979),
.B(n_310),
.Y(n_1112)
);

BUFx4f_ASAP7_75t_L g1113 ( 
.A(n_828),
.Y(n_1113)
);

HB1xp67_ASAP7_75t_L g1114 ( 
.A(n_981),
.Y(n_1114)
);

OAI21xp5_ASAP7_75t_L g1115 ( 
.A1(n_922),
.A2(n_777),
.B(n_773),
.Y(n_1115)
);

AOI21xp5_ASAP7_75t_L g1116 ( 
.A1(n_935),
.A2(n_944),
.B(n_939),
.Y(n_1116)
);

NAND3xp33_ASAP7_75t_L g1117 ( 
.A(n_926),
.B(n_340),
.C(n_338),
.Y(n_1117)
);

NOR2xp33_ASAP7_75t_L g1118 ( 
.A(n_845),
.B(n_851),
.Y(n_1118)
);

INVx1_ASAP7_75t_L g1119 ( 
.A(n_908),
.Y(n_1119)
);

INVx1_ASAP7_75t_L g1120 ( 
.A(n_912),
.Y(n_1120)
);

OAI21xp5_ASAP7_75t_L g1121 ( 
.A1(n_993),
.A2(n_777),
.B(n_773),
.Y(n_1121)
);

OAI21xp5_ASAP7_75t_L g1122 ( 
.A1(n_993),
.A2(n_707),
.B(n_706),
.Y(n_1122)
);

AOI21xp5_ASAP7_75t_L g1123 ( 
.A1(n_924),
.A2(n_582),
.B(n_604),
.Y(n_1123)
);

INVx2_ASAP7_75t_SL g1124 ( 
.A(n_835),
.Y(n_1124)
);

AOI21xp5_ASAP7_75t_L g1125 ( 
.A1(n_931),
.A2(n_582),
.B(n_577),
.Y(n_1125)
);

NOR2xp67_ASAP7_75t_L g1126 ( 
.A(n_914),
.B(n_425),
.Y(n_1126)
);

AOI22xp5_ASAP7_75t_L g1127 ( 
.A1(n_989),
.A2(n_706),
.B1(n_707),
.B2(n_315),
.Y(n_1127)
);

INVx2_ASAP7_75t_L g1128 ( 
.A(n_912),
.Y(n_1128)
);

NAND2xp5_ASAP7_75t_SL g1129 ( 
.A(n_987),
.B(n_435),
.Y(n_1129)
);

OAI22xp5_ASAP7_75t_L g1130 ( 
.A1(n_956),
.A2(n_352),
.B1(n_381),
.B2(n_362),
.Y(n_1130)
);

AOI21xp5_ASAP7_75t_L g1131 ( 
.A1(n_933),
.A2(n_582),
.B(n_577),
.Y(n_1131)
);

OR2x6_ASAP7_75t_SL g1132 ( 
.A(n_964),
.B(n_244),
.Y(n_1132)
);

AOI21xp5_ASAP7_75t_L g1133 ( 
.A1(n_982),
.A2(n_582),
.B(n_577),
.Y(n_1133)
);

NAND2xp5_ASAP7_75t_L g1134 ( 
.A(n_877),
.B(n_707),
.Y(n_1134)
);

OAI22xp5_ASAP7_75t_L g1135 ( 
.A1(n_956),
.A2(n_441),
.B1(n_359),
.B2(n_448),
.Y(n_1135)
);

INVx2_ASAP7_75t_L g1136 ( 
.A(n_917),
.Y(n_1136)
);

NAND2xp5_ASAP7_75t_L g1137 ( 
.A(n_877),
.B(n_318),
.Y(n_1137)
);

NAND2xp5_ASAP7_75t_SL g1138 ( 
.A(n_913),
.B(n_435),
.Y(n_1138)
);

INVx2_ASAP7_75t_L g1139 ( 
.A(n_917),
.Y(n_1139)
);

NAND2xp5_ASAP7_75t_L g1140 ( 
.A(n_882),
.B(n_902),
.Y(n_1140)
);

INVx1_ASAP7_75t_L g1141 ( 
.A(n_928),
.Y(n_1141)
);

AND2x2_ASAP7_75t_L g1142 ( 
.A(n_964),
.B(n_249),
.Y(n_1142)
);

AOI21xp5_ASAP7_75t_L g1143 ( 
.A1(n_870),
.A2(n_582),
.B(n_577),
.Y(n_1143)
);

AOI21xp5_ASAP7_75t_L g1144 ( 
.A1(n_870),
.A2(n_896),
.B(n_887),
.Y(n_1144)
);

NAND2x1p5_ASAP7_75t_L g1145 ( 
.A(n_880),
.B(n_386),
.Y(n_1145)
);

AOI21xp5_ASAP7_75t_L g1146 ( 
.A1(n_887),
.A2(n_897),
.B(n_896),
.Y(n_1146)
);

OAI22xp5_ASAP7_75t_L g1147 ( 
.A1(n_956),
.A2(n_419),
.B1(n_393),
.B2(n_416),
.Y(n_1147)
);

INVx2_ASAP7_75t_SL g1148 ( 
.A(n_835),
.Y(n_1148)
);

NOR3xp33_ASAP7_75t_L g1149 ( 
.A(n_966),
.B(n_438),
.C(n_437),
.Y(n_1149)
);

OAI22xp5_ASAP7_75t_L g1150 ( 
.A1(n_967),
.A2(n_408),
.B1(n_445),
.B2(n_450),
.Y(n_1150)
);

NOR3xp33_ASAP7_75t_L g1151 ( 
.A(n_966),
.B(n_438),
.C(n_437),
.Y(n_1151)
);

OA21x2_ASAP7_75t_L g1152 ( 
.A1(n_951),
.A2(n_611),
.B(n_605),
.Y(n_1152)
);

BUFx12f_ASAP7_75t_L g1153 ( 
.A(n_950),
.Y(n_1153)
);

NAND2xp5_ASAP7_75t_L g1154 ( 
.A(n_902),
.B(n_585),
.Y(n_1154)
);

INVx4_ASAP7_75t_L g1155 ( 
.A(n_957),
.Y(n_1155)
);

CKINVDCx8_ASAP7_75t_R g1156 ( 
.A(n_974),
.Y(n_1156)
);

INVx2_ASAP7_75t_L g1157 ( 
.A(n_928),
.Y(n_1157)
);

AOI21xp5_ASAP7_75t_L g1158 ( 
.A1(n_897),
.A2(n_582),
.B(n_577),
.Y(n_1158)
);

O2A1O1Ixp33_ASAP7_75t_L g1159 ( 
.A1(n_984),
.A2(n_628),
.B(n_587),
.C(n_663),
.Y(n_1159)
);

INVx2_ASAP7_75t_L g1160 ( 
.A(n_947),
.Y(n_1160)
);

NAND2xp5_ASAP7_75t_L g1161 ( 
.A(n_947),
.B(n_586),
.Y(n_1161)
);

AOI21xp5_ASAP7_75t_L g1162 ( 
.A1(n_954),
.A2(n_582),
.B(n_584),
.Y(n_1162)
);

NAND2xp5_ASAP7_75t_SL g1163 ( 
.A(n_974),
.B(n_439),
.Y(n_1163)
);

BUFx4f_ASAP7_75t_L g1164 ( 
.A(n_828),
.Y(n_1164)
);

HB1xp67_ASAP7_75t_L g1165 ( 
.A(n_830),
.Y(n_1165)
);

OAI21xp5_ASAP7_75t_L g1166 ( 
.A1(n_952),
.A2(n_611),
.B(n_605),
.Y(n_1166)
);

NAND2xp5_ASAP7_75t_L g1167 ( 
.A(n_969),
.B(n_586),
.Y(n_1167)
);

OAI22xp5_ASAP7_75t_L g1168 ( 
.A1(n_906),
.A2(n_446),
.B1(n_439),
.B2(n_450),
.Y(n_1168)
);

INVx2_ASAP7_75t_L g1169 ( 
.A(n_969),
.Y(n_1169)
);

NOR2x1_ASAP7_75t_L g1170 ( 
.A(n_940),
.B(n_587),
.Y(n_1170)
);

AOI21xp5_ASAP7_75t_L g1171 ( 
.A1(n_962),
.A2(n_582),
.B(n_584),
.Y(n_1171)
);

OAI22xp5_ASAP7_75t_L g1172 ( 
.A1(n_960),
.A2(n_446),
.B1(n_588),
.B2(n_663),
.Y(n_1172)
);

INVx4_ASAP7_75t_L g1173 ( 
.A(n_957),
.Y(n_1173)
);

OR2x6_ASAP7_75t_L g1174 ( 
.A(n_990),
.B(n_588),
.Y(n_1174)
);

NAND2xp5_ASAP7_75t_L g1175 ( 
.A(n_994),
.B(n_589),
.Y(n_1175)
);

A2O1A1Ixp33_ASAP7_75t_L g1176 ( 
.A1(n_932),
.A2(n_642),
.B(n_657),
.C(n_658),
.Y(n_1176)
);

NAND2xp5_ASAP7_75t_L g1177 ( 
.A(n_994),
.B(n_589),
.Y(n_1177)
);

NOR3xp33_ASAP7_75t_L g1178 ( 
.A(n_955),
.B(n_343),
.C(n_342),
.Y(n_1178)
);

OAI22xp5_ASAP7_75t_L g1179 ( 
.A1(n_983),
.A2(n_595),
.B1(n_598),
.B2(n_601),
.Y(n_1179)
);

AOI22xp33_ASAP7_75t_L g1180 ( 
.A1(n_876),
.A2(n_254),
.B1(n_668),
.B2(n_784),
.Y(n_1180)
);

BUFx6f_ASAP7_75t_L g1181 ( 
.A(n_983),
.Y(n_1181)
);

NOR2xp33_ASAP7_75t_L g1182 ( 
.A(n_830),
.B(n_349),
.Y(n_1182)
);

NAND2xp5_ASAP7_75t_L g1183 ( 
.A(n_920),
.B(n_595),
.Y(n_1183)
);

NAND2xp5_ASAP7_75t_L g1184 ( 
.A(n_945),
.B(n_598),
.Y(n_1184)
);

BUFx6f_ASAP7_75t_L g1185 ( 
.A(n_1091),
.Y(n_1185)
);

BUFx6f_ASAP7_75t_L g1186 ( 
.A(n_1091),
.Y(n_1186)
);

OAI21xp33_ASAP7_75t_SL g1187 ( 
.A1(n_1097),
.A2(n_976),
.B(n_952),
.Y(n_1187)
);

A2O1A1Ixp33_ASAP7_75t_L g1188 ( 
.A1(n_1065),
.A2(n_973),
.B(n_995),
.C(n_990),
.Y(n_1188)
);

CKINVDCx20_ASAP7_75t_R g1189 ( 
.A(n_1025),
.Y(n_1189)
);

BUFx2_ASAP7_75t_L g1190 ( 
.A(n_1007),
.Y(n_1190)
);

INVx2_ASAP7_75t_L g1191 ( 
.A(n_1034),
.Y(n_1191)
);

BUFx6f_ASAP7_75t_L g1192 ( 
.A(n_1091),
.Y(n_1192)
);

AOI21xp5_ASAP7_75t_L g1193 ( 
.A1(n_1002),
.A2(n_985),
.B(n_983),
.Y(n_1193)
);

OR2x2_ASAP7_75t_L g1194 ( 
.A(n_1009),
.B(n_1082),
.Y(n_1194)
);

NOR2xp33_ASAP7_75t_L g1195 ( 
.A(n_1069),
.B(n_1105),
.Y(n_1195)
);

OAI22xp5_ASAP7_75t_L g1196 ( 
.A1(n_1019),
.A2(n_1132),
.B1(n_1100),
.B2(n_1000),
.Y(n_1196)
);

INVx2_ASAP7_75t_L g1197 ( 
.A(n_1050),
.Y(n_1197)
);

OAI22xp5_ASAP7_75t_L g1198 ( 
.A1(n_1092),
.A2(n_894),
.B1(n_881),
.B2(n_976),
.Y(n_1198)
);

OAI22xp5_ASAP7_75t_L g1199 ( 
.A1(n_1105),
.A2(n_894),
.B1(n_996),
.B2(n_985),
.Y(n_1199)
);

NOR2x1_ASAP7_75t_SL g1200 ( 
.A(n_1110),
.B(n_983),
.Y(n_1200)
);

AOI21xp5_ASAP7_75t_L g1201 ( 
.A1(n_1002),
.A2(n_985),
.B(n_852),
.Y(n_1201)
);

NAND2xp5_ASAP7_75t_L g1202 ( 
.A(n_1096),
.B(n_972),
.Y(n_1202)
);

INVx1_ASAP7_75t_SL g1203 ( 
.A(n_1040),
.Y(n_1203)
);

AOI21xp5_ASAP7_75t_L g1204 ( 
.A1(n_1110),
.A2(n_985),
.B(n_852),
.Y(n_1204)
);

INVx2_ASAP7_75t_SL g1205 ( 
.A(n_1054),
.Y(n_1205)
);

BUFx3_ASAP7_75t_L g1206 ( 
.A(n_1073),
.Y(n_1206)
);

BUFx6f_ASAP7_75t_L g1207 ( 
.A(n_1181),
.Y(n_1207)
);

A2O1A1Ixp33_ASAP7_75t_L g1208 ( 
.A1(n_1118),
.A2(n_847),
.B(n_855),
.C(n_862),
.Y(n_1208)
);

INVx8_ASAP7_75t_L g1209 ( 
.A(n_1110),
.Y(n_1209)
);

AND2x4_ASAP7_75t_L g1210 ( 
.A(n_1073),
.B(n_1075),
.Y(n_1210)
);

INVx2_ASAP7_75t_L g1211 ( 
.A(n_1081),
.Y(n_1211)
);

O2A1O1Ixp5_ASAP7_75t_L g1212 ( 
.A1(n_1042),
.A2(n_1137),
.B(n_1001),
.C(n_1033),
.Y(n_1212)
);

BUFx2_ASAP7_75t_L g1213 ( 
.A(n_1015),
.Y(n_1213)
);

INVx3_ASAP7_75t_L g1214 ( 
.A(n_1063),
.Y(n_1214)
);

O2A1O1Ixp33_ASAP7_75t_L g1215 ( 
.A1(n_1020),
.A2(n_644),
.B(n_618),
.C(n_622),
.Y(n_1215)
);

AOI21xp5_ASAP7_75t_L g1216 ( 
.A1(n_1110),
.A2(n_856),
.B(n_855),
.Y(n_1216)
);

AOI22xp5_ASAP7_75t_L g1217 ( 
.A1(n_1149),
.A2(n_862),
.B1(n_856),
.B2(n_988),
.Y(n_1217)
);

AOI21xp5_ASAP7_75t_L g1218 ( 
.A1(n_1032),
.A2(n_988),
.B(n_997),
.Y(n_1218)
);

INVx4_ASAP7_75t_L g1219 ( 
.A(n_1056),
.Y(n_1219)
);

NOR2xp33_ASAP7_75t_SL g1220 ( 
.A(n_1113),
.B(n_988),
.Y(n_1220)
);

OAI22xp5_ASAP7_75t_L g1221 ( 
.A1(n_1130),
.A2(n_440),
.B1(n_253),
.B2(n_256),
.Y(n_1221)
);

INVx2_ASAP7_75t_L g1222 ( 
.A(n_1090),
.Y(n_1222)
);

INVx1_ASAP7_75t_SL g1223 ( 
.A(n_1098),
.Y(n_1223)
);

NAND2xp5_ASAP7_75t_L g1224 ( 
.A(n_1004),
.B(n_997),
.Y(n_1224)
);

NAND2xp33_ASAP7_75t_L g1225 ( 
.A(n_1056),
.B(n_988),
.Y(n_1225)
);

HB1xp67_ASAP7_75t_L g1226 ( 
.A(n_1114),
.Y(n_1226)
);

INVx1_ASAP7_75t_L g1227 ( 
.A(n_1028),
.Y(n_1227)
);

NAND2xp5_ASAP7_75t_L g1228 ( 
.A(n_1031),
.B(n_997),
.Y(n_1228)
);

AOI21xp5_ASAP7_75t_L g1229 ( 
.A1(n_1032),
.A2(n_988),
.B(n_600),
.Y(n_1229)
);

NAND2xp5_ASAP7_75t_L g1230 ( 
.A(n_1045),
.B(n_988),
.Y(n_1230)
);

AO32x1_ASAP7_75t_L g1231 ( 
.A1(n_1135),
.A2(n_638),
.A3(n_621),
.B1(n_613),
.B2(n_659),
.Y(n_1231)
);

AOI21xp5_ASAP7_75t_L g1232 ( 
.A1(n_1104),
.A2(n_600),
.B(n_584),
.Y(n_1232)
);

NAND2x1p5_ASAP7_75t_L g1233 ( 
.A(n_1155),
.B(n_1173),
.Y(n_1233)
);

NAND2xp5_ASAP7_75t_L g1234 ( 
.A(n_1060),
.B(n_601),
.Y(n_1234)
);

A2O1A1Ixp33_ASAP7_75t_L g1235 ( 
.A1(n_1126),
.A2(n_369),
.B(n_350),
.C(n_406),
.Y(n_1235)
);

NOR2xp67_ASAP7_75t_SL g1236 ( 
.A(n_1156),
.B(n_249),
.Y(n_1236)
);

AOI22xp5_ASAP7_75t_L g1237 ( 
.A1(n_1151),
.A2(n_628),
.B1(n_631),
.B2(n_618),
.Y(n_1237)
);

INVx2_ASAP7_75t_L g1238 ( 
.A(n_1128),
.Y(n_1238)
);

NAND2xp5_ASAP7_75t_L g1239 ( 
.A(n_1011),
.B(n_622),
.Y(n_1239)
);

AND2x4_ASAP7_75t_L g1240 ( 
.A(n_1073),
.B(n_116),
.Y(n_1240)
);

AND2x2_ASAP7_75t_L g1241 ( 
.A(n_1111),
.B(n_351),
.Y(n_1241)
);

NAND2xp5_ASAP7_75t_L g1242 ( 
.A(n_1012),
.B(n_630),
.Y(n_1242)
);

INVx1_ASAP7_75t_SL g1243 ( 
.A(n_1101),
.Y(n_1243)
);

BUFx6f_ASAP7_75t_L g1244 ( 
.A(n_1181),
.Y(n_1244)
);

BUFx2_ASAP7_75t_L g1245 ( 
.A(n_1064),
.Y(n_1245)
);

NOR2xp33_ASAP7_75t_L g1246 ( 
.A(n_1086),
.B(n_357),
.Y(n_1246)
);

OAI22xp5_ASAP7_75t_L g1247 ( 
.A1(n_1147),
.A2(n_443),
.B1(n_440),
.B2(n_434),
.Y(n_1247)
);

NAND2xp33_ASAP7_75t_SL g1248 ( 
.A(n_1075),
.B(n_253),
.Y(n_1248)
);

NOR3xp33_ASAP7_75t_SL g1249 ( 
.A(n_1017),
.B(n_1117),
.C(n_1150),
.Y(n_1249)
);

AOI21xp5_ASAP7_75t_L g1250 ( 
.A1(n_1104),
.A2(n_1027),
.B(n_1026),
.Y(n_1250)
);

BUFx12f_ASAP7_75t_L g1251 ( 
.A(n_1124),
.Y(n_1251)
);

O2A1O1Ixp5_ASAP7_75t_SL g1252 ( 
.A1(n_1163),
.A2(n_644),
.B(n_630),
.C(n_662),
.Y(n_1252)
);

A2O1A1Ixp33_ASAP7_75t_L g1253 ( 
.A1(n_1008),
.A2(n_401),
.B(n_396),
.C(n_395),
.Y(n_1253)
);

NAND2xp5_ASAP7_75t_L g1254 ( 
.A(n_1044),
.B(n_631),
.Y(n_1254)
);

AND2x6_ASAP7_75t_L g1255 ( 
.A(n_1013),
.B(n_613),
.Y(n_1255)
);

O2A1O1Ixp5_ASAP7_75t_L g1256 ( 
.A1(n_1051),
.A2(n_643),
.B(n_635),
.C(n_662),
.Y(n_1256)
);

AND2x6_ASAP7_75t_SL g1257 ( 
.A(n_1182),
.B(n_256),
.Y(n_1257)
);

INVxp67_ASAP7_75t_L g1258 ( 
.A(n_1043),
.Y(n_1258)
);

A2O1A1Ixp33_ASAP7_75t_L g1259 ( 
.A1(n_1008),
.A2(n_382),
.B(n_373),
.C(n_372),
.Y(n_1259)
);

AO22x1_ASAP7_75t_L g1260 ( 
.A1(n_1142),
.A2(n_430),
.B1(n_335),
.B2(n_407),
.Y(n_1260)
);

AOI21xp5_ASAP7_75t_L g1261 ( 
.A1(n_1026),
.A2(n_584),
.B(n_600),
.Y(n_1261)
);

BUFx6f_ASAP7_75t_L g1262 ( 
.A(n_1181),
.Y(n_1262)
);

O2A1O1Ixp33_ASAP7_75t_L g1263 ( 
.A1(n_1022),
.A2(n_1138),
.B(n_1129),
.C(n_1102),
.Y(n_1263)
);

NAND2xp5_ASAP7_75t_L g1264 ( 
.A(n_1103),
.B(n_635),
.Y(n_1264)
);

INVxp67_ASAP7_75t_L g1265 ( 
.A(n_1094),
.Y(n_1265)
);

NAND2xp5_ASAP7_75t_SL g1266 ( 
.A(n_1048),
.B(n_363),
.Y(n_1266)
);

INVx2_ASAP7_75t_L g1267 ( 
.A(n_1136),
.Y(n_1267)
);

INVx1_ASAP7_75t_L g1268 ( 
.A(n_1103),
.Y(n_1268)
);

NAND2xp5_ASAP7_75t_L g1269 ( 
.A(n_1016),
.B(n_642),
.Y(n_1269)
);

BUFx10_ASAP7_75t_L g1270 ( 
.A(n_1112),
.Y(n_1270)
);

INVx1_ASAP7_75t_L g1271 ( 
.A(n_1119),
.Y(n_1271)
);

O2A1O1Ixp33_ASAP7_75t_SL g1272 ( 
.A1(n_1176),
.A2(n_613),
.B(n_621),
.C(n_638),
.Y(n_1272)
);

O2A1O1Ixp33_ASAP7_75t_L g1273 ( 
.A1(n_1074),
.A2(n_659),
.B(n_658),
.C(n_657),
.Y(n_1273)
);

NOR2xp33_ASAP7_75t_L g1274 ( 
.A(n_1076),
.B(n_364),
.Y(n_1274)
);

HB1xp67_ASAP7_75t_L g1275 ( 
.A(n_1075),
.Y(n_1275)
);

NAND2xp5_ASAP7_75t_SL g1276 ( 
.A(n_1048),
.B(n_365),
.Y(n_1276)
);

NAND2xp5_ASAP7_75t_L g1277 ( 
.A(n_1006),
.B(n_643),
.Y(n_1277)
);

O2A1O1Ixp33_ASAP7_75t_L g1278 ( 
.A1(n_1168),
.A2(n_645),
.B(n_648),
.C(n_638),
.Y(n_1278)
);

HB1xp67_ASAP7_75t_L g1279 ( 
.A(n_1064),
.Y(n_1279)
);

NAND2xp5_ASAP7_75t_L g1280 ( 
.A(n_1095),
.B(n_645),
.Y(n_1280)
);

INVx1_ASAP7_75t_L g1281 ( 
.A(n_1120),
.Y(n_1281)
);

A2O1A1Ixp33_ASAP7_75t_L g1282 ( 
.A1(n_1106),
.A2(n_405),
.B(n_404),
.C(n_385),
.Y(n_1282)
);

AND2x4_ASAP7_75t_L g1283 ( 
.A(n_1112),
.B(n_119),
.Y(n_1283)
);

OAI21xp5_ASAP7_75t_L g1284 ( 
.A1(n_1024),
.A2(n_802),
.B(n_784),
.Y(n_1284)
);

AOI21xp5_ASAP7_75t_L g1285 ( 
.A1(n_1027),
.A2(n_584),
.B(n_600),
.Y(n_1285)
);

O2A1O1Ixp33_ASAP7_75t_L g1286 ( 
.A1(n_1172),
.A2(n_648),
.B(n_621),
.C(n_653),
.Y(n_1286)
);

INVx1_ASAP7_75t_L g1287 ( 
.A(n_1141),
.Y(n_1287)
);

AND2x2_ASAP7_75t_L g1288 ( 
.A(n_1068),
.B(n_394),
.Y(n_1288)
);

NAND2xp5_ASAP7_75t_L g1289 ( 
.A(n_1029),
.B(n_653),
.Y(n_1289)
);

AOI21xp5_ASAP7_75t_L g1290 ( 
.A1(n_1037),
.A2(n_600),
.B(n_655),
.Y(n_1290)
);

NAND2xp5_ASAP7_75t_L g1291 ( 
.A(n_1018),
.B(n_653),
.Y(n_1291)
);

AND2x2_ASAP7_75t_L g1292 ( 
.A(n_1068),
.B(n_402),
.Y(n_1292)
);

BUFx2_ASAP7_75t_L g1293 ( 
.A(n_1064),
.Y(n_1293)
);

NAND3xp33_ASAP7_75t_SL g1294 ( 
.A(n_1178),
.B(n_258),
.C(n_407),
.Y(n_1294)
);

INVx6_ASAP7_75t_L g1295 ( 
.A(n_1153),
.Y(n_1295)
);

NAND2xp5_ASAP7_75t_SL g1296 ( 
.A(n_1113),
.B(n_403),
.Y(n_1296)
);

NAND2xp5_ASAP7_75t_L g1297 ( 
.A(n_1021),
.B(n_653),
.Y(n_1297)
);

INVxp67_ASAP7_75t_L g1298 ( 
.A(n_1059),
.Y(n_1298)
);

OAI21xp33_ASAP7_75t_L g1299 ( 
.A1(n_1068),
.A2(n_420),
.B(n_430),
.Y(n_1299)
);

INVx2_ASAP7_75t_L g1300 ( 
.A(n_1139),
.Y(n_1300)
);

AOI22xp5_ASAP7_75t_L g1301 ( 
.A1(n_1057),
.A2(n_802),
.B1(n_784),
.B2(n_254),
.Y(n_1301)
);

OAI22xp5_ASAP7_75t_L g1302 ( 
.A1(n_1093),
.A2(n_443),
.B1(n_656),
.B2(n_655),
.Y(n_1302)
);

BUFx8_ASAP7_75t_L g1303 ( 
.A(n_1148),
.Y(n_1303)
);

BUFx3_ASAP7_75t_L g1304 ( 
.A(n_1165),
.Y(n_1304)
);

NAND2xp5_ASAP7_75t_L g1305 ( 
.A(n_1023),
.B(n_653),
.Y(n_1305)
);

BUFx3_ASAP7_75t_L g1306 ( 
.A(n_1164),
.Y(n_1306)
);

AOI21xp5_ASAP7_75t_L g1307 ( 
.A1(n_1037),
.A2(n_656),
.B(n_655),
.Y(n_1307)
);

CKINVDCx5p33_ASAP7_75t_R g1308 ( 
.A(n_1164),
.Y(n_1308)
);

INVx2_ASAP7_75t_L g1309 ( 
.A(n_1157),
.Y(n_1309)
);

NAND2xp5_ASAP7_75t_L g1310 ( 
.A(n_1061),
.B(n_1062),
.Y(n_1310)
);

A2O1A1Ixp33_ASAP7_75t_L g1311 ( 
.A1(n_1024),
.A2(n_656),
.B(n_655),
.C(n_610),
.Y(n_1311)
);

AOI21xp5_ASAP7_75t_L g1312 ( 
.A1(n_1067),
.A2(n_656),
.B(n_655),
.Y(n_1312)
);

NAND2xp5_ASAP7_75t_L g1313 ( 
.A(n_1035),
.B(n_656),
.Y(n_1313)
);

NAND2xp5_ASAP7_75t_L g1314 ( 
.A(n_1160),
.B(n_668),
.Y(n_1314)
);

NAND2xp5_ASAP7_75t_L g1315 ( 
.A(n_1071),
.B(n_668),
.Y(n_1315)
);

NAND2xp5_ASAP7_75t_SL g1316 ( 
.A(n_1057),
.B(n_254),
.Y(n_1316)
);

INVx4_ASAP7_75t_L g1317 ( 
.A(n_1155),
.Y(n_1317)
);

O2A1O1Ixp33_ASAP7_75t_L g1318 ( 
.A1(n_1046),
.A2(n_610),
.B(n_608),
.C(n_22),
.Y(n_1318)
);

NOR3xp33_ASAP7_75t_SL g1319 ( 
.A(n_1072),
.B(n_14),
.C(n_18),
.Y(n_1319)
);

AOI21xp5_ASAP7_75t_L g1320 ( 
.A1(n_1066),
.A2(n_610),
.B(n_608),
.Y(n_1320)
);

OAI21xp5_ASAP7_75t_L g1321 ( 
.A1(n_1116),
.A2(n_802),
.B(n_784),
.Y(n_1321)
);

OAI21xp33_ASAP7_75t_SL g1322 ( 
.A1(n_1099),
.A2(n_18),
.B(n_23),
.Y(n_1322)
);

AOI22xp5_ASAP7_75t_L g1323 ( 
.A1(n_1109),
.A2(n_802),
.B1(n_784),
.B2(n_254),
.Y(n_1323)
);

AOI21xp5_ASAP7_75t_L g1324 ( 
.A1(n_1038),
.A2(n_610),
.B(n_608),
.Y(n_1324)
);

INVx1_ASAP7_75t_L g1325 ( 
.A(n_1169),
.Y(n_1325)
);

NAND2xp5_ASAP7_75t_SL g1326 ( 
.A(n_1109),
.B(n_668),
.Y(n_1326)
);

NOR2xp33_ASAP7_75t_L g1327 ( 
.A(n_1003),
.B(n_25),
.Y(n_1327)
);

OAI22xp5_ASAP7_75t_L g1328 ( 
.A1(n_1077),
.A2(n_668),
.B1(n_610),
.B2(n_608),
.Y(n_1328)
);

INVx3_ASAP7_75t_L g1329 ( 
.A(n_1063),
.Y(n_1329)
);

O2A1O1Ixp33_ASAP7_75t_L g1330 ( 
.A1(n_1046),
.A2(n_608),
.B(n_27),
.C(n_31),
.Y(n_1330)
);

AOI21xp5_ASAP7_75t_L g1331 ( 
.A1(n_1038),
.A2(n_668),
.B(n_802),
.Y(n_1331)
);

OAI22xp5_ASAP7_75t_L g1332 ( 
.A1(n_1078),
.A2(n_668),
.B1(n_27),
.B2(n_32),
.Y(n_1332)
);

NAND2xp5_ASAP7_75t_L g1333 ( 
.A(n_998),
.B(n_668),
.Y(n_1333)
);

BUFx12f_ASAP7_75t_L g1334 ( 
.A(n_1173),
.Y(n_1334)
);

O2A1O1Ixp33_ASAP7_75t_L g1335 ( 
.A1(n_1036),
.A2(n_25),
.B(n_32),
.C(n_33),
.Y(n_1335)
);

INVx1_ASAP7_75t_L g1336 ( 
.A(n_1183),
.Y(n_1336)
);

AND2x2_ASAP7_75t_L g1337 ( 
.A(n_1170),
.B(n_35),
.Y(n_1337)
);

BUFx6f_ASAP7_75t_L g1338 ( 
.A(n_999),
.Y(n_1338)
);

NAND2xp5_ASAP7_75t_L g1339 ( 
.A(n_999),
.B(n_802),
.Y(n_1339)
);

AOI21xp5_ASAP7_75t_L g1340 ( 
.A1(n_1116),
.A2(n_784),
.B(n_229),
.Y(n_1340)
);

OAI22xp5_ASAP7_75t_L g1341 ( 
.A1(n_1079),
.A2(n_35),
.B1(n_38),
.B2(n_39),
.Y(n_1341)
);

INVx4_ASAP7_75t_L g1342 ( 
.A(n_1014),
.Y(n_1342)
);

AND2x2_ASAP7_75t_L g1343 ( 
.A(n_1014),
.B(n_42),
.Y(n_1343)
);

NAND2xp33_ASAP7_75t_SL g1344 ( 
.A(n_1030),
.B(n_1140),
.Y(n_1344)
);

OAI22xp5_ASAP7_75t_L g1345 ( 
.A1(n_1080),
.A2(n_43),
.B1(n_45),
.B2(n_46),
.Y(n_1345)
);

NAND3xp33_ASAP7_75t_SL g1346 ( 
.A(n_1246),
.B(n_1058),
.C(n_1005),
.Y(n_1346)
);

BUFx12f_ASAP7_75t_L g1347 ( 
.A(n_1308),
.Y(n_1347)
);

OAI22x1_ASAP7_75t_L g1348 ( 
.A1(n_1195),
.A2(n_1152),
.B1(n_1030),
.B2(n_1041),
.Y(n_1348)
);

AO31x2_ASAP7_75t_L g1349 ( 
.A1(n_1250),
.A2(n_1179),
.A3(n_1089),
.B(n_1055),
.Y(n_1349)
);

BUFx2_ASAP7_75t_L g1350 ( 
.A(n_1190),
.Y(n_1350)
);

AOI21xp5_ASAP7_75t_L g1351 ( 
.A1(n_1310),
.A2(n_1107),
.B(n_1010),
.Y(n_1351)
);

NAND2xp5_ASAP7_75t_L g1352 ( 
.A(n_1336),
.B(n_1196),
.Y(n_1352)
);

AO31x2_ASAP7_75t_L g1353 ( 
.A1(n_1218),
.A2(n_1089),
.A3(n_1055),
.B(n_1084),
.Y(n_1353)
);

AND2x2_ASAP7_75t_SL g1354 ( 
.A(n_1220),
.B(n_1152),
.Y(n_1354)
);

AND2x2_ASAP7_75t_SL g1355 ( 
.A(n_1220),
.B(n_1088),
.Y(n_1355)
);

AOI221x1_ASAP7_75t_L g1356 ( 
.A1(n_1196),
.A2(n_1084),
.B1(n_1070),
.B2(n_1115),
.C(n_1049),
.Y(n_1356)
);

NAND3xp33_ASAP7_75t_L g1357 ( 
.A(n_1249),
.B(n_1274),
.C(n_1263),
.Y(n_1357)
);

CKINVDCx8_ASAP7_75t_R g1358 ( 
.A(n_1257),
.Y(n_1358)
);

NAND3xp33_ASAP7_75t_SL g1359 ( 
.A(n_1194),
.B(n_1154),
.C(n_1127),
.Y(n_1359)
);

AND2x2_ASAP7_75t_L g1360 ( 
.A(n_1243),
.B(n_1174),
.Y(n_1360)
);

NAND2xp5_ASAP7_75t_L g1361 ( 
.A(n_1202),
.B(n_1108),
.Y(n_1361)
);

INVx5_ASAP7_75t_L g1362 ( 
.A(n_1209),
.Y(n_1362)
);

AO31x2_ASAP7_75t_L g1363 ( 
.A1(n_1302),
.A2(n_1070),
.A3(n_1049),
.B(n_1047),
.Y(n_1363)
);

A2O1A1Ixp33_ASAP7_75t_L g1364 ( 
.A1(n_1212),
.A2(n_1144),
.B(n_1146),
.C(n_1159),
.Y(n_1364)
);

NAND2xp5_ASAP7_75t_SL g1365 ( 
.A(n_1203),
.B(n_1134),
.Y(n_1365)
);

AOI21xp5_ASAP7_75t_L g1366 ( 
.A1(n_1193),
.A2(n_1083),
.B(n_1087),
.Y(n_1366)
);

INVx3_ASAP7_75t_L g1367 ( 
.A(n_1209),
.Y(n_1367)
);

O2A1O1Ixp33_ASAP7_75t_L g1368 ( 
.A1(n_1235),
.A2(n_1159),
.B(n_1184),
.C(n_1177),
.Y(n_1368)
);

OAI21xp5_ASAP7_75t_L g1369 ( 
.A1(n_1187),
.A2(n_1047),
.B(n_1085),
.Y(n_1369)
);

AOI21x1_ASAP7_75t_L g1370 ( 
.A1(n_1232),
.A2(n_1161),
.B(n_1175),
.Y(n_1370)
);

BUFx2_ASAP7_75t_L g1371 ( 
.A(n_1213),
.Y(n_1371)
);

OA21x2_ASAP7_75t_L g1372 ( 
.A1(n_1256),
.A2(n_1166),
.B(n_1121),
.Y(n_1372)
);

AO32x2_ASAP7_75t_L g1373 ( 
.A1(n_1332),
.A2(n_1174),
.A3(n_1167),
.B1(n_1145),
.B2(n_1144),
.Y(n_1373)
);

BUFx2_ASAP7_75t_L g1374 ( 
.A(n_1205),
.Y(n_1374)
);

A2O1A1Ixp33_ASAP7_75t_L g1375 ( 
.A1(n_1253),
.A2(n_1259),
.B(n_1198),
.C(n_1282),
.Y(n_1375)
);

NAND2xp5_ASAP7_75t_L g1376 ( 
.A(n_1239),
.B(n_1146),
.Y(n_1376)
);

NAND2xp5_ASAP7_75t_L g1377 ( 
.A(n_1243),
.B(n_1174),
.Y(n_1377)
);

NAND2xp5_ASAP7_75t_L g1378 ( 
.A(n_1268),
.B(n_1052),
.Y(n_1378)
);

INVxp67_ASAP7_75t_SL g1379 ( 
.A(n_1200),
.Y(n_1379)
);

CKINVDCx5p33_ASAP7_75t_R g1380 ( 
.A(n_1189),
.Y(n_1380)
);

NOR2xp67_ASAP7_75t_L g1381 ( 
.A(n_1298),
.B(n_1052),
.Y(n_1381)
);

NAND2xp5_ASAP7_75t_L g1382 ( 
.A(n_1242),
.B(n_1053),
.Y(n_1382)
);

AOI21xp5_ASAP7_75t_L g1383 ( 
.A1(n_1277),
.A2(n_1039),
.B(n_1053),
.Y(n_1383)
);

OAI22xp5_ASAP7_75t_L g1384 ( 
.A1(n_1198),
.A2(n_1145),
.B1(n_1122),
.B2(n_1180),
.Y(n_1384)
);

OAI21x1_ASAP7_75t_L g1385 ( 
.A1(n_1261),
.A2(n_1133),
.B(n_1162),
.Y(n_1385)
);

AOI21xp5_ASAP7_75t_L g1386 ( 
.A1(n_1277),
.A2(n_1188),
.B(n_1225),
.Y(n_1386)
);

NAND2xp5_ASAP7_75t_L g1387 ( 
.A(n_1254),
.B(n_1269),
.Y(n_1387)
);

CKINVDCx6p67_ASAP7_75t_R g1388 ( 
.A(n_1306),
.Y(n_1388)
);

AOI21xp5_ASAP7_75t_L g1389 ( 
.A1(n_1291),
.A2(n_1123),
.B(n_1125),
.Y(n_1389)
);

OAI21x1_ASAP7_75t_L g1390 ( 
.A1(n_1285),
.A2(n_1133),
.B(n_1162),
.Y(n_1390)
);

OAI21x1_ASAP7_75t_L g1391 ( 
.A1(n_1229),
.A2(n_1171),
.B(n_1131),
.Y(n_1391)
);

AOI21xp5_ASAP7_75t_L g1392 ( 
.A1(n_1297),
.A2(n_1305),
.B(n_1289),
.Y(n_1392)
);

O2A1O1Ixp33_ASAP7_75t_L g1393 ( 
.A1(n_1294),
.A2(n_1131),
.B(n_1125),
.C(n_1123),
.Y(n_1393)
);

AO31x2_ASAP7_75t_L g1394 ( 
.A1(n_1302),
.A2(n_1171),
.A3(n_1158),
.B(n_1143),
.Y(n_1394)
);

INVx3_ASAP7_75t_SL g1395 ( 
.A(n_1295),
.Y(n_1395)
);

CKINVDCx5p33_ASAP7_75t_R g1396 ( 
.A(n_1251),
.Y(n_1396)
);

AOI21xp5_ASAP7_75t_L g1397 ( 
.A1(n_1340),
.A2(n_1158),
.B(n_1143),
.Y(n_1397)
);

BUFx3_ASAP7_75t_L g1398 ( 
.A(n_1304),
.Y(n_1398)
);

AO31x2_ASAP7_75t_L g1399 ( 
.A1(n_1311),
.A2(n_43),
.A3(n_45),
.B(n_46),
.Y(n_1399)
);

O2A1O1Ixp33_ASAP7_75t_L g1400 ( 
.A1(n_1258),
.A2(n_47),
.B(n_50),
.C(n_53),
.Y(n_1400)
);

NAND2xp5_ASAP7_75t_L g1401 ( 
.A(n_1271),
.B(n_47),
.Y(n_1401)
);

OAI21x1_ASAP7_75t_L g1402 ( 
.A1(n_1290),
.A2(n_133),
.B(n_222),
.Y(n_1402)
);

BUFx3_ASAP7_75t_L g1403 ( 
.A(n_1206),
.Y(n_1403)
);

AOI221x1_ASAP7_75t_L g1404 ( 
.A1(n_1332),
.A2(n_50),
.B1(n_53),
.B2(n_56),
.C(n_57),
.Y(n_1404)
);

AO31x2_ASAP7_75t_L g1405 ( 
.A1(n_1331),
.A2(n_58),
.A3(n_59),
.B(n_60),
.Y(n_1405)
);

AOI21xp5_ASAP7_75t_L g1406 ( 
.A1(n_1313),
.A2(n_1208),
.B(n_1315),
.Y(n_1406)
);

OAI22xp5_ASAP7_75t_L g1407 ( 
.A1(n_1203),
.A2(n_61),
.B1(n_64),
.B2(n_67),
.Y(n_1407)
);

HB1xp67_ASAP7_75t_L g1408 ( 
.A(n_1223),
.Y(n_1408)
);

AOI211x1_ASAP7_75t_L g1409 ( 
.A1(n_1260),
.A2(n_68),
.B(n_69),
.C(n_70),
.Y(n_1409)
);

INVx1_ASAP7_75t_L g1410 ( 
.A(n_1281),
.Y(n_1410)
);

NOR2xp33_ASAP7_75t_L g1411 ( 
.A(n_1223),
.B(n_71),
.Y(n_1411)
);

AO31x2_ASAP7_75t_L g1412 ( 
.A1(n_1224),
.A2(n_72),
.A3(n_73),
.B(n_76),
.Y(n_1412)
);

AO21x2_ASAP7_75t_L g1413 ( 
.A1(n_1321),
.A2(n_157),
.B(n_221),
.Y(n_1413)
);

AOI21xp5_ASAP7_75t_L g1414 ( 
.A1(n_1209),
.A2(n_153),
.B(n_220),
.Y(n_1414)
);

AO31x2_ASAP7_75t_L g1415 ( 
.A1(n_1228),
.A2(n_78),
.A3(n_79),
.B(n_80),
.Y(n_1415)
);

AOI21xp5_ASAP7_75t_L g1416 ( 
.A1(n_1321),
.A2(n_162),
.B(n_212),
.Y(n_1416)
);

INVx1_ASAP7_75t_L g1417 ( 
.A(n_1287),
.Y(n_1417)
);

INVx1_ASAP7_75t_L g1418 ( 
.A(n_1325),
.Y(n_1418)
);

O2A1O1Ixp33_ASAP7_75t_SL g1419 ( 
.A1(n_1230),
.A2(n_158),
.B(n_211),
.C(n_208),
.Y(n_1419)
);

AO31x2_ASAP7_75t_L g1420 ( 
.A1(n_1199),
.A2(n_81),
.A3(n_82),
.B(n_84),
.Y(n_1420)
);

OAI21x1_ASAP7_75t_L g1421 ( 
.A1(n_1307),
.A2(n_125),
.B(n_127),
.Y(n_1421)
);

OAI21xp5_ASAP7_75t_L g1422 ( 
.A1(n_1312),
.A2(n_136),
.B(n_137),
.Y(n_1422)
);

O2A1O1Ixp33_ASAP7_75t_SL g1423 ( 
.A1(n_1316),
.A2(n_140),
.B(n_141),
.C(n_143),
.Y(n_1423)
);

AOI22xp33_ASAP7_75t_L g1424 ( 
.A1(n_1337),
.A2(n_146),
.B1(n_165),
.B2(n_166),
.Y(n_1424)
);

NAND2xp5_ASAP7_75t_L g1425 ( 
.A(n_1191),
.B(n_180),
.Y(n_1425)
);

NOR3xp33_ASAP7_75t_L g1426 ( 
.A(n_1296),
.B(n_1266),
.C(n_1276),
.Y(n_1426)
);

OAI21xp5_ASAP7_75t_L g1427 ( 
.A1(n_1252),
.A2(n_1320),
.B(n_1324),
.Y(n_1427)
);

OAI22xp5_ASAP7_75t_L g1428 ( 
.A1(n_1264),
.A2(n_186),
.B1(n_192),
.B2(n_200),
.Y(n_1428)
);

NAND2xp5_ASAP7_75t_L g1429 ( 
.A(n_1197),
.B(n_203),
.Y(n_1429)
);

AOI21xp5_ASAP7_75t_L g1430 ( 
.A1(n_1284),
.A2(n_1214),
.B(n_1329),
.Y(n_1430)
);

AND2x2_ASAP7_75t_L g1431 ( 
.A(n_1241),
.B(n_224),
.Y(n_1431)
);

BUFx6f_ASAP7_75t_L g1432 ( 
.A(n_1185),
.Y(n_1432)
);

NAND3xp33_ASAP7_75t_L g1433 ( 
.A(n_1322),
.B(n_1330),
.C(n_1319),
.Y(n_1433)
);

INVx2_ASAP7_75t_SL g1434 ( 
.A(n_1210),
.Y(n_1434)
);

INVx5_ASAP7_75t_L g1435 ( 
.A(n_1185),
.Y(n_1435)
);

BUFx3_ASAP7_75t_L g1436 ( 
.A(n_1210),
.Y(n_1436)
);

INVx1_ASAP7_75t_L g1437 ( 
.A(n_1211),
.Y(n_1437)
);

OAI21x1_ASAP7_75t_L g1438 ( 
.A1(n_1314),
.A2(n_1284),
.B(n_1333),
.Y(n_1438)
);

O2A1O1Ixp33_ASAP7_75t_SL g1439 ( 
.A1(n_1199),
.A2(n_1217),
.B(n_1326),
.C(n_1318),
.Y(n_1439)
);

NAND2xp5_ASAP7_75t_L g1440 ( 
.A(n_1222),
.B(n_1300),
.Y(n_1440)
);

INVx1_ASAP7_75t_L g1441 ( 
.A(n_1238),
.Y(n_1441)
);

NAND2xp5_ASAP7_75t_L g1442 ( 
.A(n_1267),
.B(n_1309),
.Y(n_1442)
);

AOI221xp5_ASAP7_75t_SL g1443 ( 
.A1(n_1345),
.A2(n_1341),
.B1(n_1335),
.B2(n_1247),
.C(n_1221),
.Y(n_1443)
);

OAI21x1_ASAP7_75t_L g1444 ( 
.A1(n_1314),
.A2(n_1204),
.B(n_1216),
.Y(n_1444)
);

AND2x6_ASAP7_75t_L g1445 ( 
.A(n_1240),
.B(n_1283),
.Y(n_1445)
);

AOI21xp33_ASAP7_75t_L g1446 ( 
.A1(n_1345),
.A2(n_1341),
.B(n_1278),
.Y(n_1446)
);

OAI22x1_ASAP7_75t_L g1447 ( 
.A1(n_1279),
.A2(n_1245),
.B1(n_1293),
.B2(n_1327),
.Y(n_1447)
);

INVx3_ASAP7_75t_L g1448 ( 
.A(n_1338),
.Y(n_1448)
);

OAI21x1_ASAP7_75t_L g1449 ( 
.A1(n_1328),
.A2(n_1286),
.B(n_1329),
.Y(n_1449)
);

INVx5_ASAP7_75t_L g1450 ( 
.A(n_1185),
.Y(n_1450)
);

AOI21xp5_ASAP7_75t_L g1451 ( 
.A1(n_1344),
.A2(n_1234),
.B(n_1280),
.Y(n_1451)
);

AO31x2_ASAP7_75t_L g1452 ( 
.A1(n_1328),
.A2(n_1231),
.A3(n_1339),
.B(n_1342),
.Y(n_1452)
);

AOI221x1_ASAP7_75t_L g1453 ( 
.A1(n_1299),
.A2(n_1221),
.B1(n_1247),
.B2(n_1248),
.C(n_1343),
.Y(n_1453)
);

OAI22xp5_ASAP7_75t_L g1454 ( 
.A1(n_1283),
.A2(n_1240),
.B1(n_1237),
.B2(n_1233),
.Y(n_1454)
);

BUFx3_ASAP7_75t_L g1455 ( 
.A(n_1303),
.Y(n_1455)
);

NAND2xp5_ASAP7_75t_L g1456 ( 
.A(n_1255),
.B(n_1338),
.Y(n_1456)
);

INVx1_ASAP7_75t_L g1457 ( 
.A(n_1226),
.Y(n_1457)
);

INVx5_ASAP7_75t_L g1458 ( 
.A(n_1186),
.Y(n_1458)
);

CKINVDCx9p33_ASAP7_75t_R g1459 ( 
.A(n_1334),
.Y(n_1459)
);

OAI21x1_ASAP7_75t_L g1460 ( 
.A1(n_1233),
.A2(n_1273),
.B(n_1215),
.Y(n_1460)
);

A2O1A1Ixp33_ASAP7_75t_L g1461 ( 
.A1(n_1265),
.A2(n_1292),
.B(n_1288),
.C(n_1236),
.Y(n_1461)
);

NAND2xp5_ASAP7_75t_L g1462 ( 
.A(n_1255),
.B(n_1338),
.Y(n_1462)
);

AOI21xp5_ASAP7_75t_L g1463 ( 
.A1(n_1231),
.A2(n_1272),
.B(n_1342),
.Y(n_1463)
);

AOI221x1_ASAP7_75t_L g1464 ( 
.A1(n_1231),
.A2(n_1186),
.B1(n_1192),
.B2(n_1207),
.C(n_1262),
.Y(n_1464)
);

NAND2xp5_ASAP7_75t_L g1465 ( 
.A(n_1255),
.B(n_1219),
.Y(n_1465)
);

BUFx6f_ASAP7_75t_L g1466 ( 
.A(n_1186),
.Y(n_1466)
);

INVx3_ASAP7_75t_L g1467 ( 
.A(n_1317),
.Y(n_1467)
);

OAI21x1_ASAP7_75t_L g1468 ( 
.A1(n_1301),
.A2(n_1323),
.B(n_1275),
.Y(n_1468)
);

NAND2xp5_ASAP7_75t_L g1469 ( 
.A(n_1219),
.B(n_1192),
.Y(n_1469)
);

AO21x2_ASAP7_75t_L g1470 ( 
.A1(n_1192),
.A2(n_1207),
.B(n_1244),
.Y(n_1470)
);

AO32x2_ASAP7_75t_L g1471 ( 
.A1(n_1270),
.A2(n_1196),
.A3(n_1332),
.B1(n_1147),
.B2(n_1135),
.Y(n_1471)
);

OAI21xp5_ASAP7_75t_L g1472 ( 
.A1(n_1270),
.A2(n_1244),
.B(n_1262),
.Y(n_1472)
);

INVx5_ASAP7_75t_L g1473 ( 
.A(n_1295),
.Y(n_1473)
);

O2A1O1Ixp33_ASAP7_75t_L g1474 ( 
.A1(n_1246),
.A2(n_904),
.B(n_1065),
.C(n_619),
.Y(n_1474)
);

AOI21xp5_ASAP7_75t_L g1475 ( 
.A1(n_1250),
.A2(n_904),
.B(n_1002),
.Y(n_1475)
);

INVx2_ASAP7_75t_L g1476 ( 
.A(n_1227),
.Y(n_1476)
);

INVx1_ASAP7_75t_SL g1477 ( 
.A(n_1203),
.Y(n_1477)
);

AOI21xp5_ASAP7_75t_L g1478 ( 
.A1(n_1250),
.A2(n_904),
.B(n_1002),
.Y(n_1478)
);

AOI21xp5_ASAP7_75t_L g1479 ( 
.A1(n_1250),
.A2(n_904),
.B(n_1002),
.Y(n_1479)
);

OR2x2_ASAP7_75t_L g1480 ( 
.A(n_1203),
.B(n_1243),
.Y(n_1480)
);

A2O1A1Ixp33_ASAP7_75t_L g1481 ( 
.A1(n_1263),
.A2(n_904),
.B(n_1092),
.C(n_1065),
.Y(n_1481)
);

OAI21x1_ASAP7_75t_L g1482 ( 
.A1(n_1201),
.A2(n_1193),
.B(n_1218),
.Y(n_1482)
);

OAI21x1_ASAP7_75t_L g1483 ( 
.A1(n_1201),
.A2(n_1193),
.B(n_1218),
.Y(n_1483)
);

INVx3_ASAP7_75t_L g1484 ( 
.A(n_1209),
.Y(n_1484)
);

AOI221xp5_ASAP7_75t_SL g1485 ( 
.A1(n_1196),
.A2(n_1065),
.B1(n_904),
.B2(n_892),
.C(n_1345),
.Y(n_1485)
);

INVx4_ASAP7_75t_L g1486 ( 
.A(n_1209),
.Y(n_1486)
);

OR2x2_ASAP7_75t_L g1487 ( 
.A(n_1203),
.B(n_1243),
.Y(n_1487)
);

AOI21x1_ASAP7_75t_L g1488 ( 
.A1(n_1218),
.A2(n_1193),
.B(n_1250),
.Y(n_1488)
);

AOI21xp5_ASAP7_75t_L g1489 ( 
.A1(n_1250),
.A2(n_904),
.B(n_1002),
.Y(n_1489)
);

INVx1_ASAP7_75t_L g1490 ( 
.A(n_1227),
.Y(n_1490)
);

NAND2xp5_ASAP7_75t_L g1491 ( 
.A(n_1336),
.B(n_904),
.Y(n_1491)
);

OAI21x1_ASAP7_75t_L g1492 ( 
.A1(n_1201),
.A2(n_1193),
.B(n_1218),
.Y(n_1492)
);

BUFx6f_ASAP7_75t_L g1493 ( 
.A(n_1185),
.Y(n_1493)
);

NAND2xp5_ASAP7_75t_SL g1494 ( 
.A(n_1203),
.B(n_904),
.Y(n_1494)
);

OAI21xp5_ASAP7_75t_L g1495 ( 
.A1(n_1212),
.A2(n_904),
.B(n_1187),
.Y(n_1495)
);

O2A1O1Ixp33_ASAP7_75t_L g1496 ( 
.A1(n_1246),
.A2(n_904),
.B(n_1065),
.C(n_619),
.Y(n_1496)
);

OAI21x1_ASAP7_75t_L g1497 ( 
.A1(n_1201),
.A2(n_1193),
.B(n_1218),
.Y(n_1497)
);

OAI21xp5_ASAP7_75t_L g1498 ( 
.A1(n_1212),
.A2(n_904),
.B(n_1187),
.Y(n_1498)
);

BUFx6f_ASAP7_75t_L g1499 ( 
.A(n_1185),
.Y(n_1499)
);

AND2x2_ASAP7_75t_L g1500 ( 
.A(n_1243),
.B(n_1009),
.Y(n_1500)
);

AOI21xp5_ASAP7_75t_L g1501 ( 
.A1(n_1250),
.A2(n_904),
.B(n_1002),
.Y(n_1501)
);

AOI21xp33_ASAP7_75t_L g1502 ( 
.A1(n_1246),
.A2(n_904),
.B(n_1118),
.Y(n_1502)
);

INVx2_ASAP7_75t_SL g1503 ( 
.A(n_1190),
.Y(n_1503)
);

NAND2xp5_ASAP7_75t_L g1504 ( 
.A(n_1336),
.B(n_904),
.Y(n_1504)
);

INVx1_ASAP7_75t_L g1505 ( 
.A(n_1227),
.Y(n_1505)
);

AO31x2_ASAP7_75t_L g1506 ( 
.A1(n_1250),
.A2(n_1218),
.A3(n_1135),
.B(n_1147),
.Y(n_1506)
);

NOR2xp33_ASAP7_75t_L g1507 ( 
.A(n_1194),
.B(n_904),
.Y(n_1507)
);

AOI22xp33_ASAP7_75t_L g1508 ( 
.A1(n_1246),
.A2(n_904),
.B1(n_1065),
.B2(n_1118),
.Y(n_1508)
);

AOI221x1_ASAP7_75t_L g1509 ( 
.A1(n_1196),
.A2(n_904),
.B1(n_1250),
.B2(n_1332),
.C(n_1065),
.Y(n_1509)
);

INVx2_ASAP7_75t_L g1510 ( 
.A(n_1227),
.Y(n_1510)
);

OAI21xp5_ASAP7_75t_L g1511 ( 
.A1(n_1212),
.A2(n_904),
.B(n_1187),
.Y(n_1511)
);

NAND2xp5_ASAP7_75t_SL g1512 ( 
.A(n_1203),
.B(n_904),
.Y(n_1512)
);

BUFx3_ASAP7_75t_L g1513 ( 
.A(n_1190),
.Y(n_1513)
);

OAI21x1_ASAP7_75t_L g1514 ( 
.A1(n_1201),
.A2(n_1193),
.B(n_1218),
.Y(n_1514)
);

BUFx6f_ASAP7_75t_L g1515 ( 
.A(n_1185),
.Y(n_1515)
);

HB1xp67_ASAP7_75t_L g1516 ( 
.A(n_1213),
.Y(n_1516)
);

BUFx2_ASAP7_75t_L g1517 ( 
.A(n_1513),
.Y(n_1517)
);

BUFx12f_ASAP7_75t_L g1518 ( 
.A(n_1396),
.Y(n_1518)
);

BUFx6f_ASAP7_75t_L g1519 ( 
.A(n_1435),
.Y(n_1519)
);

INVx1_ASAP7_75t_L g1520 ( 
.A(n_1510),
.Y(n_1520)
);

CKINVDCx5p33_ASAP7_75t_R g1521 ( 
.A(n_1380),
.Y(n_1521)
);

AOI22xp33_ASAP7_75t_L g1522 ( 
.A1(n_1508),
.A2(n_1502),
.B1(n_1357),
.B2(n_1446),
.Y(n_1522)
);

AOI22xp33_ASAP7_75t_L g1523 ( 
.A1(n_1502),
.A2(n_1357),
.B1(n_1446),
.B2(n_1507),
.Y(n_1523)
);

OAI22xp33_ASAP7_75t_L g1524 ( 
.A1(n_1404),
.A2(n_1491),
.B1(n_1504),
.B2(n_1407),
.Y(n_1524)
);

AOI22xp33_ASAP7_75t_L g1525 ( 
.A1(n_1407),
.A2(n_1433),
.B1(n_1352),
.B2(n_1491),
.Y(n_1525)
);

OAI22xp5_ASAP7_75t_L g1526 ( 
.A1(n_1504),
.A2(n_1481),
.B1(n_1496),
.B2(n_1474),
.Y(n_1526)
);

AOI22xp5_ASAP7_75t_SL g1527 ( 
.A1(n_1445),
.A2(n_1447),
.B1(n_1411),
.B2(n_1454),
.Y(n_1527)
);

NAND2x1p5_ASAP7_75t_L g1528 ( 
.A(n_1362),
.B(n_1435),
.Y(n_1528)
);

NAND2xp5_ASAP7_75t_L g1529 ( 
.A(n_1445),
.B(n_1387),
.Y(n_1529)
);

OAI22xp33_ASAP7_75t_L g1530 ( 
.A1(n_1453),
.A2(n_1352),
.B1(n_1387),
.B2(n_1509),
.Y(n_1530)
);

NAND2xp5_ASAP7_75t_L g1531 ( 
.A(n_1445),
.B(n_1494),
.Y(n_1531)
);

NAND2x1p5_ASAP7_75t_L g1532 ( 
.A(n_1362),
.B(n_1450),
.Y(n_1532)
);

BUFx2_ASAP7_75t_L g1533 ( 
.A(n_1371),
.Y(n_1533)
);

INVxp67_ASAP7_75t_SL g1534 ( 
.A(n_1376),
.Y(n_1534)
);

AOI22xp33_ASAP7_75t_SL g1535 ( 
.A1(n_1431),
.A2(n_1433),
.B1(n_1428),
.B2(n_1511),
.Y(n_1535)
);

BUFx3_ASAP7_75t_L g1536 ( 
.A(n_1403),
.Y(n_1536)
);

AOI22xp33_ASAP7_75t_L g1537 ( 
.A1(n_1512),
.A2(n_1511),
.B1(n_1498),
.B2(n_1495),
.Y(n_1537)
);

INVx6_ASAP7_75t_L g1538 ( 
.A(n_1473),
.Y(n_1538)
);

OAI22xp33_ASAP7_75t_L g1539 ( 
.A1(n_1477),
.A2(n_1487),
.B1(n_1480),
.B2(n_1401),
.Y(n_1539)
);

BUFx4f_ASAP7_75t_SL g1540 ( 
.A(n_1347),
.Y(n_1540)
);

OAI22xp33_ASAP7_75t_L g1541 ( 
.A1(n_1401),
.A2(n_1377),
.B1(n_1408),
.B2(n_1361),
.Y(n_1541)
);

OAI22xp33_ASAP7_75t_L g1542 ( 
.A1(n_1361),
.A2(n_1495),
.B1(n_1498),
.B2(n_1505),
.Y(n_1542)
);

AOI22xp33_ASAP7_75t_SL g1543 ( 
.A1(n_1428),
.A2(n_1422),
.B1(n_1384),
.B2(n_1360),
.Y(n_1543)
);

BUFx3_ASAP7_75t_L g1544 ( 
.A(n_1398),
.Y(n_1544)
);

AOI22xp33_ASAP7_75t_SL g1545 ( 
.A1(n_1422),
.A2(n_1384),
.B1(n_1473),
.B2(n_1355),
.Y(n_1545)
);

AOI22xp33_ASAP7_75t_L g1546 ( 
.A1(n_1346),
.A2(n_1426),
.B1(n_1359),
.B2(n_1376),
.Y(n_1546)
);

AOI21xp5_ASAP7_75t_L g1547 ( 
.A1(n_1475),
.A2(n_1479),
.B(n_1478),
.Y(n_1547)
);

INVx6_ASAP7_75t_L g1548 ( 
.A(n_1473),
.Y(n_1548)
);

INVx1_ASAP7_75t_L g1549 ( 
.A(n_1490),
.Y(n_1549)
);

BUFx3_ASAP7_75t_L g1550 ( 
.A(n_1350),
.Y(n_1550)
);

AOI22xp33_ASAP7_75t_L g1551 ( 
.A1(n_1424),
.A2(n_1386),
.B1(n_1485),
.B2(n_1418),
.Y(n_1551)
);

AOI22xp33_ASAP7_75t_SL g1552 ( 
.A1(n_1416),
.A2(n_1413),
.B1(n_1485),
.B2(n_1516),
.Y(n_1552)
);

BUFx12f_ASAP7_75t_L g1553 ( 
.A(n_1503),
.Y(n_1553)
);

CKINVDCx11_ASAP7_75t_R g1554 ( 
.A(n_1358),
.Y(n_1554)
);

CKINVDCx20_ASAP7_75t_R g1555 ( 
.A(n_1459),
.Y(n_1555)
);

INVx1_ASAP7_75t_L g1556 ( 
.A(n_1410),
.Y(n_1556)
);

INVx1_ASAP7_75t_L g1557 ( 
.A(n_1417),
.Y(n_1557)
);

CKINVDCx11_ASAP7_75t_R g1558 ( 
.A(n_1395),
.Y(n_1558)
);

AOI22xp33_ASAP7_75t_L g1559 ( 
.A1(n_1381),
.A2(n_1441),
.B1(n_1437),
.B2(n_1457),
.Y(n_1559)
);

NAND2x1p5_ASAP7_75t_L g1560 ( 
.A(n_1362),
.B(n_1450),
.Y(n_1560)
);

INVx5_ASAP7_75t_L g1561 ( 
.A(n_1450),
.Y(n_1561)
);

CKINVDCx6p67_ASAP7_75t_R g1562 ( 
.A(n_1455),
.Y(n_1562)
);

NAND2xp5_ASAP7_75t_L g1563 ( 
.A(n_1461),
.B(n_1374),
.Y(n_1563)
);

BUFx12f_ASAP7_75t_L g1564 ( 
.A(n_1432),
.Y(n_1564)
);

INVx1_ASAP7_75t_L g1565 ( 
.A(n_1440),
.Y(n_1565)
);

AOI21xp5_ASAP7_75t_SL g1566 ( 
.A1(n_1375),
.A2(n_1364),
.B(n_1368),
.Y(n_1566)
);

AOI22xp33_ASAP7_75t_L g1567 ( 
.A1(n_1382),
.A2(n_1365),
.B1(n_1413),
.B2(n_1489),
.Y(n_1567)
);

AOI22xp33_ASAP7_75t_L g1568 ( 
.A1(n_1382),
.A2(n_1501),
.B1(n_1378),
.B2(n_1351),
.Y(n_1568)
);

OAI22x1_ASAP7_75t_SL g1569 ( 
.A1(n_1486),
.A2(n_1434),
.B1(n_1388),
.B2(n_1458),
.Y(n_1569)
);

INVx1_ASAP7_75t_L g1570 ( 
.A(n_1440),
.Y(n_1570)
);

AOI22xp33_ASAP7_75t_L g1571 ( 
.A1(n_1414),
.A2(n_1369),
.B1(n_1443),
.B2(n_1442),
.Y(n_1571)
);

AOI22xp33_ASAP7_75t_L g1572 ( 
.A1(n_1369),
.A2(n_1443),
.B1(n_1442),
.B2(n_1451),
.Y(n_1572)
);

BUFx2_ASAP7_75t_SL g1573 ( 
.A(n_1458),
.Y(n_1573)
);

NAND2xp5_ASAP7_75t_L g1574 ( 
.A(n_1436),
.B(n_1448),
.Y(n_1574)
);

AND2x2_ASAP7_75t_L g1575 ( 
.A(n_1448),
.B(n_1472),
.Y(n_1575)
);

INVx1_ASAP7_75t_L g1576 ( 
.A(n_1470),
.Y(n_1576)
);

CKINVDCx11_ASAP7_75t_R g1577 ( 
.A(n_1432),
.Y(n_1577)
);

CKINVDCx6p67_ASAP7_75t_R g1578 ( 
.A(n_1432),
.Y(n_1578)
);

CKINVDCx14_ASAP7_75t_R g1579 ( 
.A(n_1466),
.Y(n_1579)
);

INVx1_ASAP7_75t_SL g1580 ( 
.A(n_1469),
.Y(n_1580)
);

BUFx10_ASAP7_75t_L g1581 ( 
.A(n_1466),
.Y(n_1581)
);

INVx1_ASAP7_75t_L g1582 ( 
.A(n_1470),
.Y(n_1582)
);

AOI22xp33_ASAP7_75t_L g1583 ( 
.A1(n_1348),
.A2(n_1406),
.B1(n_1383),
.B2(n_1429),
.Y(n_1583)
);

INVx1_ASAP7_75t_L g1584 ( 
.A(n_1399),
.Y(n_1584)
);

INVx1_ASAP7_75t_SL g1585 ( 
.A(n_1469),
.Y(n_1585)
);

INVx1_ASAP7_75t_L g1586 ( 
.A(n_1399),
.Y(n_1586)
);

INVx1_ASAP7_75t_L g1587 ( 
.A(n_1399),
.Y(n_1587)
);

INVx2_ASAP7_75t_SL g1588 ( 
.A(n_1466),
.Y(n_1588)
);

AOI22xp33_ASAP7_75t_L g1589 ( 
.A1(n_1425),
.A2(n_1429),
.B1(n_1392),
.B2(n_1465),
.Y(n_1589)
);

OAI22xp33_ASAP7_75t_L g1590 ( 
.A1(n_1465),
.A2(n_1456),
.B1(n_1462),
.B2(n_1464),
.Y(n_1590)
);

INVx1_ASAP7_75t_L g1591 ( 
.A(n_1456),
.Y(n_1591)
);

INVx1_ASAP7_75t_L g1592 ( 
.A(n_1462),
.Y(n_1592)
);

AOI22xp33_ASAP7_75t_L g1593 ( 
.A1(n_1425),
.A2(n_1354),
.B1(n_1409),
.B2(n_1372),
.Y(n_1593)
);

INVx8_ASAP7_75t_L g1594 ( 
.A(n_1515),
.Y(n_1594)
);

BUFx8_ASAP7_75t_L g1595 ( 
.A(n_1493),
.Y(n_1595)
);

INVx2_ASAP7_75t_L g1596 ( 
.A(n_1467),
.Y(n_1596)
);

OAI22xp5_ASAP7_75t_L g1597 ( 
.A1(n_1379),
.A2(n_1472),
.B1(n_1430),
.B2(n_1486),
.Y(n_1597)
);

CKINVDCx5p33_ASAP7_75t_R g1598 ( 
.A(n_1493),
.Y(n_1598)
);

AOI22xp33_ASAP7_75t_SL g1599 ( 
.A1(n_1421),
.A2(n_1402),
.B1(n_1460),
.B2(n_1468),
.Y(n_1599)
);

INVx2_ASAP7_75t_L g1600 ( 
.A(n_1394),
.Y(n_1600)
);

BUFx2_ASAP7_75t_L g1601 ( 
.A(n_1493),
.Y(n_1601)
);

AOI22xp33_ASAP7_75t_SL g1602 ( 
.A1(n_1400),
.A2(n_1484),
.B1(n_1367),
.B2(n_1471),
.Y(n_1602)
);

OAI22xp5_ASAP7_75t_L g1603 ( 
.A1(n_1367),
.A2(n_1484),
.B1(n_1463),
.B2(n_1499),
.Y(n_1603)
);

INVx2_ASAP7_75t_L g1604 ( 
.A(n_1394),
.Y(n_1604)
);

AOI22xp5_ASAP7_75t_L g1605 ( 
.A1(n_1439),
.A2(n_1423),
.B1(n_1419),
.B2(n_1499),
.Y(n_1605)
);

INVx1_ASAP7_75t_L g1606 ( 
.A(n_1412),
.Y(n_1606)
);

OAI22xp5_ASAP7_75t_L g1607 ( 
.A1(n_1499),
.A2(n_1515),
.B1(n_1393),
.B2(n_1427),
.Y(n_1607)
);

INVx3_ASAP7_75t_L g1608 ( 
.A(n_1515),
.Y(n_1608)
);

AOI22xp33_ASAP7_75t_L g1609 ( 
.A1(n_1372),
.A2(n_1427),
.B1(n_1389),
.B2(n_1366),
.Y(n_1609)
);

INVx5_ASAP7_75t_L g1610 ( 
.A(n_1356),
.Y(n_1610)
);

BUFx12f_ASAP7_75t_L g1611 ( 
.A(n_1420),
.Y(n_1611)
);

AND2x2_ASAP7_75t_L g1612 ( 
.A(n_1420),
.B(n_1415),
.Y(n_1612)
);

CKINVDCx11_ASAP7_75t_R g1613 ( 
.A(n_1420),
.Y(n_1613)
);

BUFx8_ASAP7_75t_L g1614 ( 
.A(n_1471),
.Y(n_1614)
);

AOI22xp33_ASAP7_75t_L g1615 ( 
.A1(n_1438),
.A2(n_1471),
.B1(n_1449),
.B2(n_1397),
.Y(n_1615)
);

AOI22xp33_ASAP7_75t_L g1616 ( 
.A1(n_1385),
.A2(n_1390),
.B1(n_1391),
.B2(n_1444),
.Y(n_1616)
);

INVx11_ASAP7_75t_L g1617 ( 
.A(n_1412),
.Y(n_1617)
);

INVx1_ASAP7_75t_L g1618 ( 
.A(n_1412),
.Y(n_1618)
);

AOI22xp33_ASAP7_75t_L g1619 ( 
.A1(n_1482),
.A2(n_1514),
.B1(n_1497),
.B2(n_1492),
.Y(n_1619)
);

AND2x4_ASAP7_75t_L g1620 ( 
.A(n_1394),
.B(n_1483),
.Y(n_1620)
);

BUFx3_ASAP7_75t_L g1621 ( 
.A(n_1405),
.Y(n_1621)
);

CKINVDCx5p33_ASAP7_75t_R g1622 ( 
.A(n_1415),
.Y(n_1622)
);

NAND2xp5_ASAP7_75t_L g1623 ( 
.A(n_1506),
.B(n_1415),
.Y(n_1623)
);

BUFx2_ASAP7_75t_R g1624 ( 
.A(n_1373),
.Y(n_1624)
);

OAI22xp5_ASAP7_75t_L g1625 ( 
.A1(n_1370),
.A2(n_1488),
.B1(n_1373),
.B2(n_1506),
.Y(n_1625)
);

BUFx6f_ASAP7_75t_L g1626 ( 
.A(n_1373),
.Y(n_1626)
);

INVx4_ASAP7_75t_L g1627 ( 
.A(n_1405),
.Y(n_1627)
);

CKINVDCx16_ASAP7_75t_R g1628 ( 
.A(n_1405),
.Y(n_1628)
);

INVx6_ASAP7_75t_L g1629 ( 
.A(n_1506),
.Y(n_1629)
);

CKINVDCx20_ASAP7_75t_R g1630 ( 
.A(n_1363),
.Y(n_1630)
);

CKINVDCx5p33_ASAP7_75t_R g1631 ( 
.A(n_1363),
.Y(n_1631)
);

INVx2_ASAP7_75t_L g1632 ( 
.A(n_1353),
.Y(n_1632)
);

AOI22xp5_ASAP7_75t_L g1633 ( 
.A1(n_1349),
.A2(n_904),
.B1(n_1118),
.B2(n_1082),
.Y(n_1633)
);

AOI22xp33_ASAP7_75t_SL g1634 ( 
.A1(n_1452),
.A2(n_904),
.B1(n_1118),
.B2(n_851),
.Y(n_1634)
);

INVx6_ASAP7_75t_L g1635 ( 
.A(n_1452),
.Y(n_1635)
);

INVx1_ASAP7_75t_SL g1636 ( 
.A(n_1452),
.Y(n_1636)
);

BUFx12f_ASAP7_75t_L g1637 ( 
.A(n_1396),
.Y(n_1637)
);

INVxp67_ASAP7_75t_L g1638 ( 
.A(n_1408),
.Y(n_1638)
);

BUFx2_ASAP7_75t_L g1639 ( 
.A(n_1513),
.Y(n_1639)
);

INVx6_ASAP7_75t_L g1640 ( 
.A(n_1473),
.Y(n_1640)
);

AOI22xp33_ASAP7_75t_L g1641 ( 
.A1(n_1508),
.A2(n_1502),
.B1(n_904),
.B2(n_1065),
.Y(n_1641)
);

AOI22xp33_ASAP7_75t_L g1642 ( 
.A1(n_1508),
.A2(n_1502),
.B1(n_904),
.B2(n_1065),
.Y(n_1642)
);

OAI22xp5_ASAP7_75t_L g1643 ( 
.A1(n_1508),
.A2(n_904),
.B1(n_964),
.B2(n_926),
.Y(n_1643)
);

AOI22xp33_ASAP7_75t_L g1644 ( 
.A1(n_1508),
.A2(n_1502),
.B1(n_904),
.B2(n_1065),
.Y(n_1644)
);

CKINVDCx6p67_ASAP7_75t_R g1645 ( 
.A(n_1473),
.Y(n_1645)
);

INVx1_ASAP7_75t_L g1646 ( 
.A(n_1476),
.Y(n_1646)
);

CKINVDCx20_ASAP7_75t_R g1647 ( 
.A(n_1380),
.Y(n_1647)
);

BUFx3_ASAP7_75t_L g1648 ( 
.A(n_1513),
.Y(n_1648)
);

OR2x2_ASAP7_75t_L g1649 ( 
.A(n_1480),
.B(n_1487),
.Y(n_1649)
);

BUFx4f_ASAP7_75t_SL g1650 ( 
.A(n_1347),
.Y(n_1650)
);

OAI21xp33_ASAP7_75t_SL g1651 ( 
.A1(n_1508),
.A2(n_904),
.B(n_1097),
.Y(n_1651)
);

CKINVDCx5p33_ASAP7_75t_R g1652 ( 
.A(n_1380),
.Y(n_1652)
);

BUFx12f_ASAP7_75t_L g1653 ( 
.A(n_1396),
.Y(n_1653)
);

AOI22xp33_ASAP7_75t_SL g1654 ( 
.A1(n_1357),
.A2(n_904),
.B1(n_1118),
.B2(n_851),
.Y(n_1654)
);

AOI22xp33_ASAP7_75t_L g1655 ( 
.A1(n_1508),
.A2(n_1502),
.B1(n_904),
.B2(n_1065),
.Y(n_1655)
);

OAI22xp5_ASAP7_75t_L g1656 ( 
.A1(n_1508),
.A2(n_904),
.B1(n_964),
.B2(n_926),
.Y(n_1656)
);

INVx2_ASAP7_75t_L g1657 ( 
.A(n_1476),
.Y(n_1657)
);

BUFx12f_ASAP7_75t_L g1658 ( 
.A(n_1396),
.Y(n_1658)
);

INVx1_ASAP7_75t_L g1659 ( 
.A(n_1476),
.Y(n_1659)
);

INVx1_ASAP7_75t_L g1660 ( 
.A(n_1476),
.Y(n_1660)
);

AOI22xp33_ASAP7_75t_L g1661 ( 
.A1(n_1508),
.A2(n_1502),
.B1(n_904),
.B2(n_1065),
.Y(n_1661)
);

BUFx2_ASAP7_75t_L g1662 ( 
.A(n_1513),
.Y(n_1662)
);

CKINVDCx20_ASAP7_75t_R g1663 ( 
.A(n_1380),
.Y(n_1663)
);

AOI22xp33_ASAP7_75t_L g1664 ( 
.A1(n_1508),
.A2(n_1502),
.B1(n_904),
.B2(n_1065),
.Y(n_1664)
);

AOI22xp33_ASAP7_75t_SL g1665 ( 
.A1(n_1357),
.A2(n_904),
.B1(n_1118),
.B2(n_851),
.Y(n_1665)
);

NAND2xp5_ASAP7_75t_L g1666 ( 
.A(n_1507),
.B(n_904),
.Y(n_1666)
);

INVx6_ASAP7_75t_L g1667 ( 
.A(n_1473),
.Y(n_1667)
);

INVx2_ASAP7_75t_L g1668 ( 
.A(n_1476),
.Y(n_1668)
);

INVx6_ASAP7_75t_L g1669 ( 
.A(n_1473),
.Y(n_1669)
);

CKINVDCx20_ASAP7_75t_R g1670 ( 
.A(n_1380),
.Y(n_1670)
);

INVx2_ASAP7_75t_L g1671 ( 
.A(n_1476),
.Y(n_1671)
);

AOI22xp33_ASAP7_75t_L g1672 ( 
.A1(n_1508),
.A2(n_1502),
.B1(n_904),
.B2(n_1065),
.Y(n_1672)
);

INVx1_ASAP7_75t_SL g1673 ( 
.A(n_1371),
.Y(n_1673)
);

AND2x2_ASAP7_75t_L g1674 ( 
.A(n_1507),
.B(n_1500),
.Y(n_1674)
);

AOI22xp33_ASAP7_75t_SL g1675 ( 
.A1(n_1357),
.A2(n_904),
.B1(n_1118),
.B2(n_851),
.Y(n_1675)
);

BUFx2_ASAP7_75t_L g1676 ( 
.A(n_1513),
.Y(n_1676)
);

HB1xp67_ASAP7_75t_L g1677 ( 
.A(n_1408),
.Y(n_1677)
);

AOI22xp33_ASAP7_75t_SL g1678 ( 
.A1(n_1357),
.A2(n_904),
.B1(n_1118),
.B2(n_851),
.Y(n_1678)
);

BUFx10_ASAP7_75t_L g1679 ( 
.A(n_1380),
.Y(n_1679)
);

INVx1_ASAP7_75t_L g1680 ( 
.A(n_1476),
.Y(n_1680)
);

NAND2xp5_ASAP7_75t_L g1681 ( 
.A(n_1507),
.B(n_904),
.Y(n_1681)
);

INVx1_ASAP7_75t_L g1682 ( 
.A(n_1476),
.Y(n_1682)
);

BUFx3_ASAP7_75t_L g1683 ( 
.A(n_1513),
.Y(n_1683)
);

BUFx8_ASAP7_75t_L g1684 ( 
.A(n_1371),
.Y(n_1684)
);

AOI22xp33_ASAP7_75t_SL g1685 ( 
.A1(n_1357),
.A2(n_904),
.B1(n_1118),
.B2(n_851),
.Y(n_1685)
);

INVx6_ASAP7_75t_L g1686 ( 
.A(n_1473),
.Y(n_1686)
);

INVx2_ASAP7_75t_L g1687 ( 
.A(n_1476),
.Y(n_1687)
);

INVx2_ASAP7_75t_L g1688 ( 
.A(n_1476),
.Y(n_1688)
);

AOI22xp33_ASAP7_75t_L g1689 ( 
.A1(n_1508),
.A2(n_1502),
.B1(n_904),
.B2(n_1065),
.Y(n_1689)
);

BUFx2_ASAP7_75t_L g1690 ( 
.A(n_1576),
.Y(n_1690)
);

INVx1_ASAP7_75t_L g1691 ( 
.A(n_1606),
.Y(n_1691)
);

INVx1_ASAP7_75t_L g1692 ( 
.A(n_1618),
.Y(n_1692)
);

AND2x2_ASAP7_75t_L g1693 ( 
.A(n_1612),
.B(n_1537),
.Y(n_1693)
);

AO21x1_ASAP7_75t_SL g1694 ( 
.A1(n_1584),
.A2(n_1587),
.B(n_1586),
.Y(n_1694)
);

OAI21x1_ASAP7_75t_L g1695 ( 
.A1(n_1547),
.A2(n_1619),
.B(n_1616),
.Y(n_1695)
);

BUFx3_ASAP7_75t_L g1696 ( 
.A(n_1536),
.Y(n_1696)
);

AND2x2_ASAP7_75t_L g1697 ( 
.A(n_1537),
.B(n_1631),
.Y(n_1697)
);

INVx2_ASAP7_75t_SL g1698 ( 
.A(n_1538),
.Y(n_1698)
);

NAND2xp5_ASAP7_75t_L g1699 ( 
.A(n_1666),
.B(n_1681),
.Y(n_1699)
);

INVx1_ASAP7_75t_L g1700 ( 
.A(n_1534),
.Y(n_1700)
);

INVx3_ASAP7_75t_L g1701 ( 
.A(n_1620),
.Y(n_1701)
);

BUFx6f_ASAP7_75t_L g1702 ( 
.A(n_1561),
.Y(n_1702)
);

NAND2xp5_ASAP7_75t_L g1703 ( 
.A(n_1649),
.B(n_1654),
.Y(n_1703)
);

INVx1_ASAP7_75t_L g1704 ( 
.A(n_1534),
.Y(n_1704)
);

HB1xp67_ASAP7_75t_L g1705 ( 
.A(n_1677),
.Y(n_1705)
);

AND2x2_ASAP7_75t_L g1706 ( 
.A(n_1628),
.B(n_1591),
.Y(n_1706)
);

INVx2_ASAP7_75t_L g1707 ( 
.A(n_1632),
.Y(n_1707)
);

INVx3_ASAP7_75t_L g1708 ( 
.A(n_1620),
.Y(n_1708)
);

HB1xp67_ASAP7_75t_L g1709 ( 
.A(n_1677),
.Y(n_1709)
);

CKINVDCx20_ASAP7_75t_R g1710 ( 
.A(n_1647),
.Y(n_1710)
);

OAI221xp5_ASAP7_75t_SL g1711 ( 
.A1(n_1641),
.A2(n_1689),
.B1(n_1644),
.B2(n_1655),
.C(n_1661),
.Y(n_1711)
);

INVx1_ASAP7_75t_L g1712 ( 
.A(n_1623),
.Y(n_1712)
);

INVx2_ASAP7_75t_L g1713 ( 
.A(n_1549),
.Y(n_1713)
);

HB1xp67_ASAP7_75t_L g1714 ( 
.A(n_1638),
.Y(n_1714)
);

INVx1_ASAP7_75t_L g1715 ( 
.A(n_1621),
.Y(n_1715)
);

INVx1_ASAP7_75t_L g1716 ( 
.A(n_1621),
.Y(n_1716)
);

INVx1_ASAP7_75t_L g1717 ( 
.A(n_1582),
.Y(n_1717)
);

NOR2xp67_ASAP7_75t_SL g1718 ( 
.A(n_1561),
.B(n_1566),
.Y(n_1718)
);

AOI21xp33_ASAP7_75t_L g1719 ( 
.A1(n_1643),
.A2(n_1656),
.B(n_1526),
.Y(n_1719)
);

BUFx2_ASAP7_75t_L g1720 ( 
.A(n_1614),
.Y(n_1720)
);

AND2x2_ASAP7_75t_L g1721 ( 
.A(n_1592),
.B(n_1634),
.Y(n_1721)
);

INVx4_ASAP7_75t_L g1722 ( 
.A(n_1561),
.Y(n_1722)
);

NAND2xp5_ASAP7_75t_SL g1723 ( 
.A(n_1665),
.B(n_1675),
.Y(n_1723)
);

INVx3_ASAP7_75t_L g1724 ( 
.A(n_1635),
.Y(n_1724)
);

INVx1_ASAP7_75t_L g1725 ( 
.A(n_1600),
.Y(n_1725)
);

INVx1_ASAP7_75t_L g1726 ( 
.A(n_1604),
.Y(n_1726)
);

BUFx2_ASAP7_75t_L g1727 ( 
.A(n_1614),
.Y(n_1727)
);

INVx1_ASAP7_75t_L g1728 ( 
.A(n_1627),
.Y(n_1728)
);

INVx1_ASAP7_75t_L g1729 ( 
.A(n_1622),
.Y(n_1729)
);

INVx2_ASAP7_75t_L g1730 ( 
.A(n_1556),
.Y(n_1730)
);

OAI21x1_ASAP7_75t_L g1731 ( 
.A1(n_1609),
.A2(n_1625),
.B(n_1615),
.Y(n_1731)
);

INVx2_ASAP7_75t_L g1732 ( 
.A(n_1557),
.Y(n_1732)
);

INVx1_ASAP7_75t_L g1733 ( 
.A(n_1626),
.Y(n_1733)
);

INVx3_ASAP7_75t_L g1734 ( 
.A(n_1635),
.Y(n_1734)
);

INVx1_ASAP7_75t_L g1735 ( 
.A(n_1626),
.Y(n_1735)
);

AND2x2_ASAP7_75t_L g1736 ( 
.A(n_1624),
.B(n_1626),
.Y(n_1736)
);

INVx1_ASAP7_75t_L g1737 ( 
.A(n_1626),
.Y(n_1737)
);

INVx1_ASAP7_75t_L g1738 ( 
.A(n_1629),
.Y(n_1738)
);

INVx2_ASAP7_75t_L g1739 ( 
.A(n_1520),
.Y(n_1739)
);

NAND2xp5_ASAP7_75t_L g1740 ( 
.A(n_1678),
.B(n_1685),
.Y(n_1740)
);

AND2x2_ASAP7_75t_L g1741 ( 
.A(n_1610),
.B(n_1630),
.Y(n_1741)
);

INVx2_ASAP7_75t_L g1742 ( 
.A(n_1646),
.Y(n_1742)
);

INVx2_ASAP7_75t_L g1743 ( 
.A(n_1659),
.Y(n_1743)
);

HB1xp67_ASAP7_75t_L g1744 ( 
.A(n_1638),
.Y(n_1744)
);

OAI21xp5_ASAP7_75t_L g1745 ( 
.A1(n_1651),
.A2(n_1642),
.B(n_1641),
.Y(n_1745)
);

INVx2_ASAP7_75t_L g1746 ( 
.A(n_1660),
.Y(n_1746)
);

INVxp67_ASAP7_75t_L g1747 ( 
.A(n_1533),
.Y(n_1747)
);

NOR2xp33_ASAP7_75t_L g1748 ( 
.A(n_1674),
.B(n_1521),
.Y(n_1748)
);

INVx2_ASAP7_75t_SL g1749 ( 
.A(n_1538),
.Y(n_1749)
);

BUFx6f_ASAP7_75t_L g1750 ( 
.A(n_1561),
.Y(n_1750)
);

INVx1_ASAP7_75t_L g1751 ( 
.A(n_1680),
.Y(n_1751)
);

INVx1_ASAP7_75t_L g1752 ( 
.A(n_1629),
.Y(n_1752)
);

INVx1_ASAP7_75t_L g1753 ( 
.A(n_1617),
.Y(n_1753)
);

INVx2_ASAP7_75t_L g1754 ( 
.A(n_1682),
.Y(n_1754)
);

INVx2_ASAP7_75t_L g1755 ( 
.A(n_1610),
.Y(n_1755)
);

OR2x6_ASAP7_75t_L g1756 ( 
.A(n_1611),
.B(n_1607),
.Y(n_1756)
);

OAI211xp5_ASAP7_75t_L g1757 ( 
.A1(n_1523),
.A2(n_1522),
.B(n_1672),
.C(n_1664),
.Y(n_1757)
);

CKINVDCx5p33_ASAP7_75t_R g1758 ( 
.A(n_1558),
.Y(n_1758)
);

INVxp67_ASAP7_75t_L g1759 ( 
.A(n_1517),
.Y(n_1759)
);

INVxp33_ASAP7_75t_L g1760 ( 
.A(n_1639),
.Y(n_1760)
);

INVx2_ASAP7_75t_L g1761 ( 
.A(n_1610),
.Y(n_1761)
);

INVx2_ASAP7_75t_L g1762 ( 
.A(n_1610),
.Y(n_1762)
);

OAI22xp5_ASAP7_75t_L g1763 ( 
.A1(n_1689),
.A2(n_1655),
.B1(n_1672),
.B2(n_1644),
.Y(n_1763)
);

OA21x2_ASAP7_75t_L g1764 ( 
.A1(n_1593),
.A2(n_1583),
.B(n_1567),
.Y(n_1764)
);

HB1xp67_ASAP7_75t_L g1765 ( 
.A(n_1580),
.Y(n_1765)
);

HB1xp67_ASAP7_75t_L g1766 ( 
.A(n_1585),
.Y(n_1766)
);

INVx1_ASAP7_75t_L g1767 ( 
.A(n_1636),
.Y(n_1767)
);

AO21x2_ASAP7_75t_L g1768 ( 
.A1(n_1530),
.A2(n_1542),
.B(n_1590),
.Y(n_1768)
);

INVx1_ASAP7_75t_L g1769 ( 
.A(n_1542),
.Y(n_1769)
);

OAI21x1_ASAP7_75t_L g1770 ( 
.A1(n_1568),
.A2(n_1589),
.B(n_1603),
.Y(n_1770)
);

BUFx3_ASAP7_75t_L g1771 ( 
.A(n_1536),
.Y(n_1771)
);

HB1xp67_ASAP7_75t_L g1772 ( 
.A(n_1575),
.Y(n_1772)
);

OR2x6_ASAP7_75t_L g1773 ( 
.A(n_1597),
.B(n_1529),
.Y(n_1773)
);

INVx2_ASAP7_75t_SL g1774 ( 
.A(n_1538),
.Y(n_1774)
);

INVx1_ASAP7_75t_L g1775 ( 
.A(n_1565),
.Y(n_1775)
);

INVx1_ASAP7_75t_L g1776 ( 
.A(n_1570),
.Y(n_1776)
);

INVx2_ASAP7_75t_SL g1777 ( 
.A(n_1548),
.Y(n_1777)
);

INVx1_ASAP7_75t_L g1778 ( 
.A(n_1530),
.Y(n_1778)
);

INVx2_ASAP7_75t_SL g1779 ( 
.A(n_1548),
.Y(n_1779)
);

CKINVDCx20_ASAP7_75t_R g1780 ( 
.A(n_1663),
.Y(n_1780)
);

OR2x2_ASAP7_75t_L g1781 ( 
.A(n_1539),
.B(n_1541),
.Y(n_1781)
);

INVx2_ASAP7_75t_SL g1782 ( 
.A(n_1548),
.Y(n_1782)
);

AND2x2_ASAP7_75t_L g1783 ( 
.A(n_1633),
.B(n_1546),
.Y(n_1783)
);

INVx1_ASAP7_75t_SL g1784 ( 
.A(n_1673),
.Y(n_1784)
);

INVx1_ASAP7_75t_L g1785 ( 
.A(n_1688),
.Y(n_1785)
);

OR2x2_ASAP7_75t_L g1786 ( 
.A(n_1539),
.B(n_1541),
.Y(n_1786)
);

AND2x2_ASAP7_75t_L g1787 ( 
.A(n_1546),
.B(n_1523),
.Y(n_1787)
);

CKINVDCx5p33_ASAP7_75t_R g1788 ( 
.A(n_1558),
.Y(n_1788)
);

INVx1_ASAP7_75t_L g1789 ( 
.A(n_1687),
.Y(n_1789)
);

INVx1_ASAP7_75t_L g1790 ( 
.A(n_1657),
.Y(n_1790)
);

INVx3_ASAP7_75t_L g1791 ( 
.A(n_1668),
.Y(n_1791)
);

INVx3_ASAP7_75t_L g1792 ( 
.A(n_1671),
.Y(n_1792)
);

AND2x2_ASAP7_75t_L g1793 ( 
.A(n_1522),
.B(n_1613),
.Y(n_1793)
);

INVxp67_ASAP7_75t_L g1794 ( 
.A(n_1662),
.Y(n_1794)
);

INVx1_ASAP7_75t_L g1795 ( 
.A(n_1613),
.Y(n_1795)
);

INVx1_ASAP7_75t_L g1796 ( 
.A(n_1568),
.Y(n_1796)
);

NAND2xp5_ASAP7_75t_L g1797 ( 
.A(n_1642),
.B(n_1661),
.Y(n_1797)
);

BUFx6f_ASAP7_75t_L g1798 ( 
.A(n_1519),
.Y(n_1798)
);

INVx1_ASAP7_75t_L g1799 ( 
.A(n_1590),
.Y(n_1799)
);

OAI21x1_ASAP7_75t_L g1800 ( 
.A1(n_1589),
.A2(n_1572),
.B(n_1593),
.Y(n_1800)
);

INVx3_ASAP7_75t_L g1801 ( 
.A(n_1528),
.Y(n_1801)
);

INVx3_ASAP7_75t_L g1802 ( 
.A(n_1528),
.Y(n_1802)
);

HB1xp67_ASAP7_75t_L g1803 ( 
.A(n_1550),
.Y(n_1803)
);

NAND2xp5_ASAP7_75t_L g1804 ( 
.A(n_1664),
.B(n_1525),
.Y(n_1804)
);

INVx1_ASAP7_75t_L g1805 ( 
.A(n_1572),
.Y(n_1805)
);

NAND2xp5_ASAP7_75t_L g1806 ( 
.A(n_1525),
.B(n_1524),
.Y(n_1806)
);

NAND2x1p5_ASAP7_75t_L g1807 ( 
.A(n_1527),
.B(n_1605),
.Y(n_1807)
);

INVx1_ASAP7_75t_L g1808 ( 
.A(n_1571),
.Y(n_1808)
);

AND2x4_ASAP7_75t_L g1809 ( 
.A(n_1531),
.B(n_1596),
.Y(n_1809)
);

OAI22xp5_ASAP7_75t_L g1810 ( 
.A1(n_1535),
.A2(n_1545),
.B1(n_1563),
.B2(n_1543),
.Y(n_1810)
);

INVx1_ASAP7_75t_L g1811 ( 
.A(n_1571),
.Y(n_1811)
);

INVx2_ASAP7_75t_SL g1812 ( 
.A(n_1640),
.Y(n_1812)
);

INVx1_ASAP7_75t_L g1813 ( 
.A(n_1552),
.Y(n_1813)
);

INVx1_ASAP7_75t_L g1814 ( 
.A(n_1559),
.Y(n_1814)
);

HB1xp67_ASAP7_75t_L g1815 ( 
.A(n_1550),
.Y(n_1815)
);

INVx1_ASAP7_75t_L g1816 ( 
.A(n_1559),
.Y(n_1816)
);

INVx1_ASAP7_75t_L g1817 ( 
.A(n_1599),
.Y(n_1817)
);

INVx1_ASAP7_75t_L g1818 ( 
.A(n_1551),
.Y(n_1818)
);

BUFx6f_ASAP7_75t_L g1819 ( 
.A(n_1519),
.Y(n_1819)
);

AOI22xp33_ASAP7_75t_L g1820 ( 
.A1(n_1524),
.A2(n_1551),
.B1(n_1602),
.B2(n_1684),
.Y(n_1820)
);

INVx1_ASAP7_75t_L g1821 ( 
.A(n_1532),
.Y(n_1821)
);

INVx1_ASAP7_75t_L g1822 ( 
.A(n_1532),
.Y(n_1822)
);

AND2x2_ASAP7_75t_L g1823 ( 
.A(n_1601),
.B(n_1608),
.Y(n_1823)
);

INVx1_ASAP7_75t_L g1824 ( 
.A(n_1560),
.Y(n_1824)
);

INVxp33_ASAP7_75t_L g1825 ( 
.A(n_1676),
.Y(n_1825)
);

INVx1_ASAP7_75t_L g1826 ( 
.A(n_1560),
.Y(n_1826)
);

INVx1_ASAP7_75t_L g1827 ( 
.A(n_1519),
.Y(n_1827)
);

NAND2xp5_ASAP7_75t_L g1828 ( 
.A(n_1574),
.B(n_1683),
.Y(n_1828)
);

INVx1_ASAP7_75t_L g1829 ( 
.A(n_1573),
.Y(n_1829)
);

AND2x2_ASAP7_75t_L g1830 ( 
.A(n_1579),
.B(n_1588),
.Y(n_1830)
);

INVxp33_ASAP7_75t_L g1831 ( 
.A(n_1648),
.Y(n_1831)
);

INVx1_ASAP7_75t_L g1832 ( 
.A(n_1581),
.Y(n_1832)
);

AOI22xp33_ASAP7_75t_L g1833 ( 
.A1(n_1684),
.A2(n_1553),
.B1(n_1683),
.B2(n_1648),
.Y(n_1833)
);

BUFx4f_ASAP7_75t_SL g1834 ( 
.A(n_1518),
.Y(n_1834)
);

INVx1_ASAP7_75t_L g1835 ( 
.A(n_1581),
.Y(n_1835)
);

INVx2_ASAP7_75t_L g1836 ( 
.A(n_1640),
.Y(n_1836)
);

NAND2xp5_ASAP7_75t_L g1837 ( 
.A(n_1700),
.B(n_1686),
.Y(n_1837)
);

OAI22xp5_ASAP7_75t_L g1838 ( 
.A1(n_1711),
.A2(n_1686),
.B1(n_1669),
.B2(n_1667),
.Y(n_1838)
);

O2A1O1Ixp33_ASAP7_75t_L g1839 ( 
.A1(n_1723),
.A2(n_1579),
.B(n_1544),
.C(n_1555),
.Y(n_1839)
);

AO32x1_ASAP7_75t_L g1840 ( 
.A1(n_1810),
.A2(n_1569),
.A3(n_1577),
.B1(n_1578),
.B2(n_1645),
.Y(n_1840)
);

AND2x4_ASAP7_75t_SL g1841 ( 
.A(n_1710),
.B(n_1679),
.Y(n_1841)
);

AND2x4_ASAP7_75t_SL g1842 ( 
.A(n_1780),
.B(n_1679),
.Y(n_1842)
);

OAI21xp5_ASAP7_75t_L g1843 ( 
.A1(n_1719),
.A2(n_1670),
.B(n_1544),
.Y(n_1843)
);

AOI22xp33_ASAP7_75t_L g1844 ( 
.A1(n_1787),
.A2(n_1540),
.B1(n_1650),
.B2(n_1667),
.Y(n_1844)
);

AND2x2_ASAP7_75t_L g1845 ( 
.A(n_1772),
.B(n_1598),
.Y(n_1845)
);

AND2x2_ASAP7_75t_L g1846 ( 
.A(n_1706),
.B(n_1577),
.Y(n_1846)
);

NOR2x1_ASAP7_75t_SL g1847 ( 
.A(n_1756),
.B(n_1564),
.Y(n_1847)
);

AND2x2_ASAP7_75t_L g1848 ( 
.A(n_1706),
.B(n_1652),
.Y(n_1848)
);

OAI21xp5_ASAP7_75t_L g1849 ( 
.A1(n_1757),
.A2(n_1640),
.B(n_1669),
.Y(n_1849)
);

NOR2xp33_ASAP7_75t_L g1850 ( 
.A(n_1787),
.B(n_1686),
.Y(n_1850)
);

CKINVDCx20_ASAP7_75t_R g1851 ( 
.A(n_1834),
.Y(n_1851)
);

AND2x2_ASAP7_75t_L g1852 ( 
.A(n_1741),
.B(n_1562),
.Y(n_1852)
);

AND2x2_ASAP7_75t_L g1853 ( 
.A(n_1795),
.B(n_1554),
.Y(n_1853)
);

AND2x4_ASAP7_75t_L g1854 ( 
.A(n_1753),
.B(n_1595),
.Y(n_1854)
);

NOR2xp33_ASAP7_75t_L g1855 ( 
.A(n_1740),
.B(n_1540),
.Y(n_1855)
);

AOI21xp5_ASAP7_75t_L g1856 ( 
.A1(n_1745),
.A2(n_1594),
.B(n_1595),
.Y(n_1856)
);

AO21x2_ASAP7_75t_L g1857 ( 
.A1(n_1695),
.A2(n_1594),
.B(n_1650),
.Y(n_1857)
);

AND2x2_ASAP7_75t_L g1858 ( 
.A(n_1795),
.B(n_1554),
.Y(n_1858)
);

INVxp67_ASAP7_75t_L g1859 ( 
.A(n_1705),
.Y(n_1859)
);

OA21x2_ASAP7_75t_L g1860 ( 
.A1(n_1731),
.A2(n_1637),
.B(n_1653),
.Y(n_1860)
);

AND2x2_ASAP7_75t_L g1861 ( 
.A(n_1697),
.B(n_1658),
.Y(n_1861)
);

AND2x2_ASAP7_75t_L g1862 ( 
.A(n_1697),
.B(n_1720),
.Y(n_1862)
);

AND2x2_ASAP7_75t_L g1863 ( 
.A(n_1720),
.B(n_1727),
.Y(n_1863)
);

A2O1A1Ixp33_ASAP7_75t_L g1864 ( 
.A1(n_1763),
.A2(n_1806),
.B(n_1783),
.C(n_1718),
.Y(n_1864)
);

OAI21xp33_ASAP7_75t_SL g1865 ( 
.A1(n_1820),
.A2(n_1793),
.B(n_1804),
.Y(n_1865)
);

OR2x2_ASAP7_75t_L g1866 ( 
.A(n_1729),
.B(n_1709),
.Y(n_1866)
);

NOR2x1_ASAP7_75t_R g1867 ( 
.A(n_1758),
.B(n_1788),
.Y(n_1867)
);

AND2x2_ASAP7_75t_L g1868 ( 
.A(n_1727),
.B(n_1693),
.Y(n_1868)
);

AOI21xp5_ASAP7_75t_L g1869 ( 
.A1(n_1770),
.A2(n_1764),
.B(n_1800),
.Y(n_1869)
);

AOI221xp5_ASAP7_75t_L g1870 ( 
.A1(n_1783),
.A2(n_1797),
.B1(n_1778),
.B2(n_1818),
.C(n_1793),
.Y(n_1870)
);

AND2x4_ASAP7_75t_L g1871 ( 
.A(n_1753),
.B(n_1809),
.Y(n_1871)
);

NOR2x1_ASAP7_75t_L g1872 ( 
.A(n_1696),
.B(n_1771),
.Y(n_1872)
);

A2O1A1Ixp33_ASAP7_75t_L g1873 ( 
.A1(n_1718),
.A2(n_1800),
.B(n_1781),
.C(n_1786),
.Y(n_1873)
);

AOI22xp5_ASAP7_75t_L g1874 ( 
.A1(n_1807),
.A2(n_1756),
.B1(n_1703),
.B2(n_1773),
.Y(n_1874)
);

AND2x4_ASAP7_75t_L g1875 ( 
.A(n_1809),
.B(n_1724),
.Y(n_1875)
);

AND2x4_ASAP7_75t_L g1876 ( 
.A(n_1809),
.B(n_1724),
.Y(n_1876)
);

O2A1O1Ixp33_ASAP7_75t_SL g1877 ( 
.A1(n_1781),
.A2(n_1786),
.B(n_1729),
.C(n_1818),
.Y(n_1877)
);

NAND2xp5_ASAP7_75t_L g1878 ( 
.A(n_1704),
.B(n_1778),
.Y(n_1878)
);

OR2x6_ASAP7_75t_L g1879 ( 
.A(n_1756),
.B(n_1773),
.Y(n_1879)
);

HB1xp67_ASAP7_75t_L g1880 ( 
.A(n_1690),
.Y(n_1880)
);

AND2x2_ASAP7_75t_L g1881 ( 
.A(n_1693),
.B(n_1736),
.Y(n_1881)
);

A2O1A1Ixp33_ASAP7_75t_L g1882 ( 
.A1(n_1813),
.A2(n_1799),
.B(n_1769),
.C(n_1808),
.Y(n_1882)
);

AND2x2_ASAP7_75t_L g1883 ( 
.A(n_1736),
.B(n_1803),
.Y(n_1883)
);

AO22x2_ASAP7_75t_L g1884 ( 
.A1(n_1715),
.A2(n_1716),
.B1(n_1799),
.B2(n_1817),
.Y(n_1884)
);

OR2x6_ASAP7_75t_L g1885 ( 
.A(n_1756),
.B(n_1773),
.Y(n_1885)
);

AOI22xp33_ASAP7_75t_L g1886 ( 
.A1(n_1768),
.A2(n_1807),
.B1(n_1699),
.B2(n_1811),
.Y(n_1886)
);

BUFx3_ASAP7_75t_L g1887 ( 
.A(n_1696),
.Y(n_1887)
);

AND2x2_ASAP7_75t_L g1888 ( 
.A(n_1815),
.B(n_1823),
.Y(n_1888)
);

BUFx2_ASAP7_75t_L g1889 ( 
.A(n_1771),
.Y(n_1889)
);

AOI22xp33_ASAP7_75t_L g1890 ( 
.A1(n_1807),
.A2(n_1808),
.B1(n_1811),
.B2(n_1813),
.Y(n_1890)
);

AO32x2_ASAP7_75t_L g1891 ( 
.A1(n_1698),
.A2(n_1779),
.A3(n_1812),
.B1(n_1777),
.B2(n_1749),
.Y(n_1891)
);

OAI21xp5_ASAP7_75t_L g1892 ( 
.A1(n_1769),
.A2(n_1796),
.B(n_1748),
.Y(n_1892)
);

AND2x2_ASAP7_75t_L g1893 ( 
.A(n_1823),
.B(n_1721),
.Y(n_1893)
);

AO32x2_ASAP7_75t_L g1894 ( 
.A1(n_1698),
.A2(n_1774),
.A3(n_1812),
.B1(n_1749),
.B2(n_1777),
.Y(n_1894)
);

OAI22xp5_ASAP7_75t_L g1895 ( 
.A1(n_1765),
.A2(n_1766),
.B1(n_1714),
.B2(n_1744),
.Y(n_1895)
);

A2O1A1Ixp33_ASAP7_75t_L g1896 ( 
.A1(n_1814),
.A2(n_1816),
.B(n_1805),
.C(n_1796),
.Y(n_1896)
);

HB1xp67_ASAP7_75t_L g1897 ( 
.A(n_1690),
.Y(n_1897)
);

NAND2xp5_ASAP7_75t_L g1898 ( 
.A(n_1704),
.B(n_1805),
.Y(n_1898)
);

BUFx2_ASAP7_75t_L g1899 ( 
.A(n_1827),
.Y(n_1899)
);

NOR2xp33_ASAP7_75t_L g1900 ( 
.A(n_1773),
.B(n_1747),
.Y(n_1900)
);

NOR2xp33_ASAP7_75t_L g1901 ( 
.A(n_1814),
.B(n_1816),
.Y(n_1901)
);

O2A1O1Ixp33_ASAP7_75t_L g1902 ( 
.A1(n_1759),
.A2(n_1794),
.B(n_1828),
.C(n_1784),
.Y(n_1902)
);

NAND2x1p5_ASAP7_75t_L g1903 ( 
.A(n_1702),
.B(n_1750),
.Y(n_1903)
);

OR2x2_ASAP7_75t_L g1904 ( 
.A(n_1713),
.B(n_1730),
.Y(n_1904)
);

AO21x2_ASAP7_75t_L g1905 ( 
.A1(n_1728),
.A2(n_1692),
.B(n_1691),
.Y(n_1905)
);

AND2x2_ASAP7_75t_L g1906 ( 
.A(n_1730),
.B(n_1732),
.Y(n_1906)
);

OAI21xp5_ASAP7_75t_L g1907 ( 
.A1(n_1760),
.A2(n_1825),
.B(n_1831),
.Y(n_1907)
);

NAND2xp5_ASAP7_75t_L g1908 ( 
.A(n_1775),
.B(n_1776),
.Y(n_1908)
);

AO32x2_ASAP7_75t_L g1909 ( 
.A1(n_1774),
.A2(n_1779),
.A3(n_1782),
.B1(n_1694),
.B2(n_1722),
.Y(n_1909)
);

AOI22xp33_ASAP7_75t_SL g1910 ( 
.A1(n_1764),
.A2(n_1758),
.B1(n_1788),
.B2(n_1702),
.Y(n_1910)
);

INVx1_ASAP7_75t_L g1911 ( 
.A(n_1717),
.Y(n_1911)
);

OR2x2_ASAP7_75t_L g1912 ( 
.A(n_1733),
.B(n_1735),
.Y(n_1912)
);

NOR2xp33_ASAP7_75t_L g1913 ( 
.A(n_1836),
.B(n_1829),
.Y(n_1913)
);

BUFx2_ASAP7_75t_R g1914 ( 
.A(n_1801),
.Y(n_1914)
);

AOI221xp5_ASAP7_75t_L g1915 ( 
.A1(n_1751),
.A2(n_1790),
.B1(n_1785),
.B2(n_1789),
.C(n_1775),
.Y(n_1915)
);

INVxp67_ASAP7_75t_SL g1916 ( 
.A(n_1691),
.Y(n_1916)
);

A2O1A1Ixp33_ASAP7_75t_SL g1917 ( 
.A1(n_1801),
.A2(n_1802),
.B(n_1826),
.C(n_1821),
.Y(n_1917)
);

NOR2x1_ASAP7_75t_SL g1918 ( 
.A(n_1694),
.B(n_1702),
.Y(n_1918)
);

INVx1_ASAP7_75t_L g1919 ( 
.A(n_1717),
.Y(n_1919)
);

AND2x2_ASAP7_75t_L g1920 ( 
.A(n_1739),
.B(n_1742),
.Y(n_1920)
);

A2O1A1Ixp33_ASAP7_75t_L g1921 ( 
.A1(n_1782),
.A2(n_1822),
.B(n_1826),
.C(n_1824),
.Y(n_1921)
);

AOI22xp33_ASAP7_75t_L g1922 ( 
.A1(n_1870),
.A2(n_1764),
.B1(n_1833),
.B2(n_1715),
.Y(n_1922)
);

OR2x2_ASAP7_75t_L g1923 ( 
.A(n_1880),
.B(n_1737),
.Y(n_1923)
);

OR2x6_ASAP7_75t_L g1924 ( 
.A(n_1879),
.B(n_1762),
.Y(n_1924)
);

INVx1_ASAP7_75t_L g1925 ( 
.A(n_1916),
.Y(n_1925)
);

HB1xp67_ASAP7_75t_L g1926 ( 
.A(n_1880),
.Y(n_1926)
);

BUFx6f_ASAP7_75t_L g1927 ( 
.A(n_1860),
.Y(n_1927)
);

INVx2_ASAP7_75t_L g1928 ( 
.A(n_1905),
.Y(n_1928)
);

INVx2_ASAP7_75t_SL g1929 ( 
.A(n_1897),
.Y(n_1929)
);

OR2x2_ASAP7_75t_L g1930 ( 
.A(n_1897),
.B(n_1859),
.Y(n_1930)
);

OR2x2_ASAP7_75t_L g1931 ( 
.A(n_1859),
.B(n_1767),
.Y(n_1931)
);

BUFx2_ASAP7_75t_SL g1932 ( 
.A(n_1854),
.Y(n_1932)
);

INVx1_ASAP7_75t_SL g1933 ( 
.A(n_1889),
.Y(n_1933)
);

INVx1_ASAP7_75t_L g1934 ( 
.A(n_1911),
.Y(n_1934)
);

AND2x2_ASAP7_75t_L g1935 ( 
.A(n_1869),
.B(n_1764),
.Y(n_1935)
);

INVx3_ASAP7_75t_L g1936 ( 
.A(n_1857),
.Y(n_1936)
);

NAND2xp5_ASAP7_75t_L g1937 ( 
.A(n_1878),
.B(n_1712),
.Y(n_1937)
);

AND2x2_ASAP7_75t_L g1938 ( 
.A(n_1884),
.B(n_1701),
.Y(n_1938)
);

INVx1_ASAP7_75t_L g1939 ( 
.A(n_1919),
.Y(n_1939)
);

AND2x4_ASAP7_75t_L g1940 ( 
.A(n_1857),
.B(n_1708),
.Y(n_1940)
);

HB1xp67_ASAP7_75t_L g1941 ( 
.A(n_1878),
.Y(n_1941)
);

AND2x2_ASAP7_75t_L g1942 ( 
.A(n_1884),
.B(n_1708),
.Y(n_1942)
);

NAND2xp5_ASAP7_75t_L g1943 ( 
.A(n_1901),
.B(n_1692),
.Y(n_1943)
);

AOI22xp33_ASAP7_75t_L g1944 ( 
.A1(n_1870),
.A2(n_1865),
.B1(n_1900),
.B2(n_1855),
.Y(n_1944)
);

OAI22xp5_ASAP7_75t_L g1945 ( 
.A1(n_1864),
.A2(n_1791),
.B1(n_1792),
.B2(n_1743),
.Y(n_1945)
);

AOI22xp33_ASAP7_75t_L g1946 ( 
.A1(n_1900),
.A2(n_1824),
.B1(n_1821),
.B2(n_1822),
.Y(n_1946)
);

BUFx2_ASAP7_75t_L g1947 ( 
.A(n_1909),
.Y(n_1947)
);

AND2x4_ASAP7_75t_L g1948 ( 
.A(n_1871),
.B(n_1875),
.Y(n_1948)
);

NAND2xp5_ASAP7_75t_SL g1949 ( 
.A(n_1874),
.B(n_1801),
.Y(n_1949)
);

AOI22xp33_ASAP7_75t_L g1950 ( 
.A1(n_1855),
.A2(n_1734),
.B1(n_1802),
.B2(n_1752),
.Y(n_1950)
);

AND2x2_ASAP7_75t_L g1951 ( 
.A(n_1909),
.B(n_1725),
.Y(n_1951)
);

NOR2x1_ASAP7_75t_L g1952 ( 
.A(n_1872),
.B(n_1746),
.Y(n_1952)
);

BUFx2_ASAP7_75t_R g1953 ( 
.A(n_1887),
.Y(n_1953)
);

AND2x2_ASAP7_75t_L g1954 ( 
.A(n_1909),
.B(n_1726),
.Y(n_1954)
);

BUFx3_ASAP7_75t_L g1955 ( 
.A(n_1903),
.Y(n_1955)
);

INVxp67_ASAP7_75t_L g1956 ( 
.A(n_1899),
.Y(n_1956)
);

NAND2xp5_ASAP7_75t_L g1957 ( 
.A(n_1901),
.B(n_1762),
.Y(n_1957)
);

NAND2xp5_ASAP7_75t_L g1958 ( 
.A(n_1898),
.B(n_1755),
.Y(n_1958)
);

AND2x2_ASAP7_75t_L g1959 ( 
.A(n_1881),
.B(n_1761),
.Y(n_1959)
);

OAI22xp5_ASAP7_75t_L g1960 ( 
.A1(n_1886),
.A2(n_1791),
.B1(n_1792),
.B2(n_1754),
.Y(n_1960)
);

OR2x2_ASAP7_75t_SL g1961 ( 
.A(n_1860),
.B(n_1754),
.Y(n_1961)
);

AOI22xp33_ASAP7_75t_L g1962 ( 
.A1(n_1892),
.A2(n_1802),
.B1(n_1752),
.B2(n_1738),
.Y(n_1962)
);

INVx2_ASAP7_75t_L g1963 ( 
.A(n_1906),
.Y(n_1963)
);

AND2x2_ASAP7_75t_L g1964 ( 
.A(n_1868),
.B(n_1761),
.Y(n_1964)
);

INVx2_ASAP7_75t_L g1965 ( 
.A(n_1904),
.Y(n_1965)
);

AND2x2_ASAP7_75t_L g1966 ( 
.A(n_1893),
.B(n_1707),
.Y(n_1966)
);

INVx1_ASAP7_75t_L g1967 ( 
.A(n_1908),
.Y(n_1967)
);

NOR3xp33_ASAP7_75t_SL g1968 ( 
.A(n_1949),
.B(n_1856),
.C(n_1945),
.Y(n_1968)
);

NAND2xp5_ASAP7_75t_L g1969 ( 
.A(n_1957),
.B(n_1895),
.Y(n_1969)
);

NAND2xp5_ASAP7_75t_L g1970 ( 
.A(n_1957),
.B(n_1895),
.Y(n_1970)
);

AND2x2_ASAP7_75t_L g1971 ( 
.A(n_1947),
.B(n_1888),
.Y(n_1971)
);

AO21x2_ASAP7_75t_L g1972 ( 
.A1(n_1928),
.A2(n_1917),
.B(n_1873),
.Y(n_1972)
);

AND2x4_ASAP7_75t_L g1973 ( 
.A(n_1940),
.B(n_1918),
.Y(n_1973)
);

INVx2_ASAP7_75t_L g1974 ( 
.A(n_1951),
.Y(n_1974)
);

INVxp67_ASAP7_75t_L g1975 ( 
.A(n_1930),
.Y(n_1975)
);

INVx4_ASAP7_75t_L g1976 ( 
.A(n_1927),
.Y(n_1976)
);

AND2x2_ASAP7_75t_L g1977 ( 
.A(n_1947),
.B(n_1862),
.Y(n_1977)
);

NAND2xp5_ASAP7_75t_L g1978 ( 
.A(n_1941),
.B(n_1920),
.Y(n_1978)
);

OR2x2_ASAP7_75t_L g1979 ( 
.A(n_1930),
.B(n_1866),
.Y(n_1979)
);

INVx1_ASAP7_75t_L g1980 ( 
.A(n_1925),
.Y(n_1980)
);

OR2x6_ASAP7_75t_L g1981 ( 
.A(n_1924),
.B(n_1879),
.Y(n_1981)
);

INVx2_ASAP7_75t_L g1982 ( 
.A(n_1951),
.Y(n_1982)
);

OAI22xp5_ASAP7_75t_L g1983 ( 
.A1(n_1944),
.A2(n_1886),
.B1(n_1890),
.B2(n_1910),
.Y(n_1983)
);

INVx2_ASAP7_75t_L g1984 ( 
.A(n_1951),
.Y(n_1984)
);

HB1xp67_ASAP7_75t_L g1985 ( 
.A(n_1926),
.Y(n_1985)
);

OAI221xp5_ASAP7_75t_L g1986 ( 
.A1(n_1946),
.A2(n_1839),
.B1(n_1843),
.B2(n_1844),
.C(n_1856),
.Y(n_1986)
);

OR2x2_ASAP7_75t_L g1987 ( 
.A(n_1929),
.B(n_1912),
.Y(n_1987)
);

OAI21xp5_ASAP7_75t_L g1988 ( 
.A1(n_1945),
.A2(n_1839),
.B(n_1910),
.Y(n_1988)
);

INVx2_ASAP7_75t_L g1989 ( 
.A(n_1954),
.Y(n_1989)
);

AO31x2_ASAP7_75t_L g1990 ( 
.A1(n_1928),
.A2(n_1921),
.A3(n_1882),
.B(n_1896),
.Y(n_1990)
);

INVx1_ASAP7_75t_L g1991 ( 
.A(n_1925),
.Y(n_1991)
);

AND2x2_ASAP7_75t_L g1992 ( 
.A(n_1964),
.B(n_1883),
.Y(n_1992)
);

NOR2x1p5_ASAP7_75t_L g1993 ( 
.A(n_1927),
.B(n_1854),
.Y(n_1993)
);

BUFx2_ASAP7_75t_L g1994 ( 
.A(n_1938),
.Y(n_1994)
);

NAND3xp33_ASAP7_75t_SL g1995 ( 
.A(n_1922),
.B(n_1902),
.C(n_1849),
.Y(n_1995)
);

NOR2x1_ASAP7_75t_SL g1996 ( 
.A(n_1924),
.B(n_1885),
.Y(n_1996)
);

INVx5_ASAP7_75t_L g1997 ( 
.A(n_1927),
.Y(n_1997)
);

INVx1_ASAP7_75t_SL g1998 ( 
.A(n_1933),
.Y(n_1998)
);

INVx2_ASAP7_75t_L g1999 ( 
.A(n_1954),
.Y(n_1999)
);

INVx1_ASAP7_75t_SL g2000 ( 
.A(n_1933),
.Y(n_2000)
);

AND2x2_ASAP7_75t_L g2001 ( 
.A(n_1964),
.B(n_1863),
.Y(n_2001)
);

INVx1_ASAP7_75t_SL g2002 ( 
.A(n_1926),
.Y(n_2002)
);

NAND2xp5_ASAP7_75t_L g2003 ( 
.A(n_1967),
.B(n_1902),
.Y(n_2003)
);

BUFx2_ASAP7_75t_SL g2004 ( 
.A(n_1929),
.Y(n_2004)
);

NOR2x1_ASAP7_75t_SL g2005 ( 
.A(n_1924),
.B(n_1885),
.Y(n_2005)
);

OAI31xp33_ASAP7_75t_L g2006 ( 
.A1(n_1960),
.A2(n_1838),
.A3(n_1877),
.B(n_1890),
.Y(n_2006)
);

INVx1_ASAP7_75t_L g2007 ( 
.A(n_1934),
.Y(n_2007)
);

INVx4_ASAP7_75t_L g2008 ( 
.A(n_1927),
.Y(n_2008)
);

INVx2_ASAP7_75t_SL g2009 ( 
.A(n_1929),
.Y(n_2009)
);

OAI22xp5_ASAP7_75t_L g2010 ( 
.A1(n_1953),
.A2(n_1914),
.B1(n_1844),
.B2(n_1885),
.Y(n_2010)
);

AND2x2_ASAP7_75t_L g2011 ( 
.A(n_1963),
.B(n_1891),
.Y(n_2011)
);

INVx1_ASAP7_75t_L g2012 ( 
.A(n_1934),
.Y(n_2012)
);

AOI22xp33_ASAP7_75t_L g2013 ( 
.A1(n_1932),
.A2(n_1850),
.B1(n_1861),
.B2(n_1876),
.Y(n_2013)
);

BUFx3_ASAP7_75t_L g2014 ( 
.A(n_1955),
.Y(n_2014)
);

AND2x2_ASAP7_75t_L g2015 ( 
.A(n_1959),
.B(n_1894),
.Y(n_2015)
);

AOI221xp5_ASAP7_75t_L g2016 ( 
.A1(n_1935),
.A2(n_1877),
.B1(n_1850),
.B2(n_1913),
.C(n_1837),
.Y(n_2016)
);

INVx2_ASAP7_75t_L g2017 ( 
.A(n_1954),
.Y(n_2017)
);

INVx1_ASAP7_75t_L g2018 ( 
.A(n_1939),
.Y(n_2018)
);

NAND3xp33_ASAP7_75t_L g2019 ( 
.A(n_1927),
.B(n_1915),
.C(n_1837),
.Y(n_2019)
);

INVx1_ASAP7_75t_L g2020 ( 
.A(n_1939),
.Y(n_2020)
);

OAI21xp5_ASAP7_75t_L g2021 ( 
.A1(n_1960),
.A2(n_1838),
.B(n_1913),
.Y(n_2021)
);

AND2x2_ASAP7_75t_L g2022 ( 
.A(n_1959),
.B(n_1894),
.Y(n_2022)
);

AND2x2_ASAP7_75t_L g2023 ( 
.A(n_1994),
.B(n_1948),
.Y(n_2023)
);

INVxp67_ASAP7_75t_L g2024 ( 
.A(n_2003),
.Y(n_2024)
);

OR2x2_ASAP7_75t_L g2025 ( 
.A(n_1994),
.B(n_1965),
.Y(n_2025)
);

OR2x2_ASAP7_75t_L g2026 ( 
.A(n_2002),
.B(n_1965),
.Y(n_2026)
);

HB1xp67_ASAP7_75t_L g2027 ( 
.A(n_1985),
.Y(n_2027)
);

INVx2_ASAP7_75t_L g2028 ( 
.A(n_1974),
.Y(n_2028)
);

NAND2xp5_ASAP7_75t_L g2029 ( 
.A(n_1969),
.B(n_1941),
.Y(n_2029)
);

AND2x2_ASAP7_75t_L g2030 ( 
.A(n_2015),
.B(n_1948),
.Y(n_2030)
);

AND2x2_ASAP7_75t_L g2031 ( 
.A(n_2015),
.B(n_1948),
.Y(n_2031)
);

INVx1_ASAP7_75t_L g2032 ( 
.A(n_2007),
.Y(n_2032)
);

INVx1_ASAP7_75t_L g2033 ( 
.A(n_2007),
.Y(n_2033)
);

NAND2xp5_ASAP7_75t_L g2034 ( 
.A(n_1970),
.B(n_1965),
.Y(n_2034)
);

NAND4xp25_ASAP7_75t_SL g2035 ( 
.A(n_2016),
.B(n_1846),
.C(n_1852),
.D(n_1858),
.Y(n_2035)
);

INVx2_ASAP7_75t_L g2036 ( 
.A(n_1974),
.Y(n_2036)
);

INVx1_ASAP7_75t_L g2037 ( 
.A(n_2012),
.Y(n_2037)
);

AND2x2_ASAP7_75t_L g2038 ( 
.A(n_2022),
.B(n_1948),
.Y(n_2038)
);

OAI33xp33_ASAP7_75t_L g2039 ( 
.A1(n_1983),
.A2(n_1943),
.A3(n_1931),
.B1(n_1967),
.B2(n_1937),
.B3(n_1958),
.Y(n_2039)
);

AND2x2_ASAP7_75t_L g2040 ( 
.A(n_2022),
.B(n_1948),
.Y(n_2040)
);

AND2x4_ASAP7_75t_SL g2041 ( 
.A(n_1968),
.B(n_1924),
.Y(n_2041)
);

INVx2_ASAP7_75t_L g2042 ( 
.A(n_1974),
.Y(n_2042)
);

OR2x2_ASAP7_75t_L g2043 ( 
.A(n_2002),
.B(n_1923),
.Y(n_2043)
);

INVx1_ASAP7_75t_L g2044 ( 
.A(n_2012),
.Y(n_2044)
);

NAND2xp5_ASAP7_75t_L g2045 ( 
.A(n_1998),
.B(n_1956),
.Y(n_2045)
);

NOR2x1_ASAP7_75t_L g2046 ( 
.A(n_1993),
.B(n_1952),
.Y(n_2046)
);

NAND2xp5_ASAP7_75t_L g2047 ( 
.A(n_1998),
.B(n_1956),
.Y(n_2047)
);

INVx1_ASAP7_75t_L g2048 ( 
.A(n_2018),
.Y(n_2048)
);

NAND2xp5_ASAP7_75t_L g2049 ( 
.A(n_2000),
.B(n_1943),
.Y(n_2049)
);

NAND2xp5_ASAP7_75t_L g2050 ( 
.A(n_2000),
.B(n_1966),
.Y(n_2050)
);

AND2x2_ASAP7_75t_L g2051 ( 
.A(n_1977),
.B(n_1924),
.Y(n_2051)
);

INVx1_ASAP7_75t_L g2052 ( 
.A(n_2018),
.Y(n_2052)
);

OR2x2_ASAP7_75t_L g2053 ( 
.A(n_1979),
.B(n_1923),
.Y(n_2053)
);

INVx1_ASAP7_75t_L g2054 ( 
.A(n_2020),
.Y(n_2054)
);

INVx1_ASAP7_75t_L g2055 ( 
.A(n_2020),
.Y(n_2055)
);

INVx1_ASAP7_75t_L g2056 ( 
.A(n_1980),
.Y(n_2056)
);

AND2x2_ASAP7_75t_L g2057 ( 
.A(n_1977),
.B(n_1924),
.Y(n_2057)
);

NAND2xp5_ASAP7_75t_L g2058 ( 
.A(n_1975),
.B(n_1966),
.Y(n_2058)
);

INVx2_ASAP7_75t_L g2059 ( 
.A(n_1982),
.Y(n_2059)
);

INVx1_ASAP7_75t_L g2060 ( 
.A(n_1980),
.Y(n_2060)
);

NOR2xp33_ASAP7_75t_SL g2061 ( 
.A(n_2006),
.B(n_1953),
.Y(n_2061)
);

INVx1_ASAP7_75t_SL g2062 ( 
.A(n_1979),
.Y(n_2062)
);

AND2x2_ASAP7_75t_L g2063 ( 
.A(n_1971),
.B(n_1938),
.Y(n_2063)
);

AND2x2_ASAP7_75t_L g2064 ( 
.A(n_1971),
.B(n_1973),
.Y(n_2064)
);

INVxp67_ASAP7_75t_L g2065 ( 
.A(n_1987),
.Y(n_2065)
);

NAND2xp5_ASAP7_75t_L g2066 ( 
.A(n_1978),
.B(n_1966),
.Y(n_2066)
);

INVx1_ASAP7_75t_L g2067 ( 
.A(n_1991),
.Y(n_2067)
);

AND2x2_ASAP7_75t_L g2068 ( 
.A(n_1973),
.B(n_1938),
.Y(n_2068)
);

AND2x4_ASAP7_75t_L g2069 ( 
.A(n_1993),
.B(n_1942),
.Y(n_2069)
);

NOR2x1_ASAP7_75t_SL g2070 ( 
.A(n_2004),
.B(n_1932),
.Y(n_2070)
);

OR2x2_ASAP7_75t_L g2071 ( 
.A(n_1987),
.B(n_1931),
.Y(n_2071)
);

AND2x2_ASAP7_75t_L g2072 ( 
.A(n_1973),
.B(n_1942),
.Y(n_2072)
);

AND2x2_ASAP7_75t_L g2073 ( 
.A(n_1973),
.B(n_1942),
.Y(n_2073)
);

AND2x4_ASAP7_75t_L g2074 ( 
.A(n_1996),
.B(n_1940),
.Y(n_2074)
);

NOR3xp33_ASAP7_75t_L g2075 ( 
.A(n_1995),
.B(n_1907),
.C(n_1936),
.Y(n_2075)
);

INVx2_ASAP7_75t_L g2076 ( 
.A(n_1982),
.Y(n_2076)
);

NAND2xp67_ASAP7_75t_L g2077 ( 
.A(n_2011),
.B(n_1841),
.Y(n_2077)
);

INVx1_ASAP7_75t_SL g2078 ( 
.A(n_2001),
.Y(n_2078)
);

OAI221xp5_ASAP7_75t_L g2079 ( 
.A1(n_1988),
.A2(n_1962),
.B1(n_1950),
.B2(n_1927),
.C(n_1853),
.Y(n_2079)
);

NAND2x1p5_ASAP7_75t_L g2080 ( 
.A(n_1997),
.B(n_1952),
.Y(n_2080)
);

AND2x2_ASAP7_75t_L g2081 ( 
.A(n_1996),
.B(n_2005),
.Y(n_2081)
);

INVx4_ASAP7_75t_L g2082 ( 
.A(n_1997),
.Y(n_2082)
);

INVx2_ASAP7_75t_SL g2083 ( 
.A(n_2023),
.Y(n_2083)
);

INVx1_ASAP7_75t_L g2084 ( 
.A(n_2032),
.Y(n_2084)
);

NAND2x1p5_ASAP7_75t_L g2085 ( 
.A(n_2046),
.B(n_1997),
.Y(n_2085)
);

INVx1_ASAP7_75t_L g2086 ( 
.A(n_2032),
.Y(n_2086)
);

INVx1_ASAP7_75t_L g2087 ( 
.A(n_2033),
.Y(n_2087)
);

INVx1_ASAP7_75t_L g2088 ( 
.A(n_2033),
.Y(n_2088)
);

NAND2xp5_ASAP7_75t_L g2089 ( 
.A(n_2024),
.B(n_2075),
.Y(n_2089)
);

INVx1_ASAP7_75t_L g2090 ( 
.A(n_2037),
.Y(n_2090)
);

INVx1_ASAP7_75t_L g2091 ( 
.A(n_2037),
.Y(n_2091)
);

INVx1_ASAP7_75t_L g2092 ( 
.A(n_2044),
.Y(n_2092)
);

INVx1_ASAP7_75t_L g2093 ( 
.A(n_2044),
.Y(n_2093)
);

NAND2xp5_ASAP7_75t_L g2094 ( 
.A(n_2029),
.B(n_1992),
.Y(n_2094)
);

INVx1_ASAP7_75t_SL g2095 ( 
.A(n_2045),
.Y(n_2095)
);

NAND2xp33_ASAP7_75t_L g2096 ( 
.A(n_2081),
.B(n_1988),
.Y(n_2096)
);

AND2x2_ASAP7_75t_L g2097 ( 
.A(n_2081),
.B(n_2005),
.Y(n_2097)
);

AND2x2_ASAP7_75t_L g2098 ( 
.A(n_2069),
.B(n_1982),
.Y(n_2098)
);

INVx2_ASAP7_75t_L g2099 ( 
.A(n_2028),
.Y(n_2099)
);

INVx2_ASAP7_75t_L g2100 ( 
.A(n_2028),
.Y(n_2100)
);

INVxp67_ASAP7_75t_L g2101 ( 
.A(n_2047),
.Y(n_2101)
);

NOR2xp67_ASAP7_75t_L g2102 ( 
.A(n_2082),
.B(n_1997),
.Y(n_2102)
);

INVx1_ASAP7_75t_L g2103 ( 
.A(n_2048),
.Y(n_2103)
);

OR2x2_ASAP7_75t_L g2104 ( 
.A(n_2053),
.B(n_2019),
.Y(n_2104)
);

NAND2xp5_ASAP7_75t_L g2105 ( 
.A(n_2062),
.B(n_2034),
.Y(n_2105)
);

INVx1_ASAP7_75t_L g2106 ( 
.A(n_2048),
.Y(n_2106)
);

INVx2_ASAP7_75t_L g2107 ( 
.A(n_2036),
.Y(n_2107)
);

NAND2xp5_ASAP7_75t_L g2108 ( 
.A(n_2049),
.B(n_1992),
.Y(n_2108)
);

NAND2x1p5_ASAP7_75t_L g2109 ( 
.A(n_2082),
.B(n_1997),
.Y(n_2109)
);

INVx2_ASAP7_75t_SL g2110 ( 
.A(n_2023),
.Y(n_2110)
);

INVx2_ASAP7_75t_L g2111 ( 
.A(n_2036),
.Y(n_2111)
);

AOI21xp33_ASAP7_75t_SL g2112 ( 
.A1(n_2079),
.A2(n_2010),
.B(n_1983),
.Y(n_2112)
);

OR2x2_ASAP7_75t_L g2113 ( 
.A(n_2053),
.B(n_2019),
.Y(n_2113)
);

AND2x2_ASAP7_75t_L g2114 ( 
.A(n_2069),
.B(n_1984),
.Y(n_2114)
);

INVx1_ASAP7_75t_L g2115 ( 
.A(n_2052),
.Y(n_2115)
);

AND2x2_ASAP7_75t_L g2116 ( 
.A(n_2069),
.B(n_1984),
.Y(n_2116)
);

OR2x2_ASAP7_75t_L g2117 ( 
.A(n_2071),
.B(n_1990),
.Y(n_2117)
);

INVx1_ASAP7_75t_L g2118 ( 
.A(n_2052),
.Y(n_2118)
);

INVx2_ASAP7_75t_L g2119 ( 
.A(n_2042),
.Y(n_2119)
);

INVx1_ASAP7_75t_L g2120 ( 
.A(n_2055),
.Y(n_2120)
);

HB1xp67_ASAP7_75t_L g2121 ( 
.A(n_2027),
.Y(n_2121)
);

OR2x2_ASAP7_75t_L g2122 ( 
.A(n_2071),
.B(n_1990),
.Y(n_2122)
);

AND2x2_ASAP7_75t_L g2123 ( 
.A(n_2064),
.B(n_1984),
.Y(n_2123)
);

NAND2x1_ASAP7_75t_L g2124 ( 
.A(n_2082),
.B(n_1976),
.Y(n_2124)
);

NAND2xp5_ASAP7_75t_L g2125 ( 
.A(n_2065),
.B(n_2001),
.Y(n_2125)
);

AOI321xp33_ASAP7_75t_L g2126 ( 
.A1(n_2035),
.A2(n_1986),
.A3(n_2010),
.B1(n_1935),
.B2(n_2013),
.C(n_2006),
.Y(n_2126)
);

INVx1_ASAP7_75t_L g2127 ( 
.A(n_2055),
.Y(n_2127)
);

INVx2_ASAP7_75t_L g2128 ( 
.A(n_2042),
.Y(n_2128)
);

AND2x2_ASAP7_75t_L g2129 ( 
.A(n_2064),
.B(n_1989),
.Y(n_2129)
);

INVx2_ASAP7_75t_L g2130 ( 
.A(n_2059),
.Y(n_2130)
);

INVx2_ASAP7_75t_L g2131 ( 
.A(n_2059),
.Y(n_2131)
);

INVx1_ASAP7_75t_L g2132 ( 
.A(n_2056),
.Y(n_2132)
);

AND2x2_ASAP7_75t_L g2133 ( 
.A(n_2051),
.B(n_1989),
.Y(n_2133)
);

AND2x2_ASAP7_75t_L g2134 ( 
.A(n_2051),
.B(n_1989),
.Y(n_2134)
);

INVx1_ASAP7_75t_L g2135 ( 
.A(n_2056),
.Y(n_2135)
);

AND2x2_ASAP7_75t_L g2136 ( 
.A(n_2057),
.B(n_1999),
.Y(n_2136)
);

INVx2_ASAP7_75t_L g2137 ( 
.A(n_2076),
.Y(n_2137)
);

INVx1_ASAP7_75t_L g2138 ( 
.A(n_2060),
.Y(n_2138)
);

NOR2xp33_ASAP7_75t_L g2139 ( 
.A(n_2077),
.B(n_1867),
.Y(n_2139)
);

INVx1_ASAP7_75t_L g2140 ( 
.A(n_2084),
.Y(n_2140)
);

NOR2xp33_ASAP7_75t_L g2141 ( 
.A(n_2112),
.B(n_2039),
.Y(n_2141)
);

OR2x2_ASAP7_75t_L g2142 ( 
.A(n_2095),
.B(n_2078),
.Y(n_2142)
);

OAI211xp5_ASAP7_75t_L g2143 ( 
.A1(n_2112),
.A2(n_2021),
.B(n_2061),
.C(n_1997),
.Y(n_2143)
);

NAND2xp5_ASAP7_75t_L g2144 ( 
.A(n_2089),
.B(n_2030),
.Y(n_2144)
);

NOR2xp33_ASAP7_75t_L g2145 ( 
.A(n_2139),
.B(n_2096),
.Y(n_2145)
);

NAND2xp5_ASAP7_75t_L g2146 ( 
.A(n_2101),
.B(n_2030),
.Y(n_2146)
);

OR2x2_ASAP7_75t_L g2147 ( 
.A(n_2105),
.B(n_2058),
.Y(n_2147)
);

AND2x2_ASAP7_75t_L g2148 ( 
.A(n_2097),
.B(n_2070),
.Y(n_2148)
);

NAND2xp5_ASAP7_75t_L g2149 ( 
.A(n_2121),
.B(n_2031),
.Y(n_2149)
);

OR2x2_ASAP7_75t_L g2150 ( 
.A(n_2104),
.B(n_2043),
.Y(n_2150)
);

NAND2xp5_ASAP7_75t_L g2151 ( 
.A(n_2104),
.B(n_2031),
.Y(n_2151)
);

AND2x4_ASAP7_75t_L g2152 ( 
.A(n_2102),
.B(n_2070),
.Y(n_2152)
);

NOR2xp33_ASAP7_75t_L g2153 ( 
.A(n_2113),
.B(n_2077),
.Y(n_2153)
);

AND2x2_ASAP7_75t_L g2154 ( 
.A(n_2097),
.B(n_2083),
.Y(n_2154)
);

INVx1_ASAP7_75t_L g2155 ( 
.A(n_2138),
.Y(n_2155)
);

NAND2xp5_ASAP7_75t_L g2156 ( 
.A(n_2113),
.B(n_2038),
.Y(n_2156)
);

AND2x2_ASAP7_75t_L g2157 ( 
.A(n_2083),
.B(n_2068),
.Y(n_2157)
);

NAND2x1_ASAP7_75t_L g2158 ( 
.A(n_2102),
.B(n_2074),
.Y(n_2158)
);

AND2x2_ASAP7_75t_L g2159 ( 
.A(n_2110),
.B(n_2068),
.Y(n_2159)
);

INVx1_ASAP7_75t_L g2160 ( 
.A(n_2084),
.Y(n_2160)
);

OR2x2_ASAP7_75t_L g2161 ( 
.A(n_2094),
.B(n_2043),
.Y(n_2161)
);

AND2x2_ASAP7_75t_L g2162 ( 
.A(n_2110),
.B(n_2072),
.Y(n_2162)
);

NAND2xp5_ASAP7_75t_L g2163 ( 
.A(n_2125),
.B(n_2038),
.Y(n_2163)
);

INVx1_ASAP7_75t_L g2164 ( 
.A(n_2086),
.Y(n_2164)
);

INVx1_ASAP7_75t_L g2165 ( 
.A(n_2086),
.Y(n_2165)
);

INVx1_ASAP7_75t_L g2166 ( 
.A(n_2138),
.Y(n_2166)
);

OR2x2_ASAP7_75t_L g2167 ( 
.A(n_2117),
.B(n_2025),
.Y(n_2167)
);

AND2x2_ASAP7_75t_L g2168 ( 
.A(n_2098),
.B(n_2072),
.Y(n_2168)
);

INVx1_ASAP7_75t_L g2169 ( 
.A(n_2087),
.Y(n_2169)
);

NOR3xp33_ASAP7_75t_L g2170 ( 
.A(n_2124),
.B(n_2008),
.C(n_1976),
.Y(n_2170)
);

INVx1_ASAP7_75t_L g2171 ( 
.A(n_2087),
.Y(n_2171)
);

NAND2xp5_ASAP7_75t_L g2172 ( 
.A(n_2108),
.B(n_2040),
.Y(n_2172)
);

AND2x2_ASAP7_75t_L g2173 ( 
.A(n_2098),
.B(n_2073),
.Y(n_2173)
);

INVx2_ASAP7_75t_SL g2174 ( 
.A(n_2124),
.Y(n_2174)
);

INVx1_ASAP7_75t_L g2175 ( 
.A(n_2088),
.Y(n_2175)
);

INVx1_ASAP7_75t_L g2176 ( 
.A(n_2088),
.Y(n_2176)
);

INVx1_ASAP7_75t_L g2177 ( 
.A(n_2090),
.Y(n_2177)
);

INVx1_ASAP7_75t_L g2178 ( 
.A(n_2090),
.Y(n_2178)
);

INVxp67_ASAP7_75t_SL g2179 ( 
.A(n_2085),
.Y(n_2179)
);

AND2x2_ASAP7_75t_L g2180 ( 
.A(n_2114),
.B(n_2116),
.Y(n_2180)
);

NOR4xp25_ASAP7_75t_L g2181 ( 
.A(n_2143),
.B(n_2126),
.C(n_2122),
.D(n_2117),
.Y(n_2181)
);

AOI221xp5_ASAP7_75t_L g2182 ( 
.A1(n_2141),
.A2(n_2021),
.B1(n_2126),
.B2(n_2122),
.C(n_2041),
.Y(n_2182)
);

INVx1_ASAP7_75t_SL g2183 ( 
.A(n_2174),
.Y(n_2183)
);

AND2x2_ASAP7_75t_L g2184 ( 
.A(n_2154),
.B(n_2073),
.Y(n_2184)
);

NAND2xp5_ASAP7_75t_L g2185 ( 
.A(n_2141),
.B(n_2091),
.Y(n_2185)
);

AND2x4_ASAP7_75t_L g2186 ( 
.A(n_2174),
.B(n_2114),
.Y(n_2186)
);

AOI32xp33_ASAP7_75t_L g2187 ( 
.A1(n_2153),
.A2(n_2041),
.A3(n_2116),
.B1(n_2074),
.B2(n_2134),
.Y(n_2187)
);

NAND3xp33_ASAP7_75t_SL g2188 ( 
.A(n_2153),
.B(n_2085),
.C(n_2109),
.Y(n_2188)
);

NAND2xp5_ASAP7_75t_L g2189 ( 
.A(n_2144),
.B(n_2133),
.Y(n_2189)
);

AOI211x1_ASAP7_75t_L g2190 ( 
.A1(n_2149),
.A2(n_2156),
.B(n_2151),
.C(n_2154),
.Y(n_2190)
);

OAI222xp33_ASAP7_75t_L g2191 ( 
.A1(n_2142),
.A2(n_2085),
.B1(n_2109),
.B2(n_1981),
.C1(n_2080),
.C2(n_2008),
.Y(n_2191)
);

INVx1_ASAP7_75t_L g2192 ( 
.A(n_2140),
.Y(n_2192)
);

AND2x2_ASAP7_75t_L g2193 ( 
.A(n_2180),
.B(n_2133),
.Y(n_2193)
);

OAI21xp33_ASAP7_75t_L g2194 ( 
.A1(n_2145),
.A2(n_2109),
.B(n_1935),
.Y(n_2194)
);

NOR2xp33_ASAP7_75t_L g2195 ( 
.A(n_2145),
.B(n_1851),
.Y(n_2195)
);

NOR2x1_ASAP7_75t_L g2196 ( 
.A(n_2152),
.B(n_2091),
.Y(n_2196)
);

OAI21xp33_ASAP7_75t_SL g2197 ( 
.A1(n_2179),
.A2(n_2136),
.B(n_2134),
.Y(n_2197)
);

INVx2_ASAP7_75t_L g2198 ( 
.A(n_2168),
.Y(n_2198)
);

INVx1_ASAP7_75t_L g2199 ( 
.A(n_2155),
.Y(n_2199)
);

NOR2xp33_ASAP7_75t_L g2200 ( 
.A(n_2146),
.B(n_1842),
.Y(n_2200)
);

INVx1_ASAP7_75t_L g2201 ( 
.A(n_2160),
.Y(n_2201)
);

AOI22xp5_ASAP7_75t_L g2202 ( 
.A1(n_2148),
.A2(n_2074),
.B1(n_1981),
.B2(n_1972),
.Y(n_2202)
);

NAND3xp33_ASAP7_75t_SL g2203 ( 
.A(n_2170),
.B(n_2080),
.C(n_2008),
.Y(n_2203)
);

XOR2x2_ASAP7_75t_L g2204 ( 
.A(n_2158),
.B(n_1847),
.Y(n_2204)
);

O2A1O1Ixp33_ASAP7_75t_L g2205 ( 
.A1(n_2150),
.A2(n_2080),
.B(n_2103),
.C(n_2135),
.Y(n_2205)
);

INVx1_ASAP7_75t_L g2206 ( 
.A(n_2164),
.Y(n_2206)
);

INVx1_ASAP7_75t_L g2207 ( 
.A(n_2165),
.Y(n_2207)
);

NAND2xp33_ASAP7_75t_L g2208 ( 
.A(n_2150),
.B(n_2148),
.Y(n_2208)
);

OAI22xp33_ASAP7_75t_SL g2209 ( 
.A1(n_2147),
.A2(n_1976),
.B1(n_2008),
.B2(n_2132),
.Y(n_2209)
);

OAI22xp5_ASAP7_75t_L g2210 ( 
.A1(n_2157),
.A2(n_1961),
.B1(n_1914),
.B2(n_2004),
.Y(n_2210)
);

INVx1_ASAP7_75t_L g2211 ( 
.A(n_2192),
.Y(n_2211)
);

INVx1_ASAP7_75t_L g2212 ( 
.A(n_2199),
.Y(n_2212)
);

INVx2_ASAP7_75t_SL g2213 ( 
.A(n_2186),
.Y(n_2213)
);

AOI221xp5_ASAP7_75t_L g2214 ( 
.A1(n_2181),
.A2(n_2175),
.B1(n_2178),
.B2(n_2177),
.C(n_2176),
.Y(n_2214)
);

NAND2xp5_ASAP7_75t_L g2215 ( 
.A(n_2185),
.B(n_2166),
.Y(n_2215)
);

NAND2xp5_ASAP7_75t_L g2216 ( 
.A(n_2190),
.B(n_2180),
.Y(n_2216)
);

OAI21xp5_ASAP7_75t_L g2217 ( 
.A1(n_2182),
.A2(n_2152),
.B(n_2169),
.Y(n_2217)
);

AOI22xp5_ASAP7_75t_L g2218 ( 
.A1(n_2208),
.A2(n_2152),
.B1(n_2157),
.B2(n_2159),
.Y(n_2218)
);

OAI22xp33_ASAP7_75t_SL g2219 ( 
.A1(n_2185),
.A2(n_2167),
.B1(n_2161),
.B2(n_2163),
.Y(n_2219)
);

INVxp67_ASAP7_75t_L g2220 ( 
.A(n_2195),
.Y(n_2220)
);

AND2x2_ASAP7_75t_L g2221 ( 
.A(n_2184),
.B(n_2159),
.Y(n_2221)
);

NAND2xp5_ASAP7_75t_L g2222 ( 
.A(n_2183),
.B(n_2168),
.Y(n_2222)
);

NOR4xp25_ASAP7_75t_SL g2223 ( 
.A(n_2194),
.B(n_2171),
.C(n_2106),
.D(n_2127),
.Y(n_2223)
);

INVx2_ASAP7_75t_L g2224 ( 
.A(n_2196),
.Y(n_2224)
);

NAND2xp5_ASAP7_75t_L g2225 ( 
.A(n_2183),
.B(n_2161),
.Y(n_2225)
);

A2O1A1Ixp33_ASAP7_75t_L g2226 ( 
.A1(n_2205),
.A2(n_2187),
.B(n_2188),
.C(n_2197),
.Y(n_2226)
);

INVx1_ASAP7_75t_L g2227 ( 
.A(n_2201),
.Y(n_2227)
);

AND2x4_ASAP7_75t_L g2228 ( 
.A(n_2186),
.B(n_2162),
.Y(n_2228)
);

A2O1A1Ixp33_ASAP7_75t_L g2229 ( 
.A1(n_2202),
.A2(n_2162),
.B(n_2173),
.C(n_2167),
.Y(n_2229)
);

OAI211xp5_ASAP7_75t_SL g2230 ( 
.A1(n_2206),
.A2(n_2207),
.B(n_2189),
.C(n_2198),
.Y(n_2230)
);

AOI22xp5_ASAP7_75t_L g2231 ( 
.A1(n_2210),
.A2(n_2173),
.B1(n_1972),
.B2(n_2172),
.Y(n_2231)
);

INVx2_ASAP7_75t_L g2232 ( 
.A(n_2193),
.Y(n_2232)
);

INVx1_ASAP7_75t_L g2233 ( 
.A(n_2209),
.Y(n_2233)
);

AND2x2_ASAP7_75t_L g2234 ( 
.A(n_2228),
.B(n_2200),
.Y(n_2234)
);

AND2x2_ASAP7_75t_L g2235 ( 
.A(n_2228),
.B(n_2221),
.Y(n_2235)
);

NAND2xp5_ASAP7_75t_SL g2236 ( 
.A(n_2219),
.B(n_2210),
.Y(n_2236)
);

INVx1_ASAP7_75t_L g2237 ( 
.A(n_2225),
.Y(n_2237)
);

NOR2xp33_ASAP7_75t_L g2238 ( 
.A(n_2220),
.B(n_2191),
.Y(n_2238)
);

NAND2xp5_ASAP7_75t_SL g2239 ( 
.A(n_2218),
.B(n_2204),
.Y(n_2239)
);

AOI211xp5_ASAP7_75t_L g2240 ( 
.A1(n_2217),
.A2(n_2203),
.B(n_1927),
.C(n_2106),
.Y(n_2240)
);

NAND3xp33_ASAP7_75t_L g2241 ( 
.A(n_2217),
.B(n_1976),
.C(n_2092),
.Y(n_2241)
);

O2A1O1Ixp33_ASAP7_75t_L g2242 ( 
.A1(n_2224),
.A2(n_2118),
.B(n_2092),
.C(n_2135),
.Y(n_2242)
);

XNOR2xp5_ASAP7_75t_L g2243 ( 
.A(n_2232),
.B(n_1848),
.Y(n_2243)
);

INVx1_ASAP7_75t_SL g2244 ( 
.A(n_2225),
.Y(n_2244)
);

OAI21xp5_ASAP7_75t_SL g2245 ( 
.A1(n_2226),
.A2(n_2136),
.B(n_2057),
.Y(n_2245)
);

OAI21xp33_ASAP7_75t_L g2246 ( 
.A1(n_2216),
.A2(n_2103),
.B(n_2093),
.Y(n_2246)
);

NAND3xp33_ASAP7_75t_L g2247 ( 
.A(n_2214),
.B(n_2115),
.C(n_2093),
.Y(n_2247)
);

NAND2xp5_ASAP7_75t_L g2248 ( 
.A(n_2213),
.B(n_2123),
.Y(n_2248)
);

INVx1_ASAP7_75t_L g2249 ( 
.A(n_2222),
.Y(n_2249)
);

NAND2xp5_ASAP7_75t_SL g2250 ( 
.A(n_2215),
.B(n_2115),
.Y(n_2250)
);

AOI211x1_ASAP7_75t_L g2251 ( 
.A1(n_2236),
.A2(n_2233),
.B(n_2215),
.C(n_2212),
.Y(n_2251)
);

INVx1_ASAP7_75t_L g2252 ( 
.A(n_2248),
.Y(n_2252)
);

HB1xp67_ASAP7_75t_L g2253 ( 
.A(n_2235),
.Y(n_2253)
);

INVx1_ASAP7_75t_SL g2254 ( 
.A(n_2244),
.Y(n_2254)
);

NOR3xp33_ASAP7_75t_L g2255 ( 
.A(n_2239),
.B(n_2230),
.C(n_2227),
.Y(n_2255)
);

NAND4xp25_ASAP7_75t_SL g2256 ( 
.A(n_2241),
.B(n_2229),
.C(n_2231),
.D(n_2211),
.Y(n_2256)
);

NAND2xp5_ASAP7_75t_SL g2257 ( 
.A(n_2240),
.B(n_2118),
.Y(n_2257)
);

OAI21xp33_ASAP7_75t_L g2258 ( 
.A1(n_2238),
.A2(n_2245),
.B(n_2249),
.Y(n_2258)
);

AND2x2_ASAP7_75t_L g2259 ( 
.A(n_2234),
.B(n_2223),
.Y(n_2259)
);

NAND2xp5_ASAP7_75t_SL g2260 ( 
.A(n_2238),
.B(n_2120),
.Y(n_2260)
);

NAND3x1_ASAP7_75t_L g2261 ( 
.A(n_2237),
.B(n_2127),
.C(n_2120),
.Y(n_2261)
);

AOI21xp33_ASAP7_75t_SL g2262 ( 
.A1(n_2243),
.A2(n_2132),
.B(n_1972),
.Y(n_2262)
);

NAND2xp5_ASAP7_75t_L g2263 ( 
.A(n_2246),
.B(n_2123),
.Y(n_2263)
);

O2A1O1Ixp33_ASAP7_75t_L g2264 ( 
.A1(n_2260),
.A2(n_2250),
.B(n_2247),
.C(n_2242),
.Y(n_2264)
);

AOI22xp5_ASAP7_75t_L g2265 ( 
.A1(n_2255),
.A2(n_2250),
.B1(n_1972),
.B2(n_2128),
.Y(n_2265)
);

INVx2_ASAP7_75t_L g2266 ( 
.A(n_2261),
.Y(n_2266)
);

OAI22xp5_ASAP7_75t_L g2267 ( 
.A1(n_2251),
.A2(n_2128),
.B1(n_2107),
.B2(n_2130),
.Y(n_2267)
);

NAND2xp5_ASAP7_75t_L g2268 ( 
.A(n_2253),
.B(n_2129),
.Y(n_2268)
);

AOI221x1_ASAP7_75t_L g2269 ( 
.A1(n_2258),
.A2(n_2137),
.B1(n_2131),
.B2(n_2100),
.C(n_2111),
.Y(n_2269)
);

O2A1O1Ixp33_ASAP7_75t_L g2270 ( 
.A1(n_2254),
.A2(n_2137),
.B(n_2131),
.C(n_2100),
.Y(n_2270)
);

AOI22xp5_ASAP7_75t_L g2271 ( 
.A1(n_2268),
.A2(n_2256),
.B1(n_2259),
.B2(n_2252),
.Y(n_2271)
);

NAND4xp25_ASAP7_75t_SL g2272 ( 
.A(n_2264),
.B(n_2265),
.C(n_2263),
.D(n_2262),
.Y(n_2272)
);

OAI21xp33_ASAP7_75t_L g2273 ( 
.A1(n_2266),
.A2(n_2263),
.B(n_2257),
.Y(n_2273)
);

OAI211xp5_ASAP7_75t_SL g2274 ( 
.A1(n_2270),
.A2(n_2137),
.B(n_2100),
.C(n_2131),
.Y(n_2274)
);

OAI211xp5_ASAP7_75t_SL g2275 ( 
.A1(n_2267),
.A2(n_2130),
.B(n_2119),
.C(n_2111),
.Y(n_2275)
);

NAND4xp75_ASAP7_75t_L g2276 ( 
.A(n_2269),
.B(n_2129),
.C(n_2119),
.D(n_2107),
.Y(n_2276)
);

INVx1_ASAP7_75t_L g2277 ( 
.A(n_2268),
.Y(n_2277)
);

NOR2xp33_ASAP7_75t_L g2278 ( 
.A(n_2273),
.B(n_2099),
.Y(n_2278)
);

AOI22xp5_ASAP7_75t_L g2279 ( 
.A1(n_2271),
.A2(n_2099),
.B1(n_2014),
.B2(n_2063),
.Y(n_2279)
);

AND2x4_ASAP7_75t_L g2280 ( 
.A(n_2277),
.B(n_2040),
.Y(n_2280)
);

NAND4xp75_ASAP7_75t_L g2281 ( 
.A(n_2272),
.B(n_1832),
.C(n_1835),
.D(n_1830),
.Y(n_2281)
);

AND3x4_ASAP7_75t_L g2282 ( 
.A(n_2276),
.B(n_2014),
.C(n_1955),
.Y(n_2282)
);

NAND4xp75_ASAP7_75t_L g2283 ( 
.A(n_2275),
.B(n_1835),
.C(n_2063),
.D(n_2009),
.Y(n_2283)
);

AOI221xp5_ASAP7_75t_L g2284 ( 
.A1(n_2278),
.A2(n_2274),
.B1(n_2060),
.B2(n_2067),
.C(n_2014),
.Y(n_2284)
);

AOI22xp5_ASAP7_75t_L g2285 ( 
.A1(n_2280),
.A2(n_1845),
.B1(n_1981),
.B2(n_2009),
.Y(n_2285)
);

AOI221xp5_ASAP7_75t_L g2286 ( 
.A1(n_2279),
.A2(n_2067),
.B1(n_2054),
.B2(n_1936),
.C(n_2050),
.Y(n_2286)
);

INVx2_ASAP7_75t_L g2287 ( 
.A(n_2285),
.Y(n_2287)
);

INVx1_ASAP7_75t_L g2288 ( 
.A(n_2287),
.Y(n_2288)
);

OAI22xp5_ASAP7_75t_L g2289 ( 
.A1(n_2288),
.A2(n_2282),
.B1(n_2281),
.B2(n_2283),
.Y(n_2289)
);

INVx1_ASAP7_75t_L g2290 ( 
.A(n_2288),
.Y(n_2290)
);

INVx1_ASAP7_75t_SL g2291 ( 
.A(n_2290),
.Y(n_2291)
);

HB1xp67_ASAP7_75t_L g2292 ( 
.A(n_2289),
.Y(n_2292)
);

OAI221xp5_ASAP7_75t_SL g2293 ( 
.A1(n_2291),
.A2(n_2284),
.B1(n_2286),
.B2(n_2026),
.C(n_2025),
.Y(n_2293)
);

AOI21xp5_ASAP7_75t_L g2294 ( 
.A1(n_2292),
.A2(n_1840),
.B(n_2066),
.Y(n_2294)
);

NAND2x1p5_ASAP7_75t_L g2295 ( 
.A(n_2294),
.B(n_1798),
.Y(n_2295)
);

XNOR2xp5_ASAP7_75t_L g2296 ( 
.A(n_2295),
.B(n_2293),
.Y(n_2296)
);

AOI22xp5_ASAP7_75t_L g2297 ( 
.A1(n_2296),
.A2(n_2076),
.B1(n_2026),
.B2(n_2017),
.Y(n_2297)
);

OAI221xp5_ASAP7_75t_R g2298 ( 
.A1(n_2297),
.A2(n_1840),
.B1(n_1961),
.B2(n_1917),
.C(n_1990),
.Y(n_2298)
);

AOI211xp5_ASAP7_75t_L g2299 ( 
.A1(n_2298),
.A2(n_1819),
.B(n_1798),
.C(n_1702),
.Y(n_2299)
);


endmodule