module fake_jpeg_18773_n_119 (n_13, n_21, n_33, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_19, n_18, n_20, n_35, n_4, n_34, n_30, n_16, n_3, n_0, n_24, n_28, n_38, n_26, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_12, n_32, n_8, n_15, n_7, n_119);

input n_13;
input n_21;
input n_33;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_35;
input n_4;
input n_34;
input n_30;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_119;

wire n_117;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_73;
wire n_84;
wire n_59;
wire n_98;
wire n_65;
wire n_110;
wire n_42;
wire n_49;
wire n_76;
wire n_88;
wire n_116;
wire n_114;
wire n_74;
wire n_103;
wire n_50;
wire n_57;
wire n_69;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_109;
wire n_113;
wire n_106;
wire n_111;
wire n_44;
wire n_75;
wire n_102;
wire n_99;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_56;
wire n_79;
wire n_67;
wire n_53;
wire n_54;
wire n_91;
wire n_93;
wire n_101;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_112;
wire n_95;
wire n_97;
wire n_62;
wire n_43;
wire n_100;
wire n_118;
wire n_82;
wire n_96;

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_34),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_25),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_8),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_17),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_29),
.Y(n_43)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_20),
.Y(n_44)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_24),
.Y(n_45)
);

INVx3_ASAP7_75t_L g46 ( 
.A(n_15),
.Y(n_46)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_36),
.Y(n_47)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_14),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g49 ( 
.A(n_13),
.B(n_6),
.Y(n_49)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_21),
.Y(n_50)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_30),
.Y(n_51)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_10),
.Y(n_52)
);

CKINVDCx5p33_ASAP7_75t_R g53 ( 
.A(n_6),
.Y(n_53)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_35),
.Y(n_54)
);

BUFx12f_ASAP7_75t_L g55 ( 
.A(n_19),
.Y(n_55)
);

BUFx24_ASAP7_75t_L g56 ( 
.A(n_53),
.Y(n_56)
);

INVx1_ASAP7_75t_SL g75 ( 
.A(n_56),
.Y(n_75)
);

INVx8_ASAP7_75t_L g57 ( 
.A(n_55),
.Y(n_57)
);

INVx5_ASAP7_75t_L g71 ( 
.A(n_57),
.Y(n_71)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_40),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g74 ( 
.A(n_58),
.Y(n_74)
);

INVx3_ASAP7_75t_L g59 ( 
.A(n_55),
.Y(n_59)
);

INVx2_ASAP7_75t_SL g67 ( 
.A(n_59),
.Y(n_67)
);

INVx8_ASAP7_75t_L g60 ( 
.A(n_55),
.Y(n_60)
);

INVx6_ASAP7_75t_L g65 ( 
.A(n_60),
.Y(n_65)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_40),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_61),
.B(n_62),
.Y(n_68)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_42),
.Y(n_62)
);

INVx8_ASAP7_75t_L g63 ( 
.A(n_42),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_63),
.B(n_54),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_SL g64 ( 
.A(n_56),
.B(n_53),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_L g88 ( 
.A(n_64),
.B(n_72),
.Y(n_88)
);

AOI22xp5_ASAP7_75t_L g66 ( 
.A1(n_63),
.A2(n_46),
.B1(n_44),
.B2(n_45),
.Y(n_66)
);

OAI22xp5_ASAP7_75t_SL g78 ( 
.A1(n_66),
.A2(n_69),
.B1(n_70),
.B2(n_75),
.Y(n_78)
);

AOI22xp33_ASAP7_75t_SL g69 ( 
.A1(n_58),
.A2(n_46),
.B1(n_52),
.B2(n_51),
.Y(n_69)
);

AOI22xp33_ASAP7_75t_SL g70 ( 
.A1(n_61),
.A2(n_48),
.B1(n_47),
.B2(n_43),
.Y(n_70)
);

CKINVDCx16_ASAP7_75t_R g72 ( 
.A(n_62),
.Y(n_72)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_73),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_SL g76 ( 
.A(n_56),
.B(n_41),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_L g90 ( 
.A(n_76),
.B(n_0),
.Y(n_90)
);

AOI22xp5_ASAP7_75t_L g92 ( 
.A1(n_78),
.A2(n_81),
.B1(n_82),
.B2(n_83),
.Y(n_92)
);

INVx4_ASAP7_75t_L g79 ( 
.A(n_65),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_79),
.B(n_80),
.Y(n_93)
);

BUFx3_ASAP7_75t_L g80 ( 
.A(n_74),
.Y(n_80)
);

AOI22xp33_ASAP7_75t_SL g81 ( 
.A1(n_65),
.A2(n_39),
.B1(n_50),
.B2(n_22),
.Y(n_81)
);

OAI22xp5_ASAP7_75t_L g82 ( 
.A1(n_69),
.A2(n_70),
.B1(n_68),
.B2(n_67),
.Y(n_82)
);

AOI22xp33_ASAP7_75t_SL g83 ( 
.A1(n_71),
.A2(n_16),
.B1(n_38),
.B2(n_37),
.Y(n_83)
);

AND2x2_ASAP7_75t_L g84 ( 
.A(n_75),
.B(n_49),
.Y(n_84)
);

MAJIxp5_ASAP7_75t_L g95 ( 
.A(n_84),
.B(n_1),
.C(n_2),
.Y(n_95)
);

BUFx2_ASAP7_75t_L g85 ( 
.A(n_74),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_85),
.B(n_89),
.Y(n_96)
);

OAI22xp5_ASAP7_75t_SL g86 ( 
.A1(n_67),
.A2(n_33),
.B1(n_11),
.B2(n_12),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_L g94 ( 
.A(n_86),
.B(n_1),
.Y(n_94)
);

HB1xp67_ASAP7_75t_L g87 ( 
.A(n_67),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_87),
.B(n_0),
.Y(n_91)
);

BUFx3_ASAP7_75t_L g89 ( 
.A(n_74),
.Y(n_89)
);

NAND3xp33_ASAP7_75t_L g101 ( 
.A(n_90),
.B(n_4),
.C(n_5),
.Y(n_101)
);

CKINVDCx16_ASAP7_75t_R g106 ( 
.A(n_91),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_SL g104 ( 
.A(n_94),
.B(n_95),
.Y(n_104)
);

MAJIxp5_ASAP7_75t_L g97 ( 
.A(n_88),
.B(n_18),
.C(n_31),
.Y(n_97)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_97),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_SL g98 ( 
.A(n_84),
.B(n_2),
.Y(n_98)
);

CKINVDCx20_ASAP7_75t_R g105 ( 
.A(n_98),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_77),
.B(n_3),
.Y(n_99)
);

AOI22xp5_ASAP7_75t_L g102 ( 
.A1(n_99),
.A2(n_100),
.B1(n_101),
.B2(n_4),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_87),
.B(n_3),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_102),
.B(n_91),
.Y(n_108)
);

OAI21xp5_ASAP7_75t_SL g107 ( 
.A1(n_106),
.A2(n_92),
.B(n_104),
.Y(n_107)
);

XOR2xp5_ASAP7_75t_L g110 ( 
.A(n_107),
.B(n_109),
.Y(n_110)
);

AND2x2_ASAP7_75t_L g111 ( 
.A(n_108),
.B(n_102),
.Y(n_111)
);

XOR2xp5_ASAP7_75t_L g109 ( 
.A(n_103),
.B(n_93),
.Y(n_109)
);

AOI22xp5_ASAP7_75t_L g112 ( 
.A1(n_111),
.A2(n_105),
.B1(n_103),
.B2(n_110),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_L g113 ( 
.A(n_112),
.B(n_96),
.Y(n_113)
);

MAJIxp5_ASAP7_75t_L g114 ( 
.A(n_113),
.B(n_83),
.C(n_81),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_L g115 ( 
.A(n_114),
.B(n_32),
.Y(n_115)
);

MAJIxp5_ASAP7_75t_L g116 ( 
.A(n_115),
.B(n_23),
.C(n_27),
.Y(n_116)
);

AOI21x1_ASAP7_75t_L g117 ( 
.A1(n_116),
.A2(n_7),
.B(n_9),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_L g118 ( 
.A(n_117),
.B(n_26),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_L g119 ( 
.A(n_118),
.B(n_28),
.Y(n_119)
);


endmodule