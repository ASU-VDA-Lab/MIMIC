module fake_netlist_1_12496_n_658 (n_44, n_81, n_69, n_22, n_57, n_52, n_26, n_50, n_33, n_73, n_49, n_80, n_60, n_41, n_35, n_65, n_9, n_10, n_19, n_74, n_7, n_29, n_45, n_62, n_36, n_47, n_37, n_34, n_5, n_23, n_8, n_16, n_13, n_70, n_17, n_63, n_14, n_71, n_56, n_42, n_24, n_78, n_6, n_4, n_40, n_79, n_38, n_64, n_46, n_31, n_58, n_32, n_0, n_84, n_55, n_12, n_75, n_72, n_43, n_76, n_68, n_27, n_53, n_67, n_77, n_20, n_2, n_54, n_83, n_28, n_48, n_11, n_25, n_30, n_59, n_3, n_18, n_66, n_1, n_82, n_15, n_61, n_21, n_51, n_39, n_658);
input n_44;
input n_81;
input n_69;
input n_22;
input n_57;
input n_52;
input n_26;
input n_50;
input n_33;
input n_73;
input n_49;
input n_80;
input n_60;
input n_41;
input n_35;
input n_65;
input n_9;
input n_10;
input n_19;
input n_74;
input n_7;
input n_29;
input n_45;
input n_62;
input n_36;
input n_47;
input n_37;
input n_34;
input n_5;
input n_23;
input n_8;
input n_16;
input n_13;
input n_70;
input n_17;
input n_63;
input n_14;
input n_71;
input n_56;
input n_42;
input n_24;
input n_78;
input n_6;
input n_4;
input n_40;
input n_79;
input n_38;
input n_64;
input n_46;
input n_31;
input n_58;
input n_32;
input n_0;
input n_84;
input n_55;
input n_12;
input n_75;
input n_72;
input n_43;
input n_76;
input n_68;
input n_27;
input n_53;
input n_67;
input n_77;
input n_20;
input n_2;
input n_54;
input n_83;
input n_28;
input n_48;
input n_11;
input n_25;
input n_30;
input n_59;
input n_3;
input n_18;
input n_66;
input n_1;
input n_82;
input n_15;
input n_61;
input n_21;
input n_51;
input n_39;
output n_658;
wire n_117;
wire n_361;
wire n_513;
wire n_185;
wire n_603;
wire n_604;
wire n_590;
wire n_407;
wire n_646;
wire n_284;
wire n_278;
wire n_500;
wire n_114;
wire n_607;
wire n_94;
wire n_125;
wire n_431;
wire n_484;
wire n_161;
wire n_496;
wire n_177;
wire n_130;
wire n_189;
wire n_311;
wire n_292;
wire n_309;
wire n_160;
wire n_612;
wire n_154;
wire n_328;
wire n_655;
wire n_468;
wire n_523;
wire n_229;
wire n_336;
wire n_464;
wire n_448;
wire n_645;
wire n_348;
wire n_252;
wire n_152;
wire n_113;
wire n_637;
wire n_353;
wire n_564;
wire n_528;
wire n_206;
wire n_288;
wire n_383;
wire n_532;
wire n_627;
wire n_544;
wire n_400;
wire n_296;
wire n_157;
wire n_202;
wire n_386;
wire n_432;
wire n_142;
wire n_232;
wire n_462;
wire n_316;
wire n_545;
wire n_211;
wire n_334;
wire n_389;
wire n_548;
wire n_436;
wire n_588;
wire n_275;
wire n_463;
wire n_131;
wire n_112;
wire n_205;
wire n_330;
wire n_587;
wire n_162;
wire n_387;
wire n_163;
wire n_476;
wire n_105;
wire n_227;
wire n_384;
wire n_434;
wire n_617;
wire n_231;
wire n_452;
wire n_518;
wire n_547;
wire n_298;
wire n_628;
wire n_411;
wire n_598;
wire n_144;
wire n_183;
wire n_489;
wire n_199;
wire n_351;
wire n_401;
wire n_100;
wire n_305;
wire n_461;
wire n_599;
wire n_228;
wire n_360;
wire n_345;
wire n_236;
wire n_340;
wire n_481;
wire n_443;
wire n_150;
wire n_373;
wire n_576;
wire n_301;
wire n_222;
wire n_234;
wire n_465;
wire n_609;
wire n_636;
wire n_366;
wire n_596;
wire n_286;
wire n_190;
wire n_246;
wire n_321;
wire n_572;
wire n_324;
wire n_392;
wire n_652;
wire n_279;
wire n_303;
wire n_437;
wire n_512;
wire n_326;
wire n_289;
wire n_333;
wire n_249;
wire n_642;
wire n_586;
wire n_244;
wire n_540;
wire n_563;
wire n_638;
wire n_141;
wire n_119;
wire n_517;
wire n_560;
wire n_479;
wire n_97;
wire n_167;
wire n_623;
wire n_593;
wire n_554;
wire n_447;
wire n_608;
wire n_171;
wire n_567;
wire n_196;
wire n_580;
wire n_192;
wire n_502;
wire n_543;
wire n_312;
wire n_455;
wire n_529;
wire n_630;
wire n_137;
wire n_511;
wire n_277;
wire n_467;
wire n_647;
wire n_367;
wire n_644;
wire n_85;
wire n_250;
wire n_314;
wire n_237;
wire n_181;
wire n_101;
wire n_255;
wire n_426;
wire n_624;
wire n_91;
wire n_108;
wire n_116;
wire n_230;
wire n_209;
wire n_274;
wire n_282;
wire n_319;
wire n_499;
wire n_417;
wire n_241;
wire n_575;
wire n_95;
wire n_238;
wire n_318;
wire n_471;
wire n_632;
wire n_293;
wire n_506;
wire n_533;
wire n_135;
wire n_393;
wire n_247;
wire n_490;
wire n_613;
wire n_648;
wire n_381;
wire n_550;
wire n_304;
wire n_399;
wire n_571;
wire n_294;
wire n_459;
wire n_313;
wire n_210;
wire n_184;
wire n_322;
wire n_310;
wire n_191;
wire n_307;
wire n_634;
wire n_610;
wire n_474;
wire n_354;
wire n_402;
wire n_413;
wire n_391;
wire n_427;
wire n_460;
wire n_478;
wire n_243;
wire n_235;
wire n_415;
wire n_394;
wire n_482;
wire n_442;
wire n_331;
wire n_485;
wire n_352;
wire n_619;
wire n_268;
wire n_174;
wire n_501;
wire n_248;
wire n_299;
wire n_89;
wire n_338;
wire n_519;
wire n_256;
wire n_551;
wire n_404;
wire n_369;
wire n_509;
wire n_651;
wire n_172;
wire n_329;
wire n_251;
wire n_635;
wire n_525;
wire n_218;
wire n_507;
wire n_605;
wire n_611;
wire n_633;
wire n_271;
wire n_626;
wire n_302;
wire n_466;
wire n_270;
wire n_362;
wire n_153;
wire n_259;
wire n_308;
wire n_546;
wire n_93;
wire n_412;
wire n_140;
wire n_207;
wire n_565;
wire n_224;
wire n_96;
wire n_219;
wire n_475;
wire n_578;
wire n_133;
wire n_149;
wire n_542;
wire n_537;
wire n_214;
wire n_204;
wire n_430;
wire n_88;
wire n_450;
wire n_579;
wire n_107;
wire n_403;
wire n_557;
wire n_516;
wire n_254;
wire n_549;
wire n_622;
wire n_262;
wire n_556;
wire n_239;
wire n_439;
wire n_601;
wire n_87;
wire n_379;
wire n_641;
wire n_614;
wire n_527;
wire n_98;
wire n_526;
wire n_276;
wire n_649;
wire n_320;
wire n_285;
wire n_195;
wire n_165;
wire n_446;
wire n_423;
wire n_342;
wire n_420;
wire n_621;
wire n_370;
wire n_589;
wire n_643;
wire n_574;
wire n_217;
wire n_139;
wire n_388;
wire n_454;
wire n_193;
wire n_273;
wire n_505;
wire n_390;
wire n_120;
wire n_514;
wire n_486;
wire n_568;
wire n_245;
wire n_357;
wire n_90;
wire n_653;
wire n_260;
wire n_539;
wire n_197;
wire n_201;
wire n_591;
wire n_317;
wire n_416;
wire n_374;
wire n_111;
wire n_536;
wire n_265;
wire n_264;
wire n_522;
wire n_200;
wire n_208;
wire n_573;
wire n_126;
wire n_178;
wire n_616;
wire n_118;
wire n_365;
wire n_541;
wire n_179;
wire n_315;
wire n_363;
wire n_409;
wire n_86;
wire n_143;
wire n_295;
wire n_654;
wire n_263;
wire n_166;
wire n_495;
wire n_186;
wire n_364;
wire n_428;
wire n_566;
wire n_376;
wire n_639;
wire n_552;
wire n_344;
wire n_136;
wire n_503;
wire n_283;
wire n_520;
wire n_435;
wire n_216;
wire n_577;
wire n_147;
wire n_148;
wire n_615;
wire n_212;
wire n_472;
wire n_92;
wire n_419;
wire n_396;
wire n_168;
wire n_477;
wire n_508;
wire n_570;
wire n_445;
wire n_398;
wire n_656;
wire n_438;
wire n_134;
wire n_640;
wire n_429;
wire n_488;
wire n_233;
wire n_106;
wire n_440;
wire n_553;
wire n_173;
wire n_422;
wire n_327;
wire n_325;
wire n_349;
wire n_498;
wire n_597;
wire n_225;
wire n_535;
wire n_530;
wire n_220;
wire n_358;
wire n_267;
wire n_221;
wire n_456;
wire n_203;
wire n_102;
wire n_449;
wire n_115;
wire n_300;
wire n_158;
wire n_524;
wire n_121;
wire n_584;
wire n_497;
wire n_339;
wire n_657;
wire n_583;
wire n_620;
wire n_240;
wire n_378;
wire n_582;
wire n_359;
wire n_346;
wire n_103;
wire n_180;
wire n_441;
wire n_104;
wire n_561;
wire n_335;
wire n_272;
wire n_594;
wire n_534;
wire n_531;
wire n_146;
wire n_397;
wire n_306;
wire n_215;
wire n_242;
wire n_155;
wire n_602;
wire n_198;
wire n_169;
wire n_424;
wire n_629;
wire n_156;
wire n_124;
wire n_569;
wire n_297;
wire n_128;
wire n_129;
wire n_410;
wire n_188;
wire n_377;
wire n_510;
wire n_343;
wire n_127;
wire n_291;
wire n_170;
wire n_504;
wire n_458;
wire n_581;
wire n_418;
wire n_493;
wire n_555;
wire n_380;
wire n_618;
wire n_356;
wire n_281;
wire n_341;
wire n_470;
wire n_600;
wire n_122;
wire n_187;
wire n_375;
wire n_138;
wire n_451;
wire n_487;
wire n_371;
wire n_323;
wire n_473;
wire n_347;
wire n_558;
wire n_258;
wire n_253;
wire n_515;
wire n_266;
wire n_213;
wire n_538;
wire n_182;
wire n_492;
wire n_592;
wire n_368;
wire n_355;
wire n_226;
wire n_382;
wire n_159;
wire n_337;
wire n_444;
wire n_176;
wire n_521;
wire n_650;
wire n_625;
wire n_469;
wire n_585;
wire n_123;
wire n_457;
wire n_595;
wire n_223;
wire n_494;
wire n_559;
wire n_480;
wire n_372;
wire n_453;
wire n_631;
wire n_194;
wire n_287;
wire n_110;
wire n_261;
wire n_606;
wire n_425;
wire n_332;
wire n_414;
wire n_562;
wire n_350;
wire n_433;
wire n_164;
wire n_421;
wire n_175;
wire n_145;
wire n_483;
wire n_408;
wire n_290;
wire n_405;
wire n_280;
wire n_99;
wire n_132;
wire n_109;
wire n_395;
wire n_406;
wire n_491;
wire n_151;
wire n_385;
wire n_257;
wire n_269;
CKINVDCx20_ASAP7_75t_R g85 ( .A(n_37), .Y(n_85) );
INVx1_ASAP7_75t_SL g86 ( .A(n_73), .Y(n_86) );
CKINVDCx5p33_ASAP7_75t_R g87 ( .A(n_39), .Y(n_87) );
INVx1_ASAP7_75t_L g88 ( .A(n_58), .Y(n_88) );
INVx1_ASAP7_75t_L g89 ( .A(n_69), .Y(n_89) );
CKINVDCx5p33_ASAP7_75t_R g90 ( .A(n_40), .Y(n_90) );
INVx1_ASAP7_75t_L g91 ( .A(n_81), .Y(n_91) );
INVx1_ASAP7_75t_L g92 ( .A(n_1), .Y(n_92) );
NOR2xp67_ASAP7_75t_L g93 ( .A(n_29), .B(n_65), .Y(n_93) );
INVx2_ASAP7_75t_SL g94 ( .A(n_22), .Y(n_94) );
INVx2_ASAP7_75t_L g95 ( .A(n_77), .Y(n_95) );
INVx1_ASAP7_75t_L g96 ( .A(n_5), .Y(n_96) );
INVx1_ASAP7_75t_L g97 ( .A(n_76), .Y(n_97) );
BUFx2_ASAP7_75t_L g98 ( .A(n_17), .Y(n_98) );
BUFx6f_ASAP7_75t_L g99 ( .A(n_17), .Y(n_99) );
BUFx3_ASAP7_75t_L g100 ( .A(n_44), .Y(n_100) );
CKINVDCx5p33_ASAP7_75t_R g101 ( .A(n_57), .Y(n_101) );
CKINVDCx16_ASAP7_75t_R g102 ( .A(n_50), .Y(n_102) );
INVx1_ASAP7_75t_L g103 ( .A(n_51), .Y(n_103) );
INVx1_ASAP7_75t_L g104 ( .A(n_9), .Y(n_104) );
INVx2_ASAP7_75t_L g105 ( .A(n_36), .Y(n_105) );
BUFx6f_ASAP7_75t_L g106 ( .A(n_71), .Y(n_106) );
CKINVDCx20_ASAP7_75t_R g107 ( .A(n_14), .Y(n_107) );
INVx2_ASAP7_75t_L g108 ( .A(n_54), .Y(n_108) );
INVx1_ASAP7_75t_L g109 ( .A(n_83), .Y(n_109) );
CKINVDCx14_ASAP7_75t_R g110 ( .A(n_11), .Y(n_110) );
INVx1_ASAP7_75t_L g111 ( .A(n_84), .Y(n_111) );
CKINVDCx5p33_ASAP7_75t_R g112 ( .A(n_8), .Y(n_112) );
INVx1_ASAP7_75t_L g113 ( .A(n_48), .Y(n_113) );
BUFx10_ASAP7_75t_L g114 ( .A(n_63), .Y(n_114) );
CKINVDCx14_ASAP7_75t_R g115 ( .A(n_9), .Y(n_115) );
INVx1_ASAP7_75t_L g116 ( .A(n_5), .Y(n_116) );
CKINVDCx5p33_ASAP7_75t_R g117 ( .A(n_80), .Y(n_117) );
CKINVDCx20_ASAP7_75t_R g118 ( .A(n_78), .Y(n_118) );
INVx1_ASAP7_75t_L g119 ( .A(n_60), .Y(n_119) );
INVx1_ASAP7_75t_L g120 ( .A(n_75), .Y(n_120) );
INVx1_ASAP7_75t_L g121 ( .A(n_0), .Y(n_121) );
INVx1_ASAP7_75t_L g122 ( .A(n_41), .Y(n_122) );
CKINVDCx20_ASAP7_75t_R g123 ( .A(n_35), .Y(n_123) );
INVx2_ASAP7_75t_L g124 ( .A(n_106), .Y(n_124) );
BUFx6f_ASAP7_75t_L g125 ( .A(n_106), .Y(n_125) );
NAND2xp5_ASAP7_75t_L g126 ( .A(n_94), .B(n_0), .Y(n_126) );
OA21x2_ASAP7_75t_L g127 ( .A1(n_95), .A2(n_42), .B(n_82), .Y(n_127) );
INVx1_ASAP7_75t_L g128 ( .A(n_88), .Y(n_128) );
NOR2xp33_ASAP7_75t_SL g129 ( .A(n_102), .B(n_20), .Y(n_129) );
NAND2xp5_ASAP7_75t_L g130 ( .A(n_94), .B(n_1), .Y(n_130) );
AND2x2_ASAP7_75t_L g131 ( .A(n_98), .B(n_2), .Y(n_131) );
INVx2_ASAP7_75t_L g132 ( .A(n_106), .Y(n_132) );
AND2x4_ASAP7_75t_L g133 ( .A(n_100), .B(n_2), .Y(n_133) );
BUFx6f_ASAP7_75t_L g134 ( .A(n_106), .Y(n_134) );
INVx3_ASAP7_75t_L g135 ( .A(n_114), .Y(n_135) );
OA22x2_ASAP7_75t_SL g136 ( .A1(n_107), .A2(n_3), .B1(n_4), .B2(n_6), .Y(n_136) );
OAI22xp5_ASAP7_75t_L g137 ( .A1(n_110), .A2(n_3), .B1(n_4), .B2(n_6), .Y(n_137) );
INVx2_ASAP7_75t_L g138 ( .A(n_106), .Y(n_138) );
CKINVDCx5p33_ASAP7_75t_R g139 ( .A(n_85), .Y(n_139) );
INVx2_ASAP7_75t_L g140 ( .A(n_95), .Y(n_140) );
NAND2xp5_ASAP7_75t_L g141 ( .A(n_92), .B(n_7), .Y(n_141) );
AND2x6_ASAP7_75t_L g142 ( .A(n_100), .B(n_45), .Y(n_142) );
AND2x4_ASAP7_75t_L g143 ( .A(n_105), .B(n_7), .Y(n_143) );
AOI22xp33_ASAP7_75t_L g144 ( .A1(n_143), .A2(n_96), .B1(n_121), .B2(n_104), .Y(n_144) );
INVx1_ASAP7_75t_L g145 ( .A(n_140), .Y(n_145) );
INVx2_ASAP7_75t_L g146 ( .A(n_124), .Y(n_146) );
OR2x2_ASAP7_75t_L g147 ( .A(n_131), .B(n_112), .Y(n_147) );
OAI22xp5_ASAP7_75t_SL g148 ( .A1(n_139), .A2(n_107), .B1(n_85), .B2(n_123), .Y(n_148) );
INVx2_ASAP7_75t_L g149 ( .A(n_124), .Y(n_149) );
NAND2xp5_ASAP7_75t_L g150 ( .A(n_135), .B(n_115), .Y(n_150) );
NOR2xp33_ASAP7_75t_L g151 ( .A(n_135), .B(n_89), .Y(n_151) );
BUFx6f_ASAP7_75t_L g152 ( .A(n_125), .Y(n_152) );
INVx1_ASAP7_75t_L g153 ( .A(n_140), .Y(n_153) );
OR2x6_ASAP7_75t_L g154 ( .A(n_137), .B(n_116), .Y(n_154) );
INVx3_ASAP7_75t_L g155 ( .A(n_143), .Y(n_155) );
BUFx3_ASAP7_75t_L g156 ( .A(n_142), .Y(n_156) );
INVx2_ASAP7_75t_L g157 ( .A(n_124), .Y(n_157) );
NOR2xp33_ASAP7_75t_L g158 ( .A(n_135), .B(n_91), .Y(n_158) );
AOI22xp5_ASAP7_75t_L g159 ( .A1(n_131), .A2(n_118), .B1(n_123), .B2(n_112), .Y(n_159) );
OR2x6_ASAP7_75t_L g160 ( .A(n_137), .B(n_99), .Y(n_160) );
NOR2xp33_ASAP7_75t_SL g161 ( .A(n_129), .B(n_118), .Y(n_161) );
NAND2xp5_ASAP7_75t_L g162 ( .A(n_135), .B(n_87), .Y(n_162) );
BUFx6f_ASAP7_75t_L g163 ( .A(n_125), .Y(n_163) );
INVx1_ASAP7_75t_L g164 ( .A(n_140), .Y(n_164) );
BUFx3_ASAP7_75t_L g165 ( .A(n_142), .Y(n_165) );
BUFx3_ASAP7_75t_L g166 ( .A(n_142), .Y(n_166) );
INVx1_ASAP7_75t_L g167 ( .A(n_143), .Y(n_167) );
INVx3_ASAP7_75t_L g168 ( .A(n_143), .Y(n_168) );
INVx1_ASAP7_75t_L g169 ( .A(n_133), .Y(n_169) );
INVx1_ASAP7_75t_L g170 ( .A(n_133), .Y(n_170) );
INVx2_ASAP7_75t_L g171 ( .A(n_125), .Y(n_171) );
INVx2_ASAP7_75t_L g172 ( .A(n_132), .Y(n_172) );
NAND2xp33_ASAP7_75t_R g173 ( .A(n_127), .B(n_87), .Y(n_173) );
INVx5_ASAP7_75t_L g174 ( .A(n_142), .Y(n_174) );
NAND2xp5_ASAP7_75t_L g175 ( .A(n_128), .B(n_90), .Y(n_175) );
NAND2xp5_ASAP7_75t_L g176 ( .A(n_175), .B(n_162), .Y(n_176) );
INVx2_ASAP7_75t_L g177 ( .A(n_146), .Y(n_177) );
AND2x2_ASAP7_75t_L g178 ( .A(n_147), .B(n_133), .Y(n_178) );
AOI22xp33_ASAP7_75t_L g179 ( .A1(n_169), .A2(n_133), .B1(n_128), .B2(n_129), .Y(n_179) );
NAND2xp5_ASAP7_75t_L g180 ( .A(n_150), .B(n_126), .Y(n_180) );
INVx2_ASAP7_75t_L g181 ( .A(n_146), .Y(n_181) );
NAND2xp5_ASAP7_75t_L g182 ( .A(n_151), .B(n_126), .Y(n_182) );
A2O1A1Ixp33_ASAP7_75t_L g183 ( .A1(n_169), .A2(n_130), .B(n_141), .C(n_97), .Y(n_183) );
NAND2xp5_ASAP7_75t_SL g184 ( .A(n_174), .B(n_90), .Y(n_184) );
INVxp67_ASAP7_75t_L g185 ( .A(n_147), .Y(n_185) );
NOR2xp33_ASAP7_75t_L g186 ( .A(n_167), .B(n_130), .Y(n_186) );
NOR2xp33_ASAP7_75t_L g187 ( .A(n_167), .B(n_141), .Y(n_187) );
NOR2xp33_ASAP7_75t_L g188 ( .A(n_155), .B(n_101), .Y(n_188) );
BUFx6f_ASAP7_75t_SL g189 ( .A(n_160), .Y(n_189) );
INVx2_ASAP7_75t_L g190 ( .A(n_149), .Y(n_190) );
AND2x4_ASAP7_75t_L g191 ( .A(n_144), .B(n_99), .Y(n_191) );
NOR2xp33_ASAP7_75t_L g192 ( .A(n_155), .B(n_101), .Y(n_192) );
NAND2xp5_ASAP7_75t_L g193 ( .A(n_158), .B(n_117), .Y(n_193) );
OR2x6_ASAP7_75t_L g194 ( .A(n_160), .B(n_154), .Y(n_194) );
INVx1_ASAP7_75t_L g195 ( .A(n_145), .Y(n_195) );
NAND2xp5_ASAP7_75t_SL g196 ( .A(n_174), .B(n_117), .Y(n_196) );
INVx1_ASAP7_75t_L g197 ( .A(n_145), .Y(n_197) );
NOR2xp67_ASAP7_75t_L g198 ( .A(n_155), .B(n_21), .Y(n_198) );
AOI21xp5_ASAP7_75t_L g199 ( .A1(n_170), .A2(n_127), .B(n_105), .Y(n_199) );
NAND2xp5_ASAP7_75t_SL g200 ( .A(n_174), .B(n_114), .Y(n_200) );
INVx2_ASAP7_75t_L g201 ( .A(n_149), .Y(n_201) );
INVx5_ASAP7_75t_L g202 ( .A(n_174), .Y(n_202) );
AOI22xp33_ASAP7_75t_L g203 ( .A1(n_170), .A2(n_142), .B1(n_99), .B2(n_127), .Y(n_203) );
INVx2_ASAP7_75t_L g204 ( .A(n_157), .Y(n_204) );
NAND2xp5_ASAP7_75t_SL g205 ( .A(n_174), .B(n_114), .Y(n_205) );
CKINVDCx5p33_ASAP7_75t_R g206 ( .A(n_148), .Y(n_206) );
INVx2_ASAP7_75t_L g207 ( .A(n_157), .Y(n_207) );
BUFx6f_ASAP7_75t_L g208 ( .A(n_156), .Y(n_208) );
NAND2xp5_ASAP7_75t_SL g209 ( .A(n_174), .B(n_86), .Y(n_209) );
INVx1_ASAP7_75t_L g210 ( .A(n_153), .Y(n_210) );
INVx1_ASAP7_75t_L g211 ( .A(n_153), .Y(n_211) );
AOI22xp33_ASAP7_75t_L g212 ( .A1(n_160), .A2(n_142), .B1(n_99), .B2(n_127), .Y(n_212) );
BUFx3_ASAP7_75t_L g213 ( .A(n_156), .Y(n_213) );
NAND2xp5_ASAP7_75t_L g214 ( .A(n_155), .B(n_142), .Y(n_214) );
NAND2xp5_ASAP7_75t_L g215 ( .A(n_168), .B(n_142), .Y(n_215) );
AOI21xp5_ASAP7_75t_L g216 ( .A1(n_215), .A2(n_156), .B(n_166), .Y(n_216) );
OAI22xp5_ASAP7_75t_L g217 ( .A1(n_194), .A2(n_159), .B1(n_168), .B2(n_160), .Y(n_217) );
INVx1_ASAP7_75t_L g218 ( .A(n_195), .Y(n_218) );
NAND2xp5_ASAP7_75t_L g219 ( .A(n_178), .B(n_168), .Y(n_219) );
NAND2xp5_ASAP7_75t_L g220 ( .A(n_178), .B(n_168), .Y(n_220) );
AOI21xp5_ASAP7_75t_L g221 ( .A1(n_215), .A2(n_165), .B(n_166), .Y(n_221) );
INVx1_ASAP7_75t_L g222 ( .A(n_195), .Y(n_222) );
A2O1A1Ixp33_ASAP7_75t_SL g223 ( .A1(n_212), .A2(n_164), .B(n_138), .C(n_132), .Y(n_223) );
NAND2xp5_ASAP7_75t_L g224 ( .A(n_180), .B(n_161), .Y(n_224) );
AOI22xp5_ASAP7_75t_L g225 ( .A1(n_185), .A2(n_160), .B1(n_159), .B2(n_154), .Y(n_225) );
OR2x6_ASAP7_75t_SL g226 ( .A(n_206), .B(n_148), .Y(n_226) );
AOI21xp5_ASAP7_75t_L g227 ( .A1(n_214), .A2(n_165), .B(n_166), .Y(n_227) );
OAI21xp33_ASAP7_75t_SL g228 ( .A1(n_194), .A2(n_154), .B(n_164), .Y(n_228) );
OAI22xp5_ASAP7_75t_L g229 ( .A1(n_194), .A2(n_154), .B1(n_165), .B2(n_173), .Y(n_229) );
INVx1_ASAP7_75t_L g230 ( .A(n_197), .Y(n_230) );
NOR2xp33_ASAP7_75t_L g231 ( .A(n_176), .B(n_154), .Y(n_231) );
AND2x2_ASAP7_75t_L g232 ( .A(n_194), .B(n_136), .Y(n_232) );
INVx5_ASAP7_75t_L g233 ( .A(n_194), .Y(n_233) );
NAND2x1p5_ASAP7_75t_L g234 ( .A(n_191), .B(n_127), .Y(n_234) );
O2A1O1Ixp33_ASAP7_75t_L g235 ( .A1(n_183), .A2(n_119), .B(n_103), .C(n_113), .Y(n_235) );
NAND2xp5_ASAP7_75t_L g236 ( .A(n_187), .B(n_142), .Y(n_236) );
NAND2xp5_ASAP7_75t_SL g237 ( .A(n_213), .B(n_109), .Y(n_237) );
AOI21xp5_ASAP7_75t_L g238 ( .A1(n_199), .A2(n_172), .B(n_171), .Y(n_238) );
O2A1O1Ixp5_ASAP7_75t_L g239 ( .A1(n_200), .A2(n_108), .B(n_111), .C(n_120), .Y(n_239) );
NAND2x1_ASAP7_75t_L g240 ( .A(n_197), .B(n_108), .Y(n_240) );
NAND2xp5_ASAP7_75t_SL g241 ( .A(n_213), .B(n_122), .Y(n_241) );
OR2x6_ASAP7_75t_L g242 ( .A(n_191), .B(n_136), .Y(n_242) );
O2A1O1Ixp5_ASAP7_75t_L g243 ( .A1(n_205), .A2(n_172), .B(n_171), .C(n_138), .Y(n_243) );
NAND2xp5_ASAP7_75t_L g244 ( .A(n_186), .B(n_8), .Y(n_244) );
INVx1_ASAP7_75t_L g245 ( .A(n_210), .Y(n_245) );
NAND2xp5_ASAP7_75t_SL g246 ( .A(n_213), .B(n_93), .Y(n_246) );
NOR2xp33_ASAP7_75t_L g247 ( .A(n_182), .B(n_10), .Y(n_247) );
AOI22xp5_ASAP7_75t_L g248 ( .A1(n_189), .A2(n_138), .B1(n_132), .B2(n_134), .Y(n_248) );
OAI21x1_ASAP7_75t_L g249 ( .A1(n_234), .A2(n_203), .B(n_198), .Y(n_249) );
OAI22xp5_ASAP7_75t_L g250 ( .A1(n_231), .A2(n_179), .B1(n_189), .B2(n_191), .Y(n_250) );
INVx1_ASAP7_75t_L g251 ( .A(n_218), .Y(n_251) );
NOR2x1_ASAP7_75t_L g252 ( .A(n_229), .B(n_191), .Y(n_252) );
AOI21x1_ASAP7_75t_L g253 ( .A1(n_238), .A2(n_198), .B(n_210), .Y(n_253) );
O2A1O1Ixp33_ASAP7_75t_SL g254 ( .A1(n_223), .A2(n_211), .B(n_209), .C(n_193), .Y(n_254) );
NAND2xp5_ASAP7_75t_SL g255 ( .A(n_233), .B(n_208), .Y(n_255) );
O2A1O1Ixp33_ASAP7_75t_SL g256 ( .A1(n_240), .A2(n_211), .B(n_184), .C(n_196), .Y(n_256) );
NAND2xp5_ASAP7_75t_L g257 ( .A(n_225), .B(n_188), .Y(n_257) );
INVx3_ASAP7_75t_L g258 ( .A(n_233), .Y(n_258) );
AO21x1_ASAP7_75t_L g259 ( .A1(n_234), .A2(n_192), .B(n_190), .Y(n_259) );
OAI21x1_ASAP7_75t_L g260 ( .A1(n_243), .A2(n_181), .B(n_207), .Y(n_260) );
INVx2_ASAP7_75t_L g261 ( .A(n_222), .Y(n_261) );
AOI22xp5_ASAP7_75t_L g262 ( .A1(n_217), .A2(n_189), .B1(n_206), .B2(n_207), .Y(n_262) );
NAND2xp5_ASAP7_75t_L g263 ( .A(n_224), .B(n_177), .Y(n_263) );
BUFx6f_ASAP7_75t_L g264 ( .A(n_233), .Y(n_264) );
AOI221xp5_ASAP7_75t_SL g265 ( .A1(n_235), .A2(n_177), .B1(n_204), .B2(n_201), .C(n_190), .Y(n_265) );
CKINVDCx11_ASAP7_75t_R g266 ( .A(n_226), .Y(n_266) );
OAI21x1_ASAP7_75t_L g267 ( .A1(n_227), .A2(n_204), .B(n_201), .Y(n_267) );
BUFx2_ASAP7_75t_L g268 ( .A(n_233), .Y(n_268) );
A2O1A1Ixp33_ASAP7_75t_L g269 ( .A1(n_228), .A2(n_181), .B(n_208), .C(n_125), .Y(n_269) );
OAI21x1_ASAP7_75t_L g270 ( .A1(n_216), .A2(n_221), .B(n_246), .Y(n_270) );
AOI221x1_ASAP7_75t_L g271 ( .A1(n_244), .A2(n_134), .B1(n_125), .B2(n_163), .C(n_152), .Y(n_271) );
BUFx8_ASAP7_75t_L g272 ( .A(n_264), .Y(n_272) );
OA21x2_ASAP7_75t_L g273 ( .A1(n_271), .A2(n_236), .B(n_230), .Y(n_273) );
AND2x2_ASAP7_75t_L g274 ( .A(n_261), .B(n_245), .Y(n_274) );
NAND2xp5_ASAP7_75t_L g275 ( .A(n_251), .B(n_219), .Y(n_275) );
AO222x2_ASAP7_75t_L g276 ( .A1(n_266), .A2(n_232), .B1(n_242), .B2(n_12), .C1(n_13), .C2(n_14), .Y(n_276) );
AND2x2_ASAP7_75t_L g277 ( .A(n_261), .B(n_242), .Y(n_277) );
INVx2_ASAP7_75t_SL g278 ( .A(n_264), .Y(n_278) );
HB1xp67_ASAP7_75t_L g279 ( .A(n_264), .Y(n_279) );
AO21x2_ASAP7_75t_L g280 ( .A1(n_269), .A2(n_247), .B(n_220), .Y(n_280) );
INVx1_ASAP7_75t_L g281 ( .A(n_251), .Y(n_281) );
AOI22xp33_ASAP7_75t_L g282 ( .A1(n_257), .A2(n_242), .B1(n_241), .B2(n_237), .Y(n_282) );
INVx1_ASAP7_75t_L g283 ( .A(n_263), .Y(n_283) );
AO31x2_ASAP7_75t_L g284 ( .A1(n_259), .A2(n_171), .A3(n_134), .B(n_125), .Y(n_284) );
INVx2_ASAP7_75t_L g285 ( .A(n_267), .Y(n_285) );
AOI21xp5_ASAP7_75t_L g286 ( .A1(n_259), .A2(n_239), .B(n_248), .Y(n_286) );
INVx1_ASAP7_75t_L g287 ( .A(n_264), .Y(n_287) );
OAI21xp5_ASAP7_75t_L g288 ( .A1(n_249), .A2(n_202), .B(n_208), .Y(n_288) );
AOI21xp5_ASAP7_75t_L g289 ( .A1(n_254), .A2(n_208), .B(n_163), .Y(n_289) );
AO21x2_ASAP7_75t_L g290 ( .A1(n_253), .A2(n_134), .B(n_11), .Y(n_290) );
INVx2_ASAP7_75t_SL g291 ( .A(n_264), .Y(n_291) );
INVx2_ASAP7_75t_L g292 ( .A(n_267), .Y(n_292) );
NAND2xp5_ASAP7_75t_SL g293 ( .A(n_252), .B(n_208), .Y(n_293) );
AOI21xp5_ASAP7_75t_L g294 ( .A1(n_271), .A2(n_163), .B(n_152), .Y(n_294) );
AOI221xp5_ASAP7_75t_L g295 ( .A1(n_276), .A2(n_250), .B1(n_262), .B2(n_265), .C(n_268), .Y(n_295) );
INVx2_ASAP7_75t_L g296 ( .A(n_292), .Y(n_296) );
AO21x2_ASAP7_75t_L g297 ( .A1(n_290), .A2(n_280), .B(n_286), .Y(n_297) );
HB1xp67_ASAP7_75t_L g298 ( .A(n_279), .Y(n_298) );
INVxp67_ASAP7_75t_SL g299 ( .A(n_292), .Y(n_299) );
INVx1_ASAP7_75t_L g300 ( .A(n_281), .Y(n_300) );
INVx2_ASAP7_75t_L g301 ( .A(n_292), .Y(n_301) );
INVx4_ASAP7_75t_L g302 ( .A(n_278), .Y(n_302) );
BUFx2_ASAP7_75t_L g303 ( .A(n_292), .Y(n_303) );
CKINVDCx5p33_ASAP7_75t_R g304 ( .A(n_272), .Y(n_304) );
INVx2_ASAP7_75t_L g305 ( .A(n_285), .Y(n_305) );
INVx1_ASAP7_75t_L g306 ( .A(n_281), .Y(n_306) );
INVx2_ASAP7_75t_L g307 ( .A(n_285), .Y(n_307) );
INVx1_ASAP7_75t_L g308 ( .A(n_285), .Y(n_308) );
OA21x2_ASAP7_75t_L g309 ( .A1(n_294), .A2(n_249), .B(n_270), .Y(n_309) );
AND2x2_ASAP7_75t_L g310 ( .A(n_277), .B(n_252), .Y(n_310) );
INVx2_ASAP7_75t_L g311 ( .A(n_284), .Y(n_311) );
INVx2_ASAP7_75t_L g312 ( .A(n_284), .Y(n_312) );
AO21x2_ASAP7_75t_L g313 ( .A1(n_290), .A2(n_253), .B(n_270), .Y(n_313) );
AND2x2_ASAP7_75t_L g314 ( .A(n_277), .B(n_268), .Y(n_314) );
INVx1_ASAP7_75t_L g315 ( .A(n_284), .Y(n_315) );
AND2x2_ASAP7_75t_L g316 ( .A(n_277), .B(n_258), .Y(n_316) );
BUFx3_ASAP7_75t_L g317 ( .A(n_272), .Y(n_317) );
INVx2_ASAP7_75t_L g318 ( .A(n_284), .Y(n_318) );
OAI21xp5_ASAP7_75t_L g319 ( .A1(n_286), .A2(n_260), .B(n_255), .Y(n_319) );
INVx1_ASAP7_75t_L g320 ( .A(n_284), .Y(n_320) );
OAI21x1_ASAP7_75t_L g321 ( .A1(n_294), .A2(n_260), .B(n_258), .Y(n_321) );
INVx1_ASAP7_75t_L g322 ( .A(n_274), .Y(n_322) );
OA21x2_ASAP7_75t_L g323 ( .A1(n_288), .A2(n_256), .B(n_134), .Y(n_323) );
BUFx6f_ASAP7_75t_L g324 ( .A(n_273), .Y(n_324) );
INVx1_ASAP7_75t_L g325 ( .A(n_284), .Y(n_325) );
AND2x4_ASAP7_75t_L g326 ( .A(n_278), .B(n_258), .Y(n_326) );
BUFx3_ASAP7_75t_L g327 ( .A(n_272), .Y(n_327) );
AND2x4_ASAP7_75t_L g328 ( .A(n_311), .B(n_284), .Y(n_328) );
NAND2xp5_ASAP7_75t_L g329 ( .A(n_322), .B(n_283), .Y(n_329) );
NAND2xp5_ASAP7_75t_SL g330 ( .A(n_304), .B(n_272), .Y(n_330) );
AND2x2_ASAP7_75t_L g331 ( .A(n_310), .B(n_274), .Y(n_331) );
AOI22xp33_ASAP7_75t_SL g332 ( .A1(n_317), .A2(n_276), .B1(n_272), .B2(n_290), .Y(n_332) );
AND2x2_ASAP7_75t_L g333 ( .A(n_310), .B(n_322), .Y(n_333) );
INVx2_ASAP7_75t_L g334 ( .A(n_296), .Y(n_334) );
AND2x2_ASAP7_75t_L g335 ( .A(n_310), .B(n_274), .Y(n_335) );
AND2x2_ASAP7_75t_L g336 ( .A(n_306), .B(n_284), .Y(n_336) );
AND2x2_ASAP7_75t_L g337 ( .A(n_306), .B(n_287), .Y(n_337) );
INVx4_ASAP7_75t_SL g338 ( .A(n_317), .Y(n_338) );
HB1xp67_ASAP7_75t_L g339 ( .A(n_303), .Y(n_339) );
INVx2_ASAP7_75t_L g340 ( .A(n_296), .Y(n_340) );
INVxp67_ASAP7_75t_SL g341 ( .A(n_299), .Y(n_341) );
AND2x2_ASAP7_75t_L g342 ( .A(n_300), .B(n_287), .Y(n_342) );
BUFx2_ASAP7_75t_L g343 ( .A(n_303), .Y(n_343) );
AND2x4_ASAP7_75t_SL g344 ( .A(n_302), .B(n_279), .Y(n_344) );
INVx2_ASAP7_75t_L g345 ( .A(n_296), .Y(n_345) );
BUFx2_ASAP7_75t_L g346 ( .A(n_303), .Y(n_346) );
INVx1_ASAP7_75t_L g347 ( .A(n_308), .Y(n_347) );
BUFx6f_ASAP7_75t_L g348 ( .A(n_324), .Y(n_348) );
AND2x2_ASAP7_75t_L g349 ( .A(n_315), .B(n_290), .Y(n_349) );
INVx1_ASAP7_75t_L g350 ( .A(n_296), .Y(n_350) );
AND2x2_ASAP7_75t_L g351 ( .A(n_315), .B(n_290), .Y(n_351) );
AND2x2_ASAP7_75t_L g352 ( .A(n_315), .B(n_280), .Y(n_352) );
NAND2xp5_ASAP7_75t_L g353 ( .A(n_316), .B(n_283), .Y(n_353) );
AND2x2_ASAP7_75t_L g354 ( .A(n_320), .B(n_280), .Y(n_354) );
NOR2x1_ASAP7_75t_L g355 ( .A(n_317), .B(n_293), .Y(n_355) );
INVx1_ASAP7_75t_L g356 ( .A(n_301), .Y(n_356) );
AND2x2_ASAP7_75t_L g357 ( .A(n_320), .B(n_280), .Y(n_357) );
INVx2_ASAP7_75t_L g358 ( .A(n_301), .Y(n_358) );
AND2x2_ASAP7_75t_L g359 ( .A(n_320), .B(n_280), .Y(n_359) );
INVx1_ASAP7_75t_L g360 ( .A(n_301), .Y(n_360) );
INVx2_ASAP7_75t_L g361 ( .A(n_301), .Y(n_361) );
NAND2xp5_ASAP7_75t_L g362 ( .A(n_316), .B(n_275), .Y(n_362) );
INVx4_ASAP7_75t_L g363 ( .A(n_317), .Y(n_363) );
INVx3_ASAP7_75t_L g364 ( .A(n_302), .Y(n_364) );
INVxp67_ASAP7_75t_L g365 ( .A(n_298), .Y(n_365) );
INVx2_ASAP7_75t_L g366 ( .A(n_305), .Y(n_366) );
INVx1_ASAP7_75t_L g367 ( .A(n_299), .Y(n_367) );
INVx2_ASAP7_75t_L g368 ( .A(n_305), .Y(n_368) );
AND2x2_ASAP7_75t_L g369 ( .A(n_314), .B(n_278), .Y(n_369) );
INVx2_ASAP7_75t_L g370 ( .A(n_305), .Y(n_370) );
OR2x2_ASAP7_75t_L g371 ( .A(n_298), .B(n_291), .Y(n_371) );
NAND2xp5_ASAP7_75t_L g372 ( .A(n_316), .B(n_275), .Y(n_372) );
INVx3_ASAP7_75t_L g373 ( .A(n_302), .Y(n_373) );
INVx1_ASAP7_75t_L g374 ( .A(n_325), .Y(n_374) );
AND2x2_ASAP7_75t_L g375 ( .A(n_314), .B(n_291), .Y(n_375) );
INVxp67_ASAP7_75t_SL g376 ( .A(n_305), .Y(n_376) );
AND2x2_ASAP7_75t_L g377 ( .A(n_314), .B(n_291), .Y(n_377) );
HB1xp67_ASAP7_75t_L g378 ( .A(n_307), .Y(n_378) );
OR2x2_ASAP7_75t_L g379 ( .A(n_325), .B(n_293), .Y(n_379) );
AND2x2_ASAP7_75t_L g380 ( .A(n_325), .B(n_288), .Y(n_380) );
AND2x2_ASAP7_75t_L g381 ( .A(n_311), .B(n_273), .Y(n_381) );
INVx2_ASAP7_75t_L g382 ( .A(n_378), .Y(n_382) );
CKINVDCx20_ASAP7_75t_R g383 ( .A(n_338), .Y(n_383) );
NAND2xp5_ASAP7_75t_L g384 ( .A(n_333), .B(n_295), .Y(n_384) );
NAND2xp5_ASAP7_75t_L g385 ( .A(n_331), .B(n_326), .Y(n_385) );
NAND2xp5_ASAP7_75t_L g386 ( .A(n_331), .B(n_326), .Y(n_386) );
AND2x4_ASAP7_75t_L g387 ( .A(n_364), .B(n_311), .Y(n_387) );
INVx2_ASAP7_75t_L g388 ( .A(n_378), .Y(n_388) );
AND2x2_ASAP7_75t_L g389 ( .A(n_335), .B(n_327), .Y(n_389) );
NAND2xp5_ASAP7_75t_L g390 ( .A(n_335), .B(n_326), .Y(n_390) );
AND2x2_ASAP7_75t_SL g391 ( .A(n_363), .B(n_302), .Y(n_391) );
AND2x4_ASAP7_75t_L g392 ( .A(n_364), .B(n_311), .Y(n_392) );
BUFx2_ASAP7_75t_L g393 ( .A(n_363), .Y(n_393) );
AND2x2_ASAP7_75t_L g394 ( .A(n_369), .B(n_327), .Y(n_394) );
AND2x2_ASAP7_75t_L g395 ( .A(n_369), .B(n_327), .Y(n_395) );
AND2x2_ASAP7_75t_L g396 ( .A(n_375), .B(n_327), .Y(n_396) );
NOR2xp33_ASAP7_75t_L g397 ( .A(n_332), .B(n_304), .Y(n_397) );
OR2x2_ASAP7_75t_L g398 ( .A(n_371), .B(n_307), .Y(n_398) );
AND2x2_ASAP7_75t_L g399 ( .A(n_375), .B(n_302), .Y(n_399) );
NAND2xp5_ASAP7_75t_L g400 ( .A(n_353), .B(n_326), .Y(n_400) );
AND2x4_ASAP7_75t_L g401 ( .A(n_364), .B(n_312), .Y(n_401) );
INVx1_ASAP7_75t_L g402 ( .A(n_342), .Y(n_402) );
NOR2xp33_ASAP7_75t_L g403 ( .A(n_332), .B(n_282), .Y(n_403) );
AND2x2_ASAP7_75t_L g404 ( .A(n_336), .B(n_312), .Y(n_404) );
OR2x2_ASAP7_75t_L g405 ( .A(n_362), .B(n_307), .Y(n_405) );
NAND2xp5_ASAP7_75t_L g406 ( .A(n_342), .B(n_326), .Y(n_406) );
INVx2_ASAP7_75t_L g407 ( .A(n_334), .Y(n_407) );
NAND2xp5_ASAP7_75t_L g408 ( .A(n_337), .B(n_312), .Y(n_408) );
OR2x2_ASAP7_75t_L g409 ( .A(n_362), .B(n_312), .Y(n_409) );
INVx2_ASAP7_75t_L g410 ( .A(n_334), .Y(n_410) );
HB1xp67_ASAP7_75t_L g411 ( .A(n_339), .Y(n_411) );
INVx1_ASAP7_75t_L g412 ( .A(n_337), .Y(n_412) );
AND2x2_ASAP7_75t_L g413 ( .A(n_377), .B(n_318), .Y(n_413) );
NAND2xp5_ASAP7_75t_L g414 ( .A(n_329), .B(n_318), .Y(n_414) );
HB1xp67_ASAP7_75t_L g415 ( .A(n_339), .Y(n_415) );
HB1xp67_ASAP7_75t_L g416 ( .A(n_341), .Y(n_416) );
NAND2xp5_ASAP7_75t_L g417 ( .A(n_329), .B(n_318), .Y(n_417) );
AND2x4_ASAP7_75t_L g418 ( .A(n_364), .B(n_297), .Y(n_418) );
INVx2_ASAP7_75t_L g419 ( .A(n_334), .Y(n_419) );
AND2x4_ASAP7_75t_L g420 ( .A(n_373), .B(n_297), .Y(n_420) );
OR2x2_ASAP7_75t_L g421 ( .A(n_372), .B(n_297), .Y(n_421) );
AND2x2_ASAP7_75t_L g422 ( .A(n_363), .B(n_297), .Y(n_422) );
INVx3_ASAP7_75t_L g423 ( .A(n_373), .Y(n_423) );
NAND2xp5_ASAP7_75t_L g424 ( .A(n_372), .B(n_282), .Y(n_424) );
AND2x2_ASAP7_75t_L g425 ( .A(n_363), .B(n_297), .Y(n_425) );
AND2x2_ASAP7_75t_L g426 ( .A(n_365), .B(n_323), .Y(n_426) );
AND2x4_ASAP7_75t_SL g427 ( .A(n_373), .B(n_324), .Y(n_427) );
OR2x2_ASAP7_75t_L g428 ( .A(n_365), .B(n_343), .Y(n_428) );
INVx2_ASAP7_75t_L g429 ( .A(n_340), .Y(n_429) );
INVx1_ASAP7_75t_L g430 ( .A(n_347), .Y(n_430) );
AND2x4_ASAP7_75t_L g431 ( .A(n_373), .B(n_324), .Y(n_431) );
NAND2xp5_ASAP7_75t_L g432 ( .A(n_336), .B(n_324), .Y(n_432) );
AND2x2_ASAP7_75t_L g433 ( .A(n_338), .B(n_323), .Y(n_433) );
AND2x2_ASAP7_75t_L g434 ( .A(n_338), .B(n_323), .Y(n_434) );
AND2x4_ASAP7_75t_L g435 ( .A(n_338), .B(n_324), .Y(n_435) );
OR2x2_ASAP7_75t_L g436 ( .A(n_343), .B(n_324), .Y(n_436) );
AND2x2_ASAP7_75t_L g437 ( .A(n_338), .B(n_323), .Y(n_437) );
AND2x2_ASAP7_75t_L g438 ( .A(n_344), .B(n_323), .Y(n_438) );
NOR2xp33_ASAP7_75t_L g439 ( .A(n_374), .B(n_10), .Y(n_439) );
OR2x2_ASAP7_75t_L g440 ( .A(n_346), .B(n_324), .Y(n_440) );
AND2x2_ASAP7_75t_L g441 ( .A(n_344), .B(n_323), .Y(n_441) );
INVx2_ASAP7_75t_L g442 ( .A(n_340), .Y(n_442) );
NOR2xp33_ASAP7_75t_L g443 ( .A(n_374), .B(n_12), .Y(n_443) );
NAND2xp5_ASAP7_75t_L g444 ( .A(n_352), .B(n_324), .Y(n_444) );
INVx1_ASAP7_75t_L g445 ( .A(n_341), .Y(n_445) );
AND2x2_ASAP7_75t_L g446 ( .A(n_380), .B(n_313), .Y(n_446) );
NAND2xp5_ASAP7_75t_L g447 ( .A(n_352), .B(n_313), .Y(n_447) );
CKINVDCx6p67_ASAP7_75t_R g448 ( .A(n_330), .Y(n_448) );
NOR2xp33_ASAP7_75t_L g449 ( .A(n_379), .B(n_13), .Y(n_449) );
AOI22xp33_ASAP7_75t_L g450 ( .A1(n_352), .A2(n_319), .B1(n_273), .B2(n_309), .Y(n_450) );
INVx1_ASAP7_75t_L g451 ( .A(n_379), .Y(n_451) );
AND2x2_ASAP7_75t_L g452 ( .A(n_380), .B(n_313), .Y(n_452) );
NAND2x1p5_ASAP7_75t_L g453 ( .A(n_391), .B(n_355), .Y(n_453) );
INVx2_ASAP7_75t_L g454 ( .A(n_416), .Y(n_454) );
AND2x2_ASAP7_75t_L g455 ( .A(n_389), .B(n_344), .Y(n_455) );
AND2x2_ASAP7_75t_L g456 ( .A(n_394), .B(n_346), .Y(n_456) );
OR2x6_ASAP7_75t_L g457 ( .A(n_393), .B(n_355), .Y(n_457) );
AND2x2_ASAP7_75t_L g458 ( .A(n_395), .B(n_380), .Y(n_458) );
AND2x2_ASAP7_75t_L g459 ( .A(n_396), .B(n_354), .Y(n_459) );
INVx2_ASAP7_75t_L g460 ( .A(n_416), .Y(n_460) );
AND2x2_ASAP7_75t_L g461 ( .A(n_399), .B(n_354), .Y(n_461) );
OR2x2_ASAP7_75t_L g462 ( .A(n_409), .B(n_367), .Y(n_462) );
NAND2xp5_ASAP7_75t_L g463 ( .A(n_446), .B(n_357), .Y(n_463) );
NAND2xp5_ASAP7_75t_L g464 ( .A(n_452), .B(n_357), .Y(n_464) );
AND2x2_ASAP7_75t_L g465 ( .A(n_413), .B(n_357), .Y(n_465) );
OR2x2_ASAP7_75t_L g466 ( .A(n_404), .B(n_367), .Y(n_466) );
AND2x2_ASAP7_75t_L g467 ( .A(n_404), .B(n_359), .Y(n_467) );
INVx1_ASAP7_75t_L g468 ( .A(n_430), .Y(n_468) );
AND3x2_ASAP7_75t_L g469 ( .A(n_397), .B(n_349), .C(n_351), .Y(n_469) );
NAND2xp5_ASAP7_75t_L g470 ( .A(n_421), .B(n_349), .Y(n_470) );
AND2x4_ASAP7_75t_L g471 ( .A(n_435), .B(n_328), .Y(n_471) );
OR2x2_ASAP7_75t_L g472 ( .A(n_408), .B(n_376), .Y(n_472) );
AND2x2_ASAP7_75t_L g473 ( .A(n_402), .B(n_349), .Y(n_473) );
AND2x4_ASAP7_75t_L g474 ( .A(n_435), .B(n_328), .Y(n_474) );
AND2x2_ASAP7_75t_L g475 ( .A(n_412), .B(n_351), .Y(n_475) );
AND2x2_ASAP7_75t_L g476 ( .A(n_385), .B(n_351), .Y(n_476) );
NAND2xp5_ASAP7_75t_L g477 ( .A(n_451), .B(n_381), .Y(n_477) );
INVx2_ASAP7_75t_SL g478 ( .A(n_391), .Y(n_478) );
NAND2xp5_ASAP7_75t_L g479 ( .A(n_447), .B(n_381), .Y(n_479) );
OR2x2_ASAP7_75t_L g480 ( .A(n_386), .B(n_376), .Y(n_480) );
NAND2xp5_ASAP7_75t_L g481 ( .A(n_414), .B(n_328), .Y(n_481) );
OR2x2_ASAP7_75t_L g482 ( .A(n_390), .B(n_350), .Y(n_482) );
NAND2xp5_ASAP7_75t_L g483 ( .A(n_417), .B(n_350), .Y(n_483) );
AND3x2_ASAP7_75t_L g484 ( .A(n_397), .B(n_360), .C(n_356), .Y(n_484) );
HB1xp67_ASAP7_75t_L g485 ( .A(n_382), .Y(n_485) );
NAND2xp5_ASAP7_75t_L g486 ( .A(n_405), .B(n_356), .Y(n_486) );
NAND2xp5_ASAP7_75t_L g487 ( .A(n_445), .B(n_360), .Y(n_487) );
AND2x4_ASAP7_75t_L g488 ( .A(n_435), .B(n_348), .Y(n_488) );
AND2x2_ASAP7_75t_L g489 ( .A(n_406), .B(n_340), .Y(n_489) );
INVx1_ASAP7_75t_L g490 ( .A(n_428), .Y(n_490) );
OR2x2_ASAP7_75t_L g491 ( .A(n_400), .B(n_345), .Y(n_491) );
AND2x2_ASAP7_75t_L g492 ( .A(n_422), .B(n_345), .Y(n_492) );
NAND2xp5_ASAP7_75t_L g493 ( .A(n_411), .B(n_358), .Y(n_493) );
AND2x2_ASAP7_75t_L g494 ( .A(n_425), .B(n_358), .Y(n_494) );
AND2x4_ASAP7_75t_L g495 ( .A(n_383), .B(n_348), .Y(n_495) );
AND2x2_ASAP7_75t_L g496 ( .A(n_415), .B(n_358), .Y(n_496) );
AND2x2_ASAP7_75t_L g497 ( .A(n_415), .B(n_361), .Y(n_497) );
AND2x4_ASAP7_75t_L g498 ( .A(n_383), .B(n_348), .Y(n_498) );
NAND2xp5_ASAP7_75t_L g499 ( .A(n_382), .B(n_361), .Y(n_499) );
BUFx3_ASAP7_75t_L g500 ( .A(n_448), .Y(n_500) );
AND2x2_ASAP7_75t_L g501 ( .A(n_432), .B(n_361), .Y(n_501) );
OR2x2_ASAP7_75t_L g502 ( .A(n_444), .B(n_370), .Y(n_502) );
NAND2xp5_ASAP7_75t_L g503 ( .A(n_388), .B(n_368), .Y(n_503) );
INVx1_ASAP7_75t_L g504 ( .A(n_398), .Y(n_504) );
NAND2xp5_ASAP7_75t_L g505 ( .A(n_388), .B(n_368), .Y(n_505) );
AND2x2_ASAP7_75t_L g506 ( .A(n_438), .B(n_368), .Y(n_506) );
INVx2_ASAP7_75t_L g507 ( .A(n_407), .Y(n_507) );
NAND2xp5_ASAP7_75t_L g508 ( .A(n_426), .B(n_370), .Y(n_508) );
INVx2_ASAP7_75t_L g509 ( .A(n_407), .Y(n_509) );
INVxp67_ASAP7_75t_L g510 ( .A(n_418), .Y(n_510) );
AND2x2_ASAP7_75t_L g511 ( .A(n_441), .B(n_370), .Y(n_511) );
INVx2_ASAP7_75t_L g512 ( .A(n_410), .Y(n_512) );
BUFx2_ASAP7_75t_L g513 ( .A(n_448), .Y(n_513) );
NOR2xp67_ASAP7_75t_SL g514 ( .A(n_423), .B(n_348), .Y(n_514) );
OR2x2_ASAP7_75t_L g515 ( .A(n_436), .B(n_366), .Y(n_515) );
INVx2_ASAP7_75t_L g516 ( .A(n_410), .Y(n_516) );
NAND2x1p5_ASAP7_75t_L g517 ( .A(n_423), .B(n_366), .Y(n_517) );
AND2x2_ASAP7_75t_L g518 ( .A(n_387), .B(n_366), .Y(n_518) );
NOR2xp33_ASAP7_75t_L g519 ( .A(n_384), .B(n_15), .Y(n_519) );
AND2x4_ASAP7_75t_L g520 ( .A(n_418), .B(n_348), .Y(n_520) );
HB1xp67_ASAP7_75t_L g521 ( .A(n_440), .Y(n_521) );
AND2x2_ASAP7_75t_L g522 ( .A(n_387), .B(n_313), .Y(n_522) );
OR2x2_ASAP7_75t_L g523 ( .A(n_419), .B(n_313), .Y(n_523) );
OAI211xp5_ASAP7_75t_L g524 ( .A1(n_403), .A2(n_319), .B(n_309), .C(n_273), .Y(n_524) );
NAND2xp5_ASAP7_75t_L g525 ( .A(n_429), .B(n_309), .Y(n_525) );
AND2x2_ASAP7_75t_L g526 ( .A(n_392), .B(n_309), .Y(n_526) );
OAI21xp5_ASAP7_75t_L g527 ( .A1(n_453), .A2(n_449), .B(n_443), .Y(n_527) );
NAND2xp5_ASAP7_75t_L g528 ( .A(n_476), .B(n_449), .Y(n_528) );
INVx1_ASAP7_75t_SL g529 ( .A(n_513), .Y(n_529) );
OAI21xp5_ASAP7_75t_L g530 ( .A1(n_453), .A2(n_443), .B(n_439), .Y(n_530) );
NAND2xp5_ASAP7_75t_L g531 ( .A(n_470), .B(n_418), .Y(n_531) );
INVx1_ASAP7_75t_SL g532 ( .A(n_521), .Y(n_532) );
OAI22xp5_ASAP7_75t_L g533 ( .A1(n_478), .A2(n_439), .B1(n_424), .B2(n_423), .Y(n_533) );
AND2x2_ASAP7_75t_L g534 ( .A(n_467), .B(n_461), .Y(n_534) );
NAND2xp5_ASAP7_75t_L g535 ( .A(n_470), .B(n_420), .Y(n_535) );
AOI22xp5_ASAP7_75t_L g536 ( .A1(n_519), .A2(n_420), .B1(n_431), .B2(n_401), .Y(n_536) );
INVx2_ASAP7_75t_SL g537 ( .A(n_500), .Y(n_537) );
INVx1_ASAP7_75t_SL g538 ( .A(n_485), .Y(n_538) );
NAND2xp5_ASAP7_75t_L g539 ( .A(n_490), .B(n_392), .Y(n_539) );
AND2x2_ASAP7_75t_SL g540 ( .A(n_455), .B(n_433), .Y(n_540) );
NAND2xp5_ASAP7_75t_L g541 ( .A(n_463), .B(n_442), .Y(n_541) );
INVx2_ASAP7_75t_L g542 ( .A(n_472), .Y(n_542) );
AND2x2_ASAP7_75t_L g543 ( .A(n_465), .B(n_401), .Y(n_543) );
NAND2xp5_ASAP7_75t_L g544 ( .A(n_473), .B(n_450), .Y(n_544) );
INVx2_ASAP7_75t_SL g545 ( .A(n_456), .Y(n_545) );
OR2x2_ASAP7_75t_L g546 ( .A(n_463), .B(n_427), .Y(n_546) );
INVx1_ASAP7_75t_L g547 ( .A(n_468), .Y(n_547) );
AND2x2_ASAP7_75t_L g548 ( .A(n_459), .B(n_437), .Y(n_548) );
AOI322xp5_ASAP7_75t_L g549 ( .A1(n_464), .A2(n_450), .A3(n_434), .B1(n_134), .B2(n_16), .C1(n_18), .C2(n_19), .Y(n_549) );
INVxp67_ASAP7_75t_L g550 ( .A(n_485), .Y(n_550) );
OR2x2_ASAP7_75t_L g551 ( .A(n_464), .B(n_309), .Y(n_551) );
AND2x4_ASAP7_75t_L g552 ( .A(n_471), .B(n_321), .Y(n_552) );
HB1xp67_ASAP7_75t_L g553 ( .A(n_454), .Y(n_553) );
NOR5xp2_ASAP7_75t_L g554 ( .A(n_524), .B(n_16), .C(n_18), .D(n_19), .E(n_309), .Y(n_554) );
HB1xp67_ASAP7_75t_L g555 ( .A(n_460), .Y(n_555) );
AOI221xp5_ASAP7_75t_L g556 ( .A1(n_510), .A2(n_289), .B1(n_163), .B2(n_152), .C(n_26), .Y(n_556) );
INVx1_ASAP7_75t_SL g557 ( .A(n_471), .Y(n_557) );
NAND2xp5_ASAP7_75t_L g558 ( .A(n_475), .B(n_321), .Y(n_558) );
INVx2_ASAP7_75t_SL g559 ( .A(n_466), .Y(n_559) );
INVx2_ASAP7_75t_L g560 ( .A(n_496), .Y(n_560) );
OAI22xp33_ASAP7_75t_L g561 ( .A1(n_457), .A2(n_273), .B1(n_289), .B2(n_25), .Y(n_561) );
AND2x2_ASAP7_75t_L g562 ( .A(n_458), .B(n_23), .Y(n_562) );
NAND2xp5_ASAP7_75t_L g563 ( .A(n_504), .B(n_24), .Y(n_563) );
OR2x2_ASAP7_75t_L g564 ( .A(n_479), .B(n_27), .Y(n_564) );
AND2x2_ASAP7_75t_L g565 ( .A(n_474), .B(n_28), .Y(n_565) );
AND2x2_ASAP7_75t_L g566 ( .A(n_474), .B(n_30), .Y(n_566) );
INVx2_ASAP7_75t_SL g567 ( .A(n_462), .Y(n_567) );
INVx1_ASAP7_75t_L g568 ( .A(n_486), .Y(n_568) );
INVx2_ASAP7_75t_L g569 ( .A(n_497), .Y(n_569) );
NAND2xp5_ASAP7_75t_L g570 ( .A(n_479), .B(n_31), .Y(n_570) );
NAND2xp5_ASAP7_75t_SL g571 ( .A(n_495), .B(n_498), .Y(n_571) );
INVx1_ASAP7_75t_L g572 ( .A(n_486), .Y(n_572) );
INVx2_ASAP7_75t_L g573 ( .A(n_518), .Y(n_573) );
AND2x2_ASAP7_75t_L g574 ( .A(n_489), .B(n_32), .Y(n_574) );
NAND2xp5_ASAP7_75t_L g575 ( .A(n_477), .B(n_33), .Y(n_575) );
NAND2xp5_ASAP7_75t_L g576 ( .A(n_477), .B(n_34), .Y(n_576) );
INVx1_ASAP7_75t_L g577 ( .A(n_482), .Y(n_577) );
INVx2_ASAP7_75t_L g578 ( .A(n_506), .Y(n_578) );
AND2x2_ASAP7_75t_L g579 ( .A(n_492), .B(n_38), .Y(n_579) );
OAI21xp5_ASAP7_75t_L g580 ( .A1(n_549), .A2(n_457), .B(n_524), .Y(n_580) );
BUFx2_ASAP7_75t_L g581 ( .A(n_529), .Y(n_581) );
INVx2_ASAP7_75t_L g582 ( .A(n_538), .Y(n_582) );
INVx2_ASAP7_75t_SL g583 ( .A(n_537), .Y(n_583) );
OAI21xp5_ASAP7_75t_L g584 ( .A1(n_533), .A2(n_457), .B(n_487), .Y(n_584) );
INVx1_ASAP7_75t_L g585 ( .A(n_568), .Y(n_585) );
NOR3xp33_ASAP7_75t_L g586 ( .A(n_533), .B(n_487), .C(n_493), .Y(n_586) );
INVx1_ASAP7_75t_L g587 ( .A(n_572), .Y(n_587) );
AOI22xp33_ASAP7_75t_L g588 ( .A1(n_544), .A2(n_469), .B1(n_522), .B2(n_481), .Y(n_588) );
OR2x2_ASAP7_75t_L g589 ( .A(n_531), .B(n_481), .Y(n_589) );
OAI32xp33_ASAP7_75t_L g590 ( .A1(n_557), .A2(n_517), .A3(n_480), .B1(n_491), .B2(n_508), .Y(n_590) );
NAND4xp25_ASAP7_75t_L g591 ( .A(n_527), .B(n_520), .C(n_526), .D(n_508), .Y(n_591) );
O2A1O1Ixp33_ASAP7_75t_L g592 ( .A1(n_527), .A2(n_493), .B(n_483), .C(n_523), .Y(n_592) );
AO22x1_ASAP7_75t_L g593 ( .A1(n_557), .A2(n_488), .B1(n_484), .B2(n_520), .Y(n_593) );
OR2x2_ASAP7_75t_L g594 ( .A(n_531), .B(n_502), .Y(n_594) );
A2O1A1Ixp33_ASAP7_75t_L g595 ( .A1(n_530), .A2(n_488), .B(n_514), .C(n_494), .Y(n_595) );
AOI32xp33_ASAP7_75t_L g596 ( .A1(n_532), .A2(n_511), .A3(n_501), .B1(n_499), .B2(n_515), .Y(n_596) );
AOI22xp33_ASAP7_75t_L g597 ( .A1(n_536), .A2(n_517), .B1(n_525), .B2(n_516), .Y(n_597) );
AOI211xp5_ASAP7_75t_SL g598 ( .A1(n_565), .A2(n_525), .B(n_505), .C(n_503), .Y(n_598) );
NAND2xp5_ASAP7_75t_L g599 ( .A(n_532), .B(n_577), .Y(n_599) );
NOR2x1_ASAP7_75t_L g600 ( .A(n_530), .B(n_505), .Y(n_600) );
NAND2xp5_ASAP7_75t_L g601 ( .A(n_535), .B(n_512), .Y(n_601) );
OAI22xp5_ASAP7_75t_L g602 ( .A1(n_540), .A2(n_503), .B1(n_507), .B2(n_509), .Y(n_602) );
OAI32xp33_ASAP7_75t_SL g603 ( .A1(n_567), .A2(n_559), .A3(n_528), .B1(n_535), .B2(n_551), .Y(n_603) );
OAI321xp33_ASAP7_75t_L g604 ( .A1(n_571), .A2(n_152), .A3(n_43), .B1(n_46), .B2(n_47), .C(n_49), .Y(n_604) );
OAI22xp5_ASAP7_75t_L g605 ( .A1(n_545), .A2(n_52), .B1(n_53), .B2(n_55), .Y(n_605) );
INVx1_ASAP7_75t_L g606 ( .A(n_547), .Y(n_606) );
CKINVDCx20_ASAP7_75t_R g607 ( .A(n_539), .Y(n_607) );
AOI21xp33_ASAP7_75t_L g608 ( .A1(n_564), .A2(n_56), .B(n_59), .Y(n_608) );
OAI221xp5_ASAP7_75t_SL g609 ( .A1(n_546), .A2(n_61), .B1(n_62), .B2(n_64), .C(n_66), .Y(n_609) );
INVx1_ASAP7_75t_L g610 ( .A(n_594), .Y(n_610) );
AOI21xp33_ASAP7_75t_L g611 ( .A1(n_580), .A2(n_563), .B(n_570), .Y(n_611) );
OAI21xp5_ASAP7_75t_L g612 ( .A1(n_600), .A2(n_550), .B(n_562), .Y(n_612) );
NAND2x1_ASAP7_75t_L g613 ( .A(n_581), .B(n_552), .Y(n_613) );
INVx1_ASAP7_75t_L g614 ( .A(n_599), .Y(n_614) );
NAND3xp33_ASAP7_75t_L g615 ( .A(n_580), .B(n_554), .C(n_576), .Y(n_615) );
NAND2xp5_ASAP7_75t_SL g616 ( .A(n_584), .B(n_561), .Y(n_616) );
NAND2xp5_ASAP7_75t_SL g617 ( .A(n_584), .B(n_566), .Y(n_617) );
AOI22xp5_ASAP7_75t_L g618 ( .A1(n_591), .A2(n_542), .B1(n_541), .B2(n_558), .Y(n_618) );
INVx1_ASAP7_75t_L g619 ( .A(n_589), .Y(n_619) );
INVx1_ASAP7_75t_L g620 ( .A(n_585), .Y(n_620) );
INVx2_ASAP7_75t_L g621 ( .A(n_582), .Y(n_621) );
NAND2xp5_ASAP7_75t_L g622 ( .A(n_586), .B(n_534), .Y(n_622) );
NAND2xp5_ASAP7_75t_L g623 ( .A(n_592), .B(n_553), .Y(n_623) );
AOI211x1_ASAP7_75t_SL g624 ( .A1(n_595), .A2(n_576), .B(n_575), .C(n_578), .Y(n_624) );
NAND2xp5_ASAP7_75t_L g625 ( .A(n_587), .B(n_555), .Y(n_625) );
NOR2xp33_ASAP7_75t_L g626 ( .A(n_583), .B(n_573), .Y(n_626) );
OAI311xp33_ASAP7_75t_L g627 ( .A1(n_597), .A2(n_556), .A3(n_574), .B1(n_579), .C1(n_548), .Y(n_627) );
OAI21x1_ASAP7_75t_L g628 ( .A1(n_602), .A2(n_560), .B(n_569), .Y(n_628) );
AOI21xp5_ASAP7_75t_L g629 ( .A1(n_593), .A2(n_543), .B(n_67), .Y(n_629) );
A2O1A1Ixp33_ASAP7_75t_L g630 ( .A1(n_596), .A2(n_68), .B(n_70), .C(n_72), .Y(n_630) );
OAI21xp5_ASAP7_75t_L g631 ( .A1(n_598), .A2(n_74), .B(n_79), .Y(n_631) );
OAI21xp5_ASAP7_75t_SL g632 ( .A1(n_598), .A2(n_202), .B(n_605), .Y(n_632) );
AOI211xp5_ASAP7_75t_L g633 ( .A1(n_605), .A2(n_202), .B(n_609), .C(n_608), .Y(n_633) );
NAND2xp5_ASAP7_75t_SL g634 ( .A(n_607), .B(n_601), .Y(n_634) );
AOI221xp5_ASAP7_75t_L g635 ( .A1(n_606), .A2(n_603), .B1(n_592), .B2(n_590), .C(n_591), .Y(n_635) );
OAI321xp33_ASAP7_75t_L g636 ( .A1(n_604), .A2(n_584), .A3(n_580), .B1(n_591), .B2(n_588), .C(n_596), .Y(n_636) );
NAND2xp5_ASAP7_75t_L g637 ( .A(n_624), .B(n_622), .Y(n_637) );
INVx1_ASAP7_75t_L g638 ( .A(n_620), .Y(n_638) );
NOR3xp33_ASAP7_75t_L g639 ( .A(n_636), .B(n_615), .C(n_632), .Y(n_639) );
AND2x2_ASAP7_75t_L g640 ( .A(n_618), .B(n_612), .Y(n_640) );
AOI21xp5_ASAP7_75t_L g641 ( .A1(n_629), .A2(n_616), .B(n_617), .Y(n_641) );
NOR2xp33_ASAP7_75t_SL g642 ( .A(n_630), .B(n_631), .Y(n_642) );
AOI21xp5_ASAP7_75t_L g643 ( .A1(n_641), .A2(n_616), .B(n_613), .Y(n_643) );
AND3x2_ASAP7_75t_L g644 ( .A(n_639), .B(n_633), .C(n_635), .Y(n_644) );
INVx2_ASAP7_75t_L g645 ( .A(n_638), .Y(n_645) );
O2A1O1Ixp5_ASAP7_75t_L g646 ( .A1(n_637), .A2(n_627), .B(n_611), .C(n_617), .Y(n_646) );
INVx1_ASAP7_75t_L g647 ( .A(n_645), .Y(n_647) );
NOR2x1_ASAP7_75t_L g648 ( .A(n_643), .B(n_640), .Y(n_648) );
AND2x2_ASAP7_75t_L g649 ( .A(n_644), .B(n_628), .Y(n_649) );
XOR2xp5_ASAP7_75t_L g650 ( .A(n_648), .B(n_647), .Y(n_650) );
OAI22xp5_ASAP7_75t_L g651 ( .A1(n_649), .A2(n_623), .B1(n_614), .B2(n_626), .Y(n_651) );
AND2x4_ASAP7_75t_L g652 ( .A(n_650), .B(n_626), .Y(n_652) );
INVx2_ASAP7_75t_L g653 ( .A(n_651), .Y(n_653) );
AOI21xp5_ASAP7_75t_L g654 ( .A1(n_653), .A2(n_646), .B(n_642), .Y(n_654) );
AOI21xp5_ASAP7_75t_L g655 ( .A1(n_654), .A2(n_652), .B(n_634), .Y(n_655) );
XNOR2x1_ASAP7_75t_L g656 ( .A(n_655), .B(n_652), .Y(n_656) );
OA21x2_ASAP7_75t_L g657 ( .A1(n_656), .A2(n_610), .B(n_619), .Y(n_657) );
OA21x2_ASAP7_75t_L g658 ( .A1(n_657), .A2(n_625), .B(n_621), .Y(n_658) );
endmodule