module fake_jpeg_362_n_148 (n_13, n_21, n_33, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_19, n_18, n_20, n_35, n_4, n_34, n_30, n_16, n_3, n_0, n_24, n_28, n_26, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_12, n_32, n_8, n_15, n_7, n_148);

input n_13;
input n_21;
input n_33;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_35;
input n_4;
input n_34;
input n_30;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_26;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_148;

wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_147;
wire n_73;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_49;
wire n_76;
wire n_127;
wire n_38;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_103;
wire n_50;
wire n_124;
wire n_141;
wire n_57;
wire n_119;
wire n_69;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_106;
wire n_111;
wire n_44;
wire n_143;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_78;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_128;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_91;
wire n_54;
wire n_93;
wire n_138;
wire n_101;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_97;
wire n_135;
wire n_62;
wire n_120;
wire n_43;
wire n_100;
wire n_118;
wire n_82;
wire n_140;
wire n_96;

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_8),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_27),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_9),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_25),
.Y(n_41)
);

BUFx12_ASAP7_75t_L g42 ( 
.A(n_23),
.Y(n_42)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_13),
.Y(n_43)
);

INVx5_ASAP7_75t_L g44 ( 
.A(n_19),
.Y(n_44)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_15),
.Y(n_45)
);

INVx11_ASAP7_75t_L g46 ( 
.A(n_6),
.Y(n_46)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_35),
.Y(n_47)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_37),
.Y(n_48)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_26),
.Y(n_49)
);

BUFx16f_ASAP7_75t_L g50 ( 
.A(n_12),
.Y(n_50)
);

INVx6_ASAP7_75t_L g51 ( 
.A(n_2),
.Y(n_51)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_3),
.Y(n_52)
);

BUFx12f_ASAP7_75t_L g53 ( 
.A(n_3),
.Y(n_53)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_43),
.Y(n_54)
);

INVx1_ASAP7_75t_SL g70 ( 
.A(n_54),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_38),
.B(n_0),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_55),
.B(n_60),
.Y(n_66)
);

INVx11_ASAP7_75t_L g56 ( 
.A(n_53),
.Y(n_56)
);

CKINVDCx6p67_ASAP7_75t_R g64 ( 
.A(n_56),
.Y(n_64)
);

BUFx5_ASAP7_75t_L g57 ( 
.A(n_50),
.Y(n_57)
);

BUFx3_ASAP7_75t_L g62 ( 
.A(n_57),
.Y(n_62)
);

BUFx12_ASAP7_75t_L g58 ( 
.A(n_50),
.Y(n_58)
);

INVx3_ASAP7_75t_L g65 ( 
.A(n_58),
.Y(n_65)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_40),
.Y(n_59)
);

INVx2_ASAP7_75t_L g63 ( 
.A(n_59),
.Y(n_63)
);

NAND2xp33_ASAP7_75t_SL g60 ( 
.A(n_50),
.B(n_0),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_52),
.B(n_1),
.Y(n_61)
);

INVx2_ASAP7_75t_L g68 ( 
.A(n_61),
.Y(n_68)
);

INVx3_ASAP7_75t_L g67 ( 
.A(n_54),
.Y(n_67)
);

INVx2_ASAP7_75t_SL g79 ( 
.A(n_67),
.Y(n_79)
);

INVx2_ASAP7_75t_L g69 ( 
.A(n_59),
.Y(n_69)
);

INVx2_ASAP7_75t_L g77 ( 
.A(n_69),
.Y(n_77)
);

INVx2_ASAP7_75t_L g71 ( 
.A(n_59),
.Y(n_71)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_71),
.Y(n_74)
);

INVx3_ASAP7_75t_L g72 ( 
.A(n_57),
.Y(n_72)
);

BUFx3_ASAP7_75t_L g80 ( 
.A(n_72),
.Y(n_80)
);

AND2x2_ASAP7_75t_SL g73 ( 
.A(n_68),
.B(n_60),
.Y(n_73)
);

INVx1_ASAP7_75t_SL g101 ( 
.A(n_73),
.Y(n_101)
);

XNOR2xp5_ASAP7_75t_L g75 ( 
.A(n_66),
.B(n_43),
.Y(n_75)
);

MAJIxp5_ASAP7_75t_L g98 ( 
.A(n_75),
.B(n_48),
.C(n_47),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_SL g76 ( 
.A(n_66),
.B(n_61),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_L g92 ( 
.A(n_76),
.B(n_81),
.Y(n_92)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_70),
.Y(n_78)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_78),
.Y(n_94)
);

CKINVDCx20_ASAP7_75t_R g81 ( 
.A(n_64),
.Y(n_81)
);

OAI22xp5_ASAP7_75t_L g82 ( 
.A1(n_63),
.A2(n_51),
.B1(n_40),
.B2(n_46),
.Y(n_82)
);

OAI22xp5_ASAP7_75t_L g90 ( 
.A1(n_82),
.A2(n_51),
.B1(n_44),
.B2(n_53),
.Y(n_90)
);

INVx8_ASAP7_75t_L g83 ( 
.A(n_64),
.Y(n_83)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_83),
.Y(n_95)
);

AOI22xp33_ASAP7_75t_SL g84 ( 
.A1(n_62),
.A2(n_56),
.B1(n_53),
.B2(n_46),
.Y(n_84)
);

AOI22xp33_ASAP7_75t_SL g99 ( 
.A1(n_84),
.A2(n_58),
.B1(n_44),
.B2(n_49),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g85 ( 
.A(n_65),
.B(n_55),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_L g93 ( 
.A(n_85),
.B(n_86),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_L g86 ( 
.A(n_64),
.B(n_41),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_75),
.B(n_45),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_L g109 ( 
.A(n_87),
.B(n_102),
.Y(n_109)
);

OAI22xp5_ASAP7_75t_SL g88 ( 
.A1(n_73),
.A2(n_84),
.B1(n_79),
.B2(n_74),
.Y(n_88)
);

AOI22xp5_ASAP7_75t_L g110 ( 
.A1(n_88),
.A2(n_90),
.B1(n_89),
.B2(n_101),
.Y(n_110)
);

AND2x4_ASAP7_75t_L g89 ( 
.A(n_73),
.B(n_58),
.Y(n_89)
);

CKINVDCx16_ASAP7_75t_R g103 ( 
.A(n_89),
.Y(n_103)
);

AOI21xp5_ASAP7_75t_L g91 ( 
.A1(n_79),
.A2(n_41),
.B(n_45),
.Y(n_91)
);

OA21x2_ASAP7_75t_L g119 ( 
.A1(n_91),
.A2(n_5),
.B(n_6),
.Y(n_119)
);

AOI21xp33_ASAP7_75t_L g96 ( 
.A1(n_83),
.A2(n_42),
.B(n_2),
.Y(n_96)
);

FAx1_ASAP7_75t_SL g118 ( 
.A(n_96),
.B(n_1),
.CI(n_4),
.CON(n_118),
.SN(n_118)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_77),
.Y(n_97)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_97),
.Y(n_104)
);

XNOR2xp5_ASAP7_75t_L g106 ( 
.A(n_98),
.B(n_58),
.Y(n_106)
);

OAI22xp5_ASAP7_75t_L g108 ( 
.A1(n_99),
.A2(n_42),
.B1(n_4),
.B2(n_5),
.Y(n_108)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_77),
.Y(n_100)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_100),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g102 ( 
.A(n_80),
.B(n_39),
.Y(n_102)
);

AND2x6_ASAP7_75t_L g105 ( 
.A(n_89),
.B(n_21),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_L g128 ( 
.A(n_105),
.B(n_112),
.Y(n_128)
);

MAJIxp5_ASAP7_75t_L g124 ( 
.A(n_106),
.B(n_111),
.C(n_113),
.Y(n_124)
);

AOI22x1_ASAP7_75t_L g107 ( 
.A1(n_88),
.A2(n_80),
.B1(n_42),
.B2(n_20),
.Y(n_107)
);

OA22x2_ASAP7_75t_L g121 ( 
.A1(n_107),
.A2(n_7),
.B1(n_8),
.B2(n_9),
.Y(n_121)
);

INVxp67_ASAP7_75t_L g131 ( 
.A(n_108),
.Y(n_131)
);

OAI22xp5_ASAP7_75t_SL g123 ( 
.A1(n_110),
.A2(n_116),
.B1(n_24),
.B2(n_32),
.Y(n_123)
);

MAJIxp5_ASAP7_75t_L g111 ( 
.A(n_101),
.B(n_17),
.C(n_34),
.Y(n_111)
);

CKINVDCx20_ASAP7_75t_R g112 ( 
.A(n_92),
.Y(n_112)
);

MAJIxp5_ASAP7_75t_L g113 ( 
.A(n_93),
.B(n_16),
.C(n_33),
.Y(n_113)
);

INVx13_ASAP7_75t_L g115 ( 
.A(n_95),
.Y(n_115)
);

INVx1_ASAP7_75t_SL g126 ( 
.A(n_115),
.Y(n_126)
);

OAI22xp5_ASAP7_75t_SL g116 ( 
.A1(n_99),
.A2(n_89),
.B1(n_94),
.B2(n_98),
.Y(n_116)
);

INVx13_ASAP7_75t_L g117 ( 
.A(n_95),
.Y(n_117)
);

BUFx5_ASAP7_75t_L g127 ( 
.A(n_117),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_L g129 ( 
.A(n_118),
.B(n_119),
.Y(n_129)
);

CKINVDCx20_ASAP7_75t_R g120 ( 
.A(n_115),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_L g133 ( 
.A(n_120),
.B(n_121),
.Y(n_133)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_104),
.Y(n_122)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_122),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_SL g135 ( 
.A(n_123),
.B(n_119),
.Y(n_135)
);

AOI21xp5_ASAP7_75t_SL g125 ( 
.A1(n_103),
.A2(n_7),
.B(n_10),
.Y(n_125)
);

AOI21xp5_ASAP7_75t_L g132 ( 
.A1(n_125),
.A2(n_130),
.B(n_107),
.Y(n_132)
);

OAI22x1_ASAP7_75t_L g130 ( 
.A1(n_103),
.A2(n_28),
.B1(n_31),
.B2(n_14),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_SL g138 ( 
.A(n_132),
.B(n_135),
.Y(n_138)
);

XOR2xp5_ASAP7_75t_L g136 ( 
.A(n_124),
.B(n_109),
.Y(n_136)
);

XOR2xp5_ASAP7_75t_L g139 ( 
.A(n_136),
.B(n_125),
.Y(n_139)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_134),
.Y(n_137)
);

AOI22xp5_ASAP7_75t_L g141 ( 
.A1(n_137),
.A2(n_139),
.B1(n_136),
.B2(n_126),
.Y(n_141)
);

AOI22xp5_ASAP7_75t_SL g140 ( 
.A1(n_138),
.A2(n_133),
.B1(n_130),
.B2(n_131),
.Y(n_140)
);

OAI22xp5_ASAP7_75t_SL g142 ( 
.A1(n_140),
.A2(n_141),
.B1(n_129),
.B2(n_131),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_SL g143 ( 
.A(n_142),
.B(n_121),
.Y(n_143)
);

OAI21xp5_ASAP7_75t_SL g144 ( 
.A1(n_143),
.A2(n_128),
.B(n_121),
.Y(n_144)
);

OAI22xp5_ASAP7_75t_SL g145 ( 
.A1(n_144),
.A2(n_118),
.B1(n_114),
.B2(n_18),
.Y(n_145)
);

AOI322xp5_ASAP7_75t_L g146 ( 
.A1(n_145),
.A2(n_117),
.A3(n_127),
.B1(n_22),
.B2(n_29),
.C1(n_30),
.C2(n_36),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_L g147 ( 
.A(n_146),
.B(n_10),
.Y(n_147)
);

XNOR2xp5_ASAP7_75t_L g148 ( 
.A(n_147),
.B(n_11),
.Y(n_148)
);


endmodule