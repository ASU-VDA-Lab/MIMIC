module fake_jpeg_9899_n_125 (n_13, n_21, n_33, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_40, n_19, n_18, n_20, n_35, n_41, n_4, n_34, n_30, n_39, n_42, n_16, n_3, n_0, n_24, n_28, n_38, n_26, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_43, n_12, n_32, n_8, n_15, n_7, n_125);

input n_13;
input n_21;
input n_33;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_42;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_43;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_125;

wire n_117;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_73;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_49;
wire n_76;
wire n_88;
wire n_116;
wire n_114;
wire n_74;
wire n_103;
wire n_50;
wire n_124;
wire n_57;
wire n_119;
wire n_69;
wire n_83;
wire n_71;
wire n_80;
wire n_81;
wire n_109;
wire n_113;
wire n_106;
wire n_111;
wire n_44;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_121;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_56;
wire n_79;
wire n_67;
wire n_53;
wire n_54;
wire n_91;
wire n_93;
wire n_101;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_97;
wire n_62;
wire n_120;
wire n_100;
wire n_118;
wire n_82;
wire n_96;

INVx1_ASAP7_75t_L g44 ( 
.A(n_29),
.Y(n_44)
);

BUFx6f_ASAP7_75t_SL g45 ( 
.A(n_21),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_26),
.Y(n_46)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_23),
.Y(n_47)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_0),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_30),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_8),
.Y(n_50)
);

BUFx12f_ASAP7_75t_L g51 ( 
.A(n_15),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_32),
.Y(n_52)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_38),
.Y(n_53)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_35),
.Y(n_54)
);

CKINVDCx5p33_ASAP7_75t_R g55 ( 
.A(n_9),
.Y(n_55)
);

BUFx12f_ASAP7_75t_L g56 ( 
.A(n_27),
.Y(n_56)
);

BUFx2_ASAP7_75t_L g57 ( 
.A(n_25),
.Y(n_57)
);

CKINVDCx20_ASAP7_75t_R g58 ( 
.A(n_33),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_37),
.Y(n_59)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_18),
.Y(n_60)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_34),
.Y(n_61)
);

BUFx5_ASAP7_75t_L g62 ( 
.A(n_14),
.Y(n_62)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_11),
.Y(n_63)
);

BUFx12f_ASAP7_75t_L g64 ( 
.A(n_45),
.Y(n_64)
);

INVx4_ASAP7_75t_L g85 ( 
.A(n_64),
.Y(n_85)
);

INVx5_ASAP7_75t_L g65 ( 
.A(n_62),
.Y(n_65)
);

INVx5_ASAP7_75t_L g88 ( 
.A(n_65),
.Y(n_88)
);

INVx8_ASAP7_75t_L g66 ( 
.A(n_57),
.Y(n_66)
);

INVx3_ASAP7_75t_SL g90 ( 
.A(n_66),
.Y(n_90)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_51),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_SL g68 ( 
.A(n_48),
.B(n_0),
.Y(n_68)
);

AND2x2_ASAP7_75t_L g81 ( 
.A(n_68),
.B(n_2),
.Y(n_81)
);

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_51),
.Y(n_69)
);

BUFx6f_ASAP7_75t_L g83 ( 
.A(n_69),
.Y(n_83)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_57),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_70),
.B(n_73),
.Y(n_74)
);

BUFx12f_ASAP7_75t_L g71 ( 
.A(n_56),
.Y(n_71)
);

BUFx2_ASAP7_75t_L g72 ( 
.A(n_56),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_L g73 ( 
.A(n_50),
.B(n_1),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_L g75 ( 
.A(n_68),
.B(n_55),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_L g94 ( 
.A(n_75),
.B(n_80),
.Y(n_94)
);

AOI22xp5_ASAP7_75t_L g76 ( 
.A1(n_67),
.A2(n_63),
.B1(n_61),
.B2(n_60),
.Y(n_76)
);

OAI22xp5_ASAP7_75t_SL g100 ( 
.A1(n_76),
.A2(n_77),
.B1(n_78),
.B2(n_82),
.Y(n_100)
);

AOI22xp5_ASAP7_75t_SL g77 ( 
.A1(n_72),
.A2(n_58),
.B1(n_54),
.B2(n_44),
.Y(n_77)
);

OAI22xp33_ASAP7_75t_SL g78 ( 
.A1(n_64),
.A2(n_59),
.B1(n_52),
.B2(n_49),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_71),
.B(n_1),
.Y(n_79)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_79),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_L g80 ( 
.A(n_69),
.B(n_2),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_L g96 ( 
.A(n_81),
.B(n_89),
.Y(n_96)
);

AOI22xp33_ASAP7_75t_L g82 ( 
.A1(n_66),
.A2(n_59),
.B1(n_52),
.B2(n_49),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_SL g84 ( 
.A(n_68),
.B(n_53),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_SL g104 ( 
.A(n_84),
.B(n_86),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_73),
.B(n_3),
.Y(n_86)
);

AOI22xp5_ASAP7_75t_SL g87 ( 
.A1(n_65),
.A2(n_47),
.B1(n_46),
.B2(n_5),
.Y(n_87)
);

OAI22xp5_ASAP7_75t_SL g101 ( 
.A1(n_87),
.A2(n_92),
.B1(n_13),
.B2(n_16),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_73),
.B(n_3),
.Y(n_89)
);

INVx2_ASAP7_75t_L g91 ( 
.A(n_65),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_L g102 ( 
.A(n_91),
.B(n_17),
.Y(n_102)
);

AOI22xp33_ASAP7_75t_SL g92 ( 
.A1(n_66),
.A2(n_4),
.B1(n_5),
.B2(n_6),
.Y(n_92)
);

AOI22xp33_ASAP7_75t_SL g93 ( 
.A1(n_88),
.A2(n_4),
.B1(n_6),
.B2(n_7),
.Y(n_93)
);

OAI21xp5_ASAP7_75t_SL g107 ( 
.A1(n_93),
.A2(n_97),
.B(n_98),
.Y(n_107)
);

OAI22xp5_ASAP7_75t_L g95 ( 
.A1(n_74),
.A2(n_24),
.B1(n_42),
.B2(n_41),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g108 ( 
.A(n_95),
.B(n_99),
.Y(n_108)
);

AND2x2_ASAP7_75t_SL g97 ( 
.A(n_90),
.B(n_7),
.Y(n_97)
);

OR2x4_ASAP7_75t_L g98 ( 
.A(n_74),
.B(n_8),
.Y(n_98)
);

AOI22xp5_ASAP7_75t_L g99 ( 
.A1(n_86),
.A2(n_9),
.B1(n_10),
.B2(n_12),
.Y(n_99)
);

AOI22xp5_ASAP7_75t_SL g103 ( 
.A1(n_82),
.A2(n_19),
.B1(n_20),
.B2(n_22),
.Y(n_103)
);

INVx4_ASAP7_75t_L g106 ( 
.A(n_85),
.Y(n_106)
);

OAI22xp5_ASAP7_75t_SL g109 ( 
.A1(n_108),
.A2(n_100),
.B1(n_103),
.B2(n_93),
.Y(n_109)
);

OAI22xp5_ASAP7_75t_SL g111 ( 
.A1(n_109),
.A2(n_110),
.B1(n_98),
.B2(n_105),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_SL g110 ( 
.A(n_107),
.B(n_104),
.Y(n_110)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_111),
.Y(n_112)
);

OAI21xp5_ASAP7_75t_L g113 ( 
.A1(n_112),
.A2(n_97),
.B(n_96),
.Y(n_113)
);

INVxp67_ASAP7_75t_L g114 ( 
.A(n_113),
.Y(n_114)
);

XNOR2xp5_ASAP7_75t_L g115 ( 
.A(n_114),
.B(n_109),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_L g116 ( 
.A(n_115),
.B(n_101),
.Y(n_116)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_116),
.Y(n_117)
);

MAJIxp5_ASAP7_75t_L g118 ( 
.A(n_117),
.B(n_28),
.C(n_31),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_L g119 ( 
.A(n_118),
.B(n_36),
.Y(n_119)
);

MAJIxp5_ASAP7_75t_L g120 ( 
.A(n_119),
.B(n_102),
.C(n_40),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_L g121 ( 
.A(n_120),
.B(n_39),
.Y(n_121)
);

OAI21x1_ASAP7_75t_SL g122 ( 
.A1(n_121),
.A2(n_43),
.B(n_83),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_SL g123 ( 
.A(n_122),
.B(n_106),
.Y(n_123)
);

NAND3xp33_ASAP7_75t_SL g124 ( 
.A(n_123),
.B(n_79),
.C(n_89),
.Y(n_124)
);

XNOR2xp5_ASAP7_75t_L g125 ( 
.A(n_124),
.B(n_94),
.Y(n_125)
);


endmodule