module fake_jpeg_122_n_244 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_244);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_244;

wire n_159;
wire n_117;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_84;
wire n_59;
wire n_98;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_223;
wire n_234;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_44;
wire n_24;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_122;
wire n_75;
wire n_37;
wire n_233;
wire n_121;
wire n_99;
wire n_130;
wire n_102;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_232;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_170;
wire n_162;
wire n_132;
wire n_133;
wire n_67;
wire n_217;
wire n_216;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_48;
wire n_35;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_118;
wire n_100;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

INVx4_ASAP7_75t_L g17 ( 
.A(n_14),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_10),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_8),
.Y(n_19)
);

NOR2xp33_ASAP7_75t_L g20 ( 
.A(n_7),
.B(n_15),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_13),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_4),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_9),
.Y(n_23)
);

INVx5_ASAP7_75t_L g24 ( 
.A(n_16),
.Y(n_24)
);

BUFx10_ASAP7_75t_L g25 ( 
.A(n_5),
.Y(n_25)
);

INVx13_ASAP7_75t_L g26 ( 
.A(n_10),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_15),
.Y(n_27)
);

INVx2_ASAP7_75t_L g28 ( 
.A(n_13),
.Y(n_28)
);

NOR2xp33_ASAP7_75t_L g29 ( 
.A(n_1),
.B(n_14),
.Y(n_29)
);

INVx13_ASAP7_75t_L g30 ( 
.A(n_1),
.Y(n_30)
);

NOR2xp33_ASAP7_75t_SL g31 ( 
.A(n_16),
.B(n_4),
.Y(n_31)
);

INVx8_ASAP7_75t_L g32 ( 
.A(n_1),
.Y(n_32)
);

BUFx10_ASAP7_75t_L g33 ( 
.A(n_9),
.Y(n_33)
);

INVx1_ASAP7_75t_SL g34 ( 
.A(n_9),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_4),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_8),
.Y(n_36)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_2),
.Y(n_37)
);

BUFx3_ASAP7_75t_L g38 ( 
.A(n_12),
.Y(n_38)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_0),
.Y(n_39)
);

INVx11_ASAP7_75t_L g40 ( 
.A(n_30),
.Y(n_40)
);

INVx11_ASAP7_75t_L g99 ( 
.A(n_40),
.Y(n_99)
);

INVx11_ASAP7_75t_L g41 ( 
.A(n_30),
.Y(n_41)
);

INVx4_ASAP7_75t_L g68 ( 
.A(n_41),
.Y(n_68)
);

BUFx3_ASAP7_75t_L g42 ( 
.A(n_32),
.Y(n_42)
);

BUFx3_ASAP7_75t_L g75 ( 
.A(n_42),
.Y(n_75)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_22),
.Y(n_43)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_43),
.Y(n_89)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_23),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g92 ( 
.A(n_44),
.Y(n_92)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_23),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g93 ( 
.A(n_45),
.Y(n_93)
);

INVx6_ASAP7_75t_SL g46 ( 
.A(n_26),
.Y(n_46)
);

CKINVDCx20_ASAP7_75t_R g85 ( 
.A(n_46),
.Y(n_85)
);

BUFx3_ASAP7_75t_L g47 ( 
.A(n_32),
.Y(n_47)
);

INVx5_ASAP7_75t_L g73 ( 
.A(n_47),
.Y(n_73)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_23),
.Y(n_48)
);

INVx8_ASAP7_75t_L g70 ( 
.A(n_48),
.Y(n_70)
);

INVx11_ASAP7_75t_L g49 ( 
.A(n_30),
.Y(n_49)
);

INVx4_ASAP7_75t_L g78 ( 
.A(n_49),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_L g50 ( 
.A(n_20),
.B(n_0),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_50),
.B(n_51),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_SL g51 ( 
.A(n_20),
.B(n_12),
.Y(n_51)
);

INVx5_ASAP7_75t_L g52 ( 
.A(n_32),
.Y(n_52)
);

INVx4_ASAP7_75t_L g88 ( 
.A(n_52),
.Y(n_88)
);

BUFx4f_ASAP7_75t_SL g53 ( 
.A(n_26),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_53),
.B(n_54),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_SL g54 ( 
.A(n_31),
.B(n_0),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_SL g55 ( 
.A(n_29),
.B(n_31),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_SL g69 ( 
.A(n_55),
.B(n_21),
.Y(n_69)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_27),
.Y(n_56)
);

INVx3_ASAP7_75t_L g77 ( 
.A(n_56),
.Y(n_77)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_28),
.Y(n_57)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_57),
.Y(n_95)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_27),
.Y(n_58)
);

INVx3_ASAP7_75t_L g91 ( 
.A(n_58),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_29),
.B(n_11),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_59),
.B(n_62),
.Y(n_67)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_27),
.Y(n_60)
);

INVx4_ASAP7_75t_L g100 ( 
.A(n_60),
.Y(n_100)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_38),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_L g86 ( 
.A(n_61),
.B(n_65),
.Y(n_86)
);

INVx4_ASAP7_75t_L g62 ( 
.A(n_17),
.Y(n_62)
);

INVx11_ASAP7_75t_L g63 ( 
.A(n_26),
.Y(n_63)
);

AOI22xp33_ASAP7_75t_SL g66 ( 
.A1(n_63),
.A2(n_64),
.B1(n_34),
.B2(n_38),
.Y(n_66)
);

INVx11_ASAP7_75t_L g64 ( 
.A(n_25),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_L g65 ( 
.A(n_28),
.B(n_2),
.Y(n_65)
);

INVxp67_ASAP7_75t_L g103 ( 
.A(n_66),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_SL g108 ( 
.A(n_69),
.B(n_98),
.Y(n_108)
);

AOI22xp33_ASAP7_75t_SL g71 ( 
.A1(n_42),
.A2(n_34),
.B1(n_17),
.B2(n_37),
.Y(n_71)
);

AOI22xp33_ASAP7_75t_SL g107 ( 
.A1(n_71),
.A2(n_74),
.B1(n_87),
.B2(n_63),
.Y(n_107)
);

AND2x4_ASAP7_75t_L g72 ( 
.A(n_65),
.B(n_57),
.Y(n_72)
);

INVx1_ASAP7_75t_SL g102 ( 
.A(n_72),
.Y(n_102)
);

AOI22xp33_ASAP7_75t_SL g74 ( 
.A1(n_47),
.A2(n_35),
.B1(n_22),
.B2(n_37),
.Y(n_74)
);

AOI22xp33_ASAP7_75t_L g76 ( 
.A1(n_44),
.A2(n_19),
.B1(n_36),
.B2(n_39),
.Y(n_76)
);

OAI22xp5_ASAP7_75t_L g111 ( 
.A1(n_76),
.A2(n_96),
.B1(n_40),
.B2(n_41),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_55),
.B(n_50),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_79),
.B(n_81),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_51),
.B(n_21),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_43),
.B(n_18),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g116 ( 
.A(n_82),
.B(n_90),
.Y(n_116)
);

MAJIxp5_ASAP7_75t_L g84 ( 
.A(n_62),
.B(n_38),
.C(n_39),
.Y(n_84)
);

MAJIxp5_ASAP7_75t_L g109 ( 
.A(n_84),
.B(n_72),
.C(n_85),
.Y(n_109)
);

AOI22xp33_ASAP7_75t_SL g87 ( 
.A1(n_52),
.A2(n_35),
.B1(n_36),
.B2(n_19),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_53),
.B(n_18),
.Y(n_90)
);

HAxp5_ASAP7_75t_SL g94 ( 
.A(n_46),
.B(n_33),
.CON(n_94),
.SN(n_94)
);

NOR2xp33_ASAP7_75t_SL g118 ( 
.A(n_94),
.B(n_25),
.Y(n_118)
);

AOI22xp5_ASAP7_75t_L g96 ( 
.A1(n_56),
.A2(n_24),
.B1(n_33),
.B2(n_25),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_53),
.B(n_24),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_97),
.B(n_60),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_SL g98 ( 
.A(n_61),
.B(n_11),
.Y(n_98)
);

XOR2xp5_ASAP7_75t_L g101 ( 
.A(n_72),
.B(n_33),
.Y(n_101)
);

XNOR2xp5_ASAP7_75t_L g142 ( 
.A(n_101),
.B(n_93),
.Y(n_142)
);

INVx2_ASAP7_75t_L g104 ( 
.A(n_89),
.Y(n_104)
);

INVx2_ASAP7_75t_L g145 ( 
.A(n_104),
.Y(n_145)
);

AOI22xp5_ASAP7_75t_L g106 ( 
.A1(n_72),
.A2(n_56),
.B1(n_58),
.B2(n_60),
.Y(n_106)
);

OAI22xp5_ASAP7_75t_SL g131 ( 
.A1(n_106),
.A2(n_124),
.B1(n_92),
.B2(n_93),
.Y(n_131)
);

AO21x1_ASAP7_75t_L g151 ( 
.A1(n_107),
.A2(n_118),
.B(n_122),
.Y(n_151)
);

AND2x2_ASAP7_75t_L g135 ( 
.A(n_109),
.B(n_111),
.Y(n_135)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_89),
.Y(n_110)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_110),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_L g112 ( 
.A(n_86),
.B(n_48),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_L g133 ( 
.A(n_112),
.B(n_113),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_L g113 ( 
.A(n_86),
.B(n_48),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_SL g114 ( 
.A(n_80),
.B(n_58),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_SL g147 ( 
.A(n_114),
.B(n_121),
.Y(n_147)
);

INVx4_ASAP7_75t_L g115 ( 
.A(n_99),
.Y(n_115)
);

INVx1_ASAP7_75t_SL g137 ( 
.A(n_115),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_L g134 ( 
.A(n_117),
.B(n_127),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_L g119 ( 
.A(n_95),
.B(n_44),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_L g138 ( 
.A(n_119),
.B(n_93),
.Y(n_138)
);

INVx1_ASAP7_75t_SL g120 ( 
.A(n_68),
.Y(n_120)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_120),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_SL g121 ( 
.A(n_80),
.B(n_45),
.Y(n_121)
);

OAI32xp33_ASAP7_75t_L g122 ( 
.A1(n_83),
.A2(n_64),
.A3(n_33),
.B1(n_25),
.B2(n_49),
.Y(n_122)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_95),
.Y(n_123)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_123),
.Y(n_140)
);

OAI22xp5_ASAP7_75t_SL g124 ( 
.A1(n_96),
.A2(n_45),
.B1(n_77),
.B2(n_91),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_SL g125 ( 
.A(n_83),
.B(n_2),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_SL g136 ( 
.A(n_125),
.B(n_126),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_L g126 ( 
.A(n_69),
.B(n_3),
.Y(n_126)
);

CKINVDCx20_ASAP7_75t_R g127 ( 
.A(n_85),
.Y(n_127)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_77),
.Y(n_128)
);

INVx2_ASAP7_75t_L g155 ( 
.A(n_128),
.Y(n_155)
);

OAI22xp5_ASAP7_75t_L g129 ( 
.A1(n_84),
.A2(n_25),
.B1(n_33),
.B2(n_6),
.Y(n_129)
);

AOI22xp33_ASAP7_75t_L g149 ( 
.A1(n_129),
.A2(n_92),
.B1(n_100),
.B2(n_99),
.Y(n_149)
);

NOR2xp33_ASAP7_75t_L g130 ( 
.A(n_67),
.B(n_8),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_L g150 ( 
.A(n_130),
.B(n_3),
.Y(n_150)
);

AOI22xp5_ASAP7_75t_L g177 ( 
.A1(n_131),
.A2(n_139),
.B1(n_149),
.B2(n_7),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_L g163 ( 
.A(n_138),
.B(n_143),
.Y(n_163)
);

OAI22xp33_ASAP7_75t_SL g139 ( 
.A1(n_102),
.A2(n_94),
.B1(n_88),
.B2(n_75),
.Y(n_139)
);

AOI32xp33_ASAP7_75t_L g141 ( 
.A1(n_112),
.A2(n_98),
.A3(n_88),
.B1(n_78),
.B2(n_68),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_L g162 ( 
.A(n_141),
.B(n_144),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_SL g169 ( 
.A(n_142),
.B(n_148),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_L g143 ( 
.A(n_113),
.B(n_91),
.Y(n_143)
);

AOI32xp33_ASAP7_75t_L g144 ( 
.A1(n_105),
.A2(n_78),
.A3(n_100),
.B1(n_73),
.B2(n_75),
.Y(n_144)
);

AOI21xp33_ASAP7_75t_L g146 ( 
.A1(n_125),
.A2(n_3),
.B(n_5),
.Y(n_146)
);

AOI21xp33_ASAP7_75t_L g164 ( 
.A1(n_146),
.A2(n_129),
.B(n_114),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_L g148 ( 
.A(n_121),
.B(n_73),
.Y(n_148)
);

NOR2xp33_ASAP7_75t_SL g160 ( 
.A(n_150),
.B(n_108),
.Y(n_160)
);

OAI32xp33_ASAP7_75t_L g153 ( 
.A1(n_102),
.A2(n_70),
.A3(n_92),
.B1(n_7),
.B2(n_5),
.Y(n_153)
);

OAI21xp5_ASAP7_75t_L g168 ( 
.A1(n_153),
.A2(n_106),
.B(n_122),
.Y(n_168)
);

NOR2xp33_ASAP7_75t_L g154 ( 
.A(n_116),
.B(n_6),
.Y(n_154)
);

CKINVDCx14_ASAP7_75t_R g159 ( 
.A(n_154),
.Y(n_159)
);

CKINVDCx20_ASAP7_75t_R g156 ( 
.A(n_134),
.Y(n_156)
);

NOR2xp33_ASAP7_75t_L g178 ( 
.A(n_156),
.B(n_160),
.Y(n_178)
);

INVxp67_ASAP7_75t_SL g157 ( 
.A(n_152),
.Y(n_157)
);

INVxp67_ASAP7_75t_L g185 ( 
.A(n_157),
.Y(n_185)
);

AOI21xp5_ASAP7_75t_L g158 ( 
.A1(n_135),
.A2(n_109),
.B(n_103),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_L g181 ( 
.A(n_158),
.B(n_161),
.Y(n_181)
);

AOI21xp5_ASAP7_75t_L g161 ( 
.A1(n_135),
.A2(n_103),
.B(n_118),
.Y(n_161)
);

NOR2xp33_ASAP7_75t_L g183 ( 
.A(n_164),
.B(n_165),
.Y(n_183)
);

CKINVDCx20_ASAP7_75t_R g165 ( 
.A(n_143),
.Y(n_165)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_132),
.Y(n_166)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_166),
.Y(n_184)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_132),
.Y(n_167)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_167),
.Y(n_186)
);

OAI22xp5_ASAP7_75t_L g191 ( 
.A1(n_168),
.A2(n_177),
.B1(n_137),
.B2(n_145),
.Y(n_191)
);

NOR3xp33_ASAP7_75t_SL g170 ( 
.A(n_136),
.B(n_127),
.C(n_110),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_SL g182 ( 
.A(n_170),
.B(n_171),
.Y(n_182)
);

NOR2xp33_ASAP7_75t_L g171 ( 
.A(n_147),
.B(n_104),
.Y(n_171)
);

A2O1A1O1Ixp25_ASAP7_75t_L g172 ( 
.A1(n_133),
.A2(n_101),
.B(n_119),
.C(n_123),
.D(n_128),
.Y(n_172)
);

NOR2xp33_ASAP7_75t_L g188 ( 
.A(n_172),
.B(n_175),
.Y(n_188)
);

OAI21xp5_ASAP7_75t_L g173 ( 
.A1(n_135),
.A2(n_111),
.B(n_120),
.Y(n_173)
);

XOR2xp5_ASAP7_75t_L g189 ( 
.A(n_173),
.B(n_131),
.Y(n_189)
);

NAND2x1_ASAP7_75t_SL g174 ( 
.A(n_151),
.B(n_115),
.Y(n_174)
);

CKINVDCx20_ASAP7_75t_R g193 ( 
.A(n_174),
.Y(n_193)
);

NOR2xp33_ASAP7_75t_L g175 ( 
.A(n_140),
.B(n_70),
.Y(n_175)
);

OAI21xp5_ASAP7_75t_SL g176 ( 
.A1(n_151),
.A2(n_124),
.B(n_6),
.Y(n_176)
);

XOR2xp5_ASAP7_75t_L g195 ( 
.A(n_176),
.B(n_155),
.Y(n_195)
);

MAJIxp5_ASAP7_75t_L g179 ( 
.A(n_158),
.B(n_142),
.C(n_133),
.Y(n_179)
);

XOR2xp5_ASAP7_75t_L g208 ( 
.A(n_179),
.B(n_189),
.Y(n_208)
);

AOI22xp5_ASAP7_75t_L g180 ( 
.A1(n_168),
.A2(n_173),
.B1(n_165),
.B2(n_162),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_L g198 ( 
.A(n_180),
.B(n_187),
.Y(n_198)
);

OAI22xp5_ASAP7_75t_SL g187 ( 
.A1(n_162),
.A2(n_148),
.B1(n_138),
.B2(n_153),
.Y(n_187)
);

NOR2xp33_ASAP7_75t_L g190 ( 
.A(n_156),
.B(n_152),
.Y(n_190)
);

NOR2xp33_ASAP7_75t_SL g209 ( 
.A(n_190),
.B(n_171),
.Y(n_209)
);

AOI22xp5_ASAP7_75t_SL g202 ( 
.A1(n_191),
.A2(n_194),
.B1(n_166),
.B2(n_167),
.Y(n_202)
);

INVx5_ASAP7_75t_L g192 ( 
.A(n_170),
.Y(n_192)
);

NOR2xp33_ASAP7_75t_L g197 ( 
.A(n_192),
.B(n_195),
.Y(n_197)
);

OAI22xp5_ASAP7_75t_L g194 ( 
.A1(n_163),
.A2(n_145),
.B1(n_155),
.B2(n_137),
.Y(n_194)
);

CKINVDCx16_ASAP7_75t_R g196 ( 
.A(n_194),
.Y(n_196)
);

NAND2xp5_ASAP7_75t_L g212 ( 
.A(n_196),
.B(n_200),
.Y(n_212)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_184),
.Y(n_199)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_199),
.Y(n_214)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_184),
.Y(n_200)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_186),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_SL g210 ( 
.A(n_201),
.B(n_202),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_L g203 ( 
.A(n_186),
.B(n_163),
.Y(n_203)
);

CKINVDCx14_ASAP7_75t_R g215 ( 
.A(n_203),
.Y(n_215)
);

CKINVDCx20_ASAP7_75t_R g204 ( 
.A(n_185),
.Y(n_204)
);

NAND2xp5_ASAP7_75t_SL g211 ( 
.A(n_204),
.B(n_205),
.Y(n_211)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_185),
.Y(n_205)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_189),
.Y(n_206)
);

XNOR2xp5_ASAP7_75t_L g219 ( 
.A(n_206),
.B(n_209),
.Y(n_219)
);

NOR2xp33_ASAP7_75t_L g207 ( 
.A(n_182),
.B(n_160),
.Y(n_207)
);

AOI322xp5_ASAP7_75t_L g216 ( 
.A1(n_207),
.A2(n_178),
.A3(n_183),
.B1(n_188),
.B2(n_192),
.C1(n_169),
.C2(n_159),
.Y(n_216)
);

MAJIxp5_ASAP7_75t_L g213 ( 
.A(n_208),
.B(n_179),
.C(n_181),
.Y(n_213)
);

MAJIxp5_ASAP7_75t_L g220 ( 
.A(n_213),
.B(n_217),
.C(n_218),
.Y(n_220)
);

NOR2xp33_ASAP7_75t_L g222 ( 
.A(n_216),
.B(n_198),
.Y(n_222)
);

MAJIxp5_ASAP7_75t_L g217 ( 
.A(n_208),
.B(n_181),
.C(n_169),
.Y(n_217)
);

MAJIxp5_ASAP7_75t_L g218 ( 
.A(n_206),
.B(n_180),
.C(n_161),
.Y(n_218)
);

NAND2xp5_ASAP7_75t_L g221 ( 
.A(n_211),
.B(n_204),
.Y(n_221)
);

NOR2xp33_ASAP7_75t_L g229 ( 
.A(n_221),
.B(n_223),
.Y(n_229)
);

AOI21xp5_ASAP7_75t_SL g232 ( 
.A1(n_222),
.A2(n_224),
.B(n_219),
.Y(n_232)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_214),
.Y(n_223)
);

OAI21xp5_ASAP7_75t_SL g224 ( 
.A1(n_210),
.A2(n_197),
.B(n_198),
.Y(n_224)
);

AOI22xp5_ASAP7_75t_L g225 ( 
.A1(n_212),
.A2(n_193),
.B1(n_195),
.B2(n_203),
.Y(n_225)
);

NOR2xp33_ASAP7_75t_L g231 ( 
.A(n_225),
.B(n_227),
.Y(n_231)
);

AOI21xp5_ASAP7_75t_L g226 ( 
.A1(n_218),
.A2(n_193),
.B(n_176),
.Y(n_226)
);

OAI21xp33_ASAP7_75t_L g228 ( 
.A1(n_226),
.A2(n_217),
.B(n_213),
.Y(n_228)
);

NOR2xp33_ASAP7_75t_L g227 ( 
.A(n_219),
.B(n_205),
.Y(n_227)
);

NAND2xp5_ASAP7_75t_L g234 ( 
.A(n_228),
.B(n_233),
.Y(n_234)
);

AOI22xp5_ASAP7_75t_SL g230 ( 
.A1(n_226),
.A2(n_187),
.B1(n_215),
.B2(n_174),
.Y(n_230)
);

MAJIxp5_ASAP7_75t_L g235 ( 
.A(n_230),
.B(n_232),
.C(n_225),
.Y(n_235)
);

NOR2xp33_ASAP7_75t_L g233 ( 
.A(n_220),
.B(n_175),
.Y(n_233)
);

AOI21xp5_ASAP7_75t_SL g240 ( 
.A1(n_235),
.A2(n_237),
.B(n_172),
.Y(n_240)
);

MAJIxp5_ASAP7_75t_L g236 ( 
.A(n_231),
.B(n_220),
.C(n_202),
.Y(n_236)
);

MAJIxp5_ASAP7_75t_L g239 ( 
.A(n_236),
.B(n_174),
.C(n_201),
.Y(n_239)
);

NAND2xp5_ASAP7_75t_L g237 ( 
.A(n_229),
.B(n_199),
.Y(n_237)
);

OAI21x1_ASAP7_75t_SL g238 ( 
.A1(n_234),
.A2(n_228),
.B(n_200),
.Y(n_238)
);

INVxp67_ASAP7_75t_L g241 ( 
.A(n_238),
.Y(n_241)
);

INVxp67_ASAP7_75t_L g242 ( 
.A(n_239),
.Y(n_242)
);

OAI21xp5_ASAP7_75t_SL g243 ( 
.A1(n_241),
.A2(n_240),
.B(n_177),
.Y(n_243)
);

XNOR2xp5_ASAP7_75t_L g244 ( 
.A(n_243),
.B(n_242),
.Y(n_244)
);


endmodule