module fake_ariane_3223_n_1932 (n_83, n_8, n_56, n_60, n_170, n_190, n_160, n_64, n_179, n_180, n_119, n_124, n_167, n_90, n_195, n_38, n_47, n_110, n_153, n_18, n_197, n_86, n_75, n_89, n_67, n_176, n_149, n_34, n_158, n_172, n_69, n_95, n_175, n_92, n_143, n_183, n_150, n_98, n_74, n_113, n_114, n_33, n_19, n_40, n_181, n_152, n_120, n_169, n_106, n_12, n_53, n_173, n_111, n_21, n_115, n_133, n_66, n_71, n_24, n_7, n_109, n_96, n_156, n_49, n_20, n_174, n_100, n_17, n_50, n_187, n_132, n_62, n_147, n_200, n_51, n_166, n_76, n_103, n_79, n_26, n_3, n_46, n_0, n_84, n_36, n_199, n_91, n_159, n_107, n_189, n_72, n_105, n_128, n_44, n_30, n_82, n_178, n_31, n_42, n_57, n_131, n_201, n_70, n_10, n_117, n_139, n_165, n_85, n_130, n_144, n_6, n_48, n_94, n_101, n_4, n_134, n_188, n_185, n_2, n_32, n_37, n_58, n_65, n_123, n_9, n_138, n_112, n_45, n_162, n_11, n_129, n_126, n_137, n_122, n_198, n_148, n_164, n_52, n_157, n_184, n_177, n_135, n_73, n_77, n_171, n_15, n_118, n_93, n_121, n_23, n_61, n_108, n_102, n_182, n_196, n_125, n_22, n_168, n_43, n_1, n_81, n_87, n_13, n_27, n_29, n_41, n_140, n_55, n_191, n_151, n_136, n_192, n_28, n_80, n_146, n_194, n_97, n_154, n_142, n_161, n_14, n_163, n_88, n_186, n_141, n_68, n_116, n_104, n_202, n_145, n_78, n_193, n_39, n_59, n_63, n_99, n_16, n_5, n_155, n_127, n_35, n_54, n_25, n_1932);

input n_83;
input n_8;
input n_56;
input n_60;
input n_170;
input n_190;
input n_160;
input n_64;
input n_179;
input n_180;
input n_119;
input n_124;
input n_167;
input n_90;
input n_195;
input n_38;
input n_47;
input n_110;
input n_153;
input n_18;
input n_197;
input n_86;
input n_75;
input n_89;
input n_67;
input n_176;
input n_149;
input n_34;
input n_158;
input n_172;
input n_69;
input n_95;
input n_175;
input n_92;
input n_143;
input n_183;
input n_150;
input n_98;
input n_74;
input n_113;
input n_114;
input n_33;
input n_19;
input n_40;
input n_181;
input n_152;
input n_120;
input n_169;
input n_106;
input n_12;
input n_53;
input n_173;
input n_111;
input n_21;
input n_115;
input n_133;
input n_66;
input n_71;
input n_24;
input n_7;
input n_109;
input n_96;
input n_156;
input n_49;
input n_20;
input n_174;
input n_100;
input n_17;
input n_50;
input n_187;
input n_132;
input n_62;
input n_147;
input n_200;
input n_51;
input n_166;
input n_76;
input n_103;
input n_79;
input n_26;
input n_3;
input n_46;
input n_0;
input n_84;
input n_36;
input n_199;
input n_91;
input n_159;
input n_107;
input n_189;
input n_72;
input n_105;
input n_128;
input n_44;
input n_30;
input n_82;
input n_178;
input n_31;
input n_42;
input n_57;
input n_131;
input n_201;
input n_70;
input n_10;
input n_117;
input n_139;
input n_165;
input n_85;
input n_130;
input n_144;
input n_6;
input n_48;
input n_94;
input n_101;
input n_4;
input n_134;
input n_188;
input n_185;
input n_2;
input n_32;
input n_37;
input n_58;
input n_65;
input n_123;
input n_9;
input n_138;
input n_112;
input n_45;
input n_162;
input n_11;
input n_129;
input n_126;
input n_137;
input n_122;
input n_198;
input n_148;
input n_164;
input n_52;
input n_157;
input n_184;
input n_177;
input n_135;
input n_73;
input n_77;
input n_171;
input n_15;
input n_118;
input n_93;
input n_121;
input n_23;
input n_61;
input n_108;
input n_102;
input n_182;
input n_196;
input n_125;
input n_22;
input n_168;
input n_43;
input n_1;
input n_81;
input n_87;
input n_13;
input n_27;
input n_29;
input n_41;
input n_140;
input n_55;
input n_191;
input n_151;
input n_136;
input n_192;
input n_28;
input n_80;
input n_146;
input n_194;
input n_97;
input n_154;
input n_142;
input n_161;
input n_14;
input n_163;
input n_88;
input n_186;
input n_141;
input n_68;
input n_116;
input n_104;
input n_202;
input n_145;
input n_78;
input n_193;
input n_39;
input n_59;
input n_63;
input n_99;
input n_16;
input n_5;
input n_155;
input n_127;
input n_35;
input n_54;
input n_25;

output n_1932;

wire n_913;
wire n_1681;
wire n_1486;
wire n_1507;
wire n_589;
wire n_1174;
wire n_1469;
wire n_691;
wire n_1353;
wire n_1355;
wire n_423;
wire n_1383;
wire n_603;
wire n_373;
wire n_1250;
wire n_1169;
wire n_789;
wire n_850;
wire n_1916;
wire n_610;
wire n_245;
wire n_1713;
wire n_319;
wire n_1436;
wire n_690;
wire n_416;
wire n_1109;
wire n_1430;
wire n_525;
wire n_1463;
wire n_1238;
wire n_1515;
wire n_817;
wire n_1837;
wire n_924;
wire n_781;
wire n_1566;
wire n_717;
wire n_952;
wire n_864;
wire n_1096;
wire n_1379;
wire n_1706;
wire n_524;
wire n_1214;
wire n_634;
wire n_1839;
wire n_1246;
wire n_1138;
wire n_214;
wire n_1853;
wire n_764;
wire n_1503;
wire n_462;
wire n_1196;
wire n_1181;
wire n_410;
wire n_1187;
wire n_1131;
wire n_1225;
wire n_737;
wire n_1298;
wire n_1745;
wire n_1366;
wire n_232;
wire n_568;
wire n_1088;
wire n_1424;
wire n_766;
wire n_1835;
wire n_1457;
wire n_377;
wire n_1682;
wire n_1836;
wire n_520;
wire n_870;
wire n_1453;
wire n_279;
wire n_958;
wire n_945;
wire n_813;
wire n_419;
wire n_270;
wire n_338;
wire n_995;
wire n_285;
wire n_1909;
wire n_1184;
wire n_1535;
wire n_500;
wire n_665;
wire n_754;
wire n_903;
wire n_871;
wire n_1073;
wire n_239;
wire n_402;
wire n_1277;
wire n_1746;
wire n_829;
wire n_1761;
wire n_1062;
wire n_339;
wire n_738;
wire n_1690;
wire n_672;
wire n_740;
wire n_1283;
wire n_1736;
wire n_1018;
wire n_259;
wire n_953;
wire n_1364;
wire n_1888;
wire n_1224;
wire n_1425;
wire n_625;
wire n_557;
wire n_1107;
wire n_1688;
wire n_989;
wire n_242;
wire n_645;
wire n_331;
wire n_559;
wire n_495;
wire n_267;
wire n_350;
wire n_381;
wire n_795;
wire n_721;
wire n_1084;
wire n_1718;
wire n_1276;
wire n_1428;
wire n_1284;
wire n_1241;
wire n_821;
wire n_561;
wire n_770;
wire n_1514;
wire n_1528;
wire n_507;
wire n_486;
wire n_901;
wire n_569;
wire n_1145;
wire n_971;
wire n_787;
wire n_1650;
wire n_1519;
wire n_1195;
wire n_1522;
wire n_518;
wire n_1207;
wire n_222;
wire n_786;
wire n_1404;
wire n_868;
wire n_1847;
wire n_1542;
wire n_1314;
wire n_1512;
wire n_1539;
wire n_884;
wire n_1851;
wire n_1415;
wire n_1034;
wire n_1652;
wire n_1676;
wire n_1085;
wire n_277;
wire n_1636;
wire n_432;
wire n_293;
wire n_823;
wire n_1900;
wire n_620;
wire n_1074;
wire n_859;
wire n_1765;
wire n_1889;
wire n_587;
wire n_693;
wire n_863;
wire n_303;
wire n_1254;
wire n_929;
wire n_206;
wire n_352;
wire n_899;
wire n_1703;
wire n_611;
wire n_1295;
wire n_1850;
wire n_365;
wire n_238;
wire n_1013;
wire n_1495;
wire n_1637;
wire n_334;
wire n_661;
wire n_1751;
wire n_300;
wire n_533;
wire n_1917;
wire n_1924;
wire n_438;
wire n_1560;
wire n_1654;
wire n_1548;
wire n_1811;
wire n_440;
wire n_273;
wire n_1396;
wire n_1230;
wire n_612;
wire n_333;
wire n_1840;
wire n_376;
wire n_512;
wire n_1597;
wire n_1771;
wire n_1544;
wire n_579;
wire n_844;
wire n_1012;
wire n_1267;
wire n_1354;
wire n_1790;
wire n_1213;
wire n_237;
wire n_780;
wire n_1918;
wire n_1021;
wire n_1443;
wire n_491;
wire n_1465;
wire n_1595;
wire n_1142;
wire n_1140;
wire n_705;
wire n_570;
wire n_260;
wire n_942;
wire n_1437;
wire n_1378;
wire n_461;
wire n_1121;
wire n_1416;
wire n_209;
wire n_490;
wire n_1461;
wire n_1391;
wire n_225;
wire n_1599;
wire n_1876;
wire n_1006;
wire n_1830;
wire n_575;
wire n_546;
wire n_503;
wire n_1112;
wire n_700;
wire n_1159;
wire n_772;
wire n_1216;
wire n_1245;
wire n_1669;
wire n_1675;
wire n_676;
wire n_1838;
wire n_1594;
wire n_680;
wire n_287;
wire n_1716;
wire n_302;
wire n_1872;
wire n_380;
wire n_1585;
wire n_1432;
wire n_249;
wire n_1108;
wire n_355;
wire n_212;
wire n_444;
wire n_851;
wire n_1590;
wire n_1351;
wire n_1274;
wire n_257;
wire n_652;
wire n_1819;
wire n_475;
wire n_947;
wire n_930;
wire n_1260;
wire n_1179;
wire n_468;
wire n_696;
wire n_1442;
wire n_482;
wire n_798;
wire n_577;
wire n_1833;
wire n_407;
wire n_1691;
wire n_916;
wire n_1386;
wire n_912;
wire n_1884;
wire n_460;
wire n_1555;
wire n_1842;
wire n_366;
wire n_762;
wire n_1253;
wire n_1468;
wire n_1661;
wire n_555;
wire n_804;
wire n_1656;
wire n_1382;
wire n_992;
wire n_966;
wire n_955;
wire n_1182;
wire n_794;
wire n_1692;
wire n_1562;
wire n_514;
wire n_418;
wire n_1376;
wire n_513;
wire n_288;
wire n_1292;
wire n_1178;
wire n_1435;
wire n_1750;
wire n_1026;
wire n_1506;
wire n_1610;
wire n_306;
wire n_203;
wire n_436;
wire n_324;
wire n_669;
wire n_931;
wire n_1491;
wire n_619;
wire n_437;
wire n_337;
wire n_274;
wire n_967;
wire n_1083;
wire n_1418;
wire n_746;
wire n_1357;
wire n_292;
wire n_1079;
wire n_1787;
wire n_1389;
wire n_615;
wire n_1139;
wire n_517;
wire n_1312;
wire n_1717;
wire n_1812;
wire n_824;
wire n_428;
wire n_892;
wire n_1880;
wire n_959;
wire n_1399;
wire n_1101;
wire n_1567;
wire n_1343;
wire n_563;
wire n_1855;
wire n_990;
wire n_1623;
wire n_1903;
wire n_867;
wire n_1226;
wire n_944;
wire n_749;
wire n_1780;
wire n_1920;
wire n_815;
wire n_542;
wire n_1340;
wire n_470;
wire n_1240;
wire n_1087;
wire n_632;
wire n_477;
wire n_650;
wire n_425;
wire n_1433;
wire n_1911;
wire n_1825;
wire n_1908;
wire n_1155;
wire n_1071;
wire n_712;
wire n_976;
wire n_909;
wire n_1392;
wire n_767;
wire n_1832;
wire n_1841;
wire n_1680;
wire n_964;
wire n_1627;
wire n_382;
wire n_489;
wire n_251;
wire n_974;
wire n_506;
wire n_1731;
wire n_799;
wire n_1147;
wire n_397;
wire n_471;
wire n_351;
wire n_965;
wire n_1914;
wire n_934;
wire n_1447;
wire n_1220;
wire n_356;
wire n_698;
wire n_1674;
wire n_307;
wire n_1209;
wire n_1020;
wire n_1563;
wire n_646;
wire n_1633;
wire n_404;
wire n_1913;
wire n_1058;
wire n_347;
wire n_1042;
wire n_1234;
wire n_479;
wire n_1578;
wire n_1455;
wire n_299;
wire n_836;
wire n_1279;
wire n_564;
wire n_205;
wire n_1029;
wire n_1247;
wire n_760;
wire n_522;
wire n_1568;
wire n_1483;
wire n_1363;
wire n_367;
wire n_1111;
wire n_970;
wire n_1689;
wire n_713;
wire n_1255;
wire n_1646;
wire n_598;
wire n_345;
wire n_1237;
wire n_927;
wire n_261;
wire n_1095;
wire n_1728;
wire n_370;
wire n_706;
wire n_286;
wire n_1401;
wire n_1419;
wire n_1531;
wire n_776;
wire n_424;
wire n_1651;
wire n_1387;
wire n_466;
wire n_1263;
wire n_346;
wire n_1817;
wire n_552;
wire n_348;
wire n_670;
wire n_1826;
wire n_379;
wire n_264;
wire n_441;
wire n_1032;
wire n_1217;
wire n_1496;
wire n_637;
wire n_1592;
wire n_327;
wire n_1259;
wire n_1177;
wire n_1231;
wire n_980;
wire n_1618;
wire n_1869;
wire n_1743;
wire n_905;
wire n_207;
wire n_720;
wire n_926;
wire n_1802;
wire n_1163;
wire n_1795;
wire n_1384;
wire n_1868;
wire n_1501;
wire n_1173;
wire n_1068;
wire n_1198;
wire n_1570;
wire n_487;
wire n_1518;
wire n_1456;
wire n_1879;
wire n_1886;
wire n_1648;
wire n_1413;
wire n_855;
wire n_808;
wire n_1365;
wire n_553;
wire n_1439;
wire n_814;
wire n_578;
wire n_1665;
wire n_1287;
wire n_405;
wire n_1611;
wire n_320;
wire n_1414;
wire n_1134;
wire n_1484;
wire n_1901;
wire n_647;
wire n_1423;
wire n_600;
wire n_481;
wire n_1053;
wire n_1609;
wire n_1906;
wire n_529;
wire n_1899;
wire n_502;
wire n_218;
wire n_1467;
wire n_247;
wire n_1828;
wire n_1798;
wire n_1304;
wire n_1608;
wire n_1744;
wire n_1105;
wire n_547;
wire n_439;
wire n_677;
wire n_604;
wire n_478;
wire n_703;
wire n_1349;
wire n_1709;
wire n_1061;
wire n_326;
wire n_681;
wire n_227;
wire n_874;
wire n_1278;
wire n_707;
wire n_983;
wire n_590;
wire n_699;
wire n_727;
wire n_301;
wire n_1726;
wire n_545;
wire n_1015;
wire n_1377;
wire n_1162;
wire n_536;
wire n_1614;
wire n_325;
wire n_1740;
wire n_1602;
wire n_688;
wire n_636;
wire n_427;
wire n_1098;
wire n_1490;
wire n_442;
wire n_777;
wire n_1553;
wire n_1080;
wire n_920;
wire n_1760;
wire n_1086;
wire n_1092;
wire n_986;
wire n_1104;
wire n_729;
wire n_887;
wire n_1122;
wire n_1205;
wire n_1408;
wire n_1693;
wire n_1132;
wire n_390;
wire n_1156;
wire n_501;
wire n_314;
wire n_1823;
wire n_1120;
wire n_1202;
wire n_627;
wire n_1188;
wire n_1498;
wire n_1371;
wire n_233;
wire n_957;
wire n_388;
wire n_1402;
wire n_1242;
wire n_1607;
wire n_1489;
wire n_1218;
wire n_221;
wire n_321;
wire n_1586;
wire n_861;
wire n_1543;
wire n_1431;
wire n_877;
wire n_1119;
wire n_1863;
wire n_1763;
wire n_1666;
wire n_1500;
wire n_616;
wire n_1055;
wire n_1395;
wire n_1346;
wire n_1189;
wire n_1089;
wire n_281;
wire n_1859;
wire n_262;
wire n_1502;
wire n_1523;
wire n_1478;
wire n_1883;
wire n_735;
wire n_297;
wire n_1005;
wire n_527;
wire n_1294;
wire n_1667;
wire n_845;
wire n_888;
wire n_1649;
wire n_1677;
wire n_1927;
wire n_1297;
wire n_551;
wire n_417;
wire n_1708;
wire n_343;
wire n_1222;
wire n_1844;
wire n_582;
wire n_755;
wire n_1097;
wire n_1219;
wire n_1711;
wire n_710;
wire n_1919;
wire n_534;
wire n_1791;
wire n_1894;
wire n_1460;
wire n_1239;
wire n_278;
wire n_560;
wire n_890;
wire n_842;
wire n_1898;
wire n_451;
wire n_745;
wire n_1741;
wire n_1572;
wire n_1907;
wire n_1793;
wire n_742;
wire n_1081;
wire n_1373;
wire n_1388;
wire n_1266;
wire n_1540;
wire n_1719;
wire n_769;
wire n_1797;
wire n_1753;
wire n_1372;
wire n_476;
wire n_832;
wire n_535;
wire n_744;
wire n_1895;
wire n_982;
wire n_1800;
wire n_915;
wire n_215;
wire n_1075;
wire n_454;
wire n_298;
wire n_1331;
wire n_1890;
wire n_1529;
wire n_1227;
wire n_655;
wire n_1734;
wire n_1860;
wire n_403;
wire n_1007;
wire n_1580;
wire n_1319;
wire n_657;
wire n_837;
wire n_812;
wire n_606;
wire n_951;
wire n_862;
wire n_1700;
wire n_659;
wire n_1332;
wire n_509;
wire n_1854;
wire n_666;
wire n_1747;
wire n_430;
wire n_1206;
wire n_1729;
wire n_722;
wire n_1508;
wire n_1532;
wire n_1171;
wire n_1030;
wire n_785;
wire n_1309;
wire n_999;
wire n_1766;
wire n_1338;
wire n_1342;
wire n_456;
wire n_1867;
wire n_852;
wire n_1394;
wire n_704;
wire n_1060;
wire n_1044;
wire n_1714;
wire n_521;
wire n_873;
wire n_1301;
wire n_1748;
wire n_1243;
wire n_1400;
wire n_342;
wire n_1466;
wire n_1527;
wire n_1513;
wire n_358;
wire n_1783;
wire n_608;
wire n_1538;
wire n_1037;
wire n_1329;
wire n_317;
wire n_1545;
wire n_1257;
wire n_1480;
wire n_1668;
wire n_1878;
wire n_1605;
wire n_1078;
wire n_266;
wire n_1897;
wire n_1161;
wire n_811;
wire n_624;
wire n_876;
wire n_791;
wire n_618;
wire n_1191;
wire n_736;
wire n_1025;
wire n_1215;
wire n_241;
wire n_1449;
wire n_687;
wire n_797;
wire n_1786;
wire n_480;
wire n_1327;
wire n_1475;
wire n_211;
wire n_642;
wire n_1804;
wire n_408;
wire n_1406;
wire n_595;
wire n_1405;
wire n_602;
wire n_1757;
wire n_592;
wire n_1499;
wire n_854;
wire n_1318;
wire n_393;
wire n_1632;
wire n_1769;
wire n_474;
wire n_1929;
wire n_805;
wire n_295;
wire n_1658;
wire n_1072;
wire n_695;
wire n_1526;
wire n_1305;
wire n_730;
wire n_386;
wire n_1596;
wire n_1281;
wire n_516;
wire n_1137;
wire n_1873;
wire n_1258;
wire n_640;
wire n_463;
wire n_1476;
wire n_1524;
wire n_1733;
wire n_1856;
wire n_943;
wire n_1118;
wire n_678;
wire n_651;
wire n_1874;
wire n_1293;
wire n_961;
wire n_469;
wire n_1046;
wire n_1807;
wire n_726;
wire n_1123;
wire n_1657;
wire n_878;
wire n_1784;
wire n_771;
wire n_1321;
wire n_752;
wire n_1488;
wire n_985;
wire n_421;
wire n_1330;
wire n_906;
wire n_1180;
wire n_1697;
wire n_283;
wire n_806;
wire n_1350;
wire n_1556;
wire n_649;
wire n_1561;
wire n_374;
wire n_1352;
wire n_1824;
wire n_643;
wire n_1492;
wire n_226;
wire n_1441;
wire n_1822;
wire n_682;
wire n_1616;
wire n_819;
wire n_586;
wire n_1324;
wire n_1429;
wire n_1778;
wire n_1776;
wire n_686;
wire n_605;
wire n_1154;
wire n_584;
wire n_1557;
wire n_1759;
wire n_1829;
wire n_1130;
wire n_1450;
wire n_349;
wire n_756;
wire n_1016;
wire n_1149;
wire n_1505;
wire n_979;
wire n_1642;
wire n_1815;
wire n_897;
wire n_949;
wire n_1493;
wire n_515;
wire n_807;
wire n_891;
wire n_885;
wire n_1659;
wire n_1864;
wire n_1887;
wire n_1208;
wire n_396;
wire n_802;
wire n_1151;
wire n_554;
wire n_960;
wire n_1256;
wire n_714;
wire n_790;
wire n_354;
wire n_725;
wire n_1577;
wire n_1448;
wire n_1009;
wire n_230;
wire n_1133;
wire n_883;
wire n_473;
wire n_1852;
wire n_801;
wire n_1286;
wire n_818;
wire n_1685;
wire n_779;
wire n_594;
wire n_1877;
wire n_1397;
wire n_1052;
wire n_272;
wire n_1333;
wire n_1306;
wire n_1849;
wire n_833;
wire n_1426;
wire n_879;
wire n_1117;
wire n_422;
wire n_1269;
wire n_1303;
wire n_1547;
wire n_1438;
wire n_1541;
wire n_597;
wire n_1047;
wire n_1472;
wire n_1593;
wire n_1050;
wire n_566;
wire n_1201;
wire n_1288;
wire n_858;
wire n_1185;
wire n_335;
wire n_1035;
wire n_1143;
wire n_344;
wire n_426;
wire n_433;
wire n_398;
wire n_210;
wire n_1090;
wire n_1367;
wire n_253;
wire n_928;
wire n_1153;
wire n_271;
wire n_465;
wire n_825;
wire n_1103;
wire n_732;
wire n_1565;
wire n_1192;
wire n_224;
wire n_894;
wire n_1380;
wire n_1624;
wire n_1801;
wire n_420;
wire n_1291;
wire n_562;
wire n_748;
wire n_510;
wire n_1045;
wire n_256;
wire n_1160;
wire n_1882;
wire n_1023;
wire n_1881;
wire n_988;
wire n_330;
wire n_914;
wire n_400;
wire n_689;
wire n_1116;
wire n_282;
wire n_328;
wire n_368;
wire n_467;
wire n_1511;
wire n_1422;
wire n_644;
wire n_1197;
wire n_276;
wire n_497;
wire n_1165;
wire n_1641;
wire n_538;
wire n_1517;
wire n_576;
wire n_843;
wire n_511;
wire n_455;
wire n_429;
wire n_588;
wire n_638;
wire n_1307;
wire n_1128;
wire n_1671;
wire n_1417;
wire n_1048;
wire n_775;
wire n_667;
wire n_1049;
wire n_869;
wire n_846;
wire n_1398;
wire n_1921;
wire n_1356;
wire n_1341;
wire n_1504;
wire n_1773;
wire n_1440;
wire n_1370;
wire n_1603;
wire n_305;
wire n_312;
wire n_728;
wire n_413;
wire n_715;
wire n_889;
wire n_1066;
wire n_1549;
wire n_935;
wire n_685;
wire n_911;
wire n_361;
wire n_623;
wire n_1712;
wire n_1403;
wire n_1065;
wire n_453;
wire n_1534;
wire n_810;
wire n_1290;
wire n_617;
wire n_543;
wire n_1362;
wire n_1559;
wire n_236;
wire n_683;
wire n_601;
wire n_565;
wire n_628;
wire n_1300;
wire n_743;
wire n_1194;
wire n_1647;
wire n_1546;
wire n_1420;
wire n_907;
wire n_1454;
wire n_660;
wire n_464;
wire n_962;
wire n_941;
wire n_1210;
wire n_847;
wire n_747;
wire n_1622;
wire n_1135;
wire n_918;
wire n_1885;
wire n_639;
wire n_452;
wire n_673;
wire n_1038;
wire n_414;
wire n_571;
wire n_1521;
wire n_1694;
wire n_284;
wire n_593;
wire n_1695;
wire n_1164;
wire n_609;
wire n_1193;
wire n_1345;
wire n_613;
wire n_1022;
wire n_1336;
wire n_1033;
wire n_1774;
wire n_409;
wire n_519;
wire n_384;
wire n_1166;
wire n_1056;
wire n_526;
wire n_1767;
wire n_1040;
wire n_674;
wire n_1158;
wire n_316;
wire n_1444;
wire n_1803;
wire n_820;
wire n_1749;
wire n_872;
wire n_1653;
wire n_254;
wire n_1157;
wire n_1584;
wire n_234;
wire n_848;
wire n_1664;
wire n_280;
wire n_629;
wire n_1739;
wire n_1814;
wire n_532;
wire n_1789;
wire n_763;
wire n_540;
wire n_216;
wire n_692;
wire n_1857;
wire n_984;
wire n_1687;
wire n_223;
wire n_1552;
wire n_750;
wire n_834;
wire n_1612;
wire n_800;
wire n_1816;
wire n_1910;
wire n_1756;
wire n_1606;
wire n_395;
wire n_621;
wire n_1587;
wire n_213;
wire n_1772;
wire n_1014;
wire n_724;
wire n_1427;
wire n_1481;
wire n_493;
wire n_1311;
wire n_1589;
wire n_1100;
wire n_585;
wire n_875;
wire n_1617;
wire n_827;
wire n_697;
wire n_622;
wire n_1626;
wire n_1335;
wire n_1715;
wire n_296;
wire n_880;
wire n_793;
wire n_1175;
wire n_751;
wire n_1027;
wire n_1070;
wire n_1621;
wire n_739;
wire n_1485;
wire n_1028;
wire n_1221;
wire n_530;
wire n_1785;
wire n_792;
wire n_1262;
wire n_580;
wire n_1579;
wire n_494;
wire n_434;
wire n_975;
wire n_229;
wire n_394;
wire n_923;
wire n_1645;
wire n_1124;
wire n_1381;
wire n_1494;
wire n_932;
wire n_1893;
wire n_1183;
wire n_1326;
wire n_1805;
wire n_981;
wire n_1110;
wire n_1758;
wire n_243;
wire n_1407;
wire n_1204;
wire n_1554;
wire n_994;
wire n_1360;
wire n_973;
wire n_268;
wire n_972;
wire n_856;
wire n_1248;
wire n_1176;
wire n_1564;
wire n_1054;
wire n_508;
wire n_1679;
wire n_1858;
wire n_353;
wire n_1678;
wire n_1482;
wire n_1361;
wire n_1601;
wire n_1057;
wire n_1834;
wire n_1011;
wire n_978;
wire n_1520;
wire n_1509;
wire n_828;
wire n_322;
wire n_1411;
wire n_1359;
wire n_558;
wire n_1721;
wire n_653;
wire n_1445;
wire n_1317;
wire n_783;
wire n_556;
wire n_1127;
wire n_1536;
wire n_1471;
wire n_1008;
wire n_332;
wire n_581;
wire n_294;
wire n_1024;
wire n_830;
wire n_987;
wire n_936;
wire n_1620;
wire n_1385;
wire n_1525;
wire n_541;
wire n_499;
wire n_1775;
wire n_788;
wire n_908;
wire n_1036;
wire n_341;
wire n_1270;
wire n_1167;
wire n_1272;
wire n_549;
wire n_591;
wire n_969;
wire n_919;
wire n_1663;
wire n_1625;
wire n_1926;
wire n_318;
wire n_1458;
wire n_244;
wire n_679;
wire n_1630;
wire n_220;
wire n_663;
wire n_1720;
wire n_443;
wire n_1412;
wire n_1738;
wire n_1550;
wire n_528;
wire n_1358;
wire n_1200;
wire n_387;
wire n_406;
wire n_826;
wire n_1922;
wire n_1735;
wire n_1788;
wire n_391;
wire n_940;
wire n_1537;
wire n_1077;
wire n_607;
wire n_956;
wire n_445;
wire n_1930;
wire n_765;
wire n_1809;
wire n_1843;
wire n_1904;
wire n_1268;
wire n_385;
wire n_917;
wire n_1271;
wire n_372;
wire n_1530;
wire n_631;
wire n_399;
wire n_1170;
wire n_1261;
wire n_702;
wire n_898;
wire n_857;
wire n_363;
wire n_1067;
wire n_968;
wire n_1323;
wire n_1235;
wire n_1462;
wire n_1064;
wire n_633;
wire n_900;
wire n_1446;
wire n_1282;
wire n_1701;
wire n_1093;
wire n_1551;
wire n_1755;
wire n_1285;
wire n_761;
wire n_733;
wire n_731;
wire n_336;
wire n_1813;
wire n_315;
wire n_311;
wire n_1452;
wire n_1573;
wire n_668;
wire n_758;
wire n_1106;
wire n_648;
wire n_784;
wire n_269;
wire n_816;
wire n_1322;
wire n_1473;
wire n_835;
wire n_446;
wire n_1076;
wire n_1348;
wire n_753;
wire n_1770;
wire n_701;
wire n_1003;
wire n_1125;
wire n_1710;
wire n_1865;
wire n_309;
wire n_1344;
wire n_1390;
wire n_485;
wire n_401;
wire n_1792;
wire n_504;
wire n_483;
wire n_435;
wire n_1141;
wire n_1629;
wire n_291;
wire n_1640;
wire n_822;
wire n_1094;
wire n_840;
wire n_1459;
wire n_1510;
wire n_1099;
wire n_839;
wire n_1754;
wire n_759;
wire n_567;
wire n_240;
wire n_369;
wire n_1727;
wire n_1575;
wire n_1848;
wire n_1892;
wire n_1172;
wire n_614;
wire n_1212;
wire n_831;
wire n_778;
wire n_1619;
wire n_323;
wire n_550;
wire n_1315;
wire n_1660;
wire n_1902;
wire n_997;
wire n_635;
wire n_694;
wire n_1643;
wire n_1320;
wire n_1113;
wire n_248;
wire n_1152;
wire n_1845;
wire n_921;
wire n_1615;
wire n_1236;
wire n_228;
wire n_1265;
wire n_1576;
wire n_1470;
wire n_671;
wire n_1533;
wire n_1806;
wire n_1409;
wire n_1148;
wire n_1588;
wire n_1684;
wire n_1673;
wire n_1334;
wire n_654;
wire n_1275;
wire n_488;
wire n_904;
wire n_505;
wire n_1696;
wire n_498;
wire n_1875;
wire n_1059;
wire n_684;
wire n_1039;
wire n_539;
wire n_1150;
wire n_977;
wire n_449;
wire n_392;
wire n_1628;
wire n_1289;
wire n_1831;
wire n_1497;
wire n_1866;
wire n_459;
wire n_1136;
wire n_1782;
wire n_458;
wire n_1190;
wire n_1600;
wire n_1144;
wire n_383;
wire n_838;
wire n_1558;
wire n_1316;
wire n_950;
wire n_1017;
wire n_711;
wire n_734;
wire n_1915;
wire n_723;
wire n_1393;
wire n_658;
wire n_630;
wire n_1369;
wire n_362;
wire n_310;
wire n_1781;
wire n_709;
wire n_809;
wire n_1686;
wire n_235;
wire n_881;
wire n_1019;
wire n_1477;
wire n_1777;
wire n_662;
wire n_641;
wire n_910;
wire n_290;
wire n_741;
wire n_939;
wire n_1410;
wire n_371;
wire n_217;
wire n_1114;
wire n_1325;
wire n_1742;
wire n_708;
wire n_308;
wire n_1223;
wire n_1768;
wire n_572;
wire n_1199;
wire n_865;
wire n_1273;
wire n_1041;
wire n_993;
wire n_1862;
wire n_948;
wire n_922;
wire n_1004;
wire n_1810;
wire n_448;
wire n_1347;
wire n_860;
wire n_1043;
wire n_255;
wire n_450;
wire n_1923;
wire n_1764;
wire n_896;
wire n_1737;
wire n_1479;
wire n_1613;
wire n_902;
wire n_1031;
wire n_1723;
wire n_1638;
wire n_853;
wire n_716;
wire n_1571;
wire n_1698;
wire n_1337;
wire n_774;
wire n_933;
wire n_1779;
wire n_596;
wire n_954;
wire n_1168;
wire n_1821;
wire n_219;
wire n_1310;
wire n_231;
wire n_656;
wire n_492;
wire n_574;
wire n_252;
wire n_664;
wire n_1591;
wire n_1229;
wire n_1683;
wire n_1896;
wire n_1732;
wire n_415;
wire n_1280;
wire n_544;
wire n_1516;
wire n_1186;
wire n_1705;
wire n_599;
wire n_768;
wire n_1091;
wire n_537;
wire n_1063;
wire n_991;
wire n_389;
wire n_1724;
wire n_1670;
wire n_1707;
wire n_1799;
wire n_1126;
wire n_1846;
wire n_1912;
wire n_938;
wire n_1891;
wire n_1328;
wire n_895;
wire n_304;
wire n_1639;
wire n_583;
wire n_1302;
wire n_1000;
wire n_313;
wire n_626;
wire n_378;
wire n_1581;
wire n_1928;
wire n_946;
wire n_757;
wire n_375;
wire n_1655;
wire n_1818;
wire n_1146;
wire n_1634;
wire n_1203;
wire n_998;
wire n_1699;
wire n_1598;
wire n_472;
wire n_937;
wire n_1474;
wire n_265;
wire n_1583;
wire n_1604;
wire n_208;
wire n_1631;
wire n_1702;
wire n_275;
wire n_1794;
wire n_1375;
wire n_204;
wire n_1232;
wire n_996;
wire n_1211;
wire n_1368;
wire n_963;
wire n_1264;
wire n_1082;
wire n_1725;
wire n_496;
wire n_1827;
wire n_866;
wire n_246;
wire n_925;
wire n_1752;
wire n_1313;
wire n_1001;
wire n_1722;
wire n_1115;
wire n_1339;
wire n_1002;
wire n_1644;
wire n_1051;
wire n_719;
wire n_263;
wire n_1102;
wire n_360;
wire n_1129;
wire n_1252;
wire n_250;
wire n_1464;
wire n_1296;
wire n_773;
wire n_1010;
wire n_882;
wire n_1249;
wire n_803;
wire n_1871;
wire n_718;
wire n_329;
wire n_1434;
wire n_340;
wire n_1905;
wire n_1569;
wire n_548;
wire n_289;
wire n_523;
wire n_1662;
wire n_457;
wire n_1299;
wire n_1870;
wire n_1925;
wire n_782;
wire n_364;
wire n_258;
wire n_431;
wire n_1861;
wire n_1228;
wire n_1931;
wire n_1244;
wire n_1796;
wire n_484;
wire n_411;
wire n_849;
wire n_1820;
wire n_357;
wire n_412;
wire n_1251;
wire n_447;
wire n_1421;
wire n_1762;
wire n_1233;
wire n_1808;
wire n_1574;
wire n_1672;
wire n_1635;
wire n_1704;
wire n_893;
wire n_1582;
wire n_841;
wire n_886;
wire n_1069;
wire n_359;
wire n_1308;
wire n_573;
wire n_796;
wire n_531;
wire n_1730;
wire n_1374;
wire n_1451;
wire n_1487;
wire n_675;

CKINVDCx20_ASAP7_75t_R g203 ( 
.A(n_6),
.Y(n_203)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_59),
.Y(n_204)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_117),
.Y(n_205)
);

CKINVDCx20_ASAP7_75t_R g206 ( 
.A(n_58),
.Y(n_206)
);

INVx2_ASAP7_75t_L g207 ( 
.A(n_116),
.Y(n_207)
);

BUFx8_ASAP7_75t_SL g208 ( 
.A(n_43),
.Y(n_208)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_97),
.Y(n_209)
);

CKINVDCx14_ASAP7_75t_R g210 ( 
.A(n_41),
.Y(n_210)
);

CKINVDCx5p33_ASAP7_75t_R g211 ( 
.A(n_159),
.Y(n_211)
);

CKINVDCx5p33_ASAP7_75t_R g212 ( 
.A(n_83),
.Y(n_212)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_29),
.Y(n_213)
);

INVx2_ASAP7_75t_L g214 ( 
.A(n_170),
.Y(n_214)
);

CKINVDCx5p33_ASAP7_75t_R g215 ( 
.A(n_42),
.Y(n_215)
);

CKINVDCx5p33_ASAP7_75t_R g216 ( 
.A(n_4),
.Y(n_216)
);

CKINVDCx5p33_ASAP7_75t_R g217 ( 
.A(n_60),
.Y(n_217)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_161),
.Y(n_218)
);

CKINVDCx20_ASAP7_75t_R g219 ( 
.A(n_88),
.Y(n_219)
);

CKINVDCx5p33_ASAP7_75t_R g220 ( 
.A(n_195),
.Y(n_220)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_102),
.Y(n_221)
);

CKINVDCx20_ASAP7_75t_R g222 ( 
.A(n_156),
.Y(n_222)
);

CKINVDCx20_ASAP7_75t_R g223 ( 
.A(n_171),
.Y(n_223)
);

CKINVDCx16_ASAP7_75t_R g224 ( 
.A(n_155),
.Y(n_224)
);

CKINVDCx5p33_ASAP7_75t_R g225 ( 
.A(n_149),
.Y(n_225)
);

BUFx10_ASAP7_75t_L g226 ( 
.A(n_152),
.Y(n_226)
);

CKINVDCx5p33_ASAP7_75t_R g227 ( 
.A(n_135),
.Y(n_227)
);

CKINVDCx20_ASAP7_75t_R g228 ( 
.A(n_175),
.Y(n_228)
);

BUFx3_ASAP7_75t_L g229 ( 
.A(n_129),
.Y(n_229)
);

INVx1_ASAP7_75t_SL g230 ( 
.A(n_168),
.Y(n_230)
);

CKINVDCx5p33_ASAP7_75t_R g231 ( 
.A(n_51),
.Y(n_231)
);

BUFx3_ASAP7_75t_L g232 ( 
.A(n_75),
.Y(n_232)
);

CKINVDCx5p33_ASAP7_75t_R g233 ( 
.A(n_84),
.Y(n_233)
);

CKINVDCx14_ASAP7_75t_R g234 ( 
.A(n_23),
.Y(n_234)
);

CKINVDCx5p33_ASAP7_75t_R g235 ( 
.A(n_60),
.Y(n_235)
);

CKINVDCx5p33_ASAP7_75t_R g236 ( 
.A(n_63),
.Y(n_236)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_160),
.Y(n_237)
);

CKINVDCx5p33_ASAP7_75t_R g238 ( 
.A(n_98),
.Y(n_238)
);

CKINVDCx5p33_ASAP7_75t_R g239 ( 
.A(n_145),
.Y(n_239)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_27),
.Y(n_240)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_163),
.Y(n_241)
);

CKINVDCx5p33_ASAP7_75t_R g242 ( 
.A(n_34),
.Y(n_242)
);

INVx1_ASAP7_75t_SL g243 ( 
.A(n_27),
.Y(n_243)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_150),
.Y(n_244)
);

CKINVDCx5p33_ASAP7_75t_R g245 ( 
.A(n_36),
.Y(n_245)
);

CKINVDCx5p33_ASAP7_75t_R g246 ( 
.A(n_130),
.Y(n_246)
);

CKINVDCx5p33_ASAP7_75t_R g247 ( 
.A(n_166),
.Y(n_247)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_196),
.Y(n_248)
);

CKINVDCx5p33_ASAP7_75t_R g249 ( 
.A(n_140),
.Y(n_249)
);

CKINVDCx5p33_ASAP7_75t_R g250 ( 
.A(n_109),
.Y(n_250)
);

CKINVDCx5p33_ASAP7_75t_R g251 ( 
.A(n_47),
.Y(n_251)
);

CKINVDCx20_ASAP7_75t_R g252 ( 
.A(n_65),
.Y(n_252)
);

BUFx3_ASAP7_75t_L g253 ( 
.A(n_108),
.Y(n_253)
);

BUFx10_ASAP7_75t_L g254 ( 
.A(n_200),
.Y(n_254)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_57),
.Y(n_255)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_99),
.Y(n_256)
);

CKINVDCx20_ASAP7_75t_R g257 ( 
.A(n_6),
.Y(n_257)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_0),
.Y(n_258)
);

BUFx6f_ASAP7_75t_L g259 ( 
.A(n_104),
.Y(n_259)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_39),
.Y(n_260)
);

CKINVDCx20_ASAP7_75t_R g261 ( 
.A(n_9),
.Y(n_261)
);

CKINVDCx5p33_ASAP7_75t_R g262 ( 
.A(n_67),
.Y(n_262)
);

CKINVDCx5p33_ASAP7_75t_R g263 ( 
.A(n_162),
.Y(n_263)
);

BUFx10_ASAP7_75t_L g264 ( 
.A(n_79),
.Y(n_264)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_11),
.Y(n_265)
);

CKINVDCx5p33_ASAP7_75t_R g266 ( 
.A(n_138),
.Y(n_266)
);

CKINVDCx5p33_ASAP7_75t_R g267 ( 
.A(n_87),
.Y(n_267)
);

CKINVDCx5p33_ASAP7_75t_R g268 ( 
.A(n_105),
.Y(n_268)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_32),
.Y(n_269)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_29),
.Y(n_270)
);

CKINVDCx5p33_ASAP7_75t_R g271 ( 
.A(n_143),
.Y(n_271)
);

INVx2_ASAP7_75t_SL g272 ( 
.A(n_183),
.Y(n_272)
);

INVx2_ASAP7_75t_SL g273 ( 
.A(n_34),
.Y(n_273)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_91),
.Y(n_274)
);

CKINVDCx14_ASAP7_75t_R g275 ( 
.A(n_131),
.Y(n_275)
);

BUFx3_ASAP7_75t_L g276 ( 
.A(n_5),
.Y(n_276)
);

CKINVDCx5p33_ASAP7_75t_R g277 ( 
.A(n_33),
.Y(n_277)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_58),
.Y(n_278)
);

CKINVDCx5p33_ASAP7_75t_R g279 ( 
.A(n_20),
.Y(n_279)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_57),
.Y(n_280)
);

CKINVDCx5p33_ASAP7_75t_R g281 ( 
.A(n_119),
.Y(n_281)
);

CKINVDCx5p33_ASAP7_75t_R g282 ( 
.A(n_123),
.Y(n_282)
);

CKINVDCx5p33_ASAP7_75t_R g283 ( 
.A(n_43),
.Y(n_283)
);

BUFx2_ASAP7_75t_L g284 ( 
.A(n_7),
.Y(n_284)
);

CKINVDCx20_ASAP7_75t_R g285 ( 
.A(n_178),
.Y(n_285)
);

CKINVDCx5p33_ASAP7_75t_R g286 ( 
.A(n_9),
.Y(n_286)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_142),
.Y(n_287)
);

INVx1_ASAP7_75t_SL g288 ( 
.A(n_146),
.Y(n_288)
);

CKINVDCx5p33_ASAP7_75t_R g289 ( 
.A(n_199),
.Y(n_289)
);

CKINVDCx5p33_ASAP7_75t_R g290 ( 
.A(n_74),
.Y(n_290)
);

INVx1_ASAP7_75t_SL g291 ( 
.A(n_148),
.Y(n_291)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_182),
.Y(n_292)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_80),
.Y(n_293)
);

INVx2_ASAP7_75t_L g294 ( 
.A(n_45),
.Y(n_294)
);

CKINVDCx5p33_ASAP7_75t_R g295 ( 
.A(n_76),
.Y(n_295)
);

CKINVDCx16_ASAP7_75t_R g296 ( 
.A(n_141),
.Y(n_296)
);

CKINVDCx5p33_ASAP7_75t_R g297 ( 
.A(n_126),
.Y(n_297)
);

BUFx6f_ASAP7_75t_L g298 ( 
.A(n_96),
.Y(n_298)
);

INVx4_ASAP7_75t_R g299 ( 
.A(n_44),
.Y(n_299)
);

CKINVDCx5p33_ASAP7_75t_R g300 ( 
.A(n_10),
.Y(n_300)
);

HB1xp67_ASAP7_75t_L g301 ( 
.A(n_95),
.Y(n_301)
);

CKINVDCx5p33_ASAP7_75t_R g302 ( 
.A(n_62),
.Y(n_302)
);

CKINVDCx5p33_ASAP7_75t_R g303 ( 
.A(n_111),
.Y(n_303)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_82),
.Y(n_304)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_100),
.Y(n_305)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_26),
.Y(n_306)
);

CKINVDCx5p33_ASAP7_75t_R g307 ( 
.A(n_89),
.Y(n_307)
);

CKINVDCx5p33_ASAP7_75t_R g308 ( 
.A(n_144),
.Y(n_308)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_21),
.Y(n_309)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_73),
.Y(n_310)
);

INVx2_ASAP7_75t_L g311 ( 
.A(n_15),
.Y(n_311)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_186),
.Y(n_312)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_106),
.Y(n_313)
);

BUFx3_ASAP7_75t_L g314 ( 
.A(n_31),
.Y(n_314)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_30),
.Y(n_315)
);

INVxp67_ASAP7_75t_SL g316 ( 
.A(n_62),
.Y(n_316)
);

CKINVDCx16_ASAP7_75t_R g317 ( 
.A(n_44),
.Y(n_317)
);

CKINVDCx5p33_ASAP7_75t_R g318 ( 
.A(n_39),
.Y(n_318)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_33),
.Y(n_319)
);

CKINVDCx5p33_ASAP7_75t_R g320 ( 
.A(n_63),
.Y(n_320)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_164),
.Y(n_321)
);

BUFx10_ASAP7_75t_L g322 ( 
.A(n_188),
.Y(n_322)
);

CKINVDCx5p33_ASAP7_75t_R g323 ( 
.A(n_179),
.Y(n_323)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_181),
.Y(n_324)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_125),
.Y(n_325)
);

CKINVDCx5p33_ASAP7_75t_R g326 ( 
.A(n_22),
.Y(n_326)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_127),
.Y(n_327)
);

CKINVDCx5p33_ASAP7_75t_R g328 ( 
.A(n_167),
.Y(n_328)
);

CKINVDCx5p33_ASAP7_75t_R g329 ( 
.A(n_197),
.Y(n_329)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_26),
.Y(n_330)
);

CKINVDCx5p33_ASAP7_75t_R g331 ( 
.A(n_86),
.Y(n_331)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_176),
.Y(n_332)
);

BUFx6f_ASAP7_75t_L g333 ( 
.A(n_0),
.Y(n_333)
);

BUFx10_ASAP7_75t_L g334 ( 
.A(n_121),
.Y(n_334)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_165),
.Y(n_335)
);

CKINVDCx5p33_ASAP7_75t_R g336 ( 
.A(n_20),
.Y(n_336)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_2),
.Y(n_337)
);

BUFx6f_ASAP7_75t_L g338 ( 
.A(n_35),
.Y(n_338)
);

BUFx6f_ASAP7_75t_L g339 ( 
.A(n_31),
.Y(n_339)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_72),
.Y(n_340)
);

CKINVDCx5p33_ASAP7_75t_R g341 ( 
.A(n_118),
.Y(n_341)
);

CKINVDCx20_ASAP7_75t_R g342 ( 
.A(n_90),
.Y(n_342)
);

CKINVDCx5p33_ASAP7_75t_R g343 ( 
.A(n_193),
.Y(n_343)
);

INVx1_ASAP7_75t_L g344 ( 
.A(n_151),
.Y(n_344)
);

CKINVDCx5p33_ASAP7_75t_R g345 ( 
.A(n_187),
.Y(n_345)
);

INVx1_ASAP7_75t_L g346 ( 
.A(n_134),
.Y(n_346)
);

CKINVDCx5p33_ASAP7_75t_R g347 ( 
.A(n_128),
.Y(n_347)
);

BUFx10_ASAP7_75t_L g348 ( 
.A(n_133),
.Y(n_348)
);

CKINVDCx5p33_ASAP7_75t_R g349 ( 
.A(n_3),
.Y(n_349)
);

CKINVDCx5p33_ASAP7_75t_R g350 ( 
.A(n_48),
.Y(n_350)
);

INVx1_ASAP7_75t_L g351 ( 
.A(n_136),
.Y(n_351)
);

INVx1_ASAP7_75t_L g352 ( 
.A(n_30),
.Y(n_352)
);

BUFx10_ASAP7_75t_L g353 ( 
.A(n_65),
.Y(n_353)
);

INVxp67_ASAP7_75t_L g354 ( 
.A(n_120),
.Y(n_354)
);

INVx1_ASAP7_75t_L g355 ( 
.A(n_48),
.Y(n_355)
);

CKINVDCx5p33_ASAP7_75t_R g356 ( 
.A(n_59),
.Y(n_356)
);

CKINVDCx5p33_ASAP7_75t_R g357 ( 
.A(n_113),
.Y(n_357)
);

BUFx10_ASAP7_75t_L g358 ( 
.A(n_45),
.Y(n_358)
);

CKINVDCx5p33_ASAP7_75t_R g359 ( 
.A(n_7),
.Y(n_359)
);

CKINVDCx5p33_ASAP7_75t_R g360 ( 
.A(n_36),
.Y(n_360)
);

CKINVDCx20_ASAP7_75t_R g361 ( 
.A(n_198),
.Y(n_361)
);

CKINVDCx20_ASAP7_75t_R g362 ( 
.A(n_40),
.Y(n_362)
);

INVx1_ASAP7_75t_L g363 ( 
.A(n_154),
.Y(n_363)
);

BUFx2_ASAP7_75t_L g364 ( 
.A(n_184),
.Y(n_364)
);

CKINVDCx5p33_ASAP7_75t_R g365 ( 
.A(n_4),
.Y(n_365)
);

INVx2_ASAP7_75t_SL g366 ( 
.A(n_94),
.Y(n_366)
);

INVx1_ASAP7_75t_SL g367 ( 
.A(n_101),
.Y(n_367)
);

CKINVDCx16_ASAP7_75t_R g368 ( 
.A(n_13),
.Y(n_368)
);

CKINVDCx5p33_ASAP7_75t_R g369 ( 
.A(n_8),
.Y(n_369)
);

CKINVDCx5p33_ASAP7_75t_R g370 ( 
.A(n_21),
.Y(n_370)
);

CKINVDCx20_ASAP7_75t_R g371 ( 
.A(n_115),
.Y(n_371)
);

INVx1_ASAP7_75t_SL g372 ( 
.A(n_81),
.Y(n_372)
);

CKINVDCx5p33_ASAP7_75t_R g373 ( 
.A(n_12),
.Y(n_373)
);

CKINVDCx5p33_ASAP7_75t_R g374 ( 
.A(n_52),
.Y(n_374)
);

CKINVDCx5p33_ASAP7_75t_R g375 ( 
.A(n_66),
.Y(n_375)
);

CKINVDCx5p33_ASAP7_75t_R g376 ( 
.A(n_24),
.Y(n_376)
);

CKINVDCx5p33_ASAP7_75t_R g377 ( 
.A(n_192),
.Y(n_377)
);

CKINVDCx5p33_ASAP7_75t_R g378 ( 
.A(n_110),
.Y(n_378)
);

CKINVDCx5p33_ASAP7_75t_R g379 ( 
.A(n_12),
.Y(n_379)
);

CKINVDCx5p33_ASAP7_75t_R g380 ( 
.A(n_46),
.Y(n_380)
);

CKINVDCx5p33_ASAP7_75t_R g381 ( 
.A(n_47),
.Y(n_381)
);

CKINVDCx5p33_ASAP7_75t_R g382 ( 
.A(n_66),
.Y(n_382)
);

BUFx3_ASAP7_75t_L g383 ( 
.A(n_69),
.Y(n_383)
);

INVx2_ASAP7_75t_L g384 ( 
.A(n_122),
.Y(n_384)
);

INVx1_ASAP7_75t_L g385 ( 
.A(n_93),
.Y(n_385)
);

INVx1_ASAP7_75t_L g386 ( 
.A(n_107),
.Y(n_386)
);

CKINVDCx5p33_ASAP7_75t_R g387 ( 
.A(n_191),
.Y(n_387)
);

INVx1_ASAP7_75t_L g388 ( 
.A(n_172),
.Y(n_388)
);

CKINVDCx5p33_ASAP7_75t_R g389 ( 
.A(n_52),
.Y(n_389)
);

CKINVDCx5p33_ASAP7_75t_R g390 ( 
.A(n_18),
.Y(n_390)
);

CKINVDCx16_ASAP7_75t_R g391 ( 
.A(n_40),
.Y(n_391)
);

HB1xp67_ASAP7_75t_L g392 ( 
.A(n_11),
.Y(n_392)
);

CKINVDCx5p33_ASAP7_75t_R g393 ( 
.A(n_112),
.Y(n_393)
);

INVx1_ASAP7_75t_L g394 ( 
.A(n_157),
.Y(n_394)
);

CKINVDCx5p33_ASAP7_75t_R g395 ( 
.A(n_194),
.Y(n_395)
);

INVx1_ASAP7_75t_L g396 ( 
.A(n_132),
.Y(n_396)
);

INVx1_ASAP7_75t_SL g397 ( 
.A(n_16),
.Y(n_397)
);

CKINVDCx5p33_ASAP7_75t_R g398 ( 
.A(n_23),
.Y(n_398)
);

INVx1_ASAP7_75t_L g399 ( 
.A(n_8),
.Y(n_399)
);

CKINVDCx5p33_ASAP7_75t_R g400 ( 
.A(n_139),
.Y(n_400)
);

CKINVDCx5p33_ASAP7_75t_R g401 ( 
.A(n_92),
.Y(n_401)
);

INVx2_ASAP7_75t_L g402 ( 
.A(n_10),
.Y(n_402)
);

CKINVDCx5p33_ASAP7_75t_R g403 ( 
.A(n_147),
.Y(n_403)
);

INVxp33_ASAP7_75t_SL g404 ( 
.A(n_392),
.Y(n_404)
);

INVx1_ASAP7_75t_L g405 ( 
.A(n_333),
.Y(n_405)
);

HB1xp67_ASAP7_75t_L g406 ( 
.A(n_284),
.Y(n_406)
);

INVx1_ASAP7_75t_L g407 ( 
.A(n_333),
.Y(n_407)
);

INVx1_ASAP7_75t_SL g408 ( 
.A(n_208),
.Y(n_408)
);

BUFx6f_ASAP7_75t_L g409 ( 
.A(n_259),
.Y(n_409)
);

INVx1_ASAP7_75t_L g410 ( 
.A(n_333),
.Y(n_410)
);

INVxp67_ASAP7_75t_L g411 ( 
.A(n_273),
.Y(n_411)
);

INVx1_ASAP7_75t_L g412 ( 
.A(n_333),
.Y(n_412)
);

NOR2xp67_ASAP7_75t_L g413 ( 
.A(n_273),
.B(n_1),
.Y(n_413)
);

NOR2xp33_ASAP7_75t_L g414 ( 
.A(n_364),
.B(n_1),
.Y(n_414)
);

CKINVDCx5p33_ASAP7_75t_R g415 ( 
.A(n_317),
.Y(n_415)
);

CKINVDCx20_ASAP7_75t_R g416 ( 
.A(n_210),
.Y(n_416)
);

INVx1_ASAP7_75t_L g417 ( 
.A(n_333),
.Y(n_417)
);

INVx1_ASAP7_75t_L g418 ( 
.A(n_338),
.Y(n_418)
);

CKINVDCx5p33_ASAP7_75t_R g419 ( 
.A(n_368),
.Y(n_419)
);

CKINVDCx5p33_ASAP7_75t_R g420 ( 
.A(n_391),
.Y(n_420)
);

INVx1_ASAP7_75t_L g421 ( 
.A(n_338),
.Y(n_421)
);

CKINVDCx20_ASAP7_75t_R g422 ( 
.A(n_234),
.Y(n_422)
);

HB1xp67_ASAP7_75t_L g423 ( 
.A(n_215),
.Y(n_423)
);

INVx1_ASAP7_75t_L g424 ( 
.A(n_338),
.Y(n_424)
);

CKINVDCx5p33_ASAP7_75t_R g425 ( 
.A(n_219),
.Y(n_425)
);

INVxp67_ASAP7_75t_SL g426 ( 
.A(n_276),
.Y(n_426)
);

NOR2xp33_ASAP7_75t_L g427 ( 
.A(n_301),
.B(n_2),
.Y(n_427)
);

CKINVDCx20_ASAP7_75t_R g428 ( 
.A(n_222),
.Y(n_428)
);

CKINVDCx5p33_ASAP7_75t_R g429 ( 
.A(n_223),
.Y(n_429)
);

CKINVDCx5p33_ASAP7_75t_R g430 ( 
.A(n_228),
.Y(n_430)
);

CKINVDCx20_ASAP7_75t_R g431 ( 
.A(n_285),
.Y(n_431)
);

INVx1_ASAP7_75t_L g432 ( 
.A(n_338),
.Y(n_432)
);

INVx1_ASAP7_75t_L g433 ( 
.A(n_338),
.Y(n_433)
);

CKINVDCx5p33_ASAP7_75t_R g434 ( 
.A(n_342),
.Y(n_434)
);

INVx1_ASAP7_75t_L g435 ( 
.A(n_339),
.Y(n_435)
);

INVx1_ASAP7_75t_L g436 ( 
.A(n_276),
.Y(n_436)
);

CKINVDCx14_ASAP7_75t_R g437 ( 
.A(n_275),
.Y(n_437)
);

CKINVDCx5p33_ASAP7_75t_R g438 ( 
.A(n_361),
.Y(n_438)
);

INVxp67_ASAP7_75t_SL g439 ( 
.A(n_314),
.Y(n_439)
);

CKINVDCx5p33_ASAP7_75t_R g440 ( 
.A(n_371),
.Y(n_440)
);

CKINVDCx20_ASAP7_75t_R g441 ( 
.A(n_203),
.Y(n_441)
);

INVx1_ASAP7_75t_L g442 ( 
.A(n_339),
.Y(n_442)
);

CKINVDCx5p33_ASAP7_75t_R g443 ( 
.A(n_262),
.Y(n_443)
);

INVx1_ASAP7_75t_L g444 ( 
.A(n_339),
.Y(n_444)
);

CKINVDCx5p33_ASAP7_75t_R g445 ( 
.A(n_277),
.Y(n_445)
);

CKINVDCx5p33_ASAP7_75t_R g446 ( 
.A(n_279),
.Y(n_446)
);

NOR2xp33_ASAP7_75t_L g447 ( 
.A(n_314),
.B(n_3),
.Y(n_447)
);

INVx1_ASAP7_75t_L g448 ( 
.A(n_339),
.Y(n_448)
);

INVx1_ASAP7_75t_L g449 ( 
.A(n_339),
.Y(n_449)
);

INVxp67_ASAP7_75t_L g450 ( 
.A(n_353),
.Y(n_450)
);

CKINVDCx5p33_ASAP7_75t_R g451 ( 
.A(n_283),
.Y(n_451)
);

INVx1_ASAP7_75t_L g452 ( 
.A(n_294),
.Y(n_452)
);

INVx1_ASAP7_75t_L g453 ( 
.A(n_294),
.Y(n_453)
);

INVx1_ASAP7_75t_L g454 ( 
.A(n_311),
.Y(n_454)
);

CKINVDCx5p33_ASAP7_75t_R g455 ( 
.A(n_286),
.Y(n_455)
);

CKINVDCx5p33_ASAP7_75t_R g456 ( 
.A(n_300),
.Y(n_456)
);

CKINVDCx5p33_ASAP7_75t_R g457 ( 
.A(n_302),
.Y(n_457)
);

CKINVDCx5p33_ASAP7_75t_R g458 ( 
.A(n_318),
.Y(n_458)
);

INVx1_ASAP7_75t_L g459 ( 
.A(n_311),
.Y(n_459)
);

INVx1_ASAP7_75t_L g460 ( 
.A(n_402),
.Y(n_460)
);

INVx1_ASAP7_75t_L g461 ( 
.A(n_402),
.Y(n_461)
);

INVx1_ASAP7_75t_L g462 ( 
.A(n_207),
.Y(n_462)
);

NOR2xp67_ASAP7_75t_L g463 ( 
.A(n_215),
.B(n_5),
.Y(n_463)
);

INVx1_ASAP7_75t_L g464 ( 
.A(n_207),
.Y(n_464)
);

INVx1_ASAP7_75t_L g465 ( 
.A(n_214),
.Y(n_465)
);

CKINVDCx5p33_ASAP7_75t_R g466 ( 
.A(n_320),
.Y(n_466)
);

CKINVDCx20_ASAP7_75t_R g467 ( 
.A(n_206),
.Y(n_467)
);

CKINVDCx5p33_ASAP7_75t_R g468 ( 
.A(n_326),
.Y(n_468)
);

INVx1_ASAP7_75t_L g469 ( 
.A(n_214),
.Y(n_469)
);

CKINVDCx20_ASAP7_75t_R g470 ( 
.A(n_252),
.Y(n_470)
);

NAND2xp5_ASAP7_75t_L g471 ( 
.A(n_205),
.B(n_13),
.Y(n_471)
);

CKINVDCx20_ASAP7_75t_R g472 ( 
.A(n_257),
.Y(n_472)
);

INVx1_ASAP7_75t_L g473 ( 
.A(n_384),
.Y(n_473)
);

CKINVDCx5p33_ASAP7_75t_R g474 ( 
.A(n_336),
.Y(n_474)
);

CKINVDCx5p33_ASAP7_75t_R g475 ( 
.A(n_216),
.Y(n_475)
);

INVxp67_ASAP7_75t_L g476 ( 
.A(n_353),
.Y(n_476)
);

INVx1_ASAP7_75t_L g477 ( 
.A(n_384),
.Y(n_477)
);

CKINVDCx5p33_ASAP7_75t_R g478 ( 
.A(n_216),
.Y(n_478)
);

NOR2xp33_ASAP7_75t_L g479 ( 
.A(n_383),
.B(n_14),
.Y(n_479)
);

CKINVDCx20_ASAP7_75t_R g480 ( 
.A(n_261),
.Y(n_480)
);

CKINVDCx20_ASAP7_75t_R g481 ( 
.A(n_362),
.Y(n_481)
);

INVx1_ASAP7_75t_L g482 ( 
.A(n_383),
.Y(n_482)
);

CKINVDCx20_ASAP7_75t_R g483 ( 
.A(n_224),
.Y(n_483)
);

INVx1_ASAP7_75t_L g484 ( 
.A(n_204),
.Y(n_484)
);

CKINVDCx5p33_ASAP7_75t_R g485 ( 
.A(n_217),
.Y(n_485)
);

INVxp67_ASAP7_75t_SL g486 ( 
.A(n_213),
.Y(n_486)
);

CKINVDCx5p33_ASAP7_75t_R g487 ( 
.A(n_217),
.Y(n_487)
);

INVx2_ASAP7_75t_L g488 ( 
.A(n_229),
.Y(n_488)
);

CKINVDCx5p33_ASAP7_75t_R g489 ( 
.A(n_231),
.Y(n_489)
);

CKINVDCx5p33_ASAP7_75t_R g490 ( 
.A(n_231),
.Y(n_490)
);

CKINVDCx5p33_ASAP7_75t_R g491 ( 
.A(n_235),
.Y(n_491)
);

INVx1_ASAP7_75t_L g492 ( 
.A(n_240),
.Y(n_492)
);

CKINVDCx20_ASAP7_75t_R g493 ( 
.A(n_296),
.Y(n_493)
);

HB1xp67_ASAP7_75t_L g494 ( 
.A(n_235),
.Y(n_494)
);

CKINVDCx5p33_ASAP7_75t_R g495 ( 
.A(n_236),
.Y(n_495)
);

INVx1_ASAP7_75t_L g496 ( 
.A(n_255),
.Y(n_496)
);

INVx1_ASAP7_75t_L g497 ( 
.A(n_258),
.Y(n_497)
);

CKINVDCx5p33_ASAP7_75t_R g498 ( 
.A(n_236),
.Y(n_498)
);

INVx1_ASAP7_75t_L g499 ( 
.A(n_260),
.Y(n_499)
);

INVx1_ASAP7_75t_L g500 ( 
.A(n_265),
.Y(n_500)
);

CKINVDCx20_ASAP7_75t_R g501 ( 
.A(n_226),
.Y(n_501)
);

CKINVDCx20_ASAP7_75t_R g502 ( 
.A(n_226),
.Y(n_502)
);

CKINVDCx5p33_ASAP7_75t_R g503 ( 
.A(n_242),
.Y(n_503)
);

CKINVDCx20_ASAP7_75t_R g504 ( 
.A(n_226),
.Y(n_504)
);

INVx2_ASAP7_75t_L g505 ( 
.A(n_229),
.Y(n_505)
);

CKINVDCx5p33_ASAP7_75t_R g506 ( 
.A(n_242),
.Y(n_506)
);

INVx1_ASAP7_75t_L g507 ( 
.A(n_405),
.Y(n_507)
);

AND2x2_ASAP7_75t_L g508 ( 
.A(n_426),
.B(n_254),
.Y(n_508)
);

INVx2_ASAP7_75t_L g509 ( 
.A(n_409),
.Y(n_509)
);

INVx3_ASAP7_75t_L g510 ( 
.A(n_409),
.Y(n_510)
);

NOR2x1_ASAP7_75t_L g511 ( 
.A(n_462),
.B(n_232),
.Y(n_511)
);

NAND2xp5_ASAP7_75t_L g512 ( 
.A(n_488),
.B(n_209),
.Y(n_512)
);

BUFx6f_ASAP7_75t_L g513 ( 
.A(n_409),
.Y(n_513)
);

OAI21x1_ASAP7_75t_L g514 ( 
.A1(n_471),
.A2(n_464),
.B(n_462),
.Y(n_514)
);

INVx2_ASAP7_75t_L g515 ( 
.A(n_409),
.Y(n_515)
);

BUFx8_ASAP7_75t_L g516 ( 
.A(n_488),
.Y(n_516)
);

INVx1_ASAP7_75t_L g517 ( 
.A(n_405),
.Y(n_517)
);

NOR2xp33_ASAP7_75t_L g518 ( 
.A(n_437),
.B(n_354),
.Y(n_518)
);

CKINVDCx20_ASAP7_75t_R g519 ( 
.A(n_441),
.Y(n_519)
);

INVx1_ASAP7_75t_L g520 ( 
.A(n_407),
.Y(n_520)
);

NAND2xp5_ASAP7_75t_L g521 ( 
.A(n_505),
.B(n_218),
.Y(n_521)
);

AND2x2_ASAP7_75t_L g522 ( 
.A(n_439),
.B(n_254),
.Y(n_522)
);

INVx2_ASAP7_75t_L g523 ( 
.A(n_409),
.Y(n_523)
);

AND2x2_ASAP7_75t_L g524 ( 
.A(n_436),
.B(n_254),
.Y(n_524)
);

INVx1_ASAP7_75t_L g525 ( 
.A(n_407),
.Y(n_525)
);

INVx2_ASAP7_75t_L g526 ( 
.A(n_410),
.Y(n_526)
);

INVx1_ASAP7_75t_L g527 ( 
.A(n_410),
.Y(n_527)
);

AND2x4_ASAP7_75t_L g528 ( 
.A(n_505),
.B(n_232),
.Y(n_528)
);

INVx1_ASAP7_75t_L g529 ( 
.A(n_412),
.Y(n_529)
);

INVx1_ASAP7_75t_L g530 ( 
.A(n_412),
.Y(n_530)
);

NAND2xp5_ASAP7_75t_SL g531 ( 
.A(n_443),
.B(n_264),
.Y(n_531)
);

AND2x2_ASAP7_75t_L g532 ( 
.A(n_482),
.B(n_484),
.Y(n_532)
);

INVx5_ASAP7_75t_L g533 ( 
.A(n_464),
.Y(n_533)
);

NAND2xp33_ASAP7_75t_L g534 ( 
.A(n_445),
.B(n_211),
.Y(n_534)
);

INVxp67_ASAP7_75t_L g535 ( 
.A(n_423),
.Y(n_535)
);

AND2x4_ASAP7_75t_L g536 ( 
.A(n_465),
.B(n_253),
.Y(n_536)
);

INVx6_ASAP7_75t_L g537 ( 
.A(n_486),
.Y(n_537)
);

INVx1_ASAP7_75t_L g538 ( 
.A(n_417),
.Y(n_538)
);

NOR2x1_ASAP7_75t_L g539 ( 
.A(n_465),
.B(n_253),
.Y(n_539)
);

CKINVDCx5p33_ASAP7_75t_R g540 ( 
.A(n_425),
.Y(n_540)
);

INVxp67_ASAP7_75t_L g541 ( 
.A(n_494),
.Y(n_541)
);

AND2x2_ASAP7_75t_L g542 ( 
.A(n_484),
.B(n_264),
.Y(n_542)
);

INVx1_ASAP7_75t_L g543 ( 
.A(n_417),
.Y(n_543)
);

BUFx6f_ASAP7_75t_L g544 ( 
.A(n_418),
.Y(n_544)
);

INVx2_ASAP7_75t_L g545 ( 
.A(n_418),
.Y(n_545)
);

NAND2xp5_ASAP7_75t_SL g546 ( 
.A(n_446),
.B(n_264),
.Y(n_546)
);

NAND2xp5_ASAP7_75t_L g547 ( 
.A(n_469),
.B(n_221),
.Y(n_547)
);

INVx2_ASAP7_75t_L g548 ( 
.A(n_421),
.Y(n_548)
);

INVx3_ASAP7_75t_L g549 ( 
.A(n_421),
.Y(n_549)
);

INVx1_ASAP7_75t_L g550 ( 
.A(n_424),
.Y(n_550)
);

INVx1_ASAP7_75t_L g551 ( 
.A(n_424),
.Y(n_551)
);

INVx3_ASAP7_75t_L g552 ( 
.A(n_432),
.Y(n_552)
);

INVx1_ASAP7_75t_L g553 ( 
.A(n_432),
.Y(n_553)
);

NAND2xp5_ASAP7_75t_L g554 ( 
.A(n_469),
.B(n_237),
.Y(n_554)
);

CKINVDCx5p33_ASAP7_75t_R g555 ( 
.A(n_429),
.Y(n_555)
);

AND2x2_ASAP7_75t_L g556 ( 
.A(n_492),
.B(n_322),
.Y(n_556)
);

INVx1_ASAP7_75t_L g557 ( 
.A(n_433),
.Y(n_557)
);

AOI22xp5_ASAP7_75t_L g558 ( 
.A1(n_404),
.A2(n_243),
.B1(n_397),
.B2(n_356),
.Y(n_558)
);

BUFx6f_ASAP7_75t_L g559 ( 
.A(n_433),
.Y(n_559)
);

INVx2_ASAP7_75t_L g560 ( 
.A(n_435),
.Y(n_560)
);

INVx1_ASAP7_75t_L g561 ( 
.A(n_435),
.Y(n_561)
);

HB1xp67_ASAP7_75t_L g562 ( 
.A(n_406),
.Y(n_562)
);

INVx2_ASAP7_75t_L g563 ( 
.A(n_442),
.Y(n_563)
);

INVx1_ASAP7_75t_L g564 ( 
.A(n_442),
.Y(n_564)
);

AND2x4_ASAP7_75t_L g565 ( 
.A(n_473),
.B(n_272),
.Y(n_565)
);

INVx1_ASAP7_75t_L g566 ( 
.A(n_444),
.Y(n_566)
);

NOR2xp33_ASAP7_75t_L g567 ( 
.A(n_451),
.B(n_272),
.Y(n_567)
);

INVx2_ASAP7_75t_L g568 ( 
.A(n_444),
.Y(n_568)
);

INVx2_ASAP7_75t_L g569 ( 
.A(n_448),
.Y(n_569)
);

INVx1_ASAP7_75t_L g570 ( 
.A(n_448),
.Y(n_570)
);

NAND2xp5_ASAP7_75t_L g571 ( 
.A(n_473),
.B(n_241),
.Y(n_571)
);

BUFx6f_ASAP7_75t_L g572 ( 
.A(n_449),
.Y(n_572)
);

OAI22xp5_ASAP7_75t_L g573 ( 
.A1(n_450),
.A2(n_365),
.B1(n_245),
.B2(n_356),
.Y(n_573)
);

NAND2xp5_ASAP7_75t_L g574 ( 
.A(n_477),
.B(n_244),
.Y(n_574)
);

BUFx6f_ASAP7_75t_L g575 ( 
.A(n_449),
.Y(n_575)
);

INVx1_ASAP7_75t_L g576 ( 
.A(n_477),
.Y(n_576)
);

CKINVDCx20_ASAP7_75t_R g577 ( 
.A(n_467),
.Y(n_577)
);

INVx2_ASAP7_75t_L g578 ( 
.A(n_452),
.Y(n_578)
);

AND2x4_ASAP7_75t_L g579 ( 
.A(n_492),
.B(n_366),
.Y(n_579)
);

BUFx6f_ASAP7_75t_L g580 ( 
.A(n_452),
.Y(n_580)
);

INVx1_ASAP7_75t_L g581 ( 
.A(n_453),
.Y(n_581)
);

BUFx6f_ASAP7_75t_L g582 ( 
.A(n_453),
.Y(n_582)
);

INVx1_ASAP7_75t_L g583 ( 
.A(n_454),
.Y(n_583)
);

AND2x4_ASAP7_75t_L g584 ( 
.A(n_497),
.B(n_499),
.Y(n_584)
);

NOR2xp33_ASAP7_75t_L g585 ( 
.A(n_455),
.B(n_366),
.Y(n_585)
);

OA21x2_ASAP7_75t_L g586 ( 
.A1(n_454),
.A2(n_256),
.B(n_248),
.Y(n_586)
);

INVx3_ASAP7_75t_L g587 ( 
.A(n_459),
.Y(n_587)
);

AND3x1_ASAP7_75t_L g588 ( 
.A(n_427),
.B(n_270),
.C(n_269),
.Y(n_588)
);

INVx2_ASAP7_75t_L g589 ( 
.A(n_549),
.Y(n_589)
);

NAND2xp5_ASAP7_75t_L g590 ( 
.A(n_542),
.B(n_456),
.Y(n_590)
);

INVx1_ASAP7_75t_L g591 ( 
.A(n_514),
.Y(n_591)
);

NAND2xp5_ASAP7_75t_L g592 ( 
.A(n_542),
.B(n_457),
.Y(n_592)
);

AOI22xp33_ASAP7_75t_L g593 ( 
.A1(n_537),
.A2(n_414),
.B1(n_413),
.B2(n_447),
.Y(n_593)
);

INVx2_ASAP7_75t_L g594 ( 
.A(n_549),
.Y(n_594)
);

BUFx4f_ASAP7_75t_L g595 ( 
.A(n_586),
.Y(n_595)
);

BUFx2_ASAP7_75t_L g596 ( 
.A(n_562),
.Y(n_596)
);

AOI22xp5_ASAP7_75t_L g597 ( 
.A1(n_588),
.A2(n_479),
.B1(n_463),
.B2(n_316),
.Y(n_597)
);

INVx2_ASAP7_75t_SL g598 ( 
.A(n_537),
.Y(n_598)
);

OR2x2_ASAP7_75t_L g599 ( 
.A(n_562),
.B(n_430),
.Y(n_599)
);

AND2x2_ASAP7_75t_SL g600 ( 
.A(n_588),
.B(n_542),
.Y(n_600)
);

NAND2xp5_ASAP7_75t_SL g601 ( 
.A(n_556),
.B(n_458),
.Y(n_601)
);

INVxp33_ASAP7_75t_L g602 ( 
.A(n_558),
.Y(n_602)
);

INVx2_ASAP7_75t_L g603 ( 
.A(n_549),
.Y(n_603)
);

NAND2xp5_ASAP7_75t_L g604 ( 
.A(n_556),
.B(n_466),
.Y(n_604)
);

INVx3_ASAP7_75t_L g605 ( 
.A(n_549),
.Y(n_605)
);

AND2x6_ASAP7_75t_L g606 ( 
.A(n_556),
.B(n_259),
.Y(n_606)
);

BUFx4f_ASAP7_75t_L g607 ( 
.A(n_586),
.Y(n_607)
);

INVx4_ASAP7_75t_L g608 ( 
.A(n_586),
.Y(n_608)
);

INVx2_ASAP7_75t_L g609 ( 
.A(n_552),
.Y(n_609)
);

INVx2_ASAP7_75t_L g610 ( 
.A(n_552),
.Y(n_610)
);

INVxp33_ASAP7_75t_SL g611 ( 
.A(n_540),
.Y(n_611)
);

INVx1_ASAP7_75t_L g612 ( 
.A(n_514),
.Y(n_612)
);

NAND2xp33_ASAP7_75t_L g613 ( 
.A(n_524),
.B(n_468),
.Y(n_613)
);

INVx1_ASAP7_75t_L g614 ( 
.A(n_514),
.Y(n_614)
);

INVx1_ASAP7_75t_L g615 ( 
.A(n_507),
.Y(n_615)
);

NOR2xp33_ASAP7_75t_L g616 ( 
.A(n_537),
.B(n_474),
.Y(n_616)
);

INVx3_ASAP7_75t_L g617 ( 
.A(n_552),
.Y(n_617)
);

OR2x6_ASAP7_75t_L g618 ( 
.A(n_537),
.B(n_497),
.Y(n_618)
);

INVx2_ASAP7_75t_L g619 ( 
.A(n_552),
.Y(n_619)
);

INVx2_ASAP7_75t_L g620 ( 
.A(n_526),
.Y(n_620)
);

INVx2_ASAP7_75t_L g621 ( 
.A(n_526),
.Y(n_621)
);

INVx2_ASAP7_75t_L g622 ( 
.A(n_526),
.Y(n_622)
);

BUFx2_ASAP7_75t_L g623 ( 
.A(n_555),
.Y(n_623)
);

INVx1_ASAP7_75t_L g624 ( 
.A(n_507),
.Y(n_624)
);

INVx2_ASAP7_75t_L g625 ( 
.A(n_545),
.Y(n_625)
);

INVxp67_ASAP7_75t_SL g626 ( 
.A(n_512),
.Y(n_626)
);

INVxp67_ASAP7_75t_SL g627 ( 
.A(n_512),
.Y(n_627)
);

NOR2xp33_ASAP7_75t_L g628 ( 
.A(n_537),
.B(n_475),
.Y(n_628)
);

INVx2_ASAP7_75t_L g629 ( 
.A(n_545),
.Y(n_629)
);

NAND2xp5_ASAP7_75t_L g630 ( 
.A(n_567),
.B(n_478),
.Y(n_630)
);

INVx2_ASAP7_75t_L g631 ( 
.A(n_545),
.Y(n_631)
);

INVx3_ASAP7_75t_L g632 ( 
.A(n_544),
.Y(n_632)
);

NAND2xp5_ASAP7_75t_L g633 ( 
.A(n_585),
.B(n_485),
.Y(n_633)
);

INVx2_ASAP7_75t_L g634 ( 
.A(n_548),
.Y(n_634)
);

OR2x6_ASAP7_75t_L g635 ( 
.A(n_524),
.B(n_499),
.Y(n_635)
);

NAND3xp33_ASAP7_75t_L g636 ( 
.A(n_586),
.B(n_489),
.C(n_487),
.Y(n_636)
);

NAND2xp5_ASAP7_75t_SL g637 ( 
.A(n_524),
.B(n_490),
.Y(n_637)
);

INVx3_ASAP7_75t_L g638 ( 
.A(n_544),
.Y(n_638)
);

INVx2_ASAP7_75t_L g639 ( 
.A(n_548),
.Y(n_639)
);

NOR2xp33_ASAP7_75t_L g640 ( 
.A(n_518),
.B(n_491),
.Y(n_640)
);

INVx2_ASAP7_75t_L g641 ( 
.A(n_548),
.Y(n_641)
);

INVx5_ASAP7_75t_L g642 ( 
.A(n_513),
.Y(n_642)
);

INVx3_ASAP7_75t_L g643 ( 
.A(n_544),
.Y(n_643)
);

OR2x6_ASAP7_75t_L g644 ( 
.A(n_579),
.B(n_500),
.Y(n_644)
);

AND3x2_ASAP7_75t_L g645 ( 
.A(n_535),
.B(n_476),
.C(n_411),
.Y(n_645)
);

AOI22xp33_ASAP7_75t_L g646 ( 
.A1(n_579),
.A2(n_278),
.B1(n_306),
.B2(n_280),
.Y(n_646)
);

INVx2_ASAP7_75t_L g647 ( 
.A(n_560),
.Y(n_647)
);

BUFx2_ASAP7_75t_L g648 ( 
.A(n_535),
.Y(n_648)
);

INVx2_ASAP7_75t_L g649 ( 
.A(n_560),
.Y(n_649)
);

INVx1_ASAP7_75t_L g650 ( 
.A(n_517),
.Y(n_650)
);

NAND2xp5_ASAP7_75t_L g651 ( 
.A(n_508),
.B(n_495),
.Y(n_651)
);

INVx2_ASAP7_75t_SL g652 ( 
.A(n_508),
.Y(n_652)
);

CKINVDCx20_ASAP7_75t_R g653 ( 
.A(n_519),
.Y(n_653)
);

INVx1_ASAP7_75t_L g654 ( 
.A(n_520),
.Y(n_654)
);

NAND2xp5_ASAP7_75t_SL g655 ( 
.A(n_508),
.B(n_498),
.Y(n_655)
);

NAND2xp5_ASAP7_75t_SL g656 ( 
.A(n_522),
.B(n_503),
.Y(n_656)
);

NOR2xp33_ASAP7_75t_L g657 ( 
.A(n_531),
.B(n_506),
.Y(n_657)
);

INVx1_ASAP7_75t_L g658 ( 
.A(n_520),
.Y(n_658)
);

INVx1_ASAP7_75t_L g659 ( 
.A(n_525),
.Y(n_659)
);

INVx1_ASAP7_75t_L g660 ( 
.A(n_525),
.Y(n_660)
);

BUFx2_ASAP7_75t_L g661 ( 
.A(n_541),
.Y(n_661)
);

BUFx3_ASAP7_75t_L g662 ( 
.A(n_516),
.Y(n_662)
);

NAND2xp5_ASAP7_75t_L g663 ( 
.A(n_522),
.B(n_500),
.Y(n_663)
);

BUFx3_ASAP7_75t_L g664 ( 
.A(n_516),
.Y(n_664)
);

NAND2xp5_ASAP7_75t_L g665 ( 
.A(n_522),
.B(n_496),
.Y(n_665)
);

NAND2xp5_ASAP7_75t_SL g666 ( 
.A(n_584),
.B(n_415),
.Y(n_666)
);

INVx2_ASAP7_75t_SL g667 ( 
.A(n_579),
.Y(n_667)
);

OR2x2_ASAP7_75t_L g668 ( 
.A(n_541),
.B(n_434),
.Y(n_668)
);

INVx1_ASAP7_75t_L g669 ( 
.A(n_527),
.Y(n_669)
);

INVx1_ASAP7_75t_SL g670 ( 
.A(n_577),
.Y(n_670)
);

CKINVDCx5p33_ASAP7_75t_R g671 ( 
.A(n_516),
.Y(n_671)
);

NAND3xp33_ASAP7_75t_L g672 ( 
.A(n_586),
.B(n_315),
.C(n_309),
.Y(n_672)
);

BUFx3_ASAP7_75t_L g673 ( 
.A(n_516),
.Y(n_673)
);

INVx1_ASAP7_75t_L g674 ( 
.A(n_527),
.Y(n_674)
);

NOR2xp33_ASAP7_75t_L g675 ( 
.A(n_546),
.B(n_419),
.Y(n_675)
);

INVx2_ASAP7_75t_SL g676 ( 
.A(n_579),
.Y(n_676)
);

BUFx3_ASAP7_75t_L g677 ( 
.A(n_584),
.Y(n_677)
);

BUFx6f_ASAP7_75t_L g678 ( 
.A(n_580),
.Y(n_678)
);

INVx1_ASAP7_75t_L g679 ( 
.A(n_529),
.Y(n_679)
);

INVx2_ASAP7_75t_L g680 ( 
.A(n_560),
.Y(n_680)
);

INVx1_ASAP7_75t_L g681 ( 
.A(n_529),
.Y(n_681)
);

BUFx3_ASAP7_75t_L g682 ( 
.A(n_584),
.Y(n_682)
);

AND2x2_ASAP7_75t_SL g683 ( 
.A(n_534),
.B(n_259),
.Y(n_683)
);

AO21x2_ASAP7_75t_L g684 ( 
.A1(n_521),
.A2(n_287),
.B(n_274),
.Y(n_684)
);

AOI22xp33_ASAP7_75t_L g685 ( 
.A1(n_565),
.A2(n_352),
.B1(n_330),
.B2(n_337),
.Y(n_685)
);

INVx2_ASAP7_75t_L g686 ( 
.A(n_563),
.Y(n_686)
);

INVx2_ASAP7_75t_L g687 ( 
.A(n_563),
.Y(n_687)
);

INVx1_ASAP7_75t_L g688 ( 
.A(n_530),
.Y(n_688)
);

NAND2xp5_ASAP7_75t_L g689 ( 
.A(n_528),
.B(n_420),
.Y(n_689)
);

OAI22xp5_ASAP7_75t_L g690 ( 
.A1(n_558),
.A2(n_373),
.B1(n_245),
.B2(n_251),
.Y(n_690)
);

AND2x2_ASAP7_75t_L g691 ( 
.A(n_532),
.B(n_459),
.Y(n_691)
);

INVx1_ASAP7_75t_L g692 ( 
.A(n_530),
.Y(n_692)
);

AND2x4_ASAP7_75t_L g693 ( 
.A(n_565),
.B(n_460),
.Y(n_693)
);

INVx2_ASAP7_75t_L g694 ( 
.A(n_563),
.Y(n_694)
);

INVx5_ASAP7_75t_L g695 ( 
.A(n_513),
.Y(n_695)
);

INVx1_ASAP7_75t_L g696 ( 
.A(n_538),
.Y(n_696)
);

INVx1_ASAP7_75t_L g697 ( 
.A(n_538),
.Y(n_697)
);

NAND2xp33_ASAP7_75t_L g698 ( 
.A(n_587),
.B(n_211),
.Y(n_698)
);

NAND2xp5_ASAP7_75t_SL g699 ( 
.A(n_573),
.B(n_438),
.Y(n_699)
);

INVx4_ASAP7_75t_L g700 ( 
.A(n_533),
.Y(n_700)
);

INVx1_ASAP7_75t_L g701 ( 
.A(n_543),
.Y(n_701)
);

BUFx2_ASAP7_75t_L g702 ( 
.A(n_573),
.Y(n_702)
);

NAND2xp5_ASAP7_75t_SL g703 ( 
.A(n_565),
.B(n_532),
.Y(n_703)
);

AND2x4_ASAP7_75t_L g704 ( 
.A(n_565),
.B(n_460),
.Y(n_704)
);

BUFx6f_ASAP7_75t_L g705 ( 
.A(n_580),
.Y(n_705)
);

NAND2xp5_ASAP7_75t_L g706 ( 
.A(n_528),
.B(n_536),
.Y(n_706)
);

INVx2_ASAP7_75t_L g707 ( 
.A(n_568),
.Y(n_707)
);

AND2x2_ASAP7_75t_L g708 ( 
.A(n_532),
.B(n_461),
.Y(n_708)
);

HB1xp67_ASAP7_75t_L g709 ( 
.A(n_536),
.Y(n_709)
);

INVx1_ASAP7_75t_L g710 ( 
.A(n_543),
.Y(n_710)
);

INVx1_ASAP7_75t_L g711 ( 
.A(n_550),
.Y(n_711)
);

CKINVDCx5p33_ASAP7_75t_R g712 ( 
.A(n_580),
.Y(n_712)
);

INVx3_ASAP7_75t_L g713 ( 
.A(n_544),
.Y(n_713)
);

NOR2xp33_ASAP7_75t_L g714 ( 
.A(n_521),
.B(n_416),
.Y(n_714)
);

NAND2xp33_ASAP7_75t_L g715 ( 
.A(n_587),
.B(n_212),
.Y(n_715)
);

BUFx6f_ASAP7_75t_L g716 ( 
.A(n_580),
.Y(n_716)
);

NAND2xp5_ASAP7_75t_SL g717 ( 
.A(n_536),
.B(n_440),
.Y(n_717)
);

OR2x6_ASAP7_75t_L g718 ( 
.A(n_536),
.B(n_461),
.Y(n_718)
);

INVx1_ASAP7_75t_L g719 ( 
.A(n_550),
.Y(n_719)
);

INVx1_ASAP7_75t_L g720 ( 
.A(n_551),
.Y(n_720)
);

OR2x6_ASAP7_75t_L g721 ( 
.A(n_547),
.B(n_319),
.Y(n_721)
);

INVx1_ASAP7_75t_L g722 ( 
.A(n_551),
.Y(n_722)
);

INVx2_ASAP7_75t_L g723 ( 
.A(n_568),
.Y(n_723)
);

INVx1_ASAP7_75t_L g724 ( 
.A(n_553),
.Y(n_724)
);

INVx1_ASAP7_75t_L g725 ( 
.A(n_553),
.Y(n_725)
);

AND2x6_ASAP7_75t_L g726 ( 
.A(n_511),
.B(n_539),
.Y(n_726)
);

NAND2xp5_ASAP7_75t_L g727 ( 
.A(n_528),
.B(n_230),
.Y(n_727)
);

INVx2_ASAP7_75t_L g728 ( 
.A(n_568),
.Y(n_728)
);

INVx2_ASAP7_75t_L g729 ( 
.A(n_569),
.Y(n_729)
);

NOR2xp33_ASAP7_75t_L g730 ( 
.A(n_576),
.B(n_422),
.Y(n_730)
);

INVx2_ASAP7_75t_L g731 ( 
.A(n_569),
.Y(n_731)
);

BUFx6f_ASAP7_75t_L g732 ( 
.A(n_580),
.Y(n_732)
);

INVx3_ASAP7_75t_L g733 ( 
.A(n_544),
.Y(n_733)
);

INVx2_ASAP7_75t_L g734 ( 
.A(n_569),
.Y(n_734)
);

INVx2_ASAP7_75t_L g735 ( 
.A(n_544),
.Y(n_735)
);

OAI21xp33_ASAP7_75t_L g736 ( 
.A1(n_576),
.A2(n_355),
.B(n_340),
.Y(n_736)
);

NAND2xp5_ASAP7_75t_L g737 ( 
.A(n_528),
.B(n_288),
.Y(n_737)
);

INVxp67_ASAP7_75t_SL g738 ( 
.A(n_547),
.Y(n_738)
);

BUFx8_ASAP7_75t_SL g739 ( 
.A(n_587),
.Y(n_739)
);

INVxp67_ASAP7_75t_L g740 ( 
.A(n_648),
.Y(n_740)
);

BUFx6f_ASAP7_75t_L g741 ( 
.A(n_682),
.Y(n_741)
);

INVx1_ASAP7_75t_L g742 ( 
.A(n_615),
.Y(n_742)
);

NAND2xp5_ASAP7_75t_SL g743 ( 
.A(n_628),
.B(n_483),
.Y(n_743)
);

NAND2xp5_ASAP7_75t_SL g744 ( 
.A(n_683),
.B(n_212),
.Y(n_744)
);

NAND2xp5_ASAP7_75t_L g745 ( 
.A(n_738),
.B(n_587),
.Y(n_745)
);

INVx1_ASAP7_75t_L g746 ( 
.A(n_624),
.Y(n_746)
);

NAND2xp5_ASAP7_75t_SL g747 ( 
.A(n_683),
.B(n_220),
.Y(n_747)
);

INVx2_ASAP7_75t_L g748 ( 
.A(n_620),
.Y(n_748)
);

NAND2xp5_ASAP7_75t_L g749 ( 
.A(n_626),
.B(n_511),
.Y(n_749)
);

O2A1O1Ixp5_ASAP7_75t_L g750 ( 
.A1(n_591),
.A2(n_583),
.B(n_581),
.C(n_574),
.Y(n_750)
);

BUFx5_ASAP7_75t_L g751 ( 
.A(n_591),
.Y(n_751)
);

NAND2xp5_ASAP7_75t_L g752 ( 
.A(n_627),
.B(n_539),
.Y(n_752)
);

INVx3_ASAP7_75t_L g753 ( 
.A(n_682),
.Y(n_753)
);

INVx2_ASAP7_75t_L g754 ( 
.A(n_621),
.Y(n_754)
);

AOI22xp5_ASAP7_75t_L g755 ( 
.A1(n_600),
.A2(n_493),
.B1(n_501),
.B2(n_502),
.Y(n_755)
);

AOI22xp5_ASAP7_75t_L g756 ( 
.A1(n_600),
.A2(n_504),
.B1(n_220),
.B2(n_347),
.Y(n_756)
);

INVx8_ASAP7_75t_L g757 ( 
.A(n_606),
.Y(n_757)
);

HB1xp67_ASAP7_75t_L g758 ( 
.A(n_596),
.Y(n_758)
);

INVxp67_ASAP7_75t_L g759 ( 
.A(n_648),
.Y(n_759)
);

NAND2xp5_ASAP7_75t_SL g760 ( 
.A(n_683),
.B(n_225),
.Y(n_760)
);

AND2x4_ASAP7_75t_L g761 ( 
.A(n_677),
.B(n_428),
.Y(n_761)
);

OAI22xp33_ASAP7_75t_L g762 ( 
.A1(n_702),
.A2(n_554),
.B1(n_571),
.B2(n_574),
.Y(n_762)
);

AO22x2_ASAP7_75t_L g763 ( 
.A1(n_636),
.A2(n_583),
.B1(n_581),
.B2(n_431),
.Y(n_763)
);

NOR2xp33_ASAP7_75t_L g764 ( 
.A(n_651),
.B(n_554),
.Y(n_764)
);

AOI22xp5_ASAP7_75t_L g765 ( 
.A1(n_600),
.A2(n_250),
.B1(n_347),
.B2(n_249),
.Y(n_765)
);

AND2x2_ASAP7_75t_L g766 ( 
.A(n_661),
.B(n_408),
.Y(n_766)
);

INVx8_ASAP7_75t_L g767 ( 
.A(n_606),
.Y(n_767)
);

BUFx6f_ASAP7_75t_L g768 ( 
.A(n_682),
.Y(n_768)
);

NAND2xp33_ASAP7_75t_L g769 ( 
.A(n_630),
.B(n_225),
.Y(n_769)
);

AND2x2_ASAP7_75t_L g770 ( 
.A(n_661),
.B(n_470),
.Y(n_770)
);

INVxp67_ASAP7_75t_SL g771 ( 
.A(n_677),
.Y(n_771)
);

INVx2_ASAP7_75t_SL g772 ( 
.A(n_668),
.Y(n_772)
);

AND2x2_ASAP7_75t_L g773 ( 
.A(n_596),
.B(n_472),
.Y(n_773)
);

INVxp67_ASAP7_75t_L g774 ( 
.A(n_616),
.Y(n_774)
);

INVx2_ASAP7_75t_SL g775 ( 
.A(n_668),
.Y(n_775)
);

NAND2xp5_ASAP7_75t_L g776 ( 
.A(n_652),
.B(n_580),
.Y(n_776)
);

NAND2xp5_ASAP7_75t_SL g777 ( 
.A(n_652),
.B(n_227),
.Y(n_777)
);

NAND2xp5_ASAP7_75t_L g778 ( 
.A(n_667),
.B(n_582),
.Y(n_778)
);

NAND2xp33_ASAP7_75t_L g779 ( 
.A(n_633),
.B(n_227),
.Y(n_779)
);

NAND2xp5_ASAP7_75t_SL g780 ( 
.A(n_590),
.B(n_233),
.Y(n_780)
);

AOI21xp5_ASAP7_75t_L g781 ( 
.A1(n_663),
.A2(n_571),
.B(n_515),
.Y(n_781)
);

INVx1_ASAP7_75t_L g782 ( 
.A(n_650),
.Y(n_782)
);

AOI22xp33_ASAP7_75t_L g783 ( 
.A1(n_702),
.A2(n_582),
.B1(n_578),
.B2(n_557),
.Y(n_783)
);

INVx1_ASAP7_75t_L g784 ( 
.A(n_654),
.Y(n_784)
);

AOI22xp5_ASAP7_75t_L g785 ( 
.A1(n_667),
.A2(n_249),
.B1(n_250),
.B2(n_401),
.Y(n_785)
);

INVx1_ASAP7_75t_L g786 ( 
.A(n_654),
.Y(n_786)
);

NAND2xp5_ASAP7_75t_L g787 ( 
.A(n_676),
.B(n_582),
.Y(n_787)
);

NAND2xp5_ASAP7_75t_SL g788 ( 
.A(n_592),
.B(n_233),
.Y(n_788)
);

NAND2xp5_ASAP7_75t_L g789 ( 
.A(n_676),
.B(n_582),
.Y(n_789)
);

BUFx2_ASAP7_75t_L g790 ( 
.A(n_653),
.Y(n_790)
);

NAND2xp33_ASAP7_75t_L g791 ( 
.A(n_604),
.B(n_238),
.Y(n_791)
);

HB1xp67_ASAP7_75t_L g792 ( 
.A(n_618),
.Y(n_792)
);

NAND2xp5_ASAP7_75t_L g793 ( 
.A(n_640),
.B(n_582),
.Y(n_793)
);

OR2x2_ASAP7_75t_L g794 ( 
.A(n_599),
.B(n_480),
.Y(n_794)
);

INVx1_ASAP7_75t_L g795 ( 
.A(n_658),
.Y(n_795)
);

AND2x2_ASAP7_75t_L g796 ( 
.A(n_623),
.B(n_481),
.Y(n_796)
);

NAND2xp5_ASAP7_75t_L g797 ( 
.A(n_598),
.B(n_582),
.Y(n_797)
);

AOI22xp5_ASAP7_75t_L g798 ( 
.A1(n_635),
.A2(n_303),
.B1(n_247),
.B2(n_401),
.Y(n_798)
);

INVx1_ASAP7_75t_L g799 ( 
.A(n_658),
.Y(n_799)
);

INVx2_ASAP7_75t_SL g800 ( 
.A(n_599),
.Y(n_800)
);

AOI22xp33_ASAP7_75t_L g801 ( 
.A1(n_602),
.A2(n_578),
.B1(n_557),
.B2(n_570),
.Y(n_801)
);

BUFx5_ASAP7_75t_L g802 ( 
.A(n_612),
.Y(n_802)
);

OR2x2_ASAP7_75t_L g803 ( 
.A(n_670),
.B(n_251),
.Y(n_803)
);

NAND2xp5_ASAP7_75t_SL g804 ( 
.A(n_595),
.B(n_238),
.Y(n_804)
);

AND2x4_ASAP7_75t_L g805 ( 
.A(n_635),
.B(n_644),
.Y(n_805)
);

NAND2x1p5_ASAP7_75t_L g806 ( 
.A(n_664),
.B(n_533),
.Y(n_806)
);

AO221x1_ASAP7_75t_L g807 ( 
.A1(n_690),
.A2(n_399),
.B1(n_259),
.B2(n_298),
.C(n_299),
.Y(n_807)
);

INVx2_ASAP7_75t_L g808 ( 
.A(n_622),
.Y(n_808)
);

AOI22x1_ASAP7_75t_L g809 ( 
.A1(n_589),
.A2(n_561),
.B1(n_564),
.B2(n_566),
.Y(n_809)
);

NOR3xp33_ASAP7_75t_L g810 ( 
.A(n_655),
.B(n_350),
.C(n_349),
.Y(n_810)
);

NAND2xp5_ASAP7_75t_L g811 ( 
.A(n_598),
.B(n_578),
.Y(n_811)
);

AOI22xp5_ASAP7_75t_L g812 ( 
.A1(n_635),
.A2(n_357),
.B1(n_239),
.B2(n_246),
.Y(n_812)
);

NAND2xp5_ASAP7_75t_SL g813 ( 
.A(n_595),
.B(n_239),
.Y(n_813)
);

INVx2_ASAP7_75t_L g814 ( 
.A(n_625),
.Y(n_814)
);

INVx4_ASAP7_75t_L g815 ( 
.A(n_618),
.Y(n_815)
);

BUFx3_ASAP7_75t_L g816 ( 
.A(n_623),
.Y(n_816)
);

INVx2_ASAP7_75t_L g817 ( 
.A(n_625),
.Y(n_817)
);

INVx1_ASAP7_75t_L g818 ( 
.A(n_659),
.Y(n_818)
);

INVx3_ASAP7_75t_L g819 ( 
.A(n_605),
.Y(n_819)
);

AOI22xp5_ASAP7_75t_L g820 ( 
.A1(n_635),
.A2(n_357),
.B1(n_246),
.B2(n_247),
.Y(n_820)
);

INVx1_ASAP7_75t_L g821 ( 
.A(n_659),
.Y(n_821)
);

INVx2_ASAP7_75t_L g822 ( 
.A(n_629),
.Y(n_822)
);

INVx1_ASAP7_75t_L g823 ( 
.A(n_660),
.Y(n_823)
);

NAND2xp5_ASAP7_75t_SL g824 ( 
.A(n_657),
.B(n_303),
.Y(n_824)
);

INVx2_ASAP7_75t_L g825 ( 
.A(n_629),
.Y(n_825)
);

AOI22xp5_ASAP7_75t_L g826 ( 
.A1(n_635),
.A2(n_606),
.B1(n_644),
.B2(n_597),
.Y(n_826)
);

INVx2_ASAP7_75t_SL g827 ( 
.A(n_645),
.Y(n_827)
);

O2A1O1Ixp33_ASAP7_75t_L g828 ( 
.A1(n_703),
.A2(n_570),
.B(n_566),
.C(n_564),
.Y(n_828)
);

AOI22xp33_ASAP7_75t_L g829 ( 
.A1(n_721),
.A2(n_322),
.B1(n_334),
.B2(n_348),
.Y(n_829)
);

AOI22xp5_ASAP7_75t_L g830 ( 
.A1(n_606),
.A2(n_377),
.B1(n_378),
.B2(n_387),
.Y(n_830)
);

NAND2xp5_ASAP7_75t_SL g831 ( 
.A(n_665),
.B(n_377),
.Y(n_831)
);

NAND2xp5_ASAP7_75t_SL g832 ( 
.A(n_597),
.B(n_378),
.Y(n_832)
);

INVx1_ASAP7_75t_L g833 ( 
.A(n_660),
.Y(n_833)
);

AND2x2_ASAP7_75t_L g834 ( 
.A(n_714),
.B(n_353),
.Y(n_834)
);

BUFx4f_ASAP7_75t_L g835 ( 
.A(n_606),
.Y(n_835)
);

NAND2xp5_ASAP7_75t_SL g836 ( 
.A(n_595),
.B(n_387),
.Y(n_836)
);

INVx2_ASAP7_75t_SL g837 ( 
.A(n_691),
.Y(n_837)
);

NAND2xp5_ASAP7_75t_L g838 ( 
.A(n_606),
.B(n_721),
.Y(n_838)
);

NOR2xp33_ASAP7_75t_L g839 ( 
.A(n_656),
.B(n_349),
.Y(n_839)
);

NAND2xp5_ASAP7_75t_L g840 ( 
.A(n_606),
.B(n_291),
.Y(n_840)
);

AOI22xp5_ASAP7_75t_L g841 ( 
.A1(n_644),
.A2(n_393),
.B1(n_395),
.B2(n_400),
.Y(n_841)
);

NOR2xp33_ASAP7_75t_L g842 ( 
.A(n_601),
.B(n_350),
.Y(n_842)
);

NAND2xp5_ASAP7_75t_L g843 ( 
.A(n_721),
.B(n_367),
.Y(n_843)
);

INVx1_ASAP7_75t_L g844 ( 
.A(n_669),
.Y(n_844)
);

INVx2_ASAP7_75t_SL g845 ( 
.A(n_691),
.Y(n_845)
);

NAND2xp5_ASAP7_75t_SL g846 ( 
.A(n_607),
.B(n_393),
.Y(n_846)
);

NAND2xp5_ASAP7_75t_L g847 ( 
.A(n_721),
.B(n_372),
.Y(n_847)
);

NAND2xp5_ASAP7_75t_L g848 ( 
.A(n_721),
.B(n_395),
.Y(n_848)
);

NAND2xp5_ASAP7_75t_SL g849 ( 
.A(n_611),
.B(n_400),
.Y(n_849)
);

NOR3xp33_ASAP7_75t_L g850 ( 
.A(n_637),
.B(n_375),
.C(n_359),
.Y(n_850)
);

NAND2xp5_ASAP7_75t_SL g851 ( 
.A(n_611),
.B(n_359),
.Y(n_851)
);

NAND2x1_ASAP7_75t_L g852 ( 
.A(n_605),
.B(n_510),
.Y(n_852)
);

INVx2_ASAP7_75t_L g853 ( 
.A(n_631),
.Y(n_853)
);

AOI22xp5_ASAP7_75t_L g854 ( 
.A1(n_644),
.A2(n_293),
.B1(n_292),
.B2(n_304),
.Y(n_854)
);

NOR2xp33_ASAP7_75t_L g855 ( 
.A(n_709),
.B(n_689),
.Y(n_855)
);

AOI22xp5_ASAP7_75t_L g856 ( 
.A1(n_644),
.A2(n_305),
.B1(n_310),
.B2(n_312),
.Y(n_856)
);

INVx2_ASAP7_75t_L g857 ( 
.A(n_631),
.Y(n_857)
);

INVx1_ASAP7_75t_L g858 ( 
.A(n_669),
.Y(n_858)
);

INVx2_ASAP7_75t_L g859 ( 
.A(n_634),
.Y(n_859)
);

INVx4_ASAP7_75t_L g860 ( 
.A(n_618),
.Y(n_860)
);

OAI22xp33_ASAP7_75t_L g861 ( 
.A1(n_718),
.A2(n_375),
.B1(n_360),
.B2(n_365),
.Y(n_861)
);

OR2x2_ASAP7_75t_L g862 ( 
.A(n_730),
.B(n_360),
.Y(n_862)
);

NAND2xp5_ASAP7_75t_L g863 ( 
.A(n_693),
.B(n_533),
.Y(n_863)
);

INVx1_ASAP7_75t_L g864 ( 
.A(n_674),
.Y(n_864)
);

NAND2xp5_ASAP7_75t_L g865 ( 
.A(n_693),
.B(n_704),
.Y(n_865)
);

NOR2xp67_ASAP7_75t_L g866 ( 
.A(n_675),
.B(n_533),
.Y(n_866)
);

NAND2xp5_ASAP7_75t_L g867 ( 
.A(n_693),
.B(n_533),
.Y(n_867)
);

NAND3xp33_ASAP7_75t_L g868 ( 
.A(n_593),
.B(n_376),
.C(n_369),
.Y(n_868)
);

INVx2_ASAP7_75t_L g869 ( 
.A(n_634),
.Y(n_869)
);

NAND2xp5_ASAP7_75t_SL g870 ( 
.A(n_607),
.B(n_313),
.Y(n_870)
);

NAND2xp5_ASAP7_75t_SL g871 ( 
.A(n_671),
.B(n_369),
.Y(n_871)
);

BUFx2_ASAP7_75t_L g872 ( 
.A(n_739),
.Y(n_872)
);

NAND2xp5_ASAP7_75t_L g873 ( 
.A(n_693),
.B(n_533),
.Y(n_873)
);

NOR2xp33_ASAP7_75t_L g874 ( 
.A(n_666),
.B(n_370),
.Y(n_874)
);

OR2x2_ASAP7_75t_L g875 ( 
.A(n_699),
.B(n_708),
.Y(n_875)
);

INVxp33_ASAP7_75t_L g876 ( 
.A(n_708),
.Y(n_876)
);

AND2x2_ASAP7_75t_L g877 ( 
.A(n_613),
.B(n_358),
.Y(n_877)
);

NOR2xp33_ASAP7_75t_L g878 ( 
.A(n_618),
.B(n_370),
.Y(n_878)
);

NAND2xp5_ASAP7_75t_L g879 ( 
.A(n_704),
.B(n_533),
.Y(n_879)
);

NOR2xp33_ASAP7_75t_L g880 ( 
.A(n_618),
.B(n_374),
.Y(n_880)
);

NAND2xp5_ASAP7_75t_L g881 ( 
.A(n_704),
.B(n_374),
.Y(n_881)
);

NAND2xp5_ASAP7_75t_L g882 ( 
.A(n_706),
.B(n_727),
.Y(n_882)
);

INVx1_ASAP7_75t_L g883 ( 
.A(n_674),
.Y(n_883)
);

NAND2xp5_ASAP7_75t_L g884 ( 
.A(n_737),
.B(n_376),
.Y(n_884)
);

NAND2xp5_ASAP7_75t_L g885 ( 
.A(n_605),
.B(n_379),
.Y(n_885)
);

AOI22xp5_ASAP7_75t_SL g886 ( 
.A1(n_671),
.A2(n_381),
.B1(n_382),
.B2(n_398),
.Y(n_886)
);

INVx2_ASAP7_75t_SL g887 ( 
.A(n_717),
.Y(n_887)
);

INVx2_ASAP7_75t_L g888 ( 
.A(n_639),
.Y(n_888)
);

NOR2xp33_ASAP7_75t_L g889 ( 
.A(n_718),
.B(n_379),
.Y(n_889)
);

NOR2xp33_ASAP7_75t_L g890 ( 
.A(n_718),
.B(n_380),
.Y(n_890)
);

AOI22xp33_ASAP7_75t_L g891 ( 
.A1(n_607),
.A2(n_322),
.B1(n_334),
.B2(n_348),
.Y(n_891)
);

NAND2xp5_ASAP7_75t_L g892 ( 
.A(n_617),
.B(n_380),
.Y(n_892)
);

INVx1_ASAP7_75t_L g893 ( 
.A(n_679),
.Y(n_893)
);

INVxp67_ASAP7_75t_L g894 ( 
.A(n_718),
.Y(n_894)
);

NAND2xp5_ASAP7_75t_L g895 ( 
.A(n_617),
.B(n_381),
.Y(n_895)
);

INVx2_ASAP7_75t_L g896 ( 
.A(n_639),
.Y(n_896)
);

NAND2xp5_ASAP7_75t_SL g897 ( 
.A(n_678),
.B(n_321),
.Y(n_897)
);

NOR2xp33_ASAP7_75t_L g898 ( 
.A(n_718),
.B(n_382),
.Y(n_898)
);

NAND2xp5_ASAP7_75t_L g899 ( 
.A(n_617),
.B(n_389),
.Y(n_899)
);

INVx2_ASAP7_75t_L g900 ( 
.A(n_641),
.Y(n_900)
);

INVx2_ASAP7_75t_L g901 ( 
.A(n_641),
.Y(n_901)
);

AOI22xp33_ASAP7_75t_L g902 ( 
.A1(n_736),
.A2(n_348),
.B1(n_334),
.B2(n_358),
.Y(n_902)
);

NAND2xp5_ASAP7_75t_L g903 ( 
.A(n_764),
.B(n_774),
.Y(n_903)
);

NAND2xp5_ASAP7_75t_L g904 ( 
.A(n_764),
.B(n_646),
.Y(n_904)
);

NAND2xp5_ASAP7_75t_L g905 ( 
.A(n_774),
.B(n_685),
.Y(n_905)
);

INVxp67_ASAP7_75t_L g906 ( 
.A(n_758),
.Y(n_906)
);

AND2x4_ASAP7_75t_L g907 ( 
.A(n_805),
.B(n_662),
.Y(n_907)
);

O2A1O1Ixp33_ASAP7_75t_L g908 ( 
.A1(n_861),
.A2(n_698),
.B(n_715),
.C(n_594),
.Y(n_908)
);

INVx4_ASAP7_75t_L g909 ( 
.A(n_805),
.Y(n_909)
);

NAND2xp5_ASAP7_75t_L g910 ( 
.A(n_762),
.B(n_712),
.Y(n_910)
);

OA22x2_ASAP7_75t_L g911 ( 
.A1(n_756),
.A2(n_736),
.B1(n_608),
.B2(n_390),
.Y(n_911)
);

AOI21xp5_ASAP7_75t_L g912 ( 
.A1(n_793),
.A2(n_614),
.B(n_612),
.Y(n_912)
);

AOI21xp5_ASAP7_75t_L g913 ( 
.A1(n_745),
.A2(n_614),
.B(n_594),
.Y(n_913)
);

AND2x4_ASAP7_75t_L g914 ( 
.A(n_894),
.B(n_662),
.Y(n_914)
);

NAND2xp5_ASAP7_75t_L g915 ( 
.A(n_762),
.B(n_712),
.Y(n_915)
);

AND2x2_ASAP7_75t_L g916 ( 
.A(n_740),
.B(n_673),
.Y(n_916)
);

INVx2_ASAP7_75t_L g917 ( 
.A(n_748),
.Y(n_917)
);

O2A1O1Ixp33_ASAP7_75t_L g918 ( 
.A1(n_861),
.A2(n_603),
.B(n_609),
.C(n_610),
.Y(n_918)
);

NOR3xp33_ASAP7_75t_L g919 ( 
.A(n_740),
.B(n_390),
.C(n_389),
.Y(n_919)
);

OAI21xp5_ASAP7_75t_L g920 ( 
.A1(n_750),
.A2(n_636),
.B(n_608),
.Y(n_920)
);

NAND2xp5_ASAP7_75t_L g921 ( 
.A(n_855),
.B(n_726),
.Y(n_921)
);

AOI21x1_ASAP7_75t_L g922 ( 
.A1(n_870),
.A2(n_681),
.B(n_679),
.Y(n_922)
);

AO21x1_ASAP7_75t_L g923 ( 
.A1(n_744),
.A2(n_608),
.B(n_681),
.Y(n_923)
);

AOI22xp33_ASAP7_75t_L g924 ( 
.A1(n_744),
.A2(n_684),
.B1(n_672),
.B2(n_726),
.Y(n_924)
);

NOR2x1p5_ASAP7_75t_L g925 ( 
.A(n_816),
.B(n_673),
.Y(n_925)
);

NAND2xp5_ASAP7_75t_L g926 ( 
.A(n_855),
.B(n_726),
.Y(n_926)
);

INVx3_ASAP7_75t_L g927 ( 
.A(n_815),
.Y(n_927)
);

INVx1_ASAP7_75t_L g928 ( 
.A(n_742),
.Y(n_928)
);

AOI22xp5_ASAP7_75t_L g929 ( 
.A1(n_771),
.A2(n_726),
.B1(n_724),
.B2(n_688),
.Y(n_929)
);

INVx3_ASAP7_75t_L g930 ( 
.A(n_815),
.Y(n_930)
);

OAI21xp5_ASAP7_75t_L g931 ( 
.A1(n_781),
.A2(n_870),
.B(n_813),
.Y(n_931)
);

NAND2xp5_ASAP7_75t_L g932 ( 
.A(n_882),
.B(n_726),
.Y(n_932)
);

NAND2xp5_ASAP7_75t_L g933 ( 
.A(n_771),
.B(n_726),
.Y(n_933)
);

NOR2xp33_ASAP7_75t_L g934 ( 
.A(n_876),
.B(n_608),
.Y(n_934)
);

NOR2xp33_ASAP7_75t_L g935 ( 
.A(n_772),
.B(n_589),
.Y(n_935)
);

NAND2xp5_ASAP7_75t_L g936 ( 
.A(n_834),
.B(n_726),
.Y(n_936)
);

NAND2xp5_ASAP7_75t_L g937 ( 
.A(n_837),
.B(n_845),
.Y(n_937)
);

CKINVDCx10_ASAP7_75t_R g938 ( 
.A(n_790),
.Y(n_938)
);

AOI21xp5_ASAP7_75t_L g939 ( 
.A1(n_804),
.A2(n_609),
.B(n_603),
.Y(n_939)
);

AOI21xp5_ASAP7_75t_L g940 ( 
.A1(n_804),
.A2(n_619),
.B(n_610),
.Y(n_940)
);

AOI21xp5_ASAP7_75t_L g941 ( 
.A1(n_813),
.A2(n_619),
.B(n_688),
.Y(n_941)
);

AOI21xp5_ASAP7_75t_L g942 ( 
.A1(n_836),
.A2(n_696),
.B(n_692),
.Y(n_942)
);

AND2x2_ASAP7_75t_L g943 ( 
.A(n_759),
.B(n_766),
.Y(n_943)
);

CKINVDCx20_ASAP7_75t_R g944 ( 
.A(n_872),
.Y(n_944)
);

NAND2xp5_ASAP7_75t_L g945 ( 
.A(n_865),
.B(n_684),
.Y(n_945)
);

CKINVDCx10_ASAP7_75t_R g946 ( 
.A(n_794),
.Y(n_946)
);

NOR2xp33_ASAP7_75t_L g947 ( 
.A(n_775),
.B(n_692),
.Y(n_947)
);

AOI21xp5_ASAP7_75t_L g948 ( 
.A1(n_836),
.A2(n_697),
.B(n_696),
.Y(n_948)
);

NAND2xp5_ASAP7_75t_L g949 ( 
.A(n_878),
.B(n_684),
.Y(n_949)
);

AND2x2_ASAP7_75t_L g950 ( 
.A(n_759),
.B(n_358),
.Y(n_950)
);

NAND2xp5_ASAP7_75t_L g951 ( 
.A(n_878),
.B(n_664),
.Y(n_951)
);

NAND2xp5_ASAP7_75t_SL g952 ( 
.A(n_826),
.B(n_751),
.Y(n_952)
);

A2O1A1Ixp33_ASAP7_75t_L g953 ( 
.A1(n_746),
.A2(n_719),
.B(n_697),
.C(n_701),
.Y(n_953)
);

NAND2xp5_ASAP7_75t_L g954 ( 
.A(n_880),
.B(n_664),
.Y(n_954)
);

AOI21xp5_ASAP7_75t_L g955 ( 
.A1(n_846),
.A2(n_710),
.B(n_701),
.Y(n_955)
);

AOI21xp5_ASAP7_75t_L g956 ( 
.A1(n_846),
.A2(n_711),
.B(n_710),
.Y(n_956)
);

AOI21xp5_ASAP7_75t_L g957 ( 
.A1(n_778),
.A2(n_719),
.B(n_711),
.Y(n_957)
);

NAND2xp5_ASAP7_75t_L g958 ( 
.A(n_880),
.B(n_720),
.Y(n_958)
);

NOR2xp33_ASAP7_75t_L g959 ( 
.A(n_875),
.B(n_720),
.Y(n_959)
);

OAI21xp33_ASAP7_75t_L g960 ( 
.A1(n_862),
.A2(n_398),
.B(n_722),
.Y(n_960)
);

AO21x1_ASAP7_75t_L g961 ( 
.A1(n_747),
.A2(n_725),
.B(n_722),
.Y(n_961)
);

NOR2xp33_ASAP7_75t_L g962 ( 
.A(n_743),
.B(n_724),
.Y(n_962)
);

OAI21xp5_ASAP7_75t_L g963 ( 
.A1(n_787),
.A2(n_672),
.B(n_725),
.Y(n_963)
);

OAI21xp5_ASAP7_75t_L g964 ( 
.A1(n_789),
.A2(n_735),
.B(n_638),
.Y(n_964)
);

HB1xp67_ASAP7_75t_L g965 ( 
.A(n_758),
.Y(n_965)
);

AOI21xp5_ASAP7_75t_L g966 ( 
.A1(n_776),
.A2(n_643),
.B(n_632),
.Y(n_966)
);

NOR2xp33_ASAP7_75t_L g967 ( 
.A(n_780),
.B(n_632),
.Y(n_967)
);

AOI21xp5_ASAP7_75t_L g968 ( 
.A1(n_797),
.A2(n_643),
.B(n_632),
.Y(n_968)
);

NAND2xp5_ASAP7_75t_L g969 ( 
.A(n_783),
.B(n_647),
.Y(n_969)
);

INVx2_ASAP7_75t_L g970 ( 
.A(n_754),
.Y(n_970)
);

AOI21xp5_ASAP7_75t_L g971 ( 
.A1(n_852),
.A2(n_643),
.B(n_638),
.Y(n_971)
);

AOI21xp5_ASAP7_75t_L g972 ( 
.A1(n_749),
.A2(n_638),
.B(n_713),
.Y(n_972)
);

INVx1_ASAP7_75t_L g973 ( 
.A(n_782),
.Y(n_973)
);

HB1xp67_ASAP7_75t_L g974 ( 
.A(n_792),
.Y(n_974)
);

NOR2xp33_ASAP7_75t_L g975 ( 
.A(n_780),
.B(n_713),
.Y(n_975)
);

NAND2xp5_ASAP7_75t_L g976 ( 
.A(n_783),
.B(n_647),
.Y(n_976)
);

BUFx12f_ASAP7_75t_L g977 ( 
.A(n_761),
.Y(n_977)
);

AOI21xp5_ASAP7_75t_L g978 ( 
.A1(n_752),
.A2(n_713),
.B(n_733),
.Y(n_978)
);

AOI21xp5_ASAP7_75t_L g979 ( 
.A1(n_784),
.A2(n_733),
.B(n_735),
.Y(n_979)
);

AOI21xp5_ASAP7_75t_L g980 ( 
.A1(n_786),
.A2(n_733),
.B(n_678),
.Y(n_980)
);

AOI21xp5_ASAP7_75t_L g981 ( 
.A1(n_795),
.A2(n_705),
.B(n_732),
.Y(n_981)
);

NAND2xp5_ASAP7_75t_L g982 ( 
.A(n_753),
.B(n_649),
.Y(n_982)
);

AOI21xp5_ASAP7_75t_L g983 ( 
.A1(n_799),
.A2(n_705),
.B(n_732),
.Y(n_983)
);

AND2x2_ASAP7_75t_L g984 ( 
.A(n_800),
.B(n_649),
.Y(n_984)
);

AOI21xp5_ASAP7_75t_L g985 ( 
.A1(n_818),
.A2(n_823),
.B(n_821),
.Y(n_985)
);

INVx2_ASAP7_75t_SL g986 ( 
.A(n_761),
.Y(n_986)
);

HB1xp67_ASAP7_75t_L g987 ( 
.A(n_792),
.Y(n_987)
);

INVx2_ASAP7_75t_L g988 ( 
.A(n_808),
.Y(n_988)
);

AOI21xp5_ASAP7_75t_L g989 ( 
.A1(n_833),
.A2(n_678),
.B(n_732),
.Y(n_989)
);

NAND2xp5_ASAP7_75t_L g990 ( 
.A(n_753),
.B(n_734),
.Y(n_990)
);

NAND2xp5_ASAP7_75t_L g991 ( 
.A(n_843),
.B(n_847),
.Y(n_991)
);

AOI21xp5_ASAP7_75t_L g992 ( 
.A1(n_844),
.A2(n_678),
.B(n_732),
.Y(n_992)
);

NAND2xp5_ASAP7_75t_SL g993 ( 
.A(n_751),
.B(n_678),
.Y(n_993)
);

NAND2xp5_ASAP7_75t_L g994 ( 
.A(n_858),
.B(n_680),
.Y(n_994)
);

AOI21xp33_ASAP7_75t_L g995 ( 
.A1(n_891),
.A2(n_734),
.B(n_686),
.Y(n_995)
);

O2A1O1Ixp33_ASAP7_75t_L g996 ( 
.A1(n_788),
.A2(n_731),
.B(n_729),
.C(n_728),
.Y(n_996)
);

NAND2xp5_ASAP7_75t_L g997 ( 
.A(n_864),
.B(n_680),
.Y(n_997)
);

CKINVDCx5p33_ASAP7_75t_R g998 ( 
.A(n_796),
.Y(n_998)
);

NOR2xp33_ASAP7_75t_L g999 ( 
.A(n_894),
.B(n_705),
.Y(n_999)
);

BUFx10_ASAP7_75t_L g1000 ( 
.A(n_889),
.Y(n_1000)
);

AND2x2_ASAP7_75t_L g1001 ( 
.A(n_770),
.B(n_686),
.Y(n_1001)
);

OAI22xp5_ASAP7_75t_L g1002 ( 
.A1(n_883),
.A2(n_732),
.B1(n_716),
.B2(n_705),
.Y(n_1002)
);

OAI21xp33_ASAP7_75t_L g1003 ( 
.A1(n_785),
.A2(n_842),
.B(n_812),
.Y(n_1003)
);

OAI321xp33_ASAP7_75t_L g1004 ( 
.A1(n_829),
.A2(n_891),
.A3(n_902),
.B1(n_868),
.B2(n_747),
.C(n_760),
.Y(n_1004)
);

OAI22xp5_ASAP7_75t_L g1005 ( 
.A1(n_893),
.A2(n_741),
.B1(n_768),
.B2(n_765),
.Y(n_1005)
);

NAND2xp5_ASAP7_75t_L g1006 ( 
.A(n_877),
.B(n_687),
.Y(n_1006)
);

NAND2xp5_ASAP7_75t_L g1007 ( 
.A(n_801),
.B(n_687),
.Y(n_1007)
);

AO21x1_ASAP7_75t_L g1008 ( 
.A1(n_760),
.A2(n_731),
.B(n_729),
.Y(n_1008)
);

BUFx6f_ASAP7_75t_L g1009 ( 
.A(n_741),
.Y(n_1009)
);

INVx2_ASAP7_75t_L g1010 ( 
.A(n_814),
.Y(n_1010)
);

NAND2xp5_ASAP7_75t_SL g1011 ( 
.A(n_751),
.B(n_705),
.Y(n_1011)
);

NAND2x1p5_ASAP7_75t_L g1012 ( 
.A(n_860),
.B(n_741),
.Y(n_1012)
);

AOI21xp5_ASAP7_75t_L g1013 ( 
.A1(n_811),
.A2(n_716),
.B(n_723),
.Y(n_1013)
);

BUFx3_ASAP7_75t_L g1014 ( 
.A(n_741),
.Y(n_1014)
);

NAND2xp5_ASAP7_75t_L g1015 ( 
.A(n_801),
.B(n_694),
.Y(n_1015)
);

NAND2xp5_ASAP7_75t_L g1016 ( 
.A(n_889),
.B(n_694),
.Y(n_1016)
);

NOR2xp33_ASAP7_75t_L g1017 ( 
.A(n_832),
.B(n_716),
.Y(n_1017)
);

NOR2xp33_ASAP7_75t_L g1018 ( 
.A(n_768),
.B(n_716),
.Y(n_1018)
);

NAND2xp5_ASAP7_75t_L g1019 ( 
.A(n_890),
.B(n_728),
.Y(n_1019)
);

INVx1_ASAP7_75t_L g1020 ( 
.A(n_828),
.Y(n_1020)
);

AOI21xp5_ASAP7_75t_L g1021 ( 
.A1(n_863),
.A2(n_873),
.B(n_867),
.Y(n_1021)
);

NAND2xp5_ASAP7_75t_L g1022 ( 
.A(n_890),
.B(n_898),
.Y(n_1022)
);

AOI21xp5_ASAP7_75t_L g1023 ( 
.A1(n_879),
.A2(n_716),
.B(n_723),
.Y(n_1023)
);

INVx4_ASAP7_75t_L g1024 ( 
.A(n_860),
.Y(n_1024)
);

NAND2xp5_ASAP7_75t_L g1025 ( 
.A(n_898),
.B(n_707),
.Y(n_1025)
);

AND2x2_ASAP7_75t_L g1026 ( 
.A(n_773),
.B(n_707),
.Y(n_1026)
);

NAND2xp5_ASAP7_75t_SL g1027 ( 
.A(n_751),
.B(n_642),
.Y(n_1027)
);

AOI21x1_ASAP7_75t_L g1028 ( 
.A1(n_897),
.A2(n_509),
.B(n_515),
.Y(n_1028)
);

NAND2xp5_ASAP7_75t_L g1029 ( 
.A(n_829),
.B(n_324),
.Y(n_1029)
);

AOI21xp5_ASAP7_75t_L g1030 ( 
.A1(n_819),
.A2(n_700),
.B(n_695),
.Y(n_1030)
);

OR2x6_ASAP7_75t_L g1031 ( 
.A(n_757),
.B(n_700),
.Y(n_1031)
);

INVx1_ASAP7_75t_L g1032 ( 
.A(n_817),
.Y(n_1032)
);

AOI21xp5_ASAP7_75t_L g1033 ( 
.A1(n_819),
.A2(n_700),
.B(n_695),
.Y(n_1033)
);

INVx1_ASAP7_75t_L g1034 ( 
.A(n_822),
.Y(n_1034)
);

O2A1O1Ixp33_ASAP7_75t_L g1035 ( 
.A1(n_777),
.A2(n_363),
.B(n_335),
.C(n_332),
.Y(n_1035)
);

OAI21xp5_ASAP7_75t_L g1036 ( 
.A1(n_809),
.A2(n_700),
.B(n_695),
.Y(n_1036)
);

INVxp67_ASAP7_75t_SL g1037 ( 
.A(n_768),
.Y(n_1037)
);

INVx2_ASAP7_75t_L g1038 ( 
.A(n_825),
.Y(n_1038)
);

OAI21x1_ASAP7_75t_L g1039 ( 
.A1(n_853),
.A2(n_859),
.B(n_857),
.Y(n_1039)
);

AOI21x1_ASAP7_75t_L g1040 ( 
.A1(n_897),
.A2(n_888),
.B(n_869),
.Y(n_1040)
);

NAND2xp5_ASAP7_75t_SL g1041 ( 
.A(n_751),
.B(n_802),
.Y(n_1041)
);

NAND2xp5_ASAP7_75t_L g1042 ( 
.A(n_884),
.B(n_768),
.Y(n_1042)
);

OAI22xp5_ASAP7_75t_L g1043 ( 
.A1(n_798),
.A2(n_385),
.B1(n_386),
.B2(n_388),
.Y(n_1043)
);

AOI21xp5_ASAP7_75t_L g1044 ( 
.A1(n_885),
.A2(n_695),
.B(n_642),
.Y(n_1044)
);

NAND2xp5_ASAP7_75t_L g1045 ( 
.A(n_848),
.B(n_325),
.Y(n_1045)
);

AOI21xp5_ASAP7_75t_L g1046 ( 
.A1(n_892),
.A2(n_695),
.B(n_642),
.Y(n_1046)
);

NAND2xp5_ASAP7_75t_L g1047 ( 
.A(n_895),
.B(n_327),
.Y(n_1047)
);

AOI21xp5_ASAP7_75t_L g1048 ( 
.A1(n_899),
.A2(n_695),
.B(n_642),
.Y(n_1048)
);

INVx1_ASAP7_75t_L g1049 ( 
.A(n_896),
.Y(n_1049)
);

A2O1A1Ixp33_ASAP7_75t_L g1050 ( 
.A1(n_839),
.A2(n_842),
.B(n_874),
.C(n_854),
.Y(n_1050)
);

NAND2xp5_ASAP7_75t_SL g1051 ( 
.A(n_751),
.B(n_642),
.Y(n_1051)
);

NAND2xp5_ASAP7_75t_SL g1052 ( 
.A(n_802),
.B(n_642),
.Y(n_1052)
);

OAI21xp5_ASAP7_75t_L g1053 ( 
.A1(n_900),
.A2(n_510),
.B(n_346),
.Y(n_1053)
);

NAND2xp5_ASAP7_75t_SL g1054 ( 
.A(n_802),
.B(n_559),
.Y(n_1054)
);

INVx2_ASAP7_75t_L g1055 ( 
.A(n_901),
.Y(n_1055)
);

AOI21xp5_ASAP7_75t_L g1056 ( 
.A1(n_831),
.A2(n_509),
.B(n_515),
.Y(n_1056)
);

NAND2xp5_ASAP7_75t_L g1057 ( 
.A(n_902),
.B(n_344),
.Y(n_1057)
);

OAI21xp5_ASAP7_75t_L g1058 ( 
.A1(n_769),
.A2(n_510),
.B(n_394),
.Y(n_1058)
);

AOI21xp5_ASAP7_75t_L g1059 ( 
.A1(n_791),
.A2(n_509),
.B(n_523),
.Y(n_1059)
);

OAI21xp5_ASAP7_75t_L g1060 ( 
.A1(n_779),
.A2(n_510),
.B(n_396),
.Y(n_1060)
);

AOI21xp5_ASAP7_75t_L g1061 ( 
.A1(n_824),
.A2(n_523),
.B(n_263),
.Y(n_1061)
);

INVx2_ASAP7_75t_L g1062 ( 
.A(n_802),
.Y(n_1062)
);

AOI21xp5_ASAP7_75t_L g1063 ( 
.A1(n_881),
.A2(n_523),
.B(n_266),
.Y(n_1063)
);

NAND2xp5_ASAP7_75t_L g1064 ( 
.A(n_856),
.B(n_351),
.Y(n_1064)
);

O2A1O1Ixp5_ASAP7_75t_L g1065 ( 
.A1(n_839),
.A2(n_575),
.B(n_572),
.C(n_559),
.Y(n_1065)
);

NAND2xp5_ASAP7_75t_L g1066 ( 
.A(n_874),
.B(n_559),
.Y(n_1066)
);

NAND2xp5_ASAP7_75t_L g1067 ( 
.A(n_820),
.B(n_559),
.Y(n_1067)
);

NAND2xp5_ASAP7_75t_L g1068 ( 
.A(n_841),
.B(n_559),
.Y(n_1068)
);

AOI21xp5_ASAP7_75t_L g1069 ( 
.A1(n_866),
.A2(n_308),
.B(n_267),
.Y(n_1069)
);

OAI21xp5_ASAP7_75t_L g1070 ( 
.A1(n_835),
.A2(n_323),
.B(n_268),
.Y(n_1070)
);

OAI22xp5_ASAP7_75t_L g1071 ( 
.A1(n_838),
.A2(n_575),
.B1(n_572),
.B2(n_559),
.Y(n_1071)
);

NAND2xp5_ASAP7_75t_SL g1072 ( 
.A(n_802),
.B(n_572),
.Y(n_1072)
);

INVx2_ASAP7_75t_L g1073 ( 
.A(n_802),
.Y(n_1073)
);

NAND2xp5_ASAP7_75t_L g1074 ( 
.A(n_763),
.B(n_572),
.Y(n_1074)
);

AOI21xp5_ASAP7_75t_L g1075 ( 
.A1(n_835),
.A2(n_307),
.B(n_271),
.Y(n_1075)
);

BUFx4f_ASAP7_75t_L g1076 ( 
.A(n_827),
.Y(n_1076)
);

INVx1_ASAP7_75t_L g1077 ( 
.A(n_763),
.Y(n_1077)
);

OAI21xp33_ASAP7_75t_L g1078 ( 
.A1(n_850),
.A2(n_328),
.B(n_281),
.Y(n_1078)
);

AOI22xp33_ASAP7_75t_L g1079 ( 
.A1(n_807),
.A2(n_575),
.B1(n_572),
.B2(n_259),
.Y(n_1079)
);

INVx1_ASAP7_75t_SL g1080 ( 
.A(n_803),
.Y(n_1080)
);

BUFx12f_ASAP7_75t_L g1081 ( 
.A(n_887),
.Y(n_1081)
);

AND2x2_ASAP7_75t_L g1082 ( 
.A(n_886),
.B(n_572),
.Y(n_1082)
);

AOI21xp5_ASAP7_75t_L g1083 ( 
.A1(n_757),
.A2(n_329),
.B(n_289),
.Y(n_1083)
);

CKINVDCx5p33_ASAP7_75t_R g1084 ( 
.A(n_755),
.Y(n_1084)
);

INVx1_ASAP7_75t_L g1085 ( 
.A(n_763),
.Y(n_1085)
);

AOI21xp5_ASAP7_75t_L g1086 ( 
.A1(n_757),
.A2(n_331),
.B(n_290),
.Y(n_1086)
);

NAND2xp5_ASAP7_75t_L g1087 ( 
.A(n_810),
.B(n_575),
.Y(n_1087)
);

AOI22xp5_ASAP7_75t_L g1088 ( 
.A1(n_1003),
.A2(n_810),
.B1(n_850),
.B2(n_851),
.Y(n_1088)
);

INVx1_ASAP7_75t_L g1089 ( 
.A(n_928),
.Y(n_1089)
);

NAND2xp5_ASAP7_75t_SL g1090 ( 
.A(n_921),
.B(n_830),
.Y(n_1090)
);

O2A1O1Ixp33_ASAP7_75t_L g1091 ( 
.A1(n_1050),
.A2(n_849),
.B(n_871),
.C(n_840),
.Y(n_1091)
);

BUFx2_ASAP7_75t_L g1092 ( 
.A(n_998),
.Y(n_1092)
);

NAND2xp5_ASAP7_75t_SL g1093 ( 
.A(n_926),
.B(n_767),
.Y(n_1093)
);

AOI21xp5_ASAP7_75t_L g1094 ( 
.A1(n_912),
.A2(n_767),
.B(n_806),
.Y(n_1094)
);

AOI21xp5_ASAP7_75t_L g1095 ( 
.A1(n_1041),
.A2(n_767),
.B(n_806),
.Y(n_1095)
);

NOR2xp33_ASAP7_75t_L g1096 ( 
.A(n_903),
.B(n_14),
.Y(n_1096)
);

A2O1A1Ixp33_ASAP7_75t_L g1097 ( 
.A1(n_1050),
.A2(n_575),
.B(n_341),
.C(n_403),
.Y(n_1097)
);

CKINVDCx5p33_ASAP7_75t_R g1098 ( 
.A(n_938),
.Y(n_1098)
);

INVxp67_ASAP7_75t_L g1099 ( 
.A(n_965),
.Y(n_1099)
);

NAND2xp5_ASAP7_75t_SL g1100 ( 
.A(n_1022),
.B(n_575),
.Y(n_1100)
);

AOI22xp5_ASAP7_75t_L g1101 ( 
.A1(n_943),
.A2(n_962),
.B1(n_904),
.B2(n_1084),
.Y(n_1101)
);

AOI221x1_ASAP7_75t_L g1102 ( 
.A1(n_910),
.A2(n_513),
.B1(n_298),
.B2(n_17),
.C(n_18),
.Y(n_1102)
);

HB1xp67_ASAP7_75t_L g1103 ( 
.A(n_965),
.Y(n_1103)
);

XOR2xp5_ASAP7_75t_L g1104 ( 
.A(n_944),
.B(n_345),
.Y(n_1104)
);

NAND3xp33_ASAP7_75t_SL g1105 ( 
.A(n_960),
.B(n_343),
.C(n_297),
.Y(n_1105)
);

O2A1O1Ixp5_ASAP7_75t_L g1106 ( 
.A1(n_931),
.A2(n_15),
.B(n_16),
.C(n_17),
.Y(n_1106)
);

BUFx12f_ASAP7_75t_L g1107 ( 
.A(n_977),
.Y(n_1107)
);

OAI22xp5_ASAP7_75t_L g1108 ( 
.A1(n_958),
.A2(n_295),
.B1(n_282),
.B2(n_298),
.Y(n_1108)
);

A2O1A1Ixp33_ASAP7_75t_L g1109 ( 
.A1(n_915),
.A2(n_298),
.B(n_513),
.C(n_25),
.Y(n_1109)
);

BUFx2_ASAP7_75t_L g1110 ( 
.A(n_906),
.Y(n_1110)
);

AOI21xp5_ASAP7_75t_L g1111 ( 
.A1(n_993),
.A2(n_513),
.B(n_202),
.Y(n_1111)
);

NAND3xp33_ASAP7_75t_SL g1112 ( 
.A(n_1078),
.B(n_1043),
.C(n_919),
.Y(n_1112)
);

AOI22xp5_ASAP7_75t_L g1113 ( 
.A1(n_947),
.A2(n_19),
.B1(n_22),
.B2(n_25),
.Y(n_1113)
);

BUFx6f_ASAP7_75t_L g1114 ( 
.A(n_909),
.Y(n_1114)
);

OAI22xp5_ASAP7_75t_L g1115 ( 
.A1(n_959),
.A2(n_19),
.B1(n_28),
.B2(n_32),
.Y(n_1115)
);

AOI21xp5_ASAP7_75t_L g1116 ( 
.A1(n_993),
.A2(n_1011),
.B(n_1054),
.Y(n_1116)
);

HB1xp67_ASAP7_75t_L g1117 ( 
.A(n_974),
.Y(n_1117)
);

INVx6_ASAP7_75t_L g1118 ( 
.A(n_907),
.Y(n_1118)
);

NAND2xp5_ASAP7_75t_L g1119 ( 
.A(n_959),
.B(n_37),
.Y(n_1119)
);

NOR2xp33_ASAP7_75t_L g1120 ( 
.A(n_991),
.B(n_38),
.Y(n_1120)
);

AND2x2_ASAP7_75t_L g1121 ( 
.A(n_1080),
.B(n_38),
.Y(n_1121)
);

AOI21xp5_ASAP7_75t_L g1122 ( 
.A1(n_1011),
.A2(n_77),
.B(n_190),
.Y(n_1122)
);

AOI21x1_ASAP7_75t_L g1123 ( 
.A1(n_949),
.A2(n_201),
.B(n_189),
.Y(n_1123)
);

INVx4_ASAP7_75t_L g1124 ( 
.A(n_907),
.Y(n_1124)
);

NAND2xp5_ASAP7_75t_L g1125 ( 
.A(n_947),
.B(n_41),
.Y(n_1125)
);

NAND2xp5_ASAP7_75t_L g1126 ( 
.A(n_905),
.B(n_42),
.Y(n_1126)
);

BUFx6f_ASAP7_75t_L g1127 ( 
.A(n_1009),
.Y(n_1127)
);

BUFx6f_ASAP7_75t_L g1128 ( 
.A(n_1009),
.Y(n_1128)
);

NAND2xp5_ASAP7_75t_SL g1129 ( 
.A(n_916),
.B(n_46),
.Y(n_1129)
);

BUFx6f_ASAP7_75t_L g1130 ( 
.A(n_1009),
.Y(n_1130)
);

AOI21x1_ASAP7_75t_L g1131 ( 
.A1(n_922),
.A2(n_1028),
.B(n_1008),
.Y(n_1131)
);

AOI22xp5_ASAP7_75t_L g1132 ( 
.A1(n_936),
.A2(n_49),
.B1(n_50),
.B2(n_51),
.Y(n_1132)
);

AOI22xp5_ASAP7_75t_L g1133 ( 
.A1(n_934),
.A2(n_49),
.B1(n_50),
.B2(n_53),
.Y(n_1133)
);

BUFx2_ASAP7_75t_L g1134 ( 
.A(n_986),
.Y(n_1134)
);

AND2x4_ASAP7_75t_L g1135 ( 
.A(n_914),
.B(n_53),
.Y(n_1135)
);

AOI22xp5_ASAP7_75t_L g1136 ( 
.A1(n_934),
.A2(n_54),
.B1(n_55),
.B2(n_56),
.Y(n_1136)
);

AND2x2_ASAP7_75t_L g1137 ( 
.A(n_1026),
.B(n_54),
.Y(n_1137)
);

BUFx2_ASAP7_75t_SL g1138 ( 
.A(n_925),
.Y(n_1138)
);

INVx2_ASAP7_75t_L g1139 ( 
.A(n_970),
.Y(n_1139)
);

NAND2xp5_ASAP7_75t_L g1140 ( 
.A(n_1001),
.B(n_55),
.Y(n_1140)
);

NOR3xp33_ASAP7_75t_SL g1141 ( 
.A(n_953),
.B(n_56),
.C(n_61),
.Y(n_1141)
);

INVx1_ASAP7_75t_L g1142 ( 
.A(n_973),
.Y(n_1142)
);

NAND2xp5_ASAP7_75t_L g1143 ( 
.A(n_974),
.B(n_61),
.Y(n_1143)
);

OAI22xp5_ASAP7_75t_L g1144 ( 
.A1(n_929),
.A2(n_64),
.B1(n_67),
.B2(n_68),
.Y(n_1144)
);

AOI21xp5_ASAP7_75t_L g1145 ( 
.A1(n_1054),
.A2(n_124),
.B(n_180),
.Y(n_1145)
);

OAI21xp5_ASAP7_75t_L g1146 ( 
.A1(n_942),
.A2(n_64),
.B(n_68),
.Y(n_1146)
);

BUFx3_ASAP7_75t_L g1147 ( 
.A(n_1076),
.Y(n_1147)
);

AOI22xp33_ASAP7_75t_L g1148 ( 
.A1(n_911),
.A2(n_69),
.B1(n_70),
.B2(n_71),
.Y(n_1148)
);

INVxp67_ASAP7_75t_L g1149 ( 
.A(n_987),
.Y(n_1149)
);

AND2x2_ASAP7_75t_L g1150 ( 
.A(n_950),
.B(n_70),
.Y(n_1150)
);

NAND2xp5_ASAP7_75t_L g1151 ( 
.A(n_987),
.B(n_71),
.Y(n_1151)
);

NAND2xp5_ASAP7_75t_L g1152 ( 
.A(n_984),
.B(n_72),
.Y(n_1152)
);

AOI21xp5_ASAP7_75t_L g1153 ( 
.A1(n_1072),
.A2(n_78),
.B(n_85),
.Y(n_1153)
);

A2O1A1Ixp33_ASAP7_75t_L g1154 ( 
.A1(n_1004),
.A2(n_908),
.B(n_985),
.C(n_1035),
.Y(n_1154)
);

NAND2xp5_ASAP7_75t_SL g1155 ( 
.A(n_952),
.B(n_103),
.Y(n_1155)
);

NOR3xp33_ASAP7_75t_SL g1156 ( 
.A(n_953),
.B(n_955),
.C(n_948),
.Y(n_1156)
);

NAND2xp5_ASAP7_75t_SL g1157 ( 
.A(n_952),
.B(n_114),
.Y(n_1157)
);

NAND2xp5_ASAP7_75t_L g1158 ( 
.A(n_935),
.B(n_137),
.Y(n_1158)
);

BUFx3_ASAP7_75t_L g1159 ( 
.A(n_1081),
.Y(n_1159)
);

OAI21xp33_ASAP7_75t_L g1160 ( 
.A1(n_935),
.A2(n_153),
.B(n_158),
.Y(n_1160)
);

NOR2xp67_ASAP7_75t_L g1161 ( 
.A(n_937),
.B(n_169),
.Y(n_1161)
);

AOI21xp5_ASAP7_75t_L g1162 ( 
.A1(n_1072),
.A2(n_173),
.B(n_174),
.Y(n_1162)
);

NOR2xp33_ASAP7_75t_L g1163 ( 
.A(n_1000),
.B(n_932),
.Y(n_1163)
);

CKINVDCx20_ASAP7_75t_R g1164 ( 
.A(n_1000),
.Y(n_1164)
);

AND2x2_ASAP7_75t_L g1165 ( 
.A(n_914),
.B(n_177),
.Y(n_1165)
);

HB1xp67_ASAP7_75t_L g1166 ( 
.A(n_933),
.Y(n_1166)
);

NOR2xp33_ASAP7_75t_R g1167 ( 
.A(n_946),
.B(n_185),
.Y(n_1167)
);

OAI21xp5_ASAP7_75t_L g1168 ( 
.A1(n_956),
.A2(n_941),
.B(n_920),
.Y(n_1168)
);

A2O1A1Ixp33_ASAP7_75t_L g1169 ( 
.A1(n_967),
.A2(n_975),
.B(n_1025),
.C(n_1019),
.Y(n_1169)
);

NOR2xp33_ASAP7_75t_L g1170 ( 
.A(n_1042),
.B(n_1006),
.Y(n_1170)
);

AOI22xp33_ASAP7_75t_L g1171 ( 
.A1(n_911),
.A2(n_1029),
.B1(n_1057),
.B2(n_1085),
.Y(n_1171)
);

NAND2xp5_ASAP7_75t_L g1172 ( 
.A(n_927),
.B(n_930),
.Y(n_1172)
);

AOI21xp5_ASAP7_75t_L g1173 ( 
.A1(n_913),
.A2(n_1073),
.B(n_1062),
.Y(n_1173)
);

NAND2xp5_ASAP7_75t_SL g1174 ( 
.A(n_1009),
.B(n_1016),
.Y(n_1174)
);

NOR2x1_ASAP7_75t_L g1175 ( 
.A(n_1014),
.B(n_1024),
.Y(n_1175)
);

NAND2xp5_ASAP7_75t_L g1176 ( 
.A(n_927),
.B(n_930),
.Y(n_1176)
);

INVx3_ASAP7_75t_L g1177 ( 
.A(n_1024),
.Y(n_1177)
);

CKINVDCx8_ASAP7_75t_R g1178 ( 
.A(n_1031),
.Y(n_1178)
);

OAI22xp5_ASAP7_75t_L g1179 ( 
.A1(n_1020),
.A2(n_1005),
.B1(n_954),
.B2(n_951),
.Y(n_1179)
);

AOI21xp5_ASAP7_75t_L g1180 ( 
.A1(n_1062),
.A2(n_1073),
.B(n_1027),
.Y(n_1180)
);

NAND2xp5_ASAP7_75t_L g1181 ( 
.A(n_945),
.B(n_1045),
.Y(n_1181)
);

AOI21xp5_ASAP7_75t_L g1182 ( 
.A1(n_1027),
.A2(n_1051),
.B(n_1052),
.Y(n_1182)
);

NAND2xp5_ASAP7_75t_L g1183 ( 
.A(n_999),
.B(n_1064),
.Y(n_1183)
);

NOR2xp33_ASAP7_75t_R g1184 ( 
.A(n_1014),
.B(n_1018),
.Y(n_1184)
);

NOR2xp33_ASAP7_75t_L g1185 ( 
.A(n_1047),
.B(n_967),
.Y(n_1185)
);

AOI21xp5_ASAP7_75t_L g1186 ( 
.A1(n_1051),
.A2(n_1052),
.B(n_957),
.Y(n_1186)
);

OAI21xp5_ASAP7_75t_L g1187 ( 
.A1(n_1021),
.A2(n_963),
.B(n_918),
.Y(n_1187)
);

AOI21xp5_ASAP7_75t_L g1188 ( 
.A1(n_939),
.A2(n_940),
.B(n_1002),
.Y(n_1188)
);

NAND2xp5_ASAP7_75t_SL g1189 ( 
.A(n_999),
.B(n_1082),
.Y(n_1189)
);

NAND2xp5_ASAP7_75t_SL g1190 ( 
.A(n_1018),
.B(n_1066),
.Y(n_1190)
);

OAI22xp5_ASAP7_75t_L g1191 ( 
.A1(n_994),
.A2(n_997),
.B1(n_975),
.B2(n_1012),
.Y(n_1191)
);

NAND2xp5_ASAP7_75t_SL g1192 ( 
.A(n_961),
.B(n_1017),
.Y(n_1192)
);

NAND2xp5_ASAP7_75t_L g1193 ( 
.A(n_1007),
.B(n_1015),
.Y(n_1193)
);

A2O1A1Ixp33_ASAP7_75t_L g1194 ( 
.A1(n_1017),
.A2(n_1058),
.B(n_1060),
.C(n_996),
.Y(n_1194)
);

CKINVDCx6p67_ASAP7_75t_R g1195 ( 
.A(n_1031),
.Y(n_1195)
);

INVxp67_ASAP7_75t_SL g1196 ( 
.A(n_969),
.Y(n_1196)
);

INVx4_ASAP7_75t_L g1197 ( 
.A(n_1012),
.Y(n_1197)
);

INVx1_ASAP7_75t_SL g1198 ( 
.A(n_1077),
.Y(n_1198)
);

AOI21xp5_ASAP7_75t_L g1199 ( 
.A1(n_981),
.A2(n_992),
.B(n_989),
.Y(n_1199)
);

A2O1A1Ixp33_ASAP7_75t_L g1200 ( 
.A1(n_1087),
.A2(n_924),
.B(n_1065),
.C(n_1067),
.Y(n_1200)
);

NAND2xp5_ASAP7_75t_SL g1201 ( 
.A(n_1070),
.B(n_1086),
.Y(n_1201)
);

INVx4_ASAP7_75t_L g1202 ( 
.A(n_1031),
.Y(n_1202)
);

AOI21xp5_ASAP7_75t_L g1203 ( 
.A1(n_983),
.A2(n_979),
.B(n_978),
.Y(n_1203)
);

CKINVDCx20_ASAP7_75t_R g1204 ( 
.A(n_1074),
.Y(n_1204)
);

NOR2xp33_ASAP7_75t_L g1205 ( 
.A(n_1032),
.B(n_1049),
.Y(n_1205)
);

AOI21xp5_ASAP7_75t_L g1206 ( 
.A1(n_972),
.A2(n_980),
.B(n_1023),
.Y(n_1206)
);

INVx1_ASAP7_75t_SL g1207 ( 
.A(n_1034),
.Y(n_1207)
);

AND2x2_ASAP7_75t_L g1208 ( 
.A(n_988),
.B(n_1038),
.Y(n_1208)
);

AOI21xp5_ASAP7_75t_L g1209 ( 
.A1(n_966),
.A2(n_1044),
.B(n_1048),
.Y(n_1209)
);

NOR2x1_ASAP7_75t_L g1210 ( 
.A(n_1083),
.B(n_1075),
.Y(n_1210)
);

INVx1_ASAP7_75t_L g1211 ( 
.A(n_1010),
.Y(n_1211)
);

NAND2xp5_ASAP7_75t_L g1212 ( 
.A(n_1037),
.B(n_976),
.Y(n_1212)
);

AOI21xp5_ASAP7_75t_L g1213 ( 
.A1(n_1046),
.A2(n_968),
.B(n_1013),
.Y(n_1213)
);

NAND2xp5_ASAP7_75t_L g1214 ( 
.A(n_1010),
.B(n_1055),
.Y(n_1214)
);

AND2x2_ASAP7_75t_L g1215 ( 
.A(n_1038),
.B(n_1055),
.Y(n_1215)
);

NAND2xp5_ASAP7_75t_L g1216 ( 
.A(n_924),
.B(n_982),
.Y(n_1216)
);

INVx2_ASAP7_75t_L g1217 ( 
.A(n_1039),
.Y(n_1217)
);

NAND2xp33_ASAP7_75t_SL g1218 ( 
.A(n_990),
.B(n_1068),
.Y(n_1218)
);

INVxp67_ASAP7_75t_SL g1219 ( 
.A(n_1071),
.Y(n_1219)
);

HB1xp67_ASAP7_75t_L g1220 ( 
.A(n_964),
.Y(n_1220)
);

AOI22xp5_ASAP7_75t_L g1221 ( 
.A1(n_1079),
.A2(n_923),
.B1(n_1053),
.B2(n_995),
.Y(n_1221)
);

INVx2_ASAP7_75t_L g1222 ( 
.A(n_1040),
.Y(n_1222)
);

O2A1O1Ixp33_ASAP7_75t_SL g1223 ( 
.A1(n_1036),
.A2(n_971),
.B(n_1030),
.C(n_1033),
.Y(n_1223)
);

INVx2_ASAP7_75t_L g1224 ( 
.A(n_1056),
.Y(n_1224)
);

AND2x2_ASAP7_75t_L g1225 ( 
.A(n_1079),
.B(n_1061),
.Y(n_1225)
);

NOR3xp33_ASAP7_75t_SL g1226 ( 
.A(n_1063),
.B(n_1059),
.C(n_1069),
.Y(n_1226)
);

NAND3xp33_ASAP7_75t_SL g1227 ( 
.A(n_1050),
.B(n_555),
.C(n_540),
.Y(n_1227)
);

OR2x6_ASAP7_75t_L g1228 ( 
.A(n_909),
.B(n_805),
.Y(n_1228)
);

A2O1A1Ixp33_ASAP7_75t_SL g1229 ( 
.A1(n_931),
.A2(n_967),
.B(n_975),
.C(n_640),
.Y(n_1229)
);

NAND2xp5_ASAP7_75t_L g1230 ( 
.A(n_903),
.B(n_764),
.Y(n_1230)
);

INVx2_ASAP7_75t_L g1231 ( 
.A(n_917),
.Y(n_1231)
);

OAI22x1_ASAP7_75t_L g1232 ( 
.A1(n_1084),
.A2(n_756),
.B1(n_702),
.B2(n_597),
.Y(n_1232)
);

INVx1_ASAP7_75t_L g1233 ( 
.A(n_1089),
.Y(n_1233)
);

NAND2xp5_ASAP7_75t_L g1234 ( 
.A(n_1230),
.B(n_1096),
.Y(n_1234)
);

AOI21xp5_ASAP7_75t_L g1235 ( 
.A1(n_1187),
.A2(n_1213),
.B(n_1223),
.Y(n_1235)
);

BUFx3_ASAP7_75t_L g1236 ( 
.A(n_1107),
.Y(n_1236)
);

AND2x2_ASAP7_75t_L g1237 ( 
.A(n_1103),
.B(n_1101),
.Y(n_1237)
);

AOI21xp5_ASAP7_75t_L g1238 ( 
.A1(n_1206),
.A2(n_1218),
.B(n_1229),
.Y(n_1238)
);

AOI21xp5_ASAP7_75t_L g1239 ( 
.A1(n_1229),
.A2(n_1203),
.B(n_1173),
.Y(n_1239)
);

NOR2xp67_ASAP7_75t_L g1240 ( 
.A(n_1099),
.B(n_1149),
.Y(n_1240)
);

OAI21x1_ASAP7_75t_L g1241 ( 
.A1(n_1131),
.A2(n_1186),
.B(n_1168),
.Y(n_1241)
);

OAI22xp33_ASAP7_75t_L g1242 ( 
.A1(n_1088),
.A2(n_1119),
.B1(n_1232),
.B2(n_1113),
.Y(n_1242)
);

AOI21xp5_ASAP7_75t_L g1243 ( 
.A1(n_1179),
.A2(n_1201),
.B(n_1194),
.Y(n_1243)
);

O2A1O1Ixp33_ASAP7_75t_SL g1244 ( 
.A1(n_1096),
.A2(n_1125),
.B(n_1097),
.C(n_1146),
.Y(n_1244)
);

OAI22xp5_ASAP7_75t_L g1245 ( 
.A1(n_1120),
.A2(n_1185),
.B1(n_1141),
.B2(n_1219),
.Y(n_1245)
);

AOI31xp67_ASAP7_75t_L g1246 ( 
.A1(n_1224),
.A2(n_1100),
.A3(n_1157),
.B(n_1155),
.Y(n_1246)
);

BUFx10_ASAP7_75t_L g1247 ( 
.A(n_1098),
.Y(n_1247)
);

NAND2xp5_ASAP7_75t_SL g1248 ( 
.A(n_1185),
.B(n_1183),
.Y(n_1248)
);

AOI21xp5_ASAP7_75t_L g1249 ( 
.A1(n_1094),
.A2(n_1190),
.B(n_1219),
.Y(n_1249)
);

OAI21xp5_ASAP7_75t_L g1250 ( 
.A1(n_1154),
.A2(n_1169),
.B(n_1090),
.Y(n_1250)
);

NAND2xp5_ASAP7_75t_L g1251 ( 
.A(n_1181),
.B(n_1170),
.Y(n_1251)
);

INVx1_ASAP7_75t_SL g1252 ( 
.A(n_1110),
.Y(n_1252)
);

AND2x2_ASAP7_75t_SL g1253 ( 
.A(n_1148),
.B(n_1135),
.Y(n_1253)
);

OAI21x1_ASAP7_75t_L g1254 ( 
.A1(n_1116),
.A2(n_1180),
.B(n_1217),
.Y(n_1254)
);

INVx1_ASAP7_75t_SL g1255 ( 
.A(n_1118),
.Y(n_1255)
);

AOI21xp5_ASAP7_75t_L g1256 ( 
.A1(n_1190),
.A2(n_1100),
.B(n_1182),
.Y(n_1256)
);

NAND2xp5_ASAP7_75t_L g1257 ( 
.A(n_1099),
.B(n_1117),
.Y(n_1257)
);

BUFx12f_ASAP7_75t_L g1258 ( 
.A(n_1092),
.Y(n_1258)
);

AND2x4_ASAP7_75t_L g1259 ( 
.A(n_1228),
.B(n_1124),
.Y(n_1259)
);

AOI22xp33_ASAP7_75t_L g1260 ( 
.A1(n_1112),
.A2(n_1204),
.B1(n_1227),
.B2(n_1148),
.Y(n_1260)
);

AOI21xp5_ASAP7_75t_SL g1261 ( 
.A1(n_1158),
.A2(n_1170),
.B(n_1191),
.Y(n_1261)
);

AO21x2_ASAP7_75t_L g1262 ( 
.A1(n_1192),
.A2(n_1221),
.B(n_1200),
.Y(n_1262)
);

AO31x2_ASAP7_75t_L g1263 ( 
.A1(n_1222),
.A2(n_1193),
.A3(n_1216),
.B(n_1102),
.Y(n_1263)
);

NAND3x1_ASAP7_75t_L g1264 ( 
.A(n_1120),
.B(n_1133),
.C(n_1136),
.Y(n_1264)
);

OAI21x1_ASAP7_75t_L g1265 ( 
.A1(n_1123),
.A2(n_1174),
.B(n_1111),
.Y(n_1265)
);

BUFx3_ASAP7_75t_L g1266 ( 
.A(n_1159),
.Y(n_1266)
);

NOR2xp33_ASAP7_75t_L g1267 ( 
.A(n_1104),
.B(n_1149),
.Y(n_1267)
);

BUFx12f_ASAP7_75t_L g1268 ( 
.A(n_1147),
.Y(n_1268)
);

AO31x2_ASAP7_75t_L g1269 ( 
.A1(n_1212),
.A2(n_1109),
.A3(n_1211),
.B(n_1205),
.Y(n_1269)
);

AOI21xp5_ASAP7_75t_L g1270 ( 
.A1(n_1090),
.A2(n_1155),
.B(n_1157),
.Y(n_1270)
);

AOI21xp5_ASAP7_75t_L g1271 ( 
.A1(n_1095),
.A2(n_1196),
.B(n_1093),
.Y(n_1271)
);

NAND2xp5_ASAP7_75t_L g1272 ( 
.A(n_1207),
.B(n_1137),
.Y(n_1272)
);

OAI21xp33_ASAP7_75t_L g1273 ( 
.A1(n_1141),
.A2(n_1132),
.B(n_1126),
.Y(n_1273)
);

NOR2xp33_ASAP7_75t_SL g1274 ( 
.A(n_1178),
.B(n_1228),
.Y(n_1274)
);

AOI21xp5_ASAP7_75t_L g1275 ( 
.A1(n_1196),
.A2(n_1093),
.B(n_1174),
.Y(n_1275)
);

OAI21xp5_ASAP7_75t_L g1276 ( 
.A1(n_1220),
.A2(n_1091),
.B(n_1156),
.Y(n_1276)
);

BUFx10_ASAP7_75t_L g1277 ( 
.A(n_1135),
.Y(n_1277)
);

NAND2xp5_ASAP7_75t_L g1278 ( 
.A(n_1163),
.B(n_1166),
.Y(n_1278)
);

AND2x4_ASAP7_75t_L g1279 ( 
.A(n_1228),
.B(n_1114),
.Y(n_1279)
);

OA21x2_ASAP7_75t_L g1280 ( 
.A1(n_1192),
.A2(n_1156),
.B(n_1220),
.Y(n_1280)
);

NOR2xp33_ASAP7_75t_SL g1281 ( 
.A(n_1160),
.B(n_1202),
.Y(n_1281)
);

OAI21x1_ASAP7_75t_SL g1282 ( 
.A1(n_1172),
.A2(n_1176),
.B(n_1143),
.Y(n_1282)
);

OAI21xp5_ASAP7_75t_L g1283 ( 
.A1(n_1106),
.A2(n_1225),
.B(n_1163),
.Y(n_1283)
);

NAND2xp5_ASAP7_75t_L g1284 ( 
.A(n_1166),
.B(n_1208),
.Y(n_1284)
);

OR2x6_ASAP7_75t_L g1285 ( 
.A(n_1138),
.B(n_1118),
.Y(n_1285)
);

AND2x2_ASAP7_75t_L g1286 ( 
.A(n_1121),
.B(n_1150),
.Y(n_1286)
);

AOI21xp5_ASAP7_75t_L g1287 ( 
.A1(n_1210),
.A2(n_1122),
.B(n_1153),
.Y(n_1287)
);

AO31x2_ASAP7_75t_L g1288 ( 
.A1(n_1205),
.A2(n_1214),
.A3(n_1231),
.B(n_1139),
.Y(n_1288)
);

AND2x2_ASAP7_75t_L g1289 ( 
.A(n_1134),
.B(n_1118),
.Y(n_1289)
);

INVx4_ASAP7_75t_L g1290 ( 
.A(n_1114),
.Y(n_1290)
);

NOR2xp33_ASAP7_75t_L g1291 ( 
.A(n_1164),
.B(n_1151),
.Y(n_1291)
);

O2A1O1Ixp33_ASAP7_75t_SL g1292 ( 
.A1(n_1129),
.A2(n_1152),
.B(n_1105),
.C(n_1140),
.Y(n_1292)
);

AOI21xp5_ASAP7_75t_L g1293 ( 
.A1(n_1145),
.A2(n_1162),
.B(n_1108),
.Y(n_1293)
);

A2O1A1Ixp33_ASAP7_75t_L g1294 ( 
.A1(n_1161),
.A2(n_1189),
.B(n_1171),
.C(n_1142),
.Y(n_1294)
);

INVx1_ASAP7_75t_L g1295 ( 
.A(n_1215),
.Y(n_1295)
);

BUFx2_ASAP7_75t_L g1296 ( 
.A(n_1184),
.Y(n_1296)
);

OR2x2_ASAP7_75t_L g1297 ( 
.A(n_1165),
.B(n_1198),
.Y(n_1297)
);

OAI21x1_ASAP7_75t_L g1298 ( 
.A1(n_1175),
.A2(n_1171),
.B(n_1177),
.Y(n_1298)
);

INVx2_ASAP7_75t_L g1299 ( 
.A(n_1127),
.Y(n_1299)
);

INVx1_ASAP7_75t_L g1300 ( 
.A(n_1127),
.Y(n_1300)
);

AOI221x1_ASAP7_75t_L g1301 ( 
.A1(n_1202),
.A2(n_1197),
.B1(n_1127),
.B2(n_1128),
.C(n_1130),
.Y(n_1301)
);

OAI21x1_ASAP7_75t_L g1302 ( 
.A1(n_1177),
.A2(n_1226),
.B(n_1195),
.Y(n_1302)
);

O2A1O1Ixp33_ASAP7_75t_SL g1303 ( 
.A1(n_1184),
.A2(n_1226),
.B(n_1127),
.C(n_1128),
.Y(n_1303)
);

NAND2xp5_ASAP7_75t_L g1304 ( 
.A(n_1128),
.B(n_1130),
.Y(n_1304)
);

AOI21xp5_ASAP7_75t_L g1305 ( 
.A1(n_1130),
.A2(n_1114),
.B(n_1167),
.Y(n_1305)
);

NAND2xp5_ASAP7_75t_L g1306 ( 
.A(n_1167),
.B(n_1230),
.Y(n_1306)
);

INVx1_ASAP7_75t_L g1307 ( 
.A(n_1089),
.Y(n_1307)
);

OA21x2_ASAP7_75t_L g1308 ( 
.A1(n_1213),
.A2(n_1209),
.B(n_1168),
.Y(n_1308)
);

OAI22xp5_ASAP7_75t_L g1309 ( 
.A1(n_1230),
.A2(n_1022),
.B1(n_1096),
.B2(n_1050),
.Y(n_1309)
);

BUFx8_ASAP7_75t_L g1310 ( 
.A(n_1107),
.Y(n_1310)
);

INVx1_ASAP7_75t_L g1311 ( 
.A(n_1089),
.Y(n_1311)
);

OAI21xp5_ASAP7_75t_L g1312 ( 
.A1(n_1230),
.A2(n_1050),
.B(n_1154),
.Y(n_1312)
);

BUFx2_ASAP7_75t_L g1313 ( 
.A(n_1092),
.Y(n_1313)
);

AOI21xp5_ASAP7_75t_L g1314 ( 
.A1(n_1187),
.A2(n_1041),
.B(n_952),
.Y(n_1314)
);

NAND2xp5_ASAP7_75t_L g1315 ( 
.A(n_1230),
.B(n_903),
.Y(n_1315)
);

OAI21x1_ASAP7_75t_L g1316 ( 
.A1(n_1209),
.A2(n_1188),
.B(n_1199),
.Y(n_1316)
);

O2A1O1Ixp33_ASAP7_75t_L g1317 ( 
.A1(n_1227),
.A2(n_1050),
.B(n_633),
.C(n_630),
.Y(n_1317)
);

AND2x2_ASAP7_75t_L g1318 ( 
.A(n_1103),
.B(n_943),
.Y(n_1318)
);

NAND2xp5_ASAP7_75t_L g1319 ( 
.A(n_1230),
.B(n_903),
.Y(n_1319)
);

INVx1_ASAP7_75t_SL g1320 ( 
.A(n_1110),
.Y(n_1320)
);

AOI21xp5_ASAP7_75t_L g1321 ( 
.A1(n_1187),
.A2(n_1041),
.B(n_952),
.Y(n_1321)
);

AOI21xp5_ASAP7_75t_L g1322 ( 
.A1(n_1187),
.A2(n_1041),
.B(n_952),
.Y(n_1322)
);

OAI21xp5_ASAP7_75t_L g1323 ( 
.A1(n_1230),
.A2(n_1050),
.B(n_1154),
.Y(n_1323)
);

BUFx2_ASAP7_75t_L g1324 ( 
.A(n_1092),
.Y(n_1324)
);

AOI22xp5_ASAP7_75t_L g1325 ( 
.A1(n_1096),
.A2(n_611),
.B1(n_770),
.B2(n_1003),
.Y(n_1325)
);

OAI21x1_ASAP7_75t_L g1326 ( 
.A1(n_1209),
.A2(n_1188),
.B(n_1199),
.Y(n_1326)
);

AOI221x1_ASAP7_75t_L g1327 ( 
.A1(n_1146),
.A2(n_1050),
.B1(n_1144),
.B2(n_1154),
.C(n_1232),
.Y(n_1327)
);

AOI22xp5_ASAP7_75t_L g1328 ( 
.A1(n_1096),
.A2(n_611),
.B1(n_770),
.B2(n_1003),
.Y(n_1328)
);

NAND2xp5_ASAP7_75t_L g1329 ( 
.A(n_1230),
.B(n_903),
.Y(n_1329)
);

AOI21xp5_ASAP7_75t_SL g1330 ( 
.A1(n_1181),
.A2(n_1050),
.B(n_958),
.Y(n_1330)
);

OAI21x1_ASAP7_75t_L g1331 ( 
.A1(n_1209),
.A2(n_1188),
.B(n_1199),
.Y(n_1331)
);

AOI21xp5_ASAP7_75t_L g1332 ( 
.A1(n_1187),
.A2(n_1041),
.B(n_952),
.Y(n_1332)
);

O2A1O1Ixp33_ASAP7_75t_SL g1333 ( 
.A1(n_1230),
.A2(n_1229),
.B(n_1050),
.C(n_903),
.Y(n_1333)
);

AO32x2_ASAP7_75t_L g1334 ( 
.A1(n_1179),
.A2(n_1115),
.A3(n_1144),
.B1(n_1191),
.B2(n_1043),
.Y(n_1334)
);

NAND2xp5_ASAP7_75t_L g1335 ( 
.A(n_1230),
.B(n_903),
.Y(n_1335)
);

A2O1A1Ixp33_ASAP7_75t_L g1336 ( 
.A1(n_1185),
.A2(n_1050),
.B(n_1003),
.C(n_1096),
.Y(n_1336)
);

NOR2xp33_ASAP7_75t_L g1337 ( 
.A(n_1230),
.B(n_611),
.Y(n_1337)
);

NAND2xp5_ASAP7_75t_L g1338 ( 
.A(n_1230),
.B(n_903),
.Y(n_1338)
);

AOI21xp5_ASAP7_75t_L g1339 ( 
.A1(n_1187),
.A2(n_1041),
.B(n_952),
.Y(n_1339)
);

AOI21xp5_ASAP7_75t_L g1340 ( 
.A1(n_1187),
.A2(n_1041),
.B(n_952),
.Y(n_1340)
);

NAND2xp5_ASAP7_75t_L g1341 ( 
.A(n_1230),
.B(n_1181),
.Y(n_1341)
);

NAND2xp5_ASAP7_75t_L g1342 ( 
.A(n_1230),
.B(n_1181),
.Y(n_1342)
);

NAND2xp5_ASAP7_75t_L g1343 ( 
.A(n_1230),
.B(n_1181),
.Y(n_1343)
);

AOI22xp33_ASAP7_75t_L g1344 ( 
.A1(n_1232),
.A2(n_602),
.B1(n_1003),
.B2(n_428),
.Y(n_1344)
);

AO31x2_ASAP7_75t_L g1345 ( 
.A1(n_1222),
.A2(n_1008),
.A3(n_923),
.B(n_1200),
.Y(n_1345)
);

OAI22xp5_ASAP7_75t_L g1346 ( 
.A1(n_1230),
.A2(n_1022),
.B1(n_1096),
.B2(n_1050),
.Y(n_1346)
);

NAND2xp5_ASAP7_75t_L g1347 ( 
.A(n_1230),
.B(n_1181),
.Y(n_1347)
);

OAI21xp5_ASAP7_75t_L g1348 ( 
.A1(n_1230),
.A2(n_1050),
.B(n_1154),
.Y(n_1348)
);

AO31x2_ASAP7_75t_L g1349 ( 
.A1(n_1222),
.A2(n_1008),
.A3(n_923),
.B(n_1200),
.Y(n_1349)
);

OAI21xp5_ASAP7_75t_L g1350 ( 
.A1(n_1230),
.A2(n_1050),
.B(n_1154),
.Y(n_1350)
);

NAND2xp5_ASAP7_75t_SL g1351 ( 
.A(n_1101),
.B(n_1022),
.Y(n_1351)
);

AOI31xp67_ASAP7_75t_L g1352 ( 
.A1(n_1224),
.A2(n_1100),
.A3(n_1157),
.B(n_1155),
.Y(n_1352)
);

O2A1O1Ixp33_ASAP7_75t_SL g1353 ( 
.A1(n_1230),
.A2(n_1229),
.B(n_1050),
.C(n_903),
.Y(n_1353)
);

AND2x4_ASAP7_75t_L g1354 ( 
.A(n_1228),
.B(n_909),
.Y(n_1354)
);

OAI21xp5_ASAP7_75t_L g1355 ( 
.A1(n_1230),
.A2(n_1050),
.B(n_1154),
.Y(n_1355)
);

NAND3xp33_ASAP7_75t_L g1356 ( 
.A(n_1096),
.B(n_1050),
.C(n_1141),
.Y(n_1356)
);

AOI221xp5_ASAP7_75t_SL g1357 ( 
.A1(n_1115),
.A2(n_1003),
.B1(n_1144),
.B2(n_1146),
.C(n_1096),
.Y(n_1357)
);

AO21x1_ASAP7_75t_L g1358 ( 
.A1(n_1185),
.A2(n_915),
.B(n_910),
.Y(n_1358)
);

AO31x2_ASAP7_75t_L g1359 ( 
.A1(n_1222),
.A2(n_1008),
.A3(n_923),
.B(n_1200),
.Y(n_1359)
);

A2O1A1Ixp33_ASAP7_75t_L g1360 ( 
.A1(n_1185),
.A2(n_1050),
.B(n_1003),
.C(n_1096),
.Y(n_1360)
);

AOI21xp5_ASAP7_75t_L g1361 ( 
.A1(n_1187),
.A2(n_1041),
.B(n_952),
.Y(n_1361)
);

AOI21xp5_ASAP7_75t_L g1362 ( 
.A1(n_1187),
.A2(n_1041),
.B(n_952),
.Y(n_1362)
);

AO31x2_ASAP7_75t_L g1363 ( 
.A1(n_1222),
.A2(n_1008),
.A3(n_923),
.B(n_1200),
.Y(n_1363)
);

NAND2xp5_ASAP7_75t_L g1364 ( 
.A(n_1230),
.B(n_1181),
.Y(n_1364)
);

NAND2xp5_ASAP7_75t_L g1365 ( 
.A(n_1230),
.B(n_1181),
.Y(n_1365)
);

AOI21xp5_ASAP7_75t_L g1366 ( 
.A1(n_1187),
.A2(n_1041),
.B(n_952),
.Y(n_1366)
);

OAI21x1_ASAP7_75t_L g1367 ( 
.A1(n_1209),
.A2(n_1188),
.B(n_1199),
.Y(n_1367)
);

INVx1_ASAP7_75t_L g1368 ( 
.A(n_1089),
.Y(n_1368)
);

AO31x2_ASAP7_75t_L g1369 ( 
.A1(n_1222),
.A2(n_1008),
.A3(n_923),
.B(n_1200),
.Y(n_1369)
);

INVx4_ASAP7_75t_L g1370 ( 
.A(n_1228),
.Y(n_1370)
);

INVx1_ASAP7_75t_L g1371 ( 
.A(n_1089),
.Y(n_1371)
);

CKINVDCx20_ASAP7_75t_R g1372 ( 
.A(n_1098),
.Y(n_1372)
);

NOR2xp33_ASAP7_75t_L g1373 ( 
.A(n_1230),
.B(n_611),
.Y(n_1373)
);

INVx3_ASAP7_75t_L g1374 ( 
.A(n_1202),
.Y(n_1374)
);

AOI22xp33_ASAP7_75t_L g1375 ( 
.A1(n_1232),
.A2(n_602),
.B1(n_1003),
.B2(n_428),
.Y(n_1375)
);

NAND3xp33_ASAP7_75t_SL g1376 ( 
.A(n_1088),
.B(n_555),
.C(n_540),
.Y(n_1376)
);

AO31x2_ASAP7_75t_L g1377 ( 
.A1(n_1222),
.A2(n_1008),
.A3(n_923),
.B(n_1200),
.Y(n_1377)
);

OAI21x1_ASAP7_75t_L g1378 ( 
.A1(n_1209),
.A2(n_1188),
.B(n_1199),
.Y(n_1378)
);

AOI22xp33_ASAP7_75t_L g1379 ( 
.A1(n_1253),
.A2(n_1356),
.B1(n_1242),
.B2(n_1344),
.Y(n_1379)
);

AOI22xp5_ASAP7_75t_L g1380 ( 
.A1(n_1337),
.A2(n_1373),
.B1(n_1264),
.B2(n_1356),
.Y(n_1380)
);

AOI22xp33_ASAP7_75t_L g1381 ( 
.A1(n_1375),
.A2(n_1273),
.B1(n_1260),
.B2(n_1245),
.Y(n_1381)
);

BUFx6f_ASAP7_75t_L g1382 ( 
.A(n_1354),
.Y(n_1382)
);

BUFx8_ASAP7_75t_SL g1383 ( 
.A(n_1372),
.Y(n_1383)
);

INVx1_ASAP7_75t_SL g1384 ( 
.A(n_1252),
.Y(n_1384)
);

OAI22xp5_ASAP7_75t_L g1385 ( 
.A1(n_1325),
.A2(n_1328),
.B1(n_1336),
.B2(n_1360),
.Y(n_1385)
);

INVx4_ASAP7_75t_L g1386 ( 
.A(n_1268),
.Y(n_1386)
);

INVx4_ASAP7_75t_L g1387 ( 
.A(n_1258),
.Y(n_1387)
);

OAI22xp33_ASAP7_75t_L g1388 ( 
.A1(n_1234),
.A2(n_1327),
.B1(n_1245),
.B2(n_1346),
.Y(n_1388)
);

BUFx2_ASAP7_75t_R g1389 ( 
.A(n_1236),
.Y(n_1389)
);

NAND2xp5_ASAP7_75t_SL g1390 ( 
.A(n_1251),
.B(n_1309),
.Y(n_1390)
);

AOI22xp33_ASAP7_75t_L g1391 ( 
.A1(n_1351),
.A2(n_1346),
.B1(n_1309),
.B2(n_1350),
.Y(n_1391)
);

INVx1_ASAP7_75t_L g1392 ( 
.A(n_1233),
.Y(n_1392)
);

BUFx3_ASAP7_75t_L g1393 ( 
.A(n_1266),
.Y(n_1393)
);

BUFx12f_ASAP7_75t_L g1394 ( 
.A(n_1310),
.Y(n_1394)
);

CKINVDCx20_ASAP7_75t_R g1395 ( 
.A(n_1310),
.Y(n_1395)
);

OAI22xp33_ASAP7_75t_L g1396 ( 
.A1(n_1312),
.A2(n_1323),
.B1(n_1348),
.B2(n_1355),
.Y(n_1396)
);

AOI22xp33_ASAP7_75t_L g1397 ( 
.A1(n_1323),
.A2(n_1237),
.B1(n_1286),
.B2(n_1251),
.Y(n_1397)
);

AOI22xp33_ASAP7_75t_L g1398 ( 
.A1(n_1376),
.A2(n_1358),
.B1(n_1248),
.B2(n_1250),
.Y(n_1398)
);

AOI22xp33_ASAP7_75t_L g1399 ( 
.A1(n_1250),
.A2(n_1347),
.B1(n_1341),
.B2(n_1365),
.Y(n_1399)
);

OAI21xp33_ASAP7_75t_L g1400 ( 
.A1(n_1317),
.A2(n_1243),
.B(n_1330),
.Y(n_1400)
);

BUFx2_ASAP7_75t_SL g1401 ( 
.A(n_1247),
.Y(n_1401)
);

NAND2xp5_ASAP7_75t_L g1402 ( 
.A(n_1315),
.B(n_1319),
.Y(n_1402)
);

AOI22xp5_ASAP7_75t_L g1403 ( 
.A1(n_1306),
.A2(n_1267),
.B1(n_1357),
.B2(n_1291),
.Y(n_1403)
);

OAI22xp5_ASAP7_75t_L g1404 ( 
.A1(n_1329),
.A2(n_1338),
.B1(n_1335),
.B2(n_1320),
.Y(n_1404)
);

INVx6_ASAP7_75t_L g1405 ( 
.A(n_1277),
.Y(n_1405)
);

AOI22xp33_ASAP7_75t_L g1406 ( 
.A1(n_1341),
.A2(n_1347),
.B1(n_1342),
.B2(n_1365),
.Y(n_1406)
);

OAI22x1_ASAP7_75t_SL g1407 ( 
.A1(n_1252),
.A2(n_1320),
.B1(n_1311),
.B2(n_1371),
.Y(n_1407)
);

AOI22xp33_ASAP7_75t_L g1408 ( 
.A1(n_1342),
.A2(n_1343),
.B1(n_1364),
.B2(n_1272),
.Y(n_1408)
);

OAI22xp33_ASAP7_75t_L g1409 ( 
.A1(n_1343),
.A2(n_1364),
.B1(n_1274),
.B2(n_1278),
.Y(n_1409)
);

BUFx2_ASAP7_75t_SL g1410 ( 
.A(n_1240),
.Y(n_1410)
);

BUFx12f_ASAP7_75t_L g1411 ( 
.A(n_1277),
.Y(n_1411)
);

CKINVDCx11_ASAP7_75t_R g1412 ( 
.A(n_1313),
.Y(n_1412)
);

BUFx2_ASAP7_75t_L g1413 ( 
.A(n_1324),
.Y(n_1413)
);

INVx1_ASAP7_75t_SL g1414 ( 
.A(n_1289),
.Y(n_1414)
);

AOI22xp33_ASAP7_75t_L g1415 ( 
.A1(n_1262),
.A2(n_1297),
.B1(n_1276),
.B2(n_1295),
.Y(n_1415)
);

BUFx2_ASAP7_75t_SL g1416 ( 
.A(n_1259),
.Y(n_1416)
);

INVx2_ASAP7_75t_L g1417 ( 
.A(n_1307),
.Y(n_1417)
);

OAI22xp33_ASAP7_75t_L g1418 ( 
.A1(n_1274),
.A2(n_1278),
.B1(n_1257),
.B2(n_1276),
.Y(n_1418)
);

CKINVDCx20_ASAP7_75t_R g1419 ( 
.A(n_1296),
.Y(n_1419)
);

AOI22xp5_ASAP7_75t_L g1420 ( 
.A1(n_1357),
.A2(n_1259),
.B1(n_1281),
.B2(n_1279),
.Y(n_1420)
);

BUFx3_ASAP7_75t_L g1421 ( 
.A(n_1285),
.Y(n_1421)
);

INVx2_ASAP7_75t_L g1422 ( 
.A(n_1368),
.Y(n_1422)
);

BUFx2_ASAP7_75t_R g1423 ( 
.A(n_1304),
.Y(n_1423)
);

BUFx10_ASAP7_75t_L g1424 ( 
.A(n_1285),
.Y(n_1424)
);

AND2x2_ASAP7_75t_L g1425 ( 
.A(n_1255),
.B(n_1370),
.Y(n_1425)
);

INVx6_ASAP7_75t_L g1426 ( 
.A(n_1370),
.Y(n_1426)
);

INVx1_ASAP7_75t_L g1427 ( 
.A(n_1284),
.Y(n_1427)
);

INVx1_ASAP7_75t_L g1428 ( 
.A(n_1288),
.Y(n_1428)
);

INVx1_ASAP7_75t_L g1429 ( 
.A(n_1288),
.Y(n_1429)
);

INVx1_ASAP7_75t_L g1430 ( 
.A(n_1300),
.Y(n_1430)
);

AOI22xp33_ASAP7_75t_L g1431 ( 
.A1(n_1280),
.A2(n_1281),
.B1(n_1283),
.B2(n_1270),
.Y(n_1431)
);

CKINVDCx5p33_ASAP7_75t_R g1432 ( 
.A(n_1255),
.Y(n_1432)
);

CKINVDCx20_ASAP7_75t_R g1433 ( 
.A(n_1290),
.Y(n_1433)
);

BUFx10_ASAP7_75t_L g1434 ( 
.A(n_1292),
.Y(n_1434)
);

AOI22xp5_ASAP7_75t_L g1435 ( 
.A1(n_1244),
.A2(n_1294),
.B1(n_1333),
.B2(n_1353),
.Y(n_1435)
);

NAND2x1p5_ASAP7_75t_L g1436 ( 
.A(n_1374),
.B(n_1298),
.Y(n_1436)
);

BUFx2_ASAP7_75t_SL g1437 ( 
.A(n_1305),
.Y(n_1437)
);

AOI22xp5_ASAP7_75t_L g1438 ( 
.A1(n_1280),
.A2(n_1374),
.B1(n_1283),
.B2(n_1299),
.Y(n_1438)
);

INVx1_ASAP7_75t_L g1439 ( 
.A(n_1282),
.Y(n_1439)
);

HB1xp67_ASAP7_75t_L g1440 ( 
.A(n_1345),
.Y(n_1440)
);

INVx6_ASAP7_75t_L g1441 ( 
.A(n_1301),
.Y(n_1441)
);

INVx1_ASAP7_75t_L g1442 ( 
.A(n_1269),
.Y(n_1442)
);

CKINVDCx11_ASAP7_75t_R g1443 ( 
.A(n_1303),
.Y(n_1443)
);

BUFx2_ASAP7_75t_L g1444 ( 
.A(n_1302),
.Y(n_1444)
);

CKINVDCx11_ASAP7_75t_R g1445 ( 
.A(n_1261),
.Y(n_1445)
);

INVx1_ASAP7_75t_L g1446 ( 
.A(n_1269),
.Y(n_1446)
);

INVx6_ASAP7_75t_L g1447 ( 
.A(n_1275),
.Y(n_1447)
);

NAND2xp5_ASAP7_75t_L g1448 ( 
.A(n_1314),
.B(n_1321),
.Y(n_1448)
);

BUFx2_ASAP7_75t_SL g1449 ( 
.A(n_1249),
.Y(n_1449)
);

CKINVDCx11_ASAP7_75t_R g1450 ( 
.A(n_1334),
.Y(n_1450)
);

CKINVDCx6p67_ASAP7_75t_R g1451 ( 
.A(n_1334),
.Y(n_1451)
);

INVxp67_ASAP7_75t_L g1452 ( 
.A(n_1256),
.Y(n_1452)
);

NAND2x1p5_ASAP7_75t_L g1453 ( 
.A(n_1271),
.B(n_1265),
.Y(n_1453)
);

NAND2x1p5_ASAP7_75t_L g1454 ( 
.A(n_1241),
.B(n_1366),
.Y(n_1454)
);

INVx6_ASAP7_75t_L g1455 ( 
.A(n_1334),
.Y(n_1455)
);

INVx6_ASAP7_75t_L g1456 ( 
.A(n_1246),
.Y(n_1456)
);

AOI22xp33_ASAP7_75t_L g1457 ( 
.A1(n_1322),
.A2(n_1362),
.B1(n_1339),
.B2(n_1340),
.Y(n_1457)
);

INVx1_ASAP7_75t_L g1458 ( 
.A(n_1263),
.Y(n_1458)
);

OAI21xp5_ASAP7_75t_SL g1459 ( 
.A1(n_1293),
.A2(n_1361),
.B(n_1332),
.Y(n_1459)
);

AOI22xp33_ASAP7_75t_SL g1460 ( 
.A1(n_1308),
.A2(n_1238),
.B1(n_1287),
.B2(n_1235),
.Y(n_1460)
);

BUFx2_ASAP7_75t_SL g1461 ( 
.A(n_1308),
.Y(n_1461)
);

CKINVDCx20_ASAP7_75t_R g1462 ( 
.A(n_1239),
.Y(n_1462)
);

INVx1_ASAP7_75t_L g1463 ( 
.A(n_1263),
.Y(n_1463)
);

INVx6_ASAP7_75t_L g1464 ( 
.A(n_1352),
.Y(n_1464)
);

BUFx6f_ASAP7_75t_L g1465 ( 
.A(n_1254),
.Y(n_1465)
);

BUFx2_ASAP7_75t_SL g1466 ( 
.A(n_1345),
.Y(n_1466)
);

CKINVDCx20_ASAP7_75t_R g1467 ( 
.A(n_1349),
.Y(n_1467)
);

NAND2xp5_ASAP7_75t_L g1468 ( 
.A(n_1349),
.B(n_1363),
.Y(n_1468)
);

OAI21xp5_ASAP7_75t_SL g1469 ( 
.A1(n_1316),
.A2(n_1326),
.B(n_1331),
.Y(n_1469)
);

INVx1_ASAP7_75t_L g1470 ( 
.A(n_1349),
.Y(n_1470)
);

AOI22xp33_ASAP7_75t_L g1471 ( 
.A1(n_1367),
.A2(n_1378),
.B1(n_1363),
.B2(n_1369),
.Y(n_1471)
);

INVx1_ASAP7_75t_L g1472 ( 
.A(n_1359),
.Y(n_1472)
);

AND2x2_ASAP7_75t_L g1473 ( 
.A(n_1359),
.B(n_1363),
.Y(n_1473)
);

CKINVDCx20_ASAP7_75t_R g1474 ( 
.A(n_1369),
.Y(n_1474)
);

AOI22xp33_ASAP7_75t_L g1475 ( 
.A1(n_1377),
.A2(n_1253),
.B1(n_1356),
.B2(n_1232),
.Y(n_1475)
);

AOI22xp33_ASAP7_75t_L g1476 ( 
.A1(n_1377),
.A2(n_1253),
.B1(n_1356),
.B2(n_1232),
.Y(n_1476)
);

OAI22xp33_ASAP7_75t_L g1477 ( 
.A1(n_1356),
.A2(n_1325),
.B1(n_1328),
.B2(n_1088),
.Y(n_1477)
);

AOI22xp33_ASAP7_75t_L g1478 ( 
.A1(n_1253),
.A2(n_1356),
.B1(n_1232),
.B2(n_1242),
.Y(n_1478)
);

AOI22xp33_ASAP7_75t_L g1479 ( 
.A1(n_1253),
.A2(n_1356),
.B1(n_1232),
.B2(n_1242),
.Y(n_1479)
);

AOI22xp33_ASAP7_75t_SL g1480 ( 
.A1(n_1253),
.A2(n_1356),
.B1(n_1245),
.B2(n_1346),
.Y(n_1480)
);

BUFx12f_ASAP7_75t_L g1481 ( 
.A(n_1310),
.Y(n_1481)
);

INVx3_ASAP7_75t_L g1482 ( 
.A(n_1354),
.Y(n_1482)
);

OAI22xp5_ASAP7_75t_L g1483 ( 
.A1(n_1325),
.A2(n_1328),
.B1(n_1356),
.B2(n_1022),
.Y(n_1483)
);

BUFx12f_ASAP7_75t_L g1484 ( 
.A(n_1310),
.Y(n_1484)
);

AOI22xp5_ASAP7_75t_L g1485 ( 
.A1(n_1337),
.A2(n_1373),
.B1(n_1253),
.B2(n_1264),
.Y(n_1485)
);

AOI22xp5_ASAP7_75t_L g1486 ( 
.A1(n_1337),
.A2(n_1373),
.B1(n_1253),
.B2(n_1264),
.Y(n_1486)
);

OAI22xp5_ASAP7_75t_L g1487 ( 
.A1(n_1325),
.A2(n_1328),
.B1(n_1356),
.B2(n_1022),
.Y(n_1487)
);

BUFx10_ASAP7_75t_L g1488 ( 
.A(n_1267),
.Y(n_1488)
);

AOI22xp33_ASAP7_75t_L g1489 ( 
.A1(n_1253),
.A2(n_1356),
.B1(n_1232),
.B2(n_1242),
.Y(n_1489)
);

AOI22xp33_ASAP7_75t_L g1490 ( 
.A1(n_1253),
.A2(n_1356),
.B1(n_1232),
.B2(n_1242),
.Y(n_1490)
);

NAND2xp5_ASAP7_75t_L g1491 ( 
.A(n_1234),
.B(n_1315),
.Y(n_1491)
);

AOI22xp33_ASAP7_75t_L g1492 ( 
.A1(n_1253),
.A2(n_1356),
.B1(n_1232),
.B2(n_1242),
.Y(n_1492)
);

OAI22xp5_ASAP7_75t_L g1493 ( 
.A1(n_1325),
.A2(n_1328),
.B1(n_1356),
.B2(n_1022),
.Y(n_1493)
);

OAI22xp5_ASAP7_75t_L g1494 ( 
.A1(n_1325),
.A2(n_1328),
.B1(n_1356),
.B2(n_1022),
.Y(n_1494)
);

AOI22xp33_ASAP7_75t_SL g1495 ( 
.A1(n_1253),
.A2(n_1356),
.B1(n_1245),
.B2(n_1346),
.Y(n_1495)
);

OAI22xp5_ASAP7_75t_L g1496 ( 
.A1(n_1325),
.A2(n_1328),
.B1(n_1356),
.B2(n_1022),
.Y(n_1496)
);

AOI22xp33_ASAP7_75t_SL g1497 ( 
.A1(n_1253),
.A2(n_1356),
.B1(n_1245),
.B2(n_1346),
.Y(n_1497)
);

AND2x2_ASAP7_75t_L g1498 ( 
.A(n_1286),
.B(n_1318),
.Y(n_1498)
);

INVx1_ASAP7_75t_SL g1499 ( 
.A(n_1252),
.Y(n_1499)
);

AOI22xp33_ASAP7_75t_SL g1500 ( 
.A1(n_1253),
.A2(n_1356),
.B1(n_1245),
.B2(n_1346),
.Y(n_1500)
);

BUFx8_ASAP7_75t_L g1501 ( 
.A(n_1268),
.Y(n_1501)
);

BUFx3_ASAP7_75t_L g1502 ( 
.A(n_1268),
.Y(n_1502)
);

INVx1_ASAP7_75t_L g1503 ( 
.A(n_1458),
.Y(n_1503)
);

INVx3_ASAP7_75t_L g1504 ( 
.A(n_1447),
.Y(n_1504)
);

BUFx2_ASAP7_75t_SL g1505 ( 
.A(n_1434),
.Y(n_1505)
);

AND2x2_ASAP7_75t_L g1506 ( 
.A(n_1451),
.B(n_1455),
.Y(n_1506)
);

AND2x2_ASAP7_75t_L g1507 ( 
.A(n_1455),
.B(n_1450),
.Y(n_1507)
);

BUFx2_ASAP7_75t_L g1508 ( 
.A(n_1444),
.Y(n_1508)
);

OA21x2_ASAP7_75t_L g1509 ( 
.A1(n_1459),
.A2(n_1469),
.B(n_1471),
.Y(n_1509)
);

INVx1_ASAP7_75t_L g1510 ( 
.A(n_1463),
.Y(n_1510)
);

O2A1O1Ixp33_ASAP7_75t_L g1511 ( 
.A1(n_1477),
.A2(n_1496),
.B(n_1493),
.C(n_1494),
.Y(n_1511)
);

INVx1_ASAP7_75t_L g1512 ( 
.A(n_1442),
.Y(n_1512)
);

INVx1_ASAP7_75t_L g1513 ( 
.A(n_1446),
.Y(n_1513)
);

INVx1_ASAP7_75t_L g1514 ( 
.A(n_1428),
.Y(n_1514)
);

INVx1_ASAP7_75t_L g1515 ( 
.A(n_1429),
.Y(n_1515)
);

INVx1_ASAP7_75t_L g1516 ( 
.A(n_1470),
.Y(n_1516)
);

INVx1_ASAP7_75t_L g1517 ( 
.A(n_1472),
.Y(n_1517)
);

INVx3_ASAP7_75t_L g1518 ( 
.A(n_1447),
.Y(n_1518)
);

INVx2_ASAP7_75t_L g1519 ( 
.A(n_1473),
.Y(n_1519)
);

INVx1_ASAP7_75t_L g1520 ( 
.A(n_1440),
.Y(n_1520)
);

AO31x2_ASAP7_75t_L g1521 ( 
.A1(n_1468),
.A2(n_1385),
.A3(n_1448),
.B(n_1430),
.Y(n_1521)
);

BUFx2_ASAP7_75t_L g1522 ( 
.A(n_1452),
.Y(n_1522)
);

INVxp67_ASAP7_75t_L g1523 ( 
.A(n_1413),
.Y(n_1523)
);

AOI21xp5_ASAP7_75t_L g1524 ( 
.A1(n_1396),
.A2(n_1400),
.B(n_1388),
.Y(n_1524)
);

INVx2_ASAP7_75t_SL g1525 ( 
.A(n_1441),
.Y(n_1525)
);

INVx1_ASAP7_75t_L g1526 ( 
.A(n_1392),
.Y(n_1526)
);

OAI21x1_ASAP7_75t_L g1527 ( 
.A1(n_1453),
.A2(n_1471),
.B(n_1454),
.Y(n_1527)
);

INVx1_ASAP7_75t_L g1528 ( 
.A(n_1417),
.Y(n_1528)
);

AOI21xp5_ASAP7_75t_L g1529 ( 
.A1(n_1396),
.A2(n_1388),
.B(n_1390),
.Y(n_1529)
);

INVx1_ASAP7_75t_L g1530 ( 
.A(n_1422),
.Y(n_1530)
);

INVx2_ASAP7_75t_SL g1531 ( 
.A(n_1441),
.Y(n_1531)
);

NAND2x1p5_ASAP7_75t_L g1532 ( 
.A(n_1438),
.B(n_1420),
.Y(n_1532)
);

AND2x2_ASAP7_75t_L g1533 ( 
.A(n_1480),
.B(n_1495),
.Y(n_1533)
);

INVx1_ASAP7_75t_L g1534 ( 
.A(n_1452),
.Y(n_1534)
);

INVx2_ASAP7_75t_SL g1535 ( 
.A(n_1441),
.Y(n_1535)
);

BUFx2_ASAP7_75t_L g1536 ( 
.A(n_1454),
.Y(n_1536)
);

AND2x2_ASAP7_75t_L g1537 ( 
.A(n_1480),
.B(n_1495),
.Y(n_1537)
);

INVx3_ASAP7_75t_L g1538 ( 
.A(n_1447),
.Y(n_1538)
);

INVx2_ASAP7_75t_SL g1539 ( 
.A(n_1436),
.Y(n_1539)
);

OR2x2_ASAP7_75t_L g1540 ( 
.A(n_1397),
.B(n_1427),
.Y(n_1540)
);

INVx1_ASAP7_75t_L g1541 ( 
.A(n_1439),
.Y(n_1541)
);

AOI22xp33_ASAP7_75t_L g1542 ( 
.A1(n_1379),
.A2(n_1479),
.B1(n_1489),
.B2(n_1490),
.Y(n_1542)
);

HB1xp67_ASAP7_75t_L g1543 ( 
.A(n_1384),
.Y(n_1543)
);

INVx1_ASAP7_75t_L g1544 ( 
.A(n_1466),
.Y(n_1544)
);

BUFx2_ASAP7_75t_L g1545 ( 
.A(n_1462),
.Y(n_1545)
);

NAND2xp5_ASAP7_75t_L g1546 ( 
.A(n_1406),
.B(n_1399),
.Y(n_1546)
);

AO21x1_ASAP7_75t_L g1547 ( 
.A1(n_1477),
.A2(n_1418),
.B(n_1409),
.Y(n_1547)
);

OAI21x1_ASAP7_75t_L g1548 ( 
.A1(n_1453),
.A2(n_1457),
.B(n_1436),
.Y(n_1548)
);

AOI22xp33_ASAP7_75t_SL g1549 ( 
.A1(n_1467),
.A2(n_1474),
.B1(n_1487),
.B2(n_1483),
.Y(n_1549)
);

OAI21x1_ASAP7_75t_L g1550 ( 
.A1(n_1457),
.A2(n_1431),
.B(n_1435),
.Y(n_1550)
);

AOI22xp33_ASAP7_75t_L g1551 ( 
.A1(n_1379),
.A2(n_1479),
.B1(n_1490),
.B2(n_1492),
.Y(n_1551)
);

A2O1A1Ixp33_ASAP7_75t_SL g1552 ( 
.A1(n_1380),
.A2(n_1403),
.B(n_1398),
.C(n_1391),
.Y(n_1552)
);

AO21x2_ASAP7_75t_L g1553 ( 
.A1(n_1409),
.A2(n_1418),
.B(n_1404),
.Y(n_1553)
);

OAI21x1_ASAP7_75t_L g1554 ( 
.A1(n_1431),
.A2(n_1391),
.B(n_1398),
.Y(n_1554)
);

OR2x2_ASAP7_75t_L g1555 ( 
.A(n_1475),
.B(n_1476),
.Y(n_1555)
);

INVx2_ASAP7_75t_SL g1556 ( 
.A(n_1425),
.Y(n_1556)
);

BUFx6f_ASAP7_75t_L g1557 ( 
.A(n_1443),
.Y(n_1557)
);

OA21x2_ASAP7_75t_L g1558 ( 
.A1(n_1475),
.A2(n_1476),
.B(n_1415),
.Y(n_1558)
);

NAND2xp5_ASAP7_75t_L g1559 ( 
.A(n_1406),
.B(n_1399),
.Y(n_1559)
);

INVx1_ASAP7_75t_L g1560 ( 
.A(n_1461),
.Y(n_1560)
);

BUFx6f_ASAP7_75t_L g1561 ( 
.A(n_1445),
.Y(n_1561)
);

INVx1_ASAP7_75t_L g1562 ( 
.A(n_1456),
.Y(n_1562)
);

INVx1_ASAP7_75t_L g1563 ( 
.A(n_1456),
.Y(n_1563)
);

INVx3_ASAP7_75t_L g1564 ( 
.A(n_1464),
.Y(n_1564)
);

INVx1_ASAP7_75t_L g1565 ( 
.A(n_1464),
.Y(n_1565)
);

HB1xp67_ASAP7_75t_L g1566 ( 
.A(n_1499),
.Y(n_1566)
);

INVx2_ASAP7_75t_SL g1567 ( 
.A(n_1426),
.Y(n_1567)
);

AND2x2_ASAP7_75t_L g1568 ( 
.A(n_1497),
.B(n_1500),
.Y(n_1568)
);

INVx1_ASAP7_75t_L g1569 ( 
.A(n_1465),
.Y(n_1569)
);

AND2x2_ASAP7_75t_L g1570 ( 
.A(n_1497),
.B(n_1500),
.Y(n_1570)
);

OAI21x1_ASAP7_75t_L g1571 ( 
.A1(n_1415),
.A2(n_1492),
.B(n_1478),
.Y(n_1571)
);

INVx1_ASAP7_75t_L g1572 ( 
.A(n_1465),
.Y(n_1572)
);

INVx2_ASAP7_75t_L g1573 ( 
.A(n_1449),
.Y(n_1573)
);

INVx1_ASAP7_75t_L g1574 ( 
.A(n_1460),
.Y(n_1574)
);

INVx1_ASAP7_75t_L g1575 ( 
.A(n_1460),
.Y(n_1575)
);

OAI21x1_ASAP7_75t_L g1576 ( 
.A1(n_1478),
.A2(n_1489),
.B(n_1482),
.Y(n_1576)
);

HB1xp67_ASAP7_75t_L g1577 ( 
.A(n_1498),
.Y(n_1577)
);

INVx1_ASAP7_75t_L g1578 ( 
.A(n_1437),
.Y(n_1578)
);

INVx3_ASAP7_75t_L g1579 ( 
.A(n_1434),
.Y(n_1579)
);

AOI222xp33_ASAP7_75t_L g1580 ( 
.A1(n_1381),
.A2(n_1407),
.B1(n_1408),
.B2(n_1402),
.C1(n_1491),
.C2(n_1414),
.Y(n_1580)
);

INVxp67_ASAP7_75t_L g1581 ( 
.A(n_1393),
.Y(n_1581)
);

AOI21x1_ASAP7_75t_L g1582 ( 
.A1(n_1410),
.A2(n_1381),
.B(n_1426),
.Y(n_1582)
);

AND2x2_ASAP7_75t_L g1583 ( 
.A(n_1408),
.B(n_1485),
.Y(n_1583)
);

INVx1_ASAP7_75t_SL g1584 ( 
.A(n_1412),
.Y(n_1584)
);

CKINVDCx11_ASAP7_75t_R g1585 ( 
.A(n_1395),
.Y(n_1585)
);

BUFx3_ASAP7_75t_L g1586 ( 
.A(n_1433),
.Y(n_1586)
);

INVx1_ASAP7_75t_L g1587 ( 
.A(n_1382),
.Y(n_1587)
);

INVx1_ASAP7_75t_L g1588 ( 
.A(n_1382),
.Y(n_1588)
);

AOI22xp33_ASAP7_75t_L g1589 ( 
.A1(n_1486),
.A2(n_1488),
.B1(n_1421),
.B2(n_1416),
.Y(n_1589)
);

INVx2_ASAP7_75t_SL g1590 ( 
.A(n_1405),
.Y(n_1590)
);

INVx2_ASAP7_75t_SL g1591 ( 
.A(n_1405),
.Y(n_1591)
);

CKINVDCx20_ASAP7_75t_R g1592 ( 
.A(n_1383),
.Y(n_1592)
);

BUFx3_ASAP7_75t_L g1593 ( 
.A(n_1419),
.Y(n_1593)
);

INVx1_ASAP7_75t_L g1594 ( 
.A(n_1424),
.Y(n_1594)
);

INVx1_ASAP7_75t_L g1595 ( 
.A(n_1432),
.Y(n_1595)
);

OA21x2_ASAP7_75t_L g1596 ( 
.A1(n_1423),
.A2(n_1488),
.B(n_1411),
.Y(n_1596)
);

OA21x2_ASAP7_75t_L g1597 ( 
.A1(n_1524),
.A2(n_1401),
.B(n_1389),
.Y(n_1597)
);

INVx1_ASAP7_75t_SL g1598 ( 
.A(n_1545),
.Y(n_1598)
);

OAI21xp5_ASAP7_75t_L g1599 ( 
.A1(n_1511),
.A2(n_1387),
.B(n_1386),
.Y(n_1599)
);

OAI211xp5_ASAP7_75t_SL g1600 ( 
.A1(n_1523),
.A2(n_1394),
.B(n_1481),
.C(n_1484),
.Y(n_1600)
);

OAI22xp5_ASAP7_75t_L g1601 ( 
.A1(n_1533),
.A2(n_1501),
.B1(n_1502),
.B2(n_1537),
.Y(n_1601)
);

NAND2xp5_ASAP7_75t_L g1602 ( 
.A(n_1543),
.B(n_1501),
.Y(n_1602)
);

AND2x2_ASAP7_75t_L g1603 ( 
.A(n_1545),
.B(n_1577),
.Y(n_1603)
);

NOR2xp33_ASAP7_75t_L g1604 ( 
.A(n_1586),
.B(n_1581),
.Y(n_1604)
);

OAI22xp5_ASAP7_75t_L g1605 ( 
.A1(n_1568),
.A2(n_1570),
.B1(n_1551),
.B2(n_1542),
.Y(n_1605)
);

OR2x6_ASAP7_75t_L g1606 ( 
.A(n_1532),
.B(n_1547),
.Y(n_1606)
);

AO32x2_ASAP7_75t_L g1607 ( 
.A1(n_1556),
.A2(n_1525),
.A3(n_1531),
.B1(n_1535),
.B2(n_1539),
.Y(n_1607)
);

INVx1_ASAP7_75t_L g1608 ( 
.A(n_1526),
.Y(n_1608)
);

A2O1A1Ixp33_ASAP7_75t_L g1609 ( 
.A1(n_1529),
.A2(n_1552),
.B(n_1549),
.C(n_1571),
.Y(n_1609)
);

HB1xp67_ASAP7_75t_L g1610 ( 
.A(n_1566),
.Y(n_1610)
);

AO32x2_ASAP7_75t_L g1611 ( 
.A1(n_1525),
.A2(n_1531),
.A3(n_1535),
.B1(n_1539),
.B2(n_1590),
.Y(n_1611)
);

OAI21x1_ASAP7_75t_L g1612 ( 
.A1(n_1548),
.A2(n_1582),
.B(n_1527),
.Y(n_1612)
);

NAND2xp5_ASAP7_75t_L g1613 ( 
.A(n_1521),
.B(n_1522),
.Y(n_1613)
);

AOI21xp5_ASAP7_75t_SL g1614 ( 
.A1(n_1553),
.A2(n_1596),
.B(n_1561),
.Y(n_1614)
);

AOI22xp5_ASAP7_75t_L g1615 ( 
.A1(n_1547),
.A2(n_1553),
.B1(n_1583),
.B2(n_1580),
.Y(n_1615)
);

AND2x2_ASAP7_75t_L g1616 ( 
.A(n_1506),
.B(n_1507),
.Y(n_1616)
);

NOR2xp33_ASAP7_75t_R g1617 ( 
.A(n_1592),
.B(n_1585),
.Y(n_1617)
);

CKINVDCx5p33_ASAP7_75t_R g1618 ( 
.A(n_1593),
.Y(n_1618)
);

A2O1A1Ixp33_ASAP7_75t_L g1619 ( 
.A1(n_1571),
.A2(n_1554),
.B(n_1583),
.C(n_1546),
.Y(n_1619)
);

AND2x2_ASAP7_75t_L g1620 ( 
.A(n_1586),
.B(n_1595),
.Y(n_1620)
);

OAI22xp5_ASAP7_75t_L g1621 ( 
.A1(n_1559),
.A2(n_1555),
.B1(n_1575),
.B2(n_1574),
.Y(n_1621)
);

OR2x6_ASAP7_75t_L g1622 ( 
.A(n_1532),
.B(n_1582),
.Y(n_1622)
);

NAND2xp5_ASAP7_75t_L g1623 ( 
.A(n_1521),
.B(n_1534),
.Y(n_1623)
);

OAI22xp5_ASAP7_75t_L g1624 ( 
.A1(n_1574),
.A2(n_1575),
.B1(n_1505),
.B2(n_1540),
.Y(n_1624)
);

NAND2xp33_ASAP7_75t_L g1625 ( 
.A(n_1579),
.B(n_1557),
.Y(n_1625)
);

AND2x2_ASAP7_75t_L g1626 ( 
.A(n_1593),
.B(n_1508),
.Y(n_1626)
);

OAI21xp5_ASAP7_75t_L g1627 ( 
.A1(n_1554),
.A2(n_1550),
.B(n_1576),
.Y(n_1627)
);

BUFx6f_ASAP7_75t_L g1628 ( 
.A(n_1561),
.Y(n_1628)
);

OAI21xp5_ASAP7_75t_L g1629 ( 
.A1(n_1550),
.A2(n_1576),
.B(n_1534),
.Y(n_1629)
);

NAND2xp5_ASAP7_75t_L g1630 ( 
.A(n_1521),
.B(n_1540),
.Y(n_1630)
);

OAI21xp5_ASAP7_75t_L g1631 ( 
.A1(n_1578),
.A2(n_1579),
.B(n_1558),
.Y(n_1631)
);

OAI22xp5_ASAP7_75t_L g1632 ( 
.A1(n_1589),
.A2(n_1558),
.B1(n_1557),
.B2(n_1596),
.Y(n_1632)
);

OA21x2_ASAP7_75t_L g1633 ( 
.A1(n_1527),
.A2(n_1560),
.B(n_1544),
.Y(n_1633)
);

AO32x2_ASAP7_75t_L g1634 ( 
.A1(n_1590),
.A2(n_1591),
.A3(n_1567),
.B1(n_1519),
.B2(n_1558),
.Y(n_1634)
);

OAI22xp5_ASAP7_75t_L g1635 ( 
.A1(n_1557),
.A2(n_1596),
.B1(n_1509),
.B2(n_1584),
.Y(n_1635)
);

OAI22xp5_ASAP7_75t_SL g1636 ( 
.A1(n_1557),
.A2(n_1596),
.B1(n_1509),
.B2(n_1591),
.Y(n_1636)
);

CKINVDCx5p33_ASAP7_75t_R g1637 ( 
.A(n_1557),
.Y(n_1637)
);

OAI21xp5_ASAP7_75t_L g1638 ( 
.A1(n_1578),
.A2(n_1573),
.B(n_1509),
.Y(n_1638)
);

AND2x2_ASAP7_75t_L g1639 ( 
.A(n_1587),
.B(n_1588),
.Y(n_1639)
);

NAND4xp25_ASAP7_75t_L g1640 ( 
.A(n_1541),
.B(n_1536),
.C(n_1565),
.D(n_1563),
.Y(n_1640)
);

OAI21xp5_ASAP7_75t_L g1641 ( 
.A1(n_1573),
.A2(n_1509),
.B(n_1504),
.Y(n_1641)
);

AND2x2_ASAP7_75t_L g1642 ( 
.A(n_1587),
.B(n_1588),
.Y(n_1642)
);

OA21x2_ASAP7_75t_L g1643 ( 
.A1(n_1560),
.A2(n_1544),
.B(n_1562),
.Y(n_1643)
);

INVxp67_ASAP7_75t_L g1644 ( 
.A(n_1594),
.Y(n_1644)
);

NAND2xp5_ASAP7_75t_L g1645 ( 
.A(n_1528),
.B(n_1530),
.Y(n_1645)
);

OR2x2_ASAP7_75t_L g1646 ( 
.A(n_1630),
.B(n_1520),
.Y(n_1646)
);

INVx1_ASAP7_75t_L g1647 ( 
.A(n_1608),
.Y(n_1647)
);

AND2x2_ASAP7_75t_L g1648 ( 
.A(n_1641),
.B(n_1638),
.Y(n_1648)
);

BUFx2_ASAP7_75t_L g1649 ( 
.A(n_1611),
.Y(n_1649)
);

AND2x2_ASAP7_75t_L g1650 ( 
.A(n_1638),
.B(n_1569),
.Y(n_1650)
);

NAND2xp5_ASAP7_75t_L g1651 ( 
.A(n_1623),
.B(n_1613),
.Y(n_1651)
);

INVxp67_ASAP7_75t_L g1652 ( 
.A(n_1643),
.Y(n_1652)
);

INVx3_ASAP7_75t_L g1653 ( 
.A(n_1633),
.Y(n_1653)
);

INVxp67_ASAP7_75t_L g1654 ( 
.A(n_1613),
.Y(n_1654)
);

INVxp67_ASAP7_75t_SL g1655 ( 
.A(n_1623),
.Y(n_1655)
);

NOR2x1_ASAP7_75t_L g1656 ( 
.A(n_1635),
.B(n_1538),
.Y(n_1656)
);

AND2x4_ASAP7_75t_L g1657 ( 
.A(n_1631),
.B(n_1564),
.Y(n_1657)
);

HB1xp67_ASAP7_75t_L g1658 ( 
.A(n_1610),
.Y(n_1658)
);

INVx2_ASAP7_75t_L g1659 ( 
.A(n_1633),
.Y(n_1659)
);

INVx5_ASAP7_75t_L g1660 ( 
.A(n_1606),
.Y(n_1660)
);

OAI22xp5_ASAP7_75t_L g1661 ( 
.A1(n_1615),
.A2(n_1538),
.B1(n_1518),
.B2(n_1536),
.Y(n_1661)
);

AOI22xp33_ASAP7_75t_L g1662 ( 
.A1(n_1605),
.A2(n_1513),
.B1(n_1512),
.B2(n_1516),
.Y(n_1662)
);

AND2x2_ASAP7_75t_L g1663 ( 
.A(n_1634),
.B(n_1572),
.Y(n_1663)
);

INVx1_ASAP7_75t_L g1664 ( 
.A(n_1645),
.Y(n_1664)
);

AOI22xp33_ASAP7_75t_L g1665 ( 
.A1(n_1605),
.A2(n_1513),
.B1(n_1512),
.B2(n_1517),
.Y(n_1665)
);

AND2x2_ASAP7_75t_L g1666 ( 
.A(n_1634),
.B(n_1631),
.Y(n_1666)
);

NOR2xp67_ASAP7_75t_L g1667 ( 
.A(n_1635),
.B(n_1518),
.Y(n_1667)
);

BUFx2_ASAP7_75t_L g1668 ( 
.A(n_1611),
.Y(n_1668)
);

INVx2_ASAP7_75t_L g1669 ( 
.A(n_1634),
.Y(n_1669)
);

AOI221xp5_ASAP7_75t_L g1670 ( 
.A1(n_1621),
.A2(n_1503),
.B1(n_1510),
.B2(n_1515),
.C(n_1514),
.Y(n_1670)
);

INVx1_ASAP7_75t_L g1671 ( 
.A(n_1607),
.Y(n_1671)
);

INVx2_ASAP7_75t_L g1672 ( 
.A(n_1607),
.Y(n_1672)
);

INVx1_ASAP7_75t_L g1673 ( 
.A(n_1607),
.Y(n_1673)
);

AND2x2_ASAP7_75t_L g1674 ( 
.A(n_1616),
.B(n_1518),
.Y(n_1674)
);

INVx3_ASAP7_75t_SL g1675 ( 
.A(n_1637),
.Y(n_1675)
);

AND2x2_ASAP7_75t_L g1676 ( 
.A(n_1649),
.B(n_1626),
.Y(n_1676)
);

INVx2_ASAP7_75t_L g1677 ( 
.A(n_1659),
.Y(n_1677)
);

NAND2xp5_ASAP7_75t_L g1678 ( 
.A(n_1651),
.B(n_1619),
.Y(n_1678)
);

AND2x2_ASAP7_75t_L g1679 ( 
.A(n_1649),
.B(n_1603),
.Y(n_1679)
);

OAI31xp33_ASAP7_75t_L g1680 ( 
.A1(n_1661),
.A2(n_1609),
.A3(n_1601),
.B(n_1624),
.Y(n_1680)
);

AND2x2_ASAP7_75t_L g1681 ( 
.A(n_1668),
.B(n_1629),
.Y(n_1681)
);

OAI33xp33_ASAP7_75t_L g1682 ( 
.A1(n_1651),
.A2(n_1621),
.A3(n_1601),
.B1(n_1624),
.B2(n_1632),
.B3(n_1636),
.Y(n_1682)
);

AND2x2_ASAP7_75t_L g1683 ( 
.A(n_1668),
.B(n_1629),
.Y(n_1683)
);

BUFx3_ASAP7_75t_L g1684 ( 
.A(n_1657),
.Y(n_1684)
);

HB1xp67_ASAP7_75t_L g1685 ( 
.A(n_1671),
.Y(n_1685)
);

AND2x2_ASAP7_75t_L g1686 ( 
.A(n_1648),
.B(n_1627),
.Y(n_1686)
);

AND2x2_ASAP7_75t_L g1687 ( 
.A(n_1648),
.B(n_1644),
.Y(n_1687)
);

AND2x4_ASAP7_75t_L g1688 ( 
.A(n_1657),
.B(n_1667),
.Y(n_1688)
);

INVx1_ASAP7_75t_L g1689 ( 
.A(n_1647),
.Y(n_1689)
);

INVxp67_ASAP7_75t_L g1690 ( 
.A(n_1658),
.Y(n_1690)
);

HB1xp67_ASAP7_75t_L g1691 ( 
.A(n_1671),
.Y(n_1691)
);

BUFx2_ASAP7_75t_L g1692 ( 
.A(n_1672),
.Y(n_1692)
);

BUFx2_ASAP7_75t_L g1693 ( 
.A(n_1672),
.Y(n_1693)
);

OA21x2_ASAP7_75t_L g1694 ( 
.A1(n_1652),
.A2(n_1612),
.B(n_1640),
.Y(n_1694)
);

NAND2xp5_ASAP7_75t_L g1695 ( 
.A(n_1655),
.B(n_1598),
.Y(n_1695)
);

INVx3_ASAP7_75t_L g1696 ( 
.A(n_1653),
.Y(n_1696)
);

AND2x2_ASAP7_75t_L g1697 ( 
.A(n_1648),
.B(n_1598),
.Y(n_1697)
);

INVx1_ASAP7_75t_L g1698 ( 
.A(n_1647),
.Y(n_1698)
);

INVx3_ASAP7_75t_L g1699 ( 
.A(n_1653),
.Y(n_1699)
);

INVxp67_ASAP7_75t_SL g1700 ( 
.A(n_1652),
.Y(n_1700)
);

OR2x6_ASAP7_75t_L g1701 ( 
.A(n_1656),
.B(n_1622),
.Y(n_1701)
);

AND2x2_ASAP7_75t_L g1702 ( 
.A(n_1666),
.B(n_1639),
.Y(n_1702)
);

AOI22xp33_ASAP7_75t_L g1703 ( 
.A1(n_1662),
.A2(n_1606),
.B1(n_1632),
.B2(n_1597),
.Y(n_1703)
);

NAND3xp33_ASAP7_75t_L g1704 ( 
.A(n_1666),
.B(n_1599),
.C(n_1614),
.Y(n_1704)
);

HB1xp67_ASAP7_75t_L g1705 ( 
.A(n_1673),
.Y(n_1705)
);

HB1xp67_ASAP7_75t_L g1706 ( 
.A(n_1673),
.Y(n_1706)
);

HB1xp67_ASAP7_75t_L g1707 ( 
.A(n_1672),
.Y(n_1707)
);

INVx4_ASAP7_75t_L g1708 ( 
.A(n_1660),
.Y(n_1708)
);

INVxp67_ASAP7_75t_SL g1709 ( 
.A(n_1653),
.Y(n_1709)
);

NAND2xp5_ASAP7_75t_SL g1710 ( 
.A(n_1656),
.B(n_1628),
.Y(n_1710)
);

AOI21xp5_ASAP7_75t_L g1711 ( 
.A1(n_1666),
.A2(n_1640),
.B(n_1622),
.Y(n_1711)
);

NAND4xp25_ASAP7_75t_SL g1712 ( 
.A(n_1670),
.B(n_1599),
.C(n_1602),
.D(n_1620),
.Y(n_1712)
);

AND2x2_ASAP7_75t_L g1713 ( 
.A(n_1663),
.B(n_1642),
.Y(n_1713)
);

INVx2_ASAP7_75t_L g1714 ( 
.A(n_1677),
.Y(n_1714)
);

BUFx2_ASAP7_75t_L g1715 ( 
.A(n_1684),
.Y(n_1715)
);

AND2x2_ASAP7_75t_L g1716 ( 
.A(n_1684),
.B(n_1669),
.Y(n_1716)
);

HB1xp67_ASAP7_75t_L g1717 ( 
.A(n_1707),
.Y(n_1717)
);

NAND2xp5_ASAP7_75t_L g1718 ( 
.A(n_1686),
.B(n_1654),
.Y(n_1718)
);

INVx1_ASAP7_75t_L g1719 ( 
.A(n_1707),
.Y(n_1719)
);

AND2x2_ASAP7_75t_L g1720 ( 
.A(n_1684),
.B(n_1669),
.Y(n_1720)
);

INVx1_ASAP7_75t_L g1721 ( 
.A(n_1689),
.Y(n_1721)
);

INVx1_ASAP7_75t_L g1722 ( 
.A(n_1689),
.Y(n_1722)
);

AND2x2_ASAP7_75t_L g1723 ( 
.A(n_1686),
.B(n_1663),
.Y(n_1723)
);

INVx1_ASAP7_75t_L g1724 ( 
.A(n_1689),
.Y(n_1724)
);

OAI31xp33_ASAP7_75t_L g1725 ( 
.A1(n_1680),
.A2(n_1661),
.A3(n_1662),
.B(n_1665),
.Y(n_1725)
);

AND2x2_ASAP7_75t_L g1726 ( 
.A(n_1686),
.B(n_1663),
.Y(n_1726)
);

INVx1_ASAP7_75t_L g1727 ( 
.A(n_1698),
.Y(n_1727)
);

BUFx2_ASAP7_75t_L g1728 ( 
.A(n_1700),
.Y(n_1728)
);

NOR2x1_ASAP7_75t_L g1729 ( 
.A(n_1712),
.B(n_1625),
.Y(n_1729)
);

INVxp67_ASAP7_75t_SL g1730 ( 
.A(n_1700),
.Y(n_1730)
);

INVx2_ASAP7_75t_SL g1731 ( 
.A(n_1688),
.Y(n_1731)
);

AND2x2_ASAP7_75t_L g1732 ( 
.A(n_1702),
.B(n_1674),
.Y(n_1732)
);

OR2x2_ASAP7_75t_L g1733 ( 
.A(n_1685),
.B(n_1646),
.Y(n_1733)
);

AND2x2_ASAP7_75t_L g1734 ( 
.A(n_1702),
.B(n_1674),
.Y(n_1734)
);

NAND2xp5_ASAP7_75t_L g1735 ( 
.A(n_1687),
.B(n_1654),
.Y(n_1735)
);

HB1xp67_ASAP7_75t_L g1736 ( 
.A(n_1691),
.Y(n_1736)
);

NAND2xp5_ASAP7_75t_L g1737 ( 
.A(n_1687),
.B(n_1664),
.Y(n_1737)
);

AND2x2_ASAP7_75t_L g1738 ( 
.A(n_1713),
.B(n_1650),
.Y(n_1738)
);

NAND2xp5_ASAP7_75t_L g1739 ( 
.A(n_1690),
.B(n_1698),
.Y(n_1739)
);

NAND2xp5_ASAP7_75t_L g1740 ( 
.A(n_1690),
.B(n_1664),
.Y(n_1740)
);

INVx3_ASAP7_75t_L g1741 ( 
.A(n_1688),
.Y(n_1741)
);

OR2x6_ASAP7_75t_SL g1742 ( 
.A(n_1704),
.B(n_1618),
.Y(n_1742)
);

INVxp67_ASAP7_75t_SL g1743 ( 
.A(n_1709),
.Y(n_1743)
);

AND2x2_ASAP7_75t_L g1744 ( 
.A(n_1729),
.B(n_1697),
.Y(n_1744)
);

AND2x2_ASAP7_75t_L g1745 ( 
.A(n_1729),
.B(n_1697),
.Y(n_1745)
);

INVxp33_ASAP7_75t_L g1746 ( 
.A(n_1729),
.Y(n_1746)
);

AND2x4_ASAP7_75t_L g1747 ( 
.A(n_1731),
.B(n_1688),
.Y(n_1747)
);

INVx1_ASAP7_75t_L g1748 ( 
.A(n_1721),
.Y(n_1748)
);

NOR2x1_ASAP7_75t_L g1749 ( 
.A(n_1728),
.B(n_1712),
.Y(n_1749)
);

INVx1_ASAP7_75t_SL g1750 ( 
.A(n_1728),
.Y(n_1750)
);

AND2x2_ASAP7_75t_L g1751 ( 
.A(n_1723),
.B(n_1676),
.Y(n_1751)
);

NAND2xp5_ASAP7_75t_L g1752 ( 
.A(n_1730),
.B(n_1691),
.Y(n_1752)
);

AND2x2_ASAP7_75t_L g1753 ( 
.A(n_1723),
.B(n_1676),
.Y(n_1753)
);

INVxp67_ASAP7_75t_L g1754 ( 
.A(n_1742),
.Y(n_1754)
);

NAND2xp5_ASAP7_75t_L g1755 ( 
.A(n_1730),
.B(n_1705),
.Y(n_1755)
);

INVx1_ASAP7_75t_L g1756 ( 
.A(n_1721),
.Y(n_1756)
);

INVx1_ASAP7_75t_SL g1757 ( 
.A(n_1728),
.Y(n_1757)
);

NOR2xp67_ASAP7_75t_L g1758 ( 
.A(n_1741),
.B(n_1704),
.Y(n_1758)
);

INVx2_ASAP7_75t_SL g1759 ( 
.A(n_1715),
.Y(n_1759)
);

OAI222xp33_ASAP7_75t_L g1760 ( 
.A1(n_1723),
.A2(n_1703),
.B1(n_1678),
.B2(n_1711),
.C1(n_1683),
.C2(n_1681),
.Y(n_1760)
);

INVx1_ASAP7_75t_L g1761 ( 
.A(n_1721),
.Y(n_1761)
);

NAND2xp5_ASAP7_75t_L g1762 ( 
.A(n_1740),
.B(n_1705),
.Y(n_1762)
);

AND2x2_ASAP7_75t_L g1763 ( 
.A(n_1723),
.B(n_1676),
.Y(n_1763)
);

INVx1_ASAP7_75t_L g1764 ( 
.A(n_1722),
.Y(n_1764)
);

AND2x2_ASAP7_75t_L g1765 ( 
.A(n_1726),
.B(n_1679),
.Y(n_1765)
);

INVx2_ASAP7_75t_L g1766 ( 
.A(n_1714),
.Y(n_1766)
);

OAI211xp5_ASAP7_75t_SL g1767 ( 
.A1(n_1725),
.A2(n_1680),
.B(n_1696),
.C(n_1699),
.Y(n_1767)
);

AND2x2_ASAP7_75t_L g1768 ( 
.A(n_1726),
.B(n_1732),
.Y(n_1768)
);

INVx1_ASAP7_75t_L g1769 ( 
.A(n_1722),
.Y(n_1769)
);

INVx1_ASAP7_75t_L g1770 ( 
.A(n_1722),
.Y(n_1770)
);

INVx2_ASAP7_75t_L g1771 ( 
.A(n_1714),
.Y(n_1771)
);

NOR2x1_ASAP7_75t_L g1772 ( 
.A(n_1715),
.B(n_1710),
.Y(n_1772)
);

INVx1_ASAP7_75t_L g1773 ( 
.A(n_1724),
.Y(n_1773)
);

INVx1_ASAP7_75t_L g1774 ( 
.A(n_1724),
.Y(n_1774)
);

INVx2_ASAP7_75t_L g1775 ( 
.A(n_1714),
.Y(n_1775)
);

OR2x2_ASAP7_75t_L g1776 ( 
.A(n_1737),
.B(n_1706),
.Y(n_1776)
);

INVx1_ASAP7_75t_L g1777 ( 
.A(n_1724),
.Y(n_1777)
);

AND2x2_ASAP7_75t_L g1778 ( 
.A(n_1726),
.B(n_1679),
.Y(n_1778)
);

NAND2xp5_ASAP7_75t_L g1779 ( 
.A(n_1740),
.B(n_1706),
.Y(n_1779)
);

INVx1_ASAP7_75t_L g1780 ( 
.A(n_1727),
.Y(n_1780)
);

INVx1_ASAP7_75t_L g1781 ( 
.A(n_1727),
.Y(n_1781)
);

NAND2xp5_ASAP7_75t_L g1782 ( 
.A(n_1736),
.B(n_1681),
.Y(n_1782)
);

NAND2xp5_ASAP7_75t_L g1783 ( 
.A(n_1736),
.B(n_1681),
.Y(n_1783)
);

NOR2x1p5_ASAP7_75t_L g1784 ( 
.A(n_1741),
.B(n_1708),
.Y(n_1784)
);

INVx1_ASAP7_75t_L g1785 ( 
.A(n_1727),
.Y(n_1785)
);

AND2x2_ASAP7_75t_L g1786 ( 
.A(n_1726),
.B(n_1679),
.Y(n_1786)
);

HB1xp67_ASAP7_75t_L g1787 ( 
.A(n_1739),
.Y(n_1787)
);

INVx2_ASAP7_75t_L g1788 ( 
.A(n_1714),
.Y(n_1788)
);

AND2x2_ASAP7_75t_L g1789 ( 
.A(n_1732),
.B(n_1734),
.Y(n_1789)
);

BUFx2_ASAP7_75t_L g1790 ( 
.A(n_1749),
.Y(n_1790)
);

INVx1_ASAP7_75t_L g1791 ( 
.A(n_1748),
.Y(n_1791)
);

OR2x2_ASAP7_75t_L g1792 ( 
.A(n_1762),
.B(n_1779),
.Y(n_1792)
);

INVx1_ASAP7_75t_L g1793 ( 
.A(n_1748),
.Y(n_1793)
);

AND2x2_ASAP7_75t_L g1794 ( 
.A(n_1749),
.B(n_1742),
.Y(n_1794)
);

INVx1_ASAP7_75t_L g1795 ( 
.A(n_1756),
.Y(n_1795)
);

HB1xp67_ASAP7_75t_L g1796 ( 
.A(n_1787),
.Y(n_1796)
);

INVx2_ASAP7_75t_L g1797 ( 
.A(n_1766),
.Y(n_1797)
);

OR2x2_ASAP7_75t_L g1798 ( 
.A(n_1762),
.B(n_1718),
.Y(n_1798)
);

NAND2xp5_ASAP7_75t_L g1799 ( 
.A(n_1750),
.B(n_1717),
.Y(n_1799)
);

AND2x2_ASAP7_75t_L g1800 ( 
.A(n_1746),
.B(n_1742),
.Y(n_1800)
);

AND2x2_ASAP7_75t_L g1801 ( 
.A(n_1744),
.B(n_1742),
.Y(n_1801)
);

INVxp67_ASAP7_75t_L g1802 ( 
.A(n_1754),
.Y(n_1802)
);

INVx1_ASAP7_75t_L g1803 ( 
.A(n_1756),
.Y(n_1803)
);

AND2x2_ASAP7_75t_L g1804 ( 
.A(n_1744),
.B(n_1738),
.Y(n_1804)
);

INVx2_ASAP7_75t_L g1805 ( 
.A(n_1766),
.Y(n_1805)
);

INVx1_ASAP7_75t_SL g1806 ( 
.A(n_1750),
.Y(n_1806)
);

OR2x2_ASAP7_75t_L g1807 ( 
.A(n_1779),
.B(n_1718),
.Y(n_1807)
);

INVx1_ASAP7_75t_L g1808 ( 
.A(n_1761),
.Y(n_1808)
);

HB1xp67_ASAP7_75t_L g1809 ( 
.A(n_1757),
.Y(n_1809)
);

AND2x2_ASAP7_75t_L g1810 ( 
.A(n_1745),
.B(n_1738),
.Y(n_1810)
);

AND2x2_ASAP7_75t_L g1811 ( 
.A(n_1745),
.B(n_1738),
.Y(n_1811)
);

OR2x2_ASAP7_75t_L g1812 ( 
.A(n_1776),
.B(n_1733),
.Y(n_1812)
);

AOI22xp33_ASAP7_75t_L g1813 ( 
.A1(n_1767),
.A2(n_1682),
.B1(n_1703),
.B2(n_1678),
.Y(n_1813)
);

NAND2xp5_ASAP7_75t_L g1814 ( 
.A(n_1757),
.B(n_1717),
.Y(n_1814)
);

HB1xp67_ASAP7_75t_L g1815 ( 
.A(n_1759),
.Y(n_1815)
);

NOR2xp33_ASAP7_75t_L g1816 ( 
.A(n_1760),
.B(n_1600),
.Y(n_1816)
);

NAND2xp5_ASAP7_75t_L g1817 ( 
.A(n_1752),
.B(n_1737),
.Y(n_1817)
);

INVx3_ASAP7_75t_L g1818 ( 
.A(n_1747),
.Y(n_1818)
);

AND2x2_ASAP7_75t_L g1819 ( 
.A(n_1768),
.B(n_1738),
.Y(n_1819)
);

INVx1_ASAP7_75t_L g1820 ( 
.A(n_1761),
.Y(n_1820)
);

INVx1_ASAP7_75t_L g1821 ( 
.A(n_1764),
.Y(n_1821)
);

INVx1_ASAP7_75t_L g1822 ( 
.A(n_1764),
.Y(n_1822)
);

INVx1_ASAP7_75t_L g1823 ( 
.A(n_1769),
.Y(n_1823)
);

OR2x2_ASAP7_75t_L g1824 ( 
.A(n_1776),
.B(n_1733),
.Y(n_1824)
);

INVx1_ASAP7_75t_L g1825 ( 
.A(n_1769),
.Y(n_1825)
);

NAND2xp5_ASAP7_75t_L g1826 ( 
.A(n_1752),
.B(n_1739),
.Y(n_1826)
);

AO22x1_ASAP7_75t_L g1827 ( 
.A1(n_1790),
.A2(n_1772),
.B1(n_1743),
.B2(n_1747),
.Y(n_1827)
);

INVx1_ASAP7_75t_L g1828 ( 
.A(n_1791),
.Y(n_1828)
);

INVx1_ASAP7_75t_L g1829 ( 
.A(n_1791),
.Y(n_1829)
);

AOI32xp33_ASAP7_75t_L g1830 ( 
.A1(n_1790),
.A2(n_1783),
.A3(n_1782),
.B1(n_1683),
.B2(n_1772),
.Y(n_1830)
);

NOR2xp33_ASAP7_75t_L g1831 ( 
.A(n_1816),
.B(n_1675),
.Y(n_1831)
);

OAI22xp5_ASAP7_75t_L g1832 ( 
.A1(n_1794),
.A2(n_1758),
.B1(n_1782),
.B2(n_1783),
.Y(n_1832)
);

INVx1_ASAP7_75t_L g1833 ( 
.A(n_1793),
.Y(n_1833)
);

INVx1_ASAP7_75t_L g1834 ( 
.A(n_1793),
.Y(n_1834)
);

NAND2xp5_ASAP7_75t_L g1835 ( 
.A(n_1806),
.B(n_1789),
.Y(n_1835)
);

INVx1_ASAP7_75t_L g1836 ( 
.A(n_1795),
.Y(n_1836)
);

NOR2xp33_ASAP7_75t_SL g1837 ( 
.A(n_1794),
.B(n_1725),
.Y(n_1837)
);

INVx1_ASAP7_75t_L g1838 ( 
.A(n_1795),
.Y(n_1838)
);

AOI22xp5_ASAP7_75t_L g1839 ( 
.A1(n_1813),
.A2(n_1682),
.B1(n_1683),
.B2(n_1758),
.Y(n_1839)
);

AOI22xp5_ASAP7_75t_L g1840 ( 
.A1(n_1801),
.A2(n_1597),
.B1(n_1711),
.B2(n_1701),
.Y(n_1840)
);

INVx1_ASAP7_75t_L g1841 ( 
.A(n_1803),
.Y(n_1841)
);

NAND4xp25_ASAP7_75t_L g1842 ( 
.A(n_1802),
.B(n_1755),
.C(n_1715),
.D(n_1768),
.Y(n_1842)
);

INVx1_ASAP7_75t_L g1843 ( 
.A(n_1803),
.Y(n_1843)
);

AOI21xp33_ASAP7_75t_L g1844 ( 
.A1(n_1800),
.A2(n_1826),
.B(n_1820),
.Y(n_1844)
);

NAND2xp5_ASAP7_75t_L g1845 ( 
.A(n_1806),
.B(n_1789),
.Y(n_1845)
);

AOI22xp5_ASAP7_75t_L g1846 ( 
.A1(n_1801),
.A2(n_1701),
.B1(n_1694),
.B2(n_1753),
.Y(n_1846)
);

INVx1_ASAP7_75t_L g1847 ( 
.A(n_1808),
.Y(n_1847)
);

NAND2xp5_ASAP7_75t_L g1848 ( 
.A(n_1796),
.B(n_1751),
.Y(n_1848)
);

OAI221xp5_ASAP7_75t_SL g1849 ( 
.A1(n_1800),
.A2(n_1755),
.B1(n_1701),
.B2(n_1765),
.C(n_1786),
.Y(n_1849)
);

INVx1_ASAP7_75t_SL g1850 ( 
.A(n_1809),
.Y(n_1850)
);

AOI21xp33_ASAP7_75t_L g1851 ( 
.A1(n_1826),
.A2(n_1759),
.B(n_1766),
.Y(n_1851)
);

AOI22xp5_ASAP7_75t_L g1852 ( 
.A1(n_1804),
.A2(n_1810),
.B1(n_1811),
.B2(n_1805),
.Y(n_1852)
);

AOI22xp5_ASAP7_75t_L g1853 ( 
.A1(n_1804),
.A2(n_1701),
.B1(n_1694),
.B2(n_1763),
.Y(n_1853)
);

INVx2_ASAP7_75t_L g1854 ( 
.A(n_1850),
.Y(n_1854)
);

AOI221xp5_ASAP7_75t_L g1855 ( 
.A1(n_1837),
.A2(n_1844),
.B1(n_1839),
.B2(n_1842),
.C(n_1832),
.Y(n_1855)
);

NOR2xp33_ASAP7_75t_L g1856 ( 
.A(n_1831),
.B(n_1792),
.Y(n_1856)
);

AOI221xp5_ASAP7_75t_L g1857 ( 
.A1(n_1842),
.A2(n_1817),
.B1(n_1805),
.B2(n_1797),
.C(n_1692),
.Y(n_1857)
);

AOI22xp5_ASAP7_75t_L g1858 ( 
.A1(n_1840),
.A2(n_1797),
.B1(n_1805),
.B2(n_1692),
.Y(n_1858)
);

NAND4xp25_ASAP7_75t_L g1859 ( 
.A(n_1830),
.B(n_1799),
.C(n_1814),
.D(n_1818),
.Y(n_1859)
);

OAI221xp5_ASAP7_75t_L g1860 ( 
.A1(n_1846),
.A2(n_1817),
.B1(n_1807),
.B2(n_1798),
.C(n_1792),
.Y(n_1860)
);

O2A1O1Ixp33_ASAP7_75t_L g1861 ( 
.A1(n_1851),
.A2(n_1849),
.B(n_1829),
.C(n_1833),
.Y(n_1861)
);

INVx2_ASAP7_75t_L g1862 ( 
.A(n_1827),
.Y(n_1862)
);

AND2x4_ASAP7_75t_L g1863 ( 
.A(n_1835),
.B(n_1818),
.Y(n_1863)
);

HB1xp67_ASAP7_75t_L g1864 ( 
.A(n_1845),
.Y(n_1864)
);

NAND2xp5_ASAP7_75t_L g1865 ( 
.A(n_1848),
.B(n_1815),
.Y(n_1865)
);

OAI22xp5_ASAP7_75t_L g1866 ( 
.A1(n_1852),
.A2(n_1810),
.B1(n_1811),
.B2(n_1818),
.Y(n_1866)
);

INVx1_ASAP7_75t_L g1867 ( 
.A(n_1828),
.Y(n_1867)
);

INVx1_ASAP7_75t_L g1868 ( 
.A(n_1834),
.Y(n_1868)
);

AOI21xp5_ASAP7_75t_L g1869 ( 
.A1(n_1836),
.A2(n_1814),
.B(n_1799),
.Y(n_1869)
);

INVxp67_ASAP7_75t_L g1870 ( 
.A(n_1838),
.Y(n_1870)
);

OAI22xp5_ASAP7_75t_L g1871 ( 
.A1(n_1853),
.A2(n_1818),
.B1(n_1731),
.B2(n_1819),
.Y(n_1871)
);

OR2x6_ASAP7_75t_L g1872 ( 
.A(n_1841),
.B(n_1617),
.Y(n_1872)
);

INVx2_ASAP7_75t_L g1873 ( 
.A(n_1843),
.Y(n_1873)
);

NOR4xp25_ASAP7_75t_SL g1874 ( 
.A(n_1847),
.B(n_1825),
.C(n_1808),
.D(n_1823),
.Y(n_1874)
);

OAI21xp5_ASAP7_75t_SL g1875 ( 
.A1(n_1855),
.A2(n_1819),
.B(n_1747),
.Y(n_1875)
);

INVx1_ASAP7_75t_L g1876 ( 
.A(n_1854),
.Y(n_1876)
);

NAND2xp5_ASAP7_75t_L g1877 ( 
.A(n_1856),
.B(n_1751),
.Y(n_1877)
);

INVx2_ASAP7_75t_SL g1878 ( 
.A(n_1872),
.Y(n_1878)
);

INVx1_ASAP7_75t_L g1879 ( 
.A(n_1867),
.Y(n_1879)
);

OR2x2_ASAP7_75t_L g1880 ( 
.A(n_1864),
.B(n_1798),
.Y(n_1880)
);

AOI22xp5_ASAP7_75t_L g1881 ( 
.A1(n_1862),
.A2(n_1797),
.B1(n_1693),
.B2(n_1692),
.Y(n_1881)
);

OR2x2_ASAP7_75t_L g1882 ( 
.A(n_1859),
.B(n_1807),
.Y(n_1882)
);

NAND2xp5_ASAP7_75t_L g1883 ( 
.A(n_1863),
.B(n_1753),
.Y(n_1883)
);

NAND2xp5_ASAP7_75t_L g1884 ( 
.A(n_1863),
.B(n_1763),
.Y(n_1884)
);

INVx1_ASAP7_75t_L g1885 ( 
.A(n_1868),
.Y(n_1885)
);

INVx1_ASAP7_75t_L g1886 ( 
.A(n_1873),
.Y(n_1886)
);

NAND3xp33_ASAP7_75t_L g1887 ( 
.A(n_1876),
.B(n_1874),
.C(n_1857),
.Y(n_1887)
);

NAND3xp33_ASAP7_75t_SL g1888 ( 
.A(n_1875),
.B(n_1861),
.C(n_1858),
.Y(n_1888)
);

NOR3xp33_ASAP7_75t_L g1889 ( 
.A(n_1878),
.B(n_1860),
.C(n_1870),
.Y(n_1889)
);

NOR3xp33_ASAP7_75t_SL g1890 ( 
.A(n_1886),
.B(n_1866),
.C(n_1865),
.Y(n_1890)
);

NAND2xp5_ASAP7_75t_L g1891 ( 
.A(n_1877),
.B(n_1869),
.Y(n_1891)
);

INVx2_ASAP7_75t_L g1892 ( 
.A(n_1880),
.Y(n_1892)
);

AND2x2_ASAP7_75t_L g1893 ( 
.A(n_1883),
.B(n_1872),
.Y(n_1893)
);

NAND2xp5_ASAP7_75t_L g1894 ( 
.A(n_1884),
.B(n_1765),
.Y(n_1894)
);

NAND4xp25_ASAP7_75t_L g1895 ( 
.A(n_1882),
.B(n_1871),
.C(n_1858),
.D(n_1812),
.Y(n_1895)
);

NAND3xp33_ASAP7_75t_L g1896 ( 
.A(n_1879),
.B(n_1821),
.C(n_1820),
.Y(n_1896)
);

AOI22xp5_ASAP7_75t_L g1897 ( 
.A1(n_1881),
.A2(n_1778),
.B1(n_1786),
.B2(n_1771),
.Y(n_1897)
);

NAND2xp5_ASAP7_75t_L g1898 ( 
.A(n_1885),
.B(n_1778),
.Y(n_1898)
);

NAND2xp5_ASAP7_75t_L g1899 ( 
.A(n_1892),
.B(n_1881),
.Y(n_1899)
);

AOI221xp5_ASAP7_75t_L g1900 ( 
.A1(n_1887),
.A2(n_1825),
.B1(n_1823),
.B2(n_1822),
.C(n_1821),
.Y(n_1900)
);

OAI211xp5_ASAP7_75t_L g1901 ( 
.A1(n_1890),
.A2(n_1743),
.B(n_1812),
.C(n_1824),
.Y(n_1901)
);

AOI222xp33_ASAP7_75t_L g1902 ( 
.A1(n_1888),
.A2(n_1822),
.B1(n_1693),
.B2(n_1788),
.C1(n_1771),
.C2(n_1775),
.Y(n_1902)
);

OAI211xp5_ASAP7_75t_L g1903 ( 
.A1(n_1895),
.A2(n_1824),
.B(n_1741),
.C(n_1731),
.Y(n_1903)
);

AOI221xp5_ASAP7_75t_L g1904 ( 
.A1(n_1889),
.A2(n_1788),
.B1(n_1771),
.B2(n_1775),
.C(n_1693),
.Y(n_1904)
);

INVx1_ASAP7_75t_L g1905 ( 
.A(n_1899),
.Y(n_1905)
);

OAI211xp5_ASAP7_75t_L g1906 ( 
.A1(n_1901),
.A2(n_1891),
.B(n_1893),
.C(n_1897),
.Y(n_1906)
);

INVx1_ASAP7_75t_L g1907 ( 
.A(n_1902),
.Y(n_1907)
);

AOI22xp5_ASAP7_75t_L g1908 ( 
.A1(n_1900),
.A2(n_1898),
.B1(n_1894),
.B2(n_1896),
.Y(n_1908)
);

OAI21xp33_ASAP7_75t_SL g1909 ( 
.A1(n_1904),
.A2(n_1784),
.B(n_1731),
.Y(n_1909)
);

NAND3xp33_ASAP7_75t_SL g1910 ( 
.A(n_1903),
.B(n_1710),
.C(n_1775),
.Y(n_1910)
);

AOI221xp5_ASAP7_75t_L g1911 ( 
.A1(n_1900),
.A2(n_1788),
.B1(n_1719),
.B2(n_1716),
.C(n_1720),
.Y(n_1911)
);

XNOR2xp5_ASAP7_75t_L g1912 ( 
.A(n_1905),
.B(n_1784),
.Y(n_1912)
);

NOR2x1_ASAP7_75t_L g1913 ( 
.A(n_1906),
.B(n_1747),
.Y(n_1913)
);

BUFx2_ASAP7_75t_L g1914 ( 
.A(n_1909),
.Y(n_1914)
);

NOR4xp75_ASAP7_75t_L g1915 ( 
.A(n_1910),
.B(n_1741),
.C(n_1735),
.D(n_1695),
.Y(n_1915)
);

AND2x2_ASAP7_75t_L g1916 ( 
.A(n_1908),
.B(n_1741),
.Y(n_1916)
);

OR2x2_ASAP7_75t_L g1917 ( 
.A(n_1914),
.B(n_1907),
.Y(n_1917)
);

HB1xp67_ASAP7_75t_L g1918 ( 
.A(n_1913),
.Y(n_1918)
);

AND2x4_ASAP7_75t_L g1919 ( 
.A(n_1916),
.B(n_1741),
.Y(n_1919)
);

XOR2x1_ASAP7_75t_L g1920 ( 
.A(n_1918),
.B(n_1912),
.Y(n_1920)
);

INVx1_ASAP7_75t_L g1921 ( 
.A(n_1920),
.Y(n_1921)
);

OAI22xp5_ASAP7_75t_SL g1922 ( 
.A1(n_1921),
.A2(n_1917),
.B1(n_1919),
.B2(n_1915),
.Y(n_1922)
);

NAND2xp5_ASAP7_75t_L g1923 ( 
.A(n_1921),
.B(n_1911),
.Y(n_1923)
);

OAI21xp33_ASAP7_75t_L g1924 ( 
.A1(n_1923),
.A2(n_1773),
.B(n_1770),
.Y(n_1924)
);

OAI22xp5_ASAP7_75t_L g1925 ( 
.A1(n_1922),
.A2(n_1785),
.B1(n_1781),
.B2(n_1780),
.Y(n_1925)
);

INVx1_ASAP7_75t_L g1926 ( 
.A(n_1925),
.Y(n_1926)
);

AOI21xp5_ASAP7_75t_L g1927 ( 
.A1(n_1924),
.A2(n_1719),
.B(n_1785),
.Y(n_1927)
);

HB1xp67_ASAP7_75t_L g1928 ( 
.A(n_1926),
.Y(n_1928)
);

AOI221xp5_ASAP7_75t_L g1929 ( 
.A1(n_1928),
.A2(n_1927),
.B1(n_1719),
.B2(n_1780),
.C(n_1777),
.Y(n_1929)
);

INVx1_ASAP7_75t_L g1930 ( 
.A(n_1929),
.Y(n_1930)
);

OAI221xp5_ASAP7_75t_R g1931 ( 
.A1(n_1930),
.A2(n_1604),
.B1(n_1777),
.B2(n_1774),
.C(n_1773),
.Y(n_1931)
);

AOI211xp5_ASAP7_75t_L g1932 ( 
.A1(n_1931),
.A2(n_1675),
.B(n_1628),
.C(n_1770),
.Y(n_1932)
);


endmodule