module fake_netlist_6_2943_n_553 (n_16, n_1, n_9, n_8, n_18, n_10, n_21, n_24, n_6, n_15, n_3, n_14, n_0, n_4, n_22, n_13, n_11, n_17, n_23, n_12, n_20, n_7, n_2, n_5, n_19, n_553);

input n_16;
input n_1;
input n_9;
input n_8;
input n_18;
input n_10;
input n_21;
input n_24;
input n_6;
input n_15;
input n_3;
input n_14;
input n_0;
input n_4;
input n_22;
input n_13;
input n_11;
input n_17;
input n_23;
input n_12;
input n_20;
input n_7;
input n_2;
input n_5;
input n_19;

output n_553;

wire n_52;
wire n_435;
wire n_91;
wire n_326;
wire n_256;
wire n_440;
wire n_507;
wire n_209;
wire n_367;
wire n_465;
wire n_63;
wire n_223;
wire n_278;
wire n_341;
wire n_362;
wire n_148;
wire n_226;
wire n_161;
wire n_208;
wire n_462;
wire n_68;
wire n_316;
wire n_419;
wire n_28;
wire n_304;
wire n_212;
wire n_50;
wire n_144;
wire n_365;
wire n_125;
wire n_168;
wire n_384;
wire n_297;
wire n_524;
wire n_342;
wire n_77;
wire n_106;
wire n_358;
wire n_160;
wire n_449;
wire n_131;
wire n_188;
wire n_310;
wire n_509;
wire n_186;
wire n_245;
wire n_368;
wire n_396;
wire n_495;
wire n_350;
wire n_78;
wire n_84;
wire n_392;
wire n_442;
wire n_480;
wire n_142;
wire n_143;
wire n_382;
wire n_180;
wire n_62;
wire n_349;
wire n_233;
wire n_255;
wire n_284;
wire n_400;
wire n_140;
wire n_337;
wire n_214;
wire n_485;
wire n_67;
wire n_443;
wire n_246;
wire n_38;
wire n_471;
wire n_289;
wire n_421;
wire n_424;
wire n_59;
wire n_181;
wire n_182;
wire n_238;
wire n_202;
wire n_320;
wire n_108;
wire n_327;
wire n_369;
wire n_280;
wire n_287;
wire n_353;
wire n_389;
wire n_415;
wire n_65;
wire n_230;
wire n_461;
wire n_141;
wire n_383;
wire n_200;
wire n_447;
wire n_176;
wire n_114;
wire n_86;
wire n_198;
wire n_104;
wire n_300;
wire n_179;
wire n_248;
wire n_222;
wire n_517;
wire n_71;
wire n_74;
wire n_229;
wire n_542;
wire n_305;
wire n_72;
wire n_532;
wire n_173;
wire n_535;
wire n_250;
wire n_372;
wire n_468;
wire n_544;
wire n_111;
wire n_504;
wire n_314;
wire n_378;
wire n_413;
wire n_377;
wire n_35;
wire n_183;
wire n_510;
wire n_79;
wire n_375;
wire n_338;
wire n_522;
wire n_466;
wire n_506;
wire n_56;
wire n_360;
wire n_119;
wire n_235;
wire n_536;
wire n_147;
wire n_191;
wire n_340;
wire n_387;
wire n_452;
wire n_39;
wire n_344;
wire n_73;
wire n_428;
wire n_432;
wire n_101;
wire n_167;
wire n_174;
wire n_127;
wire n_516;
wire n_153;
wire n_525;
wire n_156;
wire n_491;
wire n_145;
wire n_42;
wire n_133;
wire n_96;
wire n_371;
wire n_189;
wire n_405;
wire n_213;
wire n_538;
wire n_294;
wire n_302;
wire n_499;
wire n_380;
wire n_129;
wire n_197;
wire n_137;
wire n_343;
wire n_448;
wire n_494;
wire n_539;
wire n_493;
wire n_397;
wire n_155;
wire n_109;
wire n_529;
wire n_445;
wire n_425;
wire n_122;
wire n_45;
wire n_454;
wire n_34;
wire n_218;
wire n_70;
wire n_234;
wire n_37;
wire n_486;
wire n_381;
wire n_82;
wire n_27;
wire n_236;
wire n_112;
wire n_172;
wire n_472;
wire n_270;
wire n_239;
wire n_126;
wire n_414;
wire n_97;
wire n_58;
wire n_490;
wire n_290;
wire n_220;
wire n_118;
wire n_224;
wire n_48;
wire n_25;
wire n_93;
wire n_80;
wire n_196;
wire n_402;
wire n_352;
wire n_478;
wire n_460;
wire n_107;
wire n_417;
wire n_446;
wire n_498;
wire n_89;
wire n_374;
wire n_366;
wire n_407;
wire n_450;
wire n_103;
wire n_272;
wire n_526;
wire n_185;
wire n_348;
wire n_69;
wire n_376;
wire n_390;
wire n_473;
wire n_293;
wire n_31;
wire n_334;
wire n_53;
wire n_370;
wire n_44;
wire n_458;
wire n_232;
wire n_163;
wire n_46;
wire n_330;
wire n_470;
wire n_475;
wire n_298;
wire n_492;
wire n_281;
wire n_258;
wire n_551;
wire n_154;
wire n_456;
wire n_98;
wire n_260;
wire n_265;
wire n_313;
wire n_451;
wire n_279;
wire n_252;
wire n_228;
wire n_356;
wire n_166;
wire n_184;
wire n_552;
wire n_216;
wire n_455;
wire n_83;
wire n_521;
wire n_363;
wire n_395;
wire n_323;
wire n_393;
wire n_411;
wire n_503;
wire n_152;
wire n_92;
wire n_513;
wire n_321;
wire n_331;
wire n_105;
wire n_227;
wire n_132;
wire n_406;
wire n_483;
wire n_102;
wire n_204;
wire n_482;
wire n_474;
wire n_527;
wire n_261;
wire n_420;
wire n_394;
wire n_312;
wire n_32;
wire n_66;
wire n_130;
wire n_519;
wire n_541;
wire n_512;
wire n_164;
wire n_292;
wire n_100;
wire n_121;
wire n_307;
wire n_469;
wire n_433;
wire n_500;
wire n_476;
wire n_291;
wire n_219;
wire n_543;
wire n_357;
wire n_150;
wire n_264;
wire n_263;
wire n_481;
wire n_325;
wire n_329;
wire n_464;
wire n_33;
wire n_477;
wire n_549;
wire n_533;
wire n_408;
wire n_61;
wire n_237;
wire n_244;
wire n_399;
wire n_76;
wire n_243;
wire n_124;
wire n_548;
wire n_94;
wire n_282;
wire n_436;
wire n_116;
wire n_211;
wire n_523;
wire n_117;
wire n_175;
wire n_322;
wire n_409;
wire n_345;
wire n_231;
wire n_354;
wire n_40;
wire n_505;
wire n_240;
wire n_139;
wire n_319;
wire n_41;
wire n_134;
wire n_547;
wire n_537;
wire n_273;
wire n_95;
wire n_311;
wire n_403;
wire n_253;
wire n_123;
wire n_136;
wire n_546;
wire n_249;
wire n_201;
wire n_386;
wire n_159;
wire n_157;
wire n_162;
wire n_115;
wire n_487;
wire n_550;
wire n_128;
wire n_241;
wire n_30;
wire n_275;
wire n_43;
wire n_276;
wire n_441;
wire n_221;
wire n_444;
wire n_423;
wire n_146;
wire n_318;
wire n_303;
wire n_511;
wire n_467;
wire n_306;
wire n_193;
wire n_269;
wire n_359;
wire n_346;
wire n_88;
wire n_416;
wire n_530;
wire n_277;
wire n_520;
wire n_418;
wire n_113;
wire n_199;
wire n_138;
wire n_266;
wire n_296;
wire n_268;
wire n_404;
wire n_271;
wire n_439;
wire n_158;
wire n_217;
wire n_49;
wire n_210;
wire n_299;
wire n_518;
wire n_206;
wire n_453;
wire n_333;
wire n_215;
wire n_178;
wire n_247;
wire n_225;
wire n_308;
wire n_309;
wire n_355;
wire n_426;
wire n_317;
wire n_149;
wire n_431;
wire n_90;
wire n_347;
wire n_459;
wire n_54;
wire n_502;
wire n_328;
wire n_534;
wire n_488;
wire n_429;
wire n_373;
wire n_87;
wire n_195;
wire n_285;
wire n_497;
wire n_85;
wire n_99;
wire n_257;
wire n_203;
wire n_286;
wire n_254;
wire n_207;
wire n_242;
wire n_47;
wire n_29;
wire n_75;
wire n_401;
wire n_324;
wire n_335;
wire n_430;
wire n_463;
wire n_545;
wire n_489;
wire n_205;
wire n_120;
wire n_251;
wire n_301;
wire n_274;
wire n_110;
wire n_151;
wire n_412;
wire n_81;
wire n_36;
wire n_26;
wire n_55;
wire n_267;
wire n_438;
wire n_339;
wire n_434;
wire n_515;
wire n_315;
wire n_64;
wire n_288;
wire n_427;
wire n_479;
wire n_496;
wire n_422;
wire n_135;
wire n_165;
wire n_351;
wire n_437;
wire n_259;
wire n_177;
wire n_540;
wire n_514;
wire n_528;
wire n_391;
wire n_457;
wire n_364;
wire n_295;
wire n_385;
wire n_388;
wire n_190;
wire n_484;
wire n_262;
wire n_187;
wire n_501;
wire n_531;
wire n_60;
wire n_361;
wire n_508;
wire n_379;
wire n_170;
wire n_332;
wire n_336;
wire n_410;
wire n_398;
wire n_194;
wire n_171;
wire n_192;
wire n_57;
wire n_169;
wire n_51;
wire n_283;

INVx1_ASAP7_75t_L g25 ( 
.A(n_15),
.Y(n_25)
);

CKINVDCx5p33_ASAP7_75t_R g26 ( 
.A(n_15),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_13),
.Y(n_27)
);

CKINVDCx5p33_ASAP7_75t_R g28 ( 
.A(n_22),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_23),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_6),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_0),
.Y(n_31)
);

INVx2_ASAP7_75t_L g32 ( 
.A(n_18),
.Y(n_32)
);

BUFx3_ASAP7_75t_L g33 ( 
.A(n_16),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_1),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_12),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_4),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_24),
.Y(n_37)
);

NOR2xp67_ASAP7_75t_L g38 ( 
.A(n_21),
.B(n_4),
.Y(n_38)
);

CKINVDCx5p33_ASAP7_75t_R g39 ( 
.A(n_0),
.Y(n_39)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_12),
.Y(n_40)
);

CKINVDCx5p33_ASAP7_75t_R g41 ( 
.A(n_11),
.Y(n_41)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_17),
.Y(n_42)
);

BUFx3_ASAP7_75t_L g43 ( 
.A(n_17),
.Y(n_43)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_14),
.Y(n_44)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_8),
.Y(n_45)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_6),
.Y(n_46)
);

INVx2_ASAP7_75t_L g47 ( 
.A(n_3),
.Y(n_47)
);

CKINVDCx5p33_ASAP7_75t_R g48 ( 
.A(n_13),
.Y(n_48)
);

HB1xp67_ASAP7_75t_L g49 ( 
.A(n_18),
.Y(n_49)
);

INVx2_ASAP7_75t_L g50 ( 
.A(n_35),
.Y(n_50)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_35),
.Y(n_51)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_35),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_L g53 ( 
.A(n_32),
.B(n_1),
.Y(n_53)
);

INVx5_ASAP7_75t_L g54 ( 
.A(n_35),
.Y(n_54)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_35),
.Y(n_55)
);

OAI21x1_ASAP7_75t_L g56 ( 
.A1(n_32),
.A2(n_2),
.B(n_3),
.Y(n_56)
);

HB1xp67_ASAP7_75t_L g57 ( 
.A(n_49),
.Y(n_57)
);

AND2x4_ASAP7_75t_L g58 ( 
.A(n_35),
.B(n_20),
.Y(n_58)
);

INVx3_ASAP7_75t_L g59 ( 
.A(n_35),
.Y(n_59)
);

CKINVDCx16_ASAP7_75t_R g60 ( 
.A(n_37),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_L g61 ( 
.A(n_32),
.B(n_2),
.Y(n_61)
);

AND2x6_ASAP7_75t_L g62 ( 
.A(n_29),
.B(n_19),
.Y(n_62)
);

OR2x2_ASAP7_75t_L g63 ( 
.A(n_57),
.B(n_49),
.Y(n_63)
);

INVx2_ASAP7_75t_L g64 ( 
.A(n_50),
.Y(n_64)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_51),
.Y(n_65)
);

AND2x2_ASAP7_75t_L g66 ( 
.A(n_59),
.B(n_33),
.Y(n_66)
);

NAND2xp33_ASAP7_75t_L g67 ( 
.A(n_62),
.B(n_35),
.Y(n_67)
);

AOI22xp33_ASAP7_75t_L g68 ( 
.A1(n_62),
.A2(n_33),
.B1(n_43),
.B2(n_32),
.Y(n_68)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_51),
.Y(n_69)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_50),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_53),
.B(n_43),
.Y(n_71)
);

INVx3_ASAP7_75t_L g72 ( 
.A(n_58),
.Y(n_72)
);

INVx2_ASAP7_75t_L g73 ( 
.A(n_50),
.Y(n_73)
);

INVx2_ASAP7_75t_SL g74 ( 
.A(n_58),
.Y(n_74)
);

INVx1_ASAP7_75t_SL g75 ( 
.A(n_60),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_SL g76 ( 
.A(n_58),
.B(n_38),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_53),
.B(n_43),
.Y(n_77)
);

INVx2_ASAP7_75t_SL g78 ( 
.A(n_58),
.Y(n_78)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_51),
.Y(n_79)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_52),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_L g81 ( 
.A(n_59),
.B(n_33),
.Y(n_81)
);

AOI22xp5_ASAP7_75t_L g82 ( 
.A1(n_71),
.A2(n_37),
.B1(n_62),
.B2(n_39),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_L g83 ( 
.A(n_66),
.B(n_59),
.Y(n_83)
);

NAND2x1_ASAP7_75t_L g84 ( 
.A(n_68),
.B(n_62),
.Y(n_84)
);

BUFx3_ASAP7_75t_L g85 ( 
.A(n_66),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_L g86 ( 
.A(n_66),
.B(n_59),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_L g87 ( 
.A(n_74),
.B(n_59),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_SL g88 ( 
.A(n_68),
.B(n_60),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_74),
.B(n_59),
.Y(n_89)
);

AND2x2_ASAP7_75t_L g90 ( 
.A(n_71),
.B(n_61),
.Y(n_90)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_65),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_SL g92 ( 
.A(n_74),
.B(n_77),
.Y(n_92)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_65),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_L g94 ( 
.A(n_78),
.B(n_55),
.Y(n_94)
);

AOI22xp33_ASAP7_75t_L g95 ( 
.A1(n_76),
.A2(n_77),
.B1(n_62),
.B2(n_72),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_76),
.B(n_60),
.Y(n_96)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_65),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_SL g98 ( 
.A(n_78),
.B(n_63),
.Y(n_98)
);

AOI22xp33_ASAP7_75t_L g99 ( 
.A1(n_72),
.A2(n_62),
.B1(n_78),
.B2(n_67),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_SL g100 ( 
.A(n_78),
.B(n_28),
.Y(n_100)
);

INVxp67_ASAP7_75t_L g101 ( 
.A(n_63),
.Y(n_101)
);

INVx2_ASAP7_75t_L g102 ( 
.A(n_64),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_SL g103 ( 
.A(n_63),
.B(n_58),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_L g104 ( 
.A(n_69),
.B(n_55),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_L g105 ( 
.A(n_69),
.B(n_55),
.Y(n_105)
);

OAI221xp5_ASAP7_75t_L g106 ( 
.A1(n_81),
.A2(n_53),
.B1(n_61),
.B2(n_47),
.C(n_42),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_L g107 ( 
.A(n_69),
.B(n_80),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_SL g108 ( 
.A(n_72),
.B(n_58),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_SL g109 ( 
.A(n_72),
.B(n_75),
.Y(n_109)
);

OAI22xp33_ASAP7_75t_L g110 ( 
.A1(n_75),
.A2(n_57),
.B1(n_61),
.B2(n_26),
.Y(n_110)
);

AOI22xp5_ASAP7_75t_L g111 ( 
.A1(n_67),
.A2(n_62),
.B1(n_41),
.B2(n_39),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_L g112 ( 
.A(n_72),
.B(n_48),
.Y(n_112)
);

NAND3xp33_ASAP7_75t_L g113 ( 
.A(n_81),
.B(n_47),
.C(n_52),
.Y(n_113)
);

AND2x2_ASAP7_75t_L g114 ( 
.A(n_72),
.B(n_80),
.Y(n_114)
);

HB1xp67_ASAP7_75t_L g115 ( 
.A(n_79),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_L g116 ( 
.A(n_79),
.B(n_52),
.Y(n_116)
);

AOI21xp5_ASAP7_75t_L g117 ( 
.A1(n_108),
.A2(n_80),
.B(n_79),
.Y(n_117)
);

INVxp67_ASAP7_75t_SL g118 ( 
.A(n_85),
.Y(n_118)
);

A2O1A1Ixp33_ASAP7_75t_L g119 ( 
.A1(n_90),
.A2(n_56),
.B(n_47),
.C(n_25),
.Y(n_119)
);

O2A1O1Ixp33_ASAP7_75t_L g120 ( 
.A1(n_106),
.A2(n_47),
.B(n_40),
.C(n_36),
.Y(n_120)
);

INVx2_ASAP7_75t_L g121 ( 
.A(n_85),
.Y(n_121)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_85),
.Y(n_122)
);

O2A1O1Ixp33_ASAP7_75t_L g123 ( 
.A1(n_98),
.A2(n_103),
.B(n_88),
.C(n_92),
.Y(n_123)
);

NOR2x1_ASAP7_75t_L g124 ( 
.A(n_96),
.B(n_38),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_L g125 ( 
.A(n_90),
.B(n_41),
.Y(n_125)
);

AND2x2_ASAP7_75t_L g126 ( 
.A(n_101),
.B(n_33),
.Y(n_126)
);

AOI221xp5_ASAP7_75t_L g127 ( 
.A1(n_110),
.A2(n_44),
.B1(n_42),
.B2(n_40),
.C(n_46),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_L g128 ( 
.A(n_112),
.B(n_62),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_L g129 ( 
.A(n_115),
.B(n_62),
.Y(n_129)
);

AOI21xp5_ASAP7_75t_L g130 ( 
.A1(n_83),
.A2(n_73),
.B(n_70),
.Y(n_130)
);

O2A1O1Ixp33_ASAP7_75t_L g131 ( 
.A1(n_109),
.A2(n_31),
.B(n_27),
.C(n_46),
.Y(n_131)
);

AOI21xp5_ASAP7_75t_L g132 ( 
.A1(n_83),
.A2(n_73),
.B(n_70),
.Y(n_132)
);

AND2x2_ASAP7_75t_L g133 ( 
.A(n_82),
.B(n_43),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_SL g134 ( 
.A(n_82),
.B(n_29),
.Y(n_134)
);

AOI21xp5_ASAP7_75t_L g135 ( 
.A1(n_86),
.A2(n_73),
.B(n_70),
.Y(n_135)
);

AOI21xp5_ASAP7_75t_L g136 ( 
.A1(n_86),
.A2(n_89),
.B(n_87),
.Y(n_136)
);

AOI21xp5_ASAP7_75t_L g137 ( 
.A1(n_87),
.A2(n_64),
.B(n_54),
.Y(n_137)
);

AO32x1_ASAP7_75t_L g138 ( 
.A1(n_91),
.A2(n_30),
.A3(n_25),
.B1(n_27),
.B2(n_45),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_L g139 ( 
.A(n_114),
.B(n_62),
.Y(n_139)
);

AOI21xp5_ASAP7_75t_L g140 ( 
.A1(n_89),
.A2(n_64),
.B(n_54),
.Y(n_140)
);

AND2x2_ASAP7_75t_L g141 ( 
.A(n_114),
.B(n_31),
.Y(n_141)
);

AO32x1_ASAP7_75t_L g142 ( 
.A1(n_91),
.A2(n_30),
.A3(n_45),
.B1(n_44),
.B2(n_36),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_SL g143 ( 
.A(n_99),
.B(n_50),
.Y(n_143)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_93),
.Y(n_144)
);

HB1xp67_ASAP7_75t_L g145 ( 
.A(n_100),
.Y(n_145)
);

A2O1A1Ixp33_ASAP7_75t_L g146 ( 
.A1(n_84),
.A2(n_56),
.B(n_34),
.C(n_64),
.Y(n_146)
);

INVxp67_ASAP7_75t_L g147 ( 
.A(n_113),
.Y(n_147)
);

AOI22xp5_ASAP7_75t_L g148 ( 
.A1(n_95),
.A2(n_62),
.B1(n_34),
.B2(n_56),
.Y(n_148)
);

A2O1A1Ixp33_ASAP7_75t_L g149 ( 
.A1(n_84),
.A2(n_56),
.B(n_62),
.C(n_54),
.Y(n_149)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_93),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_L g151 ( 
.A(n_97),
.B(n_54),
.Y(n_151)
);

BUFx2_ASAP7_75t_L g152 ( 
.A(n_97),
.Y(n_152)
);

NOR2x1p5_ASAP7_75t_SL g153 ( 
.A(n_102),
.B(n_54),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_L g154 ( 
.A(n_94),
.B(n_107),
.Y(n_154)
);

OAI22xp5_ASAP7_75t_L g155 ( 
.A1(n_111),
.A2(n_54),
.B1(n_7),
.B2(n_8),
.Y(n_155)
);

AO21x1_ASAP7_75t_L g156 ( 
.A1(n_111),
.A2(n_5),
.B(n_7),
.Y(n_156)
);

OAI21xp5_ASAP7_75t_L g157 ( 
.A1(n_113),
.A2(n_54),
.B(n_9),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_L g158 ( 
.A(n_107),
.B(n_54),
.Y(n_158)
);

BUFx2_ASAP7_75t_L g159 ( 
.A(n_104),
.Y(n_159)
);

NOR2xp33_ASAP7_75t_R g160 ( 
.A(n_104),
.B(n_5),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_SL g161 ( 
.A(n_116),
.B(n_54),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_L g162 ( 
.A(n_116),
.B(n_54),
.Y(n_162)
);

O2A1O1Ixp33_ASAP7_75t_SL g163 ( 
.A1(n_105),
.A2(n_9),
.B(n_10),
.C(n_11),
.Y(n_163)
);

OAI21x1_ASAP7_75t_L g164 ( 
.A1(n_105),
.A2(n_10),
.B(n_14),
.Y(n_164)
);

AOI21xp5_ASAP7_75t_L g165 ( 
.A1(n_102),
.A2(n_16),
.B(n_19),
.Y(n_165)
);

A2O1A1Ixp33_ASAP7_75t_L g166 ( 
.A1(n_125),
.A2(n_123),
.B(n_120),
.C(n_134),
.Y(n_166)
);

AO31x2_ASAP7_75t_L g167 ( 
.A1(n_119),
.A2(n_102),
.A3(n_146),
.B(n_149),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_L g168 ( 
.A(n_159),
.B(n_154),
.Y(n_168)
);

AOI21xp5_ASAP7_75t_L g169 ( 
.A1(n_136),
.A2(n_118),
.B(n_139),
.Y(n_169)
);

INVx2_ASAP7_75t_L g170 ( 
.A(n_121),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_L g171 ( 
.A(n_125),
.B(n_141),
.Y(n_171)
);

NOR2xp33_ASAP7_75t_L g172 ( 
.A(n_145),
.B(n_152),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_SL g173 ( 
.A(n_121),
.B(n_124),
.Y(n_173)
);

INVx2_ASAP7_75t_SL g174 ( 
.A(n_122),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_L g175 ( 
.A(n_144),
.B(n_150),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_L g176 ( 
.A(n_147),
.B(n_133),
.Y(n_176)
);

AOI21xp5_ASAP7_75t_L g177 ( 
.A1(n_129),
.A2(n_128),
.B(n_143),
.Y(n_177)
);

AND2x4_ASAP7_75t_L g178 ( 
.A(n_153),
.B(n_126),
.Y(n_178)
);

AOI21xp5_ASAP7_75t_SL g179 ( 
.A1(n_149),
.A2(n_146),
.B(n_119),
.Y(n_179)
);

AND2x2_ASAP7_75t_L g180 ( 
.A(n_134),
.B(n_143),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_L g181 ( 
.A(n_117),
.B(n_131),
.Y(n_181)
);

OR2x2_ASAP7_75t_L g182 ( 
.A(n_155),
.B(n_161),
.Y(n_182)
);

NAND2xp33_ASAP7_75t_L g183 ( 
.A(n_157),
.B(n_148),
.Y(n_183)
);

OAI22xp5_ASAP7_75t_L g184 ( 
.A1(n_158),
.A2(n_161),
.B1(n_127),
.B2(n_151),
.Y(n_184)
);

OAI21xp5_ASAP7_75t_L g185 ( 
.A1(n_130),
.A2(n_132),
.B(n_135),
.Y(n_185)
);

AOI21xp5_ASAP7_75t_SL g186 ( 
.A1(n_162),
.A2(n_137),
.B(n_140),
.Y(n_186)
);

BUFx3_ASAP7_75t_L g187 ( 
.A(n_164),
.Y(n_187)
);

AOI221xp5_ASAP7_75t_L g188 ( 
.A1(n_156),
.A2(n_163),
.B1(n_160),
.B2(n_165),
.C(n_138),
.Y(n_188)
);

AOI21xp5_ASAP7_75t_L g189 ( 
.A1(n_138),
.A2(n_142),
.B(n_163),
.Y(n_189)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_160),
.Y(n_190)
);

AO31x2_ASAP7_75t_L g191 ( 
.A1(n_138),
.A2(n_119),
.A3(n_146),
.B(n_149),
.Y(n_191)
);

AOI21xp5_ASAP7_75t_SL g192 ( 
.A1(n_138),
.A2(n_78),
.B(n_74),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_L g193 ( 
.A(n_142),
.B(n_90),
.Y(n_193)
);

NAND3x1_ASAP7_75t_L g194 ( 
.A(n_142),
.B(n_127),
.C(n_82),
.Y(n_194)
);

AOI21xp5_ASAP7_75t_L g195 ( 
.A1(n_154),
.A2(n_74),
.B(n_78),
.Y(n_195)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_122),
.Y(n_196)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_122),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_L g198 ( 
.A(n_159),
.B(n_90),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_L g199 ( 
.A(n_159),
.B(n_90),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_L g200 ( 
.A(n_159),
.B(n_90),
.Y(n_200)
);

AND2x2_ASAP7_75t_L g201 ( 
.A(n_159),
.B(n_90),
.Y(n_201)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_122),
.Y(n_202)
);

NAND2xp5_ASAP7_75t_L g203 ( 
.A(n_159),
.B(n_90),
.Y(n_203)
);

AO31x2_ASAP7_75t_L g204 ( 
.A1(n_119),
.A2(n_146),
.A3(n_149),
.B(n_156),
.Y(n_204)
);

HB1xp67_ASAP7_75t_L g205 ( 
.A(n_141),
.Y(n_205)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_122),
.Y(n_206)
);

AND2x2_ASAP7_75t_L g207 ( 
.A(n_159),
.B(n_90),
.Y(n_207)
);

AOI21xp5_ASAP7_75t_L g208 ( 
.A1(n_154),
.A2(n_74),
.B(n_78),
.Y(n_208)
);

OAI21x1_ASAP7_75t_L g209 ( 
.A1(n_179),
.A2(n_189),
.B(n_185),
.Y(n_209)
);

BUFx6f_ASAP7_75t_L g210 ( 
.A(n_187),
.Y(n_210)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_170),
.Y(n_211)
);

OAI21x1_ASAP7_75t_SL g212 ( 
.A1(n_169),
.A2(n_177),
.B(n_171),
.Y(n_212)
);

NAND2xp5_ASAP7_75t_SL g213 ( 
.A(n_168),
.B(n_201),
.Y(n_213)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_170),
.Y(n_214)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_175),
.Y(n_215)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_180),
.Y(n_216)
);

NAND2xp5_ASAP7_75t_L g217 ( 
.A(n_201),
.B(n_207),
.Y(n_217)
);

OA21x2_ASAP7_75t_L g218 ( 
.A1(n_193),
.A2(n_166),
.B(n_188),
.Y(n_218)
);

NAND2xp5_ASAP7_75t_SL g219 ( 
.A(n_207),
.B(n_203),
.Y(n_219)
);

AO31x2_ASAP7_75t_L g220 ( 
.A1(n_166),
.A2(n_184),
.A3(n_176),
.B(n_195),
.Y(n_220)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_180),
.Y(n_221)
);

AO21x2_ASAP7_75t_L g222 ( 
.A1(n_183),
.A2(n_173),
.B(n_192),
.Y(n_222)
);

OAI21x1_ASAP7_75t_L g223 ( 
.A1(n_208),
.A2(n_186),
.B(n_173),
.Y(n_223)
);

INVx2_ASAP7_75t_L g224 ( 
.A(n_167),
.Y(n_224)
);

INVx3_ASAP7_75t_L g225 ( 
.A(n_167),
.Y(n_225)
);

INVx2_ASAP7_75t_L g226 ( 
.A(n_167),
.Y(n_226)
);

BUFx6f_ASAP7_75t_L g227 ( 
.A(n_187),
.Y(n_227)
);

NAND2xp5_ASAP7_75t_L g228 ( 
.A(n_198),
.B(n_199),
.Y(n_228)
);

AND2x2_ASAP7_75t_L g229 ( 
.A(n_205),
.B(n_200),
.Y(n_229)
);

OR2x6_ASAP7_75t_L g230 ( 
.A(n_182),
.B(n_178),
.Y(n_230)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_167),
.Y(n_231)
);

OAI21x1_ASAP7_75t_L g232 ( 
.A1(n_194),
.A2(n_181),
.B(n_182),
.Y(n_232)
);

OR2x2_ASAP7_75t_L g233 ( 
.A(n_190),
.B(n_172),
.Y(n_233)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_196),
.Y(n_234)
);

OR2x2_ASAP7_75t_L g235 ( 
.A(n_197),
.B(n_206),
.Y(n_235)
);

INVx2_ASAP7_75t_L g236 ( 
.A(n_191),
.Y(n_236)
);

BUFx6f_ASAP7_75t_L g237 ( 
.A(n_178),
.Y(n_237)
);

OR2x2_ASAP7_75t_L g238 ( 
.A(n_202),
.B(n_174),
.Y(n_238)
);

NAND2xp5_ASAP7_75t_L g239 ( 
.A(n_183),
.B(n_174),
.Y(n_239)
);

NAND2xp5_ASAP7_75t_L g240 ( 
.A(n_178),
.B(n_204),
.Y(n_240)
);

OAI21x1_ASAP7_75t_L g241 ( 
.A1(n_194),
.A2(n_191),
.B(n_204),
.Y(n_241)
);

NAND2xp5_ASAP7_75t_SL g242 ( 
.A(n_204),
.B(n_191),
.Y(n_242)
);

OAI21x1_ASAP7_75t_L g243 ( 
.A1(n_204),
.A2(n_179),
.B(n_189),
.Y(n_243)
);

OAI21x1_ASAP7_75t_L g244 ( 
.A1(n_179),
.A2(n_189),
.B(n_185),
.Y(n_244)
);

BUFx2_ASAP7_75t_L g245 ( 
.A(n_205),
.Y(n_245)
);

INVx2_ASAP7_75t_L g246 ( 
.A(n_170),
.Y(n_246)
);

CKINVDCx5p33_ASAP7_75t_R g247 ( 
.A(n_172),
.Y(n_247)
);

OAI21x1_ASAP7_75t_L g248 ( 
.A1(n_179),
.A2(n_189),
.B(n_185),
.Y(n_248)
);

OAI21x1_ASAP7_75t_L g249 ( 
.A1(n_179),
.A2(n_189),
.B(n_185),
.Y(n_249)
);

OR2x2_ASAP7_75t_L g250 ( 
.A(n_176),
.B(n_168),
.Y(n_250)
);

OAI21x1_ASAP7_75t_SL g251 ( 
.A1(n_169),
.A2(n_156),
.B(n_123),
.Y(n_251)
);

INVx2_ASAP7_75t_L g252 ( 
.A(n_170),
.Y(n_252)
);

NAND2xp5_ASAP7_75t_L g253 ( 
.A(n_215),
.B(n_228),
.Y(n_253)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_246),
.Y(n_254)
);

INVx2_ASAP7_75t_L g255 ( 
.A(n_252),
.Y(n_255)
);

NAND2xp5_ASAP7_75t_L g256 ( 
.A(n_215),
.B(n_228),
.Y(n_256)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_252),
.Y(n_257)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_211),
.Y(n_258)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_211),
.Y(n_259)
);

AND2x2_ASAP7_75t_L g260 ( 
.A(n_216),
.B(n_221),
.Y(n_260)
);

INVx2_ASAP7_75t_L g261 ( 
.A(n_225),
.Y(n_261)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_214),
.Y(n_262)
);

AO21x2_ASAP7_75t_L g263 ( 
.A1(n_212),
.A2(n_251),
.B(n_209),
.Y(n_263)
);

NAND3xp33_ASAP7_75t_SL g264 ( 
.A(n_247),
.B(n_250),
.C(n_233),
.Y(n_264)
);

INVx3_ASAP7_75t_L g265 ( 
.A(n_237),
.Y(n_265)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_214),
.Y(n_266)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_224),
.Y(n_267)
);

AND2x4_ASAP7_75t_L g268 ( 
.A(n_230),
.B(n_237),
.Y(n_268)
);

BUFx2_ASAP7_75t_L g269 ( 
.A(n_230),
.Y(n_269)
);

INVx2_ASAP7_75t_SL g270 ( 
.A(n_237),
.Y(n_270)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_216),
.Y(n_271)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_221),
.Y(n_272)
);

BUFx6f_ASAP7_75t_L g273 ( 
.A(n_227),
.Y(n_273)
);

OA21x2_ASAP7_75t_L g274 ( 
.A1(n_209),
.A2(n_249),
.B(n_248),
.Y(n_274)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_225),
.Y(n_275)
);

NAND2xp5_ASAP7_75t_L g276 ( 
.A(n_250),
.B(n_217),
.Y(n_276)
);

INVx4_ASAP7_75t_L g277 ( 
.A(n_227),
.Y(n_277)
);

AOI21x1_ASAP7_75t_L g278 ( 
.A1(n_212),
.A2(n_251),
.B(n_223),
.Y(n_278)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_224),
.Y(n_279)
);

INVx2_ASAP7_75t_L g280 ( 
.A(n_224),
.Y(n_280)
);

AND2x4_ASAP7_75t_L g281 ( 
.A(n_230),
.B(n_237),
.Y(n_281)
);

INVx2_ASAP7_75t_L g282 ( 
.A(n_226),
.Y(n_282)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_226),
.Y(n_283)
);

INVx2_ASAP7_75t_L g284 ( 
.A(n_226),
.Y(n_284)
);

NAND2xp5_ASAP7_75t_L g285 ( 
.A(n_217),
.B(n_213),
.Y(n_285)
);

BUFx2_ASAP7_75t_L g286 ( 
.A(n_230),
.Y(n_286)
);

BUFx2_ASAP7_75t_L g287 ( 
.A(n_230),
.Y(n_287)
);

INVx2_ASAP7_75t_L g288 ( 
.A(n_209),
.Y(n_288)
);

NAND2xp5_ASAP7_75t_L g289 ( 
.A(n_253),
.B(n_231),
.Y(n_289)
);

AND2x2_ASAP7_75t_L g290 ( 
.A(n_267),
.B(n_231),
.Y(n_290)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_267),
.Y(n_291)
);

AND2x2_ASAP7_75t_L g292 ( 
.A(n_267),
.B(n_241),
.Y(n_292)
);

NAND2xp5_ASAP7_75t_L g293 ( 
.A(n_253),
.B(n_239),
.Y(n_293)
);

INVxp67_ASAP7_75t_SL g294 ( 
.A(n_280),
.Y(n_294)
);

HB1xp67_ASAP7_75t_L g295 ( 
.A(n_261),
.Y(n_295)
);

BUFx3_ASAP7_75t_L g296 ( 
.A(n_268),
.Y(n_296)
);

AO21x2_ASAP7_75t_L g297 ( 
.A1(n_278),
.A2(n_249),
.B(n_244),
.Y(n_297)
);

OAI22xp33_ASAP7_75t_L g298 ( 
.A1(n_256),
.A2(n_233),
.B1(n_230),
.B2(n_235),
.Y(n_298)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_279),
.Y(n_299)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_279),
.Y(n_300)
);

AND2x2_ASAP7_75t_L g301 ( 
.A(n_280),
.B(n_241),
.Y(n_301)
);

INVxp67_ASAP7_75t_L g302 ( 
.A(n_256),
.Y(n_302)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_283),
.Y(n_303)
);

AND2x4_ASAP7_75t_L g304 ( 
.A(n_268),
.B(n_227),
.Y(n_304)
);

AND2x2_ASAP7_75t_L g305 ( 
.A(n_280),
.B(n_241),
.Y(n_305)
);

HB1xp67_ASAP7_75t_L g306 ( 
.A(n_261),
.Y(n_306)
);

HB1xp67_ASAP7_75t_L g307 ( 
.A(n_261),
.Y(n_307)
);

AND2x2_ASAP7_75t_L g308 ( 
.A(n_282),
.B(n_236),
.Y(n_308)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_283),
.Y(n_309)
);

AND2x2_ASAP7_75t_L g310 ( 
.A(n_282),
.B(n_236),
.Y(n_310)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_282),
.Y(n_311)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_284),
.Y(n_312)
);

OA21x2_ASAP7_75t_L g313 ( 
.A1(n_288),
.A2(n_249),
.B(n_248),
.Y(n_313)
);

AND2x2_ASAP7_75t_L g314 ( 
.A(n_284),
.B(n_236),
.Y(n_314)
);

INVx2_ASAP7_75t_L g315 ( 
.A(n_284),
.Y(n_315)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_291),
.Y(n_316)
);

AND2x2_ASAP7_75t_L g317 ( 
.A(n_301),
.B(n_305),
.Y(n_317)
);

AND2x2_ASAP7_75t_L g318 ( 
.A(n_301),
.B(n_274),
.Y(n_318)
);

INVx3_ASAP7_75t_L g319 ( 
.A(n_313),
.Y(n_319)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_291),
.Y(n_320)
);

INVx3_ASAP7_75t_L g321 ( 
.A(n_313),
.Y(n_321)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_291),
.Y(n_322)
);

HB1xp67_ASAP7_75t_L g323 ( 
.A(n_295),
.Y(n_323)
);

AND2x4_ASAP7_75t_L g324 ( 
.A(n_296),
.B(n_269),
.Y(n_324)
);

OR2x2_ASAP7_75t_L g325 ( 
.A(n_297),
.B(n_274),
.Y(n_325)
);

AND2x2_ASAP7_75t_L g326 ( 
.A(n_301),
.B(n_274),
.Y(n_326)
);

AND2x2_ASAP7_75t_L g327 ( 
.A(n_301),
.B(n_274),
.Y(n_327)
);

BUFx2_ASAP7_75t_SL g328 ( 
.A(n_294),
.Y(n_328)
);

NAND2xp5_ASAP7_75t_L g329 ( 
.A(n_302),
.B(n_293),
.Y(n_329)
);

AND2x4_ASAP7_75t_L g330 ( 
.A(n_296),
.B(n_269),
.Y(n_330)
);

INVx2_ASAP7_75t_L g331 ( 
.A(n_313),
.Y(n_331)
);

AND2x2_ASAP7_75t_L g332 ( 
.A(n_305),
.B(n_274),
.Y(n_332)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_292),
.Y(n_333)
);

AND2x2_ASAP7_75t_L g334 ( 
.A(n_305),
.B(n_274),
.Y(n_334)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_292),
.Y(n_335)
);

NOR2xp33_ASAP7_75t_L g336 ( 
.A(n_302),
.B(n_264),
.Y(n_336)
);

AND2x2_ASAP7_75t_L g337 ( 
.A(n_305),
.B(n_288),
.Y(n_337)
);

INVx1_ASAP7_75t_L g338 ( 
.A(n_292),
.Y(n_338)
);

INVx3_ASAP7_75t_SL g339 ( 
.A(n_304),
.Y(n_339)
);

INVx2_ASAP7_75t_L g340 ( 
.A(n_313),
.Y(n_340)
);

AND2x4_ASAP7_75t_SL g341 ( 
.A(n_304),
.B(n_281),
.Y(n_341)
);

INVx2_ASAP7_75t_SL g342 ( 
.A(n_296),
.Y(n_342)
);

AND2x2_ASAP7_75t_L g343 ( 
.A(n_292),
.B(n_288),
.Y(n_343)
);

INVx2_ASAP7_75t_L g344 ( 
.A(n_313),
.Y(n_344)
);

NAND2x1p5_ASAP7_75t_L g345 ( 
.A(n_313),
.B(n_244),
.Y(n_345)
);

NAND2xp5_ASAP7_75t_L g346 ( 
.A(n_293),
.B(n_276),
.Y(n_346)
);

OR2x2_ASAP7_75t_L g347 ( 
.A(n_297),
.B(n_288),
.Y(n_347)
);

BUFx2_ASAP7_75t_L g348 ( 
.A(n_342),
.Y(n_348)
);

OR2x2_ASAP7_75t_L g349 ( 
.A(n_317),
.B(n_297),
.Y(n_349)
);

NAND2xp5_ASAP7_75t_L g350 ( 
.A(n_329),
.B(n_289),
.Y(n_350)
);

INVx1_ASAP7_75t_L g351 ( 
.A(n_316),
.Y(n_351)
);

INVx2_ASAP7_75t_L g352 ( 
.A(n_316),
.Y(n_352)
);

INVx1_ASAP7_75t_L g353 ( 
.A(n_320),
.Y(n_353)
);

INVx1_ASAP7_75t_L g354 ( 
.A(n_320),
.Y(n_354)
);

INVx1_ASAP7_75t_L g355 ( 
.A(n_322),
.Y(n_355)
);

INVx1_ASAP7_75t_L g356 ( 
.A(n_322),
.Y(n_356)
);

INVx2_ASAP7_75t_L g357 ( 
.A(n_331),
.Y(n_357)
);

OR2x2_ASAP7_75t_L g358 ( 
.A(n_317),
.B(n_297),
.Y(n_358)
);

NAND2xp5_ASAP7_75t_L g359 ( 
.A(n_329),
.B(n_289),
.Y(n_359)
);

INVx1_ASAP7_75t_L g360 ( 
.A(n_335),
.Y(n_360)
);

NAND3xp33_ASAP7_75t_L g361 ( 
.A(n_336),
.B(n_219),
.C(n_285),
.Y(n_361)
);

INVx1_ASAP7_75t_L g362 ( 
.A(n_335),
.Y(n_362)
);

NAND2x1_ASAP7_75t_L g363 ( 
.A(n_324),
.B(n_299),
.Y(n_363)
);

AND2x2_ASAP7_75t_L g364 ( 
.A(n_317),
.B(n_296),
.Y(n_364)
);

AND2x2_ASAP7_75t_L g365 ( 
.A(n_335),
.B(n_313),
.Y(n_365)
);

AND2x2_ASAP7_75t_L g366 ( 
.A(n_318),
.B(n_297),
.Y(n_366)
);

INVx1_ASAP7_75t_L g367 ( 
.A(n_333),
.Y(n_367)
);

INVx1_ASAP7_75t_L g368 ( 
.A(n_333),
.Y(n_368)
);

INVx2_ASAP7_75t_SL g369 ( 
.A(n_341),
.Y(n_369)
);

INVx1_ASAP7_75t_L g370 ( 
.A(n_338),
.Y(n_370)
);

OR2x2_ASAP7_75t_L g371 ( 
.A(n_338),
.B(n_297),
.Y(n_371)
);

INVx1_ASAP7_75t_L g372 ( 
.A(n_323),
.Y(n_372)
);

INVx4_ASAP7_75t_L g373 ( 
.A(n_339),
.Y(n_373)
);

NAND2xp5_ASAP7_75t_L g374 ( 
.A(n_336),
.B(n_298),
.Y(n_374)
);

HB1xp67_ASAP7_75t_L g375 ( 
.A(n_323),
.Y(n_375)
);

NOR2xp33_ASAP7_75t_L g376 ( 
.A(n_346),
.B(n_264),
.Y(n_376)
);

OR2x2_ASAP7_75t_L g377 ( 
.A(n_318),
.B(n_263),
.Y(n_377)
);

AND2x2_ASAP7_75t_L g378 ( 
.A(n_318),
.B(n_269),
.Y(n_378)
);

INVx1_ASAP7_75t_L g379 ( 
.A(n_328),
.Y(n_379)
);

INVx1_ASAP7_75t_L g380 ( 
.A(n_360),
.Y(n_380)
);

AND2x2_ASAP7_75t_L g381 ( 
.A(n_366),
.B(n_326),
.Y(n_381)
);

OR2x2_ASAP7_75t_L g382 ( 
.A(n_349),
.B(n_326),
.Y(n_382)
);

NAND2xp5_ASAP7_75t_L g383 ( 
.A(n_376),
.B(n_298),
.Y(n_383)
);

INVx1_ASAP7_75t_L g384 ( 
.A(n_355),
.Y(n_384)
);

NAND2xp5_ASAP7_75t_L g385 ( 
.A(n_374),
.B(n_346),
.Y(n_385)
);

NOR2xp33_ASAP7_75t_L g386 ( 
.A(n_361),
.B(n_339),
.Y(n_386)
);

INVxp67_ASAP7_75t_L g387 ( 
.A(n_375),
.Y(n_387)
);

AND2x2_ASAP7_75t_L g388 ( 
.A(n_366),
.B(n_326),
.Y(n_388)
);

INVxp67_ASAP7_75t_L g389 ( 
.A(n_350),
.Y(n_389)
);

NAND2x1p5_ASAP7_75t_L g390 ( 
.A(n_373),
.B(n_342),
.Y(n_390)
);

AND2x2_ASAP7_75t_L g391 ( 
.A(n_364),
.B(n_327),
.Y(n_391)
);

OR2x2_ASAP7_75t_L g392 ( 
.A(n_349),
.B(n_327),
.Y(n_392)
);

INVxp67_ASAP7_75t_SL g393 ( 
.A(n_379),
.Y(n_393)
);

INVx1_ASAP7_75t_L g394 ( 
.A(n_355),
.Y(n_394)
);

AND2x2_ASAP7_75t_L g395 ( 
.A(n_364),
.B(n_327),
.Y(n_395)
);

AOI21xp33_ASAP7_75t_SL g396 ( 
.A1(n_359),
.A2(n_339),
.B(n_276),
.Y(n_396)
);

NAND2xp67_ASAP7_75t_L g397 ( 
.A(n_352),
.B(n_260),
.Y(n_397)
);

AND2x2_ASAP7_75t_L g398 ( 
.A(n_378),
.B(n_332),
.Y(n_398)
);

OR2x2_ASAP7_75t_L g399 ( 
.A(n_358),
.B(n_332),
.Y(n_399)
);

INVx1_ASAP7_75t_L g400 ( 
.A(n_360),
.Y(n_400)
);

NAND2xp5_ASAP7_75t_L g401 ( 
.A(n_378),
.B(n_324),
.Y(n_401)
);

NOR2xp33_ASAP7_75t_L g402 ( 
.A(n_369),
.B(n_339),
.Y(n_402)
);

INVx1_ASAP7_75t_L g403 ( 
.A(n_356),
.Y(n_403)
);

INVx1_ASAP7_75t_L g404 ( 
.A(n_356),
.Y(n_404)
);

AND2x2_ASAP7_75t_L g405 ( 
.A(n_358),
.B(n_332),
.Y(n_405)
);

NAND2xp5_ASAP7_75t_L g406 ( 
.A(n_372),
.B(n_324),
.Y(n_406)
);

OR2x2_ASAP7_75t_L g407 ( 
.A(n_377),
.B(n_371),
.Y(n_407)
);

NAND2xp5_ASAP7_75t_L g408 ( 
.A(n_351),
.B(n_353),
.Y(n_408)
);

INVx1_ASAP7_75t_L g409 ( 
.A(n_362),
.Y(n_409)
);

A2O1A1Ixp33_ASAP7_75t_L g410 ( 
.A1(n_363),
.A2(n_244),
.B(n_248),
.C(n_341),
.Y(n_410)
);

INVx1_ASAP7_75t_L g411 ( 
.A(n_380),
.Y(n_411)
);

INVxp67_ASAP7_75t_L g412 ( 
.A(n_387),
.Y(n_412)
);

AOI21xp33_ASAP7_75t_SL g413 ( 
.A1(n_385),
.A2(n_369),
.B(n_377),
.Y(n_413)
);

AOI21xp33_ASAP7_75t_L g414 ( 
.A1(n_383),
.A2(n_363),
.B(n_371),
.Y(n_414)
);

INVx1_ASAP7_75t_SL g415 ( 
.A(n_391),
.Y(n_415)
);

INVx1_ASAP7_75t_L g416 ( 
.A(n_380),
.Y(n_416)
);

INVx1_ASAP7_75t_L g417 ( 
.A(n_400),
.Y(n_417)
);

OAI22xp33_ASAP7_75t_L g418 ( 
.A1(n_389),
.A2(n_373),
.B1(n_287),
.B2(n_286),
.Y(n_418)
);

INVx1_ASAP7_75t_L g419 ( 
.A(n_400),
.Y(n_419)
);

INVx2_ASAP7_75t_L g420 ( 
.A(n_409),
.Y(n_420)
);

AOI21xp5_ASAP7_75t_L g421 ( 
.A1(n_410),
.A2(n_268),
.B(n_281),
.Y(n_421)
);

AOI211xp5_ASAP7_75t_L g422 ( 
.A1(n_386),
.A2(n_396),
.B(n_393),
.C(n_402),
.Y(n_422)
);

AOI22xp5_ASAP7_75t_L g423 ( 
.A1(n_406),
.A2(n_330),
.B1(n_324),
.B2(n_304),
.Y(n_423)
);

INVx1_ASAP7_75t_L g424 ( 
.A(n_384),
.Y(n_424)
);

INVx1_ASAP7_75t_L g425 ( 
.A(n_394),
.Y(n_425)
);

AOI21xp5_ASAP7_75t_L g426 ( 
.A1(n_390),
.A2(n_268),
.B(n_281),
.Y(n_426)
);

OAI22xp5_ASAP7_75t_L g427 ( 
.A1(n_401),
.A2(n_342),
.B1(n_373),
.B2(n_324),
.Y(n_427)
);

INVx1_ASAP7_75t_L g428 ( 
.A(n_403),
.Y(n_428)
);

AOI22xp33_ASAP7_75t_L g429 ( 
.A1(n_404),
.A2(n_287),
.B1(n_286),
.B2(n_285),
.Y(n_429)
);

INVx1_ASAP7_75t_L g430 ( 
.A(n_408),
.Y(n_430)
);

AND2x4_ASAP7_75t_L g431 ( 
.A(n_391),
.B(n_362),
.Y(n_431)
);

OAI22xp33_ASAP7_75t_L g432 ( 
.A1(n_382),
.A2(n_287),
.B1(n_286),
.B2(n_345),
.Y(n_432)
);

INVx1_ASAP7_75t_L g433 ( 
.A(n_407),
.Y(n_433)
);

AND2x2_ASAP7_75t_L g434 ( 
.A(n_381),
.B(n_365),
.Y(n_434)
);

INVx1_ASAP7_75t_L g435 ( 
.A(n_407),
.Y(n_435)
);

OAI21xp5_ASAP7_75t_L g436 ( 
.A1(n_390),
.A2(n_354),
.B(n_348),
.Y(n_436)
);

AND2x2_ASAP7_75t_L g437 ( 
.A(n_381),
.B(n_365),
.Y(n_437)
);

INVx1_ASAP7_75t_L g438 ( 
.A(n_382),
.Y(n_438)
);

OAI21xp5_ASAP7_75t_SL g439 ( 
.A1(n_390),
.A2(n_341),
.B(n_330),
.Y(n_439)
);

INVx1_ASAP7_75t_L g440 ( 
.A(n_411),
.Y(n_440)
);

OAI22xp5_ASAP7_75t_L g441 ( 
.A1(n_422),
.A2(n_399),
.B1(n_392),
.B2(n_324),
.Y(n_441)
);

OAI22xp5_ASAP7_75t_L g442 ( 
.A1(n_423),
.A2(n_399),
.B1(n_392),
.B2(n_330),
.Y(n_442)
);

OAI222xp33_ASAP7_75t_L g443 ( 
.A1(n_412),
.A2(n_405),
.B1(n_395),
.B2(n_348),
.C1(n_388),
.C2(n_398),
.Y(n_443)
);

AOI21xp5_ASAP7_75t_L g444 ( 
.A1(n_421),
.A2(n_330),
.B(n_341),
.Y(n_444)
);

INVx1_ASAP7_75t_L g445 ( 
.A(n_416),
.Y(n_445)
);

INVx1_ASAP7_75t_L g446 ( 
.A(n_417),
.Y(n_446)
);

OAI21xp5_ASAP7_75t_L g447 ( 
.A1(n_436),
.A2(n_368),
.B(n_367),
.Y(n_447)
);

INVx1_ASAP7_75t_L g448 ( 
.A(n_419),
.Y(n_448)
);

AOI221xp5_ASAP7_75t_L g449 ( 
.A1(n_414),
.A2(n_413),
.B1(n_430),
.B2(n_432),
.C(n_435),
.Y(n_449)
);

AOI32xp33_ASAP7_75t_L g450 ( 
.A1(n_432),
.A2(n_405),
.A3(n_395),
.B1(n_388),
.B2(n_398),
.Y(n_450)
);

AOI22xp33_ASAP7_75t_L g451 ( 
.A1(n_427),
.A2(n_330),
.B1(n_433),
.B2(n_418),
.Y(n_451)
);

O2A1O1Ixp33_ASAP7_75t_L g452 ( 
.A1(n_418),
.A2(n_439),
.B(n_424),
.C(n_425),
.Y(n_452)
);

AOI22xp5_ASAP7_75t_L g453 ( 
.A1(n_438),
.A2(n_330),
.B1(n_304),
.B2(n_281),
.Y(n_453)
);

NOR3xp33_ASAP7_75t_L g454 ( 
.A(n_426),
.B(n_245),
.C(n_229),
.Y(n_454)
);

INVx1_ASAP7_75t_L g455 ( 
.A(n_420),
.Y(n_455)
);

AOI321xp33_ASAP7_75t_L g456 ( 
.A1(n_429),
.A2(n_370),
.A3(n_368),
.B1(n_367),
.B2(n_268),
.C(n_281),
.Y(n_456)
);

OAI221xp5_ASAP7_75t_L g457 ( 
.A1(n_429),
.A2(n_428),
.B1(n_420),
.B2(n_415),
.C(n_370),
.Y(n_457)
);

AO21x1_ASAP7_75t_L g458 ( 
.A1(n_431),
.A2(n_352),
.B(n_345),
.Y(n_458)
);

AOI322xp5_ASAP7_75t_L g459 ( 
.A1(n_437),
.A2(n_434),
.A3(n_431),
.B1(n_334),
.B2(n_357),
.C1(n_343),
.C2(n_319),
.Y(n_459)
);

NOR2xp33_ASAP7_75t_L g460 ( 
.A(n_431),
.B(n_397),
.Y(n_460)
);

OAI322xp33_ASAP7_75t_L g461 ( 
.A1(n_434),
.A2(n_357),
.A3(n_325),
.B1(n_347),
.B2(n_272),
.C1(n_271),
.C2(n_345),
.Y(n_461)
);

OAI221xp5_ASAP7_75t_L g462 ( 
.A1(n_437),
.A2(n_245),
.B1(n_325),
.B2(n_345),
.C(n_229),
.Y(n_462)
);

AOI22xp5_ASAP7_75t_L g463 ( 
.A1(n_422),
.A2(n_304),
.B1(n_281),
.B2(n_268),
.Y(n_463)
);

A2O1A1Ixp33_ASAP7_75t_L g464 ( 
.A1(n_452),
.A2(n_463),
.B(n_456),
.C(n_449),
.Y(n_464)
);

NAND2xp5_ASAP7_75t_L g465 ( 
.A(n_454),
.B(n_397),
.Y(n_465)
);

AOI211x1_ASAP7_75t_L g466 ( 
.A1(n_443),
.A2(n_334),
.B(n_343),
.C(n_337),
.Y(n_466)
);

AOI21xp5_ASAP7_75t_L g467 ( 
.A1(n_441),
.A2(n_304),
.B(n_239),
.Y(n_467)
);

OAI31xp33_ASAP7_75t_SL g468 ( 
.A1(n_442),
.A2(n_334),
.A3(n_343),
.B(n_232),
.Y(n_468)
);

INVx1_ASAP7_75t_L g469 ( 
.A(n_440),
.Y(n_469)
);

AOI221xp5_ASAP7_75t_L g470 ( 
.A1(n_457),
.A2(n_271),
.B1(n_272),
.B2(n_260),
.C(n_234),
.Y(n_470)
);

OAI211xp5_ASAP7_75t_SL g471 ( 
.A1(n_450),
.A2(n_234),
.B(n_235),
.C(n_325),
.Y(n_471)
);

OAI221xp5_ASAP7_75t_L g472 ( 
.A1(n_451),
.A2(n_270),
.B1(n_347),
.B2(n_265),
.C(n_321),
.Y(n_472)
);

NAND3xp33_ASAP7_75t_L g473 ( 
.A(n_454),
.B(n_347),
.C(n_265),
.Y(n_473)
);

AND2x2_ASAP7_75t_L g474 ( 
.A(n_460),
.B(n_337),
.Y(n_474)
);

A2O1A1O1Ixp25_ASAP7_75t_L g475 ( 
.A1(n_458),
.A2(n_444),
.B(n_462),
.C(n_447),
.D(n_446),
.Y(n_475)
);

OAI31xp33_ASAP7_75t_L g476 ( 
.A1(n_443),
.A2(n_337),
.A3(n_321),
.B(n_319),
.Y(n_476)
);

AOI21xp5_ASAP7_75t_L g477 ( 
.A1(n_461),
.A2(n_270),
.B(n_232),
.Y(n_477)
);

AOI21xp5_ASAP7_75t_L g478 ( 
.A1(n_453),
.A2(n_270),
.B(n_232),
.Y(n_478)
);

OAI211xp5_ASAP7_75t_SL g479 ( 
.A1(n_459),
.A2(n_238),
.B(n_265),
.C(n_309),
.Y(n_479)
);

OAI322xp33_ASAP7_75t_L g480 ( 
.A1(n_445),
.A2(n_344),
.A3(n_340),
.B1(n_331),
.B2(n_300),
.C1(n_303),
.C2(n_299),
.Y(n_480)
);

A2O1A1Ixp33_ASAP7_75t_SL g481 ( 
.A1(n_455),
.A2(n_265),
.B(n_319),
.C(n_321),
.Y(n_481)
);

A2O1A1Ixp33_ASAP7_75t_L g482 ( 
.A1(n_448),
.A2(n_243),
.B(n_319),
.C(n_321),
.Y(n_482)
);

NAND3xp33_ASAP7_75t_L g483 ( 
.A(n_454),
.B(n_265),
.C(n_260),
.Y(n_483)
);

NAND4xp25_ASAP7_75t_L g484 ( 
.A(n_449),
.B(n_238),
.C(n_299),
.D(n_303),
.Y(n_484)
);

AOI221xp5_ASAP7_75t_L g485 ( 
.A1(n_441),
.A2(n_319),
.B1(n_321),
.B2(n_309),
.C(n_303),
.Y(n_485)
);

NOR3xp33_ASAP7_75t_L g486 ( 
.A(n_464),
.B(n_277),
.C(n_278),
.Y(n_486)
);

NOR3xp33_ASAP7_75t_L g487 ( 
.A(n_484),
.B(n_277),
.C(n_278),
.Y(n_487)
);

AOI21xp5_ASAP7_75t_L g488 ( 
.A1(n_465),
.A2(n_263),
.B(n_240),
.Y(n_488)
);

NOR3xp33_ASAP7_75t_L g489 ( 
.A(n_475),
.B(n_277),
.C(n_223),
.Y(n_489)
);

NOR4xp25_ASAP7_75t_L g490 ( 
.A(n_479),
.B(n_266),
.C(n_262),
.D(n_259),
.Y(n_490)
);

AOI221xp5_ASAP7_75t_L g491 ( 
.A1(n_485),
.A2(n_309),
.B1(n_300),
.B2(n_328),
.C(n_331),
.Y(n_491)
);

O2A1O1Ixp33_ASAP7_75t_L g492 ( 
.A1(n_476),
.A2(n_242),
.B(n_300),
.C(n_263),
.Y(n_492)
);

NOR3xp33_ASAP7_75t_L g493 ( 
.A(n_473),
.B(n_277),
.C(n_223),
.Y(n_493)
);

INVx1_ASAP7_75t_L g494 ( 
.A(n_469),
.Y(n_494)
);

NAND4xp25_ASAP7_75t_L g495 ( 
.A(n_468),
.B(n_277),
.C(n_240),
.D(n_259),
.Y(n_495)
);

NAND2xp5_ASAP7_75t_L g496 ( 
.A(n_470),
.B(n_344),
.Y(n_496)
);

AOI22xp5_ASAP7_75t_L g497 ( 
.A1(n_479),
.A2(n_344),
.B1(n_340),
.B2(n_331),
.Y(n_497)
);

INVx1_ASAP7_75t_SL g498 ( 
.A(n_474),
.Y(n_498)
);

OAI22xp5_ASAP7_75t_L g499 ( 
.A1(n_466),
.A2(n_328),
.B1(n_340),
.B2(n_344),
.Y(n_499)
);

OR3x1_ASAP7_75t_L g500 ( 
.A(n_471),
.B(n_266),
.C(n_258),
.Y(n_500)
);

AND4x1_ASAP7_75t_L g501 ( 
.A(n_486),
.B(n_489),
.C(n_487),
.D(n_490),
.Y(n_501)
);

NOR2x1_ASAP7_75t_L g502 ( 
.A(n_494),
.B(n_483),
.Y(n_502)
);

NOR3xp33_ASAP7_75t_SL g503 ( 
.A(n_495),
.B(n_472),
.C(n_478),
.Y(n_503)
);

NAND2xp5_ASAP7_75t_L g504 ( 
.A(n_498),
.B(n_467),
.Y(n_504)
);

OR2x2_ASAP7_75t_L g505 ( 
.A(n_496),
.B(n_482),
.Y(n_505)
);

NOR3xp33_ASAP7_75t_L g506 ( 
.A(n_492),
.B(n_480),
.C(n_477),
.Y(n_506)
);

INVxp67_ASAP7_75t_L g507 ( 
.A(n_488),
.Y(n_507)
);

AOI211x1_ASAP7_75t_L g508 ( 
.A1(n_500),
.A2(n_481),
.B(n_290),
.C(n_258),
.Y(n_508)
);

OAI211xp5_ASAP7_75t_SL g509 ( 
.A1(n_491),
.A2(n_262),
.B(n_312),
.C(n_311),
.Y(n_509)
);

OR2x2_ASAP7_75t_L g510 ( 
.A(n_499),
.B(n_220),
.Y(n_510)
);

INVx1_ASAP7_75t_L g511 ( 
.A(n_497),
.Y(n_511)
);

NOR2x1_ASAP7_75t_L g512 ( 
.A(n_493),
.B(n_273),
.Y(n_512)
);

NAND3xp33_ASAP7_75t_L g513 ( 
.A(n_486),
.B(n_210),
.C(n_227),
.Y(n_513)
);

NOR4xp25_ASAP7_75t_L g514 ( 
.A(n_492),
.B(n_254),
.C(n_257),
.D(n_312),
.Y(n_514)
);

NOR4xp25_ASAP7_75t_L g515 ( 
.A(n_492),
.B(n_254),
.C(n_257),
.D(n_312),
.Y(n_515)
);

INVx1_ASAP7_75t_L g516 ( 
.A(n_504),
.Y(n_516)
);

INVx1_ASAP7_75t_L g517 ( 
.A(n_502),
.Y(n_517)
);

AND4x1_ASAP7_75t_L g518 ( 
.A(n_503),
.B(n_290),
.C(n_311),
.D(n_275),
.Y(n_518)
);

NOR4xp75_ASAP7_75t_SL g519 ( 
.A(n_501),
.B(n_220),
.C(n_263),
.D(n_273),
.Y(n_519)
);

NAND4xp75_ASAP7_75t_L g520 ( 
.A(n_512),
.B(n_218),
.C(n_290),
.D(n_340),
.Y(n_520)
);

AO22x1_ASAP7_75t_L g521 ( 
.A1(n_506),
.A2(n_273),
.B1(n_210),
.B2(n_227),
.Y(n_521)
);

AOI221xp5_ASAP7_75t_L g522 ( 
.A1(n_507),
.A2(n_273),
.B1(n_210),
.B2(n_290),
.C(n_227),
.Y(n_522)
);

NAND2xp5_ASAP7_75t_SL g523 ( 
.A(n_508),
.B(n_210),
.Y(n_523)
);

INVx1_ASAP7_75t_L g524 ( 
.A(n_511),
.Y(n_524)
);

INVx5_ASAP7_75t_L g525 ( 
.A(n_513),
.Y(n_525)
);

NAND5xp2_ASAP7_75t_L g526 ( 
.A(n_505),
.B(n_515),
.C(n_514),
.D(n_509),
.E(n_510),
.Y(n_526)
);

INVx2_ASAP7_75t_L g527 ( 
.A(n_502),
.Y(n_527)
);

NAND4xp25_ASAP7_75t_L g528 ( 
.A(n_506),
.B(n_311),
.C(n_275),
.D(n_315),
.Y(n_528)
);

BUFx3_ASAP7_75t_L g529 ( 
.A(n_517),
.Y(n_529)
);

AOI21xp5_ASAP7_75t_L g530 ( 
.A1(n_527),
.A2(n_263),
.B(n_222),
.Y(n_530)
);

AOI211x1_ASAP7_75t_L g531 ( 
.A1(n_518),
.A2(n_308),
.B(n_310),
.C(n_314),
.Y(n_531)
);

NOR2x1_ASAP7_75t_L g532 ( 
.A(n_524),
.B(n_210),
.Y(n_532)
);

INVx4_ASAP7_75t_L g533 ( 
.A(n_525),
.Y(n_533)
);

NOR4xp75_ASAP7_75t_L g534 ( 
.A(n_520),
.B(n_523),
.C(n_519),
.D(n_526),
.Y(n_534)
);

NAND5xp2_ASAP7_75t_L g535 ( 
.A(n_516),
.B(n_294),
.C(n_310),
.D(n_308),
.E(n_314),
.Y(n_535)
);

INVx2_ASAP7_75t_SL g536 ( 
.A(n_533),
.Y(n_536)
);

INVx5_ASAP7_75t_L g537 ( 
.A(n_529),
.Y(n_537)
);

BUFx2_ASAP7_75t_L g538 ( 
.A(n_532),
.Y(n_538)
);

NAND2xp5_ASAP7_75t_L g539 ( 
.A(n_531),
.B(n_521),
.Y(n_539)
);

NAND2xp33_ASAP7_75t_SL g540 ( 
.A(n_534),
.B(n_525),
.Y(n_540)
);

NAND2xp5_ASAP7_75t_L g541 ( 
.A(n_530),
.B(n_525),
.Y(n_541)
);

NOR2xp33_ASAP7_75t_SL g542 ( 
.A(n_537),
.B(n_528),
.Y(n_542)
);

NAND2xp5_ASAP7_75t_L g543 ( 
.A(n_537),
.B(n_522),
.Y(n_543)
);

OAI22xp5_ASAP7_75t_SL g544 ( 
.A1(n_536),
.A2(n_535),
.B1(n_273),
.B2(n_210),
.Y(n_544)
);

INVx2_ASAP7_75t_L g545 ( 
.A(n_538),
.Y(n_545)
);

OAI22xp5_ASAP7_75t_L g546 ( 
.A1(n_539),
.A2(n_273),
.B1(n_227),
.B2(n_306),
.Y(n_546)
);

HB1xp67_ASAP7_75t_L g547 ( 
.A(n_545),
.Y(n_547)
);

OA211x2_ASAP7_75t_L g548 ( 
.A1(n_542),
.A2(n_541),
.B(n_540),
.C(n_220),
.Y(n_548)
);

OAI22xp33_ASAP7_75t_L g549 ( 
.A1(n_547),
.A2(n_543),
.B1(n_546),
.B2(n_544),
.Y(n_549)
);

AOI221xp5_ASAP7_75t_L g550 ( 
.A1(n_548),
.A2(n_273),
.B1(n_237),
.B2(n_222),
.C(n_307),
.Y(n_550)
);

NAND2xp5_ASAP7_75t_L g551 ( 
.A(n_549),
.B(n_220),
.Y(n_551)
);

OR2x6_ASAP7_75t_L g552 ( 
.A(n_551),
.B(n_550),
.Y(n_552)
);

AOI211xp5_ASAP7_75t_L g553 ( 
.A1(n_552),
.A2(n_237),
.B(n_273),
.C(n_255),
.Y(n_553)
);


endmodule