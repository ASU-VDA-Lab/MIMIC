module fake_jpeg_28594_n_77 (n_13, n_21, n_1, n_10, n_6, n_22, n_14, n_19, n_18, n_20, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_77);

input n_13;
input n_21;
input n_1;
input n_10;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_77;

wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_73;
wire n_59;
wire n_65;
wire n_42;
wire n_49;
wire n_76;
wire n_28;
wire n_38;
wire n_26;
wire n_74;
wire n_31;
wire n_29;
wire n_50;
wire n_57;
wire n_23;
wire n_69;
wire n_27;
wire n_40;
wire n_71;
wire n_30;
wire n_24;
wire n_44;
wire n_25;
wire n_75;
wire n_37;
wire n_70;
wire n_66;
wire n_61;
wire n_45;
wire n_68;
wire n_52;
wire n_58;
wire n_41;
wire n_60;
wire n_63;
wire n_34;
wire n_39;
wire n_72;
wire n_56;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_35;
wire n_48;
wire n_46;
wire n_36;
wire n_62;
wire n_43;
wire n_32;

BUFx12f_ASAP7_75t_L g23 ( 
.A(n_18),
.Y(n_23)
);

INVx2_ASAP7_75t_L g24 ( 
.A(n_12),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_3),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_3),
.Y(n_26)
);

BUFx16f_ASAP7_75t_L g27 ( 
.A(n_2),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_22),
.Y(n_28)
);

BUFx12f_ASAP7_75t_L g29 ( 
.A(n_16),
.Y(n_29)
);

BUFx8_ASAP7_75t_L g30 ( 
.A(n_13),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_21),
.Y(n_31)
);

BUFx10_ASAP7_75t_L g32 ( 
.A(n_6),
.Y(n_32)
);

INVx4_ASAP7_75t_L g33 ( 
.A(n_27),
.Y(n_33)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_33),
.Y(n_43)
);

BUFx2_ASAP7_75t_SL g34 ( 
.A(n_32),
.Y(n_34)
);

BUFx4f_ASAP7_75t_SL g48 ( 
.A(n_34),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_25),
.Y(n_35)
);

NAND2xp5_ASAP7_75t_L g42 ( 
.A(n_35),
.B(n_39),
.Y(n_42)
);

BUFx12f_ASAP7_75t_L g36 ( 
.A(n_30),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g41 ( 
.A(n_36),
.B(n_37),
.Y(n_41)
);

CKINVDCx14_ASAP7_75t_R g37 ( 
.A(n_24),
.Y(n_37)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_26),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_L g44 ( 
.A(n_38),
.B(n_28),
.Y(n_44)
);

INVx2_ASAP7_75t_L g39 ( 
.A(n_24),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g40 ( 
.A(n_23),
.B(n_0),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_44),
.B(n_47),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_L g45 ( 
.A(n_40),
.B(n_32),
.Y(n_45)
);

NAND2xp5_ASAP7_75t_L g56 ( 
.A(n_45),
.B(n_46),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_L g46 ( 
.A(n_36),
.B(n_31),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_L g47 ( 
.A(n_34),
.B(n_0),
.Y(n_47)
);

OAI22xp5_ASAP7_75t_L g49 ( 
.A1(n_35),
.A2(n_29),
.B1(n_23),
.B2(n_11),
.Y(n_49)
);

AOI22xp33_ASAP7_75t_L g51 ( 
.A1(n_49),
.A2(n_1),
.B1(n_2),
.B2(n_4),
.Y(n_51)
);

NOR2x1_ASAP7_75t_R g50 ( 
.A(n_41),
.B(n_29),
.Y(n_50)
);

AND2x2_ASAP7_75t_L g66 ( 
.A(n_50),
.B(n_55),
.Y(n_66)
);

OAI22xp5_ASAP7_75t_SL g63 ( 
.A1(n_51),
.A2(n_57),
.B1(n_9),
.B2(n_14),
.Y(n_63)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_43),
.Y(n_52)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_52),
.Y(n_64)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_42),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_53),
.B(n_60),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_SL g54 ( 
.A(n_49),
.B(n_10),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_L g61 ( 
.A(n_54),
.B(n_58),
.Y(n_61)
);

AND2x2_ASAP7_75t_L g55 ( 
.A(n_48),
.B(n_4),
.Y(n_55)
);

AOI22xp33_ASAP7_75t_L g57 ( 
.A1(n_48),
.A2(n_20),
.B1(n_7),
.B2(n_8),
.Y(n_57)
);

AND2x2_ASAP7_75t_L g58 ( 
.A(n_45),
.B(n_5),
.Y(n_58)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_43),
.Y(n_60)
);

CKINVDCx20_ASAP7_75t_R g62 ( 
.A(n_55),
.Y(n_62)
);

AOI21xp5_ASAP7_75t_L g68 ( 
.A1(n_62),
.A2(n_66),
.B(n_59),
.Y(n_68)
);

XOR2xp5_ASAP7_75t_L g69 ( 
.A(n_63),
.B(n_54),
.Y(n_69)
);

XOR2x2_ASAP7_75t_L g67 ( 
.A(n_66),
.B(n_56),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_SL g71 ( 
.A(n_67),
.B(n_68),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_L g70 ( 
.A(n_69),
.B(n_59),
.Y(n_70)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_70),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_SL g73 ( 
.A(n_72),
.B(n_65),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_L g74 ( 
.A(n_73),
.B(n_65),
.Y(n_74)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_74),
.Y(n_75)
);

AOI322xp5_ASAP7_75t_L g76 ( 
.A1(n_75),
.A2(n_71),
.A3(n_61),
.B1(n_58),
.B2(n_64),
.C1(n_17),
.C2(n_19),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_L g77 ( 
.A(n_76),
.B(n_15),
.Y(n_77)
);


endmodule