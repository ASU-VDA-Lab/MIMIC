module fake_jpeg_8062_n_136 (n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_136);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_136;

wire n_117;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_73;
wire n_14;
wire n_19;
wire n_84;
wire n_59;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_31;
wire n_29;
wire n_103;
wire n_50;
wire n_15;
wire n_124;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_30;
wire n_106;
wire n_111;
wire n_44;
wire n_24;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_20;
wire n_18;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_22;
wire n_101;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_97;
wire n_135;
wire n_36;
wire n_62;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_96;

INVx1_ASAP7_75t_L g13 ( 
.A(n_6),
.Y(n_13)
);

INVxp67_ASAP7_75t_L g14 ( 
.A(n_11),
.Y(n_14)
);

INVx1_ASAP7_75t_L g15 ( 
.A(n_1),
.Y(n_15)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_6),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_4),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_4),
.Y(n_18)
);

INVx2_ASAP7_75t_L g19 ( 
.A(n_4),
.Y(n_19)
);

INVx8_ASAP7_75t_L g20 ( 
.A(n_3),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_8),
.Y(n_21)
);

BUFx4f_ASAP7_75t_SL g22 ( 
.A(n_3),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_5),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_9),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_5),
.Y(n_25)
);

INVx3_ASAP7_75t_L g26 ( 
.A(n_11),
.Y(n_26)
);

INVx2_ASAP7_75t_L g27 ( 
.A(n_22),
.Y(n_27)
);

NOR2xp33_ASAP7_75t_L g46 ( 
.A(n_27),
.B(n_28),
.Y(n_46)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_22),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_22),
.Y(n_29)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_29),
.Y(n_37)
);

INVx2_ASAP7_75t_L g30 ( 
.A(n_19),
.Y(n_30)
);

INVx6_ASAP7_75t_L g48 ( 
.A(n_30),
.Y(n_48)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_19),
.Y(n_31)
);

NAND2xp5_ASAP7_75t_SL g42 ( 
.A(n_31),
.B(n_34),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_20),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_32),
.Y(n_40)
);

INVx2_ASAP7_75t_L g33 ( 
.A(n_20),
.Y(n_33)
);

INVx2_ASAP7_75t_L g39 ( 
.A(n_33),
.Y(n_39)
);

INVx4_ASAP7_75t_L g34 ( 
.A(n_26),
.Y(n_34)
);

INVx2_ASAP7_75t_L g35 ( 
.A(n_26),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_35),
.Y(n_43)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_27),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g51 ( 
.A(n_36),
.B(n_38),
.Y(n_51)
);

AOI22xp33_ASAP7_75t_L g38 ( 
.A1(n_34),
.A2(n_25),
.B1(n_13),
.B2(n_15),
.Y(n_38)
);

AND2x2_ASAP7_75t_L g41 ( 
.A(n_35),
.B(n_25),
.Y(n_41)
);

NAND2xp5_ASAP7_75t_L g50 ( 
.A(n_41),
.B(n_44),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_L g44 ( 
.A(n_30),
.B(n_17),
.Y(n_44)
);

NAND2xp5_ASAP7_75t_L g45 ( 
.A(n_33),
.B(n_17),
.Y(n_45)
);

NAND2xp5_ASAP7_75t_L g61 ( 
.A(n_45),
.B(n_16),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_SL g47 ( 
.A(n_32),
.B(n_18),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_47),
.B(n_18),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_32),
.Y(n_49)
);

INVx3_ASAP7_75t_L g59 ( 
.A(n_49),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_SL g68 ( 
.A(n_52),
.B(n_21),
.Y(n_68)
);

INVxp67_ASAP7_75t_L g53 ( 
.A(n_46),
.Y(n_53)
);

INVxp67_ASAP7_75t_L g66 ( 
.A(n_53),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_40),
.Y(n_54)
);

INVx3_ASAP7_75t_L g72 ( 
.A(n_54),
.Y(n_72)
);

INVx4_ASAP7_75t_L g55 ( 
.A(n_43),
.Y(n_55)
);

INVx2_ASAP7_75t_SL g75 ( 
.A(n_55),
.Y(n_75)
);

CKINVDCx16_ASAP7_75t_R g56 ( 
.A(n_45),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_56),
.B(n_58),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g57 ( 
.A(n_36),
.B(n_47),
.Y(n_57)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_57),
.Y(n_64)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_44),
.Y(n_58)
);

MAJIxp5_ASAP7_75t_L g60 ( 
.A(n_37),
.B(n_23),
.C(n_24),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_L g67 ( 
.A(n_60),
.B(n_61),
.Y(n_67)
);

BUFx24_ASAP7_75t_L g62 ( 
.A(n_43),
.Y(n_62)
);

INVxp67_ASAP7_75t_L g71 ( 
.A(n_62),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_60),
.B(n_42),
.Y(n_65)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_65),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_SL g82 ( 
.A(n_68),
.B(n_53),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_L g69 ( 
.A(n_56),
.B(n_41),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_L g78 ( 
.A(n_69),
.B(n_70),
.Y(n_78)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_61),
.Y(n_70)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_51),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_L g80 ( 
.A(n_73),
.B(n_74),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_L g74 ( 
.A(n_58),
.B(n_41),
.Y(n_74)
);

INVx2_ASAP7_75t_L g76 ( 
.A(n_62),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_76),
.B(n_55),
.Y(n_79)
);

XNOR2xp5_ASAP7_75t_SL g77 ( 
.A(n_74),
.B(n_50),
.Y(n_77)
);

XNOR2xp5_ASAP7_75t_L g92 ( 
.A(n_77),
.B(n_81),
.Y(n_92)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_79),
.Y(n_91)
);

MAJIxp5_ASAP7_75t_L g81 ( 
.A(n_69),
.B(n_50),
.C(n_37),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_SL g97 ( 
.A(n_82),
.B(n_86),
.Y(n_97)
);

OAI21xp5_ASAP7_75t_L g83 ( 
.A1(n_63),
.A2(n_13),
.B(n_16),
.Y(n_83)
);

XNOR2xp5_ASAP7_75t_L g95 ( 
.A(n_83),
.B(n_84),
.Y(n_95)
);

MAJIxp5_ASAP7_75t_L g84 ( 
.A(n_70),
.B(n_39),
.C(n_48),
.Y(n_84)
);

AOI22xp5_ASAP7_75t_L g85 ( 
.A1(n_73),
.A2(n_48),
.B1(n_39),
.B2(n_59),
.Y(n_85)
);

OAI22xp5_ASAP7_75t_L g90 ( 
.A1(n_85),
.A2(n_89),
.B1(n_75),
.B2(n_72),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_L g86 ( 
.A(n_64),
.B(n_15),
.Y(n_86)
);

MAJIxp5_ASAP7_75t_L g88 ( 
.A(n_67),
.B(n_43),
.C(n_62),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_L g94 ( 
.A(n_88),
.B(n_67),
.Y(n_94)
);

AOI22xp33_ASAP7_75t_L g89 ( 
.A1(n_75),
.A2(n_59),
.B1(n_49),
.B2(n_40),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_SL g110 ( 
.A(n_90),
.B(n_93),
.Y(n_110)
);

CKINVDCx20_ASAP7_75t_R g93 ( 
.A(n_85),
.Y(n_93)
);

MAJIxp5_ASAP7_75t_L g101 ( 
.A(n_94),
.B(n_88),
.C(n_81),
.Y(n_101)
);

AOI22xp5_ASAP7_75t_L g96 ( 
.A1(n_77),
.A2(n_66),
.B1(n_72),
.B2(n_71),
.Y(n_96)
);

OAI22xp5_ASAP7_75t_SL g106 ( 
.A1(n_96),
.A2(n_78),
.B1(n_71),
.B2(n_14),
.Y(n_106)
);

NAND3xp33_ASAP7_75t_L g98 ( 
.A(n_80),
.B(n_66),
.C(n_10),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g105 ( 
.A(n_98),
.B(n_100),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_84),
.B(n_75),
.Y(n_99)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_99),
.Y(n_102)
);

CKINVDCx20_ASAP7_75t_R g100 ( 
.A(n_83),
.Y(n_100)
);

MAJIxp5_ASAP7_75t_L g114 ( 
.A(n_101),
.B(n_103),
.C(n_107),
.Y(n_114)
);

XOR2xp5_ASAP7_75t_L g103 ( 
.A(n_92),
.B(n_94),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_91),
.B(n_87),
.Y(n_104)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_104),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_106),
.B(n_95),
.Y(n_111)
);

XOR2xp5_ASAP7_75t_L g107 ( 
.A(n_92),
.B(n_96),
.Y(n_107)
);

XNOR2xp5_ASAP7_75t_L g108 ( 
.A(n_95),
.B(n_14),
.Y(n_108)
);

XOR2xp5_ASAP7_75t_L g118 ( 
.A(n_108),
.B(n_7),
.Y(n_118)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_97),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_L g115 ( 
.A(n_109),
.B(n_54),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_L g119 ( 
.A(n_111),
.B(n_118),
.Y(n_119)
);

XNOR2xp5_ASAP7_75t_SL g112 ( 
.A(n_107),
.B(n_8),
.Y(n_112)
);

XOR2xp5_ASAP7_75t_L g121 ( 
.A(n_112),
.B(n_118),
.Y(n_121)
);

OAI322xp33_ASAP7_75t_L g113 ( 
.A1(n_102),
.A2(n_7),
.A3(n_12),
.B1(n_10),
.B2(n_9),
.C1(n_5),
.C2(n_6),
.Y(n_113)
);

AOI21xp33_ASAP7_75t_L g124 ( 
.A1(n_113),
.A2(n_105),
.B(n_12),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_L g123 ( 
.A(n_115),
.B(n_116),
.Y(n_123)
);

OAI22xp5_ASAP7_75t_L g116 ( 
.A1(n_110),
.A2(n_76),
.B1(n_54),
.B2(n_62),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_L g126 ( 
.A(n_119),
.B(n_120),
.Y(n_126)
);

CKINVDCx20_ASAP7_75t_R g120 ( 
.A(n_117),
.Y(n_120)
);

XNOR2xp5_ASAP7_75t_L g122 ( 
.A(n_114),
.B(n_103),
.Y(n_122)
);

MAJIxp5_ASAP7_75t_L g128 ( 
.A(n_122),
.B(n_114),
.C(n_108),
.Y(n_128)
);

AOI22xp5_ASAP7_75t_SL g125 ( 
.A1(n_124),
.A2(n_112),
.B1(n_1),
.B2(n_2),
.Y(n_125)
);

NOR3xp33_ASAP7_75t_L g130 ( 
.A(n_125),
.B(n_129),
.C(n_0),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_L g127 ( 
.A(n_123),
.B(n_101),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_L g131 ( 
.A(n_127),
.B(n_128),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_L g129 ( 
.A(n_121),
.B(n_0),
.Y(n_129)
);

INVxp67_ASAP7_75t_L g133 ( 
.A(n_130),
.Y(n_133)
);

AOI322xp5_ASAP7_75t_L g132 ( 
.A1(n_126),
.A2(n_121),
.A3(n_122),
.B1(n_2),
.B2(n_3),
.C1(n_0),
.C2(n_1),
.Y(n_132)
);

INVxp67_ASAP7_75t_L g134 ( 
.A(n_132),
.Y(n_134)
);

AOI21x1_ASAP7_75t_L g135 ( 
.A1(n_134),
.A2(n_131),
.B(n_128),
.Y(n_135)
);

XNOR2xp5_ASAP7_75t_L g136 ( 
.A(n_135),
.B(n_133),
.Y(n_136)
);


endmodule