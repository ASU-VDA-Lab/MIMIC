module fake_jpeg_7454_n_47 (n_13, n_1, n_10, n_6, n_14, n_19, n_18, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_47);

input n_13;
input n_1;
input n_10;
input n_6;
input n_14;
input n_19;
input n_18;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_47;

wire n_21;
wire n_33;
wire n_45;
wire n_23;
wire n_27;
wire n_22;
wire n_40;
wire n_20;
wire n_35;
wire n_46;
wire n_41;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_24;
wire n_28;
wire n_38;
wire n_26;
wire n_44;
wire n_36;
wire n_25;
wire n_31;
wire n_29;
wire n_37;
wire n_43;
wire n_32;

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_6),
.Y(n_20)
);

INVx3_ASAP7_75t_L g21 ( 
.A(n_0),
.Y(n_21)
);

INVx2_ASAP7_75t_L g22 ( 
.A(n_17),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_7),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_2),
.Y(n_24)
);

NOR2xp33_ASAP7_75t_L g25 ( 
.A(n_1),
.B(n_10),
.Y(n_25)
);

INVx3_ASAP7_75t_L g26 ( 
.A(n_24),
.Y(n_26)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_26),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_22),
.Y(n_27)
);

NAND2xp5_ASAP7_75t_L g32 ( 
.A(n_27),
.B(n_28),
.Y(n_32)
);

NOR2xp33_ASAP7_75t_SL g28 ( 
.A(n_25),
.B(n_0),
.Y(n_28)
);

NAND2xp5_ASAP7_75t_SL g29 ( 
.A(n_24),
.B(n_1),
.Y(n_29)
);

CKINVDCx16_ASAP7_75t_R g33 ( 
.A(n_29),
.Y(n_33)
);

INVx2_ASAP7_75t_L g30 ( 
.A(n_22),
.Y(n_30)
);

INVx13_ASAP7_75t_L g39 ( 
.A(n_30),
.Y(n_39)
);

INVx5_ASAP7_75t_L g31 ( 
.A(n_21),
.Y(n_31)
);

AOI22xp5_ASAP7_75t_SL g34 ( 
.A1(n_31),
.A2(n_21),
.B1(n_20),
.B2(n_23),
.Y(n_34)
);

OAI21xp5_ASAP7_75t_L g42 ( 
.A1(n_34),
.A2(n_31),
.B(n_4),
.Y(n_42)
);

AOI22xp5_ASAP7_75t_L g35 ( 
.A1(n_30),
.A2(n_12),
.B1(n_18),
.B2(n_16),
.Y(n_35)
);

MAJIxp5_ASAP7_75t_L g40 ( 
.A(n_35),
.B(n_36),
.C(n_38),
.Y(n_40)
);

AOI22xp5_ASAP7_75t_L g36 ( 
.A1(n_26),
.A2(n_2),
.B1(n_3),
.B2(n_4),
.Y(n_36)
);

MAJIxp5_ASAP7_75t_L g38 ( 
.A(n_27),
.B(n_11),
.C(n_15),
.Y(n_38)
);

CKINVDCx16_ASAP7_75t_R g41 ( 
.A(n_37),
.Y(n_41)
);

NAND2xp5_ASAP7_75t_SL g44 ( 
.A(n_41),
.B(n_42),
.Y(n_44)
);

AOI22xp5_ASAP7_75t_L g43 ( 
.A1(n_40),
.A2(n_33),
.B1(n_39),
.B2(n_35),
.Y(n_43)
);

AOI322xp5_ASAP7_75t_L g45 ( 
.A1(n_43),
.A2(n_44),
.A3(n_34),
.B1(n_39),
.B2(n_32),
.C1(n_38),
.C2(n_14),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_45),
.Y(n_46)
);

AOI322xp5_ASAP7_75t_L g47 ( 
.A1(n_46),
.A2(n_5),
.A3(n_8),
.B1(n_9),
.B2(n_13),
.C1(n_19),
.C2(n_3),
.Y(n_47)
);


endmodule