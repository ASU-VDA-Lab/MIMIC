module real_aes_17439_n_249 (n_17, n_28, n_226, n_76, n_202, n_149, n_56, n_113, n_34, n_98, n_121, n_120, n_125, n_187, n_190, n_90, n_216, n_82, n_238, n_65, n_47, n_74, n_106, n_58, n_185, n_134, n_32, n_30, n_230, n_165, n_51, n_195, n_246, n_248, n_176, n_27, n_163, n_222, n_61, n_29, n_20, n_52, n_221, n_174, n_156, n_57, n_64, n_66, n_18, n_207, n_104, n_21, n_31, n_8, n_183, n_205, n_220, n_211, n_10, n_177, n_83, n_181, n_197, n_124, n_22, n_173, n_191, n_209, n_3, n_41, n_140, n_234, n_153, n_75, n_178, n_219, n_19, n_71, n_180, n_40, n_49, n_212, n_210, n_239, n_126, n_91, n_100, n_43, n_103, n_166, n_200, n_224, n_151, n_115, n_96, n_110, n_130, n_54, n_112, n_35, n_42, n_147, n_150, n_99, n_15, n_9, n_23, n_72, n_132, n_119, n_160, n_95, n_131, n_144, n_164, n_231, n_169, n_242, n_44, n_102, n_188, n_152, n_198, n_201, n_122, n_7, n_228, n_196, n_141, n_128, n_172, n_111, n_158, n_4, n_232, n_167, n_123, n_80, n_179, n_6, n_12, n_68, n_129, n_162, n_79, n_193, n_214, n_69, n_46, n_109, n_59, n_25, n_203, n_236, n_73, n_77, n_218, n_81, n_133, n_48, n_204, n_37, n_117, n_208, n_97, n_215, n_135, n_186, n_70, n_138, n_50, n_114, n_89, n_170, n_26, n_235, n_86, n_93, n_182, n_154, n_127, n_199, n_245, n_161, n_189, n_13, n_24, n_217, n_2, n_142, n_55, n_168, n_175, n_241, n_145, n_62, n_105, n_223, n_84, n_227, n_67, n_92, n_33, n_206, n_148, n_88, n_14, n_159, n_11, n_85, n_108, n_194, n_137, n_225, n_16, n_116, n_94, n_229, n_39, n_5, n_45, n_60, n_233, n_240, n_247, n_38, n_155, n_243, n_118, n_143, n_139, n_244, n_192, n_213, n_136, n_87, n_171, n_0, n_157, n_78, n_101, n_63, n_1, n_146, n_237, n_107, n_184, n_53, n_36, n_249);
input n_17;
input n_28;
input n_226;
input n_76;
input n_202;
input n_149;
input n_56;
input n_113;
input n_34;
input n_98;
input n_121;
input n_120;
input n_125;
input n_187;
input n_190;
input n_90;
input n_216;
input n_82;
input n_238;
input n_65;
input n_47;
input n_74;
input n_106;
input n_58;
input n_185;
input n_134;
input n_32;
input n_30;
input n_230;
input n_165;
input n_51;
input n_195;
input n_246;
input n_248;
input n_176;
input n_27;
input n_163;
input n_222;
input n_61;
input n_29;
input n_20;
input n_52;
input n_221;
input n_174;
input n_156;
input n_57;
input n_64;
input n_66;
input n_18;
input n_207;
input n_104;
input n_21;
input n_31;
input n_8;
input n_183;
input n_205;
input n_220;
input n_211;
input n_10;
input n_177;
input n_83;
input n_181;
input n_197;
input n_124;
input n_22;
input n_173;
input n_191;
input n_209;
input n_3;
input n_41;
input n_140;
input n_234;
input n_153;
input n_75;
input n_178;
input n_219;
input n_19;
input n_71;
input n_180;
input n_40;
input n_49;
input n_212;
input n_210;
input n_239;
input n_126;
input n_91;
input n_100;
input n_43;
input n_103;
input n_166;
input n_200;
input n_224;
input n_151;
input n_115;
input n_96;
input n_110;
input n_130;
input n_54;
input n_112;
input n_35;
input n_42;
input n_147;
input n_150;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_132;
input n_119;
input n_160;
input n_95;
input n_131;
input n_144;
input n_164;
input n_231;
input n_169;
input n_242;
input n_44;
input n_102;
input n_188;
input n_152;
input n_198;
input n_201;
input n_122;
input n_7;
input n_228;
input n_196;
input n_141;
input n_128;
input n_172;
input n_111;
input n_158;
input n_4;
input n_232;
input n_167;
input n_123;
input n_80;
input n_179;
input n_6;
input n_12;
input n_68;
input n_129;
input n_162;
input n_79;
input n_193;
input n_214;
input n_69;
input n_46;
input n_109;
input n_59;
input n_25;
input n_203;
input n_236;
input n_73;
input n_77;
input n_218;
input n_81;
input n_133;
input n_48;
input n_204;
input n_37;
input n_117;
input n_208;
input n_97;
input n_215;
input n_135;
input n_186;
input n_70;
input n_138;
input n_50;
input n_114;
input n_89;
input n_170;
input n_26;
input n_235;
input n_86;
input n_93;
input n_182;
input n_154;
input n_127;
input n_199;
input n_245;
input n_161;
input n_189;
input n_13;
input n_24;
input n_217;
input n_2;
input n_142;
input n_55;
input n_168;
input n_175;
input n_241;
input n_145;
input n_62;
input n_105;
input n_223;
input n_84;
input n_227;
input n_67;
input n_92;
input n_33;
input n_206;
input n_148;
input n_88;
input n_14;
input n_159;
input n_11;
input n_85;
input n_108;
input n_194;
input n_137;
input n_225;
input n_16;
input n_116;
input n_94;
input n_229;
input n_39;
input n_5;
input n_45;
input n_60;
input n_233;
input n_240;
input n_247;
input n_38;
input n_155;
input n_243;
input n_118;
input n_143;
input n_139;
input n_244;
input n_192;
input n_213;
input n_136;
input n_87;
input n_171;
input n_0;
input n_157;
input n_78;
input n_101;
input n_63;
input n_1;
input n_146;
input n_237;
input n_107;
input n_184;
input n_53;
input n_36;
output n_249;
wire n_476;
wire n_599;
wire n_887;
wire n_1279;
wire n_1314;
wire n_830;
wire n_1371;
wire n_624;
wire n_618;
wire n_933;
wire n_485;
wire n_822;
wire n_750;
wire n_503;
wire n_254;
wire n_469;
wire n_1310;
wire n_1376;
wire n_592;
wire n_761;
wire n_421;
wire n_329;
wire n_919;
wire n_1217;
wire n_571;
wire n_549;
wire n_1034;
wire n_1328;
wire n_1219;
wire n_952;
wire n_1166;
wire n_752;
wire n_448;
wire n_556;
wire n_341;
wire n_593;
wire n_989;
wire n_431;
wire n_1044;
wire n_963;
wire n_551;
wire n_884;
wire n_260;
wire n_814;
wire n_944;
wire n_1283;
wire n_983;
wire n_955;
wire n_975;
wire n_941;
wire n_1313;
wire n_870;
wire n_1248;
wire n_271;
wire n_548;
wire n_572;
wire n_815;
wire n_1140;
wire n_330;
wire n_786;
wire n_512;
wire n_395;
wire n_795;
wire n_292;
wire n_1379;
wire n_400;
wire n_1160;
wire n_1287;
wire n_883;
wire n_478;
wire n_553;
wire n_744;
wire n_1367;
wire n_1325;
wire n_1225;
wire n_875;
wire n_951;
wire n_1199;
wire n_791;
wire n_976;
wire n_636;
wire n_906;
wire n_477;
wire n_595;
wire n_343;
wire n_1282;
wire n_683;
wire n_840;
wire n_570;
wire n_675;
wire n_835;
wire n_732;
wire n_784;
wire n_281;
wire n_962;
wire n_755;
wire n_409;
wire n_781;
wire n_576;
wire n_956;
wire n_1242;
wire n_796;
wire n_874;
wire n_1126;
wire n_383;
wire n_455;
wire n_682;
wire n_812;
wire n_782;
wire n_817;
wire n_760;
wire n_608;
wire n_534;
wire n_708;
wire n_1020;
wire n_885;
wire n_950;
wire n_381;
wire n_1196;
wire n_1013;
wire n_808;
wire n_1224;
wire n_688;
wire n_1042;
wire n_363;
wire n_1317;
wire n_417;
wire n_323;
wire n_690;
wire n_499;
wire n_1142;
wire n_947;
wire n_970;
wire n_1149;
wire n_368;
wire n_527;
wire n_1342;
wire n_1346;
wire n_552;
wire n_590;
wire n_1293;
wire n_432;
wire n_1131;
wire n_1008;
wire n_805;
wire n_619;
wire n_1284;
wire n_1095;
wire n_1250;
wire n_360;
wire n_859;
wire n_1304;
wire n_685;
wire n_1080;
wire n_917;
wire n_1247;
wire n_501;
wire n_488;
wire n_1380;
wire n_954;
wire n_702;
wire n_1007;
wire n_351;
wire n_898;
wire n_562;
wire n_1022;
wire n_1073;
wire n_404;
wire n_728;
wire n_1301;
wire n_1201;
wire n_997;
wire n_1105;
wire n_1243;
wire n_306;
wire n_1003;
wire n_346;
wire n_293;
wire n_749;
wire n_914;
wire n_1286;
wire n_494;
wire n_927;
wire n_723;
wire n_972;
wire n_1351;
wire n_1209;
wire n_411;
wire n_498;
wire n_765;
wire n_648;
wire n_939;
wire n_290;
wire n_928;
wire n_789;
wire n_738;
wire n_922;
wire n_1048;
wire n_787;
wire n_1214;
wire n_806;
wire n_715;
wire n_420;
wire n_1258;
wire n_873;
wire n_438;
wire n_446;
wire n_1281;
wire n_712;
wire n_266;
wire n_422;
wire n_861;
wire n_479;
wire n_825;
wire n_541;
wire n_839;
wire n_811;
wire n_558;
wire n_724;
wire n_440;
wire n_1231;
wire n_1305;
wire n_315;
wire n_1161;
wire n_686;
wire n_1299;
wire n_949;
wire n_586;
wire n_788;
wire n_441;
wire n_1045;
wire n_1339;
wire n_837;
wire n_1349;
wire n_829;
wire n_1030;
wire n_1348;
wire n_375;
wire n_597;
wire n_1036;
wire n_687;
wire n_258;
wire n_652;
wire n_500;
wire n_804;
wire n_1173;
wire n_854;
wire n_424;
wire n_877;
wire n_802;
wire n_337;
wire n_264;
wire n_480;
wire n_684;
wire n_1178;
wire n_821;
wire n_1018;
wire n_980;
wire n_1233;
wire n_1106;
wire n_1205;
wire n_838;
wire n_635;
wire n_792;
wire n_665;
wire n_991;
wire n_667;
wire n_580;
wire n_1004;
wire n_1370;
wire n_979;
wire n_445;
wire n_596;
wire n_1197;
wire n_657;
wire n_328;
wire n_1260;
wire n_355;
wire n_1129;
wire n_1285;
wire n_742;
wire n_1014;
wire n_461;
wire n_1047;
wire n_1016;
wire n_694;
wire n_1350;
wire n_894;
wire n_545;
wire n_401;
wire n_538;
wire n_537;
wire n_560;
wire n_1094;
wire n_1220;
wire n_696;
wire n_1147;
wire n_704;
wire n_453;
wire n_647;
wire n_399;
wire n_948;
wire n_700;
wire n_677;
wire n_1269;
wire n_378;
wire n_591;
wire n_1366;
wire n_678;
wire n_415;
wire n_564;
wire n_638;
wire n_510;
wire n_1361;
wire n_1358;
wire n_550;
wire n_966;
wire n_333;
wire n_1368;
wire n_994;
wire n_384;
wire n_1128;
wire n_1098;
wire n_824;
wire n_1238;
wire n_992;
wire n_813;
wire n_1338;
wire n_981;
wire n_1182;
wire n_872;
wire n_1086;
wire n_1070;
wire n_1189;
wire n_535;
wire n_882;
wire n_1210;
wire n_746;
wire n_656;
wire n_1148;
wire n_860;
wire n_748;
wire n_1261;
wire n_1062;
wire n_651;
wire n_801;
wire n_1271;
wire n_529;
wire n_504;
wire n_973;
wire n_1364;
wire n_659;
wire n_634;
wire n_903;
wire n_565;
wire n_925;
wire n_457;
wire n_1121;
wire n_1059;
wire n_493;
wire n_311;
wire n_278;
wire n_1362;
wire n_610;
wire n_1035;
wire n_620;
wire n_722;
wire n_1174;
wire n_1193;
wire n_277;
wire n_754;
wire n_508;
wire n_1141;
wire n_1112;
wire n_428;
wire n_783;
wire n_1107;
wire n_505;
wire n_600;
wire n_731;
wire n_964;
wire n_605;
wire n_406;
wire n_617;
wire n_602;
wire n_402;
wire n_733;
wire n_658;
wire n_676;
wire n_531;
wire n_1031;
wire n_807;
wire n_255;
wire n_286;
wire n_1011;
wire n_416;
wire n_895;
wire n_799;
wire n_490;
wire n_261;
wire n_391;
wire n_695;
wire n_1181;
wire n_881;
wire n_645;
wire n_1145;
wire n_557;
wire n_985;
wire n_777;
wire n_910;
wire n_642;
wire n_613;
wire n_1125;
wire n_296;
wire n_1347;
wire n_1163;
wire n_1278;
wire n_734;
wire n_735;
wire n_334;
wire n_1179;
wire n_569;
wire n_1171;
wire n_785;
wire n_1203;
wire n_1232;
wire n_471;
wire n_853;
wire n_810;
wire n_1136;
wire n_699;
wire n_1187;
wire n_1000;
wire n_649;
wire n_358;
wire n_1234;
wire n_622;
wire n_1002;
wire n_1353;
wire n_1165;
wire n_1058;
wire n_1216;
wire n_662;
wire n_850;
wire n_265;
wire n_354;
wire n_720;
wire n_1026;
wire n_492;
wire n_407;
wire n_1023;
wire n_419;
wire n_730;
wire n_643;
wire n_486;
wire n_291;
wire n_779;
wire n_481;
wire n_691;
wire n_589;
wire n_365;
wire n_526;
wire n_268;
wire n_1194;
wire n_282;
wire n_389;
wire n_701;
wire n_809;
wire n_679;
wire n_520;
wire n_926;
wire n_942;
wire n_1374;
wire n_1120;
wire n_689;
wire n_946;
wire n_300;
wire n_753;
wire n_1188;
wire n_623;
wire n_1032;
wire n_721;
wire n_1133;
wire n_313;
wire n_739;
wire n_1322;
wire n_1162;
wire n_762;
wire n_325;
wire n_1298;
wire n_442;
wire n_740;
wire n_1357;
wire n_639;
wire n_1186;
wire n_1365;
wire n_253;
wire n_459;
wire n_1172;
wire n_998;
wire n_1276;
wire n_836;
wire n_1184;
wire n_583;
wire n_347;
wire n_414;
wire n_1336;
wire n_279;
wire n_776;
wire n_1138;
wire n_890;
wire n_1306;
wire n_1266;
wire n_497;
wire n_911;
wire n_450;
wire n_473;
wire n_967;
wire n_474;
wire n_1159;
wire n_1315;
wire n_1055;
wire n_611;
wire n_380;
wire n_844;
wire n_968;
wire n_710;
wire n_1040;
wire n_307;
wire n_1102;
wire n_661;
wire n_1185;
wire n_447;
wire n_403;
wire n_1039;
wire n_1119;
wire n_574;
wire n_1069;
wire n_842;
wire n_798;
wire n_668;
wire n_862;
wire n_869;
wire n_1066;
wire n_257;
wire n_285;
wire n_1377;
wire n_800;
wire n_778;
wire n_1175;
wire n_1170;
wire n_522;
wire n_977;
wire n_943;
wire n_287;
wire n_357;
wire n_905;
wire n_386;
wire n_878;
wire n_1333;
wire n_577;
wire n_759;
wire n_1235;
wire n_299;
wire n_322;
wire n_900;
wire n_841;
wire n_318;
wire n_1218;
wire n_736;
wire n_766;
wire n_852;
wire n_1268;
wire n_1113;
wire n_1089;
wire n_1122;
wire n_908;
wire n_1123;
wire n_923;
wire n_1302;
wire n_1289;
wire n_937;
wire n_773;
wire n_353;
wire n_865;
wire n_594;
wire n_856;
wire n_1146;
wire n_374;
wire n_932;
wire n_958;
wire n_775;
wire n_763;
wire n_1093;
wire n_427;
wire n_519;
wire n_1116;
wire n_709;
wire n_388;
wire n_332;
wire n_816;
wire n_625;
wire n_953;
wire n_289;
wire n_1373;
wire n_716;
wire n_356;
wire n_584;
wire n_896;
wire n_528;
wire n_1078;
wire n_495;
wire n_1072;
wire n_370;
wire n_352;
wire n_935;
wire n_467;
wire n_1213;
wire n_1053;
wire n_263;
wire n_515;
wire n_1019;
wire n_680;
wire n_1180;
wire n_904;
wire n_920;
wire n_1117;
wire n_284;
wire n_316;
wire n_1168;
wire n_1309;
wire n_909;
wire n_523;
wire n_996;
wire n_439;
wire n_506;
wire n_606;
wire n_513;
wire n_1332;
wire n_1263;
wire n_1115;
wire n_310;
wire n_725;
wire n_960;
wire n_671;
wire n_1084;
wire n_454;
wire n_1303;
wire n_443;
wire n_1029;
wire n_345;
wire n_1207;
wire n_324;
wire n_664;
wire n_367;
wire n_267;
wire n_1017;
wire n_581;
wire n_936;
wire n_1215;
wire n_582;
wire n_641;
wire n_940;
wire n_745;
wire n_339;
wire n_1167;
wire n_1327;
wire n_609;
wire n_1006;
wire n_1259;
wire n_350;
wire n_561;
wire n_437;
wire n_405;
wire n_1223;
wire n_621;
wire n_1012;
wire n_1241;
wire n_502;
wire n_769;
wire n_434;
wire n_250;
wire n_1212;
wire n_1054;
wire n_1308;
wire n_1050;
wire n_426;
wire n_1134;
wire n_1319;
wire n_1363;
wire n_616;
wire n_880;
wire n_1103;
wire n_1274;
wire n_832;
wire n_1321;
wire n_1060;
wire n_1154;
wire n_361;
wire n_632;
wire n_1344;
wire n_714;
wire n_1331;
wire n_1222;
wire n_1041;
wire n_251;
wire n_957;
wire n_1255;
wire n_995;
wire n_1124;
wire n_1335;
wire n_912;
wire n_464;
wire n_1227;
wire n_945;
wire n_392;
wire n_288;
wire n_274;
wire n_303;
wire n_563;
wire n_891;
wire n_568;
wire n_413;
wire n_1157;
wire n_902;
wire n_1158;
wire n_1079;
wire n_1330;
wire n_1033;
wire n_1028;
wire n_366;
wire n_1083;
wire n_727;
wire n_397;
wire n_1056;
wire n_663;
wire n_588;
wire n_707;
wire n_915;
wire n_1001;
wire n_711;
wire n_864;
wire n_1169;
wire n_377;
wire n_1139;
wire n_273;
wire n_1038;
wire n_276;
wire n_1085;
wire n_295;
wire n_845;
wire n_1127;
wire n_484;
wire n_326;
wire n_893;
wire n_1068;
wire n_747;
wire n_1244;
wire n_697;
wire n_978;
wire n_847;
wire n_826;
wire n_373;
wire n_628;
wire n_487;
wire n_831;
wire n_653;
wire n_692;
wire n_1051;
wire n_1355;
wire n_309;
wire n_827;
wire n_472;
wire n_866;
wire n_452;
wire n_262;
wire n_630;
wire n_820;
wire n_1208;
wire n_612;
wire n_858;
wire n_764;
wire n_252;
wire n_741;
wire n_1090;
wire n_456;
wire n_359;
wire n_1164;
wire n_433;
wire n_627;
wire n_418;
wire n_771;
wire n_1378;
wire n_524;
wire n_705;
wire n_1191;
wire n_1206;
wire n_1270;
wire n_546;
wire n_1010;
wire n_1375;
wire n_1015;
wire n_863;
wire n_525;
wire n_1226;
wire n_644;
wire n_1150;
wire n_1341;
wire n_833;
wire n_1229;
wire n_929;
wire n_1143;
wire n_1190;
wire n_543;
wire n_305;
wire n_585;
wire n_465;
wire n_1343;
wire n_719;
wire n_1156;
wire n_988;
wire n_921;
wire n_640;
wire n_1176;
wire n_1151;
wire n_1254;
wire n_646;
wire n_650;
wire n_1211;
wire n_743;
wire n_823;
wire n_393;
wire n_294;
wire n_1101;
wire n_1076;
wire n_1251;
wire n_1104;
wire n_1061;
wire n_849;
wire n_554;
wire n_1153;
wire n_1337;
wire n_797;
wire n_1177;
wire n_758;
wire n_436;
wire n_390;
wire n_1096;
wire n_1316;
wire n_1092;
wire n_846;
wire n_631;
wire n_673;
wire n_1067;
wire n_1292;
wire n_518;
wire n_1192;
wire n_1240;
wire n_987;
wire n_362;
wire n_1065;
wire n_540;
wire n_1064;
wire n_1075;
wire n_718;
wire n_669;
wire n_1091;
wire n_423;
wire n_1221;
wire n_458;
wire n_1200;
wire n_444;
wire n_319;
wire n_364;
wire n_555;
wire n_1295;
wire n_974;
wire n_1329;
wire n_857;
wire n_376;
wire n_308;
wire n_491;
wire n_1294;
wire n_1110;
wire n_1137;
wire n_460;
wire n_317;
wire n_321;
wire n_666;
wire n_320;
wire n_660;
wire n_1359;
wire n_886;
wire n_767;
wire n_889;
wire n_379;
wire n_1021;
wire n_1297;
wire n_1046;
wire n_1109;
wire n_961;
wire n_489;
wire n_1381;
wire n_573;
wire n_1099;
wire n_626;
wire n_539;
wire n_462;
wire n_280;
wire n_615;
wire n_1118;
wire n_990;
wire n_1108;
wire n_670;
wire n_818;
wire n_918;
wire n_1272;
wire n_408;
wire n_578;
wire n_372;
wire n_892;
wire n_938;
wire n_327;
wire n_774;
wire n_559;
wire n_1049;
wire n_466;
wire n_1277;
wire n_984;
wire n_301;
wire n_726;
wire n_369;
wire n_517;
wire n_931;
wire n_780;
wire n_530;
wire n_834;
wire n_693;
wire n_496;
wire n_1257;
wire n_1082;
wire n_1360;
wire n_468;
wire n_532;
wire n_1025;
wire n_298;
wire n_924;
wire n_1264;
wire n_297;
wire n_1245;
wire n_1152;
wire n_1081;
wire n_547;
wire n_1324;
wire n_1198;
wire n_304;
wire n_1307;
wire n_993;
wire n_819;
wire n_737;
wire n_1290;
wire n_1318;
wire n_1063;
wire n_1135;
wire n_828;
wire n_770;
wire n_867;
wire n_398;
wire n_1100;
wire n_425;
wire n_879;
wire n_331;
wire n_449;
wire n_1340;
wire n_607;
wire n_629;
wire n_706;
wire n_901;
wire n_876;
wire n_655;
wire n_654;
wire n_672;
wire n_567;
wire n_916;
wire n_1354;
wire n_1334;
wire n_1291;
wire n_986;
wire n_451;
wire n_1037;
wire n_1267;
wire n_790;
wire n_1262;
wire n_410;
wire n_751;
wire n_999;
wire n_913;
wire n_1237;
wire n_1356;
wire n_768;
wire n_412;
wire n_542;
wire n_1256;
wire n_1077;
wire n_1111;
wire n_1249;
wire n_387;
wire n_1239;
wire n_969;
wire n_256;
wire n_1009;
wire n_1202;
wire n_302;
wire n_604;
wire n_848;
wire n_756;
wire n_713;
wire n_598;
wire n_269;
wire n_430;
wire n_1252;
wire n_1132;
wire n_1275;
wire n_843;
wire n_579;
wire n_533;
wire n_385;
wire n_275;
wire n_536;
wire n_470;
wire n_851;
wire n_1155;
wire n_934;
wire n_1027;
wire n_965;
wire n_1296;
wire n_382;
wire n_1043;
wire n_435;
wire n_511;
wire n_509;
wire n_1204;
wire n_930;
wire n_1265;
wire n_1057;
wire n_907;
wire n_1005;
wire n_1312;
wire n_899;
wire n_637;
wire n_544;
wire n_1087;
wire n_344;
wire n_482;
wire n_633;
wire n_971;
wire n_1052;
wire n_1071;
wire n_1311;
wire n_1273;
wire n_959;
wire n_349;
wire n_336;
wire n_1130;
wire n_794;
wire n_283;
wire n_314;
wire n_1228;
wire n_681;
wire n_982;
wire n_717;
wire n_1253;
wire n_312;
wire n_1183;
wire n_335;
wire n_516;
wire n_521;
wire n_1195;
wire n_1300;
wire n_575;
wire n_338;
wire n_1372;
wire n_698;
wire n_371;
wire n_1345;
wire n_587;
wire n_1246;
wire n_1074;
wire n_674;
wire n_888;
wire n_793;
wire n_272;
wire n_757;
wire n_803;
wire n_514;
wire n_507;
wire n_270;
wire n_614;
wire n_772;
wire n_1114;
wire n_566;
wire n_871;
wire n_1088;
wire n_1230;
wire n_1326;
wire n_340;
wire n_483;
wire n_1352;
wire n_729;
wire n_1280;
wire n_1323;
wire n_394;
wire n_1097;
wire n_703;
wire n_1369;
wire n_601;
wire n_463;
wire n_396;
wire n_1236;
wire n_342;
wire n_348;
wire n_603;
wire n_1288;
wire n_868;
wire n_1024;
wire n_259;
wire n_1144;
wire n_475;
wire n_897;
wire n_1320;
wire n_855;
wire n_429;
AOI22xp33_ASAP7_75t_SL g744 ( .A1(n_0), .A2(n_74), .B1(n_535), .B2(n_741), .Y(n_744) );
AOI22xp33_ASAP7_75t_L g758 ( .A1(n_0), .A2(n_229), .B1(n_398), .B2(n_452), .Y(n_758) );
AOI22xp33_ASAP7_75t_L g503 ( .A1(n_1), .A2(n_196), .B1(n_398), .B2(n_504), .Y(n_503) );
AOI22xp33_ASAP7_75t_L g530 ( .A1(n_1), .A2(n_66), .B1(n_330), .B2(n_531), .Y(n_530) );
INVx1_ASAP7_75t_L g347 ( .A(n_2), .Y(n_347) );
AOI22xp33_ASAP7_75t_L g394 ( .A1(n_2), .A2(n_101), .B1(n_395), .B2(n_398), .Y(n_394) );
INVx1_ASAP7_75t_L g749 ( .A(n_3), .Y(n_749) );
OAI211xp5_ASAP7_75t_L g834 ( .A1(n_4), .A2(n_835), .B(n_836), .C(n_843), .Y(n_834) );
NOR2xp33_ASAP7_75t_L g854 ( .A(n_4), .B(n_521), .Y(n_854) );
AOI22xp33_ASAP7_75t_L g781 ( .A1(n_5), .A2(n_119), .B1(n_543), .B2(n_782), .Y(n_781) );
AOI22xp33_ASAP7_75t_SL g800 ( .A1(n_5), .A2(n_125), .B1(n_452), .B2(n_801), .Y(n_800) );
AOI22xp5_ASAP7_75t_SL g1113 ( .A1(n_6), .A2(n_232), .B1(n_1097), .B2(n_1099), .Y(n_1113) );
INVx1_ASAP7_75t_L g516 ( .A(n_7), .Y(n_516) );
OAI22xp33_ASAP7_75t_L g544 ( .A1(n_7), .A2(n_69), .B1(n_545), .B2(n_551), .Y(n_544) );
AOI22xp33_ASAP7_75t_L g1035 ( .A1(n_8), .A2(n_77), .B1(n_741), .B2(n_1036), .Y(n_1035) );
AOI22xp33_ASAP7_75t_L g1055 ( .A1(n_8), .A2(n_52), .B1(n_1056), .B2(n_1057), .Y(n_1055) );
AOI22xp33_ASAP7_75t_L g566 ( .A1(n_9), .A2(n_205), .B1(n_398), .B2(n_504), .Y(n_566) );
AOI22xp33_ASAP7_75t_L g585 ( .A1(n_9), .A2(n_234), .B1(n_330), .B2(n_586), .Y(n_585) );
AOI221xp5_ASAP7_75t_L g1278 ( .A1(n_10), .A2(n_109), .B1(n_389), .B2(n_449), .C(n_572), .Y(n_1278) );
INVx1_ASAP7_75t_L g1299 ( .A(n_10), .Y(n_1299) );
INVx1_ASAP7_75t_L g900 ( .A(n_11), .Y(n_900) );
AO22x1_ASAP7_75t_L g933 ( .A1(n_11), .A2(n_143), .B1(n_379), .B2(n_841), .Y(n_933) );
INVx1_ASAP7_75t_L g259 ( .A(n_12), .Y(n_259) );
AND2x2_ASAP7_75t_L g298 ( .A(n_12), .B(n_212), .Y(n_298) );
AND2x2_ASAP7_75t_L g382 ( .A(n_12), .B(n_383), .Y(n_382) );
NOR2xp33_ASAP7_75t_L g635 ( .A(n_12), .B(n_269), .Y(n_635) );
INVx1_ASAP7_75t_L g910 ( .A(n_13), .Y(n_910) );
AOI22xp33_ASAP7_75t_L g932 ( .A1(n_13), .A2(n_99), .B1(n_390), .B2(n_839), .Y(n_932) );
AOI221xp5_ASAP7_75t_L g742 ( .A1(n_14), .A2(n_142), .B1(n_482), .B2(n_738), .C(n_743), .Y(n_742) );
AOI22xp33_ASAP7_75t_L g761 ( .A1(n_14), .A2(n_61), .B1(n_398), .B2(n_762), .Y(n_761) );
AOI22xp33_ASAP7_75t_SL g779 ( .A1(n_15), .A2(n_151), .B1(n_437), .B2(n_780), .Y(n_779) );
AOI221xp5_ASAP7_75t_L g796 ( .A1(n_15), .A2(n_19), .B1(n_392), .B2(n_797), .C(n_798), .Y(n_796) );
INVx2_ASAP7_75t_L g1092 ( .A(n_16), .Y(n_1092) );
AND2x2_ASAP7_75t_L g1095 ( .A(n_16), .B(n_1093), .Y(n_1095) );
AND2x2_ASAP7_75t_L g1100 ( .A(n_16), .B(n_105), .Y(n_1100) );
OAI22xp5_ASAP7_75t_L g579 ( .A1(n_17), .A2(n_91), .B1(n_304), .B2(n_521), .Y(n_579) );
CKINVDCx5p33_ASAP7_75t_R g735 ( .A(n_18), .Y(n_735) );
AOI22xp33_ASAP7_75t_SL g786 ( .A1(n_19), .A2(n_33), .B1(n_532), .B2(n_538), .Y(n_786) );
XOR2xp5_ASAP7_75t_L g1326 ( .A(n_20), .B(n_1327), .Y(n_1326) );
INVx1_ASAP7_75t_L g775 ( .A(n_21), .Y(n_775) );
OAI22xp33_ASAP7_75t_L g787 ( .A1(n_22), .A2(n_199), .B1(n_545), .B2(n_788), .Y(n_787) );
INVx1_ASAP7_75t_L g804 ( .A(n_22), .Y(n_804) );
XNOR2xp5_ASAP7_75t_L g442 ( .A(n_23), .B(n_443), .Y(n_442) );
AOI22xp5_ASAP7_75t_SL g1105 ( .A1(n_23), .A2(n_133), .B1(n_1097), .B2(n_1099), .Y(n_1105) );
INVx1_ASAP7_75t_L g404 ( .A(n_24), .Y(n_404) );
AOI22xp33_ASAP7_75t_SL g348 ( .A1(n_25), .A2(n_75), .B1(n_349), .B2(n_351), .Y(n_348) );
AOI221xp5_ASAP7_75t_L g385 ( .A1(n_25), .A2(n_245), .B1(n_386), .B2(n_389), .C(n_392), .Y(n_385) );
AOI22xp5_ASAP7_75t_SL g1117 ( .A1(n_26), .A2(n_225), .B1(n_1094), .B2(n_1118), .Y(n_1117) );
INVx1_ASAP7_75t_L g401 ( .A(n_27), .Y(n_401) );
OAI211xp5_ASAP7_75t_L g844 ( .A1(n_28), .A2(n_639), .B(n_845), .C(n_846), .Y(n_844) );
INVx1_ASAP7_75t_L g877 ( .A(n_28), .Y(n_877) );
AOI22xp33_ASAP7_75t_L g1279 ( .A1(n_29), .A2(n_78), .B1(n_398), .B2(n_452), .Y(n_1279) );
INVx1_ASAP7_75t_L g1304 ( .A(n_29), .Y(n_1304) );
OAI22xp5_ASAP7_75t_L g520 ( .A1(n_30), .A2(n_94), .B1(n_304), .B2(n_521), .Y(n_520) );
AOI22xp33_ASAP7_75t_L g364 ( .A1(n_31), .A2(n_245), .B1(n_349), .B2(n_351), .Y(n_364) );
AOI22xp33_ASAP7_75t_SL g425 ( .A1(n_31), .A2(n_75), .B1(n_426), .B2(n_428), .Y(n_425) );
OAI22xp5_ASAP7_75t_L g674 ( .A1(n_32), .A2(n_237), .B1(n_675), .B2(n_679), .Y(n_674) );
OAI22xp33_ASAP7_75t_L g713 ( .A1(n_32), .A2(n_237), .B1(n_714), .B2(n_717), .Y(n_713) );
A2O1A1Ixp33_ASAP7_75t_L g807 ( .A1(n_33), .A2(n_808), .B(n_809), .C(n_820), .Y(n_807) );
NAND2xp5_ASAP7_75t_SL g987 ( .A(n_34), .B(n_988), .Y(n_987) );
AOI22xp33_ASAP7_75t_L g1011 ( .A1(n_34), .A2(n_152), .B1(n_1006), .B2(n_1012), .Y(n_1011) );
XNOR2xp5_ASAP7_75t_L g555 ( .A(n_35), .B(n_556), .Y(n_555) );
AOI22xp33_ASAP7_75t_L g992 ( .A1(n_36), .A2(n_152), .B1(n_379), .B2(n_397), .Y(n_992) );
AOI22xp33_ASAP7_75t_L g1005 ( .A1(n_36), .A2(n_223), .B1(n_532), .B2(n_1006), .Y(n_1005) );
INVx1_ASAP7_75t_L g498 ( .A(n_37), .Y(n_498) );
AOI22xp5_ASAP7_75t_L g1136 ( .A1(n_38), .A2(n_165), .B1(n_1089), .B2(n_1094), .Y(n_1136) );
AOI22xp33_ASAP7_75t_L g1283 ( .A1(n_39), .A2(n_208), .B1(n_395), .B2(n_453), .Y(n_1283) );
AOI22xp33_ASAP7_75t_L g1305 ( .A1(n_39), .A2(n_109), .B1(n_862), .B2(n_1306), .Y(n_1305) );
OAI22xp5_ASAP7_75t_L g791 ( .A1(n_40), .A2(n_59), .B1(n_521), .B2(n_792), .Y(n_791) );
OAI211xp5_ASAP7_75t_L g794 ( .A1(n_40), .A2(n_506), .B(n_795), .C(n_802), .Y(n_794) );
AOI22xp33_ASAP7_75t_L g1159 ( .A1(n_41), .A2(n_93), .B1(n_1097), .B2(n_1123), .Y(n_1159) );
AOI22xp33_ASAP7_75t_L g573 ( .A1(n_42), .A2(n_159), .B1(n_398), .B2(n_511), .Y(n_573) );
AOI22xp33_ASAP7_75t_SL g589 ( .A1(n_42), .A2(n_121), .B1(n_440), .B2(n_535), .Y(n_589) );
AOI21xp33_ASAP7_75t_L g464 ( .A1(n_43), .A2(n_386), .B(n_465), .Y(n_464) );
INVx1_ASAP7_75t_L g475 ( .A(n_43), .Y(n_475) );
XNOR2x2_ASAP7_75t_L g768 ( .A(n_44), .B(n_769), .Y(n_768) );
AOI22xp5_ASAP7_75t_L g1108 ( .A1(n_44), .A2(n_87), .B1(n_1089), .B2(n_1097), .Y(n_1108) );
AOI22xp5_ASAP7_75t_L g1137 ( .A1(n_45), .A2(n_169), .B1(n_1097), .B2(n_1118), .Y(n_1137) );
AOI22xp33_ASAP7_75t_L g837 ( .A1(n_46), .A2(n_68), .B1(n_397), .B2(n_453), .Y(n_837) );
AOI22xp33_ASAP7_75t_SL g857 ( .A1(n_46), .A2(n_243), .B1(n_349), .B2(n_351), .Y(n_857) );
AOI22xp33_ASAP7_75t_SL g1041 ( .A1(n_47), .A2(n_129), .B1(n_591), .B2(n_1042), .Y(n_1041) );
INVxp67_ASAP7_75t_SL g1073 ( .A(n_47), .Y(n_1073) );
INVx1_ASAP7_75t_L g287 ( .A(n_48), .Y(n_287) );
INVx1_ASAP7_75t_L g321 ( .A(n_48), .Y(n_321) );
INVx1_ASAP7_75t_L g302 ( .A(n_49), .Y(n_302) );
AOI22xp33_ASAP7_75t_L g451 ( .A1(n_50), .A2(n_190), .B1(n_452), .B2(n_453), .Y(n_451) );
INVx1_ASAP7_75t_L g476 ( .A(n_50), .Y(n_476) );
INVx1_ASAP7_75t_L g975 ( .A(n_51), .Y(n_975) );
AOI22xp33_ASAP7_75t_L g1038 ( .A1(n_52), .A2(n_135), .B1(n_741), .B2(n_1039), .Y(n_1038) );
AOI22xp5_ASAP7_75t_L g1088 ( .A1(n_53), .A2(n_241), .B1(n_1089), .B2(n_1094), .Y(n_1088) );
AOI22xp33_ASAP7_75t_L g784 ( .A1(n_54), .A2(n_125), .B1(n_543), .B2(n_618), .Y(n_784) );
AOI221xp5_ASAP7_75t_L g810 ( .A1(n_54), .A2(n_119), .B1(n_811), .B2(n_814), .C(n_817), .Y(n_810) );
INVx1_ASAP7_75t_L g1288 ( .A(n_55), .Y(n_1288) );
INVx1_ASAP7_75t_L g253 ( .A(n_56), .Y(n_253) );
AOI221xp5_ASAP7_75t_L g447 ( .A1(n_57), .A2(n_215), .B1(n_392), .B2(n_448), .C(n_449), .Y(n_447) );
AOI22xp33_ASAP7_75t_L g477 ( .A1(n_57), .A2(n_244), .B1(n_330), .B2(n_349), .Y(n_477) );
INVx2_ASAP7_75t_L g293 ( .A(n_58), .Y(n_293) );
INVx1_ASAP7_75t_L g964 ( .A(n_60), .Y(n_964) );
AOI221xp5_ASAP7_75t_L g737 ( .A1(n_61), .A2(n_72), .B1(n_538), .B2(n_738), .C(n_739), .Y(n_737) );
AOI221xp5_ASAP7_75t_L g1333 ( .A1(n_62), .A2(n_117), .B1(n_570), .B2(n_572), .C(n_1334), .Y(n_1333) );
INVx1_ASAP7_75t_L g1371 ( .A(n_62), .Y(n_1371) );
INVx1_ASAP7_75t_L g1046 ( .A(n_63), .Y(n_1046) );
AOI22xp5_ASAP7_75t_L g1119 ( .A1(n_64), .A2(n_70), .B1(n_1089), .B2(n_1097), .Y(n_1119) );
INVx1_ASAP7_75t_L g731 ( .A(n_65), .Y(n_731) );
AOI221xp5_ASAP7_75t_L g508 ( .A1(n_66), .A2(n_187), .B1(n_389), .B2(n_392), .C(n_509), .Y(n_508) );
INVx1_ASAP7_75t_L g730 ( .A(n_67), .Y(n_730) );
AOI22xp33_ASAP7_75t_SL g861 ( .A1(n_68), .A2(n_98), .B1(n_349), .B2(n_862), .Y(n_861) );
INVx1_ASAP7_75t_L g513 ( .A(n_69), .Y(n_513) );
AOI22xp33_ASAP7_75t_L g1341 ( .A1(n_71), .A2(n_130), .B1(n_452), .B2(n_1337), .Y(n_1341) );
INVx1_ASAP7_75t_L g1359 ( .A(n_71), .Y(n_1359) );
AOI221xp5_ASAP7_75t_L g754 ( .A1(n_72), .A2(n_142), .B1(n_389), .B2(n_755), .C(n_757), .Y(n_754) );
INVx1_ASAP7_75t_L g1014 ( .A(n_73), .Y(n_1014) );
AOI221xp5_ASAP7_75t_L g763 ( .A1(n_74), .A2(n_80), .B1(n_423), .B2(n_448), .C(n_755), .Y(n_763) );
AOI221xp5_ASAP7_75t_L g1282 ( .A1(n_76), .A2(n_108), .B1(n_386), .B2(n_389), .C(n_465), .Y(n_1282) );
INVxp67_ASAP7_75t_SL g1291 ( .A(n_76), .Y(n_1291) );
INVx1_ASAP7_75t_L g1068 ( .A(n_77), .Y(n_1068) );
INVxp67_ASAP7_75t_SL g1293 ( .A(n_78), .Y(n_1293) );
AOI21xp33_ASAP7_75t_L g502 ( .A1(n_79), .A2(n_449), .B(n_465), .Y(n_502) );
AOI22xp33_ASAP7_75t_L g533 ( .A1(n_79), .A2(n_163), .B1(n_534), .B2(n_535), .Y(n_533) );
AOI22xp33_ASAP7_75t_SL g740 ( .A1(n_80), .A2(n_229), .B1(n_535), .B2(n_741), .Y(n_740) );
AOI22xp5_ASAP7_75t_L g1107 ( .A1(n_81), .A2(n_178), .B1(n_1094), .B2(n_1099), .Y(n_1107) );
OAI211xp5_ASAP7_75t_L g494 ( .A1(n_82), .A2(n_408), .B(n_495), .C(n_499), .Y(n_494) );
INVx1_ASAP7_75t_L g526 ( .A(n_82), .Y(n_526) );
CKINVDCx5p33_ASAP7_75t_R g612 ( .A(n_83), .Y(n_612) );
OAI222xp33_ASAP7_75t_L g919 ( .A1(n_84), .A2(n_197), .B1(n_920), .B2(n_922), .C1(n_924), .C2(n_926), .Y(n_919) );
INVx1_ASAP7_75t_L g937 ( .A(n_84), .Y(n_937) );
OAI22xp5_ASAP7_75t_SL g983 ( .A1(n_85), .A2(n_103), .B1(n_643), .B2(n_648), .Y(n_983) );
OAI21xp33_ASAP7_75t_L g994 ( .A1(n_85), .A2(n_551), .B(n_995), .Y(n_994) );
INVx1_ASAP7_75t_L g1028 ( .A(n_86), .Y(n_1028) );
OAI222xp33_ASAP7_75t_L g1060 ( .A1(n_86), .A2(n_123), .B1(n_1061), .B2(n_1062), .C1(n_1069), .C2(n_1075), .Y(n_1060) );
INVx1_ASAP7_75t_L g1343 ( .A(n_88), .Y(n_1343) );
INVx1_ASAP7_75t_L g560 ( .A(n_89), .Y(n_560) );
CKINVDCx5p33_ASAP7_75t_R g904 ( .A(n_90), .Y(n_904) );
OAI211xp5_ASAP7_75t_L g567 ( .A1(n_91), .A2(n_377), .B(n_568), .C(n_574), .Y(n_567) );
HB1xp67_ASAP7_75t_L g255 ( .A(n_92), .Y(n_255) );
AND2x2_ASAP7_75t_L g1090 ( .A(n_92), .B(n_253), .Y(n_1090) );
INVx1_ASAP7_75t_L g1315 ( .A(n_93), .Y(n_1315) );
AOI22xp33_ASAP7_75t_L g1322 ( .A1(n_93), .A2(n_1323), .B1(n_1325), .B2(n_1378), .Y(n_1322) );
OAI211xp5_ASAP7_75t_SL g505 ( .A1(n_94), .A2(n_506), .B(n_507), .C(n_512), .Y(n_505) );
CKINVDCx5p33_ASAP7_75t_R g734 ( .A(n_95), .Y(n_734) );
CKINVDCx5p33_ASAP7_75t_R g890 ( .A(n_96), .Y(n_890) );
CKINVDCx5p33_ASAP7_75t_R g460 ( .A(n_97), .Y(n_460) );
AOI221xp5_ASAP7_75t_SL g842 ( .A1(n_98), .A2(n_243), .B1(n_390), .B2(n_757), .C(n_815), .Y(n_842) );
INVx1_ASAP7_75t_L g906 ( .A(n_99), .Y(n_906) );
CKINVDCx5p33_ASAP7_75t_R g360 ( .A(n_100), .Y(n_360) );
INVx1_ASAP7_75t_L g363 ( .A(n_101), .Y(n_363) );
OAI211xp5_ASAP7_75t_L g977 ( .A1(n_102), .A2(n_978), .B(n_979), .C(n_980), .Y(n_977) );
INVxp33_ASAP7_75t_SL g996 ( .A(n_102), .Y(n_996) );
INVxp67_ASAP7_75t_SL g1018 ( .A(n_103), .Y(n_1018) );
CKINVDCx5p33_ASAP7_75t_R g1023 ( .A(n_104), .Y(n_1023) );
INVx1_ASAP7_75t_L g1093 ( .A(n_105), .Y(n_1093) );
AND2x2_ASAP7_75t_L g1098 ( .A(n_105), .B(n_1092), .Y(n_1098) );
CKINVDCx5p33_ASAP7_75t_R g850 ( .A(n_106), .Y(n_850) );
AOI22xp5_ASAP7_75t_L g1114 ( .A1(n_107), .A2(n_177), .B1(n_1089), .B2(n_1094), .Y(n_1114) );
INVx1_ASAP7_75t_L g1302 ( .A(n_108), .Y(n_1302) );
INVx1_ASAP7_75t_L g1346 ( .A(n_110), .Y(n_1346) );
INVx1_ASAP7_75t_L g342 ( .A(n_111), .Y(n_342) );
AOI21xp33_ASAP7_75t_L g422 ( .A1(n_111), .A2(n_386), .B(n_423), .Y(n_422) );
CKINVDCx5p33_ASAP7_75t_R g631 ( .A(n_112), .Y(n_631) );
NAND2xp5_ASAP7_75t_L g292 ( .A(n_113), .B(n_293), .Y(n_292) );
INVx2_ASAP7_75t_L g325 ( .A(n_113), .Y(n_325) );
INVx1_ASAP7_75t_L g356 ( .A(n_113), .Y(n_356) );
AOI21xp33_ASAP7_75t_L g563 ( .A1(n_114), .A2(n_564), .B(n_565), .Y(n_563) );
AOI22xp33_ASAP7_75t_L g588 ( .A1(n_114), .A2(n_159), .B1(n_534), .B2(n_535), .Y(n_588) );
OAI22xp33_ASAP7_75t_L g684 ( .A1(n_115), .A2(n_166), .B1(n_685), .B2(n_686), .Y(n_684) );
OAI22xp33_ASAP7_75t_L g692 ( .A1(n_115), .A2(n_166), .B1(n_693), .B2(n_696), .Y(n_692) );
OAI22xp5_ASAP7_75t_L g853 ( .A1(n_116), .A2(n_136), .B1(n_501), .B2(n_639), .Y(n_853) );
INVx1_ASAP7_75t_L g865 ( .A(n_116), .Y(n_865) );
INVx1_ASAP7_75t_L g1360 ( .A(n_117), .Y(n_1360) );
INVx1_ASAP7_75t_L g914 ( .A(n_118), .Y(n_914) );
NAND2xp33_ASAP7_75t_SL g954 ( .A(n_118), .B(n_390), .Y(n_954) );
NOR2xp33_ASAP7_75t_L g1377 ( .A(n_120), .B(n_281), .Y(n_1377) );
INVxp67_ASAP7_75t_SL g562 ( .A(n_121), .Y(n_562) );
OAI22xp5_ASAP7_75t_L g303 ( .A1(n_122), .A2(n_213), .B1(n_304), .B2(n_315), .Y(n_303) );
OAI211xp5_ASAP7_75t_L g376 ( .A1(n_122), .A2(n_377), .B(n_384), .C(n_400), .Y(n_376) );
INVx1_ASAP7_75t_L g1027 ( .A(n_123), .Y(n_1027) );
INVx1_ASAP7_75t_L g578 ( .A(n_124), .Y(n_578) );
CKINVDCx5p33_ASAP7_75t_R g614 ( .A(n_126), .Y(n_614) );
NOR2xp33_ASAP7_75t_L g1285 ( .A(n_127), .B(n_412), .Y(n_1285) );
INVxp67_ASAP7_75t_SL g1312 ( .A(n_127), .Y(n_1312) );
OAI211xp5_ASAP7_75t_SL g662 ( .A1(n_128), .A2(n_655), .B(n_663), .C(n_666), .Y(n_662) );
INVx1_ASAP7_75t_L g712 ( .A(n_128), .Y(n_712) );
AOI221xp5_ASAP7_75t_L g1052 ( .A1(n_129), .A2(n_238), .B1(n_572), .B2(n_1053), .C(n_1054), .Y(n_1052) );
INVx1_ASAP7_75t_L g1367 ( .A(n_130), .Y(n_1367) );
INVx1_ASAP7_75t_L g576 ( .A(n_131), .Y(n_576) );
OAI22xp33_ASAP7_75t_L g592 ( .A1(n_131), .A2(n_172), .B1(n_551), .B2(n_593), .Y(n_592) );
CKINVDCx5p33_ASAP7_75t_R g624 ( .A(n_132), .Y(n_624) );
INVx1_ASAP7_75t_L g456 ( .A(n_134), .Y(n_456) );
INVx1_ASAP7_75t_L g1064 ( .A(n_135), .Y(n_1064) );
INVx1_ASAP7_75t_L g875 ( .A(n_136), .Y(n_875) );
INVx1_ASAP7_75t_L g1158 ( .A(n_137), .Y(n_1158) );
CKINVDCx16_ASAP7_75t_R g921 ( .A(n_138), .Y(n_921) );
INVx1_ASAP7_75t_L g1284 ( .A(n_139), .Y(n_1284) );
NAND5xp2_ASAP7_75t_L g832 ( .A(n_140), .B(n_833), .C(n_855), .D(n_866), .E(n_873), .Y(n_832) );
INVx1_ASAP7_75t_L g881 ( .A(n_140), .Y(n_881) );
AOI22xp33_ASAP7_75t_SL g466 ( .A1(n_141), .A2(n_244), .B1(n_379), .B2(n_426), .Y(n_466) );
AOI22xp33_ASAP7_75t_L g481 ( .A1(n_141), .A2(n_215), .B1(n_349), .B2(n_482), .Y(n_481) );
AOI21xp5_ASAP7_75t_L g915 ( .A1(n_143), .A2(n_541), .B(n_916), .Y(n_915) );
INVx1_ASAP7_75t_L g958 ( .A(n_144), .Y(n_958) );
INVx1_ASAP7_75t_L g1287 ( .A(n_145), .Y(n_1287) );
OAI322xp33_ASAP7_75t_L g1289 ( .A1(n_145), .A2(n_551), .A3(n_603), .B1(n_1007), .B2(n_1290), .C1(n_1294), .C2(n_1300), .Y(n_1289) );
INVx1_ASAP7_75t_L g455 ( .A(n_146), .Y(n_455) );
AOI22xp5_ASAP7_75t_L g1122 ( .A1(n_147), .A2(n_173), .B1(n_1097), .B2(n_1123), .Y(n_1122) );
CKINVDCx5p33_ASAP7_75t_R g629 ( .A(n_148), .Y(n_629) );
BUFx3_ASAP7_75t_L g286 ( .A(n_149), .Y(n_286) );
INVx1_ASAP7_75t_L g1275 ( .A(n_150), .Y(n_1275) );
NAND2xp5_ASAP7_75t_L g818 ( .A(n_151), .B(n_819), .Y(n_818) );
AOI22xp5_ASAP7_75t_L g1121 ( .A1(n_153), .A2(n_188), .B1(n_1089), .B2(n_1094), .Y(n_1121) );
AOI221xp5_ASAP7_75t_L g569 ( .A1(n_154), .A2(n_234), .B1(n_389), .B2(n_570), .C(n_572), .Y(n_569) );
AOI22xp33_ASAP7_75t_L g590 ( .A1(n_154), .A2(n_205), .B1(n_538), .B2(n_591), .Y(n_590) );
INVx1_ASAP7_75t_L g1350 ( .A(n_155), .Y(n_1350) );
OAI21xp33_ASAP7_75t_L g1044 ( .A1(n_156), .A2(n_792), .B(n_1045), .Y(n_1044) );
AOI22xp5_ASAP7_75t_L g1096 ( .A1(n_157), .A2(n_202), .B1(n_1097), .B2(n_1099), .Y(n_1096) );
BUFx6f_ASAP7_75t_L g266 ( .A(n_158), .Y(n_266) );
AOI22xp33_ASAP7_75t_L g840 ( .A1(n_160), .A2(n_195), .B1(n_453), .B2(n_841), .Y(n_840) );
AOI22xp33_ASAP7_75t_L g859 ( .A1(n_160), .A2(n_189), .B1(n_535), .B2(n_860), .Y(n_859) );
INVx1_ASAP7_75t_L g750 ( .A(n_161), .Y(n_750) );
CKINVDCx5p33_ASAP7_75t_R g670 ( .A(n_162), .Y(n_670) );
AOI22xp33_ASAP7_75t_L g510 ( .A1(n_163), .A2(n_226), .B1(n_398), .B2(n_511), .Y(n_510) );
OAI21xp5_ASAP7_75t_SL g764 ( .A1(n_164), .A2(n_304), .B(n_765), .Y(n_764) );
CKINVDCx5p33_ASAP7_75t_R g1309 ( .A(n_167), .Y(n_1309) );
INVx1_ASAP7_75t_L g1047 ( .A(n_168), .Y(n_1047) );
CKINVDCx5p33_ASAP7_75t_R g608 ( .A(n_170), .Y(n_608) );
INVx1_ASAP7_75t_L g892 ( .A(n_171), .Y(n_892) );
NOR2xp33_ASAP7_75t_L g894 ( .A(n_171), .B(n_895), .Y(n_894) );
INVx1_ASAP7_75t_L g575 ( .A(n_172), .Y(n_575) );
INVx1_ASAP7_75t_L g1031 ( .A(n_174), .Y(n_1031) );
INVx1_ASAP7_75t_L g1280 ( .A(n_175), .Y(n_1280) );
OAI221xp5_ASAP7_75t_L g457 ( .A1(n_176), .A2(n_216), .B1(n_412), .B2(n_458), .C(n_459), .Y(n_457) );
OAI22xp33_ASAP7_75t_L g484 ( .A1(n_176), .A2(n_216), .B1(n_366), .B2(n_369), .Y(n_484) );
AOI21xp33_ASAP7_75t_L g991 ( .A1(n_179), .A2(n_386), .B(n_565), .Y(n_991) );
INVx1_ASAP7_75t_L g1002 ( .A(n_179), .Y(n_1002) );
INVx1_ASAP7_75t_L g671 ( .A(n_180), .Y(n_671) );
OAI211xp5_ASAP7_75t_L g699 ( .A1(n_180), .A2(n_700), .B(n_702), .C(n_704), .Y(n_699) );
XOR2x2_ASAP7_75t_L g599 ( .A(n_181), .B(n_600), .Y(n_599) );
INVx1_ASAP7_75t_L g872 ( .A(n_182), .Y(n_872) );
OAI211xp5_ASAP7_75t_L g1331 ( .A1(n_183), .A2(n_1061), .B(n_1332), .C(n_1338), .Y(n_1331) );
INVx1_ASAP7_75t_L g1374 ( .A(n_183), .Y(n_1374) );
AOI221xp5_ASAP7_75t_L g1342 ( .A1(n_184), .A2(n_230), .B1(n_389), .B2(n_449), .C(n_817), .Y(n_1342) );
INVx1_ASAP7_75t_L g1353 ( .A(n_184), .Y(n_1353) );
INVx1_ASAP7_75t_L g1348 ( .A(n_185), .Y(n_1348) );
OAI332xp33_ASAP7_75t_SL g1351 ( .A1(n_185), .A2(n_472), .A3(n_540), .B1(n_545), .B2(n_1352), .B3(n_1358), .C1(n_1363), .C2(n_1366), .Y(n_1351) );
BUFx6f_ASAP7_75t_L g265 ( .A(n_186), .Y(n_265) );
AOI22xp33_ASAP7_75t_L g537 ( .A1(n_187), .A2(n_196), .B1(n_531), .B2(n_538), .Y(n_537) );
AOI221xp5_ASAP7_75t_L g838 ( .A1(n_189), .A2(n_221), .B1(n_390), .B2(n_565), .C(n_839), .Y(n_838) );
INVx1_ASAP7_75t_L g480 ( .A(n_190), .Y(n_480) );
XOR2x2_ASAP7_75t_L g970 ( .A(n_191), .B(n_971), .Y(n_970) );
CKINVDCx5p33_ASAP7_75t_R g790 ( .A(n_192), .Y(n_790) );
AOI22xp33_ASAP7_75t_SL g986 ( .A1(n_193), .A2(n_231), .B1(n_379), .B2(n_762), .Y(n_986) );
INVx1_ASAP7_75t_L g1004 ( .A(n_193), .Y(n_1004) );
INVxp67_ASAP7_75t_SL g500 ( .A(n_194), .Y(n_500) );
AOI22xp33_ASAP7_75t_SL g542 ( .A1(n_194), .A2(n_226), .B1(n_440), .B2(n_543), .Y(n_542) );
AOI22xp33_ASAP7_75t_L g858 ( .A1(n_195), .A2(n_221), .B1(n_535), .B2(n_741), .Y(n_858) );
NOR2xp33_ASAP7_75t_R g944 ( .A(n_197), .B(n_945), .Y(n_944) );
OA22x2_ASAP7_75t_L g491 ( .A1(n_198), .A2(n_492), .B1(n_553), .B2(n_554), .Y(n_491) );
CKINVDCx16_ASAP7_75t_R g553 ( .A(n_198), .Y(n_553) );
INVx1_ASAP7_75t_L g803 ( .A(n_199), .Y(n_803) );
CKINVDCx5p33_ASAP7_75t_R g605 ( .A(n_200), .Y(n_605) );
INVx1_ASAP7_75t_L g773 ( .A(n_201), .Y(n_773) );
INVx1_ASAP7_75t_L g886 ( .A(n_202), .Y(n_886) );
OAI22xp5_ASAP7_75t_L g487 ( .A1(n_203), .A2(n_246), .B1(n_304), .B2(n_315), .Y(n_487) );
AOI22xp33_ASAP7_75t_L g1336 ( .A1(n_204), .A2(n_217), .B1(n_452), .B2(n_1337), .Y(n_1336) );
INVx1_ASAP7_75t_L g1365 ( .A(n_204), .Y(n_1365) );
AOI22xp33_ASAP7_75t_SL g1034 ( .A1(n_206), .A2(n_238), .B1(n_482), .B2(n_586), .Y(n_1034) );
INVxp67_ASAP7_75t_SL g1070 ( .A(n_206), .Y(n_1070) );
INVx1_ASAP7_75t_L g486 ( .A(n_207), .Y(n_486) );
INVxp67_ASAP7_75t_SL g1295 ( .A(n_208), .Y(n_1295) );
OAI211xp5_ASAP7_75t_L g558 ( .A1(n_209), .A2(n_408), .B(n_559), .C(n_561), .Y(n_558) );
INVx1_ASAP7_75t_L g583 ( .A(n_209), .Y(n_583) );
CKINVDCx5p33_ASAP7_75t_R g982 ( .A(n_210), .Y(n_982) );
INVx1_ASAP7_75t_L g1345 ( .A(n_211), .Y(n_1345) );
BUFx3_ASAP7_75t_L g269 ( .A(n_212), .Y(n_269) );
INVx1_ASAP7_75t_L g383 ( .A(n_212), .Y(n_383) );
CKINVDCx5p33_ASAP7_75t_R g847 ( .A(n_214), .Y(n_847) );
INVx1_ASAP7_75t_L g1355 ( .A(n_217), .Y(n_1355) );
CKINVDCx5p33_ASAP7_75t_R g621 ( .A(n_218), .Y(n_621) );
INVx1_ASAP7_75t_L g291 ( .A(n_219), .Y(n_291) );
INVx1_ASAP7_75t_L g296 ( .A(n_219), .Y(n_296) );
INVx2_ASAP7_75t_L g434 ( .A(n_219), .Y(n_434) );
XNOR2x1_ASAP7_75t_L g726 ( .A(n_220), .B(n_727), .Y(n_726) );
INVx1_ASAP7_75t_L g901 ( .A(n_222), .Y(n_901) );
AOI22xp33_ASAP7_75t_L g953 ( .A1(n_222), .A2(n_248), .B1(n_453), .B2(n_841), .Y(n_953) );
NAND2xp5_ASAP7_75t_SL g985 ( .A(n_223), .B(n_386), .Y(n_985) );
AOI22xp5_ASAP7_75t_L g1104 ( .A1(n_224), .A2(n_240), .B1(n_1089), .B2(n_1094), .Y(n_1104) );
INVx1_ASAP7_75t_L g519 ( .A(n_227), .Y(n_519) );
INVx1_ASAP7_75t_L g1156 ( .A(n_228), .Y(n_1156) );
INVxp67_ASAP7_75t_SL g1364 ( .A(n_230), .Y(n_1364) );
INVxp67_ASAP7_75t_SL g1010 ( .A(n_231), .Y(n_1010) );
OAI22xp33_ASAP7_75t_SL g365 ( .A1(n_233), .A2(n_239), .B1(n_366), .B2(n_369), .Y(n_365) );
OAI221xp5_ASAP7_75t_L g407 ( .A1(n_233), .A2(n_239), .B1(n_408), .B2(n_412), .C(n_417), .Y(n_407) );
XNOR2xp5_ASAP7_75t_L g277 ( .A(n_235), .B(n_278), .Y(n_277) );
INVx1_ASAP7_75t_L g1076 ( .A(n_236), .Y(n_1076) );
CKINVDCx5p33_ASAP7_75t_R g981 ( .A(n_242), .Y(n_981) );
OAI211xp5_ASAP7_75t_L g445 ( .A1(n_246), .A2(n_377), .B(n_446), .C(n_454), .Y(n_445) );
INVx1_ASAP7_75t_L g990 ( .A(n_247), .Y(n_990) );
INVx1_ASAP7_75t_L g911 ( .A(n_248), .Y(n_911) );
AOI21xp5_ASAP7_75t_L g249 ( .A1(n_250), .A2(n_270), .B(n_1079), .Y(n_249) );
AND2x2_ASAP7_75t_L g250 ( .A(n_251), .B(n_256), .Y(n_250) );
INVx1_ASAP7_75t_L g1321 ( .A(n_251), .Y(n_1321) );
NOR2xp33_ASAP7_75t_L g251 ( .A(n_252), .B(n_254), .Y(n_251) );
NOR2xp33_ASAP7_75t_L g1324 ( .A(n_252), .B(n_255), .Y(n_1324) );
INVx1_ASAP7_75t_L g1379 ( .A(n_252), .Y(n_1379) );
HB1xp67_ASAP7_75t_L g252 ( .A(n_253), .Y(n_252) );
INVx1_ASAP7_75t_L g254 ( .A(n_255), .Y(n_254) );
NOR2xp33_ASAP7_75t_L g1381 ( .A(n_255), .B(n_1379), .Y(n_1381) );
NAND2xp5_ASAP7_75t_L g256 ( .A(n_257), .B(n_260), .Y(n_256) );
INVx1_ASAP7_75t_L g257 ( .A(n_258), .Y(n_257) );
AND2x4_ASAP7_75t_L g689 ( .A(n_258), .B(n_690), .Y(n_689) );
NOR2xp33_ASAP7_75t_L g1320 ( .A(n_258), .B(n_1321), .Y(n_1320) );
INVx1_ASAP7_75t_L g258 ( .A(n_259), .Y(n_258) );
AND2x4_ASAP7_75t_L g393 ( .A(n_259), .B(n_269), .Y(n_393) );
AND2x4_ASAP7_75t_L g424 ( .A(n_259), .B(n_268), .Y(n_424) );
INVx1_ASAP7_75t_L g685 ( .A(n_260), .Y(n_685) );
AND2x4_ASAP7_75t_SL g1319 ( .A(n_260), .B(n_1320), .Y(n_1319) );
INVx3_ASAP7_75t_L g260 ( .A(n_261), .Y(n_260) );
OR2x6_ASAP7_75t_L g261 ( .A(n_262), .B(n_267), .Y(n_261) );
OR2x6_ASAP7_75t_L g677 ( .A(n_262), .B(n_678), .Y(n_677) );
INVxp67_ASAP7_75t_L g819 ( .A(n_262), .Y(n_819) );
INVx2_ASAP7_75t_L g262 ( .A(n_263), .Y(n_262) );
BUFx4f_ASAP7_75t_L g640 ( .A(n_263), .Y(n_640) );
INVx3_ASAP7_75t_L g654 ( .A(n_263), .Y(n_654) );
INVx3_ASAP7_75t_L g263 ( .A(n_264), .Y(n_263) );
OR2x2_ASAP7_75t_L g264 ( .A(n_265), .B(n_266), .Y(n_264) );
INVx2_ASAP7_75t_L g300 ( .A(n_265), .Y(n_300) );
INVx1_ASAP7_75t_L g313 ( .A(n_265), .Y(n_313) );
INVx2_ASAP7_75t_L g381 ( .A(n_265), .Y(n_381) );
AND2x2_ASAP7_75t_L g387 ( .A(n_265), .B(n_388), .Y(n_387) );
AND2x2_ASAP7_75t_L g391 ( .A(n_265), .B(n_266), .Y(n_391) );
NAND2x1_ASAP7_75t_L g421 ( .A(n_265), .B(n_266), .Y(n_421) );
INVx1_ASAP7_75t_L g301 ( .A(n_266), .Y(n_301) );
AND2x2_ASAP7_75t_L g380 ( .A(n_266), .B(n_381), .Y(n_380) );
INVx2_ASAP7_75t_L g388 ( .A(n_266), .Y(n_388) );
BUFx2_ASAP7_75t_L g415 ( .A(n_266), .Y(n_415) );
NAND2xp5_ASAP7_75t_L g646 ( .A(n_266), .B(n_381), .Y(n_646) );
OR2x2_ASAP7_75t_L g649 ( .A(n_266), .B(n_300), .Y(n_649) );
INVxp67_ASAP7_75t_L g267 ( .A(n_268), .Y(n_267) );
INVx1_ASAP7_75t_L g665 ( .A(n_268), .Y(n_665) );
INVx2_ASAP7_75t_L g268 ( .A(n_269), .Y(n_268) );
BUFx2_ASAP7_75t_L g669 ( .A(n_269), .Y(n_669) );
AND2x4_ASAP7_75t_L g673 ( .A(n_269), .B(n_312), .Y(n_673) );
OAI22xp5_ASAP7_75t_L g270 ( .A1(n_271), .A2(n_272), .B1(n_825), .B2(n_826), .Y(n_270) );
INVx1_ASAP7_75t_L g271 ( .A(n_272), .Y(n_271) );
AOI22xp5_ASAP7_75t_L g272 ( .A1(n_273), .A2(n_595), .B1(n_596), .B2(n_824), .Y(n_272) );
INVx2_ASAP7_75t_L g824 ( .A(n_273), .Y(n_824) );
AOI22x1_ASAP7_75t_L g273 ( .A1(n_274), .A2(n_275), .B1(n_490), .B2(n_594), .Y(n_273) );
INVx1_ASAP7_75t_L g274 ( .A(n_275), .Y(n_274) );
BUFx3_ASAP7_75t_L g275 ( .A(n_276), .Y(n_275) );
AO22x2_ASAP7_75t_L g276 ( .A1(n_277), .A2(n_441), .B1(n_442), .B2(n_489), .Y(n_276) );
INVx1_ASAP7_75t_L g489 ( .A(n_277), .Y(n_489) );
AND4x1_ASAP7_75t_L g278 ( .A(n_279), .B(n_327), .C(n_375), .D(n_435), .Y(n_278) );
AOI21xp5_ASAP7_75t_L g279 ( .A1(n_280), .A2(n_302), .B(n_303), .Y(n_279) );
AOI21xp5_ASAP7_75t_L g485 ( .A1(n_280), .A2(n_486), .B(n_487), .Y(n_485) );
AOI21xp5_ASAP7_75t_L g518 ( .A1(n_280), .A2(n_519), .B(n_520), .Y(n_518) );
AOI21xp33_ASAP7_75t_L g577 ( .A1(n_280), .A2(n_578), .B(n_579), .Y(n_577) );
AOI221xp5_ASAP7_75t_L g728 ( .A1(n_280), .A2(n_729), .B1(n_730), .B2(n_731), .C(n_732), .Y(n_728) );
AOI21xp5_ASAP7_75t_L g789 ( .A1(n_280), .A2(n_790), .B(n_791), .Y(n_789) );
AOI211x1_ASAP7_75t_L g1022 ( .A1(n_280), .A2(n_1023), .B(n_1024), .C(n_1044), .Y(n_1022) );
AOI21xp5_ASAP7_75t_L g1308 ( .A1(n_280), .A2(n_1309), .B(n_1310), .Y(n_1308) );
INVx8_ASAP7_75t_L g280 ( .A(n_281), .Y(n_280) );
AND2x4_ASAP7_75t_L g281 ( .A(n_282), .B(n_294), .Y(n_281) );
INVx1_ASAP7_75t_L g876 ( .A(n_282), .Y(n_876) );
OR2x2_ASAP7_75t_L g282 ( .A(n_283), .B(n_288), .Y(n_282) );
BUFx3_ASAP7_75t_L g1009 ( .A(n_283), .Y(n_1009) );
INVx1_ASAP7_75t_L g1357 ( .A(n_283), .Y(n_1357) );
INVx1_ASAP7_75t_L g283 ( .A(n_284), .Y(n_283) );
BUFx6f_ASAP7_75t_L g362 ( .A(n_284), .Y(n_362) );
INVx1_ASAP7_75t_L g284 ( .A(n_285), .Y(n_284) );
BUFx2_ASAP7_75t_L g346 ( .A(n_285), .Y(n_346) );
NAND2xp5_ASAP7_75t_L g285 ( .A(n_286), .B(n_287), .Y(n_285) );
BUFx6f_ASAP7_75t_L g309 ( .A(n_286), .Y(n_309) );
INVx2_ASAP7_75t_L g318 ( .A(n_286), .Y(n_318) );
AND2x4_ASAP7_75t_L g331 ( .A(n_286), .B(n_332), .Y(n_331) );
OR2x2_ASAP7_75t_L g548 ( .A(n_286), .B(n_320), .Y(n_548) );
INVx1_ASAP7_75t_L g308 ( .A(n_287), .Y(n_308) );
INVx2_ASAP7_75t_L g332 ( .A(n_287), .Y(n_332) );
OR2x2_ASAP7_75t_L g305 ( .A(n_288), .B(n_306), .Y(n_305) );
INVx1_ASAP7_75t_L g438 ( .A(n_288), .Y(n_438) );
INVx1_ASAP7_75t_L g550 ( .A(n_288), .Y(n_550) );
OR2x2_ASAP7_75t_L g288 ( .A(n_289), .B(n_292), .Y(n_288) );
OR2x2_ASAP7_75t_L g336 ( .A(n_289), .B(n_337), .Y(n_336) );
INVx1_ASAP7_75t_L g660 ( .A(n_289), .Y(n_660) );
HB1xp67_ASAP7_75t_L g723 ( .A(n_289), .Y(n_723) );
AND2x2_ASAP7_75t_SL g949 ( .A(n_289), .B(n_393), .Y(n_949) );
INVx2_ASAP7_75t_L g289 ( .A(n_290), .Y(n_289) );
BUFx2_ASAP7_75t_L g314 ( .A(n_290), .Y(n_314) );
INVx1_ASAP7_75t_L g290 ( .A(n_291), .Y(n_290) );
INVx1_ASAP7_75t_L g897 ( .A(n_292), .Y(n_897) );
INVx3_ASAP7_75t_L g323 ( .A(n_293), .Y(n_323) );
NAND2xp33_ASAP7_75t_SL g337 ( .A(n_293), .B(n_325), .Y(n_337) );
BUFx3_ASAP7_75t_L g529 ( .A(n_293), .Y(n_529) );
NAND2xp5_ASAP7_75t_L g965 ( .A(n_294), .B(n_966), .Y(n_965) );
OR2x2_ASAP7_75t_L g294 ( .A(n_295), .B(n_297), .Y(n_294) );
AND2x4_ASAP7_75t_L g333 ( .A(n_295), .B(n_322), .Y(n_333) );
INVx1_ASAP7_75t_L g295 ( .A(n_296), .Y(n_295) );
INVx1_ASAP7_75t_L g355 ( .A(n_296), .Y(n_355) );
NAND2xp5_ASAP7_75t_L g946 ( .A(n_296), .B(n_382), .Y(n_946) );
NAND2xp5_ASAP7_75t_L g297 ( .A(n_298), .B(n_299), .Y(n_297) );
NAND2xp5_ASAP7_75t_L g311 ( .A(n_298), .B(n_312), .Y(n_311) );
AND2x6_ASAP7_75t_L g399 ( .A(n_298), .B(n_390), .Y(n_399) );
INVx1_ASAP7_75t_L g416 ( .A(n_298), .Y(n_416) );
AND2x2_ASAP7_75t_L g496 ( .A(n_298), .B(n_497), .Y(n_496) );
NAND2xp5_ASAP7_75t_L g941 ( .A(n_298), .B(n_434), .Y(n_941) );
BUFx6f_ASAP7_75t_L g397 ( .A(n_299), .Y(n_397) );
AND2x2_ASAP7_75t_L g403 ( .A(n_299), .B(n_382), .Y(n_403) );
INVx3_ASAP7_75t_L g427 ( .A(n_299), .Y(n_427) );
AND2x2_ASAP7_75t_L g299 ( .A(n_300), .B(n_301), .Y(n_299) );
HB1xp67_ASAP7_75t_L g849 ( .A(n_300), .Y(n_849) );
AND2x4_ASAP7_75t_L g304 ( .A(n_305), .B(n_310), .Y(n_304) );
AND2x4_ASAP7_75t_L g792 ( .A(n_305), .B(n_310), .Y(n_792) );
INVx2_ASAP7_75t_L g874 ( .A(n_305), .Y(n_874) );
INVx3_ASAP7_75t_L g610 ( .A(n_306), .Y(n_610) );
INVx4_ASAP7_75t_L g1362 ( .A(n_306), .Y(n_1362) );
BUFx6f_ASAP7_75t_L g306 ( .A(n_307), .Y(n_306) );
BUFx3_ASAP7_75t_L g623 ( .A(n_307), .Y(n_623) );
BUFx2_ASAP7_75t_L g903 ( .A(n_307), .Y(n_903) );
NAND2x1p5_ASAP7_75t_L g307 ( .A(n_308), .B(n_309), .Y(n_307) );
BUFx2_ASAP7_75t_L g711 ( .A(n_308), .Y(n_711) );
INVx2_ASAP7_75t_L g368 ( .A(n_309), .Y(n_368) );
AND2x4_ASAP7_75t_L g536 ( .A(n_309), .B(n_374), .Y(n_536) );
BUFx2_ASAP7_75t_L g708 ( .A(n_309), .Y(n_708) );
OR2x2_ASAP7_75t_L g310 ( .A(n_311), .B(n_314), .Y(n_310) );
OR2x2_ASAP7_75t_L g936 ( .A(n_311), .B(n_314), .Y(n_936) );
INVx1_ASAP7_75t_L g312 ( .A(n_313), .Y(n_312) );
INVxp67_ASAP7_75t_L g326 ( .A(n_314), .Y(n_326) );
INVx1_ASAP7_75t_L g690 ( .A(n_314), .Y(n_690) );
INVx1_ASAP7_75t_L g870 ( .A(n_314), .Y(n_870) );
NAND2xp5_ASAP7_75t_L g959 ( .A(n_315), .B(n_960), .Y(n_959) );
OR2x2_ASAP7_75t_L g315 ( .A(n_316), .B(n_326), .Y(n_315) );
OR2x6_ASAP7_75t_L g521 ( .A(n_316), .B(n_326), .Y(n_521) );
NAND2x1p5_ASAP7_75t_L g316 ( .A(n_317), .B(n_322), .Y(n_316) );
INVx8_ASAP7_75t_L g350 ( .A(n_317), .Y(n_350) );
BUFx3_ASAP7_75t_L g532 ( .A(n_317), .Y(n_532) );
BUFx3_ASAP7_75t_L g916 ( .A(n_317), .Y(n_916) );
HB1xp67_ASAP7_75t_L g1012 ( .A(n_317), .Y(n_1012) );
AND2x4_ASAP7_75t_L g317 ( .A(n_318), .B(n_319), .Y(n_317) );
AND2x4_ASAP7_75t_L g340 ( .A(n_318), .B(n_341), .Y(n_340) );
INVx1_ASAP7_75t_L g319 ( .A(n_320), .Y(n_319) );
INVx1_ASAP7_75t_L g320 ( .A(n_321), .Y(n_320) );
INVxp67_ASAP7_75t_L g341 ( .A(n_321), .Y(n_341) );
INVx1_ASAP7_75t_L g918 ( .A(n_322), .Y(n_918) );
AND2x6_ASAP7_75t_L g925 ( .A(n_322), .B(n_367), .Y(n_925) );
AND2x2_ASAP7_75t_L g927 ( .A(n_322), .B(n_373), .Y(n_927) );
AND2x4_ASAP7_75t_L g322 ( .A(n_323), .B(n_324), .Y(n_322) );
NAND3x1_ASAP7_75t_L g354 ( .A(n_323), .B(n_355), .C(n_356), .Y(n_354) );
NAND2x1p5_ASAP7_75t_L g541 ( .A(n_323), .B(n_356), .Y(n_541) );
OR2x4_ASAP7_75t_L g695 ( .A(n_323), .B(n_548), .Y(n_695) );
INVx1_ASAP7_75t_L g698 ( .A(n_323), .Y(n_698) );
AND2x4_ASAP7_75t_L g703 ( .A(n_323), .B(n_331), .Y(n_703) );
OR2x6_ASAP7_75t_L g718 ( .A(n_323), .B(n_346), .Y(n_718) );
INVx1_ASAP7_75t_L g324 ( .A(n_325), .Y(n_324) );
AND3x4_ASAP7_75t_L g528 ( .A(n_325), .B(n_469), .C(n_529), .Y(n_528) );
HB1xp67_ASAP7_75t_L g721 ( .A(n_325), .Y(n_721) );
AND2x2_ASAP7_75t_L g907 ( .A(n_325), .B(n_529), .Y(n_907) );
NOR3xp33_ASAP7_75t_L g327 ( .A(n_328), .B(n_334), .C(n_365), .Y(n_327) );
NOR3xp33_ASAP7_75t_L g580 ( .A(n_328), .B(n_581), .C(n_592), .Y(n_580) );
NOR3xp33_ASAP7_75t_L g770 ( .A(n_328), .B(n_771), .C(n_787), .Y(n_770) );
HB1xp67_ASAP7_75t_L g328 ( .A(n_329), .Y(n_328) );
NOR3xp33_ASAP7_75t_L g470 ( .A(n_329), .B(n_471), .C(n_484), .Y(n_470) );
NOR3xp33_ASAP7_75t_L g522 ( .A(n_329), .B(n_523), .C(n_544), .Y(n_522) );
INVx3_ASAP7_75t_L g745 ( .A(n_329), .Y(n_745) );
AOI221xp5_ASAP7_75t_L g864 ( .A1(n_329), .A2(n_370), .B1(n_525), .B2(n_847), .C(n_865), .Y(n_864) );
INVx3_ASAP7_75t_L g1032 ( .A(n_329), .Y(n_1032) );
AOI221xp5_ASAP7_75t_L g1311 ( .A1(n_329), .A2(n_525), .B1(n_776), .B2(n_1280), .C(n_1312), .Y(n_1311) );
AND2x4_ASAP7_75t_L g329 ( .A(n_330), .B(n_333), .Y(n_329) );
BUFx2_ASAP7_75t_L g780 ( .A(n_330), .Y(n_780) );
BUFx2_ASAP7_75t_L g330 ( .A(n_331), .Y(n_330) );
BUFx2_ASAP7_75t_L g351 ( .A(n_331), .Y(n_351) );
INVx2_ASAP7_75t_L g483 ( .A(n_331), .Y(n_483) );
BUFx2_ASAP7_75t_L g538 ( .A(n_331), .Y(n_538) );
BUFx3_ASAP7_75t_L g1006 ( .A(n_331), .Y(n_1006) );
INVx1_ASAP7_75t_L g374 ( .A(n_332), .Y(n_374) );
NAND2x1_ASAP7_75t_L g366 ( .A(n_333), .B(n_367), .Y(n_366) );
AND2x4_ASAP7_75t_SL g370 ( .A(n_333), .B(n_371), .Y(n_370) );
AND2x4_ASAP7_75t_SL g525 ( .A(n_333), .B(n_367), .Y(n_525) );
AND2x2_ASAP7_75t_L g774 ( .A(n_333), .B(n_367), .Y(n_774) );
AND2x4_ASAP7_75t_L g776 ( .A(n_333), .B(n_371), .Y(n_776) );
OAI22xp5_ASAP7_75t_SL g334 ( .A1(n_335), .A2(n_338), .B1(n_352), .B2(n_357), .Y(n_334) );
BUFx3_ASAP7_75t_L g603 ( .A(n_335), .Y(n_603) );
BUFx4f_ASAP7_75t_L g335 ( .A(n_336), .Y(n_335) );
BUFx8_ASAP7_75t_L g472 ( .A(n_336), .Y(n_472) );
BUFx2_ASAP7_75t_L g1000 ( .A(n_336), .Y(n_1000) );
OAI221xp5_ASAP7_75t_L g338 ( .A1(n_339), .A2(n_342), .B1(n_343), .B2(n_347), .C(n_348), .Y(n_338) );
INVx3_ASAP7_75t_L g534 ( .A(n_339), .Y(n_534) );
BUFx2_ASAP7_75t_L g783 ( .A(n_339), .Y(n_783) );
OR2x6_ASAP7_75t_SL g895 ( .A(n_339), .B(n_896), .Y(n_895) );
INVx2_ASAP7_75t_L g339 ( .A(n_340), .Y(n_339) );
BUFx6f_ASAP7_75t_L g359 ( .A(n_340), .Y(n_359) );
BUFx8_ASAP7_75t_L g440 ( .A(n_340), .Y(n_440) );
BUFx6f_ASAP7_75t_L g620 ( .A(n_340), .Y(n_620) );
OAI221xp5_ASAP7_75t_L g473 ( .A1(n_343), .A2(n_474), .B1(n_475), .B2(n_476), .C(n_477), .Y(n_473) );
INVx3_ASAP7_75t_L g343 ( .A(n_344), .Y(n_343) );
BUFx2_ASAP7_75t_L g344 ( .A(n_345), .Y(n_344) );
INVx1_ASAP7_75t_L g345 ( .A(n_346), .Y(n_345) );
INVx8_ASAP7_75t_L g349 ( .A(n_350), .Y(n_349) );
INVx2_ASAP7_75t_L g437 ( .A(n_350), .Y(n_437) );
INVx3_ASAP7_75t_L g591 ( .A(n_350), .Y(n_591) );
INVx2_ASAP7_75t_L g738 ( .A(n_350), .Y(n_738) );
INVx2_ASAP7_75t_L g352 ( .A(n_353), .Y(n_352) );
CKINVDCx5p33_ASAP7_75t_R g478 ( .A(n_353), .Y(n_478) );
INVx2_ASAP7_75t_L g1007 ( .A(n_353), .Y(n_1007) );
INVx3_ASAP7_75t_L g353 ( .A(n_354), .Y(n_353) );
INVx3_ASAP7_75t_L g627 ( .A(n_354), .Y(n_627) );
OAI221xp5_ASAP7_75t_L g357 ( .A1(n_358), .A2(n_360), .B1(n_361), .B2(n_363), .C(n_364), .Y(n_357) );
INVx2_ASAP7_75t_L g358 ( .A(n_359), .Y(n_358) );
INVx2_ASAP7_75t_L g613 ( .A(n_359), .Y(n_613) );
AND2x4_ASAP7_75t_L g697 ( .A(n_359), .B(n_698), .Y(n_697) );
BUFx6f_ASAP7_75t_L g741 ( .A(n_359), .Y(n_741) );
BUFx6f_ASAP7_75t_L g860 ( .A(n_359), .Y(n_860) );
OAI211xp5_ASAP7_75t_L g417 ( .A1(n_360), .A2(n_418), .B(n_422), .C(n_425), .Y(n_417) );
OAI221xp5_ASAP7_75t_L g479 ( .A1(n_361), .A2(n_460), .B1(n_474), .B2(n_480), .C(n_481), .Y(n_479) );
OAI22xp5_ASAP7_75t_L g1290 ( .A1(n_361), .A2(n_1291), .B1(n_1292), .B2(n_1293), .Y(n_1290) );
CKINVDCx8_ASAP7_75t_R g361 ( .A(n_362), .Y(n_361) );
INVx3_ASAP7_75t_L g615 ( .A(n_362), .Y(n_615) );
INVx3_ASAP7_75t_L g630 ( .A(n_362), .Y(n_630) );
INVx3_ASAP7_75t_L g1003 ( .A(n_362), .Y(n_1003) );
INVx1_ASAP7_75t_L g1303 ( .A(n_362), .Y(n_1303) );
INVx2_ASAP7_75t_L g998 ( .A(n_366), .Y(n_998) );
INVx3_ASAP7_75t_L g367 ( .A(n_368), .Y(n_367) );
INVx1_ASAP7_75t_L g369 ( .A(n_370), .Y(n_369) );
AOI22xp33_ASAP7_75t_L g524 ( .A1(n_370), .A2(n_498), .B1(n_525), .B2(n_526), .Y(n_524) );
AOI22xp33_ASAP7_75t_L g582 ( .A1(n_370), .A2(n_525), .B1(n_560), .B2(n_583), .Y(n_582) );
AOI22xp5_ASAP7_75t_L g733 ( .A1(n_370), .A2(n_525), .B1(n_734), .B2(n_735), .Y(n_733) );
INVx2_ASAP7_75t_L g371 ( .A(n_372), .Y(n_371) );
INVx1_ASAP7_75t_L g372 ( .A(n_373), .Y(n_372) );
INVx1_ASAP7_75t_L g373 ( .A(n_374), .Y(n_373) );
OAI21xp5_ASAP7_75t_L g375 ( .A1(n_376), .A2(n_407), .B(n_430), .Y(n_375) );
INVx2_ASAP7_75t_SL g377 ( .A(n_378), .Y(n_377) );
INVx3_ASAP7_75t_L g506 ( .A(n_378), .Y(n_506) );
NAND2xp5_ASAP7_75t_R g1059 ( .A(n_378), .B(n_1031), .Y(n_1059) );
AOI22xp33_ASAP7_75t_L g1286 ( .A1(n_378), .A2(n_405), .B1(n_1287), .B2(n_1288), .Y(n_1286) );
AND2x4_ASAP7_75t_L g378 ( .A(n_379), .B(n_382), .Y(n_378) );
BUFx2_ASAP7_75t_L g1337 ( .A(n_379), .Y(n_1337) );
BUFx6f_ASAP7_75t_L g379 ( .A(n_380), .Y(n_379) );
BUFx3_ASAP7_75t_L g398 ( .A(n_380), .Y(n_398) );
INVx2_ASAP7_75t_L g429 ( .A(n_380), .Y(n_429) );
BUFx3_ASAP7_75t_L g453 ( .A(n_380), .Y(n_453) );
AND2x4_ASAP7_75t_L g405 ( .A(n_382), .B(n_406), .Y(n_405) );
AND2x4_ASAP7_75t_SL g411 ( .A(n_382), .B(n_390), .Y(n_411) );
AND2x2_ASAP7_75t_L g752 ( .A(n_382), .B(n_753), .Y(n_752) );
BUFx2_ASAP7_75t_L g852 ( .A(n_382), .Y(n_852) );
AND2x2_ASAP7_75t_L g871 ( .A(n_382), .B(n_406), .Y(n_871) );
HB1xp67_ASAP7_75t_L g678 ( .A(n_383), .Y(n_678) );
AOI21xp5_ASAP7_75t_L g384 ( .A1(n_385), .A2(n_394), .B(n_399), .Y(n_384) );
HB1xp67_ASAP7_75t_L g509 ( .A(n_386), .Y(n_509) );
INVx1_ASAP7_75t_L g571 ( .A(n_386), .Y(n_571) );
BUFx3_ASAP7_75t_L g386 ( .A(n_387), .Y(n_386) );
BUFx6f_ASAP7_75t_L g406 ( .A(n_387), .Y(n_406) );
AND2x4_ASAP7_75t_L g687 ( .A(n_387), .B(n_678), .Y(n_687) );
INVx2_ASAP7_75t_L g816 ( .A(n_387), .Y(n_816) );
BUFx2_ASAP7_75t_L g797 ( .A(n_389), .Y(n_797) );
BUFx6f_ASAP7_75t_L g389 ( .A(n_390), .Y(n_389) );
BUFx3_ASAP7_75t_L g448 ( .A(n_390), .Y(n_448) );
AND2x2_ASAP7_75t_L g664 ( .A(n_390), .B(n_665), .Y(n_664) );
BUFx3_ASAP7_75t_L g988 ( .A(n_390), .Y(n_988) );
INVx1_ASAP7_75t_L g1335 ( .A(n_390), .Y(n_1335) );
BUFx6f_ASAP7_75t_L g390 ( .A(n_391), .Y(n_390) );
INVx1_ASAP7_75t_L g813 ( .A(n_391), .Y(n_813) );
INVx4_ASAP7_75t_L g392 ( .A(n_393), .Y(n_392) );
INVx1_ASAP7_75t_SL g572 ( .A(n_393), .Y(n_572) );
NAND2xp5_ASAP7_75t_L g658 ( .A(n_393), .B(n_659), .Y(n_658) );
INVx4_ASAP7_75t_L g757 ( .A(n_393), .Y(n_757) );
NAND4xp25_ASAP7_75t_L g984 ( .A(n_393), .B(n_985), .C(n_986), .D(n_987), .Y(n_984) );
INVx2_ASAP7_75t_SL g395 ( .A(n_396), .Y(n_395) );
INVx2_ASAP7_75t_L g511 ( .A(n_396), .Y(n_511) );
INVx3_ASAP7_75t_L g396 ( .A(n_397), .Y(n_396) );
BUFx3_ASAP7_75t_L g801 ( .A(n_398), .Y(n_801) );
INVx1_ASAP7_75t_SL g1058 ( .A(n_398), .Y(n_1058) );
AOI21xp5_ASAP7_75t_L g446 ( .A1(n_399), .A2(n_447), .B(n_451), .Y(n_446) );
AOI21xp5_ASAP7_75t_L g507 ( .A1(n_399), .A2(n_508), .B(n_510), .Y(n_507) );
AOI21xp5_ASAP7_75t_L g568 ( .A1(n_399), .A2(n_569), .B(n_573), .Y(n_568) );
AOI221xp5_ASAP7_75t_L g751 ( .A1(n_399), .A2(n_730), .B1(n_752), .B2(n_754), .C(n_758), .Y(n_751) );
AOI21xp5_ASAP7_75t_L g795 ( .A1(n_399), .A2(n_796), .B(n_800), .Y(n_795) );
AOI21xp5_ASAP7_75t_L g1051 ( .A1(n_399), .A2(n_1052), .B(n_1055), .Y(n_1051) );
AOI221xp5_ASAP7_75t_L g1277 ( .A1(n_399), .A2(n_760), .B1(n_1278), .B2(n_1279), .C(n_1280), .Y(n_1277) );
INVx1_ASAP7_75t_L g1338 ( .A(n_399), .Y(n_1338) );
AOI22xp33_ASAP7_75t_L g400 ( .A1(n_401), .A2(n_402), .B1(n_404), .B2(n_405), .Y(n_400) );
AOI22xp33_ASAP7_75t_L g435 ( .A1(n_401), .A2(n_404), .B1(n_436), .B2(n_439), .Y(n_435) );
AOI22xp33_ASAP7_75t_L g574 ( .A1(n_402), .A2(n_517), .B1(n_575), .B2(n_576), .Y(n_574) );
AOI22xp5_ASAP7_75t_L g748 ( .A1(n_402), .A2(n_405), .B1(n_749), .B2(n_750), .Y(n_748) );
AOI221xp5_ASAP7_75t_SL g1281 ( .A1(n_402), .A2(n_1282), .B1(n_1283), .B2(n_1284), .C(n_1285), .Y(n_1281) );
NAND2xp5_ASAP7_75t_L g1347 ( .A(n_402), .B(n_1348), .Y(n_1347) );
BUFx6f_ASAP7_75t_L g402 ( .A(n_403), .Y(n_402) );
AOI22xp33_ASAP7_75t_L g454 ( .A1(n_403), .A2(n_405), .B1(n_455), .B2(n_456), .Y(n_454) );
INVx1_ASAP7_75t_L g515 ( .A(n_403), .Y(n_515) );
AND2x4_ASAP7_75t_L g891 ( .A(n_403), .B(n_870), .Y(n_891) );
BUFx6f_ASAP7_75t_L g517 ( .A(n_405), .Y(n_517) );
INVx1_ASAP7_75t_L g806 ( .A(n_405), .Y(n_806) );
AOI22xp33_ASAP7_75t_L g1050 ( .A1(n_405), .A2(n_514), .B1(n_1046), .B2(n_1047), .Y(n_1050) );
AOI22xp33_ASAP7_75t_L g1344 ( .A1(n_405), .A2(n_752), .B1(n_1345), .B2(n_1346), .Y(n_1344) );
INVx1_ASAP7_75t_L g450 ( .A(n_406), .Y(n_450) );
BUFx6f_ASAP7_75t_L g564 ( .A(n_406), .Y(n_564) );
INVx2_ASAP7_75t_L g756 ( .A(n_406), .Y(n_756) );
INVx2_ASAP7_75t_L g408 ( .A(n_409), .Y(n_408) );
INVx2_ASAP7_75t_L g458 ( .A(n_409), .Y(n_458) );
AOI22xp33_ASAP7_75t_L g820 ( .A1(n_409), .A2(n_413), .B1(n_773), .B2(n_775), .Y(n_820) );
INVx1_ASAP7_75t_L g1061 ( .A(n_409), .Y(n_1061) );
INVx4_ASAP7_75t_L g409 ( .A(n_410), .Y(n_409) );
INVx2_ASAP7_75t_L g410 ( .A(n_411), .Y(n_410) );
BUFx3_ASAP7_75t_L g760 ( .A(n_411), .Y(n_760) );
BUFx2_ASAP7_75t_L g1075 ( .A(n_412), .Y(n_1075) );
INVx2_ASAP7_75t_L g412 ( .A(n_413), .Y(n_412) );
NOR2x1_ASAP7_75t_L g413 ( .A(n_414), .B(n_416), .Y(n_413) );
INVx1_ASAP7_75t_L g414 ( .A(n_415), .Y(n_414) );
BUFx2_ASAP7_75t_L g497 ( .A(n_415), .Y(n_497) );
AND2x4_ASAP7_75t_L g668 ( .A(n_415), .B(n_669), .Y(n_668) );
INVx1_ASAP7_75t_L g943 ( .A(n_415), .Y(n_943) );
INVx1_ASAP7_75t_L g851 ( .A(n_416), .Y(n_851) );
INVx1_ASAP7_75t_L g418 ( .A(n_419), .Y(n_418) );
INVx2_ASAP7_75t_L g845 ( .A(n_419), .Y(n_845) );
INVx2_ASAP7_75t_L g979 ( .A(n_419), .Y(n_979) );
INVx4_ASAP7_75t_L g419 ( .A(n_420), .Y(n_419) );
BUFx4f_ASAP7_75t_L g501 ( .A(n_420), .Y(n_501) );
OR2x6_ASAP7_75t_L g955 ( .A(n_420), .B(n_956), .Y(n_955) );
BUFx4f_ASAP7_75t_L g1063 ( .A(n_420), .Y(n_1063) );
BUFx6f_ASAP7_75t_L g420 ( .A(n_421), .Y(n_420) );
BUFx3_ASAP7_75t_L g463 ( .A(n_421), .Y(n_463) );
INVx2_ASAP7_75t_L g423 ( .A(n_424), .Y(n_423) );
INVx1_ASAP7_75t_L g465 ( .A(n_424), .Y(n_465) );
INVx3_ASAP7_75t_L g565 ( .A(n_424), .Y(n_565) );
INVx2_ASAP7_75t_L g817 ( .A(n_424), .Y(n_817) );
OAI221xp5_ASAP7_75t_L g1062 ( .A1(n_424), .A2(n_1063), .B1(n_1064), .B2(n_1065), .C(n_1068), .Y(n_1062) );
INVx2_ASAP7_75t_SL g426 ( .A(n_427), .Y(n_426) );
INVx2_ASAP7_75t_L g452 ( .A(n_427), .Y(n_452) );
INVx1_ASAP7_75t_L g504 ( .A(n_427), .Y(n_504) );
INVx1_ASAP7_75t_L g762 ( .A(n_427), .Y(n_762) );
INVx2_ASAP7_75t_L g841 ( .A(n_427), .Y(n_841) );
INVx2_ASAP7_75t_L g1056 ( .A(n_427), .Y(n_1056) );
INVx1_ASAP7_75t_L g428 ( .A(n_429), .Y(n_428) );
INVx3_ASAP7_75t_L g753 ( .A(n_429), .Y(n_753) );
OAI21xp5_ASAP7_75t_SL g493 ( .A1(n_430), .A2(n_494), .B(n_505), .Y(n_493) );
OAI21xp5_ASAP7_75t_SL g557 ( .A1(n_430), .A2(n_558), .B(n_567), .Y(n_557) );
AOI21xp5_ASAP7_75t_L g746 ( .A1(n_430), .A2(n_747), .B(n_764), .Y(n_746) );
OAI21xp5_ASAP7_75t_L g1048 ( .A1(n_430), .A2(n_1049), .B(n_1060), .Y(n_1048) );
OAI21xp5_ASAP7_75t_L g1330 ( .A1(n_430), .A2(n_1331), .B(n_1339), .Y(n_1330) );
INVx2_ASAP7_75t_L g430 ( .A(n_431), .Y(n_430) );
BUFx2_ASAP7_75t_L g431 ( .A(n_432), .Y(n_431) );
NAND2xp5_ASAP7_75t_L g966 ( .A(n_432), .B(n_967), .Y(n_966) );
INVx1_ASAP7_75t_L g432 ( .A(n_433), .Y(n_432) );
OR2x6_ASAP7_75t_L g540 ( .A(n_433), .B(n_541), .Y(n_540) );
AND2x4_ASAP7_75t_L g634 ( .A(n_433), .B(n_635), .Y(n_634) );
OR2x2_ASAP7_75t_L g739 ( .A(n_433), .B(n_541), .Y(n_739) );
BUFx2_ASAP7_75t_L g433 ( .A(n_434), .Y(n_433) );
INVx2_ASAP7_75t_L g469 ( .A(n_434), .Y(n_469) );
AOI22xp33_ASAP7_75t_L g488 ( .A1(n_436), .A2(n_439), .B1(n_455), .B2(n_456), .Y(n_488) );
AOI22xp33_ASAP7_75t_L g1045 ( .A1(n_436), .A2(n_439), .B1(n_1046), .B2(n_1047), .Y(n_1045) );
NAND2xp5_ASAP7_75t_L g1314 ( .A(n_436), .B(n_1284), .Y(n_1314) );
AND2x4_ASAP7_75t_L g436 ( .A(n_437), .B(n_438), .Y(n_436) );
AND2x4_ASAP7_75t_L g766 ( .A(n_437), .B(n_438), .Y(n_766) );
AOI22xp5_ASAP7_75t_L g920 ( .A1(n_437), .A2(n_862), .B1(n_890), .B2(n_921), .Y(n_920) );
AND2x4_ASAP7_75t_L g439 ( .A(n_438), .B(n_440), .Y(n_439) );
INVx2_ASAP7_75t_L g788 ( .A(n_439), .Y(n_788) );
NAND2xp5_ASAP7_75t_L g1376 ( .A(n_439), .B(n_1345), .Y(n_1376) );
INVx2_ASAP7_75t_SL g474 ( .A(n_440), .Y(n_474) );
INVx3_ASAP7_75t_L g1354 ( .A(n_440), .Y(n_1354) );
INVx1_ASAP7_75t_L g441 ( .A(n_442), .Y(n_441) );
AND4x1_ASAP7_75t_L g443 ( .A(n_444), .B(n_470), .C(n_485), .D(n_488), .Y(n_443) );
OAI21xp5_ASAP7_75t_L g444 ( .A1(n_445), .A2(n_457), .B(n_467), .Y(n_444) );
INVx2_ASAP7_75t_SL g449 ( .A(n_450), .Y(n_449) );
OAI211xp5_ASAP7_75t_L g459 ( .A1(n_460), .A2(n_461), .B(n_464), .C(n_466), .Y(n_459) );
OAI22xp5_ASAP7_75t_L g647 ( .A1(n_461), .A2(n_612), .B1(n_621), .B2(n_648), .Y(n_647) );
OAI211xp5_ASAP7_75t_L g989 ( .A1(n_461), .A2(n_990), .B(n_991), .C(n_992), .Y(n_989) );
INVx5_ASAP7_75t_L g461 ( .A(n_462), .Y(n_461) );
INVx2_ASAP7_75t_SL g462 ( .A(n_463), .Y(n_462) );
BUFx2_ASAP7_75t_SL g655 ( .A(n_463), .Y(n_655) );
OR2x2_ASAP7_75t_L g945 ( .A(n_463), .B(n_946), .Y(n_945) );
AOI221xp5_ASAP7_75t_L g1273 ( .A1(n_467), .A2(n_1274), .B1(n_1275), .B2(n_1276), .C(n_1289), .Y(n_1273) );
BUFx2_ASAP7_75t_L g467 ( .A(n_468), .Y(n_467) );
BUFx2_ASAP7_75t_L g823 ( .A(n_468), .Y(n_823) );
AOI21x1_ASAP7_75t_L g833 ( .A1(n_468), .A2(n_834), .B(n_854), .Y(n_833) );
INVx1_ASAP7_75t_L g468 ( .A(n_469), .Y(n_468) );
OAI31xp33_ASAP7_75t_L g893 ( .A1(n_469), .A2(n_894), .A3(n_898), .B(n_919), .Y(n_893) );
OAI22xp5_ASAP7_75t_SL g471 ( .A1(n_472), .A2(n_473), .B1(n_478), .B2(n_479), .Y(n_471) );
INVx2_ASAP7_75t_L g482 ( .A(n_483), .Y(n_482) );
INVx2_ASAP7_75t_L g862 ( .A(n_483), .Y(n_862) );
INVx1_ASAP7_75t_L g594 ( .A(n_490), .Y(n_594) );
XNOR2xp5_ASAP7_75t_L g490 ( .A(n_491), .B(n_555), .Y(n_490) );
INVx1_ASAP7_75t_L g554 ( .A(n_492), .Y(n_554) );
NAND3xp33_ASAP7_75t_L g492 ( .A(n_493), .B(n_518), .C(n_522), .Y(n_492) );
NAND2xp5_ASAP7_75t_L g495 ( .A(n_496), .B(n_498), .Y(n_495) );
NAND2xp5_ASAP7_75t_L g559 ( .A(n_496), .B(n_560), .Y(n_559) );
AOI222xp33_ASAP7_75t_L g759 ( .A1(n_496), .A2(n_734), .B1(n_735), .B2(n_760), .C1(n_761), .C2(n_763), .Y(n_759) );
AOI22xp33_ASAP7_75t_L g1340 ( .A1(n_496), .A2(n_1341), .B1(n_1342), .B2(n_1343), .Y(n_1340) );
AOI22xp5_ASAP7_75t_L g846 ( .A1(n_497), .A2(n_847), .B1(n_848), .B2(n_850), .Y(n_846) );
AOI22xp33_ASAP7_75t_L g980 ( .A1(n_497), .A2(n_848), .B1(n_981), .B2(n_982), .Y(n_980) );
OAI211xp5_ASAP7_75t_L g499 ( .A1(n_500), .A2(n_501), .B(n_502), .C(n_503), .Y(n_499) );
OAI211xp5_ASAP7_75t_L g561 ( .A1(n_501), .A2(n_562), .B(n_563), .C(n_566), .Y(n_561) );
AOI22xp33_ASAP7_75t_L g512 ( .A1(n_513), .A2(n_514), .B1(n_516), .B2(n_517), .Y(n_512) );
AOI22xp33_ASAP7_75t_L g802 ( .A1(n_514), .A2(n_803), .B1(n_804), .B2(n_805), .Y(n_802) );
INVx2_ASAP7_75t_L g514 ( .A(n_515), .Y(n_514) );
INVx3_ASAP7_75t_L g729 ( .A(n_521), .Y(n_729) );
INVx5_ASAP7_75t_L g1019 ( .A(n_521), .Y(n_1019) );
NAND2xp5_ASAP7_75t_L g523 ( .A(n_524), .B(n_527), .Y(n_523) );
AOI33xp33_ASAP7_75t_L g527 ( .A1(n_528), .A2(n_530), .A3(n_533), .B1(n_537), .B2(n_539), .B3(n_542), .Y(n_527) );
AOI33xp33_ASAP7_75t_L g584 ( .A1(n_528), .A2(n_539), .A3(n_585), .B1(n_588), .B2(n_589), .B3(n_590), .Y(n_584) );
INVx1_ASAP7_75t_L g743 ( .A(n_528), .Y(n_743) );
BUFx3_ASAP7_75t_L g778 ( .A(n_528), .Y(n_778) );
AOI33xp33_ASAP7_75t_L g856 ( .A1(n_528), .A2(n_857), .A3(n_858), .B1(n_859), .B2(n_861), .B3(n_863), .Y(n_856) );
INVx3_ASAP7_75t_L g707 ( .A(n_529), .Y(n_707) );
BUFx3_ASAP7_75t_L g531 ( .A(n_532), .Y(n_531) );
INVx2_ASAP7_75t_SL g587 ( .A(n_532), .Y(n_587) );
AND2x2_ASAP7_75t_L g552 ( .A(n_534), .B(n_550), .Y(n_552) );
BUFx2_ASAP7_75t_L g1039 ( .A(n_535), .Y(n_1039) );
BUFx12f_ASAP7_75t_L g535 ( .A(n_536), .Y(n_535) );
BUFx3_ASAP7_75t_L g543 ( .A(n_536), .Y(n_543) );
AND2x4_ASAP7_75t_L g967 ( .A(n_536), .B(n_897), .Y(n_967) );
INVx5_ASAP7_75t_L g1037 ( .A(n_536), .Y(n_1037) );
INVx1_ASAP7_75t_L g1043 ( .A(n_538), .Y(n_1043) );
INVx1_ASAP7_75t_SL g539 ( .A(n_540), .Y(n_539) );
INVx1_ASAP7_75t_L g863 ( .A(n_540), .Y(n_863) );
NAND2xp5_ASAP7_75t_L g1015 ( .A(n_545), .B(n_1016), .Y(n_1015) );
OR2x6_ASAP7_75t_L g545 ( .A(n_546), .B(n_549), .Y(n_545) );
OR2x2_ASAP7_75t_L g593 ( .A(n_546), .B(n_549), .Y(n_593) );
INVx2_ASAP7_75t_SL g546 ( .A(n_547), .Y(n_546) );
INVx2_ASAP7_75t_L g547 ( .A(n_548), .Y(n_547) );
BUFx4f_ASAP7_75t_L g607 ( .A(n_548), .Y(n_607) );
OR2x4_ASAP7_75t_L g716 ( .A(n_548), .B(n_698), .Y(n_716) );
BUFx3_ASAP7_75t_L g1298 ( .A(n_548), .Y(n_1298) );
BUFx3_ASAP7_75t_L g1368 ( .A(n_548), .Y(n_1368) );
INVxp67_ASAP7_75t_L g549 ( .A(n_550), .Y(n_549) );
NAND2x1_ASAP7_75t_L g867 ( .A(n_551), .B(n_868), .Y(n_867) );
INVx2_ASAP7_75t_SL g551 ( .A(n_552), .Y(n_551) );
AOI22xp33_ASAP7_75t_L g765 ( .A1(n_552), .A2(n_749), .B1(n_750), .B2(n_766), .Y(n_765) );
NAND3xp33_ASAP7_75t_L g556 ( .A(n_557), .B(n_577), .C(n_580), .Y(n_556) );
BUFx3_ASAP7_75t_L g1054 ( .A(n_564), .Y(n_1054) );
INVx1_ASAP7_75t_L g570 ( .A(n_571), .Y(n_570) );
NAND2xp5_ASAP7_75t_L g581 ( .A(n_582), .B(n_584), .Y(n_581) );
INVx2_ASAP7_75t_L g586 ( .A(n_587), .Y(n_586) );
INVx1_ASAP7_75t_L g595 ( .A(n_596), .Y(n_595) );
XNOR2xp5_ASAP7_75t_L g596 ( .A(n_597), .B(n_767), .Y(n_596) );
AOI22xp5_ASAP7_75t_L g597 ( .A1(n_598), .A2(n_599), .B1(n_724), .B2(n_725), .Y(n_597) );
INVx1_ASAP7_75t_L g598 ( .A(n_599), .Y(n_598) );
NAND3xp33_ASAP7_75t_L g600 ( .A(n_601), .B(n_661), .C(n_691), .Y(n_600) );
NOR2xp33_ASAP7_75t_L g601 ( .A(n_602), .B(n_632), .Y(n_601) );
OAI33xp33_ASAP7_75t_L g602 ( .A1(n_603), .A2(n_604), .A3(n_611), .B1(n_616), .B2(n_625), .B3(n_628), .Y(n_602) );
OAI22xp33_ASAP7_75t_L g604 ( .A1(n_605), .A2(n_606), .B1(n_608), .B2(n_609), .Y(n_604) );
OAI22xp5_ASAP7_75t_L g636 ( .A1(n_605), .A2(n_629), .B1(n_637), .B2(n_641), .Y(n_636) );
OAI22xp33_ASAP7_75t_L g628 ( .A1(n_606), .A2(n_629), .B1(n_630), .B2(n_631), .Y(n_628) );
HB1xp67_ASAP7_75t_L g606 ( .A(n_607), .Y(n_606) );
OAI22xp5_ASAP7_75t_L g899 ( .A1(n_607), .A2(n_630), .B1(n_900), .B2(n_901), .Y(n_899) );
OAI22xp5_ASAP7_75t_L g650 ( .A1(n_608), .A2(n_631), .B1(n_641), .B2(n_648), .Y(n_650) );
INVx2_ASAP7_75t_L g609 ( .A(n_610), .Y(n_609) );
INVx3_ASAP7_75t_L g913 ( .A(n_610), .Y(n_913) );
OAI22xp5_ASAP7_75t_L g611 ( .A1(n_612), .A2(n_613), .B1(n_614), .B2(n_615), .Y(n_611) );
OAI22xp33_ASAP7_75t_L g651 ( .A1(n_614), .A2(n_624), .B1(n_652), .B2(n_655), .Y(n_651) );
OAI22xp5_ASAP7_75t_L g908 ( .A1(n_615), .A2(n_909), .B1(n_910), .B2(n_911), .Y(n_908) );
OAI22xp5_ASAP7_75t_L g616 ( .A1(n_617), .A2(n_621), .B1(n_622), .B2(n_624), .Y(n_616) );
INVx2_ASAP7_75t_L g617 ( .A(n_618), .Y(n_617) );
INVx8_ASAP7_75t_L g618 ( .A(n_619), .Y(n_618) );
OAI221xp5_ASAP7_75t_L g1008 ( .A1(n_619), .A2(n_990), .B1(n_1009), .B2(n_1010), .C(n_1011), .Y(n_1008) );
BUFx3_ASAP7_75t_L g1292 ( .A(n_619), .Y(n_1292) );
INVx5_ASAP7_75t_L g619 ( .A(n_620), .Y(n_619) );
INVx3_ASAP7_75t_L g905 ( .A(n_620), .Y(n_905) );
INVx2_ASAP7_75t_SL g909 ( .A(n_620), .Y(n_909) );
OAI22xp5_ASAP7_75t_L g1294 ( .A1(n_622), .A2(n_1295), .B1(n_1296), .B2(n_1299), .Y(n_1294) );
BUFx6f_ASAP7_75t_L g622 ( .A(n_623), .Y(n_622) );
INVx2_ASAP7_75t_L g701 ( .A(n_623), .Y(n_701) );
INVx1_ASAP7_75t_L g625 ( .A(n_626), .Y(n_625) );
BUFx2_ASAP7_75t_L g626 ( .A(n_627), .Y(n_626) );
BUFx2_ASAP7_75t_L g785 ( .A(n_627), .Y(n_785) );
BUFx2_ASAP7_75t_L g1040 ( .A(n_627), .Y(n_1040) );
OAI33xp33_ASAP7_75t_L g632 ( .A1(n_633), .A2(n_636), .A3(n_647), .B1(n_650), .B2(n_651), .B3(n_656), .Y(n_632) );
INVx4_ASAP7_75t_L g633 ( .A(n_634), .Y(n_633) );
NAND2xp5_ASAP7_75t_L g931 ( .A(n_634), .B(n_932), .Y(n_931) );
INVx2_ASAP7_75t_L g637 ( .A(n_638), .Y(n_637) );
INVx2_ASAP7_75t_SL g638 ( .A(n_639), .Y(n_638) );
INVx3_ASAP7_75t_L g639 ( .A(n_640), .Y(n_639) );
INVx4_ASAP7_75t_L g978 ( .A(n_640), .Y(n_978) );
BUFx6f_ASAP7_75t_L g1072 ( .A(n_640), .Y(n_1072) );
INVx2_ASAP7_75t_L g641 ( .A(n_642), .Y(n_641) );
INVx2_ASAP7_75t_L g642 ( .A(n_643), .Y(n_642) );
INVx4_ASAP7_75t_L g643 ( .A(n_644), .Y(n_643) );
BUFx6f_ASAP7_75t_L g808 ( .A(n_644), .Y(n_808) );
INVx8_ASAP7_75t_L g644 ( .A(n_645), .Y(n_644) );
OR2x2_ASAP7_75t_L g683 ( .A(n_645), .B(n_669), .Y(n_683) );
BUFx6f_ASAP7_75t_L g645 ( .A(n_646), .Y(n_645) );
BUFx2_ASAP7_75t_L g648 ( .A(n_649), .Y(n_648) );
INVx1_ASAP7_75t_L g952 ( .A(n_649), .Y(n_952) );
BUFx2_ASAP7_75t_L g1067 ( .A(n_649), .Y(n_1067) );
INVx2_ASAP7_75t_L g652 ( .A(n_653), .Y(n_652) );
INVx2_ASAP7_75t_SL g653 ( .A(n_654), .Y(n_653) );
INVx2_ASAP7_75t_L g656 ( .A(n_657), .Y(n_656) );
INVx1_ASAP7_75t_L g657 ( .A(n_658), .Y(n_657) );
INVx1_ASAP7_75t_L g659 ( .A(n_660), .Y(n_659) );
OAI31xp33_ASAP7_75t_SL g661 ( .A1(n_662), .A2(n_674), .A3(n_684), .B(n_688), .Y(n_661) );
INVx1_ASAP7_75t_L g663 ( .A(n_664), .Y(n_663) );
AOI22xp33_ASAP7_75t_L g666 ( .A1(n_667), .A2(n_670), .B1(n_671), .B2(n_672), .Y(n_666) );
BUFx3_ASAP7_75t_L g667 ( .A(n_668), .Y(n_667) );
AOI22xp33_ASAP7_75t_L g704 ( .A1(n_670), .A2(n_705), .B1(n_709), .B2(n_712), .Y(n_704) );
BUFx3_ASAP7_75t_L g672 ( .A(n_673), .Y(n_672) );
INVx1_ASAP7_75t_L g675 ( .A(n_676), .Y(n_675) );
INVx1_ASAP7_75t_L g676 ( .A(n_677), .Y(n_676) );
INVx2_ASAP7_75t_L g679 ( .A(n_680), .Y(n_679) );
INVx2_ASAP7_75t_L g680 ( .A(n_681), .Y(n_680) );
INVx2_ASAP7_75t_L g681 ( .A(n_682), .Y(n_681) );
INVx1_ASAP7_75t_L g682 ( .A(n_683), .Y(n_682) );
INVx3_ASAP7_75t_SL g686 ( .A(n_687), .Y(n_686) );
BUFx3_ASAP7_75t_L g688 ( .A(n_689), .Y(n_688) );
OAI31xp33_ASAP7_75t_SL g691 ( .A1(n_692), .A2(n_699), .A3(n_713), .B(n_719), .Y(n_691) );
INVx1_ASAP7_75t_L g693 ( .A(n_694), .Y(n_693) );
INVx1_ASAP7_75t_L g694 ( .A(n_695), .Y(n_694) );
INVx1_ASAP7_75t_L g696 ( .A(n_697), .Y(n_696) );
INVx2_ASAP7_75t_L g700 ( .A(n_701), .Y(n_700) );
CKINVDCx8_ASAP7_75t_R g702 ( .A(n_703), .Y(n_702) );
BUFx3_ASAP7_75t_L g705 ( .A(n_706), .Y(n_705) );
AND2x2_ASAP7_75t_L g706 ( .A(n_707), .B(n_708), .Y(n_706) );
AND2x4_ASAP7_75t_L g710 ( .A(n_707), .B(n_711), .Y(n_710) );
BUFx6f_ASAP7_75t_L g709 ( .A(n_710), .Y(n_709) );
INVx1_ASAP7_75t_L g714 ( .A(n_715), .Y(n_714) );
INVx2_ASAP7_75t_SL g715 ( .A(n_716), .Y(n_715) );
BUFx3_ASAP7_75t_L g717 ( .A(n_718), .Y(n_717) );
AND2x2_ASAP7_75t_L g719 ( .A(n_720), .B(n_722), .Y(n_719) );
INVx1_ASAP7_75t_SL g720 ( .A(n_721), .Y(n_720) );
INVx1_ASAP7_75t_L g722 ( .A(n_723), .Y(n_722) );
INVx1_ASAP7_75t_L g724 ( .A(n_725), .Y(n_724) );
INVx1_ASAP7_75t_L g725 ( .A(n_726), .Y(n_725) );
AND2x2_ASAP7_75t_L g727 ( .A(n_728), .B(n_746), .Y(n_727) );
NAND3xp33_ASAP7_75t_SL g732 ( .A(n_733), .B(n_736), .C(n_745), .Y(n_732) );
AOI22xp5_ASAP7_75t_L g736 ( .A1(n_737), .A2(n_740), .B1(n_742), .B2(n_744), .Y(n_736) );
INVx2_ASAP7_75t_L g1301 ( .A(n_741), .Y(n_1301) );
AND5x1_ASAP7_75t_L g971 ( .A(n_745), .B(n_972), .C(n_997), .D(n_1013), .E(n_1017), .Y(n_971) );
NAND3xp33_ASAP7_75t_L g747 ( .A(n_748), .B(n_751), .C(n_759), .Y(n_747) );
INVx2_ASAP7_75t_L g835 ( .A(n_752), .Y(n_835) );
AND2x4_ASAP7_75t_L g961 ( .A(n_753), .B(n_962), .Y(n_961) );
INVx1_ASAP7_75t_L g799 ( .A(n_755), .Y(n_799) );
INVx2_ASAP7_75t_L g755 ( .A(n_756), .Y(n_755) );
NAND2xp5_ASAP7_75t_L g974 ( .A(n_760), .B(n_975), .Y(n_974) );
AOI222xp33_ASAP7_75t_L g873 ( .A1(n_766), .A2(n_850), .B1(n_874), .B2(n_875), .C1(n_876), .C2(n_877), .Y(n_873) );
INVxp67_ASAP7_75t_SL g767 ( .A(n_768), .Y(n_767) );
NAND3xp33_ASAP7_75t_L g769 ( .A(n_770), .B(n_789), .C(n_793), .Y(n_769) );
NAND2xp5_ASAP7_75t_L g771 ( .A(n_772), .B(n_777), .Y(n_771) );
AOI22xp33_ASAP7_75t_L g772 ( .A1(n_773), .A2(n_774), .B1(n_775), .B2(n_776), .Y(n_772) );
AO22x1_ASAP7_75t_L g1026 ( .A1(n_774), .A2(n_776), .B1(n_1027), .B2(n_1028), .Y(n_1026) );
AOI221x1_ASAP7_75t_L g997 ( .A1(n_776), .A2(n_975), .B1(n_981), .B2(n_998), .C(n_999), .Y(n_997) );
AOI22xp33_ASAP7_75t_L g1373 ( .A1(n_776), .A2(n_998), .B1(n_1343), .B2(n_1374), .Y(n_1373) );
AOI33xp33_ASAP7_75t_L g777 ( .A1(n_778), .A2(n_779), .A3(n_781), .B1(n_784), .B2(n_785), .B3(n_786), .Y(n_777) );
AOI33xp33_ASAP7_75t_L g1033 ( .A1(n_778), .A2(n_1034), .A3(n_1035), .B1(n_1038), .B2(n_1040), .B3(n_1041), .Y(n_1033) );
INVx2_ASAP7_75t_L g782 ( .A(n_783), .Y(n_782) );
INVx2_ASAP7_75t_L g1274 ( .A(n_792), .Y(n_1274) );
OAI21xp5_ASAP7_75t_L g793 ( .A1(n_794), .A2(n_807), .B(n_821), .Y(n_793) );
INVx1_ASAP7_75t_L g798 ( .A(n_799), .Y(n_798) );
INVx1_ASAP7_75t_L g805 ( .A(n_806), .Y(n_805) );
INVx5_ASAP7_75t_L g1074 ( .A(n_808), .Y(n_1074) );
NAND2xp5_ASAP7_75t_L g809 ( .A(n_810), .B(n_818), .Y(n_809) );
INVx2_ASAP7_75t_L g811 ( .A(n_812), .Y(n_811) );
INVx1_ASAP7_75t_L g1053 ( .A(n_812), .Y(n_1053) );
BUFx2_ASAP7_75t_L g812 ( .A(n_813), .Y(n_812) );
HB1xp67_ASAP7_75t_L g814 ( .A(n_815), .Y(n_814) );
INVx2_ASAP7_75t_L g815 ( .A(n_816), .Y(n_815) );
INVx2_ASAP7_75t_L g839 ( .A(n_816), .Y(n_839) );
INVx2_ASAP7_75t_L g821 ( .A(n_822), .Y(n_821) );
INVx1_ASAP7_75t_L g822 ( .A(n_823), .Y(n_822) );
HB1xp67_ASAP7_75t_L g993 ( .A(n_823), .Y(n_993) );
INVx2_ASAP7_75t_L g825 ( .A(n_826), .Y(n_825) );
INVx1_ASAP7_75t_L g826 ( .A(n_827), .Y(n_826) );
INVx1_ASAP7_75t_L g827 ( .A(n_828), .Y(n_827) );
AO22x2_ASAP7_75t_L g828 ( .A1(n_829), .A2(n_1020), .B1(n_1077), .B2(n_1078), .Y(n_828) );
INVx1_ASAP7_75t_L g1077 ( .A(n_829), .Y(n_1077) );
XNOR2xp5_ASAP7_75t_L g829 ( .A(n_830), .B(n_970), .Y(n_829) );
OAI22xp5_ASAP7_75t_L g830 ( .A1(n_831), .A2(n_885), .B1(n_968), .B2(n_969), .Y(n_830) );
INVx1_ASAP7_75t_L g969 ( .A(n_831), .Y(n_969) );
NAND3xp33_ASAP7_75t_L g831 ( .A(n_832), .B(n_878), .C(n_882), .Y(n_831) );
INVx1_ASAP7_75t_L g879 ( .A(n_833), .Y(n_879) );
AOI22xp5_ASAP7_75t_L g836 ( .A1(n_837), .A2(n_838), .B1(n_840), .B2(n_842), .Y(n_836) );
AOI22xp5_ASAP7_75t_L g843 ( .A1(n_844), .A2(n_851), .B1(n_852), .B2(n_853), .Y(n_843) );
INVx1_ASAP7_75t_L g848 ( .A(n_849), .Y(n_848) );
AOI22xp5_ASAP7_75t_L g976 ( .A1(n_851), .A2(n_852), .B1(n_977), .B2(n_983), .Y(n_976) );
INVx1_ASAP7_75t_L g880 ( .A(n_855), .Y(n_880) );
AND2x2_ASAP7_75t_L g855 ( .A(n_856), .B(n_864), .Y(n_855) );
INVx1_ASAP7_75t_L g884 ( .A(n_866), .Y(n_884) );
NAND2xp5_ASAP7_75t_L g866 ( .A(n_867), .B(n_872), .Y(n_866) );
INVx2_ASAP7_75t_L g868 ( .A(n_869), .Y(n_868) );
AOI22xp33_ASAP7_75t_L g889 ( .A1(n_869), .A2(n_890), .B1(n_891), .B2(n_892), .Y(n_889) );
AND2x4_ASAP7_75t_L g869 ( .A(n_870), .B(n_871), .Y(n_869) );
INVx1_ASAP7_75t_L g883 ( .A(n_873), .Y(n_883) );
AOI22xp5_ASAP7_75t_L g995 ( .A1(n_874), .A2(n_876), .B1(n_982), .B2(n_996), .Y(n_995) );
OAI21xp5_ASAP7_75t_L g878 ( .A1(n_879), .A2(n_880), .B(n_881), .Y(n_878) );
OAI21xp33_ASAP7_75t_L g882 ( .A1(n_881), .A2(n_883), .B(n_884), .Y(n_882) );
INVx1_ASAP7_75t_L g968 ( .A(n_885), .Y(n_968) );
XNOR2xp5_ASAP7_75t_L g885 ( .A(n_886), .B(n_887), .Y(n_885) );
NOR2x1_ASAP7_75t_L g887 ( .A(n_888), .B(n_928), .Y(n_887) );
NAND2xp5_ASAP7_75t_L g888 ( .A(n_889), .B(n_893), .Y(n_888) );
INVx3_ASAP7_75t_L g1016 ( .A(n_891), .Y(n_1016) );
INVx2_ASAP7_75t_L g896 ( .A(n_897), .Y(n_896) );
HB1xp67_ASAP7_75t_L g923 ( .A(n_897), .Y(n_923) );
OAI221xp5_ASAP7_75t_L g898 ( .A1(n_899), .A2(n_902), .B1(n_908), .B2(n_912), .C(n_917), .Y(n_898) );
OAI221xp5_ASAP7_75t_L g902 ( .A1(n_903), .A2(n_904), .B1(n_905), .B2(n_906), .C(n_907), .Y(n_902) );
OR2x6_ASAP7_75t_L g917 ( .A(n_903), .B(n_918), .Y(n_917) );
INVx1_ASAP7_75t_L g1370 ( .A(n_903), .Y(n_1370) );
OAI211xp5_ASAP7_75t_L g950 ( .A1(n_904), .A2(n_951), .B(n_953), .C(n_954), .Y(n_950) );
OAI221xp5_ASAP7_75t_L g1001 ( .A1(n_909), .A2(n_1002), .B1(n_1003), .B2(n_1004), .C(n_1005), .Y(n_1001) );
OAI21xp5_ASAP7_75t_SL g912 ( .A1(n_913), .A2(n_914), .B(n_915), .Y(n_912) );
INVx1_ASAP7_75t_L g1307 ( .A(n_916), .Y(n_1307) );
AOI22xp5_ASAP7_75t_L g934 ( .A1(n_921), .A2(n_935), .B1(n_937), .B2(n_938), .Y(n_934) );
INVx1_ASAP7_75t_L g922 ( .A(n_923), .Y(n_922) );
INVx4_ASAP7_75t_L g924 ( .A(n_925), .Y(n_924) );
INVx2_ASAP7_75t_L g926 ( .A(n_927), .Y(n_926) );
NAND3xp33_ASAP7_75t_L g928 ( .A(n_929), .B(n_957), .C(n_963), .Y(n_928) );
NOR3xp33_ASAP7_75t_SL g929 ( .A(n_930), .B(n_944), .C(n_947), .Y(n_929) );
OAI21xp5_ASAP7_75t_SL g930 ( .A1(n_931), .A2(n_933), .B(n_934), .Y(n_930) );
INVx1_ASAP7_75t_SL g935 ( .A(n_936), .Y(n_935) );
INVx2_ASAP7_75t_SL g938 ( .A(n_939), .Y(n_938) );
NAND2x2_ASAP7_75t_L g939 ( .A(n_940), .B(n_942), .Y(n_939) );
INVx1_ASAP7_75t_L g956 ( .A(n_940), .Y(n_956) );
INVx2_ASAP7_75t_L g940 ( .A(n_941), .Y(n_940) );
INVx2_ASAP7_75t_SL g942 ( .A(n_943), .Y(n_942) );
INVx1_ASAP7_75t_L g962 ( .A(n_946), .Y(n_962) );
OAI21xp5_ASAP7_75t_L g947 ( .A1(n_948), .A2(n_950), .B(n_955), .Y(n_947) );
INVx2_ASAP7_75t_L g948 ( .A(n_949), .Y(n_948) );
INVx2_ASAP7_75t_L g951 ( .A(n_952), .Y(n_951) );
NAND2xp5_ASAP7_75t_L g957 ( .A(n_958), .B(n_959), .Y(n_957) );
INVx1_ASAP7_75t_L g960 ( .A(n_961), .Y(n_960) );
NAND2xp5_ASAP7_75t_L g963 ( .A(n_964), .B(n_965), .Y(n_963) );
AOI21xp5_ASAP7_75t_L g972 ( .A1(n_973), .A2(n_993), .B(n_994), .Y(n_972) );
NAND4xp25_ASAP7_75t_L g973 ( .A(n_974), .B(n_976), .C(n_984), .D(n_989), .Y(n_973) );
OAI22xp5_ASAP7_75t_SL g999 ( .A1(n_1000), .A2(n_1001), .B1(n_1007), .B2(n_1008), .Y(n_999) );
OAI22xp5_ASAP7_75t_L g1363 ( .A1(n_1009), .A2(n_1301), .B1(n_1364), .B2(n_1365), .Y(n_1363) );
NAND2xp5_ASAP7_75t_L g1013 ( .A(n_1014), .B(n_1015), .Y(n_1013) );
NAND2xp5_ASAP7_75t_L g1017 ( .A(n_1018), .B(n_1019), .Y(n_1017) );
NAND2xp5_ASAP7_75t_L g1030 ( .A(n_1019), .B(n_1031), .Y(n_1030) );
NAND2xp5_ASAP7_75t_L g1313 ( .A(n_1019), .B(n_1288), .Y(n_1313) );
NAND2xp5_ASAP7_75t_L g1375 ( .A(n_1019), .B(n_1346), .Y(n_1375) );
INVx2_ASAP7_75t_L g1078 ( .A(n_1020), .Y(n_1078) );
XOR2x2_ASAP7_75t_L g1020 ( .A(n_1021), .B(n_1076), .Y(n_1020) );
NAND2xp5_ASAP7_75t_SL g1021 ( .A(n_1022), .B(n_1048), .Y(n_1021) );
NAND2xp5_ASAP7_75t_L g1024 ( .A(n_1025), .B(n_1033), .Y(n_1024) );
NOR2xp33_ASAP7_75t_L g1025 ( .A(n_1026), .B(n_1029), .Y(n_1025) );
NAND2xp5_ASAP7_75t_SL g1029 ( .A(n_1030), .B(n_1032), .Y(n_1029) );
NAND4xp25_ASAP7_75t_L g1372 ( .A(n_1032), .B(n_1373), .C(n_1375), .D(n_1376), .Y(n_1372) );
INVx2_ASAP7_75t_L g1036 ( .A(n_1037), .Y(n_1036) );
INVx1_ASAP7_75t_L g1042 ( .A(n_1043), .Y(n_1042) );
NAND3xp33_ASAP7_75t_SL g1049 ( .A(n_1050), .B(n_1051), .C(n_1059), .Y(n_1049) );
INVx1_ASAP7_75t_SL g1057 ( .A(n_1058), .Y(n_1057) );
INVx2_ASAP7_75t_L g1065 ( .A(n_1066), .Y(n_1065) );
INVx4_ASAP7_75t_L g1066 ( .A(n_1067), .Y(n_1066) );
OAI22xp5_ASAP7_75t_L g1069 ( .A1(n_1070), .A2(n_1071), .B1(n_1073), .B2(n_1074), .Y(n_1069) );
INVx2_ASAP7_75t_L g1071 ( .A(n_1072), .Y(n_1071) );
OAI221xp5_ASAP7_75t_L g1079 ( .A1(n_1080), .A2(n_1266), .B1(n_1268), .B2(n_1316), .C(n_1322), .Y(n_1079) );
NOR2xp67_ASAP7_75t_SL g1080 ( .A(n_1081), .B(n_1204), .Y(n_1080) );
NAND4xp25_ASAP7_75t_L g1081 ( .A(n_1082), .B(n_1160), .C(n_1184), .D(n_1198), .Y(n_1081) );
OAI21xp5_ASAP7_75t_L g1082 ( .A1(n_1083), .A2(n_1144), .B(n_1150), .Y(n_1082) );
OAI321xp33_ASAP7_75t_L g1083 ( .A1(n_1084), .A2(n_1109), .A3(n_1120), .B1(n_1124), .B2(n_1127), .C(n_1130), .Y(n_1083) );
INVx1_ASAP7_75t_L g1084 ( .A(n_1085), .Y(n_1084) );
AND2x2_ASAP7_75t_L g1161 ( .A(n_1085), .B(n_1162), .Y(n_1161) );
AND2x2_ASAP7_75t_L g1085 ( .A(n_1086), .B(n_1101), .Y(n_1085) );
OR2x2_ASAP7_75t_L g1127 ( .A(n_1086), .B(n_1128), .Y(n_1127) );
OR2x2_ASAP7_75t_L g1173 ( .A(n_1086), .B(n_1102), .Y(n_1173) );
AND2x2_ASAP7_75t_L g1186 ( .A(n_1086), .B(n_1176), .Y(n_1186) );
NOR2xp33_ASAP7_75t_L g1250 ( .A(n_1086), .B(n_1177), .Y(n_1250) );
INVx1_ASAP7_75t_L g1086 ( .A(n_1087), .Y(n_1086) );
OR2x2_ASAP7_75t_L g1148 ( .A(n_1087), .B(n_1149), .Y(n_1148) );
OR2x2_ASAP7_75t_L g1192 ( .A(n_1087), .B(n_1103), .Y(n_1192) );
AND2x2_ASAP7_75t_L g1217 ( .A(n_1087), .B(n_1177), .Y(n_1217) );
AND2x2_ASAP7_75t_L g1222 ( .A(n_1087), .B(n_1213), .Y(n_1222) );
OR2x2_ASAP7_75t_L g1236 ( .A(n_1087), .B(n_1177), .Y(n_1236) );
NAND2xp5_ASAP7_75t_SL g1245 ( .A(n_1087), .B(n_1135), .Y(n_1245) );
OR2x2_ASAP7_75t_L g1258 ( .A(n_1087), .B(n_1135), .Y(n_1258) );
AND2x2_ASAP7_75t_L g1087 ( .A(n_1088), .B(n_1096), .Y(n_1087) );
AND2x2_ASAP7_75t_L g1167 ( .A(n_1088), .B(n_1096), .Y(n_1167) );
AND2x4_ASAP7_75t_L g1089 ( .A(n_1090), .B(n_1091), .Y(n_1089) );
AND2x6_ASAP7_75t_L g1094 ( .A(n_1090), .B(n_1095), .Y(n_1094) );
AND2x6_ASAP7_75t_L g1097 ( .A(n_1090), .B(n_1098), .Y(n_1097) );
AND2x2_ASAP7_75t_L g1099 ( .A(n_1090), .B(n_1100), .Y(n_1099) );
AND2x2_ASAP7_75t_L g1118 ( .A(n_1090), .B(n_1100), .Y(n_1118) );
AND2x2_ASAP7_75t_L g1123 ( .A(n_1090), .B(n_1100), .Y(n_1123) );
NAND2xp5_ASAP7_75t_L g1155 ( .A(n_1090), .B(n_1091), .Y(n_1155) );
AND2x2_ASAP7_75t_L g1091 ( .A(n_1092), .B(n_1093), .Y(n_1091) );
INVx2_ASAP7_75t_L g1157 ( .A(n_1094), .Y(n_1157) );
OAI21xp5_ASAP7_75t_L g1378 ( .A1(n_1100), .A2(n_1379), .B(n_1380), .Y(n_1378) );
INVx1_ASAP7_75t_L g1101 ( .A(n_1102), .Y(n_1101) );
OR2x2_ASAP7_75t_L g1102 ( .A(n_1103), .B(n_1106), .Y(n_1102) );
NAND2xp5_ASAP7_75t_L g1128 ( .A(n_1103), .B(n_1129), .Y(n_1128) );
INVx2_ASAP7_75t_L g1177 ( .A(n_1103), .Y(n_1177) );
AOI321xp33_ASAP7_75t_L g1198 ( .A1(n_1103), .A2(n_1161), .A3(n_1194), .B1(n_1199), .B2(n_1201), .C(n_1203), .Y(n_1198) );
AND2x2_ASAP7_75t_L g1213 ( .A(n_1103), .B(n_1106), .Y(n_1213) );
NAND2x1p5_ASAP7_75t_L g1103 ( .A(n_1104), .B(n_1105), .Y(n_1103) );
INVx1_ASAP7_75t_L g1129 ( .A(n_1106), .Y(n_1129) );
NOR2xp33_ASAP7_75t_L g1133 ( .A(n_1106), .B(n_1134), .Y(n_1133) );
INVx1_ASAP7_75t_L g1149 ( .A(n_1106), .Y(n_1149) );
AND2x2_ASAP7_75t_L g1176 ( .A(n_1106), .B(n_1177), .Y(n_1176) );
AND2x2_ASAP7_75t_L g1106 ( .A(n_1107), .B(n_1108), .Y(n_1106) );
INVx1_ASAP7_75t_L g1109 ( .A(n_1110), .Y(n_1109) );
AND2x2_ASAP7_75t_L g1206 ( .A(n_1110), .B(n_1164), .Y(n_1206) );
AND2x2_ASAP7_75t_L g1110 ( .A(n_1111), .B(n_1115), .Y(n_1110) );
OR2x2_ASAP7_75t_L g1132 ( .A(n_1111), .B(n_1120), .Y(n_1132) );
AND2x2_ASAP7_75t_L g1146 ( .A(n_1111), .B(n_1126), .Y(n_1146) );
AND2x2_ASAP7_75t_L g1168 ( .A(n_1111), .B(n_1120), .Y(n_1168) );
OR2x2_ASAP7_75t_L g1181 ( .A(n_1111), .B(n_1143), .Y(n_1181) );
OR2x2_ASAP7_75t_L g1195 ( .A(n_1111), .B(n_1116), .Y(n_1195) );
INVx1_ASAP7_75t_L g1211 ( .A(n_1111), .Y(n_1211) );
INVx2_ASAP7_75t_L g1234 ( .A(n_1111), .Y(n_1234) );
INVx2_ASAP7_75t_L g1111 ( .A(n_1112), .Y(n_1111) );
OR2x2_ASAP7_75t_L g1200 ( .A(n_1112), .B(n_1143), .Y(n_1200) );
NAND2xp5_ASAP7_75t_L g1112 ( .A(n_1113), .B(n_1114), .Y(n_1112) );
OR2x2_ASAP7_75t_L g1125 ( .A(n_1115), .B(n_1126), .Y(n_1125) );
INVx2_ASAP7_75t_L g1138 ( .A(n_1115), .Y(n_1138) );
AND2x2_ASAP7_75t_L g1172 ( .A(n_1115), .B(n_1164), .Y(n_1172) );
AND2x2_ASAP7_75t_L g1189 ( .A(n_1115), .B(n_1165), .Y(n_1189) );
INVx1_ASAP7_75t_L g1115 ( .A(n_1116), .Y(n_1115) );
INVx1_ASAP7_75t_L g1143 ( .A(n_1116), .Y(n_1143) );
NAND2xp5_ASAP7_75t_L g1116 ( .A(n_1117), .B(n_1119), .Y(n_1116) );
INVx3_ASAP7_75t_L g1126 ( .A(n_1120), .Y(n_1126) );
INVx1_ASAP7_75t_L g1197 ( .A(n_1120), .Y(n_1197) );
AND2x2_ASAP7_75t_L g1120 ( .A(n_1121), .B(n_1122), .Y(n_1120) );
HB1xp67_ASAP7_75t_L g1267 ( .A(n_1123), .Y(n_1267) );
INVx1_ASAP7_75t_L g1124 ( .A(n_1125), .Y(n_1124) );
OAI322xp33_ASAP7_75t_L g1229 ( .A1(n_1125), .A2(n_1127), .A3(n_1167), .B1(n_1230), .B2(n_1232), .C1(n_1233), .C2(n_1234), .Y(n_1229) );
CKINVDCx14_ASAP7_75t_R g1218 ( .A(n_1126), .Y(n_1218) );
OR2x2_ASAP7_75t_L g1240 ( .A(n_1126), .B(n_1200), .Y(n_1240) );
OR2x2_ASAP7_75t_L g1259 ( .A(n_1126), .B(n_1181), .Y(n_1259) );
OR2x2_ASAP7_75t_L g1264 ( .A(n_1126), .B(n_1142), .Y(n_1264) );
INVx1_ASAP7_75t_L g1190 ( .A(n_1127), .Y(n_1190) );
AOI21xp33_ASAP7_75t_SL g1191 ( .A1(n_1127), .A2(n_1192), .B(n_1193), .Y(n_1191) );
INVx1_ASAP7_75t_L g1139 ( .A(n_1128), .Y(n_1139) );
OR2x2_ASAP7_75t_L g1166 ( .A(n_1128), .B(n_1167), .Y(n_1166) );
NAND2xp5_ASAP7_75t_L g1230 ( .A(n_1128), .B(n_1231), .Y(n_1230) );
OR2x2_ASAP7_75t_L g1244 ( .A(n_1128), .B(n_1245), .Y(n_1244) );
AOI22xp5_ASAP7_75t_L g1130 ( .A1(n_1131), .A2(n_1133), .B1(n_1139), .B2(n_1140), .Y(n_1130) );
OAI21xp5_ASAP7_75t_L g1227 ( .A1(n_1131), .A2(n_1175), .B(n_1228), .Y(n_1227) );
CKINVDCx14_ASAP7_75t_R g1131 ( .A(n_1132), .Y(n_1131) );
NOR3xp33_ASAP7_75t_L g1203 ( .A(n_1132), .B(n_1135), .C(n_1174), .Y(n_1203) );
OR2x2_ASAP7_75t_L g1232 ( .A(n_1132), .B(n_1138), .Y(n_1232) );
NAND2xp5_ASAP7_75t_L g1134 ( .A(n_1135), .B(n_1138), .Y(n_1134) );
INVx4_ASAP7_75t_L g1141 ( .A(n_1135), .Y(n_1141) );
INVx4_ASAP7_75t_L g1165 ( .A(n_1135), .Y(n_1165) );
AND2x2_ASAP7_75t_L g1185 ( .A(n_1135), .B(n_1186), .Y(n_1185) );
NOR2xp33_ASAP7_75t_L g1251 ( .A(n_1135), .B(n_1236), .Y(n_1251) );
NOR2xp33_ASAP7_75t_L g1253 ( .A(n_1135), .B(n_1195), .Y(n_1253) );
AND2x4_ASAP7_75t_SL g1135 ( .A(n_1136), .B(n_1137), .Y(n_1135) );
AND2x2_ASAP7_75t_L g1215 ( .A(n_1139), .B(n_1165), .Y(n_1215) );
INVx1_ASAP7_75t_L g1147 ( .A(n_1140), .Y(n_1147) );
AOI21xp33_ASAP7_75t_L g1214 ( .A1(n_1140), .A2(n_1149), .B(n_1215), .Y(n_1214) );
NAND2xp5_ASAP7_75t_L g1225 ( .A(n_1140), .B(n_1197), .Y(n_1225) );
AND2x2_ASAP7_75t_L g1140 ( .A(n_1141), .B(n_1142), .Y(n_1140) );
CKINVDCx5p33_ASAP7_75t_R g1162 ( .A(n_1141), .Y(n_1162) );
NOR2xp33_ASAP7_75t_L g1228 ( .A(n_1141), .B(n_1148), .Y(n_1228) );
OR2x2_ASAP7_75t_L g1238 ( .A(n_1141), .B(n_1166), .Y(n_1238) );
AND2x2_ASAP7_75t_L g1249 ( .A(n_1141), .B(n_1250), .Y(n_1249) );
NAND2xp5_ASAP7_75t_L g1145 ( .A(n_1142), .B(n_1146), .Y(n_1145) );
AOI221xp5_ASAP7_75t_L g1205 ( .A1(n_1142), .A2(n_1177), .B1(n_1183), .B2(n_1206), .C(n_1207), .Y(n_1205) );
NOR3xp33_ASAP7_75t_L g1243 ( .A(n_1142), .B(n_1244), .C(n_1246), .Y(n_1243) );
AOI22xp33_ASAP7_75t_L g1248 ( .A1(n_1142), .A2(n_1211), .B1(n_1249), .B2(n_1251), .Y(n_1248) );
INVx1_ASAP7_75t_L g1142 ( .A(n_1143), .Y(n_1142) );
AOI21xp33_ASAP7_75t_L g1144 ( .A1(n_1145), .A2(n_1147), .B(n_1148), .Y(n_1144) );
INVx1_ASAP7_75t_L g1187 ( .A(n_1145), .Y(n_1187) );
AND2x2_ASAP7_75t_L g1171 ( .A(n_1146), .B(n_1172), .Y(n_1171) );
AOI221xp5_ASAP7_75t_L g1184 ( .A1(n_1146), .A2(n_1185), .B1(n_1187), .B2(n_1188), .C(n_1191), .Y(n_1184) );
INVx1_ASAP7_75t_L g1255 ( .A(n_1146), .Y(n_1255) );
INVx1_ASAP7_75t_L g1209 ( .A(n_1148), .Y(n_1209) );
INVx1_ASAP7_75t_L g1150 ( .A(n_1151), .Y(n_1150) );
OAI321xp33_ASAP7_75t_L g1204 ( .A1(n_1151), .A2(n_1152), .A3(n_1205), .B1(n_1216), .B2(n_1219), .C(n_1242), .Y(n_1204) );
INVx2_ASAP7_75t_L g1151 ( .A(n_1152), .Y(n_1151) );
INVx1_ASAP7_75t_L g1152 ( .A(n_1153), .Y(n_1152) );
INVx1_ASAP7_75t_L g1153 ( .A(n_1154), .Y(n_1153) );
NAND2xp5_ASAP7_75t_L g1202 ( .A(n_1154), .B(n_1165), .Y(n_1202) );
OAI221xp5_ASAP7_75t_L g1154 ( .A1(n_1155), .A2(n_1156), .B1(n_1157), .B2(n_1158), .C(n_1159), .Y(n_1154) );
O2A1O1Ixp33_ASAP7_75t_L g1160 ( .A1(n_1161), .A2(n_1163), .B(n_1168), .C(n_1169), .Y(n_1160) );
AND2x2_ASAP7_75t_L g1179 ( .A(n_1162), .B(n_1180), .Y(n_1179) );
NAND2xp5_ASAP7_75t_L g1224 ( .A(n_1162), .B(n_1199), .Y(n_1224) );
NOR2xp33_ASAP7_75t_L g1163 ( .A(n_1164), .B(n_1166), .Y(n_1163) );
AND2x2_ASAP7_75t_L g1196 ( .A(n_1164), .B(n_1197), .Y(n_1196) );
CKINVDCx5p33_ASAP7_75t_R g1164 ( .A(n_1165), .Y(n_1164) );
NAND2xp5_ASAP7_75t_SL g1208 ( .A(n_1165), .B(n_1209), .Y(n_1208) );
NAND2x1_ASAP7_75t_L g1221 ( .A(n_1165), .B(n_1222), .Y(n_1221) );
INVx1_ASAP7_75t_L g1183 ( .A(n_1166), .Y(n_1183) );
AND2x2_ASAP7_75t_L g1175 ( .A(n_1167), .B(n_1176), .Y(n_1175) );
OR2x2_ASAP7_75t_L g1241 ( .A(n_1167), .B(n_1212), .Y(n_1241) );
INVx1_ASAP7_75t_L g1246 ( .A(n_1168), .Y(n_1246) );
OAI221xp5_ASAP7_75t_L g1169 ( .A1(n_1170), .A2(n_1173), .B1(n_1174), .B2(n_1178), .C(n_1182), .Y(n_1169) );
INVx1_ASAP7_75t_L g1170 ( .A(n_1171), .Y(n_1170) );
OAI21xp5_ASAP7_75t_SL g1182 ( .A1(n_1171), .A2(n_1179), .B(n_1183), .Y(n_1182) );
INVxp67_ASAP7_75t_L g1237 ( .A(n_1172), .Y(n_1237) );
NOR2xp33_ASAP7_75t_L g1261 ( .A(n_1173), .B(n_1262), .Y(n_1261) );
OAI32xp33_ASAP7_75t_L g1263 ( .A1(n_1174), .A2(n_1181), .A3(n_1202), .B1(n_1264), .B2(n_1265), .Y(n_1263) );
INVx1_ASAP7_75t_L g1174 ( .A(n_1175), .Y(n_1174) );
INVx1_ASAP7_75t_L g1231 ( .A(n_1176), .Y(n_1231) );
NAND3xp33_ASAP7_75t_L g1233 ( .A(n_1176), .B(n_1189), .C(n_1197), .Y(n_1233) );
NAND2xp5_ASAP7_75t_L g1265 ( .A(n_1176), .B(n_1257), .Y(n_1265) );
INVx1_ASAP7_75t_L g1178 ( .A(n_1179), .Y(n_1178) );
CKINVDCx5p33_ASAP7_75t_R g1180 ( .A(n_1181), .Y(n_1180) );
OAI221xp5_ASAP7_75t_L g1207 ( .A1(n_1181), .A2(n_1208), .B1(n_1210), .B2(n_1212), .C(n_1214), .Y(n_1207) );
AND2x2_ASAP7_75t_L g1188 ( .A(n_1189), .B(n_1190), .Y(n_1188) );
NAND2xp5_ASAP7_75t_L g1193 ( .A(n_1194), .B(n_1196), .Y(n_1193) );
INVx1_ASAP7_75t_L g1194 ( .A(n_1195), .Y(n_1194) );
OR2x2_ASAP7_75t_L g1262 ( .A(n_1195), .B(n_1197), .Y(n_1262) );
OAI21xp33_ASAP7_75t_L g1247 ( .A1(n_1197), .A2(n_1248), .B(n_1252), .Y(n_1247) );
CKINVDCx5p33_ASAP7_75t_R g1199 ( .A(n_1200), .Y(n_1199) );
OAI322xp33_ASAP7_75t_L g1254 ( .A1(n_1200), .A2(n_1202), .A3(n_1241), .B1(n_1255), .B2(n_1256), .C1(n_1259), .C2(n_1260), .Y(n_1254) );
INVx1_ASAP7_75t_L g1201 ( .A(n_1202), .Y(n_1201) );
AOI21xp33_ASAP7_75t_L g1216 ( .A1(n_1206), .A2(n_1217), .B(n_1218), .Y(n_1216) );
NOR2xp33_ASAP7_75t_L g1220 ( .A(n_1210), .B(n_1221), .Y(n_1220) );
INVx1_ASAP7_75t_L g1210 ( .A(n_1211), .Y(n_1210) );
INVx1_ASAP7_75t_L g1212 ( .A(n_1213), .Y(n_1212) );
NAND2xp5_ASAP7_75t_L g1256 ( .A(n_1213), .B(n_1257), .Y(n_1256) );
CKINVDCx14_ASAP7_75t_R g1226 ( .A(n_1217), .Y(n_1226) );
NAND2xp5_ASAP7_75t_L g1252 ( .A(n_1217), .B(n_1253), .Y(n_1252) );
O2A1O1Ixp33_ASAP7_75t_L g1235 ( .A1(n_1218), .A2(n_1236), .B(n_1237), .C(n_1238), .Y(n_1235) );
NOR5xp2_ASAP7_75t_L g1219 ( .A(n_1220), .B(n_1223), .C(n_1229), .D(n_1235), .E(n_1239), .Y(n_1219) );
INVx1_ASAP7_75t_L g1260 ( .A(n_1222), .Y(n_1260) );
A2O1A1Ixp33_ASAP7_75t_L g1223 ( .A1(n_1224), .A2(n_1225), .B(n_1226), .C(n_1227), .Y(n_1223) );
NOR2xp33_ASAP7_75t_L g1239 ( .A(n_1240), .B(n_1241), .Y(n_1239) );
NOR5xp2_ASAP7_75t_L g1242 ( .A(n_1243), .B(n_1247), .C(n_1254), .D(n_1261), .E(n_1263), .Y(n_1242) );
INVx1_ASAP7_75t_L g1257 ( .A(n_1258), .Y(n_1257) );
INVx4_ASAP7_75t_L g1266 ( .A(n_1267), .Y(n_1266) );
HB1xp67_ASAP7_75t_L g1268 ( .A(n_1269), .Y(n_1268) );
INVx1_ASAP7_75t_L g1269 ( .A(n_1270), .Y(n_1269) );
INVx1_ASAP7_75t_L g1270 ( .A(n_1271), .Y(n_1270) );
XNOR2xp5_ASAP7_75t_L g1271 ( .A(n_1272), .B(n_1315), .Y(n_1271) );
NAND2xp5_ASAP7_75t_SL g1272 ( .A(n_1273), .B(n_1308), .Y(n_1272) );
AOI21xp5_ASAP7_75t_L g1349 ( .A1(n_1274), .A2(n_1350), .B(n_1351), .Y(n_1349) );
NAND3xp33_ASAP7_75t_L g1276 ( .A(n_1277), .B(n_1281), .C(n_1286), .Y(n_1276) );
INVx1_ASAP7_75t_L g1296 ( .A(n_1297), .Y(n_1296) );
INVxp67_ASAP7_75t_SL g1297 ( .A(n_1298), .Y(n_1297) );
OAI22xp33_ASAP7_75t_L g1358 ( .A1(n_1298), .A2(n_1359), .B1(n_1360), .B2(n_1361), .Y(n_1358) );
OAI221xp5_ASAP7_75t_L g1300 ( .A1(n_1301), .A2(n_1302), .B1(n_1303), .B2(n_1304), .C(n_1305), .Y(n_1300) );
INVx1_ASAP7_75t_L g1306 ( .A(n_1307), .Y(n_1306) );
NAND3xp33_ASAP7_75t_L g1310 ( .A(n_1311), .B(n_1313), .C(n_1314), .Y(n_1310) );
CKINVDCx20_ASAP7_75t_R g1316 ( .A(n_1317), .Y(n_1316) );
CKINVDCx20_ASAP7_75t_R g1317 ( .A(n_1318), .Y(n_1317) );
INVx3_ASAP7_75t_L g1318 ( .A(n_1319), .Y(n_1318) );
HB1xp67_ASAP7_75t_L g1323 ( .A(n_1324), .Y(n_1323) );
INVxp33_ASAP7_75t_SL g1325 ( .A(n_1326), .Y(n_1325) );
INVx1_ASAP7_75t_L g1327 ( .A(n_1328), .Y(n_1327) );
NOR3xp33_ASAP7_75t_L g1328 ( .A(n_1329), .B(n_1372), .C(n_1377), .Y(n_1328) );
NAND2xp5_ASAP7_75t_L g1329 ( .A(n_1330), .B(n_1349), .Y(n_1329) );
NAND2xp5_ASAP7_75t_L g1332 ( .A(n_1333), .B(n_1336), .Y(n_1332) );
INVx1_ASAP7_75t_L g1334 ( .A(n_1335), .Y(n_1334) );
NAND3xp33_ASAP7_75t_L g1339 ( .A(n_1340), .B(n_1344), .C(n_1347), .Y(n_1339) );
OAI22xp5_ASAP7_75t_L g1352 ( .A1(n_1353), .A2(n_1354), .B1(n_1355), .B2(n_1356), .Y(n_1352) );
INVx1_ASAP7_75t_L g1356 ( .A(n_1357), .Y(n_1356) );
INVx1_ASAP7_75t_L g1361 ( .A(n_1362), .Y(n_1361) );
OAI22xp5_ASAP7_75t_L g1366 ( .A1(n_1367), .A2(n_1368), .B1(n_1369), .B2(n_1371), .Y(n_1366) );
INVx1_ASAP7_75t_L g1369 ( .A(n_1370), .Y(n_1369) );
INVx1_ASAP7_75t_L g1380 ( .A(n_1381), .Y(n_1380) );
endmodule