module fake_netlist_5_1216_n_2682 (n_137, n_294, n_431, n_318, n_380, n_419, n_444, n_469, n_82, n_194, n_316, n_389, n_418, n_248, n_124, n_86, n_136, n_146, n_315, n_268, n_451, n_408, n_61, n_376, n_127, n_75, n_235, n_226, n_74, n_57, n_353, n_351, n_367, n_452, n_397, n_111, n_155, n_43, n_116, n_22, n_467, n_423, n_284, n_46, n_245, n_21, n_139, n_38, n_105, n_280, n_4, n_378, n_17, n_382, n_254, n_33, n_23, n_302, n_265, n_293, n_372, n_443, n_244, n_47, n_173, n_198, n_447, n_247, n_314, n_368, n_433, n_8, n_321, n_292, n_100, n_455, n_417, n_212, n_385, n_119, n_275, n_252, n_26, n_295, n_133, n_330, n_2, n_6, n_39, n_147, n_373, n_67, n_307, n_439, n_87, n_150, n_106, n_209, n_259, n_448, n_375, n_301, n_68, n_93, n_186, n_134, n_191, n_51, n_63, n_171, n_153, n_399, n_341, n_204, n_394, n_250, n_260, n_298, n_320, n_286, n_122, n_282, n_331, n_10, n_24, n_406, n_325, n_449, n_132, n_90, n_101, n_281, n_240, n_381, n_189, n_220, n_291, n_231, n_257, n_390, n_31, n_456, n_13, n_371, n_152, n_317, n_9, n_323, n_195, n_42, n_356, n_227, n_45, n_271, n_94, n_335, n_123, n_370, n_167, n_234, n_343, n_308, n_379, n_428, n_267, n_457, n_297, n_156, n_5, n_225, n_377, n_219, n_442, n_157, n_131, n_192, n_223, n_392, n_158, n_138, n_264, n_109, n_454, n_387, n_374, n_163, n_276, n_339, n_95, n_183, n_185, n_243, n_398, n_396, n_347, n_169, n_59, n_255, n_215, n_350, n_196, n_459, n_211, n_218, n_400, n_181, n_436, n_3, n_290, n_221, n_178, n_386, n_287, n_344, n_422, n_72, n_104, n_41, n_415, n_56, n_141, n_355, n_15, n_336, n_145, n_48, n_50, n_337, n_430, n_313, n_88, n_216, n_168, n_395, n_164, n_432, n_311, n_208, n_142, n_214, n_328, n_140, n_299, n_303, n_369, n_296, n_241, n_357, n_184, n_446, n_445, n_65, n_78, n_144, n_114, n_96, n_165, n_468, n_213, n_129, n_342, n_98, n_361, n_464, n_363, n_402, n_413, n_197, n_107, n_69, n_236, n_388, n_1, n_249, n_304, n_329, n_203, n_274, n_384, n_460, n_80, n_35, n_73, n_277, n_92, n_19, n_338, n_149, n_461, n_333, n_309, n_30, n_14, n_84, n_462, n_130, n_322, n_258, n_29, n_79, n_151, n_25, n_306, n_458, n_288, n_188, n_190, n_201, n_263, n_44, n_224, n_40, n_34, n_228, n_283, n_383, n_112, n_85, n_463, n_239, n_466, n_420, n_55, n_49, n_310, n_54, n_12, n_465, n_76, n_358, n_362, n_170, n_332, n_27, n_77, n_102, n_161, n_273, n_349, n_270, n_230, n_81, n_118, n_279, n_70, n_253, n_261, n_174, n_289, n_172, n_206, n_217, n_440, n_441, n_450, n_312, n_429, n_345, n_210, n_365, n_91, n_176, n_182, n_143, n_83, n_354, n_237, n_425, n_407, n_180, n_340, n_207, n_37, n_346, n_393, n_229, n_108, n_437, n_66, n_177, n_60, n_403, n_453, n_421, n_16, n_0, n_58, n_405, n_18, n_359, n_117, n_326, n_233, n_404, n_205, n_366, n_113, n_246, n_179, n_125, n_410, n_269, n_128, n_285, n_412, n_120, n_232, n_327, n_135, n_126, n_202, n_266, n_272, n_427, n_193, n_251, n_352, n_53, n_160, n_426, n_409, n_154, n_62, n_148, n_71, n_300, n_435, n_159, n_334, n_391, n_434, n_175, n_262, n_238, n_99, n_411, n_414, n_319, n_364, n_20, n_121, n_242, n_360, n_36, n_200, n_162, n_64, n_222, n_28, n_89, n_438, n_115, n_324, n_416, n_199, n_187, n_32, n_401, n_103, n_348, n_97, n_166, n_11, n_424, n_7, n_256, n_305, n_52, n_278, n_110, n_2682);

input n_137;
input n_294;
input n_431;
input n_318;
input n_380;
input n_419;
input n_444;
input n_469;
input n_82;
input n_194;
input n_316;
input n_389;
input n_418;
input n_248;
input n_124;
input n_86;
input n_136;
input n_146;
input n_315;
input n_268;
input n_451;
input n_408;
input n_61;
input n_376;
input n_127;
input n_75;
input n_235;
input n_226;
input n_74;
input n_57;
input n_353;
input n_351;
input n_367;
input n_452;
input n_397;
input n_111;
input n_155;
input n_43;
input n_116;
input n_22;
input n_467;
input n_423;
input n_284;
input n_46;
input n_245;
input n_21;
input n_139;
input n_38;
input n_105;
input n_280;
input n_4;
input n_378;
input n_17;
input n_382;
input n_254;
input n_33;
input n_23;
input n_302;
input n_265;
input n_293;
input n_372;
input n_443;
input n_244;
input n_47;
input n_173;
input n_198;
input n_447;
input n_247;
input n_314;
input n_368;
input n_433;
input n_8;
input n_321;
input n_292;
input n_100;
input n_455;
input n_417;
input n_212;
input n_385;
input n_119;
input n_275;
input n_252;
input n_26;
input n_295;
input n_133;
input n_330;
input n_2;
input n_6;
input n_39;
input n_147;
input n_373;
input n_67;
input n_307;
input n_439;
input n_87;
input n_150;
input n_106;
input n_209;
input n_259;
input n_448;
input n_375;
input n_301;
input n_68;
input n_93;
input n_186;
input n_134;
input n_191;
input n_51;
input n_63;
input n_171;
input n_153;
input n_399;
input n_341;
input n_204;
input n_394;
input n_250;
input n_260;
input n_298;
input n_320;
input n_286;
input n_122;
input n_282;
input n_331;
input n_10;
input n_24;
input n_406;
input n_325;
input n_449;
input n_132;
input n_90;
input n_101;
input n_281;
input n_240;
input n_381;
input n_189;
input n_220;
input n_291;
input n_231;
input n_257;
input n_390;
input n_31;
input n_456;
input n_13;
input n_371;
input n_152;
input n_317;
input n_9;
input n_323;
input n_195;
input n_42;
input n_356;
input n_227;
input n_45;
input n_271;
input n_94;
input n_335;
input n_123;
input n_370;
input n_167;
input n_234;
input n_343;
input n_308;
input n_379;
input n_428;
input n_267;
input n_457;
input n_297;
input n_156;
input n_5;
input n_225;
input n_377;
input n_219;
input n_442;
input n_157;
input n_131;
input n_192;
input n_223;
input n_392;
input n_158;
input n_138;
input n_264;
input n_109;
input n_454;
input n_387;
input n_374;
input n_163;
input n_276;
input n_339;
input n_95;
input n_183;
input n_185;
input n_243;
input n_398;
input n_396;
input n_347;
input n_169;
input n_59;
input n_255;
input n_215;
input n_350;
input n_196;
input n_459;
input n_211;
input n_218;
input n_400;
input n_181;
input n_436;
input n_3;
input n_290;
input n_221;
input n_178;
input n_386;
input n_287;
input n_344;
input n_422;
input n_72;
input n_104;
input n_41;
input n_415;
input n_56;
input n_141;
input n_355;
input n_15;
input n_336;
input n_145;
input n_48;
input n_50;
input n_337;
input n_430;
input n_313;
input n_88;
input n_216;
input n_168;
input n_395;
input n_164;
input n_432;
input n_311;
input n_208;
input n_142;
input n_214;
input n_328;
input n_140;
input n_299;
input n_303;
input n_369;
input n_296;
input n_241;
input n_357;
input n_184;
input n_446;
input n_445;
input n_65;
input n_78;
input n_144;
input n_114;
input n_96;
input n_165;
input n_468;
input n_213;
input n_129;
input n_342;
input n_98;
input n_361;
input n_464;
input n_363;
input n_402;
input n_413;
input n_197;
input n_107;
input n_69;
input n_236;
input n_388;
input n_1;
input n_249;
input n_304;
input n_329;
input n_203;
input n_274;
input n_384;
input n_460;
input n_80;
input n_35;
input n_73;
input n_277;
input n_92;
input n_19;
input n_338;
input n_149;
input n_461;
input n_333;
input n_309;
input n_30;
input n_14;
input n_84;
input n_462;
input n_130;
input n_322;
input n_258;
input n_29;
input n_79;
input n_151;
input n_25;
input n_306;
input n_458;
input n_288;
input n_188;
input n_190;
input n_201;
input n_263;
input n_44;
input n_224;
input n_40;
input n_34;
input n_228;
input n_283;
input n_383;
input n_112;
input n_85;
input n_463;
input n_239;
input n_466;
input n_420;
input n_55;
input n_49;
input n_310;
input n_54;
input n_12;
input n_465;
input n_76;
input n_358;
input n_362;
input n_170;
input n_332;
input n_27;
input n_77;
input n_102;
input n_161;
input n_273;
input n_349;
input n_270;
input n_230;
input n_81;
input n_118;
input n_279;
input n_70;
input n_253;
input n_261;
input n_174;
input n_289;
input n_172;
input n_206;
input n_217;
input n_440;
input n_441;
input n_450;
input n_312;
input n_429;
input n_345;
input n_210;
input n_365;
input n_91;
input n_176;
input n_182;
input n_143;
input n_83;
input n_354;
input n_237;
input n_425;
input n_407;
input n_180;
input n_340;
input n_207;
input n_37;
input n_346;
input n_393;
input n_229;
input n_108;
input n_437;
input n_66;
input n_177;
input n_60;
input n_403;
input n_453;
input n_421;
input n_16;
input n_0;
input n_58;
input n_405;
input n_18;
input n_359;
input n_117;
input n_326;
input n_233;
input n_404;
input n_205;
input n_366;
input n_113;
input n_246;
input n_179;
input n_125;
input n_410;
input n_269;
input n_128;
input n_285;
input n_412;
input n_120;
input n_232;
input n_327;
input n_135;
input n_126;
input n_202;
input n_266;
input n_272;
input n_427;
input n_193;
input n_251;
input n_352;
input n_53;
input n_160;
input n_426;
input n_409;
input n_154;
input n_62;
input n_148;
input n_71;
input n_300;
input n_435;
input n_159;
input n_334;
input n_391;
input n_434;
input n_175;
input n_262;
input n_238;
input n_99;
input n_411;
input n_414;
input n_319;
input n_364;
input n_20;
input n_121;
input n_242;
input n_360;
input n_36;
input n_200;
input n_162;
input n_64;
input n_222;
input n_28;
input n_89;
input n_438;
input n_115;
input n_324;
input n_416;
input n_199;
input n_187;
input n_32;
input n_401;
input n_103;
input n_348;
input n_97;
input n_166;
input n_11;
input n_424;
input n_7;
input n_256;
input n_305;
input n_52;
input n_278;
input n_110;

output n_2682;

wire n_924;
wire n_1263;
wire n_977;
wire n_1378;
wire n_2253;
wire n_2417;
wire n_611;
wire n_1126;
wire n_1423;
wire n_1729;
wire n_1166;
wire n_2380;
wire n_1751;
wire n_1508;
wire n_785;
wire n_549;
wire n_2617;
wire n_2200;
wire n_532;
wire n_1161;
wire n_1859;
wire n_1677;
wire n_1150;
wire n_2327;
wire n_1780;
wire n_1488;
wire n_667;
wire n_790;
wire n_1055;
wire n_2386;
wire n_1501;
wire n_2395;
wire n_880;
wire n_544;
wire n_1007;
wire n_2369;
wire n_552;
wire n_1528;
wire n_1370;
wire n_1292;
wire n_2347;
wire n_2520;
wire n_1198;
wire n_1360;
wire n_2388;
wire n_1099;
wire n_2568;
wire n_956;
wire n_564;
wire n_1738;
wire n_2021;
wire n_2134;
wire n_2391;
wire n_1021;
wire n_1960;
wire n_2185;
wire n_551;
wire n_2143;
wire n_2059;
wire n_1323;
wire n_1466;
wire n_688;
wire n_1695;
wire n_2487;
wire n_1353;
wire n_800;
wire n_1347;
wire n_2495;
wire n_1535;
wire n_1789;
wire n_1666;
wire n_2389;
wire n_671;
wire n_819;
wire n_1451;
wire n_1022;
wire n_2302;
wire n_915;
wire n_1545;
wire n_2374;
wire n_864;
wire n_859;
wire n_951;
wire n_1947;
wire n_1264;
wire n_2114;
wire n_2001;
wire n_1494;
wire n_625;
wire n_854;
wire n_1462;
wire n_1799;
wire n_2069;
wire n_2396;
wire n_1580;
wire n_674;
wire n_1939;
wire n_2486;
wire n_1806;
wire n_516;
wire n_933;
wire n_2244;
wire n_2257;
wire n_1152;
wire n_497;
wire n_1869;
wire n_1607;
wire n_1563;
wire n_606;
wire n_2011;
wire n_2096;
wire n_877;
wire n_2105;
wire n_2538;
wire n_2024;
wire n_2530;
wire n_1696;
wire n_2483;
wire n_755;
wire n_1118;
wire n_1686;
wire n_947;
wire n_1285;
wire n_1860;
wire n_2543;
wire n_1359;
wire n_530;
wire n_1728;
wire n_1107;
wire n_2076;
wire n_2031;
wire n_556;
wire n_2482;
wire n_2677;
wire n_1230;
wire n_668;
wire n_1896;
wire n_2165;
wire n_2147;
wire n_929;
wire n_1124;
wire n_1818;
wire n_2127;
wire n_1576;
wire n_902;
wire n_1104;
wire n_1294;
wire n_659;
wire n_1705;
wire n_2584;
wire n_1257;
wire n_2639;
wire n_1182;
wire n_579;
wire n_1698;
wire n_1261;
wire n_2329;
wire n_938;
wire n_1098;
wire n_2142;
wire n_1154;
wire n_2189;
wire n_1242;
wire n_1135;
wire n_519;
wire n_2323;
wire n_2203;
wire n_2597;
wire n_1016;
wire n_1243;
wire n_546;
wire n_2047;
wire n_1280;
wire n_1845;
wire n_2052;
wire n_2193;
wire n_2058;
wire n_2458;
wire n_2478;
wire n_731;
wire n_1483;
wire n_1314;
wire n_1512;
wire n_709;
wire n_1490;
wire n_1236;
wire n_1633;
wire n_2537;
wire n_569;
wire n_2669;
wire n_2144;
wire n_1778;
wire n_2306;
wire n_920;
wire n_2515;
wire n_1289;
wire n_1517;
wire n_2091;
wire n_2466;
wire n_2635;
wire n_2652;
wire n_2085;
wire n_1669;
wire n_2566;
wire n_976;
wire n_1949;
wire n_1449;
wire n_1946;
wire n_1566;
wire n_2032;
wire n_2587;
wire n_2149;
wire n_1078;
wire n_1670;
wire n_2672;
wire n_775;
wire n_2651;
wire n_600;
wire n_1484;
wire n_2071;
wire n_2561;
wire n_1374;
wire n_1328;
wire n_2643;
wire n_2141;
wire n_1948;
wire n_1984;
wire n_2099;
wire n_2408;
wire n_1877;
wire n_1831;
wire n_1598;
wire n_1723;
wire n_955;
wire n_1850;
wire n_1146;
wire n_882;
wire n_2384;
wire n_1097;
wire n_1749;
wire n_1036;
wire n_696;
wire n_550;
wire n_897;
wire n_798;
wire n_646;
wire n_1428;
wire n_2663;
wire n_1394;
wire n_2659;
wire n_1414;
wire n_1216;
wire n_580;
wire n_1040;
wire n_2202;
wire n_2648;
wire n_1872;
wire n_1852;
wire n_2159;
wire n_578;
wire n_926;
wire n_2180;
wire n_2249;
wire n_2353;
wire n_2439;
wire n_1931;
wire n_1218;
wire n_2632;
wire n_2276;
wire n_475;
wire n_1070;
wire n_1547;
wire n_777;
wire n_2089;
wire n_1030;
wire n_2470;
wire n_1755;
wire n_1561;
wire n_1071;
wire n_485;
wire n_1165;
wire n_1267;
wire n_496;
wire n_1801;
wire n_1391;
wire n_958;
wire n_1034;
wire n_670;
wire n_1513;
wire n_1600;
wire n_521;
wire n_663;
wire n_845;
wire n_2235;
wire n_1862;
wire n_673;
wire n_837;
wire n_1239;
wire n_528;
wire n_2300;
wire n_1796;
wire n_2551;
wire n_1587;
wire n_680;
wire n_1473;
wire n_553;
wire n_901;
wire n_2432;
wire n_813;
wire n_1521;
wire n_1284;
wire n_1590;
wire n_2174;
wire n_1748;
wire n_1672;
wire n_2506;
wire n_675;
wire n_1880;
wire n_888;
wire n_2337;
wire n_1167;
wire n_1626;
wire n_637;
wire n_2615;
wire n_1384;
wire n_1556;
wire n_1863;
wire n_1064;
wire n_858;
wire n_2079;
wire n_2238;
wire n_923;
wire n_2118;
wire n_691;
wire n_1151;
wire n_881;
wire n_1405;
wire n_2407;
wire n_1706;
wire n_1582;
wire n_1069;
wire n_1784;
wire n_1075;
wire n_1836;
wire n_1450;
wire n_1322;
wire n_2101;
wire n_1471;
wire n_1986;
wire n_2072;
wire n_1750;
wire n_1459;
wire n_889;
wire n_2358;
wire n_973;
wire n_1700;
wire n_477;
wire n_571;
wire n_1585;
wire n_1971;
wire n_1599;
wire n_2275;
wire n_2644;
wire n_1211;
wire n_1197;
wire n_1523;
wire n_1950;
wire n_1447;
wire n_907;
wire n_2251;
wire n_1377;
wire n_2370;
wire n_989;
wire n_2544;
wire n_1039;
wire n_2214;
wire n_2055;
wire n_1403;
wire n_2248;
wire n_2356;
wire n_488;
wire n_736;
wire n_892;
wire n_1000;
wire n_1202;
wire n_2620;
wire n_1278;
wire n_2622;
wire n_2062;
wire n_2668;
wire n_1002;
wire n_1463;
wire n_1581;
wire n_2100;
wire n_593;
wire n_2258;
wire n_748;
wire n_1058;
wire n_586;
wire n_1667;
wire n_838;
wire n_1053;
wire n_1224;
wire n_2557;
wire n_1926;
wire n_1248;
wire n_1331;
wire n_953;
wire n_1014;
wire n_1241;
wire n_2150;
wire n_2241;
wire n_2152;
wire n_963;
wire n_1052;
wire n_954;
wire n_627;
wire n_1385;
wire n_793;
wire n_478;
wire n_2590;
wire n_2140;
wire n_2385;
wire n_1819;
wire n_2330;
wire n_2139;
wire n_476;
wire n_1527;
wire n_2042;
wire n_534;
wire n_1882;
wire n_884;
wire n_944;
wire n_1754;
wire n_1623;
wire n_2175;
wire n_2324;
wire n_1854;
wire n_2606;
wire n_2674;
wire n_1565;
wire n_1809;
wire n_1856;
wire n_647;
wire n_1072;
wire n_2218;
wire n_2267;
wire n_857;
wire n_832;
wire n_2305;
wire n_2636;
wire n_2450;
wire n_561;
wire n_1319;
wire n_2379;
wire n_2616;
wire n_2154;
wire n_1825;
wire n_1951;
wire n_1883;
wire n_1906;
wire n_1712;
wire n_1387;
wire n_2262;
wire n_2462;
wire n_2514;
wire n_1532;
wire n_2322;
wire n_2271;
wire n_2625;
wire n_1027;
wire n_971;
wire n_1156;
wire n_794;
wire n_2331;
wire n_2293;
wire n_686;
wire n_847;
wire n_1393;
wire n_2319;
wire n_596;
wire n_1775;
wire n_2028;
wire n_1368;
wire n_558;
wire n_702;
wire n_1276;
wire n_2548;
wire n_1412;
wire n_822;
wire n_2676;
wire n_1709;
wire n_2679;
wire n_2108;
wire n_728;
wire n_1162;
wire n_1538;
wire n_1838;
wire n_1847;
wire n_1199;
wire n_1779;
wire n_2603;
wire n_1884;
wire n_2434;
wire n_2660;
wire n_1038;
wire n_1369;
wire n_520;
wire n_2611;
wire n_1841;
wire n_1660;
wire n_887;
wire n_1905;
wire n_2553;
wire n_2581;
wire n_2195;
wire n_2529;
wire n_809;
wire n_931;
wire n_1711;
wire n_599;
wire n_870;
wire n_1662;
wire n_1891;
wire n_1481;
wire n_2626;
wire n_1942;
wire n_1978;
wire n_1544;
wire n_2510;
wire n_868;
wire n_2454;
wire n_639;
wire n_914;
wire n_2120;
wire n_2546;
wire n_1629;
wire n_1293;
wire n_965;
wire n_1876;
wire n_1743;
wire n_935;
wire n_817;
wire n_1175;
wire n_1479;
wire n_1810;
wire n_2350;
wire n_1888;
wire n_2009;
wire n_759;
wire n_2222;
wire n_1892;
wire n_806;
wire n_1997;
wire n_2667;
wire n_1766;
wire n_1477;
wire n_1635;
wire n_1963;
wire n_2226;
wire n_1571;
wire n_1189;
wire n_2215;
wire n_1259;
wire n_1690;
wire n_706;
wire n_746;
wire n_1649;
wire n_747;
wire n_2064;
wire n_784;
wire n_2449;
wire n_1733;
wire n_1244;
wire n_2413;
wire n_1194;
wire n_1925;
wire n_2297;
wire n_1815;
wire n_2621;
wire n_851;
wire n_615;
wire n_1759;
wire n_843;
wire n_1788;
wire n_2177;
wire n_2491;
wire n_523;
wire n_913;
wire n_1537;
wire n_705;
wire n_865;
wire n_2227;
wire n_678;
wire n_2671;
wire n_697;
wire n_1222;
wire n_1679;
wire n_2190;
wire n_1798;
wire n_2022;
wire n_776;
wire n_1790;
wire n_2518;
wire n_1415;
wire n_2629;
wire n_2592;
wire n_525;
wire n_1260;
wire n_1746;
wire n_1647;
wire n_2181;
wire n_2479;
wire n_1829;
wire n_1464;
wire n_649;
wire n_547;
wire n_2563;
wire n_1444;
wire n_1191;
wire n_2387;
wire n_1674;
wire n_1833;
wire n_1830;
wire n_2517;
wire n_2073;
wire n_1710;
wire n_1128;
wire n_1734;
wire n_744;
wire n_590;
wire n_629;
wire n_2631;
wire n_1308;
wire n_2178;
wire n_1767;
wire n_2336;
wire n_1680;
wire n_1233;
wire n_2607;
wire n_1615;
wire n_1529;
wire n_2005;
wire n_526;
wire n_1916;
wire n_677;
wire n_1333;
wire n_2469;
wire n_1121;
wire n_604;
wire n_2007;
wire n_949;
wire n_2539;
wire n_2582;
wire n_1443;
wire n_1008;
wire n_946;
wire n_1539;
wire n_1001;
wire n_1503;
wire n_2054;
wire n_498;
wire n_1468;
wire n_1559;
wire n_1765;
wire n_1866;
wire n_689;
wire n_738;
wire n_1624;
wire n_640;
wire n_1510;
wire n_624;
wire n_1380;
wire n_1744;
wire n_2623;
wire n_1617;
wire n_1010;
wire n_1994;
wire n_1231;
wire n_739;
wire n_1279;
wire n_1406;
wire n_1195;
wire n_1839;
wire n_1837;
wire n_610;
wire n_2577;
wire n_1760;
wire n_936;
wire n_568;
wire n_1500;
wire n_1090;
wire n_757;
wire n_2342;
wire n_633;
wire n_1832;
wire n_1851;
wire n_758;
wire n_999;
wire n_2046;
wire n_1933;
wire n_2290;
wire n_1656;
wire n_1158;
wire n_2045;
wire n_1509;
wire n_1874;
wire n_2040;
wire n_563;
wire n_2060;
wire n_2613;
wire n_1987;
wire n_1145;
wire n_878;
wire n_524;
wire n_1678;
wire n_1049;
wire n_1153;
wire n_2145;
wire n_741;
wire n_1639;
wire n_1306;
wire n_1068;
wire n_1871;
wire n_2580;
wire n_2545;
wire n_1964;
wire n_1163;
wire n_906;
wire n_2039;
wire n_1207;
wire n_919;
wire n_908;
wire n_2412;
wire n_2406;
wire n_724;
wire n_1781;
wire n_2084;
wire n_2035;
wire n_658;
wire n_2061;
wire n_2378;
wire n_2509;
wire n_1740;
wire n_2398;
wire n_1362;
wire n_1586;
wire n_959;
wire n_2459;
wire n_535;
wire n_940;
wire n_1445;
wire n_1492;
wire n_2155;
wire n_2516;
wire n_1923;
wire n_1773;
wire n_592;
wire n_1169;
wire n_1596;
wire n_1692;
wire n_2666;
wire n_1017;
wire n_2481;
wire n_2171;
wire n_978;
wire n_2116;
wire n_2314;
wire n_1434;
wire n_1054;
wire n_2507;
wire n_1474;
wire n_1665;
wire n_1269;
wire n_2420;
wire n_1095;
wire n_1828;
wire n_1614;
wire n_1079;
wire n_2093;
wire n_514;
wire n_1045;
wire n_1208;
wire n_2339;
wire n_2038;
wire n_2320;
wire n_2473;
wire n_2137;
wire n_603;
wire n_1431;
wire n_2583;
wire n_484;
wire n_1593;
wire n_1033;
wire n_2299;
wire n_2540;
wire n_636;
wire n_660;
wire n_2087;
wire n_1640;
wire n_2162;
wire n_1732;
wire n_1009;
wire n_1148;
wire n_2051;
wire n_742;
wire n_2029;
wire n_750;
wire n_995;
wire n_2168;
wire n_1609;
wire n_1989;
wire n_2359;
wire n_1887;
wire n_2523;
wire n_1383;
wire n_1073;
wire n_2346;
wire n_2457;
wire n_662;
wire n_2312;
wire n_962;
wire n_1215;
wire n_1171;
wire n_1578;
wire n_723;
wire n_1920;
wire n_1065;
wire n_1592;
wire n_2536;
wire n_1336;
wire n_1721;
wire n_1959;
wire n_1758;
wire n_2338;
wire n_1574;
wire n_2399;
wire n_473;
wire n_2048;
wire n_2355;
wire n_2133;
wire n_1921;
wire n_1309;
wire n_1878;
wire n_1426;
wire n_1043;
wire n_2585;
wire n_486;
wire n_1800;
wire n_1548;
wire n_614;
wire n_1421;
wire n_2571;
wire n_1286;
wire n_1177;
wire n_1355;
wire n_974;
wire n_2565;
wire n_727;
wire n_1159;
wire n_957;
wire n_773;
wire n_2124;
wire n_743;
wire n_2081;
wire n_613;
wire n_1119;
wire n_2156;
wire n_2261;
wire n_1240;
wire n_1820;
wire n_2418;
wire n_829;
wire n_2519;
wire n_1612;
wire n_2179;
wire n_1416;
wire n_2077;
wire n_1724;
wire n_2111;
wire n_2521;
wire n_700;
wire n_1237;
wire n_573;
wire n_1420;
wire n_1132;
wire n_1366;
wire n_1300;
wire n_2595;
wire n_1127;
wire n_2277;
wire n_761;
wire n_2477;
wire n_1785;
wire n_1568;
wire n_1006;
wire n_2110;
wire n_1270;
wire n_1664;
wire n_1486;
wire n_582;
wire n_1332;
wire n_2231;
wire n_1390;
wire n_2017;
wire n_2474;
wire n_2604;
wire n_2090;
wire n_1870;
wire n_2367;
wire n_512;
wire n_1591;
wire n_2033;
wire n_1682;
wire n_1980;
wire n_2390;
wire n_2628;
wire n_1249;
wire n_652;
wire n_1111;
wire n_1365;
wire n_1927;
wire n_2132;
wire n_1349;
wire n_1093;
wire n_2400;
wire n_1031;
wire n_609;
wire n_1041;
wire n_1265;
wire n_1909;
wire n_2681;
wire n_1562;
wire n_834;
wire n_765;
wire n_2255;
wire n_2424;
wire n_2272;
wire n_893;
wire n_1015;
wire n_1140;
wire n_891;
wire n_1651;
wire n_1965;
wire n_630;
wire n_1902;
wire n_2151;
wire n_1941;
wire n_2106;
wire n_1913;
wire n_504;
wire n_1823;
wire n_511;
wire n_874;
wire n_2464;
wire n_1101;
wire n_1106;
wire n_1456;
wire n_2230;
wire n_2015;
wire n_2365;
wire n_1875;
wire n_1982;
wire n_1304;
wire n_1324;
wire n_987;
wire n_1846;
wire n_2066;
wire n_1885;
wire n_1455;
wire n_767;
wire n_993;
wire n_1903;
wire n_2490;
wire n_1407;
wire n_2452;
wire n_1551;
wire n_545;
wire n_860;
wire n_1805;
wire n_2176;
wire n_2204;
wire n_1816;
wire n_948;
wire n_1217;
wire n_2220;
wire n_2455;
wire n_628;
wire n_1849;
wire n_2410;
wire n_729;
wire n_1131;
wire n_1084;
wire n_1961;
wire n_970;
wire n_1935;
wire n_911;
wire n_1430;
wire n_2645;
wire n_2467;
wire n_513;
wire n_1094;
wire n_1354;
wire n_560;
wire n_1534;
wire n_2288;
wire n_1351;
wire n_2240;
wire n_1205;
wire n_1044;
wire n_2436;
wire n_1209;
wire n_1552;
wire n_2508;
wire n_495;
wire n_602;
wire n_574;
wire n_2593;
wire n_1435;
wire n_879;
wire n_2416;
wire n_2405;
wire n_623;
wire n_2088;
wire n_824;
wire n_1645;
wire n_2461;
wire n_490;
wire n_1327;
wire n_2243;
wire n_996;
wire n_1684;
wire n_921;
wire n_2658;
wire n_1717;
wire n_572;
wire n_815;
wire n_1795;
wire n_2128;
wire n_2578;
wire n_1821;
wire n_1381;
wire n_2555;
wire n_2662;
wire n_1611;
wire n_1037;
wire n_2368;
wire n_2656;
wire n_1080;
wire n_2301;
wire n_1274;
wire n_2554;
wire n_1316;
wire n_1708;
wire n_2419;
wire n_1438;
wire n_1082;
wire n_1840;
wire n_589;
wire n_1630;
wire n_716;
wire n_2122;
wire n_2512;
wire n_562;
wire n_1436;
wire n_1691;
wire n_952;
wire n_2534;
wire n_2092;
wire n_1229;
wire n_701;
wire n_1437;
wire n_1023;
wire n_2075;
wire n_645;
wire n_539;
wire n_803;
wire n_1092;
wire n_1776;
wire n_2198;
wire n_2610;
wire n_2661;
wire n_2572;
wire n_2281;
wire n_2131;
wire n_2216;
wire n_531;
wire n_1757;
wire n_890;
wire n_1897;
wire n_764;
wire n_1919;
wire n_1056;
wire n_1424;
wire n_960;
wire n_2308;
wire n_1893;
wire n_1290;
wire n_1123;
wire n_1467;
wire n_1047;
wire n_2053;
wire n_2163;
wire n_634;
wire n_2328;
wire n_1958;
wire n_2254;
wire n_1252;
wire n_1382;
wire n_1029;
wire n_925;
wire n_1206;
wire n_2647;
wire n_1311;
wire n_2191;
wire n_1519;
wire n_950;
wire n_2428;
wire n_1553;
wire n_2664;
wire n_1811;
wire n_2443;
wire n_2624;
wire n_1346;
wire n_1299;
wire n_2158;
wire n_1808;
wire n_1060;
wire n_1141;
wire n_2266;
wire n_2465;
wire n_2650;
wire n_912;
wire n_968;
wire n_619;
wire n_2440;
wire n_1386;
wire n_1699;
wire n_967;
wire n_1442;
wire n_2541;
wire n_1139;
wire n_515;
wire n_2333;
wire n_885;
wire n_1432;
wire n_1357;
wire n_483;
wire n_2125;
wire n_683;
wire n_1632;
wire n_1057;
wire n_1051;
wire n_1085;
wire n_1066;
wire n_721;
wire n_2402;
wire n_1157;
wire n_2403;
wire n_841;
wire n_1050;
wire n_802;
wire n_1954;
wire n_2265;
wire n_1608;
wire n_983;
wire n_1844;
wire n_1305;
wire n_873;
wire n_1826;
wire n_1112;
wire n_2304;
wire n_762;
wire n_1283;
wire n_1644;
wire n_2334;
wire n_2637;
wire n_690;
wire n_1974;
wire n_2463;
wire n_583;
wire n_2086;
wire n_2289;
wire n_1343;
wire n_2263;
wire n_1631;
wire n_1203;
wire n_2472;
wire n_821;
wire n_1763;
wire n_2341;
wire n_1966;
wire n_1768;
wire n_2294;
wire n_1179;
wire n_621;
wire n_753;
wire n_2475;
wire n_1048;
wire n_1719;
wire n_1288;
wire n_2556;
wire n_507;
wire n_2269;
wire n_2309;
wire n_2415;
wire n_2646;
wire n_1560;
wire n_1605;
wire n_2236;
wire n_1228;
wire n_2123;
wire n_972;
wire n_692;
wire n_2037;
wire n_1953;
wire n_1938;
wire n_820;
wire n_1200;
wire n_2499;
wire n_1911;
wire n_2460;
wire n_2589;
wire n_1363;
wire n_1668;
wire n_1301;
wire n_1185;
wire n_991;
wire n_828;
wire n_1967;
wire n_779;
wire n_576;
wire n_1143;
wire n_1579;
wire n_2233;
wire n_1329;
wire n_2675;
wire n_1312;
wire n_1439;
wire n_804;
wire n_537;
wire n_1688;
wire n_945;
wire n_492;
wire n_1504;
wire n_943;
wire n_992;
wire n_1932;
wire n_543;
wire n_842;
wire n_650;
wire n_984;
wire n_694;
wire n_2082;
wire n_1992;
wire n_2429;
wire n_1643;
wire n_883;
wire n_1983;
wire n_470;
wire n_1594;
wire n_1214;
wire n_1400;
wire n_1342;
wire n_900;
wire n_2362;
wire n_856;
wire n_2609;
wire n_1793;
wire n_1976;
wire n_2223;
wire n_918;
wire n_942;
wire n_2169;
wire n_1804;
wire n_1147;
wire n_1557;
wire n_1977;
wire n_2153;
wire n_2468;
wire n_1610;
wire n_1077;
wire n_1422;
wire n_2364;
wire n_2533;
wire n_540;
wire n_618;
wire n_896;
wire n_2310;
wire n_2287;
wire n_2291;
wire n_2596;
wire n_894;
wire n_1636;
wire n_2056;
wire n_1730;
wire n_831;
wire n_2280;
wire n_2192;
wire n_964;
wire n_1373;
wire n_1350;
wire n_1511;
wire n_1865;
wire n_1470;
wire n_1096;
wire n_2094;
wire n_2670;
wire n_1575;
wire n_1735;
wire n_2318;
wire n_2393;
wire n_833;
wire n_1697;
wire n_2020;
wire n_1646;
wire n_2502;
wire n_2504;
wire n_1307;
wire n_1881;
wire n_988;
wire n_2043;
wire n_1940;
wire n_814;
wire n_1549;
wire n_1934;
wire n_2311;
wire n_1201;
wire n_1114;
wire n_655;
wire n_2025;
wire n_1616;
wire n_1446;
wire n_2285;
wire n_669;
wire n_472;
wire n_1458;
wire n_1176;
wire n_1472;
wire n_2298;
wire n_2471;
wire n_1807;
wire n_1149;
wire n_2618;
wire n_1671;
wire n_635;
wire n_2559;
wire n_763;
wire n_1020;
wire n_1062;
wire n_2303;
wire n_1824;
wire n_1917;
wire n_2295;
wire n_1219;
wire n_1204;
wire n_2325;
wire n_2446;
wire n_1814;
wire n_1035;
wire n_555;
wire n_1848;
wire n_1928;
wire n_783;
wire n_2126;
wire n_1188;
wire n_2588;
wire n_1722;
wire n_661;
wire n_2441;
wire n_1802;
wire n_2600;
wire n_849;
wire n_584;
wire n_681;
wire n_1638;
wire n_1786;
wire n_2002;
wire n_2282;
wire n_510;
wire n_2371;
wire n_830;
wire n_2098;
wire n_1296;
wire n_2627;
wire n_2352;
wire n_1413;
wire n_801;
wire n_2207;
wire n_2080;
wire n_2377;
wire n_2619;
wire n_2340;
wire n_2444;
wire n_2068;
wire n_875;
wire n_1110;
wire n_1655;
wire n_2641;
wire n_749;
wire n_1895;
wire n_2574;
wire n_1134;
wire n_1358;
wire n_717;
wire n_939;
wire n_482;
wire n_2361;
wire n_1088;
wire n_588;
wire n_1173;
wire n_789;
wire n_1232;
wire n_1603;
wire n_734;
wire n_638;
wire n_2638;
wire n_866;
wire n_969;
wire n_1401;
wire n_2492;
wire n_1019;
wire n_1105;
wire n_1998;
wire n_1338;
wire n_577;
wire n_2016;
wire n_1522;
wire n_2034;
wire n_1687;
wire n_1637;
wire n_1419;
wire n_1653;
wire n_693;
wire n_2270;
wire n_1506;
wire n_2653;
wire n_836;
wire n_990;
wire n_2496;
wire n_1886;
wire n_1389;
wire n_1894;
wire n_975;
wire n_1908;
wire n_1256;
wire n_1702;
wire n_2259;
wire n_567;
wire n_1465;
wire n_778;
wire n_1122;
wire n_2608;
wire n_2657;
wire n_770;
wire n_1375;
wire n_2494;
wire n_2649;
wire n_1102;
wire n_2392;
wire n_1843;
wire n_711;
wire n_1499;
wire n_1187;
wire n_2633;
wire n_1441;
wire n_2522;
wire n_2435;
wire n_1392;
wire n_1597;
wire n_1929;
wire n_1164;
wire n_1834;
wire n_1659;
wire n_2097;
wire n_2313;
wire n_2542;
wire n_489;
wire n_1174;
wire n_2431;
wire n_2558;
wire n_1371;
wire n_617;
wire n_1303;
wire n_2206;
wire n_2063;
wire n_1572;
wire n_1968;
wire n_2564;
wire n_2252;
wire n_876;
wire n_1516;
wire n_1190;
wire n_1736;
wire n_1685;
wire n_2409;
wire n_601;
wire n_917;
wire n_1714;
wire n_966;
wire n_1116;
wire n_2000;
wire n_1661;
wire n_1212;
wire n_2074;
wire n_1541;
wire n_2576;
wire n_726;
wire n_982;
wire n_2575;
wire n_1573;
wire n_1453;
wire n_1731;
wire n_2217;
wire n_818;
wire n_2373;
wire n_1970;
wire n_861;
wire n_1713;
wire n_1183;
wire n_2307;
wire n_1658;
wire n_899;
wire n_1253;
wire n_1737;
wire n_2201;
wire n_2117;
wire n_1904;
wire n_2640;
wire n_1993;
wire n_774;
wire n_1628;
wire n_2493;
wire n_2205;
wire n_1335;
wire n_1514;
wire n_1777;
wire n_1957;
wire n_1345;
wire n_1059;
wire n_1133;
wire n_1771;
wire n_1912;
wire n_1899;
wire n_557;
wire n_1410;
wire n_1005;
wire n_607;
wire n_1003;
wire n_679;
wire n_710;
wire n_2067;
wire n_527;
wire n_707;
wire n_1168;
wire n_2219;
wire n_2437;
wire n_2148;
wire n_937;
wire n_2445;
wire n_1427;
wire n_487;
wire n_1584;
wire n_665;
wire n_1726;
wire n_1835;
wire n_1440;
wire n_2164;
wire n_1988;
wire n_2115;
wire n_1853;
wire n_1356;
wire n_1787;
wire n_2634;
wire n_910;
wire n_2232;
wire n_2212;
wire n_2602;
wire n_1657;
wire n_768;
wire n_1475;
wire n_1302;
wire n_1774;
wire n_1725;
wire n_1136;
wire n_1313;
wire n_1491;
wire n_754;
wire n_1496;
wire n_1125;
wire n_2547;
wire n_708;
wire n_529;
wire n_1812;
wire n_735;
wire n_2501;
wire n_1915;
wire n_1109;
wire n_895;
wire n_2532;
wire n_1310;
wire n_2605;
wire n_2121;
wire n_1803;
wire n_2665;
wire n_1399;
wire n_1543;
wire n_1991;
wire n_1979;
wire n_791;
wire n_732;
wire n_2224;
wire n_1533;
wire n_808;
wire n_2484;
wire n_797;
wire n_1025;
wire n_1930;
wire n_1955;
wire n_500;
wire n_1067;
wire n_1720;
wire n_2401;
wire n_2003;
wire n_1457;
wire n_766;
wire n_541;
wire n_538;
wire n_2354;
wire n_2246;
wire n_2008;
wire n_1117;
wire n_799;
wire n_2264;
wire n_687;
wire n_715;
wire n_1742;
wire n_1480;
wire n_1482;
wire n_1213;
wire n_2489;
wire n_1266;
wire n_536;
wire n_872;
wire n_2012;
wire n_594;
wire n_1291;
wire n_1297;
wire n_1753;
wire n_2283;
wire n_1782;
wire n_2245;
wire n_1155;
wire n_1418;
wire n_1972;
wire n_1524;
wire n_1689;
wire n_1485;
wire n_1011;
wire n_2184;
wire n_1184;
wire n_985;
wire n_1855;
wire n_2425;
wire n_869;
wire n_810;
wire n_827;
wire n_1703;
wire n_1352;
wire n_626;
wire n_2197;
wire n_2199;
wire n_1650;
wire n_1144;
wire n_1137;
wire n_1570;
wire n_1170;
wire n_2023;
wire n_2213;
wire n_2351;
wire n_2211;
wire n_2095;
wire n_676;
wire n_2103;
wire n_653;
wire n_2160;
wire n_642;
wire n_2228;
wire n_2527;
wire n_1602;
wire n_2498;
wire n_855;
wire n_1178;
wire n_1461;
wire n_850;
wire n_684;
wire n_2421;
wire n_2286;
wire n_664;
wire n_1999;
wire n_503;
wire n_2372;
wire n_2065;
wire n_2136;
wire n_2480;
wire n_1372;
wire n_605;
wire n_2630;
wire n_1273;
wire n_1822;
wire n_620;
wire n_643;
wire n_2363;
wire n_2430;
wire n_916;
wire n_1081;
wire n_2549;
wire n_493;
wire n_2332;
wire n_1235;
wire n_980;
wire n_698;
wire n_1115;
wire n_703;
wire n_2433;
wire n_1282;
wire n_1318;
wire n_1783;
wire n_780;
wire n_2601;
wire n_998;
wire n_2375;
wire n_2550;
wire n_1454;
wire n_1227;
wire n_1531;
wire n_840;
wire n_1334;
wire n_1907;
wire n_501;
wire n_823;
wire n_2528;
wire n_725;
wire n_2344;
wire n_1388;
wire n_1417;
wire n_1295;
wire n_2316;
wire n_672;
wire n_1985;
wire n_1898;
wire n_2107;
wire n_581;
wire n_554;
wire n_1625;
wire n_2130;
wire n_2187;
wire n_2284;
wire n_898;
wire n_2598;
wire n_1762;
wire n_1013;
wire n_1452;
wire n_718;
wire n_1120;
wire n_719;
wire n_1791;
wire n_1890;
wire n_1747;
wire n_714;
wire n_1683;
wire n_1817;
wire n_909;
wire n_1944;
wire n_1497;
wire n_1530;
wire n_2654;
wire n_997;
wire n_932;
wire n_612;
wire n_2078;
wire n_1409;
wire n_788;
wire n_1326;
wire n_1268;
wire n_559;
wire n_825;
wire n_1981;
wire n_508;
wire n_2186;
wire n_1320;
wire n_506;
wire n_1663;
wire n_737;
wire n_1718;
wire n_986;
wire n_2315;
wire n_509;
wire n_1317;
wire n_1518;
wire n_1715;
wire n_2102;
wire n_2562;
wire n_1281;
wire n_1952;
wire n_1192;
wire n_2221;
wire n_1024;
wire n_1063;
wire n_1889;
wire n_1792;
wire n_1564;
wire n_1868;
wire n_1613;
wire n_733;
wire n_1489;
wire n_1922;
wire n_1376;
wire n_941;
wire n_2326;
wire n_981;
wire n_2560;
wire n_1569;
wire n_2188;
wire n_867;
wire n_2348;
wire n_2422;
wire n_2239;
wire n_587;
wire n_792;
wire n_756;
wire n_1429;
wire n_1238;
wire n_2448;
wire n_548;
wire n_812;
wire n_2104;
wire n_518;
wire n_505;
wire n_2057;
wire n_1772;
wire n_752;
wire n_905;
wire n_1476;
wire n_1108;
wire n_782;
wire n_1100;
wire n_1861;
wire n_2129;
wire n_1395;
wire n_862;
wire n_1425;
wire n_760;
wire n_1901;
wire n_1900;
wire n_1620;
wire n_1867;
wire n_1330;
wire n_1945;
wire n_481;
wire n_1675;
wire n_1924;
wire n_2573;
wire n_1727;
wire n_1554;
wire n_1745;
wire n_769;
wire n_2497;
wire n_2006;
wire n_1995;
wire n_2411;
wire n_2138;
wire n_1046;
wire n_934;
wire n_1618;
wire n_2260;
wire n_826;
wire n_2343;
wire n_1813;
wire n_2447;
wire n_886;
wire n_2014;
wire n_1221;
wire n_2345;
wire n_654;
wire n_1172;
wire n_2535;
wire n_1341;
wire n_570;
wire n_1641;
wire n_1361;
wire n_2382;
wire n_1707;
wire n_853;
wire n_2317;
wire n_751;
wire n_2172;
wire n_1973;
wire n_786;
wire n_1083;
wire n_1142;
wire n_2376;
wire n_2488;
wire n_1129;
wire n_2579;
wire n_2476;
wire n_704;
wire n_787;
wire n_1770;
wire n_2456;
wire n_961;
wire n_2250;
wire n_2678;
wire n_1756;
wire n_771;
wire n_1716;
wire n_1225;
wire n_1520;
wire n_2451;
wire n_522;
wire n_1287;
wire n_1262;
wire n_930;
wire n_1873;
wire n_1411;
wire n_622;
wire n_1962;
wire n_1577;
wire n_2423;
wire n_1087;
wire n_2526;
wire n_994;
wire n_1701;
wire n_2194;
wire n_848;
wire n_1550;
wire n_1498;
wire n_2167;
wire n_1223;
wire n_1272;
wire n_2680;
wire n_1567;
wire n_682;
wire n_2567;
wire n_1247;
wire n_922;
wire n_816;
wire n_1648;
wire n_591;
wire n_1536;
wire n_1857;
wire n_1344;
wire n_2041;
wire n_631;
wire n_479;
wire n_1246;
wire n_1478;
wire n_1339;
wire n_1797;
wire n_1769;
wire n_839;
wire n_1210;
wire n_1364;
wire n_2357;
wire n_2183;
wire n_2673;
wire n_2360;
wire n_2292;
wire n_1250;
wire n_2173;
wire n_1842;
wire n_871;
wire n_2442;
wire n_598;
wire n_685;
wire n_928;
wire n_1367;
wire n_608;
wire n_1943;
wire n_1460;
wire n_772;
wire n_2018;
wire n_1555;
wire n_499;
wire n_2531;
wire n_1589;
wire n_517;
wire n_1086;
wire n_2570;
wire n_796;
wire n_1858;
wire n_1619;
wire n_2119;
wire n_1502;
wire n_2157;
wire n_2552;
wire n_1469;
wire n_1012;
wire n_1396;
wire n_1348;
wire n_2030;
wire n_903;
wire n_2453;
wire n_1525;
wire n_1752;
wire n_2397;
wire n_740;
wire n_2208;
wire n_1404;
wire n_1794;
wire n_2182;
wire n_1315;
wire n_2234;
wire n_1061;
wire n_1910;
wire n_1298;
wire n_1652;
wire n_2209;
wire n_2050;
wire n_1193;
wire n_1676;
wire n_1255;
wire n_1113;
wire n_2321;
wire n_1226;
wire n_1277;
wire n_722;
wire n_2591;
wire n_2146;
wire n_844;
wire n_471;
wire n_852;
wire n_1487;
wire n_1864;
wire n_1601;
wire n_1028;
wire n_781;
wire n_474;
wire n_542;
wire n_1546;
wire n_595;
wire n_502;
wire n_2612;
wire n_1337;
wire n_1495;
wire n_632;
wire n_699;
wire n_979;
wire n_1515;
wire n_1627;
wire n_1245;
wire n_846;
wire n_2427;
wire n_2438;
wire n_2505;
wire n_1673;
wire n_1321;
wire n_1975;
wire n_2296;
wire n_2070;
wire n_1937;
wire n_585;
wire n_2112;
wire n_1739;
wire n_616;
wire n_2278;
wire n_2594;
wire n_2394;
wire n_1914;
wire n_2135;
wire n_2335;
wire n_745;
wire n_2381;
wire n_1654;
wire n_2569;
wire n_2349;
wire n_1103;
wire n_648;
wire n_1379;
wire n_2196;
wire n_2170;
wire n_1076;
wire n_1091;
wire n_1408;
wire n_494;
wire n_1761;
wire n_641;
wire n_730;
wire n_2036;
wire n_1325;
wire n_1595;
wire n_2161;
wire n_575;
wire n_480;
wire n_795;
wire n_2404;
wire n_2083;
wire n_695;
wire n_656;
wire n_1606;
wire n_2503;
wire n_1220;
wire n_1694;
wire n_1540;
wire n_2485;
wire n_1936;
wire n_1956;
wire n_1642;
wire n_2279;
wire n_2655;
wire n_2027;
wire n_2642;
wire n_1130;
wire n_720;
wire n_2500;
wire n_2366;
wire n_1918;
wire n_1526;
wire n_863;
wire n_2210;
wire n_805;
wire n_1604;
wire n_2513;
wire n_2525;
wire n_1275;
wire n_1764;
wire n_712;
wire n_2414;
wire n_1583;
wire n_2426;
wire n_1042;
wire n_1402;
wire n_2049;
wire n_2273;
wire n_1493;
wire n_657;
wire n_644;
wire n_1741;
wire n_2229;
wire n_1160;
wire n_1397;
wire n_491;
wire n_1258;
wire n_1074;
wire n_2004;
wire n_1621;
wire n_2113;
wire n_566;
wire n_565;
wire n_2586;
wire n_1448;
wire n_2225;
wire n_1507;
wire n_1398;
wire n_2383;
wire n_1879;
wire n_597;
wire n_1996;
wire n_1505;
wire n_1181;
wire n_1634;
wire n_1196;
wire n_2019;
wire n_651;
wire n_1340;
wire n_2274;
wire n_811;
wire n_1558;
wire n_807;
wire n_2166;
wire n_835;
wire n_666;
wire n_1433;
wire n_1704;
wire n_2256;
wire n_1254;
wire n_1026;
wire n_2026;
wire n_1969;
wire n_1234;
wire n_2109;
wire n_1138;
wire n_2044;
wire n_927;
wire n_1089;
wire n_2013;
wire n_1990;
wire n_1004;
wire n_1186;
wire n_1032;
wire n_2614;
wire n_2511;
wire n_1681;
wire n_2010;
wire n_1018;
wire n_2242;
wire n_2247;
wire n_1693;
wire n_2599;
wire n_713;
wire n_904;
wire n_1588;
wire n_1622;
wire n_2237;
wire n_1180;
wire n_1827;
wire n_2524;
wire n_1271;
wire n_533;
wire n_1542;
wire n_1251;
wire n_2268;

BUFx3_ASAP7_75t_L g470 ( 
.A(n_450),
.Y(n_470)
);

CKINVDCx20_ASAP7_75t_R g471 ( 
.A(n_315),
.Y(n_471)
);

CKINVDCx5p33_ASAP7_75t_R g472 ( 
.A(n_405),
.Y(n_472)
);

INVx1_ASAP7_75t_L g473 ( 
.A(n_42),
.Y(n_473)
);

CKINVDCx20_ASAP7_75t_R g474 ( 
.A(n_435),
.Y(n_474)
);

INVx1_ASAP7_75t_L g475 ( 
.A(n_428),
.Y(n_475)
);

CKINVDCx20_ASAP7_75t_R g476 ( 
.A(n_444),
.Y(n_476)
);

INVx2_ASAP7_75t_L g477 ( 
.A(n_277),
.Y(n_477)
);

INVx1_ASAP7_75t_L g478 ( 
.A(n_22),
.Y(n_478)
);

INVx1_ASAP7_75t_L g479 ( 
.A(n_241),
.Y(n_479)
);

CKINVDCx5p33_ASAP7_75t_R g480 ( 
.A(n_237),
.Y(n_480)
);

CKINVDCx5p33_ASAP7_75t_R g481 ( 
.A(n_420),
.Y(n_481)
);

CKINVDCx5p33_ASAP7_75t_R g482 ( 
.A(n_39),
.Y(n_482)
);

CKINVDCx5p33_ASAP7_75t_R g483 ( 
.A(n_431),
.Y(n_483)
);

INVx1_ASAP7_75t_L g484 ( 
.A(n_256),
.Y(n_484)
);

INVx2_ASAP7_75t_SL g485 ( 
.A(n_209),
.Y(n_485)
);

BUFx3_ASAP7_75t_L g486 ( 
.A(n_257),
.Y(n_486)
);

INVx2_ASAP7_75t_L g487 ( 
.A(n_40),
.Y(n_487)
);

INVx1_ASAP7_75t_L g488 ( 
.A(n_123),
.Y(n_488)
);

BUFx2_ASAP7_75t_L g489 ( 
.A(n_463),
.Y(n_489)
);

INVx1_ASAP7_75t_L g490 ( 
.A(n_397),
.Y(n_490)
);

INVx2_ASAP7_75t_L g491 ( 
.A(n_229),
.Y(n_491)
);

BUFx3_ASAP7_75t_L g492 ( 
.A(n_44),
.Y(n_492)
);

INVx1_ASAP7_75t_L g493 ( 
.A(n_197),
.Y(n_493)
);

CKINVDCx5p33_ASAP7_75t_R g494 ( 
.A(n_196),
.Y(n_494)
);

BUFx3_ASAP7_75t_L g495 ( 
.A(n_178),
.Y(n_495)
);

CKINVDCx5p33_ASAP7_75t_R g496 ( 
.A(n_175),
.Y(n_496)
);

CKINVDCx16_ASAP7_75t_R g497 ( 
.A(n_40),
.Y(n_497)
);

CKINVDCx5p33_ASAP7_75t_R g498 ( 
.A(n_422),
.Y(n_498)
);

CKINVDCx5p33_ASAP7_75t_R g499 ( 
.A(n_79),
.Y(n_499)
);

CKINVDCx5p33_ASAP7_75t_R g500 ( 
.A(n_111),
.Y(n_500)
);

CKINVDCx5p33_ASAP7_75t_R g501 ( 
.A(n_401),
.Y(n_501)
);

CKINVDCx5p33_ASAP7_75t_R g502 ( 
.A(n_168),
.Y(n_502)
);

CKINVDCx5p33_ASAP7_75t_R g503 ( 
.A(n_313),
.Y(n_503)
);

CKINVDCx5p33_ASAP7_75t_R g504 ( 
.A(n_167),
.Y(n_504)
);

CKINVDCx5p33_ASAP7_75t_R g505 ( 
.A(n_305),
.Y(n_505)
);

CKINVDCx5p33_ASAP7_75t_R g506 ( 
.A(n_441),
.Y(n_506)
);

INVx2_ASAP7_75t_SL g507 ( 
.A(n_56),
.Y(n_507)
);

CKINVDCx5p33_ASAP7_75t_R g508 ( 
.A(n_90),
.Y(n_508)
);

CKINVDCx5p33_ASAP7_75t_R g509 ( 
.A(n_411),
.Y(n_509)
);

CKINVDCx5p33_ASAP7_75t_R g510 ( 
.A(n_416),
.Y(n_510)
);

CKINVDCx5p33_ASAP7_75t_R g511 ( 
.A(n_59),
.Y(n_511)
);

CKINVDCx5p33_ASAP7_75t_R g512 ( 
.A(n_354),
.Y(n_512)
);

BUFx2_ASAP7_75t_L g513 ( 
.A(n_298),
.Y(n_513)
);

CKINVDCx5p33_ASAP7_75t_R g514 ( 
.A(n_201),
.Y(n_514)
);

CKINVDCx5p33_ASAP7_75t_R g515 ( 
.A(n_171),
.Y(n_515)
);

CKINVDCx5p33_ASAP7_75t_R g516 ( 
.A(n_126),
.Y(n_516)
);

CKINVDCx5p33_ASAP7_75t_R g517 ( 
.A(n_227),
.Y(n_517)
);

BUFx2_ASAP7_75t_L g518 ( 
.A(n_22),
.Y(n_518)
);

CKINVDCx5p33_ASAP7_75t_R g519 ( 
.A(n_171),
.Y(n_519)
);

CKINVDCx5p33_ASAP7_75t_R g520 ( 
.A(n_252),
.Y(n_520)
);

INVx1_ASAP7_75t_L g521 ( 
.A(n_449),
.Y(n_521)
);

INVx1_ASAP7_75t_L g522 ( 
.A(n_215),
.Y(n_522)
);

INVx2_ASAP7_75t_L g523 ( 
.A(n_26),
.Y(n_523)
);

CKINVDCx5p33_ASAP7_75t_R g524 ( 
.A(n_148),
.Y(n_524)
);

CKINVDCx5p33_ASAP7_75t_R g525 ( 
.A(n_170),
.Y(n_525)
);

CKINVDCx5p33_ASAP7_75t_R g526 ( 
.A(n_122),
.Y(n_526)
);

BUFx2_ASAP7_75t_L g527 ( 
.A(n_125),
.Y(n_527)
);

CKINVDCx5p33_ASAP7_75t_R g528 ( 
.A(n_47),
.Y(n_528)
);

INVx1_ASAP7_75t_L g529 ( 
.A(n_100),
.Y(n_529)
);

CKINVDCx5p33_ASAP7_75t_R g530 ( 
.A(n_378),
.Y(n_530)
);

CKINVDCx5p33_ASAP7_75t_R g531 ( 
.A(n_436),
.Y(n_531)
);

BUFx6f_ASAP7_75t_L g532 ( 
.A(n_15),
.Y(n_532)
);

CKINVDCx5p33_ASAP7_75t_R g533 ( 
.A(n_375),
.Y(n_533)
);

CKINVDCx5p33_ASAP7_75t_R g534 ( 
.A(n_61),
.Y(n_534)
);

CKINVDCx5p33_ASAP7_75t_R g535 ( 
.A(n_340),
.Y(n_535)
);

CKINVDCx5p33_ASAP7_75t_R g536 ( 
.A(n_4),
.Y(n_536)
);

CKINVDCx5p33_ASAP7_75t_R g537 ( 
.A(n_443),
.Y(n_537)
);

INVx1_ASAP7_75t_L g538 ( 
.A(n_247),
.Y(n_538)
);

INVx2_ASAP7_75t_SL g539 ( 
.A(n_336),
.Y(n_539)
);

CKINVDCx5p33_ASAP7_75t_R g540 ( 
.A(n_185),
.Y(n_540)
);

INVx1_ASAP7_75t_L g541 ( 
.A(n_138),
.Y(n_541)
);

CKINVDCx20_ASAP7_75t_R g542 ( 
.A(n_303),
.Y(n_542)
);

INVx2_ASAP7_75t_L g543 ( 
.A(n_77),
.Y(n_543)
);

CKINVDCx16_ASAP7_75t_R g544 ( 
.A(n_54),
.Y(n_544)
);

INVx2_ASAP7_75t_SL g545 ( 
.A(n_243),
.Y(n_545)
);

CKINVDCx5p33_ASAP7_75t_R g546 ( 
.A(n_128),
.Y(n_546)
);

CKINVDCx20_ASAP7_75t_R g547 ( 
.A(n_294),
.Y(n_547)
);

CKINVDCx5p33_ASAP7_75t_R g548 ( 
.A(n_395),
.Y(n_548)
);

INVx2_ASAP7_75t_L g549 ( 
.A(n_264),
.Y(n_549)
);

CKINVDCx5p33_ASAP7_75t_R g550 ( 
.A(n_136),
.Y(n_550)
);

CKINVDCx5p33_ASAP7_75t_R g551 ( 
.A(n_3),
.Y(n_551)
);

CKINVDCx5p33_ASAP7_75t_R g552 ( 
.A(n_271),
.Y(n_552)
);

INVx1_ASAP7_75t_L g553 ( 
.A(n_41),
.Y(n_553)
);

INVx1_ASAP7_75t_L g554 ( 
.A(n_224),
.Y(n_554)
);

CKINVDCx5p33_ASAP7_75t_R g555 ( 
.A(n_286),
.Y(n_555)
);

CKINVDCx5p33_ASAP7_75t_R g556 ( 
.A(n_393),
.Y(n_556)
);

CKINVDCx5p33_ASAP7_75t_R g557 ( 
.A(n_109),
.Y(n_557)
);

CKINVDCx5p33_ASAP7_75t_R g558 ( 
.A(n_267),
.Y(n_558)
);

INVx1_ASAP7_75t_L g559 ( 
.A(n_387),
.Y(n_559)
);

INVx1_ASAP7_75t_L g560 ( 
.A(n_418),
.Y(n_560)
);

CKINVDCx5p33_ASAP7_75t_R g561 ( 
.A(n_151),
.Y(n_561)
);

CKINVDCx5p33_ASAP7_75t_R g562 ( 
.A(n_353),
.Y(n_562)
);

INVx1_ASAP7_75t_L g563 ( 
.A(n_251),
.Y(n_563)
);

CKINVDCx20_ASAP7_75t_R g564 ( 
.A(n_53),
.Y(n_564)
);

CKINVDCx5p33_ASAP7_75t_R g565 ( 
.A(n_290),
.Y(n_565)
);

INVx1_ASAP7_75t_L g566 ( 
.A(n_459),
.Y(n_566)
);

INVx1_ASAP7_75t_L g567 ( 
.A(n_59),
.Y(n_567)
);

CKINVDCx5p33_ASAP7_75t_R g568 ( 
.A(n_438),
.Y(n_568)
);

INVx1_ASAP7_75t_L g569 ( 
.A(n_20),
.Y(n_569)
);

CKINVDCx5p33_ASAP7_75t_R g570 ( 
.A(n_226),
.Y(n_570)
);

CKINVDCx5p33_ASAP7_75t_R g571 ( 
.A(n_417),
.Y(n_571)
);

INVx1_ASAP7_75t_L g572 ( 
.A(n_276),
.Y(n_572)
);

CKINVDCx5p33_ASAP7_75t_R g573 ( 
.A(n_423),
.Y(n_573)
);

INVx1_ASAP7_75t_L g574 ( 
.A(n_239),
.Y(n_574)
);

INVx2_ASAP7_75t_L g575 ( 
.A(n_338),
.Y(n_575)
);

CKINVDCx20_ASAP7_75t_R g576 ( 
.A(n_130),
.Y(n_576)
);

CKINVDCx5p33_ASAP7_75t_R g577 ( 
.A(n_49),
.Y(n_577)
);

CKINVDCx5p33_ASAP7_75t_R g578 ( 
.A(n_64),
.Y(n_578)
);

CKINVDCx20_ASAP7_75t_R g579 ( 
.A(n_413),
.Y(n_579)
);

CKINVDCx20_ASAP7_75t_R g580 ( 
.A(n_119),
.Y(n_580)
);

CKINVDCx5p33_ASAP7_75t_R g581 ( 
.A(n_385),
.Y(n_581)
);

CKINVDCx5p33_ASAP7_75t_R g582 ( 
.A(n_299),
.Y(n_582)
);

CKINVDCx5p33_ASAP7_75t_R g583 ( 
.A(n_145),
.Y(n_583)
);

CKINVDCx16_ASAP7_75t_R g584 ( 
.A(n_206),
.Y(n_584)
);

CKINVDCx5p33_ASAP7_75t_R g585 ( 
.A(n_41),
.Y(n_585)
);

CKINVDCx5p33_ASAP7_75t_R g586 ( 
.A(n_26),
.Y(n_586)
);

CKINVDCx5p33_ASAP7_75t_R g587 ( 
.A(n_137),
.Y(n_587)
);

HB1xp67_ASAP7_75t_L g588 ( 
.A(n_211),
.Y(n_588)
);

CKINVDCx5p33_ASAP7_75t_R g589 ( 
.A(n_451),
.Y(n_589)
);

BUFx2_ASAP7_75t_L g590 ( 
.A(n_371),
.Y(n_590)
);

CKINVDCx5p33_ASAP7_75t_R g591 ( 
.A(n_249),
.Y(n_591)
);

CKINVDCx5p33_ASAP7_75t_R g592 ( 
.A(n_202),
.Y(n_592)
);

CKINVDCx5p33_ASAP7_75t_R g593 ( 
.A(n_27),
.Y(n_593)
);

INVx2_ASAP7_75t_L g594 ( 
.A(n_140),
.Y(n_594)
);

INVx1_ASAP7_75t_L g595 ( 
.A(n_390),
.Y(n_595)
);

INVx1_ASAP7_75t_L g596 ( 
.A(n_181),
.Y(n_596)
);

INVx1_ASAP7_75t_SL g597 ( 
.A(n_319),
.Y(n_597)
);

CKINVDCx5p33_ASAP7_75t_R g598 ( 
.A(n_62),
.Y(n_598)
);

INVx1_ASAP7_75t_L g599 ( 
.A(n_51),
.Y(n_599)
);

INVx1_ASAP7_75t_L g600 ( 
.A(n_377),
.Y(n_600)
);

BUFx3_ASAP7_75t_L g601 ( 
.A(n_164),
.Y(n_601)
);

CKINVDCx5p33_ASAP7_75t_R g602 ( 
.A(n_349),
.Y(n_602)
);

INVx1_ASAP7_75t_L g603 ( 
.A(n_330),
.Y(n_603)
);

CKINVDCx5p33_ASAP7_75t_R g604 ( 
.A(n_242),
.Y(n_604)
);

BUFx10_ASAP7_75t_L g605 ( 
.A(n_322),
.Y(n_605)
);

CKINVDCx5p33_ASAP7_75t_R g606 ( 
.A(n_94),
.Y(n_606)
);

INVx1_ASAP7_75t_SL g607 ( 
.A(n_123),
.Y(n_607)
);

CKINVDCx5p33_ASAP7_75t_R g608 ( 
.A(n_13),
.Y(n_608)
);

BUFx2_ASAP7_75t_SL g609 ( 
.A(n_2),
.Y(n_609)
);

INVx1_ASAP7_75t_L g610 ( 
.A(n_301),
.Y(n_610)
);

CKINVDCx5p33_ASAP7_75t_R g611 ( 
.A(n_85),
.Y(n_611)
);

CKINVDCx5p33_ASAP7_75t_R g612 ( 
.A(n_45),
.Y(n_612)
);

CKINVDCx5p33_ASAP7_75t_R g613 ( 
.A(n_402),
.Y(n_613)
);

CKINVDCx16_ASAP7_75t_R g614 ( 
.A(n_152),
.Y(n_614)
);

CKINVDCx16_ASAP7_75t_R g615 ( 
.A(n_212),
.Y(n_615)
);

CKINVDCx5p33_ASAP7_75t_R g616 ( 
.A(n_445),
.Y(n_616)
);

CKINVDCx5p33_ASAP7_75t_R g617 ( 
.A(n_275),
.Y(n_617)
);

INVx1_ASAP7_75t_L g618 ( 
.A(n_312),
.Y(n_618)
);

CKINVDCx5p33_ASAP7_75t_R g619 ( 
.A(n_403),
.Y(n_619)
);

INVx1_ASAP7_75t_SL g620 ( 
.A(n_88),
.Y(n_620)
);

INVx1_ASAP7_75t_L g621 ( 
.A(n_56),
.Y(n_621)
);

CKINVDCx5p33_ASAP7_75t_R g622 ( 
.A(n_461),
.Y(n_622)
);

BUFx10_ASAP7_75t_L g623 ( 
.A(n_137),
.Y(n_623)
);

BUFx3_ASAP7_75t_L g624 ( 
.A(n_182),
.Y(n_624)
);

INVx1_ASAP7_75t_L g625 ( 
.A(n_159),
.Y(n_625)
);

INVx1_ASAP7_75t_L g626 ( 
.A(n_38),
.Y(n_626)
);

BUFx2_ASAP7_75t_L g627 ( 
.A(n_58),
.Y(n_627)
);

INVx1_ASAP7_75t_L g628 ( 
.A(n_205),
.Y(n_628)
);

INVx1_ASAP7_75t_L g629 ( 
.A(n_283),
.Y(n_629)
);

BUFx2_ASAP7_75t_L g630 ( 
.A(n_469),
.Y(n_630)
);

CKINVDCx20_ASAP7_75t_R g631 ( 
.A(n_207),
.Y(n_631)
);

BUFx10_ASAP7_75t_L g632 ( 
.A(n_108),
.Y(n_632)
);

INVx1_ASAP7_75t_L g633 ( 
.A(n_83),
.Y(n_633)
);

INVx1_ASAP7_75t_L g634 ( 
.A(n_214),
.Y(n_634)
);

CKINVDCx5p33_ASAP7_75t_R g635 ( 
.A(n_339),
.Y(n_635)
);

CKINVDCx5p33_ASAP7_75t_R g636 ( 
.A(n_363),
.Y(n_636)
);

CKINVDCx5p33_ASAP7_75t_R g637 ( 
.A(n_53),
.Y(n_637)
);

INVx1_ASAP7_75t_L g638 ( 
.A(n_284),
.Y(n_638)
);

INVx1_ASAP7_75t_L g639 ( 
.A(n_381),
.Y(n_639)
);

CKINVDCx5p33_ASAP7_75t_R g640 ( 
.A(n_213),
.Y(n_640)
);

CKINVDCx5p33_ASAP7_75t_R g641 ( 
.A(n_72),
.Y(n_641)
);

CKINVDCx5p33_ASAP7_75t_R g642 ( 
.A(n_188),
.Y(n_642)
);

BUFx10_ASAP7_75t_L g643 ( 
.A(n_145),
.Y(n_643)
);

INVx2_ASAP7_75t_L g644 ( 
.A(n_28),
.Y(n_644)
);

CKINVDCx5p33_ASAP7_75t_R g645 ( 
.A(n_272),
.Y(n_645)
);

CKINVDCx20_ASAP7_75t_R g646 ( 
.A(n_25),
.Y(n_646)
);

BUFx10_ASAP7_75t_L g647 ( 
.A(n_325),
.Y(n_647)
);

INVx1_ASAP7_75t_L g648 ( 
.A(n_238),
.Y(n_648)
);

INVx1_ASAP7_75t_L g649 ( 
.A(n_394),
.Y(n_649)
);

CKINVDCx5p33_ASAP7_75t_R g650 ( 
.A(n_115),
.Y(n_650)
);

BUFx10_ASAP7_75t_L g651 ( 
.A(n_347),
.Y(n_651)
);

BUFx6f_ASAP7_75t_L g652 ( 
.A(n_198),
.Y(n_652)
);

INVx1_ASAP7_75t_L g653 ( 
.A(n_12),
.Y(n_653)
);

INVx1_ASAP7_75t_L g654 ( 
.A(n_92),
.Y(n_654)
);

CKINVDCx5p33_ASAP7_75t_R g655 ( 
.A(n_162),
.Y(n_655)
);

INVx2_ASAP7_75t_L g656 ( 
.A(n_50),
.Y(n_656)
);

BUFx10_ASAP7_75t_L g657 ( 
.A(n_373),
.Y(n_657)
);

INVx1_ASAP7_75t_L g658 ( 
.A(n_462),
.Y(n_658)
);

CKINVDCx20_ASAP7_75t_R g659 ( 
.A(n_148),
.Y(n_659)
);

INVx1_ASAP7_75t_L g660 ( 
.A(n_174),
.Y(n_660)
);

INVx1_ASAP7_75t_L g661 ( 
.A(n_195),
.Y(n_661)
);

CKINVDCx14_ASAP7_75t_R g662 ( 
.A(n_289),
.Y(n_662)
);

INVx1_ASAP7_75t_L g663 ( 
.A(n_107),
.Y(n_663)
);

CKINVDCx20_ASAP7_75t_R g664 ( 
.A(n_159),
.Y(n_664)
);

CKINVDCx5p33_ASAP7_75t_R g665 ( 
.A(n_259),
.Y(n_665)
);

CKINVDCx20_ASAP7_75t_R g666 ( 
.A(n_76),
.Y(n_666)
);

CKINVDCx5p33_ASAP7_75t_R g667 ( 
.A(n_235),
.Y(n_667)
);

INVx1_ASAP7_75t_L g668 ( 
.A(n_84),
.Y(n_668)
);

INVx2_ASAP7_75t_L g669 ( 
.A(n_425),
.Y(n_669)
);

CKINVDCx5p33_ASAP7_75t_R g670 ( 
.A(n_16),
.Y(n_670)
);

CKINVDCx5p33_ASAP7_75t_R g671 ( 
.A(n_199),
.Y(n_671)
);

INVx1_ASAP7_75t_L g672 ( 
.A(n_295),
.Y(n_672)
);

BUFx3_ASAP7_75t_L g673 ( 
.A(n_320),
.Y(n_673)
);

INVx2_ASAP7_75t_SL g674 ( 
.A(n_404),
.Y(n_674)
);

CKINVDCx5p33_ASAP7_75t_R g675 ( 
.A(n_399),
.Y(n_675)
);

CKINVDCx5p33_ASAP7_75t_R g676 ( 
.A(n_99),
.Y(n_676)
);

CKINVDCx5p33_ASAP7_75t_R g677 ( 
.A(n_254),
.Y(n_677)
);

CKINVDCx5p33_ASAP7_75t_R g678 ( 
.A(n_155),
.Y(n_678)
);

CKINVDCx5p33_ASAP7_75t_R g679 ( 
.A(n_384),
.Y(n_679)
);

INVx1_ASAP7_75t_L g680 ( 
.A(n_292),
.Y(n_680)
);

INVx2_ASAP7_75t_L g681 ( 
.A(n_231),
.Y(n_681)
);

CKINVDCx5p33_ASAP7_75t_R g682 ( 
.A(n_454),
.Y(n_682)
);

INVx1_ASAP7_75t_L g683 ( 
.A(n_360),
.Y(n_683)
);

CKINVDCx5p33_ASAP7_75t_R g684 ( 
.A(n_466),
.Y(n_684)
);

CKINVDCx5p33_ASAP7_75t_R g685 ( 
.A(n_458),
.Y(n_685)
);

INVx2_ASAP7_75t_L g686 ( 
.A(n_194),
.Y(n_686)
);

INVx1_ASAP7_75t_L g687 ( 
.A(n_110),
.Y(n_687)
);

BUFx10_ASAP7_75t_L g688 ( 
.A(n_55),
.Y(n_688)
);

CKINVDCx5p33_ASAP7_75t_R g689 ( 
.A(n_33),
.Y(n_689)
);

INVx1_ASAP7_75t_L g690 ( 
.A(n_191),
.Y(n_690)
);

CKINVDCx5p33_ASAP7_75t_R g691 ( 
.A(n_129),
.Y(n_691)
);

CKINVDCx20_ASAP7_75t_R g692 ( 
.A(n_116),
.Y(n_692)
);

INVx2_ASAP7_75t_L g693 ( 
.A(n_204),
.Y(n_693)
);

INVx1_ASAP7_75t_L g694 ( 
.A(n_316),
.Y(n_694)
);

INVx1_ASAP7_75t_L g695 ( 
.A(n_208),
.Y(n_695)
);

INVx1_ASAP7_75t_L g696 ( 
.A(n_314),
.Y(n_696)
);

INVx1_ASAP7_75t_L g697 ( 
.A(n_125),
.Y(n_697)
);

INVx1_ASAP7_75t_L g698 ( 
.A(n_17),
.Y(n_698)
);

CKINVDCx5p33_ASAP7_75t_R g699 ( 
.A(n_306),
.Y(n_699)
);

INVx1_ASAP7_75t_L g700 ( 
.A(n_258),
.Y(n_700)
);

BUFx2_ASAP7_75t_L g701 ( 
.A(n_27),
.Y(n_701)
);

CKINVDCx5p33_ASAP7_75t_R g702 ( 
.A(n_13),
.Y(n_702)
);

CKINVDCx5p33_ASAP7_75t_R g703 ( 
.A(n_439),
.Y(n_703)
);

BUFx3_ASAP7_75t_L g704 ( 
.A(n_138),
.Y(n_704)
);

CKINVDCx5p33_ASAP7_75t_R g705 ( 
.A(n_147),
.Y(n_705)
);

INVx1_ASAP7_75t_L g706 ( 
.A(n_464),
.Y(n_706)
);

INVx1_ASAP7_75t_L g707 ( 
.A(n_261),
.Y(n_707)
);

CKINVDCx20_ASAP7_75t_R g708 ( 
.A(n_369),
.Y(n_708)
);

INVx1_ASAP7_75t_L g709 ( 
.A(n_465),
.Y(n_709)
);

CKINVDCx5p33_ASAP7_75t_R g710 ( 
.A(n_115),
.Y(n_710)
);

INVx2_ASAP7_75t_L g711 ( 
.A(n_165),
.Y(n_711)
);

CKINVDCx5p33_ASAP7_75t_R g712 ( 
.A(n_135),
.Y(n_712)
);

INVx1_ASAP7_75t_L g713 ( 
.A(n_84),
.Y(n_713)
);

CKINVDCx5p33_ASAP7_75t_R g714 ( 
.A(n_167),
.Y(n_714)
);

INVx1_ASAP7_75t_L g715 ( 
.A(n_75),
.Y(n_715)
);

CKINVDCx5p33_ASAP7_75t_R g716 ( 
.A(n_67),
.Y(n_716)
);

CKINVDCx5p33_ASAP7_75t_R g717 ( 
.A(n_291),
.Y(n_717)
);

INVx1_ASAP7_75t_L g718 ( 
.A(n_396),
.Y(n_718)
);

INVx1_ASAP7_75t_L g719 ( 
.A(n_55),
.Y(n_719)
);

CKINVDCx5p33_ASAP7_75t_R g720 ( 
.A(n_210),
.Y(n_720)
);

CKINVDCx5p33_ASAP7_75t_R g721 ( 
.A(n_18),
.Y(n_721)
);

CKINVDCx5p33_ASAP7_75t_R g722 ( 
.A(n_97),
.Y(n_722)
);

CKINVDCx5p33_ASAP7_75t_R g723 ( 
.A(n_421),
.Y(n_723)
);

INVx1_ASAP7_75t_L g724 ( 
.A(n_361),
.Y(n_724)
);

INVx1_ASAP7_75t_L g725 ( 
.A(n_356),
.Y(n_725)
);

CKINVDCx5p33_ASAP7_75t_R g726 ( 
.A(n_135),
.Y(n_726)
);

BUFx8_ASAP7_75t_SL g727 ( 
.A(n_88),
.Y(n_727)
);

CKINVDCx5p33_ASAP7_75t_R g728 ( 
.A(n_297),
.Y(n_728)
);

INVx2_ASAP7_75t_L g729 ( 
.A(n_153),
.Y(n_729)
);

INVx1_ASAP7_75t_L g730 ( 
.A(n_10),
.Y(n_730)
);

INVx2_ASAP7_75t_L g731 ( 
.A(n_343),
.Y(n_731)
);

INVx1_ASAP7_75t_L g732 ( 
.A(n_156),
.Y(n_732)
);

INVx1_ASAP7_75t_SL g733 ( 
.A(n_447),
.Y(n_733)
);

CKINVDCx5p33_ASAP7_75t_R g734 ( 
.A(n_351),
.Y(n_734)
);

INVx1_ASAP7_75t_L g735 ( 
.A(n_304),
.Y(n_735)
);

INVx1_ASAP7_75t_L g736 ( 
.A(n_448),
.Y(n_736)
);

CKINVDCx20_ASAP7_75t_R g737 ( 
.A(n_161),
.Y(n_737)
);

INVx1_ASAP7_75t_L g738 ( 
.A(n_430),
.Y(n_738)
);

INVx1_ASAP7_75t_L g739 ( 
.A(n_37),
.Y(n_739)
);

CKINVDCx5p33_ASAP7_75t_R g740 ( 
.A(n_124),
.Y(n_740)
);

INVx1_ASAP7_75t_L g741 ( 
.A(n_102),
.Y(n_741)
);

CKINVDCx5p33_ASAP7_75t_R g742 ( 
.A(n_66),
.Y(n_742)
);

CKINVDCx5p33_ASAP7_75t_R g743 ( 
.A(n_80),
.Y(n_743)
);

INVx1_ASAP7_75t_L g744 ( 
.A(n_370),
.Y(n_744)
);

CKINVDCx20_ASAP7_75t_R g745 ( 
.A(n_419),
.Y(n_745)
);

CKINVDCx5p33_ASAP7_75t_R g746 ( 
.A(n_85),
.Y(n_746)
);

INVx1_ASAP7_75t_L g747 ( 
.A(n_203),
.Y(n_747)
);

CKINVDCx5p33_ASAP7_75t_R g748 ( 
.A(n_341),
.Y(n_748)
);

CKINVDCx5p33_ASAP7_75t_R g749 ( 
.A(n_96),
.Y(n_749)
);

CKINVDCx5p33_ASAP7_75t_R g750 ( 
.A(n_233),
.Y(n_750)
);

CKINVDCx5p33_ASAP7_75t_R g751 ( 
.A(n_260),
.Y(n_751)
);

CKINVDCx5p33_ASAP7_75t_R g752 ( 
.A(n_323),
.Y(n_752)
);

INVx1_ASAP7_75t_L g753 ( 
.A(n_326),
.Y(n_753)
);

BUFx6f_ASAP7_75t_L g754 ( 
.A(n_350),
.Y(n_754)
);

INVx1_ASAP7_75t_L g755 ( 
.A(n_155),
.Y(n_755)
);

INVx1_ASAP7_75t_L g756 ( 
.A(n_218),
.Y(n_756)
);

CKINVDCx5p33_ASAP7_75t_R g757 ( 
.A(n_179),
.Y(n_757)
);

BUFx10_ASAP7_75t_L g758 ( 
.A(n_16),
.Y(n_758)
);

CKINVDCx20_ASAP7_75t_R g759 ( 
.A(n_429),
.Y(n_759)
);

CKINVDCx5p33_ASAP7_75t_R g760 ( 
.A(n_75),
.Y(n_760)
);

INVxp67_ASAP7_75t_L g761 ( 
.A(n_166),
.Y(n_761)
);

INVx1_ASAP7_75t_L g762 ( 
.A(n_165),
.Y(n_762)
);

CKINVDCx5p33_ASAP7_75t_R g763 ( 
.A(n_72),
.Y(n_763)
);

BUFx3_ASAP7_75t_L g764 ( 
.A(n_29),
.Y(n_764)
);

INVx1_ASAP7_75t_L g765 ( 
.A(n_187),
.Y(n_765)
);

CKINVDCx5p33_ASAP7_75t_R g766 ( 
.A(n_124),
.Y(n_766)
);

CKINVDCx5p33_ASAP7_75t_R g767 ( 
.A(n_70),
.Y(n_767)
);

INVx1_ASAP7_75t_L g768 ( 
.A(n_36),
.Y(n_768)
);

CKINVDCx5p33_ASAP7_75t_R g769 ( 
.A(n_380),
.Y(n_769)
);

INVx1_ASAP7_75t_L g770 ( 
.A(n_104),
.Y(n_770)
);

CKINVDCx5p33_ASAP7_75t_R g771 ( 
.A(n_246),
.Y(n_771)
);

CKINVDCx5p33_ASAP7_75t_R g772 ( 
.A(n_285),
.Y(n_772)
);

CKINVDCx5p33_ASAP7_75t_R g773 ( 
.A(n_51),
.Y(n_773)
);

CKINVDCx5p33_ASAP7_75t_R g774 ( 
.A(n_389),
.Y(n_774)
);

INVx1_ASAP7_75t_L g775 ( 
.A(n_334),
.Y(n_775)
);

CKINVDCx5p33_ASAP7_75t_R g776 ( 
.A(n_221),
.Y(n_776)
);

CKINVDCx5p33_ASAP7_75t_R g777 ( 
.A(n_184),
.Y(n_777)
);

INVx1_ASAP7_75t_L g778 ( 
.A(n_318),
.Y(n_778)
);

CKINVDCx5p33_ASAP7_75t_R g779 ( 
.A(n_268),
.Y(n_779)
);

CKINVDCx5p33_ASAP7_75t_R g780 ( 
.A(n_392),
.Y(n_780)
);

INVx3_ASAP7_75t_L g781 ( 
.A(n_410),
.Y(n_781)
);

CKINVDCx5p33_ASAP7_75t_R g782 ( 
.A(n_153),
.Y(n_782)
);

CKINVDCx5p33_ASAP7_75t_R g783 ( 
.A(n_321),
.Y(n_783)
);

CKINVDCx5p33_ASAP7_75t_R g784 ( 
.A(n_95),
.Y(n_784)
);

CKINVDCx5p33_ASAP7_75t_R g785 ( 
.A(n_100),
.Y(n_785)
);

CKINVDCx14_ASAP7_75t_R g786 ( 
.A(n_406),
.Y(n_786)
);

CKINVDCx20_ASAP7_75t_R g787 ( 
.A(n_269),
.Y(n_787)
);

CKINVDCx5p33_ASAP7_75t_R g788 ( 
.A(n_54),
.Y(n_788)
);

CKINVDCx5p33_ASAP7_75t_R g789 ( 
.A(n_412),
.Y(n_789)
);

CKINVDCx20_ASAP7_75t_R g790 ( 
.A(n_300),
.Y(n_790)
);

INVxp67_ASAP7_75t_SL g791 ( 
.A(n_44),
.Y(n_791)
);

BUFx3_ASAP7_75t_L g792 ( 
.A(n_391),
.Y(n_792)
);

CKINVDCx5p33_ASAP7_75t_R g793 ( 
.A(n_440),
.Y(n_793)
);

INVx1_ASAP7_75t_SL g794 ( 
.A(n_240),
.Y(n_794)
);

INVx1_ASAP7_75t_L g795 ( 
.A(n_359),
.Y(n_795)
);

CKINVDCx5p33_ASAP7_75t_R g796 ( 
.A(n_357),
.Y(n_796)
);

INVx1_ASAP7_75t_L g797 ( 
.A(n_255),
.Y(n_797)
);

CKINVDCx5p33_ASAP7_75t_R g798 ( 
.A(n_105),
.Y(n_798)
);

CKINVDCx5p33_ASAP7_75t_R g799 ( 
.A(n_96),
.Y(n_799)
);

CKINVDCx5p33_ASAP7_75t_R g800 ( 
.A(n_376),
.Y(n_800)
);

INVx1_ASAP7_75t_L g801 ( 
.A(n_61),
.Y(n_801)
);

CKINVDCx5p33_ASAP7_75t_R g802 ( 
.A(n_141),
.Y(n_802)
);

CKINVDCx5p33_ASAP7_75t_R g803 ( 
.A(n_68),
.Y(n_803)
);

INVx1_ASAP7_75t_L g804 ( 
.A(n_28),
.Y(n_804)
);

CKINVDCx20_ASAP7_75t_R g805 ( 
.A(n_119),
.Y(n_805)
);

INVx1_ASAP7_75t_L g806 ( 
.A(n_358),
.Y(n_806)
);

BUFx8_ASAP7_75t_SL g807 ( 
.A(n_200),
.Y(n_807)
);

CKINVDCx5p33_ASAP7_75t_R g808 ( 
.A(n_433),
.Y(n_808)
);

CKINVDCx5p33_ASAP7_75t_R g809 ( 
.A(n_142),
.Y(n_809)
);

INVx1_ASAP7_75t_L g810 ( 
.A(n_160),
.Y(n_810)
);

CKINVDCx20_ASAP7_75t_R g811 ( 
.A(n_35),
.Y(n_811)
);

INVx1_ASAP7_75t_L g812 ( 
.A(n_143),
.Y(n_812)
);

INVx2_ASAP7_75t_L g813 ( 
.A(n_263),
.Y(n_813)
);

CKINVDCx5p33_ASAP7_75t_R g814 ( 
.A(n_342),
.Y(n_814)
);

CKINVDCx20_ASAP7_75t_R g815 ( 
.A(n_7),
.Y(n_815)
);

CKINVDCx5p33_ASAP7_75t_R g816 ( 
.A(n_183),
.Y(n_816)
);

BUFx3_ASAP7_75t_L g817 ( 
.A(n_144),
.Y(n_817)
);

CKINVDCx5p33_ASAP7_75t_R g818 ( 
.A(n_57),
.Y(n_818)
);

CKINVDCx5p33_ASAP7_75t_R g819 ( 
.A(n_219),
.Y(n_819)
);

CKINVDCx20_ASAP7_75t_R g820 ( 
.A(n_149),
.Y(n_820)
);

INVx1_ASAP7_75t_SL g821 ( 
.A(n_110),
.Y(n_821)
);

CKINVDCx5p33_ASAP7_75t_R g822 ( 
.A(n_126),
.Y(n_822)
);

CKINVDCx16_ASAP7_75t_R g823 ( 
.A(n_36),
.Y(n_823)
);

INVx1_ASAP7_75t_L g824 ( 
.A(n_64),
.Y(n_824)
);

CKINVDCx5p33_ASAP7_75t_R g825 ( 
.A(n_352),
.Y(n_825)
);

CKINVDCx5p33_ASAP7_75t_R g826 ( 
.A(n_81),
.Y(n_826)
);

INVx1_ASAP7_75t_L g827 ( 
.A(n_492),
.Y(n_827)
);

INVx1_ASAP7_75t_L g828 ( 
.A(n_492),
.Y(n_828)
);

NOR2xp33_ASAP7_75t_L g829 ( 
.A(n_485),
.B(n_0),
.Y(n_829)
);

INVxp67_ASAP7_75t_SL g830 ( 
.A(n_588),
.Y(n_830)
);

INVx2_ASAP7_75t_L g831 ( 
.A(n_532),
.Y(n_831)
);

INVx1_ASAP7_75t_L g832 ( 
.A(n_601),
.Y(n_832)
);

INVx1_ASAP7_75t_L g833 ( 
.A(n_601),
.Y(n_833)
);

INVx2_ASAP7_75t_L g834 ( 
.A(n_532),
.Y(n_834)
);

INVx1_ASAP7_75t_L g835 ( 
.A(n_704),
.Y(n_835)
);

CKINVDCx14_ASAP7_75t_R g836 ( 
.A(n_662),
.Y(n_836)
);

INVx1_ASAP7_75t_L g837 ( 
.A(n_704),
.Y(n_837)
);

BUFx2_ASAP7_75t_L g838 ( 
.A(n_727),
.Y(n_838)
);

INVx1_ASAP7_75t_L g839 ( 
.A(n_764),
.Y(n_839)
);

CKINVDCx5p33_ASAP7_75t_R g840 ( 
.A(n_807),
.Y(n_840)
);

OR2x2_ASAP7_75t_L g841 ( 
.A(n_518),
.B(n_0),
.Y(n_841)
);

INVxp67_ASAP7_75t_L g842 ( 
.A(n_527),
.Y(n_842)
);

INVx2_ASAP7_75t_L g843 ( 
.A(n_532),
.Y(n_843)
);

INVx1_ASAP7_75t_L g844 ( 
.A(n_764),
.Y(n_844)
);

CKINVDCx5p33_ASAP7_75t_R g845 ( 
.A(n_540),
.Y(n_845)
);

INVx2_ASAP7_75t_L g846 ( 
.A(n_532),
.Y(n_846)
);

INVx1_ASAP7_75t_L g847 ( 
.A(n_817),
.Y(n_847)
);

CKINVDCx14_ASAP7_75t_R g848 ( 
.A(n_786),
.Y(n_848)
);

INVxp33_ASAP7_75t_SL g849 ( 
.A(n_482),
.Y(n_849)
);

INVx1_ASAP7_75t_L g850 ( 
.A(n_817),
.Y(n_850)
);

INVx1_ASAP7_75t_L g851 ( 
.A(n_532),
.Y(n_851)
);

INVxp67_ASAP7_75t_SL g852 ( 
.A(n_489),
.Y(n_852)
);

INVxp67_ASAP7_75t_SL g853 ( 
.A(n_513),
.Y(n_853)
);

INVx1_ASAP7_75t_L g854 ( 
.A(n_473),
.Y(n_854)
);

INVx1_ASAP7_75t_L g855 ( 
.A(n_478),
.Y(n_855)
);

BUFx6f_ASAP7_75t_L g856 ( 
.A(n_652),
.Y(n_856)
);

CKINVDCx20_ASAP7_75t_R g857 ( 
.A(n_564),
.Y(n_857)
);

INVx1_ASAP7_75t_L g858 ( 
.A(n_488),
.Y(n_858)
);

INVx1_ASAP7_75t_L g859 ( 
.A(n_529),
.Y(n_859)
);

INVxp67_ASAP7_75t_SL g860 ( 
.A(n_590),
.Y(n_860)
);

INVx1_ASAP7_75t_L g861 ( 
.A(n_541),
.Y(n_861)
);

INVx1_ASAP7_75t_L g862 ( 
.A(n_553),
.Y(n_862)
);

INVx1_ASAP7_75t_L g863 ( 
.A(n_567),
.Y(n_863)
);

BUFx6f_ASAP7_75t_L g864 ( 
.A(n_652),
.Y(n_864)
);

INVx1_ASAP7_75t_SL g865 ( 
.A(n_627),
.Y(n_865)
);

INVxp33_ASAP7_75t_SL g866 ( 
.A(n_482),
.Y(n_866)
);

NOR2xp33_ASAP7_75t_L g867 ( 
.A(n_485),
.B(n_1),
.Y(n_867)
);

INVx2_ASAP7_75t_L g868 ( 
.A(n_487),
.Y(n_868)
);

INVx1_ASAP7_75t_L g869 ( 
.A(n_569),
.Y(n_869)
);

INVx1_ASAP7_75t_L g870 ( 
.A(n_599),
.Y(n_870)
);

CKINVDCx5p33_ASAP7_75t_R g871 ( 
.A(n_548),
.Y(n_871)
);

INVx1_ASAP7_75t_L g872 ( 
.A(n_621),
.Y(n_872)
);

HB1xp67_ASAP7_75t_L g873 ( 
.A(n_497),
.Y(n_873)
);

INVxp67_ASAP7_75t_SL g874 ( 
.A(n_630),
.Y(n_874)
);

INVx1_ASAP7_75t_L g875 ( 
.A(n_625),
.Y(n_875)
);

INVx1_ASAP7_75t_L g876 ( 
.A(n_626),
.Y(n_876)
);

CKINVDCx16_ASAP7_75t_R g877 ( 
.A(n_544),
.Y(n_877)
);

INVx2_ASAP7_75t_L g878 ( 
.A(n_487),
.Y(n_878)
);

INVx1_ASAP7_75t_L g879 ( 
.A(n_633),
.Y(n_879)
);

HB1xp67_ASAP7_75t_L g880 ( 
.A(n_614),
.Y(n_880)
);

CKINVDCx5p33_ASAP7_75t_R g881 ( 
.A(n_552),
.Y(n_881)
);

INVx1_ASAP7_75t_L g882 ( 
.A(n_653),
.Y(n_882)
);

INVx1_ASAP7_75t_L g883 ( 
.A(n_654),
.Y(n_883)
);

CKINVDCx5p33_ASAP7_75t_R g884 ( 
.A(n_555),
.Y(n_884)
);

INVx1_ASAP7_75t_L g885 ( 
.A(n_663),
.Y(n_885)
);

HB1xp67_ASAP7_75t_L g886 ( 
.A(n_823),
.Y(n_886)
);

INVx1_ASAP7_75t_L g887 ( 
.A(n_668),
.Y(n_887)
);

INVx1_ASAP7_75t_L g888 ( 
.A(n_687),
.Y(n_888)
);

CKINVDCx5p33_ASAP7_75t_R g889 ( 
.A(n_556),
.Y(n_889)
);

INVx2_ASAP7_75t_L g890 ( 
.A(n_523),
.Y(n_890)
);

INVxp33_ASAP7_75t_SL g891 ( 
.A(n_499),
.Y(n_891)
);

INVxp33_ASAP7_75t_SL g892 ( 
.A(n_499),
.Y(n_892)
);

INVxp67_ASAP7_75t_L g893 ( 
.A(n_701),
.Y(n_893)
);

BUFx6f_ASAP7_75t_L g894 ( 
.A(n_652),
.Y(n_894)
);

INVx1_ASAP7_75t_L g895 ( 
.A(n_697),
.Y(n_895)
);

CKINVDCx5p33_ASAP7_75t_R g896 ( 
.A(n_558),
.Y(n_896)
);

INVx1_ASAP7_75t_L g897 ( 
.A(n_698),
.Y(n_897)
);

INVx1_ASAP7_75t_L g898 ( 
.A(n_713),
.Y(n_898)
);

CKINVDCx14_ASAP7_75t_R g899 ( 
.A(n_605),
.Y(n_899)
);

INVx1_ASAP7_75t_L g900 ( 
.A(n_715),
.Y(n_900)
);

INVx1_ASAP7_75t_L g901 ( 
.A(n_719),
.Y(n_901)
);

INVx1_ASAP7_75t_L g902 ( 
.A(n_730),
.Y(n_902)
);

INVxp67_ASAP7_75t_SL g903 ( 
.A(n_470),
.Y(n_903)
);

INVx1_ASAP7_75t_L g904 ( 
.A(n_732),
.Y(n_904)
);

BUFx3_ASAP7_75t_L g905 ( 
.A(n_470),
.Y(n_905)
);

INVxp33_ASAP7_75t_SL g906 ( 
.A(n_500),
.Y(n_906)
);

INVx1_ASAP7_75t_L g907 ( 
.A(n_739),
.Y(n_907)
);

INVx1_ASAP7_75t_L g908 ( 
.A(n_741),
.Y(n_908)
);

INVxp33_ASAP7_75t_SL g909 ( 
.A(n_500),
.Y(n_909)
);

INVxp67_ASAP7_75t_SL g910 ( 
.A(n_486),
.Y(n_910)
);

INVxp67_ASAP7_75t_SL g911 ( 
.A(n_486),
.Y(n_911)
);

INVx1_ASAP7_75t_L g912 ( 
.A(n_755),
.Y(n_912)
);

INVx1_ASAP7_75t_SL g913 ( 
.A(n_576),
.Y(n_913)
);

INVx1_ASAP7_75t_L g914 ( 
.A(n_762),
.Y(n_914)
);

INVx1_ASAP7_75t_L g915 ( 
.A(n_768),
.Y(n_915)
);

INVx2_ASAP7_75t_L g916 ( 
.A(n_523),
.Y(n_916)
);

INVx1_ASAP7_75t_L g917 ( 
.A(n_770),
.Y(n_917)
);

INVxp67_ASAP7_75t_L g918 ( 
.A(n_623),
.Y(n_918)
);

INVx1_ASAP7_75t_L g919 ( 
.A(n_801),
.Y(n_919)
);

INVx1_ASAP7_75t_L g920 ( 
.A(n_804),
.Y(n_920)
);

INVx1_ASAP7_75t_L g921 ( 
.A(n_810),
.Y(n_921)
);

CKINVDCx20_ASAP7_75t_R g922 ( 
.A(n_580),
.Y(n_922)
);

INVx1_ASAP7_75t_L g923 ( 
.A(n_812),
.Y(n_923)
);

INVx2_ASAP7_75t_L g924 ( 
.A(n_543),
.Y(n_924)
);

INVx1_ASAP7_75t_L g925 ( 
.A(n_824),
.Y(n_925)
);

INVx1_ASAP7_75t_L g926 ( 
.A(n_495),
.Y(n_926)
);

INVx1_ASAP7_75t_L g927 ( 
.A(n_495),
.Y(n_927)
);

INVx1_ASAP7_75t_L g928 ( 
.A(n_624),
.Y(n_928)
);

CKINVDCx5p33_ASAP7_75t_R g929 ( 
.A(n_562),
.Y(n_929)
);

CKINVDCx5p33_ASAP7_75t_R g930 ( 
.A(n_565),
.Y(n_930)
);

INVxp33_ASAP7_75t_L g931 ( 
.A(n_543),
.Y(n_931)
);

INVx1_ASAP7_75t_L g932 ( 
.A(n_624),
.Y(n_932)
);

INVxp67_ASAP7_75t_L g933 ( 
.A(n_623),
.Y(n_933)
);

INVx2_ASAP7_75t_L g934 ( 
.A(n_594),
.Y(n_934)
);

INVx1_ASAP7_75t_SL g935 ( 
.A(n_646),
.Y(n_935)
);

INVx1_ASAP7_75t_L g936 ( 
.A(n_673),
.Y(n_936)
);

INVx1_ASAP7_75t_L g937 ( 
.A(n_673),
.Y(n_937)
);

CKINVDCx14_ASAP7_75t_R g938 ( 
.A(n_605),
.Y(n_938)
);

INVx1_ASAP7_75t_L g939 ( 
.A(n_792),
.Y(n_939)
);

INVx1_ASAP7_75t_L g940 ( 
.A(n_792),
.Y(n_940)
);

INVxp67_ASAP7_75t_L g941 ( 
.A(n_623),
.Y(n_941)
);

INVx2_ASAP7_75t_L g942 ( 
.A(n_594),
.Y(n_942)
);

INVx1_ASAP7_75t_L g943 ( 
.A(n_475),
.Y(n_943)
);

INVxp33_ASAP7_75t_L g944 ( 
.A(n_644),
.Y(n_944)
);

INVx1_ASAP7_75t_L g945 ( 
.A(n_479),
.Y(n_945)
);

INVx1_ASAP7_75t_L g946 ( 
.A(n_484),
.Y(n_946)
);

INVxp33_ASAP7_75t_SL g947 ( 
.A(n_502),
.Y(n_947)
);

INVx1_ASAP7_75t_L g948 ( 
.A(n_490),
.Y(n_948)
);

INVx1_ASAP7_75t_L g949 ( 
.A(n_493),
.Y(n_949)
);

INVx2_ASAP7_75t_L g950 ( 
.A(n_644),
.Y(n_950)
);

NOR2xp67_ASAP7_75t_L g951 ( 
.A(n_781),
.B(n_1),
.Y(n_951)
);

INVx1_ASAP7_75t_L g952 ( 
.A(n_521),
.Y(n_952)
);

BUFx3_ASAP7_75t_L g953 ( 
.A(n_605),
.Y(n_953)
);

INVx1_ASAP7_75t_L g954 ( 
.A(n_522),
.Y(n_954)
);

CKINVDCx5p33_ASAP7_75t_R g955 ( 
.A(n_568),
.Y(n_955)
);

CKINVDCx5p33_ASAP7_75t_R g956 ( 
.A(n_570),
.Y(n_956)
);

INVxp67_ASAP7_75t_SL g957 ( 
.A(n_781),
.Y(n_957)
);

INVx1_ASAP7_75t_L g958 ( 
.A(n_538),
.Y(n_958)
);

INVx1_ASAP7_75t_L g959 ( 
.A(n_554),
.Y(n_959)
);

INVx1_ASAP7_75t_L g960 ( 
.A(n_559),
.Y(n_960)
);

INVx1_ASAP7_75t_L g961 ( 
.A(n_560),
.Y(n_961)
);

CKINVDCx5p33_ASAP7_75t_R g962 ( 
.A(n_571),
.Y(n_962)
);

BUFx2_ASAP7_75t_L g963 ( 
.A(n_502),
.Y(n_963)
);

INVx1_ASAP7_75t_L g964 ( 
.A(n_563),
.Y(n_964)
);

BUFx6f_ASAP7_75t_L g965 ( 
.A(n_652),
.Y(n_965)
);

INVx1_ASAP7_75t_L g966 ( 
.A(n_566),
.Y(n_966)
);

CKINVDCx5p33_ASAP7_75t_R g967 ( 
.A(n_573),
.Y(n_967)
);

CKINVDCx5p33_ASAP7_75t_R g968 ( 
.A(n_581),
.Y(n_968)
);

INVxp67_ASAP7_75t_SL g969 ( 
.A(n_781),
.Y(n_969)
);

CKINVDCx20_ASAP7_75t_R g970 ( 
.A(n_659),
.Y(n_970)
);

INVx1_ASAP7_75t_L g971 ( 
.A(n_572),
.Y(n_971)
);

INVx2_ASAP7_75t_L g972 ( 
.A(n_656),
.Y(n_972)
);

INVx1_ASAP7_75t_SL g973 ( 
.A(n_664),
.Y(n_973)
);

CKINVDCx5p33_ASAP7_75t_R g974 ( 
.A(n_582),
.Y(n_974)
);

INVx1_ASAP7_75t_L g975 ( 
.A(n_574),
.Y(n_975)
);

CKINVDCx16_ASAP7_75t_R g976 ( 
.A(n_584),
.Y(n_976)
);

INVx1_ASAP7_75t_L g977 ( 
.A(n_595),
.Y(n_977)
);

INVx1_ASAP7_75t_L g978 ( 
.A(n_596),
.Y(n_978)
);

INVx1_ASAP7_75t_L g979 ( 
.A(n_600),
.Y(n_979)
);

INVx1_ASAP7_75t_L g980 ( 
.A(n_603),
.Y(n_980)
);

INVx2_ASAP7_75t_L g981 ( 
.A(n_656),
.Y(n_981)
);

INVx1_ASAP7_75t_L g982 ( 
.A(n_610),
.Y(n_982)
);

INVxp33_ASAP7_75t_SL g983 ( 
.A(n_504),
.Y(n_983)
);

INVx1_ASAP7_75t_L g984 ( 
.A(n_618),
.Y(n_984)
);

INVx1_ASAP7_75t_L g985 ( 
.A(n_628),
.Y(n_985)
);

INVx1_ASAP7_75t_L g986 ( 
.A(n_629),
.Y(n_986)
);

CKINVDCx20_ASAP7_75t_R g987 ( 
.A(n_666),
.Y(n_987)
);

INVx1_ASAP7_75t_SL g988 ( 
.A(n_692),
.Y(n_988)
);

INVx1_ASAP7_75t_L g989 ( 
.A(n_634),
.Y(n_989)
);

INVx1_ASAP7_75t_SL g990 ( 
.A(n_737),
.Y(n_990)
);

INVx1_ASAP7_75t_L g991 ( 
.A(n_638),
.Y(n_991)
);

INVx1_ASAP7_75t_L g992 ( 
.A(n_639),
.Y(n_992)
);

INVx1_ASAP7_75t_L g993 ( 
.A(n_648),
.Y(n_993)
);

INVx1_ASAP7_75t_L g994 ( 
.A(n_649),
.Y(n_994)
);

INVx1_ASAP7_75t_L g995 ( 
.A(n_658),
.Y(n_995)
);

INVxp33_ASAP7_75t_SL g996 ( 
.A(n_504),
.Y(n_996)
);

INVxp33_ASAP7_75t_SL g997 ( 
.A(n_508),
.Y(n_997)
);

INVx1_ASAP7_75t_L g998 ( 
.A(n_660),
.Y(n_998)
);

INVxp67_ASAP7_75t_L g999 ( 
.A(n_632),
.Y(n_999)
);

INVx1_ASAP7_75t_L g1000 ( 
.A(n_661),
.Y(n_1000)
);

INVx1_ASAP7_75t_L g1001 ( 
.A(n_672),
.Y(n_1001)
);

INVxp67_ASAP7_75t_SL g1002 ( 
.A(n_680),
.Y(n_1002)
);

INVx1_ASAP7_75t_L g1003 ( 
.A(n_683),
.Y(n_1003)
);

INVx1_ASAP7_75t_L g1004 ( 
.A(n_690),
.Y(n_1004)
);

CKINVDCx20_ASAP7_75t_R g1005 ( 
.A(n_805),
.Y(n_1005)
);

INVx1_ASAP7_75t_L g1006 ( 
.A(n_694),
.Y(n_1006)
);

INVxp67_ASAP7_75t_L g1007 ( 
.A(n_632),
.Y(n_1007)
);

BUFx2_ASAP7_75t_L g1008 ( 
.A(n_508),
.Y(n_1008)
);

INVx1_ASAP7_75t_L g1009 ( 
.A(n_695),
.Y(n_1009)
);

CKINVDCx20_ASAP7_75t_R g1010 ( 
.A(n_811),
.Y(n_1010)
);

CKINVDCx14_ASAP7_75t_R g1011 ( 
.A(n_647),
.Y(n_1011)
);

INVx1_ASAP7_75t_L g1012 ( 
.A(n_696),
.Y(n_1012)
);

INVx1_ASAP7_75t_L g1013 ( 
.A(n_700),
.Y(n_1013)
);

INVx1_ASAP7_75t_L g1014 ( 
.A(n_706),
.Y(n_1014)
);

INVx1_ASAP7_75t_L g1015 ( 
.A(n_707),
.Y(n_1015)
);

BUFx3_ASAP7_75t_L g1016 ( 
.A(n_647),
.Y(n_1016)
);

INVx1_ASAP7_75t_SL g1017 ( 
.A(n_815),
.Y(n_1017)
);

INVxp67_ASAP7_75t_SL g1018 ( 
.A(n_709),
.Y(n_1018)
);

CKINVDCx20_ASAP7_75t_R g1019 ( 
.A(n_820),
.Y(n_1019)
);

CKINVDCx5p33_ASAP7_75t_R g1020 ( 
.A(n_589),
.Y(n_1020)
);

INVx1_ASAP7_75t_L g1021 ( 
.A(n_718),
.Y(n_1021)
);

INVx1_ASAP7_75t_L g1022 ( 
.A(n_724),
.Y(n_1022)
);

INVx1_ASAP7_75t_L g1023 ( 
.A(n_725),
.Y(n_1023)
);

INVx1_ASAP7_75t_L g1024 ( 
.A(n_735),
.Y(n_1024)
);

INVx1_ASAP7_75t_L g1025 ( 
.A(n_736),
.Y(n_1025)
);

INVx1_ASAP7_75t_L g1026 ( 
.A(n_738),
.Y(n_1026)
);

CKINVDCx20_ASAP7_75t_R g1027 ( 
.A(n_511),
.Y(n_1027)
);

INVx1_ASAP7_75t_L g1028 ( 
.A(n_744),
.Y(n_1028)
);

INVxp67_ASAP7_75t_SL g1029 ( 
.A(n_747),
.Y(n_1029)
);

INVx1_ASAP7_75t_L g1030 ( 
.A(n_753),
.Y(n_1030)
);

INVx1_ASAP7_75t_L g1031 ( 
.A(n_756),
.Y(n_1031)
);

INVx1_ASAP7_75t_L g1032 ( 
.A(n_765),
.Y(n_1032)
);

INVx2_ASAP7_75t_L g1033 ( 
.A(n_711),
.Y(n_1033)
);

CKINVDCx20_ASAP7_75t_R g1034 ( 
.A(n_511),
.Y(n_1034)
);

INVx2_ASAP7_75t_SL g1035 ( 
.A(n_632),
.Y(n_1035)
);

INVx1_ASAP7_75t_L g1036 ( 
.A(n_775),
.Y(n_1036)
);

INVx1_ASAP7_75t_L g1037 ( 
.A(n_778),
.Y(n_1037)
);

INVx1_ASAP7_75t_L g1038 ( 
.A(n_795),
.Y(n_1038)
);

INVx2_ASAP7_75t_L g1039 ( 
.A(n_711),
.Y(n_1039)
);

INVx1_ASAP7_75t_L g1040 ( 
.A(n_797),
.Y(n_1040)
);

INVxp33_ASAP7_75t_SL g1041 ( 
.A(n_515),
.Y(n_1041)
);

INVxp67_ASAP7_75t_L g1042 ( 
.A(n_643),
.Y(n_1042)
);

INVx2_ASAP7_75t_L g1043 ( 
.A(n_729),
.Y(n_1043)
);

INVx1_ASAP7_75t_L g1044 ( 
.A(n_806),
.Y(n_1044)
);

INVx2_ASAP7_75t_L g1045 ( 
.A(n_729),
.Y(n_1045)
);

HB1xp67_ASAP7_75t_L g1046 ( 
.A(n_515),
.Y(n_1046)
);

INVx1_ASAP7_75t_L g1047 ( 
.A(n_477),
.Y(n_1047)
);

INVx2_ASAP7_75t_L g1048 ( 
.A(n_652),
.Y(n_1048)
);

INVx1_ASAP7_75t_L g1049 ( 
.A(n_477),
.Y(n_1049)
);

CKINVDCx14_ASAP7_75t_R g1050 ( 
.A(n_647),
.Y(n_1050)
);

INVx1_ASAP7_75t_L g1051 ( 
.A(n_491),
.Y(n_1051)
);

INVx1_ASAP7_75t_L g1052 ( 
.A(n_491),
.Y(n_1052)
);

INVx1_ASAP7_75t_L g1053 ( 
.A(n_549),
.Y(n_1053)
);

INVx1_ASAP7_75t_L g1054 ( 
.A(n_549),
.Y(n_1054)
);

INVx1_ASAP7_75t_L g1055 ( 
.A(n_575),
.Y(n_1055)
);

CKINVDCx5p33_ASAP7_75t_R g1056 ( 
.A(n_591),
.Y(n_1056)
);

INVx1_ASAP7_75t_L g1057 ( 
.A(n_575),
.Y(n_1057)
);

CKINVDCx5p33_ASAP7_75t_R g1058 ( 
.A(n_592),
.Y(n_1058)
);

INVxp67_ASAP7_75t_L g1059 ( 
.A(n_643),
.Y(n_1059)
);

INVx1_ASAP7_75t_L g1060 ( 
.A(n_669),
.Y(n_1060)
);

BUFx3_ASAP7_75t_L g1061 ( 
.A(n_651),
.Y(n_1061)
);

INVx1_ASAP7_75t_L g1062 ( 
.A(n_669),
.Y(n_1062)
);

INVx1_ASAP7_75t_L g1063 ( 
.A(n_681),
.Y(n_1063)
);

CKINVDCx5p33_ASAP7_75t_R g1064 ( 
.A(n_602),
.Y(n_1064)
);

INVx1_ASAP7_75t_L g1065 ( 
.A(n_681),
.Y(n_1065)
);

INVxp33_ASAP7_75t_L g1066 ( 
.A(n_686),
.Y(n_1066)
);

INVx1_ASAP7_75t_L g1067 ( 
.A(n_686),
.Y(n_1067)
);

INVx1_ASAP7_75t_L g1068 ( 
.A(n_693),
.Y(n_1068)
);

INVx1_ASAP7_75t_L g1069 ( 
.A(n_693),
.Y(n_1069)
);

CKINVDCx20_ASAP7_75t_R g1070 ( 
.A(n_516),
.Y(n_1070)
);

INVxp67_ASAP7_75t_SL g1071 ( 
.A(n_731),
.Y(n_1071)
);

INVx2_ASAP7_75t_L g1072 ( 
.A(n_754),
.Y(n_1072)
);

INVx1_ASAP7_75t_L g1073 ( 
.A(n_731),
.Y(n_1073)
);

INVx1_ASAP7_75t_L g1074 ( 
.A(n_813),
.Y(n_1074)
);

INVx1_ASAP7_75t_L g1075 ( 
.A(n_813),
.Y(n_1075)
);

BUFx2_ASAP7_75t_L g1076 ( 
.A(n_516),
.Y(n_1076)
);

INVx1_ASAP7_75t_L g1077 ( 
.A(n_539),
.Y(n_1077)
);

CKINVDCx20_ASAP7_75t_R g1078 ( 
.A(n_519),
.Y(n_1078)
);

INVx1_ASAP7_75t_L g1079 ( 
.A(n_539),
.Y(n_1079)
);

INVx1_ASAP7_75t_L g1080 ( 
.A(n_545),
.Y(n_1080)
);

INVx1_ASAP7_75t_L g1081 ( 
.A(n_545),
.Y(n_1081)
);

INVxp33_ASAP7_75t_L g1082 ( 
.A(n_754),
.Y(n_1082)
);

BUFx6f_ASAP7_75t_SL g1083 ( 
.A(n_643),
.Y(n_1083)
);

INVx1_ASAP7_75t_L g1084 ( 
.A(n_674),
.Y(n_1084)
);

INVxp67_ASAP7_75t_SL g1085 ( 
.A(n_761),
.Y(n_1085)
);

INVxp33_ASAP7_75t_SL g1086 ( 
.A(n_519),
.Y(n_1086)
);

CKINVDCx5p33_ASAP7_75t_R g1087 ( 
.A(n_604),
.Y(n_1087)
);

INVx1_ASAP7_75t_L g1088 ( 
.A(n_674),
.Y(n_1088)
);

BUFx6f_ASAP7_75t_L g1089 ( 
.A(n_754),
.Y(n_1089)
);

BUFx6f_ASAP7_75t_L g1090 ( 
.A(n_754),
.Y(n_1090)
);

BUFx6f_ASAP7_75t_L g1091 ( 
.A(n_754),
.Y(n_1091)
);

INVx1_ASAP7_75t_L g1092 ( 
.A(n_688),
.Y(n_1092)
);

INVx1_ASAP7_75t_L g1093 ( 
.A(n_688),
.Y(n_1093)
);

INVx1_ASAP7_75t_L g1094 ( 
.A(n_688),
.Y(n_1094)
);

CKINVDCx5p33_ASAP7_75t_R g1095 ( 
.A(n_613),
.Y(n_1095)
);

INVx1_ASAP7_75t_L g1096 ( 
.A(n_758),
.Y(n_1096)
);

INVxp67_ASAP7_75t_SL g1097 ( 
.A(n_791),
.Y(n_1097)
);

INVx1_ASAP7_75t_L g1098 ( 
.A(n_758),
.Y(n_1098)
);

INVx1_ASAP7_75t_L g1099 ( 
.A(n_758),
.Y(n_1099)
);

INVx1_ASAP7_75t_L g1100 ( 
.A(n_609),
.Y(n_1100)
);

INVx1_ASAP7_75t_L g1101 ( 
.A(n_507),
.Y(n_1101)
);

BUFx5_ASAP7_75t_L g1102 ( 
.A(n_651),
.Y(n_1102)
);

INVxp67_ASAP7_75t_L g1103 ( 
.A(n_826),
.Y(n_1103)
);

INVx1_ASAP7_75t_L g1104 ( 
.A(n_507),
.Y(n_1104)
);

INVx1_ASAP7_75t_L g1105 ( 
.A(n_546),
.Y(n_1105)
);

INVxp33_ASAP7_75t_SL g1106 ( 
.A(n_524),
.Y(n_1106)
);

INVxp67_ASAP7_75t_L g1107 ( 
.A(n_826),
.Y(n_1107)
);

CKINVDCx5p33_ASAP7_75t_R g1108 ( 
.A(n_616),
.Y(n_1108)
);

INVx1_ASAP7_75t_L g1109 ( 
.A(n_550),
.Y(n_1109)
);

INVx1_ASAP7_75t_L g1110 ( 
.A(n_551),
.Y(n_1110)
);

INVxp33_ASAP7_75t_L g1111 ( 
.A(n_524),
.Y(n_1111)
);

INVx1_ASAP7_75t_L g1112 ( 
.A(n_557),
.Y(n_1112)
);

INVx1_ASAP7_75t_L g1113 ( 
.A(n_561),
.Y(n_1113)
);

NAND2xp5_ASAP7_75t_L g1114 ( 
.A(n_845),
.B(n_871),
.Y(n_1114)
);

NAND2xp5_ASAP7_75t_L g1115 ( 
.A(n_881),
.B(n_617),
.Y(n_1115)
);

BUFx6f_ASAP7_75t_L g1116 ( 
.A(n_856),
.Y(n_1116)
);

AND2x4_ASAP7_75t_L g1117 ( 
.A(n_957),
.B(n_597),
.Y(n_1117)
);

INVx1_ASAP7_75t_L g1118 ( 
.A(n_851),
.Y(n_1118)
);

BUFx12f_ASAP7_75t_L g1119 ( 
.A(n_840),
.Y(n_1119)
);

INVx1_ASAP7_75t_L g1120 ( 
.A(n_831),
.Y(n_1120)
);

BUFx2_ASAP7_75t_L g1121 ( 
.A(n_1027),
.Y(n_1121)
);

AND2x2_ASAP7_75t_L g1122 ( 
.A(n_836),
.B(n_615),
.Y(n_1122)
);

HB1xp67_ASAP7_75t_L g1123 ( 
.A(n_873),
.Y(n_1123)
);

INVx2_ASAP7_75t_L g1124 ( 
.A(n_831),
.Y(n_1124)
);

INVx2_ASAP7_75t_L g1125 ( 
.A(n_834),
.Y(n_1125)
);

INVx2_ASAP7_75t_SL g1126 ( 
.A(n_953),
.Y(n_1126)
);

BUFx6f_ASAP7_75t_L g1127 ( 
.A(n_856),
.Y(n_1127)
);

INVx2_ASAP7_75t_L g1128 ( 
.A(n_834),
.Y(n_1128)
);

INVx1_ASAP7_75t_L g1129 ( 
.A(n_843),
.Y(n_1129)
);

INVx1_ASAP7_75t_L g1130 ( 
.A(n_843),
.Y(n_1130)
);

AND2x4_ASAP7_75t_L g1131 ( 
.A(n_969),
.B(n_733),
.Y(n_1131)
);

OAI22x1_ASAP7_75t_L g1132 ( 
.A1(n_865),
.A2(n_526),
.B1(n_528),
.B2(n_525),
.Y(n_1132)
);

NAND2xp5_ASAP7_75t_L g1133 ( 
.A(n_884),
.B(n_889),
.Y(n_1133)
);

NAND2xp5_ASAP7_75t_L g1134 ( 
.A(n_896),
.B(n_619),
.Y(n_1134)
);

INVx2_ASAP7_75t_L g1135 ( 
.A(n_846),
.Y(n_1135)
);

BUFx12f_ASAP7_75t_L g1136 ( 
.A(n_929),
.Y(n_1136)
);

CKINVDCx16_ASAP7_75t_R g1137 ( 
.A(n_877),
.Y(n_1137)
);

NOR2xp33_ASAP7_75t_L g1138 ( 
.A(n_1066),
.B(n_794),
.Y(n_1138)
);

OAI22xp5_ASAP7_75t_L g1139 ( 
.A1(n_852),
.A2(n_526),
.B1(n_528),
.B2(n_525),
.Y(n_1139)
);

BUFx3_ASAP7_75t_L g1140 ( 
.A(n_905),
.Y(n_1140)
);

INVx1_ASAP7_75t_L g1141 ( 
.A(n_846),
.Y(n_1141)
);

BUFx3_ASAP7_75t_L g1142 ( 
.A(n_905),
.Y(n_1142)
);

BUFx2_ASAP7_75t_L g1143 ( 
.A(n_1027),
.Y(n_1143)
);

NOR2xp33_ASAP7_75t_L g1144 ( 
.A(n_1066),
.B(n_472),
.Y(n_1144)
);

INVx2_ASAP7_75t_L g1145 ( 
.A(n_1048),
.Y(n_1145)
);

INVx4_ASAP7_75t_L g1146 ( 
.A(n_864),
.Y(n_1146)
);

HB1xp67_ASAP7_75t_L g1147 ( 
.A(n_880),
.Y(n_1147)
);

BUFx3_ASAP7_75t_L g1148 ( 
.A(n_926),
.Y(n_1148)
);

BUFx6f_ASAP7_75t_L g1149 ( 
.A(n_864),
.Y(n_1149)
);

AND2x2_ASAP7_75t_L g1150 ( 
.A(n_903),
.B(n_651),
.Y(n_1150)
);

INVx2_ASAP7_75t_L g1151 ( 
.A(n_1048),
.Y(n_1151)
);

INVx2_ASAP7_75t_L g1152 ( 
.A(n_1072),
.Y(n_1152)
);

CKINVDCx5p33_ASAP7_75t_R g1153 ( 
.A(n_930),
.Y(n_1153)
);

INVx2_ASAP7_75t_L g1154 ( 
.A(n_1072),
.Y(n_1154)
);

INVx1_ASAP7_75t_L g1155 ( 
.A(n_943),
.Y(n_1155)
);

AND2x4_ASAP7_75t_L g1156 ( 
.A(n_1002),
.B(n_825),
.Y(n_1156)
);

AND2x2_ASAP7_75t_L g1157 ( 
.A(n_836),
.B(n_657),
.Y(n_1157)
);

BUFx3_ASAP7_75t_L g1158 ( 
.A(n_927),
.Y(n_1158)
);

AND2x2_ASAP7_75t_L g1159 ( 
.A(n_848),
.B(n_657),
.Y(n_1159)
);

BUFx2_ASAP7_75t_L g1160 ( 
.A(n_1034),
.Y(n_1160)
);

INVx1_ASAP7_75t_L g1161 ( 
.A(n_945),
.Y(n_1161)
);

OAI22x1_ASAP7_75t_R g1162 ( 
.A1(n_857),
.A2(n_970),
.B1(n_987),
.B2(n_922),
.Y(n_1162)
);

AND2x6_ASAP7_75t_L g1163 ( 
.A(n_894),
.B(n_607),
.Y(n_1163)
);

INVxp33_ASAP7_75t_L g1164 ( 
.A(n_886),
.Y(n_1164)
);

OA22x2_ASAP7_75t_SL g1165 ( 
.A1(n_853),
.A2(n_860),
.B1(n_874),
.B2(n_830),
.Y(n_1165)
);

OA21x2_ASAP7_75t_L g1166 ( 
.A1(n_1047),
.A2(n_578),
.B(n_577),
.Y(n_1166)
);

BUFx6f_ASAP7_75t_L g1167 ( 
.A(n_894),
.Y(n_1167)
);

INVx1_ASAP7_75t_L g1168 ( 
.A(n_946),
.Y(n_1168)
);

CKINVDCx6p67_ASAP7_75t_R g1169 ( 
.A(n_1083),
.Y(n_1169)
);

BUFx3_ASAP7_75t_L g1170 ( 
.A(n_928),
.Y(n_1170)
);

CKINVDCx5p33_ASAP7_75t_R g1171 ( 
.A(n_955),
.Y(n_1171)
);

BUFx6f_ASAP7_75t_L g1172 ( 
.A(n_894),
.Y(n_1172)
);

BUFx6f_ASAP7_75t_L g1173 ( 
.A(n_965),
.Y(n_1173)
);

INVx1_ASAP7_75t_L g1174 ( 
.A(n_948),
.Y(n_1174)
);

CKINVDCx5p33_ASAP7_75t_R g1175 ( 
.A(n_956),
.Y(n_1175)
);

INVx1_ASAP7_75t_L g1176 ( 
.A(n_949),
.Y(n_1176)
);

BUFx2_ASAP7_75t_L g1177 ( 
.A(n_1034),
.Y(n_1177)
);

INVx2_ASAP7_75t_L g1178 ( 
.A(n_965),
.Y(n_1178)
);

INVx1_ASAP7_75t_L g1179 ( 
.A(n_952),
.Y(n_1179)
);

CKINVDCx14_ASAP7_75t_R g1180 ( 
.A(n_899),
.Y(n_1180)
);

BUFx6f_ASAP7_75t_L g1181 ( 
.A(n_965),
.Y(n_1181)
);

BUFx6f_ASAP7_75t_L g1182 ( 
.A(n_965),
.Y(n_1182)
);

AND2x2_ASAP7_75t_L g1183 ( 
.A(n_848),
.B(n_657),
.Y(n_1183)
);

INVx2_ASAP7_75t_L g1184 ( 
.A(n_1089),
.Y(n_1184)
);

BUFx12f_ASAP7_75t_L g1185 ( 
.A(n_962),
.Y(n_1185)
);

HB1xp67_ASAP7_75t_L g1186 ( 
.A(n_913),
.Y(n_1186)
);

BUFx3_ASAP7_75t_L g1187 ( 
.A(n_932),
.Y(n_1187)
);

OA21x2_ASAP7_75t_L g1188 ( 
.A1(n_1049),
.A2(n_585),
.B(n_583),
.Y(n_1188)
);

INVx2_ASAP7_75t_L g1189 ( 
.A(n_1089),
.Y(n_1189)
);

BUFx12f_ASAP7_75t_L g1190 ( 
.A(n_967),
.Y(n_1190)
);

INVx3_ASAP7_75t_L g1191 ( 
.A(n_1089),
.Y(n_1191)
);

BUFx6f_ASAP7_75t_L g1192 ( 
.A(n_1089),
.Y(n_1192)
);

BUFx6f_ASAP7_75t_L g1193 ( 
.A(n_1090),
.Y(n_1193)
);

BUFx3_ASAP7_75t_L g1194 ( 
.A(n_936),
.Y(n_1194)
);

BUFx12f_ASAP7_75t_L g1195 ( 
.A(n_968),
.Y(n_1195)
);

AND2x2_ASAP7_75t_L g1196 ( 
.A(n_910),
.B(n_472),
.Y(n_1196)
);

BUFx2_ASAP7_75t_L g1197 ( 
.A(n_1070),
.Y(n_1197)
);

NAND2xp5_ASAP7_75t_L g1198 ( 
.A(n_974),
.B(n_622),
.Y(n_1198)
);

INVx3_ASAP7_75t_L g1199 ( 
.A(n_1090),
.Y(n_1199)
);

BUFx2_ASAP7_75t_L g1200 ( 
.A(n_1070),
.Y(n_1200)
);

AND2x2_ASAP7_75t_L g1201 ( 
.A(n_911),
.B(n_480),
.Y(n_1201)
);

INVx1_ASAP7_75t_L g1202 ( 
.A(n_954),
.Y(n_1202)
);

BUFx6f_ASAP7_75t_L g1203 ( 
.A(n_1090),
.Y(n_1203)
);

INVx1_ASAP7_75t_L g1204 ( 
.A(n_958),
.Y(n_1204)
);

AND2x2_ASAP7_75t_L g1205 ( 
.A(n_899),
.B(n_480),
.Y(n_1205)
);

BUFx6f_ASAP7_75t_L g1206 ( 
.A(n_1091),
.Y(n_1206)
);

HB1xp67_ASAP7_75t_L g1207 ( 
.A(n_935),
.Y(n_1207)
);

INVx1_ASAP7_75t_L g1208 ( 
.A(n_959),
.Y(n_1208)
);

BUFx12f_ASAP7_75t_L g1209 ( 
.A(n_1020),
.Y(n_1209)
);

INVx3_ASAP7_75t_L g1210 ( 
.A(n_1091),
.Y(n_1210)
);

AND2x2_ASAP7_75t_L g1211 ( 
.A(n_938),
.B(n_481),
.Y(n_1211)
);

BUFx3_ASAP7_75t_L g1212 ( 
.A(n_937),
.Y(n_1212)
);

BUFx8_ASAP7_75t_SL g1213 ( 
.A(n_838),
.Y(n_1213)
);

BUFx3_ASAP7_75t_L g1214 ( 
.A(n_939),
.Y(n_1214)
);

NOR2xp33_ASAP7_75t_L g1215 ( 
.A(n_829),
.B(n_481),
.Y(n_1215)
);

BUFx8_ASAP7_75t_SL g1216 ( 
.A(n_857),
.Y(n_1216)
);

BUFx3_ASAP7_75t_L g1217 ( 
.A(n_940),
.Y(n_1217)
);

BUFx6f_ASAP7_75t_L g1218 ( 
.A(n_1091),
.Y(n_1218)
);

OAI22x1_ASAP7_75t_R g1219 ( 
.A1(n_922),
.A2(n_536),
.B1(n_641),
.B2(n_534),
.Y(n_1219)
);

INVx1_ASAP7_75t_L g1220 ( 
.A(n_960),
.Y(n_1220)
);

INVx1_ASAP7_75t_L g1221 ( 
.A(n_961),
.Y(n_1221)
);

INVx2_ASAP7_75t_L g1222 ( 
.A(n_868),
.Y(n_1222)
);

AND2x2_ASAP7_75t_L g1223 ( 
.A(n_1097),
.B(n_483),
.Y(n_1223)
);

INVx3_ASAP7_75t_L g1224 ( 
.A(n_868),
.Y(n_1224)
);

NAND2xp5_ASAP7_75t_L g1225 ( 
.A(n_1056),
.B(n_635),
.Y(n_1225)
);

BUFx6f_ASAP7_75t_L g1226 ( 
.A(n_878),
.Y(n_1226)
);

INVx2_ASAP7_75t_L g1227 ( 
.A(n_878),
.Y(n_1227)
);

NAND2xp5_ASAP7_75t_L g1228 ( 
.A(n_1058),
.B(n_636),
.Y(n_1228)
);

BUFx12f_ASAP7_75t_L g1229 ( 
.A(n_1064),
.Y(n_1229)
);

BUFx6f_ASAP7_75t_L g1230 ( 
.A(n_890),
.Y(n_1230)
);

BUFx6f_ASAP7_75t_L g1231 ( 
.A(n_890),
.Y(n_1231)
);

CKINVDCx5p33_ASAP7_75t_R g1232 ( 
.A(n_1087),
.Y(n_1232)
);

NAND2xp5_ASAP7_75t_L g1233 ( 
.A(n_1095),
.B(n_665),
.Y(n_1233)
);

INVx1_ASAP7_75t_L g1234 ( 
.A(n_964),
.Y(n_1234)
);

INVx3_ASAP7_75t_L g1235 ( 
.A(n_916),
.Y(n_1235)
);

INVx2_ASAP7_75t_SL g1236 ( 
.A(n_953),
.Y(n_1236)
);

NOR2xp33_ASAP7_75t_L g1237 ( 
.A(n_829),
.B(n_483),
.Y(n_1237)
);

INVx1_ASAP7_75t_L g1238 ( 
.A(n_966),
.Y(n_1238)
);

BUFx6f_ASAP7_75t_L g1239 ( 
.A(n_924),
.Y(n_1239)
);

INVx2_ASAP7_75t_L g1240 ( 
.A(n_924),
.Y(n_1240)
);

INVx2_ASAP7_75t_L g1241 ( 
.A(n_934),
.Y(n_1241)
);

BUFx3_ASAP7_75t_L g1242 ( 
.A(n_827),
.Y(n_1242)
);

INVx1_ASAP7_75t_L g1243 ( 
.A(n_971),
.Y(n_1243)
);

AOI22xp5_ASAP7_75t_L g1244 ( 
.A1(n_866),
.A2(n_474),
.B1(n_476),
.B2(n_471),
.Y(n_1244)
);

INVx3_ASAP7_75t_L g1245 ( 
.A(n_934),
.Y(n_1245)
);

BUFx12f_ASAP7_75t_L g1246 ( 
.A(n_1108),
.Y(n_1246)
);

BUFx2_ASAP7_75t_L g1247 ( 
.A(n_1078),
.Y(n_1247)
);

INVx6_ASAP7_75t_L g1248 ( 
.A(n_1102),
.Y(n_1248)
);

INVx2_ASAP7_75t_L g1249 ( 
.A(n_942),
.Y(n_1249)
);

INVx1_ASAP7_75t_L g1250 ( 
.A(n_975),
.Y(n_1250)
);

INVx2_ASAP7_75t_L g1251 ( 
.A(n_942),
.Y(n_1251)
);

BUFx6f_ASAP7_75t_L g1252 ( 
.A(n_950),
.Y(n_1252)
);

INVx2_ASAP7_75t_L g1253 ( 
.A(n_950),
.Y(n_1253)
);

INVx5_ASAP7_75t_L g1254 ( 
.A(n_972),
.Y(n_1254)
);

AND2x2_ASAP7_75t_L g1255 ( 
.A(n_931),
.B(n_944),
.Y(n_1255)
);

BUFx3_ASAP7_75t_L g1256 ( 
.A(n_828),
.Y(n_1256)
);

INVx2_ASAP7_75t_L g1257 ( 
.A(n_972),
.Y(n_1257)
);

CKINVDCx20_ASAP7_75t_R g1258 ( 
.A(n_970),
.Y(n_1258)
);

BUFx6f_ASAP7_75t_L g1259 ( 
.A(n_981),
.Y(n_1259)
);

INVx2_ASAP7_75t_SL g1260 ( 
.A(n_1016),
.Y(n_1260)
);

BUFx6f_ASAP7_75t_L g1261 ( 
.A(n_981),
.Y(n_1261)
);

AO22x1_ASAP7_75t_L g1262 ( 
.A1(n_1111),
.A2(n_536),
.B1(n_641),
.B2(n_534),
.Y(n_1262)
);

BUFx3_ASAP7_75t_L g1263 ( 
.A(n_832),
.Y(n_1263)
);

NOR2xp33_ASAP7_75t_L g1264 ( 
.A(n_867),
.B(n_1071),
.Y(n_1264)
);

INVx1_ASAP7_75t_L g1265 ( 
.A(n_977),
.Y(n_1265)
);

INVx2_ASAP7_75t_L g1266 ( 
.A(n_1033),
.Y(n_1266)
);

INVx1_ASAP7_75t_L g1267 ( 
.A(n_978),
.Y(n_1267)
);

BUFx6f_ASAP7_75t_L g1268 ( 
.A(n_1033),
.Y(n_1268)
);

BUFx3_ASAP7_75t_L g1269 ( 
.A(n_833),
.Y(n_1269)
);

BUFx2_ASAP7_75t_L g1270 ( 
.A(n_1078),
.Y(n_1270)
);

INVx2_ASAP7_75t_L g1271 ( 
.A(n_1039),
.Y(n_1271)
);

INVx2_ASAP7_75t_L g1272 ( 
.A(n_1039),
.Y(n_1272)
);

AND2x4_ASAP7_75t_L g1273 ( 
.A(n_1018),
.B(n_825),
.Y(n_1273)
);

INVx2_ASAP7_75t_L g1274 ( 
.A(n_1043),
.Y(n_1274)
);

INVx5_ASAP7_75t_L g1275 ( 
.A(n_1043),
.Y(n_1275)
);

INVx2_ASAP7_75t_L g1276 ( 
.A(n_1045),
.Y(n_1276)
);

INVx6_ASAP7_75t_L g1277 ( 
.A(n_1102),
.Y(n_1277)
);

INVx3_ASAP7_75t_L g1278 ( 
.A(n_1045),
.Y(n_1278)
);

BUFx2_ASAP7_75t_L g1279 ( 
.A(n_1016),
.Y(n_1279)
);

NOR2xp33_ASAP7_75t_L g1280 ( 
.A(n_867),
.B(n_494),
.Y(n_1280)
);

BUFx6f_ASAP7_75t_L g1281 ( 
.A(n_854),
.Y(n_1281)
);

AND2x4_ASAP7_75t_L g1282 ( 
.A(n_1029),
.B(n_494),
.Y(n_1282)
);

INVx1_ASAP7_75t_L g1283 ( 
.A(n_979),
.Y(n_1283)
);

BUFx8_ASAP7_75t_L g1284 ( 
.A(n_1083),
.Y(n_1284)
);

INVx5_ASAP7_75t_L g1285 ( 
.A(n_1061),
.Y(n_1285)
);

HB1xp67_ASAP7_75t_L g1286 ( 
.A(n_973),
.Y(n_1286)
);

AND2x2_ASAP7_75t_L g1287 ( 
.A(n_938),
.B(n_496),
.Y(n_1287)
);

AOI22xp5_ASAP7_75t_L g1288 ( 
.A1(n_866),
.A2(n_547),
.B1(n_579),
.B2(n_542),
.Y(n_1288)
);

INVx2_ASAP7_75t_L g1289 ( 
.A(n_1051),
.Y(n_1289)
);

NAND2xp5_ASAP7_75t_L g1290 ( 
.A(n_1138),
.B(n_1102),
.Y(n_1290)
);

NAND2xp5_ASAP7_75t_L g1291 ( 
.A(n_1138),
.B(n_1102),
.Y(n_1291)
);

BUFx6f_ASAP7_75t_L g1292 ( 
.A(n_1116),
.Y(n_1292)
);

INVx2_ASAP7_75t_L g1293 ( 
.A(n_1124),
.Y(n_1293)
);

NAND2xp5_ASAP7_75t_L g1294 ( 
.A(n_1144),
.B(n_1264),
.Y(n_1294)
);

NAND2xp5_ASAP7_75t_L g1295 ( 
.A(n_1144),
.B(n_1102),
.Y(n_1295)
);

BUFx6f_ASAP7_75t_L g1296 ( 
.A(n_1116),
.Y(n_1296)
);

INVx2_ASAP7_75t_L g1297 ( 
.A(n_1124),
.Y(n_1297)
);

AND2x2_ASAP7_75t_L g1298 ( 
.A(n_1255),
.B(n_1180),
.Y(n_1298)
);

AND2x4_ASAP7_75t_L g1299 ( 
.A(n_1140),
.B(n_835),
.Y(n_1299)
);

INVx1_ASAP7_75t_L g1300 ( 
.A(n_1155),
.Y(n_1300)
);

BUFx6f_ASAP7_75t_L g1301 ( 
.A(n_1116),
.Y(n_1301)
);

NAND2xp33_ASAP7_75t_L g1302 ( 
.A(n_1163),
.B(n_841),
.Y(n_1302)
);

INVxp67_ASAP7_75t_L g1303 ( 
.A(n_1255),
.Y(n_1303)
);

INVx1_ASAP7_75t_L g1304 ( 
.A(n_1161),
.Y(n_1304)
);

INVx1_ASAP7_75t_L g1305 ( 
.A(n_1168),
.Y(n_1305)
);

NAND2xp5_ASAP7_75t_SL g1306 ( 
.A(n_1117),
.B(n_951),
.Y(n_1306)
);

BUFx2_ASAP7_75t_L g1307 ( 
.A(n_1186),
.Y(n_1307)
);

AND2x2_ASAP7_75t_L g1308 ( 
.A(n_1180),
.B(n_1011),
.Y(n_1308)
);

INVx1_ASAP7_75t_L g1309 ( 
.A(n_1174),
.Y(n_1309)
);

INVx1_ASAP7_75t_L g1310 ( 
.A(n_1176),
.Y(n_1310)
);

NAND2xp5_ASAP7_75t_L g1311 ( 
.A(n_1264),
.B(n_1011),
.Y(n_1311)
);

AND2x4_ASAP7_75t_L g1312 ( 
.A(n_1140),
.B(n_837),
.Y(n_1312)
);

NAND2xp5_ASAP7_75t_L g1313 ( 
.A(n_1117),
.B(n_1050),
.Y(n_1313)
);

INVx1_ASAP7_75t_L g1314 ( 
.A(n_1179),
.Y(n_1314)
);

AND2x2_ASAP7_75t_L g1315 ( 
.A(n_1196),
.B(n_1050),
.Y(n_1315)
);

INVx2_ASAP7_75t_L g1316 ( 
.A(n_1125),
.Y(n_1316)
);

INVx1_ASAP7_75t_L g1317 ( 
.A(n_1202),
.Y(n_1317)
);

INVx1_ASAP7_75t_L g1318 ( 
.A(n_1204),
.Y(n_1318)
);

AND2x4_ASAP7_75t_L g1319 ( 
.A(n_1142),
.B(n_839),
.Y(n_1319)
);

NAND2xp5_ASAP7_75t_L g1320 ( 
.A(n_1117),
.B(n_1082),
.Y(n_1320)
);

INVx3_ASAP7_75t_L g1321 ( 
.A(n_1127),
.Y(n_1321)
);

INVx3_ASAP7_75t_L g1322 ( 
.A(n_1127),
.Y(n_1322)
);

AND2x2_ASAP7_75t_L g1323 ( 
.A(n_1196),
.B(n_1111),
.Y(n_1323)
);

INVx2_ASAP7_75t_L g1324 ( 
.A(n_1125),
.Y(n_1324)
);

INVx1_ASAP7_75t_L g1325 ( 
.A(n_1208),
.Y(n_1325)
);

INVx2_ASAP7_75t_L g1326 ( 
.A(n_1128),
.Y(n_1326)
);

INVx1_ASAP7_75t_L g1327 ( 
.A(n_1220),
.Y(n_1327)
);

INVx1_ASAP7_75t_L g1328 ( 
.A(n_1221),
.Y(n_1328)
);

INVx1_ASAP7_75t_L g1329 ( 
.A(n_1234),
.Y(n_1329)
);

NAND2x1p5_ASAP7_75t_L g1330 ( 
.A(n_1285),
.B(n_1100),
.Y(n_1330)
);

INVx1_ASAP7_75t_L g1331 ( 
.A(n_1238),
.Y(n_1331)
);

AND2x4_ASAP7_75t_L g1332 ( 
.A(n_1142),
.B(n_844),
.Y(n_1332)
);

INVx1_ASAP7_75t_L g1333 ( 
.A(n_1243),
.Y(n_1333)
);

CKINVDCx5p33_ASAP7_75t_R g1334 ( 
.A(n_1216),
.Y(n_1334)
);

INVx2_ASAP7_75t_L g1335 ( 
.A(n_1128),
.Y(n_1335)
);

INVx1_ASAP7_75t_L g1336 ( 
.A(n_1250),
.Y(n_1336)
);

HB1xp67_ASAP7_75t_L g1337 ( 
.A(n_1207),
.Y(n_1337)
);

BUFx2_ASAP7_75t_L g1338 ( 
.A(n_1286),
.Y(n_1338)
);

BUFx6f_ASAP7_75t_L g1339 ( 
.A(n_1149),
.Y(n_1339)
);

BUFx8_ASAP7_75t_L g1340 ( 
.A(n_1121),
.Y(n_1340)
);

INVx2_ASAP7_75t_L g1341 ( 
.A(n_1135),
.Y(n_1341)
);

AND2x2_ASAP7_75t_L g1342 ( 
.A(n_1201),
.B(n_976),
.Y(n_1342)
);

NAND2xp5_ASAP7_75t_L g1343 ( 
.A(n_1131),
.B(n_1082),
.Y(n_1343)
);

INVx1_ASAP7_75t_L g1344 ( 
.A(n_1265),
.Y(n_1344)
);

INVx1_ASAP7_75t_L g1345 ( 
.A(n_1267),
.Y(n_1345)
);

AND2x2_ASAP7_75t_L g1346 ( 
.A(n_1201),
.B(n_1103),
.Y(n_1346)
);

CKINVDCx5p33_ASAP7_75t_R g1347 ( 
.A(n_1216),
.Y(n_1347)
);

INVx1_ASAP7_75t_L g1348 ( 
.A(n_1283),
.Y(n_1348)
);

BUFx6f_ASAP7_75t_L g1349 ( 
.A(n_1149),
.Y(n_1349)
);

INVx1_ASAP7_75t_L g1350 ( 
.A(n_1242),
.Y(n_1350)
);

INVx2_ASAP7_75t_L g1351 ( 
.A(n_1135),
.Y(n_1351)
);

INVx1_ASAP7_75t_L g1352 ( 
.A(n_1242),
.Y(n_1352)
);

NAND2xp5_ASAP7_75t_L g1353 ( 
.A(n_1131),
.B(n_980),
.Y(n_1353)
);

AND2x2_ASAP7_75t_L g1354 ( 
.A(n_1223),
.B(n_1107),
.Y(n_1354)
);

AND2x2_ASAP7_75t_L g1355 ( 
.A(n_1223),
.B(n_1105),
.Y(n_1355)
);

BUFx6f_ASAP7_75t_L g1356 ( 
.A(n_1149),
.Y(n_1356)
);

INVx2_ASAP7_75t_L g1357 ( 
.A(n_1145),
.Y(n_1357)
);

INVx1_ASAP7_75t_L g1358 ( 
.A(n_1256),
.Y(n_1358)
);

INVx1_ASAP7_75t_L g1359 ( 
.A(n_1256),
.Y(n_1359)
);

INVx1_ASAP7_75t_L g1360 ( 
.A(n_1263),
.Y(n_1360)
);

INVx1_ASAP7_75t_L g1361 ( 
.A(n_1263),
.Y(n_1361)
);

OAI21x1_ASAP7_75t_L g1362 ( 
.A1(n_1115),
.A2(n_1053),
.B(n_1052),
.Y(n_1362)
);

INVx2_ASAP7_75t_L g1363 ( 
.A(n_1145),
.Y(n_1363)
);

BUFx3_ASAP7_75t_L g1364 ( 
.A(n_1148),
.Y(n_1364)
);

NOR2xp33_ASAP7_75t_L g1365 ( 
.A(n_1215),
.B(n_849),
.Y(n_1365)
);

AND2x4_ASAP7_75t_L g1366 ( 
.A(n_1126),
.B(n_847),
.Y(n_1366)
);

INVx1_ASAP7_75t_L g1367 ( 
.A(n_1269),
.Y(n_1367)
);

CKINVDCx8_ASAP7_75t_R g1368 ( 
.A(n_1137),
.Y(n_1368)
);

INVx2_ASAP7_75t_L g1369 ( 
.A(n_1151),
.Y(n_1369)
);

INVx1_ASAP7_75t_SL g1370 ( 
.A(n_1258),
.Y(n_1370)
);

INVx3_ASAP7_75t_L g1371 ( 
.A(n_1149),
.Y(n_1371)
);

NOR2xp33_ASAP7_75t_L g1372 ( 
.A(n_1215),
.B(n_983),
.Y(n_1372)
);

INVx1_ASAP7_75t_L g1373 ( 
.A(n_1269),
.Y(n_1373)
);

AND2x4_ASAP7_75t_L g1374 ( 
.A(n_1148),
.B(n_1158),
.Y(n_1374)
);

CKINVDCx5p33_ASAP7_75t_R g1375 ( 
.A(n_1153),
.Y(n_1375)
);

AND2x2_ASAP7_75t_SL g1376 ( 
.A(n_1166),
.B(n_963),
.Y(n_1376)
);

NAND2xp5_ASAP7_75t_L g1377 ( 
.A(n_1131),
.B(n_982),
.Y(n_1377)
);

AND2x4_ASAP7_75t_L g1378 ( 
.A(n_1158),
.B(n_1077),
.Y(n_1378)
);

NAND2xp5_ASAP7_75t_L g1379 ( 
.A(n_1237),
.B(n_984),
.Y(n_1379)
);

NAND2xp5_ASAP7_75t_L g1380 ( 
.A(n_1237),
.B(n_985),
.Y(n_1380)
);

NAND2xp5_ASAP7_75t_L g1381 ( 
.A(n_1280),
.B(n_986),
.Y(n_1381)
);

INVx2_ASAP7_75t_L g1382 ( 
.A(n_1151),
.Y(n_1382)
);

OA21x2_ASAP7_75t_L g1383 ( 
.A1(n_1152),
.A2(n_1055),
.B(n_1054),
.Y(n_1383)
);

AND2x2_ASAP7_75t_L g1384 ( 
.A(n_1150),
.B(n_1109),
.Y(n_1384)
);

AND2x4_ASAP7_75t_L g1385 ( 
.A(n_1170),
.B(n_1079),
.Y(n_1385)
);

AND2x2_ASAP7_75t_L g1386 ( 
.A(n_1150),
.B(n_1110),
.Y(n_1386)
);

OAI22xp5_ASAP7_75t_L g1387 ( 
.A1(n_1280),
.A2(n_891),
.B1(n_906),
.B2(n_892),
.Y(n_1387)
);

INVx1_ASAP7_75t_L g1388 ( 
.A(n_1170),
.Y(n_1388)
);

INVx2_ASAP7_75t_L g1389 ( 
.A(n_1152),
.Y(n_1389)
);

INVx2_ASAP7_75t_L g1390 ( 
.A(n_1154),
.Y(n_1390)
);

INVx2_ASAP7_75t_L g1391 ( 
.A(n_1154),
.Y(n_1391)
);

INVxp67_ASAP7_75t_L g1392 ( 
.A(n_1123),
.Y(n_1392)
);

INVx1_ASAP7_75t_L g1393 ( 
.A(n_1187),
.Y(n_1393)
);

INVx1_ASAP7_75t_L g1394 ( 
.A(n_1187),
.Y(n_1394)
);

INVx1_ASAP7_75t_L g1395 ( 
.A(n_1194),
.Y(n_1395)
);

NOR2xp33_ASAP7_75t_SL g1396 ( 
.A(n_1136),
.B(n_1185),
.Y(n_1396)
);

AND2x2_ASAP7_75t_L g1397 ( 
.A(n_1279),
.B(n_1112),
.Y(n_1397)
);

INVx2_ASAP7_75t_L g1398 ( 
.A(n_1226),
.Y(n_1398)
);

INVx2_ASAP7_75t_L g1399 ( 
.A(n_1226),
.Y(n_1399)
);

HB1xp67_ASAP7_75t_L g1400 ( 
.A(n_1147),
.Y(n_1400)
);

AND2x2_ASAP7_75t_L g1401 ( 
.A(n_1126),
.B(n_1113),
.Y(n_1401)
);

NOR2xp33_ASAP7_75t_L g1402 ( 
.A(n_1156),
.B(n_891),
.Y(n_1402)
);

INVx1_ASAP7_75t_L g1403 ( 
.A(n_1194),
.Y(n_1403)
);

INVx1_ASAP7_75t_L g1404 ( 
.A(n_1212),
.Y(n_1404)
);

INVx3_ASAP7_75t_L g1405 ( 
.A(n_1167),
.Y(n_1405)
);

NAND2xp5_ASAP7_75t_L g1406 ( 
.A(n_1134),
.B(n_1198),
.Y(n_1406)
);

INVx2_ASAP7_75t_L g1407 ( 
.A(n_1226),
.Y(n_1407)
);

INVx1_ASAP7_75t_L g1408 ( 
.A(n_1212),
.Y(n_1408)
);

INVx1_ASAP7_75t_L g1409 ( 
.A(n_1214),
.Y(n_1409)
);

INVx1_ASAP7_75t_L g1410 ( 
.A(n_1214),
.Y(n_1410)
);

INVx1_ASAP7_75t_L g1411 ( 
.A(n_1217),
.Y(n_1411)
);

INVx2_ASAP7_75t_L g1412 ( 
.A(n_1226),
.Y(n_1412)
);

NAND2xp5_ASAP7_75t_L g1413 ( 
.A(n_1225),
.B(n_989),
.Y(n_1413)
);

BUFx6f_ASAP7_75t_L g1414 ( 
.A(n_1167),
.Y(n_1414)
);

AND2x2_ASAP7_75t_L g1415 ( 
.A(n_1236),
.B(n_1008),
.Y(n_1415)
);

AND2x4_ASAP7_75t_L g1416 ( 
.A(n_1236),
.B(n_850),
.Y(n_1416)
);

AND2x4_ASAP7_75t_L g1417 ( 
.A(n_1260),
.B(n_1101),
.Y(n_1417)
);

OAI21x1_ASAP7_75t_L g1418 ( 
.A1(n_1228),
.A2(n_1060),
.B(n_1057),
.Y(n_1418)
);

OA21x2_ASAP7_75t_L g1419 ( 
.A1(n_1118),
.A2(n_1063),
.B(n_1062),
.Y(n_1419)
);

INVx1_ASAP7_75t_L g1420 ( 
.A(n_1217),
.Y(n_1420)
);

INVx2_ASAP7_75t_L g1421 ( 
.A(n_1230),
.Y(n_1421)
);

AND2x2_ASAP7_75t_L g1422 ( 
.A(n_1260),
.B(n_1076),
.Y(n_1422)
);

AND2x4_ASAP7_75t_L g1423 ( 
.A(n_1285),
.B(n_1104),
.Y(n_1423)
);

BUFx2_ASAP7_75t_L g1424 ( 
.A(n_1258),
.Y(n_1424)
);

INVx1_ASAP7_75t_L g1425 ( 
.A(n_1281),
.Y(n_1425)
);

CKINVDCx5p33_ASAP7_75t_R g1426 ( 
.A(n_1153),
.Y(n_1426)
);

INVx2_ASAP7_75t_L g1427 ( 
.A(n_1230),
.Y(n_1427)
);

AND2x2_ASAP7_75t_L g1428 ( 
.A(n_1205),
.B(n_1061),
.Y(n_1428)
);

INVx1_ASAP7_75t_L g1429 ( 
.A(n_1281),
.Y(n_1429)
);

NAND2xp5_ASAP7_75t_L g1430 ( 
.A(n_1233),
.B(n_991),
.Y(n_1430)
);

NAND2xp5_ASAP7_75t_SL g1431 ( 
.A(n_1156),
.B(n_667),
.Y(n_1431)
);

INVx1_ASAP7_75t_L g1432 ( 
.A(n_1281),
.Y(n_1432)
);

NOR2xp33_ASAP7_75t_L g1433 ( 
.A(n_1156),
.B(n_892),
.Y(n_1433)
);

INVx1_ASAP7_75t_L g1434 ( 
.A(n_1281),
.Y(n_1434)
);

INVx2_ASAP7_75t_L g1435 ( 
.A(n_1230),
.Y(n_1435)
);

BUFx6f_ASAP7_75t_L g1436 ( 
.A(n_1172),
.Y(n_1436)
);

BUFx6f_ASAP7_75t_L g1437 ( 
.A(n_1172),
.Y(n_1437)
);

INVx1_ASAP7_75t_L g1438 ( 
.A(n_1231),
.Y(n_1438)
);

INVx2_ASAP7_75t_L g1439 ( 
.A(n_1231),
.Y(n_1439)
);

BUFx6f_ASAP7_75t_L g1440 ( 
.A(n_1172),
.Y(n_1440)
);

INVx1_ASAP7_75t_L g1441 ( 
.A(n_1231),
.Y(n_1441)
);

INVx1_ASAP7_75t_L g1442 ( 
.A(n_1231),
.Y(n_1442)
);

HB1xp67_ASAP7_75t_L g1443 ( 
.A(n_1273),
.Y(n_1443)
);

OAI22xp33_ASAP7_75t_L g1444 ( 
.A1(n_1294),
.A2(n_1288),
.B1(n_1244),
.B2(n_944),
.Y(n_1444)
);

OAI22xp33_ASAP7_75t_L g1445 ( 
.A1(n_1379),
.A2(n_931),
.B1(n_893),
.B2(n_842),
.Y(n_1445)
);

CKINVDCx20_ASAP7_75t_R g1446 ( 
.A(n_1368),
.Y(n_1446)
);

NOR2xp33_ASAP7_75t_L g1447 ( 
.A(n_1303),
.B(n_1114),
.Y(n_1447)
);

NAND2xp5_ASAP7_75t_L g1448 ( 
.A(n_1290),
.B(n_1273),
.Y(n_1448)
);

CKINVDCx16_ASAP7_75t_R g1449 ( 
.A(n_1337),
.Y(n_1449)
);

INVx1_ASAP7_75t_L g1450 ( 
.A(n_1300),
.Y(n_1450)
);

INVx4_ASAP7_75t_L g1451 ( 
.A(n_1374),
.Y(n_1451)
);

AOI22xp5_ASAP7_75t_L g1452 ( 
.A1(n_1365),
.A2(n_1273),
.B1(n_1282),
.B2(n_1166),
.Y(n_1452)
);

AOI21x1_ASAP7_75t_L g1453 ( 
.A1(n_1295),
.A2(n_1291),
.B(n_1406),
.Y(n_1453)
);

CKINVDCx20_ASAP7_75t_R g1454 ( 
.A(n_1375),
.Y(n_1454)
);

INVx2_ASAP7_75t_L g1455 ( 
.A(n_1293),
.Y(n_1455)
);

AOI22xp33_ASAP7_75t_SL g1456 ( 
.A1(n_1365),
.A2(n_1005),
.B1(n_1010),
.B2(n_987),
.Y(n_1456)
);

INVx2_ASAP7_75t_L g1457 ( 
.A(n_1293),
.Y(n_1457)
);

NAND2xp5_ASAP7_75t_L g1458 ( 
.A(n_1413),
.B(n_1282),
.Y(n_1458)
);

INVx1_ASAP7_75t_L g1459 ( 
.A(n_1304),
.Y(n_1459)
);

BUFx6f_ASAP7_75t_L g1460 ( 
.A(n_1383),
.Y(n_1460)
);

BUFx6f_ASAP7_75t_L g1461 ( 
.A(n_1383),
.Y(n_1461)
);

NAND2xp5_ASAP7_75t_L g1462 ( 
.A(n_1430),
.B(n_1282),
.Y(n_1462)
);

INVx2_ASAP7_75t_L g1463 ( 
.A(n_1297),
.Y(n_1463)
);

INVx1_ASAP7_75t_L g1464 ( 
.A(n_1305),
.Y(n_1464)
);

AOI22xp5_ASAP7_75t_L g1465 ( 
.A1(n_1372),
.A2(n_1166),
.B1(n_1188),
.B2(n_1133),
.Y(n_1465)
);

CKINVDCx5p33_ASAP7_75t_R g1466 ( 
.A(n_1375),
.Y(n_1466)
);

AND2x6_ASAP7_75t_L g1467 ( 
.A(n_1315),
.B(n_1157),
.Y(n_1467)
);

CKINVDCx5p33_ASAP7_75t_R g1468 ( 
.A(n_1426),
.Y(n_1468)
);

INVx2_ASAP7_75t_L g1469 ( 
.A(n_1297),
.Y(n_1469)
);

INVx1_ASAP7_75t_L g1470 ( 
.A(n_1309),
.Y(n_1470)
);

NAND3xp33_ASAP7_75t_L g1471 ( 
.A(n_1372),
.B(n_1175),
.C(n_1171),
.Y(n_1471)
);

INVx3_ASAP7_75t_L g1472 ( 
.A(n_1383),
.Y(n_1472)
);

CKINVDCx20_ASAP7_75t_R g1473 ( 
.A(n_1424),
.Y(n_1473)
);

INVx1_ASAP7_75t_L g1474 ( 
.A(n_1310),
.Y(n_1474)
);

NAND2xp5_ASAP7_75t_SL g1475 ( 
.A(n_1376),
.B(n_1171),
.Y(n_1475)
);

AOI22xp33_ASAP7_75t_L g1476 ( 
.A1(n_1376),
.A2(n_1188),
.B1(n_1163),
.B2(n_1132),
.Y(n_1476)
);

NAND2xp5_ASAP7_75t_SL g1477 ( 
.A(n_1443),
.B(n_1175),
.Y(n_1477)
);

NAND2xp5_ASAP7_75t_L g1478 ( 
.A(n_1380),
.B(n_1248),
.Y(n_1478)
);

INVx2_ASAP7_75t_L g1479 ( 
.A(n_1316),
.Y(n_1479)
);

AND2x2_ASAP7_75t_L g1480 ( 
.A(n_1323),
.B(n_1211),
.Y(n_1480)
);

NAND2xp5_ASAP7_75t_L g1481 ( 
.A(n_1381),
.B(n_1248),
.Y(n_1481)
);

INVx2_ASAP7_75t_L g1482 ( 
.A(n_1316),
.Y(n_1482)
);

INVx2_ASAP7_75t_L g1483 ( 
.A(n_1324),
.Y(n_1483)
);

INVx1_ASAP7_75t_L g1484 ( 
.A(n_1314),
.Y(n_1484)
);

INVx2_ASAP7_75t_L g1485 ( 
.A(n_1324),
.Y(n_1485)
);

INVx1_ASAP7_75t_L g1486 ( 
.A(n_1317),
.Y(n_1486)
);

BUFx3_ASAP7_75t_L g1487 ( 
.A(n_1364),
.Y(n_1487)
);

OAI22xp33_ASAP7_75t_SL g1488 ( 
.A1(n_1306),
.A2(n_1443),
.B1(n_1303),
.B2(n_1431),
.Y(n_1488)
);

NAND2xp33_ASAP7_75t_L g1489 ( 
.A(n_1311),
.B(n_1313),
.Y(n_1489)
);

BUFx3_ASAP7_75t_L g1490 ( 
.A(n_1364),
.Y(n_1490)
);

BUFx2_ASAP7_75t_L g1491 ( 
.A(n_1307),
.Y(n_1491)
);

NAND2xp5_ASAP7_75t_L g1492 ( 
.A(n_1306),
.B(n_1248),
.Y(n_1492)
);

INVx1_ASAP7_75t_L g1493 ( 
.A(n_1318),
.Y(n_1493)
);

INVx1_ASAP7_75t_L g1494 ( 
.A(n_1325),
.Y(n_1494)
);

BUFx6f_ASAP7_75t_L g1495 ( 
.A(n_1292),
.Y(n_1495)
);

INVx1_ASAP7_75t_L g1496 ( 
.A(n_1327),
.Y(n_1496)
);

INVx1_ASAP7_75t_L g1497 ( 
.A(n_1328),
.Y(n_1497)
);

INVx1_ASAP7_75t_L g1498 ( 
.A(n_1329),
.Y(n_1498)
);

INVx2_ASAP7_75t_L g1499 ( 
.A(n_1326),
.Y(n_1499)
);

INVx1_ASAP7_75t_L g1500 ( 
.A(n_1331),
.Y(n_1500)
);

NAND2xp5_ASAP7_75t_L g1501 ( 
.A(n_1320),
.B(n_1277),
.Y(n_1501)
);

INVx1_ASAP7_75t_L g1502 ( 
.A(n_1333),
.Y(n_1502)
);

INVx2_ASAP7_75t_SL g1503 ( 
.A(n_1337),
.Y(n_1503)
);

NOR2xp33_ASAP7_75t_L g1504 ( 
.A(n_1354),
.B(n_1232),
.Y(n_1504)
);

AOI22xp5_ASAP7_75t_L g1505 ( 
.A1(n_1402),
.A2(n_1188),
.B1(n_1232),
.B2(n_1163),
.Y(n_1505)
);

INVx2_ASAP7_75t_L g1506 ( 
.A(n_1326),
.Y(n_1506)
);

INVx1_ASAP7_75t_L g1507 ( 
.A(n_1336),
.Y(n_1507)
);

NAND2xp5_ASAP7_75t_SL g1508 ( 
.A(n_1402),
.B(n_1285),
.Y(n_1508)
);

NOR2x1p5_ASAP7_75t_L g1509 ( 
.A(n_1308),
.B(n_1169),
.Y(n_1509)
);

INVx4_ASAP7_75t_L g1510 ( 
.A(n_1374),
.Y(n_1510)
);

INVx2_ASAP7_75t_L g1511 ( 
.A(n_1335),
.Y(n_1511)
);

NAND2xp5_ASAP7_75t_L g1512 ( 
.A(n_1343),
.B(n_1277),
.Y(n_1512)
);

BUFx3_ASAP7_75t_L g1513 ( 
.A(n_1299),
.Y(n_1513)
);

INVx1_ASAP7_75t_L g1514 ( 
.A(n_1344),
.Y(n_1514)
);

OAI22xp33_ASAP7_75t_L g1515 ( 
.A1(n_1353),
.A2(n_821),
.B1(n_620),
.B2(n_1085),
.Y(n_1515)
);

INVx2_ASAP7_75t_L g1516 ( 
.A(n_1335),
.Y(n_1516)
);

AND2x2_ASAP7_75t_L g1517 ( 
.A(n_1415),
.B(n_1287),
.Y(n_1517)
);

INVx3_ASAP7_75t_L g1518 ( 
.A(n_1419),
.Y(n_1518)
);

NAND2xp33_ASAP7_75t_R g1519 ( 
.A(n_1338),
.B(n_1143),
.Y(n_1519)
);

INVx1_ASAP7_75t_L g1520 ( 
.A(n_1345),
.Y(n_1520)
);

AND2x2_ASAP7_75t_L g1521 ( 
.A(n_1422),
.B(n_1164),
.Y(n_1521)
);

AND2x2_ASAP7_75t_L g1522 ( 
.A(n_1346),
.B(n_1164),
.Y(n_1522)
);

NAND2xp5_ASAP7_75t_L g1523 ( 
.A(n_1355),
.B(n_1277),
.Y(n_1523)
);

AND2x2_ASAP7_75t_SL g1524 ( 
.A(n_1302),
.B(n_1433),
.Y(n_1524)
);

INVx1_ASAP7_75t_L g1525 ( 
.A(n_1348),
.Y(n_1525)
);

INVx1_ASAP7_75t_L g1526 ( 
.A(n_1378),
.Y(n_1526)
);

INVxp67_ASAP7_75t_SL g1527 ( 
.A(n_1419),
.Y(n_1527)
);

OAI22xp5_ASAP7_75t_L g1528 ( 
.A1(n_1433),
.A2(n_708),
.B1(n_745),
.B2(n_631),
.Y(n_1528)
);

INVx2_ASAP7_75t_L g1529 ( 
.A(n_1341),
.Y(n_1529)
);

INVx2_ASAP7_75t_L g1530 ( 
.A(n_1341),
.Y(n_1530)
);

INVx1_ASAP7_75t_L g1531 ( 
.A(n_1378),
.Y(n_1531)
);

BUFx8_ASAP7_75t_SL g1532 ( 
.A(n_1334),
.Y(n_1532)
);

INVx2_ASAP7_75t_L g1533 ( 
.A(n_1351),
.Y(n_1533)
);

NAND2xp5_ASAP7_75t_L g1534 ( 
.A(n_1384),
.B(n_1122),
.Y(n_1534)
);

BUFx2_ASAP7_75t_L g1535 ( 
.A(n_1400),
.Y(n_1535)
);

OAI22xp33_ASAP7_75t_L g1536 ( 
.A1(n_1377),
.A2(n_782),
.B1(n_785),
.B2(n_784),
.Y(n_1536)
);

NOR2xp33_ASAP7_75t_L g1537 ( 
.A(n_1387),
.B(n_906),
.Y(n_1537)
);

INVx1_ASAP7_75t_L g1538 ( 
.A(n_1378),
.Y(n_1538)
);

INVx1_ASAP7_75t_L g1539 ( 
.A(n_1385),
.Y(n_1539)
);

NOR2xp33_ASAP7_75t_R g1540 ( 
.A(n_1426),
.B(n_1119),
.Y(n_1540)
);

INVx1_ASAP7_75t_L g1541 ( 
.A(n_1385),
.Y(n_1541)
);

OR2x2_ASAP7_75t_L g1542 ( 
.A(n_1400),
.B(n_988),
.Y(n_1542)
);

NAND2xp5_ASAP7_75t_L g1543 ( 
.A(n_1386),
.B(n_1159),
.Y(n_1543)
);

AOI22xp33_ASAP7_75t_L g1544 ( 
.A1(n_1302),
.A2(n_1163),
.B1(n_1132),
.B2(n_1067),
.Y(n_1544)
);

OAI22xp33_ASAP7_75t_SL g1545 ( 
.A1(n_1431),
.A2(n_947),
.B1(n_996),
.B2(n_909),
.Y(n_1545)
);

INVx1_ASAP7_75t_L g1546 ( 
.A(n_1385),
.Y(n_1546)
);

NAND2xp33_ASAP7_75t_SL g1547 ( 
.A(n_1342),
.B(n_759),
.Y(n_1547)
);

NAND2xp33_ASAP7_75t_R g1548 ( 
.A(n_1397),
.B(n_1160),
.Y(n_1548)
);

BUFx3_ASAP7_75t_L g1549 ( 
.A(n_1299),
.Y(n_1549)
);

INVx1_ASAP7_75t_SL g1550 ( 
.A(n_1370),
.Y(n_1550)
);

INVx1_ASAP7_75t_L g1551 ( 
.A(n_1312),
.Y(n_1551)
);

NAND2xp33_ASAP7_75t_SL g1552 ( 
.A(n_1401),
.B(n_787),
.Y(n_1552)
);

BUFx10_ASAP7_75t_L g1553 ( 
.A(n_1334),
.Y(n_1553)
);

AOI22xp33_ASAP7_75t_L g1554 ( 
.A1(n_1419),
.A2(n_1163),
.B1(n_1068),
.B2(n_1069),
.Y(n_1554)
);

AND3x1_ASAP7_75t_L g1555 ( 
.A(n_1298),
.B(n_1035),
.C(n_1092),
.Y(n_1555)
);

NAND2xp5_ASAP7_75t_SL g1556 ( 
.A(n_1374),
.B(n_1285),
.Y(n_1556)
);

CKINVDCx5p33_ASAP7_75t_R g1557 ( 
.A(n_1347),
.Y(n_1557)
);

CKINVDCx5p33_ASAP7_75t_R g1558 ( 
.A(n_1347),
.Y(n_1558)
);

INVx2_ASAP7_75t_L g1559 ( 
.A(n_1351),
.Y(n_1559)
);

INVx3_ASAP7_75t_L g1560 ( 
.A(n_1321),
.Y(n_1560)
);

INVx2_ASAP7_75t_L g1561 ( 
.A(n_1357),
.Y(n_1561)
);

NAND2xp5_ASAP7_75t_SL g1562 ( 
.A(n_1366),
.B(n_1285),
.Y(n_1562)
);

INVx2_ASAP7_75t_L g1563 ( 
.A(n_1357),
.Y(n_1563)
);

NAND2xp5_ASAP7_75t_L g1564 ( 
.A(n_1425),
.B(n_1183),
.Y(n_1564)
);

NAND2xp5_ASAP7_75t_SL g1565 ( 
.A(n_1366),
.B(n_1136),
.Y(n_1565)
);

CKINVDCx6p67_ASAP7_75t_R g1566 ( 
.A(n_1312),
.Y(n_1566)
);

INVx1_ASAP7_75t_L g1567 ( 
.A(n_1319),
.Y(n_1567)
);

NAND2xp5_ASAP7_75t_L g1568 ( 
.A(n_1429),
.B(n_1239),
.Y(n_1568)
);

INVx1_ASAP7_75t_L g1569 ( 
.A(n_1319),
.Y(n_1569)
);

AND2x2_ASAP7_75t_L g1570 ( 
.A(n_1428),
.B(n_990),
.Y(n_1570)
);

INVx2_ASAP7_75t_L g1571 ( 
.A(n_1363),
.Y(n_1571)
);

NOR2xp33_ASAP7_75t_L g1572 ( 
.A(n_1416),
.B(n_909),
.Y(n_1572)
);

INVx2_ASAP7_75t_L g1573 ( 
.A(n_1363),
.Y(n_1573)
);

INVx1_ASAP7_75t_L g1574 ( 
.A(n_1332),
.Y(n_1574)
);

CKINVDCx5p33_ASAP7_75t_R g1575 ( 
.A(n_1340),
.Y(n_1575)
);

AND2x6_ASAP7_75t_L g1576 ( 
.A(n_1350),
.B(n_1093),
.Y(n_1576)
);

BUFx2_ASAP7_75t_L g1577 ( 
.A(n_1392),
.Y(n_1577)
);

BUFx2_ASAP7_75t_L g1578 ( 
.A(n_1392),
.Y(n_1578)
);

INVx2_ASAP7_75t_SL g1579 ( 
.A(n_1332),
.Y(n_1579)
);

INVx1_ASAP7_75t_L g1580 ( 
.A(n_1352),
.Y(n_1580)
);

INVx2_ASAP7_75t_L g1581 ( 
.A(n_1369),
.Y(n_1581)
);

BUFx6f_ASAP7_75t_L g1582 ( 
.A(n_1292),
.Y(n_1582)
);

NAND2xp5_ASAP7_75t_SL g1583 ( 
.A(n_1416),
.B(n_1185),
.Y(n_1583)
);

INVx1_ASAP7_75t_L g1584 ( 
.A(n_1358),
.Y(n_1584)
);

NAND2xp5_ASAP7_75t_L g1585 ( 
.A(n_1432),
.B(n_1239),
.Y(n_1585)
);

AOI22xp33_ASAP7_75t_L g1586 ( 
.A1(n_1369),
.A2(n_1073),
.B1(n_1074),
.B2(n_1065),
.Y(n_1586)
);

OAI22xp33_ASAP7_75t_SL g1587 ( 
.A1(n_1359),
.A2(n_996),
.B1(n_997),
.B2(n_947),
.Y(n_1587)
);

AND2x2_ASAP7_75t_L g1588 ( 
.A(n_1417),
.B(n_1017),
.Y(n_1588)
);

NAND2xp5_ASAP7_75t_L g1589 ( 
.A(n_1434),
.B(n_1239),
.Y(n_1589)
);

NOR2xp33_ASAP7_75t_L g1590 ( 
.A(n_1360),
.B(n_997),
.Y(n_1590)
);

INVx3_ASAP7_75t_L g1591 ( 
.A(n_1321),
.Y(n_1591)
);

NOR2xp33_ASAP7_75t_L g1592 ( 
.A(n_1361),
.B(n_1041),
.Y(n_1592)
);

INVx2_ASAP7_75t_L g1593 ( 
.A(n_1382),
.Y(n_1593)
);

INVx1_ASAP7_75t_L g1594 ( 
.A(n_1367),
.Y(n_1594)
);

NAND3xp33_ASAP7_75t_SL g1595 ( 
.A(n_1373),
.B(n_790),
.C(n_498),
.Y(n_1595)
);

HB1xp67_ASAP7_75t_L g1596 ( 
.A(n_1535),
.Y(n_1596)
);

INVx2_ASAP7_75t_L g1597 ( 
.A(n_1455),
.Y(n_1597)
);

BUFx6f_ASAP7_75t_L g1598 ( 
.A(n_1495),
.Y(n_1598)
);

BUFx6f_ASAP7_75t_L g1599 ( 
.A(n_1495),
.Y(n_1599)
);

INVx2_ASAP7_75t_L g1600 ( 
.A(n_1457),
.Y(n_1600)
);

INVx2_ASAP7_75t_SL g1601 ( 
.A(n_1503),
.Y(n_1601)
);

AO22x2_ASAP7_75t_L g1602 ( 
.A1(n_1475),
.A2(n_1165),
.B1(n_1139),
.B2(n_1162),
.Y(n_1602)
);

INVx3_ASAP7_75t_L g1603 ( 
.A(n_1451),
.Y(n_1603)
);

NAND2x1p5_ASAP7_75t_L g1604 ( 
.A(n_1451),
.B(n_1362),
.Y(n_1604)
);

BUFx3_ASAP7_75t_L g1605 ( 
.A(n_1491),
.Y(n_1605)
);

INVx1_ASAP7_75t_L g1606 ( 
.A(n_1450),
.Y(n_1606)
);

OR2x2_ASAP7_75t_L g1607 ( 
.A(n_1542),
.B(n_1177),
.Y(n_1607)
);

NAND2xp5_ASAP7_75t_SL g1608 ( 
.A(n_1447),
.B(n_1388),
.Y(n_1608)
);

INVx2_ASAP7_75t_SL g1609 ( 
.A(n_1588),
.Y(n_1609)
);

AND2x4_ASAP7_75t_L g1610 ( 
.A(n_1487),
.B(n_1393),
.Y(n_1610)
);

INVx1_ASAP7_75t_L g1611 ( 
.A(n_1459),
.Y(n_1611)
);

BUFx6f_ASAP7_75t_L g1612 ( 
.A(n_1495),
.Y(n_1612)
);

HB1xp67_ASAP7_75t_L g1613 ( 
.A(n_1449),
.Y(n_1613)
);

NAND2xp5_ASAP7_75t_SL g1614 ( 
.A(n_1447),
.B(n_1394),
.Y(n_1614)
);

NOR2xp33_ASAP7_75t_L g1615 ( 
.A(n_1458),
.B(n_1041),
.Y(n_1615)
);

INVx2_ASAP7_75t_SL g1616 ( 
.A(n_1521),
.Y(n_1616)
);

INVx2_ASAP7_75t_SL g1617 ( 
.A(n_1570),
.Y(n_1617)
);

OR2x2_ASAP7_75t_L g1618 ( 
.A(n_1550),
.B(n_1197),
.Y(n_1618)
);

NAND2xp5_ASAP7_75t_L g1619 ( 
.A(n_1448),
.B(n_1417),
.Y(n_1619)
);

INVx1_ASAP7_75t_L g1620 ( 
.A(n_1464),
.Y(n_1620)
);

INVx1_ASAP7_75t_L g1621 ( 
.A(n_1470),
.Y(n_1621)
);

OR2x2_ASAP7_75t_L g1622 ( 
.A(n_1522),
.B(n_1200),
.Y(n_1622)
);

INVx2_ASAP7_75t_L g1623 ( 
.A(n_1463),
.Y(n_1623)
);

NAND2xp5_ASAP7_75t_L g1624 ( 
.A(n_1462),
.B(n_1398),
.Y(n_1624)
);

INVx2_ASAP7_75t_L g1625 ( 
.A(n_1469),
.Y(n_1625)
);

NOR2xp33_ASAP7_75t_L g1626 ( 
.A(n_1504),
.B(n_1086),
.Y(n_1626)
);

INVx5_ASAP7_75t_L g1627 ( 
.A(n_1460),
.Y(n_1627)
);

INVx3_ASAP7_75t_L g1628 ( 
.A(n_1510),
.Y(n_1628)
);

AND2x2_ASAP7_75t_L g1629 ( 
.A(n_1504),
.B(n_1247),
.Y(n_1629)
);

BUFx2_ASAP7_75t_L g1630 ( 
.A(n_1473),
.Y(n_1630)
);

INVx1_ASAP7_75t_L g1631 ( 
.A(n_1474),
.Y(n_1631)
);

NAND2xp5_ASAP7_75t_L g1632 ( 
.A(n_1524),
.B(n_1398),
.Y(n_1632)
);

INVx3_ASAP7_75t_L g1633 ( 
.A(n_1510),
.Y(n_1633)
);

BUFx3_ASAP7_75t_L g1634 ( 
.A(n_1454),
.Y(n_1634)
);

NAND2xp5_ASAP7_75t_L g1635 ( 
.A(n_1524),
.B(n_1399),
.Y(n_1635)
);

AND2x4_ASAP7_75t_L g1636 ( 
.A(n_1490),
.B(n_1395),
.Y(n_1636)
);

INVx3_ASAP7_75t_L g1637 ( 
.A(n_1560),
.Y(n_1637)
);

CKINVDCx5p33_ASAP7_75t_R g1638 ( 
.A(n_1540),
.Y(n_1638)
);

INVx2_ASAP7_75t_L g1639 ( 
.A(n_1479),
.Y(n_1639)
);

INVx1_ASAP7_75t_L g1640 ( 
.A(n_1484),
.Y(n_1640)
);

INVx1_ASAP7_75t_L g1641 ( 
.A(n_1486),
.Y(n_1641)
);

BUFx2_ASAP7_75t_L g1642 ( 
.A(n_1473),
.Y(n_1642)
);

INVx2_ASAP7_75t_L g1643 ( 
.A(n_1482),
.Y(n_1643)
);

INVx1_ASAP7_75t_SL g1644 ( 
.A(n_1577),
.Y(n_1644)
);

NAND2xp5_ASAP7_75t_SL g1645 ( 
.A(n_1488),
.B(n_1403),
.Y(n_1645)
);

BUFx3_ASAP7_75t_L g1646 ( 
.A(n_1446),
.Y(n_1646)
);

NOR2xp33_ASAP7_75t_L g1647 ( 
.A(n_1444),
.B(n_1086),
.Y(n_1647)
);

INVx1_ASAP7_75t_L g1648 ( 
.A(n_1493),
.Y(n_1648)
);

INVx1_ASAP7_75t_L g1649 ( 
.A(n_1494),
.Y(n_1649)
);

INVx2_ASAP7_75t_L g1650 ( 
.A(n_1483),
.Y(n_1650)
);

INVx2_ASAP7_75t_L g1651 ( 
.A(n_1485),
.Y(n_1651)
);

BUFx6f_ASAP7_75t_L g1652 ( 
.A(n_1495),
.Y(n_1652)
);

INVx2_ASAP7_75t_SL g1653 ( 
.A(n_1578),
.Y(n_1653)
);

INVx8_ASAP7_75t_L g1654 ( 
.A(n_1576),
.Y(n_1654)
);

INVx8_ASAP7_75t_L g1655 ( 
.A(n_1576),
.Y(n_1655)
);

INVx2_ASAP7_75t_L g1656 ( 
.A(n_1499),
.Y(n_1656)
);

NAND2xp5_ASAP7_75t_SL g1657 ( 
.A(n_1543),
.B(n_1517),
.Y(n_1657)
);

AND2x2_ASAP7_75t_L g1658 ( 
.A(n_1480),
.B(n_1270),
.Y(n_1658)
);

INVx4_ASAP7_75t_L g1659 ( 
.A(n_1582),
.Y(n_1659)
);

AND2x4_ASAP7_75t_L g1660 ( 
.A(n_1513),
.B(n_1404),
.Y(n_1660)
);

AO22x2_ASAP7_75t_L g1661 ( 
.A1(n_1475),
.A2(n_1595),
.B1(n_1471),
.B2(n_1528),
.Y(n_1661)
);

NAND2xp5_ASAP7_75t_SL g1662 ( 
.A(n_1534),
.B(n_1572),
.Y(n_1662)
);

AOI22x1_ASAP7_75t_L g1663 ( 
.A1(n_1527),
.A2(n_1409),
.B1(n_1410),
.B2(n_1408),
.Y(n_1663)
);

INVx1_ASAP7_75t_L g1664 ( 
.A(n_1496),
.Y(n_1664)
);

AND2x4_ASAP7_75t_L g1665 ( 
.A(n_1549),
.B(n_1411),
.Y(n_1665)
);

HB1xp67_ASAP7_75t_L g1666 ( 
.A(n_1519),
.Y(n_1666)
);

INVx3_ASAP7_75t_L g1667 ( 
.A(n_1560),
.Y(n_1667)
);

INVx2_ASAP7_75t_L g1668 ( 
.A(n_1506),
.Y(n_1668)
);

NAND2xp5_ASAP7_75t_L g1669 ( 
.A(n_1527),
.B(n_1399),
.Y(n_1669)
);

INVx1_ASAP7_75t_SL g1670 ( 
.A(n_1466),
.Y(n_1670)
);

AND2x2_ASAP7_75t_L g1671 ( 
.A(n_1572),
.B(n_1046),
.Y(n_1671)
);

OAI22xp5_ASAP7_75t_L g1672 ( 
.A1(n_1544),
.A2(n_1476),
.B1(n_1537),
.B2(n_1452),
.Y(n_1672)
);

NAND2xp5_ASAP7_75t_SL g1673 ( 
.A(n_1545),
.B(n_1552),
.Y(n_1673)
);

BUFx2_ASAP7_75t_L g1674 ( 
.A(n_1547),
.Y(n_1674)
);

AND2x2_ASAP7_75t_L g1675 ( 
.A(n_1590),
.B(n_1190),
.Y(n_1675)
);

NOR2xp33_ASAP7_75t_L g1676 ( 
.A(n_1444),
.B(n_1106),
.Y(n_1676)
);

OR2x2_ASAP7_75t_L g1677 ( 
.A(n_1547),
.B(n_1420),
.Y(n_1677)
);

INVxp67_ASAP7_75t_L g1678 ( 
.A(n_1590),
.Y(n_1678)
);

INVxp67_ASAP7_75t_SL g1679 ( 
.A(n_1460),
.Y(n_1679)
);

BUFx4f_ASAP7_75t_L g1680 ( 
.A(n_1467),
.Y(n_1680)
);

AND2x4_ASAP7_75t_L g1681 ( 
.A(n_1579),
.B(n_1423),
.Y(n_1681)
);

AND2x4_ASAP7_75t_L g1682 ( 
.A(n_1526),
.B(n_1423),
.Y(n_1682)
);

OR2x6_ASAP7_75t_L g1683 ( 
.A(n_1565),
.B(n_1119),
.Y(n_1683)
);

NAND2xp5_ASAP7_75t_L g1684 ( 
.A(n_1478),
.B(n_1481),
.Y(n_1684)
);

BUFx3_ASAP7_75t_L g1685 ( 
.A(n_1468),
.Y(n_1685)
);

AND2x4_ASAP7_75t_L g1686 ( 
.A(n_1531),
.B(n_1418),
.Y(n_1686)
);

NAND2x1p5_ASAP7_75t_L g1687 ( 
.A(n_1582),
.B(n_1407),
.Y(n_1687)
);

AND2x2_ASAP7_75t_L g1688 ( 
.A(n_1592),
.B(n_1190),
.Y(n_1688)
);

AND2x6_ASAP7_75t_L g1689 ( 
.A(n_1460),
.B(n_1407),
.Y(n_1689)
);

INVx3_ASAP7_75t_L g1690 ( 
.A(n_1591),
.Y(n_1690)
);

NAND2xp5_ASAP7_75t_L g1691 ( 
.A(n_1523),
.B(n_1412),
.Y(n_1691)
);

BUFx6f_ASAP7_75t_L g1692 ( 
.A(n_1582),
.Y(n_1692)
);

AND2x4_ASAP7_75t_L g1693 ( 
.A(n_1538),
.B(n_1412),
.Y(n_1693)
);

INVx1_ASAP7_75t_L g1694 ( 
.A(n_1497),
.Y(n_1694)
);

NAND2xp5_ASAP7_75t_L g1695 ( 
.A(n_1465),
.B(n_1421),
.Y(n_1695)
);

AND2x4_ASAP7_75t_L g1696 ( 
.A(n_1539),
.B(n_1421),
.Y(n_1696)
);

INVx2_ASAP7_75t_L g1697 ( 
.A(n_1511),
.Y(n_1697)
);

INVx1_ASAP7_75t_L g1698 ( 
.A(n_1498),
.Y(n_1698)
);

AND2x2_ASAP7_75t_L g1699 ( 
.A(n_1592),
.B(n_1195),
.Y(n_1699)
);

INVx4_ASAP7_75t_L g1700 ( 
.A(n_1582),
.Y(n_1700)
);

NAND2xp5_ASAP7_75t_L g1701 ( 
.A(n_1489),
.B(n_1427),
.Y(n_1701)
);

NAND2xp5_ASAP7_75t_L g1702 ( 
.A(n_1453),
.B(n_1427),
.Y(n_1702)
);

BUFx6f_ASAP7_75t_L g1703 ( 
.A(n_1460),
.Y(n_1703)
);

INVx1_ASAP7_75t_L g1704 ( 
.A(n_1500),
.Y(n_1704)
);

OAI22xp5_ASAP7_75t_L g1705 ( 
.A1(n_1544),
.A2(n_1010),
.B1(n_1019),
.B2(n_1005),
.Y(n_1705)
);

AND2x4_ASAP7_75t_L g1706 ( 
.A(n_1541),
.B(n_1546),
.Y(n_1706)
);

BUFx10_ASAP7_75t_L g1707 ( 
.A(n_1537),
.Y(n_1707)
);

INVx3_ASAP7_75t_L g1708 ( 
.A(n_1591),
.Y(n_1708)
);

NOR2x1p5_ASAP7_75t_L g1709 ( 
.A(n_1566),
.B(n_1169),
.Y(n_1709)
);

NOR2xp33_ASAP7_75t_L g1710 ( 
.A(n_1477),
.B(n_1106),
.Y(n_1710)
);

INVx1_ASAP7_75t_L g1711 ( 
.A(n_1502),
.Y(n_1711)
);

INVxp67_ASAP7_75t_L g1712 ( 
.A(n_1548),
.Y(n_1712)
);

AO21x2_ASAP7_75t_L g1713 ( 
.A1(n_1505),
.A2(n_1439),
.B(n_1435),
.Y(n_1713)
);

NAND2xp5_ASAP7_75t_L g1714 ( 
.A(n_1615),
.B(n_1619),
.Y(n_1714)
);

NAND2xp5_ASAP7_75t_L g1715 ( 
.A(n_1615),
.B(n_1467),
.Y(n_1715)
);

NAND2xp5_ASAP7_75t_L g1716 ( 
.A(n_1619),
.B(n_1467),
.Y(n_1716)
);

INVx1_ASAP7_75t_L g1717 ( 
.A(n_1606),
.Y(n_1717)
);

NAND2xp5_ASAP7_75t_L g1718 ( 
.A(n_1678),
.B(n_1467),
.Y(n_1718)
);

AND2x2_ASAP7_75t_L g1719 ( 
.A(n_1671),
.B(n_1477),
.Y(n_1719)
);

NOR2xp33_ASAP7_75t_L g1720 ( 
.A(n_1678),
.B(n_1445),
.Y(n_1720)
);

NAND2xp5_ASAP7_75t_L g1721 ( 
.A(n_1662),
.B(n_1467),
.Y(n_1721)
);

INVx1_ASAP7_75t_L g1722 ( 
.A(n_1611),
.Y(n_1722)
);

NOR2xp33_ASAP7_75t_SL g1723 ( 
.A(n_1670),
.B(n_1557),
.Y(n_1723)
);

AOI22xp33_ASAP7_75t_L g1724 ( 
.A1(n_1647),
.A2(n_1476),
.B1(n_1595),
.B2(n_1514),
.Y(n_1724)
);

NOR2xp33_ASAP7_75t_L g1725 ( 
.A(n_1712),
.B(n_1445),
.Y(n_1725)
);

INVx1_ASAP7_75t_L g1726 ( 
.A(n_1620),
.Y(n_1726)
);

NAND2xp5_ASAP7_75t_L g1727 ( 
.A(n_1626),
.B(n_1507),
.Y(n_1727)
);

NAND2xp5_ASAP7_75t_L g1728 ( 
.A(n_1626),
.B(n_1520),
.Y(n_1728)
);

INVx1_ASAP7_75t_L g1729 ( 
.A(n_1621),
.Y(n_1729)
);

NAND2xp5_ASAP7_75t_L g1730 ( 
.A(n_1684),
.B(n_1657),
.Y(n_1730)
);

NAND2xp5_ASAP7_75t_L g1731 ( 
.A(n_1684),
.B(n_1525),
.Y(n_1731)
);

CKINVDCx5p33_ASAP7_75t_R g1732 ( 
.A(n_1638),
.Y(n_1732)
);

NOR2xp67_ASAP7_75t_SL g1733 ( 
.A(n_1627),
.B(n_1195),
.Y(n_1733)
);

OR2x2_ASAP7_75t_L g1734 ( 
.A(n_1622),
.B(n_1456),
.Y(n_1734)
);

NAND2xp5_ASAP7_75t_L g1735 ( 
.A(n_1679),
.B(n_1564),
.Y(n_1735)
);

OAI22xp5_ASAP7_75t_L g1736 ( 
.A1(n_1672),
.A2(n_1492),
.B1(n_1512),
.B2(n_1501),
.Y(n_1736)
);

INVx1_ASAP7_75t_L g1737 ( 
.A(n_1631),
.Y(n_1737)
);

NAND2xp5_ASAP7_75t_SL g1738 ( 
.A(n_1627),
.B(n_1554),
.Y(n_1738)
);

NOR2xp33_ASAP7_75t_L g1739 ( 
.A(n_1712),
.B(n_1456),
.Y(n_1739)
);

INVx2_ASAP7_75t_L g1740 ( 
.A(n_1703),
.Y(n_1740)
);

INVx1_ASAP7_75t_L g1741 ( 
.A(n_1640),
.Y(n_1741)
);

O2A1O1Ixp33_ASAP7_75t_L g1742 ( 
.A1(n_1672),
.A2(n_1587),
.B(n_1536),
.C(n_1515),
.Y(n_1742)
);

NAND2xp33_ASAP7_75t_SL g1743 ( 
.A(n_1674),
.B(n_1540),
.Y(n_1743)
);

NAND2xp5_ASAP7_75t_SL g1744 ( 
.A(n_1627),
.B(n_1554),
.Y(n_1744)
);

AOI22xp5_ASAP7_75t_SL g1745 ( 
.A1(n_1705),
.A2(n_1019),
.B1(n_1558),
.B2(n_1575),
.Y(n_1745)
);

NAND3xp33_ASAP7_75t_SL g1746 ( 
.A(n_1647),
.B(n_1396),
.C(n_1552),
.Y(n_1746)
);

INVx1_ASAP7_75t_L g1747 ( 
.A(n_1641),
.Y(n_1747)
);

NAND2xp5_ASAP7_75t_SL g1748 ( 
.A(n_1632),
.B(n_1461),
.Y(n_1748)
);

INVx3_ASAP7_75t_L g1749 ( 
.A(n_1603),
.Y(n_1749)
);

INVx1_ASAP7_75t_L g1750 ( 
.A(n_1648),
.Y(n_1750)
);

AOI22xp5_ASAP7_75t_L g1751 ( 
.A1(n_1676),
.A2(n_1548),
.B1(n_1574),
.B2(n_1567),
.Y(n_1751)
);

INVx1_ASAP7_75t_L g1752 ( 
.A(n_1649),
.Y(n_1752)
);

INVx1_ASAP7_75t_L g1753 ( 
.A(n_1664),
.Y(n_1753)
);

AND2x2_ASAP7_75t_L g1754 ( 
.A(n_1617),
.B(n_1551),
.Y(n_1754)
);

NAND2xp5_ASAP7_75t_L g1755 ( 
.A(n_1679),
.B(n_1580),
.Y(n_1755)
);

HB1xp67_ASAP7_75t_L g1756 ( 
.A(n_1596),
.Y(n_1756)
);

AOI22xp33_ASAP7_75t_L g1757 ( 
.A1(n_1676),
.A2(n_1584),
.B1(n_1594),
.B2(n_1576),
.Y(n_1757)
);

NOR2xp33_ASAP7_75t_L g1758 ( 
.A(n_1666),
.B(n_1644),
.Y(n_1758)
);

NOR2xp33_ASAP7_75t_SL g1759 ( 
.A(n_1670),
.B(n_1532),
.Y(n_1759)
);

A2O1A1Ixp33_ASAP7_75t_L g1760 ( 
.A1(n_1710),
.A2(n_1569),
.B(n_1583),
.C(n_1565),
.Y(n_1760)
);

OAI22xp5_ASAP7_75t_SL g1761 ( 
.A1(n_1705),
.A2(n_1555),
.B1(n_933),
.B2(n_941),
.Y(n_1761)
);

NAND2xp5_ASAP7_75t_SL g1762 ( 
.A(n_1632),
.B(n_1635),
.Y(n_1762)
);

AND2x2_ASAP7_75t_L g1763 ( 
.A(n_1629),
.B(n_1658),
.Y(n_1763)
);

AOI22xp5_ASAP7_75t_L g1764 ( 
.A1(n_1710),
.A2(n_1583),
.B1(n_1576),
.B2(n_1519),
.Y(n_1764)
);

NAND2xp5_ASAP7_75t_L g1765 ( 
.A(n_1624),
.B(n_1576),
.Y(n_1765)
);

INVx2_ASAP7_75t_L g1766 ( 
.A(n_1703),
.Y(n_1766)
);

INVx2_ASAP7_75t_L g1767 ( 
.A(n_1703),
.Y(n_1767)
);

NAND2xp5_ASAP7_75t_SL g1768 ( 
.A(n_1635),
.B(n_1461),
.Y(n_1768)
);

AND2x2_ASAP7_75t_L g1769 ( 
.A(n_1666),
.B(n_918),
.Y(n_1769)
);

INVx2_ASAP7_75t_L g1770 ( 
.A(n_1597),
.Y(n_1770)
);

INVx1_ASAP7_75t_L g1771 ( 
.A(n_1694),
.Y(n_1771)
);

OAI22xp5_ASAP7_75t_L g1772 ( 
.A1(n_1680),
.A2(n_1461),
.B1(n_1508),
.B2(n_1472),
.Y(n_1772)
);

NAND2xp5_ASAP7_75t_SL g1773 ( 
.A(n_1680),
.B(n_1461),
.Y(n_1773)
);

OAI22xp33_ASAP7_75t_L g1774 ( 
.A1(n_1609),
.A2(n_1229),
.B1(n_1246),
.B2(n_1209),
.Y(n_1774)
);

BUFx6f_ASAP7_75t_L g1775 ( 
.A(n_1598),
.Y(n_1775)
);

AOI22xp33_ASAP7_75t_L g1776 ( 
.A1(n_1661),
.A2(n_1562),
.B1(n_1508),
.B2(n_1515),
.Y(n_1776)
);

AOI22xp33_ASAP7_75t_L g1777 ( 
.A1(n_1661),
.A2(n_1562),
.B1(n_1536),
.B2(n_1556),
.Y(n_1777)
);

BUFx3_ASAP7_75t_L g1778 ( 
.A(n_1605),
.Y(n_1778)
);

NOR2xp33_ASAP7_75t_L g1779 ( 
.A(n_1644),
.B(n_1209),
.Y(n_1779)
);

AOI22xp33_ASAP7_75t_L g1780 ( 
.A1(n_1661),
.A2(n_1556),
.B1(n_1529),
.B2(n_1530),
.Y(n_1780)
);

NAND2xp5_ASAP7_75t_L g1781 ( 
.A(n_1624),
.B(n_1518),
.Y(n_1781)
);

NAND2xp5_ASAP7_75t_L g1782 ( 
.A(n_1608),
.B(n_1614),
.Y(n_1782)
);

NAND2xp5_ASAP7_75t_L g1783 ( 
.A(n_1714),
.B(n_1616),
.Y(n_1783)
);

NAND2xp5_ASAP7_75t_SL g1784 ( 
.A(n_1715),
.B(n_1727),
.Y(n_1784)
);

INVx3_ASAP7_75t_L g1785 ( 
.A(n_1749),
.Y(n_1785)
);

NAND2xp5_ASAP7_75t_L g1786 ( 
.A(n_1728),
.B(n_1698),
.Y(n_1786)
);

INVx2_ASAP7_75t_L g1787 ( 
.A(n_1770),
.Y(n_1787)
);

AND2x2_ASAP7_75t_L g1788 ( 
.A(n_1730),
.B(n_1602),
.Y(n_1788)
);

BUFx6f_ASAP7_75t_L g1789 ( 
.A(n_1775),
.Y(n_1789)
);

INVx1_ASAP7_75t_L g1790 ( 
.A(n_1717),
.Y(n_1790)
);

INVx2_ASAP7_75t_L g1791 ( 
.A(n_1770),
.Y(n_1791)
);

AOI22xp33_ASAP7_75t_L g1792 ( 
.A1(n_1739),
.A2(n_1602),
.B1(n_1673),
.B2(n_1707),
.Y(n_1792)
);

CKINVDCx5p33_ASAP7_75t_R g1793 ( 
.A(n_1732),
.Y(n_1793)
);

NOR2x1p5_ASAP7_75t_L g1794 ( 
.A(n_1746),
.B(n_1685),
.Y(n_1794)
);

CKINVDCx20_ASAP7_75t_R g1795 ( 
.A(n_1778),
.Y(n_1795)
);

INVx1_ASAP7_75t_L g1796 ( 
.A(n_1722),
.Y(n_1796)
);

NAND2xp5_ASAP7_75t_L g1797 ( 
.A(n_1731),
.B(n_1704),
.Y(n_1797)
);

AOI22xp33_ASAP7_75t_L g1798 ( 
.A1(n_1739),
.A2(n_1602),
.B1(n_1707),
.B2(n_1706),
.Y(n_1798)
);

INVxp67_ASAP7_75t_SL g1799 ( 
.A(n_1738),
.Y(n_1799)
);

INVx4_ASAP7_75t_L g1800 ( 
.A(n_1775),
.Y(n_1800)
);

AND3x1_ASAP7_75t_SL g1801 ( 
.A(n_1745),
.B(n_1219),
.C(n_1709),
.Y(n_1801)
);

INVx1_ASAP7_75t_L g1802 ( 
.A(n_1726),
.Y(n_1802)
);

BUFx4f_ASAP7_75t_L g1803 ( 
.A(n_1775),
.Y(n_1803)
);

INVx2_ASAP7_75t_L g1804 ( 
.A(n_1729),
.Y(n_1804)
);

NAND2xp5_ASAP7_75t_L g1805 ( 
.A(n_1720),
.B(n_1711),
.Y(n_1805)
);

INVx1_ASAP7_75t_L g1806 ( 
.A(n_1737),
.Y(n_1806)
);

NAND2xp5_ASAP7_75t_SL g1807 ( 
.A(n_1764),
.B(n_1677),
.Y(n_1807)
);

BUFx6f_ASAP7_75t_L g1808 ( 
.A(n_1775),
.Y(n_1808)
);

INVx1_ASAP7_75t_L g1809 ( 
.A(n_1741),
.Y(n_1809)
);

INVx2_ASAP7_75t_SL g1810 ( 
.A(n_1778),
.Y(n_1810)
);

BUFx10_ASAP7_75t_L g1811 ( 
.A(n_1779),
.Y(n_1811)
);

AND2x6_ASAP7_75t_SL g1812 ( 
.A(n_1779),
.B(n_1683),
.Y(n_1812)
);

INVx1_ASAP7_75t_L g1813 ( 
.A(n_1747),
.Y(n_1813)
);

NAND2xp5_ASAP7_75t_L g1814 ( 
.A(n_1720),
.B(n_1675),
.Y(n_1814)
);

NAND2xp5_ASAP7_75t_L g1815 ( 
.A(n_1725),
.B(n_1688),
.Y(n_1815)
);

AND2x4_ASAP7_75t_L g1816 ( 
.A(n_1750),
.B(n_1706),
.Y(n_1816)
);

INVx2_ASAP7_75t_L g1817 ( 
.A(n_1752),
.Y(n_1817)
);

INVx4_ASAP7_75t_L g1818 ( 
.A(n_1749),
.Y(n_1818)
);

BUFx2_ASAP7_75t_L g1819 ( 
.A(n_1756),
.Y(n_1819)
);

INVx3_ASAP7_75t_L g1820 ( 
.A(n_1740),
.Y(n_1820)
);

A2O1A1Ixp33_ASAP7_75t_L g1821 ( 
.A1(n_1742),
.A2(n_1699),
.B(n_1645),
.C(n_1655),
.Y(n_1821)
);

BUFx2_ASAP7_75t_L g1822 ( 
.A(n_1763),
.Y(n_1822)
);

OAI21xp5_ASAP7_75t_L g1823 ( 
.A1(n_1736),
.A2(n_1695),
.B(n_1691),
.Y(n_1823)
);

AOI22xp5_ASAP7_75t_L g1824 ( 
.A1(n_1719),
.A2(n_1246),
.B1(n_1229),
.B2(n_1613),
.Y(n_1824)
);

CKINVDCx5p33_ASAP7_75t_R g1825 ( 
.A(n_1758),
.Y(n_1825)
);

NAND2xp5_ASAP7_75t_L g1826 ( 
.A(n_1725),
.B(n_1653),
.Y(n_1826)
);

NOR2xp33_ASAP7_75t_R g1827 ( 
.A(n_1743),
.B(n_1646),
.Y(n_1827)
);

NOR2xp33_ASAP7_75t_L g1828 ( 
.A(n_1734),
.B(n_1607),
.Y(n_1828)
);

NAND2xp5_ASAP7_75t_L g1829 ( 
.A(n_1735),
.B(n_1681),
.Y(n_1829)
);

BUFx6f_ASAP7_75t_L g1830 ( 
.A(n_1740),
.Y(n_1830)
);

INVxp67_ASAP7_75t_L g1831 ( 
.A(n_1819),
.Y(n_1831)
);

INVxp67_ASAP7_75t_L g1832 ( 
.A(n_1822),
.Y(n_1832)
);

CKINVDCx16_ASAP7_75t_R g1833 ( 
.A(n_1795),
.Y(n_1833)
);

BUFx6f_ASAP7_75t_L g1834 ( 
.A(n_1803),
.Y(n_1834)
);

AOI33xp33_ASAP7_75t_L g1835 ( 
.A1(n_1792),
.A2(n_1769),
.A3(n_1099),
.B1(n_1096),
.B2(n_1098),
.B3(n_1094),
.Y(n_1835)
);

OAI21xp5_ASAP7_75t_L g1836 ( 
.A1(n_1821),
.A2(n_1716),
.B(n_1765),
.Y(n_1836)
);

AOI21xp5_ASAP7_75t_L g1837 ( 
.A1(n_1823),
.A2(n_1744),
.B(n_1738),
.Y(n_1837)
);

INVx2_ASAP7_75t_SL g1838 ( 
.A(n_1810),
.Y(n_1838)
);

INVx2_ASAP7_75t_L g1839 ( 
.A(n_1804),
.Y(n_1839)
);

AND2x2_ASAP7_75t_L g1840 ( 
.A(n_1828),
.B(n_1758),
.Y(n_1840)
);

INVx2_ASAP7_75t_L g1841 ( 
.A(n_1804),
.Y(n_1841)
);

INVx1_ASAP7_75t_L g1842 ( 
.A(n_1817),
.Y(n_1842)
);

INVx1_ASAP7_75t_L g1843 ( 
.A(n_1817),
.Y(n_1843)
);

INVx1_ASAP7_75t_L g1844 ( 
.A(n_1790),
.Y(n_1844)
);

BUFx2_ASAP7_75t_SL g1845 ( 
.A(n_1795),
.Y(n_1845)
);

O2A1O1Ixp33_ASAP7_75t_L g1846 ( 
.A1(n_1821),
.A2(n_1760),
.B(n_1774),
.C(n_1613),
.Y(n_1846)
);

AOI22xp5_ASAP7_75t_L g1847 ( 
.A1(n_1814),
.A2(n_1723),
.B1(n_1751),
.B2(n_1761),
.Y(n_1847)
);

CKINVDCx14_ASAP7_75t_R g1848 ( 
.A(n_1793),
.Y(n_1848)
);

INVx5_ASAP7_75t_L g1849 ( 
.A(n_1789),
.Y(n_1849)
);

NAND2xp5_ASAP7_75t_SL g1850 ( 
.A(n_1825),
.B(n_1760),
.Y(n_1850)
);

OAI22xp5_ASAP7_75t_L g1851 ( 
.A1(n_1786),
.A2(n_1724),
.B1(n_1757),
.B2(n_1776),
.Y(n_1851)
);

NAND2xp5_ASAP7_75t_L g1852 ( 
.A(n_1805),
.B(n_1762),
.Y(n_1852)
);

NAND2xp5_ASAP7_75t_SL g1853 ( 
.A(n_1825),
.B(n_1618),
.Y(n_1853)
);

INVx1_ASAP7_75t_L g1854 ( 
.A(n_1796),
.Y(n_1854)
);

AND2x2_ASAP7_75t_L g1855 ( 
.A(n_1788),
.B(n_1754),
.Y(n_1855)
);

INVx2_ASAP7_75t_L g1856 ( 
.A(n_1787),
.Y(n_1856)
);

NAND2xp5_ASAP7_75t_L g1857 ( 
.A(n_1797),
.B(n_1762),
.Y(n_1857)
);

O2A1O1Ixp33_ASAP7_75t_L g1858 ( 
.A1(n_1815),
.A2(n_1683),
.B(n_1782),
.C(n_1718),
.Y(n_1858)
);

NAND2xp5_ASAP7_75t_SL g1859 ( 
.A(n_1783),
.B(n_1721),
.Y(n_1859)
);

INVx1_ASAP7_75t_L g1860 ( 
.A(n_1802),
.Y(n_1860)
);

AOI21xp5_ASAP7_75t_L g1861 ( 
.A1(n_1807),
.A2(n_1744),
.B(n_1773),
.Y(n_1861)
);

AOI21xp5_ASAP7_75t_L g1862 ( 
.A1(n_1807),
.A2(n_1773),
.B(n_1772),
.Y(n_1862)
);

INVx2_ASAP7_75t_L g1863 ( 
.A(n_1787),
.Y(n_1863)
);

A2O1A1Ixp33_ASAP7_75t_L g1864 ( 
.A1(n_1784),
.A2(n_1777),
.B(n_1753),
.C(n_1771),
.Y(n_1864)
);

OR2x6_ASAP7_75t_L g1865 ( 
.A(n_1794),
.B(n_1654),
.Y(n_1865)
);

NAND2xp5_ASAP7_75t_L g1866 ( 
.A(n_1784),
.B(n_1788),
.Y(n_1866)
);

OAI22xp5_ASAP7_75t_L g1867 ( 
.A1(n_1798),
.A2(n_1755),
.B1(n_1683),
.B2(n_1669),
.Y(n_1867)
);

INVx2_ASAP7_75t_L g1868 ( 
.A(n_1791),
.Y(n_1868)
);

INVx1_ASAP7_75t_L g1869 ( 
.A(n_1806),
.Y(n_1869)
);

OR2x2_ASAP7_75t_L g1870 ( 
.A(n_1826),
.B(n_1630),
.Y(n_1870)
);

OAI22x1_ASAP7_75t_L g1871 ( 
.A1(n_1824),
.A2(n_1642),
.B1(n_1596),
.B2(n_1663),
.Y(n_1871)
);

NOR2xp33_ASAP7_75t_L g1872 ( 
.A(n_1793),
.B(n_1634),
.Y(n_1872)
);

AOI22xp5_ASAP7_75t_L g1873 ( 
.A1(n_1811),
.A2(n_1759),
.B1(n_1340),
.B2(n_1733),
.Y(n_1873)
);

INVx2_ASAP7_75t_L g1874 ( 
.A(n_1791),
.Y(n_1874)
);

NAND2xp5_ASAP7_75t_L g1875 ( 
.A(n_1799),
.B(n_1748),
.Y(n_1875)
);

INVx5_ASAP7_75t_L g1876 ( 
.A(n_1789),
.Y(n_1876)
);

INVx1_ASAP7_75t_L g1877 ( 
.A(n_1809),
.Y(n_1877)
);

OR2x6_ASAP7_75t_L g1878 ( 
.A(n_1858),
.B(n_1748),
.Y(n_1878)
);

BUFx8_ASAP7_75t_SL g1879 ( 
.A(n_1865),
.Y(n_1879)
);

AOI22xp33_ASAP7_75t_SL g1880 ( 
.A1(n_1851),
.A2(n_1811),
.B1(n_1007),
.B2(n_1042),
.Y(n_1880)
);

INVx2_ASAP7_75t_L g1881 ( 
.A(n_1839),
.Y(n_1881)
);

O2A1O1Ixp5_ASAP7_75t_L g1882 ( 
.A1(n_1850),
.A2(n_1768),
.B(n_1695),
.C(n_1702),
.Y(n_1882)
);

INVx2_ASAP7_75t_L g1883 ( 
.A(n_1841),
.Y(n_1883)
);

INVx1_ASAP7_75t_L g1884 ( 
.A(n_1844),
.Y(n_1884)
);

AND2x4_ASAP7_75t_L g1885 ( 
.A(n_1865),
.B(n_1810),
.Y(n_1885)
);

NOR2xp33_ASAP7_75t_L g1886 ( 
.A(n_1847),
.B(n_1811),
.Y(n_1886)
);

AND3x1_ASAP7_75t_SL g1887 ( 
.A(n_1854),
.B(n_1812),
.C(n_1509),
.Y(n_1887)
);

INVx1_ASAP7_75t_L g1888 ( 
.A(n_1860),
.Y(n_1888)
);

INVx6_ASAP7_75t_L g1889 ( 
.A(n_1834),
.Y(n_1889)
);

AND2x4_ASAP7_75t_L g1890 ( 
.A(n_1865),
.B(n_1830),
.Y(n_1890)
);

INVx1_ASAP7_75t_L g1891 ( 
.A(n_1869),
.Y(n_1891)
);

INVx6_ASAP7_75t_L g1892 ( 
.A(n_1834),
.Y(n_1892)
);

INVx1_ASAP7_75t_L g1893 ( 
.A(n_1877),
.Y(n_1893)
);

INVx2_ASAP7_75t_L g1894 ( 
.A(n_1842),
.Y(n_1894)
);

INVx2_ASAP7_75t_L g1895 ( 
.A(n_1843),
.Y(n_1895)
);

INVx1_ASAP7_75t_L g1896 ( 
.A(n_1866),
.Y(n_1896)
);

INVx3_ASAP7_75t_L g1897 ( 
.A(n_1834),
.Y(n_1897)
);

HB1xp67_ASAP7_75t_L g1898 ( 
.A(n_1875),
.Y(n_1898)
);

AND2x2_ASAP7_75t_L g1899 ( 
.A(n_1855),
.B(n_1813),
.Y(n_1899)
);

INVx1_ASAP7_75t_SL g1900 ( 
.A(n_1870),
.Y(n_1900)
);

NOR2xp33_ASAP7_75t_R g1901 ( 
.A(n_1848),
.B(n_1553),
.Y(n_1901)
);

AOI221xp5_ASAP7_75t_L g1902 ( 
.A1(n_1851),
.A2(n_785),
.B1(n_788),
.B2(n_784),
.C(n_782),
.Y(n_1902)
);

BUFx2_ASAP7_75t_L g1903 ( 
.A(n_1832),
.Y(n_1903)
);

INVx1_ASAP7_75t_L g1904 ( 
.A(n_1866),
.Y(n_1904)
);

INVx2_ASAP7_75t_L g1905 ( 
.A(n_1856),
.Y(n_1905)
);

INVx1_ASAP7_75t_L g1906 ( 
.A(n_1875),
.Y(n_1906)
);

NAND2xp5_ASAP7_75t_L g1907 ( 
.A(n_1852),
.B(n_1829),
.Y(n_1907)
);

OR2x6_ASAP7_75t_L g1908 ( 
.A(n_1862),
.B(n_1861),
.Y(n_1908)
);

AND2x4_ASAP7_75t_L g1909 ( 
.A(n_1838),
.B(n_1830),
.Y(n_1909)
);

AOI22xp5_ASAP7_75t_L g1910 ( 
.A1(n_1853),
.A2(n_1801),
.B1(n_1816),
.B2(n_1665),
.Y(n_1910)
);

BUFx10_ASAP7_75t_L g1911 ( 
.A(n_1872),
.Y(n_1911)
);

INVx2_ASAP7_75t_SL g1912 ( 
.A(n_1833),
.Y(n_1912)
);

AOI22xp5_ASAP7_75t_L g1913 ( 
.A1(n_1840),
.A2(n_1816),
.B1(n_1665),
.B2(n_1660),
.Y(n_1913)
);

NAND2xp5_ASAP7_75t_SL g1914 ( 
.A(n_1835),
.B(n_1816),
.Y(n_1914)
);

OR2x2_ASAP7_75t_L g1915 ( 
.A(n_1852),
.B(n_1768),
.Y(n_1915)
);

INVx1_ASAP7_75t_L g1916 ( 
.A(n_1863),
.Y(n_1916)
);

AND2x2_ASAP7_75t_L g1917 ( 
.A(n_1845),
.B(n_1820),
.Y(n_1917)
);

NOR2xp33_ASAP7_75t_L g1918 ( 
.A(n_1867),
.B(n_1831),
.Y(n_1918)
);

AOI22xp33_ASAP7_75t_L g1919 ( 
.A1(n_1867),
.A2(n_798),
.B1(n_799),
.B2(n_788),
.Y(n_1919)
);

AOI22xp33_ASAP7_75t_L g1920 ( 
.A1(n_1871),
.A2(n_799),
.B1(n_802),
.B2(n_798),
.Y(n_1920)
);

CKINVDCx11_ASAP7_75t_R g1921 ( 
.A(n_1868),
.Y(n_1921)
);

BUFx8_ASAP7_75t_SL g1922 ( 
.A(n_1874),
.Y(n_1922)
);

NOR2xp33_ASAP7_75t_L g1923 ( 
.A(n_1857),
.B(n_1859),
.Y(n_1923)
);

INVx3_ASAP7_75t_L g1924 ( 
.A(n_1849),
.Y(n_1924)
);

INVx5_ASAP7_75t_L g1925 ( 
.A(n_1849),
.Y(n_1925)
);

NAND2x1p5_ASAP7_75t_L g1926 ( 
.A(n_1849),
.B(n_1803),
.Y(n_1926)
);

AOI221xp5_ASAP7_75t_SL g1927 ( 
.A1(n_1846),
.A2(n_1059),
.B1(n_999),
.B2(n_1081),
.C(n_1080),
.Y(n_1927)
);

INVx4_ASAP7_75t_L g1928 ( 
.A(n_1876),
.Y(n_1928)
);

INVx2_ASAP7_75t_L g1929 ( 
.A(n_1876),
.Y(n_1929)
);

OAI22xp33_ASAP7_75t_L g1930 ( 
.A1(n_1873),
.A2(n_803),
.B1(n_809),
.B2(n_802),
.Y(n_1930)
);

INVx3_ASAP7_75t_L g1931 ( 
.A(n_1876),
.Y(n_1931)
);

INVx1_ASAP7_75t_L g1932 ( 
.A(n_1857),
.Y(n_1932)
);

INVx1_ASAP7_75t_L g1933 ( 
.A(n_1864),
.Y(n_1933)
);

BUFx2_ASAP7_75t_L g1934 ( 
.A(n_1876),
.Y(n_1934)
);

O2A1O1Ixp33_ASAP7_75t_SL g1935 ( 
.A1(n_1902),
.A2(n_1837),
.B(n_1836),
.C(n_1601),
.Y(n_1935)
);

INVx8_ASAP7_75t_L g1936 ( 
.A(n_1922),
.Y(n_1936)
);

AND2x2_ASAP7_75t_L g1937 ( 
.A(n_1918),
.B(n_1836),
.Y(n_1937)
);

CKINVDCx5p33_ASAP7_75t_R g1938 ( 
.A(n_1901),
.Y(n_1938)
);

NAND3xp33_ASAP7_75t_SL g1939 ( 
.A(n_1880),
.B(n_1827),
.C(n_818),
.Y(n_1939)
);

BUFx12f_ASAP7_75t_L g1940 ( 
.A(n_1911),
.Y(n_1940)
);

O2A1O1Ixp33_ASAP7_75t_L g1941 ( 
.A1(n_1930),
.A2(n_1088),
.B(n_1084),
.C(n_858),
.Y(n_1941)
);

INVx1_ASAP7_75t_SL g1942 ( 
.A(n_1921),
.Y(n_1942)
);

OAI22x1_ASAP7_75t_L g1943 ( 
.A1(n_1918),
.A2(n_1886),
.B1(n_1912),
.B2(n_1888),
.Y(n_1943)
);

OAI22xp5_ASAP7_75t_L g1944 ( 
.A1(n_1880),
.A2(n_1919),
.B1(n_1902),
.B2(n_1910),
.Y(n_1944)
);

NOR2x1_ASAP7_75t_SL g1945 ( 
.A(n_1908),
.B(n_1789),
.Y(n_1945)
);

O2A1O1Ixp33_ASAP7_75t_SL g1946 ( 
.A1(n_1930),
.A2(n_859),
.B(n_861),
.C(n_855),
.Y(n_1946)
);

O2A1O1Ixp33_ASAP7_75t_SL g1947 ( 
.A1(n_1914),
.A2(n_863),
.B(n_869),
.C(n_862),
.Y(n_1947)
);

AO31x2_ASAP7_75t_L g1948 ( 
.A1(n_1886),
.A2(n_1702),
.A3(n_1701),
.B(n_1818),
.Y(n_1948)
);

INVx2_ASAP7_75t_L g1949 ( 
.A(n_1894),
.Y(n_1949)
);

O2A1O1Ixp33_ASAP7_75t_SL g1950 ( 
.A1(n_1907),
.A2(n_872),
.B(n_875),
.C(n_870),
.Y(n_1950)
);

A2O1A1Ixp33_ASAP7_75t_L g1951 ( 
.A1(n_1919),
.A2(n_1803),
.B(n_803),
.C(n_818),
.Y(n_1951)
);

AOI21xp5_ASAP7_75t_L g1952 ( 
.A1(n_1908),
.A2(n_1655),
.B(n_1654),
.Y(n_1952)
);

AND2x4_ASAP7_75t_L g1953 ( 
.A(n_1885),
.B(n_1890),
.Y(n_1953)
);

O2A1O1Ixp33_ASAP7_75t_SL g1954 ( 
.A1(n_1907),
.A2(n_879),
.B(n_882),
.C(n_876),
.Y(n_1954)
);

INVx1_ASAP7_75t_L g1955 ( 
.A(n_1898),
.Y(n_1955)
);

AO21x1_ASAP7_75t_L g1956 ( 
.A1(n_1923),
.A2(n_1818),
.B(n_1800),
.Y(n_1956)
);

OAI21x1_ASAP7_75t_L g1957 ( 
.A1(n_1882),
.A2(n_1604),
.B(n_1701),
.Y(n_1957)
);

INVx8_ASAP7_75t_L g1958 ( 
.A(n_1879),
.Y(n_1958)
);

OAI21xp5_ASAP7_75t_L g1959 ( 
.A1(n_1927),
.A2(n_1780),
.B(n_1686),
.Y(n_1959)
);

INVx1_ASAP7_75t_L g1960 ( 
.A(n_1898),
.Y(n_1960)
);

AND2x4_ASAP7_75t_L g1961 ( 
.A(n_1885),
.B(n_1800),
.Y(n_1961)
);

OAI221xp5_ASAP7_75t_L g1962 ( 
.A1(n_1920),
.A2(n_822),
.B1(n_809),
.B2(n_593),
.C(n_598),
.Y(n_1962)
);

A2O1A1Ixp33_ASAP7_75t_L g1963 ( 
.A1(n_1920),
.A2(n_822),
.B(n_993),
.C(n_992),
.Y(n_1963)
);

OAI21x1_ASAP7_75t_L g1964 ( 
.A1(n_1882),
.A2(n_1604),
.B(n_1691),
.Y(n_1964)
);

INVx4_ASAP7_75t_L g1965 ( 
.A(n_1889),
.Y(n_1965)
);

AOI22xp33_ASAP7_75t_L g1966 ( 
.A1(n_1933),
.A2(n_885),
.B1(n_887),
.B2(n_883),
.Y(n_1966)
);

AOI221xp5_ASAP7_75t_L g1967 ( 
.A1(n_1923),
.A2(n_606),
.B1(n_608),
.B2(n_587),
.C(n_586),
.Y(n_1967)
);

INVx2_ASAP7_75t_L g1968 ( 
.A(n_1895),
.Y(n_1968)
);

AOI21xp5_ASAP7_75t_L g1969 ( 
.A1(n_1908),
.A2(n_1655),
.B(n_1654),
.Y(n_1969)
);

OAI21x1_ASAP7_75t_L g1970 ( 
.A1(n_1881),
.A2(n_1883),
.B(n_1905),
.Y(n_1970)
);

INVxp67_ASAP7_75t_SL g1971 ( 
.A(n_1906),
.Y(n_1971)
);

OAI21x1_ASAP7_75t_L g1972 ( 
.A1(n_1916),
.A2(n_1669),
.B(n_1781),
.Y(n_1972)
);

AOI22xp33_ASAP7_75t_L g1973 ( 
.A1(n_1900),
.A2(n_895),
.B1(n_897),
.B2(n_888),
.Y(n_1973)
);

AO31x2_ASAP7_75t_L g1974 ( 
.A1(n_1928),
.A2(n_1659),
.A3(n_1700),
.B(n_1075),
.Y(n_1974)
);

AO32x2_ASAP7_75t_L g1975 ( 
.A1(n_1928),
.A2(n_1713),
.A3(n_1262),
.B1(n_4),
.B2(n_2),
.Y(n_1975)
);

NOR2xp33_ASAP7_75t_L g1976 ( 
.A(n_1911),
.B(n_1532),
.Y(n_1976)
);

AOI22xp33_ASAP7_75t_L g1977 ( 
.A1(n_1878),
.A2(n_900),
.B1(n_901),
.B2(n_898),
.Y(n_1977)
);

BUFx8_ASAP7_75t_L g1978 ( 
.A(n_1903),
.Y(n_1978)
);

BUFx12f_ASAP7_75t_L g1979 ( 
.A(n_1889),
.Y(n_1979)
);

OAI21xp5_ASAP7_75t_L g1980 ( 
.A1(n_1913),
.A2(n_1686),
.B(n_1660),
.Y(n_1980)
);

INVx1_ASAP7_75t_L g1981 ( 
.A(n_1884),
.Y(n_1981)
);

INVx2_ASAP7_75t_L g1982 ( 
.A(n_1891),
.Y(n_1982)
);

A2O1A1Ixp33_ASAP7_75t_L g1983 ( 
.A1(n_1932),
.A2(n_995),
.B(n_998),
.C(n_994),
.Y(n_1983)
);

NAND2xp5_ASAP7_75t_L g1984 ( 
.A(n_1896),
.B(n_1820),
.Y(n_1984)
);

NAND2x1p5_ASAP7_75t_L g1985 ( 
.A(n_1925),
.B(n_1909),
.Y(n_1985)
);

AO32x2_ASAP7_75t_L g1986 ( 
.A1(n_1904),
.A2(n_1713),
.A3(n_6),
.B1(n_3),
.B2(n_5),
.Y(n_1986)
);

O2A1O1Ixp33_ASAP7_75t_SL g1987 ( 
.A1(n_1893),
.A2(n_904),
.B(n_907),
.C(n_902),
.Y(n_1987)
);

AOI21xp5_ASAP7_75t_L g1988 ( 
.A1(n_1925),
.A2(n_1628),
.B(n_1603),
.Y(n_1988)
);

A2O1A1Ixp33_ASAP7_75t_L g1989 ( 
.A1(n_1925),
.A2(n_1001),
.B(n_1003),
.C(n_1000),
.Y(n_1989)
);

INVx1_ASAP7_75t_L g1990 ( 
.A(n_1899),
.Y(n_1990)
);

NOR2xp33_ASAP7_75t_L g1991 ( 
.A(n_1917),
.B(n_1553),
.Y(n_1991)
);

INVxp67_ASAP7_75t_L g1992 ( 
.A(n_1909),
.Y(n_1992)
);

HB1xp67_ASAP7_75t_L g1993 ( 
.A(n_1878),
.Y(n_1993)
);

BUFx3_ASAP7_75t_L g1994 ( 
.A(n_1889),
.Y(n_1994)
);

INVx1_ASAP7_75t_L g1995 ( 
.A(n_1915),
.Y(n_1995)
);

O2A1O1Ixp33_ASAP7_75t_SL g1996 ( 
.A1(n_1929),
.A2(n_912),
.B(n_914),
.C(n_908),
.Y(n_1996)
);

A2O1A1Ixp33_ASAP7_75t_L g1997 ( 
.A1(n_1925),
.A2(n_1006),
.B(n_1009),
.C(n_1004),
.Y(n_1997)
);

AO32x2_ASAP7_75t_L g1998 ( 
.A1(n_1878),
.A2(n_7),
.A3(n_5),
.B1(n_6),
.B2(n_8),
.Y(n_1998)
);

NAND2x1p5_ASAP7_75t_L g1999 ( 
.A(n_1924),
.B(n_1785),
.Y(n_1999)
);

AOI21xp5_ASAP7_75t_L g2000 ( 
.A1(n_1926),
.A2(n_1633),
.B(n_1628),
.Y(n_2000)
);

NOR2xp33_ASAP7_75t_L g2001 ( 
.A(n_1897),
.B(n_1610),
.Y(n_2001)
);

AOI21xp33_ASAP7_75t_L g2002 ( 
.A1(n_1890),
.A2(n_1785),
.B(n_1830),
.Y(n_2002)
);

OAI21xp5_ASAP7_75t_L g2003 ( 
.A1(n_1926),
.A2(n_1013),
.B(n_1012),
.Y(n_2003)
);

O2A1O1Ixp33_ASAP7_75t_L g2004 ( 
.A1(n_1897),
.A2(n_917),
.B(n_919),
.C(n_915),
.Y(n_2004)
);

INVx2_ASAP7_75t_SL g2005 ( 
.A(n_1892),
.Y(n_2005)
);

AO31x2_ASAP7_75t_L g2006 ( 
.A1(n_1934),
.A2(n_1015),
.A3(n_1021),
.B(n_1014),
.Y(n_2006)
);

OAI22xp5_ASAP7_75t_L g2007 ( 
.A1(n_1892),
.A2(n_1785),
.B1(n_1820),
.B2(n_1830),
.Y(n_2007)
);

AO31x2_ASAP7_75t_L g2008 ( 
.A1(n_1887),
.A2(n_1023),
.A3(n_1024),
.B(n_1022),
.Y(n_2008)
);

AND2x4_ASAP7_75t_L g2009 ( 
.A(n_1924),
.B(n_1830),
.Y(n_2009)
);

A2O1A1Ixp33_ASAP7_75t_L g2010 ( 
.A1(n_1887),
.A2(n_1026),
.B(n_1028),
.C(n_1025),
.Y(n_2010)
);

NAND2xp5_ASAP7_75t_L g2011 ( 
.A(n_1892),
.B(n_1931),
.Y(n_2011)
);

INVx2_ASAP7_75t_L g2012 ( 
.A(n_1931),
.Y(n_2012)
);

INVx2_ASAP7_75t_L g2013 ( 
.A(n_1982),
.Y(n_2013)
);

INVx2_ASAP7_75t_L g2014 ( 
.A(n_1981),
.Y(n_2014)
);

INVx2_ASAP7_75t_SL g2015 ( 
.A(n_1978),
.Y(n_2015)
);

INVx3_ASAP7_75t_L g2016 ( 
.A(n_2012),
.Y(n_2016)
);

AOI21xp33_ASAP7_75t_L g2017 ( 
.A1(n_1944),
.A2(n_921),
.B(n_920),
.Y(n_2017)
);

OAI22xp5_ASAP7_75t_L g2018 ( 
.A1(n_1963),
.A2(n_612),
.B1(n_637),
.B2(n_611),
.Y(n_2018)
);

BUFx8_ASAP7_75t_L g2019 ( 
.A(n_1940),
.Y(n_2019)
);

INVx2_ASAP7_75t_L g2020 ( 
.A(n_1949),
.Y(n_2020)
);

INVx1_ASAP7_75t_L g2021 ( 
.A(n_1955),
.Y(n_2021)
);

NAND2xp5_ASAP7_75t_L g2022 ( 
.A(n_1937),
.B(n_923),
.Y(n_2022)
);

INVx1_ASAP7_75t_L g2023 ( 
.A(n_1960),
.Y(n_2023)
);

INVx1_ASAP7_75t_L g2024 ( 
.A(n_1971),
.Y(n_2024)
);

AND2x2_ASAP7_75t_L g2025 ( 
.A(n_1995),
.B(n_925),
.Y(n_2025)
);

OAI22xp5_ASAP7_75t_L g2026 ( 
.A1(n_1951),
.A2(n_655),
.B1(n_670),
.B2(n_650),
.Y(n_2026)
);

OAI22xp33_ASAP7_75t_L g2027 ( 
.A1(n_1939),
.A2(n_678),
.B1(n_689),
.B2(n_676),
.Y(n_2027)
);

OR2x6_ASAP7_75t_SL g2028 ( 
.A(n_1938),
.B(n_691),
.Y(n_2028)
);

INVx1_ASAP7_75t_L g2029 ( 
.A(n_1968),
.Y(n_2029)
);

AND2x4_ASAP7_75t_L g2030 ( 
.A(n_1953),
.B(n_1808),
.Y(n_2030)
);

AOI22xp33_ASAP7_75t_L g2031 ( 
.A1(n_1943),
.A2(n_1289),
.B1(n_705),
.B2(n_710),
.Y(n_2031)
);

CKINVDCx8_ASAP7_75t_R g2032 ( 
.A(n_1958),
.Y(n_2032)
);

OAI22xp5_ASAP7_75t_L g2033 ( 
.A1(n_1977),
.A2(n_712),
.B1(n_714),
.B2(n_702),
.Y(n_2033)
);

BUFx12f_ASAP7_75t_L g2034 ( 
.A(n_1979),
.Y(n_2034)
);

OAI22xp5_ASAP7_75t_L g2035 ( 
.A1(n_1966),
.A2(n_721),
.B1(n_722),
.B2(n_716),
.Y(n_2035)
);

OAI22xp5_ASAP7_75t_L g2036 ( 
.A1(n_1962),
.A2(n_740),
.B1(n_742),
.B2(n_726),
.Y(n_2036)
);

AND2x4_ASAP7_75t_L g2037 ( 
.A(n_1953),
.B(n_1789),
.Y(n_2037)
);

NAND2x1p5_ASAP7_75t_L g2038 ( 
.A(n_1965),
.B(n_2009),
.Y(n_2038)
);

INVx2_ASAP7_75t_SL g2039 ( 
.A(n_1936),
.Y(n_2039)
);

INVx1_ASAP7_75t_SL g2040 ( 
.A(n_2011),
.Y(n_2040)
);

NAND2x1p5_ASAP7_75t_L g2041 ( 
.A(n_2009),
.B(n_1808),
.Y(n_2041)
);

BUFx2_ASAP7_75t_L g2042 ( 
.A(n_1992),
.Y(n_2042)
);

AOI21xp33_ASAP7_75t_L g2043 ( 
.A1(n_1993),
.A2(n_1289),
.B(n_1284),
.Y(n_2043)
);

OAI22xp5_ASAP7_75t_L g2044 ( 
.A1(n_1990),
.A2(n_746),
.B1(n_749),
.B2(n_743),
.Y(n_2044)
);

INVx2_ASAP7_75t_L g2045 ( 
.A(n_1970),
.Y(n_2045)
);

CKINVDCx5p33_ASAP7_75t_R g2046 ( 
.A(n_1958),
.Y(n_2046)
);

INVx1_ASAP7_75t_L g2047 ( 
.A(n_1984),
.Y(n_2047)
);

INVx2_ASAP7_75t_L g2048 ( 
.A(n_1985),
.Y(n_2048)
);

INVx1_ASAP7_75t_L g2049 ( 
.A(n_1948),
.Y(n_2049)
);

INVx2_ASAP7_75t_SL g2050 ( 
.A(n_1936),
.Y(n_2050)
);

INVx1_ASAP7_75t_L g2051 ( 
.A(n_1948),
.Y(n_2051)
);

CKINVDCx11_ASAP7_75t_R g2052 ( 
.A(n_1942),
.Y(n_2052)
);

OAI22xp5_ASAP7_75t_L g2053 ( 
.A1(n_1998),
.A2(n_763),
.B1(n_766),
.B2(n_760),
.Y(n_2053)
);

AOI22xp5_ASAP7_75t_L g2054 ( 
.A1(n_1935),
.A2(n_773),
.B1(n_767),
.B2(n_498),
.Y(n_2054)
);

OAI221xp5_ASAP7_75t_L g2055 ( 
.A1(n_1967),
.A2(n_503),
.B1(n_505),
.B2(n_501),
.C(n_496),
.Y(n_2055)
);

BUFx6f_ASAP7_75t_L g2056 ( 
.A(n_1994),
.Y(n_2056)
);

NAND2xp5_ASAP7_75t_L g2057 ( 
.A(n_1991),
.B(n_1030),
.Y(n_2057)
);

HB1xp67_ASAP7_75t_L g2058 ( 
.A(n_1956),
.Y(n_2058)
);

AOI22xp33_ASAP7_75t_SL g2059 ( 
.A1(n_1945),
.A2(n_1284),
.B1(n_503),
.B2(n_505),
.Y(n_2059)
);

BUFx2_ASAP7_75t_L g2060 ( 
.A(n_1961),
.Y(n_2060)
);

INVx2_ASAP7_75t_SL g2061 ( 
.A(n_2005),
.Y(n_2061)
);

INVx1_ASAP7_75t_L g2062 ( 
.A(n_1986),
.Y(n_2062)
);

INVx2_ASAP7_75t_L g2063 ( 
.A(n_1999),
.Y(n_2063)
);

BUFx6f_ASAP7_75t_L g2064 ( 
.A(n_1961),
.Y(n_2064)
);

OAI211xp5_ASAP7_75t_SL g2065 ( 
.A1(n_2010),
.A2(n_1032),
.B(n_1036),
.C(n_1031),
.Y(n_2065)
);

NAND2x1p5_ASAP7_75t_L g2066 ( 
.A(n_1952),
.B(n_1808),
.Y(n_2066)
);

INVx1_ASAP7_75t_SL g2067 ( 
.A(n_2040),
.Y(n_2067)
);

NAND2xp5_ASAP7_75t_L g2068 ( 
.A(n_2047),
.B(n_2021),
.Y(n_2068)
);

INVx4_ASAP7_75t_L g2069 ( 
.A(n_2034),
.Y(n_2069)
);

BUFx3_ASAP7_75t_L g2070 ( 
.A(n_2019),
.Y(n_2070)
);

INVx1_ASAP7_75t_L g2071 ( 
.A(n_2023),
.Y(n_2071)
);

INVx1_ASAP7_75t_L g2072 ( 
.A(n_2014),
.Y(n_2072)
);

INVx2_ASAP7_75t_L g2073 ( 
.A(n_2045),
.Y(n_2073)
);

INVx2_ASAP7_75t_L g2074 ( 
.A(n_2013),
.Y(n_2074)
);

INVx1_ASAP7_75t_L g2075 ( 
.A(n_2029),
.Y(n_2075)
);

CKINVDCx20_ASAP7_75t_R g2076 ( 
.A(n_2052),
.Y(n_2076)
);

INVx2_ASAP7_75t_L g2077 ( 
.A(n_2049),
.Y(n_2077)
);

INVx3_ASAP7_75t_L g2078 ( 
.A(n_2064),
.Y(n_2078)
);

NAND2xp5_ASAP7_75t_L g2079 ( 
.A(n_2024),
.B(n_1957),
.Y(n_2079)
);

INVx2_ASAP7_75t_SL g2080 ( 
.A(n_2064),
.Y(n_2080)
);

INVx1_ASAP7_75t_L g2081 ( 
.A(n_2020),
.Y(n_2081)
);

INVx2_ASAP7_75t_L g2082 ( 
.A(n_2051),
.Y(n_2082)
);

INVx2_ASAP7_75t_L g2083 ( 
.A(n_2016),
.Y(n_2083)
);

BUFx2_ASAP7_75t_L g2084 ( 
.A(n_2058),
.Y(n_2084)
);

AO31x2_ASAP7_75t_L g2085 ( 
.A1(n_2062),
.A2(n_1969),
.A3(n_1986),
.B(n_2007),
.Y(n_2085)
);

BUFx4f_ASAP7_75t_SL g2086 ( 
.A(n_2019),
.Y(n_2086)
);

INVx2_ASAP7_75t_L g2087 ( 
.A(n_2016),
.Y(n_2087)
);

INVx1_ASAP7_75t_L g2088 ( 
.A(n_2042),
.Y(n_2088)
);

INVx3_ASAP7_75t_L g2089 ( 
.A(n_2064),
.Y(n_2089)
);

AND2x2_ASAP7_75t_L g2090 ( 
.A(n_2040),
.B(n_1998),
.Y(n_2090)
);

INVx1_ASAP7_75t_L g2091 ( 
.A(n_2048),
.Y(n_2091)
);

INVx1_ASAP7_75t_L g2092 ( 
.A(n_2025),
.Y(n_2092)
);

NAND2x1p5_ASAP7_75t_L g2093 ( 
.A(n_2063),
.B(n_1964),
.Y(n_2093)
);

AO21x1_ASAP7_75t_L g2094 ( 
.A1(n_2053),
.A2(n_1986),
.B(n_1959),
.Y(n_2094)
);

INVx1_ASAP7_75t_L g2095 ( 
.A(n_2060),
.Y(n_2095)
);

INVx1_ASAP7_75t_SL g2096 ( 
.A(n_2022),
.Y(n_2096)
);

AO21x2_ASAP7_75t_L g2097 ( 
.A1(n_2054),
.A2(n_2002),
.B(n_1972),
.Y(n_2097)
);

INVx2_ASAP7_75t_L g2098 ( 
.A(n_2077),
.Y(n_2098)
);

NAND3xp33_ASAP7_75t_L g2099 ( 
.A(n_2084),
.B(n_2031),
.C(n_2017),
.Y(n_2099)
);

INVx1_ASAP7_75t_L g2100 ( 
.A(n_2071),
.Y(n_2100)
);

OR2x6_ASAP7_75t_L g2101 ( 
.A(n_2094),
.B(n_2066),
.Y(n_2101)
);

INVx2_ASAP7_75t_L g2102 ( 
.A(n_2083),
.Y(n_2102)
);

AND2x2_ASAP7_75t_L g2103 ( 
.A(n_2078),
.B(n_2089),
.Y(n_2103)
);

AOI22xp33_ASAP7_75t_L g2104 ( 
.A1(n_2094),
.A2(n_2053),
.B1(n_2055),
.B2(n_2096),
.Y(n_2104)
);

OAI22xp5_ASAP7_75t_L g2105 ( 
.A1(n_2096),
.A2(n_2054),
.B1(n_2059),
.B2(n_2056),
.Y(n_2105)
);

AND2x4_ASAP7_75t_L g2106 ( 
.A(n_2080),
.B(n_2078),
.Y(n_2106)
);

AOI22xp33_ASAP7_75t_L g2107 ( 
.A1(n_2092),
.A2(n_2026),
.B1(n_2065),
.B2(n_2036),
.Y(n_2107)
);

OAI22xp33_ASAP7_75t_L g2108 ( 
.A1(n_2067),
.A2(n_2057),
.B1(n_2015),
.B2(n_2032),
.Y(n_2108)
);

INVxp67_ASAP7_75t_L g2109 ( 
.A(n_2084),
.Y(n_2109)
);

AOI221xp5_ASAP7_75t_L g2110 ( 
.A1(n_2092),
.A2(n_2036),
.B1(n_2027),
.B2(n_2026),
.C(n_2018),
.Y(n_2110)
);

AOI221xp5_ASAP7_75t_L g2111 ( 
.A1(n_2090),
.A2(n_2018),
.B1(n_2043),
.B2(n_2033),
.C(n_1946),
.Y(n_2111)
);

BUFx2_ASAP7_75t_L g2112 ( 
.A(n_2078),
.Y(n_2112)
);

AND2x2_ASAP7_75t_L g2113 ( 
.A(n_2078),
.B(n_2038),
.Y(n_2113)
);

OAI211xp5_ASAP7_75t_L g2114 ( 
.A1(n_2090),
.A2(n_1941),
.B(n_1973),
.C(n_2044),
.Y(n_2114)
);

AND2x4_ASAP7_75t_L g2115 ( 
.A(n_2080),
.B(n_2061),
.Y(n_2115)
);

AOI222xp33_ASAP7_75t_L g2116 ( 
.A1(n_2086),
.A2(n_2035),
.B1(n_2033),
.B2(n_2044),
.C1(n_1044),
.C2(n_1038),
.Y(n_2116)
);

INVxp67_ASAP7_75t_SL g2117 ( 
.A(n_2077),
.Y(n_2117)
);

AO21x1_ASAP7_75t_L g2118 ( 
.A1(n_2068),
.A2(n_2088),
.B(n_2071),
.Y(n_2118)
);

AOI22xp33_ASAP7_75t_L g2119 ( 
.A1(n_2097),
.A2(n_2035),
.B1(n_2003),
.B2(n_1980),
.Y(n_2119)
);

AOI21xp5_ASAP7_75t_L g2120 ( 
.A1(n_2097),
.A2(n_1947),
.B(n_1950),
.Y(n_2120)
);

INVx3_ASAP7_75t_L g2121 ( 
.A(n_2089),
.Y(n_2121)
);

AOI222xp33_ASAP7_75t_L g2122 ( 
.A1(n_2070),
.A2(n_1040),
.B1(n_1037),
.B2(n_510),
.C1(n_506),
.C2(n_512),
.Y(n_2122)
);

INVx1_ASAP7_75t_L g2123 ( 
.A(n_2075),
.Y(n_2123)
);

INVx1_ASAP7_75t_L g2124 ( 
.A(n_2100),
.Y(n_2124)
);

INVx2_ASAP7_75t_L g2125 ( 
.A(n_2098),
.Y(n_2125)
);

BUFx2_ASAP7_75t_L g2126 ( 
.A(n_2109),
.Y(n_2126)
);

INVx1_ASAP7_75t_L g2127 ( 
.A(n_2123),
.Y(n_2127)
);

AND2x2_ASAP7_75t_L g2128 ( 
.A(n_2103),
.B(n_2112),
.Y(n_2128)
);

BUFx3_ASAP7_75t_L g2129 ( 
.A(n_2115),
.Y(n_2129)
);

AND2x2_ASAP7_75t_L g2130 ( 
.A(n_2121),
.B(n_2089),
.Y(n_2130)
);

INVx3_ASAP7_75t_L g2131 ( 
.A(n_2121),
.Y(n_2131)
);

NAND2xp5_ASAP7_75t_L g2132 ( 
.A(n_2109),
.B(n_2068),
.Y(n_2132)
);

AND2x2_ASAP7_75t_L g2133 ( 
.A(n_2106),
.B(n_2089),
.Y(n_2133)
);

INVx1_ASAP7_75t_L g2134 ( 
.A(n_2117),
.Y(n_2134)
);

AND2x2_ASAP7_75t_L g2135 ( 
.A(n_2106),
.B(n_2080),
.Y(n_2135)
);

NAND2xp5_ASAP7_75t_L g2136 ( 
.A(n_2118),
.B(n_2075),
.Y(n_2136)
);

NAND2x1p5_ASAP7_75t_L g2137 ( 
.A(n_2120),
.B(n_2067),
.Y(n_2137)
);

INVx6_ASAP7_75t_L g2138 ( 
.A(n_2101),
.Y(n_2138)
);

INVx2_ASAP7_75t_L g2139 ( 
.A(n_2098),
.Y(n_2139)
);

HB1xp67_ASAP7_75t_L g2140 ( 
.A(n_2117),
.Y(n_2140)
);

AND2x4_ASAP7_75t_SL g2141 ( 
.A(n_2115),
.B(n_2076),
.Y(n_2141)
);

AND2x2_ASAP7_75t_L g2142 ( 
.A(n_2101),
.B(n_2083),
.Y(n_2142)
);

INVx1_ASAP7_75t_L g2143 ( 
.A(n_2102),
.Y(n_2143)
);

AND2x2_ASAP7_75t_L g2144 ( 
.A(n_2101),
.B(n_2113),
.Y(n_2144)
);

INVx1_ASAP7_75t_L g2145 ( 
.A(n_2099),
.Y(n_2145)
);

INVx1_ASAP7_75t_L g2146 ( 
.A(n_2104),
.Y(n_2146)
);

INVx2_ASAP7_75t_L g2147 ( 
.A(n_2105),
.Y(n_2147)
);

OAI211xp5_ASAP7_75t_L g2148 ( 
.A1(n_2104),
.A2(n_2070),
.B(n_1954),
.C(n_2079),
.Y(n_2148)
);

INVx2_ASAP7_75t_L g2149 ( 
.A(n_2108),
.Y(n_2149)
);

INVx1_ASAP7_75t_L g2150 ( 
.A(n_2108),
.Y(n_2150)
);

OA21x2_ASAP7_75t_L g2151 ( 
.A1(n_2119),
.A2(n_2082),
.B(n_2077),
.Y(n_2151)
);

INVx1_ASAP7_75t_L g2152 ( 
.A(n_2114),
.Y(n_2152)
);

INVx2_ASAP7_75t_L g2153 ( 
.A(n_2119),
.Y(n_2153)
);

INVx2_ASAP7_75t_L g2154 ( 
.A(n_2111),
.Y(n_2154)
);

NAND2xp5_ASAP7_75t_SL g2155 ( 
.A(n_2107),
.B(n_2069),
.Y(n_2155)
);

AOI211xp5_ASAP7_75t_SL g2156 ( 
.A1(n_2148),
.A2(n_2110),
.B(n_1976),
.C(n_1996),
.Y(n_2156)
);

NAND2xp5_ASAP7_75t_L g2157 ( 
.A(n_2153),
.B(n_2107),
.Y(n_2157)
);

OAI33xp33_ASAP7_75t_L g2158 ( 
.A1(n_2145),
.A2(n_2079),
.A3(n_2088),
.B1(n_2082),
.B2(n_2072),
.B3(n_2081),
.Y(n_2158)
);

OAI22xp5_ASAP7_75t_L g2159 ( 
.A1(n_2149),
.A2(n_2070),
.B1(n_2095),
.B2(n_2069),
.Y(n_2159)
);

NAND2xp5_ASAP7_75t_L g2160 ( 
.A(n_2153),
.B(n_2091),
.Y(n_2160)
);

INVxp67_ASAP7_75t_L g2161 ( 
.A(n_2150),
.Y(n_2161)
);

AOI221xp5_ASAP7_75t_L g2162 ( 
.A1(n_2145),
.A2(n_2091),
.B1(n_2095),
.B2(n_2081),
.C(n_2072),
.Y(n_2162)
);

INVx2_ASAP7_75t_L g2163 ( 
.A(n_2129),
.Y(n_2163)
);

AOI22xp33_ASAP7_75t_L g2164 ( 
.A1(n_2154),
.A2(n_2122),
.B1(n_2097),
.B2(n_2116),
.Y(n_2164)
);

AOI22xp33_ASAP7_75t_L g2165 ( 
.A1(n_2154),
.A2(n_2097),
.B1(n_2069),
.B2(n_2039),
.Y(n_2165)
);

OAI321xp33_ASAP7_75t_L g2166 ( 
.A1(n_2148),
.A2(n_2093),
.A3(n_2073),
.B1(n_2082),
.B2(n_2041),
.C(n_2074),
.Y(n_2166)
);

AND2x2_ASAP7_75t_L g2167 ( 
.A(n_2141),
.B(n_2069),
.Y(n_2167)
);

AND2x2_ASAP7_75t_L g2168 ( 
.A(n_2141),
.B(n_2056),
.Y(n_2168)
);

AOI33xp33_ASAP7_75t_L g2169 ( 
.A1(n_2152),
.A2(n_1987),
.A3(n_2050),
.B1(n_2073),
.B2(n_2074),
.B3(n_2004),
.Y(n_2169)
);

BUFx2_ASAP7_75t_L g2170 ( 
.A(n_2129),
.Y(n_2170)
);

AOI221xp5_ASAP7_75t_L g2171 ( 
.A1(n_2153),
.A2(n_2074),
.B1(n_2073),
.B2(n_2087),
.C(n_2083),
.Y(n_2171)
);

OAI31xp33_ASAP7_75t_L g2172 ( 
.A1(n_2150),
.A2(n_2093),
.A3(n_2087),
.B(n_1997),
.Y(n_2172)
);

NAND2xp5_ASAP7_75t_L g2173 ( 
.A(n_2146),
.B(n_2087),
.Y(n_2173)
);

AOI221xp5_ASAP7_75t_L g2174 ( 
.A1(n_2152),
.A2(n_509),
.B1(n_510),
.B2(n_506),
.C(n_501),
.Y(n_2174)
);

OAI31xp33_ASAP7_75t_SL g2175 ( 
.A1(n_2155),
.A2(n_2028),
.A3(n_2037),
.B(n_2030),
.Y(n_2175)
);

OAI33xp33_ASAP7_75t_L g2176 ( 
.A1(n_2146),
.A2(n_2046),
.A3(n_517),
.B1(n_512),
.B2(n_520),
.B3(n_514),
.Y(n_2176)
);

OAI321xp33_ASAP7_75t_L g2177 ( 
.A1(n_2137),
.A2(n_2093),
.A3(n_2001),
.B1(n_2056),
.B2(n_1989),
.C(n_1983),
.Y(n_2177)
);

OR2x2_ASAP7_75t_L g2178 ( 
.A(n_2161),
.B(n_2149),
.Y(n_2178)
);

NAND2xp5_ASAP7_75t_L g2179 ( 
.A(n_2169),
.B(n_2154),
.Y(n_2179)
);

BUFx2_ASAP7_75t_L g2180 ( 
.A(n_2170),
.Y(n_2180)
);

INVx2_ASAP7_75t_L g2181 ( 
.A(n_2163),
.Y(n_2181)
);

AND2x4_ASAP7_75t_L g2182 ( 
.A(n_2167),
.B(n_2141),
.Y(n_2182)
);

INVx1_ASAP7_75t_L g2183 ( 
.A(n_2173),
.Y(n_2183)
);

INVx1_ASAP7_75t_L g2184 ( 
.A(n_2160),
.Y(n_2184)
);

INVx1_ASAP7_75t_L g2185 ( 
.A(n_2157),
.Y(n_2185)
);

AND2x2_ASAP7_75t_L g2186 ( 
.A(n_2168),
.B(n_2144),
.Y(n_2186)
);

INVx1_ASAP7_75t_L g2187 ( 
.A(n_2169),
.Y(n_2187)
);

AOI22xp33_ASAP7_75t_SL g2188 ( 
.A1(n_2159),
.A2(n_2149),
.B1(n_2147),
.B2(n_2138),
.Y(n_2188)
);

NOR2x1p5_ASAP7_75t_L g2189 ( 
.A(n_2175),
.B(n_2147),
.Y(n_2189)
);

NAND2xp5_ASAP7_75t_L g2190 ( 
.A(n_2164),
.B(n_2147),
.Y(n_2190)
);

INVx1_ASAP7_75t_L g2191 ( 
.A(n_2162),
.Y(n_2191)
);

INVx2_ASAP7_75t_L g2192 ( 
.A(n_2166),
.Y(n_2192)
);

INVx2_ASAP7_75t_L g2193 ( 
.A(n_2156),
.Y(n_2193)
);

INVx1_ASAP7_75t_L g2194 ( 
.A(n_2180),
.Y(n_2194)
);

AND2x2_ASAP7_75t_L g2195 ( 
.A(n_2182),
.B(n_2144),
.Y(n_2195)
);

OAI21xp5_ASAP7_75t_L g2196 ( 
.A1(n_2188),
.A2(n_2177),
.B(n_2164),
.Y(n_2196)
);

NOR2xp33_ASAP7_75t_R g2197 ( 
.A(n_2185),
.B(n_1284),
.Y(n_2197)
);

OAI221xp5_ASAP7_75t_SL g2198 ( 
.A1(n_2193),
.A2(n_2165),
.B1(n_2172),
.B2(n_2174),
.C(n_2126),
.Y(n_2198)
);

AOI221xp5_ASAP7_75t_L g2199 ( 
.A1(n_2191),
.A2(n_2165),
.B1(n_2158),
.B2(n_2126),
.C(n_2136),
.Y(n_2199)
);

NOR2xp33_ASAP7_75t_L g2200 ( 
.A(n_2182),
.B(n_1213),
.Y(n_2200)
);

NOR2xp33_ASAP7_75t_L g2201 ( 
.A(n_2182),
.B(n_1213),
.Y(n_2201)
);

AND2x2_ASAP7_75t_L g2202 ( 
.A(n_2186),
.B(n_2129),
.Y(n_2202)
);

NAND2xp5_ASAP7_75t_L g2203 ( 
.A(n_2194),
.B(n_2193),
.Y(n_2203)
);

AND2x2_ASAP7_75t_L g2204 ( 
.A(n_2195),
.B(n_2188),
.Y(n_2204)
);

AND2x4_ASAP7_75t_L g2205 ( 
.A(n_2202),
.B(n_2181),
.Y(n_2205)
);

BUFx3_ASAP7_75t_L g2206 ( 
.A(n_2200),
.Y(n_2206)
);

OR2x2_ASAP7_75t_L g2207 ( 
.A(n_2196),
.B(n_2178),
.Y(n_2207)
);

NAND2xp5_ASAP7_75t_L g2208 ( 
.A(n_2199),
.B(n_2187),
.Y(n_2208)
);

AND2x2_ASAP7_75t_L g2209 ( 
.A(n_2201),
.B(n_2189),
.Y(n_2209)
);

INVx1_ASAP7_75t_L g2210 ( 
.A(n_2203),
.Y(n_2210)
);

NAND2xp5_ASAP7_75t_SL g2211 ( 
.A(n_2205),
.B(n_2197),
.Y(n_2211)
);

INVx1_ASAP7_75t_L g2212 ( 
.A(n_2203),
.Y(n_2212)
);

AND2x2_ASAP7_75t_L g2213 ( 
.A(n_2204),
.B(n_2181),
.Y(n_2213)
);

AOI221xp5_ASAP7_75t_L g2214 ( 
.A1(n_2208),
.A2(n_2198),
.B1(n_2190),
.B2(n_2192),
.C(n_2179),
.Y(n_2214)
);

HB1xp67_ASAP7_75t_L g2215 ( 
.A(n_2213),
.Y(n_2215)
);

NAND2xp5_ASAP7_75t_L g2216 ( 
.A(n_2210),
.B(n_2205),
.Y(n_2216)
);

INVx1_ASAP7_75t_L g2217 ( 
.A(n_2212),
.Y(n_2217)
);

INVx2_ASAP7_75t_L g2218 ( 
.A(n_2215),
.Y(n_2218)
);

AND2x2_ASAP7_75t_L g2219 ( 
.A(n_2216),
.B(n_2209),
.Y(n_2219)
);

NOR2x1_ASAP7_75t_SL g2220 ( 
.A(n_2218),
.B(n_2211),
.Y(n_2220)
);

AND2x4_ASAP7_75t_L g2221 ( 
.A(n_2219),
.B(n_2206),
.Y(n_2221)
);

INVx1_ASAP7_75t_L g2222 ( 
.A(n_2218),
.Y(n_2222)
);

OR2x2_ASAP7_75t_L g2223 ( 
.A(n_2222),
.B(n_2207),
.Y(n_2223)
);

OAI21xp5_ASAP7_75t_L g2224 ( 
.A1(n_2221),
.A2(n_2214),
.B(n_2198),
.Y(n_2224)
);

AND2x2_ASAP7_75t_L g2225 ( 
.A(n_2223),
.B(n_2221),
.Y(n_2225)
);

INVx1_ASAP7_75t_L g2226 ( 
.A(n_2224),
.Y(n_2226)
);

OAI221xp5_ASAP7_75t_L g2227 ( 
.A1(n_2224),
.A2(n_2217),
.B1(n_2192),
.B2(n_2184),
.C(n_2183),
.Y(n_2227)
);

INVx1_ASAP7_75t_L g2228 ( 
.A(n_2225),
.Y(n_2228)
);

AOI21xp33_ASAP7_75t_SL g2229 ( 
.A1(n_2226),
.A2(n_2220),
.B(n_2137),
.Y(n_2229)
);

AO21x1_ASAP7_75t_L g2230 ( 
.A1(n_2227),
.A2(n_2137),
.B(n_2134),
.Y(n_2230)
);

XNOR2x1_ASAP7_75t_L g2231 ( 
.A(n_2225),
.B(n_8),
.Y(n_2231)
);

INVx1_ASAP7_75t_L g2232 ( 
.A(n_2228),
.Y(n_2232)
);

NAND3xp33_ASAP7_75t_L g2233 ( 
.A(n_2229),
.B(n_2140),
.C(n_2171),
.Y(n_2233)
);

INVx1_ASAP7_75t_L g2234 ( 
.A(n_2231),
.Y(n_2234)
);

OAI21xp33_ASAP7_75t_SL g2235 ( 
.A1(n_2230),
.A2(n_2136),
.B(n_2140),
.Y(n_2235)
);

AO22x2_ASAP7_75t_L g2236 ( 
.A1(n_2232),
.A2(n_2134),
.B1(n_2131),
.B2(n_2125),
.Y(n_2236)
);

OA22x2_ASAP7_75t_L g2237 ( 
.A1(n_2234),
.A2(n_2131),
.B1(n_2132),
.B2(n_2142),
.Y(n_2237)
);

OAI221xp5_ASAP7_75t_L g2238 ( 
.A1(n_2235),
.A2(n_2138),
.B1(n_2137),
.B2(n_2151),
.C(n_2132),
.Y(n_2238)
);

NAND2x1_ASAP7_75t_L g2239 ( 
.A(n_2233),
.B(n_2138),
.Y(n_2239)
);

AOI21xp33_ASAP7_75t_SL g2240 ( 
.A1(n_2232),
.A2(n_9),
.B(n_10),
.Y(n_2240)
);

INVx1_ASAP7_75t_SL g2241 ( 
.A(n_2232),
.Y(n_2241)
);

NAND3x1_ASAP7_75t_SL g2242 ( 
.A(n_2235),
.B(n_2138),
.C(n_2142),
.Y(n_2242)
);

INVx1_ASAP7_75t_L g2243 ( 
.A(n_2232),
.Y(n_2243)
);

AOI22xp5_ASAP7_75t_L g2244 ( 
.A1(n_2232),
.A2(n_2138),
.B1(n_2176),
.B2(n_2142),
.Y(n_2244)
);

INVx1_ASAP7_75t_L g2245 ( 
.A(n_2232),
.Y(n_2245)
);

AOI221xp5_ASAP7_75t_L g2246 ( 
.A1(n_2235),
.A2(n_2131),
.B1(n_2127),
.B2(n_2124),
.C(n_2143),
.Y(n_2246)
);

NAND3xp33_ASAP7_75t_L g2247 ( 
.A(n_2232),
.B(n_2151),
.C(n_514),
.Y(n_2247)
);

HB1xp67_ASAP7_75t_L g2248 ( 
.A(n_2235),
.Y(n_2248)
);

NAND2xp5_ASAP7_75t_L g2249 ( 
.A(n_2232),
.B(n_2131),
.Y(n_2249)
);

XNOR2x1_ASAP7_75t_L g2250 ( 
.A(n_2241),
.B(n_9),
.Y(n_2250)
);

NAND3xp33_ASAP7_75t_L g2251 ( 
.A(n_2248),
.B(n_1636),
.C(n_1610),
.Y(n_2251)
);

AND2x2_ASAP7_75t_L g2252 ( 
.A(n_2243),
.B(n_2128),
.Y(n_2252)
);

O2A1O1Ixp33_ASAP7_75t_L g2253 ( 
.A1(n_2240),
.A2(n_1636),
.B(n_2151),
.C(n_14),
.Y(n_2253)
);

NAND3xp33_ASAP7_75t_L g2254 ( 
.A(n_2245),
.B(n_517),
.C(n_509),
.Y(n_2254)
);

NOR3xp33_ASAP7_75t_L g2255 ( 
.A(n_2242),
.B(n_2249),
.C(n_2239),
.Y(n_2255)
);

NOR2xp33_ASAP7_75t_L g2256 ( 
.A(n_2238),
.B(n_2237),
.Y(n_2256)
);

O2A1O1Ixp33_ASAP7_75t_SL g2257 ( 
.A1(n_2247),
.A2(n_2125),
.B(n_2139),
.C(n_2127),
.Y(n_2257)
);

NAND2xp5_ASAP7_75t_SL g2258 ( 
.A(n_2244),
.B(n_2125),
.Y(n_2258)
);

NAND3xp33_ASAP7_75t_L g2259 ( 
.A(n_2246),
.B(n_2236),
.C(n_530),
.Y(n_2259)
);

NAND3xp33_ASAP7_75t_SL g2260 ( 
.A(n_2241),
.B(n_530),
.C(n_520),
.Y(n_2260)
);

NOR2x1_ASAP7_75t_L g2261 ( 
.A(n_2243),
.B(n_1681),
.Y(n_2261)
);

NAND2xp5_ASAP7_75t_L g2262 ( 
.A(n_2240),
.B(n_2151),
.Y(n_2262)
);

INVx1_ASAP7_75t_L g2263 ( 
.A(n_2242),
.Y(n_2263)
);

OR2x2_ASAP7_75t_L g2264 ( 
.A(n_2249),
.B(n_2151),
.Y(n_2264)
);

NAND3xp33_ASAP7_75t_L g2265 ( 
.A(n_2248),
.B(n_533),
.C(n_531),
.Y(n_2265)
);

NAND4xp25_ASAP7_75t_L g2266 ( 
.A(n_2241),
.B(n_14),
.C(n_11),
.D(n_12),
.Y(n_2266)
);

NOR3x1_ASAP7_75t_L g2267 ( 
.A(n_2249),
.B(n_2124),
.C(n_2143),
.Y(n_2267)
);

OAI211xp5_ASAP7_75t_L g2268 ( 
.A1(n_2248),
.A2(n_533),
.B(n_535),
.C(n_531),
.Y(n_2268)
);

NOR3xp33_ASAP7_75t_L g2269 ( 
.A(n_2243),
.B(n_537),
.C(n_535),
.Y(n_2269)
);

NAND3xp33_ASAP7_75t_L g2270 ( 
.A(n_2248),
.B(n_640),
.C(n_537),
.Y(n_2270)
);

AND2x2_ASAP7_75t_L g2271 ( 
.A(n_2241),
.B(n_2128),
.Y(n_2271)
);

AOI211xp5_ASAP7_75t_L g2272 ( 
.A1(n_2241),
.A2(n_642),
.B(n_645),
.C(n_640),
.Y(n_2272)
);

OAI322xp33_ASAP7_75t_L g2273 ( 
.A1(n_2239),
.A2(n_2139),
.A3(n_2135),
.B1(n_2130),
.B2(n_2133),
.C1(n_17),
.C2(n_20),
.Y(n_2273)
);

NOR2x1_ASAP7_75t_L g2274 ( 
.A(n_2243),
.B(n_11),
.Y(n_2274)
);

NOR3xp33_ASAP7_75t_SL g2275 ( 
.A(n_2243),
.B(n_645),
.C(n_642),
.Y(n_2275)
);

AND2x4_ASAP7_75t_L g2276 ( 
.A(n_2243),
.B(n_2133),
.Y(n_2276)
);

NOR2xp33_ASAP7_75t_L g2277 ( 
.A(n_2241),
.B(n_2139),
.Y(n_2277)
);

NOR2x1_ASAP7_75t_L g2278 ( 
.A(n_2243),
.B(n_15),
.Y(n_2278)
);

AND2x2_ASAP7_75t_L g2279 ( 
.A(n_2241),
.B(n_2135),
.Y(n_2279)
);

NOR2xp33_ASAP7_75t_R g2280 ( 
.A(n_2243),
.B(n_18),
.Y(n_2280)
);

NAND4xp25_ASAP7_75t_L g2281 ( 
.A(n_2241),
.B(n_23),
.C(n_19),
.D(n_21),
.Y(n_2281)
);

NOR2x1_ASAP7_75t_L g2282 ( 
.A(n_2243),
.B(n_19),
.Y(n_2282)
);

INVx1_ASAP7_75t_L g2283 ( 
.A(n_2242),
.Y(n_2283)
);

NOR4xp25_ASAP7_75t_L g2284 ( 
.A(n_2241),
.B(n_2130),
.C(n_24),
.D(n_21),
.Y(n_2284)
);

NOR3xp33_ASAP7_75t_SL g2285 ( 
.A(n_2243),
.B(n_777),
.C(n_776),
.Y(n_2285)
);

NAND3xp33_ASAP7_75t_L g2286 ( 
.A(n_2248),
.B(n_777),
.C(n_776),
.Y(n_2286)
);

NOR2x1_ASAP7_75t_L g2287 ( 
.A(n_2243),
.B(n_23),
.Y(n_2287)
);

AND4x2_ASAP7_75t_L g2288 ( 
.A(n_2246),
.B(n_29),
.C(n_24),
.D(n_25),
.Y(n_2288)
);

NOR3xp33_ASAP7_75t_SL g2289 ( 
.A(n_2243),
.B(n_780),
.C(n_779),
.Y(n_2289)
);

NAND3xp33_ASAP7_75t_L g2290 ( 
.A(n_2248),
.B(n_780),
.C(n_779),
.Y(n_2290)
);

NOR3xp33_ASAP7_75t_L g2291 ( 
.A(n_2243),
.B(n_789),
.C(n_783),
.Y(n_2291)
);

AND2x2_ASAP7_75t_L g2292 ( 
.A(n_2241),
.B(n_2008),
.Y(n_2292)
);

NAND4xp25_ASAP7_75t_L g2293 ( 
.A(n_2241),
.B(n_32),
.C(n_30),
.D(n_31),
.Y(n_2293)
);

NAND3x1_ASAP7_75t_SL g2294 ( 
.A(n_2240),
.B(n_30),
.C(n_31),
.Y(n_2294)
);

NOR2x1_ASAP7_75t_L g2295 ( 
.A(n_2243),
.B(n_32),
.Y(n_2295)
);

AND2x2_ASAP7_75t_L g2296 ( 
.A(n_2279),
.B(n_2008),
.Y(n_2296)
);

AOI22xp33_ASAP7_75t_L g2297 ( 
.A1(n_2276),
.A2(n_789),
.B1(n_793),
.B2(n_783),
.Y(n_2297)
);

OA21x2_ASAP7_75t_L g2298 ( 
.A1(n_2263),
.A2(n_796),
.B(n_793),
.Y(n_2298)
);

INVx1_ASAP7_75t_L g2299 ( 
.A(n_2271),
.Y(n_2299)
);

INVx1_ASAP7_75t_L g2300 ( 
.A(n_2252),
.Y(n_2300)
);

OAI22xp33_ASAP7_75t_L g2301 ( 
.A1(n_2283),
.A2(n_1808),
.B1(n_800),
.B2(n_808),
.Y(n_2301)
);

AND2x2_ASAP7_75t_L g2302 ( 
.A(n_2276),
.B(n_2085),
.Y(n_2302)
);

OAI311xp33_ASAP7_75t_L g2303 ( 
.A1(n_2262),
.A2(n_35),
.A3(n_33),
.B1(n_34),
.C1(n_37),
.Y(n_2303)
);

AOI211xp5_ASAP7_75t_L g2304 ( 
.A1(n_2284),
.A2(n_800),
.B(n_808),
.C(n_796),
.Y(n_2304)
);

AND2x4_ASAP7_75t_L g2305 ( 
.A(n_2274),
.B(n_2006),
.Y(n_2305)
);

OAI22xp33_ASAP7_75t_L g2306 ( 
.A1(n_2266),
.A2(n_816),
.B1(n_819),
.B2(n_814),
.Y(n_2306)
);

INVx1_ASAP7_75t_L g2307 ( 
.A(n_2278),
.Y(n_2307)
);

NAND4xp25_ASAP7_75t_L g2308 ( 
.A(n_2255),
.B(n_2256),
.C(n_2277),
.D(n_2251),
.Y(n_2308)
);

AOI22xp5_ASAP7_75t_L g2309 ( 
.A1(n_2250),
.A2(n_816),
.B1(n_819),
.B2(n_814),
.Y(n_2309)
);

INVx1_ASAP7_75t_L g2310 ( 
.A(n_2282),
.Y(n_2310)
);

OAI221xp5_ASAP7_75t_L g2311 ( 
.A1(n_2287),
.A2(n_677),
.B1(n_679),
.B2(n_675),
.C(n_671),
.Y(n_2311)
);

OAI21xp5_ASAP7_75t_L g2312 ( 
.A1(n_2295),
.A2(n_684),
.B(n_682),
.Y(n_2312)
);

OAI221xp5_ASAP7_75t_L g2313 ( 
.A1(n_2253),
.A2(n_703),
.B1(n_717),
.B2(n_699),
.C(n_685),
.Y(n_2313)
);

HB1xp67_ASAP7_75t_L g2314 ( 
.A(n_2280),
.Y(n_2314)
);

AOI22xp33_ASAP7_75t_L g2315 ( 
.A1(n_2273),
.A2(n_723),
.B1(n_728),
.B2(n_720),
.Y(n_2315)
);

AOI22xp33_ASAP7_75t_L g2316 ( 
.A1(n_2292),
.A2(n_748),
.B1(n_750),
.B2(n_734),
.Y(n_2316)
);

AOI221xp5_ASAP7_75t_L g2317 ( 
.A1(n_2257),
.A2(n_757),
.B1(n_769),
.B2(n_752),
.C(n_751),
.Y(n_2317)
);

AND2x2_ASAP7_75t_L g2318 ( 
.A(n_2267),
.B(n_2085),
.Y(n_2318)
);

OAI21xp5_ASAP7_75t_SL g2319 ( 
.A1(n_2268),
.A2(n_34),
.B(n_38),
.Y(n_2319)
);

O2A1O1Ixp5_ASAP7_75t_L g2320 ( 
.A1(n_2258),
.A2(n_43),
.B(n_39),
.C(n_42),
.Y(n_2320)
);

INVx2_ASAP7_75t_L g2321 ( 
.A(n_2264),
.Y(n_2321)
);

AOI221xp5_ASAP7_75t_L g2322 ( 
.A1(n_2265),
.A2(n_774),
.B1(n_772),
.B2(n_771),
.C(n_46),
.Y(n_2322)
);

OAI211xp5_ASAP7_75t_L g2323 ( 
.A1(n_2281),
.A2(n_46),
.B(n_43),
.C(n_45),
.Y(n_2323)
);

OR2x2_ASAP7_75t_L g2324 ( 
.A(n_2293),
.B(n_47),
.Y(n_2324)
);

INVxp33_ASAP7_75t_SL g2325 ( 
.A(n_2270),
.Y(n_2325)
);

INVx1_ASAP7_75t_SL g2326 ( 
.A(n_2261),
.Y(n_2326)
);

INVx1_ASAP7_75t_L g2327 ( 
.A(n_2294),
.Y(n_2327)
);

NAND2xp5_ASAP7_75t_L g2328 ( 
.A(n_2275),
.B(n_48),
.Y(n_2328)
);

AOI22xp33_ASAP7_75t_SL g2329 ( 
.A1(n_2286),
.A2(n_1682),
.B1(n_50),
.B2(n_48),
.Y(n_2329)
);

AO22x2_ASAP7_75t_L g2330 ( 
.A1(n_2290),
.A2(n_57),
.B1(n_49),
.B2(n_52),
.Y(n_2330)
);

NAND4xp75_ASAP7_75t_L g2331 ( 
.A(n_2285),
.B(n_60),
.C(n_52),
.D(n_58),
.Y(n_2331)
);

OAI21xp5_ASAP7_75t_L g2332 ( 
.A1(n_2259),
.A2(n_1586),
.B(n_1682),
.Y(n_2332)
);

XNOR2xp5_ASAP7_75t_L g2333 ( 
.A(n_2289),
.B(n_60),
.Y(n_2333)
);

NAND2xp5_ASAP7_75t_L g2334 ( 
.A(n_2272),
.B(n_62),
.Y(n_2334)
);

INVxp33_ASAP7_75t_L g2335 ( 
.A(n_2269),
.Y(n_2335)
);

AND2x2_ASAP7_75t_L g2336 ( 
.A(n_2291),
.B(n_2254),
.Y(n_2336)
);

A2O1A1Ixp33_ASAP7_75t_L g2337 ( 
.A1(n_2260),
.A2(n_66),
.B(n_63),
.C(n_65),
.Y(n_2337)
);

AOI211xp5_ASAP7_75t_SL g2338 ( 
.A1(n_2288),
.A2(n_67),
.B(n_63),
.C(n_65),
.Y(n_2338)
);

AOI211xp5_ASAP7_75t_L g2339 ( 
.A1(n_2284),
.A2(n_70),
.B(n_68),
.C(n_69),
.Y(n_2339)
);

OR2x2_ASAP7_75t_L g2340 ( 
.A(n_2284),
.B(n_69),
.Y(n_2340)
);

NOR3xp33_ASAP7_75t_L g2341 ( 
.A(n_2263),
.B(n_1235),
.C(n_1224),
.Y(n_2341)
);

NOR3xp33_ASAP7_75t_L g2342 ( 
.A(n_2263),
.B(n_1235),
.C(n_1224),
.Y(n_2342)
);

OAI22xp5_ASAP7_75t_L g2343 ( 
.A1(n_2263),
.A2(n_2093),
.B1(n_1586),
.B2(n_2037),
.Y(n_2343)
);

OAI211xp5_ASAP7_75t_L g2344 ( 
.A1(n_2284),
.A2(n_74),
.B(n_71),
.C(n_73),
.Y(n_2344)
);

NAND4xp25_ASAP7_75t_L g2345 ( 
.A(n_2255),
.B(n_74),
.C(n_71),
.D(n_73),
.Y(n_2345)
);

OAI22xp5_ASAP7_75t_L g2346 ( 
.A1(n_2263),
.A2(n_2030),
.B1(n_2000),
.B2(n_1227),
.Y(n_2346)
);

INVxp67_ASAP7_75t_L g2347 ( 
.A(n_2274),
.Y(n_2347)
);

OAI221xp5_ASAP7_75t_L g2348 ( 
.A1(n_2284),
.A2(n_78),
.B1(n_76),
.B2(n_77),
.C(n_79),
.Y(n_2348)
);

NOR2xp33_ASAP7_75t_L g2349 ( 
.A(n_2273),
.B(n_78),
.Y(n_2349)
);

NOR3xp33_ASAP7_75t_L g2350 ( 
.A(n_2263),
.B(n_1235),
.C(n_1224),
.Y(n_2350)
);

NOR2x1_ASAP7_75t_L g2351 ( 
.A(n_2274),
.B(n_80),
.Y(n_2351)
);

OAI311xp33_ASAP7_75t_L g2352 ( 
.A1(n_2263),
.A2(n_83),
.A3(n_81),
.B1(n_82),
.C1(n_86),
.Y(n_2352)
);

AOI211xp5_ASAP7_75t_L g2353 ( 
.A1(n_2284),
.A2(n_87),
.B(n_82),
.C(n_86),
.Y(n_2353)
);

NAND4xp25_ASAP7_75t_SL g2354 ( 
.A(n_2253),
.B(n_90),
.C(n_87),
.D(n_89),
.Y(n_2354)
);

AOI22xp5_ASAP7_75t_L g2355 ( 
.A1(n_2276),
.A2(n_1599),
.B1(n_1612),
.B2(n_1598),
.Y(n_2355)
);

NOR2xp67_ASAP7_75t_L g2356 ( 
.A(n_2266),
.B(n_89),
.Y(n_2356)
);

NAND4xp25_ASAP7_75t_L g2357 ( 
.A(n_2255),
.B(n_93),
.C(n_91),
.D(n_92),
.Y(n_2357)
);

NAND4xp75_ASAP7_75t_L g2358 ( 
.A(n_2274),
.B(n_94),
.C(n_91),
.D(n_93),
.Y(n_2358)
);

AOI22xp5_ASAP7_75t_L g2359 ( 
.A1(n_2276),
.A2(n_1599),
.B1(n_1612),
.B2(n_1598),
.Y(n_2359)
);

AOI221xp5_ASAP7_75t_L g2360 ( 
.A1(n_2284),
.A2(n_98),
.B1(n_95),
.B2(n_97),
.C(n_99),
.Y(n_2360)
);

INVx1_ASAP7_75t_L g2361 ( 
.A(n_2279),
.Y(n_2361)
);

NAND3xp33_ASAP7_75t_L g2362 ( 
.A(n_2255),
.B(n_98),
.C(n_101),
.Y(n_2362)
);

AOI21xp5_ASAP7_75t_L g2363 ( 
.A1(n_2263),
.A2(n_1227),
.B(n_1222),
.Y(n_2363)
);

OAI322xp33_ASAP7_75t_L g2364 ( 
.A1(n_2263),
.A2(n_101),
.A3(n_102),
.B1(n_103),
.B2(n_104),
.C1(n_105),
.C2(n_106),
.Y(n_2364)
);

AOI211xp5_ASAP7_75t_L g2365 ( 
.A1(n_2284),
.A2(n_107),
.B(n_103),
.C(n_106),
.Y(n_2365)
);

INVx1_ASAP7_75t_L g2366 ( 
.A(n_2279),
.Y(n_2366)
);

NAND2xp5_ASAP7_75t_L g2367 ( 
.A(n_2276),
.B(n_108),
.Y(n_2367)
);

INVx1_ASAP7_75t_L g2368 ( 
.A(n_2279),
.Y(n_2368)
);

AOI22x1_ASAP7_75t_L g2369 ( 
.A1(n_2263),
.A2(n_112),
.B1(n_109),
.B2(n_111),
.Y(n_2369)
);

AOI322xp5_ASAP7_75t_L g2370 ( 
.A1(n_2271),
.A2(n_112),
.A3(n_113),
.B1(n_114),
.B2(n_116),
.C1(n_117),
.C2(n_118),
.Y(n_2370)
);

AND2x2_ASAP7_75t_L g2371 ( 
.A(n_2279),
.B(n_2085),
.Y(n_2371)
);

AOI22x1_ASAP7_75t_L g2372 ( 
.A1(n_2263),
.A2(n_117),
.B1(n_113),
.B2(n_114),
.Y(n_2372)
);

OAI21xp33_ASAP7_75t_L g2373 ( 
.A1(n_2271),
.A2(n_1240),
.B(n_1222),
.Y(n_2373)
);

NAND3xp33_ASAP7_75t_SL g2374 ( 
.A(n_2255),
.B(n_118),
.C(n_120),
.Y(n_2374)
);

INVx1_ASAP7_75t_L g2375 ( 
.A(n_2279),
.Y(n_2375)
);

AOI22xp5_ASAP7_75t_L g2376 ( 
.A1(n_2276),
.A2(n_1612),
.B1(n_1652),
.B2(n_1599),
.Y(n_2376)
);

OAI31xp33_ASAP7_75t_SL g2377 ( 
.A1(n_2271),
.A2(n_122),
.A3(n_120),
.B(n_121),
.Y(n_2377)
);

NAND2xp5_ASAP7_75t_L g2378 ( 
.A(n_2377),
.B(n_2351),
.Y(n_2378)
);

NAND3x1_ASAP7_75t_L g2379 ( 
.A(n_2327),
.B(n_121),
.C(n_127),
.Y(n_2379)
);

NAND3xp33_ASAP7_75t_SL g2380 ( 
.A(n_2339),
.B(n_127),
.C(n_128),
.Y(n_2380)
);

NAND3xp33_ASAP7_75t_SL g2381 ( 
.A(n_2353),
.B(n_2365),
.C(n_2360),
.Y(n_2381)
);

NAND4xp75_ASAP7_75t_L g2382 ( 
.A(n_2299),
.B(n_131),
.C(n_129),
.D(n_130),
.Y(n_2382)
);

OAI211xp5_ASAP7_75t_L g2383 ( 
.A1(n_2345),
.A2(n_133),
.B(n_131),
.C(n_132),
.Y(n_2383)
);

NAND3xp33_ASAP7_75t_L g2384 ( 
.A(n_2362),
.B(n_2357),
.C(n_2349),
.Y(n_2384)
);

NOR4xp25_ASAP7_75t_L g2385 ( 
.A(n_2303),
.B(n_134),
.C(n_132),
.D(n_133),
.Y(n_2385)
);

NAND2xp5_ASAP7_75t_L g2386 ( 
.A(n_2361),
.B(n_134),
.Y(n_2386)
);

NAND2xp5_ASAP7_75t_L g2387 ( 
.A(n_2366),
.B(n_136),
.Y(n_2387)
);

AND2x4_ASAP7_75t_L g2388 ( 
.A(n_2307),
.B(n_2310),
.Y(n_2388)
);

INVx1_ASAP7_75t_L g2389 ( 
.A(n_2340),
.Y(n_2389)
);

INVx1_ASAP7_75t_L g2390 ( 
.A(n_2367),
.Y(n_2390)
);

INVx1_ASAP7_75t_L g2391 ( 
.A(n_2358),
.Y(n_2391)
);

AND2x4_ASAP7_75t_L g2392 ( 
.A(n_2347),
.B(n_2006),
.Y(n_2392)
);

NAND3xp33_ASAP7_75t_L g2393 ( 
.A(n_2369),
.B(n_139),
.C(n_140),
.Y(n_2393)
);

AND3x2_ASAP7_75t_L g2394 ( 
.A(n_2304),
.B(n_139),
.C(n_141),
.Y(n_2394)
);

AND2x4_ASAP7_75t_L g2395 ( 
.A(n_2368),
.B(n_142),
.Y(n_2395)
);

NAND2x1p5_ASAP7_75t_L g2396 ( 
.A(n_2300),
.B(n_2375),
.Y(n_2396)
);

OAI221xp5_ASAP7_75t_L g2397 ( 
.A1(n_2348),
.A2(n_143),
.B1(n_144),
.B2(n_146),
.C(n_147),
.Y(n_2397)
);

NOR2x1_ASAP7_75t_L g2398 ( 
.A(n_2374),
.B(n_146),
.Y(n_2398)
);

INVx1_ASAP7_75t_SL g2399 ( 
.A(n_2324),
.Y(n_2399)
);

OR2x2_ASAP7_75t_L g2400 ( 
.A(n_2344),
.B(n_149),
.Y(n_2400)
);

NOR4xp25_ASAP7_75t_SL g2401 ( 
.A(n_2311),
.B(n_152),
.C(n_150),
.D(n_151),
.Y(n_2401)
);

AND2x2_ASAP7_75t_L g2402 ( 
.A(n_2338),
.B(n_2085),
.Y(n_2402)
);

NOR3xp33_ASAP7_75t_L g2403 ( 
.A(n_2308),
.B(n_1278),
.C(n_1245),
.Y(n_2403)
);

NAND4xp75_ASAP7_75t_L g2404 ( 
.A(n_2356),
.B(n_156),
.C(n_150),
.D(n_154),
.Y(n_2404)
);

NOR4xp75_ASAP7_75t_SL g2405 ( 
.A(n_2328),
.B(n_158),
.C(n_154),
.D(n_157),
.Y(n_2405)
);

AOI22xp5_ASAP7_75t_L g2406 ( 
.A1(n_2323),
.A2(n_1692),
.B1(n_1652),
.B2(n_1278),
.Y(n_2406)
);

OR2x2_ASAP7_75t_SL g2407 ( 
.A(n_2314),
.B(n_157),
.Y(n_2407)
);

AND2x4_ASAP7_75t_L g2408 ( 
.A(n_2296),
.B(n_2321),
.Y(n_2408)
);

AND2x2_ASAP7_75t_L g2409 ( 
.A(n_2371),
.B(n_2085),
.Y(n_2409)
);

NOR4xp25_ASAP7_75t_L g2410 ( 
.A(n_2315),
.B(n_161),
.C(n_158),
.D(n_160),
.Y(n_2410)
);

INVx1_ASAP7_75t_L g2411 ( 
.A(n_2333),
.Y(n_2411)
);

HB1xp67_ASAP7_75t_L g2412 ( 
.A(n_2372),
.Y(n_2412)
);

NOR2x1_ASAP7_75t_L g2413 ( 
.A(n_2364),
.B(n_2331),
.Y(n_2413)
);

INVxp33_ASAP7_75t_SL g2414 ( 
.A(n_2309),
.Y(n_2414)
);

HB1xp67_ASAP7_75t_L g2415 ( 
.A(n_2354),
.Y(n_2415)
);

AND2x2_ASAP7_75t_L g2416 ( 
.A(n_2302),
.B(n_2085),
.Y(n_2416)
);

NOR3xp33_ASAP7_75t_L g2417 ( 
.A(n_2334),
.B(n_1278),
.C(n_1245),
.Y(n_2417)
);

AND2x4_ASAP7_75t_L g2418 ( 
.A(n_2326),
.B(n_162),
.Y(n_2418)
);

NAND2x1_ASAP7_75t_L g2419 ( 
.A(n_2298),
.B(n_1652),
.Y(n_2419)
);

NOR2xp33_ASAP7_75t_L g2420 ( 
.A(n_2319),
.B(n_163),
.Y(n_2420)
);

AOI222xp33_ASAP7_75t_L g2421 ( 
.A1(n_2318),
.A2(n_2343),
.B1(n_2313),
.B2(n_2306),
.C1(n_2312),
.C2(n_2322),
.Y(n_2421)
);

NAND2xp5_ASAP7_75t_SL g2422 ( 
.A(n_2320),
.B(n_1245),
.Y(n_2422)
);

AND2x2_ASAP7_75t_SL g2423 ( 
.A(n_2298),
.B(n_163),
.Y(n_2423)
);

OR2x2_ASAP7_75t_L g2424 ( 
.A(n_2337),
.B(n_164),
.Y(n_2424)
);

NOR3xp33_ASAP7_75t_SL g2425 ( 
.A(n_2301),
.B(n_166),
.C(n_168),
.Y(n_2425)
);

INVxp33_ASAP7_75t_L g2426 ( 
.A(n_2330),
.Y(n_2426)
);

NAND2xp5_ASAP7_75t_L g2427 ( 
.A(n_2329),
.B(n_2370),
.Y(n_2427)
);

AND2x4_ASAP7_75t_L g2428 ( 
.A(n_2336),
.B(n_169),
.Y(n_2428)
);

AOI211xp5_ASAP7_75t_L g2429 ( 
.A1(n_2352),
.A2(n_172),
.B(n_169),
.C(n_170),
.Y(n_2429)
);

NAND2xp5_ASAP7_75t_L g2430 ( 
.A(n_2305),
.B(n_172),
.Y(n_2430)
);

NAND3xp33_ASAP7_75t_L g2431 ( 
.A(n_2316),
.B(n_173),
.C(n_1240),
.Y(n_2431)
);

NAND4xp75_ASAP7_75t_L g2432 ( 
.A(n_2363),
.B(n_173),
.C(n_1249),
.D(n_1241),
.Y(n_2432)
);

OAI221xp5_ASAP7_75t_L g2433 ( 
.A1(n_2332),
.A2(n_1330),
.B1(n_1633),
.B2(n_1251),
.C(n_1266),
.Y(n_2433)
);

NOR4xp75_ASAP7_75t_L g2434 ( 
.A(n_2373),
.B(n_180),
.C(n_176),
.D(n_177),
.Y(n_2434)
);

AND2x2_ASAP7_75t_L g2435 ( 
.A(n_2330),
.B(n_2085),
.Y(n_2435)
);

AOI211xp5_ASAP7_75t_L g2436 ( 
.A1(n_2335),
.A2(n_1241),
.B(n_1251),
.C(n_1249),
.Y(n_2436)
);

OAI22xp33_ASAP7_75t_L g2437 ( 
.A1(n_2355),
.A2(n_1692),
.B1(n_1767),
.B2(n_1766),
.Y(n_2437)
);

HB1xp67_ASAP7_75t_L g2438 ( 
.A(n_2305),
.Y(n_2438)
);

NAND2xp5_ASAP7_75t_L g2439 ( 
.A(n_2325),
.B(n_1253),
.Y(n_2439)
);

AND3x4_ASAP7_75t_L g2440 ( 
.A(n_2341),
.B(n_1696),
.C(n_1693),
.Y(n_2440)
);

INVx1_ASAP7_75t_L g2441 ( 
.A(n_2342),
.Y(n_2441)
);

NAND3xp33_ASAP7_75t_L g2442 ( 
.A(n_2317),
.B(n_1257),
.C(n_1253),
.Y(n_2442)
);

AND3x4_ASAP7_75t_L g2443 ( 
.A(n_2350),
.B(n_1696),
.C(n_1693),
.Y(n_2443)
);

INVx1_ASAP7_75t_L g2444 ( 
.A(n_2346),
.Y(n_2444)
);

NAND3xp33_ASAP7_75t_SL g2445 ( 
.A(n_2385),
.B(n_2297),
.C(n_2376),
.Y(n_2445)
);

OAI22xp5_ASAP7_75t_L g2446 ( 
.A1(n_2429),
.A2(n_2396),
.B1(n_2397),
.B2(n_2393),
.Y(n_2446)
);

INVx2_ASAP7_75t_L g2447 ( 
.A(n_2428),
.Y(n_2447)
);

NAND3xp33_ASAP7_75t_SL g2448 ( 
.A(n_2378),
.B(n_2401),
.C(n_2426),
.Y(n_2448)
);

NAND3xp33_ASAP7_75t_SL g2449 ( 
.A(n_2391),
.B(n_2359),
.C(n_1330),
.Y(n_2449)
);

NOR2xp33_ASAP7_75t_SL g2450 ( 
.A(n_2404),
.B(n_1257),
.Y(n_2450)
);

NAND5xp2_ASAP7_75t_L g2451 ( 
.A(n_2411),
.B(n_1687),
.C(n_189),
.D(n_190),
.E(n_192),
.Y(n_2451)
);

OAI221xp5_ASAP7_75t_L g2452 ( 
.A1(n_2383),
.A2(n_1274),
.B1(n_1272),
.B2(n_1271),
.C(n_1266),
.Y(n_2452)
);

OAI21xp5_ASAP7_75t_L g2453 ( 
.A1(n_2420),
.A2(n_1272),
.B(n_1271),
.Y(n_2453)
);

NAND3xp33_ASAP7_75t_L g2454 ( 
.A(n_2384),
.B(n_1276),
.C(n_1274),
.Y(n_2454)
);

INVx1_ASAP7_75t_L g2455 ( 
.A(n_2395),
.Y(n_2455)
);

NAND2xp5_ASAP7_75t_L g2456 ( 
.A(n_2418),
.B(n_1276),
.Y(n_2456)
);

NAND3xp33_ASAP7_75t_SL g2457 ( 
.A(n_2399),
.B(n_1129),
.C(n_1120),
.Y(n_2457)
);

NAND4xp25_ASAP7_75t_L g2458 ( 
.A(n_2413),
.B(n_1141),
.C(n_1130),
.D(n_1178),
.Y(n_2458)
);

INVx1_ASAP7_75t_L g2459 ( 
.A(n_2400),
.Y(n_2459)
);

AND2x4_ASAP7_75t_L g2460 ( 
.A(n_2398),
.B(n_186),
.Y(n_2460)
);

OR2x2_ASAP7_75t_L g2461 ( 
.A(n_2407),
.B(n_193),
.Y(n_2461)
);

OR2x2_ASAP7_75t_L g2462 ( 
.A(n_2380),
.B(n_2424),
.Y(n_2462)
);

INVx1_ASAP7_75t_L g2463 ( 
.A(n_2386),
.Y(n_2463)
);

NAND3xp33_ASAP7_75t_SL g2464 ( 
.A(n_2430),
.B(n_1623),
.C(n_1600),
.Y(n_2464)
);

INVx1_ASAP7_75t_L g2465 ( 
.A(n_2387),
.Y(n_2465)
);

NOR2xp33_ASAP7_75t_L g2466 ( 
.A(n_2412),
.B(n_216),
.Y(n_2466)
);

AOI211xp5_ASAP7_75t_L g2467 ( 
.A1(n_2410),
.A2(n_1239),
.B(n_1252),
.C(n_1259),
.Y(n_2467)
);

AOI22xp5_ASAP7_75t_L g2468 ( 
.A1(n_2388),
.A2(n_1692),
.B1(n_1625),
.B2(n_1651),
.Y(n_2468)
);

HB1xp67_ASAP7_75t_L g2469 ( 
.A(n_2382),
.Y(n_2469)
);

INVx2_ASAP7_75t_SL g2470 ( 
.A(n_2418),
.Y(n_2470)
);

AOI22xp33_ASAP7_75t_L g2471 ( 
.A1(n_2388),
.A2(n_1268),
.B1(n_1261),
.B2(n_1252),
.Y(n_2471)
);

XNOR2x1_ASAP7_75t_L g2472 ( 
.A(n_2394),
.B(n_217),
.Y(n_2472)
);

AND4x1_ASAP7_75t_L g2473 ( 
.A(n_2389),
.B(n_220),
.C(n_222),
.D(n_223),
.Y(n_2473)
);

INVx2_ASAP7_75t_SL g2474 ( 
.A(n_2428),
.Y(n_2474)
);

AOI222xp33_ASAP7_75t_L g2475 ( 
.A1(n_2402),
.A2(n_1656),
.B1(n_1668),
.B2(n_1697),
.C1(n_1650),
.C2(n_1643),
.Y(n_2475)
);

INVx1_ASAP7_75t_L g2476 ( 
.A(n_2379),
.Y(n_2476)
);

NAND2xp5_ASAP7_75t_L g2477 ( 
.A(n_2415),
.B(n_225),
.Y(n_2477)
);

INVx2_ASAP7_75t_L g2478 ( 
.A(n_2423),
.Y(n_2478)
);

XNOR2xp5_ASAP7_75t_L g2479 ( 
.A(n_2381),
.B(n_228),
.Y(n_2479)
);

NOR2x1p5_ASAP7_75t_L g2480 ( 
.A(n_2427),
.B(n_1252),
.Y(n_2480)
);

OAI211xp5_ASAP7_75t_L g2481 ( 
.A1(n_2438),
.A2(n_1268),
.B(n_1261),
.C(n_1259),
.Y(n_2481)
);

NAND2xp5_ASAP7_75t_SL g2482 ( 
.A(n_2405),
.B(n_1252),
.Y(n_2482)
);

OAI211xp5_ASAP7_75t_L g2483 ( 
.A1(n_2406),
.A2(n_1268),
.B(n_1261),
.C(n_1259),
.Y(n_2483)
);

NAND4xp25_ASAP7_75t_SL g2484 ( 
.A(n_2421),
.B(n_1988),
.C(n_1975),
.D(n_1639),
.Y(n_2484)
);

AOI221xp5_ASAP7_75t_L g2485 ( 
.A1(n_2437),
.A2(n_1268),
.B1(n_1261),
.B2(n_1259),
.C(n_1690),
.Y(n_2485)
);

NOR3xp33_ASAP7_75t_L g2486 ( 
.A(n_2390),
.B(n_1146),
.C(n_1191),
.Y(n_2486)
);

HB1xp67_ASAP7_75t_L g2487 ( 
.A(n_2434),
.Y(n_2487)
);

AOI22xp33_ASAP7_75t_SL g2488 ( 
.A1(n_2414),
.A2(n_1690),
.B1(n_1667),
.B2(n_1637),
.Y(n_2488)
);

NAND4xp25_ASAP7_75t_L g2489 ( 
.A(n_2431),
.B(n_1184),
.C(n_1189),
.D(n_1442),
.Y(n_2489)
);

INVx1_ASAP7_75t_L g2490 ( 
.A(n_2425),
.Y(n_2490)
);

AOI22xp33_ASAP7_75t_L g2491 ( 
.A1(n_2435),
.A2(n_1767),
.B1(n_1766),
.B2(n_1637),
.Y(n_2491)
);

INVx1_ASAP7_75t_SL g2492 ( 
.A(n_2408),
.Y(n_2492)
);

NAND4xp25_ASAP7_75t_L g2493 ( 
.A(n_2433),
.B(n_1189),
.C(n_1438),
.D(n_1441),
.Y(n_2493)
);

OA22x2_ASAP7_75t_L g2494 ( 
.A1(n_2440),
.A2(n_1708),
.B1(n_1667),
.B2(n_1593),
.Y(n_2494)
);

NOR4xp25_ASAP7_75t_L g2495 ( 
.A(n_2422),
.B(n_1589),
.C(n_1585),
.D(n_1568),
.Y(n_2495)
);

NOR3xp33_ASAP7_75t_L g2496 ( 
.A(n_2439),
.B(n_1146),
.C(n_1191),
.Y(n_2496)
);

AND2x2_ASAP7_75t_L g2497 ( 
.A(n_2416),
.B(n_1975),
.Y(n_2497)
);

INVx1_ASAP7_75t_L g2498 ( 
.A(n_2419),
.Y(n_2498)
);

NOR4xp25_ASAP7_75t_L g2499 ( 
.A(n_2444),
.B(n_230),
.C(n_232),
.D(n_234),
.Y(n_2499)
);

INVx1_ASAP7_75t_L g2500 ( 
.A(n_2461),
.Y(n_2500)
);

AOI21xp5_ASAP7_75t_L g2501 ( 
.A1(n_2474),
.A2(n_2441),
.B(n_2442),
.Y(n_2501)
);

OR4x1_ASAP7_75t_L g2502 ( 
.A(n_2476),
.B(n_2403),
.C(n_2432),
.D(n_2417),
.Y(n_2502)
);

HB1xp67_ASAP7_75t_L g2503 ( 
.A(n_2460),
.Y(n_2503)
);

NOR4xp25_ASAP7_75t_L g2504 ( 
.A(n_2448),
.B(n_2409),
.C(n_2443),
.D(n_2436),
.Y(n_2504)
);

INVx1_ASAP7_75t_L g2505 ( 
.A(n_2479),
.Y(n_2505)
);

OAI22xp5_ASAP7_75t_SL g2506 ( 
.A1(n_2478),
.A2(n_2392),
.B1(n_244),
.B2(n_245),
.Y(n_2506)
);

INVx2_ASAP7_75t_SL g2507 ( 
.A(n_2460),
.Y(n_2507)
);

XNOR2x1_ASAP7_75t_L g2508 ( 
.A(n_2472),
.B(n_2392),
.Y(n_2508)
);

NAND2xp5_ASAP7_75t_L g2509 ( 
.A(n_2492),
.B(n_236),
.Y(n_2509)
);

AO22x2_ASAP7_75t_L g2510 ( 
.A1(n_2470),
.A2(n_248),
.B1(n_250),
.B2(n_253),
.Y(n_2510)
);

NAND4xp75_ASAP7_75t_L g2511 ( 
.A(n_2466),
.B(n_262),
.C(n_265),
.D(n_266),
.Y(n_2511)
);

INVx2_ASAP7_75t_SL g2512 ( 
.A(n_2447),
.Y(n_2512)
);

INVx1_ASAP7_75t_L g2513 ( 
.A(n_2469),
.Y(n_2513)
);

INVx1_ASAP7_75t_L g2514 ( 
.A(n_2477),
.Y(n_2514)
);

INVx1_ASAP7_75t_L g2515 ( 
.A(n_2482),
.Y(n_2515)
);

INVx2_ASAP7_75t_L g2516 ( 
.A(n_2455),
.Y(n_2516)
);

OAI22x1_ASAP7_75t_L g2517 ( 
.A1(n_2490),
.A2(n_270),
.B1(n_273),
.B2(n_274),
.Y(n_2517)
);

INVx2_ASAP7_75t_L g2518 ( 
.A(n_2462),
.Y(n_2518)
);

INVx1_ASAP7_75t_L g2519 ( 
.A(n_2456),
.Y(n_2519)
);

NOR2xp33_ASAP7_75t_L g2520 ( 
.A(n_2446),
.B(n_278),
.Y(n_2520)
);

INVx1_ASAP7_75t_L g2521 ( 
.A(n_2487),
.Y(n_2521)
);

INVx1_ASAP7_75t_L g2522 ( 
.A(n_2494),
.Y(n_2522)
);

XNOR2x1_ASAP7_75t_L g2523 ( 
.A(n_2459),
.B(n_279),
.Y(n_2523)
);

NOR2xp33_ASAP7_75t_SL g2524 ( 
.A(n_2463),
.B(n_1146),
.Y(n_2524)
);

INVx2_ASAP7_75t_L g2525 ( 
.A(n_2480),
.Y(n_2525)
);

O2A1O1Ixp33_ASAP7_75t_L g2526 ( 
.A1(n_2498),
.A2(n_1210),
.B(n_1199),
.C(n_1191),
.Y(n_2526)
);

INVx1_ASAP7_75t_SL g2527 ( 
.A(n_2465),
.Y(n_2527)
);

INVx1_ASAP7_75t_L g2528 ( 
.A(n_2450),
.Y(n_2528)
);

HB1xp67_ASAP7_75t_L g2529 ( 
.A(n_2473),
.Y(n_2529)
);

NAND2xp5_ASAP7_75t_L g2530 ( 
.A(n_2467),
.B(n_280),
.Y(n_2530)
);

AND2x2_ASAP7_75t_L g2531 ( 
.A(n_2491),
.B(n_1974),
.Y(n_2531)
);

OA22x2_ASAP7_75t_L g2532 ( 
.A1(n_2468),
.A2(n_1516),
.B1(n_1533),
.B2(n_1559),
.Y(n_2532)
);

OAI221xp5_ASAP7_75t_L g2533 ( 
.A1(n_2499),
.A2(n_1687),
.B1(n_1708),
.B2(n_1210),
.C(n_1199),
.Y(n_2533)
);

AOI211xp5_ASAP7_75t_L g2534 ( 
.A1(n_2445),
.A2(n_2495),
.B(n_2489),
.C(n_2451),
.Y(n_2534)
);

NOR2x1p5_ASAP7_75t_L g2535 ( 
.A(n_2449),
.B(n_281),
.Y(n_2535)
);

AOI21xp5_ASAP7_75t_L g2536 ( 
.A1(n_2453),
.A2(n_1199),
.B(n_1210),
.Y(n_2536)
);

INVx3_ASAP7_75t_L g2537 ( 
.A(n_2497),
.Y(n_2537)
);

XOR2x2_ASAP7_75t_L g2538 ( 
.A(n_2464),
.B(n_282),
.Y(n_2538)
);

OAI22xp5_ASAP7_75t_L g2539 ( 
.A1(n_2488),
.A2(n_1581),
.B1(n_1573),
.B2(n_1571),
.Y(n_2539)
);

INVx1_ASAP7_75t_L g2540 ( 
.A(n_2454),
.Y(n_2540)
);

NAND3xp33_ASAP7_75t_L g2541 ( 
.A(n_2496),
.B(n_1173),
.C(n_1181),
.Y(n_2541)
);

OAI221xp5_ASAP7_75t_L g2542 ( 
.A1(n_2485),
.A2(n_287),
.B1(n_288),
.B2(n_293),
.C(n_296),
.Y(n_2542)
);

XNOR2xp5_ASAP7_75t_L g2543 ( 
.A(n_2483),
.B(n_302),
.Y(n_2543)
);

XNOR2x1_ASAP7_75t_L g2544 ( 
.A(n_2486),
.B(n_307),
.Y(n_2544)
);

INVx1_ASAP7_75t_L g2545 ( 
.A(n_2457),
.Y(n_2545)
);

OAI22xp5_ASAP7_75t_L g2546 ( 
.A1(n_2471),
.A2(n_1563),
.B1(n_1561),
.B2(n_1435),
.Y(n_2546)
);

AOI221xp5_ASAP7_75t_L g2547 ( 
.A1(n_2458),
.A2(n_1173),
.B1(n_1218),
.B2(n_1181),
.C(n_1182),
.Y(n_2547)
);

NOR2x1_ASAP7_75t_L g2548 ( 
.A(n_2481),
.B(n_1322),
.Y(n_2548)
);

NAND2x1_ASAP7_75t_L g2549 ( 
.A(n_2475),
.B(n_1689),
.Y(n_2549)
);

NOR3xp33_ASAP7_75t_L g2550 ( 
.A(n_2493),
.B(n_1439),
.C(n_309),
.Y(n_2550)
);

AOI22xp5_ASAP7_75t_L g2551 ( 
.A1(n_2484),
.A2(n_1689),
.B1(n_1322),
.B2(n_1371),
.Y(n_2551)
);

NAND4xp75_ASAP7_75t_L g2552 ( 
.A(n_2452),
.B(n_308),
.C(n_310),
.D(n_311),
.Y(n_2552)
);

NOR3xp33_ASAP7_75t_L g2553 ( 
.A(n_2448),
.B(n_317),
.C(n_324),
.Y(n_2553)
);

INVx1_ASAP7_75t_SL g2554 ( 
.A(n_2461),
.Y(n_2554)
);

AOI22xp5_ASAP7_75t_L g2555 ( 
.A1(n_2492),
.A2(n_1689),
.B1(n_1371),
.B2(n_1405),
.Y(n_2555)
);

NAND2xp5_ASAP7_75t_L g2556 ( 
.A(n_2476),
.B(n_327),
.Y(n_2556)
);

INVx1_ASAP7_75t_L g2557 ( 
.A(n_2461),
.Y(n_2557)
);

OR2x2_ASAP7_75t_L g2558 ( 
.A(n_2461),
.B(n_328),
.Y(n_2558)
);

NOR3xp33_ASAP7_75t_L g2559 ( 
.A(n_2512),
.B(n_1405),
.C(n_331),
.Y(n_2559)
);

NAND4xp25_ASAP7_75t_SL g2560 ( 
.A(n_2553),
.B(n_329),
.C(n_332),
.D(n_333),
.Y(n_2560)
);

OAI22xp5_ASAP7_75t_L g2561 ( 
.A1(n_2516),
.A2(n_1181),
.B1(n_1173),
.B2(n_1206),
.Y(n_2561)
);

BUFx2_ASAP7_75t_L g2562 ( 
.A(n_2503),
.Y(n_2562)
);

AOI22xp5_ASAP7_75t_SL g2563 ( 
.A1(n_2529),
.A2(n_2507),
.B1(n_2515),
.B2(n_2520),
.Y(n_2563)
);

AOI22xp5_ASAP7_75t_L g2564 ( 
.A1(n_2513),
.A2(n_1689),
.B1(n_1173),
.B2(n_1181),
.Y(n_2564)
);

AOI22xp33_ASAP7_75t_L g2565 ( 
.A1(n_2550),
.A2(n_1182),
.B1(n_1192),
.B2(n_1193),
.Y(n_2565)
);

OAI22xp5_ASAP7_75t_L g2566 ( 
.A1(n_2521),
.A2(n_1218),
.B1(n_1182),
.B2(n_1206),
.Y(n_2566)
);

AOI22xp5_ASAP7_75t_L g2567 ( 
.A1(n_2518),
.A2(n_1182),
.B1(n_1192),
.B2(n_1193),
.Y(n_2567)
);

NOR2x1_ASAP7_75t_L g2568 ( 
.A(n_2509),
.B(n_335),
.Y(n_2568)
);

NAND5xp2_ASAP7_75t_L g2569 ( 
.A(n_2534),
.B(n_337),
.C(n_344),
.D(n_345),
.E(n_346),
.Y(n_2569)
);

OR4x2_ASAP7_75t_L g2570 ( 
.A(n_2508),
.B(n_348),
.C(n_355),
.D(n_362),
.Y(n_2570)
);

AOI22xp33_ASAP7_75t_L g2571 ( 
.A1(n_2537),
.A2(n_1192),
.B1(n_1203),
.B2(n_1206),
.Y(n_2571)
);

INVx1_ASAP7_75t_L g2572 ( 
.A(n_2558),
.Y(n_2572)
);

INVx1_ASAP7_75t_L g2573 ( 
.A(n_2556),
.Y(n_2573)
);

OAI221xp5_ASAP7_75t_L g2574 ( 
.A1(n_2506),
.A2(n_364),
.B1(n_365),
.B2(n_366),
.C(n_367),
.Y(n_2574)
);

INVx1_ASAP7_75t_L g2575 ( 
.A(n_2538),
.Y(n_2575)
);

OAI22xp5_ASAP7_75t_L g2576 ( 
.A1(n_2527),
.A2(n_1218),
.B1(n_1192),
.B2(n_1206),
.Y(n_2576)
);

INVx3_ASAP7_75t_L g2577 ( 
.A(n_2511),
.Y(n_2577)
);

XNOR2xp5_ASAP7_75t_L g2578 ( 
.A(n_2523),
.B(n_368),
.Y(n_2578)
);

OAI22xp33_ASAP7_75t_L g2579 ( 
.A1(n_2554),
.A2(n_1203),
.B1(n_1218),
.B2(n_1193),
.Y(n_2579)
);

AND2x4_ASAP7_75t_L g2580 ( 
.A(n_2535),
.B(n_372),
.Y(n_2580)
);

AOI22xp5_ASAP7_75t_L g2581 ( 
.A1(n_2514),
.A2(n_1203),
.B1(n_1193),
.B2(n_1292),
.Y(n_2581)
);

INVx2_ASAP7_75t_L g2582 ( 
.A(n_2517),
.Y(n_2582)
);

OAI22xp5_ASAP7_75t_L g2583 ( 
.A1(n_2505),
.A2(n_1203),
.B1(n_1518),
.B2(n_1389),
.Y(n_2583)
);

NAND3xp33_ASAP7_75t_L g2584 ( 
.A(n_2500),
.B(n_1356),
.C(n_1349),
.Y(n_2584)
);

AND2x4_ASAP7_75t_L g2585 ( 
.A(n_2557),
.B(n_374),
.Y(n_2585)
);

OAI221xp5_ASAP7_75t_L g2586 ( 
.A1(n_2533),
.A2(n_379),
.B1(n_382),
.B2(n_383),
.C(n_386),
.Y(n_2586)
);

INVxp67_ASAP7_75t_L g2587 ( 
.A(n_2530),
.Y(n_2587)
);

INVx1_ASAP7_75t_L g2588 ( 
.A(n_2544),
.Y(n_2588)
);

NAND3xp33_ASAP7_75t_SL g2589 ( 
.A(n_2504),
.B(n_388),
.C(n_398),
.Y(n_2589)
);

NOR2xp33_ASAP7_75t_L g2590 ( 
.A(n_2522),
.B(n_400),
.Y(n_2590)
);

NOR4xp75_ASAP7_75t_L g2591 ( 
.A(n_2552),
.B(n_407),
.C(n_408),
.D(n_409),
.Y(n_2591)
);

OAI22xp33_ASAP7_75t_L g2592 ( 
.A1(n_2542),
.A2(n_1296),
.B1(n_1292),
.B2(n_1440),
.Y(n_2592)
);

OR4x2_ASAP7_75t_L g2593 ( 
.A(n_2502),
.B(n_414),
.C(n_415),
.D(n_424),
.Y(n_2593)
);

XOR2xp5_ASAP7_75t_L g2594 ( 
.A(n_2543),
.B(n_426),
.Y(n_2594)
);

INVx2_ASAP7_75t_L g2595 ( 
.A(n_2570),
.Y(n_2595)
);

AND2x2_ASAP7_75t_SL g2596 ( 
.A(n_2562),
.B(n_2528),
.Y(n_2596)
);

INVx2_ASAP7_75t_L g2597 ( 
.A(n_2593),
.Y(n_2597)
);

CKINVDCx5p33_ASAP7_75t_R g2598 ( 
.A(n_2563),
.Y(n_2598)
);

INVx1_ASAP7_75t_L g2599 ( 
.A(n_2578),
.Y(n_2599)
);

AND2x2_ASAP7_75t_SL g2600 ( 
.A(n_2582),
.B(n_2545),
.Y(n_2600)
);

INVx2_ASAP7_75t_L g2601 ( 
.A(n_2580),
.Y(n_2601)
);

AND2x2_ASAP7_75t_L g2602 ( 
.A(n_2580),
.B(n_2568),
.Y(n_2602)
);

INVx2_ASAP7_75t_L g2603 ( 
.A(n_2585),
.Y(n_2603)
);

INVx3_ASAP7_75t_L g2604 ( 
.A(n_2577),
.Y(n_2604)
);

OAI21x1_ASAP7_75t_SL g2605 ( 
.A1(n_2594),
.A2(n_2501),
.B(n_2525),
.Y(n_2605)
);

OR2x2_ASAP7_75t_L g2606 ( 
.A(n_2569),
.B(n_2549),
.Y(n_2606)
);

INVx1_ASAP7_75t_L g2607 ( 
.A(n_2572),
.Y(n_2607)
);

INVx2_ASAP7_75t_L g2608 ( 
.A(n_2585),
.Y(n_2608)
);

XOR2x2_ASAP7_75t_L g2609 ( 
.A(n_2591),
.B(n_2548),
.Y(n_2609)
);

AOI21xp5_ASAP7_75t_L g2610 ( 
.A1(n_2589),
.A2(n_2587),
.B(n_2573),
.Y(n_2610)
);

INVx4_ASAP7_75t_L g2611 ( 
.A(n_2575),
.Y(n_2611)
);

INVx1_ASAP7_75t_SL g2612 ( 
.A(n_2590),
.Y(n_2612)
);

XNOR2xp5_ASAP7_75t_L g2613 ( 
.A(n_2588),
.B(n_2519),
.Y(n_2613)
);

AOI22xp5_ASAP7_75t_L g2614 ( 
.A1(n_2560),
.A2(n_2540),
.B1(n_2524),
.B2(n_2551),
.Y(n_2614)
);

INVx1_ASAP7_75t_L g2615 ( 
.A(n_2584),
.Y(n_2615)
);

OAI22xp5_ASAP7_75t_L g2616 ( 
.A1(n_2574),
.A2(n_2555),
.B1(n_2541),
.B2(n_2547),
.Y(n_2616)
);

INVx3_ASAP7_75t_L g2617 ( 
.A(n_2559),
.Y(n_2617)
);

INVx2_ASAP7_75t_L g2618 ( 
.A(n_2586),
.Y(n_2618)
);

OAI22x1_ASAP7_75t_L g2619 ( 
.A1(n_2567),
.A2(n_2581),
.B1(n_2564),
.B2(n_2531),
.Y(n_2619)
);

OR2x6_ASAP7_75t_L g2620 ( 
.A(n_2603),
.B(n_2526),
.Y(n_2620)
);

AOI22xp5_ASAP7_75t_L g2621 ( 
.A1(n_2598),
.A2(n_2592),
.B1(n_2565),
.B2(n_2532),
.Y(n_2621)
);

AOI21xp5_ASAP7_75t_L g2622 ( 
.A1(n_2596),
.A2(n_2536),
.B(n_2566),
.Y(n_2622)
);

INVx1_ASAP7_75t_L g2623 ( 
.A(n_2602),
.Y(n_2623)
);

AOI21xp5_ASAP7_75t_L g2624 ( 
.A1(n_2610),
.A2(n_2579),
.B(n_2583),
.Y(n_2624)
);

OAI221xp5_ASAP7_75t_L g2625 ( 
.A1(n_2607),
.A2(n_2571),
.B1(n_2576),
.B2(n_2561),
.C(n_2539),
.Y(n_2625)
);

INVx1_ASAP7_75t_L g2626 ( 
.A(n_2608),
.Y(n_2626)
);

XNOR2xp5_ASAP7_75t_L g2627 ( 
.A(n_2613),
.B(n_2510),
.Y(n_2627)
);

AOI21xp5_ASAP7_75t_L g2628 ( 
.A1(n_2600),
.A2(n_2546),
.B(n_2510),
.Y(n_2628)
);

NOR2xp67_ASAP7_75t_SL g2629 ( 
.A(n_2604),
.B(n_2601),
.Y(n_2629)
);

INVx1_ASAP7_75t_L g2630 ( 
.A(n_2606),
.Y(n_2630)
);

INVx1_ASAP7_75t_L g2631 ( 
.A(n_2595),
.Y(n_2631)
);

INVx2_ASAP7_75t_L g2632 ( 
.A(n_2597),
.Y(n_2632)
);

INVx1_ASAP7_75t_L g2633 ( 
.A(n_2609),
.Y(n_2633)
);

CKINVDCx14_ASAP7_75t_R g2634 ( 
.A(n_2611),
.Y(n_2634)
);

AO22x2_ASAP7_75t_L g2635 ( 
.A1(n_2612),
.A2(n_427),
.B1(n_432),
.B2(n_434),
.Y(n_2635)
);

INVx1_ASAP7_75t_L g2636 ( 
.A(n_2599),
.Y(n_2636)
);

AOI21xp33_ASAP7_75t_L g2637 ( 
.A1(n_2629),
.A2(n_2605),
.B(n_2618),
.Y(n_2637)
);

NOR3xp33_ASAP7_75t_L g2638 ( 
.A(n_2634),
.B(n_2617),
.C(n_2616),
.Y(n_2638)
);

AND2x2_ASAP7_75t_L g2639 ( 
.A(n_2626),
.B(n_2614),
.Y(n_2639)
);

INVx1_ASAP7_75t_L g2640 ( 
.A(n_2627),
.Y(n_2640)
);

AOI22x1_ASAP7_75t_L g2641 ( 
.A1(n_2623),
.A2(n_2619),
.B1(n_2615),
.B2(n_446),
.Y(n_2641)
);

CKINVDCx20_ASAP7_75t_R g2642 ( 
.A(n_2633),
.Y(n_2642)
);

OAI22xp5_ASAP7_75t_SL g2643 ( 
.A1(n_2631),
.A2(n_2619),
.B1(n_442),
.B2(n_452),
.Y(n_2643)
);

AOI21xp5_ASAP7_75t_L g2644 ( 
.A1(n_2628),
.A2(n_1275),
.B(n_1254),
.Y(n_2644)
);

AOI22xp5_ASAP7_75t_L g2645 ( 
.A1(n_2632),
.A2(n_1301),
.B1(n_1440),
.B2(n_1437),
.Y(n_2645)
);

INVx1_ASAP7_75t_L g2646 ( 
.A(n_2630),
.Y(n_2646)
);

AOI22xp5_ASAP7_75t_L g2647 ( 
.A1(n_2636),
.A2(n_1301),
.B1(n_1440),
.B2(n_1437),
.Y(n_2647)
);

INVx1_ASAP7_75t_L g2648 ( 
.A(n_2620),
.Y(n_2648)
);

OAI22xp5_ASAP7_75t_SL g2649 ( 
.A1(n_2621),
.A2(n_437),
.B1(n_453),
.B2(n_455),
.Y(n_2649)
);

HB1xp67_ASAP7_75t_L g2650 ( 
.A(n_2635),
.Y(n_2650)
);

NOR3xp33_ASAP7_75t_L g2651 ( 
.A(n_2637),
.B(n_2646),
.C(n_2640),
.Y(n_2651)
);

INVx1_ASAP7_75t_L g2652 ( 
.A(n_2641),
.Y(n_2652)
);

OAI22xp5_ASAP7_75t_L g2653 ( 
.A1(n_2642),
.A2(n_2620),
.B1(n_2625),
.B2(n_2622),
.Y(n_2653)
);

INVx1_ASAP7_75t_L g2654 ( 
.A(n_2650),
.Y(n_2654)
);

AOI22xp5_ASAP7_75t_L g2655 ( 
.A1(n_2639),
.A2(n_2624),
.B1(n_1339),
.B2(n_1349),
.Y(n_2655)
);

AND3x4_ASAP7_75t_L g2656 ( 
.A(n_2638),
.B(n_2648),
.C(n_2643),
.Y(n_2656)
);

INVx1_ASAP7_75t_L g2657 ( 
.A(n_2649),
.Y(n_2657)
);

INVx2_ASAP7_75t_L g2658 ( 
.A(n_2645),
.Y(n_2658)
);

AOI22xp5_ASAP7_75t_SL g2659 ( 
.A1(n_2644),
.A2(n_456),
.B1(n_457),
.B2(n_460),
.Y(n_2659)
);

INVx3_ASAP7_75t_SL g2660 ( 
.A(n_2647),
.Y(n_2660)
);

XOR2xp5_ASAP7_75t_L g2661 ( 
.A(n_2653),
.B(n_467),
.Y(n_2661)
);

OAI22xp33_ASAP7_75t_L g2662 ( 
.A1(n_2654),
.A2(n_468),
.B1(n_1356),
.B2(n_1436),
.Y(n_2662)
);

AOI21x1_ASAP7_75t_L g2663 ( 
.A1(n_2652),
.A2(n_1391),
.B(n_1390),
.Y(n_2663)
);

AOI21xp5_ASAP7_75t_L g2664 ( 
.A1(n_2656),
.A2(n_1275),
.B(n_1254),
.Y(n_2664)
);

AOI21xp33_ASAP7_75t_SL g2665 ( 
.A1(n_2651),
.A2(n_1391),
.B(n_1390),
.Y(n_2665)
);

OAI21xp5_ASAP7_75t_SL g2666 ( 
.A1(n_2657),
.A2(n_1349),
.B(n_1414),
.Y(n_2666)
);

AOI21xp33_ASAP7_75t_L g2667 ( 
.A1(n_2658),
.A2(n_1275),
.B(n_1254),
.Y(n_2667)
);

INVx1_ASAP7_75t_L g2668 ( 
.A(n_2661),
.Y(n_2668)
);

HB1xp67_ASAP7_75t_L g2669 ( 
.A(n_2663),
.Y(n_2669)
);

INVx1_ASAP7_75t_L g2670 ( 
.A(n_2665),
.Y(n_2670)
);

NAND2xp5_ASAP7_75t_L g2671 ( 
.A(n_2666),
.B(n_2660),
.Y(n_2671)
);

OR2x6_ASAP7_75t_L g2672 ( 
.A(n_2668),
.B(n_2664),
.Y(n_2672)
);

OAI21xp5_ASAP7_75t_L g2673 ( 
.A1(n_2671),
.A2(n_2655),
.B(n_2667),
.Y(n_2673)
);

AOI22xp5_ASAP7_75t_SL g2674 ( 
.A1(n_2669),
.A2(n_2659),
.B1(n_2662),
.B2(n_1356),
.Y(n_2674)
);

NAND2xp5_ASAP7_75t_L g2675 ( 
.A(n_2670),
.B(n_1275),
.Y(n_2675)
);

HB1xp67_ASAP7_75t_L g2676 ( 
.A(n_2672),
.Y(n_2676)
);

INVx1_ASAP7_75t_L g2677 ( 
.A(n_2675),
.Y(n_2677)
);

OR2x6_ASAP7_75t_L g2678 ( 
.A(n_2676),
.B(n_2673),
.Y(n_2678)
);

OR2x6_ASAP7_75t_L g2679 ( 
.A(n_2677),
.B(n_2674),
.Y(n_2679)
);

OR2x6_ASAP7_75t_L g2680 ( 
.A(n_2676),
.B(n_1389),
.Y(n_2680)
);

AOI21xp5_ASAP7_75t_L g2681 ( 
.A1(n_2678),
.A2(n_1275),
.B(n_1254),
.Y(n_2681)
);

AOI211xp5_ASAP7_75t_L g2682 ( 
.A1(n_2681),
.A2(n_2679),
.B(n_2680),
.C(n_1356),
.Y(n_2682)
);


endmodule