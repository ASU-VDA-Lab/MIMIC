module fake_jpeg_13235_n_163 (n_13, n_21, n_33, n_1, n_45, n_10, n_23, n_27, n_6, n_22, n_47, n_14, n_40, n_19, n_18, n_20, n_35, n_48, n_46, n_41, n_4, n_34, n_30, n_39, n_42, n_16, n_3, n_0, n_24, n_28, n_38, n_26, n_44, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_43, n_12, n_32, n_8, n_15, n_7, n_163);

input n_13;
input n_21;
input n_33;
input n_1;
input n_45;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_47;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_48;
input n_46;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_42;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_44;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_43;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_163;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_51;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_84;
wire n_59;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_155;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_57;
wire n_119;
wire n_69;
wire n_83;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_106;
wire n_111;
wire n_143;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_77;
wire n_136;
wire n_61;
wire n_139;
wire n_78;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_162;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_54;
wire n_91;
wire n_93;
wire n_161;
wire n_138;
wire n_101;
wire n_149;
wire n_157;
wire n_87;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_153;
wire n_135;
wire n_62;
wire n_120;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_3),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_SL g50 ( 
.A(n_1),
.B(n_38),
.Y(n_50)
);

INVx4_ASAP7_75t_L g51 ( 
.A(n_29),
.Y(n_51)
);

INVx13_ASAP7_75t_L g52 ( 
.A(n_5),
.Y(n_52)
);

BUFx12_ASAP7_75t_L g53 ( 
.A(n_4),
.Y(n_53)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_47),
.Y(n_54)
);

INVx11_ASAP7_75t_L g55 ( 
.A(n_46),
.Y(n_55)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_26),
.Y(n_56)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_15),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_4),
.Y(n_58)
);

BUFx12_ASAP7_75t_L g59 ( 
.A(n_22),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_0),
.Y(n_60)
);

INVx13_ASAP7_75t_L g61 ( 
.A(n_0),
.Y(n_61)
);

INVx8_ASAP7_75t_L g62 ( 
.A(n_34),
.Y(n_62)
);

CKINVDCx20_ASAP7_75t_R g63 ( 
.A(n_6),
.Y(n_63)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_33),
.Y(n_64)
);

INVx5_ASAP7_75t_L g65 ( 
.A(n_36),
.Y(n_65)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_12),
.Y(n_66)
);

BUFx12f_ASAP7_75t_L g67 ( 
.A(n_11),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_30),
.B(n_31),
.Y(n_68)
);

INVx8_ASAP7_75t_L g69 ( 
.A(n_13),
.Y(n_69)
);

INVx3_ASAP7_75t_SL g70 ( 
.A(n_62),
.Y(n_70)
);

INVx2_ASAP7_75t_L g84 ( 
.A(n_70),
.Y(n_84)
);

CKINVDCx20_ASAP7_75t_R g71 ( 
.A(n_55),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_71),
.B(n_73),
.Y(n_79)
);

BUFx6f_ASAP7_75t_L g72 ( 
.A(n_64),
.Y(n_72)
);

INVx3_ASAP7_75t_L g90 ( 
.A(n_72),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_49),
.B(n_1),
.Y(n_73)
);

INVx2_ASAP7_75t_L g74 ( 
.A(n_54),
.Y(n_74)
);

INVx2_ASAP7_75t_L g88 ( 
.A(n_74),
.Y(n_88)
);

AND2x2_ASAP7_75t_L g75 ( 
.A(n_67),
.B(n_2),
.Y(n_75)
);

OAI21xp33_ASAP7_75t_L g80 ( 
.A1(n_75),
.A2(n_50),
.B(n_5),
.Y(n_80)
);

A2O1A1Ixp33_ASAP7_75t_L g76 ( 
.A1(n_68),
.A2(n_23),
.B(n_45),
.C(n_44),
.Y(n_76)
);

OR2x2_ASAP7_75t_L g86 ( 
.A(n_76),
.B(n_65),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_SL g77 ( 
.A(n_50),
.B(n_68),
.Y(n_77)
);

AND2x2_ASAP7_75t_L g83 ( 
.A(n_77),
.B(n_63),
.Y(n_83)
);

INVx11_ASAP7_75t_L g78 ( 
.A(n_52),
.Y(n_78)
);

BUFx10_ASAP7_75t_L g85 ( 
.A(n_78),
.Y(n_85)
);

OAI21xp5_ASAP7_75t_SL g106 ( 
.A1(n_80),
.A2(n_76),
.B(n_61),
.Y(n_106)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_74),
.Y(n_81)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_81),
.Y(n_96)
);

INVx2_ASAP7_75t_SL g82 ( 
.A(n_78),
.Y(n_82)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_82),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g93 ( 
.A(n_86),
.B(n_87),
.Y(n_93)
);

CKINVDCx20_ASAP7_75t_R g87 ( 
.A(n_75),
.Y(n_87)
);

INVx13_ASAP7_75t_L g89 ( 
.A(n_70),
.Y(n_89)
);

BUFx12f_ASAP7_75t_L g109 ( 
.A(n_89),
.Y(n_109)
);

OAI22xp5_ASAP7_75t_L g91 ( 
.A1(n_86),
.A2(n_72),
.B1(n_58),
.B2(n_60),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_L g128 ( 
.A(n_91),
.B(n_94),
.Y(n_128)
);

OAI22xp33_ASAP7_75t_SL g92 ( 
.A1(n_88),
.A2(n_60),
.B1(n_58),
.B2(n_64),
.Y(n_92)
);

AOI22xp33_ASAP7_75t_SL g110 ( 
.A1(n_92),
.A2(n_102),
.B1(n_108),
.B2(n_53),
.Y(n_110)
);

OAI22xp5_ASAP7_75t_L g94 ( 
.A1(n_80),
.A2(n_66),
.B1(n_51),
.B2(n_62),
.Y(n_94)
);

CKINVDCx16_ASAP7_75t_R g95 ( 
.A(n_85),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_95),
.B(n_104),
.Y(n_111)
);

INVx3_ASAP7_75t_L g97 ( 
.A(n_84),
.Y(n_97)
);

INVx2_ASAP7_75t_SL g113 ( 
.A(n_97),
.Y(n_113)
);

INVx4_ASAP7_75t_L g99 ( 
.A(n_84),
.Y(n_99)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_99),
.Y(n_123)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_90),
.Y(n_100)
);

INVxp67_ASAP7_75t_L g114 ( 
.A(n_100),
.Y(n_114)
);

MAJIxp5_ASAP7_75t_L g101 ( 
.A(n_83),
.B(n_56),
.C(n_57),
.Y(n_101)
);

MAJIxp5_ASAP7_75t_L g120 ( 
.A(n_101),
.B(n_106),
.C(n_107),
.Y(n_120)
);

OAI22xp5_ASAP7_75t_SL g102 ( 
.A1(n_90),
.A2(n_66),
.B1(n_67),
.B2(n_79),
.Y(n_102)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_82),
.Y(n_103)
);

INVxp67_ASAP7_75t_L g125 ( 
.A(n_103),
.Y(n_125)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_85),
.Y(n_104)
);

CKINVDCx20_ASAP7_75t_R g105 ( 
.A(n_85),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_L g119 ( 
.A(n_105),
.B(n_27),
.Y(n_119)
);

MAJIxp5_ASAP7_75t_L g107 ( 
.A(n_89),
.B(n_59),
.C(n_61),
.Y(n_107)
);

AOI22xp33_ASAP7_75t_SL g108 ( 
.A1(n_87),
.A2(n_69),
.B1(n_52),
.B2(n_53),
.Y(n_108)
);

INVxp67_ASAP7_75t_L g143 ( 
.A(n_110),
.Y(n_143)
);

CKINVDCx20_ASAP7_75t_R g112 ( 
.A(n_96),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_L g129 ( 
.A(n_112),
.B(n_119),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_L g115 ( 
.A(n_93),
.B(n_7),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_SL g140 ( 
.A(n_115),
.B(n_116),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_SL g116 ( 
.A(n_108),
.B(n_7),
.Y(n_116)
);

MAJIxp5_ASAP7_75t_SL g117 ( 
.A(n_98),
.B(n_8),
.C(n_9),
.Y(n_117)
);

AOI21xp5_ASAP7_75t_L g131 ( 
.A1(n_117),
.A2(n_48),
.B(n_20),
.Y(n_131)
);

NOR2x1_ASAP7_75t_L g118 ( 
.A(n_109),
.B(n_8),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_L g137 ( 
.A(n_118),
.B(n_122),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_SL g121 ( 
.A(n_109),
.B(n_10),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_L g142 ( 
.A(n_121),
.B(n_122),
.Y(n_142)
);

NOR2x1_ASAP7_75t_L g122 ( 
.A(n_109),
.B(n_10),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_92),
.B(n_14),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_L g138 ( 
.A(n_124),
.B(n_126),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_L g126 ( 
.A(n_93),
.B(n_16),
.Y(n_126)
);

XOR2xp5_ASAP7_75t_L g127 ( 
.A(n_93),
.B(n_59),
.Y(n_127)
);

MAJIxp5_ASAP7_75t_L g130 ( 
.A(n_127),
.B(n_17),
.C(n_18),
.Y(n_130)
);

XOR2xp5_ASAP7_75t_L g149 ( 
.A(n_130),
.B(n_125),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_L g146 ( 
.A(n_131),
.B(n_132),
.Y(n_146)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_123),
.Y(n_132)
);

AOI22xp33_ASAP7_75t_SL g133 ( 
.A1(n_128),
.A2(n_43),
.B1(n_21),
.B2(n_24),
.Y(n_133)
);

AOI21xp5_ASAP7_75t_L g144 ( 
.A1(n_133),
.A2(n_135),
.B(n_130),
.Y(n_144)
);

AOI22xp5_ASAP7_75t_L g134 ( 
.A1(n_110),
.A2(n_19),
.B1(n_25),
.B2(n_28),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_L g148 ( 
.A(n_134),
.B(n_136),
.Y(n_148)
);

AO21x1_ASAP7_75t_L g135 ( 
.A1(n_118),
.A2(n_32),
.B(n_35),
.Y(n_135)
);

AOI22xp5_ASAP7_75t_L g136 ( 
.A1(n_127),
.A2(n_37),
.B1(n_39),
.B2(n_40),
.Y(n_136)
);

OAI22xp5_ASAP7_75t_SL g139 ( 
.A1(n_111),
.A2(n_41),
.B1(n_42),
.B2(n_120),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_L g151 ( 
.A(n_139),
.B(n_141),
.Y(n_151)
);

BUFx3_ASAP7_75t_L g141 ( 
.A(n_113),
.Y(n_141)
);

CKINVDCx20_ASAP7_75t_R g145 ( 
.A(n_142),
.Y(n_145)
);

MAJIxp5_ASAP7_75t_L g155 ( 
.A(n_144),
.B(n_147),
.C(n_149),
.Y(n_155)
);

AOI21xp5_ASAP7_75t_L g147 ( 
.A1(n_143),
.A2(n_137),
.B(n_140),
.Y(n_147)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_141),
.Y(n_150)
);

XOR2xp5_ASAP7_75t_L g154 ( 
.A(n_150),
.B(n_114),
.Y(n_154)
);

OA21x2_ASAP7_75t_L g152 ( 
.A1(n_148),
.A2(n_143),
.B(n_138),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_L g157 ( 
.A(n_152),
.B(n_153),
.Y(n_157)
);

XOR2xp5_ASAP7_75t_L g153 ( 
.A(n_149),
.B(n_129),
.Y(n_153)
);

AOI21xp5_ASAP7_75t_L g156 ( 
.A1(n_154),
.A2(n_125),
.B(n_114),
.Y(n_156)
);

NAND2xp33_ASAP7_75t_SL g158 ( 
.A(n_156),
.B(n_146),
.Y(n_158)
);

XOR2xp5_ASAP7_75t_L g159 ( 
.A(n_158),
.B(n_157),
.Y(n_159)
);

OAI22xp5_ASAP7_75t_SL g160 ( 
.A1(n_159),
.A2(n_155),
.B1(n_133),
.B2(n_135),
.Y(n_160)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_160),
.Y(n_161)
);

NAND3xp33_ASAP7_75t_SL g162 ( 
.A(n_161),
.B(n_145),
.C(n_152),
.Y(n_162)
);

XOR2xp5_ASAP7_75t_L g163 ( 
.A(n_162),
.B(n_151),
.Y(n_163)
);


endmodule