module fake_jpeg_20298_n_311 (n_3, n_2, n_1, n_0, n_10, n_4, n_8, n_9, n_6, n_5, n_7, n_311);

input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_311;

wire n_253;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_15;
wire n_141;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_13;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_11;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_14;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_20;
wire n_18;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_12;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_208;
wire n_308;
wire n_297;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

CKINVDCx20_ASAP7_75t_R g11 ( 
.A(n_0),
.Y(n_11)
);

INVxp67_ASAP7_75t_L g12 ( 
.A(n_6),
.Y(n_12)
);

BUFx16f_ASAP7_75t_L g13 ( 
.A(n_7),
.Y(n_13)
);

INVx1_ASAP7_75t_L g14 ( 
.A(n_6),
.Y(n_14)
);

INVx1_ASAP7_75t_L g15 ( 
.A(n_9),
.Y(n_15)
);

NOR2xp33_ASAP7_75t_L g16 ( 
.A(n_6),
.B(n_8),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_4),
.Y(n_17)
);

INVx11_ASAP7_75t_L g18 ( 
.A(n_8),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_2),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_1),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_1),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_4),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_2),
.Y(n_23)
);

AND2x2_ASAP7_75t_L g24 ( 
.A(n_16),
.B(n_10),
.Y(n_24)
);

OAI21xp33_ASAP7_75t_L g44 ( 
.A1(n_24),
.A2(n_10),
.B(n_9),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_20),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_25),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g26 ( 
.A(n_16),
.B(n_10),
.Y(n_26)
);

OR2x2_ASAP7_75t_L g40 ( 
.A(n_26),
.B(n_32),
.Y(n_40)
);

INVx2_ASAP7_75t_L g27 ( 
.A(n_20),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_27),
.Y(n_43)
);

INVx3_ASAP7_75t_L g28 ( 
.A(n_13),
.Y(n_28)
);

INVx2_ASAP7_75t_L g39 ( 
.A(n_28),
.Y(n_39)
);

BUFx12f_ASAP7_75t_L g29 ( 
.A(n_20),
.Y(n_29)
);

BUFx2_ASAP7_75t_L g38 ( 
.A(n_29),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_20),
.Y(n_30)
);

INVx6_ASAP7_75t_L g41 ( 
.A(n_30),
.Y(n_41)
);

BUFx5_ASAP7_75t_L g31 ( 
.A(n_20),
.Y(n_31)
);

BUFx24_ASAP7_75t_L g37 ( 
.A(n_31),
.Y(n_37)
);

INVx2_ASAP7_75t_L g32 ( 
.A(n_13),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_13),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_33),
.Y(n_34)
);

A2O1A1Ixp33_ASAP7_75t_L g36 ( 
.A1(n_24),
.A2(n_12),
.B(n_16),
.C(n_15),
.Y(n_36)
);

AOI21xp5_ASAP7_75t_L g53 ( 
.A1(n_36),
.A2(n_24),
.B(n_26),
.Y(n_53)
);

OAI22xp5_ASAP7_75t_SL g42 ( 
.A1(n_27),
.A2(n_12),
.B1(n_15),
.B2(n_19),
.Y(n_42)
);

AOI22xp5_ASAP7_75t_L g57 ( 
.A1(n_42),
.A2(n_15),
.B1(n_11),
.B2(n_22),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_SL g55 ( 
.A(n_44),
.B(n_8),
.Y(n_55)
);

BUFx3_ASAP7_75t_L g45 ( 
.A(n_37),
.Y(n_45)
);

BUFx3_ASAP7_75t_L g63 ( 
.A(n_45),
.Y(n_63)
);

INVx3_ASAP7_75t_L g46 ( 
.A(n_39),
.Y(n_46)
);

INVx2_ASAP7_75t_L g78 ( 
.A(n_46),
.Y(n_78)
);

BUFx10_ASAP7_75t_L g47 ( 
.A(n_37),
.Y(n_47)
);

BUFx2_ASAP7_75t_L g80 ( 
.A(n_47),
.Y(n_80)
);

CKINVDCx12_ASAP7_75t_R g48 ( 
.A(n_37),
.Y(n_48)
);

CKINVDCx16_ASAP7_75t_R g73 ( 
.A(n_48),
.Y(n_73)
);

AOI22xp33_ASAP7_75t_SL g49 ( 
.A1(n_41),
.A2(n_18),
.B1(n_32),
.B2(n_15),
.Y(n_49)
);

OAI22xp5_ASAP7_75t_SL g79 ( 
.A1(n_49),
.A2(n_57),
.B1(n_60),
.B2(n_21),
.Y(n_79)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_35),
.Y(n_50)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_50),
.Y(n_70)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_43),
.Y(n_51)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_51),
.Y(n_74)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_43),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_SL g76 ( 
.A(n_52),
.B(n_53),
.Y(n_76)
);

OAI22xp5_ASAP7_75t_SL g54 ( 
.A1(n_40),
.A2(n_28),
.B1(n_30),
.B2(n_25),
.Y(n_54)
);

AOI22xp5_ASAP7_75t_L g61 ( 
.A1(n_54),
.A2(n_42),
.B1(n_41),
.B2(n_34),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_55),
.B(n_11),
.Y(n_65)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_43),
.Y(n_56)
);

INVx3_ASAP7_75t_L g62 ( 
.A(n_56),
.Y(n_62)
);

AND2x2_ASAP7_75t_L g58 ( 
.A(n_40),
.B(n_29),
.Y(n_58)
);

MAJIxp5_ASAP7_75t_L g71 ( 
.A(n_58),
.B(n_29),
.C(n_33),
.Y(n_71)
);

BUFx12f_ASAP7_75t_L g59 ( 
.A(n_37),
.Y(n_59)
);

CKINVDCx20_ASAP7_75t_R g77 ( 
.A(n_59),
.Y(n_77)
);

AOI22xp5_ASAP7_75t_SL g60 ( 
.A1(n_36),
.A2(n_19),
.B1(n_21),
.B2(n_17),
.Y(n_60)
);

OAI22xp5_ASAP7_75t_L g91 ( 
.A1(n_61),
.A2(n_66),
.B1(n_67),
.B2(n_52),
.Y(n_91)
);

NAND2xp33_ASAP7_75t_SL g64 ( 
.A(n_58),
.B(n_40),
.Y(n_64)
);

AO21x1_ASAP7_75t_L g86 ( 
.A1(n_64),
.A2(n_68),
.B(n_72),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_65),
.B(n_79),
.Y(n_82)
);

OAI22xp33_ASAP7_75t_L g66 ( 
.A1(n_57),
.A2(n_41),
.B1(n_34),
.B2(n_39),
.Y(n_66)
);

OAI22xp33_ASAP7_75t_SL g67 ( 
.A1(n_60),
.A2(n_36),
.B1(n_37),
.B2(n_11),
.Y(n_67)
);

AND2x2_ASAP7_75t_L g68 ( 
.A(n_58),
.B(n_29),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_L g69 ( 
.A(n_58),
.B(n_35),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_L g81 ( 
.A(n_69),
.B(n_75),
.Y(n_81)
);

AND2x2_ASAP7_75t_L g95 ( 
.A(n_71),
.B(n_33),
.Y(n_95)
);

AO22x2_ASAP7_75t_L g72 ( 
.A1(n_54),
.A2(n_30),
.B1(n_25),
.B2(n_31),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_L g75 ( 
.A(n_53),
.B(n_35),
.Y(n_75)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_74),
.Y(n_83)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_83),
.Y(n_112)
);

INVx2_ASAP7_75t_L g84 ( 
.A(n_62),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g119 ( 
.A(n_84),
.B(n_88),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_75),
.B(n_55),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_L g110 ( 
.A(n_85),
.B(n_92),
.Y(n_110)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_74),
.Y(n_87)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_87),
.Y(n_116)
);

AND2x6_ASAP7_75t_L g88 ( 
.A(n_76),
.B(n_48),
.Y(n_88)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_70),
.Y(n_89)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_89),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_73),
.B(n_46),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_SL g104 ( 
.A(n_90),
.B(n_95),
.Y(n_104)
);

AOI22xp5_ASAP7_75t_L g106 ( 
.A1(n_91),
.A2(n_94),
.B1(n_79),
.B2(n_72),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_65),
.B(n_46),
.Y(n_92)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_70),
.Y(n_93)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_93),
.Y(n_124)
);

OAI22xp5_ASAP7_75t_L g94 ( 
.A1(n_61),
.A2(n_51),
.B1(n_56),
.B2(n_18),
.Y(n_94)
);

INVx3_ASAP7_75t_SL g96 ( 
.A(n_63),
.Y(n_96)
);

AOI22xp33_ASAP7_75t_SL g115 ( 
.A1(n_96),
.A2(n_77),
.B1(n_78),
.B2(n_80),
.Y(n_115)
);

AND2x6_ASAP7_75t_L g97 ( 
.A(n_76),
.B(n_38),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_SL g111 ( 
.A(n_97),
.B(n_100),
.Y(n_111)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_80),
.Y(n_98)
);

CKINVDCx16_ASAP7_75t_R g122 ( 
.A(n_98),
.Y(n_122)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_80),
.Y(n_99)
);

CKINVDCx20_ASAP7_75t_R g107 ( 
.A(n_99),
.Y(n_107)
);

CKINVDCx20_ASAP7_75t_R g100 ( 
.A(n_78),
.Y(n_100)
);

MAJx2_ASAP7_75t_L g101 ( 
.A(n_88),
.B(n_64),
.C(n_68),
.Y(n_101)
);

OAI21xp5_ASAP7_75t_L g148 ( 
.A1(n_101),
.A2(n_105),
.B(n_108),
.Y(n_148)
);

INVx2_ASAP7_75t_L g102 ( 
.A(n_84),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_L g137 ( 
.A(n_102),
.B(n_93),
.Y(n_137)
);

INVxp67_ASAP7_75t_L g103 ( 
.A(n_88),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_SL g153 ( 
.A(n_103),
.B(n_59),
.Y(n_153)
);

OAI21xp5_ASAP7_75t_L g105 ( 
.A1(n_82),
.A2(n_68),
.B(n_69),
.Y(n_105)
);

OAI22xp5_ASAP7_75t_SL g150 ( 
.A1(n_106),
.A2(n_125),
.B1(n_14),
.B2(n_17),
.Y(n_150)
);

OAI21xp5_ASAP7_75t_L g108 ( 
.A1(n_82),
.A2(n_68),
.B(n_71),
.Y(n_108)
);

MAJIxp5_ASAP7_75t_L g109 ( 
.A(n_81),
.B(n_73),
.C(n_72),
.Y(n_109)
);

MAJIxp5_ASAP7_75t_L g126 ( 
.A(n_109),
.B(n_113),
.C(n_114),
.Y(n_126)
);

MAJIxp5_ASAP7_75t_L g113 ( 
.A(n_81),
.B(n_72),
.C(n_62),
.Y(n_113)
);

MAJIxp5_ASAP7_75t_L g114 ( 
.A(n_95),
.B(n_72),
.C(n_29),
.Y(n_114)
);

INVxp67_ASAP7_75t_L g149 ( 
.A(n_115),
.Y(n_149)
);

NOR2x1_ASAP7_75t_L g117 ( 
.A(n_97),
.B(n_72),
.Y(n_117)
);

OR2x2_ASAP7_75t_L g130 ( 
.A(n_117),
.B(n_86),
.Y(n_130)
);

AND2x2_ASAP7_75t_L g120 ( 
.A(n_97),
.B(n_59),
.Y(n_120)
);

AOI21xp5_ASAP7_75t_L g135 ( 
.A1(n_120),
.A2(n_99),
.B(n_98),
.Y(n_135)
);

OAI22xp5_ASAP7_75t_SL g121 ( 
.A1(n_86),
.A2(n_50),
.B1(n_17),
.B2(n_23),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_L g131 ( 
.A(n_121),
.B(n_123),
.Y(n_131)
);

AO22x1_ASAP7_75t_SL g123 ( 
.A1(n_86),
.A2(n_91),
.B1(n_94),
.B2(n_95),
.Y(n_123)
);

AOI22xp5_ASAP7_75t_L g125 ( 
.A1(n_85),
.A2(n_77),
.B1(n_18),
.B2(n_50),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_L g127 ( 
.A(n_110),
.B(n_100),
.Y(n_127)
);

CKINVDCx14_ASAP7_75t_R g164 ( 
.A(n_127),
.Y(n_164)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_110),
.B(n_92),
.Y(n_128)
);

CKINVDCx14_ASAP7_75t_R g165 ( 
.A(n_128),
.Y(n_165)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_118),
.Y(n_129)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_129),
.Y(n_172)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_130),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_L g132 ( 
.A(n_109),
.B(n_83),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_L g160 ( 
.A(n_132),
.B(n_133),
.Y(n_160)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_118),
.Y(n_133)
);

MAJIxp5_ASAP7_75t_L g134 ( 
.A(n_108),
.B(n_87),
.C(n_89),
.Y(n_134)
);

MAJIxp5_ASAP7_75t_L g171 ( 
.A(n_134),
.B(n_114),
.C(n_120),
.Y(n_171)
);

OAI21xp5_ASAP7_75t_L g168 ( 
.A1(n_135),
.A2(n_140),
.B(n_153),
.Y(n_168)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_124),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_L g174 ( 
.A(n_136),
.B(n_138),
.Y(n_174)
);

CKINVDCx20_ASAP7_75t_R g159 ( 
.A(n_137),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_L g138 ( 
.A(n_113),
.B(n_96),
.Y(n_138)
);

CKINVDCx16_ASAP7_75t_R g139 ( 
.A(n_112),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_SL g169 ( 
.A(n_139),
.B(n_154),
.Y(n_169)
);

AND2x2_ASAP7_75t_L g140 ( 
.A(n_111),
.B(n_59),
.Y(n_140)
);

CKINVDCx20_ASAP7_75t_R g141 ( 
.A(n_112),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_L g184 ( 
.A(n_141),
.B(n_143),
.Y(n_184)
);

BUFx24_ASAP7_75t_SL g142 ( 
.A(n_104),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_L g175 ( 
.A(n_142),
.B(n_122),
.Y(n_175)
);

AND2x2_ASAP7_75t_SL g143 ( 
.A(n_121),
.B(n_45),
.Y(n_143)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_124),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_L g186 ( 
.A(n_144),
.B(n_146),
.Y(n_186)
);

NOR2xp33_ASAP7_75t_L g145 ( 
.A(n_107),
.B(n_96),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_SL g173 ( 
.A(n_145),
.B(n_157),
.Y(n_173)
);

OR2x2_ASAP7_75t_L g146 ( 
.A(n_123),
.B(n_22),
.Y(n_146)
);

BUFx3_ASAP7_75t_L g147 ( 
.A(n_103),
.Y(n_147)
);

INVx2_ASAP7_75t_L g170 ( 
.A(n_147),
.Y(n_170)
);

AOI22xp5_ASAP7_75t_L g163 ( 
.A1(n_150),
.A2(n_152),
.B1(n_122),
.B2(n_117),
.Y(n_163)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_116),
.Y(n_151)
);

CKINVDCx20_ASAP7_75t_R g185 ( 
.A(n_151),
.Y(n_185)
);

OAI22xp5_ASAP7_75t_L g152 ( 
.A1(n_106),
.A2(n_18),
.B1(n_23),
.B2(n_21),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_L g154 ( 
.A(n_125),
.B(n_63),
.Y(n_154)
);

NOR2xp33_ASAP7_75t_L g155 ( 
.A(n_119),
.B(n_63),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_SL g181 ( 
.A(n_155),
.B(n_59),
.Y(n_181)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_116),
.Y(n_156)
);

CKINVDCx16_ASAP7_75t_R g166 ( 
.A(n_156),
.Y(n_166)
);

NOR2xp33_ASAP7_75t_L g157 ( 
.A(n_107),
.B(n_13),
.Y(n_157)
);

OAI21xp5_ASAP7_75t_L g158 ( 
.A1(n_101),
.A2(n_22),
.B(n_19),
.Y(n_158)
);

XOR2xp5_ASAP7_75t_L g182 ( 
.A(n_158),
.B(n_47),
.Y(n_182)
);

NAND2xp33_ASAP7_75t_SL g161 ( 
.A(n_143),
.B(n_117),
.Y(n_161)
);

AOI21xp5_ASAP7_75t_SL g188 ( 
.A1(n_161),
.A2(n_167),
.B(n_135),
.Y(n_188)
);

XNOR2xp5_ASAP7_75t_L g162 ( 
.A(n_148),
.B(n_105),
.Y(n_162)
);

XNOR2xp5_ASAP7_75t_L g210 ( 
.A(n_162),
.B(n_129),
.Y(n_210)
);

OAI22xp5_ASAP7_75t_L g194 ( 
.A1(n_163),
.A2(n_178),
.B1(n_180),
.B2(n_141),
.Y(n_194)
);

NAND2xp33_ASAP7_75t_SL g167 ( 
.A(n_143),
.B(n_120),
.Y(n_167)
);

MAJIxp5_ASAP7_75t_L g195 ( 
.A(n_171),
.B(n_126),
.C(n_132),
.Y(n_195)
);

NOR2xp33_ASAP7_75t_SL g191 ( 
.A(n_175),
.B(n_158),
.Y(n_191)
);

NOR2xp33_ASAP7_75t_L g177 ( 
.A(n_134),
.B(n_102),
.Y(n_177)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_177),
.Y(n_190)
);

AOI22xp5_ASAP7_75t_L g178 ( 
.A1(n_131),
.A2(n_123),
.B1(n_18),
.B2(n_21),
.Y(n_178)
);

OAI22xp5_ASAP7_75t_L g179 ( 
.A1(n_146),
.A2(n_14),
.B1(n_23),
.B2(n_17),
.Y(n_179)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_179),
.Y(n_202)
);

AOI22xp5_ASAP7_75t_L g180 ( 
.A1(n_131),
.A2(n_14),
.B1(n_23),
.B2(n_2),
.Y(n_180)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_181),
.Y(n_207)
);

FAx1_ASAP7_75t_SL g204 ( 
.A(n_182),
.B(n_140),
.CI(n_145),
.CON(n_204),
.SN(n_204)
);

O2A1O1Ixp33_ASAP7_75t_L g183 ( 
.A1(n_146),
.A2(n_14),
.B(n_47),
.C(n_45),
.Y(n_183)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_183),
.Y(n_189)
);

BUFx5_ASAP7_75t_L g187 ( 
.A(n_153),
.Y(n_187)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_187),
.Y(n_192)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_188),
.Y(n_217)
);

NAND2xp5_ASAP7_75t_SL g213 ( 
.A(n_191),
.B(n_196),
.Y(n_213)
);

AO22x1_ASAP7_75t_SL g193 ( 
.A1(n_161),
.A2(n_130),
.B1(n_143),
.B2(n_150),
.Y(n_193)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_193),
.Y(n_219)
);

CKINVDCx16_ASAP7_75t_R g215 ( 
.A(n_194),
.Y(n_215)
);

MAJIxp5_ASAP7_75t_L g221 ( 
.A(n_195),
.B(n_208),
.C(n_210),
.Y(n_221)
);

NOR2xp33_ASAP7_75t_SL g196 ( 
.A(n_165),
.B(n_148),
.Y(n_196)
);

OAI22xp5_ASAP7_75t_L g197 ( 
.A1(n_164),
.A2(n_170),
.B1(n_186),
.B2(n_149),
.Y(n_197)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_197),
.Y(n_224)
);

OAI22xp5_ASAP7_75t_L g198 ( 
.A1(n_170),
.A2(n_130),
.B1(n_138),
.B2(n_126),
.Y(n_198)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_198),
.Y(n_225)
);

NOR2xp33_ASAP7_75t_L g199 ( 
.A(n_173),
.B(n_159),
.Y(n_199)
);

NOR2xp33_ASAP7_75t_L g229 ( 
.A(n_199),
.B(n_201),
.Y(n_229)
);

INVxp67_ASAP7_75t_L g200 ( 
.A(n_174),
.Y(n_200)
);

OAI22xp5_ASAP7_75t_SL g218 ( 
.A1(n_200),
.A2(n_159),
.B1(n_186),
.B2(n_176),
.Y(n_218)
);

NOR2xp33_ASAP7_75t_L g201 ( 
.A(n_173),
.B(n_147),
.Y(n_201)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_174),
.Y(n_203)
);

OAI22xp5_ASAP7_75t_L g214 ( 
.A1(n_203),
.A2(n_205),
.B1(n_206),
.B2(n_211),
.Y(n_214)
);

XNOR2xp5_ASAP7_75t_L g233 ( 
.A(n_204),
.B(n_212),
.Y(n_233)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_184),
.Y(n_205)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_184),
.Y(n_206)
);

MAJIxp5_ASAP7_75t_L g208 ( 
.A(n_171),
.B(n_140),
.C(n_156),
.Y(n_208)
);

NOR2xp33_ASAP7_75t_SL g209 ( 
.A(n_162),
.B(n_136),
.Y(n_209)
);

NOR3xp33_ASAP7_75t_L g231 ( 
.A(n_209),
.B(n_189),
.C(n_202),
.Y(n_231)
);

XNOR2xp5_ASAP7_75t_SL g220 ( 
.A(n_210),
.B(n_182),
.Y(n_220)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_160),
.Y(n_211)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_160),
.Y(n_212)
);

OAI22xp5_ASAP7_75t_SL g226 ( 
.A1(n_212),
.A2(n_176),
.B1(n_185),
.B2(n_178),
.Y(n_226)
);

INVx4_ASAP7_75t_L g216 ( 
.A(n_207),
.Y(n_216)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_216),
.Y(n_239)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_218),
.Y(n_242)
);

XNOR2xp5_ASAP7_75t_L g250 ( 
.A(n_220),
.B(n_222),
.Y(n_250)
);

MAJIxp5_ASAP7_75t_L g237 ( 
.A(n_221),
.B(n_223),
.C(n_230),
.Y(n_237)
);

XOR2xp5_ASAP7_75t_L g222 ( 
.A(n_195),
.B(n_168),
.Y(n_222)
);

MAJIxp5_ASAP7_75t_L g223 ( 
.A(n_208),
.B(n_168),
.C(n_163),
.Y(n_223)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_226),
.Y(n_246)
);

XNOR2xp5_ASAP7_75t_SL g227 ( 
.A(n_204),
.B(n_167),
.Y(n_227)
);

AOI22xp5_ASAP7_75t_SL g245 ( 
.A1(n_227),
.A2(n_205),
.B1(n_193),
.B2(n_144),
.Y(n_245)
);

OAI22xp5_ASAP7_75t_SL g228 ( 
.A1(n_203),
.A2(n_185),
.B1(n_180),
.B2(n_183),
.Y(n_228)
);

AOI22xp5_ASAP7_75t_L g235 ( 
.A1(n_228),
.A2(n_234),
.B1(n_200),
.B2(n_211),
.Y(n_235)
);

MAJIxp5_ASAP7_75t_L g230 ( 
.A(n_190),
.B(n_172),
.C(n_151),
.Y(n_230)
);

NOR2xp33_ASAP7_75t_L g241 ( 
.A(n_231),
.B(n_192),
.Y(n_241)
);

XOR2xp5_ASAP7_75t_L g232 ( 
.A(n_188),
.B(n_187),
.Y(n_232)
);

MAJIxp5_ASAP7_75t_L g243 ( 
.A(n_232),
.B(n_192),
.C(n_206),
.Y(n_243)
);

NAND2xp5_ASAP7_75t_L g238 ( 
.A(n_233),
.B(n_204),
.Y(n_238)
);

OAI22xp5_ASAP7_75t_SL g234 ( 
.A1(n_189),
.A2(n_169),
.B1(n_172),
.B2(n_166),
.Y(n_234)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_235),
.Y(n_253)
);

INVxp67_ASAP7_75t_L g236 ( 
.A(n_229),
.Y(n_236)
);

NAND2xp5_ASAP7_75t_L g265 ( 
.A(n_236),
.B(n_238),
.Y(n_265)
);

INVx13_ASAP7_75t_L g240 ( 
.A(n_216),
.Y(n_240)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_240),
.Y(n_254)
);

AOI21xp5_ASAP7_75t_L g256 ( 
.A1(n_241),
.A2(n_233),
.B(n_224),
.Y(n_256)
);

XOR2xp5_ASAP7_75t_L g257 ( 
.A(n_243),
.B(n_222),
.Y(n_257)
);

NOR2xp33_ASAP7_75t_L g244 ( 
.A(n_230),
.B(n_139),
.Y(n_244)
);

NOR2xp33_ASAP7_75t_L g262 ( 
.A(n_244),
.B(n_248),
.Y(n_262)
);

XNOR2xp5_ASAP7_75t_SL g264 ( 
.A(n_245),
.B(n_243),
.Y(n_264)
);

MAJIxp5_ASAP7_75t_L g247 ( 
.A(n_221),
.B(n_133),
.C(n_137),
.Y(n_247)
);

MAJIxp5_ASAP7_75t_L g259 ( 
.A(n_247),
.B(n_220),
.C(n_227),
.Y(n_259)
);

NAND2xp5_ASAP7_75t_L g248 ( 
.A(n_213),
.B(n_193),
.Y(n_248)
);

BUFx12_ASAP7_75t_L g249 ( 
.A(n_232),
.Y(n_249)
);

XNOR2xp5_ASAP7_75t_L g261 ( 
.A(n_249),
.B(n_47),
.Y(n_261)
);

MAJIxp5_ASAP7_75t_L g251 ( 
.A(n_225),
.B(n_157),
.C(n_152),
.Y(n_251)
);

MAJIxp5_ASAP7_75t_L g267 ( 
.A(n_251),
.B(n_252),
.C(n_13),
.Y(n_267)
);

MAJIxp5_ASAP7_75t_L g252 ( 
.A(n_223),
.B(n_47),
.C(n_13),
.Y(n_252)
);

OAI21xp33_ASAP7_75t_L g255 ( 
.A1(n_242),
.A2(n_217),
.B(n_219),
.Y(n_255)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_255),
.Y(n_270)
);

CKINVDCx20_ASAP7_75t_R g279 ( 
.A(n_256),
.Y(n_279)
);

NAND2xp5_ASAP7_75t_SL g277 ( 
.A(n_257),
.B(n_259),
.Y(n_277)
);

AOI22xp5_ASAP7_75t_L g258 ( 
.A1(n_246),
.A2(n_215),
.B1(n_218),
.B2(n_214),
.Y(n_258)
);

NAND2xp5_ASAP7_75t_L g269 ( 
.A(n_258),
.B(n_260),
.Y(n_269)
);

OAI22xp5_ASAP7_75t_SL g260 ( 
.A1(n_236),
.A2(n_228),
.B1(n_38),
.B2(n_7),
.Y(n_260)
);

AND2x2_ASAP7_75t_L g271 ( 
.A(n_261),
.B(n_252),
.Y(n_271)
);

AOI22xp33_ASAP7_75t_SL g263 ( 
.A1(n_239),
.A2(n_38),
.B1(n_10),
.B2(n_9),
.Y(n_263)
);

INVxp67_ASAP7_75t_L g268 ( 
.A(n_263),
.Y(n_268)
);

MAJIxp5_ASAP7_75t_L g272 ( 
.A(n_264),
.B(n_237),
.C(n_247),
.Y(n_272)
);

XNOR2xp5_ASAP7_75t_L g266 ( 
.A(n_237),
.B(n_13),
.Y(n_266)
);

NAND2xp5_ASAP7_75t_SL g280 ( 
.A(n_266),
.B(n_267),
.Y(n_280)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_271),
.Y(n_286)
);

AND2x2_ASAP7_75t_L g291 ( 
.A(n_272),
.B(n_0),
.Y(n_291)
);

MAJIxp5_ASAP7_75t_L g273 ( 
.A(n_257),
.B(n_250),
.C(n_251),
.Y(n_273)
);

OR2x2_ASAP7_75t_L g285 ( 
.A(n_273),
.B(n_276),
.Y(n_285)
);

NOR2xp33_ASAP7_75t_L g274 ( 
.A(n_262),
.B(n_240),
.Y(n_274)
);

NAND2xp5_ASAP7_75t_L g282 ( 
.A(n_274),
.B(n_275),
.Y(n_282)
);

OAI21xp5_ASAP7_75t_SL g275 ( 
.A1(n_265),
.A2(n_249),
.B(n_9),
.Y(n_275)
);

NOR2xp33_ASAP7_75t_L g276 ( 
.A(n_254),
.B(n_249),
.Y(n_276)
);

OR2x2_ASAP7_75t_L g278 ( 
.A(n_255),
.B(n_8),
.Y(n_278)
);

NAND2xp5_ASAP7_75t_SL g288 ( 
.A(n_278),
.B(n_7),
.Y(n_288)
);

OAI21x1_ASAP7_75t_L g281 ( 
.A1(n_277),
.A2(n_264),
.B(n_259),
.Y(n_281)
);

AOI322xp5_ASAP7_75t_L g300 ( 
.A1(n_281),
.A2(n_290),
.A3(n_292),
.B1(n_3),
.B2(n_4),
.C1(n_5),
.C2(n_6),
.Y(n_300)
);

NOR2xp33_ASAP7_75t_L g283 ( 
.A(n_269),
.B(n_253),
.Y(n_283)
);

NAND2xp5_ASAP7_75t_L g296 ( 
.A(n_283),
.B(n_284),
.Y(n_296)
);

XNOR2xp5_ASAP7_75t_L g284 ( 
.A(n_280),
.B(n_267),
.Y(n_284)
);

XOR2xp5_ASAP7_75t_L g287 ( 
.A(n_271),
.B(n_263),
.Y(n_287)
);

NAND2xp5_ASAP7_75t_SL g298 ( 
.A(n_287),
.B(n_291),
.Y(n_298)
);

NAND2xp5_ASAP7_75t_L g299 ( 
.A(n_288),
.B(n_289),
.Y(n_299)
);

NOR2xp33_ASAP7_75t_L g289 ( 
.A(n_279),
.B(n_7),
.Y(n_289)
);

OAI21xp5_ASAP7_75t_L g290 ( 
.A1(n_270),
.A2(n_0),
.B(n_1),
.Y(n_290)
);

HB1xp67_ASAP7_75t_L g292 ( 
.A(n_268),
.Y(n_292)
);

MAJIxp5_ASAP7_75t_L g293 ( 
.A(n_285),
.B(n_278),
.C(n_268),
.Y(n_293)
);

HB1xp67_ASAP7_75t_L g303 ( 
.A(n_293),
.Y(n_303)
);

OAI21x1_ASAP7_75t_L g294 ( 
.A1(n_286),
.A2(n_0),
.B(n_1),
.Y(n_294)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_294),
.Y(n_301)
);

A2O1A1Ixp33_ASAP7_75t_SL g295 ( 
.A1(n_282),
.A2(n_0),
.B(n_1),
.C(n_2),
.Y(n_295)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_295),
.Y(n_302)
);

MAJIxp5_ASAP7_75t_L g297 ( 
.A(n_283),
.B(n_2),
.C(n_3),
.Y(n_297)
);

AOI21xp5_ASAP7_75t_L g304 ( 
.A1(n_297),
.A2(n_300),
.B(n_288),
.Y(n_304)
);

CKINVDCx20_ASAP7_75t_R g306 ( 
.A(n_304),
.Y(n_306)
);

AOI322xp5_ASAP7_75t_L g305 ( 
.A1(n_302),
.A2(n_298),
.A3(n_301),
.B1(n_303),
.B2(n_296),
.C1(n_295),
.C2(n_299),
.Y(n_305)
);

OAI21xp5_ASAP7_75t_SL g307 ( 
.A1(n_305),
.A2(n_3),
.B(n_4),
.Y(n_307)
);

MAJIxp5_ASAP7_75t_L g308 ( 
.A(n_307),
.B(n_306),
.C(n_4),
.Y(n_308)
);

NOR3xp33_ASAP7_75t_L g309 ( 
.A(n_308),
.B(n_3),
.C(n_5),
.Y(n_309)
);

OAI22xp5_ASAP7_75t_L g310 ( 
.A1(n_309),
.A2(n_3),
.B1(n_5),
.B2(n_6),
.Y(n_310)
);

MAJIxp5_ASAP7_75t_L g311 ( 
.A(n_310),
.B(n_5),
.C(n_293),
.Y(n_311)
);


endmodule