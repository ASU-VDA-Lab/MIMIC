module fake_jpeg_25042_n_116 (n_3, n_2, n_1, n_0, n_4, n_8, n_6, n_5, n_7, n_116);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_8;
input n_6;
input n_5;
input n_7;

output n_116;

wire n_10;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_114;
wire n_74;
wire n_31;
wire n_29;
wire n_103;
wire n_50;
wire n_15;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_109;
wire n_113;
wire n_30;
wire n_106;
wire n_111;
wire n_24;
wire n_44;
wire n_17;
wire n_25;
wire n_75;
wire n_37;
wire n_102;
wire n_99;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_18;
wire n_20;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_11;
wire n_56;
wire n_79;
wire n_12;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_22;
wire n_101;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_112;
wire n_95;
wire n_97;
wire n_9;
wire n_36;
wire n_62;
wire n_43;
wire n_32;
wire n_100;
wire n_82;
wire n_96;

CKINVDCx20_ASAP7_75t_R g9 ( 
.A(n_2),
.Y(n_9)
);

INVx1_ASAP7_75t_L g10 ( 
.A(n_1),
.Y(n_10)
);

INVx6_ASAP7_75t_L g11 ( 
.A(n_1),
.Y(n_11)
);

INVx3_ASAP7_75t_L g12 ( 
.A(n_2),
.Y(n_12)
);

INVx1_ASAP7_75t_L g13 ( 
.A(n_5),
.Y(n_13)
);

INVx1_ASAP7_75t_L g14 ( 
.A(n_5),
.Y(n_14)
);

BUFx12f_ASAP7_75t_L g15 ( 
.A(n_2),
.Y(n_15)
);

INVx2_ASAP7_75t_L g16 ( 
.A(n_1),
.Y(n_16)
);

INVx5_ASAP7_75t_L g17 ( 
.A(n_8),
.Y(n_17)
);

INVx2_ASAP7_75t_L g18 ( 
.A(n_16),
.Y(n_18)
);

INVx2_ASAP7_75t_L g32 ( 
.A(n_18),
.Y(n_32)
);

INVx3_ASAP7_75t_L g19 ( 
.A(n_15),
.Y(n_19)
);

INVx5_ASAP7_75t_L g26 ( 
.A(n_19),
.Y(n_26)
);

INVx6_ASAP7_75t_L g20 ( 
.A(n_15),
.Y(n_20)
);

AOI22xp33_ASAP7_75t_SL g33 ( 
.A1(n_20),
.A2(n_17),
.B1(n_9),
.B2(n_10),
.Y(n_33)
);

INVx3_ASAP7_75t_L g21 ( 
.A(n_15),
.Y(n_21)
);

BUFx3_ASAP7_75t_L g29 ( 
.A(n_21),
.Y(n_29)
);

INVx2_ASAP7_75t_L g22 ( 
.A(n_16),
.Y(n_22)
);

OR2x2_ASAP7_75t_L g30 ( 
.A(n_22),
.B(n_23),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_15),
.Y(n_23)
);

BUFx4f_ASAP7_75t_L g24 ( 
.A(n_11),
.Y(n_24)
);

INVx8_ASAP7_75t_L g31 ( 
.A(n_24),
.Y(n_31)
);

OA22x2_ASAP7_75t_L g25 ( 
.A1(n_19),
.A2(n_11),
.B1(n_12),
.B2(n_17),
.Y(n_25)
);

OAI22xp5_ASAP7_75t_SL g35 ( 
.A1(n_25),
.A2(n_28),
.B1(n_21),
.B2(n_10),
.Y(n_35)
);

NAND2xp5_ASAP7_75t_L g27 ( 
.A(n_22),
.B(n_12),
.Y(n_27)
);

NAND2xp5_ASAP7_75t_L g36 ( 
.A(n_27),
.B(n_32),
.Y(n_36)
);

AOI22xp33_ASAP7_75t_SL g28 ( 
.A1(n_20),
.A2(n_11),
.B1(n_17),
.B2(n_9),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_33),
.Y(n_37)
);

NAND2xp5_ASAP7_75t_SL g34 ( 
.A(n_27),
.B(n_24),
.Y(n_34)
);

NAND2xp5_ASAP7_75t_L g49 ( 
.A(n_34),
.B(n_36),
.Y(n_49)
);

OAI22xp5_ASAP7_75t_L g43 ( 
.A1(n_35),
.A2(n_28),
.B1(n_33),
.B2(n_25),
.Y(n_43)
);

BUFx3_ASAP7_75t_L g38 ( 
.A(n_32),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_L g46 ( 
.A(n_38),
.B(n_42),
.Y(n_46)
);

AND2x2_ASAP7_75t_L g39 ( 
.A(n_27),
.B(n_24),
.Y(n_39)
);

MAJIxp5_ASAP7_75t_SL g45 ( 
.A(n_39),
.B(n_30),
.C(n_25),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g40 ( 
.A(n_30),
.B(n_14),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g47 ( 
.A(n_40),
.B(n_41),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g41 ( 
.A(n_30),
.B(n_14),
.Y(n_41)
);

NAND2xp5_ASAP7_75t_L g42 ( 
.A(n_30),
.B(n_23),
.Y(n_42)
);

AOI22xp5_ASAP7_75t_L g53 ( 
.A1(n_43),
.A2(n_44),
.B1(n_35),
.B2(n_37),
.Y(n_53)
);

OAI22xp33_ASAP7_75t_SL g44 ( 
.A1(n_37),
.A2(n_25),
.B1(n_31),
.B2(n_32),
.Y(n_44)
);

NAND2xp5_ASAP7_75t_SL g55 ( 
.A(n_45),
.B(n_50),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_40),
.B(n_29),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g57 ( 
.A(n_48),
.B(n_52),
.Y(n_57)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_36),
.Y(n_50)
);

INVxp33_ASAP7_75t_SL g51 ( 
.A(n_38),
.Y(n_51)
);

INVx1_ASAP7_75t_SL g56 ( 
.A(n_51),
.Y(n_56)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_42),
.Y(n_52)
);

OAI22xp5_ASAP7_75t_L g70 ( 
.A1(n_53),
.A2(n_59),
.B1(n_26),
.B2(n_29),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_L g54 ( 
.A(n_49),
.B(n_34),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_L g71 ( 
.A(n_54),
.B(n_62),
.Y(n_71)
);

OAI22xp5_ASAP7_75t_SL g58 ( 
.A1(n_43),
.A2(n_30),
.B1(n_39),
.B2(n_31),
.Y(n_58)
);

AOI22xp5_ASAP7_75t_L g65 ( 
.A1(n_58),
.A2(n_62),
.B1(n_25),
.B2(n_26),
.Y(n_65)
);

AOI22xp5_ASAP7_75t_L g59 ( 
.A1(n_52),
.A2(n_39),
.B1(n_41),
.B2(n_31),
.Y(n_59)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_46),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_SL g63 ( 
.A(n_60),
.B(n_47),
.Y(n_63)
);

MAJIxp5_ASAP7_75t_L g61 ( 
.A(n_50),
.B(n_31),
.C(n_25),
.Y(n_61)
);

XNOR2xp5_ASAP7_75t_L g68 ( 
.A(n_61),
.B(n_29),
.Y(n_68)
);

OAI22xp5_ASAP7_75t_SL g62 ( 
.A1(n_49),
.A2(n_45),
.B1(n_47),
.B2(n_25),
.Y(n_62)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_63),
.Y(n_78)
);

INVx4_ASAP7_75t_L g64 ( 
.A(n_56),
.Y(n_64)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_64),
.Y(n_79)
);

OAI22xp5_ASAP7_75t_SL g82 ( 
.A1(n_65),
.A2(n_29),
.B1(n_13),
.B2(n_2),
.Y(n_82)
);

INVxp67_ASAP7_75t_L g66 ( 
.A(n_57),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_L g81 ( 
.A(n_66),
.B(n_70),
.Y(n_81)
);

OAI21xp5_ASAP7_75t_L g67 ( 
.A1(n_55),
.A2(n_13),
.B(n_25),
.Y(n_67)
);

AOI21xp5_ASAP7_75t_L g75 ( 
.A1(n_67),
.A2(n_55),
.B(n_54),
.Y(n_75)
);

MAJIxp5_ASAP7_75t_L g76 ( 
.A(n_68),
.B(n_61),
.C(n_26),
.Y(n_76)
);

CKINVDCx16_ASAP7_75t_R g69 ( 
.A(n_56),
.Y(n_69)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_69),
.Y(n_77)
);

INVx1_ASAP7_75t_SL g74 ( 
.A(n_71),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_60),
.B(n_26),
.Y(n_72)
);

CKINVDCx20_ASAP7_75t_R g80 ( 
.A(n_72),
.Y(n_80)
);

AOI22xp5_ASAP7_75t_SL g73 ( 
.A1(n_66),
.A2(n_58),
.B1(n_53),
.B2(n_59),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_73),
.B(n_70),
.Y(n_84)
);

XNOR2xp5_ASAP7_75t_SL g83 ( 
.A(n_75),
.B(n_67),
.Y(n_83)
);

MAJIxp5_ASAP7_75t_L g88 ( 
.A(n_76),
.B(n_68),
.C(n_65),
.Y(n_88)
);

AOI22xp5_ASAP7_75t_L g86 ( 
.A1(n_82),
.A2(n_64),
.B1(n_1),
.B2(n_3),
.Y(n_86)
);

XNOR2xp5_ASAP7_75t_SL g92 ( 
.A(n_83),
.B(n_75),
.Y(n_92)
);

AOI22xp5_ASAP7_75t_L g94 ( 
.A1(n_84),
.A2(n_86),
.B1(n_79),
.B2(n_74),
.Y(n_94)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_81),
.Y(n_85)
);

AOI21xp5_ASAP7_75t_L g96 ( 
.A1(n_85),
.A2(n_87),
.B(n_89),
.Y(n_96)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_81),
.Y(n_87)
);

XOR2xp5_ASAP7_75t_L g93 ( 
.A(n_88),
.B(n_90),
.Y(n_93)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_82),
.Y(n_89)
);

MAJIxp5_ASAP7_75t_L g90 ( 
.A(n_76),
.B(n_71),
.C(n_6),
.Y(n_90)
);

CKINVDCx20_ASAP7_75t_R g91 ( 
.A(n_80),
.Y(n_91)
);

INVx3_ASAP7_75t_L g98 ( 
.A(n_91),
.Y(n_98)
);

XOR2xp5_ASAP7_75t_L g100 ( 
.A(n_92),
.B(n_97),
.Y(n_100)
);

OR2x2_ASAP7_75t_L g103 ( 
.A(n_94),
.B(n_4),
.Y(n_103)
);

AOI321xp33_ASAP7_75t_L g95 ( 
.A1(n_83),
.A2(n_78),
.A3(n_73),
.B1(n_74),
.B2(n_77),
.C(n_6),
.Y(n_95)
);

AOI21xp5_ASAP7_75t_L g101 ( 
.A1(n_95),
.A2(n_7),
.B(n_8),
.Y(n_101)
);

XNOR2xp5_ASAP7_75t_SL g97 ( 
.A(n_90),
.B(n_88),
.Y(n_97)
);

AOI22xp5_ASAP7_75t_L g99 ( 
.A1(n_98),
.A2(n_77),
.B1(n_6),
.B2(n_4),
.Y(n_99)
);

MAJIxp5_ASAP7_75t_L g106 ( 
.A(n_99),
.B(n_102),
.C(n_0),
.Y(n_106)
);

OAI21xp5_ASAP7_75t_SL g104 ( 
.A1(n_101),
.A2(n_96),
.B(n_7),
.Y(n_104)
);

MAJIxp5_ASAP7_75t_L g102 ( 
.A(n_93),
.B(n_4),
.C(n_5),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_SL g107 ( 
.A(n_103),
.B(n_0),
.Y(n_107)
);

XNOR2xp5_ASAP7_75t_L g108 ( 
.A(n_104),
.B(n_105),
.Y(n_108)
);

AOI22xp5_ASAP7_75t_SL g105 ( 
.A1(n_100),
.A2(n_92),
.B1(n_7),
.B2(n_8),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_SL g110 ( 
.A(n_106),
.B(n_107),
.Y(n_110)
);

XNOR2xp5_ASAP7_75t_L g109 ( 
.A(n_105),
.B(n_100),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_L g111 ( 
.A(n_109),
.B(n_103),
.Y(n_111)
);

INVxp67_ASAP7_75t_L g113 ( 
.A(n_111),
.Y(n_113)
);

AOI22xp5_ASAP7_75t_SL g112 ( 
.A1(n_108),
.A2(n_0),
.B1(n_3),
.B2(n_110),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_L g114 ( 
.A(n_113),
.B(n_112),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_SL g115 ( 
.A(n_114),
.B(n_0),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_L g116 ( 
.A(n_115),
.B(n_3),
.Y(n_116)
);


endmodule