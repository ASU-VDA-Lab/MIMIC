module fake_jpeg_19760_n_79 (n_13, n_21, n_1, n_10, n_6, n_22, n_14, n_19, n_18, n_20, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_79);

input n_13;
input n_21;
input n_1;
input n_10;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_79;

wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_73;
wire n_59;
wire n_65;
wire n_42;
wire n_49;
wire n_76;
wire n_28;
wire n_38;
wire n_26;
wire n_74;
wire n_31;
wire n_29;
wire n_50;
wire n_57;
wire n_23;
wire n_69;
wire n_27;
wire n_40;
wire n_71;
wire n_30;
wire n_24;
wire n_44;
wire n_25;
wire n_75;
wire n_37;
wire n_70;
wire n_66;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_68;
wire n_52;
wire n_58;
wire n_41;
wire n_60;
wire n_63;
wire n_34;
wire n_39;
wire n_72;
wire n_56;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_35;
wire n_48;
wire n_46;
wire n_36;
wire n_62;
wire n_43;
wire n_32;

INVx1_ASAP7_75t_L g23 ( 
.A(n_0),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_3),
.Y(n_24)
);

INVx8_ASAP7_75t_L g25 ( 
.A(n_4),
.Y(n_25)
);

BUFx6f_ASAP7_75t_SL g26 ( 
.A(n_22),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_2),
.Y(n_27)
);

BUFx3_ASAP7_75t_L g28 ( 
.A(n_2),
.Y(n_28)
);

INVx13_ASAP7_75t_L g29 ( 
.A(n_15),
.Y(n_29)
);

BUFx12_ASAP7_75t_L g30 ( 
.A(n_12),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_3),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_17),
.Y(n_32)
);

BUFx12_ASAP7_75t_L g33 ( 
.A(n_16),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_20),
.Y(n_34)
);

INVx2_ASAP7_75t_L g35 ( 
.A(n_5),
.Y(n_35)
);

INVx8_ASAP7_75t_L g36 ( 
.A(n_7),
.Y(n_36)
);

NAND2xp5_ASAP7_75t_L g37 ( 
.A(n_8),
.B(n_19),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_9),
.Y(n_38)
);

BUFx3_ASAP7_75t_L g39 ( 
.A(n_11),
.Y(n_39)
);

BUFx4f_ASAP7_75t_SL g40 ( 
.A(n_18),
.Y(n_40)
);

CKINVDCx14_ASAP7_75t_R g41 ( 
.A(n_5),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_4),
.Y(n_42)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_1),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_14),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_21),
.Y(n_45)
);

BUFx4f_ASAP7_75t_SL g46 ( 
.A(n_1),
.Y(n_46)
);

BUFx12f_ASAP7_75t_L g47 ( 
.A(n_39),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_47),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_35),
.B(n_6),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_SL g58 ( 
.A(n_48),
.B(n_51),
.Y(n_58)
);

INVx2_ASAP7_75t_L g49 ( 
.A(n_28),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_49),
.B(n_50),
.Y(n_59)
);

INVx6_ASAP7_75t_L g50 ( 
.A(n_35),
.Y(n_50)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_26),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_37),
.B(n_10),
.Y(n_52)
);

INVx11_ASAP7_75t_L g53 ( 
.A(n_30),
.Y(n_53)
);

AOI22xp33_ASAP7_75t_L g54 ( 
.A1(n_36),
.A2(n_13),
.B1(n_25),
.B2(n_43),
.Y(n_54)
);

OR2x2_ASAP7_75t_L g55 ( 
.A(n_24),
.B(n_42),
.Y(n_55)
);

BUFx12f_ASAP7_75t_L g56 ( 
.A(n_32),
.Y(n_56)
);

OAI22xp5_ASAP7_75t_SL g60 ( 
.A1(n_59),
.A2(n_48),
.B1(n_37),
.B2(n_54),
.Y(n_60)
);

AOI21xp5_ASAP7_75t_L g62 ( 
.A1(n_60),
.A2(n_61),
.B(n_58),
.Y(n_62)
);

OR2x2_ASAP7_75t_L g61 ( 
.A(n_58),
.B(n_54),
.Y(n_61)
);

BUFx24_ASAP7_75t_SL g64 ( 
.A(n_62),
.Y(n_64)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_61),
.Y(n_63)
);

XNOR2xp5_ASAP7_75t_L g65 ( 
.A(n_64),
.B(n_63),
.Y(n_65)
);

MAJIxp5_ASAP7_75t_L g68 ( 
.A(n_65),
.B(n_52),
.C(n_55),
.Y(n_68)
);

AOI21xp5_ASAP7_75t_L g66 ( 
.A1(n_64),
.A2(n_38),
.B(n_34),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_L g67 ( 
.A(n_66),
.B(n_31),
.Y(n_67)
);

AOI21xp5_ASAP7_75t_L g70 ( 
.A1(n_67),
.A2(n_68),
.B(n_52),
.Y(n_70)
);

AOI22xp5_ASAP7_75t_L g69 ( 
.A1(n_67),
.A2(n_23),
.B1(n_27),
.B2(n_43),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_SL g72 ( 
.A(n_69),
.B(n_70),
.Y(n_72)
);

XNOR2xp5_ASAP7_75t_SL g71 ( 
.A(n_69),
.B(n_33),
.Y(n_71)
);

A2O1A1Ixp33_ASAP7_75t_SL g74 ( 
.A1(n_71),
.A2(n_41),
.B(n_30),
.C(n_33),
.Y(n_74)
);

NOR3xp33_ASAP7_75t_L g73 ( 
.A(n_72),
.B(n_45),
.C(n_27),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_L g75 ( 
.A(n_73),
.B(n_23),
.Y(n_75)
);

AOI311xp33_ASAP7_75t_SL g76 ( 
.A1(n_74),
.A2(n_53),
.A3(n_46),
.B(n_47),
.C(n_57),
.Y(n_76)
);

OAI21xp5_ASAP7_75t_L g77 ( 
.A1(n_75),
.A2(n_76),
.B(n_57),
.Y(n_77)
);

OAI22xp5_ASAP7_75t_SL g78 ( 
.A1(n_77),
.A2(n_40),
.B1(n_56),
.B2(n_29),
.Y(n_78)
);

XOR2xp5_ASAP7_75t_L g79 ( 
.A(n_78),
.B(n_44),
.Y(n_79)
);


endmodule