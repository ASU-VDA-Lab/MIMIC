module real_jpeg_8354_n_16 (n_5, n_4, n_8, n_0, n_12, n_319, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_3, n_10, n_9, n_16);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_319;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_16;

wire n_37;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_300;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_199;
wire n_95;
wire n_238;
wire n_67;
wire n_235;
wire n_107;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_123;
wire n_50;
wire n_186;
wire n_137;
wire n_72;
wire n_171;
wire n_151;
wire n_272;
wire n_203;
wire n_198;
wire n_23;
wire n_71;
wire n_61;
wire n_99;
wire n_80;
wire n_30;
wire n_149;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_230;
wire n_128;
wire n_202;
wire n_216;
wire n_127;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_252;
wire n_310;
wire n_83;
wire n_78;
wire n_288;
wire n_221;
wire n_104;
wire n_153;
wire n_131;
wire n_87;
wire n_40;
wire n_98;
wire n_200;
wire n_214;
wire n_113;
wire n_251;
wire n_139;
wire n_33;
wire n_175;
wire n_156;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_77;
wire n_219;
wire n_122;
wire n_19;
wire n_262;
wire n_17;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_20;
wire n_278;
wire n_314;
wire n_103;
wire n_232;
wire n_212;
wire n_284;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_213;
wire n_25;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_49;
wire n_68;
wire n_146;
wire n_286;
wire n_166;
wire n_176;
wire n_215;
wire n_312;
wire n_316;
wire n_307;
wire n_161;
wire n_207;
wire n_237;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_140;
wire n_126;
wire n_120;
wire n_155;
wire n_93;
wire n_242;
wire n_142;
wire n_76;
wire n_79;
wire n_282;
wire n_147;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_18;
wire n_145;
wire n_266;
wire n_109;
wire n_148;
wire n_196;
wire n_298;
wire n_152;
wire n_270;
wire n_159;
wire n_183;
wire n_248;
wire n_192;
wire n_90;
wire n_258;
wire n_150;
wire n_41;
wire n_74;
wire n_204;
wire n_158;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_75;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_119;
wire n_283;
wire n_181;
wire n_256;
wire n_253;
wire n_273;
wire n_54;
wire n_168;
wire n_38;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_292;
wire n_64;
wire n_291;
wire n_236;
wire n_276;
wire n_287;
wire n_174;
wire n_255;
wire n_243;
wire n_299;
wire n_56;
wire n_293;
wire n_275;
wire n_227;
wire n_229;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_45;
wire n_268;
wire n_42;
wire n_313;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_143;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_303;
wire n_100;
wire n_51;
wire n_205;
wire n_261;
wire n_86;
wire n_70;
wire n_32;
wire n_228;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_169;
wire n_88;
wire n_167;
wire n_295;
wire n_133;
wire n_257;
wire n_210;
wire n_206;
wire n_85;
wire n_96;
wire n_308;

BUFx24_ASAP7_75t_L g28 ( 
.A(n_0),
.Y(n_28)
);

BUFx12_ASAP7_75t_L g25 ( 
.A(n_1),
.Y(n_25)
);

BUFx10_ASAP7_75t_L g91 ( 
.A(n_2),
.Y(n_91)
);

BUFx12f_ASAP7_75t_L g67 ( 
.A(n_3),
.Y(n_67)
);

BUFx10_ASAP7_75t_L g62 ( 
.A(n_4),
.Y(n_62)
);

BUFx6f_ASAP7_75t_SL g46 ( 
.A(n_5),
.Y(n_46)
);

BUFx12f_ASAP7_75t_L g50 ( 
.A(n_6),
.Y(n_50)
);

OAI22xp5_ASAP7_75t_SL g53 ( 
.A1(n_7),
.A2(n_26),
.B1(n_27),
.B2(n_54),
.Y(n_53)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_7),
.Y(n_54)
);

AOI22xp5_ASAP7_75t_SL g96 ( 
.A1(n_7),
.A2(n_49),
.B1(n_51),
.B2(n_54),
.Y(n_96)
);

AOI22xp33_ASAP7_75t_SL g110 ( 
.A1(n_7),
.A2(n_31),
.B1(n_32),
.B2(n_54),
.Y(n_110)
);

AOI22xp5_ASAP7_75t_L g247 ( 
.A1(n_7),
.A2(n_54),
.B1(n_65),
.B2(n_66),
.Y(n_247)
);

AOI22xp33_ASAP7_75t_SL g159 ( 
.A1(n_8),
.A2(n_65),
.B1(n_66),
.B2(n_160),
.Y(n_159)
);

CKINVDCx20_ASAP7_75t_R g160 ( 
.A(n_8),
.Y(n_160)
);

AOI22xp33_ASAP7_75t_SL g193 ( 
.A1(n_8),
.A2(n_49),
.B1(n_51),
.B2(n_160),
.Y(n_193)
);

AOI22xp33_ASAP7_75t_SL g221 ( 
.A1(n_8),
.A2(n_26),
.B1(n_27),
.B2(n_160),
.Y(n_221)
);

AOI22xp33_ASAP7_75t_SL g270 ( 
.A1(n_8),
.A2(n_31),
.B1(n_32),
.B2(n_160),
.Y(n_270)
);

AOI21xp5_ASAP7_75t_L g166 ( 
.A1(n_9),
.A2(n_51),
.B(n_167),
.Y(n_166)
);

NOR2xp33_ASAP7_75t_L g167 ( 
.A(n_9),
.B(n_51),
.Y(n_167)
);

CKINVDCx20_ASAP7_75t_R g178 ( 
.A(n_9),
.Y(n_178)
);

OAI22xp5_ASAP7_75t_L g182 ( 
.A1(n_9),
.A2(n_89),
.B1(n_92),
.B2(n_180),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_L g226 ( 
.A(n_9),
.B(n_104),
.Y(n_226)
);

AOI21xp33_ASAP7_75t_L g244 ( 
.A1(n_9),
.A2(n_25),
.B(n_27),
.Y(n_244)
);

OAI22xp33_ASAP7_75t_SL g259 ( 
.A1(n_9),
.A2(n_31),
.B1(n_32),
.B2(n_178),
.Y(n_259)
);

AOI22xp33_ASAP7_75t_SL g141 ( 
.A1(n_10),
.A2(n_31),
.B1(n_32),
.B2(n_142),
.Y(n_141)
);

CKINVDCx20_ASAP7_75t_R g142 ( 
.A(n_10),
.Y(n_142)
);

AOI22xp33_ASAP7_75t_SL g162 ( 
.A1(n_10),
.A2(n_65),
.B1(n_66),
.B2(n_142),
.Y(n_162)
);

AOI22xp33_ASAP7_75t_SL g201 ( 
.A1(n_10),
.A2(n_49),
.B1(n_51),
.B2(n_142),
.Y(n_201)
);

AOI22xp33_ASAP7_75t_SL g257 ( 
.A1(n_10),
.A2(n_26),
.B1(n_27),
.B2(n_142),
.Y(n_257)
);

BUFx10_ASAP7_75t_L g32 ( 
.A(n_11),
.Y(n_32)
);

OAI22xp5_ASAP7_75t_SL g70 ( 
.A1(n_12),
.A2(n_49),
.B1(n_51),
.B2(n_71),
.Y(n_70)
);

CKINVDCx20_ASAP7_75t_R g71 ( 
.A(n_12),
.Y(n_71)
);

OAI22xp33_ASAP7_75t_SL g94 ( 
.A1(n_12),
.A2(n_65),
.B1(n_66),
.B2(n_71),
.Y(n_94)
);

OAI22xp5_ASAP7_75t_SL g102 ( 
.A1(n_12),
.A2(n_31),
.B1(n_32),
.B2(n_71),
.Y(n_102)
);

OAI22xp5_ASAP7_75t_L g115 ( 
.A1(n_12),
.A2(n_26),
.B1(n_27),
.B2(n_71),
.Y(n_115)
);

AOI22xp5_ASAP7_75t_SL g168 ( 
.A1(n_13),
.A2(n_49),
.B1(n_51),
.B2(n_169),
.Y(n_168)
);

CKINVDCx20_ASAP7_75t_R g169 ( 
.A(n_13),
.Y(n_169)
);

AOI22xp33_ASAP7_75t_SL g180 ( 
.A1(n_13),
.A2(n_65),
.B1(n_66),
.B2(n_169),
.Y(n_180)
);

OAI22xp5_ASAP7_75t_SL g204 ( 
.A1(n_13),
.A2(n_26),
.B1(n_27),
.B2(n_169),
.Y(n_204)
);

AOI22xp33_ASAP7_75t_L g261 ( 
.A1(n_13),
.A2(n_31),
.B1(n_32),
.B2(n_169),
.Y(n_261)
);

AOI22xp33_ASAP7_75t_SL g30 ( 
.A1(n_14),
.A2(n_31),
.B1(n_32),
.B2(n_33),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_14),
.Y(n_33)
);

AOI22xp33_ASAP7_75t_SL g77 ( 
.A1(n_14),
.A2(n_26),
.B1(n_27),
.B2(n_33),
.Y(n_77)
);

AOI22xp5_ASAP7_75t_L g138 ( 
.A1(n_14),
.A2(n_33),
.B1(n_49),
.B2(n_51),
.Y(n_138)
);

AOI22xp33_ASAP7_75t_SL g225 ( 
.A1(n_14),
.A2(n_33),
.B1(n_65),
.B2(n_66),
.Y(n_225)
);

OAI22xp33_ASAP7_75t_SL g35 ( 
.A1(n_15),
.A2(n_31),
.B1(n_32),
.B2(n_36),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_15),
.Y(n_36)
);

AOI22xp33_ASAP7_75t_L g57 ( 
.A1(n_15),
.A2(n_26),
.B1(n_27),
.B2(n_36),
.Y(n_57)
);

AOI22xp33_ASAP7_75t_L g83 ( 
.A1(n_15),
.A2(n_36),
.B1(n_49),
.B2(n_51),
.Y(n_83)
);

OAI22xp33_ASAP7_75t_SL g135 ( 
.A1(n_15),
.A2(n_36),
.B1(n_65),
.B2(n_66),
.Y(n_135)
);

XOR2xp5_ASAP7_75t_L g16 ( 
.A(n_17),
.B(n_122),
.Y(n_16)
);

NAND2xp5_ASAP7_75t_SL g17 ( 
.A(n_18),
.B(n_121),
.Y(n_17)
);

INVxp67_ASAP7_75t_L g18 ( 
.A(n_19),
.Y(n_18)
);

NOR2xp33_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_105),
.Y(n_19)
);

NAND2xp5_ASAP7_75t_L g121 ( 
.A(n_20),
.B(n_105),
.Y(n_121)
);

MAJIxp5_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_73),
.C(n_85),
.Y(n_20)
);

OAI22xp5_ASAP7_75t_SL g147 ( 
.A1(n_21),
.A2(n_73),
.B1(n_74),
.B2(n_148),
.Y(n_147)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_21),
.Y(n_148)
);

AOI22xp5_ASAP7_75t_L g21 ( 
.A1(n_22),
.A2(n_23),
.B1(n_40),
.B2(n_41),
.Y(n_21)
);

OAI22xp5_ASAP7_75t_SL g106 ( 
.A1(n_22),
.A2(n_23),
.B1(n_107),
.B2(n_108),
.Y(n_106)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_23),
.Y(n_22)
);

MAJIxp5_ASAP7_75t_L g120 ( 
.A(n_23),
.B(n_59),
.C(n_72),
.Y(n_120)
);

OAI21xp5_ASAP7_75t_L g23 ( 
.A1(n_24),
.A2(n_30),
.B(n_34),
.Y(n_23)
);

A2O1A1Ixp33_ASAP7_75t_L g38 ( 
.A1(n_24),
.A2(n_29),
.B(n_32),
.C(n_39),
.Y(n_38)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_24),
.Y(n_104)
);

OAI22xp5_ASAP7_75t_SL g109 ( 
.A1(n_24),
.A2(n_30),
.B1(n_38),
.B2(n_110),
.Y(n_109)
);

OAI22xp5_ASAP7_75t_SL g269 ( 
.A1(n_24),
.A2(n_38),
.B1(n_261),
.B2(n_270),
.Y(n_269)
);

OAI22xp5_ASAP7_75t_SL g285 ( 
.A1(n_24),
.A2(n_38),
.B1(n_141),
.B2(n_270),
.Y(n_285)
);

AOI22xp5_ASAP7_75t_L g24 ( 
.A1(n_25),
.A2(n_26),
.B1(n_27),
.B2(n_29),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_25),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_27),
.Y(n_26)
);

O2A1O1Ixp33_ASAP7_75t_L g44 ( 
.A1(n_27),
.A2(n_45),
.B(n_47),
.C(n_48),
.Y(n_44)
);

NAND2xp5_ASAP7_75t_L g47 ( 
.A(n_27),
.B(n_45),
.Y(n_47)
);

HAxp5_ASAP7_75t_SL g203 ( 
.A(n_27),
.B(n_178),
.CON(n_203),
.SN(n_203)
);

BUFx10_ASAP7_75t_L g27 ( 
.A(n_28),
.Y(n_27)
);

NOR2xp33_ASAP7_75t_L g39 ( 
.A(n_29),
.B(n_32),
.Y(n_39)
);

A2O1A1Ixp33_ASAP7_75t_L g243 ( 
.A1(n_29),
.A2(n_32),
.B(n_178),
.C(n_244),
.Y(n_243)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_32),
.Y(n_31)
);

NAND2xp5_ASAP7_75t_L g34 ( 
.A(n_35),
.B(n_37),
.Y(n_34)
);

NAND2xp5_ASAP7_75t_L g103 ( 
.A(n_35),
.B(n_104),
.Y(n_103)
);

AOI22xp5_ASAP7_75t_SL g258 ( 
.A1(n_37),
.A2(n_104),
.B1(n_259),
.B2(n_260),
.Y(n_258)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_38),
.Y(n_37)
);

OAI21xp5_ASAP7_75t_SL g100 ( 
.A1(n_38),
.A2(n_101),
.B(n_103),
.Y(n_100)
);

OAI21xp5_ASAP7_75t_SL g140 ( 
.A1(n_38),
.A2(n_141),
.B(n_143),
.Y(n_140)
);

CKINVDCx14_ASAP7_75t_R g40 ( 
.A(n_41),
.Y(n_40)
);

OAI22xp5_ASAP7_75t_L g41 ( 
.A1(n_42),
.A2(n_59),
.B1(n_60),
.B2(n_72),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g72 ( 
.A(n_42),
.Y(n_72)
);

OAI21xp5_ASAP7_75t_SL g42 ( 
.A1(n_43),
.A2(n_52),
.B(n_55),
.Y(n_42)
);

OAI22xp5_ASAP7_75t_SL g219 ( 
.A1(n_43),
.A2(n_58),
.B1(n_220),
.B2(n_221),
.Y(n_219)
);

OAI22xp5_ASAP7_75t_L g256 ( 
.A1(n_43),
.A2(n_58),
.B1(n_221),
.B2(n_257),
.Y(n_256)
);

OAI21xp5_ASAP7_75t_SL g271 ( 
.A1(n_43),
.A2(n_114),
.B(n_257),
.Y(n_271)
);

CKINVDCx16_ASAP7_75t_R g43 ( 
.A(n_44),
.Y(n_43)
);

AOI22xp5_ASAP7_75t_L g75 ( 
.A1(n_44),
.A2(n_48),
.B1(n_53),
.B2(n_76),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_SL g116 ( 
.A(n_44),
.B(n_117),
.Y(n_116)
);

AOI22xp5_ASAP7_75t_L g202 ( 
.A1(n_44),
.A2(n_48),
.B1(n_203),
.B2(n_204),
.Y(n_202)
);

AOI21xp5_ASAP7_75t_L g287 ( 
.A1(n_44),
.A2(n_56),
.B(n_115),
.Y(n_287)
);

OAI22xp5_ASAP7_75t_SL g48 ( 
.A1(n_45),
.A2(n_46),
.B1(n_49),
.B2(n_51),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_SL g209 ( 
.A(n_45),
.B(n_51),
.Y(n_209)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_46),
.Y(n_45)
);

OAI22xp5_ASAP7_75t_L g208 ( 
.A1(n_47),
.A2(n_49),
.B1(n_203),
.B2(n_209),
.Y(n_208)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_48),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_L g114 ( 
.A(n_48),
.B(n_115),
.Y(n_114)
);

INVx8_ASAP7_75t_L g51 ( 
.A(n_49),
.Y(n_51)
);

BUFx3_ASAP7_75t_L g49 ( 
.A(n_50),
.Y(n_49)
);

A2O1A1Ixp33_ASAP7_75t_SL g61 ( 
.A1(n_51),
.A2(n_62),
.B(n_63),
.C(n_64),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_51),
.B(n_62),
.Y(n_63)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_53),
.Y(n_52)
);

CKINVDCx20_ASAP7_75t_R g55 ( 
.A(n_56),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_57),
.B(n_58),
.Y(n_56)
);

INVxp67_ASAP7_75t_L g117 ( 
.A(n_57),
.Y(n_117)
);

OAI21xp5_ASAP7_75t_L g145 ( 
.A1(n_58),
.A2(n_77),
.B(n_116),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_L g191 ( 
.A(n_58),
.B(n_178),
.Y(n_191)
);

OAI22xp5_ASAP7_75t_SL g112 ( 
.A1(n_59),
.A2(n_60),
.B1(n_113),
.B2(n_118),
.Y(n_112)
);

CKINVDCx20_ASAP7_75t_R g59 ( 
.A(n_60),
.Y(n_59)
);

AOI21xp5_ASAP7_75t_SL g60 ( 
.A1(n_61),
.A2(n_64),
.B(n_69),
.Y(n_60)
);

CKINVDCx16_ASAP7_75t_R g84 ( 
.A(n_61),
.Y(n_84)
);

OAI21xp5_ASAP7_75t_SL g95 ( 
.A1(n_61),
.A2(n_96),
.B(n_97),
.Y(n_95)
);

OAI22xp5_ASAP7_75t_L g137 ( 
.A1(n_61),
.A2(n_64),
.B1(n_96),
.B2(n_138),
.Y(n_137)
);

OAI22xp5_ASAP7_75t_L g165 ( 
.A1(n_61),
.A2(n_64),
.B1(n_166),
.B2(n_168),
.Y(n_165)
);

OAI22xp5_ASAP7_75t_SL g192 ( 
.A1(n_61),
.A2(n_64),
.B1(n_168),
.B2(n_193),
.Y(n_192)
);

OAI22xp5_ASAP7_75t_L g200 ( 
.A1(n_61),
.A2(n_64),
.B1(n_193),
.B2(n_201),
.Y(n_200)
);

OAI21xp5_ASAP7_75t_SL g233 ( 
.A1(n_61),
.A2(n_79),
.B(n_201),
.Y(n_233)
);

AOI22xp5_ASAP7_75t_SL g64 ( 
.A1(n_62),
.A2(n_65),
.B1(n_66),
.B2(n_68),
.Y(n_64)
);

CKINVDCx16_ASAP7_75t_R g68 ( 
.A(n_62),
.Y(n_68)
);

INVxp67_ASAP7_75t_L g173 ( 
.A(n_63),
.Y(n_173)
);

INVxp67_ASAP7_75t_L g80 ( 
.A(n_64),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_64),
.B(n_83),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_SL g177 ( 
.A(n_64),
.B(n_178),
.Y(n_177)
);

OAI21xp5_ASAP7_75t_L g275 ( 
.A1(n_64),
.A2(n_81),
.B(n_138),
.Y(n_275)
);

NOR2xp33_ASAP7_75t_SL g90 ( 
.A(n_65),
.B(n_91),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_SL g171 ( 
.A(n_65),
.B(n_68),
.Y(n_171)
);

NOR2xp33_ASAP7_75t_SL g183 ( 
.A(n_65),
.B(n_184),
.Y(n_183)
);

CKINVDCx20_ASAP7_75t_R g65 ( 
.A(n_66),
.Y(n_65)
);

OAI22xp5_ASAP7_75t_L g170 ( 
.A1(n_66),
.A2(n_171),
.B1(n_172),
.B2(n_173),
.Y(n_170)
);

BUFx24_ASAP7_75t_L g66 ( 
.A(n_67),
.Y(n_66)
);

INVxp67_ASAP7_75t_L g69 ( 
.A(n_70),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_L g79 ( 
.A(n_70),
.B(n_80),
.Y(n_79)
);

AOI21xp5_ASAP7_75t_L g254 ( 
.A1(n_70),
.A2(n_84),
.B(n_98),
.Y(n_254)
);

CKINVDCx20_ASAP7_75t_R g73 ( 
.A(n_74),
.Y(n_73)
);

OAI21xp5_ASAP7_75t_L g130 ( 
.A1(n_74),
.A2(n_75),
.B(n_78),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_L g74 ( 
.A(n_75),
.B(n_78),
.Y(n_74)
);

CKINVDCx20_ASAP7_75t_R g76 ( 
.A(n_77),
.Y(n_76)
);

AND2x2_ASAP7_75t_L g78 ( 
.A(n_79),
.B(n_81),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_L g81 ( 
.A(n_82),
.B(n_84),
.Y(n_81)
);

INVxp67_ASAP7_75t_L g82 ( 
.A(n_83),
.Y(n_82)
);

XNOR2xp5_ASAP7_75t_L g146 ( 
.A(n_85),
.B(n_147),
.Y(n_146)
);

OAI21xp5_ASAP7_75t_L g85 ( 
.A1(n_86),
.A2(n_99),
.B(n_100),
.Y(n_85)
);

OAI22xp5_ASAP7_75t_L g126 ( 
.A1(n_86),
.A2(n_87),
.B1(n_127),
.B2(n_128),
.Y(n_126)
);

CKINVDCx20_ASAP7_75t_R g86 ( 
.A(n_87),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_L g87 ( 
.A(n_88),
.B(n_95),
.Y(n_87)
);

CKINVDCx20_ASAP7_75t_R g99 ( 
.A(n_88),
.Y(n_99)
);

AOI22xp5_ASAP7_75t_L g128 ( 
.A1(n_88),
.A2(n_99),
.B1(n_100),
.B2(n_129),
.Y(n_128)
);

OAI22xp5_ASAP7_75t_L g305 ( 
.A1(n_88),
.A2(n_95),
.B1(n_99),
.B2(n_306),
.Y(n_305)
);

AOI21xp5_ASAP7_75t_L g88 ( 
.A1(n_89),
.A2(n_92),
.B(n_93),
.Y(n_88)
);

OAI22xp5_ASAP7_75t_SL g179 ( 
.A1(n_89),
.A2(n_92),
.B1(n_159),
.B2(n_180),
.Y(n_179)
);

OAI21xp5_ASAP7_75t_L g194 ( 
.A1(n_89),
.A2(n_136),
.B(n_162),
.Y(n_194)
);

OAI21xp5_ASAP7_75t_SL g210 ( 
.A1(n_89),
.A2(n_93),
.B(n_211),
.Y(n_210)
);

OAI22xp5_ASAP7_75t_SL g246 ( 
.A1(n_89),
.A2(n_92),
.B1(n_225),
.B2(n_247),
.Y(n_246)
);

OAI21xp5_ASAP7_75t_SL g276 ( 
.A1(n_89),
.A2(n_211),
.B(n_247),
.Y(n_276)
);

CKINVDCx20_ASAP7_75t_R g89 ( 
.A(n_90),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_SL g134 ( 
.A(n_90),
.B(n_135),
.Y(n_134)
);

AOI22xp5_ASAP7_75t_SL g157 ( 
.A1(n_90),
.A2(n_91),
.B1(n_158),
.B2(n_161),
.Y(n_157)
);

CKINVDCx16_ASAP7_75t_R g92 ( 
.A(n_91),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_L g136 ( 
.A(n_91),
.B(n_94),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_L g211 ( 
.A(n_91),
.B(n_135),
.Y(n_211)
);

NOR2xp33_ASAP7_75t_L g184 ( 
.A(n_92),
.B(n_178),
.Y(n_184)
);

OAI21xp5_ASAP7_75t_L g224 ( 
.A1(n_92),
.A2(n_134),
.B(n_225),
.Y(n_224)
);

CKINVDCx20_ASAP7_75t_R g93 ( 
.A(n_94),
.Y(n_93)
);

CKINVDCx14_ASAP7_75t_R g306 ( 
.A(n_95),
.Y(n_306)
);

CKINVDCx20_ASAP7_75t_R g97 ( 
.A(n_98),
.Y(n_97)
);

CKINVDCx20_ASAP7_75t_R g129 ( 
.A(n_100),
.Y(n_129)
);

CKINVDCx20_ASAP7_75t_R g101 ( 
.A(n_102),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_SL g143 ( 
.A(n_102),
.B(n_104),
.Y(n_143)
);

XOR2xp5_ASAP7_75t_L g105 ( 
.A(n_106),
.B(n_120),
.Y(n_105)
);

CKINVDCx14_ASAP7_75t_R g107 ( 
.A(n_108),
.Y(n_107)
);

AOI22xp5_ASAP7_75t_L g108 ( 
.A1(n_109),
.A2(n_111),
.B1(n_112),
.B2(n_119),
.Y(n_108)
);

CKINVDCx20_ASAP7_75t_R g119 ( 
.A(n_109),
.Y(n_119)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_112),
.Y(n_111)
);

CKINVDCx20_ASAP7_75t_R g118 ( 
.A(n_113),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_L g113 ( 
.A(n_114),
.B(n_116),
.Y(n_113)
);

OAI21xp5_ASAP7_75t_L g122 ( 
.A1(n_123),
.A2(n_149),
.B(n_317),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_L g123 ( 
.A(n_124),
.B(n_146),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_SL g317 ( 
.A(n_124),
.B(n_146),
.Y(n_317)
);

CKINVDCx5p33_ASAP7_75t_R g124 ( 
.A(n_125),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_L g308 ( 
.A(n_125),
.B(n_309),
.Y(n_308)
);

NOR2xp33_ASAP7_75t_SL g316 ( 
.A(n_125),
.B(n_309),
.Y(n_316)
);

FAx1_ASAP7_75t_SL g125 ( 
.A(n_126),
.B(n_130),
.CI(n_131),
.CON(n_125),
.SN(n_125)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_128),
.Y(n_127)
);

MAJIxp5_ASAP7_75t_L g131 ( 
.A(n_132),
.B(n_139),
.C(n_144),
.Y(n_131)
);

XOR2xp5_ASAP7_75t_L g302 ( 
.A(n_132),
.B(n_303),
.Y(n_302)
);

NAND2xp5_ASAP7_75t_L g132 ( 
.A(n_133),
.B(n_137),
.Y(n_132)
);

XNOR2xp5_ASAP7_75t_L g288 ( 
.A(n_133),
.B(n_137),
.Y(n_288)
);

NAND2xp5_ASAP7_75t_L g133 ( 
.A(n_134),
.B(n_136),
.Y(n_133)
);

OAI22xp5_ASAP7_75t_L g303 ( 
.A1(n_139),
.A2(n_140),
.B1(n_144),
.B2(n_145),
.Y(n_303)
);

CKINVDCx20_ASAP7_75t_R g139 ( 
.A(n_140),
.Y(n_139)
);

CKINVDCx20_ASAP7_75t_R g144 ( 
.A(n_145),
.Y(n_144)
);

AOI321xp33_ASAP7_75t_L g149 ( 
.A1(n_150),
.A2(n_296),
.A3(n_308),
.B1(n_310),
.B2(n_316),
.C(n_319),
.Y(n_149)
);

NOR3xp33_ASAP7_75t_L g150 ( 
.A(n_151),
.B(n_263),
.C(n_292),
.Y(n_150)
);

AOI21xp5_ASAP7_75t_L g151 ( 
.A1(n_152),
.A2(n_237),
.B(n_262),
.Y(n_151)
);

OAI21xp5_ASAP7_75t_SL g152 ( 
.A1(n_153),
.A2(n_214),
.B(n_236),
.Y(n_152)
);

AOI21xp5_ASAP7_75t_L g153 ( 
.A1(n_154),
.A2(n_196),
.B(n_213),
.Y(n_153)
);

OAI21xp5_ASAP7_75t_SL g154 ( 
.A1(n_155),
.A2(n_187),
.B(n_195),
.Y(n_154)
);

AOI21xp5_ASAP7_75t_L g155 ( 
.A1(n_156),
.A2(n_175),
.B(n_186),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_L g156 ( 
.A(n_157),
.B(n_163),
.Y(n_156)
);

NOR2xp33_ASAP7_75t_SL g186 ( 
.A(n_157),
.B(n_163),
.Y(n_186)
);

CKINVDCx20_ASAP7_75t_R g158 ( 
.A(n_159),
.Y(n_158)
);

CKINVDCx20_ASAP7_75t_R g161 ( 
.A(n_162),
.Y(n_161)
);

AOI22xp5_ASAP7_75t_SL g163 ( 
.A1(n_164),
.A2(n_165),
.B1(n_170),
.B2(n_174),
.Y(n_163)
);

NOR2xp33_ASAP7_75t_SL g188 ( 
.A(n_164),
.B(n_174),
.Y(n_188)
);

CKINVDCx20_ASAP7_75t_R g164 ( 
.A(n_165),
.Y(n_164)
);

CKINVDCx20_ASAP7_75t_R g172 ( 
.A(n_167),
.Y(n_172)
);

CKINVDCx20_ASAP7_75t_R g174 ( 
.A(n_170),
.Y(n_174)
);

OAI21xp5_ASAP7_75t_SL g175 ( 
.A1(n_176),
.A2(n_181),
.B(n_185),
.Y(n_175)
);

NOR2xp33_ASAP7_75t_L g176 ( 
.A(n_177),
.B(n_179),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_SL g185 ( 
.A(n_177),
.B(n_179),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_SL g181 ( 
.A(n_182),
.B(n_183),
.Y(n_181)
);

NOR2xp33_ASAP7_75t_L g187 ( 
.A(n_188),
.B(n_189),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_SL g195 ( 
.A(n_188),
.B(n_189),
.Y(n_195)
);

CKINVDCx5p33_ASAP7_75t_R g189 ( 
.A(n_190),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_L g196 ( 
.A(n_190),
.B(n_197),
.Y(n_196)
);

NOR2xp33_ASAP7_75t_SL g213 ( 
.A(n_190),
.B(n_197),
.Y(n_213)
);

FAx1_ASAP7_75t_SL g190 ( 
.A(n_191),
.B(n_192),
.CI(n_194),
.CON(n_190),
.SN(n_190)
);

AOI22xp33_ASAP7_75t_SL g197 ( 
.A1(n_198),
.A2(n_199),
.B1(n_207),
.B2(n_212),
.Y(n_197)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_199),
.Y(n_198)
);

OAI22xp5_ASAP7_75t_L g199 ( 
.A1(n_200),
.A2(n_202),
.B1(n_205),
.B2(n_206),
.Y(n_199)
);

CKINVDCx20_ASAP7_75t_R g206 ( 
.A(n_200),
.Y(n_206)
);

CKINVDCx20_ASAP7_75t_R g205 ( 
.A(n_202),
.Y(n_205)
);

MAJIxp5_ASAP7_75t_L g215 ( 
.A(n_202),
.B(n_206),
.C(n_212),
.Y(n_215)
);

CKINVDCx20_ASAP7_75t_R g220 ( 
.A(n_204),
.Y(n_220)
);

CKINVDCx20_ASAP7_75t_R g212 ( 
.A(n_207),
.Y(n_212)
);

XOR2xp5_ASAP7_75t_L g207 ( 
.A(n_208),
.B(n_210),
.Y(n_207)
);

NAND2xp5_ASAP7_75t_L g232 ( 
.A(n_208),
.B(n_210),
.Y(n_232)
);

NOR2xp33_ASAP7_75t_L g214 ( 
.A(n_215),
.B(n_216),
.Y(n_214)
);

NAND2xp5_ASAP7_75t_SL g236 ( 
.A(n_215),
.B(n_216),
.Y(n_236)
);

OAI22xp5_ASAP7_75t_SL g216 ( 
.A1(n_217),
.A2(n_218),
.B1(n_230),
.B2(n_231),
.Y(n_216)
);

MAJIxp5_ASAP7_75t_L g238 ( 
.A(n_217),
.B(n_233),
.C(n_234),
.Y(n_238)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_218),
.Y(n_217)
);

AOI22xp5_ASAP7_75t_L g218 ( 
.A1(n_219),
.A2(n_222),
.B1(n_223),
.B2(n_229),
.Y(n_218)
);

CKINVDCx20_ASAP7_75t_R g229 ( 
.A(n_219),
.Y(n_229)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_223),
.Y(n_222)
);

OAI22xp5_ASAP7_75t_SL g223 ( 
.A1(n_224),
.A2(n_226),
.B1(n_227),
.B2(n_228),
.Y(n_223)
);

CKINVDCx20_ASAP7_75t_R g227 ( 
.A(n_224),
.Y(n_227)
);

CKINVDCx20_ASAP7_75t_R g228 ( 
.A(n_226),
.Y(n_228)
);

MAJIxp5_ASAP7_75t_L g248 ( 
.A(n_226),
.B(n_227),
.C(n_229),
.Y(n_248)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_231),
.Y(n_230)
);

OAI22xp5_ASAP7_75t_SL g231 ( 
.A1(n_232),
.A2(n_233),
.B1(n_234),
.B2(n_235),
.Y(n_231)
);

CKINVDCx20_ASAP7_75t_R g234 ( 
.A(n_232),
.Y(n_234)
);

CKINVDCx20_ASAP7_75t_R g235 ( 
.A(n_233),
.Y(n_235)
);

NAND2xp5_ASAP7_75t_L g237 ( 
.A(n_238),
.B(n_239),
.Y(n_237)
);

NOR2xp33_ASAP7_75t_SL g262 ( 
.A(n_238),
.B(n_239),
.Y(n_262)
);

XOR2xp5_ASAP7_75t_L g239 ( 
.A(n_240),
.B(n_251),
.Y(n_239)
);

OAI22xp5_ASAP7_75t_L g240 ( 
.A1(n_241),
.A2(n_248),
.B1(n_249),
.B2(n_250),
.Y(n_240)
);

CKINVDCx16_ASAP7_75t_R g249 ( 
.A(n_241),
.Y(n_249)
);

MAJIxp5_ASAP7_75t_L g293 ( 
.A(n_241),
.B(n_250),
.C(n_251),
.Y(n_293)
);

AOI22xp5_ASAP7_75t_L g241 ( 
.A1(n_242),
.A2(n_243),
.B1(n_245),
.B2(n_246),
.Y(n_241)
);

NAND2xp5_ASAP7_75t_L g266 ( 
.A(n_242),
.B(n_246),
.Y(n_266)
);

CKINVDCx20_ASAP7_75t_R g242 ( 
.A(n_243),
.Y(n_242)
);

CKINVDCx20_ASAP7_75t_R g245 ( 
.A(n_246),
.Y(n_245)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_248),
.Y(n_250)
);

XOR2xp5_ASAP7_75t_L g251 ( 
.A(n_252),
.B(n_258),
.Y(n_251)
);

OAI22xp5_ASAP7_75t_L g252 ( 
.A1(n_253),
.A2(n_254),
.B1(n_255),
.B2(n_256),
.Y(n_252)
);

CKINVDCx20_ASAP7_75t_R g253 ( 
.A(n_254),
.Y(n_253)
);

MAJIxp5_ASAP7_75t_L g278 ( 
.A(n_254),
.B(n_255),
.C(n_258),
.Y(n_278)
);

CKINVDCx20_ASAP7_75t_R g255 ( 
.A(n_256),
.Y(n_255)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_261),
.Y(n_260)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_263),
.Y(n_312)
);

NOR2xp33_ASAP7_75t_L g263 ( 
.A(n_264),
.B(n_279),
.Y(n_263)
);

AND2x2_ASAP7_75t_L g314 ( 
.A(n_264),
.B(n_279),
.Y(n_314)
);

MAJIxp5_ASAP7_75t_L g264 ( 
.A(n_265),
.B(n_273),
.C(n_277),
.Y(n_264)
);

XOR2xp5_ASAP7_75t_L g294 ( 
.A(n_265),
.B(n_295),
.Y(n_294)
);

XOR2xp5_ASAP7_75t_L g265 ( 
.A(n_266),
.B(n_267),
.Y(n_265)
);

MAJIxp5_ASAP7_75t_L g290 ( 
.A(n_266),
.B(n_268),
.C(n_272),
.Y(n_290)
);

OAI22xp5_ASAP7_75t_L g267 ( 
.A1(n_268),
.A2(n_269),
.B1(n_271),
.B2(n_272),
.Y(n_267)
);

CKINVDCx20_ASAP7_75t_R g268 ( 
.A(n_269),
.Y(n_268)
);

CKINVDCx20_ASAP7_75t_R g272 ( 
.A(n_271),
.Y(n_272)
);

AOI22xp5_ASAP7_75t_L g295 ( 
.A1(n_273),
.A2(n_274),
.B1(n_277),
.B2(n_278),
.Y(n_295)
);

CKINVDCx20_ASAP7_75t_R g273 ( 
.A(n_274),
.Y(n_273)
);

XOR2xp5_ASAP7_75t_L g274 ( 
.A(n_275),
.B(n_276),
.Y(n_274)
);

NAND2xp5_ASAP7_75t_L g282 ( 
.A(n_275),
.B(n_276),
.Y(n_282)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_278),
.Y(n_277)
);

OAI22xp5_ASAP7_75t_SL g279 ( 
.A1(n_280),
.A2(n_289),
.B1(n_290),
.B2(n_291),
.Y(n_279)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_280),
.Y(n_291)
);

XOR2xp5_ASAP7_75t_L g280 ( 
.A(n_281),
.B(n_288),
.Y(n_280)
);

MAJIxp5_ASAP7_75t_L g298 ( 
.A(n_281),
.B(n_288),
.C(n_289),
.Y(n_298)
);

XOR2xp5_ASAP7_75t_L g281 ( 
.A(n_282),
.B(n_283),
.Y(n_281)
);

MAJIxp5_ASAP7_75t_L g307 ( 
.A(n_282),
.B(n_284),
.C(n_287),
.Y(n_307)
);

OAI22xp5_ASAP7_75t_L g283 ( 
.A1(n_284),
.A2(n_285),
.B1(n_286),
.B2(n_287),
.Y(n_283)
);

CKINVDCx20_ASAP7_75t_R g284 ( 
.A(n_285),
.Y(n_284)
);

CKINVDCx14_ASAP7_75t_R g286 ( 
.A(n_287),
.Y(n_286)
);

CKINVDCx14_ASAP7_75t_R g289 ( 
.A(n_290),
.Y(n_289)
);

NOR2xp33_ASAP7_75t_L g292 ( 
.A(n_293),
.B(n_294),
.Y(n_292)
);

AND2x2_ASAP7_75t_L g313 ( 
.A(n_293),
.B(n_294),
.Y(n_313)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_297),
.Y(n_296)
);

OAI21xp5_ASAP7_75t_SL g310 ( 
.A1(n_297),
.A2(n_311),
.B(n_315),
.Y(n_310)
);

NOR2xp33_ASAP7_75t_L g297 ( 
.A(n_298),
.B(n_299),
.Y(n_297)
);

NAND2xp5_ASAP7_75t_SL g315 ( 
.A(n_298),
.B(n_299),
.Y(n_315)
);

XOR2xp5_ASAP7_75t_L g299 ( 
.A(n_300),
.B(n_307),
.Y(n_299)
);

OAI22xp5_ASAP7_75t_SL g300 ( 
.A1(n_301),
.A2(n_302),
.B1(n_304),
.B2(n_305),
.Y(n_300)
);

MAJIxp5_ASAP7_75t_L g309 ( 
.A(n_301),
.B(n_305),
.C(n_307),
.Y(n_309)
);

CKINVDCx14_ASAP7_75t_R g301 ( 
.A(n_302),
.Y(n_301)
);

CKINVDCx16_ASAP7_75t_R g304 ( 
.A(n_305),
.Y(n_304)
);

AOI21xp5_ASAP7_75t_L g311 ( 
.A1(n_312),
.A2(n_313),
.B(n_314),
.Y(n_311)
);


endmodule