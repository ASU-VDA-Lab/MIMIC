module real_jpeg_12587_n_6 (n_5, n_4, n_0, n_1, n_2, n_3, n_6);

input n_5;
input n_4;
input n_0;
input n_1;
input n_2;
input n_3;

output n_6;

wire n_17;
wire n_8;
wire n_43;
wire n_37;
wire n_21;
wire n_35;
wire n_33;
wire n_50;
wire n_38;
wire n_29;
wire n_49;
wire n_10;
wire n_31;
wire n_9;
wire n_52;
wire n_12;
wire n_24;
wire n_34;
wire n_28;
wire n_44;
wire n_46;
wire n_23;
wire n_11;
wire n_14;
wire n_47;
wire n_51;
wire n_45;
wire n_25;
wire n_42;
wire n_7;
wire n_22;
wire n_18;
wire n_53;
wire n_39;
wire n_36;
wire n_40;
wire n_41;
wire n_27;
wire n_26;
wire n_20;
wire n_19;
wire n_48;
wire n_32;
wire n_30;
wire n_16;
wire n_15;
wire n_13;

OAI221xp5_ASAP7_75t_SL g7 ( 
.A1(n_0),
.A2(n_8),
.B1(n_20),
.B2(n_31),
.C(n_35),
.Y(n_7)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_0),
.Y(n_17)
);

NOR2xp33_ASAP7_75t_L g18 ( 
.A(n_0),
.B(n_19),
.Y(n_18)
);

NAND2xp5_ASAP7_75t_SL g45 ( 
.A(n_0),
.B(n_1),
.Y(n_45)
);

AND2x2_ASAP7_75t_SL g13 ( 
.A(n_1),
.B(n_14),
.Y(n_13)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_1),
.Y(n_27)
);

NAND2xp5_ASAP7_75t_L g41 ( 
.A(n_1),
.B(n_28),
.Y(n_41)
);

NAND2xp5_ASAP7_75t_L g47 ( 
.A(n_1),
.B(n_9),
.Y(n_47)
);

NAND2xp5_ASAP7_75t_SL g53 ( 
.A(n_1),
.B(n_39),
.Y(n_53)
);

OR2x2_ASAP7_75t_SL g10 ( 
.A(n_2),
.B(n_11),
.Y(n_10)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_2),
.Y(n_30)
);

AND2x2_ASAP7_75t_L g44 ( 
.A(n_2),
.B(n_11),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g16 ( 
.A(n_3),
.B(n_17),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_3),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g11 ( 
.A(n_4),
.Y(n_11)
);

AO21x1_ASAP7_75t_SL g14 ( 
.A1(n_5),
.A2(n_15),
.B(n_18),
.Y(n_14)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_5),
.Y(n_24)
);

AOI22xp5_ASAP7_75t_SL g32 ( 
.A1(n_5),
.A2(n_24),
.B1(n_33),
.B2(n_34),
.Y(n_32)
);

NOR3xp33_ASAP7_75t_L g6 ( 
.A(n_7),
.B(n_46),
.C(n_50),
.Y(n_6)
);

NAND2xp5_ASAP7_75t_L g8 ( 
.A(n_9),
.B(n_12),
.Y(n_8)
);

CKINVDCx20_ASAP7_75t_R g9 ( 
.A(n_10),
.Y(n_9)
);

OR2x2_ASAP7_75t_SL g29 ( 
.A(n_11),
.B(n_30),
.Y(n_29)
);

AND2x2_ASAP7_75t_SL g39 ( 
.A(n_11),
.B(n_30),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g12 ( 
.A(n_13),
.Y(n_12)
);

OAI22xp5_ASAP7_75t_L g46 ( 
.A1(n_13),
.A2(n_47),
.B1(n_48),
.B2(n_49),
.Y(n_46)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_14),
.Y(n_48)
);

INVx1_ASAP7_75t_L g15 ( 
.A(n_16),
.Y(n_15)
);

OR2x2_ASAP7_75t_L g34 ( 
.A(n_16),
.B(n_18),
.Y(n_34)
);

NAND2xp5_ASAP7_75t_L g25 ( 
.A(n_17),
.B(n_19),
.Y(n_25)
);

NOR2xp33_ASAP7_75t_L g26 ( 
.A(n_17),
.B(n_19),
.Y(n_26)
);

NAND2xp5_ASAP7_75t_SL g20 ( 
.A(n_21),
.B(n_28),
.Y(n_20)
);

INVx1_ASAP7_75t_SL g21 ( 
.A(n_22),
.Y(n_21)
);

NOR2xp33_ASAP7_75t_L g40 ( 
.A(n_22),
.B(n_41),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_SL g22 ( 
.A(n_23),
.B(n_27),
.Y(n_22)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_23),
.Y(n_36)
);

AOI21xp5_ASAP7_75t_SL g23 ( 
.A1(n_24),
.A2(n_25),
.B(n_26),
.Y(n_23)
);

NAND2xp5_ASAP7_75t_L g38 ( 
.A(n_27),
.B(n_39),
.Y(n_38)
);

NAND2xp5_ASAP7_75t_SL g49 ( 
.A(n_27),
.B(n_44),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_29),
.Y(n_28)
);

NAND2xp5_ASAP7_75t_L g51 ( 
.A(n_31),
.B(n_52),
.Y(n_51)
);

INVx1_ASAP7_75t_SL g31 ( 
.A(n_32),
.Y(n_31)
);

INVx1_ASAP7_75t_SL g33 ( 
.A(n_34),
.Y(n_33)
);

AOI211xp5_ASAP7_75t_L g35 ( 
.A1(n_36),
.A2(n_37),
.B(n_40),
.C(n_42),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_38),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g42 ( 
.A(n_43),
.B(n_45),
.Y(n_42)
);

INVx1_ASAP7_75t_SL g43 ( 
.A(n_44),
.Y(n_43)
);

CKINVDCx16_ASAP7_75t_R g50 ( 
.A(n_51),
.Y(n_50)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_53),
.Y(n_52)
);


endmodule