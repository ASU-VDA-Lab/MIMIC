module fake_jpeg_2763_n_476 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_476);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_476;

wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_377;
wire n_291;
wire n_236;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_17;
wire n_431;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_415;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_48;
wire n_465;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_221;
wire n_256;
wire n_454;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_349;
wire n_21;
wire n_288;
wire n_393;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_429;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_474;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_305;
wire n_161;
wire n_441;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_389;
wire n_457;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_384;
wire n_168;
wire n_459;
wire n_274;
wire n_24;
wire n_467;
wire n_269;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_473;
wire n_45;
wire n_337;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_199;
wire n_260;
wire n_413;
wire n_275;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_472;
wire n_279;
wire n_154;
wire n_205;
wire n_379;
wire n_114;
wire n_444;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_469;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_183;
wire n_409;
wire n_249;
wire n_412;
wire n_217;
wire n_471;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_391;
wire n_209;
wire n_22;
wire n_138;
wire n_402;
wire n_438;
wire n_475;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

INVx2_ASAP7_75t_L g16 ( 
.A(n_8),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_5),
.Y(n_17)
);

INVx4_ASAP7_75t_L g18 ( 
.A(n_4),
.Y(n_18)
);

BUFx5_ASAP7_75t_L g19 ( 
.A(n_0),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_13),
.Y(n_20)
);

INVx6_ASAP7_75t_SL g21 ( 
.A(n_9),
.Y(n_21)
);

BUFx3_ASAP7_75t_L g22 ( 
.A(n_2),
.Y(n_22)
);

INVx8_ASAP7_75t_SL g23 ( 
.A(n_10),
.Y(n_23)
);

INVx6_ASAP7_75t_SL g24 ( 
.A(n_13),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_7),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_15),
.Y(n_26)
);

BUFx5_ASAP7_75t_L g27 ( 
.A(n_11),
.Y(n_27)
);

BUFx3_ASAP7_75t_L g28 ( 
.A(n_1),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_0),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_3),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_11),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_10),
.Y(n_32)
);

NOR2xp33_ASAP7_75t_L g33 ( 
.A(n_1),
.B(n_12),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_0),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_6),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_1),
.Y(n_36)
);

INVx8_ASAP7_75t_L g37 ( 
.A(n_6),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_9),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_2),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_13),
.Y(n_40)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_0),
.Y(n_41)
);

INVx2_ASAP7_75t_L g42 ( 
.A(n_12),
.Y(n_42)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_14),
.Y(n_43)
);

BUFx12f_ASAP7_75t_L g44 ( 
.A(n_9),
.Y(n_44)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_8),
.Y(n_45)
);

INVx6_ASAP7_75t_L g46 ( 
.A(n_2),
.Y(n_46)
);

BUFx16f_ASAP7_75t_L g47 ( 
.A(n_10),
.Y(n_47)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_15),
.Y(n_48)
);

BUFx12_ASAP7_75t_L g49 ( 
.A(n_15),
.Y(n_49)
);

BUFx16f_ASAP7_75t_L g50 ( 
.A(n_14),
.Y(n_50)
);

INVx3_ASAP7_75t_L g51 ( 
.A(n_18),
.Y(n_51)
);

INVx2_ASAP7_75t_SL g160 ( 
.A(n_51),
.Y(n_160)
);

INVx4_ASAP7_75t_SL g52 ( 
.A(n_21),
.Y(n_52)
);

INVx1_ASAP7_75t_SL g129 ( 
.A(n_52),
.Y(n_129)
);

INVx8_ASAP7_75t_L g53 ( 
.A(n_21),
.Y(n_53)
);

INVx5_ASAP7_75t_L g105 ( 
.A(n_53),
.Y(n_105)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_20),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g123 ( 
.A(n_54),
.Y(n_123)
);

INVx11_ASAP7_75t_L g55 ( 
.A(n_21),
.Y(n_55)
);

INVx4_ASAP7_75t_L g127 ( 
.A(n_55),
.Y(n_127)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_20),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g140 ( 
.A(n_56),
.Y(n_140)
);

INVx6_ASAP7_75t_L g57 ( 
.A(n_20),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g152 ( 
.A(n_57),
.Y(n_152)
);

INVx2_ASAP7_75t_SL g58 ( 
.A(n_24),
.Y(n_58)
);

INVx1_ASAP7_75t_SL g153 ( 
.A(n_58),
.Y(n_153)
);

INVx4_ASAP7_75t_L g59 ( 
.A(n_18),
.Y(n_59)
);

INVx3_ASAP7_75t_L g148 ( 
.A(n_59),
.Y(n_148)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_20),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g158 ( 
.A(n_60),
.Y(n_158)
);

BUFx5_ASAP7_75t_L g61 ( 
.A(n_24),
.Y(n_61)
);

INVx4_ASAP7_75t_L g136 ( 
.A(n_61),
.Y(n_136)
);

INVx2_ASAP7_75t_L g62 ( 
.A(n_16),
.Y(n_62)
);

INVx2_ASAP7_75t_L g121 ( 
.A(n_62),
.Y(n_121)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_26),
.Y(n_63)
);

INVx6_ASAP7_75t_L g117 ( 
.A(n_63),
.Y(n_117)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_17),
.Y(n_64)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_64),
.Y(n_114)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_17),
.Y(n_65)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_65),
.Y(n_115)
);

BUFx3_ASAP7_75t_L g66 ( 
.A(n_22),
.Y(n_66)
);

BUFx3_ASAP7_75t_L g104 ( 
.A(n_66),
.Y(n_104)
);

INVx3_ASAP7_75t_L g67 ( 
.A(n_18),
.Y(n_67)
);

BUFx2_ASAP7_75t_L g113 ( 
.A(n_67),
.Y(n_113)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_26),
.Y(n_68)
);

INVx6_ASAP7_75t_L g133 ( 
.A(n_68),
.Y(n_133)
);

INVx3_ASAP7_75t_L g69 ( 
.A(n_47),
.Y(n_69)
);

INVx2_ASAP7_75t_L g131 ( 
.A(n_69),
.Y(n_131)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_16),
.Y(n_70)
);

INVx2_ASAP7_75t_L g144 ( 
.A(n_70),
.Y(n_144)
);

BUFx5_ASAP7_75t_L g71 ( 
.A(n_24),
.Y(n_71)
);

BUFx3_ASAP7_75t_L g111 ( 
.A(n_71),
.Y(n_111)
);

INVx2_ASAP7_75t_L g72 ( 
.A(n_42),
.Y(n_72)
);

INVx2_ASAP7_75t_L g147 ( 
.A(n_72),
.Y(n_147)
);

INVx6_ASAP7_75t_L g73 ( 
.A(n_26),
.Y(n_73)
);

INVx8_ASAP7_75t_L g110 ( 
.A(n_73),
.Y(n_110)
);

BUFx6f_ASAP7_75t_L g74 ( 
.A(n_26),
.Y(n_74)
);

INVx8_ASAP7_75t_L g128 ( 
.A(n_74),
.Y(n_128)
);

BUFx3_ASAP7_75t_L g75 ( 
.A(n_22),
.Y(n_75)
);

BUFx3_ASAP7_75t_L g142 ( 
.A(n_75),
.Y(n_142)
);

BUFx3_ASAP7_75t_L g76 ( 
.A(n_22),
.Y(n_76)
);

INVx2_ASAP7_75t_L g149 ( 
.A(n_76),
.Y(n_149)
);

BUFx3_ASAP7_75t_L g77 ( 
.A(n_28),
.Y(n_77)
);

INVx2_ASAP7_75t_L g151 ( 
.A(n_77),
.Y(n_151)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_33),
.B(n_1),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_SL g150 ( 
.A(n_78),
.B(n_45),
.Y(n_150)
);

BUFx6f_ASAP7_75t_L g79 ( 
.A(n_34),
.Y(n_79)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_79),
.Y(n_126)
);

INVx2_ASAP7_75t_L g80 ( 
.A(n_42),
.Y(n_80)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_80),
.Y(n_116)
);

INVx2_ASAP7_75t_L g81 ( 
.A(n_44),
.Y(n_81)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_81),
.Y(n_119)
);

INVx2_ASAP7_75t_L g82 ( 
.A(n_44),
.Y(n_82)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_82),
.Y(n_122)
);

INVx5_ASAP7_75t_L g83 ( 
.A(n_37),
.Y(n_83)
);

CKINVDCx16_ASAP7_75t_R g103 ( 
.A(n_83),
.Y(n_103)
);

INVx3_ASAP7_75t_L g84 ( 
.A(n_47),
.Y(n_84)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_84),
.Y(n_138)
);

INVx11_ASAP7_75t_L g85 ( 
.A(n_44),
.Y(n_85)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_85),
.Y(n_139)
);

INVx3_ASAP7_75t_L g86 ( 
.A(n_47),
.Y(n_86)
);

AND2x2_ASAP7_75t_L g109 ( 
.A(n_86),
.B(n_88),
.Y(n_109)
);

CKINVDCx20_ASAP7_75t_R g87 ( 
.A(n_47),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g130 ( 
.A(n_87),
.B(n_90),
.Y(n_130)
);

INVx8_ASAP7_75t_L g88 ( 
.A(n_50),
.Y(n_88)
);

INVx2_ASAP7_75t_L g89 ( 
.A(n_44),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_SL g137 ( 
.A(n_89),
.B(n_91),
.Y(n_137)
);

BUFx3_ASAP7_75t_L g90 ( 
.A(n_28),
.Y(n_90)
);

INVx3_ASAP7_75t_L g91 ( 
.A(n_50),
.Y(n_91)
);

INVx8_ASAP7_75t_L g92 ( 
.A(n_50),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g132 ( 
.A(n_92),
.B(n_96),
.Y(n_132)
);

BUFx6f_ASAP7_75t_L g93 ( 
.A(n_34),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_L g107 ( 
.A(n_93),
.B(n_95),
.Y(n_107)
);

BUFx5_ASAP7_75t_L g94 ( 
.A(n_50),
.Y(n_94)
);

HAxp5_ASAP7_75t_SL g135 ( 
.A(n_94),
.B(n_102),
.CON(n_135),
.SN(n_135)
);

BUFx6f_ASAP7_75t_L g95 ( 
.A(n_34),
.Y(n_95)
);

CKINVDCx20_ASAP7_75t_R g96 ( 
.A(n_23),
.Y(n_96)
);

BUFx6f_ASAP7_75t_L g97 ( 
.A(n_34),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g134 ( 
.A(n_97),
.B(n_99),
.Y(n_134)
);

AOI21xp33_ASAP7_75t_SL g98 ( 
.A1(n_33),
.A2(n_2),
.B(n_3),
.Y(n_98)
);

MAJIxp5_ASAP7_75t_L g124 ( 
.A(n_98),
.B(n_29),
.C(n_30),
.Y(n_124)
);

BUFx6f_ASAP7_75t_L g99 ( 
.A(n_36),
.Y(n_99)
);

BUFx6f_ASAP7_75t_L g100 ( 
.A(n_36),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_L g146 ( 
.A(n_100),
.B(n_101),
.Y(n_146)
);

BUFx6f_ASAP7_75t_L g101 ( 
.A(n_36),
.Y(n_101)
);

HB1xp67_ASAP7_75t_L g102 ( 
.A(n_44),
.Y(n_102)
);

AOI22xp33_ASAP7_75t_L g106 ( 
.A1(n_54),
.A2(n_30),
.B1(n_48),
.B2(n_29),
.Y(n_106)
);

OAI22xp5_ASAP7_75t_L g187 ( 
.A1(n_106),
.A2(n_108),
.B1(n_112),
.B2(n_120),
.Y(n_187)
);

OAI22xp5_ASAP7_75t_L g108 ( 
.A1(n_57),
.A2(n_46),
.B1(n_36),
.B2(n_38),
.Y(n_108)
);

OAI22xp5_ASAP7_75t_L g112 ( 
.A1(n_73),
.A2(n_46),
.B1(n_38),
.B2(n_28),
.Y(n_112)
);

AOI22xp5_ASAP7_75t_SL g118 ( 
.A1(n_59),
.A2(n_38),
.B1(n_25),
.B2(n_31),
.Y(n_118)
);

OR2x2_ASAP7_75t_L g163 ( 
.A(n_118),
.B(n_150),
.Y(n_163)
);

OAI22xp5_ASAP7_75t_L g120 ( 
.A1(n_56),
.A2(n_46),
.B1(n_38),
.B2(n_48),
.Y(n_120)
);

AND2x2_ASAP7_75t_L g196 ( 
.A(n_124),
.B(n_3),
.Y(n_196)
);

OAI22xp33_ASAP7_75t_SL g125 ( 
.A1(n_60),
.A2(n_39),
.B1(n_32),
.B2(n_40),
.Y(n_125)
);

AOI22xp5_ASAP7_75t_L g204 ( 
.A1(n_125),
.A2(n_143),
.B1(n_159),
.B2(n_49),
.Y(n_204)
);

NOR2xp33_ASAP7_75t_L g141 ( 
.A(n_52),
.B(n_58),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_SL g175 ( 
.A(n_141),
.B(n_145),
.Y(n_175)
);

OAI22xp5_ASAP7_75t_L g143 ( 
.A1(n_63),
.A2(n_39),
.B1(n_32),
.B2(n_40),
.Y(n_143)
);

NOR2xp33_ASAP7_75t_L g145 ( 
.A(n_53),
.B(n_45),
.Y(n_145)
);

AOI22xp33_ASAP7_75t_L g154 ( 
.A1(n_68),
.A2(n_79),
.B1(n_101),
.B2(n_100),
.Y(n_154)
);

OAI22xp5_ASAP7_75t_SL g166 ( 
.A1(n_154),
.A2(n_25),
.B1(n_31),
.B2(n_35),
.Y(n_166)
);

AOI22xp33_ASAP7_75t_SL g155 ( 
.A1(n_55),
.A2(n_37),
.B1(n_23),
.B2(n_41),
.Y(n_155)
);

AOI22xp33_ASAP7_75t_SL g179 ( 
.A1(n_155),
.A2(n_85),
.B1(n_92),
.B2(n_88),
.Y(n_179)
);

OR2x2_ASAP7_75t_L g156 ( 
.A(n_102),
.B(n_35),
.Y(n_156)
);

CKINVDCx16_ASAP7_75t_R g173 ( 
.A(n_156),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_L g157 ( 
.A(n_99),
.B(n_43),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_L g170 ( 
.A(n_157),
.B(n_90),
.Y(n_170)
);

OAI22xp5_ASAP7_75t_L g159 ( 
.A1(n_74),
.A2(n_37),
.B1(n_43),
.B2(n_41),
.Y(n_159)
);

CKINVDCx20_ASAP7_75t_R g161 ( 
.A(n_109),
.Y(n_161)
);

NOR2xp33_ASAP7_75t_L g208 ( 
.A(n_161),
.B(n_168),
.Y(n_208)
);

INVx3_ASAP7_75t_SL g162 ( 
.A(n_128),
.Y(n_162)
);

BUFx2_ASAP7_75t_L g213 ( 
.A(n_162),
.Y(n_213)
);

AOI22xp33_ASAP7_75t_L g164 ( 
.A1(n_124),
.A2(n_97),
.B1(n_95),
.B2(n_93),
.Y(n_164)
);

OAI22xp5_ASAP7_75t_L g219 ( 
.A1(n_164),
.A2(n_174),
.B1(n_176),
.B2(n_177),
.Y(n_219)
);

INVx2_ASAP7_75t_L g165 ( 
.A(n_126),
.Y(n_165)
);

INVx2_ASAP7_75t_L g211 ( 
.A(n_165),
.Y(n_211)
);

AOI22xp5_ASAP7_75t_L g209 ( 
.A1(n_166),
.A2(n_199),
.B1(n_202),
.B2(n_204),
.Y(n_209)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_157),
.Y(n_167)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_167),
.Y(n_212)
);

CKINVDCx20_ASAP7_75t_R g168 ( 
.A(n_132),
.Y(n_168)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_126),
.Y(n_169)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_169),
.Y(n_217)
);

NOR2xp33_ASAP7_75t_L g210 ( 
.A(n_170),
.B(n_191),
.Y(n_210)
);

INVx2_ASAP7_75t_L g171 ( 
.A(n_149),
.Y(n_171)
);

INVx2_ASAP7_75t_L g224 ( 
.A(n_171),
.Y(n_224)
);

INVx2_ASAP7_75t_L g172 ( 
.A(n_149),
.Y(n_172)
);

INVx2_ASAP7_75t_L g229 ( 
.A(n_172),
.Y(n_229)
);

BUFx2_ASAP7_75t_L g174 ( 
.A(n_109),
.Y(n_174)
);

INVx2_ASAP7_75t_L g233 ( 
.A(n_174),
.Y(n_233)
);

NAND2xp5_ASAP7_75t_L g176 ( 
.A(n_107),
.B(n_77),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_L g222 ( 
.A(n_176),
.B(n_177),
.Y(n_222)
);

NAND2xp5_ASAP7_75t_L g177 ( 
.A(n_107),
.B(n_76),
.Y(n_177)
);

INVx2_ASAP7_75t_L g178 ( 
.A(n_151),
.Y(n_178)
);

INVx4_ASAP7_75t_L g227 ( 
.A(n_178),
.Y(n_227)
);

AOI22xp33_ASAP7_75t_SL g220 ( 
.A1(n_179),
.A2(n_188),
.B1(n_190),
.B2(n_195),
.Y(n_220)
);

NAND2xp5_ASAP7_75t_L g180 ( 
.A(n_134),
.B(n_146),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_L g232 ( 
.A(n_180),
.B(n_183),
.Y(n_232)
);

BUFx3_ASAP7_75t_L g181 ( 
.A(n_104),
.Y(n_181)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_181),
.Y(n_235)
);

INVx2_ASAP7_75t_L g182 ( 
.A(n_151),
.Y(n_182)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_182),
.Y(n_239)
);

NAND2xp5_ASAP7_75t_L g183 ( 
.A(n_134),
.B(n_75),
.Y(n_183)
);

BUFx5_ASAP7_75t_L g184 ( 
.A(n_131),
.Y(n_184)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_184),
.Y(n_243)
);

INVx3_ASAP7_75t_L g185 ( 
.A(n_127),
.Y(n_185)
);

INVxp67_ASAP7_75t_L g215 ( 
.A(n_185),
.Y(n_215)
);

MAJIxp5_ASAP7_75t_L g186 ( 
.A(n_114),
.B(n_66),
.C(n_27),
.Y(n_186)
);

MAJIxp5_ASAP7_75t_L g236 ( 
.A(n_186),
.B(n_196),
.C(n_136),
.Y(n_236)
);

AOI22xp33_ASAP7_75t_SL g188 ( 
.A1(n_109),
.A2(n_27),
.B1(n_19),
.B2(n_49),
.Y(n_188)
);

BUFx2_ASAP7_75t_L g189 ( 
.A(n_104),
.Y(n_189)
);

CKINVDCx16_ASAP7_75t_R g231 ( 
.A(n_189),
.Y(n_231)
);

AOI22xp33_ASAP7_75t_SL g190 ( 
.A1(n_160),
.A2(n_27),
.B1(n_19),
.B2(n_49),
.Y(n_190)
);

NAND2xp5_ASAP7_75t_L g191 ( 
.A(n_146),
.B(n_3),
.Y(n_191)
);

INVx3_ASAP7_75t_L g192 ( 
.A(n_127),
.Y(n_192)
);

NOR2xp33_ASAP7_75t_L g230 ( 
.A(n_192),
.B(n_194),
.Y(n_230)
);

HB1xp67_ASAP7_75t_L g193 ( 
.A(n_160),
.Y(n_193)
);

CKINVDCx16_ASAP7_75t_R g241 ( 
.A(n_193),
.Y(n_241)
);

NAND2xp5_ASAP7_75t_L g194 ( 
.A(n_115),
.B(n_156),
.Y(n_194)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_116),
.Y(n_195)
);

BUFx2_ASAP7_75t_L g197 ( 
.A(n_142),
.Y(n_197)
);

CKINVDCx20_ASAP7_75t_R g226 ( 
.A(n_197),
.Y(n_226)
);

INVx6_ASAP7_75t_L g198 ( 
.A(n_123),
.Y(n_198)
);

INVx8_ASAP7_75t_L g237 ( 
.A(n_198),
.Y(n_237)
);

OAI22xp5_ASAP7_75t_SL g199 ( 
.A1(n_118),
.A2(n_19),
.B1(n_49),
.B2(n_6),
.Y(n_199)
);

CKINVDCx20_ASAP7_75t_R g200 ( 
.A(n_130),
.Y(n_200)
);

AOI22xp33_ASAP7_75t_SL g223 ( 
.A1(n_200),
.A2(n_201),
.B1(n_203),
.B2(n_205),
.Y(n_223)
);

INVx2_ASAP7_75t_L g201 ( 
.A(n_121),
.Y(n_201)
);

OAI22xp5_ASAP7_75t_SL g202 ( 
.A1(n_137),
.A2(n_49),
.B1(n_5),
.B2(n_6),
.Y(n_202)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_121),
.Y(n_203)
);

CKINVDCx20_ASAP7_75t_R g205 ( 
.A(n_105),
.Y(n_205)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_144),
.Y(n_206)
);

AOI22xp33_ASAP7_75t_L g228 ( 
.A1(n_206),
.A2(n_207),
.B1(n_129),
.B2(n_153),
.Y(n_228)
);

INVx11_ASAP7_75t_L g207 ( 
.A(n_103),
.Y(n_207)
);

AOI22xp5_ASAP7_75t_L g214 ( 
.A1(n_187),
.A2(n_147),
.B1(n_144),
.B2(n_152),
.Y(n_214)
);

OAI22xp5_ASAP7_75t_SL g247 ( 
.A1(n_214),
.A2(n_216),
.B1(n_204),
.B2(n_169),
.Y(n_247)
);

AOI22xp5_ASAP7_75t_L g216 ( 
.A1(n_167),
.A2(n_147),
.B1(n_152),
.B2(n_110),
.Y(n_216)
);

OAI21xp5_ASAP7_75t_SL g218 ( 
.A1(n_161),
.A2(n_129),
.B(n_153),
.Y(n_218)
);

OAI21xp5_ASAP7_75t_SL g268 ( 
.A1(n_218),
.A2(n_196),
.B(n_195),
.Y(n_268)
);

AND2x2_ASAP7_75t_L g261 ( 
.A(n_219),
.B(n_225),
.Y(n_261)
);

AOI32xp33_ASAP7_75t_L g221 ( 
.A1(n_180),
.A2(n_136),
.A3(n_122),
.B1(n_119),
.B2(n_135),
.Y(n_221)
);

NOR2xp33_ASAP7_75t_L g245 ( 
.A(n_221),
.B(n_163),
.Y(n_245)
);

OAI22xp5_ASAP7_75t_SL g225 ( 
.A1(n_170),
.A2(n_117),
.B1(n_133),
.B2(n_158),
.Y(n_225)
);

INVxp67_ASAP7_75t_SL g260 ( 
.A(n_228),
.Y(n_260)
);

OAI22xp5_ASAP7_75t_L g234 ( 
.A1(n_183),
.A2(n_133),
.B1(n_117),
.B2(n_158),
.Y(n_234)
);

AOI22xp33_ASAP7_75t_L g262 ( 
.A1(n_234),
.A2(n_162),
.B1(n_140),
.B2(n_201),
.Y(n_262)
);

NOR2xp33_ASAP7_75t_SL g251 ( 
.A(n_236),
.B(n_186),
.Y(n_251)
);

O2A1O1Ixp33_ASAP7_75t_L g238 ( 
.A1(n_194),
.A2(n_135),
.B(n_111),
.C(n_139),
.Y(n_238)
);

OAI21xp5_ASAP7_75t_L g267 ( 
.A1(n_238),
.A2(n_242),
.B(n_202),
.Y(n_267)
);

AOI22xp33_ASAP7_75t_L g240 ( 
.A1(n_173),
.A2(n_113),
.B1(n_148),
.B2(n_123),
.Y(n_240)
);

OAI22xp33_ASAP7_75t_SL g250 ( 
.A1(n_240),
.A2(n_207),
.B1(n_165),
.B2(n_113),
.Y(n_250)
);

O2A1O1Ixp33_ASAP7_75t_L g242 ( 
.A1(n_163),
.A2(n_111),
.B(n_138),
.C(n_142),
.Y(n_242)
);

INVxp33_ASAP7_75t_L g244 ( 
.A(n_223),
.Y(n_244)
);

NOR2xp33_ASAP7_75t_L g276 ( 
.A(n_244),
.B(n_253),
.Y(n_276)
);

OAI21xp5_ASAP7_75t_SL g287 ( 
.A1(n_245),
.A2(n_254),
.B(n_268),
.Y(n_287)
);

INVx2_ASAP7_75t_L g246 ( 
.A(n_211),
.Y(n_246)
);

INVx2_ASAP7_75t_L g293 ( 
.A(n_246),
.Y(n_293)
);

AOI22xp5_ASAP7_75t_L g295 ( 
.A1(n_247),
.A2(n_248),
.B1(n_166),
.B2(n_224),
.Y(n_295)
);

OAI22xp5_ASAP7_75t_SL g248 ( 
.A1(n_209),
.A2(n_232),
.B1(n_222),
.B2(n_214),
.Y(n_248)
);

NAND2xp5_ASAP7_75t_L g249 ( 
.A(n_232),
.B(n_191),
.Y(n_249)
);

NAND2xp5_ASAP7_75t_L g275 ( 
.A(n_249),
.B(n_257),
.Y(n_275)
);

AOI22xp33_ASAP7_75t_L g281 ( 
.A1(n_250),
.A2(n_213),
.B1(n_162),
.B2(n_226),
.Y(n_281)
);

INVxp67_ASAP7_75t_L g300 ( 
.A(n_251),
.Y(n_300)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_217),
.Y(n_252)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_252),
.Y(n_282)
);

CKINVDCx20_ASAP7_75t_R g253 ( 
.A(n_215),
.Y(n_253)
);

NAND2xp67_ASAP7_75t_L g254 ( 
.A(n_238),
.B(n_185),
.Y(n_254)
);

INVxp67_ASAP7_75t_L g255 ( 
.A(n_208),
.Y(n_255)
);

NOR2xp33_ASAP7_75t_L g284 ( 
.A(n_255),
.B(n_263),
.Y(n_284)
);

NOR2xp33_ASAP7_75t_SL g256 ( 
.A(n_208),
.B(n_230),
.Y(n_256)
);

NAND2xp5_ASAP7_75t_SL g304 ( 
.A(n_256),
.B(n_273),
.Y(n_304)
);

NAND2xp5_ASAP7_75t_SL g257 ( 
.A(n_222),
.B(n_175),
.Y(n_257)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_217),
.Y(n_258)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_258),
.Y(n_288)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_211),
.Y(n_259)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_259),
.Y(n_297)
);

OAI22xp5_ASAP7_75t_L g283 ( 
.A1(n_262),
.A2(n_270),
.B1(n_216),
.B2(n_213),
.Y(n_283)
);

INVxp67_ASAP7_75t_L g263 ( 
.A(n_221),
.Y(n_263)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_239),
.Y(n_264)
);

NOR2xp33_ASAP7_75t_L g298 ( 
.A(n_264),
.B(n_266),
.Y(n_298)
);

AOI21xp5_ASAP7_75t_L g265 ( 
.A1(n_218),
.A2(n_199),
.B(n_192),
.Y(n_265)
);

AOI21xp5_ASAP7_75t_L g286 ( 
.A1(n_265),
.A2(n_242),
.B(n_226),
.Y(n_286)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_239),
.Y(n_266)
);

INVxp67_ASAP7_75t_L g303 ( 
.A(n_267),
.Y(n_303)
);

INVx1_ASAP7_75t_SL g269 ( 
.A(n_233),
.Y(n_269)
);

CKINVDCx14_ASAP7_75t_R g289 ( 
.A(n_269),
.Y(n_289)
);

AOI22xp33_ASAP7_75t_L g270 ( 
.A1(n_212),
.A2(n_206),
.B1(n_203),
.B2(n_140),
.Y(n_270)
);

BUFx8_ASAP7_75t_L g271 ( 
.A(n_213),
.Y(n_271)
);

CKINVDCx20_ASAP7_75t_R g279 ( 
.A(n_271),
.Y(n_279)
);

NAND2xp5_ASAP7_75t_L g272 ( 
.A(n_210),
.B(n_196),
.Y(n_272)
);

NAND2xp5_ASAP7_75t_L g277 ( 
.A(n_272),
.B(n_274),
.Y(n_277)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_233),
.Y(n_273)
);

NOR2xp33_ASAP7_75t_L g274 ( 
.A(n_230),
.B(n_171),
.Y(n_274)
);

XOR2xp5_ASAP7_75t_L g278 ( 
.A(n_251),
.B(n_236),
.Y(n_278)
);

MAJIxp5_ASAP7_75t_L g307 ( 
.A(n_278),
.B(n_299),
.C(n_252),
.Y(n_307)
);

OAI22xp5_ASAP7_75t_SL g280 ( 
.A1(n_261),
.A2(n_209),
.B1(n_212),
.B2(n_210),
.Y(n_280)
);

AOI22xp5_ASAP7_75t_L g310 ( 
.A1(n_280),
.A2(n_285),
.B1(n_290),
.B2(n_295),
.Y(n_310)
);

AOI22xp33_ASAP7_75t_L g329 ( 
.A1(n_281),
.A2(n_283),
.B1(n_271),
.B2(n_227),
.Y(n_329)
);

OAI22xp5_ASAP7_75t_SL g285 ( 
.A1(n_261),
.A2(n_220),
.B1(n_219),
.B2(n_238),
.Y(n_285)
);

OAI21xp5_ASAP7_75t_SL g317 ( 
.A1(n_286),
.A2(n_294),
.B(n_260),
.Y(n_317)
);

OAI22xp5_ASAP7_75t_SL g290 ( 
.A1(n_261),
.A2(n_242),
.B1(n_234),
.B2(n_225),
.Y(n_290)
);

CKINVDCx20_ASAP7_75t_R g291 ( 
.A(n_274),
.Y(n_291)
);

NOR2xp33_ASAP7_75t_L g306 ( 
.A(n_291),
.B(n_256),
.Y(n_306)
);

NOR2x1_ASAP7_75t_SL g292 ( 
.A(n_245),
.B(n_268),
.Y(n_292)
);

AO21x1_ASAP7_75t_L g313 ( 
.A1(n_292),
.A2(n_267),
.B(n_254),
.Y(n_313)
);

OAI21xp5_ASAP7_75t_SL g294 ( 
.A1(n_265),
.A2(n_235),
.B(n_105),
.Y(n_294)
);

NAND2xp5_ASAP7_75t_L g296 ( 
.A(n_249),
.B(n_229),
.Y(n_296)
);

NAND2xp5_ASAP7_75t_L g318 ( 
.A(n_296),
.B(n_302),
.Y(n_318)
);

XNOR2xp5_ASAP7_75t_L g299 ( 
.A(n_272),
.B(n_235),
.Y(n_299)
);

AOI22xp5_ASAP7_75t_L g301 ( 
.A1(n_261),
.A2(n_237),
.B1(n_128),
.B2(n_229),
.Y(n_301)
);

OAI22xp5_ASAP7_75t_SL g319 ( 
.A1(n_301),
.A2(n_262),
.B1(n_270),
.B2(n_260),
.Y(n_319)
);

NAND2xp5_ASAP7_75t_L g302 ( 
.A(n_248),
.B(n_224),
.Y(n_302)
);

CKINVDCx20_ASAP7_75t_R g305 ( 
.A(n_298),
.Y(n_305)
);

NAND2xp5_ASAP7_75t_L g333 ( 
.A(n_305),
.B(n_311),
.Y(n_333)
);

OR2x2_ASAP7_75t_L g348 ( 
.A(n_306),
.B(n_309),
.Y(n_348)
);

XNOR2xp5_ASAP7_75t_SL g354 ( 
.A(n_307),
.B(n_284),
.Y(n_354)
);

AOI32xp33_ASAP7_75t_L g308 ( 
.A1(n_303),
.A2(n_267),
.A3(n_254),
.B1(n_253),
.B2(n_258),
.Y(n_308)
);

NOR2xp33_ASAP7_75t_L g353 ( 
.A(n_308),
.B(n_331),
.Y(n_353)
);

NOR2xp33_ASAP7_75t_L g309 ( 
.A(n_291),
.B(n_259),
.Y(n_309)
);

CKINVDCx20_ASAP7_75t_R g311 ( 
.A(n_298),
.Y(n_311)
);

MAJIxp5_ASAP7_75t_L g312 ( 
.A(n_278),
.B(n_257),
.C(n_266),
.Y(n_312)
);

MAJIxp5_ASAP7_75t_L g336 ( 
.A(n_312),
.B(n_307),
.C(n_314),
.Y(n_336)
);

OAI21xp5_ASAP7_75t_SL g346 ( 
.A1(n_313),
.A2(n_317),
.B(n_321),
.Y(n_346)
);

MAJx2_ASAP7_75t_L g314 ( 
.A(n_278),
.B(n_247),
.C(n_264),
.Y(n_314)
);

XNOR2xp5_ASAP7_75t_L g342 ( 
.A(n_314),
.B(n_280),
.Y(n_342)
);

CKINVDCx20_ASAP7_75t_R g315 ( 
.A(n_289),
.Y(n_315)
);

NAND2xp5_ASAP7_75t_L g345 ( 
.A(n_315),
.B(n_326),
.Y(n_345)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_282),
.Y(n_316)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_316),
.Y(n_335)
);

AOI22xp5_ASAP7_75t_L g340 ( 
.A1(n_319),
.A2(n_332),
.B1(n_283),
.B2(n_290),
.Y(n_340)
);

NOR2xp33_ASAP7_75t_L g320 ( 
.A(n_300),
.B(n_304),
.Y(n_320)
);

NOR2xp33_ASAP7_75t_SL g356 ( 
.A(n_320),
.B(n_327),
.Y(n_356)
);

OAI21xp5_ASAP7_75t_L g321 ( 
.A1(n_287),
.A2(n_269),
.B(n_273),
.Y(n_321)
);

NAND2xp5_ASAP7_75t_L g322 ( 
.A(n_296),
.B(n_246),
.Y(n_322)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_322),
.Y(n_341)
);

INVx3_ASAP7_75t_SL g323 ( 
.A(n_293),
.Y(n_323)
);

INVx2_ASAP7_75t_L g360 ( 
.A(n_323),
.Y(n_360)
);

INVx2_ASAP7_75t_L g324 ( 
.A(n_293),
.Y(n_324)
);

INVx1_ASAP7_75t_L g343 ( 
.A(n_324),
.Y(n_343)
);

OAI21xp5_ASAP7_75t_SL g325 ( 
.A1(n_287),
.A2(n_269),
.B(n_271),
.Y(n_325)
);

AOI21xp5_ASAP7_75t_L g344 ( 
.A1(n_325),
.A2(n_286),
.B(n_294),
.Y(n_344)
);

CKINVDCx20_ASAP7_75t_R g326 ( 
.A(n_289),
.Y(n_326)
);

CKINVDCx20_ASAP7_75t_R g327 ( 
.A(n_304),
.Y(n_327)
);

CKINVDCx20_ASAP7_75t_R g334 ( 
.A(n_327),
.Y(n_334)
);

AOI22xp5_ASAP7_75t_L g328 ( 
.A1(n_285),
.A2(n_250),
.B1(n_271),
.B2(n_237),
.Y(n_328)
);

OAI22xp5_ASAP7_75t_L g347 ( 
.A1(n_328),
.A2(n_329),
.B1(n_281),
.B2(n_301),
.Y(n_347)
);

NAND2xp5_ASAP7_75t_L g330 ( 
.A(n_275),
.B(n_271),
.Y(n_330)
);

INVx1_ASAP7_75t_L g355 ( 
.A(n_330),
.Y(n_355)
);

INVxp67_ASAP7_75t_L g331 ( 
.A(n_292),
.Y(n_331)
);

OAI22xp5_ASAP7_75t_SL g332 ( 
.A1(n_295),
.A2(n_237),
.B1(n_198),
.B2(n_231),
.Y(n_332)
);

XNOR2xp5_ASAP7_75t_L g374 ( 
.A(n_336),
.B(n_342),
.Y(n_374)
);

XOR2xp5_ASAP7_75t_L g337 ( 
.A(n_312),
.B(n_299),
.Y(n_337)
);

XOR2xp5_ASAP7_75t_L g368 ( 
.A(n_337),
.B(n_354),
.Y(n_368)
);

CKINVDCx20_ASAP7_75t_R g338 ( 
.A(n_309),
.Y(n_338)
);

NAND2xp5_ASAP7_75t_SL g367 ( 
.A(n_338),
.B(n_349),
.Y(n_367)
);

MAJIxp5_ASAP7_75t_L g339 ( 
.A(n_314),
.B(n_299),
.C(n_277),
.Y(n_339)
);

MAJIxp5_ASAP7_75t_L g373 ( 
.A(n_339),
.B(n_350),
.C(n_357),
.Y(n_373)
);

OAI22xp33_ASAP7_75t_SL g372 ( 
.A1(n_340),
.A2(n_352),
.B1(n_318),
.B2(n_326),
.Y(n_372)
);

AOI21xp5_ASAP7_75t_L g364 ( 
.A1(n_344),
.A2(n_308),
.B(n_317),
.Y(n_364)
);

OAI22xp5_ASAP7_75t_L g362 ( 
.A1(n_347),
.A2(n_351),
.B1(n_356),
.B2(n_305),
.Y(n_362)
);

CKINVDCx16_ASAP7_75t_R g349 ( 
.A(n_320),
.Y(n_349)
);

MAJIxp5_ASAP7_75t_L g350 ( 
.A(n_321),
.B(n_277),
.C(n_275),
.Y(n_350)
);

OAI22xp5_ASAP7_75t_L g351 ( 
.A1(n_310),
.A2(n_284),
.B1(n_302),
.B2(n_301),
.Y(n_351)
);

CKINVDCx20_ASAP7_75t_R g352 ( 
.A(n_330),
.Y(n_352)
);

MAJIxp5_ASAP7_75t_L g357 ( 
.A(n_306),
.B(n_288),
.C(n_282),
.Y(n_357)
);

INVx1_ASAP7_75t_L g358 ( 
.A(n_322),
.Y(n_358)
);

INVx1_ASAP7_75t_L g361 ( 
.A(n_358),
.Y(n_361)
);

XNOR2xp5_ASAP7_75t_L g359 ( 
.A(n_313),
.B(n_288),
.Y(n_359)
);

XOR2xp5_ASAP7_75t_L g376 ( 
.A(n_359),
.B(n_313),
.Y(n_376)
);

AOI22xp5_ASAP7_75t_L g390 ( 
.A1(n_362),
.A2(n_370),
.B1(n_378),
.B2(n_384),
.Y(n_390)
);

NOR2xp33_ASAP7_75t_L g363 ( 
.A(n_357),
.B(n_311),
.Y(n_363)
);

NOR2xp33_ASAP7_75t_SL g401 ( 
.A(n_363),
.B(n_227),
.Y(n_401)
);

OAI21xp5_ASAP7_75t_SL g395 ( 
.A1(n_364),
.A2(n_385),
.B(n_341),
.Y(n_395)
);

CKINVDCx16_ASAP7_75t_R g365 ( 
.A(n_345),
.Y(n_365)
);

NAND2xp5_ASAP7_75t_L g389 ( 
.A(n_365),
.B(n_366),
.Y(n_389)
);

CKINVDCx20_ASAP7_75t_R g366 ( 
.A(n_345),
.Y(n_366)
);

AOI22xp5_ASAP7_75t_SL g369 ( 
.A1(n_353),
.A2(n_333),
.B1(n_334),
.B2(n_355),
.Y(n_369)
);

OAI22xp5_ASAP7_75t_SL g391 ( 
.A1(n_369),
.A2(n_358),
.B1(n_341),
.B2(n_335),
.Y(n_391)
);

OAI22xp5_ASAP7_75t_SL g370 ( 
.A1(n_340),
.A2(n_310),
.B1(n_328),
.B2(n_318),
.Y(n_370)
);

INVx1_ASAP7_75t_L g371 ( 
.A(n_333),
.Y(n_371)
);

INVx1_ASAP7_75t_L g392 ( 
.A(n_371),
.Y(n_392)
);

INVx1_ASAP7_75t_L g405 ( 
.A(n_372),
.Y(n_405)
);

XNOR2x1_ASAP7_75t_L g375 ( 
.A(n_359),
.B(n_350),
.Y(n_375)
);

XOR2xp5_ASAP7_75t_L g397 ( 
.A(n_375),
.B(n_368),
.Y(n_397)
);

XNOR2xp5_ASAP7_75t_L g387 ( 
.A(n_376),
.B(n_346),
.Y(n_387)
);

OAI22xp5_ASAP7_75t_L g377 ( 
.A1(n_348),
.A2(n_315),
.B1(n_316),
.B2(n_276),
.Y(n_377)
);

NAND2xp5_ASAP7_75t_L g393 ( 
.A(n_377),
.B(n_382),
.Y(n_393)
);

OAI22xp5_ASAP7_75t_SL g378 ( 
.A1(n_334),
.A2(n_325),
.B1(n_276),
.B2(n_323),
.Y(n_378)
);

MAJIxp5_ASAP7_75t_L g379 ( 
.A(n_336),
.B(n_297),
.C(n_241),
.Y(n_379)
);

MAJIxp5_ASAP7_75t_L g386 ( 
.A(n_379),
.B(n_380),
.C(n_381),
.Y(n_386)
);

MAJIxp5_ASAP7_75t_L g380 ( 
.A(n_337),
.B(n_354),
.C(n_339),
.Y(n_380)
);

MAJIxp5_ASAP7_75t_L g381 ( 
.A(n_342),
.B(n_297),
.C(n_241),
.Y(n_381)
);

INVx2_ASAP7_75t_L g382 ( 
.A(n_360),
.Y(n_382)
);

MAJIxp5_ASAP7_75t_L g383 ( 
.A(n_348),
.B(n_332),
.C(n_197),
.Y(n_383)
);

MAJIxp5_ASAP7_75t_L g388 ( 
.A(n_383),
.B(n_360),
.C(n_343),
.Y(n_388)
);

OAI22xp5_ASAP7_75t_SL g384 ( 
.A1(n_352),
.A2(n_323),
.B1(n_319),
.B2(n_324),
.Y(n_384)
);

OAI21xp5_ASAP7_75t_L g385 ( 
.A1(n_346),
.A2(n_344),
.B(n_355),
.Y(n_385)
);

XNOR2xp5_ASAP7_75t_SL g411 ( 
.A(n_387),
.B(n_397),
.Y(n_411)
);

XOR2xp5_ASAP7_75t_L g422 ( 
.A(n_388),
.B(n_131),
.Y(n_422)
);

AOI22xp5_ASAP7_75t_L g415 ( 
.A1(n_391),
.A2(n_402),
.B1(n_378),
.B2(n_383),
.Y(n_415)
);

CKINVDCx16_ASAP7_75t_R g394 ( 
.A(n_367),
.Y(n_394)
);

NAND2xp5_ASAP7_75t_L g407 ( 
.A(n_394),
.B(n_396),
.Y(n_407)
);

OAI21xp5_ASAP7_75t_SL g406 ( 
.A1(n_395),
.A2(n_364),
.B(n_385),
.Y(n_406)
);

NAND2xp5_ASAP7_75t_SL g396 ( 
.A(n_373),
.B(n_335),
.Y(n_396)
);

XNOR2xp5_ASAP7_75t_L g398 ( 
.A(n_380),
.B(n_343),
.Y(n_398)
);

NAND2xp5_ASAP7_75t_L g417 ( 
.A(n_398),
.B(n_399),
.Y(n_417)
);

MAJIxp5_ASAP7_75t_L g399 ( 
.A(n_379),
.B(n_279),
.C(n_243),
.Y(n_399)
);

AOI22xp5_ASAP7_75t_L g400 ( 
.A1(n_370),
.A2(n_279),
.B1(n_231),
.B2(n_243),
.Y(n_400)
);

OAI22xp5_ASAP7_75t_SL g412 ( 
.A1(n_400),
.A2(n_361),
.B1(n_382),
.B2(n_384),
.Y(n_412)
);

INVx1_ASAP7_75t_L g413 ( 
.A(n_401),
.Y(n_413)
);

OAI22xp5_ASAP7_75t_SL g402 ( 
.A1(n_369),
.A2(n_227),
.B1(n_181),
.B2(n_189),
.Y(n_402)
);

XOR2xp5_ASAP7_75t_L g403 ( 
.A(n_375),
.B(n_182),
.Y(n_403)
);

XOR2xp5_ASAP7_75t_L g414 ( 
.A(n_403),
.B(n_404),
.Y(n_414)
);

XOR2xp5_ASAP7_75t_L g404 ( 
.A(n_373),
.B(n_178),
.Y(n_404)
);

OAI21xp5_ASAP7_75t_L g426 ( 
.A1(n_406),
.A2(n_390),
.B(n_387),
.Y(n_426)
);

MAJIxp5_ASAP7_75t_L g408 ( 
.A(n_398),
.B(n_374),
.C(n_368),
.Y(n_408)
);

NAND2xp5_ASAP7_75t_L g433 ( 
.A(n_408),
.B(n_409),
.Y(n_433)
);

NOR2xp33_ASAP7_75t_L g409 ( 
.A(n_404),
.B(n_371),
.Y(n_409)
);

FAx1_ASAP7_75t_SL g410 ( 
.A(n_391),
.B(n_376),
.CI(n_366),
.CON(n_410),
.SN(n_410)
);

NOR2x1_ASAP7_75t_L g431 ( 
.A(n_410),
.B(n_392),
.Y(n_431)
);

AOI22xp5_ASAP7_75t_L g434 ( 
.A1(n_412),
.A2(n_402),
.B1(n_400),
.B2(n_110),
.Y(n_434)
);

OAI22xp5_ASAP7_75t_SL g436 ( 
.A1(n_415),
.A2(n_4),
.B1(n_5),
.B2(n_7),
.Y(n_436)
);

XOR2xp5_ASAP7_75t_L g416 ( 
.A(n_397),
.B(n_374),
.Y(n_416)
);

XNOR2xp5_ASAP7_75t_L g427 ( 
.A(n_416),
.B(n_422),
.Y(n_427)
);

NOR2xp33_ASAP7_75t_L g418 ( 
.A(n_405),
.B(n_381),
.Y(n_418)
);

INVx1_ASAP7_75t_L g424 ( 
.A(n_418),
.Y(n_424)
);

INVx1_ASAP7_75t_L g419 ( 
.A(n_389),
.Y(n_419)
);

INVx1_ASAP7_75t_L g425 ( 
.A(n_419),
.Y(n_425)
);

OAI21xp5_ASAP7_75t_SL g420 ( 
.A1(n_395),
.A2(n_361),
.B(n_172),
.Y(n_420)
);

OAI21xp5_ASAP7_75t_SL g437 ( 
.A1(n_420),
.A2(n_4),
.B(n_5),
.Y(n_437)
);

MAJIxp5_ASAP7_75t_L g421 ( 
.A(n_386),
.B(n_399),
.C(n_403),
.Y(n_421)
);

NAND2xp5_ASAP7_75t_SL g432 ( 
.A(n_421),
.B(n_408),
.Y(n_432)
);

MAJIxp5_ASAP7_75t_L g423 ( 
.A(n_421),
.B(n_386),
.C(n_388),
.Y(n_423)
);

NAND2xp5_ASAP7_75t_L g441 ( 
.A(n_423),
.B(n_429),
.Y(n_441)
);

OAI21xp5_ASAP7_75t_L g446 ( 
.A1(n_426),
.A2(n_431),
.B(n_406),
.Y(n_446)
);

XOR2xp5_ASAP7_75t_L g428 ( 
.A(n_411),
.B(n_390),
.Y(n_428)
);

XNOR2xp5_ASAP7_75t_L g450 ( 
.A(n_428),
.B(n_437),
.Y(n_450)
);

XNOR2xp5_ASAP7_75t_L g429 ( 
.A(n_417),
.B(n_393),
.Y(n_429)
);

INVx1_ASAP7_75t_L g430 ( 
.A(n_407),
.Y(n_430)
);

INVx1_ASAP7_75t_L g443 ( 
.A(n_430),
.Y(n_443)
);

NOR2xp33_ASAP7_75t_SL g440 ( 
.A(n_432),
.B(n_413),
.Y(n_440)
);

AOI22xp5_ASAP7_75t_L g445 ( 
.A1(n_434),
.A2(n_436),
.B1(n_415),
.B2(n_410),
.Y(n_445)
);

MAJIxp5_ASAP7_75t_L g435 ( 
.A(n_416),
.B(n_148),
.C(n_184),
.Y(n_435)
);

NAND2xp5_ASAP7_75t_L g442 ( 
.A(n_435),
.B(n_411),
.Y(n_442)
);

AOI21xp5_ASAP7_75t_L g438 ( 
.A1(n_423),
.A2(n_433),
.B(n_431),
.Y(n_438)
);

AOI21xp5_ASAP7_75t_L g451 ( 
.A1(n_438),
.A2(n_446),
.B(n_427),
.Y(n_451)
);

MAJIxp5_ASAP7_75t_L g439 ( 
.A(n_428),
.B(n_414),
.C(n_422),
.Y(n_439)
);

NAND2xp5_ASAP7_75t_L g452 ( 
.A(n_439),
.B(n_444),
.Y(n_452)
);

NAND2xp5_ASAP7_75t_SL g455 ( 
.A(n_440),
.B(n_447),
.Y(n_455)
);

INVx1_ASAP7_75t_L g454 ( 
.A(n_442),
.Y(n_454)
);

NAND2xp5_ASAP7_75t_L g444 ( 
.A(n_429),
.B(n_412),
.Y(n_444)
);

NAND2xp5_ASAP7_75t_L g458 ( 
.A(n_445),
.B(n_448),
.Y(n_458)
);

NOR2xp33_ASAP7_75t_SL g447 ( 
.A(n_424),
.B(n_410),
.Y(n_447)
);

NAND2xp5_ASAP7_75t_SL g448 ( 
.A(n_425),
.B(n_426),
.Y(n_448)
);

NAND2xp5_ASAP7_75t_L g449 ( 
.A(n_436),
.B(n_414),
.Y(n_449)
);

NAND2xp5_ASAP7_75t_L g459 ( 
.A(n_449),
.B(n_8),
.Y(n_459)
);

AOI21x1_ASAP7_75t_L g465 ( 
.A1(n_451),
.A2(n_457),
.B(n_11),
.Y(n_465)
);

OAI21xp5_ASAP7_75t_SL g453 ( 
.A1(n_446),
.A2(n_434),
.B(n_427),
.Y(n_453)
);

OAI21xp5_ASAP7_75t_L g461 ( 
.A1(n_453),
.A2(n_450),
.B(n_439),
.Y(n_461)
);

MAJIxp5_ASAP7_75t_L g456 ( 
.A(n_441),
.B(n_435),
.C(n_7),
.Y(n_456)
);

OR2x2_ASAP7_75t_L g466 ( 
.A(n_456),
.B(n_459),
.Y(n_466)
);

AOI21xp5_ASAP7_75t_L g457 ( 
.A1(n_443),
.A2(n_4),
.B(n_7),
.Y(n_457)
);

NAND2xp5_ASAP7_75t_L g460 ( 
.A(n_445),
.B(n_8),
.Y(n_460)
);

NAND2xp5_ASAP7_75t_SL g464 ( 
.A(n_460),
.B(n_11),
.Y(n_464)
);

OAI21x1_ASAP7_75t_L g469 ( 
.A1(n_461),
.A2(n_462),
.B(n_463),
.Y(n_469)
);

OAI21xp5_ASAP7_75t_L g462 ( 
.A1(n_451),
.A2(n_450),
.B(n_10),
.Y(n_462)
);

AND2x2_ASAP7_75t_L g463 ( 
.A(n_455),
.B(n_9),
.Y(n_463)
);

NOR2xp33_ASAP7_75t_L g467 ( 
.A(n_464),
.B(n_465),
.Y(n_467)
);

NAND2xp5_ASAP7_75t_SL g468 ( 
.A(n_466),
.B(n_454),
.Y(n_468)
);

NOR2xp33_ASAP7_75t_L g472 ( 
.A(n_468),
.B(n_470),
.Y(n_472)
);

NOR2xp33_ASAP7_75t_L g470 ( 
.A(n_463),
.B(n_452),
.Y(n_470)
);

AOI321xp33_ASAP7_75t_L g471 ( 
.A1(n_469),
.A2(n_458),
.A3(n_456),
.B1(n_14),
.B2(n_15),
.C(n_13),
.Y(n_471)
);

INVxp67_ASAP7_75t_L g473 ( 
.A(n_471),
.Y(n_473)
);

NAND2xp5_ASAP7_75t_SL g474 ( 
.A(n_473),
.B(n_472),
.Y(n_474)
);

OAI21xp33_ASAP7_75t_L g475 ( 
.A1(n_474),
.A2(n_467),
.B(n_12),
.Y(n_475)
);

XOR2xp5_ASAP7_75t_L g476 ( 
.A(n_475),
.B(n_12),
.Y(n_476)
);


endmodule