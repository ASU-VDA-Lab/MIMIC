module fake_ariane_1427_n_1236 (n_83, n_8, n_56, n_60, n_170, n_190, n_160, n_64, n_179, n_180, n_119, n_124, n_167, n_90, n_38, n_47, n_110, n_153, n_18, n_86, n_75, n_89, n_67, n_176, n_149, n_34, n_158, n_172, n_69, n_95, n_175, n_92, n_143, n_183, n_150, n_98, n_74, n_113, n_114, n_33, n_19, n_40, n_181, n_152, n_120, n_169, n_106, n_12, n_53, n_173, n_111, n_21, n_115, n_133, n_66, n_71, n_24, n_7, n_109, n_96, n_156, n_49, n_20, n_174, n_100, n_17, n_50, n_187, n_132, n_62, n_147, n_51, n_166, n_76, n_103, n_79, n_26, n_3, n_46, n_0, n_84, n_36, n_91, n_159, n_107, n_189, n_72, n_105, n_128, n_44, n_30, n_82, n_178, n_31, n_42, n_57, n_131, n_70, n_10, n_117, n_139, n_165, n_85, n_130, n_144, n_6, n_48, n_94, n_101, n_4, n_134, n_188, n_185, n_2, n_32, n_37, n_58, n_65, n_123, n_9, n_138, n_112, n_45, n_162, n_11, n_129, n_126, n_137, n_122, n_148, n_164, n_52, n_157, n_184, n_177, n_135, n_73, n_77, n_171, n_15, n_118, n_93, n_121, n_23, n_61, n_108, n_102, n_182, n_125, n_22, n_168, n_43, n_1, n_81, n_87, n_13, n_27, n_29, n_41, n_140, n_55, n_151, n_136, n_28, n_80, n_146, n_97, n_154, n_142, n_161, n_14, n_163, n_88, n_186, n_141, n_68, n_116, n_104, n_145, n_78, n_39, n_59, n_63, n_99, n_16, n_5, n_155, n_127, n_35, n_54, n_25, n_1236);

input n_83;
input n_8;
input n_56;
input n_60;
input n_170;
input n_190;
input n_160;
input n_64;
input n_179;
input n_180;
input n_119;
input n_124;
input n_167;
input n_90;
input n_38;
input n_47;
input n_110;
input n_153;
input n_18;
input n_86;
input n_75;
input n_89;
input n_67;
input n_176;
input n_149;
input n_34;
input n_158;
input n_172;
input n_69;
input n_95;
input n_175;
input n_92;
input n_143;
input n_183;
input n_150;
input n_98;
input n_74;
input n_113;
input n_114;
input n_33;
input n_19;
input n_40;
input n_181;
input n_152;
input n_120;
input n_169;
input n_106;
input n_12;
input n_53;
input n_173;
input n_111;
input n_21;
input n_115;
input n_133;
input n_66;
input n_71;
input n_24;
input n_7;
input n_109;
input n_96;
input n_156;
input n_49;
input n_20;
input n_174;
input n_100;
input n_17;
input n_50;
input n_187;
input n_132;
input n_62;
input n_147;
input n_51;
input n_166;
input n_76;
input n_103;
input n_79;
input n_26;
input n_3;
input n_46;
input n_0;
input n_84;
input n_36;
input n_91;
input n_159;
input n_107;
input n_189;
input n_72;
input n_105;
input n_128;
input n_44;
input n_30;
input n_82;
input n_178;
input n_31;
input n_42;
input n_57;
input n_131;
input n_70;
input n_10;
input n_117;
input n_139;
input n_165;
input n_85;
input n_130;
input n_144;
input n_6;
input n_48;
input n_94;
input n_101;
input n_4;
input n_134;
input n_188;
input n_185;
input n_2;
input n_32;
input n_37;
input n_58;
input n_65;
input n_123;
input n_9;
input n_138;
input n_112;
input n_45;
input n_162;
input n_11;
input n_129;
input n_126;
input n_137;
input n_122;
input n_148;
input n_164;
input n_52;
input n_157;
input n_184;
input n_177;
input n_135;
input n_73;
input n_77;
input n_171;
input n_15;
input n_118;
input n_93;
input n_121;
input n_23;
input n_61;
input n_108;
input n_102;
input n_182;
input n_125;
input n_22;
input n_168;
input n_43;
input n_1;
input n_81;
input n_87;
input n_13;
input n_27;
input n_29;
input n_41;
input n_140;
input n_55;
input n_151;
input n_136;
input n_28;
input n_80;
input n_146;
input n_97;
input n_154;
input n_142;
input n_161;
input n_14;
input n_163;
input n_88;
input n_186;
input n_141;
input n_68;
input n_116;
input n_104;
input n_145;
input n_78;
input n_39;
input n_59;
input n_63;
input n_99;
input n_16;
input n_5;
input n_155;
input n_127;
input n_35;
input n_54;
input n_25;

output n_1236;

wire n_913;
wire n_589;
wire n_1174;
wire n_691;
wire n_423;
wire n_603;
wire n_373;
wire n_1169;
wire n_789;
wire n_850;
wire n_610;
wire n_245;
wire n_319;
wire n_690;
wire n_416;
wire n_1109;
wire n_525;
wire n_817;
wire n_924;
wire n_781;
wire n_717;
wire n_952;
wire n_864;
wire n_1096;
wire n_524;
wire n_1214;
wire n_634;
wire n_1138;
wire n_214;
wire n_764;
wire n_462;
wire n_1196;
wire n_1181;
wire n_410;
wire n_1187;
wire n_1131;
wire n_1225;
wire n_737;
wire n_232;
wire n_568;
wire n_1088;
wire n_766;
wire n_377;
wire n_520;
wire n_870;
wire n_279;
wire n_945;
wire n_958;
wire n_813;
wire n_419;
wire n_270;
wire n_338;
wire n_995;
wire n_285;
wire n_1184;
wire n_202;
wire n_500;
wire n_754;
wire n_665;
wire n_903;
wire n_871;
wire n_1073;
wire n_239;
wire n_402;
wire n_829;
wire n_1062;
wire n_339;
wire n_738;
wire n_672;
wire n_740;
wire n_1018;
wire n_259;
wire n_953;
wire n_1224;
wire n_625;
wire n_557;
wire n_1107;
wire n_989;
wire n_242;
wire n_645;
wire n_331;
wire n_559;
wire n_495;
wire n_267;
wire n_350;
wire n_381;
wire n_795;
wire n_721;
wire n_1084;
wire n_200;
wire n_821;
wire n_561;
wire n_770;
wire n_507;
wire n_486;
wire n_901;
wire n_569;
wire n_1145;
wire n_971;
wire n_787;
wire n_1195;
wire n_518;
wire n_1207;
wire n_222;
wire n_786;
wire n_868;
wire n_884;
wire n_1034;
wire n_1085;
wire n_277;
wire n_432;
wire n_293;
wire n_823;
wire n_620;
wire n_1074;
wire n_859;
wire n_587;
wire n_693;
wire n_863;
wire n_303;
wire n_929;
wire n_206;
wire n_352;
wire n_899;
wire n_611;
wire n_238;
wire n_365;
wire n_1013;
wire n_334;
wire n_192;
wire n_661;
wire n_300;
wire n_533;
wire n_438;
wire n_440;
wire n_273;
wire n_1230;
wire n_612;
wire n_333;
wire n_376;
wire n_512;
wire n_579;
wire n_844;
wire n_1012;
wire n_1213;
wire n_237;
wire n_780;
wire n_1021;
wire n_491;
wire n_1142;
wire n_1140;
wire n_705;
wire n_570;
wire n_260;
wire n_942;
wire n_461;
wire n_1121;
wire n_209;
wire n_490;
wire n_225;
wire n_1006;
wire n_575;
wire n_546;
wire n_503;
wire n_1112;
wire n_700;
wire n_1159;
wire n_772;
wire n_1216;
wire n_676;
wire n_680;
wire n_287;
wire n_302;
wire n_380;
wire n_249;
wire n_1108;
wire n_355;
wire n_212;
wire n_444;
wire n_851;
wire n_257;
wire n_652;
wire n_475;
wire n_947;
wire n_930;
wire n_1179;
wire n_468;
wire n_696;
wire n_482;
wire n_798;
wire n_577;
wire n_407;
wire n_916;
wire n_912;
wire n_460;
wire n_366;
wire n_762;
wire n_555;
wire n_804;
wire n_992;
wire n_966;
wire n_955;
wire n_1182;
wire n_794;
wire n_514;
wire n_418;
wire n_513;
wire n_288;
wire n_1178;
wire n_1026;
wire n_306;
wire n_203;
wire n_436;
wire n_324;
wire n_669;
wire n_931;
wire n_619;
wire n_337;
wire n_437;
wire n_274;
wire n_967;
wire n_1083;
wire n_746;
wire n_292;
wire n_1079;
wire n_615;
wire n_1139;
wire n_517;
wire n_824;
wire n_428;
wire n_892;
wire n_959;
wire n_1101;
wire n_563;
wire n_990;
wire n_867;
wire n_1226;
wire n_944;
wire n_749;
wire n_815;
wire n_542;
wire n_470;
wire n_1087;
wire n_632;
wire n_477;
wire n_650;
wire n_425;
wire n_1155;
wire n_1071;
wire n_712;
wire n_976;
wire n_909;
wire n_767;
wire n_964;
wire n_382;
wire n_489;
wire n_251;
wire n_974;
wire n_506;
wire n_799;
wire n_1147;
wire n_397;
wire n_471;
wire n_351;
wire n_965;
wire n_934;
wire n_1220;
wire n_356;
wire n_698;
wire n_307;
wire n_1209;
wire n_1020;
wire n_646;
wire n_404;
wire n_1058;
wire n_347;
wire n_1042;
wire n_1234;
wire n_479;
wire n_299;
wire n_836;
wire n_564;
wire n_205;
wire n_1029;
wire n_760;
wire n_522;
wire n_367;
wire n_1111;
wire n_970;
wire n_713;
wire n_598;
wire n_345;
wire n_927;
wire n_261;
wire n_1095;
wire n_370;
wire n_706;
wire n_286;
wire n_776;
wire n_424;
wire n_466;
wire n_346;
wire n_348;
wire n_552;
wire n_670;
wire n_379;
wire n_264;
wire n_441;
wire n_1032;
wire n_1217;
wire n_637;
wire n_327;
wire n_1177;
wire n_1231;
wire n_980;
wire n_905;
wire n_207;
wire n_720;
wire n_926;
wire n_194;
wire n_1163;
wire n_1173;
wire n_1068;
wire n_1198;
wire n_487;
wire n_855;
wire n_808;
wire n_553;
wire n_814;
wire n_578;
wire n_405;
wire n_320;
wire n_1134;
wire n_647;
wire n_481;
wire n_600;
wire n_1053;
wire n_529;
wire n_502;
wire n_218;
wire n_247;
wire n_1105;
wire n_547;
wire n_439;
wire n_604;
wire n_677;
wire n_478;
wire n_703;
wire n_1061;
wire n_326;
wire n_681;
wire n_227;
wire n_874;
wire n_707;
wire n_983;
wire n_590;
wire n_699;
wire n_727;
wire n_301;
wire n_545;
wire n_1015;
wire n_1162;
wire n_536;
wire n_325;
wire n_688;
wire n_636;
wire n_427;
wire n_1098;
wire n_442;
wire n_777;
wire n_1080;
wire n_920;
wire n_1086;
wire n_1092;
wire n_986;
wire n_1104;
wire n_729;
wire n_887;
wire n_1122;
wire n_1205;
wire n_1132;
wire n_390;
wire n_1156;
wire n_501;
wire n_314;
wire n_1120;
wire n_1202;
wire n_627;
wire n_1188;
wire n_233;
wire n_957;
wire n_388;
wire n_1218;
wire n_321;
wire n_221;
wire n_861;
wire n_877;
wire n_1119;
wire n_616;
wire n_1055;
wire n_1189;
wire n_1089;
wire n_281;
wire n_262;
wire n_735;
wire n_297;
wire n_1005;
wire n_527;
wire n_845;
wire n_888;
wire n_551;
wire n_417;
wire n_343;
wire n_1222;
wire n_582;
wire n_755;
wire n_1097;
wire n_1219;
wire n_710;
wire n_534;
wire n_278;
wire n_560;
wire n_890;
wire n_842;
wire n_451;
wire n_745;
wire n_742;
wire n_1081;
wire n_769;
wire n_476;
wire n_832;
wire n_535;
wire n_744;
wire n_982;
wire n_915;
wire n_215;
wire n_1075;
wire n_454;
wire n_298;
wire n_1227;
wire n_655;
wire n_403;
wire n_1007;
wire n_657;
wire n_837;
wire n_812;
wire n_606;
wire n_951;
wire n_862;
wire n_659;
wire n_509;
wire n_666;
wire n_430;
wire n_1206;
wire n_722;
wire n_1171;
wire n_1030;
wire n_785;
wire n_999;
wire n_456;
wire n_852;
wire n_704;
wire n_1060;
wire n_1044;
wire n_521;
wire n_873;
wire n_342;
wire n_358;
wire n_608;
wire n_1037;
wire n_317;
wire n_1078;
wire n_266;
wire n_1161;
wire n_811;
wire n_624;
wire n_791;
wire n_876;
wire n_618;
wire n_1191;
wire n_736;
wire n_1025;
wire n_1215;
wire n_241;
wire n_687;
wire n_797;
wire n_480;
wire n_211;
wire n_642;
wire n_408;
wire n_595;
wire n_602;
wire n_592;
wire n_854;
wire n_393;
wire n_474;
wire n_805;
wire n_295;
wire n_1072;
wire n_695;
wire n_730;
wire n_386;
wire n_516;
wire n_1137;
wire n_197;
wire n_640;
wire n_463;
wire n_943;
wire n_1118;
wire n_678;
wire n_651;
wire n_961;
wire n_469;
wire n_1046;
wire n_726;
wire n_1123;
wire n_878;
wire n_771;
wire n_752;
wire n_985;
wire n_421;
wire n_906;
wire n_1180;
wire n_283;
wire n_806;
wire n_649;
wire n_374;
wire n_643;
wire n_226;
wire n_682;
wire n_819;
wire n_586;
wire n_686;
wire n_605;
wire n_1154;
wire n_584;
wire n_1130;
wire n_349;
wire n_756;
wire n_1016;
wire n_1149;
wire n_979;
wire n_897;
wire n_949;
wire n_515;
wire n_807;
wire n_891;
wire n_885;
wire n_198;
wire n_1208;
wire n_396;
wire n_802;
wire n_1151;
wire n_554;
wire n_960;
wire n_714;
wire n_790;
wire n_354;
wire n_725;
wire n_1009;
wire n_230;
wire n_1133;
wire n_883;
wire n_473;
wire n_801;
wire n_818;
wire n_779;
wire n_594;
wire n_1052;
wire n_272;
wire n_833;
wire n_879;
wire n_1117;
wire n_422;
wire n_597;
wire n_1047;
wire n_1050;
wire n_566;
wire n_1201;
wire n_858;
wire n_1185;
wire n_335;
wire n_1035;
wire n_1143;
wire n_344;
wire n_426;
wire n_433;
wire n_398;
wire n_210;
wire n_1090;
wire n_253;
wire n_928;
wire n_1153;
wire n_271;
wire n_465;
wire n_825;
wire n_1103;
wire n_732;
wire n_1192;
wire n_224;
wire n_894;
wire n_420;
wire n_562;
wire n_748;
wire n_510;
wire n_1045;
wire n_256;
wire n_1160;
wire n_1023;
wire n_988;
wire n_330;
wire n_914;
wire n_400;
wire n_689;
wire n_1116;
wire n_282;
wire n_328;
wire n_368;
wire n_467;
wire n_644;
wire n_1197;
wire n_276;
wire n_497;
wire n_1165;
wire n_538;
wire n_576;
wire n_843;
wire n_511;
wire n_455;
wire n_429;
wire n_588;
wire n_638;
wire n_1128;
wire n_1048;
wire n_775;
wire n_667;
wire n_1049;
wire n_869;
wire n_846;
wire n_305;
wire n_312;
wire n_728;
wire n_413;
wire n_715;
wire n_889;
wire n_1066;
wire n_935;
wire n_685;
wire n_911;
wire n_361;
wire n_623;
wire n_1065;
wire n_453;
wire n_810;
wire n_617;
wire n_543;
wire n_236;
wire n_601;
wire n_683;
wire n_565;
wire n_628;
wire n_743;
wire n_1194;
wire n_907;
wire n_660;
wire n_464;
wire n_962;
wire n_941;
wire n_1210;
wire n_847;
wire n_747;
wire n_1135;
wire n_918;
wire n_639;
wire n_452;
wire n_673;
wire n_1038;
wire n_414;
wire n_571;
wire n_284;
wire n_593;
wire n_1164;
wire n_609;
wire n_1193;
wire n_613;
wire n_1022;
wire n_1033;
wire n_409;
wire n_519;
wire n_384;
wire n_1166;
wire n_1056;
wire n_526;
wire n_1040;
wire n_674;
wire n_1158;
wire n_316;
wire n_820;
wire n_872;
wire n_254;
wire n_1157;
wire n_234;
wire n_848;
wire n_280;
wire n_629;
wire n_532;
wire n_763;
wire n_540;
wire n_216;
wire n_692;
wire n_984;
wire n_223;
wire n_750;
wire n_834;
wire n_800;
wire n_395;
wire n_621;
wire n_213;
wire n_1014;
wire n_724;
wire n_493;
wire n_1100;
wire n_585;
wire n_875;
wire n_827;
wire n_697;
wire n_622;
wire n_296;
wire n_880;
wire n_793;
wire n_1175;
wire n_751;
wire n_1027;
wire n_1070;
wire n_739;
wire n_1028;
wire n_1221;
wire n_530;
wire n_792;
wire n_580;
wire n_494;
wire n_434;
wire n_975;
wire n_229;
wire n_394;
wire n_923;
wire n_1124;
wire n_932;
wire n_1183;
wire n_981;
wire n_1110;
wire n_243;
wire n_1204;
wire n_994;
wire n_973;
wire n_268;
wire n_972;
wire n_856;
wire n_1176;
wire n_1054;
wire n_508;
wire n_353;
wire n_1057;
wire n_191;
wire n_978;
wire n_1011;
wire n_828;
wire n_322;
wire n_558;
wire n_653;
wire n_783;
wire n_556;
wire n_1127;
wire n_1008;
wire n_332;
wire n_581;
wire n_294;
wire n_1024;
wire n_830;
wire n_987;
wire n_936;
wire n_541;
wire n_499;
wire n_788;
wire n_908;
wire n_1036;
wire n_341;
wire n_1167;
wire n_549;
wire n_591;
wire n_969;
wire n_919;
wire n_318;
wire n_244;
wire n_679;
wire n_220;
wire n_663;
wire n_443;
wire n_528;
wire n_1200;
wire n_387;
wire n_406;
wire n_826;
wire n_391;
wire n_940;
wire n_1077;
wire n_607;
wire n_956;
wire n_445;
wire n_765;
wire n_385;
wire n_917;
wire n_372;
wire n_631;
wire n_399;
wire n_1170;
wire n_702;
wire n_898;
wire n_857;
wire n_363;
wire n_1067;
wire n_968;
wire n_1235;
wire n_1064;
wire n_633;
wire n_900;
wire n_1093;
wire n_193;
wire n_733;
wire n_761;
wire n_731;
wire n_336;
wire n_315;
wire n_311;
wire n_668;
wire n_758;
wire n_1106;
wire n_648;
wire n_784;
wire n_269;
wire n_816;
wire n_835;
wire n_446;
wire n_1076;
wire n_753;
wire n_701;
wire n_1003;
wire n_1125;
wire n_309;
wire n_401;
wire n_485;
wire n_504;
wire n_483;
wire n_435;
wire n_1141;
wire n_291;
wire n_822;
wire n_1094;
wire n_840;
wire n_1099;
wire n_839;
wire n_759;
wire n_567;
wire n_240;
wire n_369;
wire n_1172;
wire n_614;
wire n_1212;
wire n_831;
wire n_778;
wire n_323;
wire n_550;
wire n_997;
wire n_635;
wire n_694;
wire n_1113;
wire n_248;
wire n_1152;
wire n_921;
wire n_228;
wire n_671;
wire n_1148;
wire n_654;
wire n_488;
wire n_904;
wire n_505;
wire n_498;
wire n_1059;
wire n_684;
wire n_1039;
wire n_539;
wire n_1150;
wire n_977;
wire n_449;
wire n_392;
wire n_459;
wire n_1136;
wire n_458;
wire n_1190;
wire n_1144;
wire n_383;
wire n_838;
wire n_950;
wire n_1017;
wire n_711;
wire n_734;
wire n_723;
wire n_658;
wire n_630;
wire n_362;
wire n_310;
wire n_709;
wire n_809;
wire n_235;
wire n_881;
wire n_1019;
wire n_662;
wire n_641;
wire n_910;
wire n_290;
wire n_741;
wire n_939;
wire n_371;
wire n_199;
wire n_217;
wire n_1114;
wire n_708;
wire n_308;
wire n_1223;
wire n_201;
wire n_572;
wire n_1199;
wire n_865;
wire n_1041;
wire n_993;
wire n_948;
wire n_922;
wire n_1004;
wire n_448;
wire n_860;
wire n_1043;
wire n_255;
wire n_450;
wire n_896;
wire n_902;
wire n_1031;
wire n_853;
wire n_716;
wire n_196;
wire n_774;
wire n_933;
wire n_596;
wire n_954;
wire n_1168;
wire n_219;
wire n_231;
wire n_656;
wire n_492;
wire n_574;
wire n_252;
wire n_664;
wire n_1229;
wire n_415;
wire n_544;
wire n_1186;
wire n_599;
wire n_768;
wire n_1091;
wire n_537;
wire n_1063;
wire n_991;
wire n_389;
wire n_1126;
wire n_195;
wire n_938;
wire n_895;
wire n_304;
wire n_583;
wire n_1000;
wire n_313;
wire n_626;
wire n_378;
wire n_946;
wire n_757;
wire n_375;
wire n_1146;
wire n_1203;
wire n_998;
wire n_472;
wire n_937;
wire n_265;
wire n_208;
wire n_275;
wire n_204;
wire n_1232;
wire n_996;
wire n_1211;
wire n_963;
wire n_1082;
wire n_496;
wire n_866;
wire n_246;
wire n_925;
wire n_1001;
wire n_1115;
wire n_1002;
wire n_1051;
wire n_719;
wire n_263;
wire n_1102;
wire n_360;
wire n_1129;
wire n_250;
wire n_773;
wire n_1010;
wire n_882;
wire n_803;
wire n_329;
wire n_718;
wire n_340;
wire n_289;
wire n_548;
wire n_523;
wire n_457;
wire n_782;
wire n_364;
wire n_258;
wire n_431;
wire n_1228;
wire n_411;
wire n_484;
wire n_849;
wire n_357;
wire n_412;
wire n_447;
wire n_1233;
wire n_893;
wire n_841;
wire n_886;
wire n_1069;
wire n_359;
wire n_573;
wire n_796;
wire n_531;
wire n_675;

CKINVDCx5p33_ASAP7_75t_R g191 ( 
.A(n_53),
.Y(n_191)
);

CKINVDCx5p33_ASAP7_75t_R g192 ( 
.A(n_23),
.Y(n_192)
);

INVx2_ASAP7_75t_L g193 ( 
.A(n_3),
.Y(n_193)
);

CKINVDCx5p33_ASAP7_75t_R g194 ( 
.A(n_143),
.Y(n_194)
);

CKINVDCx5p33_ASAP7_75t_R g195 ( 
.A(n_134),
.Y(n_195)
);

CKINVDCx5p33_ASAP7_75t_R g196 ( 
.A(n_35),
.Y(n_196)
);

CKINVDCx5p33_ASAP7_75t_R g197 ( 
.A(n_91),
.Y(n_197)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_76),
.Y(n_198)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_162),
.Y(n_199)
);

CKINVDCx5p33_ASAP7_75t_R g200 ( 
.A(n_151),
.Y(n_200)
);

INVx1_ASAP7_75t_SL g201 ( 
.A(n_144),
.Y(n_201)
);

INVx2_ASAP7_75t_L g202 ( 
.A(n_139),
.Y(n_202)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_65),
.Y(n_203)
);

CKINVDCx5p33_ASAP7_75t_R g204 ( 
.A(n_10),
.Y(n_204)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_138),
.Y(n_205)
);

CKINVDCx5p33_ASAP7_75t_R g206 ( 
.A(n_104),
.Y(n_206)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_43),
.Y(n_207)
);

BUFx6f_ASAP7_75t_L g208 ( 
.A(n_93),
.Y(n_208)
);

CKINVDCx5p33_ASAP7_75t_R g209 ( 
.A(n_92),
.Y(n_209)
);

CKINVDCx5p33_ASAP7_75t_R g210 ( 
.A(n_18),
.Y(n_210)
);

CKINVDCx5p33_ASAP7_75t_R g211 ( 
.A(n_176),
.Y(n_211)
);

CKINVDCx5p33_ASAP7_75t_R g212 ( 
.A(n_58),
.Y(n_212)
);

CKINVDCx5p33_ASAP7_75t_R g213 ( 
.A(n_52),
.Y(n_213)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_98),
.Y(n_214)
);

BUFx6f_ASAP7_75t_L g215 ( 
.A(n_21),
.Y(n_215)
);

CKINVDCx5p33_ASAP7_75t_R g216 ( 
.A(n_13),
.Y(n_216)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_28),
.Y(n_217)
);

CKINVDCx5p33_ASAP7_75t_R g218 ( 
.A(n_186),
.Y(n_218)
);

CKINVDCx5p33_ASAP7_75t_R g219 ( 
.A(n_102),
.Y(n_219)
);

CKINVDCx5p33_ASAP7_75t_R g220 ( 
.A(n_95),
.Y(n_220)
);

CKINVDCx5p33_ASAP7_75t_R g221 ( 
.A(n_187),
.Y(n_221)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_15),
.Y(n_222)
);

CKINVDCx5p33_ASAP7_75t_R g223 ( 
.A(n_114),
.Y(n_223)
);

CKINVDCx5p33_ASAP7_75t_R g224 ( 
.A(n_167),
.Y(n_224)
);

CKINVDCx5p33_ASAP7_75t_R g225 ( 
.A(n_137),
.Y(n_225)
);

CKINVDCx5p33_ASAP7_75t_R g226 ( 
.A(n_7),
.Y(n_226)
);

CKINVDCx5p33_ASAP7_75t_R g227 ( 
.A(n_63),
.Y(n_227)
);

CKINVDCx5p33_ASAP7_75t_R g228 ( 
.A(n_41),
.Y(n_228)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_133),
.Y(n_229)
);

CKINVDCx5p33_ASAP7_75t_R g230 ( 
.A(n_41),
.Y(n_230)
);

CKINVDCx5p33_ASAP7_75t_R g231 ( 
.A(n_40),
.Y(n_231)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_171),
.Y(n_232)
);

HB1xp67_ASAP7_75t_L g233 ( 
.A(n_19),
.Y(n_233)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_136),
.Y(n_234)
);

CKINVDCx5p33_ASAP7_75t_R g235 ( 
.A(n_2),
.Y(n_235)
);

CKINVDCx20_ASAP7_75t_R g236 ( 
.A(n_154),
.Y(n_236)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_86),
.Y(n_237)
);

CKINVDCx20_ASAP7_75t_R g238 ( 
.A(n_182),
.Y(n_238)
);

CKINVDCx5p33_ASAP7_75t_R g239 ( 
.A(n_189),
.Y(n_239)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_163),
.Y(n_240)
);

CKINVDCx5p33_ASAP7_75t_R g241 ( 
.A(n_24),
.Y(n_241)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_72),
.Y(n_242)
);

CKINVDCx5p33_ASAP7_75t_R g243 ( 
.A(n_135),
.Y(n_243)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_12),
.Y(n_244)
);

CKINVDCx5p33_ASAP7_75t_R g245 ( 
.A(n_108),
.Y(n_245)
);

BUFx6f_ASAP7_75t_L g246 ( 
.A(n_19),
.Y(n_246)
);

CKINVDCx5p33_ASAP7_75t_R g247 ( 
.A(n_168),
.Y(n_247)
);

CKINVDCx5p33_ASAP7_75t_R g248 ( 
.A(n_60),
.Y(n_248)
);

CKINVDCx5p33_ASAP7_75t_R g249 ( 
.A(n_8),
.Y(n_249)
);

CKINVDCx5p33_ASAP7_75t_R g250 ( 
.A(n_57),
.Y(n_250)
);

CKINVDCx5p33_ASAP7_75t_R g251 ( 
.A(n_158),
.Y(n_251)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_10),
.Y(n_252)
);

CKINVDCx5p33_ASAP7_75t_R g253 ( 
.A(n_142),
.Y(n_253)
);

BUFx3_ASAP7_75t_L g254 ( 
.A(n_97),
.Y(n_254)
);

CKINVDCx5p33_ASAP7_75t_R g255 ( 
.A(n_69),
.Y(n_255)
);

CKINVDCx5p33_ASAP7_75t_R g256 ( 
.A(n_120),
.Y(n_256)
);

CKINVDCx5p33_ASAP7_75t_R g257 ( 
.A(n_46),
.Y(n_257)
);

CKINVDCx5p33_ASAP7_75t_R g258 ( 
.A(n_31),
.Y(n_258)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_66),
.Y(n_259)
);

CKINVDCx5p33_ASAP7_75t_R g260 ( 
.A(n_126),
.Y(n_260)
);

CKINVDCx5p33_ASAP7_75t_R g261 ( 
.A(n_90),
.Y(n_261)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_83),
.Y(n_262)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_15),
.Y(n_263)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_166),
.Y(n_264)
);

CKINVDCx5p33_ASAP7_75t_R g265 ( 
.A(n_116),
.Y(n_265)
);

CKINVDCx5p33_ASAP7_75t_R g266 ( 
.A(n_70),
.Y(n_266)
);

CKINVDCx5p33_ASAP7_75t_R g267 ( 
.A(n_152),
.Y(n_267)
);

CKINVDCx20_ASAP7_75t_R g268 ( 
.A(n_125),
.Y(n_268)
);

CKINVDCx5p33_ASAP7_75t_R g269 ( 
.A(n_147),
.Y(n_269)
);

BUFx3_ASAP7_75t_L g270 ( 
.A(n_161),
.Y(n_270)
);

CKINVDCx5p33_ASAP7_75t_R g271 ( 
.A(n_145),
.Y(n_271)
);

CKINVDCx5p33_ASAP7_75t_R g272 ( 
.A(n_94),
.Y(n_272)
);

CKINVDCx5p33_ASAP7_75t_R g273 ( 
.A(n_122),
.Y(n_273)
);

CKINVDCx5p33_ASAP7_75t_R g274 ( 
.A(n_115),
.Y(n_274)
);

BUFx3_ASAP7_75t_L g275 ( 
.A(n_42),
.Y(n_275)
);

CKINVDCx5p33_ASAP7_75t_R g276 ( 
.A(n_16),
.Y(n_276)
);

INVx1_ASAP7_75t_SL g277 ( 
.A(n_61),
.Y(n_277)
);

CKINVDCx5p33_ASAP7_75t_R g278 ( 
.A(n_112),
.Y(n_278)
);

BUFx2_ASAP7_75t_SL g279 ( 
.A(n_164),
.Y(n_279)
);

CKINVDCx5p33_ASAP7_75t_R g280 ( 
.A(n_26),
.Y(n_280)
);

CKINVDCx20_ASAP7_75t_R g281 ( 
.A(n_88),
.Y(n_281)
);

CKINVDCx5p33_ASAP7_75t_R g282 ( 
.A(n_7),
.Y(n_282)
);

CKINVDCx5p33_ASAP7_75t_R g283 ( 
.A(n_188),
.Y(n_283)
);

CKINVDCx20_ASAP7_75t_R g284 ( 
.A(n_33),
.Y(n_284)
);

CKINVDCx5p33_ASAP7_75t_R g285 ( 
.A(n_107),
.Y(n_285)
);

HB1xp67_ASAP7_75t_L g286 ( 
.A(n_87),
.Y(n_286)
);

CKINVDCx5p33_ASAP7_75t_R g287 ( 
.A(n_6),
.Y(n_287)
);

CKINVDCx5p33_ASAP7_75t_R g288 ( 
.A(n_146),
.Y(n_288)
);

CKINVDCx5p33_ASAP7_75t_R g289 ( 
.A(n_2),
.Y(n_289)
);

CKINVDCx5p33_ASAP7_75t_R g290 ( 
.A(n_160),
.Y(n_290)
);

CKINVDCx5p33_ASAP7_75t_R g291 ( 
.A(n_1),
.Y(n_291)
);

BUFx10_ASAP7_75t_L g292 ( 
.A(n_89),
.Y(n_292)
);

BUFx3_ASAP7_75t_L g293 ( 
.A(n_23),
.Y(n_293)
);

CKINVDCx5p33_ASAP7_75t_R g294 ( 
.A(n_178),
.Y(n_294)
);

CKINVDCx5p33_ASAP7_75t_R g295 ( 
.A(n_54),
.Y(n_295)
);

CKINVDCx5p33_ASAP7_75t_R g296 ( 
.A(n_11),
.Y(n_296)
);

CKINVDCx5p33_ASAP7_75t_R g297 ( 
.A(n_140),
.Y(n_297)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_29),
.Y(n_298)
);

CKINVDCx5p33_ASAP7_75t_R g299 ( 
.A(n_49),
.Y(n_299)
);

CKINVDCx5p33_ASAP7_75t_R g300 ( 
.A(n_99),
.Y(n_300)
);

CKINVDCx20_ASAP7_75t_R g301 ( 
.A(n_17),
.Y(n_301)
);

CKINVDCx5p33_ASAP7_75t_R g302 ( 
.A(n_109),
.Y(n_302)
);

CKINVDCx14_ASAP7_75t_R g303 ( 
.A(n_28),
.Y(n_303)
);

CKINVDCx5p33_ASAP7_75t_R g304 ( 
.A(n_111),
.Y(n_304)
);

CKINVDCx5p33_ASAP7_75t_R g305 ( 
.A(n_96),
.Y(n_305)
);

CKINVDCx5p33_ASAP7_75t_R g306 ( 
.A(n_25),
.Y(n_306)
);

CKINVDCx5p33_ASAP7_75t_R g307 ( 
.A(n_80),
.Y(n_307)
);

CKINVDCx5p33_ASAP7_75t_R g308 ( 
.A(n_4),
.Y(n_308)
);

CKINVDCx5p33_ASAP7_75t_R g309 ( 
.A(n_64),
.Y(n_309)
);

INVx1_ASAP7_75t_SL g310 ( 
.A(n_30),
.Y(n_310)
);

CKINVDCx5p33_ASAP7_75t_R g311 ( 
.A(n_169),
.Y(n_311)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_293),
.Y(n_312)
);

CKINVDCx5p33_ASAP7_75t_R g313 ( 
.A(n_303),
.Y(n_313)
);

CKINVDCx20_ASAP7_75t_R g314 ( 
.A(n_236),
.Y(n_314)
);

CKINVDCx20_ASAP7_75t_R g315 ( 
.A(n_238),
.Y(n_315)
);

CKINVDCx5p33_ASAP7_75t_R g316 ( 
.A(n_292),
.Y(n_316)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_293),
.Y(n_317)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_217),
.Y(n_318)
);

CKINVDCx16_ASAP7_75t_R g319 ( 
.A(n_292),
.Y(n_319)
);

CKINVDCx5p33_ASAP7_75t_R g320 ( 
.A(n_292),
.Y(n_320)
);

CKINVDCx5p33_ASAP7_75t_R g321 ( 
.A(n_191),
.Y(n_321)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_222),
.Y(n_322)
);

CKINVDCx5p33_ASAP7_75t_R g323 ( 
.A(n_191),
.Y(n_323)
);

HB1xp67_ASAP7_75t_L g324 ( 
.A(n_233),
.Y(n_324)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_244),
.Y(n_325)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_252),
.Y(n_326)
);

CKINVDCx5p33_ASAP7_75t_R g327 ( 
.A(n_194),
.Y(n_327)
);

NOR2xp33_ASAP7_75t_L g328 ( 
.A(n_286),
.B(n_198),
.Y(n_328)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_263),
.Y(n_329)
);

CKINVDCx20_ASAP7_75t_R g330 ( 
.A(n_268),
.Y(n_330)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_298),
.Y(n_331)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_193),
.Y(n_332)
);

CKINVDCx20_ASAP7_75t_R g333 ( 
.A(n_281),
.Y(n_333)
);

HB1xp67_ASAP7_75t_L g334 ( 
.A(n_192),
.Y(n_334)
);

BUFx3_ASAP7_75t_L g335 ( 
.A(n_254),
.Y(n_335)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_193),
.Y(n_336)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_215),
.Y(n_337)
);

CKINVDCx5p33_ASAP7_75t_R g338 ( 
.A(n_194),
.Y(n_338)
);

NOR2xp67_ASAP7_75t_L g339 ( 
.A(n_192),
.B(n_0),
.Y(n_339)
);

INVx2_ASAP7_75t_L g340 ( 
.A(n_215),
.Y(n_340)
);

CKINVDCx20_ASAP7_75t_R g341 ( 
.A(n_284),
.Y(n_341)
);

INVx1_ASAP7_75t_L g342 ( 
.A(n_215),
.Y(n_342)
);

INVxp67_ASAP7_75t_SL g343 ( 
.A(n_215),
.Y(n_343)
);

NOR2xp67_ASAP7_75t_L g344 ( 
.A(n_196),
.B(n_0),
.Y(n_344)
);

INVxp67_ASAP7_75t_SL g345 ( 
.A(n_215),
.Y(n_345)
);

CKINVDCx20_ASAP7_75t_R g346 ( 
.A(n_301),
.Y(n_346)
);

INVx1_ASAP7_75t_L g347 ( 
.A(n_246),
.Y(n_347)
);

INVx1_ASAP7_75t_L g348 ( 
.A(n_246),
.Y(n_348)
);

INVx1_ASAP7_75t_L g349 ( 
.A(n_246),
.Y(n_349)
);

HB1xp67_ASAP7_75t_L g350 ( 
.A(n_196),
.Y(n_350)
);

CKINVDCx20_ASAP7_75t_R g351 ( 
.A(n_254),
.Y(n_351)
);

INVx1_ASAP7_75t_L g352 ( 
.A(n_246),
.Y(n_352)
);

CKINVDCx5p33_ASAP7_75t_R g353 ( 
.A(n_195),
.Y(n_353)
);

CKINVDCx5p33_ASAP7_75t_R g354 ( 
.A(n_195),
.Y(n_354)
);

HB1xp67_ASAP7_75t_L g355 ( 
.A(n_306),
.Y(n_355)
);

CKINVDCx5p33_ASAP7_75t_R g356 ( 
.A(n_197),
.Y(n_356)
);

NOR2xp33_ASAP7_75t_L g357 ( 
.A(n_199),
.B(n_1),
.Y(n_357)
);

INVx1_ASAP7_75t_L g358 ( 
.A(n_246),
.Y(n_358)
);

INVx1_ASAP7_75t_L g359 ( 
.A(n_203),
.Y(n_359)
);

CKINVDCx5p33_ASAP7_75t_R g360 ( 
.A(n_197),
.Y(n_360)
);

CKINVDCx5p33_ASAP7_75t_R g361 ( 
.A(n_200),
.Y(n_361)
);

INVxp67_ASAP7_75t_SL g362 ( 
.A(n_270),
.Y(n_362)
);

CKINVDCx5p33_ASAP7_75t_R g363 ( 
.A(n_200),
.Y(n_363)
);

INVx2_ASAP7_75t_L g364 ( 
.A(n_270),
.Y(n_364)
);

BUFx3_ASAP7_75t_L g365 ( 
.A(n_275),
.Y(n_365)
);

CKINVDCx5p33_ASAP7_75t_R g366 ( 
.A(n_305),
.Y(n_366)
);

INVx1_ASAP7_75t_L g367 ( 
.A(n_205),
.Y(n_367)
);

INVx1_ASAP7_75t_L g368 ( 
.A(n_207),
.Y(n_368)
);

CKINVDCx20_ASAP7_75t_R g369 ( 
.A(n_275),
.Y(n_369)
);

NOR2xp67_ASAP7_75t_L g370 ( 
.A(n_306),
.B(n_3),
.Y(n_370)
);

CKINVDCx20_ASAP7_75t_R g371 ( 
.A(n_308),
.Y(n_371)
);

CKINVDCx5p33_ASAP7_75t_R g372 ( 
.A(n_305),
.Y(n_372)
);

INVxp67_ASAP7_75t_L g373 ( 
.A(n_308),
.Y(n_373)
);

INVx1_ASAP7_75t_L g374 ( 
.A(n_214),
.Y(n_374)
);

INVx1_ASAP7_75t_L g375 ( 
.A(n_229),
.Y(n_375)
);

INVx1_ASAP7_75t_L g376 ( 
.A(n_232),
.Y(n_376)
);

INVx1_ASAP7_75t_L g377 ( 
.A(n_234),
.Y(n_377)
);

CKINVDCx5p33_ASAP7_75t_R g378 ( 
.A(n_307),
.Y(n_378)
);

CKINVDCx5p33_ASAP7_75t_R g379 ( 
.A(n_307),
.Y(n_379)
);

INVx1_ASAP7_75t_L g380 ( 
.A(n_237),
.Y(n_380)
);

NAND2xp5_ASAP7_75t_L g381 ( 
.A(n_240),
.B(n_4),
.Y(n_381)
);

NOR2xp33_ASAP7_75t_L g382 ( 
.A(n_242),
.B(n_5),
.Y(n_382)
);

INVx1_ASAP7_75t_L g383 ( 
.A(n_259),
.Y(n_383)
);

CKINVDCx5p33_ASAP7_75t_R g384 ( 
.A(n_309),
.Y(n_384)
);

CKINVDCx5p33_ASAP7_75t_R g385 ( 
.A(n_309),
.Y(n_385)
);

CKINVDCx5p33_ASAP7_75t_R g386 ( 
.A(n_311),
.Y(n_386)
);

INVxp67_ASAP7_75t_L g387 ( 
.A(n_204),
.Y(n_387)
);

CKINVDCx20_ASAP7_75t_R g388 ( 
.A(n_210),
.Y(n_388)
);

INVx1_ASAP7_75t_L g389 ( 
.A(n_262),
.Y(n_389)
);

CKINVDCx5p33_ASAP7_75t_R g390 ( 
.A(n_311),
.Y(n_390)
);

CKINVDCx5p33_ASAP7_75t_R g391 ( 
.A(n_216),
.Y(n_391)
);

CKINVDCx20_ASAP7_75t_R g392 ( 
.A(n_226),
.Y(n_392)
);

INVx1_ASAP7_75t_L g393 ( 
.A(n_264),
.Y(n_393)
);

CKINVDCx11_ASAP7_75t_R g394 ( 
.A(n_310),
.Y(n_394)
);

INVxp67_ASAP7_75t_L g395 ( 
.A(n_228),
.Y(n_395)
);

INVx1_ASAP7_75t_L g396 ( 
.A(n_230),
.Y(n_396)
);

CKINVDCx5p33_ASAP7_75t_R g397 ( 
.A(n_231),
.Y(n_397)
);

NAND2xp5_ASAP7_75t_L g398 ( 
.A(n_202),
.B(n_5),
.Y(n_398)
);

INVxp67_ASAP7_75t_SL g399 ( 
.A(n_202),
.Y(n_399)
);

CKINVDCx5p33_ASAP7_75t_R g400 ( 
.A(n_235),
.Y(n_400)
);

AND2x2_ASAP7_75t_L g401 ( 
.A(n_241),
.B(n_6),
.Y(n_401)
);

INVxp67_ASAP7_75t_SL g402 ( 
.A(n_208),
.Y(n_402)
);

CKINVDCx5p33_ASAP7_75t_R g403 ( 
.A(n_394),
.Y(n_403)
);

NOR2xp33_ASAP7_75t_R g404 ( 
.A(n_321),
.B(n_206),
.Y(n_404)
);

CKINVDCx20_ASAP7_75t_R g405 ( 
.A(n_341),
.Y(n_405)
);

BUFx6f_ASAP7_75t_L g406 ( 
.A(n_340),
.Y(n_406)
);

INVx1_ASAP7_75t_L g407 ( 
.A(n_343),
.Y(n_407)
);

INVx3_ASAP7_75t_L g408 ( 
.A(n_340),
.Y(n_408)
);

INVx1_ASAP7_75t_L g409 ( 
.A(n_345),
.Y(n_409)
);

INVx2_ASAP7_75t_L g410 ( 
.A(n_337),
.Y(n_410)
);

INVx1_ASAP7_75t_L g411 ( 
.A(n_318),
.Y(n_411)
);

CKINVDCx20_ASAP7_75t_R g412 ( 
.A(n_346),
.Y(n_412)
);

CKINVDCx5p33_ASAP7_75t_R g413 ( 
.A(n_314),
.Y(n_413)
);

CKINVDCx5p33_ASAP7_75t_R g414 ( 
.A(n_315),
.Y(n_414)
);

INVx1_ASAP7_75t_L g415 ( 
.A(n_322),
.Y(n_415)
);

INVx1_ASAP7_75t_L g416 ( 
.A(n_325),
.Y(n_416)
);

INVx1_ASAP7_75t_L g417 ( 
.A(n_326),
.Y(n_417)
);

AND2x4_ASAP7_75t_L g418 ( 
.A(n_362),
.B(n_201),
.Y(n_418)
);

CKINVDCx5p33_ASAP7_75t_R g419 ( 
.A(n_330),
.Y(n_419)
);

NOR2xp67_ASAP7_75t_L g420 ( 
.A(n_316),
.B(n_209),
.Y(n_420)
);

INVx2_ASAP7_75t_L g421 ( 
.A(n_342),
.Y(n_421)
);

CKINVDCx20_ASAP7_75t_R g422 ( 
.A(n_333),
.Y(n_422)
);

CKINVDCx20_ASAP7_75t_R g423 ( 
.A(n_371),
.Y(n_423)
);

INVx1_ASAP7_75t_L g424 ( 
.A(n_329),
.Y(n_424)
);

INVx2_ASAP7_75t_L g425 ( 
.A(n_347),
.Y(n_425)
);

INVx1_ASAP7_75t_L g426 ( 
.A(n_331),
.Y(n_426)
);

INVx1_ASAP7_75t_L g427 ( 
.A(n_312),
.Y(n_427)
);

AND2x6_ASAP7_75t_L g428 ( 
.A(n_335),
.B(n_208),
.Y(n_428)
);

INVx3_ASAP7_75t_L g429 ( 
.A(n_348),
.Y(n_429)
);

BUFx6f_ASAP7_75t_L g430 ( 
.A(n_349),
.Y(n_430)
);

HB1xp67_ASAP7_75t_L g431 ( 
.A(n_391),
.Y(n_431)
);

AOI22xp5_ASAP7_75t_L g432 ( 
.A1(n_316),
.A2(n_249),
.B1(n_258),
.B2(n_276),
.Y(n_432)
);

BUFx6f_ASAP7_75t_L g433 ( 
.A(n_352),
.Y(n_433)
);

INVx1_ASAP7_75t_L g434 ( 
.A(n_317),
.Y(n_434)
);

INVx2_ASAP7_75t_L g435 ( 
.A(n_358),
.Y(n_435)
);

INVx3_ASAP7_75t_L g436 ( 
.A(n_364),
.Y(n_436)
);

INVx1_ASAP7_75t_L g437 ( 
.A(n_364),
.Y(n_437)
);

HB1xp67_ASAP7_75t_L g438 ( 
.A(n_391),
.Y(n_438)
);

INVx2_ASAP7_75t_L g439 ( 
.A(n_332),
.Y(n_439)
);

INVx1_ASAP7_75t_L g440 ( 
.A(n_402),
.Y(n_440)
);

CKINVDCx5p33_ASAP7_75t_R g441 ( 
.A(n_321),
.Y(n_441)
);

CKINVDCx5p33_ASAP7_75t_R g442 ( 
.A(n_323),
.Y(n_442)
);

INVx2_ASAP7_75t_L g443 ( 
.A(n_336),
.Y(n_443)
);

INVx1_ASAP7_75t_L g444 ( 
.A(n_359),
.Y(n_444)
);

INVx3_ASAP7_75t_L g445 ( 
.A(n_335),
.Y(n_445)
);

INVx1_ASAP7_75t_L g446 ( 
.A(n_367),
.Y(n_446)
);

HB1xp67_ASAP7_75t_L g447 ( 
.A(n_397),
.Y(n_447)
);

INVx1_ASAP7_75t_L g448 ( 
.A(n_368),
.Y(n_448)
);

INVx1_ASAP7_75t_L g449 ( 
.A(n_374),
.Y(n_449)
);

NAND2xp5_ASAP7_75t_L g450 ( 
.A(n_365),
.B(n_277),
.Y(n_450)
);

CKINVDCx5p33_ASAP7_75t_R g451 ( 
.A(n_323),
.Y(n_451)
);

INVx1_ASAP7_75t_L g452 ( 
.A(n_375),
.Y(n_452)
);

CKINVDCx5p33_ASAP7_75t_R g453 ( 
.A(n_327),
.Y(n_453)
);

CKINVDCx5p33_ASAP7_75t_R g454 ( 
.A(n_327),
.Y(n_454)
);

INVx2_ASAP7_75t_L g455 ( 
.A(n_376),
.Y(n_455)
);

NAND2xp5_ASAP7_75t_L g456 ( 
.A(n_365),
.B(n_211),
.Y(n_456)
);

CKINVDCx5p33_ASAP7_75t_R g457 ( 
.A(n_338),
.Y(n_457)
);

INVx1_ASAP7_75t_L g458 ( 
.A(n_377),
.Y(n_458)
);

CKINVDCx5p33_ASAP7_75t_R g459 ( 
.A(n_338),
.Y(n_459)
);

BUFx2_ASAP7_75t_L g460 ( 
.A(n_388),
.Y(n_460)
);

INVxp67_ASAP7_75t_L g461 ( 
.A(n_334),
.Y(n_461)
);

INVx3_ASAP7_75t_L g462 ( 
.A(n_380),
.Y(n_462)
);

INVx2_ASAP7_75t_L g463 ( 
.A(n_383),
.Y(n_463)
);

NAND2xp5_ASAP7_75t_L g464 ( 
.A(n_396),
.B(n_212),
.Y(n_464)
);

AND2x4_ASAP7_75t_L g465 ( 
.A(n_399),
.B(n_208),
.Y(n_465)
);

NAND2xp5_ASAP7_75t_L g466 ( 
.A(n_328),
.B(n_213),
.Y(n_466)
);

INVx3_ASAP7_75t_L g467 ( 
.A(n_389),
.Y(n_467)
);

AND2x6_ASAP7_75t_L g468 ( 
.A(n_393),
.B(n_208),
.Y(n_468)
);

CKINVDCx5p33_ASAP7_75t_R g469 ( 
.A(n_353),
.Y(n_469)
);

BUFx10_ASAP7_75t_L g470 ( 
.A(n_353),
.Y(n_470)
);

NAND2xp33_ASAP7_75t_SL g471 ( 
.A(n_313),
.B(n_280),
.Y(n_471)
);

INVx1_ASAP7_75t_L g472 ( 
.A(n_381),
.Y(n_472)
);

AND2x6_ASAP7_75t_L g473 ( 
.A(n_472),
.B(n_401),
.Y(n_473)
);

BUFx4f_ASAP7_75t_L g474 ( 
.A(n_418),
.Y(n_474)
);

NAND2xp5_ASAP7_75t_L g475 ( 
.A(n_445),
.B(n_320),
.Y(n_475)
);

NAND2xp5_ASAP7_75t_L g476 ( 
.A(n_445),
.B(n_320),
.Y(n_476)
);

NAND2xp5_ASAP7_75t_L g477 ( 
.A(n_445),
.B(n_319),
.Y(n_477)
);

NAND2xp5_ASAP7_75t_L g478 ( 
.A(n_418),
.B(n_354),
.Y(n_478)
);

INVx1_ASAP7_75t_L g479 ( 
.A(n_427),
.Y(n_479)
);

AND2x2_ASAP7_75t_SL g480 ( 
.A(n_418),
.B(n_401),
.Y(n_480)
);

INVx2_ASAP7_75t_L g481 ( 
.A(n_429),
.Y(n_481)
);

BUFx10_ASAP7_75t_L g482 ( 
.A(n_441),
.Y(n_482)
);

INVx1_ASAP7_75t_L g483 ( 
.A(n_434),
.Y(n_483)
);

NOR2xp33_ASAP7_75t_L g484 ( 
.A(n_464),
.B(n_354),
.Y(n_484)
);

AND2x2_ASAP7_75t_L g485 ( 
.A(n_461),
.B(n_313),
.Y(n_485)
);

NOR2xp33_ASAP7_75t_L g486 ( 
.A(n_466),
.B(n_356),
.Y(n_486)
);

NAND2xp5_ASAP7_75t_SL g487 ( 
.A(n_404),
.B(n_356),
.Y(n_487)
);

INVx1_ASAP7_75t_L g488 ( 
.A(n_437),
.Y(n_488)
);

NAND2xp33_ASAP7_75t_SL g489 ( 
.A(n_441),
.B(n_398),
.Y(n_489)
);

NOR2xp33_ASAP7_75t_SL g490 ( 
.A(n_403),
.B(n_392),
.Y(n_490)
);

INVx2_ASAP7_75t_L g491 ( 
.A(n_429),
.Y(n_491)
);

INVx2_ASAP7_75t_SL g492 ( 
.A(n_470),
.Y(n_492)
);

CKINVDCx5p33_ASAP7_75t_R g493 ( 
.A(n_413),
.Y(n_493)
);

BUFx2_ASAP7_75t_L g494 ( 
.A(n_442),
.Y(n_494)
);

NOR2xp33_ASAP7_75t_L g495 ( 
.A(n_440),
.B(n_360),
.Y(n_495)
);

INVx4_ASAP7_75t_L g496 ( 
.A(n_465),
.Y(n_496)
);

INVx5_ASAP7_75t_L g497 ( 
.A(n_428),
.Y(n_497)
);

INVx1_ASAP7_75t_L g498 ( 
.A(n_411),
.Y(n_498)
);

INVx6_ASAP7_75t_L g499 ( 
.A(n_465),
.Y(n_499)
);

INVx1_ASAP7_75t_L g500 ( 
.A(n_415),
.Y(n_500)
);

INVx2_ASAP7_75t_L g501 ( 
.A(n_429),
.Y(n_501)
);

INVx1_ASAP7_75t_L g502 ( 
.A(n_416),
.Y(n_502)
);

AND2x4_ASAP7_75t_L g503 ( 
.A(n_462),
.B(n_351),
.Y(n_503)
);

INVx1_ASAP7_75t_L g504 ( 
.A(n_417),
.Y(n_504)
);

NOR2xp33_ASAP7_75t_L g505 ( 
.A(n_407),
.B(n_360),
.Y(n_505)
);

AND2x2_ASAP7_75t_L g506 ( 
.A(n_470),
.B(n_397),
.Y(n_506)
);

BUFx6f_ASAP7_75t_L g507 ( 
.A(n_406),
.Y(n_507)
);

AND2x2_ASAP7_75t_L g508 ( 
.A(n_470),
.B(n_400),
.Y(n_508)
);

INVx1_ASAP7_75t_L g509 ( 
.A(n_424),
.Y(n_509)
);

OR2x2_ASAP7_75t_L g510 ( 
.A(n_460),
.B(n_350),
.Y(n_510)
);

NOR2xp33_ASAP7_75t_L g511 ( 
.A(n_409),
.B(n_456),
.Y(n_511)
);

OR2x6_ASAP7_75t_L g512 ( 
.A(n_431),
.B(n_324),
.Y(n_512)
);

INVx4_ASAP7_75t_SL g513 ( 
.A(n_428),
.Y(n_513)
);

NOR2xp33_ASAP7_75t_L g514 ( 
.A(n_450),
.B(n_361),
.Y(n_514)
);

INVx1_ASAP7_75t_L g515 ( 
.A(n_426),
.Y(n_515)
);

INVx3_ASAP7_75t_L g516 ( 
.A(n_436),
.Y(n_516)
);

INVx1_ASAP7_75t_L g517 ( 
.A(n_455),
.Y(n_517)
);

INVx2_ASAP7_75t_L g518 ( 
.A(n_410),
.Y(n_518)
);

BUFx10_ASAP7_75t_L g519 ( 
.A(n_442),
.Y(n_519)
);

INVx1_ASAP7_75t_L g520 ( 
.A(n_455),
.Y(n_520)
);

INVx1_ASAP7_75t_SL g521 ( 
.A(n_405),
.Y(n_521)
);

INVx4_ASAP7_75t_L g522 ( 
.A(n_465),
.Y(n_522)
);

NAND2xp5_ASAP7_75t_L g523 ( 
.A(n_462),
.B(n_361),
.Y(n_523)
);

AOI22xp33_ASAP7_75t_L g524 ( 
.A1(n_463),
.A2(n_382),
.B1(n_357),
.B2(n_339),
.Y(n_524)
);

INVx4_ASAP7_75t_SL g525 ( 
.A(n_428),
.Y(n_525)
);

NAND2xp5_ASAP7_75t_L g526 ( 
.A(n_462),
.B(n_363),
.Y(n_526)
);

INVx1_ASAP7_75t_L g527 ( 
.A(n_463),
.Y(n_527)
);

INVx2_ASAP7_75t_L g528 ( 
.A(n_410),
.Y(n_528)
);

BUFx3_ASAP7_75t_L g529 ( 
.A(n_467),
.Y(n_529)
);

INVx1_ASAP7_75t_L g530 ( 
.A(n_444),
.Y(n_530)
);

INVx5_ASAP7_75t_L g531 ( 
.A(n_428),
.Y(n_531)
);

AOI22xp33_ASAP7_75t_L g532 ( 
.A1(n_446),
.A2(n_370),
.B1(n_344),
.B2(n_279),
.Y(n_532)
);

INVx2_ASAP7_75t_L g533 ( 
.A(n_421),
.Y(n_533)
);

NAND2xp5_ASAP7_75t_SL g534 ( 
.A(n_432),
.B(n_363),
.Y(n_534)
);

INVx1_ASAP7_75t_L g535 ( 
.A(n_448),
.Y(n_535)
);

NAND2xp5_ASAP7_75t_L g536 ( 
.A(n_467),
.B(n_366),
.Y(n_536)
);

INVx2_ASAP7_75t_L g537 ( 
.A(n_421),
.Y(n_537)
);

NAND2xp5_ASAP7_75t_L g538 ( 
.A(n_467),
.B(n_366),
.Y(n_538)
);

INVx4_ASAP7_75t_L g539 ( 
.A(n_428),
.Y(n_539)
);

NAND2xp33_ASAP7_75t_SL g540 ( 
.A(n_451),
.B(n_372),
.Y(n_540)
);

BUFx6f_ASAP7_75t_L g541 ( 
.A(n_406),
.Y(n_541)
);

NAND2xp33_ASAP7_75t_L g542 ( 
.A(n_451),
.B(n_372),
.Y(n_542)
);

AOI22xp5_ASAP7_75t_L g543 ( 
.A1(n_453),
.A2(n_378),
.B1(n_379),
.B2(n_390),
.Y(n_543)
);

OAI22xp33_ASAP7_75t_L g544 ( 
.A1(n_478),
.A2(n_453),
.B1(n_469),
.B2(n_459),
.Y(n_544)
);

AOI21xp5_ASAP7_75t_L g545 ( 
.A1(n_475),
.A2(n_452),
.B(n_449),
.Y(n_545)
);

NAND2xp5_ASAP7_75t_L g546 ( 
.A(n_511),
.B(n_496),
.Y(n_546)
);

INVx1_ASAP7_75t_L g547 ( 
.A(n_499),
.Y(n_547)
);

INVx5_ASAP7_75t_L g548 ( 
.A(n_539),
.Y(n_548)
);

INVx2_ASAP7_75t_L g549 ( 
.A(n_516),
.Y(n_549)
);

INVx2_ASAP7_75t_L g550 ( 
.A(n_516),
.Y(n_550)
);

INVx1_ASAP7_75t_L g551 ( 
.A(n_499),
.Y(n_551)
);

INVx1_ASAP7_75t_L g552 ( 
.A(n_499),
.Y(n_552)
);

NAND2xp5_ASAP7_75t_L g553 ( 
.A(n_511),
.B(n_458),
.Y(n_553)
);

INVx2_ASAP7_75t_L g554 ( 
.A(n_481),
.Y(n_554)
);

NOR2xp33_ASAP7_75t_L g555 ( 
.A(n_486),
.B(n_454),
.Y(n_555)
);

INVx5_ASAP7_75t_L g556 ( 
.A(n_539),
.Y(n_556)
);

OR2x6_ASAP7_75t_L g557 ( 
.A(n_512),
.B(n_438),
.Y(n_557)
);

NAND2xp5_ASAP7_75t_L g558 ( 
.A(n_496),
.B(n_436),
.Y(n_558)
);

NAND2xp5_ASAP7_75t_L g559 ( 
.A(n_486),
.B(n_420),
.Y(n_559)
);

AOI22xp33_ASAP7_75t_L g560 ( 
.A1(n_480),
.A2(n_473),
.B1(n_474),
.B2(n_532),
.Y(n_560)
);

NOR2xp33_ASAP7_75t_L g561 ( 
.A(n_514),
.B(n_454),
.Y(n_561)
);

NOR2xp33_ASAP7_75t_L g562 ( 
.A(n_514),
.B(n_457),
.Y(n_562)
);

NAND2xp5_ASAP7_75t_SL g563 ( 
.A(n_474),
.B(n_480),
.Y(n_563)
);

NOR2xp33_ASAP7_75t_L g564 ( 
.A(n_484),
.B(n_457),
.Y(n_564)
);

AND2x2_ASAP7_75t_L g565 ( 
.A(n_485),
.B(n_459),
.Y(n_565)
);

INVx1_ASAP7_75t_L g566 ( 
.A(n_481),
.Y(n_566)
);

NOR2xp33_ASAP7_75t_L g567 ( 
.A(n_484),
.B(n_469),
.Y(n_567)
);

AOI22xp33_ASAP7_75t_L g568 ( 
.A1(n_473),
.A2(n_369),
.B1(n_355),
.B2(n_443),
.Y(n_568)
);

NAND2xp5_ASAP7_75t_SL g569 ( 
.A(n_492),
.B(n_447),
.Y(n_569)
);

NOR2xp33_ASAP7_75t_L g570 ( 
.A(n_534),
.B(n_378),
.Y(n_570)
);

NAND2xp5_ASAP7_75t_SL g571 ( 
.A(n_543),
.B(n_379),
.Y(n_571)
);

INVxp33_ASAP7_75t_L g572 ( 
.A(n_510),
.Y(n_572)
);

INVx1_ASAP7_75t_L g573 ( 
.A(n_491),
.Y(n_573)
);

NAND2xp5_ASAP7_75t_L g574 ( 
.A(n_522),
.B(n_436),
.Y(n_574)
);

INVx1_ASAP7_75t_L g575 ( 
.A(n_491),
.Y(n_575)
);

NOR2xp33_ASAP7_75t_L g576 ( 
.A(n_534),
.B(n_384),
.Y(n_576)
);

AOI22xp5_ASAP7_75t_L g577 ( 
.A1(n_473),
.A2(n_384),
.B1(n_385),
.B2(n_386),
.Y(n_577)
);

NOR2xp33_ASAP7_75t_L g578 ( 
.A(n_477),
.B(n_385),
.Y(n_578)
);

NAND2xp5_ASAP7_75t_L g579 ( 
.A(n_522),
.B(n_386),
.Y(n_579)
);

AO22x1_ASAP7_75t_L g580 ( 
.A1(n_473),
.A2(n_403),
.B1(n_413),
.B2(n_414),
.Y(n_580)
);

INVx1_ASAP7_75t_L g581 ( 
.A(n_501),
.Y(n_581)
);

NAND2xp5_ASAP7_75t_L g582 ( 
.A(n_473),
.B(n_390),
.Y(n_582)
);

NAND2xp33_ASAP7_75t_L g583 ( 
.A(n_506),
.B(n_400),
.Y(n_583)
);

NAND2xp5_ASAP7_75t_L g584 ( 
.A(n_495),
.B(n_373),
.Y(n_584)
);

OAI22xp5_ASAP7_75t_SL g585 ( 
.A1(n_521),
.A2(n_423),
.B1(n_405),
.B2(n_412),
.Y(n_585)
);

AOI22xp5_ASAP7_75t_L g586 ( 
.A1(n_489),
.A2(n_471),
.B1(n_387),
.B2(n_395),
.Y(n_586)
);

INVx2_ASAP7_75t_L g587 ( 
.A(n_501),
.Y(n_587)
);

INVx1_ASAP7_75t_L g588 ( 
.A(n_479),
.Y(n_588)
);

NAND2xp5_ASAP7_75t_L g589 ( 
.A(n_495),
.B(n_439),
.Y(n_589)
);

AOI22xp5_ASAP7_75t_L g590 ( 
.A1(n_489),
.A2(n_278),
.B1(n_248),
.B2(n_250),
.Y(n_590)
);

INVx2_ASAP7_75t_L g591 ( 
.A(n_518),
.Y(n_591)
);

AND2x4_ASAP7_75t_SL g592 ( 
.A(n_482),
.B(n_422),
.Y(n_592)
);

NAND2xp5_ASAP7_75t_L g593 ( 
.A(n_529),
.B(n_439),
.Y(n_593)
);

NAND2xp5_ASAP7_75t_L g594 ( 
.A(n_505),
.B(n_443),
.Y(n_594)
);

O2A1O1Ixp5_ASAP7_75t_L g595 ( 
.A1(n_523),
.A2(n_425),
.B(n_435),
.C(n_408),
.Y(n_595)
);

NOR2xp33_ASAP7_75t_L g596 ( 
.A(n_487),
.B(n_414),
.Y(n_596)
);

AND2x2_ASAP7_75t_SL g597 ( 
.A(n_490),
.B(n_422),
.Y(n_597)
);

NAND2xp5_ASAP7_75t_SL g598 ( 
.A(n_508),
.B(n_282),
.Y(n_598)
);

AND2x6_ASAP7_75t_L g599 ( 
.A(n_503),
.B(n_208),
.Y(n_599)
);

INVx2_ASAP7_75t_L g600 ( 
.A(n_518),
.Y(n_600)
);

INVx1_ASAP7_75t_L g601 ( 
.A(n_483),
.Y(n_601)
);

NAND2xp5_ASAP7_75t_L g602 ( 
.A(n_505),
.B(n_408),
.Y(n_602)
);

AND2x2_ASAP7_75t_SL g603 ( 
.A(n_494),
.B(n_419),
.Y(n_603)
);

INVx2_ASAP7_75t_SL g604 ( 
.A(n_503),
.Y(n_604)
);

NAND2xp5_ASAP7_75t_L g605 ( 
.A(n_529),
.B(n_408),
.Y(n_605)
);

AOI21xp5_ASAP7_75t_L g606 ( 
.A1(n_476),
.A2(n_435),
.B(n_425),
.Y(n_606)
);

NAND2xp5_ASAP7_75t_SL g607 ( 
.A(n_487),
.B(n_287),
.Y(n_607)
);

HB1xp67_ASAP7_75t_L g608 ( 
.A(n_493),
.Y(n_608)
);

NAND2xp5_ASAP7_75t_L g609 ( 
.A(n_526),
.B(n_428),
.Y(n_609)
);

NAND2xp5_ASAP7_75t_SL g610 ( 
.A(n_536),
.B(n_289),
.Y(n_610)
);

INVx2_ASAP7_75t_L g611 ( 
.A(n_528),
.Y(n_611)
);

NAND2xp5_ASAP7_75t_L g612 ( 
.A(n_538),
.B(n_291),
.Y(n_612)
);

INVx1_ASAP7_75t_L g613 ( 
.A(n_498),
.Y(n_613)
);

OR2x6_ASAP7_75t_L g614 ( 
.A(n_512),
.B(n_419),
.Y(n_614)
);

NAND2xp5_ASAP7_75t_L g615 ( 
.A(n_517),
.B(n_406),
.Y(n_615)
);

INVxp67_ASAP7_75t_SL g616 ( 
.A(n_507),
.Y(n_616)
);

NAND2xp5_ASAP7_75t_L g617 ( 
.A(n_520),
.B(n_406),
.Y(n_617)
);

INVx1_ASAP7_75t_L g618 ( 
.A(n_500),
.Y(n_618)
);

OR2x2_ASAP7_75t_L g619 ( 
.A(n_512),
.B(n_412),
.Y(n_619)
);

NOR2xp33_ASAP7_75t_L g620 ( 
.A(n_542),
.B(n_423),
.Y(n_620)
);

AND2x2_ASAP7_75t_L g621 ( 
.A(n_482),
.B(n_296),
.Y(n_621)
);

AND2x2_ASAP7_75t_SL g622 ( 
.A(n_542),
.B(n_430),
.Y(n_622)
);

BUFx3_ASAP7_75t_L g623 ( 
.A(n_519),
.Y(n_623)
);

AOI21xp5_ASAP7_75t_L g624 ( 
.A1(n_502),
.A2(n_219),
.B(n_218),
.Y(n_624)
);

INVx1_ASAP7_75t_L g625 ( 
.A(n_504),
.Y(n_625)
);

NAND2xp5_ASAP7_75t_L g626 ( 
.A(n_527),
.B(n_430),
.Y(n_626)
);

INVx1_ASAP7_75t_L g627 ( 
.A(n_509),
.Y(n_627)
);

INVx1_ASAP7_75t_L g628 ( 
.A(n_515),
.Y(n_628)
);

INVx1_ASAP7_75t_L g629 ( 
.A(n_530),
.Y(n_629)
);

OAI22xp5_ASAP7_75t_L g630 ( 
.A1(n_524),
.A2(n_299),
.B1(n_221),
.B2(n_223),
.Y(n_630)
);

NAND2xp5_ASAP7_75t_SL g631 ( 
.A(n_540),
.B(n_220),
.Y(n_631)
);

BUFx2_ASAP7_75t_L g632 ( 
.A(n_540),
.Y(n_632)
);

AOI22xp33_ASAP7_75t_L g633 ( 
.A1(n_532),
.A2(n_468),
.B1(n_433),
.B2(n_430),
.Y(n_633)
);

NAND2xp5_ASAP7_75t_L g634 ( 
.A(n_535),
.B(n_430),
.Y(n_634)
);

NAND2xp5_ASAP7_75t_L g635 ( 
.A(n_528),
.B(n_533),
.Y(n_635)
);

OAI221xp5_ASAP7_75t_L g636 ( 
.A1(n_524),
.A2(n_302),
.B1(n_225),
.B2(n_227),
.C(n_239),
.Y(n_636)
);

BUFx5_ASAP7_75t_L g637 ( 
.A(n_488),
.Y(n_637)
);

NOR2x1p5_ASAP7_75t_L g638 ( 
.A(n_519),
.B(n_224),
.Y(n_638)
);

INVx2_ASAP7_75t_L g639 ( 
.A(n_533),
.Y(n_639)
);

NAND2x1_ASAP7_75t_L g640 ( 
.A(n_507),
.B(n_468),
.Y(n_640)
);

AND2x2_ASAP7_75t_L g641 ( 
.A(n_537),
.B(n_430),
.Y(n_641)
);

NOR2xp33_ASAP7_75t_L g642 ( 
.A(n_555),
.B(n_537),
.Y(n_642)
);

AOI21xp5_ASAP7_75t_L g643 ( 
.A1(n_546),
.A2(n_541),
.B(n_507),
.Y(n_643)
);

AOI21xp5_ASAP7_75t_L g644 ( 
.A1(n_546),
.A2(n_541),
.B(n_507),
.Y(n_644)
);

NAND3xp33_ASAP7_75t_SL g645 ( 
.A(n_564),
.B(n_567),
.C(n_562),
.Y(n_645)
);

O2A1O1Ixp33_ASAP7_75t_L g646 ( 
.A1(n_561),
.A2(n_8),
.B(n_9),
.C(n_11),
.Y(n_646)
);

NAND2xp5_ASAP7_75t_L g647 ( 
.A(n_553),
.B(n_541),
.Y(n_647)
);

AOI21xp5_ASAP7_75t_L g648 ( 
.A1(n_553),
.A2(n_541),
.B(n_531),
.Y(n_648)
);

AND2x2_ASAP7_75t_L g649 ( 
.A(n_565),
.B(n_513),
.Y(n_649)
);

INVx2_ASAP7_75t_L g650 ( 
.A(n_554),
.Y(n_650)
);

NAND2xp5_ASAP7_75t_L g651 ( 
.A(n_589),
.B(n_513),
.Y(n_651)
);

AOI21xp5_ASAP7_75t_L g652 ( 
.A1(n_609),
.A2(n_531),
.B(n_497),
.Y(n_652)
);

INVx1_ASAP7_75t_L g653 ( 
.A(n_588),
.Y(n_653)
);

NOR2xp33_ASAP7_75t_L g654 ( 
.A(n_572),
.B(n_243),
.Y(n_654)
);

NAND2x1p5_ASAP7_75t_L g655 ( 
.A(n_548),
.B(n_556),
.Y(n_655)
);

INVx1_ASAP7_75t_L g656 ( 
.A(n_601),
.Y(n_656)
);

NAND2xp5_ASAP7_75t_L g657 ( 
.A(n_594),
.B(n_513),
.Y(n_657)
);

AOI21xp5_ASAP7_75t_L g658 ( 
.A1(n_605),
.A2(n_531),
.B(n_497),
.Y(n_658)
);

NAND2x1p5_ASAP7_75t_L g659 ( 
.A(n_548),
.B(n_497),
.Y(n_659)
);

CKINVDCx5p33_ASAP7_75t_R g660 ( 
.A(n_623),
.Y(n_660)
);

AND2x2_ASAP7_75t_L g661 ( 
.A(n_597),
.B(n_525),
.Y(n_661)
);

AOI21xp5_ASAP7_75t_L g662 ( 
.A1(n_548),
.A2(n_531),
.B(n_497),
.Y(n_662)
);

INVx1_ASAP7_75t_L g663 ( 
.A(n_613),
.Y(n_663)
);

NAND2xp5_ASAP7_75t_L g664 ( 
.A(n_584),
.B(n_525),
.Y(n_664)
);

AOI21xp5_ASAP7_75t_L g665 ( 
.A1(n_548),
.A2(n_272),
.B(n_247),
.Y(n_665)
);

NAND2xp5_ASAP7_75t_SL g666 ( 
.A(n_560),
.B(n_525),
.Y(n_666)
);

O2A1O1Ixp33_ASAP7_75t_L g667 ( 
.A1(n_544),
.A2(n_9),
.B(n_12),
.C(n_13),
.Y(n_667)
);

NAND2xp5_ASAP7_75t_L g668 ( 
.A(n_578),
.B(n_433),
.Y(n_668)
);

AOI21x1_ASAP7_75t_L g669 ( 
.A1(n_635),
.A2(n_606),
.B(n_626),
.Y(n_669)
);

OAI22xp5_ASAP7_75t_L g670 ( 
.A1(n_582),
.A2(n_304),
.B1(n_251),
.B2(n_253),
.Y(n_670)
);

NAND2xp5_ASAP7_75t_L g671 ( 
.A(n_559),
.B(n_433),
.Y(n_671)
);

AOI21xp5_ASAP7_75t_L g672 ( 
.A1(n_556),
.A2(n_273),
.B(n_255),
.Y(n_672)
);

AOI21xp5_ASAP7_75t_L g673 ( 
.A1(n_556),
.A2(n_274),
.B(n_256),
.Y(n_673)
);

OAI21xp5_ASAP7_75t_L g674 ( 
.A1(n_595),
.A2(n_468),
.B(n_283),
.Y(n_674)
);

NOR2xp33_ASAP7_75t_L g675 ( 
.A(n_563),
.B(n_14),
.Y(n_675)
);

AOI21xp5_ASAP7_75t_L g676 ( 
.A1(n_556),
.A2(n_271),
.B(n_257),
.Y(n_676)
);

AO21x1_ASAP7_75t_L g677 ( 
.A1(n_570),
.A2(n_433),
.B(n_468),
.Y(n_677)
);

INVx1_ASAP7_75t_L g678 ( 
.A(n_618),
.Y(n_678)
);

NAND2xp5_ASAP7_75t_L g679 ( 
.A(n_576),
.B(n_433),
.Y(n_679)
);

INVx1_ASAP7_75t_L g680 ( 
.A(n_625),
.Y(n_680)
);

AOI21xp5_ASAP7_75t_L g681 ( 
.A1(n_593),
.A2(n_545),
.B(n_558),
.Y(n_681)
);

AOI21xp5_ASAP7_75t_L g682 ( 
.A1(n_593),
.A2(n_285),
.B(n_300),
.Y(n_682)
);

NOR2xp33_ASAP7_75t_L g683 ( 
.A(n_579),
.B(n_14),
.Y(n_683)
);

OAI22xp5_ASAP7_75t_L g684 ( 
.A1(n_582),
.A2(n_245),
.B1(n_260),
.B2(n_261),
.Y(n_684)
);

AOI21xp5_ASAP7_75t_L g685 ( 
.A1(n_558),
.A2(n_288),
.B(n_297),
.Y(n_685)
);

OAI22xp5_ASAP7_75t_L g686 ( 
.A1(n_579),
.A2(n_265),
.B1(n_266),
.B2(n_267),
.Y(n_686)
);

AND2x4_ASAP7_75t_L g687 ( 
.A(n_604),
.B(n_468),
.Y(n_687)
);

AOI21xp5_ASAP7_75t_L g688 ( 
.A1(n_574),
.A2(n_295),
.B(n_294),
.Y(n_688)
);

AOI21xp5_ASAP7_75t_L g689 ( 
.A1(n_574),
.A2(n_290),
.B(n_269),
.Y(n_689)
);

AOI21xp5_ASAP7_75t_L g690 ( 
.A1(n_602),
.A2(n_468),
.B(n_85),
.Y(n_690)
);

NAND2xp5_ASAP7_75t_L g691 ( 
.A(n_627),
.B(n_16),
.Y(n_691)
);

AOI21xp5_ASAP7_75t_L g692 ( 
.A1(n_566),
.A2(n_84),
.B(n_185),
.Y(n_692)
);

NOR3xp33_ASAP7_75t_L g693 ( 
.A(n_620),
.B(n_17),
.C(n_18),
.Y(n_693)
);

NAND2xp5_ASAP7_75t_L g694 ( 
.A(n_628),
.B(n_20),
.Y(n_694)
);

INVx1_ASAP7_75t_L g695 ( 
.A(n_629),
.Y(n_695)
);

INVx3_ASAP7_75t_L g696 ( 
.A(n_640),
.Y(n_696)
);

NAND2xp5_ASAP7_75t_L g697 ( 
.A(n_612),
.B(n_20),
.Y(n_697)
);

INVx2_ASAP7_75t_L g698 ( 
.A(n_587),
.Y(n_698)
);

AND2x2_ASAP7_75t_SL g699 ( 
.A(n_622),
.B(n_603),
.Y(n_699)
);

INVx1_ASAP7_75t_L g700 ( 
.A(n_573),
.Y(n_700)
);

AOI21xp5_ASAP7_75t_L g701 ( 
.A1(n_575),
.A2(n_581),
.B(n_610),
.Y(n_701)
);

INVx3_ASAP7_75t_L g702 ( 
.A(n_549),
.Y(n_702)
);

AOI21xp5_ASAP7_75t_L g703 ( 
.A1(n_635),
.A2(n_101),
.B(n_184),
.Y(n_703)
);

OAI21xp5_ASAP7_75t_L g704 ( 
.A1(n_634),
.A2(n_100),
.B(n_183),
.Y(n_704)
);

OAI21xp33_ASAP7_75t_L g705 ( 
.A1(n_577),
.A2(n_21),
.B(n_22),
.Y(n_705)
);

OAI21xp5_ASAP7_75t_L g706 ( 
.A1(n_634),
.A2(n_82),
.B(n_181),
.Y(n_706)
);

NOR2x1p5_ASAP7_75t_SL g707 ( 
.A(n_637),
.B(n_44),
.Y(n_707)
);

NAND2xp5_ASAP7_75t_L g708 ( 
.A(n_547),
.B(n_22),
.Y(n_708)
);

AND2x2_ASAP7_75t_L g709 ( 
.A(n_557),
.B(n_24),
.Y(n_709)
);

AOI21xp5_ASAP7_75t_L g710 ( 
.A1(n_550),
.A2(n_616),
.B(n_626),
.Y(n_710)
);

OAI21xp5_ASAP7_75t_L g711 ( 
.A1(n_615),
.A2(n_105),
.B(n_180),
.Y(n_711)
);

AOI21x1_ASAP7_75t_L g712 ( 
.A1(n_615),
.A2(n_103),
.B(n_179),
.Y(n_712)
);

O2A1O1Ixp5_ASAP7_75t_L g713 ( 
.A1(n_607),
.A2(n_25),
.B(n_26),
.C(n_27),
.Y(n_713)
);

A2O1A1Ixp33_ASAP7_75t_L g714 ( 
.A1(n_596),
.A2(n_27),
.B(n_29),
.C(n_30),
.Y(n_714)
);

AOI21xp5_ASAP7_75t_L g715 ( 
.A1(n_617),
.A2(n_110),
.B(n_177),
.Y(n_715)
);

INVx1_ASAP7_75t_L g716 ( 
.A(n_551),
.Y(n_716)
);

AOI21xp5_ASAP7_75t_L g717 ( 
.A1(n_617),
.A2(n_106),
.B(n_175),
.Y(n_717)
);

OAI21xp5_ASAP7_75t_L g718 ( 
.A1(n_641),
.A2(n_81),
.B(n_174),
.Y(n_718)
);

OAI21xp5_ASAP7_75t_L g719 ( 
.A1(n_591),
.A2(n_79),
.B(n_173),
.Y(n_719)
);

HB1xp67_ASAP7_75t_L g720 ( 
.A(n_557),
.Y(n_720)
);

INVx1_ASAP7_75t_L g721 ( 
.A(n_552),
.Y(n_721)
);

O2A1O1Ixp33_ASAP7_75t_L g722 ( 
.A1(n_583),
.A2(n_31),
.B(n_32),
.C(n_33),
.Y(n_722)
);

AOI21xp5_ASAP7_75t_L g723 ( 
.A1(n_600),
.A2(n_113),
.B(n_172),
.Y(n_723)
);

OAI22xp5_ASAP7_75t_L g724 ( 
.A1(n_632),
.A2(n_32),
.B1(n_34),
.B2(n_35),
.Y(n_724)
);

NAND2xp5_ASAP7_75t_L g725 ( 
.A(n_599),
.B(n_34),
.Y(n_725)
);

O2A1O1Ixp33_ASAP7_75t_L g726 ( 
.A1(n_571),
.A2(n_36),
.B(n_37),
.C(n_38),
.Y(n_726)
);

NAND2xp5_ASAP7_75t_L g727 ( 
.A(n_599),
.B(n_36),
.Y(n_727)
);

NAND2xp5_ASAP7_75t_L g728 ( 
.A(n_599),
.B(n_37),
.Y(n_728)
);

HB1xp67_ASAP7_75t_L g729 ( 
.A(n_557),
.Y(n_729)
);

AOI21xp5_ASAP7_75t_L g730 ( 
.A1(n_611),
.A2(n_119),
.B(n_170),
.Y(n_730)
);

NAND2xp5_ASAP7_75t_SL g731 ( 
.A(n_568),
.B(n_38),
.Y(n_731)
);

OAI21xp5_ASAP7_75t_L g732 ( 
.A1(n_639),
.A2(n_118),
.B(n_165),
.Y(n_732)
);

AOI21xp5_ASAP7_75t_L g733 ( 
.A1(n_631),
.A2(n_117),
.B(n_159),
.Y(n_733)
);

AOI21xp5_ASAP7_75t_L g734 ( 
.A1(n_598),
.A2(n_78),
.B(n_157),
.Y(n_734)
);

AOI21xp5_ASAP7_75t_L g735 ( 
.A1(n_624),
.A2(n_77),
.B(n_156),
.Y(n_735)
);

AO21x1_ASAP7_75t_L g736 ( 
.A1(n_630),
.A2(n_190),
.B(n_75),
.Y(n_736)
);

NOR2xp33_ASAP7_75t_L g737 ( 
.A(n_569),
.B(n_39),
.Y(n_737)
);

AOI21xp5_ASAP7_75t_L g738 ( 
.A1(n_647),
.A2(n_586),
.B(n_621),
.Y(n_738)
);

NOR2xp33_ASAP7_75t_L g739 ( 
.A(n_645),
.B(n_608),
.Y(n_739)
);

NAND2xp5_ASAP7_75t_L g740 ( 
.A(n_645),
.B(n_599),
.Y(n_740)
);

AOI21xp5_ASAP7_75t_L g741 ( 
.A1(n_642),
.A2(n_637),
.B(n_580),
.Y(n_741)
);

AND3x4_ASAP7_75t_L g742 ( 
.A(n_693),
.B(n_592),
.C(n_614),
.Y(n_742)
);

AOI21xp5_ASAP7_75t_L g743 ( 
.A1(n_642),
.A2(n_637),
.B(n_636),
.Y(n_743)
);

OAI21x1_ASAP7_75t_L g744 ( 
.A1(n_669),
.A2(n_633),
.B(n_638),
.Y(n_744)
);

INVx1_ASAP7_75t_SL g745 ( 
.A(n_660),
.Y(n_745)
);

OAI21xp5_ASAP7_75t_L g746 ( 
.A1(n_681),
.A2(n_630),
.B(n_590),
.Y(n_746)
);

CKINVDCx16_ASAP7_75t_R g747 ( 
.A(n_720),
.Y(n_747)
);

AOI21xp5_ASAP7_75t_L g748 ( 
.A1(n_643),
.A2(n_637),
.B(n_614),
.Y(n_748)
);

INVx1_ASAP7_75t_L g749 ( 
.A(n_653),
.Y(n_749)
);

BUFx2_ASAP7_75t_L g750 ( 
.A(n_720),
.Y(n_750)
);

AOI21xp5_ASAP7_75t_L g751 ( 
.A1(n_644),
.A2(n_637),
.B(n_614),
.Y(n_751)
);

OAI21x1_ASAP7_75t_SL g752 ( 
.A1(n_736),
.A2(n_701),
.B(n_722),
.Y(n_752)
);

INVx2_ASAP7_75t_L g753 ( 
.A(n_650),
.Y(n_753)
);

INVxp67_ASAP7_75t_L g754 ( 
.A(n_737),
.Y(n_754)
);

OAI21xp5_ASAP7_75t_L g755 ( 
.A1(n_710),
.A2(n_637),
.B(n_619),
.Y(n_755)
);

OAI22x1_ASAP7_75t_L g756 ( 
.A1(n_731),
.A2(n_585),
.B1(n_40),
.B2(n_39),
.Y(n_756)
);

INVx1_ASAP7_75t_L g757 ( 
.A(n_656),
.Y(n_757)
);

OAI21x1_ASAP7_75t_L g758 ( 
.A1(n_719),
.A2(n_45),
.B(n_47),
.Y(n_758)
);

NAND2xp5_ASAP7_75t_L g759 ( 
.A(n_699),
.B(n_48),
.Y(n_759)
);

OAI21xp5_ASAP7_75t_L g760 ( 
.A1(n_697),
.A2(n_50),
.B(n_51),
.Y(n_760)
);

NOR2x1_ASAP7_75t_SL g761 ( 
.A(n_664),
.B(n_55),
.Y(n_761)
);

A2O1A1Ixp33_ASAP7_75t_L g762 ( 
.A1(n_683),
.A2(n_56),
.B(n_59),
.C(n_62),
.Y(n_762)
);

OAI21x1_ASAP7_75t_L g763 ( 
.A1(n_732),
.A2(n_67),
.B(n_68),
.Y(n_763)
);

OAI21xp5_ASAP7_75t_L g764 ( 
.A1(n_648),
.A2(n_71),
.B(n_73),
.Y(n_764)
);

BUFx12f_ASAP7_75t_L g765 ( 
.A(n_709),
.Y(n_765)
);

AOI21xp5_ASAP7_75t_L g766 ( 
.A1(n_668),
.A2(n_74),
.B(n_121),
.Y(n_766)
);

INVx3_ASAP7_75t_SL g767 ( 
.A(n_699),
.Y(n_767)
);

INVx1_ASAP7_75t_L g768 ( 
.A(n_663),
.Y(n_768)
);

INVx2_ASAP7_75t_L g769 ( 
.A(n_698),
.Y(n_769)
);

INVx1_ASAP7_75t_L g770 ( 
.A(n_678),
.Y(n_770)
);

AOI21xp5_ASAP7_75t_L g771 ( 
.A1(n_679),
.A2(n_123),
.B(n_124),
.Y(n_771)
);

AND2x2_ASAP7_75t_L g772 ( 
.A(n_680),
.B(n_127),
.Y(n_772)
);

OAI21x1_ASAP7_75t_L g773 ( 
.A1(n_704),
.A2(n_128),
.B(n_129),
.Y(n_773)
);

AND2x4_ASAP7_75t_L g774 ( 
.A(n_661),
.B(n_130),
.Y(n_774)
);

INVx1_ASAP7_75t_L g775 ( 
.A(n_695),
.Y(n_775)
);

NAND2xp5_ASAP7_75t_L g776 ( 
.A(n_683),
.B(n_649),
.Y(n_776)
);

OAI21x1_ASAP7_75t_L g777 ( 
.A1(n_706),
.A2(n_131),
.B(n_132),
.Y(n_777)
);

OAI21x1_ASAP7_75t_L g778 ( 
.A1(n_711),
.A2(n_141),
.B(n_148),
.Y(n_778)
);

CKINVDCx6p67_ASAP7_75t_R g779 ( 
.A(n_729),
.Y(n_779)
);

BUFx2_ASAP7_75t_L g780 ( 
.A(n_729),
.Y(n_780)
);

INVx1_ASAP7_75t_L g781 ( 
.A(n_700),
.Y(n_781)
);

NAND2xp5_ASAP7_75t_L g782 ( 
.A(n_737),
.B(n_149),
.Y(n_782)
);

NAND2xp5_ASAP7_75t_L g783 ( 
.A(n_675),
.B(n_150),
.Y(n_783)
);

AOI21xp5_ASAP7_75t_L g784 ( 
.A1(n_651),
.A2(n_153),
.B(n_155),
.Y(n_784)
);

OAI21xp5_ASAP7_75t_L g785 ( 
.A1(n_674),
.A2(n_671),
.B(n_682),
.Y(n_785)
);

INVx1_ASAP7_75t_L g786 ( 
.A(n_716),
.Y(n_786)
);

OAI21xp5_ASAP7_75t_L g787 ( 
.A1(n_685),
.A2(n_688),
.B(n_689),
.Y(n_787)
);

INVx2_ASAP7_75t_SL g788 ( 
.A(n_687),
.Y(n_788)
);

NAND2xp5_ASAP7_75t_L g789 ( 
.A(n_675),
.B(n_654),
.Y(n_789)
);

NOR2x1_ASAP7_75t_SL g790 ( 
.A(n_666),
.B(n_657),
.Y(n_790)
);

INVx2_ASAP7_75t_L g791 ( 
.A(n_702),
.Y(n_791)
);

NAND2xp5_ASAP7_75t_L g792 ( 
.A(n_702),
.B(n_691),
.Y(n_792)
);

OAI21x1_ASAP7_75t_L g793 ( 
.A1(n_718),
.A2(n_712),
.B(n_677),
.Y(n_793)
);

OAI21x1_ASAP7_75t_L g794 ( 
.A1(n_652),
.A2(n_703),
.B(n_690),
.Y(n_794)
);

NAND2xp5_ASAP7_75t_L g795 ( 
.A(n_694),
.B(n_721),
.Y(n_795)
);

INVx1_ASAP7_75t_L g796 ( 
.A(n_708),
.Y(n_796)
);

INVx2_ASAP7_75t_L g797 ( 
.A(n_696),
.Y(n_797)
);

AND2x2_ASAP7_75t_L g798 ( 
.A(n_693),
.B(n_687),
.Y(n_798)
);

AOI21xp5_ASAP7_75t_L g799 ( 
.A1(n_655),
.A2(n_658),
.B(n_735),
.Y(n_799)
);

NAND2x1p5_ASAP7_75t_L g800 ( 
.A(n_696),
.B(n_734),
.Y(n_800)
);

OAI21x1_ASAP7_75t_L g801 ( 
.A1(n_715),
.A2(n_717),
.B(n_692),
.Y(n_801)
);

NAND2xp5_ASAP7_75t_L g802 ( 
.A(n_686),
.B(n_705),
.Y(n_802)
);

INVx1_ASAP7_75t_L g803 ( 
.A(n_749),
.Y(n_803)
);

NAND2xp5_ASAP7_75t_L g804 ( 
.A(n_789),
.B(n_724),
.Y(n_804)
);

INVx1_ASAP7_75t_L g805 ( 
.A(n_757),
.Y(n_805)
);

NAND2xp5_ASAP7_75t_L g806 ( 
.A(n_754),
.B(n_714),
.Y(n_806)
);

INVx3_ASAP7_75t_SL g807 ( 
.A(n_745),
.Y(n_807)
);

INVx3_ASAP7_75t_L g808 ( 
.A(n_774),
.Y(n_808)
);

O2A1O1Ixp33_ASAP7_75t_L g809 ( 
.A1(n_746),
.A2(n_646),
.B(n_667),
.C(n_726),
.Y(n_809)
);

AOI221xp5_ASAP7_75t_L g810 ( 
.A1(n_756),
.A2(n_739),
.B1(n_802),
.B2(n_775),
.C(n_770),
.Y(n_810)
);

NOR2xp33_ASAP7_75t_L g811 ( 
.A(n_767),
.B(n_684),
.Y(n_811)
);

AND2x6_ASAP7_75t_L g812 ( 
.A(n_774),
.B(n_728),
.Y(n_812)
);

BUFx2_ASAP7_75t_L g813 ( 
.A(n_765),
.Y(n_813)
);

AND2x2_ASAP7_75t_L g814 ( 
.A(n_747),
.B(n_713),
.Y(n_814)
);

AOI22xp5_ASAP7_75t_L g815 ( 
.A1(n_742),
.A2(n_727),
.B1(n_725),
.B2(n_670),
.Y(n_815)
);

BUFx2_ASAP7_75t_SL g816 ( 
.A(n_774),
.Y(n_816)
);

NAND2xp5_ASAP7_75t_L g817 ( 
.A(n_739),
.B(n_676),
.Y(n_817)
);

NAND2xp5_ASAP7_75t_L g818 ( 
.A(n_767),
.B(n_768),
.Y(n_818)
);

NAND2xp5_ASAP7_75t_L g819 ( 
.A(n_776),
.B(n_673),
.Y(n_819)
);

NAND2xp5_ASAP7_75t_L g820 ( 
.A(n_750),
.B(n_780),
.Y(n_820)
);

AND2x2_ASAP7_75t_L g821 ( 
.A(n_765),
.B(n_713),
.Y(n_821)
);

INVx3_ASAP7_75t_L g822 ( 
.A(n_788),
.Y(n_822)
);

INVx1_ASAP7_75t_L g823 ( 
.A(n_781),
.Y(n_823)
);

INVx1_ASAP7_75t_L g824 ( 
.A(n_786),
.Y(n_824)
);

A2O1A1Ixp33_ASAP7_75t_SL g825 ( 
.A1(n_787),
.A2(n_733),
.B(n_730),
.C(n_723),
.Y(n_825)
);

O2A1O1Ixp33_ASAP7_75t_SL g826 ( 
.A1(n_762),
.A2(n_707),
.B(n_665),
.C(n_672),
.Y(n_826)
);

OA21x2_ASAP7_75t_L g827 ( 
.A1(n_793),
.A2(n_662),
.B(n_655),
.Y(n_827)
);

INVx3_ASAP7_75t_L g828 ( 
.A(n_788),
.Y(n_828)
);

INVx3_ASAP7_75t_L g829 ( 
.A(n_797),
.Y(n_829)
);

BUFx2_ASAP7_75t_L g830 ( 
.A(n_779),
.Y(n_830)
);

INVx1_ASAP7_75t_L g831 ( 
.A(n_753),
.Y(n_831)
);

INVx1_ASAP7_75t_L g832 ( 
.A(n_769),
.Y(n_832)
);

NAND2xp5_ASAP7_75t_L g833 ( 
.A(n_796),
.B(n_659),
.Y(n_833)
);

INVx3_ASAP7_75t_SL g834 ( 
.A(n_779),
.Y(n_834)
);

NAND2x1p5_ASAP7_75t_L g835 ( 
.A(n_798),
.B(n_659),
.Y(n_835)
);

NOR2xp33_ASAP7_75t_L g836 ( 
.A(n_798),
.B(n_795),
.Y(n_836)
);

INVx1_ASAP7_75t_L g837 ( 
.A(n_769),
.Y(n_837)
);

BUFx6f_ASAP7_75t_L g838 ( 
.A(n_797),
.Y(n_838)
);

INVx5_ASAP7_75t_L g839 ( 
.A(n_772),
.Y(n_839)
);

AND2x2_ASAP7_75t_L g840 ( 
.A(n_756),
.B(n_791),
.Y(n_840)
);

AOI22xp33_ASAP7_75t_L g841 ( 
.A1(n_742),
.A2(n_782),
.B1(n_783),
.B2(n_738),
.Y(n_841)
);

AOI21xp5_ASAP7_75t_L g842 ( 
.A1(n_743),
.A2(n_799),
.B(n_741),
.Y(n_842)
);

INVx1_ASAP7_75t_L g843 ( 
.A(n_772),
.Y(n_843)
);

NAND2xp5_ASAP7_75t_L g844 ( 
.A(n_792),
.B(n_759),
.Y(n_844)
);

AND2x4_ASAP7_75t_L g845 ( 
.A(n_755),
.B(n_748),
.Y(n_845)
);

HB1xp67_ASAP7_75t_L g846 ( 
.A(n_744),
.Y(n_846)
);

AOI22xp33_ASAP7_75t_L g847 ( 
.A1(n_760),
.A2(n_740),
.B1(n_752),
.B2(n_744),
.Y(n_847)
);

AOI21xp5_ASAP7_75t_L g848 ( 
.A1(n_785),
.A2(n_801),
.B(n_794),
.Y(n_848)
);

INVx2_ASAP7_75t_SL g849 ( 
.A(n_800),
.Y(n_849)
);

OR2x2_ASAP7_75t_L g850 ( 
.A(n_751),
.B(n_762),
.Y(n_850)
);

BUFx4_ASAP7_75t_SL g851 ( 
.A(n_761),
.Y(n_851)
);

INVx3_ASAP7_75t_SL g852 ( 
.A(n_790),
.Y(n_852)
);

INVx1_ASAP7_75t_L g853 ( 
.A(n_800),
.Y(n_853)
);

INVx1_ASAP7_75t_L g854 ( 
.A(n_778),
.Y(n_854)
);

AND2x4_ASAP7_75t_L g855 ( 
.A(n_764),
.B(n_784),
.Y(n_855)
);

AOI22xp33_ASAP7_75t_L g856 ( 
.A1(n_810),
.A2(n_804),
.B1(n_841),
.B2(n_836),
.Y(n_856)
);

AND2x2_ASAP7_75t_L g857 ( 
.A(n_836),
.B(n_777),
.Y(n_857)
);

BUFx8_ASAP7_75t_L g858 ( 
.A(n_813),
.Y(n_858)
);

INVx2_ASAP7_75t_L g859 ( 
.A(n_846),
.Y(n_859)
);

CKINVDCx11_ASAP7_75t_R g860 ( 
.A(n_807),
.Y(n_860)
);

OAI21x1_ASAP7_75t_L g861 ( 
.A1(n_848),
.A2(n_793),
.B(n_794),
.Y(n_861)
);

INVx1_ASAP7_75t_L g862 ( 
.A(n_846),
.Y(n_862)
);

INVx2_ASAP7_75t_L g863 ( 
.A(n_854),
.Y(n_863)
);

OA21x2_ASAP7_75t_L g864 ( 
.A1(n_842),
.A2(n_773),
.B(n_777),
.Y(n_864)
);

AO21x1_ASAP7_75t_L g865 ( 
.A1(n_850),
.A2(n_773),
.B(n_778),
.Y(n_865)
);

AND2x2_ASAP7_75t_L g866 ( 
.A(n_845),
.B(n_758),
.Y(n_866)
);

INVx3_ASAP7_75t_L g867 ( 
.A(n_845),
.Y(n_867)
);

AOI22xp33_ASAP7_75t_L g868 ( 
.A1(n_841),
.A2(n_758),
.B1(n_763),
.B2(n_766),
.Y(n_868)
);

OAI22xp5_ASAP7_75t_L g869 ( 
.A1(n_839),
.A2(n_771),
.B1(n_763),
.B2(n_801),
.Y(n_869)
);

INVx1_ASAP7_75t_L g870 ( 
.A(n_831),
.Y(n_870)
);

OAI22xp5_ASAP7_75t_L g871 ( 
.A1(n_839),
.A2(n_816),
.B1(n_806),
.B2(n_808),
.Y(n_871)
);

INVx1_ASAP7_75t_L g872 ( 
.A(n_832),
.Y(n_872)
);

INVx1_ASAP7_75t_L g873 ( 
.A(n_837),
.Y(n_873)
);

INVx2_ASAP7_75t_L g874 ( 
.A(n_853),
.Y(n_874)
);

INVx3_ASAP7_75t_L g875 ( 
.A(n_827),
.Y(n_875)
);

BUFx6f_ASAP7_75t_L g876 ( 
.A(n_839),
.Y(n_876)
);

INVx1_ASAP7_75t_L g877 ( 
.A(n_829),
.Y(n_877)
);

HB1xp67_ASAP7_75t_L g878 ( 
.A(n_849),
.Y(n_878)
);

INVx2_ASAP7_75t_L g879 ( 
.A(n_849),
.Y(n_879)
);

INVx1_ASAP7_75t_L g880 ( 
.A(n_829),
.Y(n_880)
);

INVx2_ASAP7_75t_L g881 ( 
.A(n_829),
.Y(n_881)
);

INVx1_ASAP7_75t_L g882 ( 
.A(n_803),
.Y(n_882)
);

BUFx2_ASAP7_75t_L g883 ( 
.A(n_839),
.Y(n_883)
);

AO21x1_ASAP7_75t_L g884 ( 
.A1(n_809),
.A2(n_855),
.B(n_817),
.Y(n_884)
);

OAI21x1_ASAP7_75t_L g885 ( 
.A1(n_847),
.A2(n_827),
.B(n_835),
.Y(n_885)
);

BUFx8_ASAP7_75t_L g886 ( 
.A(n_830),
.Y(n_886)
);

BUFx8_ASAP7_75t_SL g887 ( 
.A(n_820),
.Y(n_887)
);

INVx1_ASAP7_75t_L g888 ( 
.A(n_805),
.Y(n_888)
);

BUFx12f_ASAP7_75t_L g889 ( 
.A(n_838),
.Y(n_889)
);

INVx2_ASAP7_75t_L g890 ( 
.A(n_827),
.Y(n_890)
);

INVx2_ASAP7_75t_SL g891 ( 
.A(n_835),
.Y(n_891)
);

NAND2x1p5_ASAP7_75t_L g892 ( 
.A(n_808),
.B(n_855),
.Y(n_892)
);

BUFx3_ASAP7_75t_L g893 ( 
.A(n_812),
.Y(n_893)
);

INVx2_ASAP7_75t_L g894 ( 
.A(n_838),
.Y(n_894)
);

BUFx2_ASAP7_75t_L g895 ( 
.A(n_855),
.Y(n_895)
);

INVx1_ASAP7_75t_L g896 ( 
.A(n_823),
.Y(n_896)
);

INVx2_ASAP7_75t_L g897 ( 
.A(n_838),
.Y(n_897)
);

BUFx6f_ASAP7_75t_L g898 ( 
.A(n_812),
.Y(n_898)
);

INVx2_ASAP7_75t_L g899 ( 
.A(n_838),
.Y(n_899)
);

BUFx4f_ASAP7_75t_L g900 ( 
.A(n_812),
.Y(n_900)
);

AND2x2_ASAP7_75t_L g901 ( 
.A(n_840),
.B(n_843),
.Y(n_901)
);

INVx1_ASAP7_75t_L g902 ( 
.A(n_824),
.Y(n_902)
);

INVx2_ASAP7_75t_L g903 ( 
.A(n_819),
.Y(n_903)
);

BUFx2_ASAP7_75t_L g904 ( 
.A(n_812),
.Y(n_904)
);

AND2x2_ASAP7_75t_L g905 ( 
.A(n_847),
.B(n_814),
.Y(n_905)
);

BUFx6f_ASAP7_75t_L g906 ( 
.A(n_812),
.Y(n_906)
);

AND2x2_ASAP7_75t_L g907 ( 
.A(n_821),
.B(n_844),
.Y(n_907)
);

INVx1_ASAP7_75t_L g908 ( 
.A(n_833),
.Y(n_908)
);

BUFx2_ASAP7_75t_SL g909 ( 
.A(n_876),
.Y(n_909)
);

HB1xp67_ASAP7_75t_L g910 ( 
.A(n_859),
.Y(n_910)
);

INVx1_ASAP7_75t_L g911 ( 
.A(n_863),
.Y(n_911)
);

INVx3_ASAP7_75t_L g912 ( 
.A(n_867),
.Y(n_912)
);

INVx2_ASAP7_75t_L g913 ( 
.A(n_863),
.Y(n_913)
);

INVx2_ASAP7_75t_L g914 ( 
.A(n_863),
.Y(n_914)
);

INVx2_ASAP7_75t_L g915 ( 
.A(n_890),
.Y(n_915)
);

AND2x2_ASAP7_75t_L g916 ( 
.A(n_895),
.B(n_815),
.Y(n_916)
);

INVx1_ASAP7_75t_L g917 ( 
.A(n_903),
.Y(n_917)
);

AO21x2_ASAP7_75t_L g918 ( 
.A1(n_884),
.A2(n_825),
.B(n_826),
.Y(n_918)
);

NAND2xp5_ASAP7_75t_L g919 ( 
.A(n_903),
.B(n_818),
.Y(n_919)
);

INVx2_ASAP7_75t_L g920 ( 
.A(n_890),
.Y(n_920)
);

INVx1_ASAP7_75t_L g921 ( 
.A(n_903),
.Y(n_921)
);

AND2x2_ASAP7_75t_L g922 ( 
.A(n_895),
.B(n_811),
.Y(n_922)
);

INVx1_ASAP7_75t_L g923 ( 
.A(n_895),
.Y(n_923)
);

INVx3_ASAP7_75t_L g924 ( 
.A(n_867),
.Y(n_924)
);

HB1xp67_ASAP7_75t_L g925 ( 
.A(n_859),
.Y(n_925)
);

AO21x2_ASAP7_75t_L g926 ( 
.A1(n_884),
.A2(n_865),
.B(n_869),
.Y(n_926)
);

INVx1_ASAP7_75t_L g927 ( 
.A(n_870),
.Y(n_927)
);

INVx1_ASAP7_75t_L g928 ( 
.A(n_870),
.Y(n_928)
);

BUFx4f_ASAP7_75t_SL g929 ( 
.A(n_886),
.Y(n_929)
);

HB1xp67_ASAP7_75t_L g930 ( 
.A(n_859),
.Y(n_930)
);

NAND2xp5_ASAP7_75t_L g931 ( 
.A(n_884),
.B(n_852),
.Y(n_931)
);

INVx1_ASAP7_75t_L g932 ( 
.A(n_862),
.Y(n_932)
);

BUFx2_ASAP7_75t_L g933 ( 
.A(n_867),
.Y(n_933)
);

AO21x2_ASAP7_75t_L g934 ( 
.A1(n_865),
.A2(n_825),
.B(n_826),
.Y(n_934)
);

INVx2_ASAP7_75t_SL g935 ( 
.A(n_898),
.Y(n_935)
);

INVx1_ASAP7_75t_L g936 ( 
.A(n_862),
.Y(n_936)
);

AND2x2_ASAP7_75t_L g937 ( 
.A(n_867),
.B(n_811),
.Y(n_937)
);

NAND2xp5_ASAP7_75t_L g938 ( 
.A(n_907),
.B(n_852),
.Y(n_938)
);

OA21x2_ASAP7_75t_L g939 ( 
.A1(n_861),
.A2(n_851),
.B(n_822),
.Y(n_939)
);

AND2x2_ASAP7_75t_L g940 ( 
.A(n_937),
.B(n_867),
.Y(n_940)
);

OAI22xp33_ASAP7_75t_L g941 ( 
.A1(n_938),
.A2(n_900),
.B1(n_876),
.B2(n_883),
.Y(n_941)
);

INVx2_ASAP7_75t_L g942 ( 
.A(n_915),
.Y(n_942)
);

NOR2xp33_ASAP7_75t_L g943 ( 
.A(n_938),
.B(n_807),
.Y(n_943)
);

INVx2_ASAP7_75t_L g944 ( 
.A(n_915),
.Y(n_944)
);

INVx1_ASAP7_75t_L g945 ( 
.A(n_932),
.Y(n_945)
);

INVx1_ASAP7_75t_L g946 ( 
.A(n_932),
.Y(n_946)
);

OR2x2_ASAP7_75t_L g947 ( 
.A(n_923),
.B(n_905),
.Y(n_947)
);

AOI22xp33_ASAP7_75t_L g948 ( 
.A1(n_916),
.A2(n_856),
.B1(n_905),
.B2(n_907),
.Y(n_948)
);

AND2x2_ASAP7_75t_L g949 ( 
.A(n_937),
.B(n_905),
.Y(n_949)
);

BUFx6f_ASAP7_75t_L g950 ( 
.A(n_939),
.Y(n_950)
);

AND2x4_ASAP7_75t_L g951 ( 
.A(n_935),
.B(n_893),
.Y(n_951)
);

INVx1_ASAP7_75t_SL g952 ( 
.A(n_937),
.Y(n_952)
);

AND2x4_ASAP7_75t_L g953 ( 
.A(n_935),
.B(n_893),
.Y(n_953)
);

INVx1_ASAP7_75t_L g954 ( 
.A(n_932),
.Y(n_954)
);

INVx3_ASAP7_75t_L g955 ( 
.A(n_939),
.Y(n_955)
);

OR2x2_ASAP7_75t_L g956 ( 
.A(n_923),
.B(n_907),
.Y(n_956)
);

BUFx6f_ASAP7_75t_L g957 ( 
.A(n_939),
.Y(n_957)
);

NAND2xp5_ASAP7_75t_L g958 ( 
.A(n_936),
.B(n_882),
.Y(n_958)
);

INVx1_ASAP7_75t_L g959 ( 
.A(n_936),
.Y(n_959)
);

OR2x2_ASAP7_75t_L g960 ( 
.A(n_923),
.B(n_901),
.Y(n_960)
);

OAI221xp5_ASAP7_75t_SL g961 ( 
.A1(n_916),
.A2(n_856),
.B1(n_857),
.B2(n_868),
.C(n_904),
.Y(n_961)
);

BUFx2_ASAP7_75t_L g962 ( 
.A(n_939),
.Y(n_962)
);

AND2x4_ASAP7_75t_L g963 ( 
.A(n_935),
.B(n_893),
.Y(n_963)
);

INVx2_ASAP7_75t_SL g964 ( 
.A(n_910),
.Y(n_964)
);

AND2x2_ASAP7_75t_L g965 ( 
.A(n_933),
.B(n_866),
.Y(n_965)
);

AO21x2_ASAP7_75t_L g966 ( 
.A1(n_926),
.A2(n_865),
.B(n_869),
.Y(n_966)
);

BUFx2_ASAP7_75t_L g967 ( 
.A(n_939),
.Y(n_967)
);

NAND2xp5_ASAP7_75t_L g968 ( 
.A(n_936),
.B(n_888),
.Y(n_968)
);

INVx2_ASAP7_75t_L g969 ( 
.A(n_915),
.Y(n_969)
);

NAND2xp5_ASAP7_75t_L g970 ( 
.A(n_919),
.B(n_888),
.Y(n_970)
);

INVx2_ASAP7_75t_L g971 ( 
.A(n_915),
.Y(n_971)
);

AND2x2_ASAP7_75t_L g972 ( 
.A(n_933),
.B(n_866),
.Y(n_972)
);

INVxp67_ASAP7_75t_SL g973 ( 
.A(n_910),
.Y(n_973)
);

INVx1_ASAP7_75t_L g974 ( 
.A(n_927),
.Y(n_974)
);

INVx2_ASAP7_75t_L g975 ( 
.A(n_920),
.Y(n_975)
);

INVx3_ASAP7_75t_L g976 ( 
.A(n_939),
.Y(n_976)
);

INVx1_ASAP7_75t_L g977 ( 
.A(n_927),
.Y(n_977)
);

AND2x2_ASAP7_75t_L g978 ( 
.A(n_933),
.B(n_926),
.Y(n_978)
);

INVx1_ASAP7_75t_L g979 ( 
.A(n_928),
.Y(n_979)
);

AOI22xp5_ASAP7_75t_L g980 ( 
.A1(n_948),
.A2(n_916),
.B1(n_871),
.B2(n_931),
.Y(n_980)
);

AND2x2_ASAP7_75t_L g981 ( 
.A(n_949),
.B(n_922),
.Y(n_981)
);

NOR3xp33_ASAP7_75t_L g982 ( 
.A(n_961),
.B(n_931),
.C(n_860),
.Y(n_982)
);

NAND2xp5_ASAP7_75t_L g983 ( 
.A(n_949),
.B(n_922),
.Y(n_983)
);

NAND2xp5_ASAP7_75t_L g984 ( 
.A(n_949),
.B(n_922),
.Y(n_984)
);

INVx1_ASAP7_75t_L g985 ( 
.A(n_945),
.Y(n_985)
);

AND2x2_ASAP7_75t_L g986 ( 
.A(n_952),
.B(n_965),
.Y(n_986)
);

AND2x2_ASAP7_75t_L g987 ( 
.A(n_952),
.B(n_912),
.Y(n_987)
);

NAND2xp5_ASAP7_75t_L g988 ( 
.A(n_956),
.B(n_925),
.Y(n_988)
);

NAND2xp5_ASAP7_75t_L g989 ( 
.A(n_956),
.B(n_970),
.Y(n_989)
);

NAND2xp5_ASAP7_75t_L g990 ( 
.A(n_970),
.B(n_925),
.Y(n_990)
);

NAND2xp5_ASAP7_75t_L g991 ( 
.A(n_964),
.B(n_930),
.Y(n_991)
);

NAND2xp5_ASAP7_75t_L g992 ( 
.A(n_964),
.B(n_930),
.Y(n_992)
);

AOI221xp5_ASAP7_75t_L g993 ( 
.A1(n_961),
.A2(n_926),
.B1(n_919),
.B2(n_902),
.C(n_896),
.Y(n_993)
);

AND2x2_ASAP7_75t_SL g994 ( 
.A(n_962),
.B(n_967),
.Y(n_994)
);

OAI221xp5_ASAP7_75t_L g995 ( 
.A1(n_962),
.A2(n_967),
.B1(n_943),
.B2(n_950),
.C(n_957),
.Y(n_995)
);

NAND2xp5_ASAP7_75t_L g996 ( 
.A(n_964),
.B(n_928),
.Y(n_996)
);

NAND3xp33_ASAP7_75t_L g997 ( 
.A(n_978),
.B(n_868),
.C(n_902),
.Y(n_997)
);

NAND2xp5_ASAP7_75t_L g998 ( 
.A(n_960),
.B(n_857),
.Y(n_998)
);

NAND2xp5_ASAP7_75t_L g999 ( 
.A(n_960),
.B(n_857),
.Y(n_999)
);

AND2x2_ASAP7_75t_L g1000 ( 
.A(n_965),
.B(n_924),
.Y(n_1000)
);

NAND2xp5_ASAP7_75t_L g1001 ( 
.A(n_947),
.B(n_901),
.Y(n_1001)
);

OAI221xp5_ASAP7_75t_L g1002 ( 
.A1(n_950),
.A2(n_957),
.B1(n_882),
.B2(n_896),
.C(n_908),
.Y(n_1002)
);

AND2x2_ASAP7_75t_L g1003 ( 
.A(n_965),
.B(n_924),
.Y(n_1003)
);

NAND2xp5_ASAP7_75t_L g1004 ( 
.A(n_947),
.B(n_901),
.Y(n_1004)
);

INVx3_ASAP7_75t_L g1005 ( 
.A(n_994),
.Y(n_1005)
);

INVx1_ASAP7_75t_L g1006 ( 
.A(n_985),
.Y(n_1006)
);

INVx3_ASAP7_75t_L g1007 ( 
.A(n_994),
.Y(n_1007)
);

INVx2_ASAP7_75t_L g1008 ( 
.A(n_981),
.Y(n_1008)
);

AND2x4_ASAP7_75t_L g1009 ( 
.A(n_1000),
.B(n_978),
.Y(n_1009)
);

NAND2xp5_ASAP7_75t_L g1010 ( 
.A(n_990),
.B(n_978),
.Y(n_1010)
);

AND2x2_ASAP7_75t_L g1011 ( 
.A(n_981),
.B(n_972),
.Y(n_1011)
);

AND2x2_ASAP7_75t_L g1012 ( 
.A(n_986),
.B(n_972),
.Y(n_1012)
);

BUFx2_ASAP7_75t_L g1013 ( 
.A(n_991),
.Y(n_1013)
);

INVx1_ASAP7_75t_SL g1014 ( 
.A(n_992),
.Y(n_1014)
);

INVx1_ASAP7_75t_L g1015 ( 
.A(n_996),
.Y(n_1015)
);

INVx2_ASAP7_75t_L g1016 ( 
.A(n_1002),
.Y(n_1016)
);

INVx2_ASAP7_75t_L g1017 ( 
.A(n_987),
.Y(n_1017)
);

AND2x2_ASAP7_75t_L g1018 ( 
.A(n_986),
.B(n_972),
.Y(n_1018)
);

INVx1_ASAP7_75t_L g1019 ( 
.A(n_988),
.Y(n_1019)
);

INVx1_ASAP7_75t_L g1020 ( 
.A(n_989),
.Y(n_1020)
);

INVx2_ASAP7_75t_L g1021 ( 
.A(n_987),
.Y(n_1021)
);

INVx1_ASAP7_75t_L g1022 ( 
.A(n_1001),
.Y(n_1022)
);

AND2x2_ASAP7_75t_L g1023 ( 
.A(n_1000),
.B(n_950),
.Y(n_1023)
);

INVx2_ASAP7_75t_L g1024 ( 
.A(n_997),
.Y(n_1024)
);

AND2x2_ASAP7_75t_L g1025 ( 
.A(n_1003),
.B(n_950),
.Y(n_1025)
);

AND2x2_ASAP7_75t_L g1026 ( 
.A(n_1011),
.B(n_1005),
.Y(n_1026)
);

INVx1_ASAP7_75t_L g1027 ( 
.A(n_1006),
.Y(n_1027)
);

INVx1_ASAP7_75t_L g1028 ( 
.A(n_1006),
.Y(n_1028)
);

OR2x2_ASAP7_75t_L g1029 ( 
.A(n_1020),
.B(n_983),
.Y(n_1029)
);

INVx1_ASAP7_75t_L g1030 ( 
.A(n_1015),
.Y(n_1030)
);

INVx1_ASAP7_75t_L g1031 ( 
.A(n_1015),
.Y(n_1031)
);

AND2x2_ASAP7_75t_L g1032 ( 
.A(n_1011),
.B(n_1005),
.Y(n_1032)
);

INVx1_ASAP7_75t_L g1033 ( 
.A(n_1019),
.Y(n_1033)
);

OR2x2_ASAP7_75t_L g1034 ( 
.A(n_1020),
.B(n_984),
.Y(n_1034)
);

NAND2x1_ASAP7_75t_L g1035 ( 
.A(n_1005),
.B(n_1003),
.Y(n_1035)
);

NOR2x1_ASAP7_75t_L g1036 ( 
.A(n_1005),
.B(n_1007),
.Y(n_1036)
);

AND2x2_ASAP7_75t_L g1037 ( 
.A(n_1026),
.B(n_1005),
.Y(n_1037)
);

NOR2xp33_ASAP7_75t_SL g1038 ( 
.A(n_1036),
.B(n_1024),
.Y(n_1038)
);

AND2x2_ASAP7_75t_L g1039 ( 
.A(n_1026),
.B(n_1032),
.Y(n_1039)
);

INVx1_ASAP7_75t_L g1040 ( 
.A(n_1027),
.Y(n_1040)
);

AND2x2_ASAP7_75t_L g1041 ( 
.A(n_1032),
.B(n_1007),
.Y(n_1041)
);

INVx1_ASAP7_75t_L g1042 ( 
.A(n_1028),
.Y(n_1042)
);

OR2x2_ASAP7_75t_L g1043 ( 
.A(n_1033),
.B(n_1016),
.Y(n_1043)
);

INVx1_ASAP7_75t_L g1044 ( 
.A(n_1040),
.Y(n_1044)
);

NAND2xp5_ASAP7_75t_SL g1045 ( 
.A(n_1038),
.B(n_1007),
.Y(n_1045)
);

INVxp67_ASAP7_75t_L g1046 ( 
.A(n_1043),
.Y(n_1046)
);

INVx1_ASAP7_75t_L g1047 ( 
.A(n_1042),
.Y(n_1047)
);

INVx1_ASAP7_75t_L g1048 ( 
.A(n_1044),
.Y(n_1048)
);

NAND2xp5_ASAP7_75t_SL g1049 ( 
.A(n_1045),
.B(n_1007),
.Y(n_1049)
);

AOI32xp33_ASAP7_75t_L g1050 ( 
.A1(n_1044),
.A2(n_1024),
.A3(n_1016),
.B1(n_1043),
.B2(n_982),
.Y(n_1050)
);

INVx2_ASAP7_75t_L g1051 ( 
.A(n_1047),
.Y(n_1051)
);

INVxp67_ASAP7_75t_L g1052 ( 
.A(n_1046),
.Y(n_1052)
);

AND2x2_ASAP7_75t_L g1053 ( 
.A(n_1045),
.B(n_1039),
.Y(n_1053)
);

INVx2_ASAP7_75t_SL g1054 ( 
.A(n_1045),
.Y(n_1054)
);

INVx1_ASAP7_75t_L g1055 ( 
.A(n_1044),
.Y(n_1055)
);

AOI22xp33_ASAP7_75t_SL g1056 ( 
.A1(n_1046),
.A2(n_1024),
.B1(n_1016),
.B2(n_1037),
.Y(n_1056)
);

OAI21xp33_ASAP7_75t_L g1057 ( 
.A1(n_1045),
.A2(n_1039),
.B(n_1037),
.Y(n_1057)
);

OAI22xp5_ASAP7_75t_L g1058 ( 
.A1(n_1045),
.A2(n_995),
.B1(n_1035),
.B2(n_1041),
.Y(n_1058)
);

NAND2xp5_ASAP7_75t_L g1059 ( 
.A(n_1056),
.B(n_1030),
.Y(n_1059)
);

NAND2xp5_ASAP7_75t_L g1060 ( 
.A(n_1051),
.B(n_1031),
.Y(n_1060)
);

INVx1_ASAP7_75t_L g1061 ( 
.A(n_1048),
.Y(n_1061)
);

NOR2xp33_ASAP7_75t_L g1062 ( 
.A(n_1052),
.B(n_1054),
.Y(n_1062)
);

NAND2xp5_ASAP7_75t_L g1063 ( 
.A(n_1050),
.B(n_1041),
.Y(n_1063)
);

AOI22xp33_ASAP7_75t_L g1064 ( 
.A1(n_1055),
.A2(n_993),
.B1(n_926),
.B2(n_966),
.Y(n_1064)
);

INVx1_ASAP7_75t_L g1065 ( 
.A(n_1053),
.Y(n_1065)
);

NOR2xp33_ASAP7_75t_L g1066 ( 
.A(n_1057),
.B(n_860),
.Y(n_1066)
);

NAND2xp5_ASAP7_75t_L g1067 ( 
.A(n_1057),
.B(n_1013),
.Y(n_1067)
);

NOR2xp33_ASAP7_75t_L g1068 ( 
.A(n_1049),
.B(n_1014),
.Y(n_1068)
);

INVx1_ASAP7_75t_L g1069 ( 
.A(n_1058),
.Y(n_1069)
);

NOR2xp33_ASAP7_75t_L g1070 ( 
.A(n_1052),
.B(n_1014),
.Y(n_1070)
);

INVx1_ASAP7_75t_L g1071 ( 
.A(n_1048),
.Y(n_1071)
);

OR2x2_ASAP7_75t_L g1072 ( 
.A(n_1052),
.B(n_1029),
.Y(n_1072)
);

NAND2xp5_ASAP7_75t_SL g1073 ( 
.A(n_1054),
.B(n_1013),
.Y(n_1073)
);

NAND2xp5_ASAP7_75t_L g1074 ( 
.A(n_1056),
.B(n_1009),
.Y(n_1074)
);

OAI22x1_ASAP7_75t_L g1075 ( 
.A1(n_1054),
.A2(n_834),
.B1(n_1009),
.B2(n_980),
.Y(n_1075)
);

AOI211xp5_ASAP7_75t_L g1076 ( 
.A1(n_1063),
.A2(n_950),
.B(n_957),
.C(n_834),
.Y(n_1076)
);

AOI211xp5_ASAP7_75t_L g1077 ( 
.A1(n_1059),
.A2(n_957),
.B(n_950),
.C(n_976),
.Y(n_1077)
);

AOI22xp5_ASAP7_75t_L g1078 ( 
.A1(n_1064),
.A2(n_926),
.B1(n_966),
.B2(n_950),
.Y(n_1078)
);

AOI222xp33_ASAP7_75t_L g1079 ( 
.A1(n_1064),
.A2(n_957),
.B1(n_1010),
.B2(n_976),
.C1(n_955),
.C2(n_908),
.Y(n_1079)
);

AOI21xp33_ASAP7_75t_L g1080 ( 
.A1(n_1069),
.A2(n_1061),
.B(n_1071),
.Y(n_1080)
);

NOR2xp33_ASAP7_75t_L g1081 ( 
.A(n_1062),
.B(n_1073),
.Y(n_1081)
);

OR2x2_ASAP7_75t_L g1082 ( 
.A(n_1072),
.B(n_1034),
.Y(n_1082)
);

NAND2xp5_ASAP7_75t_SL g1083 ( 
.A(n_1066),
.B(n_1009),
.Y(n_1083)
);

OAI211xp5_ASAP7_75t_L g1084 ( 
.A1(n_1065),
.A2(n_976),
.B(n_955),
.C(n_1025),
.Y(n_1084)
);

NAND4xp25_ASAP7_75t_L g1085 ( 
.A(n_1070),
.B(n_1067),
.C(n_1068),
.D(n_1074),
.Y(n_1085)
);

NAND4xp25_ASAP7_75t_L g1086 ( 
.A(n_1060),
.B(n_1009),
.C(n_1025),
.D(n_1023),
.Y(n_1086)
);

OAI21xp33_ASAP7_75t_L g1087 ( 
.A1(n_1075),
.A2(n_1019),
.B(n_1010),
.Y(n_1087)
);

NAND2xp5_ASAP7_75t_L g1088 ( 
.A(n_1065),
.B(n_1009),
.Y(n_1088)
);

AOI22xp5_ASAP7_75t_L g1089 ( 
.A1(n_1064),
.A2(n_966),
.B1(n_957),
.B2(n_976),
.Y(n_1089)
);

AOI221xp5_ASAP7_75t_L g1090 ( 
.A1(n_1064),
.A2(n_966),
.B1(n_957),
.B2(n_955),
.C(n_918),
.Y(n_1090)
);

AOI221xp5_ASAP7_75t_L g1091 ( 
.A1(n_1064),
.A2(n_955),
.B1(n_918),
.B2(n_1022),
.C(n_934),
.Y(n_1091)
);

OAI221xp5_ASAP7_75t_SL g1092 ( 
.A1(n_1063),
.A2(n_941),
.B1(n_1004),
.B2(n_1022),
.C(n_1008),
.Y(n_1092)
);

OAI21xp5_ASAP7_75t_L g1093 ( 
.A1(n_1064),
.A2(n_1025),
.B(n_1023),
.Y(n_1093)
);

NOR3x1_ASAP7_75t_L g1094 ( 
.A(n_1069),
.B(n_887),
.C(n_998),
.Y(n_1094)
);

AOI22xp5_ASAP7_75t_L g1095 ( 
.A1(n_1078),
.A2(n_918),
.B1(n_871),
.B2(n_1023),
.Y(n_1095)
);

NOR3x1_ASAP7_75t_L g1096 ( 
.A(n_1085),
.B(n_887),
.C(n_858),
.Y(n_1096)
);

NAND2xp5_ASAP7_75t_L g1097 ( 
.A(n_1082),
.B(n_1080),
.Y(n_1097)
);

AOI22xp33_ASAP7_75t_L g1098 ( 
.A1(n_1090),
.A2(n_906),
.B1(n_898),
.B2(n_918),
.Y(n_1098)
);

NOR2x1_ASAP7_75t_L g1099 ( 
.A(n_1081),
.B(n_1008),
.Y(n_1099)
);

AOI211x1_ASAP7_75t_L g1100 ( 
.A1(n_1083),
.A2(n_1018),
.B(n_1012),
.C(n_1011),
.Y(n_1100)
);

NOR4xp25_ASAP7_75t_L g1101 ( 
.A(n_1092),
.B(n_1008),
.C(n_1017),
.D(n_1021),
.Y(n_1101)
);

NOR4xp75_ASAP7_75t_L g1102 ( 
.A(n_1088),
.B(n_1018),
.C(n_1012),
.D(n_999),
.Y(n_1102)
);

NAND2xp5_ASAP7_75t_L g1103 ( 
.A(n_1094),
.B(n_1017),
.Y(n_1103)
);

NOR3xp33_ASAP7_75t_L g1104 ( 
.A(n_1076),
.B(n_941),
.C(n_851),
.Y(n_1104)
);

NAND4xp25_ASAP7_75t_SL g1105 ( 
.A(n_1077),
.B(n_1084),
.C(n_1079),
.D(n_1091),
.Y(n_1105)
);

INVx1_ASAP7_75t_L g1106 ( 
.A(n_1087),
.Y(n_1106)
);

AOI21xp5_ASAP7_75t_L g1107 ( 
.A1(n_1089),
.A2(n_1021),
.B(n_1017),
.Y(n_1107)
);

NAND2xp5_ASAP7_75t_SL g1108 ( 
.A(n_1093),
.B(n_929),
.Y(n_1108)
);

NOR3xp33_ASAP7_75t_L g1109 ( 
.A(n_1086),
.B(n_968),
.C(n_958),
.Y(n_1109)
);

OR2x2_ASAP7_75t_L g1110 ( 
.A(n_1082),
.B(n_1012),
.Y(n_1110)
);

NAND5xp2_ASAP7_75t_L g1111 ( 
.A(n_1081),
.B(n_1018),
.C(n_858),
.D(n_929),
.E(n_886),
.Y(n_1111)
);

NAND3xp33_ASAP7_75t_L g1112 ( 
.A(n_1097),
.B(n_858),
.C(n_886),
.Y(n_1112)
);

AOI211xp5_ASAP7_75t_L g1113 ( 
.A1(n_1106),
.A2(n_1021),
.B(n_958),
.C(n_968),
.Y(n_1113)
);

NOR2xp33_ASAP7_75t_L g1114 ( 
.A(n_1111),
.B(n_858),
.Y(n_1114)
);

NOR3xp33_ASAP7_75t_L g1115 ( 
.A(n_1103),
.B(n_883),
.C(n_828),
.Y(n_1115)
);

AOI211xp5_ASAP7_75t_SL g1116 ( 
.A1(n_1110),
.A2(n_1104),
.B(n_1095),
.C(n_1096),
.Y(n_1116)
);

O2A1O1Ixp33_ASAP7_75t_L g1117 ( 
.A1(n_1101),
.A2(n_918),
.B(n_934),
.C(n_973),
.Y(n_1117)
);

NAND4xp75_ASAP7_75t_L g1118 ( 
.A(n_1099),
.B(n_858),
.C(n_886),
.D(n_946),
.Y(n_1118)
);

NAND4xp25_ASAP7_75t_L g1119 ( 
.A(n_1100),
.B(n_946),
.C(n_945),
.D(n_954),
.Y(n_1119)
);

O2A1O1Ixp33_ASAP7_75t_L g1120 ( 
.A1(n_1108),
.A2(n_934),
.B(n_973),
.C(n_864),
.Y(n_1120)
);

NAND2xp5_ASAP7_75t_SL g1121 ( 
.A(n_1098),
.B(n_886),
.Y(n_1121)
);

A2O1A1Ixp33_ASAP7_75t_L g1122 ( 
.A1(n_1107),
.A2(n_900),
.B(n_893),
.C(n_979),
.Y(n_1122)
);

OAI211xp5_ASAP7_75t_L g1123 ( 
.A1(n_1109),
.A2(n_954),
.B(n_959),
.C(n_979),
.Y(n_1123)
);

NAND3xp33_ASAP7_75t_SL g1124 ( 
.A(n_1102),
.B(n_883),
.C(n_904),
.Y(n_1124)
);

OAI221xp5_ASAP7_75t_SL g1125 ( 
.A1(n_1105),
.A2(n_904),
.B1(n_974),
.B2(n_977),
.C(n_959),
.Y(n_1125)
);

OAI211xp5_ASAP7_75t_L g1126 ( 
.A1(n_1097),
.A2(n_977),
.B(n_974),
.C(n_876),
.Y(n_1126)
);

NAND3xp33_ASAP7_75t_SL g1127 ( 
.A(n_1097),
.B(n_892),
.C(n_940),
.Y(n_1127)
);

NOR4xp25_ASAP7_75t_L g1128 ( 
.A(n_1097),
.B(n_880),
.C(n_877),
.D(n_822),
.Y(n_1128)
);

NAND2xp5_ASAP7_75t_SL g1129 ( 
.A(n_1097),
.B(n_876),
.Y(n_1129)
);

OAI211xp5_ASAP7_75t_SL g1130 ( 
.A1(n_1097),
.A2(n_924),
.B(n_912),
.C(n_934),
.Y(n_1130)
);

NAND4xp25_ASAP7_75t_L g1131 ( 
.A(n_1097),
.B(n_940),
.C(n_912),
.D(n_924),
.Y(n_1131)
);

NAND4xp25_ASAP7_75t_SL g1132 ( 
.A(n_1097),
.B(n_940),
.C(n_866),
.D(n_934),
.Y(n_1132)
);

AOI211x1_ASAP7_75t_SL g1133 ( 
.A1(n_1097),
.A2(n_897),
.B(n_894),
.C(n_899),
.Y(n_1133)
);

AOI22xp5_ASAP7_75t_L g1134 ( 
.A1(n_1097),
.A2(n_876),
.B1(n_906),
.B2(n_898),
.Y(n_1134)
);

NAND2xp5_ASAP7_75t_L g1135 ( 
.A(n_1097),
.B(n_912),
.Y(n_1135)
);

AOI22xp5_ASAP7_75t_L g1136 ( 
.A1(n_1115),
.A2(n_876),
.B1(n_906),
.B2(n_898),
.Y(n_1136)
);

INVx2_ASAP7_75t_L g1137 ( 
.A(n_1118),
.Y(n_1137)
);

INVx1_ASAP7_75t_L g1138 ( 
.A(n_1133),
.Y(n_1138)
);

INVx1_ASAP7_75t_L g1139 ( 
.A(n_1135),
.Y(n_1139)
);

INVx1_ASAP7_75t_L g1140 ( 
.A(n_1117),
.Y(n_1140)
);

OAI22xp33_ASAP7_75t_SL g1141 ( 
.A1(n_1125),
.A2(n_1129),
.B1(n_1121),
.B2(n_1114),
.Y(n_1141)
);

INVx1_ASAP7_75t_L g1142 ( 
.A(n_1113),
.Y(n_1142)
);

NOR2x1_ASAP7_75t_L g1143 ( 
.A(n_1112),
.B(n_909),
.Y(n_1143)
);

AOI22xp5_ASAP7_75t_L g1144 ( 
.A1(n_1127),
.A2(n_876),
.B1(n_906),
.B2(n_898),
.Y(n_1144)
);

NOR2xp67_ASAP7_75t_L g1145 ( 
.A(n_1132),
.B(n_912),
.Y(n_1145)
);

NOR2xp33_ASAP7_75t_SL g1146 ( 
.A(n_1124),
.B(n_889),
.Y(n_1146)
);

AOI22xp5_ASAP7_75t_L g1147 ( 
.A1(n_1134),
.A2(n_906),
.B1(n_898),
.B2(n_900),
.Y(n_1147)
);

INVx1_ASAP7_75t_L g1148 ( 
.A(n_1123),
.Y(n_1148)
);

NAND2xp5_ASAP7_75t_L g1149 ( 
.A(n_1128),
.B(n_1116),
.Y(n_1149)
);

NOR2x2_ASAP7_75t_L g1150 ( 
.A(n_1131),
.B(n_909),
.Y(n_1150)
);

INVx3_ASAP7_75t_L g1151 ( 
.A(n_1126),
.Y(n_1151)
);

INVx1_ASAP7_75t_L g1152 ( 
.A(n_1119),
.Y(n_1152)
);

INVx1_ASAP7_75t_SL g1153 ( 
.A(n_1130),
.Y(n_1153)
);

NAND2xp5_ASAP7_75t_L g1154 ( 
.A(n_1122),
.B(n_924),
.Y(n_1154)
);

INVx1_ASAP7_75t_L g1155 ( 
.A(n_1120),
.Y(n_1155)
);

NAND2xp5_ASAP7_75t_SL g1156 ( 
.A(n_1117),
.B(n_900),
.Y(n_1156)
);

NAND2xp5_ASAP7_75t_SL g1157 ( 
.A(n_1117),
.B(n_900),
.Y(n_1157)
);

HB1xp67_ASAP7_75t_L g1158 ( 
.A(n_1129),
.Y(n_1158)
);

AOI22xp5_ASAP7_75t_L g1159 ( 
.A1(n_1115),
.A2(n_906),
.B1(n_898),
.B2(n_953),
.Y(n_1159)
);

AO22x2_ASAP7_75t_L g1160 ( 
.A1(n_1140),
.A2(n_828),
.B1(n_909),
.B2(n_872),
.Y(n_1160)
);

OA222x2_ASAP7_75t_SL g1161 ( 
.A1(n_1152),
.A2(n_963),
.B1(n_953),
.B2(n_951),
.C1(n_911),
.C2(n_892),
.Y(n_1161)
);

INVx1_ASAP7_75t_L g1162 ( 
.A(n_1149),
.Y(n_1162)
);

INVx1_ASAP7_75t_SL g1163 ( 
.A(n_1158),
.Y(n_1163)
);

INVx1_ASAP7_75t_L g1164 ( 
.A(n_1138),
.Y(n_1164)
);

INVx1_ASAP7_75t_L g1165 ( 
.A(n_1142),
.Y(n_1165)
);

NAND4xp75_ASAP7_75t_L g1166 ( 
.A(n_1155),
.B(n_864),
.C(n_891),
.D(n_911),
.Y(n_1166)
);

NOR3xp33_ASAP7_75t_L g1167 ( 
.A(n_1137),
.B(n_921),
.C(n_917),
.Y(n_1167)
);

NOR3xp33_ASAP7_75t_L g1168 ( 
.A(n_1141),
.B(n_921),
.C(n_917),
.Y(n_1168)
);

OR2x2_ASAP7_75t_L g1169 ( 
.A(n_1148),
.B(n_1151),
.Y(n_1169)
);

NOR3xp33_ASAP7_75t_L g1170 ( 
.A(n_1151),
.B(n_921),
.C(n_917),
.Y(n_1170)
);

INVx2_ASAP7_75t_SL g1171 ( 
.A(n_1139),
.Y(n_1171)
);

NAND2xp5_ASAP7_75t_L g1172 ( 
.A(n_1153),
.B(n_911),
.Y(n_1172)
);

INVx1_ASAP7_75t_L g1173 ( 
.A(n_1156),
.Y(n_1173)
);

INVx1_ASAP7_75t_L g1174 ( 
.A(n_1157),
.Y(n_1174)
);

INVxp33_ASAP7_75t_L g1175 ( 
.A(n_1143),
.Y(n_1175)
);

INVx3_ASAP7_75t_SL g1176 ( 
.A(n_1150),
.Y(n_1176)
);

NOR2x1_ASAP7_75t_L g1177 ( 
.A(n_1145),
.B(n_1154),
.Y(n_1177)
);

AND2x4_ASAP7_75t_L g1178 ( 
.A(n_1159),
.B(n_963),
.Y(n_1178)
);

NAND4xp75_ASAP7_75t_L g1179 ( 
.A(n_1144),
.B(n_864),
.C(n_891),
.D(n_877),
.Y(n_1179)
);

OAI322xp33_ASAP7_75t_L g1180 ( 
.A1(n_1146),
.A2(n_880),
.A3(n_892),
.B1(n_873),
.B2(n_872),
.C1(n_913),
.C2(n_914),
.Y(n_1180)
);

NAND2xp5_ASAP7_75t_L g1181 ( 
.A(n_1136),
.B(n_1147),
.Y(n_1181)
);

NAND2xp5_ASAP7_75t_SL g1182 ( 
.A(n_1163),
.B(n_963),
.Y(n_1182)
);

INVx1_ASAP7_75t_L g1183 ( 
.A(n_1169),
.Y(n_1183)
);

INVx1_ASAP7_75t_L g1184 ( 
.A(n_1171),
.Y(n_1184)
);

HB1xp67_ASAP7_75t_L g1185 ( 
.A(n_1165),
.Y(n_1185)
);

AND2x2_ASAP7_75t_SL g1186 ( 
.A(n_1162),
.B(n_963),
.Y(n_1186)
);

AOI22xp5_ASAP7_75t_L g1187 ( 
.A1(n_1164),
.A2(n_906),
.B1(n_953),
.B2(n_951),
.Y(n_1187)
);

XNOR2x1_ASAP7_75t_L g1188 ( 
.A(n_1173),
.B(n_951),
.Y(n_1188)
);

XOR2xp5_ASAP7_75t_L g1189 ( 
.A(n_1174),
.B(n_953),
.Y(n_1189)
);

XNOR2x1_ASAP7_75t_L g1190 ( 
.A(n_1177),
.B(n_951),
.Y(n_1190)
);

INVx2_ASAP7_75t_SL g1191 ( 
.A(n_1176),
.Y(n_1191)
);

XNOR2xp5_ASAP7_75t_L g1192 ( 
.A(n_1175),
.B(n_892),
.Y(n_1192)
);

INVx1_ASAP7_75t_L g1193 ( 
.A(n_1160),
.Y(n_1193)
);

NOR2x1p5_ASAP7_75t_L g1194 ( 
.A(n_1181),
.B(n_889),
.Y(n_1194)
);

OR2x2_ASAP7_75t_L g1195 ( 
.A(n_1168),
.B(n_861),
.Y(n_1195)
);

AND2x4_ASAP7_75t_L g1196 ( 
.A(n_1170),
.B(n_861),
.Y(n_1196)
);

AOI22xp5_ASAP7_75t_L g1197 ( 
.A1(n_1185),
.A2(n_1183),
.B1(n_1191),
.B2(n_1186),
.Y(n_1197)
);

INVx2_ASAP7_75t_L g1198 ( 
.A(n_1190),
.Y(n_1198)
);

INVx1_ASAP7_75t_L g1199 ( 
.A(n_1184),
.Y(n_1199)
);

INVx1_ASAP7_75t_L g1200 ( 
.A(n_1193),
.Y(n_1200)
);

INVx1_ASAP7_75t_L g1201 ( 
.A(n_1182),
.Y(n_1201)
);

XNOR2x1_ASAP7_75t_L g1202 ( 
.A(n_1194),
.B(n_1160),
.Y(n_1202)
);

INVx1_ASAP7_75t_L g1203 ( 
.A(n_1189),
.Y(n_1203)
);

INVx1_ASAP7_75t_L g1204 ( 
.A(n_1188),
.Y(n_1204)
);

AOI22xp5_ASAP7_75t_L g1205 ( 
.A1(n_1192),
.A2(n_1166),
.B1(n_1172),
.B2(n_1167),
.Y(n_1205)
);

INVx1_ASAP7_75t_L g1206 ( 
.A(n_1196),
.Y(n_1206)
);

OAI22xp5_ASAP7_75t_L g1207 ( 
.A1(n_1187),
.A2(n_1179),
.B1(n_1178),
.B2(n_1161),
.Y(n_1207)
);

INVx1_ASAP7_75t_L g1208 ( 
.A(n_1196),
.Y(n_1208)
);

INVx1_ASAP7_75t_L g1209 ( 
.A(n_1195),
.Y(n_1209)
);

AOI22x1_ASAP7_75t_L g1210 ( 
.A1(n_1183),
.A2(n_1178),
.B1(n_1180),
.B2(n_889),
.Y(n_1210)
);

AOI22xp5_ASAP7_75t_L g1211 ( 
.A1(n_1185),
.A2(n_864),
.B1(n_873),
.B2(n_971),
.Y(n_1211)
);

OAI211xp5_ASAP7_75t_SL g1212 ( 
.A1(n_1197),
.A2(n_1199),
.B(n_1204),
.C(n_1200),
.Y(n_1212)
);

OAI22xp5_ASAP7_75t_L g1213 ( 
.A1(n_1201),
.A2(n_864),
.B1(n_975),
.B2(n_971),
.Y(n_1213)
);

OAI22xp5_ASAP7_75t_L g1214 ( 
.A1(n_1206),
.A2(n_975),
.B1(n_971),
.B2(n_969),
.Y(n_1214)
);

NOR3xp33_ASAP7_75t_L g1215 ( 
.A(n_1203),
.B(n_874),
.C(n_897),
.Y(n_1215)
);

NOR4xp25_ASAP7_75t_L g1216 ( 
.A(n_1198),
.B(n_1209),
.C(n_1208),
.D(n_1207),
.Y(n_1216)
);

OAI221xp5_ASAP7_75t_L g1217 ( 
.A1(n_1210),
.A2(n_975),
.B1(n_969),
.B2(n_944),
.C(n_942),
.Y(n_1217)
);

NOR2xp33_ASAP7_75t_L g1218 ( 
.A(n_1202),
.B(n_969),
.Y(n_1218)
);

NAND3xp33_ASAP7_75t_SL g1219 ( 
.A(n_1205),
.B(n_874),
.C(n_944),
.Y(n_1219)
);

AOI22xp5_ASAP7_75t_L g1220 ( 
.A1(n_1211),
.A2(n_942),
.B1(n_944),
.B2(n_874),
.Y(n_1220)
);

INVx1_ASAP7_75t_L g1221 ( 
.A(n_1197),
.Y(n_1221)
);

OAI21xp5_ASAP7_75t_SL g1222 ( 
.A1(n_1212),
.A2(n_878),
.B(n_875),
.Y(n_1222)
);

OAI22xp5_ASAP7_75t_L g1223 ( 
.A1(n_1221),
.A2(n_942),
.B1(n_899),
.B2(n_897),
.Y(n_1223)
);

NOR2xp33_ASAP7_75t_L g1224 ( 
.A(n_1218),
.B(n_899),
.Y(n_1224)
);

INVx1_ASAP7_75t_L g1225 ( 
.A(n_1219),
.Y(n_1225)
);

AOI22xp5_ASAP7_75t_L g1226 ( 
.A1(n_1216),
.A2(n_1215),
.B1(n_1213),
.B2(n_1217),
.Y(n_1226)
);

NAND2xp5_ASAP7_75t_L g1227 ( 
.A(n_1214),
.B(n_913),
.Y(n_1227)
);

AOI22xp5_ASAP7_75t_L g1228 ( 
.A1(n_1226),
.A2(n_1220),
.B1(n_894),
.B2(n_875),
.Y(n_1228)
);

OAI21xp5_ASAP7_75t_L g1229 ( 
.A1(n_1225),
.A2(n_885),
.B(n_914),
.Y(n_1229)
);

OR2x2_ASAP7_75t_L g1230 ( 
.A(n_1222),
.B(n_875),
.Y(n_1230)
);

AOI22xp5_ASAP7_75t_L g1231 ( 
.A1(n_1224),
.A2(n_894),
.B1(n_875),
.B2(n_891),
.Y(n_1231)
);

AOI21xp5_ASAP7_75t_SL g1232 ( 
.A1(n_1228),
.A2(n_1230),
.B(n_1229),
.Y(n_1232)
);

NAND2xp5_ASAP7_75t_L g1233 ( 
.A(n_1232),
.B(n_1231),
.Y(n_1233)
);

AOI322xp5_ASAP7_75t_L g1234 ( 
.A1(n_1233),
.A2(n_1227),
.A3(n_1223),
.B1(n_878),
.B2(n_914),
.C1(n_913),
.C2(n_920),
.Y(n_1234)
);

AOI221xp5_ASAP7_75t_L g1235 ( 
.A1(n_1234),
.A2(n_914),
.B1(n_913),
.B2(n_875),
.C(n_879),
.Y(n_1235)
);

AOI211xp5_ASAP7_75t_L g1236 ( 
.A1(n_1235),
.A2(n_879),
.B(n_885),
.C(n_881),
.Y(n_1236)
);


endmodule