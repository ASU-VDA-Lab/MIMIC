module fake_jpeg_20756_n_136 (n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_136);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_136;

wire n_117;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_73;
wire n_14;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_31;
wire n_29;
wire n_103;
wire n_50;
wire n_15;
wire n_124;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_30;
wire n_106;
wire n_111;
wire n_24;
wire n_44;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_20;
wire n_18;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_22;
wire n_101;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_97;
wire n_135;
wire n_36;
wire n_62;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_96;

NOR2xp33_ASAP7_75t_L g13 ( 
.A(n_0),
.B(n_5),
.Y(n_13)
);

BUFx3_ASAP7_75t_L g14 ( 
.A(n_12),
.Y(n_14)
);

INVx13_ASAP7_75t_L g15 ( 
.A(n_0),
.Y(n_15)
);

BUFx16f_ASAP7_75t_L g16 ( 
.A(n_0),
.Y(n_16)
);

BUFx3_ASAP7_75t_L g17 ( 
.A(n_1),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_12),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_11),
.Y(n_19)
);

INVx2_ASAP7_75t_L g20 ( 
.A(n_5),
.Y(n_20)
);

BUFx3_ASAP7_75t_L g21 ( 
.A(n_3),
.Y(n_21)
);

BUFx3_ASAP7_75t_L g22 ( 
.A(n_3),
.Y(n_22)
);

AND2x2_ASAP7_75t_L g23 ( 
.A(n_2),
.B(n_9),
.Y(n_23)
);

INVx2_ASAP7_75t_L g24 ( 
.A(n_6),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_11),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_4),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_3),
.Y(n_27)
);

BUFx2_ASAP7_75t_L g28 ( 
.A(n_15),
.Y(n_28)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_28),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_26),
.Y(n_29)
);

NOR2xp33_ASAP7_75t_L g45 ( 
.A(n_29),
.B(n_30),
.Y(n_45)
);

OR2x4_ASAP7_75t_L g30 ( 
.A(n_23),
.B(n_1),
.Y(n_30)
);

INVx11_ASAP7_75t_L g31 ( 
.A(n_16),
.Y(n_31)
);

INVx6_ASAP7_75t_L g49 ( 
.A(n_31),
.Y(n_49)
);

INVx4_ASAP7_75t_L g32 ( 
.A(n_17),
.Y(n_32)
);

INVx3_ASAP7_75t_L g43 ( 
.A(n_32),
.Y(n_43)
);

INVx4_ASAP7_75t_L g33 ( 
.A(n_17),
.Y(n_33)
);

INVx3_ASAP7_75t_L g46 ( 
.A(n_33),
.Y(n_46)
);

INVx6_ASAP7_75t_L g34 ( 
.A(n_20),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_34),
.Y(n_40)
);

INVx3_ASAP7_75t_L g35 ( 
.A(n_20),
.Y(n_35)
);

INVx2_ASAP7_75t_L g48 ( 
.A(n_35),
.Y(n_48)
);

INVx4_ASAP7_75t_L g36 ( 
.A(n_21),
.Y(n_36)
);

BUFx2_ASAP7_75t_L g39 ( 
.A(n_36),
.Y(n_39)
);

AOI22xp33_ASAP7_75t_SL g38 ( 
.A1(n_34),
.A2(n_24),
.B1(n_27),
.B2(n_18),
.Y(n_38)
);

CKINVDCx16_ASAP7_75t_R g63 ( 
.A(n_38),
.Y(n_63)
);

OAI22xp5_ASAP7_75t_L g41 ( 
.A1(n_34),
.A2(n_24),
.B1(n_27),
.B2(n_26),
.Y(n_41)
);

OAI22xp5_ASAP7_75t_L g65 ( 
.A1(n_41),
.A2(n_35),
.B1(n_19),
.B2(n_33),
.Y(n_65)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_28),
.Y(n_42)
);

INVx6_ASAP7_75t_L g62 ( 
.A(n_42),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_28),
.Y(n_44)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_44),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g47 ( 
.A(n_29),
.B(n_13),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_47),
.B(n_50),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_30),
.B(n_13),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_L g51 ( 
.A(n_45),
.B(n_23),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_L g72 ( 
.A(n_51),
.B(n_55),
.Y(n_72)
);

INVx13_ASAP7_75t_L g52 ( 
.A(n_37),
.Y(n_52)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_52),
.Y(n_75)
);

INVx3_ASAP7_75t_L g53 ( 
.A(n_48),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_53),
.B(n_60),
.Y(n_73)
);

CKINVDCx20_ASAP7_75t_R g55 ( 
.A(n_37),
.Y(n_55)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_39),
.Y(n_56)
);

AND2x2_ASAP7_75t_L g70 ( 
.A(n_56),
.B(n_49),
.Y(n_70)
);

OAI21xp5_ASAP7_75t_L g57 ( 
.A1(n_41),
.A2(n_23),
.B(n_18),
.Y(n_57)
);

AOI21xp5_ASAP7_75t_L g71 ( 
.A1(n_57),
.A2(n_25),
.B(n_2),
.Y(n_71)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_39),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g80 ( 
.A(n_58),
.Y(n_80)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_39),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_43),
.B(n_19),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_SL g74 ( 
.A(n_61),
.B(n_25),
.Y(n_74)
);

INVx13_ASAP7_75t_L g64 ( 
.A(n_42),
.Y(n_64)
);

INVxp67_ASAP7_75t_L g79 ( 
.A(n_64),
.Y(n_79)
);

AOI22xp5_ASAP7_75t_L g69 ( 
.A1(n_65),
.A2(n_46),
.B1(n_33),
.B2(n_36),
.Y(n_69)
);

O2A1O1Ixp33_ASAP7_75t_L g66 ( 
.A1(n_63),
.A2(n_46),
.B(n_43),
.C(n_36),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_L g83 ( 
.A(n_66),
.B(n_77),
.Y(n_83)
);

OAI22xp5_ASAP7_75t_SL g67 ( 
.A1(n_57),
.A2(n_65),
.B1(n_51),
.B2(n_48),
.Y(n_67)
);

OAI22xp5_ASAP7_75t_L g89 ( 
.A1(n_67),
.A2(n_69),
.B1(n_71),
.B2(n_62),
.Y(n_89)
);

NOR2xp67_ASAP7_75t_L g68 ( 
.A(n_59),
.B(n_55),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_SL g93 ( 
.A(n_68),
.B(n_74),
.Y(n_93)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_70),
.Y(n_84)
);

MAJIxp5_ASAP7_75t_L g76 ( 
.A(n_53),
.B(n_40),
.C(n_44),
.Y(n_76)
);

MAJIxp5_ASAP7_75t_L g91 ( 
.A(n_76),
.B(n_80),
.C(n_70),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_L g77 ( 
.A(n_56),
.B(n_40),
.Y(n_77)
);

BUFx2_ASAP7_75t_L g78 ( 
.A(n_64),
.Y(n_78)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_78),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_72),
.B(n_52),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g98 ( 
.A(n_81),
.B(n_82),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_SL g82 ( 
.A(n_67),
.B(n_54),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_L g86 ( 
.A(n_77),
.B(n_60),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_SL g94 ( 
.A(n_86),
.B(n_89),
.Y(n_94)
);

XNOR2xp5_ASAP7_75t_L g87 ( 
.A(n_71),
.B(n_31),
.Y(n_87)
);

XOR2xp5_ASAP7_75t_L g100 ( 
.A(n_87),
.B(n_91),
.Y(n_100)
);

OAI22xp5_ASAP7_75t_SL g88 ( 
.A1(n_69),
.A2(n_54),
.B1(n_62),
.B2(n_58),
.Y(n_88)
);

INVxp67_ASAP7_75t_L g103 ( 
.A(n_88),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_L g90 ( 
.A(n_75),
.B(n_32),
.Y(n_90)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_90),
.Y(n_95)
);

CKINVDCx20_ASAP7_75t_R g92 ( 
.A(n_73),
.Y(n_92)
);

NAND3xp33_ASAP7_75t_L g96 ( 
.A(n_92),
.B(n_8),
.C(n_10),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_SL g108 ( 
.A(n_96),
.B(n_102),
.Y(n_108)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_86),
.Y(n_97)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_97),
.Y(n_110)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_85),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_SL g106 ( 
.A(n_99),
.B(n_104),
.Y(n_106)
);

INVx2_ASAP7_75t_L g101 ( 
.A(n_91),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_101),
.B(n_70),
.Y(n_111)
);

NAND3xp33_ASAP7_75t_L g102 ( 
.A(n_93),
.B(n_9),
.C(n_10),
.Y(n_102)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_90),
.Y(n_104)
);

AOI22x1_ASAP7_75t_L g105 ( 
.A1(n_94),
.A2(n_83),
.B1(n_88),
.B2(n_87),
.Y(n_105)
);

OAI21xp5_ASAP7_75t_SL g116 ( 
.A1(n_105),
.A2(n_107),
.B(n_112),
.Y(n_116)
);

XNOR2x1_ASAP7_75t_L g107 ( 
.A(n_100),
.B(n_84),
.Y(n_107)
);

MAJIxp5_ASAP7_75t_L g109 ( 
.A(n_100),
.B(n_84),
.C(n_76),
.Y(n_109)
);

MAJIxp5_ASAP7_75t_L g115 ( 
.A(n_109),
.B(n_113),
.C(n_103),
.Y(n_115)
);

AOI21xp5_ASAP7_75t_L g117 ( 
.A1(n_111),
.A2(n_79),
.B(n_2),
.Y(n_117)
);

CKINVDCx20_ASAP7_75t_R g112 ( 
.A(n_95),
.Y(n_112)
);

MAJIxp5_ASAP7_75t_L g113 ( 
.A(n_101),
.B(n_98),
.C(n_83),
.Y(n_113)
);

A2O1A1O1Ixp25_ASAP7_75t_L g114 ( 
.A1(n_107),
.A2(n_103),
.B(n_66),
.C(n_14),
.D(n_16),
.Y(n_114)
);

OAI21xp5_ASAP7_75t_L g125 ( 
.A1(n_114),
.A2(n_117),
.B(n_118),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_L g121 ( 
.A(n_115),
.B(n_119),
.Y(n_121)
);

AOI21xp5_ASAP7_75t_L g118 ( 
.A1(n_106),
.A2(n_1),
.B(n_4),
.Y(n_118)
);

XOR2xp5_ASAP7_75t_L g119 ( 
.A(n_113),
.B(n_31),
.Y(n_119)
);

AOI221xp5_ASAP7_75t_L g120 ( 
.A1(n_105),
.A2(n_79),
.B1(n_15),
.B2(n_14),
.C(n_21),
.Y(n_120)
);

OAI22xp5_ASAP7_75t_SL g124 ( 
.A1(n_120),
.A2(n_49),
.B1(n_78),
.B2(n_16),
.Y(n_124)
);

AOI21xp5_ASAP7_75t_SL g122 ( 
.A1(n_116),
.A2(n_110),
.B(n_108),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_L g126 ( 
.A(n_122),
.B(n_123),
.Y(n_126)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_120),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_L g129 ( 
.A(n_124),
.B(n_15),
.Y(n_129)
);

XOR2xp5_ASAP7_75t_L g127 ( 
.A(n_121),
.B(n_80),
.Y(n_127)
);

OAI21xp5_ASAP7_75t_L g132 ( 
.A1(n_127),
.A2(n_4),
.B(n_22),
.Y(n_132)
);

OAI22xp5_ASAP7_75t_L g128 ( 
.A1(n_125),
.A2(n_6),
.B1(n_7),
.B2(n_8),
.Y(n_128)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_128),
.Y(n_130)
);

NOR3xp33_ASAP7_75t_L g131 ( 
.A(n_129),
.B(n_122),
.C(n_7),
.Y(n_131)
);

INVxp67_ASAP7_75t_L g134 ( 
.A(n_131),
.Y(n_134)
);

OAI21x1_ASAP7_75t_L g133 ( 
.A1(n_132),
.A2(n_126),
.B(n_22),
.Y(n_133)
);

MAJIxp5_ASAP7_75t_L g135 ( 
.A(n_133),
.B(n_130),
.C(n_127),
.Y(n_135)
);

XOR2xp5_ASAP7_75t_L g136 ( 
.A(n_135),
.B(n_134),
.Y(n_136)
);


endmodule