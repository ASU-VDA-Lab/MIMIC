module fake_netlist_6_3438_n_1903 (n_52, n_16, n_1, n_91, n_119, n_46, n_146, n_163, n_18, n_21, n_147, n_154, n_88, n_3, n_98, n_113, n_39, n_63, n_73, n_4, n_148, n_138, n_22, n_161, n_68, n_166, n_28, n_50, n_158, n_49, n_7, n_83, n_5, n_101, n_167, n_144, n_174, n_127, n_125, n_153, n_168, n_77, n_156, n_149, n_152, n_106, n_92, n_145, n_42, n_133, n_96, n_8, n_90, n_160, n_24, n_105, n_131, n_54, n_132, n_102, n_0, n_87, n_32, n_66, n_85, n_99, n_78, n_84, n_130, n_164, n_100, n_129, n_13, n_121, n_11, n_137, n_17, n_23, n_142, n_20, n_143, n_2, n_19, n_47, n_62, n_29, n_155, n_75, n_109, n_150, n_122, n_45, n_34, n_140, n_70, n_120, n_37, n_15, n_67, n_33, n_82, n_27, n_38, n_110, n_151, n_61, n_112, n_172, n_81, n_59, n_76, n_36, n_26, n_124, n_55, n_126, n_94, n_97, n_108, n_58, n_116, n_64, n_117, n_118, n_48, n_65, n_25, n_40, n_93, n_80, n_141, n_135, n_165, n_139, n_41, n_134, n_114, n_86, n_104, n_95, n_9, n_107, n_10, n_71, n_74, n_6, n_14, n_123, n_136, n_72, n_89, n_173, n_103, n_111, n_60, n_159, n_157, n_162, n_170, n_35, n_115, n_12, n_69, n_128, n_30, n_79, n_43, n_171, n_31, n_57, n_169, n_53, n_51, n_44, n_56, n_1903);

input n_52;
input n_16;
input n_1;
input n_91;
input n_119;
input n_46;
input n_146;
input n_163;
input n_18;
input n_21;
input n_147;
input n_154;
input n_88;
input n_3;
input n_98;
input n_113;
input n_39;
input n_63;
input n_73;
input n_4;
input n_148;
input n_138;
input n_22;
input n_161;
input n_68;
input n_166;
input n_28;
input n_50;
input n_158;
input n_49;
input n_7;
input n_83;
input n_5;
input n_101;
input n_167;
input n_144;
input n_174;
input n_127;
input n_125;
input n_153;
input n_168;
input n_77;
input n_156;
input n_149;
input n_152;
input n_106;
input n_92;
input n_145;
input n_42;
input n_133;
input n_96;
input n_8;
input n_90;
input n_160;
input n_24;
input n_105;
input n_131;
input n_54;
input n_132;
input n_102;
input n_0;
input n_87;
input n_32;
input n_66;
input n_85;
input n_99;
input n_78;
input n_84;
input n_130;
input n_164;
input n_100;
input n_129;
input n_13;
input n_121;
input n_11;
input n_137;
input n_17;
input n_23;
input n_142;
input n_20;
input n_143;
input n_2;
input n_19;
input n_47;
input n_62;
input n_29;
input n_155;
input n_75;
input n_109;
input n_150;
input n_122;
input n_45;
input n_34;
input n_140;
input n_70;
input n_120;
input n_37;
input n_15;
input n_67;
input n_33;
input n_82;
input n_27;
input n_38;
input n_110;
input n_151;
input n_61;
input n_112;
input n_172;
input n_81;
input n_59;
input n_76;
input n_36;
input n_26;
input n_124;
input n_55;
input n_126;
input n_94;
input n_97;
input n_108;
input n_58;
input n_116;
input n_64;
input n_117;
input n_118;
input n_48;
input n_65;
input n_25;
input n_40;
input n_93;
input n_80;
input n_141;
input n_135;
input n_165;
input n_139;
input n_41;
input n_134;
input n_114;
input n_86;
input n_104;
input n_95;
input n_9;
input n_107;
input n_10;
input n_71;
input n_74;
input n_6;
input n_14;
input n_123;
input n_136;
input n_72;
input n_89;
input n_173;
input n_103;
input n_111;
input n_60;
input n_159;
input n_157;
input n_162;
input n_170;
input n_35;
input n_115;
input n_12;
input n_69;
input n_128;
input n_30;
input n_79;
input n_43;
input n_171;
input n_31;
input n_57;
input n_169;
input n_53;
input n_51;
input n_44;
input n_56;

output n_1903;

wire n_992;
wire n_1671;
wire n_801;
wire n_1613;
wire n_1234;
wire n_1458;
wire n_1199;
wire n_1674;
wire n_741;
wire n_1027;
wire n_1351;
wire n_625;
wire n_1189;
wire n_223;
wire n_1212;
wire n_226;
wire n_208;
wire n_726;
wire n_212;
wire n_700;
wire n_1307;
wire n_1038;
wire n_578;
wire n_1581;
wire n_1003;
wire n_365;
wire n_1237;
wire n_1061;
wire n_1357;
wire n_1853;
wire n_783;
wire n_1738;
wire n_798;
wire n_188;
wire n_1575;
wire n_1854;
wire n_509;
wire n_1342;
wire n_245;
wire n_1209;
wire n_1348;
wire n_1387;
wire n_677;
wire n_1708;
wire n_805;
wire n_1151;
wire n_396;
wire n_1739;
wire n_350;
wire n_1380;
wire n_442;
wire n_480;
wire n_1402;
wire n_1691;
wire n_1688;
wire n_1009;
wire n_1743;
wire n_1160;
wire n_883;
wire n_1238;
wire n_1724;
wire n_1032;
wire n_1247;
wire n_1547;
wire n_1553;
wire n_893;
wire n_1099;
wire n_1264;
wire n_1192;
wire n_471;
wire n_1844;
wire n_424;
wire n_1700;
wire n_1555;
wire n_1415;
wire n_1370;
wire n_1786;
wire n_369;
wire n_287;
wire n_415;
wire n_830;
wire n_230;
wire n_461;
wire n_873;
wire n_383;
wire n_1285;
wire n_1371;
wire n_200;
wire n_447;
wire n_1803;
wire n_1172;
wire n_852;
wire n_229;
wire n_1590;
wire n_1532;
wire n_1393;
wire n_1517;
wire n_1867;
wire n_1704;
wire n_1078;
wire n_250;
wire n_544;
wire n_1711;
wire n_1140;
wire n_1444;
wire n_1670;
wire n_1603;
wire n_1579;
wire n_1263;
wire n_836;
wire n_375;
wire n_522;
wire n_1261;
wire n_945;
wire n_1649;
wire n_1511;
wire n_1143;
wire n_1422;
wire n_1232;
wire n_1772;
wire n_1572;
wire n_616;
wire n_658;
wire n_1874;
wire n_1119;
wire n_428;
wire n_1433;
wire n_1902;
wire n_1842;
wire n_1620;
wire n_1735;
wire n_1541;
wire n_1300;
wire n_641;
wire n_822;
wire n_693;
wire n_1313;
wire n_1056;
wire n_758;
wire n_516;
wire n_1455;
wire n_1163;
wire n_1180;
wire n_943;
wire n_1798;
wire n_1550;
wire n_491;
wire n_1591;
wire n_772;
wire n_1344;
wire n_666;
wire n_371;
wire n_940;
wire n_770;
wire n_567;
wire n_1781;
wire n_405;
wire n_213;
wire n_538;
wire n_1106;
wire n_886;
wire n_1471;
wire n_343;
wire n_953;
wire n_1094;
wire n_1345;
wire n_1820;
wire n_494;
wire n_539;
wire n_493;
wire n_454;
wire n_1421;
wire n_638;
wire n_1404;
wire n_1211;
wire n_381;
wire n_887;
wire n_1660;
wire n_1280;
wire n_713;
wire n_1400;
wire n_1467;
wire n_976;
wire n_224;
wire n_1445;
wire n_1526;
wire n_1560;
wire n_734;
wire n_1088;
wire n_1894;
wire n_196;
wire n_1231;
wire n_917;
wire n_574;
wire n_907;
wire n_1446;
wire n_659;
wire n_1815;
wire n_407;
wire n_913;
wire n_1658;
wire n_808;
wire n_867;
wire n_1230;
wire n_473;
wire n_1193;
wire n_1054;
wire n_559;
wire n_1333;
wire n_1648;
wire n_1644;
wire n_1558;
wire n_1732;
wire n_281;
wire n_551;
wire n_699;
wire n_564;
wire n_451;
wire n_824;
wire n_279;
wire n_686;
wire n_757;
wire n_594;
wire n_1641;
wire n_577;
wire n_1843;
wire n_619;
wire n_1367;
wire n_1336;
wire n_521;
wire n_572;
wire n_395;
wire n_813;
wire n_1481;
wire n_323;
wire n_606;
wire n_1441;
wire n_818;
wire n_1123;
wire n_1309;
wire n_513;
wire n_645;
wire n_1381;
wire n_331;
wire n_1699;
wire n_916;
wire n_483;
wire n_608;
wire n_261;
wire n_630;
wire n_541;
wire n_512;
wire n_433;
wire n_792;
wire n_476;
wire n_1328;
wire n_219;
wire n_264;
wire n_263;
wire n_1162;
wire n_860;
wire n_1530;
wire n_788;
wire n_939;
wire n_1543;
wire n_821;
wire n_938;
wire n_1302;
wire n_1068;
wire n_1599;
wire n_329;
wire n_982;
wire n_549;
wire n_1762;
wire n_1075;
wire n_408;
wire n_932;
wire n_237;
wire n_1876;
wire n_1895;
wire n_1697;
wire n_243;
wire n_979;
wire n_1873;
wire n_905;
wire n_1866;
wire n_1680;
wire n_175;
wire n_322;
wire n_993;
wire n_689;
wire n_354;
wire n_1330;
wire n_1413;
wire n_1605;
wire n_1278;
wire n_547;
wire n_558;
wire n_1064;
wire n_1396;
wire n_634;
wire n_966;
wire n_764;
wire n_1663;
wire n_692;
wire n_733;
wire n_1793;
wire n_1233;
wire n_1289;
wire n_487;
wire n_241;
wire n_1107;
wire n_1014;
wire n_1290;
wire n_1703;
wire n_882;
wire n_1354;
wire n_586;
wire n_423;
wire n_1875;
wire n_1865;
wire n_1701;
wire n_318;
wire n_1111;
wire n_1713;
wire n_715;
wire n_1251;
wire n_1265;
wire n_1726;
wire n_530;
wire n_1563;
wire n_277;
wire n_618;
wire n_1297;
wire n_1662;
wire n_1312;
wire n_199;
wire n_1167;
wire n_1359;
wire n_674;
wire n_871;
wire n_922;
wire n_268;
wire n_1335;
wire n_1760;
wire n_210;
wire n_1069;
wire n_1722;
wire n_1664;
wire n_612;
wire n_178;
wire n_247;
wire n_1165;
wire n_355;
wire n_702;
wire n_347;
wire n_1175;
wire n_328;
wire n_1386;
wire n_1896;
wire n_429;
wire n_1747;
wire n_1012;
wire n_195;
wire n_780;
wire n_675;
wire n_903;
wire n_1540;
wire n_1802;
wire n_1504;
wire n_286;
wire n_254;
wire n_1655;
wire n_242;
wire n_835;
wire n_928;
wire n_1214;
wire n_690;
wire n_850;
wire n_1801;
wire n_1886;
wire n_1654;
wire n_816;
wire n_1157;
wire n_1750;
wire n_1462;
wire n_1188;
wire n_1752;
wire n_877;
wire n_1813;
wire n_604;
wire n_825;
wire n_728;
wire n_1063;
wire n_1588;
wire n_267;
wire n_1124;
wire n_1624;
wire n_515;
wire n_598;
wire n_696;
wire n_1515;
wire n_961;
wire n_437;
wire n_1082;
wire n_1317;
wire n_593;
wire n_514;
wire n_687;
wire n_697;
wire n_890;
wire n_637;
wire n_295;
wire n_701;
wire n_950;
wire n_388;
wire n_190;
wire n_484;
wire n_1709;
wire n_1825;
wire n_1757;
wire n_1796;
wire n_1792;
wire n_891;
wire n_1412;
wire n_949;
wire n_1630;
wire n_678;
wire n_283;
wire n_507;
wire n_968;
wire n_909;
wire n_1369;
wire n_881;
wire n_1008;
wire n_760;
wire n_1546;
wire n_590;
wire n_362;
wire n_462;
wire n_1033;
wire n_1052;
wire n_1296;
wire n_304;
wire n_694;
wire n_1294;
wire n_1420;
wire n_1634;
wire n_297;
wire n_627;
wire n_595;
wire n_1767;
wire n_1779;
wire n_524;
wire n_1465;
wire n_342;
wire n_1858;
wire n_1044;
wire n_1712;
wire n_1391;
wire n_449;
wire n_1523;
wire n_1208;
wire n_1164;
wire n_1295;
wire n_1627;
wire n_1072;
wire n_1527;
wire n_1495;
wire n_1438;
wire n_495;
wire n_815;
wire n_1100;
wire n_585;
wire n_1487;
wire n_840;
wire n_874;
wire n_1756;
wire n_1128;
wire n_382;
wire n_673;
wire n_1071;
wire n_1067;
wire n_1565;
wire n_1493;
wire n_898;
wire n_255;
wire n_284;
wire n_865;
wire n_925;
wire n_1101;
wire n_1026;
wire n_1880;
wire n_289;
wire n_1364;
wire n_615;
wire n_1249;
wire n_1293;
wire n_1127;
wire n_1512;
wire n_1451;
wire n_320;
wire n_639;
wire n_963;
wire n_794;
wire n_727;
wire n_894;
wire n_1839;
wire n_685;
wire n_1765;
wire n_353;
wire n_605;
wire n_1514;
wire n_1863;
wire n_826;
wire n_1646;
wire n_872;
wire n_1139;
wire n_1714;
wire n_718;
wire n_1018;
wire n_1521;
wire n_1366;
wire n_542;
wire n_847;
wire n_644;
wire n_682;
wire n_851;
wire n_305;
wire n_996;
wire n_532;
wire n_1308;
wire n_1376;
wire n_1513;
wire n_413;
wire n_791;
wire n_510;
wire n_837;
wire n_1488;
wire n_1808;
wire n_948;
wire n_704;
wire n_977;
wire n_1005;
wire n_536;
wire n_1788;
wire n_622;
wire n_1469;
wire n_1838;
wire n_1835;
wire n_1766;
wire n_1776;
wire n_581;
wire n_765;
wire n_432;
wire n_987;
wire n_1492;
wire n_1340;
wire n_1771;
wire n_631;
wire n_720;
wire n_842;
wire n_1707;
wire n_1432;
wire n_843;
wire n_656;
wire n_989;
wire n_1277;
wire n_797;
wire n_1473;
wire n_1723;
wire n_1246;
wire n_1878;
wire n_899;
wire n_189;
wire n_738;
wire n_1304;
wire n_1035;
wire n_294;
wire n_499;
wire n_1426;
wire n_705;
wire n_1004;
wire n_1176;
wire n_1529;
wire n_1022;
wire n_614;
wire n_529;
wire n_425;
wire n_684;
wire n_1431;
wire n_1615;
wire n_1474;
wire n_1571;
wire n_1809;
wire n_1577;
wire n_1181;
wire n_1822;
wire n_486;
wire n_947;
wire n_1117;
wire n_1087;
wire n_1448;
wire n_648;
wire n_657;
wire n_1049;
wire n_1666;
wire n_1505;
wire n_803;
wire n_290;
wire n_1717;
wire n_926;
wire n_1817;
wire n_927;
wire n_1849;
wire n_919;
wire n_1698;
wire n_478;
wire n_929;
wire n_1228;
wire n_417;
wire n_446;
wire n_1568;
wire n_1490;
wire n_777;
wire n_1299;
wire n_272;
wire n_526;
wire n_1183;
wire n_1436;
wire n_1384;
wire n_293;
wire n_458;
wire n_1070;
wire n_998;
wire n_717;
wire n_1665;
wire n_1383;
wire n_1178;
wire n_1424;
wire n_1073;
wire n_1000;
wire n_796;
wire n_252;
wire n_1195;
wire n_1626;
wire n_1507;
wire n_184;
wire n_552;
wire n_1358;
wire n_1811;
wire n_1388;
wire n_216;
wire n_912;
wire n_1857;
wire n_1519;
wire n_745;
wire n_1284;
wire n_1604;
wire n_1142;
wire n_716;
wire n_1475;
wire n_623;
wire n_1048;
wire n_1201;
wire n_1398;
wire n_884;
wire n_1774;
wire n_1395;
wire n_731;
wire n_1502;
wire n_1659;
wire n_755;
wire n_931;
wire n_1021;
wire n_474;
wire n_527;
wire n_683;
wire n_811;
wire n_1207;
wire n_312;
wire n_1791;
wire n_1368;
wire n_1418;
wire n_958;
wire n_292;
wire n_1250;
wire n_1137;
wire n_1897;
wire n_880;
wire n_889;
wire n_1478;
wire n_589;
wire n_1310;
wire n_819;
wire n_1363;
wire n_1334;
wire n_767;
wire n_1314;
wire n_600;
wire n_964;
wire n_831;
wire n_1837;
wire n_477;
wire n_954;
wire n_864;
wire n_1110;
wire n_1410;
wire n_399;
wire n_1440;
wire n_1382;
wire n_1534;
wire n_1564;
wire n_1736;
wire n_211;
wire n_1483;
wire n_1834;
wire n_1372;
wire n_231;
wire n_1457;
wire n_505;
wire n_1719;
wire n_319;
wire n_1339;
wire n_1787;
wire n_537;
wire n_1427;
wire n_311;
wire n_1466;
wire n_403;
wire n_1080;
wire n_723;
wire n_1877;
wire n_596;
wire n_546;
wire n_562;
wire n_1141;
wire n_1268;
wire n_386;
wire n_1769;
wire n_1220;
wire n_1893;
wire n_556;
wire n_1755;
wire n_1602;
wire n_1136;
wire n_1125;
wire n_970;
wire n_642;
wire n_995;
wire n_276;
wire n_1159;
wire n_1092;
wire n_441;
wire n_221;
wire n_1060;
wire n_444;
wire n_1252;
wire n_1784;
wire n_1223;
wire n_303;
wire n_511;
wire n_193;
wire n_1286;
wire n_1775;
wire n_1773;
wire n_1053;
wire n_416;
wire n_1681;
wire n_520;
wire n_418;
wire n_1093;
wire n_1783;
wire n_1533;
wire n_1597;
wire n_266;
wire n_296;
wire n_775;
wire n_651;
wire n_1153;
wire n_439;
wire n_1618;
wire n_217;
wire n_518;
wire n_1531;
wire n_1185;
wire n_453;
wire n_215;
wire n_1745;
wire n_914;
wire n_759;
wire n_1831;
wire n_426;
wire n_317;
wire n_1653;
wire n_1679;
wire n_1625;
wire n_1453;
wire n_488;
wire n_497;
wire n_773;
wire n_1901;
wire n_920;
wire n_1374;
wire n_1315;
wire n_1647;
wire n_1224;
wire n_1614;
wire n_1459;
wire n_1892;
wire n_1135;
wire n_1179;
wire n_1169;
wire n_401;
wire n_324;
wire n_1617;
wire n_335;
wire n_1470;
wire n_463;
wire n_1243;
wire n_848;
wire n_301;
wire n_274;
wire n_1096;
wire n_1091;
wire n_1580;
wire n_1425;
wire n_1881;
wire n_1281;
wire n_1267;
wire n_1806;
wire n_983;
wire n_427;
wire n_1520;
wire n_496;
wire n_906;
wire n_1390;
wire n_688;
wire n_1077;
wire n_1733;
wire n_1419;
wire n_351;
wire n_259;
wire n_1731;
wire n_177;
wire n_1855;
wire n_1636;
wire n_1437;
wire n_1645;
wire n_1832;
wire n_385;
wire n_1687;
wire n_1439;
wire n_1323;
wire n_858;
wire n_1331;
wire n_613;
wire n_736;
wire n_501;
wire n_956;
wire n_960;
wire n_663;
wire n_856;
wire n_379;
wire n_778;
wire n_1668;
wire n_1134;
wire n_410;
wire n_1129;
wire n_554;
wire n_602;
wire n_1696;
wire n_1594;
wire n_664;
wire n_1869;
wire n_1764;
wire n_1429;
wire n_1610;
wire n_1889;
wire n_435;
wire n_793;
wire n_326;
wire n_587;
wire n_1593;
wire n_580;
wire n_762;
wire n_1030;
wire n_1202;
wire n_465;
wire n_1790;
wire n_1778;
wire n_1635;
wire n_1079;
wire n_341;
wire n_1744;
wire n_828;
wire n_607;
wire n_316;
wire n_419;
wire n_1551;
wire n_1103;
wire n_1203;
wire n_820;
wire n_951;
wire n_725;
wire n_952;
wire n_999;
wire n_358;
wire n_1254;
wire n_186;
wire n_368;
wire n_575;
wire n_994;
wire n_1508;
wire n_732;
wire n_974;
wire n_392;
wire n_724;
wire n_1020;
wire n_1042;
wire n_628;
wire n_1273;
wire n_1434;
wire n_1573;
wire n_1728;
wire n_557;
wire n_1871;
wire n_349;
wire n_617;
wire n_845;
wire n_807;
wire n_1036;
wire n_1138;
wire n_1661;
wire n_1275;
wire n_485;
wire n_1549;
wire n_443;
wire n_1510;
wire n_892;
wire n_768;
wire n_421;
wire n_1468;
wire n_1859;
wire n_238;
wire n_1095;
wire n_1595;
wire n_202;
wire n_1718;
wire n_1749;
wire n_1683;
wire n_597;
wire n_280;
wire n_1270;
wire n_1187;
wire n_610;
wire n_1403;
wire n_1669;
wire n_1852;
wire n_1024;
wire n_1768;
wire n_198;
wire n_1847;
wire n_179;
wire n_248;
wire n_517;
wire n_1667;
wire n_667;
wire n_1206;
wire n_621;
wire n_1037;
wire n_1397;
wire n_1279;
wire n_1115;
wire n_750;
wire n_901;
wire n_1499;
wire n_468;
wire n_923;
wire n_504;
wire n_1409;
wire n_1841;
wire n_1639;
wire n_1623;
wire n_183;
wire n_1015;
wire n_1503;
wire n_466;
wire n_1057;
wire n_603;
wire n_991;
wire n_1657;
wire n_235;
wire n_1126;
wire n_340;
wire n_710;
wire n_1108;
wire n_1818;
wire n_1182;
wire n_1298;
wire n_1611;
wire n_785;
wire n_746;
wire n_609;
wire n_1601;
wire n_1686;
wire n_1356;
wire n_1589;
wire n_1740;
wire n_1497;
wire n_1168;
wire n_1216;
wire n_1320;
wire n_1430;
wire n_1316;
wire n_1287;
wire n_1452;
wire n_1622;
wire n_1586;
wire n_302;
wire n_1694;
wire n_380;
wire n_1535;
wire n_1596;
wire n_1190;
wire n_1734;
wire n_397;
wire n_1262;
wire n_218;
wire n_1891;
wire n_1213;
wire n_1350;
wire n_1673;
wire n_1715;
wire n_1443;
wire n_1272;
wire n_239;
wire n_782;
wire n_1539;
wire n_490;
wire n_220;
wire n_809;
wire n_1043;
wire n_1797;
wire n_1608;
wire n_986;
wire n_1472;
wire n_1081;
wire n_402;
wire n_1870;
wire n_352;
wire n_1692;
wire n_800;
wire n_1084;
wire n_1171;
wire n_460;
wire n_1827;
wire n_1361;
wire n_1864;
wire n_1491;
wire n_662;
wire n_374;
wire n_1152;
wire n_1840;
wire n_1705;
wire n_450;
wire n_1684;
wire n_921;
wire n_1346;
wire n_711;
wire n_1642;
wire n_579;
wire n_1352;
wire n_937;
wire n_1682;
wire n_370;
wire n_1695;
wire n_1828;
wire n_650;
wire n_1046;
wire n_1145;
wire n_330;
wire n_1121;
wire n_1102;
wire n_972;
wire n_1405;
wire n_258;
wire n_1406;
wire n_456;
wire n_1332;
wire n_260;
wire n_313;
wire n_624;
wire n_962;
wire n_1041;
wire n_565;
wire n_356;
wire n_1569;
wire n_936;
wire n_1883;
wire n_1288;
wire n_1186;
wire n_1062;
wire n_885;
wire n_896;
wire n_654;
wire n_411;
wire n_1222;
wire n_599;
wire n_776;
wire n_321;
wire n_1823;
wire n_227;
wire n_1720;
wire n_204;
wire n_482;
wire n_934;
wire n_1637;
wire n_1407;
wire n_1795;
wire n_420;
wire n_1341;
wire n_394;
wire n_1456;
wire n_1845;
wire n_1489;
wire n_942;
wire n_1524;
wire n_543;
wire n_1496;
wire n_1271;
wire n_1545;
wire n_1355;
wire n_1225;
wire n_1544;
wire n_1485;
wire n_325;
wire n_1640;
wire n_804;
wire n_464;
wire n_1846;
wire n_533;
wire n_806;
wire n_959;
wire n_879;
wire n_584;
wire n_244;
wire n_1343;
wire n_1522;
wire n_548;
wire n_1782;
wire n_282;
wire n_1676;
wire n_833;
wire n_1830;
wire n_1567;
wire n_523;
wire n_1319;
wire n_707;
wire n_345;
wire n_1900;
wire n_799;
wire n_1548;
wire n_1155;
wire n_273;
wire n_1633;
wire n_787;
wire n_1416;
wire n_1528;
wire n_1146;
wire n_1086;
wire n_1066;
wire n_1282;
wire n_550;
wire n_275;
wire n_652;
wire n_560;
wire n_1484;
wire n_1321;
wire n_1241;
wire n_1672;
wire n_569;
wire n_1758;
wire n_737;
wire n_1318;
wire n_1235;
wire n_1229;
wire n_306;
wire n_1292;
wire n_1373;
wire n_346;
wire n_1029;
wire n_1447;
wire n_790;
wire n_1706;
wire n_1498;
wire n_1210;
wire n_299;
wire n_1248;
wire n_1556;
wire n_902;
wire n_333;
wire n_1047;
wire n_1385;
wire n_431;
wire n_459;
wire n_1269;
wire n_502;
wire n_672;
wire n_1257;
wire n_1751;
wire n_285;
wire n_1375;
wire n_655;
wire n_706;
wire n_1045;
wire n_1650;
wire n_786;
wire n_1794;
wire n_1236;
wire n_1559;
wire n_1725;
wire n_1872;
wire n_834;
wire n_743;
wire n_766;
wire n_430;
wire n_1741;
wire n_1325;
wire n_1002;
wire n_1746;
wire n_545;
wire n_489;
wire n_1804;
wire n_1727;
wire n_251;
wire n_1019;
wire n_636;
wire n_729;
wire n_876;
wire n_774;
wire n_1337;
wire n_660;
wire n_438;
wire n_1477;
wire n_1360;
wire n_1860;
wire n_1200;
wire n_479;
wire n_1607;
wire n_1353;
wire n_1777;
wire n_1454;
wire n_869;
wire n_1154;
wire n_1113;
wire n_1600;
wire n_646;
wire n_528;
wire n_391;
wire n_1098;
wire n_1329;
wire n_817;
wire n_262;
wire n_187;
wire n_897;
wire n_846;
wire n_841;
wire n_1476;
wire n_1001;
wire n_508;
wire n_1800;
wire n_1050;
wire n_1411;
wire n_1463;
wire n_1177;
wire n_332;
wire n_1150;
wire n_1742;
wire n_1562;
wire n_1690;
wire n_398;
wire n_1191;
wire n_1826;
wire n_566;
wire n_1023;
wire n_1882;
wire n_1076;
wire n_1118;
wire n_194;
wire n_1007;
wire n_1807;
wire n_1378;
wire n_855;
wire n_1592;
wire n_1759;
wire n_1814;
wire n_1631;
wire n_591;
wire n_1377;
wire n_1879;
wire n_256;
wire n_853;
wire n_440;
wire n_695;
wire n_1542;
wire n_875;
wire n_209;
wire n_367;
wire n_680;
wire n_1678;
wire n_661;
wire n_1716;
wire n_278;
wire n_1256;
wire n_671;
wire n_933;
wire n_740;
wire n_703;
wire n_978;
wire n_384;
wire n_1291;
wire n_1217;
wire n_751;
wire n_749;
wire n_1824;
wire n_310;
wire n_1628;
wire n_1324;
wire n_1399;
wire n_1435;
wire n_969;
wire n_988;
wire n_1065;
wire n_1401;
wire n_1255;
wire n_568;
wire n_1516;
wire n_1536;
wire n_180;
wire n_1204;
wire n_823;
wire n_1132;
wire n_643;
wire n_233;
wire n_698;
wire n_1074;
wire n_1394;
wire n_1327;
wire n_1326;
wire n_739;
wire n_400;
wire n_955;
wire n_337;
wire n_1379;
wire n_214;
wire n_246;
wire n_1338;
wire n_1097;
wire n_935;
wire n_781;
wire n_789;
wire n_1554;
wire n_1130;
wire n_181;
wire n_1810;
wire n_182;
wire n_573;
wire n_769;
wire n_676;
wire n_327;
wire n_1120;
wire n_832;
wire n_1583;
wire n_1730;
wire n_555;
wire n_389;
wire n_814;
wire n_1643;
wire n_1729;
wire n_669;
wire n_176;
wire n_300;
wire n_222;
wire n_747;
wire n_1389;
wire n_1105;
wire n_721;
wire n_1461;
wire n_742;
wire n_535;
wire n_691;
wire n_372;
wire n_314;
wire n_1408;
wire n_378;
wire n_1196;
wire n_377;
wire n_1598;
wire n_863;
wire n_601;
wire n_338;
wire n_1283;
wire n_918;
wire n_748;
wire n_506;
wire n_1114;
wire n_1785;
wire n_763;
wire n_1147;
wire n_1848;
wire n_360;
wire n_1754;
wire n_1506;
wire n_1652;
wire n_1812;
wire n_957;
wire n_895;
wire n_866;
wire n_1227;
wire n_191;
wire n_387;
wire n_452;
wire n_744;
wire n_971;
wire n_946;
wire n_344;
wire n_761;
wire n_1303;
wire n_1205;
wire n_1258;
wire n_1392;
wire n_1173;
wire n_525;
wire n_1677;
wire n_1116;
wire n_611;
wire n_1570;
wire n_1702;
wire n_1219;
wire n_1780;
wire n_1689;
wire n_1174;
wire n_1016;
wire n_1347;
wire n_795;
wire n_1501;
wire n_1221;
wire n_1245;
wire n_838;
wire n_647;
wire n_197;
wire n_844;
wire n_448;
wire n_1017;
wire n_1083;
wire n_445;
wire n_1561;
wire n_930;
wire n_888;
wire n_1112;
wire n_234;
wire n_910;
wire n_1656;
wire n_1721;
wire n_1460;
wire n_911;
wire n_1464;
wire n_236;
wire n_653;
wire n_1737;
wire n_1414;
wire n_752;
wire n_908;
wire n_944;
wire n_576;
wire n_1028;
wire n_472;
wire n_270;
wire n_414;
wire n_563;
wire n_1011;
wire n_1566;
wire n_1215;
wire n_839;
wire n_708;
wire n_668;
wire n_626;
wire n_990;
wire n_1500;
wire n_779;
wire n_1821;
wire n_1537;
wire n_1104;
wire n_854;
wire n_1058;
wire n_498;
wire n_1122;
wire n_870;
wire n_904;
wire n_1253;
wire n_709;
wire n_1266;
wire n_366;
wire n_1509;
wire n_1693;
wire n_1109;
wire n_185;
wire n_712;
wire n_348;
wire n_1276;
wire n_376;
wire n_390;
wire n_1148;
wire n_334;
wire n_1161;
wire n_1085;
wire n_232;
wire n_1239;
wire n_771;
wire n_1584;
wire n_470;
wire n_475;
wire n_924;
wire n_298;
wire n_1582;
wire n_492;
wire n_1149;
wire n_265;
wire n_1184;
wire n_228;
wire n_719;
wire n_1525;
wire n_455;
wire n_1585;
wire n_1851;
wire n_363;
wire n_1799;
wire n_1090;
wire n_592;
wire n_1816;
wire n_1518;
wire n_829;
wire n_1156;
wire n_1362;
wire n_393;
wire n_984;
wire n_1829;
wire n_503;
wire n_1450;
wire n_1638;
wire n_868;
wire n_570;
wire n_859;
wire n_406;
wire n_735;
wire n_1789;
wire n_1770;
wire n_878;
wire n_620;
wire n_519;
wire n_307;
wire n_469;
wire n_1218;
wire n_500;
wire n_1482;
wire n_981;
wire n_714;
wire n_1349;
wire n_291;
wire n_1144;
wire n_357;
wire n_985;
wire n_481;
wire n_997;
wire n_1710;
wire n_1301;
wire n_802;
wire n_561;
wire n_980;
wire n_1306;
wire n_1651;
wire n_1198;
wire n_1609;
wire n_436;
wire n_409;
wire n_1244;
wire n_1685;
wire n_1763;
wire n_1574;
wire n_240;
wire n_756;
wire n_1619;
wire n_1606;
wire n_810;
wire n_1133;
wire n_635;
wire n_1194;
wire n_1051;
wire n_253;
wire n_1552;
wire n_583;
wire n_249;
wire n_201;
wire n_1039;
wire n_1442;
wire n_1034;
wire n_1480;
wire n_1158;
wire n_754;
wire n_941;
wire n_975;
wire n_1031;
wire n_1305;
wire n_553;
wire n_849;
wire n_753;
wire n_1753;
wire n_467;
wire n_269;
wire n_359;
wire n_973;
wire n_1479;
wire n_1055;
wire n_1675;
wire n_582;
wire n_861;
wire n_857;
wire n_967;
wire n_571;
wire n_271;
wire n_404;
wire n_1884;
wire n_206;
wire n_679;
wire n_633;
wire n_1170;
wire n_665;
wire n_1629;
wire n_588;
wire n_225;
wire n_1260;
wire n_308;
wire n_309;
wire n_1819;
wire n_1010;
wire n_1040;
wire n_915;
wire n_632;
wire n_1166;
wire n_812;
wire n_1131;
wire n_1761;
wire n_534;
wire n_1578;
wire n_1006;
wire n_1861;
wire n_373;
wire n_1632;
wire n_1890;
wire n_1805;
wire n_257;
wire n_1557;
wire n_1888;
wire n_1833;
wire n_730;
wire n_1311;
wire n_1494;
wire n_670;
wire n_203;
wire n_1850;
wire n_1898;
wire n_1868;
wire n_207;
wire n_1089;
wire n_1887;
wire n_1587;
wire n_1365;
wire n_1417;
wire n_205;
wire n_1242;
wire n_1836;
wire n_681;
wire n_1226;
wire n_1274;
wire n_1486;
wire n_412;
wire n_640;
wire n_1322;
wire n_965;
wire n_1899;
wire n_1428;
wire n_1616;
wire n_1576;
wire n_1856;
wire n_1862;
wire n_339;
wire n_784;
wire n_434;
wire n_315;
wire n_288;
wire n_1059;
wire n_1197;
wire n_422;
wire n_722;
wire n_862;
wire n_540;
wire n_1423;
wire n_457;
wire n_364;
wire n_629;
wire n_1621;
wire n_1748;
wire n_900;
wire n_1449;
wire n_531;
wire n_827;
wire n_361;
wire n_1025;
wire n_336;
wire n_1885;
wire n_1013;
wire n_1259;
wire n_192;
wire n_1538;
wire n_649;
wire n_1612;
wire n_1240;

CKINVDCx5p33_ASAP7_75t_R g175 ( 
.A(n_102),
.Y(n_175)
);

CKINVDCx5p33_ASAP7_75t_R g176 ( 
.A(n_158),
.Y(n_176)
);

BUFx6f_ASAP7_75t_L g177 ( 
.A(n_140),
.Y(n_177)
);

INVx1_ASAP7_75t_SL g178 ( 
.A(n_88),
.Y(n_178)
);

CKINVDCx5p33_ASAP7_75t_R g179 ( 
.A(n_126),
.Y(n_179)
);

BUFx6f_ASAP7_75t_L g180 ( 
.A(n_67),
.Y(n_180)
);

INVx1_ASAP7_75t_SL g181 ( 
.A(n_69),
.Y(n_181)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_110),
.Y(n_182)
);

CKINVDCx20_ASAP7_75t_R g183 ( 
.A(n_141),
.Y(n_183)
);

CKINVDCx20_ASAP7_75t_R g184 ( 
.A(n_89),
.Y(n_184)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_108),
.Y(n_185)
);

CKINVDCx5p33_ASAP7_75t_R g186 ( 
.A(n_32),
.Y(n_186)
);

CKINVDCx5p33_ASAP7_75t_R g187 ( 
.A(n_46),
.Y(n_187)
);

INVx2_ASAP7_75t_L g188 ( 
.A(n_70),
.Y(n_188)
);

BUFx5_ASAP7_75t_L g189 ( 
.A(n_34),
.Y(n_189)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_107),
.Y(n_190)
);

CKINVDCx5p33_ASAP7_75t_R g191 ( 
.A(n_59),
.Y(n_191)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_123),
.Y(n_192)
);

CKINVDCx20_ASAP7_75t_R g193 ( 
.A(n_13),
.Y(n_193)
);

CKINVDCx5p33_ASAP7_75t_R g194 ( 
.A(n_48),
.Y(n_194)
);

CKINVDCx5p33_ASAP7_75t_R g195 ( 
.A(n_104),
.Y(n_195)
);

CKINVDCx5p33_ASAP7_75t_R g196 ( 
.A(n_2),
.Y(n_196)
);

CKINVDCx5p33_ASAP7_75t_R g197 ( 
.A(n_43),
.Y(n_197)
);

CKINVDCx5p33_ASAP7_75t_R g198 ( 
.A(n_42),
.Y(n_198)
);

INVx2_ASAP7_75t_L g199 ( 
.A(n_46),
.Y(n_199)
);

INVx2_ASAP7_75t_L g200 ( 
.A(n_59),
.Y(n_200)
);

CKINVDCx5p33_ASAP7_75t_R g201 ( 
.A(n_58),
.Y(n_201)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_132),
.Y(n_202)
);

CKINVDCx5p33_ASAP7_75t_R g203 ( 
.A(n_58),
.Y(n_203)
);

CKINVDCx20_ASAP7_75t_R g204 ( 
.A(n_136),
.Y(n_204)
);

CKINVDCx5p33_ASAP7_75t_R g205 ( 
.A(n_62),
.Y(n_205)
);

CKINVDCx20_ASAP7_75t_R g206 ( 
.A(n_4),
.Y(n_206)
);

CKINVDCx5p33_ASAP7_75t_R g207 ( 
.A(n_103),
.Y(n_207)
);

CKINVDCx20_ASAP7_75t_R g208 ( 
.A(n_111),
.Y(n_208)
);

CKINVDCx5p33_ASAP7_75t_R g209 ( 
.A(n_152),
.Y(n_209)
);

CKINVDCx14_ASAP7_75t_R g210 ( 
.A(n_95),
.Y(n_210)
);

CKINVDCx5p33_ASAP7_75t_R g211 ( 
.A(n_26),
.Y(n_211)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_133),
.Y(n_212)
);

CKINVDCx5p33_ASAP7_75t_R g213 ( 
.A(n_115),
.Y(n_213)
);

CKINVDCx5p33_ASAP7_75t_R g214 ( 
.A(n_48),
.Y(n_214)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_45),
.Y(n_215)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_163),
.Y(n_216)
);

CKINVDCx5p33_ASAP7_75t_R g217 ( 
.A(n_151),
.Y(n_217)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_114),
.Y(n_218)
);

CKINVDCx5p33_ASAP7_75t_R g219 ( 
.A(n_168),
.Y(n_219)
);

CKINVDCx20_ASAP7_75t_R g220 ( 
.A(n_173),
.Y(n_220)
);

CKINVDCx5p33_ASAP7_75t_R g221 ( 
.A(n_79),
.Y(n_221)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_13),
.Y(n_222)
);

CKINVDCx5p33_ASAP7_75t_R g223 ( 
.A(n_47),
.Y(n_223)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_33),
.Y(n_224)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_14),
.Y(n_225)
);

CKINVDCx5p33_ASAP7_75t_R g226 ( 
.A(n_75),
.Y(n_226)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_135),
.Y(n_227)
);

CKINVDCx5p33_ASAP7_75t_R g228 ( 
.A(n_17),
.Y(n_228)
);

CKINVDCx5p33_ASAP7_75t_R g229 ( 
.A(n_134),
.Y(n_229)
);

CKINVDCx20_ASAP7_75t_R g230 ( 
.A(n_52),
.Y(n_230)
);

CKINVDCx5p33_ASAP7_75t_R g231 ( 
.A(n_65),
.Y(n_231)
);

INVx2_ASAP7_75t_L g232 ( 
.A(n_74),
.Y(n_232)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_29),
.Y(n_233)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_76),
.Y(n_234)
);

INVx2_ASAP7_75t_SL g235 ( 
.A(n_137),
.Y(n_235)
);

CKINVDCx20_ASAP7_75t_R g236 ( 
.A(n_169),
.Y(n_236)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_155),
.Y(n_237)
);

CKINVDCx5p33_ASAP7_75t_R g238 ( 
.A(n_124),
.Y(n_238)
);

CKINVDCx5p33_ASAP7_75t_R g239 ( 
.A(n_17),
.Y(n_239)
);

CKINVDCx20_ASAP7_75t_R g240 ( 
.A(n_82),
.Y(n_240)
);

CKINVDCx16_ASAP7_75t_R g241 ( 
.A(n_159),
.Y(n_241)
);

CKINVDCx5p33_ASAP7_75t_R g242 ( 
.A(n_40),
.Y(n_242)
);

CKINVDCx5p33_ASAP7_75t_R g243 ( 
.A(n_157),
.Y(n_243)
);

CKINVDCx5p33_ASAP7_75t_R g244 ( 
.A(n_166),
.Y(n_244)
);

CKINVDCx5p33_ASAP7_75t_R g245 ( 
.A(n_4),
.Y(n_245)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_130),
.Y(n_246)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_52),
.Y(n_247)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_2),
.Y(n_248)
);

CKINVDCx5p33_ASAP7_75t_R g249 ( 
.A(n_7),
.Y(n_249)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_147),
.Y(n_250)
);

CKINVDCx5p33_ASAP7_75t_R g251 ( 
.A(n_171),
.Y(n_251)
);

INVx2_ASAP7_75t_L g252 ( 
.A(n_61),
.Y(n_252)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_146),
.Y(n_253)
);

CKINVDCx5p33_ASAP7_75t_R g254 ( 
.A(n_49),
.Y(n_254)
);

CKINVDCx5p33_ASAP7_75t_R g255 ( 
.A(n_34),
.Y(n_255)
);

CKINVDCx5p33_ASAP7_75t_R g256 ( 
.A(n_42),
.Y(n_256)
);

CKINVDCx5p33_ASAP7_75t_R g257 ( 
.A(n_56),
.Y(n_257)
);

CKINVDCx20_ASAP7_75t_R g258 ( 
.A(n_3),
.Y(n_258)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_106),
.Y(n_259)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_38),
.Y(n_260)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_66),
.Y(n_261)
);

BUFx6f_ASAP7_75t_L g262 ( 
.A(n_20),
.Y(n_262)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_40),
.Y(n_263)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_120),
.Y(n_264)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_119),
.Y(n_265)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_162),
.Y(n_266)
);

CKINVDCx5p33_ASAP7_75t_R g267 ( 
.A(n_109),
.Y(n_267)
);

CKINVDCx5p33_ASAP7_75t_R g268 ( 
.A(n_28),
.Y(n_268)
);

BUFx5_ASAP7_75t_L g269 ( 
.A(n_112),
.Y(n_269)
);

CKINVDCx5p33_ASAP7_75t_R g270 ( 
.A(n_36),
.Y(n_270)
);

CKINVDCx5p33_ASAP7_75t_R g271 ( 
.A(n_80),
.Y(n_271)
);

BUFx10_ASAP7_75t_L g272 ( 
.A(n_37),
.Y(n_272)
);

CKINVDCx5p33_ASAP7_75t_R g273 ( 
.A(n_131),
.Y(n_273)
);

CKINVDCx5p33_ASAP7_75t_R g274 ( 
.A(n_144),
.Y(n_274)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_60),
.Y(n_275)
);

CKINVDCx16_ASAP7_75t_R g276 ( 
.A(n_16),
.Y(n_276)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_14),
.Y(n_277)
);

CKINVDCx5p33_ASAP7_75t_R g278 ( 
.A(n_29),
.Y(n_278)
);

CKINVDCx5p33_ASAP7_75t_R g279 ( 
.A(n_20),
.Y(n_279)
);

CKINVDCx5p33_ASAP7_75t_R g280 ( 
.A(n_61),
.Y(n_280)
);

INVxp67_ASAP7_75t_L g281 ( 
.A(n_164),
.Y(n_281)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_128),
.Y(n_282)
);

BUFx10_ASAP7_75t_L g283 ( 
.A(n_68),
.Y(n_283)
);

INVx2_ASAP7_75t_L g284 ( 
.A(n_55),
.Y(n_284)
);

CKINVDCx5p33_ASAP7_75t_R g285 ( 
.A(n_167),
.Y(n_285)
);

BUFx5_ASAP7_75t_L g286 ( 
.A(n_150),
.Y(n_286)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_145),
.Y(n_287)
);

CKINVDCx5p33_ASAP7_75t_R g288 ( 
.A(n_138),
.Y(n_288)
);

CKINVDCx5p33_ASAP7_75t_R g289 ( 
.A(n_16),
.Y(n_289)
);

INVx2_ASAP7_75t_L g290 ( 
.A(n_143),
.Y(n_290)
);

INVx1_ASAP7_75t_SL g291 ( 
.A(n_21),
.Y(n_291)
);

CKINVDCx5p33_ASAP7_75t_R g292 ( 
.A(n_127),
.Y(n_292)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_101),
.Y(n_293)
);

CKINVDCx20_ASAP7_75t_R g294 ( 
.A(n_56),
.Y(n_294)
);

CKINVDCx5p33_ASAP7_75t_R g295 ( 
.A(n_118),
.Y(n_295)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_10),
.Y(n_296)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_0),
.Y(n_297)
);

CKINVDCx5p33_ASAP7_75t_R g298 ( 
.A(n_45),
.Y(n_298)
);

INVx1_ASAP7_75t_SL g299 ( 
.A(n_49),
.Y(n_299)
);

CKINVDCx5p33_ASAP7_75t_R g300 ( 
.A(n_77),
.Y(n_300)
);

CKINVDCx5p33_ASAP7_75t_R g301 ( 
.A(n_117),
.Y(n_301)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_43),
.Y(n_302)
);

BUFx3_ASAP7_75t_L g303 ( 
.A(n_25),
.Y(n_303)
);

CKINVDCx5p33_ASAP7_75t_R g304 ( 
.A(n_18),
.Y(n_304)
);

CKINVDCx5p33_ASAP7_75t_R g305 ( 
.A(n_60),
.Y(n_305)
);

CKINVDCx5p33_ASAP7_75t_R g306 ( 
.A(n_63),
.Y(n_306)
);

INVx1_ASAP7_75t_SL g307 ( 
.A(n_1),
.Y(n_307)
);

BUFx2_ASAP7_75t_R g308 ( 
.A(n_5),
.Y(n_308)
);

CKINVDCx5p33_ASAP7_75t_R g309 ( 
.A(n_98),
.Y(n_309)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_100),
.Y(n_310)
);

CKINVDCx20_ASAP7_75t_R g311 ( 
.A(n_50),
.Y(n_311)
);

INVx1_ASAP7_75t_SL g312 ( 
.A(n_62),
.Y(n_312)
);

INVx2_ASAP7_75t_L g313 ( 
.A(n_9),
.Y(n_313)
);

CKINVDCx5p33_ASAP7_75t_R g314 ( 
.A(n_83),
.Y(n_314)
);

CKINVDCx5p33_ASAP7_75t_R g315 ( 
.A(n_142),
.Y(n_315)
);

CKINVDCx5p33_ASAP7_75t_R g316 ( 
.A(n_36),
.Y(n_316)
);

CKINVDCx5p33_ASAP7_75t_R g317 ( 
.A(n_63),
.Y(n_317)
);

CKINVDCx5p33_ASAP7_75t_R g318 ( 
.A(n_105),
.Y(n_318)
);

BUFx6f_ASAP7_75t_L g319 ( 
.A(n_125),
.Y(n_319)
);

HB1xp67_ASAP7_75t_L g320 ( 
.A(n_39),
.Y(n_320)
);

CKINVDCx5p33_ASAP7_75t_R g321 ( 
.A(n_72),
.Y(n_321)
);

CKINVDCx5p33_ASAP7_75t_R g322 ( 
.A(n_86),
.Y(n_322)
);

CKINVDCx5p33_ASAP7_75t_R g323 ( 
.A(n_122),
.Y(n_323)
);

CKINVDCx5p33_ASAP7_75t_R g324 ( 
.A(n_37),
.Y(n_324)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_12),
.Y(n_325)
);

CKINVDCx5p33_ASAP7_75t_R g326 ( 
.A(n_10),
.Y(n_326)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_73),
.Y(n_327)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_24),
.Y(n_328)
);

BUFx5_ASAP7_75t_L g329 ( 
.A(n_156),
.Y(n_329)
);

INVx2_ASAP7_75t_L g330 ( 
.A(n_148),
.Y(n_330)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_15),
.Y(n_331)
);

CKINVDCx5p33_ASAP7_75t_R g332 ( 
.A(n_19),
.Y(n_332)
);

INVx2_ASAP7_75t_L g333 ( 
.A(n_41),
.Y(n_333)
);

CKINVDCx5p33_ASAP7_75t_R g334 ( 
.A(n_31),
.Y(n_334)
);

INVx2_ASAP7_75t_L g335 ( 
.A(n_0),
.Y(n_335)
);

CKINVDCx5p33_ASAP7_75t_R g336 ( 
.A(n_51),
.Y(n_336)
);

CKINVDCx5p33_ASAP7_75t_R g337 ( 
.A(n_94),
.Y(n_337)
);

INVx1_ASAP7_75t_L g338 ( 
.A(n_153),
.Y(n_338)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_85),
.Y(n_339)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_129),
.Y(n_340)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_11),
.Y(n_341)
);

CKINVDCx5p33_ASAP7_75t_R g342 ( 
.A(n_26),
.Y(n_342)
);

CKINVDCx5p33_ASAP7_75t_R g343 ( 
.A(n_24),
.Y(n_343)
);

CKINVDCx5p33_ASAP7_75t_R g344 ( 
.A(n_47),
.Y(n_344)
);

BUFx2_ASAP7_75t_SL g345 ( 
.A(n_87),
.Y(n_345)
);

CKINVDCx5p33_ASAP7_75t_R g346 ( 
.A(n_31),
.Y(n_346)
);

CKINVDCx5p33_ASAP7_75t_R g347 ( 
.A(n_6),
.Y(n_347)
);

CKINVDCx5p33_ASAP7_75t_R g348 ( 
.A(n_9),
.Y(n_348)
);

CKINVDCx5p33_ASAP7_75t_R g349 ( 
.A(n_176),
.Y(n_349)
);

CKINVDCx5p33_ASAP7_75t_R g350 ( 
.A(n_179),
.Y(n_350)
);

INVx1_ASAP7_75t_L g351 ( 
.A(n_189),
.Y(n_351)
);

INVx1_ASAP7_75t_L g352 ( 
.A(n_189),
.Y(n_352)
);

INVxp67_ASAP7_75t_L g353 ( 
.A(n_320),
.Y(n_353)
);

CKINVDCx5p33_ASAP7_75t_R g354 ( 
.A(n_207),
.Y(n_354)
);

INVxp67_ASAP7_75t_L g355 ( 
.A(n_272),
.Y(n_355)
);

CKINVDCx20_ASAP7_75t_R g356 ( 
.A(n_183),
.Y(n_356)
);

INVx1_ASAP7_75t_L g357 ( 
.A(n_189),
.Y(n_357)
);

CKINVDCx5p33_ASAP7_75t_R g358 ( 
.A(n_209),
.Y(n_358)
);

CKINVDCx20_ASAP7_75t_R g359 ( 
.A(n_183),
.Y(n_359)
);

INVx1_ASAP7_75t_L g360 ( 
.A(n_189),
.Y(n_360)
);

CKINVDCx16_ASAP7_75t_R g361 ( 
.A(n_276),
.Y(n_361)
);

INVx2_ASAP7_75t_L g362 ( 
.A(n_189),
.Y(n_362)
);

CKINVDCx5p33_ASAP7_75t_R g363 ( 
.A(n_213),
.Y(n_363)
);

CKINVDCx16_ASAP7_75t_R g364 ( 
.A(n_241),
.Y(n_364)
);

INVx1_ASAP7_75t_L g365 ( 
.A(n_189),
.Y(n_365)
);

INVx1_ASAP7_75t_L g366 ( 
.A(n_189),
.Y(n_366)
);

INVx1_ASAP7_75t_L g367 ( 
.A(n_262),
.Y(n_367)
);

HB1xp67_ASAP7_75t_L g368 ( 
.A(n_191),
.Y(n_368)
);

CKINVDCx20_ASAP7_75t_R g369 ( 
.A(n_184),
.Y(n_369)
);

INVxp67_ASAP7_75t_L g370 ( 
.A(n_272),
.Y(n_370)
);

CKINVDCx20_ASAP7_75t_R g371 ( 
.A(n_184),
.Y(n_371)
);

CKINVDCx5p33_ASAP7_75t_R g372 ( 
.A(n_217),
.Y(n_372)
);

NOR2xp67_ASAP7_75t_L g373 ( 
.A(n_199),
.B(n_1),
.Y(n_373)
);

CKINVDCx5p33_ASAP7_75t_R g374 ( 
.A(n_219),
.Y(n_374)
);

INVx1_ASAP7_75t_L g375 ( 
.A(n_262),
.Y(n_375)
);

CKINVDCx20_ASAP7_75t_R g376 ( 
.A(n_204),
.Y(n_376)
);

INVx1_ASAP7_75t_L g377 ( 
.A(n_262),
.Y(n_377)
);

INVx1_ASAP7_75t_L g378 ( 
.A(n_262),
.Y(n_378)
);

CKINVDCx5p33_ASAP7_75t_R g379 ( 
.A(n_221),
.Y(n_379)
);

CKINVDCx5p33_ASAP7_75t_R g380 ( 
.A(n_226),
.Y(n_380)
);

INVx1_ASAP7_75t_L g381 ( 
.A(n_262),
.Y(n_381)
);

CKINVDCx20_ASAP7_75t_R g382 ( 
.A(n_204),
.Y(n_382)
);

CKINVDCx20_ASAP7_75t_R g383 ( 
.A(n_208),
.Y(n_383)
);

CKINVDCx20_ASAP7_75t_R g384 ( 
.A(n_208),
.Y(n_384)
);

INVx1_ASAP7_75t_L g385 ( 
.A(n_199),
.Y(n_385)
);

INVx1_ASAP7_75t_L g386 ( 
.A(n_200),
.Y(n_386)
);

NOR2xp67_ASAP7_75t_L g387 ( 
.A(n_200),
.B(n_3),
.Y(n_387)
);

INVx1_ASAP7_75t_L g388 ( 
.A(n_252),
.Y(n_388)
);

INVx2_ASAP7_75t_L g389 ( 
.A(n_269),
.Y(n_389)
);

INVx1_ASAP7_75t_L g390 ( 
.A(n_252),
.Y(n_390)
);

NOR2xp67_ASAP7_75t_L g391 ( 
.A(n_284),
.B(n_5),
.Y(n_391)
);

INVx1_ASAP7_75t_L g392 ( 
.A(n_284),
.Y(n_392)
);

INVx1_ASAP7_75t_L g393 ( 
.A(n_313),
.Y(n_393)
);

INVx1_ASAP7_75t_L g394 ( 
.A(n_313),
.Y(n_394)
);

INVx2_ASAP7_75t_L g395 ( 
.A(n_269),
.Y(n_395)
);

INVxp67_ASAP7_75t_SL g396 ( 
.A(n_281),
.Y(n_396)
);

INVx1_ASAP7_75t_L g397 ( 
.A(n_333),
.Y(n_397)
);

INVxp67_ASAP7_75t_L g398 ( 
.A(n_272),
.Y(n_398)
);

INVx1_ASAP7_75t_L g399 ( 
.A(n_333),
.Y(n_399)
);

CKINVDCx5p33_ASAP7_75t_R g400 ( 
.A(n_229),
.Y(n_400)
);

CKINVDCx5p33_ASAP7_75t_R g401 ( 
.A(n_231),
.Y(n_401)
);

CKINVDCx5p33_ASAP7_75t_R g402 ( 
.A(n_238),
.Y(n_402)
);

CKINVDCx5p33_ASAP7_75t_R g403 ( 
.A(n_243),
.Y(n_403)
);

INVx1_ASAP7_75t_L g404 ( 
.A(n_335),
.Y(n_404)
);

INVxp67_ASAP7_75t_SL g405 ( 
.A(n_303),
.Y(n_405)
);

INVx1_ASAP7_75t_L g406 ( 
.A(n_335),
.Y(n_406)
);

CKINVDCx5p33_ASAP7_75t_R g407 ( 
.A(n_244),
.Y(n_407)
);

INVxp67_ASAP7_75t_SL g408 ( 
.A(n_303),
.Y(n_408)
);

CKINVDCx5p33_ASAP7_75t_R g409 ( 
.A(n_251),
.Y(n_409)
);

INVx1_ASAP7_75t_L g410 ( 
.A(n_215),
.Y(n_410)
);

INVxp67_ASAP7_75t_SL g411 ( 
.A(n_182),
.Y(n_411)
);

INVx1_ASAP7_75t_L g412 ( 
.A(n_222),
.Y(n_412)
);

CKINVDCx5p33_ASAP7_75t_R g413 ( 
.A(n_267),
.Y(n_413)
);

CKINVDCx5p33_ASAP7_75t_R g414 ( 
.A(n_271),
.Y(n_414)
);

CKINVDCx20_ASAP7_75t_R g415 ( 
.A(n_220),
.Y(n_415)
);

INVx1_ASAP7_75t_L g416 ( 
.A(n_224),
.Y(n_416)
);

INVx1_ASAP7_75t_L g417 ( 
.A(n_225),
.Y(n_417)
);

CKINVDCx20_ASAP7_75t_R g418 ( 
.A(n_220),
.Y(n_418)
);

CKINVDCx20_ASAP7_75t_R g419 ( 
.A(n_236),
.Y(n_419)
);

CKINVDCx5p33_ASAP7_75t_R g420 ( 
.A(n_273),
.Y(n_420)
);

INVx1_ASAP7_75t_L g421 ( 
.A(n_233),
.Y(n_421)
);

INVx2_ASAP7_75t_L g422 ( 
.A(n_269),
.Y(n_422)
);

CKINVDCx20_ASAP7_75t_R g423 ( 
.A(n_236),
.Y(n_423)
);

CKINVDCx20_ASAP7_75t_R g424 ( 
.A(n_240),
.Y(n_424)
);

INVxp67_ASAP7_75t_SL g425 ( 
.A(n_185),
.Y(n_425)
);

INVx1_ASAP7_75t_L g426 ( 
.A(n_247),
.Y(n_426)
);

NOR2xp33_ASAP7_75t_L g427 ( 
.A(n_235),
.B(n_6),
.Y(n_427)
);

CKINVDCx5p33_ASAP7_75t_R g428 ( 
.A(n_274),
.Y(n_428)
);

INVx3_ASAP7_75t_L g429 ( 
.A(n_177),
.Y(n_429)
);

INVx1_ASAP7_75t_L g430 ( 
.A(n_248),
.Y(n_430)
);

INVx2_ASAP7_75t_L g431 ( 
.A(n_269),
.Y(n_431)
);

CKINVDCx20_ASAP7_75t_R g432 ( 
.A(n_240),
.Y(n_432)
);

CKINVDCx5p33_ASAP7_75t_R g433 ( 
.A(n_285),
.Y(n_433)
);

NOR2xp67_ASAP7_75t_L g434 ( 
.A(n_260),
.B(n_7),
.Y(n_434)
);

INVx1_ASAP7_75t_L g435 ( 
.A(n_263),
.Y(n_435)
);

INVx1_ASAP7_75t_L g436 ( 
.A(n_275),
.Y(n_436)
);

INVx3_ASAP7_75t_L g437 ( 
.A(n_362),
.Y(n_437)
);

INVx2_ASAP7_75t_L g438 ( 
.A(n_362),
.Y(n_438)
);

INVx2_ASAP7_75t_L g439 ( 
.A(n_351),
.Y(n_439)
);

NAND2xp5_ASAP7_75t_L g440 ( 
.A(n_411),
.B(n_210),
.Y(n_440)
);

NOR2xp33_ASAP7_75t_L g441 ( 
.A(n_427),
.B(n_235),
.Y(n_441)
);

AND2x4_ASAP7_75t_L g442 ( 
.A(n_429),
.B(n_188),
.Y(n_442)
);

INVx1_ASAP7_75t_L g443 ( 
.A(n_367),
.Y(n_443)
);

INVx1_ASAP7_75t_L g444 ( 
.A(n_367),
.Y(n_444)
);

NAND2xp5_ASAP7_75t_L g445 ( 
.A(n_425),
.B(n_175),
.Y(n_445)
);

BUFx6f_ASAP7_75t_L g446 ( 
.A(n_389),
.Y(n_446)
);

BUFx8_ASAP7_75t_L g447 ( 
.A(n_410),
.Y(n_447)
);

INVx1_ASAP7_75t_L g448 ( 
.A(n_375),
.Y(n_448)
);

INVx1_ASAP7_75t_L g449 ( 
.A(n_375),
.Y(n_449)
);

AND2x2_ASAP7_75t_L g450 ( 
.A(n_405),
.B(n_188),
.Y(n_450)
);

AND3x2_ASAP7_75t_L g451 ( 
.A(n_355),
.B(n_290),
.C(n_232),
.Y(n_451)
);

INVx2_ASAP7_75t_L g452 ( 
.A(n_351),
.Y(n_452)
);

OA21x2_ASAP7_75t_L g453 ( 
.A1(n_352),
.A2(n_360),
.B(n_357),
.Y(n_453)
);

INVx1_ASAP7_75t_L g454 ( 
.A(n_377),
.Y(n_454)
);

INVx4_ASAP7_75t_L g455 ( 
.A(n_429),
.Y(n_455)
);

OA21x2_ASAP7_75t_L g456 ( 
.A1(n_352),
.A2(n_296),
.B(n_277),
.Y(n_456)
);

INVx2_ASAP7_75t_L g457 ( 
.A(n_357),
.Y(n_457)
);

BUFx6f_ASAP7_75t_L g458 ( 
.A(n_389),
.Y(n_458)
);

INVx1_ASAP7_75t_L g459 ( 
.A(n_377),
.Y(n_459)
);

INVx2_ASAP7_75t_L g460 ( 
.A(n_360),
.Y(n_460)
);

INVx2_ASAP7_75t_L g461 ( 
.A(n_365),
.Y(n_461)
);

HB1xp67_ASAP7_75t_L g462 ( 
.A(n_368),
.Y(n_462)
);

INVx1_ASAP7_75t_L g463 ( 
.A(n_378),
.Y(n_463)
);

INVxp33_ASAP7_75t_SL g464 ( 
.A(n_349),
.Y(n_464)
);

NAND2xp5_ASAP7_75t_L g465 ( 
.A(n_378),
.B(n_175),
.Y(n_465)
);

INVx2_ASAP7_75t_L g466 ( 
.A(n_365),
.Y(n_466)
);

INVx2_ASAP7_75t_L g467 ( 
.A(n_366),
.Y(n_467)
);

INVx1_ASAP7_75t_L g468 ( 
.A(n_381),
.Y(n_468)
);

INVx2_ASAP7_75t_L g469 ( 
.A(n_366),
.Y(n_469)
);

AND2x4_ASAP7_75t_L g470 ( 
.A(n_429),
.B(n_232),
.Y(n_470)
);

INVx3_ASAP7_75t_L g471 ( 
.A(n_429),
.Y(n_471)
);

INVx1_ASAP7_75t_L g472 ( 
.A(n_381),
.Y(n_472)
);

INVx1_ASAP7_75t_L g473 ( 
.A(n_395),
.Y(n_473)
);

AND2x2_ASAP7_75t_L g474 ( 
.A(n_408),
.B(n_290),
.Y(n_474)
);

AND2x6_ASAP7_75t_L g475 ( 
.A(n_395),
.B(n_330),
.Y(n_475)
);

INVx2_ASAP7_75t_L g476 ( 
.A(n_422),
.Y(n_476)
);

INVx2_ASAP7_75t_L g477 ( 
.A(n_422),
.Y(n_477)
);

INVx1_ASAP7_75t_L g478 ( 
.A(n_431),
.Y(n_478)
);

NOR2xp33_ASAP7_75t_L g479 ( 
.A(n_396),
.B(n_178),
.Y(n_479)
);

INVx3_ASAP7_75t_L g480 ( 
.A(n_431),
.Y(n_480)
);

BUFx6f_ASAP7_75t_L g481 ( 
.A(n_385),
.Y(n_481)
);

NAND2xp5_ASAP7_75t_L g482 ( 
.A(n_410),
.B(n_195),
.Y(n_482)
);

BUFx6f_ASAP7_75t_L g483 ( 
.A(n_385),
.Y(n_483)
);

INVx2_ASAP7_75t_L g484 ( 
.A(n_386),
.Y(n_484)
);

INVx1_ASAP7_75t_L g485 ( 
.A(n_386),
.Y(n_485)
);

AND2x2_ASAP7_75t_L g486 ( 
.A(n_388),
.B(n_330),
.Y(n_486)
);

CKINVDCx16_ASAP7_75t_R g487 ( 
.A(n_361),
.Y(n_487)
);

BUFx3_ASAP7_75t_L g488 ( 
.A(n_388),
.Y(n_488)
);

INVx1_ASAP7_75t_L g489 ( 
.A(n_390),
.Y(n_489)
);

INVx1_ASAP7_75t_L g490 ( 
.A(n_390),
.Y(n_490)
);

AND2x2_ASAP7_75t_L g491 ( 
.A(n_392),
.B(n_190),
.Y(n_491)
);

INVxp67_ASAP7_75t_L g492 ( 
.A(n_412),
.Y(n_492)
);

INVx2_ASAP7_75t_L g493 ( 
.A(n_392),
.Y(n_493)
);

INVx1_ASAP7_75t_L g494 ( 
.A(n_393),
.Y(n_494)
);

HB1xp67_ASAP7_75t_L g495 ( 
.A(n_370),
.Y(n_495)
);

INVx3_ASAP7_75t_L g496 ( 
.A(n_393),
.Y(n_496)
);

INVx1_ASAP7_75t_L g497 ( 
.A(n_394),
.Y(n_497)
);

INVx1_ASAP7_75t_L g498 ( 
.A(n_394),
.Y(n_498)
);

INVx1_ASAP7_75t_L g499 ( 
.A(n_397),
.Y(n_499)
);

AOI22xp5_ASAP7_75t_L g500 ( 
.A1(n_353),
.A2(n_230),
.B1(n_193),
.B2(n_206),
.Y(n_500)
);

INVx1_ASAP7_75t_L g501 ( 
.A(n_397),
.Y(n_501)
);

INVx2_ASAP7_75t_L g502 ( 
.A(n_399),
.Y(n_502)
);

INVx1_ASAP7_75t_SL g503 ( 
.A(n_356),
.Y(n_503)
);

CKINVDCx8_ASAP7_75t_R g504 ( 
.A(n_361),
.Y(n_504)
);

INVx3_ASAP7_75t_L g505 ( 
.A(n_399),
.Y(n_505)
);

AND2x2_ASAP7_75t_L g506 ( 
.A(n_404),
.B(n_192),
.Y(n_506)
);

BUFx2_ASAP7_75t_L g507 ( 
.A(n_398),
.Y(n_507)
);

OA21x2_ASAP7_75t_L g508 ( 
.A1(n_404),
.A2(n_406),
.B(n_302),
.Y(n_508)
);

HB1xp67_ASAP7_75t_L g509 ( 
.A(n_434),
.Y(n_509)
);

HB1xp67_ASAP7_75t_L g510 ( 
.A(n_373),
.Y(n_510)
);

INVxp67_ASAP7_75t_L g511 ( 
.A(n_412),
.Y(n_511)
);

NOR2xp33_ASAP7_75t_L g512 ( 
.A(n_350),
.B(n_181),
.Y(n_512)
);

INVx2_ASAP7_75t_L g513 ( 
.A(n_406),
.Y(n_513)
);

AND2x4_ASAP7_75t_L g514 ( 
.A(n_387),
.B(n_177),
.Y(n_514)
);

INVx1_ASAP7_75t_L g515 ( 
.A(n_453),
.Y(n_515)
);

XOR2xp5_ASAP7_75t_L g516 ( 
.A(n_500),
.B(n_359),
.Y(n_516)
);

BUFx3_ASAP7_75t_L g517 ( 
.A(n_453),
.Y(n_517)
);

INVx4_ASAP7_75t_L g518 ( 
.A(n_446),
.Y(n_518)
);

INVx1_ASAP7_75t_L g519 ( 
.A(n_453),
.Y(n_519)
);

NAND2xp5_ASAP7_75t_SL g520 ( 
.A(n_479),
.B(n_364),
.Y(n_520)
);

BUFx8_ASAP7_75t_SL g521 ( 
.A(n_507),
.Y(n_521)
);

NOR2xp33_ASAP7_75t_L g522 ( 
.A(n_441),
.B(n_354),
.Y(n_522)
);

NOR2xp33_ASAP7_75t_L g523 ( 
.A(n_441),
.B(n_358),
.Y(n_523)
);

INVx1_ASAP7_75t_L g524 ( 
.A(n_453),
.Y(n_524)
);

BUFx6f_ASAP7_75t_SL g525 ( 
.A(n_514),
.Y(n_525)
);

INVx3_ASAP7_75t_L g526 ( 
.A(n_446),
.Y(n_526)
);

INVx1_ASAP7_75t_L g527 ( 
.A(n_453),
.Y(n_527)
);

NOR2xp33_ASAP7_75t_L g528 ( 
.A(n_512),
.B(n_363),
.Y(n_528)
);

INVx1_ASAP7_75t_L g529 ( 
.A(n_453),
.Y(n_529)
);

INVx1_ASAP7_75t_L g530 ( 
.A(n_453),
.Y(n_530)
);

INVx4_ASAP7_75t_L g531 ( 
.A(n_446),
.Y(n_531)
);

INVx1_ASAP7_75t_L g532 ( 
.A(n_508),
.Y(n_532)
);

INVx1_ASAP7_75t_L g533 ( 
.A(n_508),
.Y(n_533)
);

BUFx4f_ASAP7_75t_L g534 ( 
.A(n_456),
.Y(n_534)
);

NAND2xp5_ASAP7_75t_SL g535 ( 
.A(n_479),
.B(n_364),
.Y(n_535)
);

NOR2xp33_ASAP7_75t_L g536 ( 
.A(n_512),
.B(n_372),
.Y(n_536)
);

INVx1_ASAP7_75t_L g537 ( 
.A(n_508),
.Y(n_537)
);

INVx4_ASAP7_75t_L g538 ( 
.A(n_446),
.Y(n_538)
);

INVx1_ASAP7_75t_L g539 ( 
.A(n_508),
.Y(n_539)
);

BUFx6f_ASAP7_75t_L g540 ( 
.A(n_446),
.Y(n_540)
);

OAI22xp33_ASAP7_75t_L g541 ( 
.A1(n_445),
.A2(n_291),
.B1(n_299),
.B2(n_307),
.Y(n_541)
);

NOR2xp33_ASAP7_75t_L g542 ( 
.A(n_440),
.B(n_374),
.Y(n_542)
);

INVx1_ASAP7_75t_L g543 ( 
.A(n_508),
.Y(n_543)
);

AOI22xp33_ASAP7_75t_L g544 ( 
.A1(n_450),
.A2(n_391),
.B1(n_297),
.B2(n_325),
.Y(n_544)
);

INVx4_ASAP7_75t_SL g545 ( 
.A(n_475),
.Y(n_545)
);

INVx8_ASAP7_75t_L g546 ( 
.A(n_475),
.Y(n_546)
);

INVx2_ASAP7_75t_L g547 ( 
.A(n_438),
.Y(n_547)
);

INVx2_ASAP7_75t_L g548 ( 
.A(n_438),
.Y(n_548)
);

AND2x4_ASAP7_75t_L g549 ( 
.A(n_491),
.B(n_202),
.Y(n_549)
);

BUFx6f_ASAP7_75t_SL g550 ( 
.A(n_514),
.Y(n_550)
);

INVx2_ASAP7_75t_L g551 ( 
.A(n_438),
.Y(n_551)
);

AOI22xp33_ASAP7_75t_SL g552 ( 
.A1(n_487),
.A2(n_230),
.B1(n_206),
.B2(n_294),
.Y(n_552)
);

BUFx3_ASAP7_75t_L g553 ( 
.A(n_456),
.Y(n_553)
);

NAND2xp5_ASAP7_75t_SL g554 ( 
.A(n_464),
.B(n_379),
.Y(n_554)
);

NAND2xp5_ASAP7_75t_L g555 ( 
.A(n_440),
.B(n_380),
.Y(n_555)
);

AOI22xp33_ASAP7_75t_L g556 ( 
.A1(n_450),
.A2(n_328),
.B1(n_331),
.B2(n_341),
.Y(n_556)
);

INVx1_ASAP7_75t_L g557 ( 
.A(n_508),
.Y(n_557)
);

INVx4_ASAP7_75t_L g558 ( 
.A(n_446),
.Y(n_558)
);

CKINVDCx5p33_ASAP7_75t_R g559 ( 
.A(n_487),
.Y(n_559)
);

INVx1_ASAP7_75t_L g560 ( 
.A(n_508),
.Y(n_560)
);

BUFx8_ASAP7_75t_SL g561 ( 
.A(n_507),
.Y(n_561)
);

NOR2x1p5_ASAP7_75t_L g562 ( 
.A(n_482),
.B(n_191),
.Y(n_562)
);

BUFx3_ASAP7_75t_L g563 ( 
.A(n_456),
.Y(n_563)
);

INVx1_ASAP7_75t_L g564 ( 
.A(n_439),
.Y(n_564)
);

NOR2xp33_ASAP7_75t_L g565 ( 
.A(n_464),
.B(n_400),
.Y(n_565)
);

INVx2_ASAP7_75t_L g566 ( 
.A(n_438),
.Y(n_566)
);

INVx2_ASAP7_75t_L g567 ( 
.A(n_476),
.Y(n_567)
);

INVx2_ASAP7_75t_L g568 ( 
.A(n_476),
.Y(n_568)
);

INVx1_ASAP7_75t_L g569 ( 
.A(n_439),
.Y(n_569)
);

OAI22xp33_ASAP7_75t_L g570 ( 
.A1(n_445),
.A2(n_312),
.B1(n_257),
.B2(n_187),
.Y(n_570)
);

AND2x2_ASAP7_75t_L g571 ( 
.A(n_450),
.B(n_416),
.Y(n_571)
);

BUFx3_ASAP7_75t_L g572 ( 
.A(n_456),
.Y(n_572)
);

INVx2_ASAP7_75t_L g573 ( 
.A(n_476),
.Y(n_573)
);

INVx1_ASAP7_75t_L g574 ( 
.A(n_439),
.Y(n_574)
);

INVx2_ASAP7_75t_L g575 ( 
.A(n_476),
.Y(n_575)
);

INVx2_ASAP7_75t_L g576 ( 
.A(n_477),
.Y(n_576)
);

AOI22xp5_ASAP7_75t_L g577 ( 
.A1(n_500),
.A2(n_294),
.B1(n_258),
.B2(n_193),
.Y(n_577)
);

AND2x2_ASAP7_75t_L g578 ( 
.A(n_450),
.B(n_416),
.Y(n_578)
);

NAND2xp5_ASAP7_75t_SL g579 ( 
.A(n_447),
.B(n_401),
.Y(n_579)
);

INVx3_ASAP7_75t_L g580 ( 
.A(n_446),
.Y(n_580)
);

INVx3_ASAP7_75t_L g581 ( 
.A(n_446),
.Y(n_581)
);

INVx2_ASAP7_75t_L g582 ( 
.A(n_477),
.Y(n_582)
);

INVx1_ASAP7_75t_L g583 ( 
.A(n_439),
.Y(n_583)
);

AOI22xp33_ASAP7_75t_L g584 ( 
.A1(n_474),
.A2(n_345),
.B1(n_180),
.B2(n_319),
.Y(n_584)
);

INVx2_ASAP7_75t_SL g585 ( 
.A(n_447),
.Y(n_585)
);

INVx2_ASAP7_75t_L g586 ( 
.A(n_477),
.Y(n_586)
);

INVx1_ASAP7_75t_L g587 ( 
.A(n_452),
.Y(n_587)
);

INVx2_ASAP7_75t_L g588 ( 
.A(n_477),
.Y(n_588)
);

INVx1_ASAP7_75t_L g589 ( 
.A(n_452),
.Y(n_589)
);

BUFx6f_ASAP7_75t_L g590 ( 
.A(n_446),
.Y(n_590)
);

AND3x2_ASAP7_75t_L g591 ( 
.A(n_507),
.B(n_216),
.C(n_212),
.Y(n_591)
);

AOI22xp33_ASAP7_75t_L g592 ( 
.A1(n_474),
.A2(n_177),
.B1(n_180),
.B2(n_319),
.Y(n_592)
);

NAND3xp33_ASAP7_75t_L g593 ( 
.A(n_456),
.B(n_421),
.C(n_417),
.Y(n_593)
);

INVx1_ASAP7_75t_L g594 ( 
.A(n_452),
.Y(n_594)
);

INVx5_ASAP7_75t_L g595 ( 
.A(n_475),
.Y(n_595)
);

BUFx2_ASAP7_75t_L g596 ( 
.A(n_495),
.Y(n_596)
);

INVx3_ASAP7_75t_L g597 ( 
.A(n_458),
.Y(n_597)
);

INVx2_ASAP7_75t_L g598 ( 
.A(n_452),
.Y(n_598)
);

NOR2xp33_ASAP7_75t_L g599 ( 
.A(n_495),
.B(n_402),
.Y(n_599)
);

BUFx2_ASAP7_75t_L g600 ( 
.A(n_462),
.Y(n_600)
);

AND2x2_ASAP7_75t_L g601 ( 
.A(n_474),
.B(n_417),
.Y(n_601)
);

INVx1_ASAP7_75t_L g602 ( 
.A(n_457),
.Y(n_602)
);

AND2x2_ASAP7_75t_L g603 ( 
.A(n_474),
.B(n_436),
.Y(n_603)
);

AOI22xp33_ASAP7_75t_SL g604 ( 
.A1(n_487),
.A2(n_311),
.B1(n_258),
.B2(n_432),
.Y(n_604)
);

INVx2_ASAP7_75t_L g605 ( 
.A(n_457),
.Y(n_605)
);

INVx1_ASAP7_75t_L g606 ( 
.A(n_457),
.Y(n_606)
);

INVx2_ASAP7_75t_L g607 ( 
.A(n_457),
.Y(n_607)
);

INVx2_ASAP7_75t_L g608 ( 
.A(n_460),
.Y(n_608)
);

NAND2xp33_ASAP7_75t_L g609 ( 
.A(n_509),
.B(n_403),
.Y(n_609)
);

BUFx6f_ASAP7_75t_L g610 ( 
.A(n_458),
.Y(n_610)
);

NAND2xp5_ASAP7_75t_SL g611 ( 
.A(n_447),
.B(n_407),
.Y(n_611)
);

INVx5_ASAP7_75t_L g612 ( 
.A(n_475),
.Y(n_612)
);

INVx1_ASAP7_75t_L g613 ( 
.A(n_460),
.Y(n_613)
);

OR2x6_ASAP7_75t_L g614 ( 
.A(n_482),
.B(n_218),
.Y(n_614)
);

NAND2xp5_ASAP7_75t_L g615 ( 
.A(n_455),
.B(n_409),
.Y(n_615)
);

BUFx2_ASAP7_75t_L g616 ( 
.A(n_462),
.Y(n_616)
);

NAND2xp5_ASAP7_75t_SL g617 ( 
.A(n_447),
.B(n_413),
.Y(n_617)
);

AOI22xp33_ASAP7_75t_L g618 ( 
.A1(n_456),
.A2(n_177),
.B1(n_180),
.B2(n_319),
.Y(n_618)
);

CKINVDCx5p33_ASAP7_75t_R g619 ( 
.A(n_504),
.Y(n_619)
);

INVx1_ASAP7_75t_L g620 ( 
.A(n_460),
.Y(n_620)
);

BUFx3_ASAP7_75t_L g621 ( 
.A(n_456),
.Y(n_621)
);

AND2x2_ASAP7_75t_SL g622 ( 
.A(n_455),
.B(n_177),
.Y(n_622)
);

AND2x2_ASAP7_75t_L g623 ( 
.A(n_491),
.B(n_436),
.Y(n_623)
);

NOR2xp33_ASAP7_75t_L g624 ( 
.A(n_465),
.B(n_414),
.Y(n_624)
);

NAND2xp33_ASAP7_75t_L g625 ( 
.A(n_509),
.B(n_420),
.Y(n_625)
);

INVx1_ASAP7_75t_L g626 ( 
.A(n_460),
.Y(n_626)
);

CKINVDCx5p33_ASAP7_75t_R g627 ( 
.A(n_504),
.Y(n_627)
);

BUFx3_ASAP7_75t_L g628 ( 
.A(n_488),
.Y(n_628)
);

INVx2_ASAP7_75t_L g629 ( 
.A(n_461),
.Y(n_629)
);

INVx2_ASAP7_75t_L g630 ( 
.A(n_461),
.Y(n_630)
);

INVx2_ASAP7_75t_L g631 ( 
.A(n_461),
.Y(n_631)
);

AND2x2_ASAP7_75t_L g632 ( 
.A(n_491),
.B(n_421),
.Y(n_632)
);

INVx2_ASAP7_75t_L g633 ( 
.A(n_461),
.Y(n_633)
);

INVx2_ASAP7_75t_L g634 ( 
.A(n_466),
.Y(n_634)
);

CKINVDCx20_ASAP7_75t_R g635 ( 
.A(n_504),
.Y(n_635)
);

INVx1_ASAP7_75t_SL g636 ( 
.A(n_503),
.Y(n_636)
);

NOR2xp33_ASAP7_75t_L g637 ( 
.A(n_465),
.B(n_428),
.Y(n_637)
);

AOI22xp5_ASAP7_75t_L g638 ( 
.A1(n_500),
.A2(n_311),
.B1(n_196),
.B2(n_348),
.Y(n_638)
);

BUFx6f_ASAP7_75t_L g639 ( 
.A(n_458),
.Y(n_639)
);

INVx1_ASAP7_75t_L g640 ( 
.A(n_466),
.Y(n_640)
);

AND2x2_ASAP7_75t_L g641 ( 
.A(n_491),
.B(n_506),
.Y(n_641)
);

NAND2xp5_ASAP7_75t_SL g642 ( 
.A(n_447),
.B(n_433),
.Y(n_642)
);

INVx1_ASAP7_75t_L g643 ( 
.A(n_466),
.Y(n_643)
);

INVx4_ASAP7_75t_L g644 ( 
.A(n_458),
.Y(n_644)
);

AND3x2_ASAP7_75t_L g645 ( 
.A(n_510),
.B(n_234),
.C(n_227),
.Y(n_645)
);

NAND2xp5_ASAP7_75t_L g646 ( 
.A(n_455),
.B(n_288),
.Y(n_646)
);

BUFx6f_ASAP7_75t_L g647 ( 
.A(n_458),
.Y(n_647)
);

INVx2_ASAP7_75t_L g648 ( 
.A(n_466),
.Y(n_648)
);

AND3x2_ASAP7_75t_L g649 ( 
.A(n_510),
.B(n_246),
.C(n_237),
.Y(n_649)
);

INVx1_ASAP7_75t_L g650 ( 
.A(n_467),
.Y(n_650)
);

AOI22xp33_ASAP7_75t_L g651 ( 
.A1(n_506),
.A2(n_180),
.B1(n_319),
.B2(n_435),
.Y(n_651)
);

INVx2_ASAP7_75t_L g652 ( 
.A(n_467),
.Y(n_652)
);

NOR2xp33_ASAP7_75t_L g653 ( 
.A(n_492),
.B(n_369),
.Y(n_653)
);

BUFx6f_ASAP7_75t_SL g654 ( 
.A(n_514),
.Y(n_654)
);

AND2x2_ASAP7_75t_L g655 ( 
.A(n_506),
.B(n_426),
.Y(n_655)
);

NAND2xp5_ASAP7_75t_L g656 ( 
.A(n_455),
.B(n_292),
.Y(n_656)
);

NAND2xp5_ASAP7_75t_SL g657 ( 
.A(n_447),
.B(n_283),
.Y(n_657)
);

INVx1_ASAP7_75t_L g658 ( 
.A(n_467),
.Y(n_658)
);

INVx2_ASAP7_75t_L g659 ( 
.A(n_467),
.Y(n_659)
);

INVx1_ASAP7_75t_SL g660 ( 
.A(n_503),
.Y(n_660)
);

NAND2xp5_ASAP7_75t_SL g661 ( 
.A(n_504),
.B(n_283),
.Y(n_661)
);

INVx2_ASAP7_75t_L g662 ( 
.A(n_469),
.Y(n_662)
);

NAND2xp5_ASAP7_75t_L g663 ( 
.A(n_455),
.B(n_295),
.Y(n_663)
);

NAND2xp5_ASAP7_75t_L g664 ( 
.A(n_455),
.B(n_300),
.Y(n_664)
);

AOI22xp33_ASAP7_75t_L g665 ( 
.A1(n_506),
.A2(n_319),
.B1(n_180),
.B2(n_435),
.Y(n_665)
);

NAND2xp5_ASAP7_75t_SL g666 ( 
.A(n_492),
.B(n_283),
.Y(n_666)
);

INVx1_ASAP7_75t_L g667 ( 
.A(n_469),
.Y(n_667)
);

INVx2_ASAP7_75t_SL g668 ( 
.A(n_571),
.Y(n_668)
);

CKINVDCx5p33_ASAP7_75t_R g669 ( 
.A(n_559),
.Y(n_669)
);

NAND2xp5_ASAP7_75t_L g670 ( 
.A(n_624),
.B(n_469),
.Y(n_670)
);

BUFx6f_ASAP7_75t_SL g671 ( 
.A(n_614),
.Y(n_671)
);

NAND2xp5_ASAP7_75t_L g672 ( 
.A(n_637),
.B(n_469),
.Y(n_672)
);

INVx2_ASAP7_75t_L g673 ( 
.A(n_547),
.Y(n_673)
);

INVx1_ASAP7_75t_L g674 ( 
.A(n_641),
.Y(n_674)
);

AND2x4_ASAP7_75t_L g675 ( 
.A(n_641),
.B(n_511),
.Y(n_675)
);

OAI22xp33_ASAP7_75t_L g676 ( 
.A1(n_577),
.A2(n_511),
.B1(n_205),
.B2(n_198),
.Y(n_676)
);

NAND2xp5_ASAP7_75t_L g677 ( 
.A(n_522),
.B(n_514),
.Y(n_677)
);

INVx2_ASAP7_75t_SL g678 ( 
.A(n_571),
.Y(n_678)
);

O2A1O1Ixp33_ASAP7_75t_L g679 ( 
.A1(n_515),
.A2(n_486),
.B(n_426),
.C(n_430),
.Y(n_679)
);

BUFx6f_ASAP7_75t_L g680 ( 
.A(n_517),
.Y(n_680)
);

NAND2xp5_ASAP7_75t_L g681 ( 
.A(n_523),
.B(n_542),
.Y(n_681)
);

INVx1_ASAP7_75t_L g682 ( 
.A(n_623),
.Y(n_682)
);

AND2x6_ASAP7_75t_SL g683 ( 
.A(n_528),
.B(n_308),
.Y(n_683)
);

AOI22xp33_ASAP7_75t_L g684 ( 
.A1(n_553),
.A2(n_486),
.B1(n_514),
.B2(n_470),
.Y(n_684)
);

OR2x6_ASAP7_75t_L g685 ( 
.A(n_600),
.B(n_430),
.Y(n_685)
);

NOR2xp33_ASAP7_75t_L g686 ( 
.A(n_536),
.B(n_195),
.Y(n_686)
);

NAND2xp5_ASAP7_75t_SL g687 ( 
.A(n_622),
.B(n_514),
.Y(n_687)
);

INVx1_ASAP7_75t_L g688 ( 
.A(n_623),
.Y(n_688)
);

A2O1A1Ixp33_ASAP7_75t_L g689 ( 
.A1(n_534),
.A2(n_442),
.B(n_470),
.C(n_339),
.Y(n_689)
);

NAND2xp5_ASAP7_75t_L g690 ( 
.A(n_515),
.B(n_458),
.Y(n_690)
);

NAND2xp5_ASAP7_75t_SL g691 ( 
.A(n_622),
.B(n_534),
.Y(n_691)
);

NAND2xp5_ASAP7_75t_L g692 ( 
.A(n_519),
.B(n_458),
.Y(n_692)
);

NAND2xp5_ASAP7_75t_L g693 ( 
.A(n_519),
.B(n_524),
.Y(n_693)
);

AOI21xp5_ASAP7_75t_L g694 ( 
.A1(n_534),
.A2(n_478),
.B(n_473),
.Y(n_694)
);

INVx2_ASAP7_75t_SL g695 ( 
.A(n_578),
.Y(n_695)
);

NAND2xp5_ASAP7_75t_SL g696 ( 
.A(n_622),
.B(n_458),
.Y(n_696)
);

OAI22xp5_ASAP7_75t_L g697 ( 
.A1(n_584),
.A2(n_282),
.B1(n_310),
.B2(n_293),
.Y(n_697)
);

NAND2xp5_ASAP7_75t_SL g698 ( 
.A(n_517),
.B(n_458),
.Y(n_698)
);

NAND2x1_ASAP7_75t_L g699 ( 
.A(n_524),
.B(n_471),
.Y(n_699)
);

CKINVDCx5p33_ASAP7_75t_R g700 ( 
.A(n_559),
.Y(n_700)
);

INVx1_ASAP7_75t_L g701 ( 
.A(n_632),
.Y(n_701)
);

NAND2xp5_ASAP7_75t_SL g702 ( 
.A(n_517),
.B(n_269),
.Y(n_702)
);

INVx1_ASAP7_75t_L g703 ( 
.A(n_632),
.Y(n_703)
);

NAND2xp5_ASAP7_75t_SL g704 ( 
.A(n_553),
.B(n_269),
.Y(n_704)
);

NAND2x1p5_ASAP7_75t_L g705 ( 
.A(n_553),
.B(n_250),
.Y(n_705)
);

AND2x2_ASAP7_75t_L g706 ( 
.A(n_578),
.B(n_601),
.Y(n_706)
);

NAND2xp5_ASAP7_75t_L g707 ( 
.A(n_527),
.B(n_442),
.Y(n_707)
);

NOR2xp33_ASAP7_75t_L g708 ( 
.A(n_555),
.B(n_186),
.Y(n_708)
);

INVx2_ASAP7_75t_L g709 ( 
.A(n_547),
.Y(n_709)
);

NAND2xp5_ASAP7_75t_L g710 ( 
.A(n_527),
.B(n_442),
.Y(n_710)
);

NAND2x1_ASAP7_75t_L g711 ( 
.A(n_529),
.B(n_471),
.Y(n_711)
);

NAND2xp5_ASAP7_75t_L g712 ( 
.A(n_529),
.B(n_442),
.Y(n_712)
);

NAND2xp5_ASAP7_75t_SL g713 ( 
.A(n_563),
.B(n_269),
.Y(n_713)
);

INVx1_ASAP7_75t_L g714 ( 
.A(n_655),
.Y(n_714)
);

NAND2xp5_ASAP7_75t_L g715 ( 
.A(n_530),
.B(n_442),
.Y(n_715)
);

NOR2xp33_ASAP7_75t_L g716 ( 
.A(n_520),
.B(n_211),
.Y(n_716)
);

NAND2xp5_ASAP7_75t_L g717 ( 
.A(n_530),
.B(n_601),
.Y(n_717)
);

NOR2xp67_ASAP7_75t_L g718 ( 
.A(n_565),
.B(n_485),
.Y(n_718)
);

NAND2xp5_ASAP7_75t_SL g719 ( 
.A(n_563),
.B(n_286),
.Y(n_719)
);

INVx1_ASAP7_75t_L g720 ( 
.A(n_655),
.Y(n_720)
);

NAND2xp5_ASAP7_75t_L g721 ( 
.A(n_603),
.B(n_442),
.Y(n_721)
);

AOI22xp5_ASAP7_75t_L g722 ( 
.A1(n_614),
.A2(n_424),
.B1(n_423),
.B2(n_419),
.Y(n_722)
);

NAND2xp5_ASAP7_75t_L g723 ( 
.A(n_603),
.B(n_470),
.Y(n_723)
);

NAND2xp33_ASAP7_75t_L g724 ( 
.A(n_618),
.B(n_592),
.Y(n_724)
);

NAND2xp33_ASAP7_75t_L g725 ( 
.A(n_585),
.B(n_286),
.Y(n_725)
);

NOR3xp33_ASAP7_75t_SL g726 ( 
.A(n_541),
.B(n_196),
.C(n_194),
.Y(n_726)
);

NAND2xp5_ASAP7_75t_L g727 ( 
.A(n_532),
.B(n_533),
.Y(n_727)
);

OR2x2_ASAP7_75t_L g728 ( 
.A(n_600),
.B(n_194),
.Y(n_728)
);

INVx1_ASAP7_75t_L g729 ( 
.A(n_628),
.Y(n_729)
);

NAND2xp5_ASAP7_75t_L g730 ( 
.A(n_532),
.B(n_470),
.Y(n_730)
);

INVx2_ASAP7_75t_L g731 ( 
.A(n_548),
.Y(n_731)
);

NAND2xp5_ASAP7_75t_L g732 ( 
.A(n_533),
.B(n_470),
.Y(n_732)
);

NAND2xp33_ASAP7_75t_L g733 ( 
.A(n_585),
.B(n_286),
.Y(n_733)
);

INVx1_ASAP7_75t_SL g734 ( 
.A(n_636),
.Y(n_734)
);

INVx2_ASAP7_75t_L g735 ( 
.A(n_551),
.Y(n_735)
);

INVx1_ASAP7_75t_L g736 ( 
.A(n_628),
.Y(n_736)
);

NAND2xp5_ASAP7_75t_SL g737 ( 
.A(n_563),
.B(n_286),
.Y(n_737)
);

NAND2xp5_ASAP7_75t_SL g738 ( 
.A(n_572),
.B(n_286),
.Y(n_738)
);

NOR2xp33_ASAP7_75t_L g739 ( 
.A(n_535),
.B(n_214),
.Y(n_739)
);

NOR2xp33_ASAP7_75t_L g740 ( 
.A(n_599),
.B(n_223),
.Y(n_740)
);

NAND2xp5_ASAP7_75t_L g741 ( 
.A(n_537),
.B(n_470),
.Y(n_741)
);

INVx2_ASAP7_75t_L g742 ( 
.A(n_551),
.Y(n_742)
);

INVx2_ASAP7_75t_L g743 ( 
.A(n_566),
.Y(n_743)
);

INVx1_ASAP7_75t_L g744 ( 
.A(n_593),
.Y(n_744)
);

NOR2xp33_ASAP7_75t_L g745 ( 
.A(n_614),
.B(n_228),
.Y(n_745)
);

INVx1_ASAP7_75t_L g746 ( 
.A(n_593),
.Y(n_746)
);

NOR3xp33_ASAP7_75t_L g747 ( 
.A(n_653),
.B(n_242),
.C(n_239),
.Y(n_747)
);

NOR2x1p5_ASAP7_75t_L g748 ( 
.A(n_619),
.B(n_197),
.Y(n_748)
);

NAND2xp5_ASAP7_75t_SL g749 ( 
.A(n_572),
.B(n_286),
.Y(n_749)
);

NAND2xp5_ASAP7_75t_L g750 ( 
.A(n_537),
.B(n_488),
.Y(n_750)
);

NOR2xp33_ASAP7_75t_L g751 ( 
.A(n_614),
.B(n_245),
.Y(n_751)
);

NAND2xp5_ASAP7_75t_L g752 ( 
.A(n_539),
.B(n_488),
.Y(n_752)
);

NOR2xp33_ASAP7_75t_L g753 ( 
.A(n_614),
.B(n_249),
.Y(n_753)
);

AOI21xp5_ASAP7_75t_L g754 ( 
.A1(n_646),
.A2(n_478),
.B(n_473),
.Y(n_754)
);

INVx1_ASAP7_75t_L g755 ( 
.A(n_539),
.Y(n_755)
);

AND2x4_ASAP7_75t_L g756 ( 
.A(n_549),
.B(n_488),
.Y(n_756)
);

INVx2_ASAP7_75t_L g757 ( 
.A(n_566),
.Y(n_757)
);

OR2x6_ASAP7_75t_L g758 ( 
.A(n_616),
.B(n_486),
.Y(n_758)
);

NAND2xp33_ASAP7_75t_L g759 ( 
.A(n_615),
.B(n_286),
.Y(n_759)
);

AOI22xp33_ASAP7_75t_L g760 ( 
.A1(n_572),
.A2(n_486),
.B1(n_287),
.B2(n_266),
.Y(n_760)
);

INVx1_ASAP7_75t_L g761 ( 
.A(n_543),
.Y(n_761)
);

AND2x4_ASAP7_75t_L g762 ( 
.A(n_549),
.B(n_451),
.Y(n_762)
);

INVx1_ASAP7_75t_L g763 ( 
.A(n_557),
.Y(n_763)
);

INVx1_ASAP7_75t_L g764 ( 
.A(n_557),
.Y(n_764)
);

NAND2xp5_ASAP7_75t_L g765 ( 
.A(n_560),
.B(n_480),
.Y(n_765)
);

NOR2xp33_ASAP7_75t_L g766 ( 
.A(n_661),
.B(n_254),
.Y(n_766)
);

NAND2xp5_ASAP7_75t_L g767 ( 
.A(n_560),
.B(n_480),
.Y(n_767)
);

NAND2xp5_ASAP7_75t_L g768 ( 
.A(n_549),
.B(n_621),
.Y(n_768)
);

NOR2xp33_ASAP7_75t_L g769 ( 
.A(n_666),
.B(n_255),
.Y(n_769)
);

NAND2xp5_ASAP7_75t_L g770 ( 
.A(n_549),
.B(n_480),
.Y(n_770)
);

NAND2xp5_ASAP7_75t_L g771 ( 
.A(n_621),
.B(n_480),
.Y(n_771)
);

NAND2xp5_ASAP7_75t_L g772 ( 
.A(n_621),
.B(n_480),
.Y(n_772)
);

INVx2_ASAP7_75t_L g773 ( 
.A(n_567),
.Y(n_773)
);

INVx1_ASAP7_75t_L g774 ( 
.A(n_564),
.Y(n_774)
);

INVx2_ASAP7_75t_SL g775 ( 
.A(n_616),
.Y(n_775)
);

AND2x4_ASAP7_75t_L g776 ( 
.A(n_562),
.B(n_451),
.Y(n_776)
);

AND2x4_ASAP7_75t_L g777 ( 
.A(n_562),
.B(n_485),
.Y(n_777)
);

AND2x2_ASAP7_75t_L g778 ( 
.A(n_596),
.B(n_660),
.Y(n_778)
);

NAND3x1_ASAP7_75t_L g779 ( 
.A(n_577),
.B(n_259),
.C(n_253),
.Y(n_779)
);

INVx2_ASAP7_75t_L g780 ( 
.A(n_567),
.Y(n_780)
);

NAND2xp5_ASAP7_75t_SL g781 ( 
.A(n_570),
.B(n_329),
.Y(n_781)
);

INVx2_ASAP7_75t_L g782 ( 
.A(n_568),
.Y(n_782)
);

AND2x4_ASAP7_75t_L g783 ( 
.A(n_545),
.B(n_485),
.Y(n_783)
);

NAND2xp5_ASAP7_75t_L g784 ( 
.A(n_526),
.B(n_480),
.Y(n_784)
);

NOR2xp33_ASAP7_75t_L g785 ( 
.A(n_554),
.B(n_256),
.Y(n_785)
);

INVx2_ASAP7_75t_L g786 ( 
.A(n_568),
.Y(n_786)
);

NAND2xp5_ASAP7_75t_SL g787 ( 
.A(n_540),
.B(n_329),
.Y(n_787)
);

NAND2xp5_ASAP7_75t_L g788 ( 
.A(n_526),
.B(n_437),
.Y(n_788)
);

NAND2xp5_ASAP7_75t_SL g789 ( 
.A(n_540),
.B(n_329),
.Y(n_789)
);

NAND2xp5_ASAP7_75t_L g790 ( 
.A(n_526),
.B(n_437),
.Y(n_790)
);

INVx2_ASAP7_75t_L g791 ( 
.A(n_573),
.Y(n_791)
);

NAND2xp5_ASAP7_75t_L g792 ( 
.A(n_526),
.B(n_437),
.Y(n_792)
);

NAND2x1_ASAP7_75t_L g793 ( 
.A(n_518),
.B(n_471),
.Y(n_793)
);

INVx2_ASAP7_75t_L g794 ( 
.A(n_573),
.Y(n_794)
);

NOR2xp33_ASAP7_75t_L g795 ( 
.A(n_609),
.B(n_268),
.Y(n_795)
);

NAND2xp33_ASAP7_75t_L g796 ( 
.A(n_651),
.B(n_329),
.Y(n_796)
);

AOI221xp5_ASAP7_75t_L g797 ( 
.A1(n_638),
.A2(n_344),
.B1(n_346),
.B2(n_347),
.C(n_348),
.Y(n_797)
);

INVx1_ASAP7_75t_L g798 ( 
.A(n_564),
.Y(n_798)
);

NAND2xp5_ASAP7_75t_L g799 ( 
.A(n_580),
.B(n_437),
.Y(n_799)
);

INVx2_ASAP7_75t_SL g800 ( 
.A(n_596),
.Y(n_800)
);

AOI221xp5_ASAP7_75t_L g801 ( 
.A1(n_638),
.A2(n_344),
.B1(n_346),
.B2(n_347),
.C(n_197),
.Y(n_801)
);

NAND2xp5_ASAP7_75t_L g802 ( 
.A(n_580),
.B(n_437),
.Y(n_802)
);

INVx1_ASAP7_75t_L g803 ( 
.A(n_569),
.Y(n_803)
);

INVx1_ASAP7_75t_L g804 ( 
.A(n_569),
.Y(n_804)
);

NOR2xp33_ASAP7_75t_L g805 ( 
.A(n_625),
.B(n_270),
.Y(n_805)
);

INVx2_ASAP7_75t_SL g806 ( 
.A(n_591),
.Y(n_806)
);

INVx2_ASAP7_75t_L g807 ( 
.A(n_575),
.Y(n_807)
);

OAI22xp33_ASAP7_75t_L g808 ( 
.A1(n_619),
.A2(n_198),
.B1(n_201),
.B2(n_203),
.Y(n_808)
);

INVx1_ASAP7_75t_L g809 ( 
.A(n_574),
.Y(n_809)
);

NAND2xp5_ASAP7_75t_SL g810 ( 
.A(n_540),
.B(n_329),
.Y(n_810)
);

AOI22xp33_ASAP7_75t_L g811 ( 
.A1(n_556),
.A2(n_265),
.B1(n_338),
.B2(n_264),
.Y(n_811)
);

BUFx3_ASAP7_75t_L g812 ( 
.A(n_546),
.Y(n_812)
);

NAND2xp5_ASAP7_75t_SL g813 ( 
.A(n_540),
.B(n_329),
.Y(n_813)
);

INVx2_ASAP7_75t_L g814 ( 
.A(n_575),
.Y(n_814)
);

NOR2xp67_ASAP7_75t_L g815 ( 
.A(n_627),
.B(n_489),
.Y(n_815)
);

NAND2x1_ASAP7_75t_L g816 ( 
.A(n_518),
.B(n_471),
.Y(n_816)
);

NOR2xp33_ASAP7_75t_L g817 ( 
.A(n_579),
.B(n_278),
.Y(n_817)
);

NAND2xp5_ASAP7_75t_SL g818 ( 
.A(n_540),
.B(n_471),
.Y(n_818)
);

INVx1_ASAP7_75t_L g819 ( 
.A(n_574),
.Y(n_819)
);

INVx1_ASAP7_75t_L g820 ( 
.A(n_583),
.Y(n_820)
);

INVx2_ASAP7_75t_SL g821 ( 
.A(n_645),
.Y(n_821)
);

NAND2xp5_ASAP7_75t_L g822 ( 
.A(n_580),
.B(n_437),
.Y(n_822)
);

AND2x4_ASAP7_75t_L g823 ( 
.A(n_545),
.B(n_489),
.Y(n_823)
);

NAND2xp5_ASAP7_75t_L g824 ( 
.A(n_580),
.B(n_471),
.Y(n_824)
);

NOR3xp33_ASAP7_75t_L g825 ( 
.A(n_552),
.B(n_298),
.C(n_279),
.Y(n_825)
);

NAND2xp5_ASAP7_75t_L g826 ( 
.A(n_581),
.B(n_473),
.Y(n_826)
);

AOI22xp33_ASAP7_75t_SL g827 ( 
.A1(n_627),
.A2(n_382),
.B1(n_415),
.B2(n_384),
.Y(n_827)
);

NAND2xp5_ASAP7_75t_SL g828 ( 
.A(n_590),
.B(n_261),
.Y(n_828)
);

NOR2xp33_ASAP7_75t_L g829 ( 
.A(n_611),
.B(n_280),
.Y(n_829)
);

NAND2xp5_ASAP7_75t_SL g830 ( 
.A(n_590),
.B(n_327),
.Y(n_830)
);

AND2x2_ASAP7_75t_L g831 ( 
.A(n_544),
.B(n_371),
.Y(n_831)
);

AOI22xp33_ASAP7_75t_L g832 ( 
.A1(n_657),
.A2(n_340),
.B1(n_475),
.B2(n_501),
.Y(n_832)
);

INVx2_ASAP7_75t_SL g833 ( 
.A(n_649),
.Y(n_833)
);

NOR2xp67_ASAP7_75t_L g834 ( 
.A(n_617),
.B(n_489),
.Y(n_834)
);

AO22x2_ASAP7_75t_L g835 ( 
.A1(n_516),
.A2(n_501),
.B1(n_499),
.B2(n_498),
.Y(n_835)
);

AOI22xp33_ASAP7_75t_L g836 ( 
.A1(n_665),
.A2(n_475),
.B1(n_498),
.B2(n_501),
.Y(n_836)
);

AOI21xp5_ASAP7_75t_L g837 ( 
.A1(n_687),
.A2(n_663),
.B(n_656),
.Y(n_837)
);

A2O1A1Ixp33_ASAP7_75t_L g838 ( 
.A1(n_681),
.A2(n_642),
.B(n_664),
.C(n_597),
.Y(n_838)
);

INVx1_ASAP7_75t_L g839 ( 
.A(n_674),
.Y(n_839)
);

NAND2xp5_ASAP7_75t_L g840 ( 
.A(n_677),
.B(n_581),
.Y(n_840)
);

AND2x2_ASAP7_75t_L g841 ( 
.A(n_778),
.B(n_604),
.Y(n_841)
);

HB1xp67_ASAP7_75t_L g842 ( 
.A(n_758),
.Y(n_842)
);

INVx3_ASAP7_75t_L g843 ( 
.A(n_783),
.Y(n_843)
);

NAND2xp5_ASAP7_75t_L g844 ( 
.A(n_686),
.B(n_581),
.Y(n_844)
);

AOI21xp5_ASAP7_75t_L g845 ( 
.A1(n_687),
.A2(n_684),
.B(n_698),
.Y(n_845)
);

AOI21xp5_ASAP7_75t_L g846 ( 
.A1(n_684),
.A2(n_531),
.B(n_518),
.Y(n_846)
);

NAND2xp5_ASAP7_75t_L g847 ( 
.A(n_686),
.B(n_581),
.Y(n_847)
);

NAND2xp5_ASAP7_75t_L g848 ( 
.A(n_706),
.B(n_597),
.Y(n_848)
);

NAND2xp5_ASAP7_75t_SL g849 ( 
.A(n_680),
.B(n_590),
.Y(n_849)
);

NOR2xp33_ASAP7_75t_L g850 ( 
.A(n_740),
.B(n_635),
.Y(n_850)
);

HB1xp67_ASAP7_75t_L g851 ( 
.A(n_758),
.Y(n_851)
);

O2A1O1Ixp5_ASAP7_75t_L g852 ( 
.A1(n_781),
.A2(n_597),
.B(n_644),
.C(n_518),
.Y(n_852)
);

NOR2xp33_ASAP7_75t_L g853 ( 
.A(n_740),
.B(n_376),
.Y(n_853)
);

AOI21xp5_ASAP7_75t_L g854 ( 
.A1(n_698),
.A2(n_538),
.B(n_531),
.Y(n_854)
);

AOI21xp5_ASAP7_75t_L g855 ( 
.A1(n_690),
.A2(n_538),
.B(n_531),
.Y(n_855)
);

BUFx2_ASAP7_75t_L g856 ( 
.A(n_734),
.Y(n_856)
);

INVx1_ASAP7_75t_L g857 ( 
.A(n_774),
.Y(n_857)
);

AND2x2_ASAP7_75t_L g858 ( 
.A(n_675),
.B(n_383),
.Y(n_858)
);

BUFx6f_ASAP7_75t_L g859 ( 
.A(n_680),
.Y(n_859)
);

NAND2xp5_ASAP7_75t_SL g860 ( 
.A(n_680),
.B(n_590),
.Y(n_860)
);

NAND2xp5_ASAP7_75t_SL g861 ( 
.A(n_680),
.B(n_590),
.Y(n_861)
);

INVx1_ASAP7_75t_L g862 ( 
.A(n_798),
.Y(n_862)
);

AOI21xp5_ASAP7_75t_L g863 ( 
.A1(n_692),
.A2(n_538),
.B(n_531),
.Y(n_863)
);

BUFx2_ASAP7_75t_L g864 ( 
.A(n_775),
.Y(n_864)
);

INVx2_ASAP7_75t_L g865 ( 
.A(n_673),
.Y(n_865)
);

AND2x2_ASAP7_75t_L g866 ( 
.A(n_675),
.B(n_418),
.Y(n_866)
);

CKINVDCx8_ASAP7_75t_R g867 ( 
.A(n_683),
.Y(n_867)
);

NAND2xp5_ASAP7_75t_L g868 ( 
.A(n_670),
.B(n_597),
.Y(n_868)
);

NOR2xp33_ASAP7_75t_L g869 ( 
.A(n_708),
.B(n_521),
.Y(n_869)
);

INVx1_ASAP7_75t_SL g870 ( 
.A(n_800),
.Y(n_870)
);

BUFx6f_ASAP7_75t_L g871 ( 
.A(n_812),
.Y(n_871)
);

AOI22xp5_ASAP7_75t_L g872 ( 
.A1(n_708),
.A2(n_525),
.B1(n_550),
.B2(n_654),
.Y(n_872)
);

NOR2xp33_ASAP7_75t_L g873 ( 
.A(n_668),
.B(n_561),
.Y(n_873)
);

AOI21xp5_ASAP7_75t_L g874 ( 
.A1(n_707),
.A2(n_558),
.B(n_538),
.Y(n_874)
);

CKINVDCx10_ASAP7_75t_R g875 ( 
.A(n_671),
.Y(n_875)
);

A2O1A1Ixp33_ASAP7_75t_L g876 ( 
.A1(n_817),
.A2(n_667),
.B(n_583),
.C(n_589),
.Y(n_876)
);

NOR2xp33_ASAP7_75t_L g877 ( 
.A(n_678),
.B(n_516),
.Y(n_877)
);

INVx3_ASAP7_75t_L g878 ( 
.A(n_783),
.Y(n_878)
);

NOR2xp33_ASAP7_75t_L g879 ( 
.A(n_695),
.B(n_525),
.Y(n_879)
);

NOR2xp67_ASAP7_75t_L g880 ( 
.A(n_795),
.B(n_301),
.Y(n_880)
);

AOI21xp5_ASAP7_75t_L g881 ( 
.A1(n_710),
.A2(n_644),
.B(n_558),
.Y(n_881)
);

NAND2xp5_ASAP7_75t_SL g882 ( 
.A(n_768),
.B(n_610),
.Y(n_882)
);

NAND2xp5_ASAP7_75t_L g883 ( 
.A(n_672),
.B(n_587),
.Y(n_883)
);

INVx2_ASAP7_75t_L g884 ( 
.A(n_709),
.Y(n_884)
);

AOI22xp5_ASAP7_75t_L g885 ( 
.A1(n_756),
.A2(n_654),
.B1(n_525),
.B2(n_550),
.Y(n_885)
);

AOI21xp5_ASAP7_75t_L g886 ( 
.A1(n_712),
.A2(n_644),
.B(n_558),
.Y(n_886)
);

INVx1_ASAP7_75t_L g887 ( 
.A(n_803),
.Y(n_887)
);

AND2x2_ASAP7_75t_L g888 ( 
.A(n_758),
.B(n_201),
.Y(n_888)
);

OAI21xp5_ASAP7_75t_L g889 ( 
.A1(n_702),
.A2(n_589),
.B(n_587),
.Y(n_889)
);

INVx1_ASAP7_75t_SL g890 ( 
.A(n_685),
.Y(n_890)
);

NAND2xp5_ASAP7_75t_L g891 ( 
.A(n_718),
.B(n_594),
.Y(n_891)
);

AND2x2_ASAP7_75t_L g892 ( 
.A(n_685),
.B(n_203),
.Y(n_892)
);

AOI21xp5_ASAP7_75t_L g893 ( 
.A1(n_715),
.A2(n_644),
.B(n_558),
.Y(n_893)
);

NAND2xp5_ASAP7_75t_L g894 ( 
.A(n_760),
.B(n_594),
.Y(n_894)
);

NAND2xp5_ASAP7_75t_SL g895 ( 
.A(n_717),
.B(n_610),
.Y(n_895)
);

BUFx3_ASAP7_75t_L g896 ( 
.A(n_685),
.Y(n_896)
);

NAND2xp5_ASAP7_75t_L g897 ( 
.A(n_760),
.B(n_602),
.Y(n_897)
);

INVx1_ASAP7_75t_SL g898 ( 
.A(n_728),
.Y(n_898)
);

A2O1A1Ixp33_ASAP7_75t_L g899 ( 
.A1(n_724),
.A2(n_496),
.B(n_505),
.C(n_620),
.Y(n_899)
);

AND2x2_ASAP7_75t_L g900 ( 
.A(n_682),
.B(n_205),
.Y(n_900)
);

INVx2_ASAP7_75t_L g901 ( 
.A(n_731),
.Y(n_901)
);

AND2x2_ASAP7_75t_L g902 ( 
.A(n_688),
.B(n_490),
.Y(n_902)
);

NAND2xp5_ASAP7_75t_L g903 ( 
.A(n_815),
.B(n_602),
.Y(n_903)
);

OAI22xp5_ASAP7_75t_L g904 ( 
.A1(n_691),
.A2(n_654),
.B1(n_550),
.B2(n_606),
.Y(n_904)
);

AND2x2_ASAP7_75t_L g905 ( 
.A(n_701),
.B(n_490),
.Y(n_905)
);

NOR2xp33_ASAP7_75t_L g906 ( 
.A(n_676),
.B(n_606),
.Y(n_906)
);

INVx2_ASAP7_75t_SL g907 ( 
.A(n_777),
.Y(n_907)
);

OAI21xp5_ASAP7_75t_L g908 ( 
.A1(n_702),
.A2(n_667),
.B(n_613),
.Y(n_908)
);

HB1xp67_ASAP7_75t_L g909 ( 
.A(n_756),
.Y(n_909)
);

BUFx6f_ASAP7_75t_L g910 ( 
.A(n_812),
.Y(n_910)
);

NAND2xp5_ASAP7_75t_L g911 ( 
.A(n_703),
.B(n_613),
.Y(n_911)
);

OAI21xp5_ASAP7_75t_L g912 ( 
.A1(n_704),
.A2(n_719),
.B(n_713),
.Y(n_912)
);

A2O1A1Ixp33_ASAP7_75t_L g913 ( 
.A1(n_744),
.A2(n_505),
.B(n_496),
.C(n_658),
.Y(n_913)
);

NAND2xp5_ASAP7_75t_L g914 ( 
.A(n_714),
.B(n_620),
.Y(n_914)
);

NAND2xp5_ASAP7_75t_L g915 ( 
.A(n_720),
.B(n_626),
.Y(n_915)
);

NAND2x1p5_ASAP7_75t_L g916 ( 
.A(n_823),
.B(n_595),
.Y(n_916)
);

AOI21xp5_ASAP7_75t_L g917 ( 
.A1(n_730),
.A2(n_546),
.B(n_610),
.Y(n_917)
);

AOI21xp5_ASAP7_75t_L g918 ( 
.A1(n_732),
.A2(n_546),
.B(n_610),
.Y(n_918)
);

AOI21xp5_ASAP7_75t_L g919 ( 
.A1(n_741),
.A2(n_693),
.B(n_771),
.Y(n_919)
);

INVx3_ASAP7_75t_L g920 ( 
.A(n_823),
.Y(n_920)
);

O2A1O1Ixp33_ASAP7_75t_L g921 ( 
.A1(n_781),
.A2(n_626),
.B(n_640),
.C(n_658),
.Y(n_921)
);

NAND2xp5_ASAP7_75t_SL g922 ( 
.A(n_746),
.B(n_610),
.Y(n_922)
);

INVx1_ASAP7_75t_L g923 ( 
.A(n_804),
.Y(n_923)
);

NAND2xp5_ASAP7_75t_L g924 ( 
.A(n_727),
.B(n_640),
.Y(n_924)
);

AOI21xp5_ASAP7_75t_L g925 ( 
.A1(n_772),
.A2(n_546),
.B(n_639),
.Y(n_925)
);

INVx4_ASAP7_75t_L g926 ( 
.A(n_762),
.Y(n_926)
);

NOR2xp33_ASAP7_75t_L g927 ( 
.A(n_676),
.B(n_643),
.Y(n_927)
);

NAND2xp5_ASAP7_75t_L g928 ( 
.A(n_721),
.B(n_643),
.Y(n_928)
);

AOI21x1_ASAP7_75t_L g929 ( 
.A1(n_704),
.A2(n_650),
.B(n_659),
.Y(n_929)
);

NAND2xp5_ASAP7_75t_L g930 ( 
.A(n_723),
.B(n_650),
.Y(n_930)
);

BUFx12f_ASAP7_75t_L g931 ( 
.A(n_669),
.Y(n_931)
);

INVx2_ASAP7_75t_SL g932 ( 
.A(n_777),
.Y(n_932)
);

A2O1A1Ixp33_ASAP7_75t_L g933 ( 
.A1(n_817),
.A2(n_505),
.B(n_496),
.C(n_498),
.Y(n_933)
);

INVx2_ASAP7_75t_L g934 ( 
.A(n_735),
.Y(n_934)
);

CKINVDCx16_ASAP7_75t_R g935 ( 
.A(n_722),
.Y(n_935)
);

INVxp33_ASAP7_75t_SL g936 ( 
.A(n_700),
.Y(n_936)
);

O2A1O1Ixp33_ASAP7_75t_L g937 ( 
.A1(n_679),
.A2(n_662),
.B(n_659),
.C(n_652),
.Y(n_937)
);

AO21x1_ASAP7_75t_L g938 ( 
.A1(n_691),
.A2(n_662),
.B(n_652),
.Y(n_938)
);

AOI21xp5_ASAP7_75t_L g939 ( 
.A1(n_765),
.A2(n_546),
.B(n_647),
.Y(n_939)
);

INVx2_ASAP7_75t_L g940 ( 
.A(n_742),
.Y(n_940)
);

NAND2xp5_ASAP7_75t_L g941 ( 
.A(n_755),
.B(n_598),
.Y(n_941)
);

A2O1A1Ixp33_ASAP7_75t_L g942 ( 
.A1(n_829),
.A2(n_648),
.B(n_634),
.C(n_633),
.Y(n_942)
);

INVx2_ASAP7_75t_L g943 ( 
.A(n_743),
.Y(n_943)
);

OAI21xp5_ASAP7_75t_L g944 ( 
.A1(n_713),
.A2(n_648),
.B(n_634),
.Y(n_944)
);

AOI21xp5_ASAP7_75t_L g945 ( 
.A1(n_767),
.A2(n_647),
.B(n_639),
.Y(n_945)
);

NAND2xp5_ASAP7_75t_L g946 ( 
.A(n_761),
.B(n_598),
.Y(n_946)
);

AOI21xp5_ASAP7_75t_L g947 ( 
.A1(n_770),
.A2(n_647),
.B(n_639),
.Y(n_947)
);

AOI21xp5_ASAP7_75t_L g948 ( 
.A1(n_696),
.A2(n_647),
.B(n_639),
.Y(n_948)
);

AOI21x1_ASAP7_75t_L g949 ( 
.A1(n_719),
.A2(n_605),
.B(n_607),
.Y(n_949)
);

NAND2xp5_ASAP7_75t_L g950 ( 
.A(n_763),
.B(n_605),
.Y(n_950)
);

AOI21xp5_ASAP7_75t_L g951 ( 
.A1(n_696),
.A2(n_647),
.B(n_639),
.Y(n_951)
);

NAND2xp5_ASAP7_75t_L g952 ( 
.A(n_764),
.B(n_607),
.Y(n_952)
);

AOI21xp5_ASAP7_75t_L g953 ( 
.A1(n_750),
.A2(n_595),
.B(n_612),
.Y(n_953)
);

AND2x2_ASAP7_75t_L g954 ( 
.A(n_716),
.B(n_490),
.Y(n_954)
);

O2A1O1Ixp33_ASAP7_75t_SL g955 ( 
.A1(n_737),
.A2(n_633),
.B(n_631),
.C(n_630),
.Y(n_955)
);

INVxp67_ASAP7_75t_SL g956 ( 
.A(n_752),
.Y(n_956)
);

INVx2_ASAP7_75t_L g957 ( 
.A(n_757),
.Y(n_957)
);

A2O1A1Ixp33_ASAP7_75t_L g958 ( 
.A1(n_829),
.A2(n_751),
.B(n_753),
.C(n_745),
.Y(n_958)
);

OAI21xp33_ASAP7_75t_L g959 ( 
.A1(n_716),
.A2(n_305),
.B(n_289),
.Y(n_959)
);

NAND2xp5_ASAP7_75t_L g960 ( 
.A(n_795),
.B(n_608),
.Y(n_960)
);

INVx3_ASAP7_75t_L g961 ( 
.A(n_699),
.Y(n_961)
);

OAI21xp5_ASAP7_75t_L g962 ( 
.A1(n_737),
.A2(n_631),
.B(n_630),
.Y(n_962)
);

AOI21xp5_ASAP7_75t_L g963 ( 
.A1(n_694),
.A2(n_612),
.B(n_595),
.Y(n_963)
);

OAI21xp5_ASAP7_75t_L g964 ( 
.A1(n_738),
.A2(n_629),
.B(n_608),
.Y(n_964)
);

AOI21xp5_ASAP7_75t_L g965 ( 
.A1(n_725),
.A2(n_612),
.B(n_595),
.Y(n_965)
);

NAND2xp5_ASAP7_75t_L g966 ( 
.A(n_805),
.B(n_629),
.Y(n_966)
);

AOI22xp5_ASAP7_75t_SL g967 ( 
.A1(n_785),
.A2(n_343),
.B1(n_336),
.B2(n_334),
.Y(n_967)
);

AOI21xp5_ASAP7_75t_L g968 ( 
.A1(n_733),
.A2(n_612),
.B(n_595),
.Y(n_968)
);

NOR2x1_ASAP7_75t_L g969 ( 
.A(n_748),
.B(n_443),
.Y(n_969)
);

O2A1O1Ixp33_ASAP7_75t_L g970 ( 
.A1(n_697),
.A2(n_749),
.B(n_738),
.C(n_808),
.Y(n_970)
);

AOI21xp5_ASAP7_75t_L g971 ( 
.A1(n_749),
.A2(n_612),
.B(n_588),
.Y(n_971)
);

INVx4_ASAP7_75t_L g972 ( 
.A(n_762),
.Y(n_972)
);

AOI21xp5_ASAP7_75t_L g973 ( 
.A1(n_711),
.A2(n_588),
.B(n_586),
.Y(n_973)
);

AOI21xp5_ASAP7_75t_L g974 ( 
.A1(n_793),
.A2(n_586),
.B(n_582),
.Y(n_974)
);

NAND2xp5_ASAP7_75t_L g975 ( 
.A(n_805),
.B(n_576),
.Y(n_975)
);

AND2x4_ASAP7_75t_L g976 ( 
.A(n_776),
.B(n_545),
.Y(n_976)
);

NOR2xp33_ASAP7_75t_L g977 ( 
.A(n_739),
.B(n_304),
.Y(n_977)
);

CKINVDCx20_ASAP7_75t_R g978 ( 
.A(n_831),
.Y(n_978)
);

NOR2xp67_ASAP7_75t_L g979 ( 
.A(n_766),
.B(n_309),
.Y(n_979)
);

AND2x4_ASAP7_75t_L g980 ( 
.A(n_776),
.B(n_545),
.Y(n_980)
);

AOI21xp5_ASAP7_75t_L g981 ( 
.A1(n_816),
.A2(n_824),
.B(n_788),
.Y(n_981)
);

NAND2xp5_ASAP7_75t_L g982 ( 
.A(n_729),
.B(n_576),
.Y(n_982)
);

A2O1A1Ixp33_ASAP7_75t_L g983 ( 
.A1(n_739),
.A2(n_582),
.B(n_496),
.C(n_505),
.Y(n_983)
);

INVx1_ASAP7_75t_L g984 ( 
.A(n_809),
.Y(n_984)
);

INVx1_ASAP7_75t_L g985 ( 
.A(n_819),
.Y(n_985)
);

AO22x1_ASAP7_75t_L g986 ( 
.A1(n_766),
.A2(n_306),
.B1(n_332),
.B2(n_326),
.Y(n_986)
);

AOI21xp33_ASAP7_75t_L g987 ( 
.A1(n_785),
.A2(n_342),
.B(n_324),
.Y(n_987)
);

NAND2xp5_ASAP7_75t_L g988 ( 
.A(n_736),
.B(n_496),
.Y(n_988)
);

INVxp67_ASAP7_75t_L g989 ( 
.A(n_745),
.Y(n_989)
);

AOI21xp5_ASAP7_75t_L g990 ( 
.A1(n_784),
.A2(n_478),
.B(n_459),
.Y(n_990)
);

AO21x1_ASAP7_75t_L g991 ( 
.A1(n_705),
.A2(n_472),
.B(n_444),
.Y(n_991)
);

AOI21x1_ASAP7_75t_L g992 ( 
.A1(n_818),
.A2(n_463),
.B(n_443),
.Y(n_992)
);

NAND2xp5_ASAP7_75t_SL g993 ( 
.A(n_834),
.B(n_705),
.Y(n_993)
);

AOI21xp5_ASAP7_75t_L g994 ( 
.A1(n_790),
.A2(n_799),
.B(n_792),
.Y(n_994)
);

INVx3_ASAP7_75t_L g995 ( 
.A(n_820),
.Y(n_995)
);

INVx4_ASAP7_75t_L g996 ( 
.A(n_671),
.Y(n_996)
);

NAND2xp5_ASAP7_75t_SL g997 ( 
.A(n_832),
.B(n_314),
.Y(n_997)
);

NAND2xp5_ASAP7_75t_L g998 ( 
.A(n_751),
.B(n_505),
.Y(n_998)
);

OAI21xp5_ASAP7_75t_L g999 ( 
.A1(n_689),
.A2(n_475),
.B(n_448),
.Y(n_999)
);

NAND2xp5_ASAP7_75t_L g1000 ( 
.A(n_753),
.B(n_505),
.Y(n_1000)
);

AOI21xp5_ASAP7_75t_L g1001 ( 
.A1(n_802),
.A2(n_459),
.B(n_443),
.Y(n_1001)
);

NAND2xp5_ASAP7_75t_L g1002 ( 
.A(n_769),
.B(n_444),
.Y(n_1002)
);

BUFx2_ASAP7_75t_L g1003 ( 
.A(n_835),
.Y(n_1003)
);

NOR2xp33_ASAP7_75t_L g1004 ( 
.A(n_808),
.B(n_316),
.Y(n_1004)
);

NAND2xp5_ASAP7_75t_L g1005 ( 
.A(n_769),
.B(n_444),
.Y(n_1005)
);

AOI21xp5_ASAP7_75t_L g1006 ( 
.A1(n_822),
.A2(n_463),
.B(n_448),
.Y(n_1006)
);

NAND2xp5_ASAP7_75t_L g1007 ( 
.A(n_836),
.B(n_448),
.Y(n_1007)
);

INVx1_ASAP7_75t_L g1008 ( 
.A(n_773),
.Y(n_1008)
);

INVx2_ASAP7_75t_L g1009 ( 
.A(n_780),
.Y(n_1009)
);

NAND2xp5_ASAP7_75t_L g1010 ( 
.A(n_836),
.B(n_449),
.Y(n_1010)
);

A2O1A1Ixp33_ASAP7_75t_L g1011 ( 
.A1(n_754),
.A2(n_494),
.B(n_497),
.C(n_499),
.Y(n_1011)
);

BUFx4f_ASAP7_75t_L g1012 ( 
.A(n_806),
.Y(n_1012)
);

INVx1_ASAP7_75t_L g1013 ( 
.A(n_782),
.Y(n_1013)
);

NAND2xp5_ASAP7_75t_L g1014 ( 
.A(n_786),
.B(n_449),
.Y(n_1014)
);

A2O1A1Ixp33_ASAP7_75t_L g1015 ( 
.A1(n_797),
.A2(n_494),
.B(n_497),
.C(n_499),
.Y(n_1015)
);

NAND2xp5_ASAP7_75t_L g1016 ( 
.A(n_791),
.B(n_449),
.Y(n_1016)
);

NAND2xp5_ASAP7_75t_L g1017 ( 
.A(n_794),
.B(n_454),
.Y(n_1017)
);

NAND2xp5_ASAP7_75t_L g1018 ( 
.A(n_807),
.B(n_454),
.Y(n_1018)
);

OR2x6_ASAP7_75t_L g1019 ( 
.A(n_821),
.B(n_494),
.Y(n_1019)
);

A2O1A1Ixp33_ASAP7_75t_L g1020 ( 
.A1(n_801),
.A2(n_497),
.B(n_317),
.C(n_513),
.Y(n_1020)
);

AOI21xp5_ASAP7_75t_L g1021 ( 
.A1(n_759),
.A2(n_463),
.B(n_454),
.Y(n_1021)
);

NAND2xp5_ASAP7_75t_L g1022 ( 
.A(n_814),
.B(n_826),
.Y(n_1022)
);

NOR2xp33_ASAP7_75t_L g1023 ( 
.A(n_825),
.B(n_315),
.Y(n_1023)
);

NAND2xp5_ASAP7_75t_L g1024 ( 
.A(n_811),
.B(n_459),
.Y(n_1024)
);

NAND2xp5_ASAP7_75t_SL g1025 ( 
.A(n_832),
.B(n_318),
.Y(n_1025)
);

AOI22xp5_ASAP7_75t_L g1026 ( 
.A1(n_747),
.A2(n_321),
.B1(n_322),
.B2(n_323),
.Y(n_1026)
);

INVx1_ASAP7_75t_L g1027 ( 
.A(n_818),
.Y(n_1027)
);

OR2x6_ASAP7_75t_L g1028 ( 
.A(n_856),
.B(n_835),
.Y(n_1028)
);

AOI21x1_ASAP7_75t_L g1029 ( 
.A1(n_922),
.A2(n_787),
.B(n_789),
.Y(n_1029)
);

NAND2xp5_ASAP7_75t_L g1030 ( 
.A(n_977),
.B(n_835),
.Y(n_1030)
);

A2O1A1Ixp33_ASAP7_75t_L g1031 ( 
.A1(n_977),
.A2(n_726),
.B(n_811),
.C(n_796),
.Y(n_1031)
);

BUFx6f_ASAP7_75t_L g1032 ( 
.A(n_859),
.Y(n_1032)
);

AND2x2_ASAP7_75t_L g1033 ( 
.A(n_841),
.B(n_898),
.Y(n_1033)
);

A2O1A1Ixp33_ASAP7_75t_L g1034 ( 
.A1(n_958),
.A2(n_813),
.B(n_789),
.C(n_810),
.Y(n_1034)
);

OAI21x1_ASAP7_75t_SL g1035 ( 
.A1(n_845),
.A2(n_833),
.B(n_468),
.Y(n_1035)
);

INVx3_ASAP7_75t_L g1036 ( 
.A(n_859),
.Y(n_1036)
);

AOI21xp5_ASAP7_75t_L g1037 ( 
.A1(n_846),
.A2(n_830),
.B(n_828),
.Y(n_1037)
);

INVx3_ASAP7_75t_L g1038 ( 
.A(n_859),
.Y(n_1038)
);

CKINVDCx5p33_ASAP7_75t_R g1039 ( 
.A(n_936),
.Y(n_1039)
);

AOI22xp5_ASAP7_75t_L g1040 ( 
.A1(n_989),
.A2(n_827),
.B1(n_779),
.B2(n_830),
.Y(n_1040)
);

NAND2xp5_ASAP7_75t_SL g1041 ( 
.A(n_989),
.B(n_337),
.Y(n_1041)
);

BUFx2_ASAP7_75t_L g1042 ( 
.A(n_858),
.Y(n_1042)
);

A2O1A1Ixp33_ASAP7_75t_L g1043 ( 
.A1(n_958),
.A2(n_813),
.B(n_810),
.C(n_787),
.Y(n_1043)
);

NAND2xp5_ASAP7_75t_SL g1044 ( 
.A(n_909),
.B(n_926),
.Y(n_1044)
);

O2A1O1Ixp33_ASAP7_75t_L g1045 ( 
.A1(n_1020),
.A2(n_828),
.B(n_472),
.C(n_468),
.Y(n_1045)
);

OAI22xp5_ASAP7_75t_L g1046 ( 
.A1(n_894),
.A2(n_513),
.B1(n_502),
.B2(n_493),
.Y(n_1046)
);

OAI22xp5_ASAP7_75t_L g1047 ( 
.A1(n_897),
.A2(n_513),
.B1(n_502),
.B2(n_493),
.Y(n_1047)
);

INVx1_ASAP7_75t_L g1048 ( 
.A(n_857),
.Y(n_1048)
);

NAND2xp5_ASAP7_75t_L g1049 ( 
.A(n_956),
.B(n_954),
.Y(n_1049)
);

A2O1A1Ixp33_ASAP7_75t_L g1050 ( 
.A1(n_970),
.A2(n_513),
.B(n_502),
.C(n_493),
.Y(n_1050)
);

INVx1_ASAP7_75t_L g1051 ( 
.A(n_862),
.Y(n_1051)
);

BUFx8_ASAP7_75t_SL g1052 ( 
.A(n_931),
.Y(n_1052)
);

AOI21xp5_ASAP7_75t_L g1053 ( 
.A1(n_840),
.A2(n_502),
.B(n_493),
.Y(n_1053)
);

NAND2x1p5_ASAP7_75t_L g1054 ( 
.A(n_859),
.B(n_472),
.Y(n_1054)
);

INVx1_ASAP7_75t_L g1055 ( 
.A(n_887),
.Y(n_1055)
);

AOI21xp5_ASAP7_75t_L g1056 ( 
.A1(n_919),
.A2(n_484),
.B(n_468),
.Y(n_1056)
);

AOI21xp5_ASAP7_75t_L g1057 ( 
.A1(n_917),
.A2(n_918),
.B(n_837),
.Y(n_1057)
);

NAND2xp5_ASAP7_75t_L g1058 ( 
.A(n_956),
.B(n_839),
.Y(n_1058)
);

AOI21xp5_ASAP7_75t_L g1059 ( 
.A1(n_912),
.A2(n_484),
.B(n_483),
.Y(n_1059)
);

INVx1_ASAP7_75t_L g1060 ( 
.A(n_923),
.Y(n_1060)
);

AND2x2_ASAP7_75t_L g1061 ( 
.A(n_850),
.B(n_853),
.Y(n_1061)
);

NAND2xp5_ASAP7_75t_L g1062 ( 
.A(n_928),
.B(n_484),
.Y(n_1062)
);

NAND2xp5_ASAP7_75t_L g1063 ( 
.A(n_930),
.B(n_484),
.Y(n_1063)
);

OAI21xp5_ASAP7_75t_L g1064 ( 
.A1(n_899),
.A2(n_475),
.B(n_483),
.Y(n_1064)
);

OAI22xp5_ASAP7_75t_L g1065 ( 
.A1(n_1020),
.A2(n_481),
.B1(n_483),
.B2(n_12),
.Y(n_1065)
);

NAND2xp5_ASAP7_75t_L g1066 ( 
.A(n_848),
.B(n_483),
.Y(n_1066)
);

O2A1O1Ixp33_ASAP7_75t_SL g1067 ( 
.A1(n_838),
.A2(n_71),
.B(n_64),
.C(n_174),
.Y(n_1067)
);

NAND2xp5_ASAP7_75t_L g1068 ( 
.A(n_906),
.B(n_927),
.Y(n_1068)
);

BUFx2_ASAP7_75t_L g1069 ( 
.A(n_866),
.Y(n_1069)
);

A2O1A1Ixp33_ASAP7_75t_L g1070 ( 
.A1(n_1023),
.A2(n_483),
.B(n_481),
.C(n_475),
.Y(n_1070)
);

AND2x4_ASAP7_75t_L g1071 ( 
.A(n_976),
.B(n_980),
.Y(n_1071)
);

AND2x4_ASAP7_75t_L g1072 ( 
.A(n_976),
.B(n_116),
.Y(n_1072)
);

O2A1O1Ixp33_ASAP7_75t_L g1073 ( 
.A1(n_987),
.A2(n_1004),
.B(n_1015),
.C(n_959),
.Y(n_1073)
);

AOI21xp5_ASAP7_75t_L g1074 ( 
.A1(n_925),
.A2(n_483),
.B(n_481),
.Y(n_1074)
);

NAND2xp5_ASAP7_75t_L g1075 ( 
.A(n_902),
.B(n_483),
.Y(n_1075)
);

INVx2_ASAP7_75t_SL g1076 ( 
.A(n_864),
.Y(n_1076)
);

OAI22xp5_ASAP7_75t_L g1077 ( 
.A1(n_906),
.A2(n_483),
.B1(n_481),
.B2(n_15),
.Y(n_1077)
);

OAI21xp5_ASAP7_75t_L g1078 ( 
.A1(n_899),
.A2(n_475),
.B(n_483),
.Y(n_1078)
);

INVx3_ASAP7_75t_L g1079 ( 
.A(n_871),
.Y(n_1079)
);

AOI21xp5_ASAP7_75t_L g1080 ( 
.A1(n_960),
.A2(n_481),
.B(n_475),
.Y(n_1080)
);

NAND2xp5_ASAP7_75t_L g1081 ( 
.A(n_905),
.B(n_481),
.Y(n_1081)
);

AO21x1_ASAP7_75t_L g1082 ( 
.A1(n_998),
.A2(n_8),
.B(n_11),
.Y(n_1082)
);

A2O1A1Ixp33_ASAP7_75t_L g1083 ( 
.A1(n_1023),
.A2(n_481),
.B(n_475),
.C(n_19),
.Y(n_1083)
);

OAI21xp33_ASAP7_75t_SL g1084 ( 
.A1(n_922),
.A2(n_8),
.B(n_18),
.Y(n_1084)
);

OR2x2_ASAP7_75t_L g1085 ( 
.A(n_853),
.B(n_481),
.Y(n_1085)
);

INVx2_ASAP7_75t_L g1086 ( 
.A(n_995),
.Y(n_1086)
);

INVx2_ASAP7_75t_L g1087 ( 
.A(n_995),
.Y(n_1087)
);

NAND2xp5_ASAP7_75t_SL g1088 ( 
.A(n_909),
.B(n_481),
.Y(n_1088)
);

INVx8_ASAP7_75t_L g1089 ( 
.A(n_980),
.Y(n_1089)
);

INVx1_ASAP7_75t_L g1090 ( 
.A(n_984),
.Y(n_1090)
);

BUFx5_ASAP7_75t_L g1091 ( 
.A(n_1027),
.Y(n_1091)
);

O2A1O1Ixp33_ASAP7_75t_SL g1092 ( 
.A1(n_933),
.A2(n_78),
.B(n_170),
.C(n_165),
.Y(n_1092)
);

AOI21xp5_ASAP7_75t_L g1093 ( 
.A1(n_966),
.A2(n_172),
.B(n_161),
.Y(n_1093)
);

AND2x2_ASAP7_75t_L g1094 ( 
.A(n_850),
.B(n_21),
.Y(n_1094)
);

AOI22xp33_ASAP7_75t_L g1095 ( 
.A1(n_1004),
.A2(n_22),
.B1(n_23),
.B2(n_25),
.Y(n_1095)
);

INVx1_ASAP7_75t_SL g1096 ( 
.A(n_870),
.Y(n_1096)
);

INVx4_ASAP7_75t_L g1097 ( 
.A(n_871),
.Y(n_1097)
);

NOR2xp33_ASAP7_75t_R g1098 ( 
.A(n_978),
.B(n_160),
.Y(n_1098)
);

NAND2xp5_ASAP7_75t_L g1099 ( 
.A(n_927),
.B(n_154),
.Y(n_1099)
);

NAND2xp5_ASAP7_75t_SL g1100 ( 
.A(n_926),
.B(n_149),
.Y(n_1100)
);

NAND2xp5_ASAP7_75t_SL g1101 ( 
.A(n_972),
.B(n_139),
.Y(n_1101)
);

AND2x2_ASAP7_75t_L g1102 ( 
.A(n_900),
.B(n_22),
.Y(n_1102)
);

OAI22xp5_ASAP7_75t_L g1103 ( 
.A1(n_1007),
.A2(n_23),
.B1(n_27),
.B2(n_28),
.Y(n_1103)
);

NAND3xp33_ASAP7_75t_SL g1104 ( 
.A(n_869),
.B(n_27),
.C(n_30),
.Y(n_1104)
);

INVx4_ASAP7_75t_L g1105 ( 
.A(n_871),
.Y(n_1105)
);

INVx2_ASAP7_75t_L g1106 ( 
.A(n_865),
.Y(n_1106)
);

O2A1O1Ixp33_ASAP7_75t_L g1107 ( 
.A1(n_1015),
.A2(n_30),
.B(n_32),
.C(n_33),
.Y(n_1107)
);

AND2x4_ASAP7_75t_L g1108 ( 
.A(n_972),
.B(n_907),
.Y(n_1108)
);

BUFx2_ASAP7_75t_L g1109 ( 
.A(n_842),
.Y(n_1109)
);

AOI21xp5_ASAP7_75t_L g1110 ( 
.A1(n_975),
.A2(n_81),
.B(n_113),
.Y(n_1110)
);

O2A1O1Ixp33_ASAP7_75t_L g1111 ( 
.A1(n_1002),
.A2(n_35),
.B(n_38),
.C(n_39),
.Y(n_1111)
);

INVx1_ASAP7_75t_L g1112 ( 
.A(n_985),
.Y(n_1112)
);

INVx2_ASAP7_75t_SL g1113 ( 
.A(n_1012),
.Y(n_1113)
);

NAND2x1p5_ASAP7_75t_L g1114 ( 
.A(n_871),
.B(n_84),
.Y(n_1114)
);

INVx1_ASAP7_75t_L g1115 ( 
.A(n_1008),
.Y(n_1115)
);

NAND2xp5_ASAP7_75t_SL g1116 ( 
.A(n_979),
.B(n_121),
.Y(n_1116)
);

BUFx2_ASAP7_75t_L g1117 ( 
.A(n_842),
.Y(n_1117)
);

AND2x2_ASAP7_75t_L g1118 ( 
.A(n_888),
.B(n_35),
.Y(n_1118)
);

AOI21xp5_ASAP7_75t_L g1119 ( 
.A1(n_939),
.A2(n_99),
.B(n_97),
.Y(n_1119)
);

CKINVDCx5p33_ASAP7_75t_R g1120 ( 
.A(n_875),
.Y(n_1120)
);

AOI21xp5_ASAP7_75t_L g1121 ( 
.A1(n_844),
.A2(n_96),
.B(n_93),
.Y(n_1121)
);

INVx3_ASAP7_75t_L g1122 ( 
.A(n_910),
.Y(n_1122)
);

INVx1_ASAP7_75t_L g1123 ( 
.A(n_1013),
.Y(n_1123)
);

NAND2xp5_ASAP7_75t_SL g1124 ( 
.A(n_877),
.B(n_92),
.Y(n_1124)
);

NAND2xp5_ASAP7_75t_L g1125 ( 
.A(n_883),
.B(n_91),
.Y(n_1125)
);

CKINVDCx14_ASAP7_75t_R g1126 ( 
.A(n_873),
.Y(n_1126)
);

INVx2_ASAP7_75t_L g1127 ( 
.A(n_884),
.Y(n_1127)
);

NOR2xp33_ASAP7_75t_L g1128 ( 
.A(n_877),
.B(n_869),
.Y(n_1128)
);

BUFx12f_ASAP7_75t_L g1129 ( 
.A(n_996),
.Y(n_1129)
);

BUFx2_ASAP7_75t_L g1130 ( 
.A(n_851),
.Y(n_1130)
);

AOI21xp5_ASAP7_75t_L g1131 ( 
.A1(n_847),
.A2(n_90),
.B(n_44),
.Y(n_1131)
);

NAND2xp5_ASAP7_75t_L g1132 ( 
.A(n_1005),
.B(n_41),
.Y(n_1132)
);

INVx4_ASAP7_75t_L g1133 ( 
.A(n_910),
.Y(n_1133)
);

NAND2xp5_ASAP7_75t_L g1134 ( 
.A(n_880),
.B(n_44),
.Y(n_1134)
);

O2A1O1Ixp33_ASAP7_75t_L g1135 ( 
.A1(n_933),
.A2(n_50),
.B(n_51),
.C(n_53),
.Y(n_1135)
);

AND2x4_ASAP7_75t_L g1136 ( 
.A(n_932),
.B(n_53),
.Y(n_1136)
);

BUFx2_ASAP7_75t_L g1137 ( 
.A(n_851),
.Y(n_1137)
);

INVx1_ASAP7_75t_L g1138 ( 
.A(n_911),
.Y(n_1138)
);

CKINVDCx5p33_ASAP7_75t_R g1139 ( 
.A(n_896),
.Y(n_1139)
);

A2O1A1Ixp33_ASAP7_75t_L g1140 ( 
.A1(n_1000),
.A2(n_54),
.B(n_55),
.C(n_57),
.Y(n_1140)
);

OR2x6_ASAP7_75t_L g1141 ( 
.A(n_996),
.B(n_1019),
.Y(n_1141)
);

INVx1_ASAP7_75t_L g1142 ( 
.A(n_914),
.Y(n_1142)
);

HB1xp67_ASAP7_75t_L g1143 ( 
.A(n_890),
.Y(n_1143)
);

AND2x2_ASAP7_75t_L g1144 ( 
.A(n_892),
.B(n_54),
.Y(n_1144)
);

NOR2xp33_ASAP7_75t_R g1145 ( 
.A(n_935),
.B(n_843),
.Y(n_1145)
);

NOR3xp33_ASAP7_75t_SL g1146 ( 
.A(n_873),
.B(n_57),
.C(n_879),
.Y(n_1146)
);

NAND2xp5_ASAP7_75t_L g1147 ( 
.A(n_915),
.B(n_924),
.Y(n_1147)
);

BUFx3_ASAP7_75t_L g1148 ( 
.A(n_1012),
.Y(n_1148)
);

NOR2xp33_ASAP7_75t_L g1149 ( 
.A(n_1003),
.B(n_1019),
.Y(n_1149)
);

BUFx6f_ASAP7_75t_L g1150 ( 
.A(n_910),
.Y(n_1150)
);

A2O1A1Ixp33_ASAP7_75t_SL g1151 ( 
.A1(n_879),
.A2(n_999),
.B(n_889),
.C(n_908),
.Y(n_1151)
);

INVx1_ASAP7_75t_L g1152 ( 
.A(n_901),
.Y(n_1152)
);

AOI21xp5_ASAP7_75t_L g1153 ( 
.A1(n_993),
.A2(n_868),
.B(n_886),
.Y(n_1153)
);

BUFx2_ASAP7_75t_SL g1154 ( 
.A(n_910),
.Y(n_1154)
);

HB1xp67_ASAP7_75t_L g1155 ( 
.A(n_1019),
.Y(n_1155)
);

NOR2xp33_ASAP7_75t_L g1156 ( 
.A(n_967),
.B(n_986),
.Y(n_1156)
);

A2O1A1Ixp33_ASAP7_75t_L g1157 ( 
.A1(n_876),
.A2(n_872),
.B(n_1024),
.C(n_993),
.Y(n_1157)
);

AOI21xp5_ASAP7_75t_L g1158 ( 
.A1(n_874),
.A2(n_881),
.B(n_893),
.Y(n_1158)
);

NAND2xp5_ASAP7_75t_L g1159 ( 
.A(n_1010),
.B(n_891),
.Y(n_1159)
);

AOI22xp5_ASAP7_75t_L g1160 ( 
.A1(n_878),
.A2(n_920),
.B1(n_1026),
.B2(n_969),
.Y(n_1160)
);

AOI22xp33_ASAP7_75t_L g1161 ( 
.A1(n_920),
.A2(n_1025),
.B1(n_997),
.B2(n_1009),
.Y(n_1161)
);

INVx4_ASAP7_75t_L g1162 ( 
.A(n_916),
.Y(n_1162)
);

OAI21x1_ASAP7_75t_L g1163 ( 
.A1(n_949),
.A2(n_929),
.B(n_951),
.Y(n_1163)
);

AOI21xp5_ASAP7_75t_L g1164 ( 
.A1(n_855),
.A2(n_863),
.B(n_854),
.Y(n_1164)
);

INVx1_ASAP7_75t_L g1165 ( 
.A(n_934),
.Y(n_1165)
);

NOR2xp33_ASAP7_75t_L g1166 ( 
.A(n_903),
.B(n_940),
.Y(n_1166)
);

O2A1O1Ixp33_ASAP7_75t_L g1167 ( 
.A1(n_913),
.A2(n_983),
.B(n_1011),
.C(n_942),
.Y(n_1167)
);

OAI21x1_ASAP7_75t_SL g1168 ( 
.A1(n_991),
.A2(n_938),
.B(n_885),
.Y(n_1168)
);

NOR2xp33_ASAP7_75t_L g1169 ( 
.A(n_943),
.B(n_957),
.Y(n_1169)
);

NAND2xp5_ASAP7_75t_L g1170 ( 
.A(n_1022),
.B(n_952),
.Y(n_1170)
);

A2O1A1Ixp33_ASAP7_75t_L g1171 ( 
.A1(n_994),
.A2(n_921),
.B(n_852),
.C(n_937),
.Y(n_1171)
);

INVx3_ASAP7_75t_L g1172 ( 
.A(n_916),
.Y(n_1172)
);

NAND2xp5_ASAP7_75t_L g1173 ( 
.A(n_941),
.B(n_946),
.Y(n_1173)
);

A2O1A1Ixp33_ASAP7_75t_L g1174 ( 
.A1(n_981),
.A2(n_913),
.B(n_948),
.C(n_882),
.Y(n_1174)
);

AO21x1_ASAP7_75t_L g1175 ( 
.A1(n_882),
.A2(n_895),
.B(n_904),
.Y(n_1175)
);

O2A1O1Ixp33_ASAP7_75t_L g1176 ( 
.A1(n_895),
.A2(n_955),
.B(n_1025),
.C(n_997),
.Y(n_1176)
);

INVx2_ASAP7_75t_L g1177 ( 
.A(n_992),
.Y(n_1177)
);

OAI22xp5_ASAP7_75t_L g1178 ( 
.A1(n_950),
.A2(n_849),
.B1(n_860),
.B2(n_861),
.Y(n_1178)
);

INVx2_ASAP7_75t_L g1179 ( 
.A(n_982),
.Y(n_1179)
);

INVxp33_ASAP7_75t_SL g1180 ( 
.A(n_988),
.Y(n_1180)
);

O2A1O1Ixp33_ASAP7_75t_L g1181 ( 
.A1(n_955),
.A2(n_1016),
.B(n_1014),
.C(n_1017),
.Y(n_1181)
);

O2A1O1Ixp33_ASAP7_75t_L g1182 ( 
.A1(n_1018),
.A2(n_849),
.B(n_860),
.C(n_861),
.Y(n_1182)
);

INVx1_ASAP7_75t_L g1183 ( 
.A(n_1001),
.Y(n_1183)
);

CKINVDCx8_ASAP7_75t_R g1184 ( 
.A(n_867),
.Y(n_1184)
);

NOR2xp33_ASAP7_75t_L g1185 ( 
.A(n_961),
.B(n_945),
.Y(n_1185)
);

NAND2xp5_ASAP7_75t_L g1186 ( 
.A(n_961),
.B(n_1006),
.Y(n_1186)
);

NAND2xp5_ASAP7_75t_L g1187 ( 
.A(n_990),
.B(n_947),
.Y(n_1187)
);

OAI21x1_ASAP7_75t_L g1188 ( 
.A1(n_944),
.A2(n_962),
.B(n_964),
.Y(n_1188)
);

AOI21xp5_ASAP7_75t_L g1189 ( 
.A1(n_1049),
.A2(n_968),
.B(n_965),
.Y(n_1189)
);

AO31x2_ASAP7_75t_L g1190 ( 
.A1(n_1175),
.A2(n_1021),
.A3(n_973),
.B(n_974),
.Y(n_1190)
);

INVx5_ASAP7_75t_L g1191 ( 
.A(n_1032),
.Y(n_1191)
);

A2O1A1Ixp33_ASAP7_75t_L g1192 ( 
.A1(n_1073),
.A2(n_971),
.B(n_953),
.C(n_963),
.Y(n_1192)
);

AO31x2_ASAP7_75t_L g1193 ( 
.A1(n_1174),
.A2(n_1171),
.A3(n_1157),
.B(n_1065),
.Y(n_1193)
);

OAI22xp33_ASAP7_75t_L g1194 ( 
.A1(n_1068),
.A2(n_1030),
.B1(n_1040),
.B2(n_1028),
.Y(n_1194)
);

AND2x2_ASAP7_75t_L g1195 ( 
.A(n_1033),
.B(n_1061),
.Y(n_1195)
);

INVxp67_ASAP7_75t_L g1196 ( 
.A(n_1143),
.Y(n_1196)
);

OAI21x1_ASAP7_75t_L g1197 ( 
.A1(n_1164),
.A2(n_1057),
.B(n_1056),
.Y(n_1197)
);

BUFx6f_ASAP7_75t_L g1198 ( 
.A(n_1150),
.Y(n_1198)
);

OAI21xp5_ASAP7_75t_L g1199 ( 
.A1(n_1068),
.A2(n_1167),
.B(n_1043),
.Y(n_1199)
);

NAND3xp33_ASAP7_75t_SL g1200 ( 
.A(n_1156),
.B(n_1128),
.C(n_1146),
.Y(n_1200)
);

INVx1_ASAP7_75t_SL g1201 ( 
.A(n_1096),
.Y(n_1201)
);

A2O1A1Ixp33_ASAP7_75t_L g1202 ( 
.A1(n_1031),
.A2(n_1099),
.B(n_1049),
.C(n_1132),
.Y(n_1202)
);

OAI21xp5_ASAP7_75t_L g1203 ( 
.A1(n_1034),
.A2(n_1176),
.B(n_1099),
.Y(n_1203)
);

OAI21x1_ASAP7_75t_L g1204 ( 
.A1(n_1074),
.A2(n_1153),
.B(n_1029),
.Y(n_1204)
);

CKINVDCx16_ASAP7_75t_R g1205 ( 
.A(n_1145),
.Y(n_1205)
);

OAI21x1_ASAP7_75t_L g1206 ( 
.A1(n_1059),
.A2(n_1037),
.B(n_1053),
.Y(n_1206)
);

INVxp67_ASAP7_75t_L g1207 ( 
.A(n_1042),
.Y(n_1207)
);

NAND2xp5_ASAP7_75t_SL g1208 ( 
.A(n_1180),
.B(n_1076),
.Y(n_1208)
);

AO31x2_ASAP7_75t_L g1209 ( 
.A1(n_1065),
.A2(n_1070),
.A3(n_1178),
.B(n_1077),
.Y(n_1209)
);

OAI21x1_ASAP7_75t_L g1210 ( 
.A1(n_1187),
.A2(n_1188),
.B(n_1078),
.Y(n_1210)
);

NAND2xp5_ASAP7_75t_SL g1211 ( 
.A(n_1094),
.B(n_1069),
.Y(n_1211)
);

OAI22xp5_ASAP7_75t_L g1212 ( 
.A1(n_1147),
.A2(n_1138),
.B1(n_1142),
.B2(n_1058),
.Y(n_1212)
);

O2A1O1Ixp33_ASAP7_75t_L g1213 ( 
.A1(n_1104),
.A2(n_1140),
.B(n_1103),
.C(n_1077),
.Y(n_1213)
);

NAND2xp5_ASAP7_75t_L g1214 ( 
.A(n_1147),
.B(n_1179),
.Y(n_1214)
);

NAND2xp5_ASAP7_75t_L g1215 ( 
.A(n_1170),
.B(n_1159),
.Y(n_1215)
);

AOI21xp5_ASAP7_75t_L g1216 ( 
.A1(n_1185),
.A2(n_1186),
.B(n_1187),
.Y(n_1216)
);

OAI22xp5_ASAP7_75t_L g1217 ( 
.A1(n_1159),
.A2(n_1095),
.B1(n_1048),
.B2(n_1060),
.Y(n_1217)
);

A2O1A1Ixp33_ASAP7_75t_L g1218 ( 
.A1(n_1131),
.A2(n_1134),
.B(n_1160),
.C(n_1166),
.Y(n_1218)
);

BUFx3_ASAP7_75t_L g1219 ( 
.A(n_1129),
.Y(n_1219)
);

A2O1A1Ixp33_ASAP7_75t_L g1220 ( 
.A1(n_1107),
.A2(n_1125),
.B(n_1084),
.C(n_1085),
.Y(n_1220)
);

BUFx6f_ASAP7_75t_L g1221 ( 
.A(n_1150),
.Y(n_1221)
);

INVx1_ASAP7_75t_L g1222 ( 
.A(n_1051),
.Y(n_1222)
);

AND2x4_ASAP7_75t_L g1223 ( 
.A(n_1071),
.B(n_1072),
.Y(n_1223)
);

O2A1O1Ixp33_ASAP7_75t_SL g1224 ( 
.A1(n_1151),
.A2(n_1124),
.B(n_1116),
.C(n_1100),
.Y(n_1224)
);

OAI21xp5_ASAP7_75t_L g1225 ( 
.A1(n_1050),
.A2(n_1080),
.B(n_1125),
.Y(n_1225)
);

AOI21xp5_ASAP7_75t_L g1226 ( 
.A1(n_1173),
.A2(n_1062),
.B(n_1063),
.Y(n_1226)
);

BUFx2_ASAP7_75t_L g1227 ( 
.A(n_1109),
.Y(n_1227)
);

OAI22xp5_ASAP7_75t_L g1228 ( 
.A1(n_1055),
.A2(n_1112),
.B1(n_1090),
.B2(n_1028),
.Y(n_1228)
);

AOI21xp5_ASAP7_75t_L g1229 ( 
.A1(n_1062),
.A2(n_1181),
.B(n_1183),
.Y(n_1229)
);

OAI21x1_ASAP7_75t_L g1230 ( 
.A1(n_1064),
.A2(n_1078),
.B(n_1066),
.Y(n_1230)
);

A2O1A1Ixp33_ASAP7_75t_L g1231 ( 
.A1(n_1182),
.A2(n_1135),
.B(n_1083),
.C(n_1121),
.Y(n_1231)
);

INVx1_ASAP7_75t_L g1232 ( 
.A(n_1115),
.Y(n_1232)
);

NAND2xp5_ASAP7_75t_L g1233 ( 
.A(n_1102),
.B(n_1169),
.Y(n_1233)
);

BUFx6f_ASAP7_75t_L g1234 ( 
.A(n_1150),
.Y(n_1234)
);

A2O1A1Ixp33_ASAP7_75t_L g1235 ( 
.A1(n_1161),
.A2(n_1110),
.B(n_1093),
.C(n_1111),
.Y(n_1235)
);

NAND2xp5_ASAP7_75t_L g1236 ( 
.A(n_1123),
.B(n_1072),
.Y(n_1236)
);

INVx2_ASAP7_75t_L g1237 ( 
.A(n_1106),
.Y(n_1237)
);

INVx3_ASAP7_75t_L g1238 ( 
.A(n_1162),
.Y(n_1238)
);

AOI221x1_ASAP7_75t_L g1239 ( 
.A1(n_1103),
.A2(n_1168),
.B1(n_1178),
.B2(n_1035),
.C(n_1119),
.Y(n_1239)
);

NAND2xp5_ASAP7_75t_L g1240 ( 
.A(n_1118),
.B(n_1108),
.Y(n_1240)
);

O2A1O1Ixp33_ASAP7_75t_SL g1241 ( 
.A1(n_1101),
.A2(n_1041),
.B(n_1088),
.C(n_1044),
.Y(n_1241)
);

OAI21x1_ASAP7_75t_L g1242 ( 
.A1(n_1064),
.A2(n_1066),
.B(n_1177),
.Y(n_1242)
);

OAI21x1_ASAP7_75t_L g1243 ( 
.A1(n_1046),
.A2(n_1047),
.B(n_1054),
.Y(n_1243)
);

AOI21xp5_ASAP7_75t_L g1244 ( 
.A1(n_1075),
.A2(n_1081),
.B(n_1067),
.Y(n_1244)
);

INVx2_ASAP7_75t_L g1245 ( 
.A(n_1127),
.Y(n_1245)
);

AOI21xp5_ASAP7_75t_L g1246 ( 
.A1(n_1092),
.A2(n_1045),
.B(n_1047),
.Y(n_1246)
);

AOI21xp5_ASAP7_75t_L g1247 ( 
.A1(n_1046),
.A2(n_1086),
.B(n_1087),
.Y(n_1247)
);

NOR2xp67_ASAP7_75t_L g1248 ( 
.A(n_1039),
.B(n_1113),
.Y(n_1248)
);

OA21x2_ASAP7_75t_L g1249 ( 
.A1(n_1082),
.A2(n_1165),
.B(n_1152),
.Y(n_1249)
);

AND2x2_ASAP7_75t_L g1250 ( 
.A(n_1144),
.B(n_1137),
.Y(n_1250)
);

A2O1A1Ixp33_ASAP7_75t_L g1251 ( 
.A1(n_1149),
.A2(n_1155),
.B(n_1108),
.C(n_1172),
.Y(n_1251)
);

NAND3xp33_ASAP7_75t_L g1252 ( 
.A(n_1126),
.B(n_1028),
.C(n_1136),
.Y(n_1252)
);

AOI22xp5_ASAP7_75t_L g1253 ( 
.A1(n_1139),
.A2(n_1141),
.B1(n_1117),
.B2(n_1130),
.Y(n_1253)
);

AND2x2_ASAP7_75t_L g1254 ( 
.A(n_1136),
.B(n_1098),
.Y(n_1254)
);

AND2x2_ASAP7_75t_L g1255 ( 
.A(n_1141),
.B(n_1148),
.Y(n_1255)
);

NOR2xp67_ASAP7_75t_L g1256 ( 
.A(n_1097),
.B(n_1105),
.Y(n_1256)
);

CKINVDCx5p33_ASAP7_75t_R g1257 ( 
.A(n_1052),
.Y(n_1257)
);

BUFx3_ASAP7_75t_L g1258 ( 
.A(n_1141),
.Y(n_1258)
);

NAND2xp5_ASAP7_75t_L g1259 ( 
.A(n_1091),
.B(n_1089),
.Y(n_1259)
);

AOI21xp5_ASAP7_75t_L g1260 ( 
.A1(n_1054),
.A2(n_1079),
.B(n_1122),
.Y(n_1260)
);

INVx2_ASAP7_75t_L g1261 ( 
.A(n_1091),
.Y(n_1261)
);

O2A1O1Ixp5_ASAP7_75t_SL g1262 ( 
.A1(n_1036),
.A2(n_1038),
.B(n_1079),
.C(n_1122),
.Y(n_1262)
);

INVx1_ASAP7_75t_L g1263 ( 
.A(n_1036),
.Y(n_1263)
);

OR2x2_ASAP7_75t_L g1264 ( 
.A(n_1089),
.B(n_1154),
.Y(n_1264)
);

INVx1_ASAP7_75t_SL g1265 ( 
.A(n_1089),
.Y(n_1265)
);

OAI22x1_ASAP7_75t_L g1266 ( 
.A1(n_1114),
.A2(n_1097),
.B1(n_1133),
.B2(n_1038),
.Y(n_1266)
);

AOI21xp5_ASAP7_75t_L g1267 ( 
.A1(n_1114),
.A2(n_1032),
.B(n_1091),
.Y(n_1267)
);

AOI221xp5_ASAP7_75t_SL g1268 ( 
.A1(n_1032),
.A2(n_1068),
.B1(n_1077),
.B2(n_1073),
.C(n_1020),
.Y(n_1268)
);

AND2x2_ASAP7_75t_L g1269 ( 
.A(n_1184),
.B(n_1120),
.Y(n_1269)
);

OAI21x1_ASAP7_75t_SL g1270 ( 
.A1(n_1091),
.A2(n_1168),
.B(n_1035),
.Y(n_1270)
);

NAND2xp5_ASAP7_75t_L g1271 ( 
.A(n_1068),
.B(n_1049),
.Y(n_1271)
);

AOI21xp5_ASAP7_75t_L g1272 ( 
.A1(n_1049),
.A2(n_681),
.B(n_837),
.Y(n_1272)
);

INVx2_ASAP7_75t_SL g1273 ( 
.A(n_1148),
.Y(n_1273)
);

NAND2xp5_ASAP7_75t_L g1274 ( 
.A(n_1068),
.B(n_1049),
.Y(n_1274)
);

NOR2xp33_ASAP7_75t_L g1275 ( 
.A(n_1061),
.B(n_681),
.Y(n_1275)
);

AO31x2_ASAP7_75t_L g1276 ( 
.A1(n_1175),
.A2(n_1174),
.A3(n_1171),
.B(n_991),
.Y(n_1276)
);

INVx4_ASAP7_75t_L g1277 ( 
.A(n_1150),
.Y(n_1277)
);

BUFx8_ASAP7_75t_L g1278 ( 
.A(n_1129),
.Y(n_1278)
);

NAND2xp5_ASAP7_75t_L g1279 ( 
.A(n_1068),
.B(n_1049),
.Y(n_1279)
);

AOI221x1_ASAP7_75t_L g1280 ( 
.A1(n_1077),
.A2(n_958),
.B1(n_1065),
.B2(n_1068),
.C(n_681),
.Y(n_1280)
);

BUFx2_ASAP7_75t_L g1281 ( 
.A(n_1042),
.Y(n_1281)
);

AND2x2_ASAP7_75t_L g1282 ( 
.A(n_1033),
.B(n_1061),
.Y(n_1282)
);

AO31x2_ASAP7_75t_L g1283 ( 
.A1(n_1175),
.A2(n_1174),
.A3(n_1171),
.B(n_991),
.Y(n_1283)
);

OAI22xp5_ASAP7_75t_L g1284 ( 
.A1(n_1068),
.A2(n_681),
.B1(n_1049),
.B2(n_760),
.Y(n_1284)
);

AND2x4_ASAP7_75t_L g1285 ( 
.A(n_1071),
.B(n_1072),
.Y(n_1285)
);

INVx2_ASAP7_75t_L g1286 ( 
.A(n_1048),
.Y(n_1286)
);

CKINVDCx5p33_ASAP7_75t_R g1287 ( 
.A(n_1039),
.Y(n_1287)
);

NAND2xp5_ASAP7_75t_L g1288 ( 
.A(n_1068),
.B(n_681),
.Y(n_1288)
);

AOI21xp5_ASAP7_75t_L g1289 ( 
.A1(n_1049),
.A2(n_681),
.B(n_837),
.Y(n_1289)
);

INVx3_ASAP7_75t_L g1290 ( 
.A(n_1071),
.Y(n_1290)
);

BUFx3_ASAP7_75t_L g1291 ( 
.A(n_1076),
.Y(n_1291)
);

NAND3x1_ASAP7_75t_L g1292 ( 
.A(n_1156),
.B(n_577),
.C(n_500),
.Y(n_1292)
);

AOI21xp5_ASAP7_75t_L g1293 ( 
.A1(n_1049),
.A2(n_681),
.B(n_837),
.Y(n_1293)
);

NAND2xp5_ASAP7_75t_L g1294 ( 
.A(n_1068),
.B(n_681),
.Y(n_1294)
);

OAI21x1_ASAP7_75t_L g1295 ( 
.A1(n_1163),
.A2(n_1158),
.B(n_1164),
.Y(n_1295)
);

NAND2xp33_ASAP7_75t_L g1296 ( 
.A(n_1068),
.B(n_681),
.Y(n_1296)
);

CKINVDCx5p33_ASAP7_75t_R g1297 ( 
.A(n_1039),
.Y(n_1297)
);

AO21x1_ASAP7_75t_L g1298 ( 
.A1(n_1073),
.A2(n_1068),
.B(n_1099),
.Y(n_1298)
);

OAI21x1_ASAP7_75t_L g1299 ( 
.A1(n_1163),
.A2(n_1158),
.B(n_1164),
.Y(n_1299)
);

INVxp67_ASAP7_75t_SL g1300 ( 
.A(n_1049),
.Y(n_1300)
);

AOI21xp5_ASAP7_75t_L g1301 ( 
.A1(n_1049),
.A2(n_681),
.B(n_837),
.Y(n_1301)
);

NAND3xp33_ASAP7_75t_SL g1302 ( 
.A(n_1061),
.B(n_681),
.C(n_853),
.Y(n_1302)
);

AO31x2_ASAP7_75t_L g1303 ( 
.A1(n_1175),
.A2(n_1174),
.A3(n_1171),
.B(n_991),
.Y(n_1303)
);

AO22x2_ASAP7_75t_L g1304 ( 
.A1(n_1077),
.A2(n_1068),
.B1(n_1065),
.B2(n_1030),
.Y(n_1304)
);

AOI221x1_ASAP7_75t_L g1305 ( 
.A1(n_1077),
.A2(n_958),
.B1(n_1065),
.B2(n_1068),
.C(n_681),
.Y(n_1305)
);

NOR2xp33_ASAP7_75t_L g1306 ( 
.A(n_1061),
.B(n_681),
.Y(n_1306)
);

NAND2x1p5_ASAP7_75t_L g1307 ( 
.A(n_1097),
.B(n_859),
.Y(n_1307)
);

INVx1_ASAP7_75t_L g1308 ( 
.A(n_1048),
.Y(n_1308)
);

NAND2xp5_ASAP7_75t_L g1309 ( 
.A(n_1068),
.B(n_681),
.Y(n_1309)
);

OAI21x1_ASAP7_75t_L g1310 ( 
.A1(n_1163),
.A2(n_1158),
.B(n_1164),
.Y(n_1310)
);

NAND2xp5_ASAP7_75t_L g1311 ( 
.A(n_1068),
.B(n_1049),
.Y(n_1311)
);

AND2x2_ASAP7_75t_L g1312 ( 
.A(n_1033),
.B(n_1061),
.Y(n_1312)
);

CKINVDCx5p33_ASAP7_75t_R g1313 ( 
.A(n_1039),
.Y(n_1313)
);

OAI21x1_ASAP7_75t_L g1314 ( 
.A1(n_1163),
.A2(n_1158),
.B(n_1164),
.Y(n_1314)
);

NAND2xp5_ASAP7_75t_L g1315 ( 
.A(n_1068),
.B(n_1049),
.Y(n_1315)
);

AO31x2_ASAP7_75t_L g1316 ( 
.A1(n_1175),
.A2(n_1174),
.A3(n_1171),
.B(n_991),
.Y(n_1316)
);

NOR2xp33_ASAP7_75t_L g1317 ( 
.A(n_1061),
.B(n_681),
.Y(n_1317)
);

OAI22xp5_ASAP7_75t_L g1318 ( 
.A1(n_1068),
.A2(n_681),
.B1(n_1049),
.B2(n_760),
.Y(n_1318)
);

OAI22xp5_ASAP7_75t_L g1319 ( 
.A1(n_1068),
.A2(n_681),
.B1(n_1049),
.B2(n_760),
.Y(n_1319)
);

NAND3xp33_ASAP7_75t_SL g1320 ( 
.A(n_1061),
.B(n_681),
.C(n_853),
.Y(n_1320)
);

OAI22xp5_ASAP7_75t_L g1321 ( 
.A1(n_1068),
.A2(n_681),
.B1(n_1049),
.B2(n_760),
.Y(n_1321)
);

A2O1A1Ixp33_ASAP7_75t_L g1322 ( 
.A1(n_1073),
.A2(n_681),
.B(n_958),
.C(n_1068),
.Y(n_1322)
);

NOR4xp25_ASAP7_75t_L g1323 ( 
.A(n_1073),
.B(n_958),
.C(n_1068),
.D(n_1111),
.Y(n_1323)
);

A2O1A1Ixp33_ASAP7_75t_L g1324 ( 
.A1(n_1073),
.A2(n_681),
.B(n_958),
.C(n_1068),
.Y(n_1324)
);

NAND2xp5_ASAP7_75t_L g1325 ( 
.A(n_1068),
.B(n_681),
.Y(n_1325)
);

INVxp67_ASAP7_75t_SL g1326 ( 
.A(n_1049),
.Y(n_1326)
);

INVxp67_ASAP7_75t_L g1327 ( 
.A(n_1033),
.Y(n_1327)
);

BUFx12f_ASAP7_75t_L g1328 ( 
.A(n_1120),
.Y(n_1328)
);

OAI21x1_ASAP7_75t_L g1329 ( 
.A1(n_1163),
.A2(n_1158),
.B(n_1164),
.Y(n_1329)
);

A2O1A1Ixp33_ASAP7_75t_L g1330 ( 
.A1(n_1073),
.A2(n_681),
.B(n_958),
.C(n_1068),
.Y(n_1330)
);

OR2x6_ASAP7_75t_L g1331 ( 
.A(n_1154),
.B(n_1089),
.Y(n_1331)
);

CKINVDCx20_ASAP7_75t_R g1332 ( 
.A(n_1052),
.Y(n_1332)
);

AOI21xp5_ASAP7_75t_L g1333 ( 
.A1(n_1049),
.A2(n_681),
.B(n_837),
.Y(n_1333)
);

INVx3_ASAP7_75t_L g1334 ( 
.A(n_1071),
.Y(n_1334)
);

AOI21xp5_ASAP7_75t_L g1335 ( 
.A1(n_1049),
.A2(n_681),
.B(n_837),
.Y(n_1335)
);

A2O1A1Ixp33_ASAP7_75t_L g1336 ( 
.A1(n_1073),
.A2(n_681),
.B(n_958),
.C(n_1068),
.Y(n_1336)
);

AOI22xp5_ASAP7_75t_L g1337 ( 
.A1(n_1061),
.A2(n_853),
.B1(n_681),
.B2(n_977),
.Y(n_1337)
);

NOR2xp33_ASAP7_75t_SL g1338 ( 
.A(n_1068),
.B(n_619),
.Y(n_1338)
);

AOI21xp5_ASAP7_75t_L g1339 ( 
.A1(n_1049),
.A2(n_681),
.B(n_837),
.Y(n_1339)
);

A2O1A1Ixp33_ASAP7_75t_L g1340 ( 
.A1(n_1073),
.A2(n_681),
.B(n_958),
.C(n_1068),
.Y(n_1340)
);

AND2x4_ASAP7_75t_L g1341 ( 
.A(n_1071),
.B(n_1072),
.Y(n_1341)
);

OAI21x1_ASAP7_75t_L g1342 ( 
.A1(n_1163),
.A2(n_1158),
.B(n_1164),
.Y(n_1342)
);

AOI22xp33_ASAP7_75t_L g1343 ( 
.A1(n_1156),
.A2(n_681),
.B1(n_977),
.B2(n_686),
.Y(n_1343)
);

OAI21xp5_ASAP7_75t_L g1344 ( 
.A1(n_1073),
.A2(n_958),
.B(n_1068),
.Y(n_1344)
);

NAND3xp33_ASAP7_75t_L g1345 ( 
.A(n_1073),
.B(n_681),
.C(n_977),
.Y(n_1345)
);

INVx6_ASAP7_75t_L g1346 ( 
.A(n_1191),
.Y(n_1346)
);

AOI22xp5_ASAP7_75t_L g1347 ( 
.A1(n_1337),
.A2(n_1343),
.B1(n_1320),
.B2(n_1302),
.Y(n_1347)
);

AOI22xp33_ASAP7_75t_L g1348 ( 
.A1(n_1345),
.A2(n_1296),
.B1(n_1200),
.B2(n_1344),
.Y(n_1348)
);

AOI22xp33_ASAP7_75t_L g1349 ( 
.A1(n_1345),
.A2(n_1344),
.B1(n_1317),
.B2(n_1275),
.Y(n_1349)
);

AOI22xp33_ASAP7_75t_L g1350 ( 
.A1(n_1306),
.A2(n_1298),
.B1(n_1194),
.B2(n_1199),
.Y(n_1350)
);

HB1xp67_ASAP7_75t_L g1351 ( 
.A(n_1261),
.Y(n_1351)
);

AOI22xp33_ASAP7_75t_L g1352 ( 
.A1(n_1199),
.A2(n_1294),
.B1(n_1309),
.B2(n_1325),
.Y(n_1352)
);

CKINVDCx6p67_ASAP7_75t_R g1353 ( 
.A(n_1328),
.Y(n_1353)
);

BUFx3_ASAP7_75t_L g1354 ( 
.A(n_1291),
.Y(n_1354)
);

INVx6_ASAP7_75t_L g1355 ( 
.A(n_1191),
.Y(n_1355)
);

AOI22xp33_ASAP7_75t_L g1356 ( 
.A1(n_1288),
.A2(n_1304),
.B1(n_1338),
.B2(n_1319),
.Y(n_1356)
);

CKINVDCx11_ASAP7_75t_R g1357 ( 
.A(n_1332),
.Y(n_1357)
);

CKINVDCx5p33_ASAP7_75t_R g1358 ( 
.A(n_1287),
.Y(n_1358)
);

AOI22xp33_ASAP7_75t_SL g1359 ( 
.A1(n_1338),
.A2(n_1284),
.B1(n_1318),
.B2(n_1319),
.Y(n_1359)
);

CKINVDCx11_ASAP7_75t_R g1360 ( 
.A(n_1205),
.Y(n_1360)
);

AND2x2_ASAP7_75t_L g1361 ( 
.A(n_1195),
.B(n_1282),
.Y(n_1361)
);

AOI22xp33_ASAP7_75t_L g1362 ( 
.A1(n_1304),
.A2(n_1321),
.B1(n_1284),
.B2(n_1318),
.Y(n_1362)
);

BUFx3_ASAP7_75t_L g1363 ( 
.A(n_1227),
.Y(n_1363)
);

INVx2_ASAP7_75t_L g1364 ( 
.A(n_1237),
.Y(n_1364)
);

AOI22xp5_ASAP7_75t_L g1365 ( 
.A1(n_1292),
.A2(n_1312),
.B1(n_1211),
.B2(n_1254),
.Y(n_1365)
);

AOI22xp33_ASAP7_75t_L g1366 ( 
.A1(n_1321),
.A2(n_1203),
.B1(n_1212),
.B2(n_1215),
.Y(n_1366)
);

AOI22xp5_ASAP7_75t_SL g1367 ( 
.A1(n_1327),
.A2(n_1233),
.B1(n_1228),
.B2(n_1258),
.Y(n_1367)
);

INVx1_ASAP7_75t_L g1368 ( 
.A(n_1222),
.Y(n_1368)
);

AOI22xp33_ASAP7_75t_L g1369 ( 
.A1(n_1203),
.A2(n_1212),
.B1(n_1274),
.B2(n_1315),
.Y(n_1369)
);

INVx2_ASAP7_75t_L g1370 ( 
.A(n_1245),
.Y(n_1370)
);

BUFx8_ASAP7_75t_SL g1371 ( 
.A(n_1257),
.Y(n_1371)
);

OAI22xp5_ASAP7_75t_L g1372 ( 
.A1(n_1300),
.A2(n_1326),
.B1(n_1274),
.B2(n_1311),
.Y(n_1372)
);

BUFx3_ASAP7_75t_L g1373 ( 
.A(n_1281),
.Y(n_1373)
);

NAND2xp5_ASAP7_75t_L g1374 ( 
.A(n_1214),
.B(n_1271),
.Y(n_1374)
);

INVx2_ASAP7_75t_L g1375 ( 
.A(n_1308),
.Y(n_1375)
);

AOI22xp33_ASAP7_75t_L g1376 ( 
.A1(n_1271),
.A2(n_1311),
.B1(n_1315),
.B2(n_1279),
.Y(n_1376)
);

CKINVDCx6p67_ASAP7_75t_R g1377 ( 
.A(n_1219),
.Y(n_1377)
);

BUFx6f_ASAP7_75t_L g1378 ( 
.A(n_1198),
.Y(n_1378)
);

OAI22xp33_ASAP7_75t_L g1379 ( 
.A1(n_1280),
.A2(n_1305),
.B1(n_1279),
.B2(n_1252),
.Y(n_1379)
);

INVx1_ASAP7_75t_L g1380 ( 
.A(n_1232),
.Y(n_1380)
);

CKINVDCx12_ASAP7_75t_R g1381 ( 
.A(n_1269),
.Y(n_1381)
);

INVx6_ASAP7_75t_L g1382 ( 
.A(n_1331),
.Y(n_1382)
);

NAND2x1p5_ASAP7_75t_L g1383 ( 
.A(n_1238),
.B(n_1265),
.Y(n_1383)
);

INVx2_ASAP7_75t_L g1384 ( 
.A(n_1249),
.Y(n_1384)
);

AOI22xp33_ASAP7_75t_L g1385 ( 
.A1(n_1217),
.A2(n_1252),
.B1(n_1228),
.B2(n_1250),
.Y(n_1385)
);

OAI22xp5_ASAP7_75t_L g1386 ( 
.A1(n_1322),
.A2(n_1324),
.B1(n_1340),
.B2(n_1330),
.Y(n_1386)
);

OAI22xp5_ASAP7_75t_L g1387 ( 
.A1(n_1336),
.A2(n_1208),
.B1(n_1240),
.B2(n_1236),
.Y(n_1387)
);

BUFx12f_ASAP7_75t_L g1388 ( 
.A(n_1278),
.Y(n_1388)
);

AOI22xp33_ASAP7_75t_L g1389 ( 
.A1(n_1217),
.A2(n_1333),
.B1(n_1301),
.B2(n_1339),
.Y(n_1389)
);

INVx1_ASAP7_75t_L g1390 ( 
.A(n_1263),
.Y(n_1390)
);

AOI22xp33_ASAP7_75t_SL g1391 ( 
.A1(n_1216),
.A2(n_1213),
.B1(n_1193),
.B2(n_1268),
.Y(n_1391)
);

CKINVDCx5p33_ASAP7_75t_R g1392 ( 
.A(n_1297),
.Y(n_1392)
);

INVx6_ASAP7_75t_L g1393 ( 
.A(n_1331),
.Y(n_1393)
);

INVx2_ASAP7_75t_R g1394 ( 
.A(n_1193),
.Y(n_1394)
);

CKINVDCx5p33_ASAP7_75t_R g1395 ( 
.A(n_1313),
.Y(n_1395)
);

BUFx8_ASAP7_75t_SL g1396 ( 
.A(n_1255),
.Y(n_1396)
);

AOI22xp5_ASAP7_75t_L g1397 ( 
.A1(n_1223),
.A2(n_1341),
.B1(n_1285),
.B2(n_1253),
.Y(n_1397)
);

INVx1_ASAP7_75t_SL g1398 ( 
.A(n_1201),
.Y(n_1398)
);

CKINVDCx5p33_ASAP7_75t_R g1399 ( 
.A(n_1278),
.Y(n_1399)
);

OAI22xp5_ASAP7_75t_L g1400 ( 
.A1(n_1251),
.A2(n_1207),
.B1(n_1202),
.B2(n_1201),
.Y(n_1400)
);

BUFx3_ASAP7_75t_L g1401 ( 
.A(n_1273),
.Y(n_1401)
);

HB1xp67_ASAP7_75t_SL g1402 ( 
.A(n_1223),
.Y(n_1402)
);

BUFx12f_ASAP7_75t_L g1403 ( 
.A(n_1198),
.Y(n_1403)
);

AOI22xp33_ASAP7_75t_L g1404 ( 
.A1(n_1272),
.A2(n_1293),
.B1(n_1289),
.B2(n_1335),
.Y(n_1404)
);

OAI22xp5_ASAP7_75t_L g1405 ( 
.A1(n_1196),
.A2(n_1218),
.B1(n_1341),
.B2(n_1285),
.Y(n_1405)
);

BUFx6f_ASAP7_75t_L g1406 ( 
.A(n_1198),
.Y(n_1406)
);

INVx6_ASAP7_75t_L g1407 ( 
.A(n_1277),
.Y(n_1407)
);

AOI22xp33_ASAP7_75t_SL g1408 ( 
.A1(n_1193),
.A2(n_1268),
.B1(n_1246),
.B2(n_1323),
.Y(n_1408)
);

BUFx2_ASAP7_75t_SL g1409 ( 
.A(n_1248),
.Y(n_1409)
);

BUFx2_ASAP7_75t_L g1410 ( 
.A(n_1221),
.Y(n_1410)
);

INVx6_ASAP7_75t_L g1411 ( 
.A(n_1277),
.Y(n_1411)
);

NAND2xp5_ASAP7_75t_L g1412 ( 
.A(n_1290),
.B(n_1334),
.Y(n_1412)
);

BUFx10_ASAP7_75t_L g1413 ( 
.A(n_1221),
.Y(n_1413)
);

INVx1_ASAP7_75t_L g1414 ( 
.A(n_1221),
.Y(n_1414)
);

AOI22xp5_ASAP7_75t_L g1415 ( 
.A1(n_1290),
.A2(n_1334),
.B1(n_1241),
.B2(n_1265),
.Y(n_1415)
);

AOI22xp33_ASAP7_75t_L g1416 ( 
.A1(n_1226),
.A2(n_1225),
.B1(n_1229),
.B2(n_1247),
.Y(n_1416)
);

BUFx6f_ASAP7_75t_L g1417 ( 
.A(n_1234),
.Y(n_1417)
);

CKINVDCx14_ASAP7_75t_R g1418 ( 
.A(n_1264),
.Y(n_1418)
);

CKINVDCx5p33_ASAP7_75t_R g1419 ( 
.A(n_1234),
.Y(n_1419)
);

NAND2xp5_ASAP7_75t_L g1420 ( 
.A(n_1259),
.B(n_1220),
.Y(n_1420)
);

AOI22xp33_ASAP7_75t_SL g1421 ( 
.A1(n_1209),
.A2(n_1230),
.B1(n_1243),
.B2(n_1238),
.Y(n_1421)
);

OAI22xp5_ASAP7_75t_L g1422 ( 
.A1(n_1231),
.A2(n_1235),
.B1(n_1267),
.B2(n_1256),
.Y(n_1422)
);

INVx1_ASAP7_75t_L g1423 ( 
.A(n_1234),
.Y(n_1423)
);

INVx2_ASAP7_75t_L g1424 ( 
.A(n_1307),
.Y(n_1424)
);

BUFx10_ASAP7_75t_L g1425 ( 
.A(n_1266),
.Y(n_1425)
);

AOI22xp33_ASAP7_75t_L g1426 ( 
.A1(n_1270),
.A2(n_1210),
.B1(n_1244),
.B2(n_1242),
.Y(n_1426)
);

INVx6_ASAP7_75t_L g1427 ( 
.A(n_1260),
.Y(n_1427)
);

AOI22xp33_ASAP7_75t_L g1428 ( 
.A1(n_1209),
.A2(n_1189),
.B1(n_1206),
.B2(n_1197),
.Y(n_1428)
);

AOI22xp33_ASAP7_75t_L g1429 ( 
.A1(n_1204),
.A2(n_1239),
.B1(n_1342),
.B2(n_1299),
.Y(n_1429)
);

AOI22xp33_ASAP7_75t_SL g1430 ( 
.A1(n_1224),
.A2(n_1316),
.B1(n_1303),
.B2(n_1283),
.Y(n_1430)
);

BUFx2_ASAP7_75t_SL g1431 ( 
.A(n_1262),
.Y(n_1431)
);

OR2x2_ASAP7_75t_L g1432 ( 
.A(n_1276),
.B(n_1303),
.Y(n_1432)
);

AOI22xp33_ASAP7_75t_L g1433 ( 
.A1(n_1295),
.A2(n_1329),
.B1(n_1314),
.B2(n_1310),
.Y(n_1433)
);

INVx1_ASAP7_75t_L g1434 ( 
.A(n_1283),
.Y(n_1434)
);

CKINVDCx11_ASAP7_75t_R g1435 ( 
.A(n_1283),
.Y(n_1435)
);

INVxp67_ASAP7_75t_L g1436 ( 
.A(n_1192),
.Y(n_1436)
);

CKINVDCx11_ASAP7_75t_R g1437 ( 
.A(n_1303),
.Y(n_1437)
);

BUFx12f_ASAP7_75t_L g1438 ( 
.A(n_1316),
.Y(n_1438)
);

CKINVDCx20_ASAP7_75t_R g1439 ( 
.A(n_1316),
.Y(n_1439)
);

INVx1_ASAP7_75t_SL g1440 ( 
.A(n_1190),
.Y(n_1440)
);

CKINVDCx6p67_ASAP7_75t_R g1441 ( 
.A(n_1190),
.Y(n_1441)
);

BUFx3_ASAP7_75t_L g1442 ( 
.A(n_1190),
.Y(n_1442)
);

INVx6_ASAP7_75t_L g1443 ( 
.A(n_1191),
.Y(n_1443)
);

AOI22xp5_ASAP7_75t_L g1444 ( 
.A1(n_1337),
.A2(n_853),
.B1(n_850),
.B2(n_681),
.Y(n_1444)
);

NAND2xp5_ASAP7_75t_L g1445 ( 
.A(n_1275),
.B(n_1306),
.Y(n_1445)
);

CKINVDCx11_ASAP7_75t_R g1446 ( 
.A(n_1328),
.Y(n_1446)
);

AOI22xp33_ASAP7_75t_L g1447 ( 
.A1(n_1343),
.A2(n_1068),
.B1(n_1345),
.B2(n_1320),
.Y(n_1447)
);

CKINVDCx11_ASAP7_75t_R g1448 ( 
.A(n_1328),
.Y(n_1448)
);

AOI22xp33_ASAP7_75t_L g1449 ( 
.A1(n_1343),
.A2(n_1068),
.B1(n_1345),
.B2(n_1320),
.Y(n_1449)
);

INVx1_ASAP7_75t_L g1450 ( 
.A(n_1286),
.Y(n_1450)
);

OAI22xp5_ASAP7_75t_L g1451 ( 
.A1(n_1343),
.A2(n_681),
.B1(n_1337),
.B2(n_1068),
.Y(n_1451)
);

BUFx3_ASAP7_75t_L g1452 ( 
.A(n_1291),
.Y(n_1452)
);

CKINVDCx6p67_ASAP7_75t_R g1453 ( 
.A(n_1328),
.Y(n_1453)
);

INVx1_ASAP7_75t_L g1454 ( 
.A(n_1286),
.Y(n_1454)
);

AOI22xp33_ASAP7_75t_SL g1455 ( 
.A1(n_1338),
.A2(n_359),
.B1(n_369),
.B2(n_356),
.Y(n_1455)
);

INVx6_ASAP7_75t_L g1456 ( 
.A(n_1191),
.Y(n_1456)
);

AOI22xp33_ASAP7_75t_L g1457 ( 
.A1(n_1343),
.A2(n_1068),
.B1(n_1345),
.B2(n_1320),
.Y(n_1457)
);

AOI22xp33_ASAP7_75t_L g1458 ( 
.A1(n_1343),
.A2(n_1068),
.B1(n_1345),
.B2(n_1320),
.Y(n_1458)
);

INVx1_ASAP7_75t_L g1459 ( 
.A(n_1286),
.Y(n_1459)
);

CKINVDCx9p33_ASAP7_75t_R g1460 ( 
.A(n_1275),
.Y(n_1460)
);

BUFx10_ASAP7_75t_L g1461 ( 
.A(n_1287),
.Y(n_1461)
);

INVx2_ASAP7_75t_SL g1462 ( 
.A(n_1291),
.Y(n_1462)
);

INVx6_ASAP7_75t_L g1463 ( 
.A(n_1191),
.Y(n_1463)
);

BUFx6f_ASAP7_75t_L g1464 ( 
.A(n_1191),
.Y(n_1464)
);

OAI22xp5_ASAP7_75t_L g1465 ( 
.A1(n_1343),
.A2(n_681),
.B1(n_1337),
.B2(n_1068),
.Y(n_1465)
);

CKINVDCx5p33_ASAP7_75t_R g1466 ( 
.A(n_1287),
.Y(n_1466)
);

AOI22xp33_ASAP7_75t_L g1467 ( 
.A1(n_1343),
.A2(n_1068),
.B1(n_1345),
.B2(n_1320),
.Y(n_1467)
);

BUFx10_ASAP7_75t_L g1468 ( 
.A(n_1287),
.Y(n_1468)
);

NAND2xp5_ASAP7_75t_L g1469 ( 
.A(n_1275),
.B(n_1306),
.Y(n_1469)
);

BUFx6f_ASAP7_75t_L g1470 ( 
.A(n_1191),
.Y(n_1470)
);

CKINVDCx20_ASAP7_75t_R g1471 ( 
.A(n_1332),
.Y(n_1471)
);

BUFx3_ASAP7_75t_L g1472 ( 
.A(n_1291),
.Y(n_1472)
);

AOI22xp33_ASAP7_75t_SL g1473 ( 
.A1(n_1451),
.A2(n_1465),
.B1(n_1386),
.B2(n_1439),
.Y(n_1473)
);

AOI22xp33_ASAP7_75t_L g1474 ( 
.A1(n_1444),
.A2(n_1455),
.B1(n_1347),
.B2(n_1457),
.Y(n_1474)
);

INVx2_ASAP7_75t_L g1475 ( 
.A(n_1384),
.Y(n_1475)
);

BUFx2_ASAP7_75t_L g1476 ( 
.A(n_1438),
.Y(n_1476)
);

AO31x2_ASAP7_75t_L g1477 ( 
.A1(n_1434),
.A2(n_1422),
.A3(n_1372),
.B(n_1420),
.Y(n_1477)
);

INVx2_ASAP7_75t_L g1478 ( 
.A(n_1432),
.Y(n_1478)
);

HB1xp67_ASAP7_75t_L g1479 ( 
.A(n_1400),
.Y(n_1479)
);

INVx6_ASAP7_75t_L g1480 ( 
.A(n_1382),
.Y(n_1480)
);

OR2x2_ASAP7_75t_L g1481 ( 
.A(n_1362),
.B(n_1356),
.Y(n_1481)
);

NOR2xp33_ASAP7_75t_L g1482 ( 
.A(n_1445),
.B(n_1469),
.Y(n_1482)
);

INVx3_ASAP7_75t_L g1483 ( 
.A(n_1427),
.Y(n_1483)
);

HB1xp67_ASAP7_75t_L g1484 ( 
.A(n_1398),
.Y(n_1484)
);

INVx2_ASAP7_75t_L g1485 ( 
.A(n_1442),
.Y(n_1485)
);

BUFx2_ASAP7_75t_L g1486 ( 
.A(n_1436),
.Y(n_1486)
);

HB1xp67_ASAP7_75t_L g1487 ( 
.A(n_1375),
.Y(n_1487)
);

INVx2_ASAP7_75t_L g1488 ( 
.A(n_1440),
.Y(n_1488)
);

INVx1_ASAP7_75t_L g1489 ( 
.A(n_1441),
.Y(n_1489)
);

AND2x2_ASAP7_75t_SL g1490 ( 
.A(n_1366),
.B(n_1362),
.Y(n_1490)
);

INVx1_ASAP7_75t_L g1491 ( 
.A(n_1394),
.Y(n_1491)
);

OR2x6_ASAP7_75t_L g1492 ( 
.A(n_1436),
.B(n_1382),
.Y(n_1492)
);

AO21x2_ASAP7_75t_L g1493 ( 
.A1(n_1379),
.A2(n_1415),
.B(n_1380),
.Y(n_1493)
);

INVx1_ASAP7_75t_L g1494 ( 
.A(n_1394),
.Y(n_1494)
);

INVx1_ASAP7_75t_L g1495 ( 
.A(n_1368),
.Y(n_1495)
);

INVx3_ASAP7_75t_L g1496 ( 
.A(n_1425),
.Y(n_1496)
);

INVx1_ASAP7_75t_L g1497 ( 
.A(n_1351),
.Y(n_1497)
);

INVx1_ASAP7_75t_L g1498 ( 
.A(n_1351),
.Y(n_1498)
);

OAI22xp5_ASAP7_75t_L g1499 ( 
.A1(n_1349),
.A2(n_1369),
.B1(n_1350),
.B2(n_1366),
.Y(n_1499)
);

INVx2_ASAP7_75t_SL g1500 ( 
.A(n_1425),
.Y(n_1500)
);

AND2x2_ASAP7_75t_L g1501 ( 
.A(n_1359),
.B(n_1356),
.Y(n_1501)
);

AND2x2_ASAP7_75t_L g1502 ( 
.A(n_1359),
.B(n_1369),
.Y(n_1502)
);

INVx1_ASAP7_75t_L g1503 ( 
.A(n_1408),
.Y(n_1503)
);

AND2x2_ASAP7_75t_L g1504 ( 
.A(n_1350),
.B(n_1348),
.Y(n_1504)
);

INVx1_ASAP7_75t_L g1505 ( 
.A(n_1408),
.Y(n_1505)
);

AOI22xp33_ASAP7_75t_L g1506 ( 
.A1(n_1455),
.A2(n_1449),
.B1(n_1467),
.B2(n_1458),
.Y(n_1506)
);

AO21x1_ASAP7_75t_SL g1507 ( 
.A1(n_1348),
.A2(n_1449),
.B(n_1457),
.Y(n_1507)
);

OA21x2_ASAP7_75t_L g1508 ( 
.A1(n_1404),
.A2(n_1389),
.B(n_1416),
.Y(n_1508)
);

NOR2xp33_ASAP7_75t_L g1509 ( 
.A(n_1361),
.B(n_1373),
.Y(n_1509)
);

INVx2_ASAP7_75t_L g1510 ( 
.A(n_1435),
.Y(n_1510)
);

NAND2xp5_ASAP7_75t_L g1511 ( 
.A(n_1376),
.B(n_1352),
.Y(n_1511)
);

INVx1_ASAP7_75t_L g1512 ( 
.A(n_1430),
.Y(n_1512)
);

INVx2_ASAP7_75t_L g1513 ( 
.A(n_1437),
.Y(n_1513)
);

BUFx3_ASAP7_75t_L g1514 ( 
.A(n_1393),
.Y(n_1514)
);

INVx1_ASAP7_75t_L g1515 ( 
.A(n_1430),
.Y(n_1515)
);

INVx1_ASAP7_75t_L g1516 ( 
.A(n_1421),
.Y(n_1516)
);

INVx1_ASAP7_75t_L g1517 ( 
.A(n_1421),
.Y(n_1517)
);

INVx1_ASAP7_75t_L g1518 ( 
.A(n_1391),
.Y(n_1518)
);

INVx2_ASAP7_75t_L g1519 ( 
.A(n_1390),
.Y(n_1519)
);

INVx1_ASAP7_75t_L g1520 ( 
.A(n_1391),
.Y(n_1520)
);

INVx1_ASAP7_75t_SL g1521 ( 
.A(n_1460),
.Y(n_1521)
);

AOI21x1_ASAP7_75t_L g1522 ( 
.A1(n_1405),
.A2(n_1387),
.B(n_1374),
.Y(n_1522)
);

NAND2xp5_ASAP7_75t_L g1523 ( 
.A(n_1376),
.B(n_1352),
.Y(n_1523)
);

BUFx2_ASAP7_75t_L g1524 ( 
.A(n_1383),
.Y(n_1524)
);

AND2x2_ASAP7_75t_L g1525 ( 
.A(n_1349),
.B(n_1447),
.Y(n_1525)
);

AOI22xp33_ASAP7_75t_SL g1526 ( 
.A1(n_1367),
.A2(n_1418),
.B1(n_1460),
.B2(n_1409),
.Y(n_1526)
);

BUFx3_ASAP7_75t_L g1527 ( 
.A(n_1346),
.Y(n_1527)
);

HB1xp67_ASAP7_75t_L g1528 ( 
.A(n_1450),
.Y(n_1528)
);

NAND2xp5_ASAP7_75t_L g1529 ( 
.A(n_1379),
.B(n_1447),
.Y(n_1529)
);

BUFx3_ASAP7_75t_L g1530 ( 
.A(n_1346),
.Y(n_1530)
);

INVx1_ASAP7_75t_L g1531 ( 
.A(n_1454),
.Y(n_1531)
);

HB1xp67_ASAP7_75t_L g1532 ( 
.A(n_1459),
.Y(n_1532)
);

AND2x2_ASAP7_75t_L g1533 ( 
.A(n_1458),
.B(n_1467),
.Y(n_1533)
);

OA21x2_ASAP7_75t_L g1534 ( 
.A1(n_1404),
.A2(n_1389),
.B(n_1416),
.Y(n_1534)
);

INVx1_ASAP7_75t_L g1535 ( 
.A(n_1431),
.Y(n_1535)
);

NAND2xp5_ASAP7_75t_L g1536 ( 
.A(n_1385),
.B(n_1370),
.Y(n_1536)
);

BUFx3_ASAP7_75t_L g1537 ( 
.A(n_1355),
.Y(n_1537)
);

AND2x2_ASAP7_75t_L g1538 ( 
.A(n_1385),
.B(n_1364),
.Y(n_1538)
);

INVx2_ASAP7_75t_L g1539 ( 
.A(n_1424),
.Y(n_1539)
);

AND2x2_ASAP7_75t_L g1540 ( 
.A(n_1365),
.B(n_1426),
.Y(n_1540)
);

INVx1_ASAP7_75t_L g1541 ( 
.A(n_1428),
.Y(n_1541)
);

INVx2_ASAP7_75t_L g1542 ( 
.A(n_1412),
.Y(n_1542)
);

INVx1_ASAP7_75t_L g1543 ( 
.A(n_1428),
.Y(n_1543)
);

HB1xp67_ASAP7_75t_L g1544 ( 
.A(n_1363),
.Y(n_1544)
);

INVx1_ASAP7_75t_L g1545 ( 
.A(n_1426),
.Y(n_1545)
);

INVx1_ASAP7_75t_L g1546 ( 
.A(n_1429),
.Y(n_1546)
);

AND2x2_ASAP7_75t_L g1547 ( 
.A(n_1418),
.B(n_1414),
.Y(n_1547)
);

OAI22xp5_ASAP7_75t_L g1548 ( 
.A1(n_1402),
.A2(n_1397),
.B1(n_1463),
.B2(n_1355),
.Y(n_1548)
);

INVx1_ASAP7_75t_L g1549 ( 
.A(n_1433),
.Y(n_1549)
);

OA21x2_ASAP7_75t_L g1550 ( 
.A1(n_1433),
.A2(n_1423),
.B(n_1410),
.Y(n_1550)
);

OAI21x1_ASAP7_75t_L g1551 ( 
.A1(n_1355),
.A2(n_1456),
.B(n_1443),
.Y(n_1551)
);

OAI21x1_ASAP7_75t_L g1552 ( 
.A1(n_1443),
.A2(n_1456),
.B(n_1463),
.Y(n_1552)
);

NOR2x1_ASAP7_75t_R g1553 ( 
.A(n_1480),
.B(n_1446),
.Y(n_1553)
);

A2O1A1Ixp33_ASAP7_75t_L g1554 ( 
.A1(n_1473),
.A2(n_1464),
.B(n_1470),
.C(n_1419),
.Y(n_1554)
);

INVx1_ASAP7_75t_L g1555 ( 
.A(n_1495),
.Y(n_1555)
);

AND2x2_ASAP7_75t_L g1556 ( 
.A(n_1547),
.B(n_1462),
.Y(n_1556)
);

NAND2xp33_ASAP7_75t_L g1557 ( 
.A(n_1474),
.B(n_1464),
.Y(n_1557)
);

NOR2x1_ASAP7_75t_SL g1558 ( 
.A(n_1492),
.B(n_1522),
.Y(n_1558)
);

OR2x2_ASAP7_75t_L g1559 ( 
.A(n_1497),
.B(n_1472),
.Y(n_1559)
);

AND2x2_ASAP7_75t_L g1560 ( 
.A(n_1547),
.B(n_1510),
.Y(n_1560)
);

OAI21xp5_ASAP7_75t_L g1561 ( 
.A1(n_1506),
.A2(n_1473),
.B(n_1499),
.Y(n_1561)
);

HB1xp67_ASAP7_75t_L g1562 ( 
.A(n_1497),
.Y(n_1562)
);

AND2x2_ASAP7_75t_L g1563 ( 
.A(n_1510),
.B(n_1406),
.Y(n_1563)
);

A2O1A1Ixp33_ASAP7_75t_L g1564 ( 
.A1(n_1499),
.A2(n_1470),
.B(n_1401),
.C(n_1452),
.Y(n_1564)
);

NOR2xp33_ASAP7_75t_L g1565 ( 
.A(n_1486),
.B(n_1479),
.Y(n_1565)
);

OR2x2_ASAP7_75t_L g1566 ( 
.A(n_1498),
.B(n_1354),
.Y(n_1566)
);

AND2x2_ASAP7_75t_L g1567 ( 
.A(n_1510),
.B(n_1406),
.Y(n_1567)
);

OR2x2_ASAP7_75t_L g1568 ( 
.A(n_1498),
.B(n_1542),
.Y(n_1568)
);

AOI22xp5_ASAP7_75t_L g1569 ( 
.A1(n_1490),
.A2(n_1381),
.B1(n_1360),
.B2(n_1388),
.Y(n_1569)
);

OAI21xp33_ASAP7_75t_L g1570 ( 
.A1(n_1529),
.A2(n_1392),
.B(n_1358),
.Y(n_1570)
);

OAI22xp5_ASAP7_75t_L g1571 ( 
.A1(n_1526),
.A2(n_1377),
.B1(n_1411),
.B2(n_1407),
.Y(n_1571)
);

NOR2xp33_ASAP7_75t_L g1572 ( 
.A(n_1486),
.B(n_1411),
.Y(n_1572)
);

AO32x1_ASAP7_75t_L g1573 ( 
.A1(n_1504),
.A2(n_1463),
.A3(n_1443),
.B1(n_1456),
.B2(n_1413),
.Y(n_1573)
);

NAND2xp5_ASAP7_75t_L g1574 ( 
.A(n_1482),
.B(n_1417),
.Y(n_1574)
);

AOI221xp5_ASAP7_75t_L g1575 ( 
.A1(n_1529),
.A2(n_1533),
.B1(n_1504),
.B2(n_1525),
.C(n_1501),
.Y(n_1575)
);

OAI21xp5_ASAP7_75t_L g1576 ( 
.A1(n_1533),
.A2(n_1466),
.B(n_1395),
.Y(n_1576)
);

AND2x2_ASAP7_75t_L g1577 ( 
.A(n_1513),
.B(n_1487),
.Y(n_1577)
);

AND2x4_ASAP7_75t_L g1578 ( 
.A(n_1489),
.B(n_1378),
.Y(n_1578)
);

AND2x4_ASAP7_75t_SL g1579 ( 
.A(n_1492),
.B(n_1468),
.Y(n_1579)
);

AO32x2_ASAP7_75t_L g1580 ( 
.A1(n_1500),
.A2(n_1378),
.A3(n_1396),
.B1(n_1403),
.B2(n_1407),
.Y(n_1580)
);

AND2x2_ASAP7_75t_L g1581 ( 
.A(n_1513),
.B(n_1461),
.Y(n_1581)
);

AND2x2_ASAP7_75t_L g1582 ( 
.A(n_1513),
.B(n_1461),
.Y(n_1582)
);

OAI21x1_ASAP7_75t_SL g1583 ( 
.A1(n_1522),
.A2(n_1448),
.B(n_1453),
.Y(n_1583)
);

AOI22xp5_ASAP7_75t_L g1584 ( 
.A1(n_1490),
.A2(n_1353),
.B1(n_1399),
.B2(n_1471),
.Y(n_1584)
);

A2O1A1Ixp33_ASAP7_75t_SL g1585 ( 
.A1(n_1483),
.A2(n_1407),
.B(n_1411),
.C(n_1470),
.Y(n_1585)
);

AND2x2_ASAP7_75t_L g1586 ( 
.A(n_1540),
.B(n_1468),
.Y(n_1586)
);

AND2x2_ASAP7_75t_L g1587 ( 
.A(n_1540),
.B(n_1509),
.Y(n_1587)
);

AO22x2_ASAP7_75t_L g1588 ( 
.A1(n_1516),
.A2(n_1357),
.B1(n_1371),
.B2(n_1517),
.Y(n_1588)
);

NAND2xp5_ASAP7_75t_L g1589 ( 
.A(n_1542),
.B(n_1525),
.Y(n_1589)
);

AOI22xp5_ASAP7_75t_L g1590 ( 
.A1(n_1490),
.A2(n_1502),
.B1(n_1501),
.B2(n_1526),
.Y(n_1590)
);

AOI21xp5_ASAP7_75t_SL g1591 ( 
.A1(n_1508),
.A2(n_1534),
.B(n_1492),
.Y(n_1591)
);

OAI22xp5_ASAP7_75t_SL g1592 ( 
.A1(n_1521),
.A2(n_1476),
.B1(n_1481),
.B2(n_1500),
.Y(n_1592)
);

OR2x6_ASAP7_75t_L g1593 ( 
.A(n_1492),
.B(n_1551),
.Y(n_1593)
);

OA21x2_ASAP7_75t_L g1594 ( 
.A1(n_1545),
.A2(n_1516),
.B(n_1517),
.Y(n_1594)
);

INVx2_ASAP7_75t_L g1595 ( 
.A(n_1519),
.Y(n_1595)
);

AND2x2_ASAP7_75t_L g1596 ( 
.A(n_1528),
.B(n_1532),
.Y(n_1596)
);

BUFx12f_ASAP7_75t_L g1597 ( 
.A(n_1500),
.Y(n_1597)
);

NAND2xp5_ASAP7_75t_L g1598 ( 
.A(n_1484),
.B(n_1502),
.Y(n_1598)
);

AND2x2_ASAP7_75t_L g1599 ( 
.A(n_1538),
.B(n_1524),
.Y(n_1599)
);

OR2x6_ASAP7_75t_L g1600 ( 
.A(n_1551),
.B(n_1552),
.Y(n_1600)
);

AND2x4_ASAP7_75t_L g1601 ( 
.A(n_1485),
.B(n_1551),
.Y(n_1601)
);

OAI21xp5_ASAP7_75t_L g1602 ( 
.A1(n_1511),
.A2(n_1523),
.B(n_1481),
.Y(n_1602)
);

AO21x1_ASAP7_75t_L g1603 ( 
.A1(n_1535),
.A2(n_1523),
.B(n_1511),
.Y(n_1603)
);

OR2x6_ASAP7_75t_L g1604 ( 
.A(n_1552),
.B(n_1548),
.Y(n_1604)
);

AND2x2_ASAP7_75t_L g1605 ( 
.A(n_1539),
.B(n_1544),
.Y(n_1605)
);

OR2x2_ASAP7_75t_L g1606 ( 
.A(n_1478),
.B(n_1477),
.Y(n_1606)
);

AND2x4_ASAP7_75t_L g1607 ( 
.A(n_1485),
.B(n_1552),
.Y(n_1607)
);

OAI22xp5_ASAP7_75t_L g1608 ( 
.A1(n_1548),
.A2(n_1536),
.B1(n_1518),
.B2(n_1520),
.Y(n_1608)
);

NOR2xp33_ASAP7_75t_L g1609 ( 
.A(n_1536),
.B(n_1496),
.Y(n_1609)
);

NOR2xp33_ASAP7_75t_L g1610 ( 
.A(n_1496),
.B(n_1518),
.Y(n_1610)
);

INVxp67_ASAP7_75t_L g1611 ( 
.A(n_1493),
.Y(n_1611)
);

AND2x2_ASAP7_75t_L g1612 ( 
.A(n_1601),
.B(n_1607),
.Y(n_1612)
);

NAND2xp5_ASAP7_75t_L g1613 ( 
.A(n_1589),
.B(n_1477),
.Y(n_1613)
);

OR2x2_ASAP7_75t_L g1614 ( 
.A(n_1606),
.B(n_1550),
.Y(n_1614)
);

AOI22xp33_ASAP7_75t_L g1615 ( 
.A1(n_1561),
.A2(n_1507),
.B1(n_1534),
.B2(n_1508),
.Y(n_1615)
);

INVx2_ASAP7_75t_L g1616 ( 
.A(n_1595),
.Y(n_1616)
);

AND2x2_ASAP7_75t_L g1617 ( 
.A(n_1601),
.B(n_1550),
.Y(n_1617)
);

AND2x4_ASAP7_75t_L g1618 ( 
.A(n_1600),
.B(n_1475),
.Y(n_1618)
);

HB1xp67_ASAP7_75t_L g1619 ( 
.A(n_1562),
.Y(n_1619)
);

NAND2xp5_ASAP7_75t_L g1620 ( 
.A(n_1594),
.B(n_1477),
.Y(n_1620)
);

NAND2xp5_ASAP7_75t_L g1621 ( 
.A(n_1594),
.B(n_1477),
.Y(n_1621)
);

INVx1_ASAP7_75t_L g1622 ( 
.A(n_1595),
.Y(n_1622)
);

AND2x2_ASAP7_75t_L g1623 ( 
.A(n_1601),
.B(n_1550),
.Y(n_1623)
);

AND2x2_ASAP7_75t_L g1624 ( 
.A(n_1607),
.B(n_1550),
.Y(n_1624)
);

NOR2x1p5_ASAP7_75t_L g1625 ( 
.A(n_1597),
.B(n_1514),
.Y(n_1625)
);

AND2x2_ASAP7_75t_L g1626 ( 
.A(n_1607),
.B(n_1545),
.Y(n_1626)
);

AND2x2_ASAP7_75t_L g1627 ( 
.A(n_1591),
.B(n_1491),
.Y(n_1627)
);

INVx2_ASAP7_75t_L g1628 ( 
.A(n_1555),
.Y(n_1628)
);

AND2x2_ASAP7_75t_L g1629 ( 
.A(n_1591),
.B(n_1494),
.Y(n_1629)
);

INVx5_ASAP7_75t_L g1630 ( 
.A(n_1593),
.Y(n_1630)
);

AND2x2_ASAP7_75t_L g1631 ( 
.A(n_1594),
.B(n_1494),
.Y(n_1631)
);

OR2x2_ASAP7_75t_L g1632 ( 
.A(n_1611),
.B(n_1541),
.Y(n_1632)
);

AND2x2_ASAP7_75t_L g1633 ( 
.A(n_1593),
.B(n_1541),
.Y(n_1633)
);

AOI22xp33_ASAP7_75t_L g1634 ( 
.A1(n_1557),
.A2(n_1507),
.B1(n_1508),
.B2(n_1534),
.Y(n_1634)
);

INVx3_ASAP7_75t_L g1635 ( 
.A(n_1593),
.Y(n_1635)
);

OAI221xp5_ASAP7_75t_L g1636 ( 
.A1(n_1557),
.A2(n_1520),
.B1(n_1503),
.B2(n_1505),
.C(n_1534),
.Y(n_1636)
);

AND2x2_ASAP7_75t_L g1637 ( 
.A(n_1611),
.B(n_1543),
.Y(n_1637)
);

INVxp67_ASAP7_75t_L g1638 ( 
.A(n_1562),
.Y(n_1638)
);

OR2x2_ASAP7_75t_L g1639 ( 
.A(n_1568),
.B(n_1549),
.Y(n_1639)
);

BUFx3_ASAP7_75t_L g1640 ( 
.A(n_1583),
.Y(n_1640)
);

BUFx3_ASAP7_75t_L g1641 ( 
.A(n_1597),
.Y(n_1641)
);

OR2x2_ASAP7_75t_L g1642 ( 
.A(n_1596),
.B(n_1488),
.Y(n_1642)
);

NAND2xp5_ASAP7_75t_L g1643 ( 
.A(n_1609),
.B(n_1477),
.Y(n_1643)
);

AOI22xp33_ASAP7_75t_L g1644 ( 
.A1(n_1575),
.A2(n_1508),
.B1(n_1503),
.B2(n_1505),
.Y(n_1644)
);

INVx1_ASAP7_75t_L g1645 ( 
.A(n_1573),
.Y(n_1645)
);

INVx1_ASAP7_75t_L g1646 ( 
.A(n_1628),
.Y(n_1646)
);

INVx1_ASAP7_75t_L g1647 ( 
.A(n_1628),
.Y(n_1647)
);

INVx2_ASAP7_75t_L g1648 ( 
.A(n_1616),
.Y(n_1648)
);

OR2x2_ASAP7_75t_L g1649 ( 
.A(n_1643),
.B(n_1598),
.Y(n_1649)
);

OAI321xp33_ASAP7_75t_L g1650 ( 
.A1(n_1636),
.A2(n_1615),
.A3(n_1590),
.B1(n_1644),
.B2(n_1554),
.C(n_1634),
.Y(n_1650)
);

NOR3xp33_ASAP7_75t_L g1651 ( 
.A(n_1636),
.B(n_1571),
.C(n_1570),
.Y(n_1651)
);

NAND2xp5_ASAP7_75t_L g1652 ( 
.A(n_1613),
.B(n_1609),
.Y(n_1652)
);

AOI33xp33_ASAP7_75t_L g1653 ( 
.A1(n_1615),
.A2(n_1587),
.A3(n_1586),
.B1(n_1584),
.B2(n_1577),
.B3(n_1569),
.Y(n_1653)
);

AOI211xp5_ASAP7_75t_SL g1654 ( 
.A1(n_1643),
.A2(n_1554),
.B(n_1564),
.C(n_1592),
.Y(n_1654)
);

AND2x2_ASAP7_75t_L g1655 ( 
.A(n_1612),
.B(n_1599),
.Y(n_1655)
);

INVx1_ASAP7_75t_L g1656 ( 
.A(n_1628),
.Y(n_1656)
);

AND3x2_ASAP7_75t_L g1657 ( 
.A(n_1638),
.B(n_1582),
.C(n_1581),
.Y(n_1657)
);

AOI22xp5_ASAP7_75t_L g1658 ( 
.A1(n_1644),
.A2(n_1602),
.B1(n_1588),
.B2(n_1608),
.Y(n_1658)
);

AND2x2_ASAP7_75t_L g1659 ( 
.A(n_1612),
.B(n_1604),
.Y(n_1659)
);

NAND2xp5_ASAP7_75t_L g1660 ( 
.A(n_1613),
.B(n_1603),
.Y(n_1660)
);

AND2x4_ASAP7_75t_L g1661 ( 
.A(n_1635),
.B(n_1604),
.Y(n_1661)
);

HB1xp67_ASAP7_75t_L g1662 ( 
.A(n_1619),
.Y(n_1662)
);

INVx4_ASAP7_75t_L g1663 ( 
.A(n_1641),
.Y(n_1663)
);

AOI22xp5_ASAP7_75t_L g1664 ( 
.A1(n_1634),
.A2(n_1588),
.B1(n_1564),
.B2(n_1565),
.Y(n_1664)
);

NAND4xp25_ASAP7_75t_L g1665 ( 
.A(n_1620),
.B(n_1565),
.C(n_1576),
.D(n_1574),
.Y(n_1665)
);

INVx1_ASAP7_75t_SL g1666 ( 
.A(n_1639),
.Y(n_1666)
);

AND2x2_ASAP7_75t_L g1667 ( 
.A(n_1612),
.B(n_1604),
.Y(n_1667)
);

OR2x2_ASAP7_75t_L g1668 ( 
.A(n_1642),
.B(n_1546),
.Y(n_1668)
);

OAI21xp5_ASAP7_75t_L g1669 ( 
.A1(n_1620),
.A2(n_1572),
.B(n_1610),
.Y(n_1669)
);

INVx1_ASAP7_75t_L g1670 ( 
.A(n_1619),
.Y(n_1670)
);

NAND2xp5_ASAP7_75t_L g1671 ( 
.A(n_1637),
.B(n_1477),
.Y(n_1671)
);

NAND2xp5_ASAP7_75t_L g1672 ( 
.A(n_1637),
.B(n_1605),
.Y(n_1672)
);

OAI33xp33_ASAP7_75t_L g1673 ( 
.A1(n_1632),
.A2(n_1515),
.A3(n_1512),
.B1(n_1559),
.B2(n_1566),
.B3(n_1531),
.Y(n_1673)
);

INVx3_ASAP7_75t_L g1674 ( 
.A(n_1618),
.Y(n_1674)
);

AND2x2_ASAP7_75t_L g1675 ( 
.A(n_1626),
.B(n_1560),
.Y(n_1675)
);

INVx1_ASAP7_75t_L g1676 ( 
.A(n_1622),
.Y(n_1676)
);

AND2x4_ASAP7_75t_L g1677 ( 
.A(n_1635),
.B(n_1558),
.Y(n_1677)
);

AOI222xp33_ASAP7_75t_L g1678 ( 
.A1(n_1645),
.A2(n_1553),
.B1(n_1512),
.B2(n_1515),
.C1(n_1588),
.C2(n_1579),
.Y(n_1678)
);

INVx2_ASAP7_75t_L g1679 ( 
.A(n_1631),
.Y(n_1679)
);

INVx1_ASAP7_75t_L g1680 ( 
.A(n_1622),
.Y(n_1680)
);

NAND2xp5_ASAP7_75t_L g1681 ( 
.A(n_1637),
.B(n_1493),
.Y(n_1681)
);

HB1xp67_ASAP7_75t_L g1682 ( 
.A(n_1626),
.Y(n_1682)
);

INVx2_ASAP7_75t_L g1683 ( 
.A(n_1679),
.Y(n_1683)
);

AND2x4_ASAP7_75t_L g1684 ( 
.A(n_1661),
.B(n_1630),
.Y(n_1684)
);

AND2x2_ASAP7_75t_L g1685 ( 
.A(n_1674),
.B(n_1617),
.Y(n_1685)
);

AOI221xp5_ASAP7_75t_L g1686 ( 
.A1(n_1650),
.A2(n_1621),
.B1(n_1645),
.B2(n_1627),
.C(n_1629),
.Y(n_1686)
);

OR2x2_ASAP7_75t_SL g1687 ( 
.A(n_1660),
.B(n_1645),
.Y(n_1687)
);

AND2x2_ASAP7_75t_L g1688 ( 
.A(n_1674),
.B(n_1617),
.Y(n_1688)
);

INVx1_ASAP7_75t_L g1689 ( 
.A(n_1676),
.Y(n_1689)
);

INVx2_ASAP7_75t_L g1690 ( 
.A(n_1679),
.Y(n_1690)
);

OR2x2_ASAP7_75t_L g1691 ( 
.A(n_1681),
.B(n_1621),
.Y(n_1691)
);

HB1xp67_ASAP7_75t_L g1692 ( 
.A(n_1662),
.Y(n_1692)
);

NOR3xp33_ASAP7_75t_SL g1693 ( 
.A(n_1650),
.B(n_1572),
.C(n_1610),
.Y(n_1693)
);

AND2x2_ASAP7_75t_L g1694 ( 
.A(n_1674),
.B(n_1617),
.Y(n_1694)
);

OR2x2_ASAP7_75t_L g1695 ( 
.A(n_1681),
.B(n_1614),
.Y(n_1695)
);

HB1xp67_ASAP7_75t_L g1696 ( 
.A(n_1676),
.Y(n_1696)
);

NAND2xp5_ASAP7_75t_L g1697 ( 
.A(n_1660),
.B(n_1631),
.Y(n_1697)
);

NOR2xp33_ASAP7_75t_L g1698 ( 
.A(n_1665),
.B(n_1556),
.Y(n_1698)
);

NOR2x1_ASAP7_75t_L g1699 ( 
.A(n_1663),
.B(n_1640),
.Y(n_1699)
);

INVx1_ASAP7_75t_L g1700 ( 
.A(n_1680),
.Y(n_1700)
);

INVx1_ASAP7_75t_L g1701 ( 
.A(n_1680),
.Y(n_1701)
);

AND2x2_ASAP7_75t_L g1702 ( 
.A(n_1674),
.B(n_1623),
.Y(n_1702)
);

INVx2_ASAP7_75t_L g1703 ( 
.A(n_1679),
.Y(n_1703)
);

INVx2_ASAP7_75t_L g1704 ( 
.A(n_1648),
.Y(n_1704)
);

AOI22xp33_ASAP7_75t_L g1705 ( 
.A1(n_1651),
.A2(n_1493),
.B1(n_1640),
.B2(n_1633),
.Y(n_1705)
);

INVx1_ASAP7_75t_L g1706 ( 
.A(n_1670),
.Y(n_1706)
);

BUFx3_ASAP7_75t_L g1707 ( 
.A(n_1663),
.Y(n_1707)
);

NOR2xp33_ASAP7_75t_L g1708 ( 
.A(n_1665),
.B(n_1640),
.Y(n_1708)
);

INVx1_ASAP7_75t_L g1709 ( 
.A(n_1670),
.Y(n_1709)
);

AND2x4_ASAP7_75t_SL g1710 ( 
.A(n_1663),
.B(n_1635),
.Y(n_1710)
);

NOR2xp33_ASAP7_75t_L g1711 ( 
.A(n_1663),
.B(n_1640),
.Y(n_1711)
);

INVx1_ASAP7_75t_L g1712 ( 
.A(n_1646),
.Y(n_1712)
);

HB1xp67_ASAP7_75t_L g1713 ( 
.A(n_1646),
.Y(n_1713)
);

AND2x2_ASAP7_75t_L g1714 ( 
.A(n_1682),
.B(n_1623),
.Y(n_1714)
);

INVx2_ASAP7_75t_L g1715 ( 
.A(n_1648),
.Y(n_1715)
);

NAND2xp5_ASAP7_75t_SL g1716 ( 
.A(n_1658),
.B(n_1630),
.Y(n_1716)
);

AND2x2_ASAP7_75t_L g1717 ( 
.A(n_1666),
.B(n_1623),
.Y(n_1717)
);

INVx2_ASAP7_75t_L g1718 ( 
.A(n_1648),
.Y(n_1718)
);

INVx1_ASAP7_75t_L g1719 ( 
.A(n_1647),
.Y(n_1719)
);

BUFx2_ASAP7_75t_L g1720 ( 
.A(n_1677),
.Y(n_1720)
);

AND2x2_ASAP7_75t_L g1721 ( 
.A(n_1666),
.B(n_1624),
.Y(n_1721)
);

OR2x2_ASAP7_75t_L g1722 ( 
.A(n_1671),
.B(n_1668),
.Y(n_1722)
);

INVx1_ASAP7_75t_L g1723 ( 
.A(n_1696),
.Y(n_1723)
);

INVx1_ASAP7_75t_L g1724 ( 
.A(n_1696),
.Y(n_1724)
);

OR2x2_ASAP7_75t_L g1725 ( 
.A(n_1722),
.B(n_1649),
.Y(n_1725)
);

INVx1_ASAP7_75t_L g1726 ( 
.A(n_1706),
.Y(n_1726)
);

NAND2xp5_ASAP7_75t_L g1727 ( 
.A(n_1697),
.B(n_1652),
.Y(n_1727)
);

AOI22xp5_ASAP7_75t_L g1728 ( 
.A1(n_1686),
.A2(n_1658),
.B1(n_1664),
.B2(n_1678),
.Y(n_1728)
);

OR2x2_ASAP7_75t_L g1729 ( 
.A(n_1722),
.B(n_1649),
.Y(n_1729)
);

HB1xp67_ASAP7_75t_L g1730 ( 
.A(n_1692),
.Y(n_1730)
);

OR2x2_ASAP7_75t_L g1731 ( 
.A(n_1722),
.B(n_1671),
.Y(n_1731)
);

OR2x2_ASAP7_75t_L g1732 ( 
.A(n_1697),
.B(n_1652),
.Y(n_1732)
);

INVx1_ASAP7_75t_L g1733 ( 
.A(n_1706),
.Y(n_1733)
);

NAND3xp33_ASAP7_75t_L g1734 ( 
.A(n_1693),
.B(n_1654),
.C(n_1664),
.Y(n_1734)
);

NAND2xp5_ASAP7_75t_L g1735 ( 
.A(n_1709),
.B(n_1668),
.Y(n_1735)
);

OR2x2_ASAP7_75t_L g1736 ( 
.A(n_1687),
.B(n_1672),
.Y(n_1736)
);

NOR2x1_ASAP7_75t_L g1737 ( 
.A(n_1699),
.B(n_1641),
.Y(n_1737)
);

INVx1_ASAP7_75t_L g1738 ( 
.A(n_1709),
.Y(n_1738)
);

NAND2xp5_ASAP7_75t_L g1739 ( 
.A(n_1686),
.B(n_1631),
.Y(n_1739)
);

OR2x2_ASAP7_75t_L g1740 ( 
.A(n_1687),
.B(n_1672),
.Y(n_1740)
);

OR2x2_ASAP7_75t_L g1741 ( 
.A(n_1687),
.B(n_1669),
.Y(n_1741)
);

OR2x2_ASAP7_75t_L g1742 ( 
.A(n_1695),
.B(n_1669),
.Y(n_1742)
);

INVxp67_ASAP7_75t_L g1743 ( 
.A(n_1708),
.Y(n_1743)
);

OR2x2_ASAP7_75t_L g1744 ( 
.A(n_1695),
.B(n_1642),
.Y(n_1744)
);

INVx1_ASAP7_75t_L g1745 ( 
.A(n_1689),
.Y(n_1745)
);

INVx1_ASAP7_75t_L g1746 ( 
.A(n_1689),
.Y(n_1746)
);

NAND2xp5_ASAP7_75t_L g1747 ( 
.A(n_1692),
.B(n_1647),
.Y(n_1747)
);

INVx1_ASAP7_75t_L g1748 ( 
.A(n_1700),
.Y(n_1748)
);

NAND2xp5_ASAP7_75t_R g1749 ( 
.A(n_1708),
.B(n_1661),
.Y(n_1749)
);

AND2x2_ASAP7_75t_L g1750 ( 
.A(n_1711),
.B(n_1659),
.Y(n_1750)
);

AND2x2_ASAP7_75t_L g1751 ( 
.A(n_1711),
.B(n_1659),
.Y(n_1751)
);

OR2x2_ASAP7_75t_L g1752 ( 
.A(n_1695),
.B(n_1642),
.Y(n_1752)
);

INVx1_ASAP7_75t_L g1753 ( 
.A(n_1700),
.Y(n_1753)
);

INVx1_ASAP7_75t_L g1754 ( 
.A(n_1701),
.Y(n_1754)
);

INVx1_ASAP7_75t_L g1755 ( 
.A(n_1701),
.Y(n_1755)
);

AND2x2_ASAP7_75t_L g1756 ( 
.A(n_1684),
.B(n_1667),
.Y(n_1756)
);

AND2x4_ASAP7_75t_L g1757 ( 
.A(n_1699),
.B(n_1707),
.Y(n_1757)
);

NAND2xp5_ASAP7_75t_L g1758 ( 
.A(n_1698),
.B(n_1656),
.Y(n_1758)
);

INVx1_ASAP7_75t_L g1759 ( 
.A(n_1713),
.Y(n_1759)
);

NAND2xp5_ASAP7_75t_L g1760 ( 
.A(n_1698),
.B(n_1656),
.Y(n_1760)
);

INVx2_ASAP7_75t_SL g1761 ( 
.A(n_1707),
.Y(n_1761)
);

AND2x2_ASAP7_75t_L g1762 ( 
.A(n_1684),
.B(n_1667),
.Y(n_1762)
);

INVx1_ASAP7_75t_L g1763 ( 
.A(n_1713),
.Y(n_1763)
);

BUFx2_ASAP7_75t_L g1764 ( 
.A(n_1707),
.Y(n_1764)
);

INVx2_ASAP7_75t_SL g1765 ( 
.A(n_1707),
.Y(n_1765)
);

NAND4xp25_ASAP7_75t_L g1766 ( 
.A(n_1734),
.B(n_1705),
.C(n_1654),
.D(n_1716),
.Y(n_1766)
);

OR2x2_ASAP7_75t_L g1767 ( 
.A(n_1736),
.B(n_1716),
.Y(n_1767)
);

INVx1_ASAP7_75t_L g1768 ( 
.A(n_1730),
.Y(n_1768)
);

INVx1_ASAP7_75t_L g1769 ( 
.A(n_1730),
.Y(n_1769)
);

INVx1_ASAP7_75t_L g1770 ( 
.A(n_1726),
.Y(n_1770)
);

INVx1_ASAP7_75t_L g1771 ( 
.A(n_1733),
.Y(n_1771)
);

INVx1_ASAP7_75t_SL g1772 ( 
.A(n_1764),
.Y(n_1772)
);

NOR2xp33_ASAP7_75t_L g1773 ( 
.A(n_1743),
.B(n_1673),
.Y(n_1773)
);

INVx1_ASAP7_75t_L g1774 ( 
.A(n_1738),
.Y(n_1774)
);

NAND4xp25_ASAP7_75t_L g1775 ( 
.A(n_1728),
.B(n_1743),
.C(n_1741),
.D(n_1705),
.Y(n_1775)
);

NAND2xp5_ASAP7_75t_SL g1776 ( 
.A(n_1737),
.B(n_1693),
.Y(n_1776)
);

INVx1_ASAP7_75t_L g1777 ( 
.A(n_1745),
.Y(n_1777)
);

NOR2xp33_ASAP7_75t_L g1778 ( 
.A(n_1739),
.B(n_1657),
.Y(n_1778)
);

INVx1_ASAP7_75t_L g1779 ( 
.A(n_1746),
.Y(n_1779)
);

NAND2xp5_ASAP7_75t_L g1780 ( 
.A(n_1740),
.B(n_1653),
.Y(n_1780)
);

INVx1_ASAP7_75t_L g1781 ( 
.A(n_1748),
.Y(n_1781)
);

NAND2xp5_ASAP7_75t_L g1782 ( 
.A(n_1758),
.B(n_1675),
.Y(n_1782)
);

INVx2_ASAP7_75t_SL g1783 ( 
.A(n_1757),
.Y(n_1783)
);

AND2x4_ASAP7_75t_L g1784 ( 
.A(n_1757),
.B(n_1710),
.Y(n_1784)
);

OR2x2_ASAP7_75t_L g1785 ( 
.A(n_1742),
.B(n_1691),
.Y(n_1785)
);

AND2x2_ASAP7_75t_L g1786 ( 
.A(n_1750),
.B(n_1684),
.Y(n_1786)
);

OR2x2_ASAP7_75t_L g1787 ( 
.A(n_1758),
.B(n_1691),
.Y(n_1787)
);

INVx1_ASAP7_75t_L g1788 ( 
.A(n_1753),
.Y(n_1788)
);

AND2x2_ASAP7_75t_L g1789 ( 
.A(n_1751),
.B(n_1684),
.Y(n_1789)
);

NAND2xp5_ASAP7_75t_L g1790 ( 
.A(n_1760),
.B(n_1675),
.Y(n_1790)
);

AND2x4_ASAP7_75t_L g1791 ( 
.A(n_1757),
.B(n_1710),
.Y(n_1791)
);

INVx2_ASAP7_75t_L g1792 ( 
.A(n_1754),
.Y(n_1792)
);

OR2x2_ASAP7_75t_L g1793 ( 
.A(n_1760),
.B(n_1691),
.Y(n_1793)
);

NAND2xp5_ASAP7_75t_L g1794 ( 
.A(n_1727),
.B(n_1678),
.Y(n_1794)
);

INVx1_ASAP7_75t_L g1795 ( 
.A(n_1755),
.Y(n_1795)
);

INVx1_ASAP7_75t_L g1796 ( 
.A(n_1723),
.Y(n_1796)
);

INVx1_ASAP7_75t_L g1797 ( 
.A(n_1724),
.Y(n_1797)
);

AND2x2_ASAP7_75t_L g1798 ( 
.A(n_1756),
.B(n_1684),
.Y(n_1798)
);

NAND2xp5_ASAP7_75t_L g1799 ( 
.A(n_1727),
.B(n_1655),
.Y(n_1799)
);

OR2x2_ASAP7_75t_L g1800 ( 
.A(n_1732),
.B(n_1725),
.Y(n_1800)
);

INVxp67_ASAP7_75t_L g1801 ( 
.A(n_1761),
.Y(n_1801)
);

OAI21xp33_ASAP7_75t_L g1802 ( 
.A1(n_1766),
.A2(n_1739),
.B(n_1749),
.Y(n_1802)
);

INVx1_ASAP7_75t_L g1803 ( 
.A(n_1792),
.Y(n_1803)
);

INVx1_ASAP7_75t_L g1804 ( 
.A(n_1792),
.Y(n_1804)
);

INVx1_ASAP7_75t_L g1805 ( 
.A(n_1768),
.Y(n_1805)
);

INVxp67_ASAP7_75t_L g1806 ( 
.A(n_1769),
.Y(n_1806)
);

NAND2xp5_ASAP7_75t_L g1807 ( 
.A(n_1772),
.B(n_1765),
.Y(n_1807)
);

NOR2xp33_ASAP7_75t_L g1808 ( 
.A(n_1775),
.B(n_1762),
.Y(n_1808)
);

INVxp67_ASAP7_75t_SL g1809 ( 
.A(n_1776),
.Y(n_1809)
);

AOI221xp5_ASAP7_75t_L g1810 ( 
.A1(n_1773),
.A2(n_1763),
.B1(n_1759),
.B2(n_1735),
.C(n_1720),
.Y(n_1810)
);

NAND2xp5_ASAP7_75t_L g1811 ( 
.A(n_1773),
.B(n_1780),
.Y(n_1811)
);

BUFx2_ASAP7_75t_L g1812 ( 
.A(n_1784),
.Y(n_1812)
);

OAI322xp33_ASAP7_75t_L g1813 ( 
.A1(n_1794),
.A2(n_1729),
.A3(n_1731),
.B1(n_1747),
.B2(n_1735),
.C1(n_1744),
.C2(n_1752),
.Y(n_1813)
);

NAND2xp5_ASAP7_75t_L g1814 ( 
.A(n_1801),
.B(n_1714),
.Y(n_1814)
);

O2A1O1Ixp33_ASAP7_75t_L g1815 ( 
.A1(n_1776),
.A2(n_1747),
.B(n_1720),
.C(n_1585),
.Y(n_1815)
);

INVx1_ASAP7_75t_L g1816 ( 
.A(n_1770),
.Y(n_1816)
);

INVx1_ASAP7_75t_L g1817 ( 
.A(n_1771),
.Y(n_1817)
);

INVx1_ASAP7_75t_SL g1818 ( 
.A(n_1784),
.Y(n_1818)
);

INVx3_ASAP7_75t_L g1819 ( 
.A(n_1784),
.Y(n_1819)
);

INVx1_ASAP7_75t_L g1820 ( 
.A(n_1774),
.Y(n_1820)
);

INVx1_ASAP7_75t_L g1821 ( 
.A(n_1777),
.Y(n_1821)
);

OAI22xp5_ASAP7_75t_L g1822 ( 
.A1(n_1778),
.A2(n_1720),
.B1(n_1630),
.B2(n_1661),
.Y(n_1822)
);

INVx2_ASAP7_75t_L g1823 ( 
.A(n_1783),
.Y(n_1823)
);

OAI221xp5_ASAP7_75t_L g1824 ( 
.A1(n_1778),
.A2(n_1641),
.B1(n_1635),
.B2(n_1630),
.C(n_1683),
.Y(n_1824)
);

AOI22xp5_ASAP7_75t_L g1825 ( 
.A1(n_1801),
.A2(n_1677),
.B1(n_1661),
.B2(n_1710),
.Y(n_1825)
);

INVx1_ASAP7_75t_L g1826 ( 
.A(n_1779),
.Y(n_1826)
);

INVx1_ASAP7_75t_L g1827 ( 
.A(n_1781),
.Y(n_1827)
);

INVx1_ASAP7_75t_L g1828 ( 
.A(n_1803),
.Y(n_1828)
);

AOI22xp33_ASAP7_75t_L g1829 ( 
.A1(n_1802),
.A2(n_1767),
.B1(n_1797),
.B2(n_1796),
.Y(n_1829)
);

AOI221xp5_ASAP7_75t_L g1830 ( 
.A1(n_1809),
.A2(n_1810),
.B1(n_1811),
.B2(n_1808),
.C(n_1813),
.Y(n_1830)
);

INVx1_ASAP7_75t_L g1831 ( 
.A(n_1804),
.Y(n_1831)
);

O2A1O1Ixp33_ASAP7_75t_L g1832 ( 
.A1(n_1809),
.A2(n_1783),
.B(n_1795),
.C(n_1788),
.Y(n_1832)
);

INVx1_ASAP7_75t_L g1833 ( 
.A(n_1823),
.Y(n_1833)
);

INVxp33_ASAP7_75t_L g1834 ( 
.A(n_1808),
.Y(n_1834)
);

OAI221xp5_ASAP7_75t_SL g1835 ( 
.A1(n_1818),
.A2(n_1785),
.B1(n_1800),
.B2(n_1787),
.C(n_1793),
.Y(n_1835)
);

AOI21xp33_ASAP7_75t_L g1836 ( 
.A1(n_1815),
.A2(n_1791),
.B(n_1798),
.Y(n_1836)
);

OAI21xp33_ASAP7_75t_L g1837 ( 
.A1(n_1807),
.A2(n_1789),
.B(n_1786),
.Y(n_1837)
);

INVx2_ASAP7_75t_L g1838 ( 
.A(n_1819),
.Y(n_1838)
);

OAI221xp5_ASAP7_75t_L g1839 ( 
.A1(n_1824),
.A2(n_1825),
.B1(n_1812),
.B2(n_1806),
.C(n_1822),
.Y(n_1839)
);

INVx1_ASAP7_75t_SL g1840 ( 
.A(n_1819),
.Y(n_1840)
);

OR2x2_ASAP7_75t_L g1841 ( 
.A(n_1814),
.B(n_1799),
.Y(n_1841)
);

INVxp67_ASAP7_75t_L g1842 ( 
.A(n_1823),
.Y(n_1842)
);

NAND2x1_ASAP7_75t_L g1843 ( 
.A(n_1805),
.B(n_1791),
.Y(n_1843)
);

AOI21xp5_ASAP7_75t_L g1844 ( 
.A1(n_1806),
.A2(n_1791),
.B(n_1790),
.Y(n_1844)
);

OAI21xp5_ASAP7_75t_L g1845 ( 
.A1(n_1816),
.A2(n_1782),
.B(n_1677),
.Y(n_1845)
);

AOI22xp33_ASAP7_75t_L g1846 ( 
.A1(n_1817),
.A2(n_1493),
.B1(n_1629),
.B2(n_1627),
.Y(n_1846)
);

OAI21xp5_ASAP7_75t_L g1847 ( 
.A1(n_1820),
.A2(n_1677),
.B(n_1629),
.Y(n_1847)
);

NAND2xp5_ASAP7_75t_L g1848 ( 
.A(n_1840),
.B(n_1821),
.Y(n_1848)
);

INVx1_ASAP7_75t_L g1849 ( 
.A(n_1833),
.Y(n_1849)
);

INVx1_ASAP7_75t_L g1850 ( 
.A(n_1842),
.Y(n_1850)
);

AND2x2_ASAP7_75t_L g1851 ( 
.A(n_1838),
.B(n_1826),
.Y(n_1851)
);

OR2x2_ASAP7_75t_L g1852 ( 
.A(n_1835),
.B(n_1827),
.Y(n_1852)
);

NAND2xp5_ASAP7_75t_L g1853 ( 
.A(n_1830),
.B(n_1717),
.Y(n_1853)
);

NAND2xp5_ASAP7_75t_L g1854 ( 
.A(n_1834),
.B(n_1717),
.Y(n_1854)
);

INVx1_ASAP7_75t_SL g1855 ( 
.A(n_1843),
.Y(n_1855)
);

INVxp67_ASAP7_75t_L g1856 ( 
.A(n_1828),
.Y(n_1856)
);

INVx1_ASAP7_75t_L g1857 ( 
.A(n_1831),
.Y(n_1857)
);

AOI21xp33_ASAP7_75t_L g1858 ( 
.A1(n_1834),
.A2(n_1641),
.B(n_1585),
.Y(n_1858)
);

NAND2xp5_ASAP7_75t_L g1859 ( 
.A(n_1844),
.B(n_1717),
.Y(n_1859)
);

NAND3xp33_ASAP7_75t_L g1860 ( 
.A(n_1852),
.B(n_1832),
.C(n_1829),
.Y(n_1860)
);

NAND2xp5_ASAP7_75t_L g1861 ( 
.A(n_1855),
.B(n_1829),
.Y(n_1861)
);

OAI22xp5_ASAP7_75t_L g1862 ( 
.A1(n_1853),
.A2(n_1839),
.B1(n_1846),
.B2(n_1841),
.Y(n_1862)
);

AOI21xp5_ASAP7_75t_L g1863 ( 
.A1(n_1854),
.A2(n_1836),
.B(n_1837),
.Y(n_1863)
);

NOR3xp33_ASAP7_75t_SL g1864 ( 
.A(n_1848),
.B(n_1845),
.C(n_1847),
.Y(n_1864)
);

INVx1_ASAP7_75t_L g1865 ( 
.A(n_1851),
.Y(n_1865)
);

NOR2x1_ASAP7_75t_L g1866 ( 
.A(n_1850),
.B(n_1849),
.Y(n_1866)
);

NAND2xp5_ASAP7_75t_L g1867 ( 
.A(n_1851),
.B(n_1846),
.Y(n_1867)
);

AOI211xp5_ASAP7_75t_L g1868 ( 
.A1(n_1858),
.A2(n_1856),
.B(n_1859),
.C(n_1857),
.Y(n_1868)
);

CKINVDCx5p33_ASAP7_75t_R g1869 ( 
.A(n_1856),
.Y(n_1869)
);

AOI321xp33_ASAP7_75t_L g1870 ( 
.A1(n_1862),
.A2(n_1627),
.A3(n_1567),
.B1(n_1563),
.B2(n_1721),
.C(n_1633),
.Y(n_1870)
);

AOI22xp5_ASAP7_75t_L g1871 ( 
.A1(n_1860),
.A2(n_1710),
.B1(n_1625),
.B2(n_1578),
.Y(n_1871)
);

AOI221x1_ASAP7_75t_L g1872 ( 
.A1(n_1861),
.A2(n_1718),
.B1(n_1715),
.B2(n_1704),
.C(n_1719),
.Y(n_1872)
);

AOI221xp5_ASAP7_75t_L g1873 ( 
.A1(n_1863),
.A2(n_1721),
.B1(n_1715),
.B2(n_1718),
.C(n_1704),
.Y(n_1873)
);

OAI22xp33_ASAP7_75t_SL g1874 ( 
.A1(n_1869),
.A2(n_1683),
.B1(n_1703),
.B2(n_1690),
.Y(n_1874)
);

NOR3xp33_ASAP7_75t_L g1875 ( 
.A(n_1868),
.B(n_1496),
.C(n_1635),
.Y(n_1875)
);

AND2x2_ASAP7_75t_SL g1876 ( 
.A(n_1875),
.B(n_1865),
.Y(n_1876)
);

AOI22xp5_ASAP7_75t_L g1877 ( 
.A1(n_1871),
.A2(n_1866),
.B1(n_1867),
.B2(n_1864),
.Y(n_1877)
);

AOI322xp5_ASAP7_75t_L g1878 ( 
.A1(n_1873),
.A2(n_1870),
.A3(n_1721),
.B1(n_1874),
.B2(n_1872),
.C1(n_1714),
.C2(n_1685),
.Y(n_1878)
);

INVx1_ASAP7_75t_L g1879 ( 
.A(n_1875),
.Y(n_1879)
);

AND2x2_ASAP7_75t_L g1880 ( 
.A(n_1875),
.B(n_1685),
.Y(n_1880)
);

INVx1_ASAP7_75t_L g1881 ( 
.A(n_1875),
.Y(n_1881)
);

AOI22xp33_ASAP7_75t_L g1882 ( 
.A1(n_1875),
.A2(n_1630),
.B1(n_1625),
.B2(n_1635),
.Y(n_1882)
);

AND2x4_ASAP7_75t_L g1883 ( 
.A(n_1879),
.B(n_1881),
.Y(n_1883)
);

NOR2xp33_ASAP7_75t_L g1884 ( 
.A(n_1877),
.B(n_1704),
.Y(n_1884)
);

INVxp67_ASAP7_75t_L g1885 ( 
.A(n_1877),
.Y(n_1885)
);

OR2x2_ASAP7_75t_L g1886 ( 
.A(n_1880),
.B(n_1683),
.Y(n_1886)
);

NAND4xp75_ASAP7_75t_L g1887 ( 
.A(n_1876),
.B(n_1685),
.C(n_1688),
.D(n_1694),
.Y(n_1887)
);

AND3x2_ASAP7_75t_L g1888 ( 
.A(n_1885),
.B(n_1878),
.C(n_1882),
.Y(n_1888)
);

AOI22xp5_ASAP7_75t_L g1889 ( 
.A1(n_1887),
.A2(n_1625),
.B1(n_1702),
.B2(n_1694),
.Y(n_1889)
);

NOR2x1_ASAP7_75t_L g1890 ( 
.A(n_1883),
.B(n_1715),
.Y(n_1890)
);

NOR2x1_ASAP7_75t_L g1891 ( 
.A(n_1890),
.B(n_1884),
.Y(n_1891)
);

INVx1_ASAP7_75t_L g1892 ( 
.A(n_1891),
.Y(n_1892)
);

XOR2x1_ASAP7_75t_L g1893 ( 
.A(n_1892),
.B(n_1888),
.Y(n_1893)
);

OAI22xp33_ASAP7_75t_L g1894 ( 
.A1(n_1892),
.A2(n_1886),
.B1(n_1889),
.B2(n_1683),
.Y(n_1894)
);

INVx2_ASAP7_75t_L g1895 ( 
.A(n_1893),
.Y(n_1895)
);

INVx2_ASAP7_75t_L g1896 ( 
.A(n_1894),
.Y(n_1896)
);

AOI22x1_ASAP7_75t_L g1897 ( 
.A1(n_1895),
.A2(n_1718),
.B1(n_1715),
.B2(n_1496),
.Y(n_1897)
);

OAI21xp5_ASAP7_75t_L g1898 ( 
.A1(n_1896),
.A2(n_1718),
.B(n_1703),
.Y(n_1898)
);

OAI22xp5_ASAP7_75t_L g1899 ( 
.A1(n_1898),
.A2(n_1703),
.B1(n_1690),
.B2(n_1712),
.Y(n_1899)
);

AOI22xp5_ASAP7_75t_L g1900 ( 
.A1(n_1899),
.A2(n_1897),
.B1(n_1703),
.B2(n_1694),
.Y(n_1900)
);

OAI22xp33_ASAP7_75t_L g1901 ( 
.A1(n_1900),
.A2(n_1690),
.B1(n_1712),
.B2(n_1719),
.Y(n_1901)
);

OAI221xp5_ASAP7_75t_R g1902 ( 
.A1(n_1901),
.A2(n_1580),
.B1(n_1702),
.B2(n_1688),
.C(n_1714),
.Y(n_1902)
);

AOI211xp5_ASAP7_75t_L g1903 ( 
.A1(n_1902),
.A2(n_1530),
.B(n_1527),
.C(n_1537),
.Y(n_1903)
);


endmodule