module fake_ariane_2602_n_2793 (n_295, n_356, n_170, n_190, n_160, n_64, n_180, n_119, n_124, n_386, n_307, n_332, n_294, n_197, n_176, n_34, n_404, n_172, n_347, n_423, n_183, n_373, n_299, n_12, n_133, n_66, n_205, n_341, n_71, n_109, n_245, n_421, n_96, n_319, n_49, n_20, n_416, n_283, n_50, n_187, n_367, n_345, n_374, n_318, n_103, n_244, n_226, n_220, n_261, n_36, n_370, n_189, n_72, n_286, n_57, n_424, n_387, n_406, n_117, n_139, n_85, n_130, n_349, n_391, n_346, n_214, n_348, n_2, n_32, n_410, n_379, n_138, n_162, n_264, n_137, n_122, n_198, n_232, n_52, n_385, n_73, n_327, n_77, n_372, n_377, n_15, n_396, n_23, n_399, n_87, n_279, n_207, n_363, n_354, n_41, n_140, n_419, n_151, n_28, n_146, n_230, n_270, n_194, n_154, n_338, n_142, n_285, n_186, n_202, n_145, n_193, n_59, n_336, n_315, n_311, n_239, n_402, n_35, n_272, n_54, n_8, n_339, n_167, n_90, n_38, n_422, n_47, n_153, n_18, n_269, n_75, n_158, n_69, n_259, n_95, n_143, n_152, n_405, n_120, n_169, n_106, n_173, n_242, n_309, n_320, n_115, n_331, n_401, n_267, n_335, n_350, n_291, n_344, n_381, n_398, n_62, n_210, n_200, n_166, n_253, n_218, n_79, n_3, n_271, n_247, n_91, n_240, n_369, n_128, n_224, n_44, n_82, n_31, n_420, n_222, n_256, n_326, n_227, n_48, n_188, n_323, n_330, n_400, n_11, n_129, n_126, n_282, n_328, n_368, n_277, n_248, n_301, n_293, n_228, n_325, n_276, n_93, n_108, n_303, n_168, n_81, n_1, n_206, n_352, n_238, n_365, n_136, n_334, n_192, n_300, n_14, n_163, n_88, n_141, n_390, n_104, n_314, n_16, n_273, n_305, n_312, n_233, n_56, n_60, n_388, n_333, n_413, n_392, n_376, n_221, n_321, n_86, n_361, n_89, n_149, n_383, n_237, n_175, n_74, n_19, n_40, n_181, n_53, n_260, n_362, n_310, n_236, n_281, n_24, n_7, n_209, n_262, n_17, n_225, n_235, n_297, n_290, n_46, n_84, n_371, n_199, n_107, n_217, n_178, n_42, n_308, n_417, n_201, n_70, n_343, n_10, n_414, n_287, n_302, n_380, n_6, n_94, n_284, n_4, n_249, n_37, n_58, n_65, n_123, n_212, n_355, n_278, n_255, n_257, n_148, n_135, n_409, n_171, n_384, n_61, n_102, n_182, n_316, n_196, n_125, n_43, n_407, n_13, n_27, n_254, n_219, n_55, n_231, n_366, n_234, n_280, n_215, n_252, n_161, n_298, n_68, n_415, n_78, n_63, n_99, n_216, n_5, n_418, n_223, n_403, n_25, n_83, n_389, n_288, n_179, n_395, n_195, n_213, n_110, n_304, n_67, n_306, n_313, n_92, n_203, n_378, n_150, n_98, n_375, n_113, n_114, n_33, n_324, n_337, n_111, n_21, n_274, n_296, n_265, n_208, n_156, n_292, n_174, n_275, n_100, n_132, n_147, n_204, n_51, n_76, n_342, n_26, n_246, n_0, n_159, n_358, n_105, n_30, n_131, n_263, n_360, n_229, n_394, n_250, n_165, n_144, n_317, n_101, n_243, n_134, n_329, n_185, n_340, n_289, n_9, n_112, n_45, n_268, n_266, n_164, n_157, n_184, n_177, n_364, n_258, n_425, n_118, n_121, n_411, n_353, n_22, n_241, n_29, n_357, n_412, n_191, n_382, n_80, n_211, n_97, n_408, n_322, n_251, n_116, n_397, n_351, n_39, n_393, n_359, n_155, n_127, n_2793);

input n_295;
input n_356;
input n_170;
input n_190;
input n_160;
input n_64;
input n_180;
input n_119;
input n_124;
input n_386;
input n_307;
input n_332;
input n_294;
input n_197;
input n_176;
input n_34;
input n_404;
input n_172;
input n_347;
input n_423;
input n_183;
input n_373;
input n_299;
input n_12;
input n_133;
input n_66;
input n_205;
input n_341;
input n_71;
input n_109;
input n_245;
input n_421;
input n_96;
input n_319;
input n_49;
input n_20;
input n_416;
input n_283;
input n_50;
input n_187;
input n_367;
input n_345;
input n_374;
input n_318;
input n_103;
input n_244;
input n_226;
input n_220;
input n_261;
input n_36;
input n_370;
input n_189;
input n_72;
input n_286;
input n_57;
input n_424;
input n_387;
input n_406;
input n_117;
input n_139;
input n_85;
input n_130;
input n_349;
input n_391;
input n_346;
input n_214;
input n_348;
input n_2;
input n_32;
input n_410;
input n_379;
input n_138;
input n_162;
input n_264;
input n_137;
input n_122;
input n_198;
input n_232;
input n_52;
input n_385;
input n_73;
input n_327;
input n_77;
input n_372;
input n_377;
input n_15;
input n_396;
input n_23;
input n_399;
input n_87;
input n_279;
input n_207;
input n_363;
input n_354;
input n_41;
input n_140;
input n_419;
input n_151;
input n_28;
input n_146;
input n_230;
input n_270;
input n_194;
input n_154;
input n_338;
input n_142;
input n_285;
input n_186;
input n_202;
input n_145;
input n_193;
input n_59;
input n_336;
input n_315;
input n_311;
input n_239;
input n_402;
input n_35;
input n_272;
input n_54;
input n_8;
input n_339;
input n_167;
input n_90;
input n_38;
input n_422;
input n_47;
input n_153;
input n_18;
input n_269;
input n_75;
input n_158;
input n_69;
input n_259;
input n_95;
input n_143;
input n_152;
input n_405;
input n_120;
input n_169;
input n_106;
input n_173;
input n_242;
input n_309;
input n_320;
input n_115;
input n_331;
input n_401;
input n_267;
input n_335;
input n_350;
input n_291;
input n_344;
input n_381;
input n_398;
input n_62;
input n_210;
input n_200;
input n_166;
input n_253;
input n_218;
input n_79;
input n_3;
input n_271;
input n_247;
input n_91;
input n_240;
input n_369;
input n_128;
input n_224;
input n_44;
input n_82;
input n_31;
input n_420;
input n_222;
input n_256;
input n_326;
input n_227;
input n_48;
input n_188;
input n_323;
input n_330;
input n_400;
input n_11;
input n_129;
input n_126;
input n_282;
input n_328;
input n_368;
input n_277;
input n_248;
input n_301;
input n_293;
input n_228;
input n_325;
input n_276;
input n_93;
input n_108;
input n_303;
input n_168;
input n_81;
input n_1;
input n_206;
input n_352;
input n_238;
input n_365;
input n_136;
input n_334;
input n_192;
input n_300;
input n_14;
input n_163;
input n_88;
input n_141;
input n_390;
input n_104;
input n_314;
input n_16;
input n_273;
input n_305;
input n_312;
input n_233;
input n_56;
input n_60;
input n_388;
input n_333;
input n_413;
input n_392;
input n_376;
input n_221;
input n_321;
input n_86;
input n_361;
input n_89;
input n_149;
input n_383;
input n_237;
input n_175;
input n_74;
input n_19;
input n_40;
input n_181;
input n_53;
input n_260;
input n_362;
input n_310;
input n_236;
input n_281;
input n_24;
input n_7;
input n_209;
input n_262;
input n_17;
input n_225;
input n_235;
input n_297;
input n_290;
input n_46;
input n_84;
input n_371;
input n_199;
input n_107;
input n_217;
input n_178;
input n_42;
input n_308;
input n_417;
input n_201;
input n_70;
input n_343;
input n_10;
input n_414;
input n_287;
input n_302;
input n_380;
input n_6;
input n_94;
input n_284;
input n_4;
input n_249;
input n_37;
input n_58;
input n_65;
input n_123;
input n_212;
input n_355;
input n_278;
input n_255;
input n_257;
input n_148;
input n_135;
input n_409;
input n_171;
input n_384;
input n_61;
input n_102;
input n_182;
input n_316;
input n_196;
input n_125;
input n_43;
input n_407;
input n_13;
input n_27;
input n_254;
input n_219;
input n_55;
input n_231;
input n_366;
input n_234;
input n_280;
input n_215;
input n_252;
input n_161;
input n_298;
input n_68;
input n_415;
input n_78;
input n_63;
input n_99;
input n_216;
input n_5;
input n_418;
input n_223;
input n_403;
input n_25;
input n_83;
input n_389;
input n_288;
input n_179;
input n_395;
input n_195;
input n_213;
input n_110;
input n_304;
input n_67;
input n_306;
input n_313;
input n_92;
input n_203;
input n_378;
input n_150;
input n_98;
input n_375;
input n_113;
input n_114;
input n_33;
input n_324;
input n_337;
input n_111;
input n_21;
input n_274;
input n_296;
input n_265;
input n_208;
input n_156;
input n_292;
input n_174;
input n_275;
input n_100;
input n_132;
input n_147;
input n_204;
input n_51;
input n_76;
input n_342;
input n_26;
input n_246;
input n_0;
input n_159;
input n_358;
input n_105;
input n_30;
input n_131;
input n_263;
input n_360;
input n_229;
input n_394;
input n_250;
input n_165;
input n_144;
input n_317;
input n_101;
input n_243;
input n_134;
input n_329;
input n_185;
input n_340;
input n_289;
input n_9;
input n_112;
input n_45;
input n_268;
input n_266;
input n_164;
input n_157;
input n_184;
input n_177;
input n_364;
input n_258;
input n_425;
input n_118;
input n_121;
input n_411;
input n_353;
input n_22;
input n_241;
input n_29;
input n_357;
input n_412;
input n_191;
input n_382;
input n_80;
input n_211;
input n_97;
input n_408;
input n_322;
input n_251;
input n_116;
input n_397;
input n_351;
input n_39;
input n_393;
input n_359;
input n_155;
input n_127;

output n_2793;

wire n_2752;
wire n_913;
wire n_1681;
wire n_2163;
wire n_1486;
wire n_1507;
wire n_1938;
wire n_589;
wire n_2484;
wire n_1174;
wire n_2346;
wire n_1469;
wire n_691;
wire n_1353;
wire n_2679;
wire n_1355;
wire n_2131;
wire n_2559;
wire n_2500;
wire n_2509;
wire n_1383;
wire n_2182;
wire n_603;
wire n_2135;
wire n_2334;
wire n_2680;
wire n_1250;
wire n_2030;
wire n_1169;
wire n_789;
wire n_850;
wire n_1916;
wire n_610;
wire n_1713;
wire n_1436;
wire n_2407;
wire n_690;
wire n_1109;
wire n_1430;
wire n_2537;
wire n_525;
wire n_2002;
wire n_1463;
wire n_2243;
wire n_1238;
wire n_2694;
wire n_2011;
wire n_2729;
wire n_1515;
wire n_817;
wire n_1837;
wire n_924;
wire n_781;
wire n_2013;
wire n_2786;
wire n_1566;
wire n_717;
wire n_2006;
wire n_952;
wire n_864;
wire n_2446;
wire n_1096;
wire n_1379;
wire n_2436;
wire n_2376;
wire n_2367;
wire n_2671;
wire n_2790;
wire n_1706;
wire n_2207;
wire n_2461;
wire n_2702;
wire n_524;
wire n_2731;
wire n_1214;
wire n_634;
wire n_1839;
wire n_1246;
wire n_1138;
wire n_2042;
wire n_2123;
wire n_1853;
wire n_2238;
wire n_1503;
wire n_764;
wire n_2529;
wire n_2374;
wire n_462;
wire n_1196;
wire n_1181;
wire n_1999;
wire n_2380;
wire n_1187;
wire n_1131;
wire n_1225;
wire n_2646;
wire n_737;
wire n_1298;
wire n_2653;
wire n_1745;
wire n_1366;
wire n_2084;
wire n_568;
wire n_2278;
wire n_1088;
wire n_1424;
wire n_766;
wire n_1835;
wire n_1457;
wire n_2482;
wire n_1682;
wire n_2750;
wire n_1836;
wire n_520;
wire n_870;
wire n_2547;
wire n_1453;
wire n_958;
wire n_945;
wire n_2554;
wire n_2248;
wire n_813;
wire n_1985;
wire n_2288;
wire n_2621;
wire n_995;
wire n_2579;
wire n_1909;
wire n_2156;
wire n_1184;
wire n_1961;
wire n_1535;
wire n_500;
wire n_665;
wire n_754;
wire n_903;
wire n_871;
wire n_2323;
wire n_1073;
wire n_1979;
wire n_1277;
wire n_2107;
wire n_1746;
wire n_1761;
wire n_829;
wire n_1062;
wire n_738;
wire n_1690;
wire n_2221;
wire n_672;
wire n_740;
wire n_1283;
wire n_2317;
wire n_1974;
wire n_1736;
wire n_1018;
wire n_2342;
wire n_2200;
wire n_2781;
wire n_2442;
wire n_2735;
wire n_953;
wire n_1364;
wire n_2390;
wire n_1888;
wire n_1224;
wire n_2109;
wire n_1425;
wire n_2634;
wire n_2709;
wire n_625;
wire n_557;
wire n_2322;
wire n_2746;
wire n_1107;
wire n_1688;
wire n_989;
wire n_1944;
wire n_645;
wire n_559;
wire n_2233;
wire n_2370;
wire n_2663;
wire n_495;
wire n_1988;
wire n_795;
wire n_721;
wire n_1084;
wire n_1718;
wire n_1276;
wire n_1936;
wire n_2149;
wire n_2277;
wire n_1428;
wire n_1284;
wire n_1241;
wire n_821;
wire n_561;
wire n_770;
wire n_1514;
wire n_2539;
wire n_1528;
wire n_507;
wire n_486;
wire n_901;
wire n_2782;
wire n_569;
wire n_2078;
wire n_1145;
wire n_971;
wire n_2359;
wire n_2201;
wire n_787;
wire n_1650;
wire n_1519;
wire n_1195;
wire n_2049;
wire n_1522;
wire n_518;
wire n_1207;
wire n_786;
wire n_1404;
wire n_868;
wire n_2232;
wire n_1847;
wire n_2458;
wire n_2779;
wire n_1542;
wire n_1314;
wire n_1512;
wire n_2227;
wire n_2301;
wire n_1539;
wire n_884;
wire n_1851;
wire n_2162;
wire n_1415;
wire n_1034;
wire n_1652;
wire n_2192;
wire n_1676;
wire n_1085;
wire n_1636;
wire n_432;
wire n_823;
wire n_1900;
wire n_620;
wire n_1074;
wire n_859;
wire n_1765;
wire n_1889;
wire n_587;
wire n_1977;
wire n_693;
wire n_863;
wire n_2650;
wire n_1254;
wire n_929;
wire n_2433;
wire n_1703;
wire n_899;
wire n_2332;
wire n_2391;
wire n_611;
wire n_1295;
wire n_2060;
wire n_1850;
wire n_2004;
wire n_1013;
wire n_1495;
wire n_1637;
wire n_2571;
wire n_2427;
wire n_661;
wire n_2098;
wire n_2616;
wire n_1751;
wire n_533;
wire n_1917;
wire n_2456;
wire n_2769;
wire n_1924;
wire n_438;
wire n_1654;
wire n_1560;
wire n_2341;
wire n_1548;
wire n_1811;
wire n_2045;
wire n_440;
wire n_2575;
wire n_2722;
wire n_1396;
wire n_1230;
wire n_612;
wire n_1840;
wire n_2739;
wire n_512;
wire n_1597;
wire n_1771;
wire n_1544;
wire n_579;
wire n_844;
wire n_1012;
wire n_1267;
wire n_2061;
wire n_2685;
wire n_2094;
wire n_2512;
wire n_1354;
wire n_1790;
wire n_1213;
wire n_2382;
wire n_2043;
wire n_780;
wire n_2349;
wire n_1918;
wire n_2788;
wire n_1021;
wire n_1443;
wire n_491;
wire n_2595;
wire n_1465;
wire n_2686;
wire n_1949;
wire n_1595;
wire n_1142;
wire n_1140;
wire n_705;
wire n_570;
wire n_2727;
wire n_942;
wire n_1437;
wire n_2077;
wire n_1378;
wire n_461;
wire n_1121;
wire n_1416;
wire n_490;
wire n_1461;
wire n_2717;
wire n_1391;
wire n_1947;
wire n_1599;
wire n_1876;
wire n_1006;
wire n_1830;
wire n_575;
wire n_546;
wire n_503;
wire n_2527;
wire n_1112;
wire n_700;
wire n_1159;
wire n_772;
wire n_1216;
wire n_2759;
wire n_1245;
wire n_2743;
wire n_1669;
wire n_1675;
wire n_2466;
wire n_676;
wire n_2038;
wire n_2263;
wire n_2568;
wire n_2116;
wire n_2271;
wire n_2145;
wire n_2326;
wire n_1838;
wire n_1594;
wire n_680;
wire n_1935;
wire n_1716;
wire n_1872;
wire n_1585;
wire n_2281;
wire n_1432;
wire n_2245;
wire n_1108;
wire n_851;
wire n_444;
wire n_1590;
wire n_1351;
wire n_2216;
wire n_1274;
wire n_2426;
wire n_652;
wire n_1819;
wire n_475;
wire n_947;
wire n_2134;
wire n_1260;
wire n_930;
wire n_1179;
wire n_468;
wire n_2703;
wire n_696;
wire n_1442;
wire n_482;
wire n_2620;
wire n_798;
wire n_1833;
wire n_577;
wire n_1691;
wire n_916;
wire n_1386;
wire n_1884;
wire n_912;
wire n_460;
wire n_1555;
wire n_1842;
wire n_2499;
wire n_2549;
wire n_762;
wire n_1253;
wire n_1468;
wire n_1661;
wire n_2791;
wire n_555;
wire n_2683;
wire n_804;
wire n_1656;
wire n_1382;
wire n_992;
wire n_966;
wire n_955;
wire n_1182;
wire n_794;
wire n_2166;
wire n_1692;
wire n_2611;
wire n_1562;
wire n_514;
wire n_2748;
wire n_2185;
wire n_2398;
wire n_1376;
wire n_513;
wire n_1292;
wire n_1178;
wire n_2015;
wire n_1972;
wire n_1435;
wire n_1750;
wire n_1026;
wire n_1506;
wire n_1610;
wire n_2202;
wire n_2072;
wire n_2415;
wire n_2693;
wire n_436;
wire n_2745;
wire n_2087;
wire n_931;
wire n_1491;
wire n_669;
wire n_2628;
wire n_619;
wire n_437;
wire n_967;
wire n_1083;
wire n_2161;
wire n_1418;
wire n_746;
wire n_1357;
wire n_1079;
wire n_1787;
wire n_2462;
wire n_1389;
wire n_2155;
wire n_2659;
wire n_615;
wire n_1139;
wire n_2439;
wire n_517;
wire n_1312;
wire n_1717;
wire n_1812;
wire n_824;
wire n_428;
wire n_2172;
wire n_2601;
wire n_892;
wire n_1880;
wire n_959;
wire n_2365;
wire n_2257;
wire n_1399;
wire n_1101;
wire n_1567;
wire n_1343;
wire n_563;
wire n_2219;
wire n_1855;
wire n_2100;
wire n_2333;
wire n_990;
wire n_1623;
wire n_1903;
wire n_867;
wire n_2147;
wire n_2435;
wire n_1226;
wire n_2224;
wire n_944;
wire n_749;
wire n_1932;
wire n_1780;
wire n_1970;
wire n_1920;
wire n_2083;
wire n_815;
wire n_542;
wire n_2167;
wire n_2293;
wire n_2753;
wire n_1340;
wire n_470;
wire n_2668;
wire n_1240;
wire n_1087;
wire n_2701;
wire n_2400;
wire n_632;
wire n_477;
wire n_650;
wire n_2388;
wire n_2273;
wire n_2712;
wire n_1433;
wire n_1911;
wire n_2567;
wire n_2557;
wire n_2695;
wire n_1825;
wire n_1908;
wire n_1155;
wire n_2598;
wire n_1071;
wire n_2755;
wire n_712;
wire n_976;
wire n_909;
wire n_1832;
wire n_767;
wire n_1392;
wire n_2682;
wire n_1841;
wire n_1680;
wire n_2066;
wire n_2302;
wire n_2762;
wire n_964;
wire n_1627;
wire n_2220;
wire n_489;
wire n_2294;
wire n_2274;
wire n_974;
wire n_506;
wire n_1731;
wire n_799;
wire n_1147;
wire n_2378;
wire n_2467;
wire n_2768;
wire n_471;
wire n_965;
wire n_1914;
wire n_2253;
wire n_934;
wire n_2213;
wire n_1447;
wire n_2363;
wire n_1220;
wire n_2019;
wire n_698;
wire n_2728;
wire n_2130;
wire n_1674;
wire n_2021;
wire n_2025;
wire n_2160;
wire n_1992;
wire n_1209;
wire n_1020;
wire n_1563;
wire n_646;
wire n_2507;
wire n_2142;
wire n_1633;
wire n_2625;
wire n_1913;
wire n_2069;
wire n_2495;
wire n_1058;
wire n_2328;
wire n_2434;
wire n_1042;
wire n_1234;
wire n_2311;
wire n_479;
wire n_1578;
wire n_2261;
wire n_1455;
wire n_2287;
wire n_836;
wire n_2223;
wire n_1279;
wire n_2473;
wire n_2144;
wire n_2511;
wire n_564;
wire n_1029;
wire n_2649;
wire n_1247;
wire n_760;
wire n_522;
wire n_2438;
wire n_1568;
wire n_1483;
wire n_1363;
wire n_2681;
wire n_1111;
wire n_970;
wire n_1689;
wire n_2535;
wire n_713;
wire n_1255;
wire n_2632;
wire n_1646;
wire n_598;
wire n_2262;
wire n_2565;
wire n_1237;
wire n_927;
wire n_1095;
wire n_1728;
wire n_2335;
wire n_2120;
wire n_706;
wire n_2631;
wire n_1401;
wire n_1419;
wire n_1531;
wire n_776;
wire n_2041;
wire n_2113;
wire n_1933;
wire n_1651;
wire n_2697;
wire n_1387;
wire n_466;
wire n_1263;
wire n_1817;
wire n_2404;
wire n_2168;
wire n_2757;
wire n_552;
wire n_2312;
wire n_670;
wire n_2677;
wire n_1826;
wire n_2483;
wire n_441;
wire n_1951;
wire n_2490;
wire n_1032;
wire n_2558;
wire n_1217;
wire n_1496;
wire n_637;
wire n_1592;
wire n_2662;
wire n_1259;
wire n_1177;
wire n_2655;
wire n_1231;
wire n_2132;
wire n_980;
wire n_1618;
wire n_1869;
wire n_1743;
wire n_905;
wire n_2718;
wire n_720;
wire n_926;
wire n_1943;
wire n_2687;
wire n_2296;
wire n_1802;
wire n_2178;
wire n_2112;
wire n_2765;
wire n_1163;
wire n_2640;
wire n_1795;
wire n_1384;
wire n_2237;
wire n_2146;
wire n_1868;
wire n_1501;
wire n_2241;
wire n_2373;
wire n_1173;
wire n_2350;
wire n_1068;
wire n_1198;
wire n_2531;
wire n_1570;
wire n_2099;
wire n_487;
wire n_1518;
wire n_1456;
wire n_1879;
wire n_1886;
wire n_1648;
wire n_2187;
wire n_1413;
wire n_2617;
wire n_2481;
wire n_2129;
wire n_855;
wire n_2327;
wire n_808;
wire n_1365;
wire n_2476;
wire n_553;
wire n_2059;
wire n_2437;
wire n_2636;
wire n_1439;
wire n_814;
wire n_578;
wire n_2074;
wire n_1665;
wire n_1287;
wire n_1611;
wire n_2122;
wire n_2399;
wire n_1414;
wire n_2067;
wire n_1134;
wire n_1484;
wire n_1901;
wire n_647;
wire n_2055;
wire n_2027;
wire n_1423;
wire n_2117;
wire n_600;
wire n_1609;
wire n_1053;
wire n_481;
wire n_1939;
wire n_2308;
wire n_2242;
wire n_1906;
wire n_1899;
wire n_529;
wire n_2195;
wire n_502;
wire n_2194;
wire n_1467;
wire n_1828;
wire n_2159;
wire n_1798;
wire n_1608;
wire n_1304;
wire n_1744;
wire n_2267;
wire n_1105;
wire n_547;
wire n_439;
wire n_677;
wire n_604;
wire n_478;
wire n_703;
wire n_1349;
wire n_1709;
wire n_1061;
wire n_2102;
wire n_681;
wire n_874;
wire n_2286;
wire n_2023;
wire n_1278;
wire n_707;
wire n_983;
wire n_2783;
wire n_2599;
wire n_699;
wire n_2075;
wire n_727;
wire n_1726;
wire n_590;
wire n_2523;
wire n_1945;
wire n_1015;
wire n_545;
wire n_2418;
wire n_1377;
wire n_1162;
wire n_536;
wire n_1614;
wire n_2031;
wire n_2496;
wire n_2118;
wire n_1740;
wire n_1602;
wire n_688;
wire n_636;
wire n_427;
wire n_1098;
wire n_1490;
wire n_2338;
wire n_442;
wire n_777;
wire n_1553;
wire n_1080;
wire n_920;
wire n_1760;
wire n_1086;
wire n_1092;
wire n_2225;
wire n_986;
wire n_1104;
wire n_1963;
wire n_887;
wire n_729;
wire n_2218;
wire n_2057;
wire n_1122;
wire n_1205;
wire n_1408;
wire n_2593;
wire n_1693;
wire n_2125;
wire n_2716;
wire n_1132;
wire n_1156;
wire n_2741;
wire n_501;
wire n_2184;
wire n_2714;
wire n_1823;
wire n_2780;
wire n_1120;
wire n_1202;
wire n_627;
wire n_2254;
wire n_1188;
wire n_1498;
wire n_1371;
wire n_2033;
wire n_2618;
wire n_1402;
wire n_957;
wire n_1242;
wire n_2754;
wire n_2707;
wire n_2774;
wire n_1607;
wire n_1489;
wire n_1218;
wire n_2756;
wire n_2217;
wire n_2226;
wire n_1586;
wire n_861;
wire n_1543;
wire n_1431;
wire n_877;
wire n_1119;
wire n_1863;
wire n_1763;
wire n_1666;
wire n_1500;
wire n_616;
wire n_2214;
wire n_1055;
wire n_1395;
wire n_1346;
wire n_2763;
wire n_2256;
wire n_1189;
wire n_1089;
wire n_1859;
wire n_2660;
wire n_1502;
wire n_1523;
wire n_2190;
wire n_1478;
wire n_2732;
wire n_1883;
wire n_2516;
wire n_2776;
wire n_2555;
wire n_1969;
wire n_2708;
wire n_735;
wire n_1005;
wire n_527;
wire n_2379;
wire n_1294;
wire n_2661;
wire n_1667;
wire n_845;
wire n_888;
wire n_2300;
wire n_1649;
wire n_2452;
wire n_1677;
wire n_2470;
wire n_1927;
wire n_1297;
wire n_551;
wire n_1708;
wire n_1222;
wire n_2284;
wire n_1844;
wire n_2283;
wire n_582;
wire n_2526;
wire n_1957;
wire n_1953;
wire n_2643;
wire n_755;
wire n_1097;
wire n_1219;
wire n_1711;
wire n_710;
wire n_1919;
wire n_534;
wire n_1791;
wire n_2508;
wire n_2124;
wire n_1894;
wire n_1460;
wire n_1239;
wire n_2594;
wire n_2266;
wire n_2449;
wire n_560;
wire n_890;
wire n_842;
wire n_1898;
wire n_451;
wire n_745;
wire n_1741;
wire n_1572;
wire n_1907;
wire n_1793;
wire n_742;
wire n_1975;
wire n_1081;
wire n_1373;
wire n_1388;
wire n_1266;
wire n_1540;
wire n_1719;
wire n_2119;
wire n_2742;
wire n_769;
wire n_1797;
wire n_2366;
wire n_2493;
wire n_1753;
wire n_1990;
wire n_1372;
wire n_476;
wire n_832;
wire n_535;
wire n_744;
wire n_1895;
wire n_2690;
wire n_2474;
wire n_2623;
wire n_982;
wire n_1800;
wire n_915;
wire n_1075;
wire n_2008;
wire n_454;
wire n_1331;
wire n_1890;
wire n_1529;
wire n_1227;
wire n_2127;
wire n_655;
wire n_1734;
wire n_1860;
wire n_2785;
wire n_2460;
wire n_1007;
wire n_1580;
wire n_1319;
wire n_657;
wire n_837;
wire n_812;
wire n_2448;
wire n_2211;
wire n_2292;
wire n_2480;
wire n_606;
wire n_951;
wire n_2772;
wire n_862;
wire n_1700;
wire n_2637;
wire n_659;
wire n_1332;
wire n_2306;
wire n_509;
wire n_1854;
wire n_666;
wire n_1747;
wire n_2071;
wire n_2424;
wire n_430;
wire n_1206;
wire n_1729;
wire n_722;
wire n_1508;
wire n_2414;
wire n_2082;
wire n_1532;
wire n_1171;
wire n_1030;
wire n_785;
wire n_2389;
wire n_1309;
wire n_999;
wire n_2280;
wire n_1766;
wire n_1338;
wire n_1342;
wire n_2737;
wire n_456;
wire n_1867;
wire n_852;
wire n_1394;
wire n_2576;
wire n_704;
wire n_1060;
wire n_1044;
wire n_1714;
wire n_2696;
wire n_521;
wire n_2140;
wire n_873;
wire n_1748;
wire n_1301;
wire n_2157;
wire n_1966;
wire n_1243;
wire n_2171;
wire n_2468;
wire n_1400;
wire n_2035;
wire n_2614;
wire n_1466;
wire n_1513;
wire n_1527;
wire n_2581;
wire n_1783;
wire n_608;
wire n_2494;
wire n_1538;
wire n_2457;
wire n_2128;
wire n_1037;
wire n_1329;
wire n_1993;
wire n_1545;
wire n_2629;
wire n_1257;
wire n_1480;
wire n_1954;
wire n_1668;
wire n_1878;
wire n_2540;
wire n_1605;
wire n_1078;
wire n_2486;
wire n_1897;
wire n_2520;
wire n_2137;
wire n_1161;
wire n_2489;
wire n_811;
wire n_624;
wire n_876;
wire n_791;
wire n_618;
wire n_1191;
wire n_2492;
wire n_736;
wire n_1025;
wire n_1215;
wire n_1449;
wire n_2337;
wire n_2265;
wire n_687;
wire n_797;
wire n_2026;
wire n_1786;
wire n_2627;
wire n_480;
wire n_1327;
wire n_1475;
wire n_642;
wire n_1804;
wire n_2106;
wire n_1406;
wire n_595;
wire n_1405;
wire n_2684;
wire n_2726;
wire n_602;
wire n_2622;
wire n_2272;
wire n_1757;
wire n_592;
wire n_1499;
wire n_1318;
wire n_854;
wire n_2091;
wire n_1632;
wire n_1769;
wire n_474;
wire n_1929;
wire n_1950;
wire n_2264;
wire n_2691;
wire n_805;
wire n_2032;
wire n_2090;
wire n_1658;
wire n_2249;
wire n_1072;
wire n_695;
wire n_1526;
wire n_1305;
wire n_730;
wire n_1596;
wire n_2348;
wire n_2656;
wire n_1281;
wire n_516;
wire n_2364;
wire n_1997;
wire n_2574;
wire n_1137;
wire n_1873;
wire n_1258;
wire n_1733;
wire n_463;
wire n_1476;
wire n_1524;
wire n_1856;
wire n_2016;
wire n_640;
wire n_2667;
wire n_2725;
wire n_943;
wire n_1118;
wire n_678;
wire n_651;
wire n_1874;
wire n_1293;
wire n_961;
wire n_469;
wire n_1807;
wire n_1046;
wire n_1123;
wire n_726;
wire n_1657;
wire n_878;
wire n_1784;
wire n_771;
wire n_1321;
wire n_752;
wire n_2307;
wire n_1488;
wire n_985;
wire n_1330;
wire n_906;
wire n_1180;
wire n_1697;
wire n_2295;
wire n_2730;
wire n_806;
wire n_1984;
wire n_1350;
wire n_1556;
wire n_1561;
wire n_649;
wire n_2412;
wire n_2720;
wire n_1352;
wire n_2405;
wire n_1824;
wire n_643;
wire n_2606;
wire n_2700;
wire n_1492;
wire n_2383;
wire n_2764;
wire n_1441;
wire n_1822;
wire n_682;
wire n_1616;
wire n_2633;
wire n_2416;
wire n_819;
wire n_2386;
wire n_1971;
wire n_1429;
wire n_1324;
wire n_2064;
wire n_2353;
wire n_586;
wire n_2528;
wire n_1778;
wire n_1776;
wire n_686;
wire n_605;
wire n_1154;
wire n_584;
wire n_1557;
wire n_1759;
wire n_1829;
wire n_2325;
wire n_1130;
wire n_1450;
wire n_756;
wire n_2022;
wire n_1016;
wire n_2298;
wire n_1149;
wire n_1505;
wire n_2408;
wire n_2698;
wire n_2320;
wire n_979;
wire n_2329;
wire n_2570;
wire n_1642;
wire n_2417;
wire n_2789;
wire n_2525;
wire n_1815;
wire n_897;
wire n_2546;
wire n_949;
wire n_2454;
wire n_1493;
wire n_515;
wire n_807;
wire n_891;
wire n_885;
wire n_1659;
wire n_2354;
wire n_1864;
wire n_2760;
wire n_1887;
wire n_1208;
wire n_1987;
wire n_2368;
wire n_802;
wire n_1151;
wire n_554;
wire n_960;
wire n_2352;
wire n_2502;
wire n_1256;
wire n_714;
wire n_2170;
wire n_790;
wire n_2244;
wire n_2143;
wire n_2393;
wire n_725;
wire n_2377;
wire n_1577;
wire n_1448;
wire n_2198;
wire n_1009;
wire n_2652;
wire n_1133;
wire n_883;
wire n_473;
wire n_1852;
wire n_801;
wire n_1286;
wire n_2612;
wire n_818;
wire n_1685;
wire n_779;
wire n_2410;
wire n_2314;
wire n_2477;
wire n_2279;
wire n_594;
wire n_2222;
wire n_1995;
wire n_1877;
wire n_1397;
wire n_1052;
wire n_1333;
wire n_1306;
wire n_1849;
wire n_2203;
wire n_2133;
wire n_2076;
wire n_833;
wire n_1426;
wire n_2250;
wire n_2497;
wire n_2247;
wire n_2230;
wire n_879;
wire n_1117;
wire n_1269;
wire n_1303;
wire n_1547;
wire n_1438;
wire n_1541;
wire n_597;
wire n_2001;
wire n_1047;
wire n_2506;
wire n_1472;
wire n_2413;
wire n_1593;
wire n_2610;
wire n_1050;
wire n_2626;
wire n_566;
wire n_2158;
wire n_2578;
wire n_2607;
wire n_2285;
wire n_1288;
wire n_2605;
wire n_1201;
wire n_858;
wire n_1185;
wire n_2475;
wire n_2173;
wire n_2715;
wire n_1035;
wire n_1143;
wire n_2665;
wire n_2070;
wire n_2136;
wire n_426;
wire n_433;
wire n_2771;
wire n_1090;
wire n_2403;
wire n_1367;
wire n_2044;
wire n_928;
wire n_1153;
wire n_465;
wire n_825;
wire n_1103;
wire n_732;
wire n_2619;
wire n_1565;
wire n_1192;
wire n_894;
wire n_1380;
wire n_1624;
wire n_1801;
wire n_1291;
wire n_562;
wire n_2020;
wire n_748;
wire n_2310;
wire n_510;
wire n_1045;
wire n_1160;
wire n_1882;
wire n_1976;
wire n_1023;
wire n_2711;
wire n_1881;
wire n_2635;
wire n_988;
wire n_914;
wire n_689;
wire n_1116;
wire n_1958;
wire n_2747;
wire n_467;
wire n_1511;
wire n_2177;
wire n_2713;
wire n_1422;
wire n_2766;
wire n_1965;
wire n_644;
wire n_1197;
wire n_2613;
wire n_497;
wire n_1165;
wire n_1641;
wire n_538;
wire n_1517;
wire n_2036;
wire n_576;
wire n_843;
wire n_511;
wire n_2647;
wire n_455;
wire n_429;
wire n_588;
wire n_638;
wire n_2003;
wire n_2533;
wire n_2210;
wire n_1307;
wire n_1128;
wire n_2053;
wire n_1671;
wire n_1417;
wire n_1048;
wire n_2343;
wire n_775;
wire n_667;
wire n_2419;
wire n_1049;
wire n_2330;
wire n_869;
wire n_846;
wire n_1398;
wire n_1921;
wire n_2777;
wire n_2450;
wire n_2411;
wire n_2234;
wire n_1341;
wire n_1356;
wire n_2309;
wire n_1504;
wire n_1955;
wire n_2110;
wire n_2431;
wire n_1773;
wire n_1440;
wire n_2666;
wire n_1370;
wire n_1603;
wire n_728;
wire n_2401;
wire n_715;
wire n_889;
wire n_1549;
wire n_1066;
wire n_2588;
wire n_2331;
wire n_935;
wire n_2478;
wire n_685;
wire n_911;
wire n_2658;
wire n_623;
wire n_2608;
wire n_1712;
wire n_1403;
wire n_1534;
wire n_453;
wire n_1065;
wire n_1948;
wire n_2767;
wire n_810;
wire n_1959;
wire n_1290;
wire n_617;
wire n_2396;
wire n_543;
wire n_1362;
wire n_1559;
wire n_2121;
wire n_2692;
wire n_601;
wire n_683;
wire n_565;
wire n_628;
wire n_1300;
wire n_1960;
wire n_2068;
wire n_743;
wire n_1194;
wire n_1647;
wire n_1546;
wire n_1420;
wire n_2553;
wire n_2645;
wire n_907;
wire n_2749;
wire n_1454;
wire n_2592;
wire n_660;
wire n_464;
wire n_2459;
wire n_962;
wire n_941;
wire n_1210;
wire n_847;
wire n_747;
wire n_1622;
wire n_1135;
wire n_2566;
wire n_2751;
wire n_1968;
wire n_918;
wire n_1885;
wire n_639;
wire n_452;
wire n_673;
wire n_2196;
wire n_1038;
wire n_2371;
wire n_1978;
wire n_571;
wire n_1521;
wire n_1694;
wire n_1940;
wire n_593;
wire n_1695;
wire n_2560;
wire n_1164;
wire n_2313;
wire n_609;
wire n_1193;
wire n_1345;
wire n_613;
wire n_1022;
wire n_1336;
wire n_1033;
wire n_1774;
wire n_519;
wire n_2609;
wire n_2561;
wire n_1166;
wire n_1056;
wire n_2007;
wire n_526;
wire n_1994;
wire n_1767;
wire n_1040;
wire n_674;
wire n_1158;
wire n_1973;
wire n_1444;
wire n_1803;
wire n_820;
wire n_1749;
wire n_1653;
wire n_872;
wire n_2303;
wire n_2669;
wire n_1157;
wire n_1584;
wire n_848;
wire n_1664;
wire n_629;
wire n_1739;
wire n_2642;
wire n_1814;
wire n_532;
wire n_2154;
wire n_2441;
wire n_2236;
wire n_1789;
wire n_763;
wire n_1986;
wire n_2174;
wire n_2688;
wire n_540;
wire n_692;
wire n_2624;
wire n_2054;
wire n_1857;
wire n_2315;
wire n_984;
wire n_1687;
wire n_2073;
wire n_2150;
wire n_1552;
wire n_750;
wire n_834;
wire n_1612;
wire n_2498;
wire n_800;
wire n_2638;
wire n_2046;
wire n_1816;
wire n_1910;
wire n_1756;
wire n_1606;
wire n_2189;
wire n_621;
wire n_2648;
wire n_1587;
wire n_2093;
wire n_2340;
wire n_2018;
wire n_2672;
wire n_1772;
wire n_2444;
wire n_2602;
wire n_1014;
wire n_724;
wire n_2204;
wire n_1427;
wire n_1481;
wire n_2040;
wire n_493;
wire n_1311;
wire n_2199;
wire n_1956;
wire n_1589;
wire n_2151;
wire n_1100;
wire n_585;
wire n_875;
wire n_1617;
wire n_2455;
wire n_827;
wire n_2600;
wire n_2231;
wire n_697;
wire n_622;
wire n_1626;
wire n_1962;
wire n_1335;
wire n_1715;
wire n_2305;
wire n_880;
wire n_793;
wire n_2114;
wire n_1175;
wire n_2289;
wire n_2530;
wire n_2299;
wire n_751;
wire n_1027;
wire n_1070;
wire n_2406;
wire n_1621;
wire n_739;
wire n_1485;
wire n_1028;
wire n_1221;
wire n_530;
wire n_1785;
wire n_792;
wire n_1262;
wire n_1942;
wire n_2180;
wire n_580;
wire n_1579;
wire n_494;
wire n_2181;
wire n_434;
wire n_2014;
wire n_975;
wire n_1645;
wire n_923;
wire n_1381;
wire n_1124;
wire n_1494;
wire n_1893;
wire n_932;
wire n_1183;
wire n_1326;
wire n_2276;
wire n_1805;
wire n_2282;
wire n_981;
wire n_2141;
wire n_1758;
wire n_1110;
wire n_2503;
wire n_2270;
wire n_2443;
wire n_2465;
wire n_1407;
wire n_1204;
wire n_1554;
wire n_994;
wire n_2428;
wire n_2586;
wire n_1360;
wire n_973;
wire n_972;
wire n_2251;
wire n_856;
wire n_2572;
wire n_1248;
wire n_1176;
wire n_1564;
wire n_2010;
wire n_1054;
wire n_508;
wire n_1679;
wire n_2126;
wire n_1952;
wire n_2425;
wire n_2394;
wire n_1858;
wire n_1678;
wire n_2589;
wire n_1482;
wire n_2356;
wire n_1361;
wire n_1601;
wire n_1057;
wire n_2487;
wire n_1834;
wire n_978;
wire n_1011;
wire n_1520;
wire n_2534;
wire n_2488;
wire n_1509;
wire n_828;
wire n_1411;
wire n_1359;
wire n_558;
wire n_1721;
wire n_2564;
wire n_2591;
wire n_653;
wire n_1445;
wire n_1317;
wire n_2050;
wire n_2197;
wire n_783;
wire n_2550;
wire n_556;
wire n_1127;
wire n_1536;
wire n_1471;
wire n_2385;
wire n_2387;
wire n_1008;
wire n_581;
wire n_1024;
wire n_830;
wire n_2291;
wire n_1980;
wire n_2518;
wire n_987;
wire n_936;
wire n_2510;
wire n_1620;
wire n_2501;
wire n_2542;
wire n_1385;
wire n_1525;
wire n_1998;
wire n_2165;
wire n_2675;
wire n_541;
wire n_499;
wire n_2604;
wire n_1775;
wire n_788;
wire n_908;
wire n_2639;
wire n_1036;
wire n_2169;
wire n_2603;
wire n_1270;
wire n_1167;
wire n_1272;
wire n_549;
wire n_2630;
wire n_591;
wire n_969;
wire n_2028;
wire n_919;
wire n_1663;
wire n_2092;
wire n_2175;
wire n_1625;
wire n_2086;
wire n_2773;
wire n_1926;
wire n_2402;
wire n_1458;
wire n_679;
wire n_1630;
wire n_663;
wire n_1720;
wire n_2409;
wire n_443;
wire n_2176;
wire n_1412;
wire n_1738;
wire n_1550;
wire n_528;
wire n_1358;
wire n_1200;
wire n_826;
wire n_2453;
wire n_2344;
wire n_1922;
wire n_1735;
wire n_1788;
wire n_940;
wire n_2392;
wire n_1537;
wire n_2138;
wire n_2065;
wire n_2543;
wire n_2321;
wire n_1077;
wire n_2597;
wire n_607;
wire n_956;
wire n_445;
wire n_1930;
wire n_1809;
wire n_765;
wire n_2787;
wire n_1843;
wire n_1904;
wire n_2000;
wire n_1268;
wire n_2676;
wire n_2758;
wire n_2395;
wire n_917;
wire n_2723;
wire n_1271;
wire n_2096;
wire n_2440;
wire n_2556;
wire n_2186;
wire n_2215;
wire n_1530;
wire n_2770;
wire n_631;
wire n_1170;
wire n_2724;
wire n_2258;
wire n_1261;
wire n_2471;
wire n_702;
wire n_857;
wire n_898;
wire n_968;
wire n_1067;
wire n_1323;
wire n_1235;
wire n_2584;
wire n_2375;
wire n_1462;
wire n_2012;
wire n_1937;
wire n_1064;
wire n_633;
wire n_900;
wire n_1446;
wire n_1282;
wire n_1701;
wire n_1093;
wire n_1551;
wire n_2039;
wire n_1755;
wire n_1285;
wire n_733;
wire n_761;
wire n_2212;
wire n_731;
wire n_1813;
wire n_2268;
wire n_1452;
wire n_1573;
wire n_2734;
wire n_668;
wire n_2569;
wire n_758;
wire n_2252;
wire n_2111;
wire n_2420;
wire n_1996;
wire n_1106;
wire n_2009;
wire n_784;
wire n_648;
wire n_816;
wire n_1322;
wire n_2583;
wire n_1473;
wire n_835;
wire n_446;
wire n_1076;
wire n_2024;
wire n_1348;
wire n_2651;
wire n_753;
wire n_2445;
wire n_2733;
wire n_1770;
wire n_701;
wire n_1003;
wire n_2469;
wire n_1125;
wire n_2103;
wire n_2358;
wire n_1710;
wire n_1865;
wire n_2522;
wire n_2641;
wire n_2463;
wire n_1344;
wire n_2355;
wire n_1390;
wire n_2580;
wire n_2699;
wire n_485;
wire n_1792;
wire n_504;
wire n_2062;
wire n_483;
wire n_435;
wire n_1141;
wire n_1629;
wire n_1640;
wire n_822;
wire n_1094;
wire n_840;
wire n_1459;
wire n_2153;
wire n_2324;
wire n_1510;
wire n_2710;
wire n_2505;
wire n_2139;
wire n_1099;
wire n_839;
wire n_1754;
wire n_759;
wire n_567;
wire n_2397;
wire n_2521;
wire n_1727;
wire n_2740;
wire n_2235;
wire n_1991;
wire n_1575;
wire n_2721;
wire n_1848;
wire n_1892;
wire n_1172;
wire n_2615;
wire n_614;
wire n_2775;
wire n_1212;
wire n_831;
wire n_778;
wire n_1619;
wire n_2351;
wire n_2260;
wire n_550;
wire n_1315;
wire n_1660;
wire n_1902;
wire n_997;
wire n_635;
wire n_2206;
wire n_2784;
wire n_2541;
wire n_694;
wire n_1643;
wire n_1320;
wire n_1113;
wire n_2347;
wire n_1152;
wire n_2657;
wire n_2447;
wire n_2034;
wire n_1845;
wire n_2538;
wire n_1934;
wire n_2101;
wire n_2577;
wire n_921;
wire n_2362;
wire n_1615;
wire n_1236;
wire n_2104;
wire n_1265;
wire n_1576;
wire n_2105;
wire n_1470;
wire n_1806;
wire n_1533;
wire n_671;
wire n_2372;
wire n_2552;
wire n_1409;
wire n_1588;
wire n_1148;
wire n_1684;
wire n_1673;
wire n_2422;
wire n_2704;
wire n_1334;
wire n_654;
wire n_2290;
wire n_2088;
wire n_1275;
wire n_488;
wire n_904;
wire n_505;
wire n_2005;
wire n_2048;
wire n_1696;
wire n_498;
wire n_1875;
wire n_1059;
wire n_684;
wire n_2429;
wire n_2108;
wire n_2736;
wire n_1039;
wire n_2246;
wire n_539;
wire n_1150;
wire n_977;
wire n_449;
wire n_2339;
wire n_1628;
wire n_1289;
wire n_1831;
wire n_2532;
wire n_2191;
wire n_1497;
wire n_1866;
wire n_2472;
wire n_2664;
wire n_2705;
wire n_2056;
wire n_459;
wire n_1136;
wire n_2515;
wire n_1782;
wire n_458;
wire n_1190;
wire n_1600;
wire n_1144;
wire n_838;
wire n_1558;
wire n_1941;
wire n_1316;
wire n_2519;
wire n_950;
wire n_1017;
wire n_711;
wire n_734;
wire n_1915;
wire n_2360;
wire n_723;
wire n_1393;
wire n_2240;
wire n_658;
wire n_630;
wire n_1369;
wire n_1781;
wire n_709;
wire n_2544;
wire n_809;
wire n_2085;
wire n_2432;
wire n_1686;
wire n_1964;
wire n_881;
wire n_1019;
wire n_1477;
wire n_1777;
wire n_2188;
wire n_1982;
wire n_2097;
wire n_662;
wire n_641;
wire n_2430;
wire n_2504;
wire n_910;
wire n_741;
wire n_1410;
wire n_939;
wire n_2297;
wire n_1114;
wire n_1325;
wire n_1742;
wire n_708;
wire n_1223;
wire n_2545;
wire n_2513;
wire n_1768;
wire n_2193;
wire n_2369;
wire n_572;
wire n_1199;
wire n_865;
wire n_1273;
wire n_1983;
wire n_1041;
wire n_2451;
wire n_2115;
wire n_993;
wire n_1862;
wire n_948;
wire n_2017;
wire n_922;
wire n_1004;
wire n_1810;
wire n_448;
wire n_2587;
wire n_1347;
wire n_860;
wire n_1043;
wire n_450;
wire n_1923;
wire n_2670;
wire n_1764;
wire n_2674;
wire n_896;
wire n_1737;
wire n_1479;
wire n_1613;
wire n_2644;
wire n_902;
wire n_1031;
wire n_1723;
wire n_1638;
wire n_853;
wire n_716;
wire n_1571;
wire n_1698;
wire n_1337;
wire n_2148;
wire n_1946;
wire n_774;
wire n_933;
wire n_1779;
wire n_2562;
wire n_596;
wire n_954;
wire n_2051;
wire n_1168;
wire n_1821;
wire n_1310;
wire n_656;
wire n_492;
wire n_574;
wire n_2673;
wire n_664;
wire n_1591;
wire n_2585;
wire n_1229;
wire n_1683;
wire n_2582;
wire n_2548;
wire n_1896;
wire n_2164;
wire n_1732;
wire n_2381;
wire n_2744;
wire n_1967;
wire n_2384;
wire n_2678;
wire n_2179;
wire n_1280;
wire n_544;
wire n_1516;
wire n_1186;
wire n_1705;
wire n_599;
wire n_768;
wire n_1091;
wire n_2052;
wire n_2485;
wire n_537;
wire n_1063;
wire n_991;
wire n_2205;
wire n_2183;
wire n_2275;
wire n_2563;
wire n_1724;
wire n_1670;
wire n_1799;
wire n_1707;
wire n_2080;
wire n_2058;
wire n_1126;
wire n_2761;
wire n_2357;
wire n_2029;
wire n_1846;
wire n_1912;
wire n_938;
wire n_1891;
wire n_1328;
wire n_895;
wire n_1639;
wire n_583;
wire n_2209;
wire n_2421;
wire n_1302;
wire n_1000;
wire n_626;
wire n_1581;
wire n_1928;
wire n_946;
wire n_757;
wire n_2047;
wire n_1655;
wire n_1818;
wire n_1146;
wire n_2792;
wire n_1634;
wire n_2596;
wire n_1203;
wire n_998;
wire n_1699;
wire n_1598;
wire n_2269;
wire n_472;
wire n_937;
wire n_1474;
wire n_2081;
wire n_2536;
wire n_2524;
wire n_1583;
wire n_1604;
wire n_1631;
wire n_1702;
wire n_1794;
wire n_1375;
wire n_1232;
wire n_996;
wire n_1211;
wire n_1368;
wire n_963;
wire n_1264;
wire n_1082;
wire n_1725;
wire n_496;
wire n_2318;
wire n_1827;
wire n_866;
wire n_925;
wire n_1752;
wire n_1313;
wire n_1001;
wire n_1722;
wire n_2361;
wire n_1115;
wire n_2229;
wire n_1339;
wire n_1002;
wire n_1644;
wire n_1051;
wire n_2551;
wire n_1102;
wire n_719;
wire n_2255;
wire n_1252;
wire n_2239;
wire n_1129;
wire n_1464;
wire n_1296;
wire n_773;
wire n_2316;
wire n_2464;
wire n_1010;
wire n_882;
wire n_2706;
wire n_2304;
wire n_1249;
wire n_803;
wire n_1871;
wire n_2514;
wire n_718;
wire n_1434;
wire n_1905;
wire n_1569;
wire n_2573;
wire n_548;
wire n_2336;
wire n_523;
wire n_1662;
wire n_457;
wire n_1299;
wire n_1870;
wire n_2063;
wire n_1925;
wire n_782;
wire n_431;
wire n_2654;
wire n_2491;
wire n_1861;
wire n_2079;
wire n_1228;
wire n_2319;
wire n_2152;
wire n_2517;
wire n_1931;
wire n_1244;
wire n_1796;
wire n_484;
wire n_2259;
wire n_849;
wire n_2095;
wire n_2719;
wire n_2738;
wire n_1820;
wire n_2590;
wire n_1251;
wire n_1989;
wire n_447;
wire n_2208;
wire n_1421;
wire n_2423;
wire n_2689;
wire n_2778;
wire n_1762;
wire n_1233;
wire n_1808;
wire n_1574;
wire n_1672;
wire n_2228;
wire n_1635;
wire n_1704;
wire n_893;
wire n_1582;
wire n_841;
wire n_2479;
wire n_886;
wire n_1069;
wire n_1981;
wire n_2037;
wire n_1308;
wire n_573;
wire n_796;
wire n_531;
wire n_2345;
wire n_1730;
wire n_1374;
wire n_1451;
wire n_2089;
wire n_1487;
wire n_675;

BUFx6f_ASAP7_75t_L g426 ( 
.A(n_388),
.Y(n_426)
);

CKINVDCx5p33_ASAP7_75t_R g427 ( 
.A(n_99),
.Y(n_427)
);

INVx1_ASAP7_75t_L g428 ( 
.A(n_265),
.Y(n_428)
);

CKINVDCx5p33_ASAP7_75t_R g429 ( 
.A(n_298),
.Y(n_429)
);

CKINVDCx20_ASAP7_75t_R g430 ( 
.A(n_368),
.Y(n_430)
);

CKINVDCx20_ASAP7_75t_R g431 ( 
.A(n_301),
.Y(n_431)
);

INVx1_ASAP7_75t_L g432 ( 
.A(n_371),
.Y(n_432)
);

CKINVDCx20_ASAP7_75t_R g433 ( 
.A(n_113),
.Y(n_433)
);

CKINVDCx5p33_ASAP7_75t_R g434 ( 
.A(n_153),
.Y(n_434)
);

BUFx2_ASAP7_75t_L g435 ( 
.A(n_133),
.Y(n_435)
);

CKINVDCx5p33_ASAP7_75t_R g436 ( 
.A(n_211),
.Y(n_436)
);

CKINVDCx5p33_ASAP7_75t_R g437 ( 
.A(n_81),
.Y(n_437)
);

CKINVDCx20_ASAP7_75t_R g438 ( 
.A(n_243),
.Y(n_438)
);

INVx1_ASAP7_75t_L g439 ( 
.A(n_167),
.Y(n_439)
);

CKINVDCx5p33_ASAP7_75t_R g440 ( 
.A(n_259),
.Y(n_440)
);

CKINVDCx5p33_ASAP7_75t_R g441 ( 
.A(n_204),
.Y(n_441)
);

CKINVDCx20_ASAP7_75t_R g442 ( 
.A(n_131),
.Y(n_442)
);

INVx1_ASAP7_75t_L g443 ( 
.A(n_334),
.Y(n_443)
);

CKINVDCx5p33_ASAP7_75t_R g444 ( 
.A(n_416),
.Y(n_444)
);

CKINVDCx5p33_ASAP7_75t_R g445 ( 
.A(n_133),
.Y(n_445)
);

INVx1_ASAP7_75t_L g446 ( 
.A(n_156),
.Y(n_446)
);

CKINVDCx5p33_ASAP7_75t_R g447 ( 
.A(n_160),
.Y(n_447)
);

BUFx10_ASAP7_75t_L g448 ( 
.A(n_325),
.Y(n_448)
);

CKINVDCx5p33_ASAP7_75t_R g449 ( 
.A(n_29),
.Y(n_449)
);

INVx1_ASAP7_75t_L g450 ( 
.A(n_315),
.Y(n_450)
);

CKINVDCx20_ASAP7_75t_R g451 ( 
.A(n_164),
.Y(n_451)
);

INVx1_ASAP7_75t_L g452 ( 
.A(n_65),
.Y(n_452)
);

INVx1_ASAP7_75t_L g453 ( 
.A(n_172),
.Y(n_453)
);

CKINVDCx5p33_ASAP7_75t_R g454 ( 
.A(n_278),
.Y(n_454)
);

CKINVDCx5p33_ASAP7_75t_R g455 ( 
.A(n_423),
.Y(n_455)
);

CKINVDCx5p33_ASAP7_75t_R g456 ( 
.A(n_287),
.Y(n_456)
);

BUFx3_ASAP7_75t_L g457 ( 
.A(n_60),
.Y(n_457)
);

CKINVDCx16_ASAP7_75t_R g458 ( 
.A(n_367),
.Y(n_458)
);

CKINVDCx5p33_ASAP7_75t_R g459 ( 
.A(n_46),
.Y(n_459)
);

INVx1_ASAP7_75t_L g460 ( 
.A(n_414),
.Y(n_460)
);

CKINVDCx5p33_ASAP7_75t_R g461 ( 
.A(n_383),
.Y(n_461)
);

INVx2_ASAP7_75t_L g462 ( 
.A(n_422),
.Y(n_462)
);

CKINVDCx20_ASAP7_75t_R g463 ( 
.A(n_62),
.Y(n_463)
);

BUFx3_ASAP7_75t_L g464 ( 
.A(n_125),
.Y(n_464)
);

CKINVDCx5p33_ASAP7_75t_R g465 ( 
.A(n_401),
.Y(n_465)
);

INVx1_ASAP7_75t_L g466 ( 
.A(n_93),
.Y(n_466)
);

INVx1_ASAP7_75t_L g467 ( 
.A(n_411),
.Y(n_467)
);

INVx1_ASAP7_75t_L g468 ( 
.A(n_282),
.Y(n_468)
);

INVx1_ASAP7_75t_L g469 ( 
.A(n_373),
.Y(n_469)
);

CKINVDCx5p33_ASAP7_75t_R g470 ( 
.A(n_74),
.Y(n_470)
);

INVx2_ASAP7_75t_SL g471 ( 
.A(n_391),
.Y(n_471)
);

INVx1_ASAP7_75t_L g472 ( 
.A(n_290),
.Y(n_472)
);

CKINVDCx5p33_ASAP7_75t_R g473 ( 
.A(n_52),
.Y(n_473)
);

INVx1_ASAP7_75t_L g474 ( 
.A(n_275),
.Y(n_474)
);

CKINVDCx5p33_ASAP7_75t_R g475 ( 
.A(n_396),
.Y(n_475)
);

CKINVDCx5p33_ASAP7_75t_R g476 ( 
.A(n_303),
.Y(n_476)
);

INVx2_ASAP7_75t_SL g477 ( 
.A(n_205),
.Y(n_477)
);

CKINVDCx5p33_ASAP7_75t_R g478 ( 
.A(n_27),
.Y(n_478)
);

INVx1_ASAP7_75t_L g479 ( 
.A(n_249),
.Y(n_479)
);

CKINVDCx5p33_ASAP7_75t_R g480 ( 
.A(n_262),
.Y(n_480)
);

CKINVDCx5p33_ASAP7_75t_R g481 ( 
.A(n_333),
.Y(n_481)
);

INVx1_ASAP7_75t_L g482 ( 
.A(n_126),
.Y(n_482)
);

CKINVDCx5p33_ASAP7_75t_R g483 ( 
.A(n_217),
.Y(n_483)
);

CKINVDCx20_ASAP7_75t_R g484 ( 
.A(n_100),
.Y(n_484)
);

CKINVDCx5p33_ASAP7_75t_R g485 ( 
.A(n_179),
.Y(n_485)
);

CKINVDCx5p33_ASAP7_75t_R g486 ( 
.A(n_51),
.Y(n_486)
);

CKINVDCx5p33_ASAP7_75t_R g487 ( 
.A(n_407),
.Y(n_487)
);

CKINVDCx5p33_ASAP7_75t_R g488 ( 
.A(n_161),
.Y(n_488)
);

INVx1_ASAP7_75t_L g489 ( 
.A(n_134),
.Y(n_489)
);

INVx1_ASAP7_75t_L g490 ( 
.A(n_369),
.Y(n_490)
);

CKINVDCx5p33_ASAP7_75t_R g491 ( 
.A(n_223),
.Y(n_491)
);

CKINVDCx5p33_ASAP7_75t_R g492 ( 
.A(n_238),
.Y(n_492)
);

INVx1_ASAP7_75t_L g493 ( 
.A(n_350),
.Y(n_493)
);

CKINVDCx5p33_ASAP7_75t_R g494 ( 
.A(n_295),
.Y(n_494)
);

CKINVDCx5p33_ASAP7_75t_R g495 ( 
.A(n_378),
.Y(n_495)
);

CKINVDCx5p33_ASAP7_75t_R g496 ( 
.A(n_323),
.Y(n_496)
);

INVx2_ASAP7_75t_L g497 ( 
.A(n_225),
.Y(n_497)
);

CKINVDCx5p33_ASAP7_75t_R g498 ( 
.A(n_145),
.Y(n_498)
);

BUFx3_ASAP7_75t_L g499 ( 
.A(n_185),
.Y(n_499)
);

INVxp67_ASAP7_75t_L g500 ( 
.A(n_178),
.Y(n_500)
);

BUFx3_ASAP7_75t_L g501 ( 
.A(n_24),
.Y(n_501)
);

INVx1_ASAP7_75t_L g502 ( 
.A(n_421),
.Y(n_502)
);

CKINVDCx5p33_ASAP7_75t_R g503 ( 
.A(n_342),
.Y(n_503)
);

INVx2_ASAP7_75t_SL g504 ( 
.A(n_320),
.Y(n_504)
);

INVx1_ASAP7_75t_L g505 ( 
.A(n_255),
.Y(n_505)
);

CKINVDCx5p33_ASAP7_75t_R g506 ( 
.A(n_45),
.Y(n_506)
);

INVx2_ASAP7_75t_L g507 ( 
.A(n_180),
.Y(n_507)
);

CKINVDCx5p33_ASAP7_75t_R g508 ( 
.A(n_181),
.Y(n_508)
);

CKINVDCx5p33_ASAP7_75t_R g509 ( 
.A(n_283),
.Y(n_509)
);

CKINVDCx5p33_ASAP7_75t_R g510 ( 
.A(n_136),
.Y(n_510)
);

CKINVDCx5p33_ASAP7_75t_R g511 ( 
.A(n_44),
.Y(n_511)
);

CKINVDCx5p33_ASAP7_75t_R g512 ( 
.A(n_349),
.Y(n_512)
);

INVx1_ASAP7_75t_L g513 ( 
.A(n_267),
.Y(n_513)
);

CKINVDCx5p33_ASAP7_75t_R g514 ( 
.A(n_176),
.Y(n_514)
);

INVx1_ASAP7_75t_L g515 ( 
.A(n_80),
.Y(n_515)
);

CKINVDCx14_ASAP7_75t_R g516 ( 
.A(n_341),
.Y(n_516)
);

BUFx3_ASAP7_75t_L g517 ( 
.A(n_165),
.Y(n_517)
);

CKINVDCx5p33_ASAP7_75t_R g518 ( 
.A(n_239),
.Y(n_518)
);

CKINVDCx5p33_ASAP7_75t_R g519 ( 
.A(n_218),
.Y(n_519)
);

INVx1_ASAP7_75t_L g520 ( 
.A(n_190),
.Y(n_520)
);

CKINVDCx5p33_ASAP7_75t_R g521 ( 
.A(n_345),
.Y(n_521)
);

CKINVDCx5p33_ASAP7_75t_R g522 ( 
.A(n_24),
.Y(n_522)
);

CKINVDCx5p33_ASAP7_75t_R g523 ( 
.A(n_269),
.Y(n_523)
);

CKINVDCx5p33_ASAP7_75t_R g524 ( 
.A(n_257),
.Y(n_524)
);

INVx1_ASAP7_75t_L g525 ( 
.A(n_173),
.Y(n_525)
);

INVx1_ASAP7_75t_L g526 ( 
.A(n_370),
.Y(n_526)
);

CKINVDCx20_ASAP7_75t_R g527 ( 
.A(n_35),
.Y(n_527)
);

CKINVDCx5p33_ASAP7_75t_R g528 ( 
.A(n_119),
.Y(n_528)
);

CKINVDCx5p33_ASAP7_75t_R g529 ( 
.A(n_284),
.Y(n_529)
);

INVx1_ASAP7_75t_L g530 ( 
.A(n_166),
.Y(n_530)
);

INVx1_ASAP7_75t_L g531 ( 
.A(n_288),
.Y(n_531)
);

CKINVDCx5p33_ASAP7_75t_R g532 ( 
.A(n_286),
.Y(n_532)
);

CKINVDCx16_ASAP7_75t_R g533 ( 
.A(n_386),
.Y(n_533)
);

BUFx2_ASAP7_75t_L g534 ( 
.A(n_372),
.Y(n_534)
);

CKINVDCx20_ASAP7_75t_R g535 ( 
.A(n_235),
.Y(n_535)
);

INVx1_ASAP7_75t_L g536 ( 
.A(n_353),
.Y(n_536)
);

CKINVDCx20_ASAP7_75t_R g537 ( 
.A(n_170),
.Y(n_537)
);

INVx1_ASAP7_75t_L g538 ( 
.A(n_335),
.Y(n_538)
);

INVx1_ASAP7_75t_L g539 ( 
.A(n_5),
.Y(n_539)
);

BUFx2_ASAP7_75t_L g540 ( 
.A(n_0),
.Y(n_540)
);

CKINVDCx20_ASAP7_75t_R g541 ( 
.A(n_310),
.Y(n_541)
);

CKINVDCx20_ASAP7_75t_R g542 ( 
.A(n_250),
.Y(n_542)
);

CKINVDCx5p33_ASAP7_75t_R g543 ( 
.A(n_65),
.Y(n_543)
);

CKINVDCx5p33_ASAP7_75t_R g544 ( 
.A(n_385),
.Y(n_544)
);

CKINVDCx5p33_ASAP7_75t_R g545 ( 
.A(n_155),
.Y(n_545)
);

INVx2_ASAP7_75t_L g546 ( 
.A(n_57),
.Y(n_546)
);

INVx1_ASAP7_75t_L g547 ( 
.A(n_242),
.Y(n_547)
);

INVx1_ASAP7_75t_L g548 ( 
.A(n_42),
.Y(n_548)
);

CKINVDCx5p33_ASAP7_75t_R g549 ( 
.A(n_256),
.Y(n_549)
);

CKINVDCx5p33_ASAP7_75t_R g550 ( 
.A(n_175),
.Y(n_550)
);

CKINVDCx5p33_ASAP7_75t_R g551 ( 
.A(n_404),
.Y(n_551)
);

CKINVDCx5p33_ASAP7_75t_R g552 ( 
.A(n_299),
.Y(n_552)
);

INVx1_ASAP7_75t_L g553 ( 
.A(n_208),
.Y(n_553)
);

BUFx3_ASAP7_75t_L g554 ( 
.A(n_354),
.Y(n_554)
);

INVx1_ASAP7_75t_L g555 ( 
.A(n_68),
.Y(n_555)
);

CKINVDCx5p33_ASAP7_75t_R g556 ( 
.A(n_158),
.Y(n_556)
);

INVx1_ASAP7_75t_L g557 ( 
.A(n_192),
.Y(n_557)
);

INVxp67_ASAP7_75t_SL g558 ( 
.A(n_330),
.Y(n_558)
);

INVx1_ASAP7_75t_L g559 ( 
.A(n_152),
.Y(n_559)
);

INVx1_ASAP7_75t_L g560 ( 
.A(n_338),
.Y(n_560)
);

CKINVDCx5p33_ASAP7_75t_R g561 ( 
.A(n_8),
.Y(n_561)
);

CKINVDCx20_ASAP7_75t_R g562 ( 
.A(n_48),
.Y(n_562)
);

CKINVDCx5p33_ASAP7_75t_R g563 ( 
.A(n_258),
.Y(n_563)
);

INVx1_ASAP7_75t_L g564 ( 
.A(n_376),
.Y(n_564)
);

INVx1_ASAP7_75t_L g565 ( 
.A(n_403),
.Y(n_565)
);

INVx3_ASAP7_75t_L g566 ( 
.A(n_121),
.Y(n_566)
);

INVx1_ASAP7_75t_L g567 ( 
.A(n_237),
.Y(n_567)
);

HB1xp67_ASAP7_75t_L g568 ( 
.A(n_232),
.Y(n_568)
);

CKINVDCx5p33_ASAP7_75t_R g569 ( 
.A(n_60),
.Y(n_569)
);

INVx1_ASAP7_75t_L g570 ( 
.A(n_181),
.Y(n_570)
);

INVxp67_ASAP7_75t_L g571 ( 
.A(n_88),
.Y(n_571)
);

CKINVDCx20_ASAP7_75t_R g572 ( 
.A(n_397),
.Y(n_572)
);

INVx1_ASAP7_75t_L g573 ( 
.A(n_38),
.Y(n_573)
);

INVx2_ASAP7_75t_L g574 ( 
.A(n_187),
.Y(n_574)
);

CKINVDCx5p33_ASAP7_75t_R g575 ( 
.A(n_99),
.Y(n_575)
);

CKINVDCx5p33_ASAP7_75t_R g576 ( 
.A(n_11),
.Y(n_576)
);

CKINVDCx5p33_ASAP7_75t_R g577 ( 
.A(n_253),
.Y(n_577)
);

CKINVDCx5p33_ASAP7_75t_R g578 ( 
.A(n_100),
.Y(n_578)
);

INVx1_ASAP7_75t_SL g579 ( 
.A(n_49),
.Y(n_579)
);

CKINVDCx5p33_ASAP7_75t_R g580 ( 
.A(n_351),
.Y(n_580)
);

BUFx10_ASAP7_75t_L g581 ( 
.A(n_218),
.Y(n_581)
);

BUFx6f_ASAP7_75t_L g582 ( 
.A(n_42),
.Y(n_582)
);

CKINVDCx5p33_ASAP7_75t_R g583 ( 
.A(n_402),
.Y(n_583)
);

CKINVDCx5p33_ASAP7_75t_R g584 ( 
.A(n_174),
.Y(n_584)
);

CKINVDCx5p33_ASAP7_75t_R g585 ( 
.A(n_21),
.Y(n_585)
);

CKINVDCx5p33_ASAP7_75t_R g586 ( 
.A(n_294),
.Y(n_586)
);

CKINVDCx5p33_ASAP7_75t_R g587 ( 
.A(n_420),
.Y(n_587)
);

INVx1_ASAP7_75t_SL g588 ( 
.A(n_313),
.Y(n_588)
);

CKINVDCx5p33_ASAP7_75t_R g589 ( 
.A(n_63),
.Y(n_589)
);

CKINVDCx5p33_ASAP7_75t_R g590 ( 
.A(n_227),
.Y(n_590)
);

BUFx3_ASAP7_75t_L g591 ( 
.A(n_115),
.Y(n_591)
);

CKINVDCx5p33_ASAP7_75t_R g592 ( 
.A(n_32),
.Y(n_592)
);

INVx1_ASAP7_75t_L g593 ( 
.A(n_410),
.Y(n_593)
);

CKINVDCx5p33_ASAP7_75t_R g594 ( 
.A(n_336),
.Y(n_594)
);

CKINVDCx5p33_ASAP7_75t_R g595 ( 
.A(n_52),
.Y(n_595)
);

CKINVDCx20_ASAP7_75t_R g596 ( 
.A(n_64),
.Y(n_596)
);

CKINVDCx5p33_ASAP7_75t_R g597 ( 
.A(n_240),
.Y(n_597)
);

CKINVDCx5p33_ASAP7_75t_R g598 ( 
.A(n_360),
.Y(n_598)
);

CKINVDCx5p33_ASAP7_75t_R g599 ( 
.A(n_130),
.Y(n_599)
);

CKINVDCx5p33_ASAP7_75t_R g600 ( 
.A(n_210),
.Y(n_600)
);

INVx1_ASAP7_75t_L g601 ( 
.A(n_209),
.Y(n_601)
);

CKINVDCx20_ASAP7_75t_R g602 ( 
.A(n_21),
.Y(n_602)
);

CKINVDCx5p33_ASAP7_75t_R g603 ( 
.A(n_405),
.Y(n_603)
);

CKINVDCx5p33_ASAP7_75t_R g604 ( 
.A(n_415),
.Y(n_604)
);

CKINVDCx5p33_ASAP7_75t_R g605 ( 
.A(n_23),
.Y(n_605)
);

CKINVDCx20_ASAP7_75t_R g606 ( 
.A(n_48),
.Y(n_606)
);

CKINVDCx5p33_ASAP7_75t_R g607 ( 
.A(n_96),
.Y(n_607)
);

INVx1_ASAP7_75t_L g608 ( 
.A(n_362),
.Y(n_608)
);

BUFx3_ASAP7_75t_L g609 ( 
.A(n_9),
.Y(n_609)
);

CKINVDCx5p33_ASAP7_75t_R g610 ( 
.A(n_314),
.Y(n_610)
);

BUFx3_ASAP7_75t_L g611 ( 
.A(n_228),
.Y(n_611)
);

CKINVDCx20_ASAP7_75t_R g612 ( 
.A(n_109),
.Y(n_612)
);

CKINVDCx5p33_ASAP7_75t_R g613 ( 
.A(n_297),
.Y(n_613)
);

CKINVDCx5p33_ASAP7_75t_R g614 ( 
.A(n_51),
.Y(n_614)
);

INVx1_ASAP7_75t_L g615 ( 
.A(n_63),
.Y(n_615)
);

INVx1_ASAP7_75t_L g616 ( 
.A(n_154),
.Y(n_616)
);

INVx1_ASAP7_75t_L g617 ( 
.A(n_58),
.Y(n_617)
);

BUFx10_ASAP7_75t_L g618 ( 
.A(n_55),
.Y(n_618)
);

CKINVDCx5p33_ASAP7_75t_R g619 ( 
.A(n_176),
.Y(n_619)
);

CKINVDCx5p33_ASAP7_75t_R g620 ( 
.A(n_153),
.Y(n_620)
);

CKINVDCx5p33_ASAP7_75t_R g621 ( 
.A(n_375),
.Y(n_621)
);

BUFx2_ASAP7_75t_L g622 ( 
.A(n_254),
.Y(n_622)
);

INVx2_ASAP7_75t_L g623 ( 
.A(n_13),
.Y(n_623)
);

CKINVDCx20_ASAP7_75t_R g624 ( 
.A(n_70),
.Y(n_624)
);

INVx1_ASAP7_75t_L g625 ( 
.A(n_56),
.Y(n_625)
);

CKINVDCx20_ASAP7_75t_R g626 ( 
.A(n_102),
.Y(n_626)
);

CKINVDCx5p33_ASAP7_75t_R g627 ( 
.A(n_185),
.Y(n_627)
);

BUFx6f_ASAP7_75t_L g628 ( 
.A(n_387),
.Y(n_628)
);

CKINVDCx5p33_ASAP7_75t_R g629 ( 
.A(n_395),
.Y(n_629)
);

INVx1_ASAP7_75t_L g630 ( 
.A(n_131),
.Y(n_630)
);

CKINVDCx5p33_ASAP7_75t_R g631 ( 
.A(n_101),
.Y(n_631)
);

INVx1_ASAP7_75t_L g632 ( 
.A(n_17),
.Y(n_632)
);

INVx4_ASAP7_75t_R g633 ( 
.A(n_393),
.Y(n_633)
);

INVx1_ASAP7_75t_L g634 ( 
.A(n_276),
.Y(n_634)
);

INVx1_ASAP7_75t_L g635 ( 
.A(n_363),
.Y(n_635)
);

INVx1_ASAP7_75t_L g636 ( 
.A(n_7),
.Y(n_636)
);

BUFx2_ASAP7_75t_L g637 ( 
.A(n_322),
.Y(n_637)
);

INVx1_ASAP7_75t_L g638 ( 
.A(n_4),
.Y(n_638)
);

CKINVDCx5p33_ASAP7_75t_R g639 ( 
.A(n_69),
.Y(n_639)
);

CKINVDCx5p33_ASAP7_75t_R g640 ( 
.A(n_263),
.Y(n_640)
);

INVx1_ASAP7_75t_SL g641 ( 
.A(n_148),
.Y(n_641)
);

BUFx3_ASAP7_75t_L g642 ( 
.A(n_419),
.Y(n_642)
);

INVx1_ASAP7_75t_L g643 ( 
.A(n_152),
.Y(n_643)
);

CKINVDCx5p33_ASAP7_75t_R g644 ( 
.A(n_180),
.Y(n_644)
);

CKINVDCx5p33_ASAP7_75t_R g645 ( 
.A(n_219),
.Y(n_645)
);

CKINVDCx20_ASAP7_75t_R g646 ( 
.A(n_161),
.Y(n_646)
);

INVx1_ASAP7_75t_L g647 ( 
.A(n_168),
.Y(n_647)
);

CKINVDCx5p33_ASAP7_75t_R g648 ( 
.A(n_245),
.Y(n_648)
);

CKINVDCx5p33_ASAP7_75t_R g649 ( 
.A(n_129),
.Y(n_649)
);

CKINVDCx5p33_ASAP7_75t_R g650 ( 
.A(n_69),
.Y(n_650)
);

CKINVDCx5p33_ASAP7_75t_R g651 ( 
.A(n_271),
.Y(n_651)
);

CKINVDCx5p33_ASAP7_75t_R g652 ( 
.A(n_214),
.Y(n_652)
);

CKINVDCx5p33_ASAP7_75t_R g653 ( 
.A(n_268),
.Y(n_653)
);

INVx1_ASAP7_75t_L g654 ( 
.A(n_346),
.Y(n_654)
);

CKINVDCx11_ASAP7_75t_R g655 ( 
.A(n_129),
.Y(n_655)
);

CKINVDCx5p33_ASAP7_75t_R g656 ( 
.A(n_226),
.Y(n_656)
);

CKINVDCx5p33_ASAP7_75t_R g657 ( 
.A(n_399),
.Y(n_657)
);

INVx1_ASAP7_75t_SL g658 ( 
.A(n_135),
.Y(n_658)
);

INVx1_ASAP7_75t_L g659 ( 
.A(n_22),
.Y(n_659)
);

CKINVDCx5p33_ASAP7_75t_R g660 ( 
.A(n_417),
.Y(n_660)
);

INVx2_ASAP7_75t_SL g661 ( 
.A(n_352),
.Y(n_661)
);

CKINVDCx20_ASAP7_75t_R g662 ( 
.A(n_306),
.Y(n_662)
);

INVx1_ASAP7_75t_SL g663 ( 
.A(n_205),
.Y(n_663)
);

CKINVDCx14_ASAP7_75t_R g664 ( 
.A(n_285),
.Y(n_664)
);

CKINVDCx14_ASAP7_75t_R g665 ( 
.A(n_27),
.Y(n_665)
);

CKINVDCx20_ASAP7_75t_R g666 ( 
.A(n_305),
.Y(n_666)
);

CKINVDCx5p33_ASAP7_75t_R g667 ( 
.A(n_337),
.Y(n_667)
);

INVx1_ASAP7_75t_L g668 ( 
.A(n_251),
.Y(n_668)
);

CKINVDCx5p33_ASAP7_75t_R g669 ( 
.A(n_304),
.Y(n_669)
);

INVx1_ASAP7_75t_L g670 ( 
.A(n_412),
.Y(n_670)
);

CKINVDCx5p33_ASAP7_75t_R g671 ( 
.A(n_34),
.Y(n_671)
);

INVx1_ASAP7_75t_L g672 ( 
.A(n_146),
.Y(n_672)
);

CKINVDCx5p33_ASAP7_75t_R g673 ( 
.A(n_379),
.Y(n_673)
);

CKINVDCx5p33_ASAP7_75t_R g674 ( 
.A(n_179),
.Y(n_674)
);

CKINVDCx5p33_ASAP7_75t_R g675 ( 
.A(n_309),
.Y(n_675)
);

INVx1_ASAP7_75t_L g676 ( 
.A(n_277),
.Y(n_676)
);

CKINVDCx5p33_ASAP7_75t_R g677 ( 
.A(n_4),
.Y(n_677)
);

CKINVDCx5p33_ASAP7_75t_R g678 ( 
.A(n_357),
.Y(n_678)
);

INVx1_ASAP7_75t_L g679 ( 
.A(n_29),
.Y(n_679)
);

INVx1_ASAP7_75t_L g680 ( 
.A(n_199),
.Y(n_680)
);

CKINVDCx5p33_ASAP7_75t_R g681 ( 
.A(n_347),
.Y(n_681)
);

CKINVDCx20_ASAP7_75t_R g682 ( 
.A(n_0),
.Y(n_682)
);

CKINVDCx20_ASAP7_75t_R g683 ( 
.A(n_62),
.Y(n_683)
);

INVx1_ASAP7_75t_L g684 ( 
.A(n_28),
.Y(n_684)
);

INVx1_ASAP7_75t_L g685 ( 
.A(n_390),
.Y(n_685)
);

CKINVDCx5p33_ASAP7_75t_R g686 ( 
.A(n_358),
.Y(n_686)
);

INVx2_ASAP7_75t_SL g687 ( 
.A(n_162),
.Y(n_687)
);

CKINVDCx5p33_ASAP7_75t_R g688 ( 
.A(n_102),
.Y(n_688)
);

CKINVDCx5p33_ASAP7_75t_R g689 ( 
.A(n_316),
.Y(n_689)
);

CKINVDCx5p33_ASAP7_75t_R g690 ( 
.A(n_151),
.Y(n_690)
);

INVx1_ASAP7_75t_L g691 ( 
.A(n_85),
.Y(n_691)
);

INVx1_ASAP7_75t_L g692 ( 
.A(n_34),
.Y(n_692)
);

CKINVDCx5p33_ASAP7_75t_R g693 ( 
.A(n_409),
.Y(n_693)
);

CKINVDCx20_ASAP7_75t_R g694 ( 
.A(n_164),
.Y(n_694)
);

CKINVDCx20_ASAP7_75t_R g695 ( 
.A(n_81),
.Y(n_695)
);

CKINVDCx20_ASAP7_75t_R g696 ( 
.A(n_55),
.Y(n_696)
);

INVx1_ASAP7_75t_L g697 ( 
.A(n_273),
.Y(n_697)
);

INVx1_ASAP7_75t_L g698 ( 
.A(n_361),
.Y(n_698)
);

CKINVDCx5p33_ASAP7_75t_R g699 ( 
.A(n_41),
.Y(n_699)
);

INVx1_ASAP7_75t_L g700 ( 
.A(n_406),
.Y(n_700)
);

BUFx3_ASAP7_75t_L g701 ( 
.A(n_326),
.Y(n_701)
);

CKINVDCx20_ASAP7_75t_R g702 ( 
.A(n_365),
.Y(n_702)
);

INVx1_ASAP7_75t_L g703 ( 
.A(n_374),
.Y(n_703)
);

CKINVDCx5p33_ASAP7_75t_R g704 ( 
.A(n_366),
.Y(n_704)
);

CKINVDCx5p33_ASAP7_75t_R g705 ( 
.A(n_45),
.Y(n_705)
);

CKINVDCx5p33_ASAP7_75t_R g706 ( 
.A(n_160),
.Y(n_706)
);

CKINVDCx5p33_ASAP7_75t_R g707 ( 
.A(n_82),
.Y(n_707)
);

INVx1_ASAP7_75t_L g708 ( 
.A(n_381),
.Y(n_708)
);

CKINVDCx5p33_ASAP7_75t_R g709 ( 
.A(n_343),
.Y(n_709)
);

INVx1_ASAP7_75t_L g710 ( 
.A(n_174),
.Y(n_710)
);

CKINVDCx5p33_ASAP7_75t_R g711 ( 
.A(n_413),
.Y(n_711)
);

INVx1_ASAP7_75t_L g712 ( 
.A(n_95),
.Y(n_712)
);

CKINVDCx5p33_ASAP7_75t_R g713 ( 
.A(n_196),
.Y(n_713)
);

CKINVDCx5p33_ASAP7_75t_R g714 ( 
.A(n_36),
.Y(n_714)
);

INVx1_ASAP7_75t_L g715 ( 
.A(n_394),
.Y(n_715)
);

CKINVDCx5p33_ASAP7_75t_R g716 ( 
.A(n_195),
.Y(n_716)
);

CKINVDCx5p33_ASAP7_75t_R g717 ( 
.A(n_32),
.Y(n_717)
);

CKINVDCx20_ASAP7_75t_R g718 ( 
.A(n_424),
.Y(n_718)
);

CKINVDCx5p33_ASAP7_75t_R g719 ( 
.A(n_355),
.Y(n_719)
);

INVx1_ASAP7_75t_L g720 ( 
.A(n_252),
.Y(n_720)
);

CKINVDCx20_ASAP7_75t_R g721 ( 
.A(n_126),
.Y(n_721)
);

INVx1_ASAP7_75t_L g722 ( 
.A(n_220),
.Y(n_722)
);

CKINVDCx20_ASAP7_75t_R g723 ( 
.A(n_344),
.Y(n_723)
);

INVx1_ASAP7_75t_SL g724 ( 
.A(n_163),
.Y(n_724)
);

INVx1_ASAP7_75t_L g725 ( 
.A(n_146),
.Y(n_725)
);

CKINVDCx5p33_ASAP7_75t_R g726 ( 
.A(n_30),
.Y(n_726)
);

CKINVDCx5p33_ASAP7_75t_R g727 ( 
.A(n_94),
.Y(n_727)
);

INVx1_ASAP7_75t_L g728 ( 
.A(n_425),
.Y(n_728)
);

CKINVDCx5p33_ASAP7_75t_R g729 ( 
.A(n_80),
.Y(n_729)
);

CKINVDCx5p33_ASAP7_75t_R g730 ( 
.A(n_339),
.Y(n_730)
);

CKINVDCx5p33_ASAP7_75t_R g731 ( 
.A(n_127),
.Y(n_731)
);

CKINVDCx5p33_ASAP7_75t_R g732 ( 
.A(n_207),
.Y(n_732)
);

INVx1_ASAP7_75t_L g733 ( 
.A(n_83),
.Y(n_733)
);

CKINVDCx5p33_ASAP7_75t_R g734 ( 
.A(n_382),
.Y(n_734)
);

INVx1_ASAP7_75t_L g735 ( 
.A(n_248),
.Y(n_735)
);

INVx1_ASAP7_75t_L g736 ( 
.A(n_359),
.Y(n_736)
);

CKINVDCx20_ASAP7_75t_R g737 ( 
.A(n_389),
.Y(n_737)
);

INVx2_ASAP7_75t_L g738 ( 
.A(n_408),
.Y(n_738)
);

CKINVDCx5p33_ASAP7_75t_R g739 ( 
.A(n_197),
.Y(n_739)
);

CKINVDCx20_ASAP7_75t_R g740 ( 
.A(n_16),
.Y(n_740)
);

CKINVDCx20_ASAP7_75t_R g741 ( 
.A(n_155),
.Y(n_741)
);

INVx1_ASAP7_75t_L g742 ( 
.A(n_380),
.Y(n_742)
);

CKINVDCx5p33_ASAP7_75t_R g743 ( 
.A(n_23),
.Y(n_743)
);

CKINVDCx5p33_ASAP7_75t_R g744 ( 
.A(n_272),
.Y(n_744)
);

INVx1_ASAP7_75t_L g745 ( 
.A(n_50),
.Y(n_745)
);

CKINVDCx5p33_ASAP7_75t_R g746 ( 
.A(n_156),
.Y(n_746)
);

CKINVDCx5p33_ASAP7_75t_R g747 ( 
.A(n_364),
.Y(n_747)
);

CKINVDCx5p33_ASAP7_75t_R g748 ( 
.A(n_280),
.Y(n_748)
);

INVx1_ASAP7_75t_L g749 ( 
.A(n_418),
.Y(n_749)
);

INVxp67_ASAP7_75t_SL g750 ( 
.A(n_33),
.Y(n_750)
);

INVx2_ASAP7_75t_L g751 ( 
.A(n_98),
.Y(n_751)
);

BUFx2_ASAP7_75t_L g752 ( 
.A(n_91),
.Y(n_752)
);

INVx1_ASAP7_75t_L g753 ( 
.A(n_96),
.Y(n_753)
);

CKINVDCx5p33_ASAP7_75t_R g754 ( 
.A(n_36),
.Y(n_754)
);

CKINVDCx5p33_ASAP7_75t_R g755 ( 
.A(n_398),
.Y(n_755)
);

INVxp67_ASAP7_75t_L g756 ( 
.A(n_261),
.Y(n_756)
);

INVx1_ASAP7_75t_L g757 ( 
.A(n_104),
.Y(n_757)
);

CKINVDCx5p33_ASAP7_75t_R g758 ( 
.A(n_340),
.Y(n_758)
);

CKINVDCx5p33_ASAP7_75t_R g759 ( 
.A(n_264),
.Y(n_759)
);

INVx1_ASAP7_75t_SL g760 ( 
.A(n_8),
.Y(n_760)
);

INVx1_ASAP7_75t_L g761 ( 
.A(n_135),
.Y(n_761)
);

INVx1_ASAP7_75t_L g762 ( 
.A(n_193),
.Y(n_762)
);

CKINVDCx5p33_ASAP7_75t_R g763 ( 
.A(n_3),
.Y(n_763)
);

CKINVDCx5p33_ASAP7_75t_R g764 ( 
.A(n_50),
.Y(n_764)
);

CKINVDCx5p33_ASAP7_75t_R g765 ( 
.A(n_125),
.Y(n_765)
);

INVx1_ASAP7_75t_L g766 ( 
.A(n_173),
.Y(n_766)
);

CKINVDCx5p33_ASAP7_75t_R g767 ( 
.A(n_64),
.Y(n_767)
);

CKINVDCx5p33_ASAP7_75t_R g768 ( 
.A(n_105),
.Y(n_768)
);

CKINVDCx20_ASAP7_75t_R g769 ( 
.A(n_18),
.Y(n_769)
);

CKINVDCx5p33_ASAP7_75t_R g770 ( 
.A(n_134),
.Y(n_770)
);

CKINVDCx5p33_ASAP7_75t_R g771 ( 
.A(n_70),
.Y(n_771)
);

CKINVDCx5p33_ASAP7_75t_R g772 ( 
.A(n_318),
.Y(n_772)
);

BUFx6f_ASAP7_75t_L g773 ( 
.A(n_302),
.Y(n_773)
);

CKINVDCx5p33_ASAP7_75t_R g774 ( 
.A(n_110),
.Y(n_774)
);

CKINVDCx5p33_ASAP7_75t_R g775 ( 
.A(n_392),
.Y(n_775)
);

INVx2_ASAP7_75t_L g776 ( 
.A(n_384),
.Y(n_776)
);

CKINVDCx20_ASAP7_75t_R g777 ( 
.A(n_111),
.Y(n_777)
);

BUFx2_ASAP7_75t_L g778 ( 
.A(n_324),
.Y(n_778)
);

INVx1_ASAP7_75t_L g779 ( 
.A(n_332),
.Y(n_779)
);

BUFx3_ASAP7_75t_L g780 ( 
.A(n_11),
.Y(n_780)
);

CKINVDCx5p33_ASAP7_75t_R g781 ( 
.A(n_71),
.Y(n_781)
);

CKINVDCx5p33_ASAP7_75t_R g782 ( 
.A(n_348),
.Y(n_782)
);

INVx1_ASAP7_75t_L g783 ( 
.A(n_400),
.Y(n_783)
);

CKINVDCx5p33_ASAP7_75t_R g784 ( 
.A(n_147),
.Y(n_784)
);

CKINVDCx5p33_ASAP7_75t_R g785 ( 
.A(n_192),
.Y(n_785)
);

INVx1_ASAP7_75t_L g786 ( 
.A(n_203),
.Y(n_786)
);

CKINVDCx5p33_ASAP7_75t_R g787 ( 
.A(n_331),
.Y(n_787)
);

INVx2_ASAP7_75t_L g788 ( 
.A(n_230),
.Y(n_788)
);

CKINVDCx5p33_ASAP7_75t_R g789 ( 
.A(n_377),
.Y(n_789)
);

INVx1_ASAP7_75t_SL g790 ( 
.A(n_1),
.Y(n_790)
);

CKINVDCx5p33_ASAP7_75t_R g791 ( 
.A(n_356),
.Y(n_791)
);

BUFx2_ASAP7_75t_L g792 ( 
.A(n_327),
.Y(n_792)
);

CKINVDCx5p33_ASAP7_75t_R g793 ( 
.A(n_169),
.Y(n_793)
);

BUFx10_ASAP7_75t_L g794 ( 
.A(n_97),
.Y(n_794)
);

CKINVDCx20_ASAP7_75t_R g795 ( 
.A(n_433),
.Y(n_795)
);

INVx1_ASAP7_75t_L g796 ( 
.A(n_566),
.Y(n_796)
);

INVx1_ASAP7_75t_L g797 ( 
.A(n_566),
.Y(n_797)
);

INVxp67_ASAP7_75t_SL g798 ( 
.A(n_566),
.Y(n_798)
);

INVx1_ASAP7_75t_L g799 ( 
.A(n_457),
.Y(n_799)
);

INVxp67_ASAP7_75t_L g800 ( 
.A(n_435),
.Y(n_800)
);

CKINVDCx5p33_ASAP7_75t_R g801 ( 
.A(n_655),
.Y(n_801)
);

INVxp33_ASAP7_75t_SL g802 ( 
.A(n_568),
.Y(n_802)
);

INVxp67_ASAP7_75t_SL g803 ( 
.A(n_457),
.Y(n_803)
);

INVxp33_ASAP7_75t_L g804 ( 
.A(n_435),
.Y(n_804)
);

INVxp33_ASAP7_75t_SL g805 ( 
.A(n_540),
.Y(n_805)
);

CKINVDCx20_ASAP7_75t_R g806 ( 
.A(n_442),
.Y(n_806)
);

BUFx3_ASAP7_75t_L g807 ( 
.A(n_534),
.Y(n_807)
);

INVx1_ASAP7_75t_L g808 ( 
.A(n_464),
.Y(n_808)
);

INVx1_ASAP7_75t_L g809 ( 
.A(n_464),
.Y(n_809)
);

INVx1_ASAP7_75t_L g810 ( 
.A(n_499),
.Y(n_810)
);

CKINVDCx5p33_ASAP7_75t_R g811 ( 
.A(n_665),
.Y(n_811)
);

CKINVDCx14_ASAP7_75t_R g812 ( 
.A(n_516),
.Y(n_812)
);

INVx1_ASAP7_75t_L g813 ( 
.A(n_499),
.Y(n_813)
);

NOR2xp33_ASAP7_75t_L g814 ( 
.A(n_534),
.B(n_1),
.Y(n_814)
);

BUFx3_ASAP7_75t_L g815 ( 
.A(n_622),
.Y(n_815)
);

CKINVDCx20_ASAP7_75t_R g816 ( 
.A(n_451),
.Y(n_816)
);

INVx1_ASAP7_75t_L g817 ( 
.A(n_501),
.Y(n_817)
);

INVx1_ASAP7_75t_L g818 ( 
.A(n_501),
.Y(n_818)
);

INVx1_ASAP7_75t_L g819 ( 
.A(n_517),
.Y(n_819)
);

INVx1_ASAP7_75t_L g820 ( 
.A(n_517),
.Y(n_820)
);

BUFx3_ASAP7_75t_L g821 ( 
.A(n_622),
.Y(n_821)
);

INVx1_ASAP7_75t_L g822 ( 
.A(n_591),
.Y(n_822)
);

INVx1_ASAP7_75t_L g823 ( 
.A(n_591),
.Y(n_823)
);

INVxp67_ASAP7_75t_SL g824 ( 
.A(n_609),
.Y(n_824)
);

CKINVDCx16_ASAP7_75t_R g825 ( 
.A(n_458),
.Y(n_825)
);

INVx2_ASAP7_75t_L g826 ( 
.A(n_582),
.Y(n_826)
);

INVx1_ASAP7_75t_L g827 ( 
.A(n_609),
.Y(n_827)
);

INVx1_ASAP7_75t_L g828 ( 
.A(n_780),
.Y(n_828)
);

CKINVDCx5p33_ASAP7_75t_R g829 ( 
.A(n_637),
.Y(n_829)
);

INVx1_ASAP7_75t_L g830 ( 
.A(n_780),
.Y(n_830)
);

INVx1_ASAP7_75t_L g831 ( 
.A(n_540),
.Y(n_831)
);

CKINVDCx14_ASAP7_75t_R g832 ( 
.A(n_664),
.Y(n_832)
);

INVx1_ASAP7_75t_L g833 ( 
.A(n_752),
.Y(n_833)
);

INVx2_ASAP7_75t_L g834 ( 
.A(n_582),
.Y(n_834)
);

CKINVDCx5p33_ASAP7_75t_R g835 ( 
.A(n_637),
.Y(n_835)
);

INVx1_ASAP7_75t_L g836 ( 
.A(n_752),
.Y(n_836)
);

INVx1_ASAP7_75t_L g837 ( 
.A(n_778),
.Y(n_837)
);

INVx1_ASAP7_75t_L g838 ( 
.A(n_778),
.Y(n_838)
);

NAND2xp5_ASAP7_75t_L g839 ( 
.A(n_792),
.B(n_2),
.Y(n_839)
);

CKINVDCx5p33_ASAP7_75t_R g840 ( 
.A(n_792),
.Y(n_840)
);

INVx1_ASAP7_75t_L g841 ( 
.A(n_439),
.Y(n_841)
);

INVxp33_ASAP7_75t_SL g842 ( 
.A(n_427),
.Y(n_842)
);

INVx1_ASAP7_75t_L g843 ( 
.A(n_439),
.Y(n_843)
);

INVx1_ASAP7_75t_L g844 ( 
.A(n_446),
.Y(n_844)
);

CKINVDCx20_ASAP7_75t_R g845 ( 
.A(n_463),
.Y(n_845)
);

INVxp33_ASAP7_75t_SL g846 ( 
.A(n_434),
.Y(n_846)
);

INVx1_ASAP7_75t_L g847 ( 
.A(n_446),
.Y(n_847)
);

INVx1_ASAP7_75t_L g848 ( 
.A(n_452),
.Y(n_848)
);

INVx1_ASAP7_75t_L g849 ( 
.A(n_452),
.Y(n_849)
);

INVx1_ASAP7_75t_L g850 ( 
.A(n_453),
.Y(n_850)
);

INVxp67_ASAP7_75t_L g851 ( 
.A(n_453),
.Y(n_851)
);

INVxp67_ASAP7_75t_SL g852 ( 
.A(n_582),
.Y(n_852)
);

INVx1_ASAP7_75t_L g853 ( 
.A(n_466),
.Y(n_853)
);

INVx1_ASAP7_75t_L g854 ( 
.A(n_466),
.Y(n_854)
);

INVxp67_ASAP7_75t_SL g855 ( 
.A(n_582),
.Y(n_855)
);

CKINVDCx5p33_ASAP7_75t_R g856 ( 
.A(n_533),
.Y(n_856)
);

INVx1_ASAP7_75t_L g857 ( 
.A(n_482),
.Y(n_857)
);

INVx1_ASAP7_75t_L g858 ( 
.A(n_482),
.Y(n_858)
);

INVx2_ASAP7_75t_L g859 ( 
.A(n_428),
.Y(n_859)
);

INVx1_ASAP7_75t_L g860 ( 
.A(n_489),
.Y(n_860)
);

INVx1_ASAP7_75t_L g861 ( 
.A(n_489),
.Y(n_861)
);

CKINVDCx16_ASAP7_75t_R g862 ( 
.A(n_581),
.Y(n_862)
);

INVx1_ASAP7_75t_L g863 ( 
.A(n_515),
.Y(n_863)
);

INVx1_ASAP7_75t_L g864 ( 
.A(n_515),
.Y(n_864)
);

INVx1_ASAP7_75t_L g865 ( 
.A(n_520),
.Y(n_865)
);

INVx1_ASAP7_75t_L g866 ( 
.A(n_520),
.Y(n_866)
);

NOR2xp67_ASAP7_75t_L g867 ( 
.A(n_477),
.B(n_2),
.Y(n_867)
);

INVx1_ASAP7_75t_L g868 ( 
.A(n_539),
.Y(n_868)
);

HB1xp67_ASAP7_75t_L g869 ( 
.A(n_436),
.Y(n_869)
);

HB1xp67_ASAP7_75t_L g870 ( 
.A(n_437),
.Y(n_870)
);

INVx1_ASAP7_75t_L g871 ( 
.A(n_539),
.Y(n_871)
);

INVx1_ASAP7_75t_L g872 ( 
.A(n_548),
.Y(n_872)
);

INVxp33_ASAP7_75t_SL g873 ( 
.A(n_441),
.Y(n_873)
);

INVx1_ASAP7_75t_L g874 ( 
.A(n_548),
.Y(n_874)
);

INVx1_ASAP7_75t_L g875 ( 
.A(n_553),
.Y(n_875)
);

BUFx6f_ASAP7_75t_L g876 ( 
.A(n_426),
.Y(n_876)
);

INVx1_ASAP7_75t_L g877 ( 
.A(n_553),
.Y(n_877)
);

INVx1_ASAP7_75t_L g878 ( 
.A(n_555),
.Y(n_878)
);

INVxp67_ASAP7_75t_L g879 ( 
.A(n_555),
.Y(n_879)
);

INVx1_ASAP7_75t_L g880 ( 
.A(n_557),
.Y(n_880)
);

INVxp33_ASAP7_75t_L g881 ( 
.A(n_507),
.Y(n_881)
);

CKINVDCx16_ASAP7_75t_R g882 ( 
.A(n_581),
.Y(n_882)
);

INVx1_ASAP7_75t_L g883 ( 
.A(n_557),
.Y(n_883)
);

INVx1_ASAP7_75t_L g884 ( 
.A(n_559),
.Y(n_884)
);

INVx1_ASAP7_75t_L g885 ( 
.A(n_559),
.Y(n_885)
);

BUFx3_ASAP7_75t_L g886 ( 
.A(n_554),
.Y(n_886)
);

INVx1_ASAP7_75t_L g887 ( 
.A(n_573),
.Y(n_887)
);

INVx1_ASAP7_75t_L g888 ( 
.A(n_573),
.Y(n_888)
);

INVx1_ASAP7_75t_L g889 ( 
.A(n_601),
.Y(n_889)
);

INVx1_ASAP7_75t_L g890 ( 
.A(n_601),
.Y(n_890)
);

INVx1_ASAP7_75t_L g891 ( 
.A(n_615),
.Y(n_891)
);

INVx1_ASAP7_75t_L g892 ( 
.A(n_615),
.Y(n_892)
);

INVx1_ASAP7_75t_L g893 ( 
.A(n_616),
.Y(n_893)
);

INVx2_ASAP7_75t_L g894 ( 
.A(n_428),
.Y(n_894)
);

INVx1_ASAP7_75t_L g895 ( 
.A(n_616),
.Y(n_895)
);

INVxp67_ASAP7_75t_SL g896 ( 
.A(n_617),
.Y(n_896)
);

INVxp33_ASAP7_75t_SL g897 ( 
.A(n_445),
.Y(n_897)
);

INVx1_ASAP7_75t_L g898 ( 
.A(n_617),
.Y(n_898)
);

INVxp67_ASAP7_75t_L g899 ( 
.A(n_636),
.Y(n_899)
);

INVx1_ASAP7_75t_L g900 ( 
.A(n_636),
.Y(n_900)
);

INVx1_ASAP7_75t_SL g901 ( 
.A(n_484),
.Y(n_901)
);

INVxp67_ASAP7_75t_L g902 ( 
.A(n_638),
.Y(n_902)
);

INVx1_ASAP7_75t_L g903 ( 
.A(n_638),
.Y(n_903)
);

CKINVDCx5p33_ASAP7_75t_R g904 ( 
.A(n_448),
.Y(n_904)
);

INVx1_ASAP7_75t_L g905 ( 
.A(n_643),
.Y(n_905)
);

INVx1_ASAP7_75t_L g906 ( 
.A(n_643),
.Y(n_906)
);

INVx1_ASAP7_75t_L g907 ( 
.A(n_647),
.Y(n_907)
);

INVx1_ASAP7_75t_L g908 ( 
.A(n_647),
.Y(n_908)
);

INVx1_ASAP7_75t_L g909 ( 
.A(n_659),
.Y(n_909)
);

INVx1_ASAP7_75t_L g910 ( 
.A(n_659),
.Y(n_910)
);

INVxp33_ASAP7_75t_SL g911 ( 
.A(n_447),
.Y(n_911)
);

INVx1_ASAP7_75t_L g912 ( 
.A(n_672),
.Y(n_912)
);

INVx2_ASAP7_75t_L g913 ( 
.A(n_432),
.Y(n_913)
);

CKINVDCx5p33_ASAP7_75t_R g914 ( 
.A(n_448),
.Y(n_914)
);

INVx1_ASAP7_75t_L g915 ( 
.A(n_672),
.Y(n_915)
);

INVx1_ASAP7_75t_L g916 ( 
.A(n_679),
.Y(n_916)
);

INVx1_ASAP7_75t_L g917 ( 
.A(n_679),
.Y(n_917)
);

INVx1_ASAP7_75t_L g918 ( 
.A(n_680),
.Y(n_918)
);

CKINVDCx5p33_ASAP7_75t_R g919 ( 
.A(n_448),
.Y(n_919)
);

INVx1_ASAP7_75t_L g920 ( 
.A(n_680),
.Y(n_920)
);

INVx1_ASAP7_75t_L g921 ( 
.A(n_684),
.Y(n_921)
);

INVxp33_ASAP7_75t_L g922 ( 
.A(n_507),
.Y(n_922)
);

INVx1_ASAP7_75t_L g923 ( 
.A(n_684),
.Y(n_923)
);

CKINVDCx5p33_ASAP7_75t_R g924 ( 
.A(n_430),
.Y(n_924)
);

CKINVDCx16_ASAP7_75t_R g925 ( 
.A(n_581),
.Y(n_925)
);

INVx1_ASAP7_75t_L g926 ( 
.A(n_691),
.Y(n_926)
);

INVx1_ASAP7_75t_L g927 ( 
.A(n_691),
.Y(n_927)
);

HB1xp67_ASAP7_75t_L g928 ( 
.A(n_449),
.Y(n_928)
);

INVx1_ASAP7_75t_L g929 ( 
.A(n_692),
.Y(n_929)
);

INVx1_ASAP7_75t_L g930 ( 
.A(n_692),
.Y(n_930)
);

INVxp67_ASAP7_75t_L g931 ( 
.A(n_710),
.Y(n_931)
);

INVx1_ASAP7_75t_L g932 ( 
.A(n_710),
.Y(n_932)
);

INVx1_ASAP7_75t_L g933 ( 
.A(n_712),
.Y(n_933)
);

INVx1_ASAP7_75t_L g934 ( 
.A(n_712),
.Y(n_934)
);

CKINVDCx20_ASAP7_75t_R g935 ( 
.A(n_527),
.Y(n_935)
);

INVx1_ASAP7_75t_L g936 ( 
.A(n_725),
.Y(n_936)
);

NOR2xp33_ASAP7_75t_L g937 ( 
.A(n_432),
.B(n_3),
.Y(n_937)
);

INVx1_ASAP7_75t_L g938 ( 
.A(n_725),
.Y(n_938)
);

INVx1_ASAP7_75t_L g939 ( 
.A(n_733),
.Y(n_939)
);

INVxp33_ASAP7_75t_L g940 ( 
.A(n_546),
.Y(n_940)
);

CKINVDCx20_ASAP7_75t_R g941 ( 
.A(n_537),
.Y(n_941)
);

CKINVDCx5p33_ASAP7_75t_R g942 ( 
.A(n_431),
.Y(n_942)
);

CKINVDCx5p33_ASAP7_75t_R g943 ( 
.A(n_438),
.Y(n_943)
);

INVx1_ASAP7_75t_L g944 ( 
.A(n_733),
.Y(n_944)
);

INVx2_ASAP7_75t_L g945 ( 
.A(n_443),
.Y(n_945)
);

INVx1_ASAP7_75t_L g946 ( 
.A(n_745),
.Y(n_946)
);

INVx2_ASAP7_75t_L g947 ( 
.A(n_443),
.Y(n_947)
);

INVx1_ASAP7_75t_L g948 ( 
.A(n_745),
.Y(n_948)
);

INVx1_ASAP7_75t_L g949 ( 
.A(n_753),
.Y(n_949)
);

CKINVDCx16_ASAP7_75t_R g950 ( 
.A(n_618),
.Y(n_950)
);

INVx1_ASAP7_75t_L g951 ( 
.A(n_753),
.Y(n_951)
);

BUFx6f_ASAP7_75t_L g952 ( 
.A(n_426),
.Y(n_952)
);

INVxp67_ASAP7_75t_SL g953 ( 
.A(n_757),
.Y(n_953)
);

INVxp67_ASAP7_75t_L g954 ( 
.A(n_757),
.Y(n_954)
);

INVx1_ASAP7_75t_L g955 ( 
.A(n_761),
.Y(n_955)
);

INVx1_ASAP7_75t_L g956 ( 
.A(n_761),
.Y(n_956)
);

CKINVDCx16_ASAP7_75t_R g957 ( 
.A(n_618),
.Y(n_957)
);

BUFx5_ASAP7_75t_L g958 ( 
.A(n_450),
.Y(n_958)
);

HB1xp67_ASAP7_75t_L g959 ( 
.A(n_459),
.Y(n_959)
);

NOR2xp67_ASAP7_75t_L g960 ( 
.A(n_477),
.B(n_5),
.Y(n_960)
);

INVxp33_ASAP7_75t_SL g961 ( 
.A(n_470),
.Y(n_961)
);

INVx1_ASAP7_75t_L g962 ( 
.A(n_762),
.Y(n_962)
);

INVx1_ASAP7_75t_L g963 ( 
.A(n_762),
.Y(n_963)
);

INVx2_ASAP7_75t_L g964 ( 
.A(n_450),
.Y(n_964)
);

CKINVDCx16_ASAP7_75t_R g965 ( 
.A(n_618),
.Y(n_965)
);

INVx1_ASAP7_75t_L g966 ( 
.A(n_766),
.Y(n_966)
);

INVxp67_ASAP7_75t_L g967 ( 
.A(n_766),
.Y(n_967)
);

INVxp33_ASAP7_75t_L g968 ( 
.A(n_546),
.Y(n_968)
);

INVx1_ASAP7_75t_L g969 ( 
.A(n_786),
.Y(n_969)
);

CKINVDCx5p33_ASAP7_75t_R g970 ( 
.A(n_535),
.Y(n_970)
);

INVxp67_ASAP7_75t_SL g971 ( 
.A(n_786),
.Y(n_971)
);

INVx1_ASAP7_75t_L g972 ( 
.A(n_525),
.Y(n_972)
);

INVxp33_ASAP7_75t_L g973 ( 
.A(n_574),
.Y(n_973)
);

INVx1_ASAP7_75t_L g974 ( 
.A(n_530),
.Y(n_974)
);

CKINVDCx5p33_ASAP7_75t_R g975 ( 
.A(n_541),
.Y(n_975)
);

INVxp67_ASAP7_75t_SL g976 ( 
.A(n_574),
.Y(n_976)
);

INVxp33_ASAP7_75t_SL g977 ( 
.A(n_473),
.Y(n_977)
);

INVx1_ASAP7_75t_L g978 ( 
.A(n_570),
.Y(n_978)
);

INVx2_ASAP7_75t_L g979 ( 
.A(n_460),
.Y(n_979)
);

INVx1_ASAP7_75t_L g980 ( 
.A(n_625),
.Y(n_980)
);

INVx1_ASAP7_75t_L g981 ( 
.A(n_630),
.Y(n_981)
);

INVx1_ASAP7_75t_L g982 ( 
.A(n_632),
.Y(n_982)
);

CKINVDCx16_ASAP7_75t_R g983 ( 
.A(n_794),
.Y(n_983)
);

INVx1_ASAP7_75t_L g984 ( 
.A(n_623),
.Y(n_984)
);

CKINVDCx5p33_ASAP7_75t_R g985 ( 
.A(n_542),
.Y(n_985)
);

INVx1_ASAP7_75t_L g986 ( 
.A(n_623),
.Y(n_986)
);

INVxp67_ASAP7_75t_SL g987 ( 
.A(n_751),
.Y(n_987)
);

INVxp33_ASAP7_75t_L g988 ( 
.A(n_751),
.Y(n_988)
);

CKINVDCx20_ASAP7_75t_R g989 ( 
.A(n_562),
.Y(n_989)
);

INVxp67_ASAP7_75t_SL g990 ( 
.A(n_687),
.Y(n_990)
);

CKINVDCx5p33_ASAP7_75t_R g991 ( 
.A(n_572),
.Y(n_991)
);

INVx1_ASAP7_75t_L g992 ( 
.A(n_687),
.Y(n_992)
);

INVxp67_ASAP7_75t_SL g993 ( 
.A(n_500),
.Y(n_993)
);

CKINVDCx5p33_ASAP7_75t_R g994 ( 
.A(n_662),
.Y(n_994)
);

INVx2_ASAP7_75t_L g995 ( 
.A(n_460),
.Y(n_995)
);

INVx1_ASAP7_75t_L g996 ( 
.A(n_467),
.Y(n_996)
);

CKINVDCx20_ASAP7_75t_R g997 ( 
.A(n_596),
.Y(n_997)
);

INVx1_ASAP7_75t_SL g998 ( 
.A(n_602),
.Y(n_998)
);

INVxp67_ASAP7_75t_SL g999 ( 
.A(n_571),
.Y(n_999)
);

INVx1_ASAP7_75t_L g1000 ( 
.A(n_467),
.Y(n_1000)
);

INVx1_ASAP7_75t_L g1001 ( 
.A(n_468),
.Y(n_1001)
);

INVxp67_ASAP7_75t_SL g1002 ( 
.A(n_554),
.Y(n_1002)
);

INVx1_ASAP7_75t_L g1003 ( 
.A(n_468),
.Y(n_1003)
);

INVxp67_ASAP7_75t_SL g1004 ( 
.A(n_611),
.Y(n_1004)
);

INVx2_ASAP7_75t_L g1005 ( 
.A(n_469),
.Y(n_1005)
);

INVx1_ASAP7_75t_L g1006 ( 
.A(n_469),
.Y(n_1006)
);

CKINVDCx16_ASAP7_75t_R g1007 ( 
.A(n_794),
.Y(n_1007)
);

CKINVDCx16_ASAP7_75t_R g1008 ( 
.A(n_794),
.Y(n_1008)
);

INVx1_ASAP7_75t_L g1009 ( 
.A(n_472),
.Y(n_1009)
);

INVx1_ASAP7_75t_L g1010 ( 
.A(n_472),
.Y(n_1010)
);

INVx1_ASAP7_75t_L g1011 ( 
.A(n_474),
.Y(n_1011)
);

INVx1_ASAP7_75t_L g1012 ( 
.A(n_474),
.Y(n_1012)
);

INVx1_ASAP7_75t_L g1013 ( 
.A(n_479),
.Y(n_1013)
);

INVx1_ASAP7_75t_L g1014 ( 
.A(n_479),
.Y(n_1014)
);

CKINVDCx16_ASAP7_75t_R g1015 ( 
.A(n_666),
.Y(n_1015)
);

INVxp67_ASAP7_75t_SL g1016 ( 
.A(n_611),
.Y(n_1016)
);

INVx1_ASAP7_75t_L g1017 ( 
.A(n_490),
.Y(n_1017)
);

INVx1_ASAP7_75t_L g1018 ( 
.A(n_490),
.Y(n_1018)
);

INVx2_ASAP7_75t_L g1019 ( 
.A(n_493),
.Y(n_1019)
);

INVxp67_ASAP7_75t_SL g1020 ( 
.A(n_642),
.Y(n_1020)
);

INVx1_ASAP7_75t_L g1021 ( 
.A(n_493),
.Y(n_1021)
);

INVx1_ASAP7_75t_L g1022 ( 
.A(n_502),
.Y(n_1022)
);

CKINVDCx20_ASAP7_75t_R g1023 ( 
.A(n_606),
.Y(n_1023)
);

INVx1_ASAP7_75t_L g1024 ( 
.A(n_502),
.Y(n_1024)
);

CKINVDCx20_ASAP7_75t_R g1025 ( 
.A(n_612),
.Y(n_1025)
);

INVx1_ASAP7_75t_L g1026 ( 
.A(n_505),
.Y(n_1026)
);

INVxp33_ASAP7_75t_SL g1027 ( 
.A(n_478),
.Y(n_1027)
);

INVxp67_ASAP7_75t_SL g1028 ( 
.A(n_642),
.Y(n_1028)
);

INVx1_ASAP7_75t_L g1029 ( 
.A(n_505),
.Y(n_1029)
);

INVx1_ASAP7_75t_L g1030 ( 
.A(n_513),
.Y(n_1030)
);

INVx2_ASAP7_75t_L g1031 ( 
.A(n_513),
.Y(n_1031)
);

INVx1_ASAP7_75t_L g1032 ( 
.A(n_531),
.Y(n_1032)
);

INVx1_ASAP7_75t_L g1033 ( 
.A(n_531),
.Y(n_1033)
);

INVxp67_ASAP7_75t_SL g1034 ( 
.A(n_701),
.Y(n_1034)
);

INVx1_ASAP7_75t_L g1035 ( 
.A(n_536),
.Y(n_1035)
);

INVxp67_ASAP7_75t_SL g1036 ( 
.A(n_701),
.Y(n_1036)
);

INVx1_ASAP7_75t_L g1037 ( 
.A(n_536),
.Y(n_1037)
);

INVx1_ASAP7_75t_L g1038 ( 
.A(n_538),
.Y(n_1038)
);

INVx1_ASAP7_75t_L g1039 ( 
.A(n_538),
.Y(n_1039)
);

INVx1_ASAP7_75t_L g1040 ( 
.A(n_547),
.Y(n_1040)
);

INVx1_ASAP7_75t_L g1041 ( 
.A(n_547),
.Y(n_1041)
);

INVx1_ASAP7_75t_L g1042 ( 
.A(n_560),
.Y(n_1042)
);

INVx1_ASAP7_75t_L g1043 ( 
.A(n_560),
.Y(n_1043)
);

INVxp67_ASAP7_75t_SL g1044 ( 
.A(n_750),
.Y(n_1044)
);

CKINVDCx5p33_ASAP7_75t_R g1045 ( 
.A(n_702),
.Y(n_1045)
);

INVx1_ASAP7_75t_L g1046 ( 
.A(n_564),
.Y(n_1046)
);

INVx1_ASAP7_75t_L g1047 ( 
.A(n_564),
.Y(n_1047)
);

INVx1_ASAP7_75t_L g1048 ( 
.A(n_565),
.Y(n_1048)
);

CKINVDCx20_ASAP7_75t_R g1049 ( 
.A(n_624),
.Y(n_1049)
);

INVx1_ASAP7_75t_L g1050 ( 
.A(n_565),
.Y(n_1050)
);

CKINVDCx5p33_ASAP7_75t_R g1051 ( 
.A(n_718),
.Y(n_1051)
);

INVxp67_ASAP7_75t_SL g1052 ( 
.A(n_567),
.Y(n_1052)
);

INVx1_ASAP7_75t_L g1053 ( 
.A(n_567),
.Y(n_1053)
);

INVx1_ASAP7_75t_L g1054 ( 
.A(n_593),
.Y(n_1054)
);

INVxp33_ASAP7_75t_SL g1055 ( 
.A(n_483),
.Y(n_1055)
);

INVxp33_ASAP7_75t_SL g1056 ( 
.A(n_485),
.Y(n_1056)
);

BUFx3_ASAP7_75t_L g1057 ( 
.A(n_593),
.Y(n_1057)
);

CKINVDCx16_ASAP7_75t_R g1058 ( 
.A(n_723),
.Y(n_1058)
);

INVx1_ASAP7_75t_L g1059 ( 
.A(n_608),
.Y(n_1059)
);

INVx3_ASAP7_75t_L g1060 ( 
.A(n_608),
.Y(n_1060)
);

INVx1_ASAP7_75t_L g1061 ( 
.A(n_635),
.Y(n_1061)
);

INVx2_ASAP7_75t_L g1062 ( 
.A(n_635),
.Y(n_1062)
);

INVx2_ASAP7_75t_L g1063 ( 
.A(n_654),
.Y(n_1063)
);

CKINVDCx20_ASAP7_75t_R g1064 ( 
.A(n_626),
.Y(n_1064)
);

CKINVDCx20_ASAP7_75t_R g1065 ( 
.A(n_646),
.Y(n_1065)
);

CKINVDCx20_ASAP7_75t_R g1066 ( 
.A(n_682),
.Y(n_1066)
);

INVx1_ASAP7_75t_L g1067 ( 
.A(n_654),
.Y(n_1067)
);

CKINVDCx20_ASAP7_75t_R g1068 ( 
.A(n_683),
.Y(n_1068)
);

INVx1_ASAP7_75t_L g1069 ( 
.A(n_668),
.Y(n_1069)
);

INVx1_ASAP7_75t_L g1070 ( 
.A(n_668),
.Y(n_1070)
);

INVx1_ASAP7_75t_L g1071 ( 
.A(n_670),
.Y(n_1071)
);

BUFx3_ASAP7_75t_L g1072 ( 
.A(n_670),
.Y(n_1072)
);

INVx1_ASAP7_75t_L g1073 ( 
.A(n_676),
.Y(n_1073)
);

INVxp33_ASAP7_75t_SL g1074 ( 
.A(n_486),
.Y(n_1074)
);

INVx1_ASAP7_75t_L g1075 ( 
.A(n_676),
.Y(n_1075)
);

CKINVDCx5p33_ASAP7_75t_R g1076 ( 
.A(n_737),
.Y(n_1076)
);

INVx1_ASAP7_75t_L g1077 ( 
.A(n_685),
.Y(n_1077)
);

BUFx6f_ASAP7_75t_L g1078 ( 
.A(n_426),
.Y(n_1078)
);

INVx1_ASAP7_75t_L g1079 ( 
.A(n_685),
.Y(n_1079)
);

INVx1_ASAP7_75t_L g1080 ( 
.A(n_697),
.Y(n_1080)
);

BUFx10_ASAP7_75t_L g1081 ( 
.A(n_471),
.Y(n_1081)
);

INVxp67_ASAP7_75t_L g1082 ( 
.A(n_488),
.Y(n_1082)
);

INVx1_ASAP7_75t_L g1083 ( 
.A(n_697),
.Y(n_1083)
);

INVxp67_ASAP7_75t_L g1084 ( 
.A(n_498),
.Y(n_1084)
);

INVx1_ASAP7_75t_L g1085 ( 
.A(n_698),
.Y(n_1085)
);

CKINVDCx5p33_ASAP7_75t_R g1086 ( 
.A(n_506),
.Y(n_1086)
);

INVx3_ASAP7_75t_L g1087 ( 
.A(n_886),
.Y(n_1087)
);

INVx1_ASAP7_75t_L g1088 ( 
.A(n_852),
.Y(n_1088)
);

BUFx3_ASAP7_75t_L g1089 ( 
.A(n_886),
.Y(n_1089)
);

NOR2xp33_ASAP7_75t_L g1090 ( 
.A(n_802),
.B(n_698),
.Y(n_1090)
);

AND2x4_ASAP7_75t_L g1091 ( 
.A(n_807),
.B(n_700),
.Y(n_1091)
);

NOR2xp33_ASAP7_75t_L g1092 ( 
.A(n_802),
.B(n_700),
.Y(n_1092)
);

INVx2_ASAP7_75t_L g1093 ( 
.A(n_826),
.Y(n_1093)
);

NAND2xp5_ASAP7_75t_L g1094 ( 
.A(n_1002),
.B(n_703),
.Y(n_1094)
);

BUFx8_ASAP7_75t_SL g1095 ( 
.A(n_795),
.Y(n_1095)
);

INVx4_ASAP7_75t_L g1096 ( 
.A(n_904),
.Y(n_1096)
);

INVx3_ASAP7_75t_L g1097 ( 
.A(n_1057),
.Y(n_1097)
);

INVx5_ASAP7_75t_L g1098 ( 
.A(n_876),
.Y(n_1098)
);

INVx2_ASAP7_75t_L g1099 ( 
.A(n_826),
.Y(n_1099)
);

INVx2_ASAP7_75t_L g1100 ( 
.A(n_834),
.Y(n_1100)
);

NAND2xp5_ASAP7_75t_L g1101 ( 
.A(n_1004),
.B(n_1016),
.Y(n_1101)
);

NOR2xp33_ASAP7_75t_SL g1102 ( 
.A(n_825),
.B(n_694),
.Y(n_1102)
);

BUFx6f_ASAP7_75t_L g1103 ( 
.A(n_876),
.Y(n_1103)
);

NOR2xp33_ASAP7_75t_L g1104 ( 
.A(n_1082),
.B(n_703),
.Y(n_1104)
);

INVx5_ASAP7_75t_L g1105 ( 
.A(n_876),
.Y(n_1105)
);

INVx1_ASAP7_75t_L g1106 ( 
.A(n_855),
.Y(n_1106)
);

CKINVDCx5p33_ASAP7_75t_R g1107 ( 
.A(n_812),
.Y(n_1107)
);

NAND2xp5_ASAP7_75t_L g1108 ( 
.A(n_1020),
.B(n_708),
.Y(n_1108)
);

BUFx3_ASAP7_75t_L g1109 ( 
.A(n_796),
.Y(n_1109)
);

AND2x4_ASAP7_75t_L g1110 ( 
.A(n_807),
.B(n_708),
.Y(n_1110)
);

BUFx8_ASAP7_75t_SL g1111 ( 
.A(n_795),
.Y(n_1111)
);

AND2x4_ASAP7_75t_L g1112 ( 
.A(n_815),
.B(n_715),
.Y(n_1112)
);

INVx2_ASAP7_75t_L g1113 ( 
.A(n_876),
.Y(n_1113)
);

NOR2xp33_ASAP7_75t_SL g1114 ( 
.A(n_856),
.B(n_695),
.Y(n_1114)
);

INVx5_ASAP7_75t_L g1115 ( 
.A(n_952),
.Y(n_1115)
);

AND2x2_ASAP7_75t_L g1116 ( 
.A(n_812),
.B(n_579),
.Y(n_1116)
);

INVx4_ASAP7_75t_L g1117 ( 
.A(n_904),
.Y(n_1117)
);

NOR2xp33_ASAP7_75t_L g1118 ( 
.A(n_1084),
.B(n_715),
.Y(n_1118)
);

NAND2xp5_ASAP7_75t_L g1119 ( 
.A(n_1028),
.B(n_720),
.Y(n_1119)
);

NOR2xp33_ASAP7_75t_L g1120 ( 
.A(n_798),
.B(n_720),
.Y(n_1120)
);

AND2x2_ASAP7_75t_L g1121 ( 
.A(n_832),
.B(n_641),
.Y(n_1121)
);

INVx4_ASAP7_75t_L g1122 ( 
.A(n_914),
.Y(n_1122)
);

BUFx6f_ASAP7_75t_L g1123 ( 
.A(n_952),
.Y(n_1123)
);

AND2x4_ASAP7_75t_L g1124 ( 
.A(n_815),
.B(n_722),
.Y(n_1124)
);

INVx5_ASAP7_75t_L g1125 ( 
.A(n_952),
.Y(n_1125)
);

INVx5_ASAP7_75t_L g1126 ( 
.A(n_952),
.Y(n_1126)
);

BUFx6f_ASAP7_75t_L g1127 ( 
.A(n_1078),
.Y(n_1127)
);

BUFx8_ASAP7_75t_L g1128 ( 
.A(n_831),
.Y(n_1128)
);

INVx5_ASAP7_75t_L g1129 ( 
.A(n_1078),
.Y(n_1129)
);

AND2x2_ASAP7_75t_L g1130 ( 
.A(n_832),
.B(n_658),
.Y(n_1130)
);

INVx3_ASAP7_75t_L g1131 ( 
.A(n_1057),
.Y(n_1131)
);

AND2x4_ASAP7_75t_L g1132 ( 
.A(n_821),
.B(n_722),
.Y(n_1132)
);

AND2x4_ASAP7_75t_L g1133 ( 
.A(n_821),
.B(n_837),
.Y(n_1133)
);

BUFx6f_ASAP7_75t_L g1134 ( 
.A(n_1078),
.Y(n_1134)
);

NAND2xp5_ASAP7_75t_L g1135 ( 
.A(n_1034),
.B(n_728),
.Y(n_1135)
);

BUFx8_ASAP7_75t_SL g1136 ( 
.A(n_806),
.Y(n_1136)
);

BUFx3_ASAP7_75t_L g1137 ( 
.A(n_797),
.Y(n_1137)
);

INVx2_ASAP7_75t_L g1138 ( 
.A(n_1078),
.Y(n_1138)
);

NAND2xp5_ASAP7_75t_L g1139 ( 
.A(n_1036),
.B(n_728),
.Y(n_1139)
);

CKINVDCx5p33_ASAP7_75t_R g1140 ( 
.A(n_924),
.Y(n_1140)
);

INVx4_ASAP7_75t_L g1141 ( 
.A(n_914),
.Y(n_1141)
);

INVx5_ASAP7_75t_L g1142 ( 
.A(n_1060),
.Y(n_1142)
);

NOR2xp33_ASAP7_75t_L g1143 ( 
.A(n_990),
.B(n_735),
.Y(n_1143)
);

NAND2xp5_ASAP7_75t_L g1144 ( 
.A(n_803),
.B(n_735),
.Y(n_1144)
);

INVx2_ASAP7_75t_L g1145 ( 
.A(n_958),
.Y(n_1145)
);

BUFx12f_ASAP7_75t_L g1146 ( 
.A(n_801),
.Y(n_1146)
);

INVx2_ASAP7_75t_L g1147 ( 
.A(n_958),
.Y(n_1147)
);

INVx2_ASAP7_75t_L g1148 ( 
.A(n_958),
.Y(n_1148)
);

INVx2_ASAP7_75t_L g1149 ( 
.A(n_958),
.Y(n_1149)
);

INVx2_ASAP7_75t_L g1150 ( 
.A(n_958),
.Y(n_1150)
);

BUFx8_ASAP7_75t_SL g1151 ( 
.A(n_806),
.Y(n_1151)
);

NAND2xp5_ASAP7_75t_L g1152 ( 
.A(n_824),
.B(n_736),
.Y(n_1152)
);

NOR2xp33_ASAP7_75t_L g1153 ( 
.A(n_1081),
.B(n_736),
.Y(n_1153)
);

INVx2_ASAP7_75t_L g1154 ( 
.A(n_958),
.Y(n_1154)
);

INVx5_ASAP7_75t_L g1155 ( 
.A(n_1060),
.Y(n_1155)
);

AND2x6_ASAP7_75t_L g1156 ( 
.A(n_1060),
.B(n_742),
.Y(n_1156)
);

NAND2xp5_ASAP7_75t_L g1157 ( 
.A(n_1081),
.B(n_742),
.Y(n_1157)
);

INVx3_ASAP7_75t_L g1158 ( 
.A(n_1072),
.Y(n_1158)
);

CKINVDCx5p33_ASAP7_75t_R g1159 ( 
.A(n_924),
.Y(n_1159)
);

INVx3_ASAP7_75t_L g1160 ( 
.A(n_1072),
.Y(n_1160)
);

INVx1_ASAP7_75t_L g1161 ( 
.A(n_972),
.Y(n_1161)
);

INVx5_ASAP7_75t_L g1162 ( 
.A(n_1081),
.Y(n_1162)
);

INVx4_ASAP7_75t_L g1163 ( 
.A(n_919),
.Y(n_1163)
);

INVx1_ASAP7_75t_L g1164 ( 
.A(n_974),
.Y(n_1164)
);

INVx1_ASAP7_75t_L g1165 ( 
.A(n_978),
.Y(n_1165)
);

INVx3_ASAP7_75t_L g1166 ( 
.A(n_859),
.Y(n_1166)
);

AND2x4_ASAP7_75t_L g1167 ( 
.A(n_838),
.B(n_749),
.Y(n_1167)
);

NAND2xp5_ASAP7_75t_L g1168 ( 
.A(n_1052),
.B(n_919),
.Y(n_1168)
);

BUFx3_ASAP7_75t_L g1169 ( 
.A(n_799),
.Y(n_1169)
);

NAND2xp5_ASAP7_75t_L g1170 ( 
.A(n_958),
.B(n_749),
.Y(n_1170)
);

INVx5_ASAP7_75t_L g1171 ( 
.A(n_859),
.Y(n_1171)
);

AND2x4_ASAP7_75t_L g1172 ( 
.A(n_833),
.B(n_779),
.Y(n_1172)
);

INVx2_ASAP7_75t_L g1173 ( 
.A(n_894),
.Y(n_1173)
);

INVx4_ASAP7_75t_L g1174 ( 
.A(n_811),
.Y(n_1174)
);

INVx1_ASAP7_75t_L g1175 ( 
.A(n_980),
.Y(n_1175)
);

NAND2xp5_ASAP7_75t_L g1176 ( 
.A(n_896),
.B(n_779),
.Y(n_1176)
);

BUFx6f_ASAP7_75t_L g1177 ( 
.A(n_894),
.Y(n_1177)
);

AND2x2_ASAP7_75t_L g1178 ( 
.A(n_881),
.B(n_663),
.Y(n_1178)
);

AND2x2_ASAP7_75t_L g1179 ( 
.A(n_881),
.B(n_724),
.Y(n_1179)
);

AND2x4_ASAP7_75t_L g1180 ( 
.A(n_836),
.B(n_783),
.Y(n_1180)
);

INVx1_ASAP7_75t_L g1181 ( 
.A(n_981),
.Y(n_1181)
);

INVx1_ASAP7_75t_L g1182 ( 
.A(n_982),
.Y(n_1182)
);

AND2x6_ASAP7_75t_L g1183 ( 
.A(n_996),
.B(n_783),
.Y(n_1183)
);

AND2x2_ASAP7_75t_L g1184 ( 
.A(n_922),
.B(n_940),
.Y(n_1184)
);

AND2x4_ASAP7_75t_L g1185 ( 
.A(n_869),
.B(n_471),
.Y(n_1185)
);

NAND2xp5_ASAP7_75t_L g1186 ( 
.A(n_953),
.B(n_526),
.Y(n_1186)
);

INVx3_ASAP7_75t_L g1187 ( 
.A(n_913),
.Y(n_1187)
);

BUFx3_ASAP7_75t_L g1188 ( 
.A(n_808),
.Y(n_1188)
);

NAND2xp5_ASAP7_75t_L g1189 ( 
.A(n_971),
.B(n_634),
.Y(n_1189)
);

CKINVDCx5p33_ASAP7_75t_R g1190 ( 
.A(n_942),
.Y(n_1190)
);

BUFx6f_ASAP7_75t_L g1191 ( 
.A(n_913),
.Y(n_1191)
);

INVx3_ASAP7_75t_L g1192 ( 
.A(n_945),
.Y(n_1192)
);

NOR2xp33_ASAP7_75t_SL g1193 ( 
.A(n_856),
.B(n_696),
.Y(n_1193)
);

INVx5_ASAP7_75t_L g1194 ( 
.A(n_945),
.Y(n_1194)
);

INVx1_ASAP7_75t_L g1195 ( 
.A(n_841),
.Y(n_1195)
);

INVx5_ASAP7_75t_L g1196 ( 
.A(n_947),
.Y(n_1196)
);

INVx2_ASAP7_75t_L g1197 ( 
.A(n_964),
.Y(n_1197)
);

NAND2xp5_ASAP7_75t_L g1198 ( 
.A(n_1044),
.B(n_504),
.Y(n_1198)
);

AND2x2_ASAP7_75t_L g1199 ( 
.A(n_922),
.B(n_760),
.Y(n_1199)
);

AND2x2_ASAP7_75t_L g1200 ( 
.A(n_940),
.B(n_790),
.Y(n_1200)
);

INVx5_ASAP7_75t_L g1201 ( 
.A(n_964),
.Y(n_1201)
);

AND2x4_ASAP7_75t_L g1202 ( 
.A(n_870),
.B(n_504),
.Y(n_1202)
);

HB1xp67_ASAP7_75t_L g1203 ( 
.A(n_829),
.Y(n_1203)
);

BUFx2_ASAP7_75t_L g1204 ( 
.A(n_1086),
.Y(n_1204)
);

INVx2_ASAP7_75t_L g1205 ( 
.A(n_979),
.Y(n_1205)
);

AND2x4_ASAP7_75t_L g1206 ( 
.A(n_928),
.B(n_661),
.Y(n_1206)
);

INVx1_ASAP7_75t_L g1207 ( 
.A(n_843),
.Y(n_1207)
);

NOR2xp33_ASAP7_75t_L g1208 ( 
.A(n_839),
.B(n_756),
.Y(n_1208)
);

NAND2xp5_ASAP7_75t_L g1209 ( 
.A(n_809),
.B(n_661),
.Y(n_1209)
);

BUFx8_ASAP7_75t_L g1210 ( 
.A(n_979),
.Y(n_1210)
);

AND2x4_ASAP7_75t_L g1211 ( 
.A(n_959),
.B(n_800),
.Y(n_1211)
);

NAND2xp5_ASAP7_75t_SL g1212 ( 
.A(n_814),
.B(n_462),
.Y(n_1212)
);

NOR2xp33_ASAP7_75t_L g1213 ( 
.A(n_829),
.B(n_462),
.Y(n_1213)
);

AND2x4_ASAP7_75t_L g1214 ( 
.A(n_993),
.B(n_497),
.Y(n_1214)
);

INVx2_ASAP7_75t_L g1215 ( 
.A(n_995),
.Y(n_1215)
);

AND2x4_ASAP7_75t_L g1216 ( 
.A(n_999),
.B(n_497),
.Y(n_1216)
);

INVx5_ASAP7_75t_L g1217 ( 
.A(n_995),
.Y(n_1217)
);

AND2x2_ASAP7_75t_L g1218 ( 
.A(n_968),
.B(n_508),
.Y(n_1218)
);

INVx1_ASAP7_75t_L g1219 ( 
.A(n_844),
.Y(n_1219)
);

BUFx6f_ASAP7_75t_L g1220 ( 
.A(n_1005),
.Y(n_1220)
);

BUFx6f_ASAP7_75t_L g1221 ( 
.A(n_1005),
.Y(n_1221)
);

AND2x4_ASAP7_75t_L g1222 ( 
.A(n_811),
.B(n_738),
.Y(n_1222)
);

BUFx6f_ASAP7_75t_L g1223 ( 
.A(n_1019),
.Y(n_1223)
);

BUFx8_ASAP7_75t_SL g1224 ( 
.A(n_816),
.Y(n_1224)
);

INVx5_ASAP7_75t_L g1225 ( 
.A(n_1019),
.Y(n_1225)
);

NAND2xp5_ASAP7_75t_L g1226 ( 
.A(n_810),
.B(n_738),
.Y(n_1226)
);

NAND2xp5_ASAP7_75t_L g1227 ( 
.A(n_813),
.B(n_776),
.Y(n_1227)
);

BUFx3_ASAP7_75t_L g1228 ( 
.A(n_817),
.Y(n_1228)
);

INVx2_ASAP7_75t_L g1229 ( 
.A(n_1031),
.Y(n_1229)
);

AND2x4_ASAP7_75t_L g1230 ( 
.A(n_1000),
.B(n_776),
.Y(n_1230)
);

INVx5_ASAP7_75t_L g1231 ( 
.A(n_1031),
.Y(n_1231)
);

NAND2xp5_ASAP7_75t_L g1232 ( 
.A(n_818),
.B(n_788),
.Y(n_1232)
);

INVx5_ASAP7_75t_L g1233 ( 
.A(n_1062),
.Y(n_1233)
);

INVx2_ASAP7_75t_L g1234 ( 
.A(n_1062),
.Y(n_1234)
);

INVx5_ASAP7_75t_L g1235 ( 
.A(n_1063),
.Y(n_1235)
);

AND2x4_ASAP7_75t_L g1236 ( 
.A(n_1001),
.B(n_788),
.Y(n_1236)
);

NAND2xp5_ASAP7_75t_L g1237 ( 
.A(n_819),
.B(n_588),
.Y(n_1237)
);

HB1xp67_ASAP7_75t_L g1238 ( 
.A(n_835),
.Y(n_1238)
);

BUFx12f_ASAP7_75t_L g1239 ( 
.A(n_942),
.Y(n_1239)
);

BUFx2_ASAP7_75t_L g1240 ( 
.A(n_1086),
.Y(n_1240)
);

NOR2xp33_ASAP7_75t_L g1241 ( 
.A(n_835),
.B(n_429),
.Y(n_1241)
);

XNOR2xp5_ASAP7_75t_L g1242 ( 
.A(n_816),
.B(n_721),
.Y(n_1242)
);

INVx1_ASAP7_75t_L g1243 ( 
.A(n_847),
.Y(n_1243)
);

BUFx3_ASAP7_75t_L g1244 ( 
.A(n_820),
.Y(n_1244)
);

INVx2_ASAP7_75t_SL g1245 ( 
.A(n_840),
.Y(n_1245)
);

INVx5_ASAP7_75t_L g1246 ( 
.A(n_1063),
.Y(n_1246)
);

INVx4_ASAP7_75t_L g1247 ( 
.A(n_840),
.Y(n_1247)
);

AND2x4_ASAP7_75t_L g1248 ( 
.A(n_1003),
.B(n_510),
.Y(n_1248)
);

NAND2xp5_ASAP7_75t_L g1249 ( 
.A(n_822),
.B(n_440),
.Y(n_1249)
);

NAND2xp5_ASAP7_75t_L g1250 ( 
.A(n_823),
.B(n_444),
.Y(n_1250)
);

NAND2xp5_ASAP7_75t_L g1251 ( 
.A(n_827),
.B(n_454),
.Y(n_1251)
);

INVx5_ASAP7_75t_L g1252 ( 
.A(n_862),
.Y(n_1252)
);

HB1xp67_ASAP7_75t_L g1253 ( 
.A(n_805),
.Y(n_1253)
);

BUFx2_ASAP7_75t_L g1254 ( 
.A(n_943),
.Y(n_1254)
);

INVx2_ASAP7_75t_SL g1255 ( 
.A(n_882),
.Y(n_1255)
);

NAND2xp5_ASAP7_75t_L g1256 ( 
.A(n_828),
.B(n_455),
.Y(n_1256)
);

NOR2xp33_ASAP7_75t_L g1257 ( 
.A(n_968),
.B(n_456),
.Y(n_1257)
);

BUFx8_ASAP7_75t_L g1258 ( 
.A(n_1006),
.Y(n_1258)
);

BUFx6f_ASAP7_75t_L g1259 ( 
.A(n_984),
.Y(n_1259)
);

AND2x4_ASAP7_75t_L g1260 ( 
.A(n_1009),
.B(n_511),
.Y(n_1260)
);

NAND2xp5_ASAP7_75t_L g1261 ( 
.A(n_830),
.B(n_461),
.Y(n_1261)
);

BUFx3_ASAP7_75t_L g1262 ( 
.A(n_1085),
.Y(n_1262)
);

NAND2xp5_ASAP7_75t_L g1263 ( 
.A(n_976),
.B(n_465),
.Y(n_1263)
);

NAND2xp5_ASAP7_75t_L g1264 ( 
.A(n_987),
.B(n_475),
.Y(n_1264)
);

BUFx12f_ASAP7_75t_L g1265 ( 
.A(n_943),
.Y(n_1265)
);

INVx1_ASAP7_75t_L g1266 ( 
.A(n_848),
.Y(n_1266)
);

NOR2xp33_ASAP7_75t_L g1267 ( 
.A(n_973),
.B(n_476),
.Y(n_1267)
);

BUFx6f_ASAP7_75t_L g1268 ( 
.A(n_986),
.Y(n_1268)
);

INVx4_ASAP7_75t_L g1269 ( 
.A(n_925),
.Y(n_1269)
);

INVx1_ASAP7_75t_L g1270 ( 
.A(n_1109),
.Y(n_1270)
);

HB1xp67_ASAP7_75t_L g1271 ( 
.A(n_1203),
.Y(n_1271)
);

INVx2_ASAP7_75t_L g1272 ( 
.A(n_1093),
.Y(n_1272)
);

INVx1_ASAP7_75t_L g1273 ( 
.A(n_1173),
.Y(n_1273)
);

INVx2_ASAP7_75t_L g1274 ( 
.A(n_1093),
.Y(n_1274)
);

AND2x6_ASAP7_75t_L g1275 ( 
.A(n_1184),
.B(n_426),
.Y(n_1275)
);

BUFx6f_ASAP7_75t_L g1276 ( 
.A(n_1177),
.Y(n_1276)
);

INVx1_ASAP7_75t_L g1277 ( 
.A(n_1173),
.Y(n_1277)
);

INVx2_ASAP7_75t_L g1278 ( 
.A(n_1099),
.Y(n_1278)
);

BUFx6f_ASAP7_75t_L g1279 ( 
.A(n_1177),
.Y(n_1279)
);

INVx2_ASAP7_75t_L g1280 ( 
.A(n_1099),
.Y(n_1280)
);

INVx2_ASAP7_75t_L g1281 ( 
.A(n_1100),
.Y(n_1281)
);

BUFx6f_ASAP7_75t_L g1282 ( 
.A(n_1177),
.Y(n_1282)
);

INVx1_ASAP7_75t_L g1283 ( 
.A(n_1109),
.Y(n_1283)
);

INVx1_ASAP7_75t_L g1284 ( 
.A(n_1137),
.Y(n_1284)
);

INVx1_ASAP7_75t_L g1285 ( 
.A(n_1137),
.Y(n_1285)
);

INVx1_ASAP7_75t_L g1286 ( 
.A(n_1169),
.Y(n_1286)
);

OR2x6_ASAP7_75t_L g1287 ( 
.A(n_1146),
.B(n_867),
.Y(n_1287)
);

AND2x2_ASAP7_75t_L g1288 ( 
.A(n_1178),
.B(n_973),
.Y(n_1288)
);

INVx1_ASAP7_75t_L g1289 ( 
.A(n_1169),
.Y(n_1289)
);

BUFx6f_ASAP7_75t_L g1290 ( 
.A(n_1177),
.Y(n_1290)
);

NAND2xp5_ASAP7_75t_L g1291 ( 
.A(n_1257),
.B(n_1010),
.Y(n_1291)
);

INVx1_ASAP7_75t_L g1292 ( 
.A(n_1188),
.Y(n_1292)
);

INVx1_ASAP7_75t_L g1293 ( 
.A(n_1188),
.Y(n_1293)
);

NAND2x1_ASAP7_75t_L g1294 ( 
.A(n_1156),
.B(n_633),
.Y(n_1294)
);

INVx1_ASAP7_75t_L g1295 ( 
.A(n_1228),
.Y(n_1295)
);

INVx1_ASAP7_75t_L g1296 ( 
.A(n_1228),
.Y(n_1296)
);

AND2x4_ASAP7_75t_L g1297 ( 
.A(n_1089),
.B(n_851),
.Y(n_1297)
);

AND2x4_ASAP7_75t_L g1298 ( 
.A(n_1089),
.B(n_879),
.Y(n_1298)
);

AND2x6_ASAP7_75t_L g1299 ( 
.A(n_1116),
.B(n_426),
.Y(n_1299)
);

NAND2xp5_ASAP7_75t_SL g1300 ( 
.A(n_1096),
.B(n_1117),
.Y(n_1300)
);

INVx3_ASAP7_75t_L g1301 ( 
.A(n_1191),
.Y(n_1301)
);

INVx1_ASAP7_75t_L g1302 ( 
.A(n_1244),
.Y(n_1302)
);

INVx1_ASAP7_75t_L g1303 ( 
.A(n_1244),
.Y(n_1303)
);

INVx3_ASAP7_75t_L g1304 ( 
.A(n_1191),
.Y(n_1304)
);

INVx1_ASAP7_75t_L g1305 ( 
.A(n_1197),
.Y(n_1305)
);

AND2x4_ASAP7_75t_L g1306 ( 
.A(n_1087),
.B(n_1097),
.Y(n_1306)
);

AND2x2_ASAP7_75t_L g1307 ( 
.A(n_1179),
.B(n_988),
.Y(n_1307)
);

INVx3_ASAP7_75t_L g1308 ( 
.A(n_1191),
.Y(n_1308)
);

BUFx6f_ASAP7_75t_L g1309 ( 
.A(n_1191),
.Y(n_1309)
);

NOR2xp33_ASAP7_75t_L g1310 ( 
.A(n_1168),
.B(n_842),
.Y(n_1310)
);

NAND2xp5_ASAP7_75t_L g1311 ( 
.A(n_1257),
.B(n_1011),
.Y(n_1311)
);

NOR2x1_ASAP7_75t_L g1312 ( 
.A(n_1174),
.B(n_1012),
.Y(n_1312)
);

INVx1_ASAP7_75t_L g1313 ( 
.A(n_1197),
.Y(n_1313)
);

CKINVDCx8_ASAP7_75t_R g1314 ( 
.A(n_1140),
.Y(n_1314)
);

AND2x2_ASAP7_75t_L g1315 ( 
.A(n_1199),
.B(n_988),
.Y(n_1315)
);

BUFx6f_ASAP7_75t_L g1316 ( 
.A(n_1220),
.Y(n_1316)
);

AND2x2_ASAP7_75t_SL g1317 ( 
.A(n_1090),
.B(n_937),
.Y(n_1317)
);

INVx1_ASAP7_75t_L g1318 ( 
.A(n_1205),
.Y(n_1318)
);

INVx1_ASAP7_75t_L g1319 ( 
.A(n_1205),
.Y(n_1319)
);

AND2x2_ASAP7_75t_L g1320 ( 
.A(n_1200),
.B(n_804),
.Y(n_1320)
);

AND2x4_ASAP7_75t_L g1321 ( 
.A(n_1087),
.B(n_1097),
.Y(n_1321)
);

INVx1_ASAP7_75t_L g1322 ( 
.A(n_1215),
.Y(n_1322)
);

INVx1_ASAP7_75t_L g1323 ( 
.A(n_1229),
.Y(n_1323)
);

INVx1_ASAP7_75t_L g1324 ( 
.A(n_1229),
.Y(n_1324)
);

INVx1_ASAP7_75t_L g1325 ( 
.A(n_1234),
.Y(n_1325)
);

NAND2xp5_ASAP7_75t_L g1326 ( 
.A(n_1267),
.B(n_1131),
.Y(n_1326)
);

INVx1_ASAP7_75t_L g1327 ( 
.A(n_1234),
.Y(n_1327)
);

BUFx6f_ASAP7_75t_L g1328 ( 
.A(n_1220),
.Y(n_1328)
);

INVx1_ASAP7_75t_L g1329 ( 
.A(n_1195),
.Y(n_1329)
);

NAND2xp5_ASAP7_75t_L g1330 ( 
.A(n_1267),
.B(n_1013),
.Y(n_1330)
);

INVx3_ASAP7_75t_L g1331 ( 
.A(n_1220),
.Y(n_1331)
);

HB1xp67_ASAP7_75t_L g1332 ( 
.A(n_1203),
.Y(n_1332)
);

INVx1_ASAP7_75t_L g1333 ( 
.A(n_1207),
.Y(n_1333)
);

INVx2_ASAP7_75t_L g1334 ( 
.A(n_1220),
.Y(n_1334)
);

INVx1_ASAP7_75t_L g1335 ( 
.A(n_1219),
.Y(n_1335)
);

CKINVDCx5p33_ASAP7_75t_R g1336 ( 
.A(n_1146),
.Y(n_1336)
);

INVx1_ASAP7_75t_L g1337 ( 
.A(n_1243),
.Y(n_1337)
);

INVx2_ASAP7_75t_L g1338 ( 
.A(n_1221),
.Y(n_1338)
);

INVx3_ASAP7_75t_L g1339 ( 
.A(n_1221),
.Y(n_1339)
);

INVx2_ASAP7_75t_L g1340 ( 
.A(n_1221),
.Y(n_1340)
);

NOR2xp33_ASAP7_75t_L g1341 ( 
.A(n_1101),
.B(n_842),
.Y(n_1341)
);

INVx3_ASAP7_75t_L g1342 ( 
.A(n_1221),
.Y(n_1342)
);

BUFx6f_ASAP7_75t_L g1343 ( 
.A(n_1223),
.Y(n_1343)
);

INVx1_ASAP7_75t_L g1344 ( 
.A(n_1266),
.Y(n_1344)
);

INVx3_ASAP7_75t_L g1345 ( 
.A(n_1223),
.Y(n_1345)
);

BUFx6f_ASAP7_75t_L g1346 ( 
.A(n_1223),
.Y(n_1346)
);

XOR2xp5_ASAP7_75t_L g1347 ( 
.A(n_1242),
.B(n_845),
.Y(n_1347)
);

INVx1_ASAP7_75t_L g1348 ( 
.A(n_1161),
.Y(n_1348)
);

HB1xp67_ASAP7_75t_L g1349 ( 
.A(n_1238),
.Y(n_1349)
);

INVx1_ASAP7_75t_L g1350 ( 
.A(n_1164),
.Y(n_1350)
);

NAND2xp5_ASAP7_75t_SL g1351 ( 
.A(n_1096),
.B(n_846),
.Y(n_1351)
);

INVx1_ASAP7_75t_L g1352 ( 
.A(n_1165),
.Y(n_1352)
);

INVx1_ASAP7_75t_L g1353 ( 
.A(n_1175),
.Y(n_1353)
);

INVx4_ASAP7_75t_L g1354 ( 
.A(n_1142),
.Y(n_1354)
);

NOR2x1_ASAP7_75t_L g1355 ( 
.A(n_1174),
.B(n_1014),
.Y(n_1355)
);

INVx3_ASAP7_75t_L g1356 ( 
.A(n_1223),
.Y(n_1356)
);

INVx1_ASAP7_75t_L g1357 ( 
.A(n_1181),
.Y(n_1357)
);

NAND2xp33_ASAP7_75t_L g1358 ( 
.A(n_1156),
.B(n_628),
.Y(n_1358)
);

INVx2_ASAP7_75t_L g1359 ( 
.A(n_1113),
.Y(n_1359)
);

INVx2_ASAP7_75t_L g1360 ( 
.A(n_1113),
.Y(n_1360)
);

INVx2_ASAP7_75t_L g1361 ( 
.A(n_1138),
.Y(n_1361)
);

INVx1_ASAP7_75t_L g1362 ( 
.A(n_1182),
.Y(n_1362)
);

AND2x2_ASAP7_75t_L g1363 ( 
.A(n_1218),
.B(n_804),
.Y(n_1363)
);

INVx1_ASAP7_75t_L g1364 ( 
.A(n_1088),
.Y(n_1364)
);

INVx1_ASAP7_75t_L g1365 ( 
.A(n_1106),
.Y(n_1365)
);

INVx2_ASAP7_75t_L g1366 ( 
.A(n_1138),
.Y(n_1366)
);

HB1xp67_ASAP7_75t_L g1367 ( 
.A(n_1238),
.Y(n_1367)
);

INVx1_ASAP7_75t_L g1368 ( 
.A(n_1262),
.Y(n_1368)
);

INVx1_ASAP7_75t_L g1369 ( 
.A(n_1262),
.Y(n_1369)
);

INVx1_ASAP7_75t_L g1370 ( 
.A(n_1170),
.Y(n_1370)
);

AND2x2_ASAP7_75t_L g1371 ( 
.A(n_1131),
.B(n_1158),
.Y(n_1371)
);

AND2x2_ASAP7_75t_L g1372 ( 
.A(n_1158),
.B(n_1017),
.Y(n_1372)
);

INVx4_ASAP7_75t_L g1373 ( 
.A(n_1142),
.Y(n_1373)
);

AND2x2_ASAP7_75t_L g1374 ( 
.A(n_1160),
.B(n_1018),
.Y(n_1374)
);

INVx1_ASAP7_75t_L g1375 ( 
.A(n_1166),
.Y(n_1375)
);

INVx1_ASAP7_75t_L g1376 ( 
.A(n_1166),
.Y(n_1376)
);

OAI21x1_ASAP7_75t_L g1377 ( 
.A1(n_1145),
.A2(n_1148),
.B(n_1147),
.Y(n_1377)
);

INVx2_ASAP7_75t_L g1378 ( 
.A(n_1145),
.Y(n_1378)
);

INVx3_ASAP7_75t_L g1379 ( 
.A(n_1103),
.Y(n_1379)
);

INVx2_ASAP7_75t_L g1380 ( 
.A(n_1147),
.Y(n_1380)
);

BUFx6f_ASAP7_75t_L g1381 ( 
.A(n_1259),
.Y(n_1381)
);

INVx1_ASAP7_75t_L g1382 ( 
.A(n_1187),
.Y(n_1382)
);

INVx1_ASAP7_75t_L g1383 ( 
.A(n_1187),
.Y(n_1383)
);

BUFx3_ASAP7_75t_L g1384 ( 
.A(n_1160),
.Y(n_1384)
);

BUFx6f_ASAP7_75t_L g1385 ( 
.A(n_1259),
.Y(n_1385)
);

NAND2xp5_ASAP7_75t_L g1386 ( 
.A(n_1208),
.B(n_1021),
.Y(n_1386)
);

INVx3_ASAP7_75t_L g1387 ( 
.A(n_1103),
.Y(n_1387)
);

BUFx6f_ASAP7_75t_L g1388 ( 
.A(n_1259),
.Y(n_1388)
);

INVx3_ASAP7_75t_L g1389 ( 
.A(n_1103),
.Y(n_1389)
);

OAI22xp5_ASAP7_75t_L g1390 ( 
.A1(n_1090),
.A2(n_805),
.B1(n_873),
.B2(n_846),
.Y(n_1390)
);

NAND2xp5_ASAP7_75t_L g1391 ( 
.A(n_1208),
.B(n_1022),
.Y(n_1391)
);

INVx3_ASAP7_75t_L g1392 ( 
.A(n_1103),
.Y(n_1392)
);

NOR2xp33_ASAP7_75t_SL g1393 ( 
.A(n_1107),
.B(n_950),
.Y(n_1393)
);

INVx1_ASAP7_75t_L g1394 ( 
.A(n_1192),
.Y(n_1394)
);

INVx1_ASAP7_75t_L g1395 ( 
.A(n_1192),
.Y(n_1395)
);

INVx2_ASAP7_75t_L g1396 ( 
.A(n_1149),
.Y(n_1396)
);

INVx3_ASAP7_75t_L g1397 ( 
.A(n_1123),
.Y(n_1397)
);

BUFx6f_ASAP7_75t_L g1398 ( 
.A(n_1259),
.Y(n_1398)
);

OAI22xp5_ASAP7_75t_SL g1399 ( 
.A1(n_1253),
.A2(n_935),
.B1(n_941),
.B2(n_845),
.Y(n_1399)
);

AND2x4_ASAP7_75t_L g1400 ( 
.A(n_1214),
.B(n_899),
.Y(n_1400)
);

BUFx6f_ASAP7_75t_L g1401 ( 
.A(n_1268),
.Y(n_1401)
);

INVx2_ASAP7_75t_L g1402 ( 
.A(n_1150),
.Y(n_1402)
);

INVx4_ASAP7_75t_L g1403 ( 
.A(n_1142),
.Y(n_1403)
);

INVx2_ASAP7_75t_L g1404 ( 
.A(n_1154),
.Y(n_1404)
);

INVx3_ASAP7_75t_L g1405 ( 
.A(n_1123),
.Y(n_1405)
);

INVx1_ASAP7_75t_L g1406 ( 
.A(n_1268),
.Y(n_1406)
);

INVx1_ASAP7_75t_L g1407 ( 
.A(n_1268),
.Y(n_1407)
);

HB1xp67_ASAP7_75t_L g1408 ( 
.A(n_1253),
.Y(n_1408)
);

NAND2xp33_ASAP7_75t_SL g1409 ( 
.A(n_1117),
.B(n_1122),
.Y(n_1409)
);

AND2x2_ASAP7_75t_L g1410 ( 
.A(n_1214),
.B(n_1216),
.Y(n_1410)
);

AND2x2_ASAP7_75t_L g1411 ( 
.A(n_1216),
.B(n_1024),
.Y(n_1411)
);

NAND2xp5_ASAP7_75t_L g1412 ( 
.A(n_1153),
.B(n_1026),
.Y(n_1412)
);

NAND2xp5_ASAP7_75t_L g1413 ( 
.A(n_1153),
.B(n_1029),
.Y(n_1413)
);

INVx1_ASAP7_75t_L g1414 ( 
.A(n_1268),
.Y(n_1414)
);

INVx1_ASAP7_75t_L g1415 ( 
.A(n_1142),
.Y(n_1415)
);

BUFx2_ASAP7_75t_L g1416 ( 
.A(n_1211),
.Y(n_1416)
);

INVx2_ASAP7_75t_L g1417 ( 
.A(n_1154),
.Y(n_1417)
);

AND2x2_ASAP7_75t_L g1418 ( 
.A(n_1230),
.B(n_1030),
.Y(n_1418)
);

INVx2_ASAP7_75t_L g1419 ( 
.A(n_1123),
.Y(n_1419)
);

HB1xp67_ASAP7_75t_L g1420 ( 
.A(n_1254),
.Y(n_1420)
);

NAND2xp5_ASAP7_75t_L g1421 ( 
.A(n_1162),
.B(n_1032),
.Y(n_1421)
);

INVx1_ASAP7_75t_L g1422 ( 
.A(n_1155),
.Y(n_1422)
);

INVx1_ASAP7_75t_L g1423 ( 
.A(n_1226),
.Y(n_1423)
);

INVx1_ASAP7_75t_SL g1424 ( 
.A(n_1288),
.Y(n_1424)
);

NAND2xp5_ASAP7_75t_L g1425 ( 
.A(n_1291),
.B(n_1092),
.Y(n_1425)
);

AOI22xp33_ASAP7_75t_L g1426 ( 
.A1(n_1317),
.A2(n_1212),
.B1(n_1213),
.B2(n_1092),
.Y(n_1426)
);

NAND3xp33_ASAP7_75t_L g1427 ( 
.A(n_1341),
.B(n_1241),
.C(n_1213),
.Y(n_1427)
);

INVx1_ASAP7_75t_L g1428 ( 
.A(n_1273),
.Y(n_1428)
);

BUFx3_ASAP7_75t_L g1429 ( 
.A(n_1306),
.Y(n_1429)
);

INVx3_ASAP7_75t_L g1430 ( 
.A(n_1276),
.Y(n_1430)
);

INVx2_ASAP7_75t_L g1431 ( 
.A(n_1272),
.Y(n_1431)
);

XNOR2xp5_ASAP7_75t_L g1432 ( 
.A(n_1347),
.B(n_1140),
.Y(n_1432)
);

NAND2xp5_ASAP7_75t_L g1433 ( 
.A(n_1311),
.B(n_1241),
.Y(n_1433)
);

INVx4_ASAP7_75t_L g1434 ( 
.A(n_1381),
.Y(n_1434)
);

NOR2xp33_ASAP7_75t_L g1435 ( 
.A(n_1310),
.B(n_1247),
.Y(n_1435)
);

INVx1_ASAP7_75t_L g1436 ( 
.A(n_1273),
.Y(n_1436)
);

NAND2xp5_ASAP7_75t_L g1437 ( 
.A(n_1330),
.B(n_1122),
.Y(n_1437)
);

NAND2xp5_ASAP7_75t_SL g1438 ( 
.A(n_1317),
.B(n_1370),
.Y(n_1438)
);

INVx1_ASAP7_75t_L g1439 ( 
.A(n_1277),
.Y(n_1439)
);

INVx2_ASAP7_75t_SL g1440 ( 
.A(n_1288),
.Y(n_1440)
);

INVx2_ASAP7_75t_L g1441 ( 
.A(n_1272),
.Y(n_1441)
);

INVx1_ASAP7_75t_L g1442 ( 
.A(n_1277),
.Y(n_1442)
);

INVx1_ASAP7_75t_L g1443 ( 
.A(n_1305),
.Y(n_1443)
);

AOI22xp33_ASAP7_75t_L g1444 ( 
.A1(n_1410),
.A2(n_1212),
.B1(n_1183),
.B2(n_1248),
.Y(n_1444)
);

INVx1_ASAP7_75t_L g1445 ( 
.A(n_1305),
.Y(n_1445)
);

INVx1_ASAP7_75t_L g1446 ( 
.A(n_1313),
.Y(n_1446)
);

INVx2_ASAP7_75t_L g1447 ( 
.A(n_1274),
.Y(n_1447)
);

OAI22xp5_ASAP7_75t_L g1448 ( 
.A1(n_1386),
.A2(n_1391),
.B1(n_1326),
.B2(n_1412),
.Y(n_1448)
);

NOR2x1p5_ASAP7_75t_L g1449 ( 
.A(n_1336),
.B(n_1269),
.Y(n_1449)
);

NOR2xp33_ASAP7_75t_L g1450 ( 
.A(n_1390),
.B(n_1247),
.Y(n_1450)
);

NAND2xp5_ASAP7_75t_SL g1451 ( 
.A(n_1370),
.B(n_1141),
.Y(n_1451)
);

BUFx3_ASAP7_75t_L g1452 ( 
.A(n_1306),
.Y(n_1452)
);

NAND2xp5_ASAP7_75t_SL g1453 ( 
.A(n_1413),
.B(n_1141),
.Y(n_1453)
);

OAI22xp33_ASAP7_75t_L g1454 ( 
.A1(n_1416),
.A2(n_1114),
.B1(n_1193),
.B2(n_1157),
.Y(n_1454)
);

INVx3_ASAP7_75t_L g1455 ( 
.A(n_1276),
.Y(n_1455)
);

INVx2_ASAP7_75t_L g1456 ( 
.A(n_1278),
.Y(n_1456)
);

INVx2_ASAP7_75t_SL g1457 ( 
.A(n_1307),
.Y(n_1457)
);

INVx4_ASAP7_75t_L g1458 ( 
.A(n_1381),
.Y(n_1458)
);

INVx2_ASAP7_75t_L g1459 ( 
.A(n_1280),
.Y(n_1459)
);

NAND2xp5_ASAP7_75t_L g1460 ( 
.A(n_1423),
.B(n_1371),
.Y(n_1460)
);

INVx1_ASAP7_75t_L g1461 ( 
.A(n_1313),
.Y(n_1461)
);

INVx1_ASAP7_75t_L g1462 ( 
.A(n_1318),
.Y(n_1462)
);

INVx2_ASAP7_75t_L g1463 ( 
.A(n_1280),
.Y(n_1463)
);

INVx1_ASAP7_75t_L g1464 ( 
.A(n_1318),
.Y(n_1464)
);

NAND3xp33_ASAP7_75t_L g1465 ( 
.A(n_1271),
.B(n_1163),
.C(n_1245),
.Y(n_1465)
);

INVx1_ASAP7_75t_L g1466 ( 
.A(n_1319),
.Y(n_1466)
);

INVx2_ASAP7_75t_L g1467 ( 
.A(n_1281),
.Y(n_1467)
);

INVx1_ASAP7_75t_L g1468 ( 
.A(n_1319),
.Y(n_1468)
);

BUFx6f_ASAP7_75t_L g1469 ( 
.A(n_1276),
.Y(n_1469)
);

NOR2xp33_ASAP7_75t_L g1470 ( 
.A(n_1416),
.B(n_1163),
.Y(n_1470)
);

NOR2xp33_ASAP7_75t_L g1471 ( 
.A(n_1408),
.B(n_1204),
.Y(n_1471)
);

NAND2xp5_ASAP7_75t_L g1472 ( 
.A(n_1371),
.B(n_1120),
.Y(n_1472)
);

NAND2xp5_ASAP7_75t_L g1473 ( 
.A(n_1372),
.B(n_1120),
.Y(n_1473)
);

NAND2xp5_ASAP7_75t_SL g1474 ( 
.A(n_1409),
.B(n_1162),
.Y(n_1474)
);

INVx2_ASAP7_75t_L g1475 ( 
.A(n_1281),
.Y(n_1475)
);

NOR2xp33_ASAP7_75t_L g1476 ( 
.A(n_1351),
.B(n_1240),
.Y(n_1476)
);

BUFx3_ASAP7_75t_L g1477 ( 
.A(n_1306),
.Y(n_1477)
);

INVx4_ASAP7_75t_L g1478 ( 
.A(n_1381),
.Y(n_1478)
);

INVx3_ASAP7_75t_L g1479 ( 
.A(n_1276),
.Y(n_1479)
);

NAND2xp5_ASAP7_75t_SL g1480 ( 
.A(n_1409),
.B(n_1162),
.Y(n_1480)
);

INVx3_ASAP7_75t_L g1481 ( 
.A(n_1276),
.Y(n_1481)
);

AND2x2_ASAP7_75t_L g1482 ( 
.A(n_1307),
.B(n_1315),
.Y(n_1482)
);

NAND2xp5_ASAP7_75t_SL g1483 ( 
.A(n_1321),
.B(n_1162),
.Y(n_1483)
);

AND2x2_ASAP7_75t_L g1484 ( 
.A(n_1315),
.B(n_1211),
.Y(n_1484)
);

INVx3_ASAP7_75t_L g1485 ( 
.A(n_1279),
.Y(n_1485)
);

NAND2xp5_ASAP7_75t_L g1486 ( 
.A(n_1372),
.B(n_1104),
.Y(n_1486)
);

NAND2xp5_ASAP7_75t_SL g1487 ( 
.A(n_1321),
.B(n_1248),
.Y(n_1487)
);

NOR2xp33_ASAP7_75t_L g1488 ( 
.A(n_1320),
.B(n_1269),
.Y(n_1488)
);

INVx1_ASAP7_75t_L g1489 ( 
.A(n_1322),
.Y(n_1489)
);

INVxp67_ASAP7_75t_SL g1490 ( 
.A(n_1384),
.Y(n_1490)
);

NAND2xp5_ASAP7_75t_SL g1491 ( 
.A(n_1321),
.B(n_1260),
.Y(n_1491)
);

AND2x2_ASAP7_75t_L g1492 ( 
.A(n_1320),
.B(n_901),
.Y(n_1492)
);

NAND2xp5_ASAP7_75t_SL g1493 ( 
.A(n_1363),
.B(n_1260),
.Y(n_1493)
);

NAND2xp5_ASAP7_75t_L g1494 ( 
.A(n_1374),
.B(n_1104),
.Y(n_1494)
);

NAND2xp33_ASAP7_75t_L g1495 ( 
.A(n_1312),
.B(n_1156),
.Y(n_1495)
);

NOR2xp33_ASAP7_75t_L g1496 ( 
.A(n_1332),
.B(n_1255),
.Y(n_1496)
);

INVx1_ASAP7_75t_L g1497 ( 
.A(n_1322),
.Y(n_1497)
);

INVx2_ASAP7_75t_SL g1498 ( 
.A(n_1420),
.Y(n_1498)
);

NAND2xp5_ASAP7_75t_SL g1499 ( 
.A(n_1363),
.B(n_1155),
.Y(n_1499)
);

NOR2xp33_ASAP7_75t_L g1500 ( 
.A(n_1349),
.B(n_873),
.Y(n_1500)
);

INVx1_ASAP7_75t_L g1501 ( 
.A(n_1323),
.Y(n_1501)
);

INVx1_ASAP7_75t_L g1502 ( 
.A(n_1323),
.Y(n_1502)
);

NAND2xp5_ASAP7_75t_L g1503 ( 
.A(n_1374),
.B(n_1118),
.Y(n_1503)
);

BUFx6f_ASAP7_75t_SL g1504 ( 
.A(n_1287),
.Y(n_1504)
);

INVx1_ASAP7_75t_L g1505 ( 
.A(n_1324),
.Y(n_1505)
);

BUFx10_ASAP7_75t_L g1506 ( 
.A(n_1336),
.Y(n_1506)
);

NAND2xp5_ASAP7_75t_SL g1507 ( 
.A(n_1381),
.B(n_1155),
.Y(n_1507)
);

BUFx6f_ASAP7_75t_SL g1508 ( 
.A(n_1287),
.Y(n_1508)
);

NAND2xp5_ASAP7_75t_SL g1509 ( 
.A(n_1381),
.B(n_1155),
.Y(n_1509)
);

INVx1_ASAP7_75t_L g1510 ( 
.A(n_1325),
.Y(n_1510)
);

INVx1_ASAP7_75t_L g1511 ( 
.A(n_1325),
.Y(n_1511)
);

INVx1_ASAP7_75t_L g1512 ( 
.A(n_1327),
.Y(n_1512)
);

INVx1_ASAP7_75t_L g1513 ( 
.A(n_1327),
.Y(n_1513)
);

INVx2_ASAP7_75t_SL g1514 ( 
.A(n_1400),
.Y(n_1514)
);

INVx1_ASAP7_75t_L g1515 ( 
.A(n_1364),
.Y(n_1515)
);

INVx2_ASAP7_75t_L g1516 ( 
.A(n_1377),
.Y(n_1516)
);

INVx1_ASAP7_75t_L g1517 ( 
.A(n_1365),
.Y(n_1517)
);

NAND3xp33_ASAP7_75t_L g1518 ( 
.A(n_1367),
.B(n_1118),
.C(n_1143),
.Y(n_1518)
);

INVx2_ASAP7_75t_L g1519 ( 
.A(n_1377),
.Y(n_1519)
);

NAND2xp5_ASAP7_75t_SL g1520 ( 
.A(n_1385),
.B(n_1252),
.Y(n_1520)
);

NAND2xp5_ASAP7_75t_L g1521 ( 
.A(n_1410),
.B(n_1143),
.Y(n_1521)
);

NAND2xp5_ASAP7_75t_SL g1522 ( 
.A(n_1385),
.B(n_1252),
.Y(n_1522)
);

INVx2_ASAP7_75t_L g1523 ( 
.A(n_1378),
.Y(n_1523)
);

BUFx6f_ASAP7_75t_SL g1524 ( 
.A(n_1287),
.Y(n_1524)
);

INVx1_ASAP7_75t_L g1525 ( 
.A(n_1375),
.Y(n_1525)
);

OR2x2_ASAP7_75t_L g1526 ( 
.A(n_1400),
.B(n_998),
.Y(n_1526)
);

INVx1_ASAP7_75t_L g1527 ( 
.A(n_1376),
.Y(n_1527)
);

AND2x2_ASAP7_75t_L g1528 ( 
.A(n_1400),
.B(n_1121),
.Y(n_1528)
);

INVx4_ASAP7_75t_L g1529 ( 
.A(n_1385),
.Y(n_1529)
);

INVx5_ASAP7_75t_L g1530 ( 
.A(n_1354),
.Y(n_1530)
);

INVx2_ASAP7_75t_L g1531 ( 
.A(n_1378),
.Y(n_1531)
);

NAND2xp5_ASAP7_75t_SL g1532 ( 
.A(n_1385),
.B(n_1252),
.Y(n_1532)
);

BUFx6f_ASAP7_75t_SL g1533 ( 
.A(n_1287),
.Y(n_1533)
);

INVx1_ASAP7_75t_L g1534 ( 
.A(n_1382),
.Y(n_1534)
);

NOR2xp33_ASAP7_75t_L g1535 ( 
.A(n_1384),
.B(n_897),
.Y(n_1535)
);

NAND2xp5_ASAP7_75t_SL g1536 ( 
.A(n_1385),
.B(n_1252),
.Y(n_1536)
);

INVx1_ASAP7_75t_L g1537 ( 
.A(n_1383),
.Y(n_1537)
);

AND2x2_ASAP7_75t_L g1538 ( 
.A(n_1297),
.B(n_1130),
.Y(n_1538)
);

NAND2xp5_ASAP7_75t_SL g1539 ( 
.A(n_1388),
.B(n_1398),
.Y(n_1539)
);

INVx3_ASAP7_75t_L g1540 ( 
.A(n_1279),
.Y(n_1540)
);

NOR2xp33_ASAP7_75t_L g1541 ( 
.A(n_1300),
.B(n_897),
.Y(n_1541)
);

NAND2xp5_ASAP7_75t_SL g1542 ( 
.A(n_1388),
.B(n_1185),
.Y(n_1542)
);

INVx2_ASAP7_75t_L g1543 ( 
.A(n_1380),
.Y(n_1543)
);

INVx2_ASAP7_75t_L g1544 ( 
.A(n_1380),
.Y(n_1544)
);

AND3x2_ASAP7_75t_L g1545 ( 
.A(n_1393),
.B(n_1102),
.C(n_1095),
.Y(n_1545)
);

AND2x2_ASAP7_75t_L g1546 ( 
.A(n_1297),
.B(n_1133),
.Y(n_1546)
);

NAND2xp5_ASAP7_75t_SL g1547 ( 
.A(n_1388),
.B(n_1398),
.Y(n_1547)
);

CKINVDCx5p33_ASAP7_75t_R g1548 ( 
.A(n_1314),
.Y(n_1548)
);

OAI22xp5_ASAP7_75t_L g1549 ( 
.A1(n_1348),
.A2(n_1176),
.B1(n_1202),
.B2(n_1185),
.Y(n_1549)
);

NOR2xp33_ASAP7_75t_L g1550 ( 
.A(n_1368),
.B(n_911),
.Y(n_1550)
);

INVx3_ASAP7_75t_L g1551 ( 
.A(n_1279),
.Y(n_1551)
);

NAND2xp33_ASAP7_75t_SL g1552 ( 
.A(n_1294),
.B(n_1107),
.Y(n_1552)
);

AOI22xp5_ASAP7_75t_L g1553 ( 
.A1(n_1297),
.A2(n_1183),
.B1(n_1206),
.B2(n_1202),
.Y(n_1553)
);

OAI22xp33_ASAP7_75t_L g1554 ( 
.A1(n_1314),
.A2(n_1159),
.B1(n_1190),
.B2(n_1189),
.Y(n_1554)
);

NAND2xp5_ASAP7_75t_L g1555 ( 
.A(n_1411),
.B(n_1198),
.Y(n_1555)
);

INVx1_ASAP7_75t_L g1556 ( 
.A(n_1394),
.Y(n_1556)
);

NAND2xp5_ASAP7_75t_SL g1557 ( 
.A(n_1398),
.B(n_1206),
.Y(n_1557)
);

INVx1_ASAP7_75t_L g1558 ( 
.A(n_1395),
.Y(n_1558)
);

OAI21xp5_ASAP7_75t_L g1559 ( 
.A1(n_1396),
.A2(n_1264),
.B(n_1263),
.Y(n_1559)
);

NAND2xp5_ASAP7_75t_SL g1560 ( 
.A(n_1398),
.B(n_1401),
.Y(n_1560)
);

NAND2xp5_ASAP7_75t_L g1561 ( 
.A(n_1411),
.B(n_1222),
.Y(n_1561)
);

AND2x6_ASAP7_75t_L g1562 ( 
.A(n_1355),
.B(n_1091),
.Y(n_1562)
);

NAND2xp5_ASAP7_75t_L g1563 ( 
.A(n_1329),
.B(n_1222),
.Y(n_1563)
);

INVx2_ASAP7_75t_L g1564 ( 
.A(n_1523),
.Y(n_1564)
);

AND2x2_ASAP7_75t_L g1565 ( 
.A(n_1492),
.B(n_1015),
.Y(n_1565)
);

XOR2xp5_ASAP7_75t_L g1566 ( 
.A(n_1432),
.B(n_1347),
.Y(n_1566)
);

XNOR2xp5_ASAP7_75t_L g1567 ( 
.A(n_1545),
.B(n_1399),
.Y(n_1567)
);

INVx1_ASAP7_75t_L g1568 ( 
.A(n_1515),
.Y(n_1568)
);

INVx1_ASAP7_75t_L g1569 ( 
.A(n_1517),
.Y(n_1569)
);

INVx1_ASAP7_75t_L g1570 ( 
.A(n_1428),
.Y(n_1570)
);

INVxp33_ASAP7_75t_L g1571 ( 
.A(n_1526),
.Y(n_1571)
);

AND2x2_ASAP7_75t_L g1572 ( 
.A(n_1484),
.B(n_1058),
.Y(n_1572)
);

NOR2xp33_ASAP7_75t_L g1573 ( 
.A(n_1433),
.B(n_1298),
.Y(n_1573)
);

NOR2xp33_ASAP7_75t_L g1574 ( 
.A(n_1425),
.B(n_1298),
.Y(n_1574)
);

OR2x6_ASAP7_75t_L g1575 ( 
.A(n_1514),
.B(n_1239),
.Y(n_1575)
);

INVx1_ASAP7_75t_L g1576 ( 
.A(n_1436),
.Y(n_1576)
);

INVx1_ASAP7_75t_L g1577 ( 
.A(n_1439),
.Y(n_1577)
);

AND2x2_ASAP7_75t_L g1578 ( 
.A(n_1528),
.B(n_970),
.Y(n_1578)
);

AND2x2_ASAP7_75t_L g1579 ( 
.A(n_1538),
.B(n_970),
.Y(n_1579)
);

XNOR2xp5_ASAP7_75t_L g1580 ( 
.A(n_1548),
.B(n_935),
.Y(n_1580)
);

XOR2xp5_ASAP7_75t_L g1581 ( 
.A(n_1548),
.B(n_941),
.Y(n_1581)
);

NAND2xp33_ASAP7_75t_R g1582 ( 
.A(n_1450),
.B(n_1159),
.Y(n_1582)
);

AND2x2_ASAP7_75t_L g1583 ( 
.A(n_1546),
.B(n_975),
.Y(n_1583)
);

NOR2xp33_ASAP7_75t_L g1584 ( 
.A(n_1438),
.B(n_1298),
.Y(n_1584)
);

INVx1_ASAP7_75t_L g1585 ( 
.A(n_1442),
.Y(n_1585)
);

XOR2x2_ASAP7_75t_L g1586 ( 
.A(n_1427),
.B(n_1095),
.Y(n_1586)
);

NOR2xp33_ASAP7_75t_L g1587 ( 
.A(n_1438),
.B(n_1369),
.Y(n_1587)
);

INVx1_ASAP7_75t_L g1588 ( 
.A(n_1443),
.Y(n_1588)
);

XOR2xp5_ASAP7_75t_L g1589 ( 
.A(n_1554),
.B(n_989),
.Y(n_1589)
);

INVx1_ASAP7_75t_L g1590 ( 
.A(n_1445),
.Y(n_1590)
);

OAI21xp5_ASAP7_75t_L g1591 ( 
.A1(n_1448),
.A2(n_1404),
.B(n_1402),
.Y(n_1591)
);

INVx1_ASAP7_75t_L g1592 ( 
.A(n_1446),
.Y(n_1592)
);

AND2x2_ASAP7_75t_L g1593 ( 
.A(n_1424),
.B(n_975),
.Y(n_1593)
);

INVx1_ASAP7_75t_L g1594 ( 
.A(n_1461),
.Y(n_1594)
);

NOR2xp33_ASAP7_75t_L g1595 ( 
.A(n_1435),
.B(n_1286),
.Y(n_1595)
);

INVx1_ASAP7_75t_L g1596 ( 
.A(n_1462),
.Y(n_1596)
);

INVx1_ASAP7_75t_L g1597 ( 
.A(n_1464),
.Y(n_1597)
);

INVx1_ASAP7_75t_L g1598 ( 
.A(n_1466),
.Y(n_1598)
);

INVx1_ASAP7_75t_L g1599 ( 
.A(n_1468),
.Y(n_1599)
);

NOR2xp33_ASAP7_75t_L g1600 ( 
.A(n_1437),
.B(n_1289),
.Y(n_1600)
);

AND2x2_ASAP7_75t_SL g1601 ( 
.A(n_1426),
.B(n_1358),
.Y(n_1601)
);

CKINVDCx20_ASAP7_75t_R g1602 ( 
.A(n_1506),
.Y(n_1602)
);

INVx1_ASAP7_75t_L g1603 ( 
.A(n_1489),
.Y(n_1603)
);

AND2x2_ASAP7_75t_SL g1604 ( 
.A(n_1434),
.B(n_1358),
.Y(n_1604)
);

INVxp67_ASAP7_75t_L g1605 ( 
.A(n_1498),
.Y(n_1605)
);

INVx1_ASAP7_75t_L g1606 ( 
.A(n_1497),
.Y(n_1606)
);

INVx1_ASAP7_75t_L g1607 ( 
.A(n_1501),
.Y(n_1607)
);

INVx1_ASAP7_75t_L g1608 ( 
.A(n_1502),
.Y(n_1608)
);

NAND2xp5_ASAP7_75t_L g1609 ( 
.A(n_1486),
.B(n_1418),
.Y(n_1609)
);

AND2x2_ASAP7_75t_L g1610 ( 
.A(n_1482),
.B(n_985),
.Y(n_1610)
);

AND2x2_ASAP7_75t_L g1611 ( 
.A(n_1471),
.B(n_985),
.Y(n_1611)
);

NOR2xp33_ASAP7_75t_L g1612 ( 
.A(n_1494),
.B(n_1292),
.Y(n_1612)
);

INVx1_ASAP7_75t_L g1613 ( 
.A(n_1505),
.Y(n_1613)
);

INVx1_ASAP7_75t_L g1614 ( 
.A(n_1510),
.Y(n_1614)
);

NOR2xp33_ASAP7_75t_L g1615 ( 
.A(n_1503),
.B(n_1488),
.Y(n_1615)
);

XOR2xp5_ASAP7_75t_L g1616 ( 
.A(n_1465),
.B(n_997),
.Y(n_1616)
);

INVx2_ASAP7_75t_L g1617 ( 
.A(n_1523),
.Y(n_1617)
);

INVx2_ASAP7_75t_L g1618 ( 
.A(n_1531),
.Y(n_1618)
);

INVxp67_ASAP7_75t_SL g1619 ( 
.A(n_1469),
.Y(n_1619)
);

OAI21xp5_ASAP7_75t_L g1620 ( 
.A1(n_1559),
.A2(n_1417),
.B(n_1404),
.Y(n_1620)
);

XOR2xp5_ASAP7_75t_L g1621 ( 
.A(n_1518),
.B(n_997),
.Y(n_1621)
);

INVx1_ASAP7_75t_L g1622 ( 
.A(n_1511),
.Y(n_1622)
);

XOR2xp5_ASAP7_75t_L g1623 ( 
.A(n_1553),
.B(n_1023),
.Y(n_1623)
);

INVx1_ASAP7_75t_L g1624 ( 
.A(n_1512),
.Y(n_1624)
);

INVx1_ASAP7_75t_L g1625 ( 
.A(n_1513),
.Y(n_1625)
);

CKINVDCx20_ASAP7_75t_R g1626 ( 
.A(n_1506),
.Y(n_1626)
);

NAND2xp5_ASAP7_75t_L g1627 ( 
.A(n_1473),
.B(n_1418),
.Y(n_1627)
);

INVxp67_ASAP7_75t_L g1628 ( 
.A(n_1561),
.Y(n_1628)
);

NOR2xp33_ASAP7_75t_L g1629 ( 
.A(n_1440),
.B(n_1293),
.Y(n_1629)
);

NOR2xp33_ASAP7_75t_L g1630 ( 
.A(n_1440),
.B(n_1295),
.Y(n_1630)
);

XOR2xp5_ASAP7_75t_L g1631 ( 
.A(n_1549),
.B(n_1023),
.Y(n_1631)
);

INVx1_ASAP7_75t_L g1632 ( 
.A(n_1525),
.Y(n_1632)
);

INVx1_ASAP7_75t_L g1633 ( 
.A(n_1527),
.Y(n_1633)
);

INVx1_ASAP7_75t_L g1634 ( 
.A(n_1534),
.Y(n_1634)
);

INVx1_ASAP7_75t_L g1635 ( 
.A(n_1537),
.Y(n_1635)
);

NAND2xp5_ASAP7_75t_L g1636 ( 
.A(n_1472),
.B(n_1299),
.Y(n_1636)
);

NAND2xp5_ASAP7_75t_L g1637 ( 
.A(n_1521),
.B(n_1299),
.Y(n_1637)
);

HB1xp67_ASAP7_75t_L g1638 ( 
.A(n_1429),
.Y(n_1638)
);

INVx1_ASAP7_75t_L g1639 ( 
.A(n_1556),
.Y(n_1639)
);

INVx1_ASAP7_75t_L g1640 ( 
.A(n_1558),
.Y(n_1640)
);

AND2x2_ASAP7_75t_L g1641 ( 
.A(n_1500),
.B(n_991),
.Y(n_1641)
);

INVx2_ASAP7_75t_L g1642 ( 
.A(n_1531),
.Y(n_1642)
);

INVx1_ASAP7_75t_L g1643 ( 
.A(n_1457),
.Y(n_1643)
);

INVxp33_ASAP7_75t_SL g1644 ( 
.A(n_1470),
.Y(n_1644)
);

AND2x2_ASAP7_75t_L g1645 ( 
.A(n_1496),
.B(n_991),
.Y(n_1645)
);

XOR2xp5_ASAP7_75t_L g1646 ( 
.A(n_1454),
.B(n_1025),
.Y(n_1646)
);

INVx2_ASAP7_75t_L g1647 ( 
.A(n_1543),
.Y(n_1647)
);

NOR2xp33_ASAP7_75t_L g1648 ( 
.A(n_1555),
.B(n_1296),
.Y(n_1648)
);

NOR2xp33_ASAP7_75t_L g1649 ( 
.A(n_1493),
.B(n_1302),
.Y(n_1649)
);

INVx1_ASAP7_75t_L g1650 ( 
.A(n_1460),
.Y(n_1650)
);

INVx1_ASAP7_75t_L g1651 ( 
.A(n_1431),
.Y(n_1651)
);

INVx2_ASAP7_75t_L g1652 ( 
.A(n_1543),
.Y(n_1652)
);

AND2x2_ASAP7_75t_L g1653 ( 
.A(n_1476),
.B(n_994),
.Y(n_1653)
);

INVxp33_ASAP7_75t_SL g1654 ( 
.A(n_1535),
.Y(n_1654)
);

CKINVDCx20_ASAP7_75t_R g1655 ( 
.A(n_1506),
.Y(n_1655)
);

INVx4_ASAP7_75t_SL g1656 ( 
.A(n_1504),
.Y(n_1656)
);

INVx1_ASAP7_75t_L g1657 ( 
.A(n_1431),
.Y(n_1657)
);

INVx1_ASAP7_75t_L g1658 ( 
.A(n_1441),
.Y(n_1658)
);

INVx1_ASAP7_75t_L g1659 ( 
.A(n_1441),
.Y(n_1659)
);

INVx1_ASAP7_75t_L g1660 ( 
.A(n_1447),
.Y(n_1660)
);

INVx1_ASAP7_75t_L g1661 ( 
.A(n_1447),
.Y(n_1661)
);

NAND2xp5_ASAP7_75t_SL g1662 ( 
.A(n_1469),
.B(n_1417),
.Y(n_1662)
);

NOR2xp33_ASAP7_75t_L g1663 ( 
.A(n_1493),
.B(n_1303),
.Y(n_1663)
);

INVx1_ASAP7_75t_L g1664 ( 
.A(n_1456),
.Y(n_1664)
);

INVx2_ASAP7_75t_L g1665 ( 
.A(n_1544),
.Y(n_1665)
);

XNOR2xp5_ASAP7_75t_L g1666 ( 
.A(n_1449),
.B(n_989),
.Y(n_1666)
);

CKINVDCx20_ASAP7_75t_R g1667 ( 
.A(n_1552),
.Y(n_1667)
);

AND2x2_ASAP7_75t_L g1668 ( 
.A(n_1563),
.B(n_994),
.Y(n_1668)
);

INVx1_ASAP7_75t_L g1669 ( 
.A(n_1459),
.Y(n_1669)
);

INVxp67_ASAP7_75t_SL g1670 ( 
.A(n_1469),
.Y(n_1670)
);

BUFx2_ASAP7_75t_L g1671 ( 
.A(n_1429),
.Y(n_1671)
);

CKINVDCx16_ASAP7_75t_R g1672 ( 
.A(n_1504),
.Y(n_1672)
);

AND2x6_ASAP7_75t_L g1673 ( 
.A(n_1452),
.B(n_1415),
.Y(n_1673)
);

BUFx4f_ASAP7_75t_L g1674 ( 
.A(n_1562),
.Y(n_1674)
);

NAND2xp5_ASAP7_75t_L g1675 ( 
.A(n_1444),
.B(n_1299),
.Y(n_1675)
);

INVx1_ASAP7_75t_L g1676 ( 
.A(n_1459),
.Y(n_1676)
);

CKINVDCx20_ASAP7_75t_R g1677 ( 
.A(n_1552),
.Y(n_1677)
);

INVx1_ASAP7_75t_L g1678 ( 
.A(n_1463),
.Y(n_1678)
);

INVx1_ASAP7_75t_L g1679 ( 
.A(n_1467),
.Y(n_1679)
);

CKINVDCx20_ASAP7_75t_R g1680 ( 
.A(n_1452),
.Y(n_1680)
);

NAND2xp5_ASAP7_75t_L g1681 ( 
.A(n_1562),
.B(n_1542),
.Y(n_1681)
);

INVx1_ASAP7_75t_L g1682 ( 
.A(n_1467),
.Y(n_1682)
);

INVx1_ASAP7_75t_L g1683 ( 
.A(n_1475),
.Y(n_1683)
);

A2O1A1Ixp33_ASAP7_75t_L g1684 ( 
.A1(n_1615),
.A2(n_1550),
.B(n_1541),
.C(n_1451),
.Y(n_1684)
);

INVx2_ASAP7_75t_L g1685 ( 
.A(n_1564),
.Y(n_1685)
);

INVx1_ASAP7_75t_L g1686 ( 
.A(n_1568),
.Y(n_1686)
);

BUFx3_ASAP7_75t_L g1687 ( 
.A(n_1626),
.Y(n_1687)
);

INVx2_ASAP7_75t_L g1688 ( 
.A(n_1617),
.Y(n_1688)
);

NOR2xp33_ASAP7_75t_L g1689 ( 
.A(n_1654),
.B(n_1487),
.Y(n_1689)
);

NAND3xp33_ASAP7_75t_L g1690 ( 
.A(n_1582),
.B(n_1190),
.C(n_1051),
.Y(n_1690)
);

NOR2xp33_ASAP7_75t_L g1691 ( 
.A(n_1644),
.B(n_1487),
.Y(n_1691)
);

NAND2xp33_ASAP7_75t_L g1692 ( 
.A(n_1650),
.B(n_1474),
.Y(n_1692)
);

NAND2xp5_ASAP7_75t_L g1693 ( 
.A(n_1615),
.B(n_1574),
.Y(n_1693)
);

NOR2xp33_ASAP7_75t_L g1694 ( 
.A(n_1573),
.B(n_1491),
.Y(n_1694)
);

NOR2xp33_ASAP7_75t_L g1695 ( 
.A(n_1573),
.B(n_1491),
.Y(n_1695)
);

AOI22xp33_ASAP7_75t_L g1696 ( 
.A1(n_1574),
.A2(n_1299),
.B1(n_1557),
.B2(n_1542),
.Y(n_1696)
);

AND2x6_ASAP7_75t_SL g1697 ( 
.A(n_1575),
.B(n_1111),
.Y(n_1697)
);

AOI22xp33_ASAP7_75t_L g1698 ( 
.A1(n_1601),
.A2(n_1299),
.B1(n_1557),
.B2(n_1167),
.Y(n_1698)
);

INVx2_ASAP7_75t_L g1699 ( 
.A(n_1618),
.Y(n_1699)
);

NAND2xp5_ASAP7_75t_L g1700 ( 
.A(n_1628),
.B(n_1477),
.Y(n_1700)
);

AOI221xp5_ASAP7_75t_L g1701 ( 
.A1(n_1641),
.A2(n_977),
.B1(n_1027),
.B2(n_961),
.C(n_911),
.Y(n_1701)
);

OAI22xp5_ASAP7_75t_SL g1702 ( 
.A1(n_1589),
.A2(n_1049),
.B1(n_1064),
.B2(n_1025),
.Y(n_1702)
);

INVx1_ASAP7_75t_L g1703 ( 
.A(n_1569),
.Y(n_1703)
);

BUFx5_ASAP7_75t_L g1704 ( 
.A(n_1673),
.Y(n_1704)
);

OAI221xp5_ASAP7_75t_L g1705 ( 
.A1(n_1582),
.A2(n_1621),
.B1(n_1611),
.B2(n_1645),
.C(n_1609),
.Y(n_1705)
);

INVx2_ASAP7_75t_L g1706 ( 
.A(n_1642),
.Y(n_1706)
);

NAND2xp5_ASAP7_75t_SL g1707 ( 
.A(n_1605),
.B(n_1477),
.Y(n_1707)
);

NOR2xp33_ASAP7_75t_L g1708 ( 
.A(n_1628),
.B(n_1453),
.Y(n_1708)
);

NAND2xp5_ASAP7_75t_L g1709 ( 
.A(n_1627),
.B(n_1045),
.Y(n_1709)
);

BUFx3_ASAP7_75t_L g1710 ( 
.A(n_1655),
.Y(n_1710)
);

NAND2xp5_ASAP7_75t_SL g1711 ( 
.A(n_1605),
.B(n_1045),
.Y(n_1711)
);

NAND2xp5_ASAP7_75t_SL g1712 ( 
.A(n_1668),
.B(n_1051),
.Y(n_1712)
);

NOR2xp33_ASAP7_75t_L g1713 ( 
.A(n_1653),
.B(n_1584),
.Y(n_1713)
);

BUFx3_ASAP7_75t_L g1714 ( 
.A(n_1602),
.Y(n_1714)
);

NAND2xp5_ASAP7_75t_L g1715 ( 
.A(n_1648),
.B(n_1076),
.Y(n_1715)
);

AOI22xp33_ASAP7_75t_L g1716 ( 
.A1(n_1601),
.A2(n_1299),
.B1(n_1167),
.B2(n_1180),
.Y(n_1716)
);

INVx1_ASAP7_75t_L g1717 ( 
.A(n_1632),
.Y(n_1717)
);

NAND2xp5_ASAP7_75t_L g1718 ( 
.A(n_1648),
.B(n_1076),
.Y(n_1718)
);

INVx2_ASAP7_75t_L g1719 ( 
.A(n_1647),
.Y(n_1719)
);

AOI22xp5_ASAP7_75t_L g1720 ( 
.A1(n_1572),
.A2(n_977),
.B1(n_1027),
.B2(n_961),
.Y(n_1720)
);

AOI22xp33_ASAP7_75t_SL g1721 ( 
.A1(n_1565),
.A2(n_1064),
.B1(n_1065),
.B2(n_1049),
.Y(n_1721)
);

INVx3_ASAP7_75t_L g1722 ( 
.A(n_1674),
.Y(n_1722)
);

NOR2xp33_ASAP7_75t_SL g1723 ( 
.A(n_1672),
.B(n_1239),
.Y(n_1723)
);

AND2x2_ASAP7_75t_L g1724 ( 
.A(n_1610),
.B(n_1133),
.Y(n_1724)
);

NAND2xp5_ASAP7_75t_SL g1725 ( 
.A(n_1595),
.B(n_1453),
.Y(n_1725)
);

OR2x2_ASAP7_75t_L g1726 ( 
.A(n_1580),
.B(n_1581),
.Y(n_1726)
);

NOR2xp33_ASAP7_75t_L g1727 ( 
.A(n_1584),
.B(n_1499),
.Y(n_1727)
);

AOI22xp33_ASAP7_75t_L g1728 ( 
.A1(n_1646),
.A2(n_1180),
.B1(n_1172),
.B2(n_1091),
.Y(n_1728)
);

BUFx2_ASAP7_75t_L g1729 ( 
.A(n_1680),
.Y(n_1729)
);

OR2x2_ASAP7_75t_L g1730 ( 
.A(n_1593),
.B(n_957),
.Y(n_1730)
);

NAND2xp5_ASAP7_75t_L g1731 ( 
.A(n_1612),
.B(n_1595),
.Y(n_1731)
);

INVx1_ASAP7_75t_L g1732 ( 
.A(n_1633),
.Y(n_1732)
);

NAND2xp5_ASAP7_75t_L g1733 ( 
.A(n_1612),
.B(n_1562),
.Y(n_1733)
);

NAND2xp5_ASAP7_75t_L g1734 ( 
.A(n_1600),
.B(n_1649),
.Y(n_1734)
);

BUFx5_ASAP7_75t_L g1735 ( 
.A(n_1673),
.Y(n_1735)
);

INVxp67_ASAP7_75t_SL g1736 ( 
.A(n_1619),
.Y(n_1736)
);

INVx1_ASAP7_75t_L g1737 ( 
.A(n_1634),
.Y(n_1737)
);

NAND2xp5_ASAP7_75t_L g1738 ( 
.A(n_1600),
.B(n_1562),
.Y(n_1738)
);

AND2x2_ASAP7_75t_SL g1739 ( 
.A(n_1674),
.B(n_1604),
.Y(n_1739)
);

OAI22xp5_ASAP7_75t_L g1740 ( 
.A1(n_1570),
.A2(n_1490),
.B1(n_1451),
.B2(n_1480),
.Y(n_1740)
);

INVx1_ASAP7_75t_L g1741 ( 
.A(n_1635),
.Y(n_1741)
);

BUFx6f_ASAP7_75t_L g1742 ( 
.A(n_1604),
.Y(n_1742)
);

NAND2xp5_ASAP7_75t_SL g1743 ( 
.A(n_1579),
.B(n_1258),
.Y(n_1743)
);

OR2x2_ASAP7_75t_L g1744 ( 
.A(n_1566),
.B(n_965),
.Y(n_1744)
);

NOR2xp33_ASAP7_75t_L g1745 ( 
.A(n_1578),
.B(n_1499),
.Y(n_1745)
);

AOI22xp5_ASAP7_75t_SL g1746 ( 
.A1(n_1631),
.A2(n_1066),
.B1(n_1068),
.B2(n_1065),
.Y(n_1746)
);

INVx2_ASAP7_75t_L g1747 ( 
.A(n_1652),
.Y(n_1747)
);

NAND2xp5_ASAP7_75t_SL g1748 ( 
.A(n_1583),
.B(n_1258),
.Y(n_1748)
);

INVx2_ASAP7_75t_L g1749 ( 
.A(n_1665),
.Y(n_1749)
);

NAND2xp5_ASAP7_75t_SL g1750 ( 
.A(n_1680),
.B(n_1210),
.Y(n_1750)
);

NAND2xp5_ASAP7_75t_L g1751 ( 
.A(n_1649),
.B(n_1663),
.Y(n_1751)
);

NOR3x1_ASAP7_75t_L g1752 ( 
.A(n_1639),
.B(n_1136),
.C(n_1111),
.Y(n_1752)
);

NAND2xp5_ASAP7_75t_L g1753 ( 
.A(n_1663),
.B(n_1562),
.Y(n_1753)
);

INVx1_ASAP7_75t_L g1754 ( 
.A(n_1640),
.Y(n_1754)
);

NAND2xp5_ASAP7_75t_L g1755 ( 
.A(n_1638),
.B(n_1562),
.Y(n_1755)
);

OAI22xp5_ASAP7_75t_L g1756 ( 
.A1(n_1576),
.A2(n_1480),
.B1(n_1474),
.B2(n_1483),
.Y(n_1756)
);

INVxp67_ASAP7_75t_SL g1757 ( 
.A(n_1619),
.Y(n_1757)
);

AND2x2_ASAP7_75t_L g1758 ( 
.A(n_1724),
.B(n_1689),
.Y(n_1758)
);

AOI22xp5_ASAP7_75t_L g1759 ( 
.A1(n_1713),
.A2(n_1265),
.B1(n_1068),
.B2(n_1066),
.Y(n_1759)
);

NOR2xp33_ASAP7_75t_SL g1760 ( 
.A(n_1723),
.B(n_1136),
.Y(n_1760)
);

NAND2xp5_ASAP7_75t_L g1761 ( 
.A(n_1731),
.B(n_1571),
.Y(n_1761)
);

BUFx2_ASAP7_75t_L g1762 ( 
.A(n_1729),
.Y(n_1762)
);

NAND2xp5_ASAP7_75t_L g1763 ( 
.A(n_1693),
.B(n_1571),
.Y(n_1763)
);

INVx2_ASAP7_75t_SL g1764 ( 
.A(n_1687),
.Y(n_1764)
);

INVx1_ASAP7_75t_SL g1765 ( 
.A(n_1726),
.Y(n_1765)
);

AOI21x1_ASAP7_75t_L g1766 ( 
.A1(n_1725),
.A2(n_1662),
.B(n_1519),
.Y(n_1766)
);

BUFx6f_ASAP7_75t_L g1767 ( 
.A(n_1739),
.Y(n_1767)
);

NAND2xp5_ASAP7_75t_L g1768 ( 
.A(n_1713),
.B(n_1623),
.Y(n_1768)
);

NAND2xp5_ASAP7_75t_L g1769 ( 
.A(n_1715),
.B(n_1629),
.Y(n_1769)
);

NAND2xp5_ASAP7_75t_L g1770 ( 
.A(n_1718),
.B(n_1629),
.Y(n_1770)
);

NAND2xp5_ASAP7_75t_L g1771 ( 
.A(n_1734),
.B(n_1630),
.Y(n_1771)
);

AOI22xp5_ASAP7_75t_L g1772 ( 
.A1(n_1691),
.A2(n_1265),
.B1(n_1616),
.B2(n_1677),
.Y(n_1772)
);

INVx1_ASAP7_75t_L g1773 ( 
.A(n_1686),
.Y(n_1773)
);

NOR2xp33_ASAP7_75t_L g1774 ( 
.A(n_1694),
.B(n_1055),
.Y(n_1774)
);

NAND2xp5_ASAP7_75t_L g1775 ( 
.A(n_1694),
.B(n_1630),
.Y(n_1775)
);

OAI22xp5_ASAP7_75t_L g1776 ( 
.A1(n_1684),
.A2(n_1602),
.B1(n_1677),
.B2(n_1585),
.Y(n_1776)
);

INVx1_ASAP7_75t_L g1777 ( 
.A(n_1703),
.Y(n_1777)
);

NAND2xp5_ASAP7_75t_L g1778 ( 
.A(n_1695),
.B(n_1577),
.Y(n_1778)
);

NAND2xp5_ASAP7_75t_SL g1779 ( 
.A(n_1751),
.B(n_1587),
.Y(n_1779)
);

OAI21xp5_ASAP7_75t_L g1780 ( 
.A1(n_1695),
.A2(n_1637),
.B(n_1636),
.Y(n_1780)
);

AOI33xp33_ASAP7_75t_L g1781 ( 
.A1(n_1701),
.A2(n_992),
.A3(n_854),
.B1(n_850),
.B2(n_857),
.B3(n_853),
.Y(n_1781)
);

OAI321xp33_ASAP7_75t_L g1782 ( 
.A1(n_1705),
.A2(n_1575),
.A3(n_967),
.B1(n_931),
.B2(n_954),
.C(n_902),
.Y(n_1782)
);

INVx2_ASAP7_75t_L g1783 ( 
.A(n_1685),
.Y(n_1783)
);

AND2x4_ASAP7_75t_L g1784 ( 
.A(n_1722),
.B(n_1656),
.Y(n_1784)
);

AOI21xp5_ASAP7_75t_L g1785 ( 
.A1(n_1692),
.A2(n_1591),
.B(n_1670),
.Y(n_1785)
);

OAI21xp5_ASAP7_75t_L g1786 ( 
.A1(n_1708),
.A2(n_1587),
.B(n_1662),
.Y(n_1786)
);

AOI22xp5_ASAP7_75t_L g1787 ( 
.A1(n_1691),
.A2(n_1666),
.B1(n_1667),
.B2(n_1586),
.Y(n_1787)
);

NAND2xp5_ASAP7_75t_L g1788 ( 
.A(n_1689),
.B(n_1588),
.Y(n_1788)
);

NAND2xp5_ASAP7_75t_L g1789 ( 
.A(n_1709),
.B(n_1590),
.Y(n_1789)
);

BUFx6f_ASAP7_75t_L g1790 ( 
.A(n_1739),
.Y(n_1790)
);

NAND2xp5_ASAP7_75t_L g1791 ( 
.A(n_1728),
.B(n_1592),
.Y(n_1791)
);

AOI21xp5_ASAP7_75t_L g1792 ( 
.A1(n_1736),
.A2(n_1670),
.B(n_1519),
.Y(n_1792)
);

A2O1A1Ixp33_ASAP7_75t_L g1793 ( 
.A1(n_1727),
.A2(n_960),
.B(n_1596),
.C(n_1594),
.Y(n_1793)
);

NAND2xp5_ASAP7_75t_SL g1794 ( 
.A(n_1738),
.B(n_1681),
.Y(n_1794)
);

INVx2_ASAP7_75t_SL g1795 ( 
.A(n_1710),
.Y(n_1795)
);

OAI21xp5_ASAP7_75t_L g1796 ( 
.A1(n_1708),
.A2(n_1733),
.B(n_1727),
.Y(n_1796)
);

BUFx6f_ASAP7_75t_L g1797 ( 
.A(n_1742),
.Y(n_1797)
);

BUFx12f_ASAP7_75t_L g1798 ( 
.A(n_1697),
.Y(n_1798)
);

NAND2xp5_ASAP7_75t_L g1799 ( 
.A(n_1728),
.B(n_1597),
.Y(n_1799)
);

NAND2xp5_ASAP7_75t_L g1800 ( 
.A(n_1745),
.B(n_1598),
.Y(n_1800)
);

NAND2xp5_ASAP7_75t_L g1801 ( 
.A(n_1745),
.B(n_1599),
.Y(n_1801)
);

NAND2xp5_ASAP7_75t_L g1802 ( 
.A(n_1720),
.B(n_1603),
.Y(n_1802)
);

AOI21x1_ASAP7_75t_L g1803 ( 
.A1(n_1756),
.A2(n_1516),
.B(n_1539),
.Y(n_1803)
);

NOR2xp33_ASAP7_75t_L g1804 ( 
.A(n_1730),
.B(n_1055),
.Y(n_1804)
);

AOI21xp5_ASAP7_75t_L g1805 ( 
.A1(n_1736),
.A2(n_1516),
.B(n_1620),
.Y(n_1805)
);

NAND2xp5_ASAP7_75t_SL g1806 ( 
.A(n_1742),
.B(n_1469),
.Y(n_1806)
);

INVx3_ASAP7_75t_SL g1807 ( 
.A(n_1764),
.Y(n_1807)
);

AOI21xp5_ASAP7_75t_L g1808 ( 
.A1(n_1785),
.A2(n_1757),
.B(n_1740),
.Y(n_1808)
);

NAND2xp5_ASAP7_75t_SL g1809 ( 
.A(n_1775),
.B(n_1742),
.Y(n_1809)
);

HB1xp67_ASAP7_75t_L g1810 ( 
.A(n_1766),
.Y(n_1810)
);

NAND2xp5_ASAP7_75t_L g1811 ( 
.A(n_1761),
.B(n_1717),
.Y(n_1811)
);

AO32x2_ASAP7_75t_L g1812 ( 
.A1(n_1776),
.A2(n_1702),
.A3(n_1478),
.B1(n_1529),
.B2(n_1458),
.Y(n_1812)
);

NAND2xp5_ASAP7_75t_L g1813 ( 
.A(n_1763),
.B(n_1732),
.Y(n_1813)
);

BUFx6f_ASAP7_75t_L g1814 ( 
.A(n_1797),
.Y(n_1814)
);

OAI22xp5_ASAP7_75t_L g1815 ( 
.A1(n_1774),
.A2(n_1771),
.B1(n_1802),
.B2(n_1770),
.Y(n_1815)
);

INVx3_ASAP7_75t_L g1816 ( 
.A(n_1767),
.Y(n_1816)
);

NOR2xp33_ASAP7_75t_L g1817 ( 
.A(n_1774),
.B(n_1804),
.Y(n_1817)
);

OAI22xp5_ASAP7_75t_L g1818 ( 
.A1(n_1769),
.A2(n_1690),
.B1(n_1716),
.B2(n_1698),
.Y(n_1818)
);

AOI21xp5_ASAP7_75t_L g1819 ( 
.A1(n_1805),
.A2(n_1757),
.B(n_1753),
.Y(n_1819)
);

AOI21xp5_ASAP7_75t_L g1820 ( 
.A1(n_1792),
.A2(n_1742),
.B(n_1547),
.Y(n_1820)
);

AOI21xp5_ASAP7_75t_L g1821 ( 
.A1(n_1779),
.A2(n_1547),
.B(n_1539),
.Y(n_1821)
);

INVx1_ASAP7_75t_L g1822 ( 
.A(n_1773),
.Y(n_1822)
);

NAND2xp5_ASAP7_75t_SL g1823 ( 
.A(n_1796),
.B(n_1704),
.Y(n_1823)
);

NAND2xp5_ASAP7_75t_L g1824 ( 
.A(n_1788),
.B(n_1737),
.Y(n_1824)
);

NAND2xp5_ASAP7_75t_L g1825 ( 
.A(n_1778),
.B(n_1758),
.Y(n_1825)
);

NOR2xp33_ASAP7_75t_L g1826 ( 
.A(n_1804),
.B(n_1151),
.Y(n_1826)
);

AOI21xp5_ASAP7_75t_L g1827 ( 
.A1(n_1793),
.A2(n_1560),
.B(n_1696),
.Y(n_1827)
);

AND2x2_ASAP7_75t_L g1828 ( 
.A(n_1768),
.B(n_1714),
.Y(n_1828)
);

NAND2xp5_ASAP7_75t_L g1829 ( 
.A(n_1800),
.B(n_1741),
.Y(n_1829)
);

NAND2xp5_ASAP7_75t_L g1830 ( 
.A(n_1801),
.B(n_1754),
.Y(n_1830)
);

INVx2_ASAP7_75t_L g1831 ( 
.A(n_1783),
.Y(n_1831)
);

NOR2xp33_ASAP7_75t_L g1832 ( 
.A(n_1795),
.B(n_1151),
.Y(n_1832)
);

NAND2xp5_ASAP7_75t_L g1833 ( 
.A(n_1789),
.B(n_1700),
.Y(n_1833)
);

INVx4_ASAP7_75t_L g1834 ( 
.A(n_1797),
.Y(n_1834)
);

AOI21x1_ASAP7_75t_L g1835 ( 
.A1(n_1803),
.A2(n_1755),
.B(n_1522),
.Y(n_1835)
);

INVx2_ASAP7_75t_L g1836 ( 
.A(n_1777),
.Y(n_1836)
);

AOI21xp5_ASAP7_75t_L g1837 ( 
.A1(n_1793),
.A2(n_1698),
.B(n_1716),
.Y(n_1837)
);

AOI22xp33_ASAP7_75t_L g1838 ( 
.A1(n_1791),
.A2(n_1224),
.B1(n_1721),
.B2(n_1748),
.Y(n_1838)
);

NOR2xp33_ASAP7_75t_L g1839 ( 
.A(n_1787),
.B(n_1224),
.Y(n_1839)
);

AND2x4_ASAP7_75t_L g1840 ( 
.A(n_1784),
.B(n_1656),
.Y(n_1840)
);

BUFx3_ASAP7_75t_L g1841 ( 
.A(n_1762),
.Y(n_1841)
);

AOI21x1_ASAP7_75t_L g1842 ( 
.A1(n_1806),
.A2(n_1794),
.B(n_1799),
.Y(n_1842)
);

AOI21xp5_ASAP7_75t_L g1843 ( 
.A1(n_1786),
.A2(n_1675),
.B(n_1455),
.Y(n_1843)
);

HB1xp67_ASAP7_75t_L g1844 ( 
.A(n_1794),
.Y(n_1844)
);

OR2x6_ASAP7_75t_SL g1845 ( 
.A(n_1760),
.B(n_1744),
.Y(n_1845)
);

OAI22xp5_ASAP7_75t_L g1846 ( 
.A1(n_1772),
.A2(n_1606),
.B1(n_1608),
.B2(n_1607),
.Y(n_1846)
);

AOI21xp5_ASAP7_75t_L g1847 ( 
.A1(n_1780),
.A2(n_1455),
.B(n_1430),
.Y(n_1847)
);

NAND2xp5_ASAP7_75t_L g1848 ( 
.A(n_1765),
.B(n_1613),
.Y(n_1848)
);

NOR2xp33_ASAP7_75t_L g1849 ( 
.A(n_1782),
.B(n_1712),
.Y(n_1849)
);

AOI22xp33_ASAP7_75t_L g1850 ( 
.A1(n_1759),
.A2(n_1743),
.B1(n_741),
.B2(n_769),
.Y(n_1850)
);

NOR2xp33_ASAP7_75t_R g1851 ( 
.A(n_1798),
.B(n_1504),
.Y(n_1851)
);

A2O1A1Ixp33_ASAP7_75t_L g1852 ( 
.A1(n_1781),
.A2(n_1622),
.B(n_1624),
.C(n_1614),
.Y(n_1852)
);

NAND3xp33_ASAP7_75t_SL g1853 ( 
.A(n_1806),
.B(n_777),
.C(n_740),
.Y(n_1853)
);

NOR2xp33_ASAP7_75t_SL g1854 ( 
.A(n_1815),
.B(n_1767),
.Y(n_1854)
);

A2O1A1Ixp33_ASAP7_75t_L g1855 ( 
.A1(n_1817),
.A2(n_1750),
.B(n_1746),
.C(n_1112),
.Y(n_1855)
);

AND2x2_ASAP7_75t_L g1856 ( 
.A(n_1825),
.B(n_1797),
.Y(n_1856)
);

BUFx2_ASAP7_75t_L g1857 ( 
.A(n_1841),
.Y(n_1857)
);

OAI21x1_ASAP7_75t_L g1858 ( 
.A1(n_1808),
.A2(n_1835),
.B(n_1819),
.Y(n_1858)
);

A2O1A1Ixp33_ASAP7_75t_L g1859 ( 
.A1(n_1817),
.A2(n_1112),
.B(n_1124),
.C(n_1110),
.Y(n_1859)
);

OAI21xp5_ASAP7_75t_L g1860 ( 
.A1(n_1837),
.A2(n_1707),
.B(n_1035),
.Y(n_1860)
);

AOI21x1_ASAP7_75t_L g1861 ( 
.A1(n_1810),
.A2(n_1827),
.B(n_1842),
.Y(n_1861)
);

INVxp67_ASAP7_75t_L g1862 ( 
.A(n_1848),
.Y(n_1862)
);

OAI21x1_ASAP7_75t_L g1863 ( 
.A1(n_1820),
.A2(n_1722),
.B(n_1455),
.Y(n_1863)
);

OAI21x1_ASAP7_75t_L g1864 ( 
.A1(n_1843),
.A2(n_1479),
.B(n_1430),
.Y(n_1864)
);

CKINVDCx20_ASAP7_75t_R g1865 ( 
.A(n_1851),
.Y(n_1865)
);

INVx1_ASAP7_75t_L g1866 ( 
.A(n_1822),
.Y(n_1866)
);

AOI21xp5_ASAP7_75t_L g1867 ( 
.A1(n_1823),
.A2(n_1790),
.B(n_1767),
.Y(n_1867)
);

A2O1A1Ixp33_ASAP7_75t_L g1868 ( 
.A1(n_1849),
.A2(n_1124),
.B(n_1132),
.C(n_1110),
.Y(n_1868)
);

BUFx6f_ASAP7_75t_L g1869 ( 
.A(n_1814),
.Y(n_1869)
);

NOR2xp33_ASAP7_75t_L g1870 ( 
.A(n_1826),
.B(n_1056),
.Y(n_1870)
);

OA22x2_ASAP7_75t_L g1871 ( 
.A1(n_1846),
.A2(n_1575),
.B1(n_1567),
.B2(n_1784),
.Y(n_1871)
);

AND3x4_ASAP7_75t_L g1872 ( 
.A(n_1840),
.B(n_1752),
.C(n_1172),
.Y(n_1872)
);

INVxp67_ASAP7_75t_L g1873 ( 
.A(n_1828),
.Y(n_1873)
);

OAI21x1_ASAP7_75t_L g1874 ( 
.A1(n_1821),
.A2(n_1481),
.B(n_1479),
.Y(n_1874)
);

NAND3x1_ASAP7_75t_L g1875 ( 
.A(n_1839),
.B(n_858),
.C(n_849),
.Y(n_1875)
);

A2O1A1Ixp33_ASAP7_75t_L g1876 ( 
.A1(n_1849),
.A2(n_1818),
.B(n_1838),
.C(n_1853),
.Y(n_1876)
);

OAI21x1_ASAP7_75t_L g1877 ( 
.A1(n_1847),
.A2(n_1485),
.B(n_1481),
.Y(n_1877)
);

NAND2xp5_ASAP7_75t_L g1878 ( 
.A(n_1824),
.B(n_1797),
.Y(n_1878)
);

OAI21xp33_ASAP7_75t_L g1879 ( 
.A1(n_1850),
.A2(n_1074),
.B(n_1056),
.Y(n_1879)
);

AOI21xp5_ASAP7_75t_L g1880 ( 
.A1(n_1809),
.A2(n_1790),
.B(n_1767),
.Y(n_1880)
);

AOI21xp5_ASAP7_75t_L g1881 ( 
.A1(n_1829),
.A2(n_1790),
.B(n_1495),
.Y(n_1881)
);

AO31x2_ASAP7_75t_L g1882 ( 
.A1(n_1831),
.A2(n_1699),
.A3(n_1706),
.B(n_1688),
.Y(n_1882)
);

NAND2xp5_ASAP7_75t_L g1883 ( 
.A(n_1833),
.B(n_1790),
.Y(n_1883)
);

NAND2xp5_ASAP7_75t_L g1884 ( 
.A(n_1830),
.B(n_1811),
.Y(n_1884)
);

NAND2xp5_ASAP7_75t_L g1885 ( 
.A(n_1813),
.B(n_1625),
.Y(n_1885)
);

AOI21x1_ASAP7_75t_L g1886 ( 
.A1(n_1810),
.A2(n_1037),
.B(n_1033),
.Y(n_1886)
);

OAI22xp5_ASAP7_75t_L g1887 ( 
.A1(n_1838),
.A2(n_1638),
.B1(n_1711),
.B2(n_1671),
.Y(n_1887)
);

OAI21xp5_ASAP7_75t_L g1888 ( 
.A1(n_1852),
.A2(n_1039),
.B(n_1038),
.Y(n_1888)
);

OR2x2_ASAP7_75t_L g1889 ( 
.A(n_1836),
.B(n_1132),
.Y(n_1889)
);

OAI22xp5_ASAP7_75t_L g1890 ( 
.A1(n_1850),
.A2(n_519),
.B1(n_522),
.B2(n_514),
.Y(n_1890)
);

BUFx5_ASAP7_75t_L g1891 ( 
.A(n_1840),
.Y(n_1891)
);

NAND2xp5_ASAP7_75t_L g1892 ( 
.A(n_1844),
.B(n_1040),
.Y(n_1892)
);

AND2x4_ASAP7_75t_L g1893 ( 
.A(n_1816),
.B(n_1656),
.Y(n_1893)
);

AOI21xp5_ASAP7_75t_L g1894 ( 
.A1(n_1844),
.A2(n_1522),
.B(n_1520),
.Y(n_1894)
);

NAND2xp5_ASAP7_75t_L g1895 ( 
.A(n_1807),
.B(n_1041),
.Y(n_1895)
);

OAI22xp5_ASAP7_75t_L g1896 ( 
.A1(n_1807),
.A2(n_1074),
.B1(n_1524),
.B2(n_1508),
.Y(n_1896)
);

NAND2xp5_ASAP7_75t_L g1897 ( 
.A(n_1814),
.B(n_1042),
.Y(n_1897)
);

AOI221x1_ASAP7_75t_L g1898 ( 
.A1(n_1834),
.A2(n_1047),
.B1(n_1048),
.B2(n_1046),
.C(n_1043),
.Y(n_1898)
);

INVx1_ASAP7_75t_L g1899 ( 
.A(n_1812),
.Y(n_1899)
);

BUFx3_ASAP7_75t_L g1900 ( 
.A(n_1845),
.Y(n_1900)
);

NAND2xp5_ASAP7_75t_L g1901 ( 
.A(n_1814),
.B(n_1834),
.Y(n_1901)
);

INVx2_ASAP7_75t_SL g1902 ( 
.A(n_1814),
.Y(n_1902)
);

AOI21xp5_ASAP7_75t_L g1903 ( 
.A1(n_1812),
.A2(n_1536),
.B(n_1532),
.Y(n_1903)
);

NOR2xp33_ASAP7_75t_L g1904 ( 
.A(n_1832),
.B(n_1128),
.Y(n_1904)
);

NAND2xp5_ASAP7_75t_L g1905 ( 
.A(n_1812),
.B(n_1050),
.Y(n_1905)
);

OAI21x1_ASAP7_75t_L g1906 ( 
.A1(n_1812),
.A2(n_1540),
.B(n_1485),
.Y(n_1906)
);

INVx2_ASAP7_75t_L g1907 ( 
.A(n_1836),
.Y(n_1907)
);

INVx2_ASAP7_75t_SL g1908 ( 
.A(n_1807),
.Y(n_1908)
);

OAI21x1_ASAP7_75t_L g1909 ( 
.A1(n_1808),
.A2(n_1551),
.B(n_1540),
.Y(n_1909)
);

INVx1_ASAP7_75t_L g1910 ( 
.A(n_1822),
.Y(n_1910)
);

NAND2xp5_ASAP7_75t_L g1911 ( 
.A(n_1815),
.B(n_1053),
.Y(n_1911)
);

AOI21xp33_ASAP7_75t_L g1912 ( 
.A1(n_1849),
.A2(n_1747),
.B(n_1719),
.Y(n_1912)
);

INVx2_ASAP7_75t_L g1913 ( 
.A(n_1836),
.Y(n_1913)
);

BUFx6f_ASAP7_75t_L g1914 ( 
.A(n_1814),
.Y(n_1914)
);

NAND2xp5_ASAP7_75t_L g1915 ( 
.A(n_1815),
.B(n_1054),
.Y(n_1915)
);

BUFx2_ASAP7_75t_SL g1916 ( 
.A(n_1865),
.Y(n_1916)
);

INVx1_ASAP7_75t_L g1917 ( 
.A(n_1866),
.Y(n_1917)
);

BUFx3_ASAP7_75t_L g1918 ( 
.A(n_1857),
.Y(n_1918)
);

AOI222xp33_ASAP7_75t_L g1919 ( 
.A1(n_1879),
.A2(n_1524),
.B1(n_1533),
.B2(n_1508),
.C1(n_550),
.C2(n_543),
.Y(n_1919)
);

NAND2xp5_ASAP7_75t_L g1920 ( 
.A(n_1884),
.B(n_1059),
.Y(n_1920)
);

INVx1_ASAP7_75t_L g1921 ( 
.A(n_1910),
.Y(n_1921)
);

INVx1_ASAP7_75t_L g1922 ( 
.A(n_1907),
.Y(n_1922)
);

INVx3_ASAP7_75t_L g1923 ( 
.A(n_1869),
.Y(n_1923)
);

NAND2xp5_ASAP7_75t_L g1924 ( 
.A(n_1905),
.B(n_1061),
.Y(n_1924)
);

A2O1A1Ixp33_ASAP7_75t_L g1925 ( 
.A1(n_1876),
.A2(n_1079),
.B(n_1067),
.C(n_1070),
.Y(n_1925)
);

AOI22xp33_ASAP7_75t_L g1926 ( 
.A1(n_1871),
.A2(n_1128),
.B1(n_1749),
.B2(n_1524),
.Y(n_1926)
);

AND2x4_ASAP7_75t_L g1927 ( 
.A(n_1908),
.B(n_1643),
.Y(n_1927)
);

BUFx6f_ASAP7_75t_L g1928 ( 
.A(n_1869),
.Y(n_1928)
);

INVx1_ASAP7_75t_L g1929 ( 
.A(n_1913),
.Y(n_1929)
);

AND2x4_ASAP7_75t_L g1930 ( 
.A(n_1856),
.B(n_860),
.Y(n_1930)
);

NOR2xp33_ASAP7_75t_L g1931 ( 
.A(n_1870),
.B(n_6),
.Y(n_1931)
);

O2A1O1Ixp5_ASAP7_75t_L g1932 ( 
.A1(n_1911),
.A2(n_861),
.B(n_864),
.C(n_863),
.Y(n_1932)
);

BUFx3_ASAP7_75t_L g1933 ( 
.A(n_1900),
.Y(n_1933)
);

OAI22xp5_ASAP7_75t_L g1934 ( 
.A1(n_1915),
.A2(n_545),
.B1(n_556),
.B2(n_528),
.Y(n_1934)
);

NAND2xp5_ASAP7_75t_L g1935 ( 
.A(n_1899),
.B(n_1069),
.Y(n_1935)
);

A2O1A1Ixp33_ASAP7_75t_L g1936 ( 
.A1(n_1855),
.A2(n_1071),
.B(n_1075),
.C(n_1073),
.Y(n_1936)
);

INVx2_ASAP7_75t_SL g1937 ( 
.A(n_1869),
.Y(n_1937)
);

BUFx3_ASAP7_75t_L g1938 ( 
.A(n_1872),
.Y(n_1938)
);

A2O1A1Ixp33_ASAP7_75t_SL g1939 ( 
.A1(n_1904),
.A2(n_865),
.B(n_868),
.C(n_866),
.Y(n_1939)
);

AND2x2_ASAP7_75t_L g1940 ( 
.A(n_1873),
.B(n_1077),
.Y(n_1940)
);

INVx3_ASAP7_75t_L g1941 ( 
.A(n_1914),
.Y(n_1941)
);

NOR2xp33_ASAP7_75t_L g1942 ( 
.A(n_1895),
.B(n_6),
.Y(n_1942)
);

INVxp67_ASAP7_75t_SL g1943 ( 
.A(n_1861),
.Y(n_1943)
);

INVx1_ASAP7_75t_L g1944 ( 
.A(n_1862),
.Y(n_1944)
);

BUFx2_ASAP7_75t_L g1945 ( 
.A(n_1901),
.Y(n_1945)
);

AOI21x1_ASAP7_75t_L g1946 ( 
.A1(n_1892),
.A2(n_872),
.B(n_871),
.Y(n_1946)
);

INVx2_ASAP7_75t_SL g1947 ( 
.A(n_1914),
.Y(n_1947)
);

INVx5_ASAP7_75t_L g1948 ( 
.A(n_1914),
.Y(n_1948)
);

INVx2_ASAP7_75t_L g1949 ( 
.A(n_1882),
.Y(n_1949)
);

INVx2_ASAP7_75t_L g1950 ( 
.A(n_1882),
.Y(n_1950)
);

NAND2xp5_ASAP7_75t_L g1951 ( 
.A(n_1878),
.B(n_1885),
.Y(n_1951)
);

A2O1A1Ixp33_ASAP7_75t_L g1952 ( 
.A1(n_1879),
.A2(n_1080),
.B(n_1083),
.C(n_558),
.Y(n_1952)
);

BUFx10_ASAP7_75t_L g1953 ( 
.A(n_1902),
.Y(n_1953)
);

INVx1_ASAP7_75t_L g1954 ( 
.A(n_1883),
.Y(n_1954)
);

NAND2xp5_ASAP7_75t_SL g1955 ( 
.A(n_1891),
.B(n_1704),
.Y(n_1955)
);

NAND2xp5_ASAP7_75t_L g1956 ( 
.A(n_1903),
.B(n_874),
.Y(n_1956)
);

OA21x2_ASAP7_75t_L g1957 ( 
.A1(n_1858),
.A2(n_877),
.B(n_875),
.Y(n_1957)
);

INVx2_ASAP7_75t_L g1958 ( 
.A(n_1882),
.Y(n_1958)
);

NAND2xp5_ASAP7_75t_L g1959 ( 
.A(n_1881),
.B(n_878),
.Y(n_1959)
);

NAND2xp5_ASAP7_75t_L g1960 ( 
.A(n_1860),
.B(n_880),
.Y(n_1960)
);

HB1xp67_ASAP7_75t_L g1961 ( 
.A(n_1897),
.Y(n_1961)
);

INVx1_ASAP7_75t_L g1962 ( 
.A(n_1889),
.Y(n_1962)
);

INVx1_ASAP7_75t_L g1963 ( 
.A(n_1886),
.Y(n_1963)
);

AND2x4_ASAP7_75t_L g1964 ( 
.A(n_1893),
.B(n_883),
.Y(n_1964)
);

INVx3_ASAP7_75t_L g1965 ( 
.A(n_1909),
.Y(n_1965)
);

AND2x2_ASAP7_75t_L g1966 ( 
.A(n_1891),
.B(n_884),
.Y(n_1966)
);

NAND2xp5_ASAP7_75t_L g1967 ( 
.A(n_1860),
.B(n_885),
.Y(n_1967)
);

INVx2_ASAP7_75t_L g1968 ( 
.A(n_1906),
.Y(n_1968)
);

AOI22xp33_ASAP7_75t_L g1969 ( 
.A1(n_1912),
.A2(n_1890),
.B1(n_1887),
.B2(n_1508),
.Y(n_1969)
);

OR2x6_ASAP7_75t_SL g1970 ( 
.A(n_1896),
.B(n_561),
.Y(n_1970)
);

AND2x2_ASAP7_75t_L g1971 ( 
.A(n_1891),
.B(n_887),
.Y(n_1971)
);

AND2x4_ASAP7_75t_L g1972 ( 
.A(n_1893),
.B(n_888),
.Y(n_1972)
);

NOR2xp67_ASAP7_75t_R g1973 ( 
.A(n_1891),
.B(n_889),
.Y(n_1973)
);

NAND2xp5_ASAP7_75t_L g1974 ( 
.A(n_1894),
.B(n_1867),
.Y(n_1974)
);

NAND2xp5_ASAP7_75t_L g1975 ( 
.A(n_1868),
.B(n_890),
.Y(n_1975)
);

INVx2_ASAP7_75t_L g1976 ( 
.A(n_1891),
.Y(n_1976)
);

AOI22xp5_ASAP7_75t_L g1977 ( 
.A1(n_1875),
.A2(n_1533),
.B1(n_1673),
.B2(n_1210),
.Y(n_1977)
);

BUFx6f_ASAP7_75t_L g1978 ( 
.A(n_1863),
.Y(n_1978)
);

AND2x2_ASAP7_75t_L g1979 ( 
.A(n_1880),
.B(n_891),
.Y(n_1979)
);

OAI22xp5_ASAP7_75t_L g1980 ( 
.A1(n_1859),
.A2(n_575),
.B1(n_576),
.B2(n_569),
.Y(n_1980)
);

INVx1_ASAP7_75t_L g1981 ( 
.A(n_1874),
.Y(n_1981)
);

INVx1_ASAP7_75t_L g1982 ( 
.A(n_1864),
.Y(n_1982)
);

AOI21xp5_ASAP7_75t_L g1983 ( 
.A1(n_1898),
.A2(n_1529),
.B(n_1509),
.Y(n_1983)
);

AND2x2_ASAP7_75t_L g1984 ( 
.A(n_1877),
.B(n_892),
.Y(n_1984)
);

CKINVDCx11_ASAP7_75t_R g1985 ( 
.A(n_1890),
.Y(n_1985)
);

INVx1_ASAP7_75t_L g1986 ( 
.A(n_1888),
.Y(n_1986)
);

INVx1_ASAP7_75t_L g1987 ( 
.A(n_1888),
.Y(n_1987)
);

A2O1A1Ixp33_ASAP7_75t_SL g1988 ( 
.A1(n_1870),
.A2(n_895),
.B(n_898),
.C(n_893),
.Y(n_1988)
);

AND2x4_ASAP7_75t_L g1989 ( 
.A(n_1857),
.B(n_900),
.Y(n_1989)
);

AND2x4_ASAP7_75t_L g1990 ( 
.A(n_1857),
.B(n_903),
.Y(n_1990)
);

OR2x6_ASAP7_75t_L g1991 ( 
.A(n_1867),
.B(n_1651),
.Y(n_1991)
);

OAI22xp5_ASAP7_75t_L g1992 ( 
.A1(n_1876),
.A2(n_584),
.B1(n_585),
.B2(n_578),
.Y(n_1992)
);

AND2x2_ASAP7_75t_L g1993 ( 
.A(n_1857),
.B(n_905),
.Y(n_1993)
);

A2O1A1Ixp33_ASAP7_75t_SL g1994 ( 
.A1(n_1870),
.A2(n_907),
.B(n_908),
.C(n_906),
.Y(n_1994)
);

INVx1_ASAP7_75t_L g1995 ( 
.A(n_1866),
.Y(n_1995)
);

INVx2_ASAP7_75t_L g1996 ( 
.A(n_1907),
.Y(n_1996)
);

NOR2xp33_ASAP7_75t_SL g1997 ( 
.A(n_1854),
.B(n_1533),
.Y(n_1997)
);

AOI22xp33_ASAP7_75t_L g1998 ( 
.A1(n_1985),
.A2(n_1236),
.B1(n_1230),
.B2(n_1679),
.Y(n_1998)
);

OAI22xp33_ASAP7_75t_L g1999 ( 
.A1(n_1997),
.A2(n_1007),
.B1(n_1008),
.B2(n_983),
.Y(n_1999)
);

AOI22xp33_ASAP7_75t_L g2000 ( 
.A1(n_1992),
.A2(n_1236),
.B1(n_1658),
.B2(n_1657),
.Y(n_2000)
);

OAI22xp5_ASAP7_75t_SL g2001 ( 
.A1(n_1931),
.A2(n_592),
.B1(n_595),
.B2(n_589),
.Y(n_2001)
);

INVx2_ASAP7_75t_L g2002 ( 
.A(n_1996),
.Y(n_2002)
);

INVx2_ASAP7_75t_L g2003 ( 
.A(n_1922),
.Y(n_2003)
);

AOI22xp33_ASAP7_75t_L g2004 ( 
.A1(n_1992),
.A2(n_1669),
.B1(n_1676),
.B2(n_1664),
.Y(n_2004)
);

INVx1_ASAP7_75t_L g2005 ( 
.A(n_1917),
.Y(n_2005)
);

BUFx6f_ASAP7_75t_L g2006 ( 
.A(n_1928),
.Y(n_2006)
);

INVx5_ASAP7_75t_L g2007 ( 
.A(n_1978),
.Y(n_2007)
);

INVx1_ASAP7_75t_L g2008 ( 
.A(n_1921),
.Y(n_2008)
);

INVx1_ASAP7_75t_L g2009 ( 
.A(n_1995),
.Y(n_2009)
);

INVx1_ASAP7_75t_L g2010 ( 
.A(n_1944),
.Y(n_2010)
);

BUFx2_ASAP7_75t_L g2011 ( 
.A(n_1918),
.Y(n_2011)
);

BUFx10_ASAP7_75t_L g2012 ( 
.A(n_1989),
.Y(n_2012)
);

INVx1_ASAP7_75t_L g2013 ( 
.A(n_1961),
.Y(n_2013)
);

OAI21xp33_ASAP7_75t_L g2014 ( 
.A1(n_1974),
.A2(n_600),
.B(n_599),
.Y(n_2014)
);

CKINVDCx5p33_ASAP7_75t_R g2015 ( 
.A(n_1916),
.Y(n_2015)
);

INVx1_ASAP7_75t_L g2016 ( 
.A(n_1954),
.Y(n_2016)
);

CKINVDCx20_ASAP7_75t_R g2017 ( 
.A(n_1933),
.Y(n_2017)
);

INVx2_ASAP7_75t_SL g2018 ( 
.A(n_1993),
.Y(n_2018)
);

AOI22xp33_ASAP7_75t_L g2019 ( 
.A1(n_1986),
.A2(n_1987),
.B1(n_1919),
.B2(n_1969),
.Y(n_2019)
);

AOI22xp33_ASAP7_75t_L g2020 ( 
.A1(n_1980),
.A2(n_1682),
.B1(n_1683),
.B2(n_1678),
.Y(n_2020)
);

AND2x2_ASAP7_75t_L g2021 ( 
.A(n_1945),
.B(n_1976),
.Y(n_2021)
);

NAND2xp5_ASAP7_75t_L g2022 ( 
.A(n_1951),
.B(n_909),
.Y(n_2022)
);

BUFx2_ASAP7_75t_SL g2023 ( 
.A(n_1989),
.Y(n_2023)
);

INVx4_ASAP7_75t_SL g2024 ( 
.A(n_1991),
.Y(n_2024)
);

INVx8_ASAP7_75t_L g2025 ( 
.A(n_1964),
.Y(n_2025)
);

NAND2xp5_ASAP7_75t_L g2026 ( 
.A(n_1951),
.B(n_1974),
.Y(n_2026)
);

AOI22xp33_ASAP7_75t_L g2027 ( 
.A1(n_1980),
.A2(n_1659),
.B1(n_1661),
.B2(n_1660),
.Y(n_2027)
);

INVx2_ASAP7_75t_L g2028 ( 
.A(n_1929),
.Y(n_2028)
);

BUFx2_ASAP7_75t_L g2029 ( 
.A(n_1923),
.Y(n_2029)
);

INVx1_ASAP7_75t_L g2030 ( 
.A(n_1962),
.Y(n_2030)
);

INVx2_ASAP7_75t_L g2031 ( 
.A(n_1949),
.Y(n_2031)
);

INVx6_ASAP7_75t_L g2032 ( 
.A(n_1953),
.Y(n_2032)
);

INVx1_ASAP7_75t_L g2033 ( 
.A(n_1935),
.Y(n_2033)
);

INVx6_ASAP7_75t_L g2034 ( 
.A(n_1953),
.Y(n_2034)
);

AOI22xp33_ASAP7_75t_SL g2035 ( 
.A1(n_1942),
.A2(n_1735),
.B1(n_1704),
.B2(n_607),
.Y(n_2035)
);

CKINVDCx6p67_ASAP7_75t_R g2036 ( 
.A(n_1970),
.Y(n_2036)
);

INVx3_ASAP7_75t_SL g2037 ( 
.A(n_1990),
.Y(n_2037)
);

CKINVDCx6p67_ASAP7_75t_R g2038 ( 
.A(n_1938),
.Y(n_2038)
);

INVx2_ASAP7_75t_L g2039 ( 
.A(n_1950),
.Y(n_2039)
);

INVx6_ASAP7_75t_L g2040 ( 
.A(n_1948),
.Y(n_2040)
);

BUFx6f_ASAP7_75t_L g2041 ( 
.A(n_1928),
.Y(n_2041)
);

INVx2_ASAP7_75t_L g2042 ( 
.A(n_1958),
.Y(n_2042)
);

INVx2_ASAP7_75t_L g2043 ( 
.A(n_1991),
.Y(n_2043)
);

BUFx2_ASAP7_75t_L g2044 ( 
.A(n_1923),
.Y(n_2044)
);

INVx1_ASAP7_75t_SL g2045 ( 
.A(n_1990),
.Y(n_2045)
);

CKINVDCx6p67_ASAP7_75t_R g2046 ( 
.A(n_1927),
.Y(n_2046)
);

INVx1_ASAP7_75t_L g2047 ( 
.A(n_1935),
.Y(n_2047)
);

INVx3_ASAP7_75t_SL g2048 ( 
.A(n_1927),
.Y(n_2048)
);

INVx8_ASAP7_75t_L g2049 ( 
.A(n_1964),
.Y(n_2049)
);

INVx1_ASAP7_75t_L g2050 ( 
.A(n_1956),
.Y(n_2050)
);

INVx1_ASAP7_75t_L g2051 ( 
.A(n_1956),
.Y(n_2051)
);

INVx1_ASAP7_75t_L g2052 ( 
.A(n_1963),
.Y(n_2052)
);

INVx2_ASAP7_75t_L g2053 ( 
.A(n_1991),
.Y(n_2053)
);

AOI22xp5_ASAP7_75t_L g2054 ( 
.A1(n_1919),
.A2(n_1673),
.B1(n_1735),
.B2(n_1704),
.Y(n_2054)
);

CKINVDCx11_ASAP7_75t_R g2055 ( 
.A(n_1930),
.Y(n_2055)
);

BUFx6f_ASAP7_75t_L g2056 ( 
.A(n_1928),
.Y(n_2056)
);

INVx6_ASAP7_75t_L g2057 ( 
.A(n_1948),
.Y(n_2057)
);

INVx1_ASAP7_75t_L g2058 ( 
.A(n_1940),
.Y(n_2058)
);

NAND2xp5_ASAP7_75t_L g2059 ( 
.A(n_2026),
.B(n_1943),
.Y(n_2059)
);

HB1xp67_ASAP7_75t_L g2060 ( 
.A(n_2026),
.Y(n_2060)
);

INVx1_ASAP7_75t_L g2061 ( 
.A(n_2052),
.Y(n_2061)
);

AOI21xp5_ASAP7_75t_L g2062 ( 
.A1(n_2014),
.A2(n_1973),
.B(n_1959),
.Y(n_2062)
);

INVx2_ASAP7_75t_L g2063 ( 
.A(n_2031),
.Y(n_2063)
);

CKINVDCx6p67_ASAP7_75t_R g2064 ( 
.A(n_2036),
.Y(n_2064)
);

INVx1_ASAP7_75t_L g2065 ( 
.A(n_2005),
.Y(n_2065)
);

AOI21x1_ASAP7_75t_SL g2066 ( 
.A1(n_2022),
.A2(n_1959),
.B(n_1924),
.Y(n_2066)
);

INVx2_ASAP7_75t_SL g2067 ( 
.A(n_2012),
.Y(n_2067)
);

BUFx2_ASAP7_75t_L g2068 ( 
.A(n_2029),
.Y(n_2068)
);

AND2x2_ASAP7_75t_L g2069 ( 
.A(n_2011),
.B(n_2021),
.Y(n_2069)
);

AND2x2_ASAP7_75t_L g2070 ( 
.A(n_2048),
.B(n_1965),
.Y(n_2070)
);

INVx2_ASAP7_75t_L g2071 ( 
.A(n_2039),
.Y(n_2071)
);

BUFx6f_ASAP7_75t_L g2072 ( 
.A(n_2006),
.Y(n_2072)
);

AND2x4_ASAP7_75t_L g2073 ( 
.A(n_2024),
.B(n_1937),
.Y(n_2073)
);

OA21x2_ASAP7_75t_L g2074 ( 
.A1(n_2042),
.A2(n_1924),
.B(n_1981),
.Y(n_2074)
);

HB1xp67_ASAP7_75t_SL g2075 ( 
.A(n_2015),
.Y(n_2075)
);

INVx2_ASAP7_75t_L g2076 ( 
.A(n_2003),
.Y(n_2076)
);

OAI22xp5_ASAP7_75t_L g2077 ( 
.A1(n_2019),
.A2(n_2035),
.B1(n_2046),
.B2(n_2018),
.Y(n_2077)
);

AOI21xp5_ASAP7_75t_L g2078 ( 
.A1(n_2050),
.A2(n_1973),
.B(n_1967),
.Y(n_2078)
);

AOI21xp5_ASAP7_75t_L g2079 ( 
.A1(n_2051),
.A2(n_1967),
.B(n_1960),
.Y(n_2079)
);

NAND2xp5_ASAP7_75t_L g2080 ( 
.A(n_2013),
.B(n_1930),
.Y(n_2080)
);

O2A1O1Ixp5_ASAP7_75t_L g2081 ( 
.A1(n_2010),
.A2(n_2016),
.B(n_2030),
.C(n_2022),
.Y(n_2081)
);

AND2x2_ASAP7_75t_L g2082 ( 
.A(n_2044),
.B(n_1965),
.Y(n_2082)
);

INVx1_ASAP7_75t_L g2083 ( 
.A(n_2008),
.Y(n_2083)
);

INVx2_ASAP7_75t_L g2084 ( 
.A(n_2028),
.Y(n_2084)
);

AND2x4_ASAP7_75t_L g2085 ( 
.A(n_2024),
.B(n_1947),
.Y(n_2085)
);

A2O1A1Ixp33_ASAP7_75t_L g2086 ( 
.A1(n_2035),
.A2(n_1977),
.B(n_1926),
.C(n_1934),
.Y(n_2086)
);

OR2x2_ASAP7_75t_L g2087 ( 
.A(n_2009),
.B(n_1982),
.Y(n_2087)
);

AOI21xp5_ASAP7_75t_L g2088 ( 
.A1(n_2043),
.A2(n_1960),
.B(n_1955),
.Y(n_2088)
);

AOI21x1_ASAP7_75t_SL g2089 ( 
.A1(n_2038),
.A2(n_1984),
.B(n_1920),
.Y(n_2089)
);

INVx2_ASAP7_75t_L g2090 ( 
.A(n_2002),
.Y(n_2090)
);

O2A1O1Ixp33_ASAP7_75t_L g2091 ( 
.A1(n_1999),
.A2(n_1934),
.B(n_1939),
.C(n_1925),
.Y(n_2091)
);

OAI22x1_ASAP7_75t_L g2092 ( 
.A1(n_2045),
.A2(n_1972),
.B1(n_1946),
.B2(n_1971),
.Y(n_2092)
);

NAND2x1p5_ASAP7_75t_L g2093 ( 
.A(n_2007),
.B(n_1948),
.Y(n_2093)
);

OR2x2_ASAP7_75t_L g2094 ( 
.A(n_2033),
.B(n_1968),
.Y(n_2094)
);

INVx1_ASAP7_75t_L g2095 ( 
.A(n_2061),
.Y(n_2095)
);

BUFx3_ASAP7_75t_L g2096 ( 
.A(n_2064),
.Y(n_2096)
);

NAND2xp5_ASAP7_75t_L g2097 ( 
.A(n_2060),
.B(n_2047),
.Y(n_2097)
);

NAND2xp5_ASAP7_75t_L g2098 ( 
.A(n_2059),
.B(n_2058),
.Y(n_2098)
);

NAND2xp5_ASAP7_75t_L g2099 ( 
.A(n_2061),
.B(n_2045),
.Y(n_2099)
);

INVx2_ASAP7_75t_L g2100 ( 
.A(n_2074),
.Y(n_2100)
);

AND2x2_ASAP7_75t_L g2101 ( 
.A(n_2068),
.B(n_2037),
.Y(n_2101)
);

CKINVDCx5p33_ASAP7_75t_R g2102 ( 
.A(n_2075),
.Y(n_2102)
);

INVx2_ASAP7_75t_L g2103 ( 
.A(n_2074),
.Y(n_2103)
);

BUFx2_ASAP7_75t_L g2104 ( 
.A(n_2082),
.Y(n_2104)
);

INVx3_ASAP7_75t_L g2105 ( 
.A(n_2093),
.Y(n_2105)
);

AND2x4_ASAP7_75t_L g2106 ( 
.A(n_2082),
.B(n_2024),
.Y(n_2106)
);

CKINVDCx16_ASAP7_75t_R g2107 ( 
.A(n_2077),
.Y(n_2107)
);

AND2x2_ASAP7_75t_L g2108 ( 
.A(n_2068),
.B(n_2023),
.Y(n_2108)
);

INVx2_ASAP7_75t_SL g2109 ( 
.A(n_2087),
.Y(n_2109)
);

BUFx3_ASAP7_75t_L g2110 ( 
.A(n_2064),
.Y(n_2110)
);

OR2x2_ASAP7_75t_L g2111 ( 
.A(n_2087),
.B(n_1957),
.Y(n_2111)
);

NOR2xp33_ASAP7_75t_R g2112 ( 
.A(n_2067),
.B(n_2017),
.Y(n_2112)
);

CKINVDCx14_ASAP7_75t_R g2113 ( 
.A(n_2069),
.Y(n_2113)
);

INVx1_ASAP7_75t_L g2114 ( 
.A(n_2065),
.Y(n_2114)
);

INVx2_ASAP7_75t_L g2115 ( 
.A(n_2074),
.Y(n_2115)
);

CKINVDCx5p33_ASAP7_75t_R g2116 ( 
.A(n_2067),
.Y(n_2116)
);

INVx2_ASAP7_75t_L g2117 ( 
.A(n_2074),
.Y(n_2117)
);

NAND3xp33_ASAP7_75t_SL g2118 ( 
.A(n_2062),
.B(n_2054),
.C(n_1998),
.Y(n_2118)
);

AND2x4_ASAP7_75t_L g2119 ( 
.A(n_2073),
.B(n_2007),
.Y(n_2119)
);

OAI222xp33_ASAP7_75t_L g2120 ( 
.A1(n_2107),
.A2(n_1999),
.B1(n_2094),
.B2(n_2078),
.C1(n_2079),
.C2(n_2084),
.Y(n_2120)
);

INVx2_ASAP7_75t_L g2121 ( 
.A(n_2100),
.Y(n_2121)
);

OR2x6_ASAP7_75t_L g2122 ( 
.A(n_2119),
.B(n_2092),
.Y(n_2122)
);

AO21x2_ASAP7_75t_L g2123 ( 
.A1(n_2100),
.A2(n_2086),
.B(n_2091),
.Y(n_2123)
);

INVx1_ASAP7_75t_L g2124 ( 
.A(n_2095),
.Y(n_2124)
);

OR2x2_ASAP7_75t_L g2125 ( 
.A(n_2097),
.B(n_2065),
.Y(n_2125)
);

OA21x2_ASAP7_75t_L g2126 ( 
.A1(n_2100),
.A2(n_2081),
.B(n_2088),
.Y(n_2126)
);

AND2x2_ASAP7_75t_L g2127 ( 
.A(n_2113),
.B(n_2070),
.Y(n_2127)
);

AND2x2_ASAP7_75t_L g2128 ( 
.A(n_2113),
.B(n_2070),
.Y(n_2128)
);

INVx1_ASAP7_75t_L g2129 ( 
.A(n_2095),
.Y(n_2129)
);

OR2x6_ASAP7_75t_L g2130 ( 
.A(n_2119),
.B(n_2092),
.Y(n_2130)
);

INVx1_ASAP7_75t_L g2131 ( 
.A(n_2114),
.Y(n_2131)
);

NAND2x1_ASAP7_75t_L g2132 ( 
.A(n_2106),
.B(n_2069),
.Y(n_2132)
);

INVx2_ASAP7_75t_L g2133 ( 
.A(n_2103),
.Y(n_2133)
);

OAI22xp5_ASAP7_75t_L g2134 ( 
.A1(n_2107),
.A2(n_2080),
.B1(n_2034),
.B2(n_2032),
.Y(n_2134)
);

INVx1_ASAP7_75t_L g2135 ( 
.A(n_2114),
.Y(n_2135)
);

NAND2xp5_ASAP7_75t_L g2136 ( 
.A(n_2098),
.B(n_2083),
.Y(n_2136)
);

INVx1_ASAP7_75t_L g2137 ( 
.A(n_2097),
.Y(n_2137)
);

HB1xp67_ASAP7_75t_L g2138 ( 
.A(n_2099),
.Y(n_2138)
);

INVx1_ASAP7_75t_L g2139 ( 
.A(n_2109),
.Y(n_2139)
);

NAND3xp33_ASAP7_75t_L g2140 ( 
.A(n_2109),
.B(n_2111),
.C(n_2004),
.Y(n_2140)
);

INVx2_ASAP7_75t_L g2141 ( 
.A(n_2103),
.Y(n_2141)
);

AND2x2_ASAP7_75t_L g2142 ( 
.A(n_2104),
.B(n_2101),
.Y(n_2142)
);

INVx1_ASAP7_75t_L g2143 ( 
.A(n_2109),
.Y(n_2143)
);

OA21x2_ASAP7_75t_L g2144 ( 
.A1(n_2103),
.A2(n_2071),
.B(n_2063),
.Y(n_2144)
);

OR2x2_ASAP7_75t_L g2145 ( 
.A(n_2098),
.B(n_2083),
.Y(n_2145)
);

BUFx6f_ASAP7_75t_L g2146 ( 
.A(n_2096),
.Y(n_2146)
);

INVx2_ASAP7_75t_L g2147 ( 
.A(n_2115),
.Y(n_2147)
);

INVx3_ASAP7_75t_L g2148 ( 
.A(n_2119),
.Y(n_2148)
);

INVx1_ASAP7_75t_L g2149 ( 
.A(n_2099),
.Y(n_2149)
);

AND2x2_ASAP7_75t_L g2150 ( 
.A(n_2104),
.B(n_2072),
.Y(n_2150)
);

AND2x2_ASAP7_75t_L g2151 ( 
.A(n_2104),
.B(n_2072),
.Y(n_2151)
);

BUFx2_ASAP7_75t_L g2152 ( 
.A(n_2142),
.Y(n_2152)
);

AND2x2_ASAP7_75t_L g2153 ( 
.A(n_2142),
.B(n_2096),
.Y(n_2153)
);

AND2x2_ASAP7_75t_L g2154 ( 
.A(n_2127),
.B(n_2096),
.Y(n_2154)
);

AND2x2_ASAP7_75t_L g2155 ( 
.A(n_2127),
.B(n_2096),
.Y(n_2155)
);

INVx2_ASAP7_75t_L g2156 ( 
.A(n_2126),
.Y(n_2156)
);

AND2x2_ASAP7_75t_L g2157 ( 
.A(n_2150),
.B(n_2105),
.Y(n_2157)
);

NOR2x1p5_ASAP7_75t_L g2158 ( 
.A(n_2146),
.B(n_2110),
.Y(n_2158)
);

HB1xp67_ASAP7_75t_L g2159 ( 
.A(n_2124),
.Y(n_2159)
);

AND2x2_ASAP7_75t_L g2160 ( 
.A(n_2128),
.B(n_2110),
.Y(n_2160)
);

AND2x2_ASAP7_75t_L g2161 ( 
.A(n_2150),
.B(n_2151),
.Y(n_2161)
);

OR2x2_ASAP7_75t_L g2162 ( 
.A(n_2125),
.B(n_2111),
.Y(n_2162)
);

INVx1_ASAP7_75t_L g2163 ( 
.A(n_2124),
.Y(n_2163)
);

AND2x2_ASAP7_75t_L g2164 ( 
.A(n_2151),
.B(n_2105),
.Y(n_2164)
);

AND2x2_ASAP7_75t_L g2165 ( 
.A(n_2148),
.B(n_2105),
.Y(n_2165)
);

AOI22xp33_ASAP7_75t_L g2166 ( 
.A1(n_2123),
.A2(n_2118),
.B1(n_2115),
.B2(n_2117),
.Y(n_2166)
);

AND2x2_ASAP7_75t_L g2167 ( 
.A(n_2128),
.B(n_2110),
.Y(n_2167)
);

INVx1_ASAP7_75t_L g2168 ( 
.A(n_2129),
.Y(n_2168)
);

INVx1_ASAP7_75t_L g2169 ( 
.A(n_2129),
.Y(n_2169)
);

INVx2_ASAP7_75t_L g2170 ( 
.A(n_2126),
.Y(n_2170)
);

OAI221xp5_ASAP7_75t_SL g2171 ( 
.A1(n_2122),
.A2(n_2111),
.B1(n_1998),
.B2(n_2110),
.C(n_2000),
.Y(n_2171)
);

AND2x2_ASAP7_75t_L g2172 ( 
.A(n_2148),
.B(n_2105),
.Y(n_2172)
);

BUFx12f_ASAP7_75t_L g2173 ( 
.A(n_2146),
.Y(n_2173)
);

NAND3xp33_ASAP7_75t_L g2174 ( 
.A(n_2166),
.B(n_2146),
.C(n_2140),
.Y(n_2174)
);

AOI22xp33_ASAP7_75t_L g2175 ( 
.A1(n_2156),
.A2(n_2123),
.B1(n_2130),
.B2(n_2122),
.Y(n_2175)
);

INVx2_ASAP7_75t_L g2176 ( 
.A(n_2156),
.Y(n_2176)
);

NAND2xp5_ASAP7_75t_L g2177 ( 
.A(n_2152),
.B(n_2123),
.Y(n_2177)
);

OAI221xp5_ASAP7_75t_L g2178 ( 
.A1(n_2171),
.A2(n_2122),
.B1(n_2130),
.B2(n_2140),
.C(n_2126),
.Y(n_2178)
);

AOI33xp33_ASAP7_75t_L g2179 ( 
.A1(n_2153),
.A2(n_2137),
.A3(n_2149),
.B1(n_2143),
.B2(n_2139),
.B3(n_2131),
.Y(n_2179)
);

INVxp67_ASAP7_75t_SL g2180 ( 
.A(n_2158),
.Y(n_2180)
);

NAND4xp25_ASAP7_75t_SL g2181 ( 
.A(n_2153),
.B(n_2101),
.C(n_2108),
.D(n_2139),
.Y(n_2181)
);

AND2x2_ASAP7_75t_L g2182 ( 
.A(n_2154),
.B(n_2146),
.Y(n_2182)
);

INVx1_ASAP7_75t_L g2183 ( 
.A(n_2159),
.Y(n_2183)
);

INVx2_ASAP7_75t_L g2184 ( 
.A(n_2156),
.Y(n_2184)
);

NAND2xp5_ASAP7_75t_L g2185 ( 
.A(n_2152),
.B(n_2137),
.Y(n_2185)
);

AND2x2_ASAP7_75t_L g2186 ( 
.A(n_2154),
.B(n_2146),
.Y(n_2186)
);

AND2x2_ASAP7_75t_L g2187 ( 
.A(n_2155),
.B(n_2146),
.Y(n_2187)
);

AND2x4_ASAP7_75t_L g2188 ( 
.A(n_2158),
.B(n_2148),
.Y(n_2188)
);

OAI31xp33_ASAP7_75t_L g2189 ( 
.A1(n_2171),
.A2(n_2120),
.A3(n_2134),
.B(n_2001),
.Y(n_2189)
);

BUFx3_ASAP7_75t_L g2190 ( 
.A(n_2173),
.Y(n_2190)
);

BUFx2_ASAP7_75t_L g2191 ( 
.A(n_2182),
.Y(n_2191)
);

HB1xp67_ASAP7_75t_L g2192 ( 
.A(n_2182),
.Y(n_2192)
);

AND2x2_ASAP7_75t_L g2193 ( 
.A(n_2186),
.B(n_2155),
.Y(n_2193)
);

BUFx2_ASAP7_75t_L g2194 ( 
.A(n_2186),
.Y(n_2194)
);

BUFx3_ASAP7_75t_L g2195 ( 
.A(n_2190),
.Y(n_2195)
);

INVx1_ASAP7_75t_L g2196 ( 
.A(n_2176),
.Y(n_2196)
);

AND2x2_ASAP7_75t_L g2197 ( 
.A(n_2187),
.B(n_2160),
.Y(n_2197)
);

INVx2_ASAP7_75t_L g2198 ( 
.A(n_2176),
.Y(n_2198)
);

AND2x2_ASAP7_75t_L g2199 ( 
.A(n_2187),
.B(n_2160),
.Y(n_2199)
);

OR2x2_ASAP7_75t_L g2200 ( 
.A(n_2191),
.B(n_2177),
.Y(n_2200)
);

HB1xp67_ASAP7_75t_L g2201 ( 
.A(n_2191),
.Y(n_2201)
);

OR2x2_ASAP7_75t_L g2202 ( 
.A(n_2194),
.B(n_2185),
.Y(n_2202)
);

OR2x2_ASAP7_75t_L g2203 ( 
.A(n_2194),
.B(n_2174),
.Y(n_2203)
);

HB1xp67_ASAP7_75t_L g2204 ( 
.A(n_2193),
.Y(n_2204)
);

INVx1_ASAP7_75t_L g2205 ( 
.A(n_2198),
.Y(n_2205)
);

NAND2xp5_ASAP7_75t_L g2206 ( 
.A(n_2192),
.B(n_2179),
.Y(n_2206)
);

AND2x2_ASAP7_75t_L g2207 ( 
.A(n_2204),
.B(n_2193),
.Y(n_2207)
);

NOR2x1p5_ASAP7_75t_L g2208 ( 
.A(n_2202),
.B(n_2195),
.Y(n_2208)
);

NAND2xp5_ASAP7_75t_L g2209 ( 
.A(n_2201),
.B(n_2197),
.Y(n_2209)
);

INVx1_ASAP7_75t_L g2210 ( 
.A(n_2205),
.Y(n_2210)
);

NAND2xp5_ASAP7_75t_L g2211 ( 
.A(n_2200),
.B(n_2197),
.Y(n_2211)
);

NAND2xp5_ASAP7_75t_L g2212 ( 
.A(n_2207),
.B(n_2199),
.Y(n_2212)
);

AOI322xp5_ASAP7_75t_L g2213 ( 
.A1(n_2210),
.A2(n_2175),
.A3(n_2206),
.B1(n_2198),
.B2(n_2196),
.C1(n_2170),
.C2(n_2184),
.Y(n_2213)
);

AND2x2_ASAP7_75t_L g2214 ( 
.A(n_2208),
.B(n_2167),
.Y(n_2214)
);

INVx1_ASAP7_75t_L g2215 ( 
.A(n_2212),
.Y(n_2215)
);

INVx1_ASAP7_75t_L g2216 ( 
.A(n_2214),
.Y(n_2216)
);

AOI22xp5_ASAP7_75t_SL g2217 ( 
.A1(n_2215),
.A2(n_2195),
.B1(n_2209),
.B2(n_2211),
.Y(n_2217)
);

OR2x2_ASAP7_75t_L g2218 ( 
.A(n_2216),
.B(n_2203),
.Y(n_2218)
);

AOI21xp33_ASAP7_75t_SL g2219 ( 
.A1(n_2218),
.A2(n_2174),
.B(n_2189),
.Y(n_2219)
);

HB1xp67_ASAP7_75t_L g2220 ( 
.A(n_2217),
.Y(n_2220)
);

INVx1_ASAP7_75t_L g2221 ( 
.A(n_2220),
.Y(n_2221)
);

AND2x2_ASAP7_75t_L g2222 ( 
.A(n_2219),
.B(n_2199),
.Y(n_2222)
);

INVx1_ASAP7_75t_L g2223 ( 
.A(n_2220),
.Y(n_2223)
);

INVx1_ASAP7_75t_L g2224 ( 
.A(n_2222),
.Y(n_2224)
);

NOR3xp33_ASAP7_75t_L g2225 ( 
.A(n_2221),
.B(n_2178),
.C(n_2184),
.Y(n_2225)
);

INVxp67_ASAP7_75t_L g2226 ( 
.A(n_2222),
.Y(n_2226)
);

NOR2xp33_ASAP7_75t_L g2227 ( 
.A(n_2223),
.B(n_2190),
.Y(n_2227)
);

INVx2_ASAP7_75t_SL g2228 ( 
.A(n_2224),
.Y(n_2228)
);

AOI21xp5_ASAP7_75t_L g2229 ( 
.A1(n_2226),
.A2(n_2180),
.B(n_2183),
.Y(n_2229)
);

INVx1_ASAP7_75t_L g2230 ( 
.A(n_2227),
.Y(n_2230)
);

NAND3xp33_ASAP7_75t_L g2231 ( 
.A(n_2228),
.B(n_2225),
.C(n_2213),
.Y(n_2231)
);

INVx1_ASAP7_75t_L g2232 ( 
.A(n_2230),
.Y(n_2232)
);

AOI211xp5_ASAP7_75t_L g2233 ( 
.A1(n_2229),
.A2(n_2183),
.B(n_2190),
.C(n_2170),
.Y(n_2233)
);

NAND2xp5_ASAP7_75t_L g2234 ( 
.A(n_2228),
.B(n_2189),
.Y(n_2234)
);

OR2x2_ASAP7_75t_L g2235 ( 
.A(n_2228),
.B(n_2170),
.Y(n_2235)
);

OAI221xp5_ASAP7_75t_SL g2236 ( 
.A1(n_2229),
.A2(n_2167),
.B1(n_2162),
.B2(n_2130),
.C(n_2122),
.Y(n_2236)
);

NAND2xp5_ASAP7_75t_SL g2237 ( 
.A(n_2228),
.B(n_2188),
.Y(n_2237)
);

NAND4xp75_ASAP7_75t_L g2238 ( 
.A(n_2228),
.B(n_912),
.C(n_915),
.D(n_910),
.Y(n_2238)
);

NAND4xp25_ASAP7_75t_L g2239 ( 
.A(n_2229),
.B(n_2188),
.C(n_1994),
.D(n_1988),
.Y(n_2239)
);

AND2x2_ASAP7_75t_L g2240 ( 
.A(n_2228),
.B(n_2188),
.Y(n_2240)
);

OAI211xp5_ASAP7_75t_L g2241 ( 
.A1(n_2228),
.A2(n_2159),
.B(n_917),
.C(n_918),
.Y(n_2241)
);

AND3x1_ASAP7_75t_L g2242 ( 
.A(n_2228),
.B(n_2161),
.C(n_2165),
.Y(n_2242)
);

AND4x1_ASAP7_75t_L g2243 ( 
.A(n_2230),
.B(n_920),
.C(n_921),
.D(n_916),
.Y(n_2243)
);

AOI211xp5_ASAP7_75t_L g2244 ( 
.A1(n_2229),
.A2(n_2188),
.B(n_2181),
.C(n_926),
.Y(n_2244)
);

NAND4xp25_ASAP7_75t_L g2245 ( 
.A(n_2231),
.B(n_1952),
.C(n_1936),
.D(n_927),
.Y(n_2245)
);

NOR3xp33_ASAP7_75t_L g2246 ( 
.A(n_2232),
.B(n_929),
.C(n_923),
.Y(n_2246)
);

NAND3xp33_ASAP7_75t_L g2247 ( 
.A(n_2243),
.B(n_932),
.C(n_930),
.Y(n_2247)
);

AOI221xp5_ASAP7_75t_L g2248 ( 
.A1(n_2234),
.A2(n_2169),
.B1(n_2168),
.B2(n_2163),
.C(n_2141),
.Y(n_2248)
);

AOI21xp5_ASAP7_75t_L g2249 ( 
.A1(n_2237),
.A2(n_2163),
.B(n_2168),
.Y(n_2249)
);

OAI211xp5_ASAP7_75t_SL g2250 ( 
.A1(n_2233),
.A2(n_934),
.B(n_936),
.C(n_933),
.Y(n_2250)
);

NOR2xp33_ASAP7_75t_L g2251 ( 
.A(n_2235),
.B(n_2102),
.Y(n_2251)
);

AOI211xp5_ASAP7_75t_L g2252 ( 
.A1(n_2240),
.A2(n_939),
.B(n_944),
.C(n_938),
.Y(n_2252)
);

OAI211xp5_ASAP7_75t_SL g2253 ( 
.A1(n_2244),
.A2(n_948),
.B(n_949),
.C(n_946),
.Y(n_2253)
);

AOI221xp5_ASAP7_75t_L g2254 ( 
.A1(n_2242),
.A2(n_2169),
.B1(n_2141),
.B2(n_2147),
.C(n_2133),
.Y(n_2254)
);

NAND3xp33_ASAP7_75t_SL g2255 ( 
.A(n_2241),
.B(n_706),
.C(n_650),
.Y(n_2255)
);

NOR4xp25_ASAP7_75t_L g2256 ( 
.A(n_2236),
.B(n_955),
.C(n_956),
.D(n_951),
.Y(n_2256)
);

AOI211xp5_ASAP7_75t_L g2257 ( 
.A1(n_2239),
.A2(n_963),
.B(n_966),
.C(n_962),
.Y(n_2257)
);

AND4x1_ASAP7_75t_L g2258 ( 
.A(n_2238),
.B(n_969),
.C(n_2161),
.D(n_1352),
.Y(n_2258)
);

NOR2x1_ASAP7_75t_L g2259 ( 
.A(n_2231),
.B(n_2161),
.Y(n_2259)
);

AOI211xp5_ASAP7_75t_L g2260 ( 
.A1(n_2231),
.A2(n_614),
.B(n_619),
.C(n_605),
.Y(n_2260)
);

NAND4xp25_ASAP7_75t_L g2261 ( 
.A(n_2231),
.B(n_2172),
.C(n_2165),
.D(n_1932),
.Y(n_2261)
);

AOI211xp5_ASAP7_75t_L g2262 ( 
.A1(n_2231),
.A2(n_627),
.B(n_631),
.C(n_620),
.Y(n_2262)
);

AND2x2_ASAP7_75t_L g2263 ( 
.A(n_2240),
.B(n_2165),
.Y(n_2263)
);

AOI211xp5_ASAP7_75t_L g2264 ( 
.A1(n_2231),
.A2(n_644),
.B(n_645),
.C(n_639),
.Y(n_2264)
);

OAI211xp5_ASAP7_75t_SL g2265 ( 
.A1(n_2237),
.A2(n_2162),
.B(n_2148),
.C(n_2173),
.Y(n_2265)
);

NOR3xp33_ASAP7_75t_L g2266 ( 
.A(n_2232),
.B(n_1237),
.C(n_652),
.Y(n_2266)
);

NOR2x1_ASAP7_75t_L g2267 ( 
.A(n_2231),
.B(n_2172),
.Y(n_2267)
);

NOR2x1_ASAP7_75t_L g2268 ( 
.A(n_2231),
.B(n_2172),
.Y(n_2268)
);

AND2x2_ASAP7_75t_L g2269 ( 
.A(n_2240),
.B(n_2157),
.Y(n_2269)
);

NAND4xp25_ASAP7_75t_L g2270 ( 
.A(n_2231),
.B(n_2157),
.C(n_2164),
.D(n_1186),
.Y(n_2270)
);

AOI221xp5_ASAP7_75t_SL g2271 ( 
.A1(n_2237),
.A2(n_2157),
.B1(n_2164),
.B2(n_2143),
.C(n_2173),
.Y(n_2271)
);

OAI211xp5_ASAP7_75t_SL g2272 ( 
.A1(n_2237),
.A2(n_1353),
.B(n_1357),
.C(n_1350),
.Y(n_2272)
);

AOI211xp5_ASAP7_75t_L g2273 ( 
.A1(n_2231),
.A2(n_671),
.B(n_674),
.C(n_649),
.Y(n_2273)
);

NAND3xp33_ASAP7_75t_L g2274 ( 
.A(n_2231),
.B(n_688),
.C(n_677),
.Y(n_2274)
);

AOI221xp5_ASAP7_75t_L g2275 ( 
.A1(n_2231),
.A2(n_2141),
.B1(n_2147),
.B2(n_2133),
.C(n_2121),
.Y(n_2275)
);

NAND3xp33_ASAP7_75t_L g2276 ( 
.A(n_2231),
.B(n_699),
.C(n_690),
.Y(n_2276)
);

NAND4xp25_ASAP7_75t_L g2277 ( 
.A(n_2231),
.B(n_2164),
.C(n_1152),
.D(n_1144),
.Y(n_2277)
);

AND4x1_ASAP7_75t_L g2278 ( 
.A(n_2231),
.B(n_1362),
.C(n_1335),
.D(n_1337),
.Y(n_2278)
);

NAND2xp5_ASAP7_75t_SL g2279 ( 
.A(n_2231),
.B(n_2112),
.Y(n_2279)
);

NOR2xp33_ASAP7_75t_L g2280 ( 
.A(n_2231),
.B(n_2133),
.Y(n_2280)
);

INVx1_ASAP7_75t_L g2281 ( 
.A(n_2242),
.Y(n_2281)
);

NAND3xp33_ASAP7_75t_L g2282 ( 
.A(n_2231),
.B(n_707),
.C(n_705),
.Y(n_2282)
);

NAND2x1_ASAP7_75t_L g2283 ( 
.A(n_2240),
.B(n_2149),
.Y(n_2283)
);

AOI221xp5_ASAP7_75t_L g2284 ( 
.A1(n_2231),
.A2(n_2147),
.B1(n_2121),
.B2(n_716),
.C(n_717),
.Y(n_2284)
);

NAND5xp2_ASAP7_75t_L g2285 ( 
.A(n_2234),
.B(n_2000),
.C(n_1966),
.D(n_1119),
.E(n_1135),
.Y(n_2285)
);

NOR2x1_ASAP7_75t_L g2286 ( 
.A(n_2231),
.B(n_2132),
.Y(n_2286)
);

AOI211xp5_ASAP7_75t_SL g2287 ( 
.A1(n_2241),
.A2(n_1344),
.B(n_1333),
.C(n_2138),
.Y(n_2287)
);

AOI21xp5_ASAP7_75t_L g2288 ( 
.A1(n_2237),
.A2(n_714),
.B(n_713),
.Y(n_2288)
);

OAI321xp33_ASAP7_75t_L g2289 ( 
.A1(n_2231),
.A2(n_2122),
.A3(n_2130),
.B1(n_2121),
.B2(n_1975),
.C(n_2118),
.Y(n_2289)
);

NAND4xp75_ASAP7_75t_L g2290 ( 
.A(n_2232),
.B(n_2126),
.C(n_1108),
.D(n_1139),
.Y(n_2290)
);

NOR2xp33_ASAP7_75t_SL g2291 ( 
.A(n_2240),
.B(n_726),
.Y(n_2291)
);

INVx2_ASAP7_75t_SL g2292 ( 
.A(n_2263),
.Y(n_2292)
);

INVx2_ASAP7_75t_L g2293 ( 
.A(n_2269),
.Y(n_2293)
);

NOR2x1_ASAP7_75t_L g2294 ( 
.A(n_2274),
.B(n_2132),
.Y(n_2294)
);

CKINVDCx6p67_ASAP7_75t_R g2295 ( 
.A(n_2279),
.Y(n_2295)
);

AOI221x1_ASAP7_75t_L g2296 ( 
.A1(n_2253),
.A2(n_2135),
.B1(n_2131),
.B2(n_2101),
.C(n_1283),
.Y(n_2296)
);

NOR3x2_ASAP7_75t_L g2297 ( 
.A(n_2257),
.B(n_729),
.C(n_727),
.Y(n_2297)
);

INVxp67_ASAP7_75t_L g2298 ( 
.A(n_2259),
.Y(n_2298)
);

AOI21xp5_ASAP7_75t_L g2299 ( 
.A1(n_2267),
.A2(n_732),
.B(n_731),
.Y(n_2299)
);

AOI22xp33_ASAP7_75t_R g2300 ( 
.A1(n_2281),
.A2(n_743),
.B1(n_746),
.B2(n_739),
.Y(n_2300)
);

NAND2xp33_ASAP7_75t_R g2301 ( 
.A(n_2288),
.B(n_754),
.Y(n_2301)
);

INVxp67_ASAP7_75t_L g2302 ( 
.A(n_2291),
.Y(n_2302)
);

AOI22xp5_ASAP7_75t_L g2303 ( 
.A1(n_2251),
.A2(n_2130),
.B1(n_2135),
.B2(n_2116),
.Y(n_2303)
);

OAI211xp5_ASAP7_75t_L g2304 ( 
.A1(n_2260),
.A2(n_764),
.B(n_765),
.C(n_763),
.Y(n_2304)
);

NAND2xp5_ASAP7_75t_L g2305 ( 
.A(n_2268),
.B(n_767),
.Y(n_2305)
);

NAND2xp33_ASAP7_75t_SL g2306 ( 
.A(n_2283),
.B(n_2112),
.Y(n_2306)
);

INVx1_ASAP7_75t_L g2307 ( 
.A(n_2286),
.Y(n_2307)
);

AOI222xp33_ASAP7_75t_L g2308 ( 
.A1(n_2280),
.A2(n_771),
.B1(n_768),
.B2(n_781),
.C1(n_774),
.C2(n_770),
.Y(n_2308)
);

OAI22xp5_ASAP7_75t_L g2309 ( 
.A1(n_2262),
.A2(n_2125),
.B1(n_2145),
.B2(n_2136),
.Y(n_2309)
);

NAND4xp25_ASAP7_75t_SL g2310 ( 
.A(n_2271),
.B(n_2108),
.C(n_2145),
.D(n_1975),
.Y(n_2310)
);

NOR2xp33_ASAP7_75t_R g2311 ( 
.A(n_2255),
.B(n_7),
.Y(n_2311)
);

INVx1_ASAP7_75t_L g2312 ( 
.A(n_2258),
.Y(n_2312)
);

NAND2xp5_ASAP7_75t_L g2313 ( 
.A(n_2264),
.B(n_784),
.Y(n_2313)
);

NOR3xp33_ASAP7_75t_L g2314 ( 
.A(n_2276),
.B(n_793),
.C(n_785),
.Y(n_2314)
);

NAND2xp5_ASAP7_75t_L g2315 ( 
.A(n_2273),
.B(n_2278),
.Y(n_2315)
);

INVx2_ASAP7_75t_L g2316 ( 
.A(n_2290),
.Y(n_2316)
);

NAND2xp5_ASAP7_75t_L g2317 ( 
.A(n_2256),
.B(n_2144),
.Y(n_2317)
);

O2A1O1Ixp33_ASAP7_75t_L g2318 ( 
.A1(n_2250),
.A2(n_1094),
.B(n_1209),
.C(n_1249),
.Y(n_2318)
);

NAND3xp33_ASAP7_75t_L g2319 ( 
.A(n_2282),
.B(n_1232),
.C(n_1227),
.Y(n_2319)
);

INVx1_ASAP7_75t_L g2320 ( 
.A(n_2247),
.Y(n_2320)
);

AOI21xp33_ASAP7_75t_L g2321 ( 
.A1(n_2284),
.A2(n_1251),
.B(n_1250),
.Y(n_2321)
);

INVx1_ASAP7_75t_L g2322 ( 
.A(n_2270),
.Y(n_2322)
);

BUFx2_ASAP7_75t_L g2323 ( 
.A(n_2277),
.Y(n_2323)
);

NAND4xp25_ASAP7_75t_SL g2324 ( 
.A(n_2248),
.B(n_2108),
.C(n_1979),
.D(n_12),
.Y(n_2324)
);

NAND4xp75_ASAP7_75t_L g2325 ( 
.A(n_2275),
.B(n_1284),
.C(n_1285),
.D(n_1270),
.Y(n_2325)
);

NAND2xp5_ASAP7_75t_L g2326 ( 
.A(n_2266),
.B(n_2144),
.Y(n_2326)
);

AND2x2_ASAP7_75t_L g2327 ( 
.A(n_2287),
.B(n_2106),
.Y(n_2327)
);

NAND2x1_ASAP7_75t_SL g2328 ( 
.A(n_2272),
.B(n_2105),
.Y(n_2328)
);

A2O1A1Ixp33_ASAP7_75t_SL g2329 ( 
.A1(n_2246),
.A2(n_1261),
.B(n_1256),
.C(n_12),
.Y(n_2329)
);

AOI322xp5_ASAP7_75t_L g2330 ( 
.A1(n_2254),
.A2(n_2117),
.A3(n_2115),
.B1(n_1972),
.B2(n_2004),
.C1(n_2106),
.C2(n_2027),
.Y(n_2330)
);

NAND3xp33_ASAP7_75t_L g2331 ( 
.A(n_2252),
.B(n_481),
.C(n_480),
.Y(n_2331)
);

NAND2xp33_ASAP7_75t_SL g2332 ( 
.A(n_2265),
.B(n_2072),
.Y(n_2332)
);

BUFx3_ASAP7_75t_L g2333 ( 
.A(n_2245),
.Y(n_2333)
);

OAI221xp5_ASAP7_75t_L g2334 ( 
.A1(n_2249),
.A2(n_2117),
.B1(n_1421),
.B2(n_2144),
.C(n_2072),
.Y(n_2334)
);

NAND2xp5_ASAP7_75t_L g2335 ( 
.A(n_2261),
.B(n_2144),
.Y(n_2335)
);

AND2x4_ASAP7_75t_L g2336 ( 
.A(n_2285),
.B(n_2119),
.Y(n_2336)
);

NAND4xp25_ASAP7_75t_SL g2337 ( 
.A(n_2289),
.B(n_13),
.C(n_9),
.D(n_10),
.Y(n_2337)
);

INVx1_ASAP7_75t_L g2338 ( 
.A(n_2259),
.Y(n_2338)
);

AOI21xp5_ASAP7_75t_SL g2339 ( 
.A1(n_2288),
.A2(n_491),
.B(n_487),
.Y(n_2339)
);

AOI22xp5_ASAP7_75t_L g2340 ( 
.A1(n_2251),
.A2(n_2106),
.B1(n_2055),
.B2(n_2119),
.Y(n_2340)
);

INVx1_ASAP7_75t_L g2341 ( 
.A(n_2259),
.Y(n_2341)
);

NAND2xp5_ASAP7_75t_L g2342 ( 
.A(n_2269),
.B(n_10),
.Y(n_2342)
);

NAND2xp5_ASAP7_75t_L g2343 ( 
.A(n_2269),
.B(n_14),
.Y(n_2343)
);

NAND3xp33_ASAP7_75t_L g2344 ( 
.A(n_2260),
.B(n_494),
.C(n_492),
.Y(n_2344)
);

NOR4xp25_ASAP7_75t_L g2345 ( 
.A(n_2281),
.B(n_16),
.C(n_14),
.D(n_15),
.Y(n_2345)
);

INVx1_ASAP7_75t_L g2346 ( 
.A(n_2259),
.Y(n_2346)
);

BUFx2_ASAP7_75t_L g2347 ( 
.A(n_2259),
.Y(n_2347)
);

BUFx6f_ASAP7_75t_L g2348 ( 
.A(n_2247),
.Y(n_2348)
);

INVx2_ASAP7_75t_L g2349 ( 
.A(n_2269),
.Y(n_2349)
);

INVx2_ASAP7_75t_L g2350 ( 
.A(n_2269),
.Y(n_2350)
);

INVx1_ASAP7_75t_SL g2351 ( 
.A(n_2259),
.Y(n_2351)
);

OAI22x1_ASAP7_75t_L g2352 ( 
.A1(n_2258),
.A2(n_2106),
.B1(n_2093),
.B2(n_18),
.Y(n_2352)
);

NOR3xp33_ASAP7_75t_L g2353 ( 
.A(n_2281),
.B(n_496),
.C(n_495),
.Y(n_2353)
);

INVx2_ASAP7_75t_L g2354 ( 
.A(n_2269),
.Y(n_2354)
);

AOI211xp5_ASAP7_75t_SL g2355 ( 
.A1(n_2281),
.A2(n_19),
.B(n_15),
.C(n_17),
.Y(n_2355)
);

NAND2xp5_ASAP7_75t_L g2356 ( 
.A(n_2269),
.B(n_19),
.Y(n_2356)
);

CKINVDCx20_ASAP7_75t_R g2357 ( 
.A(n_2279),
.Y(n_2357)
);

NAND2xp5_ASAP7_75t_L g2358 ( 
.A(n_2269),
.B(n_20),
.Y(n_2358)
);

HB1xp67_ASAP7_75t_L g2359 ( 
.A(n_2259),
.Y(n_2359)
);

AND2x2_ASAP7_75t_L g2360 ( 
.A(n_2259),
.B(n_2012),
.Y(n_2360)
);

INVx1_ASAP7_75t_L g2361 ( 
.A(n_2259),
.Y(n_2361)
);

BUFx2_ASAP7_75t_L g2362 ( 
.A(n_2259),
.Y(n_2362)
);

INVx1_ASAP7_75t_L g2363 ( 
.A(n_2259),
.Y(n_2363)
);

OAI21xp33_ASAP7_75t_SL g2364 ( 
.A1(n_2279),
.A2(n_20),
.B(n_22),
.Y(n_2364)
);

NOR2xp33_ASAP7_75t_R g2365 ( 
.A(n_2281),
.B(n_25),
.Y(n_2365)
);

AOI22xp5_ASAP7_75t_L g2366 ( 
.A1(n_2251),
.A2(n_2072),
.B1(n_2034),
.B2(n_2032),
.Y(n_2366)
);

NAND2xp5_ASAP7_75t_L g2367 ( 
.A(n_2269),
.B(n_25),
.Y(n_2367)
);

AOI22xp33_ASAP7_75t_L g2368 ( 
.A1(n_2259),
.A2(n_2094),
.B1(n_2027),
.B2(n_2020),
.Y(n_2368)
);

INVx1_ASAP7_75t_L g2369 ( 
.A(n_2259),
.Y(n_2369)
);

OAI211xp5_ASAP7_75t_SL g2370 ( 
.A1(n_2260),
.A2(n_30),
.B(n_26),
.C(n_28),
.Y(n_2370)
);

OAI21xp33_ASAP7_75t_L g2371 ( 
.A1(n_2259),
.A2(n_2020),
.B(n_509),
.Y(n_2371)
);

INVx1_ASAP7_75t_L g2372 ( 
.A(n_2259),
.Y(n_2372)
);

AND2x2_ASAP7_75t_SL g2373 ( 
.A(n_2256),
.B(n_26),
.Y(n_2373)
);

XNOR2x2_ASAP7_75t_SL g2374 ( 
.A(n_2274),
.B(n_31),
.Y(n_2374)
);

CKINVDCx5p33_ASAP7_75t_R g2375 ( 
.A(n_2281),
.Y(n_2375)
);

XOR2xp5_ASAP7_75t_L g2376 ( 
.A(n_2259),
.B(n_31),
.Y(n_2376)
);

AOI21xp5_ASAP7_75t_L g2377 ( 
.A1(n_2259),
.A2(n_512),
.B(n_503),
.Y(n_2377)
);

NOR2xp33_ASAP7_75t_L g2378 ( 
.A(n_2251),
.B(n_33),
.Y(n_2378)
);

AOI322xp5_ASAP7_75t_L g2379 ( 
.A1(n_2259),
.A2(n_2049),
.A3(n_2025),
.B1(n_2076),
.B2(n_2084),
.C1(n_2085),
.C2(n_2073),
.Y(n_2379)
);

NAND2xp33_ASAP7_75t_R g2380 ( 
.A(n_2281),
.B(n_35),
.Y(n_2380)
);

AOI221xp5_ASAP7_75t_L g2381 ( 
.A1(n_2251),
.A2(n_523),
.B1(n_524),
.B2(n_521),
.C(n_518),
.Y(n_2381)
);

A2O1A1Ixp33_ASAP7_75t_SL g2382 ( 
.A1(n_2257),
.A2(n_39),
.B(n_37),
.C(n_38),
.Y(n_2382)
);

INVx1_ASAP7_75t_L g2383 ( 
.A(n_2259),
.Y(n_2383)
);

NAND3xp33_ASAP7_75t_L g2384 ( 
.A(n_2260),
.B(n_532),
.C(n_529),
.Y(n_2384)
);

INVxp67_ASAP7_75t_L g2385 ( 
.A(n_2259),
.Y(n_2385)
);

HB1xp67_ASAP7_75t_L g2386 ( 
.A(n_2259),
.Y(n_2386)
);

INVx1_ASAP7_75t_L g2387 ( 
.A(n_2259),
.Y(n_2387)
);

NAND2xp5_ASAP7_75t_L g2388 ( 
.A(n_2269),
.B(n_37),
.Y(n_2388)
);

AOI22xp5_ASAP7_75t_L g2389 ( 
.A1(n_2251),
.A2(n_2034),
.B1(n_2032),
.B2(n_2025),
.Y(n_2389)
);

OAI322xp33_ASAP7_75t_L g2390 ( 
.A1(n_2298),
.A2(n_46),
.A3(n_44),
.B1(n_41),
.B2(n_39),
.C1(n_40),
.C2(n_43),
.Y(n_2390)
);

NOR2x1_ASAP7_75t_L g2391 ( 
.A(n_2347),
.B(n_40),
.Y(n_2391)
);

NOR2xp67_ASAP7_75t_L g2392 ( 
.A(n_2385),
.B(n_43),
.Y(n_2392)
);

NAND4xp75_ASAP7_75t_L g2393 ( 
.A(n_2338),
.B(n_53),
.C(n_47),
.D(n_49),
.Y(n_2393)
);

INVx2_ASAP7_75t_L g2394 ( 
.A(n_2373),
.Y(n_2394)
);

NAND2x1p5_ASAP7_75t_L g2395 ( 
.A(n_2351),
.B(n_2362),
.Y(n_2395)
);

AND2x4_ASAP7_75t_L g2396 ( 
.A(n_2292),
.B(n_47),
.Y(n_2396)
);

INVx1_ASAP7_75t_L g2397 ( 
.A(n_2359),
.Y(n_2397)
);

NOR3xp33_ASAP7_75t_L g2398 ( 
.A(n_2341),
.B(n_549),
.C(n_544),
.Y(n_2398)
);

NOR2x1p5_ASAP7_75t_L g2399 ( 
.A(n_2346),
.B(n_53),
.Y(n_2399)
);

NAND4xp75_ASAP7_75t_L g2400 ( 
.A(n_2361),
.B(n_57),
.C(n_54),
.D(n_56),
.Y(n_2400)
);

INVx1_ASAP7_75t_L g2401 ( 
.A(n_2386),
.Y(n_2401)
);

NAND4xp75_ASAP7_75t_L g2402 ( 
.A(n_2363),
.B(n_2372),
.C(n_2383),
.D(n_2369),
.Y(n_2402)
);

INVx1_ASAP7_75t_L g2403 ( 
.A(n_2376),
.Y(n_2403)
);

AO22x2_ASAP7_75t_L g2404 ( 
.A1(n_2387),
.A2(n_59),
.B1(n_54),
.B2(n_58),
.Y(n_2404)
);

AOI22xp5_ASAP7_75t_L g2405 ( 
.A1(n_2375),
.A2(n_2049),
.B1(n_2025),
.B2(n_1183),
.Y(n_2405)
);

NOR2x1_ASAP7_75t_L g2406 ( 
.A(n_2307),
.B(n_59),
.Y(n_2406)
);

AND2x4_ASAP7_75t_L g2407 ( 
.A(n_2360),
.B(n_61),
.Y(n_2407)
);

NAND2xp5_ASAP7_75t_L g2408 ( 
.A(n_2336),
.B(n_61),
.Y(n_2408)
);

INVx1_ASAP7_75t_L g2409 ( 
.A(n_2317),
.Y(n_2409)
);

XOR2xp5_ASAP7_75t_L g2410 ( 
.A(n_2357),
.B(n_66),
.Y(n_2410)
);

INVx1_ASAP7_75t_L g2411 ( 
.A(n_2305),
.Y(n_2411)
);

INVx2_ASAP7_75t_L g2412 ( 
.A(n_2336),
.Y(n_2412)
);

OAI22xp5_ASAP7_75t_SL g2413 ( 
.A1(n_2342),
.A2(n_68),
.B1(n_66),
.B2(n_67),
.Y(n_2413)
);

INVx2_ASAP7_75t_SL g2414 ( 
.A(n_2293),
.Y(n_2414)
);

AOI22xp5_ASAP7_75t_L g2415 ( 
.A1(n_2306),
.A2(n_2049),
.B1(n_1183),
.B2(n_1156),
.Y(n_2415)
);

INVx2_ASAP7_75t_L g2416 ( 
.A(n_2352),
.Y(n_2416)
);

NAND4xp75_ASAP7_75t_L g2417 ( 
.A(n_2349),
.B(n_72),
.C(n_67),
.D(n_71),
.Y(n_2417)
);

NOR3xp33_ASAP7_75t_L g2418 ( 
.A(n_2350),
.B(n_552),
.C(n_551),
.Y(n_2418)
);

INVx2_ASAP7_75t_L g2419 ( 
.A(n_2327),
.Y(n_2419)
);

NOR2xp67_ASAP7_75t_L g2420 ( 
.A(n_2364),
.B(n_72),
.Y(n_2420)
);

AO22x1_ASAP7_75t_L g2421 ( 
.A1(n_2354),
.A2(n_75),
.B1(n_73),
.B2(n_74),
.Y(n_2421)
);

XOR2xp5_ASAP7_75t_L g2422 ( 
.A(n_2374),
.B(n_73),
.Y(n_2422)
);

NOR2x1_ASAP7_75t_L g2423 ( 
.A(n_2331),
.B(n_75),
.Y(n_2423)
);

NAND4xp75_ASAP7_75t_L g2424 ( 
.A(n_2378),
.B(n_78),
.C(n_76),
.D(n_77),
.Y(n_2424)
);

AOI22xp33_ASAP7_75t_SL g2425 ( 
.A1(n_2365),
.A2(n_1275),
.B1(n_1156),
.B2(n_1183),
.Y(n_2425)
);

INVx1_ASAP7_75t_L g2426 ( 
.A(n_2343),
.Y(n_2426)
);

AO22x1_ASAP7_75t_L g2427 ( 
.A1(n_2314),
.A2(n_2312),
.B1(n_2358),
.B2(n_2356),
.Y(n_2427)
);

XOR2xp5_ASAP7_75t_L g2428 ( 
.A(n_2322),
.B(n_76),
.Y(n_2428)
);

AOI22xp5_ASAP7_75t_L g2429 ( 
.A1(n_2380),
.A2(n_2332),
.B1(n_2388),
.B2(n_2367),
.Y(n_2429)
);

INVx1_ASAP7_75t_L g2430 ( 
.A(n_2326),
.Y(n_2430)
);

NOR2x1_ASAP7_75t_L g2431 ( 
.A(n_2344),
.B(n_77),
.Y(n_2431)
);

INVx1_ASAP7_75t_L g2432 ( 
.A(n_2295),
.Y(n_2432)
);

INVx2_ASAP7_75t_L g2433 ( 
.A(n_2297),
.Y(n_2433)
);

NOR4xp75_ASAP7_75t_L g2434 ( 
.A(n_2315),
.B(n_82),
.C(n_78),
.D(n_79),
.Y(n_2434)
);

AOI22xp33_ASAP7_75t_SL g2435 ( 
.A1(n_2311),
.A2(n_1275),
.B1(n_773),
.B2(n_628),
.Y(n_2435)
);

NAND4xp75_ASAP7_75t_L g2436 ( 
.A(n_2299),
.B(n_84),
.C(n_79),
.D(n_83),
.Y(n_2436)
);

OR2x2_ASAP7_75t_L g2437 ( 
.A(n_2345),
.B(n_84),
.Y(n_2437)
);

NAND2xp5_ASAP7_75t_L g2438 ( 
.A(n_2302),
.B(n_85),
.Y(n_2438)
);

INVx1_ASAP7_75t_L g2439 ( 
.A(n_2313),
.Y(n_2439)
);

OR2x2_ASAP7_75t_L g2440 ( 
.A(n_2337),
.B(n_2335),
.Y(n_2440)
);

INVx2_ASAP7_75t_L g2441 ( 
.A(n_2328),
.Y(n_2441)
);

NOR2x1_ASAP7_75t_L g2442 ( 
.A(n_2384),
.B(n_86),
.Y(n_2442)
);

NAND2x1p5_ASAP7_75t_L g2443 ( 
.A(n_2333),
.B(n_1948),
.Y(n_2443)
);

INVx1_ASAP7_75t_L g2444 ( 
.A(n_2323),
.Y(n_2444)
);

NAND3xp33_ASAP7_75t_L g2445 ( 
.A(n_2300),
.B(n_773),
.C(n_628),
.Y(n_2445)
);

NAND4xp75_ASAP7_75t_L g2446 ( 
.A(n_2377),
.B(n_88),
.C(n_86),
.D(n_87),
.Y(n_2446)
);

XNOR2x1_ASAP7_75t_L g2447 ( 
.A(n_2316),
.B(n_87),
.Y(n_2447)
);

INVx1_ASAP7_75t_SL g2448 ( 
.A(n_2348),
.Y(n_2448)
);

NAND2xp5_ASAP7_75t_L g2449 ( 
.A(n_2308),
.B(n_89),
.Y(n_2449)
);

NOR3xp33_ASAP7_75t_L g2450 ( 
.A(n_2321),
.B(n_577),
.C(n_563),
.Y(n_2450)
);

OR2x2_ASAP7_75t_L g2451 ( 
.A(n_2324),
.B(n_89),
.Y(n_2451)
);

INVx1_ASAP7_75t_L g2452 ( 
.A(n_2348),
.Y(n_2452)
);

BUFx4f_ASAP7_75t_L g2453 ( 
.A(n_2348),
.Y(n_2453)
);

INVx1_ASAP7_75t_L g2454 ( 
.A(n_2318),
.Y(n_2454)
);

NAND3xp33_ASAP7_75t_L g2455 ( 
.A(n_2353),
.B(n_2355),
.C(n_2301),
.Y(n_2455)
);

OR2x2_ASAP7_75t_L g2456 ( 
.A(n_2310),
.B(n_90),
.Y(n_2456)
);

INVx1_ASAP7_75t_L g2457 ( 
.A(n_2370),
.Y(n_2457)
);

INVx1_ASAP7_75t_L g2458 ( 
.A(n_2319),
.Y(n_2458)
);

INVx1_ASAP7_75t_L g2459 ( 
.A(n_2304),
.Y(n_2459)
);

INVx1_ASAP7_75t_L g2460 ( 
.A(n_2294),
.Y(n_2460)
);

OR2x2_ASAP7_75t_L g2461 ( 
.A(n_2303),
.B(n_90),
.Y(n_2461)
);

CKINVDCx6p67_ASAP7_75t_R g2462 ( 
.A(n_2320),
.Y(n_2462)
);

NOR2x1_ASAP7_75t_L g2463 ( 
.A(n_2339),
.B(n_91),
.Y(n_2463)
);

NAND4xp75_ASAP7_75t_L g2464 ( 
.A(n_2381),
.B(n_94),
.C(n_92),
.D(n_93),
.Y(n_2464)
);

NOR2xp67_ASAP7_75t_L g2465 ( 
.A(n_2371),
.B(n_92),
.Y(n_2465)
);

INVx1_ASAP7_75t_L g2466 ( 
.A(n_2325),
.Y(n_2466)
);

NOR2xp67_ASAP7_75t_L g2467 ( 
.A(n_2340),
.B(n_95),
.Y(n_2467)
);

XOR2x1_ASAP7_75t_L g2468 ( 
.A(n_2329),
.B(n_97),
.Y(n_2468)
);

NOR2x1_ASAP7_75t_L g2469 ( 
.A(n_2334),
.B(n_98),
.Y(n_2469)
);

NOR2x1_ASAP7_75t_L g2470 ( 
.A(n_2309),
.B(n_101),
.Y(n_2470)
);

NOR3xp33_ASAP7_75t_L g2471 ( 
.A(n_2397),
.B(n_2382),
.C(n_2366),
.Y(n_2471)
);

NAND5xp2_ASAP7_75t_L g2472 ( 
.A(n_2395),
.B(n_2401),
.C(n_2432),
.D(n_2429),
.E(n_2452),
.Y(n_2472)
);

NOR2x1_ASAP7_75t_L g2473 ( 
.A(n_2402),
.B(n_2296),
.Y(n_2473)
);

NOR2x1_ASAP7_75t_L g2474 ( 
.A(n_2412),
.B(n_2460),
.Y(n_2474)
);

AND2x2_ASAP7_75t_L g2475 ( 
.A(n_2394),
.B(n_2379),
.Y(n_2475)
);

AOI211xp5_ASAP7_75t_L g2476 ( 
.A1(n_2441),
.A2(n_2389),
.B(n_2330),
.C(n_2368),
.Y(n_2476)
);

AND2x4_ASAP7_75t_L g2477 ( 
.A(n_2414),
.B(n_103),
.Y(n_2477)
);

NOR3xp33_ASAP7_75t_SL g2478 ( 
.A(n_2444),
.B(n_583),
.C(n_580),
.Y(n_2478)
);

NAND2xp5_ASAP7_75t_L g2479 ( 
.A(n_2448),
.B(n_2462),
.Y(n_2479)
);

NOR3xp33_ASAP7_75t_L g2480 ( 
.A(n_2430),
.B(n_587),
.C(n_586),
.Y(n_2480)
);

NOR3xp33_ASAP7_75t_SL g2481 ( 
.A(n_2409),
.B(n_594),
.C(n_590),
.Y(n_2481)
);

INVx2_ASAP7_75t_L g2482 ( 
.A(n_2468),
.Y(n_2482)
);

AND3x1_ASAP7_75t_L g2483 ( 
.A(n_2391),
.B(n_103),
.C(n_104),
.Y(n_2483)
);

NAND3xp33_ASAP7_75t_SL g2484 ( 
.A(n_2419),
.B(n_598),
.C(n_597),
.Y(n_2484)
);

BUFx2_ASAP7_75t_L g2485 ( 
.A(n_2406),
.Y(n_2485)
);

INVx2_ASAP7_75t_L g2486 ( 
.A(n_2399),
.Y(n_2486)
);

NOR5xp2_ASAP7_75t_L g2487 ( 
.A(n_2455),
.B(n_2445),
.C(n_2459),
.D(n_2403),
.E(n_2411),
.Y(n_2487)
);

NOR2xp67_ASAP7_75t_L g2488 ( 
.A(n_2437),
.B(n_105),
.Y(n_2488)
);

AO211x2_ASAP7_75t_L g2489 ( 
.A1(n_2408),
.A2(n_108),
.B(n_106),
.C(n_107),
.Y(n_2489)
);

INVx2_ASAP7_75t_L g2490 ( 
.A(n_2404),
.Y(n_2490)
);

OR3x2_ASAP7_75t_L g2491 ( 
.A(n_2440),
.B(n_106),
.C(n_107),
.Y(n_2491)
);

AOI21xp5_ASAP7_75t_L g2492 ( 
.A1(n_2453),
.A2(n_604),
.B(n_603),
.Y(n_2492)
);

NAND5xp2_ASAP7_75t_L g2493 ( 
.A(n_2457),
.B(n_110),
.C(n_108),
.D(n_109),
.E(n_111),
.Y(n_2493)
);

NAND4xp75_ASAP7_75t_L g2494 ( 
.A(n_2392),
.B(n_2470),
.C(n_2463),
.D(n_2420),
.Y(n_2494)
);

NOR4xp25_ASAP7_75t_L g2495 ( 
.A(n_2416),
.B(n_114),
.C(n_112),
.D(n_113),
.Y(n_2495)
);

HB1xp67_ASAP7_75t_L g2496 ( 
.A(n_2434),
.Y(n_2496)
);

AND2x4_ASAP7_75t_L g2497 ( 
.A(n_2407),
.B(n_112),
.Y(n_2497)
);

NAND4xp25_ASAP7_75t_L g2498 ( 
.A(n_2467),
.B(n_116),
.C(n_114),
.D(n_115),
.Y(n_2498)
);

NOR4xp25_ASAP7_75t_L g2499 ( 
.A(n_2426),
.B(n_118),
.C(n_116),
.D(n_117),
.Y(n_2499)
);

NAND2xp5_ASAP7_75t_L g2500 ( 
.A(n_2427),
.B(n_117),
.Y(n_2500)
);

NAND2xp5_ASAP7_75t_SL g2501 ( 
.A(n_2396),
.B(n_610),
.Y(n_2501)
);

NAND2x1p5_ASAP7_75t_L g2502 ( 
.A(n_2396),
.B(n_1507),
.Y(n_2502)
);

NAND4xp25_ASAP7_75t_SL g2503 ( 
.A(n_2451),
.B(n_120),
.C(n_118),
.D(n_119),
.Y(n_2503)
);

NAND4xp75_ASAP7_75t_L g2504 ( 
.A(n_2431),
.B(n_122),
.C(n_120),
.D(n_121),
.Y(n_2504)
);

NAND4xp75_ASAP7_75t_L g2505 ( 
.A(n_2442),
.B(n_124),
.C(n_122),
.D(n_123),
.Y(n_2505)
);

INVx2_ASAP7_75t_L g2506 ( 
.A(n_2404),
.Y(n_2506)
);

NAND2xp5_ASAP7_75t_L g2507 ( 
.A(n_2433),
.B(n_123),
.Y(n_2507)
);

INVx2_ASAP7_75t_SL g2508 ( 
.A(n_2447),
.Y(n_2508)
);

NOR2x1_ASAP7_75t_L g2509 ( 
.A(n_2422),
.B(n_2393),
.Y(n_2509)
);

NOR3xp33_ASAP7_75t_L g2510 ( 
.A(n_2439),
.B(n_621),
.C(n_613),
.Y(n_2510)
);

NOR2x1_ASAP7_75t_L g2511 ( 
.A(n_2400),
.B(n_628),
.Y(n_2511)
);

OAI211xp5_ASAP7_75t_L g2512 ( 
.A1(n_2449),
.A2(n_128),
.B(n_124),
.C(n_127),
.Y(n_2512)
);

NOR2x1p5_ASAP7_75t_L g2513 ( 
.A(n_2424),
.B(n_128),
.Y(n_2513)
);

NAND2xp5_ASAP7_75t_L g2514 ( 
.A(n_2454),
.B(n_130),
.Y(n_2514)
);

NAND4xp75_ASAP7_75t_L g2515 ( 
.A(n_2423),
.B(n_137),
.C(n_132),
.D(n_136),
.Y(n_2515)
);

NAND2xp5_ASAP7_75t_L g2516 ( 
.A(n_2410),
.B(n_132),
.Y(n_2516)
);

NOR3xp33_ASAP7_75t_L g2517 ( 
.A(n_2398),
.B(n_640),
.C(n_629),
.Y(n_2517)
);

NAND4xp25_ASAP7_75t_L g2518 ( 
.A(n_2435),
.B(n_139),
.C(n_137),
.D(n_138),
.Y(n_2518)
);

OR5x1_ASAP7_75t_L g2519 ( 
.A(n_2456),
.B(n_140),
.C(n_138),
.D(n_139),
.E(n_141),
.Y(n_2519)
);

NAND3xp33_ASAP7_75t_L g2520 ( 
.A(n_2418),
.B(n_773),
.C(n_628),
.Y(n_2520)
);

NOR3xp33_ASAP7_75t_L g2521 ( 
.A(n_2450),
.B(n_2458),
.C(n_2421),
.Y(n_2521)
);

NOR2xp33_ASAP7_75t_L g2522 ( 
.A(n_2428),
.B(n_140),
.Y(n_2522)
);

AO22x1_ASAP7_75t_L g2523 ( 
.A1(n_2438),
.A2(n_2466),
.B1(n_2469),
.B2(n_2464),
.Y(n_2523)
);

INVx1_ASAP7_75t_L g2524 ( 
.A(n_2413),
.Y(n_2524)
);

OAI211xp5_ASAP7_75t_SL g2525 ( 
.A1(n_2461),
.A2(n_143),
.B(n_141),
.C(n_142),
.Y(n_2525)
);

NOR2x1_ASAP7_75t_L g2526 ( 
.A(n_2417),
.B(n_773),
.Y(n_2526)
);

HB1xp67_ASAP7_75t_L g2527 ( 
.A(n_2436),
.Y(n_2527)
);

AND2x4_ASAP7_75t_L g2528 ( 
.A(n_2465),
.B(n_142),
.Y(n_2528)
);

NOR2x1_ASAP7_75t_L g2529 ( 
.A(n_2446),
.B(n_2390),
.Y(n_2529)
);

NAND5xp2_ASAP7_75t_L g2530 ( 
.A(n_2443),
.B(n_145),
.C(n_143),
.D(n_144),
.E(n_147),
.Y(n_2530)
);

AND2x4_ASAP7_75t_L g2531 ( 
.A(n_2405),
.B(n_144),
.Y(n_2531)
);

AND2x4_ASAP7_75t_L g2532 ( 
.A(n_2415),
.B(n_148),
.Y(n_2532)
);

NAND3xp33_ASAP7_75t_L g2533 ( 
.A(n_2425),
.B(n_773),
.C(n_651),
.Y(n_2533)
);

NAND3xp33_ASAP7_75t_L g2534 ( 
.A(n_2397),
.B(n_653),
.C(n_648),
.Y(n_2534)
);

OAI211xp5_ASAP7_75t_SL g2535 ( 
.A1(n_2397),
.A2(n_151),
.B(n_149),
.C(n_150),
.Y(n_2535)
);

NOR2xp33_ASAP7_75t_L g2536 ( 
.A(n_2395),
.B(n_149),
.Y(n_2536)
);

NOR4xp25_ASAP7_75t_L g2537 ( 
.A(n_2397),
.B(n_157),
.C(n_150),
.D(n_154),
.Y(n_2537)
);

NOR4xp25_ASAP7_75t_L g2538 ( 
.A(n_2397),
.B(n_159),
.C(n_157),
.D(n_158),
.Y(n_2538)
);

NOR3xp33_ASAP7_75t_L g2539 ( 
.A(n_2397),
.B(n_657),
.C(n_656),
.Y(n_2539)
);

BUFx2_ASAP7_75t_L g2540 ( 
.A(n_2483),
.Y(n_2540)
);

BUFx2_ASAP7_75t_L g2541 ( 
.A(n_2485),
.Y(n_2541)
);

BUFx2_ASAP7_75t_L g2542 ( 
.A(n_2474),
.Y(n_2542)
);

INVx1_ASAP7_75t_L g2543 ( 
.A(n_2479),
.Y(n_2543)
);

CKINVDCx20_ASAP7_75t_R g2544 ( 
.A(n_2496),
.Y(n_2544)
);

CKINVDCx5p33_ASAP7_75t_R g2545 ( 
.A(n_2482),
.Y(n_2545)
);

CKINVDCx5p33_ASAP7_75t_R g2546 ( 
.A(n_2508),
.Y(n_2546)
);

INVx1_ASAP7_75t_L g2547 ( 
.A(n_2494),
.Y(n_2547)
);

INVx1_ASAP7_75t_L g2548 ( 
.A(n_2488),
.Y(n_2548)
);

INVx1_ASAP7_75t_SL g2549 ( 
.A(n_2519),
.Y(n_2549)
);

INVx2_ASAP7_75t_L g2550 ( 
.A(n_2491),
.Y(n_2550)
);

INVx1_ASAP7_75t_SL g2551 ( 
.A(n_2528),
.Y(n_2551)
);

CKINVDCx5p33_ASAP7_75t_R g2552 ( 
.A(n_2486),
.Y(n_2552)
);

INVx1_ASAP7_75t_SL g2553 ( 
.A(n_2528),
.Y(n_2553)
);

NAND2xp5_ASAP7_75t_L g2554 ( 
.A(n_2490),
.B(n_159),
.Y(n_2554)
);

INVx2_ASAP7_75t_L g2555 ( 
.A(n_2506),
.Y(n_2555)
);

INVx1_ASAP7_75t_L g2556 ( 
.A(n_2477),
.Y(n_2556)
);

CKINVDCx20_ASAP7_75t_R g2557 ( 
.A(n_2500),
.Y(n_2557)
);

INVx1_ASAP7_75t_L g2558 ( 
.A(n_2477),
.Y(n_2558)
);

CKINVDCx20_ASAP7_75t_R g2559 ( 
.A(n_2527),
.Y(n_2559)
);

INVx1_ASAP7_75t_SL g2560 ( 
.A(n_2497),
.Y(n_2560)
);

AOI21xp33_ASAP7_75t_SL g2561 ( 
.A1(n_2536),
.A2(n_162),
.B(n_163),
.Y(n_2561)
);

CKINVDCx5p33_ASAP7_75t_R g2562 ( 
.A(n_2523),
.Y(n_2562)
);

AND2x4_ASAP7_75t_L g2563 ( 
.A(n_2497),
.B(n_165),
.Y(n_2563)
);

HB1xp67_ASAP7_75t_L g2564 ( 
.A(n_2473),
.Y(n_2564)
);

CKINVDCx5p33_ASAP7_75t_R g2565 ( 
.A(n_2475),
.Y(n_2565)
);

NOR2xp33_ASAP7_75t_R g2566 ( 
.A(n_2484),
.B(n_2503),
.Y(n_2566)
);

INVx2_ASAP7_75t_SL g2567 ( 
.A(n_2513),
.Y(n_2567)
);

XOR2xp5_ASAP7_75t_L g2568 ( 
.A(n_2509),
.B(n_166),
.Y(n_2568)
);

CKINVDCx5p33_ASAP7_75t_R g2569 ( 
.A(n_2524),
.Y(n_2569)
);

INVxp33_ASAP7_75t_L g2570 ( 
.A(n_2522),
.Y(n_2570)
);

CKINVDCx16_ASAP7_75t_R g2571 ( 
.A(n_2529),
.Y(n_2571)
);

CKINVDCx5p33_ASAP7_75t_R g2572 ( 
.A(n_2481),
.Y(n_2572)
);

NAND2xp5_ASAP7_75t_L g2573 ( 
.A(n_2471),
.B(n_167),
.Y(n_2573)
);

XNOR2xp5_ASAP7_75t_L g2574 ( 
.A(n_2489),
.B(n_168),
.Y(n_2574)
);

CKINVDCx5p33_ASAP7_75t_R g2575 ( 
.A(n_2478),
.Y(n_2575)
);

NAND2xp5_ASAP7_75t_L g2576 ( 
.A(n_2516),
.B(n_169),
.Y(n_2576)
);

CKINVDCx5p33_ASAP7_75t_R g2577 ( 
.A(n_2472),
.Y(n_2577)
);

AOI221xp5_ASAP7_75t_L g2578 ( 
.A1(n_2495),
.A2(n_2538),
.B1(n_2537),
.B2(n_2499),
.C(n_2525),
.Y(n_2578)
);

BUFx2_ASAP7_75t_L g2579 ( 
.A(n_2514),
.Y(n_2579)
);

CKINVDCx5p33_ASAP7_75t_R g2580 ( 
.A(n_2501),
.Y(n_2580)
);

INVx1_ASAP7_75t_SL g2581 ( 
.A(n_2507),
.Y(n_2581)
);

INVx1_ASAP7_75t_L g2582 ( 
.A(n_2502),
.Y(n_2582)
);

INVx1_ASAP7_75t_SL g2583 ( 
.A(n_2504),
.Y(n_2583)
);

INVx1_ASAP7_75t_SL g2584 ( 
.A(n_2505),
.Y(n_2584)
);

INVx1_ASAP7_75t_SL g2585 ( 
.A(n_2515),
.Y(n_2585)
);

NAND2xp5_ASAP7_75t_L g2586 ( 
.A(n_2521),
.B(n_2492),
.Y(n_2586)
);

CKINVDCx20_ASAP7_75t_R g2587 ( 
.A(n_2487),
.Y(n_2587)
);

AOI221xp5_ASAP7_75t_L g2588 ( 
.A1(n_2498),
.A2(n_669),
.B1(n_673),
.B2(n_667),
.C(n_660),
.Y(n_2588)
);

INVx3_ASAP7_75t_SL g2589 ( 
.A(n_2532),
.Y(n_2589)
);

BUFx2_ASAP7_75t_L g2590 ( 
.A(n_2526),
.Y(n_2590)
);

HB1xp67_ASAP7_75t_L g2591 ( 
.A(n_2511),
.Y(n_2591)
);

OAI21xp5_ASAP7_75t_L g2592 ( 
.A1(n_2512),
.A2(n_1294),
.B(n_1275),
.Y(n_2592)
);

INVx6_ASAP7_75t_L g2593 ( 
.A(n_2532),
.Y(n_2593)
);

INVx1_ASAP7_75t_SL g2594 ( 
.A(n_2531),
.Y(n_2594)
);

INVx1_ASAP7_75t_L g2595 ( 
.A(n_2493),
.Y(n_2595)
);

INVxp67_ASAP7_75t_SL g2596 ( 
.A(n_2539),
.Y(n_2596)
);

OAI211xp5_ASAP7_75t_SL g2597 ( 
.A1(n_2476),
.A2(n_172),
.B(n_170),
.C(n_171),
.Y(n_2597)
);

INVx2_ASAP7_75t_SL g2598 ( 
.A(n_2531),
.Y(n_2598)
);

NAND2xp5_ASAP7_75t_L g2599 ( 
.A(n_2480),
.B(n_171),
.Y(n_2599)
);

CKINVDCx6p67_ASAP7_75t_R g2600 ( 
.A(n_2530),
.Y(n_2600)
);

OAI211xp5_ASAP7_75t_L g2601 ( 
.A1(n_2517),
.A2(n_178),
.B(n_175),
.C(n_177),
.Y(n_2601)
);

INVx1_ASAP7_75t_L g2602 ( 
.A(n_2535),
.Y(n_2602)
);

NOR2x1p5_ASAP7_75t_L g2603 ( 
.A(n_2518),
.B(n_177),
.Y(n_2603)
);

NAND3x1_ASAP7_75t_L g2604 ( 
.A(n_2510),
.B(n_182),
.C(n_183),
.Y(n_2604)
);

CKINVDCx5p33_ASAP7_75t_R g2605 ( 
.A(n_2534),
.Y(n_2605)
);

OAI222xp33_ASAP7_75t_L g2606 ( 
.A1(n_2533),
.A2(n_2093),
.B1(n_183),
.B2(n_184),
.C1(n_186),
.C2(n_187),
.Y(n_2606)
);

NOR2x1p5_ASAP7_75t_L g2607 ( 
.A(n_2520),
.B(n_182),
.Y(n_2607)
);

NOR2xp33_ASAP7_75t_R g2608 ( 
.A(n_2479),
.B(n_184),
.Y(n_2608)
);

BUFx3_ASAP7_75t_L g2609 ( 
.A(n_2485),
.Y(n_2609)
);

OR2x2_ASAP7_75t_L g2610 ( 
.A(n_2472),
.B(n_186),
.Y(n_2610)
);

NAND2xp5_ASAP7_75t_L g2611 ( 
.A(n_2474),
.B(n_188),
.Y(n_2611)
);

XOR2xp5_ASAP7_75t_L g2612 ( 
.A(n_2479),
.B(n_188),
.Y(n_2612)
);

OR2x2_ASAP7_75t_L g2613 ( 
.A(n_2472),
.B(n_189),
.Y(n_2613)
);

CKINVDCx5p33_ASAP7_75t_R g2614 ( 
.A(n_2479),
.Y(n_2614)
);

INVx1_ASAP7_75t_SL g2615 ( 
.A(n_2485),
.Y(n_2615)
);

HB1xp67_ASAP7_75t_SL g2616 ( 
.A(n_2482),
.Y(n_2616)
);

INVx1_ASAP7_75t_L g2617 ( 
.A(n_2485),
.Y(n_2617)
);

O2A1O1Ixp33_ASAP7_75t_L g2618 ( 
.A1(n_2542),
.A2(n_1422),
.B(n_1415),
.C(n_1507),
.Y(n_2618)
);

AOI22xp33_ASAP7_75t_L g2619 ( 
.A1(n_2541),
.A2(n_678),
.B1(n_681),
.B2(n_675),
.Y(n_2619)
);

OAI211xp5_ASAP7_75t_L g2620 ( 
.A1(n_2577),
.A2(n_191),
.B(n_189),
.C(n_190),
.Y(n_2620)
);

XNOR2xp5_ASAP7_75t_L g2621 ( 
.A(n_2544),
.B(n_191),
.Y(n_2621)
);

AOI322xp5_ASAP7_75t_L g2622 ( 
.A1(n_2587),
.A2(n_193),
.A3(n_194),
.B1(n_195),
.B2(n_196),
.C1(n_197),
.C2(n_198),
.Y(n_2622)
);

OAI211xp5_ASAP7_75t_L g2623 ( 
.A1(n_2615),
.A2(n_199),
.B(n_194),
.C(n_198),
.Y(n_2623)
);

AOI221xp5_ASAP7_75t_L g2624 ( 
.A1(n_2609),
.A2(n_787),
.B1(n_791),
.B2(n_789),
.C(n_782),
.Y(n_2624)
);

AND2x2_ASAP7_75t_L g2625 ( 
.A(n_2571),
.B(n_2073),
.Y(n_2625)
);

INVx2_ASAP7_75t_L g2626 ( 
.A(n_2540),
.Y(n_2626)
);

INVx2_ASAP7_75t_L g2627 ( 
.A(n_2559),
.Y(n_2627)
);

OAI221xp5_ASAP7_75t_L g2628 ( 
.A1(n_2617),
.A2(n_200),
.B1(n_201),
.B2(n_202),
.C(n_203),
.Y(n_2628)
);

NAND5xp2_ASAP7_75t_L g2629 ( 
.A(n_2595),
.B(n_200),
.C(n_201),
.D(n_202),
.E(n_204),
.Y(n_2629)
);

AOI322xp5_ASAP7_75t_L g2630 ( 
.A1(n_2564),
.A2(n_206),
.A3(n_207),
.B1(n_208),
.B2(n_209),
.C1(n_210),
.C2(n_211),
.Y(n_2630)
);

AOI322xp5_ASAP7_75t_L g2631 ( 
.A1(n_2549),
.A2(n_206),
.A3(n_212),
.B1(n_213),
.B2(n_214),
.C1(n_215),
.C2(n_216),
.Y(n_2631)
);

OAI322xp33_ASAP7_75t_L g2632 ( 
.A1(n_2547),
.A2(n_212),
.A3(n_213),
.B1(n_215),
.B2(n_216),
.C1(n_217),
.C2(n_219),
.Y(n_2632)
);

NAND3xp33_ASAP7_75t_SL g2633 ( 
.A(n_2565),
.B(n_689),
.C(n_686),
.Y(n_2633)
);

NOR2x1_ASAP7_75t_L g2634 ( 
.A(n_2610),
.B(n_1301),
.Y(n_2634)
);

OR2x2_ASAP7_75t_L g2635 ( 
.A(n_2551),
.B(n_221),
.Y(n_2635)
);

NOR2xp67_ASAP7_75t_L g2636 ( 
.A(n_2574),
.B(n_2563),
.Y(n_2636)
);

XOR2x2_ASAP7_75t_L g2637 ( 
.A(n_2589),
.B(n_222),
.Y(n_2637)
);

NOR2x1_ASAP7_75t_L g2638 ( 
.A(n_2613),
.B(n_1301),
.Y(n_2638)
);

INVx2_ASAP7_75t_L g2639 ( 
.A(n_2563),
.Y(n_2639)
);

AOI22xp5_ASAP7_75t_L g2640 ( 
.A1(n_2562),
.A2(n_2614),
.B1(n_2546),
.B2(n_2545),
.Y(n_2640)
);

OAI221xp5_ASAP7_75t_L g2641 ( 
.A1(n_2555),
.A2(n_693),
.B1(n_704),
.B2(n_709),
.C(n_711),
.Y(n_2641)
);

OAI22xp5_ASAP7_75t_L g2642 ( 
.A1(n_2616),
.A2(n_730),
.B1(n_734),
.B2(n_719),
.Y(n_2642)
);

AOI322xp5_ASAP7_75t_L g2643 ( 
.A1(n_2548),
.A2(n_2085),
.A3(n_2089),
.B1(n_744),
.B2(n_775),
.C1(n_747),
.C2(n_772),
.Y(n_2643)
);

INVx1_ASAP7_75t_L g2644 ( 
.A(n_2600),
.Y(n_2644)
);

OAI22xp5_ASAP7_75t_L g2645 ( 
.A1(n_2543),
.A2(n_755),
.B1(n_758),
.B2(n_748),
.Y(n_2645)
);

BUFx3_ASAP7_75t_L g2646 ( 
.A(n_2556),
.Y(n_2646)
);

NAND3xp33_ASAP7_75t_SL g2647 ( 
.A(n_2552),
.B(n_759),
.C(n_1406),
.Y(n_2647)
);

AOI322xp5_ASAP7_75t_L g2648 ( 
.A1(n_2553),
.A2(n_2560),
.A3(n_2567),
.B1(n_2558),
.B2(n_2594),
.C1(n_2611),
.C2(n_2581),
.Y(n_2648)
);

INVx1_ASAP7_75t_L g2649 ( 
.A(n_2593),
.Y(n_2649)
);

AOI22xp5_ASAP7_75t_L g2650 ( 
.A1(n_2569),
.A2(n_2557),
.B1(n_2568),
.B2(n_2575),
.Y(n_2650)
);

AOI221xp5_ASAP7_75t_L g2651 ( 
.A1(n_2561),
.A2(n_1127),
.B1(n_1134),
.B2(n_1422),
.C(n_1301),
.Y(n_2651)
);

INVx1_ASAP7_75t_L g2652 ( 
.A(n_2593),
.Y(n_2652)
);

OAI22xp5_ASAP7_75t_L g2653 ( 
.A1(n_2573),
.A2(n_2006),
.B1(n_2056),
.B2(n_2041),
.Y(n_2653)
);

AOI322xp5_ASAP7_75t_L g2654 ( 
.A1(n_2583),
.A2(n_2085),
.A3(n_2076),
.B1(n_2053),
.B2(n_2066),
.C1(n_2007),
.C2(n_2090),
.Y(n_2654)
);

AOI22xp5_ASAP7_75t_L g2655 ( 
.A1(n_2572),
.A2(n_1275),
.B1(n_2041),
.B2(n_2006),
.Y(n_2655)
);

OAI211xp5_ASAP7_75t_SL g2656 ( 
.A1(n_2586),
.A2(n_2598),
.B(n_2584),
.C(n_2585),
.Y(n_2656)
);

AOI322xp5_ASAP7_75t_L g2657 ( 
.A1(n_2578),
.A2(n_2550),
.A3(n_2602),
.B1(n_2579),
.B2(n_2591),
.C1(n_2590),
.C2(n_2582),
.Y(n_2657)
);

INVx2_ASAP7_75t_L g2658 ( 
.A(n_2603),
.Y(n_2658)
);

AOI322xp5_ASAP7_75t_L g2659 ( 
.A1(n_2596),
.A2(n_2007),
.A3(n_2090),
.B1(n_1509),
.B2(n_1941),
.C1(n_2041),
.C2(n_2056),
.Y(n_2659)
);

NAND3xp33_ASAP7_75t_SL g2660 ( 
.A(n_2570),
.B(n_1407),
.C(n_1406),
.Y(n_2660)
);

XNOR2xp5_ASAP7_75t_L g2661 ( 
.A(n_2612),
.B(n_224),
.Y(n_2661)
);

INVx1_ASAP7_75t_L g2662 ( 
.A(n_2554),
.Y(n_2662)
);

AOI221xp5_ASAP7_75t_SL g2663 ( 
.A1(n_2588),
.A2(n_1127),
.B1(n_1134),
.B2(n_1401),
.C(n_1398),
.Y(n_2663)
);

AOI221xp5_ASAP7_75t_L g2664 ( 
.A1(n_2597),
.A2(n_1134),
.B1(n_1127),
.B2(n_1356),
.C(n_1331),
.Y(n_2664)
);

INVx2_ASAP7_75t_L g2665 ( 
.A(n_2604),
.Y(n_2665)
);

AOI221xp5_ASAP7_75t_SL g2666 ( 
.A1(n_2599),
.A2(n_1134),
.B1(n_1127),
.B2(n_1401),
.C(n_1407),
.Y(n_2666)
);

OAI211xp5_ASAP7_75t_SL g2667 ( 
.A1(n_2576),
.A2(n_1414),
.B(n_1304),
.C(n_1331),
.Y(n_2667)
);

OAI322xp33_ASAP7_75t_L g2668 ( 
.A1(n_2580),
.A2(n_1414),
.A3(n_1331),
.B1(n_1339),
.B2(n_1342),
.C1(n_1345),
.C2(n_1304),
.Y(n_2668)
);

AOI22xp5_ASAP7_75t_L g2669 ( 
.A1(n_2605),
.A2(n_1275),
.B1(n_2056),
.B2(n_2057),
.Y(n_2669)
);

AO22x2_ASAP7_75t_L g2670 ( 
.A1(n_2627),
.A2(n_2601),
.B1(n_2608),
.B2(n_2566),
.Y(n_2670)
);

OAI22xp5_ASAP7_75t_L g2671 ( 
.A1(n_2640),
.A2(n_2607),
.B1(n_2592),
.B2(n_2606),
.Y(n_2671)
);

AOI22xp5_ASAP7_75t_L g2672 ( 
.A1(n_2649),
.A2(n_1275),
.B1(n_2057),
.B2(n_2040),
.Y(n_2672)
);

INVx1_ASAP7_75t_L g2673 ( 
.A(n_2625),
.Y(n_2673)
);

AOI31xp33_ASAP7_75t_L g2674 ( 
.A1(n_2639),
.A2(n_1334),
.A3(n_1338),
.B(n_1340),
.Y(n_2674)
);

CKINVDCx20_ASAP7_75t_R g2675 ( 
.A(n_2650),
.Y(n_2675)
);

AO22x1_ASAP7_75t_L g2676 ( 
.A1(n_2652),
.A2(n_1194),
.B1(n_1246),
.B2(n_1235),
.Y(n_2676)
);

AOI22xp5_ASAP7_75t_L g2677 ( 
.A1(n_2626),
.A2(n_2057),
.B1(n_2040),
.B2(n_1530),
.Y(n_2677)
);

INVx1_ASAP7_75t_L g2678 ( 
.A(n_2646),
.Y(n_2678)
);

AOI22xp5_ASAP7_75t_L g2679 ( 
.A1(n_2644),
.A2(n_2040),
.B1(n_1530),
.B2(n_1304),
.Y(n_2679)
);

INVx1_ASAP7_75t_L g2680 ( 
.A(n_2636),
.Y(n_2680)
);

OAI22xp5_ASAP7_75t_L g2681 ( 
.A1(n_2621),
.A2(n_1530),
.B1(n_1941),
.B2(n_1233),
.Y(n_2681)
);

AOI22xp33_ASAP7_75t_L g2682 ( 
.A1(n_2656),
.A2(n_1233),
.B1(n_1171),
.B2(n_1194),
.Y(n_2682)
);

INVx1_ASAP7_75t_L g2683 ( 
.A(n_2665),
.Y(n_2683)
);

AOI22xp5_ASAP7_75t_L g2684 ( 
.A1(n_2658),
.A2(n_1530),
.B1(n_1356),
.B2(n_1342),
.Y(n_2684)
);

AO22x2_ASAP7_75t_L g2685 ( 
.A1(n_2662),
.A2(n_1356),
.B1(n_1345),
.B2(n_1342),
.Y(n_2685)
);

INVx1_ASAP7_75t_L g2686 ( 
.A(n_2661),
.Y(n_2686)
);

OAI22x1_ASAP7_75t_L g2687 ( 
.A1(n_2634),
.A2(n_1233),
.B1(n_1171),
.B2(n_1194),
.Y(n_2687)
);

OAI22x1_ASAP7_75t_L g2688 ( 
.A1(n_2638),
.A2(n_1233),
.B1(n_1171),
.B2(n_1194),
.Y(n_2688)
);

CKINVDCx20_ASAP7_75t_R g2689 ( 
.A(n_2637),
.Y(n_2689)
);

HB1xp67_ASAP7_75t_L g2690 ( 
.A(n_2635),
.Y(n_2690)
);

INVx1_ASAP7_75t_L g2691 ( 
.A(n_2629),
.Y(n_2691)
);

OAI22xp5_ASAP7_75t_L g2692 ( 
.A1(n_2620),
.A2(n_1530),
.B1(n_1246),
.B2(n_1225),
.Y(n_2692)
);

INVx2_ASAP7_75t_L g2693 ( 
.A(n_2628),
.Y(n_2693)
);

OAI22xp5_ASAP7_75t_L g2694 ( 
.A1(n_2619),
.A2(n_1217),
.B1(n_1235),
.B2(n_1231),
.Y(n_2694)
);

INVx1_ASAP7_75t_L g2695 ( 
.A(n_2633),
.Y(n_2695)
);

AOI22xp5_ASAP7_75t_L g2696 ( 
.A1(n_2623),
.A2(n_1345),
.B1(n_1339),
.B2(n_1308),
.Y(n_2696)
);

AO22x2_ASAP7_75t_L g2697 ( 
.A1(n_2642),
.A2(n_1308),
.B1(n_1339),
.B2(n_1338),
.Y(n_2697)
);

INVx1_ASAP7_75t_L g2698 ( 
.A(n_2647),
.Y(n_2698)
);

AOI22xp5_ASAP7_75t_L g2699 ( 
.A1(n_2664),
.A2(n_1308),
.B1(n_1373),
.B2(n_1354),
.Y(n_2699)
);

AO22x2_ASAP7_75t_L g2700 ( 
.A1(n_2645),
.A2(n_1340),
.B1(n_1334),
.B2(n_233),
.Y(n_2700)
);

AO22x2_ASAP7_75t_L g2701 ( 
.A1(n_2660),
.A2(n_229),
.B1(n_231),
.B2(n_234),
.Y(n_2701)
);

OA22x2_ASAP7_75t_L g2702 ( 
.A1(n_2657),
.A2(n_2655),
.B1(n_2648),
.B2(n_2653),
.Y(n_2702)
);

OAI22xp5_ASAP7_75t_L g2703 ( 
.A1(n_2641),
.A2(n_1246),
.B1(n_1235),
.B2(n_1231),
.Y(n_2703)
);

XOR2xp5_ASAP7_75t_L g2704 ( 
.A(n_2675),
.B(n_2666),
.Y(n_2704)
);

NOR3xp33_ASAP7_75t_L g2705 ( 
.A(n_2678),
.B(n_2624),
.C(n_2667),
.Y(n_2705)
);

NOR2x1p5_ASAP7_75t_L g2706 ( 
.A(n_2691),
.B(n_2663),
.Y(n_2706)
);

XNOR2xp5_ASAP7_75t_L g2707 ( 
.A(n_2689),
.B(n_2651),
.Y(n_2707)
);

NAND5xp2_ASAP7_75t_L g2708 ( 
.A(n_2680),
.B(n_2618),
.C(n_2622),
.D(n_2631),
.E(n_2630),
.Y(n_2708)
);

AOI32xp33_ASAP7_75t_L g2709 ( 
.A1(n_2683),
.A2(n_2668),
.A3(n_2632),
.B1(n_2659),
.B2(n_2669),
.Y(n_2709)
);

INVx1_ASAP7_75t_L g2710 ( 
.A(n_2690),
.Y(n_2710)
);

OAI322xp33_ASAP7_75t_L g2711 ( 
.A1(n_2673),
.A2(n_2654),
.A3(n_2643),
.B1(n_1379),
.B2(n_1405),
.C1(n_1387),
.C2(n_1389),
.Y(n_2711)
);

INVx4_ASAP7_75t_L g2712 ( 
.A(n_2702),
.Y(n_2712)
);

OAI22xp5_ASAP7_75t_L g2713 ( 
.A1(n_2670),
.A2(n_1246),
.B1(n_1171),
.B2(n_1196),
.Y(n_2713)
);

NAND5xp2_ASAP7_75t_L g2714 ( 
.A(n_2686),
.B(n_236),
.C(n_241),
.D(n_244),
.E(n_246),
.Y(n_2714)
);

NOR2xp33_ASAP7_75t_L g2715 ( 
.A(n_2695),
.B(n_247),
.Y(n_2715)
);

XNOR2xp5_ASAP7_75t_L g2716 ( 
.A(n_2670),
.B(n_260),
.Y(n_2716)
);

OAI22xp5_ASAP7_75t_L g2717 ( 
.A1(n_2698),
.A2(n_1225),
.B1(n_1196),
.B2(n_1201),
.Y(n_2717)
);

AND2x2_ASAP7_75t_L g2718 ( 
.A(n_2693),
.B(n_2063),
.Y(n_2718)
);

AOI221xp5_ASAP7_75t_L g2719 ( 
.A1(n_2671),
.A2(n_1401),
.B1(n_1235),
.B2(n_1217),
.C(n_1231),
.Y(n_2719)
);

NAND4xp25_ASAP7_75t_SL g2720 ( 
.A(n_2696),
.B(n_1983),
.C(n_270),
.D(n_274),
.Y(n_2720)
);

AOI21xp33_ASAP7_75t_L g2721 ( 
.A1(n_2687),
.A2(n_266),
.B(n_279),
.Y(n_2721)
);

NAND2xp5_ASAP7_75t_SL g2722 ( 
.A(n_2692),
.B(n_2681),
.Y(n_2722)
);

AOI211xp5_ASAP7_75t_L g2723 ( 
.A1(n_2703),
.A2(n_1401),
.B(n_1282),
.C(n_1290),
.Y(n_2723)
);

OAI222xp33_ASAP7_75t_L g2724 ( 
.A1(n_2699),
.A2(n_1217),
.B1(n_1196),
.B2(n_1225),
.C1(n_1231),
.C2(n_1201),
.Y(n_2724)
);

NAND2xp5_ASAP7_75t_L g2725 ( 
.A(n_2700),
.B(n_281),
.Y(n_2725)
);

OAI221xp5_ASAP7_75t_L g2726 ( 
.A1(n_2682),
.A2(n_1217),
.B1(n_1225),
.B2(n_1201),
.C(n_1196),
.Y(n_2726)
);

AOI22xp5_ASAP7_75t_L g2727 ( 
.A1(n_2697),
.A2(n_1354),
.B1(n_1373),
.B2(n_1403),
.Y(n_2727)
);

INVxp67_ASAP7_75t_L g2728 ( 
.A(n_2688),
.Y(n_2728)
);

NAND2xp5_ASAP7_75t_L g2729 ( 
.A(n_2710),
.B(n_2685),
.Y(n_2729)
);

NOR2xp33_ASAP7_75t_L g2730 ( 
.A(n_2712),
.B(n_2674),
.Y(n_2730)
);

AOI221xp5_ASAP7_75t_L g2731 ( 
.A1(n_2712),
.A2(n_2694),
.B1(n_2701),
.B2(n_2697),
.C(n_2676),
.Y(n_2731)
);

AOI21xp5_ASAP7_75t_L g2732 ( 
.A1(n_2704),
.A2(n_2684),
.B(n_2679),
.Y(n_2732)
);

INVx4_ASAP7_75t_L g2733 ( 
.A(n_2706),
.Y(n_2733)
);

INVx1_ASAP7_75t_L g2734 ( 
.A(n_2716),
.Y(n_2734)
);

OA22x2_ASAP7_75t_L g2735 ( 
.A1(n_2725),
.A2(n_2677),
.B1(n_2672),
.B2(n_1373),
.Y(n_2735)
);

OAI22xp33_ASAP7_75t_SL g2736 ( 
.A1(n_2728),
.A2(n_1201),
.B1(n_1379),
.B2(n_1387),
.Y(n_2736)
);

OAI21x1_ASAP7_75t_SL g2737 ( 
.A1(n_2707),
.A2(n_289),
.B(n_291),
.Y(n_2737)
);

AO22x2_ASAP7_75t_SL g2738 ( 
.A1(n_2705),
.A2(n_1359),
.B1(n_1360),
.B2(n_1361),
.Y(n_2738)
);

AOI22xp5_ASAP7_75t_L g2739 ( 
.A1(n_2718),
.A2(n_1389),
.B1(n_1405),
.B2(n_1397),
.Y(n_2739)
);

OAI21x1_ASAP7_75t_L g2740 ( 
.A1(n_2722),
.A2(n_1387),
.B(n_1379),
.Y(n_2740)
);

INVx2_ASAP7_75t_L g2741 ( 
.A(n_2715),
.Y(n_2741)
);

INVx2_ASAP7_75t_L g2742 ( 
.A(n_2727),
.Y(n_2742)
);

XNOR2xp5_ASAP7_75t_L g2743 ( 
.A(n_2723),
.B(n_292),
.Y(n_2743)
);

INVx3_ASAP7_75t_L g2744 ( 
.A(n_2708),
.Y(n_2744)
);

OAI22xp5_ASAP7_75t_L g2745 ( 
.A1(n_2709),
.A2(n_1403),
.B1(n_1405),
.B2(n_1392),
.Y(n_2745)
);

NAND2xp5_ASAP7_75t_L g2746 ( 
.A(n_2721),
.B(n_2713),
.Y(n_2746)
);

AOI22xp5_ASAP7_75t_L g2747 ( 
.A1(n_2720),
.A2(n_1389),
.B1(n_1397),
.B2(n_1392),
.Y(n_2747)
);

INVx1_ASAP7_75t_L g2748 ( 
.A(n_2711),
.Y(n_2748)
);

INVx1_ASAP7_75t_L g2749 ( 
.A(n_2744),
.Y(n_2749)
);

OAI22xp5_ASAP7_75t_L g2750 ( 
.A1(n_2733),
.A2(n_2726),
.B1(n_2717),
.B2(n_2719),
.Y(n_2750)
);

AOI22xp5_ASAP7_75t_L g2751 ( 
.A1(n_2730),
.A2(n_2714),
.B1(n_2724),
.B2(n_1392),
.Y(n_2751)
);

AOI22xp33_ASAP7_75t_L g2752 ( 
.A1(n_2741),
.A2(n_1309),
.B1(n_1346),
.B2(n_1343),
.Y(n_2752)
);

OR2x2_ASAP7_75t_L g2753 ( 
.A(n_2734),
.B(n_293),
.Y(n_2753)
);

AOI21xp5_ASAP7_75t_L g2754 ( 
.A1(n_2729),
.A2(n_1105),
.B(n_1098),
.Y(n_2754)
);

AOI22x1_ASAP7_75t_L g2755 ( 
.A1(n_2748),
.A2(n_1403),
.B1(n_1397),
.B2(n_1419),
.Y(n_2755)
);

AOI222xp33_ASAP7_75t_L g2756 ( 
.A1(n_2731),
.A2(n_1309),
.B1(n_1328),
.B2(n_1279),
.C1(n_1282),
.C2(n_1290),
.Y(n_2756)
);

XNOR2x1_ASAP7_75t_L g2757 ( 
.A(n_2746),
.B(n_296),
.Y(n_2757)
);

INVx3_ASAP7_75t_L g2758 ( 
.A(n_2742),
.Y(n_2758)
);

AOI22xp33_ASAP7_75t_L g2759 ( 
.A1(n_2737),
.A2(n_1282),
.B1(n_1309),
.B2(n_1328),
.Y(n_2759)
);

BUFx2_ASAP7_75t_L g2760 ( 
.A(n_2749),
.Y(n_2760)
);

AOI21xp5_ASAP7_75t_L g2761 ( 
.A1(n_2758),
.A2(n_2732),
.B(n_2745),
.Y(n_2761)
);

NAND2xp5_ASAP7_75t_L g2762 ( 
.A(n_2751),
.B(n_2743),
.Y(n_2762)
);

NAND2x1p5_ASAP7_75t_L g2763 ( 
.A(n_2753),
.B(n_2757),
.Y(n_2763)
);

INVx1_ASAP7_75t_L g2764 ( 
.A(n_2755),
.Y(n_2764)
);

INVx1_ASAP7_75t_L g2765 ( 
.A(n_2750),
.Y(n_2765)
);

OAI21xp5_ASAP7_75t_L g2766 ( 
.A1(n_2754),
.A2(n_2735),
.B(n_2747),
.Y(n_2766)
);

AOI21xp5_ASAP7_75t_L g2767 ( 
.A1(n_2760),
.A2(n_2736),
.B(n_2738),
.Y(n_2767)
);

AOI22xp5_ASAP7_75t_SL g2768 ( 
.A1(n_2765),
.A2(n_2759),
.B1(n_2740),
.B2(n_2739),
.Y(n_2768)
);

NAND2xp5_ASAP7_75t_L g2769 ( 
.A(n_2763),
.B(n_2756),
.Y(n_2769)
);

AOI21xp5_ASAP7_75t_L g2770 ( 
.A1(n_2762),
.A2(n_2752),
.B(n_1105),
.Y(n_2770)
);

NAND2xp5_ASAP7_75t_L g2771 ( 
.A(n_2761),
.B(n_300),
.Y(n_2771)
);

OA22x2_ASAP7_75t_L g2772 ( 
.A1(n_2766),
.A2(n_307),
.B1(n_308),
.B2(n_311),
.Y(n_2772)
);

INVx1_ASAP7_75t_L g2773 ( 
.A(n_2764),
.Y(n_2773)
);

AOI22xp33_ASAP7_75t_L g2774 ( 
.A1(n_2760),
.A2(n_1279),
.B1(n_1282),
.B2(n_1290),
.Y(n_2774)
);

OAI22xp33_ASAP7_75t_L g2775 ( 
.A1(n_2773),
.A2(n_1309),
.B1(n_1282),
.B2(n_1290),
.Y(n_2775)
);

OAI22xp5_ASAP7_75t_SL g2776 ( 
.A1(n_2769),
.A2(n_1098),
.B1(n_1115),
.B2(n_1125),
.Y(n_2776)
);

AOI22xp33_ASAP7_75t_L g2777 ( 
.A1(n_2772),
.A2(n_1290),
.B1(n_1309),
.B2(n_1316),
.Y(n_2777)
);

OAI22xp33_ASAP7_75t_L g2778 ( 
.A1(n_2771),
.A2(n_1316),
.B1(n_1328),
.B2(n_1346),
.Y(n_2778)
);

AOI22xp5_ASAP7_75t_L g2779 ( 
.A1(n_2767),
.A2(n_1328),
.B1(n_1316),
.B2(n_1343),
.Y(n_2779)
);

AOI22xp5_ASAP7_75t_L g2780 ( 
.A1(n_2770),
.A2(n_2774),
.B1(n_2768),
.B2(n_1346),
.Y(n_2780)
);

NAND3xp33_ASAP7_75t_L g2781 ( 
.A(n_2780),
.B(n_1098),
.C(n_1105),
.Y(n_2781)
);

AOI21xp5_ASAP7_75t_L g2782 ( 
.A1(n_2776),
.A2(n_1098),
.B(n_1126),
.Y(n_2782)
);

OA21x2_ASAP7_75t_L g2783 ( 
.A1(n_2777),
.A2(n_1366),
.B(n_1361),
.Y(n_2783)
);

NAND2xp5_ASAP7_75t_SL g2784 ( 
.A(n_2778),
.B(n_1105),
.Y(n_2784)
);

AOI21xp5_ASAP7_75t_L g2785 ( 
.A1(n_2775),
.A2(n_1115),
.B(n_1126),
.Y(n_2785)
);

OAI21xp5_ASAP7_75t_SL g2786 ( 
.A1(n_2779),
.A2(n_1346),
.B(n_1343),
.Y(n_2786)
);

OAI21xp5_ASAP7_75t_L g2787 ( 
.A1(n_2780),
.A2(n_1419),
.B(n_1129),
.Y(n_2787)
);

AO21x2_ASAP7_75t_L g2788 ( 
.A1(n_2787),
.A2(n_1366),
.B(n_1360),
.Y(n_2788)
);

OAI211xp5_ASAP7_75t_SL g2789 ( 
.A1(n_2784),
.A2(n_1359),
.B(n_317),
.C(n_319),
.Y(n_2789)
);

AOI221xp5_ASAP7_75t_L g2790 ( 
.A1(n_2789),
.A2(n_2782),
.B1(n_2781),
.B2(n_2785),
.C(n_2786),
.Y(n_2790)
);

AOI221xp5_ASAP7_75t_L g2791 ( 
.A1(n_2788),
.A2(n_2783),
.B1(n_1316),
.B2(n_1346),
.C(n_1343),
.Y(n_2791)
);

OA21x2_ASAP7_75t_L g2792 ( 
.A1(n_2790),
.A2(n_312),
.B(n_321),
.Y(n_2792)
);

OAI31xp33_ASAP7_75t_L g2793 ( 
.A1(n_2792),
.A2(n_2791),
.A3(n_328),
.B(n_329),
.Y(n_2793)
);


endmodule